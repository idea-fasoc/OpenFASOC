* NGSPICE file created from opamp_sample_0003.ext - technology: sky130A

.subckt opamp_sample_0003 GND VOUT VDD VN VP CS_BIAS DIFFPAIR_BIAS
X0 GND.t194 CS_BIAS.t2 CS_BIAS.t3 GND.t162 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=2
X1 VDD.t190 a_n8209_7799.t20 VOUT.t40 VDD.t97 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=1
X2 VDD.t189 a_n8209_7799.t21 VOUT.t39 VDD.t108 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=1
X3 VOUT.t112 a_n2686_8222.t8 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X4 VDD.t77 VDD.t75 VDD.t76 VDD.t50 sky130_fd_pr__pfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=1
X5 a_n2511_10356.t19 a_n2686_12578.t17 a_n2686_12578.t18 VDD.t90 sky130_fd_pr__pfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=1
X6 GND.t91 GND.t89 GND.t90 GND.t39 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=2
X7 a_n2686_12578.t6 a_n2686_12578.t5 a_n2511_10356.t18 VDD.t83 sky130_fd_pr__pfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=1
X8 VDD.t94 a_n2686_12578.t32 a_n2686_8222.t7 VDD.t93 sky130_fd_pr__pfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=1
X9 GND.t88 GND.t86 GND.t87 GND.t25 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=2
X10 GND.t193 CS_BIAS.t0 CS_BIAS.t1 GND.t132 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=2
X11 GND.t192 CS_BIAS.t40 VOUT.t111 GND.t134 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=2
X12 a_n8209_7799.t1 VN.t5 a_n1455_n3628.t7 GND.t95 sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=1
X13 VDD.t188 a_n8209_7799.t22 VOUT.t69 VDD.t105 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=1
X14 VOUT.t68 a_n8209_7799.t23 VDD.t187 VDD.t172 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=1
X15 a_n2686_12578.t10 a_n2686_12578.t9 a_n2511_10356.t17 VDD.t197 sky130_fd_pr__pfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=1
X16 CS_BIAS.t19 CS_BIAS.t18 GND.t191 GND.t136 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=2
X17 VOUT.t67 a_n8209_7799.t24 VDD.t186 VDD.t103 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=1
X18 VOUT.t113 a_n2686_8222.t8 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X19 a_n8209_7799.t2 a_n2686_12578.t33 a_n2686_8222.t2 VDD.t79 sky130_fd_pr__pfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=1
X20 VOUT.t38 a_n8209_7799.t25 VDD.t185 VDD.t152 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=1
X21 VOUT.t37 a_n8209_7799.t26 VDD.t184 VDD.t157 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=1
X22 GND.t190 CS_BIAS.t16 CS_BIAS.t17 GND.t156 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=2
X23 a_n2686_8222.t15 a_n2686_12578.t34 a_n8209_7799.t12 VDD.t197 sky130_fd_pr__pfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=1
X24 VDD.t183 a_n8209_7799.t27 VOUT.t36 VDD.t99 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=1
X25 VDD.t182 a_n8209_7799.t28 VOUT.t26 VDD.t139 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=1
X26 VOUT.t110 CS_BIAS.t41 GND.t189 GND.t143 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=2
X27 a_n2686_12578.t29 VP.t5 a_n1455_n3628.t17 GND.t100 sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=1
X28 VOUT.t25 a_n8209_7799.t29 VDD.t181 VDD.t95 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=1
X29 a_n1455_n3628.t14 DIFFPAIR_BIAS.t8 GND.t110 GND.t109 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X30 a_n1455_n3628.t10 VP.t6 a_n2686_12578.t26 GND.t98 sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=1
X31 VOUT.t24 a_n8209_7799.t30 VDD.t180 VDD.t172 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=1
X32 GND.t188 CS_BIAS.t42 VOUT.t109 GND.t151 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=2
X33 GND.t187 CS_BIAS.t43 VOUT.t108 GND.t162 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=2
X34 VDD.t199 a_n2686_12578.t35 a_n2686_8222.t9 VDD.t198 sky130_fd_pr__pfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=1
X35 DIFFPAIR_BIAS.t7 DIFFPAIR_BIAS.t6 GND.t112 GND.t111 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X36 VDD.t74 VDD.t72 VDD.t73 VDD.t30 sky130_fd_pr__pfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=1
X37 VDD.t179 a_n8209_7799.t31 VOUT.t9 VDD.t97 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=1
X38 a_n2511_10356.t16 a_n2686_12578.t21 a_n2686_12578.t22 VDD.t92 sky130_fd_pr__pfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=1
X39 VN.t4 GND.t83 GND.t85 GND.t84 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X40 GND.t82 GND.t79 GND.t81 GND.t80 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=2
X41 a_n2686_8222.t5 a_n2686_12578.t36 VDD.t89 VDD.t88 sky130_fd_pr__pfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=1
X42 GND.t78 GND.t76 GND.t77 GND.t39 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=2
X43 GND.t186 CS_BIAS.t44 VOUT.t107 GND.t148 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=2
X44 GND.t75 GND.t73 VP.t4 GND.t74 sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.5
X45 GND.t72 GND.t69 GND.t71 GND.t70 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=2
X46 VOUT.t8 a_n8209_7799.t32 VDD.t178 VDD.t162 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=1
X47 a_n2511_10356.t7 a_n2686_12578.t37 VDD.t81 VDD.t80 sky130_fd_pr__pfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=1
X48 VDD.t177 a_n8209_7799.t33 VOUT.t7 VDD.t147 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=1
X49 VOUT.t106 CS_BIAS.t45 GND.t184 GND.t115 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=2
X50 VOUT.t105 CS_BIAS.t46 GND.t183 GND.t159 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=2
X51 VDD.t176 a_n8209_7799.t34 VOUT.t59 VDD.t101 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=1
X52 GND.t185 CS_BIAS.t14 CS_BIAS.t15 GND.t148 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=2
X53 a_n2511_10356.t6 a_n2686_12578.t38 VDD.t213 VDD.t212 sky130_fd_pr__pfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=1
X54 DIFFPAIR_BIAS.t5 DIFFPAIR_BIAS.t4 GND.t114 GND.t113 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X55 CS_BIAS.t39 CS_BIAS.t38 GND.t182 GND.t123 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=2
X56 a_n8209_7799.t17 a_n2686_12578.t39 a_n2686_8222.t18 VDD.t92 sky130_fd_pr__pfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=1
X57 VOUT.t58 a_n8209_7799.t35 VDD.t175 VDD.t119 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=1
X58 a_n1455_n3628.t15 VP.t7 a_n2686_12578.t27 GND.t99 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=1
X59 VOUT.t57 a_n8209_7799.t36 VDD.t174 VDD.t152 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=1
X60 VDD.t71 VDD.t69 VDD.t70 VDD.t3 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=1
X61 GND.t68 GND.t66 VP.t3 GND.t67 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.5
X62 a_n1455_n3628.t13 DIFFPAIR_BIAS.t9 GND.t108 GND.t107 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X63 GND.t181 CS_BIAS.t47 VOUT.t104 GND.t156 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=2
X64 GND.t180 CS_BIAS.t48 VOUT.t103 GND.t154 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=2
X65 VOUT.t30 a_n8209_7799.t37 VDD.t173 VDD.t172 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=1
X66 a_n2686_12578.t20 a_n2686_12578.t19 a_n2511_10356.t15 VDD.t210 sky130_fd_pr__pfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=1
X67 a_n8209_7799.t3 VN.t6 a_n1455_n3628.t6 GND.t96 sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=1
X68 VOUT.t29 a_n8209_7799.t38 VDD.t171 VDD.t113 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=1
X69 VDD.t170 a_n8209_7799.t39 VOUT.t52 VDD.t155 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=1
X70 VDD.t68 VDD.t66 VDD.t67 VDD.t60 sky130_fd_pr__pfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=1
X71 VDD.t87 a_n2686_12578.t40 a_n2511_10356.t5 VDD.t86 sky130_fd_pr__pfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=1
X72 VN.t3 GND.t63 GND.t65 GND.t64 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X73 CS_BIAS.t37 CS_BIAS.t36 GND.t179 GND.t121 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=2
X74 VOUT.t51 a_n8209_7799.t40 VDD.t169 VDD.t157 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=1
X75 VOUT.t50 a_n8209_7799.t41 VDD.t168 VDD.t162 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=1
X76 VDD.t167 a_n8209_7799.t42 VOUT.t33 VDD.t101 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=1
X77 a_n2511_10356.t4 a_n2686_12578.t41 VDD.t85 VDD.t84 sky130_fd_pr__pfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=1
X78 VOUT.t32 a_n8209_7799.t43 VDD.t166 VDD.t95 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=1
X79 VDD.t165 a_n8209_7799.t44 VOUT.t31 VDD.t108 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=1
X80 GND.t62 GND.t60 GND.t61 GND.t29 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=1
X81 GND.t178 CS_BIAS.t49 VOUT.t102 GND.t119 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=2
X82 VOUT.t114 a_n2686_8222.t8 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X83 a_n1455_n3628.t5 VN.t7 a_n8209_7799.t15 GND.t97 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=1
X84 VDD.t164 a_n8209_7799.t45 VOUT.t35 VDD.t99 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=1
X85 GND.t59 GND.t57 GND.t58 GND.t25 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=2
X86 VDD.t65 VDD.t63 VDD.t64 VDD.t7 sky130_fd_pr__pfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=1
X87 VOUT.t34 a_n8209_7799.t46 VDD.t163 VDD.t162 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=1
X88 VDD.t161 a_n8209_7799.t47 VOUT.t43 VDD.t155 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=1
X89 VOUT.t101 CS_BIAS.t50 GND.t177 GND.t136 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=2
X90 VDD.t160 a_n8209_7799.t48 VOUT.t42 VDD.t147 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=1
X91 a_n2511_10356.t14 a_n2686_12578.t23 a_n2686_12578.t24 VDD.t211 sky130_fd_pr__pfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=1
X92 VOUT.t41 a_n8209_7799.t49 VDD.t159 VDD.t131 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=1
X93 VOUT.t54 a_n8209_7799.t50 VDD.t158 VDD.t157 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=1
X94 VDD.t156 a_n8209_7799.t51 VOUT.t53 VDD.t155 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=1
X95 VDD.t62 VDD.t59 VDD.t61 VDD.t60 sky130_fd_pr__pfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=1
X96 GND.t176 CS_BIAS.t51 VOUT.t100 GND.t129 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=2
X97 CS_BIAS.t7 CS_BIAS.t6 GND.t175 GND.t159 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=2
X98 GND.t53 GND.t51 GND.t52 GND.t12 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=2
X99 VDD.t154 a_n8209_7799.t52 VOUT.t61 VDD.t143 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=1
X100 VOUT.t60 a_n8209_7799.t53 VDD.t153 VDD.t152 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=1
X101 VOUT.t99 CS_BIAS.t52 GND.t174 GND.t141 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=2
X102 VDD.t58 VDD.t56 VDD.t57 VDD.t14 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=1
X103 a_n2511_10356.t13 a_n2686_12578.t1 a_n2686_12578.t2 VDD.t79 sky130_fd_pr__pfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=1
X104 VOUT.t98 CS_BIAS.t53 GND.t173 GND.t121 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=2
X105 VDD.t151 a_n8209_7799.t54 VOUT.t2 VDD.t139 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=1
X106 a_n2686_8222.t17 a_n2686_12578.t42 a_n8209_7799.t13 VDD.t210 sky130_fd_pr__pfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=1
X107 VDD.t150 a_n8209_7799.t55 VOUT.t1 VDD.t143 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=1
X108 GND.t56 GND.t54 VN.t2 GND.t55 sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.5
X109 VOUT.t97 CS_BIAS.t54 GND.t172 GND.t117 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=2
X110 a_n8209_7799.t4 VN.t8 a_n1455_n3628.t4 GND.t92 sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=1
X111 VDD.t55 VDD.t53 VDD.t54 VDD.t26 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=1
X112 VP.t2 GND.t48 GND.t50 GND.t49 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X113 GND.t167 CS_BIAS.t55 VOUT.t96 GND.t127 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=2
X114 VOUT.t0 a_n8209_7799.t56 VDD.t149 VDD.t127 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=1
X115 a_n2686_12578.t14 a_n2686_12578.t13 a_n2511_10356.t12 VDD.t91 sky130_fd_pr__pfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=1
X116 VDD.t148 a_n8209_7799.t57 VOUT.t21 VDD.t147 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=1
X117 VDD.t146 a_n8209_7799.t58 VOUT.t20 VDD.t122 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=1
X118 GND.t171 CS_BIAS.t4 CS_BIAS.t5 GND.t127 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=2
X119 VOUT.t95 CS_BIAS.t56 GND.t170 GND.t125 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=2
X120 GND.t169 CS_BIAS.t57 VOUT.t94 GND.t134 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=2
X121 VOUT.t45 a_n8209_7799.t59 VDD.t145 VDD.t131 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=1
X122 DIFFPAIR_BIAS.t3 DIFFPAIR_BIAS.t2 GND.t102 GND.t101 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X123 VOUT.t93 CS_BIAS.t58 GND.t168 GND.t138 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=2
X124 VOUT.t92 CS_BIAS.t59 GND.t166 GND.t123 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=2
X125 VDD.t52 VDD.t49 VDD.t51 VDD.t50 sky130_fd_pr__pfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=1
X126 VDD.t48 VDD.t45 VDD.t47 VDD.t46 sky130_fd_pr__pfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=1
X127 a_n2686_8222.t0 a_n2686_12578.t43 VDD.t1 VDD.t0 sky130_fd_pr__pfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=1
X128 VDD.t144 a_n8209_7799.t60 VOUT.t44 VDD.t143 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=1
X129 VDD.t44 VDD.t42 VDD.t43 VDD.t14 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=1
X130 VDD.t142 a_n8209_7799.t61 VOUT.t19 VDD.t115 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=1
X131 VOUT.t18 a_n8209_7799.t62 VDD.t141 VDD.t124 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=1
X132 GND.t10 GND.t7 GND.t9 GND.t8 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=1
X133 VDD.t140 a_n8209_7799.t63 VOUT.t17 VDD.t139 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=1
X134 VOUT.t115 a_n2686_8222.t8 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X135 GND.t165 CS_BIAS.t60 VOUT.t91 GND.t132 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=2
X136 VOUT.t56 a_n8209_7799.t64 VDD.t138 VDD.t127 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=1
X137 CS_BIAS.t23 CS_BIAS.t22 GND.t164 GND.t141 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=2
X138 GND.t163 CS_BIAS.t61 VOUT.t90 GND.t162 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=2
X139 a_n2686_8222.t13 a_n2686_12578.t44 VDD.t203 VDD.t202 sky130_fd_pr__pfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=1
X140 a_n1455_n3628.t19 VP.t8 a_n2686_12578.t31 GND.t195 sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=1
X141 GND.t47 GND.t45 VN.t1 GND.t46 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X142 GND.t44 GND.t42 GND.t43 GND.t1 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=2
X143 a_n1455_n3628.t12 DIFFPAIR_BIAS.t10 GND.t106 GND.t105 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X144 GND.t161 CS_BIAS.t20 CS_BIAS.t21 GND.t154 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=2
X145 VOUT.t89 CS_BIAS.t62 GND.t160 GND.t159 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=2
X146 a_n2686_12578.t16 a_n2686_12578.t15 a_n2511_10356.t11 VDD.t191 sky130_fd_pr__pfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=1
X147 GND.t41 GND.t38 GND.t40 GND.t39 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=2
X148 a_n2686_12578.t12 a_n2686_12578.t11 a_n2511_10356.t10 VDD.t82 sky130_fd_pr__pfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=1
X149 VDD.t41 VDD.t39 VDD.t40 VDD.t18 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=1
X150 VOUT.t55 a_n8209_7799.t65 VDD.t137 VDD.t103 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=1
X151 VDD.t38 VDD.t36 VDD.t37 VDD.t26 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=1
X152 VDD.t136 a_n8209_7799.t66 VOUT.t64 VDD.t117 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=1
X153 a_n2686_12578.t30 VP.t9 a_n1455_n3628.t18 GND.t95 sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=1
X154 a_n1455_n3628.t3 VN.t9 a_n8209_7799.t8 GND.t99 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=1
X155 VOUT.t63 a_n8209_7799.t67 VDD.t135 VDD.t124 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=1
X156 GND.t158 CS_BIAS.t28 CS_BIAS.t29 GND.t151 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=2
X157 VDD.t134 a_n8209_7799.t68 VOUT.t62 VDD.t122 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=1
X158 a_n2686_8222.t19 a_n2686_12578.t45 a_n8209_7799.t18 VDD.t191 sky130_fd_pr__pfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=1
X159 GND.t157 CS_BIAS.t63 VOUT.t88 GND.t156 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=2
X160 GND.t155 CS_BIAS.t64 VOUT.t87 GND.t154 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=2
X161 a_n2686_8222.t10 a_n2686_12578.t46 VDD.t201 VDD.t200 sky130_fd_pr__pfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=1
X162 VOUT.t86 CS_BIAS.t65 GND.t153 GND.t143 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=2
X163 a_n2686_12578.t28 VP.t10 a_n1455_n3628.t16 GND.t96 sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=1
X164 a_n8209_7799.t9 VN.t10 a_n1455_n3628.t2 GND.t100 sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=1
X165 VOUT.t28 a_n8209_7799.t69 VDD.t133 VDD.t119 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=1
X166 GND.t37 GND.t35 GND.t36 GND.t1 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=2
X167 a_n1455_n3628.t1 VN.t11 a_n8209_7799.t14 GND.t98 sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=1
X168 GND.t152 CS_BIAS.t66 VOUT.t85 GND.t151 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=2
X169 VDD.t35 VDD.t33 VDD.t34 VDD.t18 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=1
X170 CS_BIAS.t27 CS_BIAS.t26 GND.t150 GND.t138 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=2
X171 GND.t34 GND.t32 GND.t33 GND.t12 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=2
X172 a_n2511_10356.t9 a_n2686_12578.t7 a_n2686_12578.t8 VDD.t78 sky130_fd_pr__pfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=1
X173 a_n8209_7799.t11 a_n2686_12578.t47 a_n2686_8222.t12 VDD.t192 sky130_fd_pr__pfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=1
X174 VDD.t32 VDD.t29 VDD.t31 VDD.t30 sky130_fd_pr__pfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=1
X175 VOUT.t27 a_n8209_7799.t70 VDD.t132 VDD.t131 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=1
X176 GND.t149 CS_BIAS.t67 VOUT.t84 GND.t148 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=2
X177 VDD.t28 VDD.t25 VDD.t27 VDD.t26 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=1
X178 GND.t31 GND.t28 GND.t30 GND.t29 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=1
X179 VDD.t130 a_n8209_7799.t71 VOUT.t12 VDD.t115 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=1
X180 VDD.t129 a_n8209_7799.t72 VOUT.t11 VDD.t117 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=1
X181 VOUT.t83 CS_BIAS.t68 GND.t147 GND.t115 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=2
X182 VOUT.t116 a_n2686_8222.t8 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X183 a_n1455_n3628.t9 VP.t11 a_n2686_12578.t25 GND.t97 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=1
X184 VOUT.t10 a_n8209_7799.t73 VDD.t128 VDD.t127 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=1
X185 CS_BIAS.t13 CS_BIAS.t12 GND.t146 GND.t125 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=2
X186 VOUT.t4 a_n8209_7799.t74 VDD.t126 VDD.t113 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=1
X187 VOUT.t3 a_n8209_7799.t75 VDD.t125 VDD.t124 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=1
X188 a_n1455_n3628.t11 DIFFPAIR_BIAS.t11 GND.t104 GND.t103 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X189 VDD.t123 a_n8209_7799.t76 VOUT.t14 VDD.t122 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=1
X190 GND.t145 CS_BIAS.t10 CS_BIAS.t11 GND.t119 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=2
X191 GND.t27 GND.t24 GND.t26 GND.t25 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=2
X192 a_n8209_7799.t10 a_n2686_12578.t48 a_n2686_8222.t11 VDD.t90 sky130_fd_pr__pfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=1
X193 VDD.t24 VDD.t21 VDD.t23 VDD.t22 sky130_fd_pr__pfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=1
X194 VOUT.t13 a_n8209_7799.t77 VDD.t121 VDD.t110 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=1
X195 VOUT.t23 a_n8209_7799.t78 VDD.t120 VDD.t119 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=1
X196 VDD.t215 a_n2686_12578.t49 a_n2511_10356.t3 VDD.t214 sky130_fd_pr__pfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=1
X197 VDD.t20 VDD.t17 VDD.t19 VDD.t18 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=1
X198 a_n2686_8222.t3 a_n2686_12578.t50 a_n8209_7799.t5 VDD.t83 sky130_fd_pr__pfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=1
X199 a_n2511_10356.t8 a_n2686_12578.t3 a_n2686_12578.t4 VDD.t192 sky130_fd_pr__pfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=1
X200 VDD.t118 a_n8209_7799.t79 VOUT.t22 VDD.t117 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=1
X201 CS_BIAS.t9 CS_BIAS.t8 GND.t144 GND.t143 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=2
X202 VDD.t194 a_n2686_12578.t51 a_n2511_10356.t2 VDD.t193 sky130_fd_pr__pfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=1
X203 VDD.t207 a_n2686_12578.t52 a_n2686_8222.t16 VDD.t206 sky130_fd_pr__pfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=1
X204 VDD.t116 a_n8209_7799.t80 VOUT.t49 VDD.t115 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=1
X205 a_n8209_7799.t19 a_n2686_12578.t53 a_n2686_8222.t20 VDD.t211 sky130_fd_pr__pfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=1
X206 VP.t1 GND.t21 GND.t23 GND.t22 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X207 VOUT.t82 CS_BIAS.t69 GND.t142 GND.t141 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=2
X208 DIFFPAIR_BIAS.t1 DIFFPAIR_BIAS.t0 GND.t94 GND.t93 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X209 VOUT.t48 a_n8209_7799.t81 VDD.t114 VDD.t113 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=1
X210 VDD.t16 VDD.t13 VDD.t15 VDD.t14 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=1
X211 GND.t120 CS_BIAS.t70 VOUT.t81 GND.t119 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=2
X212 VOUT.t80 CS_BIAS.t71 GND.t118 GND.t117 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=2
X213 GND.t128 CS_BIAS.t72 VOUT.t79 GND.t127 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=2
X214 VDD.t12 VDD.t10 VDD.t11 VDD.t3 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=1
X215 VOUT.t71 a_n8209_7799.t82 VDD.t112 VDD.t110 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=1
X216 a_n2686_8222.t6 a_n2686_12578.t54 a_n8209_7799.t7 VDD.t91 sky130_fd_pr__pfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=1
X217 VOUT.t78 CS_BIAS.t73 GND.t126 GND.t125 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=2
X218 GND.t140 CS_BIAS.t34 CS_BIAS.t35 GND.t129 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=2
X219 VDD.t205 a_n2686_12578.t55 a_n2686_8222.t14 VDD.t204 sky130_fd_pr__pfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=1
X220 VOUT.t70 a_n8209_7799.t83 VDD.t111 VDD.t110 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=1
X221 VDD.t109 a_n8209_7799.t84 VOUT.t47 VDD.t108 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=1
X222 a_n2686_8222.t4 a_n2686_12578.t56 a_n8209_7799.t6 VDD.t82 sky130_fd_pr__pfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=1
X223 VOUT.t77 CS_BIAS.t74 GND.t124 GND.t123 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=2
X224 VOUT.t76 CS_BIAS.t75 GND.t139 GND.t138 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=2
X225 VOUT.t75 CS_BIAS.t76 GND.t137 GND.t136 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=2
X226 VDD.t196 a_n2686_12578.t57 a_n2511_10356.t1 VDD.t195 sky130_fd_pr__pfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=1
X227 a_n2511_10356.t0 a_n2686_12578.t58 VDD.t209 VDD.t208 sky130_fd_pr__pfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=1
X228 VDD.t9 VDD.t6 VDD.t8 VDD.t7 sky130_fd_pr__pfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=1
X229 GND.t130 CS_BIAS.t77 VOUT.t74 GND.t129 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=2
X230 VDD.t107 a_n8209_7799.t85 VOUT.t46 VDD.t105 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=1
X231 GND.t20 GND.t18 GND.t19 GND.t8 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=1
X232 VDD.t106 a_n8209_7799.t86 VOUT.t66 VDD.t105 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=1
X233 GND.t17 GND.t15 VN.t0 GND.t16 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.5
X234 VOUT.t117 a_n2686_8222.t8 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X235 GND.t135 CS_BIAS.t32 CS_BIAS.t33 GND.t134 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=2
X236 GND.t14 GND.t11 GND.t13 GND.t12 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=2
X237 VOUT.t65 a_n8209_7799.t87 VDD.t104 VDD.t103 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=1
X238 GND.t133 CS_BIAS.t78 VOUT.t73 GND.t132 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=2
X239 a_n8209_7799.t0 a_n2686_12578.t59 a_n2686_8222.t1 VDD.t78 sky130_fd_pr__pfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=1
X240 VDD.t102 a_n8209_7799.t88 VOUT.t6 VDD.t101 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=1
X241 CS_BIAS.t31 CS_BIAS.t30 GND.t131 GND.t117 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=2
X242 a_n1455_n3628.t0 VN.t12 a_n8209_7799.t16 GND.t195 sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=1
X243 VOUT.t72 CS_BIAS.t79 GND.t122 GND.t121 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=2
X244 VDD.t100 a_n8209_7799.t89 VOUT.t5 VDD.t99 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=1
X245 VDD.t98 a_n8209_7799.t90 VOUT.t16 VDD.t97 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=1
X246 a_n2686_12578.t0 VP.t12 a_n1455_n3628.t8 GND.t92 sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=1
X247 VOUT.t15 a_n8209_7799.t91 VDD.t96 VDD.t95 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=1
X248 VDD.t5 VDD.t2 VDD.t4 VDD.t3 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=1
X249 CS_BIAS.t25 CS_BIAS.t24 GND.t116 GND.t115 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=2
X250 GND.t6 GND.t4 VP.t0 GND.t5 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X251 GND.t3 GND.t0 GND.t2 GND.t1 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=2
R0 CS_BIAS.n261 CS_BIAS.n179 161.3
R1 CS_BIAS.n260 CS_BIAS.n259 161.3
R2 CS_BIAS.n258 CS_BIAS.n180 161.3
R3 CS_BIAS.n257 CS_BIAS.n256 161.3
R4 CS_BIAS.n254 CS_BIAS.n181 161.3
R5 CS_BIAS.n253 CS_BIAS.n252 161.3
R6 CS_BIAS.n251 CS_BIAS.n182 161.3
R7 CS_BIAS.n250 CS_BIAS.n249 161.3
R8 CS_BIAS.n248 CS_BIAS.n183 161.3
R9 CS_BIAS.n246 CS_BIAS.n245 161.3
R10 CS_BIAS.n244 CS_BIAS.n184 161.3
R11 CS_BIAS.n243 CS_BIAS.n242 161.3
R12 CS_BIAS.n241 CS_BIAS.n185 161.3
R13 CS_BIAS.n240 CS_BIAS.n239 161.3
R14 CS_BIAS.n238 CS_BIAS.n237 161.3
R15 CS_BIAS.n236 CS_BIAS.n187 161.3
R16 CS_BIAS.n235 CS_BIAS.n234 161.3
R17 CS_BIAS.n233 CS_BIAS.n188 161.3
R18 CS_BIAS.n232 CS_BIAS.n231 161.3
R19 CS_BIAS.n230 CS_BIAS.n189 161.3
R20 CS_BIAS.n229 CS_BIAS.n228 161.3
R21 CS_BIAS.n227 CS_BIAS.n191 161.3
R22 CS_BIAS.n226 CS_BIAS.n225 161.3
R23 CS_BIAS.n223 CS_BIAS.n192 161.3
R24 CS_BIAS.n222 CS_BIAS.n221 161.3
R25 CS_BIAS.n220 CS_BIAS.n193 161.3
R26 CS_BIAS.n219 CS_BIAS.n218 161.3
R27 CS_BIAS.n216 CS_BIAS.n194 161.3
R28 CS_BIAS.n215 CS_BIAS.n214 161.3
R29 CS_BIAS.n213 CS_BIAS.n195 161.3
R30 CS_BIAS.n212 CS_BIAS.n211 161.3
R31 CS_BIAS.n210 CS_BIAS.n196 161.3
R32 CS_BIAS.n208 CS_BIAS.n207 161.3
R33 CS_BIAS.n206 CS_BIAS.n197 161.3
R34 CS_BIAS.n205 CS_BIAS.n204 161.3
R35 CS_BIAS.n203 CS_BIAS.n198 161.3
R36 CS_BIAS.n202 CS_BIAS.n201 161.3
R37 CS_BIAS.n36 CS_BIAS.n35 161.3
R38 CS_BIAS.n37 CS_BIAS.n32 161.3
R39 CS_BIAS.n39 CS_BIAS.n38 161.3
R40 CS_BIAS.n40 CS_BIAS.n31 161.3
R41 CS_BIAS.n42 CS_BIAS.n41 161.3
R42 CS_BIAS.n44 CS_BIAS.n30 161.3
R43 CS_BIAS.n46 CS_BIAS.n45 161.3
R44 CS_BIAS.n47 CS_BIAS.n29 161.3
R45 CS_BIAS.n49 CS_BIAS.n48 161.3
R46 CS_BIAS.n50 CS_BIAS.n28 161.3
R47 CS_BIAS.n53 CS_BIAS.n52 161.3
R48 CS_BIAS.n54 CS_BIAS.n27 161.3
R49 CS_BIAS.n56 CS_BIAS.n55 161.3
R50 CS_BIAS.n57 CS_BIAS.n26 161.3
R51 CS_BIAS.n60 CS_BIAS.n59 161.3
R52 CS_BIAS.n61 CS_BIAS.n25 161.3
R53 CS_BIAS.n63 CS_BIAS.n62 161.3
R54 CS_BIAS.n64 CS_BIAS.n23 161.3
R55 CS_BIAS.n66 CS_BIAS.n65 161.3
R56 CS_BIAS.n67 CS_BIAS.n22 161.3
R57 CS_BIAS.n69 CS_BIAS.n68 161.3
R58 CS_BIAS.n70 CS_BIAS.n21 161.3
R59 CS_BIAS.n72 CS_BIAS.n71 161.3
R60 CS_BIAS.n74 CS_BIAS.n73 161.3
R61 CS_BIAS.n75 CS_BIAS.n19 161.3
R62 CS_BIAS.n77 CS_BIAS.n76 161.3
R63 CS_BIAS.n78 CS_BIAS.n18 161.3
R64 CS_BIAS.n80 CS_BIAS.n79 161.3
R65 CS_BIAS.n82 CS_BIAS.n17 161.3
R66 CS_BIAS.n84 CS_BIAS.n83 161.3
R67 CS_BIAS.n85 CS_BIAS.n16 161.3
R68 CS_BIAS.n87 CS_BIAS.n86 161.3
R69 CS_BIAS.n88 CS_BIAS.n15 161.3
R70 CS_BIAS.n91 CS_BIAS.n90 161.3
R71 CS_BIAS.n92 CS_BIAS.n14 161.3
R72 CS_BIAS.n94 CS_BIAS.n93 161.3
R73 CS_BIAS.n95 CS_BIAS.n13 161.3
R74 CS_BIAS.n117 CS_BIAS.n116 161.3
R75 CS_BIAS.n118 CS_BIAS.n113 161.3
R76 CS_BIAS.n120 CS_BIAS.n119 161.3
R77 CS_BIAS.n121 CS_BIAS.n112 161.3
R78 CS_BIAS.n123 CS_BIAS.n122 161.3
R79 CS_BIAS.n125 CS_BIAS.n111 161.3
R80 CS_BIAS.n127 CS_BIAS.n126 161.3
R81 CS_BIAS.n128 CS_BIAS.n110 161.3
R82 CS_BIAS.n130 CS_BIAS.n129 161.3
R83 CS_BIAS.n131 CS_BIAS.n109 161.3
R84 CS_BIAS.n134 CS_BIAS.n133 161.3
R85 CS_BIAS.n135 CS_BIAS.n108 161.3
R86 CS_BIAS.n137 CS_BIAS.n136 161.3
R87 CS_BIAS.n138 CS_BIAS.n107 161.3
R88 CS_BIAS.n141 CS_BIAS.n140 161.3
R89 CS_BIAS.n142 CS_BIAS.n12 161.3
R90 CS_BIAS.n144 CS_BIAS.n143 161.3
R91 CS_BIAS.n145 CS_BIAS.n10 161.3
R92 CS_BIAS.n147 CS_BIAS.n146 161.3
R93 CS_BIAS.n148 CS_BIAS.n9 161.3
R94 CS_BIAS.n150 CS_BIAS.n149 161.3
R95 CS_BIAS.n151 CS_BIAS.n8 161.3
R96 CS_BIAS.n153 CS_BIAS.n152 161.3
R97 CS_BIAS.n155 CS_BIAS.n154 161.3
R98 CS_BIAS.n156 CS_BIAS.n6 161.3
R99 CS_BIAS.n158 CS_BIAS.n157 161.3
R100 CS_BIAS.n159 CS_BIAS.n5 161.3
R101 CS_BIAS.n161 CS_BIAS.n160 161.3
R102 CS_BIAS.n163 CS_BIAS.n4 161.3
R103 CS_BIAS.n165 CS_BIAS.n164 161.3
R104 CS_BIAS.n166 CS_BIAS.n3 161.3
R105 CS_BIAS.n168 CS_BIAS.n167 161.3
R106 CS_BIAS.n169 CS_BIAS.n2 161.3
R107 CS_BIAS.n172 CS_BIAS.n171 161.3
R108 CS_BIAS.n173 CS_BIAS.n1 161.3
R109 CS_BIAS.n175 CS_BIAS.n174 161.3
R110 CS_BIAS.n176 CS_BIAS.n0 161.3
R111 CS_BIAS.n526 CS_BIAS.n444 161.3
R112 CS_BIAS.n525 CS_BIAS.n524 161.3
R113 CS_BIAS.n523 CS_BIAS.n445 161.3
R114 CS_BIAS.n522 CS_BIAS.n521 161.3
R115 CS_BIAS.n519 CS_BIAS.n446 161.3
R116 CS_BIAS.n518 CS_BIAS.n517 161.3
R117 CS_BIAS.n516 CS_BIAS.n447 161.3
R118 CS_BIAS.n515 CS_BIAS.n514 161.3
R119 CS_BIAS.n513 CS_BIAS.n448 161.3
R120 CS_BIAS.n511 CS_BIAS.n510 161.3
R121 CS_BIAS.n509 CS_BIAS.n449 161.3
R122 CS_BIAS.n508 CS_BIAS.n507 161.3
R123 CS_BIAS.n506 CS_BIAS.n450 161.3
R124 CS_BIAS.n505 CS_BIAS.n504 161.3
R125 CS_BIAS.n503 CS_BIAS.n502 161.3
R126 CS_BIAS.n501 CS_BIAS.n452 161.3
R127 CS_BIAS.n500 CS_BIAS.n499 161.3
R128 CS_BIAS.n498 CS_BIAS.n453 161.3
R129 CS_BIAS.n497 CS_BIAS.n496 161.3
R130 CS_BIAS.n494 CS_BIAS.n454 161.3
R131 CS_BIAS.n493 CS_BIAS.n492 161.3
R132 CS_BIAS.n491 CS_BIAS.n455 161.3
R133 CS_BIAS.n490 CS_BIAS.n489 161.3
R134 CS_BIAS.n487 CS_BIAS.n456 161.3
R135 CS_BIAS.n486 CS_BIAS.n485 161.3
R136 CS_BIAS.n484 CS_BIAS.n457 161.3
R137 CS_BIAS.n483 CS_BIAS.n482 161.3
R138 CS_BIAS.n480 CS_BIAS.n458 161.3
R139 CS_BIAS.n479 CS_BIAS.n478 161.3
R140 CS_BIAS.n477 CS_BIAS.n459 161.3
R141 CS_BIAS.n476 CS_BIAS.n475 161.3
R142 CS_BIAS.n474 CS_BIAS.n460 161.3
R143 CS_BIAS.n472 CS_BIAS.n471 161.3
R144 CS_BIAS.n470 CS_BIAS.n461 161.3
R145 CS_BIAS.n469 CS_BIAS.n468 161.3
R146 CS_BIAS.n467 CS_BIAS.n462 161.3
R147 CS_BIAS.n466 CS_BIAS.n465 161.3
R148 CS_BIAS.n399 CS_BIAS.n317 161.3
R149 CS_BIAS.n398 CS_BIAS.n397 161.3
R150 CS_BIAS.n396 CS_BIAS.n318 161.3
R151 CS_BIAS.n395 CS_BIAS.n394 161.3
R152 CS_BIAS.n392 CS_BIAS.n319 161.3
R153 CS_BIAS.n391 CS_BIAS.n390 161.3
R154 CS_BIAS.n389 CS_BIAS.n320 161.3
R155 CS_BIAS.n388 CS_BIAS.n387 161.3
R156 CS_BIAS.n386 CS_BIAS.n321 161.3
R157 CS_BIAS.n384 CS_BIAS.n383 161.3
R158 CS_BIAS.n382 CS_BIAS.n322 161.3
R159 CS_BIAS.n381 CS_BIAS.n380 161.3
R160 CS_BIAS.n379 CS_BIAS.n323 161.3
R161 CS_BIAS.n378 CS_BIAS.n377 161.3
R162 CS_BIAS.n376 CS_BIAS.n375 161.3
R163 CS_BIAS.n374 CS_BIAS.n325 161.3
R164 CS_BIAS.n373 CS_BIAS.n372 161.3
R165 CS_BIAS.n371 CS_BIAS.n326 161.3
R166 CS_BIAS.n370 CS_BIAS.n369 161.3
R167 CS_BIAS.n367 CS_BIAS.n327 161.3
R168 CS_BIAS.n366 CS_BIAS.n365 161.3
R169 CS_BIAS.n364 CS_BIAS.n328 161.3
R170 CS_BIAS.n363 CS_BIAS.n362 161.3
R171 CS_BIAS.n360 CS_BIAS.n329 161.3
R172 CS_BIAS.n359 CS_BIAS.n358 161.3
R173 CS_BIAS.n357 CS_BIAS.n330 161.3
R174 CS_BIAS.n356 CS_BIAS.n355 161.3
R175 CS_BIAS.n353 CS_BIAS.n331 161.3
R176 CS_BIAS.n352 CS_BIAS.n351 161.3
R177 CS_BIAS.n350 CS_BIAS.n332 161.3
R178 CS_BIAS.n349 CS_BIAS.n348 161.3
R179 CS_BIAS.n347 CS_BIAS.n333 161.3
R180 CS_BIAS.n345 CS_BIAS.n344 161.3
R181 CS_BIAS.n343 CS_BIAS.n334 161.3
R182 CS_BIAS.n342 CS_BIAS.n341 161.3
R183 CS_BIAS.n340 CS_BIAS.n335 161.3
R184 CS_BIAS.n339 CS_BIAS.n338 161.3
R185 CS_BIAS.n312 CS_BIAS.n276 161.3
R186 CS_BIAS.n311 CS_BIAS.n310 161.3
R187 CS_BIAS.n308 CS_BIAS.n277 161.3
R188 CS_BIAS.n307 CS_BIAS.n306 161.3
R189 CS_BIAS.n305 CS_BIAS.n278 161.3
R190 CS_BIAS.n304 CS_BIAS.n303 161.3
R191 CS_BIAS.n301 CS_BIAS.n279 161.3
R192 CS_BIAS.n300 CS_BIAS.n299 161.3
R193 CS_BIAS.n298 CS_BIAS.n280 161.3
R194 CS_BIAS.n297 CS_BIAS.n296 161.3
R195 CS_BIAS.n295 CS_BIAS.n281 161.3
R196 CS_BIAS.n293 CS_BIAS.n292 161.3
R197 CS_BIAS.n291 CS_BIAS.n282 161.3
R198 CS_BIAS.n290 CS_BIAS.n289 161.3
R199 CS_BIAS.n288 CS_BIAS.n283 161.3
R200 CS_BIAS.n287 CS_BIAS.n286 161.3
R201 CS_BIAS.n408 CS_BIAS.n407 161.3
R202 CS_BIAS.n441 CS_BIAS.n265 161.3
R203 CS_BIAS.n440 CS_BIAS.n439 161.3
R204 CS_BIAS.n438 CS_BIAS.n266 161.3
R205 CS_BIAS.n437 CS_BIAS.n436 161.3
R206 CS_BIAS.n434 CS_BIAS.n267 161.3
R207 CS_BIAS.n433 CS_BIAS.n432 161.3
R208 CS_BIAS.n431 CS_BIAS.n268 161.3
R209 CS_BIAS.n430 CS_BIAS.n429 161.3
R210 CS_BIAS.n428 CS_BIAS.n269 161.3
R211 CS_BIAS.n426 CS_BIAS.n425 161.3
R212 CS_BIAS.n424 CS_BIAS.n270 161.3
R213 CS_BIAS.n423 CS_BIAS.n422 161.3
R214 CS_BIAS.n421 CS_BIAS.n271 161.3
R215 CS_BIAS.n420 CS_BIAS.n419 161.3
R216 CS_BIAS.n418 CS_BIAS.n417 161.3
R217 CS_BIAS.n416 CS_BIAS.n273 161.3
R218 CS_BIAS.n415 CS_BIAS.n414 161.3
R219 CS_BIAS.n413 CS_BIAS.n274 161.3
R220 CS_BIAS.n412 CS_BIAS.n411 161.3
R221 CS_BIAS.n409 CS_BIAS.n275 161.3
R222 CS_BIAS.n200 CS_BIAS.t73 115.436
R223 CS_BIAS.n34 CS_BIAS.t12 115.436
R224 CS_BIAS.n115 CS_BIAS.t56 115.436
R225 CS_BIAS.n464 CS_BIAS.t49 115.436
R226 CS_BIAS.n337 CS_BIAS.t10 115.436
R227 CS_BIAS.n285 CS_BIAS.t70 115.436
R228 CS_BIAS.n263 CS_BIAS.n262 87.0542
R229 CS_BIAS.n97 CS_BIAS.n96 87.0542
R230 CS_BIAS.n178 CS_BIAS.n177 87.0542
R231 CS_BIAS.n528 CS_BIAS.n527 87.0542
R232 CS_BIAS.n401 CS_BIAS.n400 87.0542
R233 CS_BIAS.n443 CS_BIAS.n442 87.0542
R234 CS_BIAS.n199 CS_BIAS.t72 84.3505
R235 CS_BIAS.n209 CS_BIAS.t45 84.3505
R236 CS_BIAS.n217 CS_BIAS.t42 84.3505
R237 CS_BIAS.n224 CS_BIAS.t53 84.3505
R238 CS_BIAS.n190 CS_BIAS.t51 84.3505
R239 CS_BIAS.n186 CS_BIAS.t74 84.3505
R240 CS_BIAS.n247 CS_BIAS.t78 84.3505
R241 CS_BIAS.n255 CS_BIAS.t75 84.3505
R242 CS_BIAS.n262 CS_BIAS.t57 84.3505
R243 CS_BIAS.n96 CS_BIAS.t32 84.3505
R244 CS_BIAS.n89 CS_BIAS.t26 84.3505
R245 CS_BIAS.n81 CS_BIAS.t0 84.3505
R246 CS_BIAS.n20 CS_BIAS.t38 84.3505
R247 CS_BIAS.n24 CS_BIAS.t34 84.3505
R248 CS_BIAS.n58 CS_BIAS.t36 84.3505
R249 CS_BIAS.n51 CS_BIAS.t28 84.3505
R250 CS_BIAS.n43 CS_BIAS.t24 84.3505
R251 CS_BIAS.n33 CS_BIAS.t4 84.3505
R252 CS_BIAS.n177 CS_BIAS.t40 84.3505
R253 CS_BIAS.n170 CS_BIAS.t58 84.3505
R254 CS_BIAS.n162 CS_BIAS.t60 84.3505
R255 CS_BIAS.n7 CS_BIAS.t59 84.3505
R256 CS_BIAS.n11 CS_BIAS.t77 84.3505
R257 CS_BIAS.n139 CS_BIAS.t79 84.3505
R258 CS_BIAS.n132 CS_BIAS.t66 84.3505
R259 CS_BIAS.n124 CS_BIAS.t68 84.3505
R260 CS_BIAS.n114 CS_BIAS.t55 84.3505
R261 CS_BIAS.n463 CS_BIAS.t62 84.3505
R262 CS_BIAS.n473 CS_BIAS.t61 84.3505
R263 CS_BIAS.n481 CS_BIAS.t69 84.3505
R264 CS_BIAS.n488 CS_BIAS.t44 84.3505
R265 CS_BIAS.n495 CS_BIAS.t41 84.3505
R266 CS_BIAS.n451 CS_BIAS.t63 84.3505
R267 CS_BIAS.n512 CS_BIAS.t50 84.3505
R268 CS_BIAS.n520 CS_BIAS.t64 84.3505
R269 CS_BIAS.n527 CS_BIAS.t71 84.3505
R270 CS_BIAS.n336 CS_BIAS.t6 84.3505
R271 CS_BIAS.n346 CS_BIAS.t2 84.3505
R272 CS_BIAS.n354 CS_BIAS.t22 84.3505
R273 CS_BIAS.n361 CS_BIAS.t14 84.3505
R274 CS_BIAS.n368 CS_BIAS.t8 84.3505
R275 CS_BIAS.n324 CS_BIAS.t16 84.3505
R276 CS_BIAS.n385 CS_BIAS.t18 84.3505
R277 CS_BIAS.n393 CS_BIAS.t20 84.3505
R278 CS_BIAS.n400 CS_BIAS.t30 84.3505
R279 CS_BIAS.n442 CS_BIAS.t54 84.3505
R280 CS_BIAS.n435 CS_BIAS.t48 84.3505
R281 CS_BIAS.n427 CS_BIAS.t76 84.3505
R282 CS_BIAS.n272 CS_BIAS.t47 84.3505
R283 CS_BIAS.n410 CS_BIAS.t65 84.3505
R284 CS_BIAS.n284 CS_BIAS.t46 84.3505
R285 CS_BIAS.n294 CS_BIAS.t43 84.3505
R286 CS_BIAS.n302 CS_BIAS.t52 84.3505
R287 CS_BIAS.n309 CS_BIAS.t67 84.3505
R288 CS_BIAS.n105 CS_BIAS.n103 81.9368
R289 CS_BIAS.n315 CS_BIAS.n313 81.9368
R290 CS_BIAS.n105 CS_BIAS.n104 80.9324
R291 CS_BIAS.n106 CS_BIAS.n102 80.9324
R292 CS_BIAS.n101 CS_BIAS.n100 80.9324
R293 CS_BIAS.n99 CS_BIAS.n98 80.9324
R294 CS_BIAS.n403 CS_BIAS.n402 80.9324
R295 CS_BIAS.n405 CS_BIAS.n404 80.9324
R296 CS_BIAS.n406 CS_BIAS.n316 80.9324
R297 CS_BIAS.n315 CS_BIAS.n314 80.9324
R298 CS_BIAS.n200 CS_BIAS.n199 62.9271
R299 CS_BIAS.n34 CS_BIAS.n33 62.9271
R300 CS_BIAS.n115 CS_BIAS.n114 62.9271
R301 CS_BIAS.n464 CS_BIAS.n463 62.9271
R302 CS_BIAS.n337 CS_BIAS.n336 62.9271
R303 CS_BIAS.n285 CS_BIAS.n284 62.9271
R304 CS_BIAS.n222 CS_BIAS.n193 56.5617
R305 CS_BIAS.n236 CS_BIAS.n235 56.5617
R306 CS_BIAS.n260 CS_BIAS.n180 56.5617
R307 CS_BIAS.n94 CS_BIAS.n14 56.5617
R308 CS_BIAS.n70 CS_BIAS.n69 56.5617
R309 CS_BIAS.n56 CS_BIAS.n27 56.5617
R310 CS_BIAS.n175 CS_BIAS.n1 56.5617
R311 CS_BIAS.n151 CS_BIAS.n150 56.5617
R312 CS_BIAS.n137 CS_BIAS.n108 56.5617
R313 CS_BIAS.n486 CS_BIAS.n457 56.5617
R314 CS_BIAS.n501 CS_BIAS.n500 56.5617
R315 CS_BIAS.n525 CS_BIAS.n445 56.5617
R316 CS_BIAS.n359 CS_BIAS.n330 56.5617
R317 CS_BIAS.n374 CS_BIAS.n373 56.5617
R318 CS_BIAS.n398 CS_BIAS.n318 56.5617
R319 CS_BIAS.n440 CS_BIAS.n266 56.5617
R320 CS_BIAS.n416 CS_BIAS.n415 56.5617
R321 CS_BIAS.n307 CS_BIAS.n278 56.5617
R322 CS_BIAS.n211 CS_BIAS.n195 56.0773
R323 CS_BIAS.n242 CS_BIAS.n184 56.0773
R324 CS_BIAS.n76 CS_BIAS.n18 56.0773
R325 CS_BIAS.n45 CS_BIAS.n29 56.0773
R326 CS_BIAS.n157 CS_BIAS.n5 56.0773
R327 CS_BIAS.n126 CS_BIAS.n110 56.0773
R328 CS_BIAS.n475 CS_BIAS.n459 56.0773
R329 CS_BIAS.n507 CS_BIAS.n449 56.0773
R330 CS_BIAS.n348 CS_BIAS.n332 56.0773
R331 CS_BIAS.n380 CS_BIAS.n322 56.0773
R332 CS_BIAS.n422 CS_BIAS.n270 56.0773
R333 CS_BIAS.n296 CS_BIAS.n280 56.0773
R334 CS_BIAS.n204 CS_BIAS.n197 41.5458
R335 CS_BIAS.n249 CS_BIAS.n182 41.5458
R336 CS_BIAS.n83 CS_BIAS.n16 41.5458
R337 CS_BIAS.n38 CS_BIAS.n31 41.5458
R338 CS_BIAS.n164 CS_BIAS.n3 41.5458
R339 CS_BIAS.n119 CS_BIAS.n112 41.5458
R340 CS_BIAS.n468 CS_BIAS.n461 41.5458
R341 CS_BIAS.n514 CS_BIAS.n447 41.5458
R342 CS_BIAS.n341 CS_BIAS.n334 41.5458
R343 CS_BIAS.n387 CS_BIAS.n320 41.5458
R344 CS_BIAS.n429 CS_BIAS.n268 41.5458
R345 CS_BIAS.n289 CS_BIAS.n282 41.5458
R346 CS_BIAS.n229 CS_BIAS.n191 40.577
R347 CS_BIAS.n230 CS_BIAS.n229 40.577
R348 CS_BIAS.n64 CS_BIAS.n63 40.577
R349 CS_BIAS.n63 CS_BIAS.n25 40.577
R350 CS_BIAS.n145 CS_BIAS.n144 40.577
R351 CS_BIAS.n144 CS_BIAS.n12 40.577
R352 CS_BIAS.n493 CS_BIAS.n455 40.577
R353 CS_BIAS.n494 CS_BIAS.n493 40.577
R354 CS_BIAS.n366 CS_BIAS.n328 40.577
R355 CS_BIAS.n367 CS_BIAS.n366 40.577
R356 CS_BIAS.n409 CS_BIAS.n408 40.577
R357 CS_BIAS.n408 CS_BIAS.n276 40.577
R358 CS_BIAS.n204 CS_BIAS.n203 39.6083
R359 CS_BIAS.n253 CS_BIAS.n182 39.6083
R360 CS_BIAS.n87 CS_BIAS.n16 39.6083
R361 CS_BIAS.n38 CS_BIAS.n37 39.6083
R362 CS_BIAS.n168 CS_BIAS.n3 39.6083
R363 CS_BIAS.n119 CS_BIAS.n118 39.6083
R364 CS_BIAS.n468 CS_BIAS.n467 39.6083
R365 CS_BIAS.n518 CS_BIAS.n447 39.6083
R366 CS_BIAS.n341 CS_BIAS.n340 39.6083
R367 CS_BIAS.n391 CS_BIAS.n320 39.6083
R368 CS_BIAS.n433 CS_BIAS.n268 39.6083
R369 CS_BIAS.n289 CS_BIAS.n288 39.6083
R370 CS_BIAS.n215 CS_BIAS.n195 25.0767
R371 CS_BIAS.n242 CS_BIAS.n241 25.0767
R372 CS_BIAS.n76 CS_BIAS.n75 25.0767
R373 CS_BIAS.n49 CS_BIAS.n29 25.0767
R374 CS_BIAS.n157 CS_BIAS.n156 25.0767
R375 CS_BIAS.n130 CS_BIAS.n110 25.0767
R376 CS_BIAS.n479 CS_BIAS.n459 25.0767
R377 CS_BIAS.n507 CS_BIAS.n506 25.0767
R378 CS_BIAS.n352 CS_BIAS.n332 25.0767
R379 CS_BIAS.n380 CS_BIAS.n379 25.0767
R380 CS_BIAS.n422 CS_BIAS.n421 25.0767
R381 CS_BIAS.n300 CS_BIAS.n280 25.0767
R382 CS_BIAS.n203 CS_BIAS.n202 24.5923
R383 CS_BIAS.n211 CS_BIAS.n210 24.5923
R384 CS_BIAS.n208 CS_BIAS.n197 24.5923
R385 CS_BIAS.n218 CS_BIAS.n193 24.5923
R386 CS_BIAS.n216 CS_BIAS.n215 24.5923
R387 CS_BIAS.n225 CS_BIAS.n191 24.5923
R388 CS_BIAS.n223 CS_BIAS.n222 24.5923
R389 CS_BIAS.n235 CS_BIAS.n188 24.5923
R390 CS_BIAS.n231 CS_BIAS.n230 24.5923
R391 CS_BIAS.n241 CS_BIAS.n240 24.5923
R392 CS_BIAS.n237 CS_BIAS.n236 24.5923
R393 CS_BIAS.n249 CS_BIAS.n248 24.5923
R394 CS_BIAS.n246 CS_BIAS.n184 24.5923
R395 CS_BIAS.n256 CS_BIAS.n180 24.5923
R396 CS_BIAS.n254 CS_BIAS.n253 24.5923
R397 CS_BIAS.n261 CS_BIAS.n260 24.5923
R398 CS_BIAS.n95 CS_BIAS.n94 24.5923
R399 CS_BIAS.n90 CS_BIAS.n14 24.5923
R400 CS_BIAS.n88 CS_BIAS.n87 24.5923
R401 CS_BIAS.n83 CS_BIAS.n82 24.5923
R402 CS_BIAS.n80 CS_BIAS.n18 24.5923
R403 CS_BIAS.n75 CS_BIAS.n74 24.5923
R404 CS_BIAS.n71 CS_BIAS.n70 24.5923
R405 CS_BIAS.n69 CS_BIAS.n22 24.5923
R406 CS_BIAS.n65 CS_BIAS.n64 24.5923
R407 CS_BIAS.n59 CS_BIAS.n25 24.5923
R408 CS_BIAS.n57 CS_BIAS.n56 24.5923
R409 CS_BIAS.n52 CS_BIAS.n27 24.5923
R410 CS_BIAS.n50 CS_BIAS.n49 24.5923
R411 CS_BIAS.n45 CS_BIAS.n44 24.5923
R412 CS_BIAS.n42 CS_BIAS.n31 24.5923
R413 CS_BIAS.n37 CS_BIAS.n36 24.5923
R414 CS_BIAS.n176 CS_BIAS.n175 24.5923
R415 CS_BIAS.n171 CS_BIAS.n1 24.5923
R416 CS_BIAS.n169 CS_BIAS.n168 24.5923
R417 CS_BIAS.n164 CS_BIAS.n163 24.5923
R418 CS_BIAS.n161 CS_BIAS.n5 24.5923
R419 CS_BIAS.n156 CS_BIAS.n155 24.5923
R420 CS_BIAS.n152 CS_BIAS.n151 24.5923
R421 CS_BIAS.n150 CS_BIAS.n9 24.5923
R422 CS_BIAS.n146 CS_BIAS.n145 24.5923
R423 CS_BIAS.n140 CS_BIAS.n12 24.5923
R424 CS_BIAS.n138 CS_BIAS.n137 24.5923
R425 CS_BIAS.n133 CS_BIAS.n108 24.5923
R426 CS_BIAS.n131 CS_BIAS.n130 24.5923
R427 CS_BIAS.n126 CS_BIAS.n125 24.5923
R428 CS_BIAS.n123 CS_BIAS.n112 24.5923
R429 CS_BIAS.n118 CS_BIAS.n117 24.5923
R430 CS_BIAS.n467 CS_BIAS.n466 24.5923
R431 CS_BIAS.n472 CS_BIAS.n461 24.5923
R432 CS_BIAS.n475 CS_BIAS.n474 24.5923
R433 CS_BIAS.n480 CS_BIAS.n479 24.5923
R434 CS_BIAS.n482 CS_BIAS.n457 24.5923
R435 CS_BIAS.n487 CS_BIAS.n486 24.5923
R436 CS_BIAS.n489 CS_BIAS.n455 24.5923
R437 CS_BIAS.n496 CS_BIAS.n494 24.5923
R438 CS_BIAS.n500 CS_BIAS.n453 24.5923
R439 CS_BIAS.n502 CS_BIAS.n501 24.5923
R440 CS_BIAS.n506 CS_BIAS.n505 24.5923
R441 CS_BIAS.n511 CS_BIAS.n449 24.5923
R442 CS_BIAS.n514 CS_BIAS.n513 24.5923
R443 CS_BIAS.n519 CS_BIAS.n518 24.5923
R444 CS_BIAS.n521 CS_BIAS.n445 24.5923
R445 CS_BIAS.n526 CS_BIAS.n525 24.5923
R446 CS_BIAS.n340 CS_BIAS.n339 24.5923
R447 CS_BIAS.n345 CS_BIAS.n334 24.5923
R448 CS_BIAS.n348 CS_BIAS.n347 24.5923
R449 CS_BIAS.n353 CS_BIAS.n352 24.5923
R450 CS_BIAS.n355 CS_BIAS.n330 24.5923
R451 CS_BIAS.n360 CS_BIAS.n359 24.5923
R452 CS_BIAS.n362 CS_BIAS.n328 24.5923
R453 CS_BIAS.n369 CS_BIAS.n367 24.5923
R454 CS_BIAS.n373 CS_BIAS.n326 24.5923
R455 CS_BIAS.n375 CS_BIAS.n374 24.5923
R456 CS_BIAS.n379 CS_BIAS.n378 24.5923
R457 CS_BIAS.n384 CS_BIAS.n322 24.5923
R458 CS_BIAS.n387 CS_BIAS.n386 24.5923
R459 CS_BIAS.n392 CS_BIAS.n391 24.5923
R460 CS_BIAS.n394 CS_BIAS.n318 24.5923
R461 CS_BIAS.n399 CS_BIAS.n398 24.5923
R462 CS_BIAS.n441 CS_BIAS.n440 24.5923
R463 CS_BIAS.n434 CS_BIAS.n433 24.5923
R464 CS_BIAS.n436 CS_BIAS.n266 24.5923
R465 CS_BIAS.n426 CS_BIAS.n270 24.5923
R466 CS_BIAS.n429 CS_BIAS.n428 24.5923
R467 CS_BIAS.n417 CS_BIAS.n416 24.5923
R468 CS_BIAS.n421 CS_BIAS.n420 24.5923
R469 CS_BIAS.n411 CS_BIAS.n409 24.5923
R470 CS_BIAS.n415 CS_BIAS.n274 24.5923
R471 CS_BIAS.n288 CS_BIAS.n287 24.5923
R472 CS_BIAS.n293 CS_BIAS.n282 24.5923
R473 CS_BIAS.n296 CS_BIAS.n295 24.5923
R474 CS_BIAS.n301 CS_BIAS.n300 24.5923
R475 CS_BIAS.n303 CS_BIAS.n278 24.5923
R476 CS_BIAS.n308 CS_BIAS.n307 24.5923
R477 CS_BIAS.n310 CS_BIAS.n276 24.5923
R478 CS_BIAS.n218 CS_BIAS.n217 24.3464
R479 CS_BIAS.n237 CS_BIAS.n186 24.3464
R480 CS_BIAS.n71 CS_BIAS.n20 24.3464
R481 CS_BIAS.n52 CS_BIAS.n51 24.3464
R482 CS_BIAS.n152 CS_BIAS.n7 24.3464
R483 CS_BIAS.n133 CS_BIAS.n132 24.3464
R484 CS_BIAS.n482 CS_BIAS.n481 24.3464
R485 CS_BIAS.n502 CS_BIAS.n451 24.3464
R486 CS_BIAS.n355 CS_BIAS.n354 24.3464
R487 CS_BIAS.n375 CS_BIAS.n324 24.3464
R488 CS_BIAS.n417 CS_BIAS.n272 24.3464
R489 CS_BIAS.n303 CS_BIAS.n302 24.3464
R490 CS_BIAS.n262 CS_BIAS.n261 23.8546
R491 CS_BIAS.n96 CS_BIAS.n95 23.8546
R492 CS_BIAS.n177 CS_BIAS.n176 23.8546
R493 CS_BIAS.n527 CS_BIAS.n526 23.8546
R494 CS_BIAS.n400 CS_BIAS.n399 23.8546
R495 CS_BIAS.n442 CS_BIAS.n441 23.8546
R496 CS_BIAS.n256 CS_BIAS.n255 16.9689
R497 CS_BIAS.n90 CS_BIAS.n89 16.9689
R498 CS_BIAS.n171 CS_BIAS.n170 16.9689
R499 CS_BIAS.n521 CS_BIAS.n520 16.9689
R500 CS_BIAS.n394 CS_BIAS.n393 16.9689
R501 CS_BIAS.n436 CS_BIAS.n435 16.9689
R502 CS_BIAS.n224 CS_BIAS.n223 16.477
R503 CS_BIAS.n190 CS_BIAS.n188 16.477
R504 CS_BIAS.n24 CS_BIAS.n22 16.477
R505 CS_BIAS.n58 CS_BIAS.n57 16.477
R506 CS_BIAS.n11 CS_BIAS.n9 16.477
R507 CS_BIAS.n139 CS_BIAS.n138 16.477
R508 CS_BIAS.n488 CS_BIAS.n487 16.477
R509 CS_BIAS.n495 CS_BIAS.n453 16.477
R510 CS_BIAS.n361 CS_BIAS.n360 16.477
R511 CS_BIAS.n368 CS_BIAS.n326 16.477
R512 CS_BIAS.n410 CS_BIAS.n274 16.477
R513 CS_BIAS.n309 CS_BIAS.n308 16.477
R514 CS_BIAS.n210 CS_BIAS.n209 15.9852
R515 CS_BIAS.n247 CS_BIAS.n246 15.9852
R516 CS_BIAS.n81 CS_BIAS.n80 15.9852
R517 CS_BIAS.n44 CS_BIAS.n43 15.9852
R518 CS_BIAS.n162 CS_BIAS.n161 15.9852
R519 CS_BIAS.n125 CS_BIAS.n124 15.9852
R520 CS_BIAS.n474 CS_BIAS.n473 15.9852
R521 CS_BIAS.n512 CS_BIAS.n511 15.9852
R522 CS_BIAS.n347 CS_BIAS.n346 15.9852
R523 CS_BIAS.n385 CS_BIAS.n384 15.9852
R524 CS_BIAS.n427 CS_BIAS.n426 15.9852
R525 CS_BIAS.n295 CS_BIAS.n294 15.9852
R526 CS_BIAS.n99 CS_BIAS.n97 13.4923
R527 CS_BIAS.n403 CS_BIAS.n401 13.4923
R528 CS_BIAS.n201 CS_BIAS.n200 12.7518
R529 CS_BIAS.n35 CS_BIAS.n34 12.7518
R530 CS_BIAS.n116 CS_BIAS.n115 12.7518
R531 CS_BIAS.n465 CS_BIAS.n464 12.7518
R532 CS_BIAS.n338 CS_BIAS.n337 12.7518
R533 CS_BIAS.n286 CS_BIAS.n285 12.7518
R534 CS_BIAS.n530 CS_BIAS.n264 11.3868
R535 CS_BIAS.n530 CS_BIAS.n529 9.93702
R536 CS_BIAS.n143 CS_BIAS.n106 9.50363
R537 CS_BIAS.n407 CS_BIAS.n406 9.50363
R538 CS_BIAS.n264 CS_BIAS.n178 8.76523
R539 CS_BIAS.n529 CS_BIAS.n443 8.76523
R540 CS_BIAS.n209 CS_BIAS.n208 8.60764
R541 CS_BIAS.n248 CS_BIAS.n247 8.60764
R542 CS_BIAS.n82 CS_BIAS.n81 8.60764
R543 CS_BIAS.n43 CS_BIAS.n42 8.60764
R544 CS_BIAS.n163 CS_BIAS.n162 8.60764
R545 CS_BIAS.n124 CS_BIAS.n123 8.60764
R546 CS_BIAS.n473 CS_BIAS.n472 8.60764
R547 CS_BIAS.n513 CS_BIAS.n512 8.60764
R548 CS_BIAS.n346 CS_BIAS.n345 8.60764
R549 CS_BIAS.n386 CS_BIAS.n385 8.60764
R550 CS_BIAS.n428 CS_BIAS.n427 8.60764
R551 CS_BIAS.n294 CS_BIAS.n293 8.60764
R552 CS_BIAS.n225 CS_BIAS.n224 8.11581
R553 CS_BIAS.n231 CS_BIAS.n190 8.11581
R554 CS_BIAS.n65 CS_BIAS.n24 8.11581
R555 CS_BIAS.n59 CS_BIAS.n58 8.11581
R556 CS_BIAS.n146 CS_BIAS.n11 8.11581
R557 CS_BIAS.n140 CS_BIAS.n139 8.11581
R558 CS_BIAS.n489 CS_BIAS.n488 8.11581
R559 CS_BIAS.n496 CS_BIAS.n495 8.11581
R560 CS_BIAS.n362 CS_BIAS.n361 8.11581
R561 CS_BIAS.n369 CS_BIAS.n368 8.11581
R562 CS_BIAS.n411 CS_BIAS.n410 8.11581
R563 CS_BIAS.n310 CS_BIAS.n309 8.11581
R564 CS_BIAS.n202 CS_BIAS.n199 7.62397
R565 CS_BIAS.n255 CS_BIAS.n254 7.62397
R566 CS_BIAS.n89 CS_BIAS.n88 7.62397
R567 CS_BIAS.n36 CS_BIAS.n33 7.62397
R568 CS_BIAS.n170 CS_BIAS.n169 7.62397
R569 CS_BIAS.n117 CS_BIAS.n114 7.62397
R570 CS_BIAS.n466 CS_BIAS.n463 7.62397
R571 CS_BIAS.n520 CS_BIAS.n519 7.62397
R572 CS_BIAS.n339 CS_BIAS.n336 7.62397
R573 CS_BIAS.n393 CS_BIAS.n392 7.62397
R574 CS_BIAS.n435 CS_BIAS.n434 7.62397
R575 CS_BIAS.n287 CS_BIAS.n284 7.62397
R576 CS_BIAS.n264 CS_BIAS.n263 5.07583
R577 CS_BIAS.n529 CS_BIAS.n528 5.07583
R578 CS_BIAS CS_BIAS.n530 4.06627
R579 CS_BIAS.n103 CS_BIAS.t5 2.82907
R580 CS_BIAS.n103 CS_BIAS.t13 2.82907
R581 CS_BIAS.n104 CS_BIAS.t29 2.82907
R582 CS_BIAS.n104 CS_BIAS.t25 2.82907
R583 CS_BIAS.n102 CS_BIAS.t35 2.82907
R584 CS_BIAS.n102 CS_BIAS.t37 2.82907
R585 CS_BIAS.n100 CS_BIAS.t1 2.82907
R586 CS_BIAS.n100 CS_BIAS.t39 2.82907
R587 CS_BIAS.n98 CS_BIAS.t33 2.82907
R588 CS_BIAS.n98 CS_BIAS.t27 2.82907
R589 CS_BIAS.n402 CS_BIAS.t21 2.82907
R590 CS_BIAS.n402 CS_BIAS.t31 2.82907
R591 CS_BIAS.n404 CS_BIAS.t17 2.82907
R592 CS_BIAS.n404 CS_BIAS.t19 2.82907
R593 CS_BIAS.n316 CS_BIAS.t15 2.82907
R594 CS_BIAS.n316 CS_BIAS.t9 2.82907
R595 CS_BIAS.n314 CS_BIAS.t3 2.82907
R596 CS_BIAS.n314 CS_BIAS.t23 2.82907
R597 CS_BIAS.n313 CS_BIAS.t11 2.82907
R598 CS_BIAS.n313 CS_BIAS.t7 2.82907
R599 CS_BIAS.n101 CS_BIAS.n99 1.00481
R600 CS_BIAS.n106 CS_BIAS.n101 1.00481
R601 CS_BIAS.n106 CS_BIAS.n105 1.00481
R602 CS_BIAS.n406 CS_BIAS.n315 1.00481
R603 CS_BIAS.n406 CS_BIAS.n405 1.00481
R604 CS_BIAS.n405 CS_BIAS.n403 1.00481
R605 CS_BIAS.n263 CS_BIAS.n179 0.278335
R606 CS_BIAS.n97 CS_BIAS.n13 0.278335
R607 CS_BIAS.n178 CS_BIAS.n0 0.278335
R608 CS_BIAS.n528 CS_BIAS.n444 0.278335
R609 CS_BIAS.n401 CS_BIAS.n317 0.278335
R610 CS_BIAS.n443 CS_BIAS.n265 0.278335
R611 CS_BIAS.n217 CS_BIAS.n216 0.246418
R612 CS_BIAS.n240 CS_BIAS.n186 0.246418
R613 CS_BIAS.n74 CS_BIAS.n20 0.246418
R614 CS_BIAS.n51 CS_BIAS.n50 0.246418
R615 CS_BIAS.n155 CS_BIAS.n7 0.246418
R616 CS_BIAS.n132 CS_BIAS.n131 0.246418
R617 CS_BIAS.n481 CS_BIAS.n480 0.246418
R618 CS_BIAS.n505 CS_BIAS.n451 0.246418
R619 CS_BIAS.n354 CS_BIAS.n353 0.246418
R620 CS_BIAS.n378 CS_BIAS.n324 0.246418
R621 CS_BIAS.n420 CS_BIAS.n272 0.246418
R622 CS_BIAS.n302 CS_BIAS.n301 0.246418
R623 CS_BIAS.n259 CS_BIAS.n179 0.189894
R624 CS_BIAS.n259 CS_BIAS.n258 0.189894
R625 CS_BIAS.n258 CS_BIAS.n257 0.189894
R626 CS_BIAS.n257 CS_BIAS.n181 0.189894
R627 CS_BIAS.n252 CS_BIAS.n181 0.189894
R628 CS_BIAS.n252 CS_BIAS.n251 0.189894
R629 CS_BIAS.n251 CS_BIAS.n250 0.189894
R630 CS_BIAS.n250 CS_BIAS.n183 0.189894
R631 CS_BIAS.n245 CS_BIAS.n183 0.189894
R632 CS_BIAS.n245 CS_BIAS.n244 0.189894
R633 CS_BIAS.n244 CS_BIAS.n243 0.189894
R634 CS_BIAS.n243 CS_BIAS.n185 0.189894
R635 CS_BIAS.n239 CS_BIAS.n185 0.189894
R636 CS_BIAS.n239 CS_BIAS.n238 0.189894
R637 CS_BIAS.n238 CS_BIAS.n187 0.189894
R638 CS_BIAS.n234 CS_BIAS.n187 0.189894
R639 CS_BIAS.n234 CS_BIAS.n233 0.189894
R640 CS_BIAS.n233 CS_BIAS.n232 0.189894
R641 CS_BIAS.n232 CS_BIAS.n189 0.189894
R642 CS_BIAS.n228 CS_BIAS.n189 0.189894
R643 CS_BIAS.n228 CS_BIAS.n227 0.189894
R644 CS_BIAS.n227 CS_BIAS.n226 0.189894
R645 CS_BIAS.n226 CS_BIAS.n192 0.189894
R646 CS_BIAS.n221 CS_BIAS.n192 0.189894
R647 CS_BIAS.n221 CS_BIAS.n220 0.189894
R648 CS_BIAS.n220 CS_BIAS.n219 0.189894
R649 CS_BIAS.n219 CS_BIAS.n194 0.189894
R650 CS_BIAS.n214 CS_BIAS.n194 0.189894
R651 CS_BIAS.n214 CS_BIAS.n213 0.189894
R652 CS_BIAS.n213 CS_BIAS.n212 0.189894
R653 CS_BIAS.n212 CS_BIAS.n196 0.189894
R654 CS_BIAS.n207 CS_BIAS.n196 0.189894
R655 CS_BIAS.n207 CS_BIAS.n206 0.189894
R656 CS_BIAS.n206 CS_BIAS.n205 0.189894
R657 CS_BIAS.n205 CS_BIAS.n198 0.189894
R658 CS_BIAS.n201 CS_BIAS.n198 0.189894
R659 CS_BIAS.n93 CS_BIAS.n13 0.189894
R660 CS_BIAS.n93 CS_BIAS.n92 0.189894
R661 CS_BIAS.n92 CS_BIAS.n91 0.189894
R662 CS_BIAS.n91 CS_BIAS.n15 0.189894
R663 CS_BIAS.n86 CS_BIAS.n15 0.189894
R664 CS_BIAS.n86 CS_BIAS.n85 0.189894
R665 CS_BIAS.n85 CS_BIAS.n84 0.189894
R666 CS_BIAS.n84 CS_BIAS.n17 0.189894
R667 CS_BIAS.n79 CS_BIAS.n17 0.189894
R668 CS_BIAS.n79 CS_BIAS.n78 0.189894
R669 CS_BIAS.n78 CS_BIAS.n77 0.189894
R670 CS_BIAS.n77 CS_BIAS.n19 0.189894
R671 CS_BIAS.n73 CS_BIAS.n19 0.189894
R672 CS_BIAS.n73 CS_BIAS.n72 0.189894
R673 CS_BIAS.n72 CS_BIAS.n21 0.189894
R674 CS_BIAS.n68 CS_BIAS.n21 0.189894
R675 CS_BIAS.n68 CS_BIAS.n67 0.189894
R676 CS_BIAS.n67 CS_BIAS.n66 0.189894
R677 CS_BIAS.n66 CS_BIAS.n23 0.189894
R678 CS_BIAS.n62 CS_BIAS.n23 0.189894
R679 CS_BIAS.n62 CS_BIAS.n61 0.189894
R680 CS_BIAS.n61 CS_BIAS.n60 0.189894
R681 CS_BIAS.n60 CS_BIAS.n26 0.189894
R682 CS_BIAS.n55 CS_BIAS.n26 0.189894
R683 CS_BIAS.n55 CS_BIAS.n54 0.189894
R684 CS_BIAS.n54 CS_BIAS.n53 0.189894
R685 CS_BIAS.n53 CS_BIAS.n28 0.189894
R686 CS_BIAS.n48 CS_BIAS.n28 0.189894
R687 CS_BIAS.n48 CS_BIAS.n47 0.189894
R688 CS_BIAS.n47 CS_BIAS.n46 0.189894
R689 CS_BIAS.n46 CS_BIAS.n30 0.189894
R690 CS_BIAS.n41 CS_BIAS.n30 0.189894
R691 CS_BIAS.n41 CS_BIAS.n40 0.189894
R692 CS_BIAS.n40 CS_BIAS.n39 0.189894
R693 CS_BIAS.n39 CS_BIAS.n32 0.189894
R694 CS_BIAS.n35 CS_BIAS.n32 0.189894
R695 CS_BIAS.n142 CS_BIAS.n141 0.189894
R696 CS_BIAS.n141 CS_BIAS.n107 0.189894
R697 CS_BIAS.n136 CS_BIAS.n107 0.189894
R698 CS_BIAS.n136 CS_BIAS.n135 0.189894
R699 CS_BIAS.n135 CS_BIAS.n134 0.189894
R700 CS_BIAS.n134 CS_BIAS.n109 0.189894
R701 CS_BIAS.n129 CS_BIAS.n109 0.189894
R702 CS_BIAS.n129 CS_BIAS.n128 0.189894
R703 CS_BIAS.n128 CS_BIAS.n127 0.189894
R704 CS_BIAS.n127 CS_BIAS.n111 0.189894
R705 CS_BIAS.n122 CS_BIAS.n111 0.189894
R706 CS_BIAS.n122 CS_BIAS.n121 0.189894
R707 CS_BIAS.n121 CS_BIAS.n120 0.189894
R708 CS_BIAS.n120 CS_BIAS.n113 0.189894
R709 CS_BIAS.n116 CS_BIAS.n113 0.189894
R710 CS_BIAS.n174 CS_BIAS.n0 0.189894
R711 CS_BIAS.n174 CS_BIAS.n173 0.189894
R712 CS_BIAS.n173 CS_BIAS.n172 0.189894
R713 CS_BIAS.n172 CS_BIAS.n2 0.189894
R714 CS_BIAS.n167 CS_BIAS.n2 0.189894
R715 CS_BIAS.n167 CS_BIAS.n166 0.189894
R716 CS_BIAS.n166 CS_BIAS.n165 0.189894
R717 CS_BIAS.n165 CS_BIAS.n4 0.189894
R718 CS_BIAS.n160 CS_BIAS.n4 0.189894
R719 CS_BIAS.n160 CS_BIAS.n159 0.189894
R720 CS_BIAS.n159 CS_BIAS.n158 0.189894
R721 CS_BIAS.n158 CS_BIAS.n6 0.189894
R722 CS_BIAS.n154 CS_BIAS.n6 0.189894
R723 CS_BIAS.n154 CS_BIAS.n153 0.189894
R724 CS_BIAS.n153 CS_BIAS.n8 0.189894
R725 CS_BIAS.n149 CS_BIAS.n8 0.189894
R726 CS_BIAS.n149 CS_BIAS.n148 0.189894
R727 CS_BIAS.n148 CS_BIAS.n147 0.189894
R728 CS_BIAS.n147 CS_BIAS.n10 0.189894
R729 CS_BIAS.n465 CS_BIAS.n462 0.189894
R730 CS_BIAS.n469 CS_BIAS.n462 0.189894
R731 CS_BIAS.n470 CS_BIAS.n469 0.189894
R732 CS_BIAS.n471 CS_BIAS.n470 0.189894
R733 CS_BIAS.n471 CS_BIAS.n460 0.189894
R734 CS_BIAS.n476 CS_BIAS.n460 0.189894
R735 CS_BIAS.n477 CS_BIAS.n476 0.189894
R736 CS_BIAS.n478 CS_BIAS.n477 0.189894
R737 CS_BIAS.n478 CS_BIAS.n458 0.189894
R738 CS_BIAS.n483 CS_BIAS.n458 0.189894
R739 CS_BIAS.n484 CS_BIAS.n483 0.189894
R740 CS_BIAS.n485 CS_BIAS.n484 0.189894
R741 CS_BIAS.n485 CS_BIAS.n456 0.189894
R742 CS_BIAS.n490 CS_BIAS.n456 0.189894
R743 CS_BIAS.n491 CS_BIAS.n490 0.189894
R744 CS_BIAS.n492 CS_BIAS.n491 0.189894
R745 CS_BIAS.n492 CS_BIAS.n454 0.189894
R746 CS_BIAS.n497 CS_BIAS.n454 0.189894
R747 CS_BIAS.n498 CS_BIAS.n497 0.189894
R748 CS_BIAS.n499 CS_BIAS.n498 0.189894
R749 CS_BIAS.n499 CS_BIAS.n452 0.189894
R750 CS_BIAS.n503 CS_BIAS.n452 0.189894
R751 CS_BIAS.n504 CS_BIAS.n503 0.189894
R752 CS_BIAS.n504 CS_BIAS.n450 0.189894
R753 CS_BIAS.n508 CS_BIAS.n450 0.189894
R754 CS_BIAS.n509 CS_BIAS.n508 0.189894
R755 CS_BIAS.n510 CS_BIAS.n509 0.189894
R756 CS_BIAS.n510 CS_BIAS.n448 0.189894
R757 CS_BIAS.n515 CS_BIAS.n448 0.189894
R758 CS_BIAS.n516 CS_BIAS.n515 0.189894
R759 CS_BIAS.n517 CS_BIAS.n516 0.189894
R760 CS_BIAS.n517 CS_BIAS.n446 0.189894
R761 CS_BIAS.n522 CS_BIAS.n446 0.189894
R762 CS_BIAS.n523 CS_BIAS.n522 0.189894
R763 CS_BIAS.n524 CS_BIAS.n523 0.189894
R764 CS_BIAS.n524 CS_BIAS.n444 0.189894
R765 CS_BIAS.n338 CS_BIAS.n335 0.189894
R766 CS_BIAS.n342 CS_BIAS.n335 0.189894
R767 CS_BIAS.n343 CS_BIAS.n342 0.189894
R768 CS_BIAS.n344 CS_BIAS.n343 0.189894
R769 CS_BIAS.n344 CS_BIAS.n333 0.189894
R770 CS_BIAS.n349 CS_BIAS.n333 0.189894
R771 CS_BIAS.n350 CS_BIAS.n349 0.189894
R772 CS_BIAS.n351 CS_BIAS.n350 0.189894
R773 CS_BIAS.n351 CS_BIAS.n331 0.189894
R774 CS_BIAS.n356 CS_BIAS.n331 0.189894
R775 CS_BIAS.n357 CS_BIAS.n356 0.189894
R776 CS_BIAS.n358 CS_BIAS.n357 0.189894
R777 CS_BIAS.n358 CS_BIAS.n329 0.189894
R778 CS_BIAS.n363 CS_BIAS.n329 0.189894
R779 CS_BIAS.n364 CS_BIAS.n363 0.189894
R780 CS_BIAS.n365 CS_BIAS.n364 0.189894
R781 CS_BIAS.n365 CS_BIAS.n327 0.189894
R782 CS_BIAS.n370 CS_BIAS.n327 0.189894
R783 CS_BIAS.n371 CS_BIAS.n370 0.189894
R784 CS_BIAS.n372 CS_BIAS.n371 0.189894
R785 CS_BIAS.n372 CS_BIAS.n325 0.189894
R786 CS_BIAS.n376 CS_BIAS.n325 0.189894
R787 CS_BIAS.n377 CS_BIAS.n376 0.189894
R788 CS_BIAS.n377 CS_BIAS.n323 0.189894
R789 CS_BIAS.n381 CS_BIAS.n323 0.189894
R790 CS_BIAS.n382 CS_BIAS.n381 0.189894
R791 CS_BIAS.n383 CS_BIAS.n382 0.189894
R792 CS_BIAS.n383 CS_BIAS.n321 0.189894
R793 CS_BIAS.n388 CS_BIAS.n321 0.189894
R794 CS_BIAS.n389 CS_BIAS.n388 0.189894
R795 CS_BIAS.n390 CS_BIAS.n389 0.189894
R796 CS_BIAS.n390 CS_BIAS.n319 0.189894
R797 CS_BIAS.n395 CS_BIAS.n319 0.189894
R798 CS_BIAS.n396 CS_BIAS.n395 0.189894
R799 CS_BIAS.n397 CS_BIAS.n396 0.189894
R800 CS_BIAS.n397 CS_BIAS.n317 0.189894
R801 CS_BIAS.n286 CS_BIAS.n283 0.189894
R802 CS_BIAS.n290 CS_BIAS.n283 0.189894
R803 CS_BIAS.n291 CS_BIAS.n290 0.189894
R804 CS_BIAS.n292 CS_BIAS.n291 0.189894
R805 CS_BIAS.n292 CS_BIAS.n281 0.189894
R806 CS_BIAS.n297 CS_BIAS.n281 0.189894
R807 CS_BIAS.n298 CS_BIAS.n297 0.189894
R808 CS_BIAS.n299 CS_BIAS.n298 0.189894
R809 CS_BIAS.n299 CS_BIAS.n279 0.189894
R810 CS_BIAS.n304 CS_BIAS.n279 0.189894
R811 CS_BIAS.n305 CS_BIAS.n304 0.189894
R812 CS_BIAS.n306 CS_BIAS.n305 0.189894
R813 CS_BIAS.n306 CS_BIAS.n277 0.189894
R814 CS_BIAS.n311 CS_BIAS.n277 0.189894
R815 CS_BIAS.n312 CS_BIAS.n311 0.189894
R816 CS_BIAS.n412 CS_BIAS.n275 0.189894
R817 CS_BIAS.n413 CS_BIAS.n412 0.189894
R818 CS_BIAS.n414 CS_BIAS.n413 0.189894
R819 CS_BIAS.n414 CS_BIAS.n273 0.189894
R820 CS_BIAS.n418 CS_BIAS.n273 0.189894
R821 CS_BIAS.n419 CS_BIAS.n418 0.189894
R822 CS_BIAS.n419 CS_BIAS.n271 0.189894
R823 CS_BIAS.n423 CS_BIAS.n271 0.189894
R824 CS_BIAS.n424 CS_BIAS.n423 0.189894
R825 CS_BIAS.n425 CS_BIAS.n424 0.189894
R826 CS_BIAS.n425 CS_BIAS.n269 0.189894
R827 CS_BIAS.n430 CS_BIAS.n269 0.189894
R828 CS_BIAS.n431 CS_BIAS.n430 0.189894
R829 CS_BIAS.n432 CS_BIAS.n431 0.189894
R830 CS_BIAS.n432 CS_BIAS.n267 0.189894
R831 CS_BIAS.n437 CS_BIAS.n267 0.189894
R832 CS_BIAS.n438 CS_BIAS.n437 0.189894
R833 CS_BIAS.n439 CS_BIAS.n438 0.189894
R834 CS_BIAS.n439 CS_BIAS.n265 0.189894
R835 CS_BIAS.n143 CS_BIAS.n142 0.170955
R836 CS_BIAS.n143 CS_BIAS.n10 0.170955
R837 CS_BIAS.n407 CS_BIAS.n312 0.170955
R838 CS_BIAS.n407 CS_BIAS.n275 0.170955
R839 GND.n5482 GND.n5481 1600.64
R840 GND.n1696 GND.n1108 1156.7
R841 GND.n5834 GND.n468 800.013
R842 GND.n573 GND.n470 800.013
R843 GND.n2567 GND.n2483 800.013
R844 GND.n4406 GND.n2569 800.013
R845 GND.n1296 GND.n1239 800.013
R846 GND.n4653 GND.n1237 800.013
R847 GND.n1920 GND.n1695 800.013
R848 GND.n1831 GND.n1698 800.013
R849 GND.n5028 GND.n972 795.207
R850 GND.n5483 GND.n702 795.207
R851 GND.n5661 GND.n597 795.207
R852 GND.n4886 GND.n1109 795.207
R853 GND.n5832 GND.n472 780.793
R854 GND.n539 GND.n469 780.793
R855 GND.n4409 GND.n4408 780.793
R856 GND.n4481 GND.n2519 780.793
R857 GND.n4799 GND.n1241 780.793
R858 GND.n4801 GND.n1235 780.793
R859 GND.n1837 GND.n1697 780.793
R860 GND.n1918 GND.n1699 780.793
R861 GND.n4538 GND.n2431 766.379
R862 GND.n4540 GND.n2427 766.379
R863 GND.n2346 GND.n2345 766.379
R864 GND.n4701 GND.n1330 766.379
R865 GND.n5028 GND.n5027 585
R866 GND.n5029 GND.n5028 585
R867 GND.n5026 GND.n974 585
R868 GND.n974 GND.n973 585
R869 GND.n5025 GND.n5024 585
R870 GND.n5024 GND.n5023 585
R871 GND.n979 GND.n978 585
R872 GND.n5022 GND.n979 585
R873 GND.n5020 GND.n5019 585
R874 GND.n5021 GND.n5020 585
R875 GND.n5018 GND.n981 585
R876 GND.n981 GND.n980 585
R877 GND.n5017 GND.n5016 585
R878 GND.n5016 GND.n5015 585
R879 GND.n987 GND.n986 585
R880 GND.n5014 GND.n987 585
R881 GND.n5012 GND.n5011 585
R882 GND.n5013 GND.n5012 585
R883 GND.n5010 GND.n989 585
R884 GND.n989 GND.n988 585
R885 GND.n5009 GND.n5008 585
R886 GND.n5008 GND.n5007 585
R887 GND.n995 GND.n994 585
R888 GND.n5006 GND.n995 585
R889 GND.n5004 GND.n5003 585
R890 GND.n5005 GND.n5004 585
R891 GND.n5002 GND.n997 585
R892 GND.n997 GND.n996 585
R893 GND.n5001 GND.n5000 585
R894 GND.n5000 GND.n4999 585
R895 GND.n1003 GND.n1002 585
R896 GND.n4998 GND.n1003 585
R897 GND.n4996 GND.n4995 585
R898 GND.n4997 GND.n4996 585
R899 GND.n4994 GND.n1005 585
R900 GND.n1005 GND.n1004 585
R901 GND.n4993 GND.n4992 585
R902 GND.n4992 GND.n4991 585
R903 GND.n1011 GND.n1010 585
R904 GND.n4990 GND.n1011 585
R905 GND.n4988 GND.n4987 585
R906 GND.n4989 GND.n4988 585
R907 GND.n4986 GND.n1013 585
R908 GND.n1013 GND.n1012 585
R909 GND.n4985 GND.n4984 585
R910 GND.n4984 GND.n4983 585
R911 GND.n1019 GND.n1018 585
R912 GND.n4982 GND.n1019 585
R913 GND.n4980 GND.n4979 585
R914 GND.n4981 GND.n4980 585
R915 GND.n4978 GND.n1021 585
R916 GND.n1021 GND.n1020 585
R917 GND.n4977 GND.n4976 585
R918 GND.n4976 GND.n4975 585
R919 GND.n1027 GND.n1026 585
R920 GND.n4974 GND.n1027 585
R921 GND.n4972 GND.n4971 585
R922 GND.n4973 GND.n4972 585
R923 GND.n4970 GND.n1029 585
R924 GND.n1029 GND.n1028 585
R925 GND.n4969 GND.n4968 585
R926 GND.n4968 GND.n4967 585
R927 GND.n1035 GND.n1034 585
R928 GND.n4966 GND.n1035 585
R929 GND.n4964 GND.n4963 585
R930 GND.n4965 GND.n4964 585
R931 GND.n4962 GND.n1037 585
R932 GND.n1037 GND.n1036 585
R933 GND.n4961 GND.n4960 585
R934 GND.n4960 GND.n4959 585
R935 GND.n1043 GND.n1042 585
R936 GND.n4958 GND.n1043 585
R937 GND.n4956 GND.n4955 585
R938 GND.n4957 GND.n4956 585
R939 GND.n4954 GND.n1045 585
R940 GND.n1045 GND.n1044 585
R941 GND.n4953 GND.n4952 585
R942 GND.n4952 GND.n4951 585
R943 GND.n1051 GND.n1050 585
R944 GND.n4950 GND.n1051 585
R945 GND.n4948 GND.n4947 585
R946 GND.n4949 GND.n4948 585
R947 GND.n4946 GND.n1053 585
R948 GND.n1053 GND.n1052 585
R949 GND.n4945 GND.n4944 585
R950 GND.n4944 GND.n4943 585
R951 GND.n1059 GND.n1058 585
R952 GND.n4942 GND.n1059 585
R953 GND.n4940 GND.n4939 585
R954 GND.n4941 GND.n4940 585
R955 GND.n4938 GND.n1061 585
R956 GND.n1061 GND.n1060 585
R957 GND.n4937 GND.n4936 585
R958 GND.n4936 GND.n4935 585
R959 GND.n1067 GND.n1066 585
R960 GND.n4934 GND.n1067 585
R961 GND.n4932 GND.n4931 585
R962 GND.n4933 GND.n4932 585
R963 GND.n4930 GND.n1069 585
R964 GND.n1069 GND.n1068 585
R965 GND.n4929 GND.n4928 585
R966 GND.n4928 GND.n4927 585
R967 GND.n1075 GND.n1074 585
R968 GND.n4926 GND.n1075 585
R969 GND.n4924 GND.n4923 585
R970 GND.n4925 GND.n4924 585
R971 GND.n4922 GND.n1077 585
R972 GND.n1077 GND.n1076 585
R973 GND.n4921 GND.n4920 585
R974 GND.n4920 GND.n4919 585
R975 GND.n1083 GND.n1082 585
R976 GND.n4918 GND.n1083 585
R977 GND.n4916 GND.n4915 585
R978 GND.n4917 GND.n4916 585
R979 GND.n4914 GND.n1085 585
R980 GND.n1085 GND.n1084 585
R981 GND.n4913 GND.n4912 585
R982 GND.n4912 GND.n4911 585
R983 GND.n1091 GND.n1090 585
R984 GND.n4910 GND.n1091 585
R985 GND.n4908 GND.n4907 585
R986 GND.n4909 GND.n4908 585
R987 GND.n4906 GND.n1093 585
R988 GND.n1093 GND.n1092 585
R989 GND.n4905 GND.n4904 585
R990 GND.n4904 GND.n4903 585
R991 GND.n1099 GND.n1098 585
R992 GND.n4902 GND.n1099 585
R993 GND.n4900 GND.n4899 585
R994 GND.n4901 GND.n4900 585
R995 GND.n4898 GND.n1101 585
R996 GND.n1101 GND.n1100 585
R997 GND.n4897 GND.n4896 585
R998 GND.n4896 GND.n4895 585
R999 GND.n1107 GND.n1106 585
R1000 GND.n4894 GND.n1107 585
R1001 GND.n4892 GND.n4891 585
R1002 GND.n4893 GND.n4892 585
R1003 GND.n4890 GND.n1109 585
R1004 GND.n1109 GND.n1108 585
R1005 GND.n972 GND.n971 585
R1006 GND.n5030 GND.n972 585
R1007 GND.n5033 GND.n5032 585
R1008 GND.n5032 GND.n5031 585
R1009 GND.n969 GND.n968 585
R1010 GND.n968 GND.n967 585
R1011 GND.n5038 GND.n5037 585
R1012 GND.n5039 GND.n5038 585
R1013 GND.n966 GND.n965 585
R1014 GND.n5040 GND.n966 585
R1015 GND.n5043 GND.n5042 585
R1016 GND.n5042 GND.n5041 585
R1017 GND.n963 GND.n962 585
R1018 GND.n962 GND.n961 585
R1019 GND.n5048 GND.n5047 585
R1020 GND.n5049 GND.n5048 585
R1021 GND.n960 GND.n959 585
R1022 GND.n5050 GND.n960 585
R1023 GND.n5053 GND.n5052 585
R1024 GND.n5052 GND.n5051 585
R1025 GND.n957 GND.n956 585
R1026 GND.n956 GND.n955 585
R1027 GND.n5058 GND.n5057 585
R1028 GND.n5059 GND.n5058 585
R1029 GND.n954 GND.n953 585
R1030 GND.n5060 GND.n954 585
R1031 GND.n5063 GND.n5062 585
R1032 GND.n5062 GND.n5061 585
R1033 GND.n951 GND.n950 585
R1034 GND.n950 GND.n949 585
R1035 GND.n5068 GND.n5067 585
R1036 GND.n5069 GND.n5068 585
R1037 GND.n948 GND.n947 585
R1038 GND.n5070 GND.n948 585
R1039 GND.n5073 GND.n5072 585
R1040 GND.n5072 GND.n5071 585
R1041 GND.n945 GND.n944 585
R1042 GND.n944 GND.n943 585
R1043 GND.n5078 GND.n5077 585
R1044 GND.n5079 GND.n5078 585
R1045 GND.n942 GND.n941 585
R1046 GND.n5080 GND.n942 585
R1047 GND.n5083 GND.n5082 585
R1048 GND.n5082 GND.n5081 585
R1049 GND.n939 GND.n938 585
R1050 GND.n938 GND.n937 585
R1051 GND.n5088 GND.n5087 585
R1052 GND.n5089 GND.n5088 585
R1053 GND.n936 GND.n935 585
R1054 GND.n5090 GND.n936 585
R1055 GND.n5093 GND.n5092 585
R1056 GND.n5092 GND.n5091 585
R1057 GND.n933 GND.n932 585
R1058 GND.n932 GND.n931 585
R1059 GND.n5098 GND.n5097 585
R1060 GND.n5099 GND.n5098 585
R1061 GND.n930 GND.n929 585
R1062 GND.n5100 GND.n930 585
R1063 GND.n5103 GND.n5102 585
R1064 GND.n5102 GND.n5101 585
R1065 GND.n927 GND.n926 585
R1066 GND.n926 GND.n925 585
R1067 GND.n5108 GND.n5107 585
R1068 GND.n5109 GND.n5108 585
R1069 GND.n924 GND.n923 585
R1070 GND.n5110 GND.n924 585
R1071 GND.n5113 GND.n5112 585
R1072 GND.n5112 GND.n5111 585
R1073 GND.n921 GND.n920 585
R1074 GND.n920 GND.n919 585
R1075 GND.n5118 GND.n5117 585
R1076 GND.n5119 GND.n5118 585
R1077 GND.n918 GND.n917 585
R1078 GND.n5120 GND.n918 585
R1079 GND.n5123 GND.n5122 585
R1080 GND.n5122 GND.n5121 585
R1081 GND.n915 GND.n914 585
R1082 GND.n914 GND.n913 585
R1083 GND.n5128 GND.n5127 585
R1084 GND.n5129 GND.n5128 585
R1085 GND.n912 GND.n911 585
R1086 GND.n5130 GND.n912 585
R1087 GND.n5133 GND.n5132 585
R1088 GND.n5132 GND.n5131 585
R1089 GND.n909 GND.n908 585
R1090 GND.n908 GND.n907 585
R1091 GND.n5138 GND.n5137 585
R1092 GND.n5139 GND.n5138 585
R1093 GND.n906 GND.n905 585
R1094 GND.n5140 GND.n906 585
R1095 GND.n5143 GND.n5142 585
R1096 GND.n5142 GND.n5141 585
R1097 GND.n903 GND.n902 585
R1098 GND.n902 GND.n901 585
R1099 GND.n5148 GND.n5147 585
R1100 GND.n5149 GND.n5148 585
R1101 GND.n900 GND.n899 585
R1102 GND.n5150 GND.n900 585
R1103 GND.n5153 GND.n5152 585
R1104 GND.n5152 GND.n5151 585
R1105 GND.n897 GND.n896 585
R1106 GND.n896 GND.n895 585
R1107 GND.n5158 GND.n5157 585
R1108 GND.n5159 GND.n5158 585
R1109 GND.n894 GND.n893 585
R1110 GND.n5160 GND.n894 585
R1111 GND.n5163 GND.n5162 585
R1112 GND.n5162 GND.n5161 585
R1113 GND.n891 GND.n890 585
R1114 GND.n890 GND.n889 585
R1115 GND.n5168 GND.n5167 585
R1116 GND.n5169 GND.n5168 585
R1117 GND.n888 GND.n887 585
R1118 GND.n5170 GND.n888 585
R1119 GND.n5173 GND.n5172 585
R1120 GND.n5172 GND.n5171 585
R1121 GND.n885 GND.n884 585
R1122 GND.n884 GND.n883 585
R1123 GND.n5178 GND.n5177 585
R1124 GND.n5179 GND.n5178 585
R1125 GND.n882 GND.n881 585
R1126 GND.n5180 GND.n882 585
R1127 GND.n5183 GND.n5182 585
R1128 GND.n5182 GND.n5181 585
R1129 GND.n879 GND.n878 585
R1130 GND.n878 GND.n877 585
R1131 GND.n5188 GND.n5187 585
R1132 GND.n5189 GND.n5188 585
R1133 GND.n876 GND.n875 585
R1134 GND.n5190 GND.n876 585
R1135 GND.n5193 GND.n5192 585
R1136 GND.n5192 GND.n5191 585
R1137 GND.n873 GND.n872 585
R1138 GND.n872 GND.n871 585
R1139 GND.n5198 GND.n5197 585
R1140 GND.n5199 GND.n5198 585
R1141 GND.n870 GND.n869 585
R1142 GND.n5200 GND.n870 585
R1143 GND.n5203 GND.n5202 585
R1144 GND.n5202 GND.n5201 585
R1145 GND.n867 GND.n866 585
R1146 GND.n866 GND.n865 585
R1147 GND.n5208 GND.n5207 585
R1148 GND.n5209 GND.n5208 585
R1149 GND.n864 GND.n863 585
R1150 GND.n5210 GND.n864 585
R1151 GND.n5213 GND.n5212 585
R1152 GND.n5212 GND.n5211 585
R1153 GND.n861 GND.n860 585
R1154 GND.n860 GND.n859 585
R1155 GND.n5218 GND.n5217 585
R1156 GND.n5219 GND.n5218 585
R1157 GND.n858 GND.n857 585
R1158 GND.n5220 GND.n858 585
R1159 GND.n5223 GND.n5222 585
R1160 GND.n5222 GND.n5221 585
R1161 GND.n855 GND.n854 585
R1162 GND.n854 GND.n853 585
R1163 GND.n5228 GND.n5227 585
R1164 GND.n5229 GND.n5228 585
R1165 GND.n852 GND.n851 585
R1166 GND.n5230 GND.n852 585
R1167 GND.n5233 GND.n5232 585
R1168 GND.n5232 GND.n5231 585
R1169 GND.n849 GND.n848 585
R1170 GND.n848 GND.n847 585
R1171 GND.n5238 GND.n5237 585
R1172 GND.n5239 GND.n5238 585
R1173 GND.n846 GND.n845 585
R1174 GND.n5240 GND.n846 585
R1175 GND.n5243 GND.n5242 585
R1176 GND.n5242 GND.n5241 585
R1177 GND.n843 GND.n842 585
R1178 GND.n842 GND.n841 585
R1179 GND.n5248 GND.n5247 585
R1180 GND.n5249 GND.n5248 585
R1181 GND.n840 GND.n839 585
R1182 GND.n5250 GND.n840 585
R1183 GND.n5253 GND.n5252 585
R1184 GND.n5252 GND.n5251 585
R1185 GND.n837 GND.n836 585
R1186 GND.n836 GND.n835 585
R1187 GND.n5258 GND.n5257 585
R1188 GND.n5259 GND.n5258 585
R1189 GND.n834 GND.n833 585
R1190 GND.n5260 GND.n834 585
R1191 GND.n5263 GND.n5262 585
R1192 GND.n5262 GND.n5261 585
R1193 GND.n831 GND.n830 585
R1194 GND.n830 GND.n829 585
R1195 GND.n5268 GND.n5267 585
R1196 GND.n5269 GND.n5268 585
R1197 GND.n828 GND.n827 585
R1198 GND.n5270 GND.n828 585
R1199 GND.n5273 GND.n5272 585
R1200 GND.n5272 GND.n5271 585
R1201 GND.n825 GND.n824 585
R1202 GND.n824 GND.n823 585
R1203 GND.n5278 GND.n5277 585
R1204 GND.n5279 GND.n5278 585
R1205 GND.n822 GND.n821 585
R1206 GND.n5280 GND.n822 585
R1207 GND.n5283 GND.n5282 585
R1208 GND.n5282 GND.n5281 585
R1209 GND.n819 GND.n818 585
R1210 GND.n818 GND.n817 585
R1211 GND.n5288 GND.n5287 585
R1212 GND.n5289 GND.n5288 585
R1213 GND.n816 GND.n815 585
R1214 GND.n5290 GND.n816 585
R1215 GND.n5293 GND.n5292 585
R1216 GND.n5292 GND.n5291 585
R1217 GND.n813 GND.n812 585
R1218 GND.n812 GND.n811 585
R1219 GND.n5298 GND.n5297 585
R1220 GND.n5299 GND.n5298 585
R1221 GND.n810 GND.n809 585
R1222 GND.n5300 GND.n810 585
R1223 GND.n5303 GND.n5302 585
R1224 GND.n5302 GND.n5301 585
R1225 GND.n807 GND.n806 585
R1226 GND.n806 GND.n805 585
R1227 GND.n5308 GND.n5307 585
R1228 GND.n5309 GND.n5308 585
R1229 GND.n804 GND.n803 585
R1230 GND.n5310 GND.n804 585
R1231 GND.n5313 GND.n5312 585
R1232 GND.n5312 GND.n5311 585
R1233 GND.n801 GND.n800 585
R1234 GND.n800 GND.n799 585
R1235 GND.n5318 GND.n5317 585
R1236 GND.n5319 GND.n5318 585
R1237 GND.n798 GND.n797 585
R1238 GND.n5320 GND.n798 585
R1239 GND.n5323 GND.n5322 585
R1240 GND.n5322 GND.n5321 585
R1241 GND.n795 GND.n794 585
R1242 GND.n794 GND.n793 585
R1243 GND.n5328 GND.n5327 585
R1244 GND.n5329 GND.n5328 585
R1245 GND.n792 GND.n791 585
R1246 GND.n5330 GND.n792 585
R1247 GND.n5333 GND.n5332 585
R1248 GND.n5332 GND.n5331 585
R1249 GND.n789 GND.n788 585
R1250 GND.n788 GND.n787 585
R1251 GND.n5338 GND.n5337 585
R1252 GND.n5339 GND.n5338 585
R1253 GND.n786 GND.n785 585
R1254 GND.n5340 GND.n786 585
R1255 GND.n5343 GND.n5342 585
R1256 GND.n5342 GND.n5341 585
R1257 GND.n783 GND.n782 585
R1258 GND.n782 GND.n781 585
R1259 GND.n5348 GND.n5347 585
R1260 GND.n5349 GND.n5348 585
R1261 GND.n780 GND.n779 585
R1262 GND.n5350 GND.n780 585
R1263 GND.n5353 GND.n5352 585
R1264 GND.n5352 GND.n5351 585
R1265 GND.n777 GND.n776 585
R1266 GND.n776 GND.n775 585
R1267 GND.n5358 GND.n5357 585
R1268 GND.n5359 GND.n5358 585
R1269 GND.n774 GND.n773 585
R1270 GND.n5360 GND.n774 585
R1271 GND.n5363 GND.n5362 585
R1272 GND.n5362 GND.n5361 585
R1273 GND.n771 GND.n770 585
R1274 GND.n770 GND.n769 585
R1275 GND.n5368 GND.n5367 585
R1276 GND.n5369 GND.n5368 585
R1277 GND.n768 GND.n767 585
R1278 GND.n5370 GND.n768 585
R1279 GND.n5373 GND.n5372 585
R1280 GND.n5372 GND.n5371 585
R1281 GND.n765 GND.n764 585
R1282 GND.n764 GND.n763 585
R1283 GND.n5378 GND.n5377 585
R1284 GND.n5379 GND.n5378 585
R1285 GND.n762 GND.n761 585
R1286 GND.n5380 GND.n762 585
R1287 GND.n5383 GND.n5382 585
R1288 GND.n5382 GND.n5381 585
R1289 GND.n759 GND.n758 585
R1290 GND.n758 GND.n757 585
R1291 GND.n5388 GND.n5387 585
R1292 GND.n5389 GND.n5388 585
R1293 GND.n756 GND.n755 585
R1294 GND.n5390 GND.n756 585
R1295 GND.n5393 GND.n5392 585
R1296 GND.n5392 GND.n5391 585
R1297 GND.n753 GND.n752 585
R1298 GND.n752 GND.n751 585
R1299 GND.n5398 GND.n5397 585
R1300 GND.n5399 GND.n5398 585
R1301 GND.n750 GND.n749 585
R1302 GND.n5400 GND.n750 585
R1303 GND.n5403 GND.n5402 585
R1304 GND.n5402 GND.n5401 585
R1305 GND.n747 GND.n746 585
R1306 GND.n746 GND.n745 585
R1307 GND.n5408 GND.n5407 585
R1308 GND.n5409 GND.n5408 585
R1309 GND.n744 GND.n743 585
R1310 GND.n5410 GND.n744 585
R1311 GND.n5413 GND.n5412 585
R1312 GND.n5412 GND.n5411 585
R1313 GND.n741 GND.n740 585
R1314 GND.n740 GND.n739 585
R1315 GND.n5418 GND.n5417 585
R1316 GND.n5419 GND.n5418 585
R1317 GND.n738 GND.n737 585
R1318 GND.n5420 GND.n738 585
R1319 GND.n5423 GND.n5422 585
R1320 GND.n5422 GND.n5421 585
R1321 GND.n735 GND.n734 585
R1322 GND.n734 GND.n733 585
R1323 GND.n5428 GND.n5427 585
R1324 GND.n5429 GND.n5428 585
R1325 GND.n732 GND.n731 585
R1326 GND.n5430 GND.n732 585
R1327 GND.n5433 GND.n5432 585
R1328 GND.n5432 GND.n5431 585
R1329 GND.n729 GND.n728 585
R1330 GND.n728 GND.n727 585
R1331 GND.n5438 GND.n5437 585
R1332 GND.n5439 GND.n5438 585
R1333 GND.n726 GND.n725 585
R1334 GND.n5440 GND.n726 585
R1335 GND.n5443 GND.n5442 585
R1336 GND.n5442 GND.n5441 585
R1337 GND.n723 GND.n722 585
R1338 GND.n722 GND.n721 585
R1339 GND.n5448 GND.n5447 585
R1340 GND.n5449 GND.n5448 585
R1341 GND.n720 GND.n719 585
R1342 GND.n5450 GND.n720 585
R1343 GND.n5453 GND.n5452 585
R1344 GND.n5452 GND.n5451 585
R1345 GND.n717 GND.n716 585
R1346 GND.n716 GND.n715 585
R1347 GND.n5458 GND.n5457 585
R1348 GND.n5459 GND.n5458 585
R1349 GND.n714 GND.n713 585
R1350 GND.n5460 GND.n714 585
R1351 GND.n5463 GND.n5462 585
R1352 GND.n5462 GND.n5461 585
R1353 GND.n711 GND.n710 585
R1354 GND.n710 GND.n709 585
R1355 GND.n5468 GND.n5467 585
R1356 GND.n5469 GND.n5468 585
R1357 GND.n708 GND.n707 585
R1358 GND.n5470 GND.n708 585
R1359 GND.n5473 GND.n5472 585
R1360 GND.n5472 GND.n5471 585
R1361 GND.n705 GND.n704 585
R1362 GND.n704 GND.n703 585
R1363 GND.n5479 GND.n5478 585
R1364 GND.n5480 GND.n5479 585
R1365 GND.n5477 GND.n702 585
R1366 GND.n5481 GND.n702 585
R1367 GND.n5657 GND.n597 585
R1368 GND.n5653 GND.n597 585
R1369 GND.n5656 GND.n5655 585
R1370 GND.n5655 GND.n5654 585
R1371 GND.n601 GND.n600 585
R1372 GND.n5652 GND.n601 585
R1373 GND.n5650 GND.n5649 585
R1374 GND.n5651 GND.n5650 585
R1375 GND.n604 GND.n603 585
R1376 GND.n603 GND.n602 585
R1377 GND.n5644 GND.n5643 585
R1378 GND.n5643 GND.n5642 585
R1379 GND.n607 GND.n606 585
R1380 GND.n5641 GND.n607 585
R1381 GND.n5639 GND.n5638 585
R1382 GND.n5640 GND.n5639 585
R1383 GND.n610 GND.n609 585
R1384 GND.n609 GND.n608 585
R1385 GND.n5634 GND.n5633 585
R1386 GND.n5633 GND.n5632 585
R1387 GND.n613 GND.n612 585
R1388 GND.n5631 GND.n613 585
R1389 GND.n5629 GND.n5628 585
R1390 GND.n5630 GND.n5629 585
R1391 GND.n616 GND.n615 585
R1392 GND.n615 GND.n614 585
R1393 GND.n5624 GND.n5623 585
R1394 GND.n5623 GND.n5622 585
R1395 GND.n619 GND.n618 585
R1396 GND.n5621 GND.n619 585
R1397 GND.n5619 GND.n5618 585
R1398 GND.n5620 GND.n5619 585
R1399 GND.n622 GND.n621 585
R1400 GND.n621 GND.n620 585
R1401 GND.n5614 GND.n5613 585
R1402 GND.n5613 GND.n5612 585
R1403 GND.n625 GND.n624 585
R1404 GND.n5611 GND.n625 585
R1405 GND.n5609 GND.n5608 585
R1406 GND.n5610 GND.n5609 585
R1407 GND.n628 GND.n627 585
R1408 GND.n627 GND.n626 585
R1409 GND.n5604 GND.n5603 585
R1410 GND.n5603 GND.n5602 585
R1411 GND.n631 GND.n630 585
R1412 GND.n5601 GND.n631 585
R1413 GND.n5599 GND.n5598 585
R1414 GND.n5600 GND.n5599 585
R1415 GND.n634 GND.n633 585
R1416 GND.n633 GND.n632 585
R1417 GND.n5594 GND.n5593 585
R1418 GND.n5593 GND.n5592 585
R1419 GND.n637 GND.n636 585
R1420 GND.n5591 GND.n637 585
R1421 GND.n5589 GND.n5588 585
R1422 GND.n5590 GND.n5589 585
R1423 GND.n640 GND.n639 585
R1424 GND.n639 GND.n638 585
R1425 GND.n5584 GND.n5583 585
R1426 GND.n5583 GND.n5582 585
R1427 GND.n643 GND.n642 585
R1428 GND.n5581 GND.n643 585
R1429 GND.n5579 GND.n5578 585
R1430 GND.n5580 GND.n5579 585
R1431 GND.n646 GND.n645 585
R1432 GND.n645 GND.n644 585
R1433 GND.n5574 GND.n5573 585
R1434 GND.n5573 GND.n5572 585
R1435 GND.n649 GND.n648 585
R1436 GND.n5571 GND.n649 585
R1437 GND.n5569 GND.n5568 585
R1438 GND.n5570 GND.n5569 585
R1439 GND.n652 GND.n651 585
R1440 GND.n651 GND.n650 585
R1441 GND.n5564 GND.n5563 585
R1442 GND.n5563 GND.n5562 585
R1443 GND.n655 GND.n654 585
R1444 GND.n5561 GND.n655 585
R1445 GND.n5559 GND.n5558 585
R1446 GND.n5560 GND.n5559 585
R1447 GND.n658 GND.n657 585
R1448 GND.n657 GND.n656 585
R1449 GND.n5554 GND.n5553 585
R1450 GND.n5553 GND.n5552 585
R1451 GND.n661 GND.n660 585
R1452 GND.n5551 GND.n661 585
R1453 GND.n5549 GND.n5548 585
R1454 GND.n5550 GND.n5549 585
R1455 GND.n664 GND.n663 585
R1456 GND.n663 GND.n662 585
R1457 GND.n5544 GND.n5543 585
R1458 GND.n5543 GND.n5542 585
R1459 GND.n667 GND.n666 585
R1460 GND.n5541 GND.n667 585
R1461 GND.n5539 GND.n5538 585
R1462 GND.n5540 GND.n5539 585
R1463 GND.n670 GND.n669 585
R1464 GND.n669 GND.n668 585
R1465 GND.n5534 GND.n5533 585
R1466 GND.n5533 GND.n5532 585
R1467 GND.n673 GND.n672 585
R1468 GND.n5531 GND.n673 585
R1469 GND.n5529 GND.n5528 585
R1470 GND.n5530 GND.n5529 585
R1471 GND.n676 GND.n675 585
R1472 GND.n675 GND.n674 585
R1473 GND.n5524 GND.n5523 585
R1474 GND.n5523 GND.n5522 585
R1475 GND.n679 GND.n678 585
R1476 GND.n5521 GND.n679 585
R1477 GND.n5519 GND.n5518 585
R1478 GND.n5520 GND.n5519 585
R1479 GND.n682 GND.n681 585
R1480 GND.n681 GND.n680 585
R1481 GND.n5514 GND.n5513 585
R1482 GND.n5513 GND.n5512 585
R1483 GND.n685 GND.n684 585
R1484 GND.n5511 GND.n685 585
R1485 GND.n5509 GND.n5508 585
R1486 GND.n5510 GND.n5509 585
R1487 GND.n688 GND.n687 585
R1488 GND.n687 GND.n686 585
R1489 GND.n5504 GND.n5503 585
R1490 GND.n5503 GND.n5502 585
R1491 GND.n691 GND.n690 585
R1492 GND.n5501 GND.n691 585
R1493 GND.n5499 GND.n5498 585
R1494 GND.n5500 GND.n5499 585
R1495 GND.n694 GND.n693 585
R1496 GND.n693 GND.n692 585
R1497 GND.n5494 GND.n5493 585
R1498 GND.n5493 GND.n5492 585
R1499 GND.n697 GND.n696 585
R1500 GND.n5491 GND.n697 585
R1501 GND.n5489 GND.n5488 585
R1502 GND.n5490 GND.n5489 585
R1503 GND.n700 GND.n699 585
R1504 GND.n699 GND.n698 585
R1505 GND.n5484 GND.n5483 585
R1506 GND.n5483 GND.n5482 585
R1507 GND.n1239 GND.n1232 585
R1508 GND.n4800 GND.n1239 585
R1509 GND.n2328 GND.n1231 585
R1510 GND.n2329 GND.n2328 585
R1511 GND.n2327 GND.n1230 585
R1512 GND.n2327 GND.n2326 585
R1513 GND.n1404 GND.n1403 585
R1514 GND.n2307 GND.n1404 585
R1515 GND.n2317 GND.n1224 585
R1516 GND.n2318 GND.n2317 585
R1517 GND.n2316 GND.n1223 585
R1518 GND.n2316 GND.n2315 585
R1519 GND.n1413 GND.n1222 585
R1520 GND.n2286 GND.n1413 585
R1521 GND.n2276 GND.n2275 585
R1522 GND.n2276 GND.n1428 585
R1523 GND.n2277 GND.n1216 585
R1524 GND.n2278 GND.n2277 585
R1525 GND.n2274 GND.n1215 585
R1526 GND.n2274 GND.n2273 585
R1527 GND.n1437 GND.n1214 585
R1528 GND.n2170 GND.n1437 585
R1529 GND.n1448 GND.n1447 585
R1530 GND.n2261 GND.n1448 585
R1531 GND.n2249 GND.n1208 585
R1532 GND.n2249 GND.n2248 585
R1533 GND.n2250 GND.n1207 585
R1534 GND.n2251 GND.n2250 585
R1535 GND.n2247 GND.n1206 585
R1536 GND.n2247 GND.n2246 585
R1537 GND.n1460 GND.n1459 585
R1538 GND.n2151 GND.n1460 585
R1539 GND.n1469 GND.n1200 585
R1540 GND.n2237 GND.n1469 585
R1541 GND.n2225 GND.n1199 585
R1542 GND.n2225 GND.n2224 585
R1543 GND.n2226 GND.n1198 585
R1544 GND.n2227 GND.n2226 585
R1545 GND.n2222 GND.n1480 585
R1546 GND.n2222 GND.n2221 585
R1547 GND.n1479 GND.n1192 585
R1548 GND.n1493 GND.n1479 585
R1549 GND.n1491 GND.n1191 585
R1550 GND.n2212 GND.n1491 585
R1551 GND.n2199 GND.n1190 585
R1552 GND.n2199 GND.n2198 585
R1553 GND.n2201 GND.n2200 585
R1554 GND.n2202 GND.n2201 585
R1555 GND.n2197 GND.n1184 585
R1556 GND.n2197 GND.n2196 585
R1557 GND.n1501 GND.n1183 585
R1558 GND.n2100 GND.n1501 585
R1559 GND.n1554 GND.n1182 585
R1560 GND.n1557 GND.n1554 585
R1561 GND.n2108 GND.n1555 585
R1562 GND.n2108 GND.n2107 585
R1563 GND.n2109 GND.n1176 585
R1564 GND.n2110 GND.n2109 585
R1565 GND.n1553 GND.n1175 585
R1566 GND.n1571 GND.n1553 585
R1567 GND.n1544 GND.n1174 585
R1568 GND.n2117 GND.n1544 585
R1569 GND.n1533 GND.n1532 585
R1570 GND.n1536 GND.n1533 585
R1571 GND.n2125 GND.n1168 585
R1572 GND.n2125 GND.n2124 585
R1573 GND.n2126 GND.n1167 585
R1574 GND.n2127 GND.n2126 585
R1575 GND.n1531 GND.n1166 585
R1576 GND.n1574 GND.n1531 585
R1577 GND.n1522 GND.n1521 585
R1578 GND.n2134 GND.n1522 585
R1579 GND.n1582 GND.n1160 585
R1580 GND.n1582 GND.n1518 585
R1581 GND.n1583 GND.n1159 585
R1582 GND.n2067 GND.n1583 585
R1583 GND.n2055 GND.n1158 585
R1584 GND.n2055 GND.n2054 585
R1585 GND.n2057 GND.n2056 585
R1586 GND.n2058 GND.n2057 585
R1587 GND.n1592 GND.n1152 585
R1588 GND.n2043 GND.n1592 585
R1589 GND.n1607 GND.n1151 585
R1590 GND.n1607 GND.n1599 585
R1591 GND.n1608 GND.n1150 585
R1592 GND.n2031 GND.n1608 585
R1593 GND.n2019 GND.n1619 585
R1594 GND.n2019 GND.n2018 585
R1595 GND.n2020 GND.n1144 585
R1596 GND.n2021 GND.n2020 585
R1597 GND.n1618 GND.n1143 585
R1598 GND.n2005 GND.n1618 585
R1599 GND.n1633 GND.n1142 585
R1600 GND.n1638 GND.n1633 585
R1601 GND.n1135 GND.n1133 585
R1602 GND.n1996 GND.n1133 585
R1603 GND.n4877 GND.n4876 585
R1604 GND.n4878 GND.n4877 585
R1605 GND.n1134 GND.n1132 585
R1606 GND.n1646 GND.n1132 585
R1607 GND.n1966 GND.n1119 585
R1608 GND.n4884 GND.n1119 585
R1609 GND.n1965 GND.n1964 585
R1610 GND.n1964 GND.n1115 585
R1611 GND.n1963 GND.n1653 585
R1612 GND.n1986 GND.n1653 585
R1613 GND.n1665 GND.n1663 585
R1614 GND.n1663 GND.n1651 585
R1615 GND.n1976 GND.n1975 585
R1616 GND.n1977 GND.n1976 585
R1617 GND.n1664 GND.n1662 585
R1618 GND.n1662 GND.n1659 585
R1619 GND.n1685 GND.n1672 585
R1620 GND.n1956 GND.n1672 585
R1621 GND.n1683 GND.n1681 585
R1622 GND.n1681 GND.n1670 585
R1623 GND.n1947 GND.n1946 585
R1624 GND.n1948 GND.n1947 585
R1625 GND.n1682 GND.n1680 585
R1626 GND.n1940 GND.n1680 585
R1627 GND.n1764 GND.n1763 585
R1628 GND.n1763 GND.n1690 585
R1629 GND.n1762 GND.n1698 585
R1630 GND.n1919 GND.n1698 585
R1631 GND.n1832 GND.n1831 585
R1632 GND.n1829 GND.n1769 585
R1633 GND.n1828 GND.n1827 585
R1634 GND.n1773 GND.n1771 585
R1635 GND.n1823 GND.n1774 585
R1636 GND.n1822 GND.n1776 585
R1637 GND.n1821 GND.n1777 585
R1638 GND.n1781 GND.n1778 585
R1639 GND.n1817 GND.n1782 585
R1640 GND.n1816 GND.n1784 585
R1641 GND.n1815 GND.n1785 585
R1642 GND.n1789 GND.n1786 585
R1643 GND.n1811 GND.n1790 585
R1644 GND.n1810 GND.n1792 585
R1645 GND.n1809 GND.n1793 585
R1646 GND.n1797 GND.n1794 585
R1647 GND.n1805 GND.n1798 585
R1648 GND.n1804 GND.n1801 585
R1649 GND.n1799 GND.n1695 585
R1650 GND.n1696 GND.n1695 585
R1651 GND.n4654 GND.n4653 585
R1652 GND.n4655 GND.n1390 585
R1653 GND.n4656 GND.n1386 585
R1654 GND.n1378 GND.n1377 585
R1655 GND.n4663 GND.n1376 585
R1656 GND.n4664 GND.n1375 585
R1657 GND.n1374 GND.n1368 585
R1658 GND.n4671 GND.n1367 585
R1659 GND.n4672 GND.n1366 585
R1660 GND.n1358 GND.n1357 585
R1661 GND.n4679 GND.n1356 585
R1662 GND.n4680 GND.n1355 585
R1663 GND.n1354 GND.n1348 585
R1664 GND.n4687 GND.n1347 585
R1665 GND.n4688 GND.n1346 585
R1666 GND.n1339 GND.n1338 585
R1667 GND.n4695 GND.n1337 585
R1668 GND.n4696 GND.n1336 585
R1669 GND.n1335 GND.n1296 585
R1670 GND.n4737 GND.n1296 585
R1671 GND.n2332 GND.n1237 585
R1672 GND.n4800 GND.n1237 585
R1673 GND.n2331 GND.n2330 585
R1674 GND.n2330 GND.n2329 585
R1675 GND.n1401 GND.n1400 585
R1676 GND.n2326 GND.n1401 585
R1677 GND.n2309 GND.n2308 585
R1678 GND.n2308 GND.n2307 585
R1679 GND.n1418 GND.n1411 585
R1680 GND.n2318 GND.n1411 585
R1681 GND.n2314 GND.n2313 585
R1682 GND.n2315 GND.n2314 585
R1683 GND.n1417 GND.n1416 585
R1684 GND.n2286 GND.n1416 585
R1685 GND.n2267 GND.n2266 585
R1686 GND.n2266 GND.n1428 585
R1687 GND.n1441 GND.n1435 585
R1688 GND.n2278 GND.n1435 585
R1689 GND.n2272 GND.n2271 585
R1690 GND.n2273 GND.n2272 585
R1691 GND.n1440 GND.n1439 585
R1692 GND.n2170 GND.n1439 585
R1693 GND.n2263 GND.n2262 585
R1694 GND.n2262 GND.n2261 585
R1695 GND.n1444 GND.n1443 585
R1696 GND.n2248 GND.n1444 585
R1697 GND.n1463 GND.n1457 585
R1698 GND.n2251 GND.n1457 585
R1699 GND.n2245 GND.n2244 585
R1700 GND.n2246 GND.n2245 585
R1701 GND.n1462 GND.n1461 585
R1702 GND.n2151 GND.n1461 585
R1703 GND.n2239 GND.n2238 585
R1704 GND.n2238 GND.n2237 585
R1705 GND.n1466 GND.n1465 585
R1706 GND.n2224 GND.n1466 585
R1707 GND.n1484 GND.n1477 585
R1708 GND.n2227 GND.n1477 585
R1709 GND.n2220 GND.n2219 585
R1710 GND.n2221 GND.n2220 585
R1711 GND.n1483 GND.n1482 585
R1712 GND.n1493 GND.n1482 585
R1713 GND.n2214 GND.n2213 585
R1714 GND.n2213 GND.n2212 585
R1715 GND.n1487 GND.n1486 585
R1716 GND.n2198 GND.n1487 585
R1717 GND.n2088 GND.n1499 585
R1718 GND.n2202 GND.n1499 585
R1719 GND.n1563 GND.n1503 585
R1720 GND.n2196 GND.n1503 585
R1721 GND.n2093 GND.n2092 585
R1722 GND.n2100 GND.n2093 585
R1723 GND.n1562 GND.n1561 585
R1724 GND.n1561 GND.n1557 585
R1725 GND.n2085 GND.n1556 585
R1726 GND.n2107 GND.n1556 585
R1727 GND.n2084 GND.n1551 585
R1728 GND.n2110 GND.n1551 585
R1729 GND.n2083 GND.n1572 585
R1730 GND.n1572 GND.n1571 585
R1731 GND.n1565 GND.n1542 585
R1732 GND.n2117 GND.n1542 585
R1733 GND.n2078 GND.n2077 585
R1734 GND.n2077 GND.n1536 585
R1735 GND.n2076 GND.n1535 585
R1736 GND.n2124 GND.n1535 585
R1737 GND.n2075 GND.n1530 585
R1738 GND.n2127 GND.n1530 585
R1739 GND.n1576 GND.n1575 585
R1740 GND.n1575 GND.n1574 585
R1741 GND.n2071 GND.n1519 585
R1742 GND.n2134 GND.n1519 585
R1743 GND.n2070 GND.n2069 585
R1744 GND.n2069 GND.n1518 585
R1745 GND.n2068 GND.n1578 585
R1746 GND.n2068 GND.n2067 585
R1747 GND.n2037 GND.n1579 585
R1748 GND.n2054 GND.n1579 585
R1749 GND.n1602 GND.n1590 585
R1750 GND.n2058 GND.n1590 585
R1751 GND.n2042 GND.n2041 585
R1752 GND.n2043 GND.n2042 585
R1753 GND.n1601 GND.n1600 585
R1754 GND.n1600 GND.n1599 585
R1755 GND.n2033 GND.n2032 585
R1756 GND.n2032 GND.n2031 585
R1757 GND.n1605 GND.n1604 585
R1758 GND.n2018 GND.n1605 585
R1759 GND.n1642 GND.n1616 585
R1760 GND.n2021 GND.n1616 585
R1761 GND.n2004 GND.n2003 585
R1762 GND.n2005 GND.n2004 585
R1763 GND.n1641 GND.n1640 585
R1764 GND.n1640 GND.n1638 585
R1765 GND.n1998 GND.n1997 585
R1766 GND.n1997 GND.n1996 585
R1767 GND.n1994 GND.n1130 585
R1768 GND.n4878 GND.n1130 585
R1769 GND.n1993 GND.n1647 585
R1770 GND.n1647 GND.n1646 585
R1771 GND.n1644 GND.n1117 585
R1772 GND.n4884 GND.n1117 585
R1773 GND.n1989 GND.n1988 585
R1774 GND.n1988 GND.n1115 585
R1775 GND.n1987 GND.n1649 585
R1776 GND.n1987 GND.n1986 585
R1777 GND.n1928 GND.n1650 585
R1778 GND.n1651 GND.n1650 585
R1779 GND.n1927 GND.n1661 585
R1780 GND.n1977 GND.n1661 585
R1781 GND.n1932 GND.n1926 585
R1782 GND.n1926 GND.n1659 585
R1783 GND.n1933 GND.n1671 585
R1784 GND.n1956 GND.n1671 585
R1785 GND.n1934 GND.n1925 585
R1786 GND.n1925 GND.n1670 585
R1787 GND.n1693 GND.n1679 585
R1788 GND.n1948 GND.n1679 585
R1789 GND.n1939 GND.n1938 585
R1790 GND.n1940 GND.n1939 585
R1791 GND.n1692 GND.n1691 585
R1792 GND.n1691 GND.n1690 585
R1793 GND.n1921 GND.n1920 585
R1794 GND.n1920 GND.n1919 585
R1795 GND.n5835 GND.n5834 585
R1796 GND.n5834 GND.n5833 585
R1797 GND.n5836 GND.n464 585
R1798 GND.n464 GND.n463 585
R1799 GND.n5838 GND.n5837 585
R1800 GND.n5839 GND.n5838 585
R1801 GND.n450 GND.n449 585
R1802 GND.n453 GND.n450 585
R1803 GND.n5847 GND.n5846 585
R1804 GND.n5846 GND.n5845 585
R1805 GND.n5848 GND.n445 585
R1806 GND.n445 GND.n444 585
R1807 GND.n5850 GND.n5849 585
R1808 GND.n5851 GND.n5850 585
R1809 GND.n430 GND.n429 585
R1810 GND.n434 GND.n430 585
R1811 GND.n5859 GND.n5858 585
R1812 GND.n5858 GND.n5857 585
R1813 GND.n5860 GND.n425 585
R1814 GND.n431 GND.n425 585
R1815 GND.n5862 GND.n5861 585
R1816 GND.n5863 GND.n5862 585
R1817 GND.n410 GND.n409 585
R1818 GND.n5693 GND.n410 585
R1819 GND.n5871 GND.n5870 585
R1820 GND.n5870 GND.n5869 585
R1821 GND.n5872 GND.n405 585
R1822 GND.n5699 GND.n405 585
R1823 GND.n5874 GND.n5873 585
R1824 GND.n5875 GND.n5874 585
R1825 GND.n390 GND.n389 585
R1826 GND.n5669 GND.n390 585
R1827 GND.n5883 GND.n5882 585
R1828 GND.n5882 GND.n5881 585
R1829 GND.n5884 GND.n385 585
R1830 GND.n4251 GND.n385 585
R1831 GND.n5886 GND.n5885 585
R1832 GND.n5887 GND.n5886 585
R1833 GND.n369 GND.n368 585
R1834 GND.n4257 GND.n369 585
R1835 GND.n5895 GND.n5894 585
R1836 GND.n5894 GND.n5893 585
R1837 GND.n5896 GND.n364 585
R1838 GND.n4263 GND.n364 585
R1839 GND.n5898 GND.n5897 585
R1840 GND.n5899 GND.n5898 585
R1841 GND.n350 GND.n349 585
R1842 GND.n4269 GND.n350 585
R1843 GND.n5907 GND.n5906 585
R1844 GND.n5906 GND.n5905 585
R1845 GND.n5908 GND.n344 585
R1846 GND.n4231 GND.n344 585
R1847 GND.n5910 GND.n5909 585
R1848 GND.n5911 GND.n5910 585
R1849 GND.n345 GND.n343 585
R1850 GND.n4222 GND.n343 585
R1851 GND.n2732 GND.n2731 585
R1852 GND.n2754 GND.n2732 585
R1853 GND.n4310 GND.n4309 585
R1854 GND.n4309 GND.n4308 585
R1855 GND.n4311 GND.n323 585
R1856 GND.n5918 GND.n323 585
R1857 GND.n4313 GND.n4312 585
R1858 GND.n4314 GND.n4313 585
R1859 GND.n2727 GND.n2726 585
R1860 GND.n2726 GND.n2724 585
R1861 GND.n4208 GND.n4207 585
R1862 GND.n4207 GND.n2715 585
R1863 GND.n2706 GND.n2705 585
R1864 GND.n4323 GND.n2706 585
R1865 GND.n4329 GND.n4328 585
R1866 GND.n4328 GND.n4327 585
R1867 GND.n4330 GND.n2701 585
R1868 GND.n4201 GND.n2701 585
R1869 GND.n4332 GND.n4331 585
R1870 GND.n4333 GND.n4332 585
R1871 GND.n2685 GND.n2684 585
R1872 GND.n4183 GND.n2685 585
R1873 GND.n4341 GND.n4340 585
R1874 GND.n4340 GND.n4339 585
R1875 GND.n4342 GND.n2680 585
R1876 GND.n4176 GND.n2680 585
R1877 GND.n4344 GND.n4343 585
R1878 GND.n4345 GND.n4344 585
R1879 GND.n2664 GND.n2663 585
R1880 GND.n4168 GND.n2664 585
R1881 GND.n4353 GND.n4352 585
R1882 GND.n4352 GND.n4351 585
R1883 GND.n4354 GND.n2659 585
R1884 GND.n4161 GND.n2659 585
R1885 GND.n4356 GND.n4355 585
R1886 GND.n4357 GND.n4356 585
R1887 GND.n2644 GND.n2643 585
R1888 GND.n4153 GND.n2644 585
R1889 GND.n4365 GND.n4364 585
R1890 GND.n4364 GND.n4363 585
R1891 GND.n4366 GND.n2639 585
R1892 GND.n4146 GND.n2639 585
R1893 GND.n4368 GND.n4367 585
R1894 GND.n4369 GND.n4368 585
R1895 GND.n2623 GND.n2622 585
R1896 GND.n4138 GND.n2623 585
R1897 GND.n4377 GND.n4376 585
R1898 GND.n4376 GND.n4375 585
R1899 GND.n4378 GND.n2618 585
R1900 GND.n4131 GND.n2618 585
R1901 GND.n4380 GND.n4379 585
R1902 GND.n4381 GND.n4380 585
R1903 GND.n2602 GND.n2601 585
R1904 GND.n4123 GND.n2602 585
R1905 GND.n4389 GND.n4388 585
R1906 GND.n4388 GND.n4387 585
R1907 GND.n4390 GND.n2595 585
R1908 GND.n4116 GND.n2595 585
R1909 GND.n4392 GND.n4391 585
R1910 GND.n4393 GND.n4392 585
R1911 GND.n2596 GND.n2594 585
R1912 GND.n4108 GND.n2594 585
R1913 GND.n2578 GND.n2572 585
R1914 GND.n4399 GND.n2578 585
R1915 GND.n4404 GND.n2570 585
R1916 GND.n3988 GND.n2570 585
R1917 GND.n4406 GND.n4405 585
R1918 GND.n4407 GND.n4406 585
R1919 GND.n2569 GND.n2439 585
R1920 GND.n4529 GND.n2440 585
R1921 GND.n4528 GND.n2441 585
R1922 GND.n2504 GND.n2442 585
R1923 GND.n4521 GND.n2448 585
R1924 GND.n4520 GND.n2449 585
R1925 GND.n2507 GND.n2450 585
R1926 GND.n4513 GND.n2456 585
R1927 GND.n4512 GND.n2457 585
R1928 GND.n2509 GND.n2458 585
R1929 GND.n4505 GND.n2464 585
R1930 GND.n4504 GND.n2465 585
R1931 GND.n2512 GND.n2466 585
R1932 GND.n4497 GND.n2472 585
R1933 GND.n4496 GND.n2473 585
R1934 GND.n2514 GND.n2474 585
R1935 GND.n4489 GND.n2480 585
R1936 GND.n4488 GND.n4485 585
R1937 GND.n2483 GND.n2481 585
R1938 GND.n4483 GND.n2483 585
R1939 GND.n574 GND.n573 585
R1940 GND.n5727 GND.n569 585
R1941 GND.n5729 GND.n5728 585
R1942 GND.n5731 GND.n567 585
R1943 GND.n5733 GND.n5732 585
R1944 GND.n5734 GND.n562 585
R1945 GND.n5736 GND.n5735 585
R1946 GND.n5738 GND.n560 585
R1947 GND.n5740 GND.n5739 585
R1948 GND.n5741 GND.n555 585
R1949 GND.n5743 GND.n5742 585
R1950 GND.n5745 GND.n553 585
R1951 GND.n5747 GND.n5746 585
R1952 GND.n5748 GND.n548 585
R1953 GND.n5750 GND.n5749 585
R1954 GND.n5752 GND.n546 585
R1955 GND.n5754 GND.n5753 585
R1956 GND.n5755 GND.n544 585
R1957 GND.n5756 GND.n468 585
R1958 GND.n471 GND.n468 585
R1959 GND.n5723 GND.n470 585
R1960 GND.n5833 GND.n470 585
R1961 GND.n5722 GND.n5721 585
R1962 GND.n5721 GND.n463 585
R1963 GND.n5720 GND.n462 585
R1964 GND.n5839 GND.n462 585
R1965 GND.n579 GND.n578 585
R1966 GND.n578 GND.n453 585
R1967 GND.n5716 GND.n452 585
R1968 GND.n5845 GND.n452 585
R1969 GND.n5715 GND.n5714 585
R1970 GND.n5714 GND.n444 585
R1971 GND.n5713 GND.n443 585
R1972 GND.n5851 GND.n443 585
R1973 GND.n582 GND.n581 585
R1974 GND.n581 GND.n434 585
R1975 GND.n5709 GND.n433 585
R1976 GND.n5857 GND.n433 585
R1977 GND.n5708 GND.n5707 585
R1978 GND.n5707 GND.n431 585
R1979 GND.n5706 GND.n424 585
R1980 GND.n5863 GND.n424 585
R1981 GND.n5692 GND.n584 585
R1982 GND.n5693 GND.n5692 585
R1983 GND.n5702 GND.n413 585
R1984 GND.n5869 GND.n413 585
R1985 GND.n5701 GND.n5700 585
R1986 GND.n5700 GND.n5699 585
R1987 GND.n586 GND.n403 585
R1988 GND.n5875 GND.n403 585
R1989 GND.n4247 GND.n589 585
R1990 GND.n5669 GND.n589 585
R1991 GND.n4248 GND.n393 585
R1992 GND.n5881 GND.n393 585
R1993 GND.n4253 GND.n4252 585
R1994 GND.n4252 GND.n4251 585
R1995 GND.n4254 GND.n383 585
R1996 GND.n5887 GND.n383 585
R1997 GND.n4256 GND.n4255 585
R1998 GND.n4257 GND.n4256 585
R1999 GND.n2745 GND.n372 585
R2000 GND.n5893 GND.n372 585
R2001 GND.n4265 GND.n4264 585
R2002 GND.n4264 GND.n4263 585
R2003 GND.n4266 GND.n362 585
R2004 GND.n5899 GND.n362 585
R2005 GND.n4268 GND.n4267 585
R2006 GND.n4269 GND.n4268 585
R2007 GND.n2741 GND.n353 585
R2008 GND.n5905 GND.n353 585
R2009 GND.n4230 GND.n4229 585
R2010 GND.n4231 GND.n4230 585
R2011 GND.n2747 GND.n341 585
R2012 GND.n5911 GND.n341 585
R2013 GND.n4224 GND.n4223 585
R2014 GND.n4223 GND.n4222 585
R2015 GND.n2750 GND.n2749 585
R2016 GND.n2754 GND.n2750 585
R2017 GND.n319 GND.n317 585
R2018 GND.n4308 GND.n319 585
R2019 GND.n5920 GND.n5919 585
R2020 GND.n5919 GND.n5918 585
R2021 GND.n318 GND.n316 585
R2022 GND.n4314 GND.n318 585
R2023 GND.n4194 GND.n4193 585
R2024 GND.n4194 GND.n2724 585
R2025 GND.n4196 GND.n4195 585
R2026 GND.n4195 GND.n2715 585
R2027 GND.n4197 GND.n2714 585
R2028 GND.n4323 GND.n2714 585
R2029 GND.n4198 GND.n2709 585
R2030 GND.n4327 GND.n2709 585
R2031 GND.n4200 GND.n4199 585
R2032 GND.n4201 GND.n4200 585
R2033 GND.n2758 GND.n2699 585
R2034 GND.n4333 GND.n2699 585
R2035 GND.n4185 GND.n4184 585
R2036 GND.n4184 GND.n4183 585
R2037 GND.n2760 GND.n2688 585
R2038 GND.n4339 GND.n2688 585
R2039 GND.n4175 GND.n4174 585
R2040 GND.n4176 GND.n4175 585
R2041 GND.n2762 GND.n2678 585
R2042 GND.n4345 GND.n2678 585
R2043 GND.n4170 GND.n4169 585
R2044 GND.n4169 GND.n4168 585
R2045 GND.n2764 GND.n2667 585
R2046 GND.n4351 GND.n2667 585
R2047 GND.n4160 GND.n4159 585
R2048 GND.n4161 GND.n4160 585
R2049 GND.n2766 GND.n2657 585
R2050 GND.n4357 GND.n2657 585
R2051 GND.n4155 GND.n4154 585
R2052 GND.n4154 GND.n4153 585
R2053 GND.n2768 GND.n2647 585
R2054 GND.n4363 GND.n2647 585
R2055 GND.n4145 GND.n4144 585
R2056 GND.n4146 GND.n4145 585
R2057 GND.n2771 GND.n2637 585
R2058 GND.n4369 GND.n2637 585
R2059 GND.n4140 GND.n4139 585
R2060 GND.n4139 GND.n4138 585
R2061 GND.n2773 GND.n2626 585
R2062 GND.n4375 GND.n2626 585
R2063 GND.n4130 GND.n4129 585
R2064 GND.n4131 GND.n4130 585
R2065 GND.n2775 GND.n2616 585
R2066 GND.n4381 GND.n2616 585
R2067 GND.n4125 GND.n4124 585
R2068 GND.n4124 GND.n4123 585
R2069 GND.n2777 GND.n2605 585
R2070 GND.n4387 GND.n2605 585
R2071 GND.n4115 GND.n4114 585
R2072 GND.n4116 GND.n4115 585
R2073 GND.n2779 GND.n2592 585
R2074 GND.n4393 GND.n2592 585
R2075 GND.n4110 GND.n4109 585
R2076 GND.n4109 GND.n4108 585
R2077 GND.n2781 GND.n2577 585
R2078 GND.n4399 GND.n2577 585
R2079 GND.n3990 GND.n3989 585
R2080 GND.n3989 GND.n3988 585
R2081 GND.n3991 GND.n2567 585
R2082 GND.n4407 GND.n2567 585
R2083 GND.n4799 GND.n4798 585
R2084 GND.n4800 GND.n4799 585
R2085 GND.n1242 GND.n1240 585
R2086 GND.n2329 GND.n1240 585
R2087 GND.n2325 GND.n2324 585
R2088 GND.n2326 GND.n2325 585
R2089 GND.n1406 GND.n1405 585
R2090 GND.n2307 GND.n1405 585
R2091 GND.n2320 GND.n2319 585
R2092 GND.n2319 GND.n2318 585
R2093 GND.n1409 GND.n1408 585
R2094 GND.n2315 GND.n1409 585
R2095 GND.n2285 GND.n2284 585
R2096 GND.n2286 GND.n2285 585
R2097 GND.n1430 GND.n1429 585
R2098 GND.n1429 GND.n1428 585
R2099 GND.n2280 GND.n2279 585
R2100 GND.n2279 GND.n2278 585
R2101 GND.n1433 GND.n1432 585
R2102 GND.n2273 GND.n1433 585
R2103 GND.n2258 GND.n1450 585
R2104 GND.n2170 GND.n1450 585
R2105 GND.n2260 GND.n2259 585
R2106 GND.n2261 GND.n2260 585
R2107 GND.n1451 GND.n1449 585
R2108 GND.n2248 GND.n1449 585
R2109 GND.n2253 GND.n2252 585
R2110 GND.n2252 GND.n2251 585
R2111 GND.n1454 GND.n1453 585
R2112 GND.n2246 GND.n1454 585
R2113 GND.n2234 GND.n1471 585
R2114 GND.n2151 GND.n1471 585
R2115 GND.n2236 GND.n2235 585
R2116 GND.n2237 GND.n2236 585
R2117 GND.n1472 GND.n1470 585
R2118 GND.n2224 GND.n1470 585
R2119 GND.n2229 GND.n2228 585
R2120 GND.n2228 GND.n2227 585
R2121 GND.n1475 GND.n1474 585
R2122 GND.n2221 GND.n1475 585
R2123 GND.n2209 GND.n1494 585
R2124 GND.n1494 GND.n1493 585
R2125 GND.n2211 GND.n2210 585
R2126 GND.n2212 GND.n2211 585
R2127 GND.n1495 GND.n1492 585
R2128 GND.n2198 GND.n1492 585
R2129 GND.n2204 GND.n2203 585
R2130 GND.n2203 GND.n2202 585
R2131 GND.n1498 GND.n1497 585
R2132 GND.n2196 GND.n1498 585
R2133 GND.n2099 GND.n2098 585
R2134 GND.n2100 GND.n2099 585
R2135 GND.n2096 GND.n2094 585
R2136 GND.n2094 GND.n1557 585
R2137 GND.n2095 GND.n1550 585
R2138 GND.n2107 GND.n1550 585
R2139 GND.n2112 GND.n2111 585
R2140 GND.n2111 GND.n2110 585
R2141 GND.n2113 GND.n1546 585
R2142 GND.n1571 GND.n1546 585
R2143 GND.n2116 GND.n2115 585
R2144 GND.n2117 GND.n2116 585
R2145 GND.n1548 GND.n1545 585
R2146 GND.n1545 GND.n1536 585
R2147 GND.n1527 GND.n1526 585
R2148 GND.n2124 GND.n1527 585
R2149 GND.n2129 GND.n2128 585
R2150 GND.n2128 GND.n2127 585
R2151 GND.n2130 GND.n1524 585
R2152 GND.n1574 GND.n1524 585
R2153 GND.n2133 GND.n2132 585
R2154 GND.n2134 GND.n2133 585
R2155 GND.n1525 GND.n1523 585
R2156 GND.n1523 GND.n1518 585
R2157 GND.n2066 GND.n2065 585
R2158 GND.n2067 GND.n2066 585
R2159 GND.n1585 GND.n1584 585
R2160 GND.n2054 GND.n1584 585
R2161 GND.n2060 GND.n2059 585
R2162 GND.n2059 GND.n2058 585
R2163 GND.n1588 GND.n1587 585
R2164 GND.n2043 GND.n1588 585
R2165 GND.n2028 GND.n1610 585
R2166 GND.n1610 GND.n1599 585
R2167 GND.n2030 GND.n2029 585
R2168 GND.n2031 GND.n2030 585
R2169 GND.n1611 GND.n1609 585
R2170 GND.n2018 GND.n1609 585
R2171 GND.n2023 GND.n2022 585
R2172 GND.n2022 GND.n2021 585
R2173 GND.n1614 GND.n1613 585
R2174 GND.n2005 GND.n1614 585
R2175 GND.n1637 GND.n1636 585
R2176 GND.n1638 GND.n1637 585
R2177 GND.n1127 GND.n1126 585
R2178 GND.n1996 GND.n1127 585
R2179 GND.n4880 GND.n4879 585
R2180 GND.n4879 GND.n4878 585
R2181 GND.n4881 GND.n1121 585
R2182 GND.n1646 GND.n1121 585
R2183 GND.n4883 GND.n4882 585
R2184 GND.n4884 GND.n4883 585
R2185 GND.n1122 GND.n1120 585
R2186 GND.n1120 GND.n1115 585
R2187 GND.n1985 GND.n1984 585
R2188 GND.n1986 GND.n1985 585
R2189 GND.n1655 GND.n1654 585
R2190 GND.n1654 GND.n1651 585
R2191 GND.n1979 GND.n1978 585
R2192 GND.n1978 GND.n1977 585
R2193 GND.n1658 GND.n1657 585
R2194 GND.n1659 GND.n1658 585
R2195 GND.n1955 GND.n1954 585
R2196 GND.n1956 GND.n1955 585
R2197 GND.n1674 GND.n1673 585
R2198 GND.n1673 GND.n1670 585
R2199 GND.n1950 GND.n1949 585
R2200 GND.n1949 GND.n1948 585
R2201 GND.n1677 GND.n1676 585
R2202 GND.n1940 GND.n1677 585
R2203 GND.n1916 GND.n1700 585
R2204 GND.n1700 GND.n1690 585
R2205 GND.n1918 GND.n1917 585
R2206 GND.n1919 GND.n1918 585
R2207 GND.n1912 GND.n1699 585
R2208 GND.n1911 GND.n1910 585
R2209 GND.n1908 GND.n1702 585
R2210 GND.n1908 GND.n1696 585
R2211 GND.n1907 GND.n1906 585
R2212 GND.n1905 GND.n1904 585
R2213 GND.n1903 GND.n1707 585
R2214 GND.n1901 GND.n1900 585
R2215 GND.n1899 GND.n1708 585
R2216 GND.n1898 GND.n1897 585
R2217 GND.n1895 GND.n1713 585
R2218 GND.n1893 GND.n1892 585
R2219 GND.n1891 GND.n1714 585
R2220 GND.n1890 GND.n1889 585
R2221 GND.n1887 GND.n1719 585
R2222 GND.n1885 GND.n1884 585
R2223 GND.n1883 GND.n1720 585
R2224 GND.n1882 GND.n1881 585
R2225 GND.n1879 GND.n1725 585
R2226 GND.n1877 GND.n1876 585
R2227 GND.n1875 GND.n1726 585
R2228 GND.n1874 GND.n1873 585
R2229 GND.n1871 GND.n1734 585
R2230 GND.n1869 GND.n1868 585
R2231 GND.n1867 GND.n1735 585
R2232 GND.n1866 GND.n1865 585
R2233 GND.n1863 GND.n1740 585
R2234 GND.n1861 GND.n1860 585
R2235 GND.n1859 GND.n1741 585
R2236 GND.n1858 GND.n1857 585
R2237 GND.n1855 GND.n1746 585
R2238 GND.n1853 GND.n1852 585
R2239 GND.n1851 GND.n1747 585
R2240 GND.n1850 GND.n1849 585
R2241 GND.n1847 GND.n1752 585
R2242 GND.n1845 GND.n1844 585
R2243 GND.n1843 GND.n1753 585
R2244 GND.n1842 GND.n1758 585
R2245 GND.n1835 GND.n1761 585
R2246 GND.n1838 GND.n1837 585
R2247 GND.n4740 GND.n1235 585
R2248 GND.n4741 GND.n4739 585
R2249 GND.n1294 GND.n1290 585
R2250 GND.n4745 GND.n1289 585
R2251 GND.n4746 GND.n1288 585
R2252 GND.n4747 GND.n1287 585
R2253 GND.n4713 GND.n1285 585
R2254 GND.n4751 GND.n1284 585
R2255 GND.n4752 GND.n1283 585
R2256 GND.n4753 GND.n1282 585
R2257 GND.n4716 GND.n1280 585
R2258 GND.n4757 GND.n1279 585
R2259 GND.n4758 GND.n1278 585
R2260 GND.n4759 GND.n1277 585
R2261 GND.n4719 GND.n1275 585
R2262 GND.n4763 GND.n1274 585
R2263 GND.n4764 GND.n1273 585
R2264 GND.n4765 GND.n1272 585
R2265 GND.n4722 GND.n1270 585
R2266 GND.n4769 GND.n1269 585
R2267 GND.n4770 GND.n1268 585
R2268 GND.n4725 GND.n1262 585
R2269 GND.n4775 GND.n1261 585
R2270 GND.n4776 GND.n1260 585
R2271 GND.n4777 GND.n1259 585
R2272 GND.n4728 GND.n1257 585
R2273 GND.n4781 GND.n1256 585
R2274 GND.n4782 GND.n1255 585
R2275 GND.n4783 GND.n1254 585
R2276 GND.n4731 GND.n1252 585
R2277 GND.n4787 GND.n1251 585
R2278 GND.n4788 GND.n1250 585
R2279 GND.n4789 GND.n1249 585
R2280 GND.n4734 GND.n1247 585
R2281 GND.n4793 GND.n1246 585
R2282 GND.n4794 GND.n1245 585
R2283 GND.n4795 GND.n1241 585
R2284 GND.n4737 GND.n1241 585
R2285 GND.n4802 GND.n4801 585
R2286 GND.n4801 GND.n4800 585
R2287 GND.n1234 GND.n1229 585
R2288 GND.n2329 GND.n1234 585
R2289 GND.n4806 GND.n1228 585
R2290 GND.n2326 GND.n1228 585
R2291 GND.n4807 GND.n1227 585
R2292 GND.n2307 GND.n1227 585
R2293 GND.n4808 GND.n1226 585
R2294 GND.n2318 GND.n1226 585
R2295 GND.n1415 GND.n1221 585
R2296 GND.n2315 GND.n1415 585
R2297 GND.n4812 GND.n1220 585
R2298 GND.n2286 GND.n1220 585
R2299 GND.n4813 GND.n1219 585
R2300 GND.n1428 GND.n1219 585
R2301 GND.n4814 GND.n1218 585
R2302 GND.n2278 GND.n1218 585
R2303 GND.n1438 GND.n1213 585
R2304 GND.n2273 GND.n1438 585
R2305 GND.n4818 GND.n1212 585
R2306 GND.n2170 GND.n1212 585
R2307 GND.n4819 GND.n1211 585
R2308 GND.n2261 GND.n1211 585
R2309 GND.n4820 GND.n1210 585
R2310 GND.n2248 GND.n1210 585
R2311 GND.n1456 GND.n1205 585
R2312 GND.n2251 GND.n1456 585
R2313 GND.n4824 GND.n1204 585
R2314 GND.n2246 GND.n1204 585
R2315 GND.n4825 GND.n1203 585
R2316 GND.n2151 GND.n1203 585
R2317 GND.n4826 GND.n1202 585
R2318 GND.n2237 GND.n1202 585
R2319 GND.n2223 GND.n1197 585
R2320 GND.n2224 GND.n2223 585
R2321 GND.n4830 GND.n1196 585
R2322 GND.n2227 GND.n1196 585
R2323 GND.n4831 GND.n1195 585
R2324 GND.n2221 GND.n1195 585
R2325 GND.n4832 GND.n1194 585
R2326 GND.n1493 GND.n1194 585
R2327 GND.n1489 GND.n1189 585
R2328 GND.n2212 GND.n1489 585
R2329 GND.n4836 GND.n1188 585
R2330 GND.n2198 GND.n1188 585
R2331 GND.n4837 GND.n1187 585
R2332 GND.n2202 GND.n1187 585
R2333 GND.n4838 GND.n1186 585
R2334 GND.n2196 GND.n1186 585
R2335 GND.n1560 GND.n1181 585
R2336 GND.n2100 GND.n1560 585
R2337 GND.n4842 GND.n1180 585
R2338 GND.n1557 GND.n1180 585
R2339 GND.n4843 GND.n1179 585
R2340 GND.n2107 GND.n1179 585
R2341 GND.n4844 GND.n1178 585
R2342 GND.n2110 GND.n1178 585
R2343 GND.n1566 GND.n1173 585
R2344 GND.n1571 GND.n1566 585
R2345 GND.n4848 GND.n1172 585
R2346 GND.n2117 GND.n1172 585
R2347 GND.n4849 GND.n1171 585
R2348 GND.n1536 GND.n1171 585
R2349 GND.n4850 GND.n1170 585
R2350 GND.n2124 GND.n1170 585
R2351 GND.n1529 GND.n1165 585
R2352 GND.n2127 GND.n1529 585
R2353 GND.n4854 GND.n1164 585
R2354 GND.n1574 GND.n1164 585
R2355 GND.n4855 GND.n1163 585
R2356 GND.n2134 GND.n1163 585
R2357 GND.n4856 GND.n1162 585
R2358 GND.n1518 GND.n1162 585
R2359 GND.n1580 GND.n1157 585
R2360 GND.n2067 GND.n1580 585
R2361 GND.n4860 GND.n1156 585
R2362 GND.n2054 GND.n1156 585
R2363 GND.n4861 GND.n1155 585
R2364 GND.n2058 GND.n1155 585
R2365 GND.n4862 GND.n1154 585
R2366 GND.n2043 GND.n1154 585
R2367 GND.n1598 GND.n1149 585
R2368 GND.n1599 GND.n1598 585
R2369 GND.n4866 GND.n1148 585
R2370 GND.n2031 GND.n1148 585
R2371 GND.n4867 GND.n1147 585
R2372 GND.n2018 GND.n1147 585
R2373 GND.n4868 GND.n1146 585
R2374 GND.n2021 GND.n1146 585
R2375 GND.n1639 GND.n1141 585
R2376 GND.n2005 GND.n1639 585
R2377 GND.n4872 GND.n1140 585
R2378 GND.n1638 GND.n1140 585
R2379 GND.n4873 GND.n1139 585
R2380 GND.n1996 GND.n1139 585
R2381 GND.n4874 GND.n1129 585
R2382 GND.n4878 GND.n1129 585
R2383 GND.n1645 GND.n1138 585
R2384 GND.n1646 GND.n1645 585
R2385 GND.n1967 GND.n1116 585
R2386 GND.n4884 GND.n1116 585
R2387 GND.n1962 GND.n1961 585
R2388 GND.n1961 GND.n1115 585
R2389 GND.n1971 GND.n1652 585
R2390 GND.n1986 GND.n1652 585
R2391 GND.n1972 GND.n1960 585
R2392 GND.n1960 GND.n1651 585
R2393 GND.n1973 GND.n1660 585
R2394 GND.n1977 GND.n1660 585
R2395 GND.n1959 GND.n1958 585
R2396 GND.n1958 GND.n1659 585
R2397 GND.n1957 GND.n1668 585
R2398 GND.n1957 GND.n1956 585
R2399 GND.n1943 GND.n1669 585
R2400 GND.n1670 GND.n1669 585
R2401 GND.n1944 GND.n1678 585
R2402 GND.n1948 GND.n1678 585
R2403 GND.n1942 GND.n1941 585
R2404 GND.n1941 GND.n1940 585
R2405 GND.n1689 GND.n1688 585
R2406 GND.n1690 GND.n1689 585
R2407 GND.n1766 GND.n1697 585
R2408 GND.n1919 GND.n1697 585
R2409 GND.n5832 GND.n5831 585
R2410 GND.n5833 GND.n5832 585
R2411 GND.n460 GND.n459 585
R2412 GND.n463 GND.n460 585
R2413 GND.n5841 GND.n5840 585
R2414 GND.n5840 GND.n5839 585
R2415 GND.n5842 GND.n454 585
R2416 GND.n454 GND.n453 585
R2417 GND.n5844 GND.n5843 585
R2418 GND.n5845 GND.n5844 585
R2419 GND.n441 GND.n440 585
R2420 GND.n444 GND.n441 585
R2421 GND.n5853 GND.n5852 585
R2422 GND.n5852 GND.n5851 585
R2423 GND.n5854 GND.n435 585
R2424 GND.n435 GND.n434 585
R2425 GND.n5856 GND.n5855 585
R2426 GND.n5857 GND.n5856 585
R2427 GND.n421 GND.n420 585
R2428 GND.n431 GND.n421 585
R2429 GND.n5865 GND.n5864 585
R2430 GND.n5864 GND.n5863 585
R2431 GND.n5866 GND.n415 585
R2432 GND.n5693 GND.n415 585
R2433 GND.n5868 GND.n5867 585
R2434 GND.n5869 GND.n5868 585
R2435 GND.n401 GND.n400 585
R2436 GND.n5699 GND.n401 585
R2437 GND.n5877 GND.n5876 585
R2438 GND.n5876 GND.n5875 585
R2439 GND.n5878 GND.n395 585
R2440 GND.n5669 GND.n395 585
R2441 GND.n5880 GND.n5879 585
R2442 GND.n5881 GND.n5880 585
R2443 GND.n380 GND.n379 585
R2444 GND.n4251 GND.n380 585
R2445 GND.n5889 GND.n5888 585
R2446 GND.n5888 GND.n5887 585
R2447 GND.n5890 GND.n374 585
R2448 GND.n4257 GND.n374 585
R2449 GND.n5892 GND.n5891 585
R2450 GND.n5893 GND.n5892 585
R2451 GND.n359 GND.n358 585
R2452 GND.n4263 GND.n359 585
R2453 GND.n5901 GND.n5900 585
R2454 GND.n5900 GND.n5899 585
R2455 GND.n5902 GND.n354 585
R2456 GND.n4269 GND.n354 585
R2457 GND.n5904 GND.n5903 585
R2458 GND.n5905 GND.n5904 585
R2459 GND.n338 GND.n336 585
R2460 GND.n4231 GND.n338 585
R2461 GND.n5913 GND.n5912 585
R2462 GND.n5912 GND.n5911 585
R2463 GND.n337 GND.n335 585
R2464 GND.n4222 GND.n337 585
R2465 GND.n2753 GND.n2752 585
R2466 GND.n2754 GND.n2753 585
R2467 GND.n327 GND.n325 585
R2468 GND.n4308 GND.n325 585
R2469 GND.n5917 GND.n5916 585
R2470 GND.n5918 GND.n5917 585
R2471 GND.n326 GND.n324 585
R2472 GND.n4314 GND.n324 585
R2473 GND.n2723 GND.n2722 585
R2474 GND.n2724 GND.n2723 585
R2475 GND.n2711 GND.n333 585
R2476 GND.n2715 GND.n2711 585
R2477 GND.n4324 GND.n2712 585
R2478 GND.n4324 GND.n4323 585
R2479 GND.n4326 GND.n4325 585
R2480 GND.n4327 GND.n4326 585
R2481 GND.n2696 GND.n2695 585
R2482 GND.n4201 GND.n2696 585
R2483 GND.n4335 GND.n4334 585
R2484 GND.n4334 GND.n4333 585
R2485 GND.n4336 GND.n2690 585
R2486 GND.n4183 GND.n2690 585
R2487 GND.n4338 GND.n4337 585
R2488 GND.n4339 GND.n4338 585
R2489 GND.n2675 GND.n2674 585
R2490 GND.n4176 GND.n2675 585
R2491 GND.n4347 GND.n4346 585
R2492 GND.n4346 GND.n4345 585
R2493 GND.n4348 GND.n2669 585
R2494 GND.n4168 GND.n2669 585
R2495 GND.n4350 GND.n4349 585
R2496 GND.n4351 GND.n4350 585
R2497 GND.n2654 GND.n2653 585
R2498 GND.n4161 GND.n2654 585
R2499 GND.n4359 GND.n4358 585
R2500 GND.n4358 GND.n4357 585
R2501 GND.n4360 GND.n2648 585
R2502 GND.n4153 GND.n2648 585
R2503 GND.n4362 GND.n4361 585
R2504 GND.n4363 GND.n4362 585
R2505 GND.n2634 GND.n2633 585
R2506 GND.n4146 GND.n2634 585
R2507 GND.n4371 GND.n4370 585
R2508 GND.n4370 GND.n4369 585
R2509 GND.n4372 GND.n2628 585
R2510 GND.n4138 GND.n2628 585
R2511 GND.n4374 GND.n4373 585
R2512 GND.n4375 GND.n4374 585
R2513 GND.n2613 GND.n2612 585
R2514 GND.n4131 GND.n2613 585
R2515 GND.n4383 GND.n4382 585
R2516 GND.n4382 GND.n4381 585
R2517 GND.n4384 GND.n2607 585
R2518 GND.n4123 GND.n2607 585
R2519 GND.n4386 GND.n4385 585
R2520 GND.n4387 GND.n4386 585
R2521 GND.n2589 GND.n2588 585
R2522 GND.n4116 GND.n2589 585
R2523 GND.n4395 GND.n4394 585
R2524 GND.n4394 GND.n4393 585
R2525 GND.n4396 GND.n2580 585
R2526 GND.n4108 GND.n2580 585
R2527 GND.n4398 GND.n4397 585
R2528 GND.n4399 GND.n4398 585
R2529 GND.n2581 GND.n2579 585
R2530 GND.n3988 GND.n2579 585
R2531 GND.n2582 GND.n2519 585
R2532 GND.n4407 GND.n2519 585
R2533 GND.n4481 GND.n4480 585
R2534 GND.n4479 GND.n2518 585
R2535 GND.n4478 GND.n2517 585
R2536 GND.n4483 GND.n2517 585
R2537 GND.n4477 GND.n4476 585
R2538 GND.n4475 GND.n4474 585
R2539 GND.n4473 GND.n4472 585
R2540 GND.n4471 GND.n4470 585
R2541 GND.n4469 GND.n4468 585
R2542 GND.n4467 GND.n4466 585
R2543 GND.n4465 GND.n4464 585
R2544 GND.n4463 GND.n4462 585
R2545 GND.n4461 GND.n4460 585
R2546 GND.n4459 GND.n4458 585
R2547 GND.n4457 GND.n4456 585
R2548 GND.n4455 GND.n4454 585
R2549 GND.n4453 GND.n4452 585
R2550 GND.n4450 GND.n4449 585
R2551 GND.n4448 GND.n4447 585
R2552 GND.n4446 GND.n4445 585
R2553 GND.n4444 GND.n4443 585
R2554 GND.n4442 GND.n4441 585
R2555 GND.n4440 GND.n4439 585
R2556 GND.n4438 GND.n4437 585
R2557 GND.n4436 GND.n4435 585
R2558 GND.n4434 GND.n4433 585
R2559 GND.n4432 GND.n4431 585
R2560 GND.n4430 GND.n4429 585
R2561 GND.n4428 GND.n4427 585
R2562 GND.n4426 GND.n4425 585
R2563 GND.n4424 GND.n4423 585
R2564 GND.n4422 GND.n4421 585
R2565 GND.n4420 GND.n4419 585
R2566 GND.n4418 GND.n4417 585
R2567 GND.n4416 GND.n4415 585
R2568 GND.n4414 GND.n2559 585
R2569 GND.n2563 GND.n2560 585
R2570 GND.n4410 GND.n4409 585
R2571 GND.n540 GND.n539 585
R2572 GND.n5761 GND.n535 585
R2573 GND.n5763 GND.n5762 585
R2574 GND.n5765 GND.n533 585
R2575 GND.n5767 GND.n5766 585
R2576 GND.n5768 GND.n528 585
R2577 GND.n5770 GND.n5769 585
R2578 GND.n5772 GND.n526 585
R2579 GND.n5774 GND.n5773 585
R2580 GND.n5775 GND.n521 585
R2581 GND.n5777 GND.n5776 585
R2582 GND.n5779 GND.n519 585
R2583 GND.n5781 GND.n5780 585
R2584 GND.n5782 GND.n514 585
R2585 GND.n5784 GND.n5783 585
R2586 GND.n5786 GND.n512 585
R2587 GND.n5788 GND.n5787 585
R2588 GND.n5789 GND.n507 585
R2589 GND.n5791 GND.n5790 585
R2590 GND.n5793 GND.n505 585
R2591 GND.n5795 GND.n5794 585
R2592 GND.n5799 GND.n500 585
R2593 GND.n5801 GND.n5800 585
R2594 GND.n5803 GND.n498 585
R2595 GND.n5805 GND.n5804 585
R2596 GND.n5806 GND.n493 585
R2597 GND.n5808 GND.n5807 585
R2598 GND.n5810 GND.n491 585
R2599 GND.n5812 GND.n5811 585
R2600 GND.n5813 GND.n486 585
R2601 GND.n5815 GND.n5814 585
R2602 GND.n5817 GND.n484 585
R2603 GND.n5819 GND.n5818 585
R2604 GND.n5820 GND.n479 585
R2605 GND.n5822 GND.n5821 585
R2606 GND.n5824 GND.n477 585
R2607 GND.n5826 GND.n5825 585
R2608 GND.n5827 GND.n475 585
R2609 GND.n5828 GND.n472 585
R2610 GND.n472 GND.n471 585
R2611 GND.n5676 GND.n469 585
R2612 GND.n5833 GND.n469 585
R2613 GND.n5678 GND.n5677 585
R2614 GND.n5677 GND.n463 585
R2615 GND.n5679 GND.n461 585
R2616 GND.n5839 GND.n461 585
R2617 GND.n5681 GND.n5680 585
R2618 GND.n5680 GND.n453 585
R2619 GND.n5682 GND.n451 585
R2620 GND.n5845 GND.n451 585
R2621 GND.n5684 GND.n5683 585
R2622 GND.n5683 GND.n444 585
R2623 GND.n5685 GND.n442 585
R2624 GND.n5851 GND.n442 585
R2625 GND.n5687 GND.n5686 585
R2626 GND.n5686 GND.n434 585
R2627 GND.n5688 GND.n432 585
R2628 GND.n5857 GND.n432 585
R2629 GND.n5690 GND.n5689 585
R2630 GND.n5689 GND.n431 585
R2631 GND.n5691 GND.n423 585
R2632 GND.n5863 GND.n423 585
R2633 GND.n5695 GND.n5694 585
R2634 GND.n5694 GND.n5693 585
R2635 GND.n5696 GND.n412 585
R2636 GND.n5869 GND.n412 585
R2637 GND.n5698 GND.n5697 585
R2638 GND.n5699 GND.n5698 585
R2639 GND.n5672 GND.n402 585
R2640 GND.n5875 GND.n402 585
R2641 GND.n5671 GND.n5670 585
R2642 GND.n5670 GND.n5669 585
R2643 GND.n587 GND.n392 585
R2644 GND.n5881 GND.n392 585
R2645 GND.n4250 GND.n4249 585
R2646 GND.n4251 GND.n4250 585
R2647 GND.n4239 GND.n382 585
R2648 GND.n5887 GND.n382 585
R2649 GND.n4259 GND.n4258 585
R2650 GND.n4258 GND.n4257 585
R2651 GND.n4260 GND.n371 585
R2652 GND.n5893 GND.n371 585
R2653 GND.n4262 GND.n4261 585
R2654 GND.n4263 GND.n4262 585
R2655 GND.n4237 GND.n361 585
R2656 GND.n5899 GND.n361 585
R2657 GND.n4236 GND.n2740 585
R2658 GND.n4269 GND.n2740 585
R2659 GND.n4234 GND.n352 585
R2660 GND.n5905 GND.n352 585
R2661 GND.n4233 GND.n4232 585
R2662 GND.n4232 GND.n4231 585
R2663 GND.n2746 GND.n340 585
R2664 GND.n5911 GND.n340 585
R2665 GND.n4221 GND.n4220 585
R2666 GND.n4222 GND.n4221 585
R2667 GND.n4217 GND.n2755 585
R2668 GND.n2755 GND.n2754 585
R2669 GND.n4216 GND.n2733 585
R2670 GND.n4308 GND.n2733 585
R2671 GND.n4215 GND.n321 585
R2672 GND.n5918 GND.n321 585
R2673 GND.n4214 GND.n2725 585
R2674 GND.n4314 GND.n2725 585
R2675 GND.n4213 GND.n4212 585
R2676 GND.n4212 GND.n2724 585
R2677 GND.n4211 GND.n2756 585
R2678 GND.n4211 GND.n2715 585
R2679 GND.n4205 GND.n2713 585
R2680 GND.n4323 GND.n2713 585
R2681 GND.n4204 GND.n2708 585
R2682 GND.n4327 GND.n2708 585
R2683 GND.n4203 GND.n4202 585
R2684 GND.n4202 GND.n4201 585
R2685 GND.n2757 GND.n2698 585
R2686 GND.n4333 GND.n2698 585
R2687 GND.n4182 GND.n4181 585
R2688 GND.n4183 GND.n4182 585
R2689 GND.n4179 GND.n2687 585
R2690 GND.n4339 GND.n2687 585
R2691 GND.n4178 GND.n4177 585
R2692 GND.n4177 GND.n4176 585
R2693 GND.n2761 GND.n2677 585
R2694 GND.n4345 GND.n2677 585
R2695 GND.n4167 GND.n4166 585
R2696 GND.n4168 GND.n4167 585
R2697 GND.n4164 GND.n2666 585
R2698 GND.n4351 GND.n2666 585
R2699 GND.n4163 GND.n4162 585
R2700 GND.n4162 GND.n4161 585
R2701 GND.n2765 GND.n2656 585
R2702 GND.n4357 GND.n2656 585
R2703 GND.n4152 GND.n4151 585
R2704 GND.n4153 GND.n4152 585
R2705 GND.n4149 GND.n2646 585
R2706 GND.n4363 GND.n2646 585
R2707 GND.n4148 GND.n4147 585
R2708 GND.n4147 GND.n4146 585
R2709 GND.n2770 GND.n2636 585
R2710 GND.n4369 GND.n2636 585
R2711 GND.n4137 GND.n4136 585
R2712 GND.n4138 GND.n4137 585
R2713 GND.n4134 GND.n2625 585
R2714 GND.n4375 GND.n2625 585
R2715 GND.n4133 GND.n4132 585
R2716 GND.n4132 GND.n4131 585
R2717 GND.n2774 GND.n2615 585
R2718 GND.n4381 GND.n2615 585
R2719 GND.n4122 GND.n4121 585
R2720 GND.n4123 GND.n4122 585
R2721 GND.n4119 GND.n2604 585
R2722 GND.n4387 GND.n2604 585
R2723 GND.n4118 GND.n4117 585
R2724 GND.n4117 GND.n4116 585
R2725 GND.n2778 GND.n2591 585
R2726 GND.n4393 GND.n2591 585
R2727 GND.n2575 GND.n2574 585
R2728 GND.n4108 GND.n2575 585
R2729 GND.n4401 GND.n4400 585
R2730 GND.n4400 GND.n4399 585
R2731 GND.n4402 GND.n2564 585
R2732 GND.n3988 GND.n2564 585
R2733 GND.n4408 GND.n2565 585
R2734 GND.n4408 GND.n4407 585
R2735 GND.n3830 GND.n2870 585
R2736 GND.n2870 GND.n2838 585
R2737 GND.n3829 GND.n3828 585
R2738 GND.n3828 GND.n3827 585
R2739 GND.n2892 GND.n2891 585
R2740 GND.n3803 GND.n2892 585
R2741 GND.n3816 GND.n3815 585
R2742 GND.n3817 GND.n3816 585
R2743 GND.n3814 GND.n2903 585
R2744 GND.n3809 GND.n2903 585
R2745 GND.n3813 GND.n3812 585
R2746 GND.n3812 GND.n3811 585
R2747 GND.n2905 GND.n2904 585
R2748 GND.n3792 GND.n2905 585
R2749 GND.n3783 GND.n2987 585
R2750 GND.n2987 GND.n2986 585
R2751 GND.n3785 GND.n3784 585
R2752 GND.n3786 GND.n3785 585
R2753 GND.n3782 GND.n2984 585
R2754 GND.n2992 GND.n2984 585
R2755 GND.n3781 GND.n3780 585
R2756 GND.n3780 GND.n3779 585
R2757 GND.n2989 GND.n2988 585
R2758 GND.n3737 GND.n2989 585
R2759 GND.n3016 GND.n3015 585
R2760 GND.n3016 GND.n3001 585
R2761 GND.n3745 GND.n3744 585
R2762 GND.n3744 GND.n3743 585
R2763 GND.n3746 GND.n3013 585
R2764 GND.n3018 GND.n3013 585
R2765 GND.n3748 GND.n3747 585
R2766 GND.n3749 GND.n3748 585
R2767 GND.n3014 GND.n3012 585
R2768 GND.n3730 GND.n3012 585
R2769 GND.n3727 GND.n3726 585
R2770 GND.n3728 GND.n3727 585
R2771 GND.n3725 GND.n3024 585
R2772 GND.n3029 GND.n3024 585
R2773 GND.n3724 GND.n3723 585
R2774 GND.n3723 GND.n3722 585
R2775 GND.n3026 GND.n3025 585
R2776 GND.n3616 GND.n3026 585
R2777 GND.n3706 GND.n3705 585
R2778 GND.n3707 GND.n3706 585
R2779 GND.n3704 GND.n3039 585
R2780 GND.n3039 GND.n3036 585
R2781 GND.n3703 GND.n3702 585
R2782 GND.n3702 GND.n3701 585
R2783 GND.n3041 GND.n3040 585
R2784 GND.n3625 GND.n3041 585
R2785 GND.n3681 GND.n3680 585
R2786 GND.n3682 GND.n3681 585
R2787 GND.n3679 GND.n3054 585
R2788 GND.n3054 GND.n3051 585
R2789 GND.n3678 GND.n3677 585
R2790 GND.n3677 GND.n3676 585
R2791 GND.n3056 GND.n3055 585
R2792 GND.n3066 GND.n3056 585
R2793 GND.n3650 GND.n3649 585
R2794 GND.n3649 GND.n3065 585
R2795 GND.n3651 GND.n3076 585
R2796 GND.n3637 GND.n3076 585
R2797 GND.n3653 GND.n3652 585
R2798 GND.n3654 GND.n3653 585
R2799 GND.n3648 GND.n3075 585
R2800 GND.n3643 GND.n3075 585
R2801 GND.n3647 GND.n3646 585
R2802 GND.n3646 GND.n3645 585
R2803 GND.n3078 GND.n3077 585
R2804 GND.n3607 GND.n3078 585
R2805 GND.n3593 GND.n3592 585
R2806 GND.n3592 GND.n3591 585
R2807 GND.n3594 GND.n3093 585
R2808 GND.n3588 GND.n3093 585
R2809 GND.n3596 GND.n3595 585
R2810 GND.n3597 GND.n3596 585
R2811 GND.n3094 GND.n3092 585
R2812 GND.n3582 GND.n3092 585
R2813 GND.n3579 GND.n3578 585
R2814 GND.n3580 GND.n3579 585
R2815 GND.n3577 GND.n3098 585
R2816 GND.n3104 GND.n3098 585
R2817 GND.n3576 GND.n3575 585
R2818 GND.n3575 GND.n3574 585
R2819 GND.n3100 GND.n3099 585
R2820 GND.n3152 GND.n3100 585
R2821 GND.n3546 GND.n3545 585
R2822 GND.n3547 GND.n3546 585
R2823 GND.n3544 GND.n3114 585
R2824 GND.n3114 GND.n3111 585
R2825 GND.n3543 GND.n3542 585
R2826 GND.n3542 GND.n3541 585
R2827 GND.n3116 GND.n3115 585
R2828 GND.n3160 GND.n3116 585
R2829 GND.n3523 GND.n3522 585
R2830 GND.n3524 GND.n3523 585
R2831 GND.n3521 GND.n3130 585
R2832 GND.n3130 GND.n3126 585
R2833 GND.n3520 GND.n3519 585
R2834 GND.n3519 GND.n3518 585
R2835 GND.n3132 GND.n3131 585
R2836 GND.n3491 GND.n3132 585
R2837 GND.n3504 GND.n3503 585
R2838 GND.n3505 GND.n3504 585
R2839 GND.n3502 GND.n3143 585
R2840 GND.n3497 GND.n3143 585
R2841 GND.n3501 GND.n3500 585
R2842 GND.n3500 GND.n3499 585
R2843 GND.n3145 GND.n3144 585
R2844 GND.n3172 GND.n3145 585
R2845 GND.n3360 GND.n3359 585
R2846 GND.n3361 GND.n3360 585
R2847 GND.n3357 GND.n3181 585
R2848 GND.n3356 GND.n3355 585
R2849 GND.n3353 GND.n3202 585
R2850 GND.n3353 GND.n3178 585
R2851 GND.n3352 GND.n3351 585
R2852 GND.n3350 GND.n3349 585
R2853 GND.n3348 GND.n3204 585
R2854 GND.n3346 GND.n3345 585
R2855 GND.n3344 GND.n3205 585
R2856 GND.n3343 GND.n3342 585
R2857 GND.n3340 GND.n3206 585
R2858 GND.n3338 GND.n3337 585
R2859 GND.n3336 GND.n3207 585
R2860 GND.n3335 GND.n3334 585
R2861 GND.n3332 GND.n3208 585
R2862 GND.n3330 GND.n3329 585
R2863 GND.n3328 GND.n3209 585
R2864 GND.n3327 GND.n3326 585
R2865 GND.n3324 GND.n3210 585
R2866 GND.n3322 GND.n3321 585
R2867 GND.n3320 GND.n3211 585
R2868 GND.n3319 GND.n3318 585
R2869 GND.n3316 GND.n3212 585
R2870 GND.n3314 GND.n3313 585
R2871 GND.n3312 GND.n3213 585
R2872 GND.n3311 GND.n3310 585
R2873 GND.n3308 GND.n3214 585
R2874 GND.n3306 GND.n3305 585
R2875 GND.n3304 GND.n3215 585
R2876 GND.n3303 GND.n3302 585
R2877 GND.n3300 GND.n1267 585
R2878 GND.n3296 GND.n3295 585
R2879 GND.n3294 GND.n3219 585
R2880 GND.n3293 GND.n3292 585
R2881 GND.n3290 GND.n3289 585
R2882 GND.n3288 GND.n3287 585
R2883 GND.n3286 GND.n3224 585
R2884 GND.n3284 GND.n3283 585
R2885 GND.n3282 GND.n3225 585
R2886 GND.n3281 GND.n3280 585
R2887 GND.n3278 GND.n3226 585
R2888 GND.n3276 GND.n3275 585
R2889 GND.n3274 GND.n3227 585
R2890 GND.n3273 GND.n3272 585
R2891 GND.n3270 GND.n3228 585
R2892 GND.n3268 GND.n3267 585
R2893 GND.n3266 GND.n3229 585
R2894 GND.n3265 GND.n3264 585
R2895 GND.n3262 GND.n3230 585
R2896 GND.n3260 GND.n3259 585
R2897 GND.n3258 GND.n3231 585
R2898 GND.n3257 GND.n3256 585
R2899 GND.n3254 GND.n3232 585
R2900 GND.n3252 GND.n3251 585
R2901 GND.n3250 GND.n3233 585
R2902 GND.n3249 GND.n3248 585
R2903 GND.n3246 GND.n3234 585
R2904 GND.n3244 GND.n3243 585
R2905 GND.n3242 GND.n3235 585
R2906 GND.n3241 GND.n3240 585
R2907 GND.n2968 GND.n2967 585
R2908 GND.n2966 GND.n2965 585
R2909 GND.n2964 GND.n2963 585
R2910 GND.n2962 GND.n2961 585
R2911 GND.n2960 GND.n2959 585
R2912 GND.n2958 GND.n2957 585
R2913 GND.n2956 GND.n2955 585
R2914 GND.n2954 GND.n2953 585
R2915 GND.n2952 GND.n2951 585
R2916 GND.n2950 GND.n2949 585
R2917 GND.n2948 GND.n2947 585
R2918 GND.n2946 GND.n2945 585
R2919 GND.n2944 GND.n2943 585
R2920 GND.n2942 GND.n2941 585
R2921 GND.n2940 GND.n2939 585
R2922 GND.n2938 GND.n2937 585
R2923 GND.n2936 GND.n2935 585
R2924 GND.n2934 GND.n2933 585
R2925 GND.n2932 GND.n2931 585
R2926 GND.n2930 GND.n2929 585
R2927 GND.n2928 GND.n2927 585
R2928 GND.n2926 GND.n2925 585
R2929 GND.n2924 GND.n2923 585
R2930 GND.n2922 GND.n2921 585
R2931 GND.n2920 GND.n2919 585
R2932 GND.n2918 GND.n2917 585
R2933 GND.n2916 GND.n2915 585
R2934 GND.n2914 GND.n2913 585
R2935 GND.n2912 GND.n2911 585
R2936 GND.n3834 GND.n2536 585
R2937 GND.n3836 GND.n3835 585
R2938 GND.n3838 GND.n3837 585
R2939 GND.n3840 GND.n3839 585
R2940 GND.n3843 GND.n3842 585
R2941 GND.n3845 GND.n3844 585
R2942 GND.n3847 GND.n3846 585
R2943 GND.n3849 GND.n3848 585
R2944 GND.n3851 GND.n3850 585
R2945 GND.n3853 GND.n3852 585
R2946 GND.n3855 GND.n3854 585
R2947 GND.n3857 GND.n3856 585
R2948 GND.n3859 GND.n3858 585
R2949 GND.n3861 GND.n3860 585
R2950 GND.n3863 GND.n3862 585
R2951 GND.n3865 GND.n3864 585
R2952 GND.n3867 GND.n3866 585
R2953 GND.n3869 GND.n3868 585
R2954 GND.n3871 GND.n3870 585
R2955 GND.n3873 GND.n3872 585
R2956 GND.n3875 GND.n3874 585
R2957 GND.n3877 GND.n3876 585
R2958 GND.n3879 GND.n3878 585
R2959 GND.n3881 GND.n3880 585
R2960 GND.n3883 GND.n3882 585
R2961 GND.n3885 GND.n3884 585
R2962 GND.n3887 GND.n3886 585
R2963 GND.n3889 GND.n3888 585
R2964 GND.n3890 GND.n2871 585
R2965 GND.n3892 GND.n3891 585
R2966 GND.n3893 GND.n3892 585
R2967 GND.n2970 GND.n2969 585
R2968 GND.n2969 GND.n2838 585
R2969 GND.n2971 GND.n2894 585
R2970 GND.n3827 GND.n2894 585
R2971 GND.n3805 GND.n3804 585
R2972 GND.n3804 GND.n3803 585
R2973 GND.n3806 GND.n2902 585
R2974 GND.n3817 GND.n2902 585
R2975 GND.n3808 GND.n3807 585
R2976 GND.n3809 GND.n3808 585
R2977 GND.n2907 GND.n2906 585
R2978 GND.n3811 GND.n2906 585
R2979 GND.n3791 GND.n3790 585
R2980 GND.n3792 GND.n3791 585
R2981 GND.n3789 GND.n2979 585
R2982 GND.n2986 GND.n2979 585
R2983 GND.n3788 GND.n3787 585
R2984 GND.n3787 GND.n3786 585
R2985 GND.n2981 GND.n2980 585
R2986 GND.n2992 GND.n2981 585
R2987 GND.n3735 GND.n2991 585
R2988 GND.n3779 GND.n2991 585
R2989 GND.n3739 GND.n3738 585
R2990 GND.n3738 GND.n3737 585
R2991 GND.n3740 GND.n3020 585
R2992 GND.n3020 GND.n3001 585
R2993 GND.n3742 GND.n3741 585
R2994 GND.n3743 GND.n3742 585
R2995 GND.n3734 GND.n3019 585
R2996 GND.n3019 GND.n3018 585
R2997 GND.n3733 GND.n3010 585
R2998 GND.n3749 GND.n3010 585
R2999 GND.n3732 GND.n3731 585
R3000 GND.n3731 GND.n3730 585
R3001 GND.n3022 GND.n3021 585
R3002 GND.n3728 GND.n3022 585
R3003 GND.n3613 GND.n3612 585
R3004 GND.n3612 GND.n3029 585
R3005 GND.n3614 GND.n3028 585
R3006 GND.n3722 GND.n3028 585
R3007 GND.n3618 GND.n3617 585
R3008 GND.n3617 GND.n3616 585
R3009 GND.n3619 GND.n3037 585
R3010 GND.n3707 GND.n3037 585
R3011 GND.n3621 GND.n3620 585
R3012 GND.n3620 GND.n3036 585
R3013 GND.n3622 GND.n3043 585
R3014 GND.n3701 GND.n3043 585
R3015 GND.n3627 GND.n3626 585
R3016 GND.n3626 GND.n3625 585
R3017 GND.n3628 GND.n3052 585
R3018 GND.n3682 GND.n3052 585
R3019 GND.n3630 GND.n3629 585
R3020 GND.n3629 GND.n3051 585
R3021 GND.n3631 GND.n3058 585
R3022 GND.n3676 GND.n3058 585
R3023 GND.n3633 GND.n3632 585
R3024 GND.n3633 GND.n3066 585
R3025 GND.n3634 GND.n3611 585
R3026 GND.n3634 GND.n3065 585
R3027 GND.n3639 GND.n3638 585
R3028 GND.n3638 GND.n3637 585
R3029 GND.n3640 GND.n3073 585
R3030 GND.n3654 GND.n3073 585
R3031 GND.n3642 GND.n3641 585
R3032 GND.n3643 GND.n3642 585
R3033 GND.n3610 GND.n3080 585
R3034 GND.n3645 GND.n3080 585
R3035 GND.n3609 GND.n3608 585
R3036 GND.n3608 GND.n3607 585
R3037 GND.n3082 GND.n3081 585
R3038 GND.n3591 GND.n3082 585
R3039 GND.n3587 GND.n3586 585
R3040 GND.n3588 GND.n3587 585
R3041 GND.n3585 GND.n3090 585
R3042 GND.n3597 GND.n3090 585
R3043 GND.n3584 GND.n3583 585
R3044 GND.n3583 GND.n3582 585
R3045 GND.n3096 GND.n3095 585
R3046 GND.n3580 GND.n3096 585
R3047 GND.n3149 GND.n3148 585
R3048 GND.n3148 GND.n3104 585
R3049 GND.n3150 GND.n3103 585
R3050 GND.n3574 GND.n3103 585
R3051 GND.n3154 GND.n3153 585
R3052 GND.n3153 GND.n3152 585
R3053 GND.n3155 GND.n3112 585
R3054 GND.n3547 GND.n3112 585
R3055 GND.n3157 GND.n3156 585
R3056 GND.n3156 GND.n3111 585
R3057 GND.n3158 GND.n3118 585
R3058 GND.n3541 GND.n3118 585
R3059 GND.n3162 GND.n3161 585
R3060 GND.n3161 GND.n3160 585
R3061 GND.n3163 GND.n3128 585
R3062 GND.n3524 GND.n3128 585
R3063 GND.n3165 GND.n3164 585
R3064 GND.n3164 GND.n3126 585
R3065 GND.n3166 GND.n3134 585
R3066 GND.n3518 GND.n3134 585
R3067 GND.n3493 GND.n3492 585
R3068 GND.n3492 GND.n3491 585
R3069 GND.n3494 GND.n3142 585
R3070 GND.n3505 GND.n3142 585
R3071 GND.n3496 GND.n3495 585
R3072 GND.n3497 GND.n3496 585
R3073 GND.n3147 GND.n3146 585
R3074 GND.n3499 GND.n3146 585
R3075 GND.n3237 GND.n3236 585
R3076 GND.n3236 GND.n3172 585
R3077 GND.n3238 GND.n3179 585
R3078 GND.n3361 GND.n3179 585
R3079 GND.n5661 GND.n5660 585
R3080 GND.n5661 GND.n422 585
R3081 GND.n5662 GND.n596 585
R3082 GND.n5662 GND.n414 585
R3083 GND.n5664 GND.n5663 585
R3084 GND.n5663 GND.n411 585
R3085 GND.n5665 GND.n591 585
R3086 GND.n591 GND.n404 585
R3087 GND.n5667 GND.n5666 585
R3088 GND.n5668 GND.n5667 585
R3089 GND.n592 GND.n590 585
R3090 GND.n590 GND.n394 585
R3091 GND.n4287 GND.n4286 585
R3092 GND.n4287 GND.n391 585
R3093 GND.n4288 GND.n4282 585
R3094 GND.n4288 GND.n384 585
R3095 GND.n4290 GND.n4289 585
R3096 GND.n4289 GND.n381 585
R3097 GND.n4291 GND.n4277 585
R3098 GND.n4277 GND.n373 585
R3099 GND.n4293 GND.n4292 585
R3100 GND.n4293 GND.n370 585
R3101 GND.n4294 GND.n4276 585
R3102 GND.n4294 GND.n363 585
R3103 GND.n4296 GND.n4295 585
R3104 GND.n4295 GND.n360 585
R3105 GND.n4297 GND.n4271 585
R3106 GND.n4271 GND.n4270 585
R3107 GND.n4299 GND.n4298 585
R3108 GND.n4299 GND.n351 585
R3109 GND.n4300 GND.n2739 585
R3110 GND.n4300 GND.n342 585
R3111 GND.n4302 GND.n4301 585
R3112 GND.n4301 GND.n339 585
R3113 GND.n4304 GND.n2735 585
R3114 GND.n2751 GND.n2735 585
R3115 GND.n4306 GND.n4305 585
R3116 GND.n4307 GND.n4306 585
R3117 GND.n2737 GND.n2734 585
R3118 GND.n2734 GND.n322 585
R3119 GND.n2736 GND.n2720 585
R3120 GND.n2720 GND.n320 585
R3121 GND.n4317 GND.n4316 585
R3122 GND.n4316 GND.n4315 585
R3123 GND.n4318 GND.n2717 585
R3124 GND.n2721 GND.n2717 585
R3125 GND.n4321 GND.n4320 585
R3126 GND.n4322 GND.n4321 585
R3127 GND.n2718 GND.n2716 585
R3128 GND.n2716 GND.n2710 585
R3129 GND.n4071 GND.n4070 585
R3130 GND.n4071 GND.n2707 585
R3131 GND.n4073 GND.n4072 585
R3132 GND.n4072 GND.n2700 585
R3133 GND.n4074 GND.n4064 585
R3134 GND.n4064 GND.n2697 585
R3135 GND.n4076 GND.n4075 585
R3136 GND.n4076 GND.n2689 585
R3137 GND.n4077 GND.n4063 585
R3138 GND.n4077 GND.n2686 585
R3139 GND.n4079 GND.n4078 585
R3140 GND.n4078 GND.n2679 585
R3141 GND.n4080 GND.n4058 585
R3142 GND.n4058 GND.n2676 585
R3143 GND.n4082 GND.n4081 585
R3144 GND.n4082 GND.n2668 585
R3145 GND.n4083 GND.n4057 585
R3146 GND.n4083 GND.n2665 585
R3147 GND.n4085 GND.n4084 585
R3148 GND.n4084 GND.n2658 585
R3149 GND.n4086 GND.n4052 585
R3150 GND.n4052 GND.n2655 585
R3151 GND.n4088 GND.n4087 585
R3152 GND.n4088 GND.n2769 585
R3153 GND.n4089 GND.n4051 585
R3154 GND.n4089 GND.n2645 585
R3155 GND.n4091 GND.n4090 585
R3156 GND.n4090 GND.n2638 585
R3157 GND.n4092 GND.n4046 585
R3158 GND.n4046 GND.n2635 585
R3159 GND.n4094 GND.n4093 585
R3160 GND.n4094 GND.n2627 585
R3161 GND.n4095 GND.n4045 585
R3162 GND.n4095 GND.n2624 585
R3163 GND.n4097 GND.n4096 585
R3164 GND.n4096 GND.n2617 585
R3165 GND.n4098 GND.n4040 585
R3166 GND.n4040 GND.n2614 585
R3167 GND.n4100 GND.n4099 585
R3168 GND.n4100 GND.n2606 585
R3169 GND.n4101 GND.n4039 585
R3170 GND.n4101 GND.n2603 585
R3171 GND.n4103 GND.n4102 585
R3172 GND.n4102 GND.n2593 585
R3173 GND.n4104 GND.n2783 585
R3174 GND.n2783 GND.n2590 585
R3175 GND.n4106 GND.n4105 585
R3176 GND.n4107 GND.n4106 585
R3177 GND.n2784 GND.n2782 585
R3178 GND.n2782 GND.n2576 585
R3179 GND.n4033 GND.n4032 585
R3180 GND.n4032 GND.n2568 585
R3181 GND.n4031 GND.n2786 585
R3182 GND.n4031 GND.n2566 585
R3183 GND.n4030 GND.n4029 585
R3184 GND.n4030 GND.n2516 585
R3185 GND.n2788 GND.n2787 585
R3186 GND.n2787 GND.n2484 585
R3187 GND.n4025 GND.n4024 585
R3188 GND.n4024 GND.n4023 585
R3189 GND.n2791 GND.n2790 585
R3190 GND.n4022 GND.n2791 585
R3191 GND.n3963 GND.n3962 585
R3192 GND.n3964 GND.n3963 585
R3193 GND.n2793 GND.n2792 585
R3194 GND.n2792 GND.n2429 585
R3195 GND.n3958 GND.n3957 585
R3196 GND.n3957 GND.n2428 585
R3197 GND.n3956 GND.n2795 585
R3198 GND.n3956 GND.n3955 585
R3199 GND.n3941 GND.n2796 585
R3200 GND.n2804 GND.n2796 585
R3201 GND.n3943 GND.n3942 585
R3202 GND.n3944 GND.n3943 585
R3203 GND.n2807 GND.n2806 585
R3204 GND.n2806 GND.n2803 585
R3205 GND.n3936 GND.n3935 585
R3206 GND.n3935 GND.n3934 585
R3207 GND.n2810 GND.n2809 585
R3208 GND.n2811 GND.n2810 585
R3209 GND.n3922 GND.n3921 585
R3210 GND.n3923 GND.n3922 585
R3211 GND.n2821 GND.n2820 585
R3212 GND.n2820 GND.n2818 585
R3213 GND.n3917 GND.n3916 585
R3214 GND.n3916 GND.n3915 585
R3215 GND.n2824 GND.n2823 585
R3216 GND.n2825 GND.n2824 585
R3217 GND.n3903 GND.n3902 585
R3218 GND.n3904 GND.n3903 585
R3219 GND.n2834 GND.n2833 585
R3220 GND.n3894 GND.n2833 585
R3221 GND.n3898 GND.n3897 585
R3222 GND.n3897 GND.n3896 585
R3223 GND.n2837 GND.n2836 585
R3224 GND.n2893 GND.n2837 585
R3225 GND.n3800 GND.n3799 585
R3226 GND.n3801 GND.n3800 585
R3227 GND.n2973 GND.n2972 585
R3228 GND.n2972 GND.n2901 585
R3229 GND.n3795 GND.n3794 585
R3230 GND.n3794 GND.n3793 585
R3231 GND.n2976 GND.n2975 585
R3232 GND.n2985 GND.n2976 585
R3233 GND.n3775 GND.n2995 585
R3234 GND.n2995 GND.n2982 585
R3235 GND.n3777 GND.n3776 585
R3236 GND.n3778 GND.n3777 585
R3237 GND.n2996 GND.n2994 585
R3238 GND.n3736 GND.n2994 585
R3239 GND.n3770 GND.n3769 585
R3240 GND.n3769 GND.n3768 585
R3241 GND.n2999 GND.n2998 585
R3242 GND.n3011 GND.n2999 585
R3243 GND.n3717 GND.n3716 585
R3244 GND.n3716 GND.n3009 585
R3245 GND.n3718 GND.n3031 585
R3246 GND.n3031 GND.n3023 585
R3247 GND.n3720 GND.n3719 585
R3248 GND.n3721 GND.n3720 585
R3249 GND.n3032 GND.n3030 585
R3250 GND.n3615 GND.n3030 585
R3251 GND.n3710 GND.n3709 585
R3252 GND.n3709 GND.n3708 585
R3253 GND.n3035 GND.n3034 585
R3254 GND.n3042 GND.n3035 585
R3255 GND.n3671 GND.n3060 585
R3256 GND.n3060 GND.n3053 585
R3257 GND.n3673 GND.n3672 585
R3258 GND.n3674 GND.n3673 585
R3259 GND.n3061 GND.n3059 585
R3260 GND.n3059 GND.n3057 585
R3261 GND.n3666 GND.n3665 585
R3262 GND.n3665 GND.n3664 585
R3263 GND.n3064 GND.n3063 585
R3264 GND.n3074 GND.n3064 585
R3265 GND.n3563 GND.n3562 585
R3266 GND.n3562 GND.n3072 585
R3267 GND.n3564 GND.n3557 585
R3268 GND.n3557 GND.n3079 585
R3269 GND.n3566 GND.n3565 585
R3270 GND.n3566 GND.n3083 585
R3271 GND.n3567 GND.n3556 585
R3272 GND.n3567 GND.n3091 585
R3273 GND.n3569 GND.n3568 585
R3274 GND.n3568 GND.n3089 585
R3275 GND.n3570 GND.n3106 585
R3276 GND.n3106 GND.n3097 585
R3277 GND.n3572 GND.n3571 585
R3278 GND.n3573 GND.n3572 585
R3279 GND.n3107 GND.n3105 585
R3280 GND.n3151 GND.n3105 585
R3281 GND.n3550 GND.n3549 585
R3282 GND.n3549 GND.n3548 585
R3283 GND.n3110 GND.n3109 585
R3284 GND.n3117 GND.n3110 585
R3285 GND.n3513 GND.n3136 585
R3286 GND.n3136 GND.n3129 585
R3287 GND.n3515 GND.n3514 585
R3288 GND.n3516 GND.n3515 585
R3289 GND.n3137 GND.n3135 585
R3290 GND.n3135 GND.n3133 585
R3291 GND.n3508 GND.n3507 585
R3292 GND.n3507 GND.n3506 585
R3293 GND.n3140 GND.n3139 585
R3294 GND.n3498 GND.n3140 585
R3295 GND.n3479 GND.n3478 585
R3296 GND.n3480 GND.n3479 585
R3297 GND.n3174 GND.n3173 585
R3298 GND.n3362 GND.n3173 585
R3299 GND.n3474 GND.n3473 585
R3300 GND.n3473 GND.n3472 585
R3301 GND.n3177 GND.n3176 585
R3302 GND.n3462 GND.n3177 585
R3303 GND.n3458 GND.n3457 585
R3304 GND.n3459 GND.n3458 585
R3305 GND.n3370 GND.n3369 585
R3306 GND.n3375 GND.n3369 585
R3307 GND.n3453 GND.n3452 585
R3308 GND.n3452 GND.n3451 585
R3309 GND.n3373 GND.n3372 585
R3310 GND.n3441 GND.n3373 585
R3311 GND.n3438 GND.n3437 585
R3312 GND.n3439 GND.n3438 585
R3313 GND.n3383 GND.n3382 585
R3314 GND.n3388 GND.n3382 585
R3315 GND.n3433 GND.n3432 585
R3316 GND.n3432 GND.n3431 585
R3317 GND.n3386 GND.n3385 585
R3318 GND.n3421 GND.n3386 585
R3319 GND.n3418 GND.n3417 585
R3320 GND.n3419 GND.n3418 585
R3321 GND.n3395 GND.n3394 585
R3322 GND.n3403 GND.n3394 585
R3323 GND.n3413 GND.n3412 585
R3324 GND.n3412 GND.n3411 585
R3325 GND.n3399 GND.n3398 585
R3326 GND.n3400 GND.n3399 585
R3327 GND.n1314 GND.n1313 585
R3328 GND.n1327 GND.n1314 585
R3329 GND.n4706 GND.n4705 585
R3330 GND.n4705 GND.n4704 585
R3331 GND.n4707 GND.n1308 585
R3332 GND.n1308 GND.n1306 585
R3333 GND.n4709 GND.n4708 585
R3334 GND.n4710 GND.n4709 585
R3335 GND.n1309 GND.n1307 585
R3336 GND.n1307 GND.n1295 585
R3337 GND.n2300 GND.n2299 585
R3338 GND.n2300 GND.n1238 585
R3339 GND.n2302 GND.n2301 585
R3340 GND.n2301 GND.n1236 585
R3341 GND.n2303 GND.n1422 585
R3342 GND.n1422 GND.n1402 585
R3343 GND.n2305 GND.n2304 585
R3344 GND.n2306 GND.n2305 585
R3345 GND.n1423 GND.n1421 585
R3346 GND.n1421 GND.n1412 585
R3347 GND.n2291 GND.n2290 585
R3348 GND.n2290 GND.n1410 585
R3349 GND.n2289 GND.n1425 585
R3350 GND.n2289 GND.n1414 585
R3351 GND.n2288 GND.n1427 585
R3352 GND.n2288 GND.n2287 585
R3353 GND.n2167 GND.n1426 585
R3354 GND.n1436 GND.n1426 585
R3355 GND.n2169 GND.n2168 585
R3356 GND.n2169 GND.n1434 585
R3357 GND.n2173 GND.n2172 585
R3358 GND.n2172 GND.n2171 585
R3359 GND.n2174 GND.n2159 585
R3360 GND.n2159 GND.n1446 585
R3361 GND.n2176 GND.n2175 585
R3362 GND.n2176 GND.n1445 585
R3363 GND.n2177 GND.n2158 585
R3364 GND.n2177 GND.n1458 585
R3365 GND.n2179 GND.n2178 585
R3366 GND.n2178 GND.n1455 585
R3367 GND.n2180 GND.n2153 585
R3368 GND.n2153 GND.n2152 585
R3369 GND.n2182 GND.n2181 585
R3370 GND.n2182 GND.n1468 585
R3371 GND.n2183 GND.n2150 585
R3372 GND.n2183 GND.n1467 585
R3373 GND.n2185 GND.n2184 585
R3374 GND.n2184 GND.n1478 585
R3375 GND.n2186 GND.n2145 585
R3376 GND.n2145 GND.n1476 585
R3377 GND.n2188 GND.n2187 585
R3378 GND.n2188 GND.n1481 585
R3379 GND.n2189 GND.n2144 585
R3380 GND.n2189 GND.n1490 585
R3381 GND.n2191 GND.n2190 585
R3382 GND.n2190 GND.n1488 585
R3383 GND.n2192 GND.n1505 585
R3384 GND.n1505 GND.n1500 585
R3385 GND.n2194 GND.n2193 585
R3386 GND.n2195 GND.n2194 585
R3387 GND.n1506 GND.n1504 585
R3388 GND.n1504 GND.n1502 585
R3389 GND.n2102 GND.n1559 585
R3390 GND.n2102 GND.n2101 585
R3391 GND.n2105 GND.n2104 585
R3392 GND.n2106 GND.n2105 585
R3393 GND.n2103 GND.n1558 585
R3394 GND.n1558 GND.n1552 585
R3395 GND.n1569 GND.n1568 585
R3396 GND.n1570 GND.n1569 585
R3397 GND.n1567 GND.n1541 585
R3398 GND.n1543 GND.n1541 585
R3399 GND.n2120 GND.n2119 585
R3400 GND.n2119 GND.n2118 585
R3401 GND.n2122 GND.n2121 585
R3402 GND.n2123 GND.n2122 585
R3403 GND.n1540 GND.n1539 585
R3404 GND.n1540 GND.n1534 585
R3405 GND.n1538 GND.n1537 585
R3406 GND.n1537 GND.n1528 585
R3407 GND.n1517 GND.n1515 585
R3408 GND.n1520 GND.n1517 585
R3409 GND.n2137 GND.n2136 585
R3410 GND.n2136 GND.n2135 585
R3411 GND.n1516 GND.n1514 585
R3412 GND.n1581 GND.n1516 585
R3413 GND.n2052 GND.n2051 585
R3414 GND.n2053 GND.n2052 585
R3415 GND.n1594 GND.n1593 585
R3416 GND.n1593 GND.n1591 585
R3417 GND.n2047 GND.n2046 585
R3418 GND.n2046 GND.n1589 585
R3419 GND.n2045 GND.n1596 585
R3420 GND.n2045 GND.n2044 585
R3421 GND.n2014 GND.n1597 585
R3422 GND.n1606 GND.n1597 585
R3423 GND.n2016 GND.n2015 585
R3424 GND.n2017 GND.n2016 585
R3425 GND.n1621 GND.n1620 585
R3426 GND.n1620 GND.n1617 585
R3427 GND.n2009 GND.n2008 585
R3428 GND.n2008 GND.n1615 585
R3429 GND.n2007 GND.n1623 585
R3430 GND.n2007 GND.n2006 585
R3431 GND.n1632 GND.n1631 585
R3432 GND.n1995 GND.n1632 585
R3433 GND.n1625 GND.n1624 585
R3434 GND.n1624 GND.n1131 585
R3435 GND.n1627 GND.n1626 585
R3436 GND.n1626 GND.n1128 585
R3437 GND.n1114 GND.n1113 585
R3438 GND.n1118 GND.n1114 585
R3439 GND.n4887 GND.n4886 585
R3440 GND.n4886 GND.n4885 585
R3441 GND.n3984 GND.n2427 585
R3442 GND.n4021 GND.n2427 585
R3443 GND.n4019 GND.n4018 585
R3444 GND.n3983 GND.n3982 585
R3445 GND.n4013 GND.n4012 585
R3446 GND.n4008 GND.n4007 585
R3447 GND.n4006 GND.n4005 585
R3448 GND.n3998 GND.n3986 585
R3449 GND.n4000 GND.n3999 585
R3450 GND.n3997 GND.n3995 585
R3451 GND.n3994 GND.n2478 585
R3452 GND.n4492 GND.n2477 585
R3453 GND.n4493 GND.n2476 585
R3454 GND.n3976 GND.n2470 585
R3455 GND.n4500 GND.n2469 585
R3456 GND.n4501 GND.n2468 585
R3457 GND.n3973 GND.n2462 585
R3458 GND.n4508 GND.n2461 585
R3459 GND.n4509 GND.n2460 585
R3460 GND.n3971 GND.n2454 585
R3461 GND.n4516 GND.n2453 585
R3462 GND.n4517 GND.n2452 585
R3463 GND.n3968 GND.n2446 585
R3464 GND.n4524 GND.n2445 585
R3465 GND.n4525 GND.n2444 585
R3466 GND.n3966 GND.n2437 585
R3467 GND.n4532 GND.n2436 585
R3468 GND.n4533 GND.n2431 585
R3469 GND.n4541 GND.n4540 585
R3470 GND.n4540 GND.n4539 585
R3471 GND.n4542 GND.n2426 585
R3472 GND.n3954 GND.n2426 585
R3473 GND.n2797 GND.n2424 585
R3474 GND.n3953 GND.n2797 585
R3475 GND.n4546 GND.n2423 585
R3476 GND.n2805 GND.n2423 585
R3477 GND.n4547 GND.n2422 585
R3478 GND.n3945 GND.n2422 585
R3479 GND.n4548 GND.n2421 585
R3480 GND.n3933 GND.n2421 585
R3481 GND.n2812 GND.n2419 585
R3482 GND.n3932 GND.n2812 585
R3483 GND.n4552 GND.n2418 585
R3484 GND.n2819 GND.n2418 585
R3485 GND.n4553 GND.n2417 585
R3486 GND.n3924 GND.n2417 585
R3487 GND.n4554 GND.n2416 585
R3488 GND.n3914 GND.n2416 585
R3489 GND.n2826 GND.n2414 585
R3490 GND.n3913 GND.n2826 585
R3491 GND.n4558 GND.n2413 585
R3492 GND.n2832 GND.n2413 585
R3493 GND.n4559 GND.n2412 585
R3494 GND.n3905 GND.n2412 585
R3495 GND.n4560 GND.n2411 585
R3496 GND.n3895 GND.n2411 585
R3497 GND.n2895 GND.n2409 585
R3498 GND.n3826 GND.n2895 585
R3499 GND.n4564 GND.n2408 585
R3500 GND.n3802 GND.n2408 585
R3501 GND.n4565 GND.n2407 585
R3502 GND.n3818 GND.n2407 585
R3503 GND.n4566 GND.n2406 585
R3504 GND.n3810 GND.n2406 585
R3505 GND.n2977 GND.n2404 585
R3506 GND.n2978 GND.n2977 585
R3507 GND.n4570 GND.n2403 585
R3508 GND.n2983 GND.n2403 585
R3509 GND.n4571 GND.n2402 585
R3510 GND.n2993 GND.n2402 585
R3511 GND.n4572 GND.n2401 585
R3512 GND.n2990 GND.n2401 585
R3513 GND.n3000 GND.n2399 585
R3514 GND.n3767 GND.n3000 585
R3515 GND.n4576 GND.n2398 585
R3516 GND.n3017 GND.n2398 585
R3517 GND.n4577 GND.n2397 585
R3518 GND.n3749 GND.n2397 585
R3519 GND.n4578 GND.n2396 585
R3520 GND.n3729 GND.n2396 585
R3521 GND.n3690 GND.n2394 585
R3522 GND.n3691 GND.n3690 585
R3523 GND.n4582 GND.n2393 585
R3524 GND.n3027 GND.n2393 585
R3525 GND.n4583 GND.n2392 585
R3526 GND.n3038 GND.n2392 585
R3527 GND.n4584 GND.n2391 585
R3528 GND.n3700 GND.n2391 585
R3529 GND.n3623 GND.n2389 585
R3530 GND.n3624 GND.n3623 585
R3531 GND.n4588 GND.n2388 585
R3532 GND.n3683 GND.n2388 585
R3533 GND.n4589 GND.n2387 585
R3534 GND.n3675 GND.n2387 585
R3535 GND.n4590 GND.n2386 585
R3536 GND.n3663 GND.n2386 585
R3537 GND.n3635 GND.n2384 585
R3538 GND.n3636 GND.n3635 585
R3539 GND.n4594 GND.n2383 585
R3540 GND.n3655 GND.n2383 585
R3541 GND.n4595 GND.n2382 585
R3542 GND.n3644 GND.n2382 585
R3543 GND.n4596 GND.n2381 585
R3544 GND.n3606 GND.n2381 585
R3545 GND.n3589 GND.n2379 585
R3546 GND.n3590 GND.n3589 585
R3547 GND.n4600 GND.n2378 585
R3548 GND.n3598 GND.n2378 585
R3549 GND.n4601 GND.n2377 585
R3550 GND.n3581 GND.n2377 585
R3551 GND.n4602 GND.n2376 585
R3552 GND.n3104 GND.n2376 585
R3553 GND.n3101 GND.n2374 585
R3554 GND.n3102 GND.n3101 585
R3555 GND.n4606 GND.n2373 585
R3556 GND.n3113 GND.n2373 585
R3557 GND.n4607 GND.n2372 585
R3558 GND.n3540 GND.n2372 585
R3559 GND.n4608 GND.n2371 585
R3560 GND.n3159 GND.n2371 585
R3561 GND.n3127 GND.n2369 585
R3562 GND.n3525 GND.n3127 585
R3563 GND.n4612 GND.n2368 585
R3564 GND.n3517 GND.n2368 585
R3565 GND.n4613 GND.n2367 585
R3566 GND.n3490 GND.n2367 585
R3567 GND.n4614 GND.n2366 585
R3568 GND.n3141 GND.n2366 585
R3569 GND.n3481 GND.n2364 585
R3570 GND.n3482 GND.n3481 585
R3571 GND.n4618 GND.n2363 585
R3572 GND.n3180 GND.n2363 585
R3573 GND.n4619 GND.n2362 585
R3574 GND.n3471 GND.n2362 585
R3575 GND.n4620 GND.n2361 585
R3576 GND.n3461 GND.n2361 585
R3577 GND.n3460 GND.n2359 585
R3578 GND.n3463 GND.n3460 585
R3579 GND.n4624 GND.n2358 585
R3580 GND.n3368 GND.n2358 585
R3581 GND.n4625 GND.n2357 585
R3582 GND.n3450 GND.n2357 585
R3583 GND.n4626 GND.n2356 585
R3584 GND.n3374 GND.n2356 585
R3585 GND.n3440 GND.n2354 585
R3586 GND.n3442 GND.n3440 585
R3587 GND.n4630 GND.n2353 585
R3588 GND.n3381 GND.n2353 585
R3589 GND.n4631 GND.n2352 585
R3590 GND.n3430 GND.n2352 585
R3591 GND.n4632 GND.n2351 585
R3592 GND.n3387 GND.n2351 585
R3593 GND.n3420 GND.n2349 585
R3594 GND.n3422 GND.n3420 585
R3595 GND.n4636 GND.n2348 585
R3596 GND.n3402 GND.n2348 585
R3597 GND.n4637 GND.n2347 585
R3598 GND.n3410 GND.n2347 585
R3599 GND.n4638 GND.n2346 585
R3600 GND.n3401 GND.n2346 585
R3601 GND.n4701 GND.n4700 585
R3602 GND.n4699 GND.n1329 585
R3603 GND.n1332 GND.n1328 585
R3604 GND.n4703 GND.n1328 585
R3605 GND.n4692 GND.n1341 585
R3606 GND.n4691 GND.n1342 585
R3607 GND.n1344 GND.n1343 585
R3608 GND.n4684 GND.n1350 585
R3609 GND.n4683 GND.n1351 585
R3610 GND.n1360 GND.n1352 585
R3611 GND.n4676 GND.n1361 585
R3612 GND.n4675 GND.n1362 585
R3613 GND.n1364 GND.n1363 585
R3614 GND.n4668 GND.n1370 585
R3615 GND.n4667 GND.n1371 585
R3616 GND.n1380 GND.n1372 585
R3617 GND.n4660 GND.n1381 585
R3618 GND.n4659 GND.n1382 585
R3619 GND.n1384 GND.n1383 585
R3620 GND.n1394 GND.n1393 585
R3621 GND.n4650 GND.n1395 585
R3622 GND.n4649 GND.n1396 585
R3623 GND.n4648 GND.n1397 585
R3624 GND.n2339 GND.n1398 585
R3625 GND.n4644 GND.n2340 585
R3626 GND.n4643 GND.n2341 585
R3627 GND.n4642 GND.n2342 585
R3628 GND.n2345 GND.n2343 585
R3629 GND.n4538 GND.n4537 585
R3630 GND.n4539 GND.n4538 585
R3631 GND.n2432 GND.n2430 585
R3632 GND.n3954 GND.n2430 585
R3633 GND.n3952 GND.n3951 585
R3634 GND.n3953 GND.n3952 585
R3635 GND.n2799 GND.n2798 585
R3636 GND.n2805 GND.n2798 585
R3637 GND.n3947 GND.n3946 585
R3638 GND.n3946 GND.n3945 585
R3639 GND.n2802 GND.n2801 585
R3640 GND.n3933 GND.n2802 585
R3641 GND.n3931 GND.n3930 585
R3642 GND.n3932 GND.n3931 585
R3643 GND.n2814 GND.n2813 585
R3644 GND.n2819 GND.n2813 585
R3645 GND.n3926 GND.n3925 585
R3646 GND.n3925 GND.n3924 585
R3647 GND.n2817 GND.n2816 585
R3648 GND.n3914 GND.n2817 585
R3649 GND.n3912 GND.n3911 585
R3650 GND.n3913 GND.n3912 585
R3651 GND.n2828 GND.n2827 585
R3652 GND.n2832 GND.n2827 585
R3653 GND.n3907 GND.n3906 585
R3654 GND.n3906 GND.n3905 585
R3655 GND.n2831 GND.n2830 585
R3656 GND.n3895 GND.n2831 585
R3657 GND.n3825 GND.n3824 585
R3658 GND.n3826 GND.n3825 585
R3659 GND.n2897 GND.n2896 585
R3660 GND.n3802 GND.n2896 585
R3661 GND.n3820 GND.n3819 585
R3662 GND.n3819 GND.n3818 585
R3663 GND.n2900 GND.n2899 585
R3664 GND.n3810 GND.n2900 585
R3665 GND.n3759 GND.n3757 585
R3666 GND.n3757 GND.n2978 585
R3667 GND.n3760 GND.n3756 585
R3668 GND.n3756 GND.n2983 585
R3669 GND.n3761 GND.n3755 585
R3670 GND.n3755 GND.n2993 585
R3671 GND.n3005 GND.n3003 585
R3672 GND.n3003 GND.n2990 585
R3673 GND.n3766 GND.n3765 585
R3674 GND.n3767 GND.n3766 585
R3675 GND.n3004 GND.n3002 585
R3676 GND.n3017 GND.n3002 585
R3677 GND.n3751 GND.n3750 585
R3678 GND.n3750 GND.n3749 585
R3679 GND.n3008 GND.n3007 585
R3680 GND.n3729 GND.n3008 585
R3681 GND.n3693 GND.n3692 585
R3682 GND.n3692 GND.n3691 585
R3683 GND.n3694 GND.n3689 585
R3684 GND.n3689 GND.n3027 585
R3685 GND.n3047 GND.n3045 585
R3686 GND.n3045 GND.n3038 585
R3687 GND.n3699 GND.n3698 585
R3688 GND.n3700 GND.n3699 585
R3689 GND.n3046 GND.n3044 585
R3690 GND.n3624 GND.n3044 585
R3691 GND.n3685 GND.n3684 585
R3692 GND.n3684 GND.n3683 585
R3693 GND.n3050 GND.n3049 585
R3694 GND.n3675 GND.n3050 585
R3695 GND.n3662 GND.n3661 585
R3696 GND.n3663 GND.n3662 585
R3697 GND.n3068 GND.n3067 585
R3698 GND.n3636 GND.n3067 585
R3699 GND.n3657 GND.n3656 585
R3700 GND.n3656 GND.n3655 585
R3701 GND.n3071 GND.n3070 585
R3702 GND.n3644 GND.n3071 585
R3703 GND.n3605 GND.n3604 585
R3704 GND.n3606 GND.n3605 585
R3705 GND.n3085 GND.n3084 585
R3706 GND.n3590 GND.n3084 585
R3707 GND.n3600 GND.n3599 585
R3708 GND.n3599 GND.n3598 585
R3709 GND.n3088 GND.n3087 585
R3710 GND.n3581 GND.n3088 585
R3711 GND.n3533 GND.n3532 585
R3712 GND.n3532 GND.n3104 585
R3713 GND.n3534 GND.n3531 585
R3714 GND.n3531 GND.n3102 585
R3715 GND.n3122 GND.n3120 585
R3716 GND.n3120 GND.n3113 585
R3717 GND.n3539 GND.n3538 585
R3718 GND.n3540 GND.n3539 585
R3719 GND.n3121 GND.n3119 585
R3720 GND.n3159 GND.n3119 585
R3721 GND.n3527 GND.n3526 585
R3722 GND.n3526 GND.n3525 585
R3723 GND.n3125 GND.n3124 585
R3724 GND.n3517 GND.n3125 585
R3725 GND.n3489 GND.n3488 585
R3726 GND.n3490 GND.n3489 585
R3727 GND.n3168 GND.n3167 585
R3728 GND.n3167 GND.n3141 585
R3729 GND.n3484 GND.n3483 585
R3730 GND.n3483 GND.n3482 585
R3731 GND.n3171 GND.n3170 585
R3732 GND.n3180 GND.n3171 585
R3733 GND.n3470 GND.n3469 585
R3734 GND.n3471 GND.n3470 585
R3735 GND.n3364 GND.n3363 585
R3736 GND.n3461 GND.n3363 585
R3737 GND.n3465 GND.n3464 585
R3738 GND.n3464 GND.n3463 585
R3739 GND.n3367 GND.n3366 585
R3740 GND.n3368 GND.n3367 585
R3741 GND.n3449 GND.n3448 585
R3742 GND.n3450 GND.n3449 585
R3743 GND.n3377 GND.n3376 585
R3744 GND.n3376 GND.n3374 585
R3745 GND.n3444 GND.n3443 585
R3746 GND.n3443 GND.n3442 585
R3747 GND.n3380 GND.n3379 585
R3748 GND.n3381 GND.n3380 585
R3749 GND.n3429 GND.n3428 585
R3750 GND.n3430 GND.n3429 585
R3751 GND.n3390 GND.n3389 585
R3752 GND.n3389 GND.n3387 585
R3753 GND.n3424 GND.n3423 585
R3754 GND.n3423 GND.n3422 585
R3755 GND.n3393 GND.n3392 585
R3756 GND.n3402 GND.n3393 585
R3757 GND.n3409 GND.n3408 585
R3758 GND.n3410 GND.n3409 585
R3759 GND.n3404 GND.n1330 585
R3760 GND.n3401 GND.n1330 585
R3761 GND.n5030 GND.n5029 555.492
R3762 GND.n3892 GND.n2870 521.33
R3763 GND.n2969 GND.n2968 521.33
R3764 GND.n3240 GND.n3179 521.33
R3765 GND.n3360 GND.n3181 521.33
R3766 GND.n3220 GND.t18 347.526
R3767 GND.n2908 GND.t28 347.526
R3768 GND.n3216 GND.t7 347.526
R3769 GND.n3832 GND.t60 347.526
R3770 GND.n1264 GND.t51 291.267
R3771 GND.n1292 GND.t11 291.267
R3772 GND.n4486 GND.t35 291.267
R3773 GND.n1387 GND.t32 291.267
R3774 GND.n1802 GND.t86 291.267
R3775 GND.n2539 GND.t0 291.267
R3776 GND.n2561 GND.t42 291.267
R3777 GND.n541 GND.t38 291.267
R3778 GND.n5796 GND.t89 291.267
R3779 GND.n575 GND.t76 291.267
R3780 GND.n1727 GND.t24 291.267
R3781 GND.n1759 GND.t57 291.267
R3782 GND.n151 GND.n125 289.615
R3783 GND.n119 GND.n93 289.615
R3784 GND.n87 GND.n61 289.615
R3785 GND.n56 GND.n30 289.615
R3786 GND.n278 GND.n252 289.615
R3787 GND.n246 GND.n220 289.615
R3788 GND.n214 GND.n188 289.615
R3789 GND.n183 GND.n157 289.615
R3790 GND.n5031 GND.n5030 280.613
R3791 GND.n5031 GND.n967 280.613
R3792 GND.n5039 GND.n967 280.613
R3793 GND.n5040 GND.n5039 280.613
R3794 GND.n5041 GND.n5040 280.613
R3795 GND.n5041 GND.n961 280.613
R3796 GND.n5049 GND.n961 280.613
R3797 GND.n5050 GND.n5049 280.613
R3798 GND.n5051 GND.n5050 280.613
R3799 GND.n5051 GND.n955 280.613
R3800 GND.n5059 GND.n955 280.613
R3801 GND.n5060 GND.n5059 280.613
R3802 GND.n5061 GND.n5060 280.613
R3803 GND.n5061 GND.n949 280.613
R3804 GND.n5069 GND.n949 280.613
R3805 GND.n5070 GND.n5069 280.613
R3806 GND.n5071 GND.n5070 280.613
R3807 GND.n5071 GND.n943 280.613
R3808 GND.n5079 GND.n943 280.613
R3809 GND.n5080 GND.n5079 280.613
R3810 GND.n5081 GND.n5080 280.613
R3811 GND.n5081 GND.n937 280.613
R3812 GND.n5089 GND.n937 280.613
R3813 GND.n5090 GND.n5089 280.613
R3814 GND.n5091 GND.n5090 280.613
R3815 GND.n5091 GND.n931 280.613
R3816 GND.n5099 GND.n931 280.613
R3817 GND.n5100 GND.n5099 280.613
R3818 GND.n5101 GND.n5100 280.613
R3819 GND.n5101 GND.n925 280.613
R3820 GND.n5109 GND.n925 280.613
R3821 GND.n5110 GND.n5109 280.613
R3822 GND.n5111 GND.n5110 280.613
R3823 GND.n5111 GND.n919 280.613
R3824 GND.n5119 GND.n919 280.613
R3825 GND.n5120 GND.n5119 280.613
R3826 GND.n5121 GND.n5120 280.613
R3827 GND.n5121 GND.n913 280.613
R3828 GND.n5129 GND.n913 280.613
R3829 GND.n5130 GND.n5129 280.613
R3830 GND.n5131 GND.n5130 280.613
R3831 GND.n5131 GND.n907 280.613
R3832 GND.n5139 GND.n907 280.613
R3833 GND.n5140 GND.n5139 280.613
R3834 GND.n5141 GND.n5140 280.613
R3835 GND.n5141 GND.n901 280.613
R3836 GND.n5149 GND.n901 280.613
R3837 GND.n5150 GND.n5149 280.613
R3838 GND.n5151 GND.n5150 280.613
R3839 GND.n5151 GND.n895 280.613
R3840 GND.n5159 GND.n895 280.613
R3841 GND.n5160 GND.n5159 280.613
R3842 GND.n5161 GND.n5160 280.613
R3843 GND.n5161 GND.n889 280.613
R3844 GND.n5169 GND.n889 280.613
R3845 GND.n5170 GND.n5169 280.613
R3846 GND.n5171 GND.n5170 280.613
R3847 GND.n5171 GND.n883 280.613
R3848 GND.n5179 GND.n883 280.613
R3849 GND.n5180 GND.n5179 280.613
R3850 GND.n5181 GND.n5180 280.613
R3851 GND.n5181 GND.n877 280.613
R3852 GND.n5189 GND.n877 280.613
R3853 GND.n5190 GND.n5189 280.613
R3854 GND.n5191 GND.n5190 280.613
R3855 GND.n5191 GND.n871 280.613
R3856 GND.n5199 GND.n871 280.613
R3857 GND.n5200 GND.n5199 280.613
R3858 GND.n5201 GND.n5200 280.613
R3859 GND.n5201 GND.n865 280.613
R3860 GND.n5209 GND.n865 280.613
R3861 GND.n5210 GND.n5209 280.613
R3862 GND.n5211 GND.n5210 280.613
R3863 GND.n5211 GND.n859 280.613
R3864 GND.n5219 GND.n859 280.613
R3865 GND.n5220 GND.n5219 280.613
R3866 GND.n5221 GND.n5220 280.613
R3867 GND.n5221 GND.n853 280.613
R3868 GND.n5229 GND.n853 280.613
R3869 GND.n5230 GND.n5229 280.613
R3870 GND.n5231 GND.n5230 280.613
R3871 GND.n5231 GND.n847 280.613
R3872 GND.n5239 GND.n847 280.613
R3873 GND.n5240 GND.n5239 280.613
R3874 GND.n5241 GND.n5240 280.613
R3875 GND.n5241 GND.n841 280.613
R3876 GND.n5249 GND.n841 280.613
R3877 GND.n5250 GND.n5249 280.613
R3878 GND.n5251 GND.n5250 280.613
R3879 GND.n5251 GND.n835 280.613
R3880 GND.n5259 GND.n835 280.613
R3881 GND.n5260 GND.n5259 280.613
R3882 GND.n5261 GND.n5260 280.613
R3883 GND.n5261 GND.n829 280.613
R3884 GND.n5269 GND.n829 280.613
R3885 GND.n5270 GND.n5269 280.613
R3886 GND.n5271 GND.n5270 280.613
R3887 GND.n5271 GND.n823 280.613
R3888 GND.n5279 GND.n823 280.613
R3889 GND.n5280 GND.n5279 280.613
R3890 GND.n5281 GND.n5280 280.613
R3891 GND.n5281 GND.n817 280.613
R3892 GND.n5289 GND.n817 280.613
R3893 GND.n5290 GND.n5289 280.613
R3894 GND.n5291 GND.n5290 280.613
R3895 GND.n5291 GND.n811 280.613
R3896 GND.n5299 GND.n811 280.613
R3897 GND.n5300 GND.n5299 280.613
R3898 GND.n5301 GND.n5300 280.613
R3899 GND.n5301 GND.n805 280.613
R3900 GND.n5309 GND.n805 280.613
R3901 GND.n5310 GND.n5309 280.613
R3902 GND.n5311 GND.n5310 280.613
R3903 GND.n5311 GND.n799 280.613
R3904 GND.n5319 GND.n799 280.613
R3905 GND.n5320 GND.n5319 280.613
R3906 GND.n5321 GND.n5320 280.613
R3907 GND.n5321 GND.n793 280.613
R3908 GND.n5329 GND.n793 280.613
R3909 GND.n5330 GND.n5329 280.613
R3910 GND.n5331 GND.n5330 280.613
R3911 GND.n5331 GND.n787 280.613
R3912 GND.n5339 GND.n787 280.613
R3913 GND.n5340 GND.n5339 280.613
R3914 GND.n5341 GND.n5340 280.613
R3915 GND.n5341 GND.n781 280.613
R3916 GND.n5349 GND.n781 280.613
R3917 GND.n5350 GND.n5349 280.613
R3918 GND.n5351 GND.n5350 280.613
R3919 GND.n5351 GND.n775 280.613
R3920 GND.n5359 GND.n775 280.613
R3921 GND.n5360 GND.n5359 280.613
R3922 GND.n5361 GND.n5360 280.613
R3923 GND.n5361 GND.n769 280.613
R3924 GND.n5369 GND.n769 280.613
R3925 GND.n5370 GND.n5369 280.613
R3926 GND.n5371 GND.n5370 280.613
R3927 GND.n5371 GND.n763 280.613
R3928 GND.n5379 GND.n763 280.613
R3929 GND.n5380 GND.n5379 280.613
R3930 GND.n5381 GND.n5380 280.613
R3931 GND.n5381 GND.n757 280.613
R3932 GND.n5389 GND.n757 280.613
R3933 GND.n5390 GND.n5389 280.613
R3934 GND.n5391 GND.n5390 280.613
R3935 GND.n5391 GND.n751 280.613
R3936 GND.n5399 GND.n751 280.613
R3937 GND.n5400 GND.n5399 280.613
R3938 GND.n5401 GND.n5400 280.613
R3939 GND.n5401 GND.n745 280.613
R3940 GND.n5409 GND.n745 280.613
R3941 GND.n5410 GND.n5409 280.613
R3942 GND.n5411 GND.n5410 280.613
R3943 GND.n5411 GND.n739 280.613
R3944 GND.n5419 GND.n739 280.613
R3945 GND.n5420 GND.n5419 280.613
R3946 GND.n5421 GND.n5420 280.613
R3947 GND.n5421 GND.n733 280.613
R3948 GND.n5429 GND.n733 280.613
R3949 GND.n5430 GND.n5429 280.613
R3950 GND.n5431 GND.n5430 280.613
R3951 GND.n5431 GND.n727 280.613
R3952 GND.n5439 GND.n727 280.613
R3953 GND.n5440 GND.n5439 280.613
R3954 GND.n5441 GND.n5440 280.613
R3955 GND.n5441 GND.n721 280.613
R3956 GND.n5449 GND.n721 280.613
R3957 GND.n5450 GND.n5449 280.613
R3958 GND.n5451 GND.n5450 280.613
R3959 GND.n5451 GND.n715 280.613
R3960 GND.n5459 GND.n715 280.613
R3961 GND.n5460 GND.n5459 280.613
R3962 GND.n5461 GND.n5460 280.613
R3963 GND.n5461 GND.n709 280.613
R3964 GND.n5469 GND.n709 280.613
R3965 GND.n5470 GND.n5469 280.613
R3966 GND.n5471 GND.n5470 280.613
R3967 GND.n5471 GND.n703 280.613
R3968 GND.n5480 GND.n703 280.613
R3969 GND.n5481 GND.n5480 280.613
R3970 GND.n2336 GND.t69 279.217
R3971 GND.n4009 GND.t79 279.217
R3972 GND.n3188 GND.t56 260.649
R3973 GND.n2883 GND.t75 260.649
R3974 GND.n3354 GND.n3178 256.663
R3975 GND.n3203 GND.n3178 256.663
R3976 GND.n3347 GND.n3178 256.663
R3977 GND.n3341 GND.n3178 256.663
R3978 GND.n3339 GND.n3178 256.663
R3979 GND.n3333 GND.n3178 256.663
R3980 GND.n3331 GND.n3178 256.663
R3981 GND.n3325 GND.n3178 256.663
R3982 GND.n3323 GND.n3178 256.663
R3983 GND.n3317 GND.n3178 256.663
R3984 GND.n3315 GND.n3178 256.663
R3985 GND.n3309 GND.n3178 256.663
R3986 GND.n3307 GND.n3178 256.663
R3987 GND.n3301 GND.n3178 256.663
R3988 GND.n3299 GND.n3178 256.663
R3989 GND.n3298 GND.n1267 256.663
R3990 GND.n3297 GND.n3178 256.663
R3991 GND.n3291 GND.n3178 256.663
R3992 GND.n3223 GND.n3178 256.663
R3993 GND.n3285 GND.n3178 256.663
R3994 GND.n3279 GND.n3178 256.663
R3995 GND.n3277 GND.n3178 256.663
R3996 GND.n3271 GND.n3178 256.663
R3997 GND.n3269 GND.n3178 256.663
R3998 GND.n3263 GND.n3178 256.663
R3999 GND.n3261 GND.n3178 256.663
R4000 GND.n3255 GND.n3178 256.663
R4001 GND.n3253 GND.n3178 256.663
R4002 GND.n3247 GND.n3178 256.663
R4003 GND.n3245 GND.n3178 256.663
R4004 GND.n3239 GND.n3178 256.663
R4005 GND.n3893 GND.n2839 256.663
R4006 GND.n3893 GND.n2840 256.663
R4007 GND.n3893 GND.n2841 256.663
R4008 GND.n3893 GND.n2842 256.663
R4009 GND.n3893 GND.n2843 256.663
R4010 GND.n3893 GND.n2844 256.663
R4011 GND.n3893 GND.n2845 256.663
R4012 GND.n3893 GND.n2846 256.663
R4013 GND.n3893 GND.n2847 256.663
R4014 GND.n3893 GND.n2848 256.663
R4015 GND.n3893 GND.n2849 256.663
R4016 GND.n3893 GND.n2850 256.663
R4017 GND.n3893 GND.n2851 256.663
R4018 GND.n3893 GND.n2852 256.663
R4019 GND.n3893 GND.n2853 256.663
R4020 GND.n2854 GND.n2536 256.663
R4021 GND.n3893 GND.n2855 256.663
R4022 GND.n3893 GND.n2856 256.663
R4023 GND.n3893 GND.n2857 256.663
R4024 GND.n3893 GND.n2858 256.663
R4025 GND.n3893 GND.n2859 256.663
R4026 GND.n3893 GND.n2860 256.663
R4027 GND.n3893 GND.n2861 256.663
R4028 GND.n3893 GND.n2862 256.663
R4029 GND.n3893 GND.n2863 256.663
R4030 GND.n3893 GND.n2864 256.663
R4031 GND.n3893 GND.n2865 256.663
R4032 GND.n3893 GND.n2866 256.663
R4033 GND.n3893 GND.n2867 256.663
R4034 GND.n3893 GND.n2868 256.663
R4035 GND.n3893 GND.n2869 256.663
R4036 GND.n1830 GND.n1696 242.672
R4037 GND.n1770 GND.n1696 242.672
R4038 GND.n1775 GND.n1696 242.672
R4039 GND.n1780 GND.n1696 242.672
R4040 GND.n1783 GND.n1696 242.672
R4041 GND.n1788 GND.n1696 242.672
R4042 GND.n1791 GND.n1696 242.672
R4043 GND.n1796 GND.n1696 242.672
R4044 GND.n1800 GND.n1696 242.672
R4045 GND.n4737 GND.n1305 242.672
R4046 GND.n4737 GND.n1304 242.672
R4047 GND.n4737 GND.n1303 242.672
R4048 GND.n4737 GND.n1302 242.672
R4049 GND.n4737 GND.n1301 242.672
R4050 GND.n4737 GND.n1300 242.672
R4051 GND.n4737 GND.n1299 242.672
R4052 GND.n4737 GND.n1298 242.672
R4053 GND.n4737 GND.n1297 242.672
R4054 GND.n4483 GND.n2503 242.672
R4055 GND.n4483 GND.n2505 242.672
R4056 GND.n4483 GND.n2506 242.672
R4057 GND.n4483 GND.n2508 242.672
R4058 GND.n4483 GND.n2510 242.672
R4059 GND.n4483 GND.n2511 242.672
R4060 GND.n4483 GND.n2513 242.672
R4061 GND.n4483 GND.n2515 242.672
R4062 GND.n4484 GND.n4483 242.672
R4063 GND.n572 GND.n471 242.672
R4064 GND.n5730 GND.n471 242.672
R4065 GND.n568 GND.n471 242.672
R4066 GND.n5737 GND.n471 242.672
R4067 GND.n561 GND.n471 242.672
R4068 GND.n5744 GND.n471 242.672
R4069 GND.n554 GND.n471 242.672
R4070 GND.n5751 GND.n471 242.672
R4071 GND.n547 GND.n471 242.672
R4072 GND.n1909 GND.n1696 242.672
R4073 GND.n1703 GND.n1696 242.672
R4074 GND.n1902 GND.n1696 242.672
R4075 GND.n1896 GND.n1696 242.672
R4076 GND.n1894 GND.n1696 242.672
R4077 GND.n1888 GND.n1696 242.672
R4078 GND.n1886 GND.n1696 242.672
R4079 GND.n1880 GND.n1696 242.672
R4080 GND.n1878 GND.n1696 242.672
R4081 GND.n1872 GND.n1696 242.672
R4082 GND.n1870 GND.n1696 242.672
R4083 GND.n1864 GND.n1696 242.672
R4084 GND.n1862 GND.n1696 242.672
R4085 GND.n1856 GND.n1696 242.672
R4086 GND.n1854 GND.n1696 242.672
R4087 GND.n1848 GND.n1696 242.672
R4088 GND.n1846 GND.n1696 242.672
R4089 GND.n1757 GND.n1696 242.672
R4090 GND.n1836 GND.n1696 242.672
R4091 GND.n4738 GND.n4737 242.672
R4092 GND.n4737 GND.n4711 242.672
R4093 GND.n4737 GND.n4712 242.672
R4094 GND.n4737 GND.n4714 242.672
R4095 GND.n4737 GND.n4715 242.672
R4096 GND.n4737 GND.n4717 242.672
R4097 GND.n4737 GND.n4718 242.672
R4098 GND.n4737 GND.n4720 242.672
R4099 GND.n4737 GND.n4721 242.672
R4100 GND.n4737 GND.n4723 242.672
R4101 GND.n4737 GND.n4724 242.672
R4102 GND.n4771 GND.n1266 242.672
R4103 GND.n4737 GND.n4726 242.672
R4104 GND.n4737 GND.n4727 242.672
R4105 GND.n4737 GND.n4729 242.672
R4106 GND.n4737 GND.n4730 242.672
R4107 GND.n4737 GND.n4732 242.672
R4108 GND.n4737 GND.n4733 242.672
R4109 GND.n4737 GND.n4735 242.672
R4110 GND.n4737 GND.n4736 242.672
R4111 GND.n4483 GND.n4482 242.672
R4112 GND.n4483 GND.n2485 242.672
R4113 GND.n4483 GND.n2486 242.672
R4114 GND.n4483 GND.n2487 242.672
R4115 GND.n4483 GND.n2488 242.672
R4116 GND.n4483 GND.n2489 242.672
R4117 GND.n4483 GND.n2490 242.672
R4118 GND.n4483 GND.n2491 242.672
R4119 GND.n4451 GND.n2537 242.672
R4120 GND.n4483 GND.n2492 242.672
R4121 GND.n4483 GND.n2493 242.672
R4122 GND.n4483 GND.n2494 242.672
R4123 GND.n4483 GND.n2495 242.672
R4124 GND.n4483 GND.n2496 242.672
R4125 GND.n4483 GND.n2497 242.672
R4126 GND.n4483 GND.n2498 242.672
R4127 GND.n4483 GND.n2499 242.672
R4128 GND.n4483 GND.n2500 242.672
R4129 GND.n4483 GND.n2501 242.672
R4130 GND.n4483 GND.n2502 242.672
R4131 GND.n538 GND.n471 242.672
R4132 GND.n5764 GND.n471 242.672
R4133 GND.n534 GND.n471 242.672
R4134 GND.n5771 GND.n471 242.672
R4135 GND.n527 GND.n471 242.672
R4136 GND.n5778 GND.n471 242.672
R4137 GND.n520 GND.n471 242.672
R4138 GND.n5785 GND.n471 242.672
R4139 GND.n513 GND.n471 242.672
R4140 GND.n5792 GND.n471 242.672
R4141 GND.n506 GND.n471 242.672
R4142 GND.n5802 GND.n471 242.672
R4143 GND.n499 GND.n471 242.672
R4144 GND.n5809 GND.n471 242.672
R4145 GND.n492 GND.n471 242.672
R4146 GND.n5816 GND.n471 242.672
R4147 GND.n485 GND.n471 242.672
R4148 GND.n5823 GND.n471 242.672
R4149 GND.n478 GND.n471 242.672
R4150 GND.n4021 GND.n4020 242.672
R4151 GND.n4021 GND.n3981 242.672
R4152 GND.n4021 GND.n3980 242.672
R4153 GND.n4021 GND.n3979 242.672
R4154 GND.n4021 GND.n3978 242.672
R4155 GND.n4021 GND.n3977 242.672
R4156 GND.n4021 GND.n3975 242.672
R4157 GND.n4021 GND.n3974 242.672
R4158 GND.n4021 GND.n3972 242.672
R4159 GND.n4021 GND.n3970 242.672
R4160 GND.n4021 GND.n3969 242.672
R4161 GND.n4021 GND.n3967 242.672
R4162 GND.n4021 GND.n3965 242.672
R4163 GND.n4703 GND.n4702 242.672
R4164 GND.n4703 GND.n1315 242.672
R4165 GND.n4703 GND.n1316 242.672
R4166 GND.n4703 GND.n1317 242.672
R4167 GND.n4703 GND.n1318 242.672
R4168 GND.n4703 GND.n1319 242.672
R4169 GND.n4703 GND.n1320 242.672
R4170 GND.n4703 GND.n1321 242.672
R4171 GND.n4703 GND.n1322 242.672
R4172 GND.n4703 GND.n1323 242.672
R4173 GND.n4703 GND.n1324 242.672
R4174 GND.n4703 GND.n1325 242.672
R4175 GND.n4703 GND.n1326 242.672
R4176 GND.n475 GND.n472 240.244
R4177 GND.n5825 GND.n5824 240.244
R4178 GND.n5822 GND.n479 240.244
R4179 GND.n5818 GND.n5817 240.244
R4180 GND.n5815 GND.n486 240.244
R4181 GND.n5811 GND.n5810 240.244
R4182 GND.n5808 GND.n493 240.244
R4183 GND.n5804 GND.n5803 240.244
R4184 GND.n5801 GND.n500 240.244
R4185 GND.n5794 GND.n5793 240.244
R4186 GND.n5791 GND.n507 240.244
R4187 GND.n5787 GND.n5786 240.244
R4188 GND.n5784 GND.n514 240.244
R4189 GND.n5780 GND.n5779 240.244
R4190 GND.n5777 GND.n521 240.244
R4191 GND.n5773 GND.n5772 240.244
R4192 GND.n5770 GND.n528 240.244
R4193 GND.n5766 GND.n5765 240.244
R4194 GND.n5763 GND.n535 240.244
R4195 GND.n4408 GND.n2564 240.244
R4196 GND.n4400 GND.n2564 240.244
R4197 GND.n4400 GND.n2575 240.244
R4198 GND.n2591 GND.n2575 240.244
R4199 GND.n4117 GND.n2591 240.244
R4200 GND.n4117 GND.n2604 240.244
R4201 GND.n4122 GND.n2604 240.244
R4202 GND.n4122 GND.n2615 240.244
R4203 GND.n4132 GND.n2615 240.244
R4204 GND.n4132 GND.n2625 240.244
R4205 GND.n4137 GND.n2625 240.244
R4206 GND.n4137 GND.n2636 240.244
R4207 GND.n4147 GND.n2636 240.244
R4208 GND.n4147 GND.n2646 240.244
R4209 GND.n4152 GND.n2646 240.244
R4210 GND.n4152 GND.n2656 240.244
R4211 GND.n4162 GND.n2656 240.244
R4212 GND.n4162 GND.n2666 240.244
R4213 GND.n4167 GND.n2666 240.244
R4214 GND.n4167 GND.n2677 240.244
R4215 GND.n4177 GND.n2677 240.244
R4216 GND.n4177 GND.n2687 240.244
R4217 GND.n4182 GND.n2687 240.244
R4218 GND.n4182 GND.n2698 240.244
R4219 GND.n4202 GND.n2698 240.244
R4220 GND.n4202 GND.n2708 240.244
R4221 GND.n2713 GND.n2708 240.244
R4222 GND.n4211 GND.n2713 240.244
R4223 GND.n4212 GND.n4211 240.244
R4224 GND.n4212 GND.n2725 240.244
R4225 GND.n2725 GND.n321 240.244
R4226 GND.n2733 GND.n321 240.244
R4227 GND.n2755 GND.n2733 240.244
R4228 GND.n4221 GND.n2755 240.244
R4229 GND.n4221 GND.n340 240.244
R4230 GND.n4232 GND.n340 240.244
R4231 GND.n4232 GND.n352 240.244
R4232 GND.n2740 GND.n352 240.244
R4233 GND.n2740 GND.n361 240.244
R4234 GND.n4262 GND.n361 240.244
R4235 GND.n4262 GND.n371 240.244
R4236 GND.n4258 GND.n371 240.244
R4237 GND.n4258 GND.n382 240.244
R4238 GND.n4250 GND.n382 240.244
R4239 GND.n4250 GND.n392 240.244
R4240 GND.n5670 GND.n392 240.244
R4241 GND.n5670 GND.n402 240.244
R4242 GND.n5698 GND.n402 240.244
R4243 GND.n5698 GND.n412 240.244
R4244 GND.n5694 GND.n412 240.244
R4245 GND.n5694 GND.n423 240.244
R4246 GND.n5689 GND.n423 240.244
R4247 GND.n5689 GND.n432 240.244
R4248 GND.n5686 GND.n432 240.244
R4249 GND.n5686 GND.n442 240.244
R4250 GND.n5683 GND.n442 240.244
R4251 GND.n5683 GND.n451 240.244
R4252 GND.n5680 GND.n451 240.244
R4253 GND.n5680 GND.n461 240.244
R4254 GND.n5677 GND.n461 240.244
R4255 GND.n5677 GND.n469 240.244
R4256 GND.n2518 GND.n2517 240.244
R4257 GND.n4476 GND.n2517 240.244
R4258 GND.n4474 GND.n4473 240.244
R4259 GND.n4470 GND.n4469 240.244
R4260 GND.n4466 GND.n4465 240.244
R4261 GND.n4462 GND.n4461 240.244
R4262 GND.n4458 GND.n4457 240.244
R4263 GND.n4454 GND.n4453 240.244
R4264 GND.n4449 GND.n4448 240.244
R4265 GND.n4445 GND.n4444 240.244
R4266 GND.n4441 GND.n4440 240.244
R4267 GND.n4437 GND.n4436 240.244
R4268 GND.n4433 GND.n4432 240.244
R4269 GND.n4429 GND.n4428 240.244
R4270 GND.n4425 GND.n4424 240.244
R4271 GND.n4421 GND.n4420 240.244
R4272 GND.n4417 GND.n4416 240.244
R4273 GND.n2560 GND.n2559 240.244
R4274 GND.n2579 GND.n2519 240.244
R4275 GND.n4398 GND.n2579 240.244
R4276 GND.n4398 GND.n2580 240.244
R4277 GND.n4394 GND.n2580 240.244
R4278 GND.n4394 GND.n2589 240.244
R4279 GND.n4386 GND.n2589 240.244
R4280 GND.n4386 GND.n2607 240.244
R4281 GND.n4382 GND.n2607 240.244
R4282 GND.n4382 GND.n2613 240.244
R4283 GND.n4374 GND.n2613 240.244
R4284 GND.n4374 GND.n2628 240.244
R4285 GND.n4370 GND.n2628 240.244
R4286 GND.n4370 GND.n2634 240.244
R4287 GND.n4362 GND.n2634 240.244
R4288 GND.n4362 GND.n2648 240.244
R4289 GND.n4358 GND.n2648 240.244
R4290 GND.n4358 GND.n2654 240.244
R4291 GND.n4350 GND.n2654 240.244
R4292 GND.n4350 GND.n2669 240.244
R4293 GND.n4346 GND.n2669 240.244
R4294 GND.n4346 GND.n2675 240.244
R4295 GND.n4338 GND.n2675 240.244
R4296 GND.n4338 GND.n2690 240.244
R4297 GND.n4334 GND.n2690 240.244
R4298 GND.n4334 GND.n2696 240.244
R4299 GND.n4326 GND.n2696 240.244
R4300 GND.n4326 GND.n4324 240.244
R4301 GND.n4324 GND.n2711 240.244
R4302 GND.n2723 GND.n2711 240.244
R4303 GND.n2723 GND.n324 240.244
R4304 GND.n5917 GND.n324 240.244
R4305 GND.n5917 GND.n325 240.244
R4306 GND.n2753 GND.n325 240.244
R4307 GND.n2753 GND.n337 240.244
R4308 GND.n5912 GND.n337 240.244
R4309 GND.n5912 GND.n338 240.244
R4310 GND.n5904 GND.n338 240.244
R4311 GND.n5904 GND.n354 240.244
R4312 GND.n5900 GND.n354 240.244
R4313 GND.n5900 GND.n359 240.244
R4314 GND.n5892 GND.n359 240.244
R4315 GND.n5892 GND.n374 240.244
R4316 GND.n5888 GND.n374 240.244
R4317 GND.n5888 GND.n380 240.244
R4318 GND.n5880 GND.n380 240.244
R4319 GND.n5880 GND.n395 240.244
R4320 GND.n5876 GND.n395 240.244
R4321 GND.n5876 GND.n401 240.244
R4322 GND.n5868 GND.n401 240.244
R4323 GND.n5868 GND.n415 240.244
R4324 GND.n5864 GND.n415 240.244
R4325 GND.n5864 GND.n421 240.244
R4326 GND.n5856 GND.n421 240.244
R4327 GND.n5856 GND.n435 240.244
R4328 GND.n5852 GND.n435 240.244
R4329 GND.n5852 GND.n441 240.244
R4330 GND.n5844 GND.n441 240.244
R4331 GND.n5844 GND.n454 240.244
R4332 GND.n5840 GND.n454 240.244
R4333 GND.n5840 GND.n460 240.244
R4334 GND.n5832 GND.n460 240.244
R4335 GND.n1245 GND.n1241 240.244
R4336 GND.n4734 GND.n1246 240.244
R4337 GND.n1250 GND.n1249 240.244
R4338 GND.n4731 GND.n1251 240.244
R4339 GND.n1255 GND.n1254 240.244
R4340 GND.n4728 GND.n1256 240.244
R4341 GND.n1260 GND.n1259 240.244
R4342 GND.n4725 GND.n1261 240.244
R4343 GND.n1269 GND.n1268 240.244
R4344 GND.n4722 GND.n1272 240.244
R4345 GND.n1274 GND.n1273 240.244
R4346 GND.n4719 GND.n1277 240.244
R4347 GND.n1279 GND.n1278 240.244
R4348 GND.n4716 GND.n1282 240.244
R4349 GND.n1284 GND.n1283 240.244
R4350 GND.n4713 GND.n1287 240.244
R4351 GND.n1289 GND.n1288 240.244
R4352 GND.n4739 GND.n1294 240.244
R4353 GND.n1697 GND.n1689 240.244
R4354 GND.n1941 GND.n1689 240.244
R4355 GND.n1941 GND.n1678 240.244
R4356 GND.n1678 GND.n1669 240.244
R4357 GND.n1957 GND.n1669 240.244
R4358 GND.n1958 GND.n1957 240.244
R4359 GND.n1958 GND.n1660 240.244
R4360 GND.n1960 GND.n1660 240.244
R4361 GND.n1960 GND.n1652 240.244
R4362 GND.n1961 GND.n1652 240.244
R4363 GND.n1961 GND.n1116 240.244
R4364 GND.n1645 GND.n1116 240.244
R4365 GND.n1645 GND.n1129 240.244
R4366 GND.n1139 GND.n1129 240.244
R4367 GND.n1140 GND.n1139 240.244
R4368 GND.n1639 GND.n1140 240.244
R4369 GND.n1639 GND.n1146 240.244
R4370 GND.n1147 GND.n1146 240.244
R4371 GND.n1148 GND.n1147 240.244
R4372 GND.n1598 GND.n1148 240.244
R4373 GND.n1598 GND.n1154 240.244
R4374 GND.n1155 GND.n1154 240.244
R4375 GND.n1156 GND.n1155 240.244
R4376 GND.n1580 GND.n1156 240.244
R4377 GND.n1580 GND.n1162 240.244
R4378 GND.n1163 GND.n1162 240.244
R4379 GND.n1164 GND.n1163 240.244
R4380 GND.n1529 GND.n1164 240.244
R4381 GND.n1529 GND.n1170 240.244
R4382 GND.n1171 GND.n1170 240.244
R4383 GND.n1172 GND.n1171 240.244
R4384 GND.n1566 GND.n1172 240.244
R4385 GND.n1566 GND.n1178 240.244
R4386 GND.n1179 GND.n1178 240.244
R4387 GND.n1180 GND.n1179 240.244
R4388 GND.n1560 GND.n1180 240.244
R4389 GND.n1560 GND.n1186 240.244
R4390 GND.n1187 GND.n1186 240.244
R4391 GND.n1188 GND.n1187 240.244
R4392 GND.n1489 GND.n1188 240.244
R4393 GND.n1489 GND.n1194 240.244
R4394 GND.n1195 GND.n1194 240.244
R4395 GND.n1196 GND.n1195 240.244
R4396 GND.n2223 GND.n1196 240.244
R4397 GND.n2223 GND.n1202 240.244
R4398 GND.n1203 GND.n1202 240.244
R4399 GND.n1204 GND.n1203 240.244
R4400 GND.n1456 GND.n1204 240.244
R4401 GND.n1456 GND.n1210 240.244
R4402 GND.n1211 GND.n1210 240.244
R4403 GND.n1212 GND.n1211 240.244
R4404 GND.n1438 GND.n1212 240.244
R4405 GND.n1438 GND.n1218 240.244
R4406 GND.n1219 GND.n1218 240.244
R4407 GND.n1220 GND.n1219 240.244
R4408 GND.n1415 GND.n1220 240.244
R4409 GND.n1415 GND.n1226 240.244
R4410 GND.n1227 GND.n1226 240.244
R4411 GND.n1228 GND.n1227 240.244
R4412 GND.n1234 GND.n1228 240.244
R4413 GND.n4801 GND.n1234 240.244
R4414 GND.n1910 GND.n1908 240.244
R4415 GND.n1908 GND.n1907 240.244
R4416 GND.n1904 GND.n1903 240.244
R4417 GND.n1901 GND.n1708 240.244
R4418 GND.n1897 GND.n1895 240.244
R4419 GND.n1893 GND.n1714 240.244
R4420 GND.n1889 GND.n1887 240.244
R4421 GND.n1885 GND.n1720 240.244
R4422 GND.n1881 GND.n1879 240.244
R4423 GND.n1877 GND.n1726 240.244
R4424 GND.n1873 GND.n1871 240.244
R4425 GND.n1869 GND.n1735 240.244
R4426 GND.n1865 GND.n1863 240.244
R4427 GND.n1861 GND.n1741 240.244
R4428 GND.n1857 GND.n1855 240.244
R4429 GND.n1853 GND.n1747 240.244
R4430 GND.n1849 GND.n1847 240.244
R4431 GND.n1845 GND.n1753 240.244
R4432 GND.n1835 GND.n1758 240.244
R4433 GND.n1918 GND.n1700 240.244
R4434 GND.n1700 GND.n1677 240.244
R4435 GND.n1949 GND.n1677 240.244
R4436 GND.n1949 GND.n1673 240.244
R4437 GND.n1955 GND.n1673 240.244
R4438 GND.n1955 GND.n1658 240.244
R4439 GND.n1978 GND.n1658 240.244
R4440 GND.n1978 GND.n1654 240.244
R4441 GND.n1985 GND.n1654 240.244
R4442 GND.n1985 GND.n1120 240.244
R4443 GND.n4883 GND.n1120 240.244
R4444 GND.n4883 GND.n1121 240.244
R4445 GND.n4879 GND.n1121 240.244
R4446 GND.n4879 GND.n1127 240.244
R4447 GND.n1637 GND.n1127 240.244
R4448 GND.n1637 GND.n1614 240.244
R4449 GND.n2022 GND.n1614 240.244
R4450 GND.n2022 GND.n1609 240.244
R4451 GND.n2030 GND.n1609 240.244
R4452 GND.n2030 GND.n1610 240.244
R4453 GND.n1610 GND.n1588 240.244
R4454 GND.n2059 GND.n1588 240.244
R4455 GND.n2059 GND.n1584 240.244
R4456 GND.n2066 GND.n1584 240.244
R4457 GND.n2066 GND.n1523 240.244
R4458 GND.n2133 GND.n1523 240.244
R4459 GND.n2133 GND.n1524 240.244
R4460 GND.n2128 GND.n1524 240.244
R4461 GND.n2128 GND.n1527 240.244
R4462 GND.n1545 GND.n1527 240.244
R4463 GND.n2116 GND.n1545 240.244
R4464 GND.n2116 GND.n1546 240.244
R4465 GND.n2111 GND.n1546 240.244
R4466 GND.n2111 GND.n1550 240.244
R4467 GND.n2094 GND.n1550 240.244
R4468 GND.n2099 GND.n2094 240.244
R4469 GND.n2099 GND.n1498 240.244
R4470 GND.n2203 GND.n1498 240.244
R4471 GND.n2203 GND.n1492 240.244
R4472 GND.n2211 GND.n1492 240.244
R4473 GND.n2211 GND.n1494 240.244
R4474 GND.n1494 GND.n1475 240.244
R4475 GND.n2228 GND.n1475 240.244
R4476 GND.n2228 GND.n1470 240.244
R4477 GND.n2236 GND.n1470 240.244
R4478 GND.n2236 GND.n1471 240.244
R4479 GND.n1471 GND.n1454 240.244
R4480 GND.n2252 GND.n1454 240.244
R4481 GND.n2252 GND.n1449 240.244
R4482 GND.n2260 GND.n1449 240.244
R4483 GND.n2260 GND.n1450 240.244
R4484 GND.n1450 GND.n1433 240.244
R4485 GND.n2279 GND.n1433 240.244
R4486 GND.n2279 GND.n1429 240.244
R4487 GND.n2285 GND.n1429 240.244
R4488 GND.n2285 GND.n1409 240.244
R4489 GND.n2319 GND.n1409 240.244
R4490 GND.n2319 GND.n1405 240.244
R4491 GND.n2325 GND.n1405 240.244
R4492 GND.n2325 GND.n1240 240.244
R4493 GND.n4799 GND.n1240 240.244
R4494 GND.n544 GND.n468 240.244
R4495 GND.n5753 GND.n5752 240.244
R4496 GND.n5750 GND.n548 240.244
R4497 GND.n5746 GND.n5745 240.244
R4498 GND.n5743 GND.n555 240.244
R4499 GND.n5739 GND.n5738 240.244
R4500 GND.n5736 GND.n562 240.244
R4501 GND.n5732 GND.n5731 240.244
R4502 GND.n5729 GND.n569 240.244
R4503 GND.n3989 GND.n2567 240.244
R4504 GND.n3989 GND.n2577 240.244
R4505 GND.n4109 GND.n2577 240.244
R4506 GND.n4109 GND.n2592 240.244
R4507 GND.n4115 GND.n2592 240.244
R4508 GND.n4115 GND.n2605 240.244
R4509 GND.n4124 GND.n2605 240.244
R4510 GND.n4124 GND.n2616 240.244
R4511 GND.n4130 GND.n2616 240.244
R4512 GND.n4130 GND.n2626 240.244
R4513 GND.n4139 GND.n2626 240.244
R4514 GND.n4139 GND.n2637 240.244
R4515 GND.n4145 GND.n2637 240.244
R4516 GND.n4145 GND.n2647 240.244
R4517 GND.n4154 GND.n2647 240.244
R4518 GND.n4154 GND.n2657 240.244
R4519 GND.n4160 GND.n2657 240.244
R4520 GND.n4160 GND.n2667 240.244
R4521 GND.n4169 GND.n2667 240.244
R4522 GND.n4169 GND.n2678 240.244
R4523 GND.n4175 GND.n2678 240.244
R4524 GND.n4175 GND.n2688 240.244
R4525 GND.n4184 GND.n2688 240.244
R4526 GND.n4184 GND.n2699 240.244
R4527 GND.n4200 GND.n2699 240.244
R4528 GND.n4200 GND.n2709 240.244
R4529 GND.n2714 GND.n2709 240.244
R4530 GND.n4195 GND.n2714 240.244
R4531 GND.n4195 GND.n4194 240.244
R4532 GND.n4194 GND.n318 240.244
R4533 GND.n5919 GND.n318 240.244
R4534 GND.n5919 GND.n319 240.244
R4535 GND.n2750 GND.n319 240.244
R4536 GND.n4223 GND.n2750 240.244
R4537 GND.n4223 GND.n341 240.244
R4538 GND.n4230 GND.n341 240.244
R4539 GND.n4230 GND.n353 240.244
R4540 GND.n4268 GND.n353 240.244
R4541 GND.n4268 GND.n362 240.244
R4542 GND.n4264 GND.n362 240.244
R4543 GND.n4264 GND.n372 240.244
R4544 GND.n4256 GND.n372 240.244
R4545 GND.n4256 GND.n383 240.244
R4546 GND.n4252 GND.n383 240.244
R4547 GND.n4252 GND.n393 240.244
R4548 GND.n589 GND.n393 240.244
R4549 GND.n589 GND.n403 240.244
R4550 GND.n5700 GND.n403 240.244
R4551 GND.n5700 GND.n413 240.244
R4552 GND.n5692 GND.n413 240.244
R4553 GND.n5692 GND.n424 240.244
R4554 GND.n5707 GND.n424 240.244
R4555 GND.n5707 GND.n433 240.244
R4556 GND.n581 GND.n433 240.244
R4557 GND.n581 GND.n443 240.244
R4558 GND.n5714 GND.n443 240.244
R4559 GND.n5714 GND.n452 240.244
R4560 GND.n578 GND.n452 240.244
R4561 GND.n578 GND.n462 240.244
R4562 GND.n5721 GND.n462 240.244
R4563 GND.n5721 GND.n470 240.244
R4564 GND.n2441 GND.n2440 240.244
R4565 GND.n2504 GND.n2448 240.244
R4566 GND.n2507 GND.n2449 240.244
R4567 GND.n2457 GND.n2456 240.244
R4568 GND.n2509 GND.n2464 240.244
R4569 GND.n2512 GND.n2465 240.244
R4570 GND.n2473 GND.n2472 240.244
R4571 GND.n2514 GND.n2480 240.244
R4572 GND.n4485 GND.n2483 240.244
R4573 GND.n4406 GND.n2570 240.244
R4574 GND.n2578 GND.n2570 240.244
R4575 GND.n2594 GND.n2578 240.244
R4576 GND.n4392 GND.n2594 240.244
R4577 GND.n4392 GND.n2595 240.244
R4578 GND.n4388 GND.n2595 240.244
R4579 GND.n4388 GND.n2602 240.244
R4580 GND.n4380 GND.n2602 240.244
R4581 GND.n4380 GND.n2618 240.244
R4582 GND.n4376 GND.n2618 240.244
R4583 GND.n4376 GND.n2623 240.244
R4584 GND.n4368 GND.n2623 240.244
R4585 GND.n4368 GND.n2639 240.244
R4586 GND.n4364 GND.n2639 240.244
R4587 GND.n4364 GND.n2644 240.244
R4588 GND.n4356 GND.n2644 240.244
R4589 GND.n4356 GND.n2659 240.244
R4590 GND.n4352 GND.n2659 240.244
R4591 GND.n4352 GND.n2664 240.244
R4592 GND.n4344 GND.n2664 240.244
R4593 GND.n4344 GND.n2680 240.244
R4594 GND.n4340 GND.n2680 240.244
R4595 GND.n4340 GND.n2685 240.244
R4596 GND.n4332 GND.n2685 240.244
R4597 GND.n4332 GND.n2701 240.244
R4598 GND.n4328 GND.n2701 240.244
R4599 GND.n4328 GND.n2706 240.244
R4600 GND.n4207 GND.n2706 240.244
R4601 GND.n4207 GND.n2726 240.244
R4602 GND.n4313 GND.n2726 240.244
R4603 GND.n4313 GND.n323 240.244
R4604 GND.n4309 GND.n323 240.244
R4605 GND.n4309 GND.n2732 240.244
R4606 GND.n2732 GND.n343 240.244
R4607 GND.n5910 GND.n343 240.244
R4608 GND.n5910 GND.n344 240.244
R4609 GND.n5906 GND.n344 240.244
R4610 GND.n5906 GND.n350 240.244
R4611 GND.n5898 GND.n350 240.244
R4612 GND.n5898 GND.n364 240.244
R4613 GND.n5894 GND.n364 240.244
R4614 GND.n5894 GND.n369 240.244
R4615 GND.n5886 GND.n369 240.244
R4616 GND.n5886 GND.n385 240.244
R4617 GND.n5882 GND.n385 240.244
R4618 GND.n5882 GND.n390 240.244
R4619 GND.n5874 GND.n390 240.244
R4620 GND.n5874 GND.n405 240.244
R4621 GND.n5870 GND.n405 240.244
R4622 GND.n5870 GND.n410 240.244
R4623 GND.n5862 GND.n410 240.244
R4624 GND.n5862 GND.n425 240.244
R4625 GND.n5858 GND.n425 240.244
R4626 GND.n5858 GND.n430 240.244
R4627 GND.n5850 GND.n430 240.244
R4628 GND.n5850 GND.n445 240.244
R4629 GND.n5846 GND.n445 240.244
R4630 GND.n5846 GND.n450 240.244
R4631 GND.n5838 GND.n450 240.244
R4632 GND.n5838 GND.n464 240.244
R4633 GND.n5834 GND.n464 240.244
R4634 GND.n1336 GND.n1296 240.244
R4635 GND.n1338 GND.n1337 240.244
R4636 GND.n1347 GND.n1346 240.244
R4637 GND.n1355 GND.n1354 240.244
R4638 GND.n1357 GND.n1356 240.244
R4639 GND.n1367 GND.n1366 240.244
R4640 GND.n1375 GND.n1374 240.244
R4641 GND.n1377 GND.n1376 240.244
R4642 GND.n1390 GND.n1386 240.244
R4643 GND.n1920 GND.n1691 240.244
R4644 GND.n1939 GND.n1691 240.244
R4645 GND.n1939 GND.n1679 240.244
R4646 GND.n1925 GND.n1679 240.244
R4647 GND.n1925 GND.n1671 240.244
R4648 GND.n1926 GND.n1671 240.244
R4649 GND.n1926 GND.n1661 240.244
R4650 GND.n1661 GND.n1650 240.244
R4651 GND.n1987 GND.n1650 240.244
R4652 GND.n1988 GND.n1987 240.244
R4653 GND.n1988 GND.n1117 240.244
R4654 GND.n1647 GND.n1117 240.244
R4655 GND.n1647 GND.n1130 240.244
R4656 GND.n1997 GND.n1130 240.244
R4657 GND.n1997 GND.n1640 240.244
R4658 GND.n2004 GND.n1640 240.244
R4659 GND.n2004 GND.n1616 240.244
R4660 GND.n1616 GND.n1605 240.244
R4661 GND.n2032 GND.n1605 240.244
R4662 GND.n2032 GND.n1600 240.244
R4663 GND.n2042 GND.n1600 240.244
R4664 GND.n2042 GND.n1590 240.244
R4665 GND.n1590 GND.n1579 240.244
R4666 GND.n2068 GND.n1579 240.244
R4667 GND.n2069 GND.n2068 240.244
R4668 GND.n2069 GND.n1519 240.244
R4669 GND.n1575 GND.n1519 240.244
R4670 GND.n1575 GND.n1530 240.244
R4671 GND.n1535 GND.n1530 240.244
R4672 GND.n2077 GND.n1535 240.244
R4673 GND.n2077 GND.n1542 240.244
R4674 GND.n1572 GND.n1542 240.244
R4675 GND.n1572 GND.n1551 240.244
R4676 GND.n1556 GND.n1551 240.244
R4677 GND.n1561 GND.n1556 240.244
R4678 GND.n2093 GND.n1561 240.244
R4679 GND.n2093 GND.n1503 240.244
R4680 GND.n1503 GND.n1499 240.244
R4681 GND.n1499 GND.n1487 240.244
R4682 GND.n2213 GND.n1487 240.244
R4683 GND.n2213 GND.n1482 240.244
R4684 GND.n2220 GND.n1482 240.244
R4685 GND.n2220 GND.n1477 240.244
R4686 GND.n1477 GND.n1466 240.244
R4687 GND.n2238 GND.n1466 240.244
R4688 GND.n2238 GND.n1461 240.244
R4689 GND.n2245 GND.n1461 240.244
R4690 GND.n2245 GND.n1457 240.244
R4691 GND.n1457 GND.n1444 240.244
R4692 GND.n2262 GND.n1444 240.244
R4693 GND.n2262 GND.n1439 240.244
R4694 GND.n2272 GND.n1439 240.244
R4695 GND.n2272 GND.n1435 240.244
R4696 GND.n2266 GND.n1435 240.244
R4697 GND.n2266 GND.n1416 240.244
R4698 GND.n2314 GND.n1416 240.244
R4699 GND.n2314 GND.n1411 240.244
R4700 GND.n2308 GND.n1411 240.244
R4701 GND.n2308 GND.n1401 240.244
R4702 GND.n2330 GND.n1401 240.244
R4703 GND.n2330 GND.n1237 240.244
R4704 GND.n1829 GND.n1828 240.244
R4705 GND.n1774 GND.n1773 240.244
R4706 GND.n1777 GND.n1776 240.244
R4707 GND.n1782 GND.n1781 240.244
R4708 GND.n1785 GND.n1784 240.244
R4709 GND.n1790 GND.n1789 240.244
R4710 GND.n1793 GND.n1792 240.244
R4711 GND.n1798 GND.n1797 240.244
R4712 GND.n1801 GND.n1695 240.244
R4713 GND.n1763 GND.n1698 240.244
R4714 GND.n1763 GND.n1680 240.244
R4715 GND.n1947 GND.n1680 240.244
R4716 GND.n1947 GND.n1681 240.244
R4717 GND.n1681 GND.n1672 240.244
R4718 GND.n1672 GND.n1662 240.244
R4719 GND.n1976 GND.n1662 240.244
R4720 GND.n1976 GND.n1663 240.244
R4721 GND.n1663 GND.n1653 240.244
R4722 GND.n1964 GND.n1653 240.244
R4723 GND.n1964 GND.n1119 240.244
R4724 GND.n1132 GND.n1119 240.244
R4725 GND.n4877 GND.n1132 240.244
R4726 GND.n4877 GND.n1133 240.244
R4727 GND.n1633 GND.n1133 240.244
R4728 GND.n1633 GND.n1618 240.244
R4729 GND.n2020 GND.n1618 240.244
R4730 GND.n2020 GND.n2019 240.244
R4731 GND.n2019 GND.n1608 240.244
R4732 GND.n1608 GND.n1607 240.244
R4733 GND.n1607 GND.n1592 240.244
R4734 GND.n2057 GND.n1592 240.244
R4735 GND.n2057 GND.n2055 240.244
R4736 GND.n2055 GND.n1583 240.244
R4737 GND.n1583 GND.n1582 240.244
R4738 GND.n1582 GND.n1522 240.244
R4739 GND.n1531 GND.n1522 240.244
R4740 GND.n2126 GND.n1531 240.244
R4741 GND.n2126 GND.n2125 240.244
R4742 GND.n2125 GND.n1533 240.244
R4743 GND.n1544 GND.n1533 240.244
R4744 GND.n1553 GND.n1544 240.244
R4745 GND.n2109 GND.n1553 240.244
R4746 GND.n2109 GND.n2108 240.244
R4747 GND.n2108 GND.n1554 240.244
R4748 GND.n1554 GND.n1501 240.244
R4749 GND.n2197 GND.n1501 240.244
R4750 GND.n2201 GND.n2197 240.244
R4751 GND.n2201 GND.n2199 240.244
R4752 GND.n2199 GND.n1491 240.244
R4753 GND.n1491 GND.n1479 240.244
R4754 GND.n2222 GND.n1479 240.244
R4755 GND.n2226 GND.n2222 240.244
R4756 GND.n2226 GND.n2225 240.244
R4757 GND.n2225 GND.n1469 240.244
R4758 GND.n1469 GND.n1460 240.244
R4759 GND.n2247 GND.n1460 240.244
R4760 GND.n2250 GND.n2247 240.244
R4761 GND.n2250 GND.n2249 240.244
R4762 GND.n2249 GND.n1448 240.244
R4763 GND.n1448 GND.n1437 240.244
R4764 GND.n2274 GND.n1437 240.244
R4765 GND.n2277 GND.n2274 240.244
R4766 GND.n2277 GND.n2276 240.244
R4767 GND.n2276 GND.n1413 240.244
R4768 GND.n2316 GND.n1413 240.244
R4769 GND.n2317 GND.n2316 240.244
R4770 GND.n2317 GND.n1404 240.244
R4771 GND.n2327 GND.n1404 240.244
R4772 GND.n2328 GND.n2327 240.244
R4773 GND.n2328 GND.n1239 240.244
R4774 GND.n5032 GND.n972 240.244
R4775 GND.n5032 GND.n968 240.244
R4776 GND.n5038 GND.n968 240.244
R4777 GND.n5038 GND.n966 240.244
R4778 GND.n5042 GND.n966 240.244
R4779 GND.n5042 GND.n962 240.244
R4780 GND.n5048 GND.n962 240.244
R4781 GND.n5048 GND.n960 240.244
R4782 GND.n5052 GND.n960 240.244
R4783 GND.n5052 GND.n956 240.244
R4784 GND.n5058 GND.n956 240.244
R4785 GND.n5058 GND.n954 240.244
R4786 GND.n5062 GND.n954 240.244
R4787 GND.n5062 GND.n950 240.244
R4788 GND.n5068 GND.n950 240.244
R4789 GND.n5068 GND.n948 240.244
R4790 GND.n5072 GND.n948 240.244
R4791 GND.n5072 GND.n944 240.244
R4792 GND.n5078 GND.n944 240.244
R4793 GND.n5078 GND.n942 240.244
R4794 GND.n5082 GND.n942 240.244
R4795 GND.n5082 GND.n938 240.244
R4796 GND.n5088 GND.n938 240.244
R4797 GND.n5088 GND.n936 240.244
R4798 GND.n5092 GND.n936 240.244
R4799 GND.n5092 GND.n932 240.244
R4800 GND.n5098 GND.n932 240.244
R4801 GND.n5098 GND.n930 240.244
R4802 GND.n5102 GND.n930 240.244
R4803 GND.n5102 GND.n926 240.244
R4804 GND.n5108 GND.n926 240.244
R4805 GND.n5108 GND.n924 240.244
R4806 GND.n5112 GND.n924 240.244
R4807 GND.n5112 GND.n920 240.244
R4808 GND.n5118 GND.n920 240.244
R4809 GND.n5118 GND.n918 240.244
R4810 GND.n5122 GND.n918 240.244
R4811 GND.n5122 GND.n914 240.244
R4812 GND.n5128 GND.n914 240.244
R4813 GND.n5128 GND.n912 240.244
R4814 GND.n5132 GND.n912 240.244
R4815 GND.n5132 GND.n908 240.244
R4816 GND.n5138 GND.n908 240.244
R4817 GND.n5138 GND.n906 240.244
R4818 GND.n5142 GND.n906 240.244
R4819 GND.n5142 GND.n902 240.244
R4820 GND.n5148 GND.n902 240.244
R4821 GND.n5148 GND.n900 240.244
R4822 GND.n5152 GND.n900 240.244
R4823 GND.n5152 GND.n896 240.244
R4824 GND.n5158 GND.n896 240.244
R4825 GND.n5158 GND.n894 240.244
R4826 GND.n5162 GND.n894 240.244
R4827 GND.n5162 GND.n890 240.244
R4828 GND.n5168 GND.n890 240.244
R4829 GND.n5168 GND.n888 240.244
R4830 GND.n5172 GND.n888 240.244
R4831 GND.n5172 GND.n884 240.244
R4832 GND.n5178 GND.n884 240.244
R4833 GND.n5178 GND.n882 240.244
R4834 GND.n5182 GND.n882 240.244
R4835 GND.n5182 GND.n878 240.244
R4836 GND.n5188 GND.n878 240.244
R4837 GND.n5188 GND.n876 240.244
R4838 GND.n5192 GND.n876 240.244
R4839 GND.n5192 GND.n872 240.244
R4840 GND.n5198 GND.n872 240.244
R4841 GND.n5198 GND.n870 240.244
R4842 GND.n5202 GND.n870 240.244
R4843 GND.n5202 GND.n866 240.244
R4844 GND.n5208 GND.n866 240.244
R4845 GND.n5208 GND.n864 240.244
R4846 GND.n5212 GND.n864 240.244
R4847 GND.n5212 GND.n860 240.244
R4848 GND.n5218 GND.n860 240.244
R4849 GND.n5218 GND.n858 240.244
R4850 GND.n5222 GND.n858 240.244
R4851 GND.n5222 GND.n854 240.244
R4852 GND.n5228 GND.n854 240.244
R4853 GND.n5228 GND.n852 240.244
R4854 GND.n5232 GND.n852 240.244
R4855 GND.n5232 GND.n848 240.244
R4856 GND.n5238 GND.n848 240.244
R4857 GND.n5238 GND.n846 240.244
R4858 GND.n5242 GND.n846 240.244
R4859 GND.n5242 GND.n842 240.244
R4860 GND.n5248 GND.n842 240.244
R4861 GND.n5248 GND.n840 240.244
R4862 GND.n5252 GND.n840 240.244
R4863 GND.n5252 GND.n836 240.244
R4864 GND.n5258 GND.n836 240.244
R4865 GND.n5258 GND.n834 240.244
R4866 GND.n5262 GND.n834 240.244
R4867 GND.n5262 GND.n830 240.244
R4868 GND.n5268 GND.n830 240.244
R4869 GND.n5268 GND.n828 240.244
R4870 GND.n5272 GND.n828 240.244
R4871 GND.n5272 GND.n824 240.244
R4872 GND.n5278 GND.n824 240.244
R4873 GND.n5278 GND.n822 240.244
R4874 GND.n5282 GND.n822 240.244
R4875 GND.n5282 GND.n818 240.244
R4876 GND.n5288 GND.n818 240.244
R4877 GND.n5288 GND.n816 240.244
R4878 GND.n5292 GND.n816 240.244
R4879 GND.n5292 GND.n812 240.244
R4880 GND.n5298 GND.n812 240.244
R4881 GND.n5298 GND.n810 240.244
R4882 GND.n5302 GND.n810 240.244
R4883 GND.n5302 GND.n806 240.244
R4884 GND.n5308 GND.n806 240.244
R4885 GND.n5308 GND.n804 240.244
R4886 GND.n5312 GND.n804 240.244
R4887 GND.n5312 GND.n800 240.244
R4888 GND.n5318 GND.n800 240.244
R4889 GND.n5318 GND.n798 240.244
R4890 GND.n5322 GND.n798 240.244
R4891 GND.n5322 GND.n794 240.244
R4892 GND.n5328 GND.n794 240.244
R4893 GND.n5328 GND.n792 240.244
R4894 GND.n5332 GND.n792 240.244
R4895 GND.n5332 GND.n788 240.244
R4896 GND.n5338 GND.n788 240.244
R4897 GND.n5338 GND.n786 240.244
R4898 GND.n5342 GND.n786 240.244
R4899 GND.n5342 GND.n782 240.244
R4900 GND.n5348 GND.n782 240.244
R4901 GND.n5348 GND.n780 240.244
R4902 GND.n5352 GND.n780 240.244
R4903 GND.n5352 GND.n776 240.244
R4904 GND.n5358 GND.n776 240.244
R4905 GND.n5358 GND.n774 240.244
R4906 GND.n5362 GND.n774 240.244
R4907 GND.n5362 GND.n770 240.244
R4908 GND.n5368 GND.n770 240.244
R4909 GND.n5368 GND.n768 240.244
R4910 GND.n5372 GND.n768 240.244
R4911 GND.n5372 GND.n764 240.244
R4912 GND.n5378 GND.n764 240.244
R4913 GND.n5378 GND.n762 240.244
R4914 GND.n5382 GND.n762 240.244
R4915 GND.n5382 GND.n758 240.244
R4916 GND.n5388 GND.n758 240.244
R4917 GND.n5388 GND.n756 240.244
R4918 GND.n5392 GND.n756 240.244
R4919 GND.n5392 GND.n752 240.244
R4920 GND.n5398 GND.n752 240.244
R4921 GND.n5398 GND.n750 240.244
R4922 GND.n5402 GND.n750 240.244
R4923 GND.n5402 GND.n746 240.244
R4924 GND.n5408 GND.n746 240.244
R4925 GND.n5408 GND.n744 240.244
R4926 GND.n5412 GND.n744 240.244
R4927 GND.n5412 GND.n740 240.244
R4928 GND.n5418 GND.n740 240.244
R4929 GND.n5418 GND.n738 240.244
R4930 GND.n5422 GND.n738 240.244
R4931 GND.n5422 GND.n734 240.244
R4932 GND.n5428 GND.n734 240.244
R4933 GND.n5428 GND.n732 240.244
R4934 GND.n5432 GND.n732 240.244
R4935 GND.n5432 GND.n728 240.244
R4936 GND.n5438 GND.n728 240.244
R4937 GND.n5438 GND.n726 240.244
R4938 GND.n5442 GND.n726 240.244
R4939 GND.n5442 GND.n722 240.244
R4940 GND.n5448 GND.n722 240.244
R4941 GND.n5448 GND.n720 240.244
R4942 GND.n5452 GND.n720 240.244
R4943 GND.n5452 GND.n716 240.244
R4944 GND.n5458 GND.n716 240.244
R4945 GND.n5458 GND.n714 240.244
R4946 GND.n5462 GND.n714 240.244
R4947 GND.n5462 GND.n710 240.244
R4948 GND.n5468 GND.n710 240.244
R4949 GND.n5468 GND.n708 240.244
R4950 GND.n5472 GND.n708 240.244
R4951 GND.n5472 GND.n704 240.244
R4952 GND.n5479 GND.n704 240.244
R4953 GND.n5479 GND.n702 240.244
R4954 GND.n5483 GND.n699 240.244
R4955 GND.n5489 GND.n699 240.244
R4956 GND.n5489 GND.n697 240.244
R4957 GND.n5493 GND.n697 240.244
R4958 GND.n5493 GND.n693 240.244
R4959 GND.n5499 GND.n693 240.244
R4960 GND.n5499 GND.n691 240.244
R4961 GND.n5503 GND.n691 240.244
R4962 GND.n5503 GND.n687 240.244
R4963 GND.n5509 GND.n687 240.244
R4964 GND.n5509 GND.n685 240.244
R4965 GND.n5513 GND.n685 240.244
R4966 GND.n5513 GND.n681 240.244
R4967 GND.n5519 GND.n681 240.244
R4968 GND.n5519 GND.n679 240.244
R4969 GND.n5523 GND.n679 240.244
R4970 GND.n5523 GND.n675 240.244
R4971 GND.n5529 GND.n675 240.244
R4972 GND.n5529 GND.n673 240.244
R4973 GND.n5533 GND.n673 240.244
R4974 GND.n5533 GND.n669 240.244
R4975 GND.n5539 GND.n669 240.244
R4976 GND.n5539 GND.n667 240.244
R4977 GND.n5543 GND.n667 240.244
R4978 GND.n5543 GND.n663 240.244
R4979 GND.n5549 GND.n663 240.244
R4980 GND.n5549 GND.n661 240.244
R4981 GND.n5553 GND.n661 240.244
R4982 GND.n5553 GND.n657 240.244
R4983 GND.n5559 GND.n657 240.244
R4984 GND.n5559 GND.n655 240.244
R4985 GND.n5563 GND.n655 240.244
R4986 GND.n5563 GND.n651 240.244
R4987 GND.n5569 GND.n651 240.244
R4988 GND.n5569 GND.n649 240.244
R4989 GND.n5573 GND.n649 240.244
R4990 GND.n5573 GND.n645 240.244
R4991 GND.n5579 GND.n645 240.244
R4992 GND.n5579 GND.n643 240.244
R4993 GND.n5583 GND.n643 240.244
R4994 GND.n5583 GND.n639 240.244
R4995 GND.n5589 GND.n639 240.244
R4996 GND.n5589 GND.n637 240.244
R4997 GND.n5593 GND.n637 240.244
R4998 GND.n5593 GND.n633 240.244
R4999 GND.n5599 GND.n633 240.244
R5000 GND.n5599 GND.n631 240.244
R5001 GND.n5603 GND.n631 240.244
R5002 GND.n5603 GND.n627 240.244
R5003 GND.n5609 GND.n627 240.244
R5004 GND.n5609 GND.n625 240.244
R5005 GND.n5613 GND.n625 240.244
R5006 GND.n5613 GND.n621 240.244
R5007 GND.n5619 GND.n621 240.244
R5008 GND.n5619 GND.n619 240.244
R5009 GND.n5623 GND.n619 240.244
R5010 GND.n5623 GND.n615 240.244
R5011 GND.n5629 GND.n615 240.244
R5012 GND.n5629 GND.n613 240.244
R5013 GND.n5633 GND.n613 240.244
R5014 GND.n5633 GND.n609 240.244
R5015 GND.n5639 GND.n609 240.244
R5016 GND.n5639 GND.n607 240.244
R5017 GND.n5643 GND.n607 240.244
R5018 GND.n5643 GND.n603 240.244
R5019 GND.n5650 GND.n603 240.244
R5020 GND.n5650 GND.n601 240.244
R5021 GND.n5655 GND.n601 240.244
R5022 GND.n5655 GND.n597 240.244
R5023 GND.n4886 GND.n1114 240.244
R5024 GND.n1626 GND.n1114 240.244
R5025 GND.n1626 GND.n1624 240.244
R5026 GND.n1632 GND.n1624 240.244
R5027 GND.n2007 GND.n1632 240.244
R5028 GND.n2008 GND.n2007 240.244
R5029 GND.n2008 GND.n1620 240.244
R5030 GND.n2016 GND.n1620 240.244
R5031 GND.n2016 GND.n1597 240.244
R5032 GND.n2045 GND.n1597 240.244
R5033 GND.n2046 GND.n2045 240.244
R5034 GND.n2046 GND.n1593 240.244
R5035 GND.n2052 GND.n1593 240.244
R5036 GND.n2052 GND.n1516 240.244
R5037 GND.n2136 GND.n1516 240.244
R5038 GND.n2136 GND.n1517 240.244
R5039 GND.n1537 GND.n1517 240.244
R5040 GND.n1540 GND.n1537 240.244
R5041 GND.n2122 GND.n1540 240.244
R5042 GND.n2122 GND.n2119 240.244
R5043 GND.n2119 GND.n1541 240.244
R5044 GND.n1569 GND.n1541 240.244
R5045 GND.n1569 GND.n1558 240.244
R5046 GND.n2105 GND.n1558 240.244
R5047 GND.n2105 GND.n2102 240.244
R5048 GND.n2102 GND.n1504 240.244
R5049 GND.n2194 GND.n1504 240.244
R5050 GND.n2194 GND.n1505 240.244
R5051 GND.n2190 GND.n1505 240.244
R5052 GND.n2190 GND.n2189 240.244
R5053 GND.n2189 GND.n2188 240.244
R5054 GND.n2188 GND.n2145 240.244
R5055 GND.n2184 GND.n2145 240.244
R5056 GND.n2184 GND.n2183 240.244
R5057 GND.n2183 GND.n2182 240.244
R5058 GND.n2182 GND.n2153 240.244
R5059 GND.n2178 GND.n2153 240.244
R5060 GND.n2178 GND.n2177 240.244
R5061 GND.n2177 GND.n2176 240.244
R5062 GND.n2176 GND.n2159 240.244
R5063 GND.n2172 GND.n2159 240.244
R5064 GND.n2172 GND.n2169 240.244
R5065 GND.n2169 GND.n1426 240.244
R5066 GND.n2288 GND.n1426 240.244
R5067 GND.n2289 GND.n2288 240.244
R5068 GND.n2290 GND.n2289 240.244
R5069 GND.n2290 GND.n1421 240.244
R5070 GND.n2305 GND.n1421 240.244
R5071 GND.n2305 GND.n1422 240.244
R5072 GND.n2301 GND.n1422 240.244
R5073 GND.n2301 GND.n2300 240.244
R5074 GND.n2300 GND.n1307 240.244
R5075 GND.n4709 GND.n1307 240.244
R5076 GND.n4709 GND.n1308 240.244
R5077 GND.n4705 GND.n1308 240.244
R5078 GND.n4705 GND.n1314 240.244
R5079 GND.n3399 GND.n1314 240.244
R5080 GND.n3412 GND.n3399 240.244
R5081 GND.n3412 GND.n3394 240.244
R5082 GND.n3418 GND.n3394 240.244
R5083 GND.n3418 GND.n3386 240.244
R5084 GND.n3432 GND.n3386 240.244
R5085 GND.n3432 GND.n3382 240.244
R5086 GND.n3438 GND.n3382 240.244
R5087 GND.n3438 GND.n3373 240.244
R5088 GND.n3452 GND.n3373 240.244
R5089 GND.n3452 GND.n3369 240.244
R5090 GND.n3458 GND.n3369 240.244
R5091 GND.n3458 GND.n3177 240.244
R5092 GND.n3473 GND.n3177 240.244
R5093 GND.n3473 GND.n3173 240.244
R5094 GND.n3479 GND.n3173 240.244
R5095 GND.n3479 GND.n3140 240.244
R5096 GND.n3507 GND.n3140 240.244
R5097 GND.n3507 GND.n3135 240.244
R5098 GND.n3515 GND.n3135 240.244
R5099 GND.n3515 GND.n3136 240.244
R5100 GND.n3136 GND.n3110 240.244
R5101 GND.n3549 GND.n3110 240.244
R5102 GND.n3549 GND.n3105 240.244
R5103 GND.n3572 GND.n3105 240.244
R5104 GND.n3572 GND.n3106 240.244
R5105 GND.n3568 GND.n3106 240.244
R5106 GND.n3568 GND.n3567 240.244
R5107 GND.n3567 GND.n3566 240.244
R5108 GND.n3566 GND.n3557 240.244
R5109 GND.n3562 GND.n3557 240.244
R5110 GND.n3562 GND.n3064 240.244
R5111 GND.n3665 GND.n3064 240.244
R5112 GND.n3665 GND.n3059 240.244
R5113 GND.n3673 GND.n3059 240.244
R5114 GND.n3673 GND.n3060 240.244
R5115 GND.n3060 GND.n3035 240.244
R5116 GND.n3709 GND.n3035 240.244
R5117 GND.n3709 GND.n3030 240.244
R5118 GND.n3720 GND.n3030 240.244
R5119 GND.n3720 GND.n3031 240.244
R5120 GND.n3716 GND.n3031 240.244
R5121 GND.n3716 GND.n2999 240.244
R5122 GND.n3769 GND.n2999 240.244
R5123 GND.n3769 GND.n2994 240.244
R5124 GND.n3777 GND.n2994 240.244
R5125 GND.n3777 GND.n2995 240.244
R5126 GND.n2995 GND.n2976 240.244
R5127 GND.n3794 GND.n2976 240.244
R5128 GND.n3794 GND.n2972 240.244
R5129 GND.n3800 GND.n2972 240.244
R5130 GND.n3800 GND.n2837 240.244
R5131 GND.n3897 GND.n2837 240.244
R5132 GND.n3897 GND.n2833 240.244
R5133 GND.n3903 GND.n2833 240.244
R5134 GND.n3903 GND.n2824 240.244
R5135 GND.n3916 GND.n2824 240.244
R5136 GND.n3916 GND.n2820 240.244
R5137 GND.n3922 GND.n2820 240.244
R5138 GND.n3922 GND.n2810 240.244
R5139 GND.n3935 GND.n2810 240.244
R5140 GND.n3935 GND.n2806 240.244
R5141 GND.n3943 GND.n2806 240.244
R5142 GND.n3943 GND.n2796 240.244
R5143 GND.n3956 GND.n2796 240.244
R5144 GND.n3957 GND.n3956 240.244
R5145 GND.n3957 GND.n2792 240.244
R5146 GND.n3963 GND.n2792 240.244
R5147 GND.n3963 GND.n2791 240.244
R5148 GND.n4024 GND.n2791 240.244
R5149 GND.n4024 GND.n2787 240.244
R5150 GND.n4030 GND.n2787 240.244
R5151 GND.n4031 GND.n4030 240.244
R5152 GND.n4032 GND.n4031 240.244
R5153 GND.n4032 GND.n2782 240.244
R5154 GND.n4106 GND.n2782 240.244
R5155 GND.n4106 GND.n2783 240.244
R5156 GND.n4102 GND.n2783 240.244
R5157 GND.n4102 GND.n4101 240.244
R5158 GND.n4101 GND.n4100 240.244
R5159 GND.n4100 GND.n4040 240.244
R5160 GND.n4096 GND.n4040 240.244
R5161 GND.n4096 GND.n4095 240.244
R5162 GND.n4095 GND.n4094 240.244
R5163 GND.n4094 GND.n4046 240.244
R5164 GND.n4090 GND.n4046 240.244
R5165 GND.n4090 GND.n4089 240.244
R5166 GND.n4089 GND.n4088 240.244
R5167 GND.n4088 GND.n4052 240.244
R5168 GND.n4084 GND.n4052 240.244
R5169 GND.n4084 GND.n4083 240.244
R5170 GND.n4083 GND.n4082 240.244
R5171 GND.n4082 GND.n4058 240.244
R5172 GND.n4078 GND.n4058 240.244
R5173 GND.n4078 GND.n4077 240.244
R5174 GND.n4077 GND.n4076 240.244
R5175 GND.n4076 GND.n4064 240.244
R5176 GND.n4072 GND.n4064 240.244
R5177 GND.n4072 GND.n4071 240.244
R5178 GND.n4071 GND.n2716 240.244
R5179 GND.n4321 GND.n2716 240.244
R5180 GND.n4321 GND.n2717 240.244
R5181 GND.n4316 GND.n2717 240.244
R5182 GND.n4316 GND.n2720 240.244
R5183 GND.n2734 GND.n2720 240.244
R5184 GND.n4306 GND.n2734 240.244
R5185 GND.n4306 GND.n2735 240.244
R5186 GND.n4301 GND.n2735 240.244
R5187 GND.n4301 GND.n4300 240.244
R5188 GND.n4300 GND.n4299 240.244
R5189 GND.n4299 GND.n4271 240.244
R5190 GND.n4295 GND.n4271 240.244
R5191 GND.n4295 GND.n4294 240.244
R5192 GND.n4294 GND.n4293 240.244
R5193 GND.n4293 GND.n4277 240.244
R5194 GND.n4289 GND.n4277 240.244
R5195 GND.n4289 GND.n4288 240.244
R5196 GND.n4288 GND.n4287 240.244
R5197 GND.n4287 GND.n590 240.244
R5198 GND.n5667 GND.n590 240.244
R5199 GND.n5667 GND.n591 240.244
R5200 GND.n5663 GND.n591 240.244
R5201 GND.n5663 GND.n5662 240.244
R5202 GND.n5662 GND.n5661 240.244
R5203 GND.n5028 GND.n974 240.244
R5204 GND.n5024 GND.n974 240.244
R5205 GND.n5024 GND.n979 240.244
R5206 GND.n5020 GND.n979 240.244
R5207 GND.n5020 GND.n981 240.244
R5208 GND.n5016 GND.n981 240.244
R5209 GND.n5016 GND.n987 240.244
R5210 GND.n5012 GND.n987 240.244
R5211 GND.n5012 GND.n989 240.244
R5212 GND.n5008 GND.n989 240.244
R5213 GND.n5008 GND.n995 240.244
R5214 GND.n5004 GND.n995 240.244
R5215 GND.n5004 GND.n997 240.244
R5216 GND.n5000 GND.n997 240.244
R5217 GND.n5000 GND.n1003 240.244
R5218 GND.n4996 GND.n1003 240.244
R5219 GND.n4996 GND.n1005 240.244
R5220 GND.n4992 GND.n1005 240.244
R5221 GND.n4992 GND.n1011 240.244
R5222 GND.n4988 GND.n1011 240.244
R5223 GND.n4988 GND.n1013 240.244
R5224 GND.n4984 GND.n1013 240.244
R5225 GND.n4984 GND.n1019 240.244
R5226 GND.n4980 GND.n1019 240.244
R5227 GND.n4980 GND.n1021 240.244
R5228 GND.n4976 GND.n1021 240.244
R5229 GND.n4976 GND.n1027 240.244
R5230 GND.n4972 GND.n1027 240.244
R5231 GND.n4972 GND.n1029 240.244
R5232 GND.n4968 GND.n1029 240.244
R5233 GND.n4968 GND.n1035 240.244
R5234 GND.n4964 GND.n1035 240.244
R5235 GND.n4964 GND.n1037 240.244
R5236 GND.n4960 GND.n1037 240.244
R5237 GND.n4960 GND.n1043 240.244
R5238 GND.n4956 GND.n1043 240.244
R5239 GND.n4956 GND.n1045 240.244
R5240 GND.n4952 GND.n1045 240.244
R5241 GND.n4952 GND.n1051 240.244
R5242 GND.n4948 GND.n1051 240.244
R5243 GND.n4948 GND.n1053 240.244
R5244 GND.n4944 GND.n1053 240.244
R5245 GND.n4944 GND.n1059 240.244
R5246 GND.n4940 GND.n1059 240.244
R5247 GND.n4940 GND.n1061 240.244
R5248 GND.n4936 GND.n1061 240.244
R5249 GND.n4936 GND.n1067 240.244
R5250 GND.n4932 GND.n1067 240.244
R5251 GND.n4932 GND.n1069 240.244
R5252 GND.n4928 GND.n1069 240.244
R5253 GND.n4928 GND.n1075 240.244
R5254 GND.n4924 GND.n1075 240.244
R5255 GND.n4924 GND.n1077 240.244
R5256 GND.n4920 GND.n1077 240.244
R5257 GND.n4920 GND.n1083 240.244
R5258 GND.n4916 GND.n1083 240.244
R5259 GND.n4916 GND.n1085 240.244
R5260 GND.n4912 GND.n1085 240.244
R5261 GND.n4912 GND.n1091 240.244
R5262 GND.n4908 GND.n1091 240.244
R5263 GND.n4908 GND.n1093 240.244
R5264 GND.n4904 GND.n1093 240.244
R5265 GND.n4904 GND.n1099 240.244
R5266 GND.n4900 GND.n1099 240.244
R5267 GND.n4900 GND.n1101 240.244
R5268 GND.n4896 GND.n1101 240.244
R5269 GND.n4896 GND.n1107 240.244
R5270 GND.n4892 GND.n1107 240.244
R5271 GND.n4892 GND.n1109 240.244
R5272 GND.n3966 GND.n2436 240.244
R5273 GND.n2445 GND.n2444 240.244
R5274 GND.n3968 GND.n2452 240.244
R5275 GND.n3971 GND.n2453 240.244
R5276 GND.n2461 GND.n2460 240.244
R5277 GND.n3973 GND.n2468 240.244
R5278 GND.n3976 GND.n2469 240.244
R5279 GND.n2477 GND.n2476 240.244
R5280 GND.n3995 GND.n3994 240.244
R5281 GND.n3999 GND.n3998 240.244
R5282 GND.n4007 GND.n4006 240.244
R5283 GND.n4012 GND.n3982 240.244
R5284 GND.n4019 GND.n2427 240.244
R5285 GND.n2347 GND.n2346 240.244
R5286 GND.n2348 GND.n2347 240.244
R5287 GND.n3420 GND.n2348 240.244
R5288 GND.n3420 GND.n2351 240.244
R5289 GND.n2352 GND.n2351 240.244
R5290 GND.n2353 GND.n2352 240.244
R5291 GND.n3440 GND.n2353 240.244
R5292 GND.n3440 GND.n2356 240.244
R5293 GND.n2357 GND.n2356 240.244
R5294 GND.n2358 GND.n2357 240.244
R5295 GND.n3460 GND.n2358 240.244
R5296 GND.n3460 GND.n2361 240.244
R5297 GND.n2362 GND.n2361 240.244
R5298 GND.n2363 GND.n2362 240.244
R5299 GND.n3481 GND.n2363 240.244
R5300 GND.n3481 GND.n2366 240.244
R5301 GND.n2367 GND.n2366 240.244
R5302 GND.n2368 GND.n2367 240.244
R5303 GND.n3127 GND.n2368 240.244
R5304 GND.n3127 GND.n2371 240.244
R5305 GND.n2372 GND.n2371 240.244
R5306 GND.n2373 GND.n2372 240.244
R5307 GND.n3101 GND.n2373 240.244
R5308 GND.n3101 GND.n2376 240.244
R5309 GND.n2377 GND.n2376 240.244
R5310 GND.n2378 GND.n2377 240.244
R5311 GND.n3589 GND.n2378 240.244
R5312 GND.n3589 GND.n2381 240.244
R5313 GND.n2382 GND.n2381 240.244
R5314 GND.n2383 GND.n2382 240.244
R5315 GND.n3635 GND.n2383 240.244
R5316 GND.n3635 GND.n2386 240.244
R5317 GND.n2387 GND.n2386 240.244
R5318 GND.n2388 GND.n2387 240.244
R5319 GND.n3623 GND.n2388 240.244
R5320 GND.n3623 GND.n2391 240.244
R5321 GND.n2392 GND.n2391 240.244
R5322 GND.n2393 GND.n2392 240.244
R5323 GND.n3690 GND.n2393 240.244
R5324 GND.n3690 GND.n2396 240.244
R5325 GND.n2397 GND.n2396 240.244
R5326 GND.n2398 GND.n2397 240.244
R5327 GND.n3000 GND.n2398 240.244
R5328 GND.n3000 GND.n2401 240.244
R5329 GND.n2402 GND.n2401 240.244
R5330 GND.n2403 GND.n2402 240.244
R5331 GND.n2977 GND.n2403 240.244
R5332 GND.n2977 GND.n2406 240.244
R5333 GND.n2407 GND.n2406 240.244
R5334 GND.n2408 GND.n2407 240.244
R5335 GND.n2895 GND.n2408 240.244
R5336 GND.n2895 GND.n2411 240.244
R5337 GND.n2412 GND.n2411 240.244
R5338 GND.n2413 GND.n2412 240.244
R5339 GND.n2826 GND.n2413 240.244
R5340 GND.n2826 GND.n2416 240.244
R5341 GND.n2417 GND.n2416 240.244
R5342 GND.n2418 GND.n2417 240.244
R5343 GND.n2812 GND.n2418 240.244
R5344 GND.n2812 GND.n2421 240.244
R5345 GND.n2422 GND.n2421 240.244
R5346 GND.n2423 GND.n2422 240.244
R5347 GND.n2797 GND.n2423 240.244
R5348 GND.n2797 GND.n2426 240.244
R5349 GND.n4540 GND.n2426 240.244
R5350 GND.n1329 GND.n1328 240.244
R5351 GND.n1341 GND.n1328 240.244
R5352 GND.n1343 GND.n1342 240.244
R5353 GND.n1351 GND.n1350 240.244
R5354 GND.n1361 GND.n1360 240.244
R5355 GND.n1363 GND.n1362 240.244
R5356 GND.n1371 GND.n1370 240.244
R5357 GND.n1381 GND.n1380 240.244
R5358 GND.n1383 GND.n1382 240.244
R5359 GND.n1395 GND.n1394 240.244
R5360 GND.n1397 GND.n1396 240.244
R5361 GND.n2340 GND.n2339 240.244
R5362 GND.n2342 GND.n2341 240.244
R5363 GND.n3409 GND.n1330 240.244
R5364 GND.n3409 GND.n3393 240.244
R5365 GND.n3423 GND.n3393 240.244
R5366 GND.n3423 GND.n3389 240.244
R5367 GND.n3429 GND.n3389 240.244
R5368 GND.n3429 GND.n3380 240.244
R5369 GND.n3443 GND.n3380 240.244
R5370 GND.n3443 GND.n3376 240.244
R5371 GND.n3449 GND.n3376 240.244
R5372 GND.n3449 GND.n3367 240.244
R5373 GND.n3464 GND.n3367 240.244
R5374 GND.n3464 GND.n3363 240.244
R5375 GND.n3470 GND.n3363 240.244
R5376 GND.n3470 GND.n3171 240.244
R5377 GND.n3483 GND.n3171 240.244
R5378 GND.n3483 GND.n3167 240.244
R5379 GND.n3489 GND.n3167 240.244
R5380 GND.n3489 GND.n3125 240.244
R5381 GND.n3526 GND.n3125 240.244
R5382 GND.n3526 GND.n3119 240.244
R5383 GND.n3539 GND.n3119 240.244
R5384 GND.n3539 GND.n3120 240.244
R5385 GND.n3531 GND.n3120 240.244
R5386 GND.n3532 GND.n3531 240.244
R5387 GND.n3532 GND.n3088 240.244
R5388 GND.n3599 GND.n3088 240.244
R5389 GND.n3599 GND.n3084 240.244
R5390 GND.n3605 GND.n3084 240.244
R5391 GND.n3605 GND.n3071 240.244
R5392 GND.n3656 GND.n3071 240.244
R5393 GND.n3656 GND.n3067 240.244
R5394 GND.n3662 GND.n3067 240.244
R5395 GND.n3662 GND.n3050 240.244
R5396 GND.n3684 GND.n3050 240.244
R5397 GND.n3684 GND.n3044 240.244
R5398 GND.n3699 GND.n3044 240.244
R5399 GND.n3699 GND.n3045 240.244
R5400 GND.n3689 GND.n3045 240.244
R5401 GND.n3692 GND.n3689 240.244
R5402 GND.n3692 GND.n3008 240.244
R5403 GND.n3750 GND.n3008 240.244
R5404 GND.n3750 GND.n3002 240.244
R5405 GND.n3766 GND.n3002 240.244
R5406 GND.n3766 GND.n3003 240.244
R5407 GND.n3755 GND.n3003 240.244
R5408 GND.n3756 GND.n3755 240.244
R5409 GND.n3757 GND.n3756 240.244
R5410 GND.n3757 GND.n2900 240.244
R5411 GND.n3819 GND.n2900 240.244
R5412 GND.n3819 GND.n2896 240.244
R5413 GND.n3825 GND.n2896 240.244
R5414 GND.n3825 GND.n2831 240.244
R5415 GND.n3906 GND.n2831 240.244
R5416 GND.n3906 GND.n2827 240.244
R5417 GND.n3912 GND.n2827 240.244
R5418 GND.n3912 GND.n2817 240.244
R5419 GND.n3925 GND.n2817 240.244
R5420 GND.n3925 GND.n2813 240.244
R5421 GND.n3931 GND.n2813 240.244
R5422 GND.n3931 GND.n2802 240.244
R5423 GND.n3946 GND.n2802 240.244
R5424 GND.n3946 GND.n2798 240.244
R5425 GND.n3952 GND.n2798 240.244
R5426 GND.n3952 GND.n2430 240.244
R5427 GND.n4538 GND.n2430 240.244
R5428 GND.n3188 GND.n3187 240.132
R5429 GND.n2883 GND.n2882 240.132
R5430 GND.n2336 GND.t72 224.174
R5431 GND.n4009 GND.t81 224.174
R5432 GND.n3220 GND.t20 204.78
R5433 GND.n2908 GND.t30 204.78
R5434 GND.n3216 GND.t10 204.78
R5435 GND.n3832 GND.t61 204.78
R5436 GND.n2537 GND.n2491 199.319
R5437 GND.n2537 GND.n2492 199.319
R5438 GND.n4726 GND.n1266 199.319
R5439 GND.n4724 GND.n1266 199.319
R5440 GND.n3189 GND.n3186 186.49
R5441 GND.n2884 GND.n2881 186.49
R5442 GND.n152 GND.n151 185
R5443 GND.n150 GND.n149 185
R5444 GND.n129 GND.n128 185
R5445 GND.n144 GND.n143 185
R5446 GND.n142 GND.n141 185
R5447 GND.n133 GND.n132 185
R5448 GND.n136 GND.n135 185
R5449 GND.n120 GND.n119 185
R5450 GND.n118 GND.n117 185
R5451 GND.n97 GND.n96 185
R5452 GND.n112 GND.n111 185
R5453 GND.n110 GND.n109 185
R5454 GND.n101 GND.n100 185
R5455 GND.n104 GND.n103 185
R5456 GND.n88 GND.n87 185
R5457 GND.n86 GND.n85 185
R5458 GND.n65 GND.n64 185
R5459 GND.n80 GND.n79 185
R5460 GND.n78 GND.n77 185
R5461 GND.n69 GND.n68 185
R5462 GND.n72 GND.n71 185
R5463 GND.n57 GND.n56 185
R5464 GND.n55 GND.n54 185
R5465 GND.n34 GND.n33 185
R5466 GND.n49 GND.n48 185
R5467 GND.n47 GND.n46 185
R5468 GND.n38 GND.n37 185
R5469 GND.n41 GND.n40 185
R5470 GND.n279 GND.n278 185
R5471 GND.n277 GND.n276 185
R5472 GND.n256 GND.n255 185
R5473 GND.n271 GND.n270 185
R5474 GND.n269 GND.n268 185
R5475 GND.n260 GND.n259 185
R5476 GND.n263 GND.n262 185
R5477 GND.n247 GND.n246 185
R5478 GND.n245 GND.n244 185
R5479 GND.n224 GND.n223 185
R5480 GND.n239 GND.n238 185
R5481 GND.n237 GND.n236 185
R5482 GND.n228 GND.n227 185
R5483 GND.n231 GND.n230 185
R5484 GND.n215 GND.n214 185
R5485 GND.n213 GND.n212 185
R5486 GND.n192 GND.n191 185
R5487 GND.n207 GND.n206 185
R5488 GND.n205 GND.n204 185
R5489 GND.n196 GND.n195 185
R5490 GND.n199 GND.n198 185
R5491 GND.n184 GND.n183 185
R5492 GND.n182 GND.n181 185
R5493 GND.n161 GND.n160 185
R5494 GND.n176 GND.n175 185
R5495 GND.n174 GND.n173 185
R5496 GND.n165 GND.n164 185
R5497 GND.n168 GND.n167 185
R5498 GND.n3221 GND.t19 178.987
R5499 GND.n2909 GND.t31 178.987
R5500 GND.n2337 GND.t71 178.987
R5501 GND.n3217 GND.t9 178.987
R5502 GND.n3833 GND.t62 178.987
R5503 GND.n4010 GND.t82 178.987
R5504 GND.n5482 GND.n698 176.212
R5505 GND.n5490 GND.n698 176.212
R5506 GND.n5491 GND.n5490 176.212
R5507 GND.n5492 GND.n5491 176.212
R5508 GND.n5492 GND.n692 176.212
R5509 GND.n5500 GND.n692 176.212
R5510 GND.n5501 GND.n5500 176.212
R5511 GND.n5502 GND.n5501 176.212
R5512 GND.n5502 GND.n686 176.212
R5513 GND.n5510 GND.n686 176.212
R5514 GND.n5511 GND.n5510 176.212
R5515 GND.n5512 GND.n5511 176.212
R5516 GND.n5512 GND.n680 176.212
R5517 GND.n5520 GND.n680 176.212
R5518 GND.n5521 GND.n5520 176.212
R5519 GND.n5522 GND.n5521 176.212
R5520 GND.n5522 GND.n674 176.212
R5521 GND.n5530 GND.n674 176.212
R5522 GND.n5531 GND.n5530 176.212
R5523 GND.n5532 GND.n5531 176.212
R5524 GND.n5532 GND.n668 176.212
R5525 GND.n5540 GND.n668 176.212
R5526 GND.n5541 GND.n5540 176.212
R5527 GND.n5542 GND.n5541 176.212
R5528 GND.n5542 GND.n662 176.212
R5529 GND.n5550 GND.n662 176.212
R5530 GND.n5551 GND.n5550 176.212
R5531 GND.n5552 GND.n5551 176.212
R5532 GND.n5552 GND.n656 176.212
R5533 GND.n5560 GND.n656 176.212
R5534 GND.n5561 GND.n5560 176.212
R5535 GND.n5562 GND.n5561 176.212
R5536 GND.n5562 GND.n650 176.212
R5537 GND.n5570 GND.n650 176.212
R5538 GND.n5571 GND.n5570 176.212
R5539 GND.n5572 GND.n5571 176.212
R5540 GND.n5572 GND.n644 176.212
R5541 GND.n5580 GND.n644 176.212
R5542 GND.n5581 GND.n5580 176.212
R5543 GND.n5582 GND.n5581 176.212
R5544 GND.n5582 GND.n638 176.212
R5545 GND.n5590 GND.n638 176.212
R5546 GND.n5591 GND.n5590 176.212
R5547 GND.n5592 GND.n5591 176.212
R5548 GND.n5592 GND.n632 176.212
R5549 GND.n5600 GND.n632 176.212
R5550 GND.n5601 GND.n5600 176.212
R5551 GND.n5602 GND.n5601 176.212
R5552 GND.n5602 GND.n626 176.212
R5553 GND.n5610 GND.n626 176.212
R5554 GND.n5611 GND.n5610 176.212
R5555 GND.n5612 GND.n5611 176.212
R5556 GND.n5612 GND.n620 176.212
R5557 GND.n5620 GND.n620 176.212
R5558 GND.n5621 GND.n5620 176.212
R5559 GND.n5622 GND.n5621 176.212
R5560 GND.n5622 GND.n614 176.212
R5561 GND.n5630 GND.n614 176.212
R5562 GND.n5631 GND.n5630 176.212
R5563 GND.n5632 GND.n5631 176.212
R5564 GND.n5632 GND.n608 176.212
R5565 GND.n5640 GND.n608 176.212
R5566 GND.n5641 GND.n5640 176.212
R5567 GND.n5642 GND.n5641 176.212
R5568 GND.n5642 GND.n602 176.212
R5569 GND.n5651 GND.n602 176.212
R5570 GND.n5652 GND.n5651 176.212
R5571 GND.n5654 GND.n5652 176.212
R5572 GND.n5654 GND.n5653 176.212
R5573 GND.n3892 GND.n2871 163.367
R5574 GND.n3888 GND.n3887 163.367
R5575 GND.n3884 GND.n3883 163.367
R5576 GND.n3880 GND.n3879 163.367
R5577 GND.n3876 GND.n3875 163.367
R5578 GND.n3872 GND.n3871 163.367
R5579 GND.n3868 GND.n3867 163.367
R5580 GND.n3864 GND.n3863 163.367
R5581 GND.n3860 GND.n3859 163.367
R5582 GND.n3856 GND.n3855 163.367
R5583 GND.n3852 GND.n3851 163.367
R5584 GND.n3848 GND.n3847 163.367
R5585 GND.n3844 GND.n3843 163.367
R5586 GND.n3839 GND.n3838 163.367
R5587 GND.n3835 GND.n3834 163.367
R5588 GND.n2913 GND.n2912 163.367
R5589 GND.n2917 GND.n2916 163.367
R5590 GND.n2921 GND.n2920 163.367
R5591 GND.n2925 GND.n2924 163.367
R5592 GND.n2929 GND.n2928 163.367
R5593 GND.n2933 GND.n2932 163.367
R5594 GND.n2937 GND.n2936 163.367
R5595 GND.n2941 GND.n2940 163.367
R5596 GND.n2945 GND.n2944 163.367
R5597 GND.n2949 GND.n2948 163.367
R5598 GND.n2953 GND.n2952 163.367
R5599 GND.n2957 GND.n2956 163.367
R5600 GND.n2961 GND.n2960 163.367
R5601 GND.n2965 GND.n2964 163.367
R5602 GND.n3236 GND.n3179 163.367
R5603 GND.n3236 GND.n3146 163.367
R5604 GND.n3496 GND.n3146 163.367
R5605 GND.n3496 GND.n3142 163.367
R5606 GND.n3492 GND.n3142 163.367
R5607 GND.n3492 GND.n3134 163.367
R5608 GND.n3164 GND.n3134 163.367
R5609 GND.n3164 GND.n3128 163.367
R5610 GND.n3161 GND.n3128 163.367
R5611 GND.n3161 GND.n3118 163.367
R5612 GND.n3156 GND.n3118 163.367
R5613 GND.n3156 GND.n3112 163.367
R5614 GND.n3153 GND.n3112 163.367
R5615 GND.n3153 GND.n3103 163.367
R5616 GND.n3148 GND.n3103 163.367
R5617 GND.n3148 GND.n3096 163.367
R5618 GND.n3583 GND.n3096 163.367
R5619 GND.n3583 GND.n3090 163.367
R5620 GND.n3587 GND.n3090 163.367
R5621 GND.n3587 GND.n3082 163.367
R5622 GND.n3608 GND.n3082 163.367
R5623 GND.n3608 GND.n3080 163.367
R5624 GND.n3642 GND.n3080 163.367
R5625 GND.n3642 GND.n3073 163.367
R5626 GND.n3638 GND.n3073 163.367
R5627 GND.n3638 GND.n3634 163.367
R5628 GND.n3634 GND.n3633 163.367
R5629 GND.n3633 GND.n3058 163.367
R5630 GND.n3629 GND.n3058 163.367
R5631 GND.n3629 GND.n3052 163.367
R5632 GND.n3626 GND.n3052 163.367
R5633 GND.n3626 GND.n3043 163.367
R5634 GND.n3620 GND.n3043 163.367
R5635 GND.n3620 GND.n3037 163.367
R5636 GND.n3617 GND.n3037 163.367
R5637 GND.n3617 GND.n3028 163.367
R5638 GND.n3612 GND.n3028 163.367
R5639 GND.n3612 GND.n3022 163.367
R5640 GND.n3731 GND.n3022 163.367
R5641 GND.n3731 GND.n3010 163.367
R5642 GND.n3019 GND.n3010 163.367
R5643 GND.n3742 GND.n3019 163.367
R5644 GND.n3742 GND.n3020 163.367
R5645 GND.n3738 GND.n3020 163.367
R5646 GND.n3738 GND.n2991 163.367
R5647 GND.n2991 GND.n2981 163.367
R5648 GND.n3787 GND.n2981 163.367
R5649 GND.n3787 GND.n2979 163.367
R5650 GND.n3791 GND.n2979 163.367
R5651 GND.n3791 GND.n2906 163.367
R5652 GND.n3808 GND.n2906 163.367
R5653 GND.n3808 GND.n2902 163.367
R5654 GND.n3804 GND.n2902 163.367
R5655 GND.n3804 GND.n2894 163.367
R5656 GND.n2969 GND.n2894 163.367
R5657 GND.n3355 GND.n3353 163.367
R5658 GND.n3353 GND.n3352 163.367
R5659 GND.n3349 GND.n3348 163.367
R5660 GND.n3346 GND.n3205 163.367
R5661 GND.n3342 GND.n3340 163.367
R5662 GND.n3338 GND.n3207 163.367
R5663 GND.n3334 GND.n3332 163.367
R5664 GND.n3330 GND.n3209 163.367
R5665 GND.n3326 GND.n3324 163.367
R5666 GND.n3322 GND.n3211 163.367
R5667 GND.n3318 GND.n3316 163.367
R5668 GND.n3314 GND.n3213 163.367
R5669 GND.n3310 GND.n3308 163.367
R5670 GND.n3306 GND.n3215 163.367
R5671 GND.n3302 GND.n3300 163.367
R5672 GND.n3296 GND.n3219 163.367
R5673 GND.n3292 GND.n3290 163.367
R5674 GND.n3287 GND.n3286 163.367
R5675 GND.n3284 GND.n3225 163.367
R5676 GND.n3280 GND.n3278 163.367
R5677 GND.n3276 GND.n3227 163.367
R5678 GND.n3272 GND.n3270 163.367
R5679 GND.n3268 GND.n3229 163.367
R5680 GND.n3264 GND.n3262 163.367
R5681 GND.n3260 GND.n3231 163.367
R5682 GND.n3256 GND.n3254 163.367
R5683 GND.n3252 GND.n3233 163.367
R5684 GND.n3248 GND.n3246 163.367
R5685 GND.n3244 GND.n3235 163.367
R5686 GND.n3360 GND.n3145 163.367
R5687 GND.n3500 GND.n3145 163.367
R5688 GND.n3500 GND.n3143 163.367
R5689 GND.n3504 GND.n3143 163.367
R5690 GND.n3504 GND.n3132 163.367
R5691 GND.n3519 GND.n3132 163.367
R5692 GND.n3519 GND.n3130 163.367
R5693 GND.n3523 GND.n3130 163.367
R5694 GND.n3523 GND.n3116 163.367
R5695 GND.n3542 GND.n3116 163.367
R5696 GND.n3542 GND.n3114 163.367
R5697 GND.n3546 GND.n3114 163.367
R5698 GND.n3546 GND.n3100 163.367
R5699 GND.n3575 GND.n3100 163.367
R5700 GND.n3575 GND.n3098 163.367
R5701 GND.n3579 GND.n3098 163.367
R5702 GND.n3579 GND.n3092 163.367
R5703 GND.n3596 GND.n3092 163.367
R5704 GND.n3596 GND.n3093 163.367
R5705 GND.n3592 GND.n3093 163.367
R5706 GND.n3592 GND.n3078 163.367
R5707 GND.n3646 GND.n3078 163.367
R5708 GND.n3646 GND.n3075 163.367
R5709 GND.n3653 GND.n3075 163.367
R5710 GND.n3653 GND.n3076 163.367
R5711 GND.n3649 GND.n3076 163.367
R5712 GND.n3649 GND.n3056 163.367
R5713 GND.n3677 GND.n3056 163.367
R5714 GND.n3677 GND.n3054 163.367
R5715 GND.n3681 GND.n3054 163.367
R5716 GND.n3681 GND.n3041 163.367
R5717 GND.n3702 GND.n3041 163.367
R5718 GND.n3702 GND.n3039 163.367
R5719 GND.n3706 GND.n3039 163.367
R5720 GND.n3706 GND.n3026 163.367
R5721 GND.n3723 GND.n3026 163.367
R5722 GND.n3723 GND.n3024 163.367
R5723 GND.n3727 GND.n3024 163.367
R5724 GND.n3727 GND.n3012 163.367
R5725 GND.n3748 GND.n3012 163.367
R5726 GND.n3748 GND.n3013 163.367
R5727 GND.n3744 GND.n3013 163.367
R5728 GND.n3744 GND.n3016 163.367
R5729 GND.n3016 GND.n2989 163.367
R5730 GND.n3780 GND.n2989 163.367
R5731 GND.n3780 GND.n2984 163.367
R5732 GND.n3785 GND.n2984 163.367
R5733 GND.n3785 GND.n2987 163.367
R5734 GND.n2987 GND.n2905 163.367
R5735 GND.n3812 GND.n2905 163.367
R5736 GND.n3812 GND.n2903 163.367
R5737 GND.n3816 GND.n2903 163.367
R5738 GND.n3816 GND.n2892 163.367
R5739 GND.n3828 GND.n2892 163.367
R5740 GND.n3828 GND.n2870 163.367
R5741 GND.n2890 GND.n2889 156.462
R5742 GND.n92 GND.n60 153.042
R5743 GND.n156 GND.n155 152.079
R5744 GND.n124 GND.n123 152.079
R5745 GND.n92 GND.n91 152.079
R5746 GND.n3194 GND.n3193 152
R5747 GND.n3195 GND.n3184 152
R5748 GND.n3197 GND.n3196 152
R5749 GND.n3199 GND.n3182 152
R5750 GND.n3201 GND.n3200 152
R5751 GND.n2888 GND.n2872 152
R5752 GND.n2880 GND.n2873 152
R5753 GND.n2879 GND.n2878 152
R5754 GND.n2877 GND.n2874 152
R5755 GND.n2875 GND.t73 150.546
R5756 GND.t108 GND.n134 147.661
R5757 GND.t110 GND.n102 147.661
R5758 GND.t106 GND.n70 147.661
R5759 GND.t104 GND.n39 147.661
R5760 GND.t94 GND.n261 147.661
R5761 GND.t102 GND.n229 147.661
R5762 GND.t114 GND.n197 147.661
R5763 GND.t112 GND.n166 147.661
R5764 GND.n2855 GND.n2854 143.351
R5765 GND.n2854 GND.n2853 143.351
R5766 GND.n3299 GND.n3298 143.351
R5767 GND.n3298 GND.n3297 143.351
R5768 GND.n3191 GND.t15 130.484
R5769 GND.n3200 GND.t54 126.766
R5770 GND.n3198 GND.t63 126.766
R5771 GND.n3184 GND.t45 126.766
R5772 GND.n3192 GND.t83 126.766
R5773 GND.n2876 GND.t21 126.766
R5774 GND.n2878 GND.t4 126.766
R5775 GND.n2887 GND.t48 126.766
R5776 GND.n2889 GND.t66 126.766
R5777 GND.n1264 GND.t52 118.023
R5778 GND.n1292 GND.t13 118.023
R5779 GND.n4486 GND.t37 118.023
R5780 GND.n1387 GND.t33 118.023
R5781 GND.n1802 GND.t88 118.023
R5782 GND.n2539 GND.t3 118.023
R5783 GND.n2561 GND.t44 118.023
R5784 GND.n541 GND.t40 118.023
R5785 GND.n5796 GND.t90 118.023
R5786 GND.n575 GND.t77 118.023
R5787 GND.n1727 GND.t27 118.023
R5788 GND.n1759 GND.t59 118.023
R5789 GND.n4771 GND.n1267 110.912
R5790 GND.n4451 GND.n2536 110.912
R5791 GND.n151 GND.n150 104.615
R5792 GND.n150 GND.n128 104.615
R5793 GND.n143 GND.n128 104.615
R5794 GND.n143 GND.n142 104.615
R5795 GND.n142 GND.n132 104.615
R5796 GND.n135 GND.n132 104.615
R5797 GND.n119 GND.n118 104.615
R5798 GND.n118 GND.n96 104.615
R5799 GND.n111 GND.n96 104.615
R5800 GND.n111 GND.n110 104.615
R5801 GND.n110 GND.n100 104.615
R5802 GND.n103 GND.n100 104.615
R5803 GND.n87 GND.n86 104.615
R5804 GND.n86 GND.n64 104.615
R5805 GND.n79 GND.n64 104.615
R5806 GND.n79 GND.n78 104.615
R5807 GND.n78 GND.n68 104.615
R5808 GND.n71 GND.n68 104.615
R5809 GND.n56 GND.n55 104.615
R5810 GND.n55 GND.n33 104.615
R5811 GND.n48 GND.n33 104.615
R5812 GND.n48 GND.n47 104.615
R5813 GND.n47 GND.n37 104.615
R5814 GND.n40 GND.n37 104.615
R5815 GND.n278 GND.n277 104.615
R5816 GND.n277 GND.n255 104.615
R5817 GND.n270 GND.n255 104.615
R5818 GND.n270 GND.n269 104.615
R5819 GND.n269 GND.n259 104.615
R5820 GND.n262 GND.n259 104.615
R5821 GND.n246 GND.n245 104.615
R5822 GND.n245 GND.n223 104.615
R5823 GND.n238 GND.n223 104.615
R5824 GND.n238 GND.n237 104.615
R5825 GND.n237 GND.n227 104.615
R5826 GND.n230 GND.n227 104.615
R5827 GND.n214 GND.n213 104.615
R5828 GND.n213 GND.n191 104.615
R5829 GND.n206 GND.n191 104.615
R5830 GND.n206 GND.n205 104.615
R5831 GND.n205 GND.n195 104.615
R5832 GND.n198 GND.n195 104.615
R5833 GND.n183 GND.n182 104.615
R5834 GND.n182 GND.n160 104.615
R5835 GND.n175 GND.n160 104.615
R5836 GND.n175 GND.n174 104.615
R5837 GND.n174 GND.n164 104.615
R5838 GND.n167 GND.n164 104.615
R5839 GND.n5825 GND.n478 99.6594
R5840 GND.n5823 GND.n5822 99.6594
R5841 GND.n5818 GND.n485 99.6594
R5842 GND.n5816 GND.n5815 99.6594
R5843 GND.n5811 GND.n492 99.6594
R5844 GND.n5809 GND.n5808 99.6594
R5845 GND.n5804 GND.n499 99.6594
R5846 GND.n5802 GND.n5801 99.6594
R5847 GND.n5794 GND.n506 99.6594
R5848 GND.n5792 GND.n5791 99.6594
R5849 GND.n5787 GND.n513 99.6594
R5850 GND.n5785 GND.n5784 99.6594
R5851 GND.n5780 GND.n520 99.6594
R5852 GND.n5778 GND.n5777 99.6594
R5853 GND.n5773 GND.n527 99.6594
R5854 GND.n5771 GND.n5770 99.6594
R5855 GND.n5766 GND.n534 99.6594
R5856 GND.n5764 GND.n5763 99.6594
R5857 GND.n539 GND.n538 99.6594
R5858 GND.n4482 GND.n4481 99.6594
R5859 GND.n4476 GND.n2485 99.6594
R5860 GND.n4473 GND.n2486 99.6594
R5861 GND.n4469 GND.n2487 99.6594
R5862 GND.n4465 GND.n2488 99.6594
R5863 GND.n4461 GND.n2489 99.6594
R5864 GND.n4457 GND.n2490 99.6594
R5865 GND.n4453 GND.n2491 99.6594
R5866 GND.n4448 GND.n2493 99.6594
R5867 GND.n4444 GND.n2494 99.6594
R5868 GND.n4440 GND.n2495 99.6594
R5869 GND.n4436 GND.n2496 99.6594
R5870 GND.n4432 GND.n2497 99.6594
R5871 GND.n4428 GND.n2498 99.6594
R5872 GND.n4424 GND.n2499 99.6594
R5873 GND.n4420 GND.n2500 99.6594
R5874 GND.n4416 GND.n2501 99.6594
R5875 GND.n2560 GND.n2502 99.6594
R5876 GND.n4736 GND.n1246 99.6594
R5877 GND.n4735 GND.n1249 99.6594
R5878 GND.n4733 GND.n1251 99.6594
R5879 GND.n4732 GND.n1254 99.6594
R5880 GND.n4730 GND.n1256 99.6594
R5881 GND.n4729 GND.n1259 99.6594
R5882 GND.n4727 GND.n1261 99.6594
R5883 GND.n4724 GND.n1268 99.6594
R5884 GND.n4723 GND.n4722 99.6594
R5885 GND.n4721 GND.n1273 99.6594
R5886 GND.n4720 GND.n4719 99.6594
R5887 GND.n4718 GND.n1278 99.6594
R5888 GND.n4717 GND.n4716 99.6594
R5889 GND.n4715 GND.n1283 99.6594
R5890 GND.n4714 GND.n4713 99.6594
R5891 GND.n4712 GND.n1288 99.6594
R5892 GND.n4711 GND.n1294 99.6594
R5893 GND.n4738 GND.n1235 99.6594
R5894 GND.n1909 GND.n1699 99.6594
R5895 GND.n1907 GND.n1703 99.6594
R5896 GND.n1903 GND.n1902 99.6594
R5897 GND.n1896 GND.n1708 99.6594
R5898 GND.n1895 GND.n1894 99.6594
R5899 GND.n1888 GND.n1714 99.6594
R5900 GND.n1887 GND.n1886 99.6594
R5901 GND.n1880 GND.n1720 99.6594
R5902 GND.n1879 GND.n1878 99.6594
R5903 GND.n1872 GND.n1726 99.6594
R5904 GND.n1871 GND.n1870 99.6594
R5905 GND.n1864 GND.n1735 99.6594
R5906 GND.n1863 GND.n1862 99.6594
R5907 GND.n1856 GND.n1741 99.6594
R5908 GND.n1855 GND.n1854 99.6594
R5909 GND.n1848 GND.n1747 99.6594
R5910 GND.n1847 GND.n1846 99.6594
R5911 GND.n1757 GND.n1753 99.6594
R5912 GND.n1836 GND.n1835 99.6594
R5913 GND.n5753 GND.n547 99.6594
R5914 GND.n5751 GND.n5750 99.6594
R5915 GND.n5746 GND.n554 99.6594
R5916 GND.n5744 GND.n5743 99.6594
R5917 GND.n5739 GND.n561 99.6594
R5918 GND.n5737 GND.n5736 99.6594
R5919 GND.n5732 GND.n568 99.6594
R5920 GND.n5730 GND.n5729 99.6594
R5921 GND.n573 GND.n572 99.6594
R5922 GND.n2569 GND.n2503 99.6594
R5923 GND.n2505 GND.n2441 99.6594
R5924 GND.n2506 GND.n2448 99.6594
R5925 GND.n2508 GND.n2507 99.6594
R5926 GND.n2510 GND.n2457 99.6594
R5927 GND.n2511 GND.n2464 99.6594
R5928 GND.n2513 GND.n2512 99.6594
R5929 GND.n2515 GND.n2473 99.6594
R5930 GND.n4484 GND.n2480 99.6594
R5931 GND.n1337 GND.n1297 99.6594
R5932 GND.n1346 GND.n1298 99.6594
R5933 GND.n1354 GND.n1299 99.6594
R5934 GND.n1356 GND.n1300 99.6594
R5935 GND.n1366 GND.n1301 99.6594
R5936 GND.n1374 GND.n1302 99.6594
R5937 GND.n1376 GND.n1303 99.6594
R5938 GND.n1386 GND.n1304 99.6594
R5939 GND.n4653 GND.n1305 99.6594
R5940 GND.n1831 GND.n1830 99.6594
R5941 GND.n1828 GND.n1770 99.6594
R5942 GND.n1775 GND.n1774 99.6594
R5943 GND.n1780 GND.n1777 99.6594
R5944 GND.n1783 GND.n1782 99.6594
R5945 GND.n1788 GND.n1785 99.6594
R5946 GND.n1791 GND.n1790 99.6594
R5947 GND.n1796 GND.n1793 99.6594
R5948 GND.n1800 GND.n1798 99.6594
R5949 GND.n1830 GND.n1829 99.6594
R5950 GND.n1773 GND.n1770 99.6594
R5951 GND.n1776 GND.n1775 99.6594
R5952 GND.n1781 GND.n1780 99.6594
R5953 GND.n1784 GND.n1783 99.6594
R5954 GND.n1789 GND.n1788 99.6594
R5955 GND.n1792 GND.n1791 99.6594
R5956 GND.n1797 GND.n1796 99.6594
R5957 GND.n1801 GND.n1800 99.6594
R5958 GND.n1390 GND.n1305 99.6594
R5959 GND.n1377 GND.n1304 99.6594
R5960 GND.n1375 GND.n1303 99.6594
R5961 GND.n1367 GND.n1302 99.6594
R5962 GND.n1357 GND.n1301 99.6594
R5963 GND.n1355 GND.n1300 99.6594
R5964 GND.n1347 GND.n1299 99.6594
R5965 GND.n1338 GND.n1298 99.6594
R5966 GND.n1336 GND.n1297 99.6594
R5967 GND.n2503 GND.n2440 99.6594
R5968 GND.n2505 GND.n2504 99.6594
R5969 GND.n2506 GND.n2449 99.6594
R5970 GND.n2508 GND.n2456 99.6594
R5971 GND.n2510 GND.n2509 99.6594
R5972 GND.n2511 GND.n2465 99.6594
R5973 GND.n2513 GND.n2472 99.6594
R5974 GND.n2515 GND.n2514 99.6594
R5975 GND.n4485 GND.n4484 99.6594
R5976 GND.n572 GND.n569 99.6594
R5977 GND.n5731 GND.n5730 99.6594
R5978 GND.n568 GND.n562 99.6594
R5979 GND.n5738 GND.n5737 99.6594
R5980 GND.n561 GND.n555 99.6594
R5981 GND.n5745 GND.n5744 99.6594
R5982 GND.n554 GND.n548 99.6594
R5983 GND.n5752 GND.n5751 99.6594
R5984 GND.n547 GND.n544 99.6594
R5985 GND.n1910 GND.n1909 99.6594
R5986 GND.n1904 GND.n1703 99.6594
R5987 GND.n1902 GND.n1901 99.6594
R5988 GND.n1897 GND.n1896 99.6594
R5989 GND.n1894 GND.n1893 99.6594
R5990 GND.n1889 GND.n1888 99.6594
R5991 GND.n1886 GND.n1885 99.6594
R5992 GND.n1881 GND.n1880 99.6594
R5993 GND.n1878 GND.n1877 99.6594
R5994 GND.n1873 GND.n1872 99.6594
R5995 GND.n1870 GND.n1869 99.6594
R5996 GND.n1865 GND.n1864 99.6594
R5997 GND.n1862 GND.n1861 99.6594
R5998 GND.n1857 GND.n1856 99.6594
R5999 GND.n1854 GND.n1853 99.6594
R6000 GND.n1849 GND.n1848 99.6594
R6001 GND.n1846 GND.n1845 99.6594
R6002 GND.n1758 GND.n1757 99.6594
R6003 GND.n1837 GND.n1836 99.6594
R6004 GND.n4739 GND.n4738 99.6594
R6005 GND.n4711 GND.n1289 99.6594
R6006 GND.n4712 GND.n1287 99.6594
R6007 GND.n4714 GND.n1284 99.6594
R6008 GND.n4715 GND.n1282 99.6594
R6009 GND.n4717 GND.n1279 99.6594
R6010 GND.n4718 GND.n1277 99.6594
R6011 GND.n4720 GND.n1274 99.6594
R6012 GND.n4721 GND.n1272 99.6594
R6013 GND.n4723 GND.n1269 99.6594
R6014 GND.n4726 GND.n4725 99.6594
R6015 GND.n4727 GND.n1260 99.6594
R6016 GND.n4729 GND.n4728 99.6594
R6017 GND.n4730 GND.n1255 99.6594
R6018 GND.n4732 GND.n4731 99.6594
R6019 GND.n4733 GND.n1250 99.6594
R6020 GND.n4735 GND.n4734 99.6594
R6021 GND.n4736 GND.n1245 99.6594
R6022 GND.n4482 GND.n2518 99.6594
R6023 GND.n4474 GND.n2485 99.6594
R6024 GND.n4470 GND.n2486 99.6594
R6025 GND.n4466 GND.n2487 99.6594
R6026 GND.n4462 GND.n2488 99.6594
R6027 GND.n4458 GND.n2489 99.6594
R6028 GND.n4454 GND.n2490 99.6594
R6029 GND.n4449 GND.n2492 99.6594
R6030 GND.n4445 GND.n2493 99.6594
R6031 GND.n4441 GND.n2494 99.6594
R6032 GND.n4437 GND.n2495 99.6594
R6033 GND.n4433 GND.n2496 99.6594
R6034 GND.n4429 GND.n2497 99.6594
R6035 GND.n4425 GND.n2498 99.6594
R6036 GND.n4421 GND.n2499 99.6594
R6037 GND.n4417 GND.n2500 99.6594
R6038 GND.n2559 GND.n2501 99.6594
R6039 GND.n4409 GND.n2502 99.6594
R6040 GND.n538 GND.n535 99.6594
R6041 GND.n5765 GND.n5764 99.6594
R6042 GND.n534 GND.n528 99.6594
R6043 GND.n5772 GND.n5771 99.6594
R6044 GND.n527 GND.n521 99.6594
R6045 GND.n5779 GND.n5778 99.6594
R6046 GND.n520 GND.n514 99.6594
R6047 GND.n5786 GND.n5785 99.6594
R6048 GND.n513 GND.n507 99.6594
R6049 GND.n5793 GND.n5792 99.6594
R6050 GND.n506 GND.n500 99.6594
R6051 GND.n5803 GND.n5802 99.6594
R6052 GND.n499 GND.n493 99.6594
R6053 GND.n5810 GND.n5809 99.6594
R6054 GND.n492 GND.n486 99.6594
R6055 GND.n5817 GND.n5816 99.6594
R6056 GND.n485 GND.n479 99.6594
R6057 GND.n5824 GND.n5823 99.6594
R6058 GND.n478 GND.n475 99.6594
R6059 GND.n3965 GND.n2431 99.6594
R6060 GND.n3967 GND.n3966 99.6594
R6061 GND.n3969 GND.n2445 99.6594
R6062 GND.n3970 GND.n2452 99.6594
R6063 GND.n3972 GND.n3971 99.6594
R6064 GND.n3974 GND.n2461 99.6594
R6065 GND.n3975 GND.n2468 99.6594
R6066 GND.n3977 GND.n3976 99.6594
R6067 GND.n3978 GND.n2477 99.6594
R6068 GND.n3995 GND.n3979 99.6594
R6069 GND.n3998 GND.n3980 99.6594
R6070 GND.n4007 GND.n3981 99.6594
R6071 GND.n4020 GND.n3982 99.6594
R6072 GND.n4020 GND.n4019 99.6594
R6073 GND.n4012 GND.n3981 99.6594
R6074 GND.n4006 GND.n3980 99.6594
R6075 GND.n3999 GND.n3979 99.6594
R6076 GND.n3994 GND.n3978 99.6594
R6077 GND.n3977 GND.n2476 99.6594
R6078 GND.n3975 GND.n2469 99.6594
R6079 GND.n3974 GND.n3973 99.6594
R6080 GND.n3972 GND.n2460 99.6594
R6081 GND.n3970 GND.n2453 99.6594
R6082 GND.n3969 GND.n3968 99.6594
R6083 GND.n3967 GND.n2444 99.6594
R6084 GND.n3965 GND.n2436 99.6594
R6085 GND.n4702 GND.n4701 99.6594
R6086 GND.n1341 GND.n1315 99.6594
R6087 GND.n1343 GND.n1316 99.6594
R6088 GND.n1351 GND.n1317 99.6594
R6089 GND.n1361 GND.n1318 99.6594
R6090 GND.n1363 GND.n1319 99.6594
R6091 GND.n1371 GND.n1320 99.6594
R6092 GND.n1381 GND.n1321 99.6594
R6093 GND.n1383 GND.n1322 99.6594
R6094 GND.n1395 GND.n1323 99.6594
R6095 GND.n1397 GND.n1324 99.6594
R6096 GND.n2340 GND.n1325 99.6594
R6097 GND.n2342 GND.n1326 99.6594
R6098 GND.n4702 GND.n1329 99.6594
R6099 GND.n1342 GND.n1315 99.6594
R6100 GND.n1350 GND.n1316 99.6594
R6101 GND.n1360 GND.n1317 99.6594
R6102 GND.n1362 GND.n1318 99.6594
R6103 GND.n1370 GND.n1319 99.6594
R6104 GND.n1380 GND.n1320 99.6594
R6105 GND.n1382 GND.n1321 99.6594
R6106 GND.n1394 GND.n1322 99.6594
R6107 GND.n1396 GND.n1323 99.6594
R6108 GND.n2339 GND.n1324 99.6594
R6109 GND.n2341 GND.n1325 99.6594
R6110 GND.n2345 GND.n1326 99.6594
R6111 GND.n5653 GND.n471 91.3564
R6112 GND.n3191 GND.n3190 81.8399
R6113 GND.n3192 GND.n3185 72.8411
R6114 GND.n3198 GND.n3183 72.8411
R6115 GND.n2887 GND.n2886 72.8411
R6116 GND.n1265 GND.t53 72.836
R6117 GND.n1293 GND.t14 72.836
R6118 GND.n4487 GND.t36 72.836
R6119 GND.n1388 GND.t34 72.836
R6120 GND.n1803 GND.t87 72.836
R6121 GND.n2540 GND.t2 72.836
R6122 GND.n2562 GND.t43 72.836
R6123 GND.n542 GND.t41 72.836
R6124 GND.n5797 GND.t91 72.836
R6125 GND.n576 GND.t78 72.836
R6126 GND.n1728 GND.t26 72.836
R6127 GND.n1760 GND.t58 72.836
R6128 GND.n3888 GND.n2869 71.676
R6129 GND.n3884 GND.n2868 71.676
R6130 GND.n3880 GND.n2867 71.676
R6131 GND.n3876 GND.n2866 71.676
R6132 GND.n3872 GND.n2865 71.676
R6133 GND.n3868 GND.n2864 71.676
R6134 GND.n3864 GND.n2863 71.676
R6135 GND.n3860 GND.n2862 71.676
R6136 GND.n3856 GND.n2861 71.676
R6137 GND.n3852 GND.n2860 71.676
R6138 GND.n3848 GND.n2859 71.676
R6139 GND.n3844 GND.n2858 71.676
R6140 GND.n3839 GND.n2857 71.676
R6141 GND.n3835 GND.n2856 71.676
R6142 GND.n2912 GND.n2853 71.676
R6143 GND.n2916 GND.n2852 71.676
R6144 GND.n2920 GND.n2851 71.676
R6145 GND.n2924 GND.n2850 71.676
R6146 GND.n2928 GND.n2849 71.676
R6147 GND.n2932 GND.n2848 71.676
R6148 GND.n2936 GND.n2847 71.676
R6149 GND.n2940 GND.n2846 71.676
R6150 GND.n2944 GND.n2845 71.676
R6151 GND.n2948 GND.n2844 71.676
R6152 GND.n2952 GND.n2843 71.676
R6153 GND.n2956 GND.n2842 71.676
R6154 GND.n2960 GND.n2841 71.676
R6155 GND.n2964 GND.n2840 71.676
R6156 GND.n2968 GND.n2839 71.676
R6157 GND.n3354 GND.n3181 71.676
R6158 GND.n3352 GND.n3203 71.676
R6159 GND.n3348 GND.n3347 71.676
R6160 GND.n3341 GND.n3205 71.676
R6161 GND.n3340 GND.n3339 71.676
R6162 GND.n3333 GND.n3207 71.676
R6163 GND.n3332 GND.n3331 71.676
R6164 GND.n3325 GND.n3209 71.676
R6165 GND.n3324 GND.n3323 71.676
R6166 GND.n3317 GND.n3211 71.676
R6167 GND.n3316 GND.n3315 71.676
R6168 GND.n3309 GND.n3213 71.676
R6169 GND.n3308 GND.n3307 71.676
R6170 GND.n3301 GND.n3215 71.676
R6171 GND.n3300 GND.n3299 71.676
R6172 GND.n3291 GND.n3219 71.676
R6173 GND.n3290 GND.n3223 71.676
R6174 GND.n3286 GND.n3285 71.676
R6175 GND.n3279 GND.n3225 71.676
R6176 GND.n3278 GND.n3277 71.676
R6177 GND.n3271 GND.n3227 71.676
R6178 GND.n3270 GND.n3269 71.676
R6179 GND.n3263 GND.n3229 71.676
R6180 GND.n3262 GND.n3261 71.676
R6181 GND.n3255 GND.n3231 71.676
R6182 GND.n3254 GND.n3253 71.676
R6183 GND.n3247 GND.n3233 71.676
R6184 GND.n3246 GND.n3245 71.676
R6185 GND.n3239 GND.n3235 71.676
R6186 GND.n3355 GND.n3354 71.676
R6187 GND.n3349 GND.n3203 71.676
R6188 GND.n3347 GND.n3346 71.676
R6189 GND.n3342 GND.n3341 71.676
R6190 GND.n3339 GND.n3338 71.676
R6191 GND.n3334 GND.n3333 71.676
R6192 GND.n3331 GND.n3330 71.676
R6193 GND.n3326 GND.n3325 71.676
R6194 GND.n3323 GND.n3322 71.676
R6195 GND.n3318 GND.n3317 71.676
R6196 GND.n3315 GND.n3314 71.676
R6197 GND.n3310 GND.n3309 71.676
R6198 GND.n3307 GND.n3306 71.676
R6199 GND.n3302 GND.n3301 71.676
R6200 GND.n3297 GND.n3296 71.676
R6201 GND.n3292 GND.n3291 71.676
R6202 GND.n3287 GND.n3223 71.676
R6203 GND.n3285 GND.n3284 71.676
R6204 GND.n3280 GND.n3279 71.676
R6205 GND.n3277 GND.n3276 71.676
R6206 GND.n3272 GND.n3271 71.676
R6207 GND.n3269 GND.n3268 71.676
R6208 GND.n3264 GND.n3263 71.676
R6209 GND.n3261 GND.n3260 71.676
R6210 GND.n3256 GND.n3255 71.676
R6211 GND.n3253 GND.n3252 71.676
R6212 GND.n3248 GND.n3247 71.676
R6213 GND.n3245 GND.n3244 71.676
R6214 GND.n3240 GND.n3239 71.676
R6215 GND.n2965 GND.n2839 71.676
R6216 GND.n2961 GND.n2840 71.676
R6217 GND.n2957 GND.n2841 71.676
R6218 GND.n2953 GND.n2842 71.676
R6219 GND.n2949 GND.n2843 71.676
R6220 GND.n2945 GND.n2844 71.676
R6221 GND.n2941 GND.n2845 71.676
R6222 GND.n2937 GND.n2846 71.676
R6223 GND.n2933 GND.n2847 71.676
R6224 GND.n2929 GND.n2848 71.676
R6225 GND.n2925 GND.n2849 71.676
R6226 GND.n2921 GND.n2850 71.676
R6227 GND.n2917 GND.n2851 71.676
R6228 GND.n2913 GND.n2852 71.676
R6229 GND.n3834 GND.n2855 71.676
R6230 GND.n3838 GND.n2856 71.676
R6231 GND.n3843 GND.n2857 71.676
R6232 GND.n3847 GND.n2858 71.676
R6233 GND.n3851 GND.n2859 71.676
R6234 GND.n3855 GND.n2860 71.676
R6235 GND.n3859 GND.n2861 71.676
R6236 GND.n3863 GND.n2862 71.676
R6237 GND.n3867 GND.n2863 71.676
R6238 GND.n3871 GND.n2864 71.676
R6239 GND.n3875 GND.n2865 71.676
R6240 GND.n3879 GND.n2866 71.676
R6241 GND.n3883 GND.n2867 71.676
R6242 GND.n3887 GND.n2868 71.676
R6243 GND.n2871 GND.n2869 71.676
R6244 GND.n1919 GND.n1696 60.6121
R6245 GND.n5833 GND.n471 60.6121
R6246 GND.n3222 GND.n3221 59.5399
R6247 GND.n2910 GND.n2909 59.5399
R6248 GND.n3218 GND.n3217 59.5399
R6249 GND.n3841 GND.n3833 59.5399
R6250 GND.n3358 GND.n3201 59.1804
R6251 GND.n10 GND.t118 56.8381
R6252 GND.n19 GND.t172 56.8381
R6253 GND.n1 GND.t131 56.8381
R6254 GND.n286 GND.t169 56.8381
R6255 GND.n295 GND.t192 56.8381
R6256 GND.n305 GND.t135 56.8381
R6257 GND.n17 GND.t178 55.8337
R6258 GND.n26 GND.t120 55.8337
R6259 GND.n8 GND.t145 55.8337
R6260 GND.n293 GND.t126 55.8337
R6261 GND.n302 GND.t170 55.8337
R6262 GND.n312 GND.t146 55.8337
R6263 GND.n3189 GND.n3188 54.358
R6264 GND.n2884 GND.n2883 54.358
R6265 GND.n10 GND.n9 53.0052
R6266 GND.n12 GND.n11 53.0052
R6267 GND.n14 GND.n13 53.0052
R6268 GND.n16 GND.n15 53.0052
R6269 GND.n19 GND.n18 53.0052
R6270 GND.n21 GND.n20 53.0052
R6271 GND.n23 GND.n22 53.0052
R6272 GND.n25 GND.n24 53.0052
R6273 GND.n1 GND.n0 53.0052
R6274 GND.n3 GND.n2 53.0052
R6275 GND.n5 GND.n4 53.0052
R6276 GND.n7 GND.n6 53.0052
R6277 GND.n292 GND.n291 53.0052
R6278 GND.n290 GND.n289 53.0052
R6279 GND.n288 GND.n287 53.0052
R6280 GND.n286 GND.n285 53.0052
R6281 GND.n301 GND.n300 53.0052
R6282 GND.n299 GND.n298 53.0052
R6283 GND.n297 GND.n296 53.0052
R6284 GND.n295 GND.n294 53.0052
R6285 GND.n311 GND.n310 53.0052
R6286 GND.n309 GND.n308 53.0052
R6287 GND.n307 GND.n306 53.0052
R6288 GND.n305 GND.n304 53.0052
R6289 GND.n2875 GND.n2874 52.4801
R6290 GND.n135 GND.t108 52.3082
R6291 GND.n103 GND.t110 52.3082
R6292 GND.n71 GND.t106 52.3082
R6293 GND.n40 GND.t104 52.3082
R6294 GND.n262 GND.t94 52.3082
R6295 GND.n230 GND.t102 52.3082
R6296 GND.n198 GND.t114 52.3082
R6297 GND.n167 GND.t112 52.3082
R6298 GND.n219 GND.n187 51.4173
R6299 GND.n283 GND.n282 50.455
R6300 GND.n251 GND.n250 50.455
R6301 GND.n219 GND.n218 50.455
R6302 GND.n5029 GND.n973 48.13
R6303 GND.n5023 GND.n973 48.13
R6304 GND.n5023 GND.n5022 48.13
R6305 GND.n5022 GND.n5021 48.13
R6306 GND.n5021 GND.n980 48.13
R6307 GND.n5015 GND.n980 48.13
R6308 GND.n5015 GND.n5014 48.13
R6309 GND.n5014 GND.n5013 48.13
R6310 GND.n5013 GND.n988 48.13
R6311 GND.n5007 GND.n988 48.13
R6312 GND.n5007 GND.n5006 48.13
R6313 GND.n5006 GND.n5005 48.13
R6314 GND.n5005 GND.n996 48.13
R6315 GND.n4999 GND.n996 48.13
R6316 GND.n4999 GND.n4998 48.13
R6317 GND.n4998 GND.n4997 48.13
R6318 GND.n4997 GND.n1004 48.13
R6319 GND.n4991 GND.n1004 48.13
R6320 GND.n4991 GND.n4990 48.13
R6321 GND.n4990 GND.n4989 48.13
R6322 GND.n4989 GND.n1012 48.13
R6323 GND.n4983 GND.n1012 48.13
R6324 GND.n4983 GND.n4982 48.13
R6325 GND.n4982 GND.n4981 48.13
R6326 GND.n4981 GND.n1020 48.13
R6327 GND.n4975 GND.n1020 48.13
R6328 GND.n4975 GND.n4974 48.13
R6329 GND.n4974 GND.n4973 48.13
R6330 GND.n4973 GND.n1028 48.13
R6331 GND.n4967 GND.n1028 48.13
R6332 GND.n4967 GND.n4966 48.13
R6333 GND.n4966 GND.n4965 48.13
R6334 GND.n4965 GND.n1036 48.13
R6335 GND.n4959 GND.n1036 48.13
R6336 GND.n4959 GND.n4958 48.13
R6337 GND.n4958 GND.n4957 48.13
R6338 GND.n4957 GND.n1044 48.13
R6339 GND.n4951 GND.n1044 48.13
R6340 GND.n4951 GND.n4950 48.13
R6341 GND.n4950 GND.n4949 48.13
R6342 GND.n4949 GND.n1052 48.13
R6343 GND.n4943 GND.n1052 48.13
R6344 GND.n4943 GND.n4942 48.13
R6345 GND.n4942 GND.n4941 48.13
R6346 GND.n4941 GND.n1060 48.13
R6347 GND.n4935 GND.n1060 48.13
R6348 GND.n4935 GND.n4934 48.13
R6349 GND.n4934 GND.n4933 48.13
R6350 GND.n4933 GND.n1068 48.13
R6351 GND.n4927 GND.n1068 48.13
R6352 GND.n4927 GND.n4926 48.13
R6353 GND.n4926 GND.n4925 48.13
R6354 GND.n4925 GND.n1076 48.13
R6355 GND.n4919 GND.n1076 48.13
R6356 GND.n4919 GND.n4918 48.13
R6357 GND.n4918 GND.n4917 48.13
R6358 GND.n4917 GND.n1084 48.13
R6359 GND.n4911 GND.n1084 48.13
R6360 GND.n4911 GND.n4910 48.13
R6361 GND.n4910 GND.n4909 48.13
R6362 GND.n4909 GND.n1092 48.13
R6363 GND.n4903 GND.n1092 48.13
R6364 GND.n4903 GND.n4902 48.13
R6365 GND.n4902 GND.n4901 48.13
R6366 GND.n4901 GND.n1100 48.13
R6367 GND.n4895 GND.n1100 48.13
R6368 GND.n4895 GND.n4894 48.13
R6369 GND.n4894 GND.n4893 48.13
R6370 GND.n4893 GND.n1108 48.13
R6371 GND.n2337 GND.n2336 45.1884
R6372 GND.n1265 GND.n1264 45.1884
R6373 GND.n1293 GND.n1292 45.1884
R6374 GND.n4487 GND.n4486 45.1884
R6375 GND.n1388 GND.n1387 45.1884
R6376 GND.n1803 GND.n1802 45.1884
R6377 GND.n2540 GND.n2539 45.1884
R6378 GND.n2562 GND.n2561 45.1884
R6379 GND.n542 GND.n541 45.1884
R6380 GND.n5797 GND.n5796 45.1884
R6381 GND.n576 GND.n575 45.1884
R6382 GND.n1728 GND.n1727 45.1884
R6383 GND.n1760 GND.n1759 45.1884
R6384 GND.n4010 GND.n4009 45.1884
R6385 GND.n3831 GND.n2890 44.3322
R6386 GND.n3192 GND.n3191 44.3189
R6387 GND.n2338 GND.n2337 42.2793
R6388 GND.n4741 GND.n1293 42.2793
R6389 GND.n4488 GND.n4487 42.2793
R6390 GND.n4655 GND.n1388 42.2793
R6391 GND.n1804 GND.n1803 42.2793
R6392 GND.n2563 GND.n2562 42.2793
R6393 GND.n5761 GND.n542 42.2793
R6394 GND.n5798 GND.n5797 42.2793
R6395 GND.n5727 GND.n576 42.2793
R6396 GND.n1729 GND.n1728 42.2793
R6397 GND.n1761 GND.n1760 42.2793
R6398 GND.n4011 GND.n4010 42.2793
R6399 GND.n3190 GND.n3189 41.6274
R6400 GND.n2885 GND.n2884 41.6274
R6401 GND.n3199 GND.n3198 40.8975
R6402 GND.n2888 GND.n2887 40.8975
R6403 GND.n4771 GND.n1265 36.9518
R6404 GND.n4451 GND.n2540 36.9518
R6405 GND.n3198 GND.n3197 35.055
R6406 GND.n3193 GND.n3192 35.055
R6407 GND.n2877 GND.n2876 35.055
R6408 GND.n2887 GND.n2873 35.055
R6409 GND.n2970 GND.n2967 33.8737
R6410 GND.n3241 GND.n3238 33.8737
R6411 GND.n1919 GND.n1690 33.3036
R6412 GND.n1940 GND.n1690 33.3036
R6413 GND.n1948 GND.n1670 33.3036
R6414 GND.n1956 GND.n1670 33.3036
R6415 GND.n1956 GND.n1659 33.3036
R6416 GND.n1977 GND.n1659 33.3036
R6417 GND.n1977 GND.n1651 33.3036
R6418 GND.n1986 GND.n1651 33.3036
R6419 GND.n1295 GND.n1238 33.3036
R6420 GND.n4710 GND.n1306 33.3036
R6421 GND.n4704 GND.n1306 33.3036
R6422 GND.n3400 GND.n1327 33.3036
R6423 GND.n3964 GND.n2429 33.3036
R6424 GND.n4023 GND.n4022 33.3036
R6425 GND.n4023 GND.n2484 33.3036
R6426 GND.n2566 GND.n2516 33.3036
R6427 GND.n5857 GND.n431 33.3036
R6428 GND.n5857 GND.n434 33.3036
R6429 GND.n5851 GND.n434 33.3036
R6430 GND.n5851 GND.n444 33.3036
R6431 GND.n5845 GND.n444 33.3036
R6432 GND.n5845 GND.n453 33.3036
R6433 GND.n5839 GND.n463 33.3036
R6434 GND.n5833 GND.n463 33.3036
R6435 GND.n4885 GND.n4884 26.6429
R6436 GND.n1646 GND.n1118 26.6429
R6437 GND.n4878 GND.n1128 26.6429
R6438 GND.n1996 GND.n1131 26.6429
R6439 GND.n1995 GND.n1638 26.6429
R6440 GND.n2006 GND.n2005 26.6429
R6441 GND.n2021 GND.n1615 26.6429
R6442 GND.n2018 GND.n1617 26.6429
R6443 GND.n1606 GND.n1599 26.6429
R6444 GND.n2044 GND.n2043 26.6429
R6445 GND.n2058 GND.n1589 26.6429
R6446 GND.n2054 GND.n1591 26.6429
R6447 GND.n1581 GND.n1518 26.6429
R6448 GND.n2135 GND.n2134 26.6429
R6449 GND.n1574 GND.n1520 26.6429
R6450 GND.n2127 GND.n1528 26.6429
R6451 GND.n2124 GND.n1534 26.6429
R6452 GND.n2123 GND.n1536 26.6429
R6453 GND.n2118 GND.n2117 26.6429
R6454 GND.n1571 GND.n1543 26.6429
R6455 GND.n2107 GND.n1552 26.6429
R6456 GND.n2106 GND.n1557 26.6429
R6457 GND.n2101 GND.n2100 26.6429
R6458 GND.n2196 GND.n1502 26.6429
R6459 GND.n2198 GND.n1500 26.6429
R6460 GND.n2212 GND.n1488 26.6429
R6461 GND.n1493 GND.n1490 26.6429
R6462 GND.n2221 GND.n1481 26.6429
R6463 GND.n2227 GND.n1476 26.6429
R6464 GND.n2224 GND.n1478 26.6429
R6465 GND.n2237 GND.n1467 26.6429
R6466 GND.n2151 GND.n1468 26.6429
R6467 GND.n2251 GND.n1455 26.6429
R6468 GND.n2248 GND.n1458 26.6429
R6469 GND.n2261 GND.n1445 26.6429
R6470 GND.n2170 GND.n1446 26.6429
R6471 GND.n2278 GND.n1434 26.6429
R6472 GND.n1436 GND.n1428 26.6429
R6473 GND.n2287 GND.n2286 26.6429
R6474 GND.n2315 GND.n1414 26.6429
R6475 GND.n2318 GND.n1410 26.6429
R6476 GND.n2307 GND.n1412 26.6429
R6477 GND.n2329 GND.n1402 26.6429
R6478 GND.n4800 GND.n1236 26.6429
R6479 GND.n4407 GND.n2568 26.6429
R6480 GND.n3988 GND.n2576 26.6429
R6481 GND.n4108 GND.n2590 26.6429
R6482 GND.n4393 GND.n2593 26.6429
R6483 GND.n4116 GND.n2603 26.6429
R6484 GND.n4387 GND.n2606 26.6429
R6485 GND.n4123 GND.n2614 26.6429
R6486 GND.n4381 GND.n2617 26.6429
R6487 GND.n4375 GND.n2627 26.6429
R6488 GND.n4138 GND.n2635 26.6429
R6489 GND.n4369 GND.n2638 26.6429
R6490 GND.n4146 GND.n2645 26.6429
R6491 GND.n4153 GND.n2655 26.6429
R6492 GND.n4357 GND.n2658 26.6429
R6493 GND.n4161 GND.n2665 26.6429
R6494 GND.n4351 GND.n2668 26.6429
R6495 GND.n4168 GND.n2676 26.6429
R6496 GND.n4345 GND.n2679 26.6429
R6497 GND.n4176 GND.n2686 26.6429
R6498 GND.n4339 GND.n2689 26.6429
R6499 GND.n4333 GND.n2700 26.6429
R6500 GND.n4201 GND.n2707 26.6429
R6501 GND.n4327 GND.n2710 26.6429
R6502 GND.n4323 GND.n4322 26.6429
R6503 GND.n4315 GND.n2724 26.6429
R6504 GND.n4314 GND.n320 26.6429
R6505 GND.n5918 GND.n322 26.6429
R6506 GND.n4308 GND.n4307 26.6429
R6507 GND.n2754 GND.n2751 26.6429
R6508 GND.n4222 GND.n339 26.6429
R6509 GND.n5911 GND.n342 26.6429
R6510 GND.n4231 GND.n351 26.6429
R6511 GND.n4269 GND.n360 26.6429
R6512 GND.n5899 GND.n363 26.6429
R6513 GND.n4263 GND.n370 26.6429
R6514 GND.n5893 GND.n373 26.6429
R6515 GND.n5887 GND.n384 26.6429
R6516 GND.n4251 GND.n391 26.6429
R6517 GND.n5881 GND.n394 26.6429
R6518 GND.n5669 GND.n5668 26.6429
R6519 GND.n5875 GND.n404 26.6429
R6520 GND.n5699 GND.n411 26.6429
R6521 GND.n5869 GND.n414 26.6429
R6522 GND.n5693 GND.n422 26.6429
R6523 GND.n3221 GND.n3220 25.7944
R6524 GND.n2909 GND.n2908 25.7944
R6525 GND.n3217 GND.n3216 25.7944
R6526 GND.n3833 GND.n3832 25.7944
R6527 GND.n1940 GND.t25 22.9796
R6528 GND.n2326 GND.t12 22.9796
R6529 GND.n4399 GND.t1 22.9796
R6530 GND.n5839 GND.t39 22.9796
R6531 GND.n2017 GND.t162 21.6475
R6532 GND.t115 GND.n381 21.6475
R6533 GND.n3359 GND.n3358 21.0737
R6534 GND.n3831 GND.n3830 21.0737
R6535 GND.n1570 GND.t143 20.9814
R6536 GND.n2721 GND.t129 20.9814
R6537 GND.n4737 GND.n1295 20.6484
R6538 GND.n4483 GND.n2516 20.6484
R6539 GND.n2152 GND.t154 20.3154
R6540 GND.n2769 GND.t138 20.3154
R6541 GND.n3186 GND.t85 19.8005
R6542 GND.n3186 GND.t17 19.8005
R6543 GND.n3187 GND.t65 19.8005
R6544 GND.n3187 GND.t47 19.8005
R6545 GND.n2881 GND.t50 19.8005
R6546 GND.n2881 GND.t68 19.8005
R6547 GND.n2882 GND.t23 19.8005
R6548 GND.n2882 GND.t6 19.8005
R6549 GND.n3183 GND.n3182 19.5087
R6550 GND.n3196 GND.n3183 19.5087
R6551 GND.n3194 GND.n3185 19.5087
R6552 GND.n2886 GND.n2880 19.5087
R6553 GND.n4644 GND.n4643 19.3944
R6554 GND.n4643 GND.n4642 19.3944
R6555 GND.n4642 GND.n2343 19.3944
R6556 GND.n4700 GND.n4699 19.3944
R6557 GND.n4699 GND.n1332 19.3944
R6558 GND.n4692 GND.n1332 19.3944
R6559 GND.n4692 GND.n4691 19.3944
R6560 GND.n4691 GND.n1344 19.3944
R6561 GND.n4684 GND.n1344 19.3944
R6562 GND.n4684 GND.n4683 19.3944
R6563 GND.n4683 GND.n1352 19.3944
R6564 GND.n4676 GND.n1352 19.3944
R6565 GND.n4676 GND.n4675 19.3944
R6566 GND.n4675 GND.n1364 19.3944
R6567 GND.n4668 GND.n1364 19.3944
R6568 GND.n4668 GND.n4667 19.3944
R6569 GND.n4667 GND.n1372 19.3944
R6570 GND.n4660 GND.n1372 19.3944
R6571 GND.n4660 GND.n4659 19.3944
R6572 GND.n4659 GND.n1384 19.3944
R6573 GND.n1393 GND.n1384 19.3944
R6574 GND.n4650 GND.n1393 19.3944
R6575 GND.n4650 GND.n4649 19.3944
R6576 GND.n4649 GND.n4648 19.3944
R6577 GND.n4648 GND.n1398 19.3944
R6578 GND.n4638 GND.n4637 19.3944
R6579 GND.n4637 GND.n4636 19.3944
R6580 GND.n4636 GND.n2349 19.3944
R6581 GND.n4632 GND.n2349 19.3944
R6582 GND.n4632 GND.n4631 19.3944
R6583 GND.n4631 GND.n4630 19.3944
R6584 GND.n4630 GND.n2354 19.3944
R6585 GND.n4626 GND.n2354 19.3944
R6586 GND.n4626 GND.n4625 19.3944
R6587 GND.n4625 GND.n4624 19.3944
R6588 GND.n4624 GND.n2359 19.3944
R6589 GND.n4620 GND.n2359 19.3944
R6590 GND.n4620 GND.n4619 19.3944
R6591 GND.n4619 GND.n4618 19.3944
R6592 GND.n4618 GND.n2364 19.3944
R6593 GND.n4614 GND.n2364 19.3944
R6594 GND.n4614 GND.n4613 19.3944
R6595 GND.n4613 GND.n4612 19.3944
R6596 GND.n4612 GND.n2369 19.3944
R6597 GND.n4608 GND.n2369 19.3944
R6598 GND.n4608 GND.n4607 19.3944
R6599 GND.n4607 GND.n4606 19.3944
R6600 GND.n4606 GND.n2374 19.3944
R6601 GND.n4602 GND.n2374 19.3944
R6602 GND.n4602 GND.n4601 19.3944
R6603 GND.n4601 GND.n4600 19.3944
R6604 GND.n4600 GND.n2379 19.3944
R6605 GND.n4596 GND.n2379 19.3944
R6606 GND.n4596 GND.n4595 19.3944
R6607 GND.n4595 GND.n4594 19.3944
R6608 GND.n4594 GND.n2384 19.3944
R6609 GND.n4590 GND.n2384 19.3944
R6610 GND.n4590 GND.n4589 19.3944
R6611 GND.n4589 GND.n4588 19.3944
R6612 GND.n4588 GND.n2389 19.3944
R6613 GND.n4584 GND.n2389 19.3944
R6614 GND.n4584 GND.n4583 19.3944
R6615 GND.n4583 GND.n4582 19.3944
R6616 GND.n4582 GND.n2394 19.3944
R6617 GND.n4578 GND.n2394 19.3944
R6618 GND.n4578 GND.n4577 19.3944
R6619 GND.n4577 GND.n4576 19.3944
R6620 GND.n4576 GND.n2399 19.3944
R6621 GND.n4572 GND.n2399 19.3944
R6622 GND.n4572 GND.n4571 19.3944
R6623 GND.n4571 GND.n4570 19.3944
R6624 GND.n4570 GND.n2404 19.3944
R6625 GND.n4566 GND.n2404 19.3944
R6626 GND.n4566 GND.n4565 19.3944
R6627 GND.n4565 GND.n4564 19.3944
R6628 GND.n4564 GND.n2409 19.3944
R6629 GND.n4560 GND.n2409 19.3944
R6630 GND.n4560 GND.n4559 19.3944
R6631 GND.n4559 GND.n4558 19.3944
R6632 GND.n4558 GND.n2414 19.3944
R6633 GND.n4554 GND.n2414 19.3944
R6634 GND.n4554 GND.n4553 19.3944
R6635 GND.n4553 GND.n4552 19.3944
R6636 GND.n4552 GND.n2419 19.3944
R6637 GND.n4548 GND.n2419 19.3944
R6638 GND.n4548 GND.n4547 19.3944
R6639 GND.n4547 GND.n4546 19.3944
R6640 GND.n4546 GND.n2424 19.3944
R6641 GND.n4542 GND.n2424 19.3944
R6642 GND.n4542 GND.n4541 19.3944
R6643 GND.n1766 GND.n1688 19.3944
R6644 GND.n1942 GND.n1688 19.3944
R6645 GND.n1944 GND.n1942 19.3944
R6646 GND.n1944 GND.n1943 19.3944
R6647 GND.n1943 GND.n1668 19.3944
R6648 GND.n1959 GND.n1668 19.3944
R6649 GND.n1973 GND.n1959 19.3944
R6650 GND.n1973 GND.n1972 19.3944
R6651 GND.n1972 GND.n1971 19.3944
R6652 GND.n1971 GND.n1962 19.3944
R6653 GND.n1967 GND.n1962 19.3944
R6654 GND.n1967 GND.n1138 19.3944
R6655 GND.n4874 GND.n1138 19.3944
R6656 GND.n4874 GND.n4873 19.3944
R6657 GND.n4873 GND.n4872 19.3944
R6658 GND.n4872 GND.n1141 19.3944
R6659 GND.n4868 GND.n1141 19.3944
R6660 GND.n4868 GND.n4867 19.3944
R6661 GND.n4867 GND.n4866 19.3944
R6662 GND.n4866 GND.n1149 19.3944
R6663 GND.n4862 GND.n1149 19.3944
R6664 GND.n4862 GND.n4861 19.3944
R6665 GND.n4861 GND.n4860 19.3944
R6666 GND.n4860 GND.n1157 19.3944
R6667 GND.n4856 GND.n1157 19.3944
R6668 GND.n4856 GND.n4855 19.3944
R6669 GND.n4855 GND.n4854 19.3944
R6670 GND.n4854 GND.n1165 19.3944
R6671 GND.n4850 GND.n1165 19.3944
R6672 GND.n4850 GND.n4849 19.3944
R6673 GND.n4849 GND.n4848 19.3944
R6674 GND.n4848 GND.n1173 19.3944
R6675 GND.n4844 GND.n1173 19.3944
R6676 GND.n4844 GND.n4843 19.3944
R6677 GND.n4843 GND.n4842 19.3944
R6678 GND.n4842 GND.n1181 19.3944
R6679 GND.n4838 GND.n1181 19.3944
R6680 GND.n4838 GND.n4837 19.3944
R6681 GND.n4837 GND.n4836 19.3944
R6682 GND.n4836 GND.n1189 19.3944
R6683 GND.n4832 GND.n1189 19.3944
R6684 GND.n4832 GND.n4831 19.3944
R6685 GND.n4831 GND.n4830 19.3944
R6686 GND.n4830 GND.n1197 19.3944
R6687 GND.n4826 GND.n1197 19.3944
R6688 GND.n4826 GND.n4825 19.3944
R6689 GND.n4825 GND.n4824 19.3944
R6690 GND.n4824 GND.n1205 19.3944
R6691 GND.n4820 GND.n1205 19.3944
R6692 GND.n4820 GND.n4819 19.3944
R6693 GND.n4819 GND.n4818 19.3944
R6694 GND.n4818 GND.n1213 19.3944
R6695 GND.n4814 GND.n1213 19.3944
R6696 GND.n4814 GND.n4813 19.3944
R6697 GND.n4813 GND.n4812 19.3944
R6698 GND.n4812 GND.n1221 19.3944
R6699 GND.n4808 GND.n1221 19.3944
R6700 GND.n4808 GND.n4807 19.3944
R6701 GND.n4807 GND.n4806 19.3944
R6702 GND.n4806 GND.n1229 19.3944
R6703 GND.n4802 GND.n1229 19.3944
R6704 GND.n4795 GND.n4794 19.3944
R6705 GND.n4794 GND.n4793 19.3944
R6706 GND.n4793 GND.n1247 19.3944
R6707 GND.n4789 GND.n1247 19.3944
R6708 GND.n4789 GND.n4788 19.3944
R6709 GND.n4788 GND.n4787 19.3944
R6710 GND.n4787 GND.n1252 19.3944
R6711 GND.n4783 GND.n1252 19.3944
R6712 GND.n4783 GND.n4782 19.3944
R6713 GND.n4782 GND.n4781 19.3944
R6714 GND.n4781 GND.n1257 19.3944
R6715 GND.n4777 GND.n1257 19.3944
R6716 GND.n4777 GND.n4776 19.3944
R6717 GND.n4776 GND.n4775 19.3944
R6718 GND.n4775 GND.n1262 19.3944
R6719 GND.n4770 GND.n4769 19.3944
R6720 GND.n4769 GND.n1270 19.3944
R6721 GND.n4765 GND.n1270 19.3944
R6722 GND.n4765 GND.n4764 19.3944
R6723 GND.n4764 GND.n4763 19.3944
R6724 GND.n4763 GND.n1275 19.3944
R6725 GND.n4759 GND.n1275 19.3944
R6726 GND.n4759 GND.n4758 19.3944
R6727 GND.n4758 GND.n4757 19.3944
R6728 GND.n4757 GND.n1280 19.3944
R6729 GND.n4753 GND.n1280 19.3944
R6730 GND.n4753 GND.n4752 19.3944
R6731 GND.n4752 GND.n4751 19.3944
R6732 GND.n4751 GND.n1285 19.3944
R6733 GND.n4747 GND.n1285 19.3944
R6734 GND.n4747 GND.n4746 19.3944
R6735 GND.n4746 GND.n4745 19.3944
R6736 GND.n4745 GND.n1290 19.3944
R6737 GND.n4529 GND.n2439 19.3944
R6738 GND.n4529 GND.n4528 19.3944
R6739 GND.n4528 GND.n2442 19.3944
R6740 GND.n4521 GND.n2442 19.3944
R6741 GND.n4521 GND.n4520 19.3944
R6742 GND.n4520 GND.n2450 19.3944
R6743 GND.n4513 GND.n2450 19.3944
R6744 GND.n4513 GND.n4512 19.3944
R6745 GND.n4512 GND.n2458 19.3944
R6746 GND.n4505 GND.n2458 19.3944
R6747 GND.n4505 GND.n4504 19.3944
R6748 GND.n4504 GND.n2466 19.3944
R6749 GND.n4497 GND.n2466 19.3944
R6750 GND.n4497 GND.n4496 19.3944
R6751 GND.n4496 GND.n2474 19.3944
R6752 GND.n4489 GND.n2474 19.3944
R6753 GND.n1921 GND.n1692 19.3944
R6754 GND.n1938 GND.n1692 19.3944
R6755 GND.n1938 GND.n1693 19.3944
R6756 GND.n1934 GND.n1693 19.3944
R6757 GND.n1934 GND.n1933 19.3944
R6758 GND.n1933 GND.n1932 19.3944
R6759 GND.n1932 GND.n1927 19.3944
R6760 GND.n1928 GND.n1927 19.3944
R6761 GND.n1928 GND.n1649 19.3944
R6762 GND.n1989 GND.n1649 19.3944
R6763 GND.n1989 GND.n1644 19.3944
R6764 GND.n1993 GND.n1644 19.3944
R6765 GND.n1994 GND.n1993 19.3944
R6766 GND.n1998 GND.n1994 19.3944
R6767 GND.n1998 GND.n1641 19.3944
R6768 GND.n2003 GND.n1641 19.3944
R6769 GND.n2003 GND.n1642 19.3944
R6770 GND.n1642 GND.n1604 19.3944
R6771 GND.n2033 GND.n1604 19.3944
R6772 GND.n2033 GND.n1601 19.3944
R6773 GND.n2041 GND.n1601 19.3944
R6774 GND.n2041 GND.n1602 19.3944
R6775 GND.n2037 GND.n1602 19.3944
R6776 GND.n2037 GND.n1578 19.3944
R6777 GND.n2070 GND.n1578 19.3944
R6778 GND.n2071 GND.n2070 19.3944
R6779 GND.n2071 GND.n1576 19.3944
R6780 GND.n2075 GND.n1576 19.3944
R6781 GND.n2076 GND.n2075 19.3944
R6782 GND.n2078 GND.n2076 19.3944
R6783 GND.n2078 GND.n1565 19.3944
R6784 GND.n2083 GND.n1565 19.3944
R6785 GND.n2084 GND.n2083 19.3944
R6786 GND.n2085 GND.n2084 19.3944
R6787 GND.n2085 GND.n1562 19.3944
R6788 GND.n2092 GND.n1562 19.3944
R6789 GND.n2092 GND.n1563 19.3944
R6790 GND.n2088 GND.n1563 19.3944
R6791 GND.n2088 GND.n1486 19.3944
R6792 GND.n2214 GND.n1486 19.3944
R6793 GND.n2214 GND.n1483 19.3944
R6794 GND.n2219 GND.n1483 19.3944
R6795 GND.n2219 GND.n1484 19.3944
R6796 GND.n1484 GND.n1465 19.3944
R6797 GND.n2239 GND.n1465 19.3944
R6798 GND.n2239 GND.n1462 19.3944
R6799 GND.n2244 GND.n1462 19.3944
R6800 GND.n2244 GND.n1463 19.3944
R6801 GND.n1463 GND.n1443 19.3944
R6802 GND.n2263 GND.n1443 19.3944
R6803 GND.n2263 GND.n1440 19.3944
R6804 GND.n2271 GND.n1440 19.3944
R6805 GND.n2271 GND.n1441 19.3944
R6806 GND.n2267 GND.n1441 19.3944
R6807 GND.n2267 GND.n1417 19.3944
R6808 GND.n2313 GND.n1417 19.3944
R6809 GND.n2313 GND.n1418 19.3944
R6810 GND.n2309 GND.n1418 19.3944
R6811 GND.n2309 GND.n1400 19.3944
R6812 GND.n2331 GND.n1400 19.3944
R6813 GND.n2332 GND.n2331 19.3944
R6814 GND.n4696 GND.n1335 19.3944
R6815 GND.n4696 GND.n4695 19.3944
R6816 GND.n4695 GND.n1339 19.3944
R6817 GND.n4688 GND.n1339 19.3944
R6818 GND.n4688 GND.n4687 19.3944
R6819 GND.n4687 GND.n1348 19.3944
R6820 GND.n4680 GND.n1348 19.3944
R6821 GND.n4680 GND.n4679 19.3944
R6822 GND.n4679 GND.n1358 19.3944
R6823 GND.n4672 GND.n1358 19.3944
R6824 GND.n4672 GND.n4671 19.3944
R6825 GND.n4671 GND.n1368 19.3944
R6826 GND.n4664 GND.n1368 19.3944
R6827 GND.n4664 GND.n4663 19.3944
R6828 GND.n4663 GND.n1378 19.3944
R6829 GND.n4656 GND.n1378 19.3944
R6830 GND.n1832 GND.n1769 19.3944
R6831 GND.n1827 GND.n1769 19.3944
R6832 GND.n1827 GND.n1771 19.3944
R6833 GND.n1823 GND.n1771 19.3944
R6834 GND.n1823 GND.n1822 19.3944
R6835 GND.n1822 GND.n1821 19.3944
R6836 GND.n1821 GND.n1778 19.3944
R6837 GND.n1817 GND.n1778 19.3944
R6838 GND.n1817 GND.n1816 19.3944
R6839 GND.n1816 GND.n1815 19.3944
R6840 GND.n1815 GND.n1786 19.3944
R6841 GND.n1811 GND.n1786 19.3944
R6842 GND.n1811 GND.n1810 19.3944
R6843 GND.n1810 GND.n1809 19.3944
R6844 GND.n1809 GND.n1794 19.3944
R6845 GND.n1805 GND.n1794 19.3944
R6846 GND.n1764 GND.n1762 19.3944
R6847 GND.n1764 GND.n1682 19.3944
R6848 GND.n1946 GND.n1682 19.3944
R6849 GND.n1946 GND.n1683 19.3944
R6850 GND.n1685 GND.n1683 19.3944
R6851 GND.n1685 GND.n1664 19.3944
R6852 GND.n1975 GND.n1664 19.3944
R6853 GND.n1975 GND.n1665 19.3944
R6854 GND.n1963 GND.n1665 19.3944
R6855 GND.n1965 GND.n1963 19.3944
R6856 GND.n1966 GND.n1965 19.3944
R6857 GND.n1966 GND.n1134 19.3944
R6858 GND.n4876 GND.n1134 19.3944
R6859 GND.n4876 GND.n1135 19.3944
R6860 GND.n1142 GND.n1135 19.3944
R6861 GND.n1143 GND.n1142 19.3944
R6862 GND.n1144 GND.n1143 19.3944
R6863 GND.n1619 GND.n1144 19.3944
R6864 GND.n1619 GND.n1150 19.3944
R6865 GND.n1151 GND.n1150 19.3944
R6866 GND.n1152 GND.n1151 19.3944
R6867 GND.n2056 GND.n1152 19.3944
R6868 GND.n2056 GND.n1158 19.3944
R6869 GND.n1159 GND.n1158 19.3944
R6870 GND.n1160 GND.n1159 19.3944
R6871 GND.n1521 GND.n1160 19.3944
R6872 GND.n1521 GND.n1166 19.3944
R6873 GND.n1167 GND.n1166 19.3944
R6874 GND.n1168 GND.n1167 19.3944
R6875 GND.n1532 GND.n1168 19.3944
R6876 GND.n1532 GND.n1174 19.3944
R6877 GND.n1175 GND.n1174 19.3944
R6878 GND.n1176 GND.n1175 19.3944
R6879 GND.n1555 GND.n1176 19.3944
R6880 GND.n1555 GND.n1182 19.3944
R6881 GND.n1183 GND.n1182 19.3944
R6882 GND.n1184 GND.n1183 19.3944
R6883 GND.n2200 GND.n1184 19.3944
R6884 GND.n2200 GND.n1190 19.3944
R6885 GND.n1191 GND.n1190 19.3944
R6886 GND.n1192 GND.n1191 19.3944
R6887 GND.n1480 GND.n1192 19.3944
R6888 GND.n1480 GND.n1198 19.3944
R6889 GND.n1199 GND.n1198 19.3944
R6890 GND.n1200 GND.n1199 19.3944
R6891 GND.n1459 GND.n1200 19.3944
R6892 GND.n1459 GND.n1206 19.3944
R6893 GND.n1207 GND.n1206 19.3944
R6894 GND.n1208 GND.n1207 19.3944
R6895 GND.n1447 GND.n1208 19.3944
R6896 GND.n1447 GND.n1214 19.3944
R6897 GND.n1215 GND.n1214 19.3944
R6898 GND.n1216 GND.n1215 19.3944
R6899 GND.n2275 GND.n1216 19.3944
R6900 GND.n2275 GND.n1222 19.3944
R6901 GND.n1223 GND.n1222 19.3944
R6902 GND.n1224 GND.n1223 19.3944
R6903 GND.n1403 GND.n1224 19.3944
R6904 GND.n1403 GND.n1230 19.3944
R6905 GND.n1231 GND.n1230 19.3944
R6906 GND.n1232 GND.n1231 19.3944
R6907 GND.n5484 GND.n700 19.3944
R6908 GND.n5488 GND.n700 19.3944
R6909 GND.n5488 GND.n696 19.3944
R6910 GND.n5494 GND.n696 19.3944
R6911 GND.n5494 GND.n694 19.3944
R6912 GND.n5498 GND.n694 19.3944
R6913 GND.n5498 GND.n690 19.3944
R6914 GND.n5504 GND.n690 19.3944
R6915 GND.n5504 GND.n688 19.3944
R6916 GND.n5508 GND.n688 19.3944
R6917 GND.n5508 GND.n684 19.3944
R6918 GND.n5514 GND.n684 19.3944
R6919 GND.n5514 GND.n682 19.3944
R6920 GND.n5518 GND.n682 19.3944
R6921 GND.n5518 GND.n678 19.3944
R6922 GND.n5524 GND.n678 19.3944
R6923 GND.n5524 GND.n676 19.3944
R6924 GND.n5528 GND.n676 19.3944
R6925 GND.n5528 GND.n672 19.3944
R6926 GND.n5534 GND.n672 19.3944
R6927 GND.n5534 GND.n670 19.3944
R6928 GND.n5538 GND.n670 19.3944
R6929 GND.n5538 GND.n666 19.3944
R6930 GND.n5544 GND.n666 19.3944
R6931 GND.n5544 GND.n664 19.3944
R6932 GND.n5548 GND.n664 19.3944
R6933 GND.n5548 GND.n660 19.3944
R6934 GND.n5554 GND.n660 19.3944
R6935 GND.n5554 GND.n658 19.3944
R6936 GND.n5558 GND.n658 19.3944
R6937 GND.n5558 GND.n654 19.3944
R6938 GND.n5564 GND.n654 19.3944
R6939 GND.n5564 GND.n652 19.3944
R6940 GND.n5568 GND.n652 19.3944
R6941 GND.n5568 GND.n648 19.3944
R6942 GND.n5574 GND.n648 19.3944
R6943 GND.n5574 GND.n646 19.3944
R6944 GND.n5578 GND.n646 19.3944
R6945 GND.n5578 GND.n642 19.3944
R6946 GND.n5584 GND.n642 19.3944
R6947 GND.n5584 GND.n640 19.3944
R6948 GND.n5588 GND.n640 19.3944
R6949 GND.n5588 GND.n636 19.3944
R6950 GND.n5594 GND.n636 19.3944
R6951 GND.n5594 GND.n634 19.3944
R6952 GND.n5598 GND.n634 19.3944
R6953 GND.n5598 GND.n630 19.3944
R6954 GND.n5604 GND.n630 19.3944
R6955 GND.n5604 GND.n628 19.3944
R6956 GND.n5608 GND.n628 19.3944
R6957 GND.n5608 GND.n624 19.3944
R6958 GND.n5614 GND.n624 19.3944
R6959 GND.n5614 GND.n622 19.3944
R6960 GND.n5618 GND.n622 19.3944
R6961 GND.n5618 GND.n618 19.3944
R6962 GND.n5624 GND.n618 19.3944
R6963 GND.n5624 GND.n616 19.3944
R6964 GND.n5628 GND.n616 19.3944
R6965 GND.n5628 GND.n612 19.3944
R6966 GND.n5634 GND.n612 19.3944
R6967 GND.n5634 GND.n610 19.3944
R6968 GND.n5638 GND.n610 19.3944
R6969 GND.n5638 GND.n606 19.3944
R6970 GND.n5644 GND.n606 19.3944
R6971 GND.n5644 GND.n604 19.3944
R6972 GND.n5649 GND.n604 19.3944
R6973 GND.n5649 GND.n600 19.3944
R6974 GND.n5656 GND.n600 19.3944
R6975 GND.n5657 GND.n5656 19.3944
R6976 GND.n5033 GND.n971 19.3944
R6977 GND.n5033 GND.n969 19.3944
R6978 GND.n5037 GND.n969 19.3944
R6979 GND.n5037 GND.n965 19.3944
R6980 GND.n5043 GND.n965 19.3944
R6981 GND.n5043 GND.n963 19.3944
R6982 GND.n5047 GND.n963 19.3944
R6983 GND.n5047 GND.n959 19.3944
R6984 GND.n5053 GND.n959 19.3944
R6985 GND.n5053 GND.n957 19.3944
R6986 GND.n5057 GND.n957 19.3944
R6987 GND.n5057 GND.n953 19.3944
R6988 GND.n5063 GND.n953 19.3944
R6989 GND.n5063 GND.n951 19.3944
R6990 GND.n5067 GND.n951 19.3944
R6991 GND.n5067 GND.n947 19.3944
R6992 GND.n5073 GND.n947 19.3944
R6993 GND.n5073 GND.n945 19.3944
R6994 GND.n5077 GND.n945 19.3944
R6995 GND.n5077 GND.n941 19.3944
R6996 GND.n5083 GND.n941 19.3944
R6997 GND.n5083 GND.n939 19.3944
R6998 GND.n5087 GND.n939 19.3944
R6999 GND.n5087 GND.n935 19.3944
R7000 GND.n5093 GND.n935 19.3944
R7001 GND.n5093 GND.n933 19.3944
R7002 GND.n5097 GND.n933 19.3944
R7003 GND.n5097 GND.n929 19.3944
R7004 GND.n5103 GND.n929 19.3944
R7005 GND.n5103 GND.n927 19.3944
R7006 GND.n5107 GND.n927 19.3944
R7007 GND.n5107 GND.n923 19.3944
R7008 GND.n5113 GND.n923 19.3944
R7009 GND.n5113 GND.n921 19.3944
R7010 GND.n5117 GND.n921 19.3944
R7011 GND.n5117 GND.n917 19.3944
R7012 GND.n5123 GND.n917 19.3944
R7013 GND.n5123 GND.n915 19.3944
R7014 GND.n5127 GND.n915 19.3944
R7015 GND.n5127 GND.n911 19.3944
R7016 GND.n5133 GND.n911 19.3944
R7017 GND.n5133 GND.n909 19.3944
R7018 GND.n5137 GND.n909 19.3944
R7019 GND.n5137 GND.n905 19.3944
R7020 GND.n5143 GND.n905 19.3944
R7021 GND.n5143 GND.n903 19.3944
R7022 GND.n5147 GND.n903 19.3944
R7023 GND.n5147 GND.n899 19.3944
R7024 GND.n5153 GND.n899 19.3944
R7025 GND.n5153 GND.n897 19.3944
R7026 GND.n5157 GND.n897 19.3944
R7027 GND.n5157 GND.n893 19.3944
R7028 GND.n5163 GND.n893 19.3944
R7029 GND.n5163 GND.n891 19.3944
R7030 GND.n5167 GND.n891 19.3944
R7031 GND.n5167 GND.n887 19.3944
R7032 GND.n5173 GND.n887 19.3944
R7033 GND.n5173 GND.n885 19.3944
R7034 GND.n5177 GND.n885 19.3944
R7035 GND.n5177 GND.n881 19.3944
R7036 GND.n5183 GND.n881 19.3944
R7037 GND.n5183 GND.n879 19.3944
R7038 GND.n5187 GND.n879 19.3944
R7039 GND.n5187 GND.n875 19.3944
R7040 GND.n5193 GND.n875 19.3944
R7041 GND.n5193 GND.n873 19.3944
R7042 GND.n5197 GND.n873 19.3944
R7043 GND.n5197 GND.n869 19.3944
R7044 GND.n5203 GND.n869 19.3944
R7045 GND.n5203 GND.n867 19.3944
R7046 GND.n5207 GND.n867 19.3944
R7047 GND.n5207 GND.n863 19.3944
R7048 GND.n5213 GND.n863 19.3944
R7049 GND.n5213 GND.n861 19.3944
R7050 GND.n5217 GND.n861 19.3944
R7051 GND.n5217 GND.n857 19.3944
R7052 GND.n5223 GND.n857 19.3944
R7053 GND.n5223 GND.n855 19.3944
R7054 GND.n5227 GND.n855 19.3944
R7055 GND.n5227 GND.n851 19.3944
R7056 GND.n5233 GND.n851 19.3944
R7057 GND.n5233 GND.n849 19.3944
R7058 GND.n5237 GND.n849 19.3944
R7059 GND.n5237 GND.n845 19.3944
R7060 GND.n5243 GND.n845 19.3944
R7061 GND.n5243 GND.n843 19.3944
R7062 GND.n5247 GND.n843 19.3944
R7063 GND.n5247 GND.n839 19.3944
R7064 GND.n5253 GND.n839 19.3944
R7065 GND.n5253 GND.n837 19.3944
R7066 GND.n5257 GND.n837 19.3944
R7067 GND.n5257 GND.n833 19.3944
R7068 GND.n5263 GND.n833 19.3944
R7069 GND.n5263 GND.n831 19.3944
R7070 GND.n5267 GND.n831 19.3944
R7071 GND.n5267 GND.n827 19.3944
R7072 GND.n5273 GND.n827 19.3944
R7073 GND.n5273 GND.n825 19.3944
R7074 GND.n5277 GND.n825 19.3944
R7075 GND.n5277 GND.n821 19.3944
R7076 GND.n5283 GND.n821 19.3944
R7077 GND.n5283 GND.n819 19.3944
R7078 GND.n5287 GND.n819 19.3944
R7079 GND.n5287 GND.n815 19.3944
R7080 GND.n5293 GND.n815 19.3944
R7081 GND.n5293 GND.n813 19.3944
R7082 GND.n5297 GND.n813 19.3944
R7083 GND.n5297 GND.n809 19.3944
R7084 GND.n5303 GND.n809 19.3944
R7085 GND.n5303 GND.n807 19.3944
R7086 GND.n5307 GND.n807 19.3944
R7087 GND.n5307 GND.n803 19.3944
R7088 GND.n5313 GND.n803 19.3944
R7089 GND.n5313 GND.n801 19.3944
R7090 GND.n5317 GND.n801 19.3944
R7091 GND.n5317 GND.n797 19.3944
R7092 GND.n5323 GND.n797 19.3944
R7093 GND.n5323 GND.n795 19.3944
R7094 GND.n5327 GND.n795 19.3944
R7095 GND.n5327 GND.n791 19.3944
R7096 GND.n5333 GND.n791 19.3944
R7097 GND.n5333 GND.n789 19.3944
R7098 GND.n5337 GND.n789 19.3944
R7099 GND.n5337 GND.n785 19.3944
R7100 GND.n5343 GND.n785 19.3944
R7101 GND.n5343 GND.n783 19.3944
R7102 GND.n5347 GND.n783 19.3944
R7103 GND.n5347 GND.n779 19.3944
R7104 GND.n5353 GND.n779 19.3944
R7105 GND.n5353 GND.n777 19.3944
R7106 GND.n5357 GND.n777 19.3944
R7107 GND.n5357 GND.n773 19.3944
R7108 GND.n5363 GND.n773 19.3944
R7109 GND.n5363 GND.n771 19.3944
R7110 GND.n5367 GND.n771 19.3944
R7111 GND.n5367 GND.n767 19.3944
R7112 GND.n5373 GND.n767 19.3944
R7113 GND.n5373 GND.n765 19.3944
R7114 GND.n5377 GND.n765 19.3944
R7115 GND.n5377 GND.n761 19.3944
R7116 GND.n5383 GND.n761 19.3944
R7117 GND.n5383 GND.n759 19.3944
R7118 GND.n5387 GND.n759 19.3944
R7119 GND.n5387 GND.n755 19.3944
R7120 GND.n5393 GND.n755 19.3944
R7121 GND.n5393 GND.n753 19.3944
R7122 GND.n5397 GND.n753 19.3944
R7123 GND.n5397 GND.n749 19.3944
R7124 GND.n5403 GND.n749 19.3944
R7125 GND.n5403 GND.n747 19.3944
R7126 GND.n5407 GND.n747 19.3944
R7127 GND.n5407 GND.n743 19.3944
R7128 GND.n5413 GND.n743 19.3944
R7129 GND.n5413 GND.n741 19.3944
R7130 GND.n5417 GND.n741 19.3944
R7131 GND.n5417 GND.n737 19.3944
R7132 GND.n5423 GND.n737 19.3944
R7133 GND.n5423 GND.n735 19.3944
R7134 GND.n5427 GND.n735 19.3944
R7135 GND.n5427 GND.n731 19.3944
R7136 GND.n5433 GND.n731 19.3944
R7137 GND.n5433 GND.n729 19.3944
R7138 GND.n5437 GND.n729 19.3944
R7139 GND.n5437 GND.n725 19.3944
R7140 GND.n5443 GND.n725 19.3944
R7141 GND.n5443 GND.n723 19.3944
R7142 GND.n5447 GND.n723 19.3944
R7143 GND.n5447 GND.n719 19.3944
R7144 GND.n5453 GND.n719 19.3944
R7145 GND.n5453 GND.n717 19.3944
R7146 GND.n5457 GND.n717 19.3944
R7147 GND.n5457 GND.n713 19.3944
R7148 GND.n5463 GND.n713 19.3944
R7149 GND.n5463 GND.n711 19.3944
R7150 GND.n5467 GND.n711 19.3944
R7151 GND.n5467 GND.n707 19.3944
R7152 GND.n5473 GND.n707 19.3944
R7153 GND.n5473 GND.n705 19.3944
R7154 GND.n5478 GND.n705 19.3944
R7155 GND.n5478 GND.n5477 19.3944
R7156 GND.n4480 GND.n4479 19.3944
R7157 GND.n4479 GND.n4478 19.3944
R7158 GND.n4478 GND.n4477 19.3944
R7159 GND.n4477 GND.n4475 19.3944
R7160 GND.n4475 GND.n4472 19.3944
R7161 GND.n4472 GND.n4471 19.3944
R7162 GND.n4471 GND.n4468 19.3944
R7163 GND.n4468 GND.n4467 19.3944
R7164 GND.n4467 GND.n4464 19.3944
R7165 GND.n4464 GND.n4463 19.3944
R7166 GND.n4463 GND.n4460 19.3944
R7167 GND.n4460 GND.n4459 19.3944
R7168 GND.n4459 GND.n4456 19.3944
R7169 GND.n4456 GND.n4455 19.3944
R7170 GND.n4455 GND.n4452 19.3944
R7171 GND.n4450 GND.n4447 19.3944
R7172 GND.n4447 GND.n4446 19.3944
R7173 GND.n4446 GND.n4443 19.3944
R7174 GND.n4443 GND.n4442 19.3944
R7175 GND.n4442 GND.n4439 19.3944
R7176 GND.n4439 GND.n4438 19.3944
R7177 GND.n4438 GND.n4435 19.3944
R7178 GND.n4435 GND.n4434 19.3944
R7179 GND.n4434 GND.n4431 19.3944
R7180 GND.n4431 GND.n4430 19.3944
R7181 GND.n4430 GND.n4427 19.3944
R7182 GND.n4427 GND.n4426 19.3944
R7183 GND.n4426 GND.n4423 19.3944
R7184 GND.n4423 GND.n4422 19.3944
R7185 GND.n4422 GND.n4419 19.3944
R7186 GND.n4419 GND.n4418 19.3944
R7187 GND.n4418 GND.n4415 19.3944
R7188 GND.n4415 GND.n4414 19.3944
R7189 GND.n4402 GND.n2565 19.3944
R7190 GND.n4402 GND.n4401 19.3944
R7191 GND.n4401 GND.n2574 19.3944
R7192 GND.n2778 GND.n2574 19.3944
R7193 GND.n4118 GND.n2778 19.3944
R7194 GND.n4119 GND.n4118 19.3944
R7195 GND.n4121 GND.n4119 19.3944
R7196 GND.n4121 GND.n2774 19.3944
R7197 GND.n4133 GND.n2774 19.3944
R7198 GND.n4134 GND.n4133 19.3944
R7199 GND.n4136 GND.n4134 19.3944
R7200 GND.n4136 GND.n2770 19.3944
R7201 GND.n4148 GND.n2770 19.3944
R7202 GND.n4149 GND.n4148 19.3944
R7203 GND.n4151 GND.n4149 19.3944
R7204 GND.n4151 GND.n2765 19.3944
R7205 GND.n4163 GND.n2765 19.3944
R7206 GND.n4164 GND.n4163 19.3944
R7207 GND.n4166 GND.n4164 19.3944
R7208 GND.n4166 GND.n2761 19.3944
R7209 GND.n4178 GND.n2761 19.3944
R7210 GND.n4179 GND.n4178 19.3944
R7211 GND.n4181 GND.n4179 19.3944
R7212 GND.n4181 GND.n2757 19.3944
R7213 GND.n4203 GND.n2757 19.3944
R7214 GND.n4204 GND.n4203 19.3944
R7215 GND.n4205 GND.n4204 19.3944
R7216 GND.n4205 GND.n2756 19.3944
R7217 GND.n4213 GND.n2756 19.3944
R7218 GND.n4214 GND.n4213 19.3944
R7219 GND.n4215 GND.n4214 19.3944
R7220 GND.n4216 GND.n4215 19.3944
R7221 GND.n4217 GND.n4216 19.3944
R7222 GND.n4220 GND.n4217 19.3944
R7223 GND.n4220 GND.n2746 19.3944
R7224 GND.n4233 GND.n2746 19.3944
R7225 GND.n4234 GND.n4233 19.3944
R7226 GND.n4236 GND.n4234 19.3944
R7227 GND.n4237 GND.n4236 19.3944
R7228 GND.n4261 GND.n4237 19.3944
R7229 GND.n4261 GND.n4260 19.3944
R7230 GND.n4260 GND.n4259 19.3944
R7231 GND.n4259 GND.n4239 19.3944
R7232 GND.n4249 GND.n4239 19.3944
R7233 GND.n4249 GND.n587 19.3944
R7234 GND.n5671 GND.n587 19.3944
R7235 GND.n5672 GND.n5671 19.3944
R7236 GND.n5697 GND.n5672 19.3944
R7237 GND.n5697 GND.n5696 19.3944
R7238 GND.n5696 GND.n5695 19.3944
R7239 GND.n5695 GND.n5691 19.3944
R7240 GND.n5691 GND.n5690 19.3944
R7241 GND.n5690 GND.n5688 19.3944
R7242 GND.n5688 GND.n5687 19.3944
R7243 GND.n5687 GND.n5685 19.3944
R7244 GND.n5685 GND.n5684 19.3944
R7245 GND.n5684 GND.n5682 19.3944
R7246 GND.n5682 GND.n5681 19.3944
R7247 GND.n5681 GND.n5679 19.3944
R7248 GND.n5679 GND.n5678 19.3944
R7249 GND.n5678 GND.n5676 19.3944
R7250 GND.n4405 GND.n4404 19.3944
R7251 GND.n4404 GND.n2572 19.3944
R7252 GND.n2596 GND.n2572 19.3944
R7253 GND.n4391 GND.n2596 19.3944
R7254 GND.n4391 GND.n4390 19.3944
R7255 GND.n4390 GND.n4389 19.3944
R7256 GND.n4389 GND.n2601 19.3944
R7257 GND.n4379 GND.n2601 19.3944
R7258 GND.n4379 GND.n4378 19.3944
R7259 GND.n4378 GND.n4377 19.3944
R7260 GND.n4377 GND.n2622 19.3944
R7261 GND.n4367 GND.n2622 19.3944
R7262 GND.n4367 GND.n4366 19.3944
R7263 GND.n4366 GND.n4365 19.3944
R7264 GND.n4365 GND.n2643 19.3944
R7265 GND.n4355 GND.n2643 19.3944
R7266 GND.n4355 GND.n4354 19.3944
R7267 GND.n4354 GND.n4353 19.3944
R7268 GND.n4353 GND.n2663 19.3944
R7269 GND.n4343 GND.n2663 19.3944
R7270 GND.n4343 GND.n4342 19.3944
R7271 GND.n4342 GND.n4341 19.3944
R7272 GND.n4341 GND.n2684 19.3944
R7273 GND.n4331 GND.n2684 19.3944
R7274 GND.n4331 GND.n4330 19.3944
R7275 GND.n4330 GND.n4329 19.3944
R7276 GND.n4329 GND.n2705 19.3944
R7277 GND.n4208 GND.n2705 19.3944
R7278 GND.n4208 GND.n2727 19.3944
R7279 GND.n4312 GND.n2727 19.3944
R7280 GND.n4312 GND.n4311 19.3944
R7281 GND.n4311 GND.n4310 19.3944
R7282 GND.n4310 GND.n2731 19.3944
R7283 GND.n2731 GND.n345 19.3944
R7284 GND.n5909 GND.n345 19.3944
R7285 GND.n5909 GND.n5908 19.3944
R7286 GND.n5908 GND.n5907 19.3944
R7287 GND.n5907 GND.n349 19.3944
R7288 GND.n5897 GND.n349 19.3944
R7289 GND.n5897 GND.n5896 19.3944
R7290 GND.n5896 GND.n5895 19.3944
R7291 GND.n5895 GND.n368 19.3944
R7292 GND.n5885 GND.n368 19.3944
R7293 GND.n5885 GND.n5884 19.3944
R7294 GND.n5884 GND.n5883 19.3944
R7295 GND.n5883 GND.n389 19.3944
R7296 GND.n5873 GND.n389 19.3944
R7297 GND.n5873 GND.n5872 19.3944
R7298 GND.n5872 GND.n5871 19.3944
R7299 GND.n5871 GND.n409 19.3944
R7300 GND.n5861 GND.n409 19.3944
R7301 GND.n5861 GND.n5860 19.3944
R7302 GND.n5860 GND.n5859 19.3944
R7303 GND.n5859 GND.n429 19.3944
R7304 GND.n5849 GND.n429 19.3944
R7305 GND.n5849 GND.n5848 19.3944
R7306 GND.n5848 GND.n5847 19.3944
R7307 GND.n5847 GND.n449 19.3944
R7308 GND.n5837 GND.n449 19.3944
R7309 GND.n5837 GND.n5836 19.3944
R7310 GND.n5836 GND.n5835 19.3944
R7311 GND.n5795 GND.n505 19.3944
R7312 GND.n5790 GND.n505 19.3944
R7313 GND.n5790 GND.n5789 19.3944
R7314 GND.n5789 GND.n5788 19.3944
R7315 GND.n5788 GND.n512 19.3944
R7316 GND.n5783 GND.n512 19.3944
R7317 GND.n5783 GND.n5782 19.3944
R7318 GND.n5782 GND.n5781 19.3944
R7319 GND.n5781 GND.n519 19.3944
R7320 GND.n5776 GND.n519 19.3944
R7321 GND.n5776 GND.n5775 19.3944
R7322 GND.n5775 GND.n5774 19.3944
R7323 GND.n5774 GND.n526 19.3944
R7324 GND.n5769 GND.n526 19.3944
R7325 GND.n5769 GND.n5768 19.3944
R7326 GND.n5768 GND.n5767 19.3944
R7327 GND.n5767 GND.n533 19.3944
R7328 GND.n5762 GND.n533 19.3944
R7329 GND.n5828 GND.n5827 19.3944
R7330 GND.n5827 GND.n5826 19.3944
R7331 GND.n5826 GND.n477 19.3944
R7332 GND.n5821 GND.n477 19.3944
R7333 GND.n5821 GND.n5820 19.3944
R7334 GND.n5820 GND.n5819 19.3944
R7335 GND.n5819 GND.n484 19.3944
R7336 GND.n5814 GND.n484 19.3944
R7337 GND.n5814 GND.n5813 19.3944
R7338 GND.n5813 GND.n5812 19.3944
R7339 GND.n5812 GND.n491 19.3944
R7340 GND.n5807 GND.n491 19.3944
R7341 GND.n5807 GND.n5806 19.3944
R7342 GND.n5806 GND.n5805 19.3944
R7343 GND.n5805 GND.n498 19.3944
R7344 GND.n5800 GND.n498 19.3944
R7345 GND.n5800 GND.n5799 19.3944
R7346 GND.n5756 GND.n5755 19.3944
R7347 GND.n5755 GND.n5754 19.3944
R7348 GND.n5754 GND.n546 19.3944
R7349 GND.n5749 GND.n546 19.3944
R7350 GND.n5749 GND.n5748 19.3944
R7351 GND.n5748 GND.n5747 19.3944
R7352 GND.n5747 GND.n553 19.3944
R7353 GND.n5742 GND.n553 19.3944
R7354 GND.n5742 GND.n5741 19.3944
R7355 GND.n5741 GND.n5740 19.3944
R7356 GND.n5740 GND.n560 19.3944
R7357 GND.n5735 GND.n560 19.3944
R7358 GND.n5735 GND.n5734 19.3944
R7359 GND.n5734 GND.n5733 19.3944
R7360 GND.n5733 GND.n567 19.3944
R7361 GND.n5728 GND.n567 19.3944
R7362 GND.n3991 GND.n3990 19.3944
R7363 GND.n3990 GND.n2781 19.3944
R7364 GND.n4110 GND.n2781 19.3944
R7365 GND.n4110 GND.n2779 19.3944
R7366 GND.n4114 GND.n2779 19.3944
R7367 GND.n4114 GND.n2777 19.3944
R7368 GND.n4125 GND.n2777 19.3944
R7369 GND.n4125 GND.n2775 19.3944
R7370 GND.n4129 GND.n2775 19.3944
R7371 GND.n4129 GND.n2773 19.3944
R7372 GND.n4140 GND.n2773 19.3944
R7373 GND.n4140 GND.n2771 19.3944
R7374 GND.n4144 GND.n2771 19.3944
R7375 GND.n4144 GND.n2768 19.3944
R7376 GND.n4155 GND.n2768 19.3944
R7377 GND.n4155 GND.n2766 19.3944
R7378 GND.n4159 GND.n2766 19.3944
R7379 GND.n4159 GND.n2764 19.3944
R7380 GND.n4170 GND.n2764 19.3944
R7381 GND.n4170 GND.n2762 19.3944
R7382 GND.n4174 GND.n2762 19.3944
R7383 GND.n4174 GND.n2760 19.3944
R7384 GND.n4185 GND.n2760 19.3944
R7385 GND.n4185 GND.n2758 19.3944
R7386 GND.n4199 GND.n2758 19.3944
R7387 GND.n4199 GND.n4198 19.3944
R7388 GND.n4198 GND.n4197 19.3944
R7389 GND.n4197 GND.n4196 19.3944
R7390 GND.n4196 GND.n4193 19.3944
R7391 GND.n4193 GND.n316 19.3944
R7392 GND.n5920 GND.n316 19.3944
R7393 GND.n5920 GND.n317 19.3944
R7394 GND.n2749 GND.n317 19.3944
R7395 GND.n4224 GND.n2749 19.3944
R7396 GND.n4224 GND.n2747 19.3944
R7397 GND.n4229 GND.n2747 19.3944
R7398 GND.n4229 GND.n2741 19.3944
R7399 GND.n4267 GND.n2741 19.3944
R7400 GND.n4267 GND.n4266 19.3944
R7401 GND.n4266 GND.n4265 19.3944
R7402 GND.n4265 GND.n2745 19.3944
R7403 GND.n4255 GND.n2745 19.3944
R7404 GND.n4255 GND.n4254 19.3944
R7405 GND.n4254 GND.n4253 19.3944
R7406 GND.n4253 GND.n4248 19.3944
R7407 GND.n4248 GND.n4247 19.3944
R7408 GND.n4247 GND.n586 19.3944
R7409 GND.n5701 GND.n586 19.3944
R7410 GND.n5702 GND.n5701 19.3944
R7411 GND.n5702 GND.n584 19.3944
R7412 GND.n5706 GND.n584 19.3944
R7413 GND.n5708 GND.n5706 19.3944
R7414 GND.n5709 GND.n5708 19.3944
R7415 GND.n5709 GND.n582 19.3944
R7416 GND.n5713 GND.n582 19.3944
R7417 GND.n5715 GND.n5713 19.3944
R7418 GND.n5716 GND.n5715 19.3944
R7419 GND.n5716 GND.n579 19.3944
R7420 GND.n5720 GND.n579 19.3944
R7421 GND.n5722 GND.n5720 19.3944
R7422 GND.n5723 GND.n5722 19.3944
R7423 GND.n2582 GND.n2581 19.3944
R7424 GND.n4397 GND.n2581 19.3944
R7425 GND.n4397 GND.n4396 19.3944
R7426 GND.n4396 GND.n4395 19.3944
R7427 GND.n4395 GND.n2588 19.3944
R7428 GND.n4385 GND.n2588 19.3944
R7429 GND.n4385 GND.n4384 19.3944
R7430 GND.n4384 GND.n4383 19.3944
R7431 GND.n4383 GND.n2612 19.3944
R7432 GND.n4373 GND.n2612 19.3944
R7433 GND.n4373 GND.n4372 19.3944
R7434 GND.n4372 GND.n4371 19.3944
R7435 GND.n4371 GND.n2633 19.3944
R7436 GND.n4361 GND.n2633 19.3944
R7437 GND.n4361 GND.n4360 19.3944
R7438 GND.n4360 GND.n4359 19.3944
R7439 GND.n4359 GND.n2653 19.3944
R7440 GND.n4349 GND.n2653 19.3944
R7441 GND.n4349 GND.n4348 19.3944
R7442 GND.n4348 GND.n4347 19.3944
R7443 GND.n4347 GND.n2674 19.3944
R7444 GND.n4337 GND.n2674 19.3944
R7445 GND.n4337 GND.n4336 19.3944
R7446 GND.n4336 GND.n4335 19.3944
R7447 GND.n4335 GND.n2695 19.3944
R7448 GND.n4325 GND.n2695 19.3944
R7449 GND.n2712 GND.n333 19.3944
R7450 GND.n2722 GND.n333 19.3944
R7451 GND.n5916 GND.n326 19.3944
R7452 GND.n2752 GND.n327 19.3944
R7453 GND.n5913 GND.n335 19.3944
R7454 GND.n5913 GND.n336 19.3944
R7455 GND.n5903 GND.n336 19.3944
R7456 GND.n5903 GND.n5902 19.3944
R7457 GND.n5902 GND.n5901 19.3944
R7458 GND.n5901 GND.n358 19.3944
R7459 GND.n5891 GND.n358 19.3944
R7460 GND.n5891 GND.n5890 19.3944
R7461 GND.n5890 GND.n5889 19.3944
R7462 GND.n5889 GND.n379 19.3944
R7463 GND.n5879 GND.n379 19.3944
R7464 GND.n5879 GND.n5878 19.3944
R7465 GND.n5878 GND.n5877 19.3944
R7466 GND.n5877 GND.n400 19.3944
R7467 GND.n5867 GND.n400 19.3944
R7468 GND.n5867 GND.n5866 19.3944
R7469 GND.n5866 GND.n5865 19.3944
R7470 GND.n5865 GND.n420 19.3944
R7471 GND.n5855 GND.n420 19.3944
R7472 GND.n5855 GND.n5854 19.3944
R7473 GND.n5854 GND.n5853 19.3944
R7474 GND.n5853 GND.n440 19.3944
R7475 GND.n5843 GND.n440 19.3944
R7476 GND.n5843 GND.n5842 19.3944
R7477 GND.n5842 GND.n5841 19.3944
R7478 GND.n5841 GND.n459 19.3944
R7479 GND.n5831 GND.n459 19.3944
R7480 GND.n4887 GND.n1113 19.3944
R7481 GND.n1627 GND.n1113 19.3944
R7482 GND.n1627 GND.n1625 19.3944
R7483 GND.n1631 GND.n1625 19.3944
R7484 GND.n1631 GND.n1623 19.3944
R7485 GND.n2009 GND.n1623 19.3944
R7486 GND.n2009 GND.n1621 19.3944
R7487 GND.n2015 GND.n1621 19.3944
R7488 GND.n2015 GND.n2014 19.3944
R7489 GND.n2014 GND.n1596 19.3944
R7490 GND.n2047 GND.n1596 19.3944
R7491 GND.n2047 GND.n1594 19.3944
R7492 GND.n2051 GND.n1594 19.3944
R7493 GND.n2051 GND.n1514 19.3944
R7494 GND.n2137 GND.n1514 19.3944
R7495 GND.n2137 GND.n1515 19.3944
R7496 GND.n1539 GND.n1538 19.3944
R7497 GND.n2121 GND.n2120 19.3944
R7498 GND.n1568 GND.n1567 19.3944
R7499 GND.n2104 GND.n2103 19.3944
R7500 GND.n1559 GND.n1506 19.3944
R7501 GND.n2193 GND.n1506 19.3944
R7502 GND.n2193 GND.n2192 19.3944
R7503 GND.n2192 GND.n2191 19.3944
R7504 GND.n2191 GND.n2144 19.3944
R7505 GND.n2187 GND.n2144 19.3944
R7506 GND.n2187 GND.n2186 19.3944
R7507 GND.n2186 GND.n2185 19.3944
R7508 GND.n2185 GND.n2150 19.3944
R7509 GND.n2181 GND.n2150 19.3944
R7510 GND.n2181 GND.n2180 19.3944
R7511 GND.n2180 GND.n2179 19.3944
R7512 GND.n2179 GND.n2158 19.3944
R7513 GND.n2175 GND.n2158 19.3944
R7514 GND.n2175 GND.n2174 19.3944
R7515 GND.n2174 GND.n2173 19.3944
R7516 GND.n2173 GND.n2168 19.3944
R7517 GND.n2168 GND.n2167 19.3944
R7518 GND.n2167 GND.n1427 19.3944
R7519 GND.n1427 GND.n1425 19.3944
R7520 GND.n2291 GND.n1425 19.3944
R7521 GND.n2291 GND.n1423 19.3944
R7522 GND.n2304 GND.n1423 19.3944
R7523 GND.n2304 GND.n2303 19.3944
R7524 GND.n2303 GND.n2302 19.3944
R7525 GND.n2302 GND.n2299 19.3944
R7526 GND.n2299 GND.n1309 19.3944
R7527 GND.n4708 GND.n1309 19.3944
R7528 GND.n4708 GND.n4707 19.3944
R7529 GND.n4707 GND.n4706 19.3944
R7530 GND.n4706 GND.n1313 19.3944
R7531 GND.n3398 GND.n1313 19.3944
R7532 GND.n3413 GND.n3398 19.3944
R7533 GND.n3413 GND.n3395 19.3944
R7534 GND.n3417 GND.n3395 19.3944
R7535 GND.n3417 GND.n3385 19.3944
R7536 GND.n3433 GND.n3385 19.3944
R7537 GND.n3433 GND.n3383 19.3944
R7538 GND.n3437 GND.n3383 19.3944
R7539 GND.n3437 GND.n3372 19.3944
R7540 GND.n3453 GND.n3372 19.3944
R7541 GND.n3453 GND.n3370 19.3944
R7542 GND.n3457 GND.n3370 19.3944
R7543 GND.n3457 GND.n3176 19.3944
R7544 GND.n3474 GND.n3176 19.3944
R7545 GND.n3474 GND.n3174 19.3944
R7546 GND.n3478 GND.n3174 19.3944
R7547 GND.n3478 GND.n3139 19.3944
R7548 GND.n3508 GND.n3139 19.3944
R7549 GND.n3508 GND.n3137 19.3944
R7550 GND.n3514 GND.n3137 19.3944
R7551 GND.n3514 GND.n3513 19.3944
R7552 GND.n3513 GND.n3109 19.3944
R7553 GND.n3550 GND.n3109 19.3944
R7554 GND.n3550 GND.n3107 19.3944
R7555 GND.n3571 GND.n3107 19.3944
R7556 GND.n3571 GND.n3570 19.3944
R7557 GND.n3570 GND.n3569 19.3944
R7558 GND.n3569 GND.n3556 19.3944
R7559 GND.n3565 GND.n3556 19.3944
R7560 GND.n3565 GND.n3564 19.3944
R7561 GND.n3564 GND.n3563 19.3944
R7562 GND.n3563 GND.n3063 19.3944
R7563 GND.n3666 GND.n3063 19.3944
R7564 GND.n3666 GND.n3061 19.3944
R7565 GND.n3672 GND.n3061 19.3944
R7566 GND.n3672 GND.n3671 19.3944
R7567 GND.n3671 GND.n3034 19.3944
R7568 GND.n3710 GND.n3034 19.3944
R7569 GND.n3710 GND.n3032 19.3944
R7570 GND.n3719 GND.n3032 19.3944
R7571 GND.n3719 GND.n3718 19.3944
R7572 GND.n3718 GND.n3717 19.3944
R7573 GND.n3717 GND.n2998 19.3944
R7574 GND.n3770 GND.n2998 19.3944
R7575 GND.n3770 GND.n2996 19.3944
R7576 GND.n3776 GND.n2996 19.3944
R7577 GND.n3776 GND.n3775 19.3944
R7578 GND.n3775 GND.n2975 19.3944
R7579 GND.n3795 GND.n2975 19.3944
R7580 GND.n3795 GND.n2973 19.3944
R7581 GND.n3799 GND.n2973 19.3944
R7582 GND.n3799 GND.n2836 19.3944
R7583 GND.n3898 GND.n2836 19.3944
R7584 GND.n3898 GND.n2834 19.3944
R7585 GND.n3902 GND.n2834 19.3944
R7586 GND.n3902 GND.n2823 19.3944
R7587 GND.n3917 GND.n2823 19.3944
R7588 GND.n3917 GND.n2821 19.3944
R7589 GND.n3921 GND.n2821 19.3944
R7590 GND.n3921 GND.n2809 19.3944
R7591 GND.n3936 GND.n2809 19.3944
R7592 GND.n3936 GND.n2807 19.3944
R7593 GND.n3942 GND.n2807 19.3944
R7594 GND.n3942 GND.n3941 19.3944
R7595 GND.n3941 GND.n2795 19.3944
R7596 GND.n3958 GND.n2795 19.3944
R7597 GND.n3958 GND.n2793 19.3944
R7598 GND.n3962 GND.n2793 19.3944
R7599 GND.n3962 GND.n2790 19.3944
R7600 GND.n4025 GND.n2790 19.3944
R7601 GND.n4025 GND.n2788 19.3944
R7602 GND.n4029 GND.n2788 19.3944
R7603 GND.n4029 GND.n2786 19.3944
R7604 GND.n4033 GND.n2786 19.3944
R7605 GND.n4033 GND.n2784 19.3944
R7606 GND.n4105 GND.n2784 19.3944
R7607 GND.n4105 GND.n4104 19.3944
R7608 GND.n4104 GND.n4103 19.3944
R7609 GND.n4103 GND.n4039 19.3944
R7610 GND.n4099 GND.n4039 19.3944
R7611 GND.n4099 GND.n4098 19.3944
R7612 GND.n4098 GND.n4097 19.3944
R7613 GND.n4097 GND.n4045 19.3944
R7614 GND.n4093 GND.n4045 19.3944
R7615 GND.n4093 GND.n4092 19.3944
R7616 GND.n4092 GND.n4091 19.3944
R7617 GND.n4091 GND.n4051 19.3944
R7618 GND.n4087 GND.n4051 19.3944
R7619 GND.n4087 GND.n4086 19.3944
R7620 GND.n4086 GND.n4085 19.3944
R7621 GND.n4085 GND.n4057 19.3944
R7622 GND.n4081 GND.n4057 19.3944
R7623 GND.n4081 GND.n4080 19.3944
R7624 GND.n4080 GND.n4079 19.3944
R7625 GND.n4079 GND.n4063 19.3944
R7626 GND.n4075 GND.n4063 19.3944
R7627 GND.n4075 GND.n4074 19.3944
R7628 GND.n4074 GND.n4073 19.3944
R7629 GND.n4073 GND.n4070 19.3944
R7630 GND.n4320 GND.n2718 19.3944
R7631 GND.n4318 GND.n4317 19.3944
R7632 GND.n2737 GND.n2736 19.3944
R7633 GND.n4305 GND.n4304 19.3944
R7634 GND.n4302 GND.n2739 19.3944
R7635 GND.n4298 GND.n2739 19.3944
R7636 GND.n4298 GND.n4297 19.3944
R7637 GND.n4297 GND.n4296 19.3944
R7638 GND.n4296 GND.n4276 19.3944
R7639 GND.n4292 GND.n4276 19.3944
R7640 GND.n4292 GND.n4291 19.3944
R7641 GND.n4291 GND.n4290 19.3944
R7642 GND.n4290 GND.n4282 19.3944
R7643 GND.n4286 GND.n4282 19.3944
R7644 GND.n4286 GND.n592 19.3944
R7645 GND.n5666 GND.n592 19.3944
R7646 GND.n5666 GND.n5665 19.3944
R7647 GND.n5665 GND.n5664 19.3944
R7648 GND.n5664 GND.n596 19.3944
R7649 GND.n5660 GND.n596 19.3944
R7650 GND.n1912 GND.n1911 19.3944
R7651 GND.n1911 GND.n1702 19.3944
R7652 GND.n1906 GND.n1702 19.3944
R7653 GND.n1906 GND.n1905 19.3944
R7654 GND.n1905 GND.n1707 19.3944
R7655 GND.n1900 GND.n1707 19.3944
R7656 GND.n1900 GND.n1899 19.3944
R7657 GND.n1899 GND.n1898 19.3944
R7658 GND.n1898 GND.n1713 19.3944
R7659 GND.n1892 GND.n1713 19.3944
R7660 GND.n1892 GND.n1891 19.3944
R7661 GND.n1891 GND.n1890 19.3944
R7662 GND.n1890 GND.n1719 19.3944
R7663 GND.n1884 GND.n1719 19.3944
R7664 GND.n1884 GND.n1883 19.3944
R7665 GND.n1883 GND.n1882 19.3944
R7666 GND.n1882 GND.n1725 19.3944
R7667 GND.n1876 GND.n1875 19.3944
R7668 GND.n1875 GND.n1874 19.3944
R7669 GND.n1874 GND.n1734 19.3944
R7670 GND.n1868 GND.n1734 19.3944
R7671 GND.n1868 GND.n1867 19.3944
R7672 GND.n1867 GND.n1866 19.3944
R7673 GND.n1866 GND.n1740 19.3944
R7674 GND.n1860 GND.n1740 19.3944
R7675 GND.n1860 GND.n1859 19.3944
R7676 GND.n1859 GND.n1858 19.3944
R7677 GND.n1858 GND.n1746 19.3944
R7678 GND.n1852 GND.n1746 19.3944
R7679 GND.n1852 GND.n1851 19.3944
R7680 GND.n1851 GND.n1850 19.3944
R7681 GND.n1850 GND.n1752 19.3944
R7682 GND.n1844 GND.n1752 19.3944
R7683 GND.n1844 GND.n1843 19.3944
R7684 GND.n1843 GND.n1842 19.3944
R7685 GND.n1917 GND.n1916 19.3944
R7686 GND.n1916 GND.n1676 19.3944
R7687 GND.n1950 GND.n1676 19.3944
R7688 GND.n1950 GND.n1674 19.3944
R7689 GND.n1954 GND.n1674 19.3944
R7690 GND.n1954 GND.n1657 19.3944
R7691 GND.n1979 GND.n1657 19.3944
R7692 GND.n1979 GND.n1655 19.3944
R7693 GND.n1984 GND.n1655 19.3944
R7694 GND.n1984 GND.n1122 19.3944
R7695 GND.n4882 GND.n1122 19.3944
R7696 GND.n4882 GND.n4881 19.3944
R7697 GND.n4881 GND.n4880 19.3944
R7698 GND.n4880 GND.n1126 19.3944
R7699 GND.n1636 GND.n1126 19.3944
R7700 GND.n1636 GND.n1613 19.3944
R7701 GND.n2023 GND.n1613 19.3944
R7702 GND.n2023 GND.n1611 19.3944
R7703 GND.n2029 GND.n1611 19.3944
R7704 GND.n2029 GND.n2028 19.3944
R7705 GND.n2028 GND.n1587 19.3944
R7706 GND.n2060 GND.n1587 19.3944
R7707 GND.n2060 GND.n1585 19.3944
R7708 GND.n2065 GND.n1585 19.3944
R7709 GND.n2065 GND.n1525 19.3944
R7710 GND.n2132 GND.n1525 19.3944
R7711 GND.n2130 GND.n2129 19.3944
R7712 GND.n2129 GND.n1526 19.3944
R7713 GND.n2115 GND.n1548 19.3944
R7714 GND.n2113 GND.n2112 19.3944
R7715 GND.n2096 GND.n2095 19.3944
R7716 GND.n2098 GND.n2096 19.3944
R7717 GND.n2098 GND.n1497 19.3944
R7718 GND.n2204 GND.n1497 19.3944
R7719 GND.n2204 GND.n1495 19.3944
R7720 GND.n2210 GND.n1495 19.3944
R7721 GND.n2210 GND.n2209 19.3944
R7722 GND.n2209 GND.n1474 19.3944
R7723 GND.n2229 GND.n1474 19.3944
R7724 GND.n2229 GND.n1472 19.3944
R7725 GND.n2235 GND.n1472 19.3944
R7726 GND.n2235 GND.n2234 19.3944
R7727 GND.n2234 GND.n1453 19.3944
R7728 GND.n2253 GND.n1453 19.3944
R7729 GND.n2253 GND.n1451 19.3944
R7730 GND.n2259 GND.n1451 19.3944
R7731 GND.n2259 GND.n2258 19.3944
R7732 GND.n2258 GND.n1432 19.3944
R7733 GND.n2280 GND.n1432 19.3944
R7734 GND.n2280 GND.n1430 19.3944
R7735 GND.n2284 GND.n1430 19.3944
R7736 GND.n2284 GND.n1408 19.3944
R7737 GND.n2320 GND.n1408 19.3944
R7738 GND.n2320 GND.n1406 19.3944
R7739 GND.n2324 GND.n1406 19.3944
R7740 GND.n2324 GND.n1242 19.3944
R7741 GND.n4798 GND.n1242 19.3944
R7742 GND.n5027 GND.n5026 19.3944
R7743 GND.n5026 GND.n5025 19.3944
R7744 GND.n5025 GND.n978 19.3944
R7745 GND.n5019 GND.n978 19.3944
R7746 GND.n5019 GND.n5018 19.3944
R7747 GND.n5018 GND.n5017 19.3944
R7748 GND.n5017 GND.n986 19.3944
R7749 GND.n5011 GND.n986 19.3944
R7750 GND.n5011 GND.n5010 19.3944
R7751 GND.n5010 GND.n5009 19.3944
R7752 GND.n5009 GND.n994 19.3944
R7753 GND.n5003 GND.n994 19.3944
R7754 GND.n5003 GND.n5002 19.3944
R7755 GND.n5002 GND.n5001 19.3944
R7756 GND.n5001 GND.n1002 19.3944
R7757 GND.n4995 GND.n1002 19.3944
R7758 GND.n4995 GND.n4994 19.3944
R7759 GND.n4994 GND.n4993 19.3944
R7760 GND.n4993 GND.n1010 19.3944
R7761 GND.n4987 GND.n1010 19.3944
R7762 GND.n4987 GND.n4986 19.3944
R7763 GND.n4986 GND.n4985 19.3944
R7764 GND.n4985 GND.n1018 19.3944
R7765 GND.n4979 GND.n1018 19.3944
R7766 GND.n4979 GND.n4978 19.3944
R7767 GND.n4978 GND.n4977 19.3944
R7768 GND.n4977 GND.n1026 19.3944
R7769 GND.n4971 GND.n1026 19.3944
R7770 GND.n4971 GND.n4970 19.3944
R7771 GND.n4970 GND.n4969 19.3944
R7772 GND.n4969 GND.n1034 19.3944
R7773 GND.n4963 GND.n1034 19.3944
R7774 GND.n4963 GND.n4962 19.3944
R7775 GND.n4962 GND.n4961 19.3944
R7776 GND.n4961 GND.n1042 19.3944
R7777 GND.n4955 GND.n1042 19.3944
R7778 GND.n4955 GND.n4954 19.3944
R7779 GND.n4954 GND.n4953 19.3944
R7780 GND.n4953 GND.n1050 19.3944
R7781 GND.n4947 GND.n1050 19.3944
R7782 GND.n4947 GND.n4946 19.3944
R7783 GND.n4946 GND.n4945 19.3944
R7784 GND.n4945 GND.n1058 19.3944
R7785 GND.n4939 GND.n1058 19.3944
R7786 GND.n4939 GND.n4938 19.3944
R7787 GND.n4938 GND.n4937 19.3944
R7788 GND.n4937 GND.n1066 19.3944
R7789 GND.n4931 GND.n1066 19.3944
R7790 GND.n4931 GND.n4930 19.3944
R7791 GND.n4930 GND.n4929 19.3944
R7792 GND.n4929 GND.n1074 19.3944
R7793 GND.n4923 GND.n1074 19.3944
R7794 GND.n4923 GND.n4922 19.3944
R7795 GND.n4922 GND.n4921 19.3944
R7796 GND.n4921 GND.n1082 19.3944
R7797 GND.n4915 GND.n1082 19.3944
R7798 GND.n4915 GND.n4914 19.3944
R7799 GND.n4914 GND.n4913 19.3944
R7800 GND.n4913 GND.n1090 19.3944
R7801 GND.n4907 GND.n1090 19.3944
R7802 GND.n4907 GND.n4906 19.3944
R7803 GND.n4906 GND.n4905 19.3944
R7804 GND.n4905 GND.n1098 19.3944
R7805 GND.n4899 GND.n1098 19.3944
R7806 GND.n4899 GND.n4898 19.3944
R7807 GND.n4898 GND.n4897 19.3944
R7808 GND.n4897 GND.n1106 19.3944
R7809 GND.n4891 GND.n1106 19.3944
R7810 GND.n4891 GND.n4890 19.3944
R7811 GND.n4533 GND.n4532 19.3944
R7812 GND.n4532 GND.n2437 19.3944
R7813 GND.n4525 GND.n2437 19.3944
R7814 GND.n4525 GND.n4524 19.3944
R7815 GND.n4524 GND.n2446 19.3944
R7816 GND.n4517 GND.n2446 19.3944
R7817 GND.n4517 GND.n4516 19.3944
R7818 GND.n4516 GND.n2454 19.3944
R7819 GND.n4509 GND.n2454 19.3944
R7820 GND.n4509 GND.n4508 19.3944
R7821 GND.n4508 GND.n2462 19.3944
R7822 GND.n4501 GND.n2462 19.3944
R7823 GND.n4501 GND.n4500 19.3944
R7824 GND.n4500 GND.n2470 19.3944
R7825 GND.n4493 GND.n2470 19.3944
R7826 GND.n4493 GND.n4492 19.3944
R7827 GND.n4492 GND.n2478 19.3944
R7828 GND.n3997 GND.n2478 19.3944
R7829 GND.n4000 GND.n3997 19.3944
R7830 GND.n4000 GND.n3986 19.3944
R7831 GND.n4005 GND.n3986 19.3944
R7832 GND.n4008 GND.n4005 19.3944
R7833 GND.n4013 GND.n3983 19.3944
R7834 GND.n4018 GND.n3983 19.3944
R7835 GND.n4018 GND.n3984 19.3944
R7836 GND.n3408 GND.n3404 19.3944
R7837 GND.n3408 GND.n3392 19.3944
R7838 GND.n3424 GND.n3392 19.3944
R7839 GND.n3424 GND.n3390 19.3944
R7840 GND.n3428 GND.n3390 19.3944
R7841 GND.n3428 GND.n3379 19.3944
R7842 GND.n3444 GND.n3379 19.3944
R7843 GND.n3444 GND.n3377 19.3944
R7844 GND.n3448 GND.n3377 19.3944
R7845 GND.n3448 GND.n3366 19.3944
R7846 GND.n3465 GND.n3366 19.3944
R7847 GND.n3465 GND.n3364 19.3944
R7848 GND.n3469 GND.n3364 19.3944
R7849 GND.n3469 GND.n3170 19.3944
R7850 GND.n3484 GND.n3170 19.3944
R7851 GND.n3484 GND.n3168 19.3944
R7852 GND.n3488 GND.n3168 19.3944
R7853 GND.n3488 GND.n3124 19.3944
R7854 GND.n3527 GND.n3124 19.3944
R7855 GND.n3527 GND.n3121 19.3944
R7856 GND.n3538 GND.n3121 19.3944
R7857 GND.n3538 GND.n3122 19.3944
R7858 GND.n3534 GND.n3122 19.3944
R7859 GND.n3534 GND.n3533 19.3944
R7860 GND.n3533 GND.n3087 19.3944
R7861 GND.n3600 GND.n3087 19.3944
R7862 GND.n3600 GND.n3085 19.3944
R7863 GND.n3604 GND.n3085 19.3944
R7864 GND.n3604 GND.n3070 19.3944
R7865 GND.n3657 GND.n3070 19.3944
R7866 GND.n3657 GND.n3068 19.3944
R7867 GND.n3661 GND.n3068 19.3944
R7868 GND.n3661 GND.n3049 19.3944
R7869 GND.n3685 GND.n3049 19.3944
R7870 GND.n3685 GND.n3046 19.3944
R7871 GND.n3698 GND.n3046 19.3944
R7872 GND.n3698 GND.n3047 19.3944
R7873 GND.n3694 GND.n3047 19.3944
R7874 GND.n3694 GND.n3693 19.3944
R7875 GND.n3693 GND.n3007 19.3944
R7876 GND.n3751 GND.n3007 19.3944
R7877 GND.n3751 GND.n3004 19.3944
R7878 GND.n3765 GND.n3004 19.3944
R7879 GND.n3765 GND.n3005 19.3944
R7880 GND.n3761 GND.n3005 19.3944
R7881 GND.n3761 GND.n3760 19.3944
R7882 GND.n3760 GND.n3759 19.3944
R7883 GND.n3759 GND.n2899 19.3944
R7884 GND.n3820 GND.n2899 19.3944
R7885 GND.n3820 GND.n2897 19.3944
R7886 GND.n3824 GND.n2897 19.3944
R7887 GND.n3824 GND.n2830 19.3944
R7888 GND.n3907 GND.n2830 19.3944
R7889 GND.n3907 GND.n2828 19.3944
R7890 GND.n3911 GND.n2828 19.3944
R7891 GND.n3911 GND.n2816 19.3944
R7892 GND.n3926 GND.n2816 19.3944
R7893 GND.n3926 GND.n2814 19.3944
R7894 GND.n3930 GND.n2814 19.3944
R7895 GND.n3930 GND.n2801 19.3944
R7896 GND.n3947 GND.n2801 19.3944
R7897 GND.n3947 GND.n2799 19.3944
R7898 GND.n3951 GND.n2799 19.3944
R7899 GND.n3951 GND.n2432 19.3944
R7900 GND.n4537 GND.n2432 19.3944
R7901 GND.n4771 GND.n1262 18.4247
R7902 GND.n4452 GND.n4451 18.4247
R7903 GND.n4489 GND.n4488 18.2308
R7904 GND.n4656 GND.n4655 18.2308
R7905 GND.n1805 GND.n1804 18.2308
R7906 GND.n5728 GND.n5727 18.2308
R7907 GND.n1986 GND.t119 17.6511
R7908 GND.n2273 GND.t117 17.6511
R7909 GND.n4131 GND.t134 17.6511
R7910 GND.n431 GND.t125 17.6511
R7911 GND.n4703 GND.n1327 17.3181
R7912 GND.n4021 GND.n3964 17.3181
R7913 GND.n2202 GND.t156 16.9851
R7914 GND.n4183 GND.t123 16.9851
R7915 GND.n3401 GND.n3400 16.652
R7916 GND.n3411 GND.n3401 16.652
R7917 GND.n3411 GND.n3410 16.652
R7918 GND.n3410 GND.n3403 16.652
R7919 GND.n3403 GND.n3402 16.652
R7920 GND.n3422 GND.n3419 16.652
R7921 GND.n3422 GND.n3421 16.652
R7922 GND.n3421 GND.n3387 16.652
R7923 GND.n3431 GND.n3387 16.652
R7924 GND.n3431 GND.n3430 16.652
R7925 GND.n3430 GND.n3388 16.652
R7926 GND.n3388 GND.n3381 16.652
R7927 GND.n3439 GND.n3381 16.652
R7928 GND.n3442 GND.n3439 16.652
R7929 GND.n3442 GND.n3441 16.652
R7930 GND.n3441 GND.n3374 16.652
R7931 GND.n3451 GND.n3374 16.652
R7932 GND.n3451 GND.n3450 16.652
R7933 GND.n3375 GND.n3368 16.652
R7934 GND.n3459 GND.n3368 16.652
R7935 GND.n3463 GND.n3459 16.652
R7936 GND.n3463 GND.n3462 16.652
R7937 GND.n3462 GND.n3461 16.652
R7938 GND.n3472 GND.n3471 16.652
R7939 GND.n3482 GND.n3480 16.652
R7940 GND.n3506 GND.n3141 16.652
R7941 GND.n3573 GND.n3104 16.652
R7942 GND.n3104 GND.n3097 16.652
R7943 GND.n3598 GND.n3089 16.652
R7944 GND.n3606 GND.n3083 16.652
R7945 GND.n3655 GND.n3072 16.652
R7946 GND.n3664 GND.n3663 16.652
R7947 GND.n3675 GND.n3674 16.652
R7948 GND.n3624 GND.n3042 16.652
R7949 GND.n3615 GND.n3038 16.652
R7950 GND.n3691 GND.n3023 16.652
R7951 GND.n3749 GND.n3009 16.652
R7952 GND.n3749 GND.n3011 16.652
R7953 GND.n3778 GND.n2993 16.652
R7954 GND.n2985 GND.n2978 16.652
R7955 GND.n3818 GND.n2901 16.652
R7956 GND.n3802 GND.n2893 16.652
R7957 GND.n3896 GND.n3895 16.652
R7958 GND.n3895 GND.n3894 16.652
R7959 GND.n3905 GND.n3904 16.652
R7960 GND.n3904 GND.n2832 16.652
R7961 GND.n2832 GND.n2825 16.652
R7962 GND.n3913 GND.n2825 16.652
R7963 GND.n3915 GND.n3913 16.652
R7964 GND.n3914 GND.n2818 16.652
R7965 GND.n3924 GND.n2818 16.652
R7966 GND.n3924 GND.n3923 16.652
R7967 GND.n3923 GND.n2819 16.652
R7968 GND.n2819 GND.n2811 16.652
R7969 GND.n3932 GND.n2811 16.652
R7970 GND.n3934 GND.n3932 16.652
R7971 GND.n3934 GND.n3933 16.652
R7972 GND.n3933 GND.n2803 16.652
R7973 GND.n3945 GND.n2803 16.652
R7974 GND.n3945 GND.n3944 16.652
R7975 GND.n3944 GND.n2805 16.652
R7976 GND.n2805 GND.n2804 16.652
R7977 GND.n3955 GND.n3953 16.652
R7978 GND.n3955 GND.n3954 16.652
R7979 GND.n3954 GND.n2428 16.652
R7980 GND.n4539 GND.n2428 16.652
R7981 GND.n4539 GND.n2429 16.652
R7982 GND.n2067 GND.t141 16.319
R7983 GND.n3402 GND.t70 16.319
R7984 GND.n3953 GND.t80 16.319
R7985 GND.n5905 GND.t151 16.319
R7986 GND.n4704 GND.n4703 15.986
R7987 GND.n3180 GND.n3172 15.986
R7988 GND.n3636 GND.n3065 15.986
R7989 GND.n3683 GND.n3051 15.986
R7990 GND.n3810 GND.n3809 15.986
R7991 GND.n3827 GND.n3826 15.986
R7992 GND.n4022 GND.n4021 15.986
R7993 GND.n136 GND.n134 15.6674
R7994 GND.n104 GND.n102 15.6674
R7995 GND.n72 GND.n70 15.6674
R7996 GND.n41 GND.n39 15.6674
R7997 GND.n263 GND.n261 15.6674
R7998 GND.n231 GND.n229 15.6674
R7999 GND.n199 GND.n197 15.6674
R8000 GND.n168 GND.n166 15.6674
R8001 GND.t119 GND.n1115 15.6529
R8002 GND.n5863 GND.t125 15.6529
R8003 GND.n3548 GND.n3547 15.3199
R8004 GND.n3597 GND.n3091 15.3199
R8005 GND.n3721 GND.n3029 15.3199
R8006 GND.n3736 GND.n3001 15.3199
R8007 GND.n2876 GND.n2875 15.0827
R8008 GND.n3190 GND.n3185 15.0481
R8009 GND.n2886 GND.n2885 15.0481
R8010 GND.n3461 GND.n3178 14.9869
R8011 GND.n3471 GND.t55 14.6538
R8012 GND.n3525 GND.n3126 14.6538
R8013 GND.n3517 GND.t84 13.9878
R8014 GND.n3160 GND.n3129 13.9878
R8015 GND.t16 GND.n3117 13.9878
R8016 GND.n3607 GND.n3079 13.9878
R8017 GND.n3708 GND.n3707 13.9878
R8018 GND.n2992 GND.n2982 13.9878
R8019 GND.n4741 GND.n1290 13.5763
R8020 GND.n4414 GND.n2563 13.5763
R8021 GND.n5762 GND.n5761 13.5763
R8022 GND.n1842 GND.n1761 13.5763
R8023 GND.n3541 GND.n3540 13.3217
R8024 GND.n3151 GND.t99 13.3217
R8025 GND.n3591 GND.n3590 13.3217
R8026 GND.n3616 GND.n3027 13.3217
R8027 GND.n3768 GND.t100 13.3217
R8028 GND.n3779 GND.n2990 13.3217
R8029 GND.n3201 GND.n3182 13.1884
R8030 GND.n3196 GND.n3195 13.1884
R8031 GND.n3195 GND.n3194 13.1884
R8032 GND.n2879 GND.n2874 13.1884
R8033 GND.n2880 GND.n2879 13.1884
R8034 GND.n3197 GND.n3184 13.146
R8035 GND.n3193 GND.n3184 13.146
R8036 GND.n2878 GND.n2877 13.146
R8037 GND.n2878 GND.n2873 13.146
R8038 GND.n3358 GND.n3357 12.8005
R8039 GND.n3891 GND.n3831 12.8005
R8040 GND.n137 GND.n133 12.8005
R8041 GND.n105 GND.n101 12.8005
R8042 GND.n73 GND.n69 12.8005
R8043 GND.n42 GND.n38 12.8005
R8044 GND.n264 GND.n260 12.8005
R8045 GND.n232 GND.n228 12.8005
R8046 GND.n200 GND.n196 12.8005
R8047 GND.n169 GND.n165 12.8005
R8048 GND.n4737 GND.n4710 12.6557
R8049 GND.n3518 GND.n3133 12.6557
R8050 GND.n3654 GND.n3074 12.6557
R8051 GND.n3625 GND.n3053 12.6557
R8052 GND.n2986 GND.t74 12.6557
R8053 GND.n3793 GND.n3792 12.6557
R8054 GND.n4483 GND.n2484 12.6557
R8055 GND.n4741 GND.n4740 12.4126
R8056 GND.n4410 GND.n2563 12.4126
R8057 GND.n5761 GND.n540 12.4126
R8058 GND.n1838 GND.n1761 12.4126
R8059 GND.n141 GND.n140 12.0247
R8060 GND.n109 GND.n108 12.0247
R8061 GND.n77 GND.n76 12.0247
R8062 GND.n46 GND.n45 12.0247
R8063 GND.n268 GND.n267 12.0247
R8064 GND.n236 GND.n235 12.0247
R8065 GND.n204 GND.n203 12.0247
R8066 GND.n173 GND.n172 12.0247
R8067 GND.n3152 GND.n3102 11.9896
R8068 GND.n3582 GND.n3581 11.9896
R8069 GND.n3729 GND.n3728 11.9896
R8070 GND.n3743 GND.n3017 11.9896
R8071 GND.n3499 GND.n3498 11.3235
R8072 GND.n3498 GND.n3497 11.3235
R8073 GND.n3066 GND.n3057 11.3235
R8074 GND.n3676 GND.n3057 11.3235
R8075 GND.n3803 GND.n3801 11.3235
R8076 GND.n144 GND.n131 11.249
R8077 GND.n112 GND.n99 11.249
R8078 GND.n80 GND.n67 11.249
R8079 GND.n49 GND.n36 11.249
R8080 GND.n271 GND.n258 11.249
R8081 GND.n239 GND.n226 11.249
R8082 GND.n207 GND.n194 11.249
R8083 GND.n176 GND.n163 11.249
R8084 GND.n3450 GND.t103 10.9905
R8085 GND.t93 GND.n3914 10.9905
R8086 GND.n3574 GND.n3102 10.6575
R8087 GND.n3018 GND.n3017 10.6575
R8088 GND.n2914 GND.n2911 10.6151
R8089 GND.n2915 GND.n2914 10.6151
R8090 GND.n2919 GND.n2918 10.6151
R8091 GND.n2922 GND.n2919 10.6151
R8092 GND.n2923 GND.n2922 10.6151
R8093 GND.n2926 GND.n2923 10.6151
R8094 GND.n2927 GND.n2926 10.6151
R8095 GND.n2930 GND.n2927 10.6151
R8096 GND.n2931 GND.n2930 10.6151
R8097 GND.n2934 GND.n2931 10.6151
R8098 GND.n2935 GND.n2934 10.6151
R8099 GND.n2938 GND.n2935 10.6151
R8100 GND.n2939 GND.n2938 10.6151
R8101 GND.n2942 GND.n2939 10.6151
R8102 GND.n2943 GND.n2942 10.6151
R8103 GND.n2946 GND.n2943 10.6151
R8104 GND.n2947 GND.n2946 10.6151
R8105 GND.n2950 GND.n2947 10.6151
R8106 GND.n2951 GND.n2950 10.6151
R8107 GND.n2954 GND.n2951 10.6151
R8108 GND.n2955 GND.n2954 10.6151
R8109 GND.n2958 GND.n2955 10.6151
R8110 GND.n2959 GND.n2958 10.6151
R8111 GND.n2962 GND.n2959 10.6151
R8112 GND.n2963 GND.n2962 10.6151
R8113 GND.n2966 GND.n2963 10.6151
R8114 GND.n2967 GND.n2966 10.6151
R8115 GND.n3238 GND.n3237 10.6151
R8116 GND.n3237 GND.n3147 10.6151
R8117 GND.n3495 GND.n3147 10.6151
R8118 GND.n3495 GND.n3494 10.6151
R8119 GND.n3494 GND.n3493 10.6151
R8120 GND.n3493 GND.n3166 10.6151
R8121 GND.n3166 GND.n3165 10.6151
R8122 GND.n3165 GND.n3163 10.6151
R8123 GND.n3163 GND.n3162 10.6151
R8124 GND.n3162 GND.n3158 10.6151
R8125 GND.n3158 GND.n3157 10.6151
R8126 GND.n3157 GND.n3155 10.6151
R8127 GND.n3155 GND.n3154 10.6151
R8128 GND.n3154 GND.n3150 10.6151
R8129 GND.n3150 GND.n3149 10.6151
R8130 GND.n3149 GND.n3095 10.6151
R8131 GND.n3584 GND.n3095 10.6151
R8132 GND.n3585 GND.n3584 10.6151
R8133 GND.n3586 GND.n3585 10.6151
R8134 GND.n3586 GND.n3081 10.6151
R8135 GND.n3609 GND.n3081 10.6151
R8136 GND.n3610 GND.n3609 10.6151
R8137 GND.n3641 GND.n3610 10.6151
R8138 GND.n3641 GND.n3640 10.6151
R8139 GND.n3640 GND.n3639 10.6151
R8140 GND.n3639 GND.n3611 10.6151
R8141 GND.n3632 GND.n3611 10.6151
R8142 GND.n3632 GND.n3631 10.6151
R8143 GND.n3631 GND.n3630 10.6151
R8144 GND.n3630 GND.n3628 10.6151
R8145 GND.n3628 GND.n3627 10.6151
R8146 GND.n3627 GND.n3622 10.6151
R8147 GND.n3622 GND.n3621 10.6151
R8148 GND.n3621 GND.n3619 10.6151
R8149 GND.n3619 GND.n3618 10.6151
R8150 GND.n3618 GND.n3614 10.6151
R8151 GND.n3614 GND.n3613 10.6151
R8152 GND.n3613 GND.n3021 10.6151
R8153 GND.n3732 GND.n3021 10.6151
R8154 GND.n3733 GND.n3732 10.6151
R8155 GND.n3734 GND.n3733 10.6151
R8156 GND.n3741 GND.n3734 10.6151
R8157 GND.n3741 GND.n3740 10.6151
R8158 GND.n3740 GND.n3739 10.6151
R8159 GND.n3739 GND.n3735 10.6151
R8160 GND.n3735 GND.n2980 10.6151
R8161 GND.n3788 GND.n2980 10.6151
R8162 GND.n3789 GND.n3788 10.6151
R8163 GND.n3790 GND.n3789 10.6151
R8164 GND.n3790 GND.n2907 10.6151
R8165 GND.n3807 GND.n2907 10.6151
R8166 GND.n3807 GND.n3806 10.6151
R8167 GND.n3806 GND.n3805 10.6151
R8168 GND.n3805 GND.n2971 10.6151
R8169 GND.n2971 GND.n2970 10.6151
R8170 GND.n3295 GND.n3294 10.6151
R8171 GND.n3294 GND.n3293 10.6151
R8172 GND.n3289 GND.n3288 10.6151
R8173 GND.n3288 GND.n3224 10.6151
R8174 GND.n3283 GND.n3224 10.6151
R8175 GND.n3283 GND.n3282 10.6151
R8176 GND.n3282 GND.n3281 10.6151
R8177 GND.n3281 GND.n3226 10.6151
R8178 GND.n3275 GND.n3226 10.6151
R8179 GND.n3275 GND.n3274 10.6151
R8180 GND.n3274 GND.n3273 10.6151
R8181 GND.n3273 GND.n3228 10.6151
R8182 GND.n3267 GND.n3228 10.6151
R8183 GND.n3267 GND.n3266 10.6151
R8184 GND.n3266 GND.n3265 10.6151
R8185 GND.n3265 GND.n3230 10.6151
R8186 GND.n3259 GND.n3230 10.6151
R8187 GND.n3259 GND.n3258 10.6151
R8188 GND.n3258 GND.n3257 10.6151
R8189 GND.n3257 GND.n3232 10.6151
R8190 GND.n3251 GND.n3232 10.6151
R8191 GND.n3251 GND.n3250 10.6151
R8192 GND.n3250 GND.n3249 10.6151
R8193 GND.n3249 GND.n3234 10.6151
R8194 GND.n3243 GND.n3234 10.6151
R8195 GND.n3243 GND.n3242 10.6151
R8196 GND.n3242 GND.n3241 10.6151
R8197 GND.n3357 GND.n3356 10.6151
R8198 GND.n3356 GND.n3202 10.6151
R8199 GND.n3351 GND.n3202 10.6151
R8200 GND.n3351 GND.n3350 10.6151
R8201 GND.n3350 GND.n3204 10.6151
R8202 GND.n3345 GND.n3204 10.6151
R8203 GND.n3345 GND.n3344 10.6151
R8204 GND.n3344 GND.n3343 10.6151
R8205 GND.n3343 GND.n3206 10.6151
R8206 GND.n3337 GND.n3206 10.6151
R8207 GND.n3337 GND.n3336 10.6151
R8208 GND.n3336 GND.n3335 10.6151
R8209 GND.n3335 GND.n3208 10.6151
R8210 GND.n3329 GND.n3208 10.6151
R8211 GND.n3329 GND.n3328 10.6151
R8212 GND.n3328 GND.n3327 10.6151
R8213 GND.n3327 GND.n3210 10.6151
R8214 GND.n3321 GND.n3210 10.6151
R8215 GND.n3321 GND.n3320 10.6151
R8216 GND.n3320 GND.n3319 10.6151
R8217 GND.n3319 GND.n3212 10.6151
R8218 GND.n3313 GND.n3212 10.6151
R8219 GND.n3313 GND.n3312 10.6151
R8220 GND.n3312 GND.n3311 10.6151
R8221 GND.n3311 GND.n3214 10.6151
R8222 GND.n3305 GND.n3304 10.6151
R8223 GND.n3304 GND.n3303 10.6151
R8224 GND.n3891 GND.n3890 10.6151
R8225 GND.n3890 GND.n3889 10.6151
R8226 GND.n3889 GND.n3886 10.6151
R8227 GND.n3886 GND.n3885 10.6151
R8228 GND.n3885 GND.n3882 10.6151
R8229 GND.n3882 GND.n3881 10.6151
R8230 GND.n3881 GND.n3878 10.6151
R8231 GND.n3878 GND.n3877 10.6151
R8232 GND.n3877 GND.n3874 10.6151
R8233 GND.n3874 GND.n3873 10.6151
R8234 GND.n3873 GND.n3870 10.6151
R8235 GND.n3870 GND.n3869 10.6151
R8236 GND.n3869 GND.n3866 10.6151
R8237 GND.n3866 GND.n3865 10.6151
R8238 GND.n3865 GND.n3862 10.6151
R8239 GND.n3862 GND.n3861 10.6151
R8240 GND.n3861 GND.n3858 10.6151
R8241 GND.n3858 GND.n3857 10.6151
R8242 GND.n3857 GND.n3854 10.6151
R8243 GND.n3854 GND.n3853 10.6151
R8244 GND.n3853 GND.n3850 10.6151
R8245 GND.n3850 GND.n3849 10.6151
R8246 GND.n3849 GND.n3846 10.6151
R8247 GND.n3846 GND.n3845 10.6151
R8248 GND.n3845 GND.n3842 10.6151
R8249 GND.n3840 GND.n3837 10.6151
R8250 GND.n3837 GND.n3836 10.6151
R8251 GND.n3359 GND.n3144 10.6151
R8252 GND.n3501 GND.n3144 10.6151
R8253 GND.n3502 GND.n3501 10.6151
R8254 GND.n3503 GND.n3502 10.6151
R8255 GND.n3503 GND.n3131 10.6151
R8256 GND.n3520 GND.n3131 10.6151
R8257 GND.n3521 GND.n3520 10.6151
R8258 GND.n3522 GND.n3521 10.6151
R8259 GND.n3522 GND.n3115 10.6151
R8260 GND.n3543 GND.n3115 10.6151
R8261 GND.n3544 GND.n3543 10.6151
R8262 GND.n3545 GND.n3544 10.6151
R8263 GND.n3545 GND.n3099 10.6151
R8264 GND.n3576 GND.n3099 10.6151
R8265 GND.n3577 GND.n3576 10.6151
R8266 GND.n3578 GND.n3577 10.6151
R8267 GND.n3578 GND.n3094 10.6151
R8268 GND.n3595 GND.n3094 10.6151
R8269 GND.n3595 GND.n3594 10.6151
R8270 GND.n3594 GND.n3593 10.6151
R8271 GND.n3593 GND.n3077 10.6151
R8272 GND.n3647 GND.n3077 10.6151
R8273 GND.n3648 GND.n3647 10.6151
R8274 GND.n3652 GND.n3648 10.6151
R8275 GND.n3652 GND.n3651 10.6151
R8276 GND.n3651 GND.n3650 10.6151
R8277 GND.n3650 GND.n3055 10.6151
R8278 GND.n3678 GND.n3055 10.6151
R8279 GND.n3679 GND.n3678 10.6151
R8280 GND.n3680 GND.n3679 10.6151
R8281 GND.n3680 GND.n3040 10.6151
R8282 GND.n3703 GND.n3040 10.6151
R8283 GND.n3704 GND.n3703 10.6151
R8284 GND.n3705 GND.n3704 10.6151
R8285 GND.n3705 GND.n3025 10.6151
R8286 GND.n3724 GND.n3025 10.6151
R8287 GND.n3725 GND.n3724 10.6151
R8288 GND.n3726 GND.n3725 10.6151
R8289 GND.n3726 GND.n3014 10.6151
R8290 GND.n3747 GND.n3014 10.6151
R8291 GND.n3747 GND.n3746 10.6151
R8292 GND.n3746 GND.n3745 10.6151
R8293 GND.n3745 GND.n3015 10.6151
R8294 GND.n3015 GND.n2988 10.6151
R8295 GND.n3781 GND.n2988 10.6151
R8296 GND.n3782 GND.n3781 10.6151
R8297 GND.n3784 GND.n3782 10.6151
R8298 GND.n3784 GND.n3783 10.6151
R8299 GND.n3783 GND.n2904 10.6151
R8300 GND.n3813 GND.n2904 10.6151
R8301 GND.n3814 GND.n3813 10.6151
R8302 GND.n3815 GND.n3814 10.6151
R8303 GND.n3815 GND.n2891 10.6151
R8304 GND.n3829 GND.n2891 10.6151
R8305 GND.n3830 GND.n3829 10.6151
R8306 GND.n145 GND.n129 10.4732
R8307 GND.n113 GND.n97 10.4732
R8308 GND.n81 GND.n65 10.4732
R8309 GND.n50 GND.n34 10.4732
R8310 GND.n272 GND.n256 10.4732
R8311 GND.n240 GND.n224 10.4732
R8312 GND.n208 GND.n192 10.4732
R8313 GND.n177 GND.n161 10.4732
R8314 GND.n1948 GND.t25 10.3244
R8315 GND.n2053 GND.t141 10.3244
R8316 GND.n4270 GND.t151 10.3244
R8317 GND.t39 GND.n453 10.3244
R8318 GND.n3362 GND.n3361 9.99142
R8319 GND.n3637 GND.n3074 9.99142
R8320 GND.n3682 GND.n3053 9.99142
R8321 GND.n3896 GND.n2838 9.99142
R8322 GND.n3905 GND.t67 9.99142
R8323 GND.n149 GND.n148 9.69747
R8324 GND.n117 GND.n116 9.69747
R8325 GND.n85 GND.n84 9.69747
R8326 GND.n54 GND.n53 9.69747
R8327 GND.n276 GND.n275 9.69747
R8328 GND.n244 GND.n243 9.69747
R8329 GND.n212 GND.n211 9.69747
R8330 GND.n181 GND.n180 9.69747
R8331 GND.n2195 GND.t156 9.65839
R8332 GND.t123 GND.n2697 9.65839
R8333 GND.n155 GND.n154 9.45567
R8334 GND.n123 GND.n122 9.45567
R8335 GND.n91 GND.n90 9.45567
R8336 GND.n60 GND.n59 9.45567
R8337 GND.n282 GND.n281 9.45567
R8338 GND.n250 GND.n249 9.45567
R8339 GND.n218 GND.n217 9.45567
R8340 GND.n187 GND.n186 9.45567
R8341 GND.n3540 GND.n3111 9.32536
R8342 GND.n3590 GND.n3588 9.32536
R8343 GND.n3722 GND.n3027 9.32536
R8344 GND.n3737 GND.n2990 9.32536
R8345 GND.n971 GND.n970 9.3005
R8346 GND.n5034 GND.n5033 9.3005
R8347 GND.n5035 GND.n969 9.3005
R8348 GND.n5037 GND.n5036 9.3005
R8349 GND.n965 GND.n964 9.3005
R8350 GND.n5044 GND.n5043 9.3005
R8351 GND.n5045 GND.n963 9.3005
R8352 GND.n5047 GND.n5046 9.3005
R8353 GND.n959 GND.n958 9.3005
R8354 GND.n5054 GND.n5053 9.3005
R8355 GND.n5055 GND.n957 9.3005
R8356 GND.n5057 GND.n5056 9.3005
R8357 GND.n953 GND.n952 9.3005
R8358 GND.n5064 GND.n5063 9.3005
R8359 GND.n5065 GND.n951 9.3005
R8360 GND.n5067 GND.n5066 9.3005
R8361 GND.n947 GND.n946 9.3005
R8362 GND.n5074 GND.n5073 9.3005
R8363 GND.n5075 GND.n945 9.3005
R8364 GND.n5077 GND.n5076 9.3005
R8365 GND.n941 GND.n940 9.3005
R8366 GND.n5084 GND.n5083 9.3005
R8367 GND.n5085 GND.n939 9.3005
R8368 GND.n5087 GND.n5086 9.3005
R8369 GND.n935 GND.n934 9.3005
R8370 GND.n5094 GND.n5093 9.3005
R8371 GND.n5095 GND.n933 9.3005
R8372 GND.n5097 GND.n5096 9.3005
R8373 GND.n929 GND.n928 9.3005
R8374 GND.n5104 GND.n5103 9.3005
R8375 GND.n5105 GND.n927 9.3005
R8376 GND.n5107 GND.n5106 9.3005
R8377 GND.n923 GND.n922 9.3005
R8378 GND.n5114 GND.n5113 9.3005
R8379 GND.n5115 GND.n921 9.3005
R8380 GND.n5117 GND.n5116 9.3005
R8381 GND.n917 GND.n916 9.3005
R8382 GND.n5124 GND.n5123 9.3005
R8383 GND.n5125 GND.n915 9.3005
R8384 GND.n5127 GND.n5126 9.3005
R8385 GND.n911 GND.n910 9.3005
R8386 GND.n5134 GND.n5133 9.3005
R8387 GND.n5135 GND.n909 9.3005
R8388 GND.n5137 GND.n5136 9.3005
R8389 GND.n905 GND.n904 9.3005
R8390 GND.n5144 GND.n5143 9.3005
R8391 GND.n5145 GND.n903 9.3005
R8392 GND.n5147 GND.n5146 9.3005
R8393 GND.n899 GND.n898 9.3005
R8394 GND.n5154 GND.n5153 9.3005
R8395 GND.n5155 GND.n897 9.3005
R8396 GND.n5157 GND.n5156 9.3005
R8397 GND.n893 GND.n892 9.3005
R8398 GND.n5164 GND.n5163 9.3005
R8399 GND.n5165 GND.n891 9.3005
R8400 GND.n5167 GND.n5166 9.3005
R8401 GND.n887 GND.n886 9.3005
R8402 GND.n5174 GND.n5173 9.3005
R8403 GND.n5175 GND.n885 9.3005
R8404 GND.n5177 GND.n5176 9.3005
R8405 GND.n881 GND.n880 9.3005
R8406 GND.n5184 GND.n5183 9.3005
R8407 GND.n5185 GND.n879 9.3005
R8408 GND.n5187 GND.n5186 9.3005
R8409 GND.n875 GND.n874 9.3005
R8410 GND.n5194 GND.n5193 9.3005
R8411 GND.n5195 GND.n873 9.3005
R8412 GND.n5197 GND.n5196 9.3005
R8413 GND.n869 GND.n868 9.3005
R8414 GND.n5204 GND.n5203 9.3005
R8415 GND.n5205 GND.n867 9.3005
R8416 GND.n5207 GND.n5206 9.3005
R8417 GND.n863 GND.n862 9.3005
R8418 GND.n5214 GND.n5213 9.3005
R8419 GND.n5215 GND.n861 9.3005
R8420 GND.n5217 GND.n5216 9.3005
R8421 GND.n857 GND.n856 9.3005
R8422 GND.n5224 GND.n5223 9.3005
R8423 GND.n5225 GND.n855 9.3005
R8424 GND.n5227 GND.n5226 9.3005
R8425 GND.n851 GND.n850 9.3005
R8426 GND.n5234 GND.n5233 9.3005
R8427 GND.n5235 GND.n849 9.3005
R8428 GND.n5237 GND.n5236 9.3005
R8429 GND.n845 GND.n844 9.3005
R8430 GND.n5244 GND.n5243 9.3005
R8431 GND.n5245 GND.n843 9.3005
R8432 GND.n5247 GND.n5246 9.3005
R8433 GND.n839 GND.n838 9.3005
R8434 GND.n5254 GND.n5253 9.3005
R8435 GND.n5255 GND.n837 9.3005
R8436 GND.n5257 GND.n5256 9.3005
R8437 GND.n833 GND.n832 9.3005
R8438 GND.n5264 GND.n5263 9.3005
R8439 GND.n5265 GND.n831 9.3005
R8440 GND.n5267 GND.n5266 9.3005
R8441 GND.n827 GND.n826 9.3005
R8442 GND.n5274 GND.n5273 9.3005
R8443 GND.n5275 GND.n825 9.3005
R8444 GND.n5277 GND.n5276 9.3005
R8445 GND.n821 GND.n820 9.3005
R8446 GND.n5284 GND.n5283 9.3005
R8447 GND.n5285 GND.n819 9.3005
R8448 GND.n5287 GND.n5286 9.3005
R8449 GND.n815 GND.n814 9.3005
R8450 GND.n5294 GND.n5293 9.3005
R8451 GND.n5295 GND.n813 9.3005
R8452 GND.n5297 GND.n5296 9.3005
R8453 GND.n809 GND.n808 9.3005
R8454 GND.n5304 GND.n5303 9.3005
R8455 GND.n5305 GND.n807 9.3005
R8456 GND.n5307 GND.n5306 9.3005
R8457 GND.n803 GND.n802 9.3005
R8458 GND.n5314 GND.n5313 9.3005
R8459 GND.n5315 GND.n801 9.3005
R8460 GND.n5317 GND.n5316 9.3005
R8461 GND.n797 GND.n796 9.3005
R8462 GND.n5324 GND.n5323 9.3005
R8463 GND.n5325 GND.n795 9.3005
R8464 GND.n5327 GND.n5326 9.3005
R8465 GND.n791 GND.n790 9.3005
R8466 GND.n5334 GND.n5333 9.3005
R8467 GND.n5335 GND.n789 9.3005
R8468 GND.n5337 GND.n5336 9.3005
R8469 GND.n785 GND.n784 9.3005
R8470 GND.n5344 GND.n5343 9.3005
R8471 GND.n5345 GND.n783 9.3005
R8472 GND.n5347 GND.n5346 9.3005
R8473 GND.n779 GND.n778 9.3005
R8474 GND.n5354 GND.n5353 9.3005
R8475 GND.n5355 GND.n777 9.3005
R8476 GND.n5357 GND.n5356 9.3005
R8477 GND.n773 GND.n772 9.3005
R8478 GND.n5364 GND.n5363 9.3005
R8479 GND.n5365 GND.n771 9.3005
R8480 GND.n5367 GND.n5366 9.3005
R8481 GND.n767 GND.n766 9.3005
R8482 GND.n5374 GND.n5373 9.3005
R8483 GND.n5375 GND.n765 9.3005
R8484 GND.n5377 GND.n5376 9.3005
R8485 GND.n761 GND.n760 9.3005
R8486 GND.n5384 GND.n5383 9.3005
R8487 GND.n5385 GND.n759 9.3005
R8488 GND.n5387 GND.n5386 9.3005
R8489 GND.n755 GND.n754 9.3005
R8490 GND.n5394 GND.n5393 9.3005
R8491 GND.n5395 GND.n753 9.3005
R8492 GND.n5397 GND.n5396 9.3005
R8493 GND.n749 GND.n748 9.3005
R8494 GND.n5404 GND.n5403 9.3005
R8495 GND.n5405 GND.n747 9.3005
R8496 GND.n5407 GND.n5406 9.3005
R8497 GND.n743 GND.n742 9.3005
R8498 GND.n5414 GND.n5413 9.3005
R8499 GND.n5415 GND.n741 9.3005
R8500 GND.n5417 GND.n5416 9.3005
R8501 GND.n737 GND.n736 9.3005
R8502 GND.n5424 GND.n5423 9.3005
R8503 GND.n5425 GND.n735 9.3005
R8504 GND.n5427 GND.n5426 9.3005
R8505 GND.n731 GND.n730 9.3005
R8506 GND.n5434 GND.n5433 9.3005
R8507 GND.n5435 GND.n729 9.3005
R8508 GND.n5437 GND.n5436 9.3005
R8509 GND.n725 GND.n724 9.3005
R8510 GND.n5444 GND.n5443 9.3005
R8511 GND.n5445 GND.n723 9.3005
R8512 GND.n5447 GND.n5446 9.3005
R8513 GND.n719 GND.n718 9.3005
R8514 GND.n5454 GND.n5453 9.3005
R8515 GND.n5455 GND.n717 9.3005
R8516 GND.n5457 GND.n5456 9.3005
R8517 GND.n713 GND.n712 9.3005
R8518 GND.n5464 GND.n5463 9.3005
R8519 GND.n5465 GND.n711 9.3005
R8520 GND.n5467 GND.n5466 9.3005
R8521 GND.n707 GND.n706 9.3005
R8522 GND.n5474 GND.n5473 9.3005
R8523 GND.n5475 GND.n705 9.3005
R8524 GND.n5478 GND.n5476 9.3005
R8525 GND.n5477 GND.n701 9.3005
R8526 GND.n5486 GND.n700 9.3005
R8527 GND.n5488 GND.n5487 9.3005
R8528 GND.n696 GND.n695 9.3005
R8529 GND.n5495 GND.n5494 9.3005
R8530 GND.n5496 GND.n694 9.3005
R8531 GND.n5498 GND.n5497 9.3005
R8532 GND.n690 GND.n689 9.3005
R8533 GND.n5505 GND.n5504 9.3005
R8534 GND.n5506 GND.n688 9.3005
R8535 GND.n5508 GND.n5507 9.3005
R8536 GND.n684 GND.n683 9.3005
R8537 GND.n5515 GND.n5514 9.3005
R8538 GND.n5516 GND.n682 9.3005
R8539 GND.n5518 GND.n5517 9.3005
R8540 GND.n678 GND.n677 9.3005
R8541 GND.n5525 GND.n5524 9.3005
R8542 GND.n5526 GND.n676 9.3005
R8543 GND.n5528 GND.n5527 9.3005
R8544 GND.n672 GND.n671 9.3005
R8545 GND.n5535 GND.n5534 9.3005
R8546 GND.n5536 GND.n670 9.3005
R8547 GND.n5538 GND.n5537 9.3005
R8548 GND.n666 GND.n665 9.3005
R8549 GND.n5545 GND.n5544 9.3005
R8550 GND.n5546 GND.n664 9.3005
R8551 GND.n5548 GND.n5547 9.3005
R8552 GND.n660 GND.n659 9.3005
R8553 GND.n5555 GND.n5554 9.3005
R8554 GND.n5556 GND.n658 9.3005
R8555 GND.n5558 GND.n5557 9.3005
R8556 GND.n654 GND.n653 9.3005
R8557 GND.n5565 GND.n5564 9.3005
R8558 GND.n5566 GND.n652 9.3005
R8559 GND.n5568 GND.n5567 9.3005
R8560 GND.n648 GND.n647 9.3005
R8561 GND.n5575 GND.n5574 9.3005
R8562 GND.n5576 GND.n646 9.3005
R8563 GND.n5578 GND.n5577 9.3005
R8564 GND.n642 GND.n641 9.3005
R8565 GND.n5585 GND.n5584 9.3005
R8566 GND.n5586 GND.n640 9.3005
R8567 GND.n5588 GND.n5587 9.3005
R8568 GND.n636 GND.n635 9.3005
R8569 GND.n5595 GND.n5594 9.3005
R8570 GND.n5596 GND.n634 9.3005
R8571 GND.n5598 GND.n5597 9.3005
R8572 GND.n630 GND.n629 9.3005
R8573 GND.n5605 GND.n5604 9.3005
R8574 GND.n5606 GND.n628 9.3005
R8575 GND.n5608 GND.n5607 9.3005
R8576 GND.n624 GND.n623 9.3005
R8577 GND.n5615 GND.n5614 9.3005
R8578 GND.n5616 GND.n622 9.3005
R8579 GND.n5618 GND.n5617 9.3005
R8580 GND.n618 GND.n617 9.3005
R8581 GND.n5625 GND.n5624 9.3005
R8582 GND.n5626 GND.n616 9.3005
R8583 GND.n5628 GND.n5627 9.3005
R8584 GND.n612 GND.n611 9.3005
R8585 GND.n5635 GND.n5634 9.3005
R8586 GND.n5636 GND.n610 9.3005
R8587 GND.n5638 GND.n5637 9.3005
R8588 GND.n606 GND.n605 9.3005
R8589 GND.n5645 GND.n5644 9.3005
R8590 GND.n5646 GND.n604 9.3005
R8591 GND.n5649 GND.n5648 9.3005
R8592 GND.n5647 GND.n600 9.3005
R8593 GND.n5656 GND.n599 9.3005
R8594 GND.n5658 GND.n5657 9.3005
R8595 GND.n5485 GND.n5484 9.3005
R8596 GND.n3990 GND.n3987 9.3005
R8597 GND.n2781 GND.n2780 9.3005
R8598 GND.n4111 GND.n4110 9.3005
R8599 GND.n4112 GND.n2779 9.3005
R8600 GND.n4114 GND.n4113 9.3005
R8601 GND.n2777 GND.n2776 9.3005
R8602 GND.n4126 GND.n4125 9.3005
R8603 GND.n4127 GND.n2775 9.3005
R8604 GND.n4129 GND.n4128 9.3005
R8605 GND.n2773 GND.n2772 9.3005
R8606 GND.n4141 GND.n4140 9.3005
R8607 GND.n4142 GND.n2771 9.3005
R8608 GND.n4144 GND.n4143 9.3005
R8609 GND.n2768 GND.n2767 9.3005
R8610 GND.n4156 GND.n4155 9.3005
R8611 GND.n4157 GND.n2766 9.3005
R8612 GND.n4159 GND.n4158 9.3005
R8613 GND.n2764 GND.n2763 9.3005
R8614 GND.n4171 GND.n4170 9.3005
R8615 GND.n4172 GND.n2762 9.3005
R8616 GND.n4174 GND.n4173 9.3005
R8617 GND.n2760 GND.n2759 9.3005
R8618 GND.n4186 GND.n4185 9.3005
R8619 GND.n4187 GND.n2758 9.3005
R8620 GND.n4199 GND.n4188 9.3005
R8621 GND.n4198 GND.n4189 9.3005
R8622 GND.n4197 GND.n4190 9.3005
R8623 GND.n4196 GND.n4191 9.3005
R8624 GND.n4193 GND.n4192 9.3005
R8625 GND.n316 GND.n314 9.3005
R8626 GND.n3992 GND.n3991 9.3005
R8627 GND.n5921 GND.n5920 9.3005
R8628 GND.n317 GND.n315 9.3005
R8629 GND.n2749 GND.n2748 9.3005
R8630 GND.n4225 GND.n4224 9.3005
R8631 GND.n4226 GND.n2747 9.3005
R8632 GND.n4229 GND.n4228 9.3005
R8633 GND.n4227 GND.n2741 9.3005
R8634 GND.n4267 GND.n2742 9.3005
R8635 GND.n4266 GND.n2743 9.3005
R8636 GND.n4265 GND.n2744 9.3005
R8637 GND.n4240 GND.n2745 9.3005
R8638 GND.n4255 GND.n4241 9.3005
R8639 GND.n4254 GND.n4242 9.3005
R8640 GND.n4253 GND.n4243 9.3005
R8641 GND.n4248 GND.n4244 9.3005
R8642 GND.n4247 GND.n4246 9.3005
R8643 GND.n4245 GND.n586 9.3005
R8644 GND.n5701 GND.n585 9.3005
R8645 GND.n5703 GND.n5702 9.3005
R8646 GND.n5704 GND.n584 9.3005
R8647 GND.n5706 GND.n5705 9.3005
R8648 GND.n5708 GND.n583 9.3005
R8649 GND.n5710 GND.n5709 9.3005
R8650 GND.n5711 GND.n582 9.3005
R8651 GND.n5713 GND.n5712 9.3005
R8652 GND.n5715 GND.n580 9.3005
R8653 GND.n5717 GND.n5716 9.3005
R8654 GND.n5718 GND.n579 9.3005
R8655 GND.n5720 GND.n5719 9.3005
R8656 GND.n5722 GND.n577 9.3005
R8657 GND.n5724 GND.n5723 9.3005
R8658 GND.n5755 GND.n543 9.3005
R8659 GND.n5754 GND.n545 9.3005
R8660 GND.n549 GND.n546 9.3005
R8661 GND.n5749 GND.n550 9.3005
R8662 GND.n5748 GND.n551 9.3005
R8663 GND.n5747 GND.n552 9.3005
R8664 GND.n556 GND.n553 9.3005
R8665 GND.n5742 GND.n557 9.3005
R8666 GND.n5741 GND.n558 9.3005
R8667 GND.n5740 GND.n559 9.3005
R8668 GND.n563 GND.n560 9.3005
R8669 GND.n5735 GND.n564 9.3005
R8670 GND.n5734 GND.n565 9.3005
R8671 GND.n5733 GND.n566 9.3005
R8672 GND.n570 GND.n567 9.3005
R8673 GND.n5728 GND.n571 9.3005
R8674 GND.n5727 GND.n5726 9.3005
R8675 GND.n5725 GND.n574 9.3005
R8676 GND.n5757 GND.n5756 9.3005
R8677 GND.n5827 GND.n474 9.3005
R8678 GND.n5826 GND.n476 9.3005
R8679 GND.n480 GND.n477 9.3005
R8680 GND.n5821 GND.n481 9.3005
R8681 GND.n5820 GND.n482 9.3005
R8682 GND.n5819 GND.n483 9.3005
R8683 GND.n487 GND.n484 9.3005
R8684 GND.n5814 GND.n488 9.3005
R8685 GND.n5813 GND.n489 9.3005
R8686 GND.n5812 GND.n490 9.3005
R8687 GND.n494 GND.n491 9.3005
R8688 GND.n5807 GND.n495 9.3005
R8689 GND.n5806 GND.n496 9.3005
R8690 GND.n5805 GND.n497 9.3005
R8691 GND.n501 GND.n498 9.3005
R8692 GND.n5800 GND.n502 9.3005
R8693 GND.n5799 GND.n503 9.3005
R8694 GND.n5795 GND.n504 9.3005
R8695 GND.n508 GND.n505 9.3005
R8696 GND.n5790 GND.n509 9.3005
R8697 GND.n5789 GND.n510 9.3005
R8698 GND.n5788 GND.n511 9.3005
R8699 GND.n515 GND.n512 9.3005
R8700 GND.n5783 GND.n516 9.3005
R8701 GND.n5782 GND.n517 9.3005
R8702 GND.n5781 GND.n518 9.3005
R8703 GND.n522 GND.n519 9.3005
R8704 GND.n5776 GND.n523 9.3005
R8705 GND.n5775 GND.n524 9.3005
R8706 GND.n5774 GND.n525 9.3005
R8707 GND.n529 GND.n526 9.3005
R8708 GND.n5769 GND.n530 9.3005
R8709 GND.n5768 GND.n531 9.3005
R8710 GND.n5767 GND.n532 9.3005
R8711 GND.n536 GND.n533 9.3005
R8712 GND.n5762 GND.n537 9.3005
R8713 GND.n5761 GND.n5760 9.3005
R8714 GND.n5759 GND.n540 9.3005
R8715 GND.n5829 GND.n5828 9.3005
R8716 GND.n4404 GND.n4403 9.3005
R8717 GND.n2573 GND.n2572 9.3005
R8718 GND.n2597 GND.n2596 9.3005
R8719 GND.n4391 GND.n2598 9.3005
R8720 GND.n4390 GND.n2599 9.3005
R8721 GND.n4389 GND.n2600 9.3005
R8722 GND.n4120 GND.n2601 9.3005
R8723 GND.n4379 GND.n2619 9.3005
R8724 GND.n4378 GND.n2620 9.3005
R8725 GND.n4377 GND.n2621 9.3005
R8726 GND.n4135 GND.n2622 9.3005
R8727 GND.n4367 GND.n2640 9.3005
R8728 GND.n4366 GND.n2641 9.3005
R8729 GND.n4365 GND.n2642 9.3005
R8730 GND.n4150 GND.n2643 9.3005
R8731 GND.n4355 GND.n2660 9.3005
R8732 GND.n4354 GND.n2661 9.3005
R8733 GND.n4353 GND.n2662 9.3005
R8734 GND.n4165 GND.n2663 9.3005
R8735 GND.n4343 GND.n2681 9.3005
R8736 GND.n4342 GND.n2682 9.3005
R8737 GND.n4341 GND.n2683 9.3005
R8738 GND.n4180 GND.n2684 9.3005
R8739 GND.n4331 GND.n2702 9.3005
R8740 GND.n4330 GND.n2703 9.3005
R8741 GND.n4329 GND.n2704 9.3005
R8742 GND.n4206 GND.n2705 9.3005
R8743 GND.n4209 GND.n4208 9.3005
R8744 GND.n4210 GND.n2727 9.3005
R8745 GND.n4312 GND.n2728 9.3005
R8746 GND.n4311 GND.n2729 9.3005
R8747 GND.n4310 GND.n2730 9.3005
R8748 GND.n4218 GND.n2731 9.3005
R8749 GND.n4219 GND.n345 9.3005
R8750 GND.n5909 GND.n346 9.3005
R8751 GND.n5908 GND.n347 9.3005
R8752 GND.n5907 GND.n348 9.3005
R8753 GND.n4235 GND.n349 9.3005
R8754 GND.n5897 GND.n365 9.3005
R8755 GND.n5896 GND.n366 9.3005
R8756 GND.n5895 GND.n367 9.3005
R8757 GND.n4238 GND.n368 9.3005
R8758 GND.n5885 GND.n386 9.3005
R8759 GND.n5884 GND.n387 9.3005
R8760 GND.n5883 GND.n388 9.3005
R8761 GND.n588 GND.n389 9.3005
R8762 GND.n5873 GND.n406 9.3005
R8763 GND.n5872 GND.n407 9.3005
R8764 GND.n5871 GND.n408 9.3005
R8765 GND.n5673 GND.n409 9.3005
R8766 GND.n5861 GND.n426 9.3005
R8767 GND.n5860 GND.n427 9.3005
R8768 GND.n5859 GND.n428 9.3005
R8769 GND.n5674 GND.n429 9.3005
R8770 GND.n5849 GND.n446 9.3005
R8771 GND.n5848 GND.n447 9.3005
R8772 GND.n5847 GND.n448 9.3005
R8773 GND.n5675 GND.n449 9.3005
R8774 GND.n5837 GND.n465 9.3005
R8775 GND.n5836 GND.n466 9.3005
R8776 GND.n5835 GND.n467 9.3005
R8777 GND.n4405 GND.n2571 9.3005
R8778 GND.n4403 GND.n4402 9.3005
R8779 GND.n4401 GND.n2573 9.3005
R8780 GND.n2597 GND.n2574 9.3005
R8781 GND.n2778 GND.n2598 9.3005
R8782 GND.n4118 GND.n2599 9.3005
R8783 GND.n4119 GND.n2600 9.3005
R8784 GND.n4121 GND.n4120 9.3005
R8785 GND.n2774 GND.n2619 9.3005
R8786 GND.n4133 GND.n2620 9.3005
R8787 GND.n4134 GND.n2621 9.3005
R8788 GND.n4136 GND.n4135 9.3005
R8789 GND.n2770 GND.n2640 9.3005
R8790 GND.n4148 GND.n2641 9.3005
R8791 GND.n4149 GND.n2642 9.3005
R8792 GND.n4151 GND.n4150 9.3005
R8793 GND.n2765 GND.n2660 9.3005
R8794 GND.n4163 GND.n2661 9.3005
R8795 GND.n4164 GND.n2662 9.3005
R8796 GND.n4166 GND.n4165 9.3005
R8797 GND.n2761 GND.n2681 9.3005
R8798 GND.n4178 GND.n2682 9.3005
R8799 GND.n4179 GND.n2683 9.3005
R8800 GND.n4181 GND.n4180 9.3005
R8801 GND.n2757 GND.n2702 9.3005
R8802 GND.n4203 GND.n2703 9.3005
R8803 GND.n4204 GND.n2704 9.3005
R8804 GND.n4206 GND.n4205 9.3005
R8805 GND.n4209 GND.n2756 9.3005
R8806 GND.n4213 GND.n4210 9.3005
R8807 GND.n4214 GND.n2728 9.3005
R8808 GND.n4215 GND.n2729 9.3005
R8809 GND.n4216 GND.n2730 9.3005
R8810 GND.n4218 GND.n4217 9.3005
R8811 GND.n4220 GND.n4219 9.3005
R8812 GND.n2746 GND.n346 9.3005
R8813 GND.n4233 GND.n347 9.3005
R8814 GND.n4234 GND.n348 9.3005
R8815 GND.n4236 GND.n4235 9.3005
R8816 GND.n4237 GND.n365 9.3005
R8817 GND.n4261 GND.n366 9.3005
R8818 GND.n4260 GND.n367 9.3005
R8819 GND.n4259 GND.n4238 9.3005
R8820 GND.n4239 GND.n386 9.3005
R8821 GND.n4249 GND.n387 9.3005
R8822 GND.n587 GND.n388 9.3005
R8823 GND.n5671 GND.n588 9.3005
R8824 GND.n5672 GND.n406 9.3005
R8825 GND.n5697 GND.n407 9.3005
R8826 GND.n5696 GND.n408 9.3005
R8827 GND.n5695 GND.n5673 9.3005
R8828 GND.n5691 GND.n426 9.3005
R8829 GND.n5690 GND.n427 9.3005
R8830 GND.n5688 GND.n428 9.3005
R8831 GND.n5687 GND.n5674 9.3005
R8832 GND.n5685 GND.n446 9.3005
R8833 GND.n5684 GND.n447 9.3005
R8834 GND.n5682 GND.n448 9.3005
R8835 GND.n5681 GND.n5675 9.3005
R8836 GND.n5679 GND.n465 9.3005
R8837 GND.n5678 GND.n466 9.3005
R8838 GND.n5676 GND.n467 9.3005
R8839 GND.n2571 GND.n2565 9.3005
R8840 GND.n4414 GND.n4413 9.3005
R8841 GND.n4415 GND.n2558 9.3005
R8842 GND.n4418 GND.n2557 9.3005
R8843 GND.n4419 GND.n2556 9.3005
R8844 GND.n4422 GND.n2555 9.3005
R8845 GND.n4423 GND.n2554 9.3005
R8846 GND.n4426 GND.n2553 9.3005
R8847 GND.n4427 GND.n2552 9.3005
R8848 GND.n4430 GND.n2551 9.3005
R8849 GND.n4431 GND.n2550 9.3005
R8850 GND.n4434 GND.n2549 9.3005
R8851 GND.n4435 GND.n2548 9.3005
R8852 GND.n4438 GND.n2547 9.3005
R8853 GND.n4439 GND.n2546 9.3005
R8854 GND.n4442 GND.n2545 9.3005
R8855 GND.n4443 GND.n2544 9.3005
R8856 GND.n4446 GND.n2543 9.3005
R8857 GND.n4447 GND.n2542 9.3005
R8858 GND.n4450 GND.n2541 9.3005
R8859 GND.n4452 GND.n2535 9.3005
R8860 GND.n4455 GND.n2534 9.3005
R8861 GND.n4456 GND.n2533 9.3005
R8862 GND.n4459 GND.n2532 9.3005
R8863 GND.n4460 GND.n2531 9.3005
R8864 GND.n4463 GND.n2530 9.3005
R8865 GND.n4464 GND.n2529 9.3005
R8866 GND.n4467 GND.n2528 9.3005
R8867 GND.n4468 GND.n2527 9.3005
R8868 GND.n4471 GND.n2526 9.3005
R8869 GND.n4472 GND.n2525 9.3005
R8870 GND.n4475 GND.n2524 9.3005
R8871 GND.n4477 GND.n2523 9.3005
R8872 GND.n4478 GND.n2522 9.3005
R8873 GND.n4479 GND.n2521 9.3005
R8874 GND.n4480 GND.n2520 9.3005
R8875 GND.n4412 GND.n2563 9.3005
R8876 GND.n4411 GND.n4410 9.3005
R8877 GND.n2584 GND.n2581 9.3005
R8878 GND.n4397 GND.n2585 9.3005
R8879 GND.n4396 GND.n2586 9.3005
R8880 GND.n4395 GND.n2587 9.3005
R8881 GND.n2608 GND.n2588 9.3005
R8882 GND.n4385 GND.n2609 9.3005
R8883 GND.n4384 GND.n2610 9.3005
R8884 GND.n4383 GND.n2611 9.3005
R8885 GND.n2629 GND.n2612 9.3005
R8886 GND.n4373 GND.n2630 9.3005
R8887 GND.n4372 GND.n2631 9.3005
R8888 GND.n4371 GND.n2632 9.3005
R8889 GND.n2649 GND.n2633 9.3005
R8890 GND.n4361 GND.n2650 9.3005
R8891 GND.n4360 GND.n2651 9.3005
R8892 GND.n4359 GND.n2652 9.3005
R8893 GND.n2670 GND.n2653 9.3005
R8894 GND.n4349 GND.n2671 9.3005
R8895 GND.n4348 GND.n2672 9.3005
R8896 GND.n4347 GND.n2673 9.3005
R8897 GND.n2691 GND.n2674 9.3005
R8898 GND.n4337 GND.n2692 9.3005
R8899 GND.n4336 GND.n2693 9.3005
R8900 GND.n4335 GND.n2694 9.3005
R8901 GND.n2695 GND.n329 9.3005
R8902 GND.n336 GND.n328 9.3005
R8903 GND.n5903 GND.n355 9.3005
R8904 GND.n5902 GND.n356 9.3005
R8905 GND.n5901 GND.n357 9.3005
R8906 GND.n375 GND.n358 9.3005
R8907 GND.n5891 GND.n376 9.3005
R8908 GND.n5890 GND.n377 9.3005
R8909 GND.n5889 GND.n378 9.3005
R8910 GND.n396 GND.n379 9.3005
R8911 GND.n5879 GND.n397 9.3005
R8912 GND.n5878 GND.n398 9.3005
R8913 GND.n5877 GND.n399 9.3005
R8914 GND.n416 GND.n400 9.3005
R8915 GND.n5867 GND.n417 9.3005
R8916 GND.n5866 GND.n418 9.3005
R8917 GND.n5865 GND.n419 9.3005
R8918 GND.n436 GND.n420 9.3005
R8919 GND.n5855 GND.n437 9.3005
R8920 GND.n5854 GND.n438 9.3005
R8921 GND.n5853 GND.n439 9.3005
R8922 GND.n455 GND.n440 9.3005
R8923 GND.n5843 GND.n456 9.3005
R8924 GND.n5842 GND.n457 9.3005
R8925 GND.n5841 GND.n458 9.3005
R8926 GND.n473 GND.n459 9.3005
R8927 GND.n5831 GND.n5830 9.3005
R8928 GND.n2583 GND.n2582 9.3005
R8929 GND.n5914 GND.n333 9.3005
R8930 GND.n5914 GND.n5913 9.3005
R8931 GND.n2140 GND.n1506 9.3005
R8932 GND.n2193 GND.n2141 9.3005
R8933 GND.n2192 GND.n2142 9.3005
R8934 GND.n2191 GND.n2143 9.3005
R8935 GND.n2146 GND.n2144 9.3005
R8936 GND.n2187 GND.n2147 9.3005
R8937 GND.n2186 GND.n2148 9.3005
R8938 GND.n2185 GND.n2149 9.3005
R8939 GND.n2154 GND.n2150 9.3005
R8940 GND.n2181 GND.n2155 9.3005
R8941 GND.n2180 GND.n2156 9.3005
R8942 GND.n2179 GND.n2157 9.3005
R8943 GND.n2160 GND.n2158 9.3005
R8944 GND.n2175 GND.n2161 9.3005
R8945 GND.n2174 GND.n2162 9.3005
R8946 GND.n2173 GND.n2163 9.3005
R8947 GND.n2168 GND.n2164 9.3005
R8948 GND.n2167 GND.n2166 9.3005
R8949 GND.n2165 GND.n1427 9.3005
R8950 GND.n1425 GND.n1424 9.3005
R8951 GND.n2292 GND.n2291 9.3005
R8952 GND.n2293 GND.n1423 9.3005
R8953 GND.n2304 GND.n2294 9.3005
R8954 GND.n2303 GND.n2295 9.3005
R8955 GND.n2302 GND.n2296 9.3005
R8956 GND.n2299 GND.n2298 9.3005
R8957 GND.n2297 GND.n1309 9.3005
R8958 GND.n4708 GND.n1310 9.3005
R8959 GND.n4707 GND.n1311 9.3005
R8960 GND.n4706 GND.n1312 9.3005
R8961 GND.n3396 GND.n1313 9.3005
R8962 GND.n3398 GND.n3397 9.3005
R8963 GND.n3414 GND.n3413 9.3005
R8964 GND.n3415 GND.n3395 9.3005
R8965 GND.n3417 GND.n3416 9.3005
R8966 GND.n3385 GND.n3384 9.3005
R8967 GND.n3434 GND.n3433 9.3005
R8968 GND.n3435 GND.n3383 9.3005
R8969 GND.n3437 GND.n3436 9.3005
R8970 GND.n3372 GND.n3371 9.3005
R8971 GND.n3454 GND.n3453 9.3005
R8972 GND.n3455 GND.n3370 9.3005
R8973 GND.n3457 GND.n3456 9.3005
R8974 GND.n3176 GND.n3175 9.3005
R8975 GND.n3475 GND.n3474 9.3005
R8976 GND.n3476 GND.n3174 9.3005
R8977 GND.n3478 GND.n3477 9.3005
R8978 GND.n3139 GND.n3138 9.3005
R8979 GND.n3509 GND.n3508 9.3005
R8980 GND.n3510 GND.n3137 9.3005
R8981 GND.n3514 GND.n3511 9.3005
R8982 GND.n3513 GND.n3512 9.3005
R8983 GND.n3109 GND.n3108 9.3005
R8984 GND.n3551 GND.n3550 9.3005
R8985 GND.n3552 GND.n3107 9.3005
R8986 GND.n3571 GND.n3553 9.3005
R8987 GND.n3570 GND.n3554 9.3005
R8988 GND.n3569 GND.n3555 9.3005
R8989 GND.n3558 GND.n3556 9.3005
R8990 GND.n3565 GND.n3559 9.3005
R8991 GND.n3564 GND.n3560 9.3005
R8992 GND.n3563 GND.n3561 9.3005
R8993 GND.n3063 GND.n3062 9.3005
R8994 GND.n3667 GND.n3666 9.3005
R8995 GND.n3668 GND.n3061 9.3005
R8996 GND.n3672 GND.n3669 9.3005
R8997 GND.n3671 GND.n3670 9.3005
R8998 GND.n3034 GND.n3033 9.3005
R8999 GND.n3711 GND.n3710 9.3005
R9000 GND.n3712 GND.n3032 9.3005
R9001 GND.n3719 GND.n3713 9.3005
R9002 GND.n3718 GND.n3714 9.3005
R9003 GND.n3717 GND.n3715 9.3005
R9004 GND.n2998 GND.n2997 9.3005
R9005 GND.n3771 GND.n3770 9.3005
R9006 GND.n3772 GND.n2996 9.3005
R9007 GND.n3776 GND.n3773 9.3005
R9008 GND.n3775 GND.n3774 9.3005
R9009 GND.n2975 GND.n2974 9.3005
R9010 GND.n3796 GND.n3795 9.3005
R9011 GND.n3797 GND.n2973 9.3005
R9012 GND.n3799 GND.n3798 9.3005
R9013 GND.n2836 GND.n2835 9.3005
R9014 GND.n3899 GND.n3898 9.3005
R9015 GND.n3900 GND.n2834 9.3005
R9016 GND.n3902 GND.n3901 9.3005
R9017 GND.n2823 GND.n2822 9.3005
R9018 GND.n3918 GND.n3917 9.3005
R9019 GND.n3919 GND.n2821 9.3005
R9020 GND.n3921 GND.n3920 9.3005
R9021 GND.n2809 GND.n2808 9.3005
R9022 GND.n3937 GND.n3936 9.3005
R9023 GND.n3938 GND.n2807 9.3005
R9024 GND.n3942 GND.n3939 9.3005
R9025 GND.n3941 GND.n3940 9.3005
R9026 GND.n2795 GND.n2794 9.3005
R9027 GND.n3959 GND.n3958 9.3005
R9028 GND.n3960 GND.n2793 9.3005
R9029 GND.n3962 GND.n3961 9.3005
R9030 GND.n2790 GND.n2789 9.3005
R9031 GND.n4026 GND.n4025 9.3005
R9032 GND.n4027 GND.n2788 9.3005
R9033 GND.n4029 GND.n4028 9.3005
R9034 GND.n2786 GND.n2785 9.3005
R9035 GND.n4034 GND.n4033 9.3005
R9036 GND.n4035 GND.n2784 9.3005
R9037 GND.n4105 GND.n4036 9.3005
R9038 GND.n4104 GND.n4037 9.3005
R9039 GND.n4103 GND.n4038 9.3005
R9040 GND.n4041 GND.n4039 9.3005
R9041 GND.n4099 GND.n4042 9.3005
R9042 GND.n4098 GND.n4043 9.3005
R9043 GND.n4097 GND.n4044 9.3005
R9044 GND.n4047 GND.n4045 9.3005
R9045 GND.n4093 GND.n4048 9.3005
R9046 GND.n4092 GND.n4049 9.3005
R9047 GND.n4091 GND.n4050 9.3005
R9048 GND.n4053 GND.n4051 9.3005
R9049 GND.n4087 GND.n4054 9.3005
R9050 GND.n4086 GND.n4055 9.3005
R9051 GND.n4085 GND.n4056 9.3005
R9052 GND.n4059 GND.n4057 9.3005
R9053 GND.n4081 GND.n4060 9.3005
R9054 GND.n4080 GND.n4061 9.3005
R9055 GND.n4079 GND.n4062 9.3005
R9056 GND.n4065 GND.n4063 9.3005
R9057 GND.n4075 GND.n4066 9.3005
R9058 GND.n4074 GND.n4067 9.3005
R9059 GND.n4073 GND.n4068 9.3005
R9060 GND.n4272 GND.n2739 9.3005
R9061 GND.n4298 GND.n4273 9.3005
R9062 GND.n4297 GND.n4274 9.3005
R9063 GND.n4296 GND.n4275 9.3005
R9064 GND.n4278 GND.n4276 9.3005
R9065 GND.n4292 GND.n4279 9.3005
R9066 GND.n4291 GND.n4280 9.3005
R9067 GND.n4290 GND.n4281 9.3005
R9068 GND.n4283 GND.n4282 9.3005
R9069 GND.n4286 GND.n4285 9.3005
R9070 GND.n4284 GND.n592 9.3005
R9071 GND.n5666 GND.n593 9.3005
R9072 GND.n5665 GND.n594 9.3005
R9073 GND.n5664 GND.n595 9.3005
R9074 GND.n598 GND.n596 9.3005
R9075 GND.n5660 GND.n5659 9.3005
R9076 GND.n1842 GND.n1841 9.3005
R9077 GND.n1843 GND.n1756 9.3005
R9078 GND.n1844 GND.n1755 9.3005
R9079 GND.n1754 GND.n1752 9.3005
R9080 GND.n1850 GND.n1751 9.3005
R9081 GND.n1851 GND.n1750 9.3005
R9082 GND.n1852 GND.n1749 9.3005
R9083 GND.n1748 GND.n1746 9.3005
R9084 GND.n1858 GND.n1745 9.3005
R9085 GND.n1859 GND.n1744 9.3005
R9086 GND.n1860 GND.n1743 9.3005
R9087 GND.n1742 GND.n1740 9.3005
R9088 GND.n1866 GND.n1739 9.3005
R9089 GND.n1867 GND.n1738 9.3005
R9090 GND.n1868 GND.n1737 9.3005
R9091 GND.n1736 GND.n1734 9.3005
R9092 GND.n1874 GND.n1733 9.3005
R9093 GND.n1875 GND.n1732 9.3005
R9094 GND.n1876 GND.n1731 9.3005
R9095 GND.n1730 GND.n1725 9.3005
R9096 GND.n1882 GND.n1724 9.3005
R9097 GND.n1883 GND.n1723 9.3005
R9098 GND.n1884 GND.n1722 9.3005
R9099 GND.n1721 GND.n1719 9.3005
R9100 GND.n1890 GND.n1718 9.3005
R9101 GND.n1891 GND.n1717 9.3005
R9102 GND.n1892 GND.n1716 9.3005
R9103 GND.n1715 GND.n1713 9.3005
R9104 GND.n1898 GND.n1712 9.3005
R9105 GND.n1899 GND.n1711 9.3005
R9106 GND.n1900 GND.n1710 9.3005
R9107 GND.n1709 GND.n1707 9.3005
R9108 GND.n1905 GND.n1706 9.3005
R9109 GND.n1906 GND.n1705 9.3005
R9110 GND.n1704 GND.n1702 9.3005
R9111 GND.n1911 GND.n1701 9.3005
R9112 GND.n1913 GND.n1912 9.3005
R9113 GND.n1840 GND.n1761 9.3005
R9114 GND.n1839 GND.n1838 9.3005
R9115 GND.n1916 GND.n1915 9.3005
R9116 GND.n1676 GND.n1675 9.3005
R9117 GND.n1951 GND.n1950 9.3005
R9118 GND.n1952 GND.n1674 9.3005
R9119 GND.n1954 GND.n1953 9.3005
R9120 GND.n1657 GND.n1656 9.3005
R9121 GND.n1980 GND.n1979 9.3005
R9122 GND.n1981 GND.n1655 9.3005
R9123 GND.n1984 GND.n1983 9.3005
R9124 GND.n1982 GND.n1122 9.3005
R9125 GND.n4882 GND.n1123 9.3005
R9126 GND.n4881 GND.n1124 9.3005
R9127 GND.n4880 GND.n1125 9.3005
R9128 GND.n1634 GND.n1126 9.3005
R9129 GND.n1636 GND.n1635 9.3005
R9130 GND.n1613 GND.n1612 9.3005
R9131 GND.n2024 GND.n2023 9.3005
R9132 GND.n2025 GND.n1611 9.3005
R9133 GND.n2029 GND.n2026 9.3005
R9134 GND.n2028 GND.n2027 9.3005
R9135 GND.n1587 GND.n1586 9.3005
R9136 GND.n2061 GND.n2060 9.3005
R9137 GND.n2062 GND.n1585 9.3005
R9138 GND.n2065 GND.n2064 9.3005
R9139 GND.n2063 GND.n1525 9.3005
R9140 GND.n2098 GND.n2097 9.3005
R9141 GND.n1497 GND.n1496 9.3005
R9142 GND.n2205 GND.n2204 9.3005
R9143 GND.n2206 GND.n1495 9.3005
R9144 GND.n2210 GND.n2207 9.3005
R9145 GND.n2209 GND.n2208 9.3005
R9146 GND.n1474 GND.n1473 9.3005
R9147 GND.n2230 GND.n2229 9.3005
R9148 GND.n2231 GND.n1472 9.3005
R9149 GND.n2235 GND.n2232 9.3005
R9150 GND.n2234 GND.n2233 9.3005
R9151 GND.n1453 GND.n1452 9.3005
R9152 GND.n2254 GND.n2253 9.3005
R9153 GND.n2255 GND.n1451 9.3005
R9154 GND.n2259 GND.n2256 9.3005
R9155 GND.n2258 GND.n2257 9.3005
R9156 GND.n1432 GND.n1431 9.3005
R9157 GND.n2281 GND.n2280 9.3005
R9158 GND.n2282 GND.n1430 9.3005
R9159 GND.n2284 GND.n2283 9.3005
R9160 GND.n1408 GND.n1407 9.3005
R9161 GND.n2321 GND.n2320 9.3005
R9162 GND.n2322 GND.n1406 9.3005
R9163 GND.n2324 GND.n2323 9.3005
R9164 GND.n1243 GND.n1242 9.3005
R9165 GND.n4798 GND.n4797 9.3005
R9166 GND.n1917 GND.n1914 9.3005
R9167 GND.n2129 GND.n1511 9.3005
R9168 GND.n2096 GND.n1511 9.3005
R9169 GND.n1113 GND.n1112 9.3005
R9170 GND.n1628 GND.n1627 9.3005
R9171 GND.n1629 GND.n1625 9.3005
R9172 GND.n1631 GND.n1630 9.3005
R9173 GND.n1623 GND.n1622 9.3005
R9174 GND.n2010 GND.n2009 9.3005
R9175 GND.n2011 GND.n1621 9.3005
R9176 GND.n2015 GND.n2012 9.3005
R9177 GND.n2014 GND.n2013 9.3005
R9178 GND.n1596 GND.n1595 9.3005
R9179 GND.n2048 GND.n2047 9.3005
R9180 GND.n2049 GND.n1594 9.3005
R9181 GND.n2051 GND.n2050 9.3005
R9182 GND.n1514 GND.n1513 9.3005
R9183 GND.n2138 GND.n2137 9.3005
R9184 GND.n4888 GND.n4887 9.3005
R9185 GND.n4891 GND.n1111 9.3005
R9186 GND.n1110 GND.n1106 9.3005
R9187 GND.n4897 GND.n1105 9.3005
R9188 GND.n4898 GND.n1104 9.3005
R9189 GND.n4899 GND.n1103 9.3005
R9190 GND.n1102 GND.n1098 9.3005
R9191 GND.n4905 GND.n1097 9.3005
R9192 GND.n4906 GND.n1096 9.3005
R9193 GND.n4907 GND.n1095 9.3005
R9194 GND.n1094 GND.n1090 9.3005
R9195 GND.n4913 GND.n1089 9.3005
R9196 GND.n4914 GND.n1088 9.3005
R9197 GND.n4915 GND.n1087 9.3005
R9198 GND.n1086 GND.n1082 9.3005
R9199 GND.n4921 GND.n1081 9.3005
R9200 GND.n4922 GND.n1080 9.3005
R9201 GND.n4923 GND.n1079 9.3005
R9202 GND.n1078 GND.n1074 9.3005
R9203 GND.n4929 GND.n1073 9.3005
R9204 GND.n4930 GND.n1072 9.3005
R9205 GND.n4931 GND.n1071 9.3005
R9206 GND.n1070 GND.n1066 9.3005
R9207 GND.n4937 GND.n1065 9.3005
R9208 GND.n4938 GND.n1064 9.3005
R9209 GND.n4939 GND.n1063 9.3005
R9210 GND.n1062 GND.n1058 9.3005
R9211 GND.n4945 GND.n1057 9.3005
R9212 GND.n4946 GND.n1056 9.3005
R9213 GND.n4947 GND.n1055 9.3005
R9214 GND.n1054 GND.n1050 9.3005
R9215 GND.n4953 GND.n1049 9.3005
R9216 GND.n4954 GND.n1048 9.3005
R9217 GND.n4955 GND.n1047 9.3005
R9218 GND.n1046 GND.n1042 9.3005
R9219 GND.n4961 GND.n1041 9.3005
R9220 GND.n4962 GND.n1040 9.3005
R9221 GND.n4963 GND.n1039 9.3005
R9222 GND.n1038 GND.n1034 9.3005
R9223 GND.n4969 GND.n1033 9.3005
R9224 GND.n4970 GND.n1032 9.3005
R9225 GND.n4971 GND.n1031 9.3005
R9226 GND.n1030 GND.n1026 9.3005
R9227 GND.n4977 GND.n1025 9.3005
R9228 GND.n4978 GND.n1024 9.3005
R9229 GND.n4979 GND.n1023 9.3005
R9230 GND.n1022 GND.n1018 9.3005
R9231 GND.n4985 GND.n1017 9.3005
R9232 GND.n4986 GND.n1016 9.3005
R9233 GND.n4987 GND.n1015 9.3005
R9234 GND.n1014 GND.n1010 9.3005
R9235 GND.n4993 GND.n1009 9.3005
R9236 GND.n4994 GND.n1008 9.3005
R9237 GND.n4995 GND.n1007 9.3005
R9238 GND.n1006 GND.n1002 9.3005
R9239 GND.n5001 GND.n1001 9.3005
R9240 GND.n5002 GND.n1000 9.3005
R9241 GND.n5003 GND.n999 9.3005
R9242 GND.n998 GND.n994 9.3005
R9243 GND.n5009 GND.n993 9.3005
R9244 GND.n5010 GND.n992 9.3005
R9245 GND.n5011 GND.n991 9.3005
R9246 GND.n990 GND.n986 9.3005
R9247 GND.n5017 GND.n985 9.3005
R9248 GND.n5018 GND.n984 9.3005
R9249 GND.n5019 GND.n983 9.3005
R9250 GND.n982 GND.n978 9.3005
R9251 GND.n5025 GND.n977 9.3005
R9252 GND.n5026 GND.n976 9.3005
R9253 GND.n5027 GND.n975 9.3005
R9254 GND.n4890 GND.n4889 9.3005
R9255 GND.n3408 GND.n3407 9.3005
R9256 GND.n3392 GND.n3391 9.3005
R9257 GND.n3425 GND.n3424 9.3005
R9258 GND.n3426 GND.n3390 9.3005
R9259 GND.n3428 GND.n3427 9.3005
R9260 GND.n3379 GND.n3378 9.3005
R9261 GND.n3445 GND.n3444 9.3005
R9262 GND.n3446 GND.n3377 9.3005
R9263 GND.n3448 GND.n3447 9.3005
R9264 GND.n3366 GND.n3365 9.3005
R9265 GND.n3466 GND.n3465 9.3005
R9266 GND.n3467 GND.n3364 9.3005
R9267 GND.n3469 GND.n3468 9.3005
R9268 GND.n3170 GND.n3169 9.3005
R9269 GND.n3485 GND.n3484 9.3005
R9270 GND.n3486 GND.n3168 9.3005
R9271 GND.n3488 GND.n3487 9.3005
R9272 GND.n3124 GND.n3123 9.3005
R9273 GND.n3528 GND.n3527 9.3005
R9274 GND.n3529 GND.n3121 9.3005
R9275 GND.n3538 GND.n3537 9.3005
R9276 GND.n3536 GND.n3122 9.3005
R9277 GND.n3535 GND.n3534 9.3005
R9278 GND.n3533 GND.n3530 9.3005
R9279 GND.n3087 GND.n3086 9.3005
R9280 GND.n3601 GND.n3600 9.3005
R9281 GND.n3602 GND.n3085 9.3005
R9282 GND.n3604 GND.n3603 9.3005
R9283 GND.n3070 GND.n3069 9.3005
R9284 GND.n3658 GND.n3657 9.3005
R9285 GND.n3659 GND.n3068 9.3005
R9286 GND.n3661 GND.n3660 9.3005
R9287 GND.n3049 GND.n3048 9.3005
R9288 GND.n3686 GND.n3685 9.3005
R9289 GND.n3687 GND.n3046 9.3005
R9290 GND.n3698 GND.n3697 9.3005
R9291 GND.n3696 GND.n3047 9.3005
R9292 GND.n3695 GND.n3694 9.3005
R9293 GND.n3693 GND.n3688 9.3005
R9294 GND.n3007 GND.n3006 9.3005
R9295 GND.n3752 GND.n3751 9.3005
R9296 GND.n3753 GND.n3004 9.3005
R9297 GND.n3765 GND.n3764 9.3005
R9298 GND.n3763 GND.n3005 9.3005
R9299 GND.n3762 GND.n3761 9.3005
R9300 GND.n3760 GND.n3754 9.3005
R9301 GND.n3759 GND.n3758 9.3005
R9302 GND.n2899 GND.n2898 9.3005
R9303 GND.n3821 GND.n3820 9.3005
R9304 GND.n3822 GND.n2897 9.3005
R9305 GND.n3824 GND.n3823 9.3005
R9306 GND.n2830 GND.n2829 9.3005
R9307 GND.n3908 GND.n3907 9.3005
R9308 GND.n3909 GND.n2828 9.3005
R9309 GND.n3911 GND.n3910 9.3005
R9310 GND.n2816 GND.n2815 9.3005
R9311 GND.n3927 GND.n3926 9.3005
R9312 GND.n3928 GND.n2814 9.3005
R9313 GND.n3930 GND.n3929 9.3005
R9314 GND.n2801 GND.n2800 9.3005
R9315 GND.n3948 GND.n3947 9.3005
R9316 GND.n3949 GND.n2799 9.3005
R9317 GND.n3951 GND.n3950 9.3005
R9318 GND.n2433 GND.n2432 9.3005
R9319 GND.n4537 GND.n4536 9.3005
R9320 GND.n3406 GND.n3404 9.3005
R9321 GND.n4532 GND.n4531 9.3005
R9322 GND.n2438 GND.n2437 9.3005
R9323 GND.n4526 GND.n4525 9.3005
R9324 GND.n4524 GND.n4523 9.3005
R9325 GND.n2447 GND.n2446 9.3005
R9326 GND.n4518 GND.n4517 9.3005
R9327 GND.n4516 GND.n4515 9.3005
R9328 GND.n2455 GND.n2454 9.3005
R9329 GND.n4510 GND.n4509 9.3005
R9330 GND.n4508 GND.n4507 9.3005
R9331 GND.n2463 GND.n2462 9.3005
R9332 GND.n4502 GND.n4501 9.3005
R9333 GND.n4500 GND.n4499 9.3005
R9334 GND.n2471 GND.n2470 9.3005
R9335 GND.n4494 GND.n4493 9.3005
R9336 GND.n4492 GND.n4491 9.3005
R9337 GND.n2479 GND.n2478 9.3005
R9338 GND.n3997 GND.n3996 9.3005
R9339 GND.n4001 GND.n4000 9.3005
R9340 GND.n4002 GND.n3986 9.3005
R9341 GND.n4534 GND.n4533 9.3005
R9342 GND.n4490 GND.n4489 9.3005
R9343 GND.n2475 GND.n2474 9.3005
R9344 GND.n4496 GND.n4495 9.3005
R9345 GND.n4498 GND.n4497 9.3005
R9346 GND.n2467 GND.n2466 9.3005
R9347 GND.n4504 GND.n4503 9.3005
R9348 GND.n4506 GND.n4505 9.3005
R9349 GND.n2459 GND.n2458 9.3005
R9350 GND.n4512 GND.n4511 9.3005
R9351 GND.n4514 GND.n4513 9.3005
R9352 GND.n2451 GND.n2450 9.3005
R9353 GND.n4520 GND.n4519 9.3005
R9354 GND.n4522 GND.n4521 9.3005
R9355 GND.n2443 GND.n2442 9.3005
R9356 GND.n4528 GND.n4527 9.3005
R9357 GND.n4530 GND.n4529 9.3005
R9358 GND.n2439 GND.n2435 9.3005
R9359 GND.n4488 GND.n2482 9.3005
R9360 GND.n3993 GND.n2481 9.3005
R9361 GND.n4005 GND.n4004 9.3005
R9362 GND.n4008 GND.n3985 9.3005
R9363 GND.n4014 GND.n4013 9.3005
R9364 GND.n4015 GND.n3983 9.3005
R9365 GND.n4018 GND.n4017 9.3005
R9366 GND.n4016 GND.n3984 9.3005
R9367 GND.n4637 GND.n2344 9.3005
R9368 GND.n4636 GND.n4635 9.3005
R9369 GND.n4634 GND.n2349 9.3005
R9370 GND.n4633 GND.n4632 9.3005
R9371 GND.n4631 GND.n2350 9.3005
R9372 GND.n4630 GND.n4629 9.3005
R9373 GND.n4628 GND.n2354 9.3005
R9374 GND.n4627 GND.n4626 9.3005
R9375 GND.n4625 GND.n2355 9.3005
R9376 GND.n4624 GND.n4623 9.3005
R9377 GND.n4622 GND.n2359 9.3005
R9378 GND.n4621 GND.n4620 9.3005
R9379 GND.n4619 GND.n2360 9.3005
R9380 GND.n4618 GND.n4617 9.3005
R9381 GND.n4616 GND.n2364 9.3005
R9382 GND.n4615 GND.n4614 9.3005
R9383 GND.n4613 GND.n2365 9.3005
R9384 GND.n4612 GND.n4611 9.3005
R9385 GND.n4610 GND.n2369 9.3005
R9386 GND.n4609 GND.n4608 9.3005
R9387 GND.n4607 GND.n2370 9.3005
R9388 GND.n4606 GND.n4605 9.3005
R9389 GND.n4604 GND.n2374 9.3005
R9390 GND.n4603 GND.n4602 9.3005
R9391 GND.n4601 GND.n2375 9.3005
R9392 GND.n4600 GND.n4599 9.3005
R9393 GND.n4598 GND.n2379 9.3005
R9394 GND.n4597 GND.n4596 9.3005
R9395 GND.n4595 GND.n2380 9.3005
R9396 GND.n4594 GND.n4593 9.3005
R9397 GND.n4592 GND.n2384 9.3005
R9398 GND.n4591 GND.n4590 9.3005
R9399 GND.n4589 GND.n2385 9.3005
R9400 GND.n4588 GND.n4587 9.3005
R9401 GND.n4586 GND.n2389 9.3005
R9402 GND.n4585 GND.n4584 9.3005
R9403 GND.n4583 GND.n2390 9.3005
R9404 GND.n4582 GND.n4581 9.3005
R9405 GND.n4580 GND.n2394 9.3005
R9406 GND.n4579 GND.n4578 9.3005
R9407 GND.n4577 GND.n2395 9.3005
R9408 GND.n4576 GND.n4575 9.3005
R9409 GND.n4574 GND.n2399 9.3005
R9410 GND.n4573 GND.n4572 9.3005
R9411 GND.n4571 GND.n2400 9.3005
R9412 GND.n4570 GND.n4569 9.3005
R9413 GND.n4568 GND.n2404 9.3005
R9414 GND.n4567 GND.n4566 9.3005
R9415 GND.n4565 GND.n2405 9.3005
R9416 GND.n4564 GND.n4563 9.3005
R9417 GND.n4562 GND.n2409 9.3005
R9418 GND.n4561 GND.n4560 9.3005
R9419 GND.n4559 GND.n2410 9.3005
R9420 GND.n4558 GND.n4557 9.3005
R9421 GND.n4556 GND.n2414 9.3005
R9422 GND.n4555 GND.n4554 9.3005
R9423 GND.n4553 GND.n2415 9.3005
R9424 GND.n4552 GND.n4551 9.3005
R9425 GND.n4550 GND.n2419 9.3005
R9426 GND.n4549 GND.n4548 9.3005
R9427 GND.n4547 GND.n2420 9.3005
R9428 GND.n4546 GND.n4545 9.3005
R9429 GND.n4544 GND.n2424 9.3005
R9430 GND.n4543 GND.n4542 9.3005
R9431 GND.n4541 GND.n2425 9.3005
R9432 GND.n4639 GND.n4638 9.3005
R9433 GND.n4642 GND.n4641 9.3005
R9434 GND.n4643 GND.n2335 9.3005
R9435 GND.n4645 GND.n4644 9.3005
R9436 GND.n4646 GND.n1398 9.3005
R9437 GND.n4648 GND.n4647 9.3005
R9438 GND.n4640 GND.n2343 9.3005
R9439 GND.n2081 GND.n1565 9.3005
R9440 GND.n2083 GND.n2082 9.3005
R9441 GND.n2084 GND.n1564 9.3005
R9442 GND.n2086 GND.n2085 9.3005
R9443 GND.n2087 GND.n1562 9.3005
R9444 GND.n2092 GND.n2091 9.3005
R9445 GND.n2090 GND.n1563 9.3005
R9446 GND.n2089 GND.n2088 9.3005
R9447 GND.n1486 GND.n1485 9.3005
R9448 GND.n2215 GND.n2214 9.3005
R9449 GND.n2216 GND.n1483 9.3005
R9450 GND.n2219 GND.n2218 9.3005
R9451 GND.n2217 GND.n1484 9.3005
R9452 GND.n1465 GND.n1464 9.3005
R9453 GND.n2240 GND.n2239 9.3005
R9454 GND.n2241 GND.n1462 9.3005
R9455 GND.n2244 GND.n2243 9.3005
R9456 GND.n2242 GND.n1463 9.3005
R9457 GND.n1443 GND.n1442 9.3005
R9458 GND.n2264 GND.n2263 9.3005
R9459 GND.n2265 GND.n1440 9.3005
R9460 GND.n2271 GND.n2270 9.3005
R9461 GND.n2269 GND.n1441 9.3005
R9462 GND.n2268 GND.n2267 9.3005
R9463 GND.n1419 GND.n1417 9.3005
R9464 GND.n2313 GND.n2312 9.3005
R9465 GND.n2311 GND.n1418 9.3005
R9466 GND.n2310 GND.n2309 9.3005
R9467 GND.n1420 GND.n1400 9.3005
R9468 GND.n2331 GND.n1399 9.3005
R9469 GND.n2333 GND.n2332 9.3005
R9470 GND.n4697 GND.n4696 9.3005
R9471 GND.n4695 GND.n4694 9.3005
R9472 GND.n1340 GND.n1339 9.3005
R9473 GND.n4689 GND.n4688 9.3005
R9474 GND.n4687 GND.n4686 9.3005
R9475 GND.n1349 GND.n1348 9.3005
R9476 GND.n4681 GND.n4680 9.3005
R9477 GND.n4679 GND.n4678 9.3005
R9478 GND.n1359 GND.n1358 9.3005
R9479 GND.n4673 GND.n4672 9.3005
R9480 GND.n4671 GND.n4670 9.3005
R9481 GND.n1369 GND.n1368 9.3005
R9482 GND.n4665 GND.n4664 9.3005
R9483 GND.n4663 GND.n4662 9.3005
R9484 GND.n1379 GND.n1378 9.3005
R9485 GND.n4657 GND.n4656 9.3005
R9486 GND.n4655 GND.n1389 9.3005
R9487 GND.n4654 GND.n4652 9.3005
R9488 GND.n1335 GND.n1333 9.3005
R9489 GND.n4649 GND.n1392 9.3005
R9490 GND.n4651 GND.n4650 9.3005
R9491 GND.n1393 GND.n1391 9.3005
R9492 GND.n1385 GND.n1384 9.3005
R9493 GND.n4659 GND.n4658 9.3005
R9494 GND.n4661 GND.n4660 9.3005
R9495 GND.n1373 GND.n1372 9.3005
R9496 GND.n4667 GND.n4666 9.3005
R9497 GND.n4669 GND.n4668 9.3005
R9498 GND.n1365 GND.n1364 9.3005
R9499 GND.n4675 GND.n4674 9.3005
R9500 GND.n4677 GND.n4676 9.3005
R9501 GND.n1353 GND.n1352 9.3005
R9502 GND.n4683 GND.n4682 9.3005
R9503 GND.n4685 GND.n4684 9.3005
R9504 GND.n1345 GND.n1344 9.3005
R9505 GND.n4691 GND.n4690 9.3005
R9506 GND.n4693 GND.n4692 9.3005
R9507 GND.n1334 GND.n1332 9.3005
R9508 GND.n4699 GND.n4698 9.3005
R9509 GND.n4700 GND.n1331 9.3005
R9510 GND.n4773 GND.n1262 9.3005
R9511 GND.n4775 GND.n4774 9.3005
R9512 GND.n4776 GND.n1258 9.3005
R9513 GND.n4778 GND.n4777 9.3005
R9514 GND.n4779 GND.n1257 9.3005
R9515 GND.n4781 GND.n4780 9.3005
R9516 GND.n4782 GND.n1253 9.3005
R9517 GND.n4784 GND.n4783 9.3005
R9518 GND.n4785 GND.n1252 9.3005
R9519 GND.n4787 GND.n4786 9.3005
R9520 GND.n4788 GND.n1248 9.3005
R9521 GND.n4790 GND.n4789 9.3005
R9522 GND.n4791 GND.n1247 9.3005
R9523 GND.n4793 GND.n4792 9.3005
R9524 GND.n4794 GND.n1244 9.3005
R9525 GND.n4796 GND.n4795 9.3005
R9526 GND.n4769 GND.n4768 9.3005
R9527 GND.n4767 GND.n1270 9.3005
R9528 GND.n4766 GND.n4765 9.3005
R9529 GND.n4764 GND.n1271 9.3005
R9530 GND.n4763 GND.n4762 9.3005
R9531 GND.n4761 GND.n1275 9.3005
R9532 GND.n4760 GND.n4759 9.3005
R9533 GND.n4758 GND.n1276 9.3005
R9534 GND.n4757 GND.n4756 9.3005
R9535 GND.n4755 GND.n1280 9.3005
R9536 GND.n4754 GND.n4753 9.3005
R9537 GND.n4752 GND.n1281 9.3005
R9538 GND.n4751 GND.n4750 9.3005
R9539 GND.n4749 GND.n1285 9.3005
R9540 GND.n4748 GND.n4747 9.3005
R9541 GND.n4746 GND.n1286 9.3005
R9542 GND.n4745 GND.n4744 9.3005
R9543 GND.n4743 GND.n1290 9.3005
R9544 GND.n4742 GND.n4741 9.3005
R9545 GND.n4740 GND.n1291 9.3005
R9546 GND.n4770 GND.n1263 9.3005
R9547 GND.n1765 GND.n1764 9.3005
R9548 GND.n1684 GND.n1682 9.3005
R9549 GND.n1946 GND.n1945 9.3005
R9550 GND.n1687 GND.n1683 9.3005
R9551 GND.n1686 GND.n1685 9.3005
R9552 GND.n1666 GND.n1664 9.3005
R9553 GND.n1975 GND.n1974 9.3005
R9554 GND.n1667 GND.n1665 9.3005
R9555 GND.n1970 GND.n1963 9.3005
R9556 GND.n1969 GND.n1965 9.3005
R9557 GND.n1968 GND.n1966 9.3005
R9558 GND.n1136 GND.n1134 9.3005
R9559 GND.n4876 GND.n4875 9.3005
R9560 GND.n1137 GND.n1135 9.3005
R9561 GND.n4871 GND.n1142 9.3005
R9562 GND.n4870 GND.n1143 9.3005
R9563 GND.n4869 GND.n1144 9.3005
R9564 GND.n1619 GND.n1145 9.3005
R9565 GND.n4865 GND.n1150 9.3005
R9566 GND.n4864 GND.n1151 9.3005
R9567 GND.n4863 GND.n1152 9.3005
R9568 GND.n2056 GND.n1153 9.3005
R9569 GND.n4859 GND.n1158 9.3005
R9570 GND.n4858 GND.n1159 9.3005
R9571 GND.n4857 GND.n1160 9.3005
R9572 GND.n1521 GND.n1161 9.3005
R9573 GND.n4853 GND.n1166 9.3005
R9574 GND.n4852 GND.n1167 9.3005
R9575 GND.n4851 GND.n1168 9.3005
R9576 GND.n1532 GND.n1169 9.3005
R9577 GND.n4847 GND.n1174 9.3005
R9578 GND.n4846 GND.n1175 9.3005
R9579 GND.n4845 GND.n1176 9.3005
R9580 GND.n1555 GND.n1177 9.3005
R9581 GND.n4841 GND.n1182 9.3005
R9582 GND.n4840 GND.n1183 9.3005
R9583 GND.n4839 GND.n1184 9.3005
R9584 GND.n2200 GND.n1185 9.3005
R9585 GND.n4835 GND.n1190 9.3005
R9586 GND.n4834 GND.n1191 9.3005
R9587 GND.n4833 GND.n1192 9.3005
R9588 GND.n1480 GND.n1193 9.3005
R9589 GND.n4829 GND.n1198 9.3005
R9590 GND.n4828 GND.n1199 9.3005
R9591 GND.n4827 GND.n1200 9.3005
R9592 GND.n1459 GND.n1201 9.3005
R9593 GND.n4823 GND.n1206 9.3005
R9594 GND.n4822 GND.n1207 9.3005
R9595 GND.n4821 GND.n1208 9.3005
R9596 GND.n1447 GND.n1209 9.3005
R9597 GND.n4817 GND.n1214 9.3005
R9598 GND.n4816 GND.n1215 9.3005
R9599 GND.n4815 GND.n1216 9.3005
R9600 GND.n2275 GND.n1217 9.3005
R9601 GND.n4811 GND.n1222 9.3005
R9602 GND.n4810 GND.n1223 9.3005
R9603 GND.n4809 GND.n1224 9.3005
R9604 GND.n1403 GND.n1225 9.3005
R9605 GND.n4805 GND.n1230 9.3005
R9606 GND.n4804 GND.n1231 9.3005
R9607 GND.n4803 GND.n1232 9.3005
R9608 GND.n1767 GND.n1762 9.3005
R9609 GND.n1765 GND.n1688 9.3005
R9610 GND.n1942 GND.n1684 9.3005
R9611 GND.n1945 GND.n1944 9.3005
R9612 GND.n1943 GND.n1687 9.3005
R9613 GND.n1686 GND.n1668 9.3005
R9614 GND.n1959 GND.n1666 9.3005
R9615 GND.n1974 GND.n1973 9.3005
R9616 GND.n1972 GND.n1667 9.3005
R9617 GND.n1971 GND.n1970 9.3005
R9618 GND.n1969 GND.n1962 9.3005
R9619 GND.n1968 GND.n1967 9.3005
R9620 GND.n1138 GND.n1136 9.3005
R9621 GND.n4875 GND.n4874 9.3005
R9622 GND.n4873 GND.n1137 9.3005
R9623 GND.n4872 GND.n4871 9.3005
R9624 GND.n4870 GND.n1141 9.3005
R9625 GND.n4869 GND.n4868 9.3005
R9626 GND.n4867 GND.n1145 9.3005
R9627 GND.n4866 GND.n4865 9.3005
R9628 GND.n4864 GND.n1149 9.3005
R9629 GND.n4863 GND.n4862 9.3005
R9630 GND.n4861 GND.n1153 9.3005
R9631 GND.n4860 GND.n4859 9.3005
R9632 GND.n4858 GND.n1157 9.3005
R9633 GND.n4857 GND.n4856 9.3005
R9634 GND.n4855 GND.n1161 9.3005
R9635 GND.n4854 GND.n4853 9.3005
R9636 GND.n4852 GND.n1165 9.3005
R9637 GND.n4851 GND.n4850 9.3005
R9638 GND.n4849 GND.n1169 9.3005
R9639 GND.n4848 GND.n4847 9.3005
R9640 GND.n4846 GND.n1173 9.3005
R9641 GND.n4845 GND.n4844 9.3005
R9642 GND.n4843 GND.n1177 9.3005
R9643 GND.n4842 GND.n4841 9.3005
R9644 GND.n4840 GND.n1181 9.3005
R9645 GND.n4839 GND.n4838 9.3005
R9646 GND.n4837 GND.n1185 9.3005
R9647 GND.n4836 GND.n4835 9.3005
R9648 GND.n4834 GND.n1189 9.3005
R9649 GND.n4833 GND.n4832 9.3005
R9650 GND.n4831 GND.n1193 9.3005
R9651 GND.n4830 GND.n4829 9.3005
R9652 GND.n4828 GND.n1197 9.3005
R9653 GND.n4827 GND.n4826 9.3005
R9654 GND.n4825 GND.n1201 9.3005
R9655 GND.n4824 GND.n4823 9.3005
R9656 GND.n4822 GND.n1205 9.3005
R9657 GND.n4821 GND.n4820 9.3005
R9658 GND.n4819 GND.n1209 9.3005
R9659 GND.n4818 GND.n4817 9.3005
R9660 GND.n4816 GND.n1213 9.3005
R9661 GND.n4815 GND.n4814 9.3005
R9662 GND.n4813 GND.n1217 9.3005
R9663 GND.n4812 GND.n4811 9.3005
R9664 GND.n4810 GND.n1221 9.3005
R9665 GND.n4809 GND.n4808 9.3005
R9666 GND.n4807 GND.n1225 9.3005
R9667 GND.n4806 GND.n4805 9.3005
R9668 GND.n4804 GND.n1229 9.3005
R9669 GND.n4803 GND.n4802 9.3005
R9670 GND.n1767 GND.n1766 9.3005
R9671 GND.n1806 GND.n1805 9.3005
R9672 GND.n1807 GND.n1794 9.3005
R9673 GND.n1809 GND.n1808 9.3005
R9674 GND.n1810 GND.n1787 9.3005
R9675 GND.n1812 GND.n1811 9.3005
R9676 GND.n1813 GND.n1786 9.3005
R9677 GND.n1815 GND.n1814 9.3005
R9678 GND.n1816 GND.n1779 9.3005
R9679 GND.n1818 GND.n1817 9.3005
R9680 GND.n1819 GND.n1778 9.3005
R9681 GND.n1821 GND.n1820 9.3005
R9682 GND.n1822 GND.n1772 9.3005
R9683 GND.n1824 GND.n1823 9.3005
R9684 GND.n1825 GND.n1771 9.3005
R9685 GND.n1827 GND.n1826 9.3005
R9686 GND.n1769 GND.n1768 9.3005
R9687 GND.n1833 GND.n1832 9.3005
R9688 GND.n1804 GND.n1795 9.3005
R9689 GND.n1799 GND.n1694 9.3005
R9690 GND.n1923 GND.n1692 9.3005
R9691 GND.n1938 GND.n1937 9.3005
R9692 GND.n1936 GND.n1693 9.3005
R9693 GND.n1935 GND.n1934 9.3005
R9694 GND.n1933 GND.n1924 9.3005
R9695 GND.n1932 GND.n1931 9.3005
R9696 GND.n1930 GND.n1927 9.3005
R9697 GND.n1929 GND.n1928 9.3005
R9698 GND.n1649 GND.n1648 9.3005
R9699 GND.n1990 GND.n1989 9.3005
R9700 GND.n1991 GND.n1644 9.3005
R9701 GND.n1993 GND.n1992 9.3005
R9702 GND.n1994 GND.n1643 9.3005
R9703 GND.n1999 GND.n1998 9.3005
R9704 GND.n2000 GND.n1641 9.3005
R9705 GND.n2003 GND.n2002 9.3005
R9706 GND.n2001 GND.n1642 9.3005
R9707 GND.n1604 GND.n1603 9.3005
R9708 GND.n2034 GND.n2033 9.3005
R9709 GND.n2035 GND.n1601 9.3005
R9710 GND.n2041 GND.n2040 9.3005
R9711 GND.n2039 GND.n1602 9.3005
R9712 GND.n2038 GND.n2037 9.3005
R9713 GND.n2036 GND.n1578 9.3005
R9714 GND.n2070 GND.n1577 9.3005
R9715 GND.n2072 GND.n2071 9.3005
R9716 GND.n2073 GND.n1576 9.3005
R9717 GND.n2075 GND.n2074 9.3005
R9718 GND.n2076 GND.n1573 9.3005
R9719 GND.n2079 GND.n2078 9.3005
R9720 GND.n1922 GND.n1921 9.3005
R9721 GND.n154 GND.n153 9.3005
R9722 GND.n127 GND.n126 9.3005
R9723 GND.n148 GND.n147 9.3005
R9724 GND.n146 GND.n145 9.3005
R9725 GND.n131 GND.n130 9.3005
R9726 GND.n140 GND.n139 9.3005
R9727 GND.n138 GND.n137 9.3005
R9728 GND.n122 GND.n121 9.3005
R9729 GND.n95 GND.n94 9.3005
R9730 GND.n116 GND.n115 9.3005
R9731 GND.n114 GND.n113 9.3005
R9732 GND.n99 GND.n98 9.3005
R9733 GND.n108 GND.n107 9.3005
R9734 GND.n106 GND.n105 9.3005
R9735 GND.n90 GND.n89 9.3005
R9736 GND.n63 GND.n62 9.3005
R9737 GND.n84 GND.n83 9.3005
R9738 GND.n82 GND.n81 9.3005
R9739 GND.n67 GND.n66 9.3005
R9740 GND.n76 GND.n75 9.3005
R9741 GND.n74 GND.n73 9.3005
R9742 GND.n59 GND.n58 9.3005
R9743 GND.n32 GND.n31 9.3005
R9744 GND.n53 GND.n52 9.3005
R9745 GND.n51 GND.n50 9.3005
R9746 GND.n36 GND.n35 9.3005
R9747 GND.n45 GND.n44 9.3005
R9748 GND.n43 GND.n42 9.3005
R9749 GND.n281 GND.n280 9.3005
R9750 GND.n254 GND.n253 9.3005
R9751 GND.n275 GND.n274 9.3005
R9752 GND.n273 GND.n272 9.3005
R9753 GND.n258 GND.n257 9.3005
R9754 GND.n267 GND.n266 9.3005
R9755 GND.n265 GND.n264 9.3005
R9756 GND.n249 GND.n248 9.3005
R9757 GND.n222 GND.n221 9.3005
R9758 GND.n243 GND.n242 9.3005
R9759 GND.n241 GND.n240 9.3005
R9760 GND.n226 GND.n225 9.3005
R9761 GND.n235 GND.n234 9.3005
R9762 GND.n233 GND.n232 9.3005
R9763 GND.n217 GND.n216 9.3005
R9764 GND.n190 GND.n189 9.3005
R9765 GND.n211 GND.n210 9.3005
R9766 GND.n209 GND.n208 9.3005
R9767 GND.n194 GND.n193 9.3005
R9768 GND.n203 GND.n202 9.3005
R9769 GND.n201 GND.n200 9.3005
R9770 GND.n186 GND.n185 9.3005
R9771 GND.n159 GND.n158 9.3005
R9772 GND.n180 GND.n179 9.3005
R9773 GND.n178 GND.n177 9.3005
R9774 GND.n163 GND.n162 9.3005
R9775 GND.n172 GND.n171 9.3005
R9776 GND.n170 GND.n169 9.3005
R9777 GND.n2171 GND.t117 8.99233
R9778 GND.t134 GND.n2624 8.99233
R9779 GND.n152 GND.n127 8.92171
R9780 GND.n120 GND.n95 8.92171
R9781 GND.n88 GND.n63 8.92171
R9782 GND.n57 GND.n32 8.92171
R9783 GND.n279 GND.n254 8.92171
R9784 GND.n247 GND.n222 8.92171
R9785 GND.n215 GND.n190 8.92171
R9786 GND.n184 GND.n159 8.92171
R9787 GND.n2890 GND.n2872 8.72777
R9788 GND.n3524 GND.n3129 8.6593
R9789 GND.n3645 GND.n3079 8.6593
R9790 GND.n3708 GND.n3036 8.6593
R9791 GND.n3786 GND.n2982 8.6593
R9792 GND.t113 GND.n3643 8.32626
R9793 GND.n3701 GND.t109 8.32626
R9794 GND.n5923 GND.n5922 8.28706
R9795 GND.n2080 GND.n29 8.28706
R9796 GND.n153 GND.n125 8.14595
R9797 GND.n121 GND.n93 8.14595
R9798 GND.n89 GND.n61 8.14595
R9799 GND.n58 GND.n30 8.14595
R9800 GND.n280 GND.n252 8.14595
R9801 GND.n248 GND.n220 8.14595
R9802 GND.n216 GND.n188 8.14595
R9803 GND.n185 GND.n157 8.14595
R9804 GND.n3505 GND.t46 7.99323
R9805 GND.n3490 GND.t46 7.99323
R9806 GND.t8 GND.n3133 7.99323
R9807 GND.n3525 GND.n3524 7.99323
R9808 GND.n3581 GND.t92 7.99323
R9809 GND.n3645 GND.n3644 7.99323
R9810 GND.n3700 GND.n3036 7.99323
R9811 GND.t98 GND.n3729 7.99323
R9812 GND.n3786 GND.n2983 7.99323
R9813 GND.n4488 GND.n2481 7.75808
R9814 GND.n4655 GND.n4654 7.75808
R9815 GND.n1804 GND.n1799 7.75808
R9816 GND.n5727 GND.n574 7.75808
R9817 GND.n3548 GND.n3111 7.32717
R9818 GND.n3588 GND.n3091 7.32717
R9819 GND.n3722 GND.n3721 7.32717
R9820 GND.n3737 GND.n3736 7.32717
R9821 GND.n3793 GND.t22 7.32717
R9822 GND.n3817 GND.t5 7.32717
R9823 GND.n3200 GND.n3199 7.30353
R9824 GND.n2889 GND.n2888 7.30353
R9825 GND.n27 GND.n17 6.82809
R9826 GND.n303 GND.n293 6.82809
R9827 GND.n29 GND.n28 6.78875
R9828 GND.n5923 GND.n313 6.78875
R9829 GND.n4885 GND.n1115 6.66111
R9830 GND.n4884 GND.n1118 6.66111
R9831 GND.n1646 GND.n1128 6.66111
R9832 GND.n4878 GND.n1131 6.66111
R9833 GND.n2006 GND.n1638 6.66111
R9834 GND.n2005 GND.n1615 6.66111
R9835 GND.n2021 GND.n1617 6.66111
R9836 GND.n2018 GND.n2017 6.66111
R9837 GND.n2031 GND.n1606 6.66111
R9838 GND.n2044 GND.n1599 6.66111
R9839 GND.n2043 GND.n1589 6.66111
R9840 GND.n2058 GND.n1591 6.66111
R9841 GND.n2054 GND.n2053 6.66111
R9842 GND.n2067 GND.n1581 6.66111
R9843 GND.n2135 GND.n1518 6.66111
R9844 GND.n2134 GND.n1520 6.66111
R9845 GND.n1574 GND.n1528 6.66111
R9846 GND.n2124 GND.n2123 6.66111
R9847 GND.n2118 GND.n1536 6.66111
R9848 GND.n2117 GND.n1543 6.66111
R9849 GND.n1571 GND.n1570 6.66111
R9850 GND.n2110 GND.n1552 6.66111
R9851 GND.n2107 GND.n2106 6.66111
R9852 GND.n2101 GND.n1557 6.66111
R9853 GND.n2100 GND.n1502 6.66111
R9854 GND.n2196 GND.n2195 6.66111
R9855 GND.n2202 GND.n1500 6.66111
R9856 GND.n2198 GND.n1488 6.66111
R9857 GND.n2212 GND.n1490 6.66111
R9858 GND.n1493 GND.n1481 6.66111
R9859 GND.n2227 GND.n1478 6.66111
R9860 GND.n2224 GND.n1467 6.66111
R9861 GND.n2237 GND.n1468 6.66111
R9862 GND.n2152 GND.n2151 6.66111
R9863 GND.n2246 GND.n1455 6.66111
R9864 GND.n2251 GND.n1458 6.66111
R9865 GND.n2248 GND.n1445 6.66111
R9866 GND.n2261 GND.n1446 6.66111
R9867 GND.n2171 GND.n2170 6.66111
R9868 GND.n2273 GND.n1434 6.66111
R9869 GND.n2278 GND.n1436 6.66111
R9870 GND.n2287 GND.n1428 6.66111
R9871 GND.n2286 GND.n1414 6.66111
R9872 GND.n2315 GND.n1410 6.66111
R9873 GND.n2318 GND.n1412 6.66111
R9874 GND.n2307 GND.n2306 6.66111
R9875 GND.n2326 GND.n1402 6.66111
R9876 GND.n2329 GND.n1236 6.66111
R9877 GND.n4800 GND.n1238 6.66111
R9878 GND.n3361 GND.n3180 6.66111
R9879 GND.n3491 GND.n3490 6.66111
R9880 GND.n3637 GND.n3636 6.66111
R9881 GND.n3683 GND.n3682 6.66111
R9882 GND.n3811 GND.n3810 6.66111
R9883 GND.n4407 GND.n2566 6.66111
R9884 GND.n3988 GND.n2568 6.66111
R9885 GND.n4399 GND.n2576 6.66111
R9886 GND.n4108 GND.n4107 6.66111
R9887 GND.n4393 GND.n2590 6.66111
R9888 GND.n4116 GND.n2593 6.66111
R9889 GND.n4387 GND.n2603 6.66111
R9890 GND.n4123 GND.n2606 6.66111
R9891 GND.n4381 GND.n2614 6.66111
R9892 GND.n4131 GND.n2617 6.66111
R9893 GND.n4375 GND.n2624 6.66111
R9894 GND.n4138 GND.n2627 6.66111
R9895 GND.n4369 GND.n2635 6.66111
R9896 GND.n4146 GND.n2638 6.66111
R9897 GND.n4363 GND.n2645 6.66111
R9898 GND.n4153 GND.n2769 6.66111
R9899 GND.n4357 GND.n2655 6.66111
R9900 GND.n4161 GND.n2658 6.66111
R9901 GND.n4351 GND.n2665 6.66111
R9902 GND.n4345 GND.n2676 6.66111
R9903 GND.n4176 GND.n2679 6.66111
R9904 GND.n4339 GND.n2686 6.66111
R9905 GND.n4183 GND.n2689 6.66111
R9906 GND.n4333 GND.n2697 6.66111
R9907 GND.n4201 GND.n2700 6.66111
R9908 GND.n4327 GND.n2707 6.66111
R9909 GND.n4323 GND.n2710 6.66111
R9910 GND.n4322 GND.n2715 6.66111
R9911 GND.n2724 GND.n2721 6.66111
R9912 GND.n4315 GND.n4314 6.66111
R9913 GND.n5918 GND.n320 6.66111
R9914 GND.n4308 GND.n322 6.66111
R9915 GND.n4222 GND.n2751 6.66111
R9916 GND.n5911 GND.n339 6.66111
R9917 GND.n4231 GND.n342 6.66111
R9918 GND.n5905 GND.n351 6.66111
R9919 GND.n4270 GND.n4269 6.66111
R9920 GND.n5899 GND.n360 6.66111
R9921 GND.n4263 GND.n363 6.66111
R9922 GND.n5893 GND.n370 6.66111
R9923 GND.n4257 GND.n373 6.66111
R9924 GND.n5887 GND.n381 6.66111
R9925 GND.n4251 GND.n384 6.66111
R9926 GND.n5881 GND.n391 6.66111
R9927 GND.n5669 GND.n394 6.66111
R9928 GND.n5699 GND.n404 6.66111
R9929 GND.n5869 GND.n411 6.66111
R9930 GND.n5693 GND.n414 6.66111
R9931 GND.n5863 GND.n422 6.66111
R9932 GND.n2915 GND.n2910 6.5566
R9933 GND.n3293 GND.n3222 6.5566
R9934 GND.n3305 GND.n3218 6.5566
R9935 GND.n3841 GND.n3840 6.5566
R9936 GND.n1996 GND.t159 6.32808
R9937 GND.n2246 GND.t154 6.32808
R9938 GND.n3644 GND.t113 6.32808
R9939 GND.t109 GND.n3700 6.32808
R9940 GND.n4363 GND.t138 6.32808
R9941 GND.n5875 GND.t127 6.32808
R9942 GND.n5798 GND.n5795 6.20656
R9943 GND.n1876 GND.n1729 6.20656
R9944 GND.n3574 GND.n3573 5.99505
R9945 GND.n3580 GND.n3097 5.99505
R9946 GND.n3730 GND.n3009 5.99505
R9947 GND.n3018 GND.n3011 5.99505
R9948 GND.n155 GND.n125 5.81868
R9949 GND.n123 GND.n93 5.81868
R9950 GND.n91 GND.n61 5.81868
R9951 GND.n60 GND.n30 5.81868
R9952 GND.n282 GND.n252 5.81868
R9953 GND.n250 GND.n220 5.81868
R9954 GND.n218 GND.n188 5.81868
R9955 GND.n187 GND.n157 5.81868
R9956 GND.n2127 GND.t148 5.66202
R9957 GND.n2110 GND.t143 5.66202
R9958 GND.t103 GND.n3375 5.66202
R9959 GND.n3915 GND.t93 5.66202
R9960 GND.t129 GND.n2715 5.66202
R9961 GND.n2754 GND.t121 5.66202
R9962 GND.n2911 GND.n2536 5.62001
R9963 GND.n3295 GND.n1267 5.62001
R9964 GND.n3303 GND.n1267 5.62001
R9965 GND.n3836 GND.n2536 5.62001
R9966 GND.n4644 GND.n2338 5.4308
R9967 GND.n4013 GND.n4011 5.4308
R9968 GND.n3663 GND.n3066 5.32899
R9969 GND.n3676 GND.n3675 5.32899
R9970 GND.n3803 GND.n3802 5.32899
R9971 GND.t49 GND.n2838 5.32899
R9972 GND.n153 GND.n152 5.04292
R9973 GND.n121 GND.n120 5.04292
R9974 GND.n89 GND.n88 5.04292
R9975 GND.n58 GND.n57 5.04292
R9976 GND.n280 GND.n279 5.04292
R9977 GND.n248 GND.n247 5.04292
R9978 GND.n216 GND.n215 5.04292
R9979 GND.n185 GND.n184 5.04292
R9980 GND.n2031 GND.t162 4.99596
R9981 GND.n2221 GND.t136 4.99596
R9982 GND.n3893 GND.t67 4.99596
R9983 GND.n4168 GND.t132 4.99596
R9984 GND.n4257 GND.t115 4.99596
R9985 GND.n28 GND.n8 4.7699
R9986 GND.n313 GND.n312 4.7699
R9987 GND.n4325 GND.n334 4.74817
R9988 GND.n332 GND.n326 4.74817
R9989 GND.n5915 GND.n327 4.74817
R9990 GND.n335 GND.n331 4.74817
R9991 GND.n2712 GND.n334 4.74817
R9992 GND.n2722 GND.n332 4.74817
R9993 GND.n5916 GND.n5915 4.74817
R9994 GND.n2752 GND.n331 4.74817
R9995 GND.n1515 GND.n1512 4.74817
R9996 GND.n2121 GND.n1510 4.74817
R9997 GND.n1567 GND.n1509 4.74817
R9998 GND.n2103 GND.n1508 4.74817
R9999 GND.n1559 GND.n1507 4.74817
R10000 GND.n4069 GND.n2718 4.74817
R10001 GND.n4319 GND.n4318 4.74817
R10002 GND.n2736 GND.n2719 4.74817
R10003 GND.n4305 GND.n2738 4.74817
R10004 GND.n4303 GND.n4302 4.74817
R10005 GND.n4070 GND.n4069 4.74817
R10006 GND.n4320 GND.n4319 4.74817
R10007 GND.n4317 GND.n2719 4.74817
R10008 GND.n2738 GND.n2737 4.74817
R10009 GND.n4304 GND.n4303 4.74817
R10010 GND.n2132 GND.n2131 4.74817
R10011 GND.n1548 GND.n1547 4.74817
R10012 GND.n2114 GND.n2113 4.74817
R10013 GND.n2095 GND.n1549 4.74817
R10014 GND.n2131 GND.n2130 4.74817
R10015 GND.n1547 GND.n1526 4.74817
R10016 GND.n2115 GND.n2114 4.74817
R10017 GND.n2112 GND.n1549 4.74817
R10018 GND.n1538 GND.n1512 4.74817
R10019 GND.n1539 GND.n1510 4.74817
R10020 GND.n2120 GND.n1509 4.74817
R10021 GND.n1568 GND.n1508 4.74817
R10022 GND.n2104 GND.n1507 4.74817
R10023 GND.n27 GND.n26 4.7074
R10024 GND.n303 GND.n302 4.7074
R10025 GND.n3582 GND.n3089 4.66293
R10026 GND.n3728 GND.n3023 4.66293
R10027 GND.n4451 GND.n2538 4.6132
R10028 GND.n4772 GND.n4771 4.6132
R10029 GND.n2885 GND.n2872 4.46111
R10030 GND.n138 GND.n134 4.38594
R10031 GND.n106 GND.n102 4.38594
R10032 GND.n74 GND.n70 4.38594
R10033 GND.n43 GND.n39 4.38594
R10034 GND.n265 GND.n261 4.38594
R10035 GND.n233 GND.n229 4.38594
R10036 GND.n201 GND.n197 4.38594
R10037 GND.n170 GND.n166 4.38594
R10038 GND.n149 GND.n127 4.26717
R10039 GND.n117 GND.n95 4.26717
R10040 GND.n85 GND.n63 4.26717
R10041 GND.n54 GND.n32 4.26717
R10042 GND.n276 GND.n254 4.26717
R10043 GND.n244 GND.n222 4.26717
R10044 GND.n212 GND.n190 4.26717
R10045 GND.n181 GND.n159 4.26717
R10046 GND.n284 GND.n156 4.14478
R10047 GND.n2918 GND.n2910 4.05904
R10048 GND.n3289 GND.n3222 4.05904
R10049 GND.n3218 GND.n3214 4.05904
R10050 GND.n3842 GND.n3841 4.05904
R10051 GND.n3518 GND.n3517 3.99687
R10052 GND.n3792 GND.n2978 3.99687
R10053 GND.n3801 GND.t5 3.99687
R10054 GND.n2306 GND.t12 3.66384
R10055 GND.n3497 GND.t111 3.66384
R10056 GND.t107 GND.n3817 3.66384
R10057 GND.n4107 GND.t1 3.66384
R10058 GND.n284 GND.n283 3.60163
R10059 GND.n148 GND.n129 3.49141
R10060 GND.n116 GND.n97 3.49141
R10061 GND.n84 GND.n65 3.49141
R10062 GND.n53 GND.n34 3.49141
R10063 GND.n275 GND.n256 3.49141
R10064 GND.n243 GND.n224 3.49141
R10065 GND.n211 GND.n192 3.49141
R10066 GND.n180 GND.n161 3.49141
R10067 GND.n3482 GND.t64 3.33081
R10068 GND.n3541 GND.n3117 3.33081
R10069 GND.t99 GND.n3113 3.33081
R10070 GND.t100 GND.n3767 3.33081
R10071 GND.n3779 GND.n3778 3.33081
R10072 GND.n9 GND.t177 2.82907
R10073 GND.n9 GND.t155 2.82907
R10074 GND.n11 GND.t189 2.82907
R10075 GND.n11 GND.t157 2.82907
R10076 GND.n13 GND.t142 2.82907
R10077 GND.n13 GND.t186 2.82907
R10078 GND.n15 GND.t160 2.82907
R10079 GND.n15 GND.t163 2.82907
R10080 GND.n18 GND.t137 2.82907
R10081 GND.n18 GND.t180 2.82907
R10082 GND.n20 GND.t153 2.82907
R10083 GND.n20 GND.t181 2.82907
R10084 GND.n22 GND.t174 2.82907
R10085 GND.n22 GND.t149 2.82907
R10086 GND.n24 GND.t183 2.82907
R10087 GND.n24 GND.t187 2.82907
R10088 GND.n0 GND.t191 2.82907
R10089 GND.n0 GND.t161 2.82907
R10090 GND.n2 GND.t144 2.82907
R10091 GND.n2 GND.t190 2.82907
R10092 GND.n4 GND.t164 2.82907
R10093 GND.n4 GND.t185 2.82907
R10094 GND.n6 GND.t175 2.82907
R10095 GND.n6 GND.t194 2.82907
R10096 GND.n291 GND.t184 2.82907
R10097 GND.n291 GND.t128 2.82907
R10098 GND.n289 GND.t173 2.82907
R10099 GND.n289 GND.t188 2.82907
R10100 GND.n287 GND.t124 2.82907
R10101 GND.n287 GND.t176 2.82907
R10102 GND.n285 GND.t139 2.82907
R10103 GND.n285 GND.t133 2.82907
R10104 GND.n300 GND.t147 2.82907
R10105 GND.n300 GND.t167 2.82907
R10106 GND.n298 GND.t122 2.82907
R10107 GND.n298 GND.t152 2.82907
R10108 GND.n296 GND.t166 2.82907
R10109 GND.n296 GND.t130 2.82907
R10110 GND.n294 GND.t168 2.82907
R10111 GND.n294 GND.t165 2.82907
R10112 GND.n310 GND.t116 2.82907
R10113 GND.n310 GND.t171 2.82907
R10114 GND.n308 GND.t179 2.82907
R10115 GND.n308 GND.t158 2.82907
R10116 GND.n306 GND.t182 2.82907
R10117 GND.n306 GND.t140 2.82907
R10118 GND.n304 GND.t150 2.82907
R10119 GND.n304 GND.t193 2.82907
R10120 GND.n145 GND.n144 2.71565
R10121 GND.n113 GND.n112 2.71565
R10122 GND.n81 GND.n80 2.71565
R10123 GND.n50 GND.n49 2.71565
R10124 GND.n272 GND.n271 2.71565
R10125 GND.n240 GND.n239 2.71565
R10126 GND.n208 GND.n207 2.71565
R10127 GND.n177 GND.n176 2.71565
R10128 GND.t84 GND.n3516 2.66474
R10129 GND.n3160 GND.n3159 2.66474
R10130 GND.n3159 GND.t16 2.66474
R10131 GND.t92 GND.n3580 2.66474
R10132 GND.t195 GND.n3083 2.66474
R10133 GND.n3607 GND.n3606 2.66474
R10134 GND.n3655 GND.t95 2.66474
R10135 GND.t97 GND.n3624 2.66474
R10136 GND.n3707 GND.n3038 2.66474
R10137 GND.t96 GND.n3615 2.66474
R10138 GND.n3730 GND.t98 2.66474
R10139 GND.n2993 GND.n2992 2.66474
R10140 GND.n28 GND.n27 2.66322
R10141 GND.n313 GND.n303 2.66322
R10142 GND.t105 GND.n3151 2.33171
R10143 GND.n3152 GND.t105 2.33171
R10144 GND.n3743 GND.t101 2.33171
R10145 GND.n3768 GND.t101 2.33171
R10146 GND.n5914 GND.n334 2.27742
R10147 GND.n5914 GND.n332 2.27742
R10148 GND.n5915 GND.n5914 2.27742
R10149 GND.n5914 GND.n331 2.27742
R10150 GND.n4069 GND.n330 2.27742
R10151 GND.n4319 GND.n330 2.27742
R10152 GND.n2719 GND.n330 2.27742
R10153 GND.n2738 GND.n330 2.27742
R10154 GND.n4303 GND.n330 2.27742
R10155 GND.n2131 GND.n1511 2.27742
R10156 GND.n1547 GND.n1511 2.27742
R10157 GND.n2114 GND.n1511 2.27742
R10158 GND.n1549 GND.n1511 2.27742
R10159 GND.n2139 GND.n1512 2.27742
R10160 GND.n2139 GND.n1510 2.27742
R10161 GND.n2139 GND.n1509 2.27742
R10162 GND.n2139 GND.n1508 2.27742
R10163 GND.n2139 GND.n1507 2.27742
R10164 GND.t55 GND.n3362 1.99868
R10165 GND.n3499 GND.t64 1.99868
R10166 GND.n3491 GND.t8 1.99868
R10167 GND.n3516 GND.n3126 1.99868
R10168 GND.n3643 GND.n3072 1.99868
R10169 GND.n3701 GND.n3042 1.99868
R10170 GND.t74 GND.n2983 1.99868
R10171 GND.n2986 GND.n2985 1.99868
R10172 GND.n3811 GND.t29 1.99868
R10173 GND.n141 GND.n131 1.93989
R10174 GND.n109 GND.n99 1.93989
R10175 GND.n77 GND.n67 1.93989
R10176 GND.n46 GND.n36 1.93989
R10177 GND.n268 GND.n258 1.93989
R10178 GND.n236 GND.n226 1.93989
R10179 GND.n204 GND.n194 1.93989
R10180 GND.n173 GND.n163 1.93989
R10181 GND.t136 GND.n1476 1.66565
R10182 GND.n3472 GND.n3178 1.66565
R10183 GND.t111 GND.n3141 1.66565
R10184 GND.n3818 GND.t107 1.66565
R10185 GND.n3894 GND.n3893 1.66565
R10186 GND.t132 GND.n2668 1.66565
R10187 GND.n3547 GND.n3113 1.33262
R10188 GND.n3598 GND.n3597 1.33262
R10189 GND.t95 GND.n3654 1.33262
R10190 GND.n3625 GND.t97 1.33262
R10191 GND.n3691 GND.n3029 1.33262
R10192 GND.n3767 GND.n3001 1.33262
R10193 GND.n3826 GND.t49 1.33262
R10194 GND.n2338 GND.n1398 1.16414
R10195 GND.n4011 GND.n4008 1.16414
R10196 GND.n140 GND.n133 1.16414
R10197 GND.n108 GND.n101 1.16414
R10198 GND.n76 GND.n69 1.16414
R10199 GND.n45 GND.n38 1.16414
R10200 GND.n267 GND.n260 1.16414
R10201 GND.n235 GND.n228 1.16414
R10202 GND.n203 GND.n196 1.16414
R10203 GND.n172 GND.n165 1.16414
R10204 GND GND.n29 1.06897
R10205 GND.n17 GND.n16 1.00481
R10206 GND.n16 GND.n14 1.00481
R10207 GND.n14 GND.n12 1.00481
R10208 GND.n12 GND.n10 1.00481
R10209 GND.n26 GND.n25 1.00481
R10210 GND.n25 GND.n23 1.00481
R10211 GND.n23 GND.n21 1.00481
R10212 GND.n21 GND.n19 1.00481
R10213 GND.n8 GND.n7 1.00481
R10214 GND.n7 GND.n5 1.00481
R10215 GND.n5 GND.n3 1.00481
R10216 GND.n3 GND.n1 1.00481
R10217 GND.n288 GND.n286 1.00481
R10218 GND.n290 GND.n288 1.00481
R10219 GND.n292 GND.n290 1.00481
R10220 GND.n293 GND.n292 1.00481
R10221 GND.n297 GND.n295 1.00481
R10222 GND.n299 GND.n297 1.00481
R10223 GND.n301 GND.n299 1.00481
R10224 GND.n302 GND.n301 1.00481
R10225 GND.n307 GND.n305 1.00481
R10226 GND.n309 GND.n307 1.00481
R10227 GND.n311 GND.n309 1.00481
R10228 GND.n312 GND.n311 1.00481
R10229 GND.n1534 GND.t148 0.999592
R10230 GND.n4307 GND.t121 0.999592
R10231 GND.n4771 GND.n4770 0.970197
R10232 GND.n4451 GND.n4450 0.970197
R10233 GND.n124 GND.n92 0.962709
R10234 GND.n156 GND.n124 0.962709
R10235 GND.n251 GND.n219 0.962709
R10236 GND.n283 GND.n251 0.962709
R10237 GND.n3480 GND.n3172 0.666561
R10238 GND.n3506 GND.n3505 0.666561
R10239 GND.n3591 GND.t195 0.666561
R10240 GND.n3664 GND.n3065 0.666561
R10241 GND.n3674 GND.n3051 0.666561
R10242 GND.n3616 GND.t96 0.666561
R10243 GND.t22 GND.t29 0.666561
R10244 GND.n3809 GND.n2901 0.666561
R10245 GND.n3827 GND.n2893 0.666561
R10246 GND.n5924 GND.n5923 0.647847
R10247 GND.n5914 GND.n330 0.532625
R10248 GND.n2139 GND.n1511 0.532625
R10249 GND.n5725 GND.n5724 0.508122
R10250 GND.n1922 GND.n1694 0.508122
R10251 GND.n975 GND.n970 0.505073
R10252 GND.n5485 GND.n701 0.505073
R10253 GND.n5659 GND.n5658 0.505073
R10254 GND.n4889 GND.n4888 0.505073
R10255 GND.n5830 GND.n5829 0.495927
R10256 GND.n2583 GND.n2520 0.495927
R10257 GND.n4797 GND.n4796 0.495927
R10258 GND.n1914 GND.n1913 0.495927
R10259 GND.n4016 GND.n2425 0.48678
R10260 GND.n4640 GND.n4639 0.48678
R10261 GND.n5799 GND.n5798 0.388379
R10262 GND.n1729 GND.n1725 0.388379
R10263 GND.n137 GND.n136 0.388379
R10264 GND.n105 GND.n104 0.388379
R10265 GND.n73 GND.n72 0.388379
R10266 GND.n42 GND.n41 0.388379
R10267 GND.n264 GND.n263 0.388379
R10268 GND.n232 GND.n231 0.388379
R10269 GND.n200 GND.n199 0.388379
R10270 GND.n169 GND.n168 0.388379
R10271 GND.n5924 GND.n284 0.341877
R10272 GND.n3406 GND.n3405 0.338915
R10273 GND.n4536 GND.n4535 0.338915
R10274 GND.t159 GND.n1995 0.333531
R10275 GND.n3419 GND.t70 0.333531
R10276 GND.n2804 GND.t80 0.333531
R10277 GND.n5668 GND.t127 0.333531
R10278 GND.n5758 GND.n5757 0.293183
R10279 GND.n1834 GND.n1833 0.293183
R10280 GND.n5759 GND.n5758 0.280988
R10281 GND.n4411 GND.n2434 0.280988
R10282 GND.n1839 GND.n1834 0.280988
R10283 GND.n1291 GND.n1233 0.280988
R10284 GND.n4003 GND.n3992 0.277939
R10285 GND.n2334 GND.n2333 0.277939
R10286 GND.n2538 GND.n2535 0.229039
R10287 GND.n2541 GND.n2538 0.229039
R10288 GND.n4773 GND.n4772 0.229039
R10289 GND.n4772 GND.n1263 0.229039
R10290 GND GND.n5924 0.213018
R10291 GND.n154 GND.n126 0.155672
R10292 GND.n147 GND.n126 0.155672
R10293 GND.n147 GND.n146 0.155672
R10294 GND.n146 GND.n130 0.155672
R10295 GND.n139 GND.n130 0.155672
R10296 GND.n139 GND.n138 0.155672
R10297 GND.n122 GND.n94 0.155672
R10298 GND.n115 GND.n94 0.155672
R10299 GND.n115 GND.n114 0.155672
R10300 GND.n114 GND.n98 0.155672
R10301 GND.n107 GND.n98 0.155672
R10302 GND.n107 GND.n106 0.155672
R10303 GND.n90 GND.n62 0.155672
R10304 GND.n83 GND.n62 0.155672
R10305 GND.n83 GND.n82 0.155672
R10306 GND.n82 GND.n66 0.155672
R10307 GND.n75 GND.n66 0.155672
R10308 GND.n75 GND.n74 0.155672
R10309 GND.n59 GND.n31 0.155672
R10310 GND.n52 GND.n31 0.155672
R10311 GND.n52 GND.n51 0.155672
R10312 GND.n51 GND.n35 0.155672
R10313 GND.n44 GND.n35 0.155672
R10314 GND.n44 GND.n43 0.155672
R10315 GND.n281 GND.n253 0.155672
R10316 GND.n274 GND.n253 0.155672
R10317 GND.n274 GND.n273 0.155672
R10318 GND.n273 GND.n257 0.155672
R10319 GND.n266 GND.n257 0.155672
R10320 GND.n266 GND.n265 0.155672
R10321 GND.n249 GND.n221 0.155672
R10322 GND.n242 GND.n221 0.155672
R10323 GND.n242 GND.n241 0.155672
R10324 GND.n241 GND.n225 0.155672
R10325 GND.n234 GND.n225 0.155672
R10326 GND.n234 GND.n233 0.155672
R10327 GND.n217 GND.n189 0.155672
R10328 GND.n210 GND.n189 0.155672
R10329 GND.n210 GND.n209 0.155672
R10330 GND.n209 GND.n193 0.155672
R10331 GND.n202 GND.n193 0.155672
R10332 GND.n202 GND.n201 0.155672
R10333 GND.n186 GND.n158 0.155672
R10334 GND.n179 GND.n158 0.155672
R10335 GND.n179 GND.n178 0.155672
R10336 GND.n178 GND.n162 0.155672
R10337 GND.n171 GND.n162 0.155672
R10338 GND.n171 GND.n170 0.155672
R10339 GND.n5034 GND.n970 0.152939
R10340 GND.n5035 GND.n5034 0.152939
R10341 GND.n5036 GND.n5035 0.152939
R10342 GND.n5036 GND.n964 0.152939
R10343 GND.n5044 GND.n964 0.152939
R10344 GND.n5045 GND.n5044 0.152939
R10345 GND.n5046 GND.n5045 0.152939
R10346 GND.n5046 GND.n958 0.152939
R10347 GND.n5054 GND.n958 0.152939
R10348 GND.n5055 GND.n5054 0.152939
R10349 GND.n5056 GND.n5055 0.152939
R10350 GND.n5056 GND.n952 0.152939
R10351 GND.n5064 GND.n952 0.152939
R10352 GND.n5065 GND.n5064 0.152939
R10353 GND.n5066 GND.n5065 0.152939
R10354 GND.n5066 GND.n946 0.152939
R10355 GND.n5074 GND.n946 0.152939
R10356 GND.n5075 GND.n5074 0.152939
R10357 GND.n5076 GND.n5075 0.152939
R10358 GND.n5076 GND.n940 0.152939
R10359 GND.n5084 GND.n940 0.152939
R10360 GND.n5085 GND.n5084 0.152939
R10361 GND.n5086 GND.n5085 0.152939
R10362 GND.n5086 GND.n934 0.152939
R10363 GND.n5094 GND.n934 0.152939
R10364 GND.n5095 GND.n5094 0.152939
R10365 GND.n5096 GND.n5095 0.152939
R10366 GND.n5096 GND.n928 0.152939
R10367 GND.n5104 GND.n928 0.152939
R10368 GND.n5105 GND.n5104 0.152939
R10369 GND.n5106 GND.n5105 0.152939
R10370 GND.n5106 GND.n922 0.152939
R10371 GND.n5114 GND.n922 0.152939
R10372 GND.n5115 GND.n5114 0.152939
R10373 GND.n5116 GND.n5115 0.152939
R10374 GND.n5116 GND.n916 0.152939
R10375 GND.n5124 GND.n916 0.152939
R10376 GND.n5125 GND.n5124 0.152939
R10377 GND.n5126 GND.n5125 0.152939
R10378 GND.n5126 GND.n910 0.152939
R10379 GND.n5134 GND.n910 0.152939
R10380 GND.n5135 GND.n5134 0.152939
R10381 GND.n5136 GND.n5135 0.152939
R10382 GND.n5136 GND.n904 0.152939
R10383 GND.n5144 GND.n904 0.152939
R10384 GND.n5145 GND.n5144 0.152939
R10385 GND.n5146 GND.n5145 0.152939
R10386 GND.n5146 GND.n898 0.152939
R10387 GND.n5154 GND.n898 0.152939
R10388 GND.n5155 GND.n5154 0.152939
R10389 GND.n5156 GND.n5155 0.152939
R10390 GND.n5156 GND.n892 0.152939
R10391 GND.n5164 GND.n892 0.152939
R10392 GND.n5165 GND.n5164 0.152939
R10393 GND.n5166 GND.n5165 0.152939
R10394 GND.n5166 GND.n886 0.152939
R10395 GND.n5174 GND.n886 0.152939
R10396 GND.n5175 GND.n5174 0.152939
R10397 GND.n5176 GND.n5175 0.152939
R10398 GND.n5176 GND.n880 0.152939
R10399 GND.n5184 GND.n880 0.152939
R10400 GND.n5185 GND.n5184 0.152939
R10401 GND.n5186 GND.n5185 0.152939
R10402 GND.n5186 GND.n874 0.152939
R10403 GND.n5194 GND.n874 0.152939
R10404 GND.n5195 GND.n5194 0.152939
R10405 GND.n5196 GND.n5195 0.152939
R10406 GND.n5196 GND.n868 0.152939
R10407 GND.n5204 GND.n868 0.152939
R10408 GND.n5205 GND.n5204 0.152939
R10409 GND.n5206 GND.n5205 0.152939
R10410 GND.n5206 GND.n862 0.152939
R10411 GND.n5214 GND.n862 0.152939
R10412 GND.n5215 GND.n5214 0.152939
R10413 GND.n5216 GND.n5215 0.152939
R10414 GND.n5216 GND.n856 0.152939
R10415 GND.n5224 GND.n856 0.152939
R10416 GND.n5225 GND.n5224 0.152939
R10417 GND.n5226 GND.n5225 0.152939
R10418 GND.n5226 GND.n850 0.152939
R10419 GND.n5234 GND.n850 0.152939
R10420 GND.n5235 GND.n5234 0.152939
R10421 GND.n5236 GND.n5235 0.152939
R10422 GND.n5236 GND.n844 0.152939
R10423 GND.n5244 GND.n844 0.152939
R10424 GND.n5245 GND.n5244 0.152939
R10425 GND.n5246 GND.n5245 0.152939
R10426 GND.n5246 GND.n838 0.152939
R10427 GND.n5254 GND.n838 0.152939
R10428 GND.n5255 GND.n5254 0.152939
R10429 GND.n5256 GND.n5255 0.152939
R10430 GND.n5256 GND.n832 0.152939
R10431 GND.n5264 GND.n832 0.152939
R10432 GND.n5265 GND.n5264 0.152939
R10433 GND.n5266 GND.n5265 0.152939
R10434 GND.n5266 GND.n826 0.152939
R10435 GND.n5274 GND.n826 0.152939
R10436 GND.n5275 GND.n5274 0.152939
R10437 GND.n5276 GND.n5275 0.152939
R10438 GND.n5276 GND.n820 0.152939
R10439 GND.n5284 GND.n820 0.152939
R10440 GND.n5285 GND.n5284 0.152939
R10441 GND.n5286 GND.n5285 0.152939
R10442 GND.n5286 GND.n814 0.152939
R10443 GND.n5294 GND.n814 0.152939
R10444 GND.n5295 GND.n5294 0.152939
R10445 GND.n5296 GND.n5295 0.152939
R10446 GND.n5296 GND.n808 0.152939
R10447 GND.n5304 GND.n808 0.152939
R10448 GND.n5305 GND.n5304 0.152939
R10449 GND.n5306 GND.n5305 0.152939
R10450 GND.n5306 GND.n802 0.152939
R10451 GND.n5314 GND.n802 0.152939
R10452 GND.n5315 GND.n5314 0.152939
R10453 GND.n5316 GND.n5315 0.152939
R10454 GND.n5316 GND.n796 0.152939
R10455 GND.n5324 GND.n796 0.152939
R10456 GND.n5325 GND.n5324 0.152939
R10457 GND.n5326 GND.n5325 0.152939
R10458 GND.n5326 GND.n790 0.152939
R10459 GND.n5334 GND.n790 0.152939
R10460 GND.n5335 GND.n5334 0.152939
R10461 GND.n5336 GND.n5335 0.152939
R10462 GND.n5336 GND.n784 0.152939
R10463 GND.n5344 GND.n784 0.152939
R10464 GND.n5345 GND.n5344 0.152939
R10465 GND.n5346 GND.n5345 0.152939
R10466 GND.n5346 GND.n778 0.152939
R10467 GND.n5354 GND.n778 0.152939
R10468 GND.n5355 GND.n5354 0.152939
R10469 GND.n5356 GND.n5355 0.152939
R10470 GND.n5356 GND.n772 0.152939
R10471 GND.n5364 GND.n772 0.152939
R10472 GND.n5365 GND.n5364 0.152939
R10473 GND.n5366 GND.n5365 0.152939
R10474 GND.n5366 GND.n766 0.152939
R10475 GND.n5374 GND.n766 0.152939
R10476 GND.n5375 GND.n5374 0.152939
R10477 GND.n5376 GND.n5375 0.152939
R10478 GND.n5376 GND.n760 0.152939
R10479 GND.n5384 GND.n760 0.152939
R10480 GND.n5385 GND.n5384 0.152939
R10481 GND.n5386 GND.n5385 0.152939
R10482 GND.n5386 GND.n754 0.152939
R10483 GND.n5394 GND.n754 0.152939
R10484 GND.n5395 GND.n5394 0.152939
R10485 GND.n5396 GND.n5395 0.152939
R10486 GND.n5396 GND.n748 0.152939
R10487 GND.n5404 GND.n748 0.152939
R10488 GND.n5405 GND.n5404 0.152939
R10489 GND.n5406 GND.n5405 0.152939
R10490 GND.n5406 GND.n742 0.152939
R10491 GND.n5414 GND.n742 0.152939
R10492 GND.n5415 GND.n5414 0.152939
R10493 GND.n5416 GND.n5415 0.152939
R10494 GND.n5416 GND.n736 0.152939
R10495 GND.n5424 GND.n736 0.152939
R10496 GND.n5425 GND.n5424 0.152939
R10497 GND.n5426 GND.n5425 0.152939
R10498 GND.n5426 GND.n730 0.152939
R10499 GND.n5434 GND.n730 0.152939
R10500 GND.n5435 GND.n5434 0.152939
R10501 GND.n5436 GND.n5435 0.152939
R10502 GND.n5436 GND.n724 0.152939
R10503 GND.n5444 GND.n724 0.152939
R10504 GND.n5445 GND.n5444 0.152939
R10505 GND.n5446 GND.n5445 0.152939
R10506 GND.n5446 GND.n718 0.152939
R10507 GND.n5454 GND.n718 0.152939
R10508 GND.n5455 GND.n5454 0.152939
R10509 GND.n5456 GND.n5455 0.152939
R10510 GND.n5456 GND.n712 0.152939
R10511 GND.n5464 GND.n712 0.152939
R10512 GND.n5465 GND.n5464 0.152939
R10513 GND.n5466 GND.n5465 0.152939
R10514 GND.n5466 GND.n706 0.152939
R10515 GND.n5474 GND.n706 0.152939
R10516 GND.n5475 GND.n5474 0.152939
R10517 GND.n5476 GND.n5475 0.152939
R10518 GND.n5476 GND.n701 0.152939
R10519 GND.n5486 GND.n5485 0.152939
R10520 GND.n5487 GND.n5486 0.152939
R10521 GND.n5487 GND.n695 0.152939
R10522 GND.n5495 GND.n695 0.152939
R10523 GND.n5496 GND.n5495 0.152939
R10524 GND.n5497 GND.n5496 0.152939
R10525 GND.n5497 GND.n689 0.152939
R10526 GND.n5505 GND.n689 0.152939
R10527 GND.n5506 GND.n5505 0.152939
R10528 GND.n5507 GND.n5506 0.152939
R10529 GND.n5507 GND.n683 0.152939
R10530 GND.n5515 GND.n683 0.152939
R10531 GND.n5516 GND.n5515 0.152939
R10532 GND.n5517 GND.n5516 0.152939
R10533 GND.n5517 GND.n677 0.152939
R10534 GND.n5525 GND.n677 0.152939
R10535 GND.n5526 GND.n5525 0.152939
R10536 GND.n5527 GND.n5526 0.152939
R10537 GND.n5527 GND.n671 0.152939
R10538 GND.n5535 GND.n671 0.152939
R10539 GND.n5536 GND.n5535 0.152939
R10540 GND.n5537 GND.n5536 0.152939
R10541 GND.n5537 GND.n665 0.152939
R10542 GND.n5545 GND.n665 0.152939
R10543 GND.n5546 GND.n5545 0.152939
R10544 GND.n5547 GND.n5546 0.152939
R10545 GND.n5547 GND.n659 0.152939
R10546 GND.n5555 GND.n659 0.152939
R10547 GND.n5556 GND.n5555 0.152939
R10548 GND.n5557 GND.n5556 0.152939
R10549 GND.n5557 GND.n653 0.152939
R10550 GND.n5565 GND.n653 0.152939
R10551 GND.n5566 GND.n5565 0.152939
R10552 GND.n5567 GND.n5566 0.152939
R10553 GND.n5567 GND.n647 0.152939
R10554 GND.n5575 GND.n647 0.152939
R10555 GND.n5576 GND.n5575 0.152939
R10556 GND.n5577 GND.n5576 0.152939
R10557 GND.n5577 GND.n641 0.152939
R10558 GND.n5585 GND.n641 0.152939
R10559 GND.n5586 GND.n5585 0.152939
R10560 GND.n5587 GND.n5586 0.152939
R10561 GND.n5587 GND.n635 0.152939
R10562 GND.n5595 GND.n635 0.152939
R10563 GND.n5596 GND.n5595 0.152939
R10564 GND.n5597 GND.n5596 0.152939
R10565 GND.n5597 GND.n629 0.152939
R10566 GND.n5605 GND.n629 0.152939
R10567 GND.n5606 GND.n5605 0.152939
R10568 GND.n5607 GND.n5606 0.152939
R10569 GND.n5607 GND.n623 0.152939
R10570 GND.n5615 GND.n623 0.152939
R10571 GND.n5616 GND.n5615 0.152939
R10572 GND.n5617 GND.n5616 0.152939
R10573 GND.n5617 GND.n617 0.152939
R10574 GND.n5625 GND.n617 0.152939
R10575 GND.n5626 GND.n5625 0.152939
R10576 GND.n5627 GND.n5626 0.152939
R10577 GND.n5627 GND.n611 0.152939
R10578 GND.n5635 GND.n611 0.152939
R10579 GND.n5636 GND.n5635 0.152939
R10580 GND.n5637 GND.n5636 0.152939
R10581 GND.n5637 GND.n605 0.152939
R10582 GND.n5645 GND.n605 0.152939
R10583 GND.n5646 GND.n5645 0.152939
R10584 GND.n5648 GND.n5646 0.152939
R10585 GND.n5648 GND.n5647 0.152939
R10586 GND.n5647 GND.n599 0.152939
R10587 GND.n5658 GND.n599 0.152939
R10588 GND.n4273 GND.n4272 0.152939
R10589 GND.n4274 GND.n4273 0.152939
R10590 GND.n4275 GND.n4274 0.152939
R10591 GND.n4278 GND.n4275 0.152939
R10592 GND.n4279 GND.n4278 0.152939
R10593 GND.n4280 GND.n4279 0.152939
R10594 GND.n4281 GND.n4280 0.152939
R10595 GND.n4283 GND.n4281 0.152939
R10596 GND.n4285 GND.n4283 0.152939
R10597 GND.n4285 GND.n4284 0.152939
R10598 GND.n4284 GND.n593 0.152939
R10599 GND.n594 GND.n593 0.152939
R10600 GND.n595 GND.n594 0.152939
R10601 GND.n598 GND.n595 0.152939
R10602 GND.n5659 GND.n598 0.152939
R10603 GND.n355 GND.n328 0.152939
R10604 GND.n356 GND.n355 0.152939
R10605 GND.n357 GND.n356 0.152939
R10606 GND.n375 GND.n357 0.152939
R10607 GND.n376 GND.n375 0.152939
R10608 GND.n377 GND.n376 0.152939
R10609 GND.n378 GND.n377 0.152939
R10610 GND.n396 GND.n378 0.152939
R10611 GND.n397 GND.n396 0.152939
R10612 GND.n398 GND.n397 0.152939
R10613 GND.n399 GND.n398 0.152939
R10614 GND.n416 GND.n399 0.152939
R10615 GND.n417 GND.n416 0.152939
R10616 GND.n418 GND.n417 0.152939
R10617 GND.n419 GND.n418 0.152939
R10618 GND.n436 GND.n419 0.152939
R10619 GND.n437 GND.n436 0.152939
R10620 GND.n438 GND.n437 0.152939
R10621 GND.n439 GND.n438 0.152939
R10622 GND.n455 GND.n439 0.152939
R10623 GND.n456 GND.n455 0.152939
R10624 GND.n457 GND.n456 0.152939
R10625 GND.n458 GND.n457 0.152939
R10626 GND.n473 GND.n458 0.152939
R10627 GND.n5830 GND.n473 0.152939
R10628 GND.n3992 GND.n3987 0.152939
R10629 GND.n3987 GND.n2780 0.152939
R10630 GND.n4111 GND.n2780 0.152939
R10631 GND.n4112 GND.n4111 0.152939
R10632 GND.n4113 GND.n4112 0.152939
R10633 GND.n4113 GND.n2776 0.152939
R10634 GND.n4126 GND.n2776 0.152939
R10635 GND.n4127 GND.n4126 0.152939
R10636 GND.n4128 GND.n4127 0.152939
R10637 GND.n4128 GND.n2772 0.152939
R10638 GND.n4141 GND.n2772 0.152939
R10639 GND.n4142 GND.n4141 0.152939
R10640 GND.n4143 GND.n4142 0.152939
R10641 GND.n4143 GND.n2767 0.152939
R10642 GND.n4156 GND.n2767 0.152939
R10643 GND.n4157 GND.n4156 0.152939
R10644 GND.n4158 GND.n4157 0.152939
R10645 GND.n4158 GND.n2763 0.152939
R10646 GND.n4171 GND.n2763 0.152939
R10647 GND.n4172 GND.n4171 0.152939
R10648 GND.n4173 GND.n4172 0.152939
R10649 GND.n4173 GND.n2759 0.152939
R10650 GND.n4186 GND.n2759 0.152939
R10651 GND.n4187 GND.n4186 0.152939
R10652 GND.n4188 GND.n4187 0.152939
R10653 GND.n4189 GND.n4188 0.152939
R10654 GND.n4190 GND.n4189 0.152939
R10655 GND.n4191 GND.n4190 0.152939
R10656 GND.n4192 GND.n4191 0.152939
R10657 GND.n4192 GND.n314 0.152939
R10658 GND.n5921 GND.n315 0.152939
R10659 GND.n2748 GND.n315 0.152939
R10660 GND.n4225 GND.n2748 0.152939
R10661 GND.n4226 GND.n4225 0.152939
R10662 GND.n4228 GND.n4226 0.152939
R10663 GND.n4228 GND.n4227 0.152939
R10664 GND.n4227 GND.n2742 0.152939
R10665 GND.n2743 GND.n2742 0.152939
R10666 GND.n2744 GND.n2743 0.152939
R10667 GND.n4240 GND.n2744 0.152939
R10668 GND.n4241 GND.n4240 0.152939
R10669 GND.n4242 GND.n4241 0.152939
R10670 GND.n4243 GND.n4242 0.152939
R10671 GND.n4244 GND.n4243 0.152939
R10672 GND.n4246 GND.n4244 0.152939
R10673 GND.n4246 GND.n4245 0.152939
R10674 GND.n4245 GND.n585 0.152939
R10675 GND.n5703 GND.n585 0.152939
R10676 GND.n5704 GND.n5703 0.152939
R10677 GND.n5705 GND.n5704 0.152939
R10678 GND.n5705 GND.n583 0.152939
R10679 GND.n5710 GND.n583 0.152939
R10680 GND.n5711 GND.n5710 0.152939
R10681 GND.n5712 GND.n5711 0.152939
R10682 GND.n5712 GND.n580 0.152939
R10683 GND.n5717 GND.n580 0.152939
R10684 GND.n5718 GND.n5717 0.152939
R10685 GND.n5719 GND.n5718 0.152939
R10686 GND.n5719 GND.n577 0.152939
R10687 GND.n5724 GND.n577 0.152939
R10688 GND.n5757 GND.n543 0.152939
R10689 GND.n545 GND.n543 0.152939
R10690 GND.n549 GND.n545 0.152939
R10691 GND.n550 GND.n549 0.152939
R10692 GND.n551 GND.n550 0.152939
R10693 GND.n552 GND.n551 0.152939
R10694 GND.n556 GND.n552 0.152939
R10695 GND.n557 GND.n556 0.152939
R10696 GND.n558 GND.n557 0.152939
R10697 GND.n559 GND.n558 0.152939
R10698 GND.n563 GND.n559 0.152939
R10699 GND.n564 GND.n563 0.152939
R10700 GND.n565 GND.n564 0.152939
R10701 GND.n566 GND.n565 0.152939
R10702 GND.n570 GND.n566 0.152939
R10703 GND.n571 GND.n570 0.152939
R10704 GND.n5726 GND.n571 0.152939
R10705 GND.n5726 GND.n5725 0.152939
R10706 GND.n5829 GND.n474 0.152939
R10707 GND.n476 GND.n474 0.152939
R10708 GND.n480 GND.n476 0.152939
R10709 GND.n481 GND.n480 0.152939
R10710 GND.n482 GND.n481 0.152939
R10711 GND.n483 GND.n482 0.152939
R10712 GND.n487 GND.n483 0.152939
R10713 GND.n488 GND.n487 0.152939
R10714 GND.n489 GND.n488 0.152939
R10715 GND.n490 GND.n489 0.152939
R10716 GND.n494 GND.n490 0.152939
R10717 GND.n495 GND.n494 0.152939
R10718 GND.n496 GND.n495 0.152939
R10719 GND.n497 GND.n496 0.152939
R10720 GND.n501 GND.n497 0.152939
R10721 GND.n502 GND.n501 0.152939
R10722 GND.n503 GND.n502 0.152939
R10723 GND.n504 GND.n503 0.152939
R10724 GND.n508 GND.n504 0.152939
R10725 GND.n509 GND.n508 0.152939
R10726 GND.n510 GND.n509 0.152939
R10727 GND.n511 GND.n510 0.152939
R10728 GND.n515 GND.n511 0.152939
R10729 GND.n516 GND.n515 0.152939
R10730 GND.n517 GND.n516 0.152939
R10731 GND.n518 GND.n517 0.152939
R10732 GND.n522 GND.n518 0.152939
R10733 GND.n523 GND.n522 0.152939
R10734 GND.n524 GND.n523 0.152939
R10735 GND.n525 GND.n524 0.152939
R10736 GND.n529 GND.n525 0.152939
R10737 GND.n530 GND.n529 0.152939
R10738 GND.n531 GND.n530 0.152939
R10739 GND.n532 GND.n531 0.152939
R10740 GND.n536 GND.n532 0.152939
R10741 GND.n537 GND.n536 0.152939
R10742 GND.n5760 GND.n537 0.152939
R10743 GND.n5760 GND.n5759 0.152939
R10744 GND.n2521 GND.n2520 0.152939
R10745 GND.n2522 GND.n2521 0.152939
R10746 GND.n2523 GND.n2522 0.152939
R10747 GND.n2524 GND.n2523 0.152939
R10748 GND.n2525 GND.n2524 0.152939
R10749 GND.n2526 GND.n2525 0.152939
R10750 GND.n2527 GND.n2526 0.152939
R10751 GND.n2528 GND.n2527 0.152939
R10752 GND.n2529 GND.n2528 0.152939
R10753 GND.n2530 GND.n2529 0.152939
R10754 GND.n2531 GND.n2530 0.152939
R10755 GND.n2532 GND.n2531 0.152939
R10756 GND.n2533 GND.n2532 0.152939
R10757 GND.n2534 GND.n2533 0.152939
R10758 GND.n2535 GND.n2534 0.152939
R10759 GND.n2542 GND.n2541 0.152939
R10760 GND.n2543 GND.n2542 0.152939
R10761 GND.n2544 GND.n2543 0.152939
R10762 GND.n2545 GND.n2544 0.152939
R10763 GND.n2546 GND.n2545 0.152939
R10764 GND.n2547 GND.n2546 0.152939
R10765 GND.n2548 GND.n2547 0.152939
R10766 GND.n2549 GND.n2548 0.152939
R10767 GND.n2550 GND.n2549 0.152939
R10768 GND.n2551 GND.n2550 0.152939
R10769 GND.n2552 GND.n2551 0.152939
R10770 GND.n2553 GND.n2552 0.152939
R10771 GND.n2554 GND.n2553 0.152939
R10772 GND.n2555 GND.n2554 0.152939
R10773 GND.n2556 GND.n2555 0.152939
R10774 GND.n2557 GND.n2556 0.152939
R10775 GND.n2558 GND.n2557 0.152939
R10776 GND.n4413 GND.n2558 0.152939
R10777 GND.n4413 GND.n4412 0.152939
R10778 GND.n4412 GND.n4411 0.152939
R10779 GND.n2584 GND.n2583 0.152939
R10780 GND.n2585 GND.n2584 0.152939
R10781 GND.n2586 GND.n2585 0.152939
R10782 GND.n2587 GND.n2586 0.152939
R10783 GND.n2608 GND.n2587 0.152939
R10784 GND.n2609 GND.n2608 0.152939
R10785 GND.n2610 GND.n2609 0.152939
R10786 GND.n2611 GND.n2610 0.152939
R10787 GND.n2629 GND.n2611 0.152939
R10788 GND.n2630 GND.n2629 0.152939
R10789 GND.n2631 GND.n2630 0.152939
R10790 GND.n2632 GND.n2631 0.152939
R10791 GND.n2649 GND.n2632 0.152939
R10792 GND.n2650 GND.n2649 0.152939
R10793 GND.n2651 GND.n2650 0.152939
R10794 GND.n2652 GND.n2651 0.152939
R10795 GND.n2670 GND.n2652 0.152939
R10796 GND.n2671 GND.n2670 0.152939
R10797 GND.n2672 GND.n2671 0.152939
R10798 GND.n2673 GND.n2672 0.152939
R10799 GND.n2691 GND.n2673 0.152939
R10800 GND.n2692 GND.n2691 0.152939
R10801 GND.n2693 GND.n2692 0.152939
R10802 GND.n2694 GND.n2693 0.152939
R10803 GND.n2694 GND.n329 0.152939
R10804 GND.n2141 GND.n2140 0.152939
R10805 GND.n2142 GND.n2141 0.152939
R10806 GND.n2143 GND.n2142 0.152939
R10807 GND.n2146 GND.n2143 0.152939
R10808 GND.n2147 GND.n2146 0.152939
R10809 GND.n2148 GND.n2147 0.152939
R10810 GND.n2149 GND.n2148 0.152939
R10811 GND.n2154 GND.n2149 0.152939
R10812 GND.n2155 GND.n2154 0.152939
R10813 GND.n2156 GND.n2155 0.152939
R10814 GND.n2157 GND.n2156 0.152939
R10815 GND.n2160 GND.n2157 0.152939
R10816 GND.n2161 GND.n2160 0.152939
R10817 GND.n2162 GND.n2161 0.152939
R10818 GND.n2163 GND.n2162 0.152939
R10819 GND.n2164 GND.n2163 0.152939
R10820 GND.n2166 GND.n2164 0.152939
R10821 GND.n2166 GND.n2165 0.152939
R10822 GND.n2165 GND.n1424 0.152939
R10823 GND.n2292 GND.n1424 0.152939
R10824 GND.n2293 GND.n2292 0.152939
R10825 GND.n2294 GND.n2293 0.152939
R10826 GND.n2295 GND.n2294 0.152939
R10827 GND.n2296 GND.n2295 0.152939
R10828 GND.n2298 GND.n2296 0.152939
R10829 GND.n2298 GND.n2297 0.152939
R10830 GND.n2297 GND.n1310 0.152939
R10831 GND.n1311 GND.n1310 0.152939
R10832 GND.n1312 GND.n1311 0.152939
R10833 GND.n3396 GND.n1312 0.152939
R10834 GND.n3397 GND.n3396 0.152939
R10835 GND.n3414 GND.n3397 0.152939
R10836 GND.n3415 GND.n3414 0.152939
R10837 GND.n3416 GND.n3415 0.152939
R10838 GND.n3416 GND.n3384 0.152939
R10839 GND.n3434 GND.n3384 0.152939
R10840 GND.n3435 GND.n3434 0.152939
R10841 GND.n3436 GND.n3435 0.152939
R10842 GND.n3436 GND.n3371 0.152939
R10843 GND.n3454 GND.n3371 0.152939
R10844 GND.n3455 GND.n3454 0.152939
R10845 GND.n3456 GND.n3455 0.152939
R10846 GND.n3456 GND.n3175 0.152939
R10847 GND.n3475 GND.n3175 0.152939
R10848 GND.n3476 GND.n3475 0.152939
R10849 GND.n3477 GND.n3476 0.152939
R10850 GND.n3477 GND.n3138 0.152939
R10851 GND.n3509 GND.n3138 0.152939
R10852 GND.n3510 GND.n3509 0.152939
R10853 GND.n3511 GND.n3510 0.152939
R10854 GND.n3512 GND.n3511 0.152939
R10855 GND.n3512 GND.n3108 0.152939
R10856 GND.n3551 GND.n3108 0.152939
R10857 GND.n3552 GND.n3551 0.152939
R10858 GND.n3553 GND.n3552 0.152939
R10859 GND.n3554 GND.n3553 0.152939
R10860 GND.n3555 GND.n3554 0.152939
R10861 GND.n3558 GND.n3555 0.152939
R10862 GND.n3559 GND.n3558 0.152939
R10863 GND.n3560 GND.n3559 0.152939
R10864 GND.n3561 GND.n3560 0.152939
R10865 GND.n3561 GND.n3062 0.152939
R10866 GND.n3667 GND.n3062 0.152939
R10867 GND.n3668 GND.n3667 0.152939
R10868 GND.n3669 GND.n3668 0.152939
R10869 GND.n3670 GND.n3669 0.152939
R10870 GND.n3670 GND.n3033 0.152939
R10871 GND.n3711 GND.n3033 0.152939
R10872 GND.n3712 GND.n3711 0.152939
R10873 GND.n3713 GND.n3712 0.152939
R10874 GND.n3714 GND.n3713 0.152939
R10875 GND.n3715 GND.n3714 0.152939
R10876 GND.n3715 GND.n2997 0.152939
R10877 GND.n3771 GND.n2997 0.152939
R10878 GND.n3772 GND.n3771 0.152939
R10879 GND.n3773 GND.n3772 0.152939
R10880 GND.n3774 GND.n3773 0.152939
R10881 GND.n3774 GND.n2974 0.152939
R10882 GND.n3796 GND.n2974 0.152939
R10883 GND.n3797 GND.n3796 0.152939
R10884 GND.n3798 GND.n3797 0.152939
R10885 GND.n3798 GND.n2835 0.152939
R10886 GND.n3899 GND.n2835 0.152939
R10887 GND.n3900 GND.n3899 0.152939
R10888 GND.n3901 GND.n3900 0.152939
R10889 GND.n3901 GND.n2822 0.152939
R10890 GND.n3918 GND.n2822 0.152939
R10891 GND.n3919 GND.n3918 0.152939
R10892 GND.n3920 GND.n3919 0.152939
R10893 GND.n3920 GND.n2808 0.152939
R10894 GND.n3937 GND.n2808 0.152939
R10895 GND.n3938 GND.n3937 0.152939
R10896 GND.n3939 GND.n3938 0.152939
R10897 GND.n3940 GND.n3939 0.152939
R10898 GND.n3940 GND.n2794 0.152939
R10899 GND.n3959 GND.n2794 0.152939
R10900 GND.n3960 GND.n3959 0.152939
R10901 GND.n3961 GND.n3960 0.152939
R10902 GND.n3961 GND.n2789 0.152939
R10903 GND.n4026 GND.n2789 0.152939
R10904 GND.n4027 GND.n4026 0.152939
R10905 GND.n4028 GND.n4027 0.152939
R10906 GND.n4028 GND.n2785 0.152939
R10907 GND.n4034 GND.n2785 0.152939
R10908 GND.n4035 GND.n4034 0.152939
R10909 GND.n4036 GND.n4035 0.152939
R10910 GND.n4037 GND.n4036 0.152939
R10911 GND.n4038 GND.n4037 0.152939
R10912 GND.n4041 GND.n4038 0.152939
R10913 GND.n4042 GND.n4041 0.152939
R10914 GND.n4043 GND.n4042 0.152939
R10915 GND.n4044 GND.n4043 0.152939
R10916 GND.n4047 GND.n4044 0.152939
R10917 GND.n4048 GND.n4047 0.152939
R10918 GND.n4049 GND.n4048 0.152939
R10919 GND.n4050 GND.n4049 0.152939
R10920 GND.n4053 GND.n4050 0.152939
R10921 GND.n4054 GND.n4053 0.152939
R10922 GND.n4055 GND.n4054 0.152939
R10923 GND.n4056 GND.n4055 0.152939
R10924 GND.n4059 GND.n4056 0.152939
R10925 GND.n4060 GND.n4059 0.152939
R10926 GND.n4061 GND.n4060 0.152939
R10927 GND.n4062 GND.n4061 0.152939
R10928 GND.n4065 GND.n4062 0.152939
R10929 GND.n4066 GND.n4065 0.152939
R10930 GND.n4067 GND.n4066 0.152939
R10931 GND.n4068 GND.n4067 0.152939
R10932 GND.n2097 GND.n1496 0.152939
R10933 GND.n2205 GND.n1496 0.152939
R10934 GND.n2206 GND.n2205 0.152939
R10935 GND.n2207 GND.n2206 0.152939
R10936 GND.n2208 GND.n2207 0.152939
R10937 GND.n2208 GND.n1473 0.152939
R10938 GND.n2230 GND.n1473 0.152939
R10939 GND.n2231 GND.n2230 0.152939
R10940 GND.n2232 GND.n2231 0.152939
R10941 GND.n2233 GND.n2232 0.152939
R10942 GND.n2233 GND.n1452 0.152939
R10943 GND.n2254 GND.n1452 0.152939
R10944 GND.n2255 GND.n2254 0.152939
R10945 GND.n2256 GND.n2255 0.152939
R10946 GND.n2257 GND.n2256 0.152939
R10947 GND.n2257 GND.n1431 0.152939
R10948 GND.n2281 GND.n1431 0.152939
R10949 GND.n2282 GND.n2281 0.152939
R10950 GND.n2283 GND.n2282 0.152939
R10951 GND.n2283 GND.n1407 0.152939
R10952 GND.n2321 GND.n1407 0.152939
R10953 GND.n2322 GND.n2321 0.152939
R10954 GND.n2323 GND.n2322 0.152939
R10955 GND.n2323 GND.n1243 0.152939
R10956 GND.n4797 GND.n1243 0.152939
R10957 GND.n1913 GND.n1701 0.152939
R10958 GND.n1704 GND.n1701 0.152939
R10959 GND.n1705 GND.n1704 0.152939
R10960 GND.n1706 GND.n1705 0.152939
R10961 GND.n1709 GND.n1706 0.152939
R10962 GND.n1710 GND.n1709 0.152939
R10963 GND.n1711 GND.n1710 0.152939
R10964 GND.n1712 GND.n1711 0.152939
R10965 GND.n1715 GND.n1712 0.152939
R10966 GND.n1716 GND.n1715 0.152939
R10967 GND.n1717 GND.n1716 0.152939
R10968 GND.n1718 GND.n1717 0.152939
R10969 GND.n1721 GND.n1718 0.152939
R10970 GND.n1722 GND.n1721 0.152939
R10971 GND.n1723 GND.n1722 0.152939
R10972 GND.n1724 GND.n1723 0.152939
R10973 GND.n1730 GND.n1724 0.152939
R10974 GND.n1731 GND.n1730 0.152939
R10975 GND.n1732 GND.n1731 0.152939
R10976 GND.n1733 GND.n1732 0.152939
R10977 GND.n1736 GND.n1733 0.152939
R10978 GND.n1737 GND.n1736 0.152939
R10979 GND.n1738 GND.n1737 0.152939
R10980 GND.n1739 GND.n1738 0.152939
R10981 GND.n1742 GND.n1739 0.152939
R10982 GND.n1743 GND.n1742 0.152939
R10983 GND.n1744 GND.n1743 0.152939
R10984 GND.n1745 GND.n1744 0.152939
R10985 GND.n1748 GND.n1745 0.152939
R10986 GND.n1749 GND.n1748 0.152939
R10987 GND.n1750 GND.n1749 0.152939
R10988 GND.n1751 GND.n1750 0.152939
R10989 GND.n1754 GND.n1751 0.152939
R10990 GND.n1755 GND.n1754 0.152939
R10991 GND.n1756 GND.n1755 0.152939
R10992 GND.n1841 GND.n1756 0.152939
R10993 GND.n1841 GND.n1840 0.152939
R10994 GND.n1840 GND.n1839 0.152939
R10995 GND.n1915 GND.n1914 0.152939
R10996 GND.n1915 GND.n1675 0.152939
R10997 GND.n1951 GND.n1675 0.152939
R10998 GND.n1952 GND.n1951 0.152939
R10999 GND.n1953 GND.n1952 0.152939
R11000 GND.n1953 GND.n1656 0.152939
R11001 GND.n1980 GND.n1656 0.152939
R11002 GND.n1981 GND.n1980 0.152939
R11003 GND.n1983 GND.n1981 0.152939
R11004 GND.n1983 GND.n1982 0.152939
R11005 GND.n1982 GND.n1123 0.152939
R11006 GND.n1124 GND.n1123 0.152939
R11007 GND.n1125 GND.n1124 0.152939
R11008 GND.n1634 GND.n1125 0.152939
R11009 GND.n1635 GND.n1634 0.152939
R11010 GND.n1635 GND.n1612 0.152939
R11011 GND.n2024 GND.n1612 0.152939
R11012 GND.n2025 GND.n2024 0.152939
R11013 GND.n2026 GND.n2025 0.152939
R11014 GND.n2027 GND.n2026 0.152939
R11015 GND.n2027 GND.n1586 0.152939
R11016 GND.n2061 GND.n1586 0.152939
R11017 GND.n2062 GND.n2061 0.152939
R11018 GND.n2064 GND.n2062 0.152939
R11019 GND.n2064 GND.n2063 0.152939
R11020 GND.n4888 GND.n1112 0.152939
R11021 GND.n1628 GND.n1112 0.152939
R11022 GND.n1629 GND.n1628 0.152939
R11023 GND.n1630 GND.n1629 0.152939
R11024 GND.n1630 GND.n1622 0.152939
R11025 GND.n2010 GND.n1622 0.152939
R11026 GND.n2011 GND.n2010 0.152939
R11027 GND.n2012 GND.n2011 0.152939
R11028 GND.n2013 GND.n2012 0.152939
R11029 GND.n2013 GND.n1595 0.152939
R11030 GND.n2048 GND.n1595 0.152939
R11031 GND.n2049 GND.n2048 0.152939
R11032 GND.n2050 GND.n2049 0.152939
R11033 GND.n2050 GND.n1513 0.152939
R11034 GND.n2138 GND.n1513 0.152939
R11035 GND.n976 GND.n975 0.152939
R11036 GND.n977 GND.n976 0.152939
R11037 GND.n982 GND.n977 0.152939
R11038 GND.n983 GND.n982 0.152939
R11039 GND.n984 GND.n983 0.152939
R11040 GND.n985 GND.n984 0.152939
R11041 GND.n990 GND.n985 0.152939
R11042 GND.n991 GND.n990 0.152939
R11043 GND.n992 GND.n991 0.152939
R11044 GND.n993 GND.n992 0.152939
R11045 GND.n998 GND.n993 0.152939
R11046 GND.n999 GND.n998 0.152939
R11047 GND.n1000 GND.n999 0.152939
R11048 GND.n1001 GND.n1000 0.152939
R11049 GND.n1006 GND.n1001 0.152939
R11050 GND.n1007 GND.n1006 0.152939
R11051 GND.n1008 GND.n1007 0.152939
R11052 GND.n1009 GND.n1008 0.152939
R11053 GND.n1014 GND.n1009 0.152939
R11054 GND.n1015 GND.n1014 0.152939
R11055 GND.n1016 GND.n1015 0.152939
R11056 GND.n1017 GND.n1016 0.152939
R11057 GND.n1022 GND.n1017 0.152939
R11058 GND.n1023 GND.n1022 0.152939
R11059 GND.n1024 GND.n1023 0.152939
R11060 GND.n1025 GND.n1024 0.152939
R11061 GND.n1030 GND.n1025 0.152939
R11062 GND.n1031 GND.n1030 0.152939
R11063 GND.n1032 GND.n1031 0.152939
R11064 GND.n1033 GND.n1032 0.152939
R11065 GND.n1038 GND.n1033 0.152939
R11066 GND.n1039 GND.n1038 0.152939
R11067 GND.n1040 GND.n1039 0.152939
R11068 GND.n1041 GND.n1040 0.152939
R11069 GND.n1046 GND.n1041 0.152939
R11070 GND.n1047 GND.n1046 0.152939
R11071 GND.n1048 GND.n1047 0.152939
R11072 GND.n1049 GND.n1048 0.152939
R11073 GND.n1054 GND.n1049 0.152939
R11074 GND.n1055 GND.n1054 0.152939
R11075 GND.n1056 GND.n1055 0.152939
R11076 GND.n1057 GND.n1056 0.152939
R11077 GND.n1062 GND.n1057 0.152939
R11078 GND.n1063 GND.n1062 0.152939
R11079 GND.n1064 GND.n1063 0.152939
R11080 GND.n1065 GND.n1064 0.152939
R11081 GND.n1070 GND.n1065 0.152939
R11082 GND.n1071 GND.n1070 0.152939
R11083 GND.n1072 GND.n1071 0.152939
R11084 GND.n1073 GND.n1072 0.152939
R11085 GND.n1078 GND.n1073 0.152939
R11086 GND.n1079 GND.n1078 0.152939
R11087 GND.n1080 GND.n1079 0.152939
R11088 GND.n1081 GND.n1080 0.152939
R11089 GND.n1086 GND.n1081 0.152939
R11090 GND.n1087 GND.n1086 0.152939
R11091 GND.n1088 GND.n1087 0.152939
R11092 GND.n1089 GND.n1088 0.152939
R11093 GND.n1094 GND.n1089 0.152939
R11094 GND.n1095 GND.n1094 0.152939
R11095 GND.n1096 GND.n1095 0.152939
R11096 GND.n1097 GND.n1096 0.152939
R11097 GND.n1102 GND.n1097 0.152939
R11098 GND.n1103 GND.n1102 0.152939
R11099 GND.n1104 GND.n1103 0.152939
R11100 GND.n1105 GND.n1104 0.152939
R11101 GND.n1110 GND.n1105 0.152939
R11102 GND.n1111 GND.n1110 0.152939
R11103 GND.n4889 GND.n1111 0.152939
R11104 GND.n3407 GND.n3406 0.152939
R11105 GND.n3407 GND.n3391 0.152939
R11106 GND.n3425 GND.n3391 0.152939
R11107 GND.n3426 GND.n3425 0.152939
R11108 GND.n3427 GND.n3426 0.152939
R11109 GND.n3427 GND.n3378 0.152939
R11110 GND.n3445 GND.n3378 0.152939
R11111 GND.n3446 GND.n3445 0.152939
R11112 GND.n3447 GND.n3446 0.152939
R11113 GND.n3447 GND.n3365 0.152939
R11114 GND.n3466 GND.n3365 0.152939
R11115 GND.n3467 GND.n3466 0.152939
R11116 GND.n3468 GND.n3467 0.152939
R11117 GND.n3468 GND.n3169 0.152939
R11118 GND.n3485 GND.n3169 0.152939
R11119 GND.n3486 GND.n3485 0.152939
R11120 GND.n3487 GND.n3486 0.152939
R11121 GND.n3487 GND.n3123 0.152939
R11122 GND.n3528 GND.n3123 0.152939
R11123 GND.n3529 GND.n3528 0.152939
R11124 GND.n3537 GND.n3529 0.152939
R11125 GND.n3537 GND.n3536 0.152939
R11126 GND.n3536 GND.n3535 0.152939
R11127 GND.n3535 GND.n3530 0.152939
R11128 GND.n3530 GND.n3086 0.152939
R11129 GND.n3601 GND.n3086 0.152939
R11130 GND.n3602 GND.n3601 0.152939
R11131 GND.n3603 GND.n3602 0.152939
R11132 GND.n3603 GND.n3069 0.152939
R11133 GND.n3658 GND.n3069 0.152939
R11134 GND.n3659 GND.n3658 0.152939
R11135 GND.n3660 GND.n3659 0.152939
R11136 GND.n3660 GND.n3048 0.152939
R11137 GND.n3686 GND.n3048 0.152939
R11138 GND.n3687 GND.n3686 0.152939
R11139 GND.n3697 GND.n3687 0.152939
R11140 GND.n3697 GND.n3696 0.152939
R11141 GND.n3696 GND.n3695 0.152939
R11142 GND.n3695 GND.n3688 0.152939
R11143 GND.n3688 GND.n3006 0.152939
R11144 GND.n3752 GND.n3006 0.152939
R11145 GND.n3753 GND.n3752 0.152939
R11146 GND.n3764 GND.n3753 0.152939
R11147 GND.n3764 GND.n3763 0.152939
R11148 GND.n3763 GND.n3762 0.152939
R11149 GND.n3762 GND.n3754 0.152939
R11150 GND.n3758 GND.n3754 0.152939
R11151 GND.n3758 GND.n2898 0.152939
R11152 GND.n3821 GND.n2898 0.152939
R11153 GND.n3822 GND.n3821 0.152939
R11154 GND.n3823 GND.n3822 0.152939
R11155 GND.n3823 GND.n2829 0.152939
R11156 GND.n3908 GND.n2829 0.152939
R11157 GND.n3909 GND.n3908 0.152939
R11158 GND.n3910 GND.n3909 0.152939
R11159 GND.n3910 GND.n2815 0.152939
R11160 GND.n3927 GND.n2815 0.152939
R11161 GND.n3928 GND.n3927 0.152939
R11162 GND.n3929 GND.n3928 0.152939
R11163 GND.n3929 GND.n2800 0.152939
R11164 GND.n3948 GND.n2800 0.152939
R11165 GND.n3949 GND.n3948 0.152939
R11166 GND.n3950 GND.n3949 0.152939
R11167 GND.n3950 GND.n2433 0.152939
R11168 GND.n4536 GND.n2433 0.152939
R11169 GND.n4004 GND.n3985 0.152939
R11170 GND.n4014 GND.n3985 0.152939
R11171 GND.n4015 GND.n4014 0.152939
R11172 GND.n4017 GND.n4015 0.152939
R11173 GND.n4017 GND.n4016 0.152939
R11174 GND.n4639 GND.n2344 0.152939
R11175 GND.n4635 GND.n2344 0.152939
R11176 GND.n4635 GND.n4634 0.152939
R11177 GND.n4634 GND.n4633 0.152939
R11178 GND.n4633 GND.n2350 0.152939
R11179 GND.n4629 GND.n2350 0.152939
R11180 GND.n4629 GND.n4628 0.152939
R11181 GND.n4628 GND.n4627 0.152939
R11182 GND.n4627 GND.n2355 0.152939
R11183 GND.n4623 GND.n2355 0.152939
R11184 GND.n4623 GND.n4622 0.152939
R11185 GND.n4622 GND.n4621 0.152939
R11186 GND.n4621 GND.n2360 0.152939
R11187 GND.n4617 GND.n2360 0.152939
R11188 GND.n4617 GND.n4616 0.152939
R11189 GND.n4616 GND.n4615 0.152939
R11190 GND.n4615 GND.n2365 0.152939
R11191 GND.n4611 GND.n2365 0.152939
R11192 GND.n4611 GND.n4610 0.152939
R11193 GND.n4610 GND.n4609 0.152939
R11194 GND.n4609 GND.n2370 0.152939
R11195 GND.n4605 GND.n2370 0.152939
R11196 GND.n4605 GND.n4604 0.152939
R11197 GND.n4604 GND.n4603 0.152939
R11198 GND.n4603 GND.n2375 0.152939
R11199 GND.n4599 GND.n2375 0.152939
R11200 GND.n4599 GND.n4598 0.152939
R11201 GND.n4598 GND.n4597 0.152939
R11202 GND.n4597 GND.n2380 0.152939
R11203 GND.n4593 GND.n2380 0.152939
R11204 GND.n4593 GND.n4592 0.152939
R11205 GND.n4592 GND.n4591 0.152939
R11206 GND.n4591 GND.n2385 0.152939
R11207 GND.n4587 GND.n2385 0.152939
R11208 GND.n4587 GND.n4586 0.152939
R11209 GND.n4586 GND.n4585 0.152939
R11210 GND.n4585 GND.n2390 0.152939
R11211 GND.n4581 GND.n2390 0.152939
R11212 GND.n4581 GND.n4580 0.152939
R11213 GND.n4580 GND.n4579 0.152939
R11214 GND.n4579 GND.n2395 0.152939
R11215 GND.n4575 GND.n2395 0.152939
R11216 GND.n4575 GND.n4574 0.152939
R11217 GND.n4574 GND.n4573 0.152939
R11218 GND.n4573 GND.n2400 0.152939
R11219 GND.n4569 GND.n2400 0.152939
R11220 GND.n4569 GND.n4568 0.152939
R11221 GND.n4568 GND.n4567 0.152939
R11222 GND.n4567 GND.n2405 0.152939
R11223 GND.n4563 GND.n2405 0.152939
R11224 GND.n4563 GND.n4562 0.152939
R11225 GND.n4562 GND.n4561 0.152939
R11226 GND.n4561 GND.n2410 0.152939
R11227 GND.n4557 GND.n2410 0.152939
R11228 GND.n4557 GND.n4556 0.152939
R11229 GND.n4556 GND.n4555 0.152939
R11230 GND.n4555 GND.n2415 0.152939
R11231 GND.n4551 GND.n2415 0.152939
R11232 GND.n4551 GND.n4550 0.152939
R11233 GND.n4550 GND.n4549 0.152939
R11234 GND.n4549 GND.n2420 0.152939
R11235 GND.n4545 GND.n2420 0.152939
R11236 GND.n4545 GND.n4544 0.152939
R11237 GND.n4544 GND.n4543 0.152939
R11238 GND.n4543 GND.n2425 0.152939
R11239 GND.n4647 GND.n4646 0.152939
R11240 GND.n4646 GND.n4645 0.152939
R11241 GND.n4645 GND.n2335 0.152939
R11242 GND.n4641 GND.n2335 0.152939
R11243 GND.n4641 GND.n4640 0.152939
R11244 GND.n2082 GND.n2081 0.152939
R11245 GND.n2082 GND.n1564 0.152939
R11246 GND.n2086 GND.n1564 0.152939
R11247 GND.n2087 GND.n2086 0.152939
R11248 GND.n2091 GND.n2087 0.152939
R11249 GND.n2091 GND.n2090 0.152939
R11250 GND.n2090 GND.n2089 0.152939
R11251 GND.n2089 GND.n1485 0.152939
R11252 GND.n2215 GND.n1485 0.152939
R11253 GND.n2216 GND.n2215 0.152939
R11254 GND.n2218 GND.n2216 0.152939
R11255 GND.n2218 GND.n2217 0.152939
R11256 GND.n2217 GND.n1464 0.152939
R11257 GND.n2240 GND.n1464 0.152939
R11258 GND.n2241 GND.n2240 0.152939
R11259 GND.n2243 GND.n2241 0.152939
R11260 GND.n2243 GND.n2242 0.152939
R11261 GND.n2242 GND.n1442 0.152939
R11262 GND.n2264 GND.n1442 0.152939
R11263 GND.n2265 GND.n2264 0.152939
R11264 GND.n2270 GND.n2265 0.152939
R11265 GND.n2270 GND.n2269 0.152939
R11266 GND.n2269 GND.n2268 0.152939
R11267 GND.n2268 GND.n1419 0.152939
R11268 GND.n2312 GND.n1419 0.152939
R11269 GND.n2312 GND.n2311 0.152939
R11270 GND.n2311 GND.n2310 0.152939
R11271 GND.n2310 GND.n1420 0.152939
R11272 GND.n1420 GND.n1399 0.152939
R11273 GND.n2333 GND.n1399 0.152939
R11274 GND.n4796 GND.n1244 0.152939
R11275 GND.n4792 GND.n1244 0.152939
R11276 GND.n4792 GND.n4791 0.152939
R11277 GND.n4791 GND.n4790 0.152939
R11278 GND.n4790 GND.n1248 0.152939
R11279 GND.n4786 GND.n1248 0.152939
R11280 GND.n4786 GND.n4785 0.152939
R11281 GND.n4785 GND.n4784 0.152939
R11282 GND.n4784 GND.n1253 0.152939
R11283 GND.n4780 GND.n1253 0.152939
R11284 GND.n4780 GND.n4779 0.152939
R11285 GND.n4779 GND.n4778 0.152939
R11286 GND.n4778 GND.n1258 0.152939
R11287 GND.n4774 GND.n1258 0.152939
R11288 GND.n4774 GND.n4773 0.152939
R11289 GND.n4768 GND.n1263 0.152939
R11290 GND.n4768 GND.n4767 0.152939
R11291 GND.n4767 GND.n4766 0.152939
R11292 GND.n4766 GND.n1271 0.152939
R11293 GND.n4762 GND.n1271 0.152939
R11294 GND.n4762 GND.n4761 0.152939
R11295 GND.n4761 GND.n4760 0.152939
R11296 GND.n4760 GND.n1276 0.152939
R11297 GND.n4756 GND.n1276 0.152939
R11298 GND.n4756 GND.n4755 0.152939
R11299 GND.n4755 GND.n4754 0.152939
R11300 GND.n4754 GND.n1281 0.152939
R11301 GND.n4750 GND.n1281 0.152939
R11302 GND.n4750 GND.n4749 0.152939
R11303 GND.n4749 GND.n4748 0.152939
R11304 GND.n4748 GND.n1286 0.152939
R11305 GND.n4744 GND.n1286 0.152939
R11306 GND.n4744 GND.n4743 0.152939
R11307 GND.n4743 GND.n4742 0.152939
R11308 GND.n4742 GND.n1291 0.152939
R11309 GND.n1833 GND.n1768 0.152939
R11310 GND.n1826 GND.n1768 0.152939
R11311 GND.n1826 GND.n1825 0.152939
R11312 GND.n1825 GND.n1824 0.152939
R11313 GND.n1824 GND.n1772 0.152939
R11314 GND.n1820 GND.n1772 0.152939
R11315 GND.n1820 GND.n1819 0.152939
R11316 GND.n1819 GND.n1818 0.152939
R11317 GND.n1818 GND.n1779 0.152939
R11318 GND.n1814 GND.n1779 0.152939
R11319 GND.n1814 GND.n1813 0.152939
R11320 GND.n1813 GND.n1812 0.152939
R11321 GND.n1812 GND.n1787 0.152939
R11322 GND.n1808 GND.n1787 0.152939
R11323 GND.n1808 GND.n1807 0.152939
R11324 GND.n1807 GND.n1806 0.152939
R11325 GND.n1806 GND.n1795 0.152939
R11326 GND.n1795 GND.n1694 0.152939
R11327 GND.n1923 GND.n1922 0.152939
R11328 GND.n1937 GND.n1923 0.152939
R11329 GND.n1937 GND.n1936 0.152939
R11330 GND.n1936 GND.n1935 0.152939
R11331 GND.n1935 GND.n1924 0.152939
R11332 GND.n1931 GND.n1924 0.152939
R11333 GND.n1931 GND.n1930 0.152939
R11334 GND.n1930 GND.n1929 0.152939
R11335 GND.n1929 GND.n1648 0.152939
R11336 GND.n1990 GND.n1648 0.152939
R11337 GND.n1991 GND.n1990 0.152939
R11338 GND.n1992 GND.n1991 0.152939
R11339 GND.n1992 GND.n1643 0.152939
R11340 GND.n1999 GND.n1643 0.152939
R11341 GND.n2000 GND.n1999 0.152939
R11342 GND.n2002 GND.n2000 0.152939
R11343 GND.n2002 GND.n2001 0.152939
R11344 GND.n2001 GND.n1603 0.152939
R11345 GND.n2034 GND.n1603 0.152939
R11346 GND.n2035 GND.n2034 0.152939
R11347 GND.n2040 GND.n2035 0.152939
R11348 GND.n2040 GND.n2039 0.152939
R11349 GND.n2039 GND.n2038 0.152939
R11350 GND.n2038 GND.n2036 0.152939
R11351 GND.n2036 GND.n1577 0.152939
R11352 GND.n2072 GND.n1577 0.152939
R11353 GND.n2073 GND.n2072 0.152939
R11354 GND.n2074 GND.n2073 0.152939
R11355 GND.n2074 GND.n1573 0.152939
R11356 GND.n2079 GND.n1573 0.152939
R11357 GND.n4004 GND.n4003 0.145317
R11358 GND.n4647 GND.n2334 0.145317
R11359 GND.n2140 GND.n2139 0.107207
R11360 GND.n4068 GND.n330 0.107207
R11361 GND.n5914 GND.n328 0.0767195
R11362 GND.n5914 GND.n329 0.0767195
R11363 GND.n2097 GND.n1511 0.0767195
R11364 GND.n2063 GND.n1511 0.0767195
R11365 GND.n5922 GND.n314 0.0695946
R11366 GND.n5922 GND.n5921 0.0695946
R11367 GND.n2081 GND.n2080 0.0695946
R11368 GND.n2080 GND.n2079 0.0695946
R11369 GND.n4535 GND.n2434 0.063
R11370 GND.n3405 GND.n1233 0.063
R11371 GND.n2571 GND.n2434 0.048394
R11372 GND.n5758 GND.n467 0.048394
R11373 GND.n1834 GND.n1767 0.048394
R11374 GND.n4803 GND.n1233 0.048394
R11375 GND.n4272 GND.n330 0.0462317
R11376 GND.n2139 GND.n2138 0.0462317
R11377 GND.n4403 GND.n2571 0.0344674
R11378 GND.n4403 GND.n2573 0.0344674
R11379 GND.n2597 GND.n2573 0.0344674
R11380 GND.n2598 GND.n2597 0.0344674
R11381 GND.n2599 GND.n2598 0.0344674
R11382 GND.n2600 GND.n2599 0.0344674
R11383 GND.n4120 GND.n2600 0.0344674
R11384 GND.n4120 GND.n2619 0.0344674
R11385 GND.n2620 GND.n2619 0.0344674
R11386 GND.n2621 GND.n2620 0.0344674
R11387 GND.n4135 GND.n2621 0.0344674
R11388 GND.n4135 GND.n2640 0.0344674
R11389 GND.n2641 GND.n2640 0.0344674
R11390 GND.n2642 GND.n2641 0.0344674
R11391 GND.n4150 GND.n2642 0.0344674
R11392 GND.n4150 GND.n2660 0.0344674
R11393 GND.n2661 GND.n2660 0.0344674
R11394 GND.n2662 GND.n2661 0.0344674
R11395 GND.n4165 GND.n2662 0.0344674
R11396 GND.n4165 GND.n2681 0.0344674
R11397 GND.n2682 GND.n2681 0.0344674
R11398 GND.n2683 GND.n2682 0.0344674
R11399 GND.n4180 GND.n2683 0.0344674
R11400 GND.n4180 GND.n2702 0.0344674
R11401 GND.n2703 GND.n2702 0.0344674
R11402 GND.n2704 GND.n2703 0.0344674
R11403 GND.n4206 GND.n2704 0.0344674
R11404 GND.n4209 GND.n4206 0.0344674
R11405 GND.n4210 GND.n4209 0.0344674
R11406 GND.n4210 GND.n2728 0.0344674
R11407 GND.n2729 GND.n2728 0.0344674
R11408 GND.n2730 GND.n2729 0.0344674
R11409 GND.n4218 GND.n2730 0.0344674
R11410 GND.n4219 GND.n4218 0.0344674
R11411 GND.n4219 GND.n346 0.0344674
R11412 GND.n347 GND.n346 0.0344674
R11413 GND.n348 GND.n347 0.0344674
R11414 GND.n4235 GND.n348 0.0344674
R11415 GND.n4235 GND.n365 0.0344674
R11416 GND.n366 GND.n365 0.0344674
R11417 GND.n367 GND.n366 0.0344674
R11418 GND.n4238 GND.n367 0.0344674
R11419 GND.n4238 GND.n386 0.0344674
R11420 GND.n387 GND.n386 0.0344674
R11421 GND.n388 GND.n387 0.0344674
R11422 GND.n588 GND.n388 0.0344674
R11423 GND.n588 GND.n406 0.0344674
R11424 GND.n407 GND.n406 0.0344674
R11425 GND.n408 GND.n407 0.0344674
R11426 GND.n5673 GND.n408 0.0344674
R11427 GND.n5673 GND.n426 0.0344674
R11428 GND.n427 GND.n426 0.0344674
R11429 GND.n428 GND.n427 0.0344674
R11430 GND.n5674 GND.n428 0.0344674
R11431 GND.n5674 GND.n446 0.0344674
R11432 GND.n447 GND.n446 0.0344674
R11433 GND.n448 GND.n447 0.0344674
R11434 GND.n5675 GND.n448 0.0344674
R11435 GND.n5675 GND.n465 0.0344674
R11436 GND.n466 GND.n465 0.0344674
R11437 GND.n467 GND.n466 0.0344674
R11438 GND.n4002 GND.n4001 0.0344674
R11439 GND.n4651 GND.n1392 0.0344674
R11440 GND.n1767 GND.n1765 0.0344674
R11441 GND.n1765 GND.n1684 0.0344674
R11442 GND.n1945 GND.n1684 0.0344674
R11443 GND.n1945 GND.n1687 0.0344674
R11444 GND.n1687 GND.n1686 0.0344674
R11445 GND.n1686 GND.n1666 0.0344674
R11446 GND.n1974 GND.n1666 0.0344674
R11447 GND.n1974 GND.n1667 0.0344674
R11448 GND.n1970 GND.n1667 0.0344674
R11449 GND.n1970 GND.n1969 0.0344674
R11450 GND.n1969 GND.n1968 0.0344674
R11451 GND.n1968 GND.n1136 0.0344674
R11452 GND.n4875 GND.n1136 0.0344674
R11453 GND.n4875 GND.n1137 0.0344674
R11454 GND.n4871 GND.n1137 0.0344674
R11455 GND.n4871 GND.n4870 0.0344674
R11456 GND.n4870 GND.n4869 0.0344674
R11457 GND.n4869 GND.n1145 0.0344674
R11458 GND.n4865 GND.n1145 0.0344674
R11459 GND.n4865 GND.n4864 0.0344674
R11460 GND.n4864 GND.n4863 0.0344674
R11461 GND.n4863 GND.n1153 0.0344674
R11462 GND.n4859 GND.n1153 0.0344674
R11463 GND.n4859 GND.n4858 0.0344674
R11464 GND.n4858 GND.n4857 0.0344674
R11465 GND.n4857 GND.n1161 0.0344674
R11466 GND.n4853 GND.n1161 0.0344674
R11467 GND.n4853 GND.n4852 0.0344674
R11468 GND.n4852 GND.n4851 0.0344674
R11469 GND.n4851 GND.n1169 0.0344674
R11470 GND.n4847 GND.n1169 0.0344674
R11471 GND.n4847 GND.n4846 0.0344674
R11472 GND.n4846 GND.n4845 0.0344674
R11473 GND.n4845 GND.n1177 0.0344674
R11474 GND.n4841 GND.n1177 0.0344674
R11475 GND.n4841 GND.n4840 0.0344674
R11476 GND.n4840 GND.n4839 0.0344674
R11477 GND.n4839 GND.n1185 0.0344674
R11478 GND.n4835 GND.n1185 0.0344674
R11479 GND.n4835 GND.n4834 0.0344674
R11480 GND.n4834 GND.n4833 0.0344674
R11481 GND.n4833 GND.n1193 0.0344674
R11482 GND.n4829 GND.n1193 0.0344674
R11483 GND.n4829 GND.n4828 0.0344674
R11484 GND.n4828 GND.n4827 0.0344674
R11485 GND.n4827 GND.n1201 0.0344674
R11486 GND.n4823 GND.n1201 0.0344674
R11487 GND.n4823 GND.n4822 0.0344674
R11488 GND.n4822 GND.n4821 0.0344674
R11489 GND.n4821 GND.n1209 0.0344674
R11490 GND.n4817 GND.n1209 0.0344674
R11491 GND.n4817 GND.n4816 0.0344674
R11492 GND.n4816 GND.n4815 0.0344674
R11493 GND.n4815 GND.n1217 0.0344674
R11494 GND.n4811 GND.n1217 0.0344674
R11495 GND.n4811 GND.n4810 0.0344674
R11496 GND.n4810 GND.n4809 0.0344674
R11497 GND.n4809 GND.n1225 0.0344674
R11498 GND.n4805 GND.n1225 0.0344674
R11499 GND.n4805 GND.n4804 0.0344674
R11500 GND.n4804 GND.n4803 0.0344674
R11501 GND.n4535 GND.n4534 0.0334484
R11502 GND.n3405 GND.n1331 0.0334484
R11503 GND.n4534 GND.n2435 0.0188424
R11504 GND.n4531 GND.n4530 0.0188424
R11505 GND.n4527 GND.n2438 0.0188424
R11506 GND.n4526 GND.n2443 0.0188424
R11507 GND.n4523 GND.n4522 0.0188424
R11508 GND.n4519 GND.n2447 0.0188424
R11509 GND.n4518 GND.n2451 0.0188424
R11510 GND.n4515 GND.n4514 0.0188424
R11511 GND.n4511 GND.n2455 0.0188424
R11512 GND.n4510 GND.n2459 0.0188424
R11513 GND.n4507 GND.n4506 0.0188424
R11514 GND.n4503 GND.n2463 0.0188424
R11515 GND.n4502 GND.n2467 0.0188424
R11516 GND.n4499 GND.n4498 0.0188424
R11517 GND.n4495 GND.n2471 0.0188424
R11518 GND.n4494 GND.n2475 0.0188424
R11519 GND.n4491 GND.n4490 0.0188424
R11520 GND.n2482 GND.n2479 0.0188424
R11521 GND.n3996 GND.n3993 0.0188424
R11522 GND.n1333 GND.n1331 0.0188424
R11523 GND.n4698 GND.n4697 0.0188424
R11524 GND.n4694 GND.n1334 0.0188424
R11525 GND.n4693 GND.n1340 0.0188424
R11526 GND.n4690 GND.n4689 0.0188424
R11527 GND.n4686 GND.n1345 0.0188424
R11528 GND.n4685 GND.n1349 0.0188424
R11529 GND.n4682 GND.n4681 0.0188424
R11530 GND.n4678 GND.n1353 0.0188424
R11531 GND.n4677 GND.n1359 0.0188424
R11532 GND.n4674 GND.n4673 0.0188424
R11533 GND.n4670 GND.n1365 0.0188424
R11534 GND.n4669 GND.n1369 0.0188424
R11535 GND.n4666 GND.n4665 0.0188424
R11536 GND.n4662 GND.n1373 0.0188424
R11537 GND.n4661 GND.n1379 0.0188424
R11538 GND.n4658 GND.n4657 0.0188424
R11539 GND.n1389 GND.n1385 0.0188424
R11540 GND.n4652 GND.n1391 0.0188424
R11541 GND.n4531 GND.n2435 0.016125
R11542 GND.n4530 GND.n2438 0.016125
R11543 GND.n4527 GND.n4526 0.016125
R11544 GND.n4523 GND.n2443 0.016125
R11545 GND.n4522 GND.n2447 0.016125
R11546 GND.n4519 GND.n4518 0.016125
R11547 GND.n4515 GND.n2451 0.016125
R11548 GND.n4514 GND.n2455 0.016125
R11549 GND.n4511 GND.n4510 0.016125
R11550 GND.n4507 GND.n2459 0.016125
R11551 GND.n4506 GND.n2463 0.016125
R11552 GND.n4503 GND.n4502 0.016125
R11553 GND.n4499 GND.n2467 0.016125
R11554 GND.n4498 GND.n2471 0.016125
R11555 GND.n4495 GND.n4494 0.016125
R11556 GND.n4491 GND.n2475 0.016125
R11557 GND.n4490 GND.n2479 0.016125
R11558 GND.n3996 GND.n2482 0.016125
R11559 GND.n4001 GND.n3993 0.016125
R11560 GND.n4698 GND.n1333 0.016125
R11561 GND.n4697 GND.n1334 0.016125
R11562 GND.n4694 GND.n4693 0.016125
R11563 GND.n4690 GND.n1340 0.016125
R11564 GND.n4689 GND.n1345 0.016125
R11565 GND.n4686 GND.n4685 0.016125
R11566 GND.n4682 GND.n1349 0.016125
R11567 GND.n4681 GND.n1353 0.016125
R11568 GND.n4678 GND.n4677 0.016125
R11569 GND.n4674 GND.n1359 0.016125
R11570 GND.n4673 GND.n1365 0.016125
R11571 GND.n4670 GND.n4669 0.016125
R11572 GND.n4666 GND.n1369 0.016125
R11573 GND.n4665 GND.n1373 0.016125
R11574 GND.n4662 GND.n4661 0.016125
R11575 GND.n4658 GND.n1379 0.016125
R11576 GND.n4657 GND.n1385 0.016125
R11577 GND.n1391 GND.n1389 0.016125
R11578 GND.n4652 GND.n4651 0.016125
R11579 GND.n4003 GND.n4002 0.00219837
R11580 GND.n2334 GND.n1392 0.00219837
R11581 a_n8209_7799.n164 a_n8209_7799.t73 254.106
R11582 a_n8209_7799.n150 a_n8209_7799.t64 254.106
R11583 a_n8209_7799.n137 a_n8209_7799.t56 254.106
R11584 a_n8209_7799.n123 a_n8209_7799.t88 254.106
R11585 a_n8209_7799.n110 a_n8209_7799.t42 254.106
R11586 a_n8209_7799.n95 a_n8209_7799.t34 254.106
R11587 a_n8209_7799.n32 a_n8209_7799.t33 254.025
R11588 a_n8209_7799.n34 a_n8209_7799.t57 254.025
R11589 a_n8209_7799.n36 a_n8209_7799.t48 254.025
R11590 a_n8209_7799.n104 a_n8209_7799.t25 232.083
R11591 a_n8209_7799.n159 a_n8209_7799.t26 192.8
R11592 a_n8209_7799.n171 a_n8209_7799.t44 192.8
R11593 a_n8209_7799.n169 a_n8209_7799.t23 192.8
R11594 a_n8209_7799.n160 a_n8209_7799.t90 192.8
R11595 a_n8209_7799.n168 a_n8209_7799.t35 192.8
R11596 a_n8209_7799.n166 a_n8209_7799.t51 192.8
R11597 a_n8209_7799.n161 a_n8209_7799.t83 192.8
R11598 a_n8209_7799.n162 a_n8209_7799.t28 192.8
R11599 a_n8209_7799.n163 a_n8209_7799.t43 192.8
R11600 a_n8209_7799.n165 a_n8209_7799.t58 192.8
R11601 a_n8209_7799.n145 a_n8209_7799.t50 192.8
R11602 a_n8209_7799.n157 a_n8209_7799.t21 192.8
R11603 a_n8209_7799.n155 a_n8209_7799.t37 192.8
R11604 a_n8209_7799.n146 a_n8209_7799.t31 192.8
R11605 a_n8209_7799.n154 a_n8209_7799.t78 192.8
R11606 a_n8209_7799.n152 a_n8209_7799.t47 192.8
R11607 a_n8209_7799.n147 a_n8209_7799.t82 192.8
R11608 a_n8209_7799.n148 a_n8209_7799.t63 192.8
R11609 a_n8209_7799.n149 a_n8209_7799.t29 192.8
R11610 a_n8209_7799.n151 a_n8209_7799.t76 192.8
R11611 a_n8209_7799.n132 a_n8209_7799.t40 192.8
R11612 a_n8209_7799.n144 a_n8209_7799.t84 192.8
R11613 a_n8209_7799.n142 a_n8209_7799.t30 192.8
R11614 a_n8209_7799.n133 a_n8209_7799.t20 192.8
R11615 a_n8209_7799.n141 a_n8209_7799.t69 192.8
R11616 a_n8209_7799.n139 a_n8209_7799.t39 192.8
R11617 a_n8209_7799.n134 a_n8209_7799.t77 192.8
R11618 a_n8209_7799.n135 a_n8209_7799.t54 192.8
R11619 a_n8209_7799.n136 a_n8209_7799.t91 192.8
R11620 a_n8209_7799.n138 a_n8209_7799.t68 192.8
R11621 a_n8209_7799.n124 a_n8209_7799.t70 192.8
R11622 a_n8209_7799.n122 a_n8209_7799.t61 192.8
R11623 a_n8209_7799.n121 a_n8209_7799.t46 192.8
R11624 a_n8209_7799.n120 a_n8209_7799.t79 192.8
R11625 a_n8209_7799.n126 a_n8209_7799.t65 192.8
R11626 a_n8209_7799.n127 a_n8209_7799.t55 192.8
R11627 a_n8209_7799.n128 a_n8209_7799.t38 192.8
R11628 a_n8209_7799.n129 a_n8209_7799.t86 192.8
R11629 a_n8209_7799.n130 a_n8209_7799.t62 192.8
R11630 a_n8209_7799.n119 a_n8209_7799.t45 192.8
R11631 a_n8209_7799.n111 a_n8209_7799.t59 192.8
R11632 a_n8209_7799.n109 a_n8209_7799.t80 192.8
R11633 a_n8209_7799.n108 a_n8209_7799.t41 192.8
R11634 a_n8209_7799.n107 a_n8209_7799.t72 192.8
R11635 a_n8209_7799.n113 a_n8209_7799.t24 192.8
R11636 a_n8209_7799.n114 a_n8209_7799.t60 192.8
R11637 a_n8209_7799.n115 a_n8209_7799.t81 192.8
R11638 a_n8209_7799.n116 a_n8209_7799.t22 192.8
R11639 a_n8209_7799.n117 a_n8209_7799.t75 192.8
R11640 a_n8209_7799.n106 a_n8209_7799.t27 192.8
R11641 a_n8209_7799.n96 a_n8209_7799.t49 192.8
R11642 a_n8209_7799.n94 a_n8209_7799.t71 192.8
R11643 a_n8209_7799.n93 a_n8209_7799.t32 192.8
R11644 a_n8209_7799.n92 a_n8209_7799.t66 192.8
R11645 a_n8209_7799.n98 a_n8209_7799.t87 192.8
R11646 a_n8209_7799.n99 a_n8209_7799.t52 192.8
R11647 a_n8209_7799.n100 a_n8209_7799.t74 192.8
R11648 a_n8209_7799.n101 a_n8209_7799.t85 192.8
R11649 a_n8209_7799.n103 a_n8209_7799.t67 192.8
R11650 a_n8209_7799.n91 a_n8209_7799.t89 192.8
R11651 a_n8209_7799.n57 a_n8209_7799.n0 68.6201
R11652 a_n8209_7799.n1 a_n8209_7799.n0 39.6376
R11653 a_n8209_7799.n51 a_n8209_7799.n0 39.7274
R11654 a_n8209_7799.n56 a_n8209_7799.n0 68.6201
R11655 a_n8209_7799.n0 a_n8209_7799.n55 71.6402
R11656 a_n8209_7799.n167 a_n8209_7799.n12 161.3
R11657 a_n8209_7799.n12 a_n8209_7799.n52 68.6201
R11658 a_n8209_7799.n12 a_n8209_7799.n13 39.7274
R11659 a_n8209_7799.n12 a_n8209_7799.n54 71.4497
R11660 a_n8209_7799.n170 a_n8209_7799.n31 161.3
R11661 a_n8209_7799.n31 a_n8209_7799.n53 68.6201
R11662 a_n8209_7799.n61 a_n8209_7799.n2 68.6201
R11663 a_n8209_7799.n3 a_n8209_7799.n2 39.6376
R11664 a_n8209_7799.n48 a_n8209_7799.n2 39.7274
R11665 a_n8209_7799.n60 a_n8209_7799.n2 68.6201
R11666 a_n8209_7799.n2 a_n8209_7799.n59 71.6402
R11667 a_n8209_7799.n153 a_n8209_7799.n14 161.3
R11668 a_n8209_7799.n14 a_n8209_7799.n49 68.6201
R11669 a_n8209_7799.n14 a_n8209_7799.n15 39.7274
R11670 a_n8209_7799.n14 a_n8209_7799.n58 71.4497
R11671 a_n8209_7799.n156 a_n8209_7799.n33 161.3
R11672 a_n8209_7799.n33 a_n8209_7799.n50 68.6201
R11673 a_n8209_7799.n65 a_n8209_7799.n4 68.6201
R11674 a_n8209_7799.n5 a_n8209_7799.n4 39.6376
R11675 a_n8209_7799.n45 a_n8209_7799.n4 39.7274
R11676 a_n8209_7799.n64 a_n8209_7799.n4 68.6201
R11677 a_n8209_7799.n4 a_n8209_7799.n63 71.6402
R11678 a_n8209_7799.n140 a_n8209_7799.n16 161.3
R11679 a_n8209_7799.n16 a_n8209_7799.n46 68.6201
R11680 a_n8209_7799.n16 a_n8209_7799.n17 39.7274
R11681 a_n8209_7799.n16 a_n8209_7799.n62 71.4497
R11682 a_n8209_7799.n143 a_n8209_7799.n35 161.3
R11683 a_n8209_7799.n35 a_n8209_7799.n47 68.6201
R11684 a_n8209_7799.n10 a_n8209_7799.n68 68.6201
R11685 a_n8209_7799.n22 a_n8209_7799.n10 39.6376
R11686 a_n8209_7799.n42 a_n8209_7799.n10 39.7274
R11687 a_n8209_7799.n20 a_n8209_7799.n67 68.6201
R11688 a_n8209_7799.n21 a_n8209_7799.n20 39.6373
R11689 a_n8209_7799.n43 a_n8209_7799.n20 68.6201
R11690 a_n8209_7799.n20 a_n8209_7799.n125 161.3
R11691 a_n8209_7799.n66 a_n8209_7799.n18 68.7078
R11692 a_n8209_7799.n19 a_n8209_7799.n18 39.6376
R11693 a_n8209_7799.n44 a_n8209_7799.n18 68.6201
R11694 a_n8209_7799.n8 a_n8209_7799.n71 68.6201
R11695 a_n8209_7799.n27 a_n8209_7799.n8 39.6376
R11696 a_n8209_7799.n39 a_n8209_7799.n8 39.7274
R11697 a_n8209_7799.n25 a_n8209_7799.n70 68.6201
R11698 a_n8209_7799.n26 a_n8209_7799.n25 39.6373
R11699 a_n8209_7799.n40 a_n8209_7799.n25 68.6201
R11700 a_n8209_7799.n25 a_n8209_7799.n112 161.3
R11701 a_n8209_7799.n69 a_n8209_7799.n23 68.7078
R11702 a_n8209_7799.n24 a_n8209_7799.n23 39.6376
R11703 a_n8209_7799.n41 a_n8209_7799.n23 68.6201
R11704 a_n8209_7799.n79 a_n8209_7799.n78 74.6262
R11705 a_n8209_7799.n74 a_n8209_7799.n77 68.6201
R11706 a_n8209_7799.n76 a_n8209_7799.n75 71.8318
R11707 a_n8209_7799.n6 a_n8209_7799.n102 161.3
R11708 a_n8209_7799.n7 a_n8209_7799.n6 39.7274
R11709 a_n8209_7799.n6 a_n8209_7799.n73 68.6201
R11710 a_n8209_7799.n30 a_n8209_7799.n6 39.6373
R11711 a_n8209_7799.n37 a_n8209_7799.n6 68.6201
R11712 a_n8209_7799.n6 a_n8209_7799.n97 161.3
R11713 a_n8209_7799.n72 a_n8209_7799.n28 68.7078
R11714 a_n8209_7799.n29 a_n8209_7799.n28 39.6376
R11715 a_n8209_7799.n38 a_n8209_7799.n28 68.6201
R11716 a_n8209_7799.n87 a_n8209_7799.n85 109.74
R11717 a_n8209_7799.n82 a_n8209_7799.n80 109.74
R11718 a_n8209_7799.n89 a_n8209_7799.n88 109.166
R11719 a_n8209_7799.n87 a_n8209_7799.n86 109.166
R11720 a_n8209_7799.n82 a_n8209_7799.n81 109.166
R11721 a_n8209_7799.n84 a_n8209_7799.n83 109.166
R11722 a_n8209_7799.n181 a_n8209_7799.n180 84.3504
R11723 a_n8209_7799.n176 a_n8209_7799.n175 84.3502
R11724 a_n8209_7799.n180 a_n8209_7799.n179 84.35
R11725 a_n8209_7799.n178 a_n8209_7799.n177 84.0635
R11726 a_n8209_7799.n31 a_n8209_7799.n32 28.2026
R11727 a_n8209_7799.n33 a_n8209_7799.n34 28.2026
R11728 a_n8209_7799.n35 a_n8209_7799.n36 28.2026
R11729 a_n8209_7799.n10 a_n8209_7799.n11 28.2026
R11730 a_n8209_7799.n8 a_n8209_7799.n9 28.2026
R11731 a_n8209_7799.n105 a_n8209_7799.n104 80.6037
R11732 a_n8209_7799.n56 a_n8209_7799.n161 48.4088
R11733 a_n8209_7799.n57 a_n8209_7799.n165 47.9169
R11734 a_n8209_7799.n60 a_n8209_7799.n147 48.4088
R11735 a_n8209_7799.n61 a_n8209_7799.n151 47.9169
R11736 a_n8209_7799.n64 a_n8209_7799.n134 48.4088
R11737 a_n8209_7799.n65 a_n8209_7799.n138 47.9169
R11738 a_n8209_7799.n128 a_n8209_7799.n67 48.4088
R11739 a_n8209_7799.n119 a_n8209_7799.n68 47.9169
R11740 a_n8209_7799.n115 a_n8209_7799.n70 48.4088
R11741 a_n8209_7799.n106 a_n8209_7799.n71 47.9169
R11742 a_n8209_7799.n100 a_n8209_7799.n73 48.4088
R11743 a_n8209_7799.n91 a_n8209_7799.n77 47.9169
R11744 a_n8209_7799.n13 a_n8209_7799.n160 28.5572
R11745 a_n8209_7799.n15 a_n8209_7799.n146 28.5572
R11746 a_n8209_7799.n17 a_n8209_7799.n133 28.5572
R11747 a_n8209_7799.n125 a_n8209_7799.n66 48.9635
R11748 a_n8209_7799.n112 a_n8209_7799.n69 48.9635
R11749 a_n8209_7799.n97 a_n8209_7799.n72 48.9635
R11750 a_n8209_7799.n169 a_n8209_7799.n54 27.0108
R11751 a_n8209_7799.n155 a_n8209_7799.n58 27.0108
R11752 a_n8209_7799.n142 a_n8209_7799.n62 27.0108
R11753 a_n8209_7799.n121 a_n8209_7799.n19 41.2665
R11754 a_n8209_7799.n108 a_n8209_7799.n24 41.2665
R11755 a_n8209_7799.n93 a_n8209_7799.n29 41.2665
R11756 a_n8209_7799.n102 a_n8209_7799.n76 59.1846
R11757 a_n8209_7799.n167 a_n8209_7799.n55 58.5991
R11758 a_n8209_7799.n166 a_n8209_7799.n55 26.1378
R11759 a_n8209_7799.n153 a_n8209_7799.n59 58.5991
R11760 a_n8209_7799.n152 a_n8209_7799.n59 26.1378
R11761 a_n8209_7799.n140 a_n8209_7799.n63 58.5991
R11762 a_n8209_7799.n139 a_n8209_7799.n63 26.1378
R11763 a_n8209_7799.n127 a_n8209_7799.n21 40.5378
R11764 a_n8209_7799.n114 a_n8209_7799.n26 40.5378
R11765 a_n8209_7799.n99 a_n8209_7799.n30 40.5378
R11766 a_n8209_7799.n170 a_n8209_7799.n54 58.0115
R11767 a_n8209_7799.n1 a_n8209_7799.n163 39.8067
R11768 a_n8209_7799.n156 a_n8209_7799.n58 58.0115
R11769 a_n8209_7799.n3 a_n8209_7799.n149 39.8067
R11770 a_n8209_7799.n143 a_n8209_7799.n62 58.0115
R11771 a_n8209_7799.n5 a_n8209_7799.n136 39.8067
R11772 a_n8209_7799.n130 a_n8209_7799.n22 39.8067
R11773 a_n8209_7799.n117 a_n8209_7799.n27 39.8067
R11774 a_n8209_7799.n103 a_n8209_7799.n76 25.2628
R11775 a_n8209_7799.n165 a_n8209_7799.n164 33.0515
R11776 a_n8209_7799.n151 a_n8209_7799.n150 33.0515
R11777 a_n8209_7799.n138 a_n8209_7799.n137 33.0515
R11778 a_n8209_7799.n124 a_n8209_7799.n123 33.0515
R11779 a_n8209_7799.n111 a_n8209_7799.n110 33.0515
R11780 a_n8209_7799.n96 a_n8209_7799.n95 33.0515
R11781 a_n8209_7799.n180 a_n8209_7799.n178 30.5791
R11782 a_n8209_7799.n164 a_n8209_7799.n0 28.5514
R11783 a_n8209_7799.n150 a_n8209_7799.n2 28.5514
R11784 a_n8209_7799.n137 a_n8209_7799.n4 28.5514
R11785 a_n8209_7799.n123 a_n8209_7799.n18 28.5514
R11786 a_n8209_7799.n110 a_n8209_7799.n23 28.5514
R11787 a_n8209_7799.n95 a_n8209_7799.n28 28.5514
R11788 a_n8209_7799.n90 a_n8209_7799.n84 27.4144
R11789 a_n8209_7799.n32 a_n8209_7799.n159 33.1028
R11790 a_n8209_7799.n34 a_n8209_7799.n145 33.1028
R11791 a_n8209_7799.n36 a_n8209_7799.n132 33.1028
R11792 a_n8209_7799.t53 a_n8209_7799.n11 254.025
R11793 a_n8209_7799.t36 a_n8209_7799.n9 254.025
R11794 a_n8209_7799.n104 a_n8209_7799.n79 58.0598
R11795 a_n8209_7799.n161 a_n8209_7799.n51 28.5577
R11796 a_n8209_7799.n147 a_n8209_7799.n48 28.5577
R11797 a_n8209_7799.n134 a_n8209_7799.n45 28.5577
R11798 a_n8209_7799.n42 a_n8209_7799.n128 28.5577
R11799 a_n8209_7799.n39 a_n8209_7799.n115 28.5577
R11800 a_n8209_7799.n7 a_n8209_7799.n100 28.5577
R11801 a_n8209_7799.n52 a_n8209_7799.n160 48.4088
R11802 a_n8209_7799.n49 a_n8209_7799.n146 48.4088
R11803 a_n8209_7799.n46 a_n8209_7799.n133 48.4088
R11804 a_n8209_7799.n43 a_n8209_7799.n120 48.4088
R11805 a_n8209_7799.n40 a_n8209_7799.n107 48.4088
R11806 a_n8209_7799.n37 a_n8209_7799.n92 48.4088
R11807 a_n8209_7799.n53 a_n8209_7799.n159 47.9169
R11808 a_n8209_7799.n50 a_n8209_7799.n145 47.9169
R11809 a_n8209_7799.n47 a_n8209_7799.n132 47.9169
R11810 a_n8209_7799.n44 a_n8209_7799.n124 47.9169
R11811 a_n8209_7799.n41 a_n8209_7799.n111 47.9169
R11812 a_n8209_7799.n38 a_n8209_7799.n96 47.9169
R11813 a_n8209_7799.n90 a_n8209_7799.n89 17.7829
R11814 a_n8209_7799.n53 a_n8209_7799.n171 41.0312
R11815 a_n8209_7799.n57 a_n8209_7799.n163 41.0312
R11816 a_n8209_7799.n50 a_n8209_7799.n157 41.0312
R11817 a_n8209_7799.n61 a_n8209_7799.n149 41.0312
R11818 a_n8209_7799.n47 a_n8209_7799.n144 41.0312
R11819 a_n8209_7799.n65 a_n8209_7799.n136 41.0312
R11820 a_n8209_7799.n44 a_n8209_7799.n122 41.0312
R11821 a_n8209_7799.n68 a_n8209_7799.n130 41.0312
R11822 a_n8209_7799.n41 a_n8209_7799.n109 41.0312
R11823 a_n8209_7799.n71 a_n8209_7799.n117 41.0312
R11824 a_n8209_7799.n38 a_n8209_7799.n94 41.0312
R11825 a_n8209_7799.n77 a_n8209_7799.n103 41.0312
R11826 a_n8209_7799.n52 a_n8209_7799.n168 40.5394
R11827 a_n8209_7799.n166 a_n8209_7799.n56 40.5394
R11828 a_n8209_7799.n49 a_n8209_7799.n154 40.5394
R11829 a_n8209_7799.n152 a_n8209_7799.n60 40.5394
R11830 a_n8209_7799.n46 a_n8209_7799.n141 40.5394
R11831 a_n8209_7799.n139 a_n8209_7799.n64 40.5394
R11832 a_n8209_7799.n126 a_n8209_7799.n43 40.5394
R11833 a_n8209_7799.n67 a_n8209_7799.n127 40.5394
R11834 a_n8209_7799.n113 a_n8209_7799.n40 40.5394
R11835 a_n8209_7799.n70 a_n8209_7799.n114 40.5394
R11836 a_n8209_7799.n98 a_n8209_7799.n37 40.5394
R11837 a_n8209_7799.n73 a_n8209_7799.n99 40.5394
R11838 a_n8209_7799.n169 a_n8209_7799.n13 51.9316
R11839 a_n8209_7799.n51 a_n8209_7799.n162 51.931
R11840 a_n8209_7799.n155 a_n8209_7799.n15 51.9316
R11841 a_n8209_7799.n48 a_n8209_7799.n148 51.931
R11842 a_n8209_7799.n142 a_n8209_7799.n17 51.9316
R11843 a_n8209_7799.n45 a_n8209_7799.n135 51.931
R11844 a_n8209_7799.n66 a_n8209_7799.n121 39.872
R11845 a_n8209_7799.n129 a_n8209_7799.n42 51.931
R11846 a_n8209_7799.n69 a_n8209_7799.n108 39.872
R11847 a_n8209_7799.n116 a_n8209_7799.n39 51.931
R11848 a_n8209_7799.n72 a_n8209_7799.n93 39.872
R11849 a_n8209_7799.n101 a_n8209_7799.n7 51.931
R11850 a_n8209_7799.n176 a_n8209_7799.n174 12.3527
R11851 a_n8209_7799.n174 a_n8209_7799.n90 11.5231
R11852 a_n8209_7799.n158 a_n8209_7799.n35 9.07481
R11853 a_n8209_7799.n118 a_n8209_7799.n105 9.07481
R11854 a_n8209_7799.n1 a_n8209_7799.n162 41.266
R11855 a_n8209_7799.n3 a_n8209_7799.n148 41.266
R11856 a_n8209_7799.n5 a_n8209_7799.n135 41.266
R11857 a_n8209_7799.n22 a_n8209_7799.n129 41.266
R11858 a_n8209_7799.n27 a_n8209_7799.n116 41.266
R11859 a_n8209_7799.n102 a_n8209_7799.n101 8.60764
R11860 a_n8209_7799.n168 a_n8209_7799.n167 8.11581
R11861 a_n8209_7799.n154 a_n8209_7799.n153 8.11581
R11862 a_n8209_7799.n141 a_n8209_7799.n140 8.11581
R11863 a_n8209_7799.n21 a_n8209_7799.n126 40.5373
R11864 a_n8209_7799.n26 a_n8209_7799.n113 40.5373
R11865 a_n8209_7799.n30 a_n8209_7799.n98 40.5373
R11866 a_n8209_7799.n171 a_n8209_7799.n170 7.62397
R11867 a_n8209_7799.n157 a_n8209_7799.n156 7.62397
R11868 a_n8209_7799.n144 a_n8209_7799.n143 7.62397
R11869 a_n8209_7799.n19 a_n8209_7799.n122 39.8062
R11870 a_n8209_7799.n24 a_n8209_7799.n109 39.8062
R11871 a_n8209_7799.n29 a_n8209_7799.n94 39.8062
R11872 a_n8209_7799.n173 a_n8209_7799.n131 5.42817
R11873 a_n8209_7799.n88 a_n8209_7799.t7 5.418
R11874 a_n8209_7799.n88 a_n8209_7799.t19 5.418
R11875 a_n8209_7799.n86 a_n8209_7799.t6 5.418
R11876 a_n8209_7799.n86 a_n8209_7799.t11 5.418
R11877 a_n8209_7799.n85 a_n8209_7799.t5 5.418
R11878 a_n8209_7799.n85 a_n8209_7799.t0 5.418
R11879 a_n8209_7799.n80 a_n8209_7799.t13 5.418
R11880 a_n8209_7799.n80 a_n8209_7799.t10 5.418
R11881 a_n8209_7799.n81 a_n8209_7799.t18 5.418
R11882 a_n8209_7799.n81 a_n8209_7799.t2 5.418
R11883 a_n8209_7799.n83 a_n8209_7799.t12 5.418
R11884 a_n8209_7799.n83 a_n8209_7799.t17 5.418
R11885 a_n8209_7799.n173 a_n8209_7799.n172 5.22732
R11886 a_n8209_7799.n172 a_n8209_7799.n31 5.00473
R11887 a_n8209_7799.n158 a_n8209_7799.n33 5.00473
R11888 a_n8209_7799.n131 a_n8209_7799.n10 5.00473
R11889 a_n8209_7799.n118 a_n8209_7799.n8 5.00473
R11890 a_n8209_7799.n172 a_n8209_7799.n158 4.07058
R11891 a_n8209_7799.n131 a_n8209_7799.n118 4.07058
R11892 a_n8209_7799.n174 a_n8209_7799.n173 3.4105
R11893 a_n8209_7799.n179 a_n8209_7799.t8 3.3005
R11894 a_n8209_7799.n179 a_n8209_7799.t4 3.3005
R11895 a_n8209_7799.n177 a_n8209_7799.t14 3.3005
R11896 a_n8209_7799.n177 a_n8209_7799.t9 3.3005
R11897 a_n8209_7799.n175 a_n8209_7799.t15 3.3005
R11898 a_n8209_7799.n175 a_n8209_7799.t3 3.3005
R11899 a_n8209_7799.n181 a_n8209_7799.t16 3.3005
R11900 a_n8209_7799.t1 a_n8209_7799.n181 3.3005
R11901 a_n8209_7799.n11 a_n8209_7799.n119 33.1028
R11902 a_n8209_7799.n9 a_n8209_7799.n106 33.1028
R11903 a_n8209_7799.n79 a_n8209_7799.n91 12.7884
R11904 a_n8209_7799.n16 a_n8209_7799.n4 2.65202
R11905 a_n8209_7799.n14 a_n8209_7799.n2 2.65202
R11906 a_n8209_7799.n12 a_n8209_7799.n0 2.65202
R11907 a_n8209_7799.n89 a_n8209_7799.n87 0.573776
R11908 a_n8209_7799.n84 a_n8209_7799.n82 0.573776
R11909 a_n8209_7799.n78 a_n8209_7799.n74 0.379288
R11910 a_n8209_7799.n75 a_n8209_7799.n74 0.379288
R11911 a_n8209_7799.n178 a_n8209_7799.n176 0.287138
R11912 a_n8209_7799.n105 a_n8209_7799.n78 0.285035
R11913 a_n8209_7799.n125 a_n8209_7799.n120 0.246418
R11914 a_n8209_7799.n112 a_n8209_7799.n107 0.246418
R11915 a_n8209_7799.n97 a_n8209_7799.n92 0.246418
R11916 a_n8209_7799.n10 a_n8209_7799.n20 2.55776
R11917 a_n8209_7799.n8 a_n8209_7799.n25 2.55776
R11918 a_n8209_7799.n6 a_n8209_7799.n28 2.27323
R11919 a_n8209_7799.n25 a_n8209_7799.n23 2.27323
R11920 a_n8209_7799.n20 a_n8209_7799.n18 2.27323
R11921 a_n8209_7799.n35 a_n8209_7799.n16 2.17897
R11922 a_n8209_7799.n33 a_n8209_7799.n14 2.17897
R11923 a_n8209_7799.n31 a_n8209_7799.n12 2.17897
R11924 a_n8209_7799.n75 a_n8209_7799.n6 1.51565
R11925 VOUT.n212 VOUT.n210 103.684
R11926 VOUT.n200 VOUT.n198 103.684
R11927 VOUT.n189 VOUT.n187 103.684
R11928 VOUT.n25 VOUT.n23 103.684
R11929 VOUT.n13 VOUT.n11 103.684
R11930 VOUT.n2 VOUT.n0 103.684
R11931 VOUT.n218 VOUT.n217 103.111
R11932 VOUT.n216 VOUT.n215 103.111
R11933 VOUT.n214 VOUT.n213 103.111
R11934 VOUT.n212 VOUT.n211 103.111
R11935 VOUT.n208 VOUT.n207 103.111
R11936 VOUT.n206 VOUT.n205 103.111
R11937 VOUT.n204 VOUT.n203 103.111
R11938 VOUT.n202 VOUT.n201 103.111
R11939 VOUT.n200 VOUT.n199 103.111
R11940 VOUT.n197 VOUT.n196 103.111
R11941 VOUT.n195 VOUT.n194 103.111
R11942 VOUT.n193 VOUT.n192 103.111
R11943 VOUT.n191 VOUT.n190 103.111
R11944 VOUT.n189 VOUT.n188 103.111
R11945 VOUT.n25 VOUT.n24 103.111
R11946 VOUT.n27 VOUT.n26 103.111
R11947 VOUT.n29 VOUT.n28 103.111
R11948 VOUT.n31 VOUT.n30 103.111
R11949 VOUT.n33 VOUT.n32 103.111
R11950 VOUT.n13 VOUT.n12 103.111
R11951 VOUT.n15 VOUT.n14 103.111
R11952 VOUT.n17 VOUT.n16 103.111
R11953 VOUT.n19 VOUT.n18 103.111
R11954 VOUT.n21 VOUT.n20 103.111
R11955 VOUT.n2 VOUT.n1 103.111
R11956 VOUT.n4 VOUT.n3 103.111
R11957 VOUT.n6 VOUT.n5 103.111
R11958 VOUT.n8 VOUT.n7 103.111
R11959 VOUT.n10 VOUT.n9 103.111
R11960 VOUT.n220 VOUT.n219 103.111
R11961 VOUT.n234 VOUT.n232 81.9368
R11962 VOUT.n225 VOUT.n223 81.9368
R11963 VOUT.n254 VOUT.n252 81.9368
R11964 VOUT.n245 VOUT.n243 81.9368
R11965 VOUT.n240 VOUT.n239 80.9324
R11966 VOUT.n238 VOUT.n237 80.9324
R11967 VOUT.n236 VOUT.n235 80.9324
R11968 VOUT.n234 VOUT.n233 80.9324
R11969 VOUT.n231 VOUT.n230 80.9324
R11970 VOUT.n229 VOUT.n228 80.9324
R11971 VOUT.n227 VOUT.n226 80.9324
R11972 VOUT.n225 VOUT.n224 80.9324
R11973 VOUT.n254 VOUT.n253 80.9324
R11974 VOUT.n256 VOUT.n255 80.9324
R11975 VOUT.n258 VOUT.n257 80.9324
R11976 VOUT.n260 VOUT.n259 80.9324
R11977 VOUT.n245 VOUT.n244 80.9324
R11978 VOUT.n247 VOUT.n246 80.9324
R11979 VOUT.n249 VOUT.n248 80.9324
R11980 VOUT.n251 VOUT.n250 80.9324
R11981 VOUT.n242 VOUT.n222 8.55261
R11982 VOUT.n209 VOUT.n197 7.58994
R11983 VOUT.n22 VOUT.n10 7.58994
R11984 VOUT.n241 VOUT.n231 7.58886
R11985 VOUT.n261 VOUT.n251 7.58886
R11986 VOUT.n242 VOUT.n241 5.77257
R11987 VOUT.n262 VOUT.n261 5.77257
R11988 VOUT.n241 VOUT.n240 5.46817
R11989 VOUT.n261 VOUT.n260 5.46817
R11990 VOUT.n221 VOUT.n220 5.25266
R11991 VOUT.n209 VOUT.n208 5.25266
R11992 VOUT.n34 VOUT.n33 5.25266
R11993 VOUT.n22 VOUT.n21 5.25266
R11994 VOUT.n263 VOUT.n35 4.93275
R11995 VOUT.n222 VOUT.n221 4.78873
R11996 VOUT.n35 VOUT.n34 4.78873
R11997 VOUT.n126 VOUT.n79 4.5005
R11998 VOUT.n95 VOUT.n79 4.5005
R11999 VOUT.n90 VOUT.n74 4.5005
R12000 VOUT.n90 VOUT.n76 4.5005
R12001 VOUT.n90 VOUT.n73 4.5005
R12002 VOUT.n90 VOUT.n77 4.5005
R12003 VOUT.n90 VOUT.n72 4.5005
R12004 VOUT.n90 VOUT.t117 4.5005
R12005 VOUT.n90 VOUT.n71 4.5005
R12006 VOUT.n90 VOUT.n78 4.5005
R12007 VOUT.n90 VOUT.n79 4.5005
R12008 VOUT.n88 VOUT.n74 4.5005
R12009 VOUT.n88 VOUT.n76 4.5005
R12010 VOUT.n88 VOUT.n73 4.5005
R12011 VOUT.n88 VOUT.n77 4.5005
R12012 VOUT.n88 VOUT.n72 4.5005
R12013 VOUT.n88 VOUT.t117 4.5005
R12014 VOUT.n88 VOUT.n71 4.5005
R12015 VOUT.n88 VOUT.n78 4.5005
R12016 VOUT.n88 VOUT.n79 4.5005
R12017 VOUT.n87 VOUT.n74 4.5005
R12018 VOUT.n87 VOUT.n76 4.5005
R12019 VOUT.n87 VOUT.n73 4.5005
R12020 VOUT.n87 VOUT.n77 4.5005
R12021 VOUT.n87 VOUT.n72 4.5005
R12022 VOUT.n87 VOUT.t117 4.5005
R12023 VOUT.n87 VOUT.n71 4.5005
R12024 VOUT.n87 VOUT.n78 4.5005
R12025 VOUT.n87 VOUT.n79 4.5005
R12026 VOUT.n172 VOUT.n74 4.5005
R12027 VOUT.n172 VOUT.n76 4.5005
R12028 VOUT.n172 VOUT.n73 4.5005
R12029 VOUT.n172 VOUT.n77 4.5005
R12030 VOUT.n172 VOUT.n72 4.5005
R12031 VOUT.n172 VOUT.t117 4.5005
R12032 VOUT.n172 VOUT.n71 4.5005
R12033 VOUT.n172 VOUT.n78 4.5005
R12034 VOUT.n172 VOUT.n79 4.5005
R12035 VOUT.n170 VOUT.n74 4.5005
R12036 VOUT.n170 VOUT.n76 4.5005
R12037 VOUT.n170 VOUT.n73 4.5005
R12038 VOUT.n170 VOUT.n77 4.5005
R12039 VOUT.n170 VOUT.n72 4.5005
R12040 VOUT.n170 VOUT.t117 4.5005
R12041 VOUT.n170 VOUT.n71 4.5005
R12042 VOUT.n170 VOUT.n78 4.5005
R12043 VOUT.n168 VOUT.n74 4.5005
R12044 VOUT.n168 VOUT.n76 4.5005
R12045 VOUT.n168 VOUT.n73 4.5005
R12046 VOUT.n168 VOUT.n77 4.5005
R12047 VOUT.n168 VOUT.n72 4.5005
R12048 VOUT.n168 VOUT.t117 4.5005
R12049 VOUT.n168 VOUT.n71 4.5005
R12050 VOUT.n168 VOUT.n78 4.5005
R12051 VOUT.n98 VOUT.n74 4.5005
R12052 VOUT.n98 VOUT.n76 4.5005
R12053 VOUT.n98 VOUT.n73 4.5005
R12054 VOUT.n98 VOUT.n77 4.5005
R12055 VOUT.n98 VOUT.n72 4.5005
R12056 VOUT.n98 VOUT.t117 4.5005
R12057 VOUT.n98 VOUT.n71 4.5005
R12058 VOUT.n98 VOUT.n78 4.5005
R12059 VOUT.n98 VOUT.n79 4.5005
R12060 VOUT.n97 VOUT.n74 4.5005
R12061 VOUT.n97 VOUT.n76 4.5005
R12062 VOUT.n97 VOUT.n73 4.5005
R12063 VOUT.n97 VOUT.n77 4.5005
R12064 VOUT.n97 VOUT.n72 4.5005
R12065 VOUT.n97 VOUT.t117 4.5005
R12066 VOUT.n97 VOUT.n71 4.5005
R12067 VOUT.n97 VOUT.n78 4.5005
R12068 VOUT.n97 VOUT.n79 4.5005
R12069 VOUT.n101 VOUT.n74 4.5005
R12070 VOUT.n101 VOUT.n76 4.5005
R12071 VOUT.n101 VOUT.n73 4.5005
R12072 VOUT.n101 VOUT.n77 4.5005
R12073 VOUT.n101 VOUT.n72 4.5005
R12074 VOUT.n101 VOUT.t117 4.5005
R12075 VOUT.n101 VOUT.n71 4.5005
R12076 VOUT.n101 VOUT.n78 4.5005
R12077 VOUT.n101 VOUT.n79 4.5005
R12078 VOUT.n100 VOUT.n74 4.5005
R12079 VOUT.n100 VOUT.n76 4.5005
R12080 VOUT.n100 VOUT.n73 4.5005
R12081 VOUT.n100 VOUT.n77 4.5005
R12082 VOUT.n100 VOUT.n72 4.5005
R12083 VOUT.n100 VOUT.t117 4.5005
R12084 VOUT.n100 VOUT.n71 4.5005
R12085 VOUT.n100 VOUT.n78 4.5005
R12086 VOUT.n100 VOUT.n79 4.5005
R12087 VOUT.n83 VOUT.n74 4.5005
R12088 VOUT.n83 VOUT.n76 4.5005
R12089 VOUT.n83 VOUT.n73 4.5005
R12090 VOUT.n83 VOUT.n77 4.5005
R12091 VOUT.n83 VOUT.n72 4.5005
R12092 VOUT.n83 VOUT.t117 4.5005
R12093 VOUT.n83 VOUT.n71 4.5005
R12094 VOUT.n83 VOUT.n78 4.5005
R12095 VOUT.n83 VOUT.n79 4.5005
R12096 VOUT.n175 VOUT.n74 4.5005
R12097 VOUT.n175 VOUT.n76 4.5005
R12098 VOUT.n175 VOUT.n73 4.5005
R12099 VOUT.n175 VOUT.n77 4.5005
R12100 VOUT.n175 VOUT.n72 4.5005
R12101 VOUT.n175 VOUT.t117 4.5005
R12102 VOUT.n175 VOUT.n71 4.5005
R12103 VOUT.n175 VOUT.n78 4.5005
R12104 VOUT.n175 VOUT.n79 4.5005
R12105 VOUT.n162 VOUT.n133 4.5005
R12106 VOUT.n162 VOUT.n139 4.5005
R12107 VOUT.n120 VOUT.n109 4.5005
R12108 VOUT.n120 VOUT.n111 4.5005
R12109 VOUT.n120 VOUT.n108 4.5005
R12110 VOUT.n120 VOUT.n112 4.5005
R12111 VOUT.n120 VOUT.n107 4.5005
R12112 VOUT.n120 VOUT.t116 4.5005
R12113 VOUT.n120 VOUT.n106 4.5005
R12114 VOUT.n120 VOUT.n113 4.5005
R12115 VOUT.n162 VOUT.n120 4.5005
R12116 VOUT.n141 VOUT.n109 4.5005
R12117 VOUT.n141 VOUT.n111 4.5005
R12118 VOUT.n141 VOUT.n108 4.5005
R12119 VOUT.n141 VOUT.n112 4.5005
R12120 VOUT.n141 VOUT.n107 4.5005
R12121 VOUT.n141 VOUT.t116 4.5005
R12122 VOUT.n141 VOUT.n106 4.5005
R12123 VOUT.n141 VOUT.n113 4.5005
R12124 VOUT.n162 VOUT.n141 4.5005
R12125 VOUT.n119 VOUT.n109 4.5005
R12126 VOUT.n119 VOUT.n111 4.5005
R12127 VOUT.n119 VOUT.n108 4.5005
R12128 VOUT.n119 VOUT.n112 4.5005
R12129 VOUT.n119 VOUT.n107 4.5005
R12130 VOUT.n119 VOUT.t116 4.5005
R12131 VOUT.n119 VOUT.n106 4.5005
R12132 VOUT.n119 VOUT.n113 4.5005
R12133 VOUT.n162 VOUT.n119 4.5005
R12134 VOUT.n143 VOUT.n109 4.5005
R12135 VOUT.n143 VOUT.n111 4.5005
R12136 VOUT.n143 VOUT.n108 4.5005
R12137 VOUT.n143 VOUT.n112 4.5005
R12138 VOUT.n143 VOUT.n107 4.5005
R12139 VOUT.n143 VOUT.t116 4.5005
R12140 VOUT.n143 VOUT.n106 4.5005
R12141 VOUT.n143 VOUT.n113 4.5005
R12142 VOUT.n162 VOUT.n143 4.5005
R12143 VOUT.n109 VOUT.n104 4.5005
R12144 VOUT.n111 VOUT.n104 4.5005
R12145 VOUT.n108 VOUT.n104 4.5005
R12146 VOUT.n112 VOUT.n104 4.5005
R12147 VOUT.n107 VOUT.n104 4.5005
R12148 VOUT.t116 VOUT.n104 4.5005
R12149 VOUT.n106 VOUT.n104 4.5005
R12150 VOUT.n113 VOUT.n104 4.5005
R12151 VOUT.n165 VOUT.n109 4.5005
R12152 VOUT.n165 VOUT.n111 4.5005
R12153 VOUT.n165 VOUT.n108 4.5005
R12154 VOUT.n165 VOUT.n112 4.5005
R12155 VOUT.n165 VOUT.n107 4.5005
R12156 VOUT.n165 VOUT.t116 4.5005
R12157 VOUT.n165 VOUT.n106 4.5005
R12158 VOUT.n165 VOUT.n113 4.5005
R12159 VOUT.n163 VOUT.n109 4.5005
R12160 VOUT.n163 VOUT.n111 4.5005
R12161 VOUT.n163 VOUT.n108 4.5005
R12162 VOUT.n163 VOUT.n112 4.5005
R12163 VOUT.n163 VOUT.n107 4.5005
R12164 VOUT.n163 VOUT.t116 4.5005
R12165 VOUT.n163 VOUT.n106 4.5005
R12166 VOUT.n163 VOUT.n113 4.5005
R12167 VOUT.n163 VOUT.n162 4.5005
R12168 VOUT.n145 VOUT.n109 4.5005
R12169 VOUT.n145 VOUT.n111 4.5005
R12170 VOUT.n145 VOUT.n108 4.5005
R12171 VOUT.n145 VOUT.n112 4.5005
R12172 VOUT.n145 VOUT.n107 4.5005
R12173 VOUT.n145 VOUT.t116 4.5005
R12174 VOUT.n145 VOUT.n106 4.5005
R12175 VOUT.n145 VOUT.n113 4.5005
R12176 VOUT.n162 VOUT.n145 4.5005
R12177 VOUT.n117 VOUT.n109 4.5005
R12178 VOUT.n117 VOUT.n111 4.5005
R12179 VOUT.n117 VOUT.n108 4.5005
R12180 VOUT.n117 VOUT.n112 4.5005
R12181 VOUT.n117 VOUT.n107 4.5005
R12182 VOUT.n117 VOUT.t116 4.5005
R12183 VOUT.n117 VOUT.n106 4.5005
R12184 VOUT.n117 VOUT.n113 4.5005
R12185 VOUT.n162 VOUT.n117 4.5005
R12186 VOUT.n147 VOUT.n109 4.5005
R12187 VOUT.n147 VOUT.n111 4.5005
R12188 VOUT.n147 VOUT.n108 4.5005
R12189 VOUT.n147 VOUT.n112 4.5005
R12190 VOUT.n147 VOUT.n107 4.5005
R12191 VOUT.n147 VOUT.t116 4.5005
R12192 VOUT.n147 VOUT.n106 4.5005
R12193 VOUT.n147 VOUT.n113 4.5005
R12194 VOUT.n162 VOUT.n147 4.5005
R12195 VOUT.n116 VOUT.n109 4.5005
R12196 VOUT.n116 VOUT.n111 4.5005
R12197 VOUT.n116 VOUT.n108 4.5005
R12198 VOUT.n116 VOUT.n112 4.5005
R12199 VOUT.n116 VOUT.n107 4.5005
R12200 VOUT.n116 VOUT.t116 4.5005
R12201 VOUT.n116 VOUT.n106 4.5005
R12202 VOUT.n116 VOUT.n113 4.5005
R12203 VOUT.n162 VOUT.n116 4.5005
R12204 VOUT.n161 VOUT.n109 4.5005
R12205 VOUT.n161 VOUT.n111 4.5005
R12206 VOUT.n161 VOUT.n108 4.5005
R12207 VOUT.n161 VOUT.n112 4.5005
R12208 VOUT.n161 VOUT.n107 4.5005
R12209 VOUT.n161 VOUT.t116 4.5005
R12210 VOUT.n161 VOUT.n106 4.5005
R12211 VOUT.n161 VOUT.n113 4.5005
R12212 VOUT.n162 VOUT.n161 4.5005
R12213 VOUT.n160 VOUT.n45 4.5005
R12214 VOUT.n61 VOUT.n45 4.5005
R12215 VOUT.n56 VOUT.n40 4.5005
R12216 VOUT.n56 VOUT.n42 4.5005
R12217 VOUT.n56 VOUT.n39 4.5005
R12218 VOUT.n56 VOUT.n43 4.5005
R12219 VOUT.n56 VOUT.n38 4.5005
R12220 VOUT.n56 VOUT.t112 4.5005
R12221 VOUT.n56 VOUT.n37 4.5005
R12222 VOUT.n56 VOUT.n44 4.5005
R12223 VOUT.n56 VOUT.n45 4.5005
R12224 VOUT.n54 VOUT.n40 4.5005
R12225 VOUT.n54 VOUT.n42 4.5005
R12226 VOUT.n54 VOUT.n39 4.5005
R12227 VOUT.n54 VOUT.n43 4.5005
R12228 VOUT.n54 VOUT.n38 4.5005
R12229 VOUT.n54 VOUT.t112 4.5005
R12230 VOUT.n54 VOUT.n37 4.5005
R12231 VOUT.n54 VOUT.n44 4.5005
R12232 VOUT.n54 VOUT.n45 4.5005
R12233 VOUT.n53 VOUT.n40 4.5005
R12234 VOUT.n53 VOUT.n42 4.5005
R12235 VOUT.n53 VOUT.n39 4.5005
R12236 VOUT.n53 VOUT.n43 4.5005
R12237 VOUT.n53 VOUT.n38 4.5005
R12238 VOUT.n53 VOUT.t112 4.5005
R12239 VOUT.n53 VOUT.n37 4.5005
R12240 VOUT.n53 VOUT.n44 4.5005
R12241 VOUT.n53 VOUT.n45 4.5005
R12242 VOUT.n182 VOUT.n40 4.5005
R12243 VOUT.n182 VOUT.n42 4.5005
R12244 VOUT.n182 VOUT.n39 4.5005
R12245 VOUT.n182 VOUT.n43 4.5005
R12246 VOUT.n182 VOUT.n38 4.5005
R12247 VOUT.n182 VOUT.t112 4.5005
R12248 VOUT.n182 VOUT.n37 4.5005
R12249 VOUT.n182 VOUT.n44 4.5005
R12250 VOUT.n182 VOUT.n45 4.5005
R12251 VOUT.n180 VOUT.n40 4.5005
R12252 VOUT.n180 VOUT.n42 4.5005
R12253 VOUT.n180 VOUT.n39 4.5005
R12254 VOUT.n180 VOUT.n43 4.5005
R12255 VOUT.n180 VOUT.n38 4.5005
R12256 VOUT.n180 VOUT.t112 4.5005
R12257 VOUT.n180 VOUT.n37 4.5005
R12258 VOUT.n180 VOUT.n44 4.5005
R12259 VOUT.n178 VOUT.n40 4.5005
R12260 VOUT.n178 VOUT.n42 4.5005
R12261 VOUT.n178 VOUT.n39 4.5005
R12262 VOUT.n178 VOUT.n43 4.5005
R12263 VOUT.n178 VOUT.n38 4.5005
R12264 VOUT.n178 VOUT.t112 4.5005
R12265 VOUT.n178 VOUT.n37 4.5005
R12266 VOUT.n178 VOUT.n44 4.5005
R12267 VOUT.n64 VOUT.n40 4.5005
R12268 VOUT.n64 VOUT.n42 4.5005
R12269 VOUT.n64 VOUT.n39 4.5005
R12270 VOUT.n64 VOUT.n43 4.5005
R12271 VOUT.n64 VOUT.n38 4.5005
R12272 VOUT.n64 VOUT.t112 4.5005
R12273 VOUT.n64 VOUT.n37 4.5005
R12274 VOUT.n64 VOUT.n44 4.5005
R12275 VOUT.n64 VOUT.n45 4.5005
R12276 VOUT.n63 VOUT.n40 4.5005
R12277 VOUT.n63 VOUT.n42 4.5005
R12278 VOUT.n63 VOUT.n39 4.5005
R12279 VOUT.n63 VOUT.n43 4.5005
R12280 VOUT.n63 VOUT.n38 4.5005
R12281 VOUT.n63 VOUT.t112 4.5005
R12282 VOUT.n63 VOUT.n37 4.5005
R12283 VOUT.n63 VOUT.n44 4.5005
R12284 VOUT.n63 VOUT.n45 4.5005
R12285 VOUT.n67 VOUT.n40 4.5005
R12286 VOUT.n67 VOUT.n42 4.5005
R12287 VOUT.n67 VOUT.n39 4.5005
R12288 VOUT.n67 VOUT.n43 4.5005
R12289 VOUT.n67 VOUT.n38 4.5005
R12290 VOUT.n67 VOUT.t112 4.5005
R12291 VOUT.n67 VOUT.n37 4.5005
R12292 VOUT.n67 VOUT.n44 4.5005
R12293 VOUT.n67 VOUT.n45 4.5005
R12294 VOUT.n66 VOUT.n40 4.5005
R12295 VOUT.n66 VOUT.n42 4.5005
R12296 VOUT.n66 VOUT.n39 4.5005
R12297 VOUT.n66 VOUT.n43 4.5005
R12298 VOUT.n66 VOUT.n38 4.5005
R12299 VOUT.n66 VOUT.t112 4.5005
R12300 VOUT.n66 VOUT.n37 4.5005
R12301 VOUT.n66 VOUT.n44 4.5005
R12302 VOUT.n66 VOUT.n45 4.5005
R12303 VOUT.n49 VOUT.n40 4.5005
R12304 VOUT.n49 VOUT.n42 4.5005
R12305 VOUT.n49 VOUT.n39 4.5005
R12306 VOUT.n49 VOUT.n43 4.5005
R12307 VOUT.n49 VOUT.n38 4.5005
R12308 VOUT.n49 VOUT.t112 4.5005
R12309 VOUT.n49 VOUT.n37 4.5005
R12310 VOUT.n49 VOUT.n44 4.5005
R12311 VOUT.n49 VOUT.n45 4.5005
R12312 VOUT.n185 VOUT.n40 4.5005
R12313 VOUT.n185 VOUT.n42 4.5005
R12314 VOUT.n185 VOUT.n39 4.5005
R12315 VOUT.n185 VOUT.n43 4.5005
R12316 VOUT.n185 VOUT.n38 4.5005
R12317 VOUT.n185 VOUT.t112 4.5005
R12318 VOUT.n185 VOUT.n37 4.5005
R12319 VOUT.n185 VOUT.n44 4.5005
R12320 VOUT.n185 VOUT.n45 4.5005
R12321 VOUT.n219 VOUT.t62 4.06363
R12322 VOUT.n219 VOUT.t0 4.06363
R12323 VOUT.n217 VOUT.t2 4.06363
R12324 VOUT.n217 VOUT.t15 4.06363
R12325 VOUT.n215 VOUT.t52 4.06363
R12326 VOUT.n215 VOUT.t13 4.06363
R12327 VOUT.n213 VOUT.t40 4.06363
R12328 VOUT.n213 VOUT.t28 4.06363
R12329 VOUT.n211 VOUT.t47 4.06363
R12330 VOUT.n211 VOUT.t24 4.06363
R12331 VOUT.n210 VOUT.t42 4.06363
R12332 VOUT.n210 VOUT.t51 4.06363
R12333 VOUT.n207 VOUT.t14 4.06363
R12334 VOUT.n207 VOUT.t56 4.06363
R12335 VOUT.n205 VOUT.t17 4.06363
R12336 VOUT.n205 VOUT.t25 4.06363
R12337 VOUT.n203 VOUT.t43 4.06363
R12338 VOUT.n203 VOUT.t71 4.06363
R12339 VOUT.n201 VOUT.t9 4.06363
R12340 VOUT.n201 VOUT.t23 4.06363
R12341 VOUT.n199 VOUT.t39 4.06363
R12342 VOUT.n199 VOUT.t30 4.06363
R12343 VOUT.n198 VOUT.t21 4.06363
R12344 VOUT.n198 VOUT.t54 4.06363
R12345 VOUT.n196 VOUT.t20 4.06363
R12346 VOUT.n196 VOUT.t10 4.06363
R12347 VOUT.n194 VOUT.t26 4.06363
R12348 VOUT.n194 VOUT.t32 4.06363
R12349 VOUT.n192 VOUT.t53 4.06363
R12350 VOUT.n192 VOUT.t70 4.06363
R12351 VOUT.n190 VOUT.t16 4.06363
R12352 VOUT.n190 VOUT.t58 4.06363
R12353 VOUT.n188 VOUT.t31 4.06363
R12354 VOUT.n188 VOUT.t68 4.06363
R12355 VOUT.n187 VOUT.t7 4.06363
R12356 VOUT.n187 VOUT.t37 4.06363
R12357 VOUT.n23 VOUT.t5 4.06363
R12358 VOUT.n23 VOUT.t38 4.06363
R12359 VOUT.n24 VOUT.t46 4.06363
R12360 VOUT.n24 VOUT.t63 4.06363
R12361 VOUT.n26 VOUT.t61 4.06363
R12362 VOUT.n26 VOUT.t4 4.06363
R12363 VOUT.n28 VOUT.t64 4.06363
R12364 VOUT.n28 VOUT.t65 4.06363
R12365 VOUT.n30 VOUT.t12 4.06363
R12366 VOUT.n30 VOUT.t8 4.06363
R12367 VOUT.n32 VOUT.t59 4.06363
R12368 VOUT.n32 VOUT.t41 4.06363
R12369 VOUT.n11 VOUT.t36 4.06363
R12370 VOUT.n11 VOUT.t57 4.06363
R12371 VOUT.n12 VOUT.t69 4.06363
R12372 VOUT.n12 VOUT.t3 4.06363
R12373 VOUT.n14 VOUT.t44 4.06363
R12374 VOUT.n14 VOUT.t48 4.06363
R12375 VOUT.n16 VOUT.t11 4.06363
R12376 VOUT.n16 VOUT.t67 4.06363
R12377 VOUT.n18 VOUT.t49 4.06363
R12378 VOUT.n18 VOUT.t50 4.06363
R12379 VOUT.n20 VOUT.t33 4.06363
R12380 VOUT.n20 VOUT.t45 4.06363
R12381 VOUT.n0 VOUT.t35 4.06363
R12382 VOUT.n0 VOUT.t60 4.06363
R12383 VOUT.n1 VOUT.t66 4.06363
R12384 VOUT.n1 VOUT.t18 4.06363
R12385 VOUT.n3 VOUT.t1 4.06363
R12386 VOUT.n3 VOUT.t29 4.06363
R12387 VOUT.n5 VOUT.t22 4.06363
R12388 VOUT.n5 VOUT.t55 4.06363
R12389 VOUT.n7 VOUT.t19 4.06363
R12390 VOUT.n7 VOUT.t34 4.06363
R12391 VOUT.n9 VOUT.t6 4.06363
R12392 VOUT.n9 VOUT.t27 4.06363
R12393 VOUT.n186 VOUT 3.7135
R12394 VOUT.n263 VOUT.n262 3.60085
R12395 VOUT.n262 VOUT.n242 3.02103
R12396 VOUT.n239 VOUT.t79 2.82907
R12397 VOUT.n239 VOUT.t78 2.82907
R12398 VOUT.n237 VOUT.t109 2.82907
R12399 VOUT.n237 VOUT.t106 2.82907
R12400 VOUT.n235 VOUT.t100 2.82907
R12401 VOUT.n235 VOUT.t98 2.82907
R12402 VOUT.n233 VOUT.t73 2.82907
R12403 VOUT.n233 VOUT.t77 2.82907
R12404 VOUT.n232 VOUT.t94 2.82907
R12405 VOUT.n232 VOUT.t76 2.82907
R12406 VOUT.n230 VOUT.t96 2.82907
R12407 VOUT.n230 VOUT.t95 2.82907
R12408 VOUT.n228 VOUT.t85 2.82907
R12409 VOUT.n228 VOUT.t83 2.82907
R12410 VOUT.n226 VOUT.t74 2.82907
R12411 VOUT.n226 VOUT.t72 2.82907
R12412 VOUT.n224 VOUT.t91 2.82907
R12413 VOUT.n224 VOUT.t92 2.82907
R12414 VOUT.n223 VOUT.t111 2.82907
R12415 VOUT.n223 VOUT.t93 2.82907
R12416 VOUT.n252 VOUT.t87 2.82907
R12417 VOUT.n252 VOUT.t80 2.82907
R12418 VOUT.n253 VOUT.t88 2.82907
R12419 VOUT.n253 VOUT.t101 2.82907
R12420 VOUT.n255 VOUT.t107 2.82907
R12421 VOUT.n255 VOUT.t110 2.82907
R12422 VOUT.n257 VOUT.t90 2.82907
R12423 VOUT.n257 VOUT.t82 2.82907
R12424 VOUT.n259 VOUT.t102 2.82907
R12425 VOUT.n259 VOUT.t89 2.82907
R12426 VOUT.n243 VOUT.t103 2.82907
R12427 VOUT.n243 VOUT.t97 2.82907
R12428 VOUT.n244 VOUT.t104 2.82907
R12429 VOUT.n244 VOUT.t75 2.82907
R12430 VOUT.n246 VOUT.t84 2.82907
R12431 VOUT.n246 VOUT.t86 2.82907
R12432 VOUT.n248 VOUT.t108 2.82907
R12433 VOUT.n248 VOUT.t99 2.82907
R12434 VOUT.n250 VOUT.t81 2.82907
R12435 VOUT.n250 VOUT.t105 2.82907
R12436 VOUT.n222 VOUT.n35 2.74718
R12437 VOUT.n221 VOUT.n209 2.33778
R12438 VOUT.n34 VOUT.n22 2.33778
R12439 VOUT.n126 VOUT.n124 2.251
R12440 VOUT.n126 VOUT.n123 2.251
R12441 VOUT.n126 VOUT.n122 2.251
R12442 VOUT.n126 VOUT.n121 2.251
R12443 VOUT.n95 VOUT.n94 2.251
R12444 VOUT.n95 VOUT.n93 2.251
R12445 VOUT.n95 VOUT.n92 2.251
R12446 VOUT.n95 VOUT.n91 2.251
R12447 VOUT.n168 VOUT.n167 2.251
R12448 VOUT.n133 VOUT.n131 2.251
R12449 VOUT.n133 VOUT.n130 2.251
R12450 VOUT.n133 VOUT.n129 2.251
R12451 VOUT.n151 VOUT.n133 2.251
R12452 VOUT.n139 VOUT.n138 2.251
R12453 VOUT.n139 VOUT.n137 2.251
R12454 VOUT.n139 VOUT.n136 2.251
R12455 VOUT.n139 VOUT.n135 2.251
R12456 VOUT.n165 VOUT.n105 2.251
R12457 VOUT.n160 VOUT.n158 2.251
R12458 VOUT.n160 VOUT.n157 2.251
R12459 VOUT.n160 VOUT.n156 2.251
R12460 VOUT.n160 VOUT.n155 2.251
R12461 VOUT.n61 VOUT.n60 2.251
R12462 VOUT.n61 VOUT.n59 2.251
R12463 VOUT.n61 VOUT.n58 2.251
R12464 VOUT.n61 VOUT.n57 2.251
R12465 VOUT.n178 VOUT.n177 2.251
R12466 VOUT.n95 VOUT.n75 2.2505
R12467 VOUT.n90 VOUT.n75 2.2505
R12468 VOUT.n88 VOUT.n75 2.2505
R12469 VOUT.n87 VOUT.n75 2.2505
R12470 VOUT.n172 VOUT.n75 2.2505
R12471 VOUT.n170 VOUT.n75 2.2505
R12472 VOUT.n168 VOUT.n75 2.2505
R12473 VOUT.n98 VOUT.n75 2.2505
R12474 VOUT.n97 VOUT.n75 2.2505
R12475 VOUT.n101 VOUT.n75 2.2505
R12476 VOUT.n100 VOUT.n75 2.2505
R12477 VOUT.n83 VOUT.n75 2.2505
R12478 VOUT.n175 VOUT.n75 2.2505
R12479 VOUT.n175 VOUT.n174 2.2505
R12480 VOUT.n139 VOUT.n110 2.2505
R12481 VOUT.n120 VOUT.n110 2.2505
R12482 VOUT.n141 VOUT.n110 2.2505
R12483 VOUT.n119 VOUT.n110 2.2505
R12484 VOUT.n143 VOUT.n110 2.2505
R12485 VOUT.n110 VOUT.n104 2.2505
R12486 VOUT.n165 VOUT.n110 2.2505
R12487 VOUT.n163 VOUT.n110 2.2505
R12488 VOUT.n145 VOUT.n110 2.2505
R12489 VOUT.n117 VOUT.n110 2.2505
R12490 VOUT.n147 VOUT.n110 2.2505
R12491 VOUT.n116 VOUT.n110 2.2505
R12492 VOUT.n161 VOUT.n110 2.2505
R12493 VOUT.n161 VOUT.n114 2.2505
R12494 VOUT.n61 VOUT.n41 2.2505
R12495 VOUT.n56 VOUT.n41 2.2505
R12496 VOUT.n54 VOUT.n41 2.2505
R12497 VOUT.n53 VOUT.n41 2.2505
R12498 VOUT.n182 VOUT.n41 2.2505
R12499 VOUT.n180 VOUT.n41 2.2505
R12500 VOUT.n178 VOUT.n41 2.2505
R12501 VOUT.n64 VOUT.n41 2.2505
R12502 VOUT.n63 VOUT.n41 2.2505
R12503 VOUT.n67 VOUT.n41 2.2505
R12504 VOUT.n66 VOUT.n41 2.2505
R12505 VOUT.n49 VOUT.n41 2.2505
R12506 VOUT.n185 VOUT.n41 2.2505
R12507 VOUT.n185 VOUT.n184 2.2505
R12508 VOUT.n103 VOUT.n96 2.25024
R12509 VOUT.n103 VOUT.n89 2.25024
R12510 VOUT.n171 VOUT.n103 2.25024
R12511 VOUT.n103 VOUT.n99 2.25024
R12512 VOUT.n103 VOUT.n102 2.25024
R12513 VOUT.n103 VOUT.n70 2.25024
R12514 VOUT.n153 VOUT.n150 2.25024
R12515 VOUT.n153 VOUT.n149 2.25024
R12516 VOUT.n153 VOUT.n148 2.25024
R12517 VOUT.n153 VOUT.n115 2.25024
R12518 VOUT.n153 VOUT.n152 2.25024
R12519 VOUT.n154 VOUT.n153 2.25024
R12520 VOUT.n69 VOUT.n62 2.25024
R12521 VOUT.n69 VOUT.n55 2.25024
R12522 VOUT.n181 VOUT.n69 2.25024
R12523 VOUT.n69 VOUT.n65 2.25024
R12524 VOUT.n69 VOUT.n68 2.25024
R12525 VOUT.n69 VOUT.n36 2.25024
R12526 VOUT.n170 VOUT.n80 1.50111
R12527 VOUT.n118 VOUT.n104 1.50111
R12528 VOUT.n180 VOUT.n46 1.50111
R12529 VOUT.n126 VOUT.n125 1.501
R12530 VOUT.n133 VOUT.n132 1.501
R12531 VOUT.n160 VOUT.n159 1.501
R12532 VOUT.n174 VOUT.n85 1.12536
R12533 VOUT.n174 VOUT.n86 1.12536
R12534 VOUT.n174 VOUT.n173 1.12536
R12535 VOUT.n134 VOUT.n114 1.12536
R12536 VOUT.n140 VOUT.n114 1.12536
R12537 VOUT.n142 VOUT.n114 1.12536
R12538 VOUT.n184 VOUT.n51 1.12536
R12539 VOUT.n184 VOUT.n52 1.12536
R12540 VOUT.n184 VOUT.n183 1.12536
R12541 VOUT.n174 VOUT.n81 1.12536
R12542 VOUT.n174 VOUT.n82 1.12536
R12543 VOUT.n174 VOUT.n84 1.12536
R12544 VOUT.n164 VOUT.n114 1.12536
R12545 VOUT.n144 VOUT.n114 1.12536
R12546 VOUT.n146 VOUT.n114 1.12536
R12547 VOUT.n184 VOUT.n47 1.12536
R12548 VOUT.n184 VOUT.n48 1.12536
R12549 VOUT.n184 VOUT.n50 1.12536
R12550 VOUT.n236 VOUT.n234 1.00481
R12551 VOUT.n238 VOUT.n236 1.00481
R12552 VOUT.n240 VOUT.n238 1.00481
R12553 VOUT.n227 VOUT.n225 1.00481
R12554 VOUT.n229 VOUT.n227 1.00481
R12555 VOUT.n231 VOUT.n229 1.00481
R12556 VOUT.n260 VOUT.n258 1.00481
R12557 VOUT.n258 VOUT.n256 1.00481
R12558 VOUT.n256 VOUT.n254 1.00481
R12559 VOUT.n251 VOUT.n249 1.00481
R12560 VOUT.n249 VOUT.n247 1.00481
R12561 VOUT.n247 VOUT.n245 1.00481
R12562 VOUT.n214 VOUT.n212 0.573776
R12563 VOUT.n216 VOUT.n214 0.573776
R12564 VOUT.n218 VOUT.n216 0.573776
R12565 VOUT.n220 VOUT.n218 0.573776
R12566 VOUT.n202 VOUT.n200 0.573776
R12567 VOUT.n204 VOUT.n202 0.573776
R12568 VOUT.n206 VOUT.n204 0.573776
R12569 VOUT.n208 VOUT.n206 0.573776
R12570 VOUT.n191 VOUT.n189 0.573776
R12571 VOUT.n193 VOUT.n191 0.573776
R12572 VOUT.n195 VOUT.n193 0.573776
R12573 VOUT.n197 VOUT.n195 0.573776
R12574 VOUT.n33 VOUT.n31 0.573776
R12575 VOUT.n31 VOUT.n29 0.573776
R12576 VOUT.n29 VOUT.n27 0.573776
R12577 VOUT.n27 VOUT.n25 0.573776
R12578 VOUT.n21 VOUT.n19 0.573776
R12579 VOUT.n19 VOUT.n17 0.573776
R12580 VOUT.n17 VOUT.n15 0.573776
R12581 VOUT.n15 VOUT.n13 0.573776
R12582 VOUT.n10 VOUT.n8 0.573776
R12583 VOUT.n8 VOUT.n6 0.573776
R12584 VOUT.n6 VOUT.n4 0.573776
R12585 VOUT.n4 VOUT.n2 0.573776
R12586 VOUT.n186 VOUT.n185 0.365565
R12587 VOUT.n263 VOUT.n186 0.3624
R12588 VOUT.n128 VOUT.n127 0.0910737
R12589 VOUT.n179 VOUT.n176 0.0723685
R12590 VOUT.n133 VOUT.n128 0.0522944
R12591 VOUT.n176 VOUT.n175 0.0499135
R12592 VOUT.n127 VOUT.n126 0.0499135
R12593 VOUT.n161 VOUT.n160 0.0464294
R12594 VOUT.n169 VOUT.n166 0.0391444
R12595 VOUT.n128 VOUT.t113 0.023435
R12596 VOUT.n176 VOUT.t115 0.02262
R12597 VOUT.n127 VOUT.t114 0.02262
R12598 VOUT VOUT.n263 0.0099
R12599 VOUT.n98 VOUT.n81 0.00365111
R12600 VOUT.n101 VOUT.n82 0.00365111
R12601 VOUT.n84 VOUT.n83 0.00365111
R12602 VOUT.n126 VOUT.n85 0.00365111
R12603 VOUT.n90 VOUT.n86 0.00365111
R12604 VOUT.n173 VOUT.n87 0.00365111
R12605 VOUT.n164 VOUT.n163 0.00365111
R12606 VOUT.n144 VOUT.n117 0.00365111
R12607 VOUT.n146 VOUT.n116 0.00365111
R12608 VOUT.n134 VOUT.n133 0.00365111
R12609 VOUT.n140 VOUT.n120 0.00365111
R12610 VOUT.n142 VOUT.n119 0.00365111
R12611 VOUT.n64 VOUT.n47 0.00365111
R12612 VOUT.n67 VOUT.n48 0.00365111
R12613 VOUT.n50 VOUT.n49 0.00365111
R12614 VOUT.n160 VOUT.n51 0.00365111
R12615 VOUT.n56 VOUT.n52 0.00365111
R12616 VOUT.n183 VOUT.n53 0.00365111
R12617 VOUT.n95 VOUT.n85 0.00340054
R12618 VOUT.n88 VOUT.n86 0.00340054
R12619 VOUT.n173 VOUT.n172 0.00340054
R12620 VOUT.n168 VOUT.n81 0.00340054
R12621 VOUT.n97 VOUT.n82 0.00340054
R12622 VOUT.n100 VOUT.n84 0.00340054
R12623 VOUT.n139 VOUT.n134 0.00340054
R12624 VOUT.n141 VOUT.n140 0.00340054
R12625 VOUT.n143 VOUT.n142 0.00340054
R12626 VOUT.n165 VOUT.n164 0.00340054
R12627 VOUT.n145 VOUT.n144 0.00340054
R12628 VOUT.n147 VOUT.n146 0.00340054
R12629 VOUT.n61 VOUT.n51 0.00340054
R12630 VOUT.n54 VOUT.n52 0.00340054
R12631 VOUT.n183 VOUT.n182 0.00340054
R12632 VOUT.n178 VOUT.n47 0.00340054
R12633 VOUT.n63 VOUT.n48 0.00340054
R12634 VOUT.n66 VOUT.n50 0.00340054
R12635 VOUT.n96 VOUT.n90 0.00252698
R12636 VOUT.n89 VOUT.n87 0.00252698
R12637 VOUT.n171 VOUT.n170 0.00252698
R12638 VOUT.n99 VOUT.n97 0.00252698
R12639 VOUT.n102 VOUT.n100 0.00252698
R12640 VOUT.n175 VOUT.n70 0.00252698
R12641 VOUT.n96 VOUT.n95 0.00252698
R12642 VOUT.n89 VOUT.n88 0.00252698
R12643 VOUT.n172 VOUT.n171 0.00252698
R12644 VOUT.n99 VOUT.n98 0.00252698
R12645 VOUT.n102 VOUT.n101 0.00252698
R12646 VOUT.n83 VOUT.n70 0.00252698
R12647 VOUT.n150 VOUT.n120 0.00252698
R12648 VOUT.n149 VOUT.n119 0.00252698
R12649 VOUT.n148 VOUT.n104 0.00252698
R12650 VOUT.n145 VOUT.n115 0.00252698
R12651 VOUT.n152 VOUT.n147 0.00252698
R12652 VOUT.n161 VOUT.n154 0.00252698
R12653 VOUT.n150 VOUT.n139 0.00252698
R12654 VOUT.n149 VOUT.n141 0.00252698
R12655 VOUT.n148 VOUT.n143 0.00252698
R12656 VOUT.n163 VOUT.n115 0.00252698
R12657 VOUT.n152 VOUT.n117 0.00252698
R12658 VOUT.n154 VOUT.n116 0.00252698
R12659 VOUT.n62 VOUT.n56 0.00252698
R12660 VOUT.n55 VOUT.n53 0.00252698
R12661 VOUT.n181 VOUT.n180 0.00252698
R12662 VOUT.n65 VOUT.n63 0.00252698
R12663 VOUT.n68 VOUT.n66 0.00252698
R12664 VOUT.n185 VOUT.n36 0.00252698
R12665 VOUT.n62 VOUT.n61 0.00252698
R12666 VOUT.n55 VOUT.n54 0.00252698
R12667 VOUT.n182 VOUT.n181 0.00252698
R12668 VOUT.n65 VOUT.n64 0.00252698
R12669 VOUT.n68 VOUT.n67 0.00252698
R12670 VOUT.n49 VOUT.n36 0.00252698
R12671 VOUT.n170 VOUT.n169 0.0020275
R12672 VOUT.n169 VOUT.n168 0.0020275
R12673 VOUT.n166 VOUT.n104 0.0020275
R12674 VOUT.n166 VOUT.n165 0.0020275
R12675 VOUT.n180 VOUT.n179 0.0020275
R12676 VOUT.n179 VOUT.n178 0.0020275
R12677 VOUT.n80 VOUT.n79 0.00166668
R12678 VOUT.n162 VOUT.n118 0.00166668
R12679 VOUT.n46 VOUT.n45 0.00166668
R12680 VOUT.n184 VOUT.n46 0.00133328
R12681 VOUT.n118 VOUT.n114 0.00133328
R12682 VOUT.n174 VOUT.n80 0.00133328
R12683 VOUT.n177 VOUT.n69 0.001
R12684 VOUT.n155 VOUT.n69 0.001
R12685 VOUT.n57 VOUT.n37 0.001
R12686 VOUT.n156 VOUT.n37 0.001
R12687 VOUT.n58 VOUT.n38 0.001
R12688 VOUT.n157 VOUT.n38 0.001
R12689 VOUT.n59 VOUT.n39 0.001
R12690 VOUT.n158 VOUT.n39 0.001
R12691 VOUT.n60 VOUT.n40 0.001
R12692 VOUT.n159 VOUT.n40 0.001
R12693 VOUT.n153 VOUT.n105 0.001
R12694 VOUT.n153 VOUT.n151 0.001
R12695 VOUT.n135 VOUT.n106 0.001
R12696 VOUT.n129 VOUT.n106 0.001
R12697 VOUT.n136 VOUT.n107 0.001
R12698 VOUT.n130 VOUT.n107 0.001
R12699 VOUT.n137 VOUT.n108 0.001
R12700 VOUT.n131 VOUT.n108 0.001
R12701 VOUT.n138 VOUT.n109 0.001
R12702 VOUT.n132 VOUT.n109 0.001
R12703 VOUT.n167 VOUT.n103 0.001
R12704 VOUT.n121 VOUT.n103 0.001
R12705 VOUT.n91 VOUT.n71 0.001
R12706 VOUT.n122 VOUT.n71 0.001
R12707 VOUT.n92 VOUT.n72 0.001
R12708 VOUT.n123 VOUT.n72 0.001
R12709 VOUT.n93 VOUT.n73 0.001
R12710 VOUT.n124 VOUT.n73 0.001
R12711 VOUT.n94 VOUT.n74 0.001
R12712 VOUT.n125 VOUT.n74 0.001
R12713 VOUT.n125 VOUT.n75 0.001
R12714 VOUT.n124 VOUT.n76 0.001
R12715 VOUT.n123 VOUT.n77 0.001
R12716 VOUT.n122 VOUT.t117 0.001
R12717 VOUT.n121 VOUT.n78 0.001
R12718 VOUT.n94 VOUT.n76 0.001
R12719 VOUT.n93 VOUT.n77 0.001
R12720 VOUT.n92 VOUT.t117 0.001
R12721 VOUT.n91 VOUT.n78 0.001
R12722 VOUT.n167 VOUT.n79 0.001
R12723 VOUT.n132 VOUT.n110 0.001
R12724 VOUT.n131 VOUT.n111 0.001
R12725 VOUT.n130 VOUT.n112 0.001
R12726 VOUT.n129 VOUT.t116 0.001
R12727 VOUT.n151 VOUT.n113 0.001
R12728 VOUT.n138 VOUT.n111 0.001
R12729 VOUT.n137 VOUT.n112 0.001
R12730 VOUT.n136 VOUT.t116 0.001
R12731 VOUT.n135 VOUT.n113 0.001
R12732 VOUT.n162 VOUT.n105 0.001
R12733 VOUT.n159 VOUT.n41 0.001
R12734 VOUT.n158 VOUT.n42 0.001
R12735 VOUT.n157 VOUT.n43 0.001
R12736 VOUT.n156 VOUT.t112 0.001
R12737 VOUT.n155 VOUT.n44 0.001
R12738 VOUT.n60 VOUT.n42 0.001
R12739 VOUT.n59 VOUT.n43 0.001
R12740 VOUT.n58 VOUT.t112 0.001
R12741 VOUT.n57 VOUT.n44 0.001
R12742 VOUT.n177 VOUT.n45 0.001
R12743 VDD.n290 VDD.n254 756.745
R12744 VDD.n239 VDD.n203 756.745
R12745 VDD.n196 VDD.n160 756.745
R12746 VDD.n145 VDD.n109 756.745
R12747 VDD.n103 VDD.n67 756.745
R12748 VDD.n52 VDD.n16 756.745
R12749 VDD.n1779 VDD.n1743 756.745
R12750 VDD.n1830 VDD.n1794 756.745
R12751 VDD.n1685 VDD.n1649 756.745
R12752 VDD.n1736 VDD.n1700 756.745
R12753 VDD.n1592 VDD.n1556 756.745
R12754 VDD.n1643 VDD.n1607 756.745
R12755 VDD.n291 VDD.n290 585
R12756 VDD.n289 VDD.n256 585
R12757 VDD.n288 VDD.n287 585
R12758 VDD.n259 VDD.n257 585
R12759 VDD.n282 VDD.n281 585
R12760 VDD.n280 VDD.n279 585
R12761 VDD.n263 VDD.n262 585
R12762 VDD.n274 VDD.n273 585
R12763 VDD.n272 VDD.n271 585
R12764 VDD.n267 VDD.n266 585
R12765 VDD.n240 VDD.n239 585
R12766 VDD.n238 VDD.n205 585
R12767 VDD.n237 VDD.n236 585
R12768 VDD.n208 VDD.n206 585
R12769 VDD.n231 VDD.n230 585
R12770 VDD.n229 VDD.n228 585
R12771 VDD.n212 VDD.n211 585
R12772 VDD.n223 VDD.n222 585
R12773 VDD.n221 VDD.n220 585
R12774 VDD.n216 VDD.n215 585
R12775 VDD.n197 VDD.n196 585
R12776 VDD.n195 VDD.n162 585
R12777 VDD.n194 VDD.n193 585
R12778 VDD.n165 VDD.n163 585
R12779 VDD.n188 VDD.n187 585
R12780 VDD.n186 VDD.n185 585
R12781 VDD.n169 VDD.n168 585
R12782 VDD.n180 VDD.n179 585
R12783 VDD.n178 VDD.n177 585
R12784 VDD.n173 VDD.n172 585
R12785 VDD.n146 VDD.n145 585
R12786 VDD.n144 VDD.n111 585
R12787 VDD.n143 VDD.n142 585
R12788 VDD.n114 VDD.n112 585
R12789 VDD.n137 VDD.n136 585
R12790 VDD.n135 VDD.n134 585
R12791 VDD.n118 VDD.n117 585
R12792 VDD.n129 VDD.n128 585
R12793 VDD.n127 VDD.n126 585
R12794 VDD.n122 VDD.n121 585
R12795 VDD.n104 VDD.n103 585
R12796 VDD.n102 VDD.n69 585
R12797 VDD.n101 VDD.n100 585
R12798 VDD.n72 VDD.n70 585
R12799 VDD.n95 VDD.n94 585
R12800 VDD.n93 VDD.n92 585
R12801 VDD.n76 VDD.n75 585
R12802 VDD.n87 VDD.n86 585
R12803 VDD.n85 VDD.n84 585
R12804 VDD.n80 VDD.n79 585
R12805 VDD.n53 VDD.n52 585
R12806 VDD.n51 VDD.n18 585
R12807 VDD.n50 VDD.n49 585
R12808 VDD.n21 VDD.n19 585
R12809 VDD.n44 VDD.n43 585
R12810 VDD.n42 VDD.n41 585
R12811 VDD.n25 VDD.n24 585
R12812 VDD.n36 VDD.n35 585
R12813 VDD.n34 VDD.n33 585
R12814 VDD.n29 VDD.n28 585
R12815 VDD.n1780 VDD.n1779 585
R12816 VDD.n1778 VDD.n1745 585
R12817 VDD.n1777 VDD.n1776 585
R12818 VDD.n1748 VDD.n1746 585
R12819 VDD.n1771 VDD.n1770 585
R12820 VDD.n1769 VDD.n1768 585
R12821 VDD.n1752 VDD.n1751 585
R12822 VDD.n1763 VDD.n1762 585
R12823 VDD.n1761 VDD.n1760 585
R12824 VDD.n1756 VDD.n1755 585
R12825 VDD.n1831 VDD.n1830 585
R12826 VDD.n1829 VDD.n1796 585
R12827 VDD.n1828 VDD.n1827 585
R12828 VDD.n1799 VDD.n1797 585
R12829 VDD.n1822 VDD.n1821 585
R12830 VDD.n1820 VDD.n1819 585
R12831 VDD.n1803 VDD.n1802 585
R12832 VDD.n1814 VDD.n1813 585
R12833 VDD.n1812 VDD.n1811 585
R12834 VDD.n1807 VDD.n1806 585
R12835 VDD.n1686 VDD.n1685 585
R12836 VDD.n1684 VDD.n1651 585
R12837 VDD.n1683 VDD.n1682 585
R12838 VDD.n1654 VDD.n1652 585
R12839 VDD.n1677 VDD.n1676 585
R12840 VDD.n1675 VDD.n1674 585
R12841 VDD.n1658 VDD.n1657 585
R12842 VDD.n1669 VDD.n1668 585
R12843 VDD.n1667 VDD.n1666 585
R12844 VDD.n1662 VDD.n1661 585
R12845 VDD.n1737 VDD.n1736 585
R12846 VDD.n1735 VDD.n1702 585
R12847 VDD.n1734 VDD.n1733 585
R12848 VDD.n1705 VDD.n1703 585
R12849 VDD.n1728 VDD.n1727 585
R12850 VDD.n1726 VDD.n1725 585
R12851 VDD.n1709 VDD.n1708 585
R12852 VDD.n1720 VDD.n1719 585
R12853 VDD.n1718 VDD.n1717 585
R12854 VDD.n1713 VDD.n1712 585
R12855 VDD.n1593 VDD.n1592 585
R12856 VDD.n1591 VDD.n1558 585
R12857 VDD.n1590 VDD.n1589 585
R12858 VDD.n1561 VDD.n1559 585
R12859 VDD.n1584 VDD.n1583 585
R12860 VDD.n1582 VDD.n1581 585
R12861 VDD.n1565 VDD.n1564 585
R12862 VDD.n1576 VDD.n1575 585
R12863 VDD.n1574 VDD.n1573 585
R12864 VDD.n1569 VDD.n1568 585
R12865 VDD.n1644 VDD.n1643 585
R12866 VDD.n1642 VDD.n1609 585
R12867 VDD.n1641 VDD.n1640 585
R12868 VDD.n1612 VDD.n1610 585
R12869 VDD.n1635 VDD.n1634 585
R12870 VDD.n1633 VDD.n1632 585
R12871 VDD.n1616 VDD.n1615 585
R12872 VDD.n1627 VDD.n1626 585
R12873 VDD.n1625 VDD.n1624 585
R12874 VDD.n1620 VDD.n1619 585
R12875 VDD.n3214 VDD.n653 475.611
R12876 VDD.n432 VDD.n357 475.611
R12877 VDD.n3345 VDD.n359 475.611
R12878 VDD.n3217 VDD.n655 475.611
R12879 VDD.n2114 VDD.n1115 475.611
R12880 VDD.n2117 VDD.n2116 475.611
R12881 VDD.n1468 VDD.n1238 475.611
R12882 VDD.n1471 VDD.n1236 475.611
R12883 VDD.n1240 VDD.t13 395.726
R12884 VDD.n1265 VDD.t42 395.726
R12885 VDD.n1290 VDD.t56 395.726
R12886 VDD.n1101 VDD.t53 395.726
R12887 VDD.n1992 VDD.t25 395.726
R12888 VDD.n1952 VDD.t36 395.726
R12889 VDD.n392 VDD.t39 395.726
R12890 VDD.n406 VDD.t17 395.726
R12891 VDD.n418 VDD.t33 395.726
R12892 VDD.n733 VDD.t2 395.726
R12893 VDD.n3175 VDD.t10 395.726
R12894 VDD.n658 VDD.t69 395.726
R12895 VDD.n1082 VDD.t6 347.526
R12896 VDD.n933 VDD.t29 347.526
R12897 VDD.n1075 VDD.t63 347.526
R12898 VDD.n943 VDD.t72 347.526
R12899 VDD.n801 VDD.t21 347.526
R12900 VDD.n2608 VDD.t59 347.526
R12901 VDD.n785 VDD.t49 347.526
R12902 VDD.n2614 VDD.t66 347.526
R12903 VDD.n755 VDD.t75 347.526
R12904 VDD.n1043 VDD.t45 347.526
R12905 VDD.n1240 VDD.t16 329.483
R12906 VDD.n1265 VDD.t44 329.483
R12907 VDD.n1290 VDD.t58 329.483
R12908 VDD.n1101 VDD.t54 329.483
R12909 VDD.n1992 VDD.t27 329.483
R12910 VDD.n1952 VDD.t37 329.483
R12911 VDD.n392 VDD.t40 329.483
R12912 VDD.n406 VDD.t19 329.483
R12913 VDD.n418 VDD.t34 329.483
R12914 VDD.n733 VDD.t5 329.483
R12915 VDD.n3175 VDD.t12 329.483
R12916 VDD.n658 VDD.t71 329.483
R12917 VDD.n268 VDD.t149 329.043
R12918 VDD.n217 VDD.t160 329.043
R12919 VDD.n174 VDD.t138 329.043
R12920 VDD.n123 VDD.t148 329.043
R12921 VDD.n81 VDD.t128 329.043
R12922 VDD.n30 VDD.t177 329.043
R12923 VDD.n1757 VDD.t185 329.043
R12924 VDD.n1808 VDD.t176 329.043
R12925 VDD.n1663 VDD.t174 329.043
R12926 VDD.n1714 VDD.t167 329.043
R12927 VDD.n1570 VDD.t153 329.043
R12928 VDD.n1621 VDD.t102 329.043
R12929 VDD.n1241 VDD.t15 303.69
R12930 VDD.n1266 VDD.t43 303.69
R12931 VDD.n1291 VDD.t57 303.69
R12932 VDD.n1102 VDD.t55 303.69
R12933 VDD.n1993 VDD.t28 303.69
R12934 VDD.n1953 VDD.t38 303.69
R12935 VDD.n393 VDD.t41 303.69
R12936 VDD.n407 VDD.t20 303.69
R12937 VDD.n419 VDD.t35 303.69
R12938 VDD.n734 VDD.t4 303.69
R12939 VDD.n3176 VDD.t11 303.69
R12940 VDD.n659 VDD.t70 303.69
R12941 VDD.n3052 VDD.n765 294.147
R12942 VDD.n3004 VDD.n762 294.147
R12943 VDD.n2675 VDD.n2592 294.147
R12944 VDD.n2848 VDD.n902 294.147
R12945 VDD.n2531 VDD.n941 294.147
R12946 VDD.n2480 VDD.n2479 294.147
R12947 VDD.n2305 VDD.n1060 294.147
R12948 VDD.n2356 VDD.n1062 294.147
R12949 VDD.n2983 VDD.n763 294.147
R12950 VDD.n3055 VDD.n3054 294.147
R12951 VDD.n2794 VDD.n2593 294.147
R12952 VDD.n2846 VDD.n2595 294.147
R12953 VDD.n2589 VDD.n930 294.147
R12954 VDD.n2538 VDD.n929 294.147
R12955 VDD.n2188 VDD.n1061 294.147
R12956 VDD.n2358 VDD.n1058 294.147
R12957 VDD.n1082 VDD.t9 293.986
R12958 VDD.n933 VDD.t31 293.986
R12959 VDD.n1075 VDD.t65 293.986
R12960 VDD.n943 VDD.t73 293.986
R12961 VDD.n801 VDD.t23 293.986
R12962 VDD.n801 VDD.t24 293.986
R12963 VDD.n2608 VDD.t62 293.986
R12964 VDD.n785 VDD.t51 293.986
R12965 VDD.n2614 VDD.t68 293.986
R12966 VDD.n755 VDD.t76 293.986
R12967 VDD.n1043 VDD.t47 293.986
R12968 VDD.n1043 VDD.t48 293.986
R12969 VDD.n1083 VDD.t8 268.192
R12970 VDD.n934 VDD.t32 268.192
R12971 VDD.n1076 VDD.t64 268.192
R12972 VDD.n944 VDD.t74 268.192
R12973 VDD.n2609 VDD.t61 268.192
R12974 VDD.n786 VDD.t52 268.192
R12975 VDD.n2615 VDD.t67 268.192
R12976 VDD.n756 VDD.t77 268.192
R12977 VDD.n2985 VDD.n763 185
R12978 VDD.n3053 VDD.n763 185
R12979 VDD.n2987 VDD.n2986 185
R12980 VDD.n2986 VDD.n761 185
R12981 VDD.n2988 VDD.n792 185
R12982 VDD.n2998 VDD.n792 185
R12983 VDD.n2989 VDD.n800 185
R12984 VDD.n800 VDD.n790 185
R12985 VDD.n2991 VDD.n2990 185
R12986 VDD.n2992 VDD.n2991 185
R12987 VDD.n2953 VDD.n799 185
R12988 VDD.n799 VDD.n796 185
R12989 VDD.n2951 VDD.n2950 185
R12990 VDD.n2950 VDD.n2949 185
R12991 VDD.n803 VDD.n802 185
R12992 VDD.n804 VDD.n803 185
R12993 VDD.n2942 VDD.n2941 185
R12994 VDD.n2943 VDD.n2942 185
R12995 VDD.n2940 VDD.n813 185
R12996 VDD.n813 VDD.n810 185
R12997 VDD.n2939 VDD.n2938 185
R12998 VDD.n2938 VDD.n2937 185
R12999 VDD.n815 VDD.n814 185
R13000 VDD.n823 VDD.n815 185
R13001 VDD.n2930 VDD.n2929 185
R13002 VDD.n2931 VDD.n2930 185
R13003 VDD.n2928 VDD.n824 185
R13004 VDD.n829 VDD.n824 185
R13005 VDD.n2927 VDD.n2926 185
R13006 VDD.n2926 VDD.n2925 185
R13007 VDD.n826 VDD.n825 185
R13008 VDD.n835 VDD.n826 185
R13009 VDD.n2918 VDD.n2917 185
R13010 VDD.n2919 VDD.n2918 185
R13011 VDD.n2916 VDD.n836 185
R13012 VDD.n841 VDD.n836 185
R13013 VDD.n2915 VDD.n2914 185
R13014 VDD.n2914 VDD.n2913 185
R13015 VDD.n838 VDD.n837 185
R13016 VDD.n847 VDD.n838 185
R13017 VDD.n2906 VDD.n2905 185
R13018 VDD.n2907 VDD.n2906 185
R13019 VDD.n2904 VDD.n848 185
R13020 VDD.n2759 VDD.n848 185
R13021 VDD.n2903 VDD.n2902 185
R13022 VDD.n2902 VDD.n2901 185
R13023 VDD.n850 VDD.n849 185
R13024 VDD.n851 VDD.n850 185
R13025 VDD.n2894 VDD.n2893 185
R13026 VDD.n2895 VDD.n2894 185
R13027 VDD.n2892 VDD.n859 185
R13028 VDD.n2768 VDD.n859 185
R13029 VDD.n2891 VDD.n2890 185
R13030 VDD.n2890 VDD.n2889 185
R13031 VDD.n861 VDD.n860 185
R13032 VDD.n862 VDD.n861 185
R13033 VDD.n2882 VDD.n2881 185
R13034 VDD.n2883 VDD.n2882 185
R13035 VDD.n2880 VDD.n871 185
R13036 VDD.n871 VDD.n868 185
R13037 VDD.n2879 VDD.n2878 185
R13038 VDD.n2878 VDD.n2877 185
R13039 VDD.n873 VDD.n872 185
R13040 VDD.n882 VDD.n873 185
R13041 VDD.n2870 VDD.n2869 185
R13042 VDD.n2871 VDD.n2870 185
R13043 VDD.n2868 VDD.n883 185
R13044 VDD.n883 VDD.n879 185
R13045 VDD.n2867 VDD.n2866 185
R13046 VDD.n2866 VDD.n2865 185
R13047 VDD.n885 VDD.n884 185
R13048 VDD.n893 VDD.n885 185
R13049 VDD.n2858 VDD.n2857 185
R13050 VDD.n2859 VDD.n2858 185
R13051 VDD.n2856 VDD.n894 185
R13052 VDD.n899 VDD.n894 185
R13053 VDD.n2855 VDD.n2854 185
R13054 VDD.n2854 VDD.n2853 185
R13055 VDD.n896 VDD.n895 185
R13056 VDD.n2594 VDD.n896 185
R13057 VDD.n2846 VDD.n2845 185
R13058 VDD.n2847 VDD.n2846 185
R13059 VDD.n2844 VDD.n2595 185
R13060 VDD.n2843 VDD.n2842 185
R13061 VDD.n2840 VDD.n2596 185
R13062 VDD.n2838 VDD.n2837 185
R13063 VDD.n2836 VDD.n2597 185
R13064 VDD.n2835 VDD.n2834 185
R13065 VDD.n2832 VDD.n2598 185
R13066 VDD.n2830 VDD.n2829 185
R13067 VDD.n2828 VDD.n2599 185
R13068 VDD.n2827 VDD.n2826 185
R13069 VDD.n2824 VDD.n2600 185
R13070 VDD.n2822 VDD.n2821 185
R13071 VDD.n2820 VDD.n2601 185
R13072 VDD.n2819 VDD.n2818 185
R13073 VDD.n2816 VDD.n2602 185
R13074 VDD.n2814 VDD.n2813 185
R13075 VDD.n2812 VDD.n2603 185
R13076 VDD.n2811 VDD.n2810 185
R13077 VDD.n2808 VDD.n2604 185
R13078 VDD.n2806 VDD.n2805 185
R13079 VDD.n2804 VDD.n2605 185
R13080 VDD.n2803 VDD.n2802 185
R13081 VDD.n2800 VDD.n2606 185
R13082 VDD.n2798 VDD.n2797 185
R13083 VDD.n2796 VDD.n2607 185
R13084 VDD.n2795 VDD.n2794 185
R13085 VDD.n3056 VDD.n3055 185
R13086 VDD.n3057 VDD.n754 185
R13087 VDD.n3059 VDD.n3058 185
R13088 VDD.n3061 VDD.n752 185
R13089 VDD.n3063 VDD.n3062 185
R13090 VDD.n3064 VDD.n751 185
R13091 VDD.n3066 VDD.n3065 185
R13092 VDD.n3068 VDD.n749 185
R13093 VDD.n3070 VDD.n3069 185
R13094 VDD.n3071 VDD.n748 185
R13095 VDD.n3073 VDD.n3072 185
R13096 VDD.n3075 VDD.n746 185
R13097 VDD.n3077 VDD.n3076 185
R13098 VDD.n2962 VDD.n745 185
R13099 VDD.n2964 VDD.n2963 185
R13100 VDD.n2966 VDD.n2960 185
R13101 VDD.n2968 VDD.n2967 185
R13102 VDD.n2969 VDD.n2959 185
R13103 VDD.n2971 VDD.n2970 185
R13104 VDD.n2973 VDD.n2957 185
R13105 VDD.n2975 VDD.n2974 185
R13106 VDD.n2976 VDD.n2956 185
R13107 VDD.n2978 VDD.n2977 185
R13108 VDD.n2980 VDD.n2955 185
R13109 VDD.n2981 VDD.n2954 185
R13110 VDD.n2984 VDD.n2983 185
R13111 VDD.n3054 VDD.n758 185
R13112 VDD.n3054 VDD.n3053 185
R13113 VDD.n2728 VDD.n760 185
R13114 VDD.n761 VDD.n760 185
R13115 VDD.n2729 VDD.n791 185
R13116 VDD.n2998 VDD.n791 185
R13117 VDD.n2731 VDD.n2730 185
R13118 VDD.n2730 VDD.n790 185
R13119 VDD.n2732 VDD.n798 185
R13120 VDD.n2992 VDD.n798 185
R13121 VDD.n2734 VDD.n2733 185
R13122 VDD.n2733 VDD.n796 185
R13123 VDD.n2735 VDD.n806 185
R13124 VDD.n2949 VDD.n806 185
R13125 VDD.n2737 VDD.n2736 185
R13126 VDD.n2736 VDD.n804 185
R13127 VDD.n2738 VDD.n812 185
R13128 VDD.n2943 VDD.n812 185
R13129 VDD.n2740 VDD.n2739 185
R13130 VDD.n2739 VDD.n810 185
R13131 VDD.n2741 VDD.n817 185
R13132 VDD.n2937 VDD.n817 185
R13133 VDD.n2743 VDD.n2742 185
R13134 VDD.n2742 VDD.n823 185
R13135 VDD.n2744 VDD.n822 185
R13136 VDD.n2931 VDD.n822 185
R13137 VDD.n2746 VDD.n2745 185
R13138 VDD.n2745 VDD.n829 185
R13139 VDD.n2747 VDD.n828 185
R13140 VDD.n2925 VDD.n828 185
R13141 VDD.n2749 VDD.n2748 185
R13142 VDD.n2748 VDD.n835 185
R13143 VDD.n2750 VDD.n834 185
R13144 VDD.n2919 VDD.n834 185
R13145 VDD.n2752 VDD.n2751 185
R13146 VDD.n2751 VDD.n841 185
R13147 VDD.n2753 VDD.n840 185
R13148 VDD.n2913 VDD.n840 185
R13149 VDD.n2755 VDD.n2754 185
R13150 VDD.n2754 VDD.n847 185
R13151 VDD.n2756 VDD.n846 185
R13152 VDD.n2907 VDD.n846 185
R13153 VDD.n2758 VDD.n2757 185
R13154 VDD.n2759 VDD.n2758 185
R13155 VDD.n2727 VDD.n853 185
R13156 VDD.n2901 VDD.n853 185
R13157 VDD.n2726 VDD.n2725 185
R13158 VDD.n2725 VDD.n851 185
R13159 VDD.n2611 VDD.n858 185
R13160 VDD.n2895 VDD.n858 185
R13161 VDD.n2770 VDD.n2769 185
R13162 VDD.n2769 VDD.n2768 185
R13163 VDD.n2771 VDD.n864 185
R13164 VDD.n2889 VDD.n864 185
R13165 VDD.n2773 VDD.n2772 185
R13166 VDD.n2772 VDD.n862 185
R13167 VDD.n2774 VDD.n870 185
R13168 VDD.n2883 VDD.n870 185
R13169 VDD.n2776 VDD.n2775 185
R13170 VDD.n2775 VDD.n868 185
R13171 VDD.n2777 VDD.n875 185
R13172 VDD.n2877 VDD.n875 185
R13173 VDD.n2779 VDD.n2778 185
R13174 VDD.n2778 VDD.n882 185
R13175 VDD.n2780 VDD.n881 185
R13176 VDD.n2871 VDD.n881 185
R13177 VDD.n2782 VDD.n2781 185
R13178 VDD.n2781 VDD.n879 185
R13179 VDD.n2783 VDD.n887 185
R13180 VDD.n2865 VDD.n887 185
R13181 VDD.n2785 VDD.n2784 185
R13182 VDD.n2784 VDD.n893 185
R13183 VDD.n2786 VDD.n892 185
R13184 VDD.n2859 VDD.n892 185
R13185 VDD.n2788 VDD.n2787 185
R13186 VDD.n2787 VDD.n899 185
R13187 VDD.n2789 VDD.n898 185
R13188 VDD.n2853 VDD.n898 185
R13189 VDD.n2791 VDD.n2790 185
R13190 VDD.n2790 VDD.n2594 185
R13191 VDD.n2792 VDD.n2593 185
R13192 VDD.n2847 VDD.n2593 185
R13193 VDD.n2533 VDD.n941 185
R13194 VDD.n941 VDD.n903 185
R13195 VDD.n2535 VDD.n2534 185
R13196 VDD.n2536 VDD.n2535 185
R13197 VDD.n942 VDD.n940 185
R13198 VDD.n2474 VDD.n940 185
R13199 VDD.n2464 VDD.n955 185
R13200 VDD.n955 VDD.n947 185
R13201 VDD.n2466 VDD.n2465 185
R13202 VDD.n2467 VDD.n2466 185
R13203 VDD.n2463 VDD.n954 185
R13204 VDD.n954 VDD.n951 185
R13205 VDD.n2462 VDD.n2461 185
R13206 VDD.n2461 VDD.n2460 185
R13207 VDD.n957 VDD.n956 185
R13208 VDD.n958 VDD.n957 185
R13209 VDD.n2453 VDD.n2452 185
R13210 VDD.n2454 VDD.n2453 185
R13211 VDD.n2451 VDD.n967 185
R13212 VDD.n967 VDD.n964 185
R13213 VDD.n2450 VDD.n2449 185
R13214 VDD.n2449 VDD.n2448 185
R13215 VDD.n969 VDD.n968 185
R13216 VDD.n978 VDD.n969 185
R13217 VDD.n2441 VDD.n2440 185
R13218 VDD.n2442 VDD.n2441 185
R13219 VDD.n2439 VDD.n979 185
R13220 VDD.n979 VDD.n975 185
R13221 VDD.n2438 VDD.n2437 185
R13222 VDD.n2437 VDD.n2436 185
R13223 VDD.n981 VDD.n980 185
R13224 VDD.n2261 VDD.n981 185
R13225 VDD.n2429 VDD.n2428 185
R13226 VDD.n2430 VDD.n2429 185
R13227 VDD.n2427 VDD.n990 185
R13228 VDD.n990 VDD.n987 185
R13229 VDD.n2426 VDD.n2425 185
R13230 VDD.n2425 VDD.n2424 185
R13231 VDD.n992 VDD.n991 185
R13232 VDD.n2270 VDD.n992 185
R13233 VDD.n2417 VDD.n2416 185
R13234 VDD.n2418 VDD.n2417 185
R13235 VDD.n2415 VDD.n1001 185
R13236 VDD.n1001 VDD.n998 185
R13237 VDD.n2414 VDD.n2413 185
R13238 VDD.n2413 VDD.n2412 185
R13239 VDD.n1003 VDD.n1002 185
R13240 VDD.n1004 VDD.n1003 185
R13241 VDD.n2405 VDD.n2404 185
R13242 VDD.n2406 VDD.n2405 185
R13243 VDD.n2403 VDD.n1013 185
R13244 VDD.n1013 VDD.n1010 185
R13245 VDD.n2402 VDD.n2401 185
R13246 VDD.n2401 VDD.n2400 185
R13247 VDD.n1015 VDD.n1014 185
R13248 VDD.n1016 VDD.n1015 185
R13249 VDD.n2393 VDD.n2392 185
R13250 VDD.n2394 VDD.n2393 185
R13251 VDD.n2391 VDD.n1025 185
R13252 VDD.n1025 VDD.n1022 185
R13253 VDD.n2390 VDD.n2389 185
R13254 VDD.n2389 VDD.n2388 185
R13255 VDD.n1027 VDD.n1026 185
R13256 VDD.n1028 VDD.n1027 185
R13257 VDD.n2381 VDD.n2380 185
R13258 VDD.n2382 VDD.n2381 185
R13259 VDD.n2379 VDD.n1037 185
R13260 VDD.n1037 VDD.n1034 185
R13261 VDD.n2378 VDD.n2377 185
R13262 VDD.n2377 VDD.n2376 185
R13263 VDD.n1039 VDD.n1038 185
R13264 VDD.n1048 VDD.n1039 185
R13265 VDD.n2368 VDD.n2367 185
R13266 VDD.n2369 VDD.n2368 185
R13267 VDD.n2366 VDD.n1049 185
R13268 VDD.n1055 VDD.n1049 185
R13269 VDD.n2365 VDD.n2364 185
R13270 VDD.n2364 VDD.n2363 185
R13271 VDD.n1051 VDD.n1050 185
R13272 VDD.n1052 VDD.n1051 185
R13273 VDD.n2356 VDD.n2355 185
R13274 VDD.n2357 VDD.n2356 185
R13275 VDD.n2354 VDD.n1062 185
R13276 VDD.n2353 VDD.n2352 185
R13277 VDD.n2350 VDD.n1063 185
R13278 VDD.n2350 VDD.n1059 185
R13279 VDD.n2349 VDD.n2348 185
R13280 VDD.n2347 VDD.n2346 185
R13281 VDD.n2345 VDD.n1065 185
R13282 VDD.n2343 VDD.n2342 185
R13283 VDD.n2341 VDD.n1066 185
R13284 VDD.n2340 VDD.n2339 185
R13285 VDD.n2337 VDD.n1067 185
R13286 VDD.n2335 VDD.n2334 185
R13287 VDD.n2333 VDD.n1068 185
R13288 VDD.n2332 VDD.n2331 185
R13289 VDD.n2329 VDD.n2328 185
R13290 VDD.n2327 VDD.n2326 185
R13291 VDD.n2325 VDD.n1071 185
R13292 VDD.n2323 VDD.n2322 185
R13293 VDD.n2321 VDD.n1072 185
R13294 VDD.n2320 VDD.n2319 185
R13295 VDD.n2317 VDD.n1073 185
R13296 VDD.n2315 VDD.n2314 185
R13297 VDD.n2313 VDD.n1074 185
R13298 VDD.n2312 VDD.n2311 185
R13299 VDD.n2309 VDD.n2308 185
R13300 VDD.n2307 VDD.n2306 185
R13301 VDD.n2305 VDD.n2304 185
R13302 VDD.n2305 VDD.n1059 185
R13303 VDD.n2481 VDD.n2480 185
R13304 VDD.n2483 VDD.n2482 185
R13305 VDD.n2485 VDD.n2484 185
R13306 VDD.n2488 VDD.n2487 185
R13307 VDD.n2490 VDD.n2489 185
R13308 VDD.n2492 VDD.n2491 185
R13309 VDD.n2494 VDD.n2493 185
R13310 VDD.n2496 VDD.n2495 185
R13311 VDD.n2498 VDD.n2497 185
R13312 VDD.n2500 VDD.n2499 185
R13313 VDD.n2502 VDD.n2501 185
R13314 VDD.n2504 VDD.n2503 185
R13315 VDD.n2506 VDD.n2505 185
R13316 VDD.n2508 VDD.n2507 185
R13317 VDD.n2510 VDD.n2509 185
R13318 VDD.n2512 VDD.n2511 185
R13319 VDD.n2514 VDD.n2513 185
R13320 VDD.n2516 VDD.n2515 185
R13321 VDD.n2518 VDD.n2517 185
R13322 VDD.n2520 VDD.n2519 185
R13323 VDD.n2522 VDD.n2521 185
R13324 VDD.n2524 VDD.n2523 185
R13325 VDD.n2526 VDD.n2525 185
R13326 VDD.n2528 VDD.n2527 185
R13327 VDD.n2530 VDD.n2529 185
R13328 VDD.n2532 VDD.n2531 185
R13329 VDD.n2479 VDD.n2478 185
R13330 VDD.n2479 VDD.n903 185
R13331 VDD.n2477 VDD.n938 185
R13332 VDD.n2536 VDD.n938 185
R13333 VDD.n2476 VDD.n2475 185
R13334 VDD.n2475 VDD.n2474 185
R13335 VDD.n946 VDD.n945 185
R13336 VDD.n947 VDD.n946 185
R13337 VDD.n2243 VDD.n952 185
R13338 VDD.n2467 VDD.n952 185
R13339 VDD.n2245 VDD.n2244 185
R13340 VDD.n2244 VDD.n951 185
R13341 VDD.n2246 VDD.n959 185
R13342 VDD.n2460 VDD.n959 185
R13343 VDD.n2248 VDD.n2247 185
R13344 VDD.n2247 VDD.n958 185
R13345 VDD.n2249 VDD.n965 185
R13346 VDD.n2454 VDD.n965 185
R13347 VDD.n2251 VDD.n2250 185
R13348 VDD.n2250 VDD.n964 185
R13349 VDD.n2252 VDD.n970 185
R13350 VDD.n2448 VDD.n970 185
R13351 VDD.n2254 VDD.n2253 185
R13352 VDD.n2253 VDD.n978 185
R13353 VDD.n2255 VDD.n976 185
R13354 VDD.n2442 VDD.n976 185
R13355 VDD.n2257 VDD.n2256 185
R13356 VDD.n2256 VDD.n975 185
R13357 VDD.n2258 VDD.n982 185
R13358 VDD.n2436 VDD.n982 185
R13359 VDD.n2260 VDD.n2259 185
R13360 VDD.n2261 VDD.n2260 185
R13361 VDD.n2242 VDD.n988 185
R13362 VDD.n2430 VDD.n988 185
R13363 VDD.n2241 VDD.n2240 185
R13364 VDD.n2240 VDD.n987 185
R13365 VDD.n1079 VDD.n993 185
R13366 VDD.n2424 VDD.n993 185
R13367 VDD.n2272 VDD.n2271 185
R13368 VDD.n2271 VDD.n2270 185
R13369 VDD.n2273 VDD.n999 185
R13370 VDD.n2418 VDD.n999 185
R13371 VDD.n2275 VDD.n2274 185
R13372 VDD.n2274 VDD.n998 185
R13373 VDD.n2276 VDD.n1005 185
R13374 VDD.n2412 VDD.n1005 185
R13375 VDD.n2278 VDD.n2277 185
R13376 VDD.n2277 VDD.n1004 185
R13377 VDD.n2279 VDD.n1011 185
R13378 VDD.n2406 VDD.n1011 185
R13379 VDD.n2281 VDD.n2280 185
R13380 VDD.n2280 VDD.n1010 185
R13381 VDD.n2282 VDD.n1017 185
R13382 VDD.n2400 VDD.n1017 185
R13383 VDD.n2284 VDD.n2283 185
R13384 VDD.n2283 VDD.n1016 185
R13385 VDD.n2285 VDD.n1023 185
R13386 VDD.n2394 VDD.n1023 185
R13387 VDD.n2287 VDD.n2286 185
R13388 VDD.n2286 VDD.n1022 185
R13389 VDD.n2288 VDD.n1029 185
R13390 VDD.n2388 VDD.n1029 185
R13391 VDD.n2290 VDD.n2289 185
R13392 VDD.n2289 VDD.n1028 185
R13393 VDD.n2291 VDD.n1035 185
R13394 VDD.n2382 VDD.n1035 185
R13395 VDD.n2293 VDD.n2292 185
R13396 VDD.n2292 VDD.n1034 185
R13397 VDD.n2294 VDD.n1040 185
R13398 VDD.n2376 VDD.n1040 185
R13399 VDD.n2296 VDD.n2295 185
R13400 VDD.n2295 VDD.n1048 185
R13401 VDD.n2297 VDD.n1046 185
R13402 VDD.n2369 VDD.n1046 185
R13403 VDD.n2299 VDD.n2298 185
R13404 VDD.n2298 VDD.n1055 185
R13405 VDD.n2300 VDD.n1053 185
R13406 VDD.n2363 VDD.n1053 185
R13407 VDD.n2302 VDD.n2301 185
R13408 VDD.n2301 VDD.n1052 185
R13409 VDD.n2303 VDD.n1060 185
R13410 VDD.n2357 VDD.n1060 185
R13411 VDD.n3052 VDD.n3051 185
R13412 VDD.n3053 VDD.n3052 185
R13413 VDD.n766 VDD.n764 185
R13414 VDD.n764 VDD.n761 185
R13415 VDD.n2997 VDD.n2996 185
R13416 VDD.n2998 VDD.n2997 185
R13417 VDD.n2995 VDD.n793 185
R13418 VDD.n793 VDD.n790 185
R13419 VDD.n2994 VDD.n2993 185
R13420 VDD.n2993 VDD.n2992 185
R13421 VDD.n795 VDD.n794 185
R13422 VDD.n796 VDD.n795 185
R13423 VDD.n2948 VDD.n2947 185
R13424 VDD.n2949 VDD.n2948 185
R13425 VDD.n2946 VDD.n807 185
R13426 VDD.n807 VDD.n804 185
R13427 VDD.n2945 VDD.n2944 185
R13428 VDD.n2944 VDD.n2943 185
R13429 VDD.n809 VDD.n808 185
R13430 VDD.n810 VDD.n809 185
R13431 VDD.n2936 VDD.n2935 185
R13432 VDD.n2937 VDD.n2936 185
R13433 VDD.n2934 VDD.n818 185
R13434 VDD.n823 VDD.n818 185
R13435 VDD.n2933 VDD.n2932 185
R13436 VDD.n2932 VDD.n2931 185
R13437 VDD.n820 VDD.n819 185
R13438 VDD.n829 VDD.n820 185
R13439 VDD.n2924 VDD.n2923 185
R13440 VDD.n2925 VDD.n2924 185
R13441 VDD.n2922 VDD.n830 185
R13442 VDD.n835 VDD.n830 185
R13443 VDD.n2921 VDD.n2920 185
R13444 VDD.n2920 VDD.n2919 185
R13445 VDD.n832 VDD.n831 185
R13446 VDD.n841 VDD.n832 185
R13447 VDD.n2912 VDD.n2911 185
R13448 VDD.n2913 VDD.n2912 185
R13449 VDD.n2910 VDD.n842 185
R13450 VDD.n847 VDD.n842 185
R13451 VDD.n2909 VDD.n2908 185
R13452 VDD.n2908 VDD.n2907 185
R13453 VDD.n844 VDD.n843 185
R13454 VDD.n2759 VDD.n844 185
R13455 VDD.n2900 VDD.n2899 185
R13456 VDD.n2901 VDD.n2900 185
R13457 VDD.n2898 VDD.n854 185
R13458 VDD.n854 VDD.n851 185
R13459 VDD.n2897 VDD.n2896 185
R13460 VDD.n2896 VDD.n2895 185
R13461 VDD.n856 VDD.n855 185
R13462 VDD.n2768 VDD.n856 185
R13463 VDD.n2888 VDD.n2887 185
R13464 VDD.n2889 VDD.n2888 185
R13465 VDD.n2886 VDD.n865 185
R13466 VDD.n865 VDD.n862 185
R13467 VDD.n2885 VDD.n2884 185
R13468 VDD.n2884 VDD.n2883 185
R13469 VDD.n867 VDD.n866 185
R13470 VDD.n868 VDD.n867 185
R13471 VDD.n2876 VDD.n2875 185
R13472 VDD.n2877 VDD.n2876 185
R13473 VDD.n2874 VDD.n876 185
R13474 VDD.n882 VDD.n876 185
R13475 VDD.n2873 VDD.n2872 185
R13476 VDD.n2872 VDD.n2871 185
R13477 VDD.n878 VDD.n877 185
R13478 VDD.n879 VDD.n878 185
R13479 VDD.n2864 VDD.n2863 185
R13480 VDD.n2865 VDD.n2864 185
R13481 VDD.n2862 VDD.n888 185
R13482 VDD.n893 VDD.n888 185
R13483 VDD.n2861 VDD.n2860 185
R13484 VDD.n2860 VDD.n2859 185
R13485 VDD.n890 VDD.n889 185
R13486 VDD.n899 VDD.n890 185
R13487 VDD.n2852 VDD.n2851 185
R13488 VDD.n2853 VDD.n2852 185
R13489 VDD.n2850 VDD.n900 185
R13490 VDD.n2594 VDD.n900 185
R13491 VDD.n2849 VDD.n2848 185
R13492 VDD.n2848 VDD.n2847 185
R13493 VDD.n902 VDD.n901 185
R13494 VDD.n2628 VDD.n2627 185
R13495 VDD.n2629 VDD.n2625 185
R13496 VDD.n2625 VDD.n2591 185
R13497 VDD.n2631 VDD.n2630 185
R13498 VDD.n2633 VDD.n2624 185
R13499 VDD.n2636 VDD.n2635 185
R13500 VDD.n2637 VDD.n2623 185
R13501 VDD.n2639 VDD.n2638 185
R13502 VDD.n2641 VDD.n2622 185
R13503 VDD.n2644 VDD.n2643 185
R13504 VDD.n2645 VDD.n2621 185
R13505 VDD.n2647 VDD.n2646 185
R13506 VDD.n2649 VDD.n2620 185
R13507 VDD.n2652 VDD.n2651 185
R13508 VDD.n2653 VDD.n2619 185
R13509 VDD.n2655 VDD.n2654 185
R13510 VDD.n2657 VDD.n2618 185
R13511 VDD.n2660 VDD.n2659 185
R13512 VDD.n2661 VDD.n2617 185
R13513 VDD.n2663 VDD.n2662 185
R13514 VDD.n2665 VDD.n2616 185
R13515 VDD.n2668 VDD.n2667 185
R13516 VDD.n2669 VDD.n2613 185
R13517 VDD.n2672 VDD.n2671 185
R13518 VDD.n2674 VDD.n2612 185
R13519 VDD.n2676 VDD.n2675 185
R13520 VDD.n2675 VDD.n2591 185
R13521 VDD.n3005 VDD.n3004 185
R13522 VDD.n3006 VDD.n784 185
R13523 VDD.n3008 VDD.n3007 185
R13524 VDD.n3010 VDD.n782 185
R13525 VDD.n3012 VDD.n3011 185
R13526 VDD.n3013 VDD.n781 185
R13527 VDD.n3015 VDD.n3014 185
R13528 VDD.n3017 VDD.n779 185
R13529 VDD.n3019 VDD.n3018 185
R13530 VDD.n3020 VDD.n778 185
R13531 VDD.n3022 VDD.n3021 185
R13532 VDD.n3024 VDD.n776 185
R13533 VDD.n3026 VDD.n3025 185
R13534 VDD.n3029 VDD.n775 185
R13535 VDD.n3031 VDD.n3030 185
R13536 VDD.n3033 VDD.n773 185
R13537 VDD.n3035 VDD.n3034 185
R13538 VDD.n3036 VDD.n772 185
R13539 VDD.n3038 VDD.n3037 185
R13540 VDD.n3040 VDD.n770 185
R13541 VDD.n3042 VDD.n3041 185
R13542 VDD.n3043 VDD.n769 185
R13543 VDD.n3045 VDD.n3044 185
R13544 VDD.n3047 VDD.n767 185
R13545 VDD.n3049 VDD.n3048 185
R13546 VDD.n3050 VDD.n765 185
R13547 VDD.n3002 VDD.n762 185
R13548 VDD.n3053 VDD.n762 185
R13549 VDD.n3001 VDD.n3000 185
R13550 VDD.n3000 VDD.n761 185
R13551 VDD.n2999 VDD.n788 185
R13552 VDD.n2999 VDD.n2998 185
R13553 VDD.n2699 VDD.n789 185
R13554 VDD.n790 VDD.n789 185
R13555 VDD.n2700 VDD.n797 185
R13556 VDD.n2992 VDD.n797 185
R13557 VDD.n2702 VDD.n2701 185
R13558 VDD.n2701 VDD.n796 185
R13559 VDD.n2703 VDD.n805 185
R13560 VDD.n2949 VDD.n805 185
R13561 VDD.n2705 VDD.n2704 185
R13562 VDD.n2704 VDD.n804 185
R13563 VDD.n2706 VDD.n811 185
R13564 VDD.n2943 VDD.n811 185
R13565 VDD.n2708 VDD.n2707 185
R13566 VDD.n2707 VDD.n810 185
R13567 VDD.n2709 VDD.n816 185
R13568 VDD.n2937 VDD.n816 185
R13569 VDD.n2711 VDD.n2710 185
R13570 VDD.n2710 VDD.n823 185
R13571 VDD.n2712 VDD.n821 185
R13572 VDD.n2931 VDD.n821 185
R13573 VDD.n2714 VDD.n2713 185
R13574 VDD.n2713 VDD.n829 185
R13575 VDD.n2715 VDD.n827 185
R13576 VDD.n2925 VDD.n827 185
R13577 VDD.n2717 VDD.n2716 185
R13578 VDD.n2716 VDD.n835 185
R13579 VDD.n2718 VDD.n833 185
R13580 VDD.n2919 VDD.n833 185
R13581 VDD.n2720 VDD.n2719 185
R13582 VDD.n2719 VDD.n841 185
R13583 VDD.n2721 VDD.n839 185
R13584 VDD.n2913 VDD.n839 185
R13585 VDD.n2723 VDD.n2722 185
R13586 VDD.n2722 VDD.n847 185
R13587 VDD.n2724 VDD.n845 185
R13588 VDD.n2907 VDD.n845 185
R13589 VDD.n2761 VDD.n2760 185
R13590 VDD.n2760 VDD.n2759 185
R13591 VDD.n2762 VDD.n852 185
R13592 VDD.n2901 VDD.n852 185
R13593 VDD.n2764 VDD.n2763 185
R13594 VDD.n2763 VDD.n851 185
R13595 VDD.n2765 VDD.n857 185
R13596 VDD.n2895 VDD.n857 185
R13597 VDD.n2767 VDD.n2766 185
R13598 VDD.n2768 VDD.n2767 185
R13599 VDD.n2698 VDD.n863 185
R13600 VDD.n2889 VDD.n863 185
R13601 VDD.n2697 VDD.n2696 185
R13602 VDD.n2696 VDD.n862 185
R13603 VDD.n2695 VDD.n869 185
R13604 VDD.n2883 VDD.n869 185
R13605 VDD.n2694 VDD.n2693 185
R13606 VDD.n2693 VDD.n868 185
R13607 VDD.n2692 VDD.n874 185
R13608 VDD.n2877 VDD.n874 185
R13609 VDD.n2691 VDD.n2690 185
R13610 VDD.n2690 VDD.n882 185
R13611 VDD.n2689 VDD.n880 185
R13612 VDD.n2871 VDD.n880 185
R13613 VDD.n2688 VDD.n2687 185
R13614 VDD.n2687 VDD.n879 185
R13615 VDD.n2686 VDD.n886 185
R13616 VDD.n2865 VDD.n886 185
R13617 VDD.n2685 VDD.n2684 185
R13618 VDD.n2684 VDD.n893 185
R13619 VDD.n2683 VDD.n891 185
R13620 VDD.n2859 VDD.n891 185
R13621 VDD.n2682 VDD.n2681 185
R13622 VDD.n2681 VDD.n899 185
R13623 VDD.n2680 VDD.n897 185
R13624 VDD.n2853 VDD.n897 185
R13625 VDD.n2679 VDD.n2678 185
R13626 VDD.n2678 VDD.n2594 185
R13627 VDD.n2677 VDD.n2592 185
R13628 VDD.n2847 VDD.n2592 185
R13629 VDD.n2114 VDD.n2113 185
R13630 VDD.n2115 VDD.n2114 185
R13631 VDD.n1116 VDD.n1114 185
R13632 VDD.n1114 VDD.n1108 185
R13633 VDD.n1917 VDD.n1916 185
R13634 VDD.n1916 VDD.n1915 185
R13635 VDD.n1119 VDD.n1118 185
R13636 VDD.n1120 VDD.n1119 185
R13637 VDD.n1905 VDD.n1904 185
R13638 VDD.n1906 VDD.n1905 185
R13639 VDD.n1129 VDD.n1128 185
R13640 VDD.n1128 VDD.n1127 185
R13641 VDD.n1900 VDD.n1899 185
R13642 VDD.n1899 VDD.n1898 185
R13643 VDD.n1132 VDD.n1131 185
R13644 VDD.n1139 VDD.n1132 185
R13645 VDD.n1889 VDD.n1888 185
R13646 VDD.n1890 VDD.n1889 185
R13647 VDD.n1141 VDD.n1140 185
R13648 VDD.n1140 VDD.n1138 185
R13649 VDD.n1884 VDD.n1883 185
R13650 VDD.n1883 VDD.n1882 185
R13651 VDD.n1144 VDD.n1143 185
R13652 VDD.n1145 VDD.n1144 185
R13653 VDD.n1873 VDD.n1872 185
R13654 VDD.n1874 VDD.n1873 185
R13655 VDD.n1153 VDD.n1152 185
R13656 VDD.n1152 VDD.n1151 185
R13657 VDD.n1868 VDD.n1867 185
R13658 VDD.n1867 VDD.n1866 185
R13659 VDD.n1156 VDD.n1155 185
R13660 VDD.n1163 VDD.n1156 185
R13661 VDD.n1857 VDD.n1856 185
R13662 VDD.n1858 VDD.n1857 185
R13663 VDD.n1165 VDD.n1164 185
R13664 VDD.n1164 VDD.n1162 185
R13665 VDD.n1852 VDD.n1851 185
R13666 VDD.n1851 VDD.n1850 185
R13667 VDD.n1168 VDD.n1167 185
R13668 VDD.n1169 VDD.n1168 185
R13669 VDD.n1841 VDD.n1840 185
R13670 VDD.n1842 VDD.n1841 185
R13671 VDD.n1177 VDD.n1176 185
R13672 VDD.n1176 VDD.n1175 185
R13673 VDD.n1554 VDD.n1553 185
R13674 VDD.n1553 VDD.n1552 185
R13675 VDD.n1180 VDD.n1179 185
R13676 VDD.n1186 VDD.n1180 185
R13677 VDD.n1543 VDD.n1542 185
R13678 VDD.n1544 VDD.n1543 185
R13679 VDD.n1188 VDD.n1187 185
R13680 VDD.n1535 VDD.n1187 185
R13681 VDD.n1538 VDD.n1537 185
R13682 VDD.n1537 VDD.n1536 185
R13683 VDD.n1191 VDD.n1190 185
R13684 VDD.n1192 VDD.n1191 185
R13685 VDD.n1526 VDD.n1525 185
R13686 VDD.n1527 VDD.n1526 185
R13687 VDD.n1200 VDD.n1199 185
R13688 VDD.n1199 VDD.n1198 185
R13689 VDD.n1521 VDD.n1520 185
R13690 VDD.n1520 VDD.n1519 185
R13691 VDD.n1203 VDD.n1202 185
R13692 VDD.n1209 VDD.n1203 185
R13693 VDD.n1510 VDD.n1509 185
R13694 VDD.n1511 VDD.n1510 185
R13695 VDD.n1211 VDD.n1210 185
R13696 VDD.n1502 VDD.n1210 185
R13697 VDD.n1505 VDD.n1504 185
R13698 VDD.n1504 VDD.n1503 185
R13699 VDD.n1214 VDD.n1213 185
R13700 VDD.n1215 VDD.n1214 185
R13701 VDD.n1493 VDD.n1492 185
R13702 VDD.n1494 VDD.n1493 185
R13703 VDD.n1223 VDD.n1222 185
R13704 VDD.n1222 VDD.n1221 185
R13705 VDD.n1488 VDD.n1487 185
R13706 VDD.n1487 VDD.n1486 185
R13707 VDD.n1226 VDD.n1225 185
R13708 VDD.n1227 VDD.n1226 185
R13709 VDD.n1477 VDD.n1476 185
R13710 VDD.n1478 VDD.n1477 185
R13711 VDD.n1234 VDD.n1233 185
R13712 VDD.n1469 VDD.n1233 185
R13713 VDD.n1472 VDD.n1471 185
R13714 VDD.n1471 VDD.n1470 185
R13715 VDD.n1308 VDD.n1236 185
R13716 VDD.n1311 VDD.n1310 185
R13717 VDD.n1307 VDD.n1306 185
R13718 VDD.n1306 VDD.n1237 185
R13719 VDD.n1316 VDD.n1315 185
R13720 VDD.n1318 VDD.n1305 185
R13721 VDD.n1321 VDD.n1320 185
R13722 VDD.n1303 VDD.n1302 185
R13723 VDD.n1326 VDD.n1325 185
R13724 VDD.n1328 VDD.n1301 185
R13725 VDD.n1331 VDD.n1330 185
R13726 VDD.n1299 VDD.n1298 185
R13727 VDD.n1336 VDD.n1335 185
R13728 VDD.n1338 VDD.n1297 185
R13729 VDD.n1341 VDD.n1340 185
R13730 VDD.n1295 VDD.n1294 185
R13731 VDD.n1348 VDD.n1347 185
R13732 VDD.n1350 VDD.n1293 185
R13733 VDD.n1351 VDD.n1292 185
R13734 VDD.n1354 VDD.n1353 185
R13735 VDD.n1355 VDD.n1289 185
R13736 VDD.n1286 VDD.n1285 185
R13737 VDD.n1360 VDD.n1359 185
R13738 VDD.n1362 VDD.n1284 185
R13739 VDD.n1365 VDD.n1364 185
R13740 VDD.n1282 VDD.n1281 185
R13741 VDD.n1370 VDD.n1369 185
R13742 VDD.n1372 VDD.n1280 185
R13743 VDD.n1375 VDD.n1374 185
R13744 VDD.n1278 VDD.n1277 185
R13745 VDD.n1380 VDD.n1379 185
R13746 VDD.n1382 VDD.n1276 185
R13747 VDD.n1385 VDD.n1384 185
R13748 VDD.n1274 VDD.n1273 185
R13749 VDD.n1390 VDD.n1389 185
R13750 VDD.n1392 VDD.n1272 185
R13751 VDD.n1395 VDD.n1394 185
R13752 VDD.n1270 VDD.n1269 185
R13753 VDD.n1402 VDD.n1401 185
R13754 VDD.n1404 VDD.n1268 185
R13755 VDD.n1405 VDD.n1267 185
R13756 VDD.n1408 VDD.n1407 185
R13757 VDD.n1409 VDD.n1264 185
R13758 VDD.n1261 VDD.n1260 185
R13759 VDD.n1414 VDD.n1413 185
R13760 VDD.n1416 VDD.n1259 185
R13761 VDD.n1419 VDD.n1418 185
R13762 VDD.n1257 VDD.n1256 185
R13763 VDD.n1424 VDD.n1423 185
R13764 VDD.n1426 VDD.n1255 185
R13765 VDD.n1429 VDD.n1428 185
R13766 VDD.n1253 VDD.n1252 185
R13767 VDD.n1434 VDD.n1433 185
R13768 VDD.n1436 VDD.n1251 185
R13769 VDD.n1439 VDD.n1438 185
R13770 VDD.n1249 VDD.n1248 185
R13771 VDD.n1444 VDD.n1443 185
R13772 VDD.n1446 VDD.n1247 185
R13773 VDD.n1449 VDD.n1448 185
R13774 VDD.n1245 VDD.n1244 185
R13775 VDD.n1456 VDD.n1455 185
R13776 VDD.n1458 VDD.n1243 185
R13777 VDD.n1459 VDD.n1242 185
R13778 VDD.n1462 VDD.n1461 185
R13779 VDD.n1464 VDD.n1238 185
R13780 VDD.n1238 VDD.n1237 185
R13781 VDD.n2118 VDD.n2117 185
R13782 VDD.n2121 VDD.n1100 185
R13783 VDD.n2122 VDD.n1099 185
R13784 VDD.n2123 VDD.n1098 185
R13785 VDD.n1110 VDD.n1096 185
R13786 VDD.n2127 VDD.n1095 185
R13787 VDD.n2128 VDD.n1094 185
R13788 VDD.n2129 VDD.n1093 185
R13789 VDD.n2012 VDD.n1092 185
R13790 VDD.n2015 VDD.n2014 185
R13791 VDD.n2017 VDD.n2016 185
R13792 VDD.n2019 VDD.n2010 185
R13793 VDD.n2021 VDD.n2020 185
R13794 VDD.n2022 VDD.n2006 185
R13795 VDD.n2024 VDD.n2023 185
R13796 VDD.n2026 VDD.n2004 185
R13797 VDD.n2028 VDD.n2027 185
R13798 VDD.n2029 VDD.n2000 185
R13799 VDD.n2031 VDD.n2030 185
R13800 VDD.n2033 VDD.n1997 185
R13801 VDD.n2035 VDD.n2034 185
R13802 VDD.n1998 VDD.n1991 185
R13803 VDD.n2039 VDD.n1995 185
R13804 VDD.n2040 VDD.n1987 185
R13805 VDD.n2042 VDD.n2041 185
R13806 VDD.n2044 VDD.n1985 185
R13807 VDD.n2046 VDD.n2045 185
R13808 VDD.n2047 VDD.n1980 185
R13809 VDD.n2049 VDD.n2048 185
R13810 VDD.n2051 VDD.n1978 185
R13811 VDD.n2053 VDD.n2052 185
R13812 VDD.n2054 VDD.n1973 185
R13813 VDD.n2056 VDD.n2055 185
R13814 VDD.n2058 VDD.n1971 185
R13815 VDD.n2060 VDD.n2059 185
R13816 VDD.n2061 VDD.n1966 185
R13817 VDD.n2063 VDD.n2062 185
R13818 VDD.n2065 VDD.n1964 185
R13819 VDD.n2067 VDD.n2066 185
R13820 VDD.n2068 VDD.n1960 185
R13821 VDD.n2070 VDD.n2069 185
R13822 VDD.n2072 VDD.n1957 185
R13823 VDD.n2074 VDD.n2073 185
R13824 VDD.n1958 VDD.n1951 185
R13825 VDD.n2078 VDD.n1955 185
R13826 VDD.n2079 VDD.n1947 185
R13827 VDD.n2081 VDD.n2080 185
R13828 VDD.n2083 VDD.n1945 185
R13829 VDD.n2085 VDD.n2084 185
R13830 VDD.n2086 VDD.n1941 185
R13831 VDD.n2088 VDD.n2087 185
R13832 VDD.n2090 VDD.n1936 185
R13833 VDD.n2092 VDD.n2091 185
R13834 VDD.n1939 VDD.n1935 185
R13835 VDD.n1938 VDD.n1933 185
R13836 VDD.n2096 VDD.n1930 185
R13837 VDD.n2098 VDD.n2097 185
R13838 VDD.n2100 VDD.n1928 185
R13839 VDD.n2102 VDD.n2101 185
R13840 VDD.n2103 VDD.n1923 185
R13841 VDD.n2105 VDD.n2104 185
R13842 VDD.n2107 VDD.n1921 185
R13843 VDD.n2109 VDD.n2108 185
R13844 VDD.n2110 VDD.n1115 185
R13845 VDD.n2116 VDD.n1107 185
R13846 VDD.n2116 VDD.n2115 185
R13847 VDD.n1123 VDD.n1106 185
R13848 VDD.n1108 VDD.n1106 185
R13849 VDD.n1914 VDD.n1913 185
R13850 VDD.n1915 VDD.n1914 185
R13851 VDD.n1122 VDD.n1121 185
R13852 VDD.n1121 VDD.n1120 185
R13853 VDD.n1908 VDD.n1907 185
R13854 VDD.n1907 VDD.n1906 185
R13855 VDD.n1126 VDD.n1125 185
R13856 VDD.n1127 VDD.n1126 185
R13857 VDD.n1897 VDD.n1896 185
R13858 VDD.n1898 VDD.n1897 185
R13859 VDD.n1134 VDD.n1133 185
R13860 VDD.n1139 VDD.n1133 185
R13861 VDD.n1892 VDD.n1891 185
R13862 VDD.n1891 VDD.n1890 185
R13863 VDD.n1137 VDD.n1136 185
R13864 VDD.n1138 VDD.n1137 185
R13865 VDD.n1881 VDD.n1880 185
R13866 VDD.n1882 VDD.n1881 185
R13867 VDD.n1147 VDD.n1146 185
R13868 VDD.n1146 VDD.n1145 185
R13869 VDD.n1876 VDD.n1875 185
R13870 VDD.n1875 VDD.n1874 185
R13871 VDD.n1150 VDD.n1149 185
R13872 VDD.n1151 VDD.n1150 185
R13873 VDD.n1865 VDD.n1864 185
R13874 VDD.n1866 VDD.n1865 185
R13875 VDD.n1158 VDD.n1157 185
R13876 VDD.n1163 VDD.n1157 185
R13877 VDD.n1860 VDD.n1859 185
R13878 VDD.n1859 VDD.n1858 185
R13879 VDD.n1161 VDD.n1160 185
R13880 VDD.n1162 VDD.n1161 185
R13881 VDD.n1849 VDD.n1848 185
R13882 VDD.n1850 VDD.n1849 185
R13883 VDD.n1171 VDD.n1170 185
R13884 VDD.n1170 VDD.n1169 185
R13885 VDD.n1844 VDD.n1843 185
R13886 VDD.n1843 VDD.n1842 185
R13887 VDD.n1174 VDD.n1173 185
R13888 VDD.n1175 VDD.n1174 185
R13889 VDD.n1551 VDD.n1550 185
R13890 VDD.n1552 VDD.n1551 185
R13891 VDD.n1182 VDD.n1181 185
R13892 VDD.n1186 VDD.n1181 185
R13893 VDD.n1546 VDD.n1545 185
R13894 VDD.n1545 VDD.n1544 185
R13895 VDD.n1185 VDD.n1184 185
R13896 VDD.n1535 VDD.n1185 185
R13897 VDD.n1534 VDD.n1533 185
R13898 VDD.n1536 VDD.n1534 185
R13899 VDD.n1194 VDD.n1193 185
R13900 VDD.n1193 VDD.n1192 185
R13901 VDD.n1529 VDD.n1528 185
R13902 VDD.n1528 VDD.n1527 185
R13903 VDD.n1197 VDD.n1196 185
R13904 VDD.n1198 VDD.n1197 185
R13905 VDD.n1518 VDD.n1517 185
R13906 VDD.n1519 VDD.n1518 185
R13907 VDD.n1205 VDD.n1204 185
R13908 VDD.n1209 VDD.n1204 185
R13909 VDD.n1513 VDD.n1512 185
R13910 VDD.n1512 VDD.n1511 185
R13911 VDD.n1208 VDD.n1207 185
R13912 VDD.n1502 VDD.n1208 185
R13913 VDD.n1501 VDD.n1500 185
R13914 VDD.n1503 VDD.n1501 185
R13915 VDD.n1217 VDD.n1216 185
R13916 VDD.n1216 VDD.n1215 185
R13917 VDD.n1496 VDD.n1495 185
R13918 VDD.n1495 VDD.n1494 185
R13919 VDD.n1220 VDD.n1219 185
R13920 VDD.n1221 VDD.n1220 185
R13921 VDD.n1485 VDD.n1484 185
R13922 VDD.n1486 VDD.n1485 185
R13923 VDD.n1229 VDD.n1228 185
R13924 VDD.n1228 VDD.n1227 185
R13925 VDD.n1480 VDD.n1479 185
R13926 VDD.n1479 VDD.n1478 185
R13927 VDD.n1232 VDD.n1231 185
R13928 VDD.n1469 VDD.n1232 185
R13929 VDD.n1468 VDD.n1467 185
R13930 VDD.n1470 VDD.n1468 185
R13931 VDD.n3214 VDD.n3213 185
R13932 VDD.n3212 VDD.n694 185
R13933 VDD.n3211 VDD.n693 185
R13934 VDD.n3216 VDD.n693 185
R13935 VDD.n3210 VDD.n3209 185
R13936 VDD.n3208 VDD.n3207 185
R13937 VDD.n3206 VDD.n3205 185
R13938 VDD.n3204 VDD.n3203 185
R13939 VDD.n3202 VDD.n3201 185
R13940 VDD.n3200 VDD.n3199 185
R13941 VDD.n3198 VDD.n3197 185
R13942 VDD.n3196 VDD.n3195 185
R13943 VDD.n3194 VDD.n3193 185
R13944 VDD.n3192 VDD.n3191 185
R13945 VDD.n3190 VDD.n3189 185
R13946 VDD.n3188 VDD.n3187 185
R13947 VDD.n3186 VDD.n3185 185
R13948 VDD.n3184 VDD.n3183 185
R13949 VDD.n3182 VDD.n3181 185
R13950 VDD.n3180 VDD.n3179 185
R13951 VDD.n3178 VDD.n3177 185
R13952 VDD.n3169 VDD.n712 185
R13953 VDD.n3171 VDD.n3170 185
R13954 VDD.n3168 VDD.n3167 185
R13955 VDD.n3166 VDD.n3165 185
R13956 VDD.n3164 VDD.n3163 185
R13957 VDD.n3162 VDD.n3161 185
R13958 VDD.n3160 VDD.n3159 185
R13959 VDD.n3158 VDD.n3157 185
R13960 VDD.n3156 VDD.n3155 185
R13961 VDD.n3154 VDD.n3153 185
R13962 VDD.n3152 VDD.n3151 185
R13963 VDD.n3150 VDD.n3149 185
R13964 VDD.n3148 VDD.n3147 185
R13965 VDD.n3146 VDD.n3145 185
R13966 VDD.n3144 VDD.n3143 185
R13967 VDD.n3142 VDD.n3141 185
R13968 VDD.n3140 VDD.n3139 185
R13969 VDD.n3138 VDD.n3137 185
R13970 VDD.n3136 VDD.n3135 185
R13971 VDD.n3134 VDD.n3133 185
R13972 VDD.n3132 VDD.n3131 185
R13973 VDD.n3130 VDD.n3129 185
R13974 VDD.n3123 VDD.n732 185
R13975 VDD.n3125 VDD.n3124 185
R13976 VDD.n3122 VDD.n3121 185
R13977 VDD.n3120 VDD.n3119 185
R13978 VDD.n3118 VDD.n3117 185
R13979 VDD.n3116 VDD.n3115 185
R13980 VDD.n3114 VDD.n3113 185
R13981 VDD.n3112 VDD.n3111 185
R13982 VDD.n3110 VDD.n3109 185
R13983 VDD.n3108 VDD.n3107 185
R13984 VDD.n3106 VDD.n3105 185
R13985 VDD.n3104 VDD.n3103 185
R13986 VDD.n3102 VDD.n3101 185
R13987 VDD.n3100 VDD.n3099 185
R13988 VDD.n3098 VDD.n3097 185
R13989 VDD.n3096 VDD.n3095 185
R13990 VDD.n3094 VDD.n3093 185
R13991 VDD.n3092 VDD.n3091 185
R13992 VDD.n3090 VDD.n3089 185
R13993 VDD.n3088 VDD.n3087 185
R13994 VDD.n3086 VDD.n661 185
R13995 VDD.n3218 VDD.n3217 185
R13996 VDD.n3217 VDD.n3216 185
R13997 VDD.n3345 VDD.n3344 185
R13998 VDD.n586 VDD.n391 185
R13999 VDD.n585 VDD.n584 185
R14000 VDD.n583 VDD.n582 185
R14001 VDD.n581 VDD.n396 185
R14002 VDD.n577 VDD.n576 185
R14003 VDD.n575 VDD.n574 185
R14004 VDD.n573 VDD.n572 185
R14005 VDD.n571 VDD.n398 185
R14006 VDD.n567 VDD.n566 185
R14007 VDD.n565 VDD.n564 185
R14008 VDD.n563 VDD.n562 185
R14009 VDD.n561 VDD.n400 185
R14010 VDD.n557 VDD.n556 185
R14011 VDD.n555 VDD.n554 185
R14012 VDD.n553 VDD.n552 185
R14013 VDD.n551 VDD.n402 185
R14014 VDD.n547 VDD.n546 185
R14015 VDD.n545 VDD.n544 185
R14016 VDD.n543 VDD.n542 185
R14017 VDD.n541 VDD.n404 185
R14018 VDD.n537 VDD.n536 185
R14019 VDD.n535 VDD.n534 185
R14020 VDD.n533 VDD.n532 185
R14021 VDD.n531 VDD.n408 185
R14022 VDD.n527 VDD.n526 185
R14023 VDD.n525 VDD.n524 185
R14024 VDD.n523 VDD.n522 185
R14025 VDD.n521 VDD.n410 185
R14026 VDD.n517 VDD.n516 185
R14027 VDD.n515 VDD.n514 185
R14028 VDD.n513 VDD.n512 185
R14029 VDD.n511 VDD.n412 185
R14030 VDD.n507 VDD.n506 185
R14031 VDD.n505 VDD.n504 185
R14032 VDD.n503 VDD.n502 185
R14033 VDD.n501 VDD.n414 185
R14034 VDD.n497 VDD.n496 185
R14035 VDD.n495 VDD.n494 185
R14036 VDD.n493 VDD.n492 185
R14037 VDD.n491 VDD.n416 185
R14038 VDD.n487 VDD.n486 185
R14039 VDD.n485 VDD.n484 185
R14040 VDD.n483 VDD.n482 185
R14041 VDD.n481 VDD.n420 185
R14042 VDD.n477 VDD.n476 185
R14043 VDD.n475 VDD.n474 185
R14044 VDD.n473 VDD.n472 185
R14045 VDD.n471 VDD.n422 185
R14046 VDD.n467 VDD.n466 185
R14047 VDD.n465 VDD.n464 185
R14048 VDD.n463 VDD.n462 185
R14049 VDD.n461 VDD.n424 185
R14050 VDD.n457 VDD.n456 185
R14051 VDD.n455 VDD.n454 185
R14052 VDD.n453 VDD.n452 185
R14053 VDD.n451 VDD.n426 185
R14054 VDD.n447 VDD.n446 185
R14055 VDD.n445 VDD.n444 185
R14056 VDD.n443 VDD.n442 185
R14057 VDD.n441 VDD.n428 185
R14058 VDD.n437 VDD.n436 185
R14059 VDD.n435 VDD.n434 185
R14060 VDD.n433 VDD.n432 185
R14061 VDD.n3341 VDD.n359 185
R14062 VDD.n3348 VDD.n359 185
R14063 VDD.n3340 VDD.n358 185
R14064 VDD.n3349 VDD.n358 185
R14065 VDD.n3339 VDD.n3338 185
R14066 VDD.n3338 VDD.n350 185
R14067 VDD.n589 VDD.n349 185
R14068 VDD.n3355 VDD.n349 185
R14069 VDD.n3334 VDD.n348 185
R14070 VDD.n3356 VDD.n348 185
R14071 VDD.n3333 VDD.n347 185
R14072 VDD.n3357 VDD.n347 185
R14073 VDD.n3332 VDD.n3331 185
R14074 VDD.n3331 VDD.n346 185
R14075 VDD.n591 VDD.n338 185
R14076 VDD.n3363 VDD.n338 185
R14077 VDD.n3327 VDD.n337 185
R14078 VDD.n3364 VDD.n337 185
R14079 VDD.n3326 VDD.n336 185
R14080 VDD.n3365 VDD.n336 185
R14081 VDD.n3325 VDD.n3324 185
R14082 VDD.n3324 VDD.n328 185
R14083 VDD.n593 VDD.n327 185
R14084 VDD.n3371 VDD.n327 185
R14085 VDD.n3320 VDD.n326 185
R14086 VDD.n3372 VDD.n326 185
R14087 VDD.n3319 VDD.n325 185
R14088 VDD.n3373 VDD.n325 185
R14089 VDD.n3318 VDD.n3317 185
R14090 VDD.n3317 VDD.n324 185
R14091 VDD.n595 VDD.n316 185
R14092 VDD.n3379 VDD.n316 185
R14093 VDD.n3313 VDD.n315 185
R14094 VDD.n3380 VDD.n315 185
R14095 VDD.n3312 VDD.n314 185
R14096 VDD.n3381 VDD.n314 185
R14097 VDD.n3311 VDD.n3310 185
R14098 VDD.n3310 VDD.n307 185
R14099 VDD.n597 VDD.n306 185
R14100 VDD.n3387 VDD.n306 185
R14101 VDD.n3306 VDD.n305 185
R14102 VDD.n3388 VDD.n305 185
R14103 VDD.n3305 VDD.n304 185
R14104 VDD.n3389 VDD.n304 185
R14105 VDD.n3304 VDD.n3303 185
R14106 VDD.n3303 VDD.n303 185
R14107 VDD.n3302 VDD.n599 185
R14108 VDD.n3302 VDD.n3301 185
R14109 VDD.n3290 VDD.n601 185
R14110 VDD.n602 VDD.n601 185
R14111 VDD.n3292 VDD.n3291 185
R14112 VDD.n3293 VDD.n3292 185
R14113 VDD.n610 VDD.n609 185
R14114 VDD.n609 VDD.n608 185
R14115 VDD.n3284 VDD.n3283 185
R14116 VDD.n3283 VDD.n3282 185
R14117 VDD.n613 VDD.n612 185
R14118 VDD.n3273 VDD.n613 185
R14119 VDD.n3272 VDD.n3271 185
R14120 VDD.n3274 VDD.n3272 185
R14121 VDD.n621 VDD.n620 185
R14122 VDD.n620 VDD.n619 185
R14123 VDD.n3267 VDD.n3266 185
R14124 VDD.n3266 VDD.n3265 185
R14125 VDD.n624 VDD.n623 185
R14126 VDD.n625 VDD.n624 185
R14127 VDD.n3256 VDD.n3255 185
R14128 VDD.n3257 VDD.n3256 185
R14129 VDD.n633 VDD.n632 185
R14130 VDD.n632 VDD.n631 185
R14131 VDD.n3251 VDD.n3250 185
R14132 VDD.n3250 VDD.n3249 185
R14133 VDD.n636 VDD.n635 185
R14134 VDD.n3240 VDD.n636 185
R14135 VDD.n3239 VDD.n3238 185
R14136 VDD.n3241 VDD.n3239 185
R14137 VDD.n644 VDD.n643 185
R14138 VDD.n643 VDD.n642 185
R14139 VDD.n3234 VDD.n3233 185
R14140 VDD.n3233 VDD.n3232 185
R14141 VDD.n647 VDD.n646 185
R14142 VDD.n648 VDD.n647 185
R14143 VDD.n3223 VDD.n3222 185
R14144 VDD.n3224 VDD.n3223 185
R14145 VDD.n656 VDD.n655 185
R14146 VDD.n655 VDD.n654 185
R14147 VDD.n653 VDD.n652 185
R14148 VDD.n654 VDD.n653 185
R14149 VDD.n3226 VDD.n3225 185
R14150 VDD.n3225 VDD.n3224 185
R14151 VDD.n650 VDD.n649 185
R14152 VDD.n649 VDD.n648 185
R14153 VDD.n3231 VDD.n3230 185
R14154 VDD.n3232 VDD.n3231 185
R14155 VDD.n641 VDD.n640 185
R14156 VDD.n642 VDD.n641 185
R14157 VDD.n3243 VDD.n3242 185
R14158 VDD.n3242 VDD.n3241 185
R14159 VDD.n638 VDD.n637 185
R14160 VDD.n3240 VDD.n637 185
R14161 VDD.n3248 VDD.n3247 185
R14162 VDD.n3249 VDD.n3248 185
R14163 VDD.n630 VDD.n629 185
R14164 VDD.n631 VDD.n630 185
R14165 VDD.n3259 VDD.n3258 185
R14166 VDD.n3258 VDD.n3257 185
R14167 VDD.n627 VDD.n626 185
R14168 VDD.n626 VDD.n625 185
R14169 VDD.n3264 VDD.n3263 185
R14170 VDD.n3265 VDD.n3264 185
R14171 VDD.n618 VDD.n617 185
R14172 VDD.n619 VDD.n618 185
R14173 VDD.n3276 VDD.n3275 185
R14174 VDD.n3275 VDD.n3274 185
R14175 VDD.n615 VDD.n614 185
R14176 VDD.n3273 VDD.n614 185
R14177 VDD.n3281 VDD.n3280 185
R14178 VDD.n3282 VDD.n3281 185
R14179 VDD.n607 VDD.n606 185
R14180 VDD.n608 VDD.n607 185
R14181 VDD.n3295 VDD.n3294 185
R14182 VDD.n3294 VDD.n3293 185
R14183 VDD.n604 VDD.n603 185
R14184 VDD.n603 VDD.n602 185
R14185 VDD.n3300 VDD.n3299 185
R14186 VDD.n3301 VDD.n3300 185
R14187 VDD.n301 VDD.n299 185
R14188 VDD.n303 VDD.n301 185
R14189 VDD.n3391 VDD.n3390 185
R14190 VDD.n3390 VDD.n3389 185
R14191 VDD.n302 VDD.n300 185
R14192 VDD.n3388 VDD.n302 185
R14193 VDD.n3386 VDD.n3385 185
R14194 VDD.n3387 VDD.n3386 185
R14195 VDD.n3384 VDD.n308 185
R14196 VDD.n308 VDD.n307 185
R14197 VDD.n3383 VDD.n3382 185
R14198 VDD.n3382 VDD.n3381 185
R14199 VDD.n313 VDD.n312 185
R14200 VDD.n3380 VDD.n313 185
R14201 VDD.n3378 VDD.n3377 185
R14202 VDD.n3379 VDD.n3378 185
R14203 VDD.n3376 VDD.n317 185
R14204 VDD.n324 VDD.n317 185
R14205 VDD.n3375 VDD.n3374 185
R14206 VDD.n3374 VDD.n3373 185
R14207 VDD.n323 VDD.n322 185
R14208 VDD.n3372 VDD.n323 185
R14209 VDD.n3370 VDD.n3369 185
R14210 VDD.n3371 VDD.n3370 185
R14211 VDD.n3368 VDD.n329 185
R14212 VDD.n329 VDD.n328 185
R14213 VDD.n3367 VDD.n3366 185
R14214 VDD.n3366 VDD.n3365 185
R14215 VDD.n335 VDD.n334 185
R14216 VDD.n3364 VDD.n335 185
R14217 VDD.n3362 VDD.n3361 185
R14218 VDD.n3363 VDD.n3362 185
R14219 VDD.n3360 VDD.n339 185
R14220 VDD.n346 VDD.n339 185
R14221 VDD.n3359 VDD.n3358 185
R14222 VDD.n3358 VDD.n3357 185
R14223 VDD.n345 VDD.n344 185
R14224 VDD.n3356 VDD.n345 185
R14225 VDD.n3354 VDD.n3353 185
R14226 VDD.n3355 VDD.n3354 185
R14227 VDD.n3352 VDD.n351 185
R14228 VDD.n351 VDD.n350 185
R14229 VDD.n3351 VDD.n3350 185
R14230 VDD.n3350 VDD.n3349 185
R14231 VDD.n357 VDD.n356 185
R14232 VDD.n3348 VDD.n357 185
R14233 VDD.n932 VDD.n930 185
R14234 VDD.n930 VDD.n903 185
R14235 VDD.n2471 VDD.n939 185
R14236 VDD.n2536 VDD.n939 185
R14237 VDD.n2473 VDD.n2472 185
R14238 VDD.n2474 VDD.n2473 185
R14239 VDD.n2470 VDD.n948 185
R14240 VDD.n948 VDD.n947 185
R14241 VDD.n2469 VDD.n2468 185
R14242 VDD.n2468 VDD.n2467 185
R14243 VDD.n950 VDD.n949 185
R14244 VDD.n951 VDD.n950 185
R14245 VDD.n2459 VDD.n2458 185
R14246 VDD.n2460 VDD.n2459 185
R14247 VDD.n2457 VDD.n961 185
R14248 VDD.n961 VDD.n958 185
R14249 VDD.n2456 VDD.n2455 185
R14250 VDD.n2455 VDD.n2454 185
R14251 VDD.n963 VDD.n962 185
R14252 VDD.n964 VDD.n963 185
R14253 VDD.n2447 VDD.n2446 185
R14254 VDD.n2448 VDD.n2447 185
R14255 VDD.n2445 VDD.n972 185
R14256 VDD.n978 VDD.n972 185
R14257 VDD.n2444 VDD.n2443 185
R14258 VDD.n2443 VDD.n2442 185
R14259 VDD.n974 VDD.n973 185
R14260 VDD.n975 VDD.n974 185
R14261 VDD.n2435 VDD.n2434 185
R14262 VDD.n2436 VDD.n2435 185
R14263 VDD.n2433 VDD.n984 185
R14264 VDD.n2261 VDD.n984 185
R14265 VDD.n2432 VDD.n2431 185
R14266 VDD.n2431 VDD.n2430 185
R14267 VDD.n986 VDD.n985 185
R14268 VDD.n987 VDD.n986 185
R14269 VDD.n2423 VDD.n2422 185
R14270 VDD.n2424 VDD.n2423 185
R14271 VDD.n2421 VDD.n995 185
R14272 VDD.n2270 VDD.n995 185
R14273 VDD.n2420 VDD.n2419 185
R14274 VDD.n2419 VDD.n2418 185
R14275 VDD.n997 VDD.n996 185
R14276 VDD.n998 VDD.n997 185
R14277 VDD.n2411 VDD.n2410 185
R14278 VDD.n2412 VDD.n2411 185
R14279 VDD.n2409 VDD.n1007 185
R14280 VDD.n1007 VDD.n1004 185
R14281 VDD.n2408 VDD.n2407 185
R14282 VDD.n2407 VDD.n2406 185
R14283 VDD.n1009 VDD.n1008 185
R14284 VDD.n1010 VDD.n1009 185
R14285 VDD.n2399 VDD.n2398 185
R14286 VDD.n2400 VDD.n2399 185
R14287 VDD.n2397 VDD.n1019 185
R14288 VDD.n1019 VDD.n1016 185
R14289 VDD.n2396 VDD.n2395 185
R14290 VDD.n2395 VDD.n2394 185
R14291 VDD.n1021 VDD.n1020 185
R14292 VDD.n1022 VDD.n1021 185
R14293 VDD.n2387 VDD.n2386 185
R14294 VDD.n2388 VDD.n2387 185
R14295 VDD.n2385 VDD.n1031 185
R14296 VDD.n1031 VDD.n1028 185
R14297 VDD.n2384 VDD.n2383 185
R14298 VDD.n2383 VDD.n2382 185
R14299 VDD.n1033 VDD.n1032 185
R14300 VDD.n1034 VDD.n1033 185
R14301 VDD.n2375 VDD.n2374 185
R14302 VDD.n2376 VDD.n2375 185
R14303 VDD.n2372 VDD.n1042 185
R14304 VDD.n1048 VDD.n1042 185
R14305 VDD.n2371 VDD.n2370 185
R14306 VDD.n2370 VDD.n2369 185
R14307 VDD.n1045 VDD.n1044 185
R14308 VDD.n1055 VDD.n1045 185
R14309 VDD.n2362 VDD.n2361 185
R14310 VDD.n2363 VDD.n2362 185
R14311 VDD.n2360 VDD.n1056 185
R14312 VDD.n1056 VDD.n1052 185
R14313 VDD.n2359 VDD.n2358 185
R14314 VDD.n2358 VDD.n2357 185
R14315 VDD.n2540 VDD.n929 185
R14316 VDD.n2590 VDD.n929 185
R14317 VDD.n2542 VDD.n2541 185
R14318 VDD.n2544 VDD.n2543 185
R14319 VDD.n2546 VDD.n2545 185
R14320 VDD.n2548 VDD.n2547 185
R14321 VDD.n2550 VDD.n2549 185
R14322 VDD.n2552 VDD.n2551 185
R14323 VDD.n2554 VDD.n2553 185
R14324 VDD.n2556 VDD.n2555 185
R14325 VDD.n2558 VDD.n2557 185
R14326 VDD.n2560 VDD.n2559 185
R14327 VDD.n2562 VDD.n2561 185
R14328 VDD.n2564 VDD.n2563 185
R14329 VDD.n2566 VDD.n2565 185
R14330 VDD.n2568 VDD.n2567 185
R14331 VDD.n2570 VDD.n2569 185
R14332 VDD.n2572 VDD.n2571 185
R14333 VDD.n2574 VDD.n2573 185
R14334 VDD.n2576 VDD.n2575 185
R14335 VDD.n2578 VDD.n2577 185
R14336 VDD.n2580 VDD.n2579 185
R14337 VDD.n2582 VDD.n2581 185
R14338 VDD.n2584 VDD.n2583 185
R14339 VDD.n2586 VDD.n2585 185
R14340 VDD.n2587 VDD.n931 185
R14341 VDD.n2589 VDD.n2588 185
R14342 VDD.n2590 VDD.n2589 185
R14343 VDD.n2539 VDD.n2538 185
R14344 VDD.n2538 VDD.n903 185
R14345 VDD.n2537 VDD.n936 185
R14346 VDD.n2537 VDD.n2536 185
R14347 VDD.n2221 VDD.n937 185
R14348 VDD.n2474 VDD.n937 185
R14349 VDD.n2223 VDD.n2222 185
R14350 VDD.n2222 VDD.n947 185
R14351 VDD.n2224 VDD.n953 185
R14352 VDD.n2467 VDD.n953 185
R14353 VDD.n2226 VDD.n2225 185
R14354 VDD.n2225 VDD.n951 185
R14355 VDD.n2227 VDD.n960 185
R14356 VDD.n2460 VDD.n960 185
R14357 VDD.n2229 VDD.n2228 185
R14358 VDD.n2228 VDD.n958 185
R14359 VDD.n2230 VDD.n966 185
R14360 VDD.n2454 VDD.n966 185
R14361 VDD.n2232 VDD.n2231 185
R14362 VDD.n2231 VDD.n964 185
R14363 VDD.n2233 VDD.n971 185
R14364 VDD.n2448 VDD.n971 185
R14365 VDD.n2235 VDD.n2234 185
R14366 VDD.n2234 VDD.n978 185
R14367 VDD.n2236 VDD.n977 185
R14368 VDD.n2442 VDD.n977 185
R14369 VDD.n2238 VDD.n2237 185
R14370 VDD.n2237 VDD.n975 185
R14371 VDD.n2239 VDD.n983 185
R14372 VDD.n2436 VDD.n983 185
R14373 VDD.n2263 VDD.n2262 185
R14374 VDD.n2262 VDD.n2261 185
R14375 VDD.n2264 VDD.n989 185
R14376 VDD.n2430 VDD.n989 185
R14377 VDD.n2266 VDD.n2265 185
R14378 VDD.n2265 VDD.n987 185
R14379 VDD.n2267 VDD.n994 185
R14380 VDD.n2424 VDD.n994 185
R14381 VDD.n2269 VDD.n2268 185
R14382 VDD.n2270 VDD.n2269 185
R14383 VDD.n2220 VDD.n1000 185
R14384 VDD.n2418 VDD.n1000 185
R14385 VDD.n2219 VDD.n2218 185
R14386 VDD.n2218 VDD.n998 185
R14387 VDD.n2217 VDD.n1006 185
R14388 VDD.n2412 VDD.n1006 185
R14389 VDD.n2216 VDD.n2215 185
R14390 VDD.n2215 VDD.n1004 185
R14391 VDD.n2214 VDD.n1012 185
R14392 VDD.n2406 VDD.n1012 185
R14393 VDD.n2213 VDD.n2212 185
R14394 VDD.n2212 VDD.n1010 185
R14395 VDD.n2211 VDD.n1018 185
R14396 VDD.n2400 VDD.n1018 185
R14397 VDD.n2210 VDD.n2209 185
R14398 VDD.n2209 VDD.n1016 185
R14399 VDD.n2208 VDD.n1024 185
R14400 VDD.n2394 VDD.n1024 185
R14401 VDD.n2207 VDD.n2206 185
R14402 VDD.n2206 VDD.n1022 185
R14403 VDD.n2205 VDD.n1030 185
R14404 VDD.n2388 VDD.n1030 185
R14405 VDD.n2204 VDD.n2203 185
R14406 VDD.n2203 VDD.n1028 185
R14407 VDD.n2202 VDD.n1036 185
R14408 VDD.n2382 VDD.n1036 185
R14409 VDD.n2201 VDD.n2200 185
R14410 VDD.n2200 VDD.n1034 185
R14411 VDD.n2199 VDD.n1041 185
R14412 VDD.n2376 VDD.n1041 185
R14413 VDD.n2198 VDD.n2197 185
R14414 VDD.n2197 VDD.n1048 185
R14415 VDD.n2196 VDD.n1047 185
R14416 VDD.n2369 VDD.n1047 185
R14417 VDD.n2195 VDD.n2194 185
R14418 VDD.n2194 VDD.n1055 185
R14419 VDD.n2193 VDD.n1054 185
R14420 VDD.n2363 VDD.n1054 185
R14421 VDD.n2192 VDD.n2191 185
R14422 VDD.n2191 VDD.n1052 185
R14423 VDD.n2190 VDD.n1061 185
R14424 VDD.n2357 VDD.n1061 185
R14425 VDD.n1058 VDD.n1057 185
R14426 VDD.n1059 VDD.n1058 185
R14427 VDD.n2141 VDD.n2140 185
R14428 VDD.n2142 VDD.n2138 185
R14429 VDD.n2144 VDD.n2143 185
R14430 VDD.n2146 VDD.n2137 185
R14431 VDD.n2149 VDD.n2148 185
R14432 VDD.n2150 VDD.n2136 185
R14433 VDD.n2152 VDD.n2151 185
R14434 VDD.n2154 VDD.n2135 185
R14435 VDD.n2157 VDD.n2156 185
R14436 VDD.n2158 VDD.n2134 185
R14437 VDD.n2160 VDD.n2159 185
R14438 VDD.n2162 VDD.n2133 185
R14439 VDD.n2165 VDD.n2164 185
R14440 VDD.n2166 VDD.n1087 185
R14441 VDD.n2168 VDD.n2167 185
R14442 VDD.n2170 VDD.n1086 185
R14443 VDD.n2173 VDD.n2172 185
R14444 VDD.n2174 VDD.n1085 185
R14445 VDD.n2176 VDD.n2175 185
R14446 VDD.n2178 VDD.n1084 185
R14447 VDD.n2181 VDD.n2180 185
R14448 VDD.n2182 VDD.n1081 185
R14449 VDD.n2185 VDD.n2184 185
R14450 VDD.n2187 VDD.n1080 185
R14451 VDD.n2189 VDD.n2188 185
R14452 VDD.n2188 VDD.n1059 185
R14453 VDD.n290 VDD.n289 171.744
R14454 VDD.n289 VDD.n288 171.744
R14455 VDD.n288 VDD.n257 171.744
R14456 VDD.n281 VDD.n257 171.744
R14457 VDD.n281 VDD.n280 171.744
R14458 VDD.n280 VDD.n262 171.744
R14459 VDD.n273 VDD.n262 171.744
R14460 VDD.n273 VDD.n272 171.744
R14461 VDD.n272 VDD.n266 171.744
R14462 VDD.n239 VDD.n238 171.744
R14463 VDD.n238 VDD.n237 171.744
R14464 VDD.n237 VDD.n206 171.744
R14465 VDD.n230 VDD.n206 171.744
R14466 VDD.n230 VDD.n229 171.744
R14467 VDD.n229 VDD.n211 171.744
R14468 VDD.n222 VDD.n211 171.744
R14469 VDD.n222 VDD.n221 171.744
R14470 VDD.n221 VDD.n215 171.744
R14471 VDD.n196 VDD.n195 171.744
R14472 VDD.n195 VDD.n194 171.744
R14473 VDD.n194 VDD.n163 171.744
R14474 VDD.n187 VDD.n163 171.744
R14475 VDD.n187 VDD.n186 171.744
R14476 VDD.n186 VDD.n168 171.744
R14477 VDD.n179 VDD.n168 171.744
R14478 VDD.n179 VDD.n178 171.744
R14479 VDD.n178 VDD.n172 171.744
R14480 VDD.n145 VDD.n144 171.744
R14481 VDD.n144 VDD.n143 171.744
R14482 VDD.n143 VDD.n112 171.744
R14483 VDD.n136 VDD.n112 171.744
R14484 VDD.n136 VDD.n135 171.744
R14485 VDD.n135 VDD.n117 171.744
R14486 VDD.n128 VDD.n117 171.744
R14487 VDD.n128 VDD.n127 171.744
R14488 VDD.n127 VDD.n121 171.744
R14489 VDD.n103 VDD.n102 171.744
R14490 VDD.n102 VDD.n101 171.744
R14491 VDD.n101 VDD.n70 171.744
R14492 VDD.n94 VDD.n70 171.744
R14493 VDD.n94 VDD.n93 171.744
R14494 VDD.n93 VDD.n75 171.744
R14495 VDD.n86 VDD.n75 171.744
R14496 VDD.n86 VDD.n85 171.744
R14497 VDD.n85 VDD.n79 171.744
R14498 VDD.n52 VDD.n51 171.744
R14499 VDD.n51 VDD.n50 171.744
R14500 VDD.n50 VDD.n19 171.744
R14501 VDD.n43 VDD.n19 171.744
R14502 VDD.n43 VDD.n42 171.744
R14503 VDD.n42 VDD.n24 171.744
R14504 VDD.n35 VDD.n24 171.744
R14505 VDD.n35 VDD.n34 171.744
R14506 VDD.n34 VDD.n28 171.744
R14507 VDD.n1779 VDD.n1778 171.744
R14508 VDD.n1778 VDD.n1777 171.744
R14509 VDD.n1777 VDD.n1746 171.744
R14510 VDD.n1770 VDD.n1746 171.744
R14511 VDD.n1770 VDD.n1769 171.744
R14512 VDD.n1769 VDD.n1751 171.744
R14513 VDD.n1762 VDD.n1751 171.744
R14514 VDD.n1762 VDD.n1761 171.744
R14515 VDD.n1761 VDD.n1755 171.744
R14516 VDD.n1830 VDD.n1829 171.744
R14517 VDD.n1829 VDD.n1828 171.744
R14518 VDD.n1828 VDD.n1797 171.744
R14519 VDD.n1821 VDD.n1797 171.744
R14520 VDD.n1821 VDD.n1820 171.744
R14521 VDD.n1820 VDD.n1802 171.744
R14522 VDD.n1813 VDD.n1802 171.744
R14523 VDD.n1813 VDD.n1812 171.744
R14524 VDD.n1812 VDD.n1806 171.744
R14525 VDD.n1685 VDD.n1684 171.744
R14526 VDD.n1684 VDD.n1683 171.744
R14527 VDD.n1683 VDD.n1652 171.744
R14528 VDD.n1676 VDD.n1652 171.744
R14529 VDD.n1676 VDD.n1675 171.744
R14530 VDD.n1675 VDD.n1657 171.744
R14531 VDD.n1668 VDD.n1657 171.744
R14532 VDD.n1668 VDD.n1667 171.744
R14533 VDD.n1667 VDD.n1661 171.744
R14534 VDD.n1736 VDD.n1735 171.744
R14535 VDD.n1735 VDD.n1734 171.744
R14536 VDD.n1734 VDD.n1703 171.744
R14537 VDD.n1727 VDD.n1703 171.744
R14538 VDD.n1727 VDD.n1726 171.744
R14539 VDD.n1726 VDD.n1708 171.744
R14540 VDD.n1719 VDD.n1708 171.744
R14541 VDD.n1719 VDD.n1718 171.744
R14542 VDD.n1718 VDD.n1712 171.744
R14543 VDD.n1592 VDD.n1591 171.744
R14544 VDD.n1591 VDD.n1590 171.744
R14545 VDD.n1590 VDD.n1559 171.744
R14546 VDD.n1583 VDD.n1559 171.744
R14547 VDD.n1583 VDD.n1582 171.744
R14548 VDD.n1582 VDD.n1564 171.744
R14549 VDD.n1575 VDD.n1564 171.744
R14550 VDD.n1575 VDD.n1574 171.744
R14551 VDD.n1574 VDD.n1568 171.744
R14552 VDD.n1643 VDD.n1642 171.744
R14553 VDD.n1642 VDD.n1641 171.744
R14554 VDD.n1641 VDD.n1610 171.744
R14555 VDD.n1634 VDD.n1610 171.744
R14556 VDD.n1634 VDD.n1633 171.744
R14557 VDD.n1633 VDD.n1615 171.744
R14558 VDD.n1626 VDD.n1615 171.744
R14559 VDD.n1626 VDD.n1625 171.744
R14560 VDD.n1625 VDD.n1619 171.744
R14561 VDD.n3225 VDD.n653 146.341
R14562 VDD.n3225 VDD.n649 146.341
R14563 VDD.n3231 VDD.n649 146.341
R14564 VDD.n3231 VDD.n641 146.341
R14565 VDD.n3242 VDD.n641 146.341
R14566 VDD.n3242 VDD.n637 146.341
R14567 VDD.n3248 VDD.n637 146.341
R14568 VDD.n3248 VDD.n630 146.341
R14569 VDD.n3258 VDD.n630 146.341
R14570 VDD.n3258 VDD.n626 146.341
R14571 VDD.n3264 VDD.n626 146.341
R14572 VDD.n3264 VDD.n618 146.341
R14573 VDD.n3275 VDD.n618 146.341
R14574 VDD.n3275 VDD.n614 146.341
R14575 VDD.n3281 VDD.n614 146.341
R14576 VDD.n3281 VDD.n607 146.341
R14577 VDD.n3294 VDD.n607 146.341
R14578 VDD.n3294 VDD.n603 146.341
R14579 VDD.n3300 VDD.n603 146.341
R14580 VDD.n3300 VDD.n301 146.341
R14581 VDD.n3390 VDD.n301 146.341
R14582 VDD.n3390 VDD.n302 146.341
R14583 VDD.n3386 VDD.n302 146.341
R14584 VDD.n3386 VDD.n308 146.341
R14585 VDD.n3382 VDD.n308 146.341
R14586 VDD.n3382 VDD.n313 146.341
R14587 VDD.n3378 VDD.n313 146.341
R14588 VDD.n3378 VDD.n317 146.341
R14589 VDD.n3374 VDD.n317 146.341
R14590 VDD.n3374 VDD.n323 146.341
R14591 VDD.n3370 VDD.n323 146.341
R14592 VDD.n3370 VDD.n329 146.341
R14593 VDD.n3366 VDD.n329 146.341
R14594 VDD.n3366 VDD.n335 146.341
R14595 VDD.n3362 VDD.n335 146.341
R14596 VDD.n3362 VDD.n339 146.341
R14597 VDD.n3358 VDD.n339 146.341
R14598 VDD.n3358 VDD.n345 146.341
R14599 VDD.n3354 VDD.n345 146.341
R14600 VDD.n3354 VDD.n351 146.341
R14601 VDD.n3350 VDD.n351 146.341
R14602 VDD.n3350 VDD.n357 146.341
R14603 VDD.n436 VDD.n435 146.341
R14604 VDD.n442 VDD.n441 146.341
R14605 VDD.n446 VDD.n445 146.341
R14606 VDD.n452 VDD.n451 146.341
R14607 VDD.n456 VDD.n455 146.341
R14608 VDD.n462 VDD.n461 146.341
R14609 VDD.n466 VDD.n465 146.341
R14610 VDD.n472 VDD.n471 146.341
R14611 VDD.n476 VDD.n475 146.341
R14612 VDD.n482 VDD.n481 146.341
R14613 VDD.n486 VDD.n485 146.341
R14614 VDD.n492 VDD.n491 146.341
R14615 VDD.n496 VDD.n495 146.341
R14616 VDD.n502 VDD.n501 146.341
R14617 VDD.n506 VDD.n505 146.341
R14618 VDD.n512 VDD.n511 146.341
R14619 VDD.n516 VDD.n515 146.341
R14620 VDD.n522 VDD.n521 146.341
R14621 VDD.n526 VDD.n525 146.341
R14622 VDD.n532 VDD.n531 146.341
R14623 VDD.n536 VDD.n535 146.341
R14624 VDD.n542 VDD.n541 146.341
R14625 VDD.n546 VDD.n545 146.341
R14626 VDD.n552 VDD.n551 146.341
R14627 VDD.n556 VDD.n555 146.341
R14628 VDD.n562 VDD.n561 146.341
R14629 VDD.n566 VDD.n565 146.341
R14630 VDD.n572 VDD.n571 146.341
R14631 VDD.n576 VDD.n575 146.341
R14632 VDD.n582 VDD.n581 146.341
R14633 VDD.n584 VDD.n391 146.341
R14634 VDD.n3223 VDD.n655 146.341
R14635 VDD.n3223 VDD.n647 146.341
R14636 VDD.n3233 VDD.n647 146.341
R14637 VDD.n3233 VDD.n643 146.341
R14638 VDD.n3239 VDD.n643 146.341
R14639 VDD.n3239 VDD.n636 146.341
R14640 VDD.n3250 VDD.n636 146.341
R14641 VDD.n3250 VDD.n632 146.341
R14642 VDD.n3256 VDD.n632 146.341
R14643 VDD.n3256 VDD.n624 146.341
R14644 VDD.n3266 VDD.n624 146.341
R14645 VDD.n3266 VDD.n620 146.341
R14646 VDD.n3272 VDD.n620 146.341
R14647 VDD.n3272 VDD.n613 146.341
R14648 VDD.n3283 VDD.n613 146.341
R14649 VDD.n3283 VDD.n609 146.341
R14650 VDD.n3292 VDD.n609 146.341
R14651 VDD.n3292 VDD.n601 146.341
R14652 VDD.n3302 VDD.n601 146.341
R14653 VDD.n3303 VDD.n3302 146.341
R14654 VDD.n3303 VDD.n304 146.341
R14655 VDD.n305 VDD.n304 146.341
R14656 VDD.n306 VDD.n305 146.341
R14657 VDD.n3310 VDD.n306 146.341
R14658 VDD.n3310 VDD.n314 146.341
R14659 VDD.n315 VDD.n314 146.341
R14660 VDD.n316 VDD.n315 146.341
R14661 VDD.n3317 VDD.n316 146.341
R14662 VDD.n3317 VDD.n325 146.341
R14663 VDD.n326 VDD.n325 146.341
R14664 VDD.n327 VDD.n326 146.341
R14665 VDD.n3324 VDD.n327 146.341
R14666 VDD.n3324 VDD.n336 146.341
R14667 VDD.n337 VDD.n336 146.341
R14668 VDD.n338 VDD.n337 146.341
R14669 VDD.n3331 VDD.n338 146.341
R14670 VDD.n3331 VDD.n347 146.341
R14671 VDD.n348 VDD.n347 146.341
R14672 VDD.n349 VDD.n348 146.341
R14673 VDD.n3338 VDD.n349 146.341
R14674 VDD.n3338 VDD.n358 146.341
R14675 VDD.n359 VDD.n358 146.341
R14676 VDD.n694 VDD.n693 146.341
R14677 VDD.n3209 VDD.n693 146.341
R14678 VDD.n3207 VDD.n3206 146.341
R14679 VDD.n3203 VDD.n3202 146.341
R14680 VDD.n3199 VDD.n3198 146.341
R14681 VDD.n3195 VDD.n3194 146.341
R14682 VDD.n3191 VDD.n3190 146.341
R14683 VDD.n3187 VDD.n3186 146.341
R14684 VDD.n3183 VDD.n3182 146.341
R14685 VDD.n3179 VDD.n3178 146.341
R14686 VDD.n3170 VDD.n3169 146.341
R14687 VDD.n3167 VDD.n3166 146.341
R14688 VDD.n3163 VDD.n3162 146.341
R14689 VDD.n3159 VDD.n3158 146.341
R14690 VDD.n3155 VDD.n3154 146.341
R14691 VDD.n3151 VDD.n3150 146.341
R14692 VDD.n3147 VDD.n3146 146.341
R14693 VDD.n3143 VDD.n3142 146.341
R14694 VDD.n3139 VDD.n3138 146.341
R14695 VDD.n3135 VDD.n3134 146.341
R14696 VDD.n3131 VDD.n3130 146.341
R14697 VDD.n3124 VDD.n3123 146.341
R14698 VDD.n3121 VDD.n3120 146.341
R14699 VDD.n3117 VDD.n3116 146.341
R14700 VDD.n3113 VDD.n3112 146.341
R14701 VDD.n3109 VDD.n3108 146.341
R14702 VDD.n3105 VDD.n3104 146.341
R14703 VDD.n3101 VDD.n3100 146.341
R14704 VDD.n3097 VDD.n3096 146.341
R14705 VDD.n3093 VDD.n3092 146.341
R14706 VDD.n3089 VDD.n3088 146.341
R14707 VDD.n3217 VDD.n661 146.341
R14708 VDD.n2108 VDD.n2107 146.341
R14709 VDD.n2105 VDD.n1923 146.341
R14710 VDD.n2101 VDD.n2100 146.341
R14711 VDD.n2098 VDD.n1930 146.341
R14712 VDD.n1939 VDD.n1938 146.341
R14713 VDD.n2091 VDD.n2090 146.341
R14714 VDD.n2088 VDD.n1941 146.341
R14715 VDD.n2084 VDD.n2083 146.341
R14716 VDD.n2081 VDD.n1947 146.341
R14717 VDD.n1958 VDD.n1955 146.341
R14718 VDD.n2073 VDD.n2072 146.341
R14719 VDD.n2070 VDD.n1960 146.341
R14720 VDD.n2066 VDD.n2065 146.341
R14721 VDD.n2063 VDD.n1966 146.341
R14722 VDD.n2059 VDD.n2058 146.341
R14723 VDD.n2056 VDD.n1973 146.341
R14724 VDD.n2052 VDD.n2051 146.341
R14725 VDD.n2049 VDD.n1980 146.341
R14726 VDD.n2045 VDD.n2044 146.341
R14727 VDD.n2042 VDD.n1987 146.341
R14728 VDD.n1998 VDD.n1995 146.341
R14729 VDD.n2034 VDD.n2033 146.341
R14730 VDD.n2031 VDD.n2000 146.341
R14731 VDD.n2027 VDD.n2026 146.341
R14732 VDD.n2024 VDD.n2006 146.341
R14733 VDD.n2020 VDD.n2019 146.341
R14734 VDD.n2017 VDD.n2014 146.341
R14735 VDD.n2012 VDD.n1093 146.341
R14736 VDD.n1095 VDD.n1094 146.341
R14737 VDD.n1110 VDD.n1098 146.341
R14738 VDD.n1100 VDD.n1099 146.341
R14739 VDD.n1468 VDD.n1232 146.341
R14740 VDD.n1479 VDD.n1232 146.341
R14741 VDD.n1479 VDD.n1228 146.341
R14742 VDD.n1485 VDD.n1228 146.341
R14743 VDD.n1485 VDD.n1220 146.341
R14744 VDD.n1495 VDD.n1220 146.341
R14745 VDD.n1495 VDD.n1216 146.341
R14746 VDD.n1501 VDD.n1216 146.341
R14747 VDD.n1501 VDD.n1208 146.341
R14748 VDD.n1512 VDD.n1208 146.341
R14749 VDD.n1512 VDD.n1204 146.341
R14750 VDD.n1518 VDD.n1204 146.341
R14751 VDD.n1518 VDD.n1197 146.341
R14752 VDD.n1528 VDD.n1197 146.341
R14753 VDD.n1528 VDD.n1193 146.341
R14754 VDD.n1534 VDD.n1193 146.341
R14755 VDD.n1534 VDD.n1185 146.341
R14756 VDD.n1545 VDD.n1185 146.341
R14757 VDD.n1545 VDD.n1181 146.341
R14758 VDD.n1551 VDD.n1181 146.341
R14759 VDD.n1551 VDD.n1174 146.341
R14760 VDD.n1843 VDD.n1174 146.341
R14761 VDD.n1843 VDD.n1170 146.341
R14762 VDD.n1849 VDD.n1170 146.341
R14763 VDD.n1849 VDD.n1161 146.341
R14764 VDD.n1859 VDD.n1161 146.341
R14765 VDD.n1859 VDD.n1157 146.341
R14766 VDD.n1865 VDD.n1157 146.341
R14767 VDD.n1865 VDD.n1150 146.341
R14768 VDD.n1875 VDD.n1150 146.341
R14769 VDD.n1875 VDD.n1146 146.341
R14770 VDD.n1881 VDD.n1146 146.341
R14771 VDD.n1881 VDD.n1137 146.341
R14772 VDD.n1891 VDD.n1137 146.341
R14773 VDD.n1891 VDD.n1133 146.341
R14774 VDD.n1897 VDD.n1133 146.341
R14775 VDD.n1897 VDD.n1126 146.341
R14776 VDD.n1907 VDD.n1126 146.341
R14777 VDD.n1907 VDD.n1121 146.341
R14778 VDD.n1914 VDD.n1121 146.341
R14779 VDD.n1914 VDD.n1106 146.341
R14780 VDD.n2116 VDD.n1106 146.341
R14781 VDD.n1310 VDD.n1306 146.341
R14782 VDD.n1316 VDD.n1306 146.341
R14783 VDD.n1320 VDD.n1318 146.341
R14784 VDD.n1326 VDD.n1302 146.341
R14785 VDD.n1330 VDD.n1328 146.341
R14786 VDD.n1336 VDD.n1298 146.341
R14787 VDD.n1340 VDD.n1338 146.341
R14788 VDD.n1348 VDD.n1294 146.341
R14789 VDD.n1351 VDD.n1350 146.341
R14790 VDD.n1353 VDD.n1289 146.341
R14791 VDD.n1360 VDD.n1285 146.341
R14792 VDD.n1364 VDD.n1362 146.341
R14793 VDD.n1370 VDD.n1281 146.341
R14794 VDD.n1374 VDD.n1372 146.341
R14795 VDD.n1380 VDD.n1277 146.341
R14796 VDD.n1384 VDD.n1382 146.341
R14797 VDD.n1390 VDD.n1273 146.341
R14798 VDD.n1394 VDD.n1392 146.341
R14799 VDD.n1402 VDD.n1269 146.341
R14800 VDD.n1405 VDD.n1404 146.341
R14801 VDD.n1407 VDD.n1264 146.341
R14802 VDD.n1414 VDD.n1260 146.341
R14803 VDD.n1418 VDD.n1416 146.341
R14804 VDD.n1424 VDD.n1256 146.341
R14805 VDD.n1428 VDD.n1426 146.341
R14806 VDD.n1434 VDD.n1252 146.341
R14807 VDD.n1438 VDD.n1436 146.341
R14808 VDD.n1444 VDD.n1248 146.341
R14809 VDD.n1448 VDD.n1446 146.341
R14810 VDD.n1456 VDD.n1244 146.341
R14811 VDD.n1459 VDD.n1458 146.341
R14812 VDD.n1461 VDD.n1238 146.341
R14813 VDD.n1471 VDD.n1233 146.341
R14814 VDD.n1477 VDD.n1233 146.341
R14815 VDD.n1477 VDD.n1226 146.341
R14816 VDD.n1487 VDD.n1226 146.341
R14817 VDD.n1487 VDD.n1222 146.341
R14818 VDD.n1493 VDD.n1222 146.341
R14819 VDD.n1493 VDD.n1214 146.341
R14820 VDD.n1504 VDD.n1214 146.341
R14821 VDD.n1504 VDD.n1210 146.341
R14822 VDD.n1510 VDD.n1210 146.341
R14823 VDD.n1510 VDD.n1203 146.341
R14824 VDD.n1520 VDD.n1203 146.341
R14825 VDD.n1520 VDD.n1199 146.341
R14826 VDD.n1526 VDD.n1199 146.341
R14827 VDD.n1526 VDD.n1191 146.341
R14828 VDD.n1537 VDD.n1191 146.341
R14829 VDD.n1537 VDD.n1187 146.341
R14830 VDD.n1543 VDD.n1187 146.341
R14831 VDD.n1543 VDD.n1180 146.341
R14832 VDD.n1553 VDD.n1180 146.341
R14833 VDD.n1553 VDD.n1176 146.341
R14834 VDD.n1841 VDD.n1176 146.341
R14835 VDD.n1841 VDD.n1168 146.341
R14836 VDD.n1851 VDD.n1168 146.341
R14837 VDD.n1851 VDD.n1164 146.341
R14838 VDD.n1857 VDD.n1164 146.341
R14839 VDD.n1857 VDD.n1156 146.341
R14840 VDD.n1867 VDD.n1156 146.341
R14841 VDD.n1867 VDD.n1152 146.341
R14842 VDD.n1873 VDD.n1152 146.341
R14843 VDD.n1873 VDD.n1144 146.341
R14844 VDD.n1883 VDD.n1144 146.341
R14845 VDD.n1883 VDD.n1140 146.341
R14846 VDD.n1889 VDD.n1140 146.341
R14847 VDD.n1889 VDD.n1132 146.341
R14848 VDD.n1899 VDD.n1132 146.341
R14849 VDD.n1899 VDD.n1128 146.341
R14850 VDD.n1905 VDD.n1128 146.341
R14851 VDD.n1905 VDD.n1119 146.341
R14852 VDD.n1916 VDD.n1119 146.341
R14853 VDD.n1916 VDD.n1114 146.341
R14854 VDD.n2114 VDD.n1114 146.341
R14855 VDD.n1113 VDD.n1059 143.238
R14856 VDD.n3216 VDD.n662 143.238
R14857 VDD.n9 VDD.n7 109.74
R14858 VDD.n2 VDD.n0 109.74
R14859 VDD.n9 VDD.n8 109.166
R14860 VDD.n11 VDD.n10 109.166
R14861 VDD.n13 VDD.n12 109.166
R14862 VDD.n6 VDD.n5 109.166
R14863 VDD.n4 VDD.n3 109.166
R14864 VDD.n2 VDD.n1 109.166
R14865 VDD.n3048 VDD.n3047 99.5127
R14866 VDD.n3045 VDD.n769 99.5127
R14867 VDD.n3041 VDD.n3040 99.5127
R14868 VDD.n3038 VDD.n772 99.5127
R14869 VDD.n3034 VDD.n3033 99.5127
R14870 VDD.n3031 VDD.n775 99.5127
R14871 VDD.n3025 VDD.n3024 99.5127
R14872 VDD.n3022 VDD.n778 99.5127
R14873 VDD.n3018 VDD.n3017 99.5127
R14874 VDD.n3015 VDD.n781 99.5127
R14875 VDD.n3011 VDD.n3010 99.5127
R14876 VDD.n3008 VDD.n784 99.5127
R14877 VDD.n2678 VDD.n2592 99.5127
R14878 VDD.n2678 VDD.n897 99.5127
R14879 VDD.n2681 VDD.n897 99.5127
R14880 VDD.n2681 VDD.n891 99.5127
R14881 VDD.n2684 VDD.n891 99.5127
R14882 VDD.n2684 VDD.n886 99.5127
R14883 VDD.n2687 VDD.n886 99.5127
R14884 VDD.n2687 VDD.n880 99.5127
R14885 VDD.n2690 VDD.n880 99.5127
R14886 VDD.n2690 VDD.n874 99.5127
R14887 VDD.n2693 VDD.n874 99.5127
R14888 VDD.n2693 VDD.n869 99.5127
R14889 VDD.n2696 VDD.n869 99.5127
R14890 VDD.n2696 VDD.n863 99.5127
R14891 VDD.n2767 VDD.n863 99.5127
R14892 VDD.n2767 VDD.n857 99.5127
R14893 VDD.n2763 VDD.n857 99.5127
R14894 VDD.n2763 VDD.n852 99.5127
R14895 VDD.n2760 VDD.n852 99.5127
R14896 VDD.n2760 VDD.n845 99.5127
R14897 VDD.n2722 VDD.n845 99.5127
R14898 VDD.n2722 VDD.n839 99.5127
R14899 VDD.n2719 VDD.n839 99.5127
R14900 VDD.n2719 VDD.n833 99.5127
R14901 VDD.n2716 VDD.n833 99.5127
R14902 VDD.n2716 VDD.n827 99.5127
R14903 VDD.n2713 VDD.n827 99.5127
R14904 VDD.n2713 VDD.n821 99.5127
R14905 VDD.n2710 VDD.n821 99.5127
R14906 VDD.n2710 VDD.n816 99.5127
R14907 VDD.n2707 VDD.n816 99.5127
R14908 VDD.n2707 VDD.n811 99.5127
R14909 VDD.n2704 VDD.n811 99.5127
R14910 VDD.n2704 VDD.n805 99.5127
R14911 VDD.n2701 VDD.n805 99.5127
R14912 VDD.n2701 VDD.n797 99.5127
R14913 VDD.n797 VDD.n789 99.5127
R14914 VDD.n2999 VDD.n789 99.5127
R14915 VDD.n3000 VDD.n2999 99.5127
R14916 VDD.n3000 VDD.n762 99.5127
R14917 VDD.n2627 VDD.n2625 99.5127
R14918 VDD.n2631 VDD.n2625 99.5127
R14919 VDD.n2635 VDD.n2633 99.5127
R14920 VDD.n2639 VDD.n2623 99.5127
R14921 VDD.n2643 VDD.n2641 99.5127
R14922 VDD.n2647 VDD.n2621 99.5127
R14923 VDD.n2651 VDD.n2649 99.5127
R14924 VDD.n2655 VDD.n2619 99.5127
R14925 VDD.n2659 VDD.n2657 99.5127
R14926 VDD.n2663 VDD.n2617 99.5127
R14927 VDD.n2667 VDD.n2665 99.5127
R14928 VDD.n2672 VDD.n2613 99.5127
R14929 VDD.n2675 VDD.n2674 99.5127
R14930 VDD.n2848 VDD.n900 99.5127
R14931 VDD.n2852 VDD.n900 99.5127
R14932 VDD.n2852 VDD.n890 99.5127
R14933 VDD.n2860 VDD.n890 99.5127
R14934 VDD.n2860 VDD.n888 99.5127
R14935 VDD.n2864 VDD.n888 99.5127
R14936 VDD.n2864 VDD.n878 99.5127
R14937 VDD.n2872 VDD.n878 99.5127
R14938 VDD.n2872 VDD.n876 99.5127
R14939 VDD.n2876 VDD.n876 99.5127
R14940 VDD.n2876 VDD.n867 99.5127
R14941 VDD.n2884 VDD.n867 99.5127
R14942 VDD.n2884 VDD.n865 99.5127
R14943 VDD.n2888 VDD.n865 99.5127
R14944 VDD.n2888 VDD.n856 99.5127
R14945 VDD.n2896 VDD.n856 99.5127
R14946 VDD.n2896 VDD.n854 99.5127
R14947 VDD.n2900 VDD.n854 99.5127
R14948 VDD.n2900 VDD.n844 99.5127
R14949 VDD.n2908 VDD.n844 99.5127
R14950 VDD.n2908 VDD.n842 99.5127
R14951 VDD.n2912 VDD.n842 99.5127
R14952 VDD.n2912 VDD.n832 99.5127
R14953 VDD.n2920 VDD.n832 99.5127
R14954 VDD.n2920 VDD.n830 99.5127
R14955 VDD.n2924 VDD.n830 99.5127
R14956 VDD.n2924 VDD.n820 99.5127
R14957 VDD.n2932 VDD.n820 99.5127
R14958 VDD.n2932 VDD.n818 99.5127
R14959 VDD.n2936 VDD.n818 99.5127
R14960 VDD.n2936 VDD.n809 99.5127
R14961 VDD.n2944 VDD.n809 99.5127
R14962 VDD.n2944 VDD.n807 99.5127
R14963 VDD.n2948 VDD.n807 99.5127
R14964 VDD.n2948 VDD.n795 99.5127
R14965 VDD.n2993 VDD.n795 99.5127
R14966 VDD.n2993 VDD.n793 99.5127
R14967 VDD.n2997 VDD.n793 99.5127
R14968 VDD.n2997 VDD.n764 99.5127
R14969 VDD.n3052 VDD.n764 99.5127
R14970 VDD.n2529 VDD.n2528 99.5127
R14971 VDD.n2525 VDD.n2524 99.5127
R14972 VDD.n2521 VDD.n2520 99.5127
R14973 VDD.n2517 VDD.n2516 99.5127
R14974 VDD.n2513 VDD.n2512 99.5127
R14975 VDD.n2509 VDD.n2508 99.5127
R14976 VDD.n2505 VDD.n2504 99.5127
R14977 VDD.n2501 VDD.n2500 99.5127
R14978 VDD.n2497 VDD.n2496 99.5127
R14979 VDD.n2493 VDD.n2492 99.5127
R14980 VDD.n2489 VDD.n2488 99.5127
R14981 VDD.n2484 VDD.n2483 99.5127
R14982 VDD.n2301 VDD.n1060 99.5127
R14983 VDD.n2301 VDD.n1053 99.5127
R14984 VDD.n2298 VDD.n1053 99.5127
R14985 VDD.n2298 VDD.n1046 99.5127
R14986 VDD.n2295 VDD.n1046 99.5127
R14987 VDD.n2295 VDD.n1040 99.5127
R14988 VDD.n2292 VDD.n1040 99.5127
R14989 VDD.n2292 VDD.n1035 99.5127
R14990 VDD.n2289 VDD.n1035 99.5127
R14991 VDD.n2289 VDD.n1029 99.5127
R14992 VDD.n2286 VDD.n1029 99.5127
R14993 VDD.n2286 VDD.n1023 99.5127
R14994 VDD.n2283 VDD.n1023 99.5127
R14995 VDD.n2283 VDD.n1017 99.5127
R14996 VDD.n2280 VDD.n1017 99.5127
R14997 VDD.n2280 VDD.n1011 99.5127
R14998 VDD.n2277 VDD.n1011 99.5127
R14999 VDD.n2277 VDD.n1005 99.5127
R15000 VDD.n2274 VDD.n1005 99.5127
R15001 VDD.n2274 VDD.n999 99.5127
R15002 VDD.n2271 VDD.n999 99.5127
R15003 VDD.n2271 VDD.n993 99.5127
R15004 VDD.n2240 VDD.n993 99.5127
R15005 VDD.n2240 VDD.n988 99.5127
R15006 VDD.n2260 VDD.n988 99.5127
R15007 VDD.n2260 VDD.n982 99.5127
R15008 VDD.n2256 VDD.n982 99.5127
R15009 VDD.n2256 VDD.n976 99.5127
R15010 VDD.n2253 VDD.n976 99.5127
R15011 VDD.n2253 VDD.n970 99.5127
R15012 VDD.n2250 VDD.n970 99.5127
R15013 VDD.n2250 VDD.n965 99.5127
R15014 VDD.n2247 VDD.n965 99.5127
R15015 VDD.n2247 VDD.n959 99.5127
R15016 VDD.n2244 VDD.n959 99.5127
R15017 VDD.n2244 VDD.n952 99.5127
R15018 VDD.n952 VDD.n946 99.5127
R15019 VDD.n2475 VDD.n946 99.5127
R15020 VDD.n2475 VDD.n938 99.5127
R15021 VDD.n2479 VDD.n938 99.5127
R15022 VDD.n2352 VDD.n2350 99.5127
R15023 VDD.n2350 VDD.n2349 99.5127
R15024 VDD.n2346 VDD.n2345 99.5127
R15025 VDD.n2343 VDD.n1066 99.5127
R15026 VDD.n2339 VDD.n2337 99.5127
R15027 VDD.n2335 VDD.n1068 99.5127
R15028 VDD.n2331 VDD.n2329 99.5127
R15029 VDD.n2326 VDD.n2325 99.5127
R15030 VDD.n2323 VDD.n1072 99.5127
R15031 VDD.n2319 VDD.n2317 99.5127
R15032 VDD.n2315 VDD.n1074 99.5127
R15033 VDD.n2311 VDD.n2309 99.5127
R15034 VDD.n2306 VDD.n2305 99.5127
R15035 VDD.n2356 VDD.n1051 99.5127
R15036 VDD.n2364 VDD.n1051 99.5127
R15037 VDD.n2364 VDD.n1049 99.5127
R15038 VDD.n2368 VDD.n1049 99.5127
R15039 VDD.n2368 VDD.n1039 99.5127
R15040 VDD.n2377 VDD.n1039 99.5127
R15041 VDD.n2377 VDD.n1037 99.5127
R15042 VDD.n2381 VDD.n1037 99.5127
R15043 VDD.n2381 VDD.n1027 99.5127
R15044 VDD.n2389 VDD.n1027 99.5127
R15045 VDD.n2389 VDD.n1025 99.5127
R15046 VDD.n2393 VDD.n1025 99.5127
R15047 VDD.n2393 VDD.n1015 99.5127
R15048 VDD.n2401 VDD.n1015 99.5127
R15049 VDD.n2401 VDD.n1013 99.5127
R15050 VDD.n2405 VDD.n1013 99.5127
R15051 VDD.n2405 VDD.n1003 99.5127
R15052 VDD.n2413 VDD.n1003 99.5127
R15053 VDD.n2413 VDD.n1001 99.5127
R15054 VDD.n2417 VDD.n1001 99.5127
R15055 VDD.n2417 VDD.n992 99.5127
R15056 VDD.n2425 VDD.n992 99.5127
R15057 VDD.n2425 VDD.n990 99.5127
R15058 VDD.n2429 VDD.n990 99.5127
R15059 VDD.n2429 VDD.n981 99.5127
R15060 VDD.n2437 VDD.n981 99.5127
R15061 VDD.n2437 VDD.n979 99.5127
R15062 VDD.n2441 VDD.n979 99.5127
R15063 VDD.n2441 VDD.n969 99.5127
R15064 VDD.n2449 VDD.n969 99.5127
R15065 VDD.n2449 VDD.n967 99.5127
R15066 VDD.n2453 VDD.n967 99.5127
R15067 VDD.n2453 VDD.n957 99.5127
R15068 VDD.n2461 VDD.n957 99.5127
R15069 VDD.n2461 VDD.n954 99.5127
R15070 VDD.n2466 VDD.n954 99.5127
R15071 VDD.n2466 VDD.n955 99.5127
R15072 VDD.n955 VDD.n940 99.5127
R15073 VDD.n2535 VDD.n940 99.5127
R15074 VDD.n2535 VDD.n941 99.5127
R15075 VDD.n2981 VDD.n2980 99.5127
R15076 VDD.n2978 VDD.n2956 99.5127
R15077 VDD.n2974 VDD.n2973 99.5127
R15078 VDD.n2971 VDD.n2959 99.5127
R15079 VDD.n2967 VDD.n2966 99.5127
R15080 VDD.n2964 VDD.n2962 99.5127
R15081 VDD.n3076 VDD.n3075 99.5127
R15082 VDD.n3073 VDD.n748 99.5127
R15083 VDD.n3069 VDD.n3068 99.5127
R15084 VDD.n3066 VDD.n751 99.5127
R15085 VDD.n3062 VDD.n3061 99.5127
R15086 VDD.n3059 VDD.n754 99.5127
R15087 VDD.n2790 VDD.n2593 99.5127
R15088 VDD.n2790 VDD.n898 99.5127
R15089 VDD.n2787 VDD.n898 99.5127
R15090 VDD.n2787 VDD.n892 99.5127
R15091 VDD.n2784 VDD.n892 99.5127
R15092 VDD.n2784 VDD.n887 99.5127
R15093 VDD.n2781 VDD.n887 99.5127
R15094 VDD.n2781 VDD.n881 99.5127
R15095 VDD.n2778 VDD.n881 99.5127
R15096 VDD.n2778 VDD.n875 99.5127
R15097 VDD.n2775 VDD.n875 99.5127
R15098 VDD.n2775 VDD.n870 99.5127
R15099 VDD.n2772 VDD.n870 99.5127
R15100 VDD.n2772 VDD.n864 99.5127
R15101 VDD.n2769 VDD.n864 99.5127
R15102 VDD.n2769 VDD.n858 99.5127
R15103 VDD.n2725 VDD.n858 99.5127
R15104 VDD.n2725 VDD.n853 99.5127
R15105 VDD.n2758 VDD.n853 99.5127
R15106 VDD.n2758 VDD.n846 99.5127
R15107 VDD.n2754 VDD.n846 99.5127
R15108 VDD.n2754 VDD.n840 99.5127
R15109 VDD.n2751 VDD.n840 99.5127
R15110 VDD.n2751 VDD.n834 99.5127
R15111 VDD.n2748 VDD.n834 99.5127
R15112 VDD.n2748 VDD.n828 99.5127
R15113 VDD.n2745 VDD.n828 99.5127
R15114 VDD.n2745 VDD.n822 99.5127
R15115 VDD.n2742 VDD.n822 99.5127
R15116 VDD.n2742 VDD.n817 99.5127
R15117 VDD.n2739 VDD.n817 99.5127
R15118 VDD.n2739 VDD.n812 99.5127
R15119 VDD.n2736 VDD.n812 99.5127
R15120 VDD.n2736 VDD.n806 99.5127
R15121 VDD.n2733 VDD.n806 99.5127
R15122 VDD.n2733 VDD.n798 99.5127
R15123 VDD.n2730 VDD.n798 99.5127
R15124 VDD.n2730 VDD.n791 99.5127
R15125 VDD.n791 VDD.n760 99.5127
R15126 VDD.n3054 VDD.n760 99.5127
R15127 VDD.n2842 VDD.n2840 99.5127
R15128 VDD.n2838 VDD.n2597 99.5127
R15129 VDD.n2834 VDD.n2832 99.5127
R15130 VDD.n2830 VDD.n2599 99.5127
R15131 VDD.n2826 VDD.n2824 99.5127
R15132 VDD.n2822 VDD.n2601 99.5127
R15133 VDD.n2818 VDD.n2816 99.5127
R15134 VDD.n2814 VDD.n2603 99.5127
R15135 VDD.n2810 VDD.n2808 99.5127
R15136 VDD.n2806 VDD.n2605 99.5127
R15137 VDD.n2802 VDD.n2800 99.5127
R15138 VDD.n2798 VDD.n2607 99.5127
R15139 VDD.n2846 VDD.n896 99.5127
R15140 VDD.n2854 VDD.n896 99.5127
R15141 VDD.n2854 VDD.n894 99.5127
R15142 VDD.n2858 VDD.n894 99.5127
R15143 VDD.n2858 VDD.n885 99.5127
R15144 VDD.n2866 VDD.n885 99.5127
R15145 VDD.n2866 VDD.n883 99.5127
R15146 VDD.n2870 VDD.n883 99.5127
R15147 VDD.n2870 VDD.n873 99.5127
R15148 VDD.n2878 VDD.n873 99.5127
R15149 VDD.n2878 VDD.n871 99.5127
R15150 VDD.n2882 VDD.n871 99.5127
R15151 VDD.n2882 VDD.n861 99.5127
R15152 VDD.n2890 VDD.n861 99.5127
R15153 VDD.n2890 VDD.n859 99.5127
R15154 VDD.n2894 VDD.n859 99.5127
R15155 VDD.n2894 VDD.n850 99.5127
R15156 VDD.n2902 VDD.n850 99.5127
R15157 VDD.n2902 VDD.n848 99.5127
R15158 VDD.n2906 VDD.n848 99.5127
R15159 VDD.n2906 VDD.n838 99.5127
R15160 VDD.n2914 VDD.n838 99.5127
R15161 VDD.n2914 VDD.n836 99.5127
R15162 VDD.n2918 VDD.n836 99.5127
R15163 VDD.n2918 VDD.n826 99.5127
R15164 VDD.n2926 VDD.n826 99.5127
R15165 VDD.n2926 VDD.n824 99.5127
R15166 VDD.n2930 VDD.n824 99.5127
R15167 VDD.n2930 VDD.n815 99.5127
R15168 VDD.n2938 VDD.n815 99.5127
R15169 VDD.n2938 VDD.n813 99.5127
R15170 VDD.n2942 VDD.n813 99.5127
R15171 VDD.n2942 VDD.n803 99.5127
R15172 VDD.n2950 VDD.n803 99.5127
R15173 VDD.n2950 VDD.n799 99.5127
R15174 VDD.n2991 VDD.n799 99.5127
R15175 VDD.n2991 VDD.n800 99.5127
R15176 VDD.n800 VDD.n792 99.5127
R15177 VDD.n2986 VDD.n792 99.5127
R15178 VDD.n2986 VDD.n763 99.5127
R15179 VDD.n2589 VDD.n931 99.5127
R15180 VDD.n2585 VDD.n2584 99.5127
R15181 VDD.n2581 VDD.n2580 99.5127
R15182 VDD.n2577 VDD.n2576 99.5127
R15183 VDD.n2573 VDD.n2572 99.5127
R15184 VDD.n2569 VDD.n2568 99.5127
R15185 VDD.n2565 VDD.n2564 99.5127
R15186 VDD.n2561 VDD.n2560 99.5127
R15187 VDD.n2557 VDD.n2556 99.5127
R15188 VDD.n2553 VDD.n2552 99.5127
R15189 VDD.n2549 VDD.n2548 99.5127
R15190 VDD.n2545 VDD.n2544 99.5127
R15191 VDD.n2541 VDD.n929 99.5127
R15192 VDD.n2191 VDD.n1061 99.5127
R15193 VDD.n2191 VDD.n1054 99.5127
R15194 VDD.n2194 VDD.n1054 99.5127
R15195 VDD.n2194 VDD.n1047 99.5127
R15196 VDD.n2197 VDD.n1047 99.5127
R15197 VDD.n2197 VDD.n1041 99.5127
R15198 VDD.n2200 VDD.n1041 99.5127
R15199 VDD.n2200 VDD.n1036 99.5127
R15200 VDD.n2203 VDD.n1036 99.5127
R15201 VDD.n2203 VDD.n1030 99.5127
R15202 VDD.n2206 VDD.n1030 99.5127
R15203 VDD.n2206 VDD.n1024 99.5127
R15204 VDD.n2209 VDD.n1024 99.5127
R15205 VDD.n2209 VDD.n1018 99.5127
R15206 VDD.n2212 VDD.n1018 99.5127
R15207 VDD.n2212 VDD.n1012 99.5127
R15208 VDD.n2215 VDD.n1012 99.5127
R15209 VDD.n2215 VDD.n1006 99.5127
R15210 VDD.n2218 VDD.n1006 99.5127
R15211 VDD.n2218 VDD.n1000 99.5127
R15212 VDD.n2269 VDD.n1000 99.5127
R15213 VDD.n2269 VDD.n994 99.5127
R15214 VDD.n2265 VDD.n994 99.5127
R15215 VDD.n2265 VDD.n989 99.5127
R15216 VDD.n2262 VDD.n989 99.5127
R15217 VDD.n2262 VDD.n983 99.5127
R15218 VDD.n2237 VDD.n983 99.5127
R15219 VDD.n2237 VDD.n977 99.5127
R15220 VDD.n2234 VDD.n977 99.5127
R15221 VDD.n2234 VDD.n971 99.5127
R15222 VDD.n2231 VDD.n971 99.5127
R15223 VDD.n2231 VDD.n966 99.5127
R15224 VDD.n2228 VDD.n966 99.5127
R15225 VDD.n2228 VDD.n960 99.5127
R15226 VDD.n2225 VDD.n960 99.5127
R15227 VDD.n2225 VDD.n953 99.5127
R15228 VDD.n2222 VDD.n953 99.5127
R15229 VDD.n2222 VDD.n937 99.5127
R15230 VDD.n2537 VDD.n937 99.5127
R15231 VDD.n2538 VDD.n2537 99.5127
R15232 VDD.n2140 VDD.n1058 99.5127
R15233 VDD.n2144 VDD.n2138 99.5127
R15234 VDD.n2148 VDD.n2146 99.5127
R15235 VDD.n2152 VDD.n2136 99.5127
R15236 VDD.n2156 VDD.n2154 99.5127
R15237 VDD.n2160 VDD.n2134 99.5127
R15238 VDD.n2164 VDD.n2162 99.5127
R15239 VDD.n2168 VDD.n1087 99.5127
R15240 VDD.n2172 VDD.n2170 99.5127
R15241 VDD.n2176 VDD.n1085 99.5127
R15242 VDD.n2180 VDD.n2178 99.5127
R15243 VDD.n2185 VDD.n1081 99.5127
R15244 VDD.n2188 VDD.n2187 99.5127
R15245 VDD.n2358 VDD.n1056 99.5127
R15246 VDD.n2362 VDD.n1056 99.5127
R15247 VDD.n2362 VDD.n1045 99.5127
R15248 VDD.n2370 VDD.n1045 99.5127
R15249 VDD.n2370 VDD.n1042 99.5127
R15250 VDD.n2375 VDD.n1042 99.5127
R15251 VDD.n2375 VDD.n1033 99.5127
R15252 VDD.n2383 VDD.n1033 99.5127
R15253 VDD.n2383 VDD.n1031 99.5127
R15254 VDD.n2387 VDD.n1031 99.5127
R15255 VDD.n2387 VDD.n1021 99.5127
R15256 VDD.n2395 VDD.n1021 99.5127
R15257 VDD.n2395 VDD.n1019 99.5127
R15258 VDD.n2399 VDD.n1019 99.5127
R15259 VDD.n2399 VDD.n1009 99.5127
R15260 VDD.n2407 VDD.n1009 99.5127
R15261 VDD.n2407 VDD.n1007 99.5127
R15262 VDD.n2411 VDD.n1007 99.5127
R15263 VDD.n2411 VDD.n997 99.5127
R15264 VDD.n2419 VDD.n997 99.5127
R15265 VDD.n2419 VDD.n995 99.5127
R15266 VDD.n2423 VDD.n995 99.5127
R15267 VDD.n2423 VDD.n986 99.5127
R15268 VDD.n2431 VDD.n986 99.5127
R15269 VDD.n2431 VDD.n984 99.5127
R15270 VDD.n2435 VDD.n984 99.5127
R15271 VDD.n2435 VDD.n974 99.5127
R15272 VDD.n2443 VDD.n974 99.5127
R15273 VDD.n2443 VDD.n972 99.5127
R15274 VDD.n2447 VDD.n972 99.5127
R15275 VDD.n2447 VDD.n963 99.5127
R15276 VDD.n2455 VDD.n963 99.5127
R15277 VDD.n2455 VDD.n961 99.5127
R15278 VDD.n2459 VDD.n961 99.5127
R15279 VDD.n2459 VDD.n950 99.5127
R15280 VDD.n2468 VDD.n950 99.5127
R15281 VDD.n2468 VDD.n948 99.5127
R15282 VDD.n2473 VDD.n948 99.5127
R15283 VDD.n2473 VDD.n939 99.5127
R15284 VDD.n939 VDD.n930 99.5127
R15285 VDD.t208 VDD.t206 89.2165
R15286 VDD.t149 VDD.n266 85.8723
R15287 VDD.t160 VDD.n215 85.8723
R15288 VDD.t138 VDD.n172 85.8723
R15289 VDD.t148 VDD.n121 85.8723
R15290 VDD.t128 VDD.n79 85.8723
R15291 VDD.t177 VDD.n28 85.8723
R15292 VDD.t185 VDD.n1755 85.8723
R15293 VDD.t176 VDD.n1806 85.8723
R15294 VDD.t174 VDD.n1661 85.8723
R15295 VDD.t167 VDD.n1712 85.8723
R15296 VDD.t153 VDD.n1568 85.8723
R15297 VDD.t102 VDD.n1619 85.8723
R15298 VDD.n2952 VDD.n801 78.546
R15299 VDD.n2373 VDD.n1043 78.546
R15300 VDD.n253 VDD.n252 75.1835
R15301 VDD.n251 VDD.n250 75.1835
R15302 VDD.n249 VDD.n248 75.1835
R15303 VDD.n247 VDD.n246 75.1835
R15304 VDD.n245 VDD.n244 75.1835
R15305 VDD.n159 VDD.n158 75.1835
R15306 VDD.n157 VDD.n156 75.1835
R15307 VDD.n155 VDD.n154 75.1835
R15308 VDD.n153 VDD.n152 75.1835
R15309 VDD.n151 VDD.n150 75.1835
R15310 VDD.n66 VDD.n65 75.1835
R15311 VDD.n64 VDD.n63 75.1835
R15312 VDD.n62 VDD.n61 75.1835
R15313 VDD.n60 VDD.n59 75.1835
R15314 VDD.n58 VDD.n57 75.1835
R15315 VDD.n1785 VDD.n1784 75.1835
R15316 VDD.n1787 VDD.n1786 75.1835
R15317 VDD.n1789 VDD.n1788 75.1835
R15318 VDD.n1791 VDD.n1790 75.1835
R15319 VDD.n1793 VDD.n1792 75.1835
R15320 VDD.n1691 VDD.n1690 75.1835
R15321 VDD.n1693 VDD.n1692 75.1835
R15322 VDD.n1695 VDD.n1694 75.1835
R15323 VDD.n1697 VDD.n1696 75.1835
R15324 VDD.n1699 VDD.n1698 75.1835
R15325 VDD.n1598 VDD.n1597 75.1835
R15326 VDD.n1600 VDD.n1599 75.1835
R15327 VDD.n1602 VDD.n1601 75.1835
R15328 VDD.n1604 VDD.n1603 75.1835
R15329 VDD.n1606 VDD.n1605 75.1835
R15330 VDD.n2841 VDD.n2591 72.8958
R15331 VDD.n2839 VDD.n2591 72.8958
R15332 VDD.n2833 VDD.n2591 72.8958
R15333 VDD.n2831 VDD.n2591 72.8958
R15334 VDD.n2825 VDD.n2591 72.8958
R15335 VDD.n2823 VDD.n2591 72.8958
R15336 VDD.n2817 VDD.n2591 72.8958
R15337 VDD.n2815 VDD.n2591 72.8958
R15338 VDD.n2809 VDD.n2591 72.8958
R15339 VDD.n2807 VDD.n2591 72.8958
R15340 VDD.n2801 VDD.n2591 72.8958
R15341 VDD.n2799 VDD.n2591 72.8958
R15342 VDD.n2793 VDD.n2591 72.8958
R15343 VDD.n759 VDD.n662 72.8958
R15344 VDD.n3060 VDD.n662 72.8958
R15345 VDD.n753 VDD.n662 72.8958
R15346 VDD.n3067 VDD.n662 72.8958
R15347 VDD.n750 VDD.n662 72.8958
R15348 VDD.n3074 VDD.n662 72.8958
R15349 VDD.n747 VDD.n662 72.8958
R15350 VDD.n2965 VDD.n662 72.8958
R15351 VDD.n2961 VDD.n662 72.8958
R15352 VDD.n2972 VDD.n662 72.8958
R15353 VDD.n2958 VDD.n662 72.8958
R15354 VDD.n2979 VDD.n662 72.8958
R15355 VDD.n2982 VDD.n662 72.8958
R15356 VDD.n2351 VDD.n1059 72.8958
R15357 VDD.n1064 VDD.n1059 72.8958
R15358 VDD.n2344 VDD.n1059 72.8958
R15359 VDD.n2338 VDD.n1059 72.8958
R15360 VDD.n2336 VDD.n1059 72.8958
R15361 VDD.n2330 VDD.n1059 72.8958
R15362 VDD.n1070 VDD.n1059 72.8958
R15363 VDD.n2324 VDD.n1059 72.8958
R15364 VDD.n2318 VDD.n1059 72.8958
R15365 VDD.n2316 VDD.n1059 72.8958
R15366 VDD.n2310 VDD.n1059 72.8958
R15367 VDD.n1078 VDD.n1059 72.8958
R15368 VDD.n2590 VDD.n916 72.8958
R15369 VDD.n2590 VDD.n915 72.8958
R15370 VDD.n2590 VDD.n914 72.8958
R15371 VDD.n2590 VDD.n913 72.8958
R15372 VDD.n2590 VDD.n912 72.8958
R15373 VDD.n2590 VDD.n911 72.8958
R15374 VDD.n2590 VDD.n910 72.8958
R15375 VDD.n2590 VDD.n909 72.8958
R15376 VDD.n2590 VDD.n908 72.8958
R15377 VDD.n2590 VDD.n907 72.8958
R15378 VDD.n2590 VDD.n906 72.8958
R15379 VDD.n2590 VDD.n905 72.8958
R15380 VDD.n2590 VDD.n904 72.8958
R15381 VDD.n2626 VDD.n2591 72.8958
R15382 VDD.n2632 VDD.n2591 72.8958
R15383 VDD.n2634 VDD.n2591 72.8958
R15384 VDD.n2640 VDD.n2591 72.8958
R15385 VDD.n2642 VDD.n2591 72.8958
R15386 VDD.n2648 VDD.n2591 72.8958
R15387 VDD.n2650 VDD.n2591 72.8958
R15388 VDD.n2656 VDD.n2591 72.8958
R15389 VDD.n2658 VDD.n2591 72.8958
R15390 VDD.n2664 VDD.n2591 72.8958
R15391 VDD.n2666 VDD.n2591 72.8958
R15392 VDD.n2673 VDD.n2591 72.8958
R15393 VDD.n3003 VDD.n662 72.8958
R15394 VDD.n3009 VDD.n662 72.8958
R15395 VDD.n783 VDD.n662 72.8958
R15396 VDD.n3016 VDD.n662 72.8958
R15397 VDD.n780 VDD.n662 72.8958
R15398 VDD.n3023 VDD.n662 72.8958
R15399 VDD.n777 VDD.n662 72.8958
R15400 VDD.n3032 VDD.n662 72.8958
R15401 VDD.n774 VDD.n662 72.8958
R15402 VDD.n3039 VDD.n662 72.8958
R15403 VDD.n771 VDD.n662 72.8958
R15404 VDD.n3046 VDD.n662 72.8958
R15405 VDD.n768 VDD.n662 72.8958
R15406 VDD.n2590 VDD.n928 72.8958
R15407 VDD.n2590 VDD.n927 72.8958
R15408 VDD.n2590 VDD.n926 72.8958
R15409 VDD.n2590 VDD.n925 72.8958
R15410 VDD.n2590 VDD.n924 72.8958
R15411 VDD.n2590 VDD.n923 72.8958
R15412 VDD.n2590 VDD.n922 72.8958
R15413 VDD.n2590 VDD.n921 72.8958
R15414 VDD.n2590 VDD.n920 72.8958
R15415 VDD.n2590 VDD.n919 72.8958
R15416 VDD.n2590 VDD.n918 72.8958
R15417 VDD.n2590 VDD.n917 72.8958
R15418 VDD.n2139 VDD.n1059 72.8958
R15419 VDD.n2145 VDD.n1059 72.8958
R15420 VDD.n2147 VDD.n1059 72.8958
R15421 VDD.n2153 VDD.n1059 72.8958
R15422 VDD.n2155 VDD.n1059 72.8958
R15423 VDD.n2161 VDD.n1059 72.8958
R15424 VDD.n2163 VDD.n1059 72.8958
R15425 VDD.n2169 VDD.n1059 72.8958
R15426 VDD.n2171 VDD.n1059 72.8958
R15427 VDD.n2177 VDD.n1059 72.8958
R15428 VDD.n2179 VDD.n1059 72.8958
R15429 VDD.n2186 VDD.n1059 72.8958
R15430 VDD.n1309 VDD.n1237 66.2847
R15431 VDD.n1317 VDD.n1237 66.2847
R15432 VDD.n1319 VDD.n1237 66.2847
R15433 VDD.n1327 VDD.n1237 66.2847
R15434 VDD.n1329 VDD.n1237 66.2847
R15435 VDD.n1337 VDD.n1237 66.2847
R15436 VDD.n1339 VDD.n1237 66.2847
R15437 VDD.n1349 VDD.n1237 66.2847
R15438 VDD.n1352 VDD.n1237 66.2847
R15439 VDD.n1288 VDD.n1237 66.2847
R15440 VDD.n1361 VDD.n1237 66.2847
R15441 VDD.n1363 VDD.n1237 66.2847
R15442 VDD.n1371 VDD.n1237 66.2847
R15443 VDD.n1373 VDD.n1237 66.2847
R15444 VDD.n1381 VDD.n1237 66.2847
R15445 VDD.n1383 VDD.n1237 66.2847
R15446 VDD.n1391 VDD.n1237 66.2847
R15447 VDD.n1393 VDD.n1237 66.2847
R15448 VDD.n1403 VDD.n1237 66.2847
R15449 VDD.n1406 VDD.n1237 66.2847
R15450 VDD.n1263 VDD.n1237 66.2847
R15451 VDD.n1415 VDD.n1237 66.2847
R15452 VDD.n1417 VDD.n1237 66.2847
R15453 VDD.n1425 VDD.n1237 66.2847
R15454 VDD.n1427 VDD.n1237 66.2847
R15455 VDD.n1435 VDD.n1237 66.2847
R15456 VDD.n1437 VDD.n1237 66.2847
R15457 VDD.n1445 VDD.n1237 66.2847
R15458 VDD.n1447 VDD.n1237 66.2847
R15459 VDD.n1457 VDD.n1237 66.2847
R15460 VDD.n1460 VDD.n1237 66.2847
R15461 VDD.n1113 VDD.n1105 66.2847
R15462 VDD.n1113 VDD.n1112 66.2847
R15463 VDD.n1113 VDD.n1111 66.2847
R15464 VDD.n1113 VDD.n1109 66.2847
R15465 VDD.n2013 VDD.n1113 66.2847
R15466 VDD.n2018 VDD.n1113 66.2847
R15467 VDD.n2011 VDD.n1113 66.2847
R15468 VDD.n2025 VDD.n1113 66.2847
R15469 VDD.n2005 VDD.n1113 66.2847
R15470 VDD.n2032 VDD.n1113 66.2847
R15471 VDD.n1999 VDD.n1113 66.2847
R15472 VDD.n1994 VDD.n1113 66.2847
R15473 VDD.n2043 VDD.n1113 66.2847
R15474 VDD.n1986 VDD.n1113 66.2847
R15475 VDD.n2050 VDD.n1113 66.2847
R15476 VDD.n1979 VDD.n1113 66.2847
R15477 VDD.n2057 VDD.n1113 66.2847
R15478 VDD.n1972 VDD.n1113 66.2847
R15479 VDD.n2064 VDD.n1113 66.2847
R15480 VDD.n1965 VDD.n1113 66.2847
R15481 VDD.n2071 VDD.n1113 66.2847
R15482 VDD.n1959 VDD.n1113 66.2847
R15483 VDD.n1954 VDD.n1113 66.2847
R15484 VDD.n2082 VDD.n1113 66.2847
R15485 VDD.n1946 VDD.n1113 66.2847
R15486 VDD.n2089 VDD.n1113 66.2847
R15487 VDD.n1940 VDD.n1113 66.2847
R15488 VDD.n1937 VDD.n1113 66.2847
R15489 VDD.n2099 VDD.n1113 66.2847
R15490 VDD.n1929 VDD.n1113 66.2847
R15491 VDD.n2106 VDD.n1113 66.2847
R15492 VDD.n1922 VDD.n1113 66.2847
R15493 VDD.n3216 VDD.n3215 66.2847
R15494 VDD.n3216 VDD.n663 66.2847
R15495 VDD.n3216 VDD.n664 66.2847
R15496 VDD.n3216 VDD.n665 66.2847
R15497 VDD.n3216 VDD.n666 66.2847
R15498 VDD.n3216 VDD.n667 66.2847
R15499 VDD.n3216 VDD.n668 66.2847
R15500 VDD.n3216 VDD.n669 66.2847
R15501 VDD.n3216 VDD.n670 66.2847
R15502 VDD.n3216 VDD.n671 66.2847
R15503 VDD.n3216 VDD.n672 66.2847
R15504 VDD.n3216 VDD.n673 66.2847
R15505 VDD.n3216 VDD.n674 66.2847
R15506 VDD.n3216 VDD.n675 66.2847
R15507 VDD.n3216 VDD.n676 66.2847
R15508 VDD.n3216 VDD.n677 66.2847
R15509 VDD.n3216 VDD.n678 66.2847
R15510 VDD.n3216 VDD.n679 66.2847
R15511 VDD.n3216 VDD.n680 66.2847
R15512 VDD.n3216 VDD.n681 66.2847
R15513 VDD.n3216 VDD.n682 66.2847
R15514 VDD.n3216 VDD.n683 66.2847
R15515 VDD.n3216 VDD.n684 66.2847
R15516 VDD.n3216 VDD.n685 66.2847
R15517 VDD.n3216 VDD.n686 66.2847
R15518 VDD.n3216 VDD.n687 66.2847
R15519 VDD.n3216 VDD.n688 66.2847
R15520 VDD.n3216 VDD.n689 66.2847
R15521 VDD.n3216 VDD.n690 66.2847
R15522 VDD.n3216 VDD.n691 66.2847
R15523 VDD.n3216 VDD.n692 66.2847
R15524 VDD.n3347 VDD.n3346 66.2847
R15525 VDD.n3347 VDD.n390 66.2847
R15526 VDD.n3347 VDD.n389 66.2847
R15527 VDD.n3347 VDD.n388 66.2847
R15528 VDD.n3347 VDD.n387 66.2847
R15529 VDD.n3347 VDD.n386 66.2847
R15530 VDD.n3347 VDD.n385 66.2847
R15531 VDD.n3347 VDD.n384 66.2847
R15532 VDD.n3347 VDD.n383 66.2847
R15533 VDD.n3347 VDD.n382 66.2847
R15534 VDD.n3347 VDD.n381 66.2847
R15535 VDD.n3347 VDD.n380 66.2847
R15536 VDD.n3347 VDD.n379 66.2847
R15537 VDD.n3347 VDD.n378 66.2847
R15538 VDD.n3347 VDD.n377 66.2847
R15539 VDD.n3347 VDD.n376 66.2847
R15540 VDD.n3347 VDD.n375 66.2847
R15541 VDD.n3347 VDD.n374 66.2847
R15542 VDD.n3347 VDD.n373 66.2847
R15543 VDD.n3347 VDD.n372 66.2847
R15544 VDD.n3347 VDD.n371 66.2847
R15545 VDD.n3347 VDD.n370 66.2847
R15546 VDD.n3347 VDD.n369 66.2847
R15547 VDD.n3347 VDD.n368 66.2847
R15548 VDD.n3347 VDD.n367 66.2847
R15549 VDD.n3347 VDD.n366 66.2847
R15550 VDD.n3347 VDD.n365 66.2847
R15551 VDD.n3347 VDD.n364 66.2847
R15552 VDD.n3347 VDD.n363 66.2847
R15553 VDD.n3347 VDD.n362 66.2847
R15554 VDD.n3347 VDD.n361 66.2847
R15555 VDD.n3347 VDD.n360 66.2847
R15556 VDD.n435 VDD.n360 52.4337
R15557 VDD.n441 VDD.n361 52.4337
R15558 VDD.n445 VDD.n362 52.4337
R15559 VDD.n451 VDD.n363 52.4337
R15560 VDD.n455 VDD.n364 52.4337
R15561 VDD.n461 VDD.n365 52.4337
R15562 VDD.n465 VDD.n366 52.4337
R15563 VDD.n471 VDD.n367 52.4337
R15564 VDD.n475 VDD.n368 52.4337
R15565 VDD.n481 VDD.n369 52.4337
R15566 VDD.n485 VDD.n370 52.4337
R15567 VDD.n491 VDD.n371 52.4337
R15568 VDD.n495 VDD.n372 52.4337
R15569 VDD.n501 VDD.n373 52.4337
R15570 VDD.n505 VDD.n374 52.4337
R15571 VDD.n511 VDD.n375 52.4337
R15572 VDD.n515 VDD.n376 52.4337
R15573 VDD.n521 VDD.n377 52.4337
R15574 VDD.n525 VDD.n378 52.4337
R15575 VDD.n531 VDD.n379 52.4337
R15576 VDD.n535 VDD.n380 52.4337
R15577 VDD.n541 VDD.n381 52.4337
R15578 VDD.n545 VDD.n382 52.4337
R15579 VDD.n551 VDD.n383 52.4337
R15580 VDD.n555 VDD.n384 52.4337
R15581 VDD.n561 VDD.n385 52.4337
R15582 VDD.n565 VDD.n386 52.4337
R15583 VDD.n571 VDD.n387 52.4337
R15584 VDD.n575 VDD.n388 52.4337
R15585 VDD.n581 VDD.n389 52.4337
R15586 VDD.n584 VDD.n390 52.4337
R15587 VDD.n3346 VDD.n3345 52.4337
R15588 VDD.n3215 VDD.n3214 52.4337
R15589 VDD.n3209 VDD.n663 52.4337
R15590 VDD.n3206 VDD.n664 52.4337
R15591 VDD.n3202 VDD.n665 52.4337
R15592 VDD.n3198 VDD.n666 52.4337
R15593 VDD.n3194 VDD.n667 52.4337
R15594 VDD.n3190 VDD.n668 52.4337
R15595 VDD.n3186 VDD.n669 52.4337
R15596 VDD.n3182 VDD.n670 52.4337
R15597 VDD.n3178 VDD.n671 52.4337
R15598 VDD.n3170 VDD.n672 52.4337
R15599 VDD.n3166 VDD.n673 52.4337
R15600 VDD.n3162 VDD.n674 52.4337
R15601 VDD.n3158 VDD.n675 52.4337
R15602 VDD.n3154 VDD.n676 52.4337
R15603 VDD.n3150 VDD.n677 52.4337
R15604 VDD.n3146 VDD.n678 52.4337
R15605 VDD.n3142 VDD.n679 52.4337
R15606 VDD.n3138 VDD.n680 52.4337
R15607 VDD.n3134 VDD.n681 52.4337
R15608 VDD.n3130 VDD.n682 52.4337
R15609 VDD.n3124 VDD.n683 52.4337
R15610 VDD.n3120 VDD.n684 52.4337
R15611 VDD.n3116 VDD.n685 52.4337
R15612 VDD.n3112 VDD.n686 52.4337
R15613 VDD.n3108 VDD.n687 52.4337
R15614 VDD.n3104 VDD.n688 52.4337
R15615 VDD.n3100 VDD.n689 52.4337
R15616 VDD.n3096 VDD.n690 52.4337
R15617 VDD.n3092 VDD.n691 52.4337
R15618 VDD.n3088 VDD.n692 52.4337
R15619 VDD.n2108 VDD.n1922 52.4337
R15620 VDD.n2106 VDD.n2105 52.4337
R15621 VDD.n2101 VDD.n1929 52.4337
R15622 VDD.n2099 VDD.n2098 52.4337
R15623 VDD.n1938 VDD.n1937 52.4337
R15624 VDD.n2091 VDD.n1940 52.4337
R15625 VDD.n2089 VDD.n2088 52.4337
R15626 VDD.n2084 VDD.n1946 52.4337
R15627 VDD.n2082 VDD.n2081 52.4337
R15628 VDD.n1955 VDD.n1954 52.4337
R15629 VDD.n2073 VDD.n1959 52.4337
R15630 VDD.n2071 VDD.n2070 52.4337
R15631 VDD.n2066 VDD.n1965 52.4337
R15632 VDD.n2064 VDD.n2063 52.4337
R15633 VDD.n2059 VDD.n1972 52.4337
R15634 VDD.n2057 VDD.n2056 52.4337
R15635 VDD.n2052 VDD.n1979 52.4337
R15636 VDD.n2050 VDD.n2049 52.4337
R15637 VDD.n2045 VDD.n1986 52.4337
R15638 VDD.n2043 VDD.n2042 52.4337
R15639 VDD.n1995 VDD.n1994 52.4337
R15640 VDD.n2034 VDD.n1999 52.4337
R15641 VDD.n2032 VDD.n2031 52.4337
R15642 VDD.n2027 VDD.n2005 52.4337
R15643 VDD.n2025 VDD.n2024 52.4337
R15644 VDD.n2020 VDD.n2011 52.4337
R15645 VDD.n2018 VDD.n2017 52.4337
R15646 VDD.n2013 VDD.n2012 52.4337
R15647 VDD.n1109 VDD.n1094 52.4337
R15648 VDD.n1111 VDD.n1110 52.4337
R15649 VDD.n1112 VDD.n1099 52.4337
R15650 VDD.n2117 VDD.n1105 52.4337
R15651 VDD.n1309 VDD.n1236 52.4337
R15652 VDD.n1317 VDD.n1316 52.4337
R15653 VDD.n1320 VDD.n1319 52.4337
R15654 VDD.n1327 VDD.n1326 52.4337
R15655 VDD.n1330 VDD.n1329 52.4337
R15656 VDD.n1337 VDD.n1336 52.4337
R15657 VDD.n1340 VDD.n1339 52.4337
R15658 VDD.n1349 VDD.n1348 52.4337
R15659 VDD.n1352 VDD.n1351 52.4337
R15660 VDD.n1289 VDD.n1288 52.4337
R15661 VDD.n1361 VDD.n1360 52.4337
R15662 VDD.n1364 VDD.n1363 52.4337
R15663 VDD.n1371 VDD.n1370 52.4337
R15664 VDD.n1374 VDD.n1373 52.4337
R15665 VDD.n1381 VDD.n1380 52.4337
R15666 VDD.n1384 VDD.n1383 52.4337
R15667 VDD.n1391 VDD.n1390 52.4337
R15668 VDD.n1394 VDD.n1393 52.4337
R15669 VDD.n1403 VDD.n1402 52.4337
R15670 VDD.n1406 VDD.n1405 52.4337
R15671 VDD.n1264 VDD.n1263 52.4337
R15672 VDD.n1415 VDD.n1414 52.4337
R15673 VDD.n1418 VDD.n1417 52.4337
R15674 VDD.n1425 VDD.n1424 52.4337
R15675 VDD.n1428 VDD.n1427 52.4337
R15676 VDD.n1435 VDD.n1434 52.4337
R15677 VDD.n1438 VDD.n1437 52.4337
R15678 VDD.n1445 VDD.n1444 52.4337
R15679 VDD.n1448 VDD.n1447 52.4337
R15680 VDD.n1457 VDD.n1456 52.4337
R15681 VDD.n1460 VDD.n1459 52.4337
R15682 VDD.n1310 VDD.n1309 52.4337
R15683 VDD.n1318 VDD.n1317 52.4337
R15684 VDD.n1319 VDD.n1302 52.4337
R15685 VDD.n1328 VDD.n1327 52.4337
R15686 VDD.n1329 VDD.n1298 52.4337
R15687 VDD.n1338 VDD.n1337 52.4337
R15688 VDD.n1339 VDD.n1294 52.4337
R15689 VDD.n1350 VDD.n1349 52.4337
R15690 VDD.n1353 VDD.n1352 52.4337
R15691 VDD.n1288 VDD.n1285 52.4337
R15692 VDD.n1362 VDD.n1361 52.4337
R15693 VDD.n1363 VDD.n1281 52.4337
R15694 VDD.n1372 VDD.n1371 52.4337
R15695 VDD.n1373 VDD.n1277 52.4337
R15696 VDD.n1382 VDD.n1381 52.4337
R15697 VDD.n1383 VDD.n1273 52.4337
R15698 VDD.n1392 VDD.n1391 52.4337
R15699 VDD.n1393 VDD.n1269 52.4337
R15700 VDD.n1404 VDD.n1403 52.4337
R15701 VDD.n1407 VDD.n1406 52.4337
R15702 VDD.n1263 VDD.n1260 52.4337
R15703 VDD.n1416 VDD.n1415 52.4337
R15704 VDD.n1417 VDD.n1256 52.4337
R15705 VDD.n1426 VDD.n1425 52.4337
R15706 VDD.n1427 VDD.n1252 52.4337
R15707 VDD.n1436 VDD.n1435 52.4337
R15708 VDD.n1437 VDD.n1248 52.4337
R15709 VDD.n1446 VDD.n1445 52.4337
R15710 VDD.n1447 VDD.n1244 52.4337
R15711 VDD.n1458 VDD.n1457 52.4337
R15712 VDD.n1461 VDD.n1460 52.4337
R15713 VDD.n1105 VDD.n1100 52.4337
R15714 VDD.n1112 VDD.n1098 52.4337
R15715 VDD.n1111 VDD.n1095 52.4337
R15716 VDD.n1109 VDD.n1093 52.4337
R15717 VDD.n2014 VDD.n2013 52.4337
R15718 VDD.n2019 VDD.n2018 52.4337
R15719 VDD.n2011 VDD.n2006 52.4337
R15720 VDD.n2026 VDD.n2025 52.4337
R15721 VDD.n2005 VDD.n2000 52.4337
R15722 VDD.n2033 VDD.n2032 52.4337
R15723 VDD.n1999 VDD.n1998 52.4337
R15724 VDD.n1994 VDD.n1987 52.4337
R15725 VDD.n2044 VDD.n2043 52.4337
R15726 VDD.n1986 VDD.n1980 52.4337
R15727 VDD.n2051 VDD.n2050 52.4337
R15728 VDD.n1979 VDD.n1973 52.4337
R15729 VDD.n2058 VDD.n2057 52.4337
R15730 VDD.n1972 VDD.n1966 52.4337
R15731 VDD.n2065 VDD.n2064 52.4337
R15732 VDD.n1965 VDD.n1960 52.4337
R15733 VDD.n2072 VDD.n2071 52.4337
R15734 VDD.n1959 VDD.n1958 52.4337
R15735 VDD.n1954 VDD.n1947 52.4337
R15736 VDD.n2083 VDD.n2082 52.4337
R15737 VDD.n1946 VDD.n1941 52.4337
R15738 VDD.n2090 VDD.n2089 52.4337
R15739 VDD.n1940 VDD.n1939 52.4337
R15740 VDD.n1937 VDD.n1930 52.4337
R15741 VDD.n2100 VDD.n2099 52.4337
R15742 VDD.n1929 VDD.n1923 52.4337
R15743 VDD.n2107 VDD.n2106 52.4337
R15744 VDD.n1922 VDD.n1115 52.4337
R15745 VDD.n3215 VDD.n694 52.4337
R15746 VDD.n3207 VDD.n663 52.4337
R15747 VDD.n3203 VDD.n664 52.4337
R15748 VDD.n3199 VDD.n665 52.4337
R15749 VDD.n3195 VDD.n666 52.4337
R15750 VDD.n3191 VDD.n667 52.4337
R15751 VDD.n3187 VDD.n668 52.4337
R15752 VDD.n3183 VDD.n669 52.4337
R15753 VDD.n3179 VDD.n670 52.4337
R15754 VDD.n3169 VDD.n671 52.4337
R15755 VDD.n3167 VDD.n672 52.4337
R15756 VDD.n3163 VDD.n673 52.4337
R15757 VDD.n3159 VDD.n674 52.4337
R15758 VDD.n3155 VDD.n675 52.4337
R15759 VDD.n3151 VDD.n676 52.4337
R15760 VDD.n3147 VDD.n677 52.4337
R15761 VDD.n3143 VDD.n678 52.4337
R15762 VDD.n3139 VDD.n679 52.4337
R15763 VDD.n3135 VDD.n680 52.4337
R15764 VDD.n3131 VDD.n681 52.4337
R15765 VDD.n3123 VDD.n682 52.4337
R15766 VDD.n3121 VDD.n683 52.4337
R15767 VDD.n3117 VDD.n684 52.4337
R15768 VDD.n3113 VDD.n685 52.4337
R15769 VDD.n3109 VDD.n686 52.4337
R15770 VDD.n3105 VDD.n687 52.4337
R15771 VDD.n3101 VDD.n688 52.4337
R15772 VDD.n3097 VDD.n689 52.4337
R15773 VDD.n3093 VDD.n690 52.4337
R15774 VDD.n3089 VDD.n691 52.4337
R15775 VDD.n692 VDD.n661 52.4337
R15776 VDD.n3346 VDD.n391 52.4337
R15777 VDD.n582 VDD.n390 52.4337
R15778 VDD.n576 VDD.n389 52.4337
R15779 VDD.n572 VDD.n388 52.4337
R15780 VDD.n566 VDD.n387 52.4337
R15781 VDD.n562 VDD.n386 52.4337
R15782 VDD.n556 VDD.n385 52.4337
R15783 VDD.n552 VDD.n384 52.4337
R15784 VDD.n546 VDD.n383 52.4337
R15785 VDD.n542 VDD.n382 52.4337
R15786 VDD.n536 VDD.n381 52.4337
R15787 VDD.n532 VDD.n380 52.4337
R15788 VDD.n526 VDD.n379 52.4337
R15789 VDD.n522 VDD.n378 52.4337
R15790 VDD.n516 VDD.n377 52.4337
R15791 VDD.n512 VDD.n376 52.4337
R15792 VDD.n506 VDD.n375 52.4337
R15793 VDD.n502 VDD.n374 52.4337
R15794 VDD.n496 VDD.n373 52.4337
R15795 VDD.n492 VDD.n372 52.4337
R15796 VDD.n486 VDD.n371 52.4337
R15797 VDD.n482 VDD.n370 52.4337
R15798 VDD.n476 VDD.n369 52.4337
R15799 VDD.n472 VDD.n368 52.4337
R15800 VDD.n466 VDD.n367 52.4337
R15801 VDD.n462 VDD.n366 52.4337
R15802 VDD.n456 VDD.n365 52.4337
R15803 VDD.n452 VDD.n364 52.4337
R15804 VDD.n446 VDD.n363 52.4337
R15805 VDD.n442 VDD.n362 52.4337
R15806 VDD.n436 VDD.n361 52.4337
R15807 VDD.n432 VDD.n360 52.4337
R15808 VDD.n245 VDD.n243 42.2617
R15809 VDD.n151 VDD.n149 42.2617
R15810 VDD.n58 VDD.n56 42.2617
R15811 VDD.n1785 VDD.n1783 42.2617
R15812 VDD.n1691 VDD.n1689 42.2617
R15813 VDD.n1598 VDD.n1596 42.2617
R15814 VDD.n295 VDD.n294 41.6884
R15815 VDD.n201 VDD.n200 41.6884
R15816 VDD.n108 VDD.n107 41.6884
R15817 VDD.n1835 VDD.n1834 41.6884
R15818 VDD.n1741 VDD.n1740 41.6884
R15819 VDD.n1648 VDD.n1647 41.6884
R15820 VDD.n3048 VDD.n768 39.2114
R15821 VDD.n3046 VDD.n3045 39.2114
R15822 VDD.n3041 VDD.n771 39.2114
R15823 VDD.n3039 VDD.n3038 39.2114
R15824 VDD.n3034 VDD.n774 39.2114
R15825 VDD.n3032 VDD.n3031 39.2114
R15826 VDD.n3025 VDD.n777 39.2114
R15827 VDD.n3023 VDD.n3022 39.2114
R15828 VDD.n3018 VDD.n780 39.2114
R15829 VDD.n3016 VDD.n3015 39.2114
R15830 VDD.n3011 VDD.n783 39.2114
R15831 VDD.n3009 VDD.n3008 39.2114
R15832 VDD.n3004 VDD.n3003 39.2114
R15833 VDD.n2626 VDD.n902 39.2114
R15834 VDD.n2632 VDD.n2631 39.2114
R15835 VDD.n2635 VDD.n2634 39.2114
R15836 VDD.n2640 VDD.n2639 39.2114
R15837 VDD.n2643 VDD.n2642 39.2114
R15838 VDD.n2648 VDD.n2647 39.2114
R15839 VDD.n2651 VDD.n2650 39.2114
R15840 VDD.n2656 VDD.n2655 39.2114
R15841 VDD.n2659 VDD.n2658 39.2114
R15842 VDD.n2664 VDD.n2663 39.2114
R15843 VDD.n2667 VDD.n2666 39.2114
R15844 VDD.n2673 VDD.n2672 39.2114
R15845 VDD.n2529 VDD.n904 39.2114
R15846 VDD.n2525 VDD.n905 39.2114
R15847 VDD.n2521 VDD.n906 39.2114
R15848 VDD.n2517 VDD.n907 39.2114
R15849 VDD.n2513 VDD.n908 39.2114
R15850 VDD.n2509 VDD.n909 39.2114
R15851 VDD.n2505 VDD.n910 39.2114
R15852 VDD.n2501 VDD.n911 39.2114
R15853 VDD.n2497 VDD.n912 39.2114
R15854 VDD.n2493 VDD.n913 39.2114
R15855 VDD.n2489 VDD.n914 39.2114
R15856 VDD.n2484 VDD.n915 39.2114
R15857 VDD.n2480 VDD.n916 39.2114
R15858 VDD.n2351 VDD.n1062 39.2114
R15859 VDD.n2349 VDD.n1064 39.2114
R15860 VDD.n2345 VDD.n2344 39.2114
R15861 VDD.n2338 VDD.n1066 39.2114
R15862 VDD.n2337 VDD.n2336 39.2114
R15863 VDD.n2330 VDD.n1068 39.2114
R15864 VDD.n2329 VDD.n1070 39.2114
R15865 VDD.n2325 VDD.n2324 39.2114
R15866 VDD.n2318 VDD.n1072 39.2114
R15867 VDD.n2317 VDD.n2316 39.2114
R15868 VDD.n2310 VDD.n1074 39.2114
R15869 VDD.n2309 VDD.n1078 39.2114
R15870 VDD.n2982 VDD.n2981 39.2114
R15871 VDD.n2979 VDD.n2978 39.2114
R15872 VDD.n2974 VDD.n2958 39.2114
R15873 VDD.n2972 VDD.n2971 39.2114
R15874 VDD.n2967 VDD.n2961 39.2114
R15875 VDD.n2965 VDD.n2964 39.2114
R15876 VDD.n3076 VDD.n747 39.2114
R15877 VDD.n3074 VDD.n3073 39.2114
R15878 VDD.n3069 VDD.n750 39.2114
R15879 VDD.n3067 VDD.n3066 39.2114
R15880 VDD.n3062 VDD.n753 39.2114
R15881 VDD.n3060 VDD.n3059 39.2114
R15882 VDD.n3055 VDD.n759 39.2114
R15883 VDD.n2841 VDD.n2595 39.2114
R15884 VDD.n2840 VDD.n2839 39.2114
R15885 VDD.n2833 VDD.n2597 39.2114
R15886 VDD.n2832 VDD.n2831 39.2114
R15887 VDD.n2825 VDD.n2599 39.2114
R15888 VDD.n2824 VDD.n2823 39.2114
R15889 VDD.n2817 VDD.n2601 39.2114
R15890 VDD.n2816 VDD.n2815 39.2114
R15891 VDD.n2809 VDD.n2603 39.2114
R15892 VDD.n2808 VDD.n2807 39.2114
R15893 VDD.n2801 VDD.n2605 39.2114
R15894 VDD.n2800 VDD.n2799 39.2114
R15895 VDD.n2793 VDD.n2607 39.2114
R15896 VDD.n2842 VDD.n2841 39.2114
R15897 VDD.n2839 VDD.n2838 39.2114
R15898 VDD.n2834 VDD.n2833 39.2114
R15899 VDD.n2831 VDD.n2830 39.2114
R15900 VDD.n2826 VDD.n2825 39.2114
R15901 VDD.n2823 VDD.n2822 39.2114
R15902 VDD.n2818 VDD.n2817 39.2114
R15903 VDD.n2815 VDD.n2814 39.2114
R15904 VDD.n2810 VDD.n2809 39.2114
R15905 VDD.n2807 VDD.n2806 39.2114
R15906 VDD.n2802 VDD.n2801 39.2114
R15907 VDD.n2799 VDD.n2798 39.2114
R15908 VDD.n2794 VDD.n2793 39.2114
R15909 VDD.n759 VDD.n754 39.2114
R15910 VDD.n3061 VDD.n3060 39.2114
R15911 VDD.n753 VDD.n751 39.2114
R15912 VDD.n3068 VDD.n3067 39.2114
R15913 VDD.n750 VDD.n748 39.2114
R15914 VDD.n3075 VDD.n3074 39.2114
R15915 VDD.n2962 VDD.n747 39.2114
R15916 VDD.n2966 VDD.n2965 39.2114
R15917 VDD.n2961 VDD.n2959 39.2114
R15918 VDD.n2973 VDD.n2972 39.2114
R15919 VDD.n2958 VDD.n2956 39.2114
R15920 VDD.n2980 VDD.n2979 39.2114
R15921 VDD.n2983 VDD.n2982 39.2114
R15922 VDD.n2352 VDD.n2351 39.2114
R15923 VDD.n2346 VDD.n1064 39.2114
R15924 VDD.n2344 VDD.n2343 39.2114
R15925 VDD.n2339 VDD.n2338 39.2114
R15926 VDD.n2336 VDD.n2335 39.2114
R15927 VDD.n2331 VDD.n2330 39.2114
R15928 VDD.n2326 VDD.n1070 39.2114
R15929 VDD.n2324 VDD.n2323 39.2114
R15930 VDD.n2319 VDD.n2318 39.2114
R15931 VDD.n2316 VDD.n2315 39.2114
R15932 VDD.n2311 VDD.n2310 39.2114
R15933 VDD.n2306 VDD.n1078 39.2114
R15934 VDD.n2483 VDD.n916 39.2114
R15935 VDD.n2488 VDD.n915 39.2114
R15936 VDD.n2492 VDD.n914 39.2114
R15937 VDD.n2496 VDD.n913 39.2114
R15938 VDD.n2500 VDD.n912 39.2114
R15939 VDD.n2504 VDD.n911 39.2114
R15940 VDD.n2508 VDD.n910 39.2114
R15941 VDD.n2512 VDD.n909 39.2114
R15942 VDD.n2516 VDD.n908 39.2114
R15943 VDD.n2520 VDD.n907 39.2114
R15944 VDD.n2524 VDD.n906 39.2114
R15945 VDD.n2528 VDD.n905 39.2114
R15946 VDD.n2531 VDD.n904 39.2114
R15947 VDD.n2627 VDD.n2626 39.2114
R15948 VDD.n2633 VDD.n2632 39.2114
R15949 VDD.n2634 VDD.n2623 39.2114
R15950 VDD.n2641 VDD.n2640 39.2114
R15951 VDD.n2642 VDD.n2621 39.2114
R15952 VDD.n2649 VDD.n2648 39.2114
R15953 VDD.n2650 VDD.n2619 39.2114
R15954 VDD.n2657 VDD.n2656 39.2114
R15955 VDD.n2658 VDD.n2617 39.2114
R15956 VDD.n2665 VDD.n2664 39.2114
R15957 VDD.n2666 VDD.n2613 39.2114
R15958 VDD.n2674 VDD.n2673 39.2114
R15959 VDD.n3003 VDD.n784 39.2114
R15960 VDD.n3010 VDD.n3009 39.2114
R15961 VDD.n783 VDD.n781 39.2114
R15962 VDD.n3017 VDD.n3016 39.2114
R15963 VDD.n780 VDD.n778 39.2114
R15964 VDD.n3024 VDD.n3023 39.2114
R15965 VDD.n777 VDD.n775 39.2114
R15966 VDD.n3033 VDD.n3032 39.2114
R15967 VDD.n774 VDD.n772 39.2114
R15968 VDD.n3040 VDD.n3039 39.2114
R15969 VDD.n771 VDD.n769 39.2114
R15970 VDD.n3047 VDD.n3046 39.2114
R15971 VDD.n768 VDD.n765 39.2114
R15972 VDD.n931 VDD.n917 39.2114
R15973 VDD.n2584 VDD.n918 39.2114
R15974 VDD.n2580 VDD.n919 39.2114
R15975 VDD.n2576 VDD.n920 39.2114
R15976 VDD.n2572 VDD.n921 39.2114
R15977 VDD.n2568 VDD.n922 39.2114
R15978 VDD.n2564 VDD.n923 39.2114
R15979 VDD.n2560 VDD.n924 39.2114
R15980 VDD.n2556 VDD.n925 39.2114
R15981 VDD.n2552 VDD.n926 39.2114
R15982 VDD.n2548 VDD.n927 39.2114
R15983 VDD.n2544 VDD.n928 39.2114
R15984 VDD.n2140 VDD.n2139 39.2114
R15985 VDD.n2145 VDD.n2144 39.2114
R15986 VDD.n2148 VDD.n2147 39.2114
R15987 VDD.n2153 VDD.n2152 39.2114
R15988 VDD.n2156 VDD.n2155 39.2114
R15989 VDD.n2161 VDD.n2160 39.2114
R15990 VDD.n2164 VDD.n2163 39.2114
R15991 VDD.n2169 VDD.n2168 39.2114
R15992 VDD.n2172 VDD.n2171 39.2114
R15993 VDD.n2177 VDD.n2176 39.2114
R15994 VDD.n2180 VDD.n2179 39.2114
R15995 VDD.n2186 VDD.n2185 39.2114
R15996 VDD.n2541 VDD.n928 39.2114
R15997 VDD.n2545 VDD.n927 39.2114
R15998 VDD.n2549 VDD.n926 39.2114
R15999 VDD.n2553 VDD.n925 39.2114
R16000 VDD.n2557 VDD.n924 39.2114
R16001 VDD.n2561 VDD.n923 39.2114
R16002 VDD.n2565 VDD.n922 39.2114
R16003 VDD.n2569 VDD.n921 39.2114
R16004 VDD.n2573 VDD.n920 39.2114
R16005 VDD.n2577 VDD.n919 39.2114
R16006 VDD.n2581 VDD.n918 39.2114
R16007 VDD.n2585 VDD.n917 39.2114
R16008 VDD.n2139 VDD.n2138 39.2114
R16009 VDD.n2146 VDD.n2145 39.2114
R16010 VDD.n2147 VDD.n2136 39.2114
R16011 VDD.n2154 VDD.n2153 39.2114
R16012 VDD.n2155 VDD.n2134 39.2114
R16013 VDD.n2162 VDD.n2161 39.2114
R16014 VDD.n2163 VDD.n1087 39.2114
R16015 VDD.n2170 VDD.n2169 39.2114
R16016 VDD.n2171 VDD.n1085 39.2114
R16017 VDD.n2178 VDD.n2177 39.2114
R16018 VDD.n2179 VDD.n1081 39.2114
R16019 VDD.n2187 VDD.n2186 39.2114
R16020 VDD.n1463 VDD.n1241 37.4308
R16021 VDD.n1409 VDD.n1266 37.4308
R16022 VDD.n1355 VDD.n1291 37.4308
R16023 VDD.n1103 VDD.n1102 37.4308
R16024 VDD.n2039 VDD.n1993 37.4308
R16025 VDD.n2078 VDD.n1953 37.4308
R16026 VDD.n394 VDD.n393 37.4308
R16027 VDD.n534 VDD.n407 37.4308
R16028 VDD.n420 VDD.n419 37.4308
R16029 VDD.n3129 VDD.n734 37.4308
R16030 VDD.n3177 VDD.n3176 37.4308
R16031 VDD.n660 VDD.n659 37.4308
R16032 VDD.n2533 VDD.n2532 31.3761
R16033 VDD.n2481 VDD.n2478 31.3761
R16034 VDD.n2304 VDD.n2303 31.3761
R16035 VDD.n2355 VDD.n2354 31.3761
R16036 VDD.n2677 VDD.n2676 31.3761
R16037 VDD.n3005 VDD.n3002 31.3761
R16038 VDD.n2849 VDD.n901 31.3761
R16039 VDD.n3051 VDD.n3050 31.3761
R16040 VDD.n2985 VDD.n2984 31.3761
R16041 VDD.n3056 VDD.n758 31.3761
R16042 VDD.n2795 VDD.n2792 31.3761
R16043 VDD.n2845 VDD.n2844 31.3761
R16044 VDD.n2359 VDD.n1057 31.3761
R16045 VDD.n2588 VDD.n932 31.3761
R16046 VDD.n2540 VDD.n2539 31.3761
R16047 VDD.n2190 VDD.n2189 31.3761
R16048 VDD.n2183 VDD.n1083 30.449
R16049 VDD.n935 VDD.n934 30.449
R16050 VDD.n1077 VDD.n1076 30.449
R16051 VDD.n2486 VDD.n944 30.449
R16052 VDD.n2610 VDD.n2609 30.449
R16053 VDD.n787 VDD.n786 30.449
R16054 VDD.n2670 VDD.n2615 30.449
R16055 VDD.n757 VDD.n756 30.449
R16056 VDD.n1083 VDD.n1082 25.7944
R16057 VDD.n934 VDD.n933 25.7944
R16058 VDD.n1241 VDD.n1240 25.7944
R16059 VDD.n1266 VDD.n1265 25.7944
R16060 VDD.n1291 VDD.n1290 25.7944
R16061 VDD.n1076 VDD.n1075 25.7944
R16062 VDD.n1102 VDD.n1101 25.7944
R16063 VDD.n1993 VDD.n1992 25.7944
R16064 VDD.n1953 VDD.n1952 25.7944
R16065 VDD.n944 VDD.n943 25.7944
R16066 VDD.n2609 VDD.n2608 25.7944
R16067 VDD.n393 VDD.n392 25.7944
R16068 VDD.n407 VDD.n406 25.7944
R16069 VDD.n419 VDD.n418 25.7944
R16070 VDD.n734 VDD.n733 25.7944
R16071 VDD.n3176 VDD.n3175 25.7944
R16072 VDD.n786 VDD.n785 25.7944
R16073 VDD.n2615 VDD.n2614 25.7944
R16074 VDD.n659 VDD.n658 25.7944
R16075 VDD.n756 VDD.n755 25.7944
R16076 VDD.n1470 VDD.n1237 23.6004
R16077 VDD.n2115 VDD.n1113 23.6004
R16078 VDD.n3216 VDD.n654 23.6004
R16079 VDD.n3348 VDD.n3347 23.6004
R16080 VDD.n1467 VDD.n1231 19.3944
R16081 VDD.n1480 VDD.n1231 19.3944
R16082 VDD.n1480 VDD.n1229 19.3944
R16083 VDD.n1484 VDD.n1229 19.3944
R16084 VDD.n1484 VDD.n1219 19.3944
R16085 VDD.n1496 VDD.n1219 19.3944
R16086 VDD.n1496 VDD.n1217 19.3944
R16087 VDD.n1500 VDD.n1217 19.3944
R16088 VDD.n1500 VDD.n1207 19.3944
R16089 VDD.n1513 VDD.n1207 19.3944
R16090 VDD.n1513 VDD.n1205 19.3944
R16091 VDD.n1517 VDD.n1205 19.3944
R16092 VDD.n1517 VDD.n1196 19.3944
R16093 VDD.n1529 VDD.n1196 19.3944
R16094 VDD.n1529 VDD.n1194 19.3944
R16095 VDD.n1533 VDD.n1194 19.3944
R16096 VDD.n1533 VDD.n1184 19.3944
R16097 VDD.n1546 VDD.n1184 19.3944
R16098 VDD.n1546 VDD.n1182 19.3944
R16099 VDD.n1550 VDD.n1182 19.3944
R16100 VDD.n1550 VDD.n1173 19.3944
R16101 VDD.n1844 VDD.n1173 19.3944
R16102 VDD.n1844 VDD.n1171 19.3944
R16103 VDD.n1848 VDD.n1171 19.3944
R16104 VDD.n1848 VDD.n1160 19.3944
R16105 VDD.n1860 VDD.n1160 19.3944
R16106 VDD.n1860 VDD.n1158 19.3944
R16107 VDD.n1864 VDD.n1158 19.3944
R16108 VDD.n1864 VDD.n1149 19.3944
R16109 VDD.n1876 VDD.n1149 19.3944
R16110 VDD.n1876 VDD.n1147 19.3944
R16111 VDD.n1880 VDD.n1147 19.3944
R16112 VDD.n1880 VDD.n1136 19.3944
R16113 VDD.n1892 VDD.n1136 19.3944
R16114 VDD.n1892 VDD.n1134 19.3944
R16115 VDD.n1896 VDD.n1134 19.3944
R16116 VDD.n1896 VDD.n1125 19.3944
R16117 VDD.n1908 VDD.n1125 19.3944
R16118 VDD.n1908 VDD.n1122 19.3944
R16119 VDD.n1913 VDD.n1122 19.3944
R16120 VDD.n1913 VDD.n1123 19.3944
R16121 VDD.n1123 VDD.n1107 19.3944
R16122 VDD.n1413 VDD.n1261 19.3944
R16123 VDD.n1413 VDD.n1259 19.3944
R16124 VDD.n1419 VDD.n1259 19.3944
R16125 VDD.n1419 VDD.n1257 19.3944
R16126 VDD.n1423 VDD.n1257 19.3944
R16127 VDD.n1423 VDD.n1255 19.3944
R16128 VDD.n1429 VDD.n1255 19.3944
R16129 VDD.n1429 VDD.n1253 19.3944
R16130 VDD.n1433 VDD.n1253 19.3944
R16131 VDD.n1433 VDD.n1251 19.3944
R16132 VDD.n1439 VDD.n1251 19.3944
R16133 VDD.n1439 VDD.n1249 19.3944
R16134 VDD.n1443 VDD.n1249 19.3944
R16135 VDD.n1443 VDD.n1247 19.3944
R16136 VDD.n1449 VDD.n1247 19.3944
R16137 VDD.n1449 VDD.n1245 19.3944
R16138 VDD.n1455 VDD.n1245 19.3944
R16139 VDD.n1455 VDD.n1243 19.3944
R16140 VDD.n1243 VDD.n1242 19.3944
R16141 VDD.n1462 VDD.n1242 19.3944
R16142 VDD.n1359 VDD.n1286 19.3944
R16143 VDD.n1359 VDD.n1284 19.3944
R16144 VDD.n1365 VDD.n1284 19.3944
R16145 VDD.n1365 VDD.n1282 19.3944
R16146 VDD.n1369 VDD.n1282 19.3944
R16147 VDD.n1369 VDD.n1280 19.3944
R16148 VDD.n1375 VDD.n1280 19.3944
R16149 VDD.n1375 VDD.n1278 19.3944
R16150 VDD.n1379 VDD.n1278 19.3944
R16151 VDD.n1379 VDD.n1276 19.3944
R16152 VDD.n1385 VDD.n1276 19.3944
R16153 VDD.n1385 VDD.n1274 19.3944
R16154 VDD.n1389 VDD.n1274 19.3944
R16155 VDD.n1389 VDD.n1272 19.3944
R16156 VDD.n1395 VDD.n1272 19.3944
R16157 VDD.n1395 VDD.n1270 19.3944
R16158 VDD.n1401 VDD.n1270 19.3944
R16159 VDD.n1401 VDD.n1268 19.3944
R16160 VDD.n1268 VDD.n1267 19.3944
R16161 VDD.n1408 VDD.n1267 19.3944
R16162 VDD.n1311 VDD.n1308 19.3944
R16163 VDD.n1311 VDD.n1307 19.3944
R16164 VDD.n1315 VDD.n1307 19.3944
R16165 VDD.n1315 VDD.n1305 19.3944
R16166 VDD.n1321 VDD.n1305 19.3944
R16167 VDD.n1321 VDD.n1303 19.3944
R16168 VDD.n1325 VDD.n1303 19.3944
R16169 VDD.n1325 VDD.n1301 19.3944
R16170 VDD.n1331 VDD.n1301 19.3944
R16171 VDD.n1331 VDD.n1299 19.3944
R16172 VDD.n1335 VDD.n1299 19.3944
R16173 VDD.n1335 VDD.n1297 19.3944
R16174 VDD.n1341 VDD.n1297 19.3944
R16175 VDD.n1341 VDD.n1295 19.3944
R16176 VDD.n1347 VDD.n1295 19.3944
R16177 VDD.n1347 VDD.n1293 19.3944
R16178 VDD.n1293 VDD.n1292 19.3944
R16179 VDD.n1354 VDD.n1292 19.3944
R16180 VDD.n1472 VDD.n1234 19.3944
R16181 VDD.n1476 VDD.n1234 19.3944
R16182 VDD.n1476 VDD.n1225 19.3944
R16183 VDD.n1488 VDD.n1225 19.3944
R16184 VDD.n1488 VDD.n1223 19.3944
R16185 VDD.n1492 VDD.n1223 19.3944
R16186 VDD.n1492 VDD.n1213 19.3944
R16187 VDD.n1505 VDD.n1213 19.3944
R16188 VDD.n1505 VDD.n1211 19.3944
R16189 VDD.n1509 VDD.n1211 19.3944
R16190 VDD.n1509 VDD.n1202 19.3944
R16191 VDD.n1521 VDD.n1202 19.3944
R16192 VDD.n1521 VDD.n1200 19.3944
R16193 VDD.n1525 VDD.n1200 19.3944
R16194 VDD.n1525 VDD.n1190 19.3944
R16195 VDD.n1538 VDD.n1190 19.3944
R16196 VDD.n1538 VDD.n1188 19.3944
R16197 VDD.n1542 VDD.n1188 19.3944
R16198 VDD.n1542 VDD.n1179 19.3944
R16199 VDD.n1554 VDD.n1179 19.3944
R16200 VDD.n1554 VDD.n1177 19.3944
R16201 VDD.n1840 VDD.n1177 19.3944
R16202 VDD.n1840 VDD.n1167 19.3944
R16203 VDD.n1852 VDD.n1167 19.3944
R16204 VDD.n1852 VDD.n1165 19.3944
R16205 VDD.n1856 VDD.n1165 19.3944
R16206 VDD.n1856 VDD.n1155 19.3944
R16207 VDD.n1868 VDD.n1155 19.3944
R16208 VDD.n1868 VDD.n1153 19.3944
R16209 VDD.n1872 VDD.n1153 19.3944
R16210 VDD.n1872 VDD.n1143 19.3944
R16211 VDD.n1884 VDD.n1143 19.3944
R16212 VDD.n1884 VDD.n1141 19.3944
R16213 VDD.n1888 VDD.n1141 19.3944
R16214 VDD.n1888 VDD.n1131 19.3944
R16215 VDD.n1900 VDD.n1131 19.3944
R16216 VDD.n1900 VDD.n1129 19.3944
R16217 VDD.n1904 VDD.n1129 19.3944
R16218 VDD.n1904 VDD.n1118 19.3944
R16219 VDD.n1917 VDD.n1118 19.3944
R16220 VDD.n1917 VDD.n1116 19.3944
R16221 VDD.n2113 VDD.n1116 19.3944
R16222 VDD.n2035 VDD.n1991 19.3944
R16223 VDD.n2035 VDD.n1997 19.3944
R16224 VDD.n2030 VDD.n1997 19.3944
R16225 VDD.n2030 VDD.n2029 19.3944
R16226 VDD.n2029 VDD.n2028 19.3944
R16227 VDD.n2028 VDD.n2004 19.3944
R16228 VDD.n2023 VDD.n2004 19.3944
R16229 VDD.n2023 VDD.n2022 19.3944
R16230 VDD.n2022 VDD.n2021 19.3944
R16231 VDD.n2021 VDD.n2010 19.3944
R16232 VDD.n2016 VDD.n2015 19.3944
R16233 VDD.n2129 VDD.n1092 19.3944
R16234 VDD.n2129 VDD.n2128 19.3944
R16235 VDD.n2128 VDD.n2127 19.3944
R16236 VDD.n2127 VDD.n1096 19.3944
R16237 VDD.n2123 VDD.n1096 19.3944
R16238 VDD.n2123 VDD.n2122 19.3944
R16239 VDD.n2122 VDD.n2121 19.3944
R16240 VDD.n2074 VDD.n1951 19.3944
R16241 VDD.n2074 VDD.n1957 19.3944
R16242 VDD.n2069 VDD.n1957 19.3944
R16243 VDD.n2069 VDD.n2068 19.3944
R16244 VDD.n2068 VDD.n2067 19.3944
R16245 VDD.n2067 VDD.n1964 19.3944
R16246 VDD.n2062 VDD.n1964 19.3944
R16247 VDD.n2062 VDD.n2061 19.3944
R16248 VDD.n2061 VDD.n2060 19.3944
R16249 VDD.n2060 VDD.n1971 19.3944
R16250 VDD.n2055 VDD.n1971 19.3944
R16251 VDD.n2055 VDD.n2054 19.3944
R16252 VDD.n2054 VDD.n2053 19.3944
R16253 VDD.n2053 VDD.n1978 19.3944
R16254 VDD.n2048 VDD.n1978 19.3944
R16255 VDD.n2048 VDD.n2047 19.3944
R16256 VDD.n2047 VDD.n2046 19.3944
R16257 VDD.n2046 VDD.n1985 19.3944
R16258 VDD.n2041 VDD.n1985 19.3944
R16259 VDD.n2041 VDD.n2040 19.3944
R16260 VDD.n2110 VDD.n2109 19.3944
R16261 VDD.n2109 VDD.n1921 19.3944
R16262 VDD.n2104 VDD.n1921 19.3944
R16263 VDD.n2104 VDD.n2103 19.3944
R16264 VDD.n2103 VDD.n2102 19.3944
R16265 VDD.n2102 VDD.n1928 19.3944
R16266 VDD.n2097 VDD.n1928 19.3944
R16267 VDD.n2097 VDD.n2096 19.3944
R16268 VDD.n1935 VDD.n1933 19.3944
R16269 VDD.n2092 VDD.n1936 19.3944
R16270 VDD.n2087 VDD.n1936 19.3944
R16271 VDD.n2087 VDD.n2086 19.3944
R16272 VDD.n2086 VDD.n2085 19.3944
R16273 VDD.n2085 VDD.n1945 19.3944
R16274 VDD.n2080 VDD.n1945 19.3944
R16275 VDD.n2080 VDD.n2079 19.3944
R16276 VDD.n3222 VDD.n656 19.3944
R16277 VDD.n3222 VDD.n646 19.3944
R16278 VDD.n3234 VDD.n646 19.3944
R16279 VDD.n3234 VDD.n644 19.3944
R16280 VDD.n3238 VDD.n644 19.3944
R16281 VDD.n3238 VDD.n635 19.3944
R16282 VDD.n3251 VDD.n635 19.3944
R16283 VDD.n3251 VDD.n633 19.3944
R16284 VDD.n3255 VDD.n633 19.3944
R16285 VDD.n3255 VDD.n623 19.3944
R16286 VDD.n3267 VDD.n623 19.3944
R16287 VDD.n3267 VDD.n621 19.3944
R16288 VDD.n3271 VDD.n621 19.3944
R16289 VDD.n3271 VDD.n612 19.3944
R16290 VDD.n3284 VDD.n612 19.3944
R16291 VDD.n3284 VDD.n610 19.3944
R16292 VDD.n3291 VDD.n610 19.3944
R16293 VDD.n3291 VDD.n3290 19.3944
R16294 VDD.n3290 VDD.n599 19.3944
R16295 VDD.n3304 VDD.n599 19.3944
R16296 VDD.n3305 VDD.n3304 19.3944
R16297 VDD.n3306 VDD.n3305 19.3944
R16298 VDD.n3306 VDD.n597 19.3944
R16299 VDD.n3311 VDD.n597 19.3944
R16300 VDD.n3312 VDD.n3311 19.3944
R16301 VDD.n3313 VDD.n3312 19.3944
R16302 VDD.n3313 VDD.n595 19.3944
R16303 VDD.n3318 VDD.n595 19.3944
R16304 VDD.n3319 VDD.n3318 19.3944
R16305 VDD.n3320 VDD.n3319 19.3944
R16306 VDD.n3320 VDD.n593 19.3944
R16307 VDD.n3325 VDD.n593 19.3944
R16308 VDD.n3326 VDD.n3325 19.3944
R16309 VDD.n3327 VDD.n3326 19.3944
R16310 VDD.n3327 VDD.n591 19.3944
R16311 VDD.n3332 VDD.n591 19.3944
R16312 VDD.n3333 VDD.n3332 19.3944
R16313 VDD.n3334 VDD.n3333 19.3944
R16314 VDD.n3334 VDD.n589 19.3944
R16315 VDD.n3339 VDD.n589 19.3944
R16316 VDD.n3340 VDD.n3339 19.3944
R16317 VDD.n3341 VDD.n3340 19.3944
R16318 VDD.n537 VDD.n404 19.3944
R16319 VDD.n543 VDD.n404 19.3944
R16320 VDD.n544 VDD.n543 19.3944
R16321 VDD.n547 VDD.n544 19.3944
R16322 VDD.n547 VDD.n402 19.3944
R16323 VDD.n553 VDD.n402 19.3944
R16324 VDD.n554 VDD.n553 19.3944
R16325 VDD.n557 VDD.n554 19.3944
R16326 VDD.n557 VDD.n400 19.3944
R16327 VDD.n563 VDD.n400 19.3944
R16328 VDD.n564 VDD.n563 19.3944
R16329 VDD.n567 VDD.n564 19.3944
R16330 VDD.n567 VDD.n398 19.3944
R16331 VDD.n573 VDD.n398 19.3944
R16332 VDD.n574 VDD.n573 19.3944
R16333 VDD.n577 VDD.n574 19.3944
R16334 VDD.n577 VDD.n396 19.3944
R16335 VDD.n583 VDD.n396 19.3944
R16336 VDD.n585 VDD.n583 19.3944
R16337 VDD.n586 VDD.n585 19.3944
R16338 VDD.n484 VDD.n483 19.3944
R16339 VDD.n487 VDD.n484 19.3944
R16340 VDD.n487 VDD.n416 19.3944
R16341 VDD.n493 VDD.n416 19.3944
R16342 VDD.n494 VDD.n493 19.3944
R16343 VDD.n497 VDD.n494 19.3944
R16344 VDD.n497 VDD.n414 19.3944
R16345 VDD.n503 VDD.n414 19.3944
R16346 VDD.n504 VDD.n503 19.3944
R16347 VDD.n507 VDD.n504 19.3944
R16348 VDD.n507 VDD.n412 19.3944
R16349 VDD.n513 VDD.n412 19.3944
R16350 VDD.n514 VDD.n513 19.3944
R16351 VDD.n517 VDD.n514 19.3944
R16352 VDD.n517 VDD.n410 19.3944
R16353 VDD.n523 VDD.n410 19.3944
R16354 VDD.n524 VDD.n523 19.3944
R16355 VDD.n527 VDD.n524 19.3944
R16356 VDD.n527 VDD.n408 19.3944
R16357 VDD.n533 VDD.n408 19.3944
R16358 VDD.n434 VDD.n433 19.3944
R16359 VDD.n437 VDD.n434 19.3944
R16360 VDD.n437 VDD.n428 19.3944
R16361 VDD.n443 VDD.n428 19.3944
R16362 VDD.n444 VDD.n443 19.3944
R16363 VDD.n447 VDD.n444 19.3944
R16364 VDD.n447 VDD.n426 19.3944
R16365 VDD.n453 VDD.n426 19.3944
R16366 VDD.n454 VDD.n453 19.3944
R16367 VDD.n457 VDD.n454 19.3944
R16368 VDD.n457 VDD.n424 19.3944
R16369 VDD.n463 VDD.n424 19.3944
R16370 VDD.n464 VDD.n463 19.3944
R16371 VDD.n467 VDD.n464 19.3944
R16372 VDD.n467 VDD.n422 19.3944
R16373 VDD.n473 VDD.n422 19.3944
R16374 VDD.n474 VDD.n473 19.3944
R16375 VDD.n477 VDD.n474 19.3944
R16376 VDD.n3226 VDD.n652 19.3944
R16377 VDD.n3226 VDD.n650 19.3944
R16378 VDD.n3230 VDD.n650 19.3944
R16379 VDD.n3230 VDD.n640 19.3944
R16380 VDD.n3243 VDD.n640 19.3944
R16381 VDD.n3243 VDD.n638 19.3944
R16382 VDD.n3247 VDD.n638 19.3944
R16383 VDD.n3247 VDD.n629 19.3944
R16384 VDD.n3259 VDD.n629 19.3944
R16385 VDD.n3259 VDD.n627 19.3944
R16386 VDD.n3263 VDD.n627 19.3944
R16387 VDD.n3263 VDD.n617 19.3944
R16388 VDD.n3276 VDD.n617 19.3944
R16389 VDD.n3276 VDD.n615 19.3944
R16390 VDD.n3280 VDD.n615 19.3944
R16391 VDD.n3280 VDD.n606 19.3944
R16392 VDD.n3295 VDD.n606 19.3944
R16393 VDD.n3295 VDD.n604 19.3944
R16394 VDD.n3299 VDD.n604 19.3944
R16395 VDD.n3299 VDD.n299 19.3944
R16396 VDD.n3391 VDD.n299 19.3944
R16397 VDD.n3391 VDD.n300 19.3944
R16398 VDD.n3385 VDD.n300 19.3944
R16399 VDD.n3385 VDD.n3384 19.3944
R16400 VDD.n3384 VDD.n3383 19.3944
R16401 VDD.n3383 VDD.n312 19.3944
R16402 VDD.n3377 VDD.n312 19.3944
R16403 VDD.n3377 VDD.n3376 19.3944
R16404 VDD.n3376 VDD.n3375 19.3944
R16405 VDD.n3375 VDD.n322 19.3944
R16406 VDD.n3369 VDD.n322 19.3944
R16407 VDD.n3369 VDD.n3368 19.3944
R16408 VDD.n3368 VDD.n3367 19.3944
R16409 VDD.n3367 VDD.n334 19.3944
R16410 VDD.n3361 VDD.n334 19.3944
R16411 VDD.n3361 VDD.n3360 19.3944
R16412 VDD.n3360 VDD.n3359 19.3944
R16413 VDD.n3359 VDD.n344 19.3944
R16414 VDD.n3353 VDD.n344 19.3944
R16415 VDD.n3353 VDD.n3352 19.3944
R16416 VDD.n3352 VDD.n3351 19.3944
R16417 VDD.n3351 VDD.n356 19.3944
R16418 VDD.n3171 VDD.n712 19.3944
R16419 VDD.n3171 VDD.n3168 19.3944
R16420 VDD.n3168 VDD.n3165 19.3944
R16421 VDD.n3165 VDD.n3164 19.3944
R16422 VDD.n3164 VDD.n3161 19.3944
R16423 VDD.n3161 VDD.n3160 19.3944
R16424 VDD.n3160 VDD.n3157 19.3944
R16425 VDD.n3157 VDD.n3156 19.3944
R16426 VDD.n3156 VDD.n3153 19.3944
R16427 VDD.n3153 VDD.n3152 19.3944
R16428 VDD.n3152 VDD.n3149 19.3944
R16429 VDD.n3149 VDD.n3148 19.3944
R16430 VDD.n3148 VDD.n3145 19.3944
R16431 VDD.n3145 VDD.n3144 19.3944
R16432 VDD.n3144 VDD.n3141 19.3944
R16433 VDD.n3141 VDD.n3140 19.3944
R16434 VDD.n3140 VDD.n3137 19.3944
R16435 VDD.n3137 VDD.n3136 19.3944
R16436 VDD.n3136 VDD.n3133 19.3944
R16437 VDD.n3133 VDD.n3132 19.3944
R16438 VDD.n3213 VDD.n3212 19.3944
R16439 VDD.n3212 VDD.n3211 19.3944
R16440 VDD.n3211 VDD.n3210 19.3944
R16441 VDD.n3210 VDD.n3208 19.3944
R16442 VDD.n3208 VDD.n3205 19.3944
R16443 VDD.n3205 VDD.n3204 19.3944
R16444 VDD.n3204 VDD.n3201 19.3944
R16445 VDD.n3201 VDD.n3200 19.3944
R16446 VDD.n3197 VDD.n3196 19.3944
R16447 VDD.n3193 VDD.n3192 19.3944
R16448 VDD.n3192 VDD.n3189 19.3944
R16449 VDD.n3189 VDD.n3188 19.3944
R16450 VDD.n3188 VDD.n3185 19.3944
R16451 VDD.n3185 VDD.n3184 19.3944
R16452 VDD.n3184 VDD.n3181 19.3944
R16453 VDD.n3181 VDD.n3180 19.3944
R16454 VDD.n3125 VDD.n732 19.3944
R16455 VDD.n3125 VDD.n3122 19.3944
R16456 VDD.n3122 VDD.n3119 19.3944
R16457 VDD.n3119 VDD.n3118 19.3944
R16458 VDD.n3118 VDD.n3115 19.3944
R16459 VDD.n3115 VDD.n3114 19.3944
R16460 VDD.n3114 VDD.n3111 19.3944
R16461 VDD.n3111 VDD.n3110 19.3944
R16462 VDD.n3110 VDD.n3107 19.3944
R16463 VDD.n3107 VDD.n3106 19.3944
R16464 VDD.n3103 VDD.n3102 19.3944
R16465 VDD.n3099 VDD.n3098 19.3944
R16466 VDD.n3098 VDD.n3095 19.3944
R16467 VDD.n3095 VDD.n3094 19.3944
R16468 VDD.n3094 VDD.n3091 19.3944
R16469 VDD.n3091 VDD.n3090 19.3944
R16470 VDD.n3090 VDD.n3087 19.3944
R16471 VDD.n3087 VDD.n3086 19.3944
R16472 VDD.n1409 VDD.n1261 19.0066
R16473 VDD.n2039 VDD.n1991 19.0066
R16474 VDD.n537 VDD.n534 19.0066
R16475 VDD.n3129 VDD.n732 19.0066
R16476 VDD.n2357 VDD.n1059 16.3704
R16477 VDD.n2590 VDD.n903 16.3704
R16478 VDD.n2847 VDD.n2591 16.3704
R16479 VDD.n3053 VDD.n662 16.3704
R16480 VDD.n1470 VDD.n1469 13.6421
R16481 VDD.n1478 VDD.n1227 13.6421
R16482 VDD.n1486 VDD.n1227 13.6421
R16483 VDD.n1486 VDD.n1221 13.6421
R16484 VDD.n1494 VDD.n1221 13.6421
R16485 VDD.n1503 VDD.n1215 13.6421
R16486 VDD.n1503 VDD.n1502 13.6421
R16487 VDD.n1511 VDD.n1209 13.6421
R16488 VDD.n1519 VDD.n1198 13.6421
R16489 VDD.n1527 VDD.n1198 13.6421
R16490 VDD.n1536 VDD.n1192 13.6421
R16491 VDD.n1536 VDD.n1535 13.6421
R16492 VDD.n1544 VDD.n1186 13.6421
R16493 VDD.n1552 VDD.n1175 13.6421
R16494 VDD.n1842 VDD.n1175 13.6421
R16495 VDD.n1850 VDD.n1169 13.6421
R16496 VDD.n1858 VDD.n1162 13.6421
R16497 VDD.n1858 VDD.n1163 13.6421
R16498 VDD.n1866 VDD.n1151 13.6421
R16499 VDD.n1874 VDD.n1151 13.6421
R16500 VDD.n1882 VDD.n1145 13.6421
R16501 VDD.n1890 VDD.n1138 13.6421
R16502 VDD.n1890 VDD.n1139 13.6421
R16503 VDD.n1898 VDD.n1127 13.6421
R16504 VDD.n1906 VDD.n1127 13.6421
R16505 VDD.n1906 VDD.n1120 13.6421
R16506 VDD.n1915 VDD.n1120 13.6421
R16507 VDD.n2115 VDD.n1108 13.6421
R16508 VDD.n3224 VDD.n654 13.6421
R16509 VDD.n3232 VDD.n648 13.6421
R16510 VDD.n3232 VDD.n642 13.6421
R16511 VDD.n3241 VDD.n642 13.6421
R16512 VDD.n3241 VDD.n3240 13.6421
R16513 VDD.n3249 VDD.n631 13.6421
R16514 VDD.n3257 VDD.n631 13.6421
R16515 VDD.n3265 VDD.n625 13.6421
R16516 VDD.n3274 VDD.n619 13.6421
R16517 VDD.n3274 VDD.n3273 13.6421
R16518 VDD.n3282 VDD.n608 13.6421
R16519 VDD.n3293 VDD.n608 13.6421
R16520 VDD.n3301 VDD.n602 13.6421
R16521 VDD.n3389 VDD.n303 13.6421
R16522 VDD.n3389 VDD.n3388 13.6421
R16523 VDD.n3387 VDD.n307 13.6421
R16524 VDD.n3381 VDD.n3380 13.6421
R16525 VDD.n3380 VDD.n3379 13.6421
R16526 VDD.n3373 VDD.n324 13.6421
R16527 VDD.n3373 VDD.n3372 13.6421
R16528 VDD.n3371 VDD.n328 13.6421
R16529 VDD.n3365 VDD.n3364 13.6421
R16530 VDD.n3364 VDD.n3363 13.6421
R16531 VDD.n3357 VDD.n346 13.6421
R16532 VDD.n3357 VDD.n3356 13.6421
R16533 VDD.n3356 VDD.n3355 13.6421
R16534 VDD.n3355 VDD.n350 13.6421
R16535 VDD.n3349 VDD.n3348 13.6421
R16536 VDD.n1544 VDD.t117 13.5057
R16537 VDD.n1850 VDD.t113 13.5057
R16538 VDD.t97 VDD.n602 13.5057
R16539 VDD.t110 VDD.n307 13.5057
R16540 VDD.n1511 VDD.t131 13.2328
R16541 VDD.n1882 VDD.t99 13.2328
R16542 VDD.t157 VDD.n625 13.2328
R16543 VDD.t122 VDD.n328 13.2328
R16544 VDD.n291 VDD.n256 13.1884
R16545 VDD.n240 VDD.n205 13.1884
R16546 VDD.n197 VDD.n162 13.1884
R16547 VDD.n146 VDD.n111 13.1884
R16548 VDD.n104 VDD.n69 13.1884
R16549 VDD.n53 VDD.n18 13.1884
R16550 VDD.n1780 VDD.n1745 13.1884
R16551 VDD.n1831 VDD.n1796 13.1884
R16552 VDD.n1686 VDD.n1651 13.1884
R16553 VDD.n1737 VDD.n1702 13.1884
R16554 VDD.n1593 VDD.n1558 13.1884
R16555 VDD.n1644 VDD.n1609 13.1884
R16556 VDD.n1355 VDD.n1286 12.9944
R16557 VDD.n1355 VDD.n1354 12.9944
R16558 VDD.n2078 VDD.n1951 12.9944
R16559 VDD.n2079 VDD.n2078 12.9944
R16560 VDD.n483 VDD.n420 12.9944
R16561 VDD.n477 VDD.n420 12.9944
R16562 VDD.n3177 VDD.n712 12.9944
R16563 VDD.n3180 VDD.n3177 12.9944
R16564 VDD.n292 VDD.n254 12.8005
R16565 VDD.n287 VDD.n258 12.8005
R16566 VDD.n241 VDD.n203 12.8005
R16567 VDD.n236 VDD.n207 12.8005
R16568 VDD.n198 VDD.n160 12.8005
R16569 VDD.n193 VDD.n164 12.8005
R16570 VDD.n147 VDD.n109 12.8005
R16571 VDD.n142 VDD.n113 12.8005
R16572 VDD.n105 VDD.n67 12.8005
R16573 VDD.n100 VDD.n71 12.8005
R16574 VDD.n54 VDD.n16 12.8005
R16575 VDD.n49 VDD.n20 12.8005
R16576 VDD.n1781 VDD.n1743 12.8005
R16577 VDD.n1776 VDD.n1747 12.8005
R16578 VDD.n1832 VDD.n1794 12.8005
R16579 VDD.n1827 VDD.n1798 12.8005
R16580 VDD.n1687 VDD.n1649 12.8005
R16581 VDD.n1682 VDD.n1653 12.8005
R16582 VDD.n1738 VDD.n1700 12.8005
R16583 VDD.n1733 VDD.n1704 12.8005
R16584 VDD.n1594 VDD.n1556 12.8005
R16585 VDD.n1589 VDD.n1560 12.8005
R16586 VDD.n1645 VDD.n1607 12.8005
R16587 VDD.n1640 VDD.n1611 12.8005
R16588 VDD.n286 VDD.n259 12.0247
R16589 VDD.n235 VDD.n208 12.0247
R16590 VDD.n192 VDD.n165 12.0247
R16591 VDD.n141 VDD.n114 12.0247
R16592 VDD.n99 VDD.n72 12.0247
R16593 VDD.n48 VDD.n21 12.0247
R16594 VDD.n1775 VDD.n1748 12.0247
R16595 VDD.n1826 VDD.n1799 12.0247
R16596 VDD.n1681 VDD.n1654 12.0247
R16597 VDD.n1732 VDD.n1705 12.0247
R16598 VDD.n1588 VDD.n1561 12.0247
R16599 VDD.n1639 VDD.n1612 12.0247
R16600 VDD.n283 VDD.n282 11.249
R16601 VDD.n232 VDD.n231 11.249
R16602 VDD.n189 VDD.n188 11.249
R16603 VDD.n138 VDD.n137 11.249
R16604 VDD.n96 VDD.n95 11.249
R16605 VDD.n45 VDD.n44 11.249
R16606 VDD.n1772 VDD.n1771 11.249
R16607 VDD.n1823 VDD.n1822 11.249
R16608 VDD.n1678 VDD.n1677 11.249
R16609 VDD.n1729 VDD.n1728 11.249
R16610 VDD.n1585 VDD.n1584 11.249
R16611 VDD.n1636 VDD.n1635 11.249
R16612 VDD.n268 VDD.n267 10.7238
R16613 VDD.n217 VDD.n216 10.7238
R16614 VDD.n174 VDD.n173 10.7238
R16615 VDD.n123 VDD.n122 10.7238
R16616 VDD.n81 VDD.n80 10.7238
R16617 VDD.n30 VDD.n29 10.7238
R16618 VDD.n1757 VDD.n1756 10.7238
R16619 VDD.n1808 VDD.n1807 10.7238
R16620 VDD.n1663 VDD.n1662 10.7238
R16621 VDD.n1714 VDD.n1713 10.7238
R16622 VDD.n1570 VDD.n1569 10.7238
R16623 VDD.n1621 VDD.n1620 10.7238
R16624 VDD.n2532 VDD.n2530 10.6151
R16625 VDD.n2530 VDD.n2527 10.6151
R16626 VDD.n2527 VDD.n2526 10.6151
R16627 VDD.n2526 VDD.n2523 10.6151
R16628 VDD.n2523 VDD.n2522 10.6151
R16629 VDD.n2522 VDD.n2519 10.6151
R16630 VDD.n2519 VDD.n2518 10.6151
R16631 VDD.n2518 VDD.n2515 10.6151
R16632 VDD.n2515 VDD.n2514 10.6151
R16633 VDD.n2514 VDD.n2511 10.6151
R16634 VDD.n2511 VDD.n2510 10.6151
R16635 VDD.n2510 VDD.n2507 10.6151
R16636 VDD.n2507 VDD.n2506 10.6151
R16637 VDD.n2506 VDD.n2503 10.6151
R16638 VDD.n2503 VDD.n2502 10.6151
R16639 VDD.n2502 VDD.n2499 10.6151
R16640 VDD.n2499 VDD.n2498 10.6151
R16641 VDD.n2498 VDD.n2495 10.6151
R16642 VDD.n2495 VDD.n2494 10.6151
R16643 VDD.n2494 VDD.n2491 10.6151
R16644 VDD.n2491 VDD.n2490 10.6151
R16645 VDD.n2490 VDD.n2487 10.6151
R16646 VDD.n2485 VDD.n2482 10.6151
R16647 VDD.n2482 VDD.n2481 10.6151
R16648 VDD.n2303 VDD.n2302 10.6151
R16649 VDD.n2302 VDD.n2300 10.6151
R16650 VDD.n2300 VDD.n2299 10.6151
R16651 VDD.n2299 VDD.n2297 10.6151
R16652 VDD.n2297 VDD.n2296 10.6151
R16653 VDD.n2296 VDD.n2294 10.6151
R16654 VDD.n2294 VDD.n2293 10.6151
R16655 VDD.n2293 VDD.n2291 10.6151
R16656 VDD.n2291 VDD.n2290 10.6151
R16657 VDD.n2290 VDD.n2288 10.6151
R16658 VDD.n2288 VDD.n2287 10.6151
R16659 VDD.n2287 VDD.n2285 10.6151
R16660 VDD.n2285 VDD.n2284 10.6151
R16661 VDD.n2284 VDD.n2282 10.6151
R16662 VDD.n2282 VDD.n2281 10.6151
R16663 VDD.n2281 VDD.n2279 10.6151
R16664 VDD.n2279 VDD.n2278 10.6151
R16665 VDD.n2278 VDD.n2276 10.6151
R16666 VDD.n2276 VDD.n2275 10.6151
R16667 VDD.n2275 VDD.n2273 10.6151
R16668 VDD.n2273 VDD.n2272 10.6151
R16669 VDD.n2272 VDD.n1079 10.6151
R16670 VDD.n2241 VDD.n1079 10.6151
R16671 VDD.n2242 VDD.n2241 10.6151
R16672 VDD.n2259 VDD.n2242 10.6151
R16673 VDD.n2259 VDD.n2258 10.6151
R16674 VDD.n2258 VDD.n2257 10.6151
R16675 VDD.n2257 VDD.n2255 10.6151
R16676 VDD.n2255 VDD.n2254 10.6151
R16677 VDD.n2254 VDD.n2252 10.6151
R16678 VDD.n2252 VDD.n2251 10.6151
R16679 VDD.n2251 VDD.n2249 10.6151
R16680 VDD.n2249 VDD.n2248 10.6151
R16681 VDD.n2248 VDD.n2246 10.6151
R16682 VDD.n2246 VDD.n2245 10.6151
R16683 VDD.n2245 VDD.n2243 10.6151
R16684 VDD.n2243 VDD.n945 10.6151
R16685 VDD.n2476 VDD.n945 10.6151
R16686 VDD.n2477 VDD.n2476 10.6151
R16687 VDD.n2478 VDD.n2477 10.6151
R16688 VDD.n2354 VDD.n2353 10.6151
R16689 VDD.n2353 VDD.n1063 10.6151
R16690 VDD.n2348 VDD.n1063 10.6151
R16691 VDD.n2348 VDD.n2347 10.6151
R16692 VDD.n2347 VDD.n1065 10.6151
R16693 VDD.n2342 VDD.n1065 10.6151
R16694 VDD.n2342 VDD.n2341 10.6151
R16695 VDD.n2341 VDD.n2340 10.6151
R16696 VDD.n2340 VDD.n1067 10.6151
R16697 VDD.n2334 VDD.n1067 10.6151
R16698 VDD.n2334 VDD.n2333 10.6151
R16699 VDD.n2333 VDD.n2332 10.6151
R16700 VDD.n2328 VDD.n2327 10.6151
R16701 VDD.n2327 VDD.n1071 10.6151
R16702 VDD.n2322 VDD.n1071 10.6151
R16703 VDD.n2322 VDD.n2321 10.6151
R16704 VDD.n2321 VDD.n2320 10.6151
R16705 VDD.n2320 VDD.n1073 10.6151
R16706 VDD.n2314 VDD.n1073 10.6151
R16707 VDD.n2314 VDD.n2313 10.6151
R16708 VDD.n2313 VDD.n2312 10.6151
R16709 VDD.n2308 VDD.n2307 10.6151
R16710 VDD.n2307 VDD.n2304 10.6151
R16711 VDD.n2355 VDD.n1050 10.6151
R16712 VDD.n2365 VDD.n1050 10.6151
R16713 VDD.n2366 VDD.n2365 10.6151
R16714 VDD.n2367 VDD.n2366 10.6151
R16715 VDD.n2367 VDD.n1038 10.6151
R16716 VDD.n2378 VDD.n1038 10.6151
R16717 VDD.n2379 VDD.n2378 10.6151
R16718 VDD.n2380 VDD.n2379 10.6151
R16719 VDD.n2380 VDD.n1026 10.6151
R16720 VDD.n2390 VDD.n1026 10.6151
R16721 VDD.n2391 VDD.n2390 10.6151
R16722 VDD.n2392 VDD.n2391 10.6151
R16723 VDD.n2392 VDD.n1014 10.6151
R16724 VDD.n2402 VDD.n1014 10.6151
R16725 VDD.n2403 VDD.n2402 10.6151
R16726 VDD.n2404 VDD.n2403 10.6151
R16727 VDD.n2404 VDD.n1002 10.6151
R16728 VDD.n2414 VDD.n1002 10.6151
R16729 VDD.n2415 VDD.n2414 10.6151
R16730 VDD.n2416 VDD.n2415 10.6151
R16731 VDD.n2416 VDD.n991 10.6151
R16732 VDD.n2426 VDD.n991 10.6151
R16733 VDD.n2427 VDD.n2426 10.6151
R16734 VDD.n2428 VDD.n2427 10.6151
R16735 VDD.n2428 VDD.n980 10.6151
R16736 VDD.n2438 VDD.n980 10.6151
R16737 VDD.n2439 VDD.n2438 10.6151
R16738 VDD.n2440 VDD.n2439 10.6151
R16739 VDD.n2440 VDD.n968 10.6151
R16740 VDD.n2450 VDD.n968 10.6151
R16741 VDD.n2451 VDD.n2450 10.6151
R16742 VDD.n2452 VDD.n2451 10.6151
R16743 VDD.n2452 VDD.n956 10.6151
R16744 VDD.n2462 VDD.n956 10.6151
R16745 VDD.n2463 VDD.n2462 10.6151
R16746 VDD.n2465 VDD.n2463 10.6151
R16747 VDD.n2465 VDD.n2464 10.6151
R16748 VDD.n2464 VDD.n942 10.6151
R16749 VDD.n2534 VDD.n942 10.6151
R16750 VDD.n2534 VDD.n2533 10.6151
R16751 VDD.n2679 VDD.n2677 10.6151
R16752 VDD.n2680 VDD.n2679 10.6151
R16753 VDD.n2682 VDD.n2680 10.6151
R16754 VDD.n2683 VDD.n2682 10.6151
R16755 VDD.n2685 VDD.n2683 10.6151
R16756 VDD.n2686 VDD.n2685 10.6151
R16757 VDD.n2688 VDD.n2686 10.6151
R16758 VDD.n2689 VDD.n2688 10.6151
R16759 VDD.n2691 VDD.n2689 10.6151
R16760 VDD.n2692 VDD.n2691 10.6151
R16761 VDD.n2694 VDD.n2692 10.6151
R16762 VDD.n2695 VDD.n2694 10.6151
R16763 VDD.n2697 VDD.n2695 10.6151
R16764 VDD.n2698 VDD.n2697 10.6151
R16765 VDD.n2766 VDD.n2698 10.6151
R16766 VDD.n2766 VDD.n2765 10.6151
R16767 VDD.n2765 VDD.n2764 10.6151
R16768 VDD.n2764 VDD.n2762 10.6151
R16769 VDD.n2762 VDD.n2761 10.6151
R16770 VDD.n2761 VDD.n2724 10.6151
R16771 VDD.n2724 VDD.n2723 10.6151
R16772 VDD.n2723 VDD.n2721 10.6151
R16773 VDD.n2721 VDD.n2720 10.6151
R16774 VDD.n2720 VDD.n2718 10.6151
R16775 VDD.n2718 VDD.n2717 10.6151
R16776 VDD.n2717 VDD.n2715 10.6151
R16777 VDD.n2715 VDD.n2714 10.6151
R16778 VDD.n2714 VDD.n2712 10.6151
R16779 VDD.n2712 VDD.n2711 10.6151
R16780 VDD.n2711 VDD.n2709 10.6151
R16781 VDD.n2709 VDD.n2708 10.6151
R16782 VDD.n2708 VDD.n2706 10.6151
R16783 VDD.n2706 VDD.n2705 10.6151
R16784 VDD.n2705 VDD.n2703 10.6151
R16785 VDD.n2703 VDD.n2702 10.6151
R16786 VDD.n2702 VDD.n2700 10.6151
R16787 VDD.n2700 VDD.n2699 10.6151
R16788 VDD.n2699 VDD.n788 10.6151
R16789 VDD.n3001 VDD.n788 10.6151
R16790 VDD.n3002 VDD.n3001 10.6151
R16791 VDD.n2628 VDD.n901 10.6151
R16792 VDD.n2629 VDD.n2628 10.6151
R16793 VDD.n2630 VDD.n2629 10.6151
R16794 VDD.n2630 VDD.n2624 10.6151
R16795 VDD.n2636 VDD.n2624 10.6151
R16796 VDD.n2637 VDD.n2636 10.6151
R16797 VDD.n2638 VDD.n2637 10.6151
R16798 VDD.n2638 VDD.n2622 10.6151
R16799 VDD.n2644 VDD.n2622 10.6151
R16800 VDD.n2645 VDD.n2644 10.6151
R16801 VDD.n2646 VDD.n2645 10.6151
R16802 VDD.n2646 VDD.n2620 10.6151
R16803 VDD.n2652 VDD.n2620 10.6151
R16804 VDD.n2653 VDD.n2652 10.6151
R16805 VDD.n2654 VDD.n2653 10.6151
R16806 VDD.n2654 VDD.n2618 10.6151
R16807 VDD.n2660 VDD.n2618 10.6151
R16808 VDD.n2661 VDD.n2660 10.6151
R16809 VDD.n2662 VDD.n2661 10.6151
R16810 VDD.n2662 VDD.n2616 10.6151
R16811 VDD.n2668 VDD.n2616 10.6151
R16812 VDD.n2669 VDD.n2668 10.6151
R16813 VDD.n2671 VDD.n2612 10.6151
R16814 VDD.n2676 VDD.n2612 10.6151
R16815 VDD.n2850 VDD.n2849 10.6151
R16816 VDD.n2851 VDD.n2850 10.6151
R16817 VDD.n2851 VDD.n889 10.6151
R16818 VDD.n2861 VDD.n889 10.6151
R16819 VDD.n2862 VDD.n2861 10.6151
R16820 VDD.n2863 VDD.n2862 10.6151
R16821 VDD.n2863 VDD.n877 10.6151
R16822 VDD.n2873 VDD.n877 10.6151
R16823 VDD.n2874 VDD.n2873 10.6151
R16824 VDD.n2875 VDD.n2874 10.6151
R16825 VDD.n2875 VDD.n866 10.6151
R16826 VDD.n2885 VDD.n866 10.6151
R16827 VDD.n2886 VDD.n2885 10.6151
R16828 VDD.n2887 VDD.n2886 10.6151
R16829 VDD.n2887 VDD.n855 10.6151
R16830 VDD.n2897 VDD.n855 10.6151
R16831 VDD.n2898 VDD.n2897 10.6151
R16832 VDD.n2899 VDD.n2898 10.6151
R16833 VDD.n2899 VDD.n843 10.6151
R16834 VDD.n2909 VDD.n843 10.6151
R16835 VDD.n2910 VDD.n2909 10.6151
R16836 VDD.n2911 VDD.n2910 10.6151
R16837 VDD.n2911 VDD.n831 10.6151
R16838 VDD.n2921 VDD.n831 10.6151
R16839 VDD.n2922 VDD.n2921 10.6151
R16840 VDD.n2923 VDD.n2922 10.6151
R16841 VDD.n2923 VDD.n819 10.6151
R16842 VDD.n2933 VDD.n819 10.6151
R16843 VDD.n2934 VDD.n2933 10.6151
R16844 VDD.n2935 VDD.n2934 10.6151
R16845 VDD.n2935 VDD.n808 10.6151
R16846 VDD.n2945 VDD.n808 10.6151
R16847 VDD.n2946 VDD.n2945 10.6151
R16848 VDD.n2947 VDD.n2946 10.6151
R16849 VDD.n2947 VDD.n794 10.6151
R16850 VDD.n2994 VDD.n794 10.6151
R16851 VDD.n2995 VDD.n2994 10.6151
R16852 VDD.n2996 VDD.n2995 10.6151
R16853 VDD.n2996 VDD.n766 10.6151
R16854 VDD.n3051 VDD.n766 10.6151
R16855 VDD.n3050 VDD.n3049 10.6151
R16856 VDD.n3049 VDD.n767 10.6151
R16857 VDD.n3044 VDD.n767 10.6151
R16858 VDD.n3044 VDD.n3043 10.6151
R16859 VDD.n3043 VDD.n3042 10.6151
R16860 VDD.n3042 VDD.n770 10.6151
R16861 VDD.n3037 VDD.n770 10.6151
R16862 VDD.n3037 VDD.n3036 10.6151
R16863 VDD.n3036 VDD.n3035 10.6151
R16864 VDD.n3035 VDD.n773 10.6151
R16865 VDD.n3030 VDD.n773 10.6151
R16866 VDD.n3030 VDD.n3029 10.6151
R16867 VDD.n3026 VDD.n776 10.6151
R16868 VDD.n3021 VDD.n776 10.6151
R16869 VDD.n3021 VDD.n3020 10.6151
R16870 VDD.n3020 VDD.n3019 10.6151
R16871 VDD.n3019 VDD.n779 10.6151
R16872 VDD.n3014 VDD.n779 10.6151
R16873 VDD.n3014 VDD.n3013 10.6151
R16874 VDD.n3013 VDD.n3012 10.6151
R16875 VDD.n3012 VDD.n782 10.6151
R16876 VDD.n3007 VDD.n3006 10.6151
R16877 VDD.n3006 VDD.n3005 10.6151
R16878 VDD.n2984 VDD.n2954 10.6151
R16879 VDD.n2955 VDD.n2954 10.6151
R16880 VDD.n2977 VDD.n2955 10.6151
R16881 VDD.n2977 VDD.n2976 10.6151
R16882 VDD.n2976 VDD.n2975 10.6151
R16883 VDD.n2975 VDD.n2957 10.6151
R16884 VDD.n2970 VDD.n2957 10.6151
R16885 VDD.n2970 VDD.n2969 10.6151
R16886 VDD.n2969 VDD.n2968 10.6151
R16887 VDD.n2968 VDD.n2960 10.6151
R16888 VDD.n2963 VDD.n2960 10.6151
R16889 VDD.n2963 VDD.n745 10.6151
R16890 VDD.n3077 VDD.n746 10.6151
R16891 VDD.n3072 VDD.n746 10.6151
R16892 VDD.n3072 VDD.n3071 10.6151
R16893 VDD.n3071 VDD.n3070 10.6151
R16894 VDD.n3070 VDD.n749 10.6151
R16895 VDD.n3065 VDD.n749 10.6151
R16896 VDD.n3065 VDD.n3064 10.6151
R16897 VDD.n3064 VDD.n3063 10.6151
R16898 VDD.n3063 VDD.n752 10.6151
R16899 VDD.n3058 VDD.n3057 10.6151
R16900 VDD.n3057 VDD.n3056 10.6151
R16901 VDD.n2792 VDD.n2791 10.6151
R16902 VDD.n2791 VDD.n2789 10.6151
R16903 VDD.n2789 VDD.n2788 10.6151
R16904 VDD.n2788 VDD.n2786 10.6151
R16905 VDD.n2786 VDD.n2785 10.6151
R16906 VDD.n2785 VDD.n2783 10.6151
R16907 VDD.n2783 VDD.n2782 10.6151
R16908 VDD.n2782 VDD.n2780 10.6151
R16909 VDD.n2780 VDD.n2779 10.6151
R16910 VDD.n2779 VDD.n2777 10.6151
R16911 VDD.n2777 VDD.n2776 10.6151
R16912 VDD.n2776 VDD.n2774 10.6151
R16913 VDD.n2774 VDD.n2773 10.6151
R16914 VDD.n2773 VDD.n2771 10.6151
R16915 VDD.n2771 VDD.n2770 10.6151
R16916 VDD.n2770 VDD.n2611 10.6151
R16917 VDD.n2726 VDD.n2611 10.6151
R16918 VDD.n2727 VDD.n2726 10.6151
R16919 VDD.n2757 VDD.n2727 10.6151
R16920 VDD.n2757 VDD.n2756 10.6151
R16921 VDD.n2756 VDD.n2755 10.6151
R16922 VDD.n2755 VDD.n2753 10.6151
R16923 VDD.n2753 VDD.n2752 10.6151
R16924 VDD.n2752 VDD.n2750 10.6151
R16925 VDD.n2750 VDD.n2749 10.6151
R16926 VDD.n2749 VDD.n2747 10.6151
R16927 VDD.n2747 VDD.n2746 10.6151
R16928 VDD.n2746 VDD.n2744 10.6151
R16929 VDD.n2744 VDD.n2743 10.6151
R16930 VDD.n2743 VDD.n2741 10.6151
R16931 VDD.n2741 VDD.n2740 10.6151
R16932 VDD.n2740 VDD.n2738 10.6151
R16933 VDD.n2738 VDD.n2737 10.6151
R16934 VDD.n2737 VDD.n2735 10.6151
R16935 VDD.n2735 VDD.n2734 10.6151
R16936 VDD.n2734 VDD.n2732 10.6151
R16937 VDD.n2732 VDD.n2731 10.6151
R16938 VDD.n2731 VDD.n2729 10.6151
R16939 VDD.n2729 VDD.n2728 10.6151
R16940 VDD.n2728 VDD.n758 10.6151
R16941 VDD.n2844 VDD.n2843 10.6151
R16942 VDD.n2843 VDD.n2596 10.6151
R16943 VDD.n2837 VDD.n2596 10.6151
R16944 VDD.n2837 VDD.n2836 10.6151
R16945 VDD.n2836 VDD.n2835 10.6151
R16946 VDD.n2835 VDD.n2598 10.6151
R16947 VDD.n2829 VDD.n2598 10.6151
R16948 VDD.n2829 VDD.n2828 10.6151
R16949 VDD.n2828 VDD.n2827 10.6151
R16950 VDD.n2827 VDD.n2600 10.6151
R16951 VDD.n2821 VDD.n2600 10.6151
R16952 VDD.n2821 VDD.n2820 10.6151
R16953 VDD.n2820 VDD.n2819 10.6151
R16954 VDD.n2819 VDD.n2602 10.6151
R16955 VDD.n2813 VDD.n2602 10.6151
R16956 VDD.n2813 VDD.n2812 10.6151
R16957 VDD.n2812 VDD.n2811 10.6151
R16958 VDD.n2811 VDD.n2604 10.6151
R16959 VDD.n2805 VDD.n2604 10.6151
R16960 VDD.n2805 VDD.n2804 10.6151
R16961 VDD.n2804 VDD.n2803 10.6151
R16962 VDD.n2803 VDD.n2606 10.6151
R16963 VDD.n2797 VDD.n2796 10.6151
R16964 VDD.n2796 VDD.n2795 10.6151
R16965 VDD.n2845 VDD.n895 10.6151
R16966 VDD.n2855 VDD.n895 10.6151
R16967 VDD.n2856 VDD.n2855 10.6151
R16968 VDD.n2857 VDD.n2856 10.6151
R16969 VDD.n2857 VDD.n884 10.6151
R16970 VDD.n2867 VDD.n884 10.6151
R16971 VDD.n2868 VDD.n2867 10.6151
R16972 VDD.n2869 VDD.n2868 10.6151
R16973 VDD.n2869 VDD.n872 10.6151
R16974 VDD.n2879 VDD.n872 10.6151
R16975 VDD.n2880 VDD.n2879 10.6151
R16976 VDD.n2881 VDD.n2880 10.6151
R16977 VDD.n2881 VDD.n860 10.6151
R16978 VDD.n2891 VDD.n860 10.6151
R16979 VDD.n2892 VDD.n2891 10.6151
R16980 VDD.n2893 VDD.n2892 10.6151
R16981 VDD.n2893 VDD.n849 10.6151
R16982 VDD.n2903 VDD.n849 10.6151
R16983 VDD.n2904 VDD.n2903 10.6151
R16984 VDD.n2905 VDD.n2904 10.6151
R16985 VDD.n2905 VDD.n837 10.6151
R16986 VDD.n2915 VDD.n837 10.6151
R16987 VDD.n2916 VDD.n2915 10.6151
R16988 VDD.n2917 VDD.n2916 10.6151
R16989 VDD.n2917 VDD.n825 10.6151
R16990 VDD.n2927 VDD.n825 10.6151
R16991 VDD.n2928 VDD.n2927 10.6151
R16992 VDD.n2929 VDD.n2928 10.6151
R16993 VDD.n2929 VDD.n814 10.6151
R16994 VDD.n2939 VDD.n814 10.6151
R16995 VDD.n2940 VDD.n2939 10.6151
R16996 VDD.n2941 VDD.n2940 10.6151
R16997 VDD.n2941 VDD.n802 10.6151
R16998 VDD.n2951 VDD.n802 10.6151
R16999 VDD.n2990 VDD.n2953 10.6151
R17000 VDD.n2990 VDD.n2989 10.6151
R17001 VDD.n2989 VDD.n2988 10.6151
R17002 VDD.n2988 VDD.n2987 10.6151
R17003 VDD.n2987 VDD.n2985 10.6151
R17004 VDD.n2360 VDD.n2359 10.6151
R17005 VDD.n2361 VDD.n2360 10.6151
R17006 VDD.n2361 VDD.n1044 10.6151
R17007 VDD.n2371 VDD.n1044 10.6151
R17008 VDD.n2372 VDD.n2371 10.6151
R17009 VDD.n2374 VDD.n1032 10.6151
R17010 VDD.n2384 VDD.n1032 10.6151
R17011 VDD.n2385 VDD.n2384 10.6151
R17012 VDD.n2386 VDD.n2385 10.6151
R17013 VDD.n2386 VDD.n1020 10.6151
R17014 VDD.n2396 VDD.n1020 10.6151
R17015 VDD.n2397 VDD.n2396 10.6151
R17016 VDD.n2398 VDD.n2397 10.6151
R17017 VDD.n2398 VDD.n1008 10.6151
R17018 VDD.n2408 VDD.n1008 10.6151
R17019 VDD.n2409 VDD.n2408 10.6151
R17020 VDD.n2410 VDD.n2409 10.6151
R17021 VDD.n2410 VDD.n996 10.6151
R17022 VDD.n2420 VDD.n996 10.6151
R17023 VDD.n2421 VDD.n2420 10.6151
R17024 VDD.n2422 VDD.n2421 10.6151
R17025 VDD.n2422 VDD.n985 10.6151
R17026 VDD.n2432 VDD.n985 10.6151
R17027 VDD.n2433 VDD.n2432 10.6151
R17028 VDD.n2434 VDD.n2433 10.6151
R17029 VDD.n2434 VDD.n973 10.6151
R17030 VDD.n2444 VDD.n973 10.6151
R17031 VDD.n2445 VDD.n2444 10.6151
R17032 VDD.n2446 VDD.n2445 10.6151
R17033 VDD.n2446 VDD.n962 10.6151
R17034 VDD.n2456 VDD.n962 10.6151
R17035 VDD.n2457 VDD.n2456 10.6151
R17036 VDD.n2458 VDD.n2457 10.6151
R17037 VDD.n2458 VDD.n949 10.6151
R17038 VDD.n2469 VDD.n949 10.6151
R17039 VDD.n2470 VDD.n2469 10.6151
R17040 VDD.n2472 VDD.n2470 10.6151
R17041 VDD.n2472 VDD.n2471 10.6151
R17042 VDD.n2471 VDD.n932 10.6151
R17043 VDD.n2588 VDD.n2587 10.6151
R17044 VDD.n2587 VDD.n2586 10.6151
R17045 VDD.n2586 VDD.n2583 10.6151
R17046 VDD.n2583 VDD.n2582 10.6151
R17047 VDD.n2582 VDD.n2579 10.6151
R17048 VDD.n2579 VDD.n2578 10.6151
R17049 VDD.n2578 VDD.n2575 10.6151
R17050 VDD.n2575 VDD.n2574 10.6151
R17051 VDD.n2574 VDD.n2571 10.6151
R17052 VDD.n2571 VDD.n2570 10.6151
R17053 VDD.n2570 VDD.n2567 10.6151
R17054 VDD.n2567 VDD.n2566 10.6151
R17055 VDD.n2566 VDD.n2563 10.6151
R17056 VDD.n2563 VDD.n2562 10.6151
R17057 VDD.n2562 VDD.n2559 10.6151
R17058 VDD.n2559 VDD.n2558 10.6151
R17059 VDD.n2558 VDD.n2555 10.6151
R17060 VDD.n2555 VDD.n2554 10.6151
R17061 VDD.n2554 VDD.n2551 10.6151
R17062 VDD.n2551 VDD.n2550 10.6151
R17063 VDD.n2550 VDD.n2547 10.6151
R17064 VDD.n2547 VDD.n2546 10.6151
R17065 VDD.n2543 VDD.n2542 10.6151
R17066 VDD.n2542 VDD.n2540 10.6151
R17067 VDD.n2192 VDD.n2190 10.6151
R17068 VDD.n2193 VDD.n2192 10.6151
R17069 VDD.n2195 VDD.n2193 10.6151
R17070 VDD.n2196 VDD.n2195 10.6151
R17071 VDD.n2198 VDD.n2196 10.6151
R17072 VDD.n2199 VDD.n2198 10.6151
R17073 VDD.n2201 VDD.n2199 10.6151
R17074 VDD.n2202 VDD.n2201 10.6151
R17075 VDD.n2204 VDD.n2202 10.6151
R17076 VDD.n2205 VDD.n2204 10.6151
R17077 VDD.n2207 VDD.n2205 10.6151
R17078 VDD.n2208 VDD.n2207 10.6151
R17079 VDD.n2210 VDD.n2208 10.6151
R17080 VDD.n2211 VDD.n2210 10.6151
R17081 VDD.n2213 VDD.n2211 10.6151
R17082 VDD.n2214 VDD.n2213 10.6151
R17083 VDD.n2216 VDD.n2214 10.6151
R17084 VDD.n2217 VDD.n2216 10.6151
R17085 VDD.n2219 VDD.n2217 10.6151
R17086 VDD.n2220 VDD.n2219 10.6151
R17087 VDD.n2268 VDD.n2220 10.6151
R17088 VDD.n2268 VDD.n2267 10.6151
R17089 VDD.n2267 VDD.n2266 10.6151
R17090 VDD.n2266 VDD.n2264 10.6151
R17091 VDD.n2264 VDD.n2263 10.6151
R17092 VDD.n2263 VDD.n2239 10.6151
R17093 VDD.n2239 VDD.n2238 10.6151
R17094 VDD.n2238 VDD.n2236 10.6151
R17095 VDD.n2236 VDD.n2235 10.6151
R17096 VDD.n2235 VDD.n2233 10.6151
R17097 VDD.n2233 VDD.n2232 10.6151
R17098 VDD.n2232 VDD.n2230 10.6151
R17099 VDD.n2230 VDD.n2229 10.6151
R17100 VDD.n2229 VDD.n2227 10.6151
R17101 VDD.n2227 VDD.n2226 10.6151
R17102 VDD.n2226 VDD.n2224 10.6151
R17103 VDD.n2224 VDD.n2223 10.6151
R17104 VDD.n2223 VDD.n2221 10.6151
R17105 VDD.n2221 VDD.n936 10.6151
R17106 VDD.n2539 VDD.n936 10.6151
R17107 VDD.n2141 VDD.n1057 10.6151
R17108 VDD.n2142 VDD.n2141 10.6151
R17109 VDD.n2143 VDD.n2142 10.6151
R17110 VDD.n2143 VDD.n2137 10.6151
R17111 VDD.n2149 VDD.n2137 10.6151
R17112 VDD.n2150 VDD.n2149 10.6151
R17113 VDD.n2151 VDD.n2150 10.6151
R17114 VDD.n2151 VDD.n2135 10.6151
R17115 VDD.n2157 VDD.n2135 10.6151
R17116 VDD.n2158 VDD.n2157 10.6151
R17117 VDD.n2159 VDD.n2158 10.6151
R17118 VDD.n2159 VDD.n2133 10.6151
R17119 VDD.n2166 VDD.n2165 10.6151
R17120 VDD.n2167 VDD.n2166 10.6151
R17121 VDD.n2167 VDD.n1086 10.6151
R17122 VDD.n2173 VDD.n1086 10.6151
R17123 VDD.n2174 VDD.n2173 10.6151
R17124 VDD.n2175 VDD.n2174 10.6151
R17125 VDD.n2175 VDD.n1084 10.6151
R17126 VDD.n2181 VDD.n1084 10.6151
R17127 VDD.n2182 VDD.n2181 10.6151
R17128 VDD.n2184 VDD.n1080 10.6151
R17129 VDD.n2189 VDD.n1080 10.6151
R17130 VDD.n279 VDD.n261 10.4732
R17131 VDD.n228 VDD.n210 10.4732
R17132 VDD.n185 VDD.n167 10.4732
R17133 VDD.n134 VDD.n116 10.4732
R17134 VDD.n92 VDD.n74 10.4732
R17135 VDD.n41 VDD.n23 10.4732
R17136 VDD.n1768 VDD.n1750 10.4732
R17137 VDD.n1819 VDD.n1801 10.4732
R17138 VDD.n1674 VDD.n1656 10.4732
R17139 VDD.n1725 VDD.n1707 10.4732
R17140 VDD.n1581 VDD.n1563 10.4732
R17141 VDD.n1632 VDD.n1614 10.4732
R17142 VDD.n278 VDD.n263 9.69747
R17143 VDD.n227 VDD.n212 9.69747
R17144 VDD.n184 VDD.n169 9.69747
R17145 VDD.n133 VDD.n118 9.69747
R17146 VDD.n91 VDD.n76 9.69747
R17147 VDD.n40 VDD.n25 9.69747
R17148 VDD.n1767 VDD.n1752 9.69747
R17149 VDD.n1818 VDD.n1803 9.69747
R17150 VDD.n1673 VDD.n1658 9.69747
R17151 VDD.n1724 VDD.n1709 9.69747
R17152 VDD.n1580 VDD.n1565 9.69747
R17153 VDD.n1631 VDD.n1616 9.69747
R17154 VDD.n2094 VDD.n1069 9.61581
R17155 VDD.n3028 VDD.n3027 9.61581
R17156 VDD.n3079 VDD.n3078 9.61581
R17157 VDD.n2132 VDD.n2131 9.61581
R17158 VDD.n294 VDD.n293 9.45567
R17159 VDD.n243 VDD.n242 9.45567
R17160 VDD.n200 VDD.n199 9.45567
R17161 VDD.n149 VDD.n148 9.45567
R17162 VDD.n107 VDD.n106 9.45567
R17163 VDD.n56 VDD.n55 9.45567
R17164 VDD.n1783 VDD.n1782 9.45567
R17165 VDD.n1834 VDD.n1833 9.45567
R17166 VDD.n1689 VDD.n1688 9.45567
R17167 VDD.n1740 VDD.n1739 9.45567
R17168 VDD.n1596 VDD.n1595 9.45567
R17169 VDD.n1647 VDD.n1646 9.45567
R17170 VDD.n1209 VDD.t115 9.41319
R17171 VDD.t124 VDD.n1145 9.41319
R17172 VDD.n3265 VDD.t108 9.41319
R17173 VDD.t95 VDD.n3371 9.41319
R17174 VDD.n1840 VDD.n1839 9.3005
R17175 VDD.n1167 VDD.n1166 9.3005
R17176 VDD.n1853 VDD.n1852 9.3005
R17177 VDD.n1854 VDD.n1165 9.3005
R17178 VDD.n1856 VDD.n1855 9.3005
R17179 VDD.n1155 VDD.n1154 9.3005
R17180 VDD.n1869 VDD.n1868 9.3005
R17181 VDD.n1870 VDD.n1153 9.3005
R17182 VDD.n1872 VDD.n1871 9.3005
R17183 VDD.n1143 VDD.n1142 9.3005
R17184 VDD.n1885 VDD.n1884 9.3005
R17185 VDD.n1886 VDD.n1141 9.3005
R17186 VDD.n1888 VDD.n1887 9.3005
R17187 VDD.n1131 VDD.n1130 9.3005
R17188 VDD.n1901 VDD.n1900 9.3005
R17189 VDD.n1902 VDD.n1129 9.3005
R17190 VDD.n1904 VDD.n1903 9.3005
R17191 VDD.n1118 VDD.n1117 9.3005
R17192 VDD.n1918 VDD.n1917 9.3005
R17193 VDD.n1919 VDD.n1116 9.3005
R17194 VDD.n2113 VDD.n2112 9.3005
R17195 VDD.n2076 VDD.n1951 9.3005
R17196 VDD.n2075 VDD.n2074 9.3005
R17197 VDD.n1957 VDD.n1956 9.3005
R17198 VDD.n2069 VDD.n1961 9.3005
R17199 VDD.n2068 VDD.n1962 9.3005
R17200 VDD.n2067 VDD.n1963 9.3005
R17201 VDD.n1967 VDD.n1964 9.3005
R17202 VDD.n2062 VDD.n1968 9.3005
R17203 VDD.n2061 VDD.n1969 9.3005
R17204 VDD.n2060 VDD.n1970 9.3005
R17205 VDD.n1974 VDD.n1971 9.3005
R17206 VDD.n2055 VDD.n1975 9.3005
R17207 VDD.n2054 VDD.n1976 9.3005
R17208 VDD.n2053 VDD.n1977 9.3005
R17209 VDD.n1981 VDD.n1978 9.3005
R17210 VDD.n2048 VDD.n1982 9.3005
R17211 VDD.n2047 VDD.n1983 9.3005
R17212 VDD.n2046 VDD.n1984 9.3005
R17213 VDD.n1988 VDD.n1985 9.3005
R17214 VDD.n2041 VDD.n1989 9.3005
R17215 VDD.n2040 VDD.n1990 9.3005
R17216 VDD.n2039 VDD.n2038 9.3005
R17217 VDD.n2037 VDD.n1991 9.3005
R17218 VDD.n2036 VDD.n2035 9.3005
R17219 VDD.n1997 VDD.n1996 9.3005
R17220 VDD.n2030 VDD.n2001 9.3005
R17221 VDD.n2029 VDD.n2002 9.3005
R17222 VDD.n2028 VDD.n2003 9.3005
R17223 VDD.n2007 VDD.n2004 9.3005
R17224 VDD.n2023 VDD.n2008 9.3005
R17225 VDD.n2022 VDD.n2009 9.3005
R17226 VDD.n2021 VDD.n1088 9.3005
R17227 VDD.n2078 VDD.n2077 9.3005
R17228 VDD.n2109 VDD.n1920 9.3005
R17229 VDD.n1924 VDD.n1921 9.3005
R17230 VDD.n2104 VDD.n1925 9.3005
R17231 VDD.n2103 VDD.n1926 9.3005
R17232 VDD.n2102 VDD.n1927 9.3005
R17233 VDD.n1931 VDD.n1928 9.3005
R17234 VDD.n2097 VDD.n1932 9.3005
R17235 VDD.n1936 VDD.n1934 9.3005
R17236 VDD.n2087 VDD.n1942 9.3005
R17237 VDD.n2086 VDD.n1943 9.3005
R17238 VDD.n2085 VDD.n1944 9.3005
R17239 VDD.n1948 VDD.n1945 9.3005
R17240 VDD.n2080 VDD.n1949 9.3005
R17241 VDD.n2079 VDD.n1950 9.3005
R17242 VDD.n2111 VDD.n2110 9.3005
R17243 VDD.n270 VDD.n269 9.3005
R17244 VDD.n265 VDD.n264 9.3005
R17245 VDD.n276 VDD.n275 9.3005
R17246 VDD.n278 VDD.n277 9.3005
R17247 VDD.n261 VDD.n260 9.3005
R17248 VDD.n284 VDD.n283 9.3005
R17249 VDD.n286 VDD.n285 9.3005
R17250 VDD.n258 VDD.n255 9.3005
R17251 VDD.n293 VDD.n292 9.3005
R17252 VDD.n219 VDD.n218 9.3005
R17253 VDD.n214 VDD.n213 9.3005
R17254 VDD.n225 VDD.n224 9.3005
R17255 VDD.n227 VDD.n226 9.3005
R17256 VDD.n210 VDD.n209 9.3005
R17257 VDD.n233 VDD.n232 9.3005
R17258 VDD.n235 VDD.n234 9.3005
R17259 VDD.n207 VDD.n204 9.3005
R17260 VDD.n242 VDD.n241 9.3005
R17261 VDD.n176 VDD.n175 9.3005
R17262 VDD.n171 VDD.n170 9.3005
R17263 VDD.n182 VDD.n181 9.3005
R17264 VDD.n184 VDD.n183 9.3005
R17265 VDD.n167 VDD.n166 9.3005
R17266 VDD.n190 VDD.n189 9.3005
R17267 VDD.n192 VDD.n191 9.3005
R17268 VDD.n164 VDD.n161 9.3005
R17269 VDD.n199 VDD.n198 9.3005
R17270 VDD.n125 VDD.n124 9.3005
R17271 VDD.n120 VDD.n119 9.3005
R17272 VDD.n131 VDD.n130 9.3005
R17273 VDD.n133 VDD.n132 9.3005
R17274 VDD.n116 VDD.n115 9.3005
R17275 VDD.n139 VDD.n138 9.3005
R17276 VDD.n141 VDD.n140 9.3005
R17277 VDD.n113 VDD.n110 9.3005
R17278 VDD.n148 VDD.n147 9.3005
R17279 VDD.n83 VDD.n82 9.3005
R17280 VDD.n78 VDD.n77 9.3005
R17281 VDD.n89 VDD.n88 9.3005
R17282 VDD.n91 VDD.n90 9.3005
R17283 VDD.n74 VDD.n73 9.3005
R17284 VDD.n97 VDD.n96 9.3005
R17285 VDD.n99 VDD.n98 9.3005
R17286 VDD.n71 VDD.n68 9.3005
R17287 VDD.n106 VDD.n105 9.3005
R17288 VDD.n32 VDD.n31 9.3005
R17289 VDD.n27 VDD.n26 9.3005
R17290 VDD.n38 VDD.n37 9.3005
R17291 VDD.n40 VDD.n39 9.3005
R17292 VDD.n23 VDD.n22 9.3005
R17293 VDD.n46 VDD.n45 9.3005
R17294 VDD.n48 VDD.n47 9.3005
R17295 VDD.n20 VDD.n17 9.3005
R17296 VDD.n55 VDD.n54 9.3005
R17297 VDD.n3129 VDD.n3128 9.3005
R17298 VDD.n3132 VDD.n731 9.3005
R17299 VDD.n3133 VDD.n730 9.3005
R17300 VDD.n3136 VDD.n729 9.3005
R17301 VDD.n3137 VDD.n728 9.3005
R17302 VDD.n3140 VDD.n727 9.3005
R17303 VDD.n3141 VDD.n726 9.3005
R17304 VDD.n3144 VDD.n725 9.3005
R17305 VDD.n3145 VDD.n724 9.3005
R17306 VDD.n3148 VDD.n723 9.3005
R17307 VDD.n3149 VDD.n722 9.3005
R17308 VDD.n3152 VDD.n721 9.3005
R17309 VDD.n3153 VDD.n720 9.3005
R17310 VDD.n3156 VDD.n719 9.3005
R17311 VDD.n3157 VDD.n718 9.3005
R17312 VDD.n3160 VDD.n717 9.3005
R17313 VDD.n3161 VDD.n716 9.3005
R17314 VDD.n3164 VDD.n715 9.3005
R17315 VDD.n3165 VDD.n714 9.3005
R17316 VDD.n3168 VDD.n713 9.3005
R17317 VDD.n3172 VDD.n3171 9.3005
R17318 VDD.n3173 VDD.n712 9.3005
R17319 VDD.n3177 VDD.n3174 9.3005
R17320 VDD.n3180 VDD.n711 9.3005
R17321 VDD.n3181 VDD.n710 9.3005
R17322 VDD.n3184 VDD.n709 9.3005
R17323 VDD.n3185 VDD.n708 9.3005
R17324 VDD.n3188 VDD.n707 9.3005
R17325 VDD.n3189 VDD.n706 9.3005
R17326 VDD.n3192 VDD.n705 9.3005
R17327 VDD.n3201 VDD.n702 9.3005
R17328 VDD.n3204 VDD.n701 9.3005
R17329 VDD.n3205 VDD.n700 9.3005
R17330 VDD.n3208 VDD.n699 9.3005
R17331 VDD.n3210 VDD.n698 9.3005
R17332 VDD.n3211 VDD.n697 9.3005
R17333 VDD.n3212 VDD.n696 9.3005
R17334 VDD.n3213 VDD.n695 9.3005
R17335 VDD.n652 VDD.n651 9.3005
R17336 VDD.n3227 VDD.n3226 9.3005
R17337 VDD.n3228 VDD.n650 9.3005
R17338 VDD.n3230 VDD.n3229 9.3005
R17339 VDD.n640 VDD.n639 9.3005
R17340 VDD.n3244 VDD.n3243 9.3005
R17341 VDD.n3245 VDD.n638 9.3005
R17342 VDD.n3247 VDD.n3246 9.3005
R17343 VDD.n629 VDD.n628 9.3005
R17344 VDD.n3260 VDD.n3259 9.3005
R17345 VDD.n3261 VDD.n627 9.3005
R17346 VDD.n3263 VDD.n3262 9.3005
R17347 VDD.n617 VDD.n616 9.3005
R17348 VDD.n3277 VDD.n3276 9.3005
R17349 VDD.n3278 VDD.n615 9.3005
R17350 VDD.n3280 VDD.n3279 9.3005
R17351 VDD.n606 VDD.n605 9.3005
R17352 VDD.n3296 VDD.n3295 9.3005
R17353 VDD.n3297 VDD.n604 9.3005
R17354 VDD.n3299 VDD.n3298 9.3005
R17355 VDD.n299 VDD.n297 9.3005
R17356 VDD.n3392 VDD.n3391 9.3005
R17357 VDD.n300 VDD.n298 9.3005
R17358 VDD.n3385 VDD.n309 9.3005
R17359 VDD.n3384 VDD.n310 9.3005
R17360 VDD.n3383 VDD.n311 9.3005
R17361 VDD.n318 VDD.n312 9.3005
R17362 VDD.n3377 VDD.n319 9.3005
R17363 VDD.n3376 VDD.n320 9.3005
R17364 VDD.n3375 VDD.n321 9.3005
R17365 VDD.n330 VDD.n322 9.3005
R17366 VDD.n3369 VDD.n331 9.3005
R17367 VDD.n3368 VDD.n332 9.3005
R17368 VDD.n3367 VDD.n333 9.3005
R17369 VDD.n340 VDD.n334 9.3005
R17370 VDD.n3361 VDD.n341 9.3005
R17371 VDD.n3360 VDD.n342 9.3005
R17372 VDD.n3359 VDD.n343 9.3005
R17373 VDD.n352 VDD.n344 9.3005
R17374 VDD.n3353 VDD.n353 9.3005
R17375 VDD.n3352 VDD.n354 9.3005
R17376 VDD.n3351 VDD.n355 9.3005
R17377 VDD.n430 VDD.n356 9.3005
R17378 VDD.n434 VDD.n429 9.3005
R17379 VDD.n438 VDD.n437 9.3005
R17380 VDD.n439 VDD.n428 9.3005
R17381 VDD.n443 VDD.n440 9.3005
R17382 VDD.n444 VDD.n427 9.3005
R17383 VDD.n448 VDD.n447 9.3005
R17384 VDD.n449 VDD.n426 9.3005
R17385 VDD.n453 VDD.n450 9.3005
R17386 VDD.n454 VDD.n425 9.3005
R17387 VDD.n458 VDD.n457 9.3005
R17388 VDD.n459 VDD.n424 9.3005
R17389 VDD.n463 VDD.n460 9.3005
R17390 VDD.n464 VDD.n423 9.3005
R17391 VDD.n468 VDD.n467 9.3005
R17392 VDD.n469 VDD.n422 9.3005
R17393 VDD.n473 VDD.n470 9.3005
R17394 VDD.n474 VDD.n421 9.3005
R17395 VDD.n478 VDD.n477 9.3005
R17396 VDD.n479 VDD.n420 9.3005
R17397 VDD.n483 VDD.n480 9.3005
R17398 VDD.n484 VDD.n417 9.3005
R17399 VDD.n488 VDD.n487 9.3005
R17400 VDD.n489 VDD.n416 9.3005
R17401 VDD.n493 VDD.n490 9.3005
R17402 VDD.n494 VDD.n415 9.3005
R17403 VDD.n498 VDD.n497 9.3005
R17404 VDD.n499 VDD.n414 9.3005
R17405 VDD.n503 VDD.n500 9.3005
R17406 VDD.n504 VDD.n413 9.3005
R17407 VDD.n508 VDD.n507 9.3005
R17408 VDD.n509 VDD.n412 9.3005
R17409 VDD.n513 VDD.n510 9.3005
R17410 VDD.n514 VDD.n411 9.3005
R17411 VDD.n518 VDD.n517 9.3005
R17412 VDD.n519 VDD.n410 9.3005
R17413 VDD.n523 VDD.n520 9.3005
R17414 VDD.n524 VDD.n409 9.3005
R17415 VDD.n528 VDD.n527 9.3005
R17416 VDD.n529 VDD.n408 9.3005
R17417 VDD.n533 VDD.n530 9.3005
R17418 VDD.n534 VDD.n405 9.3005
R17419 VDD.n538 VDD.n537 9.3005
R17420 VDD.n539 VDD.n404 9.3005
R17421 VDD.n543 VDD.n540 9.3005
R17422 VDD.n544 VDD.n403 9.3005
R17423 VDD.n548 VDD.n547 9.3005
R17424 VDD.n549 VDD.n402 9.3005
R17425 VDD.n553 VDD.n550 9.3005
R17426 VDD.n554 VDD.n401 9.3005
R17427 VDD.n558 VDD.n557 9.3005
R17428 VDD.n559 VDD.n400 9.3005
R17429 VDD.n563 VDD.n560 9.3005
R17430 VDD.n564 VDD.n399 9.3005
R17431 VDD.n568 VDD.n567 9.3005
R17432 VDD.n569 VDD.n398 9.3005
R17433 VDD.n573 VDD.n570 9.3005
R17434 VDD.n574 VDD.n397 9.3005
R17435 VDD.n578 VDD.n577 9.3005
R17436 VDD.n579 VDD.n396 9.3005
R17437 VDD.n583 VDD.n580 9.3005
R17438 VDD.n585 VDD.n395 9.3005
R17439 VDD.n587 VDD.n586 9.3005
R17440 VDD.n3344 VDD.n3343 9.3005
R17441 VDD.n433 VDD.n431 9.3005
R17442 VDD.n3222 VDD.n3221 9.3005
R17443 VDD.n646 VDD.n645 9.3005
R17444 VDD.n3235 VDD.n3234 9.3005
R17445 VDD.n3236 VDD.n644 9.3005
R17446 VDD.n3238 VDD.n3237 9.3005
R17447 VDD.n635 VDD.n634 9.3005
R17448 VDD.n3252 VDD.n3251 9.3005
R17449 VDD.n3253 VDD.n633 9.3005
R17450 VDD.n3255 VDD.n3254 9.3005
R17451 VDD.n623 VDD.n622 9.3005
R17452 VDD.n3268 VDD.n3267 9.3005
R17453 VDD.n3269 VDD.n621 9.3005
R17454 VDD.n3271 VDD.n3270 9.3005
R17455 VDD.n612 VDD.n611 9.3005
R17456 VDD.n3285 VDD.n3284 9.3005
R17457 VDD.n3286 VDD.n610 9.3005
R17458 VDD.n3291 VDD.n3287 9.3005
R17459 VDD.n3290 VDD.n3289 9.3005
R17460 VDD.n3288 VDD.n599 9.3005
R17461 VDD.n3304 VDD.n600 9.3005
R17462 VDD.n3305 VDD.n598 9.3005
R17463 VDD.n3307 VDD.n3306 9.3005
R17464 VDD.n3308 VDD.n597 9.3005
R17465 VDD.n3311 VDD.n3309 9.3005
R17466 VDD.n3312 VDD.n596 9.3005
R17467 VDD.n3314 VDD.n3313 9.3005
R17468 VDD.n3315 VDD.n595 9.3005
R17469 VDD.n3318 VDD.n3316 9.3005
R17470 VDD.n3319 VDD.n594 9.3005
R17471 VDD.n3321 VDD.n3320 9.3005
R17472 VDD.n3322 VDD.n593 9.3005
R17473 VDD.n3325 VDD.n3323 9.3005
R17474 VDD.n3326 VDD.n592 9.3005
R17475 VDD.n3328 VDD.n3327 9.3005
R17476 VDD.n3329 VDD.n591 9.3005
R17477 VDD.n3332 VDD.n3330 9.3005
R17478 VDD.n3333 VDD.n590 9.3005
R17479 VDD.n3335 VDD.n3334 9.3005
R17480 VDD.n3336 VDD.n589 9.3005
R17481 VDD.n3339 VDD.n3337 9.3005
R17482 VDD.n3340 VDD.n588 9.3005
R17483 VDD.n3342 VDD.n3341 9.3005
R17484 VDD.n3220 VDD.n656 9.3005
R17485 VDD.n3219 VDD.n3218 9.3005
R17486 VDD.n3086 VDD.n657 9.3005
R17487 VDD.n3087 VDD.n3085 9.3005
R17488 VDD.n3090 VDD.n3084 9.3005
R17489 VDD.n3091 VDD.n3083 9.3005
R17490 VDD.n3094 VDD.n3082 9.3005
R17491 VDD.n3095 VDD.n3081 9.3005
R17492 VDD.n3098 VDD.n3080 9.3005
R17493 VDD.n3107 VDD.n742 9.3005
R17494 VDD.n3110 VDD.n741 9.3005
R17495 VDD.n3111 VDD.n740 9.3005
R17496 VDD.n3114 VDD.n739 9.3005
R17497 VDD.n3115 VDD.n738 9.3005
R17498 VDD.n3118 VDD.n737 9.3005
R17499 VDD.n3119 VDD.n736 9.3005
R17500 VDD.n3122 VDD.n735 9.3005
R17501 VDD.n3126 VDD.n3125 9.3005
R17502 VDD.n3127 VDD.n732 9.3005
R17503 VDD.n2130 VDD.n2129 9.3005
R17504 VDD.n2128 VDD.n1091 9.3005
R17505 VDD.n2127 VDD.n2126 9.3005
R17506 VDD.n2125 VDD.n1096 9.3005
R17507 VDD.n2124 VDD.n2123 9.3005
R17508 VDD.n2122 VDD.n1097 9.3005
R17509 VDD.n2121 VDD.n2120 9.3005
R17510 VDD.n2119 VDD.n2118 9.3005
R17511 VDD.n1231 VDD.n1230 9.3005
R17512 VDD.n1481 VDD.n1480 9.3005
R17513 VDD.n1482 VDD.n1229 9.3005
R17514 VDD.n1484 VDD.n1483 9.3005
R17515 VDD.n1219 VDD.n1218 9.3005
R17516 VDD.n1497 VDD.n1496 9.3005
R17517 VDD.n1498 VDD.n1217 9.3005
R17518 VDD.n1500 VDD.n1499 9.3005
R17519 VDD.n1207 VDD.n1206 9.3005
R17520 VDD.n1514 VDD.n1513 9.3005
R17521 VDD.n1515 VDD.n1205 9.3005
R17522 VDD.n1517 VDD.n1516 9.3005
R17523 VDD.n1196 VDD.n1195 9.3005
R17524 VDD.n1530 VDD.n1529 9.3005
R17525 VDD.n1531 VDD.n1194 9.3005
R17526 VDD.n1533 VDD.n1532 9.3005
R17527 VDD.n1184 VDD.n1183 9.3005
R17528 VDD.n1547 VDD.n1546 9.3005
R17529 VDD.n1548 VDD.n1182 9.3005
R17530 VDD.n1550 VDD.n1549 9.3005
R17531 VDD.n1173 VDD.n1172 9.3005
R17532 VDD.n1845 VDD.n1844 9.3005
R17533 VDD.n1846 VDD.n1171 9.3005
R17534 VDD.n1848 VDD.n1847 9.3005
R17535 VDD.n1160 VDD.n1159 9.3005
R17536 VDD.n1861 VDD.n1860 9.3005
R17537 VDD.n1862 VDD.n1158 9.3005
R17538 VDD.n1864 VDD.n1863 9.3005
R17539 VDD.n1149 VDD.n1148 9.3005
R17540 VDD.n1877 VDD.n1876 9.3005
R17541 VDD.n1878 VDD.n1147 9.3005
R17542 VDD.n1880 VDD.n1879 9.3005
R17543 VDD.n1136 VDD.n1135 9.3005
R17544 VDD.n1893 VDD.n1892 9.3005
R17545 VDD.n1894 VDD.n1134 9.3005
R17546 VDD.n1896 VDD.n1895 9.3005
R17547 VDD.n1125 VDD.n1124 9.3005
R17548 VDD.n1909 VDD.n1908 9.3005
R17549 VDD.n1910 VDD.n1122 9.3005
R17550 VDD.n1913 VDD.n1912 9.3005
R17551 VDD.n1911 VDD.n1123 9.3005
R17552 VDD.n1107 VDD.n1104 9.3005
R17553 VDD.n1467 VDD.n1466 9.3005
R17554 VDD.n1462 VDD.n1239 9.3005
R17555 VDD.n1452 VDD.n1242 9.3005
R17556 VDD.n1453 VDD.n1243 9.3005
R17557 VDD.n1455 VDD.n1454 9.3005
R17558 VDD.n1451 VDD.n1245 9.3005
R17559 VDD.n1450 VDD.n1449 9.3005
R17560 VDD.n1247 VDD.n1246 9.3005
R17561 VDD.n1443 VDD.n1442 9.3005
R17562 VDD.n1441 VDD.n1249 9.3005
R17563 VDD.n1440 VDD.n1439 9.3005
R17564 VDD.n1251 VDD.n1250 9.3005
R17565 VDD.n1433 VDD.n1432 9.3005
R17566 VDD.n1431 VDD.n1253 9.3005
R17567 VDD.n1430 VDD.n1429 9.3005
R17568 VDD.n1255 VDD.n1254 9.3005
R17569 VDD.n1423 VDD.n1422 9.3005
R17570 VDD.n1421 VDD.n1257 9.3005
R17571 VDD.n1420 VDD.n1419 9.3005
R17572 VDD.n1259 VDD.n1258 9.3005
R17573 VDD.n1413 VDD.n1412 9.3005
R17574 VDD.n1411 VDD.n1261 9.3005
R17575 VDD.n1410 VDD.n1409 9.3005
R17576 VDD.n1408 VDD.n1262 9.3005
R17577 VDD.n1398 VDD.n1267 9.3005
R17578 VDD.n1399 VDD.n1268 9.3005
R17579 VDD.n1401 VDD.n1400 9.3005
R17580 VDD.n1397 VDD.n1270 9.3005
R17581 VDD.n1396 VDD.n1395 9.3005
R17582 VDD.n1272 VDD.n1271 9.3005
R17583 VDD.n1389 VDD.n1388 9.3005
R17584 VDD.n1387 VDD.n1274 9.3005
R17585 VDD.n1386 VDD.n1385 9.3005
R17586 VDD.n1276 VDD.n1275 9.3005
R17587 VDD.n1379 VDD.n1378 9.3005
R17588 VDD.n1377 VDD.n1278 9.3005
R17589 VDD.n1376 VDD.n1375 9.3005
R17590 VDD.n1280 VDD.n1279 9.3005
R17591 VDD.n1369 VDD.n1368 9.3005
R17592 VDD.n1367 VDD.n1282 9.3005
R17593 VDD.n1366 VDD.n1365 9.3005
R17594 VDD.n1284 VDD.n1283 9.3005
R17595 VDD.n1359 VDD.n1358 9.3005
R17596 VDD.n1357 VDD.n1286 9.3005
R17597 VDD.n1356 VDD.n1355 9.3005
R17598 VDD.n1354 VDD.n1287 9.3005
R17599 VDD.n1344 VDD.n1292 9.3005
R17600 VDD.n1345 VDD.n1293 9.3005
R17601 VDD.n1347 VDD.n1346 9.3005
R17602 VDD.n1343 VDD.n1295 9.3005
R17603 VDD.n1342 VDD.n1341 9.3005
R17604 VDD.n1297 VDD.n1296 9.3005
R17605 VDD.n1335 VDD.n1334 9.3005
R17606 VDD.n1333 VDD.n1299 9.3005
R17607 VDD.n1332 VDD.n1331 9.3005
R17608 VDD.n1301 VDD.n1300 9.3005
R17609 VDD.n1325 VDD.n1324 9.3005
R17610 VDD.n1323 VDD.n1303 9.3005
R17611 VDD.n1322 VDD.n1321 9.3005
R17612 VDD.n1305 VDD.n1304 9.3005
R17613 VDD.n1315 VDD.n1314 9.3005
R17614 VDD.n1313 VDD.n1307 9.3005
R17615 VDD.n1312 VDD.n1311 9.3005
R17616 VDD.n1308 VDD.n1235 9.3005
R17617 VDD.n1465 VDD.n1464 9.3005
R17618 VDD.n1474 VDD.n1234 9.3005
R17619 VDD.n1476 VDD.n1475 9.3005
R17620 VDD.n1225 VDD.n1224 9.3005
R17621 VDD.n1489 VDD.n1488 9.3005
R17622 VDD.n1490 VDD.n1223 9.3005
R17623 VDD.n1492 VDD.n1491 9.3005
R17624 VDD.n1213 VDD.n1212 9.3005
R17625 VDD.n1506 VDD.n1505 9.3005
R17626 VDD.n1507 VDD.n1211 9.3005
R17627 VDD.n1509 VDD.n1508 9.3005
R17628 VDD.n1202 VDD.n1201 9.3005
R17629 VDD.n1522 VDD.n1521 9.3005
R17630 VDD.n1523 VDD.n1200 9.3005
R17631 VDD.n1525 VDD.n1524 9.3005
R17632 VDD.n1190 VDD.n1189 9.3005
R17633 VDD.n1539 VDD.n1538 9.3005
R17634 VDD.n1540 VDD.n1188 9.3005
R17635 VDD.n1542 VDD.n1541 9.3005
R17636 VDD.n1179 VDD.n1178 9.3005
R17637 VDD.n1555 VDD.n1554 9.3005
R17638 VDD.n1473 VDD.n1472 9.3005
R17639 VDD.n1838 VDD.n1177 9.3005
R17640 VDD.n1759 VDD.n1758 9.3005
R17641 VDD.n1754 VDD.n1753 9.3005
R17642 VDD.n1765 VDD.n1764 9.3005
R17643 VDD.n1767 VDD.n1766 9.3005
R17644 VDD.n1750 VDD.n1749 9.3005
R17645 VDD.n1773 VDD.n1772 9.3005
R17646 VDD.n1775 VDD.n1774 9.3005
R17647 VDD.n1747 VDD.n1744 9.3005
R17648 VDD.n1782 VDD.n1781 9.3005
R17649 VDD.n1810 VDD.n1809 9.3005
R17650 VDD.n1805 VDD.n1804 9.3005
R17651 VDD.n1816 VDD.n1815 9.3005
R17652 VDD.n1818 VDD.n1817 9.3005
R17653 VDD.n1801 VDD.n1800 9.3005
R17654 VDD.n1824 VDD.n1823 9.3005
R17655 VDD.n1826 VDD.n1825 9.3005
R17656 VDD.n1798 VDD.n1795 9.3005
R17657 VDD.n1833 VDD.n1832 9.3005
R17658 VDD.n1665 VDD.n1664 9.3005
R17659 VDD.n1660 VDD.n1659 9.3005
R17660 VDD.n1671 VDD.n1670 9.3005
R17661 VDD.n1673 VDD.n1672 9.3005
R17662 VDD.n1656 VDD.n1655 9.3005
R17663 VDD.n1679 VDD.n1678 9.3005
R17664 VDD.n1681 VDD.n1680 9.3005
R17665 VDD.n1653 VDD.n1650 9.3005
R17666 VDD.n1688 VDD.n1687 9.3005
R17667 VDD.n1716 VDD.n1715 9.3005
R17668 VDD.n1711 VDD.n1710 9.3005
R17669 VDD.n1722 VDD.n1721 9.3005
R17670 VDD.n1724 VDD.n1723 9.3005
R17671 VDD.n1707 VDD.n1706 9.3005
R17672 VDD.n1730 VDD.n1729 9.3005
R17673 VDD.n1732 VDD.n1731 9.3005
R17674 VDD.n1704 VDD.n1701 9.3005
R17675 VDD.n1739 VDD.n1738 9.3005
R17676 VDD.n1572 VDD.n1571 9.3005
R17677 VDD.n1567 VDD.n1566 9.3005
R17678 VDD.n1578 VDD.n1577 9.3005
R17679 VDD.n1580 VDD.n1579 9.3005
R17680 VDD.n1563 VDD.n1562 9.3005
R17681 VDD.n1586 VDD.n1585 9.3005
R17682 VDD.n1588 VDD.n1587 9.3005
R17683 VDD.n1560 VDD.n1557 9.3005
R17684 VDD.n1595 VDD.n1594 9.3005
R17685 VDD.n1623 VDD.n1622 9.3005
R17686 VDD.n1618 VDD.n1617 9.3005
R17687 VDD.n1629 VDD.n1628 9.3005
R17688 VDD.n1631 VDD.n1630 9.3005
R17689 VDD.n1614 VDD.n1613 9.3005
R17690 VDD.n1637 VDD.n1636 9.3005
R17691 VDD.n1639 VDD.n1638 9.3005
R17692 VDD.n1611 VDD.n1608 9.3005
R17693 VDD.n1646 VDD.n1645 9.3005
R17694 VDD.n2357 VDD.n1052 9.27678
R17695 VDD.n2363 VDD.n1052 9.27678
R17696 VDD.n2363 VDD.n1055 9.27678
R17697 VDD.n2369 VDD.n1048 9.27678
R17698 VDD.n2376 VDD.n1034 9.27678
R17699 VDD.n2382 VDD.n1034 9.27678
R17700 VDD.n2382 VDD.n1028 9.27678
R17701 VDD.n2388 VDD.n1028 9.27678
R17702 VDD.n2394 VDD.n1022 9.27678
R17703 VDD.n2400 VDD.n1016 9.27678
R17704 VDD.n2406 VDD.n1010 9.27678
R17705 VDD.n2412 VDD.n1004 9.27678
R17706 VDD.n2418 VDD.n998 9.27678
R17707 VDD.n2424 VDD.n987 9.27678
R17708 VDD.n2430 VDD.n987 9.27678
R17709 VDD.n2436 VDD.n975 9.27678
R17710 VDD.n2442 VDD.n975 9.27678
R17711 VDD.n2442 VDD.n978 9.27678
R17712 VDD.n2454 VDD.n964 9.27678
R17713 VDD.n2454 VDD.n958 9.27678
R17714 VDD.n2460 VDD.n958 9.27678
R17715 VDD.n2467 VDD.n951 9.27678
R17716 VDD.n2474 VDD.n947 9.27678
R17717 VDD.n2536 VDD.n903 9.27678
R17718 VDD.n2847 VDD.n2594 9.27678
R17719 VDD.n2853 VDD.n899 9.27678
R17720 VDD.n2859 VDD.n893 9.27678
R17721 VDD.n2865 VDD.n879 9.27678
R17722 VDD.n2871 VDD.n879 9.27678
R17723 VDD.n2871 VDD.n882 9.27678
R17724 VDD.n2883 VDD.n868 9.27678
R17725 VDD.n2883 VDD.n862 9.27678
R17726 VDD.n2889 VDD.n862 9.27678
R17727 VDD.n2895 VDD.n851 9.27678
R17728 VDD.n2901 VDD.n851 9.27678
R17729 VDD.n2907 VDD.n847 9.27678
R17730 VDD.n2913 VDD.n841 9.27678
R17731 VDD.n2919 VDD.n835 9.27678
R17732 VDD.n2925 VDD.n829 9.27678
R17733 VDD.n2931 VDD.n823 9.27678
R17734 VDD.n2937 VDD.n810 9.27678
R17735 VDD.n2943 VDD.n810 9.27678
R17736 VDD.n2943 VDD.n804 9.27678
R17737 VDD.n2949 VDD.n804 9.27678
R17738 VDD.n2992 VDD.n796 9.27678
R17739 VDD.n2998 VDD.n790 9.27678
R17740 VDD.n2998 VDD.n761 9.27678
R17741 VDD.n3053 VDD.n761 9.27678
R17742 VDD.n1186 VDD.t103 9.14036
R17743 VDD.t143 VDD.n1169 9.14036
R17744 VDD.n3301 VDD.t119 9.14036
R17745 VDD.t155 VDD.n3387 9.14036
R17746 VDD.n275 VDD.n274 8.92171
R17747 VDD.n224 VDD.n223 8.92171
R17748 VDD.n181 VDD.n180 8.92171
R17749 VDD.n130 VDD.n129 8.92171
R17750 VDD.n88 VDD.n87 8.92171
R17751 VDD.n37 VDD.n36 8.92171
R17752 VDD.n1764 VDD.n1763 8.92171
R17753 VDD.n1815 VDD.n1814 8.92171
R17754 VDD.n1670 VDD.n1669 8.92171
R17755 VDD.n1721 VDD.n1720 8.92171
R17756 VDD.n1577 VDD.n1576 8.92171
R17757 VDD.n1628 VDD.n1627 8.92171
R17758 VDD.t162 VDD.n1192 8.86753
R17759 VDD.n1163 VDD.t105 8.86753
R17760 VDD.t191 VDD.n998 8.86753
R17761 VDD.n2270 VDD.t79 8.86753
R17762 VDD.n2759 VDD.t82 8.86753
R17763 VDD.n847 VDD.t192 8.86753
R17764 VDD.n3282 VDD.t172 8.86753
R17765 VDD.n3379 VDD.t139 8.86753
R17766 VDD.t101 VDD.n1215 8.5947
R17767 VDD.n1139 VDD.t152 8.5947
R17768 VDD.n3249 VDD.t147 8.5947
R17769 VDD.n3363 VDD.t127 8.5947
R17770 VDD.n15 VDD.n14 8.35857
R17771 VDD.n2369 VDD.t7 8.32187
R17772 VDD.n2467 VDD.t30 8.32187
R17773 VDD.n2859 VDD.t60 8.32187
R17774 VDD.n2992 VDD.t50 8.32187
R17775 VDD.n271 VDD.n265 8.14595
R17776 VDD.n220 VDD.n214 8.14595
R17777 VDD.n177 VDD.n171 8.14595
R17778 VDD.n126 VDD.n120 8.14595
R17779 VDD.n84 VDD.n78 8.14595
R17780 VDD.n33 VDD.n27 8.14595
R17781 VDD.n1760 VDD.n1754 8.14595
R17782 VDD.n1811 VDD.n1805 8.14595
R17783 VDD.n1666 VDD.n1660 8.14595
R17784 VDD.n1717 VDD.n1711 8.14595
R17785 VDD.n1573 VDD.n1567 8.14595
R17786 VDD.n1624 VDD.n1618 8.14595
R17787 VDD.n3393 VDD.n3392 8.07375
R17788 VDD.n1838 VDD.n1837 8.07375
R17789 VDD.t92 VDD.n1010 8.04904
R17790 VDD.n2261 VDD.t210 8.04904
R17791 VDD.n2768 VDD.t78 8.04904
R17792 VDD.n835 VDD.t91 8.04904
R17793 VDD.n270 VDD.n267 7.3702
R17794 VDD.n219 VDD.n216 7.3702
R17795 VDD.n176 VDD.n173 7.3702
R17796 VDD.n125 VDD.n122 7.3702
R17797 VDD.n83 VDD.n80 7.3702
R17798 VDD.n32 VDD.n29 7.3702
R17799 VDD.n1759 VDD.n1756 7.3702
R17800 VDD.n1810 VDD.n1807 7.3702
R17801 VDD.n1665 VDD.n1662 7.3702
R17802 VDD.n1716 VDD.n1713 7.3702
R17803 VDD.n1572 VDD.n1569 7.3702
R17804 VDD.n1623 VDD.n1620 7.3702
R17805 VDD.n2394 VDD.t200 7.36696
R17806 VDD.n2931 VDD.t195 7.36696
R17807 VDD.n1469 VDD.t14 7.23054
R17808 VDD.t26 VDD.n1108 7.23054
R17809 VDD.t197 VDD.n1022 7.23054
R17810 VDD.n978 VDD.t90 7.23054
R17811 VDD.t83 VDD.n868 7.23054
R17812 VDD.n823 VDD.t211 7.23054
R17813 VDD.n3224 VDD.t3 7.23054
R17814 VDD.n3349 VDD.t18 7.23054
R17815 VDD.n2953 VDD.n2952 7.18099
R17816 VDD.n2373 VDD.n2372 7.18099
R17817 VDD.n202 VDD.n108 7.04468
R17818 VDD.n1742 VDD.n1648 7.04468
R17819 VDD.n1409 VDD.n1408 6.98232
R17820 VDD.n2040 VDD.n2039 6.98232
R17821 VDD.n534 VDD.n533 6.98232
R17822 VDD.n3132 VDD.n3129 6.98232
R17823 VDD.n2406 VDD.t198 6.54846
R17824 VDD.n2919 VDD.t84 6.54846
R17825 VDD.n1478 VDD.t14 6.41204
R17826 VDD.n1915 VDD.t26 6.41204
R17827 VDD.t3 VDD.n648 6.41204
R17828 VDD.t18 VDD.n350 6.41204
R17829 VDD.n1048 VDD.t46 6.27563
R17830 VDD.t22 VDD.n796 6.27563
R17831 VDD.n271 VDD.n270 5.81868
R17832 VDD.n220 VDD.n219 5.81868
R17833 VDD.n177 VDD.n176 5.81868
R17834 VDD.n126 VDD.n125 5.81868
R17835 VDD.n84 VDD.n83 5.81868
R17836 VDD.n33 VDD.n32 5.81868
R17837 VDD.n1760 VDD.n1759 5.81868
R17838 VDD.n1811 VDD.n1810 5.81868
R17839 VDD.n1666 VDD.n1665 5.81868
R17840 VDD.n1717 VDD.n1716 5.81868
R17841 VDD.n1573 VDD.n1572 5.81868
R17842 VDD.n1624 VDD.n1623 5.81868
R17843 VDD.n2487 VDD.n2486 5.77611
R17844 VDD.n2312 VDD.n1077 5.77611
R17845 VDD.n2670 VDD.n2669 5.77611
R17846 VDD.n787 VDD.n782 5.77611
R17847 VDD.n757 VDD.n752 5.77611
R17848 VDD.n2610 VDD.n2606 5.77611
R17849 VDD.n2546 VDD.n935 5.77611
R17850 VDD.n2183 VDD.n2182 5.77611
R17851 VDD.n2418 VDD.t202 5.72997
R17852 VDD.n2536 VDD.t88 5.72997
R17853 VDD.n2594 VDD.t86 5.72997
R17854 VDD.n2907 VDD.t193 5.72997
R17855 VDD.n1464 VDD.n1463 5.62474
R17856 VDD.n2118 VDD.n1103 5.62474
R17857 VDD.n3344 VDD.n394 5.62474
R17858 VDD.n3218 VDD.n660 5.62474
R17859 VDD.n7 VDD.t85 5.418
R17860 VDD.n7 VDD.t196 5.418
R17861 VDD.n8 VDD.t213 5.418
R17862 VDD.n8 VDD.t194 5.418
R17863 VDD.n10 VDD.t81 5.418
R17864 VDD.n10 VDD.t215 5.418
R17865 VDD.n12 VDD.t209 5.418
R17866 VDD.n12 VDD.t87 5.418
R17867 VDD.n5 VDD.t89 5.418
R17868 VDD.n5 VDD.t207 5.418
R17869 VDD.n3 VDD.t1 5.418
R17870 VDD.n3 VDD.t94 5.418
R17871 VDD.n1 VDD.t203 5.418
R17872 VDD.n1 VDD.t205 5.418
R17873 VDD.n0 VDD.t201 5.418
R17874 VDD.n0 VDD.t199 5.418
R17875 VDD.n2332 VDD.n1069 5.30782
R17876 VDD.n2328 VDD.n1069 5.30782
R17877 VDD.n3029 VDD.n3028 5.30782
R17878 VDD.n3028 VDD.n3026 5.30782
R17879 VDD.n3078 VDD.n745 5.30782
R17880 VDD.n3078 VDD.n3077 5.30782
R17881 VDD.n2133 VDD.n2132 5.30782
R17882 VDD.n2165 VDD.n2132 5.30782
R17883 VDD.n2448 VDD.t0 5.1843
R17884 VDD.n2877 VDD.t214 5.1843
R17885 VDD.n1494 VDD.t101 5.04789
R17886 VDD.n1898 VDD.t152 5.04789
R17887 VDD.n3240 VDD.t147 5.04789
R17888 VDD.n346 VDD.t127 5.04789
R17889 VDD.n274 VDD.n265 5.04292
R17890 VDD.n223 VDD.n214 5.04292
R17891 VDD.n180 VDD.n171 5.04292
R17892 VDD.n129 VDD.n120 5.04292
R17893 VDD.n87 VDD.n78 5.04292
R17894 VDD.n36 VDD.n27 5.04292
R17895 VDD.n1763 VDD.n1754 5.04292
R17896 VDD.n1814 VDD.n1805 5.04292
R17897 VDD.n1669 VDD.n1660 5.04292
R17898 VDD.n1720 VDD.n1711 5.04292
R17899 VDD.n1576 VDD.n1567 5.04292
R17900 VDD.n1627 VDD.n1618 5.04292
R17901 VDD.n2430 VDD.t204 4.91147
R17902 VDD.t93 VDD.n951 4.91147
R17903 VDD.t206 VDD.n2590 4.91147
R17904 VDD.n2591 VDD.t208 4.91147
R17905 VDD.n893 VDD.t80 4.91147
R17906 VDD.n2895 VDD.t212 4.91147
R17907 VDD.n2486 VDD.n2485 4.83952
R17908 VDD.n2308 VDD.n1077 4.83952
R17909 VDD.n2671 VDD.n2670 4.83952
R17910 VDD.n3007 VDD.n787 4.83952
R17911 VDD.n3058 VDD.n757 4.83952
R17912 VDD.n2797 VDD.n2610 4.83952
R17913 VDD.n2543 VDD.n935 4.83952
R17914 VDD.n2184 VDD.n2183 4.83952
R17915 VDD.n1527 VDD.t162 4.77505
R17916 VDD.n1866 VDD.t105 4.77505
R17917 VDD.n3273 VDD.t172 4.77505
R17918 VDD.n324 VDD.t139 4.77505
R17919 VDD.n2010 VDD.n1089 4.74817
R17920 VDD.n2015 VDD.n1090 4.74817
R17921 VDD.n2096 VDD.n2095 4.74817
R17922 VDD.n2093 VDD.n1935 4.74817
R17923 VDD.n2095 VDD.n1933 4.74817
R17924 VDD.n2093 VDD.n2092 4.74817
R17925 VDD.n3200 VDD.n703 4.74817
R17926 VDD.n3193 VDD.n704 4.74817
R17927 VDD.n3196 VDD.n704 4.74817
R17928 VDD.n3197 VDD.n703 4.74817
R17929 VDD.n3103 VDD.n743 4.74817
R17930 VDD.n3099 VDD.n744 4.74817
R17931 VDD.n3102 VDD.n744 4.74817
R17932 VDD.n3106 VDD.n743 4.74817
R17933 VDD.n2016 VDD.n1089 4.74817
R17934 VDD.n1092 VDD.n1090 4.74817
R17935 VDD.n296 VDD.n295 4.7074
R17936 VDD.n202 VDD.n201 4.7074
R17937 VDD.n1836 VDD.n1835 4.7074
R17938 VDD.n1742 VDD.n1741 4.7074
R17939 VDD.n1552 VDD.t103 4.50222
R17940 VDD.n1842 VDD.t143 4.50222
R17941 VDD.t119 VDD.n303 4.50222
R17942 VDD.n3388 VDD.t155 4.50222
R17943 VDD.n3393 VDD.n296 4.47685
R17944 VDD.n1837 VDD.n1836 4.47685
R17945 VDD.n2261 VDD.t204 4.36581
R17946 VDD.n2460 VDD.t93 4.36581
R17947 VDD.n2865 VDD.t80 4.36581
R17948 VDD.n2768 VDD.t212 4.36581
R17949 VDD.n275 VDD.n263 4.26717
R17950 VDD.n224 VDD.n212 4.26717
R17951 VDD.n181 VDD.n169 4.26717
R17952 VDD.n130 VDD.n118 4.26717
R17953 VDD.n88 VDD.n76 4.26717
R17954 VDD.n37 VDD.n25 4.26717
R17955 VDD.n1764 VDD.n1752 4.26717
R17956 VDD.n1815 VDD.n1803 4.26717
R17957 VDD.n1670 VDD.n1658 4.26717
R17958 VDD.n1721 VDD.n1709 4.26717
R17959 VDD.n1577 VDD.n1565 4.26717
R17960 VDD.n1628 VDD.n1616 4.26717
R17961 VDD.n1519 VDD.t115 4.22939
R17962 VDD.n1874 VDD.t124 4.22939
R17963 VDD.t108 VDD.n619 4.22939
R17964 VDD.n3372 VDD.t95 4.22939
R17965 VDD.t0 VDD.n964 4.09298
R17966 VDD.n882 VDD.t214 4.09298
R17967 VDD.n252 VDD.t96 4.06363
R17968 VDD.n252 VDD.t134 4.06363
R17969 VDD.n250 VDD.t121 4.06363
R17970 VDD.n250 VDD.t151 4.06363
R17971 VDD.n248 VDD.t133 4.06363
R17972 VDD.n248 VDD.t170 4.06363
R17973 VDD.n246 VDD.t180 4.06363
R17974 VDD.n246 VDD.t190 4.06363
R17975 VDD.n244 VDD.t169 4.06363
R17976 VDD.n244 VDD.t109 4.06363
R17977 VDD.n158 VDD.t181 4.06363
R17978 VDD.n158 VDD.t123 4.06363
R17979 VDD.n156 VDD.t112 4.06363
R17980 VDD.n156 VDD.t140 4.06363
R17981 VDD.n154 VDD.t120 4.06363
R17982 VDD.n154 VDD.t161 4.06363
R17983 VDD.n152 VDD.t173 4.06363
R17984 VDD.n152 VDD.t179 4.06363
R17985 VDD.n150 VDD.t158 4.06363
R17986 VDD.n150 VDD.t189 4.06363
R17987 VDD.n65 VDD.t166 4.06363
R17988 VDD.n65 VDD.t146 4.06363
R17989 VDD.n63 VDD.t111 4.06363
R17990 VDD.n63 VDD.t182 4.06363
R17991 VDD.n61 VDD.t175 4.06363
R17992 VDD.n61 VDD.t156 4.06363
R17993 VDD.n59 VDD.t187 4.06363
R17994 VDD.n59 VDD.t98 4.06363
R17995 VDD.n57 VDD.t184 4.06363
R17996 VDD.n57 VDD.t165 4.06363
R17997 VDD.n1784 VDD.t135 4.06363
R17998 VDD.n1784 VDD.t100 4.06363
R17999 VDD.n1786 VDD.t126 4.06363
R18000 VDD.n1786 VDD.t107 4.06363
R18001 VDD.n1788 VDD.t104 4.06363
R18002 VDD.n1788 VDD.t154 4.06363
R18003 VDD.n1790 VDD.t178 4.06363
R18004 VDD.n1790 VDD.t136 4.06363
R18005 VDD.n1792 VDD.t159 4.06363
R18006 VDD.n1792 VDD.t130 4.06363
R18007 VDD.n1690 VDD.t125 4.06363
R18008 VDD.n1690 VDD.t183 4.06363
R18009 VDD.n1692 VDD.t114 4.06363
R18010 VDD.n1692 VDD.t188 4.06363
R18011 VDD.n1694 VDD.t186 4.06363
R18012 VDD.n1694 VDD.t144 4.06363
R18013 VDD.n1696 VDD.t168 4.06363
R18014 VDD.n1696 VDD.t129 4.06363
R18015 VDD.n1698 VDD.t145 4.06363
R18016 VDD.n1698 VDD.t116 4.06363
R18017 VDD.n1597 VDD.t141 4.06363
R18018 VDD.n1597 VDD.t164 4.06363
R18019 VDD.n1599 VDD.t171 4.06363
R18020 VDD.n1599 VDD.t106 4.06363
R18021 VDD.n1601 VDD.t137 4.06363
R18022 VDD.n1601 VDD.t150 4.06363
R18023 VDD.n1603 VDD.t163 4.06363
R18024 VDD.n1603 VDD.t118 4.06363
R18025 VDD.n1605 VDD.t132 4.06363
R18026 VDD.n1605 VDD.t142 4.06363
R18027 VDD.n2270 VDD.t202 3.54731
R18028 VDD.n2474 VDD.t88 3.54731
R18029 VDD.n2853 VDD.t86 3.54731
R18030 VDD.n2759 VDD.t193 3.54731
R18031 VDD.n279 VDD.n278 3.49141
R18032 VDD.n228 VDD.n227 3.49141
R18033 VDD.n185 VDD.n184 3.49141
R18034 VDD.n134 VDD.n133 3.49141
R18035 VDD.n92 VDD.n91 3.49141
R18036 VDD.n41 VDD.n40 3.49141
R18037 VDD.n1768 VDD.n1767 3.49141
R18038 VDD.n1819 VDD.n1818 3.49141
R18039 VDD.n1674 VDD.n1673 3.49141
R18040 VDD.n1725 VDD.n1724 3.49141
R18041 VDD.n1581 VDD.n1580 3.49141
R18042 VDD.n1632 VDD.n1631 3.49141
R18043 VDD.n2952 VDD.n2951 3.43465
R18044 VDD.n2374 VDD.n2373 3.43465
R18045 VDD.n2376 VDD.t46 3.00165
R18046 VDD.n2949 VDD.t22 3.00165
R18047 VDD.t198 VDD.n1004 2.72882
R18048 VDD.n841 VDD.t84 2.72882
R18049 VDD.n282 VDD.n261 2.71565
R18050 VDD.n231 VDD.n210 2.71565
R18051 VDD.n188 VDD.n167 2.71565
R18052 VDD.n137 VDD.n116 2.71565
R18053 VDD.n95 VDD.n74 2.71565
R18054 VDD.n44 VDD.n23 2.71565
R18055 VDD.n1771 VDD.n1750 2.71565
R18056 VDD.n1822 VDD.n1801 2.71565
R18057 VDD.n1677 VDD.n1656 2.71565
R18058 VDD.n1728 VDD.n1707 2.71565
R18059 VDD.n1584 VDD.n1563 2.71565
R18060 VDD.n1635 VDD.n1614 2.71565
R18061 VDD.n269 VDD.n268 2.4129
R18062 VDD.n218 VDD.n217 2.4129
R18063 VDD.n175 VDD.n174 2.4129
R18064 VDD.n124 VDD.n123 2.4129
R18065 VDD.n82 VDD.n81 2.4129
R18066 VDD.n31 VDD.n30 2.4129
R18067 VDD.n1758 VDD.n1757 2.4129
R18068 VDD.n1809 VDD.n1808 2.4129
R18069 VDD.n1664 VDD.n1663 2.4129
R18070 VDD.n1715 VDD.n1714 2.4129
R18071 VDD.n1571 VDD.n1570 2.4129
R18072 VDD.n1622 VDD.n1621 2.4129
R18073 VDD.n296 VDD.n202 2.33778
R18074 VDD.n1836 VDD.n1742 2.33778
R18075 VDD.n2095 VDD.n2094 2.27742
R18076 VDD.n2094 VDD.n2093 2.27742
R18077 VDD.n3027 VDD.n704 2.27742
R18078 VDD.n3027 VDD.n703 2.27742
R18079 VDD.n3079 VDD.n744 2.27742
R18080 VDD.n3079 VDD.n743 2.27742
R18081 VDD.n2131 VDD.n1089 2.27742
R18082 VDD.n2131 VDD.n1090 2.27742
R18083 VDD.n2388 VDD.t197 2.04674
R18084 VDD.n2448 VDD.t90 2.04674
R18085 VDD.n2877 VDD.t83 2.04674
R18086 VDD.n2937 VDD.t211 2.04674
R18087 VDD.n283 VDD.n259 1.93989
R18088 VDD.n232 VDD.n208 1.93989
R18089 VDD.n189 VDD.n165 1.93989
R18090 VDD.n138 VDD.n114 1.93989
R18091 VDD.n96 VDD.n72 1.93989
R18092 VDD.n45 VDD.n21 1.93989
R18093 VDD.n1772 VDD.n1748 1.93989
R18094 VDD.n1823 VDD.n1799 1.93989
R18095 VDD.n1678 VDD.n1654 1.93989
R18096 VDD.n1729 VDD.n1705 1.93989
R18097 VDD.n1585 VDD.n1561 1.93989
R18098 VDD.n1636 VDD.n1612 1.93989
R18099 VDD.t200 VDD.n1016 1.91032
R18100 VDD.n829 VDD.t195 1.91032
R18101 VDD.n2400 VDD.t92 1.22824
R18102 VDD.n2436 VDD.t210 1.22824
R18103 VDD.n2889 VDD.t78 1.22824
R18104 VDD.n2925 VDD.t91 1.22824
R18105 VDD.n294 VDD.n254 1.16414
R18106 VDD.n287 VDD.n286 1.16414
R18107 VDD.n243 VDD.n203 1.16414
R18108 VDD.n236 VDD.n235 1.16414
R18109 VDD.n200 VDD.n160 1.16414
R18110 VDD.n193 VDD.n192 1.16414
R18111 VDD.n149 VDD.n109 1.16414
R18112 VDD.n142 VDD.n141 1.16414
R18113 VDD.n107 VDD.n67 1.16414
R18114 VDD.n100 VDD.n99 1.16414
R18115 VDD.n56 VDD.n16 1.16414
R18116 VDD.n49 VDD.n48 1.16414
R18117 VDD.n1783 VDD.n1743 1.16414
R18118 VDD.n1776 VDD.n1775 1.16414
R18119 VDD.n1834 VDD.n1794 1.16414
R18120 VDD.n1827 VDD.n1826 1.16414
R18121 VDD.n1689 VDD.n1649 1.16414
R18122 VDD.n1682 VDD.n1681 1.16414
R18123 VDD.n1740 VDD.n1700 1.16414
R18124 VDD.n1733 VDD.n1732 1.16414
R18125 VDD.n1596 VDD.n1556 1.16414
R18126 VDD.n1589 VDD.n1588 1.16414
R18127 VDD.n1647 VDD.n1607 1.16414
R18128 VDD.n1640 VDD.n1639 1.16414
R18129 VDD.n1837 VDD.n15 1.00254
R18130 VDD VDD.n3393 0.994707
R18131 VDD.n1463 VDD.n1462 0.970197
R18132 VDD.n2121 VDD.n1103 0.970197
R18133 VDD.n586 VDD.n394 0.970197
R18134 VDD.n3086 VDD.n660 0.970197
R18135 VDD.n1055 VDD.t7 0.955411
R18136 VDD.t30 VDD.n947 0.955411
R18137 VDD.n899 VDD.t60 0.955411
R18138 VDD.t50 VDD.n790 0.955411
R18139 VDD.n4 VDD.n2 0.728948
R18140 VDD.n11 VDD.n9 0.728948
R18141 VDD.n247 VDD.n245 0.573776
R18142 VDD.n249 VDD.n247 0.573776
R18143 VDD.n251 VDD.n249 0.573776
R18144 VDD.n253 VDD.n251 0.573776
R18145 VDD.n295 VDD.n253 0.573776
R18146 VDD.n153 VDD.n151 0.573776
R18147 VDD.n155 VDD.n153 0.573776
R18148 VDD.n157 VDD.n155 0.573776
R18149 VDD.n159 VDD.n157 0.573776
R18150 VDD.n201 VDD.n159 0.573776
R18151 VDD.n60 VDD.n58 0.573776
R18152 VDD.n62 VDD.n60 0.573776
R18153 VDD.n64 VDD.n62 0.573776
R18154 VDD.n66 VDD.n64 0.573776
R18155 VDD.n108 VDD.n66 0.573776
R18156 VDD.n1835 VDD.n1793 0.573776
R18157 VDD.n1793 VDD.n1791 0.573776
R18158 VDD.n1791 VDD.n1789 0.573776
R18159 VDD.n1789 VDD.n1787 0.573776
R18160 VDD.n1787 VDD.n1785 0.573776
R18161 VDD.n1741 VDD.n1699 0.573776
R18162 VDD.n1699 VDD.n1697 0.573776
R18163 VDD.n1697 VDD.n1695 0.573776
R18164 VDD.n1695 VDD.n1693 0.573776
R18165 VDD.n1693 VDD.n1691 0.573776
R18166 VDD.n1648 VDD.n1606 0.573776
R18167 VDD.n1606 VDD.n1604 0.573776
R18168 VDD.n1604 VDD.n1602 0.573776
R18169 VDD.n1602 VDD.n1600 0.573776
R18170 VDD.n1600 VDD.n1598 0.573776
R18171 VDD.n6 VDD.n4 0.573776
R18172 VDD.n13 VDD.n11 0.573776
R18173 VDD.n14 VDD.n6 0.49619
R18174 VDD.n14 VDD.n13 0.49619
R18175 VDD.n2112 VDD.n2111 0.495927
R18176 VDD.n695 VDD.n651 0.495927
R18177 VDD.n431 VDD.n430 0.495927
R18178 VDD.n3343 VDD.n3342 0.495927
R18179 VDD.n3220 VDD.n3219 0.495927
R18180 VDD.n2119 VDD.n1104 0.495927
R18181 VDD.n1466 VDD.n1465 0.495927
R18182 VDD.n1473 VDD.n1235 0.495927
R18183 VDD.n1502 VDD.t131 0.409748
R18184 VDD.t99 VDD.n1138 0.409748
R18185 VDD.n2412 VDD.t191 0.409748
R18186 VDD.n2424 VDD.t79 0.409748
R18187 VDD.n2901 VDD.t82 0.409748
R18188 VDD.n2913 VDD.t192 0.409748
R18189 VDD.n3257 VDD.t157 0.409748
R18190 VDD.n3365 VDD.t122 0.409748
R18191 VDD.n292 VDD.n291 0.388379
R18192 VDD.n258 VDD.n256 0.388379
R18193 VDD.n241 VDD.n240 0.388379
R18194 VDD.n207 VDD.n205 0.388379
R18195 VDD.n198 VDD.n197 0.388379
R18196 VDD.n164 VDD.n162 0.388379
R18197 VDD.n147 VDD.n146 0.388379
R18198 VDD.n113 VDD.n111 0.388379
R18199 VDD.n105 VDD.n104 0.388379
R18200 VDD.n71 VDD.n69 0.388379
R18201 VDD.n54 VDD.n53 0.388379
R18202 VDD.n20 VDD.n18 0.388379
R18203 VDD.n1781 VDD.n1780 0.388379
R18204 VDD.n1747 VDD.n1745 0.388379
R18205 VDD.n1832 VDD.n1831 0.388379
R18206 VDD.n1798 VDD.n1796 0.388379
R18207 VDD.n1687 VDD.n1686 0.388379
R18208 VDD.n1653 VDD.n1651 0.388379
R18209 VDD.n1738 VDD.n1737 0.388379
R18210 VDD.n1704 VDD.n1702 0.388379
R18211 VDD.n1594 VDD.n1593 0.388379
R18212 VDD.n1560 VDD.n1558 0.388379
R18213 VDD.n1645 VDD.n1644 0.388379
R18214 VDD.n1611 VDD.n1609 0.388379
R18215 VDD.n293 VDD.n255 0.155672
R18216 VDD.n285 VDD.n255 0.155672
R18217 VDD.n285 VDD.n284 0.155672
R18218 VDD.n284 VDD.n260 0.155672
R18219 VDD.n277 VDD.n260 0.155672
R18220 VDD.n277 VDD.n276 0.155672
R18221 VDD.n276 VDD.n264 0.155672
R18222 VDD.n269 VDD.n264 0.155672
R18223 VDD.n242 VDD.n204 0.155672
R18224 VDD.n234 VDD.n204 0.155672
R18225 VDD.n234 VDD.n233 0.155672
R18226 VDD.n233 VDD.n209 0.155672
R18227 VDD.n226 VDD.n209 0.155672
R18228 VDD.n226 VDD.n225 0.155672
R18229 VDD.n225 VDD.n213 0.155672
R18230 VDD.n218 VDD.n213 0.155672
R18231 VDD.n199 VDD.n161 0.155672
R18232 VDD.n191 VDD.n161 0.155672
R18233 VDD.n191 VDD.n190 0.155672
R18234 VDD.n190 VDD.n166 0.155672
R18235 VDD.n183 VDD.n166 0.155672
R18236 VDD.n183 VDD.n182 0.155672
R18237 VDD.n182 VDD.n170 0.155672
R18238 VDD.n175 VDD.n170 0.155672
R18239 VDD.n148 VDD.n110 0.155672
R18240 VDD.n140 VDD.n110 0.155672
R18241 VDD.n140 VDD.n139 0.155672
R18242 VDD.n139 VDD.n115 0.155672
R18243 VDD.n132 VDD.n115 0.155672
R18244 VDD.n132 VDD.n131 0.155672
R18245 VDD.n131 VDD.n119 0.155672
R18246 VDD.n124 VDD.n119 0.155672
R18247 VDD.n106 VDD.n68 0.155672
R18248 VDD.n98 VDD.n68 0.155672
R18249 VDD.n98 VDD.n97 0.155672
R18250 VDD.n97 VDD.n73 0.155672
R18251 VDD.n90 VDD.n73 0.155672
R18252 VDD.n90 VDD.n89 0.155672
R18253 VDD.n89 VDD.n77 0.155672
R18254 VDD.n82 VDD.n77 0.155672
R18255 VDD.n55 VDD.n17 0.155672
R18256 VDD.n47 VDD.n17 0.155672
R18257 VDD.n47 VDD.n46 0.155672
R18258 VDD.n46 VDD.n22 0.155672
R18259 VDD.n39 VDD.n22 0.155672
R18260 VDD.n39 VDD.n38 0.155672
R18261 VDD.n38 VDD.n26 0.155672
R18262 VDD.n31 VDD.n26 0.155672
R18263 VDD.n1782 VDD.n1744 0.155672
R18264 VDD.n1774 VDD.n1744 0.155672
R18265 VDD.n1774 VDD.n1773 0.155672
R18266 VDD.n1773 VDD.n1749 0.155672
R18267 VDD.n1766 VDD.n1749 0.155672
R18268 VDD.n1766 VDD.n1765 0.155672
R18269 VDD.n1765 VDD.n1753 0.155672
R18270 VDD.n1758 VDD.n1753 0.155672
R18271 VDD.n1833 VDD.n1795 0.155672
R18272 VDD.n1825 VDD.n1795 0.155672
R18273 VDD.n1825 VDD.n1824 0.155672
R18274 VDD.n1824 VDD.n1800 0.155672
R18275 VDD.n1817 VDD.n1800 0.155672
R18276 VDD.n1817 VDD.n1816 0.155672
R18277 VDD.n1816 VDD.n1804 0.155672
R18278 VDD.n1809 VDD.n1804 0.155672
R18279 VDD.n1688 VDD.n1650 0.155672
R18280 VDD.n1680 VDD.n1650 0.155672
R18281 VDD.n1680 VDD.n1679 0.155672
R18282 VDD.n1679 VDD.n1655 0.155672
R18283 VDD.n1672 VDD.n1655 0.155672
R18284 VDD.n1672 VDD.n1671 0.155672
R18285 VDD.n1671 VDD.n1659 0.155672
R18286 VDD.n1664 VDD.n1659 0.155672
R18287 VDD.n1739 VDD.n1701 0.155672
R18288 VDD.n1731 VDD.n1701 0.155672
R18289 VDD.n1731 VDD.n1730 0.155672
R18290 VDD.n1730 VDD.n1706 0.155672
R18291 VDD.n1723 VDD.n1706 0.155672
R18292 VDD.n1723 VDD.n1722 0.155672
R18293 VDD.n1722 VDD.n1710 0.155672
R18294 VDD.n1715 VDD.n1710 0.155672
R18295 VDD.n1595 VDD.n1557 0.155672
R18296 VDD.n1587 VDD.n1557 0.155672
R18297 VDD.n1587 VDD.n1586 0.155672
R18298 VDD.n1586 VDD.n1562 0.155672
R18299 VDD.n1579 VDD.n1562 0.155672
R18300 VDD.n1579 VDD.n1578 0.155672
R18301 VDD.n1578 VDD.n1566 0.155672
R18302 VDD.n1571 VDD.n1566 0.155672
R18303 VDD.n1646 VDD.n1608 0.155672
R18304 VDD.n1638 VDD.n1608 0.155672
R18305 VDD.n1638 VDD.n1637 0.155672
R18306 VDD.n1637 VDD.n1613 0.155672
R18307 VDD.n1630 VDD.n1613 0.155672
R18308 VDD.n1630 VDD.n1629 0.155672
R18309 VDD.n1629 VDD.n1617 0.155672
R18310 VDD.n1622 VDD.n1617 0.155672
R18311 VDD.n1839 VDD.n1166 0.152939
R18312 VDD.n1853 VDD.n1166 0.152939
R18313 VDD.n1854 VDD.n1853 0.152939
R18314 VDD.n1855 VDD.n1854 0.152939
R18315 VDD.n1855 VDD.n1154 0.152939
R18316 VDD.n1869 VDD.n1154 0.152939
R18317 VDD.n1870 VDD.n1869 0.152939
R18318 VDD.n1871 VDD.n1870 0.152939
R18319 VDD.n1871 VDD.n1142 0.152939
R18320 VDD.n1885 VDD.n1142 0.152939
R18321 VDD.n1886 VDD.n1885 0.152939
R18322 VDD.n1887 VDD.n1886 0.152939
R18323 VDD.n1887 VDD.n1130 0.152939
R18324 VDD.n1901 VDD.n1130 0.152939
R18325 VDD.n1902 VDD.n1901 0.152939
R18326 VDD.n1903 VDD.n1902 0.152939
R18327 VDD.n1903 VDD.n1117 0.152939
R18328 VDD.n1918 VDD.n1117 0.152939
R18329 VDD.n1919 VDD.n1918 0.152939
R18330 VDD.n2112 VDD.n1919 0.152939
R18331 VDD.n2111 VDD.n1920 0.152939
R18332 VDD.n1924 VDD.n1920 0.152939
R18333 VDD.n1925 VDD.n1924 0.152939
R18334 VDD.n1926 VDD.n1925 0.152939
R18335 VDD.n1927 VDD.n1926 0.152939
R18336 VDD.n1931 VDD.n1927 0.152939
R18337 VDD.n1932 VDD.n1931 0.152939
R18338 VDD.n1942 VDD.n1934 0.152939
R18339 VDD.n1943 VDD.n1942 0.152939
R18340 VDD.n1944 VDD.n1943 0.152939
R18341 VDD.n1948 VDD.n1944 0.152939
R18342 VDD.n1949 VDD.n1948 0.152939
R18343 VDD.n1950 VDD.n1949 0.152939
R18344 VDD.n2077 VDD.n1950 0.152939
R18345 VDD.n2077 VDD.n2076 0.152939
R18346 VDD.n2076 VDD.n2075 0.152939
R18347 VDD.n2075 VDD.n1956 0.152939
R18348 VDD.n1961 VDD.n1956 0.152939
R18349 VDD.n1962 VDD.n1961 0.152939
R18350 VDD.n1963 VDD.n1962 0.152939
R18351 VDD.n1967 VDD.n1963 0.152939
R18352 VDD.n1968 VDD.n1967 0.152939
R18353 VDD.n1969 VDD.n1968 0.152939
R18354 VDD.n1970 VDD.n1969 0.152939
R18355 VDD.n1974 VDD.n1970 0.152939
R18356 VDD.n1975 VDD.n1974 0.152939
R18357 VDD.n1976 VDD.n1975 0.152939
R18358 VDD.n1977 VDD.n1976 0.152939
R18359 VDD.n1981 VDD.n1977 0.152939
R18360 VDD.n1982 VDD.n1981 0.152939
R18361 VDD.n1983 VDD.n1982 0.152939
R18362 VDD.n1984 VDD.n1983 0.152939
R18363 VDD.n1988 VDD.n1984 0.152939
R18364 VDD.n1989 VDD.n1988 0.152939
R18365 VDD.n1990 VDD.n1989 0.152939
R18366 VDD.n2038 VDD.n1990 0.152939
R18367 VDD.n2038 VDD.n2037 0.152939
R18368 VDD.n2037 VDD.n2036 0.152939
R18369 VDD.n2036 VDD.n1996 0.152939
R18370 VDD.n2001 VDD.n1996 0.152939
R18371 VDD.n2002 VDD.n2001 0.152939
R18372 VDD.n2003 VDD.n2002 0.152939
R18373 VDD.n2007 VDD.n2003 0.152939
R18374 VDD.n2008 VDD.n2007 0.152939
R18375 VDD.n2009 VDD.n2008 0.152939
R18376 VDD.n2009 VDD.n1088 0.152939
R18377 VDD.n706 VDD.n705 0.152939
R18378 VDD.n707 VDD.n706 0.152939
R18379 VDD.n708 VDD.n707 0.152939
R18380 VDD.n709 VDD.n708 0.152939
R18381 VDD.n710 VDD.n709 0.152939
R18382 VDD.n711 VDD.n710 0.152939
R18383 VDD.n3174 VDD.n711 0.152939
R18384 VDD.n3174 VDD.n3173 0.152939
R18385 VDD.n3173 VDD.n3172 0.152939
R18386 VDD.n3172 VDD.n713 0.152939
R18387 VDD.n714 VDD.n713 0.152939
R18388 VDD.n715 VDD.n714 0.152939
R18389 VDD.n716 VDD.n715 0.152939
R18390 VDD.n717 VDD.n716 0.152939
R18391 VDD.n718 VDD.n717 0.152939
R18392 VDD.n719 VDD.n718 0.152939
R18393 VDD.n720 VDD.n719 0.152939
R18394 VDD.n721 VDD.n720 0.152939
R18395 VDD.n722 VDD.n721 0.152939
R18396 VDD.n723 VDD.n722 0.152939
R18397 VDD.n724 VDD.n723 0.152939
R18398 VDD.n725 VDD.n724 0.152939
R18399 VDD.n726 VDD.n725 0.152939
R18400 VDD.n727 VDD.n726 0.152939
R18401 VDD.n728 VDD.n727 0.152939
R18402 VDD.n729 VDD.n728 0.152939
R18403 VDD.n730 VDD.n729 0.152939
R18404 VDD.n731 VDD.n730 0.152939
R18405 VDD.n3128 VDD.n731 0.152939
R18406 VDD.n3128 VDD.n3127 0.152939
R18407 VDD.n3127 VDD.n3126 0.152939
R18408 VDD.n3126 VDD.n735 0.152939
R18409 VDD.n736 VDD.n735 0.152939
R18410 VDD.n737 VDD.n736 0.152939
R18411 VDD.n738 VDD.n737 0.152939
R18412 VDD.n739 VDD.n738 0.152939
R18413 VDD.n740 VDD.n739 0.152939
R18414 VDD.n741 VDD.n740 0.152939
R18415 VDD.n742 VDD.n741 0.152939
R18416 VDD.n696 VDD.n695 0.152939
R18417 VDD.n697 VDD.n696 0.152939
R18418 VDD.n698 VDD.n697 0.152939
R18419 VDD.n699 VDD.n698 0.152939
R18420 VDD.n700 VDD.n699 0.152939
R18421 VDD.n701 VDD.n700 0.152939
R18422 VDD.n702 VDD.n701 0.152939
R18423 VDD.n3227 VDD.n651 0.152939
R18424 VDD.n3228 VDD.n3227 0.152939
R18425 VDD.n3229 VDD.n3228 0.152939
R18426 VDD.n3229 VDD.n639 0.152939
R18427 VDD.n3244 VDD.n639 0.152939
R18428 VDD.n3245 VDD.n3244 0.152939
R18429 VDD.n3246 VDD.n3245 0.152939
R18430 VDD.n3246 VDD.n628 0.152939
R18431 VDD.n3260 VDD.n628 0.152939
R18432 VDD.n3261 VDD.n3260 0.152939
R18433 VDD.n3262 VDD.n3261 0.152939
R18434 VDD.n3262 VDD.n616 0.152939
R18435 VDD.n3277 VDD.n616 0.152939
R18436 VDD.n3278 VDD.n3277 0.152939
R18437 VDD.n3279 VDD.n3278 0.152939
R18438 VDD.n3279 VDD.n605 0.152939
R18439 VDD.n3296 VDD.n605 0.152939
R18440 VDD.n3297 VDD.n3296 0.152939
R18441 VDD.n3298 VDD.n3297 0.152939
R18442 VDD.n3298 VDD.n297 0.152939
R18443 VDD.n309 VDD.n298 0.152939
R18444 VDD.n310 VDD.n309 0.152939
R18445 VDD.n311 VDD.n310 0.152939
R18446 VDD.n318 VDD.n311 0.152939
R18447 VDD.n319 VDD.n318 0.152939
R18448 VDD.n320 VDD.n319 0.152939
R18449 VDD.n321 VDD.n320 0.152939
R18450 VDD.n330 VDD.n321 0.152939
R18451 VDD.n331 VDD.n330 0.152939
R18452 VDD.n332 VDD.n331 0.152939
R18453 VDD.n333 VDD.n332 0.152939
R18454 VDD.n340 VDD.n333 0.152939
R18455 VDD.n341 VDD.n340 0.152939
R18456 VDD.n342 VDD.n341 0.152939
R18457 VDD.n343 VDD.n342 0.152939
R18458 VDD.n352 VDD.n343 0.152939
R18459 VDD.n353 VDD.n352 0.152939
R18460 VDD.n354 VDD.n353 0.152939
R18461 VDD.n355 VDD.n354 0.152939
R18462 VDD.n430 VDD.n355 0.152939
R18463 VDD.n431 VDD.n429 0.152939
R18464 VDD.n438 VDD.n429 0.152939
R18465 VDD.n439 VDD.n438 0.152939
R18466 VDD.n440 VDD.n439 0.152939
R18467 VDD.n440 VDD.n427 0.152939
R18468 VDD.n448 VDD.n427 0.152939
R18469 VDD.n449 VDD.n448 0.152939
R18470 VDD.n450 VDD.n449 0.152939
R18471 VDD.n450 VDD.n425 0.152939
R18472 VDD.n458 VDD.n425 0.152939
R18473 VDD.n459 VDD.n458 0.152939
R18474 VDD.n460 VDD.n459 0.152939
R18475 VDD.n460 VDD.n423 0.152939
R18476 VDD.n468 VDD.n423 0.152939
R18477 VDD.n469 VDD.n468 0.152939
R18478 VDD.n470 VDD.n469 0.152939
R18479 VDD.n470 VDD.n421 0.152939
R18480 VDD.n478 VDD.n421 0.152939
R18481 VDD.n479 VDD.n478 0.152939
R18482 VDD.n480 VDD.n479 0.152939
R18483 VDD.n480 VDD.n417 0.152939
R18484 VDD.n488 VDD.n417 0.152939
R18485 VDD.n489 VDD.n488 0.152939
R18486 VDD.n490 VDD.n489 0.152939
R18487 VDD.n490 VDD.n415 0.152939
R18488 VDD.n498 VDD.n415 0.152939
R18489 VDD.n499 VDD.n498 0.152939
R18490 VDD.n500 VDD.n499 0.152939
R18491 VDD.n500 VDD.n413 0.152939
R18492 VDD.n508 VDD.n413 0.152939
R18493 VDD.n509 VDD.n508 0.152939
R18494 VDD.n510 VDD.n509 0.152939
R18495 VDD.n510 VDD.n411 0.152939
R18496 VDD.n518 VDD.n411 0.152939
R18497 VDD.n519 VDD.n518 0.152939
R18498 VDD.n520 VDD.n519 0.152939
R18499 VDD.n520 VDD.n409 0.152939
R18500 VDD.n528 VDD.n409 0.152939
R18501 VDD.n529 VDD.n528 0.152939
R18502 VDD.n530 VDD.n529 0.152939
R18503 VDD.n530 VDD.n405 0.152939
R18504 VDD.n538 VDD.n405 0.152939
R18505 VDD.n539 VDD.n538 0.152939
R18506 VDD.n540 VDD.n539 0.152939
R18507 VDD.n540 VDD.n403 0.152939
R18508 VDD.n548 VDD.n403 0.152939
R18509 VDD.n549 VDD.n548 0.152939
R18510 VDD.n550 VDD.n549 0.152939
R18511 VDD.n550 VDD.n401 0.152939
R18512 VDD.n558 VDD.n401 0.152939
R18513 VDD.n559 VDD.n558 0.152939
R18514 VDD.n560 VDD.n559 0.152939
R18515 VDD.n560 VDD.n399 0.152939
R18516 VDD.n568 VDD.n399 0.152939
R18517 VDD.n569 VDD.n568 0.152939
R18518 VDD.n570 VDD.n569 0.152939
R18519 VDD.n570 VDD.n397 0.152939
R18520 VDD.n578 VDD.n397 0.152939
R18521 VDD.n579 VDD.n578 0.152939
R18522 VDD.n580 VDD.n579 0.152939
R18523 VDD.n580 VDD.n395 0.152939
R18524 VDD.n587 VDD.n395 0.152939
R18525 VDD.n3343 VDD.n587 0.152939
R18526 VDD.n3221 VDD.n3220 0.152939
R18527 VDD.n3221 VDD.n645 0.152939
R18528 VDD.n3235 VDD.n645 0.152939
R18529 VDD.n3236 VDD.n3235 0.152939
R18530 VDD.n3237 VDD.n3236 0.152939
R18531 VDD.n3237 VDD.n634 0.152939
R18532 VDD.n3252 VDD.n634 0.152939
R18533 VDD.n3253 VDD.n3252 0.152939
R18534 VDD.n3254 VDD.n3253 0.152939
R18535 VDD.n3254 VDD.n622 0.152939
R18536 VDD.n3268 VDD.n622 0.152939
R18537 VDD.n3269 VDD.n3268 0.152939
R18538 VDD.n3270 VDD.n3269 0.152939
R18539 VDD.n3270 VDD.n611 0.152939
R18540 VDD.n3285 VDD.n611 0.152939
R18541 VDD.n3286 VDD.n3285 0.152939
R18542 VDD.n3287 VDD.n3286 0.152939
R18543 VDD.n3289 VDD.n3287 0.152939
R18544 VDD.n3289 VDD.n3288 0.152939
R18545 VDD.n3288 VDD.n600 0.152939
R18546 VDD.n600 VDD.n598 0.152939
R18547 VDD.n3307 VDD.n598 0.152939
R18548 VDD.n3308 VDD.n3307 0.152939
R18549 VDD.n3309 VDD.n3308 0.152939
R18550 VDD.n3309 VDD.n596 0.152939
R18551 VDD.n3314 VDD.n596 0.152939
R18552 VDD.n3315 VDD.n3314 0.152939
R18553 VDD.n3316 VDD.n3315 0.152939
R18554 VDD.n3316 VDD.n594 0.152939
R18555 VDD.n3321 VDD.n594 0.152939
R18556 VDD.n3322 VDD.n3321 0.152939
R18557 VDD.n3323 VDD.n3322 0.152939
R18558 VDD.n3323 VDD.n592 0.152939
R18559 VDD.n3328 VDD.n592 0.152939
R18560 VDD.n3329 VDD.n3328 0.152939
R18561 VDD.n3330 VDD.n3329 0.152939
R18562 VDD.n3330 VDD.n590 0.152939
R18563 VDD.n3335 VDD.n590 0.152939
R18564 VDD.n3336 VDD.n3335 0.152939
R18565 VDD.n3337 VDD.n3336 0.152939
R18566 VDD.n3337 VDD.n588 0.152939
R18567 VDD.n3342 VDD.n588 0.152939
R18568 VDD.n3081 VDD.n3080 0.152939
R18569 VDD.n3082 VDD.n3081 0.152939
R18570 VDD.n3083 VDD.n3082 0.152939
R18571 VDD.n3084 VDD.n3083 0.152939
R18572 VDD.n3085 VDD.n3084 0.152939
R18573 VDD.n3085 VDD.n657 0.152939
R18574 VDD.n3219 VDD.n657 0.152939
R18575 VDD.n2130 VDD.n1091 0.152939
R18576 VDD.n2126 VDD.n1091 0.152939
R18577 VDD.n2126 VDD.n2125 0.152939
R18578 VDD.n2125 VDD.n2124 0.152939
R18579 VDD.n2124 VDD.n1097 0.152939
R18580 VDD.n2120 VDD.n1097 0.152939
R18581 VDD.n2120 VDD.n2119 0.152939
R18582 VDD.n1466 VDD.n1230 0.152939
R18583 VDD.n1481 VDD.n1230 0.152939
R18584 VDD.n1482 VDD.n1481 0.152939
R18585 VDD.n1483 VDD.n1482 0.152939
R18586 VDD.n1483 VDD.n1218 0.152939
R18587 VDD.n1497 VDD.n1218 0.152939
R18588 VDD.n1498 VDD.n1497 0.152939
R18589 VDD.n1499 VDD.n1498 0.152939
R18590 VDD.n1499 VDD.n1206 0.152939
R18591 VDD.n1514 VDD.n1206 0.152939
R18592 VDD.n1515 VDD.n1514 0.152939
R18593 VDD.n1516 VDD.n1515 0.152939
R18594 VDD.n1516 VDD.n1195 0.152939
R18595 VDD.n1530 VDD.n1195 0.152939
R18596 VDD.n1531 VDD.n1530 0.152939
R18597 VDD.n1532 VDD.n1531 0.152939
R18598 VDD.n1532 VDD.n1183 0.152939
R18599 VDD.n1547 VDD.n1183 0.152939
R18600 VDD.n1548 VDD.n1547 0.152939
R18601 VDD.n1549 VDD.n1548 0.152939
R18602 VDD.n1549 VDD.n1172 0.152939
R18603 VDD.n1845 VDD.n1172 0.152939
R18604 VDD.n1846 VDD.n1845 0.152939
R18605 VDD.n1847 VDD.n1846 0.152939
R18606 VDD.n1847 VDD.n1159 0.152939
R18607 VDD.n1861 VDD.n1159 0.152939
R18608 VDD.n1862 VDD.n1861 0.152939
R18609 VDD.n1863 VDD.n1862 0.152939
R18610 VDD.n1863 VDD.n1148 0.152939
R18611 VDD.n1877 VDD.n1148 0.152939
R18612 VDD.n1878 VDD.n1877 0.152939
R18613 VDD.n1879 VDD.n1878 0.152939
R18614 VDD.n1879 VDD.n1135 0.152939
R18615 VDD.n1893 VDD.n1135 0.152939
R18616 VDD.n1894 VDD.n1893 0.152939
R18617 VDD.n1895 VDD.n1894 0.152939
R18618 VDD.n1895 VDD.n1124 0.152939
R18619 VDD.n1909 VDD.n1124 0.152939
R18620 VDD.n1910 VDD.n1909 0.152939
R18621 VDD.n1912 VDD.n1910 0.152939
R18622 VDD.n1912 VDD.n1911 0.152939
R18623 VDD.n1911 VDD.n1104 0.152939
R18624 VDD.n1312 VDD.n1235 0.152939
R18625 VDD.n1313 VDD.n1312 0.152939
R18626 VDD.n1314 VDD.n1313 0.152939
R18627 VDD.n1314 VDD.n1304 0.152939
R18628 VDD.n1322 VDD.n1304 0.152939
R18629 VDD.n1323 VDD.n1322 0.152939
R18630 VDD.n1324 VDD.n1323 0.152939
R18631 VDD.n1324 VDD.n1300 0.152939
R18632 VDD.n1332 VDD.n1300 0.152939
R18633 VDD.n1333 VDD.n1332 0.152939
R18634 VDD.n1334 VDD.n1333 0.152939
R18635 VDD.n1334 VDD.n1296 0.152939
R18636 VDD.n1342 VDD.n1296 0.152939
R18637 VDD.n1343 VDD.n1342 0.152939
R18638 VDD.n1346 VDD.n1343 0.152939
R18639 VDD.n1346 VDD.n1345 0.152939
R18640 VDD.n1345 VDD.n1344 0.152939
R18641 VDD.n1344 VDD.n1287 0.152939
R18642 VDD.n1356 VDD.n1287 0.152939
R18643 VDD.n1357 VDD.n1356 0.152939
R18644 VDD.n1358 VDD.n1357 0.152939
R18645 VDD.n1358 VDD.n1283 0.152939
R18646 VDD.n1366 VDD.n1283 0.152939
R18647 VDD.n1367 VDD.n1366 0.152939
R18648 VDD.n1368 VDD.n1367 0.152939
R18649 VDD.n1368 VDD.n1279 0.152939
R18650 VDD.n1376 VDD.n1279 0.152939
R18651 VDD.n1377 VDD.n1376 0.152939
R18652 VDD.n1378 VDD.n1377 0.152939
R18653 VDD.n1378 VDD.n1275 0.152939
R18654 VDD.n1386 VDD.n1275 0.152939
R18655 VDD.n1387 VDD.n1386 0.152939
R18656 VDD.n1388 VDD.n1387 0.152939
R18657 VDD.n1388 VDD.n1271 0.152939
R18658 VDD.n1396 VDD.n1271 0.152939
R18659 VDD.n1397 VDD.n1396 0.152939
R18660 VDD.n1400 VDD.n1397 0.152939
R18661 VDD.n1400 VDD.n1399 0.152939
R18662 VDD.n1399 VDD.n1398 0.152939
R18663 VDD.n1398 VDD.n1262 0.152939
R18664 VDD.n1410 VDD.n1262 0.152939
R18665 VDD.n1411 VDD.n1410 0.152939
R18666 VDD.n1412 VDD.n1411 0.152939
R18667 VDD.n1412 VDD.n1258 0.152939
R18668 VDD.n1420 VDD.n1258 0.152939
R18669 VDD.n1421 VDD.n1420 0.152939
R18670 VDD.n1422 VDD.n1421 0.152939
R18671 VDD.n1422 VDD.n1254 0.152939
R18672 VDD.n1430 VDD.n1254 0.152939
R18673 VDD.n1431 VDD.n1430 0.152939
R18674 VDD.n1432 VDD.n1431 0.152939
R18675 VDD.n1432 VDD.n1250 0.152939
R18676 VDD.n1440 VDD.n1250 0.152939
R18677 VDD.n1441 VDD.n1440 0.152939
R18678 VDD.n1442 VDD.n1441 0.152939
R18679 VDD.n1442 VDD.n1246 0.152939
R18680 VDD.n1450 VDD.n1246 0.152939
R18681 VDD.n1451 VDD.n1450 0.152939
R18682 VDD.n1454 VDD.n1451 0.152939
R18683 VDD.n1454 VDD.n1453 0.152939
R18684 VDD.n1453 VDD.n1452 0.152939
R18685 VDD.n1452 VDD.n1239 0.152939
R18686 VDD.n1465 VDD.n1239 0.152939
R18687 VDD.n1474 VDD.n1473 0.152939
R18688 VDD.n1475 VDD.n1474 0.152939
R18689 VDD.n1475 VDD.n1224 0.152939
R18690 VDD.n1489 VDD.n1224 0.152939
R18691 VDD.n1490 VDD.n1489 0.152939
R18692 VDD.n1491 VDD.n1490 0.152939
R18693 VDD.n1491 VDD.n1212 0.152939
R18694 VDD.n1506 VDD.n1212 0.152939
R18695 VDD.n1507 VDD.n1506 0.152939
R18696 VDD.n1508 VDD.n1507 0.152939
R18697 VDD.n1508 VDD.n1201 0.152939
R18698 VDD.n1522 VDD.n1201 0.152939
R18699 VDD.n1523 VDD.n1522 0.152939
R18700 VDD.n1524 VDD.n1523 0.152939
R18701 VDD.n1524 VDD.n1189 0.152939
R18702 VDD.n1539 VDD.n1189 0.152939
R18703 VDD.n1540 VDD.n1539 0.152939
R18704 VDD.n1541 VDD.n1540 0.152939
R18705 VDD.n1541 VDD.n1178 0.152939
R18706 VDD.n1555 VDD.n1178 0.152939
R18707 VDD.n1839 VDD.n1838 0.145814
R18708 VDD.n3392 VDD.n297 0.145814
R18709 VDD.n3392 VDD.n298 0.145814
R18710 VDD.n1838 VDD.n1555 0.145814
R18711 VDD.n1535 VDD.t117 0.136916
R18712 VDD.t113 VDD.n1162 0.136916
R18713 VDD.n3293 VDD.t97 0.136916
R18714 VDD.n3381 VDD.t110 0.136916
R18715 VDD.n2094 VDD.n1932 0.110256
R18716 VDD.n3027 VDD.n702 0.110256
R18717 VDD.n3080 VDD.n3079 0.110256
R18718 VDD.n2131 VDD.n2130 0.110256
R18719 VDD.n2094 VDD.n1934 0.0431829
R18720 VDD.n2131 VDD.n1088 0.0431829
R18721 VDD.n3027 VDD.n705 0.0431829
R18722 VDD.n3079 VDD.n742 0.0431829
R18723 VDD VDD.n15 0.00833333
R18724 a_n2686_8222.n171 a_n2686_8222.n157 756.745
R18725 a_n2686_8222.n191 a_n2686_8222.n177 756.745
R18726 a_n2686_8222.n96 a_n2686_8222.n82 756.745
R18727 a_n2686_8222.n115 a_n2686_8222.n101 756.745
R18728 a_n2686_8222.n133 a_n2686_8222.n119 756.745
R18729 a_n2686_8222.n152 a_n2686_8222.n138 756.745
R18730 a_n2686_8222.n58 a_n2686_8222.n44 756.745
R18731 a_n2686_8222.n78 a_n2686_8222.n64 756.745
R18732 a_n2686_8222.n172 a_n2686_8222.n171 585
R18733 a_n2686_8222.n170 a_n2686_8222.n169 585
R18734 a_n2686_8222.n160 a_n2686_8222.n159 585
R18735 a_n2686_8222.n166 a_n2686_8222.n165 585
R18736 a_n2686_8222.n164 a_n2686_8222.n163 585
R18737 a_n2686_8222.n1 a_n2686_8222.n0 585
R18738 a_n2686_8222.n29 a_n2686_8222.n162 585
R18739 a_n2686_8222.n192 a_n2686_8222.n191 585
R18740 a_n2686_8222.n190 a_n2686_8222.n189 585
R18741 a_n2686_8222.n180 a_n2686_8222.n179 585
R18742 a_n2686_8222.n186 a_n2686_8222.n185 585
R18743 a_n2686_8222.n184 a_n2686_8222.n183 585
R18744 a_n2686_8222.n3 a_n2686_8222.n2 585
R18745 a_n2686_8222.n31 a_n2686_8222.n182 585
R18746 a_n2686_8222.n97 a_n2686_8222.n96 585
R18747 a_n2686_8222.n95 a_n2686_8222.n94 585
R18748 a_n2686_8222.n85 a_n2686_8222.n84 585
R18749 a_n2686_8222.n91 a_n2686_8222.n90 585
R18750 a_n2686_8222.n89 a_n2686_8222.n88 585
R18751 a_n2686_8222.n5 a_n2686_8222.n4 585
R18752 a_n2686_8222.n33 a_n2686_8222.n87 585
R18753 a_n2686_8222.n116 a_n2686_8222.n115 585
R18754 a_n2686_8222.n114 a_n2686_8222.n113 585
R18755 a_n2686_8222.n104 a_n2686_8222.n103 585
R18756 a_n2686_8222.n110 a_n2686_8222.n109 585
R18757 a_n2686_8222.n108 a_n2686_8222.n107 585
R18758 a_n2686_8222.n7 a_n2686_8222.n6 585
R18759 a_n2686_8222.n35 a_n2686_8222.n106 585
R18760 a_n2686_8222.n134 a_n2686_8222.n133 585
R18761 a_n2686_8222.n132 a_n2686_8222.n131 585
R18762 a_n2686_8222.n122 a_n2686_8222.n121 585
R18763 a_n2686_8222.n128 a_n2686_8222.n127 585
R18764 a_n2686_8222.n126 a_n2686_8222.n125 585
R18765 a_n2686_8222.n9 a_n2686_8222.n8 585
R18766 a_n2686_8222.n37 a_n2686_8222.n124 585
R18767 a_n2686_8222.n153 a_n2686_8222.n152 585
R18768 a_n2686_8222.n151 a_n2686_8222.n150 585
R18769 a_n2686_8222.n141 a_n2686_8222.n140 585
R18770 a_n2686_8222.n147 a_n2686_8222.n146 585
R18771 a_n2686_8222.n145 a_n2686_8222.n144 585
R18772 a_n2686_8222.n11 a_n2686_8222.n10 585
R18773 a_n2686_8222.n39 a_n2686_8222.n143 585
R18774 a_n2686_8222.n59 a_n2686_8222.n58 585
R18775 a_n2686_8222.n57 a_n2686_8222.n56 585
R18776 a_n2686_8222.n47 a_n2686_8222.n46 585
R18777 a_n2686_8222.n53 a_n2686_8222.n52 585
R18778 a_n2686_8222.n51 a_n2686_8222.n50 585
R18779 a_n2686_8222.n13 a_n2686_8222.n12 585
R18780 a_n2686_8222.n41 a_n2686_8222.n49 585
R18781 a_n2686_8222.n79 a_n2686_8222.n78 585
R18782 a_n2686_8222.n77 a_n2686_8222.n76 585
R18783 a_n2686_8222.n67 a_n2686_8222.n66 585
R18784 a_n2686_8222.n73 a_n2686_8222.n72 585
R18785 a_n2686_8222.n71 a_n2686_8222.n70 585
R18786 a_n2686_8222.n15 a_n2686_8222.n14 585
R18787 a_n2686_8222.n43 a_n2686_8222.n69 585
R18788 a_n2686_8222.n171 a_n2686_8222.n170 171.744
R18789 a_n2686_8222.n170 a_n2686_8222.n159 171.744
R18790 a_n2686_8222.n165 a_n2686_8222.n159 171.744
R18791 a_n2686_8222.n165 a_n2686_8222.n164 171.744
R18792 a_n2686_8222.n164 a_n2686_8222.n0 171.744
R18793 a_n2686_8222.n162 a_n2686_8222.n0 171.744
R18794 a_n2686_8222.n191 a_n2686_8222.n190 171.744
R18795 a_n2686_8222.n190 a_n2686_8222.n179 171.744
R18796 a_n2686_8222.n185 a_n2686_8222.n179 171.744
R18797 a_n2686_8222.n185 a_n2686_8222.n184 171.744
R18798 a_n2686_8222.n184 a_n2686_8222.n2 171.744
R18799 a_n2686_8222.n182 a_n2686_8222.n2 171.744
R18800 a_n2686_8222.n96 a_n2686_8222.n95 171.744
R18801 a_n2686_8222.n95 a_n2686_8222.n84 171.744
R18802 a_n2686_8222.n90 a_n2686_8222.n84 171.744
R18803 a_n2686_8222.n90 a_n2686_8222.n89 171.744
R18804 a_n2686_8222.n89 a_n2686_8222.n4 171.744
R18805 a_n2686_8222.n87 a_n2686_8222.n4 171.744
R18806 a_n2686_8222.n115 a_n2686_8222.n114 171.744
R18807 a_n2686_8222.n114 a_n2686_8222.n103 171.744
R18808 a_n2686_8222.n109 a_n2686_8222.n103 171.744
R18809 a_n2686_8222.n109 a_n2686_8222.n108 171.744
R18810 a_n2686_8222.n108 a_n2686_8222.n6 171.744
R18811 a_n2686_8222.n106 a_n2686_8222.n6 171.744
R18812 a_n2686_8222.n133 a_n2686_8222.n132 171.744
R18813 a_n2686_8222.n132 a_n2686_8222.n121 171.744
R18814 a_n2686_8222.n127 a_n2686_8222.n121 171.744
R18815 a_n2686_8222.n127 a_n2686_8222.n126 171.744
R18816 a_n2686_8222.n126 a_n2686_8222.n8 171.744
R18817 a_n2686_8222.n124 a_n2686_8222.n8 171.744
R18818 a_n2686_8222.n152 a_n2686_8222.n151 171.744
R18819 a_n2686_8222.n151 a_n2686_8222.n140 171.744
R18820 a_n2686_8222.n146 a_n2686_8222.n140 171.744
R18821 a_n2686_8222.n146 a_n2686_8222.n145 171.744
R18822 a_n2686_8222.n145 a_n2686_8222.n10 171.744
R18823 a_n2686_8222.n143 a_n2686_8222.n10 171.744
R18824 a_n2686_8222.n58 a_n2686_8222.n57 171.744
R18825 a_n2686_8222.n57 a_n2686_8222.n46 171.744
R18826 a_n2686_8222.n52 a_n2686_8222.n46 171.744
R18827 a_n2686_8222.n52 a_n2686_8222.n51 171.744
R18828 a_n2686_8222.n51 a_n2686_8222.n12 171.744
R18829 a_n2686_8222.n49 a_n2686_8222.n12 171.744
R18830 a_n2686_8222.n78 a_n2686_8222.n77 171.744
R18831 a_n2686_8222.n77 a_n2686_8222.n66 171.744
R18832 a_n2686_8222.n72 a_n2686_8222.n66 171.744
R18833 a_n2686_8222.n72 a_n2686_8222.n71 171.744
R18834 a_n2686_8222.n71 a_n2686_8222.n14 171.744
R18835 a_n2686_8222.n69 a_n2686_8222.n14 171.744
R18836 a_n2686_8222.n162 a_n2686_8222.t11 85.8723
R18837 a_n2686_8222.n182 a_n2686_8222.t15 85.8723
R18838 a_n2686_8222.n87 a_n2686_8222.t16 85.8723
R18839 a_n2686_8222.n106 a_n2686_8222.t0 85.8723
R18840 a_n2686_8222.n124 a_n2686_8222.t14 85.8723
R18841 a_n2686_8222.n143 a_n2686_8222.t10 85.8723
R18842 a_n2686_8222.n49 a_n2686_8222.t20 85.8723
R18843 a_n2686_8222.n69 a_n2686_8222.t3 85.8723
R18844 a_n2686_8222.n17 a_n2686_8222.n175 81.2397
R18845 a_n2686_8222.n17 a_n2686_8222.n176 81.2397
R18846 a_n2686_8222.n26 a_n2686_8222.n100 81.2397
R18847 a_n2686_8222.n27 a_n2686_8222.n137 81.2397
R18848 a_n2686_8222.n16 a_n2686_8222.n62 81.2397
R18849 a_n2686_8222.n16 a_n2686_8222.n63 81.2397
R18850 a_n2686_8222.n17 a_n2686_8222.n174 38.3829
R18851 a_n2686_8222.n26 a_n2686_8222.n99 38.3829
R18852 a_n2686_8222.n16 a_n2686_8222.n61 38.3829
R18853 a_n2686_8222.n17 a_n2686_8222.n194 37.8096
R18854 a_n2686_8222.n26 a_n2686_8222.n118 37.8096
R18855 a_n2686_8222.n26 a_n2686_8222.n136 37.8096
R18856 a_n2686_8222.n27 a_n2686_8222.n155 37.8096
R18857 a_n2686_8222.n16 a_n2686_8222.n81 37.8096
R18858 a_n2686_8222.n29 a_n2686_8222.n28 5.3305
R18859 a_n2686_8222.n31 a_n2686_8222.n30 5.3305
R18860 a_n2686_8222.n33 a_n2686_8222.n32 5.3305
R18861 a_n2686_8222.n35 a_n2686_8222.n34 5.3305
R18862 a_n2686_8222.n37 a_n2686_8222.n36 5.3305
R18863 a_n2686_8222.n39 a_n2686_8222.n38 5.3305
R18864 a_n2686_8222.n41 a_n2686_8222.n40 5.3305
R18865 a_n2686_8222.n43 a_n2686_8222.n42 5.3305
R18866 a_n2686_8222.n29 a_n2686_8222.n1 12.8005
R18867 a_n2686_8222.n31 a_n2686_8222.n3 12.8005
R18868 a_n2686_8222.n33 a_n2686_8222.n5 12.8005
R18869 a_n2686_8222.n35 a_n2686_8222.n7 12.8005
R18870 a_n2686_8222.n37 a_n2686_8222.n9 12.8005
R18871 a_n2686_8222.n39 a_n2686_8222.n11 12.8005
R18872 a_n2686_8222.n41 a_n2686_8222.n13 12.8005
R18873 a_n2686_8222.n43 a_n2686_8222.n15 12.8005
R18874 a_n2686_8222.n163 a_n2686_8222.n1 12.0247
R18875 a_n2686_8222.n183 a_n2686_8222.n3 12.0247
R18876 a_n2686_8222.n88 a_n2686_8222.n5 12.0247
R18877 a_n2686_8222.n107 a_n2686_8222.n7 12.0247
R18878 a_n2686_8222.n125 a_n2686_8222.n9 12.0247
R18879 a_n2686_8222.n144 a_n2686_8222.n11 12.0247
R18880 a_n2686_8222.n50 a_n2686_8222.n13 12.0247
R18881 a_n2686_8222.n70 a_n2686_8222.n15 12.0247
R18882 a_n2686_8222.n166 a_n2686_8222.n161 11.249
R18883 a_n2686_8222.n186 a_n2686_8222.n181 11.249
R18884 a_n2686_8222.n91 a_n2686_8222.n86 11.249
R18885 a_n2686_8222.n110 a_n2686_8222.n105 11.249
R18886 a_n2686_8222.n128 a_n2686_8222.n123 11.249
R18887 a_n2686_8222.n147 a_n2686_8222.n142 11.249
R18888 a_n2686_8222.n53 a_n2686_8222.n48 11.249
R18889 a_n2686_8222.n73 a_n2686_8222.n68 11.249
R18890 a_n2686_8222.n167 a_n2686_8222.n160 10.4732
R18891 a_n2686_8222.n187 a_n2686_8222.n180 10.4732
R18892 a_n2686_8222.n92 a_n2686_8222.n85 10.4732
R18893 a_n2686_8222.n111 a_n2686_8222.n104 10.4732
R18894 a_n2686_8222.n129 a_n2686_8222.n122 10.4732
R18895 a_n2686_8222.n148 a_n2686_8222.n141 10.4732
R18896 a_n2686_8222.n54 a_n2686_8222.n47 10.4732
R18897 a_n2686_8222.n74 a_n2686_8222.n67 10.4732
R18898 a_n2686_8222.n169 a_n2686_8222.n168 9.69747
R18899 a_n2686_8222.n189 a_n2686_8222.n188 9.69747
R18900 a_n2686_8222.n94 a_n2686_8222.n93 9.69747
R18901 a_n2686_8222.n113 a_n2686_8222.n112 9.69747
R18902 a_n2686_8222.n131 a_n2686_8222.n130 9.69747
R18903 a_n2686_8222.n150 a_n2686_8222.n149 9.69747
R18904 a_n2686_8222.n56 a_n2686_8222.n55 9.69747
R18905 a_n2686_8222.n76 a_n2686_8222.n75 9.69747
R18906 a_n2686_8222.n174 a_n2686_8222.n18 9.45567
R18907 a_n2686_8222.n194 a_n2686_8222.n19 9.45567
R18908 a_n2686_8222.n99 a_n2686_8222.n20 9.45567
R18909 a_n2686_8222.n118 a_n2686_8222.n21 9.45567
R18910 a_n2686_8222.n136 a_n2686_8222.n22 9.45567
R18911 a_n2686_8222.n155 a_n2686_8222.n23 9.45567
R18912 a_n2686_8222.n61 a_n2686_8222.n24 9.45567
R18913 a_n2686_8222.n81 a_n2686_8222.n25 9.45567
R18914 a_n2686_8222.n18 a_n2686_8222.n173 9.3005
R18915 a_n2686_8222.n158 a_n2686_8222.n18 9.3005
R18916 a_n2686_8222.n168 a_n2686_8222.n18 9.3005
R18917 a_n2686_8222.n18 a_n2686_8222.n167 9.3005
R18918 a_n2686_8222.n161 a_n2686_8222.n18 9.3005
R18919 a_n2686_8222.n19 a_n2686_8222.n193 9.3005
R18920 a_n2686_8222.n178 a_n2686_8222.n19 9.3005
R18921 a_n2686_8222.n188 a_n2686_8222.n19 9.3005
R18922 a_n2686_8222.n19 a_n2686_8222.n187 9.3005
R18923 a_n2686_8222.n181 a_n2686_8222.n19 9.3005
R18924 a_n2686_8222.n20 a_n2686_8222.n98 9.3005
R18925 a_n2686_8222.n83 a_n2686_8222.n20 9.3005
R18926 a_n2686_8222.n93 a_n2686_8222.n20 9.3005
R18927 a_n2686_8222.n20 a_n2686_8222.n92 9.3005
R18928 a_n2686_8222.n86 a_n2686_8222.n20 9.3005
R18929 a_n2686_8222.n21 a_n2686_8222.n117 9.3005
R18930 a_n2686_8222.n102 a_n2686_8222.n21 9.3005
R18931 a_n2686_8222.n112 a_n2686_8222.n21 9.3005
R18932 a_n2686_8222.n21 a_n2686_8222.n111 9.3005
R18933 a_n2686_8222.n105 a_n2686_8222.n21 9.3005
R18934 a_n2686_8222.n22 a_n2686_8222.n135 9.3005
R18935 a_n2686_8222.n120 a_n2686_8222.n22 9.3005
R18936 a_n2686_8222.n130 a_n2686_8222.n22 9.3005
R18937 a_n2686_8222.n22 a_n2686_8222.n129 9.3005
R18938 a_n2686_8222.n123 a_n2686_8222.n22 9.3005
R18939 a_n2686_8222.n23 a_n2686_8222.n154 9.3005
R18940 a_n2686_8222.n139 a_n2686_8222.n23 9.3005
R18941 a_n2686_8222.n149 a_n2686_8222.n23 9.3005
R18942 a_n2686_8222.n23 a_n2686_8222.n148 9.3005
R18943 a_n2686_8222.n142 a_n2686_8222.n23 9.3005
R18944 a_n2686_8222.n24 a_n2686_8222.n60 9.3005
R18945 a_n2686_8222.n45 a_n2686_8222.n24 9.3005
R18946 a_n2686_8222.n55 a_n2686_8222.n24 9.3005
R18947 a_n2686_8222.n24 a_n2686_8222.n54 9.3005
R18948 a_n2686_8222.n48 a_n2686_8222.n24 9.3005
R18949 a_n2686_8222.n25 a_n2686_8222.n80 9.3005
R18950 a_n2686_8222.n65 a_n2686_8222.n25 9.3005
R18951 a_n2686_8222.n75 a_n2686_8222.n25 9.3005
R18952 a_n2686_8222.n25 a_n2686_8222.n74 9.3005
R18953 a_n2686_8222.n68 a_n2686_8222.n25 9.3005
R18954 a_n2686_8222.t8 a_n2686_8222.n195 9.17555
R18955 a_n2686_8222.n172 a_n2686_8222.n158 8.92171
R18956 a_n2686_8222.n192 a_n2686_8222.n178 8.92171
R18957 a_n2686_8222.n97 a_n2686_8222.n83 8.92171
R18958 a_n2686_8222.n116 a_n2686_8222.n102 8.92171
R18959 a_n2686_8222.n134 a_n2686_8222.n120 8.92171
R18960 a_n2686_8222.n153 a_n2686_8222.n139 8.92171
R18961 a_n2686_8222.n59 a_n2686_8222.n45 8.92171
R18962 a_n2686_8222.n79 a_n2686_8222.n65 8.92171
R18963 a_n2686_8222.n173 a_n2686_8222.n157 8.14595
R18964 a_n2686_8222.n193 a_n2686_8222.n177 8.14595
R18965 a_n2686_8222.n98 a_n2686_8222.n82 8.14595
R18966 a_n2686_8222.n117 a_n2686_8222.n101 8.14595
R18967 a_n2686_8222.n135 a_n2686_8222.n119 8.14595
R18968 a_n2686_8222.n154 a_n2686_8222.n138 8.14595
R18969 a_n2686_8222.n60 a_n2686_8222.n44 8.14595
R18970 a_n2686_8222.n80 a_n2686_8222.n64 8.14595
R18971 a_n2686_8222.n156 a_n2686_8222.n27 5.91753
R18972 a_n2686_8222.n174 a_n2686_8222.n157 5.81868
R18973 a_n2686_8222.n194 a_n2686_8222.n177 5.81868
R18974 a_n2686_8222.n99 a_n2686_8222.n82 5.81868
R18975 a_n2686_8222.n118 a_n2686_8222.n101 5.81868
R18976 a_n2686_8222.n136 a_n2686_8222.n119 5.81868
R18977 a_n2686_8222.n155 a_n2686_8222.n138 5.81868
R18978 a_n2686_8222.n61 a_n2686_8222.n44 5.81868
R18979 a_n2686_8222.n81 a_n2686_8222.n64 5.81868
R18980 a_n2686_8222.n175 a_n2686_8222.t2 5.418
R18981 a_n2686_8222.n175 a_n2686_8222.t17 5.418
R18982 a_n2686_8222.n176 a_n2686_8222.t18 5.418
R18983 a_n2686_8222.n176 a_n2686_8222.t19 5.418
R18984 a_n2686_8222.n100 a_n2686_8222.t7 5.418
R18985 a_n2686_8222.n100 a_n2686_8222.t5 5.418
R18986 a_n2686_8222.n137 a_n2686_8222.t9 5.418
R18987 a_n2686_8222.n137 a_n2686_8222.t13 5.418
R18988 a_n2686_8222.n62 a_n2686_8222.t12 5.418
R18989 a_n2686_8222.n62 a_n2686_8222.t6 5.418
R18990 a_n2686_8222.n63 a_n2686_8222.t1 5.418
R18991 a_n2686_8222.n63 a_n2686_8222.t4 5.418
R18992 a_n2686_8222.n173 a_n2686_8222.n172 5.04292
R18993 a_n2686_8222.n193 a_n2686_8222.n192 5.04292
R18994 a_n2686_8222.n98 a_n2686_8222.n97 5.04292
R18995 a_n2686_8222.n117 a_n2686_8222.n116 5.04292
R18996 a_n2686_8222.n135 a_n2686_8222.n134 5.04292
R18997 a_n2686_8222.n154 a_n2686_8222.n153 5.04292
R18998 a_n2686_8222.n60 a_n2686_8222.n59 5.04292
R18999 a_n2686_8222.n80 a_n2686_8222.n79 5.04292
R19000 a_n2686_8222.n169 a_n2686_8222.n158 4.26717
R19001 a_n2686_8222.n189 a_n2686_8222.n178 4.26717
R19002 a_n2686_8222.n94 a_n2686_8222.n83 4.26717
R19003 a_n2686_8222.n113 a_n2686_8222.n102 4.26717
R19004 a_n2686_8222.n131 a_n2686_8222.n120 4.26717
R19005 a_n2686_8222.n150 a_n2686_8222.n139 4.26717
R19006 a_n2686_8222.n56 a_n2686_8222.n45 4.26717
R19007 a_n2686_8222.n76 a_n2686_8222.n65 4.26717
R19008 a_n2686_8222.n195 a_n2686_8222.n156 4.20883
R19009 a_n2686_8222.n28 a_n2686_8222.t11 329.644
R19010 a_n2686_8222.n30 a_n2686_8222.t15 329.644
R19011 a_n2686_8222.n32 a_n2686_8222.t16 329.644
R19012 a_n2686_8222.n34 a_n2686_8222.t0 329.644
R19013 a_n2686_8222.n36 a_n2686_8222.t14 329.644
R19014 a_n2686_8222.n38 a_n2686_8222.t10 329.644
R19015 a_n2686_8222.n40 a_n2686_8222.t20 329.644
R19016 a_n2686_8222.n42 a_n2686_8222.t3 329.644
R19017 a_n2686_8222.n156 a_n2686_8222.n16 23.5201
R19018 a_n2686_8222.n15 a_n2686_8222.n25 10.4641
R19019 a_n2686_8222.n13 a_n2686_8222.n24 10.4641
R19020 a_n2686_8222.n11 a_n2686_8222.n23 10.4641
R19021 a_n2686_8222.n9 a_n2686_8222.n22 10.4641
R19022 a_n2686_8222.n7 a_n2686_8222.n21 10.4641
R19023 a_n2686_8222.n5 a_n2686_8222.n20 10.4641
R19024 a_n2686_8222.n3 a_n2686_8222.n19 10.4641
R19025 a_n2686_8222.n1 a_n2686_8222.n18 10.4641
R19026 a_n2686_8222.n195 a_n2686_8222.n17 6.8755
R19027 a_n2686_8222.n168 a_n2686_8222.n160 3.49141
R19028 a_n2686_8222.n188 a_n2686_8222.n180 3.49141
R19029 a_n2686_8222.n93 a_n2686_8222.n85 3.49141
R19030 a_n2686_8222.n112 a_n2686_8222.n104 3.49141
R19031 a_n2686_8222.n130 a_n2686_8222.n122 3.49141
R19032 a_n2686_8222.n149 a_n2686_8222.n141 3.49141
R19033 a_n2686_8222.n55 a_n2686_8222.n47 3.49141
R19034 a_n2686_8222.n75 a_n2686_8222.n67 3.49141
R19035 a_n2686_8222.n167 a_n2686_8222.n166 2.71565
R19036 a_n2686_8222.n187 a_n2686_8222.n186 2.71565
R19037 a_n2686_8222.n92 a_n2686_8222.n91 2.71565
R19038 a_n2686_8222.n111 a_n2686_8222.n110 2.71565
R19039 a_n2686_8222.n129 a_n2686_8222.n128 2.71565
R19040 a_n2686_8222.n148 a_n2686_8222.n147 2.71565
R19041 a_n2686_8222.n54 a_n2686_8222.n53 2.71565
R19042 a_n2686_8222.n74 a_n2686_8222.n73 2.71565
R19043 a_n2686_8222.n25 a_n2686_8222.n42 2.13947
R19044 a_n2686_8222.n24 a_n2686_8222.n40 2.13947
R19045 a_n2686_8222.n23 a_n2686_8222.n38 2.13947
R19046 a_n2686_8222.n22 a_n2686_8222.n36 2.13947
R19047 a_n2686_8222.n21 a_n2686_8222.n34 2.13947
R19048 a_n2686_8222.n20 a_n2686_8222.n32 2.13947
R19049 a_n2686_8222.n19 a_n2686_8222.n30 2.13947
R19050 a_n2686_8222.n18 a_n2686_8222.n28 2.13947
R19051 a_n2686_8222.n163 a_n2686_8222.n161 1.93989
R19052 a_n2686_8222.n183 a_n2686_8222.n181 1.93989
R19053 a_n2686_8222.n88 a_n2686_8222.n86 1.93989
R19054 a_n2686_8222.n107 a_n2686_8222.n105 1.93989
R19055 a_n2686_8222.n125 a_n2686_8222.n123 1.93989
R19056 a_n2686_8222.n144 a_n2686_8222.n142 1.93989
R19057 a_n2686_8222.n50 a_n2686_8222.n48 1.93989
R19058 a_n2686_8222.n70 a_n2686_8222.n68 1.93989
R19059 a_n2686_8222.n27 a_n2686_8222.n26 1.8755
R19060 a_n2686_12578.n118 a_n2686_12578.n98 756.745
R19061 a_n2686_12578.n89 a_n2686_12578.n69 756.745
R19062 a_n2686_12578.n166 a_n2686_12578.n146 756.745
R19063 a_n2686_12578.n195 a_n2686_12578.n175 756.745
R19064 a_n2686_12578.n119 a_n2686_12578.n118 585
R19065 a_n2686_12578.n117 a_n2686_12578.n116 585
R19066 a_n2686_12578.n101 a_n2686_12578.n100 585
R19067 a_n2686_12578.n113 a_n2686_12578.n112 585
R19068 a_n2686_12578.n111 a_n2686_12578.n110 585
R19069 a_n2686_12578.n104 a_n2686_12578.n103 585
R19070 a_n2686_12578.n107 a_n2686_12578.n106 585
R19071 a_n2686_12578.n90 a_n2686_12578.n89 585
R19072 a_n2686_12578.n88 a_n2686_12578.n87 585
R19073 a_n2686_12578.n72 a_n2686_12578.n71 585
R19074 a_n2686_12578.n84 a_n2686_12578.n83 585
R19075 a_n2686_12578.n82 a_n2686_12578.n81 585
R19076 a_n2686_12578.n75 a_n2686_12578.n74 585
R19077 a_n2686_12578.n78 a_n2686_12578.n77 585
R19078 a_n2686_12578.n167 a_n2686_12578.n166 585
R19079 a_n2686_12578.n165 a_n2686_12578.n164 585
R19080 a_n2686_12578.n149 a_n2686_12578.n148 585
R19081 a_n2686_12578.n161 a_n2686_12578.n160 585
R19082 a_n2686_12578.n159 a_n2686_12578.n158 585
R19083 a_n2686_12578.n152 a_n2686_12578.n151 585
R19084 a_n2686_12578.n155 a_n2686_12578.n154 585
R19085 a_n2686_12578.n196 a_n2686_12578.n195 585
R19086 a_n2686_12578.n194 a_n2686_12578.n193 585
R19087 a_n2686_12578.n178 a_n2686_12578.n177 585
R19088 a_n2686_12578.n190 a_n2686_12578.n189 585
R19089 a_n2686_12578.n188 a_n2686_12578.n187 585
R19090 a_n2686_12578.n181 a_n2686_12578.n180 585
R19091 a_n2686_12578.n184 a_n2686_12578.n183 585
R19092 a_n2686_12578.t24 a_n2686_12578.n105 327.601
R19093 a_n2686_12578.t6 a_n2686_12578.n76 327.601
R19094 a_n2686_12578.t18 a_n2686_12578.n153 327.601
R19095 a_n2686_12578.t10 a_n2686_12578.n182 327.601
R19096 a_n2686_12578.n144 a_n2686_12578.t9 183.883
R19097 a_n2686_12578.n136 a_n2686_12578.t17 183.883
R19098 a_n2686_12578.n228 a_n2686_12578.t38 183.883
R19099 a_n2686_12578.n233 a_n2686_12578.t57 183.883
R19100 a_n2686_12578.n220 a_n2686_12578.t58 183.883
R19101 a_n2686_12578.n225 a_n2686_12578.t49 183.883
R19102 a_n2686_12578.n212 a_n2686_12578.t43 183.883
R19103 a_n2686_12578.n217 a_n2686_12578.t52 183.883
R19104 a_n2686_12578.n204 a_n2686_12578.t46 183.883
R19105 a_n2686_12578.n209 a_n2686_12578.t55 183.883
R19106 a_n2686_12578.n10 a_n2686_12578.t5 206.089
R19107 a_n2686_12578.n8 a_n2686_12578.t34 206.089
R19108 a_n2686_12578.n12 a_n2686_12578.t50 206.089
R19109 a_n2686_12578.n118 a_n2686_12578.n117 171.744
R19110 a_n2686_12578.n117 a_n2686_12578.n100 171.744
R19111 a_n2686_12578.n112 a_n2686_12578.n100 171.744
R19112 a_n2686_12578.n112 a_n2686_12578.n111 171.744
R19113 a_n2686_12578.n111 a_n2686_12578.n103 171.744
R19114 a_n2686_12578.n106 a_n2686_12578.n103 171.744
R19115 a_n2686_12578.n89 a_n2686_12578.n88 171.744
R19116 a_n2686_12578.n88 a_n2686_12578.n71 171.744
R19117 a_n2686_12578.n83 a_n2686_12578.n71 171.744
R19118 a_n2686_12578.n83 a_n2686_12578.n82 171.744
R19119 a_n2686_12578.n82 a_n2686_12578.n74 171.744
R19120 a_n2686_12578.n77 a_n2686_12578.n74 171.744
R19121 a_n2686_12578.n166 a_n2686_12578.n165 171.744
R19122 a_n2686_12578.n165 a_n2686_12578.n148 171.744
R19123 a_n2686_12578.n160 a_n2686_12578.n148 171.744
R19124 a_n2686_12578.n160 a_n2686_12578.n159 171.744
R19125 a_n2686_12578.n159 a_n2686_12578.n151 171.744
R19126 a_n2686_12578.n154 a_n2686_12578.n151 171.744
R19127 a_n2686_12578.n195 a_n2686_12578.n194 171.744
R19128 a_n2686_12578.n194 a_n2686_12578.n177 171.744
R19129 a_n2686_12578.n189 a_n2686_12578.n177 171.744
R19130 a_n2686_12578.n189 a_n2686_12578.n188 171.744
R19131 a_n2686_12578.n188 a_n2686_12578.n180 171.744
R19132 a_n2686_12578.n183 a_n2686_12578.n180 171.744
R19133 a_n2686_12578.n17 a_n2686_12578.n5 68.6201
R19134 a_n2686_12578.n5 a_n2686_12578.n16 71.6402
R19135 a_n2686_12578.n132 a_n2686_12578.n7 161.3
R19136 a_n2686_12578.n7 a_n2686_12578.n15 68.6201
R19137 a_n2686_12578.n19 a_n2686_12578.n3 68.6201
R19138 a_n2686_12578.n3 a_n2686_12578.n18 71.6402
R19139 a_n2686_12578.n129 a_n2686_12578.n9 161.3
R19140 a_n2686_12578.n9 a_n2686_12578.n14 68.6201
R19141 a_n2686_12578.n21 a_n2686_12578.n0 68.6201
R19142 a_n2686_12578.n0 a_n2686_12578.n20 71.6402
R19143 a_n2686_12578.n237 a_n2686_12578.n11 161.3
R19144 a_n2686_12578.n11 a_n2686_12578.n13 68.6201
R19145 a_n2686_12578.n208 a_n2686_12578.n26 161.3
R19146 a_n2686_12578.n22 a_n2686_12578.n26 161.3
R19147 a_n2686_12578.n25 a_n2686_12578.n23 71.6402
R19148 a_n2686_12578.n205 a_n2686_12578.n24 161.3
R19149 a_n2686_12578.n216 a_n2686_12578.n31 161.3
R19150 a_n2686_12578.n27 a_n2686_12578.n31 161.3
R19151 a_n2686_12578.n30 a_n2686_12578.n28 71.6402
R19152 a_n2686_12578.n213 a_n2686_12578.n29 161.3
R19153 a_n2686_12578.n224 a_n2686_12578.n36 161.3
R19154 a_n2686_12578.n32 a_n2686_12578.n36 161.3
R19155 a_n2686_12578.n35 a_n2686_12578.n33 71.6402
R19156 a_n2686_12578.n221 a_n2686_12578.n34 161.3
R19157 a_n2686_12578.n232 a_n2686_12578.n41 161.3
R19158 a_n2686_12578.n37 a_n2686_12578.n41 161.3
R19159 a_n2686_12578.n40 a_n2686_12578.n38 71.6402
R19160 a_n2686_12578.n229 a_n2686_12578.n39 161.3
R19161 a_n2686_12578.n51 a_n2686_12578.n48 74.8341
R19162 a_n2686_12578.n49 a_n2686_12578.n46 68.6201
R19163 a_n2686_12578.n45 a_n2686_12578.n47 71.6402
R19164 a_n2686_12578.n138 a_n2686_12578.n42 161.3
R19165 a_n2686_12578.n140 a_n2686_12578.n42 161.3
R19166 a_n2686_12578.n44 a_n2686_12578.n141 161.3
R19167 a_n2686_12578.n142 a_n2686_12578.n44 161.3
R19168 a_n2686_12578.n143 a_n2686_12578.n43 161.3
R19169 a_n2686_12578.n134 a_n2686_12578.t21 144.601
R19170 a_n2686_12578.n139 a_n2686_12578.t15 144.601
R19171 a_n2686_12578.n137 a_n2686_12578.t1 144.601
R19172 a_n2686_12578.n135 a_n2686_12578.t19 144.601
R19173 a_n2686_12578.n230 a_n2686_12578.t51 144.601
R19174 a_n2686_12578.n231 a_n2686_12578.t41 144.601
R19175 a_n2686_12578.n222 a_n2686_12578.t40 144.601
R19176 a_n2686_12578.n223 a_n2686_12578.t37 144.601
R19177 a_n2686_12578.n214 a_n2686_12578.t32 144.601
R19178 a_n2686_12578.n215 a_n2686_12578.t36 144.601
R19179 a_n2686_12578.n206 a_n2686_12578.t35 144.601
R19180 a_n2686_12578.n207 a_n2686_12578.t44 144.601
R19181 a_n2686_12578.n126 a_n2686_12578.t7 144.601
R19182 a_n2686_12578.n130 a_n2686_12578.t11 144.601
R19183 a_n2686_12578.n128 a_n2686_12578.t3 144.601
R19184 a_n2686_12578.n127 a_n2686_12578.t13 144.601
R19185 a_n2686_12578.n124 a_n2686_12578.t39 144.601
R19186 a_n2686_12578.n133 a_n2686_12578.t45 144.601
R19187 a_n2686_12578.n131 a_n2686_12578.t33 144.601
R19188 a_n2686_12578.n125 a_n2686_12578.t42 144.601
R19189 a_n2686_12578.n67 a_n2686_12578.t59 144.601
R19190 a_n2686_12578.n238 a_n2686_12578.t56 144.601
R19191 a_n2686_12578.n236 a_n2686_12578.t47 144.601
R19192 a_n2686_12578.n68 a_n2686_12578.t54 144.601
R19193 a_n2686_12578.n106 a_n2686_12578.t24 85.8723
R19194 a_n2686_12578.n77 a_n2686_12578.t6 85.8723
R19195 a_n2686_12578.n154 a_n2686_12578.t18 85.8723
R19196 a_n2686_12578.n183 a_n2686_12578.t10 85.8723
R19197 a_n2686_12578.n241 a_n2686_12578.n240 84.3502
R19198 a_n2686_12578.n66 a_n2686_12578.n65 84.35
R19199 a_n2686_12578.n66 a_n2686_12578.n64 84.35
R19200 a_n2686_12578.n243 a_n2686_12578.n242 84.0635
R19201 a_n2686_12578.n97 a_n2686_12578.n96 81.2397
R19202 a_n2686_12578.n95 a_n2686_12578.n94 81.2397
R19203 a_n2686_12578.n172 a_n2686_12578.n171 81.2397
R19204 a_n2686_12578.n174 a_n2686_12578.n173 81.2397
R19205 a_n2686_12578.n6 a_n2686_12578.n5 28.1161
R19206 a_n2686_12578.n7 a_n2686_12578.n8 28.1161
R19207 a_n2686_12578.n4 a_n2686_12578.n3 28.1161
R19208 a_n2686_12578.n9 a_n2686_12578.n10 28.1161
R19209 a_n2686_12578.n1 a_n2686_12578.n0 28.1161
R19210 a_n2686_12578.n11 a_n2686_12578.n12 28.1161
R19211 a_n2686_12578.n210 a_n2686_12578.n209 80.6037
R19212 a_n2686_12578.n204 a_n2686_12578.n203 80.6037
R19213 a_n2686_12578.n218 a_n2686_12578.n217 80.6037
R19214 a_n2686_12578.n212 a_n2686_12578.n211 80.6037
R19215 a_n2686_12578.n226 a_n2686_12578.n225 80.6037
R19216 a_n2686_12578.n220 a_n2686_12578.n219 80.6037
R19217 a_n2686_12578.n234 a_n2686_12578.n233 80.6037
R19218 a_n2686_12578.n228 a_n2686_12578.n227 80.6037
R19219 a_n2686_12578.n136 a_n2686_12578.n50 80.6037
R19220 a_n2686_12578.n145 a_n2686_12578.n144 80.6037
R19221 a_n2686_12578.n141 a_n2686_12578.n140 56.5617
R19222 a_n2686_12578.n49 a_n2686_12578.n135 48.4088
R19223 a_n2686_12578.n19 a_n2686_12578.n127 48.4088
R19224 a_n2686_12578.n17 a_n2686_12578.n125 48.4088
R19225 a_n2686_12578.n21 a_n2686_12578.n68 48.4088
R19226 a_n2686_12578.n229 a_n2686_12578.n228 56.3158
R19227 a_n2686_12578.n233 a_n2686_12578.n232 56.3158
R19228 a_n2686_12578.n221 a_n2686_12578.n220 56.3158
R19229 a_n2686_12578.n225 a_n2686_12578.n224 56.3158
R19230 a_n2686_12578.n213 a_n2686_12578.n212 56.3158
R19231 a_n2686_12578.n217 a_n2686_12578.n216 56.3158
R19232 a_n2686_12578.n205 a_n2686_12578.n204 56.3158
R19233 a_n2686_12578.n209 a_n2686_12578.n208 56.3158
R19234 a_n2686_12578.n144 a_n2686_12578.n143 47.4702
R19235 a_n2686_12578.n138 a_n2686_12578.n47 58.5991
R19236 a_n2686_12578.n137 a_n2686_12578.n47 26.1378
R19237 a_n2686_12578.n38 a_n2686_12578.n37 58.5991
R19238 a_n2686_12578.n33 a_n2686_12578.n32 58.5991
R19239 a_n2686_12578.n28 a_n2686_12578.n27 58.5991
R19240 a_n2686_12578.n23 a_n2686_12578.n22 58.5991
R19241 a_n2686_12578.n129 a_n2686_12578.n18 58.5991
R19242 a_n2686_12578.n128 a_n2686_12578.n18 26.1378
R19243 a_n2686_12578.n132 a_n2686_12578.n16 58.5991
R19244 a_n2686_12578.n131 a_n2686_12578.n16 26.1378
R19245 a_n2686_12578.n237 a_n2686_12578.n20 58.5991
R19246 a_n2686_12578.n236 a_n2686_12578.n20 26.1378
R19247 a_n2686_12578.n95 a_n2686_12578.n93 38.3829
R19248 a_n2686_12578.n172 a_n2686_12578.n170 38.3829
R19249 a_n2686_12578.n123 a_n2686_12578.n122 37.8096
R19250 a_n2686_12578.n200 a_n2686_12578.n199 37.8096
R19251 a_n2686_12578.n242 a_n2686_12578.n66 29.8404
R19252 a_n2686_12578.n143 a_n2686_12578.n142 25.0767
R19253 a_n2686_12578.n51 a_n2686_12578.n136 59.1045
R19254 a_n2686_12578.n10 a_n2686_12578.n126 32.4972
R19255 a_n2686_12578.n4 a_n2686_12578.t23 206.089
R19256 a_n2686_12578.n8 a_n2686_12578.n124 32.4972
R19257 a_n2686_12578.n6 a_n2686_12578.t48 206.089
R19258 a_n2686_12578.n12 a_n2686_12578.n67 32.4972
R19259 a_n2686_12578.n1 a_n2686_12578.t53 206.089
R19260 a_n2686_12578.n141 a_n2686_12578.n134 24.3464
R19261 a_n2686_12578.n14 a_n2686_12578.n126 48.4088
R19262 a_n2686_12578.n15 a_n2686_12578.n124 48.4088
R19263 a_n2686_12578.n13 a_n2686_12578.n67 48.4088
R19264 a_n2686_12578.n241 a_n2686_12578.n239 23.9442
R19265 a_n2686_12578.n140 a_n2686_12578.n139 16.477
R19266 a_n2686_12578.n137 a_n2686_12578.n49 40.5394
R19267 a_n2686_12578.n230 a_n2686_12578.n229 16.477
R19268 a_n2686_12578.n232 a_n2686_12578.n231 16.477
R19269 a_n2686_12578.n222 a_n2686_12578.n221 16.477
R19270 a_n2686_12578.n224 a_n2686_12578.n223 16.477
R19271 a_n2686_12578.n214 a_n2686_12578.n213 16.477
R19272 a_n2686_12578.n216 a_n2686_12578.n215 16.477
R19273 a_n2686_12578.n206 a_n2686_12578.n205 16.477
R19274 a_n2686_12578.n208 a_n2686_12578.n207 16.477
R19275 a_n2686_12578.n14 a_n2686_12578.n130 40.5394
R19276 a_n2686_12578.n128 a_n2686_12578.n19 40.5394
R19277 a_n2686_12578.n15 a_n2686_12578.n133 40.5394
R19278 a_n2686_12578.n131 a_n2686_12578.n17 40.5394
R19279 a_n2686_12578.n13 a_n2686_12578.n238 40.5394
R19280 a_n2686_12578.n236 a_n2686_12578.n21 40.5394
R19281 a_n2686_12578.n107 a_n2686_12578.n105 16.3865
R19282 a_n2686_12578.n78 a_n2686_12578.n76 16.3865
R19283 a_n2686_12578.n155 a_n2686_12578.n153 16.3865
R19284 a_n2686_12578.n184 a_n2686_12578.n182 16.3865
R19285 a_n2686_12578.n108 a_n2686_12578.n104 12.8005
R19286 a_n2686_12578.n79 a_n2686_12578.n75 12.8005
R19287 a_n2686_12578.n156 a_n2686_12578.n152 12.8005
R19288 a_n2686_12578.n185 a_n2686_12578.n181 12.8005
R19289 a_n2686_12578.n110 a_n2686_12578.n109 12.0247
R19290 a_n2686_12578.n81 a_n2686_12578.n80 12.0247
R19291 a_n2686_12578.n158 a_n2686_12578.n157 12.0247
R19292 a_n2686_12578.n187 a_n2686_12578.n186 12.0247
R19293 a_n2686_12578.n113 a_n2686_12578.n102 11.249
R19294 a_n2686_12578.n84 a_n2686_12578.n73 11.249
R19295 a_n2686_12578.n161 a_n2686_12578.n150 11.249
R19296 a_n2686_12578.n190 a_n2686_12578.n179 11.249
R19297 a_n2686_12578.n202 a_n2686_12578.n7 10.8153
R19298 a_n2686_12578.n0 a_n2686_12578.n235 10.6108
R19299 a_n2686_12578.n114 a_n2686_12578.n101 10.4732
R19300 a_n2686_12578.n85 a_n2686_12578.n72 10.4732
R19301 a_n2686_12578.n162 a_n2686_12578.n149 10.4732
R19302 a_n2686_12578.n191 a_n2686_12578.n178 10.4732
R19303 a_n2686_12578.n116 a_n2686_12578.n115 9.69747
R19304 a_n2686_12578.n87 a_n2686_12578.n86 9.69747
R19305 a_n2686_12578.n164 a_n2686_12578.n163 9.69747
R19306 a_n2686_12578.n193 a_n2686_12578.n192 9.69747
R19307 a_n2686_12578.n122 a_n2686_12578.n121 9.45567
R19308 a_n2686_12578.n93 a_n2686_12578.n92 9.45567
R19309 a_n2686_12578.n170 a_n2686_12578.n169 9.45567
R19310 a_n2686_12578.n199 a_n2686_12578.n198 9.45567
R19311 a_n2686_12578.n201 a_n2686_12578.n145 9.30587
R19312 a_n2686_12578.n121 a_n2686_12578.n120 9.3005
R19313 a_n2686_12578.n99 a_n2686_12578.n53 9.3005
R19314 a_n2686_12578.n115 a_n2686_12578.n53 9.3005
R19315 a_n2686_12578.n52 a_n2686_12578.n114 9.3005
R19316 a_n2686_12578.n102 a_n2686_12578.n52 9.3005
R19317 a_n2686_12578.n109 a_n2686_12578.n54 9.3005
R19318 a_n2686_12578.n54 a_n2686_12578.n108 9.3005
R19319 a_n2686_12578.n92 a_n2686_12578.n91 9.3005
R19320 a_n2686_12578.n70 a_n2686_12578.n56 9.3005
R19321 a_n2686_12578.n86 a_n2686_12578.n56 9.3005
R19322 a_n2686_12578.n55 a_n2686_12578.n85 9.3005
R19323 a_n2686_12578.n73 a_n2686_12578.n55 9.3005
R19324 a_n2686_12578.n80 a_n2686_12578.n57 9.3005
R19325 a_n2686_12578.n57 a_n2686_12578.n79 9.3005
R19326 a_n2686_12578.n169 a_n2686_12578.n168 9.3005
R19327 a_n2686_12578.n147 a_n2686_12578.n59 9.3005
R19328 a_n2686_12578.n163 a_n2686_12578.n59 9.3005
R19329 a_n2686_12578.n58 a_n2686_12578.n162 9.3005
R19330 a_n2686_12578.n150 a_n2686_12578.n58 9.3005
R19331 a_n2686_12578.n157 a_n2686_12578.n60 9.3005
R19332 a_n2686_12578.n60 a_n2686_12578.n156 9.3005
R19333 a_n2686_12578.n198 a_n2686_12578.n197 9.3005
R19334 a_n2686_12578.n176 a_n2686_12578.n62 9.3005
R19335 a_n2686_12578.n192 a_n2686_12578.n62 9.3005
R19336 a_n2686_12578.n61 a_n2686_12578.n191 9.3005
R19337 a_n2686_12578.n179 a_n2686_12578.n61 9.3005
R19338 a_n2686_12578.n186 a_n2686_12578.n63 9.3005
R19339 a_n2686_12578.n63 a_n2686_12578.n185 9.3005
R19340 a_n2686_12578.n119 a_n2686_12578.n99 8.92171
R19341 a_n2686_12578.n90 a_n2686_12578.n70 8.92171
R19342 a_n2686_12578.n167 a_n2686_12578.n147 8.92171
R19343 a_n2686_12578.n196 a_n2686_12578.n176 8.92171
R19344 a_n2686_12578.n2 a_n2686_12578.n123 8.2571
R19345 a_n2686_12578.n120 a_n2686_12578.n98 8.14595
R19346 a_n2686_12578.n91 a_n2686_12578.n69 8.14595
R19347 a_n2686_12578.n168 a_n2686_12578.n146 8.14595
R19348 a_n2686_12578.n197 a_n2686_12578.n175 8.14595
R19349 a_n2686_12578.n139 a_n2686_12578.n138 8.11581
R19350 a_n2686_12578.n38 a_n2686_12578.n230 26.1378
R19351 a_n2686_12578.n231 a_n2686_12578.n37 8.11581
R19352 a_n2686_12578.n33 a_n2686_12578.n222 26.1378
R19353 a_n2686_12578.n223 a_n2686_12578.n32 8.11581
R19354 a_n2686_12578.n28 a_n2686_12578.n214 26.1378
R19355 a_n2686_12578.n215 a_n2686_12578.n27 8.11581
R19356 a_n2686_12578.n23 a_n2686_12578.n206 26.1378
R19357 a_n2686_12578.n207 a_n2686_12578.n22 8.11581
R19358 a_n2686_12578.n130 a_n2686_12578.n129 8.11581
R19359 a_n2686_12578.n133 a_n2686_12578.n132 8.11581
R19360 a_n2686_12578.n238 a_n2686_12578.n237 8.11581
R19361 a_n2686_12578.n235 a_n2686_12578.n234 7.00284
R19362 a_n2686_12578.n203 a_n2686_12578.n202 7.00284
R19363 a_n2686_12578.n3 a_n2686_12578.n2 6.60701
R19364 a_n2686_12578.n122 a_n2686_12578.n98 5.81868
R19365 a_n2686_12578.n93 a_n2686_12578.n69 5.81868
R19366 a_n2686_12578.n170 a_n2686_12578.n146 5.81868
R19367 a_n2686_12578.n199 a_n2686_12578.n175 5.81868
R19368 a_n2686_12578.n201 a_n2686_12578.n200 5.55007
R19369 a_n2686_12578.n96 a_n2686_12578.t4 5.418
R19370 a_n2686_12578.n96 a_n2686_12578.t14 5.418
R19371 a_n2686_12578.n94 a_n2686_12578.t8 5.418
R19372 a_n2686_12578.n94 a_n2686_12578.t12 5.418
R19373 a_n2686_12578.n171 a_n2686_12578.t2 5.418
R19374 a_n2686_12578.n171 a_n2686_12578.t20 5.418
R19375 a_n2686_12578.n173 a_n2686_12578.t22 5.418
R19376 a_n2686_12578.n173 a_n2686_12578.t16 5.418
R19377 a_n2686_12578.n120 a_n2686_12578.n119 5.04292
R19378 a_n2686_12578.n91 a_n2686_12578.n90 5.04292
R19379 a_n2686_12578.n168 a_n2686_12578.n167 5.04292
R19380 a_n2686_12578.n197 a_n2686_12578.n196 5.04292
R19381 a_n2686_12578.n5 a_n2686_12578.n9 4.52033
R19382 a_n2686_12578.n116 a_n2686_12578.n99 4.26717
R19383 a_n2686_12578.n87 a_n2686_12578.n70 4.26717
R19384 a_n2686_12578.n164 a_n2686_12578.n147 4.26717
R19385 a_n2686_12578.n193 a_n2686_12578.n176 4.26717
R19386 a_n2686_12578.n235 a_n2686_12578.n2 4.20883
R19387 a_n2686_12578.n54 a_n2686_12578.n105 3.71286
R19388 a_n2686_12578.n57 a_n2686_12578.n76 3.71286
R19389 a_n2686_12578.n60 a_n2686_12578.n153 3.71286
R19390 a_n2686_12578.n63 a_n2686_12578.n182 3.71286
R19391 a_n2686_12578.n115 a_n2686_12578.n101 3.49141
R19392 a_n2686_12578.n86 a_n2686_12578.n72 3.49141
R19393 a_n2686_12578.n163 a_n2686_12578.n149 3.49141
R19394 a_n2686_12578.n192 a_n2686_12578.n178 3.49141
R19395 a_n2686_12578.n239 a_n2686_12578.n11 3.45549
R19396 a_n2686_12578.n240 a_n2686_12578.t31 3.3005
R19397 a_n2686_12578.n240 a_n2686_12578.t30 3.3005
R19398 a_n2686_12578.n65 a_n2686_12578.t26 3.3005
R19399 a_n2686_12578.n65 a_n2686_12578.t29 3.3005
R19400 a_n2686_12578.n64 a_n2686_12578.t25 3.3005
R19401 a_n2686_12578.n64 a_n2686_12578.t28 3.3005
R19402 a_n2686_12578.n243 a_n2686_12578.t27 3.3005
R19403 a_n2686_12578.t0 a_n2686_12578.n243 3.3005
R19404 a_n2686_12578.n114 a_n2686_12578.n113 2.71565
R19405 a_n2686_12578.n85 a_n2686_12578.n84 2.71565
R19406 a_n2686_12578.n162 a_n2686_12578.n161 2.71565
R19407 a_n2686_12578.n191 a_n2686_12578.n190 2.71565
R19408 a_n2686_12578.n110 a_n2686_12578.n102 1.93989
R19409 a_n2686_12578.n81 a_n2686_12578.n73 1.93989
R19410 a_n2686_12578.n158 a_n2686_12578.n150 1.93989
R19411 a_n2686_12578.n187 a_n2686_12578.n179 1.93989
R19412 a_n2686_12578.n219 a_n2686_12578.n218 1.42563
R19413 a_n2686_12578.n202 a_n2686_12578.n201 1.30542
R19414 a_n2686_12578.n109 a_n2686_12578.n104 1.16414
R19415 a_n2686_12578.n80 a_n2686_12578.n75 1.16414
R19416 a_n2686_12578.n157 a_n2686_12578.n152 1.16414
R19417 a_n2686_12578.n186 a_n2686_12578.n181 1.16414
R19418 a_n2686_12578.n239 a_n2686_12578.n50 1.02746
R19419 a_n2686_12578.n211 a_n2686_12578.n210 0.96351
R19420 a_n2686_12578.n227 a_n2686_12578.n226 0.96351
R19421 a_n2686_12578.n97 a_n2686_12578.n95 0.573776
R19422 a_n2686_12578.n123 a_n2686_12578.n97 0.573776
R19423 a_n2686_12578.n200 a_n2686_12578.n174 0.573776
R19424 a_n2686_12578.n174 a_n2686_12578.n172 0.573776
R19425 a_n2686_12578.n108 a_n2686_12578.n107 0.388379
R19426 a_n2686_12578.n79 a_n2686_12578.n78 0.388379
R19427 a_n2686_12578.n156 a_n2686_12578.n155 0.388379
R19428 a_n2686_12578.n185 a_n2686_12578.n184 0.388379
R19429 a_n2686_12578.n46 a_n2686_12578.n48 0.379288
R19430 a_n2686_12578.n63 a_n2686_12578.n61 0.310845
R19431 a_n2686_12578.n62 a_n2686_12578.n61 0.310845
R19432 a_n2686_12578.n198 a_n2686_12578.n62 0.310845
R19433 a_n2686_12578.n60 a_n2686_12578.n58 0.310845
R19434 a_n2686_12578.n59 a_n2686_12578.n58 0.310845
R19435 a_n2686_12578.n169 a_n2686_12578.n59 0.310845
R19436 a_n2686_12578.n57 a_n2686_12578.n55 0.310845
R19437 a_n2686_12578.n56 a_n2686_12578.n55 0.310845
R19438 a_n2686_12578.n92 a_n2686_12578.n56 0.310845
R19439 a_n2686_12578.n54 a_n2686_12578.n52 0.310845
R19440 a_n2686_12578.n53 a_n2686_12578.n52 0.310845
R19441 a_n2686_12578.n121 a_n2686_12578.n53 0.310845
R19442 a_n2686_12578.n242 a_n2686_12578.n241 0.287138
R19443 a_n2686_12578.n203 a_n2686_12578.n24 0.285035
R19444 a_n2686_12578.n210 a_n2686_12578.n26 0.285035
R19445 a_n2686_12578.n211 a_n2686_12578.n29 0.285035
R19446 a_n2686_12578.n218 a_n2686_12578.n31 0.285035
R19447 a_n2686_12578.n219 a_n2686_12578.n34 0.285035
R19448 a_n2686_12578.n226 a_n2686_12578.n36 0.285035
R19449 a_n2686_12578.n227 a_n2686_12578.n39 0.285035
R19450 a_n2686_12578.n234 a_n2686_12578.n41 0.285035
R19451 a_n2686_12578.n145 a_n2686_12578.n43 0.285035
R19452 a_n2686_12578.n48 a_n2686_12578.n50 0.285035
R19453 a_n2686_12578.n142 a_n2686_12578.n134 0.246418
R19454 a_n2686_12578.n51 a_n2686_12578.n135 11.8807
R19455 a_n2686_12578.n45 a_n2686_12578.n46 0.379288
R19456 a_n2686_12578.n42 a_n2686_12578.n45 0.379288
R19457 a_n2686_12578.n44 a_n2686_12578.n42 0.379288
R19458 a_n2686_12578.n44 a_n2686_12578.n43 0.379288
R19459 a_n2686_12578.n41 a_n2686_12578.n40 0.379288
R19460 a_n2686_12578.n40 a_n2686_12578.n39 0.379288
R19461 a_n2686_12578.n36 a_n2686_12578.n35 0.379288
R19462 a_n2686_12578.n35 a_n2686_12578.n34 0.379288
R19463 a_n2686_12578.n31 a_n2686_12578.n30 0.379288
R19464 a_n2686_12578.n30 a_n2686_12578.n29 0.379288
R19465 a_n2686_12578.n26 a_n2686_12578.n25 0.379288
R19466 a_n2686_12578.n25 a_n2686_12578.n24 0.379288
R19467 a_n2686_12578.n4 a_n2686_12578.n127 32.4972
R19468 a_n2686_12578.n6 a_n2686_12578.n125 32.4972
R19469 a_n2686_12578.n1 a_n2686_12578.n68 32.4972
R19470 a_n2686_12578.n7 a_n2686_12578.n5 2.46351
R19471 a_n2686_12578.n9 a_n2686_12578.n3 2.46351
R19472 a_n2686_12578.n11 a_n2686_12578.n0 2.46351
R19473 a_n2511_10356.n130 a_n2511_10356.n104 756.745
R19474 a_n2511_10356.n96 a_n2511_10356.n70 756.745
R19475 a_n2511_10356.n64 a_n2511_10356.n38 756.745
R19476 a_n2511_10356.n31 a_n2511_10356.n5 756.745
R19477 a_n2511_10356.n131 a_n2511_10356.n130 585
R19478 a_n2511_10356.n129 a_n2511_10356.n128 585
R19479 a_n2511_10356.n108 a_n2511_10356.n107 585
R19480 a_n2511_10356.n123 a_n2511_10356.n122 585
R19481 a_n2511_10356.n121 a_n2511_10356.n120 585
R19482 a_n2511_10356.n112 a_n2511_10356.n111 585
R19483 a_n2511_10356.n115 a_n2511_10356.n114 585
R19484 a_n2511_10356.n97 a_n2511_10356.n96 585
R19485 a_n2511_10356.n95 a_n2511_10356.n94 585
R19486 a_n2511_10356.n74 a_n2511_10356.n73 585
R19487 a_n2511_10356.n89 a_n2511_10356.n88 585
R19488 a_n2511_10356.n87 a_n2511_10356.n86 585
R19489 a_n2511_10356.n78 a_n2511_10356.n77 585
R19490 a_n2511_10356.n81 a_n2511_10356.n80 585
R19491 a_n2511_10356.n65 a_n2511_10356.n64 585
R19492 a_n2511_10356.n63 a_n2511_10356.n62 585
R19493 a_n2511_10356.n42 a_n2511_10356.n41 585
R19494 a_n2511_10356.n57 a_n2511_10356.n56 585
R19495 a_n2511_10356.n55 a_n2511_10356.n54 585
R19496 a_n2511_10356.n46 a_n2511_10356.n45 585
R19497 a_n2511_10356.n49 a_n2511_10356.n48 585
R19498 a_n2511_10356.n32 a_n2511_10356.n31 585
R19499 a_n2511_10356.n30 a_n2511_10356.n29 585
R19500 a_n2511_10356.n9 a_n2511_10356.n8 585
R19501 a_n2511_10356.n24 a_n2511_10356.n23 585
R19502 a_n2511_10356.n22 a_n2511_10356.n21 585
R19503 a_n2511_10356.n13 a_n2511_10356.n12 585
R19504 a_n2511_10356.n16 a_n2511_10356.n15 585
R19505 a_n2511_10356.t1 a_n2511_10356.n113 327.601
R19506 a_n2511_10356.t6 a_n2511_10356.n79 327.601
R19507 a_n2511_10356.t3 a_n2511_10356.n47 327.601
R19508 a_n2511_10356.t0 a_n2511_10356.n14 327.601
R19509 a_n2511_10356.n130 a_n2511_10356.n129 171.744
R19510 a_n2511_10356.n129 a_n2511_10356.n107 171.744
R19511 a_n2511_10356.n122 a_n2511_10356.n107 171.744
R19512 a_n2511_10356.n122 a_n2511_10356.n121 171.744
R19513 a_n2511_10356.n121 a_n2511_10356.n111 171.744
R19514 a_n2511_10356.n114 a_n2511_10356.n111 171.744
R19515 a_n2511_10356.n96 a_n2511_10356.n95 171.744
R19516 a_n2511_10356.n95 a_n2511_10356.n73 171.744
R19517 a_n2511_10356.n88 a_n2511_10356.n73 171.744
R19518 a_n2511_10356.n88 a_n2511_10356.n87 171.744
R19519 a_n2511_10356.n87 a_n2511_10356.n77 171.744
R19520 a_n2511_10356.n80 a_n2511_10356.n77 171.744
R19521 a_n2511_10356.n64 a_n2511_10356.n63 171.744
R19522 a_n2511_10356.n63 a_n2511_10356.n41 171.744
R19523 a_n2511_10356.n56 a_n2511_10356.n41 171.744
R19524 a_n2511_10356.n56 a_n2511_10356.n55 171.744
R19525 a_n2511_10356.n55 a_n2511_10356.n45 171.744
R19526 a_n2511_10356.n48 a_n2511_10356.n45 171.744
R19527 a_n2511_10356.n31 a_n2511_10356.n30 171.744
R19528 a_n2511_10356.n30 a_n2511_10356.n8 171.744
R19529 a_n2511_10356.n23 a_n2511_10356.n8 171.744
R19530 a_n2511_10356.n23 a_n2511_10356.n22 171.744
R19531 a_n2511_10356.n22 a_n2511_10356.n12 171.744
R19532 a_n2511_10356.n15 a_n2511_10356.n12 171.744
R19533 a_n2511_10356.n141 a_n2511_10356.n140 109.74
R19534 a_n2511_10356.n2 a_n2511_10356.n0 109.401
R19535 a_n2511_10356.n140 a_n2511_10356.n139 109.166
R19536 a_n2511_10356.n4 a_n2511_10356.n3 109.166
R19537 a_n2511_10356.n2 a_n2511_10356.n1 109.166
R19538 a_n2511_10356.n138 a_n2511_10356.n137 109.166
R19539 a_n2511_10356.n114 a_n2511_10356.t1 85.8723
R19540 a_n2511_10356.n80 a_n2511_10356.t6 85.8723
R19541 a_n2511_10356.n48 a_n2511_10356.t3 85.8723
R19542 a_n2511_10356.n15 a_n2511_10356.t0 85.8723
R19543 a_n2511_10356.n103 a_n2511_10356.n102 81.2397
R19544 a_n2511_10356.n37 a_n2511_10356.n36 81.2397
R19545 a_n2511_10356.n37 a_n2511_10356.n35 38.3829
R19546 a_n2511_10356.n135 a_n2511_10356.n134 37.8096
R19547 a_n2511_10356.n101 a_n2511_10356.n100 37.8096
R19548 a_n2511_10356.n69 a_n2511_10356.n68 37.8096
R19549 a_n2511_10356.n115 a_n2511_10356.n113 16.3865
R19550 a_n2511_10356.n81 a_n2511_10356.n79 16.3865
R19551 a_n2511_10356.n49 a_n2511_10356.n47 16.3865
R19552 a_n2511_10356.n16 a_n2511_10356.n14 16.3865
R19553 a_n2511_10356.n136 a_n2511_10356.n4 13.2313
R19554 a_n2511_10356.n116 a_n2511_10356.n112 12.8005
R19555 a_n2511_10356.n82 a_n2511_10356.n78 12.8005
R19556 a_n2511_10356.n50 a_n2511_10356.n46 12.8005
R19557 a_n2511_10356.n17 a_n2511_10356.n13 12.8005
R19558 a_n2511_10356.n120 a_n2511_10356.n119 12.0247
R19559 a_n2511_10356.n86 a_n2511_10356.n85 12.0247
R19560 a_n2511_10356.n54 a_n2511_10356.n53 12.0247
R19561 a_n2511_10356.n21 a_n2511_10356.n20 12.0247
R19562 a_n2511_10356.n123 a_n2511_10356.n110 11.249
R19563 a_n2511_10356.n89 a_n2511_10356.n76 11.249
R19564 a_n2511_10356.n57 a_n2511_10356.n44 11.249
R19565 a_n2511_10356.n24 a_n2511_10356.n11 11.249
R19566 a_n2511_10356.n124 a_n2511_10356.n108 10.4732
R19567 a_n2511_10356.n90 a_n2511_10356.n74 10.4732
R19568 a_n2511_10356.n58 a_n2511_10356.n42 10.4732
R19569 a_n2511_10356.n25 a_n2511_10356.n9 10.4732
R19570 a_n2511_10356.n138 a_n2511_10356.n136 10.4398
R19571 a_n2511_10356.n128 a_n2511_10356.n127 9.69747
R19572 a_n2511_10356.n94 a_n2511_10356.n93 9.69747
R19573 a_n2511_10356.n62 a_n2511_10356.n61 9.69747
R19574 a_n2511_10356.n29 a_n2511_10356.n28 9.69747
R19575 a_n2511_10356.n134 a_n2511_10356.n133 9.45567
R19576 a_n2511_10356.n100 a_n2511_10356.n99 9.45567
R19577 a_n2511_10356.n68 a_n2511_10356.n67 9.45567
R19578 a_n2511_10356.n35 a_n2511_10356.n34 9.45567
R19579 a_n2511_10356.n133 a_n2511_10356.n132 9.3005
R19580 a_n2511_10356.n106 a_n2511_10356.n105 9.3005
R19581 a_n2511_10356.n127 a_n2511_10356.n126 9.3005
R19582 a_n2511_10356.n125 a_n2511_10356.n124 9.3005
R19583 a_n2511_10356.n110 a_n2511_10356.n109 9.3005
R19584 a_n2511_10356.n119 a_n2511_10356.n118 9.3005
R19585 a_n2511_10356.n117 a_n2511_10356.n116 9.3005
R19586 a_n2511_10356.n99 a_n2511_10356.n98 9.3005
R19587 a_n2511_10356.n72 a_n2511_10356.n71 9.3005
R19588 a_n2511_10356.n93 a_n2511_10356.n92 9.3005
R19589 a_n2511_10356.n91 a_n2511_10356.n90 9.3005
R19590 a_n2511_10356.n76 a_n2511_10356.n75 9.3005
R19591 a_n2511_10356.n85 a_n2511_10356.n84 9.3005
R19592 a_n2511_10356.n83 a_n2511_10356.n82 9.3005
R19593 a_n2511_10356.n67 a_n2511_10356.n66 9.3005
R19594 a_n2511_10356.n40 a_n2511_10356.n39 9.3005
R19595 a_n2511_10356.n61 a_n2511_10356.n60 9.3005
R19596 a_n2511_10356.n59 a_n2511_10356.n58 9.3005
R19597 a_n2511_10356.n44 a_n2511_10356.n43 9.3005
R19598 a_n2511_10356.n53 a_n2511_10356.n52 9.3005
R19599 a_n2511_10356.n51 a_n2511_10356.n50 9.3005
R19600 a_n2511_10356.n34 a_n2511_10356.n33 9.3005
R19601 a_n2511_10356.n7 a_n2511_10356.n6 9.3005
R19602 a_n2511_10356.n28 a_n2511_10356.n27 9.3005
R19603 a_n2511_10356.n26 a_n2511_10356.n25 9.3005
R19604 a_n2511_10356.n11 a_n2511_10356.n10 9.3005
R19605 a_n2511_10356.n20 a_n2511_10356.n19 9.3005
R19606 a_n2511_10356.n18 a_n2511_10356.n17 9.3005
R19607 a_n2511_10356.n131 a_n2511_10356.n106 8.92171
R19608 a_n2511_10356.n97 a_n2511_10356.n72 8.92171
R19609 a_n2511_10356.n65 a_n2511_10356.n40 8.92171
R19610 a_n2511_10356.n32 a_n2511_10356.n7 8.92171
R19611 a_n2511_10356.n132 a_n2511_10356.n104 8.14595
R19612 a_n2511_10356.n98 a_n2511_10356.n70 8.14595
R19613 a_n2511_10356.n66 a_n2511_10356.n38 8.14595
R19614 a_n2511_10356.n33 a_n2511_10356.n5 8.14595
R19615 a_n2511_10356.n136 a_n2511_10356.n135 5.91753
R19616 a_n2511_10356.n134 a_n2511_10356.n104 5.81868
R19617 a_n2511_10356.n100 a_n2511_10356.n70 5.81868
R19618 a_n2511_10356.n68 a_n2511_10356.n38 5.81868
R19619 a_n2511_10356.n35 a_n2511_10356.n5 5.81868
R19620 a_n2511_10356.n137 a_n2511_10356.t12 5.418
R19621 a_n2511_10356.n137 a_n2511_10356.t14 5.418
R19622 a_n2511_10356.n139 a_n2511_10356.t10 5.418
R19623 a_n2511_10356.n139 a_n2511_10356.t8 5.418
R19624 a_n2511_10356.n102 a_n2511_10356.t2 5.418
R19625 a_n2511_10356.n102 a_n2511_10356.t4 5.418
R19626 a_n2511_10356.n36 a_n2511_10356.t5 5.418
R19627 a_n2511_10356.n36 a_n2511_10356.t7 5.418
R19628 a_n2511_10356.n3 a_n2511_10356.t15 5.418
R19629 a_n2511_10356.n3 a_n2511_10356.t19 5.418
R19630 a_n2511_10356.n1 a_n2511_10356.t11 5.418
R19631 a_n2511_10356.n1 a_n2511_10356.t13 5.418
R19632 a_n2511_10356.n0 a_n2511_10356.t17 5.418
R19633 a_n2511_10356.n0 a_n2511_10356.t16 5.418
R19634 a_n2511_10356.t18 a_n2511_10356.n141 5.418
R19635 a_n2511_10356.n141 a_n2511_10356.t9 5.418
R19636 a_n2511_10356.n132 a_n2511_10356.n131 5.04292
R19637 a_n2511_10356.n98 a_n2511_10356.n97 5.04292
R19638 a_n2511_10356.n66 a_n2511_10356.n65 5.04292
R19639 a_n2511_10356.n33 a_n2511_10356.n32 5.04292
R19640 a_n2511_10356.n128 a_n2511_10356.n106 4.26717
R19641 a_n2511_10356.n94 a_n2511_10356.n72 4.26717
R19642 a_n2511_10356.n62 a_n2511_10356.n40 4.26717
R19643 a_n2511_10356.n29 a_n2511_10356.n7 4.26717
R19644 a_n2511_10356.n117 a_n2511_10356.n113 3.71286
R19645 a_n2511_10356.n83 a_n2511_10356.n79 3.71286
R19646 a_n2511_10356.n51 a_n2511_10356.n47 3.71286
R19647 a_n2511_10356.n18 a_n2511_10356.n14 3.71286
R19648 a_n2511_10356.n127 a_n2511_10356.n108 3.49141
R19649 a_n2511_10356.n93 a_n2511_10356.n74 3.49141
R19650 a_n2511_10356.n61 a_n2511_10356.n42 3.49141
R19651 a_n2511_10356.n28 a_n2511_10356.n9 3.49141
R19652 a_n2511_10356.n124 a_n2511_10356.n123 2.71565
R19653 a_n2511_10356.n90 a_n2511_10356.n89 2.71565
R19654 a_n2511_10356.n58 a_n2511_10356.n57 2.71565
R19655 a_n2511_10356.n25 a_n2511_10356.n24 2.71565
R19656 a_n2511_10356.n120 a_n2511_10356.n110 1.93989
R19657 a_n2511_10356.n86 a_n2511_10356.n76 1.93989
R19658 a_n2511_10356.n54 a_n2511_10356.n44 1.93989
R19659 a_n2511_10356.n21 a_n2511_10356.n11 1.93989
R19660 a_n2511_10356.n119 a_n2511_10356.n112 1.16414
R19661 a_n2511_10356.n85 a_n2511_10356.n78 1.16414
R19662 a_n2511_10356.n53 a_n2511_10356.n46 1.16414
R19663 a_n2511_10356.n20 a_n2511_10356.n13 1.16414
R19664 a_n2511_10356.n69 a_n2511_10356.n37 0.573776
R19665 a_n2511_10356.n103 a_n2511_10356.n101 0.573776
R19666 a_n2511_10356.n135 a_n2511_10356.n103 0.573776
R19667 a_n2511_10356.n140 a_n2511_10356.n138 0.573776
R19668 a_n2511_10356.n116 a_n2511_10356.n115 0.388379
R19669 a_n2511_10356.n82 a_n2511_10356.n81 0.388379
R19670 a_n2511_10356.n50 a_n2511_10356.n49 0.388379
R19671 a_n2511_10356.n17 a_n2511_10356.n16 0.388379
R19672 a_n2511_10356.n4 a_n2511_10356.n2 0.234655
R19673 a_n2511_10356.n133 a_n2511_10356.n105 0.155672
R19674 a_n2511_10356.n126 a_n2511_10356.n105 0.155672
R19675 a_n2511_10356.n126 a_n2511_10356.n125 0.155672
R19676 a_n2511_10356.n125 a_n2511_10356.n109 0.155672
R19677 a_n2511_10356.n118 a_n2511_10356.n109 0.155672
R19678 a_n2511_10356.n118 a_n2511_10356.n117 0.155672
R19679 a_n2511_10356.n99 a_n2511_10356.n71 0.155672
R19680 a_n2511_10356.n92 a_n2511_10356.n71 0.155672
R19681 a_n2511_10356.n92 a_n2511_10356.n91 0.155672
R19682 a_n2511_10356.n91 a_n2511_10356.n75 0.155672
R19683 a_n2511_10356.n84 a_n2511_10356.n75 0.155672
R19684 a_n2511_10356.n84 a_n2511_10356.n83 0.155672
R19685 a_n2511_10356.n67 a_n2511_10356.n39 0.155672
R19686 a_n2511_10356.n60 a_n2511_10356.n39 0.155672
R19687 a_n2511_10356.n60 a_n2511_10356.n59 0.155672
R19688 a_n2511_10356.n59 a_n2511_10356.n43 0.155672
R19689 a_n2511_10356.n52 a_n2511_10356.n43 0.155672
R19690 a_n2511_10356.n52 a_n2511_10356.n51 0.155672
R19691 a_n2511_10356.n34 a_n2511_10356.n6 0.155672
R19692 a_n2511_10356.n27 a_n2511_10356.n6 0.155672
R19693 a_n2511_10356.n27 a_n2511_10356.n26 0.155672
R19694 a_n2511_10356.n26 a_n2511_10356.n10 0.155672
R19695 a_n2511_10356.n19 a_n2511_10356.n10 0.155672
R19696 a_n2511_10356.n19 a_n2511_10356.n18 0.155672
R19697 a_n2511_10356.n101 a_n2511_10356.n69 0.155672
R19698 VN.n28 VN.t0 243.97
R19699 VN.n28 VN.n27 223.454
R19700 VN.n30 VN.n29 223.454
R19701 VN.n15 VN.t7 199.144
R19702 VN.n2 VN.t5 199.144
R19703 VN.n24 VN.t10 183.883
R19704 VN.n11 VN.t9 183.883
R19705 VN.n23 VN.n13 161.3
R19706 VN.n21 VN.n20 161.3
R19707 VN.n19 VN.n14 161.3
R19708 VN.n18 VN.n17 161.3
R19709 VN.n5 VN.n4 161.3
R19710 VN.n6 VN.n1 161.3
R19711 VN.n8 VN.n7 161.3
R19712 VN.n10 VN.n0 161.3
R19713 VN.n16 VN.t6 144.601
R19714 VN.n22 VN.t11 144.601
R19715 VN.n9 VN.t8 144.601
R19716 VN.n3 VN.t12 144.601
R19717 VN.n25 VN.n24 80.6037
R19718 VN.n12 VN.n11 80.6037
R19719 VN.n24 VN.n23 56.3158
R19720 VN.n11 VN.n10 56.3158
R19721 VN.n16 VN.n15 46.9082
R19722 VN.n3 VN.n2 46.9082
R19723 VN.n18 VN.n15 43.8991
R19724 VN.n5 VN.n2 43.8991
R19725 VN.n17 VN.n14 40.577
R19726 VN.n21 VN.n14 40.577
R19727 VN.n8 VN.n1 40.577
R19728 VN.n4 VN.n1 40.577
R19729 VN.n26 VN.n25 27.893
R19730 VN.n27 VN.t1 19.8005
R19731 VN.n27 VN.t4 19.8005
R19732 VN.n29 VN.t2 19.8005
R19733 VN.n29 VN.t3 19.8005
R19734 VN.n23 VN.n22 16.477
R19735 VN.n10 VN.n9 16.477
R19736 VN VN.n31 14.1384
R19737 VN.n26 VN.n12 11.6998
R19738 VN.n17 VN.n16 8.11581
R19739 VN.n22 VN.n21 8.11581
R19740 VN.n9 VN.n8 8.11581
R19741 VN.n4 VN.n3 8.11581
R19742 VN.n31 VN.n30 5.40567
R19743 VN.n31 VN.n26 1.188
R19744 VN.n30 VN.n28 0.716017
R19745 VN.n25 VN.n13 0.285035
R19746 VN.n12 VN.n0 0.285035
R19747 VN.n19 VN.n18 0.189894
R19748 VN.n20 VN.n19 0.189894
R19749 VN.n20 VN.n13 0.189894
R19750 VN.n7 VN.n0 0.189894
R19751 VN.n7 VN.n6 0.189894
R19752 VN.n6 VN.n5 0.189894
R19753 a_n1455_n3628.n308 a_n1455_n3628.n288 289.615
R19754 a_n1455_n3628.n335 a_n1455_n3628.n315 289.615
R19755 a_n1455_n3628.n177 a_n1455_n3628.n157 289.615
R19756 a_n1455_n3628.n281 a_n1455_n3628.n261 289.615
R19757 a_n1455_n3628.n255 a_n1455_n3628.n235 289.615
R19758 a_n1455_n3628.n229 a_n1455_n3628.n209 289.615
R19759 a_n1455_n3628.n203 a_n1455_n3628.n183 289.615
R19760 a_n1455_n3628.n69 a_n1455_n3628.n49 289.615
R19761 a_n1455_n3628.n97 a_n1455_n3628.n77 289.615
R19762 a_n1455_n3628.n123 a_n1455_n3628.n103 289.615
R19763 a_n1455_n3628.n151 a_n1455_n3628.n131 289.615
R19764 a_n1455_n3628.n344 a_n1455_n3628.n46 289.615
R19765 a_n1455_n3628.n208 a_n1455_n3628.n207 196.838
R19766 a_n1455_n3628.n286 a_n1455_n3628.n285 196.298
R19767 a_n1455_n3628.n260 a_n1455_n3628.n259 196.298
R19768 a_n1455_n3628.n234 a_n1455_n3628.n233 196.298
R19769 a_n1455_n3628.n297 a_n1455_n3628.n296 185
R19770 a_n1455_n3628.n294 a_n1455_n3628.n293 185
R19771 a_n1455_n3628.n301 a_n1455_n3628.n300 185
R19772 a_n1455_n3628.n303 a_n1455_n3628.n302 185
R19773 a_n1455_n3628.n291 a_n1455_n3628.n290 185
R19774 a_n1455_n3628.n307 a_n1455_n3628.n306 185
R19775 a_n1455_n3628.n309 a_n1455_n3628.n308 185
R19776 a_n1455_n3628.n324 a_n1455_n3628.n323 185
R19777 a_n1455_n3628.n321 a_n1455_n3628.n320 185
R19778 a_n1455_n3628.n328 a_n1455_n3628.n327 185
R19779 a_n1455_n3628.n330 a_n1455_n3628.n329 185
R19780 a_n1455_n3628.n318 a_n1455_n3628.n317 185
R19781 a_n1455_n3628.n334 a_n1455_n3628.n333 185
R19782 a_n1455_n3628.n336 a_n1455_n3628.n335 185
R19783 a_n1455_n3628.n166 a_n1455_n3628.n165 185
R19784 a_n1455_n3628.n163 a_n1455_n3628.n162 185
R19785 a_n1455_n3628.n170 a_n1455_n3628.n169 185
R19786 a_n1455_n3628.n172 a_n1455_n3628.n171 185
R19787 a_n1455_n3628.n160 a_n1455_n3628.n159 185
R19788 a_n1455_n3628.n176 a_n1455_n3628.n175 185
R19789 a_n1455_n3628.n178 a_n1455_n3628.n177 185
R19790 a_n1455_n3628.n282 a_n1455_n3628.n281 185
R19791 a_n1455_n3628.n280 a_n1455_n3628.n279 185
R19792 a_n1455_n3628.n264 a_n1455_n3628.n263 185
R19793 a_n1455_n3628.n276 a_n1455_n3628.n275 185
R19794 a_n1455_n3628.n274 a_n1455_n3628.n273 185
R19795 a_n1455_n3628.n267 a_n1455_n3628.n266 185
R19796 a_n1455_n3628.n270 a_n1455_n3628.n269 185
R19797 a_n1455_n3628.n256 a_n1455_n3628.n255 185
R19798 a_n1455_n3628.n254 a_n1455_n3628.n253 185
R19799 a_n1455_n3628.n238 a_n1455_n3628.n237 185
R19800 a_n1455_n3628.n250 a_n1455_n3628.n249 185
R19801 a_n1455_n3628.n248 a_n1455_n3628.n247 185
R19802 a_n1455_n3628.n241 a_n1455_n3628.n240 185
R19803 a_n1455_n3628.n244 a_n1455_n3628.n243 185
R19804 a_n1455_n3628.n230 a_n1455_n3628.n229 185
R19805 a_n1455_n3628.n228 a_n1455_n3628.n227 185
R19806 a_n1455_n3628.n212 a_n1455_n3628.n211 185
R19807 a_n1455_n3628.n224 a_n1455_n3628.n223 185
R19808 a_n1455_n3628.n222 a_n1455_n3628.n221 185
R19809 a_n1455_n3628.n215 a_n1455_n3628.n214 185
R19810 a_n1455_n3628.n218 a_n1455_n3628.n217 185
R19811 a_n1455_n3628.n204 a_n1455_n3628.n203 185
R19812 a_n1455_n3628.n202 a_n1455_n3628.n201 185
R19813 a_n1455_n3628.n186 a_n1455_n3628.n185 185
R19814 a_n1455_n3628.n198 a_n1455_n3628.n197 185
R19815 a_n1455_n3628.n196 a_n1455_n3628.n195 185
R19816 a_n1455_n3628.n189 a_n1455_n3628.n188 185
R19817 a_n1455_n3628.n192 a_n1455_n3628.n191 185
R19818 a_n1455_n3628.n70 a_n1455_n3628.n69 185
R19819 a_n1455_n3628.n68 a_n1455_n3628.n67 185
R19820 a_n1455_n3628.n52 a_n1455_n3628.n51 185
R19821 a_n1455_n3628.n64 a_n1455_n3628.n63 185
R19822 a_n1455_n3628.n62 a_n1455_n3628.n61 185
R19823 a_n1455_n3628.n55 a_n1455_n3628.n54 185
R19824 a_n1455_n3628.n58 a_n1455_n3628.n57 185
R19825 a_n1455_n3628.n98 a_n1455_n3628.n97 185
R19826 a_n1455_n3628.n96 a_n1455_n3628.n95 185
R19827 a_n1455_n3628.n80 a_n1455_n3628.n79 185
R19828 a_n1455_n3628.n92 a_n1455_n3628.n91 185
R19829 a_n1455_n3628.n90 a_n1455_n3628.n89 185
R19830 a_n1455_n3628.n83 a_n1455_n3628.n82 185
R19831 a_n1455_n3628.n86 a_n1455_n3628.n85 185
R19832 a_n1455_n3628.n124 a_n1455_n3628.n123 185
R19833 a_n1455_n3628.n122 a_n1455_n3628.n121 185
R19834 a_n1455_n3628.n106 a_n1455_n3628.n105 185
R19835 a_n1455_n3628.n118 a_n1455_n3628.n117 185
R19836 a_n1455_n3628.n116 a_n1455_n3628.n115 185
R19837 a_n1455_n3628.n109 a_n1455_n3628.n108 185
R19838 a_n1455_n3628.n112 a_n1455_n3628.n111 185
R19839 a_n1455_n3628.n152 a_n1455_n3628.n151 185
R19840 a_n1455_n3628.n150 a_n1455_n3628.n149 185
R19841 a_n1455_n3628.n134 a_n1455_n3628.n133 185
R19842 a_n1455_n3628.n146 a_n1455_n3628.n145 185
R19843 a_n1455_n3628.n144 a_n1455_n3628.n143 185
R19844 a_n1455_n3628.n137 a_n1455_n3628.n136 185
R19845 a_n1455_n3628.n140 a_n1455_n3628.n139 185
R19846 a_n1455_n3628.n357 a_n1455_n3628.n356 185
R19847 a_n1455_n3628.n41 a_n1455_n3628.n40 185
R19848 a_n1455_n3628.n352 a_n1455_n3628.n351 185
R19849 a_n1455_n3628.n350 a_n1455_n3628.n349 185
R19850 a_n1455_n3628.n44 a_n1455_n3628.n43 185
R19851 a_n1455_n3628.n346 a_n1455_n3628.n345 185
R19852 a_n1455_n3628.n344 a_n1455_n3628.n343 185
R19853 a_n1455_n3628.t17 a_n1455_n3628.n295 147.661
R19854 a_n1455_n3628.t9 a_n1455_n3628.n322 147.661
R19855 a_n1455_n3628.t3 a_n1455_n3628.n164 147.661
R19856 a_n1455_n3628.t13 a_n1455_n3628.n268 147.661
R19857 a_n1455_n3628.t14 a_n1455_n3628.n242 147.661
R19858 a_n1455_n3628.t12 a_n1455_n3628.n216 147.661
R19859 a_n1455_n3628.t11 a_n1455_n3628.n190 147.661
R19860 a_n1455_n3628.t2 a_n1455_n3628.n56 147.661
R19861 a_n1455_n3628.t5 a_n1455_n3628.n84 147.661
R19862 a_n1455_n3628.t18 a_n1455_n3628.n110 147.661
R19863 a_n1455_n3628.t15 a_n1455_n3628.n138 147.661
R19864 a_n1455_n3628.t7 a_n1455_n3628.n39 147.661
R19865 a_n1455_n3628.n296 a_n1455_n3628.n293 104.615
R19866 a_n1455_n3628.n301 a_n1455_n3628.n293 104.615
R19867 a_n1455_n3628.n302 a_n1455_n3628.n301 104.615
R19868 a_n1455_n3628.n302 a_n1455_n3628.n290 104.615
R19869 a_n1455_n3628.n307 a_n1455_n3628.n290 104.615
R19870 a_n1455_n3628.n308 a_n1455_n3628.n307 104.615
R19871 a_n1455_n3628.n323 a_n1455_n3628.n320 104.615
R19872 a_n1455_n3628.n328 a_n1455_n3628.n320 104.615
R19873 a_n1455_n3628.n329 a_n1455_n3628.n328 104.615
R19874 a_n1455_n3628.n329 a_n1455_n3628.n317 104.615
R19875 a_n1455_n3628.n334 a_n1455_n3628.n317 104.615
R19876 a_n1455_n3628.n335 a_n1455_n3628.n334 104.615
R19877 a_n1455_n3628.n165 a_n1455_n3628.n162 104.615
R19878 a_n1455_n3628.n170 a_n1455_n3628.n162 104.615
R19879 a_n1455_n3628.n171 a_n1455_n3628.n170 104.615
R19880 a_n1455_n3628.n171 a_n1455_n3628.n159 104.615
R19881 a_n1455_n3628.n176 a_n1455_n3628.n159 104.615
R19882 a_n1455_n3628.n177 a_n1455_n3628.n176 104.615
R19883 a_n1455_n3628.n281 a_n1455_n3628.n280 104.615
R19884 a_n1455_n3628.n280 a_n1455_n3628.n263 104.615
R19885 a_n1455_n3628.n275 a_n1455_n3628.n263 104.615
R19886 a_n1455_n3628.n275 a_n1455_n3628.n274 104.615
R19887 a_n1455_n3628.n274 a_n1455_n3628.n266 104.615
R19888 a_n1455_n3628.n269 a_n1455_n3628.n266 104.615
R19889 a_n1455_n3628.n255 a_n1455_n3628.n254 104.615
R19890 a_n1455_n3628.n254 a_n1455_n3628.n237 104.615
R19891 a_n1455_n3628.n249 a_n1455_n3628.n237 104.615
R19892 a_n1455_n3628.n249 a_n1455_n3628.n248 104.615
R19893 a_n1455_n3628.n248 a_n1455_n3628.n240 104.615
R19894 a_n1455_n3628.n243 a_n1455_n3628.n240 104.615
R19895 a_n1455_n3628.n229 a_n1455_n3628.n228 104.615
R19896 a_n1455_n3628.n228 a_n1455_n3628.n211 104.615
R19897 a_n1455_n3628.n223 a_n1455_n3628.n211 104.615
R19898 a_n1455_n3628.n223 a_n1455_n3628.n222 104.615
R19899 a_n1455_n3628.n222 a_n1455_n3628.n214 104.615
R19900 a_n1455_n3628.n217 a_n1455_n3628.n214 104.615
R19901 a_n1455_n3628.n203 a_n1455_n3628.n202 104.615
R19902 a_n1455_n3628.n202 a_n1455_n3628.n185 104.615
R19903 a_n1455_n3628.n197 a_n1455_n3628.n185 104.615
R19904 a_n1455_n3628.n197 a_n1455_n3628.n196 104.615
R19905 a_n1455_n3628.n196 a_n1455_n3628.n188 104.615
R19906 a_n1455_n3628.n191 a_n1455_n3628.n188 104.615
R19907 a_n1455_n3628.n69 a_n1455_n3628.n68 104.615
R19908 a_n1455_n3628.n68 a_n1455_n3628.n51 104.615
R19909 a_n1455_n3628.n63 a_n1455_n3628.n51 104.615
R19910 a_n1455_n3628.n63 a_n1455_n3628.n62 104.615
R19911 a_n1455_n3628.n62 a_n1455_n3628.n54 104.615
R19912 a_n1455_n3628.n57 a_n1455_n3628.n54 104.615
R19913 a_n1455_n3628.n97 a_n1455_n3628.n96 104.615
R19914 a_n1455_n3628.n96 a_n1455_n3628.n79 104.615
R19915 a_n1455_n3628.n91 a_n1455_n3628.n79 104.615
R19916 a_n1455_n3628.n91 a_n1455_n3628.n90 104.615
R19917 a_n1455_n3628.n90 a_n1455_n3628.n82 104.615
R19918 a_n1455_n3628.n85 a_n1455_n3628.n82 104.615
R19919 a_n1455_n3628.n123 a_n1455_n3628.n122 104.615
R19920 a_n1455_n3628.n122 a_n1455_n3628.n105 104.615
R19921 a_n1455_n3628.n117 a_n1455_n3628.n105 104.615
R19922 a_n1455_n3628.n117 a_n1455_n3628.n116 104.615
R19923 a_n1455_n3628.n116 a_n1455_n3628.n108 104.615
R19924 a_n1455_n3628.n111 a_n1455_n3628.n108 104.615
R19925 a_n1455_n3628.n151 a_n1455_n3628.n150 104.615
R19926 a_n1455_n3628.n150 a_n1455_n3628.n133 104.615
R19927 a_n1455_n3628.n145 a_n1455_n3628.n133 104.615
R19928 a_n1455_n3628.n145 a_n1455_n3628.n144 104.615
R19929 a_n1455_n3628.n144 a_n1455_n3628.n136 104.615
R19930 a_n1455_n3628.n139 a_n1455_n3628.n136 104.615
R19931 a_n1455_n3628.n357 a_n1455_n3628.n40 104.615
R19932 a_n1455_n3628.n351 a_n1455_n3628.n40 104.615
R19933 a_n1455_n3628.n351 a_n1455_n3628.n350 104.615
R19934 a_n1455_n3628.n350 a_n1455_n3628.n43 104.615
R19935 a_n1455_n3628.n345 a_n1455_n3628.n43 104.615
R19936 a_n1455_n3628.n345 a_n1455_n3628.n344 104.615
R19937 a_n1455_n3628.n76 a_n1455_n3628.n75 56.1363
R19938 a_n1455_n3628.n130 a_n1455_n3628.n129 56.1363
R19939 a_n1455_n3628.n314 a_n1455_n3628.n313 56.1361
R19940 a_n1455_n3628.n48 a_n1455_n3628.n47 56.1361
R19941 a_n1455_n3628.n296 a_n1455_n3628.t17 52.3082
R19942 a_n1455_n3628.n323 a_n1455_n3628.t9 52.3082
R19943 a_n1455_n3628.n165 a_n1455_n3628.t3 52.3082
R19944 a_n1455_n3628.n269 a_n1455_n3628.t13 52.3082
R19945 a_n1455_n3628.n243 a_n1455_n3628.t14 52.3082
R19946 a_n1455_n3628.n217 a_n1455_n3628.t12 52.3082
R19947 a_n1455_n3628.n191 a_n1455_n3628.t11 52.3082
R19948 a_n1455_n3628.n57 a_n1455_n3628.t2 52.3082
R19949 a_n1455_n3628.n85 a_n1455_n3628.t5 52.3082
R19950 a_n1455_n3628.n111 a_n1455_n3628.t18 52.3082
R19951 a_n1455_n3628.n139 a_n1455_n3628.t15 52.3082
R19952 a_n1455_n3628.t7 a_n1455_n3628.n357 52.3082
R19953 a_n1455_n3628.n312 a_n1455_n3628.n311 37.8096
R19954 a_n1455_n3628.n339 a_n1455_n3628.n338 37.8096
R19955 a_n1455_n3628.n181 a_n1455_n3628.n180 37.8096
R19956 a_n1455_n3628.n74 a_n1455_n3628.n73 37.8096
R19957 a_n1455_n3628.n102 a_n1455_n3628.n101 37.8096
R19958 a_n1455_n3628.n128 a_n1455_n3628.n127 37.8096
R19959 a_n1455_n3628.n156 a_n1455_n3628.n155 37.8096
R19960 a_n1455_n3628.n341 a_n1455_n3628.n340 37.8096
R19961 a_n1455_n3628.n297 a_n1455_n3628.n295 15.6674
R19962 a_n1455_n3628.n324 a_n1455_n3628.n322 15.6674
R19963 a_n1455_n3628.n166 a_n1455_n3628.n164 15.6674
R19964 a_n1455_n3628.n270 a_n1455_n3628.n268 15.6674
R19965 a_n1455_n3628.n244 a_n1455_n3628.n242 15.6674
R19966 a_n1455_n3628.n218 a_n1455_n3628.n216 15.6674
R19967 a_n1455_n3628.n192 a_n1455_n3628.n190 15.6674
R19968 a_n1455_n3628.n58 a_n1455_n3628.n56 15.6674
R19969 a_n1455_n3628.n86 a_n1455_n3628.n84 15.6674
R19970 a_n1455_n3628.n112 a_n1455_n3628.n110 15.6674
R19971 a_n1455_n3628.n140 a_n1455_n3628.n138 15.6674
R19972 a_n1455_n3628.n356 a_n1455_n3628.n39 15.6674
R19973 a_n1455_n3628.n298 a_n1455_n3628.n294 12.8005
R19974 a_n1455_n3628.n325 a_n1455_n3628.n321 12.8005
R19975 a_n1455_n3628.n167 a_n1455_n3628.n163 12.8005
R19976 a_n1455_n3628.n271 a_n1455_n3628.n267 12.8005
R19977 a_n1455_n3628.n245 a_n1455_n3628.n241 12.8005
R19978 a_n1455_n3628.n219 a_n1455_n3628.n215 12.8005
R19979 a_n1455_n3628.n193 a_n1455_n3628.n189 12.8005
R19980 a_n1455_n3628.n59 a_n1455_n3628.n55 12.8005
R19981 a_n1455_n3628.n87 a_n1455_n3628.n83 12.8005
R19982 a_n1455_n3628.n113 a_n1455_n3628.n109 12.8005
R19983 a_n1455_n3628.n141 a_n1455_n3628.n137 12.8005
R19984 a_n1455_n3628.n355 a_n1455_n3628.n41 12.8005
R19985 a_n1455_n3628.n300 a_n1455_n3628.n299 12.0247
R19986 a_n1455_n3628.n327 a_n1455_n3628.n326 12.0247
R19987 a_n1455_n3628.n169 a_n1455_n3628.n168 12.0247
R19988 a_n1455_n3628.n273 a_n1455_n3628.n272 12.0247
R19989 a_n1455_n3628.n247 a_n1455_n3628.n246 12.0247
R19990 a_n1455_n3628.n221 a_n1455_n3628.n220 12.0247
R19991 a_n1455_n3628.n195 a_n1455_n3628.n194 12.0247
R19992 a_n1455_n3628.n61 a_n1455_n3628.n60 12.0247
R19993 a_n1455_n3628.n89 a_n1455_n3628.n88 12.0247
R19994 a_n1455_n3628.n115 a_n1455_n3628.n114 12.0247
R19995 a_n1455_n3628.n143 a_n1455_n3628.n142 12.0247
R19996 a_n1455_n3628.n353 a_n1455_n3628.n352 12.0247
R19997 a_n1455_n3628.n182 a_n1455_n3628.n156 11.5057
R19998 a_n1455_n3628.n287 a_n1455_n3628.n74 11.5057
R19999 a_n1455_n3628.n303 a_n1455_n3628.n292 11.249
R20000 a_n1455_n3628.n330 a_n1455_n3628.n319 11.249
R20001 a_n1455_n3628.n172 a_n1455_n3628.n161 11.249
R20002 a_n1455_n3628.n276 a_n1455_n3628.n265 11.249
R20003 a_n1455_n3628.n250 a_n1455_n3628.n239 11.249
R20004 a_n1455_n3628.n224 a_n1455_n3628.n213 11.249
R20005 a_n1455_n3628.n198 a_n1455_n3628.n187 11.249
R20006 a_n1455_n3628.n64 a_n1455_n3628.n53 11.249
R20007 a_n1455_n3628.n92 a_n1455_n3628.n81 11.249
R20008 a_n1455_n3628.n118 a_n1455_n3628.n107 11.249
R20009 a_n1455_n3628.n146 a_n1455_n3628.n135 11.249
R20010 a_n1455_n3628.n349 a_n1455_n3628.n42 11.249
R20011 a_n1455_n3628.n304 a_n1455_n3628.n291 10.4732
R20012 a_n1455_n3628.n331 a_n1455_n3628.n318 10.4732
R20013 a_n1455_n3628.n173 a_n1455_n3628.n160 10.4732
R20014 a_n1455_n3628.n277 a_n1455_n3628.n264 10.4732
R20015 a_n1455_n3628.n251 a_n1455_n3628.n238 10.4732
R20016 a_n1455_n3628.n225 a_n1455_n3628.n212 10.4732
R20017 a_n1455_n3628.n199 a_n1455_n3628.n186 10.4732
R20018 a_n1455_n3628.n65 a_n1455_n3628.n52 10.4732
R20019 a_n1455_n3628.n93 a_n1455_n3628.n80 10.4732
R20020 a_n1455_n3628.n119 a_n1455_n3628.n106 10.4732
R20021 a_n1455_n3628.n147 a_n1455_n3628.n134 10.4732
R20022 a_n1455_n3628.n348 a_n1455_n3628.n44 10.4732
R20023 a_n1455_n3628.n306 a_n1455_n3628.n305 9.69747
R20024 a_n1455_n3628.n333 a_n1455_n3628.n332 9.69747
R20025 a_n1455_n3628.n175 a_n1455_n3628.n174 9.69747
R20026 a_n1455_n3628.n279 a_n1455_n3628.n278 9.69747
R20027 a_n1455_n3628.n253 a_n1455_n3628.n252 9.69747
R20028 a_n1455_n3628.n227 a_n1455_n3628.n226 9.69747
R20029 a_n1455_n3628.n201 a_n1455_n3628.n200 9.69747
R20030 a_n1455_n3628.n67 a_n1455_n3628.n66 9.69747
R20031 a_n1455_n3628.n95 a_n1455_n3628.n94 9.69747
R20032 a_n1455_n3628.n121 a_n1455_n3628.n120 9.69747
R20033 a_n1455_n3628.n149 a_n1455_n3628.n148 9.69747
R20034 a_n1455_n3628.n347 a_n1455_n3628.n346 9.69747
R20035 a_n1455_n3628.n1 a_n1455_n3628.n341 9.45567
R20036 a_n1455_n3628.n311 a_n1455_n3628.n5 9.45567
R20037 a_n1455_n3628.n338 a_n1455_n3628.n9 9.45567
R20038 a_n1455_n3628.n180 a_n1455_n3628.n13 9.45567
R20039 a_n1455_n3628.n285 a_n1455_n3628.n284 9.45567
R20040 a_n1455_n3628.n259 a_n1455_n3628.n258 9.45567
R20041 a_n1455_n3628.n233 a_n1455_n3628.n232 9.45567
R20042 a_n1455_n3628.n207 a_n1455_n3628.n206 9.45567
R20043 a_n1455_n3628.n73 a_n1455_n3628.n72 9.45567
R20044 a_n1455_n3628.n101 a_n1455_n3628.n100 9.45567
R20045 a_n1455_n3628.n127 a_n1455_n3628.n126 9.45567
R20046 a_n1455_n3628.n155 a_n1455_n3628.n154 9.45567
R20047 a_n1455_n3628.n5 a_n1455_n3628.n310 9.3005
R20048 a_n1455_n3628.n289 a_n1455_n3628.n5 9.3005
R20049 a_n1455_n3628.n305 a_n1455_n3628.n6 9.3005
R20050 a_n1455_n3628.n6 a_n1455_n3628.n304 9.3005
R20051 a_n1455_n3628.n292 a_n1455_n3628.n4 9.3005
R20052 a_n1455_n3628.n299 a_n1455_n3628.n4 9.3005
R20053 a_n1455_n3628.n3 a_n1455_n3628.n298 9.3005
R20054 a_n1455_n3628.n9 a_n1455_n3628.n337 9.3005
R20055 a_n1455_n3628.n316 a_n1455_n3628.n9 9.3005
R20056 a_n1455_n3628.n332 a_n1455_n3628.n10 9.3005
R20057 a_n1455_n3628.n10 a_n1455_n3628.n331 9.3005
R20058 a_n1455_n3628.n319 a_n1455_n3628.n8 9.3005
R20059 a_n1455_n3628.n326 a_n1455_n3628.n8 9.3005
R20060 a_n1455_n3628.n7 a_n1455_n3628.n325 9.3005
R20061 a_n1455_n3628.n13 a_n1455_n3628.n179 9.3005
R20062 a_n1455_n3628.n158 a_n1455_n3628.n13 9.3005
R20063 a_n1455_n3628.n174 a_n1455_n3628.n14 9.3005
R20064 a_n1455_n3628.n14 a_n1455_n3628.n173 9.3005
R20065 a_n1455_n3628.n161 a_n1455_n3628.n12 9.3005
R20066 a_n1455_n3628.n168 a_n1455_n3628.n12 9.3005
R20067 a_n1455_n3628.n11 a_n1455_n3628.n167 9.3005
R20068 a_n1455_n3628.n284 a_n1455_n3628.n283 9.3005
R20069 a_n1455_n3628.n262 a_n1455_n3628.n16 9.3005
R20070 a_n1455_n3628.n278 a_n1455_n3628.n16 9.3005
R20071 a_n1455_n3628.n15 a_n1455_n3628.n277 9.3005
R20072 a_n1455_n3628.n265 a_n1455_n3628.n15 9.3005
R20073 a_n1455_n3628.n272 a_n1455_n3628.n17 9.3005
R20074 a_n1455_n3628.n17 a_n1455_n3628.n271 9.3005
R20075 a_n1455_n3628.n258 a_n1455_n3628.n257 9.3005
R20076 a_n1455_n3628.n236 a_n1455_n3628.n19 9.3005
R20077 a_n1455_n3628.n252 a_n1455_n3628.n19 9.3005
R20078 a_n1455_n3628.n18 a_n1455_n3628.n251 9.3005
R20079 a_n1455_n3628.n239 a_n1455_n3628.n18 9.3005
R20080 a_n1455_n3628.n246 a_n1455_n3628.n20 9.3005
R20081 a_n1455_n3628.n20 a_n1455_n3628.n245 9.3005
R20082 a_n1455_n3628.n232 a_n1455_n3628.n231 9.3005
R20083 a_n1455_n3628.n210 a_n1455_n3628.n22 9.3005
R20084 a_n1455_n3628.n226 a_n1455_n3628.n22 9.3005
R20085 a_n1455_n3628.n21 a_n1455_n3628.n225 9.3005
R20086 a_n1455_n3628.n213 a_n1455_n3628.n21 9.3005
R20087 a_n1455_n3628.n220 a_n1455_n3628.n23 9.3005
R20088 a_n1455_n3628.n23 a_n1455_n3628.n219 9.3005
R20089 a_n1455_n3628.n206 a_n1455_n3628.n205 9.3005
R20090 a_n1455_n3628.n184 a_n1455_n3628.n25 9.3005
R20091 a_n1455_n3628.n200 a_n1455_n3628.n25 9.3005
R20092 a_n1455_n3628.n24 a_n1455_n3628.n199 9.3005
R20093 a_n1455_n3628.n187 a_n1455_n3628.n24 9.3005
R20094 a_n1455_n3628.n194 a_n1455_n3628.n26 9.3005
R20095 a_n1455_n3628.n26 a_n1455_n3628.n193 9.3005
R20096 a_n1455_n3628.n72 a_n1455_n3628.n71 9.3005
R20097 a_n1455_n3628.n50 a_n1455_n3628.n28 9.3005
R20098 a_n1455_n3628.n66 a_n1455_n3628.n28 9.3005
R20099 a_n1455_n3628.n27 a_n1455_n3628.n65 9.3005
R20100 a_n1455_n3628.n53 a_n1455_n3628.n27 9.3005
R20101 a_n1455_n3628.n60 a_n1455_n3628.n29 9.3005
R20102 a_n1455_n3628.n29 a_n1455_n3628.n59 9.3005
R20103 a_n1455_n3628.n100 a_n1455_n3628.n99 9.3005
R20104 a_n1455_n3628.n78 a_n1455_n3628.n31 9.3005
R20105 a_n1455_n3628.n94 a_n1455_n3628.n31 9.3005
R20106 a_n1455_n3628.n30 a_n1455_n3628.n93 9.3005
R20107 a_n1455_n3628.n81 a_n1455_n3628.n30 9.3005
R20108 a_n1455_n3628.n88 a_n1455_n3628.n32 9.3005
R20109 a_n1455_n3628.n32 a_n1455_n3628.n87 9.3005
R20110 a_n1455_n3628.n126 a_n1455_n3628.n125 9.3005
R20111 a_n1455_n3628.n104 a_n1455_n3628.n34 9.3005
R20112 a_n1455_n3628.n120 a_n1455_n3628.n34 9.3005
R20113 a_n1455_n3628.n33 a_n1455_n3628.n119 9.3005
R20114 a_n1455_n3628.n107 a_n1455_n3628.n33 9.3005
R20115 a_n1455_n3628.n114 a_n1455_n3628.n35 9.3005
R20116 a_n1455_n3628.n35 a_n1455_n3628.n113 9.3005
R20117 a_n1455_n3628.n154 a_n1455_n3628.n153 9.3005
R20118 a_n1455_n3628.n132 a_n1455_n3628.n37 9.3005
R20119 a_n1455_n3628.n148 a_n1455_n3628.n37 9.3005
R20120 a_n1455_n3628.n36 a_n1455_n3628.n147 9.3005
R20121 a_n1455_n3628.n135 a_n1455_n3628.n36 9.3005
R20122 a_n1455_n3628.n142 a_n1455_n3628.n38 9.3005
R20123 a_n1455_n3628.n38 a_n1455_n3628.n141 9.3005
R20124 a_n1455_n3628.n342 a_n1455_n3628.n1 9.3005
R20125 a_n1455_n3628.n45 a_n1455_n3628.n1 9.3005
R20126 a_n1455_n3628.n2 a_n1455_n3628.n347 9.3005
R20127 a_n1455_n3628.n348 a_n1455_n3628.n2 9.3005
R20128 a_n1455_n3628.n42 a_n1455_n3628.n0 9.3005
R20129 a_n1455_n3628.n0 a_n1455_n3628.n353 9.3005
R20130 a_n1455_n3628.n355 a_n1455_n3628.n354 9.3005
R20131 a_n1455_n3628.n309 a_n1455_n3628.n289 8.92171
R20132 a_n1455_n3628.n336 a_n1455_n3628.n316 8.92171
R20133 a_n1455_n3628.n178 a_n1455_n3628.n158 8.92171
R20134 a_n1455_n3628.n282 a_n1455_n3628.n262 8.92171
R20135 a_n1455_n3628.n256 a_n1455_n3628.n236 8.92171
R20136 a_n1455_n3628.n230 a_n1455_n3628.n210 8.92171
R20137 a_n1455_n3628.n204 a_n1455_n3628.n184 8.92171
R20138 a_n1455_n3628.n70 a_n1455_n3628.n50 8.92171
R20139 a_n1455_n3628.n98 a_n1455_n3628.n78 8.92171
R20140 a_n1455_n3628.n124 a_n1455_n3628.n104 8.92171
R20141 a_n1455_n3628.n152 a_n1455_n3628.n132 8.92171
R20142 a_n1455_n3628.n343 a_n1455_n3628.n45 8.92171
R20143 a_n1455_n3628.n310 a_n1455_n3628.n288 8.14595
R20144 a_n1455_n3628.n337 a_n1455_n3628.n315 8.14595
R20145 a_n1455_n3628.n179 a_n1455_n3628.n157 8.14595
R20146 a_n1455_n3628.n283 a_n1455_n3628.n261 8.14595
R20147 a_n1455_n3628.n257 a_n1455_n3628.n235 8.14595
R20148 a_n1455_n3628.n231 a_n1455_n3628.n209 8.14595
R20149 a_n1455_n3628.n205 a_n1455_n3628.n183 8.14595
R20150 a_n1455_n3628.n71 a_n1455_n3628.n49 8.14595
R20151 a_n1455_n3628.n99 a_n1455_n3628.n77 8.14595
R20152 a_n1455_n3628.n125 a_n1455_n3628.n103 8.14595
R20153 a_n1455_n3628.n153 a_n1455_n3628.n131 8.14595
R20154 a_n1455_n3628.n342 a_n1455_n3628.n46 8.14595
R20155 a_n1455_n3628.n311 a_n1455_n3628.n288 5.81868
R20156 a_n1455_n3628.n338 a_n1455_n3628.n315 5.81868
R20157 a_n1455_n3628.n180 a_n1455_n3628.n157 5.81868
R20158 a_n1455_n3628.n285 a_n1455_n3628.n261 5.81868
R20159 a_n1455_n3628.n259 a_n1455_n3628.n235 5.81868
R20160 a_n1455_n3628.n233 a_n1455_n3628.n209 5.81868
R20161 a_n1455_n3628.n207 a_n1455_n3628.n183 5.81868
R20162 a_n1455_n3628.n73 a_n1455_n3628.n49 5.81868
R20163 a_n1455_n3628.n101 a_n1455_n3628.n77 5.81868
R20164 a_n1455_n3628.n127 a_n1455_n3628.n103 5.81868
R20165 a_n1455_n3628.n155 a_n1455_n3628.n131 5.81868
R20166 a_n1455_n3628.n341 a_n1455_n3628.n46 5.81868
R20167 a_n1455_n3628.n182 a_n1455_n3628.n181 5.18369
R20168 a_n1455_n3628.n312 a_n1455_n3628.n287 5.18369
R20169 a_n1455_n3628.n310 a_n1455_n3628.n309 5.04292
R20170 a_n1455_n3628.n337 a_n1455_n3628.n336 5.04292
R20171 a_n1455_n3628.n179 a_n1455_n3628.n178 5.04292
R20172 a_n1455_n3628.n283 a_n1455_n3628.n282 5.04292
R20173 a_n1455_n3628.n257 a_n1455_n3628.n256 5.04292
R20174 a_n1455_n3628.n231 a_n1455_n3628.n230 5.04292
R20175 a_n1455_n3628.n205 a_n1455_n3628.n204 5.04292
R20176 a_n1455_n3628.n71 a_n1455_n3628.n70 5.04292
R20177 a_n1455_n3628.n99 a_n1455_n3628.n98 5.04292
R20178 a_n1455_n3628.n125 a_n1455_n3628.n124 5.04292
R20179 a_n1455_n3628.n153 a_n1455_n3628.n152 5.04292
R20180 a_n1455_n3628.n343 a_n1455_n3628.n342 5.04292
R20181 a_n1455_n3628.n354 a_n1455_n3628.n39 4.38594
R20182 a_n1455_n3628.n3 a_n1455_n3628.n295 4.38594
R20183 a_n1455_n3628.n7 a_n1455_n3628.n322 4.38594
R20184 a_n1455_n3628.n11 a_n1455_n3628.n164 4.38594
R20185 a_n1455_n3628.n17 a_n1455_n3628.n268 4.38594
R20186 a_n1455_n3628.n20 a_n1455_n3628.n242 4.38594
R20187 a_n1455_n3628.n23 a_n1455_n3628.n216 4.38594
R20188 a_n1455_n3628.n26 a_n1455_n3628.n190 4.38594
R20189 a_n1455_n3628.n29 a_n1455_n3628.n56 4.38594
R20190 a_n1455_n3628.n32 a_n1455_n3628.n84 4.38594
R20191 a_n1455_n3628.n35 a_n1455_n3628.n110 4.38594
R20192 a_n1455_n3628.n38 a_n1455_n3628.n138 4.38594
R20193 a_n1455_n3628.n306 a_n1455_n3628.n289 4.26717
R20194 a_n1455_n3628.n333 a_n1455_n3628.n316 4.26717
R20195 a_n1455_n3628.n175 a_n1455_n3628.n158 4.26717
R20196 a_n1455_n3628.n279 a_n1455_n3628.n262 4.26717
R20197 a_n1455_n3628.n253 a_n1455_n3628.n236 4.26717
R20198 a_n1455_n3628.n227 a_n1455_n3628.n210 4.26717
R20199 a_n1455_n3628.n201 a_n1455_n3628.n184 4.26717
R20200 a_n1455_n3628.n67 a_n1455_n3628.n50 4.26717
R20201 a_n1455_n3628.n95 a_n1455_n3628.n78 4.26717
R20202 a_n1455_n3628.n121 a_n1455_n3628.n104 4.26717
R20203 a_n1455_n3628.n149 a_n1455_n3628.n132 4.26717
R20204 a_n1455_n3628.n346 a_n1455_n3628.n45 4.26717
R20205 a_n1455_n3628.n305 a_n1455_n3628.n291 3.49141
R20206 a_n1455_n3628.n332 a_n1455_n3628.n318 3.49141
R20207 a_n1455_n3628.n174 a_n1455_n3628.n160 3.49141
R20208 a_n1455_n3628.n278 a_n1455_n3628.n264 3.49141
R20209 a_n1455_n3628.n252 a_n1455_n3628.n238 3.49141
R20210 a_n1455_n3628.n226 a_n1455_n3628.n212 3.49141
R20211 a_n1455_n3628.n200 a_n1455_n3628.n186 3.49141
R20212 a_n1455_n3628.n66 a_n1455_n3628.n52 3.49141
R20213 a_n1455_n3628.n94 a_n1455_n3628.n80 3.49141
R20214 a_n1455_n3628.n120 a_n1455_n3628.n106 3.49141
R20215 a_n1455_n3628.n148 a_n1455_n3628.n134 3.49141
R20216 a_n1455_n3628.n347 a_n1455_n3628.n44 3.49141
R20217 a_n1455_n3628.n313 a_n1455_n3628.t16 3.3005
R20218 a_n1455_n3628.n313 a_n1455_n3628.t10 3.3005
R20219 a_n1455_n3628.n47 a_n1455_n3628.t4 3.3005
R20220 a_n1455_n3628.n47 a_n1455_n3628.t0 3.3005
R20221 a_n1455_n3628.n75 a_n1455_n3628.t6 3.3005
R20222 a_n1455_n3628.n75 a_n1455_n3628.t1 3.3005
R20223 a_n1455_n3628.n129 a_n1455_n3628.t8 3.3005
R20224 a_n1455_n3628.n129 a_n1455_n3628.t19 3.3005
R20225 a_n1455_n3628.n304 a_n1455_n3628.n303 2.71565
R20226 a_n1455_n3628.n331 a_n1455_n3628.n330 2.71565
R20227 a_n1455_n3628.n173 a_n1455_n3628.n172 2.71565
R20228 a_n1455_n3628.n277 a_n1455_n3628.n276 2.71565
R20229 a_n1455_n3628.n251 a_n1455_n3628.n250 2.71565
R20230 a_n1455_n3628.n225 a_n1455_n3628.n224 2.71565
R20231 a_n1455_n3628.n199 a_n1455_n3628.n198 2.71565
R20232 a_n1455_n3628.n65 a_n1455_n3628.n64 2.71565
R20233 a_n1455_n3628.n93 a_n1455_n3628.n92 2.71565
R20234 a_n1455_n3628.n119 a_n1455_n3628.n118 2.71565
R20235 a_n1455_n3628.n147 a_n1455_n3628.n146 2.71565
R20236 a_n1455_n3628.n349 a_n1455_n3628.n348 2.71565
R20237 a_n1455_n3628.n287 a_n1455_n3628.n286 2.23674
R20238 a_n1455_n3628.n208 a_n1455_n3628.n182 1.95694
R20239 a_n1455_n3628.n300 a_n1455_n3628.n292 1.93989
R20240 a_n1455_n3628.n327 a_n1455_n3628.n319 1.93989
R20241 a_n1455_n3628.n169 a_n1455_n3628.n161 1.93989
R20242 a_n1455_n3628.n273 a_n1455_n3628.n265 1.93989
R20243 a_n1455_n3628.n247 a_n1455_n3628.n239 1.93989
R20244 a_n1455_n3628.n221 a_n1455_n3628.n213 1.93989
R20245 a_n1455_n3628.n195 a_n1455_n3628.n187 1.93989
R20246 a_n1455_n3628.n61 a_n1455_n3628.n53 1.93989
R20247 a_n1455_n3628.n89 a_n1455_n3628.n81 1.93989
R20248 a_n1455_n3628.n115 a_n1455_n3628.n107 1.93989
R20249 a_n1455_n3628.n143 a_n1455_n3628.n135 1.93989
R20250 a_n1455_n3628.n352 a_n1455_n3628.n42 1.93989
R20251 a_n1455_n3628.n299 a_n1455_n3628.n294 1.16414
R20252 a_n1455_n3628.n326 a_n1455_n3628.n321 1.16414
R20253 a_n1455_n3628.n168 a_n1455_n3628.n163 1.16414
R20254 a_n1455_n3628.n272 a_n1455_n3628.n267 1.16414
R20255 a_n1455_n3628.n246 a_n1455_n3628.n241 1.16414
R20256 a_n1455_n3628.n220 a_n1455_n3628.n215 1.16414
R20257 a_n1455_n3628.n194 a_n1455_n3628.n189 1.16414
R20258 a_n1455_n3628.n60 a_n1455_n3628.n55 1.16414
R20259 a_n1455_n3628.n88 a_n1455_n3628.n83 1.16414
R20260 a_n1455_n3628.n114 a_n1455_n3628.n109 1.16414
R20261 a_n1455_n3628.n142 a_n1455_n3628.n137 1.16414
R20262 a_n1455_n3628.n353 a_n1455_n3628.n41 1.16414
R20263 a_n1455_n3628.n260 a_n1455_n3628.n234 0.962709
R20264 a_n1455_n3628.n286 a_n1455_n3628.n260 0.962709
R20265 a_n1455_n3628.n156 a_n1455_n3628.n130 0.573776
R20266 a_n1455_n3628.n130 a_n1455_n3628.n128 0.573776
R20267 a_n1455_n3628.n102 a_n1455_n3628.n76 0.573776
R20268 a_n1455_n3628.n76 a_n1455_n3628.n74 0.573776
R20269 a_n1455_n3628.n181 a_n1455_n3628.n48 0.573776
R20270 a_n1455_n3628.n340 a_n1455_n3628.n48 0.573776
R20271 a_n1455_n3628.n339 a_n1455_n3628.n314 0.573776
R20272 a_n1455_n3628.n314 a_n1455_n3628.n312 0.573776
R20273 a_n1455_n3628.n234 a_n1455_n3628.n208 0.422738
R20274 a_n1455_n3628.n298 a_n1455_n3628.n297 0.388379
R20275 a_n1455_n3628.n325 a_n1455_n3628.n324 0.388379
R20276 a_n1455_n3628.n167 a_n1455_n3628.n166 0.388379
R20277 a_n1455_n3628.n271 a_n1455_n3628.n270 0.388379
R20278 a_n1455_n3628.n245 a_n1455_n3628.n244 0.388379
R20279 a_n1455_n3628.n219 a_n1455_n3628.n218 0.388379
R20280 a_n1455_n3628.n193 a_n1455_n3628.n192 0.388379
R20281 a_n1455_n3628.n59 a_n1455_n3628.n58 0.388379
R20282 a_n1455_n3628.n87 a_n1455_n3628.n86 0.388379
R20283 a_n1455_n3628.n113 a_n1455_n3628.n112 0.388379
R20284 a_n1455_n3628.n141 a_n1455_n3628.n140 0.388379
R20285 a_n1455_n3628.n356 a_n1455_n3628.n355 0.388379
R20286 a_n1455_n3628.n38 a_n1455_n3628.n36 0.310845
R20287 a_n1455_n3628.n37 a_n1455_n3628.n36 0.310845
R20288 a_n1455_n3628.n154 a_n1455_n3628.n37 0.310845
R20289 a_n1455_n3628.n35 a_n1455_n3628.n33 0.310845
R20290 a_n1455_n3628.n34 a_n1455_n3628.n33 0.310845
R20291 a_n1455_n3628.n126 a_n1455_n3628.n34 0.310845
R20292 a_n1455_n3628.n32 a_n1455_n3628.n30 0.310845
R20293 a_n1455_n3628.n31 a_n1455_n3628.n30 0.310845
R20294 a_n1455_n3628.n100 a_n1455_n3628.n31 0.310845
R20295 a_n1455_n3628.n29 a_n1455_n3628.n27 0.310845
R20296 a_n1455_n3628.n28 a_n1455_n3628.n27 0.310845
R20297 a_n1455_n3628.n72 a_n1455_n3628.n28 0.310845
R20298 a_n1455_n3628.n26 a_n1455_n3628.n24 0.310845
R20299 a_n1455_n3628.n25 a_n1455_n3628.n24 0.310845
R20300 a_n1455_n3628.n206 a_n1455_n3628.n25 0.310845
R20301 a_n1455_n3628.n23 a_n1455_n3628.n21 0.310845
R20302 a_n1455_n3628.n22 a_n1455_n3628.n21 0.310845
R20303 a_n1455_n3628.n232 a_n1455_n3628.n22 0.310845
R20304 a_n1455_n3628.n20 a_n1455_n3628.n18 0.310845
R20305 a_n1455_n3628.n19 a_n1455_n3628.n18 0.310845
R20306 a_n1455_n3628.n258 a_n1455_n3628.n19 0.310845
R20307 a_n1455_n3628.n17 a_n1455_n3628.n15 0.310845
R20308 a_n1455_n3628.n16 a_n1455_n3628.n15 0.310845
R20309 a_n1455_n3628.n284 a_n1455_n3628.n16 0.310845
R20310 a_n1455_n3628.n14 a_n1455_n3628.n13 0.310845
R20311 a_n1455_n3628.n14 a_n1455_n3628.n12 0.310845
R20312 a_n1455_n3628.n12 a_n1455_n3628.n11 0.310845
R20313 a_n1455_n3628.n10 a_n1455_n3628.n9 0.310845
R20314 a_n1455_n3628.n10 a_n1455_n3628.n8 0.310845
R20315 a_n1455_n3628.n8 a_n1455_n3628.n7 0.310845
R20316 a_n1455_n3628.n6 a_n1455_n3628.n5 0.310845
R20317 a_n1455_n3628.n6 a_n1455_n3628.n4 0.310845
R20318 a_n1455_n3628.n4 a_n1455_n3628.n3 0.310845
R20319 a_n1455_n3628.n2 a_n1455_n3628.n1 0.310845
R20320 a_n1455_n3628.n2 a_n1455_n3628.n0 0.310845
R20321 a_n1455_n3628.n354 a_n1455_n3628.n0 0.310845
R20322 a_n1455_n3628.n128 a_n1455_n3628.n102 0.235414
R20323 a_n1455_n3628.n340 a_n1455_n3628.n339 0.235414
R20324 VP.n30 VP.t3 243.255
R20325 VP.n29 VP.n27 224.169
R20326 VP.n29 VP.n28 223.454
R20327 VP.n15 VP.t9 199.144
R20328 VP.n2 VP.t11 199.144
R20329 VP.n24 VP.t7 183.883
R20330 VP.n11 VP.t5 183.883
R20331 VP.n18 VP.n17 161.3
R20332 VP.n19 VP.n14 161.3
R20333 VP.n21 VP.n20 161.3
R20334 VP.n23 VP.n13 161.3
R20335 VP.n10 VP.n0 161.3
R20336 VP.n8 VP.n7 161.3
R20337 VP.n6 VP.n1 161.3
R20338 VP.n5 VP.n4 161.3
R20339 VP.n22 VP.t12 144.601
R20340 VP.n16 VP.t8 144.601
R20341 VP.n3 VP.t10 144.601
R20342 VP.n9 VP.t6 144.601
R20343 VP.n25 VP.n24 80.6037
R20344 VP.n12 VP.n11 80.6037
R20345 VP.n24 VP.n23 56.3158
R20346 VP.n11 VP.n10 56.3158
R20347 VP.n16 VP.n15 46.9082
R20348 VP.n3 VP.n2 46.9082
R20349 VP.n5 VP.n2 43.8991
R20350 VP.n18 VP.n15 43.8991
R20351 VP.n21 VP.n14 40.577
R20352 VP.n17 VP.n14 40.577
R20353 VP.n4 VP.n1 40.577
R20354 VP.n8 VP.n1 40.577
R20355 VP.n26 VP.n25 28.1089
R20356 VP.n28 VP.t0 19.8005
R20357 VP.n28 VP.t2 19.8005
R20358 VP.n27 VP.t4 19.8005
R20359 VP.n27 VP.t1 19.8005
R20360 VP.n23 VP.n22 16.477
R20361 VP.n10 VP.n9 16.477
R20362 VP.n26 VP.n12 11.9157
R20363 VP VP.n31 11.8187
R20364 VP.n22 VP.n21 8.11581
R20365 VP.n17 VP.n16 8.11581
R20366 VP.n4 VP.n3 8.11581
R20367 VP.n9 VP.n8 8.11581
R20368 VP.n31 VP.n30 4.80222
R20369 VP.n31 VP.n26 0.972091
R20370 VP.n30 VP.n29 0.716017
R20371 VP.n25 VP.n13 0.285035
R20372 VP.n12 VP.n0 0.285035
R20373 VP.n20 VP.n13 0.189894
R20374 VP.n20 VP.n19 0.189894
R20375 VP.n19 VP.n18 0.189894
R20376 VP.n6 VP.n5 0.189894
R20377 VP.n7 VP.n6 0.189894
R20378 VP.n7 VP.n0 0.189894
R20379 DIFFPAIR_BIAS.n27 DIFFPAIR_BIAS.n1 289.615
R20380 DIFFPAIR_BIAS.n58 DIFFPAIR_BIAS.n32 289.615
R20381 DIFFPAIR_BIAS.n90 DIFFPAIR_BIAS.n64 289.615
R20382 DIFFPAIR_BIAS.n122 DIFFPAIR_BIAS.n96 289.615
R20383 DIFFPAIR_BIAS.n28 DIFFPAIR_BIAS.n27 185
R20384 DIFFPAIR_BIAS.n26 DIFFPAIR_BIAS.n25 185
R20385 DIFFPAIR_BIAS.n5 DIFFPAIR_BIAS.n4 185
R20386 DIFFPAIR_BIAS.n20 DIFFPAIR_BIAS.n19 185
R20387 DIFFPAIR_BIAS.n18 DIFFPAIR_BIAS.n17 185
R20388 DIFFPAIR_BIAS.n9 DIFFPAIR_BIAS.n8 185
R20389 DIFFPAIR_BIAS.n12 DIFFPAIR_BIAS.n11 185
R20390 DIFFPAIR_BIAS.n59 DIFFPAIR_BIAS.n58 185
R20391 DIFFPAIR_BIAS.n57 DIFFPAIR_BIAS.n56 185
R20392 DIFFPAIR_BIAS.n36 DIFFPAIR_BIAS.n35 185
R20393 DIFFPAIR_BIAS.n51 DIFFPAIR_BIAS.n50 185
R20394 DIFFPAIR_BIAS.n49 DIFFPAIR_BIAS.n48 185
R20395 DIFFPAIR_BIAS.n40 DIFFPAIR_BIAS.n39 185
R20396 DIFFPAIR_BIAS.n43 DIFFPAIR_BIAS.n42 185
R20397 DIFFPAIR_BIAS.n91 DIFFPAIR_BIAS.n90 185
R20398 DIFFPAIR_BIAS.n89 DIFFPAIR_BIAS.n88 185
R20399 DIFFPAIR_BIAS.n68 DIFFPAIR_BIAS.n67 185
R20400 DIFFPAIR_BIAS.n83 DIFFPAIR_BIAS.n82 185
R20401 DIFFPAIR_BIAS.n81 DIFFPAIR_BIAS.n80 185
R20402 DIFFPAIR_BIAS.n72 DIFFPAIR_BIAS.n71 185
R20403 DIFFPAIR_BIAS.n75 DIFFPAIR_BIAS.n74 185
R20404 DIFFPAIR_BIAS.n123 DIFFPAIR_BIAS.n122 185
R20405 DIFFPAIR_BIAS.n121 DIFFPAIR_BIAS.n120 185
R20406 DIFFPAIR_BIAS.n100 DIFFPAIR_BIAS.n99 185
R20407 DIFFPAIR_BIAS.n115 DIFFPAIR_BIAS.n114 185
R20408 DIFFPAIR_BIAS.n113 DIFFPAIR_BIAS.n112 185
R20409 DIFFPAIR_BIAS.n104 DIFFPAIR_BIAS.n103 185
R20410 DIFFPAIR_BIAS.n107 DIFFPAIR_BIAS.n106 185
R20411 DIFFPAIR_BIAS.n0 DIFFPAIR_BIAS.t9 178.945
R20412 DIFFPAIR_BIAS.n133 DIFFPAIR_BIAS.t10 177.018
R20413 DIFFPAIR_BIAS.n132 DIFFPAIR_BIAS.t11 177.018
R20414 DIFFPAIR_BIAS.n0 DIFFPAIR_BIAS.t8 177.018
R20415 DIFFPAIR_BIAS.t1 DIFFPAIR_BIAS.n10 147.661
R20416 DIFFPAIR_BIAS.t3 DIFFPAIR_BIAS.n41 147.661
R20417 DIFFPAIR_BIAS.t5 DIFFPAIR_BIAS.n73 147.661
R20418 DIFFPAIR_BIAS.t7 DIFFPAIR_BIAS.n105 147.661
R20419 DIFFPAIR_BIAS.n128 DIFFPAIR_BIAS.t0 132.363
R20420 DIFFPAIR_BIAS.n128 DIFFPAIR_BIAS.t2 130.436
R20421 DIFFPAIR_BIAS.n129 DIFFPAIR_BIAS.t4 130.436
R20422 DIFFPAIR_BIAS.n130 DIFFPAIR_BIAS.t6 130.436
R20423 DIFFPAIR_BIAS.n27 DIFFPAIR_BIAS.n26 104.615
R20424 DIFFPAIR_BIAS.n26 DIFFPAIR_BIAS.n4 104.615
R20425 DIFFPAIR_BIAS.n19 DIFFPAIR_BIAS.n4 104.615
R20426 DIFFPAIR_BIAS.n19 DIFFPAIR_BIAS.n18 104.615
R20427 DIFFPAIR_BIAS.n18 DIFFPAIR_BIAS.n8 104.615
R20428 DIFFPAIR_BIAS.n11 DIFFPAIR_BIAS.n8 104.615
R20429 DIFFPAIR_BIAS.n58 DIFFPAIR_BIAS.n57 104.615
R20430 DIFFPAIR_BIAS.n57 DIFFPAIR_BIAS.n35 104.615
R20431 DIFFPAIR_BIAS.n50 DIFFPAIR_BIAS.n35 104.615
R20432 DIFFPAIR_BIAS.n50 DIFFPAIR_BIAS.n49 104.615
R20433 DIFFPAIR_BIAS.n49 DIFFPAIR_BIAS.n39 104.615
R20434 DIFFPAIR_BIAS.n42 DIFFPAIR_BIAS.n39 104.615
R20435 DIFFPAIR_BIAS.n90 DIFFPAIR_BIAS.n89 104.615
R20436 DIFFPAIR_BIAS.n89 DIFFPAIR_BIAS.n67 104.615
R20437 DIFFPAIR_BIAS.n82 DIFFPAIR_BIAS.n67 104.615
R20438 DIFFPAIR_BIAS.n82 DIFFPAIR_BIAS.n81 104.615
R20439 DIFFPAIR_BIAS.n81 DIFFPAIR_BIAS.n71 104.615
R20440 DIFFPAIR_BIAS.n74 DIFFPAIR_BIAS.n71 104.615
R20441 DIFFPAIR_BIAS.n122 DIFFPAIR_BIAS.n121 104.615
R20442 DIFFPAIR_BIAS.n121 DIFFPAIR_BIAS.n99 104.615
R20443 DIFFPAIR_BIAS.n114 DIFFPAIR_BIAS.n99 104.615
R20444 DIFFPAIR_BIAS.n114 DIFFPAIR_BIAS.n113 104.615
R20445 DIFFPAIR_BIAS.n113 DIFFPAIR_BIAS.n103 104.615
R20446 DIFFPAIR_BIAS.n106 DIFFPAIR_BIAS.n103 104.615
R20447 DIFFPAIR_BIAS.n63 DIFFPAIR_BIAS.n31 95.6354
R20448 DIFFPAIR_BIAS.n63 DIFFPAIR_BIAS.n62 94.6732
R20449 DIFFPAIR_BIAS.n95 DIFFPAIR_BIAS.n94 94.6732
R20450 DIFFPAIR_BIAS.n127 DIFFPAIR_BIAS.n126 94.6732
R20451 DIFFPAIR_BIAS.n11 DIFFPAIR_BIAS.t1 52.3082
R20452 DIFFPAIR_BIAS.n42 DIFFPAIR_BIAS.t3 52.3082
R20453 DIFFPAIR_BIAS.n74 DIFFPAIR_BIAS.t5 52.3082
R20454 DIFFPAIR_BIAS.n106 DIFFPAIR_BIAS.t7 52.3082
R20455 DIFFPAIR_BIAS.n12 DIFFPAIR_BIAS.n10 15.6674
R20456 DIFFPAIR_BIAS.n43 DIFFPAIR_BIAS.n41 15.6674
R20457 DIFFPAIR_BIAS.n75 DIFFPAIR_BIAS.n73 15.6674
R20458 DIFFPAIR_BIAS.n107 DIFFPAIR_BIAS.n105 15.6674
R20459 DIFFPAIR_BIAS.n13 DIFFPAIR_BIAS.n9 12.8005
R20460 DIFFPAIR_BIAS.n44 DIFFPAIR_BIAS.n40 12.8005
R20461 DIFFPAIR_BIAS.n76 DIFFPAIR_BIAS.n72 12.8005
R20462 DIFFPAIR_BIAS.n108 DIFFPAIR_BIAS.n104 12.8005
R20463 DIFFPAIR_BIAS.n17 DIFFPAIR_BIAS.n16 12.0247
R20464 DIFFPAIR_BIAS.n48 DIFFPAIR_BIAS.n47 12.0247
R20465 DIFFPAIR_BIAS.n80 DIFFPAIR_BIAS.n79 12.0247
R20466 DIFFPAIR_BIAS.n112 DIFFPAIR_BIAS.n111 12.0247
R20467 DIFFPAIR_BIAS.n20 DIFFPAIR_BIAS.n7 11.249
R20468 DIFFPAIR_BIAS.n51 DIFFPAIR_BIAS.n38 11.249
R20469 DIFFPAIR_BIAS.n83 DIFFPAIR_BIAS.n70 11.249
R20470 DIFFPAIR_BIAS.n115 DIFFPAIR_BIAS.n102 11.249
R20471 DIFFPAIR_BIAS.n21 DIFFPAIR_BIAS.n5 10.4732
R20472 DIFFPAIR_BIAS.n52 DIFFPAIR_BIAS.n36 10.4732
R20473 DIFFPAIR_BIAS.n84 DIFFPAIR_BIAS.n68 10.4732
R20474 DIFFPAIR_BIAS.n116 DIFFPAIR_BIAS.n100 10.4732
R20475 DIFFPAIR_BIAS.n25 DIFFPAIR_BIAS.n24 9.69747
R20476 DIFFPAIR_BIAS.n56 DIFFPAIR_BIAS.n55 9.69747
R20477 DIFFPAIR_BIAS.n88 DIFFPAIR_BIAS.n87 9.69747
R20478 DIFFPAIR_BIAS.n120 DIFFPAIR_BIAS.n119 9.69747
R20479 DIFFPAIR_BIAS.n31 DIFFPAIR_BIAS.n30 9.45567
R20480 DIFFPAIR_BIAS.n62 DIFFPAIR_BIAS.n61 9.45567
R20481 DIFFPAIR_BIAS.n94 DIFFPAIR_BIAS.n93 9.45567
R20482 DIFFPAIR_BIAS.n126 DIFFPAIR_BIAS.n125 9.45567
R20483 DIFFPAIR_BIAS.n30 DIFFPAIR_BIAS.n29 9.3005
R20484 DIFFPAIR_BIAS.n3 DIFFPAIR_BIAS.n2 9.3005
R20485 DIFFPAIR_BIAS.n24 DIFFPAIR_BIAS.n23 9.3005
R20486 DIFFPAIR_BIAS.n22 DIFFPAIR_BIAS.n21 9.3005
R20487 DIFFPAIR_BIAS.n7 DIFFPAIR_BIAS.n6 9.3005
R20488 DIFFPAIR_BIAS.n16 DIFFPAIR_BIAS.n15 9.3005
R20489 DIFFPAIR_BIAS.n14 DIFFPAIR_BIAS.n13 9.3005
R20490 DIFFPAIR_BIAS.n61 DIFFPAIR_BIAS.n60 9.3005
R20491 DIFFPAIR_BIAS.n34 DIFFPAIR_BIAS.n33 9.3005
R20492 DIFFPAIR_BIAS.n55 DIFFPAIR_BIAS.n54 9.3005
R20493 DIFFPAIR_BIAS.n53 DIFFPAIR_BIAS.n52 9.3005
R20494 DIFFPAIR_BIAS.n38 DIFFPAIR_BIAS.n37 9.3005
R20495 DIFFPAIR_BIAS.n47 DIFFPAIR_BIAS.n46 9.3005
R20496 DIFFPAIR_BIAS.n45 DIFFPAIR_BIAS.n44 9.3005
R20497 DIFFPAIR_BIAS.n93 DIFFPAIR_BIAS.n92 9.3005
R20498 DIFFPAIR_BIAS.n66 DIFFPAIR_BIAS.n65 9.3005
R20499 DIFFPAIR_BIAS.n87 DIFFPAIR_BIAS.n86 9.3005
R20500 DIFFPAIR_BIAS.n85 DIFFPAIR_BIAS.n84 9.3005
R20501 DIFFPAIR_BIAS.n70 DIFFPAIR_BIAS.n69 9.3005
R20502 DIFFPAIR_BIAS.n79 DIFFPAIR_BIAS.n78 9.3005
R20503 DIFFPAIR_BIAS.n77 DIFFPAIR_BIAS.n76 9.3005
R20504 DIFFPAIR_BIAS.n125 DIFFPAIR_BIAS.n124 9.3005
R20505 DIFFPAIR_BIAS.n98 DIFFPAIR_BIAS.n97 9.3005
R20506 DIFFPAIR_BIAS.n119 DIFFPAIR_BIAS.n118 9.3005
R20507 DIFFPAIR_BIAS.n117 DIFFPAIR_BIAS.n116 9.3005
R20508 DIFFPAIR_BIAS.n102 DIFFPAIR_BIAS.n101 9.3005
R20509 DIFFPAIR_BIAS.n111 DIFFPAIR_BIAS.n110 9.3005
R20510 DIFFPAIR_BIAS.n109 DIFFPAIR_BIAS.n108 9.3005
R20511 DIFFPAIR_BIAS.n28 DIFFPAIR_BIAS.n3 8.92171
R20512 DIFFPAIR_BIAS.n59 DIFFPAIR_BIAS.n34 8.92171
R20513 DIFFPAIR_BIAS.n91 DIFFPAIR_BIAS.n66 8.92171
R20514 DIFFPAIR_BIAS.n123 DIFFPAIR_BIAS.n98 8.92171
R20515 DIFFPAIR_BIAS.n29 DIFFPAIR_BIAS.n1 8.14595
R20516 DIFFPAIR_BIAS.n60 DIFFPAIR_BIAS.n32 8.14595
R20517 DIFFPAIR_BIAS.n92 DIFFPAIR_BIAS.n64 8.14595
R20518 DIFFPAIR_BIAS.n124 DIFFPAIR_BIAS.n96 8.14595
R20519 DIFFPAIR_BIAS.n31 DIFFPAIR_BIAS.n1 5.81868
R20520 DIFFPAIR_BIAS.n62 DIFFPAIR_BIAS.n32 5.81868
R20521 DIFFPAIR_BIAS.n94 DIFFPAIR_BIAS.n64 5.81868
R20522 DIFFPAIR_BIAS.n126 DIFFPAIR_BIAS.n96 5.81868
R20523 DIFFPAIR_BIAS.n131 DIFFPAIR_BIAS.n130 5.20947
R20524 DIFFPAIR_BIAS.n29 DIFFPAIR_BIAS.n28 5.04292
R20525 DIFFPAIR_BIAS.n60 DIFFPAIR_BIAS.n59 5.04292
R20526 DIFFPAIR_BIAS.n92 DIFFPAIR_BIAS.n91 5.04292
R20527 DIFFPAIR_BIAS.n124 DIFFPAIR_BIAS.n123 5.04292
R20528 DIFFPAIR_BIAS.n131 DIFFPAIR_BIAS.n127 4.42209
R20529 DIFFPAIR_BIAS.n14 DIFFPAIR_BIAS.n10 4.38594
R20530 DIFFPAIR_BIAS.n45 DIFFPAIR_BIAS.n41 4.38594
R20531 DIFFPAIR_BIAS.n77 DIFFPAIR_BIAS.n73 4.38594
R20532 DIFFPAIR_BIAS.n109 DIFFPAIR_BIAS.n105 4.38594
R20533 DIFFPAIR_BIAS.n132 DIFFPAIR_BIAS.n131 4.28454
R20534 DIFFPAIR_BIAS.n25 DIFFPAIR_BIAS.n3 4.26717
R20535 DIFFPAIR_BIAS.n56 DIFFPAIR_BIAS.n34 4.26717
R20536 DIFFPAIR_BIAS.n88 DIFFPAIR_BIAS.n66 4.26717
R20537 DIFFPAIR_BIAS.n120 DIFFPAIR_BIAS.n98 4.26717
R20538 DIFFPAIR_BIAS.n24 DIFFPAIR_BIAS.n5 3.49141
R20539 DIFFPAIR_BIAS.n55 DIFFPAIR_BIAS.n36 3.49141
R20540 DIFFPAIR_BIAS.n87 DIFFPAIR_BIAS.n68 3.49141
R20541 DIFFPAIR_BIAS.n119 DIFFPAIR_BIAS.n100 3.49141
R20542 DIFFPAIR_BIAS.n21 DIFFPAIR_BIAS.n20 2.71565
R20543 DIFFPAIR_BIAS.n52 DIFFPAIR_BIAS.n51 2.71565
R20544 DIFFPAIR_BIAS.n84 DIFFPAIR_BIAS.n83 2.71565
R20545 DIFFPAIR_BIAS.n116 DIFFPAIR_BIAS.n115 2.71565
R20546 DIFFPAIR_BIAS.n17 DIFFPAIR_BIAS.n7 1.93989
R20547 DIFFPAIR_BIAS.n48 DIFFPAIR_BIAS.n38 1.93989
R20548 DIFFPAIR_BIAS.n80 DIFFPAIR_BIAS.n70 1.93989
R20549 DIFFPAIR_BIAS.n112 DIFFPAIR_BIAS.n102 1.93989
R20550 DIFFPAIR_BIAS.n130 DIFFPAIR_BIAS.n129 1.9266
R20551 DIFFPAIR_BIAS.n129 DIFFPAIR_BIAS.n128 1.9266
R20552 DIFFPAIR_BIAS.n133 DIFFPAIR_BIAS.n132 1.92658
R20553 DIFFPAIR_BIAS.n134 DIFFPAIR_BIAS.n133 1.29913
R20554 DIFFPAIR_BIAS.n16 DIFFPAIR_BIAS.n9 1.16414
R20555 DIFFPAIR_BIAS.n47 DIFFPAIR_BIAS.n40 1.16414
R20556 DIFFPAIR_BIAS.n79 DIFFPAIR_BIAS.n72 1.16414
R20557 DIFFPAIR_BIAS.n111 DIFFPAIR_BIAS.n104 1.16414
R20558 DIFFPAIR_BIAS.n127 DIFFPAIR_BIAS.n95 0.962709
R20559 DIFFPAIR_BIAS.n95 DIFFPAIR_BIAS.n63 0.962709
R20560 DIFFPAIR_BIAS DIFFPAIR_BIAS.n134 0.684875
R20561 DIFFPAIR_BIAS.n13 DIFFPAIR_BIAS.n12 0.388379
R20562 DIFFPAIR_BIAS.n44 DIFFPAIR_BIAS.n43 0.388379
R20563 DIFFPAIR_BIAS.n76 DIFFPAIR_BIAS.n75 0.388379
R20564 DIFFPAIR_BIAS.n108 DIFFPAIR_BIAS.n107 0.388379
R20565 DIFFPAIR_BIAS.n134 DIFFPAIR_BIAS.n0 0.337251
R20566 DIFFPAIR_BIAS.n30 DIFFPAIR_BIAS.n2 0.155672
R20567 DIFFPAIR_BIAS.n23 DIFFPAIR_BIAS.n2 0.155672
R20568 DIFFPAIR_BIAS.n23 DIFFPAIR_BIAS.n22 0.155672
R20569 DIFFPAIR_BIAS.n22 DIFFPAIR_BIAS.n6 0.155672
R20570 DIFFPAIR_BIAS.n15 DIFFPAIR_BIAS.n6 0.155672
R20571 DIFFPAIR_BIAS.n15 DIFFPAIR_BIAS.n14 0.155672
R20572 DIFFPAIR_BIAS.n61 DIFFPAIR_BIAS.n33 0.155672
R20573 DIFFPAIR_BIAS.n54 DIFFPAIR_BIAS.n33 0.155672
R20574 DIFFPAIR_BIAS.n54 DIFFPAIR_BIAS.n53 0.155672
R20575 DIFFPAIR_BIAS.n53 DIFFPAIR_BIAS.n37 0.155672
R20576 DIFFPAIR_BIAS.n46 DIFFPAIR_BIAS.n37 0.155672
R20577 DIFFPAIR_BIAS.n46 DIFFPAIR_BIAS.n45 0.155672
R20578 DIFFPAIR_BIAS.n93 DIFFPAIR_BIAS.n65 0.155672
R20579 DIFFPAIR_BIAS.n86 DIFFPAIR_BIAS.n65 0.155672
R20580 DIFFPAIR_BIAS.n86 DIFFPAIR_BIAS.n85 0.155672
R20581 DIFFPAIR_BIAS.n85 DIFFPAIR_BIAS.n69 0.155672
R20582 DIFFPAIR_BIAS.n78 DIFFPAIR_BIAS.n69 0.155672
R20583 DIFFPAIR_BIAS.n78 DIFFPAIR_BIAS.n77 0.155672
R20584 DIFFPAIR_BIAS.n125 DIFFPAIR_BIAS.n97 0.155672
R20585 DIFFPAIR_BIAS.n118 DIFFPAIR_BIAS.n97 0.155672
R20586 DIFFPAIR_BIAS.n118 DIFFPAIR_BIAS.n117 0.155672
R20587 DIFFPAIR_BIAS.n117 DIFFPAIR_BIAS.n101 0.155672
R20588 DIFFPAIR_BIAS.n110 DIFFPAIR_BIAS.n101 0.155672
R20589 DIFFPAIR_BIAS.n110 DIFFPAIR_BIAS.n109 0.155672
C0 VDD VOUT 67.65f
C1 VOUT VP 2.98653f
C2 VDD VN 0.082744f
C3 VOUT VN 0.822022f
C4 VP VN 8.176241f
C5 VOUT CS_BIAS 30.840801f
C6 VP CS_BIAS 0.306594f
C7 VN CS_BIAS 0.266289f
C8 VP DIFFPAIR_BIAS 2.16e-19
C9 VN DIFFPAIR_BIAS 2.16e-19
C10 CS_BIAS DIFFPAIR_BIAS 0.009353f
C11 DIFFPAIR_BIAS GND 32.770004f
C12 CS_BIAS GND 0.139143p
C13 VN GND 26.44436f
C14 VP GND 23.48365f
C15 VOUT GND 70.25275f
C16 VDD GND 0.370346p
C17 DIFFPAIR_BIAS.t8 GND 0.108432f
C18 DIFFPAIR_BIAS.t9 GND 0.109185f
C19 DIFFPAIR_BIAS.n0 GND 0.122922f
C20 DIFFPAIR_BIAS.n1 GND 0.001296f
C21 DIFFPAIR_BIAS.n2 GND 9.22e-19
C22 DIFFPAIR_BIAS.n3 GND 4.95e-19
C23 DIFFPAIR_BIAS.n4 GND 0.001171f
C24 DIFFPAIR_BIAS.n5 GND 5.25e-19
C25 DIFFPAIR_BIAS.n6 GND 9.22e-19
C26 DIFFPAIR_BIAS.n7 GND 4.95e-19
C27 DIFFPAIR_BIAS.n8 GND 0.001171f
C28 DIFFPAIR_BIAS.n9 GND 5.25e-19
C29 DIFFPAIR_BIAS.n10 GND 0.003945f
C30 DIFFPAIR_BIAS.t1 GND 0.001909f
C31 DIFFPAIR_BIAS.n11 GND 8.78e-19
C32 DIFFPAIR_BIAS.n12 GND 6.92e-19
C33 DIFFPAIR_BIAS.n13 GND 4.95e-19
C34 DIFFPAIR_BIAS.n14 GND 0.021937f
C35 DIFFPAIR_BIAS.n15 GND 9.22e-19
C36 DIFFPAIR_BIAS.n16 GND 4.95e-19
C37 DIFFPAIR_BIAS.n17 GND 5.25e-19
C38 DIFFPAIR_BIAS.n18 GND 0.001171f
C39 DIFFPAIR_BIAS.n19 GND 0.001171f
C40 DIFFPAIR_BIAS.n20 GND 5.25e-19
C41 DIFFPAIR_BIAS.n21 GND 4.95e-19
C42 DIFFPAIR_BIAS.n22 GND 9.22e-19
C43 DIFFPAIR_BIAS.n23 GND 9.22e-19
C44 DIFFPAIR_BIAS.n24 GND 4.95e-19
C45 DIFFPAIR_BIAS.n25 GND 5.25e-19
C46 DIFFPAIR_BIAS.n26 GND 0.001171f
C47 DIFFPAIR_BIAS.n27 GND 0.002535f
C48 DIFFPAIR_BIAS.n28 GND 5.25e-19
C49 DIFFPAIR_BIAS.n29 GND 4.95e-19
C50 DIFFPAIR_BIAS.n30 GND 0.002131f
C51 DIFFPAIR_BIAS.n31 GND 0.005461f
C52 DIFFPAIR_BIAS.n32 GND 0.001296f
C53 DIFFPAIR_BIAS.n33 GND 9.22e-19
C54 DIFFPAIR_BIAS.n34 GND 4.95e-19
C55 DIFFPAIR_BIAS.n35 GND 0.001171f
C56 DIFFPAIR_BIAS.n36 GND 5.25e-19
C57 DIFFPAIR_BIAS.n37 GND 9.22e-19
C58 DIFFPAIR_BIAS.n38 GND 4.95e-19
C59 DIFFPAIR_BIAS.n39 GND 0.001171f
C60 DIFFPAIR_BIAS.n40 GND 5.25e-19
C61 DIFFPAIR_BIAS.n41 GND 0.003945f
C62 DIFFPAIR_BIAS.t3 GND 0.001909f
C63 DIFFPAIR_BIAS.n42 GND 8.78e-19
C64 DIFFPAIR_BIAS.n43 GND 6.92e-19
C65 DIFFPAIR_BIAS.n44 GND 4.95e-19
C66 DIFFPAIR_BIAS.n45 GND 0.021937f
C67 DIFFPAIR_BIAS.n46 GND 9.22e-19
C68 DIFFPAIR_BIAS.n47 GND 4.95e-19
C69 DIFFPAIR_BIAS.n48 GND 5.25e-19
C70 DIFFPAIR_BIAS.n49 GND 0.001171f
C71 DIFFPAIR_BIAS.n50 GND 0.001171f
C72 DIFFPAIR_BIAS.n51 GND 5.25e-19
C73 DIFFPAIR_BIAS.n52 GND 4.95e-19
C74 DIFFPAIR_BIAS.n53 GND 9.22e-19
C75 DIFFPAIR_BIAS.n54 GND 9.22e-19
C76 DIFFPAIR_BIAS.n55 GND 4.95e-19
C77 DIFFPAIR_BIAS.n56 GND 5.25e-19
C78 DIFFPAIR_BIAS.n57 GND 0.001171f
C79 DIFFPAIR_BIAS.n58 GND 0.002535f
C80 DIFFPAIR_BIAS.n59 GND 5.25e-19
C81 DIFFPAIR_BIAS.n60 GND 4.95e-19
C82 DIFFPAIR_BIAS.n61 GND 0.002131f
C83 DIFFPAIR_BIAS.n62 GND 0.00491f
C84 DIFFPAIR_BIAS.n63 GND 0.11516f
C85 DIFFPAIR_BIAS.n64 GND 0.001296f
C86 DIFFPAIR_BIAS.n65 GND 9.22e-19
C87 DIFFPAIR_BIAS.n66 GND 4.95e-19
C88 DIFFPAIR_BIAS.n67 GND 0.001171f
C89 DIFFPAIR_BIAS.n68 GND 5.25e-19
C90 DIFFPAIR_BIAS.n69 GND 9.22e-19
C91 DIFFPAIR_BIAS.n70 GND 4.95e-19
C92 DIFFPAIR_BIAS.n71 GND 0.001171f
C93 DIFFPAIR_BIAS.n72 GND 5.25e-19
C94 DIFFPAIR_BIAS.n73 GND 0.003945f
C95 DIFFPAIR_BIAS.t5 GND 0.001909f
C96 DIFFPAIR_BIAS.n74 GND 8.78e-19
C97 DIFFPAIR_BIAS.n75 GND 6.92e-19
C98 DIFFPAIR_BIAS.n76 GND 4.95e-19
C99 DIFFPAIR_BIAS.n77 GND 0.021937f
C100 DIFFPAIR_BIAS.n78 GND 9.22e-19
C101 DIFFPAIR_BIAS.n79 GND 4.95e-19
C102 DIFFPAIR_BIAS.n80 GND 5.25e-19
C103 DIFFPAIR_BIAS.n81 GND 0.001171f
C104 DIFFPAIR_BIAS.n82 GND 0.001171f
C105 DIFFPAIR_BIAS.n83 GND 5.25e-19
C106 DIFFPAIR_BIAS.n84 GND 4.95e-19
C107 DIFFPAIR_BIAS.n85 GND 9.22e-19
C108 DIFFPAIR_BIAS.n86 GND 9.22e-19
C109 DIFFPAIR_BIAS.n87 GND 4.95e-19
C110 DIFFPAIR_BIAS.n88 GND 5.25e-19
C111 DIFFPAIR_BIAS.n89 GND 0.001171f
C112 DIFFPAIR_BIAS.n90 GND 0.002535f
C113 DIFFPAIR_BIAS.n91 GND 5.25e-19
C114 DIFFPAIR_BIAS.n92 GND 4.95e-19
C115 DIFFPAIR_BIAS.n93 GND 0.002131f
C116 DIFFPAIR_BIAS.n94 GND 0.00491f
C117 DIFFPAIR_BIAS.n95 GND 0.06095f
C118 DIFFPAIR_BIAS.n96 GND 0.001296f
C119 DIFFPAIR_BIAS.n97 GND 9.22e-19
C120 DIFFPAIR_BIAS.n98 GND 4.95e-19
C121 DIFFPAIR_BIAS.n99 GND 0.001171f
C122 DIFFPAIR_BIAS.n100 GND 5.25e-19
C123 DIFFPAIR_BIAS.n101 GND 9.22e-19
C124 DIFFPAIR_BIAS.n102 GND 4.95e-19
C125 DIFFPAIR_BIAS.n103 GND 0.001171f
C126 DIFFPAIR_BIAS.n104 GND 5.25e-19
C127 DIFFPAIR_BIAS.n105 GND 0.003945f
C128 DIFFPAIR_BIAS.t7 GND 0.001909f
C129 DIFFPAIR_BIAS.n106 GND 8.78e-19
C130 DIFFPAIR_BIAS.n107 GND 6.92e-19
C131 DIFFPAIR_BIAS.n108 GND 4.95e-19
C132 DIFFPAIR_BIAS.n109 GND 0.021937f
C133 DIFFPAIR_BIAS.n110 GND 9.22e-19
C134 DIFFPAIR_BIAS.n111 GND 4.95e-19
C135 DIFFPAIR_BIAS.n112 GND 5.25e-19
C136 DIFFPAIR_BIAS.n113 GND 0.001171f
C137 DIFFPAIR_BIAS.n114 GND 0.001171f
C138 DIFFPAIR_BIAS.n115 GND 5.25e-19
C139 DIFFPAIR_BIAS.n116 GND 4.95e-19
C140 DIFFPAIR_BIAS.n117 GND 9.22e-19
C141 DIFFPAIR_BIAS.n118 GND 9.22e-19
C142 DIFFPAIR_BIAS.n119 GND 4.95e-19
C143 DIFFPAIR_BIAS.n120 GND 5.25e-19
C144 DIFFPAIR_BIAS.n121 GND 0.001171f
C145 DIFFPAIR_BIAS.n122 GND 0.002535f
C146 DIFFPAIR_BIAS.n123 GND 5.25e-19
C147 DIFFPAIR_BIAS.n124 GND 4.95e-19
C148 DIFFPAIR_BIAS.n125 GND 0.002131f
C149 DIFFPAIR_BIAS.n126 GND 0.00491f
C150 DIFFPAIR_BIAS.n127 GND 0.08013f
C151 DIFFPAIR_BIAS.t6 GND 0.102337f
C152 DIFFPAIR_BIAS.t4 GND 0.102337f
C153 DIFFPAIR_BIAS.t2 GND 0.102337f
C154 DIFFPAIR_BIAS.t0 GND 0.103205f
C155 DIFFPAIR_BIAS.n128 GND 0.127236f
C156 DIFFPAIR_BIAS.n129 GND 0.068439f
C157 DIFFPAIR_BIAS.n130 GND 0.07541f
C158 DIFFPAIR_BIAS.n131 GND 0.155794f
C159 DIFFPAIR_BIAS.t11 GND 0.108432f
C160 DIFFPAIR_BIAS.n132 GND 0.063754f
C161 DIFFPAIR_BIAS.t10 GND 0.108432f
C162 DIFFPAIR_BIAS.n133 GND 0.061519f
C163 DIFFPAIR_BIAS.n134 GND 0.040079f
C164 VP.n0 GND 0.03666f
C165 VP.t6 GND 0.436296f
C166 VP.n1 GND 0.022189f
C167 VP.t11 GND 0.495129f
C168 VP.n2 GND 0.218457f
C169 VP.t10 GND 0.436296f
C170 VP.n3 GND 0.203585f
C171 VP.n4 GND 0.037464f
C172 VP.n5 GND 0.117613f
C173 VP.n6 GND 0.027473f
C174 VP.n7 GND 0.027473f
C175 VP.n8 GND 0.037464f
C176 VP.n9 GND 0.179138f
C177 VP.n10 GND 0.037684f
C178 VP.t5 GND 0.47813f
C179 VP.n11 GND 0.221639f
C180 VP.n12 GND 0.328479f
C181 VP.n13 GND 0.03666f
C182 VP.t7 GND 0.47813f
C183 VP.t12 GND 0.436296f
C184 VP.n14 GND 0.022189f
C185 VP.t9 GND 0.495129f
C186 VP.n15 GND 0.218457f
C187 VP.t8 GND 0.436296f
C188 VP.n16 GND 0.203585f
C189 VP.n17 GND 0.037464f
C190 VP.n18 GND 0.117613f
C191 VP.n19 GND 0.027473f
C192 VP.n20 GND 0.027473f
C193 VP.n21 GND 0.037464f
C194 VP.n22 GND 0.179138f
C195 VP.n23 GND 0.037684f
C196 VP.n24 GND 0.221639f
C197 VP.n25 GND 0.727079f
C198 VP.n26 GND 1.08549f
C199 VP.t4 GND 0.008469f
C200 VP.t1 GND 0.008469f
C201 VP.n27 GND 0.027849f
C202 VP.t0 GND 0.008469f
C203 VP.t2 GND 0.008469f
C204 VP.n28 GND 0.027467f
C205 VP.n29 GND 0.234421f
C206 VP.t3 GND 0.047139f
C207 VP.n30 GND 0.127921f
C208 VP.n31 GND 1.89655f
C209 a_n1455_n3628.n0 GND 0.029433f
C210 a_n1455_n3628.n1 GND 0.048734f
C211 a_n1455_n3628.n2 GND 0.029433f
C212 a_n1455_n3628.n3 GND 0.350169f
C213 a_n1455_n3628.n4 GND 0.029433f
C214 a_n1455_n3628.n5 GND 0.048734f
C215 a_n1455_n3628.n6 GND 0.029433f
C216 a_n1455_n3628.n7 GND 0.350169f
C217 a_n1455_n3628.n8 GND 0.029433f
C218 a_n1455_n3628.n9 GND 0.048734f
C219 a_n1455_n3628.n10 GND 0.029433f
C220 a_n1455_n3628.n11 GND 0.350169f
C221 a_n1455_n3628.n12 GND 0.029433f
C222 a_n1455_n3628.n13 GND 0.048734f
C223 a_n1455_n3628.n14 GND 0.029433f
C224 a_n1455_n3628.n15 GND 0.029433f
C225 a_n1455_n3628.n16 GND 0.029433f
C226 a_n1455_n3628.n17 GND 0.364885f
C227 a_n1455_n3628.n18 GND 0.029433f
C228 a_n1455_n3628.n19 GND 0.029433f
C229 a_n1455_n3628.n20 GND 0.364885f
C230 a_n1455_n3628.n21 GND 0.029433f
C231 a_n1455_n3628.n22 GND 0.029433f
C232 a_n1455_n3628.n23 GND 0.364885f
C233 a_n1455_n3628.n24 GND 0.029433f
C234 a_n1455_n3628.n25 GND 0.029433f
C235 a_n1455_n3628.n26 GND 0.364885f
C236 a_n1455_n3628.n27 GND 0.029433f
C237 a_n1455_n3628.n28 GND 0.029433f
C238 a_n1455_n3628.n29 GND 0.364885f
C239 a_n1455_n3628.n30 GND 0.029433f
C240 a_n1455_n3628.n31 GND 0.029433f
C241 a_n1455_n3628.n32 GND 0.364885f
C242 a_n1455_n3628.n33 GND 0.029433f
C243 a_n1455_n3628.n34 GND 0.029433f
C244 a_n1455_n3628.n35 GND 0.364885f
C245 a_n1455_n3628.n36 GND 0.029433f
C246 a_n1455_n3628.n37 GND 0.029433f
C247 a_n1455_n3628.n38 GND 0.364885f
C248 a_n1455_n3628.n39 GND 0.062977f
C249 a_n1455_n3628.n40 GND 0.018692f
C250 a_n1455_n3628.n41 GND 0.008373f
C251 a_n1455_n3628.n42 GND 0.007908f
C252 a_n1455_n3628.n43 GND 0.018692f
C253 a_n1455_n3628.n44 GND 0.008373f
C254 a_n1455_n3628.n45 GND 0.007908f
C255 a_n1455_n3628.n46 GND 0.020686f
C256 a_n1455_n3628.t4 GND 0.069777f
C257 a_n1455_n3628.t0 GND 0.069777f
C258 a_n1455_n3628.n47 GND 0.558309f
C259 a_n1455_n3628.n48 GND 0.347302f
C260 a_n1455_n3628.n49 GND 0.020686f
C261 a_n1455_n3628.n50 GND 0.007908f
C262 a_n1455_n3628.n51 GND 0.018692f
C263 a_n1455_n3628.n52 GND 0.008373f
C264 a_n1455_n3628.n53 GND 0.007908f
C265 a_n1455_n3628.n54 GND 0.018692f
C266 a_n1455_n3628.n55 GND 0.008373f
C267 a_n1455_n3628.n56 GND 0.062977f
C268 a_n1455_n3628.t2 GND 0.030465f
C269 a_n1455_n3628.n57 GND 0.014019f
C270 a_n1455_n3628.n58 GND 0.011041f
C271 a_n1455_n3628.n59 GND 0.007908f
C272 a_n1455_n3628.n60 GND 0.007908f
C273 a_n1455_n3628.n61 GND 0.008373f
C274 a_n1455_n3628.n62 GND 0.018692f
C275 a_n1455_n3628.n63 GND 0.018692f
C276 a_n1455_n3628.n64 GND 0.008373f
C277 a_n1455_n3628.n65 GND 0.007908f
C278 a_n1455_n3628.n66 GND 0.007908f
C279 a_n1455_n3628.n67 GND 0.008373f
C280 a_n1455_n3628.n68 GND 0.018692f
C281 a_n1455_n3628.n69 GND 0.040465f
C282 a_n1455_n3628.n70 GND 0.008373f
C283 a_n1455_n3628.n71 GND 0.007908f
C284 a_n1455_n3628.n72 GND 0.034017f
C285 a_n1455_n3628.n73 GND 0.026084f
C286 a_n1455_n3628.n74 GND 0.610154f
C287 a_n1455_n3628.t6 GND 0.069777f
C288 a_n1455_n3628.t1 GND 0.069777f
C289 a_n1455_n3628.n75 GND 0.558312f
C290 a_n1455_n3628.n76 GND 0.347298f
C291 a_n1455_n3628.n77 GND 0.020686f
C292 a_n1455_n3628.n78 GND 0.007908f
C293 a_n1455_n3628.n79 GND 0.018692f
C294 a_n1455_n3628.n80 GND 0.008373f
C295 a_n1455_n3628.n81 GND 0.007908f
C296 a_n1455_n3628.n82 GND 0.018692f
C297 a_n1455_n3628.n83 GND 0.008373f
C298 a_n1455_n3628.n84 GND 0.062977f
C299 a_n1455_n3628.t5 GND 0.030465f
C300 a_n1455_n3628.n85 GND 0.014019f
C301 a_n1455_n3628.n86 GND 0.011041f
C302 a_n1455_n3628.n87 GND 0.007908f
C303 a_n1455_n3628.n88 GND 0.007908f
C304 a_n1455_n3628.n89 GND 0.008373f
C305 a_n1455_n3628.n90 GND 0.018692f
C306 a_n1455_n3628.n91 GND 0.018692f
C307 a_n1455_n3628.n92 GND 0.008373f
C308 a_n1455_n3628.n93 GND 0.007908f
C309 a_n1455_n3628.n94 GND 0.007908f
C310 a_n1455_n3628.n95 GND 0.008373f
C311 a_n1455_n3628.n96 GND 0.018692f
C312 a_n1455_n3628.n97 GND 0.040465f
C313 a_n1455_n3628.n98 GND 0.008373f
C314 a_n1455_n3628.n99 GND 0.007908f
C315 a_n1455_n3628.n100 GND 0.034017f
C316 a_n1455_n3628.n101 GND 0.026084f
C317 a_n1455_n3628.n102 GND 0.16917f
C318 a_n1455_n3628.n103 GND 0.020686f
C319 a_n1455_n3628.n104 GND 0.007908f
C320 a_n1455_n3628.n105 GND 0.018692f
C321 a_n1455_n3628.n106 GND 0.008373f
C322 a_n1455_n3628.n107 GND 0.007908f
C323 a_n1455_n3628.n108 GND 0.018692f
C324 a_n1455_n3628.n109 GND 0.008373f
C325 a_n1455_n3628.n110 GND 0.062977f
C326 a_n1455_n3628.t18 GND 0.030465f
C327 a_n1455_n3628.n111 GND 0.014019f
C328 a_n1455_n3628.n112 GND 0.011041f
C329 a_n1455_n3628.n113 GND 0.007908f
C330 a_n1455_n3628.n114 GND 0.007908f
C331 a_n1455_n3628.n115 GND 0.008373f
C332 a_n1455_n3628.n116 GND 0.018692f
C333 a_n1455_n3628.n117 GND 0.018692f
C334 a_n1455_n3628.n118 GND 0.008373f
C335 a_n1455_n3628.n119 GND 0.007908f
C336 a_n1455_n3628.n120 GND 0.007908f
C337 a_n1455_n3628.n121 GND 0.008373f
C338 a_n1455_n3628.n122 GND 0.018692f
C339 a_n1455_n3628.n123 GND 0.040465f
C340 a_n1455_n3628.n124 GND 0.008373f
C341 a_n1455_n3628.n125 GND 0.007908f
C342 a_n1455_n3628.n126 GND 0.034017f
C343 a_n1455_n3628.n127 GND 0.026084f
C344 a_n1455_n3628.n128 GND 0.16917f
C345 a_n1455_n3628.t8 GND 0.069777f
C346 a_n1455_n3628.t19 GND 0.069777f
C347 a_n1455_n3628.n129 GND 0.558312f
C348 a_n1455_n3628.n130 GND 0.347298f
C349 a_n1455_n3628.n131 GND 0.020686f
C350 a_n1455_n3628.n132 GND 0.007908f
C351 a_n1455_n3628.n133 GND 0.018692f
C352 a_n1455_n3628.n134 GND 0.008373f
C353 a_n1455_n3628.n135 GND 0.007908f
C354 a_n1455_n3628.n136 GND 0.018692f
C355 a_n1455_n3628.n137 GND 0.008373f
C356 a_n1455_n3628.n138 GND 0.062977f
C357 a_n1455_n3628.t15 GND 0.030465f
C358 a_n1455_n3628.n139 GND 0.014019f
C359 a_n1455_n3628.n140 GND 0.011041f
C360 a_n1455_n3628.n141 GND 0.007908f
C361 a_n1455_n3628.n142 GND 0.007908f
C362 a_n1455_n3628.n143 GND 0.008373f
C363 a_n1455_n3628.n144 GND 0.018692f
C364 a_n1455_n3628.n145 GND 0.018692f
C365 a_n1455_n3628.n146 GND 0.008373f
C366 a_n1455_n3628.n147 GND 0.007908f
C367 a_n1455_n3628.n148 GND 0.007908f
C368 a_n1455_n3628.n149 GND 0.008373f
C369 a_n1455_n3628.n150 GND 0.018692f
C370 a_n1455_n3628.n151 GND 0.040465f
C371 a_n1455_n3628.n152 GND 0.008373f
C372 a_n1455_n3628.n153 GND 0.007908f
C373 a_n1455_n3628.n154 GND 0.034017f
C374 a_n1455_n3628.n155 GND 0.026084f
C375 a_n1455_n3628.n156 GND 0.610154f
C376 a_n1455_n3628.n157 GND 0.020686f
C377 a_n1455_n3628.n158 GND 0.007908f
C378 a_n1455_n3628.n159 GND 0.018692f
C379 a_n1455_n3628.n160 GND 0.008373f
C380 a_n1455_n3628.n161 GND 0.007908f
C381 a_n1455_n3628.n162 GND 0.018692f
C382 a_n1455_n3628.n163 GND 0.008373f
C383 a_n1455_n3628.n164 GND 0.062977f
C384 a_n1455_n3628.t3 GND 0.030465f
C385 a_n1455_n3628.n165 GND 0.014019f
C386 a_n1455_n3628.n166 GND 0.011041f
C387 a_n1455_n3628.n167 GND 0.007908f
C388 a_n1455_n3628.n168 GND 0.007908f
C389 a_n1455_n3628.n169 GND 0.008373f
C390 a_n1455_n3628.n170 GND 0.018692f
C391 a_n1455_n3628.n171 GND 0.018692f
C392 a_n1455_n3628.n172 GND 0.008373f
C393 a_n1455_n3628.n173 GND 0.007908f
C394 a_n1455_n3628.n174 GND 0.007908f
C395 a_n1455_n3628.n175 GND 0.008373f
C396 a_n1455_n3628.n176 GND 0.018692f
C397 a_n1455_n3628.n177 GND 0.040465f
C398 a_n1455_n3628.n178 GND 0.008373f
C399 a_n1455_n3628.n179 GND 0.007908f
C400 a_n1455_n3628.n180 GND 0.026084f
C401 a_n1455_n3628.n181 GND 0.381969f
C402 a_n1455_n3628.n182 GND 0.714807f
C403 a_n1455_n3628.n183 GND 0.020686f
C404 a_n1455_n3628.n184 GND 0.007908f
C405 a_n1455_n3628.n185 GND 0.018692f
C406 a_n1455_n3628.n186 GND 0.008373f
C407 a_n1455_n3628.n187 GND 0.007908f
C408 a_n1455_n3628.n188 GND 0.018692f
C409 a_n1455_n3628.n189 GND 0.008373f
C410 a_n1455_n3628.n190 GND 0.062977f
C411 a_n1455_n3628.t11 GND 0.030465f
C412 a_n1455_n3628.n191 GND 0.014019f
C413 a_n1455_n3628.n192 GND 0.011041f
C414 a_n1455_n3628.n193 GND 0.007908f
C415 a_n1455_n3628.n194 GND 0.007908f
C416 a_n1455_n3628.n195 GND 0.008373f
C417 a_n1455_n3628.n196 GND 0.018692f
C418 a_n1455_n3628.n197 GND 0.018692f
C419 a_n1455_n3628.n198 GND 0.008373f
C420 a_n1455_n3628.n199 GND 0.007908f
C421 a_n1455_n3628.n200 GND 0.007908f
C422 a_n1455_n3628.n201 GND 0.008373f
C423 a_n1455_n3628.n202 GND 0.018692f
C424 a_n1455_n3628.n203 GND 0.040465f
C425 a_n1455_n3628.n204 GND 0.008373f
C426 a_n1455_n3628.n205 GND 0.007908f
C427 a_n1455_n3628.n206 GND 0.034017f
C428 a_n1455_n3628.n207 GND 0.122845f
C429 a_n1455_n3628.n208 GND 0.89644f
C430 a_n1455_n3628.n209 GND 0.020686f
C431 a_n1455_n3628.n210 GND 0.007908f
C432 a_n1455_n3628.n211 GND 0.018692f
C433 a_n1455_n3628.n212 GND 0.008373f
C434 a_n1455_n3628.n213 GND 0.007908f
C435 a_n1455_n3628.n214 GND 0.018692f
C436 a_n1455_n3628.n215 GND 0.008373f
C437 a_n1455_n3628.n216 GND 0.062977f
C438 a_n1455_n3628.t12 GND 0.030465f
C439 a_n1455_n3628.n217 GND 0.014019f
C440 a_n1455_n3628.n218 GND 0.011041f
C441 a_n1455_n3628.n219 GND 0.007908f
C442 a_n1455_n3628.n220 GND 0.007908f
C443 a_n1455_n3628.n221 GND 0.008373f
C444 a_n1455_n3628.n222 GND 0.018692f
C445 a_n1455_n3628.n223 GND 0.018692f
C446 a_n1455_n3628.n224 GND 0.008373f
C447 a_n1455_n3628.n225 GND 0.007908f
C448 a_n1455_n3628.n226 GND 0.007908f
C449 a_n1455_n3628.n227 GND 0.008373f
C450 a_n1455_n3628.n228 GND 0.018692f
C451 a_n1455_n3628.n229 GND 0.040465f
C452 a_n1455_n3628.n230 GND 0.008373f
C453 a_n1455_n3628.n231 GND 0.007908f
C454 a_n1455_n3628.n232 GND 0.034017f
C455 a_n1455_n3628.n233 GND 0.121814f
C456 a_n1455_n3628.n234 GND 0.708238f
C457 a_n1455_n3628.n235 GND 0.020686f
C458 a_n1455_n3628.n236 GND 0.007908f
C459 a_n1455_n3628.n237 GND 0.018692f
C460 a_n1455_n3628.n238 GND 0.008373f
C461 a_n1455_n3628.n239 GND 0.007908f
C462 a_n1455_n3628.n240 GND 0.018692f
C463 a_n1455_n3628.n241 GND 0.008373f
C464 a_n1455_n3628.n242 GND 0.062977f
C465 a_n1455_n3628.t14 GND 0.030465f
C466 a_n1455_n3628.n243 GND 0.014019f
C467 a_n1455_n3628.n244 GND 0.011041f
C468 a_n1455_n3628.n245 GND 0.007908f
C469 a_n1455_n3628.n246 GND 0.007908f
C470 a_n1455_n3628.n247 GND 0.008373f
C471 a_n1455_n3628.n248 GND 0.018692f
C472 a_n1455_n3628.n249 GND 0.018692f
C473 a_n1455_n3628.n250 GND 0.008373f
C474 a_n1455_n3628.n251 GND 0.007908f
C475 a_n1455_n3628.n252 GND 0.007908f
C476 a_n1455_n3628.n253 GND 0.008373f
C477 a_n1455_n3628.n254 GND 0.018692f
C478 a_n1455_n3628.n255 GND 0.040465f
C479 a_n1455_n3628.n256 GND 0.008373f
C480 a_n1455_n3628.n257 GND 0.007908f
C481 a_n1455_n3628.n258 GND 0.034017f
C482 a_n1455_n3628.n259 GND 0.121814f
C483 a_n1455_n3628.n260 GND 0.933421f
C484 a_n1455_n3628.n261 GND 0.020686f
C485 a_n1455_n3628.n262 GND 0.007908f
C486 a_n1455_n3628.n263 GND 0.018692f
C487 a_n1455_n3628.n264 GND 0.008373f
C488 a_n1455_n3628.n265 GND 0.007908f
C489 a_n1455_n3628.n266 GND 0.018692f
C490 a_n1455_n3628.n267 GND 0.008373f
C491 a_n1455_n3628.n268 GND 0.062977f
C492 a_n1455_n3628.t13 GND 0.030465f
C493 a_n1455_n3628.n269 GND 0.014019f
C494 a_n1455_n3628.n270 GND 0.011041f
C495 a_n1455_n3628.n271 GND 0.007908f
C496 a_n1455_n3628.n272 GND 0.007908f
C497 a_n1455_n3628.n273 GND 0.008373f
C498 a_n1455_n3628.n274 GND 0.018692f
C499 a_n1455_n3628.n275 GND 0.018692f
C500 a_n1455_n3628.n276 GND 0.008373f
C501 a_n1455_n3628.n277 GND 0.007908f
C502 a_n1455_n3628.n278 GND 0.007908f
C503 a_n1455_n3628.n279 GND 0.008373f
C504 a_n1455_n3628.n280 GND 0.018692f
C505 a_n1455_n3628.n281 GND 0.040465f
C506 a_n1455_n3628.n282 GND 0.008373f
C507 a_n1455_n3628.n283 GND 0.007908f
C508 a_n1455_n3628.n284 GND 0.034017f
C509 a_n1455_n3628.n285 GND 0.121814f
C510 a_n1455_n3628.n286 GND 1.26754f
C511 a_n1455_n3628.n287 GND 0.80329f
C512 a_n1455_n3628.n288 GND 0.020686f
C513 a_n1455_n3628.n289 GND 0.007908f
C514 a_n1455_n3628.n290 GND 0.018692f
C515 a_n1455_n3628.n291 GND 0.008373f
C516 a_n1455_n3628.n292 GND 0.007908f
C517 a_n1455_n3628.n293 GND 0.018692f
C518 a_n1455_n3628.n294 GND 0.008373f
C519 a_n1455_n3628.n295 GND 0.062977f
C520 a_n1455_n3628.t17 GND 0.030465f
C521 a_n1455_n3628.n296 GND 0.014019f
C522 a_n1455_n3628.n297 GND 0.011041f
C523 a_n1455_n3628.n298 GND 0.007908f
C524 a_n1455_n3628.n299 GND 0.007908f
C525 a_n1455_n3628.n300 GND 0.008373f
C526 a_n1455_n3628.n301 GND 0.018692f
C527 a_n1455_n3628.n302 GND 0.018692f
C528 a_n1455_n3628.n303 GND 0.008373f
C529 a_n1455_n3628.n304 GND 0.007908f
C530 a_n1455_n3628.n305 GND 0.007908f
C531 a_n1455_n3628.n306 GND 0.008373f
C532 a_n1455_n3628.n307 GND 0.018692f
C533 a_n1455_n3628.n308 GND 0.040465f
C534 a_n1455_n3628.n309 GND 0.008373f
C535 a_n1455_n3628.n310 GND 0.007908f
C536 a_n1455_n3628.n311 GND 0.026084f
C537 a_n1455_n3628.n312 GND 0.381969f
C538 a_n1455_n3628.t16 GND 0.069777f
C539 a_n1455_n3628.t10 GND 0.069777f
C540 a_n1455_n3628.n313 GND 0.558309f
C541 a_n1455_n3628.n314 GND 0.347302f
C542 a_n1455_n3628.n315 GND 0.020686f
C543 a_n1455_n3628.n316 GND 0.007908f
C544 a_n1455_n3628.n317 GND 0.018692f
C545 a_n1455_n3628.n318 GND 0.008373f
C546 a_n1455_n3628.n319 GND 0.007908f
C547 a_n1455_n3628.n320 GND 0.018692f
C548 a_n1455_n3628.n321 GND 0.008373f
C549 a_n1455_n3628.n322 GND 0.062977f
C550 a_n1455_n3628.t9 GND 0.030465f
C551 a_n1455_n3628.n323 GND 0.014019f
C552 a_n1455_n3628.n324 GND 0.011041f
C553 a_n1455_n3628.n325 GND 0.007908f
C554 a_n1455_n3628.n326 GND 0.007908f
C555 a_n1455_n3628.n327 GND 0.008373f
C556 a_n1455_n3628.n328 GND 0.018692f
C557 a_n1455_n3628.n329 GND 0.018692f
C558 a_n1455_n3628.n330 GND 0.008373f
C559 a_n1455_n3628.n331 GND 0.007908f
C560 a_n1455_n3628.n332 GND 0.007908f
C561 a_n1455_n3628.n333 GND 0.008373f
C562 a_n1455_n3628.n334 GND 0.018692f
C563 a_n1455_n3628.n335 GND 0.040465f
C564 a_n1455_n3628.n336 GND 0.008373f
C565 a_n1455_n3628.n337 GND 0.007908f
C566 a_n1455_n3628.n338 GND 0.026084f
C567 a_n1455_n3628.n339 GND 0.16917f
C568 a_n1455_n3628.n340 GND 0.16917f
C569 a_n1455_n3628.n341 GND 0.026084f
C570 a_n1455_n3628.n342 GND 0.007908f
C571 a_n1455_n3628.n343 GND 0.008373f
C572 a_n1455_n3628.n344 GND 0.040465f
C573 a_n1455_n3628.n345 GND 0.018692f
C574 a_n1455_n3628.n346 GND 0.008373f
C575 a_n1455_n3628.n347 GND 0.007908f
C576 a_n1455_n3628.n348 GND 0.007908f
C577 a_n1455_n3628.n349 GND 0.008373f
C578 a_n1455_n3628.n350 GND 0.018692f
C579 a_n1455_n3628.n351 GND 0.018692f
C580 a_n1455_n3628.n352 GND 0.008373f
C581 a_n1455_n3628.n353 GND 0.007908f
C582 a_n1455_n3628.n354 GND 0.350169f
C583 a_n1455_n3628.n355 GND 0.007908f
C584 a_n1455_n3628.n356 GND 0.011041f
C585 a_n1455_n3628.n357 GND 0.014019f
C586 a_n1455_n3628.t7 GND 0.030465f
C587 VN.n0 GND 0.025584f
C588 VN.t9 GND 0.33368f
C589 VN.t8 GND 0.304485f
C590 VN.n1 GND 0.015486f
C591 VN.t5 GND 0.345544f
C592 VN.n2 GND 0.152458f
C593 VN.t12 GND 0.304485f
C594 VN.n3 GND 0.14208f
C595 VN.n4 GND 0.026146f
C596 VN.n5 GND 0.082081f
C597 VN.n6 GND 0.019173f
C598 VN.n7 GND 0.019173f
C599 VN.n8 GND 0.026146f
C600 VN.n9 GND 0.125018f
C601 VN.n10 GND 0.026299f
C602 VN.n11 GND 0.154679f
C603 VN.n12 GND 0.224439f
C604 VN.n13 GND 0.025584f
C605 VN.t11 GND 0.304485f
C606 VN.n14 GND 0.015486f
C607 VN.t7 GND 0.345544f
C608 VN.n15 GND 0.152458f
C609 VN.t6 GND 0.304485f
C610 VN.n16 GND 0.14208f
C611 VN.n17 GND 0.026146f
C612 VN.n18 GND 0.08208f
C613 VN.n19 GND 0.019173f
C614 VN.n20 GND 0.019173f
C615 VN.n21 GND 0.026146f
C616 VN.n22 GND 0.125018f
C617 VN.n23 GND 0.026299f
C618 VN.t10 GND 0.33368f
C619 VN.n24 GND 0.154679f
C620 VN.n25 GND 0.499734f
C621 VN.n26 GND 0.749818f
C622 VN.t0 GND 0.033099f
C623 VN.t1 GND 0.005911f
C624 VN.t4 GND 0.005911f
C625 VN.n27 GND 0.019169f
C626 VN.n28 GND 0.148811f
C627 VN.t2 GND 0.005911f
C628 VN.t3 GND 0.005911f
C629 VN.n29 GND 0.019169f
C630 VN.n30 GND 0.111701f
C631 VN.n31 GND 1.99192f
C632 a_n2511_10356.t17 GND 0.115432f
C633 a_n2511_10356.t16 GND 0.115432f
C634 a_n2511_10356.n0 GND 0.832956f
C635 a_n2511_10356.t11 GND 0.115432f
C636 a_n2511_10356.t13 GND 0.115432f
C637 a_n2511_10356.n1 GND 0.83019f
C638 a_n2511_10356.n2 GND 2.53408f
C639 a_n2511_10356.t15 GND 0.115432f
C640 a_n2511_10356.t19 GND 0.115432f
C641 a_n2511_10356.n3 GND 0.83019f
C642 a_n2511_10356.n4 GND 3.97422f
C643 a_n2511_10356.n5 GND 0.026649f
C644 a_n2511_10356.n6 GND 0.024346f
C645 a_n2511_10356.n7 GND 0.013082f
C646 a_n2511_10356.n8 GND 0.030922f
C647 a_n2511_10356.n9 GND 0.013852f
C648 a_n2511_10356.n10 GND 0.024346f
C649 a_n2511_10356.n11 GND 0.013082f
C650 a_n2511_10356.n12 GND 0.030922f
C651 a_n2511_10356.n13 GND 0.013852f
C652 a_n2511_10356.n14 GND 0.107644f
C653 a_n2511_10356.t0 GND 0.06635f
C654 a_n2511_10356.n15 GND 0.023191f
C655 a_n2511_10356.n16 GND 0.019661f
C656 a_n2511_10356.n17 GND 0.013082f
C657 a_n2511_10356.n18 GND 0.558473f
C658 a_n2511_10356.n19 GND 0.024346f
C659 a_n2511_10356.n20 GND 0.013082f
C660 a_n2511_10356.n21 GND 0.013852f
C661 a_n2511_10356.n22 GND 0.030922f
C662 a_n2511_10356.n23 GND 0.030922f
C663 a_n2511_10356.n24 GND 0.013852f
C664 a_n2511_10356.n25 GND 0.013082f
C665 a_n2511_10356.n26 GND 0.024346f
C666 a_n2511_10356.n27 GND 0.024346f
C667 a_n2511_10356.n28 GND 0.013082f
C668 a_n2511_10356.n29 GND 0.013852f
C669 a_n2511_10356.n30 GND 0.030922f
C670 a_n2511_10356.n31 GND 0.074512f
C671 a_n2511_10356.n32 GND 0.013852f
C672 a_n2511_10356.n33 GND 0.013082f
C673 a_n2511_10356.n34 GND 0.056274f
C674 a_n2511_10356.n35 GND 0.046522f
C675 a_n2511_10356.t5 GND 0.115432f
C676 a_n2511_10356.t7 GND 0.115432f
C677 a_n2511_10356.n36 GND 0.71063f
C678 a_n2511_10356.n37 GND 1.0099f
C679 a_n2511_10356.n38 GND 0.026649f
C680 a_n2511_10356.n39 GND 0.024346f
C681 a_n2511_10356.n40 GND 0.013082f
C682 a_n2511_10356.n41 GND 0.030922f
C683 a_n2511_10356.n42 GND 0.013852f
C684 a_n2511_10356.n43 GND 0.024346f
C685 a_n2511_10356.n44 GND 0.013082f
C686 a_n2511_10356.n45 GND 0.030922f
C687 a_n2511_10356.n46 GND 0.013852f
C688 a_n2511_10356.n47 GND 0.107644f
C689 a_n2511_10356.t3 GND 0.06635f
C690 a_n2511_10356.n48 GND 0.023191f
C691 a_n2511_10356.n49 GND 0.019661f
C692 a_n2511_10356.n50 GND 0.013082f
C693 a_n2511_10356.n51 GND 0.558473f
C694 a_n2511_10356.n52 GND 0.024346f
C695 a_n2511_10356.n53 GND 0.013082f
C696 a_n2511_10356.n54 GND 0.013852f
C697 a_n2511_10356.n55 GND 0.030922f
C698 a_n2511_10356.n56 GND 0.030922f
C699 a_n2511_10356.n57 GND 0.013852f
C700 a_n2511_10356.n58 GND 0.013082f
C701 a_n2511_10356.n59 GND 0.024346f
C702 a_n2511_10356.n60 GND 0.024346f
C703 a_n2511_10356.n61 GND 0.013082f
C704 a_n2511_10356.n62 GND 0.013852f
C705 a_n2511_10356.n63 GND 0.030922f
C706 a_n2511_10356.n64 GND 0.074512f
C707 a_n2511_10356.n65 GND 0.013852f
C708 a_n2511_10356.n66 GND 0.013082f
C709 a_n2511_10356.n67 GND 0.056274f
C710 a_n2511_10356.n68 GND 0.043151f
C711 a_n2511_10356.n69 GND 0.254836f
C712 a_n2511_10356.n70 GND 0.026649f
C713 a_n2511_10356.n71 GND 0.024346f
C714 a_n2511_10356.n72 GND 0.013082f
C715 a_n2511_10356.n73 GND 0.030922f
C716 a_n2511_10356.n74 GND 0.013852f
C717 a_n2511_10356.n75 GND 0.024346f
C718 a_n2511_10356.n76 GND 0.013082f
C719 a_n2511_10356.n77 GND 0.030922f
C720 a_n2511_10356.n78 GND 0.013852f
C721 a_n2511_10356.n79 GND 0.107644f
C722 a_n2511_10356.t6 GND 0.06635f
C723 a_n2511_10356.n80 GND 0.023191f
C724 a_n2511_10356.n81 GND 0.019661f
C725 a_n2511_10356.n82 GND 0.013082f
C726 a_n2511_10356.n83 GND 0.558473f
C727 a_n2511_10356.n84 GND 0.024346f
C728 a_n2511_10356.n85 GND 0.013082f
C729 a_n2511_10356.n86 GND 0.013852f
C730 a_n2511_10356.n87 GND 0.030922f
C731 a_n2511_10356.n88 GND 0.030922f
C732 a_n2511_10356.n89 GND 0.013852f
C733 a_n2511_10356.n90 GND 0.013082f
C734 a_n2511_10356.n91 GND 0.024346f
C735 a_n2511_10356.n92 GND 0.024346f
C736 a_n2511_10356.n93 GND 0.013082f
C737 a_n2511_10356.n94 GND 0.013852f
C738 a_n2511_10356.n95 GND 0.030922f
C739 a_n2511_10356.n96 GND 0.074512f
C740 a_n2511_10356.n97 GND 0.013852f
C741 a_n2511_10356.n98 GND 0.013082f
C742 a_n2511_10356.n99 GND 0.056274f
C743 a_n2511_10356.n100 GND 0.043151f
C744 a_n2511_10356.n101 GND 0.254836f
C745 a_n2511_10356.t2 GND 0.115432f
C746 a_n2511_10356.t4 GND 0.115432f
C747 a_n2511_10356.n102 GND 0.71063f
C748 a_n2511_10356.n103 GND 0.787516f
C749 a_n2511_10356.n104 GND 0.026649f
C750 a_n2511_10356.n105 GND 0.024346f
C751 a_n2511_10356.n106 GND 0.013082f
C752 a_n2511_10356.n107 GND 0.030922f
C753 a_n2511_10356.n108 GND 0.013852f
C754 a_n2511_10356.n109 GND 0.024346f
C755 a_n2511_10356.n110 GND 0.013082f
C756 a_n2511_10356.n111 GND 0.030922f
C757 a_n2511_10356.n112 GND 0.013852f
C758 a_n2511_10356.n113 GND 0.107644f
C759 a_n2511_10356.t1 GND 0.06635f
C760 a_n2511_10356.n114 GND 0.023191f
C761 a_n2511_10356.n115 GND 0.019661f
C762 a_n2511_10356.n116 GND 0.013082f
C763 a_n2511_10356.n117 GND 0.558473f
C764 a_n2511_10356.n118 GND 0.024346f
C765 a_n2511_10356.n119 GND 0.013082f
C766 a_n2511_10356.n120 GND 0.013852f
C767 a_n2511_10356.n121 GND 0.030922f
C768 a_n2511_10356.n122 GND 0.030922f
C769 a_n2511_10356.n123 GND 0.013852f
C770 a_n2511_10356.n124 GND 0.013082f
C771 a_n2511_10356.n125 GND 0.024346f
C772 a_n2511_10356.n126 GND 0.024346f
C773 a_n2511_10356.n127 GND 0.013082f
C774 a_n2511_10356.n128 GND 0.013852f
C775 a_n2511_10356.n129 GND 0.030922f
C776 a_n2511_10356.n130 GND 0.074512f
C777 a_n2511_10356.n131 GND 0.013852f
C778 a_n2511_10356.n132 GND 0.013082f
C779 a_n2511_10356.n133 GND 0.056274f
C780 a_n2511_10356.n134 GND 0.043151f
C781 a_n2511_10356.n135 GND 1.01107f
C782 a_n2511_10356.n136 GND 2.19802f
C783 a_n2511_10356.t12 GND 0.115432f
C784 a_n2511_10356.t14 GND 0.115432f
C785 a_n2511_10356.n137 GND 0.830187f
C786 a_n2511_10356.n138 GND 1.64602f
C787 a_n2511_10356.t10 GND 0.115432f
C788 a_n2511_10356.t8 GND 0.115432f
C789 a_n2511_10356.n139 GND 0.83019f
C790 a_n2511_10356.n140 GND 1.46246f
C791 a_n2511_10356.t9 GND 0.115432f
C792 a_n2511_10356.n141 GND 0.834071f
C793 a_n2511_10356.t18 GND 0.115432f
C794 a_n2686_12578.n0 GND 0.758904f
C795 a_n2686_12578.n1 GND 0.352654f
C796 a_n2686_12578.n2 GND 0.755916f
C797 a_n2686_12578.n3 GND 0.620312f
C798 a_n2686_12578.n4 GND 0.352654f
C799 a_n2686_12578.n5 GND 0.678686f
C800 a_n2686_12578.n6 GND 0.352654f
C801 a_n2686_12578.n7 GND 0.723147f
C802 a_n2686_12578.n8 GND 0.352654f
C803 a_n2686_12578.n9 GND 0.632638f
C804 a_n2686_12578.n10 GND 0.352654f
C805 a_n2686_12578.n11 GND 0.552207f
C806 a_n2686_12578.n12 GND 0.352654f
C807 a_n2686_12578.n13 GND 0.054021f
C808 a_n2686_12578.n14 GND 0.054021f
C809 a_n2686_12578.n15 GND 0.054021f
C810 a_n2686_12578.n16 GND 0.045249f
C811 a_n2686_12578.n17 GND 0.054021f
C812 a_n2686_12578.n18 GND 0.045249f
C813 a_n2686_12578.n19 GND 0.054021f
C814 a_n2686_12578.n20 GND 0.045249f
C815 a_n2686_12578.n21 GND 0.054021f
C816 a_n2686_12578.n22 GND 0.074231f
C817 a_n2686_12578.n23 GND 0.045249f
C818 a_n2686_12578.n24 GND 0.061445f
C819 a_n2686_12578.n25 GND 0.092095f
C820 a_n2686_12578.n26 GND 0.107492f
C821 a_n2686_12578.n27 GND 0.074231f
C822 a_n2686_12578.n28 GND 0.045249f
C823 a_n2686_12578.n29 GND 0.061445f
C824 a_n2686_12578.n30 GND 0.092095f
C825 a_n2686_12578.n31 GND 0.107492f
C826 a_n2686_12578.n32 GND 0.074231f
C827 a_n2686_12578.n33 GND 0.045249f
C828 a_n2686_12578.n34 GND 0.061445f
C829 a_n2686_12578.n35 GND 0.092095f
C830 a_n2686_12578.n36 GND 0.107492f
C831 a_n2686_12578.n37 GND 0.074231f
C832 a_n2686_12578.n38 GND 0.045249f
C833 a_n2686_12578.n39 GND 0.061445f
C834 a_n2686_12578.n40 GND 0.092095f
C835 a_n2686_12578.n41 GND 0.107492f
C836 a_n2686_12578.n42 GND 0.092095f
C837 a_n2686_12578.n43 GND 0.061445f
C838 a_n2686_12578.n44 GND 0.092095f
C839 a_n2686_12578.n45 GND 0.092095f
C840 a_n2686_12578.n46 GND 0.092095f
C841 a_n2686_12578.n47 GND 0.045249f
C842 a_n2686_12578.n48 GND 0.107492f
C843 a_n2686_12578.n49 GND 0.054021f
C844 a_n2686_12578.n50 GND 0.123121f
C845 a_n2686_12578.n51 GND 0.041966f
C846 a_n2686_12578.n52 GND 0.035927f
C847 a_n2686_12578.n53 GND 0.035927f
C848 a_n2686_12578.n54 GND 0.430029f
C849 a_n2686_12578.n55 GND 0.035927f
C850 a_n2686_12578.n56 GND 0.035927f
C851 a_n2686_12578.n57 GND 0.430029f
C852 a_n2686_12578.n58 GND 0.035927f
C853 a_n2686_12578.n59 GND 0.035927f
C854 a_n2686_12578.n60 GND 0.430029f
C855 a_n2686_12578.n61 GND 0.035927f
C856 a_n2686_12578.n62 GND 0.035927f
C857 a_n2686_12578.n63 GND 0.430029f
C858 a_n2686_12578.t27 GND 0.085171f
C859 a_n2686_12578.t25 GND 0.085171f
C860 a_n2686_12578.t28 GND 0.085171f
C861 a_n2686_12578.n64 GND 0.745023f
C862 a_n2686_12578.t26 GND 0.085171f
C863 a_n2686_12578.t29 GND 0.085171f
C864 a_n2686_12578.n65 GND 0.745023f
C865 a_n2686_12578.n66 GND 2.15627f
C866 a_n2686_12578.t50 GND 0.842114f
C867 a_n2686_12578.t59 GND 0.731265f
C868 a_n2686_12578.n67 GND 0.398404f
C869 a_n2686_12578.t56 GND 0.731265f
C870 a_n2686_12578.t47 GND 0.731265f
C871 a_n2686_12578.t54 GND 0.731265f
C872 a_n2686_12578.n68 GND 0.398404f
C873 a_n2686_12578.t53 GND 0.842114f
C874 a_n2686_12578.n69 GND 0.019663f
C875 a_n2686_12578.n70 GND 0.009653f
C876 a_n2686_12578.n71 GND 0.022816f
C877 a_n2686_12578.n72 GND 0.01022f
C878 a_n2686_12578.n73 GND 0.009653f
C879 a_n2686_12578.n74 GND 0.022816f
C880 a_n2686_12578.n75 GND 0.01022f
C881 a_n2686_12578.n76 GND 0.079425f
C882 a_n2686_12578.t6 GND 0.048956f
C883 a_n2686_12578.n77 GND 0.017112f
C884 a_n2686_12578.n78 GND 0.014506f
C885 a_n2686_12578.n79 GND 0.009653f
C886 a_n2686_12578.n80 GND 0.009653f
C887 a_n2686_12578.n81 GND 0.01022f
C888 a_n2686_12578.n82 GND 0.022816f
C889 a_n2686_12578.n83 GND 0.022816f
C890 a_n2686_12578.n84 GND 0.01022f
C891 a_n2686_12578.n85 GND 0.009653f
C892 a_n2686_12578.n86 GND 0.009653f
C893 a_n2686_12578.n87 GND 0.01022f
C894 a_n2686_12578.n88 GND 0.022816f
C895 a_n2686_12578.n89 GND 0.054978f
C896 a_n2686_12578.n90 GND 0.01022f
C897 a_n2686_12578.n91 GND 0.009653f
C898 a_n2686_12578.n92 GND 0.041521f
C899 a_n2686_12578.n93 GND 0.034326f
C900 a_n2686_12578.t8 GND 0.085171f
C901 a_n2686_12578.t12 GND 0.085171f
C902 a_n2686_12578.n94 GND 0.524334f
C903 a_n2686_12578.n95 GND 0.745148f
C904 a_n2686_12578.t4 GND 0.085171f
C905 a_n2686_12578.t14 GND 0.085171f
C906 a_n2686_12578.n96 GND 0.524334f
C907 a_n2686_12578.n97 GND 0.581063f
C908 a_n2686_12578.n98 GND 0.019663f
C909 a_n2686_12578.n99 GND 0.009653f
C910 a_n2686_12578.n100 GND 0.022816f
C911 a_n2686_12578.n101 GND 0.01022f
C912 a_n2686_12578.n102 GND 0.009653f
C913 a_n2686_12578.n103 GND 0.022816f
C914 a_n2686_12578.n104 GND 0.01022f
C915 a_n2686_12578.n105 GND 0.079425f
C916 a_n2686_12578.t24 GND 0.048956f
C917 a_n2686_12578.n106 GND 0.017112f
C918 a_n2686_12578.n107 GND 0.014506f
C919 a_n2686_12578.n108 GND 0.009653f
C920 a_n2686_12578.n109 GND 0.009653f
C921 a_n2686_12578.n110 GND 0.01022f
C922 a_n2686_12578.n111 GND 0.022816f
C923 a_n2686_12578.n112 GND 0.022816f
C924 a_n2686_12578.n113 GND 0.01022f
C925 a_n2686_12578.n114 GND 0.009653f
C926 a_n2686_12578.n115 GND 0.009653f
C927 a_n2686_12578.n116 GND 0.01022f
C928 a_n2686_12578.n117 GND 0.022816f
C929 a_n2686_12578.n118 GND 0.054978f
C930 a_n2686_12578.n119 GND 0.01022f
C931 a_n2686_12578.n120 GND 0.009653f
C932 a_n2686_12578.n121 GND 0.041521f
C933 a_n2686_12578.n122 GND 0.031838f
C934 a_n2686_12578.n123 GND 0.693228f
C935 a_n2686_12578.t41 GND 0.731265f
C936 a_n2686_12578.t51 GND 0.731265f
C937 a_n2686_12578.t38 GND 0.80138f
C938 a_n2686_12578.t37 GND 0.731265f
C939 a_n2686_12578.t40 GND 0.731265f
C940 a_n2686_12578.t58 GND 0.80138f
C941 a_n2686_12578.t36 GND 0.731265f
C942 a_n2686_12578.t32 GND 0.731265f
C943 a_n2686_12578.t43 GND 0.80138f
C944 a_n2686_12578.t44 GND 0.731265f
C945 a_n2686_12578.t35 GND 0.731265f
C946 a_n2686_12578.t46 GND 0.80138f
C947 a_n2686_12578.t34 GND 0.842114f
C948 a_n2686_12578.t39 GND 0.731265f
C949 a_n2686_12578.n124 GND 0.398404f
C950 a_n2686_12578.t45 GND 0.731265f
C951 a_n2686_12578.t33 GND 0.731265f
C952 a_n2686_12578.t42 GND 0.731265f
C953 a_n2686_12578.n125 GND 0.398404f
C954 a_n2686_12578.t48 GND 0.842114f
C955 a_n2686_12578.t5 GND 0.842114f
C956 a_n2686_12578.t7 GND 0.731265f
C957 a_n2686_12578.n126 GND 0.398404f
C958 a_n2686_12578.t11 GND 0.731265f
C959 a_n2686_12578.t3 GND 0.731265f
C960 a_n2686_12578.t13 GND 0.731265f
C961 a_n2686_12578.n127 GND 0.398404f
C962 a_n2686_12578.t23 GND 0.842114f
C963 a_n2686_12578.n128 GND 0.381069f
C964 a_n2686_12578.n129 GND 0.074231f
C965 a_n2686_12578.n130 GND 0.337772f
C966 a_n2686_12578.n131 GND 0.381069f
C967 a_n2686_12578.n132 GND 0.074231f
C968 a_n2686_12578.n133 GND 0.337772f
C969 a_n2686_12578.t9 GND 0.80138f
C970 a_n2686_12578.t21 GND 0.731265f
C971 a_n2686_12578.n134 GND 0.300249f
C972 a_n2686_12578.t15 GND 0.731265f
C973 a_n2686_12578.t1 GND 0.731265f
C974 a_n2686_12578.t19 GND 0.731265f
C975 a_n2686_12578.n135 GND 0.37178f
C976 a_n2686_12578.t17 GND 0.80138f
C977 a_n2686_12578.n136 GND 0.378046f
C978 a_n2686_12578.n137 GND 0.381069f
C979 a_n2686_12578.n138 GND 0.074231f
C980 a_n2686_12578.n139 GND 0.300249f
C981 a_n2686_12578.n140 GND 0.063218f
C982 a_n2686_12578.n141 GND 0.056324f
C983 a_n2686_12578.n142 GND 0.044455f
C984 a_n2686_12578.n143 GND 0.051105f
C985 a_n2686_12578.n144 GND 0.367987f
C986 a_n2686_12578.n145 GND 0.406786f
C987 a_n2686_12578.n146 GND 0.019663f
C988 a_n2686_12578.n147 GND 0.009653f
C989 a_n2686_12578.n148 GND 0.022816f
C990 a_n2686_12578.n149 GND 0.01022f
C991 a_n2686_12578.n150 GND 0.009653f
C992 a_n2686_12578.n151 GND 0.022816f
C993 a_n2686_12578.n152 GND 0.01022f
C994 a_n2686_12578.n153 GND 0.079425f
C995 a_n2686_12578.t18 GND 0.048956f
C996 a_n2686_12578.n154 GND 0.017112f
C997 a_n2686_12578.n155 GND 0.014506f
C998 a_n2686_12578.n156 GND 0.009653f
C999 a_n2686_12578.n157 GND 0.009653f
C1000 a_n2686_12578.n158 GND 0.01022f
C1001 a_n2686_12578.n159 GND 0.022816f
C1002 a_n2686_12578.n160 GND 0.022816f
C1003 a_n2686_12578.n161 GND 0.01022f
C1004 a_n2686_12578.n162 GND 0.009653f
C1005 a_n2686_12578.n163 GND 0.009653f
C1006 a_n2686_12578.n164 GND 0.01022f
C1007 a_n2686_12578.n165 GND 0.022816f
C1008 a_n2686_12578.n166 GND 0.054978f
C1009 a_n2686_12578.n167 GND 0.01022f
C1010 a_n2686_12578.n168 GND 0.009653f
C1011 a_n2686_12578.n169 GND 0.041521f
C1012 a_n2686_12578.n170 GND 0.034326f
C1013 a_n2686_12578.t2 GND 0.085171f
C1014 a_n2686_12578.t20 GND 0.085171f
C1015 a_n2686_12578.n171 GND 0.524334f
C1016 a_n2686_12578.n172 GND 0.745148f
C1017 a_n2686_12578.t22 GND 0.085171f
C1018 a_n2686_12578.t16 GND 0.085171f
C1019 a_n2686_12578.n173 GND 0.524334f
C1020 a_n2686_12578.n174 GND 0.581063f
C1021 a_n2686_12578.n175 GND 0.019663f
C1022 a_n2686_12578.n176 GND 0.009653f
C1023 a_n2686_12578.n177 GND 0.022816f
C1024 a_n2686_12578.n178 GND 0.01022f
C1025 a_n2686_12578.n179 GND 0.009653f
C1026 a_n2686_12578.n180 GND 0.022816f
C1027 a_n2686_12578.n181 GND 0.01022f
C1028 a_n2686_12578.n182 GND 0.079425f
C1029 a_n2686_12578.t10 GND 0.048956f
C1030 a_n2686_12578.n183 GND 0.017112f
C1031 a_n2686_12578.n184 GND 0.014506f
C1032 a_n2686_12578.n185 GND 0.009653f
C1033 a_n2686_12578.n186 GND 0.009653f
C1034 a_n2686_12578.n187 GND 0.01022f
C1035 a_n2686_12578.n188 GND 0.022816f
C1036 a_n2686_12578.n189 GND 0.022816f
C1037 a_n2686_12578.n190 GND 0.01022f
C1038 a_n2686_12578.n191 GND 0.009653f
C1039 a_n2686_12578.n192 GND 0.009653f
C1040 a_n2686_12578.n193 GND 0.01022f
C1041 a_n2686_12578.n194 GND 0.022816f
C1042 a_n2686_12578.n195 GND 0.054978f
C1043 a_n2686_12578.n196 GND 0.01022f
C1044 a_n2686_12578.n197 GND 0.009653f
C1045 a_n2686_12578.n198 GND 0.041521f
C1046 a_n2686_12578.n199 GND 0.031838f
C1047 a_n2686_12578.n200 GND 0.60505f
C1048 a_n2686_12578.n201 GND 0.540369f
C1049 a_n2686_12578.n202 GND 0.722296f
C1050 a_n2686_12578.n203 GND 0.370438f
C1051 a_n2686_12578.n204 GND 0.371483f
C1052 a_n2686_12578.n205 GND 0.063161f
C1053 a_n2686_12578.n206 GND 0.343545f
C1054 a_n2686_12578.n207 GND 0.300249f
C1055 a_n2686_12578.n208 GND 0.063161f
C1056 a_n2686_12578.t55 GND 0.80138f
C1057 a_n2686_12578.n209 GND 0.371483f
C1058 a_n2686_12578.n210 GND 0.120419f
C1059 a_n2686_12578.n211 GND 0.120419f
C1060 a_n2686_12578.n212 GND 0.371483f
C1061 a_n2686_12578.n213 GND 0.063161f
C1062 a_n2686_12578.n214 GND 0.343545f
C1063 a_n2686_12578.n215 GND 0.300249f
C1064 a_n2686_12578.n216 GND 0.063161f
C1065 a_n2686_12578.t52 GND 0.80138f
C1066 a_n2686_12578.n217 GND 0.371483f
C1067 a_n2686_12578.n218 GND 0.155055f
C1068 a_n2686_12578.n219 GND 0.155055f
C1069 a_n2686_12578.n220 GND 0.371483f
C1070 a_n2686_12578.n221 GND 0.063161f
C1071 a_n2686_12578.n222 GND 0.343545f
C1072 a_n2686_12578.n223 GND 0.300249f
C1073 a_n2686_12578.n224 GND 0.063161f
C1074 a_n2686_12578.t49 GND 0.80138f
C1075 a_n2686_12578.n225 GND 0.371483f
C1076 a_n2686_12578.n226 GND 0.120419f
C1077 a_n2686_12578.n227 GND 0.120419f
C1078 a_n2686_12578.n228 GND 0.371483f
C1079 a_n2686_12578.n229 GND 0.063161f
C1080 a_n2686_12578.n230 GND 0.343545f
C1081 a_n2686_12578.n231 GND 0.300249f
C1082 a_n2686_12578.n232 GND 0.063161f
C1083 a_n2686_12578.t57 GND 0.80138f
C1084 a_n2686_12578.n233 GND 0.371483f
C1085 a_n2686_12578.n234 GND 0.370438f
C1086 a_n2686_12578.n235 GND 0.919537f
C1087 a_n2686_12578.n236 GND 0.381069f
C1088 a_n2686_12578.n237 GND 0.074231f
C1089 a_n2686_12578.n238 GND 0.337772f
C1090 a_n2686_12578.n239 GND 2.6988f
C1091 a_n2686_12578.t31 GND 0.085171f
C1092 a_n2686_12578.t30 GND 0.085171f
C1093 a_n2686_12578.n240 GND 0.745025f
C1094 a_n2686_12578.n241 GND 2.84719f
C1095 a_n2686_12578.n242 GND 2.02113f
C1096 a_n2686_12578.n243 GND 0.743834f
C1097 a_n2686_12578.t0 GND 0.085171f
C1098 a_n2686_8222.n0 GND 0.013106f
C1099 a_n2686_8222.n1 GND 0.011416f
C1100 a_n2686_8222.n2 GND 0.013106f
C1101 a_n2686_8222.n3 GND 0.011416f
C1102 a_n2686_8222.n4 GND 0.013106f
C1103 a_n2686_8222.n5 GND 0.011416f
C1104 a_n2686_8222.n6 GND 0.013106f
C1105 a_n2686_8222.n7 GND 0.011416f
C1106 a_n2686_8222.n8 GND 0.013106f
C1107 a_n2686_8222.n9 GND 0.011416f
C1108 a_n2686_8222.n10 GND 0.013106f
C1109 a_n2686_8222.n11 GND 0.011416f
C1110 a_n2686_8222.n12 GND 0.013106f
C1111 a_n2686_8222.n13 GND 0.011416f
C1112 a_n2686_8222.n14 GND 0.013106f
C1113 a_n2686_8222.n15 GND 0.011416f
C1114 a_n2686_8222.n16 GND 1.7145f
C1115 a_n2686_8222.n17 GND 1.15064f
C1116 a_n2686_8222.n18 GND 0.31216f
C1117 a_n2686_8222.n19 GND 0.31216f
C1118 a_n2686_8222.n20 GND 0.31216f
C1119 a_n2686_8222.n21 GND 0.31216f
C1120 a_n2686_8222.n22 GND 0.31216f
C1121 a_n2686_8222.n23 GND 0.31216f
C1122 a_n2686_8222.n24 GND 0.31216f
C1123 a_n2686_8222.n25 GND 0.31216f
C1124 a_n2686_8222.n26 GND 0.644082f
C1125 a_n2686_8222.n27 GND 0.762343f
C1126 a_n2686_8222.n28 GND 0.045343f
C1127 a_n2686_8222.n29 GND 0.013878f
C1128 a_n2686_8222.n30 GND 0.045343f
C1129 a_n2686_8222.n31 GND 0.013878f
C1130 a_n2686_8222.n32 GND 0.045343f
C1131 a_n2686_8222.n33 GND 0.013878f
C1132 a_n2686_8222.n34 GND 0.045343f
C1133 a_n2686_8222.n35 GND 0.013878f
C1134 a_n2686_8222.n36 GND 0.045343f
C1135 a_n2686_8222.n37 GND 0.013878f
C1136 a_n2686_8222.n38 GND 0.045343f
C1137 a_n2686_8222.n39 GND 0.013878f
C1138 a_n2686_8222.n40 GND 0.045343f
C1139 a_n2686_8222.n41 GND 0.013878f
C1140 a_n2686_8222.n42 GND 0.045343f
C1141 a_n2686_8222.n43 GND 0.013878f
C1142 a_n2686_8222.t8 GND 98.2232f
C1143 a_n2686_8222.n44 GND 0.011295f
C1144 a_n2686_8222.n45 GND 0.005545f
C1145 a_n2686_8222.n46 GND 0.013106f
C1146 a_n2686_8222.n47 GND 0.005871f
C1147 a_n2686_8222.n48 GND 0.005545f
C1148 a_n2686_8222.t20 GND 0.028406f
C1149 a_n2686_8222.n49 GND 0.00983f
C1150 a_n2686_8222.n50 GND 0.005871f
C1151 a_n2686_8222.n51 GND 0.013106f
C1152 a_n2686_8222.n52 GND 0.013106f
C1153 a_n2686_8222.n53 GND 0.005871f
C1154 a_n2686_8222.n54 GND 0.005545f
C1155 a_n2686_8222.n55 GND 0.005545f
C1156 a_n2686_8222.n56 GND 0.005871f
C1157 a_n2686_8222.n57 GND 0.013106f
C1158 a_n2686_8222.n58 GND 0.031582f
C1159 a_n2686_8222.n59 GND 0.005871f
C1160 a_n2686_8222.n60 GND 0.005545f
C1161 a_n2686_8222.n61 GND 0.019719f
C1162 a_n2686_8222.t12 GND 0.048927f
C1163 a_n2686_8222.t6 GND 0.048927f
C1164 a_n2686_8222.n62 GND 0.301206f
C1165 a_n2686_8222.t1 GND 0.048927f
C1166 a_n2686_8222.t4 GND 0.048927f
C1167 a_n2686_8222.n63 GND 0.301206f
C1168 a_n2686_8222.n64 GND 0.011295f
C1169 a_n2686_8222.n65 GND 0.005545f
C1170 a_n2686_8222.n66 GND 0.013106f
C1171 a_n2686_8222.n67 GND 0.005871f
C1172 a_n2686_8222.n68 GND 0.005545f
C1173 a_n2686_8222.t3 GND 0.028406f
C1174 a_n2686_8222.n69 GND 0.00983f
C1175 a_n2686_8222.n70 GND 0.005871f
C1176 a_n2686_8222.n71 GND 0.013106f
C1177 a_n2686_8222.n72 GND 0.013106f
C1178 a_n2686_8222.n73 GND 0.005871f
C1179 a_n2686_8222.n74 GND 0.005545f
C1180 a_n2686_8222.n75 GND 0.005545f
C1181 a_n2686_8222.n76 GND 0.005871f
C1182 a_n2686_8222.n77 GND 0.013106f
C1183 a_n2686_8222.n78 GND 0.031582f
C1184 a_n2686_8222.n79 GND 0.005871f
C1185 a_n2686_8222.n80 GND 0.005545f
C1186 a_n2686_8222.n81 GND 0.01829f
C1187 a_n2686_8222.n82 GND 0.011295f
C1188 a_n2686_8222.n83 GND 0.005545f
C1189 a_n2686_8222.n84 GND 0.013106f
C1190 a_n2686_8222.n85 GND 0.005871f
C1191 a_n2686_8222.n86 GND 0.005545f
C1192 a_n2686_8222.t16 GND 0.028406f
C1193 a_n2686_8222.n87 GND 0.00983f
C1194 a_n2686_8222.n88 GND 0.005871f
C1195 a_n2686_8222.n89 GND 0.013106f
C1196 a_n2686_8222.n90 GND 0.013106f
C1197 a_n2686_8222.n91 GND 0.005871f
C1198 a_n2686_8222.n92 GND 0.005545f
C1199 a_n2686_8222.n93 GND 0.005545f
C1200 a_n2686_8222.n94 GND 0.005871f
C1201 a_n2686_8222.n95 GND 0.013106f
C1202 a_n2686_8222.n96 GND 0.031582f
C1203 a_n2686_8222.n97 GND 0.005871f
C1204 a_n2686_8222.n98 GND 0.005545f
C1205 a_n2686_8222.n99 GND 0.019719f
C1206 a_n2686_8222.t7 GND 0.048927f
C1207 a_n2686_8222.t5 GND 0.048927f
C1208 a_n2686_8222.n100 GND 0.301206f
C1209 a_n2686_8222.n101 GND 0.011295f
C1210 a_n2686_8222.n102 GND 0.005545f
C1211 a_n2686_8222.n103 GND 0.013106f
C1212 a_n2686_8222.n104 GND 0.005871f
C1213 a_n2686_8222.n105 GND 0.005545f
C1214 a_n2686_8222.t0 GND 0.028406f
C1215 a_n2686_8222.n106 GND 0.00983f
C1216 a_n2686_8222.n107 GND 0.005871f
C1217 a_n2686_8222.n108 GND 0.013106f
C1218 a_n2686_8222.n109 GND 0.013106f
C1219 a_n2686_8222.n110 GND 0.005871f
C1220 a_n2686_8222.n111 GND 0.005545f
C1221 a_n2686_8222.n112 GND 0.005545f
C1222 a_n2686_8222.n113 GND 0.005871f
C1223 a_n2686_8222.n114 GND 0.013106f
C1224 a_n2686_8222.n115 GND 0.031582f
C1225 a_n2686_8222.n116 GND 0.005871f
C1226 a_n2686_8222.n117 GND 0.005545f
C1227 a_n2686_8222.n118 GND 0.01829f
C1228 a_n2686_8222.n119 GND 0.011295f
C1229 a_n2686_8222.n120 GND 0.005545f
C1230 a_n2686_8222.n121 GND 0.013106f
C1231 a_n2686_8222.n122 GND 0.005871f
C1232 a_n2686_8222.n123 GND 0.005545f
C1233 a_n2686_8222.t14 GND 0.028406f
C1234 a_n2686_8222.n124 GND 0.00983f
C1235 a_n2686_8222.n125 GND 0.005871f
C1236 a_n2686_8222.n126 GND 0.013106f
C1237 a_n2686_8222.n127 GND 0.013106f
C1238 a_n2686_8222.n128 GND 0.005871f
C1239 a_n2686_8222.n129 GND 0.005545f
C1240 a_n2686_8222.n130 GND 0.005545f
C1241 a_n2686_8222.n131 GND 0.005871f
C1242 a_n2686_8222.n132 GND 0.013106f
C1243 a_n2686_8222.n133 GND 0.031582f
C1244 a_n2686_8222.n134 GND 0.005871f
C1245 a_n2686_8222.n135 GND 0.005545f
C1246 a_n2686_8222.n136 GND 0.01829f
C1247 a_n2686_8222.t9 GND 0.048927f
C1248 a_n2686_8222.t13 GND 0.048927f
C1249 a_n2686_8222.n137 GND 0.301206f
C1250 a_n2686_8222.n138 GND 0.011295f
C1251 a_n2686_8222.n139 GND 0.005545f
C1252 a_n2686_8222.n140 GND 0.013106f
C1253 a_n2686_8222.n141 GND 0.005871f
C1254 a_n2686_8222.n142 GND 0.005545f
C1255 a_n2686_8222.t10 GND 0.028406f
C1256 a_n2686_8222.n143 GND 0.00983f
C1257 a_n2686_8222.n144 GND 0.005871f
C1258 a_n2686_8222.n145 GND 0.013106f
C1259 a_n2686_8222.n146 GND 0.013106f
C1260 a_n2686_8222.n147 GND 0.005871f
C1261 a_n2686_8222.n148 GND 0.005545f
C1262 a_n2686_8222.n149 GND 0.005545f
C1263 a_n2686_8222.n150 GND 0.005871f
C1264 a_n2686_8222.n151 GND 0.013106f
C1265 a_n2686_8222.n152 GND 0.031582f
C1266 a_n2686_8222.n153 GND 0.005871f
C1267 a_n2686_8222.n154 GND 0.005545f
C1268 a_n2686_8222.n155 GND 0.01829f
C1269 a_n2686_8222.n156 GND 1.23733f
C1270 a_n2686_8222.n157 GND 0.011295f
C1271 a_n2686_8222.n158 GND 0.005545f
C1272 a_n2686_8222.n159 GND 0.013106f
C1273 a_n2686_8222.n160 GND 0.005871f
C1274 a_n2686_8222.n161 GND 0.005545f
C1275 a_n2686_8222.t11 GND 0.028406f
C1276 a_n2686_8222.n162 GND 0.00983f
C1277 a_n2686_8222.n163 GND 0.005871f
C1278 a_n2686_8222.n164 GND 0.013106f
C1279 a_n2686_8222.n165 GND 0.013106f
C1280 a_n2686_8222.n166 GND 0.005871f
C1281 a_n2686_8222.n167 GND 0.005545f
C1282 a_n2686_8222.n168 GND 0.005545f
C1283 a_n2686_8222.n169 GND 0.005871f
C1284 a_n2686_8222.n170 GND 0.013106f
C1285 a_n2686_8222.n171 GND 0.031582f
C1286 a_n2686_8222.n172 GND 0.005871f
C1287 a_n2686_8222.n173 GND 0.005545f
C1288 a_n2686_8222.n174 GND 0.019719f
C1289 a_n2686_8222.t2 GND 0.048927f
C1290 a_n2686_8222.t17 GND 0.048927f
C1291 a_n2686_8222.n175 GND 0.301206f
C1292 a_n2686_8222.t18 GND 0.048927f
C1293 a_n2686_8222.t19 GND 0.048927f
C1294 a_n2686_8222.n176 GND 0.301206f
C1295 a_n2686_8222.n177 GND 0.011295f
C1296 a_n2686_8222.n178 GND 0.005545f
C1297 a_n2686_8222.n179 GND 0.013106f
C1298 a_n2686_8222.n180 GND 0.005871f
C1299 a_n2686_8222.n181 GND 0.005545f
C1300 a_n2686_8222.t15 GND 0.028406f
C1301 a_n2686_8222.n182 GND 0.00983f
C1302 a_n2686_8222.n183 GND 0.005871f
C1303 a_n2686_8222.n184 GND 0.013106f
C1304 a_n2686_8222.n185 GND 0.013106f
C1305 a_n2686_8222.n186 GND 0.005871f
C1306 a_n2686_8222.n187 GND 0.005545f
C1307 a_n2686_8222.n188 GND 0.005545f
C1308 a_n2686_8222.n189 GND 0.005871f
C1309 a_n2686_8222.n190 GND 0.013106f
C1310 a_n2686_8222.n191 GND 0.031582f
C1311 a_n2686_8222.n192 GND 0.005871f
C1312 a_n2686_8222.n193 GND 0.005545f
C1313 a_n2686_8222.n194 GND 0.01829f
C1314 a_n2686_8222.n195 GND 1.73078f
C1315 VDD.t201 GND 0.021885f
C1316 VDD.t199 GND 0.021885f
C1317 VDD.n0 GND 0.158137f
C1318 VDD.t203 GND 0.021885f
C1319 VDD.t205 GND 0.021885f
C1320 VDD.n1 GND 0.157401f
C1321 VDD.n2 GND 0.286508f
C1322 VDD.t1 GND 0.021885f
C1323 VDD.t94 GND 0.021885f
C1324 VDD.n3 GND 0.157401f
C1325 VDD.n4 GND 0.146379f
C1326 VDD.t89 GND 0.021885f
C1327 VDD.t207 GND 0.021885f
C1328 VDD.n5 GND 0.157401f
C1329 VDD.n6 GND 0.132531f
C1330 VDD.t85 GND 0.021885f
C1331 VDD.t196 GND 0.021885f
C1332 VDD.n7 GND 0.158137f
C1333 VDD.t213 GND 0.021885f
C1334 VDD.t194 GND 0.021885f
C1335 VDD.n8 GND 0.157401f
C1336 VDD.n9 GND 0.286508f
C1337 VDD.t81 GND 0.021885f
C1338 VDD.t215 GND 0.021885f
C1339 VDD.n10 GND 0.157401f
C1340 VDD.n11 GND 0.146379f
C1341 VDD.t209 GND 0.021885f
C1342 VDD.t87 GND 0.021885f
C1343 VDD.n12 GND 0.157401f
C1344 VDD.n13 GND 0.132531f
C1345 VDD.n14 GND 0.091271f
C1346 VDD.n15 GND 2.31548f
C1347 VDD.n16 GND 0.004974f
C1348 VDD.n17 GND 0.004616f
C1349 VDD.n18 GND 0.002553f
C1350 VDD.n19 GND 0.005863f
C1351 VDD.n20 GND 0.00248f
C1352 VDD.n21 GND 0.002626f
C1353 VDD.n22 GND 0.004616f
C1354 VDD.n23 GND 0.00248f
C1355 VDD.n24 GND 0.005863f
C1356 VDD.n25 GND 0.002626f
C1357 VDD.n26 GND 0.004616f
C1358 VDD.n27 GND 0.00248f
C1359 VDD.n28 GND 0.004397f
C1360 VDD.n29 GND 0.00441f
C1361 VDD.t177 GND 0.012595f
C1362 VDD.n30 GND 0.028025f
C1363 VDD.n31 GND 0.145847f
C1364 VDD.n32 GND 0.00248f
C1365 VDD.n33 GND 0.002626f
C1366 VDD.n34 GND 0.005863f
C1367 VDD.n35 GND 0.005863f
C1368 VDD.n36 GND 0.002626f
C1369 VDD.n37 GND 0.00248f
C1370 VDD.n38 GND 0.004616f
C1371 VDD.n39 GND 0.004616f
C1372 VDD.n40 GND 0.00248f
C1373 VDD.n41 GND 0.002626f
C1374 VDD.n42 GND 0.005863f
C1375 VDD.n43 GND 0.005863f
C1376 VDD.n44 GND 0.002626f
C1377 VDD.n45 GND 0.00248f
C1378 VDD.n46 GND 0.004616f
C1379 VDD.n47 GND 0.004616f
C1380 VDD.n48 GND 0.00248f
C1381 VDD.n49 GND 0.002626f
C1382 VDD.n50 GND 0.005863f
C1383 VDD.n51 GND 0.005863f
C1384 VDD.n52 GND 0.013861f
C1385 VDD.n53 GND 0.002553f
C1386 VDD.n54 GND 0.00248f
C1387 VDD.n55 GND 0.011931f
C1388 VDD.n56 GND 0.008658f
C1389 VDD.t184 GND 0.029181f
C1390 VDD.t165 GND 0.029181f
C1391 VDD.n57 GND 0.20055f
C1392 VDD.n58 GND 0.195838f
C1393 VDD.t187 GND 0.029181f
C1394 VDD.t98 GND 0.029181f
C1395 VDD.n59 GND 0.20055f
C1396 VDD.n60 GND 0.152908f
C1397 VDD.t175 GND 0.029181f
C1398 VDD.t156 GND 0.029181f
C1399 VDD.n61 GND 0.20055f
C1400 VDD.n62 GND 0.152908f
C1401 VDD.t111 GND 0.029181f
C1402 VDD.t182 GND 0.029181f
C1403 VDD.n63 GND 0.20055f
C1404 VDD.n64 GND 0.152908f
C1405 VDD.t166 GND 0.029181f
C1406 VDD.t146 GND 0.029181f
C1407 VDD.n65 GND 0.20055f
C1408 VDD.n66 GND 0.152908f
C1409 VDD.n67 GND 0.004974f
C1410 VDD.n68 GND 0.004616f
C1411 VDD.n69 GND 0.002553f
C1412 VDD.n70 GND 0.005863f
C1413 VDD.n71 GND 0.00248f
C1414 VDD.n72 GND 0.002626f
C1415 VDD.n73 GND 0.004616f
C1416 VDD.n74 GND 0.00248f
C1417 VDD.n75 GND 0.005863f
C1418 VDD.n76 GND 0.002626f
C1419 VDD.n77 GND 0.004616f
C1420 VDD.n78 GND 0.00248f
C1421 VDD.n79 GND 0.004397f
C1422 VDD.n80 GND 0.00441f
C1423 VDD.t128 GND 0.012595f
C1424 VDD.n81 GND 0.028025f
C1425 VDD.n82 GND 0.145847f
C1426 VDD.n83 GND 0.00248f
C1427 VDD.n84 GND 0.002626f
C1428 VDD.n85 GND 0.005863f
C1429 VDD.n86 GND 0.005863f
C1430 VDD.n87 GND 0.002626f
C1431 VDD.n88 GND 0.00248f
C1432 VDD.n89 GND 0.004616f
C1433 VDD.n90 GND 0.004616f
C1434 VDD.n91 GND 0.00248f
C1435 VDD.n92 GND 0.002626f
C1436 VDD.n93 GND 0.005863f
C1437 VDD.n94 GND 0.005863f
C1438 VDD.n95 GND 0.002626f
C1439 VDD.n96 GND 0.00248f
C1440 VDD.n97 GND 0.004616f
C1441 VDD.n98 GND 0.004616f
C1442 VDD.n99 GND 0.00248f
C1443 VDD.n100 GND 0.002626f
C1444 VDD.n101 GND 0.005863f
C1445 VDD.n102 GND 0.005863f
C1446 VDD.n103 GND 0.013861f
C1447 VDD.n104 GND 0.002553f
C1448 VDD.n105 GND 0.00248f
C1449 VDD.n106 GND 0.011931f
C1450 VDD.n107 GND 0.008068f
C1451 VDD.n108 GND 0.117377f
C1452 VDD.n109 GND 0.004974f
C1453 VDD.n110 GND 0.004616f
C1454 VDD.n111 GND 0.002553f
C1455 VDD.n112 GND 0.005863f
C1456 VDD.n113 GND 0.00248f
C1457 VDD.n114 GND 0.002626f
C1458 VDD.n115 GND 0.004616f
C1459 VDD.n116 GND 0.00248f
C1460 VDD.n117 GND 0.005863f
C1461 VDD.n118 GND 0.002626f
C1462 VDD.n119 GND 0.004616f
C1463 VDD.n120 GND 0.00248f
C1464 VDD.n121 GND 0.004397f
C1465 VDD.n122 GND 0.00441f
C1466 VDD.t148 GND 0.012595f
C1467 VDD.n123 GND 0.028025f
C1468 VDD.n124 GND 0.145847f
C1469 VDD.n125 GND 0.00248f
C1470 VDD.n126 GND 0.002626f
C1471 VDD.n127 GND 0.005863f
C1472 VDD.n128 GND 0.005863f
C1473 VDD.n129 GND 0.002626f
C1474 VDD.n130 GND 0.00248f
C1475 VDD.n131 GND 0.004616f
C1476 VDD.n132 GND 0.004616f
C1477 VDD.n133 GND 0.00248f
C1478 VDD.n134 GND 0.002626f
C1479 VDD.n135 GND 0.005863f
C1480 VDD.n136 GND 0.005863f
C1481 VDD.n137 GND 0.002626f
C1482 VDD.n138 GND 0.00248f
C1483 VDD.n139 GND 0.004616f
C1484 VDD.n140 GND 0.004616f
C1485 VDD.n141 GND 0.00248f
C1486 VDD.n142 GND 0.002626f
C1487 VDD.n143 GND 0.005863f
C1488 VDD.n144 GND 0.005863f
C1489 VDD.n145 GND 0.013861f
C1490 VDD.n146 GND 0.002553f
C1491 VDD.n147 GND 0.00248f
C1492 VDD.n148 GND 0.011931f
C1493 VDD.n149 GND 0.008658f
C1494 VDD.t158 GND 0.029181f
C1495 VDD.t189 GND 0.029181f
C1496 VDD.n150 GND 0.20055f
C1497 VDD.n151 GND 0.195838f
C1498 VDD.t173 GND 0.029181f
C1499 VDD.t179 GND 0.029181f
C1500 VDD.n152 GND 0.20055f
C1501 VDD.n153 GND 0.152908f
C1502 VDD.t120 GND 0.029181f
C1503 VDD.t161 GND 0.029181f
C1504 VDD.n154 GND 0.20055f
C1505 VDD.n155 GND 0.152908f
C1506 VDD.t112 GND 0.029181f
C1507 VDD.t140 GND 0.029181f
C1508 VDD.n156 GND 0.20055f
C1509 VDD.n157 GND 0.152908f
C1510 VDD.t181 GND 0.029181f
C1511 VDD.t123 GND 0.029181f
C1512 VDD.n158 GND 0.20055f
C1513 VDD.n159 GND 0.152908f
C1514 VDD.n160 GND 0.004974f
C1515 VDD.n161 GND 0.004616f
C1516 VDD.n162 GND 0.002553f
C1517 VDD.n163 GND 0.005863f
C1518 VDD.n164 GND 0.00248f
C1519 VDD.n165 GND 0.002626f
C1520 VDD.n166 GND 0.004616f
C1521 VDD.n167 GND 0.00248f
C1522 VDD.n168 GND 0.005863f
C1523 VDD.n169 GND 0.002626f
C1524 VDD.n170 GND 0.004616f
C1525 VDD.n171 GND 0.00248f
C1526 VDD.n172 GND 0.004397f
C1527 VDD.n173 GND 0.00441f
C1528 VDD.t138 GND 0.012595f
C1529 VDD.n174 GND 0.028025f
C1530 VDD.n175 GND 0.145847f
C1531 VDD.n176 GND 0.00248f
C1532 VDD.n177 GND 0.002626f
C1533 VDD.n178 GND 0.005863f
C1534 VDD.n179 GND 0.005863f
C1535 VDD.n180 GND 0.002626f
C1536 VDD.n181 GND 0.00248f
C1537 VDD.n182 GND 0.004616f
C1538 VDD.n183 GND 0.004616f
C1539 VDD.n184 GND 0.00248f
C1540 VDD.n185 GND 0.002626f
C1541 VDD.n186 GND 0.005863f
C1542 VDD.n187 GND 0.005863f
C1543 VDD.n188 GND 0.002626f
C1544 VDD.n189 GND 0.00248f
C1545 VDD.n190 GND 0.004616f
C1546 VDD.n191 GND 0.004616f
C1547 VDD.n192 GND 0.00248f
C1548 VDD.n193 GND 0.002626f
C1549 VDD.n194 GND 0.005863f
C1550 VDD.n195 GND 0.005863f
C1551 VDD.n196 GND 0.013861f
C1552 VDD.n197 GND 0.002553f
C1553 VDD.n198 GND 0.00248f
C1554 VDD.n199 GND 0.011931f
C1555 VDD.n200 GND 0.008068f
C1556 VDD.n201 GND 0.06915f
C1557 VDD.n202 GND 0.376011f
C1558 VDD.n203 GND 0.004974f
C1559 VDD.n204 GND 0.004616f
C1560 VDD.n205 GND 0.002553f
C1561 VDD.n206 GND 0.005863f
C1562 VDD.n207 GND 0.00248f
C1563 VDD.n208 GND 0.002626f
C1564 VDD.n209 GND 0.004616f
C1565 VDD.n210 GND 0.00248f
C1566 VDD.n211 GND 0.005863f
C1567 VDD.n212 GND 0.002626f
C1568 VDD.n213 GND 0.004616f
C1569 VDD.n214 GND 0.00248f
C1570 VDD.n215 GND 0.004397f
C1571 VDD.n216 GND 0.00441f
C1572 VDD.t160 GND 0.012595f
C1573 VDD.n217 GND 0.028025f
C1574 VDD.n218 GND 0.145847f
C1575 VDD.n219 GND 0.00248f
C1576 VDD.n220 GND 0.002626f
C1577 VDD.n221 GND 0.005863f
C1578 VDD.n222 GND 0.005863f
C1579 VDD.n223 GND 0.002626f
C1580 VDD.n224 GND 0.00248f
C1581 VDD.n225 GND 0.004616f
C1582 VDD.n226 GND 0.004616f
C1583 VDD.n227 GND 0.00248f
C1584 VDD.n228 GND 0.002626f
C1585 VDD.n229 GND 0.005863f
C1586 VDD.n230 GND 0.005863f
C1587 VDD.n231 GND 0.002626f
C1588 VDD.n232 GND 0.00248f
C1589 VDD.n233 GND 0.004616f
C1590 VDD.n234 GND 0.004616f
C1591 VDD.n235 GND 0.00248f
C1592 VDD.n236 GND 0.002626f
C1593 VDD.n237 GND 0.005863f
C1594 VDD.n238 GND 0.005863f
C1595 VDD.n239 GND 0.013861f
C1596 VDD.n240 GND 0.002553f
C1597 VDD.n241 GND 0.00248f
C1598 VDD.n242 GND 0.011931f
C1599 VDD.n243 GND 0.008658f
C1600 VDD.t169 GND 0.029181f
C1601 VDD.t109 GND 0.029181f
C1602 VDD.n244 GND 0.20055f
C1603 VDD.n245 GND 0.195838f
C1604 VDD.t180 GND 0.029181f
C1605 VDD.t190 GND 0.029181f
C1606 VDD.n246 GND 0.20055f
C1607 VDD.n247 GND 0.152908f
C1608 VDD.t133 GND 0.029181f
C1609 VDD.t170 GND 0.029181f
C1610 VDD.n248 GND 0.20055f
C1611 VDD.n249 GND 0.152908f
C1612 VDD.t121 GND 0.029181f
C1613 VDD.t151 GND 0.029181f
C1614 VDD.n250 GND 0.20055f
C1615 VDD.n251 GND 0.152908f
C1616 VDD.t96 GND 0.029181f
C1617 VDD.t134 GND 0.029181f
C1618 VDD.n252 GND 0.20055f
C1619 VDD.n253 GND 0.152908f
C1620 VDD.n254 GND 0.004974f
C1621 VDD.n255 GND 0.004616f
C1622 VDD.n256 GND 0.002553f
C1623 VDD.n257 GND 0.005863f
C1624 VDD.n258 GND 0.00248f
C1625 VDD.n259 GND 0.002626f
C1626 VDD.n260 GND 0.004616f
C1627 VDD.n261 GND 0.00248f
C1628 VDD.n262 GND 0.005863f
C1629 VDD.n263 GND 0.002626f
C1630 VDD.n264 GND 0.004616f
C1631 VDD.n265 GND 0.00248f
C1632 VDD.n266 GND 0.004397f
C1633 VDD.n267 GND 0.00441f
C1634 VDD.t149 GND 0.012595f
C1635 VDD.n268 GND 0.028025f
C1636 VDD.n269 GND 0.145847f
C1637 VDD.n270 GND 0.00248f
C1638 VDD.n271 GND 0.002626f
C1639 VDD.n272 GND 0.005863f
C1640 VDD.n273 GND 0.005863f
C1641 VDD.n274 GND 0.002626f
C1642 VDD.n275 GND 0.00248f
C1643 VDD.n276 GND 0.004616f
C1644 VDD.n277 GND 0.004616f
C1645 VDD.n278 GND 0.00248f
C1646 VDD.n279 GND 0.002626f
C1647 VDD.n280 GND 0.005863f
C1648 VDD.n281 GND 0.005863f
C1649 VDD.n282 GND 0.002626f
C1650 VDD.n283 GND 0.00248f
C1651 VDD.n284 GND 0.004616f
C1652 VDD.n285 GND 0.004616f
C1653 VDD.n286 GND 0.00248f
C1654 VDD.n287 GND 0.002626f
C1655 VDD.n288 GND 0.005863f
C1656 VDD.n289 GND 0.005863f
C1657 VDD.n290 GND 0.013861f
C1658 VDD.n291 GND 0.002553f
C1659 VDD.n292 GND 0.00248f
C1660 VDD.n293 GND 0.011931f
C1661 VDD.n294 GND 0.008068f
C1662 VDD.n295 GND 0.06915f
C1663 VDD.n296 GND 0.322101f
C1664 VDD.n297 GND 0.009033f
C1665 VDD.n298 GND 0.009033f
C1666 VDD.n299 GND 0.007295f
C1667 VDD.n300 GND 0.007295f
C1668 VDD.n301 GND 0.009064f
C1669 VDD.n302 GND 0.009064f
C1670 VDD.n303 GND 0.511885f
C1671 VDD.n304 GND 0.009064f
C1672 VDD.n305 GND 0.009064f
C1673 VDD.n306 GND 0.009064f
C1674 VDD.n307 GND 0.765903f
C1675 VDD.n308 GND 0.009064f
C1676 VDD.n309 GND 0.009064f
C1677 VDD.n310 GND 0.009064f
C1678 VDD.n311 GND 0.009064f
C1679 VDD.n312 GND 0.007295f
C1680 VDD.n313 GND 0.009064f
C1681 VDD.t110 GND 0.384876f
C1682 VDD.n314 GND 0.009064f
C1683 VDD.n315 GND 0.009064f
C1684 VDD.n316 GND 0.009064f
C1685 VDD.t139 GND 0.384876f
C1686 VDD.n317 GND 0.009064f
C1687 VDD.n318 GND 0.009064f
C1688 VDD.n319 GND 0.009064f
C1689 VDD.n320 GND 0.009064f
C1690 VDD.n321 GND 0.009064f
C1691 VDD.n322 GND 0.007295f
C1692 VDD.n323 GND 0.009064f
C1693 VDD.n324 GND 0.519582f
C1694 VDD.n325 GND 0.009064f
C1695 VDD.n326 GND 0.009064f
C1696 VDD.n327 GND 0.009064f
C1697 VDD.n328 GND 0.758205f
C1698 VDD.n329 GND 0.009064f
C1699 VDD.n330 GND 0.009064f
C1700 VDD.n331 GND 0.009064f
C1701 VDD.n332 GND 0.009064f
C1702 VDD.n333 GND 0.009064f
C1703 VDD.n334 GND 0.007295f
C1704 VDD.n335 GND 0.009064f
C1705 VDD.t122 GND 0.384876f
C1706 VDD.n336 GND 0.009064f
C1707 VDD.n337 GND 0.009064f
C1708 VDD.n338 GND 0.009064f
C1709 VDD.t127 GND 0.384876f
C1710 VDD.n339 GND 0.009064f
C1711 VDD.n340 GND 0.009064f
C1712 VDD.n341 GND 0.009064f
C1713 VDD.n342 GND 0.009064f
C1714 VDD.n343 GND 0.009064f
C1715 VDD.n344 GND 0.007295f
C1716 VDD.n345 GND 0.009064f
C1717 VDD.n346 GND 0.52728f
C1718 VDD.n347 GND 0.009064f
C1719 VDD.n348 GND 0.009064f
C1720 VDD.n349 GND 0.009064f
C1721 VDD.n350 GND 0.565767f
C1722 VDD.n351 GND 0.009064f
C1723 VDD.n352 GND 0.009064f
C1724 VDD.n353 GND 0.009064f
C1725 VDD.n354 GND 0.009064f
C1726 VDD.n355 GND 0.009064f
C1727 VDD.n356 GND 0.006055f
C1728 VDD.n357 GND 0.020998f
C1729 VDD.t18 GND 0.384876f
C1730 VDD.n358 GND 0.009064f
C1731 VDD.n359 GND 0.020998f
C1732 VDD.n391 GND 0.009064f
C1733 VDD.t41 GND 0.111507f
C1734 VDD.t40 GND 0.123568f
C1735 VDD.t39 GND 0.30702f
C1736 VDD.n392 GND 0.203209f
C1737 VDD.n393 GND 0.158699f
C1738 VDD.n394 GND 0.011271f
C1739 VDD.n395 GND 0.009064f
C1740 VDD.n396 GND 0.007295f
C1741 VDD.n397 GND 0.009064f
C1742 VDD.n398 GND 0.007295f
C1743 VDD.n399 GND 0.009064f
C1744 VDD.n400 GND 0.007295f
C1745 VDD.n401 GND 0.009064f
C1746 VDD.n402 GND 0.007295f
C1747 VDD.n403 GND 0.009064f
C1748 VDD.n404 GND 0.007295f
C1749 VDD.n405 GND 0.009064f
C1750 VDD.t20 GND 0.111507f
C1751 VDD.t19 GND 0.123568f
C1752 VDD.t17 GND 0.30702f
C1753 VDD.n406 GND 0.203209f
C1754 VDD.n407 GND 0.158699f
C1755 VDD.n408 GND 0.007295f
C1756 VDD.n409 GND 0.009064f
C1757 VDD.n410 GND 0.007295f
C1758 VDD.n411 GND 0.009064f
C1759 VDD.n412 GND 0.007295f
C1760 VDD.n413 GND 0.009064f
C1761 VDD.n414 GND 0.007295f
C1762 VDD.n415 GND 0.009064f
C1763 VDD.n416 GND 0.007295f
C1764 VDD.n417 GND 0.009064f
C1765 VDD.t35 GND 0.111507f
C1766 VDD.t34 GND 0.123568f
C1767 VDD.t33 GND 0.30702f
C1768 VDD.n418 GND 0.203209f
C1769 VDD.n419 GND 0.158699f
C1770 VDD.n420 GND 0.014919f
C1771 VDD.n421 GND 0.009064f
C1772 VDD.n422 GND 0.007295f
C1773 VDD.n423 GND 0.009064f
C1774 VDD.n424 GND 0.007295f
C1775 VDD.n425 GND 0.009064f
C1776 VDD.n426 GND 0.007295f
C1777 VDD.n427 GND 0.009064f
C1778 VDD.n428 GND 0.007295f
C1779 VDD.n429 GND 0.009064f
C1780 VDD.n430 GND 0.020998f
C1781 VDD.n431 GND 0.021239f
C1782 VDD.n432 GND 0.021239f
C1783 VDD.n433 GND 0.006055f
C1784 VDD.n434 GND 0.007295f
C1785 VDD.n435 GND 0.009064f
C1786 VDD.n436 GND 0.009064f
C1787 VDD.n437 GND 0.007295f
C1788 VDD.n438 GND 0.009064f
C1789 VDD.n439 GND 0.009064f
C1790 VDD.n440 GND 0.009064f
C1791 VDD.n441 GND 0.009064f
C1792 VDD.n442 GND 0.009064f
C1793 VDD.n443 GND 0.007295f
C1794 VDD.n444 GND 0.007295f
C1795 VDD.n445 GND 0.009064f
C1796 VDD.n446 GND 0.009064f
C1797 VDD.n447 GND 0.007295f
C1798 VDD.n448 GND 0.009064f
C1799 VDD.n449 GND 0.009064f
C1800 VDD.n450 GND 0.009064f
C1801 VDD.n451 GND 0.009064f
C1802 VDD.n452 GND 0.009064f
C1803 VDD.n453 GND 0.007295f
C1804 VDD.n454 GND 0.007295f
C1805 VDD.n455 GND 0.009064f
C1806 VDD.n456 GND 0.009064f
C1807 VDD.n457 GND 0.007295f
C1808 VDD.n458 GND 0.009064f
C1809 VDD.n459 GND 0.009064f
C1810 VDD.n460 GND 0.009064f
C1811 VDD.n461 GND 0.009064f
C1812 VDD.n462 GND 0.009064f
C1813 VDD.n463 GND 0.007295f
C1814 VDD.n464 GND 0.007295f
C1815 VDD.n465 GND 0.009064f
C1816 VDD.n466 GND 0.009064f
C1817 VDD.n467 GND 0.007295f
C1818 VDD.n468 GND 0.009064f
C1819 VDD.n469 GND 0.009064f
C1820 VDD.n470 GND 0.009064f
C1821 VDD.n471 GND 0.009064f
C1822 VDD.n472 GND 0.009064f
C1823 VDD.n473 GND 0.007295f
C1824 VDD.n474 GND 0.007295f
C1825 VDD.n475 GND 0.009064f
C1826 VDD.n476 GND 0.009064f
C1827 VDD.n477 GND 0.006091f
C1828 VDD.n478 GND 0.009064f
C1829 VDD.n479 GND 0.009064f
C1830 VDD.n480 GND 0.009064f
C1831 VDD.n481 GND 0.009064f
C1832 VDD.n482 GND 0.009064f
C1833 VDD.n483 GND 0.006091f
C1834 VDD.n484 GND 0.007295f
C1835 VDD.n485 GND 0.009064f
C1836 VDD.n486 GND 0.009064f
C1837 VDD.n487 GND 0.007295f
C1838 VDD.n488 GND 0.009064f
C1839 VDD.n489 GND 0.009064f
C1840 VDD.n490 GND 0.009064f
C1841 VDD.n491 GND 0.009064f
C1842 VDD.n492 GND 0.009064f
C1843 VDD.n493 GND 0.007295f
C1844 VDD.n494 GND 0.007295f
C1845 VDD.n495 GND 0.009064f
C1846 VDD.n496 GND 0.009064f
C1847 VDD.n497 GND 0.007295f
C1848 VDD.n498 GND 0.009064f
C1849 VDD.n499 GND 0.009064f
C1850 VDD.n500 GND 0.009064f
C1851 VDD.n501 GND 0.009064f
C1852 VDD.n502 GND 0.009064f
C1853 VDD.n503 GND 0.007295f
C1854 VDD.n504 GND 0.007295f
C1855 VDD.n505 GND 0.009064f
C1856 VDD.n506 GND 0.009064f
C1857 VDD.n507 GND 0.007295f
C1858 VDD.n508 GND 0.009064f
C1859 VDD.n509 GND 0.009064f
C1860 VDD.n510 GND 0.009064f
C1861 VDD.n511 GND 0.009064f
C1862 VDD.n512 GND 0.009064f
C1863 VDD.n513 GND 0.007295f
C1864 VDD.n514 GND 0.007295f
C1865 VDD.n515 GND 0.009064f
C1866 VDD.n516 GND 0.009064f
C1867 VDD.n517 GND 0.007295f
C1868 VDD.n518 GND 0.009064f
C1869 VDD.n519 GND 0.009064f
C1870 VDD.n520 GND 0.009064f
C1871 VDD.n521 GND 0.009064f
C1872 VDD.n522 GND 0.009064f
C1873 VDD.n523 GND 0.007295f
C1874 VDD.n524 GND 0.007295f
C1875 VDD.n525 GND 0.009064f
C1876 VDD.n526 GND 0.009064f
C1877 VDD.n527 GND 0.007295f
C1878 VDD.n528 GND 0.009064f
C1879 VDD.n529 GND 0.009064f
C1880 VDD.n530 GND 0.009064f
C1881 VDD.n531 GND 0.009064f
C1882 VDD.n532 GND 0.009064f
C1883 VDD.n533 GND 0.004961f
C1884 VDD.n534 GND 0.014919f
C1885 VDD.n535 GND 0.009064f
C1886 VDD.n536 GND 0.009064f
C1887 VDD.n537 GND 0.007222f
C1888 VDD.n538 GND 0.009064f
C1889 VDD.n539 GND 0.009064f
C1890 VDD.n540 GND 0.009064f
C1891 VDD.n541 GND 0.009064f
C1892 VDD.n542 GND 0.009064f
C1893 VDD.n543 GND 0.007295f
C1894 VDD.n544 GND 0.007295f
C1895 VDD.n545 GND 0.009064f
C1896 VDD.n546 GND 0.009064f
C1897 VDD.n547 GND 0.007295f
C1898 VDD.n548 GND 0.009064f
C1899 VDD.n549 GND 0.009064f
C1900 VDD.n550 GND 0.009064f
C1901 VDD.n551 GND 0.009064f
C1902 VDD.n552 GND 0.009064f
C1903 VDD.n553 GND 0.007295f
C1904 VDD.n554 GND 0.007295f
C1905 VDD.n555 GND 0.009064f
C1906 VDD.n556 GND 0.009064f
C1907 VDD.n557 GND 0.007295f
C1908 VDD.n558 GND 0.009064f
C1909 VDD.n559 GND 0.009064f
C1910 VDD.n560 GND 0.009064f
C1911 VDD.n561 GND 0.009064f
C1912 VDD.n562 GND 0.009064f
C1913 VDD.n563 GND 0.007295f
C1914 VDD.n564 GND 0.007295f
C1915 VDD.n565 GND 0.009064f
C1916 VDD.n566 GND 0.009064f
C1917 VDD.n567 GND 0.007295f
C1918 VDD.n568 GND 0.009064f
C1919 VDD.n569 GND 0.009064f
C1920 VDD.n570 GND 0.009064f
C1921 VDD.n571 GND 0.009064f
C1922 VDD.n572 GND 0.009064f
C1923 VDD.n573 GND 0.007295f
C1924 VDD.n574 GND 0.007295f
C1925 VDD.n575 GND 0.009064f
C1926 VDD.n576 GND 0.009064f
C1927 VDD.n577 GND 0.007295f
C1928 VDD.n578 GND 0.009064f
C1929 VDD.n579 GND 0.009064f
C1930 VDD.n580 GND 0.009064f
C1931 VDD.n581 GND 0.009064f
C1932 VDD.n582 GND 0.009064f
C1933 VDD.n583 GND 0.007295f
C1934 VDD.n584 GND 0.009064f
C1935 VDD.n585 GND 0.007295f
C1936 VDD.n586 GND 0.00383f
C1937 VDD.n587 GND 0.009064f
C1938 VDD.n588 GND 0.009064f
C1939 VDD.n589 GND 0.007295f
C1940 VDD.n590 GND 0.009064f
C1941 VDD.n591 GND 0.007295f
C1942 VDD.n592 GND 0.009064f
C1943 VDD.n593 GND 0.007295f
C1944 VDD.n594 GND 0.009064f
C1945 VDD.n595 GND 0.007295f
C1946 VDD.n596 GND 0.009064f
C1947 VDD.n597 GND 0.007295f
C1948 VDD.n598 GND 0.009064f
C1949 VDD.n599 GND 0.007295f
C1950 VDD.n600 GND 0.009064f
C1951 VDD.n601 GND 0.009064f
C1952 VDD.n602 GND 0.765903f
C1953 VDD.t119 GND 0.384876f
C1954 VDD.n603 GND 0.009064f
C1955 VDD.n604 GND 0.007295f
C1956 VDD.n605 GND 0.009064f
C1957 VDD.n606 GND 0.007295f
C1958 VDD.n607 GND 0.009064f
C1959 VDD.n608 GND 0.769751f
C1960 VDD.n609 GND 0.009064f
C1961 VDD.n610 GND 0.007295f
C1962 VDD.n611 GND 0.009064f
C1963 VDD.n612 GND 0.007295f
C1964 VDD.n613 GND 0.009064f
C1965 VDD.t172 GND 0.384876f
C1966 VDD.n614 GND 0.009064f
C1967 VDD.n615 GND 0.007295f
C1968 VDD.n616 GND 0.009064f
C1969 VDD.n617 GND 0.007295f
C1970 VDD.n618 GND 0.009064f
C1971 VDD.n619 GND 0.504187f
C1972 VDD.n620 GND 0.009064f
C1973 VDD.n621 GND 0.007295f
C1974 VDD.n622 GND 0.009064f
C1975 VDD.n623 GND 0.007295f
C1976 VDD.n624 GND 0.009064f
C1977 VDD.n625 GND 0.758205f
C1978 VDD.t108 GND 0.384876f
C1979 VDD.n626 GND 0.009064f
C1980 VDD.n627 GND 0.007295f
C1981 VDD.n628 GND 0.009064f
C1982 VDD.n629 GND 0.007295f
C1983 VDD.n630 GND 0.009064f
C1984 VDD.n631 GND 0.769751f
C1985 VDD.n632 GND 0.009064f
C1986 VDD.n633 GND 0.007295f
C1987 VDD.n634 GND 0.009064f
C1988 VDD.n635 GND 0.007295f
C1989 VDD.n636 GND 0.009064f
C1990 VDD.t147 GND 0.384876f
C1991 VDD.n637 GND 0.009064f
C1992 VDD.n638 GND 0.007295f
C1993 VDD.n639 GND 0.009064f
C1994 VDD.n640 GND 0.007295f
C1995 VDD.n641 GND 0.009064f
C1996 VDD.n642 GND 0.769751f
C1997 VDD.n643 GND 0.009064f
C1998 VDD.n644 GND 0.007295f
C1999 VDD.n645 GND 0.009064f
C2000 VDD.n646 GND 0.007295f
C2001 VDD.n647 GND 0.009064f
C2002 VDD.n648 GND 0.565767f
C2003 VDD.n649 GND 0.009064f
C2004 VDD.n650 GND 0.007295f
C2005 VDD.n651 GND 0.020998f
C2006 VDD.n652 GND 0.006055f
C2007 VDD.n653 GND 0.020998f
C2008 VDD.n654 GND 1.05071f
C2009 VDD.n655 GND 0.020998f
C2010 VDD.n656 GND 0.006055f
C2011 VDD.n657 GND 0.009064f
C2012 VDD.t70 GND 0.111507f
C2013 VDD.t71 GND 0.123568f
C2014 VDD.t69 GND 0.30702f
C2015 VDD.n658 GND 0.203209f
C2016 VDD.n659 GND 0.158699f
C2017 VDD.n660 GND 0.011271f
C2018 VDD.n661 GND 0.009064f
C2019 VDD.n662 GND 4.50305f
C2020 VDD.n693 GND 0.009064f
C2021 VDD.n694 GND 0.009064f
C2022 VDD.n695 GND 0.021239f
C2023 VDD.n696 GND 0.009064f
C2024 VDD.n697 GND 0.009064f
C2025 VDD.n698 GND 0.009064f
C2026 VDD.n699 GND 0.009064f
C2027 VDD.n700 GND 0.009064f
C2028 VDD.n701 GND 0.009064f
C2029 VDD.n702 GND 0.007795f
C2030 VDD.n705 GND 0.005801f
C2031 VDD.n706 GND 0.009064f
C2032 VDD.n707 GND 0.009064f
C2033 VDD.n708 GND 0.009064f
C2034 VDD.n709 GND 0.009064f
C2035 VDD.n710 GND 0.009064f
C2036 VDD.n711 GND 0.009064f
C2037 VDD.n712 GND 0.006091f
C2038 VDD.n713 GND 0.009064f
C2039 VDD.n714 GND 0.009064f
C2040 VDD.n715 GND 0.009064f
C2041 VDD.n716 GND 0.009064f
C2042 VDD.n717 GND 0.009064f
C2043 VDD.n718 GND 0.009064f
C2044 VDD.n719 GND 0.009064f
C2045 VDD.n720 GND 0.009064f
C2046 VDD.n721 GND 0.009064f
C2047 VDD.n722 GND 0.009064f
C2048 VDD.n723 GND 0.009064f
C2049 VDD.n724 GND 0.009064f
C2050 VDD.n725 GND 0.009064f
C2051 VDD.n726 GND 0.009064f
C2052 VDD.n727 GND 0.009064f
C2053 VDD.n728 GND 0.009064f
C2054 VDD.n729 GND 0.009064f
C2055 VDD.n730 GND 0.009064f
C2056 VDD.n731 GND 0.009064f
C2057 VDD.n732 GND 0.007222f
C2058 VDD.t4 GND 0.111507f
C2059 VDD.t5 GND 0.123568f
C2060 VDD.t2 GND 0.30702f
C2061 VDD.n733 GND 0.203209f
C2062 VDD.n734 GND 0.158699f
C2063 VDD.n735 GND 0.009064f
C2064 VDD.n736 GND 0.009064f
C2065 VDD.n737 GND 0.009064f
C2066 VDD.n738 GND 0.009064f
C2067 VDD.n739 GND 0.009064f
C2068 VDD.n740 GND 0.009064f
C2069 VDD.n741 GND 0.009064f
C2070 VDD.n742 GND 0.005801f
C2071 VDD.n745 GND 0.004622f
C2072 VDD.n746 GND 0.006163f
C2073 VDD.n748 GND 0.006163f
C2074 VDD.n749 GND 0.006163f
C2075 VDD.n751 GND 0.006163f
C2076 VDD.n752 GND 0.004758f
C2077 VDD.n754 GND 0.006163f
C2078 VDD.t77 GND 0.0788f
C2079 VDD.t76 GND 0.089602f
C2080 VDD.t75 GND 0.235114f
C2081 VDD.n755 GND 0.156988f
C2082 VDD.n756 GND 0.126426f
C2083 VDD.n757 GND 0.008808f
C2084 VDD.n758 GND 0.014446f
C2085 VDD.n760 GND 0.006163f
C2086 VDD.n761 GND 0.523431f
C2087 VDD.n762 GND 0.013688f
C2088 VDD.n763 GND 0.013688f
C2089 VDD.n764 GND 0.006163f
C2090 VDD.n765 GND 0.014409f
C2091 VDD.n766 GND 0.006163f
C2092 VDD.n767 GND 0.006163f
C2093 VDD.n769 GND 0.006163f
C2094 VDD.n770 GND 0.006163f
C2095 VDD.n772 GND 0.006163f
C2096 VDD.n773 GND 0.006163f
C2097 VDD.n775 GND 0.006163f
C2098 VDD.n776 GND 0.006163f
C2099 VDD.n778 GND 0.006163f
C2100 VDD.n779 GND 0.006163f
C2101 VDD.n781 GND 0.006163f
C2102 VDD.n782 GND 0.004758f
C2103 VDD.n784 GND 0.006163f
C2104 VDD.t52 GND 0.0788f
C2105 VDD.t51 GND 0.089602f
C2106 VDD.t49 GND 0.235114f
C2107 VDD.n785 GND 0.156988f
C2108 VDD.n786 GND 0.126426f
C2109 VDD.n787 GND 0.008808f
C2110 VDD.n788 GND 0.006163f
C2111 VDD.n789 GND 0.006163f
C2112 VDD.n790 GND 0.288657f
C2113 VDD.n791 GND 0.006163f
C2114 VDD.n792 GND 0.006163f
C2115 VDD.n793 GND 0.006163f
C2116 VDD.n794 GND 0.006163f
C2117 VDD.n795 GND 0.006163f
C2118 VDD.n796 GND 0.438758f
C2119 VDD.n797 GND 0.006163f
C2120 VDD.n798 GND 0.006163f
C2121 VDD.t50 GND 0.261715f
C2122 VDD.n799 GND 0.006163f
C2123 VDD.n800 GND 0.006163f
C2124 VDD.t23 GND 0.089602f
C2125 VDD.t21 GND 0.235114f
C2126 VDD.t24 GND 0.089602f
C2127 VDD.n801 GND 0.284066f
C2128 VDD.n802 GND 0.006163f
C2129 VDD.n803 GND 0.006163f
C2130 VDD.n804 GND 0.523431f
C2131 VDD.n805 GND 0.006163f
C2132 VDD.n806 GND 0.006163f
C2133 VDD.t22 GND 0.261715f
C2134 VDD.n807 GND 0.006163f
C2135 VDD.n808 GND 0.006163f
C2136 VDD.n809 GND 0.006163f
C2137 VDD.n810 GND 0.523431f
C2138 VDD.n811 GND 0.006163f
C2139 VDD.n812 GND 0.006163f
C2140 VDD.n813 GND 0.006163f
C2141 VDD.n814 GND 0.006163f
C2142 VDD.n815 GND 0.006163f
C2143 VDD.t211 GND 0.261715f
C2144 VDD.n816 GND 0.006163f
C2145 VDD.n817 GND 0.006163f
C2146 VDD.n818 GND 0.006163f
C2147 VDD.n819 GND 0.006163f
C2148 VDD.n820 GND 0.006163f
C2149 VDD.t195 GND 0.261715f
C2150 VDD.n821 GND 0.006163f
C2151 VDD.n822 GND 0.006163f
C2152 VDD.n823 GND 0.4657f
C2153 VDD.n824 GND 0.006163f
C2154 VDD.n825 GND 0.006163f
C2155 VDD.n826 GND 0.006163f
C2156 VDD.t91 GND 0.261715f
C2157 VDD.n827 GND 0.006163f
C2158 VDD.n828 GND 0.006163f
C2159 VDD.n829 GND 0.315598f
C2160 VDD.n830 GND 0.006163f
C2161 VDD.n831 GND 0.006163f
C2162 VDD.n832 GND 0.006163f
C2163 VDD.t84 GND 0.261715f
C2164 VDD.n833 GND 0.006163f
C2165 VDD.n834 GND 0.006163f
C2166 VDD.n835 GND 0.488792f
C2167 VDD.n836 GND 0.006163f
C2168 VDD.n837 GND 0.006163f
C2169 VDD.n838 GND 0.006163f
C2170 VDD.t192 GND 0.261715f
C2171 VDD.n839 GND 0.006163f
C2172 VDD.n840 GND 0.006163f
C2173 VDD.n841 GND 0.338691f
C2174 VDD.n842 GND 0.006163f
C2175 VDD.n843 GND 0.006163f
C2176 VDD.n844 GND 0.006163f
C2177 VDD.t193 GND 0.261715f
C2178 VDD.n845 GND 0.006163f
C2179 VDD.n846 GND 0.006163f
C2180 VDD.n847 GND 0.511885f
C2181 VDD.n848 GND 0.006163f
C2182 VDD.n849 GND 0.006163f
C2183 VDD.n850 GND 0.006163f
C2184 VDD.n851 GND 0.523431f
C2185 VDD.n852 GND 0.006163f
C2186 VDD.n853 GND 0.006163f
C2187 VDD.t82 GND 0.261715f
C2188 VDD.n854 GND 0.006163f
C2189 VDD.n855 GND 0.006163f
C2190 VDD.n856 GND 0.006163f
C2191 VDD.t212 GND 0.261715f
C2192 VDD.n857 GND 0.006163f
C2193 VDD.n858 GND 0.006163f
C2194 VDD.n859 GND 0.006163f
C2195 VDD.n860 GND 0.006163f
C2196 VDD.n861 GND 0.006163f
C2197 VDD.n862 GND 0.523431f
C2198 VDD.n863 GND 0.006163f
C2199 VDD.n864 GND 0.006163f
C2200 VDD.t78 GND 0.261715f
C2201 VDD.n865 GND 0.006163f
C2202 VDD.n866 GND 0.006163f
C2203 VDD.n867 GND 0.006163f
C2204 VDD.n868 GND 0.4657f
C2205 VDD.n869 GND 0.006163f
C2206 VDD.n870 GND 0.006163f
C2207 VDD.n871 GND 0.006163f
C2208 VDD.n872 GND 0.006163f
C2209 VDD.n873 GND 0.006163f
C2210 VDD.t214 GND 0.261715f
C2211 VDD.n874 GND 0.006163f
C2212 VDD.n875 GND 0.006163f
C2213 VDD.t83 GND 0.261715f
C2214 VDD.n876 GND 0.006163f
C2215 VDD.n877 GND 0.006163f
C2216 VDD.n878 GND 0.006163f
C2217 VDD.n879 GND 0.523431f
C2218 VDD.n880 GND 0.006163f
C2219 VDD.n881 GND 0.006163f
C2220 VDD.n882 GND 0.377178f
C2221 VDD.n883 GND 0.006163f
C2222 VDD.n884 GND 0.006163f
C2223 VDD.n885 GND 0.006163f
C2224 VDD.t80 GND 0.261715f
C2225 VDD.n886 GND 0.006163f
C2226 VDD.n887 GND 0.006163f
C2227 VDD.n888 GND 0.006163f
C2228 VDD.n889 GND 0.006163f
C2229 VDD.n890 GND 0.006163f
C2230 VDD.t60 GND 0.261715f
C2231 VDD.n891 GND 0.006163f
C2232 VDD.n892 GND 0.006163f
C2233 VDD.n893 GND 0.400271f
C2234 VDD.n894 GND 0.006163f
C2235 VDD.n895 GND 0.006163f
C2236 VDD.n896 GND 0.006163f
C2237 VDD.t86 GND 0.261715f
C2238 VDD.n897 GND 0.006163f
C2239 VDD.n898 GND 0.006163f
C2240 VDD.n899 GND 0.288657f
C2241 VDD.n900 GND 0.006163f
C2242 VDD.n901 GND 0.014409f
C2243 VDD.n902 GND 0.014409f
C2244 VDD.n903 GND 0.723566f
C2245 VDD.n929 GND 0.014409f
C2246 VDD.n930 GND 0.013688f
C2247 VDD.n931 GND 0.006163f
C2248 VDD.n932 GND 0.013688f
C2249 VDD.t32 GND 0.0788f
C2250 VDD.t31 GND 0.089602f
C2251 VDD.t29 GND 0.235114f
C2252 VDD.n933 GND 0.156988f
C2253 VDD.n934 GND 0.126426f
C2254 VDD.n935 GND 0.008808f
C2255 VDD.n936 GND 0.006163f
C2256 VDD.n937 GND 0.006163f
C2257 VDD.t88 GND 0.261715f
C2258 VDD.n938 GND 0.006163f
C2259 VDD.n939 GND 0.006163f
C2260 VDD.n940 GND 0.006163f
C2261 VDD.n941 GND 0.013688f
C2262 VDD.n942 GND 0.006163f
C2263 VDD.t74 GND 0.0788f
C2264 VDD.t73 GND 0.089602f
C2265 VDD.t72 GND 0.235114f
C2266 VDD.n943 GND 0.156988f
C2267 VDD.n944 GND 0.126426f
C2268 VDD.n945 GND 0.006163f
C2269 VDD.n946 GND 0.006163f
C2270 VDD.n947 GND 0.288657f
C2271 VDD.n948 GND 0.006163f
C2272 VDD.n949 GND 0.006163f
C2273 VDD.n950 GND 0.006163f
C2274 VDD.n951 GND 0.400271f
C2275 VDD.n952 GND 0.006163f
C2276 VDD.n953 GND 0.006163f
C2277 VDD.t30 GND 0.261715f
C2278 VDD.n954 GND 0.006163f
C2279 VDD.n955 GND 0.006163f
C2280 VDD.n956 GND 0.006163f
C2281 VDD.n957 GND 0.006163f
C2282 VDD.n958 GND 0.523431f
C2283 VDD.n959 GND 0.006163f
C2284 VDD.n960 GND 0.006163f
C2285 VDD.t93 GND 0.261715f
C2286 VDD.n961 GND 0.006163f
C2287 VDD.n962 GND 0.006163f
C2288 VDD.n963 GND 0.006163f
C2289 VDD.n964 GND 0.377178f
C2290 VDD.n965 GND 0.006163f
C2291 VDD.n966 GND 0.006163f
C2292 VDD.n967 GND 0.006163f
C2293 VDD.n968 GND 0.006163f
C2294 VDD.n969 GND 0.006163f
C2295 VDD.t90 GND 0.261715f
C2296 VDD.n970 GND 0.006163f
C2297 VDD.n971 GND 0.006163f
C2298 VDD.t0 GND 0.261715f
C2299 VDD.n972 GND 0.006163f
C2300 VDD.n973 GND 0.006163f
C2301 VDD.n974 GND 0.006163f
C2302 VDD.n975 GND 0.523431f
C2303 VDD.n976 GND 0.006163f
C2304 VDD.n977 GND 0.006163f
C2305 VDD.n978 GND 0.4657f
C2306 VDD.n979 GND 0.006163f
C2307 VDD.n980 GND 0.006163f
C2308 VDD.n981 GND 0.006163f
C2309 VDD.t210 GND 0.261715f
C2310 VDD.n982 GND 0.006163f
C2311 VDD.n983 GND 0.006163f
C2312 VDD.n984 GND 0.006163f
C2313 VDD.n985 GND 0.006163f
C2314 VDD.n986 GND 0.006163f
C2315 VDD.n987 GND 0.523431f
C2316 VDD.n988 GND 0.006163f
C2317 VDD.n989 GND 0.006163f
C2318 VDD.t204 GND 0.261715f
C2319 VDD.n990 GND 0.006163f
C2320 VDD.n991 GND 0.006163f
C2321 VDD.n992 GND 0.006163f
C2322 VDD.t79 GND 0.261715f
C2323 VDD.n993 GND 0.006163f
C2324 VDD.n994 GND 0.006163f
C2325 VDD.n995 GND 0.006163f
C2326 VDD.n996 GND 0.006163f
C2327 VDD.n997 GND 0.006163f
C2328 VDD.n998 GND 0.511885f
C2329 VDD.n999 GND 0.006163f
C2330 VDD.n1000 GND 0.006163f
C2331 VDD.t202 GND 0.261715f
C2332 VDD.n1001 GND 0.006163f
C2333 VDD.n1002 GND 0.006163f
C2334 VDD.n1003 GND 0.006163f
C2335 VDD.n1004 GND 0.338691f
C2336 VDD.n1005 GND 0.006163f
C2337 VDD.n1006 GND 0.006163f
C2338 VDD.t191 GND 0.261715f
C2339 VDD.n1007 GND 0.006163f
C2340 VDD.n1008 GND 0.006163f
C2341 VDD.n1009 GND 0.006163f
C2342 VDD.n1010 GND 0.488792f
C2343 VDD.n1011 GND 0.006163f
C2344 VDD.n1012 GND 0.006163f
C2345 VDD.t198 GND 0.261715f
C2346 VDD.n1013 GND 0.006163f
C2347 VDD.n1014 GND 0.006163f
C2348 VDD.n1015 GND 0.006163f
C2349 VDD.n1016 GND 0.315598f
C2350 VDD.n1017 GND 0.006163f
C2351 VDD.n1018 GND 0.006163f
C2352 VDD.t92 GND 0.261715f
C2353 VDD.n1019 GND 0.006163f
C2354 VDD.n1020 GND 0.006163f
C2355 VDD.n1021 GND 0.006163f
C2356 VDD.n1022 GND 0.4657f
C2357 VDD.n1023 GND 0.006163f
C2358 VDD.n1024 GND 0.006163f
C2359 VDD.t200 GND 0.261715f
C2360 VDD.n1025 GND 0.006163f
C2361 VDD.n1026 GND 0.006163f
C2362 VDD.n1027 GND 0.006163f
C2363 VDD.n1028 GND 0.523431f
C2364 VDD.n1029 GND 0.006163f
C2365 VDD.n1030 GND 0.006163f
C2366 VDD.t197 GND 0.261715f
C2367 VDD.n1031 GND 0.006163f
C2368 VDD.n1032 GND 0.006163f
C2369 VDD.n1033 GND 0.006163f
C2370 VDD.n1034 GND 0.523431f
C2371 VDD.n1035 GND 0.006163f
C2372 VDD.n1036 GND 0.006163f
C2373 VDD.n1037 GND 0.006163f
C2374 VDD.n1038 GND 0.006163f
C2375 VDD.n1039 GND 0.006163f
C2376 VDD.t46 GND 0.261715f
C2377 VDD.n1040 GND 0.006163f
C2378 VDD.n1041 GND 0.006163f
C2379 VDD.n1042 GND 0.006163f
C2380 VDD.t47 GND 0.089602f
C2381 VDD.t45 GND 0.235114f
C2382 VDD.t48 GND 0.089602f
C2383 VDD.n1043 GND 0.284066f
C2384 VDD.n1044 GND 0.006163f
C2385 VDD.n1045 GND 0.006163f
C2386 VDD.t7 GND 0.261715f
C2387 VDD.n1046 GND 0.006163f
C2388 VDD.n1047 GND 0.006163f
C2389 VDD.n1048 GND 0.438758f
C2390 VDD.n1049 GND 0.006163f
C2391 VDD.n1050 GND 0.006163f
C2392 VDD.n1051 GND 0.006163f
C2393 VDD.n1052 GND 0.523431f
C2394 VDD.n1053 GND 0.006163f
C2395 VDD.n1054 GND 0.006163f
C2396 VDD.n1055 GND 0.288657f
C2397 VDD.n1056 GND 0.006163f
C2398 VDD.n1057 GND 0.014409f
C2399 VDD.n1058 GND 0.014409f
C2400 VDD.n1059 GND 4.50305f
C2401 VDD.n1060 GND 0.013688f
C2402 VDD.n1061 GND 0.013688f
C2403 VDD.n1062 GND 0.014409f
C2404 VDD.n1063 GND 0.006163f
C2405 VDD.n1065 GND 0.006163f
C2406 VDD.n1066 GND 0.006163f
C2407 VDD.n1067 GND 0.006163f
C2408 VDD.n1068 GND 0.006163f
C2409 VDD.n1069 GND 0.012195f
C2410 VDD.n1071 GND 0.006163f
C2411 VDD.n1072 GND 0.006163f
C2412 VDD.n1073 GND 0.006163f
C2413 VDD.n1074 GND 0.006163f
C2414 VDD.t64 GND 0.0788f
C2415 VDD.t65 GND 0.089602f
C2416 VDD.t63 GND 0.235114f
C2417 VDD.n1075 GND 0.156988f
C2418 VDD.n1076 GND 0.126426f
C2419 VDD.n1077 GND 0.008808f
C2420 VDD.n1079 GND 0.006163f
C2421 VDD.n1080 GND 0.006163f
C2422 VDD.n1081 GND 0.006163f
C2423 VDD.t8 GND 0.0788f
C2424 VDD.t9 GND 0.089602f
C2425 VDD.t6 GND 0.235114f
C2426 VDD.n1082 GND 0.156988f
C2427 VDD.n1083 GND 0.126426f
C2428 VDD.n1084 GND 0.006163f
C2429 VDD.n1085 GND 0.006163f
C2430 VDD.n1086 GND 0.006163f
C2431 VDD.n1087 GND 0.006163f
C2432 VDD.n1088 GND 0.005801f
C2433 VDD.n1091 GND 0.009064f
C2434 VDD.n1092 GND 0.007295f
C2435 VDD.n1093 GND 0.009064f
C2436 VDD.n1094 GND 0.009064f
C2437 VDD.n1095 GND 0.009064f
C2438 VDD.n1096 GND 0.007295f
C2439 VDD.n1097 GND 0.009064f
C2440 VDD.n1098 GND 0.009064f
C2441 VDD.n1099 GND 0.009064f
C2442 VDD.n1100 GND 0.009064f
C2443 VDD.t55 GND 0.111507f
C2444 VDD.t54 GND 0.123568f
C2445 VDD.t53 GND 0.30702f
C2446 VDD.n1101 GND 0.203209f
C2447 VDD.n1102 GND 0.158699f
C2448 VDD.n1103 GND 0.011271f
C2449 VDD.n1104 GND 0.020998f
C2450 VDD.n1106 GND 0.009064f
C2451 VDD.n1107 GND 0.006055f
C2452 VDD.n1108 GND 0.58886f
C2453 VDD.n1110 GND 0.009064f
C2454 VDD.n1113 GND 4.70703f
C2455 VDD.n1114 GND 0.009064f
C2456 VDD.n1115 GND 0.021239f
C2457 VDD.n1116 GND 0.007295f
C2458 VDD.n1117 GND 0.009064f
C2459 VDD.n1118 GND 0.007295f
C2460 VDD.n1119 GND 0.009064f
C2461 VDD.n1120 GND 0.769751f
C2462 VDD.n1121 GND 0.009064f
C2463 VDD.n1122 GND 0.007295f
C2464 VDD.n1123 GND 0.007295f
C2465 VDD.n1124 GND 0.009064f
C2466 VDD.n1125 GND 0.007295f
C2467 VDD.n1126 GND 0.009064f
C2468 VDD.n1127 GND 0.769751f
C2469 VDD.n1128 GND 0.009064f
C2470 VDD.n1129 GND 0.007295f
C2471 VDD.n1130 GND 0.009064f
C2472 VDD.n1131 GND 0.007295f
C2473 VDD.n1132 GND 0.009064f
C2474 VDD.t152 GND 0.384876f
C2475 VDD.n1133 GND 0.009064f
C2476 VDD.n1134 GND 0.007295f
C2477 VDD.n1135 GND 0.009064f
C2478 VDD.n1136 GND 0.007295f
C2479 VDD.n1137 GND 0.009064f
C2480 VDD.n1138 GND 0.396422f
C2481 VDD.n1139 GND 0.627347f
C2482 VDD.n1140 GND 0.009064f
C2483 VDD.n1141 GND 0.007295f
C2484 VDD.n1142 GND 0.009064f
C2485 VDD.n1143 GND 0.007295f
C2486 VDD.n1144 GND 0.009064f
C2487 VDD.n1145 GND 0.65044f
C2488 VDD.n1146 GND 0.009064f
C2489 VDD.n1147 GND 0.007295f
C2490 VDD.n1148 GND 0.009064f
C2491 VDD.n1149 GND 0.007295f
C2492 VDD.n1150 GND 0.009064f
C2493 VDD.n1151 GND 0.769751f
C2494 VDD.t124 GND 0.384876f
C2495 VDD.n1152 GND 0.009064f
C2496 VDD.n1153 GND 0.007295f
C2497 VDD.n1154 GND 0.009064f
C2498 VDD.n1155 GND 0.007295f
C2499 VDD.n1156 GND 0.009064f
C2500 VDD.t105 GND 0.384876f
C2501 VDD.n1157 GND 0.009064f
C2502 VDD.n1158 GND 0.007295f
C2503 VDD.n1159 GND 0.009064f
C2504 VDD.n1160 GND 0.007295f
C2505 VDD.n1161 GND 0.009064f
C2506 VDD.n1162 GND 0.388724f
C2507 VDD.n1163 GND 0.635045f
C2508 VDD.n1164 GND 0.009064f
C2509 VDD.n1165 GND 0.007295f
C2510 VDD.n1166 GND 0.009064f
C2511 VDD.n1167 GND 0.007295f
C2512 VDD.n1168 GND 0.009064f
C2513 VDD.n1169 GND 0.642742f
C2514 VDD.n1170 GND 0.009064f
C2515 VDD.n1171 GND 0.007295f
C2516 VDD.n1172 GND 0.009064f
C2517 VDD.n1173 GND 0.007295f
C2518 VDD.n1174 GND 0.009064f
C2519 VDD.n1175 GND 0.769751f
C2520 VDD.t143 GND 0.384876f
C2521 VDD.n1176 GND 0.009064f
C2522 VDD.n1177 GND 0.007295f
C2523 VDD.n1178 GND 0.009064f
C2524 VDD.n1179 GND 0.007295f
C2525 VDD.n1180 GND 0.009064f
C2526 VDD.t103 GND 0.384876f
C2527 VDD.n1181 GND 0.009064f
C2528 VDD.n1182 GND 0.007295f
C2529 VDD.n1183 GND 0.009064f
C2530 VDD.n1184 GND 0.007295f
C2531 VDD.n1185 GND 0.009064f
C2532 VDD.t117 GND 0.384876f
C2533 VDD.n1186 GND 0.642742f
C2534 VDD.n1187 GND 0.009064f
C2535 VDD.n1188 GND 0.007295f
C2536 VDD.n1189 GND 0.009064f
C2537 VDD.n1190 GND 0.007295f
C2538 VDD.n1191 GND 0.009064f
C2539 VDD.n1192 GND 0.635045f
C2540 VDD.n1193 GND 0.009064f
C2541 VDD.n1194 GND 0.007295f
C2542 VDD.n1195 GND 0.009064f
C2543 VDD.n1196 GND 0.007295f
C2544 VDD.n1197 GND 0.009064f
C2545 VDD.n1198 GND 0.769751f
C2546 VDD.t162 GND 0.384876f
C2547 VDD.n1199 GND 0.009064f
C2548 VDD.n1200 GND 0.007295f
C2549 VDD.n1201 GND 0.009064f
C2550 VDD.n1202 GND 0.007295f
C2551 VDD.n1203 GND 0.009064f
C2552 VDD.t115 GND 0.384876f
C2553 VDD.n1204 GND 0.009064f
C2554 VDD.n1205 GND 0.007295f
C2555 VDD.n1206 GND 0.009064f
C2556 VDD.n1207 GND 0.007295f
C2557 VDD.n1208 GND 0.009064f
C2558 VDD.t131 GND 0.384876f
C2559 VDD.n1209 GND 0.65044f
C2560 VDD.n1210 GND 0.009064f
C2561 VDD.n1211 GND 0.007295f
C2562 VDD.n1212 GND 0.009064f
C2563 VDD.n1213 GND 0.007295f
C2564 VDD.n1214 GND 0.009064f
C2565 VDD.n1215 GND 0.627347f
C2566 VDD.n1216 GND 0.009064f
C2567 VDD.n1217 GND 0.007295f
C2568 VDD.n1218 GND 0.009064f
C2569 VDD.n1219 GND 0.007295f
C2570 VDD.n1220 GND 0.009064f
C2571 VDD.n1221 GND 0.769751f
C2572 VDD.t101 GND 0.384876f
C2573 VDD.n1222 GND 0.009064f
C2574 VDD.n1223 GND 0.007295f
C2575 VDD.n1224 GND 0.009064f
C2576 VDD.n1225 GND 0.007295f
C2577 VDD.n1226 GND 0.009064f
C2578 VDD.n1227 GND 0.769751f
C2579 VDD.n1228 GND 0.009064f
C2580 VDD.n1229 GND 0.007295f
C2581 VDD.n1230 GND 0.009064f
C2582 VDD.n1231 GND 0.007295f
C2583 VDD.n1232 GND 0.009064f
C2584 VDD.t14 GND 0.384876f
C2585 VDD.n1233 GND 0.009064f
C2586 VDD.n1234 GND 0.007295f
C2587 VDD.n1235 GND 0.021239f
C2588 VDD.n1236 GND 0.021239f
C2589 VDD.n1237 GND 1.73579f
C2590 VDD.n1238 GND 0.021239f
C2591 VDD.n1239 GND 0.009064f
C2592 VDD.t15 GND 0.111507f
C2593 VDD.t16 GND 0.123568f
C2594 VDD.t13 GND 0.30702f
C2595 VDD.n1240 GND 0.203209f
C2596 VDD.n1241 GND 0.158699f
C2597 VDD.n1242 GND 0.007295f
C2598 VDD.n1243 GND 0.007295f
C2599 VDD.n1244 GND 0.009064f
C2600 VDD.n1245 GND 0.007295f
C2601 VDD.n1246 GND 0.009064f
C2602 VDD.n1247 GND 0.007295f
C2603 VDD.n1248 GND 0.009064f
C2604 VDD.n1249 GND 0.007295f
C2605 VDD.n1250 GND 0.009064f
C2606 VDD.n1251 GND 0.007295f
C2607 VDD.n1252 GND 0.009064f
C2608 VDD.n1253 GND 0.007295f
C2609 VDD.n1254 GND 0.009064f
C2610 VDD.n1255 GND 0.007295f
C2611 VDD.n1256 GND 0.009064f
C2612 VDD.n1257 GND 0.007295f
C2613 VDD.n1258 GND 0.009064f
C2614 VDD.n1259 GND 0.007295f
C2615 VDD.n1260 GND 0.009064f
C2616 VDD.n1261 GND 0.007222f
C2617 VDD.n1262 GND 0.009064f
C2618 VDD.n1264 GND 0.009064f
C2619 VDD.t43 GND 0.111507f
C2620 VDD.t44 GND 0.123568f
C2621 VDD.t42 GND 0.30702f
C2622 VDD.n1265 GND 0.203209f
C2623 VDD.n1266 GND 0.158699f
C2624 VDD.n1267 GND 0.007295f
C2625 VDD.n1268 GND 0.007295f
C2626 VDD.n1269 GND 0.009064f
C2627 VDD.n1270 GND 0.007295f
C2628 VDD.n1271 GND 0.009064f
C2629 VDD.n1272 GND 0.007295f
C2630 VDD.n1273 GND 0.009064f
C2631 VDD.n1274 GND 0.007295f
C2632 VDD.n1275 GND 0.009064f
C2633 VDD.n1276 GND 0.007295f
C2634 VDD.n1277 GND 0.009064f
C2635 VDD.n1278 GND 0.007295f
C2636 VDD.n1279 GND 0.009064f
C2637 VDD.n1280 GND 0.007295f
C2638 VDD.n1281 GND 0.009064f
C2639 VDD.n1282 GND 0.007295f
C2640 VDD.n1283 GND 0.009064f
C2641 VDD.n1284 GND 0.007295f
C2642 VDD.n1285 GND 0.009064f
C2643 VDD.n1286 GND 0.006091f
C2644 VDD.n1287 GND 0.009064f
C2645 VDD.n1289 GND 0.009064f
C2646 VDD.t57 GND 0.111507f
C2647 VDD.t58 GND 0.123568f
C2648 VDD.t56 GND 0.30702f
C2649 VDD.n1290 GND 0.203209f
C2650 VDD.n1291 GND 0.158699f
C2651 VDD.n1292 GND 0.007295f
C2652 VDD.n1293 GND 0.007295f
C2653 VDD.n1294 GND 0.009064f
C2654 VDD.n1295 GND 0.007295f
C2655 VDD.n1296 GND 0.009064f
C2656 VDD.n1297 GND 0.007295f
C2657 VDD.n1298 GND 0.009064f
C2658 VDD.n1299 GND 0.007295f
C2659 VDD.n1300 GND 0.009064f
C2660 VDD.n1301 GND 0.007295f
C2661 VDD.n1302 GND 0.009064f
C2662 VDD.n1303 GND 0.007295f
C2663 VDD.n1304 GND 0.009064f
C2664 VDD.n1305 GND 0.007295f
C2665 VDD.n1306 GND 0.009064f
C2666 VDD.n1307 GND 0.007295f
C2667 VDD.n1308 GND 0.006055f
C2668 VDD.n1310 GND 0.009064f
C2669 VDD.n1311 GND 0.007295f
C2670 VDD.n1312 GND 0.009064f
C2671 VDD.n1313 GND 0.009064f
C2672 VDD.n1314 GND 0.009064f
C2673 VDD.n1315 GND 0.007295f
C2674 VDD.n1316 GND 0.009064f
C2675 VDD.n1318 GND 0.009064f
C2676 VDD.n1320 GND 0.009064f
C2677 VDD.n1321 GND 0.007295f
C2678 VDD.n1322 GND 0.009064f
C2679 VDD.n1323 GND 0.009064f
C2680 VDD.n1324 GND 0.009064f
C2681 VDD.n1325 GND 0.007295f
C2682 VDD.n1326 GND 0.009064f
C2683 VDD.n1328 GND 0.009064f
C2684 VDD.n1330 GND 0.009064f
C2685 VDD.n1331 GND 0.007295f
C2686 VDD.n1332 GND 0.009064f
C2687 VDD.n1333 GND 0.009064f
C2688 VDD.n1334 GND 0.009064f
C2689 VDD.n1335 GND 0.007295f
C2690 VDD.n1336 GND 0.009064f
C2691 VDD.n1338 GND 0.009064f
C2692 VDD.n1340 GND 0.009064f
C2693 VDD.n1341 GND 0.007295f
C2694 VDD.n1342 GND 0.009064f
C2695 VDD.n1343 GND 0.009064f
C2696 VDD.n1344 GND 0.009064f
C2697 VDD.n1345 GND 0.009064f
C2698 VDD.n1346 GND 0.009064f
C2699 VDD.n1347 GND 0.007295f
C2700 VDD.n1348 GND 0.009064f
C2701 VDD.n1350 GND 0.009064f
C2702 VDD.n1351 GND 0.009064f
C2703 VDD.n1353 GND 0.009064f
C2704 VDD.n1354 GND 0.006091f
C2705 VDD.n1355 GND 0.014919f
C2706 VDD.n1356 GND 0.009064f
C2707 VDD.n1357 GND 0.009064f
C2708 VDD.n1358 GND 0.009064f
C2709 VDD.n1359 GND 0.007295f
C2710 VDD.n1360 GND 0.009064f
C2711 VDD.n1362 GND 0.009064f
C2712 VDD.n1364 GND 0.009064f
C2713 VDD.n1365 GND 0.007295f
C2714 VDD.n1366 GND 0.009064f
C2715 VDD.n1367 GND 0.009064f
C2716 VDD.n1368 GND 0.009064f
C2717 VDD.n1369 GND 0.007295f
C2718 VDD.n1370 GND 0.009064f
C2719 VDD.n1372 GND 0.009064f
C2720 VDD.n1374 GND 0.009064f
C2721 VDD.n1375 GND 0.007295f
C2722 VDD.n1376 GND 0.009064f
C2723 VDD.n1377 GND 0.009064f
C2724 VDD.n1378 GND 0.009064f
C2725 VDD.n1379 GND 0.007295f
C2726 VDD.n1380 GND 0.009064f
C2727 VDD.n1382 GND 0.009064f
C2728 VDD.n1384 GND 0.009064f
C2729 VDD.n1385 GND 0.007295f
C2730 VDD.n1386 GND 0.009064f
C2731 VDD.n1387 GND 0.009064f
C2732 VDD.n1388 GND 0.009064f
C2733 VDD.n1389 GND 0.007295f
C2734 VDD.n1390 GND 0.009064f
C2735 VDD.n1392 GND 0.009064f
C2736 VDD.n1394 GND 0.009064f
C2737 VDD.n1395 GND 0.007295f
C2738 VDD.n1396 GND 0.009064f
C2739 VDD.n1397 GND 0.009064f
C2740 VDD.n1398 GND 0.009064f
C2741 VDD.n1399 GND 0.009064f
C2742 VDD.n1400 GND 0.009064f
C2743 VDD.n1401 GND 0.007295f
C2744 VDD.n1402 GND 0.009064f
C2745 VDD.n1404 GND 0.009064f
C2746 VDD.n1405 GND 0.009064f
C2747 VDD.n1407 GND 0.009064f
C2748 VDD.n1408 GND 0.004961f
C2749 VDD.n1409 GND 0.014919f
C2750 VDD.n1410 GND 0.009064f
C2751 VDD.n1411 GND 0.009064f
C2752 VDD.n1412 GND 0.009064f
C2753 VDD.n1413 GND 0.007295f
C2754 VDD.n1414 GND 0.009064f
C2755 VDD.n1416 GND 0.009064f
C2756 VDD.n1418 GND 0.009064f
C2757 VDD.n1419 GND 0.007295f
C2758 VDD.n1420 GND 0.009064f
C2759 VDD.n1421 GND 0.009064f
C2760 VDD.n1422 GND 0.009064f
C2761 VDD.n1423 GND 0.007295f
C2762 VDD.n1424 GND 0.009064f
C2763 VDD.n1426 GND 0.009064f
C2764 VDD.n1428 GND 0.009064f
C2765 VDD.n1429 GND 0.007295f
C2766 VDD.n1430 GND 0.009064f
C2767 VDD.n1431 GND 0.009064f
C2768 VDD.n1432 GND 0.009064f
C2769 VDD.n1433 GND 0.007295f
C2770 VDD.n1434 GND 0.009064f
C2771 VDD.n1436 GND 0.009064f
C2772 VDD.n1438 GND 0.009064f
C2773 VDD.n1439 GND 0.007295f
C2774 VDD.n1440 GND 0.009064f
C2775 VDD.n1441 GND 0.009064f
C2776 VDD.n1442 GND 0.009064f
C2777 VDD.n1443 GND 0.007295f
C2778 VDD.n1444 GND 0.009064f
C2779 VDD.n1446 GND 0.009064f
C2780 VDD.n1448 GND 0.009064f
C2781 VDD.n1449 GND 0.007295f
C2782 VDD.n1450 GND 0.009064f
C2783 VDD.n1451 GND 0.009064f
C2784 VDD.n1452 GND 0.009064f
C2785 VDD.n1453 GND 0.009064f
C2786 VDD.n1454 GND 0.009064f
C2787 VDD.n1455 GND 0.007295f
C2788 VDD.n1456 GND 0.009064f
C2789 VDD.n1458 GND 0.009064f
C2790 VDD.n1459 GND 0.009064f
C2791 VDD.n1461 GND 0.009064f
C2792 VDD.n1462 GND 0.00383f
C2793 VDD.n1463 GND 0.011271f
C2794 VDD.n1464 GND 0.003465f
C2795 VDD.n1465 GND 0.021239f
C2796 VDD.n1466 GND 0.020998f
C2797 VDD.n1467 GND 0.006055f
C2798 VDD.n1468 GND 0.020998f
C2799 VDD.n1469 GND 0.58886f
C2800 VDD.n1470 GND 1.05071f
C2801 VDD.n1471 GND 0.020998f
C2802 VDD.n1472 GND 0.006055f
C2803 VDD.n1473 GND 0.020998f
C2804 VDD.n1474 GND 0.009064f
C2805 VDD.n1475 GND 0.009064f
C2806 VDD.n1476 GND 0.007295f
C2807 VDD.n1477 GND 0.009064f
C2808 VDD.n1478 GND 0.565767f
C2809 VDD.n1479 GND 0.009064f
C2810 VDD.n1480 GND 0.007295f
C2811 VDD.n1481 GND 0.009064f
C2812 VDD.n1482 GND 0.009064f
C2813 VDD.n1483 GND 0.009064f
C2814 VDD.n1484 GND 0.007295f
C2815 VDD.n1485 GND 0.009064f
C2816 VDD.n1486 GND 0.769751f
C2817 VDD.n1487 GND 0.009064f
C2818 VDD.n1488 GND 0.007295f
C2819 VDD.n1489 GND 0.009064f
C2820 VDD.n1490 GND 0.009064f
C2821 VDD.n1491 GND 0.009064f
C2822 VDD.n1492 GND 0.007295f
C2823 VDD.n1493 GND 0.009064f
C2824 VDD.n1494 GND 0.52728f
C2825 VDD.n1495 GND 0.009064f
C2826 VDD.n1496 GND 0.007295f
C2827 VDD.n1497 GND 0.009064f
C2828 VDD.n1498 GND 0.009064f
C2829 VDD.n1499 GND 0.009064f
C2830 VDD.n1500 GND 0.007295f
C2831 VDD.n1501 GND 0.009064f
C2832 VDD.n1502 GND 0.396422f
C2833 VDD.n1503 GND 0.769751f
C2834 VDD.n1504 GND 0.009064f
C2835 VDD.n1505 GND 0.007295f
C2836 VDD.n1506 GND 0.009064f
C2837 VDD.n1507 GND 0.009064f
C2838 VDD.n1508 GND 0.009064f
C2839 VDD.n1509 GND 0.007295f
C2840 VDD.n1510 GND 0.009064f
C2841 VDD.n1511 GND 0.758205f
C2842 VDD.n1512 GND 0.009064f
C2843 VDD.n1513 GND 0.007295f
C2844 VDD.n1514 GND 0.009064f
C2845 VDD.n1515 GND 0.009064f
C2846 VDD.n1516 GND 0.009064f
C2847 VDD.n1517 GND 0.007295f
C2848 VDD.n1518 GND 0.009064f
C2849 VDD.n1519 GND 0.504187f
C2850 VDD.n1520 GND 0.009064f
C2851 VDD.n1521 GND 0.007295f
C2852 VDD.n1522 GND 0.009064f
C2853 VDD.n1523 GND 0.009064f
C2854 VDD.n1524 GND 0.009064f
C2855 VDD.n1525 GND 0.007295f
C2856 VDD.n1526 GND 0.009064f
C2857 VDD.n1527 GND 0.519582f
C2858 VDD.n1528 GND 0.009064f
C2859 VDD.n1529 GND 0.007295f
C2860 VDD.n1530 GND 0.009064f
C2861 VDD.n1531 GND 0.009064f
C2862 VDD.n1532 GND 0.009064f
C2863 VDD.n1533 GND 0.007295f
C2864 VDD.n1534 GND 0.009064f
C2865 VDD.n1535 GND 0.388724f
C2866 VDD.n1536 GND 0.769751f
C2867 VDD.n1537 GND 0.009064f
C2868 VDD.n1538 GND 0.007295f
C2869 VDD.n1539 GND 0.009064f
C2870 VDD.n1540 GND 0.009064f
C2871 VDD.n1541 GND 0.009064f
C2872 VDD.n1542 GND 0.007295f
C2873 VDD.n1543 GND 0.009064f
C2874 VDD.n1544 GND 0.765903f
C2875 VDD.n1545 GND 0.009064f
C2876 VDD.n1546 GND 0.007295f
C2877 VDD.n1547 GND 0.009064f
C2878 VDD.n1548 GND 0.009064f
C2879 VDD.n1549 GND 0.009064f
C2880 VDD.n1550 GND 0.007295f
C2881 VDD.n1551 GND 0.009064f
C2882 VDD.n1552 GND 0.511885f
C2883 VDD.n1553 GND 0.009064f
C2884 VDD.n1554 GND 0.007295f
C2885 VDD.n1555 GND 0.009033f
C2886 VDD.n1556 GND 0.004974f
C2887 VDD.n1557 GND 0.004616f
C2888 VDD.n1558 GND 0.002553f
C2889 VDD.n1559 GND 0.005863f
C2890 VDD.n1560 GND 0.00248f
C2891 VDD.n1561 GND 0.002626f
C2892 VDD.n1562 GND 0.004616f
C2893 VDD.n1563 GND 0.00248f
C2894 VDD.n1564 GND 0.005863f
C2895 VDD.n1565 GND 0.002626f
C2896 VDD.n1566 GND 0.004616f
C2897 VDD.n1567 GND 0.00248f
C2898 VDD.n1568 GND 0.004397f
C2899 VDD.n1569 GND 0.00441f
C2900 VDD.t153 GND 0.012595f
C2901 VDD.n1570 GND 0.028025f
C2902 VDD.n1571 GND 0.145847f
C2903 VDD.n1572 GND 0.00248f
C2904 VDD.n1573 GND 0.002626f
C2905 VDD.n1574 GND 0.005863f
C2906 VDD.n1575 GND 0.005863f
C2907 VDD.n1576 GND 0.002626f
C2908 VDD.n1577 GND 0.00248f
C2909 VDD.n1578 GND 0.004616f
C2910 VDD.n1579 GND 0.004616f
C2911 VDD.n1580 GND 0.00248f
C2912 VDD.n1581 GND 0.002626f
C2913 VDD.n1582 GND 0.005863f
C2914 VDD.n1583 GND 0.005863f
C2915 VDD.n1584 GND 0.002626f
C2916 VDD.n1585 GND 0.00248f
C2917 VDD.n1586 GND 0.004616f
C2918 VDD.n1587 GND 0.004616f
C2919 VDD.n1588 GND 0.00248f
C2920 VDD.n1589 GND 0.002626f
C2921 VDD.n1590 GND 0.005863f
C2922 VDD.n1591 GND 0.005863f
C2923 VDD.n1592 GND 0.013861f
C2924 VDD.n1593 GND 0.002553f
C2925 VDD.n1594 GND 0.00248f
C2926 VDD.n1595 GND 0.011931f
C2927 VDD.n1596 GND 0.008658f
C2928 VDD.t141 GND 0.029181f
C2929 VDD.t164 GND 0.029181f
C2930 VDD.n1597 GND 0.20055f
C2931 VDD.n1598 GND 0.195838f
C2932 VDD.t171 GND 0.029181f
C2933 VDD.t106 GND 0.029181f
C2934 VDD.n1599 GND 0.20055f
C2935 VDD.n1600 GND 0.152908f
C2936 VDD.t137 GND 0.029181f
C2937 VDD.t150 GND 0.029181f
C2938 VDD.n1601 GND 0.20055f
C2939 VDD.n1602 GND 0.152908f
C2940 VDD.t163 GND 0.029181f
C2941 VDD.t118 GND 0.029181f
C2942 VDD.n1603 GND 0.20055f
C2943 VDD.n1604 GND 0.152908f
C2944 VDD.t132 GND 0.029181f
C2945 VDD.t142 GND 0.029181f
C2946 VDD.n1605 GND 0.20055f
C2947 VDD.n1606 GND 0.152908f
C2948 VDD.n1607 GND 0.004974f
C2949 VDD.n1608 GND 0.004616f
C2950 VDD.n1609 GND 0.002553f
C2951 VDD.n1610 GND 0.005863f
C2952 VDD.n1611 GND 0.00248f
C2953 VDD.n1612 GND 0.002626f
C2954 VDD.n1613 GND 0.004616f
C2955 VDD.n1614 GND 0.00248f
C2956 VDD.n1615 GND 0.005863f
C2957 VDD.n1616 GND 0.002626f
C2958 VDD.n1617 GND 0.004616f
C2959 VDD.n1618 GND 0.00248f
C2960 VDD.n1619 GND 0.004397f
C2961 VDD.n1620 GND 0.00441f
C2962 VDD.t102 GND 0.012595f
C2963 VDD.n1621 GND 0.028025f
C2964 VDD.n1622 GND 0.145847f
C2965 VDD.n1623 GND 0.00248f
C2966 VDD.n1624 GND 0.002626f
C2967 VDD.n1625 GND 0.005863f
C2968 VDD.n1626 GND 0.005863f
C2969 VDD.n1627 GND 0.002626f
C2970 VDD.n1628 GND 0.00248f
C2971 VDD.n1629 GND 0.004616f
C2972 VDD.n1630 GND 0.004616f
C2973 VDD.n1631 GND 0.00248f
C2974 VDD.n1632 GND 0.002626f
C2975 VDD.n1633 GND 0.005863f
C2976 VDD.n1634 GND 0.005863f
C2977 VDD.n1635 GND 0.002626f
C2978 VDD.n1636 GND 0.00248f
C2979 VDD.n1637 GND 0.004616f
C2980 VDD.n1638 GND 0.004616f
C2981 VDD.n1639 GND 0.00248f
C2982 VDD.n1640 GND 0.002626f
C2983 VDD.n1641 GND 0.005863f
C2984 VDD.n1642 GND 0.005863f
C2985 VDD.n1643 GND 0.013861f
C2986 VDD.n1644 GND 0.002553f
C2987 VDD.n1645 GND 0.00248f
C2988 VDD.n1646 GND 0.011931f
C2989 VDD.n1647 GND 0.008068f
C2990 VDD.n1648 GND 0.117377f
C2991 VDD.n1649 GND 0.004974f
C2992 VDD.n1650 GND 0.004616f
C2993 VDD.n1651 GND 0.002553f
C2994 VDD.n1652 GND 0.005863f
C2995 VDD.n1653 GND 0.00248f
C2996 VDD.n1654 GND 0.002626f
C2997 VDD.n1655 GND 0.004616f
C2998 VDD.n1656 GND 0.00248f
C2999 VDD.n1657 GND 0.005863f
C3000 VDD.n1658 GND 0.002626f
C3001 VDD.n1659 GND 0.004616f
C3002 VDD.n1660 GND 0.00248f
C3003 VDD.n1661 GND 0.004397f
C3004 VDD.n1662 GND 0.00441f
C3005 VDD.t174 GND 0.012595f
C3006 VDD.n1663 GND 0.028025f
C3007 VDD.n1664 GND 0.145847f
C3008 VDD.n1665 GND 0.00248f
C3009 VDD.n1666 GND 0.002626f
C3010 VDD.n1667 GND 0.005863f
C3011 VDD.n1668 GND 0.005863f
C3012 VDD.n1669 GND 0.002626f
C3013 VDD.n1670 GND 0.00248f
C3014 VDD.n1671 GND 0.004616f
C3015 VDD.n1672 GND 0.004616f
C3016 VDD.n1673 GND 0.00248f
C3017 VDD.n1674 GND 0.002626f
C3018 VDD.n1675 GND 0.005863f
C3019 VDD.n1676 GND 0.005863f
C3020 VDD.n1677 GND 0.002626f
C3021 VDD.n1678 GND 0.00248f
C3022 VDD.n1679 GND 0.004616f
C3023 VDD.n1680 GND 0.004616f
C3024 VDD.n1681 GND 0.00248f
C3025 VDD.n1682 GND 0.002626f
C3026 VDD.n1683 GND 0.005863f
C3027 VDD.n1684 GND 0.005863f
C3028 VDD.n1685 GND 0.013861f
C3029 VDD.n1686 GND 0.002553f
C3030 VDD.n1687 GND 0.00248f
C3031 VDD.n1688 GND 0.011931f
C3032 VDD.n1689 GND 0.008658f
C3033 VDD.t125 GND 0.029181f
C3034 VDD.t183 GND 0.029181f
C3035 VDD.n1690 GND 0.20055f
C3036 VDD.n1691 GND 0.195838f
C3037 VDD.t114 GND 0.029181f
C3038 VDD.t188 GND 0.029181f
C3039 VDD.n1692 GND 0.20055f
C3040 VDD.n1693 GND 0.152908f
C3041 VDD.t186 GND 0.029181f
C3042 VDD.t144 GND 0.029181f
C3043 VDD.n1694 GND 0.20055f
C3044 VDD.n1695 GND 0.152908f
C3045 VDD.t168 GND 0.029181f
C3046 VDD.t129 GND 0.029181f
C3047 VDD.n1696 GND 0.20055f
C3048 VDD.n1697 GND 0.152908f
C3049 VDD.t145 GND 0.029181f
C3050 VDD.t116 GND 0.029181f
C3051 VDD.n1698 GND 0.20055f
C3052 VDD.n1699 GND 0.152908f
C3053 VDD.n1700 GND 0.004974f
C3054 VDD.n1701 GND 0.004616f
C3055 VDD.n1702 GND 0.002553f
C3056 VDD.n1703 GND 0.005863f
C3057 VDD.n1704 GND 0.00248f
C3058 VDD.n1705 GND 0.002626f
C3059 VDD.n1706 GND 0.004616f
C3060 VDD.n1707 GND 0.00248f
C3061 VDD.n1708 GND 0.005863f
C3062 VDD.n1709 GND 0.002626f
C3063 VDD.n1710 GND 0.004616f
C3064 VDD.n1711 GND 0.00248f
C3065 VDD.n1712 GND 0.004397f
C3066 VDD.n1713 GND 0.00441f
C3067 VDD.t167 GND 0.012595f
C3068 VDD.n1714 GND 0.028025f
C3069 VDD.n1715 GND 0.145847f
C3070 VDD.n1716 GND 0.00248f
C3071 VDD.n1717 GND 0.002626f
C3072 VDD.n1718 GND 0.005863f
C3073 VDD.n1719 GND 0.005863f
C3074 VDD.n1720 GND 0.002626f
C3075 VDD.n1721 GND 0.00248f
C3076 VDD.n1722 GND 0.004616f
C3077 VDD.n1723 GND 0.004616f
C3078 VDD.n1724 GND 0.00248f
C3079 VDD.n1725 GND 0.002626f
C3080 VDD.n1726 GND 0.005863f
C3081 VDD.n1727 GND 0.005863f
C3082 VDD.n1728 GND 0.002626f
C3083 VDD.n1729 GND 0.00248f
C3084 VDD.n1730 GND 0.004616f
C3085 VDD.n1731 GND 0.004616f
C3086 VDD.n1732 GND 0.00248f
C3087 VDD.n1733 GND 0.002626f
C3088 VDD.n1734 GND 0.005863f
C3089 VDD.n1735 GND 0.005863f
C3090 VDD.n1736 GND 0.013861f
C3091 VDD.n1737 GND 0.002553f
C3092 VDD.n1738 GND 0.00248f
C3093 VDD.n1739 GND 0.011931f
C3094 VDD.n1740 GND 0.008068f
C3095 VDD.n1741 GND 0.06915f
C3096 VDD.n1742 GND 0.376011f
C3097 VDD.n1743 GND 0.004974f
C3098 VDD.n1744 GND 0.004616f
C3099 VDD.n1745 GND 0.002553f
C3100 VDD.n1746 GND 0.005863f
C3101 VDD.n1747 GND 0.00248f
C3102 VDD.n1748 GND 0.002626f
C3103 VDD.n1749 GND 0.004616f
C3104 VDD.n1750 GND 0.00248f
C3105 VDD.n1751 GND 0.005863f
C3106 VDD.n1752 GND 0.002626f
C3107 VDD.n1753 GND 0.004616f
C3108 VDD.n1754 GND 0.00248f
C3109 VDD.n1755 GND 0.004397f
C3110 VDD.n1756 GND 0.00441f
C3111 VDD.t185 GND 0.012595f
C3112 VDD.n1757 GND 0.028025f
C3113 VDD.n1758 GND 0.145847f
C3114 VDD.n1759 GND 0.00248f
C3115 VDD.n1760 GND 0.002626f
C3116 VDD.n1761 GND 0.005863f
C3117 VDD.n1762 GND 0.005863f
C3118 VDD.n1763 GND 0.002626f
C3119 VDD.n1764 GND 0.00248f
C3120 VDD.n1765 GND 0.004616f
C3121 VDD.n1766 GND 0.004616f
C3122 VDD.n1767 GND 0.00248f
C3123 VDD.n1768 GND 0.002626f
C3124 VDD.n1769 GND 0.005863f
C3125 VDD.n1770 GND 0.005863f
C3126 VDD.n1771 GND 0.002626f
C3127 VDD.n1772 GND 0.00248f
C3128 VDD.n1773 GND 0.004616f
C3129 VDD.n1774 GND 0.004616f
C3130 VDD.n1775 GND 0.00248f
C3131 VDD.n1776 GND 0.002626f
C3132 VDD.n1777 GND 0.005863f
C3133 VDD.n1778 GND 0.005863f
C3134 VDD.n1779 GND 0.013861f
C3135 VDD.n1780 GND 0.002553f
C3136 VDD.n1781 GND 0.00248f
C3137 VDD.n1782 GND 0.011931f
C3138 VDD.n1783 GND 0.008658f
C3139 VDD.t135 GND 0.029181f
C3140 VDD.t100 GND 0.029181f
C3141 VDD.n1784 GND 0.20055f
C3142 VDD.n1785 GND 0.195838f
C3143 VDD.t126 GND 0.029181f
C3144 VDD.t107 GND 0.029181f
C3145 VDD.n1786 GND 0.20055f
C3146 VDD.n1787 GND 0.152908f
C3147 VDD.t104 GND 0.029181f
C3148 VDD.t154 GND 0.029181f
C3149 VDD.n1788 GND 0.20055f
C3150 VDD.n1789 GND 0.152908f
C3151 VDD.t178 GND 0.029181f
C3152 VDD.t136 GND 0.029181f
C3153 VDD.n1790 GND 0.20055f
C3154 VDD.n1791 GND 0.152908f
C3155 VDD.t159 GND 0.029181f
C3156 VDD.t130 GND 0.029181f
C3157 VDD.n1792 GND 0.20055f
C3158 VDD.n1793 GND 0.152908f
C3159 VDD.n1794 GND 0.004974f
C3160 VDD.n1795 GND 0.004616f
C3161 VDD.n1796 GND 0.002553f
C3162 VDD.n1797 GND 0.005863f
C3163 VDD.n1798 GND 0.00248f
C3164 VDD.n1799 GND 0.002626f
C3165 VDD.n1800 GND 0.004616f
C3166 VDD.n1801 GND 0.00248f
C3167 VDD.n1802 GND 0.005863f
C3168 VDD.n1803 GND 0.002626f
C3169 VDD.n1804 GND 0.004616f
C3170 VDD.n1805 GND 0.00248f
C3171 VDD.n1806 GND 0.004397f
C3172 VDD.n1807 GND 0.00441f
C3173 VDD.t176 GND 0.012595f
C3174 VDD.n1808 GND 0.028025f
C3175 VDD.n1809 GND 0.145847f
C3176 VDD.n1810 GND 0.00248f
C3177 VDD.n1811 GND 0.002626f
C3178 VDD.n1812 GND 0.005863f
C3179 VDD.n1813 GND 0.005863f
C3180 VDD.n1814 GND 0.002626f
C3181 VDD.n1815 GND 0.00248f
C3182 VDD.n1816 GND 0.004616f
C3183 VDD.n1817 GND 0.004616f
C3184 VDD.n1818 GND 0.00248f
C3185 VDD.n1819 GND 0.002626f
C3186 VDD.n1820 GND 0.005863f
C3187 VDD.n1821 GND 0.005863f
C3188 VDD.n1822 GND 0.002626f
C3189 VDD.n1823 GND 0.00248f
C3190 VDD.n1824 GND 0.004616f
C3191 VDD.n1825 GND 0.004616f
C3192 VDD.n1826 GND 0.00248f
C3193 VDD.n1827 GND 0.002626f
C3194 VDD.n1828 GND 0.005863f
C3195 VDD.n1829 GND 0.005863f
C3196 VDD.n1830 GND 0.013861f
C3197 VDD.n1831 GND 0.002553f
C3198 VDD.n1832 GND 0.00248f
C3199 VDD.n1833 GND 0.011931f
C3200 VDD.n1834 GND 0.008068f
C3201 VDD.n1835 GND 0.06915f
C3202 VDD.n1836 GND 0.322101f
C3203 VDD.n1837 GND 1.9344f
C3204 VDD.n1838 GND 0.200692f
C3205 VDD.n1839 GND 0.009033f
C3206 VDD.n1840 GND 0.007295f
C3207 VDD.n1841 GND 0.009064f
C3208 VDD.n1842 GND 0.511885f
C3209 VDD.n1843 GND 0.009064f
C3210 VDD.n1844 GND 0.007295f
C3211 VDD.n1845 GND 0.009064f
C3212 VDD.n1846 GND 0.009064f
C3213 VDD.n1847 GND 0.009064f
C3214 VDD.n1848 GND 0.007295f
C3215 VDD.n1849 GND 0.009064f
C3216 VDD.t113 GND 0.384876f
C3217 VDD.n1850 GND 0.765903f
C3218 VDD.n1851 GND 0.009064f
C3219 VDD.n1852 GND 0.007295f
C3220 VDD.n1853 GND 0.009064f
C3221 VDD.n1854 GND 0.009064f
C3222 VDD.n1855 GND 0.009064f
C3223 VDD.n1856 GND 0.007295f
C3224 VDD.n1857 GND 0.009064f
C3225 VDD.n1858 GND 0.769751f
C3226 VDD.n1859 GND 0.009064f
C3227 VDD.n1860 GND 0.007295f
C3228 VDD.n1861 GND 0.009064f
C3229 VDD.n1862 GND 0.009064f
C3230 VDD.n1863 GND 0.009064f
C3231 VDD.n1864 GND 0.007295f
C3232 VDD.n1865 GND 0.009064f
C3233 VDD.n1866 GND 0.519582f
C3234 VDD.n1867 GND 0.009064f
C3235 VDD.n1868 GND 0.007295f
C3236 VDD.n1869 GND 0.009064f
C3237 VDD.n1870 GND 0.009064f
C3238 VDD.n1871 GND 0.009064f
C3239 VDD.n1872 GND 0.007295f
C3240 VDD.n1873 GND 0.009064f
C3241 VDD.n1874 GND 0.504187f
C3242 VDD.n1875 GND 0.009064f
C3243 VDD.n1876 GND 0.007295f
C3244 VDD.n1877 GND 0.009064f
C3245 VDD.n1878 GND 0.009064f
C3246 VDD.n1879 GND 0.009064f
C3247 VDD.n1880 GND 0.007295f
C3248 VDD.n1881 GND 0.009064f
C3249 VDD.t99 GND 0.384876f
C3250 VDD.n1882 GND 0.758205f
C3251 VDD.n1883 GND 0.009064f
C3252 VDD.n1884 GND 0.007295f
C3253 VDD.n1885 GND 0.009064f
C3254 VDD.n1886 GND 0.009064f
C3255 VDD.n1887 GND 0.009064f
C3256 VDD.n1888 GND 0.007295f
C3257 VDD.n1889 GND 0.009064f
C3258 VDD.n1890 GND 0.769751f
C3259 VDD.n1891 GND 0.009064f
C3260 VDD.n1892 GND 0.007295f
C3261 VDD.n1893 GND 0.009064f
C3262 VDD.n1894 GND 0.009064f
C3263 VDD.n1895 GND 0.009064f
C3264 VDD.n1896 GND 0.007295f
C3265 VDD.n1897 GND 0.009064f
C3266 VDD.n1898 GND 0.52728f
C3267 VDD.n1899 GND 0.009064f
C3268 VDD.n1900 GND 0.007295f
C3269 VDD.n1901 GND 0.009064f
C3270 VDD.n1902 GND 0.009064f
C3271 VDD.n1903 GND 0.009064f
C3272 VDD.n1904 GND 0.007295f
C3273 VDD.n1905 GND 0.009064f
C3274 VDD.n1906 GND 0.769751f
C3275 VDD.n1907 GND 0.009064f
C3276 VDD.n1908 GND 0.007295f
C3277 VDD.n1909 GND 0.009064f
C3278 VDD.n1910 GND 0.009064f
C3279 VDD.n1911 GND 0.009064f
C3280 VDD.n1912 GND 0.009064f
C3281 VDD.n1913 GND 0.007295f
C3282 VDD.n1914 GND 0.009064f
C3283 VDD.t26 GND 0.384876f
C3284 VDD.n1915 GND 0.565767f
C3285 VDD.n1916 GND 0.009064f
C3286 VDD.n1917 GND 0.007295f
C3287 VDD.n1918 GND 0.009064f
C3288 VDD.n1919 GND 0.009064f
C3289 VDD.n1920 GND 0.009064f
C3290 VDD.n1921 GND 0.007295f
C3291 VDD.n1923 GND 0.009064f
C3292 VDD.n1924 GND 0.009064f
C3293 VDD.n1925 GND 0.009064f
C3294 VDD.n1926 GND 0.009064f
C3295 VDD.n1927 GND 0.009064f
C3296 VDD.n1928 GND 0.007295f
C3297 VDD.n1930 GND 0.009064f
C3298 VDD.n1931 GND 0.009064f
C3299 VDD.n1932 GND 0.007795f
C3300 VDD.n1933 GND 0.007295f
C3301 VDD.n1934 GND 0.005801f
C3302 VDD.n1935 GND 0.007295f
C3303 VDD.n1936 GND 0.007295f
C3304 VDD.n1938 GND 0.009064f
C3305 VDD.n1939 GND 0.009064f
C3306 VDD.n1941 GND 0.009064f
C3307 VDD.n1942 GND 0.009064f
C3308 VDD.n1943 GND 0.009064f
C3309 VDD.n1944 GND 0.009064f
C3310 VDD.n1945 GND 0.007295f
C3311 VDD.n1947 GND 0.009064f
C3312 VDD.n1948 GND 0.009064f
C3313 VDD.n1949 GND 0.009064f
C3314 VDD.n1950 GND 0.009064f
C3315 VDD.n1951 GND 0.006091f
C3316 VDD.t38 GND 0.111507f
C3317 VDD.t37 GND 0.123568f
C3318 VDD.t36 GND 0.30702f
C3319 VDD.n1952 GND 0.203209f
C3320 VDD.n1953 GND 0.158699f
C3321 VDD.n1955 GND 0.009064f
C3322 VDD.n1956 GND 0.009064f
C3323 VDD.n1957 GND 0.007295f
C3324 VDD.n1958 GND 0.009064f
C3325 VDD.n1960 GND 0.009064f
C3326 VDD.n1961 GND 0.009064f
C3327 VDD.n1962 GND 0.009064f
C3328 VDD.n1963 GND 0.009064f
C3329 VDD.n1964 GND 0.007295f
C3330 VDD.n1966 GND 0.009064f
C3331 VDD.n1967 GND 0.009064f
C3332 VDD.n1968 GND 0.009064f
C3333 VDD.n1969 GND 0.009064f
C3334 VDD.n1970 GND 0.009064f
C3335 VDD.n1971 GND 0.007295f
C3336 VDD.n1973 GND 0.009064f
C3337 VDD.n1974 GND 0.009064f
C3338 VDD.n1975 GND 0.009064f
C3339 VDD.n1976 GND 0.009064f
C3340 VDD.n1977 GND 0.009064f
C3341 VDD.n1978 GND 0.007295f
C3342 VDD.n1980 GND 0.009064f
C3343 VDD.n1981 GND 0.009064f
C3344 VDD.n1982 GND 0.009064f
C3345 VDD.n1983 GND 0.009064f
C3346 VDD.n1984 GND 0.009064f
C3347 VDD.n1985 GND 0.007295f
C3348 VDD.n1987 GND 0.009064f
C3349 VDD.n1988 GND 0.009064f
C3350 VDD.n1989 GND 0.009064f
C3351 VDD.n1990 GND 0.009064f
C3352 VDD.n1991 GND 0.007222f
C3353 VDD.t28 GND 0.111507f
C3354 VDD.t27 GND 0.123568f
C3355 VDD.t25 GND 0.30702f
C3356 VDD.n1992 GND 0.203209f
C3357 VDD.n1993 GND 0.158699f
C3358 VDD.n1995 GND 0.009064f
C3359 VDD.n1996 GND 0.009064f
C3360 VDD.n1997 GND 0.007295f
C3361 VDD.n1998 GND 0.009064f
C3362 VDD.n2000 GND 0.009064f
C3363 VDD.n2001 GND 0.009064f
C3364 VDD.n2002 GND 0.009064f
C3365 VDD.n2003 GND 0.009064f
C3366 VDD.n2004 GND 0.007295f
C3367 VDD.n2006 GND 0.009064f
C3368 VDD.n2007 GND 0.009064f
C3369 VDD.n2008 GND 0.009064f
C3370 VDD.n2009 GND 0.009064f
C3371 VDD.n2010 GND 0.007295f
C3372 VDD.n2012 GND 0.009064f
C3373 VDD.n2014 GND 0.009064f
C3374 VDD.n2015 GND 0.007295f
C3375 VDD.n2016 GND 0.007295f
C3376 VDD.n2017 GND 0.009064f
C3377 VDD.n2019 GND 0.009064f
C3378 VDD.n2020 GND 0.009064f
C3379 VDD.n2021 GND 0.007295f
C3380 VDD.n2022 GND 0.007295f
C3381 VDD.n2023 GND 0.007295f
C3382 VDD.n2024 GND 0.009064f
C3383 VDD.n2026 GND 0.009064f
C3384 VDD.n2027 GND 0.009064f
C3385 VDD.n2028 GND 0.007295f
C3386 VDD.n2029 GND 0.007295f
C3387 VDD.n2030 GND 0.007295f
C3388 VDD.n2031 GND 0.009064f
C3389 VDD.n2033 GND 0.009064f
C3390 VDD.n2034 GND 0.009064f
C3391 VDD.n2035 GND 0.007295f
C3392 VDD.n2036 GND 0.009064f
C3393 VDD.n2037 GND 0.009064f
C3394 VDD.n2038 GND 0.009064f
C3395 VDD.n2039 GND 0.014919f
C3396 VDD.n2040 GND 0.004961f
C3397 VDD.n2041 GND 0.007295f
C3398 VDD.n2042 GND 0.009064f
C3399 VDD.n2044 GND 0.009064f
C3400 VDD.n2045 GND 0.009064f
C3401 VDD.n2046 GND 0.007295f
C3402 VDD.n2047 GND 0.007295f
C3403 VDD.n2048 GND 0.007295f
C3404 VDD.n2049 GND 0.009064f
C3405 VDD.n2051 GND 0.009064f
C3406 VDD.n2052 GND 0.009064f
C3407 VDD.n2053 GND 0.007295f
C3408 VDD.n2054 GND 0.007295f
C3409 VDD.n2055 GND 0.007295f
C3410 VDD.n2056 GND 0.009064f
C3411 VDD.n2058 GND 0.009064f
C3412 VDD.n2059 GND 0.009064f
C3413 VDD.n2060 GND 0.007295f
C3414 VDD.n2061 GND 0.007295f
C3415 VDD.n2062 GND 0.007295f
C3416 VDD.n2063 GND 0.009064f
C3417 VDD.n2065 GND 0.009064f
C3418 VDD.n2066 GND 0.009064f
C3419 VDD.n2067 GND 0.007295f
C3420 VDD.n2068 GND 0.007295f
C3421 VDD.n2069 GND 0.007295f
C3422 VDD.n2070 GND 0.009064f
C3423 VDD.n2072 GND 0.009064f
C3424 VDD.n2073 GND 0.009064f
C3425 VDD.n2074 GND 0.007295f
C3426 VDD.n2075 GND 0.009064f
C3427 VDD.n2076 GND 0.009064f
C3428 VDD.n2077 GND 0.009064f
C3429 VDD.n2078 GND 0.014919f
C3430 VDD.n2079 GND 0.006091f
C3431 VDD.n2080 GND 0.007295f
C3432 VDD.n2081 GND 0.009064f
C3433 VDD.n2083 GND 0.009064f
C3434 VDD.n2084 GND 0.009064f
C3435 VDD.n2085 GND 0.007295f
C3436 VDD.n2086 GND 0.007295f
C3437 VDD.n2087 GND 0.007295f
C3438 VDD.n2088 GND 0.009064f
C3439 VDD.n2090 GND 0.009064f
C3440 VDD.n2091 GND 0.009064f
C3441 VDD.n2092 GND 0.007295f
C3442 VDD.n2094 GND 0.459657f
C3443 VDD.n2096 GND 0.007295f
C3444 VDD.n2097 GND 0.007295f
C3445 VDD.n2098 GND 0.009064f
C3446 VDD.n2100 GND 0.009064f
C3447 VDD.n2101 GND 0.009064f
C3448 VDD.n2102 GND 0.007295f
C3449 VDD.n2103 GND 0.007295f
C3450 VDD.n2104 GND 0.007295f
C3451 VDD.n2105 GND 0.009064f
C3452 VDD.n2107 GND 0.009064f
C3453 VDD.n2108 GND 0.009064f
C3454 VDD.n2109 GND 0.007295f
C3455 VDD.n2110 GND 0.006055f
C3456 VDD.n2111 GND 0.021239f
C3457 VDD.n2112 GND 0.020998f
C3458 VDD.n2113 GND 0.006055f
C3459 VDD.n2114 GND 0.020998f
C3460 VDD.n2115 GND 1.05071f
C3461 VDD.n2116 GND 0.020998f
C3462 VDD.n2117 GND 0.021239f
C3463 VDD.n2118 GND 0.003465f
C3464 VDD.n2119 GND 0.021239f
C3465 VDD.n2120 GND 0.009064f
C3466 VDD.n2121 GND 0.00383f
C3467 VDD.n2122 GND 0.007295f
C3468 VDD.n2123 GND 0.007295f
C3469 VDD.n2124 GND 0.009064f
C3470 VDD.n2125 GND 0.009064f
C3471 VDD.n2126 GND 0.009064f
C3472 VDD.n2127 GND 0.007295f
C3473 VDD.n2128 GND 0.007295f
C3474 VDD.n2129 GND 0.007295f
C3475 VDD.n2130 GND 0.007795f
C3476 VDD.n2131 GND 0.459657f
C3477 VDD.n2132 GND 0.012195f
C3478 VDD.n2133 GND 0.004622f
C3479 VDD.n2134 GND 0.006163f
C3480 VDD.n2135 GND 0.006163f
C3481 VDD.n2136 GND 0.006163f
C3482 VDD.n2137 GND 0.006163f
C3483 VDD.n2138 GND 0.006163f
C3484 VDD.n2140 GND 0.006163f
C3485 VDD.n2141 GND 0.006163f
C3486 VDD.n2142 GND 0.006163f
C3487 VDD.n2143 GND 0.006163f
C3488 VDD.n2144 GND 0.006163f
C3489 VDD.n2146 GND 0.006163f
C3490 VDD.n2148 GND 0.006163f
C3491 VDD.n2149 GND 0.006163f
C3492 VDD.n2150 GND 0.006163f
C3493 VDD.n2151 GND 0.006163f
C3494 VDD.n2152 GND 0.006163f
C3495 VDD.n2154 GND 0.006163f
C3496 VDD.n2156 GND 0.006163f
C3497 VDD.n2157 GND 0.006163f
C3498 VDD.n2158 GND 0.006163f
C3499 VDD.n2159 GND 0.006163f
C3500 VDD.n2160 GND 0.006163f
C3501 VDD.n2162 GND 0.006163f
C3502 VDD.n2164 GND 0.006163f
C3503 VDD.n2165 GND 0.004622f
C3504 VDD.n2166 GND 0.006163f
C3505 VDD.n2167 GND 0.006163f
C3506 VDD.n2168 GND 0.006163f
C3507 VDD.n2170 GND 0.006163f
C3508 VDD.n2172 GND 0.006163f
C3509 VDD.n2173 GND 0.006163f
C3510 VDD.n2174 GND 0.006163f
C3511 VDD.n2175 GND 0.006163f
C3512 VDD.n2176 GND 0.006163f
C3513 VDD.n2178 GND 0.006163f
C3514 VDD.n2180 GND 0.006163f
C3515 VDD.n2181 GND 0.006163f
C3516 VDD.n2182 GND 0.004758f
C3517 VDD.n2183 GND 0.008808f
C3518 VDD.n2184 GND 0.004487f
C3519 VDD.n2185 GND 0.006163f
C3520 VDD.n2187 GND 0.006163f
C3521 VDD.n2188 GND 0.014409f
C3522 VDD.n2189 GND 0.014409f
C3523 VDD.n2190 GND 0.013688f
C3524 VDD.n2191 GND 0.006163f
C3525 VDD.n2192 GND 0.006163f
C3526 VDD.n2193 GND 0.006163f
C3527 VDD.n2194 GND 0.006163f
C3528 VDD.n2195 GND 0.006163f
C3529 VDD.n2196 GND 0.006163f
C3530 VDD.n2197 GND 0.006163f
C3531 VDD.n2198 GND 0.006163f
C3532 VDD.n2199 GND 0.006163f
C3533 VDD.n2200 GND 0.006163f
C3534 VDD.n2201 GND 0.006163f
C3535 VDD.n2202 GND 0.006163f
C3536 VDD.n2203 GND 0.006163f
C3537 VDD.n2204 GND 0.006163f
C3538 VDD.n2205 GND 0.006163f
C3539 VDD.n2206 GND 0.006163f
C3540 VDD.n2207 GND 0.006163f
C3541 VDD.n2208 GND 0.006163f
C3542 VDD.n2209 GND 0.006163f
C3543 VDD.n2210 GND 0.006163f
C3544 VDD.n2211 GND 0.006163f
C3545 VDD.n2212 GND 0.006163f
C3546 VDD.n2213 GND 0.006163f
C3547 VDD.n2214 GND 0.006163f
C3548 VDD.n2215 GND 0.006163f
C3549 VDD.n2216 GND 0.006163f
C3550 VDD.n2217 GND 0.006163f
C3551 VDD.n2218 GND 0.006163f
C3552 VDD.n2219 GND 0.006163f
C3553 VDD.n2220 GND 0.006163f
C3554 VDD.n2221 GND 0.006163f
C3555 VDD.n2222 GND 0.006163f
C3556 VDD.n2223 GND 0.006163f
C3557 VDD.n2224 GND 0.006163f
C3558 VDD.n2225 GND 0.006163f
C3559 VDD.n2226 GND 0.006163f
C3560 VDD.n2227 GND 0.006163f
C3561 VDD.n2228 GND 0.006163f
C3562 VDD.n2229 GND 0.006163f
C3563 VDD.n2230 GND 0.006163f
C3564 VDD.n2231 GND 0.006163f
C3565 VDD.n2232 GND 0.006163f
C3566 VDD.n2233 GND 0.006163f
C3567 VDD.n2234 GND 0.006163f
C3568 VDD.n2235 GND 0.006163f
C3569 VDD.n2236 GND 0.006163f
C3570 VDD.n2237 GND 0.006163f
C3571 VDD.n2238 GND 0.006163f
C3572 VDD.n2239 GND 0.006163f
C3573 VDD.n2240 GND 0.006163f
C3574 VDD.n2241 GND 0.006163f
C3575 VDD.n2242 GND 0.006163f
C3576 VDD.n2243 GND 0.006163f
C3577 VDD.n2244 GND 0.006163f
C3578 VDD.n2245 GND 0.006163f
C3579 VDD.n2246 GND 0.006163f
C3580 VDD.n2247 GND 0.006163f
C3581 VDD.n2248 GND 0.006163f
C3582 VDD.n2249 GND 0.006163f
C3583 VDD.n2250 GND 0.006163f
C3584 VDD.n2251 GND 0.006163f
C3585 VDD.n2252 GND 0.006163f
C3586 VDD.n2253 GND 0.006163f
C3587 VDD.n2254 GND 0.006163f
C3588 VDD.n2255 GND 0.006163f
C3589 VDD.n2256 GND 0.006163f
C3590 VDD.n2257 GND 0.006163f
C3591 VDD.n2258 GND 0.006163f
C3592 VDD.n2259 GND 0.006163f
C3593 VDD.n2260 GND 0.006163f
C3594 VDD.n2261 GND 0.350237f
C3595 VDD.n2262 GND 0.006163f
C3596 VDD.n2263 GND 0.006163f
C3597 VDD.n2264 GND 0.006163f
C3598 VDD.n2265 GND 0.006163f
C3599 VDD.n2266 GND 0.006163f
C3600 VDD.n2267 GND 0.006163f
C3601 VDD.n2268 GND 0.006163f
C3602 VDD.n2269 GND 0.006163f
C3603 VDD.n2270 GND 0.350237f
C3604 VDD.n2271 GND 0.006163f
C3605 VDD.n2272 GND 0.006163f
C3606 VDD.n2273 GND 0.006163f
C3607 VDD.n2274 GND 0.006163f
C3608 VDD.n2275 GND 0.006163f
C3609 VDD.n2276 GND 0.006163f
C3610 VDD.n2277 GND 0.006163f
C3611 VDD.n2278 GND 0.006163f
C3612 VDD.n2279 GND 0.006163f
C3613 VDD.n2280 GND 0.006163f
C3614 VDD.n2281 GND 0.006163f
C3615 VDD.n2282 GND 0.006163f
C3616 VDD.n2283 GND 0.006163f
C3617 VDD.n2284 GND 0.006163f
C3618 VDD.n2285 GND 0.006163f
C3619 VDD.n2286 GND 0.006163f
C3620 VDD.n2287 GND 0.006163f
C3621 VDD.n2288 GND 0.006163f
C3622 VDD.n2289 GND 0.006163f
C3623 VDD.n2290 GND 0.006163f
C3624 VDD.n2291 GND 0.006163f
C3625 VDD.n2292 GND 0.006163f
C3626 VDD.n2293 GND 0.006163f
C3627 VDD.n2294 GND 0.006163f
C3628 VDD.n2295 GND 0.006163f
C3629 VDD.n2296 GND 0.006163f
C3630 VDD.n2297 GND 0.006163f
C3631 VDD.n2298 GND 0.006163f
C3632 VDD.n2299 GND 0.006163f
C3633 VDD.n2300 GND 0.006163f
C3634 VDD.n2301 GND 0.006163f
C3635 VDD.n2302 GND 0.006163f
C3636 VDD.n2303 GND 0.013688f
C3637 VDD.n2304 GND 0.014409f
C3638 VDD.n2305 GND 0.014409f
C3639 VDD.n2306 GND 0.006163f
C3640 VDD.n2307 GND 0.006163f
C3641 VDD.n2308 GND 0.004487f
C3642 VDD.n2309 GND 0.006163f
C3643 VDD.n2311 GND 0.006163f
C3644 VDD.n2312 GND 0.004758f
C3645 VDD.n2313 GND 0.006163f
C3646 VDD.n2314 GND 0.006163f
C3647 VDD.n2315 GND 0.006163f
C3648 VDD.n2317 GND 0.006163f
C3649 VDD.n2319 GND 0.006163f
C3650 VDD.n2320 GND 0.006163f
C3651 VDD.n2321 GND 0.006163f
C3652 VDD.n2322 GND 0.006163f
C3653 VDD.n2323 GND 0.006163f
C3654 VDD.n2325 GND 0.006163f
C3655 VDD.n2326 GND 0.006163f
C3656 VDD.n2327 GND 0.006163f
C3657 VDD.n2328 GND 0.004622f
C3658 VDD.n2329 GND 0.006163f
C3659 VDD.n2331 GND 0.006163f
C3660 VDD.n2332 GND 0.004622f
C3661 VDD.n2333 GND 0.006163f
C3662 VDD.n2334 GND 0.006163f
C3663 VDD.n2335 GND 0.006163f
C3664 VDD.n2337 GND 0.006163f
C3665 VDD.n2339 GND 0.006163f
C3666 VDD.n2340 GND 0.006163f
C3667 VDD.n2341 GND 0.006163f
C3668 VDD.n2342 GND 0.006163f
C3669 VDD.n2343 GND 0.006163f
C3670 VDD.n2345 GND 0.006163f
C3671 VDD.n2346 GND 0.006163f
C3672 VDD.n2347 GND 0.006163f
C3673 VDD.n2348 GND 0.006163f
C3674 VDD.n2349 GND 0.006163f
C3675 VDD.n2350 GND 0.006163f
C3676 VDD.n2352 GND 0.006163f
C3677 VDD.n2353 GND 0.006163f
C3678 VDD.n2354 GND 0.014409f
C3679 VDD.n2355 GND 0.013688f
C3680 VDD.n2356 GND 0.013688f
C3681 VDD.n2357 GND 0.723566f
C3682 VDD.n2358 GND 0.013688f
C3683 VDD.n2359 GND 0.013688f
C3684 VDD.n2360 GND 0.006163f
C3685 VDD.n2361 GND 0.006163f
C3686 VDD.n2362 GND 0.006163f
C3687 VDD.n2363 GND 0.523431f
C3688 VDD.n2364 GND 0.006163f
C3689 VDD.n2365 GND 0.006163f
C3690 VDD.n2366 GND 0.006163f
C3691 VDD.n2367 GND 0.006163f
C3692 VDD.n2368 GND 0.006163f
C3693 VDD.n2369 GND 0.49649f
C3694 VDD.n2370 GND 0.006163f
C3695 VDD.n2371 GND 0.006163f
C3696 VDD.n2372 GND 0.005166f
C3697 VDD.n2373 GND 0.017854f
C3698 VDD.n2374 GND 0.004079f
C3699 VDD.n2375 GND 0.006163f
C3700 VDD.n2376 GND 0.346388f
C3701 VDD.n2377 GND 0.006163f
C3702 VDD.n2378 GND 0.006163f
C3703 VDD.n2379 GND 0.006163f
C3704 VDD.n2380 GND 0.006163f
C3705 VDD.n2381 GND 0.006163f
C3706 VDD.n2382 GND 0.523431f
C3707 VDD.n2383 GND 0.006163f
C3708 VDD.n2384 GND 0.006163f
C3709 VDD.n2385 GND 0.006163f
C3710 VDD.n2386 GND 0.006163f
C3711 VDD.n2387 GND 0.006163f
C3712 VDD.n2388 GND 0.319447f
C3713 VDD.n2389 GND 0.006163f
C3714 VDD.n2390 GND 0.006163f
C3715 VDD.n2391 GND 0.006163f
C3716 VDD.n2392 GND 0.006163f
C3717 VDD.n2393 GND 0.006163f
C3718 VDD.n2394 GND 0.469548f
C3719 VDD.n2395 GND 0.006163f
C3720 VDD.n2396 GND 0.006163f
C3721 VDD.n2397 GND 0.006163f
C3722 VDD.n2398 GND 0.006163f
C3723 VDD.n2399 GND 0.006163f
C3724 VDD.n2400 GND 0.296354f
C3725 VDD.n2401 GND 0.006163f
C3726 VDD.n2402 GND 0.006163f
C3727 VDD.n2403 GND 0.006163f
C3728 VDD.n2404 GND 0.006163f
C3729 VDD.n2405 GND 0.006163f
C3730 VDD.n2406 GND 0.446456f
C3731 VDD.n2407 GND 0.006163f
C3732 VDD.n2408 GND 0.006163f
C3733 VDD.n2409 GND 0.006163f
C3734 VDD.n2410 GND 0.006163f
C3735 VDD.n2411 GND 0.006163f
C3736 VDD.n2412 GND 0.273262f
C3737 VDD.n2413 GND 0.006163f
C3738 VDD.n2414 GND 0.006163f
C3739 VDD.n2415 GND 0.006163f
C3740 VDD.n2416 GND 0.006163f
C3741 VDD.n2417 GND 0.006163f
C3742 VDD.n2418 GND 0.423363f
C3743 VDD.n2419 GND 0.006163f
C3744 VDD.n2420 GND 0.006163f
C3745 VDD.n2421 GND 0.006163f
C3746 VDD.n2422 GND 0.006163f
C3747 VDD.n2423 GND 0.006163f
C3748 VDD.n2424 GND 0.273262f
C3749 VDD.n2425 GND 0.006163f
C3750 VDD.n2426 GND 0.006163f
C3751 VDD.n2427 GND 0.006163f
C3752 VDD.n2428 GND 0.006163f
C3753 VDD.n2429 GND 0.006163f
C3754 VDD.n2430 GND 0.400271f
C3755 VDD.n2431 GND 0.006163f
C3756 VDD.n2432 GND 0.006163f
C3757 VDD.n2433 GND 0.006163f
C3758 VDD.n2434 GND 0.006163f
C3759 VDD.n2435 GND 0.006163f
C3760 VDD.n2436 GND 0.296354f
C3761 VDD.n2437 GND 0.006163f
C3762 VDD.n2438 GND 0.006163f
C3763 VDD.n2439 GND 0.006163f
C3764 VDD.n2440 GND 0.006163f
C3765 VDD.n2441 GND 0.006163f
C3766 VDD.n2442 GND 0.523431f
C3767 VDD.n2443 GND 0.006163f
C3768 VDD.n2444 GND 0.006163f
C3769 VDD.n2445 GND 0.006163f
C3770 VDD.n2446 GND 0.006163f
C3771 VDD.n2447 GND 0.006163f
C3772 VDD.n2448 GND 0.203984f
C3773 VDD.n2449 GND 0.006163f
C3774 VDD.n2450 GND 0.006163f
C3775 VDD.n2451 GND 0.006163f
C3776 VDD.n2452 GND 0.006163f
C3777 VDD.n2453 GND 0.006163f
C3778 VDD.n2454 GND 0.523431f
C3779 VDD.n2455 GND 0.006163f
C3780 VDD.n2456 GND 0.006163f
C3781 VDD.n2457 GND 0.006163f
C3782 VDD.n2458 GND 0.006163f
C3783 VDD.n2459 GND 0.006163f
C3784 VDD.n2460 GND 0.384876f
C3785 VDD.n2461 GND 0.006163f
C3786 VDD.n2462 GND 0.006163f
C3787 VDD.n2463 GND 0.006163f
C3788 VDD.n2464 GND 0.006163f
C3789 VDD.n2465 GND 0.006163f
C3790 VDD.n2466 GND 0.006163f
C3791 VDD.n2467 GND 0.49649f
C3792 VDD.n2468 GND 0.006163f
C3793 VDD.n2469 GND 0.006163f
C3794 VDD.n2470 GND 0.006163f
C3795 VDD.n2471 GND 0.006163f
C3796 VDD.n2472 GND 0.006163f
C3797 VDD.n2473 GND 0.006163f
C3798 VDD.n2474 GND 0.361783f
C3799 VDD.n2475 GND 0.006163f
C3800 VDD.n2476 GND 0.006163f
C3801 VDD.n2477 GND 0.006163f
C3802 VDD.n2478 GND 0.014446f
C3803 VDD.n2479 GND 0.013688f
C3804 VDD.n2480 GND 0.014409f
C3805 VDD.n2481 GND 0.013651f
C3806 VDD.n2482 GND 0.006163f
C3807 VDD.n2483 GND 0.006163f
C3808 VDD.n2484 GND 0.006163f
C3809 VDD.n2485 GND 0.004487f
C3810 VDD.n2486 GND 0.008808f
C3811 VDD.n2487 GND 0.004758f
C3812 VDD.n2488 GND 0.006163f
C3813 VDD.n2489 GND 0.006163f
C3814 VDD.n2490 GND 0.006163f
C3815 VDD.n2491 GND 0.006163f
C3816 VDD.n2492 GND 0.006163f
C3817 VDD.n2493 GND 0.006163f
C3818 VDD.n2494 GND 0.006163f
C3819 VDD.n2495 GND 0.006163f
C3820 VDD.n2496 GND 0.006163f
C3821 VDD.n2497 GND 0.006163f
C3822 VDD.n2498 GND 0.006163f
C3823 VDD.n2499 GND 0.006163f
C3824 VDD.n2500 GND 0.006163f
C3825 VDD.n2501 GND 0.006163f
C3826 VDD.n2502 GND 0.006163f
C3827 VDD.n2503 GND 0.006163f
C3828 VDD.n2504 GND 0.006163f
C3829 VDD.n2505 GND 0.006163f
C3830 VDD.n2506 GND 0.006163f
C3831 VDD.n2507 GND 0.006163f
C3832 VDD.n2508 GND 0.006163f
C3833 VDD.n2509 GND 0.006163f
C3834 VDD.n2510 GND 0.006163f
C3835 VDD.n2511 GND 0.006163f
C3836 VDD.n2512 GND 0.006163f
C3837 VDD.n2513 GND 0.006163f
C3838 VDD.n2514 GND 0.006163f
C3839 VDD.n2515 GND 0.006163f
C3840 VDD.n2516 GND 0.006163f
C3841 VDD.n2517 GND 0.006163f
C3842 VDD.n2518 GND 0.006163f
C3843 VDD.n2519 GND 0.006163f
C3844 VDD.n2520 GND 0.006163f
C3845 VDD.n2521 GND 0.006163f
C3846 VDD.n2522 GND 0.006163f
C3847 VDD.n2523 GND 0.006163f
C3848 VDD.n2524 GND 0.006163f
C3849 VDD.n2525 GND 0.006163f
C3850 VDD.n2526 GND 0.006163f
C3851 VDD.n2527 GND 0.006163f
C3852 VDD.n2528 GND 0.006163f
C3853 VDD.n2529 GND 0.006163f
C3854 VDD.n2530 GND 0.006163f
C3855 VDD.n2531 GND 0.014409f
C3856 VDD.n2532 GND 0.014409f
C3857 VDD.n2533 GND 0.013688f
C3858 VDD.n2534 GND 0.006163f
C3859 VDD.n2535 GND 0.006163f
C3860 VDD.n2536 GND 0.423363f
C3861 VDD.n2537 GND 0.006163f
C3862 VDD.n2538 GND 0.013688f
C3863 VDD.n2539 GND 0.014446f
C3864 VDD.n2540 GND 0.013651f
C3865 VDD.n2541 GND 0.006163f
C3866 VDD.n2542 GND 0.006163f
C3867 VDD.n2543 GND 0.004487f
C3868 VDD.n2544 GND 0.006163f
C3869 VDD.n2545 GND 0.006163f
C3870 VDD.n2546 GND 0.004758f
C3871 VDD.n2547 GND 0.006163f
C3872 VDD.n2548 GND 0.006163f
C3873 VDD.n2549 GND 0.006163f
C3874 VDD.n2550 GND 0.006163f
C3875 VDD.n2551 GND 0.006163f
C3876 VDD.n2552 GND 0.006163f
C3877 VDD.n2553 GND 0.006163f
C3878 VDD.n2554 GND 0.006163f
C3879 VDD.n2555 GND 0.006163f
C3880 VDD.n2556 GND 0.006163f
C3881 VDD.n2557 GND 0.006163f
C3882 VDD.n2558 GND 0.006163f
C3883 VDD.n2559 GND 0.006163f
C3884 VDD.n2560 GND 0.006163f
C3885 VDD.n2561 GND 0.006163f
C3886 VDD.n2562 GND 0.006163f
C3887 VDD.n2563 GND 0.006163f
C3888 VDD.n2564 GND 0.006163f
C3889 VDD.n2565 GND 0.006163f
C3890 VDD.n2566 GND 0.006163f
C3891 VDD.n2567 GND 0.006163f
C3892 VDD.n2568 GND 0.006163f
C3893 VDD.n2569 GND 0.006163f
C3894 VDD.n2570 GND 0.006163f
C3895 VDD.n2571 GND 0.006163f
C3896 VDD.n2572 GND 0.006163f
C3897 VDD.n2573 GND 0.006163f
C3898 VDD.n2574 GND 0.006163f
C3899 VDD.n2575 GND 0.006163f
C3900 VDD.n2576 GND 0.006163f
C3901 VDD.n2577 GND 0.006163f
C3902 VDD.n2578 GND 0.006163f
C3903 VDD.n2579 GND 0.006163f
C3904 VDD.n2580 GND 0.006163f
C3905 VDD.n2581 GND 0.006163f
C3906 VDD.n2582 GND 0.006163f
C3907 VDD.n2583 GND 0.006163f
C3908 VDD.n2584 GND 0.006163f
C3909 VDD.n2585 GND 0.006163f
C3910 VDD.n2586 GND 0.006163f
C3911 VDD.n2587 GND 0.006163f
C3912 VDD.n2588 GND 0.014409f
C3913 VDD.n2589 GND 0.014409f
C3914 VDD.n2590 GND 0.600406f
C3915 VDD.t206 GND 2.65564f
C3916 VDD.t208 GND 2.65564f
C3917 VDD.n2591 GND 0.600406f
C3918 VDD.n2592 GND 0.013688f
C3919 VDD.n2593 GND 0.013688f
C3920 VDD.n2594 GND 0.423363f
C3921 VDD.n2595 GND 0.014409f
C3922 VDD.n2596 GND 0.006163f
C3923 VDD.n2597 GND 0.006163f
C3924 VDD.n2598 GND 0.006163f
C3925 VDD.n2599 GND 0.006163f
C3926 VDD.n2600 GND 0.006163f
C3927 VDD.n2601 GND 0.006163f
C3928 VDD.n2602 GND 0.006163f
C3929 VDD.n2603 GND 0.006163f
C3930 VDD.n2604 GND 0.006163f
C3931 VDD.n2605 GND 0.006163f
C3932 VDD.n2606 GND 0.004758f
C3933 VDD.n2607 GND 0.006163f
C3934 VDD.t61 GND 0.0788f
C3935 VDD.t62 GND 0.089602f
C3936 VDD.t59 GND 0.235114f
C3937 VDD.n2608 GND 0.156988f
C3938 VDD.n2609 GND 0.126426f
C3939 VDD.n2610 GND 0.008808f
C3940 VDD.n2611 GND 0.006163f
C3941 VDD.n2612 GND 0.006163f
C3942 VDD.n2613 GND 0.006163f
C3943 VDD.t67 GND 0.0788f
C3944 VDD.t68 GND 0.089602f
C3945 VDD.t66 GND 0.235114f
C3946 VDD.n2614 GND 0.156988f
C3947 VDD.n2615 GND 0.126426f
C3948 VDD.n2616 GND 0.006163f
C3949 VDD.n2617 GND 0.006163f
C3950 VDD.n2618 GND 0.006163f
C3951 VDD.n2619 GND 0.006163f
C3952 VDD.n2620 GND 0.006163f
C3953 VDD.n2621 GND 0.006163f
C3954 VDD.n2622 GND 0.006163f
C3955 VDD.n2623 GND 0.006163f
C3956 VDD.n2624 GND 0.006163f
C3957 VDD.n2625 GND 0.006163f
C3958 VDD.n2627 GND 0.006163f
C3959 VDD.n2628 GND 0.006163f
C3960 VDD.n2629 GND 0.006163f
C3961 VDD.n2630 GND 0.006163f
C3962 VDD.n2631 GND 0.006163f
C3963 VDD.n2633 GND 0.006163f
C3964 VDD.n2635 GND 0.006163f
C3965 VDD.n2636 GND 0.006163f
C3966 VDD.n2637 GND 0.006163f
C3967 VDD.n2638 GND 0.006163f
C3968 VDD.n2639 GND 0.006163f
C3969 VDD.n2641 GND 0.006163f
C3970 VDD.n2643 GND 0.006163f
C3971 VDD.n2644 GND 0.006163f
C3972 VDD.n2645 GND 0.006163f
C3973 VDD.n2646 GND 0.006163f
C3974 VDD.n2647 GND 0.006163f
C3975 VDD.n2649 GND 0.006163f
C3976 VDD.n2651 GND 0.006163f
C3977 VDD.n2652 GND 0.006163f
C3978 VDD.n2653 GND 0.006163f
C3979 VDD.n2654 GND 0.006163f
C3980 VDD.n2655 GND 0.006163f
C3981 VDD.n2657 GND 0.006163f
C3982 VDD.n2659 GND 0.006163f
C3983 VDD.n2660 GND 0.006163f
C3984 VDD.n2661 GND 0.006163f
C3985 VDD.n2662 GND 0.006163f
C3986 VDD.n2663 GND 0.006163f
C3987 VDD.n2665 GND 0.006163f
C3988 VDD.n2667 GND 0.006163f
C3989 VDD.n2668 GND 0.006163f
C3990 VDD.n2669 GND 0.004758f
C3991 VDD.n2670 GND 0.008808f
C3992 VDD.n2671 GND 0.004487f
C3993 VDD.n2672 GND 0.006163f
C3994 VDD.n2674 GND 0.006163f
C3995 VDD.n2675 GND 0.014409f
C3996 VDD.n2676 GND 0.014409f
C3997 VDD.n2677 GND 0.013688f
C3998 VDD.n2678 GND 0.006163f
C3999 VDD.n2679 GND 0.006163f
C4000 VDD.n2680 GND 0.006163f
C4001 VDD.n2681 GND 0.006163f
C4002 VDD.n2682 GND 0.006163f
C4003 VDD.n2683 GND 0.006163f
C4004 VDD.n2684 GND 0.006163f
C4005 VDD.n2685 GND 0.006163f
C4006 VDD.n2686 GND 0.006163f
C4007 VDD.n2687 GND 0.006163f
C4008 VDD.n2688 GND 0.006163f
C4009 VDD.n2689 GND 0.006163f
C4010 VDD.n2690 GND 0.006163f
C4011 VDD.n2691 GND 0.006163f
C4012 VDD.n2692 GND 0.006163f
C4013 VDD.n2693 GND 0.006163f
C4014 VDD.n2694 GND 0.006163f
C4015 VDD.n2695 GND 0.006163f
C4016 VDD.n2696 GND 0.006163f
C4017 VDD.n2697 GND 0.006163f
C4018 VDD.n2698 GND 0.006163f
C4019 VDD.n2699 GND 0.006163f
C4020 VDD.n2700 GND 0.006163f
C4021 VDD.n2701 GND 0.006163f
C4022 VDD.n2702 GND 0.006163f
C4023 VDD.n2703 GND 0.006163f
C4024 VDD.n2704 GND 0.006163f
C4025 VDD.n2705 GND 0.006163f
C4026 VDD.n2706 GND 0.006163f
C4027 VDD.n2707 GND 0.006163f
C4028 VDD.n2708 GND 0.006163f
C4029 VDD.n2709 GND 0.006163f
C4030 VDD.n2710 GND 0.006163f
C4031 VDD.n2711 GND 0.006163f
C4032 VDD.n2712 GND 0.006163f
C4033 VDD.n2713 GND 0.006163f
C4034 VDD.n2714 GND 0.006163f
C4035 VDD.n2715 GND 0.006163f
C4036 VDD.n2716 GND 0.006163f
C4037 VDD.n2717 GND 0.006163f
C4038 VDD.n2718 GND 0.006163f
C4039 VDD.n2719 GND 0.006163f
C4040 VDD.n2720 GND 0.006163f
C4041 VDD.n2721 GND 0.006163f
C4042 VDD.n2722 GND 0.006163f
C4043 VDD.n2723 GND 0.006163f
C4044 VDD.n2724 GND 0.006163f
C4045 VDD.n2725 GND 0.006163f
C4046 VDD.n2726 GND 0.006163f
C4047 VDD.n2727 GND 0.006163f
C4048 VDD.n2728 GND 0.006163f
C4049 VDD.n2729 GND 0.006163f
C4050 VDD.n2730 GND 0.006163f
C4051 VDD.n2731 GND 0.006163f
C4052 VDD.n2732 GND 0.006163f
C4053 VDD.n2733 GND 0.006163f
C4054 VDD.n2734 GND 0.006163f
C4055 VDD.n2735 GND 0.006163f
C4056 VDD.n2736 GND 0.006163f
C4057 VDD.n2737 GND 0.006163f
C4058 VDD.n2738 GND 0.006163f
C4059 VDD.n2739 GND 0.006163f
C4060 VDD.n2740 GND 0.006163f
C4061 VDD.n2741 GND 0.006163f
C4062 VDD.n2742 GND 0.006163f
C4063 VDD.n2743 GND 0.006163f
C4064 VDD.n2744 GND 0.006163f
C4065 VDD.n2745 GND 0.006163f
C4066 VDD.n2746 GND 0.006163f
C4067 VDD.n2747 GND 0.006163f
C4068 VDD.n2748 GND 0.006163f
C4069 VDD.n2749 GND 0.006163f
C4070 VDD.n2750 GND 0.006163f
C4071 VDD.n2751 GND 0.006163f
C4072 VDD.n2752 GND 0.006163f
C4073 VDD.n2753 GND 0.006163f
C4074 VDD.n2754 GND 0.006163f
C4075 VDD.n2755 GND 0.006163f
C4076 VDD.n2756 GND 0.006163f
C4077 VDD.n2757 GND 0.006163f
C4078 VDD.n2758 GND 0.006163f
C4079 VDD.n2759 GND 0.350237f
C4080 VDD.n2760 GND 0.006163f
C4081 VDD.n2761 GND 0.006163f
C4082 VDD.n2762 GND 0.006163f
C4083 VDD.n2763 GND 0.006163f
C4084 VDD.n2764 GND 0.006163f
C4085 VDD.n2765 GND 0.006163f
C4086 VDD.n2766 GND 0.006163f
C4087 VDD.n2767 GND 0.006163f
C4088 VDD.n2768 GND 0.350237f
C4089 VDD.n2769 GND 0.006163f
C4090 VDD.n2770 GND 0.006163f
C4091 VDD.n2771 GND 0.006163f
C4092 VDD.n2772 GND 0.006163f
C4093 VDD.n2773 GND 0.006163f
C4094 VDD.n2774 GND 0.006163f
C4095 VDD.n2775 GND 0.006163f
C4096 VDD.n2776 GND 0.006163f
C4097 VDD.n2777 GND 0.006163f
C4098 VDD.n2778 GND 0.006163f
C4099 VDD.n2779 GND 0.006163f
C4100 VDD.n2780 GND 0.006163f
C4101 VDD.n2781 GND 0.006163f
C4102 VDD.n2782 GND 0.006163f
C4103 VDD.n2783 GND 0.006163f
C4104 VDD.n2784 GND 0.006163f
C4105 VDD.n2785 GND 0.006163f
C4106 VDD.n2786 GND 0.006163f
C4107 VDD.n2787 GND 0.006163f
C4108 VDD.n2788 GND 0.006163f
C4109 VDD.n2789 GND 0.006163f
C4110 VDD.n2790 GND 0.006163f
C4111 VDD.n2791 GND 0.006163f
C4112 VDD.n2792 GND 0.013688f
C4113 VDD.n2794 GND 0.014409f
C4114 VDD.n2795 GND 0.014409f
C4115 VDD.n2796 GND 0.006163f
C4116 VDD.n2797 GND 0.004487f
C4117 VDD.n2798 GND 0.006163f
C4118 VDD.n2800 GND 0.006163f
C4119 VDD.n2802 GND 0.006163f
C4120 VDD.n2803 GND 0.006163f
C4121 VDD.n2804 GND 0.006163f
C4122 VDD.n2805 GND 0.006163f
C4123 VDD.n2806 GND 0.006163f
C4124 VDD.n2808 GND 0.006163f
C4125 VDD.n2810 GND 0.006163f
C4126 VDD.n2811 GND 0.006163f
C4127 VDD.n2812 GND 0.006163f
C4128 VDD.n2813 GND 0.006163f
C4129 VDD.n2814 GND 0.006163f
C4130 VDD.n2816 GND 0.006163f
C4131 VDD.n2818 GND 0.006163f
C4132 VDD.n2819 GND 0.006163f
C4133 VDD.n2820 GND 0.006163f
C4134 VDD.n2821 GND 0.006163f
C4135 VDD.n2822 GND 0.006163f
C4136 VDD.n2824 GND 0.006163f
C4137 VDD.n2826 GND 0.006163f
C4138 VDD.n2827 GND 0.006163f
C4139 VDD.n2828 GND 0.006163f
C4140 VDD.n2829 GND 0.006163f
C4141 VDD.n2830 GND 0.006163f
C4142 VDD.n2832 GND 0.006163f
C4143 VDD.n2834 GND 0.006163f
C4144 VDD.n2835 GND 0.006163f
C4145 VDD.n2836 GND 0.006163f
C4146 VDD.n2837 GND 0.006163f
C4147 VDD.n2838 GND 0.006163f
C4148 VDD.n2840 GND 0.006163f
C4149 VDD.n2842 GND 0.006163f
C4150 VDD.n2843 GND 0.006163f
C4151 VDD.n2844 GND 0.014409f
C4152 VDD.n2845 GND 0.013688f
C4153 VDD.n2846 GND 0.013688f
C4154 VDD.n2847 GND 0.723566f
C4155 VDD.n2848 GND 0.013688f
C4156 VDD.n2849 GND 0.013688f
C4157 VDD.n2850 GND 0.006163f
C4158 VDD.n2851 GND 0.006163f
C4159 VDD.n2852 GND 0.006163f
C4160 VDD.n2853 GND 0.361783f
C4161 VDD.n2854 GND 0.006163f
C4162 VDD.n2855 GND 0.006163f
C4163 VDD.n2856 GND 0.006163f
C4164 VDD.n2857 GND 0.006163f
C4165 VDD.n2858 GND 0.006163f
C4166 VDD.n2859 GND 0.49649f
C4167 VDD.n2860 GND 0.006163f
C4168 VDD.n2861 GND 0.006163f
C4169 VDD.n2862 GND 0.006163f
C4170 VDD.n2863 GND 0.006163f
C4171 VDD.n2864 GND 0.006163f
C4172 VDD.n2865 GND 0.384876f
C4173 VDD.n2866 GND 0.006163f
C4174 VDD.n2867 GND 0.006163f
C4175 VDD.n2868 GND 0.006163f
C4176 VDD.n2869 GND 0.006163f
C4177 VDD.n2870 GND 0.006163f
C4178 VDD.n2871 GND 0.523431f
C4179 VDD.n2872 GND 0.006163f
C4180 VDD.n2873 GND 0.006163f
C4181 VDD.n2874 GND 0.006163f
C4182 VDD.n2875 GND 0.006163f
C4183 VDD.n2876 GND 0.006163f
C4184 VDD.n2877 GND 0.203984f
C4185 VDD.n2878 GND 0.006163f
C4186 VDD.n2879 GND 0.006163f
C4187 VDD.n2880 GND 0.006163f
C4188 VDD.n2881 GND 0.006163f
C4189 VDD.n2882 GND 0.006163f
C4190 VDD.n2883 GND 0.523431f
C4191 VDD.n2884 GND 0.006163f
C4192 VDD.n2885 GND 0.006163f
C4193 VDD.n2886 GND 0.006163f
C4194 VDD.n2887 GND 0.006163f
C4195 VDD.n2888 GND 0.006163f
C4196 VDD.n2889 GND 0.296354f
C4197 VDD.n2890 GND 0.006163f
C4198 VDD.n2891 GND 0.006163f
C4199 VDD.n2892 GND 0.006163f
C4200 VDD.n2893 GND 0.006163f
C4201 VDD.n2894 GND 0.006163f
C4202 VDD.n2895 GND 0.400271f
C4203 VDD.n2896 GND 0.006163f
C4204 VDD.n2897 GND 0.006163f
C4205 VDD.n2898 GND 0.006163f
C4206 VDD.n2899 GND 0.006163f
C4207 VDD.n2900 GND 0.006163f
C4208 VDD.n2901 GND 0.273262f
C4209 VDD.n2902 GND 0.006163f
C4210 VDD.n2903 GND 0.006163f
C4211 VDD.n2904 GND 0.006163f
C4212 VDD.n2905 GND 0.006163f
C4213 VDD.n2906 GND 0.006163f
C4214 VDD.n2907 GND 0.423363f
C4215 VDD.n2908 GND 0.006163f
C4216 VDD.n2909 GND 0.006163f
C4217 VDD.n2910 GND 0.006163f
C4218 VDD.n2911 GND 0.006163f
C4219 VDD.n2912 GND 0.006163f
C4220 VDD.n2913 GND 0.273262f
C4221 VDD.n2914 GND 0.006163f
C4222 VDD.n2915 GND 0.006163f
C4223 VDD.n2916 GND 0.006163f
C4224 VDD.n2917 GND 0.006163f
C4225 VDD.n2918 GND 0.006163f
C4226 VDD.n2919 GND 0.446456f
C4227 VDD.n2920 GND 0.006163f
C4228 VDD.n2921 GND 0.006163f
C4229 VDD.n2922 GND 0.006163f
C4230 VDD.n2923 GND 0.006163f
C4231 VDD.n2924 GND 0.006163f
C4232 VDD.n2925 GND 0.296354f
C4233 VDD.n2926 GND 0.006163f
C4234 VDD.n2927 GND 0.006163f
C4235 VDD.n2928 GND 0.006163f
C4236 VDD.n2929 GND 0.006163f
C4237 VDD.n2930 GND 0.006163f
C4238 VDD.n2931 GND 0.469548f
C4239 VDD.n2932 GND 0.006163f
C4240 VDD.n2933 GND 0.006163f
C4241 VDD.n2934 GND 0.006163f
C4242 VDD.n2935 GND 0.006163f
C4243 VDD.n2936 GND 0.006163f
C4244 VDD.n2937 GND 0.319447f
C4245 VDD.n2938 GND 0.006163f
C4246 VDD.n2939 GND 0.006163f
C4247 VDD.n2940 GND 0.006163f
C4248 VDD.n2941 GND 0.006163f
C4249 VDD.n2942 GND 0.006163f
C4250 VDD.n2943 GND 0.523431f
C4251 VDD.n2944 GND 0.006163f
C4252 VDD.n2945 GND 0.006163f
C4253 VDD.n2946 GND 0.006163f
C4254 VDD.n2947 GND 0.006163f
C4255 VDD.n2948 GND 0.006163f
C4256 VDD.n2949 GND 0.346388f
C4257 VDD.n2950 GND 0.006163f
C4258 VDD.n2951 GND 0.004079f
C4259 VDD.n2952 GND 0.017854f
C4260 VDD.n2953 GND 0.005166f
C4261 VDD.n2954 GND 0.006163f
C4262 VDD.n2955 GND 0.006163f
C4263 VDD.n2956 GND 0.006163f
C4264 VDD.n2957 GND 0.006163f
C4265 VDD.n2959 GND 0.006163f
C4266 VDD.n2960 GND 0.006163f
C4267 VDD.n2962 GND 0.006163f
C4268 VDD.n2963 GND 0.006163f
C4269 VDD.n2964 GND 0.006163f
C4270 VDD.n2966 GND 0.006163f
C4271 VDD.n2967 GND 0.006163f
C4272 VDD.n2968 GND 0.006163f
C4273 VDD.n2969 GND 0.006163f
C4274 VDD.n2970 GND 0.006163f
C4275 VDD.n2971 GND 0.006163f
C4276 VDD.n2973 GND 0.006163f
C4277 VDD.n2974 GND 0.006163f
C4278 VDD.n2975 GND 0.006163f
C4279 VDD.n2976 GND 0.006163f
C4280 VDD.n2977 GND 0.006163f
C4281 VDD.n2978 GND 0.006163f
C4282 VDD.n2980 GND 0.006163f
C4283 VDD.n2981 GND 0.006163f
C4284 VDD.n2983 GND 0.014409f
C4285 VDD.n2984 GND 0.014409f
C4286 VDD.n2985 GND 0.013688f
C4287 VDD.n2986 GND 0.006163f
C4288 VDD.n2987 GND 0.006163f
C4289 VDD.n2988 GND 0.006163f
C4290 VDD.n2989 GND 0.006163f
C4291 VDD.n2990 GND 0.006163f
C4292 VDD.n2991 GND 0.006163f
C4293 VDD.n2992 GND 0.49649f
C4294 VDD.n2993 GND 0.006163f
C4295 VDD.n2994 GND 0.006163f
C4296 VDD.n2995 GND 0.006163f
C4297 VDD.n2996 GND 0.006163f
C4298 VDD.n2997 GND 0.006163f
C4299 VDD.n2998 GND 0.523431f
C4300 VDD.n2999 GND 0.006163f
C4301 VDD.n3000 GND 0.006163f
C4302 VDD.n3001 GND 0.006163f
C4303 VDD.n3002 GND 0.014446f
C4304 VDD.n3004 GND 0.014409f
C4305 VDD.n3005 GND 0.013651f
C4306 VDD.n3006 GND 0.006163f
C4307 VDD.n3007 GND 0.004487f
C4308 VDD.n3008 GND 0.006163f
C4309 VDD.n3010 GND 0.006163f
C4310 VDD.n3011 GND 0.006163f
C4311 VDD.n3012 GND 0.006163f
C4312 VDD.n3013 GND 0.006163f
C4313 VDD.n3014 GND 0.006163f
C4314 VDD.n3015 GND 0.006163f
C4315 VDD.n3017 GND 0.006163f
C4316 VDD.n3018 GND 0.006163f
C4317 VDD.n3019 GND 0.006163f
C4318 VDD.n3020 GND 0.006163f
C4319 VDD.n3021 GND 0.006163f
C4320 VDD.n3022 GND 0.006163f
C4321 VDD.n3024 GND 0.006163f
C4322 VDD.n3025 GND 0.006163f
C4323 VDD.n3026 GND 0.004622f
C4324 VDD.n3027 GND 0.463254f
C4325 VDD.n3028 GND 0.008598f
C4326 VDD.n3029 GND 0.004622f
C4327 VDD.n3030 GND 0.006163f
C4328 VDD.n3031 GND 0.006163f
C4329 VDD.n3033 GND 0.006163f
C4330 VDD.n3034 GND 0.006163f
C4331 VDD.n3035 GND 0.006163f
C4332 VDD.n3036 GND 0.006163f
C4333 VDD.n3037 GND 0.006163f
C4334 VDD.n3038 GND 0.006163f
C4335 VDD.n3040 GND 0.006163f
C4336 VDD.n3041 GND 0.006163f
C4337 VDD.n3042 GND 0.006163f
C4338 VDD.n3043 GND 0.006163f
C4339 VDD.n3044 GND 0.006163f
C4340 VDD.n3045 GND 0.006163f
C4341 VDD.n3047 GND 0.006163f
C4342 VDD.n3048 GND 0.006163f
C4343 VDD.n3049 GND 0.006163f
C4344 VDD.n3050 GND 0.014409f
C4345 VDD.n3051 GND 0.013688f
C4346 VDD.n3052 GND 0.013688f
C4347 VDD.n3053 GND 0.723566f
C4348 VDD.n3054 GND 0.013688f
C4349 VDD.n3055 GND 0.014409f
C4350 VDD.n3056 GND 0.013651f
C4351 VDD.n3057 GND 0.006163f
C4352 VDD.n3058 GND 0.004487f
C4353 VDD.n3059 GND 0.006163f
C4354 VDD.n3061 GND 0.006163f
C4355 VDD.n3062 GND 0.006163f
C4356 VDD.n3063 GND 0.006163f
C4357 VDD.n3064 GND 0.006163f
C4358 VDD.n3065 GND 0.006163f
C4359 VDD.n3066 GND 0.006163f
C4360 VDD.n3068 GND 0.006163f
C4361 VDD.n3069 GND 0.006163f
C4362 VDD.n3070 GND 0.006163f
C4363 VDD.n3071 GND 0.006163f
C4364 VDD.n3072 GND 0.006163f
C4365 VDD.n3073 GND 0.006163f
C4366 VDD.n3075 GND 0.006163f
C4367 VDD.n3076 GND 0.006163f
C4368 VDD.n3077 GND 0.004622f
C4369 VDD.n3078 GND 0.008598f
C4370 VDD.n3079 GND 0.463254f
C4371 VDD.n3080 GND 0.007795f
C4372 VDD.n3081 GND 0.009064f
C4373 VDD.n3082 GND 0.009064f
C4374 VDD.n3083 GND 0.009064f
C4375 VDD.n3084 GND 0.009064f
C4376 VDD.n3085 GND 0.009064f
C4377 VDD.n3086 GND 0.00383f
C4378 VDD.n3087 GND 0.007295f
C4379 VDD.n3088 GND 0.009064f
C4380 VDD.n3089 GND 0.009064f
C4381 VDD.n3090 GND 0.007295f
C4382 VDD.n3091 GND 0.007295f
C4383 VDD.n3092 GND 0.009064f
C4384 VDD.n3093 GND 0.009064f
C4385 VDD.n3094 GND 0.007295f
C4386 VDD.n3095 GND 0.007295f
C4387 VDD.n3096 GND 0.009064f
C4388 VDD.n3097 GND 0.009064f
C4389 VDD.n3098 GND 0.007295f
C4390 VDD.n3099 GND 0.007295f
C4391 VDD.n3100 GND 0.009064f
C4392 VDD.n3101 GND 0.009064f
C4393 VDD.n3102 GND 0.007295f
C4394 VDD.n3103 GND 0.007295f
C4395 VDD.n3104 GND 0.009064f
C4396 VDD.n3105 GND 0.009064f
C4397 VDD.n3106 GND 0.007295f
C4398 VDD.n3107 GND 0.007295f
C4399 VDD.n3108 GND 0.009064f
C4400 VDD.n3109 GND 0.009064f
C4401 VDD.n3110 GND 0.007295f
C4402 VDD.n3111 GND 0.007295f
C4403 VDD.n3112 GND 0.009064f
C4404 VDD.n3113 GND 0.009064f
C4405 VDD.n3114 GND 0.007295f
C4406 VDD.n3115 GND 0.007295f
C4407 VDD.n3116 GND 0.009064f
C4408 VDD.n3117 GND 0.009064f
C4409 VDD.n3118 GND 0.007295f
C4410 VDD.n3119 GND 0.007295f
C4411 VDD.n3120 GND 0.009064f
C4412 VDD.n3121 GND 0.009064f
C4413 VDD.n3122 GND 0.007295f
C4414 VDD.n3123 GND 0.009064f
C4415 VDD.n3124 GND 0.009064f
C4416 VDD.n3125 GND 0.007295f
C4417 VDD.n3126 GND 0.009064f
C4418 VDD.n3127 GND 0.009064f
C4419 VDD.n3128 GND 0.009064f
C4420 VDD.n3129 GND 0.014919f
C4421 VDD.n3130 GND 0.009064f
C4422 VDD.n3131 GND 0.009064f
C4423 VDD.n3132 GND 0.004961f
C4424 VDD.n3133 GND 0.007295f
C4425 VDD.n3134 GND 0.009064f
C4426 VDD.n3135 GND 0.009064f
C4427 VDD.n3136 GND 0.007295f
C4428 VDD.n3137 GND 0.007295f
C4429 VDD.n3138 GND 0.009064f
C4430 VDD.n3139 GND 0.009064f
C4431 VDD.n3140 GND 0.007295f
C4432 VDD.n3141 GND 0.007295f
C4433 VDD.n3142 GND 0.009064f
C4434 VDD.n3143 GND 0.009064f
C4435 VDD.n3144 GND 0.007295f
C4436 VDD.n3145 GND 0.007295f
C4437 VDD.n3146 GND 0.009064f
C4438 VDD.n3147 GND 0.009064f
C4439 VDD.n3148 GND 0.007295f
C4440 VDD.n3149 GND 0.007295f
C4441 VDD.n3150 GND 0.009064f
C4442 VDD.n3151 GND 0.009064f
C4443 VDD.n3152 GND 0.007295f
C4444 VDD.n3153 GND 0.007295f
C4445 VDD.n3154 GND 0.009064f
C4446 VDD.n3155 GND 0.009064f
C4447 VDD.n3156 GND 0.007295f
C4448 VDD.n3157 GND 0.007295f
C4449 VDD.n3158 GND 0.009064f
C4450 VDD.n3159 GND 0.009064f
C4451 VDD.n3160 GND 0.007295f
C4452 VDD.n3161 GND 0.007295f
C4453 VDD.n3162 GND 0.009064f
C4454 VDD.n3163 GND 0.009064f
C4455 VDD.n3164 GND 0.007295f
C4456 VDD.n3165 GND 0.007295f
C4457 VDD.n3166 GND 0.009064f
C4458 VDD.n3167 GND 0.009064f
C4459 VDD.n3168 GND 0.007295f
C4460 VDD.n3169 GND 0.009064f
C4461 VDD.n3170 GND 0.009064f
C4462 VDD.n3171 GND 0.007295f
C4463 VDD.n3172 GND 0.009064f
C4464 VDD.n3173 GND 0.009064f
C4465 VDD.n3174 GND 0.009064f
C4466 VDD.t11 GND 0.111507f
C4467 VDD.t12 GND 0.123568f
C4468 VDD.t10 GND 0.30702f
C4469 VDD.n3175 GND 0.203209f
C4470 VDD.n3176 GND 0.158699f
C4471 VDD.n3177 GND 0.014919f
C4472 VDD.n3178 GND 0.009064f
C4473 VDD.n3179 GND 0.009064f
C4474 VDD.n3180 GND 0.006091f
C4475 VDD.n3181 GND 0.007295f
C4476 VDD.n3182 GND 0.009064f
C4477 VDD.n3183 GND 0.009064f
C4478 VDD.n3184 GND 0.007295f
C4479 VDD.n3185 GND 0.007295f
C4480 VDD.n3186 GND 0.009064f
C4481 VDD.n3187 GND 0.009064f
C4482 VDD.n3188 GND 0.007295f
C4483 VDD.n3189 GND 0.007295f
C4484 VDD.n3190 GND 0.009064f
C4485 VDD.n3191 GND 0.009064f
C4486 VDD.n3192 GND 0.007295f
C4487 VDD.n3193 GND 0.007295f
C4488 VDD.n3194 GND 0.009064f
C4489 VDD.n3195 GND 0.009064f
C4490 VDD.n3196 GND 0.007295f
C4491 VDD.n3197 GND 0.007295f
C4492 VDD.n3198 GND 0.009064f
C4493 VDD.n3199 GND 0.009064f
C4494 VDD.n3200 GND 0.007295f
C4495 VDD.n3201 GND 0.007295f
C4496 VDD.n3202 GND 0.009064f
C4497 VDD.n3203 GND 0.009064f
C4498 VDD.n3204 GND 0.007295f
C4499 VDD.n3205 GND 0.007295f
C4500 VDD.n3206 GND 0.009064f
C4501 VDD.n3207 GND 0.009064f
C4502 VDD.n3208 GND 0.007295f
C4503 VDD.n3209 GND 0.009064f
C4504 VDD.n3210 GND 0.007295f
C4505 VDD.n3211 GND 0.007295f
C4506 VDD.n3212 GND 0.007295f
C4507 VDD.n3213 GND 0.006055f
C4508 VDD.n3214 GND 0.021239f
C4509 VDD.n3216 GND 4.70703f
C4510 VDD.n3217 GND 0.021239f
C4511 VDD.n3218 GND 0.003465f
C4512 VDD.n3219 GND 0.021239f
C4513 VDD.n3220 GND 0.020998f
C4514 VDD.n3221 GND 0.009064f
C4515 VDD.n3222 GND 0.007295f
C4516 VDD.n3223 GND 0.009064f
C4517 VDD.t3 GND 0.384876f
C4518 VDD.n3224 GND 0.58886f
C4519 VDD.n3225 GND 0.009064f
C4520 VDD.n3226 GND 0.007295f
C4521 VDD.n3227 GND 0.009064f
C4522 VDD.n3228 GND 0.009064f
C4523 VDD.n3229 GND 0.009064f
C4524 VDD.n3230 GND 0.007295f
C4525 VDD.n3231 GND 0.009064f
C4526 VDD.n3232 GND 0.769751f
C4527 VDD.n3233 GND 0.009064f
C4528 VDD.n3234 GND 0.007295f
C4529 VDD.n3235 GND 0.009064f
C4530 VDD.n3236 GND 0.009064f
C4531 VDD.n3237 GND 0.009064f
C4532 VDD.n3238 GND 0.007295f
C4533 VDD.n3239 GND 0.009064f
C4534 VDD.n3240 GND 0.52728f
C4535 VDD.n3241 GND 0.769751f
C4536 VDD.n3242 GND 0.009064f
C4537 VDD.n3243 GND 0.007295f
C4538 VDD.n3244 GND 0.009064f
C4539 VDD.n3245 GND 0.009064f
C4540 VDD.n3246 GND 0.009064f
C4541 VDD.n3247 GND 0.007295f
C4542 VDD.n3248 GND 0.009064f
C4543 VDD.n3249 GND 0.627347f
C4544 VDD.n3250 GND 0.009064f
C4545 VDD.n3251 GND 0.007295f
C4546 VDD.n3252 GND 0.009064f
C4547 VDD.n3253 GND 0.009064f
C4548 VDD.n3254 GND 0.009064f
C4549 VDD.n3255 GND 0.007295f
C4550 VDD.n3256 GND 0.009064f
C4551 VDD.t157 GND 0.384876f
C4552 VDD.n3257 GND 0.396422f
C4553 VDD.n3258 GND 0.009064f
C4554 VDD.n3259 GND 0.007295f
C4555 VDD.n3260 GND 0.009064f
C4556 VDD.n3261 GND 0.009064f
C4557 VDD.n3262 GND 0.009064f
C4558 VDD.n3263 GND 0.007295f
C4559 VDD.n3264 GND 0.009064f
C4560 VDD.n3265 GND 0.65044f
C4561 VDD.n3266 GND 0.009064f
C4562 VDD.n3267 GND 0.007295f
C4563 VDD.n3268 GND 0.009064f
C4564 VDD.n3269 GND 0.009064f
C4565 VDD.n3270 GND 0.009064f
C4566 VDD.n3271 GND 0.007295f
C4567 VDD.n3272 GND 0.009064f
C4568 VDD.n3273 GND 0.519582f
C4569 VDD.n3274 GND 0.769751f
C4570 VDD.n3275 GND 0.009064f
C4571 VDD.n3276 GND 0.007295f
C4572 VDD.n3277 GND 0.009064f
C4573 VDD.n3278 GND 0.009064f
C4574 VDD.n3279 GND 0.009064f
C4575 VDD.n3280 GND 0.007295f
C4576 VDD.n3281 GND 0.009064f
C4577 VDD.n3282 GND 0.635045f
C4578 VDD.n3283 GND 0.009064f
C4579 VDD.n3284 GND 0.007295f
C4580 VDD.n3285 GND 0.009064f
C4581 VDD.n3286 GND 0.009064f
C4582 VDD.n3287 GND 0.009064f
C4583 VDD.n3288 GND 0.009064f
C4584 VDD.n3289 GND 0.009064f
C4585 VDD.n3290 GND 0.007295f
C4586 VDD.n3291 GND 0.007295f
C4587 VDD.n3292 GND 0.009064f
C4588 VDD.t97 GND 0.384876f
C4589 VDD.n3293 GND 0.388724f
C4590 VDD.n3294 GND 0.009064f
C4591 VDD.n3295 GND 0.007295f
C4592 VDD.n3296 GND 0.009064f
C4593 VDD.n3297 GND 0.009064f
C4594 VDD.n3298 GND 0.009064f
C4595 VDD.n3299 GND 0.007295f
C4596 VDD.n3300 GND 0.009064f
C4597 VDD.n3301 GND 0.642742f
C4598 VDD.n3302 GND 0.009064f
C4599 VDD.n3303 GND 0.009064f
C4600 VDD.n3304 GND 0.007295f
C4601 VDD.n3305 GND 0.007295f
C4602 VDD.n3306 GND 0.007295f
C4603 VDD.n3307 GND 0.009064f
C4604 VDD.n3308 GND 0.009064f
C4605 VDD.n3309 GND 0.009064f
C4606 VDD.n3310 GND 0.009064f
C4607 VDD.n3311 GND 0.007295f
C4608 VDD.n3312 GND 0.007295f
C4609 VDD.n3313 GND 0.007295f
C4610 VDD.n3314 GND 0.009064f
C4611 VDD.n3315 GND 0.009064f
C4612 VDD.n3316 GND 0.009064f
C4613 VDD.n3317 GND 0.009064f
C4614 VDD.n3318 GND 0.007295f
C4615 VDD.n3319 GND 0.007295f
C4616 VDD.n3320 GND 0.007295f
C4617 VDD.n3321 GND 0.009064f
C4618 VDD.n3322 GND 0.009064f
C4619 VDD.n3323 GND 0.009064f
C4620 VDD.n3324 GND 0.009064f
C4621 VDD.n3325 GND 0.007295f
C4622 VDD.n3326 GND 0.007295f
C4623 VDD.n3327 GND 0.007295f
C4624 VDD.n3328 GND 0.009064f
C4625 VDD.n3329 GND 0.009064f
C4626 VDD.n3330 GND 0.009064f
C4627 VDD.n3331 GND 0.009064f
C4628 VDD.n3332 GND 0.007295f
C4629 VDD.n3333 GND 0.007295f
C4630 VDD.n3334 GND 0.007295f
C4631 VDD.n3335 GND 0.009064f
C4632 VDD.n3336 GND 0.009064f
C4633 VDD.n3337 GND 0.009064f
C4634 VDD.n3338 GND 0.009064f
C4635 VDD.n3339 GND 0.007295f
C4636 VDD.n3340 GND 0.007295f
C4637 VDD.n3341 GND 0.006055f
C4638 VDD.n3342 GND 0.020998f
C4639 VDD.n3343 GND 0.021239f
C4640 VDD.n3344 GND 0.003465f
C4641 VDD.n3345 GND 0.021239f
C4642 VDD.n3347 GND 1.73579f
C4643 VDD.n3348 GND 1.05071f
C4644 VDD.n3349 GND 0.58886f
C4645 VDD.n3350 GND 0.009064f
C4646 VDD.n3351 GND 0.007295f
C4647 VDD.n3352 GND 0.007295f
C4648 VDD.n3353 GND 0.007295f
C4649 VDD.n3354 GND 0.009064f
C4650 VDD.n3355 GND 0.769751f
C4651 VDD.n3356 GND 0.769751f
C4652 VDD.n3357 GND 0.769751f
C4653 VDD.n3358 GND 0.009064f
C4654 VDD.n3359 GND 0.007295f
C4655 VDD.n3360 GND 0.007295f
C4656 VDD.n3361 GND 0.007295f
C4657 VDD.n3362 GND 0.009064f
C4658 VDD.n3363 GND 0.627347f
C4659 VDD.n3364 GND 0.769751f
C4660 VDD.n3365 GND 0.396422f
C4661 VDD.n3366 GND 0.009064f
C4662 VDD.n3367 GND 0.007295f
C4663 VDD.n3368 GND 0.007295f
C4664 VDD.n3369 GND 0.007295f
C4665 VDD.n3370 GND 0.009064f
C4666 VDD.n3371 GND 0.65044f
C4667 VDD.t95 GND 0.384876f
C4668 VDD.n3372 GND 0.504187f
C4669 VDD.n3373 GND 0.769751f
C4670 VDD.n3374 GND 0.009064f
C4671 VDD.n3375 GND 0.007295f
C4672 VDD.n3376 GND 0.007295f
C4673 VDD.n3377 GND 0.007295f
C4674 VDD.n3378 GND 0.009064f
C4675 VDD.n3379 GND 0.635045f
C4676 VDD.n3380 GND 0.769751f
C4677 VDD.n3381 GND 0.388724f
C4678 VDD.n3382 GND 0.009064f
C4679 VDD.n3383 GND 0.007295f
C4680 VDD.n3384 GND 0.007295f
C4681 VDD.n3385 GND 0.007295f
C4682 VDD.n3386 GND 0.009064f
C4683 VDD.n3387 GND 0.642742f
C4684 VDD.t155 GND 0.384876f
C4685 VDD.n3388 GND 0.511885f
C4686 VDD.n3389 GND 0.769751f
C4687 VDD.n3390 GND 0.009064f
C4688 VDD.n3391 GND 0.007295f
C4689 VDD.n3392 GND 0.200692f
C4690 VDD.n3393 GND 1.92438f
C4691 VOUT.t35 GND 0.049715f
C4692 VOUT.t60 GND 0.049715f
C4693 VOUT.n0 GND 0.385563f
C4694 VOUT.t66 GND 0.049715f
C4695 VOUT.t18 GND 0.049715f
C4696 VOUT.n1 GND 0.384224f
C4697 VOUT.n2 GND 0.476712f
C4698 VOUT.t1 GND 0.049715f
C4699 VOUT.t29 GND 0.049715f
C4700 VOUT.n3 GND 0.384224f
C4701 VOUT.n4 GND 0.235858f
C4702 VOUT.t22 GND 0.049715f
C4703 VOUT.t55 GND 0.049715f
C4704 VOUT.n5 GND 0.384224f
C4705 VOUT.n6 GND 0.235858f
C4706 VOUT.t19 GND 0.049715f
C4707 VOUT.t34 GND 0.049715f
C4708 VOUT.n7 GND 0.384224f
C4709 VOUT.n8 GND 0.235858f
C4710 VOUT.t6 GND 0.049715f
C4711 VOUT.t27 GND 0.049715f
C4712 VOUT.n9 GND 0.384224f
C4713 VOUT.n10 GND 0.406983f
C4714 VOUT.t36 GND 0.049715f
C4715 VOUT.t57 GND 0.049715f
C4716 VOUT.n11 GND 0.385563f
C4717 VOUT.t69 GND 0.049715f
C4718 VOUT.t3 GND 0.049715f
C4719 VOUT.n12 GND 0.384224f
C4720 VOUT.n13 GND 0.476712f
C4721 VOUT.t44 GND 0.049715f
C4722 VOUT.t48 GND 0.049715f
C4723 VOUT.n14 GND 0.384224f
C4724 VOUT.n15 GND 0.235858f
C4725 VOUT.t11 GND 0.049715f
C4726 VOUT.t67 GND 0.049715f
C4727 VOUT.n16 GND 0.384224f
C4728 VOUT.n17 GND 0.235858f
C4729 VOUT.t49 GND 0.049715f
C4730 VOUT.t50 GND 0.049715f
C4731 VOUT.n18 GND 0.384224f
C4732 VOUT.n19 GND 0.235858f
C4733 VOUT.t33 GND 0.049715f
C4734 VOUT.t45 GND 0.049715f
C4735 VOUT.n20 GND 0.384224f
C4736 VOUT.n21 GND 0.327356f
C4737 VOUT.n22 GND 0.665002f
C4738 VOUT.t5 GND 0.049715f
C4739 VOUT.t38 GND 0.049715f
C4740 VOUT.n23 GND 0.385563f
C4741 VOUT.t46 GND 0.049715f
C4742 VOUT.t63 GND 0.049715f
C4743 VOUT.n24 GND 0.384224f
C4744 VOUT.n25 GND 0.476712f
C4745 VOUT.t61 GND 0.049715f
C4746 VOUT.t4 GND 0.049715f
C4747 VOUT.n26 GND 0.384224f
C4748 VOUT.n27 GND 0.235858f
C4749 VOUT.t64 GND 0.049715f
C4750 VOUT.t65 GND 0.049715f
C4751 VOUT.n28 GND 0.384224f
C4752 VOUT.n29 GND 0.235858f
C4753 VOUT.t12 GND 0.049715f
C4754 VOUT.t8 GND 0.049715f
C4755 VOUT.n30 GND 0.384224f
C4756 VOUT.n31 GND 0.235858f
C4757 VOUT.t59 GND 0.049715f
C4758 VOUT.t41 GND 0.049715f
C4759 VOUT.n32 GND 0.384224f
C4760 VOUT.n33 GND 0.327356f
C4761 VOUT.n34 GND 0.600494f
C4762 VOUT.n35 GND 7.1915f
C4763 VOUT.n37 GND 0.705049f
C4764 VOUT.n38 GND 0.528787f
C4765 VOUT.n39 GND 0.705049f
C4766 VOUT.n40 GND 0.705049f
C4767 VOUT.n41 GND 1.89821f
C4768 VOUT.n42 GND 0.705049f
C4769 VOUT.n43 GND 0.705049f
C4770 VOUT.t112 GND 0.881311f
C4771 VOUT.n44 GND 0.705049f
C4772 VOUT.n45 GND 0.705049f
C4773 VOUT.n49 GND 0.705049f
C4774 VOUT.n53 GND 0.705049f
C4775 VOUT.n54 GND 0.705049f
C4776 VOUT.n56 GND 0.705049f
C4777 VOUT.n61 GND 0.705049f
C4778 VOUT.n63 GND 0.705049f
C4779 VOUT.n64 GND 0.705049f
C4780 VOUT.n66 GND 0.705049f
C4781 VOUT.n67 GND 0.705049f
C4782 VOUT.n69 GND 0.705049f
C4783 VOUT.t115 GND 11.7813f
C4784 VOUT.n71 GND 0.705049f
C4785 VOUT.n72 GND 0.528787f
C4786 VOUT.n73 GND 0.705049f
C4787 VOUT.n74 GND 0.705049f
C4788 VOUT.n75 GND 1.89821f
C4789 VOUT.n76 GND 0.705049f
C4790 VOUT.n77 GND 0.705049f
C4791 VOUT.t117 GND 0.881311f
C4792 VOUT.n78 GND 0.705049f
C4793 VOUT.n79 GND 0.705049f
C4794 VOUT.n83 GND 0.705049f
C4795 VOUT.n87 GND 0.705049f
C4796 VOUT.n88 GND 0.705049f
C4797 VOUT.n90 GND 0.705049f
C4798 VOUT.n95 GND 0.705049f
C4799 VOUT.n97 GND 0.705049f
C4800 VOUT.n98 GND 0.705049f
C4801 VOUT.n100 GND 0.705049f
C4802 VOUT.n101 GND 0.705049f
C4803 VOUT.n103 GND 0.705049f
C4804 VOUT.n104 GND 0.528787f
C4805 VOUT.n106 GND 0.705049f
C4806 VOUT.n107 GND 0.528787f
C4807 VOUT.n108 GND 0.705049f
C4808 VOUT.n109 GND 0.705049f
C4809 VOUT.n110 GND 1.89821f
C4810 VOUT.n111 GND 0.705049f
C4811 VOUT.n112 GND 0.705049f
C4812 VOUT.t116 GND 0.881311f
C4813 VOUT.n113 GND 0.705049f
C4814 VOUT.n114 GND 1.89821f
C4815 VOUT.n116 GND 0.705049f
C4816 VOUT.n117 GND 0.705049f
C4817 VOUT.n119 GND 0.705049f
C4818 VOUT.n120 GND 0.705049f
C4819 VOUT.t113 GND 11.589299f
C4820 VOUT.t114 GND 11.7813f
C4821 VOUT.n126 GND 2.21184f
C4822 VOUT.n127 GND 9.010241f
C4823 VOUT.n128 GND 9.387259f
C4824 VOUT.n133 GND 2.39602f
C4825 VOUT.n139 GND 0.705049f
C4826 VOUT.n141 GND 0.705049f
C4827 VOUT.n143 GND 0.705049f
C4828 VOUT.n145 GND 0.705049f
C4829 VOUT.n147 GND 0.705049f
C4830 VOUT.n153 GND 0.705049f
C4831 VOUT.n160 GND 1.29349f
C4832 VOUT.n161 GND 1.29349f
C4833 VOUT.n162 GND 0.705049f
C4834 VOUT.n163 GND 0.705049f
C4835 VOUT.n165 GND 0.528787f
C4836 VOUT.n166 GND 0.452858f
C4837 VOUT.n168 GND 0.528787f
C4838 VOUT.n169 GND 0.452858f
C4839 VOUT.n170 GND 0.528787f
C4840 VOUT.n172 GND 0.705049f
C4841 VOUT.n174 GND 1.89821f
C4842 VOUT.n175 GND 2.21184f
C4843 VOUT.n176 GND 8.287099f
C4844 VOUT.n178 GND 0.528787f
C4845 VOUT.n179 GND 1.3606f
C4846 VOUT.n180 GND 0.528787f
C4847 VOUT.n182 GND 0.705049f
C4848 VOUT.n184 GND 1.89821f
C4849 VOUT.n185 GND 3.52915f
C4850 VOUT.n186 GND 2.36321f
C4851 VOUT.t7 GND 0.049715f
C4852 VOUT.t37 GND 0.049715f
C4853 VOUT.n187 GND 0.385563f
C4854 VOUT.t31 GND 0.049715f
C4855 VOUT.t68 GND 0.049715f
C4856 VOUT.n188 GND 0.384224f
C4857 VOUT.n189 GND 0.476712f
C4858 VOUT.t16 GND 0.049715f
C4859 VOUT.t58 GND 0.049715f
C4860 VOUT.n190 GND 0.384224f
C4861 VOUT.n191 GND 0.235858f
C4862 VOUT.t53 GND 0.049715f
C4863 VOUT.t70 GND 0.049715f
C4864 VOUT.n192 GND 0.384224f
C4865 VOUT.n193 GND 0.235858f
C4866 VOUT.t26 GND 0.049715f
C4867 VOUT.t32 GND 0.049715f
C4868 VOUT.n194 GND 0.384224f
C4869 VOUT.n195 GND 0.235858f
C4870 VOUT.t20 GND 0.049715f
C4871 VOUT.t10 GND 0.049715f
C4872 VOUT.n196 GND 0.384224f
C4873 VOUT.n197 GND 0.406983f
C4874 VOUT.t21 GND 0.049715f
C4875 VOUT.t54 GND 0.049715f
C4876 VOUT.n198 GND 0.385563f
C4877 VOUT.t39 GND 0.049715f
C4878 VOUT.t30 GND 0.049715f
C4879 VOUT.n199 GND 0.384224f
C4880 VOUT.n200 GND 0.476712f
C4881 VOUT.t9 GND 0.049715f
C4882 VOUT.t23 GND 0.049715f
C4883 VOUT.n201 GND 0.384224f
C4884 VOUT.n202 GND 0.235858f
C4885 VOUT.t43 GND 0.049715f
C4886 VOUT.t71 GND 0.049715f
C4887 VOUT.n203 GND 0.384224f
C4888 VOUT.n204 GND 0.235858f
C4889 VOUT.t17 GND 0.049715f
C4890 VOUT.t25 GND 0.049715f
C4891 VOUT.n205 GND 0.384224f
C4892 VOUT.n206 GND 0.235858f
C4893 VOUT.t14 GND 0.049715f
C4894 VOUT.t56 GND 0.049715f
C4895 VOUT.n207 GND 0.384224f
C4896 VOUT.n208 GND 0.327356f
C4897 VOUT.n209 GND 0.665002f
C4898 VOUT.t42 GND 0.049715f
C4899 VOUT.t51 GND 0.049715f
C4900 VOUT.n210 GND 0.385563f
C4901 VOUT.t47 GND 0.049715f
C4902 VOUT.t24 GND 0.049715f
C4903 VOUT.n211 GND 0.384224f
C4904 VOUT.n212 GND 0.476712f
C4905 VOUT.t40 GND 0.049715f
C4906 VOUT.t28 GND 0.049715f
C4907 VOUT.n213 GND 0.384224f
C4908 VOUT.n214 GND 0.235858f
C4909 VOUT.t52 GND 0.049715f
C4910 VOUT.t13 GND 0.049715f
C4911 VOUT.n215 GND 0.384224f
C4912 VOUT.n216 GND 0.235858f
C4913 VOUT.t2 GND 0.049715f
C4914 VOUT.t15 GND 0.049715f
C4915 VOUT.n217 GND 0.384224f
C4916 VOUT.n218 GND 0.235858f
C4917 VOUT.t62 GND 0.049715f
C4918 VOUT.t0 GND 0.049715f
C4919 VOUT.n219 GND 0.384222f
C4920 VOUT.n220 GND 0.327357f
C4921 VOUT.n221 GND 0.600494f
C4922 VOUT.n222 GND 10.1415f
C4923 VOUT.t111 GND 0.043501f
C4924 VOUT.t93 GND 0.043501f
C4925 VOUT.n223 GND 0.3877f
C4926 VOUT.t91 GND 0.043501f
C4927 VOUT.t92 GND 0.043501f
C4928 VOUT.n224 GND 0.384387f
C4929 VOUT.n225 GND 0.530906f
C4930 VOUT.t74 GND 0.043501f
C4931 VOUT.t72 GND 0.043501f
C4932 VOUT.n226 GND 0.384387f
C4933 VOUT.n227 GND 0.263942f
C4934 VOUT.t85 GND 0.043501f
C4935 VOUT.t83 GND 0.043501f
C4936 VOUT.n228 GND 0.384387f
C4937 VOUT.n229 GND 0.263942f
C4938 VOUT.t96 GND 0.043501f
C4939 VOUT.t95 GND 0.043501f
C4940 VOUT.n230 GND 0.384387f
C4941 VOUT.n231 GND 0.416694f
C4942 VOUT.t94 GND 0.043501f
C4943 VOUT.t76 GND 0.043501f
C4944 VOUT.n232 GND 0.3877f
C4945 VOUT.t73 GND 0.043501f
C4946 VOUT.t77 GND 0.043501f
C4947 VOUT.n233 GND 0.384387f
C4948 VOUT.n234 GND 0.530906f
C4949 VOUT.t100 GND 0.043501f
C4950 VOUT.t98 GND 0.043501f
C4951 VOUT.n235 GND 0.384387f
C4952 VOUT.n236 GND 0.263942f
C4953 VOUT.t109 GND 0.043501f
C4954 VOUT.t106 GND 0.043501f
C4955 VOUT.n237 GND 0.384387f
C4956 VOUT.n238 GND 0.263942f
C4957 VOUT.t79 GND 0.043501f
C4958 VOUT.t78 GND 0.043501f
C4959 VOUT.n239 GND 0.384387f
C4960 VOUT.n240 GND 0.348682f
C4961 VOUT.n241 GND 0.88321f
C4962 VOUT.n242 GND 10.3764f
C4963 VOUT.t103 GND 0.043501f
C4964 VOUT.t97 GND 0.043501f
C4965 VOUT.n243 GND 0.3877f
C4966 VOUT.t104 GND 0.043501f
C4967 VOUT.t75 GND 0.043501f
C4968 VOUT.n244 GND 0.384387f
C4969 VOUT.n245 GND 0.530906f
C4970 VOUT.t84 GND 0.043501f
C4971 VOUT.t86 GND 0.043501f
C4972 VOUT.n246 GND 0.384387f
C4973 VOUT.n247 GND 0.263942f
C4974 VOUT.t108 GND 0.043501f
C4975 VOUT.t99 GND 0.043501f
C4976 VOUT.n248 GND 0.384387f
C4977 VOUT.n249 GND 0.263942f
C4978 VOUT.t81 GND 0.043501f
C4979 VOUT.t105 GND 0.043501f
C4980 VOUT.n250 GND 0.384387f
C4981 VOUT.n251 GND 0.416694f
C4982 VOUT.t87 GND 0.043501f
C4983 VOUT.t80 GND 0.043501f
C4984 VOUT.n252 GND 0.3877f
C4985 VOUT.t88 GND 0.043501f
C4986 VOUT.t101 GND 0.043501f
C4987 VOUT.n253 GND 0.384387f
C4988 VOUT.n254 GND 0.530906f
C4989 VOUT.t107 GND 0.043501f
C4990 VOUT.t110 GND 0.043501f
C4991 VOUT.n255 GND 0.384387f
C4992 VOUT.n256 GND 0.263942f
C4993 VOUT.t90 GND 0.043501f
C4994 VOUT.t82 GND 0.043501f
C4995 VOUT.n257 GND 0.384387f
C4996 VOUT.n258 GND 0.263942f
C4997 VOUT.t102 GND 0.043501f
C4998 VOUT.t89 GND 0.043501f
C4999 VOUT.n259 GND 0.384387f
C5000 VOUT.n260 GND 0.348682f
C5001 VOUT.n261 GND 0.88321f
C5002 VOUT.n262 GND 6.35633f
C5003 VOUT.n263 GND 7.11697f
C5004 a_n8209_7799.n0 GND 0.676161f
C5005 a_n8209_7799.n1 GND 0.04032f
C5006 a_n8209_7799.n2 GND 0.676161f
C5007 a_n8209_7799.n3 GND 0.04032f
C5008 a_n8209_7799.n4 GND 0.676161f
C5009 a_n8209_7799.n5 GND 0.04032f
C5010 a_n8209_7799.n6 GND 0.506037f
C5011 a_n8209_7799.n7 GND 0.0382f
C5012 a_n8209_7799.n8 GND 0.5638f
C5013 a_n8209_7799.n9 GND 0.40251f
C5014 a_n8209_7799.n10 GND 0.5638f
C5015 a_n8209_7799.n11 GND 0.40251f
C5016 a_n8209_7799.n12 GND 0.337358f
C5017 a_n8209_7799.n13 GND 0.0382f
C5018 a_n8209_7799.n14 GND 0.337358f
C5019 a_n8209_7799.n15 GND 0.0382f
C5020 a_n8209_7799.n16 GND 0.337358f
C5021 a_n8209_7799.n17 GND 0.0382f
C5022 a_n8209_7799.n18 GND 0.465312f
C5023 a_n8209_7799.n19 GND 0.04032f
C5024 a_n8209_7799.n20 GND 0.337358f
C5025 a_n8209_7799.n21 GND 0.040328f
C5026 a_n8209_7799.n22 GND 0.04032f
C5027 a_n8209_7799.n23 GND 0.465312f
C5028 a_n8209_7799.n24 GND 0.04032f
C5029 a_n8209_7799.n25 GND 0.337358f
C5030 a_n8209_7799.n26 GND 0.040328f
C5031 a_n8209_7799.n27 GND 0.04032f
C5032 a_n8209_7799.n28 GND 0.465312f
C5033 a_n8209_7799.n29 GND 0.04032f
C5034 a_n8209_7799.n30 GND 0.040328f
C5035 a_n8209_7799.n31 GND 0.352951f
C5036 a_n8209_7799.n32 GND 0.40251f
C5037 a_n8209_7799.n33 GND 0.352951f
C5038 a_n8209_7799.n34 GND 0.40251f
C5039 a_n8209_7799.n35 GND 0.490143f
C5040 a_n8209_7799.n36 GND 0.40251f
C5041 a_n8209_7799.n37 GND 0.049472f
C5042 a_n8209_7799.n38 GND 0.049654f
C5043 a_n8209_7799.n39 GND 0.0382f
C5044 a_n8209_7799.n40 GND 0.049472f
C5045 a_n8209_7799.n41 GND 0.049654f
C5046 a_n8209_7799.n42 GND 0.0382f
C5047 a_n8209_7799.n43 GND 0.049472f
C5048 a_n8209_7799.n44 GND 0.049654f
C5049 a_n8209_7799.n45 GND 0.0382f
C5050 a_n8209_7799.n46 GND 0.049472f
C5051 a_n8209_7799.n47 GND 0.049654f
C5052 a_n8209_7799.n48 GND 0.0382f
C5053 a_n8209_7799.n49 GND 0.049472f
C5054 a_n8209_7799.n50 GND 0.049654f
C5055 a_n8209_7799.n51 GND 0.0382f
C5056 a_n8209_7799.n52 GND 0.049472f
C5057 a_n8209_7799.n53 GND 0.049654f
C5058 a_n8209_7799.n54 GND 0.04172f
C5059 a_n8209_7799.n55 GND 0.041439f
C5060 a_n8209_7799.n56 GND 0.049472f
C5061 a_n8209_7799.n57 GND 0.049654f
C5062 a_n8209_7799.n58 GND 0.04172f
C5063 a_n8209_7799.n59 GND 0.041439f
C5064 a_n8209_7799.n60 GND 0.049472f
C5065 a_n8209_7799.n61 GND 0.049654f
C5066 a_n8209_7799.n62 GND 0.04172f
C5067 a_n8209_7799.n63 GND 0.041439f
C5068 a_n8209_7799.n64 GND 0.049472f
C5069 a_n8209_7799.n65 GND 0.049654f
C5070 a_n8209_7799.n66 GND 0.049022f
C5071 a_n8209_7799.n67 GND 0.049472f
C5072 a_n8209_7799.n68 GND 0.049654f
C5073 a_n8209_7799.n69 GND 0.049022f
C5074 a_n8209_7799.n70 GND 0.049472f
C5075 a_n8209_7799.n71 GND 0.049654f
C5076 a_n8209_7799.n72 GND 0.049022f
C5077 a_n8209_7799.n73 GND 0.049472f
C5078 a_n8209_7799.n74 GND 0.084339f
C5079 a_n8209_7799.n75 GND 0.084339f
C5080 a_n8209_7799.n76 GND 0.041185f
C5081 a_n8209_7799.n77 GND 0.049654f
C5082 a_n8209_7799.n78 GND 0.09844f
C5083 a_n8209_7799.n79 GND 0.037513f
C5084 a_n8209_7799.t16 GND 0.077998f
C5085 a_n8209_7799.t13 GND 0.077998f
C5086 a_n8209_7799.t10 GND 0.077998f
C5087 a_n8209_7799.n80 GND 0.563586f
C5088 a_n8209_7799.t18 GND 0.077998f
C5089 a_n8209_7799.t2 GND 0.077998f
C5090 a_n8209_7799.n81 GND 0.560966f
C5091 a_n8209_7799.n82 GND 0.988196f
C5092 a_n8209_7799.t12 GND 0.077998f
C5093 a_n8209_7799.t17 GND 0.077998f
C5094 a_n8209_7799.n83 GND 0.560966f
C5095 a_n8209_7799.n84 GND 2.2129f
C5096 a_n8209_7799.t5 GND 0.077998f
C5097 a_n8209_7799.t0 GND 0.077998f
C5098 a_n8209_7799.n85 GND 0.563588f
C5099 a_n8209_7799.t6 GND 0.077998f
C5100 a_n8209_7799.t11 GND 0.077998f
C5101 a_n8209_7799.n86 GND 0.560966f
C5102 a_n8209_7799.n87 GND 0.988193f
C5103 a_n8209_7799.t7 GND 0.077998f
C5104 a_n8209_7799.t19 GND 0.077998f
C5105 a_n8209_7799.n88 GND 0.560966f
C5106 a_n8209_7799.n89 GND 1.52644f
C5107 a_n8209_7799.n90 GND 4.74367f
C5108 a_n8209_7799.t89 GND 0.906042f
C5109 a_n8209_7799.n91 GND 0.42016f
C5110 a_n8209_7799.t67 GND 0.906042f
C5111 a_n8209_7799.t85 GND 0.906042f
C5112 a_n8209_7799.t52 GND 0.906042f
C5113 a_n8209_7799.t87 GND 0.906042f
C5114 a_n8209_7799.t66 GND 0.906042f
C5115 a_n8209_7799.n92 GND 0.379389f
C5116 a_n8209_7799.t32 GND 0.906042f
C5117 a_n8209_7799.n93 GND 0.442425f
C5118 a_n8209_7799.t71 GND 0.906042f
C5119 a_n8209_7799.n94 GND 0.442404f
C5120 a_n8209_7799.t49 GND 0.906042f
C5121 a_n8209_7799.t34 GND 1.0071f
C5122 a_n8209_7799.n95 GND 0.404292f
C5123 a_n8209_7799.n96 GND 0.443169f
C5124 a_n8209_7799.n97 GND 0.065188f
C5125 a_n8209_7799.n98 GND 0.442485f
C5126 a_n8209_7799.n99 GND 0.442485f
C5127 a_n8209_7799.t74 GND 0.906042f
C5128 a_n8209_7799.n100 GND 0.444016f
C5129 a_n8209_7799.n101 GND 0.399993f
C5130 a_n8209_7799.n102 GND 0.067999f
C5131 a_n8209_7799.n103 GND 0.427356f
C5132 a_n8209_7799.t25 GND 0.970253f
C5133 a_n8209_7799.n104 GND 0.424702f
C5134 a_n8209_7799.n105 GND 0.265193f
C5135 a_n8209_7799.t27 GND 0.906042f
C5136 a_n8209_7799.n106 GND 0.443181f
C5137 a_n8209_7799.t75 GND 0.906042f
C5138 a_n8209_7799.t22 GND 0.906042f
C5139 a_n8209_7799.t60 GND 0.906042f
C5140 a_n8209_7799.t24 GND 0.906042f
C5141 a_n8209_7799.t72 GND 0.906042f
C5142 a_n8209_7799.n107 GND 0.379389f
C5143 a_n8209_7799.t41 GND 0.906042f
C5144 a_n8209_7799.n108 GND 0.442425f
C5145 a_n8209_7799.t80 GND 0.906042f
C5146 a_n8209_7799.n109 GND 0.442404f
C5147 a_n8209_7799.t59 GND 0.906042f
C5148 a_n8209_7799.t42 GND 1.0071f
C5149 a_n8209_7799.n110 GND 0.404292f
C5150 a_n8209_7799.n111 GND 0.443169f
C5151 a_n8209_7799.n112 GND 0.065188f
C5152 a_n8209_7799.n113 GND 0.442485f
C5153 a_n8209_7799.n114 GND 0.442485f
C5154 a_n8209_7799.t81 GND 0.906042f
C5155 a_n8209_7799.n115 GND 0.444016f
C5156 a_n8209_7799.n116 GND 0.453809f
C5157 a_n8209_7799.n117 GND 0.442404f
C5158 a_n8209_7799.t36 GND 1.00694f
C5159 a_n8209_7799.n118 GND 0.745335f
C5160 a_n8209_7799.t45 GND 0.906042f
C5161 a_n8209_7799.n119 GND 0.443181f
C5162 a_n8209_7799.t62 GND 0.906042f
C5163 a_n8209_7799.t86 GND 0.906042f
C5164 a_n8209_7799.t55 GND 0.906042f
C5165 a_n8209_7799.t65 GND 0.906042f
C5166 a_n8209_7799.t79 GND 0.906042f
C5167 a_n8209_7799.n120 GND 0.379389f
C5168 a_n8209_7799.t46 GND 0.906042f
C5169 a_n8209_7799.n121 GND 0.442425f
C5170 a_n8209_7799.t61 GND 0.906042f
C5171 a_n8209_7799.n122 GND 0.442404f
C5172 a_n8209_7799.t70 GND 0.906042f
C5173 a_n8209_7799.t88 GND 1.0071f
C5174 a_n8209_7799.n123 GND 0.404292f
C5175 a_n8209_7799.n124 GND 0.443169f
C5176 a_n8209_7799.n125 GND 0.065188f
C5177 a_n8209_7799.n126 GND 0.442485f
C5178 a_n8209_7799.n127 GND 0.442485f
C5179 a_n8209_7799.t38 GND 0.906042f
C5180 a_n8209_7799.n128 GND 0.444016f
C5181 a_n8209_7799.n129 GND 0.453809f
C5182 a_n8209_7799.n130 GND 0.442404f
C5183 a_n8209_7799.t53 GND 1.00694f
C5184 a_n8209_7799.n131 GND 1.24603f
C5185 a_n8209_7799.t48 GND 1.00694f
C5186 a_n8209_7799.t40 GND 0.906042f
C5187 a_n8209_7799.n132 GND 0.443181f
C5188 a_n8209_7799.t84 GND 0.906042f
C5189 a_n8209_7799.t30 GND 0.906042f
C5190 a_n8209_7799.t20 GND 0.906042f
C5191 a_n8209_7799.n133 GND 0.444016f
C5192 a_n8209_7799.t69 GND 0.906042f
C5193 a_n8209_7799.t39 GND 0.906042f
C5194 a_n8209_7799.t77 GND 0.906042f
C5195 a_n8209_7799.n134 GND 0.444016f
C5196 a_n8209_7799.t54 GND 0.906042f
C5197 a_n8209_7799.n135 GND 0.453809f
C5198 a_n8209_7799.t91 GND 0.906042f
C5199 a_n8209_7799.n136 GND 0.442404f
C5200 a_n8209_7799.t68 GND 0.906042f
C5201 a_n8209_7799.t56 GND 1.0071f
C5202 a_n8209_7799.n137 GND 0.404292f
C5203 a_n8209_7799.n138 GND 0.443169f
C5204 a_n8209_7799.n139 GND 0.427765f
C5205 a_n8209_7799.n140 GND 0.06798f
C5206 a_n8209_7799.n141 GND 0.388114f
C5207 a_n8209_7799.n142 GND 0.439397f
C5208 a_n8209_7799.n143 GND 0.067946f
C5209 a_n8209_7799.n144 GND 0.387471f
C5210 a_n8209_7799.t57 GND 1.00694f
C5211 a_n8209_7799.t50 GND 0.906042f
C5212 a_n8209_7799.n145 GND 0.443181f
C5213 a_n8209_7799.t21 GND 0.906042f
C5214 a_n8209_7799.t37 GND 0.906042f
C5215 a_n8209_7799.t31 GND 0.906042f
C5216 a_n8209_7799.n146 GND 0.444016f
C5217 a_n8209_7799.t78 GND 0.906042f
C5218 a_n8209_7799.t47 GND 0.906042f
C5219 a_n8209_7799.t82 GND 0.906042f
C5220 a_n8209_7799.n147 GND 0.444016f
C5221 a_n8209_7799.t63 GND 0.906042f
C5222 a_n8209_7799.n148 GND 0.453809f
C5223 a_n8209_7799.t29 GND 0.906042f
C5224 a_n8209_7799.n149 GND 0.442404f
C5225 a_n8209_7799.t76 GND 0.906042f
C5226 a_n8209_7799.t64 GND 1.0071f
C5227 a_n8209_7799.n150 GND 0.404292f
C5228 a_n8209_7799.n151 GND 0.443169f
C5229 a_n8209_7799.n152 GND 0.427765f
C5230 a_n8209_7799.n153 GND 0.06798f
C5231 a_n8209_7799.n154 GND 0.388114f
C5232 a_n8209_7799.n155 GND 0.439397f
C5233 a_n8209_7799.n156 GND 0.067946f
C5234 a_n8209_7799.n157 GND 0.387471f
C5235 a_n8209_7799.n158 GND 0.745335f
C5236 a_n8209_7799.t33 GND 1.00694f
C5237 a_n8209_7799.t26 GND 0.906042f
C5238 a_n8209_7799.n159 GND 0.443181f
C5239 a_n8209_7799.t44 GND 0.906042f
C5240 a_n8209_7799.t23 GND 0.906042f
C5241 a_n8209_7799.t90 GND 0.906042f
C5242 a_n8209_7799.n160 GND 0.444016f
C5243 a_n8209_7799.t35 GND 0.906042f
C5244 a_n8209_7799.t51 GND 0.906042f
C5245 a_n8209_7799.t83 GND 0.906042f
C5246 a_n8209_7799.n161 GND 0.444016f
C5247 a_n8209_7799.t28 GND 0.906042f
C5248 a_n8209_7799.n162 GND 0.453809f
C5249 a_n8209_7799.t43 GND 0.906042f
C5250 a_n8209_7799.n163 GND 0.442404f
C5251 a_n8209_7799.t58 GND 0.906042f
C5252 a_n8209_7799.t73 GND 1.0071f
C5253 a_n8209_7799.n164 GND 0.404292f
C5254 a_n8209_7799.n165 GND 0.443169f
C5255 a_n8209_7799.n166 GND 0.427765f
C5256 a_n8209_7799.n167 GND 0.06798f
C5257 a_n8209_7799.n168 GND 0.388114f
C5258 a_n8209_7799.n169 GND 0.439397f
C5259 a_n8209_7799.n170 GND 0.067946f
C5260 a_n8209_7799.n171 GND 0.387471f
C5261 a_n8209_7799.n172 GND 1.03812f
C5262 a_n8209_7799.n173 GND 11.029f
C5263 a_n8209_7799.n174 GND 3.6885f
C5264 a_n8209_7799.t15 GND 0.077998f
C5265 a_n8209_7799.t3 GND 0.077998f
C5266 a_n8209_7799.n175 GND 0.682285f
C5267 a_n8209_7799.n176 GND 0.733606f
C5268 a_n8209_7799.t14 GND 0.077998f
C5269 a_n8209_7799.t9 GND 0.077998f
C5270 a_n8209_7799.n177 GND 0.681194f
C5271 a_n8209_7799.n178 GND 1.89394f
C5272 a_n8209_7799.t8 GND 0.077998f
C5273 a_n8209_7799.t4 GND 0.077998f
C5274 a_n8209_7799.n179 GND 0.682283f
C5275 a_n8209_7799.n180 GND 2.0167f
C5276 a_n8209_7799.n181 GND 0.682282f
C5277 a_n8209_7799.t1 GND 0.077998f
C5278 CS_BIAS.n0 GND 0.007821f
C5279 CS_BIAS.t40 GND 0.221674f
C5280 CS_BIAS.n1 GND 0.009773f
C5281 CS_BIAS.n2 GND 0.005932f
C5282 CS_BIAS.t58 GND 0.221674f
C5283 CS_BIAS.n3 GND 0.004799f
C5284 CS_BIAS.n4 GND 0.005932f
C5285 CS_BIAS.t60 GND 0.221674f
C5286 CS_BIAS.n5 GND 0.010086f
C5287 CS_BIAS.n6 GND 0.005932f
C5288 CS_BIAS.t59 GND 0.221674f
C5289 CS_BIAS.n7 GND 0.083017f
C5290 CS_BIAS.n8 GND 0.005932f
C5291 CS_BIAS.n9 GND 0.009209f
C5292 CS_BIAS.n10 GND 0.005904f
C5293 CS_BIAS.t77 GND 0.221674f
C5294 CS_BIAS.n11 GND 0.083017f
C5295 CS_BIAS.n12 GND 0.011729f
C5296 CS_BIAS.n13 GND 0.007821f
C5297 CS_BIAS.t32 GND 0.221674f
C5298 CS_BIAS.n14 GND 0.009773f
C5299 CS_BIAS.n15 GND 0.005932f
C5300 CS_BIAS.t26 GND 0.221674f
C5301 CS_BIAS.n16 GND 0.004799f
C5302 CS_BIAS.n17 GND 0.005932f
C5303 CS_BIAS.t0 GND 0.221674f
C5304 CS_BIAS.n18 GND 0.010086f
C5305 CS_BIAS.n19 GND 0.005932f
C5306 CS_BIAS.t38 GND 0.221674f
C5307 CS_BIAS.n20 GND 0.083017f
C5308 CS_BIAS.n21 GND 0.005932f
C5309 CS_BIAS.n22 GND 0.009209f
C5310 CS_BIAS.n23 GND 0.005932f
C5311 CS_BIAS.t34 GND 0.221674f
C5312 CS_BIAS.n24 GND 0.083017f
C5313 CS_BIAS.n25 GND 0.011729f
C5314 CS_BIAS.n26 GND 0.005932f
C5315 CS_BIAS.t36 GND 0.221674f
C5316 CS_BIAS.n27 GND 0.007311f
C5317 CS_BIAS.n28 GND 0.005932f
C5318 CS_BIAS.t28 GND 0.221674f
C5319 CS_BIAS.n29 GND 0.007058f
C5320 CS_BIAS.n30 GND 0.005932f
C5321 CS_BIAS.t24 GND 0.221674f
C5322 CS_BIAS.n31 GND 0.011666f
C5323 CS_BIAS.n32 GND 0.005932f
C5324 CS_BIAS.t4 GND 0.221674f
C5325 CS_BIAS.n33 GND 0.096202f
C5326 CS_BIAS.t12 GND 0.252039f
C5327 CS_BIAS.n34 GND 0.097593f
C5328 CS_BIAS.n35 GND 0.044363f
C5329 CS_BIAS.n36 GND 0.007254f
C5330 CS_BIAS.n37 GND 0.011784f
C5331 CS_BIAS.n38 GND 0.004799f
C5332 CS_BIAS.n39 GND 0.005932f
C5333 CS_BIAS.n40 GND 0.005932f
C5334 CS_BIAS.n41 GND 0.005932f
C5335 CS_BIAS.n42 GND 0.007471f
C5336 CS_BIAS.n43 GND 0.083017f
C5337 CS_BIAS.n44 GND 0.0091f
C5338 CS_BIAS.n45 GND 0.010086f
C5339 CS_BIAS.n46 GND 0.005932f
C5340 CS_BIAS.n47 GND 0.005932f
C5341 CS_BIAS.n48 GND 0.005932f
C5342 CS_BIAS.n49 GND 0.011104f
C5343 CS_BIAS.n50 GND 0.005625f
C5344 CS_BIAS.n51 GND 0.083017f
C5345 CS_BIAS.n52 GND 0.010947f
C5346 CS_BIAS.n53 GND 0.005932f
C5347 CS_BIAS.n54 GND 0.005932f
C5348 CS_BIAS.n55 GND 0.005932f
C5349 CS_BIAS.n56 GND 0.009937f
C5350 CS_BIAS.n57 GND 0.009209f
C5351 CS_BIAS.n58 GND 0.083017f
C5352 CS_BIAS.n59 GND 0.007362f
C5353 CS_BIAS.n60 GND 0.005932f
C5354 CS_BIAS.n61 GND 0.005932f
C5355 CS_BIAS.n62 GND 0.005932f
C5356 CS_BIAS.n63 GND 0.004791f
C5357 CS_BIAS.n64 GND 0.011729f
C5358 CS_BIAS.n65 GND 0.007362f
C5359 CS_BIAS.n66 GND 0.005932f
C5360 CS_BIAS.n67 GND 0.005932f
C5361 CS_BIAS.n68 GND 0.005932f
C5362 CS_BIAS.n69 GND 0.009937f
C5363 CS_BIAS.n70 GND 0.007311f
C5364 CS_BIAS.n71 GND 0.010947f
C5365 CS_BIAS.n72 GND 0.005932f
C5366 CS_BIAS.n73 GND 0.005932f
C5367 CS_BIAS.n74 GND 0.005625f
C5368 CS_BIAS.n75 GND 0.011104f
C5369 CS_BIAS.n76 GND 0.007058f
C5370 CS_BIAS.n77 GND 0.005932f
C5371 CS_BIAS.n78 GND 0.005932f
C5372 CS_BIAS.n79 GND 0.005932f
C5373 CS_BIAS.n80 GND 0.0091f
C5374 CS_BIAS.n81 GND 0.083017f
C5375 CS_BIAS.n82 GND 0.007471f
C5376 CS_BIAS.n83 GND 0.011666f
C5377 CS_BIAS.n84 GND 0.005932f
C5378 CS_BIAS.n85 GND 0.005932f
C5379 CS_BIAS.n86 GND 0.005932f
C5380 CS_BIAS.n87 GND 0.011784f
C5381 CS_BIAS.n88 GND 0.007254f
C5382 CS_BIAS.n89 GND 0.083017f
C5383 CS_BIAS.n90 GND 0.009318f
C5384 CS_BIAS.n91 GND 0.005932f
C5385 CS_BIAS.n92 GND 0.005932f
C5386 CS_BIAS.n93 GND 0.005932f
C5387 CS_BIAS.n94 GND 0.007475f
C5388 CS_BIAS.n95 GND 0.010838f
C5389 CS_BIAS.n96 GND 0.102559f
C5390 CS_BIAS.n97 GND 0.063147f
C5391 CS_BIAS.t33 GND 0.012802f
C5392 CS_BIAS.t27 GND 0.012802f
C5393 CS_BIAS.n98 GND 0.11312f
C5394 CS_BIAS.n99 GND 0.122649f
C5395 CS_BIAS.t1 GND 0.012802f
C5396 CS_BIAS.t39 GND 0.012802f
C5397 CS_BIAS.n100 GND 0.11312f
C5398 CS_BIAS.n101 GND 0.077675f
C5399 CS_BIAS.t35 GND 0.012802f
C5400 CS_BIAS.t37 GND 0.012802f
C5401 CS_BIAS.n102 GND 0.11312f
C5402 CS_BIAS.t5 GND 0.012802f
C5403 CS_BIAS.t13 GND 0.012802f
C5404 CS_BIAS.n103 GND 0.114095f
C5405 CS_BIAS.t29 GND 0.012802f
C5406 CS_BIAS.t25 GND 0.012802f
C5407 CS_BIAS.n104 GND 0.11312f
C5408 CS_BIAS.n105 GND 0.156239f
C5409 CS_BIAS.n106 GND 0.11314f
C5410 CS_BIAS.n107 GND 0.005932f
C5411 CS_BIAS.t79 GND 0.221674f
C5412 CS_BIAS.n108 GND 0.007311f
C5413 CS_BIAS.n109 GND 0.005932f
C5414 CS_BIAS.t66 GND 0.221674f
C5415 CS_BIAS.n110 GND 0.007058f
C5416 CS_BIAS.n111 GND 0.005932f
C5417 CS_BIAS.t68 GND 0.221674f
C5418 CS_BIAS.n112 GND 0.011666f
C5419 CS_BIAS.n113 GND 0.005932f
C5420 CS_BIAS.t55 GND 0.221674f
C5421 CS_BIAS.n114 GND 0.096202f
C5422 CS_BIAS.t56 GND 0.252039f
C5423 CS_BIAS.n115 GND 0.097593f
C5424 CS_BIAS.n116 GND 0.044363f
C5425 CS_BIAS.n117 GND 0.007254f
C5426 CS_BIAS.n118 GND 0.011784f
C5427 CS_BIAS.n119 GND 0.004799f
C5428 CS_BIAS.n120 GND 0.005932f
C5429 CS_BIAS.n121 GND 0.005932f
C5430 CS_BIAS.n122 GND 0.005932f
C5431 CS_BIAS.n123 GND 0.007471f
C5432 CS_BIAS.n124 GND 0.083017f
C5433 CS_BIAS.n125 GND 0.0091f
C5434 CS_BIAS.n126 GND 0.010086f
C5435 CS_BIAS.n127 GND 0.005932f
C5436 CS_BIAS.n128 GND 0.005932f
C5437 CS_BIAS.n129 GND 0.005932f
C5438 CS_BIAS.n130 GND 0.011104f
C5439 CS_BIAS.n131 GND 0.005625f
C5440 CS_BIAS.n132 GND 0.083017f
C5441 CS_BIAS.n133 GND 0.010947f
C5442 CS_BIAS.n134 GND 0.005932f
C5443 CS_BIAS.n135 GND 0.005932f
C5444 CS_BIAS.n136 GND 0.005932f
C5445 CS_BIAS.n137 GND 0.009937f
C5446 CS_BIAS.n138 GND 0.009209f
C5447 CS_BIAS.n139 GND 0.083017f
C5448 CS_BIAS.n140 GND 0.007362f
C5449 CS_BIAS.n141 GND 0.005932f
C5450 CS_BIAS.n142 GND 0.005904f
C5451 CS_BIAS.n143 GND 0.042885f
C5452 CS_BIAS.n144 GND 0.004791f
C5453 CS_BIAS.n145 GND 0.011729f
C5454 CS_BIAS.n146 GND 0.007362f
C5455 CS_BIAS.n147 GND 0.005932f
C5456 CS_BIAS.n148 GND 0.005932f
C5457 CS_BIAS.n149 GND 0.005932f
C5458 CS_BIAS.n150 GND 0.009937f
C5459 CS_BIAS.n151 GND 0.007311f
C5460 CS_BIAS.n152 GND 0.010947f
C5461 CS_BIAS.n153 GND 0.005932f
C5462 CS_BIAS.n154 GND 0.005932f
C5463 CS_BIAS.n155 GND 0.005625f
C5464 CS_BIAS.n156 GND 0.011104f
C5465 CS_BIAS.n157 GND 0.007058f
C5466 CS_BIAS.n158 GND 0.005932f
C5467 CS_BIAS.n159 GND 0.005932f
C5468 CS_BIAS.n160 GND 0.005932f
C5469 CS_BIAS.n161 GND 0.0091f
C5470 CS_BIAS.n162 GND 0.083017f
C5471 CS_BIAS.n163 GND 0.007471f
C5472 CS_BIAS.n164 GND 0.011666f
C5473 CS_BIAS.n165 GND 0.005932f
C5474 CS_BIAS.n166 GND 0.005932f
C5475 CS_BIAS.n167 GND 0.005932f
C5476 CS_BIAS.n168 GND 0.011784f
C5477 CS_BIAS.n169 GND 0.007254f
C5478 CS_BIAS.n170 GND 0.083017f
C5479 CS_BIAS.n171 GND 0.009318f
C5480 CS_BIAS.n172 GND 0.005932f
C5481 CS_BIAS.n173 GND 0.005932f
C5482 CS_BIAS.n174 GND 0.005932f
C5483 CS_BIAS.n175 GND 0.007475f
C5484 CS_BIAS.n176 GND 0.010838f
C5485 CS_BIAS.n177 GND 0.102559f
C5486 CS_BIAS.n178 GND 0.038082f
C5487 CS_BIAS.n179 GND 0.007821f
C5488 CS_BIAS.t57 GND 0.221674f
C5489 CS_BIAS.n180 GND 0.009773f
C5490 CS_BIAS.n181 GND 0.005932f
C5491 CS_BIAS.t75 GND 0.221674f
C5492 CS_BIAS.n182 GND 0.004799f
C5493 CS_BIAS.n183 GND 0.005932f
C5494 CS_BIAS.t78 GND 0.221674f
C5495 CS_BIAS.n184 GND 0.010086f
C5496 CS_BIAS.n185 GND 0.005932f
C5497 CS_BIAS.t74 GND 0.221674f
C5498 CS_BIAS.n186 GND 0.083017f
C5499 CS_BIAS.n187 GND 0.005932f
C5500 CS_BIAS.n188 GND 0.009209f
C5501 CS_BIAS.n189 GND 0.005932f
C5502 CS_BIAS.t51 GND 0.221674f
C5503 CS_BIAS.n190 GND 0.083017f
C5504 CS_BIAS.n191 GND 0.011729f
C5505 CS_BIAS.n192 GND 0.005932f
C5506 CS_BIAS.t53 GND 0.221674f
C5507 CS_BIAS.n193 GND 0.007311f
C5508 CS_BIAS.n194 GND 0.005932f
C5509 CS_BIAS.t42 GND 0.221674f
C5510 CS_BIAS.n195 GND 0.007058f
C5511 CS_BIAS.n196 GND 0.005932f
C5512 CS_BIAS.t45 GND 0.221674f
C5513 CS_BIAS.n197 GND 0.011666f
C5514 CS_BIAS.n198 GND 0.005932f
C5515 CS_BIAS.t72 GND 0.221674f
C5516 CS_BIAS.n199 GND 0.096202f
C5517 CS_BIAS.t73 GND 0.252039f
C5518 CS_BIAS.n200 GND 0.097593f
C5519 CS_BIAS.n201 GND 0.044363f
C5520 CS_BIAS.n202 GND 0.007254f
C5521 CS_BIAS.n203 GND 0.011784f
C5522 CS_BIAS.n204 GND 0.004799f
C5523 CS_BIAS.n205 GND 0.005932f
C5524 CS_BIAS.n206 GND 0.005932f
C5525 CS_BIAS.n207 GND 0.005932f
C5526 CS_BIAS.n208 GND 0.007471f
C5527 CS_BIAS.n209 GND 0.083017f
C5528 CS_BIAS.n210 GND 0.0091f
C5529 CS_BIAS.n211 GND 0.010086f
C5530 CS_BIAS.n212 GND 0.005932f
C5531 CS_BIAS.n213 GND 0.005932f
C5532 CS_BIAS.n214 GND 0.005932f
C5533 CS_BIAS.n215 GND 0.011104f
C5534 CS_BIAS.n216 GND 0.005625f
C5535 CS_BIAS.n217 GND 0.083017f
C5536 CS_BIAS.n218 GND 0.010947f
C5537 CS_BIAS.n219 GND 0.005932f
C5538 CS_BIAS.n220 GND 0.005932f
C5539 CS_BIAS.n221 GND 0.005932f
C5540 CS_BIAS.n222 GND 0.009937f
C5541 CS_BIAS.n223 GND 0.009209f
C5542 CS_BIAS.n224 GND 0.083017f
C5543 CS_BIAS.n225 GND 0.007362f
C5544 CS_BIAS.n226 GND 0.005932f
C5545 CS_BIAS.n227 GND 0.005932f
C5546 CS_BIAS.n228 GND 0.005932f
C5547 CS_BIAS.n229 GND 0.004791f
C5548 CS_BIAS.n230 GND 0.011729f
C5549 CS_BIAS.n231 GND 0.007362f
C5550 CS_BIAS.n232 GND 0.005932f
C5551 CS_BIAS.n233 GND 0.005932f
C5552 CS_BIAS.n234 GND 0.005932f
C5553 CS_BIAS.n235 GND 0.009937f
C5554 CS_BIAS.n236 GND 0.007311f
C5555 CS_BIAS.n237 GND 0.010947f
C5556 CS_BIAS.n238 GND 0.005932f
C5557 CS_BIAS.n239 GND 0.005932f
C5558 CS_BIAS.n240 GND 0.005625f
C5559 CS_BIAS.n241 GND 0.011104f
C5560 CS_BIAS.n242 GND 0.007058f
C5561 CS_BIAS.n243 GND 0.005932f
C5562 CS_BIAS.n244 GND 0.005932f
C5563 CS_BIAS.n245 GND 0.005932f
C5564 CS_BIAS.n246 GND 0.0091f
C5565 CS_BIAS.n247 GND 0.083017f
C5566 CS_BIAS.n248 GND 0.007471f
C5567 CS_BIAS.n249 GND 0.011666f
C5568 CS_BIAS.n250 GND 0.005932f
C5569 CS_BIAS.n251 GND 0.005932f
C5570 CS_BIAS.n252 GND 0.005932f
C5571 CS_BIAS.n253 GND 0.011784f
C5572 CS_BIAS.n254 GND 0.007254f
C5573 CS_BIAS.n255 GND 0.083017f
C5574 CS_BIAS.n256 GND 0.009318f
C5575 CS_BIAS.n257 GND 0.005932f
C5576 CS_BIAS.n258 GND 0.005932f
C5577 CS_BIAS.n259 GND 0.005932f
C5578 CS_BIAS.n260 GND 0.007475f
C5579 CS_BIAS.n261 GND 0.010838f
C5580 CS_BIAS.n262 GND 0.102559f
C5581 CS_BIAS.n263 GND 0.021424f
C5582 CS_BIAS.n264 GND 0.273162f
C5583 CS_BIAS.n265 GND 0.007821f
C5584 CS_BIAS.t54 GND 0.221674f
C5585 CS_BIAS.n266 GND 0.009773f
C5586 CS_BIAS.n267 GND 0.005932f
C5587 CS_BIAS.t48 GND 0.221674f
C5588 CS_BIAS.n268 GND 0.004799f
C5589 CS_BIAS.n269 GND 0.005932f
C5590 CS_BIAS.t76 GND 0.221674f
C5591 CS_BIAS.n270 GND 0.010086f
C5592 CS_BIAS.n271 GND 0.005932f
C5593 CS_BIAS.t47 GND 0.221674f
C5594 CS_BIAS.n272 GND 0.083017f
C5595 CS_BIAS.n273 GND 0.005932f
C5596 CS_BIAS.n274 GND 0.009209f
C5597 CS_BIAS.n275 GND 0.005904f
C5598 CS_BIAS.n276 GND 0.011729f
C5599 CS_BIAS.n277 GND 0.005932f
C5600 CS_BIAS.t67 GND 0.221674f
C5601 CS_BIAS.n278 GND 0.007311f
C5602 CS_BIAS.n279 GND 0.005932f
C5603 CS_BIAS.t52 GND 0.221674f
C5604 CS_BIAS.n280 GND 0.007058f
C5605 CS_BIAS.n281 GND 0.005932f
C5606 CS_BIAS.t43 GND 0.221674f
C5607 CS_BIAS.n282 GND 0.011666f
C5608 CS_BIAS.n283 GND 0.005932f
C5609 CS_BIAS.t46 GND 0.221674f
C5610 CS_BIAS.n284 GND 0.096202f
C5611 CS_BIAS.t70 GND 0.252039f
C5612 CS_BIAS.n285 GND 0.097593f
C5613 CS_BIAS.n286 GND 0.044363f
C5614 CS_BIAS.n287 GND 0.007254f
C5615 CS_BIAS.n288 GND 0.011784f
C5616 CS_BIAS.n289 GND 0.004799f
C5617 CS_BIAS.n290 GND 0.005932f
C5618 CS_BIAS.n291 GND 0.005932f
C5619 CS_BIAS.n292 GND 0.005932f
C5620 CS_BIAS.n293 GND 0.007471f
C5621 CS_BIAS.n294 GND 0.083017f
C5622 CS_BIAS.n295 GND 0.0091f
C5623 CS_BIAS.n296 GND 0.010086f
C5624 CS_BIAS.n297 GND 0.005932f
C5625 CS_BIAS.n298 GND 0.005932f
C5626 CS_BIAS.n299 GND 0.005932f
C5627 CS_BIAS.n300 GND 0.011104f
C5628 CS_BIAS.n301 GND 0.005625f
C5629 CS_BIAS.n302 GND 0.083017f
C5630 CS_BIAS.n303 GND 0.010947f
C5631 CS_BIAS.n304 GND 0.005932f
C5632 CS_BIAS.n305 GND 0.005932f
C5633 CS_BIAS.n306 GND 0.005932f
C5634 CS_BIAS.n307 GND 0.009937f
C5635 CS_BIAS.n308 GND 0.009209f
C5636 CS_BIAS.n309 GND 0.083017f
C5637 CS_BIAS.n310 GND 0.007362f
C5638 CS_BIAS.n311 GND 0.005932f
C5639 CS_BIAS.n312 GND 0.005904f
C5640 CS_BIAS.t11 GND 0.012802f
C5641 CS_BIAS.t7 GND 0.012802f
C5642 CS_BIAS.n313 GND 0.114095f
C5643 CS_BIAS.t3 GND 0.012802f
C5644 CS_BIAS.t23 GND 0.012802f
C5645 CS_BIAS.n314 GND 0.11312f
C5646 CS_BIAS.n315 GND 0.156239f
C5647 CS_BIAS.t15 GND 0.012802f
C5648 CS_BIAS.t9 GND 0.012802f
C5649 CS_BIAS.n316 GND 0.11312f
C5650 CS_BIAS.n317 GND 0.007821f
C5651 CS_BIAS.t30 GND 0.221674f
C5652 CS_BIAS.n318 GND 0.009773f
C5653 CS_BIAS.n319 GND 0.005932f
C5654 CS_BIAS.t20 GND 0.221674f
C5655 CS_BIAS.n320 GND 0.004799f
C5656 CS_BIAS.n321 GND 0.005932f
C5657 CS_BIAS.t18 GND 0.221674f
C5658 CS_BIAS.n322 GND 0.010086f
C5659 CS_BIAS.n323 GND 0.005932f
C5660 CS_BIAS.t16 GND 0.221674f
C5661 CS_BIAS.n324 GND 0.083017f
C5662 CS_BIAS.n325 GND 0.005932f
C5663 CS_BIAS.n326 GND 0.009209f
C5664 CS_BIAS.n327 GND 0.005932f
C5665 CS_BIAS.n328 GND 0.011729f
C5666 CS_BIAS.n329 GND 0.005932f
C5667 CS_BIAS.t14 GND 0.221674f
C5668 CS_BIAS.n330 GND 0.007311f
C5669 CS_BIAS.n331 GND 0.005932f
C5670 CS_BIAS.t22 GND 0.221674f
C5671 CS_BIAS.n332 GND 0.007058f
C5672 CS_BIAS.n333 GND 0.005932f
C5673 CS_BIAS.t2 GND 0.221674f
C5674 CS_BIAS.n334 GND 0.011666f
C5675 CS_BIAS.n335 GND 0.005932f
C5676 CS_BIAS.t6 GND 0.221674f
C5677 CS_BIAS.n336 GND 0.096202f
C5678 CS_BIAS.t10 GND 0.252039f
C5679 CS_BIAS.n337 GND 0.097593f
C5680 CS_BIAS.n338 GND 0.044363f
C5681 CS_BIAS.n339 GND 0.007254f
C5682 CS_BIAS.n340 GND 0.011784f
C5683 CS_BIAS.n341 GND 0.004799f
C5684 CS_BIAS.n342 GND 0.005932f
C5685 CS_BIAS.n343 GND 0.005932f
C5686 CS_BIAS.n344 GND 0.005932f
C5687 CS_BIAS.n345 GND 0.007471f
C5688 CS_BIAS.n346 GND 0.083017f
C5689 CS_BIAS.n347 GND 0.0091f
C5690 CS_BIAS.n348 GND 0.010086f
C5691 CS_BIAS.n349 GND 0.005932f
C5692 CS_BIAS.n350 GND 0.005932f
C5693 CS_BIAS.n351 GND 0.005932f
C5694 CS_BIAS.n352 GND 0.011104f
C5695 CS_BIAS.n353 GND 0.005625f
C5696 CS_BIAS.n354 GND 0.083017f
C5697 CS_BIAS.n355 GND 0.010947f
C5698 CS_BIAS.n356 GND 0.005932f
C5699 CS_BIAS.n357 GND 0.005932f
C5700 CS_BIAS.n358 GND 0.005932f
C5701 CS_BIAS.n359 GND 0.009937f
C5702 CS_BIAS.n360 GND 0.009209f
C5703 CS_BIAS.n361 GND 0.083017f
C5704 CS_BIAS.n362 GND 0.007362f
C5705 CS_BIAS.n363 GND 0.005932f
C5706 CS_BIAS.n364 GND 0.005932f
C5707 CS_BIAS.n365 GND 0.005932f
C5708 CS_BIAS.n366 GND 0.004791f
C5709 CS_BIAS.n367 GND 0.011729f
C5710 CS_BIAS.t8 GND 0.221674f
C5711 CS_BIAS.n368 GND 0.083017f
C5712 CS_BIAS.n369 GND 0.007362f
C5713 CS_BIAS.n370 GND 0.005932f
C5714 CS_BIAS.n371 GND 0.005932f
C5715 CS_BIAS.n372 GND 0.005932f
C5716 CS_BIAS.n373 GND 0.009937f
C5717 CS_BIAS.n374 GND 0.007311f
C5718 CS_BIAS.n375 GND 0.010947f
C5719 CS_BIAS.n376 GND 0.005932f
C5720 CS_BIAS.n377 GND 0.005932f
C5721 CS_BIAS.n378 GND 0.005625f
C5722 CS_BIAS.n379 GND 0.011104f
C5723 CS_BIAS.n380 GND 0.007058f
C5724 CS_BIAS.n381 GND 0.005932f
C5725 CS_BIAS.n382 GND 0.005932f
C5726 CS_BIAS.n383 GND 0.005932f
C5727 CS_BIAS.n384 GND 0.0091f
C5728 CS_BIAS.n385 GND 0.083017f
C5729 CS_BIAS.n386 GND 0.007471f
C5730 CS_BIAS.n387 GND 0.011666f
C5731 CS_BIAS.n388 GND 0.005932f
C5732 CS_BIAS.n389 GND 0.005932f
C5733 CS_BIAS.n390 GND 0.005932f
C5734 CS_BIAS.n391 GND 0.011784f
C5735 CS_BIAS.n392 GND 0.007254f
C5736 CS_BIAS.n393 GND 0.083017f
C5737 CS_BIAS.n394 GND 0.009318f
C5738 CS_BIAS.n395 GND 0.005932f
C5739 CS_BIAS.n396 GND 0.005932f
C5740 CS_BIAS.n397 GND 0.005932f
C5741 CS_BIAS.n398 GND 0.007475f
C5742 CS_BIAS.n399 GND 0.010838f
C5743 CS_BIAS.n400 GND 0.102559f
C5744 CS_BIAS.n401 GND 0.063147f
C5745 CS_BIAS.t21 GND 0.012802f
C5746 CS_BIAS.t31 GND 0.012802f
C5747 CS_BIAS.n402 GND 0.11312f
C5748 CS_BIAS.n403 GND 0.122649f
C5749 CS_BIAS.t17 GND 0.012802f
C5750 CS_BIAS.t19 GND 0.012802f
C5751 CS_BIAS.n404 GND 0.11312f
C5752 CS_BIAS.n405 GND 0.077675f
C5753 CS_BIAS.n406 GND 0.11314f
C5754 CS_BIAS.n407 GND 0.042885f
C5755 CS_BIAS.n408 GND 0.004791f
C5756 CS_BIAS.n409 GND 0.011729f
C5757 CS_BIAS.t65 GND 0.221674f
C5758 CS_BIAS.n410 GND 0.083017f
C5759 CS_BIAS.n411 GND 0.007362f
C5760 CS_BIAS.n412 GND 0.005932f
C5761 CS_BIAS.n413 GND 0.005932f
C5762 CS_BIAS.n414 GND 0.005932f
C5763 CS_BIAS.n415 GND 0.009937f
C5764 CS_BIAS.n416 GND 0.007311f
C5765 CS_BIAS.n417 GND 0.010947f
C5766 CS_BIAS.n418 GND 0.005932f
C5767 CS_BIAS.n419 GND 0.005932f
C5768 CS_BIAS.n420 GND 0.005625f
C5769 CS_BIAS.n421 GND 0.011104f
C5770 CS_BIAS.n422 GND 0.007058f
C5771 CS_BIAS.n423 GND 0.005932f
C5772 CS_BIAS.n424 GND 0.005932f
C5773 CS_BIAS.n425 GND 0.005932f
C5774 CS_BIAS.n426 GND 0.0091f
C5775 CS_BIAS.n427 GND 0.083017f
C5776 CS_BIAS.n428 GND 0.007471f
C5777 CS_BIAS.n429 GND 0.011666f
C5778 CS_BIAS.n430 GND 0.005932f
C5779 CS_BIAS.n431 GND 0.005932f
C5780 CS_BIAS.n432 GND 0.005932f
C5781 CS_BIAS.n433 GND 0.011784f
C5782 CS_BIAS.n434 GND 0.007254f
C5783 CS_BIAS.n435 GND 0.083017f
C5784 CS_BIAS.n436 GND 0.009318f
C5785 CS_BIAS.n437 GND 0.005932f
C5786 CS_BIAS.n438 GND 0.005932f
C5787 CS_BIAS.n439 GND 0.005932f
C5788 CS_BIAS.n440 GND 0.007475f
C5789 CS_BIAS.n441 GND 0.010838f
C5790 CS_BIAS.n442 GND 0.102559f
C5791 CS_BIAS.n443 GND 0.038082f
C5792 CS_BIAS.n444 GND 0.007821f
C5793 CS_BIAS.t71 GND 0.221674f
C5794 CS_BIAS.n445 GND 0.009773f
C5795 CS_BIAS.n446 GND 0.005932f
C5796 CS_BIAS.t64 GND 0.221674f
C5797 CS_BIAS.n447 GND 0.004799f
C5798 CS_BIAS.n448 GND 0.005932f
C5799 CS_BIAS.t50 GND 0.221674f
C5800 CS_BIAS.n449 GND 0.010086f
C5801 CS_BIAS.n450 GND 0.005932f
C5802 CS_BIAS.t63 GND 0.221674f
C5803 CS_BIAS.n451 GND 0.083017f
C5804 CS_BIAS.n452 GND 0.005932f
C5805 CS_BIAS.n453 GND 0.009209f
C5806 CS_BIAS.n454 GND 0.005932f
C5807 CS_BIAS.n455 GND 0.011729f
C5808 CS_BIAS.n456 GND 0.005932f
C5809 CS_BIAS.t44 GND 0.221674f
C5810 CS_BIAS.n457 GND 0.007311f
C5811 CS_BIAS.n458 GND 0.005932f
C5812 CS_BIAS.t69 GND 0.221674f
C5813 CS_BIAS.n459 GND 0.007058f
C5814 CS_BIAS.n460 GND 0.005932f
C5815 CS_BIAS.t61 GND 0.221674f
C5816 CS_BIAS.n461 GND 0.011666f
C5817 CS_BIAS.n462 GND 0.005932f
C5818 CS_BIAS.t62 GND 0.221674f
C5819 CS_BIAS.n463 GND 0.096202f
C5820 CS_BIAS.t49 GND 0.252039f
C5821 CS_BIAS.n464 GND 0.097593f
C5822 CS_BIAS.n465 GND 0.044363f
C5823 CS_BIAS.n466 GND 0.007254f
C5824 CS_BIAS.n467 GND 0.011784f
C5825 CS_BIAS.n468 GND 0.004799f
C5826 CS_BIAS.n469 GND 0.005932f
C5827 CS_BIAS.n470 GND 0.005932f
C5828 CS_BIAS.n471 GND 0.005932f
C5829 CS_BIAS.n472 GND 0.007471f
C5830 CS_BIAS.n473 GND 0.083017f
C5831 CS_BIAS.n474 GND 0.0091f
C5832 CS_BIAS.n475 GND 0.010086f
C5833 CS_BIAS.n476 GND 0.005932f
C5834 CS_BIAS.n477 GND 0.005932f
C5835 CS_BIAS.n478 GND 0.005932f
C5836 CS_BIAS.n479 GND 0.011104f
C5837 CS_BIAS.n480 GND 0.005625f
C5838 CS_BIAS.n481 GND 0.083017f
C5839 CS_BIAS.n482 GND 0.010947f
C5840 CS_BIAS.n483 GND 0.005932f
C5841 CS_BIAS.n484 GND 0.005932f
C5842 CS_BIAS.n485 GND 0.005932f
C5843 CS_BIAS.n486 GND 0.009937f
C5844 CS_BIAS.n487 GND 0.009209f
C5845 CS_BIAS.n488 GND 0.083017f
C5846 CS_BIAS.n489 GND 0.007362f
C5847 CS_BIAS.n490 GND 0.005932f
C5848 CS_BIAS.n491 GND 0.005932f
C5849 CS_BIAS.n492 GND 0.005932f
C5850 CS_BIAS.n493 GND 0.004791f
C5851 CS_BIAS.n494 GND 0.011729f
C5852 CS_BIAS.t41 GND 0.221674f
C5853 CS_BIAS.n495 GND 0.083017f
C5854 CS_BIAS.n496 GND 0.007362f
C5855 CS_BIAS.n497 GND 0.005932f
C5856 CS_BIAS.n498 GND 0.005932f
C5857 CS_BIAS.n499 GND 0.005932f
C5858 CS_BIAS.n500 GND 0.009937f
C5859 CS_BIAS.n501 GND 0.007311f
C5860 CS_BIAS.n502 GND 0.010947f
C5861 CS_BIAS.n503 GND 0.005932f
C5862 CS_BIAS.n504 GND 0.005932f
C5863 CS_BIAS.n505 GND 0.005625f
C5864 CS_BIAS.n506 GND 0.011104f
C5865 CS_BIAS.n507 GND 0.007058f
C5866 CS_BIAS.n508 GND 0.005932f
C5867 CS_BIAS.n509 GND 0.005932f
C5868 CS_BIAS.n510 GND 0.005932f
C5869 CS_BIAS.n511 GND 0.0091f
C5870 CS_BIAS.n512 GND 0.083017f
C5871 CS_BIAS.n513 GND 0.007471f
C5872 CS_BIAS.n514 GND 0.011666f
C5873 CS_BIAS.n515 GND 0.005932f
C5874 CS_BIAS.n516 GND 0.005932f
C5875 CS_BIAS.n517 GND 0.005932f
C5876 CS_BIAS.n518 GND 0.011784f
C5877 CS_BIAS.n519 GND 0.007254f
C5878 CS_BIAS.n520 GND 0.083017f
C5879 CS_BIAS.n521 GND 0.009318f
C5880 CS_BIAS.n522 GND 0.005932f
C5881 CS_BIAS.n523 GND 0.005932f
C5882 CS_BIAS.n524 GND 0.005932f
C5883 CS_BIAS.n525 GND 0.007475f
C5884 CS_BIAS.n526 GND 0.010838f
C5885 CS_BIAS.n527 GND 0.102559f
C5886 CS_BIAS.n528 GND 0.021424f
C5887 CS_BIAS.n529 GND 0.162707f
C5888 CS_BIAS.n530 GND 3.03503f
.ends

