* NGSPICE file created from diff_pair_sample_0390.ext - technology: sky130A

.subckt diff_pair_sample_0390 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t1 VP.t0 VTAIL.t2 w_n2502_n2372# sky130_fd_pr__pfet_01v8 ad=2.7378 pd=14.82 as=2.7378 ps=14.82 w=7.02 l=3.5
X1 B.t11 B.t9 B.t10 w_n2502_n2372# sky130_fd_pr__pfet_01v8 ad=2.7378 pd=14.82 as=0 ps=0 w=7.02 l=3.5
X2 VDD1.t0 VP.t1 VTAIL.t3 w_n2502_n2372# sky130_fd_pr__pfet_01v8 ad=2.7378 pd=14.82 as=2.7378 ps=14.82 w=7.02 l=3.5
X3 B.t8 B.t6 B.t7 w_n2502_n2372# sky130_fd_pr__pfet_01v8 ad=2.7378 pd=14.82 as=0 ps=0 w=7.02 l=3.5
X4 B.t5 B.t3 B.t4 w_n2502_n2372# sky130_fd_pr__pfet_01v8 ad=2.7378 pd=14.82 as=0 ps=0 w=7.02 l=3.5
X5 VDD2.t1 VN.t0 VTAIL.t1 w_n2502_n2372# sky130_fd_pr__pfet_01v8 ad=2.7378 pd=14.82 as=2.7378 ps=14.82 w=7.02 l=3.5
X6 B.t2 B.t0 B.t1 w_n2502_n2372# sky130_fd_pr__pfet_01v8 ad=2.7378 pd=14.82 as=0 ps=0 w=7.02 l=3.5
X7 VDD2.t0 VN.t1 VTAIL.t0 w_n2502_n2372# sky130_fd_pr__pfet_01v8 ad=2.7378 pd=14.82 as=2.7378 ps=14.82 w=7.02 l=3.5
R0 VP.n0 VP.t1 130.454
R1 VP.n0 VP.t0 87.1839
R2 VP VP.n0 0.526373
R3 VTAIL.n1 VTAIL.t1 73.554
R4 VTAIL.n2 VTAIL.t3 73.5538
R5 VTAIL.n3 VTAIL.t0 73.5538
R6 VTAIL.n0 VTAIL.t2 73.5538
R7 VTAIL.n1 VTAIL.n0 25.0221
R8 VTAIL.n3 VTAIL.n2 21.7203
R9 VTAIL.n2 VTAIL.n1 2.12119
R10 VTAIL VTAIL.n0 1.35395
R11 VTAIL VTAIL.n3 0.767741
R12 VDD1 VDD1.t1 127.897
R13 VDD1 VDD1.t0 91.1162
R14 B.n276 B.n85 585
R15 B.n275 B.n274 585
R16 B.n273 B.n86 585
R17 B.n272 B.n271 585
R18 B.n270 B.n87 585
R19 B.n269 B.n268 585
R20 B.n267 B.n88 585
R21 B.n266 B.n265 585
R22 B.n264 B.n89 585
R23 B.n263 B.n262 585
R24 B.n261 B.n90 585
R25 B.n260 B.n259 585
R26 B.n258 B.n91 585
R27 B.n257 B.n256 585
R28 B.n255 B.n92 585
R29 B.n254 B.n253 585
R30 B.n252 B.n93 585
R31 B.n251 B.n250 585
R32 B.n249 B.n94 585
R33 B.n248 B.n247 585
R34 B.n246 B.n95 585
R35 B.n245 B.n244 585
R36 B.n243 B.n96 585
R37 B.n242 B.n241 585
R38 B.n240 B.n97 585
R39 B.n239 B.n238 585
R40 B.n237 B.n98 585
R41 B.n235 B.n234 585
R42 B.n233 B.n101 585
R43 B.n232 B.n231 585
R44 B.n230 B.n102 585
R45 B.n229 B.n228 585
R46 B.n227 B.n103 585
R47 B.n226 B.n225 585
R48 B.n224 B.n104 585
R49 B.n223 B.n222 585
R50 B.n221 B.n105 585
R51 B.n220 B.n219 585
R52 B.n215 B.n106 585
R53 B.n214 B.n213 585
R54 B.n212 B.n107 585
R55 B.n211 B.n210 585
R56 B.n209 B.n108 585
R57 B.n208 B.n207 585
R58 B.n206 B.n109 585
R59 B.n205 B.n204 585
R60 B.n203 B.n110 585
R61 B.n202 B.n201 585
R62 B.n200 B.n111 585
R63 B.n199 B.n198 585
R64 B.n197 B.n112 585
R65 B.n196 B.n195 585
R66 B.n194 B.n113 585
R67 B.n193 B.n192 585
R68 B.n191 B.n114 585
R69 B.n190 B.n189 585
R70 B.n188 B.n115 585
R71 B.n187 B.n186 585
R72 B.n185 B.n116 585
R73 B.n184 B.n183 585
R74 B.n182 B.n117 585
R75 B.n181 B.n180 585
R76 B.n179 B.n118 585
R77 B.n178 B.n177 585
R78 B.n278 B.n277 585
R79 B.n279 B.n84 585
R80 B.n281 B.n280 585
R81 B.n282 B.n83 585
R82 B.n284 B.n283 585
R83 B.n285 B.n82 585
R84 B.n287 B.n286 585
R85 B.n288 B.n81 585
R86 B.n290 B.n289 585
R87 B.n291 B.n80 585
R88 B.n293 B.n292 585
R89 B.n294 B.n79 585
R90 B.n296 B.n295 585
R91 B.n297 B.n78 585
R92 B.n299 B.n298 585
R93 B.n300 B.n77 585
R94 B.n302 B.n301 585
R95 B.n303 B.n76 585
R96 B.n305 B.n304 585
R97 B.n306 B.n75 585
R98 B.n308 B.n307 585
R99 B.n309 B.n74 585
R100 B.n311 B.n310 585
R101 B.n312 B.n73 585
R102 B.n314 B.n313 585
R103 B.n315 B.n72 585
R104 B.n317 B.n316 585
R105 B.n318 B.n71 585
R106 B.n320 B.n319 585
R107 B.n321 B.n70 585
R108 B.n323 B.n322 585
R109 B.n324 B.n69 585
R110 B.n326 B.n325 585
R111 B.n327 B.n68 585
R112 B.n329 B.n328 585
R113 B.n330 B.n67 585
R114 B.n332 B.n331 585
R115 B.n333 B.n66 585
R116 B.n335 B.n334 585
R117 B.n336 B.n65 585
R118 B.n338 B.n337 585
R119 B.n339 B.n64 585
R120 B.n341 B.n340 585
R121 B.n342 B.n63 585
R122 B.n344 B.n343 585
R123 B.n345 B.n62 585
R124 B.n347 B.n346 585
R125 B.n348 B.n61 585
R126 B.n350 B.n349 585
R127 B.n351 B.n60 585
R128 B.n353 B.n352 585
R129 B.n354 B.n59 585
R130 B.n356 B.n355 585
R131 B.n357 B.n58 585
R132 B.n359 B.n358 585
R133 B.n360 B.n57 585
R134 B.n362 B.n361 585
R135 B.n363 B.n56 585
R136 B.n365 B.n364 585
R137 B.n366 B.n55 585
R138 B.n368 B.n367 585
R139 B.n369 B.n54 585
R140 B.n466 B.n17 585
R141 B.n465 B.n464 585
R142 B.n463 B.n18 585
R143 B.n462 B.n461 585
R144 B.n460 B.n19 585
R145 B.n459 B.n458 585
R146 B.n457 B.n20 585
R147 B.n456 B.n455 585
R148 B.n454 B.n21 585
R149 B.n453 B.n452 585
R150 B.n451 B.n22 585
R151 B.n450 B.n449 585
R152 B.n448 B.n23 585
R153 B.n447 B.n446 585
R154 B.n445 B.n24 585
R155 B.n444 B.n443 585
R156 B.n442 B.n25 585
R157 B.n441 B.n440 585
R158 B.n439 B.n26 585
R159 B.n438 B.n437 585
R160 B.n436 B.n27 585
R161 B.n435 B.n434 585
R162 B.n433 B.n28 585
R163 B.n432 B.n431 585
R164 B.n430 B.n29 585
R165 B.n429 B.n428 585
R166 B.n427 B.n30 585
R167 B.n426 B.n425 585
R168 B.n424 B.n31 585
R169 B.n423 B.n422 585
R170 B.n421 B.n35 585
R171 B.n420 B.n419 585
R172 B.n418 B.n36 585
R173 B.n417 B.n416 585
R174 B.n415 B.n37 585
R175 B.n414 B.n413 585
R176 B.n412 B.n38 585
R177 B.n410 B.n409 585
R178 B.n408 B.n41 585
R179 B.n407 B.n406 585
R180 B.n405 B.n42 585
R181 B.n404 B.n403 585
R182 B.n402 B.n43 585
R183 B.n401 B.n400 585
R184 B.n399 B.n44 585
R185 B.n398 B.n397 585
R186 B.n396 B.n45 585
R187 B.n395 B.n394 585
R188 B.n393 B.n46 585
R189 B.n392 B.n391 585
R190 B.n390 B.n47 585
R191 B.n389 B.n388 585
R192 B.n387 B.n48 585
R193 B.n386 B.n385 585
R194 B.n384 B.n49 585
R195 B.n383 B.n382 585
R196 B.n381 B.n50 585
R197 B.n380 B.n379 585
R198 B.n378 B.n51 585
R199 B.n377 B.n376 585
R200 B.n375 B.n52 585
R201 B.n374 B.n373 585
R202 B.n372 B.n53 585
R203 B.n371 B.n370 585
R204 B.n468 B.n467 585
R205 B.n469 B.n16 585
R206 B.n471 B.n470 585
R207 B.n472 B.n15 585
R208 B.n474 B.n473 585
R209 B.n475 B.n14 585
R210 B.n477 B.n476 585
R211 B.n478 B.n13 585
R212 B.n480 B.n479 585
R213 B.n481 B.n12 585
R214 B.n483 B.n482 585
R215 B.n484 B.n11 585
R216 B.n486 B.n485 585
R217 B.n487 B.n10 585
R218 B.n489 B.n488 585
R219 B.n490 B.n9 585
R220 B.n492 B.n491 585
R221 B.n493 B.n8 585
R222 B.n495 B.n494 585
R223 B.n496 B.n7 585
R224 B.n498 B.n497 585
R225 B.n499 B.n6 585
R226 B.n501 B.n500 585
R227 B.n502 B.n5 585
R228 B.n504 B.n503 585
R229 B.n505 B.n4 585
R230 B.n507 B.n506 585
R231 B.n508 B.n3 585
R232 B.n510 B.n509 585
R233 B.n511 B.n0 585
R234 B.n2 B.n1 585
R235 B.n134 B.n133 585
R236 B.n136 B.n135 585
R237 B.n137 B.n132 585
R238 B.n139 B.n138 585
R239 B.n140 B.n131 585
R240 B.n142 B.n141 585
R241 B.n143 B.n130 585
R242 B.n145 B.n144 585
R243 B.n146 B.n129 585
R244 B.n148 B.n147 585
R245 B.n149 B.n128 585
R246 B.n151 B.n150 585
R247 B.n152 B.n127 585
R248 B.n154 B.n153 585
R249 B.n155 B.n126 585
R250 B.n157 B.n156 585
R251 B.n158 B.n125 585
R252 B.n160 B.n159 585
R253 B.n161 B.n124 585
R254 B.n163 B.n162 585
R255 B.n164 B.n123 585
R256 B.n166 B.n165 585
R257 B.n167 B.n122 585
R258 B.n169 B.n168 585
R259 B.n170 B.n121 585
R260 B.n172 B.n171 585
R261 B.n173 B.n120 585
R262 B.n175 B.n174 585
R263 B.n176 B.n119 585
R264 B.n177 B.n176 482.89
R265 B.n277 B.n276 482.89
R266 B.n371 B.n54 482.89
R267 B.n468 B.n17 482.89
R268 B.n216 B.t3 257.432
R269 B.n99 B.t9 257.432
R270 B.n39 B.t6 257.432
R271 B.n32 B.t0 257.432
R272 B.n513 B.n512 256.663
R273 B.n512 B.n511 235.042
R274 B.n512 B.n2 235.042
R275 B.n99 B.t10 188.149
R276 B.n39 B.t8 188.149
R277 B.n216 B.t4 188.143
R278 B.n32 B.t2 188.143
R279 B.n177 B.n118 163.367
R280 B.n181 B.n118 163.367
R281 B.n182 B.n181 163.367
R282 B.n183 B.n182 163.367
R283 B.n183 B.n116 163.367
R284 B.n187 B.n116 163.367
R285 B.n188 B.n187 163.367
R286 B.n189 B.n188 163.367
R287 B.n189 B.n114 163.367
R288 B.n193 B.n114 163.367
R289 B.n194 B.n193 163.367
R290 B.n195 B.n194 163.367
R291 B.n195 B.n112 163.367
R292 B.n199 B.n112 163.367
R293 B.n200 B.n199 163.367
R294 B.n201 B.n200 163.367
R295 B.n201 B.n110 163.367
R296 B.n205 B.n110 163.367
R297 B.n206 B.n205 163.367
R298 B.n207 B.n206 163.367
R299 B.n207 B.n108 163.367
R300 B.n211 B.n108 163.367
R301 B.n212 B.n211 163.367
R302 B.n213 B.n212 163.367
R303 B.n213 B.n106 163.367
R304 B.n220 B.n106 163.367
R305 B.n221 B.n220 163.367
R306 B.n222 B.n221 163.367
R307 B.n222 B.n104 163.367
R308 B.n226 B.n104 163.367
R309 B.n227 B.n226 163.367
R310 B.n228 B.n227 163.367
R311 B.n228 B.n102 163.367
R312 B.n232 B.n102 163.367
R313 B.n233 B.n232 163.367
R314 B.n234 B.n233 163.367
R315 B.n234 B.n98 163.367
R316 B.n239 B.n98 163.367
R317 B.n240 B.n239 163.367
R318 B.n241 B.n240 163.367
R319 B.n241 B.n96 163.367
R320 B.n245 B.n96 163.367
R321 B.n246 B.n245 163.367
R322 B.n247 B.n246 163.367
R323 B.n247 B.n94 163.367
R324 B.n251 B.n94 163.367
R325 B.n252 B.n251 163.367
R326 B.n253 B.n252 163.367
R327 B.n253 B.n92 163.367
R328 B.n257 B.n92 163.367
R329 B.n258 B.n257 163.367
R330 B.n259 B.n258 163.367
R331 B.n259 B.n90 163.367
R332 B.n263 B.n90 163.367
R333 B.n264 B.n263 163.367
R334 B.n265 B.n264 163.367
R335 B.n265 B.n88 163.367
R336 B.n269 B.n88 163.367
R337 B.n270 B.n269 163.367
R338 B.n271 B.n270 163.367
R339 B.n271 B.n86 163.367
R340 B.n275 B.n86 163.367
R341 B.n276 B.n275 163.367
R342 B.n367 B.n54 163.367
R343 B.n367 B.n366 163.367
R344 B.n366 B.n365 163.367
R345 B.n365 B.n56 163.367
R346 B.n361 B.n56 163.367
R347 B.n361 B.n360 163.367
R348 B.n360 B.n359 163.367
R349 B.n359 B.n58 163.367
R350 B.n355 B.n58 163.367
R351 B.n355 B.n354 163.367
R352 B.n354 B.n353 163.367
R353 B.n353 B.n60 163.367
R354 B.n349 B.n60 163.367
R355 B.n349 B.n348 163.367
R356 B.n348 B.n347 163.367
R357 B.n347 B.n62 163.367
R358 B.n343 B.n62 163.367
R359 B.n343 B.n342 163.367
R360 B.n342 B.n341 163.367
R361 B.n341 B.n64 163.367
R362 B.n337 B.n64 163.367
R363 B.n337 B.n336 163.367
R364 B.n336 B.n335 163.367
R365 B.n335 B.n66 163.367
R366 B.n331 B.n66 163.367
R367 B.n331 B.n330 163.367
R368 B.n330 B.n329 163.367
R369 B.n329 B.n68 163.367
R370 B.n325 B.n68 163.367
R371 B.n325 B.n324 163.367
R372 B.n324 B.n323 163.367
R373 B.n323 B.n70 163.367
R374 B.n319 B.n70 163.367
R375 B.n319 B.n318 163.367
R376 B.n318 B.n317 163.367
R377 B.n317 B.n72 163.367
R378 B.n313 B.n72 163.367
R379 B.n313 B.n312 163.367
R380 B.n312 B.n311 163.367
R381 B.n311 B.n74 163.367
R382 B.n307 B.n74 163.367
R383 B.n307 B.n306 163.367
R384 B.n306 B.n305 163.367
R385 B.n305 B.n76 163.367
R386 B.n301 B.n76 163.367
R387 B.n301 B.n300 163.367
R388 B.n300 B.n299 163.367
R389 B.n299 B.n78 163.367
R390 B.n295 B.n78 163.367
R391 B.n295 B.n294 163.367
R392 B.n294 B.n293 163.367
R393 B.n293 B.n80 163.367
R394 B.n289 B.n80 163.367
R395 B.n289 B.n288 163.367
R396 B.n288 B.n287 163.367
R397 B.n287 B.n82 163.367
R398 B.n283 B.n82 163.367
R399 B.n283 B.n282 163.367
R400 B.n282 B.n281 163.367
R401 B.n281 B.n84 163.367
R402 B.n277 B.n84 163.367
R403 B.n464 B.n17 163.367
R404 B.n464 B.n463 163.367
R405 B.n463 B.n462 163.367
R406 B.n462 B.n19 163.367
R407 B.n458 B.n19 163.367
R408 B.n458 B.n457 163.367
R409 B.n457 B.n456 163.367
R410 B.n456 B.n21 163.367
R411 B.n452 B.n21 163.367
R412 B.n452 B.n451 163.367
R413 B.n451 B.n450 163.367
R414 B.n450 B.n23 163.367
R415 B.n446 B.n23 163.367
R416 B.n446 B.n445 163.367
R417 B.n445 B.n444 163.367
R418 B.n444 B.n25 163.367
R419 B.n440 B.n25 163.367
R420 B.n440 B.n439 163.367
R421 B.n439 B.n438 163.367
R422 B.n438 B.n27 163.367
R423 B.n434 B.n27 163.367
R424 B.n434 B.n433 163.367
R425 B.n433 B.n432 163.367
R426 B.n432 B.n29 163.367
R427 B.n428 B.n29 163.367
R428 B.n428 B.n427 163.367
R429 B.n427 B.n426 163.367
R430 B.n426 B.n31 163.367
R431 B.n422 B.n31 163.367
R432 B.n422 B.n421 163.367
R433 B.n421 B.n420 163.367
R434 B.n420 B.n36 163.367
R435 B.n416 B.n36 163.367
R436 B.n416 B.n415 163.367
R437 B.n415 B.n414 163.367
R438 B.n414 B.n38 163.367
R439 B.n409 B.n38 163.367
R440 B.n409 B.n408 163.367
R441 B.n408 B.n407 163.367
R442 B.n407 B.n42 163.367
R443 B.n403 B.n42 163.367
R444 B.n403 B.n402 163.367
R445 B.n402 B.n401 163.367
R446 B.n401 B.n44 163.367
R447 B.n397 B.n44 163.367
R448 B.n397 B.n396 163.367
R449 B.n396 B.n395 163.367
R450 B.n395 B.n46 163.367
R451 B.n391 B.n46 163.367
R452 B.n391 B.n390 163.367
R453 B.n390 B.n389 163.367
R454 B.n389 B.n48 163.367
R455 B.n385 B.n48 163.367
R456 B.n385 B.n384 163.367
R457 B.n384 B.n383 163.367
R458 B.n383 B.n50 163.367
R459 B.n379 B.n50 163.367
R460 B.n379 B.n378 163.367
R461 B.n378 B.n377 163.367
R462 B.n377 B.n52 163.367
R463 B.n373 B.n52 163.367
R464 B.n373 B.n372 163.367
R465 B.n372 B.n371 163.367
R466 B.n469 B.n468 163.367
R467 B.n470 B.n469 163.367
R468 B.n470 B.n15 163.367
R469 B.n474 B.n15 163.367
R470 B.n475 B.n474 163.367
R471 B.n476 B.n475 163.367
R472 B.n476 B.n13 163.367
R473 B.n480 B.n13 163.367
R474 B.n481 B.n480 163.367
R475 B.n482 B.n481 163.367
R476 B.n482 B.n11 163.367
R477 B.n486 B.n11 163.367
R478 B.n487 B.n486 163.367
R479 B.n488 B.n487 163.367
R480 B.n488 B.n9 163.367
R481 B.n492 B.n9 163.367
R482 B.n493 B.n492 163.367
R483 B.n494 B.n493 163.367
R484 B.n494 B.n7 163.367
R485 B.n498 B.n7 163.367
R486 B.n499 B.n498 163.367
R487 B.n500 B.n499 163.367
R488 B.n500 B.n5 163.367
R489 B.n504 B.n5 163.367
R490 B.n505 B.n504 163.367
R491 B.n506 B.n505 163.367
R492 B.n506 B.n3 163.367
R493 B.n510 B.n3 163.367
R494 B.n511 B.n510 163.367
R495 B.n134 B.n2 163.367
R496 B.n135 B.n134 163.367
R497 B.n135 B.n132 163.367
R498 B.n139 B.n132 163.367
R499 B.n140 B.n139 163.367
R500 B.n141 B.n140 163.367
R501 B.n141 B.n130 163.367
R502 B.n145 B.n130 163.367
R503 B.n146 B.n145 163.367
R504 B.n147 B.n146 163.367
R505 B.n147 B.n128 163.367
R506 B.n151 B.n128 163.367
R507 B.n152 B.n151 163.367
R508 B.n153 B.n152 163.367
R509 B.n153 B.n126 163.367
R510 B.n157 B.n126 163.367
R511 B.n158 B.n157 163.367
R512 B.n159 B.n158 163.367
R513 B.n159 B.n124 163.367
R514 B.n163 B.n124 163.367
R515 B.n164 B.n163 163.367
R516 B.n165 B.n164 163.367
R517 B.n165 B.n122 163.367
R518 B.n169 B.n122 163.367
R519 B.n170 B.n169 163.367
R520 B.n171 B.n170 163.367
R521 B.n171 B.n120 163.367
R522 B.n175 B.n120 163.367
R523 B.n176 B.n175 163.367
R524 B.n100 B.t11 113.871
R525 B.n40 B.t7 113.871
R526 B.n217 B.t5 113.864
R527 B.n33 B.t1 113.864
R528 B.n217 B.n216 74.2793
R529 B.n100 B.n99 74.2793
R530 B.n40 B.n39 74.2793
R531 B.n33 B.n32 74.2793
R532 B.n218 B.n217 59.5399
R533 B.n236 B.n100 59.5399
R534 B.n411 B.n40 59.5399
R535 B.n34 B.n33 59.5399
R536 B.n467 B.n466 31.3761
R537 B.n370 B.n369 31.3761
R538 B.n278 B.n85 31.3761
R539 B.n178 B.n119 31.3761
R540 B B.n513 18.0485
R541 B.n467 B.n16 10.6151
R542 B.n471 B.n16 10.6151
R543 B.n472 B.n471 10.6151
R544 B.n473 B.n472 10.6151
R545 B.n473 B.n14 10.6151
R546 B.n477 B.n14 10.6151
R547 B.n478 B.n477 10.6151
R548 B.n479 B.n478 10.6151
R549 B.n479 B.n12 10.6151
R550 B.n483 B.n12 10.6151
R551 B.n484 B.n483 10.6151
R552 B.n485 B.n484 10.6151
R553 B.n485 B.n10 10.6151
R554 B.n489 B.n10 10.6151
R555 B.n490 B.n489 10.6151
R556 B.n491 B.n490 10.6151
R557 B.n491 B.n8 10.6151
R558 B.n495 B.n8 10.6151
R559 B.n496 B.n495 10.6151
R560 B.n497 B.n496 10.6151
R561 B.n497 B.n6 10.6151
R562 B.n501 B.n6 10.6151
R563 B.n502 B.n501 10.6151
R564 B.n503 B.n502 10.6151
R565 B.n503 B.n4 10.6151
R566 B.n507 B.n4 10.6151
R567 B.n508 B.n507 10.6151
R568 B.n509 B.n508 10.6151
R569 B.n509 B.n0 10.6151
R570 B.n466 B.n465 10.6151
R571 B.n465 B.n18 10.6151
R572 B.n461 B.n18 10.6151
R573 B.n461 B.n460 10.6151
R574 B.n460 B.n459 10.6151
R575 B.n459 B.n20 10.6151
R576 B.n455 B.n20 10.6151
R577 B.n455 B.n454 10.6151
R578 B.n454 B.n453 10.6151
R579 B.n453 B.n22 10.6151
R580 B.n449 B.n22 10.6151
R581 B.n449 B.n448 10.6151
R582 B.n448 B.n447 10.6151
R583 B.n447 B.n24 10.6151
R584 B.n443 B.n24 10.6151
R585 B.n443 B.n442 10.6151
R586 B.n442 B.n441 10.6151
R587 B.n441 B.n26 10.6151
R588 B.n437 B.n26 10.6151
R589 B.n437 B.n436 10.6151
R590 B.n436 B.n435 10.6151
R591 B.n435 B.n28 10.6151
R592 B.n431 B.n28 10.6151
R593 B.n431 B.n430 10.6151
R594 B.n430 B.n429 10.6151
R595 B.n429 B.n30 10.6151
R596 B.n425 B.n424 10.6151
R597 B.n424 B.n423 10.6151
R598 B.n423 B.n35 10.6151
R599 B.n419 B.n35 10.6151
R600 B.n419 B.n418 10.6151
R601 B.n418 B.n417 10.6151
R602 B.n417 B.n37 10.6151
R603 B.n413 B.n37 10.6151
R604 B.n413 B.n412 10.6151
R605 B.n410 B.n41 10.6151
R606 B.n406 B.n41 10.6151
R607 B.n406 B.n405 10.6151
R608 B.n405 B.n404 10.6151
R609 B.n404 B.n43 10.6151
R610 B.n400 B.n43 10.6151
R611 B.n400 B.n399 10.6151
R612 B.n399 B.n398 10.6151
R613 B.n398 B.n45 10.6151
R614 B.n394 B.n45 10.6151
R615 B.n394 B.n393 10.6151
R616 B.n393 B.n392 10.6151
R617 B.n392 B.n47 10.6151
R618 B.n388 B.n47 10.6151
R619 B.n388 B.n387 10.6151
R620 B.n387 B.n386 10.6151
R621 B.n386 B.n49 10.6151
R622 B.n382 B.n49 10.6151
R623 B.n382 B.n381 10.6151
R624 B.n381 B.n380 10.6151
R625 B.n380 B.n51 10.6151
R626 B.n376 B.n51 10.6151
R627 B.n376 B.n375 10.6151
R628 B.n375 B.n374 10.6151
R629 B.n374 B.n53 10.6151
R630 B.n370 B.n53 10.6151
R631 B.n369 B.n368 10.6151
R632 B.n368 B.n55 10.6151
R633 B.n364 B.n55 10.6151
R634 B.n364 B.n363 10.6151
R635 B.n363 B.n362 10.6151
R636 B.n362 B.n57 10.6151
R637 B.n358 B.n57 10.6151
R638 B.n358 B.n357 10.6151
R639 B.n357 B.n356 10.6151
R640 B.n356 B.n59 10.6151
R641 B.n352 B.n59 10.6151
R642 B.n352 B.n351 10.6151
R643 B.n351 B.n350 10.6151
R644 B.n350 B.n61 10.6151
R645 B.n346 B.n61 10.6151
R646 B.n346 B.n345 10.6151
R647 B.n345 B.n344 10.6151
R648 B.n344 B.n63 10.6151
R649 B.n340 B.n63 10.6151
R650 B.n340 B.n339 10.6151
R651 B.n339 B.n338 10.6151
R652 B.n338 B.n65 10.6151
R653 B.n334 B.n65 10.6151
R654 B.n334 B.n333 10.6151
R655 B.n333 B.n332 10.6151
R656 B.n332 B.n67 10.6151
R657 B.n328 B.n67 10.6151
R658 B.n328 B.n327 10.6151
R659 B.n327 B.n326 10.6151
R660 B.n326 B.n69 10.6151
R661 B.n322 B.n69 10.6151
R662 B.n322 B.n321 10.6151
R663 B.n321 B.n320 10.6151
R664 B.n320 B.n71 10.6151
R665 B.n316 B.n71 10.6151
R666 B.n316 B.n315 10.6151
R667 B.n315 B.n314 10.6151
R668 B.n314 B.n73 10.6151
R669 B.n310 B.n73 10.6151
R670 B.n310 B.n309 10.6151
R671 B.n309 B.n308 10.6151
R672 B.n308 B.n75 10.6151
R673 B.n304 B.n75 10.6151
R674 B.n304 B.n303 10.6151
R675 B.n303 B.n302 10.6151
R676 B.n302 B.n77 10.6151
R677 B.n298 B.n77 10.6151
R678 B.n298 B.n297 10.6151
R679 B.n297 B.n296 10.6151
R680 B.n296 B.n79 10.6151
R681 B.n292 B.n79 10.6151
R682 B.n292 B.n291 10.6151
R683 B.n291 B.n290 10.6151
R684 B.n290 B.n81 10.6151
R685 B.n286 B.n81 10.6151
R686 B.n286 B.n285 10.6151
R687 B.n285 B.n284 10.6151
R688 B.n284 B.n83 10.6151
R689 B.n280 B.n83 10.6151
R690 B.n280 B.n279 10.6151
R691 B.n279 B.n278 10.6151
R692 B.n133 B.n1 10.6151
R693 B.n136 B.n133 10.6151
R694 B.n137 B.n136 10.6151
R695 B.n138 B.n137 10.6151
R696 B.n138 B.n131 10.6151
R697 B.n142 B.n131 10.6151
R698 B.n143 B.n142 10.6151
R699 B.n144 B.n143 10.6151
R700 B.n144 B.n129 10.6151
R701 B.n148 B.n129 10.6151
R702 B.n149 B.n148 10.6151
R703 B.n150 B.n149 10.6151
R704 B.n150 B.n127 10.6151
R705 B.n154 B.n127 10.6151
R706 B.n155 B.n154 10.6151
R707 B.n156 B.n155 10.6151
R708 B.n156 B.n125 10.6151
R709 B.n160 B.n125 10.6151
R710 B.n161 B.n160 10.6151
R711 B.n162 B.n161 10.6151
R712 B.n162 B.n123 10.6151
R713 B.n166 B.n123 10.6151
R714 B.n167 B.n166 10.6151
R715 B.n168 B.n167 10.6151
R716 B.n168 B.n121 10.6151
R717 B.n172 B.n121 10.6151
R718 B.n173 B.n172 10.6151
R719 B.n174 B.n173 10.6151
R720 B.n174 B.n119 10.6151
R721 B.n179 B.n178 10.6151
R722 B.n180 B.n179 10.6151
R723 B.n180 B.n117 10.6151
R724 B.n184 B.n117 10.6151
R725 B.n185 B.n184 10.6151
R726 B.n186 B.n185 10.6151
R727 B.n186 B.n115 10.6151
R728 B.n190 B.n115 10.6151
R729 B.n191 B.n190 10.6151
R730 B.n192 B.n191 10.6151
R731 B.n192 B.n113 10.6151
R732 B.n196 B.n113 10.6151
R733 B.n197 B.n196 10.6151
R734 B.n198 B.n197 10.6151
R735 B.n198 B.n111 10.6151
R736 B.n202 B.n111 10.6151
R737 B.n203 B.n202 10.6151
R738 B.n204 B.n203 10.6151
R739 B.n204 B.n109 10.6151
R740 B.n208 B.n109 10.6151
R741 B.n209 B.n208 10.6151
R742 B.n210 B.n209 10.6151
R743 B.n210 B.n107 10.6151
R744 B.n214 B.n107 10.6151
R745 B.n215 B.n214 10.6151
R746 B.n219 B.n215 10.6151
R747 B.n223 B.n105 10.6151
R748 B.n224 B.n223 10.6151
R749 B.n225 B.n224 10.6151
R750 B.n225 B.n103 10.6151
R751 B.n229 B.n103 10.6151
R752 B.n230 B.n229 10.6151
R753 B.n231 B.n230 10.6151
R754 B.n231 B.n101 10.6151
R755 B.n235 B.n101 10.6151
R756 B.n238 B.n237 10.6151
R757 B.n238 B.n97 10.6151
R758 B.n242 B.n97 10.6151
R759 B.n243 B.n242 10.6151
R760 B.n244 B.n243 10.6151
R761 B.n244 B.n95 10.6151
R762 B.n248 B.n95 10.6151
R763 B.n249 B.n248 10.6151
R764 B.n250 B.n249 10.6151
R765 B.n250 B.n93 10.6151
R766 B.n254 B.n93 10.6151
R767 B.n255 B.n254 10.6151
R768 B.n256 B.n255 10.6151
R769 B.n256 B.n91 10.6151
R770 B.n260 B.n91 10.6151
R771 B.n261 B.n260 10.6151
R772 B.n262 B.n261 10.6151
R773 B.n262 B.n89 10.6151
R774 B.n266 B.n89 10.6151
R775 B.n267 B.n266 10.6151
R776 B.n268 B.n267 10.6151
R777 B.n268 B.n87 10.6151
R778 B.n272 B.n87 10.6151
R779 B.n273 B.n272 10.6151
R780 B.n274 B.n273 10.6151
R781 B.n274 B.n85 10.6151
R782 B.n34 B.n30 9.36635
R783 B.n411 B.n410 9.36635
R784 B.n219 B.n218 9.36635
R785 B.n237 B.n236 9.36635
R786 B.n513 B.n0 8.11757
R787 B.n513 B.n1 8.11757
R788 B.n425 B.n34 1.24928
R789 B.n412 B.n411 1.24928
R790 B.n218 B.n105 1.24928
R791 B.n236 B.n235 1.24928
R792 VN VN.t0 130.362
R793 VN VN.t1 87.7098
R794 VDD2.n0 VDD2.t0 126.547
R795 VDD2.n0 VDD2.t1 90.2326
R796 VDD2 VDD2.n0 0.884121
C0 w_n2502_n2372# VP 3.7621f
C1 VN VP 4.95105f
C2 w_n2502_n2372# VTAIL 2.09147f
C3 VTAIL VN 1.8567f
C4 VDD1 VP 2.01819f
C5 VP B 1.67716f
C6 w_n2502_n2372# VDD2 1.57902f
C7 VDD2 VN 1.79765f
C8 VDD1 VTAIL 3.98581f
C9 VTAIL B 2.81384f
C10 VDD2 VDD1 0.784143f
C11 VDD2 B 1.46243f
C12 w_n2502_n2372# VN 3.44145f
C13 VTAIL VP 1.87088f
C14 w_n2502_n2372# VDD1 1.542f
C15 VDD2 VP 0.370906f
C16 VDD1 VN 0.14887f
C17 w_n2502_n2372# B 8.38889f
C18 VN B 1.14639f
C19 VDD2 VTAIL 4.04408f
C20 VDD1 B 1.42433f
C21 VDD2 VSUBS 0.760013f
C22 VDD1 VSUBS 4.293912f
C23 VTAIL VSUBS 0.633609f
C24 VN VSUBS 5.7874f
C25 VP VSUBS 1.658737f
C26 B VSUBS 4.148643f
C27 w_n2502_n2372# VSUBS 73.828995f
C28 VDD2.t0 VSUBS 1.02968f
C29 VDD2.t1 VSUBS 0.734898f
C30 VDD2.n0 VSUBS 2.11712f
C31 VN.t1 VSUBS 2.24125f
C32 VN.t0 VSUBS 2.87824f
C33 B.n0 VSUBS 0.006248f
C34 B.n1 VSUBS 0.006248f
C35 B.n2 VSUBS 0.009241f
C36 B.n3 VSUBS 0.007082f
C37 B.n4 VSUBS 0.007082f
C38 B.n5 VSUBS 0.007082f
C39 B.n6 VSUBS 0.007082f
C40 B.n7 VSUBS 0.007082f
C41 B.n8 VSUBS 0.007082f
C42 B.n9 VSUBS 0.007082f
C43 B.n10 VSUBS 0.007082f
C44 B.n11 VSUBS 0.007082f
C45 B.n12 VSUBS 0.007082f
C46 B.n13 VSUBS 0.007082f
C47 B.n14 VSUBS 0.007082f
C48 B.n15 VSUBS 0.007082f
C49 B.n16 VSUBS 0.007082f
C50 B.n17 VSUBS 0.016832f
C51 B.n18 VSUBS 0.007082f
C52 B.n19 VSUBS 0.007082f
C53 B.n20 VSUBS 0.007082f
C54 B.n21 VSUBS 0.007082f
C55 B.n22 VSUBS 0.007082f
C56 B.n23 VSUBS 0.007082f
C57 B.n24 VSUBS 0.007082f
C58 B.n25 VSUBS 0.007082f
C59 B.n26 VSUBS 0.007082f
C60 B.n27 VSUBS 0.007082f
C61 B.n28 VSUBS 0.007082f
C62 B.n29 VSUBS 0.007082f
C63 B.n30 VSUBS 0.006665f
C64 B.n31 VSUBS 0.007082f
C65 B.t1 VSUBS 0.21403f
C66 B.t2 VSUBS 0.239986f
C67 B.t0 VSUBS 1.18379f
C68 B.n32 VSUBS 0.141795f
C69 B.n33 VSUBS 0.075843f
C70 B.n34 VSUBS 0.016407f
C71 B.n35 VSUBS 0.007082f
C72 B.n36 VSUBS 0.007082f
C73 B.n37 VSUBS 0.007082f
C74 B.n38 VSUBS 0.007082f
C75 B.t7 VSUBS 0.214029f
C76 B.t8 VSUBS 0.239984f
C77 B.t6 VSUBS 1.18379f
C78 B.n39 VSUBS 0.141797f
C79 B.n40 VSUBS 0.075844f
C80 B.n41 VSUBS 0.007082f
C81 B.n42 VSUBS 0.007082f
C82 B.n43 VSUBS 0.007082f
C83 B.n44 VSUBS 0.007082f
C84 B.n45 VSUBS 0.007082f
C85 B.n46 VSUBS 0.007082f
C86 B.n47 VSUBS 0.007082f
C87 B.n48 VSUBS 0.007082f
C88 B.n49 VSUBS 0.007082f
C89 B.n50 VSUBS 0.007082f
C90 B.n51 VSUBS 0.007082f
C91 B.n52 VSUBS 0.007082f
C92 B.n53 VSUBS 0.007082f
C93 B.n54 VSUBS 0.015451f
C94 B.n55 VSUBS 0.007082f
C95 B.n56 VSUBS 0.007082f
C96 B.n57 VSUBS 0.007082f
C97 B.n58 VSUBS 0.007082f
C98 B.n59 VSUBS 0.007082f
C99 B.n60 VSUBS 0.007082f
C100 B.n61 VSUBS 0.007082f
C101 B.n62 VSUBS 0.007082f
C102 B.n63 VSUBS 0.007082f
C103 B.n64 VSUBS 0.007082f
C104 B.n65 VSUBS 0.007082f
C105 B.n66 VSUBS 0.007082f
C106 B.n67 VSUBS 0.007082f
C107 B.n68 VSUBS 0.007082f
C108 B.n69 VSUBS 0.007082f
C109 B.n70 VSUBS 0.007082f
C110 B.n71 VSUBS 0.007082f
C111 B.n72 VSUBS 0.007082f
C112 B.n73 VSUBS 0.007082f
C113 B.n74 VSUBS 0.007082f
C114 B.n75 VSUBS 0.007082f
C115 B.n76 VSUBS 0.007082f
C116 B.n77 VSUBS 0.007082f
C117 B.n78 VSUBS 0.007082f
C118 B.n79 VSUBS 0.007082f
C119 B.n80 VSUBS 0.007082f
C120 B.n81 VSUBS 0.007082f
C121 B.n82 VSUBS 0.007082f
C122 B.n83 VSUBS 0.007082f
C123 B.n84 VSUBS 0.007082f
C124 B.n85 VSUBS 0.015961f
C125 B.n86 VSUBS 0.007082f
C126 B.n87 VSUBS 0.007082f
C127 B.n88 VSUBS 0.007082f
C128 B.n89 VSUBS 0.007082f
C129 B.n90 VSUBS 0.007082f
C130 B.n91 VSUBS 0.007082f
C131 B.n92 VSUBS 0.007082f
C132 B.n93 VSUBS 0.007082f
C133 B.n94 VSUBS 0.007082f
C134 B.n95 VSUBS 0.007082f
C135 B.n96 VSUBS 0.007082f
C136 B.n97 VSUBS 0.007082f
C137 B.n98 VSUBS 0.007082f
C138 B.t11 VSUBS 0.214029f
C139 B.t10 VSUBS 0.239984f
C140 B.t9 VSUBS 1.18379f
C141 B.n99 VSUBS 0.141797f
C142 B.n100 VSUBS 0.075844f
C143 B.n101 VSUBS 0.007082f
C144 B.n102 VSUBS 0.007082f
C145 B.n103 VSUBS 0.007082f
C146 B.n104 VSUBS 0.007082f
C147 B.n105 VSUBS 0.003957f
C148 B.n106 VSUBS 0.007082f
C149 B.n107 VSUBS 0.007082f
C150 B.n108 VSUBS 0.007082f
C151 B.n109 VSUBS 0.007082f
C152 B.n110 VSUBS 0.007082f
C153 B.n111 VSUBS 0.007082f
C154 B.n112 VSUBS 0.007082f
C155 B.n113 VSUBS 0.007082f
C156 B.n114 VSUBS 0.007082f
C157 B.n115 VSUBS 0.007082f
C158 B.n116 VSUBS 0.007082f
C159 B.n117 VSUBS 0.007082f
C160 B.n118 VSUBS 0.007082f
C161 B.n119 VSUBS 0.015451f
C162 B.n120 VSUBS 0.007082f
C163 B.n121 VSUBS 0.007082f
C164 B.n122 VSUBS 0.007082f
C165 B.n123 VSUBS 0.007082f
C166 B.n124 VSUBS 0.007082f
C167 B.n125 VSUBS 0.007082f
C168 B.n126 VSUBS 0.007082f
C169 B.n127 VSUBS 0.007082f
C170 B.n128 VSUBS 0.007082f
C171 B.n129 VSUBS 0.007082f
C172 B.n130 VSUBS 0.007082f
C173 B.n131 VSUBS 0.007082f
C174 B.n132 VSUBS 0.007082f
C175 B.n133 VSUBS 0.007082f
C176 B.n134 VSUBS 0.007082f
C177 B.n135 VSUBS 0.007082f
C178 B.n136 VSUBS 0.007082f
C179 B.n137 VSUBS 0.007082f
C180 B.n138 VSUBS 0.007082f
C181 B.n139 VSUBS 0.007082f
C182 B.n140 VSUBS 0.007082f
C183 B.n141 VSUBS 0.007082f
C184 B.n142 VSUBS 0.007082f
C185 B.n143 VSUBS 0.007082f
C186 B.n144 VSUBS 0.007082f
C187 B.n145 VSUBS 0.007082f
C188 B.n146 VSUBS 0.007082f
C189 B.n147 VSUBS 0.007082f
C190 B.n148 VSUBS 0.007082f
C191 B.n149 VSUBS 0.007082f
C192 B.n150 VSUBS 0.007082f
C193 B.n151 VSUBS 0.007082f
C194 B.n152 VSUBS 0.007082f
C195 B.n153 VSUBS 0.007082f
C196 B.n154 VSUBS 0.007082f
C197 B.n155 VSUBS 0.007082f
C198 B.n156 VSUBS 0.007082f
C199 B.n157 VSUBS 0.007082f
C200 B.n158 VSUBS 0.007082f
C201 B.n159 VSUBS 0.007082f
C202 B.n160 VSUBS 0.007082f
C203 B.n161 VSUBS 0.007082f
C204 B.n162 VSUBS 0.007082f
C205 B.n163 VSUBS 0.007082f
C206 B.n164 VSUBS 0.007082f
C207 B.n165 VSUBS 0.007082f
C208 B.n166 VSUBS 0.007082f
C209 B.n167 VSUBS 0.007082f
C210 B.n168 VSUBS 0.007082f
C211 B.n169 VSUBS 0.007082f
C212 B.n170 VSUBS 0.007082f
C213 B.n171 VSUBS 0.007082f
C214 B.n172 VSUBS 0.007082f
C215 B.n173 VSUBS 0.007082f
C216 B.n174 VSUBS 0.007082f
C217 B.n175 VSUBS 0.007082f
C218 B.n176 VSUBS 0.015451f
C219 B.n177 VSUBS 0.016832f
C220 B.n178 VSUBS 0.016832f
C221 B.n179 VSUBS 0.007082f
C222 B.n180 VSUBS 0.007082f
C223 B.n181 VSUBS 0.007082f
C224 B.n182 VSUBS 0.007082f
C225 B.n183 VSUBS 0.007082f
C226 B.n184 VSUBS 0.007082f
C227 B.n185 VSUBS 0.007082f
C228 B.n186 VSUBS 0.007082f
C229 B.n187 VSUBS 0.007082f
C230 B.n188 VSUBS 0.007082f
C231 B.n189 VSUBS 0.007082f
C232 B.n190 VSUBS 0.007082f
C233 B.n191 VSUBS 0.007082f
C234 B.n192 VSUBS 0.007082f
C235 B.n193 VSUBS 0.007082f
C236 B.n194 VSUBS 0.007082f
C237 B.n195 VSUBS 0.007082f
C238 B.n196 VSUBS 0.007082f
C239 B.n197 VSUBS 0.007082f
C240 B.n198 VSUBS 0.007082f
C241 B.n199 VSUBS 0.007082f
C242 B.n200 VSUBS 0.007082f
C243 B.n201 VSUBS 0.007082f
C244 B.n202 VSUBS 0.007082f
C245 B.n203 VSUBS 0.007082f
C246 B.n204 VSUBS 0.007082f
C247 B.n205 VSUBS 0.007082f
C248 B.n206 VSUBS 0.007082f
C249 B.n207 VSUBS 0.007082f
C250 B.n208 VSUBS 0.007082f
C251 B.n209 VSUBS 0.007082f
C252 B.n210 VSUBS 0.007082f
C253 B.n211 VSUBS 0.007082f
C254 B.n212 VSUBS 0.007082f
C255 B.n213 VSUBS 0.007082f
C256 B.n214 VSUBS 0.007082f
C257 B.n215 VSUBS 0.007082f
C258 B.t5 VSUBS 0.21403f
C259 B.t4 VSUBS 0.239986f
C260 B.t3 VSUBS 1.18379f
C261 B.n216 VSUBS 0.141795f
C262 B.n217 VSUBS 0.075843f
C263 B.n218 VSUBS 0.016407f
C264 B.n219 VSUBS 0.006665f
C265 B.n220 VSUBS 0.007082f
C266 B.n221 VSUBS 0.007082f
C267 B.n222 VSUBS 0.007082f
C268 B.n223 VSUBS 0.007082f
C269 B.n224 VSUBS 0.007082f
C270 B.n225 VSUBS 0.007082f
C271 B.n226 VSUBS 0.007082f
C272 B.n227 VSUBS 0.007082f
C273 B.n228 VSUBS 0.007082f
C274 B.n229 VSUBS 0.007082f
C275 B.n230 VSUBS 0.007082f
C276 B.n231 VSUBS 0.007082f
C277 B.n232 VSUBS 0.007082f
C278 B.n233 VSUBS 0.007082f
C279 B.n234 VSUBS 0.007082f
C280 B.n235 VSUBS 0.003957f
C281 B.n236 VSUBS 0.016407f
C282 B.n237 VSUBS 0.006665f
C283 B.n238 VSUBS 0.007082f
C284 B.n239 VSUBS 0.007082f
C285 B.n240 VSUBS 0.007082f
C286 B.n241 VSUBS 0.007082f
C287 B.n242 VSUBS 0.007082f
C288 B.n243 VSUBS 0.007082f
C289 B.n244 VSUBS 0.007082f
C290 B.n245 VSUBS 0.007082f
C291 B.n246 VSUBS 0.007082f
C292 B.n247 VSUBS 0.007082f
C293 B.n248 VSUBS 0.007082f
C294 B.n249 VSUBS 0.007082f
C295 B.n250 VSUBS 0.007082f
C296 B.n251 VSUBS 0.007082f
C297 B.n252 VSUBS 0.007082f
C298 B.n253 VSUBS 0.007082f
C299 B.n254 VSUBS 0.007082f
C300 B.n255 VSUBS 0.007082f
C301 B.n256 VSUBS 0.007082f
C302 B.n257 VSUBS 0.007082f
C303 B.n258 VSUBS 0.007082f
C304 B.n259 VSUBS 0.007082f
C305 B.n260 VSUBS 0.007082f
C306 B.n261 VSUBS 0.007082f
C307 B.n262 VSUBS 0.007082f
C308 B.n263 VSUBS 0.007082f
C309 B.n264 VSUBS 0.007082f
C310 B.n265 VSUBS 0.007082f
C311 B.n266 VSUBS 0.007082f
C312 B.n267 VSUBS 0.007082f
C313 B.n268 VSUBS 0.007082f
C314 B.n269 VSUBS 0.007082f
C315 B.n270 VSUBS 0.007082f
C316 B.n271 VSUBS 0.007082f
C317 B.n272 VSUBS 0.007082f
C318 B.n273 VSUBS 0.007082f
C319 B.n274 VSUBS 0.007082f
C320 B.n275 VSUBS 0.007082f
C321 B.n276 VSUBS 0.016832f
C322 B.n277 VSUBS 0.015451f
C323 B.n278 VSUBS 0.016322f
C324 B.n279 VSUBS 0.007082f
C325 B.n280 VSUBS 0.007082f
C326 B.n281 VSUBS 0.007082f
C327 B.n282 VSUBS 0.007082f
C328 B.n283 VSUBS 0.007082f
C329 B.n284 VSUBS 0.007082f
C330 B.n285 VSUBS 0.007082f
C331 B.n286 VSUBS 0.007082f
C332 B.n287 VSUBS 0.007082f
C333 B.n288 VSUBS 0.007082f
C334 B.n289 VSUBS 0.007082f
C335 B.n290 VSUBS 0.007082f
C336 B.n291 VSUBS 0.007082f
C337 B.n292 VSUBS 0.007082f
C338 B.n293 VSUBS 0.007082f
C339 B.n294 VSUBS 0.007082f
C340 B.n295 VSUBS 0.007082f
C341 B.n296 VSUBS 0.007082f
C342 B.n297 VSUBS 0.007082f
C343 B.n298 VSUBS 0.007082f
C344 B.n299 VSUBS 0.007082f
C345 B.n300 VSUBS 0.007082f
C346 B.n301 VSUBS 0.007082f
C347 B.n302 VSUBS 0.007082f
C348 B.n303 VSUBS 0.007082f
C349 B.n304 VSUBS 0.007082f
C350 B.n305 VSUBS 0.007082f
C351 B.n306 VSUBS 0.007082f
C352 B.n307 VSUBS 0.007082f
C353 B.n308 VSUBS 0.007082f
C354 B.n309 VSUBS 0.007082f
C355 B.n310 VSUBS 0.007082f
C356 B.n311 VSUBS 0.007082f
C357 B.n312 VSUBS 0.007082f
C358 B.n313 VSUBS 0.007082f
C359 B.n314 VSUBS 0.007082f
C360 B.n315 VSUBS 0.007082f
C361 B.n316 VSUBS 0.007082f
C362 B.n317 VSUBS 0.007082f
C363 B.n318 VSUBS 0.007082f
C364 B.n319 VSUBS 0.007082f
C365 B.n320 VSUBS 0.007082f
C366 B.n321 VSUBS 0.007082f
C367 B.n322 VSUBS 0.007082f
C368 B.n323 VSUBS 0.007082f
C369 B.n324 VSUBS 0.007082f
C370 B.n325 VSUBS 0.007082f
C371 B.n326 VSUBS 0.007082f
C372 B.n327 VSUBS 0.007082f
C373 B.n328 VSUBS 0.007082f
C374 B.n329 VSUBS 0.007082f
C375 B.n330 VSUBS 0.007082f
C376 B.n331 VSUBS 0.007082f
C377 B.n332 VSUBS 0.007082f
C378 B.n333 VSUBS 0.007082f
C379 B.n334 VSUBS 0.007082f
C380 B.n335 VSUBS 0.007082f
C381 B.n336 VSUBS 0.007082f
C382 B.n337 VSUBS 0.007082f
C383 B.n338 VSUBS 0.007082f
C384 B.n339 VSUBS 0.007082f
C385 B.n340 VSUBS 0.007082f
C386 B.n341 VSUBS 0.007082f
C387 B.n342 VSUBS 0.007082f
C388 B.n343 VSUBS 0.007082f
C389 B.n344 VSUBS 0.007082f
C390 B.n345 VSUBS 0.007082f
C391 B.n346 VSUBS 0.007082f
C392 B.n347 VSUBS 0.007082f
C393 B.n348 VSUBS 0.007082f
C394 B.n349 VSUBS 0.007082f
C395 B.n350 VSUBS 0.007082f
C396 B.n351 VSUBS 0.007082f
C397 B.n352 VSUBS 0.007082f
C398 B.n353 VSUBS 0.007082f
C399 B.n354 VSUBS 0.007082f
C400 B.n355 VSUBS 0.007082f
C401 B.n356 VSUBS 0.007082f
C402 B.n357 VSUBS 0.007082f
C403 B.n358 VSUBS 0.007082f
C404 B.n359 VSUBS 0.007082f
C405 B.n360 VSUBS 0.007082f
C406 B.n361 VSUBS 0.007082f
C407 B.n362 VSUBS 0.007082f
C408 B.n363 VSUBS 0.007082f
C409 B.n364 VSUBS 0.007082f
C410 B.n365 VSUBS 0.007082f
C411 B.n366 VSUBS 0.007082f
C412 B.n367 VSUBS 0.007082f
C413 B.n368 VSUBS 0.007082f
C414 B.n369 VSUBS 0.015451f
C415 B.n370 VSUBS 0.016832f
C416 B.n371 VSUBS 0.016832f
C417 B.n372 VSUBS 0.007082f
C418 B.n373 VSUBS 0.007082f
C419 B.n374 VSUBS 0.007082f
C420 B.n375 VSUBS 0.007082f
C421 B.n376 VSUBS 0.007082f
C422 B.n377 VSUBS 0.007082f
C423 B.n378 VSUBS 0.007082f
C424 B.n379 VSUBS 0.007082f
C425 B.n380 VSUBS 0.007082f
C426 B.n381 VSUBS 0.007082f
C427 B.n382 VSUBS 0.007082f
C428 B.n383 VSUBS 0.007082f
C429 B.n384 VSUBS 0.007082f
C430 B.n385 VSUBS 0.007082f
C431 B.n386 VSUBS 0.007082f
C432 B.n387 VSUBS 0.007082f
C433 B.n388 VSUBS 0.007082f
C434 B.n389 VSUBS 0.007082f
C435 B.n390 VSUBS 0.007082f
C436 B.n391 VSUBS 0.007082f
C437 B.n392 VSUBS 0.007082f
C438 B.n393 VSUBS 0.007082f
C439 B.n394 VSUBS 0.007082f
C440 B.n395 VSUBS 0.007082f
C441 B.n396 VSUBS 0.007082f
C442 B.n397 VSUBS 0.007082f
C443 B.n398 VSUBS 0.007082f
C444 B.n399 VSUBS 0.007082f
C445 B.n400 VSUBS 0.007082f
C446 B.n401 VSUBS 0.007082f
C447 B.n402 VSUBS 0.007082f
C448 B.n403 VSUBS 0.007082f
C449 B.n404 VSUBS 0.007082f
C450 B.n405 VSUBS 0.007082f
C451 B.n406 VSUBS 0.007082f
C452 B.n407 VSUBS 0.007082f
C453 B.n408 VSUBS 0.007082f
C454 B.n409 VSUBS 0.007082f
C455 B.n410 VSUBS 0.006665f
C456 B.n411 VSUBS 0.016407f
C457 B.n412 VSUBS 0.003957f
C458 B.n413 VSUBS 0.007082f
C459 B.n414 VSUBS 0.007082f
C460 B.n415 VSUBS 0.007082f
C461 B.n416 VSUBS 0.007082f
C462 B.n417 VSUBS 0.007082f
C463 B.n418 VSUBS 0.007082f
C464 B.n419 VSUBS 0.007082f
C465 B.n420 VSUBS 0.007082f
C466 B.n421 VSUBS 0.007082f
C467 B.n422 VSUBS 0.007082f
C468 B.n423 VSUBS 0.007082f
C469 B.n424 VSUBS 0.007082f
C470 B.n425 VSUBS 0.003957f
C471 B.n426 VSUBS 0.007082f
C472 B.n427 VSUBS 0.007082f
C473 B.n428 VSUBS 0.007082f
C474 B.n429 VSUBS 0.007082f
C475 B.n430 VSUBS 0.007082f
C476 B.n431 VSUBS 0.007082f
C477 B.n432 VSUBS 0.007082f
C478 B.n433 VSUBS 0.007082f
C479 B.n434 VSUBS 0.007082f
C480 B.n435 VSUBS 0.007082f
C481 B.n436 VSUBS 0.007082f
C482 B.n437 VSUBS 0.007082f
C483 B.n438 VSUBS 0.007082f
C484 B.n439 VSUBS 0.007082f
C485 B.n440 VSUBS 0.007082f
C486 B.n441 VSUBS 0.007082f
C487 B.n442 VSUBS 0.007082f
C488 B.n443 VSUBS 0.007082f
C489 B.n444 VSUBS 0.007082f
C490 B.n445 VSUBS 0.007082f
C491 B.n446 VSUBS 0.007082f
C492 B.n447 VSUBS 0.007082f
C493 B.n448 VSUBS 0.007082f
C494 B.n449 VSUBS 0.007082f
C495 B.n450 VSUBS 0.007082f
C496 B.n451 VSUBS 0.007082f
C497 B.n452 VSUBS 0.007082f
C498 B.n453 VSUBS 0.007082f
C499 B.n454 VSUBS 0.007082f
C500 B.n455 VSUBS 0.007082f
C501 B.n456 VSUBS 0.007082f
C502 B.n457 VSUBS 0.007082f
C503 B.n458 VSUBS 0.007082f
C504 B.n459 VSUBS 0.007082f
C505 B.n460 VSUBS 0.007082f
C506 B.n461 VSUBS 0.007082f
C507 B.n462 VSUBS 0.007082f
C508 B.n463 VSUBS 0.007082f
C509 B.n464 VSUBS 0.007082f
C510 B.n465 VSUBS 0.007082f
C511 B.n466 VSUBS 0.016832f
C512 B.n467 VSUBS 0.015451f
C513 B.n468 VSUBS 0.015451f
C514 B.n469 VSUBS 0.007082f
C515 B.n470 VSUBS 0.007082f
C516 B.n471 VSUBS 0.007082f
C517 B.n472 VSUBS 0.007082f
C518 B.n473 VSUBS 0.007082f
C519 B.n474 VSUBS 0.007082f
C520 B.n475 VSUBS 0.007082f
C521 B.n476 VSUBS 0.007082f
C522 B.n477 VSUBS 0.007082f
C523 B.n478 VSUBS 0.007082f
C524 B.n479 VSUBS 0.007082f
C525 B.n480 VSUBS 0.007082f
C526 B.n481 VSUBS 0.007082f
C527 B.n482 VSUBS 0.007082f
C528 B.n483 VSUBS 0.007082f
C529 B.n484 VSUBS 0.007082f
C530 B.n485 VSUBS 0.007082f
C531 B.n486 VSUBS 0.007082f
C532 B.n487 VSUBS 0.007082f
C533 B.n488 VSUBS 0.007082f
C534 B.n489 VSUBS 0.007082f
C535 B.n490 VSUBS 0.007082f
C536 B.n491 VSUBS 0.007082f
C537 B.n492 VSUBS 0.007082f
C538 B.n493 VSUBS 0.007082f
C539 B.n494 VSUBS 0.007082f
C540 B.n495 VSUBS 0.007082f
C541 B.n496 VSUBS 0.007082f
C542 B.n497 VSUBS 0.007082f
C543 B.n498 VSUBS 0.007082f
C544 B.n499 VSUBS 0.007082f
C545 B.n500 VSUBS 0.007082f
C546 B.n501 VSUBS 0.007082f
C547 B.n502 VSUBS 0.007082f
C548 B.n503 VSUBS 0.007082f
C549 B.n504 VSUBS 0.007082f
C550 B.n505 VSUBS 0.007082f
C551 B.n506 VSUBS 0.007082f
C552 B.n507 VSUBS 0.007082f
C553 B.n508 VSUBS 0.007082f
C554 B.n509 VSUBS 0.007082f
C555 B.n510 VSUBS 0.007082f
C556 B.n511 VSUBS 0.009241f
C557 B.n512 VSUBS 0.009844f
C558 B.n513 VSUBS 0.019576f
C559 VDD1.t0 VSUBS 1.09257f
C560 VDD1.t1 VSUBS 1.55886f
C561 VTAIL.t2 VSUBS 1.20024f
C562 VTAIL.n0 VSUBS 2.09823f
C563 VTAIL.t1 VSUBS 1.20024f
C564 VTAIL.n1 VSUBS 2.16202f
C565 VTAIL.t3 VSUBS 1.20024f
C566 VTAIL.n2 VSUBS 1.88749f
C567 VTAIL.t0 VSUBS 1.20024f
C568 VTAIL.n3 VSUBS 1.77495f
C569 VP.t1 VSUBS 3.71745f
C570 VP.t0 VSUBS 2.88985f
C571 VP.n0 VSUBS 4.05744f
.ends

