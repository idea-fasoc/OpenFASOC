* NGSPICE file created from diff_pair_sample_1513.ext - technology: sky130A

.subckt diff_pair_sample_1513 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t15 VN.t0 VDD2.t5 w_n4280_n1136# sky130_fd_pr__pfet_01v8 ad=0.3276 pd=2.46 as=0.1386 ps=1.17 w=0.84 l=2.98
X1 VDD1.t7 VP.t0 VTAIL.t1 w_n4280_n1136# sky130_fd_pr__pfet_01v8 ad=0.1386 pd=1.17 as=0.3276 ps=2.46 w=0.84 l=2.98
X2 VTAIL.t2 VP.t1 VDD1.t6 w_n4280_n1136# sky130_fd_pr__pfet_01v8 ad=0.3276 pd=2.46 as=0.1386 ps=1.17 w=0.84 l=2.98
X3 VDD2.t0 VN.t1 VTAIL.t14 w_n4280_n1136# sky130_fd_pr__pfet_01v8 ad=0.1386 pd=1.17 as=0.1386 ps=1.17 w=0.84 l=2.98
X4 VDD2.t1 VN.t2 VTAIL.t13 w_n4280_n1136# sky130_fd_pr__pfet_01v8 ad=0.1386 pd=1.17 as=0.3276 ps=2.46 w=0.84 l=2.98
X5 B.t11 B.t9 B.t10 w_n4280_n1136# sky130_fd_pr__pfet_01v8 ad=0.3276 pd=2.46 as=0 ps=0 w=0.84 l=2.98
X6 VDD1.t5 VP.t2 VTAIL.t3 w_n4280_n1136# sky130_fd_pr__pfet_01v8 ad=0.1386 pd=1.17 as=0.3276 ps=2.46 w=0.84 l=2.98
X7 VTAIL.t4 VP.t3 VDD1.t4 w_n4280_n1136# sky130_fd_pr__pfet_01v8 ad=0.1386 pd=1.17 as=0.1386 ps=1.17 w=0.84 l=2.98
X8 B.t8 B.t6 B.t7 w_n4280_n1136# sky130_fd_pr__pfet_01v8 ad=0.3276 pd=2.46 as=0 ps=0 w=0.84 l=2.98
X9 B.t5 B.t3 B.t4 w_n4280_n1136# sky130_fd_pr__pfet_01v8 ad=0.3276 pd=2.46 as=0 ps=0 w=0.84 l=2.98
X10 VTAIL.t12 VN.t3 VDD2.t3 w_n4280_n1136# sky130_fd_pr__pfet_01v8 ad=0.1386 pd=1.17 as=0.1386 ps=1.17 w=0.84 l=2.98
X11 VDD1.t3 VP.t4 VTAIL.t0 w_n4280_n1136# sky130_fd_pr__pfet_01v8 ad=0.1386 pd=1.17 as=0.1386 ps=1.17 w=0.84 l=2.98
X12 VTAIL.t6 VP.t5 VDD1.t2 w_n4280_n1136# sky130_fd_pr__pfet_01v8 ad=0.1386 pd=1.17 as=0.1386 ps=1.17 w=0.84 l=2.98
X13 VDD1.t1 VP.t6 VTAIL.t5 w_n4280_n1136# sky130_fd_pr__pfet_01v8 ad=0.1386 pd=1.17 as=0.1386 ps=1.17 w=0.84 l=2.98
X14 VDD2.t4 VN.t4 VTAIL.t11 w_n4280_n1136# sky130_fd_pr__pfet_01v8 ad=0.1386 pd=1.17 as=0.1386 ps=1.17 w=0.84 l=2.98
X15 VTAIL.t7 VP.t7 VDD1.t0 w_n4280_n1136# sky130_fd_pr__pfet_01v8 ad=0.3276 pd=2.46 as=0.1386 ps=1.17 w=0.84 l=2.98
X16 VTAIL.t10 VN.t5 VDD2.t2 w_n4280_n1136# sky130_fd_pr__pfet_01v8 ad=0.3276 pd=2.46 as=0.1386 ps=1.17 w=0.84 l=2.98
X17 B.t2 B.t0 B.t1 w_n4280_n1136# sky130_fd_pr__pfet_01v8 ad=0.3276 pd=2.46 as=0 ps=0 w=0.84 l=2.98
X18 VDD2.t6 VN.t6 VTAIL.t9 w_n4280_n1136# sky130_fd_pr__pfet_01v8 ad=0.1386 pd=1.17 as=0.3276 ps=2.46 w=0.84 l=2.98
X19 VTAIL.t8 VN.t7 VDD2.t7 w_n4280_n1136# sky130_fd_pr__pfet_01v8 ad=0.1386 pd=1.17 as=0.1386 ps=1.17 w=0.84 l=2.98
R0 VN.n60 VN.n59 161.3
R1 VN.n58 VN.n32 161.3
R2 VN.n57 VN.n56 161.3
R3 VN.n55 VN.n33 161.3
R4 VN.n54 VN.n53 161.3
R5 VN.n52 VN.n34 161.3
R6 VN.n50 VN.n49 161.3
R7 VN.n48 VN.n35 161.3
R8 VN.n47 VN.n46 161.3
R9 VN.n45 VN.n36 161.3
R10 VN.n44 VN.n43 161.3
R11 VN.n42 VN.n37 161.3
R12 VN.n41 VN.n40 161.3
R13 VN.n29 VN.n28 161.3
R14 VN.n27 VN.n1 161.3
R15 VN.n26 VN.n25 161.3
R16 VN.n24 VN.n2 161.3
R17 VN.n23 VN.n22 161.3
R18 VN.n21 VN.n3 161.3
R19 VN.n19 VN.n18 161.3
R20 VN.n17 VN.n4 161.3
R21 VN.n16 VN.n15 161.3
R22 VN.n14 VN.n5 161.3
R23 VN.n13 VN.n12 161.3
R24 VN.n11 VN.n6 161.3
R25 VN.n10 VN.n9 161.3
R26 VN.n30 VN.n0 67.3751
R27 VN.n61 VN.n31 67.3751
R28 VN.n8 VN.n7 66.4586
R29 VN.n39 VN.n38 66.4586
R30 VN.n26 VN.n2 56.5617
R31 VN.n57 VN.n33 56.5617
R32 VN VN.n61 44.5436
R33 VN.n14 VN.n13 40.577
R34 VN.n15 VN.n14 40.577
R35 VN.n45 VN.n44 40.577
R36 VN.n46 VN.n45 40.577
R37 VN.n38 VN.t2 38.6352
R38 VN.n7 VN.t0 38.6352
R39 VN.n9 VN.n6 24.5923
R40 VN.n13 VN.n6 24.5923
R41 VN.n15 VN.n4 24.5923
R42 VN.n19 VN.n4 24.5923
R43 VN.n22 VN.n21 24.5923
R44 VN.n22 VN.n2 24.5923
R45 VN.n27 VN.n26 24.5923
R46 VN.n28 VN.n27 24.5923
R47 VN.n44 VN.n37 24.5923
R48 VN.n40 VN.n37 24.5923
R49 VN.n53 VN.n33 24.5923
R50 VN.n53 VN.n52 24.5923
R51 VN.n50 VN.n35 24.5923
R52 VN.n46 VN.n35 24.5923
R53 VN.n59 VN.n58 24.5923
R54 VN.n58 VN.n57 24.5923
R55 VN.n28 VN.n0 22.8709
R56 VN.n59 VN.n31 22.8709
R57 VN.n21 VN.n20 16.9689
R58 VN.n52 VN.n51 16.9689
R59 VN.n9 VN.n8 7.62397
R60 VN.n20 VN.n19 7.62397
R61 VN.n40 VN.n39 7.62397
R62 VN.n51 VN.n50 7.62397
R63 VN.n8 VN.t1 6.79379
R64 VN.n20 VN.t7 6.79379
R65 VN.n0 VN.t6 6.79379
R66 VN.n39 VN.t3 6.79379
R67 VN.n51 VN.t4 6.79379
R68 VN.n31 VN.t5 6.79379
R69 VN.n41 VN.n38 5.33858
R70 VN.n10 VN.n7 5.33858
R71 VN.n61 VN.n60 0.354861
R72 VN.n30 VN.n29 0.354861
R73 VN VN.n30 0.267071
R74 VN.n60 VN.n32 0.189894
R75 VN.n56 VN.n32 0.189894
R76 VN.n56 VN.n55 0.189894
R77 VN.n55 VN.n54 0.189894
R78 VN.n54 VN.n34 0.189894
R79 VN.n49 VN.n34 0.189894
R80 VN.n49 VN.n48 0.189894
R81 VN.n48 VN.n47 0.189894
R82 VN.n47 VN.n36 0.189894
R83 VN.n43 VN.n36 0.189894
R84 VN.n43 VN.n42 0.189894
R85 VN.n42 VN.n41 0.189894
R86 VN.n11 VN.n10 0.189894
R87 VN.n12 VN.n11 0.189894
R88 VN.n12 VN.n5 0.189894
R89 VN.n16 VN.n5 0.189894
R90 VN.n17 VN.n16 0.189894
R91 VN.n18 VN.n17 0.189894
R92 VN.n18 VN.n3 0.189894
R93 VN.n23 VN.n3 0.189894
R94 VN.n24 VN.n23 0.189894
R95 VN.n25 VN.n24 0.189894
R96 VN.n25 VN.n1 0.189894
R97 VN.n29 VN.n1 0.189894
R98 VDD2.n2 VDD2.n1 638.4
R99 VDD2.n2 VDD2.n0 638.4
R100 VDD2 VDD2.n5 638.399
R101 VDD2.n4 VDD2.n3 637.029
R102 VDD2.n5 VDD2.t3 38.6969
R103 VDD2.n5 VDD2.t1 38.6969
R104 VDD2.n3 VDD2.t2 38.6969
R105 VDD2.n3 VDD2.t4 38.6969
R106 VDD2.n1 VDD2.t7 38.6969
R107 VDD2.n1 VDD2.t6 38.6969
R108 VDD2.n0 VDD2.t5 38.6969
R109 VDD2.n0 VDD2.t0 38.6969
R110 VDD2.n4 VDD2.n2 37.28
R111 VDD2 VDD2.n4 1.48541
R112 VTAIL.n14 VTAIL.t1 659.048
R113 VTAIL.n11 VTAIL.t7 659.048
R114 VTAIL.n10 VTAIL.t13 659.048
R115 VTAIL.n7 VTAIL.t10 659.048
R116 VTAIL.n15 VTAIL.t9 659.047
R117 VTAIL.n2 VTAIL.t15 659.047
R118 VTAIL.n3 VTAIL.t3 659.047
R119 VTAIL.n6 VTAIL.t2 659.047
R120 VTAIL.n13 VTAIL.n12 620.351
R121 VTAIL.n9 VTAIL.n8 620.351
R122 VTAIL.n1 VTAIL.n0 620.351
R123 VTAIL.n5 VTAIL.n4 620.351
R124 VTAIL.n0 VTAIL.t14 38.6969
R125 VTAIL.n0 VTAIL.t8 38.6969
R126 VTAIL.n4 VTAIL.t0 38.6969
R127 VTAIL.n4 VTAIL.t4 38.6969
R128 VTAIL.n12 VTAIL.t5 38.6969
R129 VTAIL.n12 VTAIL.t6 38.6969
R130 VTAIL.n8 VTAIL.t11 38.6969
R131 VTAIL.n8 VTAIL.t12 38.6969
R132 VTAIL.n15 VTAIL.n14 15.9445
R133 VTAIL.n7 VTAIL.n6 15.9445
R134 VTAIL.n9 VTAIL.n7 2.85395
R135 VTAIL.n10 VTAIL.n9 2.85395
R136 VTAIL.n13 VTAIL.n11 2.85395
R137 VTAIL.n14 VTAIL.n13 2.85395
R138 VTAIL.n6 VTAIL.n5 2.85395
R139 VTAIL.n5 VTAIL.n3 2.85395
R140 VTAIL.n2 VTAIL.n1 2.85395
R141 VTAIL VTAIL.n15 2.79576
R142 VTAIL.n11 VTAIL.n10 0.470328
R143 VTAIL.n3 VTAIL.n2 0.470328
R144 VTAIL VTAIL.n1 0.0586897
R145 VP.n21 VP.n20 161.3
R146 VP.n22 VP.n17 161.3
R147 VP.n24 VP.n23 161.3
R148 VP.n25 VP.n16 161.3
R149 VP.n27 VP.n26 161.3
R150 VP.n28 VP.n15 161.3
R151 VP.n30 VP.n29 161.3
R152 VP.n32 VP.n14 161.3
R153 VP.n34 VP.n33 161.3
R154 VP.n35 VP.n13 161.3
R155 VP.n37 VP.n36 161.3
R156 VP.n38 VP.n12 161.3
R157 VP.n40 VP.n39 161.3
R158 VP.n73 VP.n72 161.3
R159 VP.n71 VP.n1 161.3
R160 VP.n70 VP.n69 161.3
R161 VP.n68 VP.n2 161.3
R162 VP.n67 VP.n66 161.3
R163 VP.n65 VP.n3 161.3
R164 VP.n63 VP.n62 161.3
R165 VP.n61 VP.n4 161.3
R166 VP.n60 VP.n59 161.3
R167 VP.n58 VP.n5 161.3
R168 VP.n57 VP.n56 161.3
R169 VP.n55 VP.n6 161.3
R170 VP.n54 VP.n53 161.3
R171 VP.n51 VP.n7 161.3
R172 VP.n50 VP.n49 161.3
R173 VP.n48 VP.n8 161.3
R174 VP.n47 VP.n46 161.3
R175 VP.n45 VP.n9 161.3
R176 VP.n44 VP.n43 161.3
R177 VP.n42 VP.n10 67.3751
R178 VP.n74 VP.n0 67.3751
R179 VP.n41 VP.n11 67.3751
R180 VP.n19 VP.n18 66.4586
R181 VP.n46 VP.n8 56.5617
R182 VP.n70 VP.n2 56.5617
R183 VP.n37 VP.n13 56.5617
R184 VP.n42 VP.n41 44.3783
R185 VP.n58 VP.n57 40.577
R186 VP.n59 VP.n58 40.577
R187 VP.n26 VP.n25 40.577
R188 VP.n25 VP.n24 40.577
R189 VP.n18 VP.t7 38.6349
R190 VP.n45 VP.n44 24.5923
R191 VP.n46 VP.n45 24.5923
R192 VP.n50 VP.n8 24.5923
R193 VP.n51 VP.n50 24.5923
R194 VP.n53 VP.n6 24.5923
R195 VP.n57 VP.n6 24.5923
R196 VP.n59 VP.n4 24.5923
R197 VP.n63 VP.n4 24.5923
R198 VP.n66 VP.n65 24.5923
R199 VP.n66 VP.n2 24.5923
R200 VP.n71 VP.n70 24.5923
R201 VP.n72 VP.n71 24.5923
R202 VP.n38 VP.n37 24.5923
R203 VP.n39 VP.n38 24.5923
R204 VP.n26 VP.n15 24.5923
R205 VP.n30 VP.n15 24.5923
R206 VP.n33 VP.n32 24.5923
R207 VP.n33 VP.n13 24.5923
R208 VP.n20 VP.n17 24.5923
R209 VP.n24 VP.n17 24.5923
R210 VP.n44 VP.n10 22.8709
R211 VP.n72 VP.n0 22.8709
R212 VP.n39 VP.n11 22.8709
R213 VP.n52 VP.n51 16.9689
R214 VP.n65 VP.n64 16.9689
R215 VP.n32 VP.n31 16.9689
R216 VP.n53 VP.n52 7.62397
R217 VP.n64 VP.n63 7.62397
R218 VP.n31 VP.n30 7.62397
R219 VP.n20 VP.n19 7.62397
R220 VP.n10 VP.t1 6.79379
R221 VP.n52 VP.t4 6.79379
R222 VP.n64 VP.t3 6.79379
R223 VP.n0 VP.t2 6.79379
R224 VP.n11 VP.t0 6.79379
R225 VP.n31 VP.t5 6.79379
R226 VP.n19 VP.t6 6.79379
R227 VP.n21 VP.n18 5.33854
R228 VP.n41 VP.n40 0.354861
R229 VP.n43 VP.n42 0.354861
R230 VP.n74 VP.n73 0.354861
R231 VP VP.n74 0.267071
R232 VP.n22 VP.n21 0.189894
R233 VP.n23 VP.n22 0.189894
R234 VP.n23 VP.n16 0.189894
R235 VP.n27 VP.n16 0.189894
R236 VP.n28 VP.n27 0.189894
R237 VP.n29 VP.n28 0.189894
R238 VP.n29 VP.n14 0.189894
R239 VP.n34 VP.n14 0.189894
R240 VP.n35 VP.n34 0.189894
R241 VP.n36 VP.n35 0.189894
R242 VP.n36 VP.n12 0.189894
R243 VP.n40 VP.n12 0.189894
R244 VP.n43 VP.n9 0.189894
R245 VP.n47 VP.n9 0.189894
R246 VP.n48 VP.n47 0.189894
R247 VP.n49 VP.n48 0.189894
R248 VP.n49 VP.n7 0.189894
R249 VP.n54 VP.n7 0.189894
R250 VP.n55 VP.n54 0.189894
R251 VP.n56 VP.n55 0.189894
R252 VP.n56 VP.n5 0.189894
R253 VP.n60 VP.n5 0.189894
R254 VP.n61 VP.n60 0.189894
R255 VP.n62 VP.n61 0.189894
R256 VP.n62 VP.n3 0.189894
R257 VP.n67 VP.n3 0.189894
R258 VP.n68 VP.n67 0.189894
R259 VP.n69 VP.n68 0.189894
R260 VP.n69 VP.n1 0.189894
R261 VP.n73 VP.n1 0.189894
R262 VDD1 VDD1.n0 638.514
R263 VDD1.n3 VDD1.n2 638.4
R264 VDD1.n3 VDD1.n1 638.4
R265 VDD1.n5 VDD1.n4 637.029
R266 VDD1.n4 VDD1.t2 38.6969
R267 VDD1.n4 VDD1.t7 38.6969
R268 VDD1.n0 VDD1.t0 38.6969
R269 VDD1.n0 VDD1.t1 38.6969
R270 VDD1.n2 VDD1.t4 38.6969
R271 VDD1.n2 VDD1.t5 38.6969
R272 VDD1.n1 VDD1.t6 38.6969
R273 VDD1.n1 VDD1.t3 38.6969
R274 VDD1.n5 VDD1.n3 37.863
R275 VDD1 VDD1.n5 1.36903
R276 B.n117 B.t7 713.879
R277 B.n111 B.t4 713.879
R278 B.n43 B.t2 713.879
R279 B.n36 B.t11 713.879
R280 B.n118 B.t8 649.684
R281 B.n112 B.t5 649.684
R282 B.n44 B.t1 649.684
R283 B.n37 B.t10 649.684
R284 B.n275 B.n274 585
R285 B.n273 B.n106 585
R286 B.n272 B.n271 585
R287 B.n270 B.n107 585
R288 B.n269 B.n268 585
R289 B.n267 B.n108 585
R290 B.n266 B.n265 585
R291 B.n264 B.n109 585
R292 B.n263 B.n262 585
R293 B.n260 B.n110 585
R294 B.n259 B.n258 585
R295 B.n257 B.n113 585
R296 B.n256 B.n255 585
R297 B.n254 B.n114 585
R298 B.n253 B.n252 585
R299 B.n251 B.n115 585
R300 B.n250 B.n249 585
R301 B.n248 B.n116 585
R302 B.n246 B.n245 585
R303 B.n244 B.n119 585
R304 B.n243 B.n242 585
R305 B.n241 B.n120 585
R306 B.n240 B.n239 585
R307 B.n238 B.n121 585
R308 B.n237 B.n236 585
R309 B.n235 B.n122 585
R310 B.n234 B.n233 585
R311 B.n276 B.n105 585
R312 B.n278 B.n277 585
R313 B.n279 B.n104 585
R314 B.n281 B.n280 585
R315 B.n282 B.n103 585
R316 B.n284 B.n283 585
R317 B.n285 B.n102 585
R318 B.n287 B.n286 585
R319 B.n288 B.n101 585
R320 B.n290 B.n289 585
R321 B.n291 B.n100 585
R322 B.n293 B.n292 585
R323 B.n294 B.n99 585
R324 B.n296 B.n295 585
R325 B.n297 B.n98 585
R326 B.n299 B.n298 585
R327 B.n300 B.n97 585
R328 B.n302 B.n301 585
R329 B.n303 B.n96 585
R330 B.n305 B.n304 585
R331 B.n306 B.n95 585
R332 B.n308 B.n307 585
R333 B.n309 B.n94 585
R334 B.n311 B.n310 585
R335 B.n312 B.n93 585
R336 B.n314 B.n313 585
R337 B.n315 B.n92 585
R338 B.n317 B.n316 585
R339 B.n318 B.n91 585
R340 B.n320 B.n319 585
R341 B.n321 B.n90 585
R342 B.n323 B.n322 585
R343 B.n324 B.n89 585
R344 B.n326 B.n325 585
R345 B.n327 B.n88 585
R346 B.n329 B.n328 585
R347 B.n330 B.n87 585
R348 B.n332 B.n331 585
R349 B.n333 B.n86 585
R350 B.n335 B.n334 585
R351 B.n336 B.n85 585
R352 B.n338 B.n337 585
R353 B.n339 B.n84 585
R354 B.n341 B.n340 585
R355 B.n342 B.n83 585
R356 B.n344 B.n343 585
R357 B.n345 B.n82 585
R358 B.n347 B.n346 585
R359 B.n348 B.n81 585
R360 B.n350 B.n349 585
R361 B.n351 B.n80 585
R362 B.n353 B.n352 585
R363 B.n354 B.n79 585
R364 B.n356 B.n355 585
R365 B.n357 B.n78 585
R366 B.n359 B.n358 585
R367 B.n360 B.n77 585
R368 B.n362 B.n361 585
R369 B.n363 B.n76 585
R370 B.n365 B.n364 585
R371 B.n366 B.n75 585
R372 B.n368 B.n367 585
R373 B.n369 B.n74 585
R374 B.n371 B.n370 585
R375 B.n372 B.n73 585
R376 B.n374 B.n373 585
R377 B.n375 B.n72 585
R378 B.n377 B.n376 585
R379 B.n378 B.n71 585
R380 B.n380 B.n379 585
R381 B.n381 B.n70 585
R382 B.n383 B.n382 585
R383 B.n384 B.n69 585
R384 B.n386 B.n385 585
R385 B.n387 B.n68 585
R386 B.n389 B.n388 585
R387 B.n390 B.n67 585
R388 B.n392 B.n391 585
R389 B.n393 B.n66 585
R390 B.n395 B.n394 585
R391 B.n396 B.n65 585
R392 B.n398 B.n397 585
R393 B.n399 B.n64 585
R394 B.n401 B.n400 585
R395 B.n402 B.n63 585
R396 B.n404 B.n403 585
R397 B.n405 B.n62 585
R398 B.n407 B.n406 585
R399 B.n408 B.n61 585
R400 B.n410 B.n409 585
R401 B.n411 B.n60 585
R402 B.n413 B.n412 585
R403 B.n414 B.n59 585
R404 B.n416 B.n415 585
R405 B.n417 B.n58 585
R406 B.n419 B.n418 585
R407 B.n420 B.n57 585
R408 B.n422 B.n421 585
R409 B.n423 B.n56 585
R410 B.n425 B.n424 585
R411 B.n426 B.n55 585
R412 B.n428 B.n427 585
R413 B.n429 B.n54 585
R414 B.n431 B.n430 585
R415 B.n432 B.n53 585
R416 B.n434 B.n433 585
R417 B.n435 B.n52 585
R418 B.n437 B.n436 585
R419 B.n438 B.n51 585
R420 B.n440 B.n439 585
R421 B.n441 B.n50 585
R422 B.n443 B.n442 585
R423 B.n444 B.n49 585
R424 B.n446 B.n445 585
R425 B.n487 B.n30 585
R426 B.n486 B.n485 585
R427 B.n484 B.n31 585
R428 B.n483 B.n482 585
R429 B.n481 B.n32 585
R430 B.n480 B.n479 585
R431 B.n478 B.n33 585
R432 B.n477 B.n476 585
R433 B.n475 B.n34 585
R434 B.n474 B.n473 585
R435 B.n472 B.n35 585
R436 B.n471 B.n470 585
R437 B.n469 B.n39 585
R438 B.n468 B.n467 585
R439 B.n466 B.n40 585
R440 B.n465 B.n464 585
R441 B.n463 B.n41 585
R442 B.n462 B.n461 585
R443 B.n459 B.n42 585
R444 B.n458 B.n457 585
R445 B.n456 B.n45 585
R446 B.n455 B.n454 585
R447 B.n453 B.n46 585
R448 B.n452 B.n451 585
R449 B.n450 B.n47 585
R450 B.n449 B.n448 585
R451 B.n447 B.n48 585
R452 B.n489 B.n488 585
R453 B.n490 B.n29 585
R454 B.n492 B.n491 585
R455 B.n493 B.n28 585
R456 B.n495 B.n494 585
R457 B.n496 B.n27 585
R458 B.n498 B.n497 585
R459 B.n499 B.n26 585
R460 B.n501 B.n500 585
R461 B.n502 B.n25 585
R462 B.n504 B.n503 585
R463 B.n505 B.n24 585
R464 B.n507 B.n506 585
R465 B.n508 B.n23 585
R466 B.n510 B.n509 585
R467 B.n511 B.n22 585
R468 B.n513 B.n512 585
R469 B.n514 B.n21 585
R470 B.n516 B.n515 585
R471 B.n517 B.n20 585
R472 B.n519 B.n518 585
R473 B.n520 B.n19 585
R474 B.n522 B.n521 585
R475 B.n523 B.n18 585
R476 B.n525 B.n524 585
R477 B.n526 B.n17 585
R478 B.n528 B.n527 585
R479 B.n529 B.n16 585
R480 B.n531 B.n530 585
R481 B.n532 B.n15 585
R482 B.n534 B.n533 585
R483 B.n535 B.n14 585
R484 B.n537 B.n536 585
R485 B.n538 B.n13 585
R486 B.n540 B.n539 585
R487 B.n541 B.n12 585
R488 B.n543 B.n542 585
R489 B.n544 B.n11 585
R490 B.n546 B.n545 585
R491 B.n547 B.n10 585
R492 B.n549 B.n548 585
R493 B.n550 B.n9 585
R494 B.n552 B.n551 585
R495 B.n553 B.n8 585
R496 B.n555 B.n554 585
R497 B.n556 B.n7 585
R498 B.n558 B.n557 585
R499 B.n559 B.n6 585
R500 B.n561 B.n560 585
R501 B.n562 B.n5 585
R502 B.n564 B.n563 585
R503 B.n565 B.n4 585
R504 B.n567 B.n566 585
R505 B.n568 B.n3 585
R506 B.n570 B.n569 585
R507 B.n571 B.n0 585
R508 B.n2 B.n1 585
R509 B.n151 B.n150 585
R510 B.n153 B.n152 585
R511 B.n154 B.n149 585
R512 B.n156 B.n155 585
R513 B.n157 B.n148 585
R514 B.n159 B.n158 585
R515 B.n160 B.n147 585
R516 B.n162 B.n161 585
R517 B.n163 B.n146 585
R518 B.n165 B.n164 585
R519 B.n166 B.n145 585
R520 B.n168 B.n167 585
R521 B.n169 B.n144 585
R522 B.n171 B.n170 585
R523 B.n172 B.n143 585
R524 B.n174 B.n173 585
R525 B.n175 B.n142 585
R526 B.n177 B.n176 585
R527 B.n178 B.n141 585
R528 B.n180 B.n179 585
R529 B.n181 B.n140 585
R530 B.n183 B.n182 585
R531 B.n184 B.n139 585
R532 B.n186 B.n185 585
R533 B.n187 B.n138 585
R534 B.n189 B.n188 585
R535 B.n190 B.n137 585
R536 B.n192 B.n191 585
R537 B.n193 B.n136 585
R538 B.n195 B.n194 585
R539 B.n196 B.n135 585
R540 B.n198 B.n197 585
R541 B.n199 B.n134 585
R542 B.n201 B.n200 585
R543 B.n202 B.n133 585
R544 B.n204 B.n203 585
R545 B.n205 B.n132 585
R546 B.n207 B.n206 585
R547 B.n208 B.n131 585
R548 B.n210 B.n209 585
R549 B.n211 B.n130 585
R550 B.n213 B.n212 585
R551 B.n214 B.n129 585
R552 B.n216 B.n215 585
R553 B.n217 B.n128 585
R554 B.n219 B.n218 585
R555 B.n220 B.n127 585
R556 B.n222 B.n221 585
R557 B.n223 B.n126 585
R558 B.n225 B.n224 585
R559 B.n226 B.n125 585
R560 B.n228 B.n227 585
R561 B.n229 B.n124 585
R562 B.n231 B.n230 585
R563 B.n232 B.n123 585
R564 B.n233 B.n232 559.769
R565 B.n276 B.n275 559.769
R566 B.n445 B.n48 559.769
R567 B.n488 B.n487 559.769
R568 B.n573 B.n572 256.663
R569 B.n572 B.n571 235.042
R570 B.n572 B.n2 235.042
R571 B.n117 B.t6 209.466
R572 B.n111 B.t3 209.466
R573 B.n43 B.t0 209.466
R574 B.n36 B.t9 209.466
R575 B.n233 B.n122 163.367
R576 B.n237 B.n122 163.367
R577 B.n238 B.n237 163.367
R578 B.n239 B.n238 163.367
R579 B.n239 B.n120 163.367
R580 B.n243 B.n120 163.367
R581 B.n244 B.n243 163.367
R582 B.n245 B.n244 163.367
R583 B.n245 B.n116 163.367
R584 B.n250 B.n116 163.367
R585 B.n251 B.n250 163.367
R586 B.n252 B.n251 163.367
R587 B.n252 B.n114 163.367
R588 B.n256 B.n114 163.367
R589 B.n257 B.n256 163.367
R590 B.n258 B.n257 163.367
R591 B.n258 B.n110 163.367
R592 B.n263 B.n110 163.367
R593 B.n264 B.n263 163.367
R594 B.n265 B.n264 163.367
R595 B.n265 B.n108 163.367
R596 B.n269 B.n108 163.367
R597 B.n270 B.n269 163.367
R598 B.n271 B.n270 163.367
R599 B.n271 B.n106 163.367
R600 B.n275 B.n106 163.367
R601 B.n445 B.n444 163.367
R602 B.n444 B.n443 163.367
R603 B.n443 B.n50 163.367
R604 B.n439 B.n50 163.367
R605 B.n439 B.n438 163.367
R606 B.n438 B.n437 163.367
R607 B.n437 B.n52 163.367
R608 B.n433 B.n52 163.367
R609 B.n433 B.n432 163.367
R610 B.n432 B.n431 163.367
R611 B.n431 B.n54 163.367
R612 B.n427 B.n54 163.367
R613 B.n427 B.n426 163.367
R614 B.n426 B.n425 163.367
R615 B.n425 B.n56 163.367
R616 B.n421 B.n56 163.367
R617 B.n421 B.n420 163.367
R618 B.n420 B.n419 163.367
R619 B.n419 B.n58 163.367
R620 B.n415 B.n58 163.367
R621 B.n415 B.n414 163.367
R622 B.n414 B.n413 163.367
R623 B.n413 B.n60 163.367
R624 B.n409 B.n60 163.367
R625 B.n409 B.n408 163.367
R626 B.n408 B.n407 163.367
R627 B.n407 B.n62 163.367
R628 B.n403 B.n62 163.367
R629 B.n403 B.n402 163.367
R630 B.n402 B.n401 163.367
R631 B.n401 B.n64 163.367
R632 B.n397 B.n64 163.367
R633 B.n397 B.n396 163.367
R634 B.n396 B.n395 163.367
R635 B.n395 B.n66 163.367
R636 B.n391 B.n66 163.367
R637 B.n391 B.n390 163.367
R638 B.n390 B.n389 163.367
R639 B.n389 B.n68 163.367
R640 B.n385 B.n68 163.367
R641 B.n385 B.n384 163.367
R642 B.n384 B.n383 163.367
R643 B.n383 B.n70 163.367
R644 B.n379 B.n70 163.367
R645 B.n379 B.n378 163.367
R646 B.n378 B.n377 163.367
R647 B.n377 B.n72 163.367
R648 B.n373 B.n72 163.367
R649 B.n373 B.n372 163.367
R650 B.n372 B.n371 163.367
R651 B.n371 B.n74 163.367
R652 B.n367 B.n74 163.367
R653 B.n367 B.n366 163.367
R654 B.n366 B.n365 163.367
R655 B.n365 B.n76 163.367
R656 B.n361 B.n76 163.367
R657 B.n361 B.n360 163.367
R658 B.n360 B.n359 163.367
R659 B.n359 B.n78 163.367
R660 B.n355 B.n78 163.367
R661 B.n355 B.n354 163.367
R662 B.n354 B.n353 163.367
R663 B.n353 B.n80 163.367
R664 B.n349 B.n80 163.367
R665 B.n349 B.n348 163.367
R666 B.n348 B.n347 163.367
R667 B.n347 B.n82 163.367
R668 B.n343 B.n82 163.367
R669 B.n343 B.n342 163.367
R670 B.n342 B.n341 163.367
R671 B.n341 B.n84 163.367
R672 B.n337 B.n84 163.367
R673 B.n337 B.n336 163.367
R674 B.n336 B.n335 163.367
R675 B.n335 B.n86 163.367
R676 B.n331 B.n86 163.367
R677 B.n331 B.n330 163.367
R678 B.n330 B.n329 163.367
R679 B.n329 B.n88 163.367
R680 B.n325 B.n88 163.367
R681 B.n325 B.n324 163.367
R682 B.n324 B.n323 163.367
R683 B.n323 B.n90 163.367
R684 B.n319 B.n90 163.367
R685 B.n319 B.n318 163.367
R686 B.n318 B.n317 163.367
R687 B.n317 B.n92 163.367
R688 B.n313 B.n92 163.367
R689 B.n313 B.n312 163.367
R690 B.n312 B.n311 163.367
R691 B.n311 B.n94 163.367
R692 B.n307 B.n94 163.367
R693 B.n307 B.n306 163.367
R694 B.n306 B.n305 163.367
R695 B.n305 B.n96 163.367
R696 B.n301 B.n96 163.367
R697 B.n301 B.n300 163.367
R698 B.n300 B.n299 163.367
R699 B.n299 B.n98 163.367
R700 B.n295 B.n98 163.367
R701 B.n295 B.n294 163.367
R702 B.n294 B.n293 163.367
R703 B.n293 B.n100 163.367
R704 B.n289 B.n100 163.367
R705 B.n289 B.n288 163.367
R706 B.n288 B.n287 163.367
R707 B.n287 B.n102 163.367
R708 B.n283 B.n102 163.367
R709 B.n283 B.n282 163.367
R710 B.n282 B.n281 163.367
R711 B.n281 B.n104 163.367
R712 B.n277 B.n104 163.367
R713 B.n277 B.n276 163.367
R714 B.n487 B.n486 163.367
R715 B.n486 B.n31 163.367
R716 B.n482 B.n31 163.367
R717 B.n482 B.n481 163.367
R718 B.n481 B.n480 163.367
R719 B.n480 B.n33 163.367
R720 B.n476 B.n33 163.367
R721 B.n476 B.n475 163.367
R722 B.n475 B.n474 163.367
R723 B.n474 B.n35 163.367
R724 B.n470 B.n35 163.367
R725 B.n470 B.n469 163.367
R726 B.n469 B.n468 163.367
R727 B.n468 B.n40 163.367
R728 B.n464 B.n40 163.367
R729 B.n464 B.n463 163.367
R730 B.n463 B.n462 163.367
R731 B.n462 B.n42 163.367
R732 B.n457 B.n42 163.367
R733 B.n457 B.n456 163.367
R734 B.n456 B.n455 163.367
R735 B.n455 B.n46 163.367
R736 B.n451 B.n46 163.367
R737 B.n451 B.n450 163.367
R738 B.n450 B.n449 163.367
R739 B.n449 B.n48 163.367
R740 B.n488 B.n29 163.367
R741 B.n492 B.n29 163.367
R742 B.n493 B.n492 163.367
R743 B.n494 B.n493 163.367
R744 B.n494 B.n27 163.367
R745 B.n498 B.n27 163.367
R746 B.n499 B.n498 163.367
R747 B.n500 B.n499 163.367
R748 B.n500 B.n25 163.367
R749 B.n504 B.n25 163.367
R750 B.n505 B.n504 163.367
R751 B.n506 B.n505 163.367
R752 B.n506 B.n23 163.367
R753 B.n510 B.n23 163.367
R754 B.n511 B.n510 163.367
R755 B.n512 B.n511 163.367
R756 B.n512 B.n21 163.367
R757 B.n516 B.n21 163.367
R758 B.n517 B.n516 163.367
R759 B.n518 B.n517 163.367
R760 B.n518 B.n19 163.367
R761 B.n522 B.n19 163.367
R762 B.n523 B.n522 163.367
R763 B.n524 B.n523 163.367
R764 B.n524 B.n17 163.367
R765 B.n528 B.n17 163.367
R766 B.n529 B.n528 163.367
R767 B.n530 B.n529 163.367
R768 B.n530 B.n15 163.367
R769 B.n534 B.n15 163.367
R770 B.n535 B.n534 163.367
R771 B.n536 B.n535 163.367
R772 B.n536 B.n13 163.367
R773 B.n540 B.n13 163.367
R774 B.n541 B.n540 163.367
R775 B.n542 B.n541 163.367
R776 B.n542 B.n11 163.367
R777 B.n546 B.n11 163.367
R778 B.n547 B.n546 163.367
R779 B.n548 B.n547 163.367
R780 B.n548 B.n9 163.367
R781 B.n552 B.n9 163.367
R782 B.n553 B.n552 163.367
R783 B.n554 B.n553 163.367
R784 B.n554 B.n7 163.367
R785 B.n558 B.n7 163.367
R786 B.n559 B.n558 163.367
R787 B.n560 B.n559 163.367
R788 B.n560 B.n5 163.367
R789 B.n564 B.n5 163.367
R790 B.n565 B.n564 163.367
R791 B.n566 B.n565 163.367
R792 B.n566 B.n3 163.367
R793 B.n570 B.n3 163.367
R794 B.n571 B.n570 163.367
R795 B.n150 B.n2 163.367
R796 B.n153 B.n150 163.367
R797 B.n154 B.n153 163.367
R798 B.n155 B.n154 163.367
R799 B.n155 B.n148 163.367
R800 B.n159 B.n148 163.367
R801 B.n160 B.n159 163.367
R802 B.n161 B.n160 163.367
R803 B.n161 B.n146 163.367
R804 B.n165 B.n146 163.367
R805 B.n166 B.n165 163.367
R806 B.n167 B.n166 163.367
R807 B.n167 B.n144 163.367
R808 B.n171 B.n144 163.367
R809 B.n172 B.n171 163.367
R810 B.n173 B.n172 163.367
R811 B.n173 B.n142 163.367
R812 B.n177 B.n142 163.367
R813 B.n178 B.n177 163.367
R814 B.n179 B.n178 163.367
R815 B.n179 B.n140 163.367
R816 B.n183 B.n140 163.367
R817 B.n184 B.n183 163.367
R818 B.n185 B.n184 163.367
R819 B.n185 B.n138 163.367
R820 B.n189 B.n138 163.367
R821 B.n190 B.n189 163.367
R822 B.n191 B.n190 163.367
R823 B.n191 B.n136 163.367
R824 B.n195 B.n136 163.367
R825 B.n196 B.n195 163.367
R826 B.n197 B.n196 163.367
R827 B.n197 B.n134 163.367
R828 B.n201 B.n134 163.367
R829 B.n202 B.n201 163.367
R830 B.n203 B.n202 163.367
R831 B.n203 B.n132 163.367
R832 B.n207 B.n132 163.367
R833 B.n208 B.n207 163.367
R834 B.n209 B.n208 163.367
R835 B.n209 B.n130 163.367
R836 B.n213 B.n130 163.367
R837 B.n214 B.n213 163.367
R838 B.n215 B.n214 163.367
R839 B.n215 B.n128 163.367
R840 B.n219 B.n128 163.367
R841 B.n220 B.n219 163.367
R842 B.n221 B.n220 163.367
R843 B.n221 B.n126 163.367
R844 B.n225 B.n126 163.367
R845 B.n226 B.n225 163.367
R846 B.n227 B.n226 163.367
R847 B.n227 B.n124 163.367
R848 B.n231 B.n124 163.367
R849 B.n232 B.n231 163.367
R850 B.n118 B.n117 64.1944
R851 B.n112 B.n111 64.1944
R852 B.n44 B.n43 64.1944
R853 B.n37 B.n36 64.1944
R854 B.n247 B.n118 59.5399
R855 B.n261 B.n112 59.5399
R856 B.n460 B.n44 59.5399
R857 B.n38 B.n37 59.5399
R858 B.n274 B.n105 36.3712
R859 B.n489 B.n30 36.3712
R860 B.n447 B.n446 36.3712
R861 B.n234 B.n123 36.3712
R862 B B.n573 18.0485
R863 B.n490 B.n489 10.6151
R864 B.n491 B.n490 10.6151
R865 B.n491 B.n28 10.6151
R866 B.n495 B.n28 10.6151
R867 B.n496 B.n495 10.6151
R868 B.n497 B.n496 10.6151
R869 B.n497 B.n26 10.6151
R870 B.n501 B.n26 10.6151
R871 B.n502 B.n501 10.6151
R872 B.n503 B.n502 10.6151
R873 B.n503 B.n24 10.6151
R874 B.n507 B.n24 10.6151
R875 B.n508 B.n507 10.6151
R876 B.n509 B.n508 10.6151
R877 B.n509 B.n22 10.6151
R878 B.n513 B.n22 10.6151
R879 B.n514 B.n513 10.6151
R880 B.n515 B.n514 10.6151
R881 B.n515 B.n20 10.6151
R882 B.n519 B.n20 10.6151
R883 B.n520 B.n519 10.6151
R884 B.n521 B.n520 10.6151
R885 B.n521 B.n18 10.6151
R886 B.n525 B.n18 10.6151
R887 B.n526 B.n525 10.6151
R888 B.n527 B.n526 10.6151
R889 B.n527 B.n16 10.6151
R890 B.n531 B.n16 10.6151
R891 B.n532 B.n531 10.6151
R892 B.n533 B.n532 10.6151
R893 B.n533 B.n14 10.6151
R894 B.n537 B.n14 10.6151
R895 B.n538 B.n537 10.6151
R896 B.n539 B.n538 10.6151
R897 B.n539 B.n12 10.6151
R898 B.n543 B.n12 10.6151
R899 B.n544 B.n543 10.6151
R900 B.n545 B.n544 10.6151
R901 B.n545 B.n10 10.6151
R902 B.n549 B.n10 10.6151
R903 B.n550 B.n549 10.6151
R904 B.n551 B.n550 10.6151
R905 B.n551 B.n8 10.6151
R906 B.n555 B.n8 10.6151
R907 B.n556 B.n555 10.6151
R908 B.n557 B.n556 10.6151
R909 B.n557 B.n6 10.6151
R910 B.n561 B.n6 10.6151
R911 B.n562 B.n561 10.6151
R912 B.n563 B.n562 10.6151
R913 B.n563 B.n4 10.6151
R914 B.n567 B.n4 10.6151
R915 B.n568 B.n567 10.6151
R916 B.n569 B.n568 10.6151
R917 B.n569 B.n0 10.6151
R918 B.n485 B.n30 10.6151
R919 B.n485 B.n484 10.6151
R920 B.n484 B.n483 10.6151
R921 B.n483 B.n32 10.6151
R922 B.n479 B.n32 10.6151
R923 B.n479 B.n478 10.6151
R924 B.n478 B.n477 10.6151
R925 B.n477 B.n34 10.6151
R926 B.n473 B.n472 10.6151
R927 B.n472 B.n471 10.6151
R928 B.n471 B.n39 10.6151
R929 B.n467 B.n39 10.6151
R930 B.n467 B.n466 10.6151
R931 B.n466 B.n465 10.6151
R932 B.n465 B.n41 10.6151
R933 B.n461 B.n41 10.6151
R934 B.n459 B.n458 10.6151
R935 B.n458 B.n45 10.6151
R936 B.n454 B.n45 10.6151
R937 B.n454 B.n453 10.6151
R938 B.n453 B.n452 10.6151
R939 B.n452 B.n47 10.6151
R940 B.n448 B.n47 10.6151
R941 B.n448 B.n447 10.6151
R942 B.n446 B.n49 10.6151
R943 B.n442 B.n49 10.6151
R944 B.n442 B.n441 10.6151
R945 B.n441 B.n440 10.6151
R946 B.n440 B.n51 10.6151
R947 B.n436 B.n51 10.6151
R948 B.n436 B.n435 10.6151
R949 B.n435 B.n434 10.6151
R950 B.n434 B.n53 10.6151
R951 B.n430 B.n53 10.6151
R952 B.n430 B.n429 10.6151
R953 B.n429 B.n428 10.6151
R954 B.n428 B.n55 10.6151
R955 B.n424 B.n55 10.6151
R956 B.n424 B.n423 10.6151
R957 B.n423 B.n422 10.6151
R958 B.n422 B.n57 10.6151
R959 B.n418 B.n57 10.6151
R960 B.n418 B.n417 10.6151
R961 B.n417 B.n416 10.6151
R962 B.n416 B.n59 10.6151
R963 B.n412 B.n59 10.6151
R964 B.n412 B.n411 10.6151
R965 B.n411 B.n410 10.6151
R966 B.n410 B.n61 10.6151
R967 B.n406 B.n61 10.6151
R968 B.n406 B.n405 10.6151
R969 B.n405 B.n404 10.6151
R970 B.n404 B.n63 10.6151
R971 B.n400 B.n63 10.6151
R972 B.n400 B.n399 10.6151
R973 B.n399 B.n398 10.6151
R974 B.n398 B.n65 10.6151
R975 B.n394 B.n65 10.6151
R976 B.n394 B.n393 10.6151
R977 B.n393 B.n392 10.6151
R978 B.n392 B.n67 10.6151
R979 B.n388 B.n67 10.6151
R980 B.n388 B.n387 10.6151
R981 B.n387 B.n386 10.6151
R982 B.n386 B.n69 10.6151
R983 B.n382 B.n69 10.6151
R984 B.n382 B.n381 10.6151
R985 B.n381 B.n380 10.6151
R986 B.n380 B.n71 10.6151
R987 B.n376 B.n71 10.6151
R988 B.n376 B.n375 10.6151
R989 B.n375 B.n374 10.6151
R990 B.n374 B.n73 10.6151
R991 B.n370 B.n73 10.6151
R992 B.n370 B.n369 10.6151
R993 B.n369 B.n368 10.6151
R994 B.n368 B.n75 10.6151
R995 B.n364 B.n75 10.6151
R996 B.n364 B.n363 10.6151
R997 B.n363 B.n362 10.6151
R998 B.n362 B.n77 10.6151
R999 B.n358 B.n77 10.6151
R1000 B.n358 B.n357 10.6151
R1001 B.n357 B.n356 10.6151
R1002 B.n356 B.n79 10.6151
R1003 B.n352 B.n79 10.6151
R1004 B.n352 B.n351 10.6151
R1005 B.n351 B.n350 10.6151
R1006 B.n350 B.n81 10.6151
R1007 B.n346 B.n81 10.6151
R1008 B.n346 B.n345 10.6151
R1009 B.n345 B.n344 10.6151
R1010 B.n344 B.n83 10.6151
R1011 B.n340 B.n83 10.6151
R1012 B.n340 B.n339 10.6151
R1013 B.n339 B.n338 10.6151
R1014 B.n338 B.n85 10.6151
R1015 B.n334 B.n85 10.6151
R1016 B.n334 B.n333 10.6151
R1017 B.n333 B.n332 10.6151
R1018 B.n332 B.n87 10.6151
R1019 B.n328 B.n87 10.6151
R1020 B.n328 B.n327 10.6151
R1021 B.n327 B.n326 10.6151
R1022 B.n326 B.n89 10.6151
R1023 B.n322 B.n89 10.6151
R1024 B.n322 B.n321 10.6151
R1025 B.n321 B.n320 10.6151
R1026 B.n320 B.n91 10.6151
R1027 B.n316 B.n91 10.6151
R1028 B.n316 B.n315 10.6151
R1029 B.n315 B.n314 10.6151
R1030 B.n314 B.n93 10.6151
R1031 B.n310 B.n93 10.6151
R1032 B.n310 B.n309 10.6151
R1033 B.n309 B.n308 10.6151
R1034 B.n308 B.n95 10.6151
R1035 B.n304 B.n95 10.6151
R1036 B.n304 B.n303 10.6151
R1037 B.n303 B.n302 10.6151
R1038 B.n302 B.n97 10.6151
R1039 B.n298 B.n97 10.6151
R1040 B.n298 B.n297 10.6151
R1041 B.n297 B.n296 10.6151
R1042 B.n296 B.n99 10.6151
R1043 B.n292 B.n99 10.6151
R1044 B.n292 B.n291 10.6151
R1045 B.n291 B.n290 10.6151
R1046 B.n290 B.n101 10.6151
R1047 B.n286 B.n101 10.6151
R1048 B.n286 B.n285 10.6151
R1049 B.n285 B.n284 10.6151
R1050 B.n284 B.n103 10.6151
R1051 B.n280 B.n103 10.6151
R1052 B.n280 B.n279 10.6151
R1053 B.n279 B.n278 10.6151
R1054 B.n278 B.n105 10.6151
R1055 B.n151 B.n1 10.6151
R1056 B.n152 B.n151 10.6151
R1057 B.n152 B.n149 10.6151
R1058 B.n156 B.n149 10.6151
R1059 B.n157 B.n156 10.6151
R1060 B.n158 B.n157 10.6151
R1061 B.n158 B.n147 10.6151
R1062 B.n162 B.n147 10.6151
R1063 B.n163 B.n162 10.6151
R1064 B.n164 B.n163 10.6151
R1065 B.n164 B.n145 10.6151
R1066 B.n168 B.n145 10.6151
R1067 B.n169 B.n168 10.6151
R1068 B.n170 B.n169 10.6151
R1069 B.n170 B.n143 10.6151
R1070 B.n174 B.n143 10.6151
R1071 B.n175 B.n174 10.6151
R1072 B.n176 B.n175 10.6151
R1073 B.n176 B.n141 10.6151
R1074 B.n180 B.n141 10.6151
R1075 B.n181 B.n180 10.6151
R1076 B.n182 B.n181 10.6151
R1077 B.n182 B.n139 10.6151
R1078 B.n186 B.n139 10.6151
R1079 B.n187 B.n186 10.6151
R1080 B.n188 B.n187 10.6151
R1081 B.n188 B.n137 10.6151
R1082 B.n192 B.n137 10.6151
R1083 B.n193 B.n192 10.6151
R1084 B.n194 B.n193 10.6151
R1085 B.n194 B.n135 10.6151
R1086 B.n198 B.n135 10.6151
R1087 B.n199 B.n198 10.6151
R1088 B.n200 B.n199 10.6151
R1089 B.n200 B.n133 10.6151
R1090 B.n204 B.n133 10.6151
R1091 B.n205 B.n204 10.6151
R1092 B.n206 B.n205 10.6151
R1093 B.n206 B.n131 10.6151
R1094 B.n210 B.n131 10.6151
R1095 B.n211 B.n210 10.6151
R1096 B.n212 B.n211 10.6151
R1097 B.n212 B.n129 10.6151
R1098 B.n216 B.n129 10.6151
R1099 B.n217 B.n216 10.6151
R1100 B.n218 B.n217 10.6151
R1101 B.n218 B.n127 10.6151
R1102 B.n222 B.n127 10.6151
R1103 B.n223 B.n222 10.6151
R1104 B.n224 B.n223 10.6151
R1105 B.n224 B.n125 10.6151
R1106 B.n228 B.n125 10.6151
R1107 B.n229 B.n228 10.6151
R1108 B.n230 B.n229 10.6151
R1109 B.n230 B.n123 10.6151
R1110 B.n235 B.n234 10.6151
R1111 B.n236 B.n235 10.6151
R1112 B.n236 B.n121 10.6151
R1113 B.n240 B.n121 10.6151
R1114 B.n241 B.n240 10.6151
R1115 B.n242 B.n241 10.6151
R1116 B.n242 B.n119 10.6151
R1117 B.n246 B.n119 10.6151
R1118 B.n249 B.n248 10.6151
R1119 B.n249 B.n115 10.6151
R1120 B.n253 B.n115 10.6151
R1121 B.n254 B.n253 10.6151
R1122 B.n255 B.n254 10.6151
R1123 B.n255 B.n113 10.6151
R1124 B.n259 B.n113 10.6151
R1125 B.n260 B.n259 10.6151
R1126 B.n262 B.n109 10.6151
R1127 B.n266 B.n109 10.6151
R1128 B.n267 B.n266 10.6151
R1129 B.n268 B.n267 10.6151
R1130 B.n268 B.n107 10.6151
R1131 B.n272 B.n107 10.6151
R1132 B.n273 B.n272 10.6151
R1133 B.n274 B.n273 10.6151
R1134 B.n573 B.n0 8.11757
R1135 B.n573 B.n1 8.11757
R1136 B.n473 B.n38 6.5566
R1137 B.n461 B.n460 6.5566
R1138 B.n248 B.n247 6.5566
R1139 B.n261 B.n260 6.5566
R1140 B.n38 B.n34 4.05904
R1141 B.n460 B.n459 4.05904
R1142 B.n247 B.n246 4.05904
R1143 B.n262 B.n261 4.05904
C0 w_n4280_n1136# B 7.67957f
C1 VN B 1.14185f
C2 VP B 2.07583f
C3 VTAIL w_n4280_n1136# 1.67183f
C4 VN VTAIL 2.56866f
C5 VTAIL VP 2.58276f
C6 VDD1 VDD2 1.97622f
C7 VN w_n4280_n1136# 8.640559f
C8 VP w_n4280_n1136# 9.188991f
C9 VN VP 6.06439f
C10 VDD1 B 1.46398f
C11 VDD2 B 1.57273f
C12 VDD1 VTAIL 4.69096f
C13 VTAIL VDD2 4.74793f
C14 VDD1 w_n4280_n1136# 1.7714f
C15 VDD2 w_n4280_n1136# 1.90089f
C16 VDD1 VN 0.160258f
C17 VDD1 VP 1.46554f
C18 VN VDD2 1.06f
C19 VTAIL B 1.21521f
C20 VDD2 VP 0.570173f
C21 VDD2 VSUBS 1.196887f
C22 VDD1 VSUBS 1.893034f
C23 VTAIL VSUBS 0.588258f
C24 VN VSUBS 7.77965f
C25 VP VSUBS 3.357004f
C26 B VSUBS 4.20822f
C27 w_n4280_n1136# VSUBS 62.8133f
C28 B.n0 VSUBS 0.011501f
C29 B.n1 VSUBS 0.011501f
C30 B.n2 VSUBS 0.017009f
C31 B.n3 VSUBS 0.013034f
C32 B.n4 VSUBS 0.013034f
C33 B.n5 VSUBS 0.013034f
C34 B.n6 VSUBS 0.013034f
C35 B.n7 VSUBS 0.013034f
C36 B.n8 VSUBS 0.013034f
C37 B.n9 VSUBS 0.013034f
C38 B.n10 VSUBS 0.013034f
C39 B.n11 VSUBS 0.013034f
C40 B.n12 VSUBS 0.013034f
C41 B.n13 VSUBS 0.013034f
C42 B.n14 VSUBS 0.013034f
C43 B.n15 VSUBS 0.013034f
C44 B.n16 VSUBS 0.013034f
C45 B.n17 VSUBS 0.013034f
C46 B.n18 VSUBS 0.013034f
C47 B.n19 VSUBS 0.013034f
C48 B.n20 VSUBS 0.013034f
C49 B.n21 VSUBS 0.013034f
C50 B.n22 VSUBS 0.013034f
C51 B.n23 VSUBS 0.013034f
C52 B.n24 VSUBS 0.013034f
C53 B.n25 VSUBS 0.013034f
C54 B.n26 VSUBS 0.013034f
C55 B.n27 VSUBS 0.013034f
C56 B.n28 VSUBS 0.013034f
C57 B.n29 VSUBS 0.013034f
C58 B.n30 VSUBS 0.033671f
C59 B.n31 VSUBS 0.013034f
C60 B.n32 VSUBS 0.013034f
C61 B.n33 VSUBS 0.013034f
C62 B.n34 VSUBS 0.009009f
C63 B.n35 VSUBS 0.013034f
C64 B.t10 VSUBS 0.030125f
C65 B.t11 VSUBS 0.035949f
C66 B.t9 VSUBS 0.235822f
C67 B.n36 VSUBS 0.118422f
C68 B.n37 VSUBS 0.083355f
C69 B.n38 VSUBS 0.030199f
C70 B.n39 VSUBS 0.013034f
C71 B.n40 VSUBS 0.013034f
C72 B.n41 VSUBS 0.013034f
C73 B.n42 VSUBS 0.013034f
C74 B.t1 VSUBS 0.030125f
C75 B.t2 VSUBS 0.035949f
C76 B.t0 VSUBS 0.235822f
C77 B.n43 VSUBS 0.118422f
C78 B.n44 VSUBS 0.083355f
C79 B.n45 VSUBS 0.013034f
C80 B.n46 VSUBS 0.013034f
C81 B.n47 VSUBS 0.013034f
C82 B.n48 VSUBS 0.033671f
C83 B.n49 VSUBS 0.013034f
C84 B.n50 VSUBS 0.013034f
C85 B.n51 VSUBS 0.013034f
C86 B.n52 VSUBS 0.013034f
C87 B.n53 VSUBS 0.013034f
C88 B.n54 VSUBS 0.013034f
C89 B.n55 VSUBS 0.013034f
C90 B.n56 VSUBS 0.013034f
C91 B.n57 VSUBS 0.013034f
C92 B.n58 VSUBS 0.013034f
C93 B.n59 VSUBS 0.013034f
C94 B.n60 VSUBS 0.013034f
C95 B.n61 VSUBS 0.013034f
C96 B.n62 VSUBS 0.013034f
C97 B.n63 VSUBS 0.013034f
C98 B.n64 VSUBS 0.013034f
C99 B.n65 VSUBS 0.013034f
C100 B.n66 VSUBS 0.013034f
C101 B.n67 VSUBS 0.013034f
C102 B.n68 VSUBS 0.013034f
C103 B.n69 VSUBS 0.013034f
C104 B.n70 VSUBS 0.013034f
C105 B.n71 VSUBS 0.013034f
C106 B.n72 VSUBS 0.013034f
C107 B.n73 VSUBS 0.013034f
C108 B.n74 VSUBS 0.013034f
C109 B.n75 VSUBS 0.013034f
C110 B.n76 VSUBS 0.013034f
C111 B.n77 VSUBS 0.013034f
C112 B.n78 VSUBS 0.013034f
C113 B.n79 VSUBS 0.013034f
C114 B.n80 VSUBS 0.013034f
C115 B.n81 VSUBS 0.013034f
C116 B.n82 VSUBS 0.013034f
C117 B.n83 VSUBS 0.013034f
C118 B.n84 VSUBS 0.013034f
C119 B.n85 VSUBS 0.013034f
C120 B.n86 VSUBS 0.013034f
C121 B.n87 VSUBS 0.013034f
C122 B.n88 VSUBS 0.013034f
C123 B.n89 VSUBS 0.013034f
C124 B.n90 VSUBS 0.013034f
C125 B.n91 VSUBS 0.013034f
C126 B.n92 VSUBS 0.013034f
C127 B.n93 VSUBS 0.013034f
C128 B.n94 VSUBS 0.013034f
C129 B.n95 VSUBS 0.013034f
C130 B.n96 VSUBS 0.013034f
C131 B.n97 VSUBS 0.013034f
C132 B.n98 VSUBS 0.013034f
C133 B.n99 VSUBS 0.013034f
C134 B.n100 VSUBS 0.013034f
C135 B.n101 VSUBS 0.013034f
C136 B.n102 VSUBS 0.013034f
C137 B.n103 VSUBS 0.013034f
C138 B.n104 VSUBS 0.013034f
C139 B.n105 VSUBS 0.033266f
C140 B.n106 VSUBS 0.013034f
C141 B.n107 VSUBS 0.013034f
C142 B.n108 VSUBS 0.013034f
C143 B.n109 VSUBS 0.013034f
C144 B.n110 VSUBS 0.013034f
C145 B.t5 VSUBS 0.030125f
C146 B.t4 VSUBS 0.035949f
C147 B.t3 VSUBS 0.235822f
C148 B.n111 VSUBS 0.118422f
C149 B.n112 VSUBS 0.083355f
C150 B.n113 VSUBS 0.013034f
C151 B.n114 VSUBS 0.013034f
C152 B.n115 VSUBS 0.013034f
C153 B.n116 VSUBS 0.013034f
C154 B.t8 VSUBS 0.030125f
C155 B.t7 VSUBS 0.035949f
C156 B.t6 VSUBS 0.235822f
C157 B.n117 VSUBS 0.118422f
C158 B.n118 VSUBS 0.083355f
C159 B.n119 VSUBS 0.013034f
C160 B.n120 VSUBS 0.013034f
C161 B.n121 VSUBS 0.013034f
C162 B.n122 VSUBS 0.013034f
C163 B.n123 VSUBS 0.031883f
C164 B.n124 VSUBS 0.013034f
C165 B.n125 VSUBS 0.013034f
C166 B.n126 VSUBS 0.013034f
C167 B.n127 VSUBS 0.013034f
C168 B.n128 VSUBS 0.013034f
C169 B.n129 VSUBS 0.013034f
C170 B.n130 VSUBS 0.013034f
C171 B.n131 VSUBS 0.013034f
C172 B.n132 VSUBS 0.013034f
C173 B.n133 VSUBS 0.013034f
C174 B.n134 VSUBS 0.013034f
C175 B.n135 VSUBS 0.013034f
C176 B.n136 VSUBS 0.013034f
C177 B.n137 VSUBS 0.013034f
C178 B.n138 VSUBS 0.013034f
C179 B.n139 VSUBS 0.013034f
C180 B.n140 VSUBS 0.013034f
C181 B.n141 VSUBS 0.013034f
C182 B.n142 VSUBS 0.013034f
C183 B.n143 VSUBS 0.013034f
C184 B.n144 VSUBS 0.013034f
C185 B.n145 VSUBS 0.013034f
C186 B.n146 VSUBS 0.013034f
C187 B.n147 VSUBS 0.013034f
C188 B.n148 VSUBS 0.013034f
C189 B.n149 VSUBS 0.013034f
C190 B.n150 VSUBS 0.013034f
C191 B.n151 VSUBS 0.013034f
C192 B.n152 VSUBS 0.013034f
C193 B.n153 VSUBS 0.013034f
C194 B.n154 VSUBS 0.013034f
C195 B.n155 VSUBS 0.013034f
C196 B.n156 VSUBS 0.013034f
C197 B.n157 VSUBS 0.013034f
C198 B.n158 VSUBS 0.013034f
C199 B.n159 VSUBS 0.013034f
C200 B.n160 VSUBS 0.013034f
C201 B.n161 VSUBS 0.013034f
C202 B.n162 VSUBS 0.013034f
C203 B.n163 VSUBS 0.013034f
C204 B.n164 VSUBS 0.013034f
C205 B.n165 VSUBS 0.013034f
C206 B.n166 VSUBS 0.013034f
C207 B.n167 VSUBS 0.013034f
C208 B.n168 VSUBS 0.013034f
C209 B.n169 VSUBS 0.013034f
C210 B.n170 VSUBS 0.013034f
C211 B.n171 VSUBS 0.013034f
C212 B.n172 VSUBS 0.013034f
C213 B.n173 VSUBS 0.013034f
C214 B.n174 VSUBS 0.013034f
C215 B.n175 VSUBS 0.013034f
C216 B.n176 VSUBS 0.013034f
C217 B.n177 VSUBS 0.013034f
C218 B.n178 VSUBS 0.013034f
C219 B.n179 VSUBS 0.013034f
C220 B.n180 VSUBS 0.013034f
C221 B.n181 VSUBS 0.013034f
C222 B.n182 VSUBS 0.013034f
C223 B.n183 VSUBS 0.013034f
C224 B.n184 VSUBS 0.013034f
C225 B.n185 VSUBS 0.013034f
C226 B.n186 VSUBS 0.013034f
C227 B.n187 VSUBS 0.013034f
C228 B.n188 VSUBS 0.013034f
C229 B.n189 VSUBS 0.013034f
C230 B.n190 VSUBS 0.013034f
C231 B.n191 VSUBS 0.013034f
C232 B.n192 VSUBS 0.013034f
C233 B.n193 VSUBS 0.013034f
C234 B.n194 VSUBS 0.013034f
C235 B.n195 VSUBS 0.013034f
C236 B.n196 VSUBS 0.013034f
C237 B.n197 VSUBS 0.013034f
C238 B.n198 VSUBS 0.013034f
C239 B.n199 VSUBS 0.013034f
C240 B.n200 VSUBS 0.013034f
C241 B.n201 VSUBS 0.013034f
C242 B.n202 VSUBS 0.013034f
C243 B.n203 VSUBS 0.013034f
C244 B.n204 VSUBS 0.013034f
C245 B.n205 VSUBS 0.013034f
C246 B.n206 VSUBS 0.013034f
C247 B.n207 VSUBS 0.013034f
C248 B.n208 VSUBS 0.013034f
C249 B.n209 VSUBS 0.013034f
C250 B.n210 VSUBS 0.013034f
C251 B.n211 VSUBS 0.013034f
C252 B.n212 VSUBS 0.013034f
C253 B.n213 VSUBS 0.013034f
C254 B.n214 VSUBS 0.013034f
C255 B.n215 VSUBS 0.013034f
C256 B.n216 VSUBS 0.013034f
C257 B.n217 VSUBS 0.013034f
C258 B.n218 VSUBS 0.013034f
C259 B.n219 VSUBS 0.013034f
C260 B.n220 VSUBS 0.013034f
C261 B.n221 VSUBS 0.013034f
C262 B.n222 VSUBS 0.013034f
C263 B.n223 VSUBS 0.013034f
C264 B.n224 VSUBS 0.013034f
C265 B.n225 VSUBS 0.013034f
C266 B.n226 VSUBS 0.013034f
C267 B.n227 VSUBS 0.013034f
C268 B.n228 VSUBS 0.013034f
C269 B.n229 VSUBS 0.013034f
C270 B.n230 VSUBS 0.013034f
C271 B.n231 VSUBS 0.013034f
C272 B.n232 VSUBS 0.031883f
C273 B.n233 VSUBS 0.033671f
C274 B.n234 VSUBS 0.033671f
C275 B.n235 VSUBS 0.013034f
C276 B.n236 VSUBS 0.013034f
C277 B.n237 VSUBS 0.013034f
C278 B.n238 VSUBS 0.013034f
C279 B.n239 VSUBS 0.013034f
C280 B.n240 VSUBS 0.013034f
C281 B.n241 VSUBS 0.013034f
C282 B.n242 VSUBS 0.013034f
C283 B.n243 VSUBS 0.013034f
C284 B.n244 VSUBS 0.013034f
C285 B.n245 VSUBS 0.013034f
C286 B.n246 VSUBS 0.009009f
C287 B.n247 VSUBS 0.030199f
C288 B.n248 VSUBS 0.010542f
C289 B.n249 VSUBS 0.013034f
C290 B.n250 VSUBS 0.013034f
C291 B.n251 VSUBS 0.013034f
C292 B.n252 VSUBS 0.013034f
C293 B.n253 VSUBS 0.013034f
C294 B.n254 VSUBS 0.013034f
C295 B.n255 VSUBS 0.013034f
C296 B.n256 VSUBS 0.013034f
C297 B.n257 VSUBS 0.013034f
C298 B.n258 VSUBS 0.013034f
C299 B.n259 VSUBS 0.013034f
C300 B.n260 VSUBS 0.010542f
C301 B.n261 VSUBS 0.030199f
C302 B.n262 VSUBS 0.009009f
C303 B.n263 VSUBS 0.013034f
C304 B.n264 VSUBS 0.013034f
C305 B.n265 VSUBS 0.013034f
C306 B.n266 VSUBS 0.013034f
C307 B.n267 VSUBS 0.013034f
C308 B.n268 VSUBS 0.013034f
C309 B.n269 VSUBS 0.013034f
C310 B.n270 VSUBS 0.013034f
C311 B.n271 VSUBS 0.013034f
C312 B.n272 VSUBS 0.013034f
C313 B.n273 VSUBS 0.013034f
C314 B.n274 VSUBS 0.032288f
C315 B.n275 VSUBS 0.033671f
C316 B.n276 VSUBS 0.031883f
C317 B.n277 VSUBS 0.013034f
C318 B.n278 VSUBS 0.013034f
C319 B.n279 VSUBS 0.013034f
C320 B.n280 VSUBS 0.013034f
C321 B.n281 VSUBS 0.013034f
C322 B.n282 VSUBS 0.013034f
C323 B.n283 VSUBS 0.013034f
C324 B.n284 VSUBS 0.013034f
C325 B.n285 VSUBS 0.013034f
C326 B.n286 VSUBS 0.013034f
C327 B.n287 VSUBS 0.013034f
C328 B.n288 VSUBS 0.013034f
C329 B.n289 VSUBS 0.013034f
C330 B.n290 VSUBS 0.013034f
C331 B.n291 VSUBS 0.013034f
C332 B.n292 VSUBS 0.013034f
C333 B.n293 VSUBS 0.013034f
C334 B.n294 VSUBS 0.013034f
C335 B.n295 VSUBS 0.013034f
C336 B.n296 VSUBS 0.013034f
C337 B.n297 VSUBS 0.013034f
C338 B.n298 VSUBS 0.013034f
C339 B.n299 VSUBS 0.013034f
C340 B.n300 VSUBS 0.013034f
C341 B.n301 VSUBS 0.013034f
C342 B.n302 VSUBS 0.013034f
C343 B.n303 VSUBS 0.013034f
C344 B.n304 VSUBS 0.013034f
C345 B.n305 VSUBS 0.013034f
C346 B.n306 VSUBS 0.013034f
C347 B.n307 VSUBS 0.013034f
C348 B.n308 VSUBS 0.013034f
C349 B.n309 VSUBS 0.013034f
C350 B.n310 VSUBS 0.013034f
C351 B.n311 VSUBS 0.013034f
C352 B.n312 VSUBS 0.013034f
C353 B.n313 VSUBS 0.013034f
C354 B.n314 VSUBS 0.013034f
C355 B.n315 VSUBS 0.013034f
C356 B.n316 VSUBS 0.013034f
C357 B.n317 VSUBS 0.013034f
C358 B.n318 VSUBS 0.013034f
C359 B.n319 VSUBS 0.013034f
C360 B.n320 VSUBS 0.013034f
C361 B.n321 VSUBS 0.013034f
C362 B.n322 VSUBS 0.013034f
C363 B.n323 VSUBS 0.013034f
C364 B.n324 VSUBS 0.013034f
C365 B.n325 VSUBS 0.013034f
C366 B.n326 VSUBS 0.013034f
C367 B.n327 VSUBS 0.013034f
C368 B.n328 VSUBS 0.013034f
C369 B.n329 VSUBS 0.013034f
C370 B.n330 VSUBS 0.013034f
C371 B.n331 VSUBS 0.013034f
C372 B.n332 VSUBS 0.013034f
C373 B.n333 VSUBS 0.013034f
C374 B.n334 VSUBS 0.013034f
C375 B.n335 VSUBS 0.013034f
C376 B.n336 VSUBS 0.013034f
C377 B.n337 VSUBS 0.013034f
C378 B.n338 VSUBS 0.013034f
C379 B.n339 VSUBS 0.013034f
C380 B.n340 VSUBS 0.013034f
C381 B.n341 VSUBS 0.013034f
C382 B.n342 VSUBS 0.013034f
C383 B.n343 VSUBS 0.013034f
C384 B.n344 VSUBS 0.013034f
C385 B.n345 VSUBS 0.013034f
C386 B.n346 VSUBS 0.013034f
C387 B.n347 VSUBS 0.013034f
C388 B.n348 VSUBS 0.013034f
C389 B.n349 VSUBS 0.013034f
C390 B.n350 VSUBS 0.013034f
C391 B.n351 VSUBS 0.013034f
C392 B.n352 VSUBS 0.013034f
C393 B.n353 VSUBS 0.013034f
C394 B.n354 VSUBS 0.013034f
C395 B.n355 VSUBS 0.013034f
C396 B.n356 VSUBS 0.013034f
C397 B.n357 VSUBS 0.013034f
C398 B.n358 VSUBS 0.013034f
C399 B.n359 VSUBS 0.013034f
C400 B.n360 VSUBS 0.013034f
C401 B.n361 VSUBS 0.013034f
C402 B.n362 VSUBS 0.013034f
C403 B.n363 VSUBS 0.013034f
C404 B.n364 VSUBS 0.013034f
C405 B.n365 VSUBS 0.013034f
C406 B.n366 VSUBS 0.013034f
C407 B.n367 VSUBS 0.013034f
C408 B.n368 VSUBS 0.013034f
C409 B.n369 VSUBS 0.013034f
C410 B.n370 VSUBS 0.013034f
C411 B.n371 VSUBS 0.013034f
C412 B.n372 VSUBS 0.013034f
C413 B.n373 VSUBS 0.013034f
C414 B.n374 VSUBS 0.013034f
C415 B.n375 VSUBS 0.013034f
C416 B.n376 VSUBS 0.013034f
C417 B.n377 VSUBS 0.013034f
C418 B.n378 VSUBS 0.013034f
C419 B.n379 VSUBS 0.013034f
C420 B.n380 VSUBS 0.013034f
C421 B.n381 VSUBS 0.013034f
C422 B.n382 VSUBS 0.013034f
C423 B.n383 VSUBS 0.013034f
C424 B.n384 VSUBS 0.013034f
C425 B.n385 VSUBS 0.013034f
C426 B.n386 VSUBS 0.013034f
C427 B.n387 VSUBS 0.013034f
C428 B.n388 VSUBS 0.013034f
C429 B.n389 VSUBS 0.013034f
C430 B.n390 VSUBS 0.013034f
C431 B.n391 VSUBS 0.013034f
C432 B.n392 VSUBS 0.013034f
C433 B.n393 VSUBS 0.013034f
C434 B.n394 VSUBS 0.013034f
C435 B.n395 VSUBS 0.013034f
C436 B.n396 VSUBS 0.013034f
C437 B.n397 VSUBS 0.013034f
C438 B.n398 VSUBS 0.013034f
C439 B.n399 VSUBS 0.013034f
C440 B.n400 VSUBS 0.013034f
C441 B.n401 VSUBS 0.013034f
C442 B.n402 VSUBS 0.013034f
C443 B.n403 VSUBS 0.013034f
C444 B.n404 VSUBS 0.013034f
C445 B.n405 VSUBS 0.013034f
C446 B.n406 VSUBS 0.013034f
C447 B.n407 VSUBS 0.013034f
C448 B.n408 VSUBS 0.013034f
C449 B.n409 VSUBS 0.013034f
C450 B.n410 VSUBS 0.013034f
C451 B.n411 VSUBS 0.013034f
C452 B.n412 VSUBS 0.013034f
C453 B.n413 VSUBS 0.013034f
C454 B.n414 VSUBS 0.013034f
C455 B.n415 VSUBS 0.013034f
C456 B.n416 VSUBS 0.013034f
C457 B.n417 VSUBS 0.013034f
C458 B.n418 VSUBS 0.013034f
C459 B.n419 VSUBS 0.013034f
C460 B.n420 VSUBS 0.013034f
C461 B.n421 VSUBS 0.013034f
C462 B.n422 VSUBS 0.013034f
C463 B.n423 VSUBS 0.013034f
C464 B.n424 VSUBS 0.013034f
C465 B.n425 VSUBS 0.013034f
C466 B.n426 VSUBS 0.013034f
C467 B.n427 VSUBS 0.013034f
C468 B.n428 VSUBS 0.013034f
C469 B.n429 VSUBS 0.013034f
C470 B.n430 VSUBS 0.013034f
C471 B.n431 VSUBS 0.013034f
C472 B.n432 VSUBS 0.013034f
C473 B.n433 VSUBS 0.013034f
C474 B.n434 VSUBS 0.013034f
C475 B.n435 VSUBS 0.013034f
C476 B.n436 VSUBS 0.013034f
C477 B.n437 VSUBS 0.013034f
C478 B.n438 VSUBS 0.013034f
C479 B.n439 VSUBS 0.013034f
C480 B.n440 VSUBS 0.013034f
C481 B.n441 VSUBS 0.013034f
C482 B.n442 VSUBS 0.013034f
C483 B.n443 VSUBS 0.013034f
C484 B.n444 VSUBS 0.013034f
C485 B.n445 VSUBS 0.031883f
C486 B.n446 VSUBS 0.031883f
C487 B.n447 VSUBS 0.033671f
C488 B.n448 VSUBS 0.013034f
C489 B.n449 VSUBS 0.013034f
C490 B.n450 VSUBS 0.013034f
C491 B.n451 VSUBS 0.013034f
C492 B.n452 VSUBS 0.013034f
C493 B.n453 VSUBS 0.013034f
C494 B.n454 VSUBS 0.013034f
C495 B.n455 VSUBS 0.013034f
C496 B.n456 VSUBS 0.013034f
C497 B.n457 VSUBS 0.013034f
C498 B.n458 VSUBS 0.013034f
C499 B.n459 VSUBS 0.009009f
C500 B.n460 VSUBS 0.030199f
C501 B.n461 VSUBS 0.010542f
C502 B.n462 VSUBS 0.013034f
C503 B.n463 VSUBS 0.013034f
C504 B.n464 VSUBS 0.013034f
C505 B.n465 VSUBS 0.013034f
C506 B.n466 VSUBS 0.013034f
C507 B.n467 VSUBS 0.013034f
C508 B.n468 VSUBS 0.013034f
C509 B.n469 VSUBS 0.013034f
C510 B.n470 VSUBS 0.013034f
C511 B.n471 VSUBS 0.013034f
C512 B.n472 VSUBS 0.013034f
C513 B.n473 VSUBS 0.010542f
C514 B.n474 VSUBS 0.013034f
C515 B.n475 VSUBS 0.013034f
C516 B.n476 VSUBS 0.013034f
C517 B.n477 VSUBS 0.013034f
C518 B.n478 VSUBS 0.013034f
C519 B.n479 VSUBS 0.013034f
C520 B.n480 VSUBS 0.013034f
C521 B.n481 VSUBS 0.013034f
C522 B.n482 VSUBS 0.013034f
C523 B.n483 VSUBS 0.013034f
C524 B.n484 VSUBS 0.013034f
C525 B.n485 VSUBS 0.013034f
C526 B.n486 VSUBS 0.013034f
C527 B.n487 VSUBS 0.033671f
C528 B.n488 VSUBS 0.031883f
C529 B.n489 VSUBS 0.031883f
C530 B.n490 VSUBS 0.013034f
C531 B.n491 VSUBS 0.013034f
C532 B.n492 VSUBS 0.013034f
C533 B.n493 VSUBS 0.013034f
C534 B.n494 VSUBS 0.013034f
C535 B.n495 VSUBS 0.013034f
C536 B.n496 VSUBS 0.013034f
C537 B.n497 VSUBS 0.013034f
C538 B.n498 VSUBS 0.013034f
C539 B.n499 VSUBS 0.013034f
C540 B.n500 VSUBS 0.013034f
C541 B.n501 VSUBS 0.013034f
C542 B.n502 VSUBS 0.013034f
C543 B.n503 VSUBS 0.013034f
C544 B.n504 VSUBS 0.013034f
C545 B.n505 VSUBS 0.013034f
C546 B.n506 VSUBS 0.013034f
C547 B.n507 VSUBS 0.013034f
C548 B.n508 VSUBS 0.013034f
C549 B.n509 VSUBS 0.013034f
C550 B.n510 VSUBS 0.013034f
C551 B.n511 VSUBS 0.013034f
C552 B.n512 VSUBS 0.013034f
C553 B.n513 VSUBS 0.013034f
C554 B.n514 VSUBS 0.013034f
C555 B.n515 VSUBS 0.013034f
C556 B.n516 VSUBS 0.013034f
C557 B.n517 VSUBS 0.013034f
C558 B.n518 VSUBS 0.013034f
C559 B.n519 VSUBS 0.013034f
C560 B.n520 VSUBS 0.013034f
C561 B.n521 VSUBS 0.013034f
C562 B.n522 VSUBS 0.013034f
C563 B.n523 VSUBS 0.013034f
C564 B.n524 VSUBS 0.013034f
C565 B.n525 VSUBS 0.013034f
C566 B.n526 VSUBS 0.013034f
C567 B.n527 VSUBS 0.013034f
C568 B.n528 VSUBS 0.013034f
C569 B.n529 VSUBS 0.013034f
C570 B.n530 VSUBS 0.013034f
C571 B.n531 VSUBS 0.013034f
C572 B.n532 VSUBS 0.013034f
C573 B.n533 VSUBS 0.013034f
C574 B.n534 VSUBS 0.013034f
C575 B.n535 VSUBS 0.013034f
C576 B.n536 VSUBS 0.013034f
C577 B.n537 VSUBS 0.013034f
C578 B.n538 VSUBS 0.013034f
C579 B.n539 VSUBS 0.013034f
C580 B.n540 VSUBS 0.013034f
C581 B.n541 VSUBS 0.013034f
C582 B.n542 VSUBS 0.013034f
C583 B.n543 VSUBS 0.013034f
C584 B.n544 VSUBS 0.013034f
C585 B.n545 VSUBS 0.013034f
C586 B.n546 VSUBS 0.013034f
C587 B.n547 VSUBS 0.013034f
C588 B.n548 VSUBS 0.013034f
C589 B.n549 VSUBS 0.013034f
C590 B.n550 VSUBS 0.013034f
C591 B.n551 VSUBS 0.013034f
C592 B.n552 VSUBS 0.013034f
C593 B.n553 VSUBS 0.013034f
C594 B.n554 VSUBS 0.013034f
C595 B.n555 VSUBS 0.013034f
C596 B.n556 VSUBS 0.013034f
C597 B.n557 VSUBS 0.013034f
C598 B.n558 VSUBS 0.013034f
C599 B.n559 VSUBS 0.013034f
C600 B.n560 VSUBS 0.013034f
C601 B.n561 VSUBS 0.013034f
C602 B.n562 VSUBS 0.013034f
C603 B.n563 VSUBS 0.013034f
C604 B.n564 VSUBS 0.013034f
C605 B.n565 VSUBS 0.013034f
C606 B.n566 VSUBS 0.013034f
C607 B.n567 VSUBS 0.013034f
C608 B.n568 VSUBS 0.013034f
C609 B.n569 VSUBS 0.013034f
C610 B.n570 VSUBS 0.013034f
C611 B.n571 VSUBS 0.017009f
C612 B.n572 VSUBS 0.018119f
C613 B.n573 VSUBS 0.036031f
C614 VDD1.t0 VSUBS 0.012729f
C615 VDD1.t1 VSUBS 0.012729f
C616 VDD1.n0 VSUBS 0.035325f
C617 VDD1.t6 VSUBS 0.012729f
C618 VDD1.t3 VSUBS 0.012729f
C619 VDD1.n1 VSUBS 0.035237f
C620 VDD1.t4 VSUBS 0.012729f
C621 VDD1.t5 VSUBS 0.012729f
C622 VDD1.n2 VSUBS 0.035237f
C623 VDD1.n3 VSUBS 2.17266f
C624 VDD1.t2 VSUBS 0.012729f
C625 VDD1.t7 VSUBS 0.012729f
C626 VDD1.n4 VSUBS 0.034368f
C627 VDD1.n5 VSUBS 1.69867f
C628 VP.t2 VSUBS 0.300387f
C629 VP.n0 VSUBS 0.521916f
C630 VP.n1 VSUBS 0.070991f
C631 VP.n2 VSUBS 0.114981f
C632 VP.n3 VSUBS 0.070991f
C633 VP.t3 VSUBS 0.300387f
C634 VP.n4 VSUBS 0.131646f
C635 VP.n5 VSUBS 0.070991f
C636 VP.n6 VSUBS 0.131646f
C637 VP.n7 VSUBS 0.070991f
C638 VP.t4 VSUBS 0.300387f
C639 VP.n8 VSUBS 0.114981f
C640 VP.n9 VSUBS 0.070991f
C641 VP.t1 VSUBS 0.300387f
C642 VP.n10 VSUBS 0.521916f
C643 VP.t0 VSUBS 0.300387f
C644 VP.n11 VSUBS 0.521916f
C645 VP.n12 VSUBS 0.070991f
C646 VP.n13 VSUBS 0.114981f
C647 VP.n14 VSUBS 0.070991f
C648 VP.t5 VSUBS 0.300387f
C649 VP.n15 VSUBS 0.131646f
C650 VP.n16 VSUBS 0.070991f
C651 VP.n17 VSUBS 0.131646f
C652 VP.t7 VSUBS 0.88545f
C653 VP.n18 VSUBS 0.495848f
C654 VP.t6 VSUBS 0.300387f
C655 VP.n19 VSUBS 0.442827f
C656 VP.n20 VSUBS 0.086803f
C657 VP.n21 VSUBS 0.762167f
C658 VP.n22 VSUBS 0.070991f
C659 VP.n23 VSUBS 0.070991f
C660 VP.n24 VSUBS 0.14035f
C661 VP.n25 VSUBS 0.057337f
C662 VP.n26 VSUBS 0.14035f
C663 VP.n27 VSUBS 0.070991f
C664 VP.n28 VSUBS 0.070991f
C665 VP.n29 VSUBS 0.070991f
C666 VP.n30 VSUBS 0.086803f
C667 VP.n31 VSUBS 0.230993f
C668 VP.n32 VSUBS 0.111499f
C669 VP.n33 VSUBS 0.131646f
C670 VP.n34 VSUBS 0.070991f
C671 VP.n35 VSUBS 0.070991f
C672 VP.n36 VSUBS 0.070991f
C673 VP.n37 VSUBS 0.091411f
C674 VP.n38 VSUBS 0.131646f
C675 VP.n39 VSUBS 0.127096f
C676 VP.n40 VSUBS 0.114559f
C677 VP.n41 VSUBS 3.35213f
C678 VP.n42 VSUBS 3.4098f
C679 VP.n43 VSUBS 0.114559f
C680 VP.n44 VSUBS 0.127096f
C681 VP.n45 VSUBS 0.131646f
C682 VP.n46 VSUBS 0.091411f
C683 VP.n47 VSUBS 0.070991f
C684 VP.n48 VSUBS 0.070991f
C685 VP.n49 VSUBS 0.070991f
C686 VP.n50 VSUBS 0.131646f
C687 VP.n51 VSUBS 0.111499f
C688 VP.n52 VSUBS 0.230993f
C689 VP.n53 VSUBS 0.086803f
C690 VP.n54 VSUBS 0.070991f
C691 VP.n55 VSUBS 0.070991f
C692 VP.n56 VSUBS 0.070991f
C693 VP.n57 VSUBS 0.14035f
C694 VP.n58 VSUBS 0.057337f
C695 VP.n59 VSUBS 0.14035f
C696 VP.n60 VSUBS 0.070991f
C697 VP.n61 VSUBS 0.070991f
C698 VP.n62 VSUBS 0.070991f
C699 VP.n63 VSUBS 0.086803f
C700 VP.n64 VSUBS 0.230993f
C701 VP.n65 VSUBS 0.111499f
C702 VP.n66 VSUBS 0.131646f
C703 VP.n67 VSUBS 0.070991f
C704 VP.n68 VSUBS 0.070991f
C705 VP.n69 VSUBS 0.070991f
C706 VP.n70 VSUBS 0.091411f
C707 VP.n71 VSUBS 0.131646f
C708 VP.n72 VSUBS 0.127096f
C709 VP.n73 VSUBS 0.114559f
C710 VP.n74 VSUBS 0.13784f
C711 VTAIL.t14 VSUBS 0.026667f
C712 VTAIL.t8 VSUBS 0.026667f
C713 VTAIL.n0 VSUBS 0.064574f
C714 VTAIL.n1 VSUBS 0.613691f
C715 VTAIL.t15 VSUBS 0.130806f
C716 VTAIL.n2 VSUBS 0.673473f
C717 VTAIL.t3 VSUBS 0.130806f
C718 VTAIL.n3 VSUBS 0.673473f
C719 VTAIL.t0 VSUBS 0.026667f
C720 VTAIL.t4 VSUBS 0.026667f
C721 VTAIL.n4 VSUBS 0.064574f
C722 VTAIL.n5 VSUBS 0.975532f
C723 VTAIL.t2 VSUBS 0.130806f
C724 VTAIL.n6 VSUBS 1.62148f
C725 VTAIL.t10 VSUBS 0.130806f
C726 VTAIL.n7 VSUBS 1.62148f
C727 VTAIL.t11 VSUBS 0.026667f
C728 VTAIL.t12 VSUBS 0.026667f
C729 VTAIL.n8 VSUBS 0.064574f
C730 VTAIL.n9 VSUBS 0.975532f
C731 VTAIL.t13 VSUBS 0.130806f
C732 VTAIL.n10 VSUBS 0.673473f
C733 VTAIL.t7 VSUBS 0.130806f
C734 VTAIL.n11 VSUBS 0.673473f
C735 VTAIL.t5 VSUBS 0.026667f
C736 VTAIL.t6 VSUBS 0.026667f
C737 VTAIL.n12 VSUBS 0.064574f
C738 VTAIL.n13 VSUBS 0.975532f
C739 VTAIL.t1 VSUBS 0.130806f
C740 VTAIL.n14 VSUBS 1.62148f
C741 VTAIL.t9 VSUBS 0.130806f
C742 VTAIL.n15 VSUBS 1.61394f
C743 VDD2.t5 VSUBS 0.012923f
C744 VDD2.t0 VSUBS 0.012923f
C745 VDD2.n0 VSUBS 0.035776f
C746 VDD2.t7 VSUBS 0.012923f
C747 VDD2.t6 VSUBS 0.012923f
C748 VDD2.n1 VSUBS 0.035776f
C749 VDD2.n2 VSUBS 2.16535f
C750 VDD2.t2 VSUBS 0.012923f
C751 VDD2.t4 VSUBS 0.012923f
C752 VDD2.n3 VSUBS 0.034894f
C753 VDD2.n4 VSUBS 1.7006f
C754 VDD2.t3 VSUBS 0.012923f
C755 VDD2.t1 VSUBS 0.012923f
C756 VDD2.n5 VSUBS 0.035774f
C757 VN.t6 VSUBS 0.258545f
C758 VN.n0 VSUBS 0.449216f
C759 VN.n1 VSUBS 0.061102f
C760 VN.n2 VSUBS 0.098964f
C761 VN.n3 VSUBS 0.061102f
C762 VN.t7 VSUBS 0.258545f
C763 VN.n4 VSUBS 0.113308f
C764 VN.n5 VSUBS 0.061102f
C765 VN.n6 VSUBS 0.113308f
C766 VN.t0 VSUBS 0.762114f
C767 VN.n7 VSUBS 0.426778f
C768 VN.t1 VSUBS 0.258545f
C769 VN.n8 VSUBS 0.381144f
C770 VN.n9 VSUBS 0.074711f
C771 VN.n10 VSUBS 0.656f
C772 VN.n11 VSUBS 0.061102f
C773 VN.n12 VSUBS 0.061102f
C774 VN.n13 VSUBS 0.1208f
C775 VN.n14 VSUBS 0.04935f
C776 VN.n15 VSUBS 0.1208f
C777 VN.n16 VSUBS 0.061102f
C778 VN.n17 VSUBS 0.061102f
C779 VN.n18 VSUBS 0.061102f
C780 VN.n19 VSUBS 0.074711f
C781 VN.n20 VSUBS 0.198817f
C782 VN.n21 VSUBS 0.095968f
C783 VN.n22 VSUBS 0.113308f
C784 VN.n23 VSUBS 0.061102f
C785 VN.n24 VSUBS 0.061102f
C786 VN.n25 VSUBS 0.061102f
C787 VN.n26 VSUBS 0.078678f
C788 VN.n27 VSUBS 0.113308f
C789 VN.n28 VSUBS 0.109393f
C790 VN.n29 VSUBS 0.098602f
C791 VN.n30 VSUBS 0.11864f
C792 VN.t5 VSUBS 0.258545f
C793 VN.n31 VSUBS 0.449216f
C794 VN.n32 VSUBS 0.061102f
C795 VN.n33 VSUBS 0.098964f
C796 VN.n34 VSUBS 0.061102f
C797 VN.t4 VSUBS 0.258545f
C798 VN.n35 VSUBS 0.113308f
C799 VN.n36 VSUBS 0.061102f
C800 VN.n37 VSUBS 0.113308f
C801 VN.t2 VSUBS 0.762114f
C802 VN.n38 VSUBS 0.426778f
C803 VN.t3 VSUBS 0.258545f
C804 VN.n39 VSUBS 0.381144f
C805 VN.n40 VSUBS 0.074711f
C806 VN.n41 VSUBS 0.656f
C807 VN.n42 VSUBS 0.061102f
C808 VN.n43 VSUBS 0.061102f
C809 VN.n44 VSUBS 0.1208f
C810 VN.n45 VSUBS 0.04935f
C811 VN.n46 VSUBS 0.1208f
C812 VN.n47 VSUBS 0.061102f
C813 VN.n48 VSUBS 0.061102f
C814 VN.n49 VSUBS 0.061102f
C815 VN.n50 VSUBS 0.074711f
C816 VN.n51 VSUBS 0.198817f
C817 VN.n52 VSUBS 0.095968f
C818 VN.n53 VSUBS 0.113308f
C819 VN.n54 VSUBS 0.061102f
C820 VN.n55 VSUBS 0.061102f
C821 VN.n56 VSUBS 0.061102f
C822 VN.n57 VSUBS 0.078678f
C823 VN.n58 VSUBS 0.113308f
C824 VN.n59 VSUBS 0.109393f
C825 VN.n60 VSUBS 0.098602f
C826 VN.n61 VSUBS 2.91127f
.ends

