* NGSPICE file created from diff_pair_sample_1444.ext - technology: sky130A

.subckt diff_pair_sample_1444 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t19 VP.t0 VDD1.t2 B.t4 sky130_fd_pr__nfet_01v8 ad=0.58245 pd=3.86 as=0.58245 ps=3.86 w=3.53 l=3.26
X1 VDD2.t9 VN.t0 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=1.3767 pd=7.84 as=0.58245 ps=3.86 w=3.53 l=3.26
X2 VDD1.t7 VP.t1 VTAIL.t18 B.t8 sky130_fd_pr__nfet_01v8 ad=0.58245 pd=3.86 as=1.3767 ps=7.84 w=3.53 l=3.26
X3 VDD1.t3 VP.t2 VTAIL.t17 B.t1 sky130_fd_pr__nfet_01v8 ad=0.58245 pd=3.86 as=0.58245 ps=3.86 w=3.53 l=3.26
X4 B.t23 B.t21 B.t22 B.t15 sky130_fd_pr__nfet_01v8 ad=1.3767 pd=7.84 as=0 ps=0 w=3.53 l=3.26
X5 VDD1.t0 VP.t3 VTAIL.t16 B.t0 sky130_fd_pr__nfet_01v8 ad=1.3767 pd=7.84 as=0.58245 ps=3.86 w=3.53 l=3.26
X6 B.t20 B.t18 B.t19 B.t11 sky130_fd_pr__nfet_01v8 ad=1.3767 pd=7.84 as=0 ps=0 w=3.53 l=3.26
X7 VDD2.t8 VN.t1 VTAIL.t9 B.t9 sky130_fd_pr__nfet_01v8 ad=0.58245 pd=3.86 as=1.3767 ps=7.84 w=3.53 l=3.26
X8 VDD2.t7 VN.t2 VTAIL.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=0.58245 pd=3.86 as=0.58245 ps=3.86 w=3.53 l=3.26
X9 VTAIL.t15 VP.t4 VDD1.t6 B.t7 sky130_fd_pr__nfet_01v8 ad=0.58245 pd=3.86 as=0.58245 ps=3.86 w=3.53 l=3.26
X10 VTAIL.t7 VN.t3 VDD2.t6 B.t7 sky130_fd_pr__nfet_01v8 ad=0.58245 pd=3.86 as=0.58245 ps=3.86 w=3.53 l=3.26
X11 VDD2.t5 VN.t4 VTAIL.t8 B.t8 sky130_fd_pr__nfet_01v8 ad=0.58245 pd=3.86 as=1.3767 ps=7.84 w=3.53 l=3.26
X12 VTAIL.t14 VP.t5 VDD1.t9 B.t2 sky130_fd_pr__nfet_01v8 ad=0.58245 pd=3.86 as=0.58245 ps=3.86 w=3.53 l=3.26
X13 B.t17 B.t14 B.t16 B.t15 sky130_fd_pr__nfet_01v8 ad=1.3767 pd=7.84 as=0 ps=0 w=3.53 l=3.26
X14 VDD1.t5 VP.t6 VTAIL.t13 B.t9 sky130_fd_pr__nfet_01v8 ad=0.58245 pd=3.86 as=1.3767 ps=7.84 w=3.53 l=3.26
X15 VTAIL.t2 VN.t5 VDD2.t4 B.t2 sky130_fd_pr__nfet_01v8 ad=0.58245 pd=3.86 as=0.58245 ps=3.86 w=3.53 l=3.26
X16 VDD2.t3 VN.t6 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=1.3767 pd=7.84 as=0.58245 ps=3.86 w=3.53 l=3.26
X17 VDD1.t8 VP.t7 VTAIL.t12 B.t3 sky130_fd_pr__nfet_01v8 ad=1.3767 pd=7.84 as=0.58245 ps=3.86 w=3.53 l=3.26
X18 VDD2.t2 VN.t7 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=0.58245 pd=3.86 as=0.58245 ps=3.86 w=3.53 l=3.26
X19 VDD1.t1 VP.t8 VTAIL.t11 B.t5 sky130_fd_pr__nfet_01v8 ad=0.58245 pd=3.86 as=0.58245 ps=3.86 w=3.53 l=3.26
X20 VTAIL.t10 VP.t9 VDD1.t4 B.t6 sky130_fd_pr__nfet_01v8 ad=0.58245 pd=3.86 as=0.58245 ps=3.86 w=3.53 l=3.26
X21 VTAIL.t4 VN.t8 VDD2.t1 B.t4 sky130_fd_pr__nfet_01v8 ad=0.58245 pd=3.86 as=0.58245 ps=3.86 w=3.53 l=3.26
X22 B.t13 B.t10 B.t12 B.t11 sky130_fd_pr__nfet_01v8 ad=1.3767 pd=7.84 as=0 ps=0 w=3.53 l=3.26
X23 VTAIL.t6 VN.t9 VDD2.t0 B.t6 sky130_fd_pr__nfet_01v8 ad=0.58245 pd=3.86 as=0.58245 ps=3.86 w=3.53 l=3.26
R0 VP.n32 VP.n31 161.3
R1 VP.n33 VP.n28 161.3
R2 VP.n35 VP.n34 161.3
R3 VP.n36 VP.n27 161.3
R4 VP.n38 VP.n37 161.3
R5 VP.n39 VP.n26 161.3
R6 VP.n41 VP.n40 161.3
R7 VP.n42 VP.n25 161.3
R8 VP.n44 VP.n43 161.3
R9 VP.n45 VP.n24 161.3
R10 VP.n47 VP.n46 161.3
R11 VP.n48 VP.n23 161.3
R12 VP.n50 VP.n49 161.3
R13 VP.n51 VP.n22 161.3
R14 VP.n53 VP.n52 161.3
R15 VP.n55 VP.n54 161.3
R16 VP.n56 VP.n20 161.3
R17 VP.n58 VP.n57 161.3
R18 VP.n59 VP.n19 161.3
R19 VP.n61 VP.n60 161.3
R20 VP.n62 VP.n18 161.3
R21 VP.n64 VP.n63 161.3
R22 VP.n111 VP.n110 161.3
R23 VP.n109 VP.n1 161.3
R24 VP.n108 VP.n107 161.3
R25 VP.n106 VP.n2 161.3
R26 VP.n105 VP.n104 161.3
R27 VP.n103 VP.n3 161.3
R28 VP.n102 VP.n101 161.3
R29 VP.n100 VP.n99 161.3
R30 VP.n98 VP.n5 161.3
R31 VP.n97 VP.n96 161.3
R32 VP.n95 VP.n6 161.3
R33 VP.n94 VP.n93 161.3
R34 VP.n92 VP.n7 161.3
R35 VP.n91 VP.n90 161.3
R36 VP.n89 VP.n8 161.3
R37 VP.n88 VP.n87 161.3
R38 VP.n86 VP.n9 161.3
R39 VP.n85 VP.n84 161.3
R40 VP.n83 VP.n10 161.3
R41 VP.n82 VP.n81 161.3
R42 VP.n80 VP.n11 161.3
R43 VP.n79 VP.n78 161.3
R44 VP.n77 VP.n76 161.3
R45 VP.n75 VP.n13 161.3
R46 VP.n74 VP.n73 161.3
R47 VP.n72 VP.n14 161.3
R48 VP.n71 VP.n70 161.3
R49 VP.n69 VP.n15 161.3
R50 VP.n68 VP.n67 161.3
R51 VP.n66 VP.n16 81.2593
R52 VP.n112 VP.n0 81.2593
R53 VP.n65 VP.n17 81.2593
R54 VP.n30 VP.n29 70.1236
R55 VP.n30 VP.t7 58.0018
R56 VP.n85 VP.n10 56.5193
R57 VP.n93 VP.n6 56.5193
R58 VP.n46 VP.n23 56.5193
R59 VP.n38 VP.n27 56.5193
R60 VP.n74 VP.n14 51.663
R61 VP.n104 VP.n2 51.663
R62 VP.n57 VP.n19 51.663
R63 VP.n66 VP.n65 50.2986
R64 VP.n70 VP.n14 29.3238
R65 VP.n108 VP.n2 29.3238
R66 VP.n61 VP.n19 29.3238
R67 VP.n8 VP.t2 26.0965
R68 VP.n16 VP.t3 26.0965
R69 VP.n12 VP.t4 26.0965
R70 VP.n4 VP.t5 26.0965
R71 VP.n0 VP.t1 26.0965
R72 VP.n25 VP.t8 26.0965
R73 VP.n17 VP.t6 26.0965
R74 VP.n21 VP.t9 26.0965
R75 VP.n29 VP.t0 26.0965
R76 VP.n69 VP.n68 24.4675
R77 VP.n70 VP.n69 24.4675
R78 VP.n75 VP.n74 24.4675
R79 VP.n76 VP.n75 24.4675
R80 VP.n80 VP.n79 24.4675
R81 VP.n81 VP.n80 24.4675
R82 VP.n81 VP.n10 24.4675
R83 VP.n86 VP.n85 24.4675
R84 VP.n87 VP.n86 24.4675
R85 VP.n87 VP.n8 24.4675
R86 VP.n91 VP.n8 24.4675
R87 VP.n92 VP.n91 24.4675
R88 VP.n93 VP.n92 24.4675
R89 VP.n97 VP.n6 24.4675
R90 VP.n98 VP.n97 24.4675
R91 VP.n99 VP.n98 24.4675
R92 VP.n103 VP.n102 24.4675
R93 VP.n104 VP.n103 24.4675
R94 VP.n109 VP.n108 24.4675
R95 VP.n110 VP.n109 24.4675
R96 VP.n62 VP.n61 24.4675
R97 VP.n63 VP.n62 24.4675
R98 VP.n50 VP.n23 24.4675
R99 VP.n51 VP.n50 24.4675
R100 VP.n52 VP.n51 24.4675
R101 VP.n56 VP.n55 24.4675
R102 VP.n57 VP.n56 24.4675
R103 VP.n39 VP.n38 24.4675
R104 VP.n40 VP.n39 24.4675
R105 VP.n40 VP.n25 24.4675
R106 VP.n44 VP.n25 24.4675
R107 VP.n45 VP.n44 24.4675
R108 VP.n46 VP.n45 24.4675
R109 VP.n33 VP.n32 24.4675
R110 VP.n34 VP.n33 24.4675
R111 VP.n34 VP.n27 24.4675
R112 VP.n76 VP.n12 20.0634
R113 VP.n102 VP.n4 20.0634
R114 VP.n55 VP.n21 20.0634
R115 VP.n68 VP.n16 8.80862
R116 VP.n110 VP.n0 8.80862
R117 VP.n63 VP.n17 8.80862
R118 VP.n31 VP.n30 4.46391
R119 VP.n79 VP.n12 4.40456
R120 VP.n99 VP.n4 4.40456
R121 VP.n52 VP.n21 4.40456
R122 VP.n32 VP.n29 4.40456
R123 VP.n65 VP.n64 0.354971
R124 VP.n67 VP.n66 0.354971
R125 VP.n112 VP.n111 0.354971
R126 VP VP.n112 0.26696
R127 VP.n31 VP.n28 0.189894
R128 VP.n35 VP.n28 0.189894
R129 VP.n36 VP.n35 0.189894
R130 VP.n37 VP.n36 0.189894
R131 VP.n37 VP.n26 0.189894
R132 VP.n41 VP.n26 0.189894
R133 VP.n42 VP.n41 0.189894
R134 VP.n43 VP.n42 0.189894
R135 VP.n43 VP.n24 0.189894
R136 VP.n47 VP.n24 0.189894
R137 VP.n48 VP.n47 0.189894
R138 VP.n49 VP.n48 0.189894
R139 VP.n49 VP.n22 0.189894
R140 VP.n53 VP.n22 0.189894
R141 VP.n54 VP.n53 0.189894
R142 VP.n54 VP.n20 0.189894
R143 VP.n58 VP.n20 0.189894
R144 VP.n59 VP.n58 0.189894
R145 VP.n60 VP.n59 0.189894
R146 VP.n60 VP.n18 0.189894
R147 VP.n64 VP.n18 0.189894
R148 VP.n67 VP.n15 0.189894
R149 VP.n71 VP.n15 0.189894
R150 VP.n72 VP.n71 0.189894
R151 VP.n73 VP.n72 0.189894
R152 VP.n73 VP.n13 0.189894
R153 VP.n77 VP.n13 0.189894
R154 VP.n78 VP.n77 0.189894
R155 VP.n78 VP.n11 0.189894
R156 VP.n82 VP.n11 0.189894
R157 VP.n83 VP.n82 0.189894
R158 VP.n84 VP.n83 0.189894
R159 VP.n84 VP.n9 0.189894
R160 VP.n88 VP.n9 0.189894
R161 VP.n89 VP.n88 0.189894
R162 VP.n90 VP.n89 0.189894
R163 VP.n90 VP.n7 0.189894
R164 VP.n94 VP.n7 0.189894
R165 VP.n95 VP.n94 0.189894
R166 VP.n96 VP.n95 0.189894
R167 VP.n96 VP.n5 0.189894
R168 VP.n100 VP.n5 0.189894
R169 VP.n101 VP.n100 0.189894
R170 VP.n101 VP.n3 0.189894
R171 VP.n105 VP.n3 0.189894
R172 VP.n106 VP.n105 0.189894
R173 VP.n107 VP.n106 0.189894
R174 VP.n107 VP.n1 0.189894
R175 VP.n111 VP.n1 0.189894
R176 VDD1.n1 VDD1.t8 85.0341
R177 VDD1.n3 VDD1.t0 85.0341
R178 VDD1.n5 VDD1.n4 78.5959
R179 VDD1.n1 VDD1.n0 76.3303
R180 VDD1.n7 VDD1.n6 76.3302
R181 VDD1.n3 VDD1.n2 76.3301
R182 VDD1.n7 VDD1.n5 43.5893
R183 VDD1.n6 VDD1.t4 5.60957
R184 VDD1.n6 VDD1.t5 5.60957
R185 VDD1.n0 VDD1.t2 5.60957
R186 VDD1.n0 VDD1.t1 5.60957
R187 VDD1.n4 VDD1.t9 5.60957
R188 VDD1.n4 VDD1.t7 5.60957
R189 VDD1.n2 VDD1.t6 5.60957
R190 VDD1.n2 VDD1.t3 5.60957
R191 VDD1 VDD1.n7 2.26343
R192 VDD1 VDD1.n1 0.832397
R193 VDD1.n5 VDD1.n3 0.718861
R194 VTAIL.n11 VTAIL.t8 65.2605
R195 VTAIL.n17 VTAIL.t9 65.2605
R196 VTAIL.n2 VTAIL.t18 65.2605
R197 VTAIL.n16 VTAIL.t13 65.2605
R198 VTAIL.n15 VTAIL.n14 59.6516
R199 VTAIL.n13 VTAIL.n12 59.6516
R200 VTAIL.n10 VTAIL.n9 59.6516
R201 VTAIL.n8 VTAIL.n7 59.6516
R202 VTAIL.n19 VTAIL.n18 59.6513
R203 VTAIL.n1 VTAIL.n0 59.6513
R204 VTAIL.n4 VTAIL.n3 59.6513
R205 VTAIL.n6 VTAIL.n5 59.6513
R206 VTAIL.n8 VTAIL.n6 21.5996
R207 VTAIL.n17 VTAIL.n16 18.5048
R208 VTAIL.n18 VTAIL.t5 5.60957
R209 VTAIL.n18 VTAIL.t6 5.60957
R210 VTAIL.n0 VTAIL.t3 5.60957
R211 VTAIL.n0 VTAIL.t4 5.60957
R212 VTAIL.n3 VTAIL.t17 5.60957
R213 VTAIL.n3 VTAIL.t14 5.60957
R214 VTAIL.n5 VTAIL.t16 5.60957
R215 VTAIL.n5 VTAIL.t15 5.60957
R216 VTAIL.n14 VTAIL.t11 5.60957
R217 VTAIL.n14 VTAIL.t10 5.60957
R218 VTAIL.n12 VTAIL.t12 5.60957
R219 VTAIL.n12 VTAIL.t19 5.60957
R220 VTAIL.n9 VTAIL.t1 5.60957
R221 VTAIL.n9 VTAIL.t2 5.60957
R222 VTAIL.n7 VTAIL.t0 5.60957
R223 VTAIL.n7 VTAIL.t7 5.60957
R224 VTAIL.n10 VTAIL.n8 3.09533
R225 VTAIL.n11 VTAIL.n10 3.09533
R226 VTAIL.n15 VTAIL.n13 3.09533
R227 VTAIL.n16 VTAIL.n15 3.09533
R228 VTAIL.n6 VTAIL.n4 3.09533
R229 VTAIL.n4 VTAIL.n2 3.09533
R230 VTAIL.n19 VTAIL.n17 3.09533
R231 VTAIL VTAIL.n1 2.37981
R232 VTAIL.n13 VTAIL.n11 2.01774
R233 VTAIL.n2 VTAIL.n1 2.01774
R234 VTAIL VTAIL.n19 0.716017
R235 B.n797 B.n796 585
R236 B.n798 B.n797 585
R237 B.n238 B.n152 585
R238 B.n237 B.n236 585
R239 B.n235 B.n234 585
R240 B.n233 B.n232 585
R241 B.n231 B.n230 585
R242 B.n229 B.n228 585
R243 B.n227 B.n226 585
R244 B.n225 B.n224 585
R245 B.n223 B.n222 585
R246 B.n221 B.n220 585
R247 B.n219 B.n218 585
R248 B.n217 B.n216 585
R249 B.n215 B.n214 585
R250 B.n213 B.n212 585
R251 B.n211 B.n210 585
R252 B.n209 B.n208 585
R253 B.n207 B.n206 585
R254 B.n205 B.n204 585
R255 B.n203 B.n202 585
R256 B.n201 B.n200 585
R257 B.n199 B.n198 585
R258 B.n197 B.n196 585
R259 B.n195 B.n194 585
R260 B.n193 B.n192 585
R261 B.n191 B.n190 585
R262 B.n188 B.n187 585
R263 B.n186 B.n185 585
R264 B.n184 B.n183 585
R265 B.n182 B.n181 585
R266 B.n180 B.n179 585
R267 B.n178 B.n177 585
R268 B.n176 B.n175 585
R269 B.n174 B.n173 585
R270 B.n172 B.n171 585
R271 B.n170 B.n169 585
R272 B.n168 B.n167 585
R273 B.n166 B.n165 585
R274 B.n164 B.n163 585
R275 B.n162 B.n161 585
R276 B.n160 B.n159 585
R277 B.n131 B.n130 585
R278 B.n801 B.n800 585
R279 B.n795 B.n153 585
R280 B.n153 B.n128 585
R281 B.n794 B.n127 585
R282 B.n805 B.n127 585
R283 B.n793 B.n126 585
R284 B.n806 B.n126 585
R285 B.n792 B.n125 585
R286 B.n807 B.n125 585
R287 B.n791 B.n790 585
R288 B.n790 B.n121 585
R289 B.n789 B.n120 585
R290 B.n813 B.n120 585
R291 B.n788 B.n119 585
R292 B.n814 B.n119 585
R293 B.n787 B.n118 585
R294 B.n815 B.n118 585
R295 B.n786 B.n785 585
R296 B.n785 B.n117 585
R297 B.n784 B.n113 585
R298 B.n821 B.n113 585
R299 B.n783 B.n112 585
R300 B.n822 B.n112 585
R301 B.n782 B.n111 585
R302 B.n823 B.n111 585
R303 B.n781 B.n780 585
R304 B.n780 B.n107 585
R305 B.n779 B.n106 585
R306 B.n829 B.n106 585
R307 B.n778 B.n105 585
R308 B.n830 B.n105 585
R309 B.n777 B.n104 585
R310 B.n831 B.n104 585
R311 B.n776 B.n775 585
R312 B.n775 B.n100 585
R313 B.n774 B.n99 585
R314 B.n837 B.n99 585
R315 B.n773 B.n98 585
R316 B.n838 B.n98 585
R317 B.n772 B.n97 585
R318 B.n839 B.n97 585
R319 B.n771 B.n770 585
R320 B.n770 B.n93 585
R321 B.n769 B.n92 585
R322 B.n845 B.n92 585
R323 B.n768 B.n91 585
R324 B.n846 B.n91 585
R325 B.n767 B.n90 585
R326 B.n847 B.n90 585
R327 B.n766 B.n765 585
R328 B.n765 B.n86 585
R329 B.n764 B.n85 585
R330 B.n853 B.n85 585
R331 B.n763 B.n84 585
R332 B.n854 B.n84 585
R333 B.n762 B.n83 585
R334 B.n855 B.n83 585
R335 B.n761 B.n760 585
R336 B.n760 B.n79 585
R337 B.n759 B.n78 585
R338 B.n861 B.n78 585
R339 B.n758 B.n77 585
R340 B.n862 B.n77 585
R341 B.n757 B.n76 585
R342 B.n863 B.n76 585
R343 B.n756 B.n755 585
R344 B.n755 B.n75 585
R345 B.n754 B.n71 585
R346 B.n869 B.n71 585
R347 B.n753 B.n70 585
R348 B.n870 B.n70 585
R349 B.n752 B.n69 585
R350 B.n871 B.n69 585
R351 B.n751 B.n750 585
R352 B.n750 B.n65 585
R353 B.n749 B.n64 585
R354 B.n877 B.n64 585
R355 B.n748 B.n63 585
R356 B.n878 B.n63 585
R357 B.n747 B.n62 585
R358 B.n879 B.n62 585
R359 B.n746 B.n745 585
R360 B.n745 B.n58 585
R361 B.n744 B.n57 585
R362 B.n885 B.n57 585
R363 B.n743 B.n56 585
R364 B.n886 B.n56 585
R365 B.n742 B.n55 585
R366 B.n887 B.n55 585
R367 B.n741 B.n740 585
R368 B.n740 B.n51 585
R369 B.n739 B.n50 585
R370 B.n893 B.n50 585
R371 B.n738 B.n49 585
R372 B.n894 B.n49 585
R373 B.n737 B.n48 585
R374 B.n895 B.n48 585
R375 B.n736 B.n735 585
R376 B.n735 B.n44 585
R377 B.n734 B.n43 585
R378 B.n901 B.n43 585
R379 B.n733 B.n42 585
R380 B.n902 B.n42 585
R381 B.n732 B.n41 585
R382 B.n903 B.n41 585
R383 B.n731 B.n730 585
R384 B.n730 B.n37 585
R385 B.n729 B.n36 585
R386 B.n909 B.n36 585
R387 B.n728 B.n35 585
R388 B.n910 B.n35 585
R389 B.n727 B.n34 585
R390 B.n911 B.n34 585
R391 B.n726 B.n725 585
R392 B.n725 B.n30 585
R393 B.n724 B.n29 585
R394 B.n917 B.n29 585
R395 B.n723 B.n28 585
R396 B.n918 B.n28 585
R397 B.n722 B.n27 585
R398 B.n919 B.n27 585
R399 B.n721 B.n720 585
R400 B.n720 B.n23 585
R401 B.n719 B.n22 585
R402 B.n925 B.n22 585
R403 B.n718 B.n21 585
R404 B.n926 B.n21 585
R405 B.n717 B.n20 585
R406 B.n927 B.n20 585
R407 B.n716 B.n715 585
R408 B.n715 B.n19 585
R409 B.n714 B.n15 585
R410 B.n933 B.n15 585
R411 B.n713 B.n14 585
R412 B.n934 B.n14 585
R413 B.n712 B.n13 585
R414 B.n935 B.n13 585
R415 B.n711 B.n710 585
R416 B.n710 B.n12 585
R417 B.n709 B.n708 585
R418 B.n709 B.n8 585
R419 B.n707 B.n7 585
R420 B.n942 B.n7 585
R421 B.n706 B.n6 585
R422 B.n943 B.n6 585
R423 B.n705 B.n5 585
R424 B.n944 B.n5 585
R425 B.n704 B.n703 585
R426 B.n703 B.n4 585
R427 B.n702 B.n239 585
R428 B.n702 B.n701 585
R429 B.n692 B.n240 585
R430 B.n241 B.n240 585
R431 B.n694 B.n693 585
R432 B.n695 B.n694 585
R433 B.n691 B.n246 585
R434 B.n246 B.n245 585
R435 B.n690 B.n689 585
R436 B.n689 B.n688 585
R437 B.n248 B.n247 585
R438 B.n681 B.n248 585
R439 B.n680 B.n679 585
R440 B.n682 B.n680 585
R441 B.n678 B.n253 585
R442 B.n253 B.n252 585
R443 B.n677 B.n676 585
R444 B.n676 B.n675 585
R445 B.n255 B.n254 585
R446 B.n256 B.n255 585
R447 B.n668 B.n667 585
R448 B.n669 B.n668 585
R449 B.n666 B.n261 585
R450 B.n261 B.n260 585
R451 B.n665 B.n664 585
R452 B.n664 B.n663 585
R453 B.n263 B.n262 585
R454 B.n264 B.n263 585
R455 B.n656 B.n655 585
R456 B.n657 B.n656 585
R457 B.n654 B.n268 585
R458 B.n272 B.n268 585
R459 B.n653 B.n652 585
R460 B.n652 B.n651 585
R461 B.n270 B.n269 585
R462 B.n271 B.n270 585
R463 B.n644 B.n643 585
R464 B.n645 B.n644 585
R465 B.n642 B.n277 585
R466 B.n277 B.n276 585
R467 B.n641 B.n640 585
R468 B.n640 B.n639 585
R469 B.n279 B.n278 585
R470 B.n280 B.n279 585
R471 B.n632 B.n631 585
R472 B.n633 B.n632 585
R473 B.n630 B.n285 585
R474 B.n285 B.n284 585
R475 B.n629 B.n628 585
R476 B.n628 B.n627 585
R477 B.n287 B.n286 585
R478 B.n288 B.n287 585
R479 B.n620 B.n619 585
R480 B.n621 B.n620 585
R481 B.n618 B.n293 585
R482 B.n293 B.n292 585
R483 B.n617 B.n616 585
R484 B.n616 B.n615 585
R485 B.n295 B.n294 585
R486 B.n296 B.n295 585
R487 B.n608 B.n607 585
R488 B.n609 B.n608 585
R489 B.n606 B.n301 585
R490 B.n301 B.n300 585
R491 B.n605 B.n604 585
R492 B.n604 B.n603 585
R493 B.n303 B.n302 585
R494 B.n304 B.n303 585
R495 B.n596 B.n595 585
R496 B.n597 B.n596 585
R497 B.n594 B.n309 585
R498 B.n309 B.n308 585
R499 B.n593 B.n592 585
R500 B.n592 B.n591 585
R501 B.n311 B.n310 585
R502 B.n584 B.n311 585
R503 B.n583 B.n582 585
R504 B.n585 B.n583 585
R505 B.n581 B.n316 585
R506 B.n316 B.n315 585
R507 B.n580 B.n579 585
R508 B.n579 B.n578 585
R509 B.n318 B.n317 585
R510 B.n319 B.n318 585
R511 B.n571 B.n570 585
R512 B.n572 B.n571 585
R513 B.n569 B.n324 585
R514 B.n324 B.n323 585
R515 B.n568 B.n567 585
R516 B.n567 B.n566 585
R517 B.n326 B.n325 585
R518 B.n327 B.n326 585
R519 B.n559 B.n558 585
R520 B.n560 B.n559 585
R521 B.n557 B.n331 585
R522 B.n335 B.n331 585
R523 B.n556 B.n555 585
R524 B.n555 B.n554 585
R525 B.n333 B.n332 585
R526 B.n334 B.n333 585
R527 B.n547 B.n546 585
R528 B.n548 B.n547 585
R529 B.n545 B.n340 585
R530 B.n340 B.n339 585
R531 B.n544 B.n543 585
R532 B.n543 B.n542 585
R533 B.n342 B.n341 585
R534 B.n343 B.n342 585
R535 B.n535 B.n534 585
R536 B.n536 B.n535 585
R537 B.n533 B.n348 585
R538 B.n348 B.n347 585
R539 B.n532 B.n531 585
R540 B.n531 B.n530 585
R541 B.n350 B.n349 585
R542 B.n351 B.n350 585
R543 B.n523 B.n522 585
R544 B.n524 B.n523 585
R545 B.n521 B.n356 585
R546 B.n356 B.n355 585
R547 B.n520 B.n519 585
R548 B.n519 B.n518 585
R549 B.n358 B.n357 585
R550 B.n511 B.n358 585
R551 B.n510 B.n509 585
R552 B.n512 B.n510 585
R553 B.n508 B.n363 585
R554 B.n363 B.n362 585
R555 B.n507 B.n506 585
R556 B.n506 B.n505 585
R557 B.n365 B.n364 585
R558 B.n366 B.n365 585
R559 B.n498 B.n497 585
R560 B.n499 B.n498 585
R561 B.n496 B.n371 585
R562 B.n371 B.n370 585
R563 B.n495 B.n494 585
R564 B.n494 B.n493 585
R565 B.n373 B.n372 585
R566 B.n374 B.n373 585
R567 B.n489 B.n488 585
R568 B.n377 B.n376 585
R569 B.n485 B.n484 585
R570 B.n486 B.n485 585
R571 B.n483 B.n398 585
R572 B.n482 B.n481 585
R573 B.n480 B.n479 585
R574 B.n478 B.n477 585
R575 B.n476 B.n475 585
R576 B.n474 B.n473 585
R577 B.n472 B.n471 585
R578 B.n470 B.n469 585
R579 B.n468 B.n467 585
R580 B.n466 B.n465 585
R581 B.n464 B.n463 585
R582 B.n462 B.n461 585
R583 B.n460 B.n459 585
R584 B.n458 B.n457 585
R585 B.n456 B.n455 585
R586 B.n454 B.n453 585
R587 B.n452 B.n451 585
R588 B.n450 B.n449 585
R589 B.n448 B.n447 585
R590 B.n446 B.n445 585
R591 B.n444 B.n443 585
R592 B.n442 B.n441 585
R593 B.n440 B.n439 585
R594 B.n437 B.n436 585
R595 B.n435 B.n434 585
R596 B.n433 B.n432 585
R597 B.n431 B.n430 585
R598 B.n429 B.n428 585
R599 B.n427 B.n426 585
R600 B.n425 B.n424 585
R601 B.n423 B.n422 585
R602 B.n421 B.n420 585
R603 B.n419 B.n418 585
R604 B.n417 B.n416 585
R605 B.n415 B.n414 585
R606 B.n413 B.n412 585
R607 B.n411 B.n410 585
R608 B.n409 B.n408 585
R609 B.n407 B.n406 585
R610 B.n405 B.n404 585
R611 B.n490 B.n375 585
R612 B.n375 B.n374 585
R613 B.n492 B.n491 585
R614 B.n493 B.n492 585
R615 B.n369 B.n368 585
R616 B.n370 B.n369 585
R617 B.n501 B.n500 585
R618 B.n500 B.n499 585
R619 B.n502 B.n367 585
R620 B.n367 B.n366 585
R621 B.n504 B.n503 585
R622 B.n505 B.n504 585
R623 B.n361 B.n360 585
R624 B.n362 B.n361 585
R625 B.n514 B.n513 585
R626 B.n513 B.n512 585
R627 B.n515 B.n359 585
R628 B.n511 B.n359 585
R629 B.n517 B.n516 585
R630 B.n518 B.n517 585
R631 B.n354 B.n353 585
R632 B.n355 B.n354 585
R633 B.n526 B.n525 585
R634 B.n525 B.n524 585
R635 B.n527 B.n352 585
R636 B.n352 B.n351 585
R637 B.n529 B.n528 585
R638 B.n530 B.n529 585
R639 B.n346 B.n345 585
R640 B.n347 B.n346 585
R641 B.n538 B.n537 585
R642 B.n537 B.n536 585
R643 B.n539 B.n344 585
R644 B.n344 B.n343 585
R645 B.n541 B.n540 585
R646 B.n542 B.n541 585
R647 B.n338 B.n337 585
R648 B.n339 B.n338 585
R649 B.n550 B.n549 585
R650 B.n549 B.n548 585
R651 B.n551 B.n336 585
R652 B.n336 B.n334 585
R653 B.n553 B.n552 585
R654 B.n554 B.n553 585
R655 B.n330 B.n329 585
R656 B.n335 B.n330 585
R657 B.n562 B.n561 585
R658 B.n561 B.n560 585
R659 B.n563 B.n328 585
R660 B.n328 B.n327 585
R661 B.n565 B.n564 585
R662 B.n566 B.n565 585
R663 B.n322 B.n321 585
R664 B.n323 B.n322 585
R665 B.n574 B.n573 585
R666 B.n573 B.n572 585
R667 B.n575 B.n320 585
R668 B.n320 B.n319 585
R669 B.n577 B.n576 585
R670 B.n578 B.n577 585
R671 B.n314 B.n313 585
R672 B.n315 B.n314 585
R673 B.n587 B.n586 585
R674 B.n586 B.n585 585
R675 B.n588 B.n312 585
R676 B.n584 B.n312 585
R677 B.n590 B.n589 585
R678 B.n591 B.n590 585
R679 B.n307 B.n306 585
R680 B.n308 B.n307 585
R681 B.n599 B.n598 585
R682 B.n598 B.n597 585
R683 B.n600 B.n305 585
R684 B.n305 B.n304 585
R685 B.n602 B.n601 585
R686 B.n603 B.n602 585
R687 B.n299 B.n298 585
R688 B.n300 B.n299 585
R689 B.n611 B.n610 585
R690 B.n610 B.n609 585
R691 B.n612 B.n297 585
R692 B.n297 B.n296 585
R693 B.n614 B.n613 585
R694 B.n615 B.n614 585
R695 B.n291 B.n290 585
R696 B.n292 B.n291 585
R697 B.n623 B.n622 585
R698 B.n622 B.n621 585
R699 B.n624 B.n289 585
R700 B.n289 B.n288 585
R701 B.n626 B.n625 585
R702 B.n627 B.n626 585
R703 B.n283 B.n282 585
R704 B.n284 B.n283 585
R705 B.n635 B.n634 585
R706 B.n634 B.n633 585
R707 B.n636 B.n281 585
R708 B.n281 B.n280 585
R709 B.n638 B.n637 585
R710 B.n639 B.n638 585
R711 B.n275 B.n274 585
R712 B.n276 B.n275 585
R713 B.n647 B.n646 585
R714 B.n646 B.n645 585
R715 B.n648 B.n273 585
R716 B.n273 B.n271 585
R717 B.n650 B.n649 585
R718 B.n651 B.n650 585
R719 B.n267 B.n266 585
R720 B.n272 B.n267 585
R721 B.n659 B.n658 585
R722 B.n658 B.n657 585
R723 B.n660 B.n265 585
R724 B.n265 B.n264 585
R725 B.n662 B.n661 585
R726 B.n663 B.n662 585
R727 B.n259 B.n258 585
R728 B.n260 B.n259 585
R729 B.n671 B.n670 585
R730 B.n670 B.n669 585
R731 B.n672 B.n257 585
R732 B.n257 B.n256 585
R733 B.n674 B.n673 585
R734 B.n675 B.n674 585
R735 B.n251 B.n250 585
R736 B.n252 B.n251 585
R737 B.n684 B.n683 585
R738 B.n683 B.n682 585
R739 B.n685 B.n249 585
R740 B.n681 B.n249 585
R741 B.n687 B.n686 585
R742 B.n688 B.n687 585
R743 B.n244 B.n243 585
R744 B.n245 B.n244 585
R745 B.n697 B.n696 585
R746 B.n696 B.n695 585
R747 B.n698 B.n242 585
R748 B.n242 B.n241 585
R749 B.n700 B.n699 585
R750 B.n701 B.n700 585
R751 B.n3 B.n0 585
R752 B.n4 B.n3 585
R753 B.n941 B.n1 585
R754 B.n942 B.n941 585
R755 B.n940 B.n939 585
R756 B.n940 B.n8 585
R757 B.n938 B.n9 585
R758 B.n12 B.n9 585
R759 B.n937 B.n936 585
R760 B.n936 B.n935 585
R761 B.n11 B.n10 585
R762 B.n934 B.n11 585
R763 B.n932 B.n931 585
R764 B.n933 B.n932 585
R765 B.n930 B.n16 585
R766 B.n19 B.n16 585
R767 B.n929 B.n928 585
R768 B.n928 B.n927 585
R769 B.n18 B.n17 585
R770 B.n926 B.n18 585
R771 B.n924 B.n923 585
R772 B.n925 B.n924 585
R773 B.n922 B.n24 585
R774 B.n24 B.n23 585
R775 B.n921 B.n920 585
R776 B.n920 B.n919 585
R777 B.n26 B.n25 585
R778 B.n918 B.n26 585
R779 B.n916 B.n915 585
R780 B.n917 B.n916 585
R781 B.n914 B.n31 585
R782 B.n31 B.n30 585
R783 B.n913 B.n912 585
R784 B.n912 B.n911 585
R785 B.n33 B.n32 585
R786 B.n910 B.n33 585
R787 B.n908 B.n907 585
R788 B.n909 B.n908 585
R789 B.n906 B.n38 585
R790 B.n38 B.n37 585
R791 B.n905 B.n904 585
R792 B.n904 B.n903 585
R793 B.n40 B.n39 585
R794 B.n902 B.n40 585
R795 B.n900 B.n899 585
R796 B.n901 B.n900 585
R797 B.n898 B.n45 585
R798 B.n45 B.n44 585
R799 B.n897 B.n896 585
R800 B.n896 B.n895 585
R801 B.n47 B.n46 585
R802 B.n894 B.n47 585
R803 B.n892 B.n891 585
R804 B.n893 B.n892 585
R805 B.n890 B.n52 585
R806 B.n52 B.n51 585
R807 B.n889 B.n888 585
R808 B.n888 B.n887 585
R809 B.n54 B.n53 585
R810 B.n886 B.n54 585
R811 B.n884 B.n883 585
R812 B.n885 B.n884 585
R813 B.n882 B.n59 585
R814 B.n59 B.n58 585
R815 B.n881 B.n880 585
R816 B.n880 B.n879 585
R817 B.n61 B.n60 585
R818 B.n878 B.n61 585
R819 B.n876 B.n875 585
R820 B.n877 B.n876 585
R821 B.n874 B.n66 585
R822 B.n66 B.n65 585
R823 B.n873 B.n872 585
R824 B.n872 B.n871 585
R825 B.n68 B.n67 585
R826 B.n870 B.n68 585
R827 B.n868 B.n867 585
R828 B.n869 B.n868 585
R829 B.n866 B.n72 585
R830 B.n75 B.n72 585
R831 B.n865 B.n864 585
R832 B.n864 B.n863 585
R833 B.n74 B.n73 585
R834 B.n862 B.n74 585
R835 B.n860 B.n859 585
R836 B.n861 B.n860 585
R837 B.n858 B.n80 585
R838 B.n80 B.n79 585
R839 B.n857 B.n856 585
R840 B.n856 B.n855 585
R841 B.n82 B.n81 585
R842 B.n854 B.n82 585
R843 B.n852 B.n851 585
R844 B.n853 B.n852 585
R845 B.n850 B.n87 585
R846 B.n87 B.n86 585
R847 B.n849 B.n848 585
R848 B.n848 B.n847 585
R849 B.n89 B.n88 585
R850 B.n846 B.n89 585
R851 B.n844 B.n843 585
R852 B.n845 B.n844 585
R853 B.n842 B.n94 585
R854 B.n94 B.n93 585
R855 B.n841 B.n840 585
R856 B.n840 B.n839 585
R857 B.n96 B.n95 585
R858 B.n838 B.n96 585
R859 B.n836 B.n835 585
R860 B.n837 B.n836 585
R861 B.n834 B.n101 585
R862 B.n101 B.n100 585
R863 B.n833 B.n832 585
R864 B.n832 B.n831 585
R865 B.n103 B.n102 585
R866 B.n830 B.n103 585
R867 B.n828 B.n827 585
R868 B.n829 B.n828 585
R869 B.n826 B.n108 585
R870 B.n108 B.n107 585
R871 B.n825 B.n824 585
R872 B.n824 B.n823 585
R873 B.n110 B.n109 585
R874 B.n822 B.n110 585
R875 B.n820 B.n819 585
R876 B.n821 B.n820 585
R877 B.n818 B.n114 585
R878 B.n117 B.n114 585
R879 B.n817 B.n816 585
R880 B.n816 B.n815 585
R881 B.n116 B.n115 585
R882 B.n814 B.n116 585
R883 B.n812 B.n811 585
R884 B.n813 B.n812 585
R885 B.n810 B.n122 585
R886 B.n122 B.n121 585
R887 B.n809 B.n808 585
R888 B.n808 B.n807 585
R889 B.n124 B.n123 585
R890 B.n806 B.n124 585
R891 B.n804 B.n803 585
R892 B.n805 B.n804 585
R893 B.n802 B.n129 585
R894 B.n129 B.n128 585
R895 B.n945 B.n944 585
R896 B.n943 B.n2 585
R897 B.n800 B.n129 492.5
R898 B.n797 B.n153 492.5
R899 B.n404 B.n373 492.5
R900 B.n488 B.n375 492.5
R901 B.n798 B.n151 256.663
R902 B.n798 B.n150 256.663
R903 B.n798 B.n149 256.663
R904 B.n798 B.n148 256.663
R905 B.n798 B.n147 256.663
R906 B.n798 B.n146 256.663
R907 B.n798 B.n145 256.663
R908 B.n798 B.n144 256.663
R909 B.n798 B.n143 256.663
R910 B.n798 B.n142 256.663
R911 B.n798 B.n141 256.663
R912 B.n798 B.n140 256.663
R913 B.n798 B.n139 256.663
R914 B.n798 B.n138 256.663
R915 B.n798 B.n137 256.663
R916 B.n798 B.n136 256.663
R917 B.n798 B.n135 256.663
R918 B.n798 B.n134 256.663
R919 B.n798 B.n133 256.663
R920 B.n798 B.n132 256.663
R921 B.n799 B.n798 256.663
R922 B.n487 B.n486 256.663
R923 B.n486 B.n378 256.663
R924 B.n486 B.n379 256.663
R925 B.n486 B.n380 256.663
R926 B.n486 B.n381 256.663
R927 B.n486 B.n382 256.663
R928 B.n486 B.n383 256.663
R929 B.n486 B.n384 256.663
R930 B.n486 B.n385 256.663
R931 B.n486 B.n386 256.663
R932 B.n486 B.n387 256.663
R933 B.n486 B.n388 256.663
R934 B.n486 B.n389 256.663
R935 B.n486 B.n390 256.663
R936 B.n486 B.n391 256.663
R937 B.n486 B.n392 256.663
R938 B.n486 B.n393 256.663
R939 B.n486 B.n394 256.663
R940 B.n486 B.n395 256.663
R941 B.n486 B.n396 256.663
R942 B.n486 B.n397 256.663
R943 B.n947 B.n946 256.663
R944 B.n157 B.t18 234.96
R945 B.n154 B.t10 234.96
R946 B.n402 B.t14 234.96
R947 B.n399 B.t21 234.96
R948 B.n159 B.n131 163.367
R949 B.n163 B.n162 163.367
R950 B.n167 B.n166 163.367
R951 B.n171 B.n170 163.367
R952 B.n175 B.n174 163.367
R953 B.n179 B.n178 163.367
R954 B.n183 B.n182 163.367
R955 B.n187 B.n186 163.367
R956 B.n192 B.n191 163.367
R957 B.n196 B.n195 163.367
R958 B.n200 B.n199 163.367
R959 B.n204 B.n203 163.367
R960 B.n208 B.n207 163.367
R961 B.n212 B.n211 163.367
R962 B.n216 B.n215 163.367
R963 B.n220 B.n219 163.367
R964 B.n224 B.n223 163.367
R965 B.n228 B.n227 163.367
R966 B.n232 B.n231 163.367
R967 B.n236 B.n235 163.367
R968 B.n797 B.n152 163.367
R969 B.n494 B.n373 163.367
R970 B.n494 B.n371 163.367
R971 B.n498 B.n371 163.367
R972 B.n498 B.n365 163.367
R973 B.n506 B.n365 163.367
R974 B.n506 B.n363 163.367
R975 B.n510 B.n363 163.367
R976 B.n510 B.n358 163.367
R977 B.n519 B.n358 163.367
R978 B.n519 B.n356 163.367
R979 B.n523 B.n356 163.367
R980 B.n523 B.n350 163.367
R981 B.n531 B.n350 163.367
R982 B.n531 B.n348 163.367
R983 B.n535 B.n348 163.367
R984 B.n535 B.n342 163.367
R985 B.n543 B.n342 163.367
R986 B.n543 B.n340 163.367
R987 B.n547 B.n340 163.367
R988 B.n547 B.n333 163.367
R989 B.n555 B.n333 163.367
R990 B.n555 B.n331 163.367
R991 B.n559 B.n331 163.367
R992 B.n559 B.n326 163.367
R993 B.n567 B.n326 163.367
R994 B.n567 B.n324 163.367
R995 B.n571 B.n324 163.367
R996 B.n571 B.n318 163.367
R997 B.n579 B.n318 163.367
R998 B.n579 B.n316 163.367
R999 B.n583 B.n316 163.367
R1000 B.n583 B.n311 163.367
R1001 B.n592 B.n311 163.367
R1002 B.n592 B.n309 163.367
R1003 B.n596 B.n309 163.367
R1004 B.n596 B.n303 163.367
R1005 B.n604 B.n303 163.367
R1006 B.n604 B.n301 163.367
R1007 B.n608 B.n301 163.367
R1008 B.n608 B.n295 163.367
R1009 B.n616 B.n295 163.367
R1010 B.n616 B.n293 163.367
R1011 B.n620 B.n293 163.367
R1012 B.n620 B.n287 163.367
R1013 B.n628 B.n287 163.367
R1014 B.n628 B.n285 163.367
R1015 B.n632 B.n285 163.367
R1016 B.n632 B.n279 163.367
R1017 B.n640 B.n279 163.367
R1018 B.n640 B.n277 163.367
R1019 B.n644 B.n277 163.367
R1020 B.n644 B.n270 163.367
R1021 B.n652 B.n270 163.367
R1022 B.n652 B.n268 163.367
R1023 B.n656 B.n268 163.367
R1024 B.n656 B.n263 163.367
R1025 B.n664 B.n263 163.367
R1026 B.n664 B.n261 163.367
R1027 B.n668 B.n261 163.367
R1028 B.n668 B.n255 163.367
R1029 B.n676 B.n255 163.367
R1030 B.n676 B.n253 163.367
R1031 B.n680 B.n253 163.367
R1032 B.n680 B.n248 163.367
R1033 B.n689 B.n248 163.367
R1034 B.n689 B.n246 163.367
R1035 B.n694 B.n246 163.367
R1036 B.n694 B.n240 163.367
R1037 B.n702 B.n240 163.367
R1038 B.n703 B.n702 163.367
R1039 B.n703 B.n5 163.367
R1040 B.n6 B.n5 163.367
R1041 B.n7 B.n6 163.367
R1042 B.n709 B.n7 163.367
R1043 B.n710 B.n709 163.367
R1044 B.n710 B.n13 163.367
R1045 B.n14 B.n13 163.367
R1046 B.n15 B.n14 163.367
R1047 B.n715 B.n15 163.367
R1048 B.n715 B.n20 163.367
R1049 B.n21 B.n20 163.367
R1050 B.n22 B.n21 163.367
R1051 B.n720 B.n22 163.367
R1052 B.n720 B.n27 163.367
R1053 B.n28 B.n27 163.367
R1054 B.n29 B.n28 163.367
R1055 B.n725 B.n29 163.367
R1056 B.n725 B.n34 163.367
R1057 B.n35 B.n34 163.367
R1058 B.n36 B.n35 163.367
R1059 B.n730 B.n36 163.367
R1060 B.n730 B.n41 163.367
R1061 B.n42 B.n41 163.367
R1062 B.n43 B.n42 163.367
R1063 B.n735 B.n43 163.367
R1064 B.n735 B.n48 163.367
R1065 B.n49 B.n48 163.367
R1066 B.n50 B.n49 163.367
R1067 B.n740 B.n50 163.367
R1068 B.n740 B.n55 163.367
R1069 B.n56 B.n55 163.367
R1070 B.n57 B.n56 163.367
R1071 B.n745 B.n57 163.367
R1072 B.n745 B.n62 163.367
R1073 B.n63 B.n62 163.367
R1074 B.n64 B.n63 163.367
R1075 B.n750 B.n64 163.367
R1076 B.n750 B.n69 163.367
R1077 B.n70 B.n69 163.367
R1078 B.n71 B.n70 163.367
R1079 B.n755 B.n71 163.367
R1080 B.n755 B.n76 163.367
R1081 B.n77 B.n76 163.367
R1082 B.n78 B.n77 163.367
R1083 B.n760 B.n78 163.367
R1084 B.n760 B.n83 163.367
R1085 B.n84 B.n83 163.367
R1086 B.n85 B.n84 163.367
R1087 B.n765 B.n85 163.367
R1088 B.n765 B.n90 163.367
R1089 B.n91 B.n90 163.367
R1090 B.n92 B.n91 163.367
R1091 B.n770 B.n92 163.367
R1092 B.n770 B.n97 163.367
R1093 B.n98 B.n97 163.367
R1094 B.n99 B.n98 163.367
R1095 B.n775 B.n99 163.367
R1096 B.n775 B.n104 163.367
R1097 B.n105 B.n104 163.367
R1098 B.n106 B.n105 163.367
R1099 B.n780 B.n106 163.367
R1100 B.n780 B.n111 163.367
R1101 B.n112 B.n111 163.367
R1102 B.n113 B.n112 163.367
R1103 B.n785 B.n113 163.367
R1104 B.n785 B.n118 163.367
R1105 B.n119 B.n118 163.367
R1106 B.n120 B.n119 163.367
R1107 B.n790 B.n120 163.367
R1108 B.n790 B.n125 163.367
R1109 B.n126 B.n125 163.367
R1110 B.n127 B.n126 163.367
R1111 B.n153 B.n127 163.367
R1112 B.n485 B.n377 163.367
R1113 B.n485 B.n398 163.367
R1114 B.n481 B.n480 163.367
R1115 B.n477 B.n476 163.367
R1116 B.n473 B.n472 163.367
R1117 B.n469 B.n468 163.367
R1118 B.n465 B.n464 163.367
R1119 B.n461 B.n460 163.367
R1120 B.n457 B.n456 163.367
R1121 B.n453 B.n452 163.367
R1122 B.n449 B.n448 163.367
R1123 B.n445 B.n444 163.367
R1124 B.n441 B.n440 163.367
R1125 B.n436 B.n435 163.367
R1126 B.n432 B.n431 163.367
R1127 B.n428 B.n427 163.367
R1128 B.n424 B.n423 163.367
R1129 B.n420 B.n419 163.367
R1130 B.n416 B.n415 163.367
R1131 B.n412 B.n411 163.367
R1132 B.n408 B.n407 163.367
R1133 B.n492 B.n375 163.367
R1134 B.n492 B.n369 163.367
R1135 B.n500 B.n369 163.367
R1136 B.n500 B.n367 163.367
R1137 B.n504 B.n367 163.367
R1138 B.n504 B.n361 163.367
R1139 B.n513 B.n361 163.367
R1140 B.n513 B.n359 163.367
R1141 B.n517 B.n359 163.367
R1142 B.n517 B.n354 163.367
R1143 B.n525 B.n354 163.367
R1144 B.n525 B.n352 163.367
R1145 B.n529 B.n352 163.367
R1146 B.n529 B.n346 163.367
R1147 B.n537 B.n346 163.367
R1148 B.n537 B.n344 163.367
R1149 B.n541 B.n344 163.367
R1150 B.n541 B.n338 163.367
R1151 B.n549 B.n338 163.367
R1152 B.n549 B.n336 163.367
R1153 B.n553 B.n336 163.367
R1154 B.n553 B.n330 163.367
R1155 B.n561 B.n330 163.367
R1156 B.n561 B.n328 163.367
R1157 B.n565 B.n328 163.367
R1158 B.n565 B.n322 163.367
R1159 B.n573 B.n322 163.367
R1160 B.n573 B.n320 163.367
R1161 B.n577 B.n320 163.367
R1162 B.n577 B.n314 163.367
R1163 B.n586 B.n314 163.367
R1164 B.n586 B.n312 163.367
R1165 B.n590 B.n312 163.367
R1166 B.n590 B.n307 163.367
R1167 B.n598 B.n307 163.367
R1168 B.n598 B.n305 163.367
R1169 B.n602 B.n305 163.367
R1170 B.n602 B.n299 163.367
R1171 B.n610 B.n299 163.367
R1172 B.n610 B.n297 163.367
R1173 B.n614 B.n297 163.367
R1174 B.n614 B.n291 163.367
R1175 B.n622 B.n291 163.367
R1176 B.n622 B.n289 163.367
R1177 B.n626 B.n289 163.367
R1178 B.n626 B.n283 163.367
R1179 B.n634 B.n283 163.367
R1180 B.n634 B.n281 163.367
R1181 B.n638 B.n281 163.367
R1182 B.n638 B.n275 163.367
R1183 B.n646 B.n275 163.367
R1184 B.n646 B.n273 163.367
R1185 B.n650 B.n273 163.367
R1186 B.n650 B.n267 163.367
R1187 B.n658 B.n267 163.367
R1188 B.n658 B.n265 163.367
R1189 B.n662 B.n265 163.367
R1190 B.n662 B.n259 163.367
R1191 B.n670 B.n259 163.367
R1192 B.n670 B.n257 163.367
R1193 B.n674 B.n257 163.367
R1194 B.n674 B.n251 163.367
R1195 B.n683 B.n251 163.367
R1196 B.n683 B.n249 163.367
R1197 B.n687 B.n249 163.367
R1198 B.n687 B.n244 163.367
R1199 B.n696 B.n244 163.367
R1200 B.n696 B.n242 163.367
R1201 B.n700 B.n242 163.367
R1202 B.n700 B.n3 163.367
R1203 B.n945 B.n3 163.367
R1204 B.n941 B.n2 163.367
R1205 B.n941 B.n940 163.367
R1206 B.n940 B.n9 163.367
R1207 B.n936 B.n9 163.367
R1208 B.n936 B.n11 163.367
R1209 B.n932 B.n11 163.367
R1210 B.n932 B.n16 163.367
R1211 B.n928 B.n16 163.367
R1212 B.n928 B.n18 163.367
R1213 B.n924 B.n18 163.367
R1214 B.n924 B.n24 163.367
R1215 B.n920 B.n24 163.367
R1216 B.n920 B.n26 163.367
R1217 B.n916 B.n26 163.367
R1218 B.n916 B.n31 163.367
R1219 B.n912 B.n31 163.367
R1220 B.n912 B.n33 163.367
R1221 B.n908 B.n33 163.367
R1222 B.n908 B.n38 163.367
R1223 B.n904 B.n38 163.367
R1224 B.n904 B.n40 163.367
R1225 B.n900 B.n40 163.367
R1226 B.n900 B.n45 163.367
R1227 B.n896 B.n45 163.367
R1228 B.n896 B.n47 163.367
R1229 B.n892 B.n47 163.367
R1230 B.n892 B.n52 163.367
R1231 B.n888 B.n52 163.367
R1232 B.n888 B.n54 163.367
R1233 B.n884 B.n54 163.367
R1234 B.n884 B.n59 163.367
R1235 B.n880 B.n59 163.367
R1236 B.n880 B.n61 163.367
R1237 B.n876 B.n61 163.367
R1238 B.n876 B.n66 163.367
R1239 B.n872 B.n66 163.367
R1240 B.n872 B.n68 163.367
R1241 B.n868 B.n68 163.367
R1242 B.n868 B.n72 163.367
R1243 B.n864 B.n72 163.367
R1244 B.n864 B.n74 163.367
R1245 B.n860 B.n74 163.367
R1246 B.n860 B.n80 163.367
R1247 B.n856 B.n80 163.367
R1248 B.n856 B.n82 163.367
R1249 B.n852 B.n82 163.367
R1250 B.n852 B.n87 163.367
R1251 B.n848 B.n87 163.367
R1252 B.n848 B.n89 163.367
R1253 B.n844 B.n89 163.367
R1254 B.n844 B.n94 163.367
R1255 B.n840 B.n94 163.367
R1256 B.n840 B.n96 163.367
R1257 B.n836 B.n96 163.367
R1258 B.n836 B.n101 163.367
R1259 B.n832 B.n101 163.367
R1260 B.n832 B.n103 163.367
R1261 B.n828 B.n103 163.367
R1262 B.n828 B.n108 163.367
R1263 B.n824 B.n108 163.367
R1264 B.n824 B.n110 163.367
R1265 B.n820 B.n110 163.367
R1266 B.n820 B.n114 163.367
R1267 B.n816 B.n114 163.367
R1268 B.n816 B.n116 163.367
R1269 B.n812 B.n116 163.367
R1270 B.n812 B.n122 163.367
R1271 B.n808 B.n122 163.367
R1272 B.n808 B.n124 163.367
R1273 B.n804 B.n124 163.367
R1274 B.n804 B.n129 163.367
R1275 B.n486 B.n374 151.165
R1276 B.n798 B.n128 151.165
R1277 B.n154 B.t12 144.716
R1278 B.n402 B.t17 144.716
R1279 B.n157 B.t19 144.714
R1280 B.n399 B.t23 144.714
R1281 B.n493 B.n374 84.9522
R1282 B.n493 B.n370 84.9522
R1283 B.n499 B.n370 84.9522
R1284 B.n499 B.n366 84.9522
R1285 B.n505 B.n366 84.9522
R1286 B.n505 B.n362 84.9522
R1287 B.n512 B.n362 84.9522
R1288 B.n512 B.n511 84.9522
R1289 B.n518 B.n355 84.9522
R1290 B.n524 B.n355 84.9522
R1291 B.n524 B.n351 84.9522
R1292 B.n530 B.n351 84.9522
R1293 B.n530 B.n347 84.9522
R1294 B.n536 B.n347 84.9522
R1295 B.n536 B.n343 84.9522
R1296 B.n542 B.n343 84.9522
R1297 B.n542 B.n339 84.9522
R1298 B.n548 B.n339 84.9522
R1299 B.n548 B.n334 84.9522
R1300 B.n554 B.n334 84.9522
R1301 B.n554 B.n335 84.9522
R1302 B.n560 B.n327 84.9522
R1303 B.n566 B.n327 84.9522
R1304 B.n566 B.n323 84.9522
R1305 B.n572 B.n323 84.9522
R1306 B.n572 B.n319 84.9522
R1307 B.n578 B.n319 84.9522
R1308 B.n578 B.n315 84.9522
R1309 B.n585 B.n315 84.9522
R1310 B.n585 B.n584 84.9522
R1311 B.n591 B.n308 84.9522
R1312 B.n597 B.n308 84.9522
R1313 B.n597 B.n304 84.9522
R1314 B.n603 B.n304 84.9522
R1315 B.n603 B.n300 84.9522
R1316 B.n609 B.n300 84.9522
R1317 B.n609 B.n296 84.9522
R1318 B.n615 B.n296 84.9522
R1319 B.n615 B.n292 84.9522
R1320 B.n621 B.n292 84.9522
R1321 B.n627 B.n288 84.9522
R1322 B.n627 B.n284 84.9522
R1323 B.n633 B.n284 84.9522
R1324 B.n633 B.n280 84.9522
R1325 B.n639 B.n280 84.9522
R1326 B.n639 B.n276 84.9522
R1327 B.n645 B.n276 84.9522
R1328 B.n645 B.n271 84.9522
R1329 B.n651 B.n271 84.9522
R1330 B.n651 B.n272 84.9522
R1331 B.n657 B.n264 84.9522
R1332 B.n663 B.n264 84.9522
R1333 B.n663 B.n260 84.9522
R1334 B.n669 B.n260 84.9522
R1335 B.n669 B.n256 84.9522
R1336 B.n675 B.n256 84.9522
R1337 B.n675 B.n252 84.9522
R1338 B.n682 B.n252 84.9522
R1339 B.n682 B.n681 84.9522
R1340 B.n688 B.n245 84.9522
R1341 B.n695 B.n245 84.9522
R1342 B.n695 B.n241 84.9522
R1343 B.n701 B.n241 84.9522
R1344 B.n701 B.n4 84.9522
R1345 B.n944 B.n4 84.9522
R1346 B.n944 B.n943 84.9522
R1347 B.n943 B.n942 84.9522
R1348 B.n942 B.n8 84.9522
R1349 B.n12 B.n8 84.9522
R1350 B.n935 B.n12 84.9522
R1351 B.n935 B.n934 84.9522
R1352 B.n934 B.n933 84.9522
R1353 B.n927 B.n19 84.9522
R1354 B.n927 B.n926 84.9522
R1355 B.n926 B.n925 84.9522
R1356 B.n925 B.n23 84.9522
R1357 B.n919 B.n23 84.9522
R1358 B.n919 B.n918 84.9522
R1359 B.n918 B.n917 84.9522
R1360 B.n917 B.n30 84.9522
R1361 B.n911 B.n30 84.9522
R1362 B.n910 B.n909 84.9522
R1363 B.n909 B.n37 84.9522
R1364 B.n903 B.n37 84.9522
R1365 B.n903 B.n902 84.9522
R1366 B.n902 B.n901 84.9522
R1367 B.n901 B.n44 84.9522
R1368 B.n895 B.n44 84.9522
R1369 B.n895 B.n894 84.9522
R1370 B.n894 B.n893 84.9522
R1371 B.n893 B.n51 84.9522
R1372 B.n887 B.n886 84.9522
R1373 B.n886 B.n885 84.9522
R1374 B.n885 B.n58 84.9522
R1375 B.n879 B.n58 84.9522
R1376 B.n879 B.n878 84.9522
R1377 B.n878 B.n877 84.9522
R1378 B.n877 B.n65 84.9522
R1379 B.n871 B.n65 84.9522
R1380 B.n871 B.n870 84.9522
R1381 B.n870 B.n869 84.9522
R1382 B.n863 B.n75 84.9522
R1383 B.n863 B.n862 84.9522
R1384 B.n862 B.n861 84.9522
R1385 B.n861 B.n79 84.9522
R1386 B.n855 B.n79 84.9522
R1387 B.n855 B.n854 84.9522
R1388 B.n854 B.n853 84.9522
R1389 B.n853 B.n86 84.9522
R1390 B.n847 B.n86 84.9522
R1391 B.n846 B.n845 84.9522
R1392 B.n845 B.n93 84.9522
R1393 B.n839 B.n93 84.9522
R1394 B.n839 B.n838 84.9522
R1395 B.n838 B.n837 84.9522
R1396 B.n837 B.n100 84.9522
R1397 B.n831 B.n100 84.9522
R1398 B.n831 B.n830 84.9522
R1399 B.n830 B.n829 84.9522
R1400 B.n829 B.n107 84.9522
R1401 B.n823 B.n107 84.9522
R1402 B.n823 B.n822 84.9522
R1403 B.n822 B.n821 84.9522
R1404 B.n815 B.n117 84.9522
R1405 B.n815 B.n814 84.9522
R1406 B.n814 B.n813 84.9522
R1407 B.n813 B.n121 84.9522
R1408 B.n807 B.n121 84.9522
R1409 B.n807 B.n806 84.9522
R1410 B.n806 B.n805 84.9522
R1411 B.n805 B.n128 84.9522
R1412 B.n584 B.t7 79.9551
R1413 B.n657 B.t2 79.9551
R1414 B.n911 B.t4 79.9551
R1415 B.n75 B.t6 79.9551
R1416 B.n155 B.t13 75.0918
R1417 B.n403 B.t16 75.0918
R1418 B.n158 B.t20 75.0889
R1419 B.n400 B.t22 75.0889
R1420 B.n800 B.n799 71.676
R1421 B.n159 B.n132 71.676
R1422 B.n163 B.n133 71.676
R1423 B.n167 B.n134 71.676
R1424 B.n171 B.n135 71.676
R1425 B.n175 B.n136 71.676
R1426 B.n179 B.n137 71.676
R1427 B.n183 B.n138 71.676
R1428 B.n187 B.n139 71.676
R1429 B.n192 B.n140 71.676
R1430 B.n196 B.n141 71.676
R1431 B.n200 B.n142 71.676
R1432 B.n204 B.n143 71.676
R1433 B.n208 B.n144 71.676
R1434 B.n212 B.n145 71.676
R1435 B.n216 B.n146 71.676
R1436 B.n220 B.n147 71.676
R1437 B.n224 B.n148 71.676
R1438 B.n228 B.n149 71.676
R1439 B.n232 B.n150 71.676
R1440 B.n236 B.n151 71.676
R1441 B.n152 B.n151 71.676
R1442 B.n235 B.n150 71.676
R1443 B.n231 B.n149 71.676
R1444 B.n227 B.n148 71.676
R1445 B.n223 B.n147 71.676
R1446 B.n219 B.n146 71.676
R1447 B.n215 B.n145 71.676
R1448 B.n211 B.n144 71.676
R1449 B.n207 B.n143 71.676
R1450 B.n203 B.n142 71.676
R1451 B.n199 B.n141 71.676
R1452 B.n195 B.n140 71.676
R1453 B.n191 B.n139 71.676
R1454 B.n186 B.n138 71.676
R1455 B.n182 B.n137 71.676
R1456 B.n178 B.n136 71.676
R1457 B.n174 B.n135 71.676
R1458 B.n170 B.n134 71.676
R1459 B.n166 B.n133 71.676
R1460 B.n162 B.n132 71.676
R1461 B.n799 B.n131 71.676
R1462 B.n488 B.n487 71.676
R1463 B.n398 B.n378 71.676
R1464 B.n480 B.n379 71.676
R1465 B.n476 B.n380 71.676
R1466 B.n472 B.n381 71.676
R1467 B.n468 B.n382 71.676
R1468 B.n464 B.n383 71.676
R1469 B.n460 B.n384 71.676
R1470 B.n456 B.n385 71.676
R1471 B.n452 B.n386 71.676
R1472 B.n448 B.n387 71.676
R1473 B.n444 B.n388 71.676
R1474 B.n440 B.n389 71.676
R1475 B.n435 B.n390 71.676
R1476 B.n431 B.n391 71.676
R1477 B.n427 B.n392 71.676
R1478 B.n423 B.n393 71.676
R1479 B.n419 B.n394 71.676
R1480 B.n415 B.n395 71.676
R1481 B.n411 B.n396 71.676
R1482 B.n407 B.n397 71.676
R1483 B.n487 B.n377 71.676
R1484 B.n481 B.n378 71.676
R1485 B.n477 B.n379 71.676
R1486 B.n473 B.n380 71.676
R1487 B.n469 B.n381 71.676
R1488 B.n465 B.n382 71.676
R1489 B.n461 B.n383 71.676
R1490 B.n457 B.n384 71.676
R1491 B.n453 B.n385 71.676
R1492 B.n449 B.n386 71.676
R1493 B.n445 B.n387 71.676
R1494 B.n441 B.n388 71.676
R1495 B.n436 B.n389 71.676
R1496 B.n432 B.n390 71.676
R1497 B.n428 B.n391 71.676
R1498 B.n424 B.n392 71.676
R1499 B.n420 B.n393 71.676
R1500 B.n416 B.n394 71.676
R1501 B.n412 B.n395 71.676
R1502 B.n408 B.n396 71.676
R1503 B.n404 B.n397 71.676
R1504 B.n946 B.n945 71.676
R1505 B.n946 B.n2 71.676
R1506 B.n158 B.n157 69.6247
R1507 B.n155 B.n154 69.6247
R1508 B.n403 B.n402 69.6247
R1509 B.n400 B.n399 69.6247
R1510 B.n189 B.n158 59.5399
R1511 B.n156 B.n155 59.5399
R1512 B.n438 B.n403 59.5399
R1513 B.n401 B.n400 59.5399
R1514 B.n511 B.t15 52.4707
R1515 B.n560 B.t0 52.4707
R1516 B.n681 B.t8 52.4707
R1517 B.n19 B.t3 52.4707
R1518 B.n847 B.t9 52.4707
R1519 B.n117 B.t11 52.4707
R1520 B.n621 B.t1 42.4764
R1521 B.t1 B.n288 42.4764
R1522 B.t5 B.n51 42.4764
R1523 B.n887 B.t5 42.4764
R1524 B.n518 B.t15 32.482
R1525 B.n335 B.t0 32.482
R1526 B.n688 B.t8 32.482
R1527 B.n933 B.t3 32.482
R1528 B.t9 B.n846 32.482
R1529 B.n821 B.t11 32.482
R1530 B.n490 B.n489 32.0005
R1531 B.n405 B.n372 32.0005
R1532 B.n796 B.n795 32.0005
R1533 B.n802 B.n801 32.0005
R1534 B B.n947 18.0485
R1535 B.n491 B.n490 10.6151
R1536 B.n491 B.n368 10.6151
R1537 B.n501 B.n368 10.6151
R1538 B.n502 B.n501 10.6151
R1539 B.n503 B.n502 10.6151
R1540 B.n503 B.n360 10.6151
R1541 B.n514 B.n360 10.6151
R1542 B.n515 B.n514 10.6151
R1543 B.n516 B.n515 10.6151
R1544 B.n516 B.n353 10.6151
R1545 B.n526 B.n353 10.6151
R1546 B.n527 B.n526 10.6151
R1547 B.n528 B.n527 10.6151
R1548 B.n528 B.n345 10.6151
R1549 B.n538 B.n345 10.6151
R1550 B.n539 B.n538 10.6151
R1551 B.n540 B.n539 10.6151
R1552 B.n540 B.n337 10.6151
R1553 B.n550 B.n337 10.6151
R1554 B.n551 B.n550 10.6151
R1555 B.n552 B.n551 10.6151
R1556 B.n552 B.n329 10.6151
R1557 B.n562 B.n329 10.6151
R1558 B.n563 B.n562 10.6151
R1559 B.n564 B.n563 10.6151
R1560 B.n564 B.n321 10.6151
R1561 B.n574 B.n321 10.6151
R1562 B.n575 B.n574 10.6151
R1563 B.n576 B.n575 10.6151
R1564 B.n576 B.n313 10.6151
R1565 B.n587 B.n313 10.6151
R1566 B.n588 B.n587 10.6151
R1567 B.n589 B.n588 10.6151
R1568 B.n589 B.n306 10.6151
R1569 B.n599 B.n306 10.6151
R1570 B.n600 B.n599 10.6151
R1571 B.n601 B.n600 10.6151
R1572 B.n601 B.n298 10.6151
R1573 B.n611 B.n298 10.6151
R1574 B.n612 B.n611 10.6151
R1575 B.n613 B.n612 10.6151
R1576 B.n613 B.n290 10.6151
R1577 B.n623 B.n290 10.6151
R1578 B.n624 B.n623 10.6151
R1579 B.n625 B.n624 10.6151
R1580 B.n625 B.n282 10.6151
R1581 B.n635 B.n282 10.6151
R1582 B.n636 B.n635 10.6151
R1583 B.n637 B.n636 10.6151
R1584 B.n637 B.n274 10.6151
R1585 B.n647 B.n274 10.6151
R1586 B.n648 B.n647 10.6151
R1587 B.n649 B.n648 10.6151
R1588 B.n649 B.n266 10.6151
R1589 B.n659 B.n266 10.6151
R1590 B.n660 B.n659 10.6151
R1591 B.n661 B.n660 10.6151
R1592 B.n661 B.n258 10.6151
R1593 B.n671 B.n258 10.6151
R1594 B.n672 B.n671 10.6151
R1595 B.n673 B.n672 10.6151
R1596 B.n673 B.n250 10.6151
R1597 B.n684 B.n250 10.6151
R1598 B.n685 B.n684 10.6151
R1599 B.n686 B.n685 10.6151
R1600 B.n686 B.n243 10.6151
R1601 B.n697 B.n243 10.6151
R1602 B.n698 B.n697 10.6151
R1603 B.n699 B.n698 10.6151
R1604 B.n699 B.n0 10.6151
R1605 B.n489 B.n376 10.6151
R1606 B.n484 B.n376 10.6151
R1607 B.n484 B.n483 10.6151
R1608 B.n483 B.n482 10.6151
R1609 B.n482 B.n479 10.6151
R1610 B.n479 B.n478 10.6151
R1611 B.n478 B.n475 10.6151
R1612 B.n475 B.n474 10.6151
R1613 B.n474 B.n471 10.6151
R1614 B.n471 B.n470 10.6151
R1615 B.n470 B.n467 10.6151
R1616 B.n467 B.n466 10.6151
R1617 B.n466 B.n463 10.6151
R1618 B.n463 B.n462 10.6151
R1619 B.n462 B.n459 10.6151
R1620 B.n459 B.n458 10.6151
R1621 B.n455 B.n454 10.6151
R1622 B.n454 B.n451 10.6151
R1623 B.n451 B.n450 10.6151
R1624 B.n450 B.n447 10.6151
R1625 B.n447 B.n446 10.6151
R1626 B.n446 B.n443 10.6151
R1627 B.n443 B.n442 10.6151
R1628 B.n442 B.n439 10.6151
R1629 B.n437 B.n434 10.6151
R1630 B.n434 B.n433 10.6151
R1631 B.n433 B.n430 10.6151
R1632 B.n430 B.n429 10.6151
R1633 B.n429 B.n426 10.6151
R1634 B.n426 B.n425 10.6151
R1635 B.n425 B.n422 10.6151
R1636 B.n422 B.n421 10.6151
R1637 B.n421 B.n418 10.6151
R1638 B.n418 B.n417 10.6151
R1639 B.n417 B.n414 10.6151
R1640 B.n414 B.n413 10.6151
R1641 B.n413 B.n410 10.6151
R1642 B.n410 B.n409 10.6151
R1643 B.n409 B.n406 10.6151
R1644 B.n406 B.n405 10.6151
R1645 B.n495 B.n372 10.6151
R1646 B.n496 B.n495 10.6151
R1647 B.n497 B.n496 10.6151
R1648 B.n497 B.n364 10.6151
R1649 B.n507 B.n364 10.6151
R1650 B.n508 B.n507 10.6151
R1651 B.n509 B.n508 10.6151
R1652 B.n509 B.n357 10.6151
R1653 B.n520 B.n357 10.6151
R1654 B.n521 B.n520 10.6151
R1655 B.n522 B.n521 10.6151
R1656 B.n522 B.n349 10.6151
R1657 B.n532 B.n349 10.6151
R1658 B.n533 B.n532 10.6151
R1659 B.n534 B.n533 10.6151
R1660 B.n534 B.n341 10.6151
R1661 B.n544 B.n341 10.6151
R1662 B.n545 B.n544 10.6151
R1663 B.n546 B.n545 10.6151
R1664 B.n546 B.n332 10.6151
R1665 B.n556 B.n332 10.6151
R1666 B.n557 B.n556 10.6151
R1667 B.n558 B.n557 10.6151
R1668 B.n558 B.n325 10.6151
R1669 B.n568 B.n325 10.6151
R1670 B.n569 B.n568 10.6151
R1671 B.n570 B.n569 10.6151
R1672 B.n570 B.n317 10.6151
R1673 B.n580 B.n317 10.6151
R1674 B.n581 B.n580 10.6151
R1675 B.n582 B.n581 10.6151
R1676 B.n582 B.n310 10.6151
R1677 B.n593 B.n310 10.6151
R1678 B.n594 B.n593 10.6151
R1679 B.n595 B.n594 10.6151
R1680 B.n595 B.n302 10.6151
R1681 B.n605 B.n302 10.6151
R1682 B.n606 B.n605 10.6151
R1683 B.n607 B.n606 10.6151
R1684 B.n607 B.n294 10.6151
R1685 B.n617 B.n294 10.6151
R1686 B.n618 B.n617 10.6151
R1687 B.n619 B.n618 10.6151
R1688 B.n619 B.n286 10.6151
R1689 B.n629 B.n286 10.6151
R1690 B.n630 B.n629 10.6151
R1691 B.n631 B.n630 10.6151
R1692 B.n631 B.n278 10.6151
R1693 B.n641 B.n278 10.6151
R1694 B.n642 B.n641 10.6151
R1695 B.n643 B.n642 10.6151
R1696 B.n643 B.n269 10.6151
R1697 B.n653 B.n269 10.6151
R1698 B.n654 B.n653 10.6151
R1699 B.n655 B.n654 10.6151
R1700 B.n655 B.n262 10.6151
R1701 B.n665 B.n262 10.6151
R1702 B.n666 B.n665 10.6151
R1703 B.n667 B.n666 10.6151
R1704 B.n667 B.n254 10.6151
R1705 B.n677 B.n254 10.6151
R1706 B.n678 B.n677 10.6151
R1707 B.n679 B.n678 10.6151
R1708 B.n679 B.n247 10.6151
R1709 B.n690 B.n247 10.6151
R1710 B.n691 B.n690 10.6151
R1711 B.n693 B.n691 10.6151
R1712 B.n693 B.n692 10.6151
R1713 B.n692 B.n239 10.6151
R1714 B.n704 B.n239 10.6151
R1715 B.n705 B.n704 10.6151
R1716 B.n706 B.n705 10.6151
R1717 B.n707 B.n706 10.6151
R1718 B.n708 B.n707 10.6151
R1719 B.n711 B.n708 10.6151
R1720 B.n712 B.n711 10.6151
R1721 B.n713 B.n712 10.6151
R1722 B.n714 B.n713 10.6151
R1723 B.n716 B.n714 10.6151
R1724 B.n717 B.n716 10.6151
R1725 B.n718 B.n717 10.6151
R1726 B.n719 B.n718 10.6151
R1727 B.n721 B.n719 10.6151
R1728 B.n722 B.n721 10.6151
R1729 B.n723 B.n722 10.6151
R1730 B.n724 B.n723 10.6151
R1731 B.n726 B.n724 10.6151
R1732 B.n727 B.n726 10.6151
R1733 B.n728 B.n727 10.6151
R1734 B.n729 B.n728 10.6151
R1735 B.n731 B.n729 10.6151
R1736 B.n732 B.n731 10.6151
R1737 B.n733 B.n732 10.6151
R1738 B.n734 B.n733 10.6151
R1739 B.n736 B.n734 10.6151
R1740 B.n737 B.n736 10.6151
R1741 B.n738 B.n737 10.6151
R1742 B.n739 B.n738 10.6151
R1743 B.n741 B.n739 10.6151
R1744 B.n742 B.n741 10.6151
R1745 B.n743 B.n742 10.6151
R1746 B.n744 B.n743 10.6151
R1747 B.n746 B.n744 10.6151
R1748 B.n747 B.n746 10.6151
R1749 B.n748 B.n747 10.6151
R1750 B.n749 B.n748 10.6151
R1751 B.n751 B.n749 10.6151
R1752 B.n752 B.n751 10.6151
R1753 B.n753 B.n752 10.6151
R1754 B.n754 B.n753 10.6151
R1755 B.n756 B.n754 10.6151
R1756 B.n757 B.n756 10.6151
R1757 B.n758 B.n757 10.6151
R1758 B.n759 B.n758 10.6151
R1759 B.n761 B.n759 10.6151
R1760 B.n762 B.n761 10.6151
R1761 B.n763 B.n762 10.6151
R1762 B.n764 B.n763 10.6151
R1763 B.n766 B.n764 10.6151
R1764 B.n767 B.n766 10.6151
R1765 B.n768 B.n767 10.6151
R1766 B.n769 B.n768 10.6151
R1767 B.n771 B.n769 10.6151
R1768 B.n772 B.n771 10.6151
R1769 B.n773 B.n772 10.6151
R1770 B.n774 B.n773 10.6151
R1771 B.n776 B.n774 10.6151
R1772 B.n777 B.n776 10.6151
R1773 B.n778 B.n777 10.6151
R1774 B.n779 B.n778 10.6151
R1775 B.n781 B.n779 10.6151
R1776 B.n782 B.n781 10.6151
R1777 B.n783 B.n782 10.6151
R1778 B.n784 B.n783 10.6151
R1779 B.n786 B.n784 10.6151
R1780 B.n787 B.n786 10.6151
R1781 B.n788 B.n787 10.6151
R1782 B.n789 B.n788 10.6151
R1783 B.n791 B.n789 10.6151
R1784 B.n792 B.n791 10.6151
R1785 B.n793 B.n792 10.6151
R1786 B.n794 B.n793 10.6151
R1787 B.n795 B.n794 10.6151
R1788 B.n939 B.n1 10.6151
R1789 B.n939 B.n938 10.6151
R1790 B.n938 B.n937 10.6151
R1791 B.n937 B.n10 10.6151
R1792 B.n931 B.n10 10.6151
R1793 B.n931 B.n930 10.6151
R1794 B.n930 B.n929 10.6151
R1795 B.n929 B.n17 10.6151
R1796 B.n923 B.n17 10.6151
R1797 B.n923 B.n922 10.6151
R1798 B.n922 B.n921 10.6151
R1799 B.n921 B.n25 10.6151
R1800 B.n915 B.n25 10.6151
R1801 B.n915 B.n914 10.6151
R1802 B.n914 B.n913 10.6151
R1803 B.n913 B.n32 10.6151
R1804 B.n907 B.n32 10.6151
R1805 B.n907 B.n906 10.6151
R1806 B.n906 B.n905 10.6151
R1807 B.n905 B.n39 10.6151
R1808 B.n899 B.n39 10.6151
R1809 B.n899 B.n898 10.6151
R1810 B.n898 B.n897 10.6151
R1811 B.n897 B.n46 10.6151
R1812 B.n891 B.n46 10.6151
R1813 B.n891 B.n890 10.6151
R1814 B.n890 B.n889 10.6151
R1815 B.n889 B.n53 10.6151
R1816 B.n883 B.n53 10.6151
R1817 B.n883 B.n882 10.6151
R1818 B.n882 B.n881 10.6151
R1819 B.n881 B.n60 10.6151
R1820 B.n875 B.n60 10.6151
R1821 B.n875 B.n874 10.6151
R1822 B.n874 B.n873 10.6151
R1823 B.n873 B.n67 10.6151
R1824 B.n867 B.n67 10.6151
R1825 B.n867 B.n866 10.6151
R1826 B.n866 B.n865 10.6151
R1827 B.n865 B.n73 10.6151
R1828 B.n859 B.n73 10.6151
R1829 B.n859 B.n858 10.6151
R1830 B.n858 B.n857 10.6151
R1831 B.n857 B.n81 10.6151
R1832 B.n851 B.n81 10.6151
R1833 B.n851 B.n850 10.6151
R1834 B.n850 B.n849 10.6151
R1835 B.n849 B.n88 10.6151
R1836 B.n843 B.n88 10.6151
R1837 B.n843 B.n842 10.6151
R1838 B.n842 B.n841 10.6151
R1839 B.n841 B.n95 10.6151
R1840 B.n835 B.n95 10.6151
R1841 B.n835 B.n834 10.6151
R1842 B.n834 B.n833 10.6151
R1843 B.n833 B.n102 10.6151
R1844 B.n827 B.n102 10.6151
R1845 B.n827 B.n826 10.6151
R1846 B.n826 B.n825 10.6151
R1847 B.n825 B.n109 10.6151
R1848 B.n819 B.n109 10.6151
R1849 B.n819 B.n818 10.6151
R1850 B.n818 B.n817 10.6151
R1851 B.n817 B.n115 10.6151
R1852 B.n811 B.n115 10.6151
R1853 B.n811 B.n810 10.6151
R1854 B.n810 B.n809 10.6151
R1855 B.n809 B.n123 10.6151
R1856 B.n803 B.n123 10.6151
R1857 B.n803 B.n802 10.6151
R1858 B.n801 B.n130 10.6151
R1859 B.n160 B.n130 10.6151
R1860 B.n161 B.n160 10.6151
R1861 B.n164 B.n161 10.6151
R1862 B.n165 B.n164 10.6151
R1863 B.n168 B.n165 10.6151
R1864 B.n169 B.n168 10.6151
R1865 B.n172 B.n169 10.6151
R1866 B.n173 B.n172 10.6151
R1867 B.n176 B.n173 10.6151
R1868 B.n177 B.n176 10.6151
R1869 B.n180 B.n177 10.6151
R1870 B.n181 B.n180 10.6151
R1871 B.n184 B.n181 10.6151
R1872 B.n185 B.n184 10.6151
R1873 B.n188 B.n185 10.6151
R1874 B.n193 B.n190 10.6151
R1875 B.n194 B.n193 10.6151
R1876 B.n197 B.n194 10.6151
R1877 B.n198 B.n197 10.6151
R1878 B.n201 B.n198 10.6151
R1879 B.n202 B.n201 10.6151
R1880 B.n205 B.n202 10.6151
R1881 B.n206 B.n205 10.6151
R1882 B.n210 B.n209 10.6151
R1883 B.n213 B.n210 10.6151
R1884 B.n214 B.n213 10.6151
R1885 B.n217 B.n214 10.6151
R1886 B.n218 B.n217 10.6151
R1887 B.n221 B.n218 10.6151
R1888 B.n222 B.n221 10.6151
R1889 B.n225 B.n222 10.6151
R1890 B.n226 B.n225 10.6151
R1891 B.n229 B.n226 10.6151
R1892 B.n230 B.n229 10.6151
R1893 B.n233 B.n230 10.6151
R1894 B.n234 B.n233 10.6151
R1895 B.n237 B.n234 10.6151
R1896 B.n238 B.n237 10.6151
R1897 B.n796 B.n238 10.6151
R1898 B.n947 B.n0 8.11757
R1899 B.n947 B.n1 8.11757
R1900 B.n455 B.n401 6.5566
R1901 B.n439 B.n438 6.5566
R1902 B.n190 B.n189 6.5566
R1903 B.n206 B.n156 6.5566
R1904 B.n591 B.t7 4.99766
R1905 B.n272 B.t2 4.99766
R1906 B.t4 B.n910 4.99766
R1907 B.n869 B.t6 4.99766
R1908 B.n458 B.n401 4.05904
R1909 B.n438 B.n437 4.05904
R1910 B.n189 B.n188 4.05904
R1911 B.n209 B.n156 4.05904
R1912 VN.n96 VN.n95 161.3
R1913 VN.n94 VN.n50 161.3
R1914 VN.n93 VN.n92 161.3
R1915 VN.n91 VN.n51 161.3
R1916 VN.n90 VN.n89 161.3
R1917 VN.n88 VN.n52 161.3
R1918 VN.n87 VN.n86 161.3
R1919 VN.n85 VN.n84 161.3
R1920 VN.n83 VN.n54 161.3
R1921 VN.n82 VN.n81 161.3
R1922 VN.n80 VN.n55 161.3
R1923 VN.n79 VN.n78 161.3
R1924 VN.n77 VN.n56 161.3
R1925 VN.n76 VN.n75 161.3
R1926 VN.n74 VN.n57 161.3
R1927 VN.n73 VN.n72 161.3
R1928 VN.n71 VN.n58 161.3
R1929 VN.n70 VN.n69 161.3
R1930 VN.n68 VN.n59 161.3
R1931 VN.n67 VN.n66 161.3
R1932 VN.n65 VN.n60 161.3
R1933 VN.n64 VN.n63 161.3
R1934 VN.n47 VN.n46 161.3
R1935 VN.n45 VN.n1 161.3
R1936 VN.n44 VN.n43 161.3
R1937 VN.n42 VN.n2 161.3
R1938 VN.n41 VN.n40 161.3
R1939 VN.n39 VN.n3 161.3
R1940 VN.n38 VN.n37 161.3
R1941 VN.n36 VN.n35 161.3
R1942 VN.n34 VN.n5 161.3
R1943 VN.n33 VN.n32 161.3
R1944 VN.n31 VN.n6 161.3
R1945 VN.n30 VN.n29 161.3
R1946 VN.n28 VN.n7 161.3
R1947 VN.n27 VN.n26 161.3
R1948 VN.n25 VN.n8 161.3
R1949 VN.n24 VN.n23 161.3
R1950 VN.n22 VN.n9 161.3
R1951 VN.n21 VN.n20 161.3
R1952 VN.n19 VN.n10 161.3
R1953 VN.n18 VN.n17 161.3
R1954 VN.n16 VN.n11 161.3
R1955 VN.n15 VN.n14 161.3
R1956 VN.n48 VN.n0 81.2593
R1957 VN.n97 VN.n49 81.2593
R1958 VN.n13 VN.n12 70.1236
R1959 VN.n62 VN.n61 70.1236
R1960 VN.n62 VN.t4 58.0019
R1961 VN.n13 VN.t0 58.0019
R1962 VN.n21 VN.n10 56.5193
R1963 VN.n29 VN.n6 56.5193
R1964 VN.n70 VN.n59 56.5193
R1965 VN.n78 VN.n55 56.5193
R1966 VN.n40 VN.n2 51.663
R1967 VN.n89 VN.n51 51.663
R1968 VN VN.n97 50.4639
R1969 VN.n44 VN.n2 29.3238
R1970 VN.n93 VN.n51 29.3238
R1971 VN.n8 VN.t2 26.0965
R1972 VN.n12 VN.t8 26.0965
R1973 VN.n4 VN.t9 26.0965
R1974 VN.n0 VN.t1 26.0965
R1975 VN.n57 VN.t7 26.0965
R1976 VN.n61 VN.t5 26.0965
R1977 VN.n53 VN.t3 26.0965
R1978 VN.n49 VN.t6 26.0965
R1979 VN.n16 VN.n15 24.4675
R1980 VN.n17 VN.n16 24.4675
R1981 VN.n17 VN.n10 24.4675
R1982 VN.n22 VN.n21 24.4675
R1983 VN.n23 VN.n22 24.4675
R1984 VN.n23 VN.n8 24.4675
R1985 VN.n27 VN.n8 24.4675
R1986 VN.n28 VN.n27 24.4675
R1987 VN.n29 VN.n28 24.4675
R1988 VN.n33 VN.n6 24.4675
R1989 VN.n34 VN.n33 24.4675
R1990 VN.n35 VN.n34 24.4675
R1991 VN.n39 VN.n38 24.4675
R1992 VN.n40 VN.n39 24.4675
R1993 VN.n45 VN.n44 24.4675
R1994 VN.n46 VN.n45 24.4675
R1995 VN.n66 VN.n59 24.4675
R1996 VN.n66 VN.n65 24.4675
R1997 VN.n65 VN.n64 24.4675
R1998 VN.n78 VN.n77 24.4675
R1999 VN.n77 VN.n76 24.4675
R2000 VN.n76 VN.n57 24.4675
R2001 VN.n72 VN.n57 24.4675
R2002 VN.n72 VN.n71 24.4675
R2003 VN.n71 VN.n70 24.4675
R2004 VN.n89 VN.n88 24.4675
R2005 VN.n88 VN.n87 24.4675
R2006 VN.n84 VN.n83 24.4675
R2007 VN.n83 VN.n82 24.4675
R2008 VN.n82 VN.n55 24.4675
R2009 VN.n95 VN.n94 24.4675
R2010 VN.n94 VN.n93 24.4675
R2011 VN.n38 VN.n4 20.0634
R2012 VN.n87 VN.n53 20.0634
R2013 VN.n46 VN.n0 8.80862
R2014 VN.n95 VN.n49 8.80862
R2015 VN.n63 VN.n62 4.46393
R2016 VN.n14 VN.n13 4.46393
R2017 VN.n15 VN.n12 4.40456
R2018 VN.n35 VN.n4 4.40456
R2019 VN.n64 VN.n61 4.40456
R2020 VN.n84 VN.n53 4.40456
R2021 VN.n97 VN.n96 0.354971
R2022 VN.n48 VN.n47 0.354971
R2023 VN VN.n48 0.26696
R2024 VN.n96 VN.n50 0.189894
R2025 VN.n92 VN.n50 0.189894
R2026 VN.n92 VN.n91 0.189894
R2027 VN.n91 VN.n90 0.189894
R2028 VN.n90 VN.n52 0.189894
R2029 VN.n86 VN.n52 0.189894
R2030 VN.n86 VN.n85 0.189894
R2031 VN.n85 VN.n54 0.189894
R2032 VN.n81 VN.n54 0.189894
R2033 VN.n81 VN.n80 0.189894
R2034 VN.n80 VN.n79 0.189894
R2035 VN.n79 VN.n56 0.189894
R2036 VN.n75 VN.n56 0.189894
R2037 VN.n75 VN.n74 0.189894
R2038 VN.n74 VN.n73 0.189894
R2039 VN.n73 VN.n58 0.189894
R2040 VN.n69 VN.n58 0.189894
R2041 VN.n69 VN.n68 0.189894
R2042 VN.n68 VN.n67 0.189894
R2043 VN.n67 VN.n60 0.189894
R2044 VN.n63 VN.n60 0.189894
R2045 VN.n14 VN.n11 0.189894
R2046 VN.n18 VN.n11 0.189894
R2047 VN.n19 VN.n18 0.189894
R2048 VN.n20 VN.n19 0.189894
R2049 VN.n20 VN.n9 0.189894
R2050 VN.n24 VN.n9 0.189894
R2051 VN.n25 VN.n24 0.189894
R2052 VN.n26 VN.n25 0.189894
R2053 VN.n26 VN.n7 0.189894
R2054 VN.n30 VN.n7 0.189894
R2055 VN.n31 VN.n30 0.189894
R2056 VN.n32 VN.n31 0.189894
R2057 VN.n32 VN.n5 0.189894
R2058 VN.n36 VN.n5 0.189894
R2059 VN.n37 VN.n36 0.189894
R2060 VN.n37 VN.n3 0.189894
R2061 VN.n41 VN.n3 0.189894
R2062 VN.n42 VN.n41 0.189894
R2063 VN.n43 VN.n42 0.189894
R2064 VN.n43 VN.n1 0.189894
R2065 VN.n47 VN.n1 0.189894
R2066 VDD2.n1 VDD2.t9 85.0341
R2067 VDD2.n4 VDD2.t3 81.9393
R2068 VDD2.n3 VDD2.n2 78.5959
R2069 VDD2 VDD2.n7 78.5932
R2070 VDD2.n6 VDD2.n5 76.3303
R2071 VDD2.n1 VDD2.n0 76.3301
R2072 VDD2.n4 VDD2.n3 41.4588
R2073 VDD2.n7 VDD2.t4 5.60957
R2074 VDD2.n7 VDD2.t5 5.60957
R2075 VDD2.n5 VDD2.t6 5.60957
R2076 VDD2.n5 VDD2.t2 5.60957
R2077 VDD2.n2 VDD2.t0 5.60957
R2078 VDD2.n2 VDD2.t8 5.60957
R2079 VDD2.n0 VDD2.t1 5.60957
R2080 VDD2.n0 VDD2.t7 5.60957
R2081 VDD2.n6 VDD2.n4 3.09533
R2082 VDD2 VDD2.n6 0.832397
R2083 VDD2.n3 VDD2.n1 0.718861
C0 VN VDD2 3.64861f
C1 VDD1 VN 0.15962f
C2 VN VP 7.81468f
C3 VDD2 VTAIL 7.2048f
C4 VDD1 VTAIL 7.14727f
C5 VDD1 VDD2 2.60402f
C6 VP VTAIL 5.287971f
C7 VP VDD2 0.672856f
C8 VDD1 VP 4.15803f
C9 VN VTAIL 5.27383f
C10 VDD2 B 6.587092f
C11 VDD1 B 6.479705f
C12 VTAIL B 4.737021f
C13 VN B 20.519428f
C14 VP B 18.984869f
C15 VDD2.t9 B 0.788957f
C16 VDD2.t1 B 0.078693f
C17 VDD2.t7 B 0.078693f
C18 VDD2.n0 B 0.604684f
C19 VDD2.n1 B 1.10231f
C20 VDD2.t0 B 0.078693f
C21 VDD2.t8 B 0.078693f
C22 VDD2.n2 B 0.62529f
C23 VDD2.n3 B 3.07304f
C24 VDD2.t3 B 0.768606f
C25 VDD2.n4 B 3.02982f
C26 VDD2.t6 B 0.078693f
C27 VDD2.t2 B 0.078693f
C28 VDD2.n5 B 0.604685f
C29 VDD2.n6 B 0.572812f
C30 VDD2.t4 B 0.078693f
C31 VDD2.t5 B 0.078693f
C32 VDD2.n7 B 0.625248f
C33 VN.t1 B 0.693762f
C34 VN.n0 B 0.361505f
C35 VN.n1 B 0.023755f
C36 VN.n2 B 0.023572f
C37 VN.n3 B 0.023755f
C38 VN.t9 B 0.693762f
C39 VN.n4 B 0.277226f
C40 VN.n5 B 0.023755f
C41 VN.n6 B 0.031701f
C42 VN.n7 B 0.023755f
C43 VN.t2 B 0.693762f
C44 VN.n8 B 0.299641f
C45 VN.n9 B 0.023755f
C46 VN.n10 B 0.031701f
C47 VN.n11 B 0.023755f
C48 VN.t8 B 0.693762f
C49 VN.n12 B 0.350092f
C50 VN.t0 B 0.936499f
C51 VN.n13 B 0.347861f
C52 VN.n14 B 0.279825f
C53 VN.n15 B 0.02635f
C54 VN.n16 B 0.044273f
C55 VN.n17 B 0.044273f
C56 VN.n18 B 0.023755f
C57 VN.n19 B 0.023755f
C58 VN.n20 B 0.023755f
C59 VN.n21 B 0.037659f
C60 VN.n22 B 0.044273f
C61 VN.n23 B 0.044273f
C62 VN.n24 B 0.023755f
C63 VN.n25 B 0.023755f
C64 VN.n26 B 0.023755f
C65 VN.n27 B 0.044273f
C66 VN.n28 B 0.044273f
C67 VN.n29 B 0.037659f
C68 VN.n30 B 0.023755f
C69 VN.n31 B 0.023755f
C70 VN.n32 B 0.023755f
C71 VN.n33 B 0.044273f
C72 VN.n34 B 0.044273f
C73 VN.n35 B 0.02635f
C74 VN.n36 B 0.023755f
C75 VN.n37 B 0.023755f
C76 VN.n38 B 0.040339f
C77 VN.n39 B 0.044273f
C78 VN.n40 B 0.042893f
C79 VN.n41 B 0.023755f
C80 VN.n42 B 0.023755f
C81 VN.n43 B 0.023755f
C82 VN.n44 B 0.047169f
C83 VN.n45 B 0.044273f
C84 VN.n46 B 0.030284f
C85 VN.n47 B 0.03834f
C86 VN.n48 B 0.061996f
C87 VN.t6 B 0.693762f
C88 VN.n49 B 0.361505f
C89 VN.n50 B 0.023755f
C90 VN.n51 B 0.023572f
C91 VN.n52 B 0.023755f
C92 VN.t3 B 0.693762f
C93 VN.n53 B 0.277226f
C94 VN.n54 B 0.023755f
C95 VN.n55 B 0.031701f
C96 VN.n56 B 0.023755f
C97 VN.t7 B 0.693762f
C98 VN.n57 B 0.299641f
C99 VN.n58 B 0.023755f
C100 VN.n59 B 0.031701f
C101 VN.n60 B 0.023755f
C102 VN.t5 B 0.693762f
C103 VN.n61 B 0.350092f
C104 VN.t4 B 0.936499f
C105 VN.n62 B 0.347861f
C106 VN.n63 B 0.279825f
C107 VN.n64 B 0.02635f
C108 VN.n65 B 0.044273f
C109 VN.n66 B 0.044273f
C110 VN.n67 B 0.023755f
C111 VN.n68 B 0.023755f
C112 VN.n69 B 0.023755f
C113 VN.n70 B 0.037659f
C114 VN.n71 B 0.044273f
C115 VN.n72 B 0.044273f
C116 VN.n73 B 0.023755f
C117 VN.n74 B 0.023755f
C118 VN.n75 B 0.023755f
C119 VN.n76 B 0.044273f
C120 VN.n77 B 0.044273f
C121 VN.n78 B 0.037659f
C122 VN.n79 B 0.023755f
C123 VN.n80 B 0.023755f
C124 VN.n81 B 0.023755f
C125 VN.n82 B 0.044273f
C126 VN.n83 B 0.044273f
C127 VN.n84 B 0.02635f
C128 VN.n85 B 0.023755f
C129 VN.n86 B 0.023755f
C130 VN.n87 B 0.040339f
C131 VN.n88 B 0.044273f
C132 VN.n89 B 0.042893f
C133 VN.n90 B 0.023755f
C134 VN.n91 B 0.023755f
C135 VN.n92 B 0.023755f
C136 VN.n93 B 0.047169f
C137 VN.n94 B 0.044273f
C138 VN.n95 B 0.030284f
C139 VN.n96 B 0.03834f
C140 VN.n97 B 1.37498f
C141 VTAIL.t3 B 0.093015f
C142 VTAIL.t4 B 0.093015f
C143 VTAIL.n0 B 0.645167f
C144 VTAIL.n1 B 0.751797f
C145 VTAIL.t18 B 0.829584f
C146 VTAIL.n2 B 0.897937f
C147 VTAIL.t17 B 0.093015f
C148 VTAIL.t14 B 0.093015f
C149 VTAIL.n3 B 0.645167f
C150 VTAIL.n4 B 0.944455f
C151 VTAIL.t16 B 0.093015f
C152 VTAIL.t15 B 0.093015f
C153 VTAIL.n5 B 0.645167f
C154 VTAIL.n6 B 2.05689f
C155 VTAIL.t0 B 0.093015f
C156 VTAIL.t7 B 0.093015f
C157 VTAIL.n7 B 0.645171f
C158 VTAIL.n8 B 2.05688f
C159 VTAIL.t1 B 0.093015f
C160 VTAIL.t2 B 0.093015f
C161 VTAIL.n9 B 0.645171f
C162 VTAIL.n10 B 0.944452f
C163 VTAIL.t8 B 0.829589f
C164 VTAIL.n11 B 0.897932f
C165 VTAIL.t12 B 0.093015f
C166 VTAIL.t19 B 0.093015f
C167 VTAIL.n12 B 0.645171f
C168 VTAIL.n13 B 0.828672f
C169 VTAIL.t11 B 0.093015f
C170 VTAIL.t10 B 0.093015f
C171 VTAIL.n14 B 0.645171f
C172 VTAIL.n15 B 0.944452f
C173 VTAIL.t13 B 0.829584f
C174 VTAIL.n16 B 1.79363f
C175 VTAIL.t9 B 0.829584f
C176 VTAIL.n17 B 1.79363f
C177 VTAIL.t5 B 0.093015f
C178 VTAIL.t6 B 0.093015f
C179 VTAIL.n18 B 0.645167f
C180 VTAIL.n19 B 0.688813f
C181 VDD1.t8 B 0.812084f
C182 VDD1.t2 B 0.081f
C183 VDD1.t1 B 0.081f
C184 VDD1.n0 B 0.622409f
C185 VDD1.n1 B 1.14429f
C186 VDD1.t0 B 0.812081f
C187 VDD1.t6 B 0.081f
C188 VDD1.t3 B 0.081f
C189 VDD1.n2 B 0.622407f
C190 VDD1.n3 B 1.13461f
C191 VDD1.t9 B 0.081f
C192 VDD1.t7 B 0.081f
C193 VDD1.n4 B 0.643617f
C194 VDD1.n5 B 3.31994f
C195 VDD1.t4 B 0.081f
C196 VDD1.t5 B 0.081f
C197 VDD1.n6 B 0.622406f
C198 VDD1.n7 B 3.22859f
C199 VP.t1 B 0.720127f
C200 VP.n0 B 0.375243f
C201 VP.n1 B 0.024658f
C202 VP.n2 B 0.024468f
C203 VP.n3 B 0.024658f
C204 VP.t5 B 0.720127f
C205 VP.n4 B 0.287762f
C206 VP.n5 B 0.024658f
C207 VP.n6 B 0.032906f
C208 VP.n7 B 0.024658f
C209 VP.t2 B 0.720127f
C210 VP.n8 B 0.311029f
C211 VP.n9 B 0.024658f
C212 VP.n10 B 0.032906f
C213 VP.n11 B 0.024658f
C214 VP.t4 B 0.720127f
C215 VP.n12 B 0.287762f
C216 VP.n13 B 0.024658f
C217 VP.n14 B 0.024468f
C218 VP.n15 B 0.024658f
C219 VP.t3 B 0.720127f
C220 VP.n16 B 0.375243f
C221 VP.t6 B 0.720127f
C222 VP.n17 B 0.375243f
C223 VP.n18 B 0.024658f
C224 VP.n19 B 0.024468f
C225 VP.n20 B 0.024658f
C226 VP.t9 B 0.720127f
C227 VP.n21 B 0.287762f
C228 VP.n22 B 0.024658f
C229 VP.n23 B 0.032906f
C230 VP.n24 B 0.024658f
C231 VP.t8 B 0.720127f
C232 VP.n25 B 0.311029f
C233 VP.n26 B 0.024658f
C234 VP.n27 B 0.032906f
C235 VP.n28 B 0.024658f
C236 VP.t0 B 0.720127f
C237 VP.n29 B 0.363396f
C238 VP.t7 B 0.972088f
C239 VP.n30 B 0.361081f
C240 VP.n31 B 0.29046f
C241 VP.n32 B 0.027351f
C242 VP.n33 B 0.045956f
C243 VP.n34 B 0.045956f
C244 VP.n35 B 0.024658f
C245 VP.n36 B 0.024658f
C246 VP.n37 B 0.024658f
C247 VP.n38 B 0.03909f
C248 VP.n39 B 0.045956f
C249 VP.n40 B 0.045956f
C250 VP.n41 B 0.024658f
C251 VP.n42 B 0.024658f
C252 VP.n43 B 0.024658f
C253 VP.n44 B 0.045956f
C254 VP.n45 B 0.045956f
C255 VP.n46 B 0.03909f
C256 VP.n47 B 0.024658f
C257 VP.n48 B 0.024658f
C258 VP.n49 B 0.024658f
C259 VP.n50 B 0.045956f
C260 VP.n51 B 0.045956f
C261 VP.n52 B 0.027351f
C262 VP.n53 B 0.024658f
C263 VP.n54 B 0.024658f
C264 VP.n55 B 0.041872f
C265 VP.n56 B 0.045956f
C266 VP.n57 B 0.044523f
C267 VP.n58 B 0.024658f
C268 VP.n59 B 0.024658f
C269 VP.n60 B 0.024658f
C270 VP.n61 B 0.048962f
C271 VP.n62 B 0.045956f
C272 VP.n63 B 0.031435f
C273 VP.n64 B 0.039797f
C274 VP.n65 B 1.41715f
C275 VP.n66 B 1.43478f
C276 VP.n67 B 0.039797f
C277 VP.n68 B 0.031435f
C278 VP.n69 B 0.045956f
C279 VP.n70 B 0.048962f
C280 VP.n71 B 0.024658f
C281 VP.n72 B 0.024658f
C282 VP.n73 B 0.024658f
C283 VP.n74 B 0.044523f
C284 VP.n75 B 0.045956f
C285 VP.n76 B 0.041872f
C286 VP.n77 B 0.024658f
C287 VP.n78 B 0.024658f
C288 VP.n79 B 0.027351f
C289 VP.n80 B 0.045956f
C290 VP.n81 B 0.045956f
C291 VP.n82 B 0.024658f
C292 VP.n83 B 0.024658f
C293 VP.n84 B 0.024658f
C294 VP.n85 B 0.03909f
C295 VP.n86 B 0.045956f
C296 VP.n87 B 0.045956f
C297 VP.n88 B 0.024658f
C298 VP.n89 B 0.024658f
C299 VP.n90 B 0.024658f
C300 VP.n91 B 0.045956f
C301 VP.n92 B 0.045956f
C302 VP.n93 B 0.03909f
C303 VP.n94 B 0.024658f
C304 VP.n95 B 0.024658f
C305 VP.n96 B 0.024658f
C306 VP.n97 B 0.045956f
C307 VP.n98 B 0.045956f
C308 VP.n99 B 0.027351f
C309 VP.n100 B 0.024658f
C310 VP.n101 B 0.024658f
C311 VP.n102 B 0.041872f
C312 VP.n103 B 0.045956f
C313 VP.n104 B 0.044523f
C314 VP.n105 B 0.024658f
C315 VP.n106 B 0.024658f
C316 VP.n107 B 0.024658f
C317 VP.n108 B 0.048962f
C318 VP.n109 B 0.045956f
C319 VP.n110 B 0.031435f
C320 VP.n111 B 0.039797f
C321 VP.n112 B 0.064352f
.ends

