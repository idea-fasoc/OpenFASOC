* NGSPICE file created from diff_pair_sample_0144.ext - technology: sky130A

.subckt diff_pair_sample_0144 VTAIL VN VP B VDD2 VDD1
X0 B.t23 B.t21 B.t22 B.t15 sky130_fd_pr__nfet_01v8 ad=0.7293 pd=4.52 as=0 ps=0 w=1.87 l=2.76
X1 VTAIL.t19 VP.t0 VDD1.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=0.30855 pd=2.2 as=0.30855 ps=2.2 w=1.87 l=2.76
X2 VDD1.t8 VP.t1 VTAIL.t18 B.t4 sky130_fd_pr__nfet_01v8 ad=0.7293 pd=4.52 as=0.30855 ps=2.2 w=1.87 l=2.76
X3 VDD2.t9 VN.t0 VTAIL.t9 B.t3 sky130_fd_pr__nfet_01v8 ad=0.7293 pd=4.52 as=0.30855 ps=2.2 w=1.87 l=2.76
X4 VDD1.t1 VP.t2 VTAIL.t17 B.t5 sky130_fd_pr__nfet_01v8 ad=0.30855 pd=2.2 as=0.30855 ps=2.2 w=1.87 l=2.76
X5 VDD1.t5 VP.t3 VTAIL.t16 B.t3 sky130_fd_pr__nfet_01v8 ad=0.7293 pd=4.52 as=0.30855 ps=2.2 w=1.87 l=2.76
X6 VDD1.t4 VP.t4 VTAIL.t15 B.t8 sky130_fd_pr__nfet_01v8 ad=0.30855 pd=2.2 as=0.7293 ps=4.52 w=1.87 l=2.76
X7 B.t20 B.t18 B.t19 B.t11 sky130_fd_pr__nfet_01v8 ad=0.7293 pd=4.52 as=0 ps=0 w=1.87 l=2.76
X8 VDD2.t8 VN.t1 VTAIL.t7 B.t5 sky130_fd_pr__nfet_01v8 ad=0.30855 pd=2.2 as=0.30855 ps=2.2 w=1.87 l=2.76
X9 VDD2.t7 VN.t2 VTAIL.t0 B.t4 sky130_fd_pr__nfet_01v8 ad=0.7293 pd=4.52 as=0.30855 ps=2.2 w=1.87 l=2.76
X10 B.t17 B.t14 B.t16 B.t15 sky130_fd_pr__nfet_01v8 ad=0.7293 pd=4.52 as=0 ps=0 w=1.87 l=2.76
X11 VDD2.t6 VN.t3 VTAIL.t5 B.t8 sky130_fd_pr__nfet_01v8 ad=0.30855 pd=2.2 as=0.7293 ps=4.52 w=1.87 l=2.76
X12 VDD1.t6 VP.t5 VTAIL.t14 B.t9 sky130_fd_pr__nfet_01v8 ad=0.30855 pd=2.2 as=0.7293 ps=4.52 w=1.87 l=2.76
X13 VTAIL.t13 VP.t6 VDD1.t0 B.t7 sky130_fd_pr__nfet_01v8 ad=0.30855 pd=2.2 as=0.30855 ps=2.2 w=1.87 l=2.76
X14 VTAIL.t12 VP.t7 VDD1.t7 B.t1 sky130_fd_pr__nfet_01v8 ad=0.30855 pd=2.2 as=0.30855 ps=2.2 w=1.87 l=2.76
X15 VDD2.t5 VN.t4 VTAIL.t8 B.t9 sky130_fd_pr__nfet_01v8 ad=0.30855 pd=2.2 as=0.7293 ps=4.52 w=1.87 l=2.76
X16 VTAIL.t6 VN.t5 VDD2.t4 B.t2 sky130_fd_pr__nfet_01v8 ad=0.30855 pd=2.2 as=0.30855 ps=2.2 w=1.87 l=2.76
X17 VTAIL.t4 VN.t6 VDD2.t3 B.t1 sky130_fd_pr__nfet_01v8 ad=0.30855 pd=2.2 as=0.30855 ps=2.2 w=1.87 l=2.76
X18 B.t13 B.t10 B.t12 B.t11 sky130_fd_pr__nfet_01v8 ad=0.7293 pd=4.52 as=0 ps=0 w=1.87 l=2.76
X19 VTAIL.t3 VN.t7 VDD2.t2 B.t7 sky130_fd_pr__nfet_01v8 ad=0.30855 pd=2.2 as=0.30855 ps=2.2 w=1.87 l=2.76
X20 VDD2.t1 VN.t8 VTAIL.t2 B.t0 sky130_fd_pr__nfet_01v8 ad=0.30855 pd=2.2 as=0.30855 ps=2.2 w=1.87 l=2.76
X21 VTAIL.t1 VN.t9 VDD2.t0 B.t6 sky130_fd_pr__nfet_01v8 ad=0.30855 pd=2.2 as=0.30855 ps=2.2 w=1.87 l=2.76
X22 VTAIL.t11 VP.t8 VDD1.t9 B.t6 sky130_fd_pr__nfet_01v8 ad=0.30855 pd=2.2 as=0.30855 ps=2.2 w=1.87 l=2.76
X23 VDD1.t3 VP.t9 VTAIL.t10 B.t0 sky130_fd_pr__nfet_01v8 ad=0.30855 pd=2.2 as=0.30855 ps=2.2 w=1.87 l=2.76
R0 B.n611 B.n135 585
R1 B.n135 B.n114 585
R2 B.n613 B.n612 585
R3 B.n615 B.n134 585
R4 B.n618 B.n617 585
R5 B.n619 B.n133 585
R6 B.n621 B.n620 585
R7 B.n623 B.n132 585
R8 B.n626 B.n625 585
R9 B.n627 B.n131 585
R10 B.n629 B.n628 585
R11 B.n631 B.n130 585
R12 B.n634 B.n633 585
R13 B.n636 B.n127 585
R14 B.n638 B.n637 585
R15 B.n640 B.n126 585
R16 B.n643 B.n642 585
R17 B.n644 B.n125 585
R18 B.n646 B.n645 585
R19 B.n648 B.n124 585
R20 B.n651 B.n650 585
R21 B.n652 B.n121 585
R22 B.n655 B.n654 585
R23 B.n657 B.n120 585
R24 B.n660 B.n659 585
R25 B.n661 B.n119 585
R26 B.n663 B.n662 585
R27 B.n665 B.n118 585
R28 B.n668 B.n667 585
R29 B.n669 B.n117 585
R30 B.n671 B.n670 585
R31 B.n673 B.n116 585
R32 B.n676 B.n675 585
R33 B.n677 B.n115 585
R34 B.n610 B.n113 585
R35 B.n680 B.n113 585
R36 B.n609 B.n112 585
R37 B.n681 B.n112 585
R38 B.n608 B.n111 585
R39 B.n682 B.n111 585
R40 B.n607 B.n606 585
R41 B.n606 B.n107 585
R42 B.n605 B.n106 585
R43 B.n688 B.n106 585
R44 B.n604 B.n105 585
R45 B.n689 B.n105 585
R46 B.n603 B.n104 585
R47 B.n690 B.n104 585
R48 B.n602 B.n601 585
R49 B.n601 B.n103 585
R50 B.n600 B.n99 585
R51 B.n696 B.n99 585
R52 B.n599 B.n98 585
R53 B.n697 B.n98 585
R54 B.n598 B.n97 585
R55 B.n698 B.n97 585
R56 B.n597 B.n596 585
R57 B.n596 B.n93 585
R58 B.n595 B.n92 585
R59 B.n704 B.n92 585
R60 B.n594 B.n91 585
R61 B.n705 B.n91 585
R62 B.n593 B.n90 585
R63 B.n706 B.n90 585
R64 B.n592 B.n591 585
R65 B.n591 B.n86 585
R66 B.n590 B.n85 585
R67 B.n712 B.n85 585
R68 B.n589 B.n84 585
R69 B.n713 B.n84 585
R70 B.n588 B.n83 585
R71 B.n714 B.n83 585
R72 B.n587 B.n586 585
R73 B.n586 B.n79 585
R74 B.n585 B.n78 585
R75 B.t8 B.n78 585
R76 B.n584 B.n77 585
R77 B.n720 B.n77 585
R78 B.n583 B.n76 585
R79 B.n721 B.n76 585
R80 B.n582 B.n581 585
R81 B.n581 B.n72 585
R82 B.n580 B.n71 585
R83 B.n727 B.n71 585
R84 B.n579 B.n70 585
R85 B.n728 B.n70 585
R86 B.n578 B.n69 585
R87 B.n729 B.n69 585
R88 B.n577 B.n576 585
R89 B.n576 B.n65 585
R90 B.n575 B.n64 585
R91 B.n735 B.n64 585
R92 B.n574 B.n63 585
R93 B.n736 B.n63 585
R94 B.n573 B.n62 585
R95 B.n737 B.n62 585
R96 B.n572 B.n571 585
R97 B.n571 B.n58 585
R98 B.n570 B.n57 585
R99 B.n743 B.n57 585
R100 B.n569 B.n56 585
R101 B.n744 B.n56 585
R102 B.n568 B.n55 585
R103 B.n745 B.n55 585
R104 B.n567 B.n566 585
R105 B.n566 B.n51 585
R106 B.n565 B.n50 585
R107 B.n751 B.n50 585
R108 B.n564 B.n49 585
R109 B.n752 B.n49 585
R110 B.n563 B.n48 585
R111 B.n753 B.n48 585
R112 B.n562 B.n561 585
R113 B.n561 B.n44 585
R114 B.n560 B.n43 585
R115 B.n759 B.n43 585
R116 B.n559 B.n42 585
R117 B.n760 B.n42 585
R118 B.n558 B.n41 585
R119 B.n761 B.n41 585
R120 B.n557 B.n556 585
R121 B.n556 B.n37 585
R122 B.n555 B.n36 585
R123 B.n767 B.n36 585
R124 B.n554 B.n35 585
R125 B.n768 B.n35 585
R126 B.n553 B.n34 585
R127 B.n769 B.n34 585
R128 B.n552 B.n551 585
R129 B.n551 B.n33 585
R130 B.n550 B.n29 585
R131 B.n775 B.n29 585
R132 B.n549 B.n28 585
R133 B.n776 B.n28 585
R134 B.n548 B.n27 585
R135 B.n777 B.n27 585
R136 B.n547 B.n546 585
R137 B.n546 B.n23 585
R138 B.n545 B.n22 585
R139 B.n783 B.n22 585
R140 B.n544 B.n21 585
R141 B.n784 B.n21 585
R142 B.n543 B.n20 585
R143 B.n785 B.n20 585
R144 B.n542 B.n541 585
R145 B.n541 B.n16 585
R146 B.n540 B.n15 585
R147 B.n791 B.n15 585
R148 B.n539 B.n14 585
R149 B.n792 B.n14 585
R150 B.n538 B.n13 585
R151 B.n793 B.n13 585
R152 B.n537 B.n536 585
R153 B.n536 B.n12 585
R154 B.n535 B.n534 585
R155 B.n535 B.n8 585
R156 B.n533 B.n7 585
R157 B.n800 B.n7 585
R158 B.n532 B.n6 585
R159 B.n801 B.n6 585
R160 B.n531 B.n5 585
R161 B.n802 B.n5 585
R162 B.n530 B.n529 585
R163 B.n529 B.n4 585
R164 B.n528 B.n136 585
R165 B.n528 B.n527 585
R166 B.n518 B.n137 585
R167 B.n138 B.n137 585
R168 B.n520 B.n519 585
R169 B.n521 B.n520 585
R170 B.n517 B.n143 585
R171 B.n143 B.n142 585
R172 B.n516 B.n515 585
R173 B.n515 B.n514 585
R174 B.n145 B.n144 585
R175 B.n146 B.n145 585
R176 B.n507 B.n506 585
R177 B.n508 B.n507 585
R178 B.n505 B.n151 585
R179 B.n151 B.n150 585
R180 B.n504 B.n503 585
R181 B.n503 B.n502 585
R182 B.n153 B.n152 585
R183 B.n154 B.n153 585
R184 B.n495 B.n494 585
R185 B.n496 B.n495 585
R186 B.n493 B.n159 585
R187 B.n159 B.n158 585
R188 B.n492 B.n491 585
R189 B.n491 B.n490 585
R190 B.n161 B.n160 585
R191 B.n483 B.n161 585
R192 B.n482 B.n481 585
R193 B.n484 B.n482 585
R194 B.n480 B.n166 585
R195 B.n166 B.n165 585
R196 B.n479 B.n478 585
R197 B.n478 B.n477 585
R198 B.n168 B.n167 585
R199 B.n169 B.n168 585
R200 B.n470 B.n469 585
R201 B.n471 B.n470 585
R202 B.n468 B.n174 585
R203 B.n174 B.n173 585
R204 B.n467 B.n466 585
R205 B.n466 B.n465 585
R206 B.n176 B.n175 585
R207 B.n177 B.n176 585
R208 B.n458 B.n457 585
R209 B.n459 B.n458 585
R210 B.n456 B.n182 585
R211 B.n182 B.n181 585
R212 B.n455 B.n454 585
R213 B.n454 B.n453 585
R214 B.n184 B.n183 585
R215 B.n185 B.n184 585
R216 B.n446 B.n445 585
R217 B.n447 B.n446 585
R218 B.n444 B.n190 585
R219 B.n190 B.n189 585
R220 B.n443 B.n442 585
R221 B.n442 B.n441 585
R222 B.n192 B.n191 585
R223 B.n193 B.n192 585
R224 B.n434 B.n433 585
R225 B.n435 B.n434 585
R226 B.n432 B.n197 585
R227 B.n201 B.n197 585
R228 B.n431 B.n430 585
R229 B.n430 B.n429 585
R230 B.n199 B.n198 585
R231 B.n200 B.n199 585
R232 B.n422 B.n421 585
R233 B.n423 B.n422 585
R234 B.n420 B.n206 585
R235 B.n206 B.n205 585
R236 B.n419 B.n418 585
R237 B.n418 B.n417 585
R238 B.n208 B.n207 585
R239 B.n209 B.n208 585
R240 B.n410 B.n409 585
R241 B.n411 B.n410 585
R242 B.n408 B.n214 585
R243 B.n214 B.n213 585
R244 B.n407 B.n406 585
R245 B.n406 B.t3 585
R246 B.n216 B.n215 585
R247 B.n217 B.n216 585
R248 B.n399 B.n398 585
R249 B.n400 B.n399 585
R250 B.n397 B.n222 585
R251 B.n222 B.n221 585
R252 B.n396 B.n395 585
R253 B.n395 B.n394 585
R254 B.n224 B.n223 585
R255 B.n225 B.n224 585
R256 B.n387 B.n386 585
R257 B.n388 B.n387 585
R258 B.n385 B.n230 585
R259 B.n230 B.n229 585
R260 B.n384 B.n383 585
R261 B.n383 B.n382 585
R262 B.n232 B.n231 585
R263 B.n233 B.n232 585
R264 B.n375 B.n374 585
R265 B.n376 B.n375 585
R266 B.n373 B.n238 585
R267 B.n238 B.n237 585
R268 B.n372 B.n371 585
R269 B.n371 B.n370 585
R270 B.n240 B.n239 585
R271 B.n363 B.n240 585
R272 B.n362 B.n361 585
R273 B.n364 B.n362 585
R274 B.n360 B.n245 585
R275 B.n245 B.n244 585
R276 B.n359 B.n358 585
R277 B.n358 B.n357 585
R278 B.n247 B.n246 585
R279 B.n248 B.n247 585
R280 B.n350 B.n349 585
R281 B.n351 B.n350 585
R282 B.n348 B.n253 585
R283 B.n253 B.n252 585
R284 B.n347 B.n346 585
R285 B.n346 B.n345 585
R286 B.n342 B.n257 585
R287 B.n341 B.n340 585
R288 B.n338 B.n258 585
R289 B.n338 B.n256 585
R290 B.n337 B.n336 585
R291 B.n335 B.n334 585
R292 B.n333 B.n260 585
R293 B.n331 B.n330 585
R294 B.n329 B.n261 585
R295 B.n328 B.n327 585
R296 B.n325 B.n262 585
R297 B.n323 B.n322 585
R298 B.n321 B.n263 585
R299 B.n319 B.n318 585
R300 B.n316 B.n266 585
R301 B.n314 B.n313 585
R302 B.n312 B.n267 585
R303 B.n311 B.n310 585
R304 B.n308 B.n268 585
R305 B.n306 B.n305 585
R306 B.n304 B.n269 585
R307 B.n303 B.n302 585
R308 B.n300 B.n299 585
R309 B.n298 B.n297 585
R310 B.n296 B.n274 585
R311 B.n294 B.n293 585
R312 B.n292 B.n275 585
R313 B.n291 B.n290 585
R314 B.n288 B.n276 585
R315 B.n286 B.n285 585
R316 B.n284 B.n277 585
R317 B.n283 B.n282 585
R318 B.n280 B.n278 585
R319 B.n255 B.n254 585
R320 B.n344 B.n343 585
R321 B.n345 B.n344 585
R322 B.n251 B.n250 585
R323 B.n252 B.n251 585
R324 B.n353 B.n352 585
R325 B.n352 B.n351 585
R326 B.n354 B.n249 585
R327 B.n249 B.n248 585
R328 B.n356 B.n355 585
R329 B.n357 B.n356 585
R330 B.n243 B.n242 585
R331 B.n244 B.n243 585
R332 B.n366 B.n365 585
R333 B.n365 B.n364 585
R334 B.n367 B.n241 585
R335 B.n363 B.n241 585
R336 B.n369 B.n368 585
R337 B.n370 B.n369 585
R338 B.n236 B.n235 585
R339 B.n237 B.n236 585
R340 B.n378 B.n377 585
R341 B.n377 B.n376 585
R342 B.n379 B.n234 585
R343 B.n234 B.n233 585
R344 B.n381 B.n380 585
R345 B.n382 B.n381 585
R346 B.n228 B.n227 585
R347 B.n229 B.n228 585
R348 B.n390 B.n389 585
R349 B.n389 B.n388 585
R350 B.n391 B.n226 585
R351 B.n226 B.n225 585
R352 B.n393 B.n392 585
R353 B.n394 B.n393 585
R354 B.n220 B.n219 585
R355 B.n221 B.n220 585
R356 B.n402 B.n401 585
R357 B.n401 B.n400 585
R358 B.n403 B.n218 585
R359 B.n218 B.n217 585
R360 B.n405 B.n404 585
R361 B.t3 B.n405 585
R362 B.n212 B.n211 585
R363 B.n213 B.n212 585
R364 B.n413 B.n412 585
R365 B.n412 B.n411 585
R366 B.n414 B.n210 585
R367 B.n210 B.n209 585
R368 B.n416 B.n415 585
R369 B.n417 B.n416 585
R370 B.n204 B.n203 585
R371 B.n205 B.n204 585
R372 B.n425 B.n424 585
R373 B.n424 B.n423 585
R374 B.n426 B.n202 585
R375 B.n202 B.n200 585
R376 B.n428 B.n427 585
R377 B.n429 B.n428 585
R378 B.n196 B.n195 585
R379 B.n201 B.n196 585
R380 B.n437 B.n436 585
R381 B.n436 B.n435 585
R382 B.n438 B.n194 585
R383 B.n194 B.n193 585
R384 B.n440 B.n439 585
R385 B.n441 B.n440 585
R386 B.n188 B.n187 585
R387 B.n189 B.n188 585
R388 B.n449 B.n448 585
R389 B.n448 B.n447 585
R390 B.n450 B.n186 585
R391 B.n186 B.n185 585
R392 B.n452 B.n451 585
R393 B.n453 B.n452 585
R394 B.n180 B.n179 585
R395 B.n181 B.n180 585
R396 B.n461 B.n460 585
R397 B.n460 B.n459 585
R398 B.n462 B.n178 585
R399 B.n178 B.n177 585
R400 B.n464 B.n463 585
R401 B.n465 B.n464 585
R402 B.n172 B.n171 585
R403 B.n173 B.n172 585
R404 B.n473 B.n472 585
R405 B.n472 B.n471 585
R406 B.n474 B.n170 585
R407 B.n170 B.n169 585
R408 B.n476 B.n475 585
R409 B.n477 B.n476 585
R410 B.n164 B.n163 585
R411 B.n165 B.n164 585
R412 B.n486 B.n485 585
R413 B.n485 B.n484 585
R414 B.n487 B.n162 585
R415 B.n483 B.n162 585
R416 B.n489 B.n488 585
R417 B.n490 B.n489 585
R418 B.n157 B.n156 585
R419 B.n158 B.n157 585
R420 B.n498 B.n497 585
R421 B.n497 B.n496 585
R422 B.n499 B.n155 585
R423 B.n155 B.n154 585
R424 B.n501 B.n500 585
R425 B.n502 B.n501 585
R426 B.n149 B.n148 585
R427 B.n150 B.n149 585
R428 B.n510 B.n509 585
R429 B.n509 B.n508 585
R430 B.n511 B.n147 585
R431 B.n147 B.n146 585
R432 B.n513 B.n512 585
R433 B.n514 B.n513 585
R434 B.n141 B.n140 585
R435 B.n142 B.n141 585
R436 B.n523 B.n522 585
R437 B.n522 B.n521 585
R438 B.n524 B.n139 585
R439 B.n139 B.n138 585
R440 B.n526 B.n525 585
R441 B.n527 B.n526 585
R442 B.n3 B.n0 585
R443 B.n4 B.n3 585
R444 B.n799 B.n1 585
R445 B.n800 B.n799 585
R446 B.n798 B.n797 585
R447 B.n798 B.n8 585
R448 B.n796 B.n9 585
R449 B.n12 B.n9 585
R450 B.n795 B.n794 585
R451 B.n794 B.n793 585
R452 B.n11 B.n10 585
R453 B.n792 B.n11 585
R454 B.n790 B.n789 585
R455 B.n791 B.n790 585
R456 B.n788 B.n17 585
R457 B.n17 B.n16 585
R458 B.n787 B.n786 585
R459 B.n786 B.n785 585
R460 B.n19 B.n18 585
R461 B.n784 B.n19 585
R462 B.n782 B.n781 585
R463 B.n783 B.n782 585
R464 B.n780 B.n24 585
R465 B.n24 B.n23 585
R466 B.n779 B.n778 585
R467 B.n778 B.n777 585
R468 B.n26 B.n25 585
R469 B.n776 B.n26 585
R470 B.n774 B.n773 585
R471 B.n775 B.n774 585
R472 B.n772 B.n30 585
R473 B.n33 B.n30 585
R474 B.n771 B.n770 585
R475 B.n770 B.n769 585
R476 B.n32 B.n31 585
R477 B.n768 B.n32 585
R478 B.n766 B.n765 585
R479 B.n767 B.n766 585
R480 B.n764 B.n38 585
R481 B.n38 B.n37 585
R482 B.n763 B.n762 585
R483 B.n762 B.n761 585
R484 B.n40 B.n39 585
R485 B.n760 B.n40 585
R486 B.n758 B.n757 585
R487 B.n759 B.n758 585
R488 B.n756 B.n45 585
R489 B.n45 B.n44 585
R490 B.n755 B.n754 585
R491 B.n754 B.n753 585
R492 B.n47 B.n46 585
R493 B.n752 B.n47 585
R494 B.n750 B.n749 585
R495 B.n751 B.n750 585
R496 B.n748 B.n52 585
R497 B.n52 B.n51 585
R498 B.n747 B.n746 585
R499 B.n746 B.n745 585
R500 B.n54 B.n53 585
R501 B.n744 B.n54 585
R502 B.n742 B.n741 585
R503 B.n743 B.n742 585
R504 B.n740 B.n59 585
R505 B.n59 B.n58 585
R506 B.n739 B.n738 585
R507 B.n738 B.n737 585
R508 B.n61 B.n60 585
R509 B.n736 B.n61 585
R510 B.n734 B.n733 585
R511 B.n735 B.n734 585
R512 B.n732 B.n66 585
R513 B.n66 B.n65 585
R514 B.n731 B.n730 585
R515 B.n730 B.n729 585
R516 B.n68 B.n67 585
R517 B.n728 B.n68 585
R518 B.n726 B.n725 585
R519 B.n727 B.n726 585
R520 B.n724 B.n73 585
R521 B.n73 B.n72 585
R522 B.n723 B.n722 585
R523 B.n722 B.n721 585
R524 B.n75 B.n74 585
R525 B.n720 B.n75 585
R526 B.n719 B.n718 585
R527 B.t8 B.n719 585
R528 B.n717 B.n80 585
R529 B.n80 B.n79 585
R530 B.n716 B.n715 585
R531 B.n715 B.n714 585
R532 B.n82 B.n81 585
R533 B.n713 B.n82 585
R534 B.n711 B.n710 585
R535 B.n712 B.n711 585
R536 B.n709 B.n87 585
R537 B.n87 B.n86 585
R538 B.n708 B.n707 585
R539 B.n707 B.n706 585
R540 B.n89 B.n88 585
R541 B.n705 B.n89 585
R542 B.n703 B.n702 585
R543 B.n704 B.n703 585
R544 B.n701 B.n94 585
R545 B.n94 B.n93 585
R546 B.n700 B.n699 585
R547 B.n699 B.n698 585
R548 B.n96 B.n95 585
R549 B.n697 B.n96 585
R550 B.n695 B.n694 585
R551 B.n696 B.n695 585
R552 B.n693 B.n100 585
R553 B.n103 B.n100 585
R554 B.n692 B.n691 585
R555 B.n691 B.n690 585
R556 B.n102 B.n101 585
R557 B.n689 B.n102 585
R558 B.n687 B.n686 585
R559 B.n688 B.n687 585
R560 B.n685 B.n108 585
R561 B.n108 B.n107 585
R562 B.n684 B.n683 585
R563 B.n683 B.n682 585
R564 B.n110 B.n109 585
R565 B.n681 B.n110 585
R566 B.n679 B.n678 585
R567 B.n680 B.n679 585
R568 B.n803 B.n802 585
R569 B.n801 B.n2 585
R570 B.n679 B.n115 540.549
R571 B.n135 B.n113 540.549
R572 B.n346 B.n255 540.549
R573 B.n344 B.n257 540.549
R574 B.n614 B.n114 256.663
R575 B.n616 B.n114 256.663
R576 B.n622 B.n114 256.663
R577 B.n624 B.n114 256.663
R578 B.n630 B.n114 256.663
R579 B.n632 B.n114 256.663
R580 B.n639 B.n114 256.663
R581 B.n641 B.n114 256.663
R582 B.n647 B.n114 256.663
R583 B.n649 B.n114 256.663
R584 B.n656 B.n114 256.663
R585 B.n658 B.n114 256.663
R586 B.n664 B.n114 256.663
R587 B.n666 B.n114 256.663
R588 B.n672 B.n114 256.663
R589 B.n674 B.n114 256.663
R590 B.n339 B.n256 256.663
R591 B.n259 B.n256 256.663
R592 B.n332 B.n256 256.663
R593 B.n326 B.n256 256.663
R594 B.n324 B.n256 256.663
R595 B.n317 B.n256 256.663
R596 B.n315 B.n256 256.663
R597 B.n309 B.n256 256.663
R598 B.n307 B.n256 256.663
R599 B.n301 B.n256 256.663
R600 B.n273 B.n256 256.663
R601 B.n295 B.n256 256.663
R602 B.n289 B.n256 256.663
R603 B.n287 B.n256 256.663
R604 B.n281 B.n256 256.663
R605 B.n279 B.n256 256.663
R606 B.n805 B.n804 256.663
R607 B.n122 B.t21 224.606
R608 B.n128 B.t14 224.606
R609 B.n270 B.t18 224.606
R610 B.n264 B.t10 224.606
R611 B.n345 B.n256 204.76
R612 B.n680 B.n114 204.76
R613 B.n128 B.t16 180.424
R614 B.n270 B.t20 180.424
R615 B.n122 B.t22 180.424
R616 B.n264 B.t13 180.424
R617 B.n675 B.n673 163.367
R618 B.n671 B.n117 163.367
R619 B.n667 B.n665 163.367
R620 B.n663 B.n119 163.367
R621 B.n659 B.n657 163.367
R622 B.n655 B.n121 163.367
R623 B.n650 B.n648 163.367
R624 B.n646 B.n125 163.367
R625 B.n642 B.n640 163.367
R626 B.n638 B.n127 163.367
R627 B.n633 B.n631 163.367
R628 B.n629 B.n131 163.367
R629 B.n625 B.n623 163.367
R630 B.n621 B.n133 163.367
R631 B.n617 B.n615 163.367
R632 B.n613 B.n135 163.367
R633 B.n346 B.n253 163.367
R634 B.n350 B.n253 163.367
R635 B.n350 B.n247 163.367
R636 B.n358 B.n247 163.367
R637 B.n358 B.n245 163.367
R638 B.n362 B.n245 163.367
R639 B.n362 B.n240 163.367
R640 B.n371 B.n240 163.367
R641 B.n371 B.n238 163.367
R642 B.n375 B.n238 163.367
R643 B.n375 B.n232 163.367
R644 B.n383 B.n232 163.367
R645 B.n383 B.n230 163.367
R646 B.n387 B.n230 163.367
R647 B.n387 B.n224 163.367
R648 B.n395 B.n224 163.367
R649 B.n395 B.n222 163.367
R650 B.n399 B.n222 163.367
R651 B.n399 B.n216 163.367
R652 B.n406 B.n216 163.367
R653 B.n406 B.n214 163.367
R654 B.n410 B.n214 163.367
R655 B.n410 B.n208 163.367
R656 B.n418 B.n208 163.367
R657 B.n418 B.n206 163.367
R658 B.n422 B.n206 163.367
R659 B.n422 B.n199 163.367
R660 B.n430 B.n199 163.367
R661 B.n430 B.n197 163.367
R662 B.n434 B.n197 163.367
R663 B.n434 B.n192 163.367
R664 B.n442 B.n192 163.367
R665 B.n442 B.n190 163.367
R666 B.n446 B.n190 163.367
R667 B.n446 B.n184 163.367
R668 B.n454 B.n184 163.367
R669 B.n454 B.n182 163.367
R670 B.n458 B.n182 163.367
R671 B.n458 B.n176 163.367
R672 B.n466 B.n176 163.367
R673 B.n466 B.n174 163.367
R674 B.n470 B.n174 163.367
R675 B.n470 B.n168 163.367
R676 B.n478 B.n168 163.367
R677 B.n478 B.n166 163.367
R678 B.n482 B.n166 163.367
R679 B.n482 B.n161 163.367
R680 B.n491 B.n161 163.367
R681 B.n491 B.n159 163.367
R682 B.n495 B.n159 163.367
R683 B.n495 B.n153 163.367
R684 B.n503 B.n153 163.367
R685 B.n503 B.n151 163.367
R686 B.n507 B.n151 163.367
R687 B.n507 B.n145 163.367
R688 B.n515 B.n145 163.367
R689 B.n515 B.n143 163.367
R690 B.n520 B.n143 163.367
R691 B.n520 B.n137 163.367
R692 B.n528 B.n137 163.367
R693 B.n529 B.n528 163.367
R694 B.n529 B.n5 163.367
R695 B.n6 B.n5 163.367
R696 B.n7 B.n6 163.367
R697 B.n535 B.n7 163.367
R698 B.n536 B.n535 163.367
R699 B.n536 B.n13 163.367
R700 B.n14 B.n13 163.367
R701 B.n15 B.n14 163.367
R702 B.n541 B.n15 163.367
R703 B.n541 B.n20 163.367
R704 B.n21 B.n20 163.367
R705 B.n22 B.n21 163.367
R706 B.n546 B.n22 163.367
R707 B.n546 B.n27 163.367
R708 B.n28 B.n27 163.367
R709 B.n29 B.n28 163.367
R710 B.n551 B.n29 163.367
R711 B.n551 B.n34 163.367
R712 B.n35 B.n34 163.367
R713 B.n36 B.n35 163.367
R714 B.n556 B.n36 163.367
R715 B.n556 B.n41 163.367
R716 B.n42 B.n41 163.367
R717 B.n43 B.n42 163.367
R718 B.n561 B.n43 163.367
R719 B.n561 B.n48 163.367
R720 B.n49 B.n48 163.367
R721 B.n50 B.n49 163.367
R722 B.n566 B.n50 163.367
R723 B.n566 B.n55 163.367
R724 B.n56 B.n55 163.367
R725 B.n57 B.n56 163.367
R726 B.n571 B.n57 163.367
R727 B.n571 B.n62 163.367
R728 B.n63 B.n62 163.367
R729 B.n64 B.n63 163.367
R730 B.n576 B.n64 163.367
R731 B.n576 B.n69 163.367
R732 B.n70 B.n69 163.367
R733 B.n71 B.n70 163.367
R734 B.n581 B.n71 163.367
R735 B.n581 B.n76 163.367
R736 B.n77 B.n76 163.367
R737 B.n78 B.n77 163.367
R738 B.n586 B.n78 163.367
R739 B.n586 B.n83 163.367
R740 B.n84 B.n83 163.367
R741 B.n85 B.n84 163.367
R742 B.n591 B.n85 163.367
R743 B.n591 B.n90 163.367
R744 B.n91 B.n90 163.367
R745 B.n92 B.n91 163.367
R746 B.n596 B.n92 163.367
R747 B.n596 B.n97 163.367
R748 B.n98 B.n97 163.367
R749 B.n99 B.n98 163.367
R750 B.n601 B.n99 163.367
R751 B.n601 B.n104 163.367
R752 B.n105 B.n104 163.367
R753 B.n106 B.n105 163.367
R754 B.n606 B.n106 163.367
R755 B.n606 B.n111 163.367
R756 B.n112 B.n111 163.367
R757 B.n113 B.n112 163.367
R758 B.n340 B.n338 163.367
R759 B.n338 B.n337 163.367
R760 B.n334 B.n333 163.367
R761 B.n331 B.n261 163.367
R762 B.n327 B.n325 163.367
R763 B.n323 B.n263 163.367
R764 B.n318 B.n316 163.367
R765 B.n314 B.n267 163.367
R766 B.n310 B.n308 163.367
R767 B.n306 B.n269 163.367
R768 B.n302 B.n300 163.367
R769 B.n297 B.n296 163.367
R770 B.n294 B.n275 163.367
R771 B.n290 B.n288 163.367
R772 B.n286 B.n277 163.367
R773 B.n282 B.n280 163.367
R774 B.n344 B.n251 163.367
R775 B.n352 B.n251 163.367
R776 B.n352 B.n249 163.367
R777 B.n356 B.n249 163.367
R778 B.n356 B.n243 163.367
R779 B.n365 B.n243 163.367
R780 B.n365 B.n241 163.367
R781 B.n369 B.n241 163.367
R782 B.n369 B.n236 163.367
R783 B.n377 B.n236 163.367
R784 B.n377 B.n234 163.367
R785 B.n381 B.n234 163.367
R786 B.n381 B.n228 163.367
R787 B.n389 B.n228 163.367
R788 B.n389 B.n226 163.367
R789 B.n393 B.n226 163.367
R790 B.n393 B.n220 163.367
R791 B.n401 B.n220 163.367
R792 B.n401 B.n218 163.367
R793 B.n405 B.n218 163.367
R794 B.n405 B.n212 163.367
R795 B.n412 B.n212 163.367
R796 B.n412 B.n210 163.367
R797 B.n416 B.n210 163.367
R798 B.n416 B.n204 163.367
R799 B.n424 B.n204 163.367
R800 B.n424 B.n202 163.367
R801 B.n428 B.n202 163.367
R802 B.n428 B.n196 163.367
R803 B.n436 B.n196 163.367
R804 B.n436 B.n194 163.367
R805 B.n440 B.n194 163.367
R806 B.n440 B.n188 163.367
R807 B.n448 B.n188 163.367
R808 B.n448 B.n186 163.367
R809 B.n452 B.n186 163.367
R810 B.n452 B.n180 163.367
R811 B.n460 B.n180 163.367
R812 B.n460 B.n178 163.367
R813 B.n464 B.n178 163.367
R814 B.n464 B.n172 163.367
R815 B.n472 B.n172 163.367
R816 B.n472 B.n170 163.367
R817 B.n476 B.n170 163.367
R818 B.n476 B.n164 163.367
R819 B.n485 B.n164 163.367
R820 B.n485 B.n162 163.367
R821 B.n489 B.n162 163.367
R822 B.n489 B.n157 163.367
R823 B.n497 B.n157 163.367
R824 B.n497 B.n155 163.367
R825 B.n501 B.n155 163.367
R826 B.n501 B.n149 163.367
R827 B.n509 B.n149 163.367
R828 B.n509 B.n147 163.367
R829 B.n513 B.n147 163.367
R830 B.n513 B.n141 163.367
R831 B.n522 B.n141 163.367
R832 B.n522 B.n139 163.367
R833 B.n526 B.n139 163.367
R834 B.n526 B.n3 163.367
R835 B.n803 B.n3 163.367
R836 B.n799 B.n2 163.367
R837 B.n799 B.n798 163.367
R838 B.n798 B.n9 163.367
R839 B.n794 B.n9 163.367
R840 B.n794 B.n11 163.367
R841 B.n790 B.n11 163.367
R842 B.n790 B.n17 163.367
R843 B.n786 B.n17 163.367
R844 B.n786 B.n19 163.367
R845 B.n782 B.n19 163.367
R846 B.n782 B.n24 163.367
R847 B.n778 B.n24 163.367
R848 B.n778 B.n26 163.367
R849 B.n774 B.n26 163.367
R850 B.n774 B.n30 163.367
R851 B.n770 B.n30 163.367
R852 B.n770 B.n32 163.367
R853 B.n766 B.n32 163.367
R854 B.n766 B.n38 163.367
R855 B.n762 B.n38 163.367
R856 B.n762 B.n40 163.367
R857 B.n758 B.n40 163.367
R858 B.n758 B.n45 163.367
R859 B.n754 B.n45 163.367
R860 B.n754 B.n47 163.367
R861 B.n750 B.n47 163.367
R862 B.n750 B.n52 163.367
R863 B.n746 B.n52 163.367
R864 B.n746 B.n54 163.367
R865 B.n742 B.n54 163.367
R866 B.n742 B.n59 163.367
R867 B.n738 B.n59 163.367
R868 B.n738 B.n61 163.367
R869 B.n734 B.n61 163.367
R870 B.n734 B.n66 163.367
R871 B.n730 B.n66 163.367
R872 B.n730 B.n68 163.367
R873 B.n726 B.n68 163.367
R874 B.n726 B.n73 163.367
R875 B.n722 B.n73 163.367
R876 B.n722 B.n75 163.367
R877 B.n719 B.n75 163.367
R878 B.n719 B.n80 163.367
R879 B.n715 B.n80 163.367
R880 B.n715 B.n82 163.367
R881 B.n711 B.n82 163.367
R882 B.n711 B.n87 163.367
R883 B.n707 B.n87 163.367
R884 B.n707 B.n89 163.367
R885 B.n703 B.n89 163.367
R886 B.n703 B.n94 163.367
R887 B.n699 B.n94 163.367
R888 B.n699 B.n96 163.367
R889 B.n695 B.n96 163.367
R890 B.n695 B.n100 163.367
R891 B.n691 B.n100 163.367
R892 B.n691 B.n102 163.367
R893 B.n687 B.n102 163.367
R894 B.n687 B.n108 163.367
R895 B.n683 B.n108 163.367
R896 B.n683 B.n110 163.367
R897 B.n679 B.n110 163.367
R898 B.n129 B.t17 120.498
R899 B.n271 B.t19 120.498
R900 B.n123 B.t23 120.498
R901 B.n265 B.t12 120.498
R902 B.n345 B.n252 104.689
R903 B.n351 B.n252 104.689
R904 B.n351 B.n248 104.689
R905 B.n357 B.n248 104.689
R906 B.n357 B.n244 104.689
R907 B.n364 B.n244 104.689
R908 B.n364 B.n363 104.689
R909 B.n370 B.n237 104.689
R910 B.n376 B.n237 104.689
R911 B.n376 B.n233 104.689
R912 B.n382 B.n233 104.689
R913 B.n382 B.n229 104.689
R914 B.n388 B.n229 104.689
R915 B.n388 B.n225 104.689
R916 B.n394 B.n225 104.689
R917 B.n394 B.n221 104.689
R918 B.n400 B.n221 104.689
R919 B.n400 B.n217 104.689
R920 B.t3 B.n217 104.689
R921 B.t3 B.n213 104.689
R922 B.n411 B.n213 104.689
R923 B.n411 B.n209 104.689
R924 B.n417 B.n209 104.689
R925 B.n417 B.n205 104.689
R926 B.n423 B.n205 104.689
R927 B.n423 B.n200 104.689
R928 B.n429 B.n200 104.689
R929 B.n429 B.n201 104.689
R930 B.n435 B.n193 104.689
R931 B.n441 B.n193 104.689
R932 B.n441 B.n189 104.689
R933 B.n447 B.n189 104.689
R934 B.n447 B.n185 104.689
R935 B.n453 B.n185 104.689
R936 B.n453 B.n181 104.689
R937 B.n459 B.n181 104.689
R938 B.n465 B.n177 104.689
R939 B.n465 B.n173 104.689
R940 B.n471 B.n173 104.689
R941 B.n471 B.n169 104.689
R942 B.n477 B.n169 104.689
R943 B.n477 B.n165 104.689
R944 B.n484 B.n165 104.689
R945 B.n484 B.n483 104.689
R946 B.n490 B.n158 104.689
R947 B.n496 B.n158 104.689
R948 B.n496 B.n154 104.689
R949 B.n502 B.n154 104.689
R950 B.n502 B.n150 104.689
R951 B.n508 B.n150 104.689
R952 B.n508 B.n146 104.689
R953 B.n514 B.n146 104.689
R954 B.n521 B.n142 104.689
R955 B.n521 B.n138 104.689
R956 B.n527 B.n138 104.689
R957 B.n527 B.n4 104.689
R958 B.n802 B.n4 104.689
R959 B.n802 B.n801 104.689
R960 B.n801 B.n800 104.689
R961 B.n800 B.n8 104.689
R962 B.n12 B.n8 104.689
R963 B.n793 B.n12 104.689
R964 B.n793 B.n792 104.689
R965 B.n791 B.n16 104.689
R966 B.n785 B.n16 104.689
R967 B.n785 B.n784 104.689
R968 B.n784 B.n783 104.689
R969 B.n783 B.n23 104.689
R970 B.n777 B.n23 104.689
R971 B.n777 B.n776 104.689
R972 B.n776 B.n775 104.689
R973 B.n769 B.n33 104.689
R974 B.n769 B.n768 104.689
R975 B.n768 B.n767 104.689
R976 B.n767 B.n37 104.689
R977 B.n761 B.n37 104.689
R978 B.n761 B.n760 104.689
R979 B.n760 B.n759 104.689
R980 B.n759 B.n44 104.689
R981 B.n753 B.n752 104.689
R982 B.n752 B.n751 104.689
R983 B.n751 B.n51 104.689
R984 B.n745 B.n51 104.689
R985 B.n745 B.n744 104.689
R986 B.n744 B.n743 104.689
R987 B.n743 B.n58 104.689
R988 B.n737 B.n58 104.689
R989 B.n736 B.n735 104.689
R990 B.n735 B.n65 104.689
R991 B.n729 B.n65 104.689
R992 B.n729 B.n728 104.689
R993 B.n728 B.n727 104.689
R994 B.n727 B.n72 104.689
R995 B.n721 B.n72 104.689
R996 B.n721 B.n720 104.689
R997 B.n720 B.t8 104.689
R998 B.t8 B.n79 104.689
R999 B.n714 B.n79 104.689
R1000 B.n714 B.n713 104.689
R1001 B.n713 B.n712 104.689
R1002 B.n712 B.n86 104.689
R1003 B.n706 B.n86 104.689
R1004 B.n706 B.n705 104.689
R1005 B.n705 B.n704 104.689
R1006 B.n704 B.n93 104.689
R1007 B.n698 B.n93 104.689
R1008 B.n698 B.n697 104.689
R1009 B.n697 B.n696 104.689
R1010 B.n690 B.n103 104.689
R1011 B.n690 B.n689 104.689
R1012 B.n689 B.n688 104.689
R1013 B.n688 B.n107 104.689
R1014 B.n682 B.n107 104.689
R1015 B.n682 B.n681 104.689
R1016 B.n681 B.n680 104.689
R1017 B.n435 B.t7 95.4519
R1018 B.n737 B.t2 95.4519
R1019 B.t5 B.n177 86.2146
R1020 B.t0 B.n44 86.2146
R1021 B.n490 B.t6 76.9774
R1022 B.n775 B.t1 76.9774
R1023 B.n363 B.t11 73.8983
R1024 B.n103 B.t15 73.8983
R1025 B.n674 B.n115 71.676
R1026 B.n673 B.n672 71.676
R1027 B.n666 B.n117 71.676
R1028 B.n665 B.n664 71.676
R1029 B.n658 B.n119 71.676
R1030 B.n657 B.n656 71.676
R1031 B.n649 B.n121 71.676
R1032 B.n648 B.n647 71.676
R1033 B.n641 B.n125 71.676
R1034 B.n640 B.n639 71.676
R1035 B.n632 B.n127 71.676
R1036 B.n631 B.n630 71.676
R1037 B.n624 B.n131 71.676
R1038 B.n623 B.n622 71.676
R1039 B.n616 B.n133 71.676
R1040 B.n615 B.n614 71.676
R1041 B.n614 B.n613 71.676
R1042 B.n617 B.n616 71.676
R1043 B.n622 B.n621 71.676
R1044 B.n625 B.n624 71.676
R1045 B.n630 B.n629 71.676
R1046 B.n633 B.n632 71.676
R1047 B.n639 B.n638 71.676
R1048 B.n642 B.n641 71.676
R1049 B.n647 B.n646 71.676
R1050 B.n650 B.n649 71.676
R1051 B.n656 B.n655 71.676
R1052 B.n659 B.n658 71.676
R1053 B.n664 B.n663 71.676
R1054 B.n667 B.n666 71.676
R1055 B.n672 B.n671 71.676
R1056 B.n675 B.n674 71.676
R1057 B.n339 B.n257 71.676
R1058 B.n337 B.n259 71.676
R1059 B.n333 B.n332 71.676
R1060 B.n326 B.n261 71.676
R1061 B.n325 B.n324 71.676
R1062 B.n317 B.n263 71.676
R1063 B.n316 B.n315 71.676
R1064 B.n309 B.n267 71.676
R1065 B.n308 B.n307 71.676
R1066 B.n301 B.n269 71.676
R1067 B.n300 B.n273 71.676
R1068 B.n296 B.n295 71.676
R1069 B.n289 B.n275 71.676
R1070 B.n288 B.n287 71.676
R1071 B.n281 B.n277 71.676
R1072 B.n280 B.n279 71.676
R1073 B.n340 B.n339 71.676
R1074 B.n334 B.n259 71.676
R1075 B.n332 B.n331 71.676
R1076 B.n327 B.n326 71.676
R1077 B.n324 B.n323 71.676
R1078 B.n318 B.n317 71.676
R1079 B.n315 B.n314 71.676
R1080 B.n310 B.n309 71.676
R1081 B.n307 B.n306 71.676
R1082 B.n302 B.n301 71.676
R1083 B.n297 B.n273 71.676
R1084 B.n295 B.n294 71.676
R1085 B.n290 B.n289 71.676
R1086 B.n287 B.n286 71.676
R1087 B.n282 B.n281 71.676
R1088 B.n279 B.n255 71.676
R1089 B.n804 B.n803 71.676
R1090 B.n804 B.n2 71.676
R1091 B.t9 B.n142 67.7402
R1092 B.n792 B.t4 67.7402
R1093 B.n123 B.n122 59.9278
R1094 B.n129 B.n128 59.9278
R1095 B.n271 B.n270 59.9278
R1096 B.n265 B.n264 59.9278
R1097 B.n653 B.n123 59.5399
R1098 B.n635 B.n129 59.5399
R1099 B.n272 B.n271 59.5399
R1100 B.n320 B.n265 59.5399
R1101 B.n514 B.t9 36.9494
R1102 B.t4 B.n791 36.9494
R1103 B.n343 B.n342 35.1225
R1104 B.n347 B.n254 35.1225
R1105 B.n611 B.n610 35.1225
R1106 B.n678 B.n677 35.1225
R1107 B.n370 B.t11 30.7913
R1108 B.n696 B.t15 30.7913
R1109 B.n483 B.t6 27.7122
R1110 B.n33 B.t1 27.7122
R1111 B.n459 B.t5 18.475
R1112 B.n753 B.t0 18.475
R1113 B B.n805 18.0485
R1114 B.n343 B.n250 10.6151
R1115 B.n353 B.n250 10.6151
R1116 B.n354 B.n353 10.6151
R1117 B.n355 B.n354 10.6151
R1118 B.n355 B.n242 10.6151
R1119 B.n366 B.n242 10.6151
R1120 B.n367 B.n366 10.6151
R1121 B.n368 B.n367 10.6151
R1122 B.n368 B.n235 10.6151
R1123 B.n378 B.n235 10.6151
R1124 B.n379 B.n378 10.6151
R1125 B.n380 B.n379 10.6151
R1126 B.n380 B.n227 10.6151
R1127 B.n390 B.n227 10.6151
R1128 B.n391 B.n390 10.6151
R1129 B.n392 B.n391 10.6151
R1130 B.n392 B.n219 10.6151
R1131 B.n402 B.n219 10.6151
R1132 B.n403 B.n402 10.6151
R1133 B.n404 B.n403 10.6151
R1134 B.n404 B.n211 10.6151
R1135 B.n413 B.n211 10.6151
R1136 B.n414 B.n413 10.6151
R1137 B.n415 B.n414 10.6151
R1138 B.n415 B.n203 10.6151
R1139 B.n425 B.n203 10.6151
R1140 B.n426 B.n425 10.6151
R1141 B.n427 B.n426 10.6151
R1142 B.n427 B.n195 10.6151
R1143 B.n437 B.n195 10.6151
R1144 B.n438 B.n437 10.6151
R1145 B.n439 B.n438 10.6151
R1146 B.n439 B.n187 10.6151
R1147 B.n449 B.n187 10.6151
R1148 B.n450 B.n449 10.6151
R1149 B.n451 B.n450 10.6151
R1150 B.n451 B.n179 10.6151
R1151 B.n461 B.n179 10.6151
R1152 B.n462 B.n461 10.6151
R1153 B.n463 B.n462 10.6151
R1154 B.n463 B.n171 10.6151
R1155 B.n473 B.n171 10.6151
R1156 B.n474 B.n473 10.6151
R1157 B.n475 B.n474 10.6151
R1158 B.n475 B.n163 10.6151
R1159 B.n486 B.n163 10.6151
R1160 B.n487 B.n486 10.6151
R1161 B.n488 B.n487 10.6151
R1162 B.n488 B.n156 10.6151
R1163 B.n498 B.n156 10.6151
R1164 B.n499 B.n498 10.6151
R1165 B.n500 B.n499 10.6151
R1166 B.n500 B.n148 10.6151
R1167 B.n510 B.n148 10.6151
R1168 B.n511 B.n510 10.6151
R1169 B.n512 B.n511 10.6151
R1170 B.n512 B.n140 10.6151
R1171 B.n523 B.n140 10.6151
R1172 B.n524 B.n523 10.6151
R1173 B.n525 B.n524 10.6151
R1174 B.n525 B.n0 10.6151
R1175 B.n342 B.n341 10.6151
R1176 B.n341 B.n258 10.6151
R1177 B.n336 B.n258 10.6151
R1178 B.n336 B.n335 10.6151
R1179 B.n335 B.n260 10.6151
R1180 B.n330 B.n260 10.6151
R1181 B.n330 B.n329 10.6151
R1182 B.n329 B.n328 10.6151
R1183 B.n328 B.n262 10.6151
R1184 B.n322 B.n262 10.6151
R1185 B.n322 B.n321 10.6151
R1186 B.n319 B.n266 10.6151
R1187 B.n313 B.n266 10.6151
R1188 B.n313 B.n312 10.6151
R1189 B.n312 B.n311 10.6151
R1190 B.n311 B.n268 10.6151
R1191 B.n305 B.n268 10.6151
R1192 B.n305 B.n304 10.6151
R1193 B.n304 B.n303 10.6151
R1194 B.n299 B.n298 10.6151
R1195 B.n298 B.n274 10.6151
R1196 B.n293 B.n274 10.6151
R1197 B.n293 B.n292 10.6151
R1198 B.n292 B.n291 10.6151
R1199 B.n291 B.n276 10.6151
R1200 B.n285 B.n276 10.6151
R1201 B.n285 B.n284 10.6151
R1202 B.n284 B.n283 10.6151
R1203 B.n283 B.n278 10.6151
R1204 B.n278 B.n254 10.6151
R1205 B.n348 B.n347 10.6151
R1206 B.n349 B.n348 10.6151
R1207 B.n349 B.n246 10.6151
R1208 B.n359 B.n246 10.6151
R1209 B.n360 B.n359 10.6151
R1210 B.n361 B.n360 10.6151
R1211 B.n361 B.n239 10.6151
R1212 B.n372 B.n239 10.6151
R1213 B.n373 B.n372 10.6151
R1214 B.n374 B.n373 10.6151
R1215 B.n374 B.n231 10.6151
R1216 B.n384 B.n231 10.6151
R1217 B.n385 B.n384 10.6151
R1218 B.n386 B.n385 10.6151
R1219 B.n386 B.n223 10.6151
R1220 B.n396 B.n223 10.6151
R1221 B.n397 B.n396 10.6151
R1222 B.n398 B.n397 10.6151
R1223 B.n398 B.n215 10.6151
R1224 B.n407 B.n215 10.6151
R1225 B.n408 B.n407 10.6151
R1226 B.n409 B.n408 10.6151
R1227 B.n409 B.n207 10.6151
R1228 B.n419 B.n207 10.6151
R1229 B.n420 B.n419 10.6151
R1230 B.n421 B.n420 10.6151
R1231 B.n421 B.n198 10.6151
R1232 B.n431 B.n198 10.6151
R1233 B.n432 B.n431 10.6151
R1234 B.n433 B.n432 10.6151
R1235 B.n433 B.n191 10.6151
R1236 B.n443 B.n191 10.6151
R1237 B.n444 B.n443 10.6151
R1238 B.n445 B.n444 10.6151
R1239 B.n445 B.n183 10.6151
R1240 B.n455 B.n183 10.6151
R1241 B.n456 B.n455 10.6151
R1242 B.n457 B.n456 10.6151
R1243 B.n457 B.n175 10.6151
R1244 B.n467 B.n175 10.6151
R1245 B.n468 B.n467 10.6151
R1246 B.n469 B.n468 10.6151
R1247 B.n469 B.n167 10.6151
R1248 B.n479 B.n167 10.6151
R1249 B.n480 B.n479 10.6151
R1250 B.n481 B.n480 10.6151
R1251 B.n481 B.n160 10.6151
R1252 B.n492 B.n160 10.6151
R1253 B.n493 B.n492 10.6151
R1254 B.n494 B.n493 10.6151
R1255 B.n494 B.n152 10.6151
R1256 B.n504 B.n152 10.6151
R1257 B.n505 B.n504 10.6151
R1258 B.n506 B.n505 10.6151
R1259 B.n506 B.n144 10.6151
R1260 B.n516 B.n144 10.6151
R1261 B.n517 B.n516 10.6151
R1262 B.n519 B.n517 10.6151
R1263 B.n519 B.n518 10.6151
R1264 B.n518 B.n136 10.6151
R1265 B.n530 B.n136 10.6151
R1266 B.n531 B.n530 10.6151
R1267 B.n532 B.n531 10.6151
R1268 B.n533 B.n532 10.6151
R1269 B.n534 B.n533 10.6151
R1270 B.n537 B.n534 10.6151
R1271 B.n538 B.n537 10.6151
R1272 B.n539 B.n538 10.6151
R1273 B.n540 B.n539 10.6151
R1274 B.n542 B.n540 10.6151
R1275 B.n543 B.n542 10.6151
R1276 B.n544 B.n543 10.6151
R1277 B.n545 B.n544 10.6151
R1278 B.n547 B.n545 10.6151
R1279 B.n548 B.n547 10.6151
R1280 B.n549 B.n548 10.6151
R1281 B.n550 B.n549 10.6151
R1282 B.n552 B.n550 10.6151
R1283 B.n553 B.n552 10.6151
R1284 B.n554 B.n553 10.6151
R1285 B.n555 B.n554 10.6151
R1286 B.n557 B.n555 10.6151
R1287 B.n558 B.n557 10.6151
R1288 B.n559 B.n558 10.6151
R1289 B.n560 B.n559 10.6151
R1290 B.n562 B.n560 10.6151
R1291 B.n563 B.n562 10.6151
R1292 B.n564 B.n563 10.6151
R1293 B.n565 B.n564 10.6151
R1294 B.n567 B.n565 10.6151
R1295 B.n568 B.n567 10.6151
R1296 B.n569 B.n568 10.6151
R1297 B.n570 B.n569 10.6151
R1298 B.n572 B.n570 10.6151
R1299 B.n573 B.n572 10.6151
R1300 B.n574 B.n573 10.6151
R1301 B.n575 B.n574 10.6151
R1302 B.n577 B.n575 10.6151
R1303 B.n578 B.n577 10.6151
R1304 B.n579 B.n578 10.6151
R1305 B.n580 B.n579 10.6151
R1306 B.n582 B.n580 10.6151
R1307 B.n583 B.n582 10.6151
R1308 B.n584 B.n583 10.6151
R1309 B.n585 B.n584 10.6151
R1310 B.n587 B.n585 10.6151
R1311 B.n588 B.n587 10.6151
R1312 B.n589 B.n588 10.6151
R1313 B.n590 B.n589 10.6151
R1314 B.n592 B.n590 10.6151
R1315 B.n593 B.n592 10.6151
R1316 B.n594 B.n593 10.6151
R1317 B.n595 B.n594 10.6151
R1318 B.n597 B.n595 10.6151
R1319 B.n598 B.n597 10.6151
R1320 B.n599 B.n598 10.6151
R1321 B.n600 B.n599 10.6151
R1322 B.n602 B.n600 10.6151
R1323 B.n603 B.n602 10.6151
R1324 B.n604 B.n603 10.6151
R1325 B.n605 B.n604 10.6151
R1326 B.n607 B.n605 10.6151
R1327 B.n608 B.n607 10.6151
R1328 B.n609 B.n608 10.6151
R1329 B.n610 B.n609 10.6151
R1330 B.n797 B.n1 10.6151
R1331 B.n797 B.n796 10.6151
R1332 B.n796 B.n795 10.6151
R1333 B.n795 B.n10 10.6151
R1334 B.n789 B.n10 10.6151
R1335 B.n789 B.n788 10.6151
R1336 B.n788 B.n787 10.6151
R1337 B.n787 B.n18 10.6151
R1338 B.n781 B.n18 10.6151
R1339 B.n781 B.n780 10.6151
R1340 B.n780 B.n779 10.6151
R1341 B.n779 B.n25 10.6151
R1342 B.n773 B.n25 10.6151
R1343 B.n773 B.n772 10.6151
R1344 B.n772 B.n771 10.6151
R1345 B.n771 B.n31 10.6151
R1346 B.n765 B.n31 10.6151
R1347 B.n765 B.n764 10.6151
R1348 B.n764 B.n763 10.6151
R1349 B.n763 B.n39 10.6151
R1350 B.n757 B.n39 10.6151
R1351 B.n757 B.n756 10.6151
R1352 B.n756 B.n755 10.6151
R1353 B.n755 B.n46 10.6151
R1354 B.n749 B.n46 10.6151
R1355 B.n749 B.n748 10.6151
R1356 B.n748 B.n747 10.6151
R1357 B.n747 B.n53 10.6151
R1358 B.n741 B.n53 10.6151
R1359 B.n741 B.n740 10.6151
R1360 B.n740 B.n739 10.6151
R1361 B.n739 B.n60 10.6151
R1362 B.n733 B.n60 10.6151
R1363 B.n733 B.n732 10.6151
R1364 B.n732 B.n731 10.6151
R1365 B.n731 B.n67 10.6151
R1366 B.n725 B.n67 10.6151
R1367 B.n725 B.n724 10.6151
R1368 B.n724 B.n723 10.6151
R1369 B.n723 B.n74 10.6151
R1370 B.n718 B.n74 10.6151
R1371 B.n718 B.n717 10.6151
R1372 B.n717 B.n716 10.6151
R1373 B.n716 B.n81 10.6151
R1374 B.n710 B.n81 10.6151
R1375 B.n710 B.n709 10.6151
R1376 B.n709 B.n708 10.6151
R1377 B.n708 B.n88 10.6151
R1378 B.n702 B.n88 10.6151
R1379 B.n702 B.n701 10.6151
R1380 B.n701 B.n700 10.6151
R1381 B.n700 B.n95 10.6151
R1382 B.n694 B.n95 10.6151
R1383 B.n694 B.n693 10.6151
R1384 B.n693 B.n692 10.6151
R1385 B.n692 B.n101 10.6151
R1386 B.n686 B.n101 10.6151
R1387 B.n686 B.n685 10.6151
R1388 B.n685 B.n684 10.6151
R1389 B.n684 B.n109 10.6151
R1390 B.n678 B.n109 10.6151
R1391 B.n677 B.n676 10.6151
R1392 B.n676 B.n116 10.6151
R1393 B.n670 B.n116 10.6151
R1394 B.n670 B.n669 10.6151
R1395 B.n669 B.n668 10.6151
R1396 B.n668 B.n118 10.6151
R1397 B.n662 B.n118 10.6151
R1398 B.n662 B.n661 10.6151
R1399 B.n661 B.n660 10.6151
R1400 B.n660 B.n120 10.6151
R1401 B.n654 B.n120 10.6151
R1402 B.n652 B.n651 10.6151
R1403 B.n651 B.n124 10.6151
R1404 B.n645 B.n124 10.6151
R1405 B.n645 B.n644 10.6151
R1406 B.n644 B.n643 10.6151
R1407 B.n643 B.n126 10.6151
R1408 B.n637 B.n126 10.6151
R1409 B.n637 B.n636 10.6151
R1410 B.n634 B.n130 10.6151
R1411 B.n628 B.n130 10.6151
R1412 B.n628 B.n627 10.6151
R1413 B.n627 B.n626 10.6151
R1414 B.n626 B.n132 10.6151
R1415 B.n620 B.n132 10.6151
R1416 B.n620 B.n619 10.6151
R1417 B.n619 B.n618 10.6151
R1418 B.n618 B.n134 10.6151
R1419 B.n612 B.n134 10.6151
R1420 B.n612 B.n611 10.6151
R1421 B.n201 B.t7 9.23773
R1422 B.t2 B.n736 9.23773
R1423 B.n805 B.n0 8.11757
R1424 B.n805 B.n1 8.11757
R1425 B.n320 B.n319 6.5566
R1426 B.n303 B.n272 6.5566
R1427 B.n653 B.n652 6.5566
R1428 B.n636 B.n635 6.5566
R1429 B.n321 B.n320 4.05904
R1430 B.n299 B.n272 4.05904
R1431 B.n654 B.n653 4.05904
R1432 B.n635 B.n634 4.05904
R1433 VP.n25 VP.n22 161.3
R1434 VP.n27 VP.n26 161.3
R1435 VP.n28 VP.n21 161.3
R1436 VP.n30 VP.n29 161.3
R1437 VP.n31 VP.n20 161.3
R1438 VP.n34 VP.n33 161.3
R1439 VP.n35 VP.n19 161.3
R1440 VP.n37 VP.n36 161.3
R1441 VP.n38 VP.n18 161.3
R1442 VP.n40 VP.n39 161.3
R1443 VP.n41 VP.n17 161.3
R1444 VP.n43 VP.n42 161.3
R1445 VP.n45 VP.n16 161.3
R1446 VP.n47 VP.n46 161.3
R1447 VP.n48 VP.n15 161.3
R1448 VP.n50 VP.n49 161.3
R1449 VP.n51 VP.n14 161.3
R1450 VP.n53 VP.n52 161.3
R1451 VP.n95 VP.n94 161.3
R1452 VP.n93 VP.n1 161.3
R1453 VP.n92 VP.n91 161.3
R1454 VP.n90 VP.n2 161.3
R1455 VP.n89 VP.n88 161.3
R1456 VP.n87 VP.n3 161.3
R1457 VP.n85 VP.n84 161.3
R1458 VP.n83 VP.n4 161.3
R1459 VP.n82 VP.n81 161.3
R1460 VP.n80 VP.n5 161.3
R1461 VP.n79 VP.n78 161.3
R1462 VP.n77 VP.n6 161.3
R1463 VP.n76 VP.n75 161.3
R1464 VP.n73 VP.n7 161.3
R1465 VP.n72 VP.n71 161.3
R1466 VP.n70 VP.n8 161.3
R1467 VP.n69 VP.n68 161.3
R1468 VP.n67 VP.n9 161.3
R1469 VP.n65 VP.n64 161.3
R1470 VP.n63 VP.n10 161.3
R1471 VP.n62 VP.n61 161.3
R1472 VP.n60 VP.n11 161.3
R1473 VP.n59 VP.n58 161.3
R1474 VP.n57 VP.n12 161.3
R1475 VP.n56 VP.n55 69.0258
R1476 VP.n96 VP.n0 69.0258
R1477 VP.n54 VP.n13 69.0258
R1478 VP.n24 VP.n23 56.938
R1479 VP.n72 VP.n8 56.5193
R1480 VP.n81 VP.n80 56.5193
R1481 VP.n39 VP.n38 56.5193
R1482 VP.n30 VP.n21 56.5193
R1483 VP.n61 VP.n60 51.663
R1484 VP.n92 VP.n2 51.663
R1485 VP.n50 VP.n15 51.663
R1486 VP.n23 VP.t1 48.2125
R1487 VP.n56 VP.n54 46.3895
R1488 VP.n60 VP.n59 29.3238
R1489 VP.n93 VP.n92 29.3238
R1490 VP.n51 VP.n50 29.3238
R1491 VP.n59 VP.n12 24.4675
R1492 VP.n61 VP.n10 24.4675
R1493 VP.n65 VP.n10 24.4675
R1494 VP.n68 VP.n67 24.4675
R1495 VP.n68 VP.n8 24.4675
R1496 VP.n73 VP.n72 24.4675
R1497 VP.n75 VP.n73 24.4675
R1498 VP.n79 VP.n6 24.4675
R1499 VP.n80 VP.n79 24.4675
R1500 VP.n81 VP.n4 24.4675
R1501 VP.n85 VP.n4 24.4675
R1502 VP.n88 VP.n87 24.4675
R1503 VP.n88 VP.n2 24.4675
R1504 VP.n94 VP.n93 24.4675
R1505 VP.n52 VP.n51 24.4675
R1506 VP.n39 VP.n17 24.4675
R1507 VP.n43 VP.n17 24.4675
R1508 VP.n46 VP.n45 24.4675
R1509 VP.n46 VP.n15 24.4675
R1510 VP.n31 VP.n30 24.4675
R1511 VP.n33 VP.n31 24.4675
R1512 VP.n37 VP.n19 24.4675
R1513 VP.n38 VP.n37 24.4675
R1514 VP.n26 VP.n25 24.4675
R1515 VP.n26 VP.n21 24.4675
R1516 VP.n55 VP.n12 21.0421
R1517 VP.n94 VP.n0 21.0421
R1518 VP.n52 VP.n13 21.0421
R1519 VP.n67 VP.n66 16.6381
R1520 VP.n86 VP.n85 16.6381
R1521 VP.n44 VP.n43 16.6381
R1522 VP.n25 VP.n24 16.6381
R1523 VP.n55 VP.t3 16.3291
R1524 VP.n66 VP.t6 16.3291
R1525 VP.n74 VP.t2 16.3291
R1526 VP.n86 VP.t8 16.3291
R1527 VP.n0 VP.t5 16.3291
R1528 VP.n13 VP.t4 16.3291
R1529 VP.n44 VP.t0 16.3291
R1530 VP.n32 VP.t9 16.3291
R1531 VP.n24 VP.t7 16.3291
R1532 VP.n75 VP.n74 12.234
R1533 VP.n74 VP.n6 12.234
R1534 VP.n33 VP.n32 12.234
R1535 VP.n32 VP.n19 12.234
R1536 VP.n66 VP.n65 7.82994
R1537 VP.n87 VP.n86 7.82994
R1538 VP.n45 VP.n44 7.82994
R1539 VP.n23 VP.n22 5.4582
R1540 VP.n54 VP.n53 0.354971
R1541 VP.n57 VP.n56 0.354971
R1542 VP.n96 VP.n95 0.354971
R1543 VP VP.n96 0.26696
R1544 VP.n27 VP.n22 0.189894
R1545 VP.n28 VP.n27 0.189894
R1546 VP.n29 VP.n28 0.189894
R1547 VP.n29 VP.n20 0.189894
R1548 VP.n34 VP.n20 0.189894
R1549 VP.n35 VP.n34 0.189894
R1550 VP.n36 VP.n35 0.189894
R1551 VP.n36 VP.n18 0.189894
R1552 VP.n40 VP.n18 0.189894
R1553 VP.n41 VP.n40 0.189894
R1554 VP.n42 VP.n41 0.189894
R1555 VP.n42 VP.n16 0.189894
R1556 VP.n47 VP.n16 0.189894
R1557 VP.n48 VP.n47 0.189894
R1558 VP.n49 VP.n48 0.189894
R1559 VP.n49 VP.n14 0.189894
R1560 VP.n53 VP.n14 0.189894
R1561 VP.n58 VP.n57 0.189894
R1562 VP.n58 VP.n11 0.189894
R1563 VP.n62 VP.n11 0.189894
R1564 VP.n63 VP.n62 0.189894
R1565 VP.n64 VP.n63 0.189894
R1566 VP.n64 VP.n9 0.189894
R1567 VP.n69 VP.n9 0.189894
R1568 VP.n70 VP.n69 0.189894
R1569 VP.n71 VP.n70 0.189894
R1570 VP.n71 VP.n7 0.189894
R1571 VP.n76 VP.n7 0.189894
R1572 VP.n77 VP.n76 0.189894
R1573 VP.n78 VP.n77 0.189894
R1574 VP.n78 VP.n5 0.189894
R1575 VP.n82 VP.n5 0.189894
R1576 VP.n83 VP.n82 0.189894
R1577 VP.n84 VP.n83 0.189894
R1578 VP.n84 VP.n3 0.189894
R1579 VP.n89 VP.n3 0.189894
R1580 VP.n90 VP.n89 0.189894
R1581 VP.n91 VP.n90 0.189894
R1582 VP.n91 VP.n1 0.189894
R1583 VP.n95 VP.n1 0.189894
R1584 VDD1.n2 VDD1.n0 289.615
R1585 VDD1.n11 VDD1.n9 289.615
R1586 VDD1.n3 VDD1.n2 185
R1587 VDD1.n12 VDD1.n11 185
R1588 VDD1.t8 VDD1.n1 164.876
R1589 VDD1.t5 VDD1.n10 164.876
R1590 VDD1.n19 VDD1.n18 105.111
R1591 VDD1.n21 VDD1.n20 103.168
R1592 VDD1.n8 VDD1.n7 103.168
R1593 VDD1.n17 VDD1.n16 103.168
R1594 VDD1.n8 VDD1.n6 55.2128
R1595 VDD1.n17 VDD1.n15 55.2128
R1596 VDD1.n2 VDD1.t8 52.3082
R1597 VDD1.n11 VDD1.t5 52.3082
R1598 VDD1.n21 VDD1.n19 39.8953
R1599 VDD1.n3 VDD1.n1 14.7318
R1600 VDD1.n12 VDD1.n10 14.7318
R1601 VDD1.n4 VDD1.n0 12.8005
R1602 VDD1.n13 VDD1.n9 12.8005
R1603 VDD1.n20 VDD1.t2 10.5887
R1604 VDD1.n20 VDD1.t4 10.5887
R1605 VDD1.n7 VDD1.t7 10.5887
R1606 VDD1.n7 VDD1.t3 10.5887
R1607 VDD1.n18 VDD1.t9 10.5887
R1608 VDD1.n18 VDD1.t6 10.5887
R1609 VDD1.n16 VDD1.t0 10.5887
R1610 VDD1.n16 VDD1.t1 10.5887
R1611 VDD1.n6 VDD1.n5 9.45567
R1612 VDD1.n15 VDD1.n14 9.45567
R1613 VDD1.n5 VDD1.n4 9.3005
R1614 VDD1.n14 VDD1.n13 9.3005
R1615 VDD1.n5 VDD1.n1 5.62509
R1616 VDD1.n14 VDD1.n10 5.62509
R1617 VDD1 VDD1.n21 1.94016
R1618 VDD1.n6 VDD1.n0 1.16414
R1619 VDD1.n15 VDD1.n9 1.16414
R1620 VDD1 VDD1.n8 0.724638
R1621 VDD1.n19 VDD1.n17 0.611102
R1622 VDD1.n4 VDD1.n3 0.388379
R1623 VDD1.n13 VDD1.n12 0.388379
R1624 VTAIL.n40 VTAIL.n38 289.615
R1625 VTAIL.n4 VTAIL.n2 289.615
R1626 VTAIL.n32 VTAIL.n30 289.615
R1627 VTAIL.n20 VTAIL.n18 289.615
R1628 VTAIL.n41 VTAIL.n40 185
R1629 VTAIL.n5 VTAIL.n4 185
R1630 VTAIL.n33 VTAIL.n32 185
R1631 VTAIL.n21 VTAIL.n20 185
R1632 VTAIL.t5 VTAIL.n39 164.876
R1633 VTAIL.t14 VTAIL.n3 164.876
R1634 VTAIL.t15 VTAIL.n31 164.876
R1635 VTAIL.t8 VTAIL.n19 164.876
R1636 VTAIL.n29 VTAIL.n28 86.4898
R1637 VTAIL.n27 VTAIL.n26 86.4898
R1638 VTAIL.n17 VTAIL.n16 86.4898
R1639 VTAIL.n15 VTAIL.n14 86.4898
R1640 VTAIL.n47 VTAIL.n46 86.4897
R1641 VTAIL.n1 VTAIL.n0 86.4897
R1642 VTAIL.n11 VTAIL.n10 86.4897
R1643 VTAIL.n13 VTAIL.n12 86.4897
R1644 VTAIL.n40 VTAIL.t5 52.3082
R1645 VTAIL.n4 VTAIL.t14 52.3082
R1646 VTAIL.n32 VTAIL.t15 52.3082
R1647 VTAIL.n20 VTAIL.t8 52.3082
R1648 VTAIL.n45 VTAIL.n44 35.8702
R1649 VTAIL.n9 VTAIL.n8 35.8702
R1650 VTAIL.n37 VTAIL.n36 35.8702
R1651 VTAIL.n25 VTAIL.n24 35.8702
R1652 VTAIL.n15 VTAIL.n13 19.3065
R1653 VTAIL.n45 VTAIL.n37 16.6427
R1654 VTAIL.n41 VTAIL.n39 14.7318
R1655 VTAIL.n5 VTAIL.n3 14.7318
R1656 VTAIL.n33 VTAIL.n31 14.7318
R1657 VTAIL.n21 VTAIL.n19 14.7318
R1658 VTAIL.n42 VTAIL.n38 12.8005
R1659 VTAIL.n6 VTAIL.n2 12.8005
R1660 VTAIL.n34 VTAIL.n30 12.8005
R1661 VTAIL.n22 VTAIL.n18 12.8005
R1662 VTAIL.n46 VTAIL.t2 10.5887
R1663 VTAIL.n46 VTAIL.t6 10.5887
R1664 VTAIL.n0 VTAIL.t0 10.5887
R1665 VTAIL.n0 VTAIL.t4 10.5887
R1666 VTAIL.n10 VTAIL.t17 10.5887
R1667 VTAIL.n10 VTAIL.t11 10.5887
R1668 VTAIL.n12 VTAIL.t16 10.5887
R1669 VTAIL.n12 VTAIL.t13 10.5887
R1670 VTAIL.n28 VTAIL.t10 10.5887
R1671 VTAIL.n28 VTAIL.t19 10.5887
R1672 VTAIL.n26 VTAIL.t18 10.5887
R1673 VTAIL.n26 VTAIL.t12 10.5887
R1674 VTAIL.n16 VTAIL.t7 10.5887
R1675 VTAIL.n16 VTAIL.t1 10.5887
R1676 VTAIL.n14 VTAIL.t9 10.5887
R1677 VTAIL.n14 VTAIL.t3 10.5887
R1678 VTAIL.n44 VTAIL.n43 9.45567
R1679 VTAIL.n8 VTAIL.n7 9.45567
R1680 VTAIL.n36 VTAIL.n35 9.45567
R1681 VTAIL.n24 VTAIL.n23 9.45567
R1682 VTAIL.n43 VTAIL.n42 9.3005
R1683 VTAIL.n7 VTAIL.n6 9.3005
R1684 VTAIL.n35 VTAIL.n34 9.3005
R1685 VTAIL.n23 VTAIL.n22 9.3005
R1686 VTAIL.n43 VTAIL.n39 5.62509
R1687 VTAIL.n7 VTAIL.n3 5.62509
R1688 VTAIL.n35 VTAIL.n31 5.62509
R1689 VTAIL.n23 VTAIL.n19 5.62509
R1690 VTAIL.n17 VTAIL.n15 2.66429
R1691 VTAIL.n25 VTAIL.n17 2.66429
R1692 VTAIL.n29 VTAIL.n27 2.66429
R1693 VTAIL.n37 VTAIL.n29 2.66429
R1694 VTAIL.n13 VTAIL.n11 2.66429
R1695 VTAIL.n11 VTAIL.n9 2.66429
R1696 VTAIL.n47 VTAIL.n45 2.66429
R1697 VTAIL VTAIL.n1 2.05653
R1698 VTAIL.n27 VTAIL.n25 1.80222
R1699 VTAIL.n9 VTAIL.n1 1.80222
R1700 VTAIL.n44 VTAIL.n38 1.16414
R1701 VTAIL.n8 VTAIL.n2 1.16414
R1702 VTAIL.n36 VTAIL.n30 1.16414
R1703 VTAIL.n24 VTAIL.n18 1.16414
R1704 VTAIL VTAIL.n47 0.608259
R1705 VTAIL.n42 VTAIL.n41 0.388379
R1706 VTAIL.n6 VTAIL.n5 0.388379
R1707 VTAIL.n34 VTAIL.n33 0.388379
R1708 VTAIL.n22 VTAIL.n21 0.388379
R1709 VN.n82 VN.n81 161.3
R1710 VN.n80 VN.n43 161.3
R1711 VN.n79 VN.n78 161.3
R1712 VN.n77 VN.n44 161.3
R1713 VN.n76 VN.n75 161.3
R1714 VN.n74 VN.n45 161.3
R1715 VN.n72 VN.n71 161.3
R1716 VN.n70 VN.n46 161.3
R1717 VN.n69 VN.n68 161.3
R1718 VN.n67 VN.n47 161.3
R1719 VN.n66 VN.n65 161.3
R1720 VN.n64 VN.n48 161.3
R1721 VN.n63 VN.n62 161.3
R1722 VN.n61 VN.n49 161.3
R1723 VN.n60 VN.n59 161.3
R1724 VN.n58 VN.n51 161.3
R1725 VN.n57 VN.n56 161.3
R1726 VN.n55 VN.n52 161.3
R1727 VN.n40 VN.n39 161.3
R1728 VN.n38 VN.n1 161.3
R1729 VN.n37 VN.n36 161.3
R1730 VN.n35 VN.n2 161.3
R1731 VN.n34 VN.n33 161.3
R1732 VN.n32 VN.n3 161.3
R1733 VN.n30 VN.n29 161.3
R1734 VN.n28 VN.n4 161.3
R1735 VN.n27 VN.n26 161.3
R1736 VN.n25 VN.n5 161.3
R1737 VN.n24 VN.n23 161.3
R1738 VN.n22 VN.n6 161.3
R1739 VN.n21 VN.n20 161.3
R1740 VN.n18 VN.n7 161.3
R1741 VN.n17 VN.n16 161.3
R1742 VN.n15 VN.n8 161.3
R1743 VN.n14 VN.n13 161.3
R1744 VN.n12 VN.n9 161.3
R1745 VN.n41 VN.n0 69.0258
R1746 VN.n83 VN.n42 69.0258
R1747 VN.n11 VN.n10 56.938
R1748 VN.n54 VN.n53 56.938
R1749 VN.n17 VN.n8 56.5193
R1750 VN.n26 VN.n25 56.5193
R1751 VN.n60 VN.n51 56.5193
R1752 VN.n68 VN.n67 56.5193
R1753 VN.n37 VN.n2 51.663
R1754 VN.n79 VN.n44 51.663
R1755 VN.n53 VN.t4 48.2127
R1756 VN.n10 VN.t2 48.2127
R1757 VN VN.n83 46.5548
R1758 VN.n38 VN.n37 29.3238
R1759 VN.n80 VN.n79 29.3238
R1760 VN.n13 VN.n12 24.4675
R1761 VN.n13 VN.n8 24.4675
R1762 VN.n18 VN.n17 24.4675
R1763 VN.n20 VN.n18 24.4675
R1764 VN.n24 VN.n6 24.4675
R1765 VN.n25 VN.n24 24.4675
R1766 VN.n26 VN.n4 24.4675
R1767 VN.n30 VN.n4 24.4675
R1768 VN.n33 VN.n32 24.4675
R1769 VN.n33 VN.n2 24.4675
R1770 VN.n39 VN.n38 24.4675
R1771 VN.n56 VN.n51 24.4675
R1772 VN.n56 VN.n55 24.4675
R1773 VN.n67 VN.n66 24.4675
R1774 VN.n66 VN.n48 24.4675
R1775 VN.n62 VN.n61 24.4675
R1776 VN.n61 VN.n60 24.4675
R1777 VN.n75 VN.n44 24.4675
R1778 VN.n75 VN.n74 24.4675
R1779 VN.n72 VN.n46 24.4675
R1780 VN.n68 VN.n46 24.4675
R1781 VN.n81 VN.n80 24.4675
R1782 VN.n39 VN.n0 21.0421
R1783 VN.n81 VN.n42 21.0421
R1784 VN.n12 VN.n11 16.6381
R1785 VN.n31 VN.n30 16.6381
R1786 VN.n55 VN.n54 16.6381
R1787 VN.n73 VN.n72 16.6381
R1788 VN.n11 VN.t6 16.3291
R1789 VN.n19 VN.t8 16.3291
R1790 VN.n31 VN.t5 16.3291
R1791 VN.n0 VN.t3 16.3291
R1792 VN.n54 VN.t9 16.3291
R1793 VN.n50 VN.t1 16.3291
R1794 VN.n73 VN.t7 16.3291
R1795 VN.n42 VN.t0 16.3291
R1796 VN.n20 VN.n19 12.234
R1797 VN.n19 VN.n6 12.234
R1798 VN.n50 VN.n48 12.234
R1799 VN.n62 VN.n50 12.234
R1800 VN.n32 VN.n31 7.82994
R1801 VN.n74 VN.n73 7.82994
R1802 VN.n53 VN.n52 5.45824
R1803 VN.n10 VN.n9 5.45823
R1804 VN.n83 VN.n82 0.354971
R1805 VN.n41 VN.n40 0.354971
R1806 VN VN.n41 0.26696
R1807 VN.n82 VN.n43 0.189894
R1808 VN.n78 VN.n43 0.189894
R1809 VN.n78 VN.n77 0.189894
R1810 VN.n77 VN.n76 0.189894
R1811 VN.n76 VN.n45 0.189894
R1812 VN.n71 VN.n45 0.189894
R1813 VN.n71 VN.n70 0.189894
R1814 VN.n70 VN.n69 0.189894
R1815 VN.n69 VN.n47 0.189894
R1816 VN.n65 VN.n47 0.189894
R1817 VN.n65 VN.n64 0.189894
R1818 VN.n64 VN.n63 0.189894
R1819 VN.n63 VN.n49 0.189894
R1820 VN.n59 VN.n49 0.189894
R1821 VN.n59 VN.n58 0.189894
R1822 VN.n58 VN.n57 0.189894
R1823 VN.n57 VN.n52 0.189894
R1824 VN.n14 VN.n9 0.189894
R1825 VN.n15 VN.n14 0.189894
R1826 VN.n16 VN.n15 0.189894
R1827 VN.n16 VN.n7 0.189894
R1828 VN.n21 VN.n7 0.189894
R1829 VN.n22 VN.n21 0.189894
R1830 VN.n23 VN.n22 0.189894
R1831 VN.n23 VN.n5 0.189894
R1832 VN.n27 VN.n5 0.189894
R1833 VN.n28 VN.n27 0.189894
R1834 VN.n29 VN.n28 0.189894
R1835 VN.n29 VN.n3 0.189894
R1836 VN.n34 VN.n3 0.189894
R1837 VN.n35 VN.n34 0.189894
R1838 VN.n36 VN.n35 0.189894
R1839 VN.n36 VN.n1 0.189894
R1840 VN.n40 VN.n1 0.189894
R1841 VDD2.n13 VDD2.n11 289.615
R1842 VDD2.n2 VDD2.n0 289.615
R1843 VDD2.n14 VDD2.n13 185
R1844 VDD2.n3 VDD2.n2 185
R1845 VDD2.t9 VDD2.n12 164.876
R1846 VDD2.t7 VDD2.n1 164.876
R1847 VDD2.n10 VDD2.n9 105.111
R1848 VDD2 VDD2.n21 105.109
R1849 VDD2.n20 VDD2.n19 103.168
R1850 VDD2.n8 VDD2.n7 103.168
R1851 VDD2.n8 VDD2.n6 55.2128
R1852 VDD2.n18 VDD2.n17 52.549
R1853 VDD2.n13 VDD2.t9 52.3082
R1854 VDD2.n2 VDD2.t7 52.3082
R1855 VDD2.n18 VDD2.n10 37.9804
R1856 VDD2.n14 VDD2.n12 14.7318
R1857 VDD2.n3 VDD2.n1 14.7318
R1858 VDD2.n15 VDD2.n11 12.8005
R1859 VDD2.n4 VDD2.n0 12.8005
R1860 VDD2.n21 VDD2.t0 10.5887
R1861 VDD2.n21 VDD2.t5 10.5887
R1862 VDD2.n19 VDD2.t2 10.5887
R1863 VDD2.n19 VDD2.t8 10.5887
R1864 VDD2.n9 VDD2.t4 10.5887
R1865 VDD2.n9 VDD2.t6 10.5887
R1866 VDD2.n7 VDD2.t3 10.5887
R1867 VDD2.n7 VDD2.t1 10.5887
R1868 VDD2.n17 VDD2.n16 9.45567
R1869 VDD2.n6 VDD2.n5 9.45567
R1870 VDD2.n16 VDD2.n15 9.3005
R1871 VDD2.n5 VDD2.n4 9.3005
R1872 VDD2.n16 VDD2.n12 5.62509
R1873 VDD2.n5 VDD2.n1 5.62509
R1874 VDD2.n20 VDD2.n18 2.66429
R1875 VDD2.n17 VDD2.n11 1.16414
R1876 VDD2.n6 VDD2.n0 1.16414
R1877 VDD2 VDD2.n20 0.724638
R1878 VDD2.n10 VDD2.n8 0.611102
R1879 VDD2.n15 VDD2.n14 0.388379
R1880 VDD2.n4 VDD2.n3 0.388379
C0 VTAIL VDD1 5.89437f
C1 VDD2 VDD1 2.27792f
C2 VTAIL VP 3.65911f
C3 VTAIL VN 3.64498f
C4 VDD2 VP 0.611399f
C5 VDD2 VN 2.12513f
C6 VP VDD1 2.57203f
C7 VN VDD1 0.160425f
C8 VN VP 6.77157f
C9 VDD2 VTAIL 5.94878f
C10 VDD2 B 5.739356f
C11 VDD1 B 5.61038f
C12 VTAIL B 3.749026f
C13 VN B 18.12801f
C14 VP B 16.49141f
C15 VDD2.n0 B 0.04082f
C16 VDD2.n1 B 0.095702f
C17 VDD2.t7 B 0.067825f
C18 VDD2.n2 B 0.070591f
C19 VDD2.n3 B 0.019698f
C20 VDD2.n4 B 0.015989f
C21 VDD2.n5 B 0.188335f
C22 VDD2.n6 B 0.08062f
C23 VDD2.t3 B 0.04397f
C24 VDD2.t1 B 0.04397f
C25 VDD2.n7 B 0.282298f
C26 VDD2.n8 B 0.82869f
C27 VDD2.t4 B 0.04397f
C28 VDD2.t6 B 0.04397f
C29 VDD2.n9 B 0.294602f
C30 VDD2.n10 B 2.807f
C31 VDD2.n11 B 0.04082f
C32 VDD2.n12 B 0.095702f
C33 VDD2.t9 B 0.067825f
C34 VDD2.n13 B 0.070591f
C35 VDD2.n14 B 0.019698f
C36 VDD2.n15 B 0.015989f
C37 VDD2.n16 B 0.188335f
C38 VDD2.n17 B 0.065321f
C39 VDD2.n18 B 2.57002f
C40 VDD2.t2 B 0.04397f
C41 VDD2.t8 B 0.04397f
C42 VDD2.n19 B 0.282299f
C43 VDD2.n20 B 0.536626f
C44 VDD2.t0 B 0.04397f
C45 VDD2.t5 B 0.04397f
C46 VDD2.n21 B 0.294574f
C47 VN.t3 B 0.346187f
C48 VN.n0 B 0.27614f
C49 VN.n1 B 0.029126f
C50 VN.n2 B 0.052591f
C51 VN.n3 B 0.029126f
C52 VN.t5 B 0.346187f
C53 VN.n4 B 0.054284f
C54 VN.n5 B 0.029126f
C55 VN.n6 B 0.040883f
C56 VN.n7 B 0.029126f
C57 VN.n8 B 0.038869f
C58 VN.n9 B 0.306292f
C59 VN.t6 B 0.346187f
C60 VN.t2 B 0.579935f
C61 VN.n10 B 0.253561f
C62 VN.n11 B 0.260704f
C63 VN.n12 B 0.045707f
C64 VN.n13 B 0.054284f
C65 VN.n14 B 0.029126f
C66 VN.n15 B 0.029126f
C67 VN.n16 B 0.029126f
C68 VN.n17 B 0.046174f
C69 VN.n18 B 0.054284f
C70 VN.t8 B 0.346187f
C71 VN.n19 B 0.167227f
C72 VN.n20 B 0.040883f
C73 VN.n21 B 0.029126f
C74 VN.n22 B 0.029126f
C75 VN.n23 B 0.029126f
C76 VN.n24 B 0.054284f
C77 VN.n25 B 0.046174f
C78 VN.n26 B 0.038869f
C79 VN.n27 B 0.029126f
C80 VN.n28 B 0.029126f
C81 VN.n29 B 0.029126f
C82 VN.n30 B 0.045707f
C83 VN.n31 B 0.167227f
C84 VN.n32 B 0.03606f
C85 VN.n33 B 0.054284f
C86 VN.n34 B 0.029126f
C87 VN.n35 B 0.029126f
C88 VN.n36 B 0.029126f
C89 VN.n37 B 0.028902f
C90 VN.n38 B 0.057834f
C91 VN.n39 B 0.050532f
C92 VN.n40 B 0.047009f
C93 VN.n41 B 0.057035f
C94 VN.t0 B 0.346187f
C95 VN.n42 B 0.27614f
C96 VN.n43 B 0.029126f
C97 VN.n44 B 0.052591f
C98 VN.n45 B 0.029126f
C99 VN.t7 B 0.346187f
C100 VN.n46 B 0.054284f
C101 VN.n47 B 0.029126f
C102 VN.n48 B 0.040883f
C103 VN.n49 B 0.029126f
C104 VN.t1 B 0.346187f
C105 VN.n50 B 0.167227f
C106 VN.n51 B 0.038869f
C107 VN.n52 B 0.306292f
C108 VN.t9 B 0.346187f
C109 VN.t4 B 0.579935f
C110 VN.n53 B 0.253561f
C111 VN.n54 B 0.260704f
C112 VN.n55 B 0.045707f
C113 VN.n56 B 0.054284f
C114 VN.n57 B 0.029126f
C115 VN.n58 B 0.029126f
C116 VN.n59 B 0.029126f
C117 VN.n60 B 0.046174f
C118 VN.n61 B 0.054284f
C119 VN.n62 B 0.040883f
C120 VN.n63 B 0.029126f
C121 VN.n64 B 0.029126f
C122 VN.n65 B 0.029126f
C123 VN.n66 B 0.054284f
C124 VN.n67 B 0.046174f
C125 VN.n68 B 0.038869f
C126 VN.n69 B 0.029126f
C127 VN.n70 B 0.029126f
C128 VN.n71 B 0.029126f
C129 VN.n72 B 0.045707f
C130 VN.n73 B 0.167227f
C131 VN.n74 B 0.03606f
C132 VN.n75 B 0.054284f
C133 VN.n76 B 0.029126f
C134 VN.n77 B 0.029126f
C135 VN.n78 B 0.029126f
C136 VN.n79 B 0.028902f
C137 VN.n80 B 0.057834f
C138 VN.n81 B 0.050532f
C139 VN.n82 B 0.047009f
C140 VN.n83 B 1.48103f
C141 VTAIL.t0 B 0.055355f
C142 VTAIL.t4 B 0.055355f
C143 VTAIL.n0 B 0.305345f
C144 VTAIL.n1 B 0.731405f
C145 VTAIL.n2 B 0.051389f
C146 VTAIL.n3 B 0.12048f
C147 VTAIL.t14 B 0.085385f
C148 VTAIL.n4 B 0.088868f
C149 VTAIL.n5 B 0.024798f
C150 VTAIL.n6 B 0.020129f
C151 VTAIL.n7 B 0.237098f
C152 VTAIL.n8 B 0.056436f
C153 VTAIL.n9 B 0.576492f
C154 VTAIL.t17 B 0.055355f
C155 VTAIL.t11 B 0.055355f
C156 VTAIL.n10 B 0.305345f
C157 VTAIL.n11 B 0.908817f
C158 VTAIL.t16 B 0.055355f
C159 VTAIL.t13 B 0.055355f
C160 VTAIL.n12 B 0.305345f
C161 VTAIL.n13 B 1.93376f
C162 VTAIL.t9 B 0.055355f
C163 VTAIL.t3 B 0.055355f
C164 VTAIL.n14 B 0.305347f
C165 VTAIL.n15 B 1.93376f
C166 VTAIL.t7 B 0.055355f
C167 VTAIL.t1 B 0.055355f
C168 VTAIL.n16 B 0.305347f
C169 VTAIL.n17 B 0.908815f
C170 VTAIL.n18 B 0.051389f
C171 VTAIL.n19 B 0.12048f
C172 VTAIL.t8 B 0.085385f
C173 VTAIL.n20 B 0.088868f
C174 VTAIL.n21 B 0.024798f
C175 VTAIL.n22 B 0.020129f
C176 VTAIL.n23 B 0.237098f
C177 VTAIL.n24 B 0.056436f
C178 VTAIL.n25 B 0.576492f
C179 VTAIL.t18 B 0.055355f
C180 VTAIL.t12 B 0.055355f
C181 VTAIL.n26 B 0.305347f
C182 VTAIL.n27 B 0.804761f
C183 VTAIL.t10 B 0.055355f
C184 VTAIL.t19 B 0.055355f
C185 VTAIL.n28 B 0.305347f
C186 VTAIL.n29 B 0.908815f
C187 VTAIL.n30 B 0.051389f
C188 VTAIL.n31 B 0.12048f
C189 VTAIL.t15 B 0.085385f
C190 VTAIL.n32 B 0.088868f
C191 VTAIL.n33 B 0.024798f
C192 VTAIL.n34 B 0.020129f
C193 VTAIL.n35 B 0.237098f
C194 VTAIL.n36 B 0.056436f
C195 VTAIL.n37 B 1.38397f
C196 VTAIL.n38 B 0.051389f
C197 VTAIL.n39 B 0.12048f
C198 VTAIL.t5 B 0.085385f
C199 VTAIL.n40 B 0.088868f
C200 VTAIL.n41 B 0.024798f
C201 VTAIL.n42 B 0.020129f
C202 VTAIL.n43 B 0.237098f
C203 VTAIL.n44 B 0.056436f
C204 VTAIL.n45 B 1.38397f
C205 VTAIL.t2 B 0.055355f
C206 VTAIL.t6 B 0.055355f
C207 VTAIL.n46 B 0.305345f
C208 VTAIL.n47 B 0.660649f
C209 VDD1.n0 B 0.042349f
C210 VDD1.n1 B 0.099288f
C211 VDD1.t8 B 0.070366f
C212 VDD1.n2 B 0.073237f
C213 VDD1.n3 B 0.020436f
C214 VDD1.n4 B 0.016588f
C215 VDD1.n5 B 0.195393f
C216 VDD1.n6 B 0.083642f
C217 VDD1.t7 B 0.045618f
C218 VDD1.t3 B 0.045618f
C219 VDD1.n7 B 0.292878f
C220 VDD1.n8 B 0.869864f
C221 VDD1.n9 B 0.042349f
C222 VDD1.n10 B 0.099288f
C223 VDD1.t5 B 0.070366f
C224 VDD1.n11 B 0.073237f
C225 VDD1.n12 B 0.020436f
C226 VDD1.n13 B 0.016588f
C227 VDD1.n14 B 0.195393f
C228 VDD1.n15 B 0.083642f
C229 VDD1.t0 B 0.045618f
C230 VDD1.t1 B 0.045618f
C231 VDD1.n16 B 0.292877f
C232 VDD1.n17 B 0.859744f
C233 VDD1.t9 B 0.045618f
C234 VDD1.t6 B 0.045618f
C235 VDD1.n18 B 0.305642f
C236 VDD1.n19 B 3.06012f
C237 VDD1.t2 B 0.045618f
C238 VDD1.t4 B 0.045618f
C239 VDD1.n20 B 0.292878f
C240 VDD1.n21 B 2.99349f
C241 VP.t5 B 0.363996f
C242 VP.n0 B 0.290346f
C243 VP.n1 B 0.030624f
C244 VP.n2 B 0.055296f
C245 VP.n3 B 0.030624f
C246 VP.t8 B 0.363996f
C247 VP.n4 B 0.057076f
C248 VP.n5 B 0.030624f
C249 VP.n6 B 0.042987f
C250 VP.n7 B 0.030624f
C251 VP.n8 B 0.040869f
C252 VP.n9 B 0.030624f
C253 VP.t6 B 0.363996f
C254 VP.n10 B 0.057076f
C255 VP.n11 B 0.030624f
C256 VP.n12 B 0.053131f
C257 VP.t4 B 0.363996f
C258 VP.n13 B 0.290346f
C259 VP.n14 B 0.030624f
C260 VP.n15 B 0.055296f
C261 VP.n16 B 0.030624f
C262 VP.t0 B 0.363996f
C263 VP.n17 B 0.057076f
C264 VP.n18 B 0.030624f
C265 VP.n19 B 0.042987f
C266 VP.n20 B 0.030624f
C267 VP.n21 B 0.040869f
C268 VP.n22 B 0.322049f
C269 VP.t7 B 0.363996f
C270 VP.t1 B 0.609768f
C271 VP.n23 B 0.266606f
C272 VP.n24 B 0.274115f
C273 VP.n25 B 0.048059f
C274 VP.n26 B 0.057076f
C275 VP.n27 B 0.030624f
C276 VP.n28 B 0.030624f
C277 VP.n29 B 0.030624f
C278 VP.n30 B 0.048549f
C279 VP.n31 B 0.057076f
C280 VP.t9 B 0.363996f
C281 VP.n32 B 0.17583f
C282 VP.n33 B 0.042987f
C283 VP.n34 B 0.030624f
C284 VP.n35 B 0.030624f
C285 VP.n36 B 0.030624f
C286 VP.n37 B 0.057076f
C287 VP.n38 B 0.048549f
C288 VP.n39 B 0.040869f
C289 VP.n40 B 0.030624f
C290 VP.n41 B 0.030624f
C291 VP.n42 B 0.030624f
C292 VP.n43 B 0.048059f
C293 VP.n44 B 0.17583f
C294 VP.n45 B 0.037915f
C295 VP.n46 B 0.057076f
C296 VP.n47 B 0.030624f
C297 VP.n48 B 0.030624f
C298 VP.n49 B 0.030624f
C299 VP.n50 B 0.030388f
C300 VP.n51 B 0.06081f
C301 VP.n52 B 0.053131f
C302 VP.n53 B 0.049427f
C303 VP.n54 B 1.54434f
C304 VP.t3 B 0.363996f
C305 VP.n55 B 0.290346f
C306 VP.n56 B 1.56807f
C307 VP.n57 B 0.049427f
C308 VP.n58 B 0.030624f
C309 VP.n59 B 0.06081f
C310 VP.n60 B 0.030388f
C311 VP.n61 B 0.055296f
C312 VP.n62 B 0.030624f
C313 VP.n63 B 0.030624f
C314 VP.n64 B 0.030624f
C315 VP.n65 B 0.037915f
C316 VP.n66 B 0.17583f
C317 VP.n67 B 0.048059f
C318 VP.n68 B 0.057076f
C319 VP.n69 B 0.030624f
C320 VP.n70 B 0.030624f
C321 VP.n71 B 0.030624f
C322 VP.n72 B 0.048549f
C323 VP.n73 B 0.057076f
C324 VP.t2 B 0.363996f
C325 VP.n74 B 0.17583f
C326 VP.n75 B 0.042987f
C327 VP.n76 B 0.030624f
C328 VP.n77 B 0.030624f
C329 VP.n78 B 0.030624f
C330 VP.n79 B 0.057076f
C331 VP.n80 B 0.048549f
C332 VP.n81 B 0.040869f
C333 VP.n82 B 0.030624f
C334 VP.n83 B 0.030624f
C335 VP.n84 B 0.030624f
C336 VP.n85 B 0.048059f
C337 VP.n86 B 0.17583f
C338 VP.n87 B 0.037915f
C339 VP.n88 B 0.057076f
C340 VP.n89 B 0.030624f
C341 VP.n90 B 0.030624f
C342 VP.n91 B 0.030624f
C343 VP.n92 B 0.030388f
C344 VP.n93 B 0.06081f
C345 VP.n94 B 0.053131f
C346 VP.n95 B 0.049427f
C347 VP.n96 B 0.059969f
.ends

