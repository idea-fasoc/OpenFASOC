* NGSPICE file created from diff_pair_sample_0731.ext - technology: sky130A

.subckt diff_pair_sample_0731 VTAIL VN VP B VDD2 VDD1
X0 B.t20 B.t18 B.t19 B.t12 sky130_fd_pr__nfet_01v8 ad=4.4655 pd=23.68 as=0 ps=0 w=11.45 l=0.49
X1 VTAIL.t17 VP.t0 VDD1.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=1.88925 pd=11.78 as=1.88925 ps=11.78 w=11.45 l=0.49
X2 VDD1.t7 VP.t1 VTAIL.t16 B.t3 sky130_fd_pr__nfet_01v8 ad=1.88925 pd=11.78 as=1.88925 ps=11.78 w=11.45 l=0.49
X3 VDD2.t9 VN.t0 VTAIL.t3 B.t2 sky130_fd_pr__nfet_01v8 ad=1.88925 pd=11.78 as=1.88925 ps=11.78 w=11.45 l=0.49
X4 B.t17 B.t15 B.t16 B.t8 sky130_fd_pr__nfet_01v8 ad=4.4655 pd=23.68 as=0 ps=0 w=11.45 l=0.49
X5 B.t14 B.t11 B.t13 B.t12 sky130_fd_pr__nfet_01v8 ad=4.4655 pd=23.68 as=0 ps=0 w=11.45 l=0.49
X6 B.t10 B.t7 B.t9 B.t8 sky130_fd_pr__nfet_01v8 ad=4.4655 pd=23.68 as=0 ps=0 w=11.45 l=0.49
X7 VTAIL.t2 VN.t1 VDD2.t8 B.t4 sky130_fd_pr__nfet_01v8 ad=1.88925 pd=11.78 as=1.88925 ps=11.78 w=11.45 l=0.49
X8 VDD1.t8 VP.t2 VTAIL.t15 B.t6 sky130_fd_pr__nfet_01v8 ad=1.88925 pd=11.78 as=4.4655 ps=23.68 w=11.45 l=0.49
X9 VDD2.t7 VN.t2 VTAIL.t6 B.t5 sky130_fd_pr__nfet_01v8 ad=4.4655 pd=23.68 as=1.88925 ps=11.78 w=11.45 l=0.49
X10 VDD2.t6 VN.t3 VTAIL.t1 B.t3 sky130_fd_pr__nfet_01v8 ad=1.88925 pd=11.78 as=1.88925 ps=11.78 w=11.45 l=0.49
X11 VDD2.t5 VN.t4 VTAIL.t4 B.t6 sky130_fd_pr__nfet_01v8 ad=1.88925 pd=11.78 as=4.4655 ps=23.68 w=11.45 l=0.49
X12 VDD2.t4 VN.t5 VTAIL.t5 B.t0 sky130_fd_pr__nfet_01v8 ad=4.4655 pd=23.68 as=1.88925 ps=11.78 w=11.45 l=0.49
X13 VTAIL.t14 VP.t3 VDD1.t5 B.t22 sky130_fd_pr__nfet_01v8 ad=1.88925 pd=11.78 as=1.88925 ps=11.78 w=11.45 l=0.49
X14 VTAIL.t18 VN.t6 VDD2.t3 B.t22 sky130_fd_pr__nfet_01v8 ad=1.88925 pd=11.78 as=1.88925 ps=11.78 w=11.45 l=0.49
X15 VDD2.t2 VN.t7 VTAIL.t7 B.t21 sky130_fd_pr__nfet_01v8 ad=1.88925 pd=11.78 as=4.4655 ps=23.68 w=11.45 l=0.49
X16 VTAIL.t0 VN.t8 VDD2.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=1.88925 pd=11.78 as=1.88925 ps=11.78 w=11.45 l=0.49
X17 VDD1.t4 VP.t4 VTAIL.t13 B.t21 sky130_fd_pr__nfet_01v8 ad=1.88925 pd=11.78 as=4.4655 ps=23.68 w=11.45 l=0.49
X18 VTAIL.t19 VN.t9 VDD2.t0 B.t23 sky130_fd_pr__nfet_01v8 ad=1.88925 pd=11.78 as=1.88925 ps=11.78 w=11.45 l=0.49
X19 VDD1.t3 VP.t5 VTAIL.t12 B.t2 sky130_fd_pr__nfet_01v8 ad=1.88925 pd=11.78 as=1.88925 ps=11.78 w=11.45 l=0.49
X20 VDD1.t9 VP.t6 VTAIL.t11 B.t5 sky130_fd_pr__nfet_01v8 ad=4.4655 pd=23.68 as=1.88925 ps=11.78 w=11.45 l=0.49
X21 VDD1.t6 VP.t7 VTAIL.t10 B.t0 sky130_fd_pr__nfet_01v8 ad=4.4655 pd=23.68 as=1.88925 ps=11.78 w=11.45 l=0.49
X22 VTAIL.t9 VP.t8 VDD1.t0 B.t4 sky130_fd_pr__nfet_01v8 ad=1.88925 pd=11.78 as=1.88925 ps=11.78 w=11.45 l=0.49
X23 VTAIL.t8 VP.t9 VDD1.t2 B.t23 sky130_fd_pr__nfet_01v8 ad=1.88925 pd=11.78 as=1.88925 ps=11.78 w=11.45 l=0.49
R0 B.n66 B.t7 769.808
R1 B.n72 B.t15 769.808
R2 B.n166 B.t18 769.808
R3 B.n158 B.t11 769.808
R4 B.n464 B.n463 585
R5 B.n466 B.n94 585
R6 B.n469 B.n468 585
R7 B.n470 B.n93 585
R8 B.n472 B.n471 585
R9 B.n474 B.n92 585
R10 B.n477 B.n476 585
R11 B.n478 B.n91 585
R12 B.n480 B.n479 585
R13 B.n482 B.n90 585
R14 B.n485 B.n484 585
R15 B.n486 B.n89 585
R16 B.n488 B.n487 585
R17 B.n490 B.n88 585
R18 B.n493 B.n492 585
R19 B.n494 B.n87 585
R20 B.n496 B.n495 585
R21 B.n498 B.n86 585
R22 B.n501 B.n500 585
R23 B.n502 B.n85 585
R24 B.n504 B.n503 585
R25 B.n506 B.n84 585
R26 B.n509 B.n508 585
R27 B.n510 B.n83 585
R28 B.n512 B.n511 585
R29 B.n514 B.n82 585
R30 B.n517 B.n516 585
R31 B.n518 B.n81 585
R32 B.n520 B.n519 585
R33 B.n522 B.n80 585
R34 B.n525 B.n524 585
R35 B.n526 B.n79 585
R36 B.n528 B.n527 585
R37 B.n530 B.n78 585
R38 B.n533 B.n532 585
R39 B.n534 B.n77 585
R40 B.n536 B.n535 585
R41 B.n538 B.n76 585
R42 B.n540 B.n539 585
R43 B.n542 B.n541 585
R44 B.n545 B.n544 585
R45 B.n546 B.n71 585
R46 B.n548 B.n547 585
R47 B.n550 B.n70 585
R48 B.n553 B.n552 585
R49 B.n554 B.n69 585
R50 B.n556 B.n555 585
R51 B.n558 B.n68 585
R52 B.n561 B.n560 585
R53 B.n562 B.n65 585
R54 B.n565 B.n564 585
R55 B.n567 B.n64 585
R56 B.n570 B.n569 585
R57 B.n571 B.n63 585
R58 B.n573 B.n572 585
R59 B.n575 B.n62 585
R60 B.n578 B.n577 585
R61 B.n579 B.n61 585
R62 B.n581 B.n580 585
R63 B.n583 B.n60 585
R64 B.n586 B.n585 585
R65 B.n587 B.n59 585
R66 B.n589 B.n588 585
R67 B.n591 B.n58 585
R68 B.n594 B.n593 585
R69 B.n595 B.n57 585
R70 B.n597 B.n596 585
R71 B.n599 B.n56 585
R72 B.n602 B.n601 585
R73 B.n603 B.n55 585
R74 B.n605 B.n604 585
R75 B.n607 B.n54 585
R76 B.n610 B.n609 585
R77 B.n611 B.n53 585
R78 B.n613 B.n612 585
R79 B.n615 B.n52 585
R80 B.n618 B.n617 585
R81 B.n619 B.n51 585
R82 B.n621 B.n620 585
R83 B.n623 B.n50 585
R84 B.n626 B.n625 585
R85 B.n627 B.n49 585
R86 B.n629 B.n628 585
R87 B.n631 B.n48 585
R88 B.n634 B.n633 585
R89 B.n635 B.n47 585
R90 B.n637 B.n636 585
R91 B.n639 B.n46 585
R92 B.n642 B.n641 585
R93 B.n643 B.n45 585
R94 B.n462 B.n43 585
R95 B.n646 B.n43 585
R96 B.n461 B.n42 585
R97 B.n647 B.n42 585
R98 B.n460 B.n41 585
R99 B.n648 B.n41 585
R100 B.n459 B.n458 585
R101 B.n458 B.n37 585
R102 B.n457 B.n36 585
R103 B.n654 B.n36 585
R104 B.n456 B.n35 585
R105 B.n655 B.n35 585
R106 B.n455 B.n34 585
R107 B.n656 B.n34 585
R108 B.n454 B.n453 585
R109 B.n453 B.n30 585
R110 B.n452 B.n29 585
R111 B.n662 B.n29 585
R112 B.n451 B.n28 585
R113 B.n663 B.n28 585
R114 B.n450 B.n27 585
R115 B.n664 B.n27 585
R116 B.n449 B.n448 585
R117 B.n448 B.n23 585
R118 B.n447 B.n22 585
R119 B.n670 B.n22 585
R120 B.n446 B.n21 585
R121 B.n671 B.n21 585
R122 B.n445 B.n20 585
R123 B.n672 B.n20 585
R124 B.n444 B.n443 585
R125 B.n443 B.n16 585
R126 B.n442 B.n15 585
R127 B.n678 B.n15 585
R128 B.n441 B.n14 585
R129 B.n679 B.n14 585
R130 B.n440 B.n13 585
R131 B.n680 B.n13 585
R132 B.n439 B.n438 585
R133 B.n438 B.n12 585
R134 B.n437 B.n436 585
R135 B.n437 B.n8 585
R136 B.n435 B.n7 585
R137 B.n687 B.n7 585
R138 B.n434 B.n6 585
R139 B.n688 B.n6 585
R140 B.n433 B.n5 585
R141 B.n689 B.n5 585
R142 B.n432 B.n431 585
R143 B.n431 B.n4 585
R144 B.n430 B.n95 585
R145 B.n430 B.n429 585
R146 B.n419 B.n96 585
R147 B.n422 B.n96 585
R148 B.n421 B.n420 585
R149 B.n423 B.n421 585
R150 B.n418 B.n100 585
R151 B.n104 B.n100 585
R152 B.n417 B.n416 585
R153 B.n416 B.n415 585
R154 B.n102 B.n101 585
R155 B.n103 B.n102 585
R156 B.n408 B.n407 585
R157 B.n409 B.n408 585
R158 B.n406 B.n109 585
R159 B.n109 B.n108 585
R160 B.n405 B.n404 585
R161 B.n404 B.n403 585
R162 B.n111 B.n110 585
R163 B.n112 B.n111 585
R164 B.n396 B.n395 585
R165 B.n397 B.n396 585
R166 B.n394 B.n117 585
R167 B.n117 B.n116 585
R168 B.n393 B.n392 585
R169 B.n392 B.n391 585
R170 B.n119 B.n118 585
R171 B.n120 B.n119 585
R172 B.n384 B.n383 585
R173 B.n385 B.n384 585
R174 B.n382 B.n125 585
R175 B.n125 B.n124 585
R176 B.n381 B.n380 585
R177 B.n380 B.n379 585
R178 B.n127 B.n126 585
R179 B.n128 B.n127 585
R180 B.n372 B.n371 585
R181 B.n373 B.n372 585
R182 B.n370 B.n133 585
R183 B.n133 B.n132 585
R184 B.n369 B.n368 585
R185 B.n368 B.n367 585
R186 B.n364 B.n137 585
R187 B.n363 B.n362 585
R188 B.n360 B.n138 585
R189 B.n360 B.n136 585
R190 B.n359 B.n358 585
R191 B.n357 B.n356 585
R192 B.n355 B.n140 585
R193 B.n353 B.n352 585
R194 B.n351 B.n141 585
R195 B.n350 B.n349 585
R196 B.n347 B.n142 585
R197 B.n345 B.n344 585
R198 B.n343 B.n143 585
R199 B.n342 B.n341 585
R200 B.n339 B.n144 585
R201 B.n337 B.n336 585
R202 B.n335 B.n145 585
R203 B.n334 B.n333 585
R204 B.n331 B.n146 585
R205 B.n329 B.n328 585
R206 B.n327 B.n147 585
R207 B.n326 B.n325 585
R208 B.n323 B.n148 585
R209 B.n321 B.n320 585
R210 B.n319 B.n149 585
R211 B.n318 B.n317 585
R212 B.n315 B.n150 585
R213 B.n313 B.n312 585
R214 B.n311 B.n151 585
R215 B.n310 B.n309 585
R216 B.n307 B.n152 585
R217 B.n305 B.n304 585
R218 B.n303 B.n153 585
R219 B.n302 B.n301 585
R220 B.n299 B.n154 585
R221 B.n297 B.n296 585
R222 B.n295 B.n155 585
R223 B.n294 B.n293 585
R224 B.n291 B.n156 585
R225 B.n289 B.n288 585
R226 B.n287 B.n157 585
R227 B.n285 B.n284 585
R228 B.n282 B.n160 585
R229 B.n280 B.n279 585
R230 B.n278 B.n161 585
R231 B.n277 B.n276 585
R232 B.n274 B.n162 585
R233 B.n272 B.n271 585
R234 B.n270 B.n163 585
R235 B.n269 B.n268 585
R236 B.n266 B.n164 585
R237 B.n264 B.n263 585
R238 B.n262 B.n165 585
R239 B.n261 B.n260 585
R240 B.n258 B.n169 585
R241 B.n256 B.n255 585
R242 B.n254 B.n170 585
R243 B.n253 B.n252 585
R244 B.n250 B.n171 585
R245 B.n248 B.n247 585
R246 B.n246 B.n172 585
R247 B.n245 B.n244 585
R248 B.n242 B.n173 585
R249 B.n240 B.n239 585
R250 B.n238 B.n174 585
R251 B.n237 B.n236 585
R252 B.n234 B.n175 585
R253 B.n232 B.n231 585
R254 B.n230 B.n176 585
R255 B.n229 B.n228 585
R256 B.n226 B.n177 585
R257 B.n224 B.n223 585
R258 B.n222 B.n178 585
R259 B.n221 B.n220 585
R260 B.n218 B.n179 585
R261 B.n216 B.n215 585
R262 B.n214 B.n180 585
R263 B.n213 B.n212 585
R264 B.n210 B.n181 585
R265 B.n208 B.n207 585
R266 B.n206 B.n182 585
R267 B.n205 B.n204 585
R268 B.n202 B.n183 585
R269 B.n200 B.n199 585
R270 B.n198 B.n184 585
R271 B.n197 B.n196 585
R272 B.n194 B.n185 585
R273 B.n192 B.n191 585
R274 B.n190 B.n186 585
R275 B.n189 B.n188 585
R276 B.n135 B.n134 585
R277 B.n136 B.n135 585
R278 B.n366 B.n365 585
R279 B.n367 B.n366 585
R280 B.n131 B.n130 585
R281 B.n132 B.n131 585
R282 B.n375 B.n374 585
R283 B.n374 B.n373 585
R284 B.n376 B.n129 585
R285 B.n129 B.n128 585
R286 B.n378 B.n377 585
R287 B.n379 B.n378 585
R288 B.n123 B.n122 585
R289 B.n124 B.n123 585
R290 B.n387 B.n386 585
R291 B.n386 B.n385 585
R292 B.n388 B.n121 585
R293 B.n121 B.n120 585
R294 B.n390 B.n389 585
R295 B.n391 B.n390 585
R296 B.n115 B.n114 585
R297 B.n116 B.n115 585
R298 B.n399 B.n398 585
R299 B.n398 B.n397 585
R300 B.n400 B.n113 585
R301 B.n113 B.n112 585
R302 B.n402 B.n401 585
R303 B.n403 B.n402 585
R304 B.n107 B.n106 585
R305 B.n108 B.n107 585
R306 B.n411 B.n410 585
R307 B.n410 B.n409 585
R308 B.n412 B.n105 585
R309 B.n105 B.n103 585
R310 B.n414 B.n413 585
R311 B.n415 B.n414 585
R312 B.n99 B.n98 585
R313 B.n104 B.n99 585
R314 B.n425 B.n424 585
R315 B.n424 B.n423 585
R316 B.n426 B.n97 585
R317 B.n422 B.n97 585
R318 B.n428 B.n427 585
R319 B.n429 B.n428 585
R320 B.n3 B.n0 585
R321 B.n4 B.n3 585
R322 B.n686 B.n1 585
R323 B.n687 B.n686 585
R324 B.n685 B.n684 585
R325 B.n685 B.n8 585
R326 B.n683 B.n9 585
R327 B.n12 B.n9 585
R328 B.n682 B.n681 585
R329 B.n681 B.n680 585
R330 B.n11 B.n10 585
R331 B.n679 B.n11 585
R332 B.n677 B.n676 585
R333 B.n678 B.n677 585
R334 B.n675 B.n17 585
R335 B.n17 B.n16 585
R336 B.n674 B.n673 585
R337 B.n673 B.n672 585
R338 B.n19 B.n18 585
R339 B.n671 B.n19 585
R340 B.n669 B.n668 585
R341 B.n670 B.n669 585
R342 B.n667 B.n24 585
R343 B.n24 B.n23 585
R344 B.n666 B.n665 585
R345 B.n665 B.n664 585
R346 B.n26 B.n25 585
R347 B.n663 B.n26 585
R348 B.n661 B.n660 585
R349 B.n662 B.n661 585
R350 B.n659 B.n31 585
R351 B.n31 B.n30 585
R352 B.n658 B.n657 585
R353 B.n657 B.n656 585
R354 B.n33 B.n32 585
R355 B.n655 B.n33 585
R356 B.n653 B.n652 585
R357 B.n654 B.n653 585
R358 B.n651 B.n38 585
R359 B.n38 B.n37 585
R360 B.n650 B.n649 585
R361 B.n649 B.n648 585
R362 B.n40 B.n39 585
R363 B.n647 B.n40 585
R364 B.n645 B.n644 585
R365 B.n646 B.n645 585
R366 B.n690 B.n689 585
R367 B.n688 B.n2 585
R368 B.n645 B.n45 478.086
R369 B.n464 B.n43 478.086
R370 B.n368 B.n135 478.086
R371 B.n366 B.n137 478.086
R372 B.n72 B.t16 288.721
R373 B.n166 B.t20 288.721
R374 B.n66 B.t9 288.719
R375 B.n158 B.t14 288.719
R376 B.n73 B.t17 272.817
R377 B.n167 B.t19 272.817
R378 B.n67 B.t10 272.817
R379 B.n159 B.t13 272.817
R380 B.n465 B.n44 256.663
R381 B.n467 B.n44 256.663
R382 B.n473 B.n44 256.663
R383 B.n475 B.n44 256.663
R384 B.n481 B.n44 256.663
R385 B.n483 B.n44 256.663
R386 B.n489 B.n44 256.663
R387 B.n491 B.n44 256.663
R388 B.n497 B.n44 256.663
R389 B.n499 B.n44 256.663
R390 B.n505 B.n44 256.663
R391 B.n507 B.n44 256.663
R392 B.n513 B.n44 256.663
R393 B.n515 B.n44 256.663
R394 B.n521 B.n44 256.663
R395 B.n523 B.n44 256.663
R396 B.n529 B.n44 256.663
R397 B.n531 B.n44 256.663
R398 B.n537 B.n44 256.663
R399 B.n75 B.n44 256.663
R400 B.n543 B.n44 256.663
R401 B.n549 B.n44 256.663
R402 B.n551 B.n44 256.663
R403 B.n557 B.n44 256.663
R404 B.n559 B.n44 256.663
R405 B.n566 B.n44 256.663
R406 B.n568 B.n44 256.663
R407 B.n574 B.n44 256.663
R408 B.n576 B.n44 256.663
R409 B.n582 B.n44 256.663
R410 B.n584 B.n44 256.663
R411 B.n590 B.n44 256.663
R412 B.n592 B.n44 256.663
R413 B.n598 B.n44 256.663
R414 B.n600 B.n44 256.663
R415 B.n606 B.n44 256.663
R416 B.n608 B.n44 256.663
R417 B.n614 B.n44 256.663
R418 B.n616 B.n44 256.663
R419 B.n622 B.n44 256.663
R420 B.n624 B.n44 256.663
R421 B.n630 B.n44 256.663
R422 B.n632 B.n44 256.663
R423 B.n638 B.n44 256.663
R424 B.n640 B.n44 256.663
R425 B.n361 B.n136 256.663
R426 B.n139 B.n136 256.663
R427 B.n354 B.n136 256.663
R428 B.n348 B.n136 256.663
R429 B.n346 B.n136 256.663
R430 B.n340 B.n136 256.663
R431 B.n338 B.n136 256.663
R432 B.n332 B.n136 256.663
R433 B.n330 B.n136 256.663
R434 B.n324 B.n136 256.663
R435 B.n322 B.n136 256.663
R436 B.n316 B.n136 256.663
R437 B.n314 B.n136 256.663
R438 B.n308 B.n136 256.663
R439 B.n306 B.n136 256.663
R440 B.n300 B.n136 256.663
R441 B.n298 B.n136 256.663
R442 B.n292 B.n136 256.663
R443 B.n290 B.n136 256.663
R444 B.n283 B.n136 256.663
R445 B.n281 B.n136 256.663
R446 B.n275 B.n136 256.663
R447 B.n273 B.n136 256.663
R448 B.n267 B.n136 256.663
R449 B.n265 B.n136 256.663
R450 B.n259 B.n136 256.663
R451 B.n257 B.n136 256.663
R452 B.n251 B.n136 256.663
R453 B.n249 B.n136 256.663
R454 B.n243 B.n136 256.663
R455 B.n241 B.n136 256.663
R456 B.n235 B.n136 256.663
R457 B.n233 B.n136 256.663
R458 B.n227 B.n136 256.663
R459 B.n225 B.n136 256.663
R460 B.n219 B.n136 256.663
R461 B.n217 B.n136 256.663
R462 B.n211 B.n136 256.663
R463 B.n209 B.n136 256.663
R464 B.n203 B.n136 256.663
R465 B.n201 B.n136 256.663
R466 B.n195 B.n136 256.663
R467 B.n193 B.n136 256.663
R468 B.n187 B.n136 256.663
R469 B.n692 B.n691 256.663
R470 B.n641 B.n639 163.367
R471 B.n637 B.n47 163.367
R472 B.n633 B.n631 163.367
R473 B.n629 B.n49 163.367
R474 B.n625 B.n623 163.367
R475 B.n621 B.n51 163.367
R476 B.n617 B.n615 163.367
R477 B.n613 B.n53 163.367
R478 B.n609 B.n607 163.367
R479 B.n605 B.n55 163.367
R480 B.n601 B.n599 163.367
R481 B.n597 B.n57 163.367
R482 B.n593 B.n591 163.367
R483 B.n589 B.n59 163.367
R484 B.n585 B.n583 163.367
R485 B.n581 B.n61 163.367
R486 B.n577 B.n575 163.367
R487 B.n573 B.n63 163.367
R488 B.n569 B.n567 163.367
R489 B.n565 B.n65 163.367
R490 B.n560 B.n558 163.367
R491 B.n556 B.n69 163.367
R492 B.n552 B.n550 163.367
R493 B.n548 B.n71 163.367
R494 B.n544 B.n542 163.367
R495 B.n539 B.n538 163.367
R496 B.n536 B.n77 163.367
R497 B.n532 B.n530 163.367
R498 B.n528 B.n79 163.367
R499 B.n524 B.n522 163.367
R500 B.n520 B.n81 163.367
R501 B.n516 B.n514 163.367
R502 B.n512 B.n83 163.367
R503 B.n508 B.n506 163.367
R504 B.n504 B.n85 163.367
R505 B.n500 B.n498 163.367
R506 B.n496 B.n87 163.367
R507 B.n492 B.n490 163.367
R508 B.n488 B.n89 163.367
R509 B.n484 B.n482 163.367
R510 B.n480 B.n91 163.367
R511 B.n476 B.n474 163.367
R512 B.n472 B.n93 163.367
R513 B.n468 B.n466 163.367
R514 B.n368 B.n133 163.367
R515 B.n372 B.n133 163.367
R516 B.n372 B.n127 163.367
R517 B.n380 B.n127 163.367
R518 B.n380 B.n125 163.367
R519 B.n384 B.n125 163.367
R520 B.n384 B.n119 163.367
R521 B.n392 B.n119 163.367
R522 B.n392 B.n117 163.367
R523 B.n396 B.n117 163.367
R524 B.n396 B.n111 163.367
R525 B.n404 B.n111 163.367
R526 B.n404 B.n109 163.367
R527 B.n408 B.n109 163.367
R528 B.n408 B.n102 163.367
R529 B.n416 B.n102 163.367
R530 B.n416 B.n100 163.367
R531 B.n421 B.n100 163.367
R532 B.n421 B.n96 163.367
R533 B.n430 B.n96 163.367
R534 B.n431 B.n430 163.367
R535 B.n431 B.n5 163.367
R536 B.n6 B.n5 163.367
R537 B.n7 B.n6 163.367
R538 B.n437 B.n7 163.367
R539 B.n438 B.n437 163.367
R540 B.n438 B.n13 163.367
R541 B.n14 B.n13 163.367
R542 B.n15 B.n14 163.367
R543 B.n443 B.n15 163.367
R544 B.n443 B.n20 163.367
R545 B.n21 B.n20 163.367
R546 B.n22 B.n21 163.367
R547 B.n448 B.n22 163.367
R548 B.n448 B.n27 163.367
R549 B.n28 B.n27 163.367
R550 B.n29 B.n28 163.367
R551 B.n453 B.n29 163.367
R552 B.n453 B.n34 163.367
R553 B.n35 B.n34 163.367
R554 B.n36 B.n35 163.367
R555 B.n458 B.n36 163.367
R556 B.n458 B.n41 163.367
R557 B.n42 B.n41 163.367
R558 B.n43 B.n42 163.367
R559 B.n362 B.n360 163.367
R560 B.n360 B.n359 163.367
R561 B.n356 B.n355 163.367
R562 B.n353 B.n141 163.367
R563 B.n349 B.n347 163.367
R564 B.n345 B.n143 163.367
R565 B.n341 B.n339 163.367
R566 B.n337 B.n145 163.367
R567 B.n333 B.n331 163.367
R568 B.n329 B.n147 163.367
R569 B.n325 B.n323 163.367
R570 B.n321 B.n149 163.367
R571 B.n317 B.n315 163.367
R572 B.n313 B.n151 163.367
R573 B.n309 B.n307 163.367
R574 B.n305 B.n153 163.367
R575 B.n301 B.n299 163.367
R576 B.n297 B.n155 163.367
R577 B.n293 B.n291 163.367
R578 B.n289 B.n157 163.367
R579 B.n284 B.n282 163.367
R580 B.n280 B.n161 163.367
R581 B.n276 B.n274 163.367
R582 B.n272 B.n163 163.367
R583 B.n268 B.n266 163.367
R584 B.n264 B.n165 163.367
R585 B.n260 B.n258 163.367
R586 B.n256 B.n170 163.367
R587 B.n252 B.n250 163.367
R588 B.n248 B.n172 163.367
R589 B.n244 B.n242 163.367
R590 B.n240 B.n174 163.367
R591 B.n236 B.n234 163.367
R592 B.n232 B.n176 163.367
R593 B.n228 B.n226 163.367
R594 B.n224 B.n178 163.367
R595 B.n220 B.n218 163.367
R596 B.n216 B.n180 163.367
R597 B.n212 B.n210 163.367
R598 B.n208 B.n182 163.367
R599 B.n204 B.n202 163.367
R600 B.n200 B.n184 163.367
R601 B.n196 B.n194 163.367
R602 B.n192 B.n186 163.367
R603 B.n188 B.n135 163.367
R604 B.n366 B.n131 163.367
R605 B.n374 B.n131 163.367
R606 B.n374 B.n129 163.367
R607 B.n378 B.n129 163.367
R608 B.n378 B.n123 163.367
R609 B.n386 B.n123 163.367
R610 B.n386 B.n121 163.367
R611 B.n390 B.n121 163.367
R612 B.n390 B.n115 163.367
R613 B.n398 B.n115 163.367
R614 B.n398 B.n113 163.367
R615 B.n402 B.n113 163.367
R616 B.n402 B.n107 163.367
R617 B.n410 B.n107 163.367
R618 B.n410 B.n105 163.367
R619 B.n414 B.n105 163.367
R620 B.n414 B.n99 163.367
R621 B.n424 B.n99 163.367
R622 B.n424 B.n97 163.367
R623 B.n428 B.n97 163.367
R624 B.n428 B.n3 163.367
R625 B.n690 B.n3 163.367
R626 B.n686 B.n2 163.367
R627 B.n686 B.n685 163.367
R628 B.n685 B.n9 163.367
R629 B.n681 B.n9 163.367
R630 B.n681 B.n11 163.367
R631 B.n677 B.n11 163.367
R632 B.n677 B.n17 163.367
R633 B.n673 B.n17 163.367
R634 B.n673 B.n19 163.367
R635 B.n669 B.n19 163.367
R636 B.n669 B.n24 163.367
R637 B.n665 B.n24 163.367
R638 B.n665 B.n26 163.367
R639 B.n661 B.n26 163.367
R640 B.n661 B.n31 163.367
R641 B.n657 B.n31 163.367
R642 B.n657 B.n33 163.367
R643 B.n653 B.n33 163.367
R644 B.n653 B.n38 163.367
R645 B.n649 B.n38 163.367
R646 B.n649 B.n40 163.367
R647 B.n645 B.n40 163.367
R648 B.n367 B.n136 84.8435
R649 B.n646 B.n44 84.8435
R650 B.n640 B.n45 71.676
R651 B.n639 B.n638 71.676
R652 B.n632 B.n47 71.676
R653 B.n631 B.n630 71.676
R654 B.n624 B.n49 71.676
R655 B.n623 B.n622 71.676
R656 B.n616 B.n51 71.676
R657 B.n615 B.n614 71.676
R658 B.n608 B.n53 71.676
R659 B.n607 B.n606 71.676
R660 B.n600 B.n55 71.676
R661 B.n599 B.n598 71.676
R662 B.n592 B.n57 71.676
R663 B.n591 B.n590 71.676
R664 B.n584 B.n59 71.676
R665 B.n583 B.n582 71.676
R666 B.n576 B.n61 71.676
R667 B.n575 B.n574 71.676
R668 B.n568 B.n63 71.676
R669 B.n567 B.n566 71.676
R670 B.n559 B.n65 71.676
R671 B.n558 B.n557 71.676
R672 B.n551 B.n69 71.676
R673 B.n550 B.n549 71.676
R674 B.n543 B.n71 71.676
R675 B.n542 B.n75 71.676
R676 B.n538 B.n537 71.676
R677 B.n531 B.n77 71.676
R678 B.n530 B.n529 71.676
R679 B.n523 B.n79 71.676
R680 B.n522 B.n521 71.676
R681 B.n515 B.n81 71.676
R682 B.n514 B.n513 71.676
R683 B.n507 B.n83 71.676
R684 B.n506 B.n505 71.676
R685 B.n499 B.n85 71.676
R686 B.n498 B.n497 71.676
R687 B.n491 B.n87 71.676
R688 B.n490 B.n489 71.676
R689 B.n483 B.n89 71.676
R690 B.n482 B.n481 71.676
R691 B.n475 B.n91 71.676
R692 B.n474 B.n473 71.676
R693 B.n467 B.n93 71.676
R694 B.n466 B.n465 71.676
R695 B.n465 B.n464 71.676
R696 B.n468 B.n467 71.676
R697 B.n473 B.n472 71.676
R698 B.n476 B.n475 71.676
R699 B.n481 B.n480 71.676
R700 B.n484 B.n483 71.676
R701 B.n489 B.n488 71.676
R702 B.n492 B.n491 71.676
R703 B.n497 B.n496 71.676
R704 B.n500 B.n499 71.676
R705 B.n505 B.n504 71.676
R706 B.n508 B.n507 71.676
R707 B.n513 B.n512 71.676
R708 B.n516 B.n515 71.676
R709 B.n521 B.n520 71.676
R710 B.n524 B.n523 71.676
R711 B.n529 B.n528 71.676
R712 B.n532 B.n531 71.676
R713 B.n537 B.n536 71.676
R714 B.n539 B.n75 71.676
R715 B.n544 B.n543 71.676
R716 B.n549 B.n548 71.676
R717 B.n552 B.n551 71.676
R718 B.n557 B.n556 71.676
R719 B.n560 B.n559 71.676
R720 B.n566 B.n565 71.676
R721 B.n569 B.n568 71.676
R722 B.n574 B.n573 71.676
R723 B.n577 B.n576 71.676
R724 B.n582 B.n581 71.676
R725 B.n585 B.n584 71.676
R726 B.n590 B.n589 71.676
R727 B.n593 B.n592 71.676
R728 B.n598 B.n597 71.676
R729 B.n601 B.n600 71.676
R730 B.n606 B.n605 71.676
R731 B.n609 B.n608 71.676
R732 B.n614 B.n613 71.676
R733 B.n617 B.n616 71.676
R734 B.n622 B.n621 71.676
R735 B.n625 B.n624 71.676
R736 B.n630 B.n629 71.676
R737 B.n633 B.n632 71.676
R738 B.n638 B.n637 71.676
R739 B.n641 B.n640 71.676
R740 B.n361 B.n137 71.676
R741 B.n359 B.n139 71.676
R742 B.n355 B.n354 71.676
R743 B.n348 B.n141 71.676
R744 B.n347 B.n346 71.676
R745 B.n340 B.n143 71.676
R746 B.n339 B.n338 71.676
R747 B.n332 B.n145 71.676
R748 B.n331 B.n330 71.676
R749 B.n324 B.n147 71.676
R750 B.n323 B.n322 71.676
R751 B.n316 B.n149 71.676
R752 B.n315 B.n314 71.676
R753 B.n308 B.n151 71.676
R754 B.n307 B.n306 71.676
R755 B.n300 B.n153 71.676
R756 B.n299 B.n298 71.676
R757 B.n292 B.n155 71.676
R758 B.n291 B.n290 71.676
R759 B.n283 B.n157 71.676
R760 B.n282 B.n281 71.676
R761 B.n275 B.n161 71.676
R762 B.n274 B.n273 71.676
R763 B.n267 B.n163 71.676
R764 B.n266 B.n265 71.676
R765 B.n259 B.n165 71.676
R766 B.n258 B.n257 71.676
R767 B.n251 B.n170 71.676
R768 B.n250 B.n249 71.676
R769 B.n243 B.n172 71.676
R770 B.n242 B.n241 71.676
R771 B.n235 B.n174 71.676
R772 B.n234 B.n233 71.676
R773 B.n227 B.n176 71.676
R774 B.n226 B.n225 71.676
R775 B.n219 B.n178 71.676
R776 B.n218 B.n217 71.676
R777 B.n211 B.n180 71.676
R778 B.n210 B.n209 71.676
R779 B.n203 B.n182 71.676
R780 B.n202 B.n201 71.676
R781 B.n195 B.n184 71.676
R782 B.n194 B.n193 71.676
R783 B.n187 B.n186 71.676
R784 B.n362 B.n361 71.676
R785 B.n356 B.n139 71.676
R786 B.n354 B.n353 71.676
R787 B.n349 B.n348 71.676
R788 B.n346 B.n345 71.676
R789 B.n341 B.n340 71.676
R790 B.n338 B.n337 71.676
R791 B.n333 B.n332 71.676
R792 B.n330 B.n329 71.676
R793 B.n325 B.n324 71.676
R794 B.n322 B.n321 71.676
R795 B.n317 B.n316 71.676
R796 B.n314 B.n313 71.676
R797 B.n309 B.n308 71.676
R798 B.n306 B.n305 71.676
R799 B.n301 B.n300 71.676
R800 B.n298 B.n297 71.676
R801 B.n293 B.n292 71.676
R802 B.n290 B.n289 71.676
R803 B.n284 B.n283 71.676
R804 B.n281 B.n280 71.676
R805 B.n276 B.n275 71.676
R806 B.n273 B.n272 71.676
R807 B.n268 B.n267 71.676
R808 B.n265 B.n264 71.676
R809 B.n260 B.n259 71.676
R810 B.n257 B.n256 71.676
R811 B.n252 B.n251 71.676
R812 B.n249 B.n248 71.676
R813 B.n244 B.n243 71.676
R814 B.n241 B.n240 71.676
R815 B.n236 B.n235 71.676
R816 B.n233 B.n232 71.676
R817 B.n228 B.n227 71.676
R818 B.n225 B.n224 71.676
R819 B.n220 B.n219 71.676
R820 B.n217 B.n216 71.676
R821 B.n212 B.n211 71.676
R822 B.n209 B.n208 71.676
R823 B.n204 B.n203 71.676
R824 B.n201 B.n200 71.676
R825 B.n196 B.n195 71.676
R826 B.n193 B.n192 71.676
R827 B.n188 B.n187 71.676
R828 B.n691 B.n690 71.676
R829 B.n691 B.n2 71.676
R830 B.n563 B.n67 59.5399
R831 B.n74 B.n73 59.5399
R832 B.n168 B.n167 59.5399
R833 B.n286 B.n159 59.5399
R834 B.n367 B.n132 44.724
R835 B.n373 B.n132 44.724
R836 B.n373 B.n128 44.724
R837 B.n379 B.n128 44.724
R838 B.n385 B.n124 44.724
R839 B.n385 B.n120 44.724
R840 B.n391 B.n120 44.724
R841 B.n391 B.n116 44.724
R842 B.n397 B.n116 44.724
R843 B.n403 B.n112 44.724
R844 B.n409 B.n108 44.724
R845 B.n415 B.n103 44.724
R846 B.n415 B.n104 44.724
R847 B.n423 B.n422 44.724
R848 B.n429 B.n4 44.724
R849 B.n689 B.n4 44.724
R850 B.n689 B.n688 44.724
R851 B.n688 B.n687 44.724
R852 B.n687 B.n8 44.724
R853 B.n680 B.n12 44.724
R854 B.n679 B.n678 44.724
R855 B.n678 B.n16 44.724
R856 B.n672 B.n671 44.724
R857 B.n670 B.n23 44.724
R858 B.n664 B.n663 44.724
R859 B.n663 B.n662 44.724
R860 B.n662 B.n30 44.724
R861 B.n656 B.n30 44.724
R862 B.n656 B.n655 44.724
R863 B.n654 B.n37 44.724
R864 B.n648 B.n37 44.724
R865 B.n648 B.n647 44.724
R866 B.n647 B.n646 44.724
R867 B.t0 B.n112 42.7509
R868 B.t21 B.n23 42.7509
R869 B.n409 B.t3 38.8047
R870 B.n672 B.t2 38.8047
R871 B.n423 B.t1 32.2277
R872 B.n680 B.t23 32.2277
R873 B.n365 B.n364 31.0639
R874 B.n369 B.n134 31.0639
R875 B.n463 B.n462 31.0639
R876 B.n644 B.n643 31.0639
R877 B.n422 B.t6 30.9123
R878 B.n12 B.t5 30.9123
R879 B.t12 B.n124 25.6507
R880 B.n655 B.t8 25.6507
R881 B.t22 B.n108 24.3353
R882 B.n671 B.t4 24.3353
R883 B.n403 B.t22 20.3891
R884 B.t4 B.n670 20.3891
R885 B.n379 B.t12 19.0737
R886 B.t8 B.n654 19.0737
R887 B B.n692 18.0485
R888 B.n67 B.n66 15.9035
R889 B.n73 B.n72 15.9035
R890 B.n167 B.n166 15.9035
R891 B.n159 B.n158 15.9035
R892 B.n429 B.t6 13.8122
R893 B.t5 B.n8 13.8122
R894 B.n104 B.t1 12.4968
R895 B.t23 B.n679 12.4968
R896 B.n365 B.n130 10.6151
R897 B.n375 B.n130 10.6151
R898 B.n376 B.n375 10.6151
R899 B.n377 B.n376 10.6151
R900 B.n377 B.n122 10.6151
R901 B.n387 B.n122 10.6151
R902 B.n388 B.n387 10.6151
R903 B.n389 B.n388 10.6151
R904 B.n389 B.n114 10.6151
R905 B.n399 B.n114 10.6151
R906 B.n400 B.n399 10.6151
R907 B.n401 B.n400 10.6151
R908 B.n401 B.n106 10.6151
R909 B.n411 B.n106 10.6151
R910 B.n412 B.n411 10.6151
R911 B.n413 B.n412 10.6151
R912 B.n413 B.n98 10.6151
R913 B.n425 B.n98 10.6151
R914 B.n426 B.n425 10.6151
R915 B.n427 B.n426 10.6151
R916 B.n427 B.n0 10.6151
R917 B.n364 B.n363 10.6151
R918 B.n363 B.n138 10.6151
R919 B.n358 B.n138 10.6151
R920 B.n358 B.n357 10.6151
R921 B.n357 B.n140 10.6151
R922 B.n352 B.n140 10.6151
R923 B.n352 B.n351 10.6151
R924 B.n351 B.n350 10.6151
R925 B.n350 B.n142 10.6151
R926 B.n344 B.n142 10.6151
R927 B.n344 B.n343 10.6151
R928 B.n343 B.n342 10.6151
R929 B.n342 B.n144 10.6151
R930 B.n336 B.n144 10.6151
R931 B.n336 B.n335 10.6151
R932 B.n335 B.n334 10.6151
R933 B.n334 B.n146 10.6151
R934 B.n328 B.n146 10.6151
R935 B.n328 B.n327 10.6151
R936 B.n327 B.n326 10.6151
R937 B.n326 B.n148 10.6151
R938 B.n320 B.n148 10.6151
R939 B.n320 B.n319 10.6151
R940 B.n319 B.n318 10.6151
R941 B.n318 B.n150 10.6151
R942 B.n312 B.n150 10.6151
R943 B.n312 B.n311 10.6151
R944 B.n311 B.n310 10.6151
R945 B.n310 B.n152 10.6151
R946 B.n304 B.n152 10.6151
R947 B.n304 B.n303 10.6151
R948 B.n303 B.n302 10.6151
R949 B.n302 B.n154 10.6151
R950 B.n296 B.n154 10.6151
R951 B.n296 B.n295 10.6151
R952 B.n295 B.n294 10.6151
R953 B.n294 B.n156 10.6151
R954 B.n288 B.n156 10.6151
R955 B.n288 B.n287 10.6151
R956 B.n285 B.n160 10.6151
R957 B.n279 B.n160 10.6151
R958 B.n279 B.n278 10.6151
R959 B.n278 B.n277 10.6151
R960 B.n277 B.n162 10.6151
R961 B.n271 B.n162 10.6151
R962 B.n271 B.n270 10.6151
R963 B.n270 B.n269 10.6151
R964 B.n269 B.n164 10.6151
R965 B.n263 B.n262 10.6151
R966 B.n262 B.n261 10.6151
R967 B.n261 B.n169 10.6151
R968 B.n255 B.n169 10.6151
R969 B.n255 B.n254 10.6151
R970 B.n254 B.n253 10.6151
R971 B.n253 B.n171 10.6151
R972 B.n247 B.n171 10.6151
R973 B.n247 B.n246 10.6151
R974 B.n246 B.n245 10.6151
R975 B.n245 B.n173 10.6151
R976 B.n239 B.n173 10.6151
R977 B.n239 B.n238 10.6151
R978 B.n238 B.n237 10.6151
R979 B.n237 B.n175 10.6151
R980 B.n231 B.n175 10.6151
R981 B.n231 B.n230 10.6151
R982 B.n230 B.n229 10.6151
R983 B.n229 B.n177 10.6151
R984 B.n223 B.n177 10.6151
R985 B.n223 B.n222 10.6151
R986 B.n222 B.n221 10.6151
R987 B.n221 B.n179 10.6151
R988 B.n215 B.n179 10.6151
R989 B.n215 B.n214 10.6151
R990 B.n214 B.n213 10.6151
R991 B.n213 B.n181 10.6151
R992 B.n207 B.n181 10.6151
R993 B.n207 B.n206 10.6151
R994 B.n206 B.n205 10.6151
R995 B.n205 B.n183 10.6151
R996 B.n199 B.n183 10.6151
R997 B.n199 B.n198 10.6151
R998 B.n198 B.n197 10.6151
R999 B.n197 B.n185 10.6151
R1000 B.n191 B.n185 10.6151
R1001 B.n191 B.n190 10.6151
R1002 B.n190 B.n189 10.6151
R1003 B.n189 B.n134 10.6151
R1004 B.n370 B.n369 10.6151
R1005 B.n371 B.n370 10.6151
R1006 B.n371 B.n126 10.6151
R1007 B.n381 B.n126 10.6151
R1008 B.n382 B.n381 10.6151
R1009 B.n383 B.n382 10.6151
R1010 B.n383 B.n118 10.6151
R1011 B.n393 B.n118 10.6151
R1012 B.n394 B.n393 10.6151
R1013 B.n395 B.n394 10.6151
R1014 B.n395 B.n110 10.6151
R1015 B.n405 B.n110 10.6151
R1016 B.n406 B.n405 10.6151
R1017 B.n407 B.n406 10.6151
R1018 B.n407 B.n101 10.6151
R1019 B.n417 B.n101 10.6151
R1020 B.n418 B.n417 10.6151
R1021 B.n420 B.n418 10.6151
R1022 B.n420 B.n419 10.6151
R1023 B.n419 B.n95 10.6151
R1024 B.n432 B.n95 10.6151
R1025 B.n433 B.n432 10.6151
R1026 B.n434 B.n433 10.6151
R1027 B.n435 B.n434 10.6151
R1028 B.n436 B.n435 10.6151
R1029 B.n439 B.n436 10.6151
R1030 B.n440 B.n439 10.6151
R1031 B.n441 B.n440 10.6151
R1032 B.n442 B.n441 10.6151
R1033 B.n444 B.n442 10.6151
R1034 B.n445 B.n444 10.6151
R1035 B.n446 B.n445 10.6151
R1036 B.n447 B.n446 10.6151
R1037 B.n449 B.n447 10.6151
R1038 B.n450 B.n449 10.6151
R1039 B.n451 B.n450 10.6151
R1040 B.n452 B.n451 10.6151
R1041 B.n454 B.n452 10.6151
R1042 B.n455 B.n454 10.6151
R1043 B.n456 B.n455 10.6151
R1044 B.n457 B.n456 10.6151
R1045 B.n459 B.n457 10.6151
R1046 B.n460 B.n459 10.6151
R1047 B.n461 B.n460 10.6151
R1048 B.n462 B.n461 10.6151
R1049 B.n684 B.n1 10.6151
R1050 B.n684 B.n683 10.6151
R1051 B.n683 B.n682 10.6151
R1052 B.n682 B.n10 10.6151
R1053 B.n676 B.n10 10.6151
R1054 B.n676 B.n675 10.6151
R1055 B.n675 B.n674 10.6151
R1056 B.n674 B.n18 10.6151
R1057 B.n668 B.n18 10.6151
R1058 B.n668 B.n667 10.6151
R1059 B.n667 B.n666 10.6151
R1060 B.n666 B.n25 10.6151
R1061 B.n660 B.n25 10.6151
R1062 B.n660 B.n659 10.6151
R1063 B.n659 B.n658 10.6151
R1064 B.n658 B.n32 10.6151
R1065 B.n652 B.n32 10.6151
R1066 B.n652 B.n651 10.6151
R1067 B.n651 B.n650 10.6151
R1068 B.n650 B.n39 10.6151
R1069 B.n644 B.n39 10.6151
R1070 B.n643 B.n642 10.6151
R1071 B.n642 B.n46 10.6151
R1072 B.n636 B.n46 10.6151
R1073 B.n636 B.n635 10.6151
R1074 B.n635 B.n634 10.6151
R1075 B.n634 B.n48 10.6151
R1076 B.n628 B.n48 10.6151
R1077 B.n628 B.n627 10.6151
R1078 B.n627 B.n626 10.6151
R1079 B.n626 B.n50 10.6151
R1080 B.n620 B.n50 10.6151
R1081 B.n620 B.n619 10.6151
R1082 B.n619 B.n618 10.6151
R1083 B.n618 B.n52 10.6151
R1084 B.n612 B.n52 10.6151
R1085 B.n612 B.n611 10.6151
R1086 B.n611 B.n610 10.6151
R1087 B.n610 B.n54 10.6151
R1088 B.n604 B.n54 10.6151
R1089 B.n604 B.n603 10.6151
R1090 B.n603 B.n602 10.6151
R1091 B.n602 B.n56 10.6151
R1092 B.n596 B.n56 10.6151
R1093 B.n596 B.n595 10.6151
R1094 B.n595 B.n594 10.6151
R1095 B.n594 B.n58 10.6151
R1096 B.n588 B.n58 10.6151
R1097 B.n588 B.n587 10.6151
R1098 B.n587 B.n586 10.6151
R1099 B.n586 B.n60 10.6151
R1100 B.n580 B.n60 10.6151
R1101 B.n580 B.n579 10.6151
R1102 B.n579 B.n578 10.6151
R1103 B.n578 B.n62 10.6151
R1104 B.n572 B.n62 10.6151
R1105 B.n572 B.n571 10.6151
R1106 B.n571 B.n570 10.6151
R1107 B.n570 B.n64 10.6151
R1108 B.n564 B.n64 10.6151
R1109 B.n562 B.n561 10.6151
R1110 B.n561 B.n68 10.6151
R1111 B.n555 B.n68 10.6151
R1112 B.n555 B.n554 10.6151
R1113 B.n554 B.n553 10.6151
R1114 B.n553 B.n70 10.6151
R1115 B.n547 B.n70 10.6151
R1116 B.n547 B.n546 10.6151
R1117 B.n546 B.n545 10.6151
R1118 B.n541 B.n540 10.6151
R1119 B.n540 B.n76 10.6151
R1120 B.n535 B.n76 10.6151
R1121 B.n535 B.n534 10.6151
R1122 B.n534 B.n533 10.6151
R1123 B.n533 B.n78 10.6151
R1124 B.n527 B.n78 10.6151
R1125 B.n527 B.n526 10.6151
R1126 B.n526 B.n525 10.6151
R1127 B.n525 B.n80 10.6151
R1128 B.n519 B.n80 10.6151
R1129 B.n519 B.n518 10.6151
R1130 B.n518 B.n517 10.6151
R1131 B.n517 B.n82 10.6151
R1132 B.n511 B.n82 10.6151
R1133 B.n511 B.n510 10.6151
R1134 B.n510 B.n509 10.6151
R1135 B.n509 B.n84 10.6151
R1136 B.n503 B.n84 10.6151
R1137 B.n503 B.n502 10.6151
R1138 B.n502 B.n501 10.6151
R1139 B.n501 B.n86 10.6151
R1140 B.n495 B.n86 10.6151
R1141 B.n495 B.n494 10.6151
R1142 B.n494 B.n493 10.6151
R1143 B.n493 B.n88 10.6151
R1144 B.n487 B.n88 10.6151
R1145 B.n487 B.n486 10.6151
R1146 B.n486 B.n485 10.6151
R1147 B.n485 B.n90 10.6151
R1148 B.n479 B.n90 10.6151
R1149 B.n479 B.n478 10.6151
R1150 B.n478 B.n477 10.6151
R1151 B.n477 B.n92 10.6151
R1152 B.n471 B.n92 10.6151
R1153 B.n471 B.n470 10.6151
R1154 B.n470 B.n469 10.6151
R1155 B.n469 B.n94 10.6151
R1156 B.n463 B.n94 10.6151
R1157 B.n287 B.n286 9.36635
R1158 B.n263 B.n168 9.36635
R1159 B.n564 B.n563 9.36635
R1160 B.n541 B.n74 9.36635
R1161 B.n692 B.n0 8.11757
R1162 B.n692 B.n1 8.11757
R1163 B.t3 B.n103 5.91978
R1164 B.t2 B.n16 5.91978
R1165 B.n397 B.t0 1.97359
R1166 B.n664 B.t21 1.97359
R1167 B.n286 B.n285 1.24928
R1168 B.n168 B.n164 1.24928
R1169 B.n563 B.n562 1.24928
R1170 B.n545 B.n74 1.24928
R1171 VP.n5 VP.t6 664.797
R1172 VP.n16 VP.t7 643.814
R1173 VP.n17 VP.t3 643.814
R1174 VP.n1 VP.t1 643.814
R1175 VP.n23 VP.t0 643.814
R1176 VP.n24 VP.t2 643.814
R1177 VP.n13 VP.t4 643.814
R1178 VP.n12 VP.t8 643.814
R1179 VP.n4 VP.t5 643.814
R1180 VP.n6 VP.t9 643.814
R1181 VP.n25 VP.n24 161.3
R1182 VP.n8 VP.n7 161.3
R1183 VP.n9 VP.n4 161.3
R1184 VP.n11 VP.n10 161.3
R1185 VP.n12 VP.n3 161.3
R1186 VP.n14 VP.n13 161.3
R1187 VP.n23 VP.n0 161.3
R1188 VP.n22 VP.n21 161.3
R1189 VP.n20 VP.n1 161.3
R1190 VP.n19 VP.n18 161.3
R1191 VP.n17 VP.n2 161.3
R1192 VP.n16 VP.n15 161.3
R1193 VP.n8 VP.n5 70.4033
R1194 VP.n17 VP.n16 48.2005
R1195 VP.n24 VP.n23 48.2005
R1196 VP.n13 VP.n12 48.2005
R1197 VP.n15 VP.n14 41.2353
R1198 VP.n18 VP.n1 37.246
R1199 VP.n22 VP.n1 37.246
R1200 VP.n11 VP.n4 37.246
R1201 VP.n7 VP.n4 37.246
R1202 VP.n6 VP.n5 20.9576
R1203 VP.n18 VP.n17 10.955
R1204 VP.n23 VP.n22 10.955
R1205 VP.n12 VP.n11 10.955
R1206 VP.n7 VP.n6 10.955
R1207 VP.n9 VP.n8 0.189894
R1208 VP.n10 VP.n9 0.189894
R1209 VP.n10 VP.n3 0.189894
R1210 VP.n14 VP.n3 0.189894
R1211 VP.n15 VP.n2 0.189894
R1212 VP.n19 VP.n2 0.189894
R1213 VP.n20 VP.n19 0.189894
R1214 VP.n21 VP.n20 0.189894
R1215 VP.n21 VP.n0 0.189894
R1216 VP.n25 VP.n0 0.189894
R1217 VP VP.n25 0.0516364
R1218 VDD1.n56 VDD1.n0 289.615
R1219 VDD1.n119 VDD1.n63 289.615
R1220 VDD1.n57 VDD1.n56 185
R1221 VDD1.n55 VDD1.n54 185
R1222 VDD1.n4 VDD1.n3 185
R1223 VDD1.n49 VDD1.n48 185
R1224 VDD1.n47 VDD1.n46 185
R1225 VDD1.n8 VDD1.n7 185
R1226 VDD1.n12 VDD1.n10 185
R1227 VDD1.n41 VDD1.n40 185
R1228 VDD1.n39 VDD1.n38 185
R1229 VDD1.n14 VDD1.n13 185
R1230 VDD1.n33 VDD1.n32 185
R1231 VDD1.n31 VDD1.n30 185
R1232 VDD1.n18 VDD1.n17 185
R1233 VDD1.n25 VDD1.n24 185
R1234 VDD1.n23 VDD1.n22 185
R1235 VDD1.n84 VDD1.n83 185
R1236 VDD1.n86 VDD1.n85 185
R1237 VDD1.n79 VDD1.n78 185
R1238 VDD1.n92 VDD1.n91 185
R1239 VDD1.n94 VDD1.n93 185
R1240 VDD1.n75 VDD1.n74 185
R1241 VDD1.n101 VDD1.n100 185
R1242 VDD1.n102 VDD1.n73 185
R1243 VDD1.n104 VDD1.n103 185
R1244 VDD1.n71 VDD1.n70 185
R1245 VDD1.n110 VDD1.n109 185
R1246 VDD1.n112 VDD1.n111 185
R1247 VDD1.n67 VDD1.n66 185
R1248 VDD1.n118 VDD1.n117 185
R1249 VDD1.n120 VDD1.n119 185
R1250 VDD1.n21 VDD1.t9 149.524
R1251 VDD1.n82 VDD1.t6 149.524
R1252 VDD1.n56 VDD1.n55 104.615
R1253 VDD1.n55 VDD1.n3 104.615
R1254 VDD1.n48 VDD1.n3 104.615
R1255 VDD1.n48 VDD1.n47 104.615
R1256 VDD1.n47 VDD1.n7 104.615
R1257 VDD1.n12 VDD1.n7 104.615
R1258 VDD1.n40 VDD1.n12 104.615
R1259 VDD1.n40 VDD1.n39 104.615
R1260 VDD1.n39 VDD1.n13 104.615
R1261 VDD1.n32 VDD1.n13 104.615
R1262 VDD1.n32 VDD1.n31 104.615
R1263 VDD1.n31 VDD1.n17 104.615
R1264 VDD1.n24 VDD1.n17 104.615
R1265 VDD1.n24 VDD1.n23 104.615
R1266 VDD1.n85 VDD1.n84 104.615
R1267 VDD1.n85 VDD1.n78 104.615
R1268 VDD1.n92 VDD1.n78 104.615
R1269 VDD1.n93 VDD1.n92 104.615
R1270 VDD1.n93 VDD1.n74 104.615
R1271 VDD1.n101 VDD1.n74 104.615
R1272 VDD1.n102 VDD1.n101 104.615
R1273 VDD1.n103 VDD1.n102 104.615
R1274 VDD1.n103 VDD1.n70 104.615
R1275 VDD1.n110 VDD1.n70 104.615
R1276 VDD1.n111 VDD1.n110 104.615
R1277 VDD1.n111 VDD1.n66 104.615
R1278 VDD1.n118 VDD1.n66 104.615
R1279 VDD1.n119 VDD1.n118 104.615
R1280 VDD1.n127 VDD1.n126 63.5342
R1281 VDD1.n62 VDD1.n61 63.0596
R1282 VDD1.n129 VDD1.n128 63.0594
R1283 VDD1.n125 VDD1.n124 63.0594
R1284 VDD1.n23 VDD1.t9 52.3082
R1285 VDD1.n84 VDD1.t6 52.3082
R1286 VDD1.n62 VDD1.n60 50.5407
R1287 VDD1.n125 VDD1.n123 50.5407
R1288 VDD1.n129 VDD1.n127 37.8802
R1289 VDD1.n10 VDD1.n8 13.1884
R1290 VDD1.n104 VDD1.n71 13.1884
R1291 VDD1.n46 VDD1.n45 12.8005
R1292 VDD1.n42 VDD1.n41 12.8005
R1293 VDD1.n105 VDD1.n73 12.8005
R1294 VDD1.n109 VDD1.n108 12.8005
R1295 VDD1.n49 VDD1.n6 12.0247
R1296 VDD1.n38 VDD1.n11 12.0247
R1297 VDD1.n100 VDD1.n99 12.0247
R1298 VDD1.n112 VDD1.n69 12.0247
R1299 VDD1.n50 VDD1.n4 11.249
R1300 VDD1.n37 VDD1.n14 11.249
R1301 VDD1.n98 VDD1.n75 11.249
R1302 VDD1.n113 VDD1.n67 11.249
R1303 VDD1.n54 VDD1.n53 10.4732
R1304 VDD1.n34 VDD1.n33 10.4732
R1305 VDD1.n95 VDD1.n94 10.4732
R1306 VDD1.n117 VDD1.n116 10.4732
R1307 VDD1.n22 VDD1.n21 10.2747
R1308 VDD1.n83 VDD1.n82 10.2747
R1309 VDD1.n57 VDD1.n2 9.69747
R1310 VDD1.n30 VDD1.n16 9.69747
R1311 VDD1.n91 VDD1.n77 9.69747
R1312 VDD1.n120 VDD1.n65 9.69747
R1313 VDD1.n60 VDD1.n59 9.45567
R1314 VDD1.n123 VDD1.n122 9.45567
R1315 VDD1.n20 VDD1.n19 9.3005
R1316 VDD1.n27 VDD1.n26 9.3005
R1317 VDD1.n29 VDD1.n28 9.3005
R1318 VDD1.n16 VDD1.n15 9.3005
R1319 VDD1.n35 VDD1.n34 9.3005
R1320 VDD1.n37 VDD1.n36 9.3005
R1321 VDD1.n11 VDD1.n9 9.3005
R1322 VDD1.n43 VDD1.n42 9.3005
R1323 VDD1.n59 VDD1.n58 9.3005
R1324 VDD1.n2 VDD1.n1 9.3005
R1325 VDD1.n53 VDD1.n52 9.3005
R1326 VDD1.n51 VDD1.n50 9.3005
R1327 VDD1.n6 VDD1.n5 9.3005
R1328 VDD1.n45 VDD1.n44 9.3005
R1329 VDD1.n122 VDD1.n121 9.3005
R1330 VDD1.n65 VDD1.n64 9.3005
R1331 VDD1.n116 VDD1.n115 9.3005
R1332 VDD1.n114 VDD1.n113 9.3005
R1333 VDD1.n69 VDD1.n68 9.3005
R1334 VDD1.n108 VDD1.n107 9.3005
R1335 VDD1.n81 VDD1.n80 9.3005
R1336 VDD1.n88 VDD1.n87 9.3005
R1337 VDD1.n90 VDD1.n89 9.3005
R1338 VDD1.n77 VDD1.n76 9.3005
R1339 VDD1.n96 VDD1.n95 9.3005
R1340 VDD1.n98 VDD1.n97 9.3005
R1341 VDD1.n99 VDD1.n72 9.3005
R1342 VDD1.n106 VDD1.n105 9.3005
R1343 VDD1.n58 VDD1.n0 8.92171
R1344 VDD1.n29 VDD1.n18 8.92171
R1345 VDD1.n90 VDD1.n79 8.92171
R1346 VDD1.n121 VDD1.n63 8.92171
R1347 VDD1.n26 VDD1.n25 8.14595
R1348 VDD1.n87 VDD1.n86 8.14595
R1349 VDD1.n22 VDD1.n20 7.3702
R1350 VDD1.n83 VDD1.n81 7.3702
R1351 VDD1.n25 VDD1.n20 5.81868
R1352 VDD1.n86 VDD1.n81 5.81868
R1353 VDD1.n60 VDD1.n0 5.04292
R1354 VDD1.n26 VDD1.n18 5.04292
R1355 VDD1.n87 VDD1.n79 5.04292
R1356 VDD1.n123 VDD1.n63 5.04292
R1357 VDD1.n58 VDD1.n57 4.26717
R1358 VDD1.n30 VDD1.n29 4.26717
R1359 VDD1.n91 VDD1.n90 4.26717
R1360 VDD1.n121 VDD1.n120 4.26717
R1361 VDD1.n54 VDD1.n2 3.49141
R1362 VDD1.n33 VDD1.n16 3.49141
R1363 VDD1.n94 VDD1.n77 3.49141
R1364 VDD1.n117 VDD1.n65 3.49141
R1365 VDD1.n21 VDD1.n19 2.84303
R1366 VDD1.n82 VDD1.n80 2.84303
R1367 VDD1.n53 VDD1.n4 2.71565
R1368 VDD1.n34 VDD1.n14 2.71565
R1369 VDD1.n95 VDD1.n75 2.71565
R1370 VDD1.n116 VDD1.n67 2.71565
R1371 VDD1.n50 VDD1.n49 1.93989
R1372 VDD1.n38 VDD1.n37 1.93989
R1373 VDD1.n100 VDD1.n98 1.93989
R1374 VDD1.n113 VDD1.n112 1.93989
R1375 VDD1.n128 VDD1.t0 1.72976
R1376 VDD1.n128 VDD1.t4 1.72976
R1377 VDD1.n61 VDD1.t2 1.72976
R1378 VDD1.n61 VDD1.t3 1.72976
R1379 VDD1.n126 VDD1.t1 1.72976
R1380 VDD1.n126 VDD1.t8 1.72976
R1381 VDD1.n124 VDD1.t5 1.72976
R1382 VDD1.n124 VDD1.t7 1.72976
R1383 VDD1.n46 VDD1.n6 1.16414
R1384 VDD1.n41 VDD1.n11 1.16414
R1385 VDD1.n99 VDD1.n73 1.16414
R1386 VDD1.n109 VDD1.n69 1.16414
R1387 VDD1 VDD1.n129 0.472483
R1388 VDD1.n45 VDD1.n8 0.388379
R1389 VDD1.n42 VDD1.n10 0.388379
R1390 VDD1.n105 VDD1.n104 0.388379
R1391 VDD1.n108 VDD1.n71 0.388379
R1392 VDD1 VDD1.n62 0.235414
R1393 VDD1.n59 VDD1.n1 0.155672
R1394 VDD1.n52 VDD1.n1 0.155672
R1395 VDD1.n52 VDD1.n51 0.155672
R1396 VDD1.n51 VDD1.n5 0.155672
R1397 VDD1.n44 VDD1.n5 0.155672
R1398 VDD1.n44 VDD1.n43 0.155672
R1399 VDD1.n43 VDD1.n9 0.155672
R1400 VDD1.n36 VDD1.n9 0.155672
R1401 VDD1.n36 VDD1.n35 0.155672
R1402 VDD1.n35 VDD1.n15 0.155672
R1403 VDD1.n28 VDD1.n15 0.155672
R1404 VDD1.n28 VDD1.n27 0.155672
R1405 VDD1.n27 VDD1.n19 0.155672
R1406 VDD1.n88 VDD1.n80 0.155672
R1407 VDD1.n89 VDD1.n88 0.155672
R1408 VDD1.n89 VDD1.n76 0.155672
R1409 VDD1.n96 VDD1.n76 0.155672
R1410 VDD1.n97 VDD1.n96 0.155672
R1411 VDD1.n97 VDD1.n72 0.155672
R1412 VDD1.n106 VDD1.n72 0.155672
R1413 VDD1.n107 VDD1.n106 0.155672
R1414 VDD1.n107 VDD1.n68 0.155672
R1415 VDD1.n114 VDD1.n68 0.155672
R1416 VDD1.n115 VDD1.n114 0.155672
R1417 VDD1.n115 VDD1.n64 0.155672
R1418 VDD1.n122 VDD1.n64 0.155672
R1419 VDD1.n127 VDD1.n125 0.121878
R1420 VTAIL.n256 VTAIL.n200 289.615
R1421 VTAIL.n58 VTAIL.n2 289.615
R1422 VTAIL.n194 VTAIL.n138 289.615
R1423 VTAIL.n128 VTAIL.n72 289.615
R1424 VTAIL.n221 VTAIL.n220 185
R1425 VTAIL.n223 VTAIL.n222 185
R1426 VTAIL.n216 VTAIL.n215 185
R1427 VTAIL.n229 VTAIL.n228 185
R1428 VTAIL.n231 VTAIL.n230 185
R1429 VTAIL.n212 VTAIL.n211 185
R1430 VTAIL.n238 VTAIL.n237 185
R1431 VTAIL.n239 VTAIL.n210 185
R1432 VTAIL.n241 VTAIL.n240 185
R1433 VTAIL.n208 VTAIL.n207 185
R1434 VTAIL.n247 VTAIL.n246 185
R1435 VTAIL.n249 VTAIL.n248 185
R1436 VTAIL.n204 VTAIL.n203 185
R1437 VTAIL.n255 VTAIL.n254 185
R1438 VTAIL.n257 VTAIL.n256 185
R1439 VTAIL.n23 VTAIL.n22 185
R1440 VTAIL.n25 VTAIL.n24 185
R1441 VTAIL.n18 VTAIL.n17 185
R1442 VTAIL.n31 VTAIL.n30 185
R1443 VTAIL.n33 VTAIL.n32 185
R1444 VTAIL.n14 VTAIL.n13 185
R1445 VTAIL.n40 VTAIL.n39 185
R1446 VTAIL.n41 VTAIL.n12 185
R1447 VTAIL.n43 VTAIL.n42 185
R1448 VTAIL.n10 VTAIL.n9 185
R1449 VTAIL.n49 VTAIL.n48 185
R1450 VTAIL.n51 VTAIL.n50 185
R1451 VTAIL.n6 VTAIL.n5 185
R1452 VTAIL.n57 VTAIL.n56 185
R1453 VTAIL.n59 VTAIL.n58 185
R1454 VTAIL.n195 VTAIL.n194 185
R1455 VTAIL.n193 VTAIL.n192 185
R1456 VTAIL.n142 VTAIL.n141 185
R1457 VTAIL.n187 VTAIL.n186 185
R1458 VTAIL.n185 VTAIL.n184 185
R1459 VTAIL.n146 VTAIL.n145 185
R1460 VTAIL.n150 VTAIL.n148 185
R1461 VTAIL.n179 VTAIL.n178 185
R1462 VTAIL.n177 VTAIL.n176 185
R1463 VTAIL.n152 VTAIL.n151 185
R1464 VTAIL.n171 VTAIL.n170 185
R1465 VTAIL.n169 VTAIL.n168 185
R1466 VTAIL.n156 VTAIL.n155 185
R1467 VTAIL.n163 VTAIL.n162 185
R1468 VTAIL.n161 VTAIL.n160 185
R1469 VTAIL.n129 VTAIL.n128 185
R1470 VTAIL.n127 VTAIL.n126 185
R1471 VTAIL.n76 VTAIL.n75 185
R1472 VTAIL.n121 VTAIL.n120 185
R1473 VTAIL.n119 VTAIL.n118 185
R1474 VTAIL.n80 VTAIL.n79 185
R1475 VTAIL.n84 VTAIL.n82 185
R1476 VTAIL.n113 VTAIL.n112 185
R1477 VTAIL.n111 VTAIL.n110 185
R1478 VTAIL.n86 VTAIL.n85 185
R1479 VTAIL.n105 VTAIL.n104 185
R1480 VTAIL.n103 VTAIL.n102 185
R1481 VTAIL.n90 VTAIL.n89 185
R1482 VTAIL.n97 VTAIL.n96 185
R1483 VTAIL.n95 VTAIL.n94 185
R1484 VTAIL.n219 VTAIL.t7 149.524
R1485 VTAIL.n21 VTAIL.t15 149.524
R1486 VTAIL.n159 VTAIL.t13 149.524
R1487 VTAIL.n93 VTAIL.t4 149.524
R1488 VTAIL.n222 VTAIL.n221 104.615
R1489 VTAIL.n222 VTAIL.n215 104.615
R1490 VTAIL.n229 VTAIL.n215 104.615
R1491 VTAIL.n230 VTAIL.n229 104.615
R1492 VTAIL.n230 VTAIL.n211 104.615
R1493 VTAIL.n238 VTAIL.n211 104.615
R1494 VTAIL.n239 VTAIL.n238 104.615
R1495 VTAIL.n240 VTAIL.n239 104.615
R1496 VTAIL.n240 VTAIL.n207 104.615
R1497 VTAIL.n247 VTAIL.n207 104.615
R1498 VTAIL.n248 VTAIL.n247 104.615
R1499 VTAIL.n248 VTAIL.n203 104.615
R1500 VTAIL.n255 VTAIL.n203 104.615
R1501 VTAIL.n256 VTAIL.n255 104.615
R1502 VTAIL.n24 VTAIL.n23 104.615
R1503 VTAIL.n24 VTAIL.n17 104.615
R1504 VTAIL.n31 VTAIL.n17 104.615
R1505 VTAIL.n32 VTAIL.n31 104.615
R1506 VTAIL.n32 VTAIL.n13 104.615
R1507 VTAIL.n40 VTAIL.n13 104.615
R1508 VTAIL.n41 VTAIL.n40 104.615
R1509 VTAIL.n42 VTAIL.n41 104.615
R1510 VTAIL.n42 VTAIL.n9 104.615
R1511 VTAIL.n49 VTAIL.n9 104.615
R1512 VTAIL.n50 VTAIL.n49 104.615
R1513 VTAIL.n50 VTAIL.n5 104.615
R1514 VTAIL.n57 VTAIL.n5 104.615
R1515 VTAIL.n58 VTAIL.n57 104.615
R1516 VTAIL.n194 VTAIL.n193 104.615
R1517 VTAIL.n193 VTAIL.n141 104.615
R1518 VTAIL.n186 VTAIL.n141 104.615
R1519 VTAIL.n186 VTAIL.n185 104.615
R1520 VTAIL.n185 VTAIL.n145 104.615
R1521 VTAIL.n150 VTAIL.n145 104.615
R1522 VTAIL.n178 VTAIL.n150 104.615
R1523 VTAIL.n178 VTAIL.n177 104.615
R1524 VTAIL.n177 VTAIL.n151 104.615
R1525 VTAIL.n170 VTAIL.n151 104.615
R1526 VTAIL.n170 VTAIL.n169 104.615
R1527 VTAIL.n169 VTAIL.n155 104.615
R1528 VTAIL.n162 VTAIL.n155 104.615
R1529 VTAIL.n162 VTAIL.n161 104.615
R1530 VTAIL.n128 VTAIL.n127 104.615
R1531 VTAIL.n127 VTAIL.n75 104.615
R1532 VTAIL.n120 VTAIL.n75 104.615
R1533 VTAIL.n120 VTAIL.n119 104.615
R1534 VTAIL.n119 VTAIL.n79 104.615
R1535 VTAIL.n84 VTAIL.n79 104.615
R1536 VTAIL.n112 VTAIL.n84 104.615
R1537 VTAIL.n112 VTAIL.n111 104.615
R1538 VTAIL.n111 VTAIL.n85 104.615
R1539 VTAIL.n104 VTAIL.n85 104.615
R1540 VTAIL.n104 VTAIL.n103 104.615
R1541 VTAIL.n103 VTAIL.n89 104.615
R1542 VTAIL.n96 VTAIL.n89 104.615
R1543 VTAIL.n96 VTAIL.n95 104.615
R1544 VTAIL.n221 VTAIL.t7 52.3082
R1545 VTAIL.n23 VTAIL.t15 52.3082
R1546 VTAIL.n161 VTAIL.t13 52.3082
R1547 VTAIL.n95 VTAIL.t4 52.3082
R1548 VTAIL.n137 VTAIL.n136 46.3808
R1549 VTAIL.n135 VTAIL.n134 46.3808
R1550 VTAIL.n71 VTAIL.n70 46.3808
R1551 VTAIL.n69 VTAIL.n68 46.3808
R1552 VTAIL.n263 VTAIL.n262 46.3806
R1553 VTAIL.n1 VTAIL.n0 46.3806
R1554 VTAIL.n65 VTAIL.n64 46.3806
R1555 VTAIL.n67 VTAIL.n66 46.3806
R1556 VTAIL.n261 VTAIL.n260 33.155
R1557 VTAIL.n63 VTAIL.n62 33.155
R1558 VTAIL.n199 VTAIL.n198 33.155
R1559 VTAIL.n133 VTAIL.n132 33.155
R1560 VTAIL.n69 VTAIL.n67 23.6514
R1561 VTAIL.n261 VTAIL.n199 22.9445
R1562 VTAIL.n241 VTAIL.n208 13.1884
R1563 VTAIL.n43 VTAIL.n10 13.1884
R1564 VTAIL.n148 VTAIL.n146 13.1884
R1565 VTAIL.n82 VTAIL.n80 13.1884
R1566 VTAIL.n242 VTAIL.n210 12.8005
R1567 VTAIL.n246 VTAIL.n245 12.8005
R1568 VTAIL.n44 VTAIL.n12 12.8005
R1569 VTAIL.n48 VTAIL.n47 12.8005
R1570 VTAIL.n184 VTAIL.n183 12.8005
R1571 VTAIL.n180 VTAIL.n179 12.8005
R1572 VTAIL.n118 VTAIL.n117 12.8005
R1573 VTAIL.n114 VTAIL.n113 12.8005
R1574 VTAIL.n237 VTAIL.n236 12.0247
R1575 VTAIL.n249 VTAIL.n206 12.0247
R1576 VTAIL.n39 VTAIL.n38 12.0247
R1577 VTAIL.n51 VTAIL.n8 12.0247
R1578 VTAIL.n187 VTAIL.n144 12.0247
R1579 VTAIL.n176 VTAIL.n149 12.0247
R1580 VTAIL.n121 VTAIL.n78 12.0247
R1581 VTAIL.n110 VTAIL.n83 12.0247
R1582 VTAIL.n235 VTAIL.n212 11.249
R1583 VTAIL.n250 VTAIL.n204 11.249
R1584 VTAIL.n37 VTAIL.n14 11.249
R1585 VTAIL.n52 VTAIL.n6 11.249
R1586 VTAIL.n188 VTAIL.n142 11.249
R1587 VTAIL.n175 VTAIL.n152 11.249
R1588 VTAIL.n122 VTAIL.n76 11.249
R1589 VTAIL.n109 VTAIL.n86 11.249
R1590 VTAIL.n232 VTAIL.n231 10.4732
R1591 VTAIL.n254 VTAIL.n253 10.4732
R1592 VTAIL.n34 VTAIL.n33 10.4732
R1593 VTAIL.n56 VTAIL.n55 10.4732
R1594 VTAIL.n192 VTAIL.n191 10.4732
R1595 VTAIL.n172 VTAIL.n171 10.4732
R1596 VTAIL.n126 VTAIL.n125 10.4732
R1597 VTAIL.n106 VTAIL.n105 10.4732
R1598 VTAIL.n220 VTAIL.n219 10.2747
R1599 VTAIL.n22 VTAIL.n21 10.2747
R1600 VTAIL.n160 VTAIL.n159 10.2747
R1601 VTAIL.n94 VTAIL.n93 10.2747
R1602 VTAIL.n228 VTAIL.n214 9.69747
R1603 VTAIL.n257 VTAIL.n202 9.69747
R1604 VTAIL.n30 VTAIL.n16 9.69747
R1605 VTAIL.n59 VTAIL.n4 9.69747
R1606 VTAIL.n195 VTAIL.n140 9.69747
R1607 VTAIL.n168 VTAIL.n154 9.69747
R1608 VTAIL.n129 VTAIL.n74 9.69747
R1609 VTAIL.n102 VTAIL.n88 9.69747
R1610 VTAIL.n260 VTAIL.n259 9.45567
R1611 VTAIL.n62 VTAIL.n61 9.45567
R1612 VTAIL.n198 VTAIL.n197 9.45567
R1613 VTAIL.n132 VTAIL.n131 9.45567
R1614 VTAIL.n259 VTAIL.n258 9.3005
R1615 VTAIL.n202 VTAIL.n201 9.3005
R1616 VTAIL.n253 VTAIL.n252 9.3005
R1617 VTAIL.n251 VTAIL.n250 9.3005
R1618 VTAIL.n206 VTAIL.n205 9.3005
R1619 VTAIL.n245 VTAIL.n244 9.3005
R1620 VTAIL.n218 VTAIL.n217 9.3005
R1621 VTAIL.n225 VTAIL.n224 9.3005
R1622 VTAIL.n227 VTAIL.n226 9.3005
R1623 VTAIL.n214 VTAIL.n213 9.3005
R1624 VTAIL.n233 VTAIL.n232 9.3005
R1625 VTAIL.n235 VTAIL.n234 9.3005
R1626 VTAIL.n236 VTAIL.n209 9.3005
R1627 VTAIL.n243 VTAIL.n242 9.3005
R1628 VTAIL.n61 VTAIL.n60 9.3005
R1629 VTAIL.n4 VTAIL.n3 9.3005
R1630 VTAIL.n55 VTAIL.n54 9.3005
R1631 VTAIL.n53 VTAIL.n52 9.3005
R1632 VTAIL.n8 VTAIL.n7 9.3005
R1633 VTAIL.n47 VTAIL.n46 9.3005
R1634 VTAIL.n20 VTAIL.n19 9.3005
R1635 VTAIL.n27 VTAIL.n26 9.3005
R1636 VTAIL.n29 VTAIL.n28 9.3005
R1637 VTAIL.n16 VTAIL.n15 9.3005
R1638 VTAIL.n35 VTAIL.n34 9.3005
R1639 VTAIL.n37 VTAIL.n36 9.3005
R1640 VTAIL.n38 VTAIL.n11 9.3005
R1641 VTAIL.n45 VTAIL.n44 9.3005
R1642 VTAIL.n158 VTAIL.n157 9.3005
R1643 VTAIL.n165 VTAIL.n164 9.3005
R1644 VTAIL.n167 VTAIL.n166 9.3005
R1645 VTAIL.n154 VTAIL.n153 9.3005
R1646 VTAIL.n173 VTAIL.n172 9.3005
R1647 VTAIL.n175 VTAIL.n174 9.3005
R1648 VTAIL.n149 VTAIL.n147 9.3005
R1649 VTAIL.n181 VTAIL.n180 9.3005
R1650 VTAIL.n197 VTAIL.n196 9.3005
R1651 VTAIL.n140 VTAIL.n139 9.3005
R1652 VTAIL.n191 VTAIL.n190 9.3005
R1653 VTAIL.n189 VTAIL.n188 9.3005
R1654 VTAIL.n144 VTAIL.n143 9.3005
R1655 VTAIL.n183 VTAIL.n182 9.3005
R1656 VTAIL.n92 VTAIL.n91 9.3005
R1657 VTAIL.n99 VTAIL.n98 9.3005
R1658 VTAIL.n101 VTAIL.n100 9.3005
R1659 VTAIL.n88 VTAIL.n87 9.3005
R1660 VTAIL.n107 VTAIL.n106 9.3005
R1661 VTAIL.n109 VTAIL.n108 9.3005
R1662 VTAIL.n83 VTAIL.n81 9.3005
R1663 VTAIL.n115 VTAIL.n114 9.3005
R1664 VTAIL.n131 VTAIL.n130 9.3005
R1665 VTAIL.n74 VTAIL.n73 9.3005
R1666 VTAIL.n125 VTAIL.n124 9.3005
R1667 VTAIL.n123 VTAIL.n122 9.3005
R1668 VTAIL.n78 VTAIL.n77 9.3005
R1669 VTAIL.n117 VTAIL.n116 9.3005
R1670 VTAIL.n227 VTAIL.n216 8.92171
R1671 VTAIL.n258 VTAIL.n200 8.92171
R1672 VTAIL.n29 VTAIL.n18 8.92171
R1673 VTAIL.n60 VTAIL.n2 8.92171
R1674 VTAIL.n196 VTAIL.n138 8.92171
R1675 VTAIL.n167 VTAIL.n156 8.92171
R1676 VTAIL.n130 VTAIL.n72 8.92171
R1677 VTAIL.n101 VTAIL.n90 8.92171
R1678 VTAIL.n224 VTAIL.n223 8.14595
R1679 VTAIL.n26 VTAIL.n25 8.14595
R1680 VTAIL.n164 VTAIL.n163 8.14595
R1681 VTAIL.n98 VTAIL.n97 8.14595
R1682 VTAIL.n220 VTAIL.n218 7.3702
R1683 VTAIL.n22 VTAIL.n20 7.3702
R1684 VTAIL.n160 VTAIL.n158 7.3702
R1685 VTAIL.n94 VTAIL.n92 7.3702
R1686 VTAIL.n223 VTAIL.n218 5.81868
R1687 VTAIL.n25 VTAIL.n20 5.81868
R1688 VTAIL.n163 VTAIL.n158 5.81868
R1689 VTAIL.n97 VTAIL.n92 5.81868
R1690 VTAIL.n224 VTAIL.n216 5.04292
R1691 VTAIL.n260 VTAIL.n200 5.04292
R1692 VTAIL.n26 VTAIL.n18 5.04292
R1693 VTAIL.n62 VTAIL.n2 5.04292
R1694 VTAIL.n198 VTAIL.n138 5.04292
R1695 VTAIL.n164 VTAIL.n156 5.04292
R1696 VTAIL.n132 VTAIL.n72 5.04292
R1697 VTAIL.n98 VTAIL.n90 5.04292
R1698 VTAIL.n228 VTAIL.n227 4.26717
R1699 VTAIL.n258 VTAIL.n257 4.26717
R1700 VTAIL.n30 VTAIL.n29 4.26717
R1701 VTAIL.n60 VTAIL.n59 4.26717
R1702 VTAIL.n196 VTAIL.n195 4.26717
R1703 VTAIL.n168 VTAIL.n167 4.26717
R1704 VTAIL.n130 VTAIL.n129 4.26717
R1705 VTAIL.n102 VTAIL.n101 4.26717
R1706 VTAIL.n231 VTAIL.n214 3.49141
R1707 VTAIL.n254 VTAIL.n202 3.49141
R1708 VTAIL.n33 VTAIL.n16 3.49141
R1709 VTAIL.n56 VTAIL.n4 3.49141
R1710 VTAIL.n192 VTAIL.n140 3.49141
R1711 VTAIL.n171 VTAIL.n154 3.49141
R1712 VTAIL.n126 VTAIL.n74 3.49141
R1713 VTAIL.n105 VTAIL.n88 3.49141
R1714 VTAIL.n219 VTAIL.n217 2.84303
R1715 VTAIL.n21 VTAIL.n19 2.84303
R1716 VTAIL.n159 VTAIL.n157 2.84303
R1717 VTAIL.n93 VTAIL.n91 2.84303
R1718 VTAIL.n232 VTAIL.n212 2.71565
R1719 VTAIL.n253 VTAIL.n204 2.71565
R1720 VTAIL.n34 VTAIL.n14 2.71565
R1721 VTAIL.n55 VTAIL.n6 2.71565
R1722 VTAIL.n191 VTAIL.n142 2.71565
R1723 VTAIL.n172 VTAIL.n152 2.71565
R1724 VTAIL.n125 VTAIL.n76 2.71565
R1725 VTAIL.n106 VTAIL.n86 2.71565
R1726 VTAIL.n237 VTAIL.n235 1.93989
R1727 VTAIL.n250 VTAIL.n249 1.93989
R1728 VTAIL.n39 VTAIL.n37 1.93989
R1729 VTAIL.n52 VTAIL.n51 1.93989
R1730 VTAIL.n188 VTAIL.n187 1.93989
R1731 VTAIL.n176 VTAIL.n175 1.93989
R1732 VTAIL.n122 VTAIL.n121 1.93989
R1733 VTAIL.n110 VTAIL.n109 1.93989
R1734 VTAIL.n262 VTAIL.t3 1.72976
R1735 VTAIL.n262 VTAIL.t2 1.72976
R1736 VTAIL.n0 VTAIL.t6 1.72976
R1737 VTAIL.n0 VTAIL.t19 1.72976
R1738 VTAIL.n64 VTAIL.t16 1.72976
R1739 VTAIL.n64 VTAIL.t17 1.72976
R1740 VTAIL.n66 VTAIL.t10 1.72976
R1741 VTAIL.n66 VTAIL.t14 1.72976
R1742 VTAIL.n136 VTAIL.t12 1.72976
R1743 VTAIL.n136 VTAIL.t9 1.72976
R1744 VTAIL.n134 VTAIL.t11 1.72976
R1745 VTAIL.n134 VTAIL.t8 1.72976
R1746 VTAIL.n70 VTAIL.t1 1.72976
R1747 VTAIL.n70 VTAIL.t0 1.72976
R1748 VTAIL.n68 VTAIL.t5 1.72976
R1749 VTAIL.n68 VTAIL.t18 1.72976
R1750 VTAIL.n236 VTAIL.n210 1.16414
R1751 VTAIL.n246 VTAIL.n206 1.16414
R1752 VTAIL.n38 VTAIL.n12 1.16414
R1753 VTAIL.n48 VTAIL.n8 1.16414
R1754 VTAIL.n184 VTAIL.n144 1.16414
R1755 VTAIL.n179 VTAIL.n149 1.16414
R1756 VTAIL.n118 VTAIL.n78 1.16414
R1757 VTAIL.n113 VTAIL.n83 1.16414
R1758 VTAIL.n135 VTAIL.n133 0.823776
R1759 VTAIL.n63 VTAIL.n1 0.823776
R1760 VTAIL.n71 VTAIL.n69 0.707397
R1761 VTAIL.n133 VTAIL.n71 0.707397
R1762 VTAIL.n137 VTAIL.n135 0.707397
R1763 VTAIL.n199 VTAIL.n137 0.707397
R1764 VTAIL.n67 VTAIL.n65 0.707397
R1765 VTAIL.n65 VTAIL.n63 0.707397
R1766 VTAIL.n263 VTAIL.n261 0.707397
R1767 VTAIL VTAIL.n1 0.588862
R1768 VTAIL.n242 VTAIL.n241 0.388379
R1769 VTAIL.n245 VTAIL.n208 0.388379
R1770 VTAIL.n44 VTAIL.n43 0.388379
R1771 VTAIL.n47 VTAIL.n10 0.388379
R1772 VTAIL.n183 VTAIL.n146 0.388379
R1773 VTAIL.n180 VTAIL.n148 0.388379
R1774 VTAIL.n117 VTAIL.n80 0.388379
R1775 VTAIL.n114 VTAIL.n82 0.388379
R1776 VTAIL.n225 VTAIL.n217 0.155672
R1777 VTAIL.n226 VTAIL.n225 0.155672
R1778 VTAIL.n226 VTAIL.n213 0.155672
R1779 VTAIL.n233 VTAIL.n213 0.155672
R1780 VTAIL.n234 VTAIL.n233 0.155672
R1781 VTAIL.n234 VTAIL.n209 0.155672
R1782 VTAIL.n243 VTAIL.n209 0.155672
R1783 VTAIL.n244 VTAIL.n243 0.155672
R1784 VTAIL.n244 VTAIL.n205 0.155672
R1785 VTAIL.n251 VTAIL.n205 0.155672
R1786 VTAIL.n252 VTAIL.n251 0.155672
R1787 VTAIL.n252 VTAIL.n201 0.155672
R1788 VTAIL.n259 VTAIL.n201 0.155672
R1789 VTAIL.n27 VTAIL.n19 0.155672
R1790 VTAIL.n28 VTAIL.n27 0.155672
R1791 VTAIL.n28 VTAIL.n15 0.155672
R1792 VTAIL.n35 VTAIL.n15 0.155672
R1793 VTAIL.n36 VTAIL.n35 0.155672
R1794 VTAIL.n36 VTAIL.n11 0.155672
R1795 VTAIL.n45 VTAIL.n11 0.155672
R1796 VTAIL.n46 VTAIL.n45 0.155672
R1797 VTAIL.n46 VTAIL.n7 0.155672
R1798 VTAIL.n53 VTAIL.n7 0.155672
R1799 VTAIL.n54 VTAIL.n53 0.155672
R1800 VTAIL.n54 VTAIL.n3 0.155672
R1801 VTAIL.n61 VTAIL.n3 0.155672
R1802 VTAIL.n197 VTAIL.n139 0.155672
R1803 VTAIL.n190 VTAIL.n139 0.155672
R1804 VTAIL.n190 VTAIL.n189 0.155672
R1805 VTAIL.n189 VTAIL.n143 0.155672
R1806 VTAIL.n182 VTAIL.n143 0.155672
R1807 VTAIL.n182 VTAIL.n181 0.155672
R1808 VTAIL.n181 VTAIL.n147 0.155672
R1809 VTAIL.n174 VTAIL.n147 0.155672
R1810 VTAIL.n174 VTAIL.n173 0.155672
R1811 VTAIL.n173 VTAIL.n153 0.155672
R1812 VTAIL.n166 VTAIL.n153 0.155672
R1813 VTAIL.n166 VTAIL.n165 0.155672
R1814 VTAIL.n165 VTAIL.n157 0.155672
R1815 VTAIL.n131 VTAIL.n73 0.155672
R1816 VTAIL.n124 VTAIL.n73 0.155672
R1817 VTAIL.n124 VTAIL.n123 0.155672
R1818 VTAIL.n123 VTAIL.n77 0.155672
R1819 VTAIL.n116 VTAIL.n77 0.155672
R1820 VTAIL.n116 VTAIL.n115 0.155672
R1821 VTAIL.n115 VTAIL.n81 0.155672
R1822 VTAIL.n108 VTAIL.n81 0.155672
R1823 VTAIL.n108 VTAIL.n107 0.155672
R1824 VTAIL.n107 VTAIL.n87 0.155672
R1825 VTAIL.n100 VTAIL.n87 0.155672
R1826 VTAIL.n100 VTAIL.n99 0.155672
R1827 VTAIL.n99 VTAIL.n91 0.155672
R1828 VTAIL VTAIL.n263 0.119034
R1829 VN.n2 VN.t2 664.797
R1830 VN.n14 VN.t4 664.797
R1831 VN.n3 VN.t9 643.814
R1832 VN.n1 VN.t0 643.814
R1833 VN.n9 VN.t1 643.814
R1834 VN.n10 VN.t7 643.814
R1835 VN.n15 VN.t8 643.814
R1836 VN.n13 VN.t3 643.814
R1837 VN.n21 VN.t6 643.814
R1838 VN.n22 VN.t5 643.814
R1839 VN.n11 VN.n10 161.3
R1840 VN.n23 VN.n22 161.3
R1841 VN.n21 VN.n12 161.3
R1842 VN.n20 VN.n19 161.3
R1843 VN.n18 VN.n13 161.3
R1844 VN.n17 VN.n16 161.3
R1845 VN.n9 VN.n0 161.3
R1846 VN.n8 VN.n7 161.3
R1847 VN.n6 VN.n1 161.3
R1848 VN.n5 VN.n4 161.3
R1849 VN.n17 VN.n14 70.4033
R1850 VN.n5 VN.n2 70.4033
R1851 VN.n10 VN.n9 48.2005
R1852 VN.n22 VN.n21 48.2005
R1853 VN VN.n23 41.616
R1854 VN.n4 VN.n1 37.246
R1855 VN.n8 VN.n1 37.246
R1856 VN.n16 VN.n13 37.246
R1857 VN.n20 VN.n13 37.246
R1858 VN.n15 VN.n14 20.9576
R1859 VN.n3 VN.n2 20.9576
R1860 VN.n4 VN.n3 10.955
R1861 VN.n9 VN.n8 10.955
R1862 VN.n16 VN.n15 10.955
R1863 VN.n21 VN.n20 10.955
R1864 VN.n23 VN.n12 0.189894
R1865 VN.n19 VN.n12 0.189894
R1866 VN.n19 VN.n18 0.189894
R1867 VN.n18 VN.n17 0.189894
R1868 VN.n6 VN.n5 0.189894
R1869 VN.n7 VN.n6 0.189894
R1870 VN.n7 VN.n0 0.189894
R1871 VN.n11 VN.n0 0.189894
R1872 VN VN.n11 0.0516364
R1873 VDD2.n121 VDD2.n65 289.615
R1874 VDD2.n56 VDD2.n0 289.615
R1875 VDD2.n122 VDD2.n121 185
R1876 VDD2.n120 VDD2.n119 185
R1877 VDD2.n69 VDD2.n68 185
R1878 VDD2.n114 VDD2.n113 185
R1879 VDD2.n112 VDD2.n111 185
R1880 VDD2.n73 VDD2.n72 185
R1881 VDD2.n77 VDD2.n75 185
R1882 VDD2.n106 VDD2.n105 185
R1883 VDD2.n104 VDD2.n103 185
R1884 VDD2.n79 VDD2.n78 185
R1885 VDD2.n98 VDD2.n97 185
R1886 VDD2.n96 VDD2.n95 185
R1887 VDD2.n83 VDD2.n82 185
R1888 VDD2.n90 VDD2.n89 185
R1889 VDD2.n88 VDD2.n87 185
R1890 VDD2.n21 VDD2.n20 185
R1891 VDD2.n23 VDD2.n22 185
R1892 VDD2.n16 VDD2.n15 185
R1893 VDD2.n29 VDD2.n28 185
R1894 VDD2.n31 VDD2.n30 185
R1895 VDD2.n12 VDD2.n11 185
R1896 VDD2.n38 VDD2.n37 185
R1897 VDD2.n39 VDD2.n10 185
R1898 VDD2.n41 VDD2.n40 185
R1899 VDD2.n8 VDD2.n7 185
R1900 VDD2.n47 VDD2.n46 185
R1901 VDD2.n49 VDD2.n48 185
R1902 VDD2.n4 VDD2.n3 185
R1903 VDD2.n55 VDD2.n54 185
R1904 VDD2.n57 VDD2.n56 185
R1905 VDD2.n86 VDD2.t4 149.524
R1906 VDD2.n19 VDD2.t7 149.524
R1907 VDD2.n121 VDD2.n120 104.615
R1908 VDD2.n120 VDD2.n68 104.615
R1909 VDD2.n113 VDD2.n68 104.615
R1910 VDD2.n113 VDD2.n112 104.615
R1911 VDD2.n112 VDD2.n72 104.615
R1912 VDD2.n77 VDD2.n72 104.615
R1913 VDD2.n105 VDD2.n77 104.615
R1914 VDD2.n105 VDD2.n104 104.615
R1915 VDD2.n104 VDD2.n78 104.615
R1916 VDD2.n97 VDD2.n78 104.615
R1917 VDD2.n97 VDD2.n96 104.615
R1918 VDD2.n96 VDD2.n82 104.615
R1919 VDD2.n89 VDD2.n82 104.615
R1920 VDD2.n89 VDD2.n88 104.615
R1921 VDD2.n22 VDD2.n21 104.615
R1922 VDD2.n22 VDD2.n15 104.615
R1923 VDD2.n29 VDD2.n15 104.615
R1924 VDD2.n30 VDD2.n29 104.615
R1925 VDD2.n30 VDD2.n11 104.615
R1926 VDD2.n38 VDD2.n11 104.615
R1927 VDD2.n39 VDD2.n38 104.615
R1928 VDD2.n40 VDD2.n39 104.615
R1929 VDD2.n40 VDD2.n7 104.615
R1930 VDD2.n47 VDD2.n7 104.615
R1931 VDD2.n48 VDD2.n47 104.615
R1932 VDD2.n48 VDD2.n3 104.615
R1933 VDD2.n55 VDD2.n3 104.615
R1934 VDD2.n56 VDD2.n55 104.615
R1935 VDD2.n64 VDD2.n63 63.5342
R1936 VDD2 VDD2.n129 63.5314
R1937 VDD2.n128 VDD2.n127 63.0596
R1938 VDD2.n62 VDD2.n61 63.0594
R1939 VDD2.n88 VDD2.t4 52.3082
R1940 VDD2.n21 VDD2.t7 52.3082
R1941 VDD2.n62 VDD2.n60 50.5407
R1942 VDD2.n126 VDD2.n125 49.8338
R1943 VDD2.n126 VDD2.n64 36.9437
R1944 VDD2.n75 VDD2.n73 13.1884
R1945 VDD2.n41 VDD2.n8 13.1884
R1946 VDD2.n111 VDD2.n110 12.8005
R1947 VDD2.n107 VDD2.n106 12.8005
R1948 VDD2.n42 VDD2.n10 12.8005
R1949 VDD2.n46 VDD2.n45 12.8005
R1950 VDD2.n114 VDD2.n71 12.0247
R1951 VDD2.n103 VDD2.n76 12.0247
R1952 VDD2.n37 VDD2.n36 12.0247
R1953 VDD2.n49 VDD2.n6 12.0247
R1954 VDD2.n115 VDD2.n69 11.249
R1955 VDD2.n102 VDD2.n79 11.249
R1956 VDD2.n35 VDD2.n12 11.249
R1957 VDD2.n50 VDD2.n4 11.249
R1958 VDD2.n119 VDD2.n118 10.4732
R1959 VDD2.n99 VDD2.n98 10.4732
R1960 VDD2.n32 VDD2.n31 10.4732
R1961 VDD2.n54 VDD2.n53 10.4732
R1962 VDD2.n87 VDD2.n86 10.2747
R1963 VDD2.n20 VDD2.n19 10.2747
R1964 VDD2.n122 VDD2.n67 9.69747
R1965 VDD2.n95 VDD2.n81 9.69747
R1966 VDD2.n28 VDD2.n14 9.69747
R1967 VDD2.n57 VDD2.n2 9.69747
R1968 VDD2.n125 VDD2.n124 9.45567
R1969 VDD2.n60 VDD2.n59 9.45567
R1970 VDD2.n85 VDD2.n84 9.3005
R1971 VDD2.n92 VDD2.n91 9.3005
R1972 VDD2.n94 VDD2.n93 9.3005
R1973 VDD2.n81 VDD2.n80 9.3005
R1974 VDD2.n100 VDD2.n99 9.3005
R1975 VDD2.n102 VDD2.n101 9.3005
R1976 VDD2.n76 VDD2.n74 9.3005
R1977 VDD2.n108 VDD2.n107 9.3005
R1978 VDD2.n124 VDD2.n123 9.3005
R1979 VDD2.n67 VDD2.n66 9.3005
R1980 VDD2.n118 VDD2.n117 9.3005
R1981 VDD2.n116 VDD2.n115 9.3005
R1982 VDD2.n71 VDD2.n70 9.3005
R1983 VDD2.n110 VDD2.n109 9.3005
R1984 VDD2.n59 VDD2.n58 9.3005
R1985 VDD2.n2 VDD2.n1 9.3005
R1986 VDD2.n53 VDD2.n52 9.3005
R1987 VDD2.n51 VDD2.n50 9.3005
R1988 VDD2.n6 VDD2.n5 9.3005
R1989 VDD2.n45 VDD2.n44 9.3005
R1990 VDD2.n18 VDD2.n17 9.3005
R1991 VDD2.n25 VDD2.n24 9.3005
R1992 VDD2.n27 VDD2.n26 9.3005
R1993 VDD2.n14 VDD2.n13 9.3005
R1994 VDD2.n33 VDD2.n32 9.3005
R1995 VDD2.n35 VDD2.n34 9.3005
R1996 VDD2.n36 VDD2.n9 9.3005
R1997 VDD2.n43 VDD2.n42 9.3005
R1998 VDD2.n123 VDD2.n65 8.92171
R1999 VDD2.n94 VDD2.n83 8.92171
R2000 VDD2.n27 VDD2.n16 8.92171
R2001 VDD2.n58 VDD2.n0 8.92171
R2002 VDD2.n91 VDD2.n90 8.14595
R2003 VDD2.n24 VDD2.n23 8.14595
R2004 VDD2.n87 VDD2.n85 7.3702
R2005 VDD2.n20 VDD2.n18 7.3702
R2006 VDD2.n90 VDD2.n85 5.81868
R2007 VDD2.n23 VDD2.n18 5.81868
R2008 VDD2.n125 VDD2.n65 5.04292
R2009 VDD2.n91 VDD2.n83 5.04292
R2010 VDD2.n24 VDD2.n16 5.04292
R2011 VDD2.n60 VDD2.n0 5.04292
R2012 VDD2.n123 VDD2.n122 4.26717
R2013 VDD2.n95 VDD2.n94 4.26717
R2014 VDD2.n28 VDD2.n27 4.26717
R2015 VDD2.n58 VDD2.n57 4.26717
R2016 VDD2.n119 VDD2.n67 3.49141
R2017 VDD2.n98 VDD2.n81 3.49141
R2018 VDD2.n31 VDD2.n14 3.49141
R2019 VDD2.n54 VDD2.n2 3.49141
R2020 VDD2.n86 VDD2.n84 2.84303
R2021 VDD2.n19 VDD2.n17 2.84303
R2022 VDD2.n118 VDD2.n69 2.71565
R2023 VDD2.n99 VDD2.n79 2.71565
R2024 VDD2.n32 VDD2.n12 2.71565
R2025 VDD2.n53 VDD2.n4 2.71565
R2026 VDD2.n115 VDD2.n114 1.93989
R2027 VDD2.n103 VDD2.n102 1.93989
R2028 VDD2.n37 VDD2.n35 1.93989
R2029 VDD2.n50 VDD2.n49 1.93989
R2030 VDD2.n129 VDD2.t1 1.72976
R2031 VDD2.n129 VDD2.t5 1.72976
R2032 VDD2.n127 VDD2.t3 1.72976
R2033 VDD2.n127 VDD2.t6 1.72976
R2034 VDD2.n63 VDD2.t8 1.72976
R2035 VDD2.n63 VDD2.t2 1.72976
R2036 VDD2.n61 VDD2.t0 1.72976
R2037 VDD2.n61 VDD2.t9 1.72976
R2038 VDD2.n111 VDD2.n71 1.16414
R2039 VDD2.n106 VDD2.n76 1.16414
R2040 VDD2.n36 VDD2.n10 1.16414
R2041 VDD2.n46 VDD2.n6 1.16414
R2042 VDD2.n128 VDD2.n126 0.707397
R2043 VDD2.n110 VDD2.n73 0.388379
R2044 VDD2.n107 VDD2.n75 0.388379
R2045 VDD2.n42 VDD2.n41 0.388379
R2046 VDD2.n45 VDD2.n8 0.388379
R2047 VDD2 VDD2.n128 0.235414
R2048 VDD2.n124 VDD2.n66 0.155672
R2049 VDD2.n117 VDD2.n66 0.155672
R2050 VDD2.n117 VDD2.n116 0.155672
R2051 VDD2.n116 VDD2.n70 0.155672
R2052 VDD2.n109 VDD2.n70 0.155672
R2053 VDD2.n109 VDD2.n108 0.155672
R2054 VDD2.n108 VDD2.n74 0.155672
R2055 VDD2.n101 VDD2.n74 0.155672
R2056 VDD2.n101 VDD2.n100 0.155672
R2057 VDD2.n100 VDD2.n80 0.155672
R2058 VDD2.n93 VDD2.n80 0.155672
R2059 VDD2.n93 VDD2.n92 0.155672
R2060 VDD2.n92 VDD2.n84 0.155672
R2061 VDD2.n25 VDD2.n17 0.155672
R2062 VDD2.n26 VDD2.n25 0.155672
R2063 VDD2.n26 VDD2.n13 0.155672
R2064 VDD2.n33 VDD2.n13 0.155672
R2065 VDD2.n34 VDD2.n33 0.155672
R2066 VDD2.n34 VDD2.n9 0.155672
R2067 VDD2.n43 VDD2.n9 0.155672
R2068 VDD2.n44 VDD2.n43 0.155672
R2069 VDD2.n44 VDD2.n5 0.155672
R2070 VDD2.n51 VDD2.n5 0.155672
R2071 VDD2.n52 VDD2.n51 0.155672
R2072 VDD2.n52 VDD2.n1 0.155672
R2073 VDD2.n59 VDD2.n1 0.155672
R2074 VDD2.n64 VDD2.n62 0.121878
C0 VDD2 VDD1 0.841757f
C1 VDD1 VP 5.3832f
C2 VDD2 VN 5.22169f
C3 VDD1 VTAIL 16.039598f
C4 VP VN 5.18731f
C5 VDD2 VP 0.31479f
C6 VTAIL VN 4.96208f
C7 VDD2 VTAIL 16.0718f
C8 VP VTAIL 4.97673f
C9 VDD1 VN 0.148521f
C10 VDD2 B 4.642199f
C11 VDD1 B 4.54203f
C12 VTAIL B 6.101159f
C13 VN B 8.5063f
C14 VP B 6.451479f
C15 VDD2.n0 B 0.037117f
C16 VDD2.n1 B 0.026281f
C17 VDD2.n2 B 0.014122f
C18 VDD2.n3 B 0.03338f
C19 VDD2.n4 B 0.014953f
C20 VDD2.n5 B 0.026281f
C21 VDD2.n6 B 0.014122f
C22 VDD2.n7 B 0.03338f
C23 VDD2.n8 B 0.014538f
C24 VDD2.n9 B 0.026281f
C25 VDD2.n10 B 0.014953f
C26 VDD2.n11 B 0.03338f
C27 VDD2.n12 B 0.014953f
C28 VDD2.n13 B 0.026281f
C29 VDD2.n14 B 0.014122f
C30 VDD2.n15 B 0.03338f
C31 VDD2.n16 B 0.014953f
C32 VDD2.n17 B 1.26153f
C33 VDD2.n18 B 0.014122f
C34 VDD2.t7 B 0.056298f
C35 VDD2.n19 B 0.183932f
C36 VDD2.n20 B 0.023597f
C37 VDD2.n21 B 0.025035f
C38 VDD2.n22 B 0.03338f
C39 VDD2.n23 B 0.014953f
C40 VDD2.n24 B 0.014122f
C41 VDD2.n25 B 0.026281f
C42 VDD2.n26 B 0.026281f
C43 VDD2.n27 B 0.014122f
C44 VDD2.n28 B 0.014953f
C45 VDD2.n29 B 0.03338f
C46 VDD2.n30 B 0.03338f
C47 VDD2.n31 B 0.014953f
C48 VDD2.n32 B 0.014122f
C49 VDD2.n33 B 0.026281f
C50 VDD2.n34 B 0.026281f
C51 VDD2.n35 B 0.014122f
C52 VDD2.n36 B 0.014122f
C53 VDD2.n37 B 0.014953f
C54 VDD2.n38 B 0.03338f
C55 VDD2.n39 B 0.03338f
C56 VDD2.n40 B 0.03338f
C57 VDD2.n41 B 0.014538f
C58 VDD2.n42 B 0.014122f
C59 VDD2.n43 B 0.026281f
C60 VDD2.n44 B 0.026281f
C61 VDD2.n45 B 0.014122f
C62 VDD2.n46 B 0.014953f
C63 VDD2.n47 B 0.03338f
C64 VDD2.n48 B 0.03338f
C65 VDD2.n49 B 0.014953f
C66 VDD2.n50 B 0.014122f
C67 VDD2.n51 B 0.026281f
C68 VDD2.n52 B 0.026281f
C69 VDD2.n53 B 0.014122f
C70 VDD2.n54 B 0.014953f
C71 VDD2.n55 B 0.03338f
C72 VDD2.n56 B 0.072575f
C73 VDD2.n57 B 0.014953f
C74 VDD2.n58 B 0.014122f
C75 VDD2.n59 B 0.062542f
C76 VDD2.n60 B 0.060387f
C77 VDD2.t0 B 0.237792f
C78 VDD2.t9 B 0.237792f
C79 VDD2.n61 B 2.11364f
C80 VDD2.n62 B 0.400951f
C81 VDD2.t8 B 0.237792f
C82 VDD2.t2 B 0.237792f
C83 VDD2.n63 B 2.11609f
C84 VDD2.n64 B 1.84655f
C85 VDD2.n65 B 0.037117f
C86 VDD2.n66 B 0.026281f
C87 VDD2.n67 B 0.014122f
C88 VDD2.n68 B 0.03338f
C89 VDD2.n69 B 0.014953f
C90 VDD2.n70 B 0.026281f
C91 VDD2.n71 B 0.014122f
C92 VDD2.n72 B 0.03338f
C93 VDD2.n73 B 0.014538f
C94 VDD2.n74 B 0.026281f
C95 VDD2.n75 B 0.014538f
C96 VDD2.n76 B 0.014122f
C97 VDD2.n77 B 0.03338f
C98 VDD2.n78 B 0.03338f
C99 VDD2.n79 B 0.014953f
C100 VDD2.n80 B 0.026281f
C101 VDD2.n81 B 0.014122f
C102 VDD2.n82 B 0.03338f
C103 VDD2.n83 B 0.014953f
C104 VDD2.n84 B 1.26153f
C105 VDD2.n85 B 0.014122f
C106 VDD2.t4 B 0.056298f
C107 VDD2.n86 B 0.183933f
C108 VDD2.n87 B 0.023597f
C109 VDD2.n88 B 0.025035f
C110 VDD2.n89 B 0.03338f
C111 VDD2.n90 B 0.014953f
C112 VDD2.n91 B 0.014122f
C113 VDD2.n92 B 0.026281f
C114 VDD2.n93 B 0.026281f
C115 VDD2.n94 B 0.014122f
C116 VDD2.n95 B 0.014953f
C117 VDD2.n96 B 0.03338f
C118 VDD2.n97 B 0.03338f
C119 VDD2.n98 B 0.014953f
C120 VDD2.n99 B 0.014122f
C121 VDD2.n100 B 0.026281f
C122 VDD2.n101 B 0.026281f
C123 VDD2.n102 B 0.014122f
C124 VDD2.n103 B 0.014953f
C125 VDD2.n104 B 0.03338f
C126 VDD2.n105 B 0.03338f
C127 VDD2.n106 B 0.014953f
C128 VDD2.n107 B 0.014122f
C129 VDD2.n108 B 0.026281f
C130 VDD2.n109 B 0.026281f
C131 VDD2.n110 B 0.014122f
C132 VDD2.n111 B 0.014953f
C133 VDD2.n112 B 0.03338f
C134 VDD2.n113 B 0.03338f
C135 VDD2.n114 B 0.014953f
C136 VDD2.n115 B 0.014122f
C137 VDD2.n116 B 0.026281f
C138 VDD2.n117 B 0.026281f
C139 VDD2.n118 B 0.014122f
C140 VDD2.n119 B 0.014953f
C141 VDD2.n120 B 0.03338f
C142 VDD2.n121 B 0.072575f
C143 VDD2.n122 B 0.014953f
C144 VDD2.n123 B 0.014122f
C145 VDD2.n124 B 0.062542f
C146 VDD2.n125 B 0.058827f
C147 VDD2.n126 B 2.1359f
C148 VDD2.t3 B 0.237792f
C149 VDD2.t6 B 0.237792f
C150 VDD2.n127 B 2.11365f
C151 VDD2.n128 B 0.295602f
C152 VDD2.t1 B 0.237792f
C153 VDD2.t5 B 0.237792f
C154 VDD2.n129 B 2.11607f
C155 VN.n0 B 0.047924f
C156 VN.t0 B 0.767556f
C157 VN.n1 B 0.31782f
C158 VN.t2 B 0.777421f
C159 VN.n2 B 0.302981f
C160 VN.t9 B 0.767556f
C161 VN.n3 B 0.314717f
C162 VN.n4 B 0.010875f
C163 VN.n5 B 0.151404f
C164 VN.n6 B 0.047924f
C165 VN.n7 B 0.047924f
C166 VN.n8 B 0.010875f
C167 VN.t1 B 0.767556f
C168 VN.n9 B 0.314717f
C169 VN.t7 B 0.767556f
C170 VN.n10 B 0.312501f
C171 VN.n11 B 0.037139f
C172 VN.n12 B 0.047924f
C173 VN.t3 B 0.767556f
C174 VN.n13 B 0.31782f
C175 VN.t4 B 0.777421f
C176 VN.n14 B 0.302981f
C177 VN.t8 B 0.767556f
C178 VN.n15 B 0.314717f
C179 VN.n16 B 0.010875f
C180 VN.n17 B 0.151404f
C181 VN.n18 B 0.047924f
C182 VN.n19 B 0.047924f
C183 VN.n20 B 0.010875f
C184 VN.t6 B 0.767556f
C185 VN.n21 B 0.314717f
C186 VN.t5 B 0.767556f
C187 VN.n22 B 0.312501f
C188 VN.n23 B 1.94961f
C189 VTAIL.t6 B 0.248466f
C190 VTAIL.t19 B 0.248466f
C191 VTAIL.n0 B 2.12929f
C192 VTAIL.n1 B 0.392356f
C193 VTAIL.n2 B 0.038783f
C194 VTAIL.n3 B 0.027461f
C195 VTAIL.n4 B 0.014756f
C196 VTAIL.n5 B 0.034878f
C197 VTAIL.n6 B 0.015624f
C198 VTAIL.n7 B 0.027461f
C199 VTAIL.n8 B 0.014756f
C200 VTAIL.n9 B 0.034878f
C201 VTAIL.n10 B 0.01519f
C202 VTAIL.n11 B 0.027461f
C203 VTAIL.n12 B 0.015624f
C204 VTAIL.n13 B 0.034878f
C205 VTAIL.n14 B 0.015624f
C206 VTAIL.n15 B 0.027461f
C207 VTAIL.n16 B 0.014756f
C208 VTAIL.n17 B 0.034878f
C209 VTAIL.n18 B 0.015624f
C210 VTAIL.n19 B 1.31815f
C211 VTAIL.n20 B 0.014756f
C212 VTAIL.t15 B 0.058826f
C213 VTAIL.n21 B 0.192189f
C214 VTAIL.n22 B 0.024656f
C215 VTAIL.n23 B 0.026159f
C216 VTAIL.n24 B 0.034878f
C217 VTAIL.n25 B 0.015624f
C218 VTAIL.n26 B 0.014756f
C219 VTAIL.n27 B 0.027461f
C220 VTAIL.n28 B 0.027461f
C221 VTAIL.n29 B 0.014756f
C222 VTAIL.n30 B 0.015624f
C223 VTAIL.n31 B 0.034878f
C224 VTAIL.n32 B 0.034878f
C225 VTAIL.n33 B 0.015624f
C226 VTAIL.n34 B 0.014756f
C227 VTAIL.n35 B 0.027461f
C228 VTAIL.n36 B 0.027461f
C229 VTAIL.n37 B 0.014756f
C230 VTAIL.n38 B 0.014756f
C231 VTAIL.n39 B 0.015624f
C232 VTAIL.n40 B 0.034878f
C233 VTAIL.n41 B 0.034878f
C234 VTAIL.n42 B 0.034878f
C235 VTAIL.n43 B 0.01519f
C236 VTAIL.n44 B 0.014756f
C237 VTAIL.n45 B 0.027461f
C238 VTAIL.n46 B 0.027461f
C239 VTAIL.n47 B 0.014756f
C240 VTAIL.n48 B 0.015624f
C241 VTAIL.n49 B 0.034878f
C242 VTAIL.n50 B 0.034878f
C243 VTAIL.n51 B 0.015624f
C244 VTAIL.n52 B 0.014756f
C245 VTAIL.n53 B 0.027461f
C246 VTAIL.n54 B 0.027461f
C247 VTAIL.n55 B 0.014756f
C248 VTAIL.n56 B 0.015624f
C249 VTAIL.n57 B 0.034878f
C250 VTAIL.n58 B 0.075833f
C251 VTAIL.n59 B 0.015624f
C252 VTAIL.n60 B 0.014756f
C253 VTAIL.n61 B 0.065349f
C254 VTAIL.n62 B 0.042522f
C255 VTAIL.n63 B 0.159908f
C256 VTAIL.t16 B 0.248466f
C257 VTAIL.t17 B 0.248466f
C258 VTAIL.n64 B 2.12929f
C259 VTAIL.n65 B 0.392547f
C260 VTAIL.t10 B 0.248466f
C261 VTAIL.t14 B 0.248466f
C262 VTAIL.n66 B 2.12929f
C263 VTAIL.n67 B 1.70151f
C264 VTAIL.t5 B 0.248466f
C265 VTAIL.t18 B 0.248466f
C266 VTAIL.n68 B 2.1293f
C267 VTAIL.n69 B 1.7015f
C268 VTAIL.t1 B 0.248466f
C269 VTAIL.t0 B 0.248466f
C270 VTAIL.n70 B 2.1293f
C271 VTAIL.n71 B 0.392535f
C272 VTAIL.n72 B 0.038783f
C273 VTAIL.n73 B 0.027461f
C274 VTAIL.n74 B 0.014756f
C275 VTAIL.n75 B 0.034878f
C276 VTAIL.n76 B 0.015624f
C277 VTAIL.n77 B 0.027461f
C278 VTAIL.n78 B 0.014756f
C279 VTAIL.n79 B 0.034878f
C280 VTAIL.n80 B 0.01519f
C281 VTAIL.n81 B 0.027461f
C282 VTAIL.n82 B 0.01519f
C283 VTAIL.n83 B 0.014756f
C284 VTAIL.n84 B 0.034878f
C285 VTAIL.n85 B 0.034878f
C286 VTAIL.n86 B 0.015624f
C287 VTAIL.n87 B 0.027461f
C288 VTAIL.n88 B 0.014756f
C289 VTAIL.n89 B 0.034878f
C290 VTAIL.n90 B 0.015624f
C291 VTAIL.n91 B 1.31815f
C292 VTAIL.n92 B 0.014756f
C293 VTAIL.t4 B 0.058826f
C294 VTAIL.n93 B 0.192189f
C295 VTAIL.n94 B 0.024656f
C296 VTAIL.n95 B 0.026159f
C297 VTAIL.n96 B 0.034878f
C298 VTAIL.n97 B 0.015624f
C299 VTAIL.n98 B 0.014756f
C300 VTAIL.n99 B 0.027461f
C301 VTAIL.n100 B 0.027461f
C302 VTAIL.n101 B 0.014756f
C303 VTAIL.n102 B 0.015624f
C304 VTAIL.n103 B 0.034878f
C305 VTAIL.n104 B 0.034878f
C306 VTAIL.n105 B 0.015624f
C307 VTAIL.n106 B 0.014756f
C308 VTAIL.n107 B 0.027461f
C309 VTAIL.n108 B 0.027461f
C310 VTAIL.n109 B 0.014756f
C311 VTAIL.n110 B 0.015624f
C312 VTAIL.n111 B 0.034878f
C313 VTAIL.n112 B 0.034878f
C314 VTAIL.n113 B 0.015624f
C315 VTAIL.n114 B 0.014756f
C316 VTAIL.n115 B 0.027461f
C317 VTAIL.n116 B 0.027461f
C318 VTAIL.n117 B 0.014756f
C319 VTAIL.n118 B 0.015624f
C320 VTAIL.n119 B 0.034878f
C321 VTAIL.n120 B 0.034878f
C322 VTAIL.n121 B 0.015624f
C323 VTAIL.n122 B 0.014756f
C324 VTAIL.n123 B 0.027461f
C325 VTAIL.n124 B 0.027461f
C326 VTAIL.n125 B 0.014756f
C327 VTAIL.n126 B 0.015624f
C328 VTAIL.n127 B 0.034878f
C329 VTAIL.n128 B 0.075833f
C330 VTAIL.n129 B 0.015624f
C331 VTAIL.n130 B 0.014756f
C332 VTAIL.n131 B 0.065349f
C333 VTAIL.n132 B 0.042522f
C334 VTAIL.n133 B 0.159908f
C335 VTAIL.t11 B 0.248466f
C336 VTAIL.t8 B 0.248466f
C337 VTAIL.n134 B 2.1293f
C338 VTAIL.n135 B 0.402832f
C339 VTAIL.t12 B 0.248466f
C340 VTAIL.t9 B 0.248466f
C341 VTAIL.n136 B 2.1293f
C342 VTAIL.n137 B 0.392535f
C343 VTAIL.n138 B 0.038783f
C344 VTAIL.n139 B 0.027461f
C345 VTAIL.n140 B 0.014756f
C346 VTAIL.n141 B 0.034878f
C347 VTAIL.n142 B 0.015624f
C348 VTAIL.n143 B 0.027461f
C349 VTAIL.n144 B 0.014756f
C350 VTAIL.n145 B 0.034878f
C351 VTAIL.n146 B 0.01519f
C352 VTAIL.n147 B 0.027461f
C353 VTAIL.n148 B 0.01519f
C354 VTAIL.n149 B 0.014756f
C355 VTAIL.n150 B 0.034878f
C356 VTAIL.n151 B 0.034878f
C357 VTAIL.n152 B 0.015624f
C358 VTAIL.n153 B 0.027461f
C359 VTAIL.n154 B 0.014756f
C360 VTAIL.n155 B 0.034878f
C361 VTAIL.n156 B 0.015624f
C362 VTAIL.n157 B 1.31815f
C363 VTAIL.n158 B 0.014756f
C364 VTAIL.t13 B 0.058826f
C365 VTAIL.n159 B 0.192189f
C366 VTAIL.n160 B 0.024656f
C367 VTAIL.n161 B 0.026159f
C368 VTAIL.n162 B 0.034878f
C369 VTAIL.n163 B 0.015624f
C370 VTAIL.n164 B 0.014756f
C371 VTAIL.n165 B 0.027461f
C372 VTAIL.n166 B 0.027461f
C373 VTAIL.n167 B 0.014756f
C374 VTAIL.n168 B 0.015624f
C375 VTAIL.n169 B 0.034878f
C376 VTAIL.n170 B 0.034878f
C377 VTAIL.n171 B 0.015624f
C378 VTAIL.n172 B 0.014756f
C379 VTAIL.n173 B 0.027461f
C380 VTAIL.n174 B 0.027461f
C381 VTAIL.n175 B 0.014756f
C382 VTAIL.n176 B 0.015624f
C383 VTAIL.n177 B 0.034878f
C384 VTAIL.n178 B 0.034878f
C385 VTAIL.n179 B 0.015624f
C386 VTAIL.n180 B 0.014756f
C387 VTAIL.n181 B 0.027461f
C388 VTAIL.n182 B 0.027461f
C389 VTAIL.n183 B 0.014756f
C390 VTAIL.n184 B 0.015624f
C391 VTAIL.n185 B 0.034878f
C392 VTAIL.n186 B 0.034878f
C393 VTAIL.n187 B 0.015624f
C394 VTAIL.n188 B 0.014756f
C395 VTAIL.n189 B 0.027461f
C396 VTAIL.n190 B 0.027461f
C397 VTAIL.n191 B 0.014756f
C398 VTAIL.n192 B 0.015624f
C399 VTAIL.n193 B 0.034878f
C400 VTAIL.n194 B 0.075833f
C401 VTAIL.n195 B 0.015624f
C402 VTAIL.n196 B 0.014756f
C403 VTAIL.n197 B 0.065349f
C404 VTAIL.n198 B 0.042522f
C405 VTAIL.n199 B 1.39602f
C406 VTAIL.n200 B 0.038783f
C407 VTAIL.n201 B 0.027461f
C408 VTAIL.n202 B 0.014756f
C409 VTAIL.n203 B 0.034878f
C410 VTAIL.n204 B 0.015624f
C411 VTAIL.n205 B 0.027461f
C412 VTAIL.n206 B 0.014756f
C413 VTAIL.n207 B 0.034878f
C414 VTAIL.n208 B 0.01519f
C415 VTAIL.n209 B 0.027461f
C416 VTAIL.n210 B 0.015624f
C417 VTAIL.n211 B 0.034878f
C418 VTAIL.n212 B 0.015624f
C419 VTAIL.n213 B 0.027461f
C420 VTAIL.n214 B 0.014756f
C421 VTAIL.n215 B 0.034878f
C422 VTAIL.n216 B 0.015624f
C423 VTAIL.n217 B 1.31815f
C424 VTAIL.n218 B 0.014756f
C425 VTAIL.t7 B 0.058826f
C426 VTAIL.n219 B 0.192189f
C427 VTAIL.n220 B 0.024656f
C428 VTAIL.n221 B 0.026159f
C429 VTAIL.n222 B 0.034878f
C430 VTAIL.n223 B 0.015624f
C431 VTAIL.n224 B 0.014756f
C432 VTAIL.n225 B 0.027461f
C433 VTAIL.n226 B 0.027461f
C434 VTAIL.n227 B 0.014756f
C435 VTAIL.n228 B 0.015624f
C436 VTAIL.n229 B 0.034878f
C437 VTAIL.n230 B 0.034878f
C438 VTAIL.n231 B 0.015624f
C439 VTAIL.n232 B 0.014756f
C440 VTAIL.n233 B 0.027461f
C441 VTAIL.n234 B 0.027461f
C442 VTAIL.n235 B 0.014756f
C443 VTAIL.n236 B 0.014756f
C444 VTAIL.n237 B 0.015624f
C445 VTAIL.n238 B 0.034878f
C446 VTAIL.n239 B 0.034878f
C447 VTAIL.n240 B 0.034878f
C448 VTAIL.n241 B 0.01519f
C449 VTAIL.n242 B 0.014756f
C450 VTAIL.n243 B 0.027461f
C451 VTAIL.n244 B 0.027461f
C452 VTAIL.n245 B 0.014756f
C453 VTAIL.n246 B 0.015624f
C454 VTAIL.n247 B 0.034878f
C455 VTAIL.n248 B 0.034878f
C456 VTAIL.n249 B 0.015624f
C457 VTAIL.n250 B 0.014756f
C458 VTAIL.n251 B 0.027461f
C459 VTAIL.n252 B 0.027461f
C460 VTAIL.n253 B 0.014756f
C461 VTAIL.n254 B 0.015624f
C462 VTAIL.n255 B 0.034878f
C463 VTAIL.n256 B 0.075833f
C464 VTAIL.n257 B 0.015624f
C465 VTAIL.n258 B 0.014756f
C466 VTAIL.n259 B 0.065349f
C467 VTAIL.n260 B 0.042522f
C468 VTAIL.n261 B 1.39602f
C469 VTAIL.t3 B 0.248466f
C470 VTAIL.t2 B 0.248466f
C471 VTAIL.n262 B 2.12929f
C472 VTAIL.n263 B 0.340486f
C473 VDD1.n0 B 0.037122f
C474 VDD1.n1 B 0.026284f
C475 VDD1.n2 B 0.014124f
C476 VDD1.n3 B 0.033384f
C477 VDD1.n4 B 0.014955f
C478 VDD1.n5 B 0.026284f
C479 VDD1.n6 B 0.014124f
C480 VDD1.n7 B 0.033384f
C481 VDD1.n8 B 0.01454f
C482 VDD1.n9 B 0.026284f
C483 VDD1.n10 B 0.01454f
C484 VDD1.n11 B 0.014124f
C485 VDD1.n12 B 0.033384f
C486 VDD1.n13 B 0.033384f
C487 VDD1.n14 B 0.014955f
C488 VDD1.n15 B 0.026284f
C489 VDD1.n16 B 0.014124f
C490 VDD1.n17 B 0.033384f
C491 VDD1.n18 B 0.014955f
C492 VDD1.n19 B 1.2617f
C493 VDD1.n20 B 0.014124f
C494 VDD1.t9 B 0.056306f
C495 VDD1.n21 B 0.183958f
C496 VDD1.n22 B 0.0236f
C497 VDD1.n23 B 0.025038f
C498 VDD1.n24 B 0.033384f
C499 VDD1.n25 B 0.014955f
C500 VDD1.n26 B 0.014124f
C501 VDD1.n27 B 0.026284f
C502 VDD1.n28 B 0.026284f
C503 VDD1.n29 B 0.014124f
C504 VDD1.n30 B 0.014955f
C505 VDD1.n31 B 0.033384f
C506 VDD1.n32 B 0.033384f
C507 VDD1.n33 B 0.014955f
C508 VDD1.n34 B 0.014124f
C509 VDD1.n35 B 0.026284f
C510 VDD1.n36 B 0.026284f
C511 VDD1.n37 B 0.014124f
C512 VDD1.n38 B 0.014955f
C513 VDD1.n39 B 0.033384f
C514 VDD1.n40 B 0.033384f
C515 VDD1.n41 B 0.014955f
C516 VDD1.n42 B 0.014124f
C517 VDD1.n43 B 0.026284f
C518 VDD1.n44 B 0.026284f
C519 VDD1.n45 B 0.014124f
C520 VDD1.n46 B 0.014955f
C521 VDD1.n47 B 0.033384f
C522 VDD1.n48 B 0.033384f
C523 VDD1.n49 B 0.014955f
C524 VDD1.n50 B 0.014124f
C525 VDD1.n51 B 0.026284f
C526 VDD1.n52 B 0.026284f
C527 VDD1.n53 B 0.014124f
C528 VDD1.n54 B 0.014955f
C529 VDD1.n55 B 0.033384f
C530 VDD1.n56 B 0.072585f
C531 VDD1.n57 B 0.014955f
C532 VDD1.n58 B 0.014124f
C533 VDD1.n59 B 0.06255f
C534 VDD1.n60 B 0.060395f
C535 VDD1.t2 B 0.237824f
C536 VDD1.t3 B 0.237824f
C537 VDD1.n61 B 2.11394f
C538 VDD1.n62 B 0.405593f
C539 VDD1.n63 B 0.037122f
C540 VDD1.n64 B 0.026284f
C541 VDD1.n65 B 0.014124f
C542 VDD1.n66 B 0.033384f
C543 VDD1.n67 B 0.014955f
C544 VDD1.n68 B 0.026284f
C545 VDD1.n69 B 0.014124f
C546 VDD1.n70 B 0.033384f
C547 VDD1.n71 B 0.01454f
C548 VDD1.n72 B 0.026284f
C549 VDD1.n73 B 0.014955f
C550 VDD1.n74 B 0.033384f
C551 VDD1.n75 B 0.014955f
C552 VDD1.n76 B 0.026284f
C553 VDD1.n77 B 0.014124f
C554 VDD1.n78 B 0.033384f
C555 VDD1.n79 B 0.014955f
C556 VDD1.n80 B 1.2617f
C557 VDD1.n81 B 0.014124f
C558 VDD1.t6 B 0.056306f
C559 VDD1.n82 B 0.183958f
C560 VDD1.n83 B 0.0236f
C561 VDD1.n84 B 0.025038f
C562 VDD1.n85 B 0.033384f
C563 VDD1.n86 B 0.014955f
C564 VDD1.n87 B 0.014124f
C565 VDD1.n88 B 0.026284f
C566 VDD1.n89 B 0.026284f
C567 VDD1.n90 B 0.014124f
C568 VDD1.n91 B 0.014955f
C569 VDD1.n92 B 0.033384f
C570 VDD1.n93 B 0.033384f
C571 VDD1.n94 B 0.014955f
C572 VDD1.n95 B 0.014124f
C573 VDD1.n96 B 0.026284f
C574 VDD1.n97 B 0.026284f
C575 VDD1.n98 B 0.014124f
C576 VDD1.n99 B 0.014124f
C577 VDD1.n100 B 0.014955f
C578 VDD1.n101 B 0.033384f
C579 VDD1.n102 B 0.033384f
C580 VDD1.n103 B 0.033384f
C581 VDD1.n104 B 0.01454f
C582 VDD1.n105 B 0.014124f
C583 VDD1.n106 B 0.026284f
C584 VDD1.n107 B 0.026284f
C585 VDD1.n108 B 0.014124f
C586 VDD1.n109 B 0.014955f
C587 VDD1.n110 B 0.033384f
C588 VDD1.n111 B 0.033384f
C589 VDD1.n112 B 0.014955f
C590 VDD1.n113 B 0.014124f
C591 VDD1.n114 B 0.026284f
C592 VDD1.n115 B 0.026284f
C593 VDD1.n116 B 0.014124f
C594 VDD1.n117 B 0.014955f
C595 VDD1.n118 B 0.033384f
C596 VDD1.n119 B 0.072585f
C597 VDD1.n120 B 0.014955f
C598 VDD1.n121 B 0.014124f
C599 VDD1.n122 B 0.06255f
C600 VDD1.n123 B 0.060395f
C601 VDD1.t5 B 0.237824f
C602 VDD1.t7 B 0.237824f
C603 VDD1.n124 B 2.11393f
C604 VDD1.n125 B 0.401006f
C605 VDD1.t1 B 0.237824f
C606 VDD1.t8 B 0.237824f
C607 VDD1.n126 B 2.11638f
C608 VDD1.n127 B 1.92249f
C609 VDD1.t0 B 0.237824f
C610 VDD1.t4 B 0.237824f
C611 VDD1.n128 B 2.11393f
C612 VDD1.n129 B 2.37239f
C613 VP.n0 B 0.048759f
C614 VP.t1 B 0.780941f
C615 VP.n1 B 0.323362f
C616 VP.n2 B 0.048759f
C617 VP.n3 B 0.048759f
C618 VP.t4 B 0.780941f
C619 VP.t8 B 0.780941f
C620 VP.t5 B 0.780941f
C621 VP.n4 B 0.323362f
C622 VP.t6 B 0.790978f
C623 VP.n5 B 0.308264f
C624 VP.t9 B 0.780941f
C625 VP.n6 B 0.320205f
C626 VP.n7 B 0.011065f
C627 VP.n8 B 0.154044f
C628 VP.n9 B 0.048759f
C629 VP.n10 B 0.048759f
C630 VP.n11 B 0.011065f
C631 VP.n12 B 0.320205f
C632 VP.n13 B 0.31795f
C633 VP.n14 B 1.95157f
C634 VP.n15 B 1.99407f
C635 VP.t7 B 0.780941f
C636 VP.n16 B 0.31795f
C637 VP.t3 B 0.780941f
C638 VP.n17 B 0.320205f
C639 VP.n18 B 0.011065f
C640 VP.n19 B 0.048759f
C641 VP.n20 B 0.048759f
C642 VP.n21 B 0.048759f
C643 VP.n22 B 0.011065f
C644 VP.t0 B 0.780941f
C645 VP.n23 B 0.320205f
C646 VP.t2 B 0.780941f
C647 VP.n24 B 0.31795f
C648 VP.n25 B 0.037787f
.ends

