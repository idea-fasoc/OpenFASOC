* NGSPICE file created from diff_pair_sample_1153.ext - technology: sky130A

.subckt diff_pair_sample_1153 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t9 VN.t0 VDD2.t3 w_n4330_n1874# sky130_fd_pr__pfet_01v8 ad=0.74745 pd=4.86 as=0.74745 ps=4.86 w=4.53 l=3.87
X1 VDD1.t5 VP.t0 VTAIL.t10 w_n4330_n1874# sky130_fd_pr__pfet_01v8 ad=1.7667 pd=9.84 as=0.74745 ps=4.86 w=4.53 l=3.87
X2 B.t11 B.t9 B.t10 w_n4330_n1874# sky130_fd_pr__pfet_01v8 ad=1.7667 pd=9.84 as=0 ps=0 w=4.53 l=3.87
X3 VDD1.t4 VP.t1 VTAIL.t0 w_n4330_n1874# sky130_fd_pr__pfet_01v8 ad=0.74745 pd=4.86 as=1.7667 ps=9.84 w=4.53 l=3.87
X4 B.t8 B.t6 B.t7 w_n4330_n1874# sky130_fd_pr__pfet_01v8 ad=1.7667 pd=9.84 as=0 ps=0 w=4.53 l=3.87
X5 VDD1.t3 VP.t2 VTAIL.t11 w_n4330_n1874# sky130_fd_pr__pfet_01v8 ad=0.74745 pd=4.86 as=1.7667 ps=9.84 w=4.53 l=3.87
X6 B.t5 B.t3 B.t4 w_n4330_n1874# sky130_fd_pr__pfet_01v8 ad=1.7667 pd=9.84 as=0 ps=0 w=4.53 l=3.87
X7 VDD1.t2 VP.t3 VTAIL.t1 w_n4330_n1874# sky130_fd_pr__pfet_01v8 ad=1.7667 pd=9.84 as=0.74745 ps=4.86 w=4.53 l=3.87
X8 VDD2.t2 VN.t1 VTAIL.t8 w_n4330_n1874# sky130_fd_pr__pfet_01v8 ad=0.74745 pd=4.86 as=1.7667 ps=9.84 w=4.53 l=3.87
X9 VDD2.t5 VN.t2 VTAIL.t7 w_n4330_n1874# sky130_fd_pr__pfet_01v8 ad=1.7667 pd=9.84 as=0.74745 ps=4.86 w=4.53 l=3.87
X10 VTAIL.t2 VP.t4 VDD1.t1 w_n4330_n1874# sky130_fd_pr__pfet_01v8 ad=0.74745 pd=4.86 as=0.74745 ps=4.86 w=4.53 l=3.87
X11 VTAIL.t6 VN.t3 VDD2.t0 w_n4330_n1874# sky130_fd_pr__pfet_01v8 ad=0.74745 pd=4.86 as=0.74745 ps=4.86 w=4.53 l=3.87
X12 B.t2 B.t0 B.t1 w_n4330_n1874# sky130_fd_pr__pfet_01v8 ad=1.7667 pd=9.84 as=0 ps=0 w=4.53 l=3.87
X13 VDD2.t1 VN.t4 VTAIL.t5 w_n4330_n1874# sky130_fd_pr__pfet_01v8 ad=0.74745 pd=4.86 as=1.7667 ps=9.84 w=4.53 l=3.87
X14 VTAIL.t3 VP.t5 VDD1.t0 w_n4330_n1874# sky130_fd_pr__pfet_01v8 ad=0.74745 pd=4.86 as=0.74745 ps=4.86 w=4.53 l=3.87
X15 VDD2.t4 VN.t5 VTAIL.t4 w_n4330_n1874# sky130_fd_pr__pfet_01v8 ad=1.7667 pd=9.84 as=0.74745 ps=4.86 w=4.53 l=3.87
R0 VN.n37 VN.n20 161.3
R1 VN.n36 VN.n35 161.3
R2 VN.n34 VN.n21 161.3
R3 VN.n33 VN.n32 161.3
R4 VN.n31 VN.n22 161.3
R5 VN.n30 VN.n29 161.3
R6 VN.n28 VN.n23 161.3
R7 VN.n27 VN.n26 161.3
R8 VN.n17 VN.n0 161.3
R9 VN.n16 VN.n15 161.3
R10 VN.n14 VN.n1 161.3
R11 VN.n13 VN.n12 161.3
R12 VN.n11 VN.n2 161.3
R13 VN.n10 VN.n9 161.3
R14 VN.n8 VN.n3 161.3
R15 VN.n7 VN.n6 161.3
R16 VN.n5 VN.n4 62.8742
R17 VN.n25 VN.n24 62.8742
R18 VN.n4 VN.t2 60.3918
R19 VN.n24 VN.t1 60.3918
R20 VN.n19 VN.n18 60.1615
R21 VN.n39 VN.n38 60.1615
R22 VN.n12 VN.n11 55.0624
R23 VN.n32 VN.n31 55.0624
R24 VN VN.n39 48.2769
R25 VN.n5 VN.t3 28.2106
R26 VN.n18 VN.t4 28.2106
R27 VN.n25 VN.t0 28.2106
R28 VN.n38 VN.t5 28.2106
R29 VN.n12 VN.n1 25.9244
R30 VN.n32 VN.n21 25.9244
R31 VN.n6 VN.n3 24.4675
R32 VN.n10 VN.n3 24.4675
R33 VN.n11 VN.n10 24.4675
R34 VN.n16 VN.n1 24.4675
R35 VN.n17 VN.n16 24.4675
R36 VN.n31 VN.n30 24.4675
R37 VN.n30 VN.n23 24.4675
R38 VN.n26 VN.n23 24.4675
R39 VN.n37 VN.n36 24.4675
R40 VN.n36 VN.n21 24.4675
R41 VN.n18 VN.n17 22.0208
R42 VN.n38 VN.n37 22.0208
R43 VN.n6 VN.n5 12.234
R44 VN.n26 VN.n25 12.234
R45 VN.n27 VN.n24 2.62187
R46 VN.n7 VN.n4 2.62187
R47 VN.n39 VN.n20 0.417535
R48 VN.n19 VN.n0 0.417535
R49 VN VN.n19 0.394291
R50 VN.n35 VN.n20 0.189894
R51 VN.n35 VN.n34 0.189894
R52 VN.n34 VN.n33 0.189894
R53 VN.n33 VN.n22 0.189894
R54 VN.n29 VN.n22 0.189894
R55 VN.n29 VN.n28 0.189894
R56 VN.n28 VN.n27 0.189894
R57 VN.n8 VN.n7 0.189894
R58 VN.n9 VN.n8 0.189894
R59 VN.n9 VN.n2 0.189894
R60 VN.n13 VN.n2 0.189894
R61 VN.n14 VN.n13 0.189894
R62 VN.n15 VN.n14 0.189894
R63 VN.n15 VN.n0 0.189894
R64 VDD2.n43 VDD2.n25 756.745
R65 VDD2.n18 VDD2.n0 756.745
R66 VDD2.n44 VDD2.n43 585
R67 VDD2.n42 VDD2.n41 585
R68 VDD2.n29 VDD2.n28 585
R69 VDD2.n36 VDD2.n35 585
R70 VDD2.n34 VDD2.n33 585
R71 VDD2.n9 VDD2.n8 585
R72 VDD2.n11 VDD2.n10 585
R73 VDD2.n4 VDD2.n3 585
R74 VDD2.n17 VDD2.n16 585
R75 VDD2.n19 VDD2.n18 585
R76 VDD2.n32 VDD2.t4 328.587
R77 VDD2.n7 VDD2.t5 328.587
R78 VDD2.n43 VDD2.n42 171.744
R79 VDD2.n42 VDD2.n28 171.744
R80 VDD2.n35 VDD2.n28 171.744
R81 VDD2.n35 VDD2.n34 171.744
R82 VDD2.n10 VDD2.n9 171.744
R83 VDD2.n10 VDD2.n3 171.744
R84 VDD2.n17 VDD2.n3 171.744
R85 VDD2.n18 VDD2.n17 171.744
R86 VDD2.n24 VDD2.n23 104.347
R87 VDD2 VDD2.n49 104.344
R88 VDD2.n34 VDD2.t4 85.8723
R89 VDD2.n9 VDD2.t5 85.8723
R90 VDD2.n24 VDD2.n22 50.9425
R91 VDD2.n48 VDD2.n47 48.2823
R92 VDD2.n48 VDD2.n24 39.3877
R93 VDD2.n33 VDD2.n32 16.3651
R94 VDD2.n8 VDD2.n7 16.3651
R95 VDD2.n36 VDD2.n31 12.8005
R96 VDD2.n11 VDD2.n6 12.8005
R97 VDD2.n37 VDD2.n29 12.0247
R98 VDD2.n12 VDD2.n4 12.0247
R99 VDD2.n41 VDD2.n40 11.249
R100 VDD2.n16 VDD2.n15 11.249
R101 VDD2.n44 VDD2.n27 10.4732
R102 VDD2.n19 VDD2.n2 10.4732
R103 VDD2.n45 VDD2.n25 9.69747
R104 VDD2.n20 VDD2.n0 9.69747
R105 VDD2.n47 VDD2.n46 9.45567
R106 VDD2.n22 VDD2.n21 9.45567
R107 VDD2.n46 VDD2.n45 9.3005
R108 VDD2.n27 VDD2.n26 9.3005
R109 VDD2.n40 VDD2.n39 9.3005
R110 VDD2.n38 VDD2.n37 9.3005
R111 VDD2.n31 VDD2.n30 9.3005
R112 VDD2.n21 VDD2.n20 9.3005
R113 VDD2.n2 VDD2.n1 9.3005
R114 VDD2.n15 VDD2.n14 9.3005
R115 VDD2.n13 VDD2.n12 9.3005
R116 VDD2.n6 VDD2.n5 9.3005
R117 VDD2.n49 VDD2.t3 7.176
R118 VDD2.n49 VDD2.t2 7.176
R119 VDD2.n23 VDD2.t0 7.176
R120 VDD2.n23 VDD2.t1 7.176
R121 VDD2.n47 VDD2.n25 4.26717
R122 VDD2.n22 VDD2.n0 4.26717
R123 VDD2.n32 VDD2.n30 3.73474
R124 VDD2.n7 VDD2.n5 3.73474
R125 VDD2.n45 VDD2.n44 3.49141
R126 VDD2.n20 VDD2.n19 3.49141
R127 VDD2 VDD2.n48 2.77421
R128 VDD2.n41 VDD2.n27 2.71565
R129 VDD2.n16 VDD2.n2 2.71565
R130 VDD2.n40 VDD2.n29 1.93989
R131 VDD2.n15 VDD2.n4 1.93989
R132 VDD2.n37 VDD2.n36 1.16414
R133 VDD2.n12 VDD2.n11 1.16414
R134 VDD2.n33 VDD2.n31 0.388379
R135 VDD2.n8 VDD2.n6 0.388379
R136 VDD2.n46 VDD2.n26 0.155672
R137 VDD2.n39 VDD2.n26 0.155672
R138 VDD2.n39 VDD2.n38 0.155672
R139 VDD2.n38 VDD2.n30 0.155672
R140 VDD2.n13 VDD2.n5 0.155672
R141 VDD2.n14 VDD2.n13 0.155672
R142 VDD2.n14 VDD2.n1 0.155672
R143 VDD2.n21 VDD2.n1 0.155672
R144 VTAIL.n98 VTAIL.n80 756.745
R145 VTAIL.n20 VTAIL.n2 756.745
R146 VTAIL.n74 VTAIL.n56 756.745
R147 VTAIL.n48 VTAIL.n30 756.745
R148 VTAIL.n89 VTAIL.n88 585
R149 VTAIL.n91 VTAIL.n90 585
R150 VTAIL.n84 VTAIL.n83 585
R151 VTAIL.n97 VTAIL.n96 585
R152 VTAIL.n99 VTAIL.n98 585
R153 VTAIL.n11 VTAIL.n10 585
R154 VTAIL.n13 VTAIL.n12 585
R155 VTAIL.n6 VTAIL.n5 585
R156 VTAIL.n19 VTAIL.n18 585
R157 VTAIL.n21 VTAIL.n20 585
R158 VTAIL.n75 VTAIL.n74 585
R159 VTAIL.n73 VTAIL.n72 585
R160 VTAIL.n60 VTAIL.n59 585
R161 VTAIL.n67 VTAIL.n66 585
R162 VTAIL.n65 VTAIL.n64 585
R163 VTAIL.n49 VTAIL.n48 585
R164 VTAIL.n47 VTAIL.n46 585
R165 VTAIL.n34 VTAIL.n33 585
R166 VTAIL.n41 VTAIL.n40 585
R167 VTAIL.n39 VTAIL.n38 585
R168 VTAIL.n87 VTAIL.t5 328.587
R169 VTAIL.n9 VTAIL.t11 328.587
R170 VTAIL.n63 VTAIL.t0 328.587
R171 VTAIL.n37 VTAIL.t8 328.587
R172 VTAIL.n90 VTAIL.n89 171.744
R173 VTAIL.n90 VTAIL.n83 171.744
R174 VTAIL.n97 VTAIL.n83 171.744
R175 VTAIL.n98 VTAIL.n97 171.744
R176 VTAIL.n12 VTAIL.n11 171.744
R177 VTAIL.n12 VTAIL.n5 171.744
R178 VTAIL.n19 VTAIL.n5 171.744
R179 VTAIL.n20 VTAIL.n19 171.744
R180 VTAIL.n74 VTAIL.n73 171.744
R181 VTAIL.n73 VTAIL.n59 171.744
R182 VTAIL.n66 VTAIL.n59 171.744
R183 VTAIL.n66 VTAIL.n65 171.744
R184 VTAIL.n48 VTAIL.n47 171.744
R185 VTAIL.n47 VTAIL.n33 171.744
R186 VTAIL.n40 VTAIL.n33 171.744
R187 VTAIL.n40 VTAIL.n39 171.744
R188 VTAIL.n55 VTAIL.n54 86.8192
R189 VTAIL.n29 VTAIL.n28 86.8192
R190 VTAIL.n1 VTAIL.n0 86.8191
R191 VTAIL.n27 VTAIL.n26 86.8191
R192 VTAIL.n89 VTAIL.t5 85.8723
R193 VTAIL.n11 VTAIL.t11 85.8723
R194 VTAIL.n65 VTAIL.t0 85.8723
R195 VTAIL.n39 VTAIL.t8 85.8723
R196 VTAIL.n103 VTAIL.n102 31.6035
R197 VTAIL.n25 VTAIL.n24 31.6035
R198 VTAIL.n79 VTAIL.n78 31.6035
R199 VTAIL.n53 VTAIL.n52 31.6035
R200 VTAIL.n29 VTAIL.n27 23.5134
R201 VTAIL.n103 VTAIL.n79 19.8927
R202 VTAIL.n88 VTAIL.n87 16.3651
R203 VTAIL.n10 VTAIL.n9 16.3651
R204 VTAIL.n64 VTAIL.n63 16.3651
R205 VTAIL.n38 VTAIL.n37 16.3651
R206 VTAIL.n91 VTAIL.n86 12.8005
R207 VTAIL.n13 VTAIL.n8 12.8005
R208 VTAIL.n67 VTAIL.n62 12.8005
R209 VTAIL.n41 VTAIL.n36 12.8005
R210 VTAIL.n92 VTAIL.n84 12.0247
R211 VTAIL.n14 VTAIL.n6 12.0247
R212 VTAIL.n68 VTAIL.n60 12.0247
R213 VTAIL.n42 VTAIL.n34 12.0247
R214 VTAIL.n96 VTAIL.n95 11.249
R215 VTAIL.n18 VTAIL.n17 11.249
R216 VTAIL.n72 VTAIL.n71 11.249
R217 VTAIL.n46 VTAIL.n45 11.249
R218 VTAIL.n99 VTAIL.n82 10.4732
R219 VTAIL.n21 VTAIL.n4 10.4732
R220 VTAIL.n75 VTAIL.n58 10.4732
R221 VTAIL.n49 VTAIL.n32 10.4732
R222 VTAIL.n100 VTAIL.n80 9.69747
R223 VTAIL.n22 VTAIL.n2 9.69747
R224 VTAIL.n76 VTAIL.n56 9.69747
R225 VTAIL.n50 VTAIL.n30 9.69747
R226 VTAIL.n102 VTAIL.n101 9.45567
R227 VTAIL.n24 VTAIL.n23 9.45567
R228 VTAIL.n78 VTAIL.n77 9.45567
R229 VTAIL.n52 VTAIL.n51 9.45567
R230 VTAIL.n101 VTAIL.n100 9.3005
R231 VTAIL.n82 VTAIL.n81 9.3005
R232 VTAIL.n95 VTAIL.n94 9.3005
R233 VTAIL.n93 VTAIL.n92 9.3005
R234 VTAIL.n86 VTAIL.n85 9.3005
R235 VTAIL.n23 VTAIL.n22 9.3005
R236 VTAIL.n4 VTAIL.n3 9.3005
R237 VTAIL.n17 VTAIL.n16 9.3005
R238 VTAIL.n15 VTAIL.n14 9.3005
R239 VTAIL.n8 VTAIL.n7 9.3005
R240 VTAIL.n77 VTAIL.n76 9.3005
R241 VTAIL.n58 VTAIL.n57 9.3005
R242 VTAIL.n71 VTAIL.n70 9.3005
R243 VTAIL.n69 VTAIL.n68 9.3005
R244 VTAIL.n62 VTAIL.n61 9.3005
R245 VTAIL.n51 VTAIL.n50 9.3005
R246 VTAIL.n32 VTAIL.n31 9.3005
R247 VTAIL.n45 VTAIL.n44 9.3005
R248 VTAIL.n43 VTAIL.n42 9.3005
R249 VTAIL.n36 VTAIL.n35 9.3005
R250 VTAIL.n0 VTAIL.t7 7.176
R251 VTAIL.n0 VTAIL.t6 7.176
R252 VTAIL.n26 VTAIL.t10 7.176
R253 VTAIL.n26 VTAIL.t2 7.176
R254 VTAIL.n54 VTAIL.t1 7.176
R255 VTAIL.n54 VTAIL.t3 7.176
R256 VTAIL.n28 VTAIL.t4 7.176
R257 VTAIL.n28 VTAIL.t9 7.176
R258 VTAIL.n102 VTAIL.n80 4.26717
R259 VTAIL.n24 VTAIL.n2 4.26717
R260 VTAIL.n78 VTAIL.n56 4.26717
R261 VTAIL.n52 VTAIL.n30 4.26717
R262 VTAIL.n87 VTAIL.n85 3.73474
R263 VTAIL.n9 VTAIL.n7 3.73474
R264 VTAIL.n63 VTAIL.n61 3.73474
R265 VTAIL.n37 VTAIL.n35 3.73474
R266 VTAIL.n53 VTAIL.n29 3.62119
R267 VTAIL.n79 VTAIL.n55 3.62119
R268 VTAIL.n27 VTAIL.n25 3.62119
R269 VTAIL.n100 VTAIL.n99 3.49141
R270 VTAIL.n22 VTAIL.n21 3.49141
R271 VTAIL.n76 VTAIL.n75 3.49141
R272 VTAIL.n50 VTAIL.n49 3.49141
R273 VTAIL.n96 VTAIL.n82 2.71565
R274 VTAIL.n18 VTAIL.n4 2.71565
R275 VTAIL.n72 VTAIL.n58 2.71565
R276 VTAIL.n46 VTAIL.n32 2.71565
R277 VTAIL VTAIL.n103 2.65783
R278 VTAIL.n55 VTAIL.n53 2.28067
R279 VTAIL.n25 VTAIL.n1 2.28067
R280 VTAIL.n95 VTAIL.n84 1.93989
R281 VTAIL.n17 VTAIL.n6 1.93989
R282 VTAIL.n71 VTAIL.n60 1.93989
R283 VTAIL.n45 VTAIL.n34 1.93989
R284 VTAIL.n92 VTAIL.n91 1.16414
R285 VTAIL.n14 VTAIL.n13 1.16414
R286 VTAIL.n68 VTAIL.n67 1.16414
R287 VTAIL.n42 VTAIL.n41 1.16414
R288 VTAIL VTAIL.n1 0.963862
R289 VTAIL.n88 VTAIL.n86 0.388379
R290 VTAIL.n10 VTAIL.n8 0.388379
R291 VTAIL.n64 VTAIL.n62 0.388379
R292 VTAIL.n38 VTAIL.n36 0.388379
R293 VTAIL.n93 VTAIL.n85 0.155672
R294 VTAIL.n94 VTAIL.n93 0.155672
R295 VTAIL.n94 VTAIL.n81 0.155672
R296 VTAIL.n101 VTAIL.n81 0.155672
R297 VTAIL.n15 VTAIL.n7 0.155672
R298 VTAIL.n16 VTAIL.n15 0.155672
R299 VTAIL.n16 VTAIL.n3 0.155672
R300 VTAIL.n23 VTAIL.n3 0.155672
R301 VTAIL.n77 VTAIL.n57 0.155672
R302 VTAIL.n70 VTAIL.n57 0.155672
R303 VTAIL.n70 VTAIL.n69 0.155672
R304 VTAIL.n69 VTAIL.n61 0.155672
R305 VTAIL.n51 VTAIL.n31 0.155672
R306 VTAIL.n44 VTAIL.n31 0.155672
R307 VTAIL.n44 VTAIL.n43 0.155672
R308 VTAIL.n43 VTAIL.n35 0.155672
R309 VP.n15 VP.n14 161.3
R310 VP.n16 VP.n11 161.3
R311 VP.n18 VP.n17 161.3
R312 VP.n19 VP.n10 161.3
R313 VP.n21 VP.n20 161.3
R314 VP.n22 VP.n9 161.3
R315 VP.n24 VP.n23 161.3
R316 VP.n25 VP.n8 161.3
R317 VP.n54 VP.n0 161.3
R318 VP.n53 VP.n52 161.3
R319 VP.n51 VP.n1 161.3
R320 VP.n50 VP.n49 161.3
R321 VP.n48 VP.n2 161.3
R322 VP.n47 VP.n46 161.3
R323 VP.n45 VP.n3 161.3
R324 VP.n44 VP.n43 161.3
R325 VP.n41 VP.n4 161.3
R326 VP.n40 VP.n39 161.3
R327 VP.n38 VP.n5 161.3
R328 VP.n37 VP.n36 161.3
R329 VP.n35 VP.n6 161.3
R330 VP.n34 VP.n33 161.3
R331 VP.n32 VP.n7 161.3
R332 VP.n31 VP.n30 161.3
R333 VP.n13 VP.n12 62.8743
R334 VP.n12 VP.t3 60.3914
R335 VP.n29 VP.n28 60.1615
R336 VP.n56 VP.n55 60.1615
R337 VP.n27 VP.n26 60.1615
R338 VP.n36 VP.n35 55.0624
R339 VP.n49 VP.n48 55.0624
R340 VP.n20 VP.n19 55.0624
R341 VP.n28 VP.n27 48.2388
R342 VP.n29 VP.t0 28.2106
R343 VP.n42 VP.t4 28.2106
R344 VP.n55 VP.t2 28.2106
R345 VP.n26 VP.t1 28.2106
R346 VP.n13 VP.t5 28.2106
R347 VP.n35 VP.n34 25.9244
R348 VP.n49 VP.n1 25.9244
R349 VP.n20 VP.n9 25.9244
R350 VP.n30 VP.n7 24.4675
R351 VP.n34 VP.n7 24.4675
R352 VP.n36 VP.n5 24.4675
R353 VP.n40 VP.n5 24.4675
R354 VP.n41 VP.n40 24.4675
R355 VP.n43 VP.n3 24.4675
R356 VP.n47 VP.n3 24.4675
R357 VP.n48 VP.n47 24.4675
R358 VP.n53 VP.n1 24.4675
R359 VP.n54 VP.n53 24.4675
R360 VP.n24 VP.n9 24.4675
R361 VP.n25 VP.n24 24.4675
R362 VP.n14 VP.n11 24.4675
R363 VP.n18 VP.n11 24.4675
R364 VP.n19 VP.n18 24.4675
R365 VP.n30 VP.n29 22.0208
R366 VP.n55 VP.n54 22.0208
R367 VP.n26 VP.n25 22.0208
R368 VP.n42 VP.n41 12.234
R369 VP.n43 VP.n42 12.234
R370 VP.n14 VP.n13 12.234
R371 VP.n15 VP.n12 2.62184
R372 VP.n27 VP.n8 0.417535
R373 VP.n31 VP.n28 0.417535
R374 VP.n56 VP.n0 0.417535
R375 VP VP.n56 0.394291
R376 VP.n16 VP.n15 0.189894
R377 VP.n17 VP.n16 0.189894
R378 VP.n17 VP.n10 0.189894
R379 VP.n21 VP.n10 0.189894
R380 VP.n22 VP.n21 0.189894
R381 VP.n23 VP.n22 0.189894
R382 VP.n23 VP.n8 0.189894
R383 VP.n32 VP.n31 0.189894
R384 VP.n33 VP.n32 0.189894
R385 VP.n33 VP.n6 0.189894
R386 VP.n37 VP.n6 0.189894
R387 VP.n38 VP.n37 0.189894
R388 VP.n39 VP.n38 0.189894
R389 VP.n39 VP.n4 0.189894
R390 VP.n44 VP.n4 0.189894
R391 VP.n45 VP.n44 0.189894
R392 VP.n46 VP.n45 0.189894
R393 VP.n46 VP.n2 0.189894
R394 VP.n50 VP.n2 0.189894
R395 VP.n51 VP.n50 0.189894
R396 VP.n52 VP.n51 0.189894
R397 VP.n52 VP.n0 0.189894
R398 VDD1.n18 VDD1.n0 756.745
R399 VDD1.n41 VDD1.n23 756.745
R400 VDD1.n19 VDD1.n18 585
R401 VDD1.n17 VDD1.n16 585
R402 VDD1.n4 VDD1.n3 585
R403 VDD1.n11 VDD1.n10 585
R404 VDD1.n9 VDD1.n8 585
R405 VDD1.n32 VDD1.n31 585
R406 VDD1.n34 VDD1.n33 585
R407 VDD1.n27 VDD1.n26 585
R408 VDD1.n40 VDD1.n39 585
R409 VDD1.n42 VDD1.n41 585
R410 VDD1.n7 VDD1.t2 328.587
R411 VDD1.n30 VDD1.t5 328.587
R412 VDD1.n18 VDD1.n17 171.744
R413 VDD1.n17 VDD1.n3 171.744
R414 VDD1.n10 VDD1.n3 171.744
R415 VDD1.n10 VDD1.n9 171.744
R416 VDD1.n33 VDD1.n32 171.744
R417 VDD1.n33 VDD1.n26 171.744
R418 VDD1.n40 VDD1.n26 171.744
R419 VDD1.n41 VDD1.n40 171.744
R420 VDD1.n47 VDD1.n46 104.347
R421 VDD1.n49 VDD1.n48 103.498
R422 VDD1.n9 VDD1.t2 85.8723
R423 VDD1.n32 VDD1.t5 85.8723
R424 VDD1 VDD1.n22 51.056
R425 VDD1.n47 VDD1.n45 50.9425
R426 VDD1.n49 VDD1.n47 41.7811
R427 VDD1.n8 VDD1.n7 16.3651
R428 VDD1.n31 VDD1.n30 16.3651
R429 VDD1.n11 VDD1.n6 12.8005
R430 VDD1.n34 VDD1.n29 12.8005
R431 VDD1.n12 VDD1.n4 12.0247
R432 VDD1.n35 VDD1.n27 12.0247
R433 VDD1.n16 VDD1.n15 11.249
R434 VDD1.n39 VDD1.n38 11.249
R435 VDD1.n19 VDD1.n2 10.4732
R436 VDD1.n42 VDD1.n25 10.4732
R437 VDD1.n20 VDD1.n0 9.69747
R438 VDD1.n43 VDD1.n23 9.69747
R439 VDD1.n22 VDD1.n21 9.45567
R440 VDD1.n45 VDD1.n44 9.45567
R441 VDD1.n21 VDD1.n20 9.3005
R442 VDD1.n2 VDD1.n1 9.3005
R443 VDD1.n15 VDD1.n14 9.3005
R444 VDD1.n13 VDD1.n12 9.3005
R445 VDD1.n6 VDD1.n5 9.3005
R446 VDD1.n44 VDD1.n43 9.3005
R447 VDD1.n25 VDD1.n24 9.3005
R448 VDD1.n38 VDD1.n37 9.3005
R449 VDD1.n36 VDD1.n35 9.3005
R450 VDD1.n29 VDD1.n28 9.3005
R451 VDD1.n48 VDD1.t0 7.176
R452 VDD1.n48 VDD1.t4 7.176
R453 VDD1.n46 VDD1.t1 7.176
R454 VDD1.n46 VDD1.t3 7.176
R455 VDD1.n22 VDD1.n0 4.26717
R456 VDD1.n45 VDD1.n23 4.26717
R457 VDD1.n7 VDD1.n5 3.73474
R458 VDD1.n30 VDD1.n28 3.73474
R459 VDD1.n20 VDD1.n19 3.49141
R460 VDD1.n43 VDD1.n42 3.49141
R461 VDD1.n16 VDD1.n2 2.71565
R462 VDD1.n39 VDD1.n25 2.71565
R463 VDD1.n15 VDD1.n4 1.93989
R464 VDD1.n38 VDD1.n27 1.93989
R465 VDD1.n12 VDD1.n11 1.16414
R466 VDD1.n35 VDD1.n34 1.16414
R467 VDD1 VDD1.n49 0.847483
R468 VDD1.n8 VDD1.n6 0.388379
R469 VDD1.n31 VDD1.n29 0.388379
R470 VDD1.n21 VDD1.n1 0.155672
R471 VDD1.n14 VDD1.n1 0.155672
R472 VDD1.n14 VDD1.n13 0.155672
R473 VDD1.n13 VDD1.n5 0.155672
R474 VDD1.n36 VDD1.n28 0.155672
R475 VDD1.n37 VDD1.n36 0.155672
R476 VDD1.n37 VDD1.n24 0.155672
R477 VDD1.n44 VDD1.n24 0.155672
R478 B.n333 B.n118 585
R479 B.n332 B.n331 585
R480 B.n330 B.n119 585
R481 B.n329 B.n328 585
R482 B.n327 B.n120 585
R483 B.n326 B.n325 585
R484 B.n324 B.n121 585
R485 B.n323 B.n322 585
R486 B.n321 B.n122 585
R487 B.n320 B.n319 585
R488 B.n318 B.n123 585
R489 B.n317 B.n316 585
R490 B.n315 B.n124 585
R491 B.n314 B.n313 585
R492 B.n312 B.n125 585
R493 B.n311 B.n310 585
R494 B.n309 B.n126 585
R495 B.n308 B.n307 585
R496 B.n306 B.n127 585
R497 B.n305 B.n304 585
R498 B.n302 B.n128 585
R499 B.n301 B.n300 585
R500 B.n299 B.n131 585
R501 B.n298 B.n297 585
R502 B.n296 B.n132 585
R503 B.n295 B.n294 585
R504 B.n293 B.n133 585
R505 B.n292 B.n291 585
R506 B.n290 B.n134 585
R507 B.n288 B.n287 585
R508 B.n286 B.n137 585
R509 B.n285 B.n284 585
R510 B.n283 B.n138 585
R511 B.n282 B.n281 585
R512 B.n280 B.n139 585
R513 B.n279 B.n278 585
R514 B.n277 B.n140 585
R515 B.n276 B.n275 585
R516 B.n274 B.n141 585
R517 B.n273 B.n272 585
R518 B.n271 B.n142 585
R519 B.n270 B.n269 585
R520 B.n268 B.n143 585
R521 B.n267 B.n266 585
R522 B.n265 B.n144 585
R523 B.n264 B.n263 585
R524 B.n262 B.n145 585
R525 B.n261 B.n260 585
R526 B.n259 B.n146 585
R527 B.n335 B.n334 585
R528 B.n336 B.n117 585
R529 B.n338 B.n337 585
R530 B.n339 B.n116 585
R531 B.n341 B.n340 585
R532 B.n342 B.n115 585
R533 B.n344 B.n343 585
R534 B.n345 B.n114 585
R535 B.n347 B.n346 585
R536 B.n348 B.n113 585
R537 B.n350 B.n349 585
R538 B.n351 B.n112 585
R539 B.n353 B.n352 585
R540 B.n354 B.n111 585
R541 B.n356 B.n355 585
R542 B.n357 B.n110 585
R543 B.n359 B.n358 585
R544 B.n360 B.n109 585
R545 B.n362 B.n361 585
R546 B.n363 B.n108 585
R547 B.n365 B.n364 585
R548 B.n366 B.n107 585
R549 B.n368 B.n367 585
R550 B.n369 B.n106 585
R551 B.n371 B.n370 585
R552 B.n372 B.n105 585
R553 B.n374 B.n373 585
R554 B.n375 B.n104 585
R555 B.n377 B.n376 585
R556 B.n378 B.n103 585
R557 B.n380 B.n379 585
R558 B.n381 B.n102 585
R559 B.n383 B.n382 585
R560 B.n384 B.n101 585
R561 B.n386 B.n385 585
R562 B.n387 B.n100 585
R563 B.n389 B.n388 585
R564 B.n390 B.n99 585
R565 B.n392 B.n391 585
R566 B.n393 B.n98 585
R567 B.n395 B.n394 585
R568 B.n396 B.n97 585
R569 B.n398 B.n397 585
R570 B.n399 B.n96 585
R571 B.n401 B.n400 585
R572 B.n402 B.n95 585
R573 B.n404 B.n403 585
R574 B.n405 B.n94 585
R575 B.n407 B.n406 585
R576 B.n408 B.n93 585
R577 B.n410 B.n409 585
R578 B.n411 B.n92 585
R579 B.n413 B.n412 585
R580 B.n414 B.n91 585
R581 B.n416 B.n415 585
R582 B.n417 B.n90 585
R583 B.n419 B.n418 585
R584 B.n420 B.n89 585
R585 B.n422 B.n421 585
R586 B.n423 B.n88 585
R587 B.n425 B.n424 585
R588 B.n426 B.n87 585
R589 B.n428 B.n427 585
R590 B.n429 B.n86 585
R591 B.n431 B.n430 585
R592 B.n432 B.n85 585
R593 B.n434 B.n433 585
R594 B.n435 B.n84 585
R595 B.n437 B.n436 585
R596 B.n438 B.n83 585
R597 B.n440 B.n439 585
R598 B.n441 B.n82 585
R599 B.n443 B.n442 585
R600 B.n444 B.n81 585
R601 B.n446 B.n445 585
R602 B.n447 B.n80 585
R603 B.n449 B.n448 585
R604 B.n450 B.n79 585
R605 B.n452 B.n451 585
R606 B.n453 B.n78 585
R607 B.n455 B.n454 585
R608 B.n456 B.n77 585
R609 B.n458 B.n457 585
R610 B.n459 B.n76 585
R611 B.n461 B.n460 585
R612 B.n462 B.n75 585
R613 B.n464 B.n463 585
R614 B.n465 B.n74 585
R615 B.n467 B.n466 585
R616 B.n468 B.n73 585
R617 B.n470 B.n469 585
R618 B.n471 B.n72 585
R619 B.n473 B.n472 585
R620 B.n474 B.n71 585
R621 B.n476 B.n475 585
R622 B.n477 B.n70 585
R623 B.n479 B.n478 585
R624 B.n480 B.n69 585
R625 B.n482 B.n481 585
R626 B.n483 B.n68 585
R627 B.n485 B.n484 585
R628 B.n486 B.n67 585
R629 B.n488 B.n487 585
R630 B.n489 B.n66 585
R631 B.n491 B.n490 585
R632 B.n492 B.n65 585
R633 B.n494 B.n493 585
R634 B.n495 B.n64 585
R635 B.n497 B.n496 585
R636 B.n498 B.n63 585
R637 B.n500 B.n499 585
R638 B.n501 B.n62 585
R639 B.n503 B.n502 585
R640 B.n504 B.n61 585
R641 B.n506 B.n505 585
R642 B.n507 B.n60 585
R643 B.n582 B.n581 585
R644 B.n580 B.n31 585
R645 B.n579 B.n578 585
R646 B.n577 B.n32 585
R647 B.n576 B.n575 585
R648 B.n574 B.n33 585
R649 B.n573 B.n572 585
R650 B.n571 B.n34 585
R651 B.n570 B.n569 585
R652 B.n568 B.n35 585
R653 B.n567 B.n566 585
R654 B.n565 B.n36 585
R655 B.n564 B.n563 585
R656 B.n562 B.n37 585
R657 B.n561 B.n560 585
R658 B.n559 B.n38 585
R659 B.n558 B.n557 585
R660 B.n556 B.n39 585
R661 B.n555 B.n554 585
R662 B.n553 B.n40 585
R663 B.n552 B.n551 585
R664 B.n550 B.n41 585
R665 B.n549 B.n548 585
R666 B.n547 B.n45 585
R667 B.n546 B.n545 585
R668 B.n544 B.n46 585
R669 B.n543 B.n542 585
R670 B.n541 B.n47 585
R671 B.n540 B.n539 585
R672 B.n537 B.n48 585
R673 B.n536 B.n535 585
R674 B.n534 B.n51 585
R675 B.n533 B.n532 585
R676 B.n531 B.n52 585
R677 B.n530 B.n529 585
R678 B.n528 B.n53 585
R679 B.n527 B.n526 585
R680 B.n525 B.n54 585
R681 B.n524 B.n523 585
R682 B.n522 B.n55 585
R683 B.n521 B.n520 585
R684 B.n519 B.n56 585
R685 B.n518 B.n517 585
R686 B.n516 B.n57 585
R687 B.n515 B.n514 585
R688 B.n513 B.n58 585
R689 B.n512 B.n511 585
R690 B.n510 B.n59 585
R691 B.n509 B.n508 585
R692 B.n583 B.n30 585
R693 B.n585 B.n584 585
R694 B.n586 B.n29 585
R695 B.n588 B.n587 585
R696 B.n589 B.n28 585
R697 B.n591 B.n590 585
R698 B.n592 B.n27 585
R699 B.n594 B.n593 585
R700 B.n595 B.n26 585
R701 B.n597 B.n596 585
R702 B.n598 B.n25 585
R703 B.n600 B.n599 585
R704 B.n601 B.n24 585
R705 B.n603 B.n602 585
R706 B.n604 B.n23 585
R707 B.n606 B.n605 585
R708 B.n607 B.n22 585
R709 B.n609 B.n608 585
R710 B.n610 B.n21 585
R711 B.n612 B.n611 585
R712 B.n613 B.n20 585
R713 B.n615 B.n614 585
R714 B.n616 B.n19 585
R715 B.n618 B.n617 585
R716 B.n619 B.n18 585
R717 B.n621 B.n620 585
R718 B.n622 B.n17 585
R719 B.n624 B.n623 585
R720 B.n625 B.n16 585
R721 B.n627 B.n626 585
R722 B.n628 B.n15 585
R723 B.n630 B.n629 585
R724 B.n631 B.n14 585
R725 B.n633 B.n632 585
R726 B.n634 B.n13 585
R727 B.n636 B.n635 585
R728 B.n637 B.n12 585
R729 B.n639 B.n638 585
R730 B.n640 B.n11 585
R731 B.n642 B.n641 585
R732 B.n643 B.n10 585
R733 B.n645 B.n644 585
R734 B.n646 B.n9 585
R735 B.n648 B.n647 585
R736 B.n649 B.n8 585
R737 B.n651 B.n650 585
R738 B.n652 B.n7 585
R739 B.n654 B.n653 585
R740 B.n655 B.n6 585
R741 B.n657 B.n656 585
R742 B.n658 B.n5 585
R743 B.n660 B.n659 585
R744 B.n661 B.n4 585
R745 B.n663 B.n662 585
R746 B.n664 B.n3 585
R747 B.n666 B.n665 585
R748 B.n667 B.n0 585
R749 B.n2 B.n1 585
R750 B.n175 B.n174 585
R751 B.n177 B.n176 585
R752 B.n178 B.n173 585
R753 B.n180 B.n179 585
R754 B.n181 B.n172 585
R755 B.n183 B.n182 585
R756 B.n184 B.n171 585
R757 B.n186 B.n185 585
R758 B.n187 B.n170 585
R759 B.n189 B.n188 585
R760 B.n190 B.n169 585
R761 B.n192 B.n191 585
R762 B.n193 B.n168 585
R763 B.n195 B.n194 585
R764 B.n196 B.n167 585
R765 B.n198 B.n197 585
R766 B.n199 B.n166 585
R767 B.n201 B.n200 585
R768 B.n202 B.n165 585
R769 B.n204 B.n203 585
R770 B.n205 B.n164 585
R771 B.n207 B.n206 585
R772 B.n208 B.n163 585
R773 B.n210 B.n209 585
R774 B.n211 B.n162 585
R775 B.n213 B.n212 585
R776 B.n214 B.n161 585
R777 B.n216 B.n215 585
R778 B.n217 B.n160 585
R779 B.n219 B.n218 585
R780 B.n220 B.n159 585
R781 B.n222 B.n221 585
R782 B.n223 B.n158 585
R783 B.n225 B.n224 585
R784 B.n226 B.n157 585
R785 B.n228 B.n227 585
R786 B.n229 B.n156 585
R787 B.n231 B.n230 585
R788 B.n232 B.n155 585
R789 B.n234 B.n233 585
R790 B.n235 B.n154 585
R791 B.n237 B.n236 585
R792 B.n238 B.n153 585
R793 B.n240 B.n239 585
R794 B.n241 B.n152 585
R795 B.n243 B.n242 585
R796 B.n244 B.n151 585
R797 B.n246 B.n245 585
R798 B.n247 B.n150 585
R799 B.n249 B.n248 585
R800 B.n250 B.n149 585
R801 B.n252 B.n251 585
R802 B.n253 B.n148 585
R803 B.n255 B.n254 585
R804 B.n256 B.n147 585
R805 B.n258 B.n257 585
R806 B.n257 B.n146 492.5
R807 B.n335 B.n118 492.5
R808 B.n509 B.n60 492.5
R809 B.n583 B.n582 492.5
R810 B.n129 B.t7 324.442
R811 B.n49 B.t11 324.442
R812 B.n135 B.t4 324.442
R813 B.n42 B.t2 324.442
R814 B.n669 B.n668 256.663
R815 B.n130 B.t8 242.988
R816 B.n50 B.t10 242.988
R817 B.n136 B.t5 242.987
R818 B.n43 B.t1 242.987
R819 B.n135 B.t3 237.607
R820 B.n129 B.t6 237.607
R821 B.n49 B.t9 237.607
R822 B.n42 B.t0 237.607
R823 B.n668 B.n667 235.042
R824 B.n668 B.n2 235.042
R825 B.n261 B.n146 163.367
R826 B.n262 B.n261 163.367
R827 B.n263 B.n262 163.367
R828 B.n263 B.n144 163.367
R829 B.n267 B.n144 163.367
R830 B.n268 B.n267 163.367
R831 B.n269 B.n268 163.367
R832 B.n269 B.n142 163.367
R833 B.n273 B.n142 163.367
R834 B.n274 B.n273 163.367
R835 B.n275 B.n274 163.367
R836 B.n275 B.n140 163.367
R837 B.n279 B.n140 163.367
R838 B.n280 B.n279 163.367
R839 B.n281 B.n280 163.367
R840 B.n281 B.n138 163.367
R841 B.n285 B.n138 163.367
R842 B.n286 B.n285 163.367
R843 B.n287 B.n286 163.367
R844 B.n287 B.n134 163.367
R845 B.n292 B.n134 163.367
R846 B.n293 B.n292 163.367
R847 B.n294 B.n293 163.367
R848 B.n294 B.n132 163.367
R849 B.n298 B.n132 163.367
R850 B.n299 B.n298 163.367
R851 B.n300 B.n299 163.367
R852 B.n300 B.n128 163.367
R853 B.n305 B.n128 163.367
R854 B.n306 B.n305 163.367
R855 B.n307 B.n306 163.367
R856 B.n307 B.n126 163.367
R857 B.n311 B.n126 163.367
R858 B.n312 B.n311 163.367
R859 B.n313 B.n312 163.367
R860 B.n313 B.n124 163.367
R861 B.n317 B.n124 163.367
R862 B.n318 B.n317 163.367
R863 B.n319 B.n318 163.367
R864 B.n319 B.n122 163.367
R865 B.n323 B.n122 163.367
R866 B.n324 B.n323 163.367
R867 B.n325 B.n324 163.367
R868 B.n325 B.n120 163.367
R869 B.n329 B.n120 163.367
R870 B.n330 B.n329 163.367
R871 B.n331 B.n330 163.367
R872 B.n331 B.n118 163.367
R873 B.n505 B.n60 163.367
R874 B.n505 B.n504 163.367
R875 B.n504 B.n503 163.367
R876 B.n503 B.n62 163.367
R877 B.n499 B.n62 163.367
R878 B.n499 B.n498 163.367
R879 B.n498 B.n497 163.367
R880 B.n497 B.n64 163.367
R881 B.n493 B.n64 163.367
R882 B.n493 B.n492 163.367
R883 B.n492 B.n491 163.367
R884 B.n491 B.n66 163.367
R885 B.n487 B.n66 163.367
R886 B.n487 B.n486 163.367
R887 B.n486 B.n485 163.367
R888 B.n485 B.n68 163.367
R889 B.n481 B.n68 163.367
R890 B.n481 B.n480 163.367
R891 B.n480 B.n479 163.367
R892 B.n479 B.n70 163.367
R893 B.n475 B.n70 163.367
R894 B.n475 B.n474 163.367
R895 B.n474 B.n473 163.367
R896 B.n473 B.n72 163.367
R897 B.n469 B.n72 163.367
R898 B.n469 B.n468 163.367
R899 B.n468 B.n467 163.367
R900 B.n467 B.n74 163.367
R901 B.n463 B.n74 163.367
R902 B.n463 B.n462 163.367
R903 B.n462 B.n461 163.367
R904 B.n461 B.n76 163.367
R905 B.n457 B.n76 163.367
R906 B.n457 B.n456 163.367
R907 B.n456 B.n455 163.367
R908 B.n455 B.n78 163.367
R909 B.n451 B.n78 163.367
R910 B.n451 B.n450 163.367
R911 B.n450 B.n449 163.367
R912 B.n449 B.n80 163.367
R913 B.n445 B.n80 163.367
R914 B.n445 B.n444 163.367
R915 B.n444 B.n443 163.367
R916 B.n443 B.n82 163.367
R917 B.n439 B.n82 163.367
R918 B.n439 B.n438 163.367
R919 B.n438 B.n437 163.367
R920 B.n437 B.n84 163.367
R921 B.n433 B.n84 163.367
R922 B.n433 B.n432 163.367
R923 B.n432 B.n431 163.367
R924 B.n431 B.n86 163.367
R925 B.n427 B.n86 163.367
R926 B.n427 B.n426 163.367
R927 B.n426 B.n425 163.367
R928 B.n425 B.n88 163.367
R929 B.n421 B.n88 163.367
R930 B.n421 B.n420 163.367
R931 B.n420 B.n419 163.367
R932 B.n419 B.n90 163.367
R933 B.n415 B.n90 163.367
R934 B.n415 B.n414 163.367
R935 B.n414 B.n413 163.367
R936 B.n413 B.n92 163.367
R937 B.n409 B.n92 163.367
R938 B.n409 B.n408 163.367
R939 B.n408 B.n407 163.367
R940 B.n407 B.n94 163.367
R941 B.n403 B.n94 163.367
R942 B.n403 B.n402 163.367
R943 B.n402 B.n401 163.367
R944 B.n401 B.n96 163.367
R945 B.n397 B.n96 163.367
R946 B.n397 B.n396 163.367
R947 B.n396 B.n395 163.367
R948 B.n395 B.n98 163.367
R949 B.n391 B.n98 163.367
R950 B.n391 B.n390 163.367
R951 B.n390 B.n389 163.367
R952 B.n389 B.n100 163.367
R953 B.n385 B.n100 163.367
R954 B.n385 B.n384 163.367
R955 B.n384 B.n383 163.367
R956 B.n383 B.n102 163.367
R957 B.n379 B.n102 163.367
R958 B.n379 B.n378 163.367
R959 B.n378 B.n377 163.367
R960 B.n377 B.n104 163.367
R961 B.n373 B.n104 163.367
R962 B.n373 B.n372 163.367
R963 B.n372 B.n371 163.367
R964 B.n371 B.n106 163.367
R965 B.n367 B.n106 163.367
R966 B.n367 B.n366 163.367
R967 B.n366 B.n365 163.367
R968 B.n365 B.n108 163.367
R969 B.n361 B.n108 163.367
R970 B.n361 B.n360 163.367
R971 B.n360 B.n359 163.367
R972 B.n359 B.n110 163.367
R973 B.n355 B.n110 163.367
R974 B.n355 B.n354 163.367
R975 B.n354 B.n353 163.367
R976 B.n353 B.n112 163.367
R977 B.n349 B.n112 163.367
R978 B.n349 B.n348 163.367
R979 B.n348 B.n347 163.367
R980 B.n347 B.n114 163.367
R981 B.n343 B.n114 163.367
R982 B.n343 B.n342 163.367
R983 B.n342 B.n341 163.367
R984 B.n341 B.n116 163.367
R985 B.n337 B.n116 163.367
R986 B.n337 B.n336 163.367
R987 B.n336 B.n335 163.367
R988 B.n582 B.n31 163.367
R989 B.n578 B.n31 163.367
R990 B.n578 B.n577 163.367
R991 B.n577 B.n576 163.367
R992 B.n576 B.n33 163.367
R993 B.n572 B.n33 163.367
R994 B.n572 B.n571 163.367
R995 B.n571 B.n570 163.367
R996 B.n570 B.n35 163.367
R997 B.n566 B.n35 163.367
R998 B.n566 B.n565 163.367
R999 B.n565 B.n564 163.367
R1000 B.n564 B.n37 163.367
R1001 B.n560 B.n37 163.367
R1002 B.n560 B.n559 163.367
R1003 B.n559 B.n558 163.367
R1004 B.n558 B.n39 163.367
R1005 B.n554 B.n39 163.367
R1006 B.n554 B.n553 163.367
R1007 B.n553 B.n552 163.367
R1008 B.n552 B.n41 163.367
R1009 B.n548 B.n41 163.367
R1010 B.n548 B.n547 163.367
R1011 B.n547 B.n546 163.367
R1012 B.n546 B.n46 163.367
R1013 B.n542 B.n46 163.367
R1014 B.n542 B.n541 163.367
R1015 B.n541 B.n540 163.367
R1016 B.n540 B.n48 163.367
R1017 B.n535 B.n48 163.367
R1018 B.n535 B.n534 163.367
R1019 B.n534 B.n533 163.367
R1020 B.n533 B.n52 163.367
R1021 B.n529 B.n52 163.367
R1022 B.n529 B.n528 163.367
R1023 B.n528 B.n527 163.367
R1024 B.n527 B.n54 163.367
R1025 B.n523 B.n54 163.367
R1026 B.n523 B.n522 163.367
R1027 B.n522 B.n521 163.367
R1028 B.n521 B.n56 163.367
R1029 B.n517 B.n56 163.367
R1030 B.n517 B.n516 163.367
R1031 B.n516 B.n515 163.367
R1032 B.n515 B.n58 163.367
R1033 B.n511 B.n58 163.367
R1034 B.n511 B.n510 163.367
R1035 B.n510 B.n509 163.367
R1036 B.n584 B.n583 163.367
R1037 B.n584 B.n29 163.367
R1038 B.n588 B.n29 163.367
R1039 B.n589 B.n588 163.367
R1040 B.n590 B.n589 163.367
R1041 B.n590 B.n27 163.367
R1042 B.n594 B.n27 163.367
R1043 B.n595 B.n594 163.367
R1044 B.n596 B.n595 163.367
R1045 B.n596 B.n25 163.367
R1046 B.n600 B.n25 163.367
R1047 B.n601 B.n600 163.367
R1048 B.n602 B.n601 163.367
R1049 B.n602 B.n23 163.367
R1050 B.n606 B.n23 163.367
R1051 B.n607 B.n606 163.367
R1052 B.n608 B.n607 163.367
R1053 B.n608 B.n21 163.367
R1054 B.n612 B.n21 163.367
R1055 B.n613 B.n612 163.367
R1056 B.n614 B.n613 163.367
R1057 B.n614 B.n19 163.367
R1058 B.n618 B.n19 163.367
R1059 B.n619 B.n618 163.367
R1060 B.n620 B.n619 163.367
R1061 B.n620 B.n17 163.367
R1062 B.n624 B.n17 163.367
R1063 B.n625 B.n624 163.367
R1064 B.n626 B.n625 163.367
R1065 B.n626 B.n15 163.367
R1066 B.n630 B.n15 163.367
R1067 B.n631 B.n630 163.367
R1068 B.n632 B.n631 163.367
R1069 B.n632 B.n13 163.367
R1070 B.n636 B.n13 163.367
R1071 B.n637 B.n636 163.367
R1072 B.n638 B.n637 163.367
R1073 B.n638 B.n11 163.367
R1074 B.n642 B.n11 163.367
R1075 B.n643 B.n642 163.367
R1076 B.n644 B.n643 163.367
R1077 B.n644 B.n9 163.367
R1078 B.n648 B.n9 163.367
R1079 B.n649 B.n648 163.367
R1080 B.n650 B.n649 163.367
R1081 B.n650 B.n7 163.367
R1082 B.n654 B.n7 163.367
R1083 B.n655 B.n654 163.367
R1084 B.n656 B.n655 163.367
R1085 B.n656 B.n5 163.367
R1086 B.n660 B.n5 163.367
R1087 B.n661 B.n660 163.367
R1088 B.n662 B.n661 163.367
R1089 B.n662 B.n3 163.367
R1090 B.n666 B.n3 163.367
R1091 B.n667 B.n666 163.367
R1092 B.n174 B.n2 163.367
R1093 B.n177 B.n174 163.367
R1094 B.n178 B.n177 163.367
R1095 B.n179 B.n178 163.367
R1096 B.n179 B.n172 163.367
R1097 B.n183 B.n172 163.367
R1098 B.n184 B.n183 163.367
R1099 B.n185 B.n184 163.367
R1100 B.n185 B.n170 163.367
R1101 B.n189 B.n170 163.367
R1102 B.n190 B.n189 163.367
R1103 B.n191 B.n190 163.367
R1104 B.n191 B.n168 163.367
R1105 B.n195 B.n168 163.367
R1106 B.n196 B.n195 163.367
R1107 B.n197 B.n196 163.367
R1108 B.n197 B.n166 163.367
R1109 B.n201 B.n166 163.367
R1110 B.n202 B.n201 163.367
R1111 B.n203 B.n202 163.367
R1112 B.n203 B.n164 163.367
R1113 B.n207 B.n164 163.367
R1114 B.n208 B.n207 163.367
R1115 B.n209 B.n208 163.367
R1116 B.n209 B.n162 163.367
R1117 B.n213 B.n162 163.367
R1118 B.n214 B.n213 163.367
R1119 B.n215 B.n214 163.367
R1120 B.n215 B.n160 163.367
R1121 B.n219 B.n160 163.367
R1122 B.n220 B.n219 163.367
R1123 B.n221 B.n220 163.367
R1124 B.n221 B.n158 163.367
R1125 B.n225 B.n158 163.367
R1126 B.n226 B.n225 163.367
R1127 B.n227 B.n226 163.367
R1128 B.n227 B.n156 163.367
R1129 B.n231 B.n156 163.367
R1130 B.n232 B.n231 163.367
R1131 B.n233 B.n232 163.367
R1132 B.n233 B.n154 163.367
R1133 B.n237 B.n154 163.367
R1134 B.n238 B.n237 163.367
R1135 B.n239 B.n238 163.367
R1136 B.n239 B.n152 163.367
R1137 B.n243 B.n152 163.367
R1138 B.n244 B.n243 163.367
R1139 B.n245 B.n244 163.367
R1140 B.n245 B.n150 163.367
R1141 B.n249 B.n150 163.367
R1142 B.n250 B.n249 163.367
R1143 B.n251 B.n250 163.367
R1144 B.n251 B.n148 163.367
R1145 B.n255 B.n148 163.367
R1146 B.n256 B.n255 163.367
R1147 B.n257 B.n256 163.367
R1148 B.n136 B.n135 81.455
R1149 B.n130 B.n129 81.455
R1150 B.n50 B.n49 81.455
R1151 B.n43 B.n42 81.455
R1152 B.n289 B.n136 59.5399
R1153 B.n303 B.n130 59.5399
R1154 B.n538 B.n50 59.5399
R1155 B.n44 B.n43 59.5399
R1156 B.n581 B.n30 32.0005
R1157 B.n508 B.n507 32.0005
R1158 B.n334 B.n333 32.0005
R1159 B.n259 B.n258 32.0005
R1160 B B.n669 18.0485
R1161 B.n585 B.n30 10.6151
R1162 B.n586 B.n585 10.6151
R1163 B.n587 B.n586 10.6151
R1164 B.n587 B.n28 10.6151
R1165 B.n591 B.n28 10.6151
R1166 B.n592 B.n591 10.6151
R1167 B.n593 B.n592 10.6151
R1168 B.n593 B.n26 10.6151
R1169 B.n597 B.n26 10.6151
R1170 B.n598 B.n597 10.6151
R1171 B.n599 B.n598 10.6151
R1172 B.n599 B.n24 10.6151
R1173 B.n603 B.n24 10.6151
R1174 B.n604 B.n603 10.6151
R1175 B.n605 B.n604 10.6151
R1176 B.n605 B.n22 10.6151
R1177 B.n609 B.n22 10.6151
R1178 B.n610 B.n609 10.6151
R1179 B.n611 B.n610 10.6151
R1180 B.n611 B.n20 10.6151
R1181 B.n615 B.n20 10.6151
R1182 B.n616 B.n615 10.6151
R1183 B.n617 B.n616 10.6151
R1184 B.n617 B.n18 10.6151
R1185 B.n621 B.n18 10.6151
R1186 B.n622 B.n621 10.6151
R1187 B.n623 B.n622 10.6151
R1188 B.n623 B.n16 10.6151
R1189 B.n627 B.n16 10.6151
R1190 B.n628 B.n627 10.6151
R1191 B.n629 B.n628 10.6151
R1192 B.n629 B.n14 10.6151
R1193 B.n633 B.n14 10.6151
R1194 B.n634 B.n633 10.6151
R1195 B.n635 B.n634 10.6151
R1196 B.n635 B.n12 10.6151
R1197 B.n639 B.n12 10.6151
R1198 B.n640 B.n639 10.6151
R1199 B.n641 B.n640 10.6151
R1200 B.n641 B.n10 10.6151
R1201 B.n645 B.n10 10.6151
R1202 B.n646 B.n645 10.6151
R1203 B.n647 B.n646 10.6151
R1204 B.n647 B.n8 10.6151
R1205 B.n651 B.n8 10.6151
R1206 B.n652 B.n651 10.6151
R1207 B.n653 B.n652 10.6151
R1208 B.n653 B.n6 10.6151
R1209 B.n657 B.n6 10.6151
R1210 B.n658 B.n657 10.6151
R1211 B.n659 B.n658 10.6151
R1212 B.n659 B.n4 10.6151
R1213 B.n663 B.n4 10.6151
R1214 B.n664 B.n663 10.6151
R1215 B.n665 B.n664 10.6151
R1216 B.n665 B.n0 10.6151
R1217 B.n581 B.n580 10.6151
R1218 B.n580 B.n579 10.6151
R1219 B.n579 B.n32 10.6151
R1220 B.n575 B.n32 10.6151
R1221 B.n575 B.n574 10.6151
R1222 B.n574 B.n573 10.6151
R1223 B.n573 B.n34 10.6151
R1224 B.n569 B.n34 10.6151
R1225 B.n569 B.n568 10.6151
R1226 B.n568 B.n567 10.6151
R1227 B.n567 B.n36 10.6151
R1228 B.n563 B.n36 10.6151
R1229 B.n563 B.n562 10.6151
R1230 B.n562 B.n561 10.6151
R1231 B.n561 B.n38 10.6151
R1232 B.n557 B.n38 10.6151
R1233 B.n557 B.n556 10.6151
R1234 B.n556 B.n555 10.6151
R1235 B.n555 B.n40 10.6151
R1236 B.n551 B.n550 10.6151
R1237 B.n550 B.n549 10.6151
R1238 B.n549 B.n45 10.6151
R1239 B.n545 B.n45 10.6151
R1240 B.n545 B.n544 10.6151
R1241 B.n544 B.n543 10.6151
R1242 B.n543 B.n47 10.6151
R1243 B.n539 B.n47 10.6151
R1244 B.n537 B.n536 10.6151
R1245 B.n536 B.n51 10.6151
R1246 B.n532 B.n51 10.6151
R1247 B.n532 B.n531 10.6151
R1248 B.n531 B.n530 10.6151
R1249 B.n530 B.n53 10.6151
R1250 B.n526 B.n53 10.6151
R1251 B.n526 B.n525 10.6151
R1252 B.n525 B.n524 10.6151
R1253 B.n524 B.n55 10.6151
R1254 B.n520 B.n55 10.6151
R1255 B.n520 B.n519 10.6151
R1256 B.n519 B.n518 10.6151
R1257 B.n518 B.n57 10.6151
R1258 B.n514 B.n57 10.6151
R1259 B.n514 B.n513 10.6151
R1260 B.n513 B.n512 10.6151
R1261 B.n512 B.n59 10.6151
R1262 B.n508 B.n59 10.6151
R1263 B.n507 B.n506 10.6151
R1264 B.n506 B.n61 10.6151
R1265 B.n502 B.n61 10.6151
R1266 B.n502 B.n501 10.6151
R1267 B.n501 B.n500 10.6151
R1268 B.n500 B.n63 10.6151
R1269 B.n496 B.n63 10.6151
R1270 B.n496 B.n495 10.6151
R1271 B.n495 B.n494 10.6151
R1272 B.n494 B.n65 10.6151
R1273 B.n490 B.n65 10.6151
R1274 B.n490 B.n489 10.6151
R1275 B.n489 B.n488 10.6151
R1276 B.n488 B.n67 10.6151
R1277 B.n484 B.n67 10.6151
R1278 B.n484 B.n483 10.6151
R1279 B.n483 B.n482 10.6151
R1280 B.n482 B.n69 10.6151
R1281 B.n478 B.n69 10.6151
R1282 B.n478 B.n477 10.6151
R1283 B.n477 B.n476 10.6151
R1284 B.n476 B.n71 10.6151
R1285 B.n472 B.n71 10.6151
R1286 B.n472 B.n471 10.6151
R1287 B.n471 B.n470 10.6151
R1288 B.n470 B.n73 10.6151
R1289 B.n466 B.n73 10.6151
R1290 B.n466 B.n465 10.6151
R1291 B.n465 B.n464 10.6151
R1292 B.n464 B.n75 10.6151
R1293 B.n460 B.n75 10.6151
R1294 B.n460 B.n459 10.6151
R1295 B.n459 B.n458 10.6151
R1296 B.n458 B.n77 10.6151
R1297 B.n454 B.n77 10.6151
R1298 B.n454 B.n453 10.6151
R1299 B.n453 B.n452 10.6151
R1300 B.n452 B.n79 10.6151
R1301 B.n448 B.n79 10.6151
R1302 B.n448 B.n447 10.6151
R1303 B.n447 B.n446 10.6151
R1304 B.n446 B.n81 10.6151
R1305 B.n442 B.n81 10.6151
R1306 B.n442 B.n441 10.6151
R1307 B.n441 B.n440 10.6151
R1308 B.n440 B.n83 10.6151
R1309 B.n436 B.n83 10.6151
R1310 B.n436 B.n435 10.6151
R1311 B.n435 B.n434 10.6151
R1312 B.n434 B.n85 10.6151
R1313 B.n430 B.n85 10.6151
R1314 B.n430 B.n429 10.6151
R1315 B.n429 B.n428 10.6151
R1316 B.n428 B.n87 10.6151
R1317 B.n424 B.n87 10.6151
R1318 B.n424 B.n423 10.6151
R1319 B.n423 B.n422 10.6151
R1320 B.n422 B.n89 10.6151
R1321 B.n418 B.n89 10.6151
R1322 B.n418 B.n417 10.6151
R1323 B.n417 B.n416 10.6151
R1324 B.n416 B.n91 10.6151
R1325 B.n412 B.n91 10.6151
R1326 B.n412 B.n411 10.6151
R1327 B.n411 B.n410 10.6151
R1328 B.n410 B.n93 10.6151
R1329 B.n406 B.n93 10.6151
R1330 B.n406 B.n405 10.6151
R1331 B.n405 B.n404 10.6151
R1332 B.n404 B.n95 10.6151
R1333 B.n400 B.n95 10.6151
R1334 B.n400 B.n399 10.6151
R1335 B.n399 B.n398 10.6151
R1336 B.n398 B.n97 10.6151
R1337 B.n394 B.n97 10.6151
R1338 B.n394 B.n393 10.6151
R1339 B.n393 B.n392 10.6151
R1340 B.n392 B.n99 10.6151
R1341 B.n388 B.n99 10.6151
R1342 B.n388 B.n387 10.6151
R1343 B.n387 B.n386 10.6151
R1344 B.n386 B.n101 10.6151
R1345 B.n382 B.n101 10.6151
R1346 B.n382 B.n381 10.6151
R1347 B.n381 B.n380 10.6151
R1348 B.n380 B.n103 10.6151
R1349 B.n376 B.n103 10.6151
R1350 B.n376 B.n375 10.6151
R1351 B.n375 B.n374 10.6151
R1352 B.n374 B.n105 10.6151
R1353 B.n370 B.n105 10.6151
R1354 B.n370 B.n369 10.6151
R1355 B.n369 B.n368 10.6151
R1356 B.n368 B.n107 10.6151
R1357 B.n364 B.n107 10.6151
R1358 B.n364 B.n363 10.6151
R1359 B.n363 B.n362 10.6151
R1360 B.n362 B.n109 10.6151
R1361 B.n358 B.n109 10.6151
R1362 B.n358 B.n357 10.6151
R1363 B.n357 B.n356 10.6151
R1364 B.n356 B.n111 10.6151
R1365 B.n352 B.n111 10.6151
R1366 B.n352 B.n351 10.6151
R1367 B.n351 B.n350 10.6151
R1368 B.n350 B.n113 10.6151
R1369 B.n346 B.n113 10.6151
R1370 B.n346 B.n345 10.6151
R1371 B.n345 B.n344 10.6151
R1372 B.n344 B.n115 10.6151
R1373 B.n340 B.n115 10.6151
R1374 B.n340 B.n339 10.6151
R1375 B.n339 B.n338 10.6151
R1376 B.n338 B.n117 10.6151
R1377 B.n334 B.n117 10.6151
R1378 B.n175 B.n1 10.6151
R1379 B.n176 B.n175 10.6151
R1380 B.n176 B.n173 10.6151
R1381 B.n180 B.n173 10.6151
R1382 B.n181 B.n180 10.6151
R1383 B.n182 B.n181 10.6151
R1384 B.n182 B.n171 10.6151
R1385 B.n186 B.n171 10.6151
R1386 B.n187 B.n186 10.6151
R1387 B.n188 B.n187 10.6151
R1388 B.n188 B.n169 10.6151
R1389 B.n192 B.n169 10.6151
R1390 B.n193 B.n192 10.6151
R1391 B.n194 B.n193 10.6151
R1392 B.n194 B.n167 10.6151
R1393 B.n198 B.n167 10.6151
R1394 B.n199 B.n198 10.6151
R1395 B.n200 B.n199 10.6151
R1396 B.n200 B.n165 10.6151
R1397 B.n204 B.n165 10.6151
R1398 B.n205 B.n204 10.6151
R1399 B.n206 B.n205 10.6151
R1400 B.n206 B.n163 10.6151
R1401 B.n210 B.n163 10.6151
R1402 B.n211 B.n210 10.6151
R1403 B.n212 B.n211 10.6151
R1404 B.n212 B.n161 10.6151
R1405 B.n216 B.n161 10.6151
R1406 B.n217 B.n216 10.6151
R1407 B.n218 B.n217 10.6151
R1408 B.n218 B.n159 10.6151
R1409 B.n222 B.n159 10.6151
R1410 B.n223 B.n222 10.6151
R1411 B.n224 B.n223 10.6151
R1412 B.n224 B.n157 10.6151
R1413 B.n228 B.n157 10.6151
R1414 B.n229 B.n228 10.6151
R1415 B.n230 B.n229 10.6151
R1416 B.n230 B.n155 10.6151
R1417 B.n234 B.n155 10.6151
R1418 B.n235 B.n234 10.6151
R1419 B.n236 B.n235 10.6151
R1420 B.n236 B.n153 10.6151
R1421 B.n240 B.n153 10.6151
R1422 B.n241 B.n240 10.6151
R1423 B.n242 B.n241 10.6151
R1424 B.n242 B.n151 10.6151
R1425 B.n246 B.n151 10.6151
R1426 B.n247 B.n246 10.6151
R1427 B.n248 B.n247 10.6151
R1428 B.n248 B.n149 10.6151
R1429 B.n252 B.n149 10.6151
R1430 B.n253 B.n252 10.6151
R1431 B.n254 B.n253 10.6151
R1432 B.n254 B.n147 10.6151
R1433 B.n258 B.n147 10.6151
R1434 B.n260 B.n259 10.6151
R1435 B.n260 B.n145 10.6151
R1436 B.n264 B.n145 10.6151
R1437 B.n265 B.n264 10.6151
R1438 B.n266 B.n265 10.6151
R1439 B.n266 B.n143 10.6151
R1440 B.n270 B.n143 10.6151
R1441 B.n271 B.n270 10.6151
R1442 B.n272 B.n271 10.6151
R1443 B.n272 B.n141 10.6151
R1444 B.n276 B.n141 10.6151
R1445 B.n277 B.n276 10.6151
R1446 B.n278 B.n277 10.6151
R1447 B.n278 B.n139 10.6151
R1448 B.n282 B.n139 10.6151
R1449 B.n283 B.n282 10.6151
R1450 B.n284 B.n283 10.6151
R1451 B.n284 B.n137 10.6151
R1452 B.n288 B.n137 10.6151
R1453 B.n291 B.n290 10.6151
R1454 B.n291 B.n133 10.6151
R1455 B.n295 B.n133 10.6151
R1456 B.n296 B.n295 10.6151
R1457 B.n297 B.n296 10.6151
R1458 B.n297 B.n131 10.6151
R1459 B.n301 B.n131 10.6151
R1460 B.n302 B.n301 10.6151
R1461 B.n304 B.n127 10.6151
R1462 B.n308 B.n127 10.6151
R1463 B.n309 B.n308 10.6151
R1464 B.n310 B.n309 10.6151
R1465 B.n310 B.n125 10.6151
R1466 B.n314 B.n125 10.6151
R1467 B.n315 B.n314 10.6151
R1468 B.n316 B.n315 10.6151
R1469 B.n316 B.n123 10.6151
R1470 B.n320 B.n123 10.6151
R1471 B.n321 B.n320 10.6151
R1472 B.n322 B.n321 10.6151
R1473 B.n322 B.n121 10.6151
R1474 B.n326 B.n121 10.6151
R1475 B.n327 B.n326 10.6151
R1476 B.n328 B.n327 10.6151
R1477 B.n328 B.n119 10.6151
R1478 B.n332 B.n119 10.6151
R1479 B.n333 B.n332 10.6151
R1480 B.n669 B.n0 8.11757
R1481 B.n669 B.n1 8.11757
R1482 B.n551 B.n44 6.5566
R1483 B.n539 B.n538 6.5566
R1484 B.n290 B.n289 6.5566
R1485 B.n303 B.n302 6.5566
R1486 B.n44 B.n40 4.05904
R1487 B.n538 B.n537 4.05904
R1488 B.n289 B.n288 4.05904
R1489 B.n304 B.n303 4.05904
C0 w_n4330_n1874# VN 8.389589f
C1 B VDD1 1.81823f
C2 B VTAIL 2.33107f
C3 w_n4330_n1874# VDD1 2.08927f
C4 VDD2 VN 2.95885f
C5 VP VN 6.7863f
C6 w_n4330_n1874# VTAIL 2.07228f
C7 VDD2 VDD1 1.90251f
C8 VP VDD1 3.36972f
C9 VDD2 VTAIL 5.8951f
C10 VP VTAIL 4.02808f
C11 B w_n4330_n1874# 9.36026f
C12 VN VDD1 0.156539f
C13 VN VTAIL 4.0137f
C14 B VDD2 1.92296f
C15 VP B 2.32492f
C16 VTAIL VDD1 5.83361f
C17 w_n4330_n1874# VDD2 2.21463f
C18 VP w_n4330_n1874# 8.952731f
C19 B VN 1.37806f
C20 VP VDD2 0.569979f
C21 VDD2 VSUBS 1.884245f
C22 VDD1 VSUBS 2.036315f
C23 VTAIL VSUBS 0.78966f
C24 VN VSUBS 6.95462f
C25 VP VSUBS 3.393653f
C26 B VSUBS 4.947911f
C27 w_n4330_n1874# VSUBS 0.101894p
C28 B.n0 VSUBS 0.008598f
C29 B.n1 VSUBS 0.008598f
C30 B.n2 VSUBS 0.012716f
C31 B.n3 VSUBS 0.009745f
C32 B.n4 VSUBS 0.009745f
C33 B.n5 VSUBS 0.009745f
C34 B.n6 VSUBS 0.009745f
C35 B.n7 VSUBS 0.009745f
C36 B.n8 VSUBS 0.009745f
C37 B.n9 VSUBS 0.009745f
C38 B.n10 VSUBS 0.009745f
C39 B.n11 VSUBS 0.009745f
C40 B.n12 VSUBS 0.009745f
C41 B.n13 VSUBS 0.009745f
C42 B.n14 VSUBS 0.009745f
C43 B.n15 VSUBS 0.009745f
C44 B.n16 VSUBS 0.009745f
C45 B.n17 VSUBS 0.009745f
C46 B.n18 VSUBS 0.009745f
C47 B.n19 VSUBS 0.009745f
C48 B.n20 VSUBS 0.009745f
C49 B.n21 VSUBS 0.009745f
C50 B.n22 VSUBS 0.009745f
C51 B.n23 VSUBS 0.009745f
C52 B.n24 VSUBS 0.009745f
C53 B.n25 VSUBS 0.009745f
C54 B.n26 VSUBS 0.009745f
C55 B.n27 VSUBS 0.009745f
C56 B.n28 VSUBS 0.009745f
C57 B.n29 VSUBS 0.009745f
C58 B.n30 VSUBS 0.021854f
C59 B.n31 VSUBS 0.009745f
C60 B.n32 VSUBS 0.009745f
C61 B.n33 VSUBS 0.009745f
C62 B.n34 VSUBS 0.009745f
C63 B.n35 VSUBS 0.009745f
C64 B.n36 VSUBS 0.009745f
C65 B.n37 VSUBS 0.009745f
C66 B.n38 VSUBS 0.009745f
C67 B.n39 VSUBS 0.009745f
C68 B.n40 VSUBS 0.006735f
C69 B.n41 VSUBS 0.009745f
C70 B.t1 VSUBS 0.090882f
C71 B.t2 VSUBS 0.133791f
C72 B.t0 VSUBS 1.18479f
C73 B.n42 VSUBS 0.224765f
C74 B.n43 VSUBS 0.184812f
C75 B.n44 VSUBS 0.022577f
C76 B.n45 VSUBS 0.009745f
C77 B.n46 VSUBS 0.009745f
C78 B.n47 VSUBS 0.009745f
C79 B.n48 VSUBS 0.009745f
C80 B.t10 VSUBS 0.090884f
C81 B.t11 VSUBS 0.133793f
C82 B.t9 VSUBS 1.18479f
C83 B.n49 VSUBS 0.224763f
C84 B.n50 VSUBS 0.18481f
C85 B.n51 VSUBS 0.009745f
C86 B.n52 VSUBS 0.009745f
C87 B.n53 VSUBS 0.009745f
C88 B.n54 VSUBS 0.009745f
C89 B.n55 VSUBS 0.009745f
C90 B.n56 VSUBS 0.009745f
C91 B.n57 VSUBS 0.009745f
C92 B.n58 VSUBS 0.009745f
C93 B.n59 VSUBS 0.009745f
C94 B.n60 VSUBS 0.021854f
C95 B.n61 VSUBS 0.009745f
C96 B.n62 VSUBS 0.009745f
C97 B.n63 VSUBS 0.009745f
C98 B.n64 VSUBS 0.009745f
C99 B.n65 VSUBS 0.009745f
C100 B.n66 VSUBS 0.009745f
C101 B.n67 VSUBS 0.009745f
C102 B.n68 VSUBS 0.009745f
C103 B.n69 VSUBS 0.009745f
C104 B.n70 VSUBS 0.009745f
C105 B.n71 VSUBS 0.009745f
C106 B.n72 VSUBS 0.009745f
C107 B.n73 VSUBS 0.009745f
C108 B.n74 VSUBS 0.009745f
C109 B.n75 VSUBS 0.009745f
C110 B.n76 VSUBS 0.009745f
C111 B.n77 VSUBS 0.009745f
C112 B.n78 VSUBS 0.009745f
C113 B.n79 VSUBS 0.009745f
C114 B.n80 VSUBS 0.009745f
C115 B.n81 VSUBS 0.009745f
C116 B.n82 VSUBS 0.009745f
C117 B.n83 VSUBS 0.009745f
C118 B.n84 VSUBS 0.009745f
C119 B.n85 VSUBS 0.009745f
C120 B.n86 VSUBS 0.009745f
C121 B.n87 VSUBS 0.009745f
C122 B.n88 VSUBS 0.009745f
C123 B.n89 VSUBS 0.009745f
C124 B.n90 VSUBS 0.009745f
C125 B.n91 VSUBS 0.009745f
C126 B.n92 VSUBS 0.009745f
C127 B.n93 VSUBS 0.009745f
C128 B.n94 VSUBS 0.009745f
C129 B.n95 VSUBS 0.009745f
C130 B.n96 VSUBS 0.009745f
C131 B.n97 VSUBS 0.009745f
C132 B.n98 VSUBS 0.009745f
C133 B.n99 VSUBS 0.009745f
C134 B.n100 VSUBS 0.009745f
C135 B.n101 VSUBS 0.009745f
C136 B.n102 VSUBS 0.009745f
C137 B.n103 VSUBS 0.009745f
C138 B.n104 VSUBS 0.009745f
C139 B.n105 VSUBS 0.009745f
C140 B.n106 VSUBS 0.009745f
C141 B.n107 VSUBS 0.009745f
C142 B.n108 VSUBS 0.009745f
C143 B.n109 VSUBS 0.009745f
C144 B.n110 VSUBS 0.009745f
C145 B.n111 VSUBS 0.009745f
C146 B.n112 VSUBS 0.009745f
C147 B.n113 VSUBS 0.009745f
C148 B.n114 VSUBS 0.009745f
C149 B.n115 VSUBS 0.009745f
C150 B.n116 VSUBS 0.009745f
C151 B.n117 VSUBS 0.009745f
C152 B.n118 VSUBS 0.023144f
C153 B.n119 VSUBS 0.009745f
C154 B.n120 VSUBS 0.009745f
C155 B.n121 VSUBS 0.009745f
C156 B.n122 VSUBS 0.009745f
C157 B.n123 VSUBS 0.009745f
C158 B.n124 VSUBS 0.009745f
C159 B.n125 VSUBS 0.009745f
C160 B.n126 VSUBS 0.009745f
C161 B.n127 VSUBS 0.009745f
C162 B.n128 VSUBS 0.009745f
C163 B.t8 VSUBS 0.090884f
C164 B.t7 VSUBS 0.133793f
C165 B.t6 VSUBS 1.18479f
C166 B.n129 VSUBS 0.224763f
C167 B.n130 VSUBS 0.18481f
C168 B.n131 VSUBS 0.009745f
C169 B.n132 VSUBS 0.009745f
C170 B.n133 VSUBS 0.009745f
C171 B.n134 VSUBS 0.009745f
C172 B.t5 VSUBS 0.090882f
C173 B.t4 VSUBS 0.133791f
C174 B.t3 VSUBS 1.18479f
C175 B.n135 VSUBS 0.224765f
C176 B.n136 VSUBS 0.184812f
C177 B.n137 VSUBS 0.009745f
C178 B.n138 VSUBS 0.009745f
C179 B.n139 VSUBS 0.009745f
C180 B.n140 VSUBS 0.009745f
C181 B.n141 VSUBS 0.009745f
C182 B.n142 VSUBS 0.009745f
C183 B.n143 VSUBS 0.009745f
C184 B.n144 VSUBS 0.009745f
C185 B.n145 VSUBS 0.009745f
C186 B.n146 VSUBS 0.023144f
C187 B.n147 VSUBS 0.009745f
C188 B.n148 VSUBS 0.009745f
C189 B.n149 VSUBS 0.009745f
C190 B.n150 VSUBS 0.009745f
C191 B.n151 VSUBS 0.009745f
C192 B.n152 VSUBS 0.009745f
C193 B.n153 VSUBS 0.009745f
C194 B.n154 VSUBS 0.009745f
C195 B.n155 VSUBS 0.009745f
C196 B.n156 VSUBS 0.009745f
C197 B.n157 VSUBS 0.009745f
C198 B.n158 VSUBS 0.009745f
C199 B.n159 VSUBS 0.009745f
C200 B.n160 VSUBS 0.009745f
C201 B.n161 VSUBS 0.009745f
C202 B.n162 VSUBS 0.009745f
C203 B.n163 VSUBS 0.009745f
C204 B.n164 VSUBS 0.009745f
C205 B.n165 VSUBS 0.009745f
C206 B.n166 VSUBS 0.009745f
C207 B.n167 VSUBS 0.009745f
C208 B.n168 VSUBS 0.009745f
C209 B.n169 VSUBS 0.009745f
C210 B.n170 VSUBS 0.009745f
C211 B.n171 VSUBS 0.009745f
C212 B.n172 VSUBS 0.009745f
C213 B.n173 VSUBS 0.009745f
C214 B.n174 VSUBS 0.009745f
C215 B.n175 VSUBS 0.009745f
C216 B.n176 VSUBS 0.009745f
C217 B.n177 VSUBS 0.009745f
C218 B.n178 VSUBS 0.009745f
C219 B.n179 VSUBS 0.009745f
C220 B.n180 VSUBS 0.009745f
C221 B.n181 VSUBS 0.009745f
C222 B.n182 VSUBS 0.009745f
C223 B.n183 VSUBS 0.009745f
C224 B.n184 VSUBS 0.009745f
C225 B.n185 VSUBS 0.009745f
C226 B.n186 VSUBS 0.009745f
C227 B.n187 VSUBS 0.009745f
C228 B.n188 VSUBS 0.009745f
C229 B.n189 VSUBS 0.009745f
C230 B.n190 VSUBS 0.009745f
C231 B.n191 VSUBS 0.009745f
C232 B.n192 VSUBS 0.009745f
C233 B.n193 VSUBS 0.009745f
C234 B.n194 VSUBS 0.009745f
C235 B.n195 VSUBS 0.009745f
C236 B.n196 VSUBS 0.009745f
C237 B.n197 VSUBS 0.009745f
C238 B.n198 VSUBS 0.009745f
C239 B.n199 VSUBS 0.009745f
C240 B.n200 VSUBS 0.009745f
C241 B.n201 VSUBS 0.009745f
C242 B.n202 VSUBS 0.009745f
C243 B.n203 VSUBS 0.009745f
C244 B.n204 VSUBS 0.009745f
C245 B.n205 VSUBS 0.009745f
C246 B.n206 VSUBS 0.009745f
C247 B.n207 VSUBS 0.009745f
C248 B.n208 VSUBS 0.009745f
C249 B.n209 VSUBS 0.009745f
C250 B.n210 VSUBS 0.009745f
C251 B.n211 VSUBS 0.009745f
C252 B.n212 VSUBS 0.009745f
C253 B.n213 VSUBS 0.009745f
C254 B.n214 VSUBS 0.009745f
C255 B.n215 VSUBS 0.009745f
C256 B.n216 VSUBS 0.009745f
C257 B.n217 VSUBS 0.009745f
C258 B.n218 VSUBS 0.009745f
C259 B.n219 VSUBS 0.009745f
C260 B.n220 VSUBS 0.009745f
C261 B.n221 VSUBS 0.009745f
C262 B.n222 VSUBS 0.009745f
C263 B.n223 VSUBS 0.009745f
C264 B.n224 VSUBS 0.009745f
C265 B.n225 VSUBS 0.009745f
C266 B.n226 VSUBS 0.009745f
C267 B.n227 VSUBS 0.009745f
C268 B.n228 VSUBS 0.009745f
C269 B.n229 VSUBS 0.009745f
C270 B.n230 VSUBS 0.009745f
C271 B.n231 VSUBS 0.009745f
C272 B.n232 VSUBS 0.009745f
C273 B.n233 VSUBS 0.009745f
C274 B.n234 VSUBS 0.009745f
C275 B.n235 VSUBS 0.009745f
C276 B.n236 VSUBS 0.009745f
C277 B.n237 VSUBS 0.009745f
C278 B.n238 VSUBS 0.009745f
C279 B.n239 VSUBS 0.009745f
C280 B.n240 VSUBS 0.009745f
C281 B.n241 VSUBS 0.009745f
C282 B.n242 VSUBS 0.009745f
C283 B.n243 VSUBS 0.009745f
C284 B.n244 VSUBS 0.009745f
C285 B.n245 VSUBS 0.009745f
C286 B.n246 VSUBS 0.009745f
C287 B.n247 VSUBS 0.009745f
C288 B.n248 VSUBS 0.009745f
C289 B.n249 VSUBS 0.009745f
C290 B.n250 VSUBS 0.009745f
C291 B.n251 VSUBS 0.009745f
C292 B.n252 VSUBS 0.009745f
C293 B.n253 VSUBS 0.009745f
C294 B.n254 VSUBS 0.009745f
C295 B.n255 VSUBS 0.009745f
C296 B.n256 VSUBS 0.009745f
C297 B.n257 VSUBS 0.021854f
C298 B.n258 VSUBS 0.021854f
C299 B.n259 VSUBS 0.023144f
C300 B.n260 VSUBS 0.009745f
C301 B.n261 VSUBS 0.009745f
C302 B.n262 VSUBS 0.009745f
C303 B.n263 VSUBS 0.009745f
C304 B.n264 VSUBS 0.009745f
C305 B.n265 VSUBS 0.009745f
C306 B.n266 VSUBS 0.009745f
C307 B.n267 VSUBS 0.009745f
C308 B.n268 VSUBS 0.009745f
C309 B.n269 VSUBS 0.009745f
C310 B.n270 VSUBS 0.009745f
C311 B.n271 VSUBS 0.009745f
C312 B.n272 VSUBS 0.009745f
C313 B.n273 VSUBS 0.009745f
C314 B.n274 VSUBS 0.009745f
C315 B.n275 VSUBS 0.009745f
C316 B.n276 VSUBS 0.009745f
C317 B.n277 VSUBS 0.009745f
C318 B.n278 VSUBS 0.009745f
C319 B.n279 VSUBS 0.009745f
C320 B.n280 VSUBS 0.009745f
C321 B.n281 VSUBS 0.009745f
C322 B.n282 VSUBS 0.009745f
C323 B.n283 VSUBS 0.009745f
C324 B.n284 VSUBS 0.009745f
C325 B.n285 VSUBS 0.009745f
C326 B.n286 VSUBS 0.009745f
C327 B.n287 VSUBS 0.009745f
C328 B.n288 VSUBS 0.006735f
C329 B.n289 VSUBS 0.022577f
C330 B.n290 VSUBS 0.007882f
C331 B.n291 VSUBS 0.009745f
C332 B.n292 VSUBS 0.009745f
C333 B.n293 VSUBS 0.009745f
C334 B.n294 VSUBS 0.009745f
C335 B.n295 VSUBS 0.009745f
C336 B.n296 VSUBS 0.009745f
C337 B.n297 VSUBS 0.009745f
C338 B.n298 VSUBS 0.009745f
C339 B.n299 VSUBS 0.009745f
C340 B.n300 VSUBS 0.009745f
C341 B.n301 VSUBS 0.009745f
C342 B.n302 VSUBS 0.007882f
C343 B.n303 VSUBS 0.022577f
C344 B.n304 VSUBS 0.006735f
C345 B.n305 VSUBS 0.009745f
C346 B.n306 VSUBS 0.009745f
C347 B.n307 VSUBS 0.009745f
C348 B.n308 VSUBS 0.009745f
C349 B.n309 VSUBS 0.009745f
C350 B.n310 VSUBS 0.009745f
C351 B.n311 VSUBS 0.009745f
C352 B.n312 VSUBS 0.009745f
C353 B.n313 VSUBS 0.009745f
C354 B.n314 VSUBS 0.009745f
C355 B.n315 VSUBS 0.009745f
C356 B.n316 VSUBS 0.009745f
C357 B.n317 VSUBS 0.009745f
C358 B.n318 VSUBS 0.009745f
C359 B.n319 VSUBS 0.009745f
C360 B.n320 VSUBS 0.009745f
C361 B.n321 VSUBS 0.009745f
C362 B.n322 VSUBS 0.009745f
C363 B.n323 VSUBS 0.009745f
C364 B.n324 VSUBS 0.009745f
C365 B.n325 VSUBS 0.009745f
C366 B.n326 VSUBS 0.009745f
C367 B.n327 VSUBS 0.009745f
C368 B.n328 VSUBS 0.009745f
C369 B.n329 VSUBS 0.009745f
C370 B.n330 VSUBS 0.009745f
C371 B.n331 VSUBS 0.009745f
C372 B.n332 VSUBS 0.009745f
C373 B.n333 VSUBS 0.021969f
C374 B.n334 VSUBS 0.023029f
C375 B.n335 VSUBS 0.021854f
C376 B.n336 VSUBS 0.009745f
C377 B.n337 VSUBS 0.009745f
C378 B.n338 VSUBS 0.009745f
C379 B.n339 VSUBS 0.009745f
C380 B.n340 VSUBS 0.009745f
C381 B.n341 VSUBS 0.009745f
C382 B.n342 VSUBS 0.009745f
C383 B.n343 VSUBS 0.009745f
C384 B.n344 VSUBS 0.009745f
C385 B.n345 VSUBS 0.009745f
C386 B.n346 VSUBS 0.009745f
C387 B.n347 VSUBS 0.009745f
C388 B.n348 VSUBS 0.009745f
C389 B.n349 VSUBS 0.009745f
C390 B.n350 VSUBS 0.009745f
C391 B.n351 VSUBS 0.009745f
C392 B.n352 VSUBS 0.009745f
C393 B.n353 VSUBS 0.009745f
C394 B.n354 VSUBS 0.009745f
C395 B.n355 VSUBS 0.009745f
C396 B.n356 VSUBS 0.009745f
C397 B.n357 VSUBS 0.009745f
C398 B.n358 VSUBS 0.009745f
C399 B.n359 VSUBS 0.009745f
C400 B.n360 VSUBS 0.009745f
C401 B.n361 VSUBS 0.009745f
C402 B.n362 VSUBS 0.009745f
C403 B.n363 VSUBS 0.009745f
C404 B.n364 VSUBS 0.009745f
C405 B.n365 VSUBS 0.009745f
C406 B.n366 VSUBS 0.009745f
C407 B.n367 VSUBS 0.009745f
C408 B.n368 VSUBS 0.009745f
C409 B.n369 VSUBS 0.009745f
C410 B.n370 VSUBS 0.009745f
C411 B.n371 VSUBS 0.009745f
C412 B.n372 VSUBS 0.009745f
C413 B.n373 VSUBS 0.009745f
C414 B.n374 VSUBS 0.009745f
C415 B.n375 VSUBS 0.009745f
C416 B.n376 VSUBS 0.009745f
C417 B.n377 VSUBS 0.009745f
C418 B.n378 VSUBS 0.009745f
C419 B.n379 VSUBS 0.009745f
C420 B.n380 VSUBS 0.009745f
C421 B.n381 VSUBS 0.009745f
C422 B.n382 VSUBS 0.009745f
C423 B.n383 VSUBS 0.009745f
C424 B.n384 VSUBS 0.009745f
C425 B.n385 VSUBS 0.009745f
C426 B.n386 VSUBS 0.009745f
C427 B.n387 VSUBS 0.009745f
C428 B.n388 VSUBS 0.009745f
C429 B.n389 VSUBS 0.009745f
C430 B.n390 VSUBS 0.009745f
C431 B.n391 VSUBS 0.009745f
C432 B.n392 VSUBS 0.009745f
C433 B.n393 VSUBS 0.009745f
C434 B.n394 VSUBS 0.009745f
C435 B.n395 VSUBS 0.009745f
C436 B.n396 VSUBS 0.009745f
C437 B.n397 VSUBS 0.009745f
C438 B.n398 VSUBS 0.009745f
C439 B.n399 VSUBS 0.009745f
C440 B.n400 VSUBS 0.009745f
C441 B.n401 VSUBS 0.009745f
C442 B.n402 VSUBS 0.009745f
C443 B.n403 VSUBS 0.009745f
C444 B.n404 VSUBS 0.009745f
C445 B.n405 VSUBS 0.009745f
C446 B.n406 VSUBS 0.009745f
C447 B.n407 VSUBS 0.009745f
C448 B.n408 VSUBS 0.009745f
C449 B.n409 VSUBS 0.009745f
C450 B.n410 VSUBS 0.009745f
C451 B.n411 VSUBS 0.009745f
C452 B.n412 VSUBS 0.009745f
C453 B.n413 VSUBS 0.009745f
C454 B.n414 VSUBS 0.009745f
C455 B.n415 VSUBS 0.009745f
C456 B.n416 VSUBS 0.009745f
C457 B.n417 VSUBS 0.009745f
C458 B.n418 VSUBS 0.009745f
C459 B.n419 VSUBS 0.009745f
C460 B.n420 VSUBS 0.009745f
C461 B.n421 VSUBS 0.009745f
C462 B.n422 VSUBS 0.009745f
C463 B.n423 VSUBS 0.009745f
C464 B.n424 VSUBS 0.009745f
C465 B.n425 VSUBS 0.009745f
C466 B.n426 VSUBS 0.009745f
C467 B.n427 VSUBS 0.009745f
C468 B.n428 VSUBS 0.009745f
C469 B.n429 VSUBS 0.009745f
C470 B.n430 VSUBS 0.009745f
C471 B.n431 VSUBS 0.009745f
C472 B.n432 VSUBS 0.009745f
C473 B.n433 VSUBS 0.009745f
C474 B.n434 VSUBS 0.009745f
C475 B.n435 VSUBS 0.009745f
C476 B.n436 VSUBS 0.009745f
C477 B.n437 VSUBS 0.009745f
C478 B.n438 VSUBS 0.009745f
C479 B.n439 VSUBS 0.009745f
C480 B.n440 VSUBS 0.009745f
C481 B.n441 VSUBS 0.009745f
C482 B.n442 VSUBS 0.009745f
C483 B.n443 VSUBS 0.009745f
C484 B.n444 VSUBS 0.009745f
C485 B.n445 VSUBS 0.009745f
C486 B.n446 VSUBS 0.009745f
C487 B.n447 VSUBS 0.009745f
C488 B.n448 VSUBS 0.009745f
C489 B.n449 VSUBS 0.009745f
C490 B.n450 VSUBS 0.009745f
C491 B.n451 VSUBS 0.009745f
C492 B.n452 VSUBS 0.009745f
C493 B.n453 VSUBS 0.009745f
C494 B.n454 VSUBS 0.009745f
C495 B.n455 VSUBS 0.009745f
C496 B.n456 VSUBS 0.009745f
C497 B.n457 VSUBS 0.009745f
C498 B.n458 VSUBS 0.009745f
C499 B.n459 VSUBS 0.009745f
C500 B.n460 VSUBS 0.009745f
C501 B.n461 VSUBS 0.009745f
C502 B.n462 VSUBS 0.009745f
C503 B.n463 VSUBS 0.009745f
C504 B.n464 VSUBS 0.009745f
C505 B.n465 VSUBS 0.009745f
C506 B.n466 VSUBS 0.009745f
C507 B.n467 VSUBS 0.009745f
C508 B.n468 VSUBS 0.009745f
C509 B.n469 VSUBS 0.009745f
C510 B.n470 VSUBS 0.009745f
C511 B.n471 VSUBS 0.009745f
C512 B.n472 VSUBS 0.009745f
C513 B.n473 VSUBS 0.009745f
C514 B.n474 VSUBS 0.009745f
C515 B.n475 VSUBS 0.009745f
C516 B.n476 VSUBS 0.009745f
C517 B.n477 VSUBS 0.009745f
C518 B.n478 VSUBS 0.009745f
C519 B.n479 VSUBS 0.009745f
C520 B.n480 VSUBS 0.009745f
C521 B.n481 VSUBS 0.009745f
C522 B.n482 VSUBS 0.009745f
C523 B.n483 VSUBS 0.009745f
C524 B.n484 VSUBS 0.009745f
C525 B.n485 VSUBS 0.009745f
C526 B.n486 VSUBS 0.009745f
C527 B.n487 VSUBS 0.009745f
C528 B.n488 VSUBS 0.009745f
C529 B.n489 VSUBS 0.009745f
C530 B.n490 VSUBS 0.009745f
C531 B.n491 VSUBS 0.009745f
C532 B.n492 VSUBS 0.009745f
C533 B.n493 VSUBS 0.009745f
C534 B.n494 VSUBS 0.009745f
C535 B.n495 VSUBS 0.009745f
C536 B.n496 VSUBS 0.009745f
C537 B.n497 VSUBS 0.009745f
C538 B.n498 VSUBS 0.009745f
C539 B.n499 VSUBS 0.009745f
C540 B.n500 VSUBS 0.009745f
C541 B.n501 VSUBS 0.009745f
C542 B.n502 VSUBS 0.009745f
C543 B.n503 VSUBS 0.009745f
C544 B.n504 VSUBS 0.009745f
C545 B.n505 VSUBS 0.009745f
C546 B.n506 VSUBS 0.009745f
C547 B.n507 VSUBS 0.021854f
C548 B.n508 VSUBS 0.023144f
C549 B.n509 VSUBS 0.023144f
C550 B.n510 VSUBS 0.009745f
C551 B.n511 VSUBS 0.009745f
C552 B.n512 VSUBS 0.009745f
C553 B.n513 VSUBS 0.009745f
C554 B.n514 VSUBS 0.009745f
C555 B.n515 VSUBS 0.009745f
C556 B.n516 VSUBS 0.009745f
C557 B.n517 VSUBS 0.009745f
C558 B.n518 VSUBS 0.009745f
C559 B.n519 VSUBS 0.009745f
C560 B.n520 VSUBS 0.009745f
C561 B.n521 VSUBS 0.009745f
C562 B.n522 VSUBS 0.009745f
C563 B.n523 VSUBS 0.009745f
C564 B.n524 VSUBS 0.009745f
C565 B.n525 VSUBS 0.009745f
C566 B.n526 VSUBS 0.009745f
C567 B.n527 VSUBS 0.009745f
C568 B.n528 VSUBS 0.009745f
C569 B.n529 VSUBS 0.009745f
C570 B.n530 VSUBS 0.009745f
C571 B.n531 VSUBS 0.009745f
C572 B.n532 VSUBS 0.009745f
C573 B.n533 VSUBS 0.009745f
C574 B.n534 VSUBS 0.009745f
C575 B.n535 VSUBS 0.009745f
C576 B.n536 VSUBS 0.009745f
C577 B.n537 VSUBS 0.006735f
C578 B.n538 VSUBS 0.022577f
C579 B.n539 VSUBS 0.007882f
C580 B.n540 VSUBS 0.009745f
C581 B.n541 VSUBS 0.009745f
C582 B.n542 VSUBS 0.009745f
C583 B.n543 VSUBS 0.009745f
C584 B.n544 VSUBS 0.009745f
C585 B.n545 VSUBS 0.009745f
C586 B.n546 VSUBS 0.009745f
C587 B.n547 VSUBS 0.009745f
C588 B.n548 VSUBS 0.009745f
C589 B.n549 VSUBS 0.009745f
C590 B.n550 VSUBS 0.009745f
C591 B.n551 VSUBS 0.007882f
C592 B.n552 VSUBS 0.009745f
C593 B.n553 VSUBS 0.009745f
C594 B.n554 VSUBS 0.009745f
C595 B.n555 VSUBS 0.009745f
C596 B.n556 VSUBS 0.009745f
C597 B.n557 VSUBS 0.009745f
C598 B.n558 VSUBS 0.009745f
C599 B.n559 VSUBS 0.009745f
C600 B.n560 VSUBS 0.009745f
C601 B.n561 VSUBS 0.009745f
C602 B.n562 VSUBS 0.009745f
C603 B.n563 VSUBS 0.009745f
C604 B.n564 VSUBS 0.009745f
C605 B.n565 VSUBS 0.009745f
C606 B.n566 VSUBS 0.009745f
C607 B.n567 VSUBS 0.009745f
C608 B.n568 VSUBS 0.009745f
C609 B.n569 VSUBS 0.009745f
C610 B.n570 VSUBS 0.009745f
C611 B.n571 VSUBS 0.009745f
C612 B.n572 VSUBS 0.009745f
C613 B.n573 VSUBS 0.009745f
C614 B.n574 VSUBS 0.009745f
C615 B.n575 VSUBS 0.009745f
C616 B.n576 VSUBS 0.009745f
C617 B.n577 VSUBS 0.009745f
C618 B.n578 VSUBS 0.009745f
C619 B.n579 VSUBS 0.009745f
C620 B.n580 VSUBS 0.009745f
C621 B.n581 VSUBS 0.023144f
C622 B.n582 VSUBS 0.023144f
C623 B.n583 VSUBS 0.021854f
C624 B.n584 VSUBS 0.009745f
C625 B.n585 VSUBS 0.009745f
C626 B.n586 VSUBS 0.009745f
C627 B.n587 VSUBS 0.009745f
C628 B.n588 VSUBS 0.009745f
C629 B.n589 VSUBS 0.009745f
C630 B.n590 VSUBS 0.009745f
C631 B.n591 VSUBS 0.009745f
C632 B.n592 VSUBS 0.009745f
C633 B.n593 VSUBS 0.009745f
C634 B.n594 VSUBS 0.009745f
C635 B.n595 VSUBS 0.009745f
C636 B.n596 VSUBS 0.009745f
C637 B.n597 VSUBS 0.009745f
C638 B.n598 VSUBS 0.009745f
C639 B.n599 VSUBS 0.009745f
C640 B.n600 VSUBS 0.009745f
C641 B.n601 VSUBS 0.009745f
C642 B.n602 VSUBS 0.009745f
C643 B.n603 VSUBS 0.009745f
C644 B.n604 VSUBS 0.009745f
C645 B.n605 VSUBS 0.009745f
C646 B.n606 VSUBS 0.009745f
C647 B.n607 VSUBS 0.009745f
C648 B.n608 VSUBS 0.009745f
C649 B.n609 VSUBS 0.009745f
C650 B.n610 VSUBS 0.009745f
C651 B.n611 VSUBS 0.009745f
C652 B.n612 VSUBS 0.009745f
C653 B.n613 VSUBS 0.009745f
C654 B.n614 VSUBS 0.009745f
C655 B.n615 VSUBS 0.009745f
C656 B.n616 VSUBS 0.009745f
C657 B.n617 VSUBS 0.009745f
C658 B.n618 VSUBS 0.009745f
C659 B.n619 VSUBS 0.009745f
C660 B.n620 VSUBS 0.009745f
C661 B.n621 VSUBS 0.009745f
C662 B.n622 VSUBS 0.009745f
C663 B.n623 VSUBS 0.009745f
C664 B.n624 VSUBS 0.009745f
C665 B.n625 VSUBS 0.009745f
C666 B.n626 VSUBS 0.009745f
C667 B.n627 VSUBS 0.009745f
C668 B.n628 VSUBS 0.009745f
C669 B.n629 VSUBS 0.009745f
C670 B.n630 VSUBS 0.009745f
C671 B.n631 VSUBS 0.009745f
C672 B.n632 VSUBS 0.009745f
C673 B.n633 VSUBS 0.009745f
C674 B.n634 VSUBS 0.009745f
C675 B.n635 VSUBS 0.009745f
C676 B.n636 VSUBS 0.009745f
C677 B.n637 VSUBS 0.009745f
C678 B.n638 VSUBS 0.009745f
C679 B.n639 VSUBS 0.009745f
C680 B.n640 VSUBS 0.009745f
C681 B.n641 VSUBS 0.009745f
C682 B.n642 VSUBS 0.009745f
C683 B.n643 VSUBS 0.009745f
C684 B.n644 VSUBS 0.009745f
C685 B.n645 VSUBS 0.009745f
C686 B.n646 VSUBS 0.009745f
C687 B.n647 VSUBS 0.009745f
C688 B.n648 VSUBS 0.009745f
C689 B.n649 VSUBS 0.009745f
C690 B.n650 VSUBS 0.009745f
C691 B.n651 VSUBS 0.009745f
C692 B.n652 VSUBS 0.009745f
C693 B.n653 VSUBS 0.009745f
C694 B.n654 VSUBS 0.009745f
C695 B.n655 VSUBS 0.009745f
C696 B.n656 VSUBS 0.009745f
C697 B.n657 VSUBS 0.009745f
C698 B.n658 VSUBS 0.009745f
C699 B.n659 VSUBS 0.009745f
C700 B.n660 VSUBS 0.009745f
C701 B.n661 VSUBS 0.009745f
C702 B.n662 VSUBS 0.009745f
C703 B.n663 VSUBS 0.009745f
C704 B.n664 VSUBS 0.009745f
C705 B.n665 VSUBS 0.009745f
C706 B.n666 VSUBS 0.009745f
C707 B.n667 VSUBS 0.012716f
C708 B.n668 VSUBS 0.013546f
C709 B.n669 VSUBS 0.026938f
C710 VDD1.n0 VSUBS 0.029324f
C711 VDD1.n1 VSUBS 0.027981f
C712 VDD1.n2 VSUBS 0.015036f
C713 VDD1.n3 VSUBS 0.035539f
C714 VDD1.n4 VSUBS 0.01592f
C715 VDD1.n5 VSUBS 0.453734f
C716 VDD1.n6 VSUBS 0.015036f
C717 VDD1.t2 VSUBS 0.077041f
C718 VDD1.n7 VSUBS 0.112188f
C719 VDD1.n8 VSUBS 0.022515f
C720 VDD1.n9 VSUBS 0.026654f
C721 VDD1.n10 VSUBS 0.035539f
C722 VDD1.n11 VSUBS 0.01592f
C723 VDD1.n12 VSUBS 0.015036f
C724 VDD1.n13 VSUBS 0.027981f
C725 VDD1.n14 VSUBS 0.027981f
C726 VDD1.n15 VSUBS 0.015036f
C727 VDD1.n16 VSUBS 0.01592f
C728 VDD1.n17 VSUBS 0.035539f
C729 VDD1.n18 VSUBS 0.081194f
C730 VDD1.n19 VSUBS 0.01592f
C731 VDD1.n20 VSUBS 0.015036f
C732 VDD1.n21 VSUBS 0.06353f
C733 VDD1.n22 VSUBS 0.076389f
C734 VDD1.n23 VSUBS 0.029324f
C735 VDD1.n24 VSUBS 0.027981f
C736 VDD1.n25 VSUBS 0.015036f
C737 VDD1.n26 VSUBS 0.035539f
C738 VDD1.n27 VSUBS 0.01592f
C739 VDD1.n28 VSUBS 0.453734f
C740 VDD1.n29 VSUBS 0.015036f
C741 VDD1.t5 VSUBS 0.077041f
C742 VDD1.n30 VSUBS 0.112188f
C743 VDD1.n31 VSUBS 0.022515f
C744 VDD1.n32 VSUBS 0.026654f
C745 VDD1.n33 VSUBS 0.035539f
C746 VDD1.n34 VSUBS 0.01592f
C747 VDD1.n35 VSUBS 0.015036f
C748 VDD1.n36 VSUBS 0.027981f
C749 VDD1.n37 VSUBS 0.027981f
C750 VDD1.n38 VSUBS 0.015036f
C751 VDD1.n39 VSUBS 0.01592f
C752 VDD1.n40 VSUBS 0.035539f
C753 VDD1.n41 VSUBS 0.081194f
C754 VDD1.n42 VSUBS 0.01592f
C755 VDD1.n43 VSUBS 0.015036f
C756 VDD1.n44 VSUBS 0.06353f
C757 VDD1.n45 VSUBS 0.075228f
C758 VDD1.t1 VSUBS 0.100165f
C759 VDD1.t3 VSUBS 0.100165f
C760 VDD1.n46 VSUBS 0.616382f
C761 VDD1.n47 VSUBS 3.45248f
C762 VDD1.t0 VSUBS 0.100165f
C763 VDD1.t4 VSUBS 0.100165f
C764 VDD1.n48 VSUBS 0.609624f
C765 VDD1.n49 VSUBS 3.06476f
C766 VP.n0 VSUBS 0.07897f
C767 VP.t2 VSUBS 1.91086f
C768 VP.n1 VSUBS 0.080284f
C769 VP.n2 VSUBS 0.041983f
C770 VP.n3 VSUBS 0.078246f
C771 VP.n4 VSUBS 0.041983f
C772 VP.t4 VSUBS 1.91086f
C773 VP.n5 VSUBS 0.078246f
C774 VP.n6 VSUBS 0.041983f
C775 VP.n7 VSUBS 0.078246f
C776 VP.n8 VSUBS 0.07897f
C777 VP.t1 VSUBS 1.91086f
C778 VP.n9 VSUBS 0.080284f
C779 VP.n10 VSUBS 0.041983f
C780 VP.n11 VSUBS 0.078246f
C781 VP.t3 VSUBS 2.47402f
C782 VP.n12 VSUBS 0.880757f
C783 VP.t5 VSUBS 1.91086f
C784 VP.n13 VSUBS 0.877897f
C785 VP.n14 VSUBS 0.058931f
C786 VP.n15 VSUBS 0.551261f
C787 VP.n16 VSUBS 0.041983f
C788 VP.n17 VSUBS 0.041983f
C789 VP.n18 VSUBS 0.078246f
C790 VP.n19 VSUBS 0.072661f
C791 VP.n20 VSUBS 0.047875f
C792 VP.n21 VSUBS 0.041983f
C793 VP.n22 VSUBS 0.041983f
C794 VP.n23 VSUBS 0.041983f
C795 VP.n24 VSUBS 0.078246f
C796 VP.n25 VSUBS 0.074383f
C797 VP.n26 VSUBS 0.911998f
C798 VP.n27 VSUBS 2.31697f
C799 VP.n28 VSUBS 2.34825f
C800 VP.t0 VSUBS 1.91086f
C801 VP.n29 VSUBS 0.911998f
C802 VP.n30 VSUBS 0.074383f
C803 VP.n31 VSUBS 0.07897f
C804 VP.n32 VSUBS 0.041983f
C805 VP.n33 VSUBS 0.041983f
C806 VP.n34 VSUBS 0.080284f
C807 VP.n35 VSUBS 0.047875f
C808 VP.n36 VSUBS 0.072661f
C809 VP.n37 VSUBS 0.041983f
C810 VP.n38 VSUBS 0.041983f
C811 VP.n39 VSUBS 0.041983f
C812 VP.n40 VSUBS 0.078246f
C813 VP.n41 VSUBS 0.058931f
C814 VP.n42 VSUBS 0.726177f
C815 VP.n43 VSUBS 0.058931f
C816 VP.n44 VSUBS 0.041983f
C817 VP.n45 VSUBS 0.041983f
C818 VP.n46 VSUBS 0.041983f
C819 VP.n47 VSUBS 0.078246f
C820 VP.n48 VSUBS 0.072661f
C821 VP.n49 VSUBS 0.047875f
C822 VP.n50 VSUBS 0.041983f
C823 VP.n51 VSUBS 0.041983f
C824 VP.n52 VSUBS 0.041983f
C825 VP.n53 VSUBS 0.078246f
C826 VP.n54 VSUBS 0.074383f
C827 VP.n55 VSUBS 0.911998f
C828 VP.n56 VSUBS 0.127705f
C829 VTAIL.t7 VSUBS 0.133329f
C830 VTAIL.t6 VSUBS 0.133329f
C831 VTAIL.n0 VSUBS 0.706792f
C832 VTAIL.n1 VSUBS 0.995273f
C833 VTAIL.n2 VSUBS 0.039032f
C834 VTAIL.n3 VSUBS 0.037245f
C835 VTAIL.n4 VSUBS 0.020014f
C836 VTAIL.n5 VSUBS 0.047306f
C837 VTAIL.n6 VSUBS 0.021191f
C838 VTAIL.n7 VSUBS 0.603962f
C839 VTAIL.n8 VSUBS 0.020014f
C840 VTAIL.t11 VSUBS 0.102548f
C841 VTAIL.n9 VSUBS 0.149333f
C842 VTAIL.n10 VSUBS 0.029969f
C843 VTAIL.n11 VSUBS 0.03548f
C844 VTAIL.n12 VSUBS 0.047306f
C845 VTAIL.n13 VSUBS 0.021191f
C846 VTAIL.n14 VSUBS 0.020014f
C847 VTAIL.n15 VSUBS 0.037245f
C848 VTAIL.n16 VSUBS 0.037245f
C849 VTAIL.n17 VSUBS 0.020014f
C850 VTAIL.n18 VSUBS 0.021191f
C851 VTAIL.n19 VSUBS 0.047306f
C852 VTAIL.n20 VSUBS 0.108077f
C853 VTAIL.n21 VSUBS 0.021191f
C854 VTAIL.n22 VSUBS 0.020014f
C855 VTAIL.n23 VSUBS 0.084565f
C856 VTAIL.n24 VSUBS 0.054017f
C857 VTAIL.n25 VSUBS 0.739132f
C858 VTAIL.t10 VSUBS 0.133329f
C859 VTAIL.t2 VSUBS 0.133329f
C860 VTAIL.n26 VSUBS 0.706792f
C861 VTAIL.n27 VSUBS 2.88421f
C862 VTAIL.t4 VSUBS 0.133329f
C863 VTAIL.t9 VSUBS 0.133329f
C864 VTAIL.n28 VSUBS 0.706797f
C865 VTAIL.n29 VSUBS 2.8842f
C866 VTAIL.n30 VSUBS 0.039032f
C867 VTAIL.n31 VSUBS 0.037245f
C868 VTAIL.n32 VSUBS 0.020014f
C869 VTAIL.n33 VSUBS 0.047306f
C870 VTAIL.n34 VSUBS 0.021191f
C871 VTAIL.n35 VSUBS 0.603962f
C872 VTAIL.n36 VSUBS 0.020014f
C873 VTAIL.t8 VSUBS 0.102548f
C874 VTAIL.n37 VSUBS 0.149333f
C875 VTAIL.n38 VSUBS 0.029969f
C876 VTAIL.n39 VSUBS 0.03548f
C877 VTAIL.n40 VSUBS 0.047306f
C878 VTAIL.n41 VSUBS 0.021191f
C879 VTAIL.n42 VSUBS 0.020014f
C880 VTAIL.n43 VSUBS 0.037245f
C881 VTAIL.n44 VSUBS 0.037245f
C882 VTAIL.n45 VSUBS 0.020014f
C883 VTAIL.n46 VSUBS 0.021191f
C884 VTAIL.n47 VSUBS 0.047306f
C885 VTAIL.n48 VSUBS 0.108077f
C886 VTAIL.n49 VSUBS 0.021191f
C887 VTAIL.n50 VSUBS 0.020014f
C888 VTAIL.n51 VSUBS 0.084565f
C889 VTAIL.n52 VSUBS 0.054017f
C890 VTAIL.n53 VSUBS 0.739132f
C891 VTAIL.t1 VSUBS 0.133329f
C892 VTAIL.t3 VSUBS 0.133329f
C893 VTAIL.n54 VSUBS 0.706797f
C894 VTAIL.n55 VSUBS 1.31418f
C895 VTAIL.n56 VSUBS 0.039032f
C896 VTAIL.n57 VSUBS 0.037245f
C897 VTAIL.n58 VSUBS 0.020014f
C898 VTAIL.n59 VSUBS 0.047306f
C899 VTAIL.n60 VSUBS 0.021191f
C900 VTAIL.n61 VSUBS 0.603962f
C901 VTAIL.n62 VSUBS 0.020014f
C902 VTAIL.t0 VSUBS 0.102548f
C903 VTAIL.n63 VSUBS 0.149333f
C904 VTAIL.n64 VSUBS 0.029969f
C905 VTAIL.n65 VSUBS 0.03548f
C906 VTAIL.n66 VSUBS 0.047306f
C907 VTAIL.n67 VSUBS 0.021191f
C908 VTAIL.n68 VSUBS 0.020014f
C909 VTAIL.n69 VSUBS 0.037245f
C910 VTAIL.n70 VSUBS 0.037245f
C911 VTAIL.n71 VSUBS 0.020014f
C912 VTAIL.n72 VSUBS 0.021191f
C913 VTAIL.n73 VSUBS 0.047306f
C914 VTAIL.n74 VSUBS 0.108077f
C915 VTAIL.n75 VSUBS 0.021191f
C916 VTAIL.n76 VSUBS 0.020014f
C917 VTAIL.n77 VSUBS 0.084565f
C918 VTAIL.n78 VSUBS 0.054017f
C919 VTAIL.n79 VSUBS 1.87462f
C920 VTAIL.n80 VSUBS 0.039032f
C921 VTAIL.n81 VSUBS 0.037245f
C922 VTAIL.n82 VSUBS 0.020014f
C923 VTAIL.n83 VSUBS 0.047306f
C924 VTAIL.n84 VSUBS 0.021191f
C925 VTAIL.n85 VSUBS 0.603962f
C926 VTAIL.n86 VSUBS 0.020014f
C927 VTAIL.t5 VSUBS 0.102548f
C928 VTAIL.n87 VSUBS 0.149333f
C929 VTAIL.n88 VSUBS 0.029969f
C930 VTAIL.n89 VSUBS 0.03548f
C931 VTAIL.n90 VSUBS 0.047306f
C932 VTAIL.n91 VSUBS 0.021191f
C933 VTAIL.n92 VSUBS 0.020014f
C934 VTAIL.n93 VSUBS 0.037245f
C935 VTAIL.n94 VSUBS 0.037245f
C936 VTAIL.n95 VSUBS 0.020014f
C937 VTAIL.n96 VSUBS 0.021191f
C938 VTAIL.n97 VSUBS 0.047306f
C939 VTAIL.n98 VSUBS 0.108077f
C940 VTAIL.n99 VSUBS 0.021191f
C941 VTAIL.n100 VSUBS 0.020014f
C942 VTAIL.n101 VSUBS 0.084565f
C943 VTAIL.n102 VSUBS 0.054017f
C944 VTAIL.n103 VSUBS 1.759f
C945 VDD2.n0 VSUBS 0.02907f
C946 VDD2.n1 VSUBS 0.02774f
C947 VDD2.n2 VSUBS 0.014906f
C948 VDD2.n3 VSUBS 0.035232f
C949 VDD2.n4 VSUBS 0.015783f
C950 VDD2.n5 VSUBS 0.449818f
C951 VDD2.n6 VSUBS 0.014906f
C952 VDD2.t5 VSUBS 0.076376f
C953 VDD2.n7 VSUBS 0.11122f
C954 VDD2.n8 VSUBS 0.02232f
C955 VDD2.n9 VSUBS 0.026424f
C956 VDD2.n10 VSUBS 0.035232f
C957 VDD2.n11 VSUBS 0.015783f
C958 VDD2.n12 VSUBS 0.014906f
C959 VDD2.n13 VSUBS 0.02774f
C960 VDD2.n14 VSUBS 0.02774f
C961 VDD2.n15 VSUBS 0.014906f
C962 VDD2.n16 VSUBS 0.015783f
C963 VDD2.n17 VSUBS 0.035232f
C964 VDD2.n18 VSUBS 0.080493f
C965 VDD2.n19 VSUBS 0.015783f
C966 VDD2.n20 VSUBS 0.014906f
C967 VDD2.n21 VSUBS 0.062982f
C968 VDD2.n22 VSUBS 0.074578f
C969 VDD2.t0 VSUBS 0.099301f
C970 VDD2.t1 VSUBS 0.099301f
C971 VDD2.n23 VSUBS 0.611061f
C972 VDD2.n24 VSUBS 3.25694f
C973 VDD2.n25 VSUBS 0.02907f
C974 VDD2.n26 VSUBS 0.02774f
C975 VDD2.n27 VSUBS 0.014906f
C976 VDD2.n28 VSUBS 0.035232f
C977 VDD2.n29 VSUBS 0.015783f
C978 VDD2.n30 VSUBS 0.449818f
C979 VDD2.n31 VSUBS 0.014906f
C980 VDD2.t4 VSUBS 0.076376f
C981 VDD2.n32 VSUBS 0.11122f
C982 VDD2.n33 VSUBS 0.02232f
C983 VDD2.n34 VSUBS 0.026424f
C984 VDD2.n35 VSUBS 0.035232f
C985 VDD2.n36 VSUBS 0.015783f
C986 VDD2.n37 VSUBS 0.014906f
C987 VDD2.n38 VSUBS 0.02774f
C988 VDD2.n39 VSUBS 0.02774f
C989 VDD2.n40 VSUBS 0.014906f
C990 VDD2.n41 VSUBS 0.015783f
C991 VDD2.n42 VSUBS 0.035232f
C992 VDD2.n43 VSUBS 0.080493f
C993 VDD2.n44 VSUBS 0.015783f
C994 VDD2.n45 VSUBS 0.014906f
C995 VDD2.n46 VSUBS 0.062982f
C996 VDD2.n47 VSUBS 0.059394f
C997 VDD2.n48 VSUBS 2.58067f
C998 VDD2.t3 VSUBS 0.099301f
C999 VDD2.t2 VSUBS 0.099301f
C1000 VDD2.n49 VSUBS 0.611031f
C1001 VN.n0 VSUBS 0.068592f
C1002 VN.t4 VSUBS 1.65973f
C1003 VN.n1 VSUBS 0.069733f
C1004 VN.n2 VSUBS 0.036465f
C1005 VN.n3 VSUBS 0.067963f
C1006 VN.t2 VSUBS 2.14888f
C1007 VN.n4 VSUBS 0.765003f
C1008 VN.t3 VSUBS 1.65973f
C1009 VN.n5 VSUBS 0.762522f
C1010 VN.n6 VSUBS 0.051186f
C1011 VN.n7 VSUBS 0.478812f
C1012 VN.n8 VSUBS 0.036465f
C1013 VN.n9 VSUBS 0.036465f
C1014 VN.n10 VSUBS 0.067963f
C1015 VN.n11 VSUBS 0.063112f
C1016 VN.n12 VSUBS 0.041583f
C1017 VN.n13 VSUBS 0.036465f
C1018 VN.n14 VSUBS 0.036465f
C1019 VN.n15 VSUBS 0.036465f
C1020 VN.n16 VSUBS 0.067963f
C1021 VN.n17 VSUBS 0.064607f
C1022 VN.n18 VSUBS 0.792142f
C1023 VN.n19 VSUBS 0.110922f
C1024 VN.n20 VSUBS 0.068592f
C1025 VN.t5 VSUBS 1.65973f
C1026 VN.n21 VSUBS 0.069733f
C1027 VN.n22 VSUBS 0.036465f
C1028 VN.n23 VSUBS 0.067963f
C1029 VN.t1 VSUBS 2.14888f
C1030 VN.n24 VSUBS 0.765003f
C1031 VN.t0 VSUBS 1.65973f
C1032 VN.n25 VSUBS 0.762522f
C1033 VN.n26 VSUBS 0.051186f
C1034 VN.n27 VSUBS 0.478812f
C1035 VN.n28 VSUBS 0.036465f
C1036 VN.n29 VSUBS 0.036465f
C1037 VN.n30 VSUBS 0.067963f
C1038 VN.n31 VSUBS 0.063112f
C1039 VN.n32 VSUBS 0.041583f
C1040 VN.n33 VSUBS 0.036465f
C1041 VN.n34 VSUBS 0.036465f
C1042 VN.n35 VSUBS 0.036465f
C1043 VN.n36 VSUBS 0.067963f
C1044 VN.n37 VSUBS 0.064607f
C1045 VN.n38 VSUBS 0.792142f
C1046 VN.n39 VSUBS 2.02228f
.ends

