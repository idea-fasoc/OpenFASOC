* NGSPICE file created from diff_pair_sample_1762.ext - technology: sky130A

.subckt diff_pair_sample_1762 VTAIL VN VP B VDD2 VDD1
X0 B.t22 B.t20 B.t21 B.t17 sky130_fd_pr__nfet_01v8 ad=1.8135 pd=10.08 as=0 ps=0 w=4.65 l=1.43
X1 VDD2.t9 VN.t0 VTAIL.t15 B.t2 sky130_fd_pr__nfet_01v8 ad=0.76725 pd=4.98 as=1.8135 ps=10.08 w=4.65 l=1.43
X2 B.t19 B.t16 B.t18 B.t17 sky130_fd_pr__nfet_01v8 ad=1.8135 pd=10.08 as=0 ps=0 w=4.65 l=1.43
X3 VTAIL.t1 VP.t0 VDD1.t9 B.t7 sky130_fd_pr__nfet_01v8 ad=0.76725 pd=4.98 as=0.76725 ps=4.98 w=4.65 l=1.43
X4 VDD1.t8 VP.t1 VTAIL.t0 B.t3 sky130_fd_pr__nfet_01v8 ad=1.8135 pd=10.08 as=0.76725 ps=4.98 w=4.65 l=1.43
X5 VDD1.t7 VP.t2 VTAIL.t4 B.t1 sky130_fd_pr__nfet_01v8 ad=1.8135 pd=10.08 as=0.76725 ps=4.98 w=4.65 l=1.43
X6 VTAIL.t3 VP.t3 VDD1.t6 B.t0 sky130_fd_pr__nfet_01v8 ad=0.76725 pd=4.98 as=0.76725 ps=4.98 w=4.65 l=1.43
X7 VDD2.t8 VN.t1 VTAIL.t9 B.t23 sky130_fd_pr__nfet_01v8 ad=0.76725 pd=4.98 as=0.76725 ps=4.98 w=4.65 l=1.43
X8 B.t15 B.t13 B.t14 B.t10 sky130_fd_pr__nfet_01v8 ad=1.8135 pd=10.08 as=0 ps=0 w=4.65 l=1.43
X9 VDD1.t5 VP.t4 VTAIL.t17 B.t6 sky130_fd_pr__nfet_01v8 ad=0.76725 pd=4.98 as=1.8135 ps=10.08 w=4.65 l=1.43
X10 VDD1.t4 VP.t5 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=0.76725 pd=4.98 as=1.8135 ps=10.08 w=4.65 l=1.43
X11 VTAIL.t19 VP.t6 VDD1.t3 B.t8 sky130_fd_pr__nfet_01v8 ad=0.76725 pd=4.98 as=0.76725 ps=4.98 w=4.65 l=1.43
X12 VDD1.t2 VP.t7 VTAIL.t5 B.t23 sky130_fd_pr__nfet_01v8 ad=0.76725 pd=4.98 as=0.76725 ps=4.98 w=4.65 l=1.43
X13 VTAIL.t16 VN.t2 VDD2.t7 B.t7 sky130_fd_pr__nfet_01v8 ad=0.76725 pd=4.98 as=0.76725 ps=4.98 w=4.65 l=1.43
X14 VDD2.t6 VN.t3 VTAIL.t7 B.t6 sky130_fd_pr__nfet_01v8 ad=0.76725 pd=4.98 as=1.8135 ps=10.08 w=4.65 l=1.43
X15 B.t12 B.t9 B.t11 B.t10 sky130_fd_pr__nfet_01v8 ad=1.8135 pd=10.08 as=0 ps=0 w=4.65 l=1.43
X16 VDD1.t1 VP.t8 VTAIL.t18 B.t4 sky130_fd_pr__nfet_01v8 ad=0.76725 pd=4.98 as=0.76725 ps=4.98 w=4.65 l=1.43
X17 VTAIL.t10 VN.t4 VDD2.t5 B.t0 sky130_fd_pr__nfet_01v8 ad=0.76725 pd=4.98 as=0.76725 ps=4.98 w=4.65 l=1.43
X18 VTAIL.t11 VN.t5 VDD2.t4 B.t5 sky130_fd_pr__nfet_01v8 ad=0.76725 pd=4.98 as=0.76725 ps=4.98 w=4.65 l=1.43
X19 VTAIL.t6 VP.t9 VDD1.t0 B.t5 sky130_fd_pr__nfet_01v8 ad=0.76725 pd=4.98 as=0.76725 ps=4.98 w=4.65 l=1.43
X20 VDD2.t3 VN.t6 VTAIL.t13 B.t4 sky130_fd_pr__nfet_01v8 ad=0.76725 pd=4.98 as=0.76725 ps=4.98 w=4.65 l=1.43
X21 VTAIL.t14 VN.t7 VDD2.t2 B.t8 sky130_fd_pr__nfet_01v8 ad=0.76725 pd=4.98 as=0.76725 ps=4.98 w=4.65 l=1.43
X22 VDD2.t1 VN.t8 VTAIL.t8 B.t3 sky130_fd_pr__nfet_01v8 ad=1.8135 pd=10.08 as=0.76725 ps=4.98 w=4.65 l=1.43
X23 VDD2.t0 VN.t9 VTAIL.t12 B.t1 sky130_fd_pr__nfet_01v8 ad=1.8135 pd=10.08 as=0.76725 ps=4.98 w=4.65 l=1.43
R0 B.n572 B.n571 585
R1 B.n198 B.n98 585
R2 B.n197 B.n196 585
R3 B.n195 B.n194 585
R4 B.n193 B.n192 585
R5 B.n191 B.n190 585
R6 B.n189 B.n188 585
R7 B.n187 B.n186 585
R8 B.n185 B.n184 585
R9 B.n183 B.n182 585
R10 B.n181 B.n180 585
R11 B.n179 B.n178 585
R12 B.n177 B.n176 585
R13 B.n175 B.n174 585
R14 B.n173 B.n172 585
R15 B.n171 B.n170 585
R16 B.n169 B.n168 585
R17 B.n167 B.n166 585
R18 B.n165 B.n164 585
R19 B.n163 B.n162 585
R20 B.n161 B.n160 585
R21 B.n159 B.n158 585
R22 B.n157 B.n156 585
R23 B.n155 B.n154 585
R24 B.n153 B.n152 585
R25 B.n151 B.n150 585
R26 B.n149 B.n148 585
R27 B.n147 B.n146 585
R28 B.n145 B.n144 585
R29 B.n143 B.n142 585
R30 B.n141 B.n140 585
R31 B.n139 B.n138 585
R32 B.n137 B.n136 585
R33 B.n135 B.n134 585
R34 B.n133 B.n132 585
R35 B.n131 B.n130 585
R36 B.n129 B.n128 585
R37 B.n127 B.n126 585
R38 B.n125 B.n124 585
R39 B.n123 B.n122 585
R40 B.n121 B.n120 585
R41 B.n119 B.n118 585
R42 B.n117 B.n116 585
R43 B.n115 B.n114 585
R44 B.n113 B.n112 585
R45 B.n111 B.n110 585
R46 B.n109 B.n108 585
R47 B.n107 B.n106 585
R48 B.n74 B.n73 585
R49 B.n577 B.n576 585
R50 B.n570 B.n99 585
R51 B.n99 B.n71 585
R52 B.n569 B.n70 585
R53 B.n581 B.n70 585
R54 B.n568 B.n69 585
R55 B.n582 B.n69 585
R56 B.n567 B.n68 585
R57 B.n583 B.n68 585
R58 B.n566 B.n565 585
R59 B.n565 B.n64 585
R60 B.n564 B.n63 585
R61 B.n589 B.n63 585
R62 B.n563 B.n62 585
R63 B.n590 B.n62 585
R64 B.n562 B.n61 585
R65 B.n591 B.n61 585
R66 B.n561 B.n560 585
R67 B.n560 B.n57 585
R68 B.n559 B.n56 585
R69 B.n597 B.n56 585
R70 B.n558 B.n55 585
R71 B.n598 B.n55 585
R72 B.n557 B.n54 585
R73 B.n599 B.n54 585
R74 B.n556 B.n555 585
R75 B.n555 B.n50 585
R76 B.n554 B.n49 585
R77 B.n605 B.n49 585
R78 B.n553 B.n48 585
R79 B.n606 B.n48 585
R80 B.n552 B.n47 585
R81 B.n607 B.n47 585
R82 B.n551 B.n550 585
R83 B.n550 B.n43 585
R84 B.n549 B.n42 585
R85 B.n613 B.n42 585
R86 B.n548 B.n41 585
R87 B.n614 B.n41 585
R88 B.n547 B.n40 585
R89 B.n615 B.n40 585
R90 B.n546 B.n545 585
R91 B.n545 B.n36 585
R92 B.n544 B.n35 585
R93 B.n621 B.n35 585
R94 B.n543 B.n34 585
R95 B.n622 B.n34 585
R96 B.n542 B.n33 585
R97 B.n623 B.n33 585
R98 B.n541 B.n540 585
R99 B.n540 B.n32 585
R100 B.n539 B.n28 585
R101 B.n629 B.n28 585
R102 B.n538 B.n27 585
R103 B.n630 B.n27 585
R104 B.n537 B.n26 585
R105 B.n631 B.n26 585
R106 B.n536 B.n535 585
R107 B.n535 B.n22 585
R108 B.n534 B.n21 585
R109 B.n637 B.n21 585
R110 B.n533 B.n20 585
R111 B.n638 B.n20 585
R112 B.n532 B.n19 585
R113 B.n639 B.n19 585
R114 B.n531 B.n530 585
R115 B.n530 B.n15 585
R116 B.n529 B.n14 585
R117 B.n645 B.n14 585
R118 B.n528 B.n13 585
R119 B.n646 B.n13 585
R120 B.n527 B.n12 585
R121 B.n647 B.n12 585
R122 B.n526 B.n525 585
R123 B.n525 B.n8 585
R124 B.n524 B.n7 585
R125 B.n653 B.n7 585
R126 B.n523 B.n6 585
R127 B.n654 B.n6 585
R128 B.n522 B.n5 585
R129 B.n655 B.n5 585
R130 B.n521 B.n520 585
R131 B.n520 B.n4 585
R132 B.n519 B.n199 585
R133 B.n519 B.n518 585
R134 B.n509 B.n200 585
R135 B.n201 B.n200 585
R136 B.n511 B.n510 585
R137 B.n512 B.n511 585
R138 B.n508 B.n205 585
R139 B.n209 B.n205 585
R140 B.n507 B.n506 585
R141 B.n506 B.n505 585
R142 B.n207 B.n206 585
R143 B.n208 B.n207 585
R144 B.n498 B.n497 585
R145 B.n499 B.n498 585
R146 B.n496 B.n214 585
R147 B.n214 B.n213 585
R148 B.n495 B.n494 585
R149 B.n494 B.n493 585
R150 B.n216 B.n215 585
R151 B.n217 B.n216 585
R152 B.n486 B.n485 585
R153 B.n487 B.n486 585
R154 B.n484 B.n222 585
R155 B.n222 B.n221 585
R156 B.n483 B.n482 585
R157 B.n482 B.n481 585
R158 B.n224 B.n223 585
R159 B.n474 B.n224 585
R160 B.n473 B.n472 585
R161 B.n475 B.n473 585
R162 B.n471 B.n229 585
R163 B.n229 B.n228 585
R164 B.n470 B.n469 585
R165 B.n469 B.n468 585
R166 B.n231 B.n230 585
R167 B.n232 B.n231 585
R168 B.n461 B.n460 585
R169 B.n462 B.n461 585
R170 B.n459 B.n237 585
R171 B.n237 B.n236 585
R172 B.n458 B.n457 585
R173 B.n457 B.n456 585
R174 B.n239 B.n238 585
R175 B.n240 B.n239 585
R176 B.n449 B.n448 585
R177 B.n450 B.n449 585
R178 B.n447 B.n244 585
R179 B.n248 B.n244 585
R180 B.n446 B.n445 585
R181 B.n445 B.n444 585
R182 B.n246 B.n245 585
R183 B.n247 B.n246 585
R184 B.n437 B.n436 585
R185 B.n438 B.n437 585
R186 B.n435 B.n253 585
R187 B.n253 B.n252 585
R188 B.n434 B.n433 585
R189 B.n433 B.n432 585
R190 B.n255 B.n254 585
R191 B.n256 B.n255 585
R192 B.n425 B.n424 585
R193 B.n426 B.n425 585
R194 B.n423 B.n261 585
R195 B.n261 B.n260 585
R196 B.n422 B.n421 585
R197 B.n421 B.n420 585
R198 B.n263 B.n262 585
R199 B.n264 B.n263 585
R200 B.n413 B.n412 585
R201 B.n414 B.n413 585
R202 B.n411 B.n269 585
R203 B.n269 B.n268 585
R204 B.n410 B.n409 585
R205 B.n409 B.n408 585
R206 B.n271 B.n270 585
R207 B.n272 B.n271 585
R208 B.n404 B.n403 585
R209 B.n275 B.n274 585
R210 B.n400 B.n399 585
R211 B.n401 B.n400 585
R212 B.n398 B.n300 585
R213 B.n397 B.n396 585
R214 B.n395 B.n394 585
R215 B.n393 B.n392 585
R216 B.n391 B.n390 585
R217 B.n389 B.n388 585
R218 B.n387 B.n386 585
R219 B.n385 B.n384 585
R220 B.n383 B.n382 585
R221 B.n381 B.n380 585
R222 B.n379 B.n378 585
R223 B.n377 B.n376 585
R224 B.n375 B.n374 585
R225 B.n373 B.n372 585
R226 B.n371 B.n370 585
R227 B.n369 B.n368 585
R228 B.n367 B.n366 585
R229 B.n364 B.n363 585
R230 B.n362 B.n361 585
R231 B.n360 B.n359 585
R232 B.n358 B.n357 585
R233 B.n356 B.n355 585
R234 B.n354 B.n353 585
R235 B.n352 B.n351 585
R236 B.n350 B.n349 585
R237 B.n348 B.n347 585
R238 B.n346 B.n345 585
R239 B.n343 B.n342 585
R240 B.n341 B.n340 585
R241 B.n339 B.n338 585
R242 B.n337 B.n336 585
R243 B.n335 B.n334 585
R244 B.n333 B.n332 585
R245 B.n331 B.n330 585
R246 B.n329 B.n328 585
R247 B.n327 B.n326 585
R248 B.n325 B.n324 585
R249 B.n323 B.n322 585
R250 B.n321 B.n320 585
R251 B.n319 B.n318 585
R252 B.n317 B.n316 585
R253 B.n315 B.n314 585
R254 B.n313 B.n312 585
R255 B.n311 B.n310 585
R256 B.n309 B.n308 585
R257 B.n307 B.n306 585
R258 B.n305 B.n299 585
R259 B.n401 B.n299 585
R260 B.n405 B.n273 585
R261 B.n273 B.n272 585
R262 B.n407 B.n406 585
R263 B.n408 B.n407 585
R264 B.n267 B.n266 585
R265 B.n268 B.n267 585
R266 B.n416 B.n415 585
R267 B.n415 B.n414 585
R268 B.n417 B.n265 585
R269 B.n265 B.n264 585
R270 B.n419 B.n418 585
R271 B.n420 B.n419 585
R272 B.n259 B.n258 585
R273 B.n260 B.n259 585
R274 B.n428 B.n427 585
R275 B.n427 B.n426 585
R276 B.n429 B.n257 585
R277 B.n257 B.n256 585
R278 B.n431 B.n430 585
R279 B.n432 B.n431 585
R280 B.n251 B.n250 585
R281 B.n252 B.n251 585
R282 B.n440 B.n439 585
R283 B.n439 B.n438 585
R284 B.n441 B.n249 585
R285 B.n249 B.n247 585
R286 B.n443 B.n442 585
R287 B.n444 B.n443 585
R288 B.n243 B.n242 585
R289 B.n248 B.n243 585
R290 B.n452 B.n451 585
R291 B.n451 B.n450 585
R292 B.n453 B.n241 585
R293 B.n241 B.n240 585
R294 B.n455 B.n454 585
R295 B.n456 B.n455 585
R296 B.n235 B.n234 585
R297 B.n236 B.n235 585
R298 B.n464 B.n463 585
R299 B.n463 B.n462 585
R300 B.n465 B.n233 585
R301 B.n233 B.n232 585
R302 B.n467 B.n466 585
R303 B.n468 B.n467 585
R304 B.n227 B.n226 585
R305 B.n228 B.n227 585
R306 B.n477 B.n476 585
R307 B.n476 B.n475 585
R308 B.n478 B.n225 585
R309 B.n474 B.n225 585
R310 B.n480 B.n479 585
R311 B.n481 B.n480 585
R312 B.n220 B.n219 585
R313 B.n221 B.n220 585
R314 B.n489 B.n488 585
R315 B.n488 B.n487 585
R316 B.n490 B.n218 585
R317 B.n218 B.n217 585
R318 B.n492 B.n491 585
R319 B.n493 B.n492 585
R320 B.n212 B.n211 585
R321 B.n213 B.n212 585
R322 B.n501 B.n500 585
R323 B.n500 B.n499 585
R324 B.n502 B.n210 585
R325 B.n210 B.n208 585
R326 B.n504 B.n503 585
R327 B.n505 B.n504 585
R328 B.n204 B.n203 585
R329 B.n209 B.n204 585
R330 B.n514 B.n513 585
R331 B.n513 B.n512 585
R332 B.n515 B.n202 585
R333 B.n202 B.n201 585
R334 B.n517 B.n516 585
R335 B.n518 B.n517 585
R336 B.n2 B.n0 585
R337 B.n4 B.n2 585
R338 B.n3 B.n1 585
R339 B.n654 B.n3 585
R340 B.n652 B.n651 585
R341 B.n653 B.n652 585
R342 B.n650 B.n9 585
R343 B.n9 B.n8 585
R344 B.n649 B.n648 585
R345 B.n648 B.n647 585
R346 B.n11 B.n10 585
R347 B.n646 B.n11 585
R348 B.n644 B.n643 585
R349 B.n645 B.n644 585
R350 B.n642 B.n16 585
R351 B.n16 B.n15 585
R352 B.n641 B.n640 585
R353 B.n640 B.n639 585
R354 B.n18 B.n17 585
R355 B.n638 B.n18 585
R356 B.n636 B.n635 585
R357 B.n637 B.n636 585
R358 B.n634 B.n23 585
R359 B.n23 B.n22 585
R360 B.n633 B.n632 585
R361 B.n632 B.n631 585
R362 B.n25 B.n24 585
R363 B.n630 B.n25 585
R364 B.n628 B.n627 585
R365 B.n629 B.n628 585
R366 B.n626 B.n29 585
R367 B.n32 B.n29 585
R368 B.n625 B.n624 585
R369 B.n624 B.n623 585
R370 B.n31 B.n30 585
R371 B.n622 B.n31 585
R372 B.n620 B.n619 585
R373 B.n621 B.n620 585
R374 B.n618 B.n37 585
R375 B.n37 B.n36 585
R376 B.n617 B.n616 585
R377 B.n616 B.n615 585
R378 B.n39 B.n38 585
R379 B.n614 B.n39 585
R380 B.n612 B.n611 585
R381 B.n613 B.n612 585
R382 B.n610 B.n44 585
R383 B.n44 B.n43 585
R384 B.n609 B.n608 585
R385 B.n608 B.n607 585
R386 B.n46 B.n45 585
R387 B.n606 B.n46 585
R388 B.n604 B.n603 585
R389 B.n605 B.n604 585
R390 B.n602 B.n51 585
R391 B.n51 B.n50 585
R392 B.n601 B.n600 585
R393 B.n600 B.n599 585
R394 B.n53 B.n52 585
R395 B.n598 B.n53 585
R396 B.n596 B.n595 585
R397 B.n597 B.n596 585
R398 B.n594 B.n58 585
R399 B.n58 B.n57 585
R400 B.n593 B.n592 585
R401 B.n592 B.n591 585
R402 B.n60 B.n59 585
R403 B.n590 B.n60 585
R404 B.n588 B.n587 585
R405 B.n589 B.n588 585
R406 B.n586 B.n65 585
R407 B.n65 B.n64 585
R408 B.n585 B.n584 585
R409 B.n584 B.n583 585
R410 B.n67 B.n66 585
R411 B.n582 B.n67 585
R412 B.n580 B.n579 585
R413 B.n581 B.n580 585
R414 B.n578 B.n72 585
R415 B.n72 B.n71 585
R416 B.n657 B.n656 585
R417 B.n656 B.n655 585
R418 B.n403 B.n273 492.5
R419 B.n576 B.n72 492.5
R420 B.n299 B.n271 492.5
R421 B.n572 B.n99 492.5
R422 B.n303 B.t13 283.536
R423 B.n301 B.t9 283.536
R424 B.n103 B.t20 283.536
R425 B.n100 B.t16 283.536
R426 B.n574 B.n573 256.663
R427 B.n574 B.n97 256.663
R428 B.n574 B.n96 256.663
R429 B.n574 B.n95 256.663
R430 B.n574 B.n94 256.663
R431 B.n574 B.n93 256.663
R432 B.n574 B.n92 256.663
R433 B.n574 B.n91 256.663
R434 B.n574 B.n90 256.663
R435 B.n574 B.n89 256.663
R436 B.n574 B.n88 256.663
R437 B.n574 B.n87 256.663
R438 B.n574 B.n86 256.663
R439 B.n574 B.n85 256.663
R440 B.n574 B.n84 256.663
R441 B.n574 B.n83 256.663
R442 B.n574 B.n82 256.663
R443 B.n574 B.n81 256.663
R444 B.n574 B.n80 256.663
R445 B.n574 B.n79 256.663
R446 B.n574 B.n78 256.663
R447 B.n574 B.n77 256.663
R448 B.n574 B.n76 256.663
R449 B.n574 B.n75 256.663
R450 B.n575 B.n574 256.663
R451 B.n402 B.n401 256.663
R452 B.n401 B.n276 256.663
R453 B.n401 B.n277 256.663
R454 B.n401 B.n278 256.663
R455 B.n401 B.n279 256.663
R456 B.n401 B.n280 256.663
R457 B.n401 B.n281 256.663
R458 B.n401 B.n282 256.663
R459 B.n401 B.n283 256.663
R460 B.n401 B.n284 256.663
R461 B.n401 B.n285 256.663
R462 B.n401 B.n286 256.663
R463 B.n401 B.n287 256.663
R464 B.n401 B.n288 256.663
R465 B.n401 B.n289 256.663
R466 B.n401 B.n290 256.663
R467 B.n401 B.n291 256.663
R468 B.n401 B.n292 256.663
R469 B.n401 B.n293 256.663
R470 B.n401 B.n294 256.663
R471 B.n401 B.n295 256.663
R472 B.n401 B.n296 256.663
R473 B.n401 B.n297 256.663
R474 B.n401 B.n298 256.663
R475 B.n303 B.t15 190.133
R476 B.n100 B.t18 190.133
R477 B.n301 B.t12 190.133
R478 B.n103 B.t21 190.133
R479 B.n407 B.n273 163.367
R480 B.n407 B.n267 163.367
R481 B.n415 B.n267 163.367
R482 B.n415 B.n265 163.367
R483 B.n419 B.n265 163.367
R484 B.n419 B.n259 163.367
R485 B.n427 B.n259 163.367
R486 B.n427 B.n257 163.367
R487 B.n431 B.n257 163.367
R488 B.n431 B.n251 163.367
R489 B.n439 B.n251 163.367
R490 B.n439 B.n249 163.367
R491 B.n443 B.n249 163.367
R492 B.n443 B.n243 163.367
R493 B.n451 B.n243 163.367
R494 B.n451 B.n241 163.367
R495 B.n455 B.n241 163.367
R496 B.n455 B.n235 163.367
R497 B.n463 B.n235 163.367
R498 B.n463 B.n233 163.367
R499 B.n467 B.n233 163.367
R500 B.n467 B.n227 163.367
R501 B.n476 B.n227 163.367
R502 B.n476 B.n225 163.367
R503 B.n480 B.n225 163.367
R504 B.n480 B.n220 163.367
R505 B.n488 B.n220 163.367
R506 B.n488 B.n218 163.367
R507 B.n492 B.n218 163.367
R508 B.n492 B.n212 163.367
R509 B.n500 B.n212 163.367
R510 B.n500 B.n210 163.367
R511 B.n504 B.n210 163.367
R512 B.n504 B.n204 163.367
R513 B.n513 B.n204 163.367
R514 B.n513 B.n202 163.367
R515 B.n517 B.n202 163.367
R516 B.n517 B.n2 163.367
R517 B.n656 B.n2 163.367
R518 B.n656 B.n3 163.367
R519 B.n652 B.n3 163.367
R520 B.n652 B.n9 163.367
R521 B.n648 B.n9 163.367
R522 B.n648 B.n11 163.367
R523 B.n644 B.n11 163.367
R524 B.n644 B.n16 163.367
R525 B.n640 B.n16 163.367
R526 B.n640 B.n18 163.367
R527 B.n636 B.n18 163.367
R528 B.n636 B.n23 163.367
R529 B.n632 B.n23 163.367
R530 B.n632 B.n25 163.367
R531 B.n628 B.n25 163.367
R532 B.n628 B.n29 163.367
R533 B.n624 B.n29 163.367
R534 B.n624 B.n31 163.367
R535 B.n620 B.n31 163.367
R536 B.n620 B.n37 163.367
R537 B.n616 B.n37 163.367
R538 B.n616 B.n39 163.367
R539 B.n612 B.n39 163.367
R540 B.n612 B.n44 163.367
R541 B.n608 B.n44 163.367
R542 B.n608 B.n46 163.367
R543 B.n604 B.n46 163.367
R544 B.n604 B.n51 163.367
R545 B.n600 B.n51 163.367
R546 B.n600 B.n53 163.367
R547 B.n596 B.n53 163.367
R548 B.n596 B.n58 163.367
R549 B.n592 B.n58 163.367
R550 B.n592 B.n60 163.367
R551 B.n588 B.n60 163.367
R552 B.n588 B.n65 163.367
R553 B.n584 B.n65 163.367
R554 B.n584 B.n67 163.367
R555 B.n580 B.n67 163.367
R556 B.n580 B.n72 163.367
R557 B.n400 B.n275 163.367
R558 B.n400 B.n300 163.367
R559 B.n396 B.n395 163.367
R560 B.n392 B.n391 163.367
R561 B.n388 B.n387 163.367
R562 B.n384 B.n383 163.367
R563 B.n380 B.n379 163.367
R564 B.n376 B.n375 163.367
R565 B.n372 B.n371 163.367
R566 B.n368 B.n367 163.367
R567 B.n363 B.n362 163.367
R568 B.n359 B.n358 163.367
R569 B.n355 B.n354 163.367
R570 B.n351 B.n350 163.367
R571 B.n347 B.n346 163.367
R572 B.n342 B.n341 163.367
R573 B.n338 B.n337 163.367
R574 B.n334 B.n333 163.367
R575 B.n330 B.n329 163.367
R576 B.n326 B.n325 163.367
R577 B.n322 B.n321 163.367
R578 B.n318 B.n317 163.367
R579 B.n314 B.n313 163.367
R580 B.n310 B.n309 163.367
R581 B.n306 B.n299 163.367
R582 B.n409 B.n271 163.367
R583 B.n409 B.n269 163.367
R584 B.n413 B.n269 163.367
R585 B.n413 B.n263 163.367
R586 B.n421 B.n263 163.367
R587 B.n421 B.n261 163.367
R588 B.n425 B.n261 163.367
R589 B.n425 B.n255 163.367
R590 B.n433 B.n255 163.367
R591 B.n433 B.n253 163.367
R592 B.n437 B.n253 163.367
R593 B.n437 B.n246 163.367
R594 B.n445 B.n246 163.367
R595 B.n445 B.n244 163.367
R596 B.n449 B.n244 163.367
R597 B.n449 B.n239 163.367
R598 B.n457 B.n239 163.367
R599 B.n457 B.n237 163.367
R600 B.n461 B.n237 163.367
R601 B.n461 B.n231 163.367
R602 B.n469 B.n231 163.367
R603 B.n469 B.n229 163.367
R604 B.n473 B.n229 163.367
R605 B.n473 B.n224 163.367
R606 B.n482 B.n224 163.367
R607 B.n482 B.n222 163.367
R608 B.n486 B.n222 163.367
R609 B.n486 B.n216 163.367
R610 B.n494 B.n216 163.367
R611 B.n494 B.n214 163.367
R612 B.n498 B.n214 163.367
R613 B.n498 B.n207 163.367
R614 B.n506 B.n207 163.367
R615 B.n506 B.n205 163.367
R616 B.n511 B.n205 163.367
R617 B.n511 B.n200 163.367
R618 B.n519 B.n200 163.367
R619 B.n520 B.n519 163.367
R620 B.n520 B.n5 163.367
R621 B.n6 B.n5 163.367
R622 B.n7 B.n6 163.367
R623 B.n525 B.n7 163.367
R624 B.n525 B.n12 163.367
R625 B.n13 B.n12 163.367
R626 B.n14 B.n13 163.367
R627 B.n530 B.n14 163.367
R628 B.n530 B.n19 163.367
R629 B.n20 B.n19 163.367
R630 B.n21 B.n20 163.367
R631 B.n535 B.n21 163.367
R632 B.n535 B.n26 163.367
R633 B.n27 B.n26 163.367
R634 B.n28 B.n27 163.367
R635 B.n540 B.n28 163.367
R636 B.n540 B.n33 163.367
R637 B.n34 B.n33 163.367
R638 B.n35 B.n34 163.367
R639 B.n545 B.n35 163.367
R640 B.n545 B.n40 163.367
R641 B.n41 B.n40 163.367
R642 B.n42 B.n41 163.367
R643 B.n550 B.n42 163.367
R644 B.n550 B.n47 163.367
R645 B.n48 B.n47 163.367
R646 B.n49 B.n48 163.367
R647 B.n555 B.n49 163.367
R648 B.n555 B.n54 163.367
R649 B.n55 B.n54 163.367
R650 B.n56 B.n55 163.367
R651 B.n560 B.n56 163.367
R652 B.n560 B.n61 163.367
R653 B.n62 B.n61 163.367
R654 B.n63 B.n62 163.367
R655 B.n565 B.n63 163.367
R656 B.n565 B.n68 163.367
R657 B.n69 B.n68 163.367
R658 B.n70 B.n69 163.367
R659 B.n99 B.n70 163.367
R660 B.n106 B.n74 163.367
R661 B.n110 B.n109 163.367
R662 B.n114 B.n113 163.367
R663 B.n118 B.n117 163.367
R664 B.n122 B.n121 163.367
R665 B.n126 B.n125 163.367
R666 B.n130 B.n129 163.367
R667 B.n134 B.n133 163.367
R668 B.n138 B.n137 163.367
R669 B.n142 B.n141 163.367
R670 B.n146 B.n145 163.367
R671 B.n150 B.n149 163.367
R672 B.n154 B.n153 163.367
R673 B.n158 B.n157 163.367
R674 B.n162 B.n161 163.367
R675 B.n166 B.n165 163.367
R676 B.n170 B.n169 163.367
R677 B.n174 B.n173 163.367
R678 B.n178 B.n177 163.367
R679 B.n182 B.n181 163.367
R680 B.n186 B.n185 163.367
R681 B.n190 B.n189 163.367
R682 B.n194 B.n193 163.367
R683 B.n196 B.n98 163.367
R684 B.n304 B.t14 156
R685 B.n101 B.t19 156
R686 B.n302 B.t11 156
R687 B.n104 B.t22 156
R688 B.n401 B.n272 149.623
R689 B.n574 B.n71 149.623
R690 B.n408 B.n272 75.3657
R691 B.n408 B.n268 75.3657
R692 B.n414 B.n268 75.3657
R693 B.n414 B.n264 75.3657
R694 B.n420 B.n264 75.3657
R695 B.n426 B.n260 75.3657
R696 B.n426 B.n256 75.3657
R697 B.n432 B.n256 75.3657
R698 B.n432 B.n252 75.3657
R699 B.n438 B.n252 75.3657
R700 B.n438 B.n247 75.3657
R701 B.n444 B.n247 75.3657
R702 B.n444 B.n248 75.3657
R703 B.n450 B.n240 75.3657
R704 B.n456 B.n240 75.3657
R705 B.n456 B.n236 75.3657
R706 B.n462 B.n236 75.3657
R707 B.n468 B.n232 75.3657
R708 B.n468 B.n228 75.3657
R709 B.n475 B.n228 75.3657
R710 B.n475 B.n474 75.3657
R711 B.n481 B.n221 75.3657
R712 B.n487 B.n221 75.3657
R713 B.n487 B.n217 75.3657
R714 B.n493 B.n217 75.3657
R715 B.n499 B.n213 75.3657
R716 B.n499 B.n208 75.3657
R717 B.n505 B.n208 75.3657
R718 B.n505 B.n209 75.3657
R719 B.n512 B.n201 75.3657
R720 B.n518 B.n201 75.3657
R721 B.n518 B.n4 75.3657
R722 B.n655 B.n4 75.3657
R723 B.n655 B.n654 75.3657
R724 B.n654 B.n653 75.3657
R725 B.n653 B.n8 75.3657
R726 B.n647 B.n8 75.3657
R727 B.n646 B.n645 75.3657
R728 B.n645 B.n15 75.3657
R729 B.n639 B.n15 75.3657
R730 B.n639 B.n638 75.3657
R731 B.n637 B.n22 75.3657
R732 B.n631 B.n22 75.3657
R733 B.n631 B.n630 75.3657
R734 B.n630 B.n629 75.3657
R735 B.n623 B.n32 75.3657
R736 B.n623 B.n622 75.3657
R737 B.n622 B.n621 75.3657
R738 B.n621 B.n36 75.3657
R739 B.n615 B.n614 75.3657
R740 B.n614 B.n613 75.3657
R741 B.n613 B.n43 75.3657
R742 B.n607 B.n43 75.3657
R743 B.n606 B.n605 75.3657
R744 B.n605 B.n50 75.3657
R745 B.n599 B.n50 75.3657
R746 B.n599 B.n598 75.3657
R747 B.n598 B.n597 75.3657
R748 B.n597 B.n57 75.3657
R749 B.n591 B.n57 75.3657
R750 B.n591 B.n590 75.3657
R751 B.n589 B.n64 75.3657
R752 B.n583 B.n64 75.3657
R753 B.n583 B.n582 75.3657
R754 B.n582 B.n581 75.3657
R755 B.n581 B.n71 75.3657
R756 B.n403 B.n402 71.676
R757 B.n300 B.n276 71.676
R758 B.n395 B.n277 71.676
R759 B.n391 B.n278 71.676
R760 B.n387 B.n279 71.676
R761 B.n383 B.n280 71.676
R762 B.n379 B.n281 71.676
R763 B.n375 B.n282 71.676
R764 B.n371 B.n283 71.676
R765 B.n367 B.n284 71.676
R766 B.n362 B.n285 71.676
R767 B.n358 B.n286 71.676
R768 B.n354 B.n287 71.676
R769 B.n350 B.n288 71.676
R770 B.n346 B.n289 71.676
R771 B.n341 B.n290 71.676
R772 B.n337 B.n291 71.676
R773 B.n333 B.n292 71.676
R774 B.n329 B.n293 71.676
R775 B.n325 B.n294 71.676
R776 B.n321 B.n295 71.676
R777 B.n317 B.n296 71.676
R778 B.n313 B.n297 71.676
R779 B.n309 B.n298 71.676
R780 B.n576 B.n575 71.676
R781 B.n106 B.n75 71.676
R782 B.n110 B.n76 71.676
R783 B.n114 B.n77 71.676
R784 B.n118 B.n78 71.676
R785 B.n122 B.n79 71.676
R786 B.n126 B.n80 71.676
R787 B.n130 B.n81 71.676
R788 B.n134 B.n82 71.676
R789 B.n138 B.n83 71.676
R790 B.n142 B.n84 71.676
R791 B.n146 B.n85 71.676
R792 B.n150 B.n86 71.676
R793 B.n154 B.n87 71.676
R794 B.n158 B.n88 71.676
R795 B.n162 B.n89 71.676
R796 B.n166 B.n90 71.676
R797 B.n170 B.n91 71.676
R798 B.n174 B.n92 71.676
R799 B.n178 B.n93 71.676
R800 B.n182 B.n94 71.676
R801 B.n186 B.n95 71.676
R802 B.n190 B.n96 71.676
R803 B.n194 B.n97 71.676
R804 B.n573 B.n98 71.676
R805 B.n573 B.n572 71.676
R806 B.n196 B.n97 71.676
R807 B.n193 B.n96 71.676
R808 B.n189 B.n95 71.676
R809 B.n185 B.n94 71.676
R810 B.n181 B.n93 71.676
R811 B.n177 B.n92 71.676
R812 B.n173 B.n91 71.676
R813 B.n169 B.n90 71.676
R814 B.n165 B.n89 71.676
R815 B.n161 B.n88 71.676
R816 B.n157 B.n87 71.676
R817 B.n153 B.n86 71.676
R818 B.n149 B.n85 71.676
R819 B.n145 B.n84 71.676
R820 B.n141 B.n83 71.676
R821 B.n137 B.n82 71.676
R822 B.n133 B.n81 71.676
R823 B.n129 B.n80 71.676
R824 B.n125 B.n79 71.676
R825 B.n121 B.n78 71.676
R826 B.n117 B.n77 71.676
R827 B.n113 B.n76 71.676
R828 B.n109 B.n75 71.676
R829 B.n575 B.n74 71.676
R830 B.n402 B.n275 71.676
R831 B.n396 B.n276 71.676
R832 B.n392 B.n277 71.676
R833 B.n388 B.n278 71.676
R834 B.n384 B.n279 71.676
R835 B.n380 B.n280 71.676
R836 B.n376 B.n281 71.676
R837 B.n372 B.n282 71.676
R838 B.n368 B.n283 71.676
R839 B.n363 B.n284 71.676
R840 B.n359 B.n285 71.676
R841 B.n355 B.n286 71.676
R842 B.n351 B.n287 71.676
R843 B.n347 B.n288 71.676
R844 B.n342 B.n289 71.676
R845 B.n338 B.n290 71.676
R846 B.n334 B.n291 71.676
R847 B.n330 B.n292 71.676
R848 B.n326 B.n293 71.676
R849 B.n322 B.n294 71.676
R850 B.n318 B.n295 71.676
R851 B.n314 B.n296 71.676
R852 B.n310 B.n297 71.676
R853 B.n306 B.n298 71.676
R854 B.n450 B.t3 67.6076
R855 B.n607 B.t2 67.6076
R856 B.n209 B.t6 60.9577
R857 B.t1 B.n646 60.9577
R858 B.n344 B.n304 59.5399
R859 B.n365 B.n302 59.5399
R860 B.n105 B.n104 59.5399
R861 B.n102 B.n101 59.5399
R862 B.n420 B.t10 54.3078
R863 B.t7 B.n232 54.3078
R864 B.t5 B.n36 54.3078
R865 B.t17 B.n589 54.3078
R866 B.n493 B.t0 47.6579
R867 B.t8 B.n637 47.6579
R868 B.n481 B.t23 41.0081
R869 B.n629 B.t4 41.0081
R870 B.n474 B.t23 34.3582
R871 B.n32 B.t4 34.3582
R872 B.n304 B.n303 34.1338
R873 B.n302 B.n301 34.1338
R874 B.n104 B.n103 34.1338
R875 B.n101 B.n100 34.1338
R876 B.n578 B.n577 32.0005
R877 B.n571 B.n570 32.0005
R878 B.n305 B.n270 32.0005
R879 B.n405 B.n404 32.0005
R880 B.t0 B.n213 27.7083
R881 B.n638 B.t8 27.7083
R882 B.t10 B.n260 21.0584
R883 B.n462 B.t7 21.0584
R884 B.n615 B.t5 21.0584
R885 B.n590 B.t17 21.0584
R886 B B.n657 18.0485
R887 B.n512 B.t6 14.4086
R888 B.n647 B.t1 14.4086
R889 B.n577 B.n73 10.6151
R890 B.n107 B.n73 10.6151
R891 B.n108 B.n107 10.6151
R892 B.n111 B.n108 10.6151
R893 B.n112 B.n111 10.6151
R894 B.n115 B.n112 10.6151
R895 B.n116 B.n115 10.6151
R896 B.n119 B.n116 10.6151
R897 B.n120 B.n119 10.6151
R898 B.n123 B.n120 10.6151
R899 B.n124 B.n123 10.6151
R900 B.n127 B.n124 10.6151
R901 B.n128 B.n127 10.6151
R902 B.n131 B.n128 10.6151
R903 B.n132 B.n131 10.6151
R904 B.n135 B.n132 10.6151
R905 B.n136 B.n135 10.6151
R906 B.n139 B.n136 10.6151
R907 B.n140 B.n139 10.6151
R908 B.n144 B.n143 10.6151
R909 B.n147 B.n144 10.6151
R910 B.n148 B.n147 10.6151
R911 B.n151 B.n148 10.6151
R912 B.n152 B.n151 10.6151
R913 B.n155 B.n152 10.6151
R914 B.n156 B.n155 10.6151
R915 B.n159 B.n156 10.6151
R916 B.n160 B.n159 10.6151
R917 B.n164 B.n163 10.6151
R918 B.n167 B.n164 10.6151
R919 B.n168 B.n167 10.6151
R920 B.n171 B.n168 10.6151
R921 B.n172 B.n171 10.6151
R922 B.n175 B.n172 10.6151
R923 B.n176 B.n175 10.6151
R924 B.n179 B.n176 10.6151
R925 B.n180 B.n179 10.6151
R926 B.n183 B.n180 10.6151
R927 B.n184 B.n183 10.6151
R928 B.n187 B.n184 10.6151
R929 B.n188 B.n187 10.6151
R930 B.n191 B.n188 10.6151
R931 B.n192 B.n191 10.6151
R932 B.n195 B.n192 10.6151
R933 B.n197 B.n195 10.6151
R934 B.n198 B.n197 10.6151
R935 B.n571 B.n198 10.6151
R936 B.n410 B.n270 10.6151
R937 B.n411 B.n410 10.6151
R938 B.n412 B.n411 10.6151
R939 B.n412 B.n262 10.6151
R940 B.n422 B.n262 10.6151
R941 B.n423 B.n422 10.6151
R942 B.n424 B.n423 10.6151
R943 B.n424 B.n254 10.6151
R944 B.n434 B.n254 10.6151
R945 B.n435 B.n434 10.6151
R946 B.n436 B.n435 10.6151
R947 B.n436 B.n245 10.6151
R948 B.n446 B.n245 10.6151
R949 B.n447 B.n446 10.6151
R950 B.n448 B.n447 10.6151
R951 B.n448 B.n238 10.6151
R952 B.n458 B.n238 10.6151
R953 B.n459 B.n458 10.6151
R954 B.n460 B.n459 10.6151
R955 B.n460 B.n230 10.6151
R956 B.n470 B.n230 10.6151
R957 B.n471 B.n470 10.6151
R958 B.n472 B.n471 10.6151
R959 B.n472 B.n223 10.6151
R960 B.n483 B.n223 10.6151
R961 B.n484 B.n483 10.6151
R962 B.n485 B.n484 10.6151
R963 B.n485 B.n215 10.6151
R964 B.n495 B.n215 10.6151
R965 B.n496 B.n495 10.6151
R966 B.n497 B.n496 10.6151
R967 B.n497 B.n206 10.6151
R968 B.n507 B.n206 10.6151
R969 B.n508 B.n507 10.6151
R970 B.n510 B.n508 10.6151
R971 B.n510 B.n509 10.6151
R972 B.n509 B.n199 10.6151
R973 B.n521 B.n199 10.6151
R974 B.n522 B.n521 10.6151
R975 B.n523 B.n522 10.6151
R976 B.n524 B.n523 10.6151
R977 B.n526 B.n524 10.6151
R978 B.n527 B.n526 10.6151
R979 B.n528 B.n527 10.6151
R980 B.n529 B.n528 10.6151
R981 B.n531 B.n529 10.6151
R982 B.n532 B.n531 10.6151
R983 B.n533 B.n532 10.6151
R984 B.n534 B.n533 10.6151
R985 B.n536 B.n534 10.6151
R986 B.n537 B.n536 10.6151
R987 B.n538 B.n537 10.6151
R988 B.n539 B.n538 10.6151
R989 B.n541 B.n539 10.6151
R990 B.n542 B.n541 10.6151
R991 B.n543 B.n542 10.6151
R992 B.n544 B.n543 10.6151
R993 B.n546 B.n544 10.6151
R994 B.n547 B.n546 10.6151
R995 B.n548 B.n547 10.6151
R996 B.n549 B.n548 10.6151
R997 B.n551 B.n549 10.6151
R998 B.n552 B.n551 10.6151
R999 B.n553 B.n552 10.6151
R1000 B.n554 B.n553 10.6151
R1001 B.n556 B.n554 10.6151
R1002 B.n557 B.n556 10.6151
R1003 B.n558 B.n557 10.6151
R1004 B.n559 B.n558 10.6151
R1005 B.n561 B.n559 10.6151
R1006 B.n562 B.n561 10.6151
R1007 B.n563 B.n562 10.6151
R1008 B.n564 B.n563 10.6151
R1009 B.n566 B.n564 10.6151
R1010 B.n567 B.n566 10.6151
R1011 B.n568 B.n567 10.6151
R1012 B.n569 B.n568 10.6151
R1013 B.n570 B.n569 10.6151
R1014 B.n404 B.n274 10.6151
R1015 B.n399 B.n274 10.6151
R1016 B.n399 B.n398 10.6151
R1017 B.n398 B.n397 10.6151
R1018 B.n397 B.n394 10.6151
R1019 B.n394 B.n393 10.6151
R1020 B.n393 B.n390 10.6151
R1021 B.n390 B.n389 10.6151
R1022 B.n389 B.n386 10.6151
R1023 B.n386 B.n385 10.6151
R1024 B.n385 B.n382 10.6151
R1025 B.n382 B.n381 10.6151
R1026 B.n381 B.n378 10.6151
R1027 B.n378 B.n377 10.6151
R1028 B.n377 B.n374 10.6151
R1029 B.n374 B.n373 10.6151
R1030 B.n373 B.n370 10.6151
R1031 B.n370 B.n369 10.6151
R1032 B.n369 B.n366 10.6151
R1033 B.n364 B.n361 10.6151
R1034 B.n361 B.n360 10.6151
R1035 B.n360 B.n357 10.6151
R1036 B.n357 B.n356 10.6151
R1037 B.n356 B.n353 10.6151
R1038 B.n353 B.n352 10.6151
R1039 B.n352 B.n349 10.6151
R1040 B.n349 B.n348 10.6151
R1041 B.n348 B.n345 10.6151
R1042 B.n343 B.n340 10.6151
R1043 B.n340 B.n339 10.6151
R1044 B.n339 B.n336 10.6151
R1045 B.n336 B.n335 10.6151
R1046 B.n335 B.n332 10.6151
R1047 B.n332 B.n331 10.6151
R1048 B.n331 B.n328 10.6151
R1049 B.n328 B.n327 10.6151
R1050 B.n327 B.n324 10.6151
R1051 B.n324 B.n323 10.6151
R1052 B.n323 B.n320 10.6151
R1053 B.n320 B.n319 10.6151
R1054 B.n319 B.n316 10.6151
R1055 B.n316 B.n315 10.6151
R1056 B.n315 B.n312 10.6151
R1057 B.n312 B.n311 10.6151
R1058 B.n311 B.n308 10.6151
R1059 B.n308 B.n307 10.6151
R1060 B.n307 B.n305 10.6151
R1061 B.n406 B.n405 10.6151
R1062 B.n406 B.n266 10.6151
R1063 B.n416 B.n266 10.6151
R1064 B.n417 B.n416 10.6151
R1065 B.n418 B.n417 10.6151
R1066 B.n418 B.n258 10.6151
R1067 B.n428 B.n258 10.6151
R1068 B.n429 B.n428 10.6151
R1069 B.n430 B.n429 10.6151
R1070 B.n430 B.n250 10.6151
R1071 B.n440 B.n250 10.6151
R1072 B.n441 B.n440 10.6151
R1073 B.n442 B.n441 10.6151
R1074 B.n442 B.n242 10.6151
R1075 B.n452 B.n242 10.6151
R1076 B.n453 B.n452 10.6151
R1077 B.n454 B.n453 10.6151
R1078 B.n454 B.n234 10.6151
R1079 B.n464 B.n234 10.6151
R1080 B.n465 B.n464 10.6151
R1081 B.n466 B.n465 10.6151
R1082 B.n466 B.n226 10.6151
R1083 B.n477 B.n226 10.6151
R1084 B.n478 B.n477 10.6151
R1085 B.n479 B.n478 10.6151
R1086 B.n479 B.n219 10.6151
R1087 B.n489 B.n219 10.6151
R1088 B.n490 B.n489 10.6151
R1089 B.n491 B.n490 10.6151
R1090 B.n491 B.n211 10.6151
R1091 B.n501 B.n211 10.6151
R1092 B.n502 B.n501 10.6151
R1093 B.n503 B.n502 10.6151
R1094 B.n503 B.n203 10.6151
R1095 B.n514 B.n203 10.6151
R1096 B.n515 B.n514 10.6151
R1097 B.n516 B.n515 10.6151
R1098 B.n516 B.n0 10.6151
R1099 B.n651 B.n1 10.6151
R1100 B.n651 B.n650 10.6151
R1101 B.n650 B.n649 10.6151
R1102 B.n649 B.n10 10.6151
R1103 B.n643 B.n10 10.6151
R1104 B.n643 B.n642 10.6151
R1105 B.n642 B.n641 10.6151
R1106 B.n641 B.n17 10.6151
R1107 B.n635 B.n17 10.6151
R1108 B.n635 B.n634 10.6151
R1109 B.n634 B.n633 10.6151
R1110 B.n633 B.n24 10.6151
R1111 B.n627 B.n24 10.6151
R1112 B.n627 B.n626 10.6151
R1113 B.n626 B.n625 10.6151
R1114 B.n625 B.n30 10.6151
R1115 B.n619 B.n30 10.6151
R1116 B.n619 B.n618 10.6151
R1117 B.n618 B.n617 10.6151
R1118 B.n617 B.n38 10.6151
R1119 B.n611 B.n38 10.6151
R1120 B.n611 B.n610 10.6151
R1121 B.n610 B.n609 10.6151
R1122 B.n609 B.n45 10.6151
R1123 B.n603 B.n45 10.6151
R1124 B.n603 B.n602 10.6151
R1125 B.n602 B.n601 10.6151
R1126 B.n601 B.n52 10.6151
R1127 B.n595 B.n52 10.6151
R1128 B.n595 B.n594 10.6151
R1129 B.n594 B.n593 10.6151
R1130 B.n593 B.n59 10.6151
R1131 B.n587 B.n59 10.6151
R1132 B.n587 B.n586 10.6151
R1133 B.n586 B.n585 10.6151
R1134 B.n585 B.n66 10.6151
R1135 B.n579 B.n66 10.6151
R1136 B.n579 B.n578 10.6151
R1137 B.n140 B.n105 9.36635
R1138 B.n163 B.n102 9.36635
R1139 B.n366 B.n365 9.36635
R1140 B.n344 B.n343 9.36635
R1141 B.n248 B.t3 7.75869
R1142 B.t2 B.n606 7.75869
R1143 B.n657 B.n0 2.81026
R1144 B.n657 B.n1 2.81026
R1145 B.n143 B.n105 1.24928
R1146 B.n160 B.n102 1.24928
R1147 B.n365 B.n364 1.24928
R1148 B.n345 B.n344 1.24928
R1149 VN.n27 VN.n26 172.555
R1150 VN.n55 VN.n54 172.555
R1151 VN.n53 VN.n28 161.3
R1152 VN.n52 VN.n51 161.3
R1153 VN.n50 VN.n29 161.3
R1154 VN.n49 VN.n48 161.3
R1155 VN.n47 VN.n30 161.3
R1156 VN.n46 VN.n45 161.3
R1157 VN.n44 VN.n32 161.3
R1158 VN.n43 VN.n42 161.3
R1159 VN.n41 VN.n33 161.3
R1160 VN.n40 VN.n39 161.3
R1161 VN.n38 VN.n35 161.3
R1162 VN.n25 VN.n0 161.3
R1163 VN.n24 VN.n23 161.3
R1164 VN.n22 VN.n1 161.3
R1165 VN.n21 VN.n20 161.3
R1166 VN.n18 VN.n2 161.3
R1167 VN.n17 VN.n16 161.3
R1168 VN.n15 VN.n3 161.3
R1169 VN.n14 VN.n13 161.3
R1170 VN.n11 VN.n4 161.3
R1171 VN.n10 VN.n9 161.3
R1172 VN.n8 VN.n5 161.3
R1173 VN.n7 VN.t9 107.415
R1174 VN.n37 VN.t3 107.415
R1175 VN.n6 VN.t7 78.3676
R1176 VN.n12 VN.t6 78.3676
R1177 VN.n19 VN.t5 78.3676
R1178 VN.n26 VN.t0 78.3676
R1179 VN.n36 VN.t4 78.3676
R1180 VN.n34 VN.t1 78.3676
R1181 VN.n31 VN.t2 78.3676
R1182 VN.n54 VN.t8 78.3676
R1183 VN.n7 VN.n6 65.4496
R1184 VN.n37 VN.n36 65.4496
R1185 VN.n11 VN.n10 53.1199
R1186 VN.n18 VN.n17 53.1199
R1187 VN.n41 VN.n40 53.1199
R1188 VN.n47 VN.n46 53.1199
R1189 VN.n24 VN.n1 51.1773
R1190 VN.n52 VN.n29 51.1773
R1191 VN VN.n55 41.5251
R1192 VN.n25 VN.n24 29.8095
R1193 VN.n53 VN.n52 29.8095
R1194 VN.n13 VN.n11 27.8669
R1195 VN.n17 VN.n3 27.8669
R1196 VN.n42 VN.n41 27.8669
R1197 VN.n46 VN.n32 27.8669
R1198 VN.n38 VN.n37 27.1884
R1199 VN.n8 VN.n7 27.1884
R1200 VN.n10 VN.n5 24.4675
R1201 VN.n20 VN.n18 24.4675
R1202 VN.n40 VN.n35 24.4675
R1203 VN.n48 VN.n47 24.4675
R1204 VN.n19 VN.n1 23.9782
R1205 VN.n31 VN.n29 23.9782
R1206 VN.n26 VN.n25 13.2127
R1207 VN.n54 VN.n53 13.2127
R1208 VN.n13 VN.n12 12.234
R1209 VN.n12 VN.n3 12.234
R1210 VN.n34 VN.n32 12.234
R1211 VN.n42 VN.n34 12.234
R1212 VN.n6 VN.n5 0.48984
R1213 VN.n20 VN.n19 0.48984
R1214 VN.n36 VN.n35 0.48984
R1215 VN.n48 VN.n31 0.48984
R1216 VN.n55 VN.n28 0.189894
R1217 VN.n51 VN.n28 0.189894
R1218 VN.n51 VN.n50 0.189894
R1219 VN.n50 VN.n49 0.189894
R1220 VN.n49 VN.n30 0.189894
R1221 VN.n45 VN.n30 0.189894
R1222 VN.n45 VN.n44 0.189894
R1223 VN.n44 VN.n43 0.189894
R1224 VN.n43 VN.n33 0.189894
R1225 VN.n39 VN.n33 0.189894
R1226 VN.n39 VN.n38 0.189894
R1227 VN.n9 VN.n8 0.189894
R1228 VN.n9 VN.n4 0.189894
R1229 VN.n14 VN.n4 0.189894
R1230 VN.n15 VN.n14 0.189894
R1231 VN.n16 VN.n15 0.189894
R1232 VN.n16 VN.n2 0.189894
R1233 VN.n21 VN.n2 0.189894
R1234 VN.n22 VN.n21 0.189894
R1235 VN.n23 VN.n22 0.189894
R1236 VN.n23 VN.n0 0.189894
R1237 VN.n27 VN.n0 0.189894
R1238 VN VN.n27 0.0516364
R1239 VTAIL.n104 VTAIL.n86 289.615
R1240 VTAIL.n20 VTAIL.n2 289.615
R1241 VTAIL.n80 VTAIL.n62 289.615
R1242 VTAIL.n52 VTAIL.n34 289.615
R1243 VTAIL.n95 VTAIL.n94 185
R1244 VTAIL.n97 VTAIL.n96 185
R1245 VTAIL.n90 VTAIL.n89 185
R1246 VTAIL.n103 VTAIL.n102 185
R1247 VTAIL.n105 VTAIL.n104 185
R1248 VTAIL.n11 VTAIL.n10 185
R1249 VTAIL.n13 VTAIL.n12 185
R1250 VTAIL.n6 VTAIL.n5 185
R1251 VTAIL.n19 VTAIL.n18 185
R1252 VTAIL.n21 VTAIL.n20 185
R1253 VTAIL.n81 VTAIL.n80 185
R1254 VTAIL.n79 VTAIL.n78 185
R1255 VTAIL.n66 VTAIL.n65 185
R1256 VTAIL.n73 VTAIL.n72 185
R1257 VTAIL.n71 VTAIL.n70 185
R1258 VTAIL.n53 VTAIL.n52 185
R1259 VTAIL.n51 VTAIL.n50 185
R1260 VTAIL.n38 VTAIL.n37 185
R1261 VTAIL.n45 VTAIL.n44 185
R1262 VTAIL.n43 VTAIL.n42 185
R1263 VTAIL.n93 VTAIL.t15 147.714
R1264 VTAIL.n9 VTAIL.t17 147.714
R1265 VTAIL.n69 VTAIL.t2 147.714
R1266 VTAIL.n41 VTAIL.t7 147.714
R1267 VTAIL.n96 VTAIL.n95 104.615
R1268 VTAIL.n96 VTAIL.n89 104.615
R1269 VTAIL.n103 VTAIL.n89 104.615
R1270 VTAIL.n104 VTAIL.n103 104.615
R1271 VTAIL.n12 VTAIL.n11 104.615
R1272 VTAIL.n12 VTAIL.n5 104.615
R1273 VTAIL.n19 VTAIL.n5 104.615
R1274 VTAIL.n20 VTAIL.n19 104.615
R1275 VTAIL.n80 VTAIL.n79 104.615
R1276 VTAIL.n79 VTAIL.n65 104.615
R1277 VTAIL.n72 VTAIL.n65 104.615
R1278 VTAIL.n72 VTAIL.n71 104.615
R1279 VTAIL.n52 VTAIL.n51 104.615
R1280 VTAIL.n51 VTAIL.n37 104.615
R1281 VTAIL.n44 VTAIL.n37 104.615
R1282 VTAIL.n44 VTAIL.n43 104.615
R1283 VTAIL.n61 VTAIL.n60 55.7085
R1284 VTAIL.n59 VTAIL.n58 55.7085
R1285 VTAIL.n33 VTAIL.n32 55.7085
R1286 VTAIL.n31 VTAIL.n30 55.7085
R1287 VTAIL.n111 VTAIL.n110 55.7083
R1288 VTAIL.n1 VTAIL.n0 55.7083
R1289 VTAIL.n27 VTAIL.n26 55.7083
R1290 VTAIL.n29 VTAIL.n28 55.7083
R1291 VTAIL.n95 VTAIL.t15 52.3082
R1292 VTAIL.n11 VTAIL.t17 52.3082
R1293 VTAIL.n71 VTAIL.t2 52.3082
R1294 VTAIL.n43 VTAIL.t7 52.3082
R1295 VTAIL.n109 VTAIL.n108 33.9308
R1296 VTAIL.n25 VTAIL.n24 33.9308
R1297 VTAIL.n85 VTAIL.n84 33.9308
R1298 VTAIL.n57 VTAIL.n56 33.9308
R1299 VTAIL.n31 VTAIL.n29 19.41
R1300 VTAIL.n109 VTAIL.n85 17.8927
R1301 VTAIL.n94 VTAIL.n93 15.6631
R1302 VTAIL.n10 VTAIL.n9 15.6631
R1303 VTAIL.n70 VTAIL.n69 15.6631
R1304 VTAIL.n42 VTAIL.n41 15.6631
R1305 VTAIL.n97 VTAIL.n92 12.8005
R1306 VTAIL.n13 VTAIL.n8 12.8005
R1307 VTAIL.n73 VTAIL.n68 12.8005
R1308 VTAIL.n45 VTAIL.n40 12.8005
R1309 VTAIL.n98 VTAIL.n90 12.0247
R1310 VTAIL.n14 VTAIL.n6 12.0247
R1311 VTAIL.n74 VTAIL.n66 12.0247
R1312 VTAIL.n46 VTAIL.n38 12.0247
R1313 VTAIL.n102 VTAIL.n101 11.249
R1314 VTAIL.n18 VTAIL.n17 11.249
R1315 VTAIL.n78 VTAIL.n77 11.249
R1316 VTAIL.n50 VTAIL.n49 11.249
R1317 VTAIL.n105 VTAIL.n88 10.4732
R1318 VTAIL.n21 VTAIL.n4 10.4732
R1319 VTAIL.n81 VTAIL.n64 10.4732
R1320 VTAIL.n53 VTAIL.n36 10.4732
R1321 VTAIL.n106 VTAIL.n86 9.69747
R1322 VTAIL.n22 VTAIL.n2 9.69747
R1323 VTAIL.n82 VTAIL.n62 9.69747
R1324 VTAIL.n54 VTAIL.n34 9.69747
R1325 VTAIL.n108 VTAIL.n107 9.45567
R1326 VTAIL.n24 VTAIL.n23 9.45567
R1327 VTAIL.n84 VTAIL.n83 9.45567
R1328 VTAIL.n56 VTAIL.n55 9.45567
R1329 VTAIL.n107 VTAIL.n106 9.3005
R1330 VTAIL.n88 VTAIL.n87 9.3005
R1331 VTAIL.n101 VTAIL.n100 9.3005
R1332 VTAIL.n99 VTAIL.n98 9.3005
R1333 VTAIL.n92 VTAIL.n91 9.3005
R1334 VTAIL.n23 VTAIL.n22 9.3005
R1335 VTAIL.n4 VTAIL.n3 9.3005
R1336 VTAIL.n17 VTAIL.n16 9.3005
R1337 VTAIL.n15 VTAIL.n14 9.3005
R1338 VTAIL.n8 VTAIL.n7 9.3005
R1339 VTAIL.n83 VTAIL.n82 9.3005
R1340 VTAIL.n64 VTAIL.n63 9.3005
R1341 VTAIL.n77 VTAIL.n76 9.3005
R1342 VTAIL.n75 VTAIL.n74 9.3005
R1343 VTAIL.n68 VTAIL.n67 9.3005
R1344 VTAIL.n55 VTAIL.n54 9.3005
R1345 VTAIL.n36 VTAIL.n35 9.3005
R1346 VTAIL.n49 VTAIL.n48 9.3005
R1347 VTAIL.n47 VTAIL.n46 9.3005
R1348 VTAIL.n40 VTAIL.n39 9.3005
R1349 VTAIL.n93 VTAIL.n91 4.39059
R1350 VTAIL.n9 VTAIL.n7 4.39059
R1351 VTAIL.n69 VTAIL.n67 4.39059
R1352 VTAIL.n41 VTAIL.n39 4.39059
R1353 VTAIL.n108 VTAIL.n86 4.26717
R1354 VTAIL.n24 VTAIL.n2 4.26717
R1355 VTAIL.n84 VTAIL.n62 4.26717
R1356 VTAIL.n56 VTAIL.n34 4.26717
R1357 VTAIL.n110 VTAIL.t13 4.25856
R1358 VTAIL.n110 VTAIL.t11 4.25856
R1359 VTAIL.n0 VTAIL.t12 4.25856
R1360 VTAIL.n0 VTAIL.t14 4.25856
R1361 VTAIL.n26 VTAIL.t5 4.25856
R1362 VTAIL.n26 VTAIL.t3 4.25856
R1363 VTAIL.n28 VTAIL.t0 4.25856
R1364 VTAIL.n28 VTAIL.t1 4.25856
R1365 VTAIL.n60 VTAIL.t18 4.25856
R1366 VTAIL.n60 VTAIL.t6 4.25856
R1367 VTAIL.n58 VTAIL.t4 4.25856
R1368 VTAIL.n58 VTAIL.t19 4.25856
R1369 VTAIL.n32 VTAIL.t9 4.25856
R1370 VTAIL.n32 VTAIL.t10 4.25856
R1371 VTAIL.n30 VTAIL.t8 4.25856
R1372 VTAIL.n30 VTAIL.t16 4.25856
R1373 VTAIL.n106 VTAIL.n105 3.49141
R1374 VTAIL.n22 VTAIL.n21 3.49141
R1375 VTAIL.n82 VTAIL.n81 3.49141
R1376 VTAIL.n54 VTAIL.n53 3.49141
R1377 VTAIL.n102 VTAIL.n88 2.71565
R1378 VTAIL.n18 VTAIL.n4 2.71565
R1379 VTAIL.n78 VTAIL.n64 2.71565
R1380 VTAIL.n50 VTAIL.n36 2.71565
R1381 VTAIL.n101 VTAIL.n90 1.93989
R1382 VTAIL.n17 VTAIL.n6 1.93989
R1383 VTAIL.n77 VTAIL.n66 1.93989
R1384 VTAIL.n49 VTAIL.n38 1.93989
R1385 VTAIL.n33 VTAIL.n31 1.51774
R1386 VTAIL.n57 VTAIL.n33 1.51774
R1387 VTAIL.n61 VTAIL.n59 1.51774
R1388 VTAIL.n85 VTAIL.n61 1.51774
R1389 VTAIL.n29 VTAIL.n27 1.51774
R1390 VTAIL.n27 VTAIL.n25 1.51774
R1391 VTAIL.n111 VTAIL.n109 1.51774
R1392 VTAIL.n59 VTAIL.n57 1.22895
R1393 VTAIL.n25 VTAIL.n1 1.22895
R1394 VTAIL VTAIL.n1 1.19662
R1395 VTAIL.n98 VTAIL.n97 1.16414
R1396 VTAIL.n14 VTAIL.n13 1.16414
R1397 VTAIL.n74 VTAIL.n73 1.16414
R1398 VTAIL.n46 VTAIL.n45 1.16414
R1399 VTAIL.n94 VTAIL.n92 0.388379
R1400 VTAIL.n10 VTAIL.n8 0.388379
R1401 VTAIL.n70 VTAIL.n68 0.388379
R1402 VTAIL.n42 VTAIL.n40 0.388379
R1403 VTAIL VTAIL.n111 0.321621
R1404 VTAIL.n99 VTAIL.n91 0.155672
R1405 VTAIL.n100 VTAIL.n99 0.155672
R1406 VTAIL.n100 VTAIL.n87 0.155672
R1407 VTAIL.n107 VTAIL.n87 0.155672
R1408 VTAIL.n15 VTAIL.n7 0.155672
R1409 VTAIL.n16 VTAIL.n15 0.155672
R1410 VTAIL.n16 VTAIL.n3 0.155672
R1411 VTAIL.n23 VTAIL.n3 0.155672
R1412 VTAIL.n83 VTAIL.n63 0.155672
R1413 VTAIL.n76 VTAIL.n63 0.155672
R1414 VTAIL.n76 VTAIL.n75 0.155672
R1415 VTAIL.n75 VTAIL.n67 0.155672
R1416 VTAIL.n55 VTAIL.n35 0.155672
R1417 VTAIL.n48 VTAIL.n35 0.155672
R1418 VTAIL.n48 VTAIL.n47 0.155672
R1419 VTAIL.n47 VTAIL.n39 0.155672
R1420 VDD2.n45 VDD2.n27 289.615
R1421 VDD2.n18 VDD2.n0 289.615
R1422 VDD2.n46 VDD2.n45 185
R1423 VDD2.n44 VDD2.n43 185
R1424 VDD2.n31 VDD2.n30 185
R1425 VDD2.n38 VDD2.n37 185
R1426 VDD2.n36 VDD2.n35 185
R1427 VDD2.n9 VDD2.n8 185
R1428 VDD2.n11 VDD2.n10 185
R1429 VDD2.n4 VDD2.n3 185
R1430 VDD2.n17 VDD2.n16 185
R1431 VDD2.n19 VDD2.n18 185
R1432 VDD2.n34 VDD2.t1 147.714
R1433 VDD2.n7 VDD2.t0 147.714
R1434 VDD2.n45 VDD2.n44 104.615
R1435 VDD2.n44 VDD2.n30 104.615
R1436 VDD2.n37 VDD2.n30 104.615
R1437 VDD2.n37 VDD2.n36 104.615
R1438 VDD2.n10 VDD2.n9 104.615
R1439 VDD2.n10 VDD2.n3 104.615
R1440 VDD2.n17 VDD2.n3 104.615
R1441 VDD2.n18 VDD2.n17 104.615
R1442 VDD2.n26 VDD2.n25 73.4697
R1443 VDD2 VDD2.n53 73.4668
R1444 VDD2.n52 VDD2.n51 72.3872
R1445 VDD2.n24 VDD2.n23 72.3871
R1446 VDD2.n36 VDD2.t1 52.3082
R1447 VDD2.n9 VDD2.t0 52.3082
R1448 VDD2.n24 VDD2.n22 52.1268
R1449 VDD2.n50 VDD2.n49 50.6096
R1450 VDD2.n50 VDD2.n26 34.9308
R1451 VDD2.n35 VDD2.n34 15.6631
R1452 VDD2.n8 VDD2.n7 15.6631
R1453 VDD2.n38 VDD2.n33 12.8005
R1454 VDD2.n11 VDD2.n6 12.8005
R1455 VDD2.n39 VDD2.n31 12.0247
R1456 VDD2.n12 VDD2.n4 12.0247
R1457 VDD2.n43 VDD2.n42 11.249
R1458 VDD2.n16 VDD2.n15 11.249
R1459 VDD2.n46 VDD2.n29 10.4732
R1460 VDD2.n19 VDD2.n2 10.4732
R1461 VDD2.n47 VDD2.n27 9.69747
R1462 VDD2.n20 VDD2.n0 9.69747
R1463 VDD2.n49 VDD2.n48 9.45567
R1464 VDD2.n22 VDD2.n21 9.45567
R1465 VDD2.n48 VDD2.n47 9.3005
R1466 VDD2.n29 VDD2.n28 9.3005
R1467 VDD2.n42 VDD2.n41 9.3005
R1468 VDD2.n40 VDD2.n39 9.3005
R1469 VDD2.n33 VDD2.n32 9.3005
R1470 VDD2.n21 VDD2.n20 9.3005
R1471 VDD2.n2 VDD2.n1 9.3005
R1472 VDD2.n15 VDD2.n14 9.3005
R1473 VDD2.n13 VDD2.n12 9.3005
R1474 VDD2.n6 VDD2.n5 9.3005
R1475 VDD2.n34 VDD2.n32 4.39059
R1476 VDD2.n7 VDD2.n5 4.39059
R1477 VDD2.n49 VDD2.n27 4.26717
R1478 VDD2.n22 VDD2.n0 4.26717
R1479 VDD2.n53 VDD2.t5 4.25856
R1480 VDD2.n53 VDD2.t6 4.25856
R1481 VDD2.n51 VDD2.t7 4.25856
R1482 VDD2.n51 VDD2.t8 4.25856
R1483 VDD2.n25 VDD2.t4 4.25856
R1484 VDD2.n25 VDD2.t9 4.25856
R1485 VDD2.n23 VDD2.t2 4.25856
R1486 VDD2.n23 VDD2.t3 4.25856
R1487 VDD2.n47 VDD2.n46 3.49141
R1488 VDD2.n20 VDD2.n19 3.49141
R1489 VDD2.n43 VDD2.n29 2.71565
R1490 VDD2.n16 VDD2.n2 2.71565
R1491 VDD2.n42 VDD2.n31 1.93989
R1492 VDD2.n15 VDD2.n4 1.93989
R1493 VDD2.n52 VDD2.n50 1.51774
R1494 VDD2.n39 VDD2.n38 1.16414
R1495 VDD2.n12 VDD2.n11 1.16414
R1496 VDD2 VDD2.n52 0.438
R1497 VDD2.n35 VDD2.n33 0.388379
R1498 VDD2.n8 VDD2.n6 0.388379
R1499 VDD2.n26 VDD2.n24 0.324464
R1500 VDD2.n48 VDD2.n28 0.155672
R1501 VDD2.n41 VDD2.n28 0.155672
R1502 VDD2.n41 VDD2.n40 0.155672
R1503 VDD2.n40 VDD2.n32 0.155672
R1504 VDD2.n13 VDD2.n5 0.155672
R1505 VDD2.n14 VDD2.n13 0.155672
R1506 VDD2.n14 VDD2.n1 0.155672
R1507 VDD2.n21 VDD2.n1 0.155672
R1508 VP.n36 VP.n7 172.555
R1509 VP.n62 VP.n61 172.555
R1510 VP.n35 VP.n34 172.555
R1511 VP.n16 VP.n13 161.3
R1512 VP.n18 VP.n17 161.3
R1513 VP.n19 VP.n12 161.3
R1514 VP.n22 VP.n21 161.3
R1515 VP.n23 VP.n11 161.3
R1516 VP.n25 VP.n24 161.3
R1517 VP.n26 VP.n10 161.3
R1518 VP.n29 VP.n28 161.3
R1519 VP.n30 VP.n9 161.3
R1520 VP.n32 VP.n31 161.3
R1521 VP.n33 VP.n8 161.3
R1522 VP.n60 VP.n0 161.3
R1523 VP.n59 VP.n58 161.3
R1524 VP.n57 VP.n1 161.3
R1525 VP.n56 VP.n55 161.3
R1526 VP.n53 VP.n2 161.3
R1527 VP.n52 VP.n51 161.3
R1528 VP.n50 VP.n3 161.3
R1529 VP.n49 VP.n48 161.3
R1530 VP.n46 VP.n4 161.3
R1531 VP.n45 VP.n44 161.3
R1532 VP.n43 VP.n5 161.3
R1533 VP.n42 VP.n41 161.3
R1534 VP.n39 VP.n6 161.3
R1535 VP.n38 VP.n37 161.3
R1536 VP.n15 VP.t2 107.415
R1537 VP.n7 VP.t1 78.3676
R1538 VP.n40 VP.t0 78.3676
R1539 VP.n47 VP.t7 78.3676
R1540 VP.n54 VP.t3 78.3676
R1541 VP.n61 VP.t4 78.3676
R1542 VP.n34 VP.t5 78.3676
R1543 VP.n27 VP.t9 78.3676
R1544 VP.n20 VP.t8 78.3676
R1545 VP.n14 VP.t6 78.3676
R1546 VP.n15 VP.n14 65.4496
R1547 VP.n46 VP.n45 53.1199
R1548 VP.n53 VP.n52 53.1199
R1549 VP.n26 VP.n25 53.1199
R1550 VP.n19 VP.n18 53.1199
R1551 VP.n41 VP.n39 51.1773
R1552 VP.n59 VP.n1 51.1773
R1553 VP.n32 VP.n9 51.1773
R1554 VP.n36 VP.n35 41.1444
R1555 VP.n39 VP.n38 29.8095
R1556 VP.n60 VP.n59 29.8095
R1557 VP.n33 VP.n32 29.8095
R1558 VP.n48 VP.n46 27.8669
R1559 VP.n52 VP.n3 27.8669
R1560 VP.n25 VP.n11 27.8669
R1561 VP.n21 VP.n19 27.8669
R1562 VP.n16 VP.n15 27.1884
R1563 VP.n45 VP.n5 24.4675
R1564 VP.n55 VP.n53 24.4675
R1565 VP.n28 VP.n26 24.4675
R1566 VP.n18 VP.n13 24.4675
R1567 VP.n41 VP.n40 23.9782
R1568 VP.n54 VP.n1 23.9782
R1569 VP.n27 VP.n9 23.9782
R1570 VP.n38 VP.n7 13.2127
R1571 VP.n61 VP.n60 13.2127
R1572 VP.n34 VP.n33 13.2127
R1573 VP.n48 VP.n47 12.234
R1574 VP.n47 VP.n3 12.234
R1575 VP.n21 VP.n20 12.234
R1576 VP.n20 VP.n11 12.234
R1577 VP.n40 VP.n5 0.48984
R1578 VP.n55 VP.n54 0.48984
R1579 VP.n28 VP.n27 0.48984
R1580 VP.n14 VP.n13 0.48984
R1581 VP.n17 VP.n16 0.189894
R1582 VP.n17 VP.n12 0.189894
R1583 VP.n22 VP.n12 0.189894
R1584 VP.n23 VP.n22 0.189894
R1585 VP.n24 VP.n23 0.189894
R1586 VP.n24 VP.n10 0.189894
R1587 VP.n29 VP.n10 0.189894
R1588 VP.n30 VP.n29 0.189894
R1589 VP.n31 VP.n30 0.189894
R1590 VP.n31 VP.n8 0.189894
R1591 VP.n35 VP.n8 0.189894
R1592 VP.n37 VP.n36 0.189894
R1593 VP.n37 VP.n6 0.189894
R1594 VP.n42 VP.n6 0.189894
R1595 VP.n43 VP.n42 0.189894
R1596 VP.n44 VP.n43 0.189894
R1597 VP.n44 VP.n4 0.189894
R1598 VP.n49 VP.n4 0.189894
R1599 VP.n50 VP.n49 0.189894
R1600 VP.n51 VP.n50 0.189894
R1601 VP.n51 VP.n2 0.189894
R1602 VP.n56 VP.n2 0.189894
R1603 VP.n57 VP.n56 0.189894
R1604 VP.n58 VP.n57 0.189894
R1605 VP.n58 VP.n0 0.189894
R1606 VP.n62 VP.n0 0.189894
R1607 VP VP.n62 0.0516364
R1608 VDD1.n18 VDD1.n0 289.615
R1609 VDD1.n43 VDD1.n25 289.615
R1610 VDD1.n19 VDD1.n18 185
R1611 VDD1.n17 VDD1.n16 185
R1612 VDD1.n4 VDD1.n3 185
R1613 VDD1.n11 VDD1.n10 185
R1614 VDD1.n9 VDD1.n8 185
R1615 VDD1.n34 VDD1.n33 185
R1616 VDD1.n36 VDD1.n35 185
R1617 VDD1.n29 VDD1.n28 185
R1618 VDD1.n42 VDD1.n41 185
R1619 VDD1.n44 VDD1.n43 185
R1620 VDD1.n7 VDD1.t7 147.714
R1621 VDD1.n32 VDD1.t8 147.714
R1622 VDD1.n18 VDD1.n17 104.615
R1623 VDD1.n17 VDD1.n3 104.615
R1624 VDD1.n10 VDD1.n3 104.615
R1625 VDD1.n10 VDD1.n9 104.615
R1626 VDD1.n35 VDD1.n34 104.615
R1627 VDD1.n35 VDD1.n28 104.615
R1628 VDD1.n42 VDD1.n28 104.615
R1629 VDD1.n43 VDD1.n42 104.615
R1630 VDD1.n51 VDD1.n50 73.4697
R1631 VDD1.n24 VDD1.n23 72.3872
R1632 VDD1.n53 VDD1.n52 72.3871
R1633 VDD1.n49 VDD1.n48 72.3871
R1634 VDD1.n9 VDD1.t7 52.3082
R1635 VDD1.n34 VDD1.t8 52.3082
R1636 VDD1.n24 VDD1.n22 52.1268
R1637 VDD1.n49 VDD1.n47 52.1268
R1638 VDD1.n53 VDD1.n51 36.2724
R1639 VDD1.n8 VDD1.n7 15.6631
R1640 VDD1.n33 VDD1.n32 15.6631
R1641 VDD1.n11 VDD1.n6 12.8005
R1642 VDD1.n36 VDD1.n31 12.8005
R1643 VDD1.n12 VDD1.n4 12.0247
R1644 VDD1.n37 VDD1.n29 12.0247
R1645 VDD1.n16 VDD1.n15 11.249
R1646 VDD1.n41 VDD1.n40 11.249
R1647 VDD1.n19 VDD1.n2 10.4732
R1648 VDD1.n44 VDD1.n27 10.4732
R1649 VDD1.n20 VDD1.n0 9.69747
R1650 VDD1.n45 VDD1.n25 9.69747
R1651 VDD1.n22 VDD1.n21 9.45567
R1652 VDD1.n47 VDD1.n46 9.45567
R1653 VDD1.n21 VDD1.n20 9.3005
R1654 VDD1.n2 VDD1.n1 9.3005
R1655 VDD1.n15 VDD1.n14 9.3005
R1656 VDD1.n13 VDD1.n12 9.3005
R1657 VDD1.n6 VDD1.n5 9.3005
R1658 VDD1.n46 VDD1.n45 9.3005
R1659 VDD1.n27 VDD1.n26 9.3005
R1660 VDD1.n40 VDD1.n39 9.3005
R1661 VDD1.n38 VDD1.n37 9.3005
R1662 VDD1.n31 VDD1.n30 9.3005
R1663 VDD1.n7 VDD1.n5 4.39059
R1664 VDD1.n32 VDD1.n30 4.39059
R1665 VDD1.n22 VDD1.n0 4.26717
R1666 VDD1.n47 VDD1.n25 4.26717
R1667 VDD1.n52 VDD1.t0 4.25856
R1668 VDD1.n52 VDD1.t4 4.25856
R1669 VDD1.n23 VDD1.t3 4.25856
R1670 VDD1.n23 VDD1.t1 4.25856
R1671 VDD1.n50 VDD1.t6 4.25856
R1672 VDD1.n50 VDD1.t5 4.25856
R1673 VDD1.n48 VDD1.t9 4.25856
R1674 VDD1.n48 VDD1.t2 4.25856
R1675 VDD1.n20 VDD1.n19 3.49141
R1676 VDD1.n45 VDD1.n44 3.49141
R1677 VDD1.n16 VDD1.n2 2.71565
R1678 VDD1.n41 VDD1.n27 2.71565
R1679 VDD1.n15 VDD1.n4 1.93989
R1680 VDD1.n40 VDD1.n29 1.93989
R1681 VDD1.n12 VDD1.n11 1.16414
R1682 VDD1.n37 VDD1.n36 1.16414
R1683 VDD1 VDD1.n53 1.08024
R1684 VDD1 VDD1.n24 0.438
R1685 VDD1.n8 VDD1.n6 0.388379
R1686 VDD1.n33 VDD1.n31 0.388379
R1687 VDD1.n51 VDD1.n49 0.324464
R1688 VDD1.n21 VDD1.n1 0.155672
R1689 VDD1.n14 VDD1.n1 0.155672
R1690 VDD1.n14 VDD1.n13 0.155672
R1691 VDD1.n13 VDD1.n5 0.155672
R1692 VDD1.n38 VDD1.n30 0.155672
R1693 VDD1.n39 VDD1.n38 0.155672
R1694 VDD1.n39 VDD1.n26 0.155672
R1695 VDD1.n46 VDD1.n26 0.155672
C0 VTAIL VDD2 6.40751f
C1 VTAIL VDD1 6.36345f
C2 VP VTAIL 4.42534f
C3 VN VDD2 3.82358f
C4 VN VDD1 0.154617f
C5 VP VN 5.31116f
C6 VDD2 VDD1 1.41218f
C7 VN VTAIL 4.41111f
C8 VP VDD2 0.437957f
C9 VP VDD1 4.10421f
C10 VDD2 B 4.524367f
C11 VDD1 B 4.493844f
C12 VTAIL B 4.147271f
C13 VN B 11.85238f
C14 VP B 10.359131f
C15 VDD1.n0 B 0.033085f
C16 VDD1.n1 B 0.023425f
C17 VDD1.n2 B 0.012588f
C18 VDD1.n3 B 0.029753f
C19 VDD1.n4 B 0.013328f
C20 VDD1.n5 B 0.411059f
C21 VDD1.n6 B 0.012588f
C22 VDD1.t7 B 0.048876f
C23 VDD1.n7 B 0.093232f
C24 VDD1.n8 B 0.017559f
C25 VDD1.n9 B 0.022315f
C26 VDD1.n10 B 0.029753f
C27 VDD1.n11 B 0.013328f
C28 VDD1.n12 B 0.012588f
C29 VDD1.n13 B 0.023425f
C30 VDD1.n14 B 0.023425f
C31 VDD1.n15 B 0.012588f
C32 VDD1.n16 B 0.013328f
C33 VDD1.n17 B 0.029753f
C34 VDD1.n18 B 0.06469f
C35 VDD1.n19 B 0.013328f
C36 VDD1.n20 B 0.012588f
C37 VDD1.n21 B 0.057027f
C38 VDD1.n22 B 0.057159f
C39 VDD1.t3 B 0.086078f
C40 VDD1.t1 B 0.086078f
C41 VDD1.n23 B 0.693436f
C42 VDD1.n24 B 0.489354f
C43 VDD1.n25 B 0.033085f
C44 VDD1.n26 B 0.023425f
C45 VDD1.n27 B 0.012588f
C46 VDD1.n28 B 0.029753f
C47 VDD1.n29 B 0.013328f
C48 VDD1.n30 B 0.411059f
C49 VDD1.n31 B 0.012588f
C50 VDD1.t8 B 0.048876f
C51 VDD1.n32 B 0.093232f
C52 VDD1.n33 B 0.017559f
C53 VDD1.n34 B 0.022315f
C54 VDD1.n35 B 0.029753f
C55 VDD1.n36 B 0.013328f
C56 VDD1.n37 B 0.012588f
C57 VDD1.n38 B 0.023425f
C58 VDD1.n39 B 0.023425f
C59 VDD1.n40 B 0.012588f
C60 VDD1.n41 B 0.013328f
C61 VDD1.n42 B 0.029753f
C62 VDD1.n43 B 0.06469f
C63 VDD1.n44 B 0.013328f
C64 VDD1.n45 B 0.012588f
C65 VDD1.n46 B 0.057027f
C66 VDD1.n47 B 0.057159f
C67 VDD1.t9 B 0.086078f
C68 VDD1.t2 B 0.086078f
C69 VDD1.n48 B 0.693433f
C70 VDD1.n49 B 0.482463f
C71 VDD1.t6 B 0.086078f
C72 VDD1.t5 B 0.086078f
C73 VDD1.n50 B 0.6992f
C74 VDD1.n51 B 1.81279f
C75 VDD1.t0 B 0.086078f
C76 VDD1.t4 B 0.086078f
C77 VDD1.n52 B 0.693433f
C78 VDD1.n53 B 1.97116f
C79 VP.n0 B 0.034247f
C80 VP.t4 B 0.592453f
C81 VP.n1 B 0.061551f
C82 VP.n2 B 0.034247f
C83 VP.n3 B 0.051376f
C84 VP.n4 B 0.034247f
C85 VP.n5 B 0.032946f
C86 VP.n6 B 0.034247f
C87 VP.t1 B 0.592453f
C88 VP.n7 B 0.315695f
C89 VP.n8 B 0.034247f
C90 VP.t5 B 0.592453f
C91 VP.n9 B 0.061551f
C92 VP.n10 B 0.034247f
C93 VP.n11 B 0.051376f
C94 VP.n12 B 0.034247f
C95 VP.n13 B 0.032946f
C96 VP.t2 B 0.690651f
C97 VP.t6 B 0.592453f
C98 VP.n14 B 0.291067f
C99 VP.n15 B 0.321147f
C100 VP.n16 B 0.18437f
C101 VP.n17 B 0.034247f
C102 VP.n18 B 0.060766f
C103 VP.n19 B 0.03592f
C104 VP.t8 B 0.592453f
C105 VP.n20 B 0.244247f
C106 VP.n21 B 0.051376f
C107 VP.n22 B 0.034247f
C108 VP.n23 B 0.034247f
C109 VP.n24 B 0.034247f
C110 VP.n25 B 0.03592f
C111 VP.n26 B 0.060766f
C112 VP.t9 B 0.592453f
C113 VP.n27 B 0.244247f
C114 VP.n28 B 0.032946f
C115 VP.n29 B 0.034247f
C116 VP.n30 B 0.034247f
C117 VP.n31 B 0.034247f
C118 VP.n32 B 0.033406f
C119 VP.n33 B 0.053736f
C120 VP.n34 B 0.315695f
C121 VP.n35 B 1.37062f
C122 VP.n36 B 1.40054f
C123 VP.n37 B 0.034247f
C124 VP.n38 B 0.053736f
C125 VP.n39 B 0.033406f
C126 VP.t0 B 0.592453f
C127 VP.n40 B 0.244247f
C128 VP.n41 B 0.061551f
C129 VP.n42 B 0.034247f
C130 VP.n43 B 0.034247f
C131 VP.n44 B 0.034247f
C132 VP.n45 B 0.060766f
C133 VP.n46 B 0.03592f
C134 VP.t7 B 0.592453f
C135 VP.n47 B 0.244247f
C136 VP.n48 B 0.051376f
C137 VP.n49 B 0.034247f
C138 VP.n50 B 0.034247f
C139 VP.n51 B 0.034247f
C140 VP.n52 B 0.03592f
C141 VP.n53 B 0.060766f
C142 VP.t3 B 0.592453f
C143 VP.n54 B 0.244247f
C144 VP.n55 B 0.032946f
C145 VP.n56 B 0.034247f
C146 VP.n57 B 0.034247f
C147 VP.n58 B 0.034247f
C148 VP.n59 B 0.033406f
C149 VP.n60 B 0.053736f
C150 VP.n61 B 0.315695f
C151 VP.n62 B 0.031526f
C152 VDD2.n0 B 0.032406f
C153 VDD2.n1 B 0.022945f
C154 VDD2.n2 B 0.01233f
C155 VDD2.n3 B 0.029143f
C156 VDD2.n4 B 0.013055f
C157 VDD2.n5 B 0.402632f
C158 VDD2.n6 B 0.01233f
C159 VDD2.t0 B 0.047874f
C160 VDD2.n7 B 0.091321f
C161 VDD2.n8 B 0.017199f
C162 VDD2.n9 B 0.021857f
C163 VDD2.n10 B 0.029143f
C164 VDD2.n11 B 0.013055f
C165 VDD2.n12 B 0.01233f
C166 VDD2.n13 B 0.022945f
C167 VDD2.n14 B 0.022945f
C168 VDD2.n15 B 0.01233f
C169 VDD2.n16 B 0.013055f
C170 VDD2.n17 B 0.029143f
C171 VDD2.n18 B 0.063363f
C172 VDD2.n19 B 0.013055f
C173 VDD2.n20 B 0.01233f
C174 VDD2.n21 B 0.055858f
C175 VDD2.n22 B 0.055987f
C176 VDD2.t2 B 0.084314f
C177 VDD2.t3 B 0.084314f
C178 VDD2.n23 B 0.679217f
C179 VDD2.n24 B 0.472573f
C180 VDD2.t4 B 0.084314f
C181 VDD2.t9 B 0.084314f
C182 VDD2.n25 B 0.684866f
C183 VDD2.n26 B 1.69303f
C184 VDD2.n27 B 0.032406f
C185 VDD2.n28 B 0.022945f
C186 VDD2.n29 B 0.01233f
C187 VDD2.n30 B 0.029143f
C188 VDD2.n31 B 0.013055f
C189 VDD2.n32 B 0.402632f
C190 VDD2.n33 B 0.01233f
C191 VDD2.t1 B 0.047874f
C192 VDD2.n34 B 0.091321f
C193 VDD2.n35 B 0.017199f
C194 VDD2.n36 B 0.021857f
C195 VDD2.n37 B 0.029143f
C196 VDD2.n38 B 0.013055f
C197 VDD2.n39 B 0.01233f
C198 VDD2.n40 B 0.022945f
C199 VDD2.n41 B 0.022945f
C200 VDD2.n42 B 0.01233f
C201 VDD2.n43 B 0.013055f
C202 VDD2.n44 B 0.029143f
C203 VDD2.n45 B 0.063363f
C204 VDD2.n46 B 0.013055f
C205 VDD2.n47 B 0.01233f
C206 VDD2.n48 B 0.055858f
C207 VDD2.n49 B 0.051389f
C208 VDD2.n50 B 1.7039f
C209 VDD2.t7 B 0.084314f
C210 VDD2.t8 B 0.084314f
C211 VDD2.n51 B 0.67922f
C212 VDD2.n52 B 0.325945f
C213 VDD2.t5 B 0.084314f
C214 VDD2.t6 B 0.084314f
C215 VDD2.n53 B 0.684841f
C216 VTAIL.t12 B 0.104152f
C217 VTAIL.t14 B 0.104152f
C218 VTAIL.n0 B 0.77355f
C219 VTAIL.n1 B 0.472511f
C220 VTAIL.n2 B 0.040031f
C221 VTAIL.n3 B 0.028344f
C222 VTAIL.n4 B 0.015231f
C223 VTAIL.n5 B 0.036f
C224 VTAIL.n6 B 0.016127f
C225 VTAIL.n7 B 0.497369f
C226 VTAIL.n8 B 0.015231f
C227 VTAIL.t17 B 0.059139f
C228 VTAIL.n9 B 0.112808f
C229 VTAIL.n10 B 0.021245f
C230 VTAIL.n11 B 0.027f
C231 VTAIL.n12 B 0.036f
C232 VTAIL.n13 B 0.016127f
C233 VTAIL.n14 B 0.015231f
C234 VTAIL.n15 B 0.028344f
C235 VTAIL.n16 B 0.028344f
C236 VTAIL.n17 B 0.015231f
C237 VTAIL.n18 B 0.016127f
C238 VTAIL.n19 B 0.036f
C239 VTAIL.n20 B 0.078273f
C240 VTAIL.n21 B 0.016127f
C241 VTAIL.n22 B 0.015231f
C242 VTAIL.n23 B 0.069001f
C243 VTAIL.n24 B 0.043936f
C244 VTAIL.n25 B 0.276944f
C245 VTAIL.t5 B 0.104152f
C246 VTAIL.t3 B 0.104152f
C247 VTAIL.n26 B 0.77355f
C248 VTAIL.n27 B 0.528215f
C249 VTAIL.t0 B 0.104152f
C250 VTAIL.t1 B 0.104152f
C251 VTAIL.n28 B 0.77355f
C252 VTAIL.n29 B 1.41792f
C253 VTAIL.t8 B 0.104152f
C254 VTAIL.t16 B 0.104152f
C255 VTAIL.n30 B 0.773556f
C256 VTAIL.n31 B 1.41791f
C257 VTAIL.t9 B 0.104152f
C258 VTAIL.t10 B 0.104152f
C259 VTAIL.n32 B 0.773556f
C260 VTAIL.n33 B 0.52821f
C261 VTAIL.n34 B 0.040031f
C262 VTAIL.n35 B 0.028344f
C263 VTAIL.n36 B 0.015231f
C264 VTAIL.n37 B 0.036f
C265 VTAIL.n38 B 0.016127f
C266 VTAIL.n39 B 0.497369f
C267 VTAIL.n40 B 0.015231f
C268 VTAIL.t7 B 0.059139f
C269 VTAIL.n41 B 0.112808f
C270 VTAIL.n42 B 0.021245f
C271 VTAIL.n43 B 0.027f
C272 VTAIL.n44 B 0.036f
C273 VTAIL.n45 B 0.016127f
C274 VTAIL.n46 B 0.015231f
C275 VTAIL.n47 B 0.028344f
C276 VTAIL.n48 B 0.028344f
C277 VTAIL.n49 B 0.015231f
C278 VTAIL.n50 B 0.016127f
C279 VTAIL.n51 B 0.036f
C280 VTAIL.n52 B 0.078273f
C281 VTAIL.n53 B 0.016127f
C282 VTAIL.n54 B 0.015231f
C283 VTAIL.n55 B 0.069001f
C284 VTAIL.n56 B 0.043936f
C285 VTAIL.n57 B 0.276944f
C286 VTAIL.t4 B 0.104152f
C287 VTAIL.t19 B 0.104152f
C288 VTAIL.n58 B 0.773556f
C289 VTAIL.n59 B 0.501834f
C290 VTAIL.t18 B 0.104152f
C291 VTAIL.t6 B 0.104152f
C292 VTAIL.n60 B 0.773556f
C293 VTAIL.n61 B 0.52821f
C294 VTAIL.n62 B 0.040031f
C295 VTAIL.n63 B 0.028344f
C296 VTAIL.n64 B 0.015231f
C297 VTAIL.n65 B 0.036f
C298 VTAIL.n66 B 0.016127f
C299 VTAIL.n67 B 0.497369f
C300 VTAIL.n68 B 0.015231f
C301 VTAIL.t2 B 0.059139f
C302 VTAIL.n69 B 0.112808f
C303 VTAIL.n70 B 0.021245f
C304 VTAIL.n71 B 0.027f
C305 VTAIL.n72 B 0.036f
C306 VTAIL.n73 B 0.016127f
C307 VTAIL.n74 B 0.015231f
C308 VTAIL.n75 B 0.028344f
C309 VTAIL.n76 B 0.028344f
C310 VTAIL.n77 B 0.015231f
C311 VTAIL.n78 B 0.016127f
C312 VTAIL.n79 B 0.036f
C313 VTAIL.n80 B 0.078273f
C314 VTAIL.n81 B 0.016127f
C315 VTAIL.n82 B 0.015231f
C316 VTAIL.n83 B 0.069001f
C317 VTAIL.n84 B 0.043936f
C318 VTAIL.n85 B 1.05445f
C319 VTAIL.n86 B 0.040031f
C320 VTAIL.n87 B 0.028344f
C321 VTAIL.n88 B 0.015231f
C322 VTAIL.n89 B 0.036f
C323 VTAIL.n90 B 0.016127f
C324 VTAIL.n91 B 0.497369f
C325 VTAIL.n92 B 0.015231f
C326 VTAIL.t15 B 0.059139f
C327 VTAIL.n93 B 0.112808f
C328 VTAIL.n94 B 0.021245f
C329 VTAIL.n95 B 0.027f
C330 VTAIL.n96 B 0.036f
C331 VTAIL.n97 B 0.016127f
C332 VTAIL.n98 B 0.015231f
C333 VTAIL.n99 B 0.028344f
C334 VTAIL.n100 B 0.028344f
C335 VTAIL.n101 B 0.015231f
C336 VTAIL.n102 B 0.016127f
C337 VTAIL.n103 B 0.036f
C338 VTAIL.n104 B 0.078273f
C339 VTAIL.n105 B 0.016127f
C340 VTAIL.n106 B 0.015231f
C341 VTAIL.n107 B 0.069001f
C342 VTAIL.n108 B 0.043936f
C343 VTAIL.n109 B 1.05445f
C344 VTAIL.t13 B 0.104152f
C345 VTAIL.t11 B 0.104152f
C346 VTAIL.n110 B 0.77355f
C347 VTAIL.n111 B 0.418972f
C348 VN.n0 B 0.033387f
C349 VN.t0 B 0.577559f
C350 VN.n1 B 0.060004f
C351 VN.n2 B 0.033387f
C352 VN.n3 B 0.050085f
C353 VN.n4 B 0.033387f
C354 VN.n5 B 0.032118f
C355 VN.t9 B 0.673288f
C356 VN.t7 B 0.577559f
C357 VN.n6 B 0.283749f
C358 VN.n7 B 0.313073f
C359 VN.n8 B 0.179734f
C360 VN.n9 B 0.033387f
C361 VN.n10 B 0.059239f
C362 VN.n11 B 0.035017f
C363 VN.t6 B 0.577559f
C364 VN.n12 B 0.238106f
C365 VN.n13 B 0.050085f
C366 VN.n14 B 0.033387f
C367 VN.n15 B 0.033387f
C368 VN.n16 B 0.033387f
C369 VN.n17 B 0.035017f
C370 VN.n18 B 0.059239f
C371 VN.t5 B 0.577559f
C372 VN.n19 B 0.238106f
C373 VN.n20 B 0.032118f
C374 VN.n21 B 0.033387f
C375 VN.n22 B 0.033387f
C376 VN.n23 B 0.033387f
C377 VN.n24 B 0.032567f
C378 VN.n25 B 0.052385f
C379 VN.n26 B 0.307758f
C380 VN.n27 B 0.030733f
C381 VN.n28 B 0.033387f
C382 VN.t8 B 0.577559f
C383 VN.n29 B 0.060004f
C384 VN.n30 B 0.033387f
C385 VN.t2 B 0.577559f
C386 VN.n31 B 0.238106f
C387 VN.n32 B 0.050085f
C388 VN.n33 B 0.033387f
C389 VN.t1 B 0.577559f
C390 VN.n34 B 0.238106f
C391 VN.n35 B 0.032118f
C392 VN.t3 B 0.673288f
C393 VN.t4 B 0.577559f
C394 VN.n36 B 0.283749f
C395 VN.n37 B 0.313073f
C396 VN.n38 B 0.179734f
C397 VN.n39 B 0.033387f
C398 VN.n40 B 0.059239f
C399 VN.n41 B 0.035017f
C400 VN.n42 B 0.050085f
C401 VN.n43 B 0.033387f
C402 VN.n44 B 0.033387f
C403 VN.n45 B 0.033387f
C404 VN.n46 B 0.035017f
C405 VN.n47 B 0.059239f
C406 VN.n48 B 0.032118f
C407 VN.n49 B 0.033387f
C408 VN.n50 B 0.033387f
C409 VN.n51 B 0.033387f
C410 VN.n52 B 0.032567f
C411 VN.n53 B 0.052385f
C412 VN.n54 B 0.307758f
C413 VN.n55 B 1.35811f
.ends

