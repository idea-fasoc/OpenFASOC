* NGSPICE file created from diff_pair_sample_0041.ext - technology: sky130A

.subckt diff_pair_sample_0041 VTAIL VN VP B VDD2 VDD1
X0 B.t11 B.t9 B.t10 w_n2314_n4716# sky130_fd_pr__pfet_01v8 ad=7.3086 pd=38.26 as=0 ps=0 w=18.74 l=1.91
X1 VTAIL.t7 VN.t0 VDD2.t0 w_n2314_n4716# sky130_fd_pr__pfet_01v8 ad=7.3086 pd=38.26 as=3.0921 ps=19.07 w=18.74 l=1.91
X2 VDD2.t2 VN.t1 VTAIL.t6 w_n2314_n4716# sky130_fd_pr__pfet_01v8 ad=3.0921 pd=19.07 as=7.3086 ps=38.26 w=18.74 l=1.91
X3 VDD1.t3 VP.t0 VTAIL.t1 w_n2314_n4716# sky130_fd_pr__pfet_01v8 ad=3.0921 pd=19.07 as=7.3086 ps=38.26 w=18.74 l=1.91
X4 VDD1.t2 VP.t1 VTAIL.t3 w_n2314_n4716# sky130_fd_pr__pfet_01v8 ad=3.0921 pd=19.07 as=7.3086 ps=38.26 w=18.74 l=1.91
X5 VTAIL.t0 VP.t2 VDD1.t1 w_n2314_n4716# sky130_fd_pr__pfet_01v8 ad=7.3086 pd=38.26 as=3.0921 ps=19.07 w=18.74 l=1.91
X6 VDD2.t1 VN.t2 VTAIL.t5 w_n2314_n4716# sky130_fd_pr__pfet_01v8 ad=3.0921 pd=19.07 as=7.3086 ps=38.26 w=18.74 l=1.91
X7 VTAIL.t4 VN.t3 VDD2.t3 w_n2314_n4716# sky130_fd_pr__pfet_01v8 ad=7.3086 pd=38.26 as=3.0921 ps=19.07 w=18.74 l=1.91
X8 B.t8 B.t6 B.t7 w_n2314_n4716# sky130_fd_pr__pfet_01v8 ad=7.3086 pd=38.26 as=0 ps=0 w=18.74 l=1.91
X9 B.t5 B.t3 B.t4 w_n2314_n4716# sky130_fd_pr__pfet_01v8 ad=7.3086 pd=38.26 as=0 ps=0 w=18.74 l=1.91
X10 B.t2 B.t0 B.t1 w_n2314_n4716# sky130_fd_pr__pfet_01v8 ad=7.3086 pd=38.26 as=0 ps=0 w=18.74 l=1.91
X11 VTAIL.t2 VP.t3 VDD1.t0 w_n2314_n4716# sky130_fd_pr__pfet_01v8 ad=7.3086 pd=38.26 as=3.0921 ps=19.07 w=18.74 l=1.91
R0 B.n526 B.n525 585
R1 B.n527 B.n86 585
R2 B.n529 B.n528 585
R3 B.n530 B.n85 585
R4 B.n532 B.n531 585
R5 B.n533 B.n84 585
R6 B.n535 B.n534 585
R7 B.n536 B.n83 585
R8 B.n538 B.n537 585
R9 B.n539 B.n82 585
R10 B.n541 B.n540 585
R11 B.n542 B.n81 585
R12 B.n544 B.n543 585
R13 B.n545 B.n80 585
R14 B.n547 B.n546 585
R15 B.n548 B.n79 585
R16 B.n550 B.n549 585
R17 B.n551 B.n78 585
R18 B.n553 B.n552 585
R19 B.n554 B.n77 585
R20 B.n556 B.n555 585
R21 B.n557 B.n76 585
R22 B.n559 B.n558 585
R23 B.n560 B.n75 585
R24 B.n562 B.n561 585
R25 B.n563 B.n74 585
R26 B.n565 B.n564 585
R27 B.n566 B.n73 585
R28 B.n568 B.n567 585
R29 B.n569 B.n72 585
R30 B.n571 B.n570 585
R31 B.n572 B.n71 585
R32 B.n574 B.n573 585
R33 B.n575 B.n70 585
R34 B.n577 B.n576 585
R35 B.n578 B.n69 585
R36 B.n580 B.n579 585
R37 B.n581 B.n68 585
R38 B.n583 B.n582 585
R39 B.n584 B.n67 585
R40 B.n586 B.n585 585
R41 B.n587 B.n66 585
R42 B.n589 B.n588 585
R43 B.n590 B.n65 585
R44 B.n592 B.n591 585
R45 B.n593 B.n64 585
R46 B.n595 B.n594 585
R47 B.n596 B.n63 585
R48 B.n598 B.n597 585
R49 B.n599 B.n62 585
R50 B.n601 B.n600 585
R51 B.n602 B.n61 585
R52 B.n604 B.n603 585
R53 B.n605 B.n60 585
R54 B.n607 B.n606 585
R55 B.n608 B.n59 585
R56 B.n610 B.n609 585
R57 B.n611 B.n58 585
R58 B.n613 B.n612 585
R59 B.n614 B.n57 585
R60 B.n616 B.n615 585
R61 B.n618 B.n54 585
R62 B.n620 B.n619 585
R63 B.n621 B.n53 585
R64 B.n623 B.n622 585
R65 B.n624 B.n52 585
R66 B.n626 B.n625 585
R67 B.n627 B.n51 585
R68 B.n629 B.n628 585
R69 B.n630 B.n47 585
R70 B.n632 B.n631 585
R71 B.n633 B.n46 585
R72 B.n635 B.n634 585
R73 B.n636 B.n45 585
R74 B.n638 B.n637 585
R75 B.n639 B.n44 585
R76 B.n641 B.n640 585
R77 B.n642 B.n43 585
R78 B.n644 B.n643 585
R79 B.n645 B.n42 585
R80 B.n647 B.n646 585
R81 B.n648 B.n41 585
R82 B.n650 B.n649 585
R83 B.n651 B.n40 585
R84 B.n653 B.n652 585
R85 B.n654 B.n39 585
R86 B.n656 B.n655 585
R87 B.n657 B.n38 585
R88 B.n659 B.n658 585
R89 B.n660 B.n37 585
R90 B.n662 B.n661 585
R91 B.n663 B.n36 585
R92 B.n665 B.n664 585
R93 B.n666 B.n35 585
R94 B.n668 B.n667 585
R95 B.n669 B.n34 585
R96 B.n671 B.n670 585
R97 B.n672 B.n33 585
R98 B.n674 B.n673 585
R99 B.n675 B.n32 585
R100 B.n677 B.n676 585
R101 B.n678 B.n31 585
R102 B.n680 B.n679 585
R103 B.n681 B.n30 585
R104 B.n683 B.n682 585
R105 B.n684 B.n29 585
R106 B.n686 B.n685 585
R107 B.n687 B.n28 585
R108 B.n689 B.n688 585
R109 B.n690 B.n27 585
R110 B.n692 B.n691 585
R111 B.n693 B.n26 585
R112 B.n695 B.n694 585
R113 B.n696 B.n25 585
R114 B.n698 B.n697 585
R115 B.n699 B.n24 585
R116 B.n701 B.n700 585
R117 B.n702 B.n23 585
R118 B.n704 B.n703 585
R119 B.n705 B.n22 585
R120 B.n707 B.n706 585
R121 B.n708 B.n21 585
R122 B.n710 B.n709 585
R123 B.n711 B.n20 585
R124 B.n713 B.n712 585
R125 B.n714 B.n19 585
R126 B.n716 B.n715 585
R127 B.n717 B.n18 585
R128 B.n719 B.n718 585
R129 B.n720 B.n17 585
R130 B.n722 B.n721 585
R131 B.n723 B.n16 585
R132 B.n524 B.n87 585
R133 B.n523 B.n522 585
R134 B.n521 B.n88 585
R135 B.n520 B.n519 585
R136 B.n518 B.n89 585
R137 B.n517 B.n516 585
R138 B.n515 B.n90 585
R139 B.n514 B.n513 585
R140 B.n512 B.n91 585
R141 B.n511 B.n510 585
R142 B.n509 B.n92 585
R143 B.n508 B.n507 585
R144 B.n506 B.n93 585
R145 B.n505 B.n504 585
R146 B.n503 B.n94 585
R147 B.n502 B.n501 585
R148 B.n500 B.n95 585
R149 B.n499 B.n498 585
R150 B.n497 B.n96 585
R151 B.n496 B.n495 585
R152 B.n494 B.n97 585
R153 B.n493 B.n492 585
R154 B.n491 B.n98 585
R155 B.n490 B.n489 585
R156 B.n488 B.n99 585
R157 B.n487 B.n486 585
R158 B.n485 B.n100 585
R159 B.n484 B.n483 585
R160 B.n482 B.n101 585
R161 B.n481 B.n480 585
R162 B.n479 B.n102 585
R163 B.n478 B.n477 585
R164 B.n476 B.n103 585
R165 B.n475 B.n474 585
R166 B.n473 B.n104 585
R167 B.n472 B.n471 585
R168 B.n470 B.n105 585
R169 B.n469 B.n468 585
R170 B.n467 B.n106 585
R171 B.n466 B.n465 585
R172 B.n464 B.n107 585
R173 B.n463 B.n462 585
R174 B.n461 B.n108 585
R175 B.n460 B.n459 585
R176 B.n458 B.n109 585
R177 B.n457 B.n456 585
R178 B.n455 B.n110 585
R179 B.n454 B.n453 585
R180 B.n452 B.n111 585
R181 B.n451 B.n450 585
R182 B.n449 B.n112 585
R183 B.n448 B.n447 585
R184 B.n446 B.n113 585
R185 B.n445 B.n444 585
R186 B.n443 B.n114 585
R187 B.n442 B.n441 585
R188 B.n440 B.n115 585
R189 B.n241 B.n240 585
R190 B.n242 B.n185 585
R191 B.n244 B.n243 585
R192 B.n245 B.n184 585
R193 B.n247 B.n246 585
R194 B.n248 B.n183 585
R195 B.n250 B.n249 585
R196 B.n251 B.n182 585
R197 B.n253 B.n252 585
R198 B.n254 B.n181 585
R199 B.n256 B.n255 585
R200 B.n257 B.n180 585
R201 B.n259 B.n258 585
R202 B.n260 B.n179 585
R203 B.n262 B.n261 585
R204 B.n263 B.n178 585
R205 B.n265 B.n264 585
R206 B.n266 B.n177 585
R207 B.n268 B.n267 585
R208 B.n269 B.n176 585
R209 B.n271 B.n270 585
R210 B.n272 B.n175 585
R211 B.n274 B.n273 585
R212 B.n275 B.n174 585
R213 B.n277 B.n276 585
R214 B.n278 B.n173 585
R215 B.n280 B.n279 585
R216 B.n281 B.n172 585
R217 B.n283 B.n282 585
R218 B.n284 B.n171 585
R219 B.n286 B.n285 585
R220 B.n287 B.n170 585
R221 B.n289 B.n288 585
R222 B.n290 B.n169 585
R223 B.n292 B.n291 585
R224 B.n293 B.n168 585
R225 B.n295 B.n294 585
R226 B.n296 B.n167 585
R227 B.n298 B.n297 585
R228 B.n299 B.n166 585
R229 B.n301 B.n300 585
R230 B.n302 B.n165 585
R231 B.n304 B.n303 585
R232 B.n305 B.n164 585
R233 B.n307 B.n306 585
R234 B.n308 B.n163 585
R235 B.n310 B.n309 585
R236 B.n311 B.n162 585
R237 B.n313 B.n312 585
R238 B.n314 B.n161 585
R239 B.n316 B.n315 585
R240 B.n317 B.n160 585
R241 B.n319 B.n318 585
R242 B.n320 B.n159 585
R243 B.n322 B.n321 585
R244 B.n323 B.n158 585
R245 B.n325 B.n324 585
R246 B.n326 B.n157 585
R247 B.n328 B.n327 585
R248 B.n329 B.n156 585
R249 B.n331 B.n330 585
R250 B.n333 B.n332 585
R251 B.n334 B.n152 585
R252 B.n336 B.n335 585
R253 B.n337 B.n151 585
R254 B.n339 B.n338 585
R255 B.n340 B.n150 585
R256 B.n342 B.n341 585
R257 B.n343 B.n149 585
R258 B.n345 B.n344 585
R259 B.n346 B.n146 585
R260 B.n349 B.n348 585
R261 B.n350 B.n145 585
R262 B.n352 B.n351 585
R263 B.n353 B.n144 585
R264 B.n355 B.n354 585
R265 B.n356 B.n143 585
R266 B.n358 B.n357 585
R267 B.n359 B.n142 585
R268 B.n361 B.n360 585
R269 B.n362 B.n141 585
R270 B.n364 B.n363 585
R271 B.n365 B.n140 585
R272 B.n367 B.n366 585
R273 B.n368 B.n139 585
R274 B.n370 B.n369 585
R275 B.n371 B.n138 585
R276 B.n373 B.n372 585
R277 B.n374 B.n137 585
R278 B.n376 B.n375 585
R279 B.n377 B.n136 585
R280 B.n379 B.n378 585
R281 B.n380 B.n135 585
R282 B.n382 B.n381 585
R283 B.n383 B.n134 585
R284 B.n385 B.n384 585
R285 B.n386 B.n133 585
R286 B.n388 B.n387 585
R287 B.n389 B.n132 585
R288 B.n391 B.n390 585
R289 B.n392 B.n131 585
R290 B.n394 B.n393 585
R291 B.n395 B.n130 585
R292 B.n397 B.n396 585
R293 B.n398 B.n129 585
R294 B.n400 B.n399 585
R295 B.n401 B.n128 585
R296 B.n403 B.n402 585
R297 B.n404 B.n127 585
R298 B.n406 B.n405 585
R299 B.n407 B.n126 585
R300 B.n409 B.n408 585
R301 B.n410 B.n125 585
R302 B.n412 B.n411 585
R303 B.n413 B.n124 585
R304 B.n415 B.n414 585
R305 B.n416 B.n123 585
R306 B.n418 B.n417 585
R307 B.n419 B.n122 585
R308 B.n421 B.n420 585
R309 B.n422 B.n121 585
R310 B.n424 B.n423 585
R311 B.n425 B.n120 585
R312 B.n427 B.n426 585
R313 B.n428 B.n119 585
R314 B.n430 B.n429 585
R315 B.n431 B.n118 585
R316 B.n433 B.n432 585
R317 B.n434 B.n117 585
R318 B.n436 B.n435 585
R319 B.n437 B.n116 585
R320 B.n439 B.n438 585
R321 B.n239 B.n186 585
R322 B.n238 B.n237 585
R323 B.n236 B.n187 585
R324 B.n235 B.n234 585
R325 B.n233 B.n188 585
R326 B.n232 B.n231 585
R327 B.n230 B.n189 585
R328 B.n229 B.n228 585
R329 B.n227 B.n190 585
R330 B.n226 B.n225 585
R331 B.n224 B.n191 585
R332 B.n223 B.n222 585
R333 B.n221 B.n192 585
R334 B.n220 B.n219 585
R335 B.n218 B.n193 585
R336 B.n217 B.n216 585
R337 B.n215 B.n194 585
R338 B.n214 B.n213 585
R339 B.n212 B.n195 585
R340 B.n211 B.n210 585
R341 B.n209 B.n196 585
R342 B.n208 B.n207 585
R343 B.n206 B.n197 585
R344 B.n205 B.n204 585
R345 B.n203 B.n198 585
R346 B.n202 B.n201 585
R347 B.n200 B.n199 585
R348 B.n2 B.n0 585
R349 B.n765 B.n1 585
R350 B.n764 B.n763 585
R351 B.n762 B.n3 585
R352 B.n761 B.n760 585
R353 B.n759 B.n4 585
R354 B.n758 B.n757 585
R355 B.n756 B.n5 585
R356 B.n755 B.n754 585
R357 B.n753 B.n6 585
R358 B.n752 B.n751 585
R359 B.n750 B.n7 585
R360 B.n749 B.n748 585
R361 B.n747 B.n8 585
R362 B.n746 B.n745 585
R363 B.n744 B.n9 585
R364 B.n743 B.n742 585
R365 B.n741 B.n10 585
R366 B.n740 B.n739 585
R367 B.n738 B.n11 585
R368 B.n737 B.n736 585
R369 B.n735 B.n12 585
R370 B.n734 B.n733 585
R371 B.n732 B.n13 585
R372 B.n731 B.n730 585
R373 B.n729 B.n14 585
R374 B.n728 B.n727 585
R375 B.n726 B.n15 585
R376 B.n725 B.n724 585
R377 B.n767 B.n766 585
R378 B.n147 B.t5 540.288
R379 B.n55 B.t7 540.288
R380 B.n153 B.t2 540.288
R381 B.n48 B.t10 540.288
R382 B.n241 B.n186 516.524
R383 B.n724 B.n723 516.524
R384 B.n440 B.n439 516.524
R385 B.n525 B.n524 516.524
R386 B.n148 B.t4 496.846
R387 B.n56 B.t8 496.846
R388 B.n154 B.t1 496.846
R389 B.n49 B.t11 496.846
R390 B.n147 B.t3 443.156
R391 B.n153 B.t0 443.156
R392 B.n48 B.t9 443.156
R393 B.n55 B.t6 443.156
R394 B.n237 B.n186 163.367
R395 B.n237 B.n236 163.367
R396 B.n236 B.n235 163.367
R397 B.n235 B.n188 163.367
R398 B.n231 B.n188 163.367
R399 B.n231 B.n230 163.367
R400 B.n230 B.n229 163.367
R401 B.n229 B.n190 163.367
R402 B.n225 B.n190 163.367
R403 B.n225 B.n224 163.367
R404 B.n224 B.n223 163.367
R405 B.n223 B.n192 163.367
R406 B.n219 B.n192 163.367
R407 B.n219 B.n218 163.367
R408 B.n218 B.n217 163.367
R409 B.n217 B.n194 163.367
R410 B.n213 B.n194 163.367
R411 B.n213 B.n212 163.367
R412 B.n212 B.n211 163.367
R413 B.n211 B.n196 163.367
R414 B.n207 B.n196 163.367
R415 B.n207 B.n206 163.367
R416 B.n206 B.n205 163.367
R417 B.n205 B.n198 163.367
R418 B.n201 B.n198 163.367
R419 B.n201 B.n200 163.367
R420 B.n200 B.n2 163.367
R421 B.n766 B.n2 163.367
R422 B.n766 B.n765 163.367
R423 B.n765 B.n764 163.367
R424 B.n764 B.n3 163.367
R425 B.n760 B.n3 163.367
R426 B.n760 B.n759 163.367
R427 B.n759 B.n758 163.367
R428 B.n758 B.n5 163.367
R429 B.n754 B.n5 163.367
R430 B.n754 B.n753 163.367
R431 B.n753 B.n752 163.367
R432 B.n752 B.n7 163.367
R433 B.n748 B.n7 163.367
R434 B.n748 B.n747 163.367
R435 B.n747 B.n746 163.367
R436 B.n746 B.n9 163.367
R437 B.n742 B.n9 163.367
R438 B.n742 B.n741 163.367
R439 B.n741 B.n740 163.367
R440 B.n740 B.n11 163.367
R441 B.n736 B.n11 163.367
R442 B.n736 B.n735 163.367
R443 B.n735 B.n734 163.367
R444 B.n734 B.n13 163.367
R445 B.n730 B.n13 163.367
R446 B.n730 B.n729 163.367
R447 B.n729 B.n728 163.367
R448 B.n728 B.n15 163.367
R449 B.n724 B.n15 163.367
R450 B.n242 B.n241 163.367
R451 B.n243 B.n242 163.367
R452 B.n243 B.n184 163.367
R453 B.n247 B.n184 163.367
R454 B.n248 B.n247 163.367
R455 B.n249 B.n248 163.367
R456 B.n249 B.n182 163.367
R457 B.n253 B.n182 163.367
R458 B.n254 B.n253 163.367
R459 B.n255 B.n254 163.367
R460 B.n255 B.n180 163.367
R461 B.n259 B.n180 163.367
R462 B.n260 B.n259 163.367
R463 B.n261 B.n260 163.367
R464 B.n261 B.n178 163.367
R465 B.n265 B.n178 163.367
R466 B.n266 B.n265 163.367
R467 B.n267 B.n266 163.367
R468 B.n267 B.n176 163.367
R469 B.n271 B.n176 163.367
R470 B.n272 B.n271 163.367
R471 B.n273 B.n272 163.367
R472 B.n273 B.n174 163.367
R473 B.n277 B.n174 163.367
R474 B.n278 B.n277 163.367
R475 B.n279 B.n278 163.367
R476 B.n279 B.n172 163.367
R477 B.n283 B.n172 163.367
R478 B.n284 B.n283 163.367
R479 B.n285 B.n284 163.367
R480 B.n285 B.n170 163.367
R481 B.n289 B.n170 163.367
R482 B.n290 B.n289 163.367
R483 B.n291 B.n290 163.367
R484 B.n291 B.n168 163.367
R485 B.n295 B.n168 163.367
R486 B.n296 B.n295 163.367
R487 B.n297 B.n296 163.367
R488 B.n297 B.n166 163.367
R489 B.n301 B.n166 163.367
R490 B.n302 B.n301 163.367
R491 B.n303 B.n302 163.367
R492 B.n303 B.n164 163.367
R493 B.n307 B.n164 163.367
R494 B.n308 B.n307 163.367
R495 B.n309 B.n308 163.367
R496 B.n309 B.n162 163.367
R497 B.n313 B.n162 163.367
R498 B.n314 B.n313 163.367
R499 B.n315 B.n314 163.367
R500 B.n315 B.n160 163.367
R501 B.n319 B.n160 163.367
R502 B.n320 B.n319 163.367
R503 B.n321 B.n320 163.367
R504 B.n321 B.n158 163.367
R505 B.n325 B.n158 163.367
R506 B.n326 B.n325 163.367
R507 B.n327 B.n326 163.367
R508 B.n327 B.n156 163.367
R509 B.n331 B.n156 163.367
R510 B.n332 B.n331 163.367
R511 B.n332 B.n152 163.367
R512 B.n336 B.n152 163.367
R513 B.n337 B.n336 163.367
R514 B.n338 B.n337 163.367
R515 B.n338 B.n150 163.367
R516 B.n342 B.n150 163.367
R517 B.n343 B.n342 163.367
R518 B.n344 B.n343 163.367
R519 B.n344 B.n146 163.367
R520 B.n349 B.n146 163.367
R521 B.n350 B.n349 163.367
R522 B.n351 B.n350 163.367
R523 B.n351 B.n144 163.367
R524 B.n355 B.n144 163.367
R525 B.n356 B.n355 163.367
R526 B.n357 B.n356 163.367
R527 B.n357 B.n142 163.367
R528 B.n361 B.n142 163.367
R529 B.n362 B.n361 163.367
R530 B.n363 B.n362 163.367
R531 B.n363 B.n140 163.367
R532 B.n367 B.n140 163.367
R533 B.n368 B.n367 163.367
R534 B.n369 B.n368 163.367
R535 B.n369 B.n138 163.367
R536 B.n373 B.n138 163.367
R537 B.n374 B.n373 163.367
R538 B.n375 B.n374 163.367
R539 B.n375 B.n136 163.367
R540 B.n379 B.n136 163.367
R541 B.n380 B.n379 163.367
R542 B.n381 B.n380 163.367
R543 B.n381 B.n134 163.367
R544 B.n385 B.n134 163.367
R545 B.n386 B.n385 163.367
R546 B.n387 B.n386 163.367
R547 B.n387 B.n132 163.367
R548 B.n391 B.n132 163.367
R549 B.n392 B.n391 163.367
R550 B.n393 B.n392 163.367
R551 B.n393 B.n130 163.367
R552 B.n397 B.n130 163.367
R553 B.n398 B.n397 163.367
R554 B.n399 B.n398 163.367
R555 B.n399 B.n128 163.367
R556 B.n403 B.n128 163.367
R557 B.n404 B.n403 163.367
R558 B.n405 B.n404 163.367
R559 B.n405 B.n126 163.367
R560 B.n409 B.n126 163.367
R561 B.n410 B.n409 163.367
R562 B.n411 B.n410 163.367
R563 B.n411 B.n124 163.367
R564 B.n415 B.n124 163.367
R565 B.n416 B.n415 163.367
R566 B.n417 B.n416 163.367
R567 B.n417 B.n122 163.367
R568 B.n421 B.n122 163.367
R569 B.n422 B.n421 163.367
R570 B.n423 B.n422 163.367
R571 B.n423 B.n120 163.367
R572 B.n427 B.n120 163.367
R573 B.n428 B.n427 163.367
R574 B.n429 B.n428 163.367
R575 B.n429 B.n118 163.367
R576 B.n433 B.n118 163.367
R577 B.n434 B.n433 163.367
R578 B.n435 B.n434 163.367
R579 B.n435 B.n116 163.367
R580 B.n439 B.n116 163.367
R581 B.n441 B.n440 163.367
R582 B.n441 B.n114 163.367
R583 B.n445 B.n114 163.367
R584 B.n446 B.n445 163.367
R585 B.n447 B.n446 163.367
R586 B.n447 B.n112 163.367
R587 B.n451 B.n112 163.367
R588 B.n452 B.n451 163.367
R589 B.n453 B.n452 163.367
R590 B.n453 B.n110 163.367
R591 B.n457 B.n110 163.367
R592 B.n458 B.n457 163.367
R593 B.n459 B.n458 163.367
R594 B.n459 B.n108 163.367
R595 B.n463 B.n108 163.367
R596 B.n464 B.n463 163.367
R597 B.n465 B.n464 163.367
R598 B.n465 B.n106 163.367
R599 B.n469 B.n106 163.367
R600 B.n470 B.n469 163.367
R601 B.n471 B.n470 163.367
R602 B.n471 B.n104 163.367
R603 B.n475 B.n104 163.367
R604 B.n476 B.n475 163.367
R605 B.n477 B.n476 163.367
R606 B.n477 B.n102 163.367
R607 B.n481 B.n102 163.367
R608 B.n482 B.n481 163.367
R609 B.n483 B.n482 163.367
R610 B.n483 B.n100 163.367
R611 B.n487 B.n100 163.367
R612 B.n488 B.n487 163.367
R613 B.n489 B.n488 163.367
R614 B.n489 B.n98 163.367
R615 B.n493 B.n98 163.367
R616 B.n494 B.n493 163.367
R617 B.n495 B.n494 163.367
R618 B.n495 B.n96 163.367
R619 B.n499 B.n96 163.367
R620 B.n500 B.n499 163.367
R621 B.n501 B.n500 163.367
R622 B.n501 B.n94 163.367
R623 B.n505 B.n94 163.367
R624 B.n506 B.n505 163.367
R625 B.n507 B.n506 163.367
R626 B.n507 B.n92 163.367
R627 B.n511 B.n92 163.367
R628 B.n512 B.n511 163.367
R629 B.n513 B.n512 163.367
R630 B.n513 B.n90 163.367
R631 B.n517 B.n90 163.367
R632 B.n518 B.n517 163.367
R633 B.n519 B.n518 163.367
R634 B.n519 B.n88 163.367
R635 B.n523 B.n88 163.367
R636 B.n524 B.n523 163.367
R637 B.n723 B.n722 163.367
R638 B.n722 B.n17 163.367
R639 B.n718 B.n17 163.367
R640 B.n718 B.n717 163.367
R641 B.n717 B.n716 163.367
R642 B.n716 B.n19 163.367
R643 B.n712 B.n19 163.367
R644 B.n712 B.n711 163.367
R645 B.n711 B.n710 163.367
R646 B.n710 B.n21 163.367
R647 B.n706 B.n21 163.367
R648 B.n706 B.n705 163.367
R649 B.n705 B.n704 163.367
R650 B.n704 B.n23 163.367
R651 B.n700 B.n23 163.367
R652 B.n700 B.n699 163.367
R653 B.n699 B.n698 163.367
R654 B.n698 B.n25 163.367
R655 B.n694 B.n25 163.367
R656 B.n694 B.n693 163.367
R657 B.n693 B.n692 163.367
R658 B.n692 B.n27 163.367
R659 B.n688 B.n27 163.367
R660 B.n688 B.n687 163.367
R661 B.n687 B.n686 163.367
R662 B.n686 B.n29 163.367
R663 B.n682 B.n29 163.367
R664 B.n682 B.n681 163.367
R665 B.n681 B.n680 163.367
R666 B.n680 B.n31 163.367
R667 B.n676 B.n31 163.367
R668 B.n676 B.n675 163.367
R669 B.n675 B.n674 163.367
R670 B.n674 B.n33 163.367
R671 B.n670 B.n33 163.367
R672 B.n670 B.n669 163.367
R673 B.n669 B.n668 163.367
R674 B.n668 B.n35 163.367
R675 B.n664 B.n35 163.367
R676 B.n664 B.n663 163.367
R677 B.n663 B.n662 163.367
R678 B.n662 B.n37 163.367
R679 B.n658 B.n37 163.367
R680 B.n658 B.n657 163.367
R681 B.n657 B.n656 163.367
R682 B.n656 B.n39 163.367
R683 B.n652 B.n39 163.367
R684 B.n652 B.n651 163.367
R685 B.n651 B.n650 163.367
R686 B.n650 B.n41 163.367
R687 B.n646 B.n41 163.367
R688 B.n646 B.n645 163.367
R689 B.n645 B.n644 163.367
R690 B.n644 B.n43 163.367
R691 B.n640 B.n43 163.367
R692 B.n640 B.n639 163.367
R693 B.n639 B.n638 163.367
R694 B.n638 B.n45 163.367
R695 B.n634 B.n45 163.367
R696 B.n634 B.n633 163.367
R697 B.n633 B.n632 163.367
R698 B.n632 B.n47 163.367
R699 B.n628 B.n47 163.367
R700 B.n628 B.n627 163.367
R701 B.n627 B.n626 163.367
R702 B.n626 B.n52 163.367
R703 B.n622 B.n52 163.367
R704 B.n622 B.n621 163.367
R705 B.n621 B.n620 163.367
R706 B.n620 B.n54 163.367
R707 B.n615 B.n54 163.367
R708 B.n615 B.n614 163.367
R709 B.n614 B.n613 163.367
R710 B.n613 B.n58 163.367
R711 B.n609 B.n58 163.367
R712 B.n609 B.n608 163.367
R713 B.n608 B.n607 163.367
R714 B.n607 B.n60 163.367
R715 B.n603 B.n60 163.367
R716 B.n603 B.n602 163.367
R717 B.n602 B.n601 163.367
R718 B.n601 B.n62 163.367
R719 B.n597 B.n62 163.367
R720 B.n597 B.n596 163.367
R721 B.n596 B.n595 163.367
R722 B.n595 B.n64 163.367
R723 B.n591 B.n64 163.367
R724 B.n591 B.n590 163.367
R725 B.n590 B.n589 163.367
R726 B.n589 B.n66 163.367
R727 B.n585 B.n66 163.367
R728 B.n585 B.n584 163.367
R729 B.n584 B.n583 163.367
R730 B.n583 B.n68 163.367
R731 B.n579 B.n68 163.367
R732 B.n579 B.n578 163.367
R733 B.n578 B.n577 163.367
R734 B.n577 B.n70 163.367
R735 B.n573 B.n70 163.367
R736 B.n573 B.n572 163.367
R737 B.n572 B.n571 163.367
R738 B.n571 B.n72 163.367
R739 B.n567 B.n72 163.367
R740 B.n567 B.n566 163.367
R741 B.n566 B.n565 163.367
R742 B.n565 B.n74 163.367
R743 B.n561 B.n74 163.367
R744 B.n561 B.n560 163.367
R745 B.n560 B.n559 163.367
R746 B.n559 B.n76 163.367
R747 B.n555 B.n76 163.367
R748 B.n555 B.n554 163.367
R749 B.n554 B.n553 163.367
R750 B.n553 B.n78 163.367
R751 B.n549 B.n78 163.367
R752 B.n549 B.n548 163.367
R753 B.n548 B.n547 163.367
R754 B.n547 B.n80 163.367
R755 B.n543 B.n80 163.367
R756 B.n543 B.n542 163.367
R757 B.n542 B.n541 163.367
R758 B.n541 B.n82 163.367
R759 B.n537 B.n82 163.367
R760 B.n537 B.n536 163.367
R761 B.n536 B.n535 163.367
R762 B.n535 B.n84 163.367
R763 B.n531 B.n84 163.367
R764 B.n531 B.n530 163.367
R765 B.n530 B.n529 163.367
R766 B.n529 B.n86 163.367
R767 B.n525 B.n86 163.367
R768 B.n347 B.n148 59.5399
R769 B.n155 B.n154 59.5399
R770 B.n50 B.n49 59.5399
R771 B.n617 B.n56 59.5399
R772 B.n148 B.n147 43.4429
R773 B.n154 B.n153 43.4429
R774 B.n49 B.n48 43.4429
R775 B.n56 B.n55 43.4429
R776 B.n725 B.n16 33.5615
R777 B.n526 B.n87 33.5615
R778 B.n438 B.n115 33.5615
R779 B.n240 B.n239 33.5615
R780 B B.n767 18.0485
R781 B.n721 B.n16 10.6151
R782 B.n721 B.n720 10.6151
R783 B.n720 B.n719 10.6151
R784 B.n719 B.n18 10.6151
R785 B.n715 B.n18 10.6151
R786 B.n715 B.n714 10.6151
R787 B.n714 B.n713 10.6151
R788 B.n713 B.n20 10.6151
R789 B.n709 B.n20 10.6151
R790 B.n709 B.n708 10.6151
R791 B.n708 B.n707 10.6151
R792 B.n707 B.n22 10.6151
R793 B.n703 B.n22 10.6151
R794 B.n703 B.n702 10.6151
R795 B.n702 B.n701 10.6151
R796 B.n701 B.n24 10.6151
R797 B.n697 B.n24 10.6151
R798 B.n697 B.n696 10.6151
R799 B.n696 B.n695 10.6151
R800 B.n695 B.n26 10.6151
R801 B.n691 B.n26 10.6151
R802 B.n691 B.n690 10.6151
R803 B.n690 B.n689 10.6151
R804 B.n689 B.n28 10.6151
R805 B.n685 B.n28 10.6151
R806 B.n685 B.n684 10.6151
R807 B.n684 B.n683 10.6151
R808 B.n683 B.n30 10.6151
R809 B.n679 B.n30 10.6151
R810 B.n679 B.n678 10.6151
R811 B.n678 B.n677 10.6151
R812 B.n677 B.n32 10.6151
R813 B.n673 B.n32 10.6151
R814 B.n673 B.n672 10.6151
R815 B.n672 B.n671 10.6151
R816 B.n671 B.n34 10.6151
R817 B.n667 B.n34 10.6151
R818 B.n667 B.n666 10.6151
R819 B.n666 B.n665 10.6151
R820 B.n665 B.n36 10.6151
R821 B.n661 B.n36 10.6151
R822 B.n661 B.n660 10.6151
R823 B.n660 B.n659 10.6151
R824 B.n659 B.n38 10.6151
R825 B.n655 B.n38 10.6151
R826 B.n655 B.n654 10.6151
R827 B.n654 B.n653 10.6151
R828 B.n653 B.n40 10.6151
R829 B.n649 B.n40 10.6151
R830 B.n649 B.n648 10.6151
R831 B.n648 B.n647 10.6151
R832 B.n647 B.n42 10.6151
R833 B.n643 B.n42 10.6151
R834 B.n643 B.n642 10.6151
R835 B.n642 B.n641 10.6151
R836 B.n641 B.n44 10.6151
R837 B.n637 B.n44 10.6151
R838 B.n637 B.n636 10.6151
R839 B.n636 B.n635 10.6151
R840 B.n635 B.n46 10.6151
R841 B.n631 B.n630 10.6151
R842 B.n630 B.n629 10.6151
R843 B.n629 B.n51 10.6151
R844 B.n625 B.n51 10.6151
R845 B.n625 B.n624 10.6151
R846 B.n624 B.n623 10.6151
R847 B.n623 B.n53 10.6151
R848 B.n619 B.n53 10.6151
R849 B.n619 B.n618 10.6151
R850 B.n616 B.n57 10.6151
R851 B.n612 B.n57 10.6151
R852 B.n612 B.n611 10.6151
R853 B.n611 B.n610 10.6151
R854 B.n610 B.n59 10.6151
R855 B.n606 B.n59 10.6151
R856 B.n606 B.n605 10.6151
R857 B.n605 B.n604 10.6151
R858 B.n604 B.n61 10.6151
R859 B.n600 B.n61 10.6151
R860 B.n600 B.n599 10.6151
R861 B.n599 B.n598 10.6151
R862 B.n598 B.n63 10.6151
R863 B.n594 B.n63 10.6151
R864 B.n594 B.n593 10.6151
R865 B.n593 B.n592 10.6151
R866 B.n592 B.n65 10.6151
R867 B.n588 B.n65 10.6151
R868 B.n588 B.n587 10.6151
R869 B.n587 B.n586 10.6151
R870 B.n586 B.n67 10.6151
R871 B.n582 B.n67 10.6151
R872 B.n582 B.n581 10.6151
R873 B.n581 B.n580 10.6151
R874 B.n580 B.n69 10.6151
R875 B.n576 B.n69 10.6151
R876 B.n576 B.n575 10.6151
R877 B.n575 B.n574 10.6151
R878 B.n574 B.n71 10.6151
R879 B.n570 B.n71 10.6151
R880 B.n570 B.n569 10.6151
R881 B.n569 B.n568 10.6151
R882 B.n568 B.n73 10.6151
R883 B.n564 B.n73 10.6151
R884 B.n564 B.n563 10.6151
R885 B.n563 B.n562 10.6151
R886 B.n562 B.n75 10.6151
R887 B.n558 B.n75 10.6151
R888 B.n558 B.n557 10.6151
R889 B.n557 B.n556 10.6151
R890 B.n556 B.n77 10.6151
R891 B.n552 B.n77 10.6151
R892 B.n552 B.n551 10.6151
R893 B.n551 B.n550 10.6151
R894 B.n550 B.n79 10.6151
R895 B.n546 B.n79 10.6151
R896 B.n546 B.n545 10.6151
R897 B.n545 B.n544 10.6151
R898 B.n544 B.n81 10.6151
R899 B.n540 B.n81 10.6151
R900 B.n540 B.n539 10.6151
R901 B.n539 B.n538 10.6151
R902 B.n538 B.n83 10.6151
R903 B.n534 B.n83 10.6151
R904 B.n534 B.n533 10.6151
R905 B.n533 B.n532 10.6151
R906 B.n532 B.n85 10.6151
R907 B.n528 B.n85 10.6151
R908 B.n528 B.n527 10.6151
R909 B.n527 B.n526 10.6151
R910 B.n442 B.n115 10.6151
R911 B.n443 B.n442 10.6151
R912 B.n444 B.n443 10.6151
R913 B.n444 B.n113 10.6151
R914 B.n448 B.n113 10.6151
R915 B.n449 B.n448 10.6151
R916 B.n450 B.n449 10.6151
R917 B.n450 B.n111 10.6151
R918 B.n454 B.n111 10.6151
R919 B.n455 B.n454 10.6151
R920 B.n456 B.n455 10.6151
R921 B.n456 B.n109 10.6151
R922 B.n460 B.n109 10.6151
R923 B.n461 B.n460 10.6151
R924 B.n462 B.n461 10.6151
R925 B.n462 B.n107 10.6151
R926 B.n466 B.n107 10.6151
R927 B.n467 B.n466 10.6151
R928 B.n468 B.n467 10.6151
R929 B.n468 B.n105 10.6151
R930 B.n472 B.n105 10.6151
R931 B.n473 B.n472 10.6151
R932 B.n474 B.n473 10.6151
R933 B.n474 B.n103 10.6151
R934 B.n478 B.n103 10.6151
R935 B.n479 B.n478 10.6151
R936 B.n480 B.n479 10.6151
R937 B.n480 B.n101 10.6151
R938 B.n484 B.n101 10.6151
R939 B.n485 B.n484 10.6151
R940 B.n486 B.n485 10.6151
R941 B.n486 B.n99 10.6151
R942 B.n490 B.n99 10.6151
R943 B.n491 B.n490 10.6151
R944 B.n492 B.n491 10.6151
R945 B.n492 B.n97 10.6151
R946 B.n496 B.n97 10.6151
R947 B.n497 B.n496 10.6151
R948 B.n498 B.n497 10.6151
R949 B.n498 B.n95 10.6151
R950 B.n502 B.n95 10.6151
R951 B.n503 B.n502 10.6151
R952 B.n504 B.n503 10.6151
R953 B.n504 B.n93 10.6151
R954 B.n508 B.n93 10.6151
R955 B.n509 B.n508 10.6151
R956 B.n510 B.n509 10.6151
R957 B.n510 B.n91 10.6151
R958 B.n514 B.n91 10.6151
R959 B.n515 B.n514 10.6151
R960 B.n516 B.n515 10.6151
R961 B.n516 B.n89 10.6151
R962 B.n520 B.n89 10.6151
R963 B.n521 B.n520 10.6151
R964 B.n522 B.n521 10.6151
R965 B.n522 B.n87 10.6151
R966 B.n240 B.n185 10.6151
R967 B.n244 B.n185 10.6151
R968 B.n245 B.n244 10.6151
R969 B.n246 B.n245 10.6151
R970 B.n246 B.n183 10.6151
R971 B.n250 B.n183 10.6151
R972 B.n251 B.n250 10.6151
R973 B.n252 B.n251 10.6151
R974 B.n252 B.n181 10.6151
R975 B.n256 B.n181 10.6151
R976 B.n257 B.n256 10.6151
R977 B.n258 B.n257 10.6151
R978 B.n258 B.n179 10.6151
R979 B.n262 B.n179 10.6151
R980 B.n263 B.n262 10.6151
R981 B.n264 B.n263 10.6151
R982 B.n264 B.n177 10.6151
R983 B.n268 B.n177 10.6151
R984 B.n269 B.n268 10.6151
R985 B.n270 B.n269 10.6151
R986 B.n270 B.n175 10.6151
R987 B.n274 B.n175 10.6151
R988 B.n275 B.n274 10.6151
R989 B.n276 B.n275 10.6151
R990 B.n276 B.n173 10.6151
R991 B.n280 B.n173 10.6151
R992 B.n281 B.n280 10.6151
R993 B.n282 B.n281 10.6151
R994 B.n282 B.n171 10.6151
R995 B.n286 B.n171 10.6151
R996 B.n287 B.n286 10.6151
R997 B.n288 B.n287 10.6151
R998 B.n288 B.n169 10.6151
R999 B.n292 B.n169 10.6151
R1000 B.n293 B.n292 10.6151
R1001 B.n294 B.n293 10.6151
R1002 B.n294 B.n167 10.6151
R1003 B.n298 B.n167 10.6151
R1004 B.n299 B.n298 10.6151
R1005 B.n300 B.n299 10.6151
R1006 B.n300 B.n165 10.6151
R1007 B.n304 B.n165 10.6151
R1008 B.n305 B.n304 10.6151
R1009 B.n306 B.n305 10.6151
R1010 B.n306 B.n163 10.6151
R1011 B.n310 B.n163 10.6151
R1012 B.n311 B.n310 10.6151
R1013 B.n312 B.n311 10.6151
R1014 B.n312 B.n161 10.6151
R1015 B.n316 B.n161 10.6151
R1016 B.n317 B.n316 10.6151
R1017 B.n318 B.n317 10.6151
R1018 B.n318 B.n159 10.6151
R1019 B.n322 B.n159 10.6151
R1020 B.n323 B.n322 10.6151
R1021 B.n324 B.n323 10.6151
R1022 B.n324 B.n157 10.6151
R1023 B.n328 B.n157 10.6151
R1024 B.n329 B.n328 10.6151
R1025 B.n330 B.n329 10.6151
R1026 B.n334 B.n333 10.6151
R1027 B.n335 B.n334 10.6151
R1028 B.n335 B.n151 10.6151
R1029 B.n339 B.n151 10.6151
R1030 B.n340 B.n339 10.6151
R1031 B.n341 B.n340 10.6151
R1032 B.n341 B.n149 10.6151
R1033 B.n345 B.n149 10.6151
R1034 B.n346 B.n345 10.6151
R1035 B.n348 B.n145 10.6151
R1036 B.n352 B.n145 10.6151
R1037 B.n353 B.n352 10.6151
R1038 B.n354 B.n353 10.6151
R1039 B.n354 B.n143 10.6151
R1040 B.n358 B.n143 10.6151
R1041 B.n359 B.n358 10.6151
R1042 B.n360 B.n359 10.6151
R1043 B.n360 B.n141 10.6151
R1044 B.n364 B.n141 10.6151
R1045 B.n365 B.n364 10.6151
R1046 B.n366 B.n365 10.6151
R1047 B.n366 B.n139 10.6151
R1048 B.n370 B.n139 10.6151
R1049 B.n371 B.n370 10.6151
R1050 B.n372 B.n371 10.6151
R1051 B.n372 B.n137 10.6151
R1052 B.n376 B.n137 10.6151
R1053 B.n377 B.n376 10.6151
R1054 B.n378 B.n377 10.6151
R1055 B.n378 B.n135 10.6151
R1056 B.n382 B.n135 10.6151
R1057 B.n383 B.n382 10.6151
R1058 B.n384 B.n383 10.6151
R1059 B.n384 B.n133 10.6151
R1060 B.n388 B.n133 10.6151
R1061 B.n389 B.n388 10.6151
R1062 B.n390 B.n389 10.6151
R1063 B.n390 B.n131 10.6151
R1064 B.n394 B.n131 10.6151
R1065 B.n395 B.n394 10.6151
R1066 B.n396 B.n395 10.6151
R1067 B.n396 B.n129 10.6151
R1068 B.n400 B.n129 10.6151
R1069 B.n401 B.n400 10.6151
R1070 B.n402 B.n401 10.6151
R1071 B.n402 B.n127 10.6151
R1072 B.n406 B.n127 10.6151
R1073 B.n407 B.n406 10.6151
R1074 B.n408 B.n407 10.6151
R1075 B.n408 B.n125 10.6151
R1076 B.n412 B.n125 10.6151
R1077 B.n413 B.n412 10.6151
R1078 B.n414 B.n413 10.6151
R1079 B.n414 B.n123 10.6151
R1080 B.n418 B.n123 10.6151
R1081 B.n419 B.n418 10.6151
R1082 B.n420 B.n419 10.6151
R1083 B.n420 B.n121 10.6151
R1084 B.n424 B.n121 10.6151
R1085 B.n425 B.n424 10.6151
R1086 B.n426 B.n425 10.6151
R1087 B.n426 B.n119 10.6151
R1088 B.n430 B.n119 10.6151
R1089 B.n431 B.n430 10.6151
R1090 B.n432 B.n431 10.6151
R1091 B.n432 B.n117 10.6151
R1092 B.n436 B.n117 10.6151
R1093 B.n437 B.n436 10.6151
R1094 B.n438 B.n437 10.6151
R1095 B.n239 B.n238 10.6151
R1096 B.n238 B.n187 10.6151
R1097 B.n234 B.n187 10.6151
R1098 B.n234 B.n233 10.6151
R1099 B.n233 B.n232 10.6151
R1100 B.n232 B.n189 10.6151
R1101 B.n228 B.n189 10.6151
R1102 B.n228 B.n227 10.6151
R1103 B.n227 B.n226 10.6151
R1104 B.n226 B.n191 10.6151
R1105 B.n222 B.n191 10.6151
R1106 B.n222 B.n221 10.6151
R1107 B.n221 B.n220 10.6151
R1108 B.n220 B.n193 10.6151
R1109 B.n216 B.n193 10.6151
R1110 B.n216 B.n215 10.6151
R1111 B.n215 B.n214 10.6151
R1112 B.n214 B.n195 10.6151
R1113 B.n210 B.n195 10.6151
R1114 B.n210 B.n209 10.6151
R1115 B.n209 B.n208 10.6151
R1116 B.n208 B.n197 10.6151
R1117 B.n204 B.n197 10.6151
R1118 B.n204 B.n203 10.6151
R1119 B.n203 B.n202 10.6151
R1120 B.n202 B.n199 10.6151
R1121 B.n199 B.n0 10.6151
R1122 B.n763 B.n1 10.6151
R1123 B.n763 B.n762 10.6151
R1124 B.n762 B.n761 10.6151
R1125 B.n761 B.n4 10.6151
R1126 B.n757 B.n4 10.6151
R1127 B.n757 B.n756 10.6151
R1128 B.n756 B.n755 10.6151
R1129 B.n755 B.n6 10.6151
R1130 B.n751 B.n6 10.6151
R1131 B.n751 B.n750 10.6151
R1132 B.n750 B.n749 10.6151
R1133 B.n749 B.n8 10.6151
R1134 B.n745 B.n8 10.6151
R1135 B.n745 B.n744 10.6151
R1136 B.n744 B.n743 10.6151
R1137 B.n743 B.n10 10.6151
R1138 B.n739 B.n10 10.6151
R1139 B.n739 B.n738 10.6151
R1140 B.n738 B.n737 10.6151
R1141 B.n737 B.n12 10.6151
R1142 B.n733 B.n12 10.6151
R1143 B.n733 B.n732 10.6151
R1144 B.n732 B.n731 10.6151
R1145 B.n731 B.n14 10.6151
R1146 B.n727 B.n14 10.6151
R1147 B.n727 B.n726 10.6151
R1148 B.n726 B.n725 10.6151
R1149 B.n50 B.n46 9.36635
R1150 B.n617 B.n616 9.36635
R1151 B.n330 B.n155 9.36635
R1152 B.n348 B.n347 9.36635
R1153 B.n767 B.n0 2.81026
R1154 B.n767 B.n1 2.81026
R1155 B.n631 B.n50 1.24928
R1156 B.n618 B.n617 1.24928
R1157 B.n333 B.n155 1.24928
R1158 B.n347 B.n346 1.24928
R1159 VN.n0 VN.t0 271.589
R1160 VN.n1 VN.t2 271.589
R1161 VN.n0 VN.t1 271.07
R1162 VN.n1 VN.t3 271.07
R1163 VN VN.n1 57.0854
R1164 VN VN.n0 7.60439
R1165 VDD2.n2 VDD2.n0 116.465
R1166 VDD2.n2 VDD2.n1 70.8013
R1167 VDD2.n1 VDD2.t3 1.73502
R1168 VDD2.n1 VDD2.t1 1.73502
R1169 VDD2.n0 VDD2.t0 1.73502
R1170 VDD2.n0 VDD2.t2 1.73502
R1171 VDD2 VDD2.n2 0.0586897
R1172 VTAIL.n830 VTAIL.n829 756.745
R1173 VTAIL.n102 VTAIL.n101 756.745
R1174 VTAIL.n206 VTAIL.n205 756.745
R1175 VTAIL.n310 VTAIL.n309 756.745
R1176 VTAIL.n726 VTAIL.n725 756.745
R1177 VTAIL.n622 VTAIL.n621 756.745
R1178 VTAIL.n518 VTAIL.n517 756.745
R1179 VTAIL.n414 VTAIL.n413 756.745
R1180 VTAIL.n763 VTAIL.n762 585
R1181 VTAIL.n765 VTAIL.n764 585
R1182 VTAIL.n758 VTAIL.n757 585
R1183 VTAIL.n771 VTAIL.n770 585
R1184 VTAIL.n773 VTAIL.n772 585
R1185 VTAIL.n754 VTAIL.n753 585
R1186 VTAIL.n780 VTAIL.n779 585
R1187 VTAIL.n781 VTAIL.n752 585
R1188 VTAIL.n783 VTAIL.n782 585
R1189 VTAIL.n750 VTAIL.n749 585
R1190 VTAIL.n789 VTAIL.n788 585
R1191 VTAIL.n791 VTAIL.n790 585
R1192 VTAIL.n746 VTAIL.n745 585
R1193 VTAIL.n797 VTAIL.n796 585
R1194 VTAIL.n799 VTAIL.n798 585
R1195 VTAIL.n742 VTAIL.n741 585
R1196 VTAIL.n805 VTAIL.n804 585
R1197 VTAIL.n807 VTAIL.n806 585
R1198 VTAIL.n738 VTAIL.n737 585
R1199 VTAIL.n813 VTAIL.n812 585
R1200 VTAIL.n815 VTAIL.n814 585
R1201 VTAIL.n734 VTAIL.n733 585
R1202 VTAIL.n821 VTAIL.n820 585
R1203 VTAIL.n823 VTAIL.n822 585
R1204 VTAIL.n730 VTAIL.n729 585
R1205 VTAIL.n829 VTAIL.n828 585
R1206 VTAIL.n35 VTAIL.n34 585
R1207 VTAIL.n37 VTAIL.n36 585
R1208 VTAIL.n30 VTAIL.n29 585
R1209 VTAIL.n43 VTAIL.n42 585
R1210 VTAIL.n45 VTAIL.n44 585
R1211 VTAIL.n26 VTAIL.n25 585
R1212 VTAIL.n52 VTAIL.n51 585
R1213 VTAIL.n53 VTAIL.n24 585
R1214 VTAIL.n55 VTAIL.n54 585
R1215 VTAIL.n22 VTAIL.n21 585
R1216 VTAIL.n61 VTAIL.n60 585
R1217 VTAIL.n63 VTAIL.n62 585
R1218 VTAIL.n18 VTAIL.n17 585
R1219 VTAIL.n69 VTAIL.n68 585
R1220 VTAIL.n71 VTAIL.n70 585
R1221 VTAIL.n14 VTAIL.n13 585
R1222 VTAIL.n77 VTAIL.n76 585
R1223 VTAIL.n79 VTAIL.n78 585
R1224 VTAIL.n10 VTAIL.n9 585
R1225 VTAIL.n85 VTAIL.n84 585
R1226 VTAIL.n87 VTAIL.n86 585
R1227 VTAIL.n6 VTAIL.n5 585
R1228 VTAIL.n93 VTAIL.n92 585
R1229 VTAIL.n95 VTAIL.n94 585
R1230 VTAIL.n2 VTAIL.n1 585
R1231 VTAIL.n101 VTAIL.n100 585
R1232 VTAIL.n139 VTAIL.n138 585
R1233 VTAIL.n141 VTAIL.n140 585
R1234 VTAIL.n134 VTAIL.n133 585
R1235 VTAIL.n147 VTAIL.n146 585
R1236 VTAIL.n149 VTAIL.n148 585
R1237 VTAIL.n130 VTAIL.n129 585
R1238 VTAIL.n156 VTAIL.n155 585
R1239 VTAIL.n157 VTAIL.n128 585
R1240 VTAIL.n159 VTAIL.n158 585
R1241 VTAIL.n126 VTAIL.n125 585
R1242 VTAIL.n165 VTAIL.n164 585
R1243 VTAIL.n167 VTAIL.n166 585
R1244 VTAIL.n122 VTAIL.n121 585
R1245 VTAIL.n173 VTAIL.n172 585
R1246 VTAIL.n175 VTAIL.n174 585
R1247 VTAIL.n118 VTAIL.n117 585
R1248 VTAIL.n181 VTAIL.n180 585
R1249 VTAIL.n183 VTAIL.n182 585
R1250 VTAIL.n114 VTAIL.n113 585
R1251 VTAIL.n189 VTAIL.n188 585
R1252 VTAIL.n191 VTAIL.n190 585
R1253 VTAIL.n110 VTAIL.n109 585
R1254 VTAIL.n197 VTAIL.n196 585
R1255 VTAIL.n199 VTAIL.n198 585
R1256 VTAIL.n106 VTAIL.n105 585
R1257 VTAIL.n205 VTAIL.n204 585
R1258 VTAIL.n243 VTAIL.n242 585
R1259 VTAIL.n245 VTAIL.n244 585
R1260 VTAIL.n238 VTAIL.n237 585
R1261 VTAIL.n251 VTAIL.n250 585
R1262 VTAIL.n253 VTAIL.n252 585
R1263 VTAIL.n234 VTAIL.n233 585
R1264 VTAIL.n260 VTAIL.n259 585
R1265 VTAIL.n261 VTAIL.n232 585
R1266 VTAIL.n263 VTAIL.n262 585
R1267 VTAIL.n230 VTAIL.n229 585
R1268 VTAIL.n269 VTAIL.n268 585
R1269 VTAIL.n271 VTAIL.n270 585
R1270 VTAIL.n226 VTAIL.n225 585
R1271 VTAIL.n277 VTAIL.n276 585
R1272 VTAIL.n279 VTAIL.n278 585
R1273 VTAIL.n222 VTAIL.n221 585
R1274 VTAIL.n285 VTAIL.n284 585
R1275 VTAIL.n287 VTAIL.n286 585
R1276 VTAIL.n218 VTAIL.n217 585
R1277 VTAIL.n293 VTAIL.n292 585
R1278 VTAIL.n295 VTAIL.n294 585
R1279 VTAIL.n214 VTAIL.n213 585
R1280 VTAIL.n301 VTAIL.n300 585
R1281 VTAIL.n303 VTAIL.n302 585
R1282 VTAIL.n210 VTAIL.n209 585
R1283 VTAIL.n309 VTAIL.n308 585
R1284 VTAIL.n725 VTAIL.n724 585
R1285 VTAIL.n626 VTAIL.n625 585
R1286 VTAIL.n719 VTAIL.n718 585
R1287 VTAIL.n717 VTAIL.n716 585
R1288 VTAIL.n630 VTAIL.n629 585
R1289 VTAIL.n711 VTAIL.n710 585
R1290 VTAIL.n709 VTAIL.n708 585
R1291 VTAIL.n634 VTAIL.n633 585
R1292 VTAIL.n703 VTAIL.n702 585
R1293 VTAIL.n701 VTAIL.n700 585
R1294 VTAIL.n638 VTAIL.n637 585
R1295 VTAIL.n695 VTAIL.n694 585
R1296 VTAIL.n693 VTAIL.n692 585
R1297 VTAIL.n642 VTAIL.n641 585
R1298 VTAIL.n687 VTAIL.n686 585
R1299 VTAIL.n685 VTAIL.n684 585
R1300 VTAIL.n646 VTAIL.n645 585
R1301 VTAIL.n650 VTAIL.n648 585
R1302 VTAIL.n679 VTAIL.n678 585
R1303 VTAIL.n677 VTAIL.n676 585
R1304 VTAIL.n652 VTAIL.n651 585
R1305 VTAIL.n671 VTAIL.n670 585
R1306 VTAIL.n669 VTAIL.n668 585
R1307 VTAIL.n656 VTAIL.n655 585
R1308 VTAIL.n663 VTAIL.n662 585
R1309 VTAIL.n661 VTAIL.n660 585
R1310 VTAIL.n621 VTAIL.n620 585
R1311 VTAIL.n522 VTAIL.n521 585
R1312 VTAIL.n615 VTAIL.n614 585
R1313 VTAIL.n613 VTAIL.n612 585
R1314 VTAIL.n526 VTAIL.n525 585
R1315 VTAIL.n607 VTAIL.n606 585
R1316 VTAIL.n605 VTAIL.n604 585
R1317 VTAIL.n530 VTAIL.n529 585
R1318 VTAIL.n599 VTAIL.n598 585
R1319 VTAIL.n597 VTAIL.n596 585
R1320 VTAIL.n534 VTAIL.n533 585
R1321 VTAIL.n591 VTAIL.n590 585
R1322 VTAIL.n589 VTAIL.n588 585
R1323 VTAIL.n538 VTAIL.n537 585
R1324 VTAIL.n583 VTAIL.n582 585
R1325 VTAIL.n581 VTAIL.n580 585
R1326 VTAIL.n542 VTAIL.n541 585
R1327 VTAIL.n546 VTAIL.n544 585
R1328 VTAIL.n575 VTAIL.n574 585
R1329 VTAIL.n573 VTAIL.n572 585
R1330 VTAIL.n548 VTAIL.n547 585
R1331 VTAIL.n567 VTAIL.n566 585
R1332 VTAIL.n565 VTAIL.n564 585
R1333 VTAIL.n552 VTAIL.n551 585
R1334 VTAIL.n559 VTAIL.n558 585
R1335 VTAIL.n557 VTAIL.n556 585
R1336 VTAIL.n517 VTAIL.n516 585
R1337 VTAIL.n418 VTAIL.n417 585
R1338 VTAIL.n511 VTAIL.n510 585
R1339 VTAIL.n509 VTAIL.n508 585
R1340 VTAIL.n422 VTAIL.n421 585
R1341 VTAIL.n503 VTAIL.n502 585
R1342 VTAIL.n501 VTAIL.n500 585
R1343 VTAIL.n426 VTAIL.n425 585
R1344 VTAIL.n495 VTAIL.n494 585
R1345 VTAIL.n493 VTAIL.n492 585
R1346 VTAIL.n430 VTAIL.n429 585
R1347 VTAIL.n487 VTAIL.n486 585
R1348 VTAIL.n485 VTAIL.n484 585
R1349 VTAIL.n434 VTAIL.n433 585
R1350 VTAIL.n479 VTAIL.n478 585
R1351 VTAIL.n477 VTAIL.n476 585
R1352 VTAIL.n438 VTAIL.n437 585
R1353 VTAIL.n442 VTAIL.n440 585
R1354 VTAIL.n471 VTAIL.n470 585
R1355 VTAIL.n469 VTAIL.n468 585
R1356 VTAIL.n444 VTAIL.n443 585
R1357 VTAIL.n463 VTAIL.n462 585
R1358 VTAIL.n461 VTAIL.n460 585
R1359 VTAIL.n448 VTAIL.n447 585
R1360 VTAIL.n455 VTAIL.n454 585
R1361 VTAIL.n453 VTAIL.n452 585
R1362 VTAIL.n413 VTAIL.n412 585
R1363 VTAIL.n314 VTAIL.n313 585
R1364 VTAIL.n407 VTAIL.n406 585
R1365 VTAIL.n405 VTAIL.n404 585
R1366 VTAIL.n318 VTAIL.n317 585
R1367 VTAIL.n399 VTAIL.n398 585
R1368 VTAIL.n397 VTAIL.n396 585
R1369 VTAIL.n322 VTAIL.n321 585
R1370 VTAIL.n391 VTAIL.n390 585
R1371 VTAIL.n389 VTAIL.n388 585
R1372 VTAIL.n326 VTAIL.n325 585
R1373 VTAIL.n383 VTAIL.n382 585
R1374 VTAIL.n381 VTAIL.n380 585
R1375 VTAIL.n330 VTAIL.n329 585
R1376 VTAIL.n375 VTAIL.n374 585
R1377 VTAIL.n373 VTAIL.n372 585
R1378 VTAIL.n334 VTAIL.n333 585
R1379 VTAIL.n338 VTAIL.n336 585
R1380 VTAIL.n367 VTAIL.n366 585
R1381 VTAIL.n365 VTAIL.n364 585
R1382 VTAIL.n340 VTAIL.n339 585
R1383 VTAIL.n359 VTAIL.n358 585
R1384 VTAIL.n357 VTAIL.n356 585
R1385 VTAIL.n344 VTAIL.n343 585
R1386 VTAIL.n351 VTAIL.n350 585
R1387 VTAIL.n349 VTAIL.n348 585
R1388 VTAIL.n761 VTAIL.t6 329.036
R1389 VTAIL.n33 VTAIL.t7 329.036
R1390 VTAIL.n137 VTAIL.t3 329.036
R1391 VTAIL.n241 VTAIL.t0 329.036
R1392 VTAIL.n659 VTAIL.t1 329.036
R1393 VTAIL.n555 VTAIL.t2 329.036
R1394 VTAIL.n451 VTAIL.t5 329.036
R1395 VTAIL.n347 VTAIL.t4 329.036
R1396 VTAIL.n764 VTAIL.n763 171.744
R1397 VTAIL.n764 VTAIL.n757 171.744
R1398 VTAIL.n771 VTAIL.n757 171.744
R1399 VTAIL.n772 VTAIL.n771 171.744
R1400 VTAIL.n772 VTAIL.n753 171.744
R1401 VTAIL.n780 VTAIL.n753 171.744
R1402 VTAIL.n781 VTAIL.n780 171.744
R1403 VTAIL.n782 VTAIL.n781 171.744
R1404 VTAIL.n782 VTAIL.n749 171.744
R1405 VTAIL.n789 VTAIL.n749 171.744
R1406 VTAIL.n790 VTAIL.n789 171.744
R1407 VTAIL.n790 VTAIL.n745 171.744
R1408 VTAIL.n797 VTAIL.n745 171.744
R1409 VTAIL.n798 VTAIL.n797 171.744
R1410 VTAIL.n798 VTAIL.n741 171.744
R1411 VTAIL.n805 VTAIL.n741 171.744
R1412 VTAIL.n806 VTAIL.n805 171.744
R1413 VTAIL.n806 VTAIL.n737 171.744
R1414 VTAIL.n813 VTAIL.n737 171.744
R1415 VTAIL.n814 VTAIL.n813 171.744
R1416 VTAIL.n814 VTAIL.n733 171.744
R1417 VTAIL.n821 VTAIL.n733 171.744
R1418 VTAIL.n822 VTAIL.n821 171.744
R1419 VTAIL.n822 VTAIL.n729 171.744
R1420 VTAIL.n829 VTAIL.n729 171.744
R1421 VTAIL.n36 VTAIL.n35 171.744
R1422 VTAIL.n36 VTAIL.n29 171.744
R1423 VTAIL.n43 VTAIL.n29 171.744
R1424 VTAIL.n44 VTAIL.n43 171.744
R1425 VTAIL.n44 VTAIL.n25 171.744
R1426 VTAIL.n52 VTAIL.n25 171.744
R1427 VTAIL.n53 VTAIL.n52 171.744
R1428 VTAIL.n54 VTAIL.n53 171.744
R1429 VTAIL.n54 VTAIL.n21 171.744
R1430 VTAIL.n61 VTAIL.n21 171.744
R1431 VTAIL.n62 VTAIL.n61 171.744
R1432 VTAIL.n62 VTAIL.n17 171.744
R1433 VTAIL.n69 VTAIL.n17 171.744
R1434 VTAIL.n70 VTAIL.n69 171.744
R1435 VTAIL.n70 VTAIL.n13 171.744
R1436 VTAIL.n77 VTAIL.n13 171.744
R1437 VTAIL.n78 VTAIL.n77 171.744
R1438 VTAIL.n78 VTAIL.n9 171.744
R1439 VTAIL.n85 VTAIL.n9 171.744
R1440 VTAIL.n86 VTAIL.n85 171.744
R1441 VTAIL.n86 VTAIL.n5 171.744
R1442 VTAIL.n93 VTAIL.n5 171.744
R1443 VTAIL.n94 VTAIL.n93 171.744
R1444 VTAIL.n94 VTAIL.n1 171.744
R1445 VTAIL.n101 VTAIL.n1 171.744
R1446 VTAIL.n140 VTAIL.n139 171.744
R1447 VTAIL.n140 VTAIL.n133 171.744
R1448 VTAIL.n147 VTAIL.n133 171.744
R1449 VTAIL.n148 VTAIL.n147 171.744
R1450 VTAIL.n148 VTAIL.n129 171.744
R1451 VTAIL.n156 VTAIL.n129 171.744
R1452 VTAIL.n157 VTAIL.n156 171.744
R1453 VTAIL.n158 VTAIL.n157 171.744
R1454 VTAIL.n158 VTAIL.n125 171.744
R1455 VTAIL.n165 VTAIL.n125 171.744
R1456 VTAIL.n166 VTAIL.n165 171.744
R1457 VTAIL.n166 VTAIL.n121 171.744
R1458 VTAIL.n173 VTAIL.n121 171.744
R1459 VTAIL.n174 VTAIL.n173 171.744
R1460 VTAIL.n174 VTAIL.n117 171.744
R1461 VTAIL.n181 VTAIL.n117 171.744
R1462 VTAIL.n182 VTAIL.n181 171.744
R1463 VTAIL.n182 VTAIL.n113 171.744
R1464 VTAIL.n189 VTAIL.n113 171.744
R1465 VTAIL.n190 VTAIL.n189 171.744
R1466 VTAIL.n190 VTAIL.n109 171.744
R1467 VTAIL.n197 VTAIL.n109 171.744
R1468 VTAIL.n198 VTAIL.n197 171.744
R1469 VTAIL.n198 VTAIL.n105 171.744
R1470 VTAIL.n205 VTAIL.n105 171.744
R1471 VTAIL.n244 VTAIL.n243 171.744
R1472 VTAIL.n244 VTAIL.n237 171.744
R1473 VTAIL.n251 VTAIL.n237 171.744
R1474 VTAIL.n252 VTAIL.n251 171.744
R1475 VTAIL.n252 VTAIL.n233 171.744
R1476 VTAIL.n260 VTAIL.n233 171.744
R1477 VTAIL.n261 VTAIL.n260 171.744
R1478 VTAIL.n262 VTAIL.n261 171.744
R1479 VTAIL.n262 VTAIL.n229 171.744
R1480 VTAIL.n269 VTAIL.n229 171.744
R1481 VTAIL.n270 VTAIL.n269 171.744
R1482 VTAIL.n270 VTAIL.n225 171.744
R1483 VTAIL.n277 VTAIL.n225 171.744
R1484 VTAIL.n278 VTAIL.n277 171.744
R1485 VTAIL.n278 VTAIL.n221 171.744
R1486 VTAIL.n285 VTAIL.n221 171.744
R1487 VTAIL.n286 VTAIL.n285 171.744
R1488 VTAIL.n286 VTAIL.n217 171.744
R1489 VTAIL.n293 VTAIL.n217 171.744
R1490 VTAIL.n294 VTAIL.n293 171.744
R1491 VTAIL.n294 VTAIL.n213 171.744
R1492 VTAIL.n301 VTAIL.n213 171.744
R1493 VTAIL.n302 VTAIL.n301 171.744
R1494 VTAIL.n302 VTAIL.n209 171.744
R1495 VTAIL.n309 VTAIL.n209 171.744
R1496 VTAIL.n725 VTAIL.n625 171.744
R1497 VTAIL.n718 VTAIL.n625 171.744
R1498 VTAIL.n718 VTAIL.n717 171.744
R1499 VTAIL.n717 VTAIL.n629 171.744
R1500 VTAIL.n710 VTAIL.n629 171.744
R1501 VTAIL.n710 VTAIL.n709 171.744
R1502 VTAIL.n709 VTAIL.n633 171.744
R1503 VTAIL.n702 VTAIL.n633 171.744
R1504 VTAIL.n702 VTAIL.n701 171.744
R1505 VTAIL.n701 VTAIL.n637 171.744
R1506 VTAIL.n694 VTAIL.n637 171.744
R1507 VTAIL.n694 VTAIL.n693 171.744
R1508 VTAIL.n693 VTAIL.n641 171.744
R1509 VTAIL.n686 VTAIL.n641 171.744
R1510 VTAIL.n686 VTAIL.n685 171.744
R1511 VTAIL.n685 VTAIL.n645 171.744
R1512 VTAIL.n650 VTAIL.n645 171.744
R1513 VTAIL.n678 VTAIL.n650 171.744
R1514 VTAIL.n678 VTAIL.n677 171.744
R1515 VTAIL.n677 VTAIL.n651 171.744
R1516 VTAIL.n670 VTAIL.n651 171.744
R1517 VTAIL.n670 VTAIL.n669 171.744
R1518 VTAIL.n669 VTAIL.n655 171.744
R1519 VTAIL.n662 VTAIL.n655 171.744
R1520 VTAIL.n662 VTAIL.n661 171.744
R1521 VTAIL.n621 VTAIL.n521 171.744
R1522 VTAIL.n614 VTAIL.n521 171.744
R1523 VTAIL.n614 VTAIL.n613 171.744
R1524 VTAIL.n613 VTAIL.n525 171.744
R1525 VTAIL.n606 VTAIL.n525 171.744
R1526 VTAIL.n606 VTAIL.n605 171.744
R1527 VTAIL.n605 VTAIL.n529 171.744
R1528 VTAIL.n598 VTAIL.n529 171.744
R1529 VTAIL.n598 VTAIL.n597 171.744
R1530 VTAIL.n597 VTAIL.n533 171.744
R1531 VTAIL.n590 VTAIL.n533 171.744
R1532 VTAIL.n590 VTAIL.n589 171.744
R1533 VTAIL.n589 VTAIL.n537 171.744
R1534 VTAIL.n582 VTAIL.n537 171.744
R1535 VTAIL.n582 VTAIL.n581 171.744
R1536 VTAIL.n581 VTAIL.n541 171.744
R1537 VTAIL.n546 VTAIL.n541 171.744
R1538 VTAIL.n574 VTAIL.n546 171.744
R1539 VTAIL.n574 VTAIL.n573 171.744
R1540 VTAIL.n573 VTAIL.n547 171.744
R1541 VTAIL.n566 VTAIL.n547 171.744
R1542 VTAIL.n566 VTAIL.n565 171.744
R1543 VTAIL.n565 VTAIL.n551 171.744
R1544 VTAIL.n558 VTAIL.n551 171.744
R1545 VTAIL.n558 VTAIL.n557 171.744
R1546 VTAIL.n517 VTAIL.n417 171.744
R1547 VTAIL.n510 VTAIL.n417 171.744
R1548 VTAIL.n510 VTAIL.n509 171.744
R1549 VTAIL.n509 VTAIL.n421 171.744
R1550 VTAIL.n502 VTAIL.n421 171.744
R1551 VTAIL.n502 VTAIL.n501 171.744
R1552 VTAIL.n501 VTAIL.n425 171.744
R1553 VTAIL.n494 VTAIL.n425 171.744
R1554 VTAIL.n494 VTAIL.n493 171.744
R1555 VTAIL.n493 VTAIL.n429 171.744
R1556 VTAIL.n486 VTAIL.n429 171.744
R1557 VTAIL.n486 VTAIL.n485 171.744
R1558 VTAIL.n485 VTAIL.n433 171.744
R1559 VTAIL.n478 VTAIL.n433 171.744
R1560 VTAIL.n478 VTAIL.n477 171.744
R1561 VTAIL.n477 VTAIL.n437 171.744
R1562 VTAIL.n442 VTAIL.n437 171.744
R1563 VTAIL.n470 VTAIL.n442 171.744
R1564 VTAIL.n470 VTAIL.n469 171.744
R1565 VTAIL.n469 VTAIL.n443 171.744
R1566 VTAIL.n462 VTAIL.n443 171.744
R1567 VTAIL.n462 VTAIL.n461 171.744
R1568 VTAIL.n461 VTAIL.n447 171.744
R1569 VTAIL.n454 VTAIL.n447 171.744
R1570 VTAIL.n454 VTAIL.n453 171.744
R1571 VTAIL.n413 VTAIL.n313 171.744
R1572 VTAIL.n406 VTAIL.n313 171.744
R1573 VTAIL.n406 VTAIL.n405 171.744
R1574 VTAIL.n405 VTAIL.n317 171.744
R1575 VTAIL.n398 VTAIL.n317 171.744
R1576 VTAIL.n398 VTAIL.n397 171.744
R1577 VTAIL.n397 VTAIL.n321 171.744
R1578 VTAIL.n390 VTAIL.n321 171.744
R1579 VTAIL.n390 VTAIL.n389 171.744
R1580 VTAIL.n389 VTAIL.n325 171.744
R1581 VTAIL.n382 VTAIL.n325 171.744
R1582 VTAIL.n382 VTAIL.n381 171.744
R1583 VTAIL.n381 VTAIL.n329 171.744
R1584 VTAIL.n374 VTAIL.n329 171.744
R1585 VTAIL.n374 VTAIL.n373 171.744
R1586 VTAIL.n373 VTAIL.n333 171.744
R1587 VTAIL.n338 VTAIL.n333 171.744
R1588 VTAIL.n366 VTAIL.n338 171.744
R1589 VTAIL.n366 VTAIL.n365 171.744
R1590 VTAIL.n365 VTAIL.n339 171.744
R1591 VTAIL.n358 VTAIL.n339 171.744
R1592 VTAIL.n358 VTAIL.n357 171.744
R1593 VTAIL.n357 VTAIL.n343 171.744
R1594 VTAIL.n350 VTAIL.n343 171.744
R1595 VTAIL.n350 VTAIL.n349 171.744
R1596 VTAIL.n763 VTAIL.t6 85.8723
R1597 VTAIL.n35 VTAIL.t7 85.8723
R1598 VTAIL.n139 VTAIL.t3 85.8723
R1599 VTAIL.n243 VTAIL.t0 85.8723
R1600 VTAIL.n661 VTAIL.t1 85.8723
R1601 VTAIL.n557 VTAIL.t2 85.8723
R1602 VTAIL.n453 VTAIL.t5 85.8723
R1603 VTAIL.n349 VTAIL.t4 85.8723
R1604 VTAIL.n831 VTAIL.n830 34.5126
R1605 VTAIL.n103 VTAIL.n102 34.5126
R1606 VTAIL.n207 VTAIL.n206 34.5126
R1607 VTAIL.n311 VTAIL.n310 34.5126
R1608 VTAIL.n727 VTAIL.n726 34.5126
R1609 VTAIL.n623 VTAIL.n622 34.5126
R1610 VTAIL.n519 VTAIL.n518 34.5126
R1611 VTAIL.n415 VTAIL.n414 34.5126
R1612 VTAIL.n831 VTAIL.n727 30.4531
R1613 VTAIL.n415 VTAIL.n311 30.4531
R1614 VTAIL.n783 VTAIL.n750 13.1884
R1615 VTAIL.n55 VTAIL.n22 13.1884
R1616 VTAIL.n159 VTAIL.n126 13.1884
R1617 VTAIL.n263 VTAIL.n230 13.1884
R1618 VTAIL.n648 VTAIL.n646 13.1884
R1619 VTAIL.n544 VTAIL.n542 13.1884
R1620 VTAIL.n440 VTAIL.n438 13.1884
R1621 VTAIL.n336 VTAIL.n334 13.1884
R1622 VTAIL.n784 VTAIL.n752 12.8005
R1623 VTAIL.n788 VTAIL.n787 12.8005
R1624 VTAIL.n828 VTAIL.n728 12.8005
R1625 VTAIL.n56 VTAIL.n24 12.8005
R1626 VTAIL.n60 VTAIL.n59 12.8005
R1627 VTAIL.n100 VTAIL.n0 12.8005
R1628 VTAIL.n160 VTAIL.n128 12.8005
R1629 VTAIL.n164 VTAIL.n163 12.8005
R1630 VTAIL.n204 VTAIL.n104 12.8005
R1631 VTAIL.n264 VTAIL.n232 12.8005
R1632 VTAIL.n268 VTAIL.n267 12.8005
R1633 VTAIL.n308 VTAIL.n208 12.8005
R1634 VTAIL.n724 VTAIL.n624 12.8005
R1635 VTAIL.n684 VTAIL.n683 12.8005
R1636 VTAIL.n680 VTAIL.n679 12.8005
R1637 VTAIL.n620 VTAIL.n520 12.8005
R1638 VTAIL.n580 VTAIL.n579 12.8005
R1639 VTAIL.n576 VTAIL.n575 12.8005
R1640 VTAIL.n516 VTAIL.n416 12.8005
R1641 VTAIL.n476 VTAIL.n475 12.8005
R1642 VTAIL.n472 VTAIL.n471 12.8005
R1643 VTAIL.n412 VTAIL.n312 12.8005
R1644 VTAIL.n372 VTAIL.n371 12.8005
R1645 VTAIL.n368 VTAIL.n367 12.8005
R1646 VTAIL.n779 VTAIL.n778 12.0247
R1647 VTAIL.n791 VTAIL.n748 12.0247
R1648 VTAIL.n827 VTAIL.n730 12.0247
R1649 VTAIL.n51 VTAIL.n50 12.0247
R1650 VTAIL.n63 VTAIL.n20 12.0247
R1651 VTAIL.n99 VTAIL.n2 12.0247
R1652 VTAIL.n155 VTAIL.n154 12.0247
R1653 VTAIL.n167 VTAIL.n124 12.0247
R1654 VTAIL.n203 VTAIL.n106 12.0247
R1655 VTAIL.n259 VTAIL.n258 12.0247
R1656 VTAIL.n271 VTAIL.n228 12.0247
R1657 VTAIL.n307 VTAIL.n210 12.0247
R1658 VTAIL.n723 VTAIL.n626 12.0247
R1659 VTAIL.n687 VTAIL.n644 12.0247
R1660 VTAIL.n676 VTAIL.n649 12.0247
R1661 VTAIL.n619 VTAIL.n522 12.0247
R1662 VTAIL.n583 VTAIL.n540 12.0247
R1663 VTAIL.n572 VTAIL.n545 12.0247
R1664 VTAIL.n515 VTAIL.n418 12.0247
R1665 VTAIL.n479 VTAIL.n436 12.0247
R1666 VTAIL.n468 VTAIL.n441 12.0247
R1667 VTAIL.n411 VTAIL.n314 12.0247
R1668 VTAIL.n375 VTAIL.n332 12.0247
R1669 VTAIL.n364 VTAIL.n337 12.0247
R1670 VTAIL.n777 VTAIL.n754 11.249
R1671 VTAIL.n792 VTAIL.n746 11.249
R1672 VTAIL.n824 VTAIL.n823 11.249
R1673 VTAIL.n49 VTAIL.n26 11.249
R1674 VTAIL.n64 VTAIL.n18 11.249
R1675 VTAIL.n96 VTAIL.n95 11.249
R1676 VTAIL.n153 VTAIL.n130 11.249
R1677 VTAIL.n168 VTAIL.n122 11.249
R1678 VTAIL.n200 VTAIL.n199 11.249
R1679 VTAIL.n257 VTAIL.n234 11.249
R1680 VTAIL.n272 VTAIL.n226 11.249
R1681 VTAIL.n304 VTAIL.n303 11.249
R1682 VTAIL.n720 VTAIL.n719 11.249
R1683 VTAIL.n688 VTAIL.n642 11.249
R1684 VTAIL.n675 VTAIL.n652 11.249
R1685 VTAIL.n616 VTAIL.n615 11.249
R1686 VTAIL.n584 VTAIL.n538 11.249
R1687 VTAIL.n571 VTAIL.n548 11.249
R1688 VTAIL.n512 VTAIL.n511 11.249
R1689 VTAIL.n480 VTAIL.n434 11.249
R1690 VTAIL.n467 VTAIL.n444 11.249
R1691 VTAIL.n408 VTAIL.n407 11.249
R1692 VTAIL.n376 VTAIL.n330 11.249
R1693 VTAIL.n363 VTAIL.n340 11.249
R1694 VTAIL.n762 VTAIL.n761 10.7239
R1695 VTAIL.n34 VTAIL.n33 10.7239
R1696 VTAIL.n138 VTAIL.n137 10.7239
R1697 VTAIL.n242 VTAIL.n241 10.7239
R1698 VTAIL.n660 VTAIL.n659 10.7239
R1699 VTAIL.n556 VTAIL.n555 10.7239
R1700 VTAIL.n452 VTAIL.n451 10.7239
R1701 VTAIL.n348 VTAIL.n347 10.7239
R1702 VTAIL.n774 VTAIL.n773 10.4732
R1703 VTAIL.n796 VTAIL.n795 10.4732
R1704 VTAIL.n820 VTAIL.n732 10.4732
R1705 VTAIL.n46 VTAIL.n45 10.4732
R1706 VTAIL.n68 VTAIL.n67 10.4732
R1707 VTAIL.n92 VTAIL.n4 10.4732
R1708 VTAIL.n150 VTAIL.n149 10.4732
R1709 VTAIL.n172 VTAIL.n171 10.4732
R1710 VTAIL.n196 VTAIL.n108 10.4732
R1711 VTAIL.n254 VTAIL.n253 10.4732
R1712 VTAIL.n276 VTAIL.n275 10.4732
R1713 VTAIL.n300 VTAIL.n212 10.4732
R1714 VTAIL.n716 VTAIL.n628 10.4732
R1715 VTAIL.n692 VTAIL.n691 10.4732
R1716 VTAIL.n672 VTAIL.n671 10.4732
R1717 VTAIL.n612 VTAIL.n524 10.4732
R1718 VTAIL.n588 VTAIL.n587 10.4732
R1719 VTAIL.n568 VTAIL.n567 10.4732
R1720 VTAIL.n508 VTAIL.n420 10.4732
R1721 VTAIL.n484 VTAIL.n483 10.4732
R1722 VTAIL.n464 VTAIL.n463 10.4732
R1723 VTAIL.n404 VTAIL.n316 10.4732
R1724 VTAIL.n380 VTAIL.n379 10.4732
R1725 VTAIL.n360 VTAIL.n359 10.4732
R1726 VTAIL.n770 VTAIL.n756 9.69747
R1727 VTAIL.n799 VTAIL.n744 9.69747
R1728 VTAIL.n819 VTAIL.n734 9.69747
R1729 VTAIL.n42 VTAIL.n28 9.69747
R1730 VTAIL.n71 VTAIL.n16 9.69747
R1731 VTAIL.n91 VTAIL.n6 9.69747
R1732 VTAIL.n146 VTAIL.n132 9.69747
R1733 VTAIL.n175 VTAIL.n120 9.69747
R1734 VTAIL.n195 VTAIL.n110 9.69747
R1735 VTAIL.n250 VTAIL.n236 9.69747
R1736 VTAIL.n279 VTAIL.n224 9.69747
R1737 VTAIL.n299 VTAIL.n214 9.69747
R1738 VTAIL.n715 VTAIL.n630 9.69747
R1739 VTAIL.n695 VTAIL.n640 9.69747
R1740 VTAIL.n668 VTAIL.n654 9.69747
R1741 VTAIL.n611 VTAIL.n526 9.69747
R1742 VTAIL.n591 VTAIL.n536 9.69747
R1743 VTAIL.n564 VTAIL.n550 9.69747
R1744 VTAIL.n507 VTAIL.n422 9.69747
R1745 VTAIL.n487 VTAIL.n432 9.69747
R1746 VTAIL.n460 VTAIL.n446 9.69747
R1747 VTAIL.n403 VTAIL.n318 9.69747
R1748 VTAIL.n383 VTAIL.n328 9.69747
R1749 VTAIL.n356 VTAIL.n342 9.69747
R1750 VTAIL.n826 VTAIL.n728 9.45567
R1751 VTAIL.n98 VTAIL.n0 9.45567
R1752 VTAIL.n202 VTAIL.n104 9.45567
R1753 VTAIL.n306 VTAIL.n208 9.45567
R1754 VTAIL.n722 VTAIL.n624 9.45567
R1755 VTAIL.n618 VTAIL.n520 9.45567
R1756 VTAIL.n514 VTAIL.n416 9.45567
R1757 VTAIL.n410 VTAIL.n312 9.45567
R1758 VTAIL.n809 VTAIL.n808 9.3005
R1759 VTAIL.n811 VTAIL.n810 9.3005
R1760 VTAIL.n736 VTAIL.n735 9.3005
R1761 VTAIL.n817 VTAIL.n816 9.3005
R1762 VTAIL.n819 VTAIL.n818 9.3005
R1763 VTAIL.n732 VTAIL.n731 9.3005
R1764 VTAIL.n825 VTAIL.n824 9.3005
R1765 VTAIL.n827 VTAIL.n826 9.3005
R1766 VTAIL.n803 VTAIL.n802 9.3005
R1767 VTAIL.n801 VTAIL.n800 9.3005
R1768 VTAIL.n744 VTAIL.n743 9.3005
R1769 VTAIL.n795 VTAIL.n794 9.3005
R1770 VTAIL.n793 VTAIL.n792 9.3005
R1771 VTAIL.n748 VTAIL.n747 9.3005
R1772 VTAIL.n787 VTAIL.n786 9.3005
R1773 VTAIL.n760 VTAIL.n759 9.3005
R1774 VTAIL.n767 VTAIL.n766 9.3005
R1775 VTAIL.n769 VTAIL.n768 9.3005
R1776 VTAIL.n756 VTAIL.n755 9.3005
R1777 VTAIL.n775 VTAIL.n774 9.3005
R1778 VTAIL.n777 VTAIL.n776 9.3005
R1779 VTAIL.n778 VTAIL.n751 9.3005
R1780 VTAIL.n785 VTAIL.n784 9.3005
R1781 VTAIL.n740 VTAIL.n739 9.3005
R1782 VTAIL.n81 VTAIL.n80 9.3005
R1783 VTAIL.n83 VTAIL.n82 9.3005
R1784 VTAIL.n8 VTAIL.n7 9.3005
R1785 VTAIL.n89 VTAIL.n88 9.3005
R1786 VTAIL.n91 VTAIL.n90 9.3005
R1787 VTAIL.n4 VTAIL.n3 9.3005
R1788 VTAIL.n97 VTAIL.n96 9.3005
R1789 VTAIL.n99 VTAIL.n98 9.3005
R1790 VTAIL.n75 VTAIL.n74 9.3005
R1791 VTAIL.n73 VTAIL.n72 9.3005
R1792 VTAIL.n16 VTAIL.n15 9.3005
R1793 VTAIL.n67 VTAIL.n66 9.3005
R1794 VTAIL.n65 VTAIL.n64 9.3005
R1795 VTAIL.n20 VTAIL.n19 9.3005
R1796 VTAIL.n59 VTAIL.n58 9.3005
R1797 VTAIL.n32 VTAIL.n31 9.3005
R1798 VTAIL.n39 VTAIL.n38 9.3005
R1799 VTAIL.n41 VTAIL.n40 9.3005
R1800 VTAIL.n28 VTAIL.n27 9.3005
R1801 VTAIL.n47 VTAIL.n46 9.3005
R1802 VTAIL.n49 VTAIL.n48 9.3005
R1803 VTAIL.n50 VTAIL.n23 9.3005
R1804 VTAIL.n57 VTAIL.n56 9.3005
R1805 VTAIL.n12 VTAIL.n11 9.3005
R1806 VTAIL.n185 VTAIL.n184 9.3005
R1807 VTAIL.n187 VTAIL.n186 9.3005
R1808 VTAIL.n112 VTAIL.n111 9.3005
R1809 VTAIL.n193 VTAIL.n192 9.3005
R1810 VTAIL.n195 VTAIL.n194 9.3005
R1811 VTAIL.n108 VTAIL.n107 9.3005
R1812 VTAIL.n201 VTAIL.n200 9.3005
R1813 VTAIL.n203 VTAIL.n202 9.3005
R1814 VTAIL.n179 VTAIL.n178 9.3005
R1815 VTAIL.n177 VTAIL.n176 9.3005
R1816 VTAIL.n120 VTAIL.n119 9.3005
R1817 VTAIL.n171 VTAIL.n170 9.3005
R1818 VTAIL.n169 VTAIL.n168 9.3005
R1819 VTAIL.n124 VTAIL.n123 9.3005
R1820 VTAIL.n163 VTAIL.n162 9.3005
R1821 VTAIL.n136 VTAIL.n135 9.3005
R1822 VTAIL.n143 VTAIL.n142 9.3005
R1823 VTAIL.n145 VTAIL.n144 9.3005
R1824 VTAIL.n132 VTAIL.n131 9.3005
R1825 VTAIL.n151 VTAIL.n150 9.3005
R1826 VTAIL.n153 VTAIL.n152 9.3005
R1827 VTAIL.n154 VTAIL.n127 9.3005
R1828 VTAIL.n161 VTAIL.n160 9.3005
R1829 VTAIL.n116 VTAIL.n115 9.3005
R1830 VTAIL.n289 VTAIL.n288 9.3005
R1831 VTAIL.n291 VTAIL.n290 9.3005
R1832 VTAIL.n216 VTAIL.n215 9.3005
R1833 VTAIL.n297 VTAIL.n296 9.3005
R1834 VTAIL.n299 VTAIL.n298 9.3005
R1835 VTAIL.n212 VTAIL.n211 9.3005
R1836 VTAIL.n305 VTAIL.n304 9.3005
R1837 VTAIL.n307 VTAIL.n306 9.3005
R1838 VTAIL.n283 VTAIL.n282 9.3005
R1839 VTAIL.n281 VTAIL.n280 9.3005
R1840 VTAIL.n224 VTAIL.n223 9.3005
R1841 VTAIL.n275 VTAIL.n274 9.3005
R1842 VTAIL.n273 VTAIL.n272 9.3005
R1843 VTAIL.n228 VTAIL.n227 9.3005
R1844 VTAIL.n267 VTAIL.n266 9.3005
R1845 VTAIL.n240 VTAIL.n239 9.3005
R1846 VTAIL.n247 VTAIL.n246 9.3005
R1847 VTAIL.n249 VTAIL.n248 9.3005
R1848 VTAIL.n236 VTAIL.n235 9.3005
R1849 VTAIL.n255 VTAIL.n254 9.3005
R1850 VTAIL.n257 VTAIL.n256 9.3005
R1851 VTAIL.n258 VTAIL.n231 9.3005
R1852 VTAIL.n265 VTAIL.n264 9.3005
R1853 VTAIL.n220 VTAIL.n219 9.3005
R1854 VTAIL.n723 VTAIL.n722 9.3005
R1855 VTAIL.n721 VTAIL.n720 9.3005
R1856 VTAIL.n628 VTAIL.n627 9.3005
R1857 VTAIL.n715 VTAIL.n714 9.3005
R1858 VTAIL.n713 VTAIL.n712 9.3005
R1859 VTAIL.n632 VTAIL.n631 9.3005
R1860 VTAIL.n707 VTAIL.n706 9.3005
R1861 VTAIL.n705 VTAIL.n704 9.3005
R1862 VTAIL.n636 VTAIL.n635 9.3005
R1863 VTAIL.n699 VTAIL.n698 9.3005
R1864 VTAIL.n697 VTAIL.n696 9.3005
R1865 VTAIL.n640 VTAIL.n639 9.3005
R1866 VTAIL.n691 VTAIL.n690 9.3005
R1867 VTAIL.n689 VTAIL.n688 9.3005
R1868 VTAIL.n644 VTAIL.n643 9.3005
R1869 VTAIL.n683 VTAIL.n682 9.3005
R1870 VTAIL.n681 VTAIL.n680 9.3005
R1871 VTAIL.n649 VTAIL.n647 9.3005
R1872 VTAIL.n675 VTAIL.n674 9.3005
R1873 VTAIL.n673 VTAIL.n672 9.3005
R1874 VTAIL.n654 VTAIL.n653 9.3005
R1875 VTAIL.n667 VTAIL.n666 9.3005
R1876 VTAIL.n665 VTAIL.n664 9.3005
R1877 VTAIL.n658 VTAIL.n657 9.3005
R1878 VTAIL.n554 VTAIL.n553 9.3005
R1879 VTAIL.n561 VTAIL.n560 9.3005
R1880 VTAIL.n563 VTAIL.n562 9.3005
R1881 VTAIL.n550 VTAIL.n549 9.3005
R1882 VTAIL.n569 VTAIL.n568 9.3005
R1883 VTAIL.n571 VTAIL.n570 9.3005
R1884 VTAIL.n545 VTAIL.n543 9.3005
R1885 VTAIL.n577 VTAIL.n576 9.3005
R1886 VTAIL.n603 VTAIL.n602 9.3005
R1887 VTAIL.n528 VTAIL.n527 9.3005
R1888 VTAIL.n609 VTAIL.n608 9.3005
R1889 VTAIL.n611 VTAIL.n610 9.3005
R1890 VTAIL.n524 VTAIL.n523 9.3005
R1891 VTAIL.n617 VTAIL.n616 9.3005
R1892 VTAIL.n619 VTAIL.n618 9.3005
R1893 VTAIL.n601 VTAIL.n600 9.3005
R1894 VTAIL.n532 VTAIL.n531 9.3005
R1895 VTAIL.n595 VTAIL.n594 9.3005
R1896 VTAIL.n593 VTAIL.n592 9.3005
R1897 VTAIL.n536 VTAIL.n535 9.3005
R1898 VTAIL.n587 VTAIL.n586 9.3005
R1899 VTAIL.n585 VTAIL.n584 9.3005
R1900 VTAIL.n540 VTAIL.n539 9.3005
R1901 VTAIL.n579 VTAIL.n578 9.3005
R1902 VTAIL.n450 VTAIL.n449 9.3005
R1903 VTAIL.n457 VTAIL.n456 9.3005
R1904 VTAIL.n459 VTAIL.n458 9.3005
R1905 VTAIL.n446 VTAIL.n445 9.3005
R1906 VTAIL.n465 VTAIL.n464 9.3005
R1907 VTAIL.n467 VTAIL.n466 9.3005
R1908 VTAIL.n441 VTAIL.n439 9.3005
R1909 VTAIL.n473 VTAIL.n472 9.3005
R1910 VTAIL.n499 VTAIL.n498 9.3005
R1911 VTAIL.n424 VTAIL.n423 9.3005
R1912 VTAIL.n505 VTAIL.n504 9.3005
R1913 VTAIL.n507 VTAIL.n506 9.3005
R1914 VTAIL.n420 VTAIL.n419 9.3005
R1915 VTAIL.n513 VTAIL.n512 9.3005
R1916 VTAIL.n515 VTAIL.n514 9.3005
R1917 VTAIL.n497 VTAIL.n496 9.3005
R1918 VTAIL.n428 VTAIL.n427 9.3005
R1919 VTAIL.n491 VTAIL.n490 9.3005
R1920 VTAIL.n489 VTAIL.n488 9.3005
R1921 VTAIL.n432 VTAIL.n431 9.3005
R1922 VTAIL.n483 VTAIL.n482 9.3005
R1923 VTAIL.n481 VTAIL.n480 9.3005
R1924 VTAIL.n436 VTAIL.n435 9.3005
R1925 VTAIL.n475 VTAIL.n474 9.3005
R1926 VTAIL.n346 VTAIL.n345 9.3005
R1927 VTAIL.n353 VTAIL.n352 9.3005
R1928 VTAIL.n355 VTAIL.n354 9.3005
R1929 VTAIL.n342 VTAIL.n341 9.3005
R1930 VTAIL.n361 VTAIL.n360 9.3005
R1931 VTAIL.n363 VTAIL.n362 9.3005
R1932 VTAIL.n337 VTAIL.n335 9.3005
R1933 VTAIL.n369 VTAIL.n368 9.3005
R1934 VTAIL.n395 VTAIL.n394 9.3005
R1935 VTAIL.n320 VTAIL.n319 9.3005
R1936 VTAIL.n401 VTAIL.n400 9.3005
R1937 VTAIL.n403 VTAIL.n402 9.3005
R1938 VTAIL.n316 VTAIL.n315 9.3005
R1939 VTAIL.n409 VTAIL.n408 9.3005
R1940 VTAIL.n411 VTAIL.n410 9.3005
R1941 VTAIL.n393 VTAIL.n392 9.3005
R1942 VTAIL.n324 VTAIL.n323 9.3005
R1943 VTAIL.n387 VTAIL.n386 9.3005
R1944 VTAIL.n385 VTAIL.n384 9.3005
R1945 VTAIL.n328 VTAIL.n327 9.3005
R1946 VTAIL.n379 VTAIL.n378 9.3005
R1947 VTAIL.n377 VTAIL.n376 9.3005
R1948 VTAIL.n332 VTAIL.n331 9.3005
R1949 VTAIL.n371 VTAIL.n370 9.3005
R1950 VTAIL.n769 VTAIL.n758 8.92171
R1951 VTAIL.n800 VTAIL.n742 8.92171
R1952 VTAIL.n816 VTAIL.n815 8.92171
R1953 VTAIL.n41 VTAIL.n30 8.92171
R1954 VTAIL.n72 VTAIL.n14 8.92171
R1955 VTAIL.n88 VTAIL.n87 8.92171
R1956 VTAIL.n145 VTAIL.n134 8.92171
R1957 VTAIL.n176 VTAIL.n118 8.92171
R1958 VTAIL.n192 VTAIL.n191 8.92171
R1959 VTAIL.n249 VTAIL.n238 8.92171
R1960 VTAIL.n280 VTAIL.n222 8.92171
R1961 VTAIL.n296 VTAIL.n295 8.92171
R1962 VTAIL.n712 VTAIL.n711 8.92171
R1963 VTAIL.n696 VTAIL.n638 8.92171
R1964 VTAIL.n667 VTAIL.n656 8.92171
R1965 VTAIL.n608 VTAIL.n607 8.92171
R1966 VTAIL.n592 VTAIL.n534 8.92171
R1967 VTAIL.n563 VTAIL.n552 8.92171
R1968 VTAIL.n504 VTAIL.n503 8.92171
R1969 VTAIL.n488 VTAIL.n430 8.92171
R1970 VTAIL.n459 VTAIL.n448 8.92171
R1971 VTAIL.n400 VTAIL.n399 8.92171
R1972 VTAIL.n384 VTAIL.n326 8.92171
R1973 VTAIL.n355 VTAIL.n344 8.92171
R1974 VTAIL.n766 VTAIL.n765 8.14595
R1975 VTAIL.n804 VTAIL.n803 8.14595
R1976 VTAIL.n812 VTAIL.n736 8.14595
R1977 VTAIL.n38 VTAIL.n37 8.14595
R1978 VTAIL.n76 VTAIL.n75 8.14595
R1979 VTAIL.n84 VTAIL.n8 8.14595
R1980 VTAIL.n142 VTAIL.n141 8.14595
R1981 VTAIL.n180 VTAIL.n179 8.14595
R1982 VTAIL.n188 VTAIL.n112 8.14595
R1983 VTAIL.n246 VTAIL.n245 8.14595
R1984 VTAIL.n284 VTAIL.n283 8.14595
R1985 VTAIL.n292 VTAIL.n216 8.14595
R1986 VTAIL.n708 VTAIL.n632 8.14595
R1987 VTAIL.n700 VTAIL.n699 8.14595
R1988 VTAIL.n664 VTAIL.n663 8.14595
R1989 VTAIL.n604 VTAIL.n528 8.14595
R1990 VTAIL.n596 VTAIL.n595 8.14595
R1991 VTAIL.n560 VTAIL.n559 8.14595
R1992 VTAIL.n500 VTAIL.n424 8.14595
R1993 VTAIL.n492 VTAIL.n491 8.14595
R1994 VTAIL.n456 VTAIL.n455 8.14595
R1995 VTAIL.n396 VTAIL.n320 8.14595
R1996 VTAIL.n388 VTAIL.n387 8.14595
R1997 VTAIL.n352 VTAIL.n351 8.14595
R1998 VTAIL.n762 VTAIL.n760 7.3702
R1999 VTAIL.n807 VTAIL.n740 7.3702
R2000 VTAIL.n811 VTAIL.n738 7.3702
R2001 VTAIL.n34 VTAIL.n32 7.3702
R2002 VTAIL.n79 VTAIL.n12 7.3702
R2003 VTAIL.n83 VTAIL.n10 7.3702
R2004 VTAIL.n138 VTAIL.n136 7.3702
R2005 VTAIL.n183 VTAIL.n116 7.3702
R2006 VTAIL.n187 VTAIL.n114 7.3702
R2007 VTAIL.n242 VTAIL.n240 7.3702
R2008 VTAIL.n287 VTAIL.n220 7.3702
R2009 VTAIL.n291 VTAIL.n218 7.3702
R2010 VTAIL.n707 VTAIL.n634 7.3702
R2011 VTAIL.n703 VTAIL.n636 7.3702
R2012 VTAIL.n660 VTAIL.n658 7.3702
R2013 VTAIL.n603 VTAIL.n530 7.3702
R2014 VTAIL.n599 VTAIL.n532 7.3702
R2015 VTAIL.n556 VTAIL.n554 7.3702
R2016 VTAIL.n499 VTAIL.n426 7.3702
R2017 VTAIL.n495 VTAIL.n428 7.3702
R2018 VTAIL.n452 VTAIL.n450 7.3702
R2019 VTAIL.n395 VTAIL.n322 7.3702
R2020 VTAIL.n391 VTAIL.n324 7.3702
R2021 VTAIL.n348 VTAIL.n346 7.3702
R2022 VTAIL.n808 VTAIL.n807 6.59444
R2023 VTAIL.n808 VTAIL.n738 6.59444
R2024 VTAIL.n80 VTAIL.n79 6.59444
R2025 VTAIL.n80 VTAIL.n10 6.59444
R2026 VTAIL.n184 VTAIL.n183 6.59444
R2027 VTAIL.n184 VTAIL.n114 6.59444
R2028 VTAIL.n288 VTAIL.n287 6.59444
R2029 VTAIL.n288 VTAIL.n218 6.59444
R2030 VTAIL.n704 VTAIL.n634 6.59444
R2031 VTAIL.n704 VTAIL.n703 6.59444
R2032 VTAIL.n600 VTAIL.n530 6.59444
R2033 VTAIL.n600 VTAIL.n599 6.59444
R2034 VTAIL.n496 VTAIL.n426 6.59444
R2035 VTAIL.n496 VTAIL.n495 6.59444
R2036 VTAIL.n392 VTAIL.n322 6.59444
R2037 VTAIL.n392 VTAIL.n391 6.59444
R2038 VTAIL.n765 VTAIL.n760 5.81868
R2039 VTAIL.n804 VTAIL.n740 5.81868
R2040 VTAIL.n812 VTAIL.n811 5.81868
R2041 VTAIL.n37 VTAIL.n32 5.81868
R2042 VTAIL.n76 VTAIL.n12 5.81868
R2043 VTAIL.n84 VTAIL.n83 5.81868
R2044 VTAIL.n141 VTAIL.n136 5.81868
R2045 VTAIL.n180 VTAIL.n116 5.81868
R2046 VTAIL.n188 VTAIL.n187 5.81868
R2047 VTAIL.n245 VTAIL.n240 5.81868
R2048 VTAIL.n284 VTAIL.n220 5.81868
R2049 VTAIL.n292 VTAIL.n291 5.81868
R2050 VTAIL.n708 VTAIL.n707 5.81868
R2051 VTAIL.n700 VTAIL.n636 5.81868
R2052 VTAIL.n663 VTAIL.n658 5.81868
R2053 VTAIL.n604 VTAIL.n603 5.81868
R2054 VTAIL.n596 VTAIL.n532 5.81868
R2055 VTAIL.n559 VTAIL.n554 5.81868
R2056 VTAIL.n500 VTAIL.n499 5.81868
R2057 VTAIL.n492 VTAIL.n428 5.81868
R2058 VTAIL.n455 VTAIL.n450 5.81868
R2059 VTAIL.n396 VTAIL.n395 5.81868
R2060 VTAIL.n388 VTAIL.n324 5.81868
R2061 VTAIL.n351 VTAIL.n346 5.81868
R2062 VTAIL.n766 VTAIL.n758 5.04292
R2063 VTAIL.n803 VTAIL.n742 5.04292
R2064 VTAIL.n815 VTAIL.n736 5.04292
R2065 VTAIL.n38 VTAIL.n30 5.04292
R2066 VTAIL.n75 VTAIL.n14 5.04292
R2067 VTAIL.n87 VTAIL.n8 5.04292
R2068 VTAIL.n142 VTAIL.n134 5.04292
R2069 VTAIL.n179 VTAIL.n118 5.04292
R2070 VTAIL.n191 VTAIL.n112 5.04292
R2071 VTAIL.n246 VTAIL.n238 5.04292
R2072 VTAIL.n283 VTAIL.n222 5.04292
R2073 VTAIL.n295 VTAIL.n216 5.04292
R2074 VTAIL.n711 VTAIL.n632 5.04292
R2075 VTAIL.n699 VTAIL.n638 5.04292
R2076 VTAIL.n664 VTAIL.n656 5.04292
R2077 VTAIL.n607 VTAIL.n528 5.04292
R2078 VTAIL.n595 VTAIL.n534 5.04292
R2079 VTAIL.n560 VTAIL.n552 5.04292
R2080 VTAIL.n503 VTAIL.n424 5.04292
R2081 VTAIL.n491 VTAIL.n430 5.04292
R2082 VTAIL.n456 VTAIL.n448 5.04292
R2083 VTAIL.n399 VTAIL.n320 5.04292
R2084 VTAIL.n387 VTAIL.n326 5.04292
R2085 VTAIL.n352 VTAIL.n344 5.04292
R2086 VTAIL.n770 VTAIL.n769 4.26717
R2087 VTAIL.n800 VTAIL.n799 4.26717
R2088 VTAIL.n816 VTAIL.n734 4.26717
R2089 VTAIL.n42 VTAIL.n41 4.26717
R2090 VTAIL.n72 VTAIL.n71 4.26717
R2091 VTAIL.n88 VTAIL.n6 4.26717
R2092 VTAIL.n146 VTAIL.n145 4.26717
R2093 VTAIL.n176 VTAIL.n175 4.26717
R2094 VTAIL.n192 VTAIL.n110 4.26717
R2095 VTAIL.n250 VTAIL.n249 4.26717
R2096 VTAIL.n280 VTAIL.n279 4.26717
R2097 VTAIL.n296 VTAIL.n214 4.26717
R2098 VTAIL.n712 VTAIL.n630 4.26717
R2099 VTAIL.n696 VTAIL.n695 4.26717
R2100 VTAIL.n668 VTAIL.n667 4.26717
R2101 VTAIL.n608 VTAIL.n526 4.26717
R2102 VTAIL.n592 VTAIL.n591 4.26717
R2103 VTAIL.n564 VTAIL.n563 4.26717
R2104 VTAIL.n504 VTAIL.n422 4.26717
R2105 VTAIL.n488 VTAIL.n487 4.26717
R2106 VTAIL.n460 VTAIL.n459 4.26717
R2107 VTAIL.n400 VTAIL.n318 4.26717
R2108 VTAIL.n384 VTAIL.n383 4.26717
R2109 VTAIL.n356 VTAIL.n355 4.26717
R2110 VTAIL.n773 VTAIL.n756 3.49141
R2111 VTAIL.n796 VTAIL.n744 3.49141
R2112 VTAIL.n820 VTAIL.n819 3.49141
R2113 VTAIL.n45 VTAIL.n28 3.49141
R2114 VTAIL.n68 VTAIL.n16 3.49141
R2115 VTAIL.n92 VTAIL.n91 3.49141
R2116 VTAIL.n149 VTAIL.n132 3.49141
R2117 VTAIL.n172 VTAIL.n120 3.49141
R2118 VTAIL.n196 VTAIL.n195 3.49141
R2119 VTAIL.n253 VTAIL.n236 3.49141
R2120 VTAIL.n276 VTAIL.n224 3.49141
R2121 VTAIL.n300 VTAIL.n299 3.49141
R2122 VTAIL.n716 VTAIL.n715 3.49141
R2123 VTAIL.n692 VTAIL.n640 3.49141
R2124 VTAIL.n671 VTAIL.n654 3.49141
R2125 VTAIL.n612 VTAIL.n611 3.49141
R2126 VTAIL.n588 VTAIL.n536 3.49141
R2127 VTAIL.n567 VTAIL.n550 3.49141
R2128 VTAIL.n508 VTAIL.n507 3.49141
R2129 VTAIL.n484 VTAIL.n432 3.49141
R2130 VTAIL.n463 VTAIL.n446 3.49141
R2131 VTAIL.n404 VTAIL.n403 3.49141
R2132 VTAIL.n380 VTAIL.n328 3.49141
R2133 VTAIL.n359 VTAIL.n342 3.49141
R2134 VTAIL.n774 VTAIL.n754 2.71565
R2135 VTAIL.n795 VTAIL.n746 2.71565
R2136 VTAIL.n823 VTAIL.n732 2.71565
R2137 VTAIL.n46 VTAIL.n26 2.71565
R2138 VTAIL.n67 VTAIL.n18 2.71565
R2139 VTAIL.n95 VTAIL.n4 2.71565
R2140 VTAIL.n150 VTAIL.n130 2.71565
R2141 VTAIL.n171 VTAIL.n122 2.71565
R2142 VTAIL.n199 VTAIL.n108 2.71565
R2143 VTAIL.n254 VTAIL.n234 2.71565
R2144 VTAIL.n275 VTAIL.n226 2.71565
R2145 VTAIL.n303 VTAIL.n212 2.71565
R2146 VTAIL.n719 VTAIL.n628 2.71565
R2147 VTAIL.n691 VTAIL.n642 2.71565
R2148 VTAIL.n672 VTAIL.n652 2.71565
R2149 VTAIL.n615 VTAIL.n524 2.71565
R2150 VTAIL.n587 VTAIL.n538 2.71565
R2151 VTAIL.n568 VTAIL.n548 2.71565
R2152 VTAIL.n511 VTAIL.n420 2.71565
R2153 VTAIL.n483 VTAIL.n434 2.71565
R2154 VTAIL.n464 VTAIL.n444 2.71565
R2155 VTAIL.n407 VTAIL.n316 2.71565
R2156 VTAIL.n379 VTAIL.n330 2.71565
R2157 VTAIL.n360 VTAIL.n340 2.71565
R2158 VTAIL.n659 VTAIL.n657 2.41282
R2159 VTAIL.n555 VTAIL.n553 2.41282
R2160 VTAIL.n451 VTAIL.n449 2.41282
R2161 VTAIL.n347 VTAIL.n345 2.41282
R2162 VTAIL.n761 VTAIL.n759 2.41282
R2163 VTAIL.n33 VTAIL.n31 2.41282
R2164 VTAIL.n137 VTAIL.n135 2.41282
R2165 VTAIL.n241 VTAIL.n239 2.41282
R2166 VTAIL.n779 VTAIL.n777 1.93989
R2167 VTAIL.n792 VTAIL.n791 1.93989
R2168 VTAIL.n824 VTAIL.n730 1.93989
R2169 VTAIL.n51 VTAIL.n49 1.93989
R2170 VTAIL.n64 VTAIL.n63 1.93989
R2171 VTAIL.n96 VTAIL.n2 1.93989
R2172 VTAIL.n155 VTAIL.n153 1.93989
R2173 VTAIL.n168 VTAIL.n167 1.93989
R2174 VTAIL.n200 VTAIL.n106 1.93989
R2175 VTAIL.n259 VTAIL.n257 1.93989
R2176 VTAIL.n272 VTAIL.n271 1.93989
R2177 VTAIL.n304 VTAIL.n210 1.93989
R2178 VTAIL.n720 VTAIL.n626 1.93989
R2179 VTAIL.n688 VTAIL.n687 1.93989
R2180 VTAIL.n676 VTAIL.n675 1.93989
R2181 VTAIL.n616 VTAIL.n522 1.93989
R2182 VTAIL.n584 VTAIL.n583 1.93989
R2183 VTAIL.n572 VTAIL.n571 1.93989
R2184 VTAIL.n512 VTAIL.n418 1.93989
R2185 VTAIL.n480 VTAIL.n479 1.93989
R2186 VTAIL.n468 VTAIL.n467 1.93989
R2187 VTAIL.n408 VTAIL.n314 1.93989
R2188 VTAIL.n376 VTAIL.n375 1.93989
R2189 VTAIL.n364 VTAIL.n363 1.93989
R2190 VTAIL.n519 VTAIL.n415 1.93153
R2191 VTAIL.n727 VTAIL.n623 1.93153
R2192 VTAIL.n311 VTAIL.n207 1.93153
R2193 VTAIL.n778 VTAIL.n752 1.16414
R2194 VTAIL.n788 VTAIL.n748 1.16414
R2195 VTAIL.n828 VTAIL.n827 1.16414
R2196 VTAIL.n50 VTAIL.n24 1.16414
R2197 VTAIL.n60 VTAIL.n20 1.16414
R2198 VTAIL.n100 VTAIL.n99 1.16414
R2199 VTAIL.n154 VTAIL.n128 1.16414
R2200 VTAIL.n164 VTAIL.n124 1.16414
R2201 VTAIL.n204 VTAIL.n203 1.16414
R2202 VTAIL.n258 VTAIL.n232 1.16414
R2203 VTAIL.n268 VTAIL.n228 1.16414
R2204 VTAIL.n308 VTAIL.n307 1.16414
R2205 VTAIL.n724 VTAIL.n723 1.16414
R2206 VTAIL.n684 VTAIL.n644 1.16414
R2207 VTAIL.n679 VTAIL.n649 1.16414
R2208 VTAIL.n620 VTAIL.n619 1.16414
R2209 VTAIL.n580 VTAIL.n540 1.16414
R2210 VTAIL.n575 VTAIL.n545 1.16414
R2211 VTAIL.n516 VTAIL.n515 1.16414
R2212 VTAIL.n476 VTAIL.n436 1.16414
R2213 VTAIL.n471 VTAIL.n441 1.16414
R2214 VTAIL.n412 VTAIL.n411 1.16414
R2215 VTAIL.n372 VTAIL.n332 1.16414
R2216 VTAIL.n367 VTAIL.n337 1.16414
R2217 VTAIL VTAIL.n103 1.02421
R2218 VTAIL VTAIL.n831 0.907828
R2219 VTAIL.n623 VTAIL.n519 0.470328
R2220 VTAIL.n207 VTAIL.n103 0.470328
R2221 VTAIL.n784 VTAIL.n783 0.388379
R2222 VTAIL.n787 VTAIL.n750 0.388379
R2223 VTAIL.n830 VTAIL.n728 0.388379
R2224 VTAIL.n56 VTAIL.n55 0.388379
R2225 VTAIL.n59 VTAIL.n22 0.388379
R2226 VTAIL.n102 VTAIL.n0 0.388379
R2227 VTAIL.n160 VTAIL.n159 0.388379
R2228 VTAIL.n163 VTAIL.n126 0.388379
R2229 VTAIL.n206 VTAIL.n104 0.388379
R2230 VTAIL.n264 VTAIL.n263 0.388379
R2231 VTAIL.n267 VTAIL.n230 0.388379
R2232 VTAIL.n310 VTAIL.n208 0.388379
R2233 VTAIL.n726 VTAIL.n624 0.388379
R2234 VTAIL.n683 VTAIL.n646 0.388379
R2235 VTAIL.n680 VTAIL.n648 0.388379
R2236 VTAIL.n622 VTAIL.n520 0.388379
R2237 VTAIL.n579 VTAIL.n542 0.388379
R2238 VTAIL.n576 VTAIL.n544 0.388379
R2239 VTAIL.n518 VTAIL.n416 0.388379
R2240 VTAIL.n475 VTAIL.n438 0.388379
R2241 VTAIL.n472 VTAIL.n440 0.388379
R2242 VTAIL.n414 VTAIL.n312 0.388379
R2243 VTAIL.n371 VTAIL.n334 0.388379
R2244 VTAIL.n368 VTAIL.n336 0.388379
R2245 VTAIL.n767 VTAIL.n759 0.155672
R2246 VTAIL.n768 VTAIL.n767 0.155672
R2247 VTAIL.n768 VTAIL.n755 0.155672
R2248 VTAIL.n775 VTAIL.n755 0.155672
R2249 VTAIL.n776 VTAIL.n775 0.155672
R2250 VTAIL.n776 VTAIL.n751 0.155672
R2251 VTAIL.n785 VTAIL.n751 0.155672
R2252 VTAIL.n786 VTAIL.n785 0.155672
R2253 VTAIL.n786 VTAIL.n747 0.155672
R2254 VTAIL.n793 VTAIL.n747 0.155672
R2255 VTAIL.n794 VTAIL.n793 0.155672
R2256 VTAIL.n794 VTAIL.n743 0.155672
R2257 VTAIL.n801 VTAIL.n743 0.155672
R2258 VTAIL.n802 VTAIL.n801 0.155672
R2259 VTAIL.n802 VTAIL.n739 0.155672
R2260 VTAIL.n809 VTAIL.n739 0.155672
R2261 VTAIL.n810 VTAIL.n809 0.155672
R2262 VTAIL.n810 VTAIL.n735 0.155672
R2263 VTAIL.n817 VTAIL.n735 0.155672
R2264 VTAIL.n818 VTAIL.n817 0.155672
R2265 VTAIL.n818 VTAIL.n731 0.155672
R2266 VTAIL.n825 VTAIL.n731 0.155672
R2267 VTAIL.n826 VTAIL.n825 0.155672
R2268 VTAIL.n39 VTAIL.n31 0.155672
R2269 VTAIL.n40 VTAIL.n39 0.155672
R2270 VTAIL.n40 VTAIL.n27 0.155672
R2271 VTAIL.n47 VTAIL.n27 0.155672
R2272 VTAIL.n48 VTAIL.n47 0.155672
R2273 VTAIL.n48 VTAIL.n23 0.155672
R2274 VTAIL.n57 VTAIL.n23 0.155672
R2275 VTAIL.n58 VTAIL.n57 0.155672
R2276 VTAIL.n58 VTAIL.n19 0.155672
R2277 VTAIL.n65 VTAIL.n19 0.155672
R2278 VTAIL.n66 VTAIL.n65 0.155672
R2279 VTAIL.n66 VTAIL.n15 0.155672
R2280 VTAIL.n73 VTAIL.n15 0.155672
R2281 VTAIL.n74 VTAIL.n73 0.155672
R2282 VTAIL.n74 VTAIL.n11 0.155672
R2283 VTAIL.n81 VTAIL.n11 0.155672
R2284 VTAIL.n82 VTAIL.n81 0.155672
R2285 VTAIL.n82 VTAIL.n7 0.155672
R2286 VTAIL.n89 VTAIL.n7 0.155672
R2287 VTAIL.n90 VTAIL.n89 0.155672
R2288 VTAIL.n90 VTAIL.n3 0.155672
R2289 VTAIL.n97 VTAIL.n3 0.155672
R2290 VTAIL.n98 VTAIL.n97 0.155672
R2291 VTAIL.n143 VTAIL.n135 0.155672
R2292 VTAIL.n144 VTAIL.n143 0.155672
R2293 VTAIL.n144 VTAIL.n131 0.155672
R2294 VTAIL.n151 VTAIL.n131 0.155672
R2295 VTAIL.n152 VTAIL.n151 0.155672
R2296 VTAIL.n152 VTAIL.n127 0.155672
R2297 VTAIL.n161 VTAIL.n127 0.155672
R2298 VTAIL.n162 VTAIL.n161 0.155672
R2299 VTAIL.n162 VTAIL.n123 0.155672
R2300 VTAIL.n169 VTAIL.n123 0.155672
R2301 VTAIL.n170 VTAIL.n169 0.155672
R2302 VTAIL.n170 VTAIL.n119 0.155672
R2303 VTAIL.n177 VTAIL.n119 0.155672
R2304 VTAIL.n178 VTAIL.n177 0.155672
R2305 VTAIL.n178 VTAIL.n115 0.155672
R2306 VTAIL.n185 VTAIL.n115 0.155672
R2307 VTAIL.n186 VTAIL.n185 0.155672
R2308 VTAIL.n186 VTAIL.n111 0.155672
R2309 VTAIL.n193 VTAIL.n111 0.155672
R2310 VTAIL.n194 VTAIL.n193 0.155672
R2311 VTAIL.n194 VTAIL.n107 0.155672
R2312 VTAIL.n201 VTAIL.n107 0.155672
R2313 VTAIL.n202 VTAIL.n201 0.155672
R2314 VTAIL.n247 VTAIL.n239 0.155672
R2315 VTAIL.n248 VTAIL.n247 0.155672
R2316 VTAIL.n248 VTAIL.n235 0.155672
R2317 VTAIL.n255 VTAIL.n235 0.155672
R2318 VTAIL.n256 VTAIL.n255 0.155672
R2319 VTAIL.n256 VTAIL.n231 0.155672
R2320 VTAIL.n265 VTAIL.n231 0.155672
R2321 VTAIL.n266 VTAIL.n265 0.155672
R2322 VTAIL.n266 VTAIL.n227 0.155672
R2323 VTAIL.n273 VTAIL.n227 0.155672
R2324 VTAIL.n274 VTAIL.n273 0.155672
R2325 VTAIL.n274 VTAIL.n223 0.155672
R2326 VTAIL.n281 VTAIL.n223 0.155672
R2327 VTAIL.n282 VTAIL.n281 0.155672
R2328 VTAIL.n282 VTAIL.n219 0.155672
R2329 VTAIL.n289 VTAIL.n219 0.155672
R2330 VTAIL.n290 VTAIL.n289 0.155672
R2331 VTAIL.n290 VTAIL.n215 0.155672
R2332 VTAIL.n297 VTAIL.n215 0.155672
R2333 VTAIL.n298 VTAIL.n297 0.155672
R2334 VTAIL.n298 VTAIL.n211 0.155672
R2335 VTAIL.n305 VTAIL.n211 0.155672
R2336 VTAIL.n306 VTAIL.n305 0.155672
R2337 VTAIL.n722 VTAIL.n721 0.155672
R2338 VTAIL.n721 VTAIL.n627 0.155672
R2339 VTAIL.n714 VTAIL.n627 0.155672
R2340 VTAIL.n714 VTAIL.n713 0.155672
R2341 VTAIL.n713 VTAIL.n631 0.155672
R2342 VTAIL.n706 VTAIL.n631 0.155672
R2343 VTAIL.n706 VTAIL.n705 0.155672
R2344 VTAIL.n705 VTAIL.n635 0.155672
R2345 VTAIL.n698 VTAIL.n635 0.155672
R2346 VTAIL.n698 VTAIL.n697 0.155672
R2347 VTAIL.n697 VTAIL.n639 0.155672
R2348 VTAIL.n690 VTAIL.n639 0.155672
R2349 VTAIL.n690 VTAIL.n689 0.155672
R2350 VTAIL.n689 VTAIL.n643 0.155672
R2351 VTAIL.n682 VTAIL.n643 0.155672
R2352 VTAIL.n682 VTAIL.n681 0.155672
R2353 VTAIL.n681 VTAIL.n647 0.155672
R2354 VTAIL.n674 VTAIL.n647 0.155672
R2355 VTAIL.n674 VTAIL.n673 0.155672
R2356 VTAIL.n673 VTAIL.n653 0.155672
R2357 VTAIL.n666 VTAIL.n653 0.155672
R2358 VTAIL.n666 VTAIL.n665 0.155672
R2359 VTAIL.n665 VTAIL.n657 0.155672
R2360 VTAIL.n618 VTAIL.n617 0.155672
R2361 VTAIL.n617 VTAIL.n523 0.155672
R2362 VTAIL.n610 VTAIL.n523 0.155672
R2363 VTAIL.n610 VTAIL.n609 0.155672
R2364 VTAIL.n609 VTAIL.n527 0.155672
R2365 VTAIL.n602 VTAIL.n527 0.155672
R2366 VTAIL.n602 VTAIL.n601 0.155672
R2367 VTAIL.n601 VTAIL.n531 0.155672
R2368 VTAIL.n594 VTAIL.n531 0.155672
R2369 VTAIL.n594 VTAIL.n593 0.155672
R2370 VTAIL.n593 VTAIL.n535 0.155672
R2371 VTAIL.n586 VTAIL.n535 0.155672
R2372 VTAIL.n586 VTAIL.n585 0.155672
R2373 VTAIL.n585 VTAIL.n539 0.155672
R2374 VTAIL.n578 VTAIL.n539 0.155672
R2375 VTAIL.n578 VTAIL.n577 0.155672
R2376 VTAIL.n577 VTAIL.n543 0.155672
R2377 VTAIL.n570 VTAIL.n543 0.155672
R2378 VTAIL.n570 VTAIL.n569 0.155672
R2379 VTAIL.n569 VTAIL.n549 0.155672
R2380 VTAIL.n562 VTAIL.n549 0.155672
R2381 VTAIL.n562 VTAIL.n561 0.155672
R2382 VTAIL.n561 VTAIL.n553 0.155672
R2383 VTAIL.n514 VTAIL.n513 0.155672
R2384 VTAIL.n513 VTAIL.n419 0.155672
R2385 VTAIL.n506 VTAIL.n419 0.155672
R2386 VTAIL.n506 VTAIL.n505 0.155672
R2387 VTAIL.n505 VTAIL.n423 0.155672
R2388 VTAIL.n498 VTAIL.n423 0.155672
R2389 VTAIL.n498 VTAIL.n497 0.155672
R2390 VTAIL.n497 VTAIL.n427 0.155672
R2391 VTAIL.n490 VTAIL.n427 0.155672
R2392 VTAIL.n490 VTAIL.n489 0.155672
R2393 VTAIL.n489 VTAIL.n431 0.155672
R2394 VTAIL.n482 VTAIL.n431 0.155672
R2395 VTAIL.n482 VTAIL.n481 0.155672
R2396 VTAIL.n481 VTAIL.n435 0.155672
R2397 VTAIL.n474 VTAIL.n435 0.155672
R2398 VTAIL.n474 VTAIL.n473 0.155672
R2399 VTAIL.n473 VTAIL.n439 0.155672
R2400 VTAIL.n466 VTAIL.n439 0.155672
R2401 VTAIL.n466 VTAIL.n465 0.155672
R2402 VTAIL.n465 VTAIL.n445 0.155672
R2403 VTAIL.n458 VTAIL.n445 0.155672
R2404 VTAIL.n458 VTAIL.n457 0.155672
R2405 VTAIL.n457 VTAIL.n449 0.155672
R2406 VTAIL.n410 VTAIL.n409 0.155672
R2407 VTAIL.n409 VTAIL.n315 0.155672
R2408 VTAIL.n402 VTAIL.n315 0.155672
R2409 VTAIL.n402 VTAIL.n401 0.155672
R2410 VTAIL.n401 VTAIL.n319 0.155672
R2411 VTAIL.n394 VTAIL.n319 0.155672
R2412 VTAIL.n394 VTAIL.n393 0.155672
R2413 VTAIL.n393 VTAIL.n323 0.155672
R2414 VTAIL.n386 VTAIL.n323 0.155672
R2415 VTAIL.n386 VTAIL.n385 0.155672
R2416 VTAIL.n385 VTAIL.n327 0.155672
R2417 VTAIL.n378 VTAIL.n327 0.155672
R2418 VTAIL.n378 VTAIL.n377 0.155672
R2419 VTAIL.n377 VTAIL.n331 0.155672
R2420 VTAIL.n370 VTAIL.n331 0.155672
R2421 VTAIL.n370 VTAIL.n369 0.155672
R2422 VTAIL.n369 VTAIL.n335 0.155672
R2423 VTAIL.n362 VTAIL.n335 0.155672
R2424 VTAIL.n362 VTAIL.n361 0.155672
R2425 VTAIL.n361 VTAIL.n341 0.155672
R2426 VTAIL.n354 VTAIL.n341 0.155672
R2427 VTAIL.n354 VTAIL.n353 0.155672
R2428 VTAIL.n353 VTAIL.n345 0.155672
R2429 VP.n2 VP.t3 271.589
R2430 VP.n2 VP.t0 271.07
R2431 VP.n4 VP.t2 236.458
R2432 VP.n11 VP.t1 236.458
R2433 VP.n10 VP.n0 161.3
R2434 VP.n9 VP.n8 161.3
R2435 VP.n7 VP.n1 161.3
R2436 VP.n6 VP.n5 161.3
R2437 VP.n4 VP.n3 92.7103
R2438 VP.n12 VP.n11 92.7103
R2439 VP.n3 VP.n2 56.8066
R2440 VP.n9 VP.n1 56.5617
R2441 VP.n5 VP.n1 24.5923
R2442 VP.n10 VP.n9 24.5923
R2443 VP.n5 VP.n4 18.1985
R2444 VP.n11 VP.n10 18.1985
R2445 VP.n6 VP.n3 0.278335
R2446 VP.n12 VP.n0 0.278335
R2447 VP.n7 VP.n6 0.189894
R2448 VP.n8 VP.n7 0.189894
R2449 VP.n8 VP.n0 0.189894
R2450 VP VP.n12 0.153485
R2451 VDD1 VDD1.n1 116.99
R2452 VDD1 VDD1.n0 70.8595
R2453 VDD1.n0 VDD1.t0 1.73502
R2454 VDD1.n0 VDD1.t3 1.73502
R2455 VDD1.n1 VDD1.t1 1.73502
R2456 VDD1.n1 VDD1.t2 1.73502
C0 VTAIL VDD2 7.26233f
C1 B w_n2314_n4716# 10.2865f
C2 VN w_n2314_n4716# 3.9227f
C3 B VP 1.54768f
C4 w_n2314_n4716# VDD1 1.50125f
C5 VP VN 6.94259f
C6 w_n2314_n4716# VDD2 1.54193f
C7 VP VDD1 6.98767f
C8 VTAIL w_n2314_n4716# 5.53004f
C9 VP VDD2 0.350857f
C10 VP VTAIL 6.341f
C11 B VN 1.06014f
C12 B VDD1 1.3225f
C13 VN VDD1 0.148834f
C14 B VDD2 1.36335f
C15 B VTAIL 6.71562f
C16 VN VDD2 6.78621f
C17 VN VTAIL 6.32689f
C18 VDD1 VDD2 0.8613f
C19 VP w_n2314_n4716# 4.218431f
C20 VTAIL VDD1 7.21275f
C21 VDD2 VSUBS 0.998586f
C22 VDD1 VSUBS 6.21816f
C23 VTAIL VSUBS 1.465255f
C24 VN VSUBS 5.52201f
C25 VP VSUBS 2.176818f
C26 B VSUBS 4.246814f
C27 w_n2314_n4716# VSUBS 0.13337p
C28 VDD1.t0 VSUBS 0.393268f
C29 VDD1.t3 VSUBS 0.393268f
C30 VDD1.n0 VSUBS 3.30437f
C31 VDD1.t1 VSUBS 0.393268f
C32 VDD1.t2 VSUBS 0.393268f
C33 VDD1.n1 VSUBS 4.25163f
C34 VP.n0 VSUBS 0.047452f
C35 VP.t1 VSUBS 3.54633f
C36 VP.n1 VSUBS 0.052323f
C37 VP.t0 VSUBS 3.72675f
C38 VP.t3 VSUBS 3.72948f
C39 VP.n2 VSUBS 4.443491f
C40 VP.n3 VSUBS 2.2626f
C41 VP.t2 VSUBS 3.54633f
C42 VP.n4 VSUBS 1.33782f
C43 VP.n5 VSUBS 0.05818f
C44 VP.n6 VSUBS 0.047452f
C45 VP.n7 VSUBS 0.035994f
C46 VP.n8 VSUBS 0.035994f
C47 VP.n9 VSUBS 0.052323f
C48 VP.n10 VSUBS 0.05818f
C49 VP.n11 VSUBS 1.33782f
C50 VP.n12 VSUBS 0.044756f
C51 VTAIL.n0 VSUBS 0.012258f
C52 VTAIL.n1 VSUBS 0.027683f
C53 VTAIL.n2 VSUBS 0.012401f
C54 VTAIL.n3 VSUBS 0.021795f
C55 VTAIL.n4 VSUBS 0.011712f
C56 VTAIL.n5 VSUBS 0.027683f
C57 VTAIL.n6 VSUBS 0.012401f
C58 VTAIL.n7 VSUBS 0.021795f
C59 VTAIL.n8 VSUBS 0.011712f
C60 VTAIL.n9 VSUBS 0.027683f
C61 VTAIL.n10 VSUBS 0.012401f
C62 VTAIL.n11 VSUBS 0.021795f
C63 VTAIL.n12 VSUBS 0.011712f
C64 VTAIL.n13 VSUBS 0.027683f
C65 VTAIL.n14 VSUBS 0.012401f
C66 VTAIL.n15 VSUBS 0.021795f
C67 VTAIL.n16 VSUBS 0.011712f
C68 VTAIL.n17 VSUBS 0.027683f
C69 VTAIL.n18 VSUBS 0.012401f
C70 VTAIL.n19 VSUBS 0.021795f
C71 VTAIL.n20 VSUBS 0.011712f
C72 VTAIL.n21 VSUBS 0.027683f
C73 VTAIL.n22 VSUBS 0.012056f
C74 VTAIL.n23 VSUBS 0.021795f
C75 VTAIL.n24 VSUBS 0.012401f
C76 VTAIL.n25 VSUBS 0.027683f
C77 VTAIL.n26 VSUBS 0.012401f
C78 VTAIL.n27 VSUBS 0.021795f
C79 VTAIL.n28 VSUBS 0.011712f
C80 VTAIL.n29 VSUBS 0.027683f
C81 VTAIL.n30 VSUBS 0.012401f
C82 VTAIL.n31 VSUBS 1.71454f
C83 VTAIL.n32 VSUBS 0.011712f
C84 VTAIL.t7 VSUBS 0.060149f
C85 VTAIL.n33 VSUBS 0.238073f
C86 VTAIL.n34 VSUBS 0.020824f
C87 VTAIL.n35 VSUBS 0.020762f
C88 VTAIL.n36 VSUBS 0.027683f
C89 VTAIL.n37 VSUBS 0.012401f
C90 VTAIL.n38 VSUBS 0.011712f
C91 VTAIL.n39 VSUBS 0.021795f
C92 VTAIL.n40 VSUBS 0.021795f
C93 VTAIL.n41 VSUBS 0.011712f
C94 VTAIL.n42 VSUBS 0.012401f
C95 VTAIL.n43 VSUBS 0.027683f
C96 VTAIL.n44 VSUBS 0.027683f
C97 VTAIL.n45 VSUBS 0.012401f
C98 VTAIL.n46 VSUBS 0.011712f
C99 VTAIL.n47 VSUBS 0.021795f
C100 VTAIL.n48 VSUBS 0.021795f
C101 VTAIL.n49 VSUBS 0.011712f
C102 VTAIL.n50 VSUBS 0.011712f
C103 VTAIL.n51 VSUBS 0.012401f
C104 VTAIL.n52 VSUBS 0.027683f
C105 VTAIL.n53 VSUBS 0.027683f
C106 VTAIL.n54 VSUBS 0.027683f
C107 VTAIL.n55 VSUBS 0.012056f
C108 VTAIL.n56 VSUBS 0.011712f
C109 VTAIL.n57 VSUBS 0.021795f
C110 VTAIL.n58 VSUBS 0.021795f
C111 VTAIL.n59 VSUBS 0.011712f
C112 VTAIL.n60 VSUBS 0.012401f
C113 VTAIL.n61 VSUBS 0.027683f
C114 VTAIL.n62 VSUBS 0.027683f
C115 VTAIL.n63 VSUBS 0.012401f
C116 VTAIL.n64 VSUBS 0.011712f
C117 VTAIL.n65 VSUBS 0.021795f
C118 VTAIL.n66 VSUBS 0.021795f
C119 VTAIL.n67 VSUBS 0.011712f
C120 VTAIL.n68 VSUBS 0.012401f
C121 VTAIL.n69 VSUBS 0.027683f
C122 VTAIL.n70 VSUBS 0.027683f
C123 VTAIL.n71 VSUBS 0.012401f
C124 VTAIL.n72 VSUBS 0.011712f
C125 VTAIL.n73 VSUBS 0.021795f
C126 VTAIL.n74 VSUBS 0.021795f
C127 VTAIL.n75 VSUBS 0.011712f
C128 VTAIL.n76 VSUBS 0.012401f
C129 VTAIL.n77 VSUBS 0.027683f
C130 VTAIL.n78 VSUBS 0.027683f
C131 VTAIL.n79 VSUBS 0.012401f
C132 VTAIL.n80 VSUBS 0.011712f
C133 VTAIL.n81 VSUBS 0.021795f
C134 VTAIL.n82 VSUBS 0.021795f
C135 VTAIL.n83 VSUBS 0.011712f
C136 VTAIL.n84 VSUBS 0.012401f
C137 VTAIL.n85 VSUBS 0.027683f
C138 VTAIL.n86 VSUBS 0.027683f
C139 VTAIL.n87 VSUBS 0.012401f
C140 VTAIL.n88 VSUBS 0.011712f
C141 VTAIL.n89 VSUBS 0.021795f
C142 VTAIL.n90 VSUBS 0.021795f
C143 VTAIL.n91 VSUBS 0.011712f
C144 VTAIL.n92 VSUBS 0.012401f
C145 VTAIL.n93 VSUBS 0.027683f
C146 VTAIL.n94 VSUBS 0.027683f
C147 VTAIL.n95 VSUBS 0.012401f
C148 VTAIL.n96 VSUBS 0.011712f
C149 VTAIL.n97 VSUBS 0.021795f
C150 VTAIL.n98 VSUBS 0.054547f
C151 VTAIL.n99 VSUBS 0.011712f
C152 VTAIL.n100 VSUBS 0.012401f
C153 VTAIL.n101 VSUBS 0.061041f
C154 VTAIL.n102 VSUBS 0.04014f
C155 VTAIL.n103 VSUBS 0.125525f
C156 VTAIL.n104 VSUBS 0.012258f
C157 VTAIL.n105 VSUBS 0.027683f
C158 VTAIL.n106 VSUBS 0.012401f
C159 VTAIL.n107 VSUBS 0.021795f
C160 VTAIL.n108 VSUBS 0.011712f
C161 VTAIL.n109 VSUBS 0.027683f
C162 VTAIL.n110 VSUBS 0.012401f
C163 VTAIL.n111 VSUBS 0.021795f
C164 VTAIL.n112 VSUBS 0.011712f
C165 VTAIL.n113 VSUBS 0.027683f
C166 VTAIL.n114 VSUBS 0.012401f
C167 VTAIL.n115 VSUBS 0.021795f
C168 VTAIL.n116 VSUBS 0.011712f
C169 VTAIL.n117 VSUBS 0.027683f
C170 VTAIL.n118 VSUBS 0.012401f
C171 VTAIL.n119 VSUBS 0.021795f
C172 VTAIL.n120 VSUBS 0.011712f
C173 VTAIL.n121 VSUBS 0.027683f
C174 VTAIL.n122 VSUBS 0.012401f
C175 VTAIL.n123 VSUBS 0.021795f
C176 VTAIL.n124 VSUBS 0.011712f
C177 VTAIL.n125 VSUBS 0.027683f
C178 VTAIL.n126 VSUBS 0.012056f
C179 VTAIL.n127 VSUBS 0.021795f
C180 VTAIL.n128 VSUBS 0.012401f
C181 VTAIL.n129 VSUBS 0.027683f
C182 VTAIL.n130 VSUBS 0.012401f
C183 VTAIL.n131 VSUBS 0.021795f
C184 VTAIL.n132 VSUBS 0.011712f
C185 VTAIL.n133 VSUBS 0.027683f
C186 VTAIL.n134 VSUBS 0.012401f
C187 VTAIL.n135 VSUBS 1.71454f
C188 VTAIL.n136 VSUBS 0.011712f
C189 VTAIL.t3 VSUBS 0.060149f
C190 VTAIL.n137 VSUBS 0.238073f
C191 VTAIL.n138 VSUBS 0.020824f
C192 VTAIL.n139 VSUBS 0.020762f
C193 VTAIL.n140 VSUBS 0.027683f
C194 VTAIL.n141 VSUBS 0.012401f
C195 VTAIL.n142 VSUBS 0.011712f
C196 VTAIL.n143 VSUBS 0.021795f
C197 VTAIL.n144 VSUBS 0.021795f
C198 VTAIL.n145 VSUBS 0.011712f
C199 VTAIL.n146 VSUBS 0.012401f
C200 VTAIL.n147 VSUBS 0.027683f
C201 VTAIL.n148 VSUBS 0.027683f
C202 VTAIL.n149 VSUBS 0.012401f
C203 VTAIL.n150 VSUBS 0.011712f
C204 VTAIL.n151 VSUBS 0.021795f
C205 VTAIL.n152 VSUBS 0.021795f
C206 VTAIL.n153 VSUBS 0.011712f
C207 VTAIL.n154 VSUBS 0.011712f
C208 VTAIL.n155 VSUBS 0.012401f
C209 VTAIL.n156 VSUBS 0.027683f
C210 VTAIL.n157 VSUBS 0.027683f
C211 VTAIL.n158 VSUBS 0.027683f
C212 VTAIL.n159 VSUBS 0.012056f
C213 VTAIL.n160 VSUBS 0.011712f
C214 VTAIL.n161 VSUBS 0.021795f
C215 VTAIL.n162 VSUBS 0.021795f
C216 VTAIL.n163 VSUBS 0.011712f
C217 VTAIL.n164 VSUBS 0.012401f
C218 VTAIL.n165 VSUBS 0.027683f
C219 VTAIL.n166 VSUBS 0.027683f
C220 VTAIL.n167 VSUBS 0.012401f
C221 VTAIL.n168 VSUBS 0.011712f
C222 VTAIL.n169 VSUBS 0.021795f
C223 VTAIL.n170 VSUBS 0.021795f
C224 VTAIL.n171 VSUBS 0.011712f
C225 VTAIL.n172 VSUBS 0.012401f
C226 VTAIL.n173 VSUBS 0.027683f
C227 VTAIL.n174 VSUBS 0.027683f
C228 VTAIL.n175 VSUBS 0.012401f
C229 VTAIL.n176 VSUBS 0.011712f
C230 VTAIL.n177 VSUBS 0.021795f
C231 VTAIL.n178 VSUBS 0.021795f
C232 VTAIL.n179 VSUBS 0.011712f
C233 VTAIL.n180 VSUBS 0.012401f
C234 VTAIL.n181 VSUBS 0.027683f
C235 VTAIL.n182 VSUBS 0.027683f
C236 VTAIL.n183 VSUBS 0.012401f
C237 VTAIL.n184 VSUBS 0.011712f
C238 VTAIL.n185 VSUBS 0.021795f
C239 VTAIL.n186 VSUBS 0.021795f
C240 VTAIL.n187 VSUBS 0.011712f
C241 VTAIL.n188 VSUBS 0.012401f
C242 VTAIL.n189 VSUBS 0.027683f
C243 VTAIL.n190 VSUBS 0.027683f
C244 VTAIL.n191 VSUBS 0.012401f
C245 VTAIL.n192 VSUBS 0.011712f
C246 VTAIL.n193 VSUBS 0.021795f
C247 VTAIL.n194 VSUBS 0.021795f
C248 VTAIL.n195 VSUBS 0.011712f
C249 VTAIL.n196 VSUBS 0.012401f
C250 VTAIL.n197 VSUBS 0.027683f
C251 VTAIL.n198 VSUBS 0.027683f
C252 VTAIL.n199 VSUBS 0.012401f
C253 VTAIL.n200 VSUBS 0.011712f
C254 VTAIL.n201 VSUBS 0.021795f
C255 VTAIL.n202 VSUBS 0.054547f
C256 VTAIL.n203 VSUBS 0.011712f
C257 VTAIL.n204 VSUBS 0.012401f
C258 VTAIL.n205 VSUBS 0.061041f
C259 VTAIL.n206 VSUBS 0.04014f
C260 VTAIL.n207 VSUBS 0.189246f
C261 VTAIL.n208 VSUBS 0.012258f
C262 VTAIL.n209 VSUBS 0.027683f
C263 VTAIL.n210 VSUBS 0.012401f
C264 VTAIL.n211 VSUBS 0.021795f
C265 VTAIL.n212 VSUBS 0.011712f
C266 VTAIL.n213 VSUBS 0.027683f
C267 VTAIL.n214 VSUBS 0.012401f
C268 VTAIL.n215 VSUBS 0.021795f
C269 VTAIL.n216 VSUBS 0.011712f
C270 VTAIL.n217 VSUBS 0.027683f
C271 VTAIL.n218 VSUBS 0.012401f
C272 VTAIL.n219 VSUBS 0.021795f
C273 VTAIL.n220 VSUBS 0.011712f
C274 VTAIL.n221 VSUBS 0.027683f
C275 VTAIL.n222 VSUBS 0.012401f
C276 VTAIL.n223 VSUBS 0.021795f
C277 VTAIL.n224 VSUBS 0.011712f
C278 VTAIL.n225 VSUBS 0.027683f
C279 VTAIL.n226 VSUBS 0.012401f
C280 VTAIL.n227 VSUBS 0.021795f
C281 VTAIL.n228 VSUBS 0.011712f
C282 VTAIL.n229 VSUBS 0.027683f
C283 VTAIL.n230 VSUBS 0.012056f
C284 VTAIL.n231 VSUBS 0.021795f
C285 VTAIL.n232 VSUBS 0.012401f
C286 VTAIL.n233 VSUBS 0.027683f
C287 VTAIL.n234 VSUBS 0.012401f
C288 VTAIL.n235 VSUBS 0.021795f
C289 VTAIL.n236 VSUBS 0.011712f
C290 VTAIL.n237 VSUBS 0.027683f
C291 VTAIL.n238 VSUBS 0.012401f
C292 VTAIL.n239 VSUBS 1.71454f
C293 VTAIL.n240 VSUBS 0.011712f
C294 VTAIL.t0 VSUBS 0.060149f
C295 VTAIL.n241 VSUBS 0.238073f
C296 VTAIL.n242 VSUBS 0.020824f
C297 VTAIL.n243 VSUBS 0.020762f
C298 VTAIL.n244 VSUBS 0.027683f
C299 VTAIL.n245 VSUBS 0.012401f
C300 VTAIL.n246 VSUBS 0.011712f
C301 VTAIL.n247 VSUBS 0.021795f
C302 VTAIL.n248 VSUBS 0.021795f
C303 VTAIL.n249 VSUBS 0.011712f
C304 VTAIL.n250 VSUBS 0.012401f
C305 VTAIL.n251 VSUBS 0.027683f
C306 VTAIL.n252 VSUBS 0.027683f
C307 VTAIL.n253 VSUBS 0.012401f
C308 VTAIL.n254 VSUBS 0.011712f
C309 VTAIL.n255 VSUBS 0.021795f
C310 VTAIL.n256 VSUBS 0.021795f
C311 VTAIL.n257 VSUBS 0.011712f
C312 VTAIL.n258 VSUBS 0.011712f
C313 VTAIL.n259 VSUBS 0.012401f
C314 VTAIL.n260 VSUBS 0.027683f
C315 VTAIL.n261 VSUBS 0.027683f
C316 VTAIL.n262 VSUBS 0.027683f
C317 VTAIL.n263 VSUBS 0.012056f
C318 VTAIL.n264 VSUBS 0.011712f
C319 VTAIL.n265 VSUBS 0.021795f
C320 VTAIL.n266 VSUBS 0.021795f
C321 VTAIL.n267 VSUBS 0.011712f
C322 VTAIL.n268 VSUBS 0.012401f
C323 VTAIL.n269 VSUBS 0.027683f
C324 VTAIL.n270 VSUBS 0.027683f
C325 VTAIL.n271 VSUBS 0.012401f
C326 VTAIL.n272 VSUBS 0.011712f
C327 VTAIL.n273 VSUBS 0.021795f
C328 VTAIL.n274 VSUBS 0.021795f
C329 VTAIL.n275 VSUBS 0.011712f
C330 VTAIL.n276 VSUBS 0.012401f
C331 VTAIL.n277 VSUBS 0.027683f
C332 VTAIL.n278 VSUBS 0.027683f
C333 VTAIL.n279 VSUBS 0.012401f
C334 VTAIL.n280 VSUBS 0.011712f
C335 VTAIL.n281 VSUBS 0.021795f
C336 VTAIL.n282 VSUBS 0.021795f
C337 VTAIL.n283 VSUBS 0.011712f
C338 VTAIL.n284 VSUBS 0.012401f
C339 VTAIL.n285 VSUBS 0.027683f
C340 VTAIL.n286 VSUBS 0.027683f
C341 VTAIL.n287 VSUBS 0.012401f
C342 VTAIL.n288 VSUBS 0.011712f
C343 VTAIL.n289 VSUBS 0.021795f
C344 VTAIL.n290 VSUBS 0.021795f
C345 VTAIL.n291 VSUBS 0.011712f
C346 VTAIL.n292 VSUBS 0.012401f
C347 VTAIL.n293 VSUBS 0.027683f
C348 VTAIL.n294 VSUBS 0.027683f
C349 VTAIL.n295 VSUBS 0.012401f
C350 VTAIL.n296 VSUBS 0.011712f
C351 VTAIL.n297 VSUBS 0.021795f
C352 VTAIL.n298 VSUBS 0.021795f
C353 VTAIL.n299 VSUBS 0.011712f
C354 VTAIL.n300 VSUBS 0.012401f
C355 VTAIL.n301 VSUBS 0.027683f
C356 VTAIL.n302 VSUBS 0.027683f
C357 VTAIL.n303 VSUBS 0.012401f
C358 VTAIL.n304 VSUBS 0.011712f
C359 VTAIL.n305 VSUBS 0.021795f
C360 VTAIL.n306 VSUBS 0.054547f
C361 VTAIL.n307 VSUBS 0.011712f
C362 VTAIL.n308 VSUBS 0.012401f
C363 VTAIL.n309 VSUBS 0.061041f
C364 VTAIL.n310 VSUBS 0.04014f
C365 VTAIL.n311 VSUBS 1.7225f
C366 VTAIL.n312 VSUBS 0.012258f
C367 VTAIL.n313 VSUBS 0.027683f
C368 VTAIL.n314 VSUBS 0.012401f
C369 VTAIL.n315 VSUBS 0.021795f
C370 VTAIL.n316 VSUBS 0.011712f
C371 VTAIL.n317 VSUBS 0.027683f
C372 VTAIL.n318 VSUBS 0.012401f
C373 VTAIL.n319 VSUBS 0.021795f
C374 VTAIL.n320 VSUBS 0.011712f
C375 VTAIL.n321 VSUBS 0.027683f
C376 VTAIL.n322 VSUBS 0.012401f
C377 VTAIL.n323 VSUBS 0.021795f
C378 VTAIL.n324 VSUBS 0.011712f
C379 VTAIL.n325 VSUBS 0.027683f
C380 VTAIL.n326 VSUBS 0.012401f
C381 VTAIL.n327 VSUBS 0.021795f
C382 VTAIL.n328 VSUBS 0.011712f
C383 VTAIL.n329 VSUBS 0.027683f
C384 VTAIL.n330 VSUBS 0.012401f
C385 VTAIL.n331 VSUBS 0.021795f
C386 VTAIL.n332 VSUBS 0.011712f
C387 VTAIL.n333 VSUBS 0.027683f
C388 VTAIL.n334 VSUBS 0.012056f
C389 VTAIL.n335 VSUBS 0.021795f
C390 VTAIL.n336 VSUBS 0.012056f
C391 VTAIL.n337 VSUBS 0.011712f
C392 VTAIL.n338 VSUBS 0.027683f
C393 VTAIL.n339 VSUBS 0.027683f
C394 VTAIL.n340 VSUBS 0.012401f
C395 VTAIL.n341 VSUBS 0.021795f
C396 VTAIL.n342 VSUBS 0.011712f
C397 VTAIL.n343 VSUBS 0.027683f
C398 VTAIL.n344 VSUBS 0.012401f
C399 VTAIL.n345 VSUBS 1.71454f
C400 VTAIL.n346 VSUBS 0.011712f
C401 VTAIL.t4 VSUBS 0.060149f
C402 VTAIL.n347 VSUBS 0.238073f
C403 VTAIL.n348 VSUBS 0.020824f
C404 VTAIL.n349 VSUBS 0.020762f
C405 VTAIL.n350 VSUBS 0.027683f
C406 VTAIL.n351 VSUBS 0.012401f
C407 VTAIL.n352 VSUBS 0.011712f
C408 VTAIL.n353 VSUBS 0.021795f
C409 VTAIL.n354 VSUBS 0.021795f
C410 VTAIL.n355 VSUBS 0.011712f
C411 VTAIL.n356 VSUBS 0.012401f
C412 VTAIL.n357 VSUBS 0.027683f
C413 VTAIL.n358 VSUBS 0.027683f
C414 VTAIL.n359 VSUBS 0.012401f
C415 VTAIL.n360 VSUBS 0.011712f
C416 VTAIL.n361 VSUBS 0.021795f
C417 VTAIL.n362 VSUBS 0.021795f
C418 VTAIL.n363 VSUBS 0.011712f
C419 VTAIL.n364 VSUBS 0.012401f
C420 VTAIL.n365 VSUBS 0.027683f
C421 VTAIL.n366 VSUBS 0.027683f
C422 VTAIL.n367 VSUBS 0.012401f
C423 VTAIL.n368 VSUBS 0.011712f
C424 VTAIL.n369 VSUBS 0.021795f
C425 VTAIL.n370 VSUBS 0.021795f
C426 VTAIL.n371 VSUBS 0.011712f
C427 VTAIL.n372 VSUBS 0.012401f
C428 VTAIL.n373 VSUBS 0.027683f
C429 VTAIL.n374 VSUBS 0.027683f
C430 VTAIL.n375 VSUBS 0.012401f
C431 VTAIL.n376 VSUBS 0.011712f
C432 VTAIL.n377 VSUBS 0.021795f
C433 VTAIL.n378 VSUBS 0.021795f
C434 VTAIL.n379 VSUBS 0.011712f
C435 VTAIL.n380 VSUBS 0.012401f
C436 VTAIL.n381 VSUBS 0.027683f
C437 VTAIL.n382 VSUBS 0.027683f
C438 VTAIL.n383 VSUBS 0.012401f
C439 VTAIL.n384 VSUBS 0.011712f
C440 VTAIL.n385 VSUBS 0.021795f
C441 VTAIL.n386 VSUBS 0.021795f
C442 VTAIL.n387 VSUBS 0.011712f
C443 VTAIL.n388 VSUBS 0.012401f
C444 VTAIL.n389 VSUBS 0.027683f
C445 VTAIL.n390 VSUBS 0.027683f
C446 VTAIL.n391 VSUBS 0.012401f
C447 VTAIL.n392 VSUBS 0.011712f
C448 VTAIL.n393 VSUBS 0.021795f
C449 VTAIL.n394 VSUBS 0.021795f
C450 VTAIL.n395 VSUBS 0.011712f
C451 VTAIL.n396 VSUBS 0.012401f
C452 VTAIL.n397 VSUBS 0.027683f
C453 VTAIL.n398 VSUBS 0.027683f
C454 VTAIL.n399 VSUBS 0.012401f
C455 VTAIL.n400 VSUBS 0.011712f
C456 VTAIL.n401 VSUBS 0.021795f
C457 VTAIL.n402 VSUBS 0.021795f
C458 VTAIL.n403 VSUBS 0.011712f
C459 VTAIL.n404 VSUBS 0.012401f
C460 VTAIL.n405 VSUBS 0.027683f
C461 VTAIL.n406 VSUBS 0.027683f
C462 VTAIL.n407 VSUBS 0.012401f
C463 VTAIL.n408 VSUBS 0.011712f
C464 VTAIL.n409 VSUBS 0.021795f
C465 VTAIL.n410 VSUBS 0.054547f
C466 VTAIL.n411 VSUBS 0.011712f
C467 VTAIL.n412 VSUBS 0.012401f
C468 VTAIL.n413 VSUBS 0.061041f
C469 VTAIL.n414 VSUBS 0.04014f
C470 VTAIL.n415 VSUBS 1.7225f
C471 VTAIL.n416 VSUBS 0.012258f
C472 VTAIL.n417 VSUBS 0.027683f
C473 VTAIL.n418 VSUBS 0.012401f
C474 VTAIL.n419 VSUBS 0.021795f
C475 VTAIL.n420 VSUBS 0.011712f
C476 VTAIL.n421 VSUBS 0.027683f
C477 VTAIL.n422 VSUBS 0.012401f
C478 VTAIL.n423 VSUBS 0.021795f
C479 VTAIL.n424 VSUBS 0.011712f
C480 VTAIL.n425 VSUBS 0.027683f
C481 VTAIL.n426 VSUBS 0.012401f
C482 VTAIL.n427 VSUBS 0.021795f
C483 VTAIL.n428 VSUBS 0.011712f
C484 VTAIL.n429 VSUBS 0.027683f
C485 VTAIL.n430 VSUBS 0.012401f
C486 VTAIL.n431 VSUBS 0.021795f
C487 VTAIL.n432 VSUBS 0.011712f
C488 VTAIL.n433 VSUBS 0.027683f
C489 VTAIL.n434 VSUBS 0.012401f
C490 VTAIL.n435 VSUBS 0.021795f
C491 VTAIL.n436 VSUBS 0.011712f
C492 VTAIL.n437 VSUBS 0.027683f
C493 VTAIL.n438 VSUBS 0.012056f
C494 VTAIL.n439 VSUBS 0.021795f
C495 VTAIL.n440 VSUBS 0.012056f
C496 VTAIL.n441 VSUBS 0.011712f
C497 VTAIL.n442 VSUBS 0.027683f
C498 VTAIL.n443 VSUBS 0.027683f
C499 VTAIL.n444 VSUBS 0.012401f
C500 VTAIL.n445 VSUBS 0.021795f
C501 VTAIL.n446 VSUBS 0.011712f
C502 VTAIL.n447 VSUBS 0.027683f
C503 VTAIL.n448 VSUBS 0.012401f
C504 VTAIL.n449 VSUBS 1.71454f
C505 VTAIL.n450 VSUBS 0.011712f
C506 VTAIL.t5 VSUBS 0.060149f
C507 VTAIL.n451 VSUBS 0.238073f
C508 VTAIL.n452 VSUBS 0.020824f
C509 VTAIL.n453 VSUBS 0.020762f
C510 VTAIL.n454 VSUBS 0.027683f
C511 VTAIL.n455 VSUBS 0.012401f
C512 VTAIL.n456 VSUBS 0.011712f
C513 VTAIL.n457 VSUBS 0.021795f
C514 VTAIL.n458 VSUBS 0.021795f
C515 VTAIL.n459 VSUBS 0.011712f
C516 VTAIL.n460 VSUBS 0.012401f
C517 VTAIL.n461 VSUBS 0.027683f
C518 VTAIL.n462 VSUBS 0.027683f
C519 VTAIL.n463 VSUBS 0.012401f
C520 VTAIL.n464 VSUBS 0.011712f
C521 VTAIL.n465 VSUBS 0.021795f
C522 VTAIL.n466 VSUBS 0.021795f
C523 VTAIL.n467 VSUBS 0.011712f
C524 VTAIL.n468 VSUBS 0.012401f
C525 VTAIL.n469 VSUBS 0.027683f
C526 VTAIL.n470 VSUBS 0.027683f
C527 VTAIL.n471 VSUBS 0.012401f
C528 VTAIL.n472 VSUBS 0.011712f
C529 VTAIL.n473 VSUBS 0.021795f
C530 VTAIL.n474 VSUBS 0.021795f
C531 VTAIL.n475 VSUBS 0.011712f
C532 VTAIL.n476 VSUBS 0.012401f
C533 VTAIL.n477 VSUBS 0.027683f
C534 VTAIL.n478 VSUBS 0.027683f
C535 VTAIL.n479 VSUBS 0.012401f
C536 VTAIL.n480 VSUBS 0.011712f
C537 VTAIL.n481 VSUBS 0.021795f
C538 VTAIL.n482 VSUBS 0.021795f
C539 VTAIL.n483 VSUBS 0.011712f
C540 VTAIL.n484 VSUBS 0.012401f
C541 VTAIL.n485 VSUBS 0.027683f
C542 VTAIL.n486 VSUBS 0.027683f
C543 VTAIL.n487 VSUBS 0.012401f
C544 VTAIL.n488 VSUBS 0.011712f
C545 VTAIL.n489 VSUBS 0.021795f
C546 VTAIL.n490 VSUBS 0.021795f
C547 VTAIL.n491 VSUBS 0.011712f
C548 VTAIL.n492 VSUBS 0.012401f
C549 VTAIL.n493 VSUBS 0.027683f
C550 VTAIL.n494 VSUBS 0.027683f
C551 VTAIL.n495 VSUBS 0.012401f
C552 VTAIL.n496 VSUBS 0.011712f
C553 VTAIL.n497 VSUBS 0.021795f
C554 VTAIL.n498 VSUBS 0.021795f
C555 VTAIL.n499 VSUBS 0.011712f
C556 VTAIL.n500 VSUBS 0.012401f
C557 VTAIL.n501 VSUBS 0.027683f
C558 VTAIL.n502 VSUBS 0.027683f
C559 VTAIL.n503 VSUBS 0.012401f
C560 VTAIL.n504 VSUBS 0.011712f
C561 VTAIL.n505 VSUBS 0.021795f
C562 VTAIL.n506 VSUBS 0.021795f
C563 VTAIL.n507 VSUBS 0.011712f
C564 VTAIL.n508 VSUBS 0.012401f
C565 VTAIL.n509 VSUBS 0.027683f
C566 VTAIL.n510 VSUBS 0.027683f
C567 VTAIL.n511 VSUBS 0.012401f
C568 VTAIL.n512 VSUBS 0.011712f
C569 VTAIL.n513 VSUBS 0.021795f
C570 VTAIL.n514 VSUBS 0.054547f
C571 VTAIL.n515 VSUBS 0.011712f
C572 VTAIL.n516 VSUBS 0.012401f
C573 VTAIL.n517 VSUBS 0.061041f
C574 VTAIL.n518 VSUBS 0.04014f
C575 VTAIL.n519 VSUBS 0.189246f
C576 VTAIL.n520 VSUBS 0.012258f
C577 VTAIL.n521 VSUBS 0.027683f
C578 VTAIL.n522 VSUBS 0.012401f
C579 VTAIL.n523 VSUBS 0.021795f
C580 VTAIL.n524 VSUBS 0.011712f
C581 VTAIL.n525 VSUBS 0.027683f
C582 VTAIL.n526 VSUBS 0.012401f
C583 VTAIL.n527 VSUBS 0.021795f
C584 VTAIL.n528 VSUBS 0.011712f
C585 VTAIL.n529 VSUBS 0.027683f
C586 VTAIL.n530 VSUBS 0.012401f
C587 VTAIL.n531 VSUBS 0.021795f
C588 VTAIL.n532 VSUBS 0.011712f
C589 VTAIL.n533 VSUBS 0.027683f
C590 VTAIL.n534 VSUBS 0.012401f
C591 VTAIL.n535 VSUBS 0.021795f
C592 VTAIL.n536 VSUBS 0.011712f
C593 VTAIL.n537 VSUBS 0.027683f
C594 VTAIL.n538 VSUBS 0.012401f
C595 VTAIL.n539 VSUBS 0.021795f
C596 VTAIL.n540 VSUBS 0.011712f
C597 VTAIL.n541 VSUBS 0.027683f
C598 VTAIL.n542 VSUBS 0.012056f
C599 VTAIL.n543 VSUBS 0.021795f
C600 VTAIL.n544 VSUBS 0.012056f
C601 VTAIL.n545 VSUBS 0.011712f
C602 VTAIL.n546 VSUBS 0.027683f
C603 VTAIL.n547 VSUBS 0.027683f
C604 VTAIL.n548 VSUBS 0.012401f
C605 VTAIL.n549 VSUBS 0.021795f
C606 VTAIL.n550 VSUBS 0.011712f
C607 VTAIL.n551 VSUBS 0.027683f
C608 VTAIL.n552 VSUBS 0.012401f
C609 VTAIL.n553 VSUBS 1.71454f
C610 VTAIL.n554 VSUBS 0.011712f
C611 VTAIL.t2 VSUBS 0.060149f
C612 VTAIL.n555 VSUBS 0.238073f
C613 VTAIL.n556 VSUBS 0.020824f
C614 VTAIL.n557 VSUBS 0.020762f
C615 VTAIL.n558 VSUBS 0.027683f
C616 VTAIL.n559 VSUBS 0.012401f
C617 VTAIL.n560 VSUBS 0.011712f
C618 VTAIL.n561 VSUBS 0.021795f
C619 VTAIL.n562 VSUBS 0.021795f
C620 VTAIL.n563 VSUBS 0.011712f
C621 VTAIL.n564 VSUBS 0.012401f
C622 VTAIL.n565 VSUBS 0.027683f
C623 VTAIL.n566 VSUBS 0.027683f
C624 VTAIL.n567 VSUBS 0.012401f
C625 VTAIL.n568 VSUBS 0.011712f
C626 VTAIL.n569 VSUBS 0.021795f
C627 VTAIL.n570 VSUBS 0.021795f
C628 VTAIL.n571 VSUBS 0.011712f
C629 VTAIL.n572 VSUBS 0.012401f
C630 VTAIL.n573 VSUBS 0.027683f
C631 VTAIL.n574 VSUBS 0.027683f
C632 VTAIL.n575 VSUBS 0.012401f
C633 VTAIL.n576 VSUBS 0.011712f
C634 VTAIL.n577 VSUBS 0.021795f
C635 VTAIL.n578 VSUBS 0.021795f
C636 VTAIL.n579 VSUBS 0.011712f
C637 VTAIL.n580 VSUBS 0.012401f
C638 VTAIL.n581 VSUBS 0.027683f
C639 VTAIL.n582 VSUBS 0.027683f
C640 VTAIL.n583 VSUBS 0.012401f
C641 VTAIL.n584 VSUBS 0.011712f
C642 VTAIL.n585 VSUBS 0.021795f
C643 VTAIL.n586 VSUBS 0.021795f
C644 VTAIL.n587 VSUBS 0.011712f
C645 VTAIL.n588 VSUBS 0.012401f
C646 VTAIL.n589 VSUBS 0.027683f
C647 VTAIL.n590 VSUBS 0.027683f
C648 VTAIL.n591 VSUBS 0.012401f
C649 VTAIL.n592 VSUBS 0.011712f
C650 VTAIL.n593 VSUBS 0.021795f
C651 VTAIL.n594 VSUBS 0.021795f
C652 VTAIL.n595 VSUBS 0.011712f
C653 VTAIL.n596 VSUBS 0.012401f
C654 VTAIL.n597 VSUBS 0.027683f
C655 VTAIL.n598 VSUBS 0.027683f
C656 VTAIL.n599 VSUBS 0.012401f
C657 VTAIL.n600 VSUBS 0.011712f
C658 VTAIL.n601 VSUBS 0.021795f
C659 VTAIL.n602 VSUBS 0.021795f
C660 VTAIL.n603 VSUBS 0.011712f
C661 VTAIL.n604 VSUBS 0.012401f
C662 VTAIL.n605 VSUBS 0.027683f
C663 VTAIL.n606 VSUBS 0.027683f
C664 VTAIL.n607 VSUBS 0.012401f
C665 VTAIL.n608 VSUBS 0.011712f
C666 VTAIL.n609 VSUBS 0.021795f
C667 VTAIL.n610 VSUBS 0.021795f
C668 VTAIL.n611 VSUBS 0.011712f
C669 VTAIL.n612 VSUBS 0.012401f
C670 VTAIL.n613 VSUBS 0.027683f
C671 VTAIL.n614 VSUBS 0.027683f
C672 VTAIL.n615 VSUBS 0.012401f
C673 VTAIL.n616 VSUBS 0.011712f
C674 VTAIL.n617 VSUBS 0.021795f
C675 VTAIL.n618 VSUBS 0.054547f
C676 VTAIL.n619 VSUBS 0.011712f
C677 VTAIL.n620 VSUBS 0.012401f
C678 VTAIL.n621 VSUBS 0.061041f
C679 VTAIL.n622 VSUBS 0.04014f
C680 VTAIL.n623 VSUBS 0.189246f
C681 VTAIL.n624 VSUBS 0.012258f
C682 VTAIL.n625 VSUBS 0.027683f
C683 VTAIL.n626 VSUBS 0.012401f
C684 VTAIL.n627 VSUBS 0.021795f
C685 VTAIL.n628 VSUBS 0.011712f
C686 VTAIL.n629 VSUBS 0.027683f
C687 VTAIL.n630 VSUBS 0.012401f
C688 VTAIL.n631 VSUBS 0.021795f
C689 VTAIL.n632 VSUBS 0.011712f
C690 VTAIL.n633 VSUBS 0.027683f
C691 VTAIL.n634 VSUBS 0.012401f
C692 VTAIL.n635 VSUBS 0.021795f
C693 VTAIL.n636 VSUBS 0.011712f
C694 VTAIL.n637 VSUBS 0.027683f
C695 VTAIL.n638 VSUBS 0.012401f
C696 VTAIL.n639 VSUBS 0.021795f
C697 VTAIL.n640 VSUBS 0.011712f
C698 VTAIL.n641 VSUBS 0.027683f
C699 VTAIL.n642 VSUBS 0.012401f
C700 VTAIL.n643 VSUBS 0.021795f
C701 VTAIL.n644 VSUBS 0.011712f
C702 VTAIL.n645 VSUBS 0.027683f
C703 VTAIL.n646 VSUBS 0.012056f
C704 VTAIL.n647 VSUBS 0.021795f
C705 VTAIL.n648 VSUBS 0.012056f
C706 VTAIL.n649 VSUBS 0.011712f
C707 VTAIL.n650 VSUBS 0.027683f
C708 VTAIL.n651 VSUBS 0.027683f
C709 VTAIL.n652 VSUBS 0.012401f
C710 VTAIL.n653 VSUBS 0.021795f
C711 VTAIL.n654 VSUBS 0.011712f
C712 VTAIL.n655 VSUBS 0.027683f
C713 VTAIL.n656 VSUBS 0.012401f
C714 VTAIL.n657 VSUBS 1.71454f
C715 VTAIL.n658 VSUBS 0.011712f
C716 VTAIL.t1 VSUBS 0.060149f
C717 VTAIL.n659 VSUBS 0.238073f
C718 VTAIL.n660 VSUBS 0.020824f
C719 VTAIL.n661 VSUBS 0.020762f
C720 VTAIL.n662 VSUBS 0.027683f
C721 VTAIL.n663 VSUBS 0.012401f
C722 VTAIL.n664 VSUBS 0.011712f
C723 VTAIL.n665 VSUBS 0.021795f
C724 VTAIL.n666 VSUBS 0.021795f
C725 VTAIL.n667 VSUBS 0.011712f
C726 VTAIL.n668 VSUBS 0.012401f
C727 VTAIL.n669 VSUBS 0.027683f
C728 VTAIL.n670 VSUBS 0.027683f
C729 VTAIL.n671 VSUBS 0.012401f
C730 VTAIL.n672 VSUBS 0.011712f
C731 VTAIL.n673 VSUBS 0.021795f
C732 VTAIL.n674 VSUBS 0.021795f
C733 VTAIL.n675 VSUBS 0.011712f
C734 VTAIL.n676 VSUBS 0.012401f
C735 VTAIL.n677 VSUBS 0.027683f
C736 VTAIL.n678 VSUBS 0.027683f
C737 VTAIL.n679 VSUBS 0.012401f
C738 VTAIL.n680 VSUBS 0.011712f
C739 VTAIL.n681 VSUBS 0.021795f
C740 VTAIL.n682 VSUBS 0.021795f
C741 VTAIL.n683 VSUBS 0.011712f
C742 VTAIL.n684 VSUBS 0.012401f
C743 VTAIL.n685 VSUBS 0.027683f
C744 VTAIL.n686 VSUBS 0.027683f
C745 VTAIL.n687 VSUBS 0.012401f
C746 VTAIL.n688 VSUBS 0.011712f
C747 VTAIL.n689 VSUBS 0.021795f
C748 VTAIL.n690 VSUBS 0.021795f
C749 VTAIL.n691 VSUBS 0.011712f
C750 VTAIL.n692 VSUBS 0.012401f
C751 VTAIL.n693 VSUBS 0.027683f
C752 VTAIL.n694 VSUBS 0.027683f
C753 VTAIL.n695 VSUBS 0.012401f
C754 VTAIL.n696 VSUBS 0.011712f
C755 VTAIL.n697 VSUBS 0.021795f
C756 VTAIL.n698 VSUBS 0.021795f
C757 VTAIL.n699 VSUBS 0.011712f
C758 VTAIL.n700 VSUBS 0.012401f
C759 VTAIL.n701 VSUBS 0.027683f
C760 VTAIL.n702 VSUBS 0.027683f
C761 VTAIL.n703 VSUBS 0.012401f
C762 VTAIL.n704 VSUBS 0.011712f
C763 VTAIL.n705 VSUBS 0.021795f
C764 VTAIL.n706 VSUBS 0.021795f
C765 VTAIL.n707 VSUBS 0.011712f
C766 VTAIL.n708 VSUBS 0.012401f
C767 VTAIL.n709 VSUBS 0.027683f
C768 VTAIL.n710 VSUBS 0.027683f
C769 VTAIL.n711 VSUBS 0.012401f
C770 VTAIL.n712 VSUBS 0.011712f
C771 VTAIL.n713 VSUBS 0.021795f
C772 VTAIL.n714 VSUBS 0.021795f
C773 VTAIL.n715 VSUBS 0.011712f
C774 VTAIL.n716 VSUBS 0.012401f
C775 VTAIL.n717 VSUBS 0.027683f
C776 VTAIL.n718 VSUBS 0.027683f
C777 VTAIL.n719 VSUBS 0.012401f
C778 VTAIL.n720 VSUBS 0.011712f
C779 VTAIL.n721 VSUBS 0.021795f
C780 VTAIL.n722 VSUBS 0.054547f
C781 VTAIL.n723 VSUBS 0.011712f
C782 VTAIL.n724 VSUBS 0.012401f
C783 VTAIL.n725 VSUBS 0.061041f
C784 VTAIL.n726 VSUBS 0.04014f
C785 VTAIL.n727 VSUBS 1.7225f
C786 VTAIL.n728 VSUBS 0.012258f
C787 VTAIL.n729 VSUBS 0.027683f
C788 VTAIL.n730 VSUBS 0.012401f
C789 VTAIL.n731 VSUBS 0.021795f
C790 VTAIL.n732 VSUBS 0.011712f
C791 VTAIL.n733 VSUBS 0.027683f
C792 VTAIL.n734 VSUBS 0.012401f
C793 VTAIL.n735 VSUBS 0.021795f
C794 VTAIL.n736 VSUBS 0.011712f
C795 VTAIL.n737 VSUBS 0.027683f
C796 VTAIL.n738 VSUBS 0.012401f
C797 VTAIL.n739 VSUBS 0.021795f
C798 VTAIL.n740 VSUBS 0.011712f
C799 VTAIL.n741 VSUBS 0.027683f
C800 VTAIL.n742 VSUBS 0.012401f
C801 VTAIL.n743 VSUBS 0.021795f
C802 VTAIL.n744 VSUBS 0.011712f
C803 VTAIL.n745 VSUBS 0.027683f
C804 VTAIL.n746 VSUBS 0.012401f
C805 VTAIL.n747 VSUBS 0.021795f
C806 VTAIL.n748 VSUBS 0.011712f
C807 VTAIL.n749 VSUBS 0.027683f
C808 VTAIL.n750 VSUBS 0.012056f
C809 VTAIL.n751 VSUBS 0.021795f
C810 VTAIL.n752 VSUBS 0.012401f
C811 VTAIL.n753 VSUBS 0.027683f
C812 VTAIL.n754 VSUBS 0.012401f
C813 VTAIL.n755 VSUBS 0.021795f
C814 VTAIL.n756 VSUBS 0.011712f
C815 VTAIL.n757 VSUBS 0.027683f
C816 VTAIL.n758 VSUBS 0.012401f
C817 VTAIL.n759 VSUBS 1.71454f
C818 VTAIL.n760 VSUBS 0.011712f
C819 VTAIL.t6 VSUBS 0.060149f
C820 VTAIL.n761 VSUBS 0.238073f
C821 VTAIL.n762 VSUBS 0.020824f
C822 VTAIL.n763 VSUBS 0.020762f
C823 VTAIL.n764 VSUBS 0.027683f
C824 VTAIL.n765 VSUBS 0.012401f
C825 VTAIL.n766 VSUBS 0.011712f
C826 VTAIL.n767 VSUBS 0.021795f
C827 VTAIL.n768 VSUBS 0.021795f
C828 VTAIL.n769 VSUBS 0.011712f
C829 VTAIL.n770 VSUBS 0.012401f
C830 VTAIL.n771 VSUBS 0.027683f
C831 VTAIL.n772 VSUBS 0.027683f
C832 VTAIL.n773 VSUBS 0.012401f
C833 VTAIL.n774 VSUBS 0.011712f
C834 VTAIL.n775 VSUBS 0.021795f
C835 VTAIL.n776 VSUBS 0.021795f
C836 VTAIL.n777 VSUBS 0.011712f
C837 VTAIL.n778 VSUBS 0.011712f
C838 VTAIL.n779 VSUBS 0.012401f
C839 VTAIL.n780 VSUBS 0.027683f
C840 VTAIL.n781 VSUBS 0.027683f
C841 VTAIL.n782 VSUBS 0.027683f
C842 VTAIL.n783 VSUBS 0.012056f
C843 VTAIL.n784 VSUBS 0.011712f
C844 VTAIL.n785 VSUBS 0.021795f
C845 VTAIL.n786 VSUBS 0.021795f
C846 VTAIL.n787 VSUBS 0.011712f
C847 VTAIL.n788 VSUBS 0.012401f
C848 VTAIL.n789 VSUBS 0.027683f
C849 VTAIL.n790 VSUBS 0.027683f
C850 VTAIL.n791 VSUBS 0.012401f
C851 VTAIL.n792 VSUBS 0.011712f
C852 VTAIL.n793 VSUBS 0.021795f
C853 VTAIL.n794 VSUBS 0.021795f
C854 VTAIL.n795 VSUBS 0.011712f
C855 VTAIL.n796 VSUBS 0.012401f
C856 VTAIL.n797 VSUBS 0.027683f
C857 VTAIL.n798 VSUBS 0.027683f
C858 VTAIL.n799 VSUBS 0.012401f
C859 VTAIL.n800 VSUBS 0.011712f
C860 VTAIL.n801 VSUBS 0.021795f
C861 VTAIL.n802 VSUBS 0.021795f
C862 VTAIL.n803 VSUBS 0.011712f
C863 VTAIL.n804 VSUBS 0.012401f
C864 VTAIL.n805 VSUBS 0.027683f
C865 VTAIL.n806 VSUBS 0.027683f
C866 VTAIL.n807 VSUBS 0.012401f
C867 VTAIL.n808 VSUBS 0.011712f
C868 VTAIL.n809 VSUBS 0.021795f
C869 VTAIL.n810 VSUBS 0.021795f
C870 VTAIL.n811 VSUBS 0.011712f
C871 VTAIL.n812 VSUBS 0.012401f
C872 VTAIL.n813 VSUBS 0.027683f
C873 VTAIL.n814 VSUBS 0.027683f
C874 VTAIL.n815 VSUBS 0.012401f
C875 VTAIL.n816 VSUBS 0.011712f
C876 VTAIL.n817 VSUBS 0.021795f
C877 VTAIL.n818 VSUBS 0.021795f
C878 VTAIL.n819 VSUBS 0.011712f
C879 VTAIL.n820 VSUBS 0.012401f
C880 VTAIL.n821 VSUBS 0.027683f
C881 VTAIL.n822 VSUBS 0.027683f
C882 VTAIL.n823 VSUBS 0.012401f
C883 VTAIL.n824 VSUBS 0.011712f
C884 VTAIL.n825 VSUBS 0.021795f
C885 VTAIL.n826 VSUBS 0.054547f
C886 VTAIL.n827 VSUBS 0.011712f
C887 VTAIL.n828 VSUBS 0.012401f
C888 VTAIL.n829 VSUBS 0.061041f
C889 VTAIL.n830 VSUBS 0.04014f
C890 VTAIL.n831 VSUBS 1.6506f
C891 VDD2.t0 VSUBS 0.393215f
C892 VDD2.t2 VSUBS 0.393215f
C893 VDD2.n0 VSUBS 4.22394f
C894 VDD2.t3 VSUBS 0.393215f
C895 VDD2.t1 VSUBS 0.393215f
C896 VDD2.n1 VSUBS 3.30336f
C897 VDD2.n2 VSUBS 4.82891f
C898 VN.t0 VSUBS 3.64549f
C899 VN.t1 VSUBS 3.64282f
C900 VN.n0 VSUBS 2.48979f
C901 VN.t2 VSUBS 3.64549f
C902 VN.t3 VSUBS 3.64282f
C903 VN.n1 VSUBS 4.36127f
C904 B.n0 VSUBS 0.004093f
C905 B.n1 VSUBS 0.004093f
C906 B.n2 VSUBS 0.006473f
C907 B.n3 VSUBS 0.006473f
C908 B.n4 VSUBS 0.006473f
C909 B.n5 VSUBS 0.006473f
C910 B.n6 VSUBS 0.006473f
C911 B.n7 VSUBS 0.006473f
C912 B.n8 VSUBS 0.006473f
C913 B.n9 VSUBS 0.006473f
C914 B.n10 VSUBS 0.006473f
C915 B.n11 VSUBS 0.006473f
C916 B.n12 VSUBS 0.006473f
C917 B.n13 VSUBS 0.006473f
C918 B.n14 VSUBS 0.006473f
C919 B.n15 VSUBS 0.006473f
C920 B.n16 VSUBS 0.015556f
C921 B.n17 VSUBS 0.006473f
C922 B.n18 VSUBS 0.006473f
C923 B.n19 VSUBS 0.006473f
C924 B.n20 VSUBS 0.006473f
C925 B.n21 VSUBS 0.006473f
C926 B.n22 VSUBS 0.006473f
C927 B.n23 VSUBS 0.006473f
C928 B.n24 VSUBS 0.006473f
C929 B.n25 VSUBS 0.006473f
C930 B.n26 VSUBS 0.006473f
C931 B.n27 VSUBS 0.006473f
C932 B.n28 VSUBS 0.006473f
C933 B.n29 VSUBS 0.006473f
C934 B.n30 VSUBS 0.006473f
C935 B.n31 VSUBS 0.006473f
C936 B.n32 VSUBS 0.006473f
C937 B.n33 VSUBS 0.006473f
C938 B.n34 VSUBS 0.006473f
C939 B.n35 VSUBS 0.006473f
C940 B.n36 VSUBS 0.006473f
C941 B.n37 VSUBS 0.006473f
C942 B.n38 VSUBS 0.006473f
C943 B.n39 VSUBS 0.006473f
C944 B.n40 VSUBS 0.006473f
C945 B.n41 VSUBS 0.006473f
C946 B.n42 VSUBS 0.006473f
C947 B.n43 VSUBS 0.006473f
C948 B.n44 VSUBS 0.006473f
C949 B.n45 VSUBS 0.006473f
C950 B.n46 VSUBS 0.006092f
C951 B.n47 VSUBS 0.006473f
C952 B.t11 VSUBS 0.341047f
C953 B.t10 VSUBS 0.3652f
C954 B.t9 VSUBS 1.42997f
C955 B.n48 VSUBS 0.530412f
C956 B.n49 VSUBS 0.309613f
C957 B.n50 VSUBS 0.014996f
C958 B.n51 VSUBS 0.006473f
C959 B.n52 VSUBS 0.006473f
C960 B.n53 VSUBS 0.006473f
C961 B.n54 VSUBS 0.006473f
C962 B.t8 VSUBS 0.341051f
C963 B.t7 VSUBS 0.365203f
C964 B.t6 VSUBS 1.42997f
C965 B.n55 VSUBS 0.530409f
C966 B.n56 VSUBS 0.309609f
C967 B.n57 VSUBS 0.006473f
C968 B.n58 VSUBS 0.006473f
C969 B.n59 VSUBS 0.006473f
C970 B.n60 VSUBS 0.006473f
C971 B.n61 VSUBS 0.006473f
C972 B.n62 VSUBS 0.006473f
C973 B.n63 VSUBS 0.006473f
C974 B.n64 VSUBS 0.006473f
C975 B.n65 VSUBS 0.006473f
C976 B.n66 VSUBS 0.006473f
C977 B.n67 VSUBS 0.006473f
C978 B.n68 VSUBS 0.006473f
C979 B.n69 VSUBS 0.006473f
C980 B.n70 VSUBS 0.006473f
C981 B.n71 VSUBS 0.006473f
C982 B.n72 VSUBS 0.006473f
C983 B.n73 VSUBS 0.006473f
C984 B.n74 VSUBS 0.006473f
C985 B.n75 VSUBS 0.006473f
C986 B.n76 VSUBS 0.006473f
C987 B.n77 VSUBS 0.006473f
C988 B.n78 VSUBS 0.006473f
C989 B.n79 VSUBS 0.006473f
C990 B.n80 VSUBS 0.006473f
C991 B.n81 VSUBS 0.006473f
C992 B.n82 VSUBS 0.006473f
C993 B.n83 VSUBS 0.006473f
C994 B.n84 VSUBS 0.006473f
C995 B.n85 VSUBS 0.006473f
C996 B.n86 VSUBS 0.006473f
C997 B.n87 VSUBS 0.016028f
C998 B.n88 VSUBS 0.006473f
C999 B.n89 VSUBS 0.006473f
C1000 B.n90 VSUBS 0.006473f
C1001 B.n91 VSUBS 0.006473f
C1002 B.n92 VSUBS 0.006473f
C1003 B.n93 VSUBS 0.006473f
C1004 B.n94 VSUBS 0.006473f
C1005 B.n95 VSUBS 0.006473f
C1006 B.n96 VSUBS 0.006473f
C1007 B.n97 VSUBS 0.006473f
C1008 B.n98 VSUBS 0.006473f
C1009 B.n99 VSUBS 0.006473f
C1010 B.n100 VSUBS 0.006473f
C1011 B.n101 VSUBS 0.006473f
C1012 B.n102 VSUBS 0.006473f
C1013 B.n103 VSUBS 0.006473f
C1014 B.n104 VSUBS 0.006473f
C1015 B.n105 VSUBS 0.006473f
C1016 B.n106 VSUBS 0.006473f
C1017 B.n107 VSUBS 0.006473f
C1018 B.n108 VSUBS 0.006473f
C1019 B.n109 VSUBS 0.006473f
C1020 B.n110 VSUBS 0.006473f
C1021 B.n111 VSUBS 0.006473f
C1022 B.n112 VSUBS 0.006473f
C1023 B.n113 VSUBS 0.006473f
C1024 B.n114 VSUBS 0.006473f
C1025 B.n115 VSUBS 0.015284f
C1026 B.n116 VSUBS 0.006473f
C1027 B.n117 VSUBS 0.006473f
C1028 B.n118 VSUBS 0.006473f
C1029 B.n119 VSUBS 0.006473f
C1030 B.n120 VSUBS 0.006473f
C1031 B.n121 VSUBS 0.006473f
C1032 B.n122 VSUBS 0.006473f
C1033 B.n123 VSUBS 0.006473f
C1034 B.n124 VSUBS 0.006473f
C1035 B.n125 VSUBS 0.006473f
C1036 B.n126 VSUBS 0.006473f
C1037 B.n127 VSUBS 0.006473f
C1038 B.n128 VSUBS 0.006473f
C1039 B.n129 VSUBS 0.006473f
C1040 B.n130 VSUBS 0.006473f
C1041 B.n131 VSUBS 0.006473f
C1042 B.n132 VSUBS 0.006473f
C1043 B.n133 VSUBS 0.006473f
C1044 B.n134 VSUBS 0.006473f
C1045 B.n135 VSUBS 0.006473f
C1046 B.n136 VSUBS 0.006473f
C1047 B.n137 VSUBS 0.006473f
C1048 B.n138 VSUBS 0.006473f
C1049 B.n139 VSUBS 0.006473f
C1050 B.n140 VSUBS 0.006473f
C1051 B.n141 VSUBS 0.006473f
C1052 B.n142 VSUBS 0.006473f
C1053 B.n143 VSUBS 0.006473f
C1054 B.n144 VSUBS 0.006473f
C1055 B.n145 VSUBS 0.006473f
C1056 B.n146 VSUBS 0.006473f
C1057 B.t4 VSUBS 0.341051f
C1058 B.t5 VSUBS 0.365203f
C1059 B.t3 VSUBS 1.42997f
C1060 B.n147 VSUBS 0.530409f
C1061 B.n148 VSUBS 0.309609f
C1062 B.n149 VSUBS 0.006473f
C1063 B.n150 VSUBS 0.006473f
C1064 B.n151 VSUBS 0.006473f
C1065 B.n152 VSUBS 0.006473f
C1066 B.t1 VSUBS 0.341047f
C1067 B.t2 VSUBS 0.3652f
C1068 B.t0 VSUBS 1.42997f
C1069 B.n153 VSUBS 0.530412f
C1070 B.n154 VSUBS 0.309613f
C1071 B.n155 VSUBS 0.014996f
C1072 B.n156 VSUBS 0.006473f
C1073 B.n157 VSUBS 0.006473f
C1074 B.n158 VSUBS 0.006473f
C1075 B.n159 VSUBS 0.006473f
C1076 B.n160 VSUBS 0.006473f
C1077 B.n161 VSUBS 0.006473f
C1078 B.n162 VSUBS 0.006473f
C1079 B.n163 VSUBS 0.006473f
C1080 B.n164 VSUBS 0.006473f
C1081 B.n165 VSUBS 0.006473f
C1082 B.n166 VSUBS 0.006473f
C1083 B.n167 VSUBS 0.006473f
C1084 B.n168 VSUBS 0.006473f
C1085 B.n169 VSUBS 0.006473f
C1086 B.n170 VSUBS 0.006473f
C1087 B.n171 VSUBS 0.006473f
C1088 B.n172 VSUBS 0.006473f
C1089 B.n173 VSUBS 0.006473f
C1090 B.n174 VSUBS 0.006473f
C1091 B.n175 VSUBS 0.006473f
C1092 B.n176 VSUBS 0.006473f
C1093 B.n177 VSUBS 0.006473f
C1094 B.n178 VSUBS 0.006473f
C1095 B.n179 VSUBS 0.006473f
C1096 B.n180 VSUBS 0.006473f
C1097 B.n181 VSUBS 0.006473f
C1098 B.n182 VSUBS 0.006473f
C1099 B.n183 VSUBS 0.006473f
C1100 B.n184 VSUBS 0.006473f
C1101 B.n185 VSUBS 0.006473f
C1102 B.n186 VSUBS 0.015284f
C1103 B.n187 VSUBS 0.006473f
C1104 B.n188 VSUBS 0.006473f
C1105 B.n189 VSUBS 0.006473f
C1106 B.n190 VSUBS 0.006473f
C1107 B.n191 VSUBS 0.006473f
C1108 B.n192 VSUBS 0.006473f
C1109 B.n193 VSUBS 0.006473f
C1110 B.n194 VSUBS 0.006473f
C1111 B.n195 VSUBS 0.006473f
C1112 B.n196 VSUBS 0.006473f
C1113 B.n197 VSUBS 0.006473f
C1114 B.n198 VSUBS 0.006473f
C1115 B.n199 VSUBS 0.006473f
C1116 B.n200 VSUBS 0.006473f
C1117 B.n201 VSUBS 0.006473f
C1118 B.n202 VSUBS 0.006473f
C1119 B.n203 VSUBS 0.006473f
C1120 B.n204 VSUBS 0.006473f
C1121 B.n205 VSUBS 0.006473f
C1122 B.n206 VSUBS 0.006473f
C1123 B.n207 VSUBS 0.006473f
C1124 B.n208 VSUBS 0.006473f
C1125 B.n209 VSUBS 0.006473f
C1126 B.n210 VSUBS 0.006473f
C1127 B.n211 VSUBS 0.006473f
C1128 B.n212 VSUBS 0.006473f
C1129 B.n213 VSUBS 0.006473f
C1130 B.n214 VSUBS 0.006473f
C1131 B.n215 VSUBS 0.006473f
C1132 B.n216 VSUBS 0.006473f
C1133 B.n217 VSUBS 0.006473f
C1134 B.n218 VSUBS 0.006473f
C1135 B.n219 VSUBS 0.006473f
C1136 B.n220 VSUBS 0.006473f
C1137 B.n221 VSUBS 0.006473f
C1138 B.n222 VSUBS 0.006473f
C1139 B.n223 VSUBS 0.006473f
C1140 B.n224 VSUBS 0.006473f
C1141 B.n225 VSUBS 0.006473f
C1142 B.n226 VSUBS 0.006473f
C1143 B.n227 VSUBS 0.006473f
C1144 B.n228 VSUBS 0.006473f
C1145 B.n229 VSUBS 0.006473f
C1146 B.n230 VSUBS 0.006473f
C1147 B.n231 VSUBS 0.006473f
C1148 B.n232 VSUBS 0.006473f
C1149 B.n233 VSUBS 0.006473f
C1150 B.n234 VSUBS 0.006473f
C1151 B.n235 VSUBS 0.006473f
C1152 B.n236 VSUBS 0.006473f
C1153 B.n237 VSUBS 0.006473f
C1154 B.n238 VSUBS 0.006473f
C1155 B.n239 VSUBS 0.015284f
C1156 B.n240 VSUBS 0.015556f
C1157 B.n241 VSUBS 0.015556f
C1158 B.n242 VSUBS 0.006473f
C1159 B.n243 VSUBS 0.006473f
C1160 B.n244 VSUBS 0.006473f
C1161 B.n245 VSUBS 0.006473f
C1162 B.n246 VSUBS 0.006473f
C1163 B.n247 VSUBS 0.006473f
C1164 B.n248 VSUBS 0.006473f
C1165 B.n249 VSUBS 0.006473f
C1166 B.n250 VSUBS 0.006473f
C1167 B.n251 VSUBS 0.006473f
C1168 B.n252 VSUBS 0.006473f
C1169 B.n253 VSUBS 0.006473f
C1170 B.n254 VSUBS 0.006473f
C1171 B.n255 VSUBS 0.006473f
C1172 B.n256 VSUBS 0.006473f
C1173 B.n257 VSUBS 0.006473f
C1174 B.n258 VSUBS 0.006473f
C1175 B.n259 VSUBS 0.006473f
C1176 B.n260 VSUBS 0.006473f
C1177 B.n261 VSUBS 0.006473f
C1178 B.n262 VSUBS 0.006473f
C1179 B.n263 VSUBS 0.006473f
C1180 B.n264 VSUBS 0.006473f
C1181 B.n265 VSUBS 0.006473f
C1182 B.n266 VSUBS 0.006473f
C1183 B.n267 VSUBS 0.006473f
C1184 B.n268 VSUBS 0.006473f
C1185 B.n269 VSUBS 0.006473f
C1186 B.n270 VSUBS 0.006473f
C1187 B.n271 VSUBS 0.006473f
C1188 B.n272 VSUBS 0.006473f
C1189 B.n273 VSUBS 0.006473f
C1190 B.n274 VSUBS 0.006473f
C1191 B.n275 VSUBS 0.006473f
C1192 B.n276 VSUBS 0.006473f
C1193 B.n277 VSUBS 0.006473f
C1194 B.n278 VSUBS 0.006473f
C1195 B.n279 VSUBS 0.006473f
C1196 B.n280 VSUBS 0.006473f
C1197 B.n281 VSUBS 0.006473f
C1198 B.n282 VSUBS 0.006473f
C1199 B.n283 VSUBS 0.006473f
C1200 B.n284 VSUBS 0.006473f
C1201 B.n285 VSUBS 0.006473f
C1202 B.n286 VSUBS 0.006473f
C1203 B.n287 VSUBS 0.006473f
C1204 B.n288 VSUBS 0.006473f
C1205 B.n289 VSUBS 0.006473f
C1206 B.n290 VSUBS 0.006473f
C1207 B.n291 VSUBS 0.006473f
C1208 B.n292 VSUBS 0.006473f
C1209 B.n293 VSUBS 0.006473f
C1210 B.n294 VSUBS 0.006473f
C1211 B.n295 VSUBS 0.006473f
C1212 B.n296 VSUBS 0.006473f
C1213 B.n297 VSUBS 0.006473f
C1214 B.n298 VSUBS 0.006473f
C1215 B.n299 VSUBS 0.006473f
C1216 B.n300 VSUBS 0.006473f
C1217 B.n301 VSUBS 0.006473f
C1218 B.n302 VSUBS 0.006473f
C1219 B.n303 VSUBS 0.006473f
C1220 B.n304 VSUBS 0.006473f
C1221 B.n305 VSUBS 0.006473f
C1222 B.n306 VSUBS 0.006473f
C1223 B.n307 VSUBS 0.006473f
C1224 B.n308 VSUBS 0.006473f
C1225 B.n309 VSUBS 0.006473f
C1226 B.n310 VSUBS 0.006473f
C1227 B.n311 VSUBS 0.006473f
C1228 B.n312 VSUBS 0.006473f
C1229 B.n313 VSUBS 0.006473f
C1230 B.n314 VSUBS 0.006473f
C1231 B.n315 VSUBS 0.006473f
C1232 B.n316 VSUBS 0.006473f
C1233 B.n317 VSUBS 0.006473f
C1234 B.n318 VSUBS 0.006473f
C1235 B.n319 VSUBS 0.006473f
C1236 B.n320 VSUBS 0.006473f
C1237 B.n321 VSUBS 0.006473f
C1238 B.n322 VSUBS 0.006473f
C1239 B.n323 VSUBS 0.006473f
C1240 B.n324 VSUBS 0.006473f
C1241 B.n325 VSUBS 0.006473f
C1242 B.n326 VSUBS 0.006473f
C1243 B.n327 VSUBS 0.006473f
C1244 B.n328 VSUBS 0.006473f
C1245 B.n329 VSUBS 0.006473f
C1246 B.n330 VSUBS 0.006092f
C1247 B.n331 VSUBS 0.006473f
C1248 B.n332 VSUBS 0.006473f
C1249 B.n333 VSUBS 0.003617f
C1250 B.n334 VSUBS 0.006473f
C1251 B.n335 VSUBS 0.006473f
C1252 B.n336 VSUBS 0.006473f
C1253 B.n337 VSUBS 0.006473f
C1254 B.n338 VSUBS 0.006473f
C1255 B.n339 VSUBS 0.006473f
C1256 B.n340 VSUBS 0.006473f
C1257 B.n341 VSUBS 0.006473f
C1258 B.n342 VSUBS 0.006473f
C1259 B.n343 VSUBS 0.006473f
C1260 B.n344 VSUBS 0.006473f
C1261 B.n345 VSUBS 0.006473f
C1262 B.n346 VSUBS 0.003617f
C1263 B.n347 VSUBS 0.014996f
C1264 B.n348 VSUBS 0.006092f
C1265 B.n349 VSUBS 0.006473f
C1266 B.n350 VSUBS 0.006473f
C1267 B.n351 VSUBS 0.006473f
C1268 B.n352 VSUBS 0.006473f
C1269 B.n353 VSUBS 0.006473f
C1270 B.n354 VSUBS 0.006473f
C1271 B.n355 VSUBS 0.006473f
C1272 B.n356 VSUBS 0.006473f
C1273 B.n357 VSUBS 0.006473f
C1274 B.n358 VSUBS 0.006473f
C1275 B.n359 VSUBS 0.006473f
C1276 B.n360 VSUBS 0.006473f
C1277 B.n361 VSUBS 0.006473f
C1278 B.n362 VSUBS 0.006473f
C1279 B.n363 VSUBS 0.006473f
C1280 B.n364 VSUBS 0.006473f
C1281 B.n365 VSUBS 0.006473f
C1282 B.n366 VSUBS 0.006473f
C1283 B.n367 VSUBS 0.006473f
C1284 B.n368 VSUBS 0.006473f
C1285 B.n369 VSUBS 0.006473f
C1286 B.n370 VSUBS 0.006473f
C1287 B.n371 VSUBS 0.006473f
C1288 B.n372 VSUBS 0.006473f
C1289 B.n373 VSUBS 0.006473f
C1290 B.n374 VSUBS 0.006473f
C1291 B.n375 VSUBS 0.006473f
C1292 B.n376 VSUBS 0.006473f
C1293 B.n377 VSUBS 0.006473f
C1294 B.n378 VSUBS 0.006473f
C1295 B.n379 VSUBS 0.006473f
C1296 B.n380 VSUBS 0.006473f
C1297 B.n381 VSUBS 0.006473f
C1298 B.n382 VSUBS 0.006473f
C1299 B.n383 VSUBS 0.006473f
C1300 B.n384 VSUBS 0.006473f
C1301 B.n385 VSUBS 0.006473f
C1302 B.n386 VSUBS 0.006473f
C1303 B.n387 VSUBS 0.006473f
C1304 B.n388 VSUBS 0.006473f
C1305 B.n389 VSUBS 0.006473f
C1306 B.n390 VSUBS 0.006473f
C1307 B.n391 VSUBS 0.006473f
C1308 B.n392 VSUBS 0.006473f
C1309 B.n393 VSUBS 0.006473f
C1310 B.n394 VSUBS 0.006473f
C1311 B.n395 VSUBS 0.006473f
C1312 B.n396 VSUBS 0.006473f
C1313 B.n397 VSUBS 0.006473f
C1314 B.n398 VSUBS 0.006473f
C1315 B.n399 VSUBS 0.006473f
C1316 B.n400 VSUBS 0.006473f
C1317 B.n401 VSUBS 0.006473f
C1318 B.n402 VSUBS 0.006473f
C1319 B.n403 VSUBS 0.006473f
C1320 B.n404 VSUBS 0.006473f
C1321 B.n405 VSUBS 0.006473f
C1322 B.n406 VSUBS 0.006473f
C1323 B.n407 VSUBS 0.006473f
C1324 B.n408 VSUBS 0.006473f
C1325 B.n409 VSUBS 0.006473f
C1326 B.n410 VSUBS 0.006473f
C1327 B.n411 VSUBS 0.006473f
C1328 B.n412 VSUBS 0.006473f
C1329 B.n413 VSUBS 0.006473f
C1330 B.n414 VSUBS 0.006473f
C1331 B.n415 VSUBS 0.006473f
C1332 B.n416 VSUBS 0.006473f
C1333 B.n417 VSUBS 0.006473f
C1334 B.n418 VSUBS 0.006473f
C1335 B.n419 VSUBS 0.006473f
C1336 B.n420 VSUBS 0.006473f
C1337 B.n421 VSUBS 0.006473f
C1338 B.n422 VSUBS 0.006473f
C1339 B.n423 VSUBS 0.006473f
C1340 B.n424 VSUBS 0.006473f
C1341 B.n425 VSUBS 0.006473f
C1342 B.n426 VSUBS 0.006473f
C1343 B.n427 VSUBS 0.006473f
C1344 B.n428 VSUBS 0.006473f
C1345 B.n429 VSUBS 0.006473f
C1346 B.n430 VSUBS 0.006473f
C1347 B.n431 VSUBS 0.006473f
C1348 B.n432 VSUBS 0.006473f
C1349 B.n433 VSUBS 0.006473f
C1350 B.n434 VSUBS 0.006473f
C1351 B.n435 VSUBS 0.006473f
C1352 B.n436 VSUBS 0.006473f
C1353 B.n437 VSUBS 0.006473f
C1354 B.n438 VSUBS 0.015556f
C1355 B.n439 VSUBS 0.015556f
C1356 B.n440 VSUBS 0.015284f
C1357 B.n441 VSUBS 0.006473f
C1358 B.n442 VSUBS 0.006473f
C1359 B.n443 VSUBS 0.006473f
C1360 B.n444 VSUBS 0.006473f
C1361 B.n445 VSUBS 0.006473f
C1362 B.n446 VSUBS 0.006473f
C1363 B.n447 VSUBS 0.006473f
C1364 B.n448 VSUBS 0.006473f
C1365 B.n449 VSUBS 0.006473f
C1366 B.n450 VSUBS 0.006473f
C1367 B.n451 VSUBS 0.006473f
C1368 B.n452 VSUBS 0.006473f
C1369 B.n453 VSUBS 0.006473f
C1370 B.n454 VSUBS 0.006473f
C1371 B.n455 VSUBS 0.006473f
C1372 B.n456 VSUBS 0.006473f
C1373 B.n457 VSUBS 0.006473f
C1374 B.n458 VSUBS 0.006473f
C1375 B.n459 VSUBS 0.006473f
C1376 B.n460 VSUBS 0.006473f
C1377 B.n461 VSUBS 0.006473f
C1378 B.n462 VSUBS 0.006473f
C1379 B.n463 VSUBS 0.006473f
C1380 B.n464 VSUBS 0.006473f
C1381 B.n465 VSUBS 0.006473f
C1382 B.n466 VSUBS 0.006473f
C1383 B.n467 VSUBS 0.006473f
C1384 B.n468 VSUBS 0.006473f
C1385 B.n469 VSUBS 0.006473f
C1386 B.n470 VSUBS 0.006473f
C1387 B.n471 VSUBS 0.006473f
C1388 B.n472 VSUBS 0.006473f
C1389 B.n473 VSUBS 0.006473f
C1390 B.n474 VSUBS 0.006473f
C1391 B.n475 VSUBS 0.006473f
C1392 B.n476 VSUBS 0.006473f
C1393 B.n477 VSUBS 0.006473f
C1394 B.n478 VSUBS 0.006473f
C1395 B.n479 VSUBS 0.006473f
C1396 B.n480 VSUBS 0.006473f
C1397 B.n481 VSUBS 0.006473f
C1398 B.n482 VSUBS 0.006473f
C1399 B.n483 VSUBS 0.006473f
C1400 B.n484 VSUBS 0.006473f
C1401 B.n485 VSUBS 0.006473f
C1402 B.n486 VSUBS 0.006473f
C1403 B.n487 VSUBS 0.006473f
C1404 B.n488 VSUBS 0.006473f
C1405 B.n489 VSUBS 0.006473f
C1406 B.n490 VSUBS 0.006473f
C1407 B.n491 VSUBS 0.006473f
C1408 B.n492 VSUBS 0.006473f
C1409 B.n493 VSUBS 0.006473f
C1410 B.n494 VSUBS 0.006473f
C1411 B.n495 VSUBS 0.006473f
C1412 B.n496 VSUBS 0.006473f
C1413 B.n497 VSUBS 0.006473f
C1414 B.n498 VSUBS 0.006473f
C1415 B.n499 VSUBS 0.006473f
C1416 B.n500 VSUBS 0.006473f
C1417 B.n501 VSUBS 0.006473f
C1418 B.n502 VSUBS 0.006473f
C1419 B.n503 VSUBS 0.006473f
C1420 B.n504 VSUBS 0.006473f
C1421 B.n505 VSUBS 0.006473f
C1422 B.n506 VSUBS 0.006473f
C1423 B.n507 VSUBS 0.006473f
C1424 B.n508 VSUBS 0.006473f
C1425 B.n509 VSUBS 0.006473f
C1426 B.n510 VSUBS 0.006473f
C1427 B.n511 VSUBS 0.006473f
C1428 B.n512 VSUBS 0.006473f
C1429 B.n513 VSUBS 0.006473f
C1430 B.n514 VSUBS 0.006473f
C1431 B.n515 VSUBS 0.006473f
C1432 B.n516 VSUBS 0.006473f
C1433 B.n517 VSUBS 0.006473f
C1434 B.n518 VSUBS 0.006473f
C1435 B.n519 VSUBS 0.006473f
C1436 B.n520 VSUBS 0.006473f
C1437 B.n521 VSUBS 0.006473f
C1438 B.n522 VSUBS 0.006473f
C1439 B.n523 VSUBS 0.006473f
C1440 B.n524 VSUBS 0.015284f
C1441 B.n525 VSUBS 0.015556f
C1442 B.n526 VSUBS 0.014812f
C1443 B.n527 VSUBS 0.006473f
C1444 B.n528 VSUBS 0.006473f
C1445 B.n529 VSUBS 0.006473f
C1446 B.n530 VSUBS 0.006473f
C1447 B.n531 VSUBS 0.006473f
C1448 B.n532 VSUBS 0.006473f
C1449 B.n533 VSUBS 0.006473f
C1450 B.n534 VSUBS 0.006473f
C1451 B.n535 VSUBS 0.006473f
C1452 B.n536 VSUBS 0.006473f
C1453 B.n537 VSUBS 0.006473f
C1454 B.n538 VSUBS 0.006473f
C1455 B.n539 VSUBS 0.006473f
C1456 B.n540 VSUBS 0.006473f
C1457 B.n541 VSUBS 0.006473f
C1458 B.n542 VSUBS 0.006473f
C1459 B.n543 VSUBS 0.006473f
C1460 B.n544 VSUBS 0.006473f
C1461 B.n545 VSUBS 0.006473f
C1462 B.n546 VSUBS 0.006473f
C1463 B.n547 VSUBS 0.006473f
C1464 B.n548 VSUBS 0.006473f
C1465 B.n549 VSUBS 0.006473f
C1466 B.n550 VSUBS 0.006473f
C1467 B.n551 VSUBS 0.006473f
C1468 B.n552 VSUBS 0.006473f
C1469 B.n553 VSUBS 0.006473f
C1470 B.n554 VSUBS 0.006473f
C1471 B.n555 VSUBS 0.006473f
C1472 B.n556 VSUBS 0.006473f
C1473 B.n557 VSUBS 0.006473f
C1474 B.n558 VSUBS 0.006473f
C1475 B.n559 VSUBS 0.006473f
C1476 B.n560 VSUBS 0.006473f
C1477 B.n561 VSUBS 0.006473f
C1478 B.n562 VSUBS 0.006473f
C1479 B.n563 VSUBS 0.006473f
C1480 B.n564 VSUBS 0.006473f
C1481 B.n565 VSUBS 0.006473f
C1482 B.n566 VSUBS 0.006473f
C1483 B.n567 VSUBS 0.006473f
C1484 B.n568 VSUBS 0.006473f
C1485 B.n569 VSUBS 0.006473f
C1486 B.n570 VSUBS 0.006473f
C1487 B.n571 VSUBS 0.006473f
C1488 B.n572 VSUBS 0.006473f
C1489 B.n573 VSUBS 0.006473f
C1490 B.n574 VSUBS 0.006473f
C1491 B.n575 VSUBS 0.006473f
C1492 B.n576 VSUBS 0.006473f
C1493 B.n577 VSUBS 0.006473f
C1494 B.n578 VSUBS 0.006473f
C1495 B.n579 VSUBS 0.006473f
C1496 B.n580 VSUBS 0.006473f
C1497 B.n581 VSUBS 0.006473f
C1498 B.n582 VSUBS 0.006473f
C1499 B.n583 VSUBS 0.006473f
C1500 B.n584 VSUBS 0.006473f
C1501 B.n585 VSUBS 0.006473f
C1502 B.n586 VSUBS 0.006473f
C1503 B.n587 VSUBS 0.006473f
C1504 B.n588 VSUBS 0.006473f
C1505 B.n589 VSUBS 0.006473f
C1506 B.n590 VSUBS 0.006473f
C1507 B.n591 VSUBS 0.006473f
C1508 B.n592 VSUBS 0.006473f
C1509 B.n593 VSUBS 0.006473f
C1510 B.n594 VSUBS 0.006473f
C1511 B.n595 VSUBS 0.006473f
C1512 B.n596 VSUBS 0.006473f
C1513 B.n597 VSUBS 0.006473f
C1514 B.n598 VSUBS 0.006473f
C1515 B.n599 VSUBS 0.006473f
C1516 B.n600 VSUBS 0.006473f
C1517 B.n601 VSUBS 0.006473f
C1518 B.n602 VSUBS 0.006473f
C1519 B.n603 VSUBS 0.006473f
C1520 B.n604 VSUBS 0.006473f
C1521 B.n605 VSUBS 0.006473f
C1522 B.n606 VSUBS 0.006473f
C1523 B.n607 VSUBS 0.006473f
C1524 B.n608 VSUBS 0.006473f
C1525 B.n609 VSUBS 0.006473f
C1526 B.n610 VSUBS 0.006473f
C1527 B.n611 VSUBS 0.006473f
C1528 B.n612 VSUBS 0.006473f
C1529 B.n613 VSUBS 0.006473f
C1530 B.n614 VSUBS 0.006473f
C1531 B.n615 VSUBS 0.006473f
C1532 B.n616 VSUBS 0.006092f
C1533 B.n617 VSUBS 0.014996f
C1534 B.n618 VSUBS 0.003617f
C1535 B.n619 VSUBS 0.006473f
C1536 B.n620 VSUBS 0.006473f
C1537 B.n621 VSUBS 0.006473f
C1538 B.n622 VSUBS 0.006473f
C1539 B.n623 VSUBS 0.006473f
C1540 B.n624 VSUBS 0.006473f
C1541 B.n625 VSUBS 0.006473f
C1542 B.n626 VSUBS 0.006473f
C1543 B.n627 VSUBS 0.006473f
C1544 B.n628 VSUBS 0.006473f
C1545 B.n629 VSUBS 0.006473f
C1546 B.n630 VSUBS 0.006473f
C1547 B.n631 VSUBS 0.003617f
C1548 B.n632 VSUBS 0.006473f
C1549 B.n633 VSUBS 0.006473f
C1550 B.n634 VSUBS 0.006473f
C1551 B.n635 VSUBS 0.006473f
C1552 B.n636 VSUBS 0.006473f
C1553 B.n637 VSUBS 0.006473f
C1554 B.n638 VSUBS 0.006473f
C1555 B.n639 VSUBS 0.006473f
C1556 B.n640 VSUBS 0.006473f
C1557 B.n641 VSUBS 0.006473f
C1558 B.n642 VSUBS 0.006473f
C1559 B.n643 VSUBS 0.006473f
C1560 B.n644 VSUBS 0.006473f
C1561 B.n645 VSUBS 0.006473f
C1562 B.n646 VSUBS 0.006473f
C1563 B.n647 VSUBS 0.006473f
C1564 B.n648 VSUBS 0.006473f
C1565 B.n649 VSUBS 0.006473f
C1566 B.n650 VSUBS 0.006473f
C1567 B.n651 VSUBS 0.006473f
C1568 B.n652 VSUBS 0.006473f
C1569 B.n653 VSUBS 0.006473f
C1570 B.n654 VSUBS 0.006473f
C1571 B.n655 VSUBS 0.006473f
C1572 B.n656 VSUBS 0.006473f
C1573 B.n657 VSUBS 0.006473f
C1574 B.n658 VSUBS 0.006473f
C1575 B.n659 VSUBS 0.006473f
C1576 B.n660 VSUBS 0.006473f
C1577 B.n661 VSUBS 0.006473f
C1578 B.n662 VSUBS 0.006473f
C1579 B.n663 VSUBS 0.006473f
C1580 B.n664 VSUBS 0.006473f
C1581 B.n665 VSUBS 0.006473f
C1582 B.n666 VSUBS 0.006473f
C1583 B.n667 VSUBS 0.006473f
C1584 B.n668 VSUBS 0.006473f
C1585 B.n669 VSUBS 0.006473f
C1586 B.n670 VSUBS 0.006473f
C1587 B.n671 VSUBS 0.006473f
C1588 B.n672 VSUBS 0.006473f
C1589 B.n673 VSUBS 0.006473f
C1590 B.n674 VSUBS 0.006473f
C1591 B.n675 VSUBS 0.006473f
C1592 B.n676 VSUBS 0.006473f
C1593 B.n677 VSUBS 0.006473f
C1594 B.n678 VSUBS 0.006473f
C1595 B.n679 VSUBS 0.006473f
C1596 B.n680 VSUBS 0.006473f
C1597 B.n681 VSUBS 0.006473f
C1598 B.n682 VSUBS 0.006473f
C1599 B.n683 VSUBS 0.006473f
C1600 B.n684 VSUBS 0.006473f
C1601 B.n685 VSUBS 0.006473f
C1602 B.n686 VSUBS 0.006473f
C1603 B.n687 VSUBS 0.006473f
C1604 B.n688 VSUBS 0.006473f
C1605 B.n689 VSUBS 0.006473f
C1606 B.n690 VSUBS 0.006473f
C1607 B.n691 VSUBS 0.006473f
C1608 B.n692 VSUBS 0.006473f
C1609 B.n693 VSUBS 0.006473f
C1610 B.n694 VSUBS 0.006473f
C1611 B.n695 VSUBS 0.006473f
C1612 B.n696 VSUBS 0.006473f
C1613 B.n697 VSUBS 0.006473f
C1614 B.n698 VSUBS 0.006473f
C1615 B.n699 VSUBS 0.006473f
C1616 B.n700 VSUBS 0.006473f
C1617 B.n701 VSUBS 0.006473f
C1618 B.n702 VSUBS 0.006473f
C1619 B.n703 VSUBS 0.006473f
C1620 B.n704 VSUBS 0.006473f
C1621 B.n705 VSUBS 0.006473f
C1622 B.n706 VSUBS 0.006473f
C1623 B.n707 VSUBS 0.006473f
C1624 B.n708 VSUBS 0.006473f
C1625 B.n709 VSUBS 0.006473f
C1626 B.n710 VSUBS 0.006473f
C1627 B.n711 VSUBS 0.006473f
C1628 B.n712 VSUBS 0.006473f
C1629 B.n713 VSUBS 0.006473f
C1630 B.n714 VSUBS 0.006473f
C1631 B.n715 VSUBS 0.006473f
C1632 B.n716 VSUBS 0.006473f
C1633 B.n717 VSUBS 0.006473f
C1634 B.n718 VSUBS 0.006473f
C1635 B.n719 VSUBS 0.006473f
C1636 B.n720 VSUBS 0.006473f
C1637 B.n721 VSUBS 0.006473f
C1638 B.n722 VSUBS 0.006473f
C1639 B.n723 VSUBS 0.015556f
C1640 B.n724 VSUBS 0.015284f
C1641 B.n725 VSUBS 0.015284f
C1642 B.n726 VSUBS 0.006473f
C1643 B.n727 VSUBS 0.006473f
C1644 B.n728 VSUBS 0.006473f
C1645 B.n729 VSUBS 0.006473f
C1646 B.n730 VSUBS 0.006473f
C1647 B.n731 VSUBS 0.006473f
C1648 B.n732 VSUBS 0.006473f
C1649 B.n733 VSUBS 0.006473f
C1650 B.n734 VSUBS 0.006473f
C1651 B.n735 VSUBS 0.006473f
C1652 B.n736 VSUBS 0.006473f
C1653 B.n737 VSUBS 0.006473f
C1654 B.n738 VSUBS 0.006473f
C1655 B.n739 VSUBS 0.006473f
C1656 B.n740 VSUBS 0.006473f
C1657 B.n741 VSUBS 0.006473f
C1658 B.n742 VSUBS 0.006473f
C1659 B.n743 VSUBS 0.006473f
C1660 B.n744 VSUBS 0.006473f
C1661 B.n745 VSUBS 0.006473f
C1662 B.n746 VSUBS 0.006473f
C1663 B.n747 VSUBS 0.006473f
C1664 B.n748 VSUBS 0.006473f
C1665 B.n749 VSUBS 0.006473f
C1666 B.n750 VSUBS 0.006473f
C1667 B.n751 VSUBS 0.006473f
C1668 B.n752 VSUBS 0.006473f
C1669 B.n753 VSUBS 0.006473f
C1670 B.n754 VSUBS 0.006473f
C1671 B.n755 VSUBS 0.006473f
C1672 B.n756 VSUBS 0.006473f
C1673 B.n757 VSUBS 0.006473f
C1674 B.n758 VSUBS 0.006473f
C1675 B.n759 VSUBS 0.006473f
C1676 B.n760 VSUBS 0.006473f
C1677 B.n761 VSUBS 0.006473f
C1678 B.n762 VSUBS 0.006473f
C1679 B.n763 VSUBS 0.006473f
C1680 B.n764 VSUBS 0.006473f
C1681 B.n765 VSUBS 0.006473f
C1682 B.n766 VSUBS 0.006473f
C1683 B.n767 VSUBS 0.014656f
.ends

