* NGSPICE file created from diff_pair_sample_0213.ext - technology: sky130A

.subckt diff_pair_sample_0213 VTAIL VN VP B VDD2 VDD1
X0 B.t11 B.t9 B.t10 w_n1880_n1732# sky130_fd_pr__pfet_01v8 ad=1.4898 pd=8.42 as=0 ps=0 w=3.82 l=0.58
X1 VDD1.t7 VP.t0 VTAIL.t10 w_n1880_n1732# sky130_fd_pr__pfet_01v8 ad=0.6303 pd=4.15 as=0.6303 ps=4.15 w=3.82 l=0.58
X2 VTAIL.t8 VP.t1 VDD1.t6 w_n1880_n1732# sky130_fd_pr__pfet_01v8 ad=0.6303 pd=4.15 as=0.6303 ps=4.15 w=3.82 l=0.58
X3 VTAIL.t12 VP.t2 VDD1.t5 w_n1880_n1732# sky130_fd_pr__pfet_01v8 ad=1.4898 pd=8.42 as=0.6303 ps=4.15 w=3.82 l=0.58
X4 VDD2.t7 VN.t0 VTAIL.t6 w_n1880_n1732# sky130_fd_pr__pfet_01v8 ad=0.6303 pd=4.15 as=0.6303 ps=4.15 w=3.82 l=0.58
X5 B.t8 B.t6 B.t7 w_n1880_n1732# sky130_fd_pr__pfet_01v8 ad=1.4898 pd=8.42 as=0 ps=0 w=3.82 l=0.58
X6 VTAIL.t13 VP.t3 VDD1.t4 w_n1880_n1732# sky130_fd_pr__pfet_01v8 ad=0.6303 pd=4.15 as=0.6303 ps=4.15 w=3.82 l=0.58
X7 VDD2.t6 VN.t1 VTAIL.t4 w_n1880_n1732# sky130_fd_pr__pfet_01v8 ad=0.6303 pd=4.15 as=1.4898 ps=8.42 w=3.82 l=0.58
X8 VDD1.t3 VP.t4 VTAIL.t11 w_n1880_n1732# sky130_fd_pr__pfet_01v8 ad=0.6303 pd=4.15 as=1.4898 ps=8.42 w=3.82 l=0.58
X9 VDD2.t5 VN.t2 VTAIL.t5 w_n1880_n1732# sky130_fd_pr__pfet_01v8 ad=0.6303 pd=4.15 as=1.4898 ps=8.42 w=3.82 l=0.58
X10 VDD1.t2 VP.t5 VTAIL.t9 w_n1880_n1732# sky130_fd_pr__pfet_01v8 ad=0.6303 pd=4.15 as=1.4898 ps=8.42 w=3.82 l=0.58
X11 VTAIL.t3 VN.t3 VDD2.t4 w_n1880_n1732# sky130_fd_pr__pfet_01v8 ad=1.4898 pd=8.42 as=0.6303 ps=4.15 w=3.82 l=0.58
X12 B.t5 B.t3 B.t4 w_n1880_n1732# sky130_fd_pr__pfet_01v8 ad=1.4898 pd=8.42 as=0 ps=0 w=3.82 l=0.58
X13 VTAIL.t2 VN.t4 VDD2.t3 w_n1880_n1732# sky130_fd_pr__pfet_01v8 ad=0.6303 pd=4.15 as=0.6303 ps=4.15 w=3.82 l=0.58
X14 VTAIL.t1 VN.t5 VDD2.t2 w_n1880_n1732# sky130_fd_pr__pfet_01v8 ad=0.6303 pd=4.15 as=0.6303 ps=4.15 w=3.82 l=0.58
X15 VTAIL.t15 VP.t6 VDD1.t1 w_n1880_n1732# sky130_fd_pr__pfet_01v8 ad=1.4898 pd=8.42 as=0.6303 ps=4.15 w=3.82 l=0.58
X16 VDD1.t0 VP.t7 VTAIL.t14 w_n1880_n1732# sky130_fd_pr__pfet_01v8 ad=0.6303 pd=4.15 as=0.6303 ps=4.15 w=3.82 l=0.58
X17 B.t2 B.t0 B.t1 w_n1880_n1732# sky130_fd_pr__pfet_01v8 ad=1.4898 pd=8.42 as=0 ps=0 w=3.82 l=0.58
X18 VDD2.t1 VN.t6 VTAIL.t0 w_n1880_n1732# sky130_fd_pr__pfet_01v8 ad=0.6303 pd=4.15 as=0.6303 ps=4.15 w=3.82 l=0.58
X19 VTAIL.t7 VN.t7 VDD2.t0 w_n1880_n1732# sky130_fd_pr__pfet_01v8 ad=1.4898 pd=8.42 as=0.6303 ps=4.15 w=3.82 l=0.58
R0 B.n197 B.n196 585
R1 B.n195 B.n62 585
R2 B.n194 B.n193 585
R3 B.n192 B.n63 585
R4 B.n191 B.n190 585
R5 B.n189 B.n64 585
R6 B.n188 B.n187 585
R7 B.n186 B.n65 585
R8 B.n185 B.n184 585
R9 B.n183 B.n66 585
R10 B.n182 B.n181 585
R11 B.n180 B.n67 585
R12 B.n179 B.n178 585
R13 B.n177 B.n68 585
R14 B.n176 B.n175 585
R15 B.n174 B.n69 585
R16 B.n173 B.n172 585
R17 B.n171 B.n70 585
R18 B.n170 B.n169 585
R19 B.n165 B.n71 585
R20 B.n164 B.n163 585
R21 B.n162 B.n72 585
R22 B.n161 B.n160 585
R23 B.n159 B.n73 585
R24 B.n158 B.n157 585
R25 B.n156 B.n74 585
R26 B.n155 B.n154 585
R27 B.n152 B.n75 585
R28 B.n151 B.n150 585
R29 B.n149 B.n78 585
R30 B.n148 B.n147 585
R31 B.n146 B.n79 585
R32 B.n145 B.n144 585
R33 B.n143 B.n80 585
R34 B.n142 B.n141 585
R35 B.n140 B.n81 585
R36 B.n139 B.n138 585
R37 B.n137 B.n82 585
R38 B.n136 B.n135 585
R39 B.n134 B.n83 585
R40 B.n133 B.n132 585
R41 B.n131 B.n84 585
R42 B.n130 B.n129 585
R43 B.n128 B.n85 585
R44 B.n127 B.n126 585
R45 B.n198 B.n61 585
R46 B.n200 B.n199 585
R47 B.n201 B.n60 585
R48 B.n203 B.n202 585
R49 B.n204 B.n59 585
R50 B.n206 B.n205 585
R51 B.n207 B.n58 585
R52 B.n209 B.n208 585
R53 B.n210 B.n57 585
R54 B.n212 B.n211 585
R55 B.n213 B.n56 585
R56 B.n215 B.n214 585
R57 B.n216 B.n55 585
R58 B.n218 B.n217 585
R59 B.n219 B.n54 585
R60 B.n221 B.n220 585
R61 B.n222 B.n53 585
R62 B.n224 B.n223 585
R63 B.n225 B.n52 585
R64 B.n227 B.n226 585
R65 B.n228 B.n51 585
R66 B.n230 B.n229 585
R67 B.n231 B.n50 585
R68 B.n233 B.n232 585
R69 B.n234 B.n49 585
R70 B.n236 B.n235 585
R71 B.n237 B.n48 585
R72 B.n239 B.n238 585
R73 B.n240 B.n47 585
R74 B.n242 B.n241 585
R75 B.n243 B.n46 585
R76 B.n245 B.n244 585
R77 B.n246 B.n45 585
R78 B.n248 B.n247 585
R79 B.n249 B.n44 585
R80 B.n251 B.n250 585
R81 B.n252 B.n43 585
R82 B.n254 B.n253 585
R83 B.n255 B.n42 585
R84 B.n257 B.n256 585
R85 B.n258 B.n41 585
R86 B.n260 B.n259 585
R87 B.n261 B.n40 585
R88 B.n263 B.n262 585
R89 B.n332 B.n331 585
R90 B.n330 B.n13 585
R91 B.n329 B.n328 585
R92 B.n327 B.n14 585
R93 B.n326 B.n325 585
R94 B.n324 B.n15 585
R95 B.n323 B.n322 585
R96 B.n321 B.n16 585
R97 B.n320 B.n319 585
R98 B.n318 B.n17 585
R99 B.n317 B.n316 585
R100 B.n315 B.n18 585
R101 B.n314 B.n313 585
R102 B.n312 B.n19 585
R103 B.n311 B.n310 585
R104 B.n309 B.n20 585
R105 B.n308 B.n307 585
R106 B.n306 B.n21 585
R107 B.n304 B.n303 585
R108 B.n302 B.n24 585
R109 B.n301 B.n300 585
R110 B.n299 B.n25 585
R111 B.n298 B.n297 585
R112 B.n296 B.n26 585
R113 B.n295 B.n294 585
R114 B.n293 B.n27 585
R115 B.n292 B.n291 585
R116 B.n290 B.n289 585
R117 B.n288 B.n31 585
R118 B.n287 B.n286 585
R119 B.n285 B.n32 585
R120 B.n284 B.n283 585
R121 B.n282 B.n33 585
R122 B.n281 B.n280 585
R123 B.n279 B.n34 585
R124 B.n278 B.n277 585
R125 B.n276 B.n35 585
R126 B.n275 B.n274 585
R127 B.n273 B.n36 585
R128 B.n272 B.n271 585
R129 B.n270 B.n37 585
R130 B.n269 B.n268 585
R131 B.n267 B.n38 585
R132 B.n266 B.n265 585
R133 B.n264 B.n39 585
R134 B.n333 B.n12 585
R135 B.n335 B.n334 585
R136 B.n336 B.n11 585
R137 B.n338 B.n337 585
R138 B.n339 B.n10 585
R139 B.n341 B.n340 585
R140 B.n342 B.n9 585
R141 B.n344 B.n343 585
R142 B.n345 B.n8 585
R143 B.n347 B.n346 585
R144 B.n348 B.n7 585
R145 B.n350 B.n349 585
R146 B.n351 B.n6 585
R147 B.n353 B.n352 585
R148 B.n354 B.n5 585
R149 B.n356 B.n355 585
R150 B.n357 B.n4 585
R151 B.n359 B.n358 585
R152 B.n360 B.n3 585
R153 B.n362 B.n361 585
R154 B.n363 B.n0 585
R155 B.n2 B.n1 585
R156 B.n97 B.n96 585
R157 B.n98 B.n95 585
R158 B.n100 B.n99 585
R159 B.n101 B.n94 585
R160 B.n103 B.n102 585
R161 B.n104 B.n93 585
R162 B.n106 B.n105 585
R163 B.n107 B.n92 585
R164 B.n109 B.n108 585
R165 B.n110 B.n91 585
R166 B.n112 B.n111 585
R167 B.n113 B.n90 585
R168 B.n115 B.n114 585
R169 B.n116 B.n89 585
R170 B.n118 B.n117 585
R171 B.n119 B.n88 585
R172 B.n121 B.n120 585
R173 B.n122 B.n87 585
R174 B.n124 B.n123 585
R175 B.n125 B.n86 585
R176 B.n126 B.n125 473.281
R177 B.n196 B.n61 473.281
R178 B.n262 B.n39 473.281
R179 B.n333 B.n332 473.281
R180 B.n76 B.t6 363.474
R181 B.n166 B.t9 363.474
R182 B.n28 B.t3 363.474
R183 B.n22 B.t0 363.474
R184 B.n365 B.n364 256.663
R185 B.n166 B.t10 249.787
R186 B.n28 B.t5 249.787
R187 B.n76 B.t7 249.786
R188 B.n22 B.t2 249.786
R189 B.n364 B.n363 235.042
R190 B.n364 B.n2 235.042
R191 B.n167 B.t11 232.138
R192 B.n29 B.t4 232.138
R193 B.n77 B.t8 232.138
R194 B.n23 B.t1 232.138
R195 B.n126 B.n85 163.367
R196 B.n130 B.n85 163.367
R197 B.n131 B.n130 163.367
R198 B.n132 B.n131 163.367
R199 B.n132 B.n83 163.367
R200 B.n136 B.n83 163.367
R201 B.n137 B.n136 163.367
R202 B.n138 B.n137 163.367
R203 B.n138 B.n81 163.367
R204 B.n142 B.n81 163.367
R205 B.n143 B.n142 163.367
R206 B.n144 B.n143 163.367
R207 B.n144 B.n79 163.367
R208 B.n148 B.n79 163.367
R209 B.n149 B.n148 163.367
R210 B.n150 B.n149 163.367
R211 B.n150 B.n75 163.367
R212 B.n155 B.n75 163.367
R213 B.n156 B.n155 163.367
R214 B.n157 B.n156 163.367
R215 B.n157 B.n73 163.367
R216 B.n161 B.n73 163.367
R217 B.n162 B.n161 163.367
R218 B.n163 B.n162 163.367
R219 B.n163 B.n71 163.367
R220 B.n170 B.n71 163.367
R221 B.n171 B.n170 163.367
R222 B.n172 B.n171 163.367
R223 B.n172 B.n69 163.367
R224 B.n176 B.n69 163.367
R225 B.n177 B.n176 163.367
R226 B.n178 B.n177 163.367
R227 B.n178 B.n67 163.367
R228 B.n182 B.n67 163.367
R229 B.n183 B.n182 163.367
R230 B.n184 B.n183 163.367
R231 B.n184 B.n65 163.367
R232 B.n188 B.n65 163.367
R233 B.n189 B.n188 163.367
R234 B.n190 B.n189 163.367
R235 B.n190 B.n63 163.367
R236 B.n194 B.n63 163.367
R237 B.n195 B.n194 163.367
R238 B.n196 B.n195 163.367
R239 B.n262 B.n261 163.367
R240 B.n261 B.n260 163.367
R241 B.n260 B.n41 163.367
R242 B.n256 B.n41 163.367
R243 B.n256 B.n255 163.367
R244 B.n255 B.n254 163.367
R245 B.n254 B.n43 163.367
R246 B.n250 B.n43 163.367
R247 B.n250 B.n249 163.367
R248 B.n249 B.n248 163.367
R249 B.n248 B.n45 163.367
R250 B.n244 B.n45 163.367
R251 B.n244 B.n243 163.367
R252 B.n243 B.n242 163.367
R253 B.n242 B.n47 163.367
R254 B.n238 B.n47 163.367
R255 B.n238 B.n237 163.367
R256 B.n237 B.n236 163.367
R257 B.n236 B.n49 163.367
R258 B.n232 B.n49 163.367
R259 B.n232 B.n231 163.367
R260 B.n231 B.n230 163.367
R261 B.n230 B.n51 163.367
R262 B.n226 B.n51 163.367
R263 B.n226 B.n225 163.367
R264 B.n225 B.n224 163.367
R265 B.n224 B.n53 163.367
R266 B.n220 B.n53 163.367
R267 B.n220 B.n219 163.367
R268 B.n219 B.n218 163.367
R269 B.n218 B.n55 163.367
R270 B.n214 B.n55 163.367
R271 B.n214 B.n213 163.367
R272 B.n213 B.n212 163.367
R273 B.n212 B.n57 163.367
R274 B.n208 B.n57 163.367
R275 B.n208 B.n207 163.367
R276 B.n207 B.n206 163.367
R277 B.n206 B.n59 163.367
R278 B.n202 B.n59 163.367
R279 B.n202 B.n201 163.367
R280 B.n201 B.n200 163.367
R281 B.n200 B.n61 163.367
R282 B.n332 B.n13 163.367
R283 B.n328 B.n13 163.367
R284 B.n328 B.n327 163.367
R285 B.n327 B.n326 163.367
R286 B.n326 B.n15 163.367
R287 B.n322 B.n15 163.367
R288 B.n322 B.n321 163.367
R289 B.n321 B.n320 163.367
R290 B.n320 B.n17 163.367
R291 B.n316 B.n17 163.367
R292 B.n316 B.n315 163.367
R293 B.n315 B.n314 163.367
R294 B.n314 B.n19 163.367
R295 B.n310 B.n19 163.367
R296 B.n310 B.n309 163.367
R297 B.n309 B.n308 163.367
R298 B.n308 B.n21 163.367
R299 B.n303 B.n21 163.367
R300 B.n303 B.n302 163.367
R301 B.n302 B.n301 163.367
R302 B.n301 B.n25 163.367
R303 B.n297 B.n25 163.367
R304 B.n297 B.n296 163.367
R305 B.n296 B.n295 163.367
R306 B.n295 B.n27 163.367
R307 B.n291 B.n27 163.367
R308 B.n291 B.n290 163.367
R309 B.n290 B.n31 163.367
R310 B.n286 B.n31 163.367
R311 B.n286 B.n285 163.367
R312 B.n285 B.n284 163.367
R313 B.n284 B.n33 163.367
R314 B.n280 B.n33 163.367
R315 B.n280 B.n279 163.367
R316 B.n279 B.n278 163.367
R317 B.n278 B.n35 163.367
R318 B.n274 B.n35 163.367
R319 B.n274 B.n273 163.367
R320 B.n273 B.n272 163.367
R321 B.n272 B.n37 163.367
R322 B.n268 B.n37 163.367
R323 B.n268 B.n267 163.367
R324 B.n267 B.n266 163.367
R325 B.n266 B.n39 163.367
R326 B.n334 B.n333 163.367
R327 B.n334 B.n11 163.367
R328 B.n338 B.n11 163.367
R329 B.n339 B.n338 163.367
R330 B.n340 B.n339 163.367
R331 B.n340 B.n9 163.367
R332 B.n344 B.n9 163.367
R333 B.n345 B.n344 163.367
R334 B.n346 B.n345 163.367
R335 B.n346 B.n7 163.367
R336 B.n350 B.n7 163.367
R337 B.n351 B.n350 163.367
R338 B.n352 B.n351 163.367
R339 B.n352 B.n5 163.367
R340 B.n356 B.n5 163.367
R341 B.n357 B.n356 163.367
R342 B.n358 B.n357 163.367
R343 B.n358 B.n3 163.367
R344 B.n362 B.n3 163.367
R345 B.n363 B.n362 163.367
R346 B.n96 B.n2 163.367
R347 B.n96 B.n95 163.367
R348 B.n100 B.n95 163.367
R349 B.n101 B.n100 163.367
R350 B.n102 B.n101 163.367
R351 B.n102 B.n93 163.367
R352 B.n106 B.n93 163.367
R353 B.n107 B.n106 163.367
R354 B.n108 B.n107 163.367
R355 B.n108 B.n91 163.367
R356 B.n112 B.n91 163.367
R357 B.n113 B.n112 163.367
R358 B.n114 B.n113 163.367
R359 B.n114 B.n89 163.367
R360 B.n118 B.n89 163.367
R361 B.n119 B.n118 163.367
R362 B.n120 B.n119 163.367
R363 B.n120 B.n87 163.367
R364 B.n124 B.n87 163.367
R365 B.n125 B.n124 163.367
R366 B.n153 B.n77 59.5399
R367 B.n168 B.n167 59.5399
R368 B.n30 B.n29 59.5399
R369 B.n305 B.n23 59.5399
R370 B.n331 B.n12 30.7517
R371 B.n264 B.n263 30.7517
R372 B.n198 B.n197 30.7517
R373 B.n127 B.n86 30.7517
R374 B B.n365 18.0485
R375 B.n77 B.n76 17.649
R376 B.n167 B.n166 17.649
R377 B.n29 B.n28 17.649
R378 B.n23 B.n22 17.649
R379 B.n335 B.n12 10.6151
R380 B.n336 B.n335 10.6151
R381 B.n337 B.n336 10.6151
R382 B.n337 B.n10 10.6151
R383 B.n341 B.n10 10.6151
R384 B.n342 B.n341 10.6151
R385 B.n343 B.n342 10.6151
R386 B.n343 B.n8 10.6151
R387 B.n347 B.n8 10.6151
R388 B.n348 B.n347 10.6151
R389 B.n349 B.n348 10.6151
R390 B.n349 B.n6 10.6151
R391 B.n353 B.n6 10.6151
R392 B.n354 B.n353 10.6151
R393 B.n355 B.n354 10.6151
R394 B.n355 B.n4 10.6151
R395 B.n359 B.n4 10.6151
R396 B.n360 B.n359 10.6151
R397 B.n361 B.n360 10.6151
R398 B.n361 B.n0 10.6151
R399 B.n331 B.n330 10.6151
R400 B.n330 B.n329 10.6151
R401 B.n329 B.n14 10.6151
R402 B.n325 B.n14 10.6151
R403 B.n325 B.n324 10.6151
R404 B.n324 B.n323 10.6151
R405 B.n323 B.n16 10.6151
R406 B.n319 B.n16 10.6151
R407 B.n319 B.n318 10.6151
R408 B.n318 B.n317 10.6151
R409 B.n317 B.n18 10.6151
R410 B.n313 B.n18 10.6151
R411 B.n313 B.n312 10.6151
R412 B.n312 B.n311 10.6151
R413 B.n311 B.n20 10.6151
R414 B.n307 B.n20 10.6151
R415 B.n307 B.n306 10.6151
R416 B.n304 B.n24 10.6151
R417 B.n300 B.n24 10.6151
R418 B.n300 B.n299 10.6151
R419 B.n299 B.n298 10.6151
R420 B.n298 B.n26 10.6151
R421 B.n294 B.n26 10.6151
R422 B.n294 B.n293 10.6151
R423 B.n293 B.n292 10.6151
R424 B.n289 B.n288 10.6151
R425 B.n288 B.n287 10.6151
R426 B.n287 B.n32 10.6151
R427 B.n283 B.n32 10.6151
R428 B.n283 B.n282 10.6151
R429 B.n282 B.n281 10.6151
R430 B.n281 B.n34 10.6151
R431 B.n277 B.n34 10.6151
R432 B.n277 B.n276 10.6151
R433 B.n276 B.n275 10.6151
R434 B.n275 B.n36 10.6151
R435 B.n271 B.n36 10.6151
R436 B.n271 B.n270 10.6151
R437 B.n270 B.n269 10.6151
R438 B.n269 B.n38 10.6151
R439 B.n265 B.n38 10.6151
R440 B.n265 B.n264 10.6151
R441 B.n263 B.n40 10.6151
R442 B.n259 B.n40 10.6151
R443 B.n259 B.n258 10.6151
R444 B.n258 B.n257 10.6151
R445 B.n257 B.n42 10.6151
R446 B.n253 B.n42 10.6151
R447 B.n253 B.n252 10.6151
R448 B.n252 B.n251 10.6151
R449 B.n251 B.n44 10.6151
R450 B.n247 B.n44 10.6151
R451 B.n247 B.n246 10.6151
R452 B.n246 B.n245 10.6151
R453 B.n245 B.n46 10.6151
R454 B.n241 B.n46 10.6151
R455 B.n241 B.n240 10.6151
R456 B.n240 B.n239 10.6151
R457 B.n239 B.n48 10.6151
R458 B.n235 B.n48 10.6151
R459 B.n235 B.n234 10.6151
R460 B.n234 B.n233 10.6151
R461 B.n233 B.n50 10.6151
R462 B.n229 B.n50 10.6151
R463 B.n229 B.n228 10.6151
R464 B.n228 B.n227 10.6151
R465 B.n227 B.n52 10.6151
R466 B.n223 B.n52 10.6151
R467 B.n223 B.n222 10.6151
R468 B.n222 B.n221 10.6151
R469 B.n221 B.n54 10.6151
R470 B.n217 B.n54 10.6151
R471 B.n217 B.n216 10.6151
R472 B.n216 B.n215 10.6151
R473 B.n215 B.n56 10.6151
R474 B.n211 B.n56 10.6151
R475 B.n211 B.n210 10.6151
R476 B.n210 B.n209 10.6151
R477 B.n209 B.n58 10.6151
R478 B.n205 B.n58 10.6151
R479 B.n205 B.n204 10.6151
R480 B.n204 B.n203 10.6151
R481 B.n203 B.n60 10.6151
R482 B.n199 B.n60 10.6151
R483 B.n199 B.n198 10.6151
R484 B.n97 B.n1 10.6151
R485 B.n98 B.n97 10.6151
R486 B.n99 B.n98 10.6151
R487 B.n99 B.n94 10.6151
R488 B.n103 B.n94 10.6151
R489 B.n104 B.n103 10.6151
R490 B.n105 B.n104 10.6151
R491 B.n105 B.n92 10.6151
R492 B.n109 B.n92 10.6151
R493 B.n110 B.n109 10.6151
R494 B.n111 B.n110 10.6151
R495 B.n111 B.n90 10.6151
R496 B.n115 B.n90 10.6151
R497 B.n116 B.n115 10.6151
R498 B.n117 B.n116 10.6151
R499 B.n117 B.n88 10.6151
R500 B.n121 B.n88 10.6151
R501 B.n122 B.n121 10.6151
R502 B.n123 B.n122 10.6151
R503 B.n123 B.n86 10.6151
R504 B.n128 B.n127 10.6151
R505 B.n129 B.n128 10.6151
R506 B.n129 B.n84 10.6151
R507 B.n133 B.n84 10.6151
R508 B.n134 B.n133 10.6151
R509 B.n135 B.n134 10.6151
R510 B.n135 B.n82 10.6151
R511 B.n139 B.n82 10.6151
R512 B.n140 B.n139 10.6151
R513 B.n141 B.n140 10.6151
R514 B.n141 B.n80 10.6151
R515 B.n145 B.n80 10.6151
R516 B.n146 B.n145 10.6151
R517 B.n147 B.n146 10.6151
R518 B.n147 B.n78 10.6151
R519 B.n151 B.n78 10.6151
R520 B.n152 B.n151 10.6151
R521 B.n154 B.n74 10.6151
R522 B.n158 B.n74 10.6151
R523 B.n159 B.n158 10.6151
R524 B.n160 B.n159 10.6151
R525 B.n160 B.n72 10.6151
R526 B.n164 B.n72 10.6151
R527 B.n165 B.n164 10.6151
R528 B.n169 B.n165 10.6151
R529 B.n173 B.n70 10.6151
R530 B.n174 B.n173 10.6151
R531 B.n175 B.n174 10.6151
R532 B.n175 B.n68 10.6151
R533 B.n179 B.n68 10.6151
R534 B.n180 B.n179 10.6151
R535 B.n181 B.n180 10.6151
R536 B.n181 B.n66 10.6151
R537 B.n185 B.n66 10.6151
R538 B.n186 B.n185 10.6151
R539 B.n187 B.n186 10.6151
R540 B.n187 B.n64 10.6151
R541 B.n191 B.n64 10.6151
R542 B.n192 B.n191 10.6151
R543 B.n193 B.n192 10.6151
R544 B.n193 B.n62 10.6151
R545 B.n197 B.n62 10.6151
R546 B.n365 B.n0 8.11757
R547 B.n365 B.n1 8.11757
R548 B.n305 B.n304 6.5566
R549 B.n292 B.n30 6.5566
R550 B.n154 B.n153 6.5566
R551 B.n169 B.n168 6.5566
R552 B.n306 B.n305 4.05904
R553 B.n289 B.n30 4.05904
R554 B.n153 B.n152 4.05904
R555 B.n168 B.n70 4.05904
R556 VP.n4 VP.t6 253.126
R557 VP.n11 VP.t2 226.458
R558 VP.n1 VP.t7 226.458
R559 VP.n16 VP.t1 226.458
R560 VP.n18 VP.t4 226.458
R561 VP.n8 VP.t5 226.458
R562 VP.n6 VP.t3 226.458
R563 VP.n5 VP.t0 226.458
R564 VP.n19 VP.n18 161.3
R565 VP.n6 VP.n3 161.3
R566 VP.n7 VP.n2 161.3
R567 VP.n9 VP.n8 161.3
R568 VP.n17 VP.n0 161.3
R569 VP.n16 VP.n15 161.3
R570 VP.n14 VP.n1 161.3
R571 VP.n13 VP.n12 161.3
R572 VP.n11 VP.n10 161.3
R573 VP.n16 VP.n1 48.2005
R574 VP.n6 VP.n5 48.2005
R575 VP.n12 VP.n11 47.4702
R576 VP.n18 VP.n17 47.4702
R577 VP.n8 VP.n7 47.4702
R578 VP.n4 VP.n3 45.1192
R579 VP.n10 VP.n9 35.2581
R580 VP.n5 VP.n4 13.6377
R581 VP.n12 VP.n1 0.730803
R582 VP.n17 VP.n16 0.730803
R583 VP.n7 VP.n6 0.730803
R584 VP.n3 VP.n2 0.189894
R585 VP.n9 VP.n2 0.189894
R586 VP.n13 VP.n10 0.189894
R587 VP.n14 VP.n13 0.189894
R588 VP.n15 VP.n14 0.189894
R589 VP.n15 VP.n0 0.189894
R590 VP.n19 VP.n0 0.189894
R591 VP VP.n19 0.0516364
R592 VTAIL.n162 VTAIL.n148 756.745
R593 VTAIL.n16 VTAIL.n2 756.745
R594 VTAIL.n36 VTAIL.n22 756.745
R595 VTAIL.n58 VTAIL.n44 756.745
R596 VTAIL.n142 VTAIL.n128 756.745
R597 VTAIL.n120 VTAIL.n106 756.745
R598 VTAIL.n100 VTAIL.n86 756.745
R599 VTAIL.n78 VTAIL.n64 756.745
R600 VTAIL.n155 VTAIL.n154 585
R601 VTAIL.n152 VTAIL.n151 585
R602 VTAIL.n161 VTAIL.n160 585
R603 VTAIL.n163 VTAIL.n162 585
R604 VTAIL.n9 VTAIL.n8 585
R605 VTAIL.n6 VTAIL.n5 585
R606 VTAIL.n15 VTAIL.n14 585
R607 VTAIL.n17 VTAIL.n16 585
R608 VTAIL.n29 VTAIL.n28 585
R609 VTAIL.n26 VTAIL.n25 585
R610 VTAIL.n35 VTAIL.n34 585
R611 VTAIL.n37 VTAIL.n36 585
R612 VTAIL.n51 VTAIL.n50 585
R613 VTAIL.n48 VTAIL.n47 585
R614 VTAIL.n57 VTAIL.n56 585
R615 VTAIL.n59 VTAIL.n58 585
R616 VTAIL.n143 VTAIL.n142 585
R617 VTAIL.n141 VTAIL.n140 585
R618 VTAIL.n132 VTAIL.n131 585
R619 VTAIL.n135 VTAIL.n134 585
R620 VTAIL.n121 VTAIL.n120 585
R621 VTAIL.n119 VTAIL.n118 585
R622 VTAIL.n110 VTAIL.n109 585
R623 VTAIL.n113 VTAIL.n112 585
R624 VTAIL.n101 VTAIL.n100 585
R625 VTAIL.n99 VTAIL.n98 585
R626 VTAIL.n90 VTAIL.n89 585
R627 VTAIL.n93 VTAIL.n92 585
R628 VTAIL.n79 VTAIL.n78 585
R629 VTAIL.n77 VTAIL.n76 585
R630 VTAIL.n68 VTAIL.n67 585
R631 VTAIL.n71 VTAIL.n70 585
R632 VTAIL.t5 VTAIL.n153 330.707
R633 VTAIL.t3 VTAIL.n7 330.707
R634 VTAIL.t11 VTAIL.n27 330.707
R635 VTAIL.t12 VTAIL.n49 330.707
R636 VTAIL.t9 VTAIL.n133 330.707
R637 VTAIL.t15 VTAIL.n111 330.707
R638 VTAIL.t4 VTAIL.n91 330.707
R639 VTAIL.t7 VTAIL.n69 330.707
R640 VTAIL.n154 VTAIL.n151 171.744
R641 VTAIL.n161 VTAIL.n151 171.744
R642 VTAIL.n162 VTAIL.n161 171.744
R643 VTAIL.n8 VTAIL.n5 171.744
R644 VTAIL.n15 VTAIL.n5 171.744
R645 VTAIL.n16 VTAIL.n15 171.744
R646 VTAIL.n28 VTAIL.n25 171.744
R647 VTAIL.n35 VTAIL.n25 171.744
R648 VTAIL.n36 VTAIL.n35 171.744
R649 VTAIL.n50 VTAIL.n47 171.744
R650 VTAIL.n57 VTAIL.n47 171.744
R651 VTAIL.n58 VTAIL.n57 171.744
R652 VTAIL.n142 VTAIL.n141 171.744
R653 VTAIL.n141 VTAIL.n131 171.744
R654 VTAIL.n134 VTAIL.n131 171.744
R655 VTAIL.n120 VTAIL.n119 171.744
R656 VTAIL.n119 VTAIL.n109 171.744
R657 VTAIL.n112 VTAIL.n109 171.744
R658 VTAIL.n100 VTAIL.n99 171.744
R659 VTAIL.n99 VTAIL.n89 171.744
R660 VTAIL.n92 VTAIL.n89 171.744
R661 VTAIL.n78 VTAIL.n77 171.744
R662 VTAIL.n77 VTAIL.n67 171.744
R663 VTAIL.n70 VTAIL.n67 171.744
R664 VTAIL.n127 VTAIL.n126 96.5017
R665 VTAIL.n85 VTAIL.n84 96.5017
R666 VTAIL.n1 VTAIL.n0 96.5015
R667 VTAIL.n43 VTAIL.n42 96.5015
R668 VTAIL.n154 VTAIL.t5 85.8723
R669 VTAIL.n8 VTAIL.t3 85.8723
R670 VTAIL.n28 VTAIL.t11 85.8723
R671 VTAIL.n50 VTAIL.t12 85.8723
R672 VTAIL.n134 VTAIL.t9 85.8723
R673 VTAIL.n112 VTAIL.t15 85.8723
R674 VTAIL.n92 VTAIL.t4 85.8723
R675 VTAIL.n70 VTAIL.t7 85.8723
R676 VTAIL.n167 VTAIL.n166 31.7975
R677 VTAIL.n21 VTAIL.n20 31.7975
R678 VTAIL.n41 VTAIL.n40 31.7975
R679 VTAIL.n63 VTAIL.n62 31.7975
R680 VTAIL.n147 VTAIL.n146 31.7975
R681 VTAIL.n125 VTAIL.n124 31.7975
R682 VTAIL.n105 VTAIL.n104 31.7975
R683 VTAIL.n83 VTAIL.n82 31.7975
R684 VTAIL.n167 VTAIL.n147 16.4445
R685 VTAIL.n83 VTAIL.n63 16.4445
R686 VTAIL.n155 VTAIL.n153 16.3201
R687 VTAIL.n9 VTAIL.n7 16.3201
R688 VTAIL.n29 VTAIL.n27 16.3201
R689 VTAIL.n51 VTAIL.n49 16.3201
R690 VTAIL.n135 VTAIL.n133 16.3201
R691 VTAIL.n113 VTAIL.n111 16.3201
R692 VTAIL.n93 VTAIL.n91 16.3201
R693 VTAIL.n71 VTAIL.n69 16.3201
R694 VTAIL.n156 VTAIL.n152 12.8005
R695 VTAIL.n10 VTAIL.n6 12.8005
R696 VTAIL.n30 VTAIL.n26 12.8005
R697 VTAIL.n52 VTAIL.n48 12.8005
R698 VTAIL.n136 VTAIL.n132 12.8005
R699 VTAIL.n114 VTAIL.n110 12.8005
R700 VTAIL.n94 VTAIL.n90 12.8005
R701 VTAIL.n72 VTAIL.n68 12.8005
R702 VTAIL.n160 VTAIL.n159 12.0247
R703 VTAIL.n14 VTAIL.n13 12.0247
R704 VTAIL.n34 VTAIL.n33 12.0247
R705 VTAIL.n56 VTAIL.n55 12.0247
R706 VTAIL.n140 VTAIL.n139 12.0247
R707 VTAIL.n118 VTAIL.n117 12.0247
R708 VTAIL.n98 VTAIL.n97 12.0247
R709 VTAIL.n76 VTAIL.n75 12.0247
R710 VTAIL.n163 VTAIL.n150 11.249
R711 VTAIL.n17 VTAIL.n4 11.249
R712 VTAIL.n37 VTAIL.n24 11.249
R713 VTAIL.n59 VTAIL.n46 11.249
R714 VTAIL.n143 VTAIL.n130 11.249
R715 VTAIL.n121 VTAIL.n108 11.249
R716 VTAIL.n101 VTAIL.n88 11.249
R717 VTAIL.n79 VTAIL.n66 11.249
R718 VTAIL.n164 VTAIL.n148 10.4732
R719 VTAIL.n18 VTAIL.n2 10.4732
R720 VTAIL.n38 VTAIL.n22 10.4732
R721 VTAIL.n60 VTAIL.n44 10.4732
R722 VTAIL.n144 VTAIL.n128 10.4732
R723 VTAIL.n122 VTAIL.n106 10.4732
R724 VTAIL.n102 VTAIL.n86 10.4732
R725 VTAIL.n80 VTAIL.n64 10.4732
R726 VTAIL.n166 VTAIL.n165 9.45567
R727 VTAIL.n20 VTAIL.n19 9.45567
R728 VTAIL.n40 VTAIL.n39 9.45567
R729 VTAIL.n62 VTAIL.n61 9.45567
R730 VTAIL.n146 VTAIL.n145 9.45567
R731 VTAIL.n124 VTAIL.n123 9.45567
R732 VTAIL.n104 VTAIL.n103 9.45567
R733 VTAIL.n82 VTAIL.n81 9.45567
R734 VTAIL.n165 VTAIL.n164 9.3005
R735 VTAIL.n150 VTAIL.n149 9.3005
R736 VTAIL.n159 VTAIL.n158 9.3005
R737 VTAIL.n157 VTAIL.n156 9.3005
R738 VTAIL.n19 VTAIL.n18 9.3005
R739 VTAIL.n4 VTAIL.n3 9.3005
R740 VTAIL.n13 VTAIL.n12 9.3005
R741 VTAIL.n11 VTAIL.n10 9.3005
R742 VTAIL.n39 VTAIL.n38 9.3005
R743 VTAIL.n24 VTAIL.n23 9.3005
R744 VTAIL.n33 VTAIL.n32 9.3005
R745 VTAIL.n31 VTAIL.n30 9.3005
R746 VTAIL.n61 VTAIL.n60 9.3005
R747 VTAIL.n46 VTAIL.n45 9.3005
R748 VTAIL.n55 VTAIL.n54 9.3005
R749 VTAIL.n53 VTAIL.n52 9.3005
R750 VTAIL.n145 VTAIL.n144 9.3005
R751 VTAIL.n130 VTAIL.n129 9.3005
R752 VTAIL.n139 VTAIL.n138 9.3005
R753 VTAIL.n137 VTAIL.n136 9.3005
R754 VTAIL.n123 VTAIL.n122 9.3005
R755 VTAIL.n108 VTAIL.n107 9.3005
R756 VTAIL.n117 VTAIL.n116 9.3005
R757 VTAIL.n115 VTAIL.n114 9.3005
R758 VTAIL.n103 VTAIL.n102 9.3005
R759 VTAIL.n88 VTAIL.n87 9.3005
R760 VTAIL.n97 VTAIL.n96 9.3005
R761 VTAIL.n95 VTAIL.n94 9.3005
R762 VTAIL.n81 VTAIL.n80 9.3005
R763 VTAIL.n66 VTAIL.n65 9.3005
R764 VTAIL.n75 VTAIL.n74 9.3005
R765 VTAIL.n73 VTAIL.n72 9.3005
R766 VTAIL.n0 VTAIL.t6 8.50966
R767 VTAIL.n0 VTAIL.t1 8.50966
R768 VTAIL.n42 VTAIL.t14 8.50966
R769 VTAIL.n42 VTAIL.t8 8.50966
R770 VTAIL.n126 VTAIL.t10 8.50966
R771 VTAIL.n126 VTAIL.t13 8.50966
R772 VTAIL.n84 VTAIL.t0 8.50966
R773 VTAIL.n84 VTAIL.t2 8.50966
R774 VTAIL.n157 VTAIL.n153 3.78097
R775 VTAIL.n11 VTAIL.n7 3.78097
R776 VTAIL.n31 VTAIL.n27 3.78097
R777 VTAIL.n53 VTAIL.n49 3.78097
R778 VTAIL.n137 VTAIL.n133 3.78097
R779 VTAIL.n115 VTAIL.n111 3.78097
R780 VTAIL.n95 VTAIL.n91 3.78097
R781 VTAIL.n73 VTAIL.n69 3.78097
R782 VTAIL.n166 VTAIL.n148 3.49141
R783 VTAIL.n20 VTAIL.n2 3.49141
R784 VTAIL.n40 VTAIL.n22 3.49141
R785 VTAIL.n62 VTAIL.n44 3.49141
R786 VTAIL.n146 VTAIL.n128 3.49141
R787 VTAIL.n124 VTAIL.n106 3.49141
R788 VTAIL.n104 VTAIL.n86 3.49141
R789 VTAIL.n82 VTAIL.n64 3.49141
R790 VTAIL.n164 VTAIL.n163 2.71565
R791 VTAIL.n18 VTAIL.n17 2.71565
R792 VTAIL.n38 VTAIL.n37 2.71565
R793 VTAIL.n60 VTAIL.n59 2.71565
R794 VTAIL.n144 VTAIL.n143 2.71565
R795 VTAIL.n122 VTAIL.n121 2.71565
R796 VTAIL.n102 VTAIL.n101 2.71565
R797 VTAIL.n80 VTAIL.n79 2.71565
R798 VTAIL.n160 VTAIL.n150 1.93989
R799 VTAIL.n14 VTAIL.n4 1.93989
R800 VTAIL.n34 VTAIL.n24 1.93989
R801 VTAIL.n56 VTAIL.n46 1.93989
R802 VTAIL.n140 VTAIL.n130 1.93989
R803 VTAIL.n118 VTAIL.n108 1.93989
R804 VTAIL.n98 VTAIL.n88 1.93989
R805 VTAIL.n76 VTAIL.n66 1.93989
R806 VTAIL.n159 VTAIL.n152 1.16414
R807 VTAIL.n13 VTAIL.n6 1.16414
R808 VTAIL.n33 VTAIL.n26 1.16414
R809 VTAIL.n55 VTAIL.n48 1.16414
R810 VTAIL.n139 VTAIL.n132 1.16414
R811 VTAIL.n117 VTAIL.n110 1.16414
R812 VTAIL.n97 VTAIL.n90 1.16414
R813 VTAIL.n75 VTAIL.n68 1.16414
R814 VTAIL.n85 VTAIL.n83 0.784983
R815 VTAIL.n105 VTAIL.n85 0.784983
R816 VTAIL.n127 VTAIL.n125 0.784983
R817 VTAIL.n147 VTAIL.n127 0.784983
R818 VTAIL.n63 VTAIL.n43 0.784983
R819 VTAIL.n43 VTAIL.n41 0.784983
R820 VTAIL.n21 VTAIL.n1 0.784983
R821 VTAIL VTAIL.n167 0.726793
R822 VTAIL.n125 VTAIL.n105 0.470328
R823 VTAIL.n41 VTAIL.n21 0.470328
R824 VTAIL.n156 VTAIL.n155 0.388379
R825 VTAIL.n10 VTAIL.n9 0.388379
R826 VTAIL.n30 VTAIL.n29 0.388379
R827 VTAIL.n52 VTAIL.n51 0.388379
R828 VTAIL.n136 VTAIL.n135 0.388379
R829 VTAIL.n114 VTAIL.n113 0.388379
R830 VTAIL.n94 VTAIL.n93 0.388379
R831 VTAIL.n72 VTAIL.n71 0.388379
R832 VTAIL.n158 VTAIL.n157 0.155672
R833 VTAIL.n158 VTAIL.n149 0.155672
R834 VTAIL.n165 VTAIL.n149 0.155672
R835 VTAIL.n12 VTAIL.n11 0.155672
R836 VTAIL.n12 VTAIL.n3 0.155672
R837 VTAIL.n19 VTAIL.n3 0.155672
R838 VTAIL.n32 VTAIL.n31 0.155672
R839 VTAIL.n32 VTAIL.n23 0.155672
R840 VTAIL.n39 VTAIL.n23 0.155672
R841 VTAIL.n54 VTAIL.n53 0.155672
R842 VTAIL.n54 VTAIL.n45 0.155672
R843 VTAIL.n61 VTAIL.n45 0.155672
R844 VTAIL.n145 VTAIL.n129 0.155672
R845 VTAIL.n138 VTAIL.n129 0.155672
R846 VTAIL.n138 VTAIL.n137 0.155672
R847 VTAIL.n123 VTAIL.n107 0.155672
R848 VTAIL.n116 VTAIL.n107 0.155672
R849 VTAIL.n116 VTAIL.n115 0.155672
R850 VTAIL.n103 VTAIL.n87 0.155672
R851 VTAIL.n96 VTAIL.n87 0.155672
R852 VTAIL.n96 VTAIL.n95 0.155672
R853 VTAIL.n81 VTAIL.n65 0.155672
R854 VTAIL.n74 VTAIL.n65 0.155672
R855 VTAIL.n74 VTAIL.n73 0.155672
R856 VTAIL VTAIL.n1 0.0586897
R857 VDD1 VDD1.n0 113.63
R858 VDD1.n3 VDD1.n2 113.517
R859 VDD1.n3 VDD1.n1 113.517
R860 VDD1.n5 VDD1.n4 113.18
R861 VDD1.n5 VDD1.n3 31.1216
R862 VDD1.n4 VDD1.t4 8.50966
R863 VDD1.n4 VDD1.t2 8.50966
R864 VDD1.n0 VDD1.t1 8.50966
R865 VDD1.n0 VDD1.t7 8.50966
R866 VDD1.n2 VDD1.t6 8.50966
R867 VDD1.n2 VDD1.t3 8.50966
R868 VDD1.n1 VDD1.t5 8.50966
R869 VDD1.n1 VDD1.t0 8.50966
R870 VDD1 VDD1.n5 0.334552
R871 VN.n2 VN.t3 253.126
R872 VN.n10 VN.t1 253.126
R873 VN.n1 VN.t0 226.458
R874 VN.n4 VN.t5 226.458
R875 VN.n6 VN.t2 226.458
R876 VN.n9 VN.t4 226.458
R877 VN.n12 VN.t6 226.458
R878 VN.n14 VN.t7 226.458
R879 VN.n7 VN.n6 161.3
R880 VN.n15 VN.n14 161.3
R881 VN.n13 VN.n8 161.3
R882 VN.n12 VN.n11 161.3
R883 VN.n5 VN.n0 161.3
R884 VN.n4 VN.n3 161.3
R885 VN.n4 VN.n1 48.2005
R886 VN.n12 VN.n9 48.2005
R887 VN.n6 VN.n5 47.4702
R888 VN.n14 VN.n13 47.4702
R889 VN.n11 VN.n10 45.1192
R890 VN.n3 VN.n2 45.1192
R891 VN VN.n15 35.6388
R892 VN.n2 VN.n1 13.6377
R893 VN.n10 VN.n9 13.6377
R894 VN.n5 VN.n4 0.730803
R895 VN.n13 VN.n12 0.730803
R896 VN.n15 VN.n8 0.189894
R897 VN.n11 VN.n8 0.189894
R898 VN.n3 VN.n0 0.189894
R899 VN.n7 VN.n0 0.189894
R900 VN VN.n7 0.0516364
R901 VDD2.n2 VDD2.n1 113.517
R902 VDD2.n2 VDD2.n0 113.517
R903 VDD2 VDD2.n5 113.514
R904 VDD2.n4 VDD2.n3 113.18
R905 VDD2.n4 VDD2.n2 30.5386
R906 VDD2.n5 VDD2.t3 8.50966
R907 VDD2.n5 VDD2.t6 8.50966
R908 VDD2.n3 VDD2.t0 8.50966
R909 VDD2.n3 VDD2.t1 8.50966
R910 VDD2.n1 VDD2.t2 8.50966
R911 VDD2.n1 VDD2.t5 8.50966
R912 VDD2.n0 VDD2.t4 8.50966
R913 VDD2.n0 VDD2.t7 8.50966
R914 VDD2 VDD2.n4 0.450931
C0 B VTAIL 1.56537f
C1 VN VDD1 0.152829f
C2 VDD2 VP 0.309871f
C3 B VP 1.04989f
C4 VTAIL VDD1 5.21049f
C5 VTAIL VN 1.94538f
C6 VDD2 w_n1880_n1732# 1.06185f
C7 VDD1 VP 1.99508f
C8 B w_n1880_n1732# 4.72758f
C9 VN VP 3.68092f
C10 w_n1880_n1732# VDD1 1.03236f
C11 VTAIL VP 1.95948f
C12 w_n1880_n1732# VN 3.09384f
C13 VDD2 B 0.845432f
C14 w_n1880_n1732# VTAIL 2.12859f
C15 VDD2 VDD1 0.767187f
C16 VDD2 VN 1.83883f
C17 B VDD1 0.812415f
C18 w_n1880_n1732# VP 3.33082f
C19 B VN 0.661746f
C20 VDD2 VTAIL 5.25136f
C21 VDD2 VSUBS 0.833517f
C22 VDD1 VSUBS 1.101911f
C23 VTAIL VSUBS 0.388234f
C24 VN VSUBS 3.21262f
C25 VP VSUBS 1.109954f
C26 B VSUBS 1.958536f
C27 w_n1880_n1732# VSUBS 41.036602f
C28 VDD2.t4 VSUBS 0.06159f
C29 VDD2.t7 VSUBS 0.06159f
C30 VDD2.n0 VSUBS 0.355494f
C31 VDD2.t2 VSUBS 0.06159f
C32 VDD2.t5 VSUBS 0.06159f
C33 VDD2.n1 VSUBS 0.355494f
C34 VDD2.n2 VSUBS 1.55224f
C35 VDD2.t0 VSUBS 0.06159f
C36 VDD2.t1 VSUBS 0.06159f
C37 VDD2.n3 VSUBS 0.354406f
C38 VDD2.n4 VSUBS 1.41836f
C39 VDD2.t3 VSUBS 0.06159f
C40 VDD2.t6 VSUBS 0.06159f
C41 VDD2.n5 VSUBS 0.35548f
C42 VN.n0 VSUBS 0.04391f
C43 VN.t0 VSUBS 0.287634f
C44 VN.n1 VSUBS 0.165087f
C45 VN.t3 VSUBS 0.304005f
C46 VN.n2 VSUBS 0.140067f
C47 VN.n3 VSUBS 0.183128f
C48 VN.t5 VSUBS 0.287634f
C49 VN.n4 VSUBS 0.155463f
C50 VN.n5 VSUBS 0.009964f
C51 VN.t2 VSUBS 0.287634f
C52 VN.n6 VSUBS 0.155192f
C53 VN.n7 VSUBS 0.034029f
C54 VN.n8 VSUBS 0.04391f
C55 VN.t4 VSUBS 0.287634f
C56 VN.n9 VSUBS 0.165087f
C57 VN.t6 VSUBS 0.287634f
C58 VN.t1 VSUBS 0.304005f
C59 VN.n10 VSUBS 0.140067f
C60 VN.n11 VSUBS 0.183128f
C61 VN.n12 VSUBS 0.155463f
C62 VN.n13 VSUBS 0.009964f
C63 VN.t7 VSUBS 0.287634f
C64 VN.n14 VSUBS 0.155192f
C65 VN.n15 VSUBS 1.35614f
C66 VDD1.t1 VSUBS 0.059581f
C67 VDD1.t7 VSUBS 0.059581f
C68 VDD1.n0 VSUBS 0.344275f
C69 VDD1.t5 VSUBS 0.059581f
C70 VDD1.t0 VSUBS 0.059581f
C71 VDD1.n1 VSUBS 0.343896f
C72 VDD1.t6 VSUBS 0.059581f
C73 VDD1.t3 VSUBS 0.059581f
C74 VDD1.n2 VSUBS 0.343896f
C75 VDD1.n3 VSUBS 1.544f
C76 VDD1.t4 VSUBS 0.059581f
C77 VDD1.t2 VSUBS 0.059581f
C78 VDD1.n4 VSUBS 0.342843f
C79 VDD1.n5 VSUBS 1.3952f
C80 VTAIL.t6 VSUBS 0.06315f
C81 VTAIL.t1 VSUBS 0.06315f
C82 VTAIL.n0 VSUBS 0.31382f
C83 VTAIL.n1 VSUBS 0.368659f
C84 VTAIL.n2 VSUBS 0.021657f
C85 VTAIL.n3 VSUBS 0.02092f
C86 VTAIL.n4 VSUBS 0.011241f
C87 VTAIL.n5 VSUBS 0.02657f
C88 VTAIL.n6 VSUBS 0.011903f
C89 VTAIL.n7 VSUBS 0.079616f
C90 VTAIL.t3 VSUBS 0.058072f
C91 VTAIL.n8 VSUBS 0.019928f
C92 VTAIL.n9 VSUBS 0.016712f
C93 VTAIL.n10 VSUBS 0.011241f
C94 VTAIL.n11 VSUBS 0.271287f
C95 VTAIL.n12 VSUBS 0.02092f
C96 VTAIL.n13 VSUBS 0.011241f
C97 VTAIL.n14 VSUBS 0.011903f
C98 VTAIL.n15 VSUBS 0.02657f
C99 VTAIL.n16 VSUBS 0.059797f
C100 VTAIL.n17 VSUBS 0.011903f
C101 VTAIL.n18 VSUBS 0.011241f
C102 VTAIL.n19 VSUBS 0.047783f
C103 VTAIL.n20 VSUBS 0.029853f
C104 VTAIL.n21 VSUBS 0.102095f
C105 VTAIL.n22 VSUBS 0.021657f
C106 VTAIL.n23 VSUBS 0.02092f
C107 VTAIL.n24 VSUBS 0.011241f
C108 VTAIL.n25 VSUBS 0.02657f
C109 VTAIL.n26 VSUBS 0.011903f
C110 VTAIL.n27 VSUBS 0.079616f
C111 VTAIL.t11 VSUBS 0.058072f
C112 VTAIL.n28 VSUBS 0.019928f
C113 VTAIL.n29 VSUBS 0.016712f
C114 VTAIL.n30 VSUBS 0.011241f
C115 VTAIL.n31 VSUBS 0.271287f
C116 VTAIL.n32 VSUBS 0.02092f
C117 VTAIL.n33 VSUBS 0.011241f
C118 VTAIL.n34 VSUBS 0.011903f
C119 VTAIL.n35 VSUBS 0.02657f
C120 VTAIL.n36 VSUBS 0.059797f
C121 VTAIL.n37 VSUBS 0.011903f
C122 VTAIL.n38 VSUBS 0.011241f
C123 VTAIL.n39 VSUBS 0.047783f
C124 VTAIL.n40 VSUBS 0.029853f
C125 VTAIL.n41 VSUBS 0.102095f
C126 VTAIL.t14 VSUBS 0.06315f
C127 VTAIL.t8 VSUBS 0.06315f
C128 VTAIL.n42 VSUBS 0.31382f
C129 VTAIL.n43 VSUBS 0.417616f
C130 VTAIL.n44 VSUBS 0.021657f
C131 VTAIL.n45 VSUBS 0.02092f
C132 VTAIL.n46 VSUBS 0.011241f
C133 VTAIL.n47 VSUBS 0.02657f
C134 VTAIL.n48 VSUBS 0.011903f
C135 VTAIL.n49 VSUBS 0.079616f
C136 VTAIL.t12 VSUBS 0.058072f
C137 VTAIL.n50 VSUBS 0.019928f
C138 VTAIL.n51 VSUBS 0.016712f
C139 VTAIL.n52 VSUBS 0.011241f
C140 VTAIL.n53 VSUBS 0.271287f
C141 VTAIL.n54 VSUBS 0.02092f
C142 VTAIL.n55 VSUBS 0.011241f
C143 VTAIL.n56 VSUBS 0.011903f
C144 VTAIL.n57 VSUBS 0.02657f
C145 VTAIL.n58 VSUBS 0.059797f
C146 VTAIL.n59 VSUBS 0.011903f
C147 VTAIL.n60 VSUBS 0.011241f
C148 VTAIL.n61 VSUBS 0.047783f
C149 VTAIL.n62 VSUBS 0.029853f
C150 VTAIL.n63 VSUBS 0.629454f
C151 VTAIL.n64 VSUBS 0.021657f
C152 VTAIL.n65 VSUBS 0.02092f
C153 VTAIL.n66 VSUBS 0.011241f
C154 VTAIL.n67 VSUBS 0.02657f
C155 VTAIL.n68 VSUBS 0.011903f
C156 VTAIL.n69 VSUBS 0.079616f
C157 VTAIL.t7 VSUBS 0.058072f
C158 VTAIL.n70 VSUBS 0.019928f
C159 VTAIL.n71 VSUBS 0.016712f
C160 VTAIL.n72 VSUBS 0.011241f
C161 VTAIL.n73 VSUBS 0.271287f
C162 VTAIL.n74 VSUBS 0.02092f
C163 VTAIL.n75 VSUBS 0.011241f
C164 VTAIL.n76 VSUBS 0.011903f
C165 VTAIL.n77 VSUBS 0.02657f
C166 VTAIL.n78 VSUBS 0.059797f
C167 VTAIL.n79 VSUBS 0.011903f
C168 VTAIL.n80 VSUBS 0.011241f
C169 VTAIL.n81 VSUBS 0.047783f
C170 VTAIL.n82 VSUBS 0.029853f
C171 VTAIL.n83 VSUBS 0.629454f
C172 VTAIL.t0 VSUBS 0.06315f
C173 VTAIL.t2 VSUBS 0.06315f
C174 VTAIL.n84 VSUBS 0.313822f
C175 VTAIL.n85 VSUBS 0.417614f
C176 VTAIL.n86 VSUBS 0.021657f
C177 VTAIL.n87 VSUBS 0.02092f
C178 VTAIL.n88 VSUBS 0.011241f
C179 VTAIL.n89 VSUBS 0.02657f
C180 VTAIL.n90 VSUBS 0.011903f
C181 VTAIL.n91 VSUBS 0.079616f
C182 VTAIL.t4 VSUBS 0.058072f
C183 VTAIL.n92 VSUBS 0.019928f
C184 VTAIL.n93 VSUBS 0.016712f
C185 VTAIL.n94 VSUBS 0.011241f
C186 VTAIL.n95 VSUBS 0.271287f
C187 VTAIL.n96 VSUBS 0.02092f
C188 VTAIL.n97 VSUBS 0.011241f
C189 VTAIL.n98 VSUBS 0.011903f
C190 VTAIL.n99 VSUBS 0.02657f
C191 VTAIL.n100 VSUBS 0.059797f
C192 VTAIL.n101 VSUBS 0.011903f
C193 VTAIL.n102 VSUBS 0.011241f
C194 VTAIL.n103 VSUBS 0.047783f
C195 VTAIL.n104 VSUBS 0.029853f
C196 VTAIL.n105 VSUBS 0.102095f
C197 VTAIL.n106 VSUBS 0.021657f
C198 VTAIL.n107 VSUBS 0.02092f
C199 VTAIL.n108 VSUBS 0.011241f
C200 VTAIL.n109 VSUBS 0.02657f
C201 VTAIL.n110 VSUBS 0.011903f
C202 VTAIL.n111 VSUBS 0.079616f
C203 VTAIL.t15 VSUBS 0.058072f
C204 VTAIL.n112 VSUBS 0.019928f
C205 VTAIL.n113 VSUBS 0.016712f
C206 VTAIL.n114 VSUBS 0.011241f
C207 VTAIL.n115 VSUBS 0.271287f
C208 VTAIL.n116 VSUBS 0.02092f
C209 VTAIL.n117 VSUBS 0.011241f
C210 VTAIL.n118 VSUBS 0.011903f
C211 VTAIL.n119 VSUBS 0.02657f
C212 VTAIL.n120 VSUBS 0.059797f
C213 VTAIL.n121 VSUBS 0.011903f
C214 VTAIL.n122 VSUBS 0.011241f
C215 VTAIL.n123 VSUBS 0.047783f
C216 VTAIL.n124 VSUBS 0.029853f
C217 VTAIL.n125 VSUBS 0.102095f
C218 VTAIL.t10 VSUBS 0.06315f
C219 VTAIL.t13 VSUBS 0.06315f
C220 VTAIL.n126 VSUBS 0.313822f
C221 VTAIL.n127 VSUBS 0.417614f
C222 VTAIL.n128 VSUBS 0.021657f
C223 VTAIL.n129 VSUBS 0.02092f
C224 VTAIL.n130 VSUBS 0.011241f
C225 VTAIL.n131 VSUBS 0.02657f
C226 VTAIL.n132 VSUBS 0.011903f
C227 VTAIL.n133 VSUBS 0.079616f
C228 VTAIL.t9 VSUBS 0.058072f
C229 VTAIL.n134 VSUBS 0.019928f
C230 VTAIL.n135 VSUBS 0.016712f
C231 VTAIL.n136 VSUBS 0.011241f
C232 VTAIL.n137 VSUBS 0.271287f
C233 VTAIL.n138 VSUBS 0.02092f
C234 VTAIL.n139 VSUBS 0.011241f
C235 VTAIL.n140 VSUBS 0.011903f
C236 VTAIL.n141 VSUBS 0.02657f
C237 VTAIL.n142 VSUBS 0.059797f
C238 VTAIL.n143 VSUBS 0.011903f
C239 VTAIL.n144 VSUBS 0.011241f
C240 VTAIL.n145 VSUBS 0.047783f
C241 VTAIL.n146 VSUBS 0.029853f
C242 VTAIL.n147 VSUBS 0.629454f
C243 VTAIL.n148 VSUBS 0.021657f
C244 VTAIL.n149 VSUBS 0.02092f
C245 VTAIL.n150 VSUBS 0.011241f
C246 VTAIL.n151 VSUBS 0.02657f
C247 VTAIL.n152 VSUBS 0.011903f
C248 VTAIL.n153 VSUBS 0.079616f
C249 VTAIL.t5 VSUBS 0.058072f
C250 VTAIL.n154 VSUBS 0.019928f
C251 VTAIL.n155 VSUBS 0.016712f
C252 VTAIL.n156 VSUBS 0.011241f
C253 VTAIL.n157 VSUBS 0.271287f
C254 VTAIL.n158 VSUBS 0.02092f
C255 VTAIL.n159 VSUBS 0.011241f
C256 VTAIL.n160 VSUBS 0.011903f
C257 VTAIL.n161 VSUBS 0.02657f
C258 VTAIL.n162 VSUBS 0.059797f
C259 VTAIL.n163 VSUBS 0.011903f
C260 VTAIL.n164 VSUBS 0.011241f
C261 VTAIL.n165 VSUBS 0.047783f
C262 VTAIL.n166 VSUBS 0.029853f
C263 VTAIL.n167 VSUBS 0.625532f
C264 VP.n0 VSUBS 0.045616f
C265 VP.t7 VSUBS 0.298806f
C266 VP.n1 VSUBS 0.161501f
C267 VP.n2 VSUBS 0.045616f
C268 VP.t5 VSUBS 0.298806f
C269 VP.t3 VSUBS 0.298806f
C270 VP.n3 VSUBS 0.19024f
C271 VP.t0 VSUBS 0.298806f
C272 VP.t6 VSUBS 0.315814f
C273 VP.n4 VSUBS 0.145508f
C274 VP.n5 VSUBS 0.1715f
C275 VP.n6 VSUBS 0.161501f
C276 VP.n7 VSUBS 0.010351f
C277 VP.n8 VSUBS 0.16122f
C278 VP.n9 VSUBS 1.37851f
C279 VP.n10 VSUBS 1.42515f
C280 VP.t2 VSUBS 0.298806f
C281 VP.n11 VSUBS 0.16122f
C282 VP.n12 VSUBS 0.010351f
C283 VP.n13 VSUBS 0.045616f
C284 VP.n14 VSUBS 0.045616f
C285 VP.n15 VSUBS 0.045616f
C286 VP.t1 VSUBS 0.298806f
C287 VP.n16 VSUBS 0.161501f
C288 VP.n17 VSUBS 0.010351f
C289 VP.t4 VSUBS 0.298806f
C290 VP.n18 VSUBS 0.16122f
C291 VP.n19 VSUBS 0.035351f
C292 B.n0 VSUBS 0.006564f
C293 B.n1 VSUBS 0.006564f
C294 B.n2 VSUBS 0.009708f
C295 B.n3 VSUBS 0.007439f
C296 B.n4 VSUBS 0.007439f
C297 B.n5 VSUBS 0.007439f
C298 B.n6 VSUBS 0.007439f
C299 B.n7 VSUBS 0.007439f
C300 B.n8 VSUBS 0.007439f
C301 B.n9 VSUBS 0.007439f
C302 B.n10 VSUBS 0.007439f
C303 B.n11 VSUBS 0.007439f
C304 B.n12 VSUBS 0.016181f
C305 B.n13 VSUBS 0.007439f
C306 B.n14 VSUBS 0.007439f
C307 B.n15 VSUBS 0.007439f
C308 B.n16 VSUBS 0.007439f
C309 B.n17 VSUBS 0.007439f
C310 B.n18 VSUBS 0.007439f
C311 B.n19 VSUBS 0.007439f
C312 B.n20 VSUBS 0.007439f
C313 B.n21 VSUBS 0.007439f
C314 B.t1 VSUBS 0.058426f
C315 B.t2 VSUBS 0.065468f
C316 B.t0 VSUBS 0.104255f
C317 B.n22 VSUBS 0.120431f
C318 B.n23 VSUBS 0.110278f
C319 B.n24 VSUBS 0.007439f
C320 B.n25 VSUBS 0.007439f
C321 B.n26 VSUBS 0.007439f
C322 B.n27 VSUBS 0.007439f
C323 B.t4 VSUBS 0.058427f
C324 B.t5 VSUBS 0.065469f
C325 B.t3 VSUBS 0.104255f
C326 B.n28 VSUBS 0.12043f
C327 B.n29 VSUBS 0.110277f
C328 B.n30 VSUBS 0.017236f
C329 B.n31 VSUBS 0.007439f
C330 B.n32 VSUBS 0.007439f
C331 B.n33 VSUBS 0.007439f
C332 B.n34 VSUBS 0.007439f
C333 B.n35 VSUBS 0.007439f
C334 B.n36 VSUBS 0.007439f
C335 B.n37 VSUBS 0.007439f
C336 B.n38 VSUBS 0.007439f
C337 B.n39 VSUBS 0.017296f
C338 B.n40 VSUBS 0.007439f
C339 B.n41 VSUBS 0.007439f
C340 B.n42 VSUBS 0.007439f
C341 B.n43 VSUBS 0.007439f
C342 B.n44 VSUBS 0.007439f
C343 B.n45 VSUBS 0.007439f
C344 B.n46 VSUBS 0.007439f
C345 B.n47 VSUBS 0.007439f
C346 B.n48 VSUBS 0.007439f
C347 B.n49 VSUBS 0.007439f
C348 B.n50 VSUBS 0.007439f
C349 B.n51 VSUBS 0.007439f
C350 B.n52 VSUBS 0.007439f
C351 B.n53 VSUBS 0.007439f
C352 B.n54 VSUBS 0.007439f
C353 B.n55 VSUBS 0.007439f
C354 B.n56 VSUBS 0.007439f
C355 B.n57 VSUBS 0.007439f
C356 B.n58 VSUBS 0.007439f
C357 B.n59 VSUBS 0.007439f
C358 B.n60 VSUBS 0.007439f
C359 B.n61 VSUBS 0.016181f
C360 B.n62 VSUBS 0.007439f
C361 B.n63 VSUBS 0.007439f
C362 B.n64 VSUBS 0.007439f
C363 B.n65 VSUBS 0.007439f
C364 B.n66 VSUBS 0.007439f
C365 B.n67 VSUBS 0.007439f
C366 B.n68 VSUBS 0.007439f
C367 B.n69 VSUBS 0.007439f
C368 B.n70 VSUBS 0.005142f
C369 B.n71 VSUBS 0.007439f
C370 B.n72 VSUBS 0.007439f
C371 B.n73 VSUBS 0.007439f
C372 B.n74 VSUBS 0.007439f
C373 B.n75 VSUBS 0.007439f
C374 B.t8 VSUBS 0.058426f
C375 B.t7 VSUBS 0.065468f
C376 B.t6 VSUBS 0.104255f
C377 B.n76 VSUBS 0.120431f
C378 B.n77 VSUBS 0.110278f
C379 B.n78 VSUBS 0.007439f
C380 B.n79 VSUBS 0.007439f
C381 B.n80 VSUBS 0.007439f
C382 B.n81 VSUBS 0.007439f
C383 B.n82 VSUBS 0.007439f
C384 B.n83 VSUBS 0.007439f
C385 B.n84 VSUBS 0.007439f
C386 B.n85 VSUBS 0.007439f
C387 B.n86 VSUBS 0.016181f
C388 B.n87 VSUBS 0.007439f
C389 B.n88 VSUBS 0.007439f
C390 B.n89 VSUBS 0.007439f
C391 B.n90 VSUBS 0.007439f
C392 B.n91 VSUBS 0.007439f
C393 B.n92 VSUBS 0.007439f
C394 B.n93 VSUBS 0.007439f
C395 B.n94 VSUBS 0.007439f
C396 B.n95 VSUBS 0.007439f
C397 B.n96 VSUBS 0.007439f
C398 B.n97 VSUBS 0.007439f
C399 B.n98 VSUBS 0.007439f
C400 B.n99 VSUBS 0.007439f
C401 B.n100 VSUBS 0.007439f
C402 B.n101 VSUBS 0.007439f
C403 B.n102 VSUBS 0.007439f
C404 B.n103 VSUBS 0.007439f
C405 B.n104 VSUBS 0.007439f
C406 B.n105 VSUBS 0.007439f
C407 B.n106 VSUBS 0.007439f
C408 B.n107 VSUBS 0.007439f
C409 B.n108 VSUBS 0.007439f
C410 B.n109 VSUBS 0.007439f
C411 B.n110 VSUBS 0.007439f
C412 B.n111 VSUBS 0.007439f
C413 B.n112 VSUBS 0.007439f
C414 B.n113 VSUBS 0.007439f
C415 B.n114 VSUBS 0.007439f
C416 B.n115 VSUBS 0.007439f
C417 B.n116 VSUBS 0.007439f
C418 B.n117 VSUBS 0.007439f
C419 B.n118 VSUBS 0.007439f
C420 B.n119 VSUBS 0.007439f
C421 B.n120 VSUBS 0.007439f
C422 B.n121 VSUBS 0.007439f
C423 B.n122 VSUBS 0.007439f
C424 B.n123 VSUBS 0.007439f
C425 B.n124 VSUBS 0.007439f
C426 B.n125 VSUBS 0.016181f
C427 B.n126 VSUBS 0.017296f
C428 B.n127 VSUBS 0.017296f
C429 B.n128 VSUBS 0.007439f
C430 B.n129 VSUBS 0.007439f
C431 B.n130 VSUBS 0.007439f
C432 B.n131 VSUBS 0.007439f
C433 B.n132 VSUBS 0.007439f
C434 B.n133 VSUBS 0.007439f
C435 B.n134 VSUBS 0.007439f
C436 B.n135 VSUBS 0.007439f
C437 B.n136 VSUBS 0.007439f
C438 B.n137 VSUBS 0.007439f
C439 B.n138 VSUBS 0.007439f
C440 B.n139 VSUBS 0.007439f
C441 B.n140 VSUBS 0.007439f
C442 B.n141 VSUBS 0.007439f
C443 B.n142 VSUBS 0.007439f
C444 B.n143 VSUBS 0.007439f
C445 B.n144 VSUBS 0.007439f
C446 B.n145 VSUBS 0.007439f
C447 B.n146 VSUBS 0.007439f
C448 B.n147 VSUBS 0.007439f
C449 B.n148 VSUBS 0.007439f
C450 B.n149 VSUBS 0.007439f
C451 B.n150 VSUBS 0.007439f
C452 B.n151 VSUBS 0.007439f
C453 B.n152 VSUBS 0.005142f
C454 B.n153 VSUBS 0.017236f
C455 B.n154 VSUBS 0.006017f
C456 B.n155 VSUBS 0.007439f
C457 B.n156 VSUBS 0.007439f
C458 B.n157 VSUBS 0.007439f
C459 B.n158 VSUBS 0.007439f
C460 B.n159 VSUBS 0.007439f
C461 B.n160 VSUBS 0.007439f
C462 B.n161 VSUBS 0.007439f
C463 B.n162 VSUBS 0.007439f
C464 B.n163 VSUBS 0.007439f
C465 B.n164 VSUBS 0.007439f
C466 B.n165 VSUBS 0.007439f
C467 B.t11 VSUBS 0.058427f
C468 B.t10 VSUBS 0.065469f
C469 B.t9 VSUBS 0.104255f
C470 B.n166 VSUBS 0.12043f
C471 B.n167 VSUBS 0.110277f
C472 B.n168 VSUBS 0.017236f
C473 B.n169 VSUBS 0.006017f
C474 B.n170 VSUBS 0.007439f
C475 B.n171 VSUBS 0.007439f
C476 B.n172 VSUBS 0.007439f
C477 B.n173 VSUBS 0.007439f
C478 B.n174 VSUBS 0.007439f
C479 B.n175 VSUBS 0.007439f
C480 B.n176 VSUBS 0.007439f
C481 B.n177 VSUBS 0.007439f
C482 B.n178 VSUBS 0.007439f
C483 B.n179 VSUBS 0.007439f
C484 B.n180 VSUBS 0.007439f
C485 B.n181 VSUBS 0.007439f
C486 B.n182 VSUBS 0.007439f
C487 B.n183 VSUBS 0.007439f
C488 B.n184 VSUBS 0.007439f
C489 B.n185 VSUBS 0.007439f
C490 B.n186 VSUBS 0.007439f
C491 B.n187 VSUBS 0.007439f
C492 B.n188 VSUBS 0.007439f
C493 B.n189 VSUBS 0.007439f
C494 B.n190 VSUBS 0.007439f
C495 B.n191 VSUBS 0.007439f
C496 B.n192 VSUBS 0.007439f
C497 B.n193 VSUBS 0.007439f
C498 B.n194 VSUBS 0.007439f
C499 B.n195 VSUBS 0.007439f
C500 B.n196 VSUBS 0.017296f
C501 B.n197 VSUBS 0.016363f
C502 B.n198 VSUBS 0.017114f
C503 B.n199 VSUBS 0.007439f
C504 B.n200 VSUBS 0.007439f
C505 B.n201 VSUBS 0.007439f
C506 B.n202 VSUBS 0.007439f
C507 B.n203 VSUBS 0.007439f
C508 B.n204 VSUBS 0.007439f
C509 B.n205 VSUBS 0.007439f
C510 B.n206 VSUBS 0.007439f
C511 B.n207 VSUBS 0.007439f
C512 B.n208 VSUBS 0.007439f
C513 B.n209 VSUBS 0.007439f
C514 B.n210 VSUBS 0.007439f
C515 B.n211 VSUBS 0.007439f
C516 B.n212 VSUBS 0.007439f
C517 B.n213 VSUBS 0.007439f
C518 B.n214 VSUBS 0.007439f
C519 B.n215 VSUBS 0.007439f
C520 B.n216 VSUBS 0.007439f
C521 B.n217 VSUBS 0.007439f
C522 B.n218 VSUBS 0.007439f
C523 B.n219 VSUBS 0.007439f
C524 B.n220 VSUBS 0.007439f
C525 B.n221 VSUBS 0.007439f
C526 B.n222 VSUBS 0.007439f
C527 B.n223 VSUBS 0.007439f
C528 B.n224 VSUBS 0.007439f
C529 B.n225 VSUBS 0.007439f
C530 B.n226 VSUBS 0.007439f
C531 B.n227 VSUBS 0.007439f
C532 B.n228 VSUBS 0.007439f
C533 B.n229 VSUBS 0.007439f
C534 B.n230 VSUBS 0.007439f
C535 B.n231 VSUBS 0.007439f
C536 B.n232 VSUBS 0.007439f
C537 B.n233 VSUBS 0.007439f
C538 B.n234 VSUBS 0.007439f
C539 B.n235 VSUBS 0.007439f
C540 B.n236 VSUBS 0.007439f
C541 B.n237 VSUBS 0.007439f
C542 B.n238 VSUBS 0.007439f
C543 B.n239 VSUBS 0.007439f
C544 B.n240 VSUBS 0.007439f
C545 B.n241 VSUBS 0.007439f
C546 B.n242 VSUBS 0.007439f
C547 B.n243 VSUBS 0.007439f
C548 B.n244 VSUBS 0.007439f
C549 B.n245 VSUBS 0.007439f
C550 B.n246 VSUBS 0.007439f
C551 B.n247 VSUBS 0.007439f
C552 B.n248 VSUBS 0.007439f
C553 B.n249 VSUBS 0.007439f
C554 B.n250 VSUBS 0.007439f
C555 B.n251 VSUBS 0.007439f
C556 B.n252 VSUBS 0.007439f
C557 B.n253 VSUBS 0.007439f
C558 B.n254 VSUBS 0.007439f
C559 B.n255 VSUBS 0.007439f
C560 B.n256 VSUBS 0.007439f
C561 B.n257 VSUBS 0.007439f
C562 B.n258 VSUBS 0.007439f
C563 B.n259 VSUBS 0.007439f
C564 B.n260 VSUBS 0.007439f
C565 B.n261 VSUBS 0.007439f
C566 B.n262 VSUBS 0.016181f
C567 B.n263 VSUBS 0.016181f
C568 B.n264 VSUBS 0.017296f
C569 B.n265 VSUBS 0.007439f
C570 B.n266 VSUBS 0.007439f
C571 B.n267 VSUBS 0.007439f
C572 B.n268 VSUBS 0.007439f
C573 B.n269 VSUBS 0.007439f
C574 B.n270 VSUBS 0.007439f
C575 B.n271 VSUBS 0.007439f
C576 B.n272 VSUBS 0.007439f
C577 B.n273 VSUBS 0.007439f
C578 B.n274 VSUBS 0.007439f
C579 B.n275 VSUBS 0.007439f
C580 B.n276 VSUBS 0.007439f
C581 B.n277 VSUBS 0.007439f
C582 B.n278 VSUBS 0.007439f
C583 B.n279 VSUBS 0.007439f
C584 B.n280 VSUBS 0.007439f
C585 B.n281 VSUBS 0.007439f
C586 B.n282 VSUBS 0.007439f
C587 B.n283 VSUBS 0.007439f
C588 B.n284 VSUBS 0.007439f
C589 B.n285 VSUBS 0.007439f
C590 B.n286 VSUBS 0.007439f
C591 B.n287 VSUBS 0.007439f
C592 B.n288 VSUBS 0.007439f
C593 B.n289 VSUBS 0.005142f
C594 B.n290 VSUBS 0.007439f
C595 B.n291 VSUBS 0.007439f
C596 B.n292 VSUBS 0.006017f
C597 B.n293 VSUBS 0.007439f
C598 B.n294 VSUBS 0.007439f
C599 B.n295 VSUBS 0.007439f
C600 B.n296 VSUBS 0.007439f
C601 B.n297 VSUBS 0.007439f
C602 B.n298 VSUBS 0.007439f
C603 B.n299 VSUBS 0.007439f
C604 B.n300 VSUBS 0.007439f
C605 B.n301 VSUBS 0.007439f
C606 B.n302 VSUBS 0.007439f
C607 B.n303 VSUBS 0.007439f
C608 B.n304 VSUBS 0.006017f
C609 B.n305 VSUBS 0.017236f
C610 B.n306 VSUBS 0.005142f
C611 B.n307 VSUBS 0.007439f
C612 B.n308 VSUBS 0.007439f
C613 B.n309 VSUBS 0.007439f
C614 B.n310 VSUBS 0.007439f
C615 B.n311 VSUBS 0.007439f
C616 B.n312 VSUBS 0.007439f
C617 B.n313 VSUBS 0.007439f
C618 B.n314 VSUBS 0.007439f
C619 B.n315 VSUBS 0.007439f
C620 B.n316 VSUBS 0.007439f
C621 B.n317 VSUBS 0.007439f
C622 B.n318 VSUBS 0.007439f
C623 B.n319 VSUBS 0.007439f
C624 B.n320 VSUBS 0.007439f
C625 B.n321 VSUBS 0.007439f
C626 B.n322 VSUBS 0.007439f
C627 B.n323 VSUBS 0.007439f
C628 B.n324 VSUBS 0.007439f
C629 B.n325 VSUBS 0.007439f
C630 B.n326 VSUBS 0.007439f
C631 B.n327 VSUBS 0.007439f
C632 B.n328 VSUBS 0.007439f
C633 B.n329 VSUBS 0.007439f
C634 B.n330 VSUBS 0.007439f
C635 B.n331 VSUBS 0.017296f
C636 B.n332 VSUBS 0.017296f
C637 B.n333 VSUBS 0.016181f
C638 B.n334 VSUBS 0.007439f
C639 B.n335 VSUBS 0.007439f
C640 B.n336 VSUBS 0.007439f
C641 B.n337 VSUBS 0.007439f
C642 B.n338 VSUBS 0.007439f
C643 B.n339 VSUBS 0.007439f
C644 B.n340 VSUBS 0.007439f
C645 B.n341 VSUBS 0.007439f
C646 B.n342 VSUBS 0.007439f
C647 B.n343 VSUBS 0.007439f
C648 B.n344 VSUBS 0.007439f
C649 B.n345 VSUBS 0.007439f
C650 B.n346 VSUBS 0.007439f
C651 B.n347 VSUBS 0.007439f
C652 B.n348 VSUBS 0.007439f
C653 B.n349 VSUBS 0.007439f
C654 B.n350 VSUBS 0.007439f
C655 B.n351 VSUBS 0.007439f
C656 B.n352 VSUBS 0.007439f
C657 B.n353 VSUBS 0.007439f
C658 B.n354 VSUBS 0.007439f
C659 B.n355 VSUBS 0.007439f
C660 B.n356 VSUBS 0.007439f
C661 B.n357 VSUBS 0.007439f
C662 B.n358 VSUBS 0.007439f
C663 B.n359 VSUBS 0.007439f
C664 B.n360 VSUBS 0.007439f
C665 B.n361 VSUBS 0.007439f
C666 B.n362 VSUBS 0.007439f
C667 B.n363 VSUBS 0.009708f
C668 B.n364 VSUBS 0.010341f
C669 B.n365 VSUBS 0.020565f
.ends

