* NGSPICE file created from diff_pair_sample_0904.ext - technology: sky130A

.subckt diff_pair_sample_0904 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t1 VP.t0 VTAIL.t2 w_n1610_n3824# sky130_fd_pr__pfet_01v8 ad=5.5692 pd=29.34 as=5.5692 ps=29.34 w=14.28 l=1.27
X1 VDD1.t0 VP.t1 VTAIL.t3 w_n1610_n3824# sky130_fd_pr__pfet_01v8 ad=5.5692 pd=29.34 as=5.5692 ps=29.34 w=14.28 l=1.27
X2 B.t11 B.t9 B.t10 w_n1610_n3824# sky130_fd_pr__pfet_01v8 ad=5.5692 pd=29.34 as=0 ps=0 w=14.28 l=1.27
X3 B.t8 B.t6 B.t7 w_n1610_n3824# sky130_fd_pr__pfet_01v8 ad=5.5692 pd=29.34 as=0 ps=0 w=14.28 l=1.27
X4 VDD2.t1 VN.t0 VTAIL.t1 w_n1610_n3824# sky130_fd_pr__pfet_01v8 ad=5.5692 pd=29.34 as=5.5692 ps=29.34 w=14.28 l=1.27
X5 B.t5 B.t3 B.t4 w_n1610_n3824# sky130_fd_pr__pfet_01v8 ad=5.5692 pd=29.34 as=0 ps=0 w=14.28 l=1.27
X6 B.t2 B.t0 B.t1 w_n1610_n3824# sky130_fd_pr__pfet_01v8 ad=5.5692 pd=29.34 as=0 ps=0 w=14.28 l=1.27
X7 VDD2.t0 VN.t1 VTAIL.t0 w_n1610_n3824# sky130_fd_pr__pfet_01v8 ad=5.5692 pd=29.34 as=5.5692 ps=29.34 w=14.28 l=1.27
R0 VP.n0 VP.t1 425.375
R1 VP.n0 VP.t0 382.517
R2 VP VP.n0 0.146778
R3 VTAIL.n306 VTAIL.n234 756.745
R4 VTAIL.n72 VTAIL.n0 756.745
R5 VTAIL.n228 VTAIL.n156 756.745
R6 VTAIL.n150 VTAIL.n78 756.745
R7 VTAIL.n258 VTAIL.n257 585
R8 VTAIL.n263 VTAIL.n262 585
R9 VTAIL.n265 VTAIL.n264 585
R10 VTAIL.n254 VTAIL.n253 585
R11 VTAIL.n271 VTAIL.n270 585
R12 VTAIL.n273 VTAIL.n272 585
R13 VTAIL.n250 VTAIL.n249 585
R14 VTAIL.n280 VTAIL.n279 585
R15 VTAIL.n281 VTAIL.n248 585
R16 VTAIL.n283 VTAIL.n282 585
R17 VTAIL.n246 VTAIL.n245 585
R18 VTAIL.n289 VTAIL.n288 585
R19 VTAIL.n291 VTAIL.n290 585
R20 VTAIL.n242 VTAIL.n241 585
R21 VTAIL.n297 VTAIL.n296 585
R22 VTAIL.n299 VTAIL.n298 585
R23 VTAIL.n238 VTAIL.n237 585
R24 VTAIL.n305 VTAIL.n304 585
R25 VTAIL.n307 VTAIL.n306 585
R26 VTAIL.n24 VTAIL.n23 585
R27 VTAIL.n29 VTAIL.n28 585
R28 VTAIL.n31 VTAIL.n30 585
R29 VTAIL.n20 VTAIL.n19 585
R30 VTAIL.n37 VTAIL.n36 585
R31 VTAIL.n39 VTAIL.n38 585
R32 VTAIL.n16 VTAIL.n15 585
R33 VTAIL.n46 VTAIL.n45 585
R34 VTAIL.n47 VTAIL.n14 585
R35 VTAIL.n49 VTAIL.n48 585
R36 VTAIL.n12 VTAIL.n11 585
R37 VTAIL.n55 VTAIL.n54 585
R38 VTAIL.n57 VTAIL.n56 585
R39 VTAIL.n8 VTAIL.n7 585
R40 VTAIL.n63 VTAIL.n62 585
R41 VTAIL.n65 VTAIL.n64 585
R42 VTAIL.n4 VTAIL.n3 585
R43 VTAIL.n71 VTAIL.n70 585
R44 VTAIL.n73 VTAIL.n72 585
R45 VTAIL.n229 VTAIL.n228 585
R46 VTAIL.n227 VTAIL.n226 585
R47 VTAIL.n160 VTAIL.n159 585
R48 VTAIL.n221 VTAIL.n220 585
R49 VTAIL.n219 VTAIL.n218 585
R50 VTAIL.n164 VTAIL.n163 585
R51 VTAIL.n213 VTAIL.n212 585
R52 VTAIL.n211 VTAIL.n210 585
R53 VTAIL.n168 VTAIL.n167 585
R54 VTAIL.n205 VTAIL.n204 585
R55 VTAIL.n203 VTAIL.n170 585
R56 VTAIL.n202 VTAIL.n201 585
R57 VTAIL.n173 VTAIL.n171 585
R58 VTAIL.n196 VTAIL.n195 585
R59 VTAIL.n194 VTAIL.n193 585
R60 VTAIL.n177 VTAIL.n176 585
R61 VTAIL.n188 VTAIL.n187 585
R62 VTAIL.n186 VTAIL.n185 585
R63 VTAIL.n181 VTAIL.n180 585
R64 VTAIL.n151 VTAIL.n150 585
R65 VTAIL.n149 VTAIL.n148 585
R66 VTAIL.n82 VTAIL.n81 585
R67 VTAIL.n143 VTAIL.n142 585
R68 VTAIL.n141 VTAIL.n140 585
R69 VTAIL.n86 VTAIL.n85 585
R70 VTAIL.n135 VTAIL.n134 585
R71 VTAIL.n133 VTAIL.n132 585
R72 VTAIL.n90 VTAIL.n89 585
R73 VTAIL.n127 VTAIL.n126 585
R74 VTAIL.n125 VTAIL.n92 585
R75 VTAIL.n124 VTAIL.n123 585
R76 VTAIL.n95 VTAIL.n93 585
R77 VTAIL.n118 VTAIL.n117 585
R78 VTAIL.n116 VTAIL.n115 585
R79 VTAIL.n99 VTAIL.n98 585
R80 VTAIL.n110 VTAIL.n109 585
R81 VTAIL.n108 VTAIL.n107 585
R82 VTAIL.n103 VTAIL.n102 585
R83 VTAIL.n259 VTAIL.t0 329.036
R84 VTAIL.n25 VTAIL.t2 329.036
R85 VTAIL.n104 VTAIL.t1 329.036
R86 VTAIL.n182 VTAIL.t3 329.036
R87 VTAIL.n263 VTAIL.n257 171.744
R88 VTAIL.n264 VTAIL.n263 171.744
R89 VTAIL.n264 VTAIL.n253 171.744
R90 VTAIL.n271 VTAIL.n253 171.744
R91 VTAIL.n272 VTAIL.n271 171.744
R92 VTAIL.n272 VTAIL.n249 171.744
R93 VTAIL.n280 VTAIL.n249 171.744
R94 VTAIL.n281 VTAIL.n280 171.744
R95 VTAIL.n282 VTAIL.n281 171.744
R96 VTAIL.n282 VTAIL.n245 171.744
R97 VTAIL.n289 VTAIL.n245 171.744
R98 VTAIL.n290 VTAIL.n289 171.744
R99 VTAIL.n290 VTAIL.n241 171.744
R100 VTAIL.n297 VTAIL.n241 171.744
R101 VTAIL.n298 VTAIL.n297 171.744
R102 VTAIL.n298 VTAIL.n237 171.744
R103 VTAIL.n305 VTAIL.n237 171.744
R104 VTAIL.n306 VTAIL.n305 171.744
R105 VTAIL.n29 VTAIL.n23 171.744
R106 VTAIL.n30 VTAIL.n29 171.744
R107 VTAIL.n30 VTAIL.n19 171.744
R108 VTAIL.n37 VTAIL.n19 171.744
R109 VTAIL.n38 VTAIL.n37 171.744
R110 VTAIL.n38 VTAIL.n15 171.744
R111 VTAIL.n46 VTAIL.n15 171.744
R112 VTAIL.n47 VTAIL.n46 171.744
R113 VTAIL.n48 VTAIL.n47 171.744
R114 VTAIL.n48 VTAIL.n11 171.744
R115 VTAIL.n55 VTAIL.n11 171.744
R116 VTAIL.n56 VTAIL.n55 171.744
R117 VTAIL.n56 VTAIL.n7 171.744
R118 VTAIL.n63 VTAIL.n7 171.744
R119 VTAIL.n64 VTAIL.n63 171.744
R120 VTAIL.n64 VTAIL.n3 171.744
R121 VTAIL.n71 VTAIL.n3 171.744
R122 VTAIL.n72 VTAIL.n71 171.744
R123 VTAIL.n228 VTAIL.n227 171.744
R124 VTAIL.n227 VTAIL.n159 171.744
R125 VTAIL.n220 VTAIL.n159 171.744
R126 VTAIL.n220 VTAIL.n219 171.744
R127 VTAIL.n219 VTAIL.n163 171.744
R128 VTAIL.n212 VTAIL.n163 171.744
R129 VTAIL.n212 VTAIL.n211 171.744
R130 VTAIL.n211 VTAIL.n167 171.744
R131 VTAIL.n204 VTAIL.n167 171.744
R132 VTAIL.n204 VTAIL.n203 171.744
R133 VTAIL.n203 VTAIL.n202 171.744
R134 VTAIL.n202 VTAIL.n171 171.744
R135 VTAIL.n195 VTAIL.n171 171.744
R136 VTAIL.n195 VTAIL.n194 171.744
R137 VTAIL.n194 VTAIL.n176 171.744
R138 VTAIL.n187 VTAIL.n176 171.744
R139 VTAIL.n187 VTAIL.n186 171.744
R140 VTAIL.n186 VTAIL.n180 171.744
R141 VTAIL.n150 VTAIL.n149 171.744
R142 VTAIL.n149 VTAIL.n81 171.744
R143 VTAIL.n142 VTAIL.n81 171.744
R144 VTAIL.n142 VTAIL.n141 171.744
R145 VTAIL.n141 VTAIL.n85 171.744
R146 VTAIL.n134 VTAIL.n85 171.744
R147 VTAIL.n134 VTAIL.n133 171.744
R148 VTAIL.n133 VTAIL.n89 171.744
R149 VTAIL.n126 VTAIL.n89 171.744
R150 VTAIL.n126 VTAIL.n125 171.744
R151 VTAIL.n125 VTAIL.n124 171.744
R152 VTAIL.n124 VTAIL.n93 171.744
R153 VTAIL.n117 VTAIL.n93 171.744
R154 VTAIL.n117 VTAIL.n116 171.744
R155 VTAIL.n116 VTAIL.n98 171.744
R156 VTAIL.n109 VTAIL.n98 171.744
R157 VTAIL.n109 VTAIL.n108 171.744
R158 VTAIL.n108 VTAIL.n102 171.744
R159 VTAIL.t0 VTAIL.n257 85.8723
R160 VTAIL.t2 VTAIL.n23 85.8723
R161 VTAIL.t3 VTAIL.n180 85.8723
R162 VTAIL.t1 VTAIL.n102 85.8723
R163 VTAIL.n311 VTAIL.n310 32.1853
R164 VTAIL.n77 VTAIL.n76 32.1853
R165 VTAIL.n233 VTAIL.n232 32.1853
R166 VTAIL.n155 VTAIL.n154 32.1853
R167 VTAIL.n155 VTAIL.n77 27.4358
R168 VTAIL.n311 VTAIL.n233 26.0565
R169 VTAIL.n283 VTAIL.n248 13.1884
R170 VTAIL.n49 VTAIL.n14 13.1884
R171 VTAIL.n205 VTAIL.n170 13.1884
R172 VTAIL.n127 VTAIL.n92 13.1884
R173 VTAIL.n279 VTAIL.n278 12.8005
R174 VTAIL.n284 VTAIL.n246 12.8005
R175 VTAIL.n45 VTAIL.n44 12.8005
R176 VTAIL.n50 VTAIL.n12 12.8005
R177 VTAIL.n206 VTAIL.n168 12.8005
R178 VTAIL.n201 VTAIL.n172 12.8005
R179 VTAIL.n128 VTAIL.n90 12.8005
R180 VTAIL.n123 VTAIL.n94 12.8005
R181 VTAIL.n277 VTAIL.n250 12.0247
R182 VTAIL.n288 VTAIL.n287 12.0247
R183 VTAIL.n43 VTAIL.n16 12.0247
R184 VTAIL.n54 VTAIL.n53 12.0247
R185 VTAIL.n210 VTAIL.n209 12.0247
R186 VTAIL.n200 VTAIL.n173 12.0247
R187 VTAIL.n132 VTAIL.n131 12.0247
R188 VTAIL.n122 VTAIL.n95 12.0247
R189 VTAIL.n274 VTAIL.n273 11.249
R190 VTAIL.n291 VTAIL.n244 11.249
R191 VTAIL.n40 VTAIL.n39 11.249
R192 VTAIL.n57 VTAIL.n10 11.249
R193 VTAIL.n213 VTAIL.n166 11.249
R194 VTAIL.n197 VTAIL.n196 11.249
R195 VTAIL.n135 VTAIL.n88 11.249
R196 VTAIL.n119 VTAIL.n118 11.249
R197 VTAIL.n259 VTAIL.n258 10.7239
R198 VTAIL.n25 VTAIL.n24 10.7239
R199 VTAIL.n182 VTAIL.n181 10.7239
R200 VTAIL.n104 VTAIL.n103 10.7239
R201 VTAIL.n270 VTAIL.n252 10.4732
R202 VTAIL.n292 VTAIL.n242 10.4732
R203 VTAIL.n36 VTAIL.n18 10.4732
R204 VTAIL.n58 VTAIL.n8 10.4732
R205 VTAIL.n214 VTAIL.n164 10.4732
R206 VTAIL.n193 VTAIL.n175 10.4732
R207 VTAIL.n136 VTAIL.n86 10.4732
R208 VTAIL.n115 VTAIL.n97 10.4732
R209 VTAIL.n269 VTAIL.n254 9.69747
R210 VTAIL.n296 VTAIL.n295 9.69747
R211 VTAIL.n35 VTAIL.n20 9.69747
R212 VTAIL.n62 VTAIL.n61 9.69747
R213 VTAIL.n218 VTAIL.n217 9.69747
R214 VTAIL.n192 VTAIL.n177 9.69747
R215 VTAIL.n140 VTAIL.n139 9.69747
R216 VTAIL.n114 VTAIL.n99 9.69747
R217 VTAIL.n310 VTAIL.n309 9.45567
R218 VTAIL.n76 VTAIL.n75 9.45567
R219 VTAIL.n232 VTAIL.n231 9.45567
R220 VTAIL.n154 VTAIL.n153 9.45567
R221 VTAIL.n236 VTAIL.n235 9.3005
R222 VTAIL.n309 VTAIL.n308 9.3005
R223 VTAIL.n301 VTAIL.n300 9.3005
R224 VTAIL.n240 VTAIL.n239 9.3005
R225 VTAIL.n295 VTAIL.n294 9.3005
R226 VTAIL.n293 VTAIL.n292 9.3005
R227 VTAIL.n244 VTAIL.n243 9.3005
R228 VTAIL.n287 VTAIL.n286 9.3005
R229 VTAIL.n285 VTAIL.n284 9.3005
R230 VTAIL.n261 VTAIL.n260 9.3005
R231 VTAIL.n256 VTAIL.n255 9.3005
R232 VTAIL.n267 VTAIL.n266 9.3005
R233 VTAIL.n269 VTAIL.n268 9.3005
R234 VTAIL.n252 VTAIL.n251 9.3005
R235 VTAIL.n275 VTAIL.n274 9.3005
R236 VTAIL.n277 VTAIL.n276 9.3005
R237 VTAIL.n278 VTAIL.n247 9.3005
R238 VTAIL.n303 VTAIL.n302 9.3005
R239 VTAIL.n2 VTAIL.n1 9.3005
R240 VTAIL.n75 VTAIL.n74 9.3005
R241 VTAIL.n67 VTAIL.n66 9.3005
R242 VTAIL.n6 VTAIL.n5 9.3005
R243 VTAIL.n61 VTAIL.n60 9.3005
R244 VTAIL.n59 VTAIL.n58 9.3005
R245 VTAIL.n10 VTAIL.n9 9.3005
R246 VTAIL.n53 VTAIL.n52 9.3005
R247 VTAIL.n51 VTAIL.n50 9.3005
R248 VTAIL.n27 VTAIL.n26 9.3005
R249 VTAIL.n22 VTAIL.n21 9.3005
R250 VTAIL.n33 VTAIL.n32 9.3005
R251 VTAIL.n35 VTAIL.n34 9.3005
R252 VTAIL.n18 VTAIL.n17 9.3005
R253 VTAIL.n41 VTAIL.n40 9.3005
R254 VTAIL.n43 VTAIL.n42 9.3005
R255 VTAIL.n44 VTAIL.n13 9.3005
R256 VTAIL.n69 VTAIL.n68 9.3005
R257 VTAIL.n158 VTAIL.n157 9.3005
R258 VTAIL.n225 VTAIL.n224 9.3005
R259 VTAIL.n223 VTAIL.n222 9.3005
R260 VTAIL.n162 VTAIL.n161 9.3005
R261 VTAIL.n217 VTAIL.n216 9.3005
R262 VTAIL.n215 VTAIL.n214 9.3005
R263 VTAIL.n166 VTAIL.n165 9.3005
R264 VTAIL.n209 VTAIL.n208 9.3005
R265 VTAIL.n207 VTAIL.n206 9.3005
R266 VTAIL.n172 VTAIL.n169 9.3005
R267 VTAIL.n200 VTAIL.n199 9.3005
R268 VTAIL.n198 VTAIL.n197 9.3005
R269 VTAIL.n175 VTAIL.n174 9.3005
R270 VTAIL.n192 VTAIL.n191 9.3005
R271 VTAIL.n190 VTAIL.n189 9.3005
R272 VTAIL.n179 VTAIL.n178 9.3005
R273 VTAIL.n184 VTAIL.n183 9.3005
R274 VTAIL.n231 VTAIL.n230 9.3005
R275 VTAIL.n106 VTAIL.n105 9.3005
R276 VTAIL.n101 VTAIL.n100 9.3005
R277 VTAIL.n112 VTAIL.n111 9.3005
R278 VTAIL.n114 VTAIL.n113 9.3005
R279 VTAIL.n97 VTAIL.n96 9.3005
R280 VTAIL.n120 VTAIL.n119 9.3005
R281 VTAIL.n122 VTAIL.n121 9.3005
R282 VTAIL.n94 VTAIL.n91 9.3005
R283 VTAIL.n153 VTAIL.n152 9.3005
R284 VTAIL.n80 VTAIL.n79 9.3005
R285 VTAIL.n147 VTAIL.n146 9.3005
R286 VTAIL.n145 VTAIL.n144 9.3005
R287 VTAIL.n84 VTAIL.n83 9.3005
R288 VTAIL.n139 VTAIL.n138 9.3005
R289 VTAIL.n137 VTAIL.n136 9.3005
R290 VTAIL.n88 VTAIL.n87 9.3005
R291 VTAIL.n131 VTAIL.n130 9.3005
R292 VTAIL.n129 VTAIL.n128 9.3005
R293 VTAIL.n266 VTAIL.n265 8.92171
R294 VTAIL.n299 VTAIL.n240 8.92171
R295 VTAIL.n32 VTAIL.n31 8.92171
R296 VTAIL.n65 VTAIL.n6 8.92171
R297 VTAIL.n221 VTAIL.n162 8.92171
R298 VTAIL.n189 VTAIL.n188 8.92171
R299 VTAIL.n143 VTAIL.n84 8.92171
R300 VTAIL.n111 VTAIL.n110 8.92171
R301 VTAIL.n262 VTAIL.n256 8.14595
R302 VTAIL.n300 VTAIL.n238 8.14595
R303 VTAIL.n310 VTAIL.n234 8.14595
R304 VTAIL.n28 VTAIL.n22 8.14595
R305 VTAIL.n66 VTAIL.n4 8.14595
R306 VTAIL.n76 VTAIL.n0 8.14595
R307 VTAIL.n232 VTAIL.n156 8.14595
R308 VTAIL.n222 VTAIL.n160 8.14595
R309 VTAIL.n185 VTAIL.n179 8.14595
R310 VTAIL.n154 VTAIL.n78 8.14595
R311 VTAIL.n144 VTAIL.n82 8.14595
R312 VTAIL.n107 VTAIL.n101 8.14595
R313 VTAIL.n261 VTAIL.n258 7.3702
R314 VTAIL.n304 VTAIL.n303 7.3702
R315 VTAIL.n308 VTAIL.n307 7.3702
R316 VTAIL.n27 VTAIL.n24 7.3702
R317 VTAIL.n70 VTAIL.n69 7.3702
R318 VTAIL.n74 VTAIL.n73 7.3702
R319 VTAIL.n230 VTAIL.n229 7.3702
R320 VTAIL.n226 VTAIL.n225 7.3702
R321 VTAIL.n184 VTAIL.n181 7.3702
R322 VTAIL.n152 VTAIL.n151 7.3702
R323 VTAIL.n148 VTAIL.n147 7.3702
R324 VTAIL.n106 VTAIL.n103 7.3702
R325 VTAIL.n304 VTAIL.n236 6.59444
R326 VTAIL.n307 VTAIL.n236 6.59444
R327 VTAIL.n70 VTAIL.n2 6.59444
R328 VTAIL.n73 VTAIL.n2 6.59444
R329 VTAIL.n229 VTAIL.n158 6.59444
R330 VTAIL.n226 VTAIL.n158 6.59444
R331 VTAIL.n151 VTAIL.n80 6.59444
R332 VTAIL.n148 VTAIL.n80 6.59444
R333 VTAIL.n262 VTAIL.n261 5.81868
R334 VTAIL.n303 VTAIL.n238 5.81868
R335 VTAIL.n308 VTAIL.n234 5.81868
R336 VTAIL.n28 VTAIL.n27 5.81868
R337 VTAIL.n69 VTAIL.n4 5.81868
R338 VTAIL.n74 VTAIL.n0 5.81868
R339 VTAIL.n230 VTAIL.n156 5.81868
R340 VTAIL.n225 VTAIL.n160 5.81868
R341 VTAIL.n185 VTAIL.n184 5.81868
R342 VTAIL.n152 VTAIL.n78 5.81868
R343 VTAIL.n147 VTAIL.n82 5.81868
R344 VTAIL.n107 VTAIL.n106 5.81868
R345 VTAIL.n265 VTAIL.n256 5.04292
R346 VTAIL.n300 VTAIL.n299 5.04292
R347 VTAIL.n31 VTAIL.n22 5.04292
R348 VTAIL.n66 VTAIL.n65 5.04292
R349 VTAIL.n222 VTAIL.n221 5.04292
R350 VTAIL.n188 VTAIL.n179 5.04292
R351 VTAIL.n144 VTAIL.n143 5.04292
R352 VTAIL.n110 VTAIL.n101 5.04292
R353 VTAIL.n266 VTAIL.n254 4.26717
R354 VTAIL.n296 VTAIL.n240 4.26717
R355 VTAIL.n32 VTAIL.n20 4.26717
R356 VTAIL.n62 VTAIL.n6 4.26717
R357 VTAIL.n218 VTAIL.n162 4.26717
R358 VTAIL.n189 VTAIL.n177 4.26717
R359 VTAIL.n140 VTAIL.n84 4.26717
R360 VTAIL.n111 VTAIL.n99 4.26717
R361 VTAIL.n270 VTAIL.n269 3.49141
R362 VTAIL.n295 VTAIL.n242 3.49141
R363 VTAIL.n36 VTAIL.n35 3.49141
R364 VTAIL.n61 VTAIL.n8 3.49141
R365 VTAIL.n217 VTAIL.n164 3.49141
R366 VTAIL.n193 VTAIL.n192 3.49141
R367 VTAIL.n139 VTAIL.n86 3.49141
R368 VTAIL.n115 VTAIL.n114 3.49141
R369 VTAIL.n273 VTAIL.n252 2.71565
R370 VTAIL.n292 VTAIL.n291 2.71565
R371 VTAIL.n39 VTAIL.n18 2.71565
R372 VTAIL.n58 VTAIL.n57 2.71565
R373 VTAIL.n214 VTAIL.n213 2.71565
R374 VTAIL.n196 VTAIL.n175 2.71565
R375 VTAIL.n136 VTAIL.n135 2.71565
R376 VTAIL.n118 VTAIL.n97 2.71565
R377 VTAIL.n183 VTAIL.n182 2.41282
R378 VTAIL.n105 VTAIL.n104 2.41282
R379 VTAIL.n260 VTAIL.n259 2.41282
R380 VTAIL.n26 VTAIL.n25 2.41282
R381 VTAIL.n274 VTAIL.n250 1.93989
R382 VTAIL.n288 VTAIL.n244 1.93989
R383 VTAIL.n40 VTAIL.n16 1.93989
R384 VTAIL.n54 VTAIL.n10 1.93989
R385 VTAIL.n210 VTAIL.n166 1.93989
R386 VTAIL.n197 VTAIL.n173 1.93989
R387 VTAIL.n132 VTAIL.n88 1.93989
R388 VTAIL.n119 VTAIL.n95 1.93989
R389 VTAIL.n279 VTAIL.n277 1.16414
R390 VTAIL.n287 VTAIL.n246 1.16414
R391 VTAIL.n45 VTAIL.n43 1.16414
R392 VTAIL.n53 VTAIL.n12 1.16414
R393 VTAIL.n209 VTAIL.n168 1.16414
R394 VTAIL.n201 VTAIL.n200 1.16414
R395 VTAIL.n131 VTAIL.n90 1.16414
R396 VTAIL.n123 VTAIL.n122 1.16414
R397 VTAIL.n233 VTAIL.n155 1.15998
R398 VTAIL VTAIL.n77 0.873345
R399 VTAIL.n278 VTAIL.n248 0.388379
R400 VTAIL.n284 VTAIL.n283 0.388379
R401 VTAIL.n44 VTAIL.n14 0.388379
R402 VTAIL.n50 VTAIL.n49 0.388379
R403 VTAIL.n206 VTAIL.n205 0.388379
R404 VTAIL.n172 VTAIL.n170 0.388379
R405 VTAIL.n128 VTAIL.n127 0.388379
R406 VTAIL.n94 VTAIL.n92 0.388379
R407 VTAIL VTAIL.n311 0.287138
R408 VTAIL.n260 VTAIL.n255 0.155672
R409 VTAIL.n267 VTAIL.n255 0.155672
R410 VTAIL.n268 VTAIL.n267 0.155672
R411 VTAIL.n268 VTAIL.n251 0.155672
R412 VTAIL.n275 VTAIL.n251 0.155672
R413 VTAIL.n276 VTAIL.n275 0.155672
R414 VTAIL.n276 VTAIL.n247 0.155672
R415 VTAIL.n285 VTAIL.n247 0.155672
R416 VTAIL.n286 VTAIL.n285 0.155672
R417 VTAIL.n286 VTAIL.n243 0.155672
R418 VTAIL.n293 VTAIL.n243 0.155672
R419 VTAIL.n294 VTAIL.n293 0.155672
R420 VTAIL.n294 VTAIL.n239 0.155672
R421 VTAIL.n301 VTAIL.n239 0.155672
R422 VTAIL.n302 VTAIL.n301 0.155672
R423 VTAIL.n302 VTAIL.n235 0.155672
R424 VTAIL.n309 VTAIL.n235 0.155672
R425 VTAIL.n26 VTAIL.n21 0.155672
R426 VTAIL.n33 VTAIL.n21 0.155672
R427 VTAIL.n34 VTAIL.n33 0.155672
R428 VTAIL.n34 VTAIL.n17 0.155672
R429 VTAIL.n41 VTAIL.n17 0.155672
R430 VTAIL.n42 VTAIL.n41 0.155672
R431 VTAIL.n42 VTAIL.n13 0.155672
R432 VTAIL.n51 VTAIL.n13 0.155672
R433 VTAIL.n52 VTAIL.n51 0.155672
R434 VTAIL.n52 VTAIL.n9 0.155672
R435 VTAIL.n59 VTAIL.n9 0.155672
R436 VTAIL.n60 VTAIL.n59 0.155672
R437 VTAIL.n60 VTAIL.n5 0.155672
R438 VTAIL.n67 VTAIL.n5 0.155672
R439 VTAIL.n68 VTAIL.n67 0.155672
R440 VTAIL.n68 VTAIL.n1 0.155672
R441 VTAIL.n75 VTAIL.n1 0.155672
R442 VTAIL.n231 VTAIL.n157 0.155672
R443 VTAIL.n224 VTAIL.n157 0.155672
R444 VTAIL.n224 VTAIL.n223 0.155672
R445 VTAIL.n223 VTAIL.n161 0.155672
R446 VTAIL.n216 VTAIL.n161 0.155672
R447 VTAIL.n216 VTAIL.n215 0.155672
R448 VTAIL.n215 VTAIL.n165 0.155672
R449 VTAIL.n208 VTAIL.n165 0.155672
R450 VTAIL.n208 VTAIL.n207 0.155672
R451 VTAIL.n207 VTAIL.n169 0.155672
R452 VTAIL.n199 VTAIL.n169 0.155672
R453 VTAIL.n199 VTAIL.n198 0.155672
R454 VTAIL.n198 VTAIL.n174 0.155672
R455 VTAIL.n191 VTAIL.n174 0.155672
R456 VTAIL.n191 VTAIL.n190 0.155672
R457 VTAIL.n190 VTAIL.n178 0.155672
R458 VTAIL.n183 VTAIL.n178 0.155672
R459 VTAIL.n153 VTAIL.n79 0.155672
R460 VTAIL.n146 VTAIL.n79 0.155672
R461 VTAIL.n146 VTAIL.n145 0.155672
R462 VTAIL.n145 VTAIL.n83 0.155672
R463 VTAIL.n138 VTAIL.n83 0.155672
R464 VTAIL.n138 VTAIL.n137 0.155672
R465 VTAIL.n137 VTAIL.n87 0.155672
R466 VTAIL.n130 VTAIL.n87 0.155672
R467 VTAIL.n130 VTAIL.n129 0.155672
R468 VTAIL.n129 VTAIL.n91 0.155672
R469 VTAIL.n121 VTAIL.n91 0.155672
R470 VTAIL.n121 VTAIL.n120 0.155672
R471 VTAIL.n120 VTAIL.n96 0.155672
R472 VTAIL.n113 VTAIL.n96 0.155672
R473 VTAIL.n113 VTAIL.n112 0.155672
R474 VTAIL.n112 VTAIL.n100 0.155672
R475 VTAIL.n105 VTAIL.n100 0.155672
R476 VDD1.n72 VDD1.n0 756.745
R477 VDD1.n149 VDD1.n77 756.745
R478 VDD1.n73 VDD1.n72 585
R479 VDD1.n71 VDD1.n70 585
R480 VDD1.n4 VDD1.n3 585
R481 VDD1.n65 VDD1.n64 585
R482 VDD1.n63 VDD1.n62 585
R483 VDD1.n8 VDD1.n7 585
R484 VDD1.n57 VDD1.n56 585
R485 VDD1.n55 VDD1.n54 585
R486 VDD1.n12 VDD1.n11 585
R487 VDD1.n49 VDD1.n48 585
R488 VDD1.n47 VDD1.n14 585
R489 VDD1.n46 VDD1.n45 585
R490 VDD1.n17 VDD1.n15 585
R491 VDD1.n40 VDD1.n39 585
R492 VDD1.n38 VDD1.n37 585
R493 VDD1.n21 VDD1.n20 585
R494 VDD1.n32 VDD1.n31 585
R495 VDD1.n30 VDD1.n29 585
R496 VDD1.n25 VDD1.n24 585
R497 VDD1.n101 VDD1.n100 585
R498 VDD1.n106 VDD1.n105 585
R499 VDD1.n108 VDD1.n107 585
R500 VDD1.n97 VDD1.n96 585
R501 VDD1.n114 VDD1.n113 585
R502 VDD1.n116 VDD1.n115 585
R503 VDD1.n93 VDD1.n92 585
R504 VDD1.n123 VDD1.n122 585
R505 VDD1.n124 VDD1.n91 585
R506 VDD1.n126 VDD1.n125 585
R507 VDD1.n89 VDD1.n88 585
R508 VDD1.n132 VDD1.n131 585
R509 VDD1.n134 VDD1.n133 585
R510 VDD1.n85 VDD1.n84 585
R511 VDD1.n140 VDD1.n139 585
R512 VDD1.n142 VDD1.n141 585
R513 VDD1.n81 VDD1.n80 585
R514 VDD1.n148 VDD1.n147 585
R515 VDD1.n150 VDD1.n149 585
R516 VDD1.n102 VDD1.t1 329.036
R517 VDD1.n26 VDD1.t0 329.036
R518 VDD1.n72 VDD1.n71 171.744
R519 VDD1.n71 VDD1.n3 171.744
R520 VDD1.n64 VDD1.n3 171.744
R521 VDD1.n64 VDD1.n63 171.744
R522 VDD1.n63 VDD1.n7 171.744
R523 VDD1.n56 VDD1.n7 171.744
R524 VDD1.n56 VDD1.n55 171.744
R525 VDD1.n55 VDD1.n11 171.744
R526 VDD1.n48 VDD1.n11 171.744
R527 VDD1.n48 VDD1.n47 171.744
R528 VDD1.n47 VDD1.n46 171.744
R529 VDD1.n46 VDD1.n15 171.744
R530 VDD1.n39 VDD1.n15 171.744
R531 VDD1.n39 VDD1.n38 171.744
R532 VDD1.n38 VDD1.n20 171.744
R533 VDD1.n31 VDD1.n20 171.744
R534 VDD1.n31 VDD1.n30 171.744
R535 VDD1.n30 VDD1.n24 171.744
R536 VDD1.n106 VDD1.n100 171.744
R537 VDD1.n107 VDD1.n106 171.744
R538 VDD1.n107 VDD1.n96 171.744
R539 VDD1.n114 VDD1.n96 171.744
R540 VDD1.n115 VDD1.n114 171.744
R541 VDD1.n115 VDD1.n92 171.744
R542 VDD1.n123 VDD1.n92 171.744
R543 VDD1.n124 VDD1.n123 171.744
R544 VDD1.n125 VDD1.n124 171.744
R545 VDD1.n125 VDD1.n88 171.744
R546 VDD1.n132 VDD1.n88 171.744
R547 VDD1.n133 VDD1.n132 171.744
R548 VDD1.n133 VDD1.n84 171.744
R549 VDD1.n140 VDD1.n84 171.744
R550 VDD1.n141 VDD1.n140 171.744
R551 VDD1.n141 VDD1.n80 171.744
R552 VDD1.n148 VDD1.n80 171.744
R553 VDD1.n149 VDD1.n148 171.744
R554 VDD1 VDD1.n153 88.4622
R555 VDD1.t0 VDD1.n24 85.8723
R556 VDD1.t1 VDD1.n100 85.8723
R557 VDD1 VDD1.n76 49.2672
R558 VDD1.n49 VDD1.n14 13.1884
R559 VDD1.n126 VDD1.n91 13.1884
R560 VDD1.n50 VDD1.n12 12.8005
R561 VDD1.n45 VDD1.n16 12.8005
R562 VDD1.n122 VDD1.n121 12.8005
R563 VDD1.n127 VDD1.n89 12.8005
R564 VDD1.n54 VDD1.n53 12.0247
R565 VDD1.n44 VDD1.n17 12.0247
R566 VDD1.n120 VDD1.n93 12.0247
R567 VDD1.n131 VDD1.n130 12.0247
R568 VDD1.n57 VDD1.n10 11.249
R569 VDD1.n41 VDD1.n40 11.249
R570 VDD1.n117 VDD1.n116 11.249
R571 VDD1.n134 VDD1.n87 11.249
R572 VDD1.n26 VDD1.n25 10.7239
R573 VDD1.n102 VDD1.n101 10.7239
R574 VDD1.n58 VDD1.n8 10.4732
R575 VDD1.n37 VDD1.n19 10.4732
R576 VDD1.n113 VDD1.n95 10.4732
R577 VDD1.n135 VDD1.n85 10.4732
R578 VDD1.n62 VDD1.n61 9.69747
R579 VDD1.n36 VDD1.n21 9.69747
R580 VDD1.n112 VDD1.n97 9.69747
R581 VDD1.n139 VDD1.n138 9.69747
R582 VDD1.n76 VDD1.n75 9.45567
R583 VDD1.n153 VDD1.n152 9.45567
R584 VDD1.n2 VDD1.n1 9.3005
R585 VDD1.n69 VDD1.n68 9.3005
R586 VDD1.n67 VDD1.n66 9.3005
R587 VDD1.n6 VDD1.n5 9.3005
R588 VDD1.n61 VDD1.n60 9.3005
R589 VDD1.n59 VDD1.n58 9.3005
R590 VDD1.n10 VDD1.n9 9.3005
R591 VDD1.n53 VDD1.n52 9.3005
R592 VDD1.n51 VDD1.n50 9.3005
R593 VDD1.n16 VDD1.n13 9.3005
R594 VDD1.n44 VDD1.n43 9.3005
R595 VDD1.n42 VDD1.n41 9.3005
R596 VDD1.n19 VDD1.n18 9.3005
R597 VDD1.n36 VDD1.n35 9.3005
R598 VDD1.n34 VDD1.n33 9.3005
R599 VDD1.n23 VDD1.n22 9.3005
R600 VDD1.n28 VDD1.n27 9.3005
R601 VDD1.n75 VDD1.n74 9.3005
R602 VDD1.n79 VDD1.n78 9.3005
R603 VDD1.n152 VDD1.n151 9.3005
R604 VDD1.n144 VDD1.n143 9.3005
R605 VDD1.n83 VDD1.n82 9.3005
R606 VDD1.n138 VDD1.n137 9.3005
R607 VDD1.n136 VDD1.n135 9.3005
R608 VDD1.n87 VDD1.n86 9.3005
R609 VDD1.n130 VDD1.n129 9.3005
R610 VDD1.n128 VDD1.n127 9.3005
R611 VDD1.n104 VDD1.n103 9.3005
R612 VDD1.n99 VDD1.n98 9.3005
R613 VDD1.n110 VDD1.n109 9.3005
R614 VDD1.n112 VDD1.n111 9.3005
R615 VDD1.n95 VDD1.n94 9.3005
R616 VDD1.n118 VDD1.n117 9.3005
R617 VDD1.n120 VDD1.n119 9.3005
R618 VDD1.n121 VDD1.n90 9.3005
R619 VDD1.n146 VDD1.n145 9.3005
R620 VDD1.n65 VDD1.n6 8.92171
R621 VDD1.n33 VDD1.n32 8.92171
R622 VDD1.n109 VDD1.n108 8.92171
R623 VDD1.n142 VDD1.n83 8.92171
R624 VDD1.n76 VDD1.n0 8.14595
R625 VDD1.n66 VDD1.n4 8.14595
R626 VDD1.n29 VDD1.n23 8.14595
R627 VDD1.n105 VDD1.n99 8.14595
R628 VDD1.n143 VDD1.n81 8.14595
R629 VDD1.n153 VDD1.n77 8.14595
R630 VDD1.n74 VDD1.n73 7.3702
R631 VDD1.n70 VDD1.n69 7.3702
R632 VDD1.n28 VDD1.n25 7.3702
R633 VDD1.n104 VDD1.n101 7.3702
R634 VDD1.n147 VDD1.n146 7.3702
R635 VDD1.n151 VDD1.n150 7.3702
R636 VDD1.n73 VDD1.n2 6.59444
R637 VDD1.n70 VDD1.n2 6.59444
R638 VDD1.n147 VDD1.n79 6.59444
R639 VDD1.n150 VDD1.n79 6.59444
R640 VDD1.n74 VDD1.n0 5.81868
R641 VDD1.n69 VDD1.n4 5.81868
R642 VDD1.n29 VDD1.n28 5.81868
R643 VDD1.n105 VDD1.n104 5.81868
R644 VDD1.n146 VDD1.n81 5.81868
R645 VDD1.n151 VDD1.n77 5.81868
R646 VDD1.n66 VDD1.n65 5.04292
R647 VDD1.n32 VDD1.n23 5.04292
R648 VDD1.n108 VDD1.n99 5.04292
R649 VDD1.n143 VDD1.n142 5.04292
R650 VDD1.n62 VDD1.n6 4.26717
R651 VDD1.n33 VDD1.n21 4.26717
R652 VDD1.n109 VDD1.n97 4.26717
R653 VDD1.n139 VDD1.n83 4.26717
R654 VDD1.n61 VDD1.n8 3.49141
R655 VDD1.n37 VDD1.n36 3.49141
R656 VDD1.n113 VDD1.n112 3.49141
R657 VDD1.n138 VDD1.n85 3.49141
R658 VDD1.n58 VDD1.n57 2.71565
R659 VDD1.n40 VDD1.n19 2.71565
R660 VDD1.n116 VDD1.n95 2.71565
R661 VDD1.n135 VDD1.n134 2.71565
R662 VDD1.n27 VDD1.n26 2.41282
R663 VDD1.n103 VDD1.n102 2.41282
R664 VDD1.n54 VDD1.n10 1.93989
R665 VDD1.n41 VDD1.n17 1.93989
R666 VDD1.n117 VDD1.n93 1.93989
R667 VDD1.n131 VDD1.n87 1.93989
R668 VDD1.n53 VDD1.n12 1.16414
R669 VDD1.n45 VDD1.n44 1.16414
R670 VDD1.n122 VDD1.n120 1.16414
R671 VDD1.n130 VDD1.n89 1.16414
R672 VDD1.n50 VDD1.n49 0.388379
R673 VDD1.n16 VDD1.n14 0.388379
R674 VDD1.n121 VDD1.n91 0.388379
R675 VDD1.n127 VDD1.n126 0.388379
R676 VDD1.n75 VDD1.n1 0.155672
R677 VDD1.n68 VDD1.n1 0.155672
R678 VDD1.n68 VDD1.n67 0.155672
R679 VDD1.n67 VDD1.n5 0.155672
R680 VDD1.n60 VDD1.n5 0.155672
R681 VDD1.n60 VDD1.n59 0.155672
R682 VDD1.n59 VDD1.n9 0.155672
R683 VDD1.n52 VDD1.n9 0.155672
R684 VDD1.n52 VDD1.n51 0.155672
R685 VDD1.n51 VDD1.n13 0.155672
R686 VDD1.n43 VDD1.n13 0.155672
R687 VDD1.n43 VDD1.n42 0.155672
R688 VDD1.n42 VDD1.n18 0.155672
R689 VDD1.n35 VDD1.n18 0.155672
R690 VDD1.n35 VDD1.n34 0.155672
R691 VDD1.n34 VDD1.n22 0.155672
R692 VDD1.n27 VDD1.n22 0.155672
R693 VDD1.n103 VDD1.n98 0.155672
R694 VDD1.n110 VDD1.n98 0.155672
R695 VDD1.n111 VDD1.n110 0.155672
R696 VDD1.n111 VDD1.n94 0.155672
R697 VDD1.n118 VDD1.n94 0.155672
R698 VDD1.n119 VDD1.n118 0.155672
R699 VDD1.n119 VDD1.n90 0.155672
R700 VDD1.n128 VDD1.n90 0.155672
R701 VDD1.n129 VDD1.n128 0.155672
R702 VDD1.n129 VDD1.n86 0.155672
R703 VDD1.n136 VDD1.n86 0.155672
R704 VDD1.n137 VDD1.n136 0.155672
R705 VDD1.n137 VDD1.n82 0.155672
R706 VDD1.n144 VDD1.n82 0.155672
R707 VDD1.n145 VDD1.n144 0.155672
R708 VDD1.n145 VDD1.n78 0.155672
R709 VDD1.n152 VDD1.n78 0.155672
R710 B.n336 B.n335 585
R711 B.n334 B.n87 585
R712 B.n333 B.n332 585
R713 B.n331 B.n88 585
R714 B.n330 B.n329 585
R715 B.n328 B.n89 585
R716 B.n327 B.n326 585
R717 B.n325 B.n90 585
R718 B.n324 B.n323 585
R719 B.n322 B.n91 585
R720 B.n321 B.n320 585
R721 B.n319 B.n92 585
R722 B.n318 B.n317 585
R723 B.n316 B.n93 585
R724 B.n315 B.n314 585
R725 B.n313 B.n94 585
R726 B.n312 B.n311 585
R727 B.n310 B.n95 585
R728 B.n309 B.n308 585
R729 B.n307 B.n96 585
R730 B.n306 B.n305 585
R731 B.n304 B.n97 585
R732 B.n303 B.n302 585
R733 B.n301 B.n98 585
R734 B.n300 B.n299 585
R735 B.n298 B.n99 585
R736 B.n297 B.n296 585
R737 B.n295 B.n100 585
R738 B.n294 B.n293 585
R739 B.n292 B.n101 585
R740 B.n291 B.n290 585
R741 B.n289 B.n102 585
R742 B.n288 B.n287 585
R743 B.n286 B.n103 585
R744 B.n285 B.n284 585
R745 B.n283 B.n104 585
R746 B.n282 B.n281 585
R747 B.n280 B.n105 585
R748 B.n279 B.n278 585
R749 B.n277 B.n106 585
R750 B.n276 B.n275 585
R751 B.n274 B.n107 585
R752 B.n273 B.n272 585
R753 B.n271 B.n108 585
R754 B.n270 B.n269 585
R755 B.n268 B.n109 585
R756 B.n267 B.n266 585
R757 B.n265 B.n110 585
R758 B.n263 B.n262 585
R759 B.n261 B.n113 585
R760 B.n260 B.n259 585
R761 B.n258 B.n114 585
R762 B.n257 B.n256 585
R763 B.n255 B.n115 585
R764 B.n254 B.n253 585
R765 B.n252 B.n116 585
R766 B.n251 B.n250 585
R767 B.n249 B.n117 585
R768 B.n248 B.n247 585
R769 B.n243 B.n118 585
R770 B.n242 B.n241 585
R771 B.n240 B.n119 585
R772 B.n239 B.n238 585
R773 B.n237 B.n120 585
R774 B.n236 B.n235 585
R775 B.n234 B.n121 585
R776 B.n233 B.n232 585
R777 B.n231 B.n122 585
R778 B.n230 B.n229 585
R779 B.n228 B.n123 585
R780 B.n227 B.n226 585
R781 B.n225 B.n124 585
R782 B.n224 B.n223 585
R783 B.n222 B.n125 585
R784 B.n221 B.n220 585
R785 B.n219 B.n126 585
R786 B.n218 B.n217 585
R787 B.n216 B.n127 585
R788 B.n215 B.n214 585
R789 B.n213 B.n128 585
R790 B.n212 B.n211 585
R791 B.n210 B.n129 585
R792 B.n209 B.n208 585
R793 B.n207 B.n130 585
R794 B.n206 B.n205 585
R795 B.n204 B.n131 585
R796 B.n203 B.n202 585
R797 B.n201 B.n132 585
R798 B.n200 B.n199 585
R799 B.n198 B.n133 585
R800 B.n197 B.n196 585
R801 B.n195 B.n134 585
R802 B.n194 B.n193 585
R803 B.n192 B.n135 585
R804 B.n191 B.n190 585
R805 B.n189 B.n136 585
R806 B.n188 B.n187 585
R807 B.n186 B.n137 585
R808 B.n185 B.n184 585
R809 B.n183 B.n138 585
R810 B.n182 B.n181 585
R811 B.n180 B.n139 585
R812 B.n179 B.n178 585
R813 B.n177 B.n140 585
R814 B.n176 B.n175 585
R815 B.n174 B.n141 585
R816 B.n337 B.n86 585
R817 B.n339 B.n338 585
R818 B.n340 B.n85 585
R819 B.n342 B.n341 585
R820 B.n343 B.n84 585
R821 B.n345 B.n344 585
R822 B.n346 B.n83 585
R823 B.n348 B.n347 585
R824 B.n349 B.n82 585
R825 B.n351 B.n350 585
R826 B.n352 B.n81 585
R827 B.n354 B.n353 585
R828 B.n355 B.n80 585
R829 B.n357 B.n356 585
R830 B.n358 B.n79 585
R831 B.n360 B.n359 585
R832 B.n361 B.n78 585
R833 B.n363 B.n362 585
R834 B.n364 B.n77 585
R835 B.n366 B.n365 585
R836 B.n367 B.n76 585
R837 B.n369 B.n368 585
R838 B.n370 B.n75 585
R839 B.n372 B.n371 585
R840 B.n373 B.n74 585
R841 B.n375 B.n374 585
R842 B.n376 B.n73 585
R843 B.n378 B.n377 585
R844 B.n379 B.n72 585
R845 B.n381 B.n380 585
R846 B.n382 B.n71 585
R847 B.n384 B.n383 585
R848 B.n385 B.n70 585
R849 B.n387 B.n386 585
R850 B.n388 B.n69 585
R851 B.n390 B.n389 585
R852 B.n550 B.n549 585
R853 B.n548 B.n11 585
R854 B.n547 B.n546 585
R855 B.n545 B.n12 585
R856 B.n544 B.n543 585
R857 B.n542 B.n13 585
R858 B.n541 B.n540 585
R859 B.n539 B.n14 585
R860 B.n538 B.n537 585
R861 B.n536 B.n15 585
R862 B.n535 B.n534 585
R863 B.n533 B.n16 585
R864 B.n532 B.n531 585
R865 B.n530 B.n17 585
R866 B.n529 B.n528 585
R867 B.n527 B.n18 585
R868 B.n526 B.n525 585
R869 B.n524 B.n19 585
R870 B.n523 B.n522 585
R871 B.n521 B.n20 585
R872 B.n520 B.n519 585
R873 B.n518 B.n21 585
R874 B.n517 B.n516 585
R875 B.n515 B.n22 585
R876 B.n514 B.n513 585
R877 B.n512 B.n23 585
R878 B.n511 B.n510 585
R879 B.n509 B.n24 585
R880 B.n508 B.n507 585
R881 B.n506 B.n25 585
R882 B.n505 B.n504 585
R883 B.n503 B.n26 585
R884 B.n502 B.n501 585
R885 B.n500 B.n27 585
R886 B.n499 B.n498 585
R887 B.n497 B.n28 585
R888 B.n496 B.n495 585
R889 B.n494 B.n29 585
R890 B.n493 B.n492 585
R891 B.n491 B.n30 585
R892 B.n490 B.n489 585
R893 B.n488 B.n31 585
R894 B.n487 B.n486 585
R895 B.n485 B.n32 585
R896 B.n484 B.n483 585
R897 B.n482 B.n33 585
R898 B.n481 B.n480 585
R899 B.n479 B.n34 585
R900 B.n478 B.n477 585
R901 B.n476 B.n35 585
R902 B.n475 B.n474 585
R903 B.n473 B.n39 585
R904 B.n472 B.n471 585
R905 B.n470 B.n40 585
R906 B.n469 B.n468 585
R907 B.n467 B.n41 585
R908 B.n466 B.n465 585
R909 B.n464 B.n42 585
R910 B.n462 B.n461 585
R911 B.n460 B.n45 585
R912 B.n459 B.n458 585
R913 B.n457 B.n46 585
R914 B.n456 B.n455 585
R915 B.n454 B.n47 585
R916 B.n453 B.n452 585
R917 B.n451 B.n48 585
R918 B.n450 B.n449 585
R919 B.n448 B.n49 585
R920 B.n447 B.n446 585
R921 B.n445 B.n50 585
R922 B.n444 B.n443 585
R923 B.n442 B.n51 585
R924 B.n441 B.n440 585
R925 B.n439 B.n52 585
R926 B.n438 B.n437 585
R927 B.n436 B.n53 585
R928 B.n435 B.n434 585
R929 B.n433 B.n54 585
R930 B.n432 B.n431 585
R931 B.n430 B.n55 585
R932 B.n429 B.n428 585
R933 B.n427 B.n56 585
R934 B.n426 B.n425 585
R935 B.n424 B.n57 585
R936 B.n423 B.n422 585
R937 B.n421 B.n58 585
R938 B.n420 B.n419 585
R939 B.n418 B.n59 585
R940 B.n417 B.n416 585
R941 B.n415 B.n60 585
R942 B.n414 B.n413 585
R943 B.n412 B.n61 585
R944 B.n411 B.n410 585
R945 B.n409 B.n62 585
R946 B.n408 B.n407 585
R947 B.n406 B.n63 585
R948 B.n405 B.n404 585
R949 B.n403 B.n64 585
R950 B.n402 B.n401 585
R951 B.n400 B.n65 585
R952 B.n399 B.n398 585
R953 B.n397 B.n66 585
R954 B.n396 B.n395 585
R955 B.n394 B.n67 585
R956 B.n393 B.n392 585
R957 B.n391 B.n68 585
R958 B.n551 B.n10 585
R959 B.n553 B.n552 585
R960 B.n554 B.n9 585
R961 B.n556 B.n555 585
R962 B.n557 B.n8 585
R963 B.n559 B.n558 585
R964 B.n560 B.n7 585
R965 B.n562 B.n561 585
R966 B.n563 B.n6 585
R967 B.n565 B.n564 585
R968 B.n566 B.n5 585
R969 B.n568 B.n567 585
R970 B.n569 B.n4 585
R971 B.n571 B.n570 585
R972 B.n572 B.n3 585
R973 B.n574 B.n573 585
R974 B.n575 B.n0 585
R975 B.n2 B.n1 585
R976 B.n150 B.n149 585
R977 B.n152 B.n151 585
R978 B.n153 B.n148 585
R979 B.n155 B.n154 585
R980 B.n156 B.n147 585
R981 B.n158 B.n157 585
R982 B.n159 B.n146 585
R983 B.n161 B.n160 585
R984 B.n162 B.n145 585
R985 B.n164 B.n163 585
R986 B.n165 B.n144 585
R987 B.n167 B.n166 585
R988 B.n168 B.n143 585
R989 B.n170 B.n169 585
R990 B.n171 B.n142 585
R991 B.n173 B.n172 585
R992 B.n174 B.n173 521.33
R993 B.n335 B.n86 521.33
R994 B.n389 B.n68 521.33
R995 B.n551 B.n550 521.33
R996 B.n244 B.t3 475.45
R997 B.n111 B.t6 475.45
R998 B.n43 B.t9 475.45
R999 B.n36 B.t0 475.45
R1000 B.n111 B.t7 447.957
R1001 B.n43 B.t11 447.957
R1002 B.n244 B.t4 447.957
R1003 B.n36 B.t2 447.957
R1004 B.n112 B.t8 416.926
R1005 B.n44 B.t10 416.926
R1006 B.n245 B.t5 416.926
R1007 B.n37 B.t1 416.926
R1008 B.n577 B.n576 256.663
R1009 B.n576 B.n575 235.042
R1010 B.n576 B.n2 235.042
R1011 B.n175 B.n174 163.367
R1012 B.n175 B.n140 163.367
R1013 B.n179 B.n140 163.367
R1014 B.n180 B.n179 163.367
R1015 B.n181 B.n180 163.367
R1016 B.n181 B.n138 163.367
R1017 B.n185 B.n138 163.367
R1018 B.n186 B.n185 163.367
R1019 B.n187 B.n186 163.367
R1020 B.n187 B.n136 163.367
R1021 B.n191 B.n136 163.367
R1022 B.n192 B.n191 163.367
R1023 B.n193 B.n192 163.367
R1024 B.n193 B.n134 163.367
R1025 B.n197 B.n134 163.367
R1026 B.n198 B.n197 163.367
R1027 B.n199 B.n198 163.367
R1028 B.n199 B.n132 163.367
R1029 B.n203 B.n132 163.367
R1030 B.n204 B.n203 163.367
R1031 B.n205 B.n204 163.367
R1032 B.n205 B.n130 163.367
R1033 B.n209 B.n130 163.367
R1034 B.n210 B.n209 163.367
R1035 B.n211 B.n210 163.367
R1036 B.n211 B.n128 163.367
R1037 B.n215 B.n128 163.367
R1038 B.n216 B.n215 163.367
R1039 B.n217 B.n216 163.367
R1040 B.n217 B.n126 163.367
R1041 B.n221 B.n126 163.367
R1042 B.n222 B.n221 163.367
R1043 B.n223 B.n222 163.367
R1044 B.n223 B.n124 163.367
R1045 B.n227 B.n124 163.367
R1046 B.n228 B.n227 163.367
R1047 B.n229 B.n228 163.367
R1048 B.n229 B.n122 163.367
R1049 B.n233 B.n122 163.367
R1050 B.n234 B.n233 163.367
R1051 B.n235 B.n234 163.367
R1052 B.n235 B.n120 163.367
R1053 B.n239 B.n120 163.367
R1054 B.n240 B.n239 163.367
R1055 B.n241 B.n240 163.367
R1056 B.n241 B.n118 163.367
R1057 B.n248 B.n118 163.367
R1058 B.n249 B.n248 163.367
R1059 B.n250 B.n249 163.367
R1060 B.n250 B.n116 163.367
R1061 B.n254 B.n116 163.367
R1062 B.n255 B.n254 163.367
R1063 B.n256 B.n255 163.367
R1064 B.n256 B.n114 163.367
R1065 B.n260 B.n114 163.367
R1066 B.n261 B.n260 163.367
R1067 B.n262 B.n261 163.367
R1068 B.n262 B.n110 163.367
R1069 B.n267 B.n110 163.367
R1070 B.n268 B.n267 163.367
R1071 B.n269 B.n268 163.367
R1072 B.n269 B.n108 163.367
R1073 B.n273 B.n108 163.367
R1074 B.n274 B.n273 163.367
R1075 B.n275 B.n274 163.367
R1076 B.n275 B.n106 163.367
R1077 B.n279 B.n106 163.367
R1078 B.n280 B.n279 163.367
R1079 B.n281 B.n280 163.367
R1080 B.n281 B.n104 163.367
R1081 B.n285 B.n104 163.367
R1082 B.n286 B.n285 163.367
R1083 B.n287 B.n286 163.367
R1084 B.n287 B.n102 163.367
R1085 B.n291 B.n102 163.367
R1086 B.n292 B.n291 163.367
R1087 B.n293 B.n292 163.367
R1088 B.n293 B.n100 163.367
R1089 B.n297 B.n100 163.367
R1090 B.n298 B.n297 163.367
R1091 B.n299 B.n298 163.367
R1092 B.n299 B.n98 163.367
R1093 B.n303 B.n98 163.367
R1094 B.n304 B.n303 163.367
R1095 B.n305 B.n304 163.367
R1096 B.n305 B.n96 163.367
R1097 B.n309 B.n96 163.367
R1098 B.n310 B.n309 163.367
R1099 B.n311 B.n310 163.367
R1100 B.n311 B.n94 163.367
R1101 B.n315 B.n94 163.367
R1102 B.n316 B.n315 163.367
R1103 B.n317 B.n316 163.367
R1104 B.n317 B.n92 163.367
R1105 B.n321 B.n92 163.367
R1106 B.n322 B.n321 163.367
R1107 B.n323 B.n322 163.367
R1108 B.n323 B.n90 163.367
R1109 B.n327 B.n90 163.367
R1110 B.n328 B.n327 163.367
R1111 B.n329 B.n328 163.367
R1112 B.n329 B.n88 163.367
R1113 B.n333 B.n88 163.367
R1114 B.n334 B.n333 163.367
R1115 B.n335 B.n334 163.367
R1116 B.n389 B.n388 163.367
R1117 B.n388 B.n387 163.367
R1118 B.n387 B.n70 163.367
R1119 B.n383 B.n70 163.367
R1120 B.n383 B.n382 163.367
R1121 B.n382 B.n381 163.367
R1122 B.n381 B.n72 163.367
R1123 B.n377 B.n72 163.367
R1124 B.n377 B.n376 163.367
R1125 B.n376 B.n375 163.367
R1126 B.n375 B.n74 163.367
R1127 B.n371 B.n74 163.367
R1128 B.n371 B.n370 163.367
R1129 B.n370 B.n369 163.367
R1130 B.n369 B.n76 163.367
R1131 B.n365 B.n76 163.367
R1132 B.n365 B.n364 163.367
R1133 B.n364 B.n363 163.367
R1134 B.n363 B.n78 163.367
R1135 B.n359 B.n78 163.367
R1136 B.n359 B.n358 163.367
R1137 B.n358 B.n357 163.367
R1138 B.n357 B.n80 163.367
R1139 B.n353 B.n80 163.367
R1140 B.n353 B.n352 163.367
R1141 B.n352 B.n351 163.367
R1142 B.n351 B.n82 163.367
R1143 B.n347 B.n82 163.367
R1144 B.n347 B.n346 163.367
R1145 B.n346 B.n345 163.367
R1146 B.n345 B.n84 163.367
R1147 B.n341 B.n84 163.367
R1148 B.n341 B.n340 163.367
R1149 B.n340 B.n339 163.367
R1150 B.n339 B.n86 163.367
R1151 B.n550 B.n11 163.367
R1152 B.n546 B.n11 163.367
R1153 B.n546 B.n545 163.367
R1154 B.n545 B.n544 163.367
R1155 B.n544 B.n13 163.367
R1156 B.n540 B.n13 163.367
R1157 B.n540 B.n539 163.367
R1158 B.n539 B.n538 163.367
R1159 B.n538 B.n15 163.367
R1160 B.n534 B.n15 163.367
R1161 B.n534 B.n533 163.367
R1162 B.n533 B.n532 163.367
R1163 B.n532 B.n17 163.367
R1164 B.n528 B.n17 163.367
R1165 B.n528 B.n527 163.367
R1166 B.n527 B.n526 163.367
R1167 B.n526 B.n19 163.367
R1168 B.n522 B.n19 163.367
R1169 B.n522 B.n521 163.367
R1170 B.n521 B.n520 163.367
R1171 B.n520 B.n21 163.367
R1172 B.n516 B.n21 163.367
R1173 B.n516 B.n515 163.367
R1174 B.n515 B.n514 163.367
R1175 B.n514 B.n23 163.367
R1176 B.n510 B.n23 163.367
R1177 B.n510 B.n509 163.367
R1178 B.n509 B.n508 163.367
R1179 B.n508 B.n25 163.367
R1180 B.n504 B.n25 163.367
R1181 B.n504 B.n503 163.367
R1182 B.n503 B.n502 163.367
R1183 B.n502 B.n27 163.367
R1184 B.n498 B.n27 163.367
R1185 B.n498 B.n497 163.367
R1186 B.n497 B.n496 163.367
R1187 B.n496 B.n29 163.367
R1188 B.n492 B.n29 163.367
R1189 B.n492 B.n491 163.367
R1190 B.n491 B.n490 163.367
R1191 B.n490 B.n31 163.367
R1192 B.n486 B.n31 163.367
R1193 B.n486 B.n485 163.367
R1194 B.n485 B.n484 163.367
R1195 B.n484 B.n33 163.367
R1196 B.n480 B.n33 163.367
R1197 B.n480 B.n479 163.367
R1198 B.n479 B.n478 163.367
R1199 B.n478 B.n35 163.367
R1200 B.n474 B.n35 163.367
R1201 B.n474 B.n473 163.367
R1202 B.n473 B.n472 163.367
R1203 B.n472 B.n40 163.367
R1204 B.n468 B.n40 163.367
R1205 B.n468 B.n467 163.367
R1206 B.n467 B.n466 163.367
R1207 B.n466 B.n42 163.367
R1208 B.n461 B.n42 163.367
R1209 B.n461 B.n460 163.367
R1210 B.n460 B.n459 163.367
R1211 B.n459 B.n46 163.367
R1212 B.n455 B.n46 163.367
R1213 B.n455 B.n454 163.367
R1214 B.n454 B.n453 163.367
R1215 B.n453 B.n48 163.367
R1216 B.n449 B.n48 163.367
R1217 B.n449 B.n448 163.367
R1218 B.n448 B.n447 163.367
R1219 B.n447 B.n50 163.367
R1220 B.n443 B.n50 163.367
R1221 B.n443 B.n442 163.367
R1222 B.n442 B.n441 163.367
R1223 B.n441 B.n52 163.367
R1224 B.n437 B.n52 163.367
R1225 B.n437 B.n436 163.367
R1226 B.n436 B.n435 163.367
R1227 B.n435 B.n54 163.367
R1228 B.n431 B.n54 163.367
R1229 B.n431 B.n430 163.367
R1230 B.n430 B.n429 163.367
R1231 B.n429 B.n56 163.367
R1232 B.n425 B.n56 163.367
R1233 B.n425 B.n424 163.367
R1234 B.n424 B.n423 163.367
R1235 B.n423 B.n58 163.367
R1236 B.n419 B.n58 163.367
R1237 B.n419 B.n418 163.367
R1238 B.n418 B.n417 163.367
R1239 B.n417 B.n60 163.367
R1240 B.n413 B.n60 163.367
R1241 B.n413 B.n412 163.367
R1242 B.n412 B.n411 163.367
R1243 B.n411 B.n62 163.367
R1244 B.n407 B.n62 163.367
R1245 B.n407 B.n406 163.367
R1246 B.n406 B.n405 163.367
R1247 B.n405 B.n64 163.367
R1248 B.n401 B.n64 163.367
R1249 B.n401 B.n400 163.367
R1250 B.n400 B.n399 163.367
R1251 B.n399 B.n66 163.367
R1252 B.n395 B.n66 163.367
R1253 B.n395 B.n394 163.367
R1254 B.n394 B.n393 163.367
R1255 B.n393 B.n68 163.367
R1256 B.n552 B.n551 163.367
R1257 B.n552 B.n9 163.367
R1258 B.n556 B.n9 163.367
R1259 B.n557 B.n556 163.367
R1260 B.n558 B.n557 163.367
R1261 B.n558 B.n7 163.367
R1262 B.n562 B.n7 163.367
R1263 B.n563 B.n562 163.367
R1264 B.n564 B.n563 163.367
R1265 B.n564 B.n5 163.367
R1266 B.n568 B.n5 163.367
R1267 B.n569 B.n568 163.367
R1268 B.n570 B.n569 163.367
R1269 B.n570 B.n3 163.367
R1270 B.n574 B.n3 163.367
R1271 B.n575 B.n574 163.367
R1272 B.n150 B.n2 163.367
R1273 B.n151 B.n150 163.367
R1274 B.n151 B.n148 163.367
R1275 B.n155 B.n148 163.367
R1276 B.n156 B.n155 163.367
R1277 B.n157 B.n156 163.367
R1278 B.n157 B.n146 163.367
R1279 B.n161 B.n146 163.367
R1280 B.n162 B.n161 163.367
R1281 B.n163 B.n162 163.367
R1282 B.n163 B.n144 163.367
R1283 B.n167 B.n144 163.367
R1284 B.n168 B.n167 163.367
R1285 B.n169 B.n168 163.367
R1286 B.n169 B.n142 163.367
R1287 B.n173 B.n142 163.367
R1288 B.n246 B.n245 59.5399
R1289 B.n264 B.n112 59.5399
R1290 B.n463 B.n44 59.5399
R1291 B.n38 B.n37 59.5399
R1292 B.n549 B.n10 33.8737
R1293 B.n391 B.n390 33.8737
R1294 B.n337 B.n336 33.8737
R1295 B.n172 B.n141 33.8737
R1296 B.n245 B.n244 31.0308
R1297 B.n112 B.n111 31.0308
R1298 B.n44 B.n43 31.0308
R1299 B.n37 B.n36 31.0308
R1300 B B.n577 18.0485
R1301 B.n553 B.n10 10.6151
R1302 B.n554 B.n553 10.6151
R1303 B.n555 B.n554 10.6151
R1304 B.n555 B.n8 10.6151
R1305 B.n559 B.n8 10.6151
R1306 B.n560 B.n559 10.6151
R1307 B.n561 B.n560 10.6151
R1308 B.n561 B.n6 10.6151
R1309 B.n565 B.n6 10.6151
R1310 B.n566 B.n565 10.6151
R1311 B.n567 B.n566 10.6151
R1312 B.n567 B.n4 10.6151
R1313 B.n571 B.n4 10.6151
R1314 B.n572 B.n571 10.6151
R1315 B.n573 B.n572 10.6151
R1316 B.n573 B.n0 10.6151
R1317 B.n549 B.n548 10.6151
R1318 B.n548 B.n547 10.6151
R1319 B.n547 B.n12 10.6151
R1320 B.n543 B.n12 10.6151
R1321 B.n543 B.n542 10.6151
R1322 B.n542 B.n541 10.6151
R1323 B.n541 B.n14 10.6151
R1324 B.n537 B.n14 10.6151
R1325 B.n537 B.n536 10.6151
R1326 B.n536 B.n535 10.6151
R1327 B.n535 B.n16 10.6151
R1328 B.n531 B.n16 10.6151
R1329 B.n531 B.n530 10.6151
R1330 B.n530 B.n529 10.6151
R1331 B.n529 B.n18 10.6151
R1332 B.n525 B.n18 10.6151
R1333 B.n525 B.n524 10.6151
R1334 B.n524 B.n523 10.6151
R1335 B.n523 B.n20 10.6151
R1336 B.n519 B.n20 10.6151
R1337 B.n519 B.n518 10.6151
R1338 B.n518 B.n517 10.6151
R1339 B.n517 B.n22 10.6151
R1340 B.n513 B.n22 10.6151
R1341 B.n513 B.n512 10.6151
R1342 B.n512 B.n511 10.6151
R1343 B.n511 B.n24 10.6151
R1344 B.n507 B.n24 10.6151
R1345 B.n507 B.n506 10.6151
R1346 B.n506 B.n505 10.6151
R1347 B.n505 B.n26 10.6151
R1348 B.n501 B.n26 10.6151
R1349 B.n501 B.n500 10.6151
R1350 B.n500 B.n499 10.6151
R1351 B.n499 B.n28 10.6151
R1352 B.n495 B.n28 10.6151
R1353 B.n495 B.n494 10.6151
R1354 B.n494 B.n493 10.6151
R1355 B.n493 B.n30 10.6151
R1356 B.n489 B.n30 10.6151
R1357 B.n489 B.n488 10.6151
R1358 B.n488 B.n487 10.6151
R1359 B.n487 B.n32 10.6151
R1360 B.n483 B.n32 10.6151
R1361 B.n483 B.n482 10.6151
R1362 B.n482 B.n481 10.6151
R1363 B.n481 B.n34 10.6151
R1364 B.n477 B.n476 10.6151
R1365 B.n476 B.n475 10.6151
R1366 B.n475 B.n39 10.6151
R1367 B.n471 B.n39 10.6151
R1368 B.n471 B.n470 10.6151
R1369 B.n470 B.n469 10.6151
R1370 B.n469 B.n41 10.6151
R1371 B.n465 B.n41 10.6151
R1372 B.n465 B.n464 10.6151
R1373 B.n462 B.n45 10.6151
R1374 B.n458 B.n45 10.6151
R1375 B.n458 B.n457 10.6151
R1376 B.n457 B.n456 10.6151
R1377 B.n456 B.n47 10.6151
R1378 B.n452 B.n47 10.6151
R1379 B.n452 B.n451 10.6151
R1380 B.n451 B.n450 10.6151
R1381 B.n450 B.n49 10.6151
R1382 B.n446 B.n49 10.6151
R1383 B.n446 B.n445 10.6151
R1384 B.n445 B.n444 10.6151
R1385 B.n444 B.n51 10.6151
R1386 B.n440 B.n51 10.6151
R1387 B.n440 B.n439 10.6151
R1388 B.n439 B.n438 10.6151
R1389 B.n438 B.n53 10.6151
R1390 B.n434 B.n53 10.6151
R1391 B.n434 B.n433 10.6151
R1392 B.n433 B.n432 10.6151
R1393 B.n432 B.n55 10.6151
R1394 B.n428 B.n55 10.6151
R1395 B.n428 B.n427 10.6151
R1396 B.n427 B.n426 10.6151
R1397 B.n426 B.n57 10.6151
R1398 B.n422 B.n57 10.6151
R1399 B.n422 B.n421 10.6151
R1400 B.n421 B.n420 10.6151
R1401 B.n420 B.n59 10.6151
R1402 B.n416 B.n59 10.6151
R1403 B.n416 B.n415 10.6151
R1404 B.n415 B.n414 10.6151
R1405 B.n414 B.n61 10.6151
R1406 B.n410 B.n61 10.6151
R1407 B.n410 B.n409 10.6151
R1408 B.n409 B.n408 10.6151
R1409 B.n408 B.n63 10.6151
R1410 B.n404 B.n63 10.6151
R1411 B.n404 B.n403 10.6151
R1412 B.n403 B.n402 10.6151
R1413 B.n402 B.n65 10.6151
R1414 B.n398 B.n65 10.6151
R1415 B.n398 B.n397 10.6151
R1416 B.n397 B.n396 10.6151
R1417 B.n396 B.n67 10.6151
R1418 B.n392 B.n67 10.6151
R1419 B.n392 B.n391 10.6151
R1420 B.n390 B.n69 10.6151
R1421 B.n386 B.n69 10.6151
R1422 B.n386 B.n385 10.6151
R1423 B.n385 B.n384 10.6151
R1424 B.n384 B.n71 10.6151
R1425 B.n380 B.n71 10.6151
R1426 B.n380 B.n379 10.6151
R1427 B.n379 B.n378 10.6151
R1428 B.n378 B.n73 10.6151
R1429 B.n374 B.n73 10.6151
R1430 B.n374 B.n373 10.6151
R1431 B.n373 B.n372 10.6151
R1432 B.n372 B.n75 10.6151
R1433 B.n368 B.n75 10.6151
R1434 B.n368 B.n367 10.6151
R1435 B.n367 B.n366 10.6151
R1436 B.n366 B.n77 10.6151
R1437 B.n362 B.n77 10.6151
R1438 B.n362 B.n361 10.6151
R1439 B.n361 B.n360 10.6151
R1440 B.n360 B.n79 10.6151
R1441 B.n356 B.n79 10.6151
R1442 B.n356 B.n355 10.6151
R1443 B.n355 B.n354 10.6151
R1444 B.n354 B.n81 10.6151
R1445 B.n350 B.n81 10.6151
R1446 B.n350 B.n349 10.6151
R1447 B.n349 B.n348 10.6151
R1448 B.n348 B.n83 10.6151
R1449 B.n344 B.n83 10.6151
R1450 B.n344 B.n343 10.6151
R1451 B.n343 B.n342 10.6151
R1452 B.n342 B.n85 10.6151
R1453 B.n338 B.n85 10.6151
R1454 B.n338 B.n337 10.6151
R1455 B.n149 B.n1 10.6151
R1456 B.n152 B.n149 10.6151
R1457 B.n153 B.n152 10.6151
R1458 B.n154 B.n153 10.6151
R1459 B.n154 B.n147 10.6151
R1460 B.n158 B.n147 10.6151
R1461 B.n159 B.n158 10.6151
R1462 B.n160 B.n159 10.6151
R1463 B.n160 B.n145 10.6151
R1464 B.n164 B.n145 10.6151
R1465 B.n165 B.n164 10.6151
R1466 B.n166 B.n165 10.6151
R1467 B.n166 B.n143 10.6151
R1468 B.n170 B.n143 10.6151
R1469 B.n171 B.n170 10.6151
R1470 B.n172 B.n171 10.6151
R1471 B.n176 B.n141 10.6151
R1472 B.n177 B.n176 10.6151
R1473 B.n178 B.n177 10.6151
R1474 B.n178 B.n139 10.6151
R1475 B.n182 B.n139 10.6151
R1476 B.n183 B.n182 10.6151
R1477 B.n184 B.n183 10.6151
R1478 B.n184 B.n137 10.6151
R1479 B.n188 B.n137 10.6151
R1480 B.n189 B.n188 10.6151
R1481 B.n190 B.n189 10.6151
R1482 B.n190 B.n135 10.6151
R1483 B.n194 B.n135 10.6151
R1484 B.n195 B.n194 10.6151
R1485 B.n196 B.n195 10.6151
R1486 B.n196 B.n133 10.6151
R1487 B.n200 B.n133 10.6151
R1488 B.n201 B.n200 10.6151
R1489 B.n202 B.n201 10.6151
R1490 B.n202 B.n131 10.6151
R1491 B.n206 B.n131 10.6151
R1492 B.n207 B.n206 10.6151
R1493 B.n208 B.n207 10.6151
R1494 B.n208 B.n129 10.6151
R1495 B.n212 B.n129 10.6151
R1496 B.n213 B.n212 10.6151
R1497 B.n214 B.n213 10.6151
R1498 B.n214 B.n127 10.6151
R1499 B.n218 B.n127 10.6151
R1500 B.n219 B.n218 10.6151
R1501 B.n220 B.n219 10.6151
R1502 B.n220 B.n125 10.6151
R1503 B.n224 B.n125 10.6151
R1504 B.n225 B.n224 10.6151
R1505 B.n226 B.n225 10.6151
R1506 B.n226 B.n123 10.6151
R1507 B.n230 B.n123 10.6151
R1508 B.n231 B.n230 10.6151
R1509 B.n232 B.n231 10.6151
R1510 B.n232 B.n121 10.6151
R1511 B.n236 B.n121 10.6151
R1512 B.n237 B.n236 10.6151
R1513 B.n238 B.n237 10.6151
R1514 B.n238 B.n119 10.6151
R1515 B.n242 B.n119 10.6151
R1516 B.n243 B.n242 10.6151
R1517 B.n247 B.n243 10.6151
R1518 B.n251 B.n117 10.6151
R1519 B.n252 B.n251 10.6151
R1520 B.n253 B.n252 10.6151
R1521 B.n253 B.n115 10.6151
R1522 B.n257 B.n115 10.6151
R1523 B.n258 B.n257 10.6151
R1524 B.n259 B.n258 10.6151
R1525 B.n259 B.n113 10.6151
R1526 B.n263 B.n113 10.6151
R1527 B.n266 B.n265 10.6151
R1528 B.n266 B.n109 10.6151
R1529 B.n270 B.n109 10.6151
R1530 B.n271 B.n270 10.6151
R1531 B.n272 B.n271 10.6151
R1532 B.n272 B.n107 10.6151
R1533 B.n276 B.n107 10.6151
R1534 B.n277 B.n276 10.6151
R1535 B.n278 B.n277 10.6151
R1536 B.n278 B.n105 10.6151
R1537 B.n282 B.n105 10.6151
R1538 B.n283 B.n282 10.6151
R1539 B.n284 B.n283 10.6151
R1540 B.n284 B.n103 10.6151
R1541 B.n288 B.n103 10.6151
R1542 B.n289 B.n288 10.6151
R1543 B.n290 B.n289 10.6151
R1544 B.n290 B.n101 10.6151
R1545 B.n294 B.n101 10.6151
R1546 B.n295 B.n294 10.6151
R1547 B.n296 B.n295 10.6151
R1548 B.n296 B.n99 10.6151
R1549 B.n300 B.n99 10.6151
R1550 B.n301 B.n300 10.6151
R1551 B.n302 B.n301 10.6151
R1552 B.n302 B.n97 10.6151
R1553 B.n306 B.n97 10.6151
R1554 B.n307 B.n306 10.6151
R1555 B.n308 B.n307 10.6151
R1556 B.n308 B.n95 10.6151
R1557 B.n312 B.n95 10.6151
R1558 B.n313 B.n312 10.6151
R1559 B.n314 B.n313 10.6151
R1560 B.n314 B.n93 10.6151
R1561 B.n318 B.n93 10.6151
R1562 B.n319 B.n318 10.6151
R1563 B.n320 B.n319 10.6151
R1564 B.n320 B.n91 10.6151
R1565 B.n324 B.n91 10.6151
R1566 B.n325 B.n324 10.6151
R1567 B.n326 B.n325 10.6151
R1568 B.n326 B.n89 10.6151
R1569 B.n330 B.n89 10.6151
R1570 B.n331 B.n330 10.6151
R1571 B.n332 B.n331 10.6151
R1572 B.n332 B.n87 10.6151
R1573 B.n336 B.n87 10.6151
R1574 B.n38 B.n34 9.36635
R1575 B.n463 B.n462 9.36635
R1576 B.n247 B.n246 9.36635
R1577 B.n265 B.n264 9.36635
R1578 B.n577 B.n0 8.11757
R1579 B.n577 B.n1 8.11757
R1580 B.n477 B.n38 1.24928
R1581 B.n464 B.n463 1.24928
R1582 B.n246 B.n117 1.24928
R1583 B.n264 B.n263 1.24928
R1584 VN VN.t0 425.661
R1585 VN VN.t1 382.664
R1586 VDD2.n149 VDD2.n77 756.745
R1587 VDD2.n72 VDD2.n0 756.745
R1588 VDD2.n150 VDD2.n149 585
R1589 VDD2.n148 VDD2.n147 585
R1590 VDD2.n81 VDD2.n80 585
R1591 VDD2.n142 VDD2.n141 585
R1592 VDD2.n140 VDD2.n139 585
R1593 VDD2.n85 VDD2.n84 585
R1594 VDD2.n134 VDD2.n133 585
R1595 VDD2.n132 VDD2.n131 585
R1596 VDD2.n89 VDD2.n88 585
R1597 VDD2.n126 VDD2.n125 585
R1598 VDD2.n124 VDD2.n91 585
R1599 VDD2.n123 VDD2.n122 585
R1600 VDD2.n94 VDD2.n92 585
R1601 VDD2.n117 VDD2.n116 585
R1602 VDD2.n115 VDD2.n114 585
R1603 VDD2.n98 VDD2.n97 585
R1604 VDD2.n109 VDD2.n108 585
R1605 VDD2.n107 VDD2.n106 585
R1606 VDD2.n102 VDD2.n101 585
R1607 VDD2.n24 VDD2.n23 585
R1608 VDD2.n29 VDD2.n28 585
R1609 VDD2.n31 VDD2.n30 585
R1610 VDD2.n20 VDD2.n19 585
R1611 VDD2.n37 VDD2.n36 585
R1612 VDD2.n39 VDD2.n38 585
R1613 VDD2.n16 VDD2.n15 585
R1614 VDD2.n46 VDD2.n45 585
R1615 VDD2.n47 VDD2.n14 585
R1616 VDD2.n49 VDD2.n48 585
R1617 VDD2.n12 VDD2.n11 585
R1618 VDD2.n55 VDD2.n54 585
R1619 VDD2.n57 VDD2.n56 585
R1620 VDD2.n8 VDD2.n7 585
R1621 VDD2.n63 VDD2.n62 585
R1622 VDD2.n65 VDD2.n64 585
R1623 VDD2.n4 VDD2.n3 585
R1624 VDD2.n71 VDD2.n70 585
R1625 VDD2.n73 VDD2.n72 585
R1626 VDD2.n25 VDD2.t0 329.036
R1627 VDD2.n103 VDD2.t1 329.036
R1628 VDD2.n149 VDD2.n148 171.744
R1629 VDD2.n148 VDD2.n80 171.744
R1630 VDD2.n141 VDD2.n80 171.744
R1631 VDD2.n141 VDD2.n140 171.744
R1632 VDD2.n140 VDD2.n84 171.744
R1633 VDD2.n133 VDD2.n84 171.744
R1634 VDD2.n133 VDD2.n132 171.744
R1635 VDD2.n132 VDD2.n88 171.744
R1636 VDD2.n125 VDD2.n88 171.744
R1637 VDD2.n125 VDD2.n124 171.744
R1638 VDD2.n124 VDD2.n123 171.744
R1639 VDD2.n123 VDD2.n92 171.744
R1640 VDD2.n116 VDD2.n92 171.744
R1641 VDD2.n116 VDD2.n115 171.744
R1642 VDD2.n115 VDD2.n97 171.744
R1643 VDD2.n108 VDD2.n97 171.744
R1644 VDD2.n108 VDD2.n107 171.744
R1645 VDD2.n107 VDD2.n101 171.744
R1646 VDD2.n29 VDD2.n23 171.744
R1647 VDD2.n30 VDD2.n29 171.744
R1648 VDD2.n30 VDD2.n19 171.744
R1649 VDD2.n37 VDD2.n19 171.744
R1650 VDD2.n38 VDD2.n37 171.744
R1651 VDD2.n38 VDD2.n15 171.744
R1652 VDD2.n46 VDD2.n15 171.744
R1653 VDD2.n47 VDD2.n46 171.744
R1654 VDD2.n48 VDD2.n47 171.744
R1655 VDD2.n48 VDD2.n11 171.744
R1656 VDD2.n55 VDD2.n11 171.744
R1657 VDD2.n56 VDD2.n55 171.744
R1658 VDD2.n56 VDD2.n7 171.744
R1659 VDD2.n63 VDD2.n7 171.744
R1660 VDD2.n64 VDD2.n63 171.744
R1661 VDD2.n64 VDD2.n3 171.744
R1662 VDD2.n71 VDD2.n3 171.744
R1663 VDD2.n72 VDD2.n71 171.744
R1664 VDD2.n154 VDD2.n76 87.5925
R1665 VDD2.t1 VDD2.n101 85.8723
R1666 VDD2.t0 VDD2.n23 85.8723
R1667 VDD2.n154 VDD2.n153 48.8641
R1668 VDD2.n126 VDD2.n91 13.1884
R1669 VDD2.n49 VDD2.n14 13.1884
R1670 VDD2.n127 VDD2.n89 12.8005
R1671 VDD2.n122 VDD2.n93 12.8005
R1672 VDD2.n45 VDD2.n44 12.8005
R1673 VDD2.n50 VDD2.n12 12.8005
R1674 VDD2.n131 VDD2.n130 12.0247
R1675 VDD2.n121 VDD2.n94 12.0247
R1676 VDD2.n43 VDD2.n16 12.0247
R1677 VDD2.n54 VDD2.n53 12.0247
R1678 VDD2.n134 VDD2.n87 11.249
R1679 VDD2.n118 VDD2.n117 11.249
R1680 VDD2.n40 VDD2.n39 11.249
R1681 VDD2.n57 VDD2.n10 11.249
R1682 VDD2.n103 VDD2.n102 10.7239
R1683 VDD2.n25 VDD2.n24 10.7239
R1684 VDD2.n135 VDD2.n85 10.4732
R1685 VDD2.n114 VDD2.n96 10.4732
R1686 VDD2.n36 VDD2.n18 10.4732
R1687 VDD2.n58 VDD2.n8 10.4732
R1688 VDD2.n139 VDD2.n138 9.69747
R1689 VDD2.n113 VDD2.n98 9.69747
R1690 VDD2.n35 VDD2.n20 9.69747
R1691 VDD2.n62 VDD2.n61 9.69747
R1692 VDD2.n153 VDD2.n152 9.45567
R1693 VDD2.n76 VDD2.n75 9.45567
R1694 VDD2.n79 VDD2.n78 9.3005
R1695 VDD2.n146 VDD2.n145 9.3005
R1696 VDD2.n144 VDD2.n143 9.3005
R1697 VDD2.n83 VDD2.n82 9.3005
R1698 VDD2.n138 VDD2.n137 9.3005
R1699 VDD2.n136 VDD2.n135 9.3005
R1700 VDD2.n87 VDD2.n86 9.3005
R1701 VDD2.n130 VDD2.n129 9.3005
R1702 VDD2.n128 VDD2.n127 9.3005
R1703 VDD2.n93 VDD2.n90 9.3005
R1704 VDD2.n121 VDD2.n120 9.3005
R1705 VDD2.n119 VDD2.n118 9.3005
R1706 VDD2.n96 VDD2.n95 9.3005
R1707 VDD2.n113 VDD2.n112 9.3005
R1708 VDD2.n111 VDD2.n110 9.3005
R1709 VDD2.n100 VDD2.n99 9.3005
R1710 VDD2.n105 VDD2.n104 9.3005
R1711 VDD2.n152 VDD2.n151 9.3005
R1712 VDD2.n2 VDD2.n1 9.3005
R1713 VDD2.n75 VDD2.n74 9.3005
R1714 VDD2.n67 VDD2.n66 9.3005
R1715 VDD2.n6 VDD2.n5 9.3005
R1716 VDD2.n61 VDD2.n60 9.3005
R1717 VDD2.n59 VDD2.n58 9.3005
R1718 VDD2.n10 VDD2.n9 9.3005
R1719 VDD2.n53 VDD2.n52 9.3005
R1720 VDD2.n51 VDD2.n50 9.3005
R1721 VDD2.n27 VDD2.n26 9.3005
R1722 VDD2.n22 VDD2.n21 9.3005
R1723 VDD2.n33 VDD2.n32 9.3005
R1724 VDD2.n35 VDD2.n34 9.3005
R1725 VDD2.n18 VDD2.n17 9.3005
R1726 VDD2.n41 VDD2.n40 9.3005
R1727 VDD2.n43 VDD2.n42 9.3005
R1728 VDD2.n44 VDD2.n13 9.3005
R1729 VDD2.n69 VDD2.n68 9.3005
R1730 VDD2.n142 VDD2.n83 8.92171
R1731 VDD2.n110 VDD2.n109 8.92171
R1732 VDD2.n32 VDD2.n31 8.92171
R1733 VDD2.n65 VDD2.n6 8.92171
R1734 VDD2.n153 VDD2.n77 8.14595
R1735 VDD2.n143 VDD2.n81 8.14595
R1736 VDD2.n106 VDD2.n100 8.14595
R1737 VDD2.n28 VDD2.n22 8.14595
R1738 VDD2.n66 VDD2.n4 8.14595
R1739 VDD2.n76 VDD2.n0 8.14595
R1740 VDD2.n151 VDD2.n150 7.3702
R1741 VDD2.n147 VDD2.n146 7.3702
R1742 VDD2.n105 VDD2.n102 7.3702
R1743 VDD2.n27 VDD2.n24 7.3702
R1744 VDD2.n70 VDD2.n69 7.3702
R1745 VDD2.n74 VDD2.n73 7.3702
R1746 VDD2.n150 VDD2.n79 6.59444
R1747 VDD2.n147 VDD2.n79 6.59444
R1748 VDD2.n70 VDD2.n2 6.59444
R1749 VDD2.n73 VDD2.n2 6.59444
R1750 VDD2.n151 VDD2.n77 5.81868
R1751 VDD2.n146 VDD2.n81 5.81868
R1752 VDD2.n106 VDD2.n105 5.81868
R1753 VDD2.n28 VDD2.n27 5.81868
R1754 VDD2.n69 VDD2.n4 5.81868
R1755 VDD2.n74 VDD2.n0 5.81868
R1756 VDD2.n143 VDD2.n142 5.04292
R1757 VDD2.n109 VDD2.n100 5.04292
R1758 VDD2.n31 VDD2.n22 5.04292
R1759 VDD2.n66 VDD2.n65 5.04292
R1760 VDD2.n139 VDD2.n83 4.26717
R1761 VDD2.n110 VDD2.n98 4.26717
R1762 VDD2.n32 VDD2.n20 4.26717
R1763 VDD2.n62 VDD2.n6 4.26717
R1764 VDD2.n138 VDD2.n85 3.49141
R1765 VDD2.n114 VDD2.n113 3.49141
R1766 VDD2.n36 VDD2.n35 3.49141
R1767 VDD2.n61 VDD2.n8 3.49141
R1768 VDD2.n135 VDD2.n134 2.71565
R1769 VDD2.n117 VDD2.n96 2.71565
R1770 VDD2.n39 VDD2.n18 2.71565
R1771 VDD2.n58 VDD2.n57 2.71565
R1772 VDD2.n104 VDD2.n103 2.41282
R1773 VDD2.n26 VDD2.n25 2.41282
R1774 VDD2.n131 VDD2.n87 1.93989
R1775 VDD2.n118 VDD2.n94 1.93989
R1776 VDD2.n40 VDD2.n16 1.93989
R1777 VDD2.n54 VDD2.n10 1.93989
R1778 VDD2.n130 VDD2.n89 1.16414
R1779 VDD2.n122 VDD2.n121 1.16414
R1780 VDD2.n45 VDD2.n43 1.16414
R1781 VDD2.n53 VDD2.n12 1.16414
R1782 VDD2 VDD2.n154 0.403517
R1783 VDD2.n127 VDD2.n126 0.388379
R1784 VDD2.n93 VDD2.n91 0.388379
R1785 VDD2.n44 VDD2.n14 0.388379
R1786 VDD2.n50 VDD2.n49 0.388379
R1787 VDD2.n152 VDD2.n78 0.155672
R1788 VDD2.n145 VDD2.n78 0.155672
R1789 VDD2.n145 VDD2.n144 0.155672
R1790 VDD2.n144 VDD2.n82 0.155672
R1791 VDD2.n137 VDD2.n82 0.155672
R1792 VDD2.n137 VDD2.n136 0.155672
R1793 VDD2.n136 VDD2.n86 0.155672
R1794 VDD2.n129 VDD2.n86 0.155672
R1795 VDD2.n129 VDD2.n128 0.155672
R1796 VDD2.n128 VDD2.n90 0.155672
R1797 VDD2.n120 VDD2.n90 0.155672
R1798 VDD2.n120 VDD2.n119 0.155672
R1799 VDD2.n119 VDD2.n95 0.155672
R1800 VDD2.n112 VDD2.n95 0.155672
R1801 VDD2.n112 VDD2.n111 0.155672
R1802 VDD2.n111 VDD2.n99 0.155672
R1803 VDD2.n104 VDD2.n99 0.155672
R1804 VDD2.n26 VDD2.n21 0.155672
R1805 VDD2.n33 VDD2.n21 0.155672
R1806 VDD2.n34 VDD2.n33 0.155672
R1807 VDD2.n34 VDD2.n17 0.155672
R1808 VDD2.n41 VDD2.n17 0.155672
R1809 VDD2.n42 VDD2.n41 0.155672
R1810 VDD2.n42 VDD2.n13 0.155672
R1811 VDD2.n51 VDD2.n13 0.155672
R1812 VDD2.n52 VDD2.n51 0.155672
R1813 VDD2.n52 VDD2.n9 0.155672
R1814 VDD2.n59 VDD2.n9 0.155672
R1815 VDD2.n60 VDD2.n59 0.155672
R1816 VDD2.n60 VDD2.n5 0.155672
R1817 VDD2.n67 VDD2.n5 0.155672
R1818 VDD2.n68 VDD2.n67 0.155672
R1819 VDD2.n68 VDD2.n1 0.155672
R1820 VDD2.n75 VDD2.n1 0.155672
C0 B VDD1 1.68415f
C1 VDD2 VDD1 0.521295f
C2 VN VDD1 0.147846f
C3 B VDD2 1.70282f
C4 VN B 0.854257f
C5 w_n1610_n3824# VDD1 1.79709f
C6 VN VDD2 2.80469f
C7 B w_n1610_n3824# 8.009851f
C8 VDD2 w_n1610_n3824# 1.80743f
C9 VDD1 VTAIL 5.84546f
C10 VN w_n1610_n3824# 2.15023f
C11 B VTAIL 3.47896f
C12 VP VDD1 2.93065f
C13 VDD2 VTAIL 5.884f
C14 VN VTAIL 2.27868f
C15 VP B 1.18137f
C16 VP VDD2 0.278001f
C17 VP VN 5.25249f
C18 w_n1610_n3824# VTAIL 3.1677f
C19 VP w_n1610_n3824# 2.35244f
C20 VP VTAIL 2.29321f
C21 VDD2 VSUBS 0.861528f
C22 VDD1 VSUBS 3.512096f
C23 VTAIL VSUBS 0.924632f
C24 VN VSUBS 8.17344f
C25 VP VSUBS 1.375117f
C26 B VSUBS 3.104628f
C27 w_n1610_n3824# VSUBS 75.5605f
C28 VDD2.n0 VSUBS 0.023176f
C29 VDD2.n1 VSUBS 0.020233f
C30 VDD2.n2 VSUBS 0.010872f
C31 VDD2.n3 VSUBS 0.025698f
C32 VDD2.n4 VSUBS 0.011512f
C33 VDD2.n5 VSUBS 0.020233f
C34 VDD2.n6 VSUBS 0.010872f
C35 VDD2.n7 VSUBS 0.025698f
C36 VDD2.n8 VSUBS 0.011512f
C37 VDD2.n9 VSUBS 0.020233f
C38 VDD2.n10 VSUBS 0.010872f
C39 VDD2.n11 VSUBS 0.025698f
C40 VDD2.n12 VSUBS 0.011512f
C41 VDD2.n13 VSUBS 0.020233f
C42 VDD2.n14 VSUBS 0.011192f
C43 VDD2.n15 VSUBS 0.025698f
C44 VDD2.n16 VSUBS 0.011512f
C45 VDD2.n17 VSUBS 0.020233f
C46 VDD2.n18 VSUBS 0.010872f
C47 VDD2.n19 VSUBS 0.025698f
C48 VDD2.n20 VSUBS 0.011512f
C49 VDD2.n21 VSUBS 0.020233f
C50 VDD2.n22 VSUBS 0.010872f
C51 VDD2.n23 VSUBS 0.019274f
C52 VDD2.n24 VSUBS 0.019332f
C53 VDD2.t0 VSUBS 0.055531f
C54 VDD2.n25 VSUBS 0.180204f
C55 VDD2.n26 VSUBS 1.19625f
C56 VDD2.n27 VSUBS 0.010872f
C57 VDD2.n28 VSUBS 0.011512f
C58 VDD2.n29 VSUBS 0.025698f
C59 VDD2.n30 VSUBS 0.025698f
C60 VDD2.n31 VSUBS 0.011512f
C61 VDD2.n32 VSUBS 0.010872f
C62 VDD2.n33 VSUBS 0.020233f
C63 VDD2.n34 VSUBS 0.020233f
C64 VDD2.n35 VSUBS 0.010872f
C65 VDD2.n36 VSUBS 0.011512f
C66 VDD2.n37 VSUBS 0.025698f
C67 VDD2.n38 VSUBS 0.025698f
C68 VDD2.n39 VSUBS 0.011512f
C69 VDD2.n40 VSUBS 0.010872f
C70 VDD2.n41 VSUBS 0.020233f
C71 VDD2.n42 VSUBS 0.020233f
C72 VDD2.n43 VSUBS 0.010872f
C73 VDD2.n44 VSUBS 0.010872f
C74 VDD2.n45 VSUBS 0.011512f
C75 VDD2.n46 VSUBS 0.025698f
C76 VDD2.n47 VSUBS 0.025698f
C77 VDD2.n48 VSUBS 0.025698f
C78 VDD2.n49 VSUBS 0.011192f
C79 VDD2.n50 VSUBS 0.010872f
C80 VDD2.n51 VSUBS 0.020233f
C81 VDD2.n52 VSUBS 0.020233f
C82 VDD2.n53 VSUBS 0.010872f
C83 VDD2.n54 VSUBS 0.011512f
C84 VDD2.n55 VSUBS 0.025698f
C85 VDD2.n56 VSUBS 0.025698f
C86 VDD2.n57 VSUBS 0.011512f
C87 VDD2.n58 VSUBS 0.010872f
C88 VDD2.n59 VSUBS 0.020233f
C89 VDD2.n60 VSUBS 0.020233f
C90 VDD2.n61 VSUBS 0.010872f
C91 VDD2.n62 VSUBS 0.011512f
C92 VDD2.n63 VSUBS 0.025698f
C93 VDD2.n64 VSUBS 0.025698f
C94 VDD2.n65 VSUBS 0.011512f
C95 VDD2.n66 VSUBS 0.010872f
C96 VDD2.n67 VSUBS 0.020233f
C97 VDD2.n68 VSUBS 0.020233f
C98 VDD2.n69 VSUBS 0.010872f
C99 VDD2.n70 VSUBS 0.011512f
C100 VDD2.n71 VSUBS 0.025698f
C101 VDD2.n72 VSUBS 0.06543f
C102 VDD2.n73 VSUBS 0.011512f
C103 VDD2.n74 VSUBS 0.010872f
C104 VDD2.n75 VSUBS 0.046768f
C105 VDD2.n76 VSUBS 0.591711f
C106 VDD2.n77 VSUBS 0.023176f
C107 VDD2.n78 VSUBS 0.020233f
C108 VDD2.n79 VSUBS 0.010872f
C109 VDD2.n80 VSUBS 0.025698f
C110 VDD2.n81 VSUBS 0.011512f
C111 VDD2.n82 VSUBS 0.020233f
C112 VDD2.n83 VSUBS 0.010872f
C113 VDD2.n84 VSUBS 0.025698f
C114 VDD2.n85 VSUBS 0.011512f
C115 VDD2.n86 VSUBS 0.020233f
C116 VDD2.n87 VSUBS 0.010872f
C117 VDD2.n88 VSUBS 0.025698f
C118 VDD2.n89 VSUBS 0.011512f
C119 VDD2.n90 VSUBS 0.020233f
C120 VDD2.n91 VSUBS 0.011192f
C121 VDD2.n92 VSUBS 0.025698f
C122 VDD2.n93 VSUBS 0.010872f
C123 VDD2.n94 VSUBS 0.011512f
C124 VDD2.n95 VSUBS 0.020233f
C125 VDD2.n96 VSUBS 0.010872f
C126 VDD2.n97 VSUBS 0.025698f
C127 VDD2.n98 VSUBS 0.011512f
C128 VDD2.n99 VSUBS 0.020233f
C129 VDD2.n100 VSUBS 0.010872f
C130 VDD2.n101 VSUBS 0.019274f
C131 VDD2.n102 VSUBS 0.019332f
C132 VDD2.t1 VSUBS 0.055531f
C133 VDD2.n103 VSUBS 0.180204f
C134 VDD2.n104 VSUBS 1.19625f
C135 VDD2.n105 VSUBS 0.010872f
C136 VDD2.n106 VSUBS 0.011512f
C137 VDD2.n107 VSUBS 0.025698f
C138 VDD2.n108 VSUBS 0.025698f
C139 VDD2.n109 VSUBS 0.011512f
C140 VDD2.n110 VSUBS 0.010872f
C141 VDD2.n111 VSUBS 0.020233f
C142 VDD2.n112 VSUBS 0.020233f
C143 VDD2.n113 VSUBS 0.010872f
C144 VDD2.n114 VSUBS 0.011512f
C145 VDD2.n115 VSUBS 0.025698f
C146 VDD2.n116 VSUBS 0.025698f
C147 VDD2.n117 VSUBS 0.011512f
C148 VDD2.n118 VSUBS 0.010872f
C149 VDD2.n119 VSUBS 0.020233f
C150 VDD2.n120 VSUBS 0.020233f
C151 VDD2.n121 VSUBS 0.010872f
C152 VDD2.n122 VSUBS 0.011512f
C153 VDD2.n123 VSUBS 0.025698f
C154 VDD2.n124 VSUBS 0.025698f
C155 VDD2.n125 VSUBS 0.025698f
C156 VDD2.n126 VSUBS 0.011192f
C157 VDD2.n127 VSUBS 0.010872f
C158 VDD2.n128 VSUBS 0.020233f
C159 VDD2.n129 VSUBS 0.020233f
C160 VDD2.n130 VSUBS 0.010872f
C161 VDD2.n131 VSUBS 0.011512f
C162 VDD2.n132 VSUBS 0.025698f
C163 VDD2.n133 VSUBS 0.025698f
C164 VDD2.n134 VSUBS 0.011512f
C165 VDD2.n135 VSUBS 0.010872f
C166 VDD2.n136 VSUBS 0.020233f
C167 VDD2.n137 VSUBS 0.020233f
C168 VDD2.n138 VSUBS 0.010872f
C169 VDD2.n139 VSUBS 0.011512f
C170 VDD2.n140 VSUBS 0.025698f
C171 VDD2.n141 VSUBS 0.025698f
C172 VDD2.n142 VSUBS 0.011512f
C173 VDD2.n143 VSUBS 0.010872f
C174 VDD2.n144 VSUBS 0.020233f
C175 VDD2.n145 VSUBS 0.020233f
C176 VDD2.n146 VSUBS 0.010872f
C177 VDD2.n147 VSUBS 0.011512f
C178 VDD2.n148 VSUBS 0.025698f
C179 VDD2.n149 VSUBS 0.06543f
C180 VDD2.n150 VSUBS 0.011512f
C181 VDD2.n151 VSUBS 0.010872f
C182 VDD2.n152 VSUBS 0.046768f
C183 VDD2.n153 VSUBS 0.047018f
C184 VDD2.n154 VSUBS 2.45179f
C185 VN.t1 VSUBS 3.02839f
C186 VN.t0 VSUBS 3.35655f
C187 B.n0 VSUBS 0.005826f
C188 B.n1 VSUBS 0.005826f
C189 B.n2 VSUBS 0.008616f
C190 B.n3 VSUBS 0.006603f
C191 B.n4 VSUBS 0.006603f
C192 B.n5 VSUBS 0.006603f
C193 B.n6 VSUBS 0.006603f
C194 B.n7 VSUBS 0.006603f
C195 B.n8 VSUBS 0.006603f
C196 B.n9 VSUBS 0.006603f
C197 B.n10 VSUBS 0.015524f
C198 B.n11 VSUBS 0.006603f
C199 B.n12 VSUBS 0.006603f
C200 B.n13 VSUBS 0.006603f
C201 B.n14 VSUBS 0.006603f
C202 B.n15 VSUBS 0.006603f
C203 B.n16 VSUBS 0.006603f
C204 B.n17 VSUBS 0.006603f
C205 B.n18 VSUBS 0.006603f
C206 B.n19 VSUBS 0.006603f
C207 B.n20 VSUBS 0.006603f
C208 B.n21 VSUBS 0.006603f
C209 B.n22 VSUBS 0.006603f
C210 B.n23 VSUBS 0.006603f
C211 B.n24 VSUBS 0.006603f
C212 B.n25 VSUBS 0.006603f
C213 B.n26 VSUBS 0.006603f
C214 B.n27 VSUBS 0.006603f
C215 B.n28 VSUBS 0.006603f
C216 B.n29 VSUBS 0.006603f
C217 B.n30 VSUBS 0.006603f
C218 B.n31 VSUBS 0.006603f
C219 B.n32 VSUBS 0.006603f
C220 B.n33 VSUBS 0.006603f
C221 B.n34 VSUBS 0.006214f
C222 B.n35 VSUBS 0.006603f
C223 B.t1 VSUBS 0.248188f
C224 B.t2 VSUBS 0.265613f
C225 B.t0 VSUBS 0.729591f
C226 B.n36 VSUBS 0.381196f
C227 B.n37 VSUBS 0.260963f
C228 B.n38 VSUBS 0.015298f
C229 B.n39 VSUBS 0.006603f
C230 B.n40 VSUBS 0.006603f
C231 B.n41 VSUBS 0.006603f
C232 B.n42 VSUBS 0.006603f
C233 B.t10 VSUBS 0.248191f
C234 B.t11 VSUBS 0.265616f
C235 B.t9 VSUBS 0.729591f
C236 B.n43 VSUBS 0.381194f
C237 B.n44 VSUBS 0.26096f
C238 B.n45 VSUBS 0.006603f
C239 B.n46 VSUBS 0.006603f
C240 B.n47 VSUBS 0.006603f
C241 B.n48 VSUBS 0.006603f
C242 B.n49 VSUBS 0.006603f
C243 B.n50 VSUBS 0.006603f
C244 B.n51 VSUBS 0.006603f
C245 B.n52 VSUBS 0.006603f
C246 B.n53 VSUBS 0.006603f
C247 B.n54 VSUBS 0.006603f
C248 B.n55 VSUBS 0.006603f
C249 B.n56 VSUBS 0.006603f
C250 B.n57 VSUBS 0.006603f
C251 B.n58 VSUBS 0.006603f
C252 B.n59 VSUBS 0.006603f
C253 B.n60 VSUBS 0.006603f
C254 B.n61 VSUBS 0.006603f
C255 B.n62 VSUBS 0.006603f
C256 B.n63 VSUBS 0.006603f
C257 B.n64 VSUBS 0.006603f
C258 B.n65 VSUBS 0.006603f
C259 B.n66 VSUBS 0.006603f
C260 B.n67 VSUBS 0.006603f
C261 B.n68 VSUBS 0.01613f
C262 B.n69 VSUBS 0.006603f
C263 B.n70 VSUBS 0.006603f
C264 B.n71 VSUBS 0.006603f
C265 B.n72 VSUBS 0.006603f
C266 B.n73 VSUBS 0.006603f
C267 B.n74 VSUBS 0.006603f
C268 B.n75 VSUBS 0.006603f
C269 B.n76 VSUBS 0.006603f
C270 B.n77 VSUBS 0.006603f
C271 B.n78 VSUBS 0.006603f
C272 B.n79 VSUBS 0.006603f
C273 B.n80 VSUBS 0.006603f
C274 B.n81 VSUBS 0.006603f
C275 B.n82 VSUBS 0.006603f
C276 B.n83 VSUBS 0.006603f
C277 B.n84 VSUBS 0.006603f
C278 B.n85 VSUBS 0.006603f
C279 B.n86 VSUBS 0.015524f
C280 B.n87 VSUBS 0.006603f
C281 B.n88 VSUBS 0.006603f
C282 B.n89 VSUBS 0.006603f
C283 B.n90 VSUBS 0.006603f
C284 B.n91 VSUBS 0.006603f
C285 B.n92 VSUBS 0.006603f
C286 B.n93 VSUBS 0.006603f
C287 B.n94 VSUBS 0.006603f
C288 B.n95 VSUBS 0.006603f
C289 B.n96 VSUBS 0.006603f
C290 B.n97 VSUBS 0.006603f
C291 B.n98 VSUBS 0.006603f
C292 B.n99 VSUBS 0.006603f
C293 B.n100 VSUBS 0.006603f
C294 B.n101 VSUBS 0.006603f
C295 B.n102 VSUBS 0.006603f
C296 B.n103 VSUBS 0.006603f
C297 B.n104 VSUBS 0.006603f
C298 B.n105 VSUBS 0.006603f
C299 B.n106 VSUBS 0.006603f
C300 B.n107 VSUBS 0.006603f
C301 B.n108 VSUBS 0.006603f
C302 B.n109 VSUBS 0.006603f
C303 B.n110 VSUBS 0.006603f
C304 B.t8 VSUBS 0.248191f
C305 B.t7 VSUBS 0.265616f
C306 B.t6 VSUBS 0.729591f
C307 B.n111 VSUBS 0.381194f
C308 B.n112 VSUBS 0.26096f
C309 B.n113 VSUBS 0.006603f
C310 B.n114 VSUBS 0.006603f
C311 B.n115 VSUBS 0.006603f
C312 B.n116 VSUBS 0.006603f
C313 B.n117 VSUBS 0.00369f
C314 B.n118 VSUBS 0.006603f
C315 B.n119 VSUBS 0.006603f
C316 B.n120 VSUBS 0.006603f
C317 B.n121 VSUBS 0.006603f
C318 B.n122 VSUBS 0.006603f
C319 B.n123 VSUBS 0.006603f
C320 B.n124 VSUBS 0.006603f
C321 B.n125 VSUBS 0.006603f
C322 B.n126 VSUBS 0.006603f
C323 B.n127 VSUBS 0.006603f
C324 B.n128 VSUBS 0.006603f
C325 B.n129 VSUBS 0.006603f
C326 B.n130 VSUBS 0.006603f
C327 B.n131 VSUBS 0.006603f
C328 B.n132 VSUBS 0.006603f
C329 B.n133 VSUBS 0.006603f
C330 B.n134 VSUBS 0.006603f
C331 B.n135 VSUBS 0.006603f
C332 B.n136 VSUBS 0.006603f
C333 B.n137 VSUBS 0.006603f
C334 B.n138 VSUBS 0.006603f
C335 B.n139 VSUBS 0.006603f
C336 B.n140 VSUBS 0.006603f
C337 B.n141 VSUBS 0.01613f
C338 B.n142 VSUBS 0.006603f
C339 B.n143 VSUBS 0.006603f
C340 B.n144 VSUBS 0.006603f
C341 B.n145 VSUBS 0.006603f
C342 B.n146 VSUBS 0.006603f
C343 B.n147 VSUBS 0.006603f
C344 B.n148 VSUBS 0.006603f
C345 B.n149 VSUBS 0.006603f
C346 B.n150 VSUBS 0.006603f
C347 B.n151 VSUBS 0.006603f
C348 B.n152 VSUBS 0.006603f
C349 B.n153 VSUBS 0.006603f
C350 B.n154 VSUBS 0.006603f
C351 B.n155 VSUBS 0.006603f
C352 B.n156 VSUBS 0.006603f
C353 B.n157 VSUBS 0.006603f
C354 B.n158 VSUBS 0.006603f
C355 B.n159 VSUBS 0.006603f
C356 B.n160 VSUBS 0.006603f
C357 B.n161 VSUBS 0.006603f
C358 B.n162 VSUBS 0.006603f
C359 B.n163 VSUBS 0.006603f
C360 B.n164 VSUBS 0.006603f
C361 B.n165 VSUBS 0.006603f
C362 B.n166 VSUBS 0.006603f
C363 B.n167 VSUBS 0.006603f
C364 B.n168 VSUBS 0.006603f
C365 B.n169 VSUBS 0.006603f
C366 B.n170 VSUBS 0.006603f
C367 B.n171 VSUBS 0.006603f
C368 B.n172 VSUBS 0.015524f
C369 B.n173 VSUBS 0.015524f
C370 B.n174 VSUBS 0.01613f
C371 B.n175 VSUBS 0.006603f
C372 B.n176 VSUBS 0.006603f
C373 B.n177 VSUBS 0.006603f
C374 B.n178 VSUBS 0.006603f
C375 B.n179 VSUBS 0.006603f
C376 B.n180 VSUBS 0.006603f
C377 B.n181 VSUBS 0.006603f
C378 B.n182 VSUBS 0.006603f
C379 B.n183 VSUBS 0.006603f
C380 B.n184 VSUBS 0.006603f
C381 B.n185 VSUBS 0.006603f
C382 B.n186 VSUBS 0.006603f
C383 B.n187 VSUBS 0.006603f
C384 B.n188 VSUBS 0.006603f
C385 B.n189 VSUBS 0.006603f
C386 B.n190 VSUBS 0.006603f
C387 B.n191 VSUBS 0.006603f
C388 B.n192 VSUBS 0.006603f
C389 B.n193 VSUBS 0.006603f
C390 B.n194 VSUBS 0.006603f
C391 B.n195 VSUBS 0.006603f
C392 B.n196 VSUBS 0.006603f
C393 B.n197 VSUBS 0.006603f
C394 B.n198 VSUBS 0.006603f
C395 B.n199 VSUBS 0.006603f
C396 B.n200 VSUBS 0.006603f
C397 B.n201 VSUBS 0.006603f
C398 B.n202 VSUBS 0.006603f
C399 B.n203 VSUBS 0.006603f
C400 B.n204 VSUBS 0.006603f
C401 B.n205 VSUBS 0.006603f
C402 B.n206 VSUBS 0.006603f
C403 B.n207 VSUBS 0.006603f
C404 B.n208 VSUBS 0.006603f
C405 B.n209 VSUBS 0.006603f
C406 B.n210 VSUBS 0.006603f
C407 B.n211 VSUBS 0.006603f
C408 B.n212 VSUBS 0.006603f
C409 B.n213 VSUBS 0.006603f
C410 B.n214 VSUBS 0.006603f
C411 B.n215 VSUBS 0.006603f
C412 B.n216 VSUBS 0.006603f
C413 B.n217 VSUBS 0.006603f
C414 B.n218 VSUBS 0.006603f
C415 B.n219 VSUBS 0.006603f
C416 B.n220 VSUBS 0.006603f
C417 B.n221 VSUBS 0.006603f
C418 B.n222 VSUBS 0.006603f
C419 B.n223 VSUBS 0.006603f
C420 B.n224 VSUBS 0.006603f
C421 B.n225 VSUBS 0.006603f
C422 B.n226 VSUBS 0.006603f
C423 B.n227 VSUBS 0.006603f
C424 B.n228 VSUBS 0.006603f
C425 B.n229 VSUBS 0.006603f
C426 B.n230 VSUBS 0.006603f
C427 B.n231 VSUBS 0.006603f
C428 B.n232 VSUBS 0.006603f
C429 B.n233 VSUBS 0.006603f
C430 B.n234 VSUBS 0.006603f
C431 B.n235 VSUBS 0.006603f
C432 B.n236 VSUBS 0.006603f
C433 B.n237 VSUBS 0.006603f
C434 B.n238 VSUBS 0.006603f
C435 B.n239 VSUBS 0.006603f
C436 B.n240 VSUBS 0.006603f
C437 B.n241 VSUBS 0.006603f
C438 B.n242 VSUBS 0.006603f
C439 B.n243 VSUBS 0.006603f
C440 B.t5 VSUBS 0.248188f
C441 B.t4 VSUBS 0.265613f
C442 B.t3 VSUBS 0.729591f
C443 B.n244 VSUBS 0.381196f
C444 B.n245 VSUBS 0.260963f
C445 B.n246 VSUBS 0.015298f
C446 B.n247 VSUBS 0.006214f
C447 B.n248 VSUBS 0.006603f
C448 B.n249 VSUBS 0.006603f
C449 B.n250 VSUBS 0.006603f
C450 B.n251 VSUBS 0.006603f
C451 B.n252 VSUBS 0.006603f
C452 B.n253 VSUBS 0.006603f
C453 B.n254 VSUBS 0.006603f
C454 B.n255 VSUBS 0.006603f
C455 B.n256 VSUBS 0.006603f
C456 B.n257 VSUBS 0.006603f
C457 B.n258 VSUBS 0.006603f
C458 B.n259 VSUBS 0.006603f
C459 B.n260 VSUBS 0.006603f
C460 B.n261 VSUBS 0.006603f
C461 B.n262 VSUBS 0.006603f
C462 B.n263 VSUBS 0.00369f
C463 B.n264 VSUBS 0.015298f
C464 B.n265 VSUBS 0.006214f
C465 B.n266 VSUBS 0.006603f
C466 B.n267 VSUBS 0.006603f
C467 B.n268 VSUBS 0.006603f
C468 B.n269 VSUBS 0.006603f
C469 B.n270 VSUBS 0.006603f
C470 B.n271 VSUBS 0.006603f
C471 B.n272 VSUBS 0.006603f
C472 B.n273 VSUBS 0.006603f
C473 B.n274 VSUBS 0.006603f
C474 B.n275 VSUBS 0.006603f
C475 B.n276 VSUBS 0.006603f
C476 B.n277 VSUBS 0.006603f
C477 B.n278 VSUBS 0.006603f
C478 B.n279 VSUBS 0.006603f
C479 B.n280 VSUBS 0.006603f
C480 B.n281 VSUBS 0.006603f
C481 B.n282 VSUBS 0.006603f
C482 B.n283 VSUBS 0.006603f
C483 B.n284 VSUBS 0.006603f
C484 B.n285 VSUBS 0.006603f
C485 B.n286 VSUBS 0.006603f
C486 B.n287 VSUBS 0.006603f
C487 B.n288 VSUBS 0.006603f
C488 B.n289 VSUBS 0.006603f
C489 B.n290 VSUBS 0.006603f
C490 B.n291 VSUBS 0.006603f
C491 B.n292 VSUBS 0.006603f
C492 B.n293 VSUBS 0.006603f
C493 B.n294 VSUBS 0.006603f
C494 B.n295 VSUBS 0.006603f
C495 B.n296 VSUBS 0.006603f
C496 B.n297 VSUBS 0.006603f
C497 B.n298 VSUBS 0.006603f
C498 B.n299 VSUBS 0.006603f
C499 B.n300 VSUBS 0.006603f
C500 B.n301 VSUBS 0.006603f
C501 B.n302 VSUBS 0.006603f
C502 B.n303 VSUBS 0.006603f
C503 B.n304 VSUBS 0.006603f
C504 B.n305 VSUBS 0.006603f
C505 B.n306 VSUBS 0.006603f
C506 B.n307 VSUBS 0.006603f
C507 B.n308 VSUBS 0.006603f
C508 B.n309 VSUBS 0.006603f
C509 B.n310 VSUBS 0.006603f
C510 B.n311 VSUBS 0.006603f
C511 B.n312 VSUBS 0.006603f
C512 B.n313 VSUBS 0.006603f
C513 B.n314 VSUBS 0.006603f
C514 B.n315 VSUBS 0.006603f
C515 B.n316 VSUBS 0.006603f
C516 B.n317 VSUBS 0.006603f
C517 B.n318 VSUBS 0.006603f
C518 B.n319 VSUBS 0.006603f
C519 B.n320 VSUBS 0.006603f
C520 B.n321 VSUBS 0.006603f
C521 B.n322 VSUBS 0.006603f
C522 B.n323 VSUBS 0.006603f
C523 B.n324 VSUBS 0.006603f
C524 B.n325 VSUBS 0.006603f
C525 B.n326 VSUBS 0.006603f
C526 B.n327 VSUBS 0.006603f
C527 B.n328 VSUBS 0.006603f
C528 B.n329 VSUBS 0.006603f
C529 B.n330 VSUBS 0.006603f
C530 B.n331 VSUBS 0.006603f
C531 B.n332 VSUBS 0.006603f
C532 B.n333 VSUBS 0.006603f
C533 B.n334 VSUBS 0.006603f
C534 B.n335 VSUBS 0.01613f
C535 B.n336 VSUBS 0.015378f
C536 B.n337 VSUBS 0.016277f
C537 B.n338 VSUBS 0.006603f
C538 B.n339 VSUBS 0.006603f
C539 B.n340 VSUBS 0.006603f
C540 B.n341 VSUBS 0.006603f
C541 B.n342 VSUBS 0.006603f
C542 B.n343 VSUBS 0.006603f
C543 B.n344 VSUBS 0.006603f
C544 B.n345 VSUBS 0.006603f
C545 B.n346 VSUBS 0.006603f
C546 B.n347 VSUBS 0.006603f
C547 B.n348 VSUBS 0.006603f
C548 B.n349 VSUBS 0.006603f
C549 B.n350 VSUBS 0.006603f
C550 B.n351 VSUBS 0.006603f
C551 B.n352 VSUBS 0.006603f
C552 B.n353 VSUBS 0.006603f
C553 B.n354 VSUBS 0.006603f
C554 B.n355 VSUBS 0.006603f
C555 B.n356 VSUBS 0.006603f
C556 B.n357 VSUBS 0.006603f
C557 B.n358 VSUBS 0.006603f
C558 B.n359 VSUBS 0.006603f
C559 B.n360 VSUBS 0.006603f
C560 B.n361 VSUBS 0.006603f
C561 B.n362 VSUBS 0.006603f
C562 B.n363 VSUBS 0.006603f
C563 B.n364 VSUBS 0.006603f
C564 B.n365 VSUBS 0.006603f
C565 B.n366 VSUBS 0.006603f
C566 B.n367 VSUBS 0.006603f
C567 B.n368 VSUBS 0.006603f
C568 B.n369 VSUBS 0.006603f
C569 B.n370 VSUBS 0.006603f
C570 B.n371 VSUBS 0.006603f
C571 B.n372 VSUBS 0.006603f
C572 B.n373 VSUBS 0.006603f
C573 B.n374 VSUBS 0.006603f
C574 B.n375 VSUBS 0.006603f
C575 B.n376 VSUBS 0.006603f
C576 B.n377 VSUBS 0.006603f
C577 B.n378 VSUBS 0.006603f
C578 B.n379 VSUBS 0.006603f
C579 B.n380 VSUBS 0.006603f
C580 B.n381 VSUBS 0.006603f
C581 B.n382 VSUBS 0.006603f
C582 B.n383 VSUBS 0.006603f
C583 B.n384 VSUBS 0.006603f
C584 B.n385 VSUBS 0.006603f
C585 B.n386 VSUBS 0.006603f
C586 B.n387 VSUBS 0.006603f
C587 B.n388 VSUBS 0.006603f
C588 B.n389 VSUBS 0.015524f
C589 B.n390 VSUBS 0.015524f
C590 B.n391 VSUBS 0.01613f
C591 B.n392 VSUBS 0.006603f
C592 B.n393 VSUBS 0.006603f
C593 B.n394 VSUBS 0.006603f
C594 B.n395 VSUBS 0.006603f
C595 B.n396 VSUBS 0.006603f
C596 B.n397 VSUBS 0.006603f
C597 B.n398 VSUBS 0.006603f
C598 B.n399 VSUBS 0.006603f
C599 B.n400 VSUBS 0.006603f
C600 B.n401 VSUBS 0.006603f
C601 B.n402 VSUBS 0.006603f
C602 B.n403 VSUBS 0.006603f
C603 B.n404 VSUBS 0.006603f
C604 B.n405 VSUBS 0.006603f
C605 B.n406 VSUBS 0.006603f
C606 B.n407 VSUBS 0.006603f
C607 B.n408 VSUBS 0.006603f
C608 B.n409 VSUBS 0.006603f
C609 B.n410 VSUBS 0.006603f
C610 B.n411 VSUBS 0.006603f
C611 B.n412 VSUBS 0.006603f
C612 B.n413 VSUBS 0.006603f
C613 B.n414 VSUBS 0.006603f
C614 B.n415 VSUBS 0.006603f
C615 B.n416 VSUBS 0.006603f
C616 B.n417 VSUBS 0.006603f
C617 B.n418 VSUBS 0.006603f
C618 B.n419 VSUBS 0.006603f
C619 B.n420 VSUBS 0.006603f
C620 B.n421 VSUBS 0.006603f
C621 B.n422 VSUBS 0.006603f
C622 B.n423 VSUBS 0.006603f
C623 B.n424 VSUBS 0.006603f
C624 B.n425 VSUBS 0.006603f
C625 B.n426 VSUBS 0.006603f
C626 B.n427 VSUBS 0.006603f
C627 B.n428 VSUBS 0.006603f
C628 B.n429 VSUBS 0.006603f
C629 B.n430 VSUBS 0.006603f
C630 B.n431 VSUBS 0.006603f
C631 B.n432 VSUBS 0.006603f
C632 B.n433 VSUBS 0.006603f
C633 B.n434 VSUBS 0.006603f
C634 B.n435 VSUBS 0.006603f
C635 B.n436 VSUBS 0.006603f
C636 B.n437 VSUBS 0.006603f
C637 B.n438 VSUBS 0.006603f
C638 B.n439 VSUBS 0.006603f
C639 B.n440 VSUBS 0.006603f
C640 B.n441 VSUBS 0.006603f
C641 B.n442 VSUBS 0.006603f
C642 B.n443 VSUBS 0.006603f
C643 B.n444 VSUBS 0.006603f
C644 B.n445 VSUBS 0.006603f
C645 B.n446 VSUBS 0.006603f
C646 B.n447 VSUBS 0.006603f
C647 B.n448 VSUBS 0.006603f
C648 B.n449 VSUBS 0.006603f
C649 B.n450 VSUBS 0.006603f
C650 B.n451 VSUBS 0.006603f
C651 B.n452 VSUBS 0.006603f
C652 B.n453 VSUBS 0.006603f
C653 B.n454 VSUBS 0.006603f
C654 B.n455 VSUBS 0.006603f
C655 B.n456 VSUBS 0.006603f
C656 B.n457 VSUBS 0.006603f
C657 B.n458 VSUBS 0.006603f
C658 B.n459 VSUBS 0.006603f
C659 B.n460 VSUBS 0.006603f
C660 B.n461 VSUBS 0.006603f
C661 B.n462 VSUBS 0.006214f
C662 B.n463 VSUBS 0.015298f
C663 B.n464 VSUBS 0.00369f
C664 B.n465 VSUBS 0.006603f
C665 B.n466 VSUBS 0.006603f
C666 B.n467 VSUBS 0.006603f
C667 B.n468 VSUBS 0.006603f
C668 B.n469 VSUBS 0.006603f
C669 B.n470 VSUBS 0.006603f
C670 B.n471 VSUBS 0.006603f
C671 B.n472 VSUBS 0.006603f
C672 B.n473 VSUBS 0.006603f
C673 B.n474 VSUBS 0.006603f
C674 B.n475 VSUBS 0.006603f
C675 B.n476 VSUBS 0.006603f
C676 B.n477 VSUBS 0.00369f
C677 B.n478 VSUBS 0.006603f
C678 B.n479 VSUBS 0.006603f
C679 B.n480 VSUBS 0.006603f
C680 B.n481 VSUBS 0.006603f
C681 B.n482 VSUBS 0.006603f
C682 B.n483 VSUBS 0.006603f
C683 B.n484 VSUBS 0.006603f
C684 B.n485 VSUBS 0.006603f
C685 B.n486 VSUBS 0.006603f
C686 B.n487 VSUBS 0.006603f
C687 B.n488 VSUBS 0.006603f
C688 B.n489 VSUBS 0.006603f
C689 B.n490 VSUBS 0.006603f
C690 B.n491 VSUBS 0.006603f
C691 B.n492 VSUBS 0.006603f
C692 B.n493 VSUBS 0.006603f
C693 B.n494 VSUBS 0.006603f
C694 B.n495 VSUBS 0.006603f
C695 B.n496 VSUBS 0.006603f
C696 B.n497 VSUBS 0.006603f
C697 B.n498 VSUBS 0.006603f
C698 B.n499 VSUBS 0.006603f
C699 B.n500 VSUBS 0.006603f
C700 B.n501 VSUBS 0.006603f
C701 B.n502 VSUBS 0.006603f
C702 B.n503 VSUBS 0.006603f
C703 B.n504 VSUBS 0.006603f
C704 B.n505 VSUBS 0.006603f
C705 B.n506 VSUBS 0.006603f
C706 B.n507 VSUBS 0.006603f
C707 B.n508 VSUBS 0.006603f
C708 B.n509 VSUBS 0.006603f
C709 B.n510 VSUBS 0.006603f
C710 B.n511 VSUBS 0.006603f
C711 B.n512 VSUBS 0.006603f
C712 B.n513 VSUBS 0.006603f
C713 B.n514 VSUBS 0.006603f
C714 B.n515 VSUBS 0.006603f
C715 B.n516 VSUBS 0.006603f
C716 B.n517 VSUBS 0.006603f
C717 B.n518 VSUBS 0.006603f
C718 B.n519 VSUBS 0.006603f
C719 B.n520 VSUBS 0.006603f
C720 B.n521 VSUBS 0.006603f
C721 B.n522 VSUBS 0.006603f
C722 B.n523 VSUBS 0.006603f
C723 B.n524 VSUBS 0.006603f
C724 B.n525 VSUBS 0.006603f
C725 B.n526 VSUBS 0.006603f
C726 B.n527 VSUBS 0.006603f
C727 B.n528 VSUBS 0.006603f
C728 B.n529 VSUBS 0.006603f
C729 B.n530 VSUBS 0.006603f
C730 B.n531 VSUBS 0.006603f
C731 B.n532 VSUBS 0.006603f
C732 B.n533 VSUBS 0.006603f
C733 B.n534 VSUBS 0.006603f
C734 B.n535 VSUBS 0.006603f
C735 B.n536 VSUBS 0.006603f
C736 B.n537 VSUBS 0.006603f
C737 B.n538 VSUBS 0.006603f
C738 B.n539 VSUBS 0.006603f
C739 B.n540 VSUBS 0.006603f
C740 B.n541 VSUBS 0.006603f
C741 B.n542 VSUBS 0.006603f
C742 B.n543 VSUBS 0.006603f
C743 B.n544 VSUBS 0.006603f
C744 B.n545 VSUBS 0.006603f
C745 B.n546 VSUBS 0.006603f
C746 B.n547 VSUBS 0.006603f
C747 B.n548 VSUBS 0.006603f
C748 B.n549 VSUBS 0.01613f
C749 B.n550 VSUBS 0.01613f
C750 B.n551 VSUBS 0.015524f
C751 B.n552 VSUBS 0.006603f
C752 B.n553 VSUBS 0.006603f
C753 B.n554 VSUBS 0.006603f
C754 B.n555 VSUBS 0.006603f
C755 B.n556 VSUBS 0.006603f
C756 B.n557 VSUBS 0.006603f
C757 B.n558 VSUBS 0.006603f
C758 B.n559 VSUBS 0.006603f
C759 B.n560 VSUBS 0.006603f
C760 B.n561 VSUBS 0.006603f
C761 B.n562 VSUBS 0.006603f
C762 B.n563 VSUBS 0.006603f
C763 B.n564 VSUBS 0.006603f
C764 B.n565 VSUBS 0.006603f
C765 B.n566 VSUBS 0.006603f
C766 B.n567 VSUBS 0.006603f
C767 B.n568 VSUBS 0.006603f
C768 B.n569 VSUBS 0.006603f
C769 B.n570 VSUBS 0.006603f
C770 B.n571 VSUBS 0.006603f
C771 B.n572 VSUBS 0.006603f
C772 B.n573 VSUBS 0.006603f
C773 B.n574 VSUBS 0.006603f
C774 B.n575 VSUBS 0.008616f
C775 B.n576 VSUBS 0.009179f
C776 B.n577 VSUBS 0.018252f
C777 VDD1.n0 VSUBS 0.022979f
C778 VDD1.n1 VSUBS 0.020061f
C779 VDD1.n2 VSUBS 0.01078f
C780 VDD1.n3 VSUBS 0.025479f
C781 VDD1.n4 VSUBS 0.011414f
C782 VDD1.n5 VSUBS 0.020061f
C783 VDD1.n6 VSUBS 0.01078f
C784 VDD1.n7 VSUBS 0.025479f
C785 VDD1.n8 VSUBS 0.011414f
C786 VDD1.n9 VSUBS 0.020061f
C787 VDD1.n10 VSUBS 0.01078f
C788 VDD1.n11 VSUBS 0.025479f
C789 VDD1.n12 VSUBS 0.011414f
C790 VDD1.n13 VSUBS 0.020061f
C791 VDD1.n14 VSUBS 0.011097f
C792 VDD1.n15 VSUBS 0.025479f
C793 VDD1.n16 VSUBS 0.01078f
C794 VDD1.n17 VSUBS 0.011414f
C795 VDD1.n18 VSUBS 0.020061f
C796 VDD1.n19 VSUBS 0.01078f
C797 VDD1.n20 VSUBS 0.025479f
C798 VDD1.n21 VSUBS 0.011414f
C799 VDD1.n22 VSUBS 0.020061f
C800 VDD1.n23 VSUBS 0.01078f
C801 VDD1.n24 VSUBS 0.01911f
C802 VDD1.n25 VSUBS 0.019167f
C803 VDD1.t0 VSUBS 0.055058f
C804 VDD1.n26 VSUBS 0.178669f
C805 VDD1.n27 VSUBS 1.18606f
C806 VDD1.n28 VSUBS 0.01078f
C807 VDD1.n29 VSUBS 0.011414f
C808 VDD1.n30 VSUBS 0.025479f
C809 VDD1.n31 VSUBS 0.025479f
C810 VDD1.n32 VSUBS 0.011414f
C811 VDD1.n33 VSUBS 0.01078f
C812 VDD1.n34 VSUBS 0.020061f
C813 VDD1.n35 VSUBS 0.020061f
C814 VDD1.n36 VSUBS 0.01078f
C815 VDD1.n37 VSUBS 0.011414f
C816 VDD1.n38 VSUBS 0.025479f
C817 VDD1.n39 VSUBS 0.025479f
C818 VDD1.n40 VSUBS 0.011414f
C819 VDD1.n41 VSUBS 0.01078f
C820 VDD1.n42 VSUBS 0.020061f
C821 VDD1.n43 VSUBS 0.020061f
C822 VDD1.n44 VSUBS 0.01078f
C823 VDD1.n45 VSUBS 0.011414f
C824 VDD1.n46 VSUBS 0.025479f
C825 VDD1.n47 VSUBS 0.025479f
C826 VDD1.n48 VSUBS 0.025479f
C827 VDD1.n49 VSUBS 0.011097f
C828 VDD1.n50 VSUBS 0.01078f
C829 VDD1.n51 VSUBS 0.020061f
C830 VDD1.n52 VSUBS 0.020061f
C831 VDD1.n53 VSUBS 0.01078f
C832 VDD1.n54 VSUBS 0.011414f
C833 VDD1.n55 VSUBS 0.025479f
C834 VDD1.n56 VSUBS 0.025479f
C835 VDD1.n57 VSUBS 0.011414f
C836 VDD1.n58 VSUBS 0.01078f
C837 VDD1.n59 VSUBS 0.020061f
C838 VDD1.n60 VSUBS 0.020061f
C839 VDD1.n61 VSUBS 0.01078f
C840 VDD1.n62 VSUBS 0.011414f
C841 VDD1.n63 VSUBS 0.025479f
C842 VDD1.n64 VSUBS 0.025479f
C843 VDD1.n65 VSUBS 0.011414f
C844 VDD1.n66 VSUBS 0.01078f
C845 VDD1.n67 VSUBS 0.020061f
C846 VDD1.n68 VSUBS 0.020061f
C847 VDD1.n69 VSUBS 0.01078f
C848 VDD1.n70 VSUBS 0.011414f
C849 VDD1.n71 VSUBS 0.025479f
C850 VDD1.n72 VSUBS 0.064873f
C851 VDD1.n73 VSUBS 0.011414f
C852 VDD1.n74 VSUBS 0.01078f
C853 VDD1.n75 VSUBS 0.046369f
C854 VDD1.n76 VSUBS 0.047146f
C855 VDD1.n77 VSUBS 0.022979f
C856 VDD1.n78 VSUBS 0.020061f
C857 VDD1.n79 VSUBS 0.01078f
C858 VDD1.n80 VSUBS 0.025479f
C859 VDD1.n81 VSUBS 0.011414f
C860 VDD1.n82 VSUBS 0.020061f
C861 VDD1.n83 VSUBS 0.01078f
C862 VDD1.n84 VSUBS 0.025479f
C863 VDD1.n85 VSUBS 0.011414f
C864 VDD1.n86 VSUBS 0.020061f
C865 VDD1.n87 VSUBS 0.01078f
C866 VDD1.n88 VSUBS 0.025479f
C867 VDD1.n89 VSUBS 0.011414f
C868 VDD1.n90 VSUBS 0.020061f
C869 VDD1.n91 VSUBS 0.011097f
C870 VDD1.n92 VSUBS 0.025479f
C871 VDD1.n93 VSUBS 0.011414f
C872 VDD1.n94 VSUBS 0.020061f
C873 VDD1.n95 VSUBS 0.01078f
C874 VDD1.n96 VSUBS 0.025479f
C875 VDD1.n97 VSUBS 0.011414f
C876 VDD1.n98 VSUBS 0.020061f
C877 VDD1.n99 VSUBS 0.01078f
C878 VDD1.n100 VSUBS 0.01911f
C879 VDD1.n101 VSUBS 0.019167f
C880 VDD1.t1 VSUBS 0.055058f
C881 VDD1.n102 VSUBS 0.178669f
C882 VDD1.n103 VSUBS 1.18606f
C883 VDD1.n104 VSUBS 0.01078f
C884 VDD1.n105 VSUBS 0.011414f
C885 VDD1.n106 VSUBS 0.025479f
C886 VDD1.n107 VSUBS 0.025479f
C887 VDD1.n108 VSUBS 0.011414f
C888 VDD1.n109 VSUBS 0.01078f
C889 VDD1.n110 VSUBS 0.020061f
C890 VDD1.n111 VSUBS 0.020061f
C891 VDD1.n112 VSUBS 0.01078f
C892 VDD1.n113 VSUBS 0.011414f
C893 VDD1.n114 VSUBS 0.025479f
C894 VDD1.n115 VSUBS 0.025479f
C895 VDD1.n116 VSUBS 0.011414f
C896 VDD1.n117 VSUBS 0.01078f
C897 VDD1.n118 VSUBS 0.020061f
C898 VDD1.n119 VSUBS 0.020061f
C899 VDD1.n120 VSUBS 0.01078f
C900 VDD1.n121 VSUBS 0.01078f
C901 VDD1.n122 VSUBS 0.011414f
C902 VDD1.n123 VSUBS 0.025479f
C903 VDD1.n124 VSUBS 0.025479f
C904 VDD1.n125 VSUBS 0.025479f
C905 VDD1.n126 VSUBS 0.011097f
C906 VDD1.n127 VSUBS 0.01078f
C907 VDD1.n128 VSUBS 0.020061f
C908 VDD1.n129 VSUBS 0.020061f
C909 VDD1.n130 VSUBS 0.01078f
C910 VDD1.n131 VSUBS 0.011414f
C911 VDD1.n132 VSUBS 0.025479f
C912 VDD1.n133 VSUBS 0.025479f
C913 VDD1.n134 VSUBS 0.011414f
C914 VDD1.n135 VSUBS 0.01078f
C915 VDD1.n136 VSUBS 0.020061f
C916 VDD1.n137 VSUBS 0.020061f
C917 VDD1.n138 VSUBS 0.01078f
C918 VDD1.n139 VSUBS 0.011414f
C919 VDD1.n140 VSUBS 0.025479f
C920 VDD1.n141 VSUBS 0.025479f
C921 VDD1.n142 VSUBS 0.011414f
C922 VDD1.n143 VSUBS 0.01078f
C923 VDD1.n144 VSUBS 0.020061f
C924 VDD1.n145 VSUBS 0.020061f
C925 VDD1.n146 VSUBS 0.01078f
C926 VDD1.n147 VSUBS 0.011414f
C927 VDD1.n148 VSUBS 0.025479f
C928 VDD1.n149 VSUBS 0.064873f
C929 VDD1.n150 VSUBS 0.011414f
C930 VDD1.n151 VSUBS 0.01078f
C931 VDD1.n152 VSUBS 0.046369f
C932 VDD1.n153 VSUBS 0.618196f
C933 VTAIL.n0 VSUBS 0.032448f
C934 VTAIL.n1 VSUBS 0.028327f
C935 VTAIL.n2 VSUBS 0.015222f
C936 VTAIL.n3 VSUBS 0.035978f
C937 VTAIL.n4 VSUBS 0.016117f
C938 VTAIL.n5 VSUBS 0.028327f
C939 VTAIL.n6 VSUBS 0.015222f
C940 VTAIL.n7 VSUBS 0.035978f
C941 VTAIL.n8 VSUBS 0.016117f
C942 VTAIL.n9 VSUBS 0.028327f
C943 VTAIL.n10 VSUBS 0.015222f
C944 VTAIL.n11 VSUBS 0.035978f
C945 VTAIL.n12 VSUBS 0.016117f
C946 VTAIL.n13 VSUBS 0.028327f
C947 VTAIL.n14 VSUBS 0.015669f
C948 VTAIL.n15 VSUBS 0.035978f
C949 VTAIL.n16 VSUBS 0.016117f
C950 VTAIL.n17 VSUBS 0.028327f
C951 VTAIL.n18 VSUBS 0.015222f
C952 VTAIL.n19 VSUBS 0.035978f
C953 VTAIL.n20 VSUBS 0.016117f
C954 VTAIL.n21 VSUBS 0.028327f
C955 VTAIL.n22 VSUBS 0.015222f
C956 VTAIL.n23 VSUBS 0.026984f
C957 VTAIL.n24 VSUBS 0.027065f
C958 VTAIL.t2 VSUBS 0.077744f
C959 VTAIL.n25 VSUBS 0.25229f
C960 VTAIL.n26 VSUBS 1.67478f
C961 VTAIL.n27 VSUBS 0.015222f
C962 VTAIL.n28 VSUBS 0.016117f
C963 VTAIL.n29 VSUBS 0.035978f
C964 VTAIL.n30 VSUBS 0.035978f
C965 VTAIL.n31 VSUBS 0.016117f
C966 VTAIL.n32 VSUBS 0.015222f
C967 VTAIL.n33 VSUBS 0.028327f
C968 VTAIL.n34 VSUBS 0.028327f
C969 VTAIL.n35 VSUBS 0.015222f
C970 VTAIL.n36 VSUBS 0.016117f
C971 VTAIL.n37 VSUBS 0.035978f
C972 VTAIL.n38 VSUBS 0.035978f
C973 VTAIL.n39 VSUBS 0.016117f
C974 VTAIL.n40 VSUBS 0.015222f
C975 VTAIL.n41 VSUBS 0.028327f
C976 VTAIL.n42 VSUBS 0.028327f
C977 VTAIL.n43 VSUBS 0.015222f
C978 VTAIL.n44 VSUBS 0.015222f
C979 VTAIL.n45 VSUBS 0.016117f
C980 VTAIL.n46 VSUBS 0.035978f
C981 VTAIL.n47 VSUBS 0.035978f
C982 VTAIL.n48 VSUBS 0.035978f
C983 VTAIL.n49 VSUBS 0.015669f
C984 VTAIL.n50 VSUBS 0.015222f
C985 VTAIL.n51 VSUBS 0.028327f
C986 VTAIL.n52 VSUBS 0.028327f
C987 VTAIL.n53 VSUBS 0.015222f
C988 VTAIL.n54 VSUBS 0.016117f
C989 VTAIL.n55 VSUBS 0.035978f
C990 VTAIL.n56 VSUBS 0.035978f
C991 VTAIL.n57 VSUBS 0.016117f
C992 VTAIL.n58 VSUBS 0.015222f
C993 VTAIL.n59 VSUBS 0.028327f
C994 VTAIL.n60 VSUBS 0.028327f
C995 VTAIL.n61 VSUBS 0.015222f
C996 VTAIL.n62 VSUBS 0.016117f
C997 VTAIL.n63 VSUBS 0.035978f
C998 VTAIL.n64 VSUBS 0.035978f
C999 VTAIL.n65 VSUBS 0.016117f
C1000 VTAIL.n66 VSUBS 0.015222f
C1001 VTAIL.n67 VSUBS 0.028327f
C1002 VTAIL.n68 VSUBS 0.028327f
C1003 VTAIL.n69 VSUBS 0.015222f
C1004 VTAIL.n70 VSUBS 0.016117f
C1005 VTAIL.n71 VSUBS 0.035978f
C1006 VTAIL.n72 VSUBS 0.091604f
C1007 VTAIL.n73 VSUBS 0.016117f
C1008 VTAIL.n74 VSUBS 0.015222f
C1009 VTAIL.n75 VSUBS 0.065476f
C1010 VTAIL.n76 VSUBS 0.046267f
C1011 VTAIL.n77 VSUBS 1.86407f
C1012 VTAIL.n78 VSUBS 0.032448f
C1013 VTAIL.n79 VSUBS 0.028327f
C1014 VTAIL.n80 VSUBS 0.015222f
C1015 VTAIL.n81 VSUBS 0.035978f
C1016 VTAIL.n82 VSUBS 0.016117f
C1017 VTAIL.n83 VSUBS 0.028327f
C1018 VTAIL.n84 VSUBS 0.015222f
C1019 VTAIL.n85 VSUBS 0.035978f
C1020 VTAIL.n86 VSUBS 0.016117f
C1021 VTAIL.n87 VSUBS 0.028327f
C1022 VTAIL.n88 VSUBS 0.015222f
C1023 VTAIL.n89 VSUBS 0.035978f
C1024 VTAIL.n90 VSUBS 0.016117f
C1025 VTAIL.n91 VSUBS 0.028327f
C1026 VTAIL.n92 VSUBS 0.015669f
C1027 VTAIL.n93 VSUBS 0.035978f
C1028 VTAIL.n94 VSUBS 0.015222f
C1029 VTAIL.n95 VSUBS 0.016117f
C1030 VTAIL.n96 VSUBS 0.028327f
C1031 VTAIL.n97 VSUBS 0.015222f
C1032 VTAIL.n98 VSUBS 0.035978f
C1033 VTAIL.n99 VSUBS 0.016117f
C1034 VTAIL.n100 VSUBS 0.028327f
C1035 VTAIL.n101 VSUBS 0.015222f
C1036 VTAIL.n102 VSUBS 0.026984f
C1037 VTAIL.n103 VSUBS 0.027065f
C1038 VTAIL.t1 VSUBS 0.077744f
C1039 VTAIL.n104 VSUBS 0.25229f
C1040 VTAIL.n105 VSUBS 1.67478f
C1041 VTAIL.n106 VSUBS 0.015222f
C1042 VTAIL.n107 VSUBS 0.016117f
C1043 VTAIL.n108 VSUBS 0.035978f
C1044 VTAIL.n109 VSUBS 0.035978f
C1045 VTAIL.n110 VSUBS 0.016117f
C1046 VTAIL.n111 VSUBS 0.015222f
C1047 VTAIL.n112 VSUBS 0.028327f
C1048 VTAIL.n113 VSUBS 0.028327f
C1049 VTAIL.n114 VSUBS 0.015222f
C1050 VTAIL.n115 VSUBS 0.016117f
C1051 VTAIL.n116 VSUBS 0.035978f
C1052 VTAIL.n117 VSUBS 0.035978f
C1053 VTAIL.n118 VSUBS 0.016117f
C1054 VTAIL.n119 VSUBS 0.015222f
C1055 VTAIL.n120 VSUBS 0.028327f
C1056 VTAIL.n121 VSUBS 0.028327f
C1057 VTAIL.n122 VSUBS 0.015222f
C1058 VTAIL.n123 VSUBS 0.016117f
C1059 VTAIL.n124 VSUBS 0.035978f
C1060 VTAIL.n125 VSUBS 0.035978f
C1061 VTAIL.n126 VSUBS 0.035978f
C1062 VTAIL.n127 VSUBS 0.015669f
C1063 VTAIL.n128 VSUBS 0.015222f
C1064 VTAIL.n129 VSUBS 0.028327f
C1065 VTAIL.n130 VSUBS 0.028327f
C1066 VTAIL.n131 VSUBS 0.015222f
C1067 VTAIL.n132 VSUBS 0.016117f
C1068 VTAIL.n133 VSUBS 0.035978f
C1069 VTAIL.n134 VSUBS 0.035978f
C1070 VTAIL.n135 VSUBS 0.016117f
C1071 VTAIL.n136 VSUBS 0.015222f
C1072 VTAIL.n137 VSUBS 0.028327f
C1073 VTAIL.n138 VSUBS 0.028327f
C1074 VTAIL.n139 VSUBS 0.015222f
C1075 VTAIL.n140 VSUBS 0.016117f
C1076 VTAIL.n141 VSUBS 0.035978f
C1077 VTAIL.n142 VSUBS 0.035978f
C1078 VTAIL.n143 VSUBS 0.016117f
C1079 VTAIL.n144 VSUBS 0.015222f
C1080 VTAIL.n145 VSUBS 0.028327f
C1081 VTAIL.n146 VSUBS 0.028327f
C1082 VTAIL.n147 VSUBS 0.015222f
C1083 VTAIL.n148 VSUBS 0.016117f
C1084 VTAIL.n149 VSUBS 0.035978f
C1085 VTAIL.n150 VSUBS 0.091604f
C1086 VTAIL.n151 VSUBS 0.016117f
C1087 VTAIL.n152 VSUBS 0.015222f
C1088 VTAIL.n153 VSUBS 0.065476f
C1089 VTAIL.n154 VSUBS 0.046267f
C1090 VTAIL.n155 VSUBS 1.89023f
C1091 VTAIL.n156 VSUBS 0.032448f
C1092 VTAIL.n157 VSUBS 0.028327f
C1093 VTAIL.n158 VSUBS 0.015222f
C1094 VTAIL.n159 VSUBS 0.035978f
C1095 VTAIL.n160 VSUBS 0.016117f
C1096 VTAIL.n161 VSUBS 0.028327f
C1097 VTAIL.n162 VSUBS 0.015222f
C1098 VTAIL.n163 VSUBS 0.035978f
C1099 VTAIL.n164 VSUBS 0.016117f
C1100 VTAIL.n165 VSUBS 0.028327f
C1101 VTAIL.n166 VSUBS 0.015222f
C1102 VTAIL.n167 VSUBS 0.035978f
C1103 VTAIL.n168 VSUBS 0.016117f
C1104 VTAIL.n169 VSUBS 0.028327f
C1105 VTAIL.n170 VSUBS 0.015669f
C1106 VTAIL.n171 VSUBS 0.035978f
C1107 VTAIL.n172 VSUBS 0.015222f
C1108 VTAIL.n173 VSUBS 0.016117f
C1109 VTAIL.n174 VSUBS 0.028327f
C1110 VTAIL.n175 VSUBS 0.015222f
C1111 VTAIL.n176 VSUBS 0.035978f
C1112 VTAIL.n177 VSUBS 0.016117f
C1113 VTAIL.n178 VSUBS 0.028327f
C1114 VTAIL.n179 VSUBS 0.015222f
C1115 VTAIL.n180 VSUBS 0.026984f
C1116 VTAIL.n181 VSUBS 0.027065f
C1117 VTAIL.t3 VSUBS 0.077744f
C1118 VTAIL.n182 VSUBS 0.25229f
C1119 VTAIL.n183 VSUBS 1.67478f
C1120 VTAIL.n184 VSUBS 0.015222f
C1121 VTAIL.n185 VSUBS 0.016117f
C1122 VTAIL.n186 VSUBS 0.035978f
C1123 VTAIL.n187 VSUBS 0.035978f
C1124 VTAIL.n188 VSUBS 0.016117f
C1125 VTAIL.n189 VSUBS 0.015222f
C1126 VTAIL.n190 VSUBS 0.028327f
C1127 VTAIL.n191 VSUBS 0.028327f
C1128 VTAIL.n192 VSUBS 0.015222f
C1129 VTAIL.n193 VSUBS 0.016117f
C1130 VTAIL.n194 VSUBS 0.035978f
C1131 VTAIL.n195 VSUBS 0.035978f
C1132 VTAIL.n196 VSUBS 0.016117f
C1133 VTAIL.n197 VSUBS 0.015222f
C1134 VTAIL.n198 VSUBS 0.028327f
C1135 VTAIL.n199 VSUBS 0.028327f
C1136 VTAIL.n200 VSUBS 0.015222f
C1137 VTAIL.n201 VSUBS 0.016117f
C1138 VTAIL.n202 VSUBS 0.035978f
C1139 VTAIL.n203 VSUBS 0.035978f
C1140 VTAIL.n204 VSUBS 0.035978f
C1141 VTAIL.n205 VSUBS 0.015669f
C1142 VTAIL.n206 VSUBS 0.015222f
C1143 VTAIL.n207 VSUBS 0.028327f
C1144 VTAIL.n208 VSUBS 0.028327f
C1145 VTAIL.n209 VSUBS 0.015222f
C1146 VTAIL.n210 VSUBS 0.016117f
C1147 VTAIL.n211 VSUBS 0.035978f
C1148 VTAIL.n212 VSUBS 0.035978f
C1149 VTAIL.n213 VSUBS 0.016117f
C1150 VTAIL.n214 VSUBS 0.015222f
C1151 VTAIL.n215 VSUBS 0.028327f
C1152 VTAIL.n216 VSUBS 0.028327f
C1153 VTAIL.n217 VSUBS 0.015222f
C1154 VTAIL.n218 VSUBS 0.016117f
C1155 VTAIL.n219 VSUBS 0.035978f
C1156 VTAIL.n220 VSUBS 0.035978f
C1157 VTAIL.n221 VSUBS 0.016117f
C1158 VTAIL.n222 VSUBS 0.015222f
C1159 VTAIL.n223 VSUBS 0.028327f
C1160 VTAIL.n224 VSUBS 0.028327f
C1161 VTAIL.n225 VSUBS 0.015222f
C1162 VTAIL.n226 VSUBS 0.016117f
C1163 VTAIL.n227 VSUBS 0.035978f
C1164 VTAIL.n228 VSUBS 0.091604f
C1165 VTAIL.n229 VSUBS 0.016117f
C1166 VTAIL.n230 VSUBS 0.015222f
C1167 VTAIL.n231 VSUBS 0.065476f
C1168 VTAIL.n232 VSUBS 0.046267f
C1169 VTAIL.n233 VSUBS 1.76434f
C1170 VTAIL.n234 VSUBS 0.032448f
C1171 VTAIL.n235 VSUBS 0.028327f
C1172 VTAIL.n236 VSUBS 0.015222f
C1173 VTAIL.n237 VSUBS 0.035978f
C1174 VTAIL.n238 VSUBS 0.016117f
C1175 VTAIL.n239 VSUBS 0.028327f
C1176 VTAIL.n240 VSUBS 0.015222f
C1177 VTAIL.n241 VSUBS 0.035978f
C1178 VTAIL.n242 VSUBS 0.016117f
C1179 VTAIL.n243 VSUBS 0.028327f
C1180 VTAIL.n244 VSUBS 0.015222f
C1181 VTAIL.n245 VSUBS 0.035978f
C1182 VTAIL.n246 VSUBS 0.016117f
C1183 VTAIL.n247 VSUBS 0.028327f
C1184 VTAIL.n248 VSUBS 0.015669f
C1185 VTAIL.n249 VSUBS 0.035978f
C1186 VTAIL.n250 VSUBS 0.016117f
C1187 VTAIL.n251 VSUBS 0.028327f
C1188 VTAIL.n252 VSUBS 0.015222f
C1189 VTAIL.n253 VSUBS 0.035978f
C1190 VTAIL.n254 VSUBS 0.016117f
C1191 VTAIL.n255 VSUBS 0.028327f
C1192 VTAIL.n256 VSUBS 0.015222f
C1193 VTAIL.n257 VSUBS 0.026984f
C1194 VTAIL.n258 VSUBS 0.027065f
C1195 VTAIL.t0 VSUBS 0.077744f
C1196 VTAIL.n259 VSUBS 0.25229f
C1197 VTAIL.n260 VSUBS 1.67478f
C1198 VTAIL.n261 VSUBS 0.015222f
C1199 VTAIL.n262 VSUBS 0.016117f
C1200 VTAIL.n263 VSUBS 0.035978f
C1201 VTAIL.n264 VSUBS 0.035978f
C1202 VTAIL.n265 VSUBS 0.016117f
C1203 VTAIL.n266 VSUBS 0.015222f
C1204 VTAIL.n267 VSUBS 0.028327f
C1205 VTAIL.n268 VSUBS 0.028327f
C1206 VTAIL.n269 VSUBS 0.015222f
C1207 VTAIL.n270 VSUBS 0.016117f
C1208 VTAIL.n271 VSUBS 0.035978f
C1209 VTAIL.n272 VSUBS 0.035978f
C1210 VTAIL.n273 VSUBS 0.016117f
C1211 VTAIL.n274 VSUBS 0.015222f
C1212 VTAIL.n275 VSUBS 0.028327f
C1213 VTAIL.n276 VSUBS 0.028327f
C1214 VTAIL.n277 VSUBS 0.015222f
C1215 VTAIL.n278 VSUBS 0.015222f
C1216 VTAIL.n279 VSUBS 0.016117f
C1217 VTAIL.n280 VSUBS 0.035978f
C1218 VTAIL.n281 VSUBS 0.035978f
C1219 VTAIL.n282 VSUBS 0.035978f
C1220 VTAIL.n283 VSUBS 0.015669f
C1221 VTAIL.n284 VSUBS 0.015222f
C1222 VTAIL.n285 VSUBS 0.028327f
C1223 VTAIL.n286 VSUBS 0.028327f
C1224 VTAIL.n287 VSUBS 0.015222f
C1225 VTAIL.n288 VSUBS 0.016117f
C1226 VTAIL.n289 VSUBS 0.035978f
C1227 VTAIL.n290 VSUBS 0.035978f
C1228 VTAIL.n291 VSUBS 0.016117f
C1229 VTAIL.n292 VSUBS 0.015222f
C1230 VTAIL.n293 VSUBS 0.028327f
C1231 VTAIL.n294 VSUBS 0.028327f
C1232 VTAIL.n295 VSUBS 0.015222f
C1233 VTAIL.n296 VSUBS 0.016117f
C1234 VTAIL.n297 VSUBS 0.035978f
C1235 VTAIL.n298 VSUBS 0.035978f
C1236 VTAIL.n299 VSUBS 0.016117f
C1237 VTAIL.n300 VSUBS 0.015222f
C1238 VTAIL.n301 VSUBS 0.028327f
C1239 VTAIL.n302 VSUBS 0.028327f
C1240 VTAIL.n303 VSUBS 0.015222f
C1241 VTAIL.n304 VSUBS 0.016117f
C1242 VTAIL.n305 VSUBS 0.035978f
C1243 VTAIL.n306 VSUBS 0.091604f
C1244 VTAIL.n307 VSUBS 0.016117f
C1245 VTAIL.n308 VSUBS 0.015222f
C1246 VTAIL.n309 VSUBS 0.065476f
C1247 VTAIL.n310 VSUBS 0.046267f
C1248 VTAIL.n311 VSUBS 1.68467f
C1249 VP.t1 VSUBS 3.45227f
C1250 VP.t0 VSUBS 3.11904f
C1251 VP.n0 VSUBS 6.27857f
.ends

