* NGSPICE file created from diff_pair_sample_1218.ext - technology: sky130A

.subckt diff_pair_sample_1218 VTAIL VN VP B VDD2 VDD1
X0 B.t11 B.t9 B.t10 w_n2866_n3224# sky130_fd_pr__pfet_01v8 ad=4.3992 pd=23.34 as=0 ps=0 w=11.28 l=2.83
X1 VTAIL.t5 VN.t0 VDD2.t0 w_n2866_n3224# sky130_fd_pr__pfet_01v8 ad=4.3992 pd=23.34 as=1.8612 ps=11.61 w=11.28 l=2.83
X2 VDD1.t3 VP.t0 VTAIL.t0 w_n2866_n3224# sky130_fd_pr__pfet_01v8 ad=1.8612 pd=11.61 as=4.3992 ps=23.34 w=11.28 l=2.83
X3 B.t8 B.t6 B.t7 w_n2866_n3224# sky130_fd_pr__pfet_01v8 ad=4.3992 pd=23.34 as=0 ps=0 w=11.28 l=2.83
X4 VDD2.t1 VN.t1 VTAIL.t4 w_n2866_n3224# sky130_fd_pr__pfet_01v8 ad=1.8612 pd=11.61 as=4.3992 ps=23.34 w=11.28 l=2.83
X5 VTAIL.t7 VP.t1 VDD1.t2 w_n2866_n3224# sky130_fd_pr__pfet_01v8 ad=4.3992 pd=23.34 as=1.8612 ps=11.61 w=11.28 l=2.83
X6 VTAIL.t3 VN.t2 VDD2.t3 w_n2866_n3224# sky130_fd_pr__pfet_01v8 ad=4.3992 pd=23.34 as=1.8612 ps=11.61 w=11.28 l=2.83
X7 B.t5 B.t3 B.t4 w_n2866_n3224# sky130_fd_pr__pfet_01v8 ad=4.3992 pd=23.34 as=0 ps=0 w=11.28 l=2.83
X8 VDD1.t1 VP.t2 VTAIL.t6 w_n2866_n3224# sky130_fd_pr__pfet_01v8 ad=1.8612 pd=11.61 as=4.3992 ps=23.34 w=11.28 l=2.83
X9 B.t2 B.t0 B.t1 w_n2866_n3224# sky130_fd_pr__pfet_01v8 ad=4.3992 pd=23.34 as=0 ps=0 w=11.28 l=2.83
X10 VDD2.t2 VN.t3 VTAIL.t2 w_n2866_n3224# sky130_fd_pr__pfet_01v8 ad=1.8612 pd=11.61 as=4.3992 ps=23.34 w=11.28 l=2.83
X11 VTAIL.t1 VP.t3 VDD1.t0 w_n2866_n3224# sky130_fd_pr__pfet_01v8 ad=4.3992 pd=23.34 as=1.8612 ps=11.61 w=11.28 l=2.83
R0 B.n470 B.n469 585
R1 B.n471 B.n68 585
R2 B.n473 B.n472 585
R3 B.n474 B.n67 585
R4 B.n476 B.n475 585
R5 B.n477 B.n66 585
R6 B.n479 B.n478 585
R7 B.n480 B.n65 585
R8 B.n482 B.n481 585
R9 B.n483 B.n64 585
R10 B.n485 B.n484 585
R11 B.n486 B.n63 585
R12 B.n488 B.n487 585
R13 B.n489 B.n62 585
R14 B.n491 B.n490 585
R15 B.n492 B.n61 585
R16 B.n494 B.n493 585
R17 B.n495 B.n60 585
R18 B.n497 B.n496 585
R19 B.n498 B.n59 585
R20 B.n500 B.n499 585
R21 B.n501 B.n58 585
R22 B.n503 B.n502 585
R23 B.n504 B.n57 585
R24 B.n506 B.n505 585
R25 B.n507 B.n56 585
R26 B.n509 B.n508 585
R27 B.n510 B.n55 585
R28 B.n512 B.n511 585
R29 B.n513 B.n54 585
R30 B.n515 B.n514 585
R31 B.n516 B.n53 585
R32 B.n518 B.n517 585
R33 B.n519 B.n52 585
R34 B.n521 B.n520 585
R35 B.n522 B.n51 585
R36 B.n524 B.n523 585
R37 B.n525 B.n50 585
R38 B.n527 B.n526 585
R39 B.n528 B.n47 585
R40 B.n531 B.n530 585
R41 B.n532 B.n46 585
R42 B.n534 B.n533 585
R43 B.n535 B.n45 585
R44 B.n537 B.n536 585
R45 B.n538 B.n44 585
R46 B.n540 B.n539 585
R47 B.n541 B.n43 585
R48 B.n543 B.n542 585
R49 B.n545 B.n544 585
R50 B.n546 B.n39 585
R51 B.n548 B.n547 585
R52 B.n549 B.n38 585
R53 B.n551 B.n550 585
R54 B.n552 B.n37 585
R55 B.n554 B.n553 585
R56 B.n555 B.n36 585
R57 B.n557 B.n556 585
R58 B.n558 B.n35 585
R59 B.n560 B.n559 585
R60 B.n561 B.n34 585
R61 B.n563 B.n562 585
R62 B.n564 B.n33 585
R63 B.n566 B.n565 585
R64 B.n567 B.n32 585
R65 B.n569 B.n568 585
R66 B.n570 B.n31 585
R67 B.n572 B.n571 585
R68 B.n573 B.n30 585
R69 B.n575 B.n574 585
R70 B.n576 B.n29 585
R71 B.n578 B.n577 585
R72 B.n579 B.n28 585
R73 B.n581 B.n580 585
R74 B.n582 B.n27 585
R75 B.n584 B.n583 585
R76 B.n585 B.n26 585
R77 B.n587 B.n586 585
R78 B.n588 B.n25 585
R79 B.n590 B.n589 585
R80 B.n591 B.n24 585
R81 B.n593 B.n592 585
R82 B.n594 B.n23 585
R83 B.n596 B.n595 585
R84 B.n597 B.n22 585
R85 B.n599 B.n598 585
R86 B.n600 B.n21 585
R87 B.n602 B.n601 585
R88 B.n603 B.n20 585
R89 B.n468 B.n69 585
R90 B.n467 B.n466 585
R91 B.n465 B.n70 585
R92 B.n464 B.n463 585
R93 B.n462 B.n71 585
R94 B.n461 B.n460 585
R95 B.n459 B.n72 585
R96 B.n458 B.n457 585
R97 B.n456 B.n73 585
R98 B.n455 B.n454 585
R99 B.n453 B.n74 585
R100 B.n452 B.n451 585
R101 B.n450 B.n75 585
R102 B.n449 B.n448 585
R103 B.n447 B.n76 585
R104 B.n446 B.n445 585
R105 B.n444 B.n77 585
R106 B.n443 B.n442 585
R107 B.n441 B.n78 585
R108 B.n440 B.n439 585
R109 B.n438 B.n79 585
R110 B.n437 B.n436 585
R111 B.n435 B.n80 585
R112 B.n434 B.n433 585
R113 B.n432 B.n81 585
R114 B.n431 B.n430 585
R115 B.n429 B.n82 585
R116 B.n428 B.n427 585
R117 B.n426 B.n83 585
R118 B.n425 B.n424 585
R119 B.n423 B.n84 585
R120 B.n422 B.n421 585
R121 B.n420 B.n85 585
R122 B.n419 B.n418 585
R123 B.n417 B.n86 585
R124 B.n416 B.n415 585
R125 B.n414 B.n87 585
R126 B.n413 B.n412 585
R127 B.n411 B.n88 585
R128 B.n410 B.n409 585
R129 B.n408 B.n89 585
R130 B.n407 B.n406 585
R131 B.n405 B.n90 585
R132 B.n404 B.n403 585
R133 B.n402 B.n91 585
R134 B.n401 B.n400 585
R135 B.n399 B.n92 585
R136 B.n398 B.n397 585
R137 B.n396 B.n93 585
R138 B.n395 B.n394 585
R139 B.n393 B.n94 585
R140 B.n392 B.n391 585
R141 B.n390 B.n95 585
R142 B.n389 B.n388 585
R143 B.n387 B.n96 585
R144 B.n386 B.n385 585
R145 B.n384 B.n97 585
R146 B.n383 B.n382 585
R147 B.n381 B.n98 585
R148 B.n380 B.n379 585
R149 B.n378 B.n99 585
R150 B.n377 B.n376 585
R151 B.n375 B.n100 585
R152 B.n374 B.n373 585
R153 B.n372 B.n101 585
R154 B.n371 B.n370 585
R155 B.n369 B.n102 585
R156 B.n368 B.n367 585
R157 B.n366 B.n103 585
R158 B.n365 B.n364 585
R159 B.n363 B.n104 585
R160 B.n362 B.n361 585
R161 B.n360 B.n105 585
R162 B.n225 B.n154 585
R163 B.n227 B.n226 585
R164 B.n228 B.n153 585
R165 B.n230 B.n229 585
R166 B.n231 B.n152 585
R167 B.n233 B.n232 585
R168 B.n234 B.n151 585
R169 B.n236 B.n235 585
R170 B.n237 B.n150 585
R171 B.n239 B.n238 585
R172 B.n240 B.n149 585
R173 B.n242 B.n241 585
R174 B.n243 B.n148 585
R175 B.n245 B.n244 585
R176 B.n246 B.n147 585
R177 B.n248 B.n247 585
R178 B.n249 B.n146 585
R179 B.n251 B.n250 585
R180 B.n252 B.n145 585
R181 B.n254 B.n253 585
R182 B.n255 B.n144 585
R183 B.n257 B.n256 585
R184 B.n258 B.n143 585
R185 B.n260 B.n259 585
R186 B.n261 B.n142 585
R187 B.n263 B.n262 585
R188 B.n264 B.n141 585
R189 B.n266 B.n265 585
R190 B.n267 B.n140 585
R191 B.n269 B.n268 585
R192 B.n270 B.n139 585
R193 B.n272 B.n271 585
R194 B.n273 B.n138 585
R195 B.n275 B.n274 585
R196 B.n276 B.n137 585
R197 B.n278 B.n277 585
R198 B.n279 B.n136 585
R199 B.n281 B.n280 585
R200 B.n282 B.n135 585
R201 B.n284 B.n283 585
R202 B.n286 B.n285 585
R203 B.n287 B.n131 585
R204 B.n289 B.n288 585
R205 B.n290 B.n130 585
R206 B.n292 B.n291 585
R207 B.n293 B.n129 585
R208 B.n295 B.n294 585
R209 B.n296 B.n128 585
R210 B.n298 B.n297 585
R211 B.n300 B.n125 585
R212 B.n302 B.n301 585
R213 B.n303 B.n124 585
R214 B.n305 B.n304 585
R215 B.n306 B.n123 585
R216 B.n308 B.n307 585
R217 B.n309 B.n122 585
R218 B.n311 B.n310 585
R219 B.n312 B.n121 585
R220 B.n314 B.n313 585
R221 B.n315 B.n120 585
R222 B.n317 B.n316 585
R223 B.n318 B.n119 585
R224 B.n320 B.n319 585
R225 B.n321 B.n118 585
R226 B.n323 B.n322 585
R227 B.n324 B.n117 585
R228 B.n326 B.n325 585
R229 B.n327 B.n116 585
R230 B.n329 B.n328 585
R231 B.n330 B.n115 585
R232 B.n332 B.n331 585
R233 B.n333 B.n114 585
R234 B.n335 B.n334 585
R235 B.n336 B.n113 585
R236 B.n338 B.n337 585
R237 B.n339 B.n112 585
R238 B.n341 B.n340 585
R239 B.n342 B.n111 585
R240 B.n344 B.n343 585
R241 B.n345 B.n110 585
R242 B.n347 B.n346 585
R243 B.n348 B.n109 585
R244 B.n350 B.n349 585
R245 B.n351 B.n108 585
R246 B.n353 B.n352 585
R247 B.n354 B.n107 585
R248 B.n356 B.n355 585
R249 B.n357 B.n106 585
R250 B.n359 B.n358 585
R251 B.n224 B.n223 585
R252 B.n222 B.n155 585
R253 B.n221 B.n220 585
R254 B.n219 B.n156 585
R255 B.n218 B.n217 585
R256 B.n216 B.n157 585
R257 B.n215 B.n214 585
R258 B.n213 B.n158 585
R259 B.n212 B.n211 585
R260 B.n210 B.n159 585
R261 B.n209 B.n208 585
R262 B.n207 B.n160 585
R263 B.n206 B.n205 585
R264 B.n204 B.n161 585
R265 B.n203 B.n202 585
R266 B.n201 B.n162 585
R267 B.n200 B.n199 585
R268 B.n198 B.n163 585
R269 B.n197 B.n196 585
R270 B.n195 B.n164 585
R271 B.n194 B.n193 585
R272 B.n192 B.n165 585
R273 B.n191 B.n190 585
R274 B.n189 B.n166 585
R275 B.n188 B.n187 585
R276 B.n186 B.n167 585
R277 B.n185 B.n184 585
R278 B.n183 B.n168 585
R279 B.n182 B.n181 585
R280 B.n180 B.n169 585
R281 B.n179 B.n178 585
R282 B.n177 B.n170 585
R283 B.n176 B.n175 585
R284 B.n174 B.n171 585
R285 B.n173 B.n172 585
R286 B.n2 B.n0 585
R287 B.n657 B.n1 585
R288 B.n656 B.n655 585
R289 B.n654 B.n3 585
R290 B.n653 B.n652 585
R291 B.n651 B.n4 585
R292 B.n650 B.n649 585
R293 B.n648 B.n5 585
R294 B.n647 B.n646 585
R295 B.n645 B.n6 585
R296 B.n644 B.n643 585
R297 B.n642 B.n7 585
R298 B.n641 B.n640 585
R299 B.n639 B.n8 585
R300 B.n638 B.n637 585
R301 B.n636 B.n9 585
R302 B.n635 B.n634 585
R303 B.n633 B.n10 585
R304 B.n632 B.n631 585
R305 B.n630 B.n11 585
R306 B.n629 B.n628 585
R307 B.n627 B.n12 585
R308 B.n626 B.n625 585
R309 B.n624 B.n13 585
R310 B.n623 B.n622 585
R311 B.n621 B.n14 585
R312 B.n620 B.n619 585
R313 B.n618 B.n15 585
R314 B.n617 B.n616 585
R315 B.n615 B.n16 585
R316 B.n614 B.n613 585
R317 B.n612 B.n17 585
R318 B.n611 B.n610 585
R319 B.n609 B.n18 585
R320 B.n608 B.n607 585
R321 B.n606 B.n19 585
R322 B.n605 B.n604 585
R323 B.n659 B.n658 585
R324 B.n225 B.n224 463.671
R325 B.n604 B.n603 463.671
R326 B.n358 B.n105 463.671
R327 B.n470 B.n69 463.671
R328 B.n126 B.t11 423.793
R329 B.n48 B.t4 423.793
R330 B.n132 B.t2 423.793
R331 B.n40 B.t7 423.793
R332 B.n127 B.t10 362.509
R333 B.n49 B.t5 362.509
R334 B.n133 B.t1 362.509
R335 B.n41 B.t8 362.509
R336 B.n126 B.t9 304.43
R337 B.n132 B.t0 304.43
R338 B.n40 B.t6 304.43
R339 B.n48 B.t3 304.43
R340 B.n224 B.n155 163.367
R341 B.n220 B.n155 163.367
R342 B.n220 B.n219 163.367
R343 B.n219 B.n218 163.367
R344 B.n218 B.n157 163.367
R345 B.n214 B.n157 163.367
R346 B.n214 B.n213 163.367
R347 B.n213 B.n212 163.367
R348 B.n212 B.n159 163.367
R349 B.n208 B.n159 163.367
R350 B.n208 B.n207 163.367
R351 B.n207 B.n206 163.367
R352 B.n206 B.n161 163.367
R353 B.n202 B.n161 163.367
R354 B.n202 B.n201 163.367
R355 B.n201 B.n200 163.367
R356 B.n200 B.n163 163.367
R357 B.n196 B.n163 163.367
R358 B.n196 B.n195 163.367
R359 B.n195 B.n194 163.367
R360 B.n194 B.n165 163.367
R361 B.n190 B.n165 163.367
R362 B.n190 B.n189 163.367
R363 B.n189 B.n188 163.367
R364 B.n188 B.n167 163.367
R365 B.n184 B.n167 163.367
R366 B.n184 B.n183 163.367
R367 B.n183 B.n182 163.367
R368 B.n182 B.n169 163.367
R369 B.n178 B.n169 163.367
R370 B.n178 B.n177 163.367
R371 B.n177 B.n176 163.367
R372 B.n176 B.n171 163.367
R373 B.n172 B.n171 163.367
R374 B.n172 B.n2 163.367
R375 B.n658 B.n2 163.367
R376 B.n658 B.n657 163.367
R377 B.n657 B.n656 163.367
R378 B.n656 B.n3 163.367
R379 B.n652 B.n3 163.367
R380 B.n652 B.n651 163.367
R381 B.n651 B.n650 163.367
R382 B.n650 B.n5 163.367
R383 B.n646 B.n5 163.367
R384 B.n646 B.n645 163.367
R385 B.n645 B.n644 163.367
R386 B.n644 B.n7 163.367
R387 B.n640 B.n7 163.367
R388 B.n640 B.n639 163.367
R389 B.n639 B.n638 163.367
R390 B.n638 B.n9 163.367
R391 B.n634 B.n9 163.367
R392 B.n634 B.n633 163.367
R393 B.n633 B.n632 163.367
R394 B.n632 B.n11 163.367
R395 B.n628 B.n11 163.367
R396 B.n628 B.n627 163.367
R397 B.n627 B.n626 163.367
R398 B.n626 B.n13 163.367
R399 B.n622 B.n13 163.367
R400 B.n622 B.n621 163.367
R401 B.n621 B.n620 163.367
R402 B.n620 B.n15 163.367
R403 B.n616 B.n15 163.367
R404 B.n616 B.n615 163.367
R405 B.n615 B.n614 163.367
R406 B.n614 B.n17 163.367
R407 B.n610 B.n17 163.367
R408 B.n610 B.n609 163.367
R409 B.n609 B.n608 163.367
R410 B.n608 B.n19 163.367
R411 B.n604 B.n19 163.367
R412 B.n226 B.n225 163.367
R413 B.n226 B.n153 163.367
R414 B.n230 B.n153 163.367
R415 B.n231 B.n230 163.367
R416 B.n232 B.n231 163.367
R417 B.n232 B.n151 163.367
R418 B.n236 B.n151 163.367
R419 B.n237 B.n236 163.367
R420 B.n238 B.n237 163.367
R421 B.n238 B.n149 163.367
R422 B.n242 B.n149 163.367
R423 B.n243 B.n242 163.367
R424 B.n244 B.n243 163.367
R425 B.n244 B.n147 163.367
R426 B.n248 B.n147 163.367
R427 B.n249 B.n248 163.367
R428 B.n250 B.n249 163.367
R429 B.n250 B.n145 163.367
R430 B.n254 B.n145 163.367
R431 B.n255 B.n254 163.367
R432 B.n256 B.n255 163.367
R433 B.n256 B.n143 163.367
R434 B.n260 B.n143 163.367
R435 B.n261 B.n260 163.367
R436 B.n262 B.n261 163.367
R437 B.n262 B.n141 163.367
R438 B.n266 B.n141 163.367
R439 B.n267 B.n266 163.367
R440 B.n268 B.n267 163.367
R441 B.n268 B.n139 163.367
R442 B.n272 B.n139 163.367
R443 B.n273 B.n272 163.367
R444 B.n274 B.n273 163.367
R445 B.n274 B.n137 163.367
R446 B.n278 B.n137 163.367
R447 B.n279 B.n278 163.367
R448 B.n280 B.n279 163.367
R449 B.n280 B.n135 163.367
R450 B.n284 B.n135 163.367
R451 B.n285 B.n284 163.367
R452 B.n285 B.n131 163.367
R453 B.n289 B.n131 163.367
R454 B.n290 B.n289 163.367
R455 B.n291 B.n290 163.367
R456 B.n291 B.n129 163.367
R457 B.n295 B.n129 163.367
R458 B.n296 B.n295 163.367
R459 B.n297 B.n296 163.367
R460 B.n297 B.n125 163.367
R461 B.n302 B.n125 163.367
R462 B.n303 B.n302 163.367
R463 B.n304 B.n303 163.367
R464 B.n304 B.n123 163.367
R465 B.n308 B.n123 163.367
R466 B.n309 B.n308 163.367
R467 B.n310 B.n309 163.367
R468 B.n310 B.n121 163.367
R469 B.n314 B.n121 163.367
R470 B.n315 B.n314 163.367
R471 B.n316 B.n315 163.367
R472 B.n316 B.n119 163.367
R473 B.n320 B.n119 163.367
R474 B.n321 B.n320 163.367
R475 B.n322 B.n321 163.367
R476 B.n322 B.n117 163.367
R477 B.n326 B.n117 163.367
R478 B.n327 B.n326 163.367
R479 B.n328 B.n327 163.367
R480 B.n328 B.n115 163.367
R481 B.n332 B.n115 163.367
R482 B.n333 B.n332 163.367
R483 B.n334 B.n333 163.367
R484 B.n334 B.n113 163.367
R485 B.n338 B.n113 163.367
R486 B.n339 B.n338 163.367
R487 B.n340 B.n339 163.367
R488 B.n340 B.n111 163.367
R489 B.n344 B.n111 163.367
R490 B.n345 B.n344 163.367
R491 B.n346 B.n345 163.367
R492 B.n346 B.n109 163.367
R493 B.n350 B.n109 163.367
R494 B.n351 B.n350 163.367
R495 B.n352 B.n351 163.367
R496 B.n352 B.n107 163.367
R497 B.n356 B.n107 163.367
R498 B.n357 B.n356 163.367
R499 B.n358 B.n357 163.367
R500 B.n362 B.n105 163.367
R501 B.n363 B.n362 163.367
R502 B.n364 B.n363 163.367
R503 B.n364 B.n103 163.367
R504 B.n368 B.n103 163.367
R505 B.n369 B.n368 163.367
R506 B.n370 B.n369 163.367
R507 B.n370 B.n101 163.367
R508 B.n374 B.n101 163.367
R509 B.n375 B.n374 163.367
R510 B.n376 B.n375 163.367
R511 B.n376 B.n99 163.367
R512 B.n380 B.n99 163.367
R513 B.n381 B.n380 163.367
R514 B.n382 B.n381 163.367
R515 B.n382 B.n97 163.367
R516 B.n386 B.n97 163.367
R517 B.n387 B.n386 163.367
R518 B.n388 B.n387 163.367
R519 B.n388 B.n95 163.367
R520 B.n392 B.n95 163.367
R521 B.n393 B.n392 163.367
R522 B.n394 B.n393 163.367
R523 B.n394 B.n93 163.367
R524 B.n398 B.n93 163.367
R525 B.n399 B.n398 163.367
R526 B.n400 B.n399 163.367
R527 B.n400 B.n91 163.367
R528 B.n404 B.n91 163.367
R529 B.n405 B.n404 163.367
R530 B.n406 B.n405 163.367
R531 B.n406 B.n89 163.367
R532 B.n410 B.n89 163.367
R533 B.n411 B.n410 163.367
R534 B.n412 B.n411 163.367
R535 B.n412 B.n87 163.367
R536 B.n416 B.n87 163.367
R537 B.n417 B.n416 163.367
R538 B.n418 B.n417 163.367
R539 B.n418 B.n85 163.367
R540 B.n422 B.n85 163.367
R541 B.n423 B.n422 163.367
R542 B.n424 B.n423 163.367
R543 B.n424 B.n83 163.367
R544 B.n428 B.n83 163.367
R545 B.n429 B.n428 163.367
R546 B.n430 B.n429 163.367
R547 B.n430 B.n81 163.367
R548 B.n434 B.n81 163.367
R549 B.n435 B.n434 163.367
R550 B.n436 B.n435 163.367
R551 B.n436 B.n79 163.367
R552 B.n440 B.n79 163.367
R553 B.n441 B.n440 163.367
R554 B.n442 B.n441 163.367
R555 B.n442 B.n77 163.367
R556 B.n446 B.n77 163.367
R557 B.n447 B.n446 163.367
R558 B.n448 B.n447 163.367
R559 B.n448 B.n75 163.367
R560 B.n452 B.n75 163.367
R561 B.n453 B.n452 163.367
R562 B.n454 B.n453 163.367
R563 B.n454 B.n73 163.367
R564 B.n458 B.n73 163.367
R565 B.n459 B.n458 163.367
R566 B.n460 B.n459 163.367
R567 B.n460 B.n71 163.367
R568 B.n464 B.n71 163.367
R569 B.n465 B.n464 163.367
R570 B.n466 B.n465 163.367
R571 B.n466 B.n69 163.367
R572 B.n603 B.n602 163.367
R573 B.n602 B.n21 163.367
R574 B.n598 B.n21 163.367
R575 B.n598 B.n597 163.367
R576 B.n597 B.n596 163.367
R577 B.n596 B.n23 163.367
R578 B.n592 B.n23 163.367
R579 B.n592 B.n591 163.367
R580 B.n591 B.n590 163.367
R581 B.n590 B.n25 163.367
R582 B.n586 B.n25 163.367
R583 B.n586 B.n585 163.367
R584 B.n585 B.n584 163.367
R585 B.n584 B.n27 163.367
R586 B.n580 B.n27 163.367
R587 B.n580 B.n579 163.367
R588 B.n579 B.n578 163.367
R589 B.n578 B.n29 163.367
R590 B.n574 B.n29 163.367
R591 B.n574 B.n573 163.367
R592 B.n573 B.n572 163.367
R593 B.n572 B.n31 163.367
R594 B.n568 B.n31 163.367
R595 B.n568 B.n567 163.367
R596 B.n567 B.n566 163.367
R597 B.n566 B.n33 163.367
R598 B.n562 B.n33 163.367
R599 B.n562 B.n561 163.367
R600 B.n561 B.n560 163.367
R601 B.n560 B.n35 163.367
R602 B.n556 B.n35 163.367
R603 B.n556 B.n555 163.367
R604 B.n555 B.n554 163.367
R605 B.n554 B.n37 163.367
R606 B.n550 B.n37 163.367
R607 B.n550 B.n549 163.367
R608 B.n549 B.n548 163.367
R609 B.n548 B.n39 163.367
R610 B.n544 B.n39 163.367
R611 B.n544 B.n543 163.367
R612 B.n543 B.n43 163.367
R613 B.n539 B.n43 163.367
R614 B.n539 B.n538 163.367
R615 B.n538 B.n537 163.367
R616 B.n537 B.n45 163.367
R617 B.n533 B.n45 163.367
R618 B.n533 B.n532 163.367
R619 B.n532 B.n531 163.367
R620 B.n531 B.n47 163.367
R621 B.n526 B.n47 163.367
R622 B.n526 B.n525 163.367
R623 B.n525 B.n524 163.367
R624 B.n524 B.n51 163.367
R625 B.n520 B.n51 163.367
R626 B.n520 B.n519 163.367
R627 B.n519 B.n518 163.367
R628 B.n518 B.n53 163.367
R629 B.n514 B.n53 163.367
R630 B.n514 B.n513 163.367
R631 B.n513 B.n512 163.367
R632 B.n512 B.n55 163.367
R633 B.n508 B.n55 163.367
R634 B.n508 B.n507 163.367
R635 B.n507 B.n506 163.367
R636 B.n506 B.n57 163.367
R637 B.n502 B.n57 163.367
R638 B.n502 B.n501 163.367
R639 B.n501 B.n500 163.367
R640 B.n500 B.n59 163.367
R641 B.n496 B.n59 163.367
R642 B.n496 B.n495 163.367
R643 B.n495 B.n494 163.367
R644 B.n494 B.n61 163.367
R645 B.n490 B.n61 163.367
R646 B.n490 B.n489 163.367
R647 B.n489 B.n488 163.367
R648 B.n488 B.n63 163.367
R649 B.n484 B.n63 163.367
R650 B.n484 B.n483 163.367
R651 B.n483 B.n482 163.367
R652 B.n482 B.n65 163.367
R653 B.n478 B.n65 163.367
R654 B.n478 B.n477 163.367
R655 B.n477 B.n476 163.367
R656 B.n476 B.n67 163.367
R657 B.n472 B.n67 163.367
R658 B.n472 B.n471 163.367
R659 B.n471 B.n470 163.367
R660 B.n127 B.n126 61.2853
R661 B.n133 B.n132 61.2853
R662 B.n41 B.n40 61.2853
R663 B.n49 B.n48 61.2853
R664 B.n299 B.n127 59.5399
R665 B.n134 B.n133 59.5399
R666 B.n42 B.n41 59.5399
R667 B.n529 B.n49 59.5399
R668 B.n469 B.n468 30.1273
R669 B.n605 B.n20 30.1273
R670 B.n360 B.n359 30.1273
R671 B.n223 B.n154 30.1273
R672 B B.n659 18.0485
R673 B.n601 B.n20 10.6151
R674 B.n601 B.n600 10.6151
R675 B.n600 B.n599 10.6151
R676 B.n599 B.n22 10.6151
R677 B.n595 B.n22 10.6151
R678 B.n595 B.n594 10.6151
R679 B.n594 B.n593 10.6151
R680 B.n593 B.n24 10.6151
R681 B.n589 B.n24 10.6151
R682 B.n589 B.n588 10.6151
R683 B.n588 B.n587 10.6151
R684 B.n587 B.n26 10.6151
R685 B.n583 B.n26 10.6151
R686 B.n583 B.n582 10.6151
R687 B.n582 B.n581 10.6151
R688 B.n581 B.n28 10.6151
R689 B.n577 B.n28 10.6151
R690 B.n577 B.n576 10.6151
R691 B.n576 B.n575 10.6151
R692 B.n575 B.n30 10.6151
R693 B.n571 B.n30 10.6151
R694 B.n571 B.n570 10.6151
R695 B.n570 B.n569 10.6151
R696 B.n569 B.n32 10.6151
R697 B.n565 B.n32 10.6151
R698 B.n565 B.n564 10.6151
R699 B.n564 B.n563 10.6151
R700 B.n563 B.n34 10.6151
R701 B.n559 B.n34 10.6151
R702 B.n559 B.n558 10.6151
R703 B.n558 B.n557 10.6151
R704 B.n557 B.n36 10.6151
R705 B.n553 B.n36 10.6151
R706 B.n553 B.n552 10.6151
R707 B.n552 B.n551 10.6151
R708 B.n551 B.n38 10.6151
R709 B.n547 B.n38 10.6151
R710 B.n547 B.n546 10.6151
R711 B.n546 B.n545 10.6151
R712 B.n542 B.n541 10.6151
R713 B.n541 B.n540 10.6151
R714 B.n540 B.n44 10.6151
R715 B.n536 B.n44 10.6151
R716 B.n536 B.n535 10.6151
R717 B.n535 B.n534 10.6151
R718 B.n534 B.n46 10.6151
R719 B.n530 B.n46 10.6151
R720 B.n528 B.n527 10.6151
R721 B.n527 B.n50 10.6151
R722 B.n523 B.n50 10.6151
R723 B.n523 B.n522 10.6151
R724 B.n522 B.n521 10.6151
R725 B.n521 B.n52 10.6151
R726 B.n517 B.n52 10.6151
R727 B.n517 B.n516 10.6151
R728 B.n516 B.n515 10.6151
R729 B.n515 B.n54 10.6151
R730 B.n511 B.n54 10.6151
R731 B.n511 B.n510 10.6151
R732 B.n510 B.n509 10.6151
R733 B.n509 B.n56 10.6151
R734 B.n505 B.n56 10.6151
R735 B.n505 B.n504 10.6151
R736 B.n504 B.n503 10.6151
R737 B.n503 B.n58 10.6151
R738 B.n499 B.n58 10.6151
R739 B.n499 B.n498 10.6151
R740 B.n498 B.n497 10.6151
R741 B.n497 B.n60 10.6151
R742 B.n493 B.n60 10.6151
R743 B.n493 B.n492 10.6151
R744 B.n492 B.n491 10.6151
R745 B.n491 B.n62 10.6151
R746 B.n487 B.n62 10.6151
R747 B.n487 B.n486 10.6151
R748 B.n486 B.n485 10.6151
R749 B.n485 B.n64 10.6151
R750 B.n481 B.n64 10.6151
R751 B.n481 B.n480 10.6151
R752 B.n480 B.n479 10.6151
R753 B.n479 B.n66 10.6151
R754 B.n475 B.n66 10.6151
R755 B.n475 B.n474 10.6151
R756 B.n474 B.n473 10.6151
R757 B.n473 B.n68 10.6151
R758 B.n469 B.n68 10.6151
R759 B.n361 B.n360 10.6151
R760 B.n361 B.n104 10.6151
R761 B.n365 B.n104 10.6151
R762 B.n366 B.n365 10.6151
R763 B.n367 B.n366 10.6151
R764 B.n367 B.n102 10.6151
R765 B.n371 B.n102 10.6151
R766 B.n372 B.n371 10.6151
R767 B.n373 B.n372 10.6151
R768 B.n373 B.n100 10.6151
R769 B.n377 B.n100 10.6151
R770 B.n378 B.n377 10.6151
R771 B.n379 B.n378 10.6151
R772 B.n379 B.n98 10.6151
R773 B.n383 B.n98 10.6151
R774 B.n384 B.n383 10.6151
R775 B.n385 B.n384 10.6151
R776 B.n385 B.n96 10.6151
R777 B.n389 B.n96 10.6151
R778 B.n390 B.n389 10.6151
R779 B.n391 B.n390 10.6151
R780 B.n391 B.n94 10.6151
R781 B.n395 B.n94 10.6151
R782 B.n396 B.n395 10.6151
R783 B.n397 B.n396 10.6151
R784 B.n397 B.n92 10.6151
R785 B.n401 B.n92 10.6151
R786 B.n402 B.n401 10.6151
R787 B.n403 B.n402 10.6151
R788 B.n403 B.n90 10.6151
R789 B.n407 B.n90 10.6151
R790 B.n408 B.n407 10.6151
R791 B.n409 B.n408 10.6151
R792 B.n409 B.n88 10.6151
R793 B.n413 B.n88 10.6151
R794 B.n414 B.n413 10.6151
R795 B.n415 B.n414 10.6151
R796 B.n415 B.n86 10.6151
R797 B.n419 B.n86 10.6151
R798 B.n420 B.n419 10.6151
R799 B.n421 B.n420 10.6151
R800 B.n421 B.n84 10.6151
R801 B.n425 B.n84 10.6151
R802 B.n426 B.n425 10.6151
R803 B.n427 B.n426 10.6151
R804 B.n427 B.n82 10.6151
R805 B.n431 B.n82 10.6151
R806 B.n432 B.n431 10.6151
R807 B.n433 B.n432 10.6151
R808 B.n433 B.n80 10.6151
R809 B.n437 B.n80 10.6151
R810 B.n438 B.n437 10.6151
R811 B.n439 B.n438 10.6151
R812 B.n439 B.n78 10.6151
R813 B.n443 B.n78 10.6151
R814 B.n444 B.n443 10.6151
R815 B.n445 B.n444 10.6151
R816 B.n445 B.n76 10.6151
R817 B.n449 B.n76 10.6151
R818 B.n450 B.n449 10.6151
R819 B.n451 B.n450 10.6151
R820 B.n451 B.n74 10.6151
R821 B.n455 B.n74 10.6151
R822 B.n456 B.n455 10.6151
R823 B.n457 B.n456 10.6151
R824 B.n457 B.n72 10.6151
R825 B.n461 B.n72 10.6151
R826 B.n462 B.n461 10.6151
R827 B.n463 B.n462 10.6151
R828 B.n463 B.n70 10.6151
R829 B.n467 B.n70 10.6151
R830 B.n468 B.n467 10.6151
R831 B.n227 B.n154 10.6151
R832 B.n228 B.n227 10.6151
R833 B.n229 B.n228 10.6151
R834 B.n229 B.n152 10.6151
R835 B.n233 B.n152 10.6151
R836 B.n234 B.n233 10.6151
R837 B.n235 B.n234 10.6151
R838 B.n235 B.n150 10.6151
R839 B.n239 B.n150 10.6151
R840 B.n240 B.n239 10.6151
R841 B.n241 B.n240 10.6151
R842 B.n241 B.n148 10.6151
R843 B.n245 B.n148 10.6151
R844 B.n246 B.n245 10.6151
R845 B.n247 B.n246 10.6151
R846 B.n247 B.n146 10.6151
R847 B.n251 B.n146 10.6151
R848 B.n252 B.n251 10.6151
R849 B.n253 B.n252 10.6151
R850 B.n253 B.n144 10.6151
R851 B.n257 B.n144 10.6151
R852 B.n258 B.n257 10.6151
R853 B.n259 B.n258 10.6151
R854 B.n259 B.n142 10.6151
R855 B.n263 B.n142 10.6151
R856 B.n264 B.n263 10.6151
R857 B.n265 B.n264 10.6151
R858 B.n265 B.n140 10.6151
R859 B.n269 B.n140 10.6151
R860 B.n270 B.n269 10.6151
R861 B.n271 B.n270 10.6151
R862 B.n271 B.n138 10.6151
R863 B.n275 B.n138 10.6151
R864 B.n276 B.n275 10.6151
R865 B.n277 B.n276 10.6151
R866 B.n277 B.n136 10.6151
R867 B.n281 B.n136 10.6151
R868 B.n282 B.n281 10.6151
R869 B.n283 B.n282 10.6151
R870 B.n287 B.n286 10.6151
R871 B.n288 B.n287 10.6151
R872 B.n288 B.n130 10.6151
R873 B.n292 B.n130 10.6151
R874 B.n293 B.n292 10.6151
R875 B.n294 B.n293 10.6151
R876 B.n294 B.n128 10.6151
R877 B.n298 B.n128 10.6151
R878 B.n301 B.n300 10.6151
R879 B.n301 B.n124 10.6151
R880 B.n305 B.n124 10.6151
R881 B.n306 B.n305 10.6151
R882 B.n307 B.n306 10.6151
R883 B.n307 B.n122 10.6151
R884 B.n311 B.n122 10.6151
R885 B.n312 B.n311 10.6151
R886 B.n313 B.n312 10.6151
R887 B.n313 B.n120 10.6151
R888 B.n317 B.n120 10.6151
R889 B.n318 B.n317 10.6151
R890 B.n319 B.n318 10.6151
R891 B.n319 B.n118 10.6151
R892 B.n323 B.n118 10.6151
R893 B.n324 B.n323 10.6151
R894 B.n325 B.n324 10.6151
R895 B.n325 B.n116 10.6151
R896 B.n329 B.n116 10.6151
R897 B.n330 B.n329 10.6151
R898 B.n331 B.n330 10.6151
R899 B.n331 B.n114 10.6151
R900 B.n335 B.n114 10.6151
R901 B.n336 B.n335 10.6151
R902 B.n337 B.n336 10.6151
R903 B.n337 B.n112 10.6151
R904 B.n341 B.n112 10.6151
R905 B.n342 B.n341 10.6151
R906 B.n343 B.n342 10.6151
R907 B.n343 B.n110 10.6151
R908 B.n347 B.n110 10.6151
R909 B.n348 B.n347 10.6151
R910 B.n349 B.n348 10.6151
R911 B.n349 B.n108 10.6151
R912 B.n353 B.n108 10.6151
R913 B.n354 B.n353 10.6151
R914 B.n355 B.n354 10.6151
R915 B.n355 B.n106 10.6151
R916 B.n359 B.n106 10.6151
R917 B.n223 B.n222 10.6151
R918 B.n222 B.n221 10.6151
R919 B.n221 B.n156 10.6151
R920 B.n217 B.n156 10.6151
R921 B.n217 B.n216 10.6151
R922 B.n216 B.n215 10.6151
R923 B.n215 B.n158 10.6151
R924 B.n211 B.n158 10.6151
R925 B.n211 B.n210 10.6151
R926 B.n210 B.n209 10.6151
R927 B.n209 B.n160 10.6151
R928 B.n205 B.n160 10.6151
R929 B.n205 B.n204 10.6151
R930 B.n204 B.n203 10.6151
R931 B.n203 B.n162 10.6151
R932 B.n199 B.n162 10.6151
R933 B.n199 B.n198 10.6151
R934 B.n198 B.n197 10.6151
R935 B.n197 B.n164 10.6151
R936 B.n193 B.n164 10.6151
R937 B.n193 B.n192 10.6151
R938 B.n192 B.n191 10.6151
R939 B.n191 B.n166 10.6151
R940 B.n187 B.n166 10.6151
R941 B.n187 B.n186 10.6151
R942 B.n186 B.n185 10.6151
R943 B.n185 B.n168 10.6151
R944 B.n181 B.n168 10.6151
R945 B.n181 B.n180 10.6151
R946 B.n180 B.n179 10.6151
R947 B.n179 B.n170 10.6151
R948 B.n175 B.n170 10.6151
R949 B.n175 B.n174 10.6151
R950 B.n174 B.n173 10.6151
R951 B.n173 B.n0 10.6151
R952 B.n655 B.n1 10.6151
R953 B.n655 B.n654 10.6151
R954 B.n654 B.n653 10.6151
R955 B.n653 B.n4 10.6151
R956 B.n649 B.n4 10.6151
R957 B.n649 B.n648 10.6151
R958 B.n648 B.n647 10.6151
R959 B.n647 B.n6 10.6151
R960 B.n643 B.n6 10.6151
R961 B.n643 B.n642 10.6151
R962 B.n642 B.n641 10.6151
R963 B.n641 B.n8 10.6151
R964 B.n637 B.n8 10.6151
R965 B.n637 B.n636 10.6151
R966 B.n636 B.n635 10.6151
R967 B.n635 B.n10 10.6151
R968 B.n631 B.n10 10.6151
R969 B.n631 B.n630 10.6151
R970 B.n630 B.n629 10.6151
R971 B.n629 B.n12 10.6151
R972 B.n625 B.n12 10.6151
R973 B.n625 B.n624 10.6151
R974 B.n624 B.n623 10.6151
R975 B.n623 B.n14 10.6151
R976 B.n619 B.n14 10.6151
R977 B.n619 B.n618 10.6151
R978 B.n618 B.n617 10.6151
R979 B.n617 B.n16 10.6151
R980 B.n613 B.n16 10.6151
R981 B.n613 B.n612 10.6151
R982 B.n612 B.n611 10.6151
R983 B.n611 B.n18 10.6151
R984 B.n607 B.n18 10.6151
R985 B.n607 B.n606 10.6151
R986 B.n606 B.n605 10.6151
R987 B.n542 B.n42 6.5566
R988 B.n530 B.n529 6.5566
R989 B.n286 B.n134 6.5566
R990 B.n299 B.n298 6.5566
R991 B.n545 B.n42 4.05904
R992 B.n529 B.n528 4.05904
R993 B.n283 B.n134 4.05904
R994 B.n300 B.n299 4.05904
R995 B.n659 B.n0 2.81026
R996 B.n659 B.n1 2.81026
R997 VN.n0 VN.t2 131.362
R998 VN.n1 VN.t1 131.362
R999 VN.n0 VN.t3 130.466
R1000 VN.n1 VN.t0 130.466
R1001 VN VN.n1 50.1996
R1002 VN VN.n0 3.45334
R1003 VDD2.n2 VDD2.n0 114.067
R1004 VDD2.n2 VDD2.n1 72.4555
R1005 VDD2.n1 VDD2.t0 2.88215
R1006 VDD2.n1 VDD2.t1 2.88215
R1007 VDD2.n0 VDD2.t3 2.88215
R1008 VDD2.n0 VDD2.t2 2.88215
R1009 VDD2 VDD2.n2 0.0586897
R1010 VTAIL.n490 VTAIL.n434 756.745
R1011 VTAIL.n56 VTAIL.n0 756.745
R1012 VTAIL.n118 VTAIL.n62 756.745
R1013 VTAIL.n180 VTAIL.n124 756.745
R1014 VTAIL.n428 VTAIL.n372 756.745
R1015 VTAIL.n366 VTAIL.n310 756.745
R1016 VTAIL.n304 VTAIL.n248 756.745
R1017 VTAIL.n242 VTAIL.n186 756.745
R1018 VTAIL.n455 VTAIL.n454 585
R1019 VTAIL.n457 VTAIL.n456 585
R1020 VTAIL.n450 VTAIL.n449 585
R1021 VTAIL.n463 VTAIL.n462 585
R1022 VTAIL.n465 VTAIL.n464 585
R1023 VTAIL.n446 VTAIL.n445 585
R1024 VTAIL.n472 VTAIL.n471 585
R1025 VTAIL.n473 VTAIL.n444 585
R1026 VTAIL.n475 VTAIL.n474 585
R1027 VTAIL.n442 VTAIL.n441 585
R1028 VTAIL.n481 VTAIL.n480 585
R1029 VTAIL.n483 VTAIL.n482 585
R1030 VTAIL.n438 VTAIL.n437 585
R1031 VTAIL.n489 VTAIL.n488 585
R1032 VTAIL.n491 VTAIL.n490 585
R1033 VTAIL.n21 VTAIL.n20 585
R1034 VTAIL.n23 VTAIL.n22 585
R1035 VTAIL.n16 VTAIL.n15 585
R1036 VTAIL.n29 VTAIL.n28 585
R1037 VTAIL.n31 VTAIL.n30 585
R1038 VTAIL.n12 VTAIL.n11 585
R1039 VTAIL.n38 VTAIL.n37 585
R1040 VTAIL.n39 VTAIL.n10 585
R1041 VTAIL.n41 VTAIL.n40 585
R1042 VTAIL.n8 VTAIL.n7 585
R1043 VTAIL.n47 VTAIL.n46 585
R1044 VTAIL.n49 VTAIL.n48 585
R1045 VTAIL.n4 VTAIL.n3 585
R1046 VTAIL.n55 VTAIL.n54 585
R1047 VTAIL.n57 VTAIL.n56 585
R1048 VTAIL.n83 VTAIL.n82 585
R1049 VTAIL.n85 VTAIL.n84 585
R1050 VTAIL.n78 VTAIL.n77 585
R1051 VTAIL.n91 VTAIL.n90 585
R1052 VTAIL.n93 VTAIL.n92 585
R1053 VTAIL.n74 VTAIL.n73 585
R1054 VTAIL.n100 VTAIL.n99 585
R1055 VTAIL.n101 VTAIL.n72 585
R1056 VTAIL.n103 VTAIL.n102 585
R1057 VTAIL.n70 VTAIL.n69 585
R1058 VTAIL.n109 VTAIL.n108 585
R1059 VTAIL.n111 VTAIL.n110 585
R1060 VTAIL.n66 VTAIL.n65 585
R1061 VTAIL.n117 VTAIL.n116 585
R1062 VTAIL.n119 VTAIL.n118 585
R1063 VTAIL.n145 VTAIL.n144 585
R1064 VTAIL.n147 VTAIL.n146 585
R1065 VTAIL.n140 VTAIL.n139 585
R1066 VTAIL.n153 VTAIL.n152 585
R1067 VTAIL.n155 VTAIL.n154 585
R1068 VTAIL.n136 VTAIL.n135 585
R1069 VTAIL.n162 VTAIL.n161 585
R1070 VTAIL.n163 VTAIL.n134 585
R1071 VTAIL.n165 VTAIL.n164 585
R1072 VTAIL.n132 VTAIL.n131 585
R1073 VTAIL.n171 VTAIL.n170 585
R1074 VTAIL.n173 VTAIL.n172 585
R1075 VTAIL.n128 VTAIL.n127 585
R1076 VTAIL.n179 VTAIL.n178 585
R1077 VTAIL.n181 VTAIL.n180 585
R1078 VTAIL.n429 VTAIL.n428 585
R1079 VTAIL.n427 VTAIL.n426 585
R1080 VTAIL.n376 VTAIL.n375 585
R1081 VTAIL.n421 VTAIL.n420 585
R1082 VTAIL.n419 VTAIL.n418 585
R1083 VTAIL.n380 VTAIL.n379 585
R1084 VTAIL.n384 VTAIL.n382 585
R1085 VTAIL.n413 VTAIL.n412 585
R1086 VTAIL.n411 VTAIL.n410 585
R1087 VTAIL.n386 VTAIL.n385 585
R1088 VTAIL.n405 VTAIL.n404 585
R1089 VTAIL.n403 VTAIL.n402 585
R1090 VTAIL.n390 VTAIL.n389 585
R1091 VTAIL.n397 VTAIL.n396 585
R1092 VTAIL.n395 VTAIL.n394 585
R1093 VTAIL.n367 VTAIL.n366 585
R1094 VTAIL.n365 VTAIL.n364 585
R1095 VTAIL.n314 VTAIL.n313 585
R1096 VTAIL.n359 VTAIL.n358 585
R1097 VTAIL.n357 VTAIL.n356 585
R1098 VTAIL.n318 VTAIL.n317 585
R1099 VTAIL.n322 VTAIL.n320 585
R1100 VTAIL.n351 VTAIL.n350 585
R1101 VTAIL.n349 VTAIL.n348 585
R1102 VTAIL.n324 VTAIL.n323 585
R1103 VTAIL.n343 VTAIL.n342 585
R1104 VTAIL.n341 VTAIL.n340 585
R1105 VTAIL.n328 VTAIL.n327 585
R1106 VTAIL.n335 VTAIL.n334 585
R1107 VTAIL.n333 VTAIL.n332 585
R1108 VTAIL.n305 VTAIL.n304 585
R1109 VTAIL.n303 VTAIL.n302 585
R1110 VTAIL.n252 VTAIL.n251 585
R1111 VTAIL.n297 VTAIL.n296 585
R1112 VTAIL.n295 VTAIL.n294 585
R1113 VTAIL.n256 VTAIL.n255 585
R1114 VTAIL.n260 VTAIL.n258 585
R1115 VTAIL.n289 VTAIL.n288 585
R1116 VTAIL.n287 VTAIL.n286 585
R1117 VTAIL.n262 VTAIL.n261 585
R1118 VTAIL.n281 VTAIL.n280 585
R1119 VTAIL.n279 VTAIL.n278 585
R1120 VTAIL.n266 VTAIL.n265 585
R1121 VTAIL.n273 VTAIL.n272 585
R1122 VTAIL.n271 VTAIL.n270 585
R1123 VTAIL.n243 VTAIL.n242 585
R1124 VTAIL.n241 VTAIL.n240 585
R1125 VTAIL.n190 VTAIL.n189 585
R1126 VTAIL.n235 VTAIL.n234 585
R1127 VTAIL.n233 VTAIL.n232 585
R1128 VTAIL.n194 VTAIL.n193 585
R1129 VTAIL.n198 VTAIL.n196 585
R1130 VTAIL.n227 VTAIL.n226 585
R1131 VTAIL.n225 VTAIL.n224 585
R1132 VTAIL.n200 VTAIL.n199 585
R1133 VTAIL.n219 VTAIL.n218 585
R1134 VTAIL.n217 VTAIL.n216 585
R1135 VTAIL.n204 VTAIL.n203 585
R1136 VTAIL.n211 VTAIL.n210 585
R1137 VTAIL.n209 VTAIL.n208 585
R1138 VTAIL.n453 VTAIL.t2 329.036
R1139 VTAIL.n19 VTAIL.t3 329.036
R1140 VTAIL.n81 VTAIL.t6 329.036
R1141 VTAIL.n143 VTAIL.t1 329.036
R1142 VTAIL.n393 VTAIL.t0 329.036
R1143 VTAIL.n331 VTAIL.t7 329.036
R1144 VTAIL.n269 VTAIL.t4 329.036
R1145 VTAIL.n207 VTAIL.t5 329.036
R1146 VTAIL.n456 VTAIL.n455 171.744
R1147 VTAIL.n456 VTAIL.n449 171.744
R1148 VTAIL.n463 VTAIL.n449 171.744
R1149 VTAIL.n464 VTAIL.n463 171.744
R1150 VTAIL.n464 VTAIL.n445 171.744
R1151 VTAIL.n472 VTAIL.n445 171.744
R1152 VTAIL.n473 VTAIL.n472 171.744
R1153 VTAIL.n474 VTAIL.n473 171.744
R1154 VTAIL.n474 VTAIL.n441 171.744
R1155 VTAIL.n481 VTAIL.n441 171.744
R1156 VTAIL.n482 VTAIL.n481 171.744
R1157 VTAIL.n482 VTAIL.n437 171.744
R1158 VTAIL.n489 VTAIL.n437 171.744
R1159 VTAIL.n490 VTAIL.n489 171.744
R1160 VTAIL.n22 VTAIL.n21 171.744
R1161 VTAIL.n22 VTAIL.n15 171.744
R1162 VTAIL.n29 VTAIL.n15 171.744
R1163 VTAIL.n30 VTAIL.n29 171.744
R1164 VTAIL.n30 VTAIL.n11 171.744
R1165 VTAIL.n38 VTAIL.n11 171.744
R1166 VTAIL.n39 VTAIL.n38 171.744
R1167 VTAIL.n40 VTAIL.n39 171.744
R1168 VTAIL.n40 VTAIL.n7 171.744
R1169 VTAIL.n47 VTAIL.n7 171.744
R1170 VTAIL.n48 VTAIL.n47 171.744
R1171 VTAIL.n48 VTAIL.n3 171.744
R1172 VTAIL.n55 VTAIL.n3 171.744
R1173 VTAIL.n56 VTAIL.n55 171.744
R1174 VTAIL.n84 VTAIL.n83 171.744
R1175 VTAIL.n84 VTAIL.n77 171.744
R1176 VTAIL.n91 VTAIL.n77 171.744
R1177 VTAIL.n92 VTAIL.n91 171.744
R1178 VTAIL.n92 VTAIL.n73 171.744
R1179 VTAIL.n100 VTAIL.n73 171.744
R1180 VTAIL.n101 VTAIL.n100 171.744
R1181 VTAIL.n102 VTAIL.n101 171.744
R1182 VTAIL.n102 VTAIL.n69 171.744
R1183 VTAIL.n109 VTAIL.n69 171.744
R1184 VTAIL.n110 VTAIL.n109 171.744
R1185 VTAIL.n110 VTAIL.n65 171.744
R1186 VTAIL.n117 VTAIL.n65 171.744
R1187 VTAIL.n118 VTAIL.n117 171.744
R1188 VTAIL.n146 VTAIL.n145 171.744
R1189 VTAIL.n146 VTAIL.n139 171.744
R1190 VTAIL.n153 VTAIL.n139 171.744
R1191 VTAIL.n154 VTAIL.n153 171.744
R1192 VTAIL.n154 VTAIL.n135 171.744
R1193 VTAIL.n162 VTAIL.n135 171.744
R1194 VTAIL.n163 VTAIL.n162 171.744
R1195 VTAIL.n164 VTAIL.n163 171.744
R1196 VTAIL.n164 VTAIL.n131 171.744
R1197 VTAIL.n171 VTAIL.n131 171.744
R1198 VTAIL.n172 VTAIL.n171 171.744
R1199 VTAIL.n172 VTAIL.n127 171.744
R1200 VTAIL.n179 VTAIL.n127 171.744
R1201 VTAIL.n180 VTAIL.n179 171.744
R1202 VTAIL.n428 VTAIL.n427 171.744
R1203 VTAIL.n427 VTAIL.n375 171.744
R1204 VTAIL.n420 VTAIL.n375 171.744
R1205 VTAIL.n420 VTAIL.n419 171.744
R1206 VTAIL.n419 VTAIL.n379 171.744
R1207 VTAIL.n384 VTAIL.n379 171.744
R1208 VTAIL.n412 VTAIL.n384 171.744
R1209 VTAIL.n412 VTAIL.n411 171.744
R1210 VTAIL.n411 VTAIL.n385 171.744
R1211 VTAIL.n404 VTAIL.n385 171.744
R1212 VTAIL.n404 VTAIL.n403 171.744
R1213 VTAIL.n403 VTAIL.n389 171.744
R1214 VTAIL.n396 VTAIL.n389 171.744
R1215 VTAIL.n396 VTAIL.n395 171.744
R1216 VTAIL.n366 VTAIL.n365 171.744
R1217 VTAIL.n365 VTAIL.n313 171.744
R1218 VTAIL.n358 VTAIL.n313 171.744
R1219 VTAIL.n358 VTAIL.n357 171.744
R1220 VTAIL.n357 VTAIL.n317 171.744
R1221 VTAIL.n322 VTAIL.n317 171.744
R1222 VTAIL.n350 VTAIL.n322 171.744
R1223 VTAIL.n350 VTAIL.n349 171.744
R1224 VTAIL.n349 VTAIL.n323 171.744
R1225 VTAIL.n342 VTAIL.n323 171.744
R1226 VTAIL.n342 VTAIL.n341 171.744
R1227 VTAIL.n341 VTAIL.n327 171.744
R1228 VTAIL.n334 VTAIL.n327 171.744
R1229 VTAIL.n334 VTAIL.n333 171.744
R1230 VTAIL.n304 VTAIL.n303 171.744
R1231 VTAIL.n303 VTAIL.n251 171.744
R1232 VTAIL.n296 VTAIL.n251 171.744
R1233 VTAIL.n296 VTAIL.n295 171.744
R1234 VTAIL.n295 VTAIL.n255 171.744
R1235 VTAIL.n260 VTAIL.n255 171.744
R1236 VTAIL.n288 VTAIL.n260 171.744
R1237 VTAIL.n288 VTAIL.n287 171.744
R1238 VTAIL.n287 VTAIL.n261 171.744
R1239 VTAIL.n280 VTAIL.n261 171.744
R1240 VTAIL.n280 VTAIL.n279 171.744
R1241 VTAIL.n279 VTAIL.n265 171.744
R1242 VTAIL.n272 VTAIL.n265 171.744
R1243 VTAIL.n272 VTAIL.n271 171.744
R1244 VTAIL.n242 VTAIL.n241 171.744
R1245 VTAIL.n241 VTAIL.n189 171.744
R1246 VTAIL.n234 VTAIL.n189 171.744
R1247 VTAIL.n234 VTAIL.n233 171.744
R1248 VTAIL.n233 VTAIL.n193 171.744
R1249 VTAIL.n198 VTAIL.n193 171.744
R1250 VTAIL.n226 VTAIL.n198 171.744
R1251 VTAIL.n226 VTAIL.n225 171.744
R1252 VTAIL.n225 VTAIL.n199 171.744
R1253 VTAIL.n218 VTAIL.n199 171.744
R1254 VTAIL.n218 VTAIL.n217 171.744
R1255 VTAIL.n217 VTAIL.n203 171.744
R1256 VTAIL.n210 VTAIL.n203 171.744
R1257 VTAIL.n210 VTAIL.n209 171.744
R1258 VTAIL.n455 VTAIL.t2 85.8723
R1259 VTAIL.n21 VTAIL.t3 85.8723
R1260 VTAIL.n83 VTAIL.t6 85.8723
R1261 VTAIL.n145 VTAIL.t1 85.8723
R1262 VTAIL.n395 VTAIL.t0 85.8723
R1263 VTAIL.n333 VTAIL.t7 85.8723
R1264 VTAIL.n271 VTAIL.t4 85.8723
R1265 VTAIL.n209 VTAIL.t5 85.8723
R1266 VTAIL.n495 VTAIL.n494 29.8581
R1267 VTAIL.n61 VTAIL.n60 29.8581
R1268 VTAIL.n123 VTAIL.n122 29.8581
R1269 VTAIL.n185 VTAIL.n184 29.8581
R1270 VTAIL.n433 VTAIL.n432 29.8581
R1271 VTAIL.n371 VTAIL.n370 29.8581
R1272 VTAIL.n309 VTAIL.n308 29.8581
R1273 VTAIL.n247 VTAIL.n246 29.8581
R1274 VTAIL.n495 VTAIL.n433 24.8152
R1275 VTAIL.n247 VTAIL.n185 24.8152
R1276 VTAIL.n475 VTAIL.n442 13.1884
R1277 VTAIL.n41 VTAIL.n8 13.1884
R1278 VTAIL.n103 VTAIL.n70 13.1884
R1279 VTAIL.n165 VTAIL.n132 13.1884
R1280 VTAIL.n382 VTAIL.n380 13.1884
R1281 VTAIL.n320 VTAIL.n318 13.1884
R1282 VTAIL.n258 VTAIL.n256 13.1884
R1283 VTAIL.n196 VTAIL.n194 13.1884
R1284 VTAIL.n476 VTAIL.n444 12.8005
R1285 VTAIL.n480 VTAIL.n479 12.8005
R1286 VTAIL.n42 VTAIL.n10 12.8005
R1287 VTAIL.n46 VTAIL.n45 12.8005
R1288 VTAIL.n104 VTAIL.n72 12.8005
R1289 VTAIL.n108 VTAIL.n107 12.8005
R1290 VTAIL.n166 VTAIL.n134 12.8005
R1291 VTAIL.n170 VTAIL.n169 12.8005
R1292 VTAIL.n418 VTAIL.n417 12.8005
R1293 VTAIL.n414 VTAIL.n413 12.8005
R1294 VTAIL.n356 VTAIL.n355 12.8005
R1295 VTAIL.n352 VTAIL.n351 12.8005
R1296 VTAIL.n294 VTAIL.n293 12.8005
R1297 VTAIL.n290 VTAIL.n289 12.8005
R1298 VTAIL.n232 VTAIL.n231 12.8005
R1299 VTAIL.n228 VTAIL.n227 12.8005
R1300 VTAIL.n471 VTAIL.n470 12.0247
R1301 VTAIL.n483 VTAIL.n440 12.0247
R1302 VTAIL.n37 VTAIL.n36 12.0247
R1303 VTAIL.n49 VTAIL.n6 12.0247
R1304 VTAIL.n99 VTAIL.n98 12.0247
R1305 VTAIL.n111 VTAIL.n68 12.0247
R1306 VTAIL.n161 VTAIL.n160 12.0247
R1307 VTAIL.n173 VTAIL.n130 12.0247
R1308 VTAIL.n421 VTAIL.n378 12.0247
R1309 VTAIL.n410 VTAIL.n383 12.0247
R1310 VTAIL.n359 VTAIL.n316 12.0247
R1311 VTAIL.n348 VTAIL.n321 12.0247
R1312 VTAIL.n297 VTAIL.n254 12.0247
R1313 VTAIL.n286 VTAIL.n259 12.0247
R1314 VTAIL.n235 VTAIL.n192 12.0247
R1315 VTAIL.n224 VTAIL.n197 12.0247
R1316 VTAIL.n469 VTAIL.n446 11.249
R1317 VTAIL.n484 VTAIL.n438 11.249
R1318 VTAIL.n35 VTAIL.n12 11.249
R1319 VTAIL.n50 VTAIL.n4 11.249
R1320 VTAIL.n97 VTAIL.n74 11.249
R1321 VTAIL.n112 VTAIL.n66 11.249
R1322 VTAIL.n159 VTAIL.n136 11.249
R1323 VTAIL.n174 VTAIL.n128 11.249
R1324 VTAIL.n422 VTAIL.n376 11.249
R1325 VTAIL.n409 VTAIL.n386 11.249
R1326 VTAIL.n360 VTAIL.n314 11.249
R1327 VTAIL.n347 VTAIL.n324 11.249
R1328 VTAIL.n298 VTAIL.n252 11.249
R1329 VTAIL.n285 VTAIL.n262 11.249
R1330 VTAIL.n236 VTAIL.n190 11.249
R1331 VTAIL.n223 VTAIL.n200 11.249
R1332 VTAIL.n454 VTAIL.n453 10.7239
R1333 VTAIL.n20 VTAIL.n19 10.7239
R1334 VTAIL.n82 VTAIL.n81 10.7239
R1335 VTAIL.n144 VTAIL.n143 10.7239
R1336 VTAIL.n394 VTAIL.n393 10.7239
R1337 VTAIL.n332 VTAIL.n331 10.7239
R1338 VTAIL.n270 VTAIL.n269 10.7239
R1339 VTAIL.n208 VTAIL.n207 10.7239
R1340 VTAIL.n466 VTAIL.n465 10.4732
R1341 VTAIL.n488 VTAIL.n487 10.4732
R1342 VTAIL.n32 VTAIL.n31 10.4732
R1343 VTAIL.n54 VTAIL.n53 10.4732
R1344 VTAIL.n94 VTAIL.n93 10.4732
R1345 VTAIL.n116 VTAIL.n115 10.4732
R1346 VTAIL.n156 VTAIL.n155 10.4732
R1347 VTAIL.n178 VTAIL.n177 10.4732
R1348 VTAIL.n426 VTAIL.n425 10.4732
R1349 VTAIL.n406 VTAIL.n405 10.4732
R1350 VTAIL.n364 VTAIL.n363 10.4732
R1351 VTAIL.n344 VTAIL.n343 10.4732
R1352 VTAIL.n302 VTAIL.n301 10.4732
R1353 VTAIL.n282 VTAIL.n281 10.4732
R1354 VTAIL.n240 VTAIL.n239 10.4732
R1355 VTAIL.n220 VTAIL.n219 10.4732
R1356 VTAIL.n462 VTAIL.n448 9.69747
R1357 VTAIL.n491 VTAIL.n436 9.69747
R1358 VTAIL.n28 VTAIL.n14 9.69747
R1359 VTAIL.n57 VTAIL.n2 9.69747
R1360 VTAIL.n90 VTAIL.n76 9.69747
R1361 VTAIL.n119 VTAIL.n64 9.69747
R1362 VTAIL.n152 VTAIL.n138 9.69747
R1363 VTAIL.n181 VTAIL.n126 9.69747
R1364 VTAIL.n429 VTAIL.n374 9.69747
R1365 VTAIL.n402 VTAIL.n388 9.69747
R1366 VTAIL.n367 VTAIL.n312 9.69747
R1367 VTAIL.n340 VTAIL.n326 9.69747
R1368 VTAIL.n305 VTAIL.n250 9.69747
R1369 VTAIL.n278 VTAIL.n264 9.69747
R1370 VTAIL.n243 VTAIL.n188 9.69747
R1371 VTAIL.n216 VTAIL.n202 9.69747
R1372 VTAIL.n494 VTAIL.n493 9.45567
R1373 VTAIL.n60 VTAIL.n59 9.45567
R1374 VTAIL.n122 VTAIL.n121 9.45567
R1375 VTAIL.n184 VTAIL.n183 9.45567
R1376 VTAIL.n432 VTAIL.n431 9.45567
R1377 VTAIL.n370 VTAIL.n369 9.45567
R1378 VTAIL.n308 VTAIL.n307 9.45567
R1379 VTAIL.n246 VTAIL.n245 9.45567
R1380 VTAIL.n493 VTAIL.n492 9.3005
R1381 VTAIL.n436 VTAIL.n435 9.3005
R1382 VTAIL.n487 VTAIL.n486 9.3005
R1383 VTAIL.n485 VTAIL.n484 9.3005
R1384 VTAIL.n440 VTAIL.n439 9.3005
R1385 VTAIL.n479 VTAIL.n478 9.3005
R1386 VTAIL.n452 VTAIL.n451 9.3005
R1387 VTAIL.n459 VTAIL.n458 9.3005
R1388 VTAIL.n461 VTAIL.n460 9.3005
R1389 VTAIL.n448 VTAIL.n447 9.3005
R1390 VTAIL.n467 VTAIL.n466 9.3005
R1391 VTAIL.n469 VTAIL.n468 9.3005
R1392 VTAIL.n470 VTAIL.n443 9.3005
R1393 VTAIL.n477 VTAIL.n476 9.3005
R1394 VTAIL.n59 VTAIL.n58 9.3005
R1395 VTAIL.n2 VTAIL.n1 9.3005
R1396 VTAIL.n53 VTAIL.n52 9.3005
R1397 VTAIL.n51 VTAIL.n50 9.3005
R1398 VTAIL.n6 VTAIL.n5 9.3005
R1399 VTAIL.n45 VTAIL.n44 9.3005
R1400 VTAIL.n18 VTAIL.n17 9.3005
R1401 VTAIL.n25 VTAIL.n24 9.3005
R1402 VTAIL.n27 VTAIL.n26 9.3005
R1403 VTAIL.n14 VTAIL.n13 9.3005
R1404 VTAIL.n33 VTAIL.n32 9.3005
R1405 VTAIL.n35 VTAIL.n34 9.3005
R1406 VTAIL.n36 VTAIL.n9 9.3005
R1407 VTAIL.n43 VTAIL.n42 9.3005
R1408 VTAIL.n121 VTAIL.n120 9.3005
R1409 VTAIL.n64 VTAIL.n63 9.3005
R1410 VTAIL.n115 VTAIL.n114 9.3005
R1411 VTAIL.n113 VTAIL.n112 9.3005
R1412 VTAIL.n68 VTAIL.n67 9.3005
R1413 VTAIL.n107 VTAIL.n106 9.3005
R1414 VTAIL.n80 VTAIL.n79 9.3005
R1415 VTAIL.n87 VTAIL.n86 9.3005
R1416 VTAIL.n89 VTAIL.n88 9.3005
R1417 VTAIL.n76 VTAIL.n75 9.3005
R1418 VTAIL.n95 VTAIL.n94 9.3005
R1419 VTAIL.n97 VTAIL.n96 9.3005
R1420 VTAIL.n98 VTAIL.n71 9.3005
R1421 VTAIL.n105 VTAIL.n104 9.3005
R1422 VTAIL.n183 VTAIL.n182 9.3005
R1423 VTAIL.n126 VTAIL.n125 9.3005
R1424 VTAIL.n177 VTAIL.n176 9.3005
R1425 VTAIL.n175 VTAIL.n174 9.3005
R1426 VTAIL.n130 VTAIL.n129 9.3005
R1427 VTAIL.n169 VTAIL.n168 9.3005
R1428 VTAIL.n142 VTAIL.n141 9.3005
R1429 VTAIL.n149 VTAIL.n148 9.3005
R1430 VTAIL.n151 VTAIL.n150 9.3005
R1431 VTAIL.n138 VTAIL.n137 9.3005
R1432 VTAIL.n157 VTAIL.n156 9.3005
R1433 VTAIL.n159 VTAIL.n158 9.3005
R1434 VTAIL.n160 VTAIL.n133 9.3005
R1435 VTAIL.n167 VTAIL.n166 9.3005
R1436 VTAIL.n392 VTAIL.n391 9.3005
R1437 VTAIL.n399 VTAIL.n398 9.3005
R1438 VTAIL.n401 VTAIL.n400 9.3005
R1439 VTAIL.n388 VTAIL.n387 9.3005
R1440 VTAIL.n407 VTAIL.n406 9.3005
R1441 VTAIL.n409 VTAIL.n408 9.3005
R1442 VTAIL.n383 VTAIL.n381 9.3005
R1443 VTAIL.n415 VTAIL.n414 9.3005
R1444 VTAIL.n431 VTAIL.n430 9.3005
R1445 VTAIL.n374 VTAIL.n373 9.3005
R1446 VTAIL.n425 VTAIL.n424 9.3005
R1447 VTAIL.n423 VTAIL.n422 9.3005
R1448 VTAIL.n378 VTAIL.n377 9.3005
R1449 VTAIL.n417 VTAIL.n416 9.3005
R1450 VTAIL.n330 VTAIL.n329 9.3005
R1451 VTAIL.n337 VTAIL.n336 9.3005
R1452 VTAIL.n339 VTAIL.n338 9.3005
R1453 VTAIL.n326 VTAIL.n325 9.3005
R1454 VTAIL.n345 VTAIL.n344 9.3005
R1455 VTAIL.n347 VTAIL.n346 9.3005
R1456 VTAIL.n321 VTAIL.n319 9.3005
R1457 VTAIL.n353 VTAIL.n352 9.3005
R1458 VTAIL.n369 VTAIL.n368 9.3005
R1459 VTAIL.n312 VTAIL.n311 9.3005
R1460 VTAIL.n363 VTAIL.n362 9.3005
R1461 VTAIL.n361 VTAIL.n360 9.3005
R1462 VTAIL.n316 VTAIL.n315 9.3005
R1463 VTAIL.n355 VTAIL.n354 9.3005
R1464 VTAIL.n268 VTAIL.n267 9.3005
R1465 VTAIL.n275 VTAIL.n274 9.3005
R1466 VTAIL.n277 VTAIL.n276 9.3005
R1467 VTAIL.n264 VTAIL.n263 9.3005
R1468 VTAIL.n283 VTAIL.n282 9.3005
R1469 VTAIL.n285 VTAIL.n284 9.3005
R1470 VTAIL.n259 VTAIL.n257 9.3005
R1471 VTAIL.n291 VTAIL.n290 9.3005
R1472 VTAIL.n307 VTAIL.n306 9.3005
R1473 VTAIL.n250 VTAIL.n249 9.3005
R1474 VTAIL.n301 VTAIL.n300 9.3005
R1475 VTAIL.n299 VTAIL.n298 9.3005
R1476 VTAIL.n254 VTAIL.n253 9.3005
R1477 VTAIL.n293 VTAIL.n292 9.3005
R1478 VTAIL.n206 VTAIL.n205 9.3005
R1479 VTAIL.n213 VTAIL.n212 9.3005
R1480 VTAIL.n215 VTAIL.n214 9.3005
R1481 VTAIL.n202 VTAIL.n201 9.3005
R1482 VTAIL.n221 VTAIL.n220 9.3005
R1483 VTAIL.n223 VTAIL.n222 9.3005
R1484 VTAIL.n197 VTAIL.n195 9.3005
R1485 VTAIL.n229 VTAIL.n228 9.3005
R1486 VTAIL.n245 VTAIL.n244 9.3005
R1487 VTAIL.n188 VTAIL.n187 9.3005
R1488 VTAIL.n239 VTAIL.n238 9.3005
R1489 VTAIL.n237 VTAIL.n236 9.3005
R1490 VTAIL.n192 VTAIL.n191 9.3005
R1491 VTAIL.n231 VTAIL.n230 9.3005
R1492 VTAIL.n461 VTAIL.n450 8.92171
R1493 VTAIL.n492 VTAIL.n434 8.92171
R1494 VTAIL.n27 VTAIL.n16 8.92171
R1495 VTAIL.n58 VTAIL.n0 8.92171
R1496 VTAIL.n89 VTAIL.n78 8.92171
R1497 VTAIL.n120 VTAIL.n62 8.92171
R1498 VTAIL.n151 VTAIL.n140 8.92171
R1499 VTAIL.n182 VTAIL.n124 8.92171
R1500 VTAIL.n430 VTAIL.n372 8.92171
R1501 VTAIL.n401 VTAIL.n390 8.92171
R1502 VTAIL.n368 VTAIL.n310 8.92171
R1503 VTAIL.n339 VTAIL.n328 8.92171
R1504 VTAIL.n306 VTAIL.n248 8.92171
R1505 VTAIL.n277 VTAIL.n266 8.92171
R1506 VTAIL.n244 VTAIL.n186 8.92171
R1507 VTAIL.n215 VTAIL.n204 8.92171
R1508 VTAIL.n458 VTAIL.n457 8.14595
R1509 VTAIL.n24 VTAIL.n23 8.14595
R1510 VTAIL.n86 VTAIL.n85 8.14595
R1511 VTAIL.n148 VTAIL.n147 8.14595
R1512 VTAIL.n398 VTAIL.n397 8.14595
R1513 VTAIL.n336 VTAIL.n335 8.14595
R1514 VTAIL.n274 VTAIL.n273 8.14595
R1515 VTAIL.n212 VTAIL.n211 8.14595
R1516 VTAIL.n454 VTAIL.n452 7.3702
R1517 VTAIL.n20 VTAIL.n18 7.3702
R1518 VTAIL.n82 VTAIL.n80 7.3702
R1519 VTAIL.n144 VTAIL.n142 7.3702
R1520 VTAIL.n394 VTAIL.n392 7.3702
R1521 VTAIL.n332 VTAIL.n330 7.3702
R1522 VTAIL.n270 VTAIL.n268 7.3702
R1523 VTAIL.n208 VTAIL.n206 7.3702
R1524 VTAIL.n457 VTAIL.n452 5.81868
R1525 VTAIL.n23 VTAIL.n18 5.81868
R1526 VTAIL.n85 VTAIL.n80 5.81868
R1527 VTAIL.n147 VTAIL.n142 5.81868
R1528 VTAIL.n397 VTAIL.n392 5.81868
R1529 VTAIL.n335 VTAIL.n330 5.81868
R1530 VTAIL.n273 VTAIL.n268 5.81868
R1531 VTAIL.n211 VTAIL.n206 5.81868
R1532 VTAIL.n458 VTAIL.n450 5.04292
R1533 VTAIL.n494 VTAIL.n434 5.04292
R1534 VTAIL.n24 VTAIL.n16 5.04292
R1535 VTAIL.n60 VTAIL.n0 5.04292
R1536 VTAIL.n86 VTAIL.n78 5.04292
R1537 VTAIL.n122 VTAIL.n62 5.04292
R1538 VTAIL.n148 VTAIL.n140 5.04292
R1539 VTAIL.n184 VTAIL.n124 5.04292
R1540 VTAIL.n432 VTAIL.n372 5.04292
R1541 VTAIL.n398 VTAIL.n390 5.04292
R1542 VTAIL.n370 VTAIL.n310 5.04292
R1543 VTAIL.n336 VTAIL.n328 5.04292
R1544 VTAIL.n308 VTAIL.n248 5.04292
R1545 VTAIL.n274 VTAIL.n266 5.04292
R1546 VTAIL.n246 VTAIL.n186 5.04292
R1547 VTAIL.n212 VTAIL.n204 5.04292
R1548 VTAIL.n462 VTAIL.n461 4.26717
R1549 VTAIL.n492 VTAIL.n491 4.26717
R1550 VTAIL.n28 VTAIL.n27 4.26717
R1551 VTAIL.n58 VTAIL.n57 4.26717
R1552 VTAIL.n90 VTAIL.n89 4.26717
R1553 VTAIL.n120 VTAIL.n119 4.26717
R1554 VTAIL.n152 VTAIL.n151 4.26717
R1555 VTAIL.n182 VTAIL.n181 4.26717
R1556 VTAIL.n430 VTAIL.n429 4.26717
R1557 VTAIL.n402 VTAIL.n401 4.26717
R1558 VTAIL.n368 VTAIL.n367 4.26717
R1559 VTAIL.n340 VTAIL.n339 4.26717
R1560 VTAIL.n306 VTAIL.n305 4.26717
R1561 VTAIL.n278 VTAIL.n277 4.26717
R1562 VTAIL.n244 VTAIL.n243 4.26717
R1563 VTAIL.n216 VTAIL.n215 4.26717
R1564 VTAIL.n465 VTAIL.n448 3.49141
R1565 VTAIL.n488 VTAIL.n436 3.49141
R1566 VTAIL.n31 VTAIL.n14 3.49141
R1567 VTAIL.n54 VTAIL.n2 3.49141
R1568 VTAIL.n93 VTAIL.n76 3.49141
R1569 VTAIL.n116 VTAIL.n64 3.49141
R1570 VTAIL.n155 VTAIL.n138 3.49141
R1571 VTAIL.n178 VTAIL.n126 3.49141
R1572 VTAIL.n426 VTAIL.n374 3.49141
R1573 VTAIL.n405 VTAIL.n388 3.49141
R1574 VTAIL.n364 VTAIL.n312 3.49141
R1575 VTAIL.n343 VTAIL.n326 3.49141
R1576 VTAIL.n302 VTAIL.n250 3.49141
R1577 VTAIL.n281 VTAIL.n264 3.49141
R1578 VTAIL.n240 VTAIL.n188 3.49141
R1579 VTAIL.n219 VTAIL.n202 3.49141
R1580 VTAIL.n309 VTAIL.n247 2.72464
R1581 VTAIL.n433 VTAIL.n371 2.72464
R1582 VTAIL.n185 VTAIL.n123 2.72464
R1583 VTAIL.n466 VTAIL.n446 2.71565
R1584 VTAIL.n487 VTAIL.n438 2.71565
R1585 VTAIL.n32 VTAIL.n12 2.71565
R1586 VTAIL.n53 VTAIL.n4 2.71565
R1587 VTAIL.n94 VTAIL.n74 2.71565
R1588 VTAIL.n115 VTAIL.n66 2.71565
R1589 VTAIL.n156 VTAIL.n136 2.71565
R1590 VTAIL.n177 VTAIL.n128 2.71565
R1591 VTAIL.n425 VTAIL.n376 2.71565
R1592 VTAIL.n406 VTAIL.n386 2.71565
R1593 VTAIL.n363 VTAIL.n314 2.71565
R1594 VTAIL.n344 VTAIL.n324 2.71565
R1595 VTAIL.n301 VTAIL.n252 2.71565
R1596 VTAIL.n282 VTAIL.n262 2.71565
R1597 VTAIL.n239 VTAIL.n190 2.71565
R1598 VTAIL.n220 VTAIL.n200 2.71565
R1599 VTAIL.n453 VTAIL.n451 2.41282
R1600 VTAIL.n19 VTAIL.n17 2.41282
R1601 VTAIL.n81 VTAIL.n79 2.41282
R1602 VTAIL.n143 VTAIL.n141 2.41282
R1603 VTAIL.n393 VTAIL.n391 2.41282
R1604 VTAIL.n331 VTAIL.n329 2.41282
R1605 VTAIL.n269 VTAIL.n267 2.41282
R1606 VTAIL.n207 VTAIL.n205 2.41282
R1607 VTAIL.n471 VTAIL.n469 1.93989
R1608 VTAIL.n484 VTAIL.n483 1.93989
R1609 VTAIL.n37 VTAIL.n35 1.93989
R1610 VTAIL.n50 VTAIL.n49 1.93989
R1611 VTAIL.n99 VTAIL.n97 1.93989
R1612 VTAIL.n112 VTAIL.n111 1.93989
R1613 VTAIL.n161 VTAIL.n159 1.93989
R1614 VTAIL.n174 VTAIL.n173 1.93989
R1615 VTAIL.n422 VTAIL.n421 1.93989
R1616 VTAIL.n410 VTAIL.n409 1.93989
R1617 VTAIL.n360 VTAIL.n359 1.93989
R1618 VTAIL.n348 VTAIL.n347 1.93989
R1619 VTAIL.n298 VTAIL.n297 1.93989
R1620 VTAIL.n286 VTAIL.n285 1.93989
R1621 VTAIL.n236 VTAIL.n235 1.93989
R1622 VTAIL.n224 VTAIL.n223 1.93989
R1623 VTAIL VTAIL.n61 1.42076
R1624 VTAIL VTAIL.n495 1.30438
R1625 VTAIL.n470 VTAIL.n444 1.16414
R1626 VTAIL.n480 VTAIL.n440 1.16414
R1627 VTAIL.n36 VTAIL.n10 1.16414
R1628 VTAIL.n46 VTAIL.n6 1.16414
R1629 VTAIL.n98 VTAIL.n72 1.16414
R1630 VTAIL.n108 VTAIL.n68 1.16414
R1631 VTAIL.n160 VTAIL.n134 1.16414
R1632 VTAIL.n170 VTAIL.n130 1.16414
R1633 VTAIL.n418 VTAIL.n378 1.16414
R1634 VTAIL.n413 VTAIL.n383 1.16414
R1635 VTAIL.n356 VTAIL.n316 1.16414
R1636 VTAIL.n351 VTAIL.n321 1.16414
R1637 VTAIL.n294 VTAIL.n254 1.16414
R1638 VTAIL.n289 VTAIL.n259 1.16414
R1639 VTAIL.n232 VTAIL.n192 1.16414
R1640 VTAIL.n227 VTAIL.n197 1.16414
R1641 VTAIL.n371 VTAIL.n309 0.470328
R1642 VTAIL.n123 VTAIL.n61 0.470328
R1643 VTAIL.n476 VTAIL.n475 0.388379
R1644 VTAIL.n479 VTAIL.n442 0.388379
R1645 VTAIL.n42 VTAIL.n41 0.388379
R1646 VTAIL.n45 VTAIL.n8 0.388379
R1647 VTAIL.n104 VTAIL.n103 0.388379
R1648 VTAIL.n107 VTAIL.n70 0.388379
R1649 VTAIL.n166 VTAIL.n165 0.388379
R1650 VTAIL.n169 VTAIL.n132 0.388379
R1651 VTAIL.n417 VTAIL.n380 0.388379
R1652 VTAIL.n414 VTAIL.n382 0.388379
R1653 VTAIL.n355 VTAIL.n318 0.388379
R1654 VTAIL.n352 VTAIL.n320 0.388379
R1655 VTAIL.n293 VTAIL.n256 0.388379
R1656 VTAIL.n290 VTAIL.n258 0.388379
R1657 VTAIL.n231 VTAIL.n194 0.388379
R1658 VTAIL.n228 VTAIL.n196 0.388379
R1659 VTAIL.n459 VTAIL.n451 0.155672
R1660 VTAIL.n460 VTAIL.n459 0.155672
R1661 VTAIL.n460 VTAIL.n447 0.155672
R1662 VTAIL.n467 VTAIL.n447 0.155672
R1663 VTAIL.n468 VTAIL.n467 0.155672
R1664 VTAIL.n468 VTAIL.n443 0.155672
R1665 VTAIL.n477 VTAIL.n443 0.155672
R1666 VTAIL.n478 VTAIL.n477 0.155672
R1667 VTAIL.n478 VTAIL.n439 0.155672
R1668 VTAIL.n485 VTAIL.n439 0.155672
R1669 VTAIL.n486 VTAIL.n485 0.155672
R1670 VTAIL.n486 VTAIL.n435 0.155672
R1671 VTAIL.n493 VTAIL.n435 0.155672
R1672 VTAIL.n25 VTAIL.n17 0.155672
R1673 VTAIL.n26 VTAIL.n25 0.155672
R1674 VTAIL.n26 VTAIL.n13 0.155672
R1675 VTAIL.n33 VTAIL.n13 0.155672
R1676 VTAIL.n34 VTAIL.n33 0.155672
R1677 VTAIL.n34 VTAIL.n9 0.155672
R1678 VTAIL.n43 VTAIL.n9 0.155672
R1679 VTAIL.n44 VTAIL.n43 0.155672
R1680 VTAIL.n44 VTAIL.n5 0.155672
R1681 VTAIL.n51 VTAIL.n5 0.155672
R1682 VTAIL.n52 VTAIL.n51 0.155672
R1683 VTAIL.n52 VTAIL.n1 0.155672
R1684 VTAIL.n59 VTAIL.n1 0.155672
R1685 VTAIL.n87 VTAIL.n79 0.155672
R1686 VTAIL.n88 VTAIL.n87 0.155672
R1687 VTAIL.n88 VTAIL.n75 0.155672
R1688 VTAIL.n95 VTAIL.n75 0.155672
R1689 VTAIL.n96 VTAIL.n95 0.155672
R1690 VTAIL.n96 VTAIL.n71 0.155672
R1691 VTAIL.n105 VTAIL.n71 0.155672
R1692 VTAIL.n106 VTAIL.n105 0.155672
R1693 VTAIL.n106 VTAIL.n67 0.155672
R1694 VTAIL.n113 VTAIL.n67 0.155672
R1695 VTAIL.n114 VTAIL.n113 0.155672
R1696 VTAIL.n114 VTAIL.n63 0.155672
R1697 VTAIL.n121 VTAIL.n63 0.155672
R1698 VTAIL.n149 VTAIL.n141 0.155672
R1699 VTAIL.n150 VTAIL.n149 0.155672
R1700 VTAIL.n150 VTAIL.n137 0.155672
R1701 VTAIL.n157 VTAIL.n137 0.155672
R1702 VTAIL.n158 VTAIL.n157 0.155672
R1703 VTAIL.n158 VTAIL.n133 0.155672
R1704 VTAIL.n167 VTAIL.n133 0.155672
R1705 VTAIL.n168 VTAIL.n167 0.155672
R1706 VTAIL.n168 VTAIL.n129 0.155672
R1707 VTAIL.n175 VTAIL.n129 0.155672
R1708 VTAIL.n176 VTAIL.n175 0.155672
R1709 VTAIL.n176 VTAIL.n125 0.155672
R1710 VTAIL.n183 VTAIL.n125 0.155672
R1711 VTAIL.n431 VTAIL.n373 0.155672
R1712 VTAIL.n424 VTAIL.n373 0.155672
R1713 VTAIL.n424 VTAIL.n423 0.155672
R1714 VTAIL.n423 VTAIL.n377 0.155672
R1715 VTAIL.n416 VTAIL.n377 0.155672
R1716 VTAIL.n416 VTAIL.n415 0.155672
R1717 VTAIL.n415 VTAIL.n381 0.155672
R1718 VTAIL.n408 VTAIL.n381 0.155672
R1719 VTAIL.n408 VTAIL.n407 0.155672
R1720 VTAIL.n407 VTAIL.n387 0.155672
R1721 VTAIL.n400 VTAIL.n387 0.155672
R1722 VTAIL.n400 VTAIL.n399 0.155672
R1723 VTAIL.n399 VTAIL.n391 0.155672
R1724 VTAIL.n369 VTAIL.n311 0.155672
R1725 VTAIL.n362 VTAIL.n311 0.155672
R1726 VTAIL.n362 VTAIL.n361 0.155672
R1727 VTAIL.n361 VTAIL.n315 0.155672
R1728 VTAIL.n354 VTAIL.n315 0.155672
R1729 VTAIL.n354 VTAIL.n353 0.155672
R1730 VTAIL.n353 VTAIL.n319 0.155672
R1731 VTAIL.n346 VTAIL.n319 0.155672
R1732 VTAIL.n346 VTAIL.n345 0.155672
R1733 VTAIL.n345 VTAIL.n325 0.155672
R1734 VTAIL.n338 VTAIL.n325 0.155672
R1735 VTAIL.n338 VTAIL.n337 0.155672
R1736 VTAIL.n337 VTAIL.n329 0.155672
R1737 VTAIL.n307 VTAIL.n249 0.155672
R1738 VTAIL.n300 VTAIL.n249 0.155672
R1739 VTAIL.n300 VTAIL.n299 0.155672
R1740 VTAIL.n299 VTAIL.n253 0.155672
R1741 VTAIL.n292 VTAIL.n253 0.155672
R1742 VTAIL.n292 VTAIL.n291 0.155672
R1743 VTAIL.n291 VTAIL.n257 0.155672
R1744 VTAIL.n284 VTAIL.n257 0.155672
R1745 VTAIL.n284 VTAIL.n283 0.155672
R1746 VTAIL.n283 VTAIL.n263 0.155672
R1747 VTAIL.n276 VTAIL.n263 0.155672
R1748 VTAIL.n276 VTAIL.n275 0.155672
R1749 VTAIL.n275 VTAIL.n267 0.155672
R1750 VTAIL.n245 VTAIL.n187 0.155672
R1751 VTAIL.n238 VTAIL.n187 0.155672
R1752 VTAIL.n238 VTAIL.n237 0.155672
R1753 VTAIL.n237 VTAIL.n191 0.155672
R1754 VTAIL.n230 VTAIL.n191 0.155672
R1755 VTAIL.n230 VTAIL.n229 0.155672
R1756 VTAIL.n229 VTAIL.n195 0.155672
R1757 VTAIL.n222 VTAIL.n195 0.155672
R1758 VTAIL.n222 VTAIL.n221 0.155672
R1759 VTAIL.n221 VTAIL.n201 0.155672
R1760 VTAIL.n214 VTAIL.n201 0.155672
R1761 VTAIL.n214 VTAIL.n213 0.155672
R1762 VTAIL.n213 VTAIL.n205 0.155672
R1763 VP.n16 VP.n0 161.3
R1764 VP.n15 VP.n14 161.3
R1765 VP.n13 VP.n1 161.3
R1766 VP.n12 VP.n11 161.3
R1767 VP.n10 VP.n2 161.3
R1768 VP.n9 VP.n8 161.3
R1769 VP.n7 VP.n3 161.3
R1770 VP.n4 VP.t1 131.362
R1771 VP.n4 VP.t0 130.466
R1772 VP.n6 VP.n5 106.974
R1773 VP.n18 VP.n17 106.974
R1774 VP.n5 VP.t3 96.0599
R1775 VP.n17 VP.t2 96.0599
R1776 VP.n6 VP.n4 49.9207
R1777 VP.n11 VP.n10 40.577
R1778 VP.n11 VP.n1 40.577
R1779 VP.n9 VP.n3 24.5923
R1780 VP.n10 VP.n9 24.5923
R1781 VP.n15 VP.n1 24.5923
R1782 VP.n16 VP.n15 24.5923
R1783 VP.n5 VP.n3 3.93519
R1784 VP.n17 VP.n16 3.93519
R1785 VP.n7 VP.n6 0.278335
R1786 VP.n18 VP.n0 0.278335
R1787 VP.n8 VP.n7 0.189894
R1788 VP.n8 VP.n2 0.189894
R1789 VP.n12 VP.n2 0.189894
R1790 VP.n13 VP.n12 0.189894
R1791 VP.n14 VP.n13 0.189894
R1792 VP.n14 VP.n0 0.189894
R1793 VP VP.n18 0.153485
R1794 VDD1 VDD1.n1 114.591
R1795 VDD1 VDD1.n0 72.5137
R1796 VDD1.n0 VDD1.t2 2.88215
R1797 VDD1.n0 VDD1.t3 2.88215
R1798 VDD1.n1 VDD1.t0 2.88215
R1799 VDD1.n1 VDD1.t1 2.88215
C0 VDD2 w_n2866_n3224# 1.53625f
C1 w_n2866_n3224# VP 5.24585f
C2 w_n2866_n3224# VN 4.87683f
C3 w_n2866_n3224# B 9.32702f
C4 VTAIL VDD1 5.2841f
C5 VDD2 VDD1 1.07745f
C6 VDD1 VP 4.81337f
C7 VN VDD1 0.14938f
C8 VDD2 VTAIL 5.33985f
C9 VTAIL VP 4.54137f
C10 B VDD1 1.28232f
C11 VN VTAIL 4.52726f
C12 VDD2 VP 0.409113f
C13 VDD2 VN 4.55443f
C14 VN VP 6.21827f
C15 w_n2866_n3224# VDD1 1.47503f
C16 VTAIL B 4.80827f
C17 VDD2 B 1.33829f
C18 B VP 1.76132f
C19 VN B 1.14788f
C20 w_n2866_n3224# VTAIL 3.81986f
C21 VDD2 VSUBS 0.970204f
C22 VDD1 VSUBS 5.78311f
C23 VTAIL VSUBS 1.207754f
C24 VN VSUBS 5.54626f
C25 VP VSUBS 2.371798f
C26 B VSUBS 4.413948f
C27 w_n2866_n3224# VSUBS 0.113872p
C28 VDD1.t2 VSUBS 0.243137f
C29 VDD1.t3 VSUBS 0.243137f
C30 VDD1.n0 VSUBS 1.86828f
C31 VDD1.t0 VSUBS 0.243137f
C32 VDD1.t1 VSUBS 0.243137f
C33 VDD1.n1 VSUBS 2.60746f
C34 VP.n0 VSUBS 0.043473f
C35 VP.t2 VSUBS 2.86291f
C36 VP.n1 VSUBS 0.065194f
C37 VP.n2 VSUBS 0.032976f
C38 VP.n3 VSUBS 0.035792f
C39 VP.t0 VSUBS 3.18844f
C40 VP.t1 VSUBS 3.19662f
C41 VP.n4 VSUBS 3.82139f
C42 VP.t3 VSUBS 2.86291f
C43 VP.n5 VSUBS 1.12252f
C44 VP.n6 VSUBS 1.81646f
C45 VP.n7 VSUBS 0.043473f
C46 VP.n8 VSUBS 0.032976f
C47 VP.n9 VSUBS 0.061151f
C48 VP.n10 VSUBS 0.065194f
C49 VP.n11 VSUBS 0.026634f
C50 VP.n12 VSUBS 0.032976f
C51 VP.n13 VSUBS 0.032976f
C52 VP.n14 VSUBS 0.032976f
C53 VP.n15 VSUBS 0.061151f
C54 VP.n16 VSUBS 0.035792f
C55 VP.n17 VSUBS 1.12252f
C56 VP.n18 VSUBS 0.061113f
C57 VTAIL.n0 VSUBS 0.024673f
C58 VTAIL.n1 VSUBS 0.02403f
C59 VTAIL.n2 VSUBS 0.012913f
C60 VTAIL.n3 VSUBS 0.03052f
C61 VTAIL.n4 VSUBS 0.013672f
C62 VTAIL.n5 VSUBS 0.02403f
C63 VTAIL.n6 VSUBS 0.012913f
C64 VTAIL.n7 VSUBS 0.03052f
C65 VTAIL.n8 VSUBS 0.013292f
C66 VTAIL.n9 VSUBS 0.02403f
C67 VTAIL.n10 VSUBS 0.013672f
C68 VTAIL.n11 VSUBS 0.03052f
C69 VTAIL.n12 VSUBS 0.013672f
C70 VTAIL.n13 VSUBS 0.02403f
C71 VTAIL.n14 VSUBS 0.012913f
C72 VTAIL.n15 VSUBS 0.03052f
C73 VTAIL.n16 VSUBS 0.013672f
C74 VTAIL.n17 VSUBS 1.10484f
C75 VTAIL.n18 VSUBS 0.012913f
C76 VTAIL.t3 VSUBS 0.06571f
C77 VTAIL.n19 VSUBS 0.181425f
C78 VTAIL.n20 VSUBS 0.022959f
C79 VTAIL.n21 VSUBS 0.02289f
C80 VTAIL.n22 VSUBS 0.03052f
C81 VTAIL.n23 VSUBS 0.013672f
C82 VTAIL.n24 VSUBS 0.012913f
C83 VTAIL.n25 VSUBS 0.02403f
C84 VTAIL.n26 VSUBS 0.02403f
C85 VTAIL.n27 VSUBS 0.012913f
C86 VTAIL.n28 VSUBS 0.013672f
C87 VTAIL.n29 VSUBS 0.03052f
C88 VTAIL.n30 VSUBS 0.03052f
C89 VTAIL.n31 VSUBS 0.013672f
C90 VTAIL.n32 VSUBS 0.012913f
C91 VTAIL.n33 VSUBS 0.02403f
C92 VTAIL.n34 VSUBS 0.02403f
C93 VTAIL.n35 VSUBS 0.012913f
C94 VTAIL.n36 VSUBS 0.012913f
C95 VTAIL.n37 VSUBS 0.013672f
C96 VTAIL.n38 VSUBS 0.03052f
C97 VTAIL.n39 VSUBS 0.03052f
C98 VTAIL.n40 VSUBS 0.03052f
C99 VTAIL.n41 VSUBS 0.013292f
C100 VTAIL.n42 VSUBS 0.012913f
C101 VTAIL.n43 VSUBS 0.02403f
C102 VTAIL.n44 VSUBS 0.02403f
C103 VTAIL.n45 VSUBS 0.012913f
C104 VTAIL.n46 VSUBS 0.013672f
C105 VTAIL.n47 VSUBS 0.03052f
C106 VTAIL.n48 VSUBS 0.03052f
C107 VTAIL.n49 VSUBS 0.013672f
C108 VTAIL.n50 VSUBS 0.012913f
C109 VTAIL.n51 VSUBS 0.02403f
C110 VTAIL.n52 VSUBS 0.02403f
C111 VTAIL.n53 VSUBS 0.012913f
C112 VTAIL.n54 VSUBS 0.013672f
C113 VTAIL.n55 VSUBS 0.03052f
C114 VTAIL.n56 VSUBS 0.067993f
C115 VTAIL.n57 VSUBS 0.013672f
C116 VTAIL.n58 VSUBS 0.012913f
C117 VTAIL.n59 VSUBS 0.051604f
C118 VTAIL.n60 VSUBS 0.033806f
C119 VTAIL.n61 VSUBS 0.164651f
C120 VTAIL.n62 VSUBS 0.024673f
C121 VTAIL.n63 VSUBS 0.02403f
C122 VTAIL.n64 VSUBS 0.012913f
C123 VTAIL.n65 VSUBS 0.03052f
C124 VTAIL.n66 VSUBS 0.013672f
C125 VTAIL.n67 VSUBS 0.02403f
C126 VTAIL.n68 VSUBS 0.012913f
C127 VTAIL.n69 VSUBS 0.03052f
C128 VTAIL.n70 VSUBS 0.013292f
C129 VTAIL.n71 VSUBS 0.02403f
C130 VTAIL.n72 VSUBS 0.013672f
C131 VTAIL.n73 VSUBS 0.03052f
C132 VTAIL.n74 VSUBS 0.013672f
C133 VTAIL.n75 VSUBS 0.02403f
C134 VTAIL.n76 VSUBS 0.012913f
C135 VTAIL.n77 VSUBS 0.03052f
C136 VTAIL.n78 VSUBS 0.013672f
C137 VTAIL.n79 VSUBS 1.10484f
C138 VTAIL.n80 VSUBS 0.012913f
C139 VTAIL.t6 VSUBS 0.06571f
C140 VTAIL.n81 VSUBS 0.181425f
C141 VTAIL.n82 VSUBS 0.022959f
C142 VTAIL.n83 VSUBS 0.02289f
C143 VTAIL.n84 VSUBS 0.03052f
C144 VTAIL.n85 VSUBS 0.013672f
C145 VTAIL.n86 VSUBS 0.012913f
C146 VTAIL.n87 VSUBS 0.02403f
C147 VTAIL.n88 VSUBS 0.02403f
C148 VTAIL.n89 VSUBS 0.012913f
C149 VTAIL.n90 VSUBS 0.013672f
C150 VTAIL.n91 VSUBS 0.03052f
C151 VTAIL.n92 VSUBS 0.03052f
C152 VTAIL.n93 VSUBS 0.013672f
C153 VTAIL.n94 VSUBS 0.012913f
C154 VTAIL.n95 VSUBS 0.02403f
C155 VTAIL.n96 VSUBS 0.02403f
C156 VTAIL.n97 VSUBS 0.012913f
C157 VTAIL.n98 VSUBS 0.012913f
C158 VTAIL.n99 VSUBS 0.013672f
C159 VTAIL.n100 VSUBS 0.03052f
C160 VTAIL.n101 VSUBS 0.03052f
C161 VTAIL.n102 VSUBS 0.03052f
C162 VTAIL.n103 VSUBS 0.013292f
C163 VTAIL.n104 VSUBS 0.012913f
C164 VTAIL.n105 VSUBS 0.02403f
C165 VTAIL.n106 VSUBS 0.02403f
C166 VTAIL.n107 VSUBS 0.012913f
C167 VTAIL.n108 VSUBS 0.013672f
C168 VTAIL.n109 VSUBS 0.03052f
C169 VTAIL.n110 VSUBS 0.03052f
C170 VTAIL.n111 VSUBS 0.013672f
C171 VTAIL.n112 VSUBS 0.012913f
C172 VTAIL.n113 VSUBS 0.02403f
C173 VTAIL.n114 VSUBS 0.02403f
C174 VTAIL.n115 VSUBS 0.012913f
C175 VTAIL.n116 VSUBS 0.013672f
C176 VTAIL.n117 VSUBS 0.03052f
C177 VTAIL.n118 VSUBS 0.067993f
C178 VTAIL.n119 VSUBS 0.013672f
C179 VTAIL.n120 VSUBS 0.012913f
C180 VTAIL.n121 VSUBS 0.051604f
C181 VTAIL.n122 VSUBS 0.033806f
C182 VTAIL.n123 VSUBS 0.265609f
C183 VTAIL.n124 VSUBS 0.024673f
C184 VTAIL.n125 VSUBS 0.02403f
C185 VTAIL.n126 VSUBS 0.012913f
C186 VTAIL.n127 VSUBS 0.03052f
C187 VTAIL.n128 VSUBS 0.013672f
C188 VTAIL.n129 VSUBS 0.02403f
C189 VTAIL.n130 VSUBS 0.012913f
C190 VTAIL.n131 VSUBS 0.03052f
C191 VTAIL.n132 VSUBS 0.013292f
C192 VTAIL.n133 VSUBS 0.02403f
C193 VTAIL.n134 VSUBS 0.013672f
C194 VTAIL.n135 VSUBS 0.03052f
C195 VTAIL.n136 VSUBS 0.013672f
C196 VTAIL.n137 VSUBS 0.02403f
C197 VTAIL.n138 VSUBS 0.012913f
C198 VTAIL.n139 VSUBS 0.03052f
C199 VTAIL.n140 VSUBS 0.013672f
C200 VTAIL.n141 VSUBS 1.10484f
C201 VTAIL.n142 VSUBS 0.012913f
C202 VTAIL.t1 VSUBS 0.06571f
C203 VTAIL.n143 VSUBS 0.181425f
C204 VTAIL.n144 VSUBS 0.022959f
C205 VTAIL.n145 VSUBS 0.02289f
C206 VTAIL.n146 VSUBS 0.03052f
C207 VTAIL.n147 VSUBS 0.013672f
C208 VTAIL.n148 VSUBS 0.012913f
C209 VTAIL.n149 VSUBS 0.02403f
C210 VTAIL.n150 VSUBS 0.02403f
C211 VTAIL.n151 VSUBS 0.012913f
C212 VTAIL.n152 VSUBS 0.013672f
C213 VTAIL.n153 VSUBS 0.03052f
C214 VTAIL.n154 VSUBS 0.03052f
C215 VTAIL.n155 VSUBS 0.013672f
C216 VTAIL.n156 VSUBS 0.012913f
C217 VTAIL.n157 VSUBS 0.02403f
C218 VTAIL.n158 VSUBS 0.02403f
C219 VTAIL.n159 VSUBS 0.012913f
C220 VTAIL.n160 VSUBS 0.012913f
C221 VTAIL.n161 VSUBS 0.013672f
C222 VTAIL.n162 VSUBS 0.03052f
C223 VTAIL.n163 VSUBS 0.03052f
C224 VTAIL.n164 VSUBS 0.03052f
C225 VTAIL.n165 VSUBS 0.013292f
C226 VTAIL.n166 VSUBS 0.012913f
C227 VTAIL.n167 VSUBS 0.02403f
C228 VTAIL.n168 VSUBS 0.02403f
C229 VTAIL.n169 VSUBS 0.012913f
C230 VTAIL.n170 VSUBS 0.013672f
C231 VTAIL.n171 VSUBS 0.03052f
C232 VTAIL.n172 VSUBS 0.03052f
C233 VTAIL.n173 VSUBS 0.013672f
C234 VTAIL.n174 VSUBS 0.012913f
C235 VTAIL.n175 VSUBS 0.02403f
C236 VTAIL.n176 VSUBS 0.02403f
C237 VTAIL.n177 VSUBS 0.012913f
C238 VTAIL.n178 VSUBS 0.013672f
C239 VTAIL.n179 VSUBS 0.03052f
C240 VTAIL.n180 VSUBS 0.067993f
C241 VTAIL.n181 VSUBS 0.013672f
C242 VTAIL.n182 VSUBS 0.012913f
C243 VTAIL.n183 VSUBS 0.051604f
C244 VTAIL.n184 VSUBS 0.033806f
C245 VTAIL.n185 VSUBS 1.5195f
C246 VTAIL.n186 VSUBS 0.024673f
C247 VTAIL.n187 VSUBS 0.02403f
C248 VTAIL.n188 VSUBS 0.012913f
C249 VTAIL.n189 VSUBS 0.03052f
C250 VTAIL.n190 VSUBS 0.013672f
C251 VTAIL.n191 VSUBS 0.02403f
C252 VTAIL.n192 VSUBS 0.012913f
C253 VTAIL.n193 VSUBS 0.03052f
C254 VTAIL.n194 VSUBS 0.013292f
C255 VTAIL.n195 VSUBS 0.02403f
C256 VTAIL.n196 VSUBS 0.013292f
C257 VTAIL.n197 VSUBS 0.012913f
C258 VTAIL.n198 VSUBS 0.03052f
C259 VTAIL.n199 VSUBS 0.03052f
C260 VTAIL.n200 VSUBS 0.013672f
C261 VTAIL.n201 VSUBS 0.02403f
C262 VTAIL.n202 VSUBS 0.012913f
C263 VTAIL.n203 VSUBS 0.03052f
C264 VTAIL.n204 VSUBS 0.013672f
C265 VTAIL.n205 VSUBS 1.10484f
C266 VTAIL.n206 VSUBS 0.012913f
C267 VTAIL.t5 VSUBS 0.06571f
C268 VTAIL.n207 VSUBS 0.181425f
C269 VTAIL.n208 VSUBS 0.022959f
C270 VTAIL.n209 VSUBS 0.02289f
C271 VTAIL.n210 VSUBS 0.03052f
C272 VTAIL.n211 VSUBS 0.013672f
C273 VTAIL.n212 VSUBS 0.012913f
C274 VTAIL.n213 VSUBS 0.02403f
C275 VTAIL.n214 VSUBS 0.02403f
C276 VTAIL.n215 VSUBS 0.012913f
C277 VTAIL.n216 VSUBS 0.013672f
C278 VTAIL.n217 VSUBS 0.03052f
C279 VTAIL.n218 VSUBS 0.03052f
C280 VTAIL.n219 VSUBS 0.013672f
C281 VTAIL.n220 VSUBS 0.012913f
C282 VTAIL.n221 VSUBS 0.02403f
C283 VTAIL.n222 VSUBS 0.02403f
C284 VTAIL.n223 VSUBS 0.012913f
C285 VTAIL.n224 VSUBS 0.013672f
C286 VTAIL.n225 VSUBS 0.03052f
C287 VTAIL.n226 VSUBS 0.03052f
C288 VTAIL.n227 VSUBS 0.013672f
C289 VTAIL.n228 VSUBS 0.012913f
C290 VTAIL.n229 VSUBS 0.02403f
C291 VTAIL.n230 VSUBS 0.02403f
C292 VTAIL.n231 VSUBS 0.012913f
C293 VTAIL.n232 VSUBS 0.013672f
C294 VTAIL.n233 VSUBS 0.03052f
C295 VTAIL.n234 VSUBS 0.03052f
C296 VTAIL.n235 VSUBS 0.013672f
C297 VTAIL.n236 VSUBS 0.012913f
C298 VTAIL.n237 VSUBS 0.02403f
C299 VTAIL.n238 VSUBS 0.02403f
C300 VTAIL.n239 VSUBS 0.012913f
C301 VTAIL.n240 VSUBS 0.013672f
C302 VTAIL.n241 VSUBS 0.03052f
C303 VTAIL.n242 VSUBS 0.067993f
C304 VTAIL.n243 VSUBS 0.013672f
C305 VTAIL.n244 VSUBS 0.012913f
C306 VTAIL.n245 VSUBS 0.051604f
C307 VTAIL.n246 VSUBS 0.033806f
C308 VTAIL.n247 VSUBS 1.5195f
C309 VTAIL.n248 VSUBS 0.024673f
C310 VTAIL.n249 VSUBS 0.02403f
C311 VTAIL.n250 VSUBS 0.012913f
C312 VTAIL.n251 VSUBS 0.03052f
C313 VTAIL.n252 VSUBS 0.013672f
C314 VTAIL.n253 VSUBS 0.02403f
C315 VTAIL.n254 VSUBS 0.012913f
C316 VTAIL.n255 VSUBS 0.03052f
C317 VTAIL.n256 VSUBS 0.013292f
C318 VTAIL.n257 VSUBS 0.02403f
C319 VTAIL.n258 VSUBS 0.013292f
C320 VTAIL.n259 VSUBS 0.012913f
C321 VTAIL.n260 VSUBS 0.03052f
C322 VTAIL.n261 VSUBS 0.03052f
C323 VTAIL.n262 VSUBS 0.013672f
C324 VTAIL.n263 VSUBS 0.02403f
C325 VTAIL.n264 VSUBS 0.012913f
C326 VTAIL.n265 VSUBS 0.03052f
C327 VTAIL.n266 VSUBS 0.013672f
C328 VTAIL.n267 VSUBS 1.10484f
C329 VTAIL.n268 VSUBS 0.012913f
C330 VTAIL.t4 VSUBS 0.06571f
C331 VTAIL.n269 VSUBS 0.181425f
C332 VTAIL.n270 VSUBS 0.022959f
C333 VTAIL.n271 VSUBS 0.02289f
C334 VTAIL.n272 VSUBS 0.03052f
C335 VTAIL.n273 VSUBS 0.013672f
C336 VTAIL.n274 VSUBS 0.012913f
C337 VTAIL.n275 VSUBS 0.02403f
C338 VTAIL.n276 VSUBS 0.02403f
C339 VTAIL.n277 VSUBS 0.012913f
C340 VTAIL.n278 VSUBS 0.013672f
C341 VTAIL.n279 VSUBS 0.03052f
C342 VTAIL.n280 VSUBS 0.03052f
C343 VTAIL.n281 VSUBS 0.013672f
C344 VTAIL.n282 VSUBS 0.012913f
C345 VTAIL.n283 VSUBS 0.02403f
C346 VTAIL.n284 VSUBS 0.02403f
C347 VTAIL.n285 VSUBS 0.012913f
C348 VTAIL.n286 VSUBS 0.013672f
C349 VTAIL.n287 VSUBS 0.03052f
C350 VTAIL.n288 VSUBS 0.03052f
C351 VTAIL.n289 VSUBS 0.013672f
C352 VTAIL.n290 VSUBS 0.012913f
C353 VTAIL.n291 VSUBS 0.02403f
C354 VTAIL.n292 VSUBS 0.02403f
C355 VTAIL.n293 VSUBS 0.012913f
C356 VTAIL.n294 VSUBS 0.013672f
C357 VTAIL.n295 VSUBS 0.03052f
C358 VTAIL.n296 VSUBS 0.03052f
C359 VTAIL.n297 VSUBS 0.013672f
C360 VTAIL.n298 VSUBS 0.012913f
C361 VTAIL.n299 VSUBS 0.02403f
C362 VTAIL.n300 VSUBS 0.02403f
C363 VTAIL.n301 VSUBS 0.012913f
C364 VTAIL.n302 VSUBS 0.013672f
C365 VTAIL.n303 VSUBS 0.03052f
C366 VTAIL.n304 VSUBS 0.067993f
C367 VTAIL.n305 VSUBS 0.013672f
C368 VTAIL.n306 VSUBS 0.012913f
C369 VTAIL.n307 VSUBS 0.051604f
C370 VTAIL.n308 VSUBS 0.033806f
C371 VTAIL.n309 VSUBS 0.265609f
C372 VTAIL.n310 VSUBS 0.024673f
C373 VTAIL.n311 VSUBS 0.02403f
C374 VTAIL.n312 VSUBS 0.012913f
C375 VTAIL.n313 VSUBS 0.03052f
C376 VTAIL.n314 VSUBS 0.013672f
C377 VTAIL.n315 VSUBS 0.02403f
C378 VTAIL.n316 VSUBS 0.012913f
C379 VTAIL.n317 VSUBS 0.03052f
C380 VTAIL.n318 VSUBS 0.013292f
C381 VTAIL.n319 VSUBS 0.02403f
C382 VTAIL.n320 VSUBS 0.013292f
C383 VTAIL.n321 VSUBS 0.012913f
C384 VTAIL.n322 VSUBS 0.03052f
C385 VTAIL.n323 VSUBS 0.03052f
C386 VTAIL.n324 VSUBS 0.013672f
C387 VTAIL.n325 VSUBS 0.02403f
C388 VTAIL.n326 VSUBS 0.012913f
C389 VTAIL.n327 VSUBS 0.03052f
C390 VTAIL.n328 VSUBS 0.013672f
C391 VTAIL.n329 VSUBS 1.10484f
C392 VTAIL.n330 VSUBS 0.012913f
C393 VTAIL.t7 VSUBS 0.06571f
C394 VTAIL.n331 VSUBS 0.181425f
C395 VTAIL.n332 VSUBS 0.022959f
C396 VTAIL.n333 VSUBS 0.02289f
C397 VTAIL.n334 VSUBS 0.03052f
C398 VTAIL.n335 VSUBS 0.013672f
C399 VTAIL.n336 VSUBS 0.012913f
C400 VTAIL.n337 VSUBS 0.02403f
C401 VTAIL.n338 VSUBS 0.02403f
C402 VTAIL.n339 VSUBS 0.012913f
C403 VTAIL.n340 VSUBS 0.013672f
C404 VTAIL.n341 VSUBS 0.03052f
C405 VTAIL.n342 VSUBS 0.03052f
C406 VTAIL.n343 VSUBS 0.013672f
C407 VTAIL.n344 VSUBS 0.012913f
C408 VTAIL.n345 VSUBS 0.02403f
C409 VTAIL.n346 VSUBS 0.02403f
C410 VTAIL.n347 VSUBS 0.012913f
C411 VTAIL.n348 VSUBS 0.013672f
C412 VTAIL.n349 VSUBS 0.03052f
C413 VTAIL.n350 VSUBS 0.03052f
C414 VTAIL.n351 VSUBS 0.013672f
C415 VTAIL.n352 VSUBS 0.012913f
C416 VTAIL.n353 VSUBS 0.02403f
C417 VTAIL.n354 VSUBS 0.02403f
C418 VTAIL.n355 VSUBS 0.012913f
C419 VTAIL.n356 VSUBS 0.013672f
C420 VTAIL.n357 VSUBS 0.03052f
C421 VTAIL.n358 VSUBS 0.03052f
C422 VTAIL.n359 VSUBS 0.013672f
C423 VTAIL.n360 VSUBS 0.012913f
C424 VTAIL.n361 VSUBS 0.02403f
C425 VTAIL.n362 VSUBS 0.02403f
C426 VTAIL.n363 VSUBS 0.012913f
C427 VTAIL.n364 VSUBS 0.013672f
C428 VTAIL.n365 VSUBS 0.03052f
C429 VTAIL.n366 VSUBS 0.067993f
C430 VTAIL.n367 VSUBS 0.013672f
C431 VTAIL.n368 VSUBS 0.012913f
C432 VTAIL.n369 VSUBS 0.051604f
C433 VTAIL.n370 VSUBS 0.033806f
C434 VTAIL.n371 VSUBS 0.265609f
C435 VTAIL.n372 VSUBS 0.024673f
C436 VTAIL.n373 VSUBS 0.02403f
C437 VTAIL.n374 VSUBS 0.012913f
C438 VTAIL.n375 VSUBS 0.03052f
C439 VTAIL.n376 VSUBS 0.013672f
C440 VTAIL.n377 VSUBS 0.02403f
C441 VTAIL.n378 VSUBS 0.012913f
C442 VTAIL.n379 VSUBS 0.03052f
C443 VTAIL.n380 VSUBS 0.013292f
C444 VTAIL.n381 VSUBS 0.02403f
C445 VTAIL.n382 VSUBS 0.013292f
C446 VTAIL.n383 VSUBS 0.012913f
C447 VTAIL.n384 VSUBS 0.03052f
C448 VTAIL.n385 VSUBS 0.03052f
C449 VTAIL.n386 VSUBS 0.013672f
C450 VTAIL.n387 VSUBS 0.02403f
C451 VTAIL.n388 VSUBS 0.012913f
C452 VTAIL.n389 VSUBS 0.03052f
C453 VTAIL.n390 VSUBS 0.013672f
C454 VTAIL.n391 VSUBS 1.10484f
C455 VTAIL.n392 VSUBS 0.012913f
C456 VTAIL.t0 VSUBS 0.06571f
C457 VTAIL.n393 VSUBS 0.181425f
C458 VTAIL.n394 VSUBS 0.022959f
C459 VTAIL.n395 VSUBS 0.02289f
C460 VTAIL.n396 VSUBS 0.03052f
C461 VTAIL.n397 VSUBS 0.013672f
C462 VTAIL.n398 VSUBS 0.012913f
C463 VTAIL.n399 VSUBS 0.02403f
C464 VTAIL.n400 VSUBS 0.02403f
C465 VTAIL.n401 VSUBS 0.012913f
C466 VTAIL.n402 VSUBS 0.013672f
C467 VTAIL.n403 VSUBS 0.03052f
C468 VTAIL.n404 VSUBS 0.03052f
C469 VTAIL.n405 VSUBS 0.013672f
C470 VTAIL.n406 VSUBS 0.012913f
C471 VTAIL.n407 VSUBS 0.02403f
C472 VTAIL.n408 VSUBS 0.02403f
C473 VTAIL.n409 VSUBS 0.012913f
C474 VTAIL.n410 VSUBS 0.013672f
C475 VTAIL.n411 VSUBS 0.03052f
C476 VTAIL.n412 VSUBS 0.03052f
C477 VTAIL.n413 VSUBS 0.013672f
C478 VTAIL.n414 VSUBS 0.012913f
C479 VTAIL.n415 VSUBS 0.02403f
C480 VTAIL.n416 VSUBS 0.02403f
C481 VTAIL.n417 VSUBS 0.012913f
C482 VTAIL.n418 VSUBS 0.013672f
C483 VTAIL.n419 VSUBS 0.03052f
C484 VTAIL.n420 VSUBS 0.03052f
C485 VTAIL.n421 VSUBS 0.013672f
C486 VTAIL.n422 VSUBS 0.012913f
C487 VTAIL.n423 VSUBS 0.02403f
C488 VTAIL.n424 VSUBS 0.02403f
C489 VTAIL.n425 VSUBS 0.012913f
C490 VTAIL.n426 VSUBS 0.013672f
C491 VTAIL.n427 VSUBS 0.03052f
C492 VTAIL.n428 VSUBS 0.067993f
C493 VTAIL.n429 VSUBS 0.013672f
C494 VTAIL.n430 VSUBS 0.012913f
C495 VTAIL.n431 VSUBS 0.051604f
C496 VTAIL.n432 VSUBS 0.033806f
C497 VTAIL.n433 VSUBS 1.5195f
C498 VTAIL.n434 VSUBS 0.024673f
C499 VTAIL.n435 VSUBS 0.02403f
C500 VTAIL.n436 VSUBS 0.012913f
C501 VTAIL.n437 VSUBS 0.03052f
C502 VTAIL.n438 VSUBS 0.013672f
C503 VTAIL.n439 VSUBS 0.02403f
C504 VTAIL.n440 VSUBS 0.012913f
C505 VTAIL.n441 VSUBS 0.03052f
C506 VTAIL.n442 VSUBS 0.013292f
C507 VTAIL.n443 VSUBS 0.02403f
C508 VTAIL.n444 VSUBS 0.013672f
C509 VTAIL.n445 VSUBS 0.03052f
C510 VTAIL.n446 VSUBS 0.013672f
C511 VTAIL.n447 VSUBS 0.02403f
C512 VTAIL.n448 VSUBS 0.012913f
C513 VTAIL.n449 VSUBS 0.03052f
C514 VTAIL.n450 VSUBS 0.013672f
C515 VTAIL.n451 VSUBS 1.10484f
C516 VTAIL.n452 VSUBS 0.012913f
C517 VTAIL.t2 VSUBS 0.06571f
C518 VTAIL.n453 VSUBS 0.181425f
C519 VTAIL.n454 VSUBS 0.022959f
C520 VTAIL.n455 VSUBS 0.02289f
C521 VTAIL.n456 VSUBS 0.03052f
C522 VTAIL.n457 VSUBS 0.013672f
C523 VTAIL.n458 VSUBS 0.012913f
C524 VTAIL.n459 VSUBS 0.02403f
C525 VTAIL.n460 VSUBS 0.02403f
C526 VTAIL.n461 VSUBS 0.012913f
C527 VTAIL.n462 VSUBS 0.013672f
C528 VTAIL.n463 VSUBS 0.03052f
C529 VTAIL.n464 VSUBS 0.03052f
C530 VTAIL.n465 VSUBS 0.013672f
C531 VTAIL.n466 VSUBS 0.012913f
C532 VTAIL.n467 VSUBS 0.02403f
C533 VTAIL.n468 VSUBS 0.02403f
C534 VTAIL.n469 VSUBS 0.012913f
C535 VTAIL.n470 VSUBS 0.012913f
C536 VTAIL.n471 VSUBS 0.013672f
C537 VTAIL.n472 VSUBS 0.03052f
C538 VTAIL.n473 VSUBS 0.03052f
C539 VTAIL.n474 VSUBS 0.03052f
C540 VTAIL.n475 VSUBS 0.013292f
C541 VTAIL.n476 VSUBS 0.012913f
C542 VTAIL.n477 VSUBS 0.02403f
C543 VTAIL.n478 VSUBS 0.02403f
C544 VTAIL.n479 VSUBS 0.012913f
C545 VTAIL.n480 VSUBS 0.013672f
C546 VTAIL.n481 VSUBS 0.03052f
C547 VTAIL.n482 VSUBS 0.03052f
C548 VTAIL.n483 VSUBS 0.013672f
C549 VTAIL.n484 VSUBS 0.012913f
C550 VTAIL.n485 VSUBS 0.02403f
C551 VTAIL.n486 VSUBS 0.02403f
C552 VTAIL.n487 VSUBS 0.012913f
C553 VTAIL.n488 VSUBS 0.013672f
C554 VTAIL.n489 VSUBS 0.03052f
C555 VTAIL.n490 VSUBS 0.067993f
C556 VTAIL.n491 VSUBS 0.013672f
C557 VTAIL.n492 VSUBS 0.012913f
C558 VTAIL.n493 VSUBS 0.051604f
C559 VTAIL.n494 VSUBS 0.033806f
C560 VTAIL.n495 VSUBS 1.40953f
C561 VDD2.t3 VSUBS 0.240723f
C562 VDD2.t2 VSUBS 0.240723f
C563 VDD2.n0 VSUBS 2.55619f
C564 VDD2.t0 VSUBS 0.240723f
C565 VDD2.t1 VSUBS 0.240723f
C566 VDD2.n1 VSUBS 1.84912f
C567 VDD2.n2 VSUBS 4.28893f
C568 VN.t2 VSUBS 3.11244f
C569 VN.t3 VSUBS 3.10447f
C570 VN.n0 VSUBS 1.93781f
C571 VN.t1 VSUBS 3.11244f
C572 VN.t0 VSUBS 3.10447f
C573 VN.n1 VSUBS 3.73776f
C574 B.n0 VSUBS 0.004235f
C575 B.n1 VSUBS 0.004235f
C576 B.n2 VSUBS 0.006697f
C577 B.n3 VSUBS 0.006697f
C578 B.n4 VSUBS 0.006697f
C579 B.n5 VSUBS 0.006697f
C580 B.n6 VSUBS 0.006697f
C581 B.n7 VSUBS 0.006697f
C582 B.n8 VSUBS 0.006697f
C583 B.n9 VSUBS 0.006697f
C584 B.n10 VSUBS 0.006697f
C585 B.n11 VSUBS 0.006697f
C586 B.n12 VSUBS 0.006697f
C587 B.n13 VSUBS 0.006697f
C588 B.n14 VSUBS 0.006697f
C589 B.n15 VSUBS 0.006697f
C590 B.n16 VSUBS 0.006697f
C591 B.n17 VSUBS 0.006697f
C592 B.n18 VSUBS 0.006697f
C593 B.n19 VSUBS 0.006697f
C594 B.n20 VSUBS 0.015427f
C595 B.n21 VSUBS 0.006697f
C596 B.n22 VSUBS 0.006697f
C597 B.n23 VSUBS 0.006697f
C598 B.n24 VSUBS 0.006697f
C599 B.n25 VSUBS 0.006697f
C600 B.n26 VSUBS 0.006697f
C601 B.n27 VSUBS 0.006697f
C602 B.n28 VSUBS 0.006697f
C603 B.n29 VSUBS 0.006697f
C604 B.n30 VSUBS 0.006697f
C605 B.n31 VSUBS 0.006697f
C606 B.n32 VSUBS 0.006697f
C607 B.n33 VSUBS 0.006697f
C608 B.n34 VSUBS 0.006697f
C609 B.n35 VSUBS 0.006697f
C610 B.n36 VSUBS 0.006697f
C611 B.n37 VSUBS 0.006697f
C612 B.n38 VSUBS 0.006697f
C613 B.n39 VSUBS 0.006697f
C614 B.t8 VSUBS 0.186515f
C615 B.t7 VSUBS 0.218733f
C616 B.t6 VSUBS 1.40416f
C617 B.n40 VSUBS 0.350392f
C618 B.n41 VSUBS 0.232342f
C619 B.n42 VSUBS 0.015517f
C620 B.n43 VSUBS 0.006697f
C621 B.n44 VSUBS 0.006697f
C622 B.n45 VSUBS 0.006697f
C623 B.n46 VSUBS 0.006697f
C624 B.n47 VSUBS 0.006697f
C625 B.t5 VSUBS 0.186518f
C626 B.t4 VSUBS 0.218735f
C627 B.t3 VSUBS 1.40416f
C628 B.n48 VSUBS 0.35039f
C629 B.n49 VSUBS 0.232339f
C630 B.n50 VSUBS 0.006697f
C631 B.n51 VSUBS 0.006697f
C632 B.n52 VSUBS 0.006697f
C633 B.n53 VSUBS 0.006697f
C634 B.n54 VSUBS 0.006697f
C635 B.n55 VSUBS 0.006697f
C636 B.n56 VSUBS 0.006697f
C637 B.n57 VSUBS 0.006697f
C638 B.n58 VSUBS 0.006697f
C639 B.n59 VSUBS 0.006697f
C640 B.n60 VSUBS 0.006697f
C641 B.n61 VSUBS 0.006697f
C642 B.n62 VSUBS 0.006697f
C643 B.n63 VSUBS 0.006697f
C644 B.n64 VSUBS 0.006697f
C645 B.n65 VSUBS 0.006697f
C646 B.n66 VSUBS 0.006697f
C647 B.n67 VSUBS 0.006697f
C648 B.n68 VSUBS 0.006697f
C649 B.n69 VSUBS 0.014318f
C650 B.n70 VSUBS 0.006697f
C651 B.n71 VSUBS 0.006697f
C652 B.n72 VSUBS 0.006697f
C653 B.n73 VSUBS 0.006697f
C654 B.n74 VSUBS 0.006697f
C655 B.n75 VSUBS 0.006697f
C656 B.n76 VSUBS 0.006697f
C657 B.n77 VSUBS 0.006697f
C658 B.n78 VSUBS 0.006697f
C659 B.n79 VSUBS 0.006697f
C660 B.n80 VSUBS 0.006697f
C661 B.n81 VSUBS 0.006697f
C662 B.n82 VSUBS 0.006697f
C663 B.n83 VSUBS 0.006697f
C664 B.n84 VSUBS 0.006697f
C665 B.n85 VSUBS 0.006697f
C666 B.n86 VSUBS 0.006697f
C667 B.n87 VSUBS 0.006697f
C668 B.n88 VSUBS 0.006697f
C669 B.n89 VSUBS 0.006697f
C670 B.n90 VSUBS 0.006697f
C671 B.n91 VSUBS 0.006697f
C672 B.n92 VSUBS 0.006697f
C673 B.n93 VSUBS 0.006697f
C674 B.n94 VSUBS 0.006697f
C675 B.n95 VSUBS 0.006697f
C676 B.n96 VSUBS 0.006697f
C677 B.n97 VSUBS 0.006697f
C678 B.n98 VSUBS 0.006697f
C679 B.n99 VSUBS 0.006697f
C680 B.n100 VSUBS 0.006697f
C681 B.n101 VSUBS 0.006697f
C682 B.n102 VSUBS 0.006697f
C683 B.n103 VSUBS 0.006697f
C684 B.n104 VSUBS 0.006697f
C685 B.n105 VSUBS 0.014318f
C686 B.n106 VSUBS 0.006697f
C687 B.n107 VSUBS 0.006697f
C688 B.n108 VSUBS 0.006697f
C689 B.n109 VSUBS 0.006697f
C690 B.n110 VSUBS 0.006697f
C691 B.n111 VSUBS 0.006697f
C692 B.n112 VSUBS 0.006697f
C693 B.n113 VSUBS 0.006697f
C694 B.n114 VSUBS 0.006697f
C695 B.n115 VSUBS 0.006697f
C696 B.n116 VSUBS 0.006697f
C697 B.n117 VSUBS 0.006697f
C698 B.n118 VSUBS 0.006697f
C699 B.n119 VSUBS 0.006697f
C700 B.n120 VSUBS 0.006697f
C701 B.n121 VSUBS 0.006697f
C702 B.n122 VSUBS 0.006697f
C703 B.n123 VSUBS 0.006697f
C704 B.n124 VSUBS 0.006697f
C705 B.n125 VSUBS 0.006697f
C706 B.t10 VSUBS 0.186518f
C707 B.t11 VSUBS 0.218735f
C708 B.t9 VSUBS 1.40416f
C709 B.n126 VSUBS 0.35039f
C710 B.n127 VSUBS 0.232339f
C711 B.n128 VSUBS 0.006697f
C712 B.n129 VSUBS 0.006697f
C713 B.n130 VSUBS 0.006697f
C714 B.n131 VSUBS 0.006697f
C715 B.t1 VSUBS 0.186515f
C716 B.t2 VSUBS 0.218733f
C717 B.t0 VSUBS 1.40416f
C718 B.n132 VSUBS 0.350392f
C719 B.n133 VSUBS 0.232342f
C720 B.n134 VSUBS 0.015517f
C721 B.n135 VSUBS 0.006697f
C722 B.n136 VSUBS 0.006697f
C723 B.n137 VSUBS 0.006697f
C724 B.n138 VSUBS 0.006697f
C725 B.n139 VSUBS 0.006697f
C726 B.n140 VSUBS 0.006697f
C727 B.n141 VSUBS 0.006697f
C728 B.n142 VSUBS 0.006697f
C729 B.n143 VSUBS 0.006697f
C730 B.n144 VSUBS 0.006697f
C731 B.n145 VSUBS 0.006697f
C732 B.n146 VSUBS 0.006697f
C733 B.n147 VSUBS 0.006697f
C734 B.n148 VSUBS 0.006697f
C735 B.n149 VSUBS 0.006697f
C736 B.n150 VSUBS 0.006697f
C737 B.n151 VSUBS 0.006697f
C738 B.n152 VSUBS 0.006697f
C739 B.n153 VSUBS 0.006697f
C740 B.n154 VSUBS 0.015427f
C741 B.n155 VSUBS 0.006697f
C742 B.n156 VSUBS 0.006697f
C743 B.n157 VSUBS 0.006697f
C744 B.n158 VSUBS 0.006697f
C745 B.n159 VSUBS 0.006697f
C746 B.n160 VSUBS 0.006697f
C747 B.n161 VSUBS 0.006697f
C748 B.n162 VSUBS 0.006697f
C749 B.n163 VSUBS 0.006697f
C750 B.n164 VSUBS 0.006697f
C751 B.n165 VSUBS 0.006697f
C752 B.n166 VSUBS 0.006697f
C753 B.n167 VSUBS 0.006697f
C754 B.n168 VSUBS 0.006697f
C755 B.n169 VSUBS 0.006697f
C756 B.n170 VSUBS 0.006697f
C757 B.n171 VSUBS 0.006697f
C758 B.n172 VSUBS 0.006697f
C759 B.n173 VSUBS 0.006697f
C760 B.n174 VSUBS 0.006697f
C761 B.n175 VSUBS 0.006697f
C762 B.n176 VSUBS 0.006697f
C763 B.n177 VSUBS 0.006697f
C764 B.n178 VSUBS 0.006697f
C765 B.n179 VSUBS 0.006697f
C766 B.n180 VSUBS 0.006697f
C767 B.n181 VSUBS 0.006697f
C768 B.n182 VSUBS 0.006697f
C769 B.n183 VSUBS 0.006697f
C770 B.n184 VSUBS 0.006697f
C771 B.n185 VSUBS 0.006697f
C772 B.n186 VSUBS 0.006697f
C773 B.n187 VSUBS 0.006697f
C774 B.n188 VSUBS 0.006697f
C775 B.n189 VSUBS 0.006697f
C776 B.n190 VSUBS 0.006697f
C777 B.n191 VSUBS 0.006697f
C778 B.n192 VSUBS 0.006697f
C779 B.n193 VSUBS 0.006697f
C780 B.n194 VSUBS 0.006697f
C781 B.n195 VSUBS 0.006697f
C782 B.n196 VSUBS 0.006697f
C783 B.n197 VSUBS 0.006697f
C784 B.n198 VSUBS 0.006697f
C785 B.n199 VSUBS 0.006697f
C786 B.n200 VSUBS 0.006697f
C787 B.n201 VSUBS 0.006697f
C788 B.n202 VSUBS 0.006697f
C789 B.n203 VSUBS 0.006697f
C790 B.n204 VSUBS 0.006697f
C791 B.n205 VSUBS 0.006697f
C792 B.n206 VSUBS 0.006697f
C793 B.n207 VSUBS 0.006697f
C794 B.n208 VSUBS 0.006697f
C795 B.n209 VSUBS 0.006697f
C796 B.n210 VSUBS 0.006697f
C797 B.n211 VSUBS 0.006697f
C798 B.n212 VSUBS 0.006697f
C799 B.n213 VSUBS 0.006697f
C800 B.n214 VSUBS 0.006697f
C801 B.n215 VSUBS 0.006697f
C802 B.n216 VSUBS 0.006697f
C803 B.n217 VSUBS 0.006697f
C804 B.n218 VSUBS 0.006697f
C805 B.n219 VSUBS 0.006697f
C806 B.n220 VSUBS 0.006697f
C807 B.n221 VSUBS 0.006697f
C808 B.n222 VSUBS 0.006697f
C809 B.n223 VSUBS 0.014318f
C810 B.n224 VSUBS 0.014318f
C811 B.n225 VSUBS 0.015427f
C812 B.n226 VSUBS 0.006697f
C813 B.n227 VSUBS 0.006697f
C814 B.n228 VSUBS 0.006697f
C815 B.n229 VSUBS 0.006697f
C816 B.n230 VSUBS 0.006697f
C817 B.n231 VSUBS 0.006697f
C818 B.n232 VSUBS 0.006697f
C819 B.n233 VSUBS 0.006697f
C820 B.n234 VSUBS 0.006697f
C821 B.n235 VSUBS 0.006697f
C822 B.n236 VSUBS 0.006697f
C823 B.n237 VSUBS 0.006697f
C824 B.n238 VSUBS 0.006697f
C825 B.n239 VSUBS 0.006697f
C826 B.n240 VSUBS 0.006697f
C827 B.n241 VSUBS 0.006697f
C828 B.n242 VSUBS 0.006697f
C829 B.n243 VSUBS 0.006697f
C830 B.n244 VSUBS 0.006697f
C831 B.n245 VSUBS 0.006697f
C832 B.n246 VSUBS 0.006697f
C833 B.n247 VSUBS 0.006697f
C834 B.n248 VSUBS 0.006697f
C835 B.n249 VSUBS 0.006697f
C836 B.n250 VSUBS 0.006697f
C837 B.n251 VSUBS 0.006697f
C838 B.n252 VSUBS 0.006697f
C839 B.n253 VSUBS 0.006697f
C840 B.n254 VSUBS 0.006697f
C841 B.n255 VSUBS 0.006697f
C842 B.n256 VSUBS 0.006697f
C843 B.n257 VSUBS 0.006697f
C844 B.n258 VSUBS 0.006697f
C845 B.n259 VSUBS 0.006697f
C846 B.n260 VSUBS 0.006697f
C847 B.n261 VSUBS 0.006697f
C848 B.n262 VSUBS 0.006697f
C849 B.n263 VSUBS 0.006697f
C850 B.n264 VSUBS 0.006697f
C851 B.n265 VSUBS 0.006697f
C852 B.n266 VSUBS 0.006697f
C853 B.n267 VSUBS 0.006697f
C854 B.n268 VSUBS 0.006697f
C855 B.n269 VSUBS 0.006697f
C856 B.n270 VSUBS 0.006697f
C857 B.n271 VSUBS 0.006697f
C858 B.n272 VSUBS 0.006697f
C859 B.n273 VSUBS 0.006697f
C860 B.n274 VSUBS 0.006697f
C861 B.n275 VSUBS 0.006697f
C862 B.n276 VSUBS 0.006697f
C863 B.n277 VSUBS 0.006697f
C864 B.n278 VSUBS 0.006697f
C865 B.n279 VSUBS 0.006697f
C866 B.n280 VSUBS 0.006697f
C867 B.n281 VSUBS 0.006697f
C868 B.n282 VSUBS 0.006697f
C869 B.n283 VSUBS 0.004629f
C870 B.n284 VSUBS 0.006697f
C871 B.n285 VSUBS 0.006697f
C872 B.n286 VSUBS 0.005417f
C873 B.n287 VSUBS 0.006697f
C874 B.n288 VSUBS 0.006697f
C875 B.n289 VSUBS 0.006697f
C876 B.n290 VSUBS 0.006697f
C877 B.n291 VSUBS 0.006697f
C878 B.n292 VSUBS 0.006697f
C879 B.n293 VSUBS 0.006697f
C880 B.n294 VSUBS 0.006697f
C881 B.n295 VSUBS 0.006697f
C882 B.n296 VSUBS 0.006697f
C883 B.n297 VSUBS 0.006697f
C884 B.n298 VSUBS 0.005417f
C885 B.n299 VSUBS 0.015517f
C886 B.n300 VSUBS 0.004629f
C887 B.n301 VSUBS 0.006697f
C888 B.n302 VSUBS 0.006697f
C889 B.n303 VSUBS 0.006697f
C890 B.n304 VSUBS 0.006697f
C891 B.n305 VSUBS 0.006697f
C892 B.n306 VSUBS 0.006697f
C893 B.n307 VSUBS 0.006697f
C894 B.n308 VSUBS 0.006697f
C895 B.n309 VSUBS 0.006697f
C896 B.n310 VSUBS 0.006697f
C897 B.n311 VSUBS 0.006697f
C898 B.n312 VSUBS 0.006697f
C899 B.n313 VSUBS 0.006697f
C900 B.n314 VSUBS 0.006697f
C901 B.n315 VSUBS 0.006697f
C902 B.n316 VSUBS 0.006697f
C903 B.n317 VSUBS 0.006697f
C904 B.n318 VSUBS 0.006697f
C905 B.n319 VSUBS 0.006697f
C906 B.n320 VSUBS 0.006697f
C907 B.n321 VSUBS 0.006697f
C908 B.n322 VSUBS 0.006697f
C909 B.n323 VSUBS 0.006697f
C910 B.n324 VSUBS 0.006697f
C911 B.n325 VSUBS 0.006697f
C912 B.n326 VSUBS 0.006697f
C913 B.n327 VSUBS 0.006697f
C914 B.n328 VSUBS 0.006697f
C915 B.n329 VSUBS 0.006697f
C916 B.n330 VSUBS 0.006697f
C917 B.n331 VSUBS 0.006697f
C918 B.n332 VSUBS 0.006697f
C919 B.n333 VSUBS 0.006697f
C920 B.n334 VSUBS 0.006697f
C921 B.n335 VSUBS 0.006697f
C922 B.n336 VSUBS 0.006697f
C923 B.n337 VSUBS 0.006697f
C924 B.n338 VSUBS 0.006697f
C925 B.n339 VSUBS 0.006697f
C926 B.n340 VSUBS 0.006697f
C927 B.n341 VSUBS 0.006697f
C928 B.n342 VSUBS 0.006697f
C929 B.n343 VSUBS 0.006697f
C930 B.n344 VSUBS 0.006697f
C931 B.n345 VSUBS 0.006697f
C932 B.n346 VSUBS 0.006697f
C933 B.n347 VSUBS 0.006697f
C934 B.n348 VSUBS 0.006697f
C935 B.n349 VSUBS 0.006697f
C936 B.n350 VSUBS 0.006697f
C937 B.n351 VSUBS 0.006697f
C938 B.n352 VSUBS 0.006697f
C939 B.n353 VSUBS 0.006697f
C940 B.n354 VSUBS 0.006697f
C941 B.n355 VSUBS 0.006697f
C942 B.n356 VSUBS 0.006697f
C943 B.n357 VSUBS 0.006697f
C944 B.n358 VSUBS 0.015427f
C945 B.n359 VSUBS 0.015427f
C946 B.n360 VSUBS 0.014318f
C947 B.n361 VSUBS 0.006697f
C948 B.n362 VSUBS 0.006697f
C949 B.n363 VSUBS 0.006697f
C950 B.n364 VSUBS 0.006697f
C951 B.n365 VSUBS 0.006697f
C952 B.n366 VSUBS 0.006697f
C953 B.n367 VSUBS 0.006697f
C954 B.n368 VSUBS 0.006697f
C955 B.n369 VSUBS 0.006697f
C956 B.n370 VSUBS 0.006697f
C957 B.n371 VSUBS 0.006697f
C958 B.n372 VSUBS 0.006697f
C959 B.n373 VSUBS 0.006697f
C960 B.n374 VSUBS 0.006697f
C961 B.n375 VSUBS 0.006697f
C962 B.n376 VSUBS 0.006697f
C963 B.n377 VSUBS 0.006697f
C964 B.n378 VSUBS 0.006697f
C965 B.n379 VSUBS 0.006697f
C966 B.n380 VSUBS 0.006697f
C967 B.n381 VSUBS 0.006697f
C968 B.n382 VSUBS 0.006697f
C969 B.n383 VSUBS 0.006697f
C970 B.n384 VSUBS 0.006697f
C971 B.n385 VSUBS 0.006697f
C972 B.n386 VSUBS 0.006697f
C973 B.n387 VSUBS 0.006697f
C974 B.n388 VSUBS 0.006697f
C975 B.n389 VSUBS 0.006697f
C976 B.n390 VSUBS 0.006697f
C977 B.n391 VSUBS 0.006697f
C978 B.n392 VSUBS 0.006697f
C979 B.n393 VSUBS 0.006697f
C980 B.n394 VSUBS 0.006697f
C981 B.n395 VSUBS 0.006697f
C982 B.n396 VSUBS 0.006697f
C983 B.n397 VSUBS 0.006697f
C984 B.n398 VSUBS 0.006697f
C985 B.n399 VSUBS 0.006697f
C986 B.n400 VSUBS 0.006697f
C987 B.n401 VSUBS 0.006697f
C988 B.n402 VSUBS 0.006697f
C989 B.n403 VSUBS 0.006697f
C990 B.n404 VSUBS 0.006697f
C991 B.n405 VSUBS 0.006697f
C992 B.n406 VSUBS 0.006697f
C993 B.n407 VSUBS 0.006697f
C994 B.n408 VSUBS 0.006697f
C995 B.n409 VSUBS 0.006697f
C996 B.n410 VSUBS 0.006697f
C997 B.n411 VSUBS 0.006697f
C998 B.n412 VSUBS 0.006697f
C999 B.n413 VSUBS 0.006697f
C1000 B.n414 VSUBS 0.006697f
C1001 B.n415 VSUBS 0.006697f
C1002 B.n416 VSUBS 0.006697f
C1003 B.n417 VSUBS 0.006697f
C1004 B.n418 VSUBS 0.006697f
C1005 B.n419 VSUBS 0.006697f
C1006 B.n420 VSUBS 0.006697f
C1007 B.n421 VSUBS 0.006697f
C1008 B.n422 VSUBS 0.006697f
C1009 B.n423 VSUBS 0.006697f
C1010 B.n424 VSUBS 0.006697f
C1011 B.n425 VSUBS 0.006697f
C1012 B.n426 VSUBS 0.006697f
C1013 B.n427 VSUBS 0.006697f
C1014 B.n428 VSUBS 0.006697f
C1015 B.n429 VSUBS 0.006697f
C1016 B.n430 VSUBS 0.006697f
C1017 B.n431 VSUBS 0.006697f
C1018 B.n432 VSUBS 0.006697f
C1019 B.n433 VSUBS 0.006697f
C1020 B.n434 VSUBS 0.006697f
C1021 B.n435 VSUBS 0.006697f
C1022 B.n436 VSUBS 0.006697f
C1023 B.n437 VSUBS 0.006697f
C1024 B.n438 VSUBS 0.006697f
C1025 B.n439 VSUBS 0.006697f
C1026 B.n440 VSUBS 0.006697f
C1027 B.n441 VSUBS 0.006697f
C1028 B.n442 VSUBS 0.006697f
C1029 B.n443 VSUBS 0.006697f
C1030 B.n444 VSUBS 0.006697f
C1031 B.n445 VSUBS 0.006697f
C1032 B.n446 VSUBS 0.006697f
C1033 B.n447 VSUBS 0.006697f
C1034 B.n448 VSUBS 0.006697f
C1035 B.n449 VSUBS 0.006697f
C1036 B.n450 VSUBS 0.006697f
C1037 B.n451 VSUBS 0.006697f
C1038 B.n452 VSUBS 0.006697f
C1039 B.n453 VSUBS 0.006697f
C1040 B.n454 VSUBS 0.006697f
C1041 B.n455 VSUBS 0.006697f
C1042 B.n456 VSUBS 0.006697f
C1043 B.n457 VSUBS 0.006697f
C1044 B.n458 VSUBS 0.006697f
C1045 B.n459 VSUBS 0.006697f
C1046 B.n460 VSUBS 0.006697f
C1047 B.n461 VSUBS 0.006697f
C1048 B.n462 VSUBS 0.006697f
C1049 B.n463 VSUBS 0.006697f
C1050 B.n464 VSUBS 0.006697f
C1051 B.n465 VSUBS 0.006697f
C1052 B.n466 VSUBS 0.006697f
C1053 B.n467 VSUBS 0.006697f
C1054 B.n468 VSUBS 0.015176f
C1055 B.n469 VSUBS 0.014569f
C1056 B.n470 VSUBS 0.015427f
C1057 B.n471 VSUBS 0.006697f
C1058 B.n472 VSUBS 0.006697f
C1059 B.n473 VSUBS 0.006697f
C1060 B.n474 VSUBS 0.006697f
C1061 B.n475 VSUBS 0.006697f
C1062 B.n476 VSUBS 0.006697f
C1063 B.n477 VSUBS 0.006697f
C1064 B.n478 VSUBS 0.006697f
C1065 B.n479 VSUBS 0.006697f
C1066 B.n480 VSUBS 0.006697f
C1067 B.n481 VSUBS 0.006697f
C1068 B.n482 VSUBS 0.006697f
C1069 B.n483 VSUBS 0.006697f
C1070 B.n484 VSUBS 0.006697f
C1071 B.n485 VSUBS 0.006697f
C1072 B.n486 VSUBS 0.006697f
C1073 B.n487 VSUBS 0.006697f
C1074 B.n488 VSUBS 0.006697f
C1075 B.n489 VSUBS 0.006697f
C1076 B.n490 VSUBS 0.006697f
C1077 B.n491 VSUBS 0.006697f
C1078 B.n492 VSUBS 0.006697f
C1079 B.n493 VSUBS 0.006697f
C1080 B.n494 VSUBS 0.006697f
C1081 B.n495 VSUBS 0.006697f
C1082 B.n496 VSUBS 0.006697f
C1083 B.n497 VSUBS 0.006697f
C1084 B.n498 VSUBS 0.006697f
C1085 B.n499 VSUBS 0.006697f
C1086 B.n500 VSUBS 0.006697f
C1087 B.n501 VSUBS 0.006697f
C1088 B.n502 VSUBS 0.006697f
C1089 B.n503 VSUBS 0.006697f
C1090 B.n504 VSUBS 0.006697f
C1091 B.n505 VSUBS 0.006697f
C1092 B.n506 VSUBS 0.006697f
C1093 B.n507 VSUBS 0.006697f
C1094 B.n508 VSUBS 0.006697f
C1095 B.n509 VSUBS 0.006697f
C1096 B.n510 VSUBS 0.006697f
C1097 B.n511 VSUBS 0.006697f
C1098 B.n512 VSUBS 0.006697f
C1099 B.n513 VSUBS 0.006697f
C1100 B.n514 VSUBS 0.006697f
C1101 B.n515 VSUBS 0.006697f
C1102 B.n516 VSUBS 0.006697f
C1103 B.n517 VSUBS 0.006697f
C1104 B.n518 VSUBS 0.006697f
C1105 B.n519 VSUBS 0.006697f
C1106 B.n520 VSUBS 0.006697f
C1107 B.n521 VSUBS 0.006697f
C1108 B.n522 VSUBS 0.006697f
C1109 B.n523 VSUBS 0.006697f
C1110 B.n524 VSUBS 0.006697f
C1111 B.n525 VSUBS 0.006697f
C1112 B.n526 VSUBS 0.006697f
C1113 B.n527 VSUBS 0.006697f
C1114 B.n528 VSUBS 0.004629f
C1115 B.n529 VSUBS 0.015517f
C1116 B.n530 VSUBS 0.005417f
C1117 B.n531 VSUBS 0.006697f
C1118 B.n532 VSUBS 0.006697f
C1119 B.n533 VSUBS 0.006697f
C1120 B.n534 VSUBS 0.006697f
C1121 B.n535 VSUBS 0.006697f
C1122 B.n536 VSUBS 0.006697f
C1123 B.n537 VSUBS 0.006697f
C1124 B.n538 VSUBS 0.006697f
C1125 B.n539 VSUBS 0.006697f
C1126 B.n540 VSUBS 0.006697f
C1127 B.n541 VSUBS 0.006697f
C1128 B.n542 VSUBS 0.005417f
C1129 B.n543 VSUBS 0.006697f
C1130 B.n544 VSUBS 0.006697f
C1131 B.n545 VSUBS 0.004629f
C1132 B.n546 VSUBS 0.006697f
C1133 B.n547 VSUBS 0.006697f
C1134 B.n548 VSUBS 0.006697f
C1135 B.n549 VSUBS 0.006697f
C1136 B.n550 VSUBS 0.006697f
C1137 B.n551 VSUBS 0.006697f
C1138 B.n552 VSUBS 0.006697f
C1139 B.n553 VSUBS 0.006697f
C1140 B.n554 VSUBS 0.006697f
C1141 B.n555 VSUBS 0.006697f
C1142 B.n556 VSUBS 0.006697f
C1143 B.n557 VSUBS 0.006697f
C1144 B.n558 VSUBS 0.006697f
C1145 B.n559 VSUBS 0.006697f
C1146 B.n560 VSUBS 0.006697f
C1147 B.n561 VSUBS 0.006697f
C1148 B.n562 VSUBS 0.006697f
C1149 B.n563 VSUBS 0.006697f
C1150 B.n564 VSUBS 0.006697f
C1151 B.n565 VSUBS 0.006697f
C1152 B.n566 VSUBS 0.006697f
C1153 B.n567 VSUBS 0.006697f
C1154 B.n568 VSUBS 0.006697f
C1155 B.n569 VSUBS 0.006697f
C1156 B.n570 VSUBS 0.006697f
C1157 B.n571 VSUBS 0.006697f
C1158 B.n572 VSUBS 0.006697f
C1159 B.n573 VSUBS 0.006697f
C1160 B.n574 VSUBS 0.006697f
C1161 B.n575 VSUBS 0.006697f
C1162 B.n576 VSUBS 0.006697f
C1163 B.n577 VSUBS 0.006697f
C1164 B.n578 VSUBS 0.006697f
C1165 B.n579 VSUBS 0.006697f
C1166 B.n580 VSUBS 0.006697f
C1167 B.n581 VSUBS 0.006697f
C1168 B.n582 VSUBS 0.006697f
C1169 B.n583 VSUBS 0.006697f
C1170 B.n584 VSUBS 0.006697f
C1171 B.n585 VSUBS 0.006697f
C1172 B.n586 VSUBS 0.006697f
C1173 B.n587 VSUBS 0.006697f
C1174 B.n588 VSUBS 0.006697f
C1175 B.n589 VSUBS 0.006697f
C1176 B.n590 VSUBS 0.006697f
C1177 B.n591 VSUBS 0.006697f
C1178 B.n592 VSUBS 0.006697f
C1179 B.n593 VSUBS 0.006697f
C1180 B.n594 VSUBS 0.006697f
C1181 B.n595 VSUBS 0.006697f
C1182 B.n596 VSUBS 0.006697f
C1183 B.n597 VSUBS 0.006697f
C1184 B.n598 VSUBS 0.006697f
C1185 B.n599 VSUBS 0.006697f
C1186 B.n600 VSUBS 0.006697f
C1187 B.n601 VSUBS 0.006697f
C1188 B.n602 VSUBS 0.006697f
C1189 B.n603 VSUBS 0.015427f
C1190 B.n604 VSUBS 0.014318f
C1191 B.n605 VSUBS 0.014318f
C1192 B.n606 VSUBS 0.006697f
C1193 B.n607 VSUBS 0.006697f
C1194 B.n608 VSUBS 0.006697f
C1195 B.n609 VSUBS 0.006697f
C1196 B.n610 VSUBS 0.006697f
C1197 B.n611 VSUBS 0.006697f
C1198 B.n612 VSUBS 0.006697f
C1199 B.n613 VSUBS 0.006697f
C1200 B.n614 VSUBS 0.006697f
C1201 B.n615 VSUBS 0.006697f
C1202 B.n616 VSUBS 0.006697f
C1203 B.n617 VSUBS 0.006697f
C1204 B.n618 VSUBS 0.006697f
C1205 B.n619 VSUBS 0.006697f
C1206 B.n620 VSUBS 0.006697f
C1207 B.n621 VSUBS 0.006697f
C1208 B.n622 VSUBS 0.006697f
C1209 B.n623 VSUBS 0.006697f
C1210 B.n624 VSUBS 0.006697f
C1211 B.n625 VSUBS 0.006697f
C1212 B.n626 VSUBS 0.006697f
C1213 B.n627 VSUBS 0.006697f
C1214 B.n628 VSUBS 0.006697f
C1215 B.n629 VSUBS 0.006697f
C1216 B.n630 VSUBS 0.006697f
C1217 B.n631 VSUBS 0.006697f
C1218 B.n632 VSUBS 0.006697f
C1219 B.n633 VSUBS 0.006697f
C1220 B.n634 VSUBS 0.006697f
C1221 B.n635 VSUBS 0.006697f
C1222 B.n636 VSUBS 0.006697f
C1223 B.n637 VSUBS 0.006697f
C1224 B.n638 VSUBS 0.006697f
C1225 B.n639 VSUBS 0.006697f
C1226 B.n640 VSUBS 0.006697f
C1227 B.n641 VSUBS 0.006697f
C1228 B.n642 VSUBS 0.006697f
C1229 B.n643 VSUBS 0.006697f
C1230 B.n644 VSUBS 0.006697f
C1231 B.n645 VSUBS 0.006697f
C1232 B.n646 VSUBS 0.006697f
C1233 B.n647 VSUBS 0.006697f
C1234 B.n648 VSUBS 0.006697f
C1235 B.n649 VSUBS 0.006697f
C1236 B.n650 VSUBS 0.006697f
C1237 B.n651 VSUBS 0.006697f
C1238 B.n652 VSUBS 0.006697f
C1239 B.n653 VSUBS 0.006697f
C1240 B.n654 VSUBS 0.006697f
C1241 B.n655 VSUBS 0.006697f
C1242 B.n656 VSUBS 0.006697f
C1243 B.n657 VSUBS 0.006697f
C1244 B.n658 VSUBS 0.006697f
C1245 B.n659 VSUBS 0.015165f
.ends

