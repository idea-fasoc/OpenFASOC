* NGSPICE file created from diff_pair_sample_0641.ext - technology: sky130A

.subckt diff_pair_sample_0641 VTAIL VN VP B VDD2 VDD1
X0 B.t23 B.t21 B.t22 B.t15 sky130_fd_pr__nfet_01v8 ad=5.1753 pd=27.32 as=0 ps=0 w=13.27 l=1.58
X1 VTAIL.t19 VP.t0 VDD1.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=2.18955 pd=13.6 as=2.18955 ps=13.6 w=13.27 l=1.58
X2 VDD2.t9 VN.t0 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=5.1753 pd=27.32 as=2.18955 ps=13.6 w=13.27 l=1.58
X3 VDD2.t8 VN.t1 VTAIL.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=5.1753 pd=27.32 as=2.18955 ps=13.6 w=13.27 l=1.58
X4 VDD1.t4 VP.t1 VTAIL.t18 B.t3 sky130_fd_pr__nfet_01v8 ad=2.18955 pd=13.6 as=5.1753 ps=27.32 w=13.27 l=1.58
X5 VDD1.t1 VP.t2 VTAIL.t17 B.t5 sky130_fd_pr__nfet_01v8 ad=2.18955 pd=13.6 as=2.18955 ps=13.6 w=13.27 l=1.58
X6 VTAIL.t16 VP.t3 VDD1.t5 B.t4 sky130_fd_pr__nfet_01v8 ad=2.18955 pd=13.6 as=2.18955 ps=13.6 w=13.27 l=1.58
X7 VTAIL.t9 VN.t2 VDD2.t7 B.t8 sky130_fd_pr__nfet_01v8 ad=2.18955 pd=13.6 as=2.18955 ps=13.6 w=13.27 l=1.58
X8 VTAIL.t15 VP.t4 VDD1.t6 B.t9 sky130_fd_pr__nfet_01v8 ad=2.18955 pd=13.6 as=2.18955 ps=13.6 w=13.27 l=1.58
X9 VDD1.t8 VP.t5 VTAIL.t14 B.t7 sky130_fd_pr__nfet_01v8 ad=5.1753 pd=27.32 as=2.18955 ps=13.6 w=13.27 l=1.58
X10 VTAIL.t7 VN.t3 VDD2.t6 B.t9 sky130_fd_pr__nfet_01v8 ad=2.18955 pd=13.6 as=2.18955 ps=13.6 w=13.27 l=1.58
X11 VTAIL.t6 VN.t4 VDD2.t5 B.t4 sky130_fd_pr__nfet_01v8 ad=2.18955 pd=13.6 as=2.18955 ps=13.6 w=13.27 l=1.58
X12 VDD1.t0 VP.t6 VTAIL.t13 B.t0 sky130_fd_pr__nfet_01v8 ad=5.1753 pd=27.32 as=2.18955 ps=13.6 w=13.27 l=1.58
X13 VDD2.t4 VN.t5 VTAIL.t2 B.t3 sky130_fd_pr__nfet_01v8 ad=2.18955 pd=13.6 as=5.1753 ps=27.32 w=13.27 l=1.58
X14 VDD2.t3 VN.t6 VTAIL.t4 B.t6 sky130_fd_pr__nfet_01v8 ad=2.18955 pd=13.6 as=5.1753 ps=27.32 w=13.27 l=1.58
X15 VDD1.t7 VP.t7 VTAIL.t12 B.t1 sky130_fd_pr__nfet_01v8 ad=2.18955 pd=13.6 as=2.18955 ps=13.6 w=13.27 l=1.58
X16 VTAIL.t3 VN.t7 VDD2.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=2.18955 pd=13.6 as=2.18955 ps=13.6 w=13.27 l=1.58
X17 B.t20 B.t18 B.t19 B.t11 sky130_fd_pr__nfet_01v8 ad=5.1753 pd=27.32 as=0 ps=0 w=13.27 l=1.58
X18 VTAIL.t11 VP.t8 VDD1.t3 B.t8 sky130_fd_pr__nfet_01v8 ad=2.18955 pd=13.6 as=2.18955 ps=13.6 w=13.27 l=1.58
X19 VDD1.t9 VP.t9 VTAIL.t10 B.t6 sky130_fd_pr__nfet_01v8 ad=2.18955 pd=13.6 as=5.1753 ps=27.32 w=13.27 l=1.58
X20 B.t17 B.t14 B.t16 B.t15 sky130_fd_pr__nfet_01v8 ad=5.1753 pd=27.32 as=0 ps=0 w=13.27 l=1.58
X21 VDD2.t1 VN.t8 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=2.18955 pd=13.6 as=2.18955 ps=13.6 w=13.27 l=1.58
X22 VDD2.t0 VN.t9 VTAIL.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=2.18955 pd=13.6 as=2.18955 ps=13.6 w=13.27 l=1.58
X23 B.t13 B.t10 B.t12 B.t11 sky130_fd_pr__nfet_01v8 ad=5.1753 pd=27.32 as=0 ps=0 w=13.27 l=1.58
R0 B.n651 B.n650 585
R1 B.n653 B.n133 585
R2 B.n656 B.n655 585
R3 B.n657 B.n132 585
R4 B.n659 B.n658 585
R5 B.n661 B.n131 585
R6 B.n664 B.n663 585
R7 B.n665 B.n130 585
R8 B.n667 B.n666 585
R9 B.n669 B.n129 585
R10 B.n672 B.n671 585
R11 B.n673 B.n128 585
R12 B.n675 B.n674 585
R13 B.n677 B.n127 585
R14 B.n680 B.n679 585
R15 B.n681 B.n126 585
R16 B.n683 B.n682 585
R17 B.n685 B.n125 585
R18 B.n688 B.n687 585
R19 B.n689 B.n124 585
R20 B.n691 B.n690 585
R21 B.n693 B.n123 585
R22 B.n696 B.n695 585
R23 B.n697 B.n122 585
R24 B.n699 B.n698 585
R25 B.n701 B.n121 585
R26 B.n704 B.n703 585
R27 B.n705 B.n120 585
R28 B.n707 B.n706 585
R29 B.n709 B.n119 585
R30 B.n712 B.n711 585
R31 B.n713 B.n118 585
R32 B.n715 B.n714 585
R33 B.n717 B.n117 585
R34 B.n720 B.n719 585
R35 B.n721 B.n116 585
R36 B.n723 B.n722 585
R37 B.n725 B.n115 585
R38 B.n728 B.n727 585
R39 B.n729 B.n114 585
R40 B.n731 B.n730 585
R41 B.n733 B.n113 585
R42 B.n736 B.n735 585
R43 B.n737 B.n109 585
R44 B.n739 B.n738 585
R45 B.n741 B.n108 585
R46 B.n744 B.n743 585
R47 B.n745 B.n107 585
R48 B.n747 B.n746 585
R49 B.n749 B.n106 585
R50 B.n752 B.n751 585
R51 B.n753 B.n105 585
R52 B.n755 B.n754 585
R53 B.n757 B.n104 585
R54 B.n760 B.n759 585
R55 B.n762 B.n101 585
R56 B.n764 B.n763 585
R57 B.n766 B.n100 585
R58 B.n769 B.n768 585
R59 B.n770 B.n99 585
R60 B.n772 B.n771 585
R61 B.n774 B.n98 585
R62 B.n777 B.n776 585
R63 B.n778 B.n97 585
R64 B.n780 B.n779 585
R65 B.n782 B.n96 585
R66 B.n785 B.n784 585
R67 B.n786 B.n95 585
R68 B.n788 B.n787 585
R69 B.n790 B.n94 585
R70 B.n793 B.n792 585
R71 B.n794 B.n93 585
R72 B.n796 B.n795 585
R73 B.n798 B.n92 585
R74 B.n801 B.n800 585
R75 B.n802 B.n91 585
R76 B.n804 B.n803 585
R77 B.n806 B.n90 585
R78 B.n809 B.n808 585
R79 B.n810 B.n89 585
R80 B.n812 B.n811 585
R81 B.n814 B.n88 585
R82 B.n817 B.n816 585
R83 B.n818 B.n87 585
R84 B.n820 B.n819 585
R85 B.n822 B.n86 585
R86 B.n825 B.n824 585
R87 B.n826 B.n85 585
R88 B.n828 B.n827 585
R89 B.n830 B.n84 585
R90 B.n833 B.n832 585
R91 B.n834 B.n83 585
R92 B.n836 B.n835 585
R93 B.n838 B.n82 585
R94 B.n841 B.n840 585
R95 B.n842 B.n81 585
R96 B.n844 B.n843 585
R97 B.n846 B.n80 585
R98 B.n849 B.n848 585
R99 B.n850 B.n79 585
R100 B.n649 B.n77 585
R101 B.n853 B.n77 585
R102 B.n648 B.n76 585
R103 B.n854 B.n76 585
R104 B.n647 B.n75 585
R105 B.n855 B.n75 585
R106 B.n646 B.n645 585
R107 B.n645 B.n71 585
R108 B.n644 B.n70 585
R109 B.n861 B.n70 585
R110 B.n643 B.n69 585
R111 B.n862 B.n69 585
R112 B.n642 B.n68 585
R113 B.n863 B.n68 585
R114 B.n641 B.n640 585
R115 B.n640 B.n64 585
R116 B.n639 B.n63 585
R117 B.n869 B.n63 585
R118 B.n638 B.n62 585
R119 B.n870 B.n62 585
R120 B.n637 B.n61 585
R121 B.n871 B.n61 585
R122 B.n636 B.n635 585
R123 B.n635 B.n57 585
R124 B.n634 B.n56 585
R125 B.n877 B.n56 585
R126 B.n633 B.n55 585
R127 B.n878 B.n55 585
R128 B.n632 B.n54 585
R129 B.n879 B.n54 585
R130 B.n631 B.n630 585
R131 B.n630 B.n53 585
R132 B.n629 B.n49 585
R133 B.n885 B.n49 585
R134 B.n628 B.n48 585
R135 B.n886 B.n48 585
R136 B.n627 B.n47 585
R137 B.n887 B.n47 585
R138 B.n626 B.n625 585
R139 B.n625 B.n43 585
R140 B.n624 B.n42 585
R141 B.n893 B.n42 585
R142 B.n623 B.n41 585
R143 B.n894 B.n41 585
R144 B.n622 B.n40 585
R145 B.n895 B.n40 585
R146 B.n621 B.n620 585
R147 B.n620 B.n36 585
R148 B.n619 B.n35 585
R149 B.n901 B.n35 585
R150 B.n618 B.n34 585
R151 B.n902 B.n34 585
R152 B.n617 B.n33 585
R153 B.n903 B.n33 585
R154 B.n616 B.n615 585
R155 B.n615 B.n29 585
R156 B.n614 B.n28 585
R157 B.n909 B.n28 585
R158 B.n613 B.n27 585
R159 B.n910 B.n27 585
R160 B.n612 B.n26 585
R161 B.n911 B.n26 585
R162 B.n611 B.n610 585
R163 B.n610 B.n25 585
R164 B.n609 B.n21 585
R165 B.n917 B.n21 585
R166 B.n608 B.n20 585
R167 B.n918 B.n20 585
R168 B.n607 B.n19 585
R169 B.n919 B.n19 585
R170 B.n606 B.n605 585
R171 B.n605 B.n15 585
R172 B.n604 B.n14 585
R173 B.n925 B.n14 585
R174 B.n603 B.n13 585
R175 B.n926 B.n13 585
R176 B.n602 B.n12 585
R177 B.n927 B.n12 585
R178 B.n601 B.n600 585
R179 B.n600 B.n8 585
R180 B.n599 B.n7 585
R181 B.n933 B.n7 585
R182 B.n598 B.n6 585
R183 B.n934 B.n6 585
R184 B.n597 B.n5 585
R185 B.n935 B.n5 585
R186 B.n596 B.n595 585
R187 B.n595 B.n4 585
R188 B.n594 B.n134 585
R189 B.n594 B.n593 585
R190 B.n584 B.n135 585
R191 B.n136 B.n135 585
R192 B.n586 B.n585 585
R193 B.n587 B.n586 585
R194 B.n583 B.n140 585
R195 B.n144 B.n140 585
R196 B.n582 B.n581 585
R197 B.n581 B.n580 585
R198 B.n142 B.n141 585
R199 B.n143 B.n142 585
R200 B.n573 B.n572 585
R201 B.n574 B.n573 585
R202 B.n571 B.n149 585
R203 B.n149 B.n148 585
R204 B.n570 B.n569 585
R205 B.n569 B.n568 585
R206 B.n151 B.n150 585
R207 B.n561 B.n151 585
R208 B.n560 B.n559 585
R209 B.n562 B.n560 585
R210 B.n558 B.n156 585
R211 B.n156 B.n155 585
R212 B.n557 B.n556 585
R213 B.n556 B.n555 585
R214 B.n158 B.n157 585
R215 B.n159 B.n158 585
R216 B.n548 B.n547 585
R217 B.n549 B.n548 585
R218 B.n546 B.n164 585
R219 B.n164 B.n163 585
R220 B.n545 B.n544 585
R221 B.n544 B.n543 585
R222 B.n166 B.n165 585
R223 B.n167 B.n166 585
R224 B.n536 B.n535 585
R225 B.n537 B.n536 585
R226 B.n534 B.n172 585
R227 B.n172 B.n171 585
R228 B.n533 B.n532 585
R229 B.n532 B.n531 585
R230 B.n174 B.n173 585
R231 B.n175 B.n174 585
R232 B.n524 B.n523 585
R233 B.n525 B.n524 585
R234 B.n522 B.n180 585
R235 B.n180 B.n179 585
R236 B.n521 B.n520 585
R237 B.n520 B.n519 585
R238 B.n182 B.n181 585
R239 B.n512 B.n182 585
R240 B.n511 B.n510 585
R241 B.n513 B.n511 585
R242 B.n509 B.n187 585
R243 B.n187 B.n186 585
R244 B.n508 B.n507 585
R245 B.n507 B.n506 585
R246 B.n189 B.n188 585
R247 B.n190 B.n189 585
R248 B.n499 B.n498 585
R249 B.n500 B.n499 585
R250 B.n497 B.n195 585
R251 B.n195 B.n194 585
R252 B.n496 B.n495 585
R253 B.n495 B.n494 585
R254 B.n197 B.n196 585
R255 B.n198 B.n197 585
R256 B.n487 B.n486 585
R257 B.n488 B.n487 585
R258 B.n485 B.n203 585
R259 B.n203 B.n202 585
R260 B.n484 B.n483 585
R261 B.n483 B.n482 585
R262 B.n205 B.n204 585
R263 B.n206 B.n205 585
R264 B.n475 B.n474 585
R265 B.n476 B.n475 585
R266 B.n473 B.n211 585
R267 B.n211 B.n210 585
R268 B.n472 B.n471 585
R269 B.n471 B.n470 585
R270 B.n467 B.n215 585
R271 B.n466 B.n465 585
R272 B.n463 B.n216 585
R273 B.n463 B.n214 585
R274 B.n462 B.n461 585
R275 B.n460 B.n459 585
R276 B.n458 B.n218 585
R277 B.n456 B.n455 585
R278 B.n454 B.n219 585
R279 B.n453 B.n452 585
R280 B.n450 B.n220 585
R281 B.n448 B.n447 585
R282 B.n446 B.n221 585
R283 B.n445 B.n444 585
R284 B.n442 B.n222 585
R285 B.n440 B.n439 585
R286 B.n438 B.n223 585
R287 B.n437 B.n436 585
R288 B.n434 B.n224 585
R289 B.n432 B.n431 585
R290 B.n430 B.n225 585
R291 B.n429 B.n428 585
R292 B.n426 B.n226 585
R293 B.n424 B.n423 585
R294 B.n422 B.n227 585
R295 B.n421 B.n420 585
R296 B.n418 B.n228 585
R297 B.n416 B.n415 585
R298 B.n414 B.n229 585
R299 B.n413 B.n412 585
R300 B.n410 B.n230 585
R301 B.n408 B.n407 585
R302 B.n406 B.n231 585
R303 B.n405 B.n404 585
R304 B.n402 B.n232 585
R305 B.n400 B.n399 585
R306 B.n398 B.n233 585
R307 B.n397 B.n396 585
R308 B.n394 B.n234 585
R309 B.n392 B.n391 585
R310 B.n390 B.n235 585
R311 B.n389 B.n388 585
R312 B.n386 B.n236 585
R313 B.n384 B.n383 585
R314 B.n382 B.n237 585
R315 B.n381 B.n380 585
R316 B.n378 B.n377 585
R317 B.n376 B.n375 585
R318 B.n374 B.n242 585
R319 B.n372 B.n371 585
R320 B.n370 B.n243 585
R321 B.n369 B.n368 585
R322 B.n366 B.n244 585
R323 B.n364 B.n363 585
R324 B.n362 B.n245 585
R325 B.n361 B.n360 585
R326 B.n358 B.n357 585
R327 B.n356 B.n355 585
R328 B.n354 B.n250 585
R329 B.n352 B.n351 585
R330 B.n350 B.n251 585
R331 B.n349 B.n348 585
R332 B.n346 B.n252 585
R333 B.n344 B.n343 585
R334 B.n342 B.n253 585
R335 B.n341 B.n340 585
R336 B.n338 B.n254 585
R337 B.n336 B.n335 585
R338 B.n334 B.n255 585
R339 B.n333 B.n332 585
R340 B.n330 B.n256 585
R341 B.n328 B.n327 585
R342 B.n326 B.n257 585
R343 B.n325 B.n324 585
R344 B.n322 B.n258 585
R345 B.n320 B.n319 585
R346 B.n318 B.n259 585
R347 B.n317 B.n316 585
R348 B.n314 B.n260 585
R349 B.n312 B.n311 585
R350 B.n310 B.n261 585
R351 B.n309 B.n308 585
R352 B.n306 B.n262 585
R353 B.n304 B.n303 585
R354 B.n302 B.n263 585
R355 B.n301 B.n300 585
R356 B.n298 B.n264 585
R357 B.n296 B.n295 585
R358 B.n294 B.n265 585
R359 B.n293 B.n292 585
R360 B.n290 B.n266 585
R361 B.n288 B.n287 585
R362 B.n286 B.n267 585
R363 B.n285 B.n284 585
R364 B.n282 B.n268 585
R365 B.n280 B.n279 585
R366 B.n278 B.n269 585
R367 B.n277 B.n276 585
R368 B.n274 B.n270 585
R369 B.n272 B.n271 585
R370 B.n213 B.n212 585
R371 B.n214 B.n213 585
R372 B.n469 B.n468 585
R373 B.n470 B.n469 585
R374 B.n209 B.n208 585
R375 B.n210 B.n209 585
R376 B.n478 B.n477 585
R377 B.n477 B.n476 585
R378 B.n479 B.n207 585
R379 B.n207 B.n206 585
R380 B.n481 B.n480 585
R381 B.n482 B.n481 585
R382 B.n201 B.n200 585
R383 B.n202 B.n201 585
R384 B.n490 B.n489 585
R385 B.n489 B.n488 585
R386 B.n491 B.n199 585
R387 B.n199 B.n198 585
R388 B.n493 B.n492 585
R389 B.n494 B.n493 585
R390 B.n193 B.n192 585
R391 B.n194 B.n193 585
R392 B.n502 B.n501 585
R393 B.n501 B.n500 585
R394 B.n503 B.n191 585
R395 B.n191 B.n190 585
R396 B.n505 B.n504 585
R397 B.n506 B.n505 585
R398 B.n185 B.n184 585
R399 B.n186 B.n185 585
R400 B.n515 B.n514 585
R401 B.n514 B.n513 585
R402 B.n516 B.n183 585
R403 B.n512 B.n183 585
R404 B.n518 B.n517 585
R405 B.n519 B.n518 585
R406 B.n178 B.n177 585
R407 B.n179 B.n178 585
R408 B.n527 B.n526 585
R409 B.n526 B.n525 585
R410 B.n528 B.n176 585
R411 B.n176 B.n175 585
R412 B.n530 B.n529 585
R413 B.n531 B.n530 585
R414 B.n170 B.n169 585
R415 B.n171 B.n170 585
R416 B.n539 B.n538 585
R417 B.n538 B.n537 585
R418 B.n540 B.n168 585
R419 B.n168 B.n167 585
R420 B.n542 B.n541 585
R421 B.n543 B.n542 585
R422 B.n162 B.n161 585
R423 B.n163 B.n162 585
R424 B.n551 B.n550 585
R425 B.n550 B.n549 585
R426 B.n552 B.n160 585
R427 B.n160 B.n159 585
R428 B.n554 B.n553 585
R429 B.n555 B.n554 585
R430 B.n154 B.n153 585
R431 B.n155 B.n154 585
R432 B.n564 B.n563 585
R433 B.n563 B.n562 585
R434 B.n565 B.n152 585
R435 B.n561 B.n152 585
R436 B.n567 B.n566 585
R437 B.n568 B.n567 585
R438 B.n147 B.n146 585
R439 B.n148 B.n147 585
R440 B.n576 B.n575 585
R441 B.n575 B.n574 585
R442 B.n577 B.n145 585
R443 B.n145 B.n143 585
R444 B.n579 B.n578 585
R445 B.n580 B.n579 585
R446 B.n139 B.n138 585
R447 B.n144 B.n139 585
R448 B.n589 B.n588 585
R449 B.n588 B.n587 585
R450 B.n590 B.n137 585
R451 B.n137 B.n136 585
R452 B.n592 B.n591 585
R453 B.n593 B.n592 585
R454 B.n2 B.n0 585
R455 B.n4 B.n2 585
R456 B.n3 B.n1 585
R457 B.n934 B.n3 585
R458 B.n932 B.n931 585
R459 B.n933 B.n932 585
R460 B.n930 B.n9 585
R461 B.n9 B.n8 585
R462 B.n929 B.n928 585
R463 B.n928 B.n927 585
R464 B.n11 B.n10 585
R465 B.n926 B.n11 585
R466 B.n924 B.n923 585
R467 B.n925 B.n924 585
R468 B.n922 B.n16 585
R469 B.n16 B.n15 585
R470 B.n921 B.n920 585
R471 B.n920 B.n919 585
R472 B.n18 B.n17 585
R473 B.n918 B.n18 585
R474 B.n916 B.n915 585
R475 B.n917 B.n916 585
R476 B.n914 B.n22 585
R477 B.n25 B.n22 585
R478 B.n913 B.n912 585
R479 B.n912 B.n911 585
R480 B.n24 B.n23 585
R481 B.n910 B.n24 585
R482 B.n908 B.n907 585
R483 B.n909 B.n908 585
R484 B.n906 B.n30 585
R485 B.n30 B.n29 585
R486 B.n905 B.n904 585
R487 B.n904 B.n903 585
R488 B.n32 B.n31 585
R489 B.n902 B.n32 585
R490 B.n900 B.n899 585
R491 B.n901 B.n900 585
R492 B.n898 B.n37 585
R493 B.n37 B.n36 585
R494 B.n897 B.n896 585
R495 B.n896 B.n895 585
R496 B.n39 B.n38 585
R497 B.n894 B.n39 585
R498 B.n892 B.n891 585
R499 B.n893 B.n892 585
R500 B.n890 B.n44 585
R501 B.n44 B.n43 585
R502 B.n889 B.n888 585
R503 B.n888 B.n887 585
R504 B.n46 B.n45 585
R505 B.n886 B.n46 585
R506 B.n884 B.n883 585
R507 B.n885 B.n884 585
R508 B.n882 B.n50 585
R509 B.n53 B.n50 585
R510 B.n881 B.n880 585
R511 B.n880 B.n879 585
R512 B.n52 B.n51 585
R513 B.n878 B.n52 585
R514 B.n876 B.n875 585
R515 B.n877 B.n876 585
R516 B.n874 B.n58 585
R517 B.n58 B.n57 585
R518 B.n873 B.n872 585
R519 B.n872 B.n871 585
R520 B.n60 B.n59 585
R521 B.n870 B.n60 585
R522 B.n868 B.n867 585
R523 B.n869 B.n868 585
R524 B.n866 B.n65 585
R525 B.n65 B.n64 585
R526 B.n865 B.n864 585
R527 B.n864 B.n863 585
R528 B.n67 B.n66 585
R529 B.n862 B.n67 585
R530 B.n860 B.n859 585
R531 B.n861 B.n860 585
R532 B.n858 B.n72 585
R533 B.n72 B.n71 585
R534 B.n857 B.n856 585
R535 B.n856 B.n855 585
R536 B.n74 B.n73 585
R537 B.n854 B.n74 585
R538 B.n852 B.n851 585
R539 B.n853 B.n852 585
R540 B.n937 B.n936 585
R541 B.n936 B.n935 585
R542 B.n469 B.n215 492.5
R543 B.n852 B.n79 492.5
R544 B.n471 B.n213 492.5
R545 B.n651 B.n77 492.5
R546 B.n246 B.t14 408.135
R547 B.n238 B.t21 408.135
R548 B.n102 B.t18 408.135
R549 B.n110 B.t10 408.135
R550 B.n246 B.t17 340.729
R551 B.n110 B.t12 340.729
R552 B.n238 B.t23 340.729
R553 B.n102 B.t19 340.729
R554 B.n247 B.t16 303.688
R555 B.n111 B.t13 303.688
R556 B.n239 B.t22 303.688
R557 B.n103 B.t20 303.688
R558 B.n652 B.n78 256.663
R559 B.n654 B.n78 256.663
R560 B.n660 B.n78 256.663
R561 B.n662 B.n78 256.663
R562 B.n668 B.n78 256.663
R563 B.n670 B.n78 256.663
R564 B.n676 B.n78 256.663
R565 B.n678 B.n78 256.663
R566 B.n684 B.n78 256.663
R567 B.n686 B.n78 256.663
R568 B.n692 B.n78 256.663
R569 B.n694 B.n78 256.663
R570 B.n700 B.n78 256.663
R571 B.n702 B.n78 256.663
R572 B.n708 B.n78 256.663
R573 B.n710 B.n78 256.663
R574 B.n716 B.n78 256.663
R575 B.n718 B.n78 256.663
R576 B.n724 B.n78 256.663
R577 B.n726 B.n78 256.663
R578 B.n732 B.n78 256.663
R579 B.n734 B.n78 256.663
R580 B.n740 B.n78 256.663
R581 B.n742 B.n78 256.663
R582 B.n748 B.n78 256.663
R583 B.n750 B.n78 256.663
R584 B.n756 B.n78 256.663
R585 B.n758 B.n78 256.663
R586 B.n765 B.n78 256.663
R587 B.n767 B.n78 256.663
R588 B.n773 B.n78 256.663
R589 B.n775 B.n78 256.663
R590 B.n781 B.n78 256.663
R591 B.n783 B.n78 256.663
R592 B.n789 B.n78 256.663
R593 B.n791 B.n78 256.663
R594 B.n797 B.n78 256.663
R595 B.n799 B.n78 256.663
R596 B.n805 B.n78 256.663
R597 B.n807 B.n78 256.663
R598 B.n813 B.n78 256.663
R599 B.n815 B.n78 256.663
R600 B.n821 B.n78 256.663
R601 B.n823 B.n78 256.663
R602 B.n829 B.n78 256.663
R603 B.n831 B.n78 256.663
R604 B.n837 B.n78 256.663
R605 B.n839 B.n78 256.663
R606 B.n845 B.n78 256.663
R607 B.n847 B.n78 256.663
R608 B.n464 B.n214 256.663
R609 B.n217 B.n214 256.663
R610 B.n457 B.n214 256.663
R611 B.n451 B.n214 256.663
R612 B.n449 B.n214 256.663
R613 B.n443 B.n214 256.663
R614 B.n441 B.n214 256.663
R615 B.n435 B.n214 256.663
R616 B.n433 B.n214 256.663
R617 B.n427 B.n214 256.663
R618 B.n425 B.n214 256.663
R619 B.n419 B.n214 256.663
R620 B.n417 B.n214 256.663
R621 B.n411 B.n214 256.663
R622 B.n409 B.n214 256.663
R623 B.n403 B.n214 256.663
R624 B.n401 B.n214 256.663
R625 B.n395 B.n214 256.663
R626 B.n393 B.n214 256.663
R627 B.n387 B.n214 256.663
R628 B.n385 B.n214 256.663
R629 B.n379 B.n214 256.663
R630 B.n241 B.n214 256.663
R631 B.n373 B.n214 256.663
R632 B.n367 B.n214 256.663
R633 B.n365 B.n214 256.663
R634 B.n359 B.n214 256.663
R635 B.n249 B.n214 256.663
R636 B.n353 B.n214 256.663
R637 B.n347 B.n214 256.663
R638 B.n345 B.n214 256.663
R639 B.n339 B.n214 256.663
R640 B.n337 B.n214 256.663
R641 B.n331 B.n214 256.663
R642 B.n329 B.n214 256.663
R643 B.n323 B.n214 256.663
R644 B.n321 B.n214 256.663
R645 B.n315 B.n214 256.663
R646 B.n313 B.n214 256.663
R647 B.n307 B.n214 256.663
R648 B.n305 B.n214 256.663
R649 B.n299 B.n214 256.663
R650 B.n297 B.n214 256.663
R651 B.n291 B.n214 256.663
R652 B.n289 B.n214 256.663
R653 B.n283 B.n214 256.663
R654 B.n281 B.n214 256.663
R655 B.n275 B.n214 256.663
R656 B.n273 B.n214 256.663
R657 B.n469 B.n209 163.367
R658 B.n477 B.n209 163.367
R659 B.n477 B.n207 163.367
R660 B.n481 B.n207 163.367
R661 B.n481 B.n201 163.367
R662 B.n489 B.n201 163.367
R663 B.n489 B.n199 163.367
R664 B.n493 B.n199 163.367
R665 B.n493 B.n193 163.367
R666 B.n501 B.n193 163.367
R667 B.n501 B.n191 163.367
R668 B.n505 B.n191 163.367
R669 B.n505 B.n185 163.367
R670 B.n514 B.n185 163.367
R671 B.n514 B.n183 163.367
R672 B.n518 B.n183 163.367
R673 B.n518 B.n178 163.367
R674 B.n526 B.n178 163.367
R675 B.n526 B.n176 163.367
R676 B.n530 B.n176 163.367
R677 B.n530 B.n170 163.367
R678 B.n538 B.n170 163.367
R679 B.n538 B.n168 163.367
R680 B.n542 B.n168 163.367
R681 B.n542 B.n162 163.367
R682 B.n550 B.n162 163.367
R683 B.n550 B.n160 163.367
R684 B.n554 B.n160 163.367
R685 B.n554 B.n154 163.367
R686 B.n563 B.n154 163.367
R687 B.n563 B.n152 163.367
R688 B.n567 B.n152 163.367
R689 B.n567 B.n147 163.367
R690 B.n575 B.n147 163.367
R691 B.n575 B.n145 163.367
R692 B.n579 B.n145 163.367
R693 B.n579 B.n139 163.367
R694 B.n588 B.n139 163.367
R695 B.n588 B.n137 163.367
R696 B.n592 B.n137 163.367
R697 B.n592 B.n2 163.367
R698 B.n936 B.n2 163.367
R699 B.n936 B.n3 163.367
R700 B.n932 B.n3 163.367
R701 B.n932 B.n9 163.367
R702 B.n928 B.n9 163.367
R703 B.n928 B.n11 163.367
R704 B.n924 B.n11 163.367
R705 B.n924 B.n16 163.367
R706 B.n920 B.n16 163.367
R707 B.n920 B.n18 163.367
R708 B.n916 B.n18 163.367
R709 B.n916 B.n22 163.367
R710 B.n912 B.n22 163.367
R711 B.n912 B.n24 163.367
R712 B.n908 B.n24 163.367
R713 B.n908 B.n30 163.367
R714 B.n904 B.n30 163.367
R715 B.n904 B.n32 163.367
R716 B.n900 B.n32 163.367
R717 B.n900 B.n37 163.367
R718 B.n896 B.n37 163.367
R719 B.n896 B.n39 163.367
R720 B.n892 B.n39 163.367
R721 B.n892 B.n44 163.367
R722 B.n888 B.n44 163.367
R723 B.n888 B.n46 163.367
R724 B.n884 B.n46 163.367
R725 B.n884 B.n50 163.367
R726 B.n880 B.n50 163.367
R727 B.n880 B.n52 163.367
R728 B.n876 B.n52 163.367
R729 B.n876 B.n58 163.367
R730 B.n872 B.n58 163.367
R731 B.n872 B.n60 163.367
R732 B.n868 B.n60 163.367
R733 B.n868 B.n65 163.367
R734 B.n864 B.n65 163.367
R735 B.n864 B.n67 163.367
R736 B.n860 B.n67 163.367
R737 B.n860 B.n72 163.367
R738 B.n856 B.n72 163.367
R739 B.n856 B.n74 163.367
R740 B.n852 B.n74 163.367
R741 B.n465 B.n463 163.367
R742 B.n463 B.n462 163.367
R743 B.n459 B.n458 163.367
R744 B.n456 B.n219 163.367
R745 B.n452 B.n450 163.367
R746 B.n448 B.n221 163.367
R747 B.n444 B.n442 163.367
R748 B.n440 B.n223 163.367
R749 B.n436 B.n434 163.367
R750 B.n432 B.n225 163.367
R751 B.n428 B.n426 163.367
R752 B.n424 B.n227 163.367
R753 B.n420 B.n418 163.367
R754 B.n416 B.n229 163.367
R755 B.n412 B.n410 163.367
R756 B.n408 B.n231 163.367
R757 B.n404 B.n402 163.367
R758 B.n400 B.n233 163.367
R759 B.n396 B.n394 163.367
R760 B.n392 B.n235 163.367
R761 B.n388 B.n386 163.367
R762 B.n384 B.n237 163.367
R763 B.n380 B.n378 163.367
R764 B.n375 B.n374 163.367
R765 B.n372 B.n243 163.367
R766 B.n368 B.n366 163.367
R767 B.n364 B.n245 163.367
R768 B.n360 B.n358 163.367
R769 B.n355 B.n354 163.367
R770 B.n352 B.n251 163.367
R771 B.n348 B.n346 163.367
R772 B.n344 B.n253 163.367
R773 B.n340 B.n338 163.367
R774 B.n336 B.n255 163.367
R775 B.n332 B.n330 163.367
R776 B.n328 B.n257 163.367
R777 B.n324 B.n322 163.367
R778 B.n320 B.n259 163.367
R779 B.n316 B.n314 163.367
R780 B.n312 B.n261 163.367
R781 B.n308 B.n306 163.367
R782 B.n304 B.n263 163.367
R783 B.n300 B.n298 163.367
R784 B.n296 B.n265 163.367
R785 B.n292 B.n290 163.367
R786 B.n288 B.n267 163.367
R787 B.n284 B.n282 163.367
R788 B.n280 B.n269 163.367
R789 B.n276 B.n274 163.367
R790 B.n272 B.n213 163.367
R791 B.n471 B.n211 163.367
R792 B.n475 B.n211 163.367
R793 B.n475 B.n205 163.367
R794 B.n483 B.n205 163.367
R795 B.n483 B.n203 163.367
R796 B.n487 B.n203 163.367
R797 B.n487 B.n197 163.367
R798 B.n495 B.n197 163.367
R799 B.n495 B.n195 163.367
R800 B.n499 B.n195 163.367
R801 B.n499 B.n189 163.367
R802 B.n507 B.n189 163.367
R803 B.n507 B.n187 163.367
R804 B.n511 B.n187 163.367
R805 B.n511 B.n182 163.367
R806 B.n520 B.n182 163.367
R807 B.n520 B.n180 163.367
R808 B.n524 B.n180 163.367
R809 B.n524 B.n174 163.367
R810 B.n532 B.n174 163.367
R811 B.n532 B.n172 163.367
R812 B.n536 B.n172 163.367
R813 B.n536 B.n166 163.367
R814 B.n544 B.n166 163.367
R815 B.n544 B.n164 163.367
R816 B.n548 B.n164 163.367
R817 B.n548 B.n158 163.367
R818 B.n556 B.n158 163.367
R819 B.n556 B.n156 163.367
R820 B.n560 B.n156 163.367
R821 B.n560 B.n151 163.367
R822 B.n569 B.n151 163.367
R823 B.n569 B.n149 163.367
R824 B.n573 B.n149 163.367
R825 B.n573 B.n142 163.367
R826 B.n581 B.n142 163.367
R827 B.n581 B.n140 163.367
R828 B.n586 B.n140 163.367
R829 B.n586 B.n135 163.367
R830 B.n594 B.n135 163.367
R831 B.n595 B.n594 163.367
R832 B.n595 B.n5 163.367
R833 B.n6 B.n5 163.367
R834 B.n7 B.n6 163.367
R835 B.n600 B.n7 163.367
R836 B.n600 B.n12 163.367
R837 B.n13 B.n12 163.367
R838 B.n14 B.n13 163.367
R839 B.n605 B.n14 163.367
R840 B.n605 B.n19 163.367
R841 B.n20 B.n19 163.367
R842 B.n21 B.n20 163.367
R843 B.n610 B.n21 163.367
R844 B.n610 B.n26 163.367
R845 B.n27 B.n26 163.367
R846 B.n28 B.n27 163.367
R847 B.n615 B.n28 163.367
R848 B.n615 B.n33 163.367
R849 B.n34 B.n33 163.367
R850 B.n35 B.n34 163.367
R851 B.n620 B.n35 163.367
R852 B.n620 B.n40 163.367
R853 B.n41 B.n40 163.367
R854 B.n42 B.n41 163.367
R855 B.n625 B.n42 163.367
R856 B.n625 B.n47 163.367
R857 B.n48 B.n47 163.367
R858 B.n49 B.n48 163.367
R859 B.n630 B.n49 163.367
R860 B.n630 B.n54 163.367
R861 B.n55 B.n54 163.367
R862 B.n56 B.n55 163.367
R863 B.n635 B.n56 163.367
R864 B.n635 B.n61 163.367
R865 B.n62 B.n61 163.367
R866 B.n63 B.n62 163.367
R867 B.n640 B.n63 163.367
R868 B.n640 B.n68 163.367
R869 B.n69 B.n68 163.367
R870 B.n70 B.n69 163.367
R871 B.n645 B.n70 163.367
R872 B.n645 B.n75 163.367
R873 B.n76 B.n75 163.367
R874 B.n77 B.n76 163.367
R875 B.n848 B.n846 163.367
R876 B.n844 B.n81 163.367
R877 B.n840 B.n838 163.367
R878 B.n836 B.n83 163.367
R879 B.n832 B.n830 163.367
R880 B.n828 B.n85 163.367
R881 B.n824 B.n822 163.367
R882 B.n820 B.n87 163.367
R883 B.n816 B.n814 163.367
R884 B.n812 B.n89 163.367
R885 B.n808 B.n806 163.367
R886 B.n804 B.n91 163.367
R887 B.n800 B.n798 163.367
R888 B.n796 B.n93 163.367
R889 B.n792 B.n790 163.367
R890 B.n788 B.n95 163.367
R891 B.n784 B.n782 163.367
R892 B.n780 B.n97 163.367
R893 B.n776 B.n774 163.367
R894 B.n772 B.n99 163.367
R895 B.n768 B.n766 163.367
R896 B.n764 B.n101 163.367
R897 B.n759 B.n757 163.367
R898 B.n755 B.n105 163.367
R899 B.n751 B.n749 163.367
R900 B.n747 B.n107 163.367
R901 B.n743 B.n741 163.367
R902 B.n739 B.n109 163.367
R903 B.n735 B.n733 163.367
R904 B.n731 B.n114 163.367
R905 B.n727 B.n725 163.367
R906 B.n723 B.n116 163.367
R907 B.n719 B.n717 163.367
R908 B.n715 B.n118 163.367
R909 B.n711 B.n709 163.367
R910 B.n707 B.n120 163.367
R911 B.n703 B.n701 163.367
R912 B.n699 B.n122 163.367
R913 B.n695 B.n693 163.367
R914 B.n691 B.n124 163.367
R915 B.n687 B.n685 163.367
R916 B.n683 B.n126 163.367
R917 B.n679 B.n677 163.367
R918 B.n675 B.n128 163.367
R919 B.n671 B.n669 163.367
R920 B.n667 B.n130 163.367
R921 B.n663 B.n661 163.367
R922 B.n659 B.n132 163.367
R923 B.n655 B.n653 163.367
R924 B.n464 B.n215 71.676
R925 B.n462 B.n217 71.676
R926 B.n458 B.n457 71.676
R927 B.n451 B.n219 71.676
R928 B.n450 B.n449 71.676
R929 B.n443 B.n221 71.676
R930 B.n442 B.n441 71.676
R931 B.n435 B.n223 71.676
R932 B.n434 B.n433 71.676
R933 B.n427 B.n225 71.676
R934 B.n426 B.n425 71.676
R935 B.n419 B.n227 71.676
R936 B.n418 B.n417 71.676
R937 B.n411 B.n229 71.676
R938 B.n410 B.n409 71.676
R939 B.n403 B.n231 71.676
R940 B.n402 B.n401 71.676
R941 B.n395 B.n233 71.676
R942 B.n394 B.n393 71.676
R943 B.n387 B.n235 71.676
R944 B.n386 B.n385 71.676
R945 B.n379 B.n237 71.676
R946 B.n378 B.n241 71.676
R947 B.n374 B.n373 71.676
R948 B.n367 B.n243 71.676
R949 B.n366 B.n365 71.676
R950 B.n359 B.n245 71.676
R951 B.n358 B.n249 71.676
R952 B.n354 B.n353 71.676
R953 B.n347 B.n251 71.676
R954 B.n346 B.n345 71.676
R955 B.n339 B.n253 71.676
R956 B.n338 B.n337 71.676
R957 B.n331 B.n255 71.676
R958 B.n330 B.n329 71.676
R959 B.n323 B.n257 71.676
R960 B.n322 B.n321 71.676
R961 B.n315 B.n259 71.676
R962 B.n314 B.n313 71.676
R963 B.n307 B.n261 71.676
R964 B.n306 B.n305 71.676
R965 B.n299 B.n263 71.676
R966 B.n298 B.n297 71.676
R967 B.n291 B.n265 71.676
R968 B.n290 B.n289 71.676
R969 B.n283 B.n267 71.676
R970 B.n282 B.n281 71.676
R971 B.n275 B.n269 71.676
R972 B.n274 B.n273 71.676
R973 B.n847 B.n79 71.676
R974 B.n846 B.n845 71.676
R975 B.n839 B.n81 71.676
R976 B.n838 B.n837 71.676
R977 B.n831 B.n83 71.676
R978 B.n830 B.n829 71.676
R979 B.n823 B.n85 71.676
R980 B.n822 B.n821 71.676
R981 B.n815 B.n87 71.676
R982 B.n814 B.n813 71.676
R983 B.n807 B.n89 71.676
R984 B.n806 B.n805 71.676
R985 B.n799 B.n91 71.676
R986 B.n798 B.n797 71.676
R987 B.n791 B.n93 71.676
R988 B.n790 B.n789 71.676
R989 B.n783 B.n95 71.676
R990 B.n782 B.n781 71.676
R991 B.n775 B.n97 71.676
R992 B.n774 B.n773 71.676
R993 B.n767 B.n99 71.676
R994 B.n766 B.n765 71.676
R995 B.n758 B.n101 71.676
R996 B.n757 B.n756 71.676
R997 B.n750 B.n105 71.676
R998 B.n749 B.n748 71.676
R999 B.n742 B.n107 71.676
R1000 B.n741 B.n740 71.676
R1001 B.n734 B.n109 71.676
R1002 B.n733 B.n732 71.676
R1003 B.n726 B.n114 71.676
R1004 B.n725 B.n724 71.676
R1005 B.n718 B.n116 71.676
R1006 B.n717 B.n716 71.676
R1007 B.n710 B.n118 71.676
R1008 B.n709 B.n708 71.676
R1009 B.n702 B.n120 71.676
R1010 B.n701 B.n700 71.676
R1011 B.n694 B.n122 71.676
R1012 B.n693 B.n692 71.676
R1013 B.n686 B.n124 71.676
R1014 B.n685 B.n684 71.676
R1015 B.n678 B.n126 71.676
R1016 B.n677 B.n676 71.676
R1017 B.n670 B.n128 71.676
R1018 B.n669 B.n668 71.676
R1019 B.n662 B.n130 71.676
R1020 B.n661 B.n660 71.676
R1021 B.n654 B.n132 71.676
R1022 B.n653 B.n652 71.676
R1023 B.n652 B.n651 71.676
R1024 B.n655 B.n654 71.676
R1025 B.n660 B.n659 71.676
R1026 B.n663 B.n662 71.676
R1027 B.n668 B.n667 71.676
R1028 B.n671 B.n670 71.676
R1029 B.n676 B.n675 71.676
R1030 B.n679 B.n678 71.676
R1031 B.n684 B.n683 71.676
R1032 B.n687 B.n686 71.676
R1033 B.n692 B.n691 71.676
R1034 B.n695 B.n694 71.676
R1035 B.n700 B.n699 71.676
R1036 B.n703 B.n702 71.676
R1037 B.n708 B.n707 71.676
R1038 B.n711 B.n710 71.676
R1039 B.n716 B.n715 71.676
R1040 B.n719 B.n718 71.676
R1041 B.n724 B.n723 71.676
R1042 B.n727 B.n726 71.676
R1043 B.n732 B.n731 71.676
R1044 B.n735 B.n734 71.676
R1045 B.n740 B.n739 71.676
R1046 B.n743 B.n742 71.676
R1047 B.n748 B.n747 71.676
R1048 B.n751 B.n750 71.676
R1049 B.n756 B.n755 71.676
R1050 B.n759 B.n758 71.676
R1051 B.n765 B.n764 71.676
R1052 B.n768 B.n767 71.676
R1053 B.n773 B.n772 71.676
R1054 B.n776 B.n775 71.676
R1055 B.n781 B.n780 71.676
R1056 B.n784 B.n783 71.676
R1057 B.n789 B.n788 71.676
R1058 B.n792 B.n791 71.676
R1059 B.n797 B.n796 71.676
R1060 B.n800 B.n799 71.676
R1061 B.n805 B.n804 71.676
R1062 B.n808 B.n807 71.676
R1063 B.n813 B.n812 71.676
R1064 B.n816 B.n815 71.676
R1065 B.n821 B.n820 71.676
R1066 B.n824 B.n823 71.676
R1067 B.n829 B.n828 71.676
R1068 B.n832 B.n831 71.676
R1069 B.n837 B.n836 71.676
R1070 B.n840 B.n839 71.676
R1071 B.n845 B.n844 71.676
R1072 B.n848 B.n847 71.676
R1073 B.n465 B.n464 71.676
R1074 B.n459 B.n217 71.676
R1075 B.n457 B.n456 71.676
R1076 B.n452 B.n451 71.676
R1077 B.n449 B.n448 71.676
R1078 B.n444 B.n443 71.676
R1079 B.n441 B.n440 71.676
R1080 B.n436 B.n435 71.676
R1081 B.n433 B.n432 71.676
R1082 B.n428 B.n427 71.676
R1083 B.n425 B.n424 71.676
R1084 B.n420 B.n419 71.676
R1085 B.n417 B.n416 71.676
R1086 B.n412 B.n411 71.676
R1087 B.n409 B.n408 71.676
R1088 B.n404 B.n403 71.676
R1089 B.n401 B.n400 71.676
R1090 B.n396 B.n395 71.676
R1091 B.n393 B.n392 71.676
R1092 B.n388 B.n387 71.676
R1093 B.n385 B.n384 71.676
R1094 B.n380 B.n379 71.676
R1095 B.n375 B.n241 71.676
R1096 B.n373 B.n372 71.676
R1097 B.n368 B.n367 71.676
R1098 B.n365 B.n364 71.676
R1099 B.n360 B.n359 71.676
R1100 B.n355 B.n249 71.676
R1101 B.n353 B.n352 71.676
R1102 B.n348 B.n347 71.676
R1103 B.n345 B.n344 71.676
R1104 B.n340 B.n339 71.676
R1105 B.n337 B.n336 71.676
R1106 B.n332 B.n331 71.676
R1107 B.n329 B.n328 71.676
R1108 B.n324 B.n323 71.676
R1109 B.n321 B.n320 71.676
R1110 B.n316 B.n315 71.676
R1111 B.n313 B.n312 71.676
R1112 B.n308 B.n307 71.676
R1113 B.n305 B.n304 71.676
R1114 B.n300 B.n299 71.676
R1115 B.n297 B.n296 71.676
R1116 B.n292 B.n291 71.676
R1117 B.n289 B.n288 71.676
R1118 B.n284 B.n283 71.676
R1119 B.n281 B.n280 71.676
R1120 B.n276 B.n275 71.676
R1121 B.n273 B.n272 71.676
R1122 B.n470 B.n214 65.8404
R1123 B.n853 B.n78 65.8404
R1124 B.n248 B.n247 59.5399
R1125 B.n240 B.n239 59.5399
R1126 B.n761 B.n103 59.5399
R1127 B.n112 B.n111 59.5399
R1128 B.n470 B.n210 40.3348
R1129 B.n476 B.n210 40.3348
R1130 B.n476 B.n206 40.3348
R1131 B.n482 B.n206 40.3348
R1132 B.n482 B.n202 40.3348
R1133 B.n488 B.n202 40.3348
R1134 B.n494 B.n198 40.3348
R1135 B.n494 B.n194 40.3348
R1136 B.n500 B.n194 40.3348
R1137 B.n500 B.n190 40.3348
R1138 B.n506 B.n190 40.3348
R1139 B.n506 B.n186 40.3348
R1140 B.n513 B.n186 40.3348
R1141 B.n513 B.n512 40.3348
R1142 B.n519 B.n179 40.3348
R1143 B.n525 B.n179 40.3348
R1144 B.n525 B.n175 40.3348
R1145 B.n531 B.n175 40.3348
R1146 B.n537 B.n171 40.3348
R1147 B.n537 B.n167 40.3348
R1148 B.n543 B.n167 40.3348
R1149 B.n543 B.n163 40.3348
R1150 B.n549 B.n163 40.3348
R1151 B.n555 B.n159 40.3348
R1152 B.n555 B.n155 40.3348
R1153 B.n562 B.n155 40.3348
R1154 B.n562 B.n561 40.3348
R1155 B.n568 B.n148 40.3348
R1156 B.n574 B.n148 40.3348
R1157 B.n574 B.n143 40.3348
R1158 B.n580 B.n143 40.3348
R1159 B.n580 B.n144 40.3348
R1160 B.n587 B.n136 40.3348
R1161 B.n593 B.n136 40.3348
R1162 B.n593 B.n4 40.3348
R1163 B.n935 B.n4 40.3348
R1164 B.n935 B.n934 40.3348
R1165 B.n934 B.n933 40.3348
R1166 B.n933 B.n8 40.3348
R1167 B.n927 B.n8 40.3348
R1168 B.n926 B.n925 40.3348
R1169 B.n925 B.n15 40.3348
R1170 B.n919 B.n15 40.3348
R1171 B.n919 B.n918 40.3348
R1172 B.n918 B.n917 40.3348
R1173 B.n911 B.n25 40.3348
R1174 B.n911 B.n910 40.3348
R1175 B.n910 B.n909 40.3348
R1176 B.n909 B.n29 40.3348
R1177 B.n903 B.n902 40.3348
R1178 B.n902 B.n901 40.3348
R1179 B.n901 B.n36 40.3348
R1180 B.n895 B.n36 40.3348
R1181 B.n895 B.n894 40.3348
R1182 B.n893 B.n43 40.3348
R1183 B.n887 B.n43 40.3348
R1184 B.n887 B.n886 40.3348
R1185 B.n886 B.n885 40.3348
R1186 B.n879 B.n53 40.3348
R1187 B.n879 B.n878 40.3348
R1188 B.n878 B.n877 40.3348
R1189 B.n877 B.n57 40.3348
R1190 B.n871 B.n57 40.3348
R1191 B.n871 B.n870 40.3348
R1192 B.n870 B.n869 40.3348
R1193 B.n869 B.n64 40.3348
R1194 B.n863 B.n862 40.3348
R1195 B.n862 B.n861 40.3348
R1196 B.n861 B.n71 40.3348
R1197 B.n855 B.n71 40.3348
R1198 B.n855 B.n854 40.3348
R1199 B.n854 B.n853 40.3348
R1200 B.n561 B.t8 39.1485
R1201 B.n25 B.t2 39.1485
R1202 B.n247 B.n246 37.0429
R1203 B.n239 B.n238 37.0429
R1204 B.n103 B.n102 37.0429
R1205 B.n111 B.n110 37.0429
R1206 B.n519 B.t0 35.5896
R1207 B.n885 B.t6 35.5896
R1208 B.n851 B.n850 32.0005
R1209 B.n650 B.n649 32.0005
R1210 B.n472 B.n212 32.0005
R1211 B.n468 B.n467 32.0005
R1212 B.n531 B.t4 29.6581
R1213 B.t9 B.n893 29.6581
R1214 B.t15 B.n198 28.4718
R1215 B.t11 B.n64 28.4718
R1216 B.t5 B.n159 26.0992
R1217 B.t1 B.n29 26.0992
R1218 B.n144 B.t3 23.7266
R1219 B.t7 B.n926 23.7266
R1220 B B.n937 18.0485
R1221 B.n587 B.t3 16.6087
R1222 B.n927 B.t7 16.6087
R1223 B.n549 B.t5 14.2361
R1224 B.n903 B.t1 14.2361
R1225 B.n488 B.t15 11.8635
R1226 B.n863 B.t11 11.8635
R1227 B.t4 B.n171 10.6772
R1228 B.n894 B.t9 10.6772
R1229 B.n850 B.n849 10.6151
R1230 B.n849 B.n80 10.6151
R1231 B.n843 B.n80 10.6151
R1232 B.n843 B.n842 10.6151
R1233 B.n842 B.n841 10.6151
R1234 B.n841 B.n82 10.6151
R1235 B.n835 B.n82 10.6151
R1236 B.n835 B.n834 10.6151
R1237 B.n834 B.n833 10.6151
R1238 B.n833 B.n84 10.6151
R1239 B.n827 B.n84 10.6151
R1240 B.n827 B.n826 10.6151
R1241 B.n826 B.n825 10.6151
R1242 B.n825 B.n86 10.6151
R1243 B.n819 B.n86 10.6151
R1244 B.n819 B.n818 10.6151
R1245 B.n818 B.n817 10.6151
R1246 B.n817 B.n88 10.6151
R1247 B.n811 B.n88 10.6151
R1248 B.n811 B.n810 10.6151
R1249 B.n810 B.n809 10.6151
R1250 B.n809 B.n90 10.6151
R1251 B.n803 B.n90 10.6151
R1252 B.n803 B.n802 10.6151
R1253 B.n802 B.n801 10.6151
R1254 B.n801 B.n92 10.6151
R1255 B.n795 B.n92 10.6151
R1256 B.n795 B.n794 10.6151
R1257 B.n794 B.n793 10.6151
R1258 B.n793 B.n94 10.6151
R1259 B.n787 B.n94 10.6151
R1260 B.n787 B.n786 10.6151
R1261 B.n786 B.n785 10.6151
R1262 B.n785 B.n96 10.6151
R1263 B.n779 B.n96 10.6151
R1264 B.n779 B.n778 10.6151
R1265 B.n778 B.n777 10.6151
R1266 B.n777 B.n98 10.6151
R1267 B.n771 B.n98 10.6151
R1268 B.n771 B.n770 10.6151
R1269 B.n770 B.n769 10.6151
R1270 B.n769 B.n100 10.6151
R1271 B.n763 B.n100 10.6151
R1272 B.n763 B.n762 10.6151
R1273 B.n760 B.n104 10.6151
R1274 B.n754 B.n104 10.6151
R1275 B.n754 B.n753 10.6151
R1276 B.n753 B.n752 10.6151
R1277 B.n752 B.n106 10.6151
R1278 B.n746 B.n106 10.6151
R1279 B.n746 B.n745 10.6151
R1280 B.n745 B.n744 10.6151
R1281 B.n744 B.n108 10.6151
R1282 B.n738 B.n737 10.6151
R1283 B.n737 B.n736 10.6151
R1284 B.n736 B.n113 10.6151
R1285 B.n730 B.n113 10.6151
R1286 B.n730 B.n729 10.6151
R1287 B.n729 B.n728 10.6151
R1288 B.n728 B.n115 10.6151
R1289 B.n722 B.n115 10.6151
R1290 B.n722 B.n721 10.6151
R1291 B.n721 B.n720 10.6151
R1292 B.n720 B.n117 10.6151
R1293 B.n714 B.n117 10.6151
R1294 B.n714 B.n713 10.6151
R1295 B.n713 B.n712 10.6151
R1296 B.n712 B.n119 10.6151
R1297 B.n706 B.n119 10.6151
R1298 B.n706 B.n705 10.6151
R1299 B.n705 B.n704 10.6151
R1300 B.n704 B.n121 10.6151
R1301 B.n698 B.n121 10.6151
R1302 B.n698 B.n697 10.6151
R1303 B.n697 B.n696 10.6151
R1304 B.n696 B.n123 10.6151
R1305 B.n690 B.n123 10.6151
R1306 B.n690 B.n689 10.6151
R1307 B.n689 B.n688 10.6151
R1308 B.n688 B.n125 10.6151
R1309 B.n682 B.n125 10.6151
R1310 B.n682 B.n681 10.6151
R1311 B.n681 B.n680 10.6151
R1312 B.n680 B.n127 10.6151
R1313 B.n674 B.n127 10.6151
R1314 B.n674 B.n673 10.6151
R1315 B.n673 B.n672 10.6151
R1316 B.n672 B.n129 10.6151
R1317 B.n666 B.n129 10.6151
R1318 B.n666 B.n665 10.6151
R1319 B.n665 B.n664 10.6151
R1320 B.n664 B.n131 10.6151
R1321 B.n658 B.n131 10.6151
R1322 B.n658 B.n657 10.6151
R1323 B.n657 B.n656 10.6151
R1324 B.n656 B.n133 10.6151
R1325 B.n650 B.n133 10.6151
R1326 B.n473 B.n472 10.6151
R1327 B.n474 B.n473 10.6151
R1328 B.n474 B.n204 10.6151
R1329 B.n484 B.n204 10.6151
R1330 B.n485 B.n484 10.6151
R1331 B.n486 B.n485 10.6151
R1332 B.n486 B.n196 10.6151
R1333 B.n496 B.n196 10.6151
R1334 B.n497 B.n496 10.6151
R1335 B.n498 B.n497 10.6151
R1336 B.n498 B.n188 10.6151
R1337 B.n508 B.n188 10.6151
R1338 B.n509 B.n508 10.6151
R1339 B.n510 B.n509 10.6151
R1340 B.n510 B.n181 10.6151
R1341 B.n521 B.n181 10.6151
R1342 B.n522 B.n521 10.6151
R1343 B.n523 B.n522 10.6151
R1344 B.n523 B.n173 10.6151
R1345 B.n533 B.n173 10.6151
R1346 B.n534 B.n533 10.6151
R1347 B.n535 B.n534 10.6151
R1348 B.n535 B.n165 10.6151
R1349 B.n545 B.n165 10.6151
R1350 B.n546 B.n545 10.6151
R1351 B.n547 B.n546 10.6151
R1352 B.n547 B.n157 10.6151
R1353 B.n557 B.n157 10.6151
R1354 B.n558 B.n557 10.6151
R1355 B.n559 B.n558 10.6151
R1356 B.n559 B.n150 10.6151
R1357 B.n570 B.n150 10.6151
R1358 B.n571 B.n570 10.6151
R1359 B.n572 B.n571 10.6151
R1360 B.n572 B.n141 10.6151
R1361 B.n582 B.n141 10.6151
R1362 B.n583 B.n582 10.6151
R1363 B.n585 B.n583 10.6151
R1364 B.n585 B.n584 10.6151
R1365 B.n584 B.n134 10.6151
R1366 B.n596 B.n134 10.6151
R1367 B.n597 B.n596 10.6151
R1368 B.n598 B.n597 10.6151
R1369 B.n599 B.n598 10.6151
R1370 B.n601 B.n599 10.6151
R1371 B.n602 B.n601 10.6151
R1372 B.n603 B.n602 10.6151
R1373 B.n604 B.n603 10.6151
R1374 B.n606 B.n604 10.6151
R1375 B.n607 B.n606 10.6151
R1376 B.n608 B.n607 10.6151
R1377 B.n609 B.n608 10.6151
R1378 B.n611 B.n609 10.6151
R1379 B.n612 B.n611 10.6151
R1380 B.n613 B.n612 10.6151
R1381 B.n614 B.n613 10.6151
R1382 B.n616 B.n614 10.6151
R1383 B.n617 B.n616 10.6151
R1384 B.n618 B.n617 10.6151
R1385 B.n619 B.n618 10.6151
R1386 B.n621 B.n619 10.6151
R1387 B.n622 B.n621 10.6151
R1388 B.n623 B.n622 10.6151
R1389 B.n624 B.n623 10.6151
R1390 B.n626 B.n624 10.6151
R1391 B.n627 B.n626 10.6151
R1392 B.n628 B.n627 10.6151
R1393 B.n629 B.n628 10.6151
R1394 B.n631 B.n629 10.6151
R1395 B.n632 B.n631 10.6151
R1396 B.n633 B.n632 10.6151
R1397 B.n634 B.n633 10.6151
R1398 B.n636 B.n634 10.6151
R1399 B.n637 B.n636 10.6151
R1400 B.n638 B.n637 10.6151
R1401 B.n639 B.n638 10.6151
R1402 B.n641 B.n639 10.6151
R1403 B.n642 B.n641 10.6151
R1404 B.n643 B.n642 10.6151
R1405 B.n644 B.n643 10.6151
R1406 B.n646 B.n644 10.6151
R1407 B.n647 B.n646 10.6151
R1408 B.n648 B.n647 10.6151
R1409 B.n649 B.n648 10.6151
R1410 B.n467 B.n466 10.6151
R1411 B.n466 B.n216 10.6151
R1412 B.n461 B.n216 10.6151
R1413 B.n461 B.n460 10.6151
R1414 B.n460 B.n218 10.6151
R1415 B.n455 B.n218 10.6151
R1416 B.n455 B.n454 10.6151
R1417 B.n454 B.n453 10.6151
R1418 B.n453 B.n220 10.6151
R1419 B.n447 B.n220 10.6151
R1420 B.n447 B.n446 10.6151
R1421 B.n446 B.n445 10.6151
R1422 B.n445 B.n222 10.6151
R1423 B.n439 B.n222 10.6151
R1424 B.n439 B.n438 10.6151
R1425 B.n438 B.n437 10.6151
R1426 B.n437 B.n224 10.6151
R1427 B.n431 B.n224 10.6151
R1428 B.n431 B.n430 10.6151
R1429 B.n430 B.n429 10.6151
R1430 B.n429 B.n226 10.6151
R1431 B.n423 B.n226 10.6151
R1432 B.n423 B.n422 10.6151
R1433 B.n422 B.n421 10.6151
R1434 B.n421 B.n228 10.6151
R1435 B.n415 B.n228 10.6151
R1436 B.n415 B.n414 10.6151
R1437 B.n414 B.n413 10.6151
R1438 B.n413 B.n230 10.6151
R1439 B.n407 B.n230 10.6151
R1440 B.n407 B.n406 10.6151
R1441 B.n406 B.n405 10.6151
R1442 B.n405 B.n232 10.6151
R1443 B.n399 B.n232 10.6151
R1444 B.n399 B.n398 10.6151
R1445 B.n398 B.n397 10.6151
R1446 B.n397 B.n234 10.6151
R1447 B.n391 B.n234 10.6151
R1448 B.n391 B.n390 10.6151
R1449 B.n390 B.n389 10.6151
R1450 B.n389 B.n236 10.6151
R1451 B.n383 B.n236 10.6151
R1452 B.n383 B.n382 10.6151
R1453 B.n382 B.n381 10.6151
R1454 B.n377 B.n376 10.6151
R1455 B.n376 B.n242 10.6151
R1456 B.n371 B.n242 10.6151
R1457 B.n371 B.n370 10.6151
R1458 B.n370 B.n369 10.6151
R1459 B.n369 B.n244 10.6151
R1460 B.n363 B.n244 10.6151
R1461 B.n363 B.n362 10.6151
R1462 B.n362 B.n361 10.6151
R1463 B.n357 B.n356 10.6151
R1464 B.n356 B.n250 10.6151
R1465 B.n351 B.n250 10.6151
R1466 B.n351 B.n350 10.6151
R1467 B.n350 B.n349 10.6151
R1468 B.n349 B.n252 10.6151
R1469 B.n343 B.n252 10.6151
R1470 B.n343 B.n342 10.6151
R1471 B.n342 B.n341 10.6151
R1472 B.n341 B.n254 10.6151
R1473 B.n335 B.n254 10.6151
R1474 B.n335 B.n334 10.6151
R1475 B.n334 B.n333 10.6151
R1476 B.n333 B.n256 10.6151
R1477 B.n327 B.n256 10.6151
R1478 B.n327 B.n326 10.6151
R1479 B.n326 B.n325 10.6151
R1480 B.n325 B.n258 10.6151
R1481 B.n319 B.n258 10.6151
R1482 B.n319 B.n318 10.6151
R1483 B.n318 B.n317 10.6151
R1484 B.n317 B.n260 10.6151
R1485 B.n311 B.n260 10.6151
R1486 B.n311 B.n310 10.6151
R1487 B.n310 B.n309 10.6151
R1488 B.n309 B.n262 10.6151
R1489 B.n303 B.n262 10.6151
R1490 B.n303 B.n302 10.6151
R1491 B.n302 B.n301 10.6151
R1492 B.n301 B.n264 10.6151
R1493 B.n295 B.n264 10.6151
R1494 B.n295 B.n294 10.6151
R1495 B.n294 B.n293 10.6151
R1496 B.n293 B.n266 10.6151
R1497 B.n287 B.n266 10.6151
R1498 B.n287 B.n286 10.6151
R1499 B.n286 B.n285 10.6151
R1500 B.n285 B.n268 10.6151
R1501 B.n279 B.n268 10.6151
R1502 B.n279 B.n278 10.6151
R1503 B.n278 B.n277 10.6151
R1504 B.n277 B.n270 10.6151
R1505 B.n271 B.n270 10.6151
R1506 B.n271 B.n212 10.6151
R1507 B.n468 B.n208 10.6151
R1508 B.n478 B.n208 10.6151
R1509 B.n479 B.n478 10.6151
R1510 B.n480 B.n479 10.6151
R1511 B.n480 B.n200 10.6151
R1512 B.n490 B.n200 10.6151
R1513 B.n491 B.n490 10.6151
R1514 B.n492 B.n491 10.6151
R1515 B.n492 B.n192 10.6151
R1516 B.n502 B.n192 10.6151
R1517 B.n503 B.n502 10.6151
R1518 B.n504 B.n503 10.6151
R1519 B.n504 B.n184 10.6151
R1520 B.n515 B.n184 10.6151
R1521 B.n516 B.n515 10.6151
R1522 B.n517 B.n516 10.6151
R1523 B.n517 B.n177 10.6151
R1524 B.n527 B.n177 10.6151
R1525 B.n528 B.n527 10.6151
R1526 B.n529 B.n528 10.6151
R1527 B.n529 B.n169 10.6151
R1528 B.n539 B.n169 10.6151
R1529 B.n540 B.n539 10.6151
R1530 B.n541 B.n540 10.6151
R1531 B.n541 B.n161 10.6151
R1532 B.n551 B.n161 10.6151
R1533 B.n552 B.n551 10.6151
R1534 B.n553 B.n552 10.6151
R1535 B.n553 B.n153 10.6151
R1536 B.n564 B.n153 10.6151
R1537 B.n565 B.n564 10.6151
R1538 B.n566 B.n565 10.6151
R1539 B.n566 B.n146 10.6151
R1540 B.n576 B.n146 10.6151
R1541 B.n577 B.n576 10.6151
R1542 B.n578 B.n577 10.6151
R1543 B.n578 B.n138 10.6151
R1544 B.n589 B.n138 10.6151
R1545 B.n590 B.n589 10.6151
R1546 B.n591 B.n590 10.6151
R1547 B.n591 B.n0 10.6151
R1548 B.n931 B.n1 10.6151
R1549 B.n931 B.n930 10.6151
R1550 B.n930 B.n929 10.6151
R1551 B.n929 B.n10 10.6151
R1552 B.n923 B.n10 10.6151
R1553 B.n923 B.n922 10.6151
R1554 B.n922 B.n921 10.6151
R1555 B.n921 B.n17 10.6151
R1556 B.n915 B.n17 10.6151
R1557 B.n915 B.n914 10.6151
R1558 B.n914 B.n913 10.6151
R1559 B.n913 B.n23 10.6151
R1560 B.n907 B.n23 10.6151
R1561 B.n907 B.n906 10.6151
R1562 B.n906 B.n905 10.6151
R1563 B.n905 B.n31 10.6151
R1564 B.n899 B.n31 10.6151
R1565 B.n899 B.n898 10.6151
R1566 B.n898 B.n897 10.6151
R1567 B.n897 B.n38 10.6151
R1568 B.n891 B.n38 10.6151
R1569 B.n891 B.n890 10.6151
R1570 B.n890 B.n889 10.6151
R1571 B.n889 B.n45 10.6151
R1572 B.n883 B.n45 10.6151
R1573 B.n883 B.n882 10.6151
R1574 B.n882 B.n881 10.6151
R1575 B.n881 B.n51 10.6151
R1576 B.n875 B.n51 10.6151
R1577 B.n875 B.n874 10.6151
R1578 B.n874 B.n873 10.6151
R1579 B.n873 B.n59 10.6151
R1580 B.n867 B.n59 10.6151
R1581 B.n867 B.n866 10.6151
R1582 B.n866 B.n865 10.6151
R1583 B.n865 B.n66 10.6151
R1584 B.n859 B.n66 10.6151
R1585 B.n859 B.n858 10.6151
R1586 B.n858 B.n857 10.6151
R1587 B.n857 B.n73 10.6151
R1588 B.n851 B.n73 10.6151
R1589 B.n762 B.n761 9.36635
R1590 B.n738 B.n112 9.36635
R1591 B.n381 B.n240 9.36635
R1592 B.n357 B.n248 9.36635
R1593 B.n512 B.t0 4.74571
R1594 B.n53 B.t6 4.74571
R1595 B.n937 B.n0 2.81026
R1596 B.n937 B.n1 2.81026
R1597 B.n761 B.n760 1.24928
R1598 B.n112 B.n108 1.24928
R1599 B.n377 B.n240 1.24928
R1600 B.n361 B.n248 1.24928
R1601 B.n568 B.t8 1.1868
R1602 B.n917 B.t2 1.1868
R1603 VP.n14 VP.t5 232.237
R1604 VP.n39 VP.t6 202.411
R1605 VP.n46 VP.t3 202.411
R1606 VP.n53 VP.t2 202.411
R1607 VP.n60 VP.t8 202.411
R1608 VP.n67 VP.t1 202.411
R1609 VP.n36 VP.t9 202.411
R1610 VP.n29 VP.t4 202.411
R1611 VP.n22 VP.t7 202.411
R1612 VP.n15 VP.t0 202.411
R1613 VP.n39 VP.n38 182.343
R1614 VP.n68 VP.n67 182.343
R1615 VP.n37 VP.n36 182.343
R1616 VP.n17 VP.n16 161.3
R1617 VP.n18 VP.n13 161.3
R1618 VP.n20 VP.n19 161.3
R1619 VP.n21 VP.n12 161.3
R1620 VP.n24 VP.n23 161.3
R1621 VP.n25 VP.n11 161.3
R1622 VP.n27 VP.n26 161.3
R1623 VP.n28 VP.n10 161.3
R1624 VP.n31 VP.n30 161.3
R1625 VP.n32 VP.n9 161.3
R1626 VP.n34 VP.n33 161.3
R1627 VP.n35 VP.n8 161.3
R1628 VP.n66 VP.n0 161.3
R1629 VP.n65 VP.n64 161.3
R1630 VP.n63 VP.n1 161.3
R1631 VP.n62 VP.n61 161.3
R1632 VP.n59 VP.n2 161.3
R1633 VP.n58 VP.n57 161.3
R1634 VP.n56 VP.n3 161.3
R1635 VP.n55 VP.n54 161.3
R1636 VP.n52 VP.n4 161.3
R1637 VP.n51 VP.n50 161.3
R1638 VP.n49 VP.n5 161.3
R1639 VP.n48 VP.n47 161.3
R1640 VP.n45 VP.n6 161.3
R1641 VP.n44 VP.n43 161.3
R1642 VP.n42 VP.n7 161.3
R1643 VP.n41 VP.n40 161.3
R1644 VP.n15 VP.n14 59.0939
R1645 VP.n51 VP.n5 56.5193
R1646 VP.n58 VP.n3 56.5193
R1647 VP.n27 VP.n11 56.5193
R1648 VP.n20 VP.n13 56.5193
R1649 VP.n44 VP.n7 51.663
R1650 VP.n65 VP.n1 51.663
R1651 VP.n34 VP.n9 51.663
R1652 VP.n38 VP.n37 48.3755
R1653 VP.n45 VP.n44 29.3238
R1654 VP.n61 VP.n1 29.3238
R1655 VP.n30 VP.n9 29.3238
R1656 VP.n40 VP.n7 24.4675
R1657 VP.n47 VP.n5 24.4675
R1658 VP.n52 VP.n51 24.4675
R1659 VP.n54 VP.n3 24.4675
R1660 VP.n59 VP.n58 24.4675
R1661 VP.n66 VP.n65 24.4675
R1662 VP.n35 VP.n34 24.4675
R1663 VP.n28 VP.n27 24.4675
R1664 VP.n21 VP.n20 24.4675
R1665 VP.n23 VP.n11 24.4675
R1666 VP.n16 VP.n13 24.4675
R1667 VP.n17 VP.n14 18.5156
R1668 VP.n46 VP.n45 16.6381
R1669 VP.n61 VP.n60 16.6381
R1670 VP.n30 VP.n29 16.6381
R1671 VP.n53 VP.n52 12.234
R1672 VP.n54 VP.n53 12.234
R1673 VP.n22 VP.n21 12.234
R1674 VP.n23 VP.n22 12.234
R1675 VP.n47 VP.n46 7.82994
R1676 VP.n60 VP.n59 7.82994
R1677 VP.n29 VP.n28 7.82994
R1678 VP.n16 VP.n15 7.82994
R1679 VP.n40 VP.n39 3.42588
R1680 VP.n67 VP.n66 3.42588
R1681 VP.n36 VP.n35 3.42588
R1682 VP.n18 VP.n17 0.189894
R1683 VP.n19 VP.n18 0.189894
R1684 VP.n19 VP.n12 0.189894
R1685 VP.n24 VP.n12 0.189894
R1686 VP.n25 VP.n24 0.189894
R1687 VP.n26 VP.n25 0.189894
R1688 VP.n26 VP.n10 0.189894
R1689 VP.n31 VP.n10 0.189894
R1690 VP.n32 VP.n31 0.189894
R1691 VP.n33 VP.n32 0.189894
R1692 VP.n33 VP.n8 0.189894
R1693 VP.n37 VP.n8 0.189894
R1694 VP.n41 VP.n38 0.189894
R1695 VP.n42 VP.n41 0.189894
R1696 VP.n43 VP.n42 0.189894
R1697 VP.n43 VP.n6 0.189894
R1698 VP.n48 VP.n6 0.189894
R1699 VP.n49 VP.n48 0.189894
R1700 VP.n50 VP.n49 0.189894
R1701 VP.n50 VP.n4 0.189894
R1702 VP.n55 VP.n4 0.189894
R1703 VP.n56 VP.n55 0.189894
R1704 VP.n57 VP.n56 0.189894
R1705 VP.n57 VP.n2 0.189894
R1706 VP.n62 VP.n2 0.189894
R1707 VP.n63 VP.n62 0.189894
R1708 VP.n64 VP.n63 0.189894
R1709 VP.n64 VP.n0 0.189894
R1710 VP.n68 VP.n0 0.189894
R1711 VP VP.n68 0.0516364
R1712 VDD1.n66 VDD1.n0 214.453
R1713 VDD1.n139 VDD1.n73 214.453
R1714 VDD1.n67 VDD1.n66 185
R1715 VDD1.n65 VDD1.n64 185
R1716 VDD1.n4 VDD1.n3 185
R1717 VDD1.n59 VDD1.n58 185
R1718 VDD1.n57 VDD1.n56 185
R1719 VDD1.n8 VDD1.n7 185
R1720 VDD1.n51 VDD1.n50 185
R1721 VDD1.n49 VDD1.n48 185
R1722 VDD1.n12 VDD1.n11 185
R1723 VDD1.n43 VDD1.n42 185
R1724 VDD1.n41 VDD1.n40 185
R1725 VDD1.n16 VDD1.n15 185
R1726 VDD1.n35 VDD1.n34 185
R1727 VDD1.n33 VDD1.n32 185
R1728 VDD1.n20 VDD1.n19 185
R1729 VDD1.n27 VDD1.n26 185
R1730 VDD1.n25 VDD1.n24 185
R1731 VDD1.n98 VDD1.n97 185
R1732 VDD1.n100 VDD1.n99 185
R1733 VDD1.n93 VDD1.n92 185
R1734 VDD1.n106 VDD1.n105 185
R1735 VDD1.n108 VDD1.n107 185
R1736 VDD1.n89 VDD1.n88 185
R1737 VDD1.n114 VDD1.n113 185
R1738 VDD1.n116 VDD1.n115 185
R1739 VDD1.n85 VDD1.n84 185
R1740 VDD1.n122 VDD1.n121 185
R1741 VDD1.n124 VDD1.n123 185
R1742 VDD1.n81 VDD1.n80 185
R1743 VDD1.n130 VDD1.n129 185
R1744 VDD1.n132 VDD1.n131 185
R1745 VDD1.n77 VDD1.n76 185
R1746 VDD1.n138 VDD1.n137 185
R1747 VDD1.n140 VDD1.n139 185
R1748 VDD1.n96 VDD1.t0 147.659
R1749 VDD1.n23 VDD1.t8 147.659
R1750 VDD1.n66 VDD1.n65 104.615
R1751 VDD1.n65 VDD1.n3 104.615
R1752 VDD1.n58 VDD1.n3 104.615
R1753 VDD1.n58 VDD1.n57 104.615
R1754 VDD1.n57 VDD1.n7 104.615
R1755 VDD1.n50 VDD1.n7 104.615
R1756 VDD1.n50 VDD1.n49 104.615
R1757 VDD1.n49 VDD1.n11 104.615
R1758 VDD1.n42 VDD1.n11 104.615
R1759 VDD1.n42 VDD1.n41 104.615
R1760 VDD1.n41 VDD1.n15 104.615
R1761 VDD1.n34 VDD1.n15 104.615
R1762 VDD1.n34 VDD1.n33 104.615
R1763 VDD1.n33 VDD1.n19 104.615
R1764 VDD1.n26 VDD1.n19 104.615
R1765 VDD1.n26 VDD1.n25 104.615
R1766 VDD1.n99 VDD1.n98 104.615
R1767 VDD1.n99 VDD1.n92 104.615
R1768 VDD1.n106 VDD1.n92 104.615
R1769 VDD1.n107 VDD1.n106 104.615
R1770 VDD1.n107 VDD1.n88 104.615
R1771 VDD1.n114 VDD1.n88 104.615
R1772 VDD1.n115 VDD1.n114 104.615
R1773 VDD1.n115 VDD1.n84 104.615
R1774 VDD1.n122 VDD1.n84 104.615
R1775 VDD1.n123 VDD1.n122 104.615
R1776 VDD1.n123 VDD1.n80 104.615
R1777 VDD1.n130 VDD1.n80 104.615
R1778 VDD1.n131 VDD1.n130 104.615
R1779 VDD1.n131 VDD1.n76 104.615
R1780 VDD1.n138 VDD1.n76 104.615
R1781 VDD1.n139 VDD1.n138 104.615
R1782 VDD1.n147 VDD1.n146 63.6566
R1783 VDD1.n72 VDD1.n71 62.4772
R1784 VDD1.n149 VDD1.n148 62.477
R1785 VDD1.n145 VDD1.n144 62.477
R1786 VDD1.n25 VDD1.t8 52.3082
R1787 VDD1.n98 VDD1.t0 52.3082
R1788 VDD1.n72 VDD1.n70 51.8683
R1789 VDD1.n145 VDD1.n143 51.8683
R1790 VDD1.n149 VDD1.n147 44.3824
R1791 VDD1.n24 VDD1.n23 15.6677
R1792 VDD1.n97 VDD1.n96 15.6677
R1793 VDD1.n68 VDD1.n67 12.8005
R1794 VDD1.n27 VDD1.n22 12.8005
R1795 VDD1.n100 VDD1.n95 12.8005
R1796 VDD1.n141 VDD1.n140 12.8005
R1797 VDD1.n64 VDD1.n2 12.0247
R1798 VDD1.n28 VDD1.n20 12.0247
R1799 VDD1.n101 VDD1.n93 12.0247
R1800 VDD1.n137 VDD1.n75 12.0247
R1801 VDD1.n63 VDD1.n4 11.249
R1802 VDD1.n32 VDD1.n31 11.249
R1803 VDD1.n105 VDD1.n104 11.249
R1804 VDD1.n136 VDD1.n77 11.249
R1805 VDD1.n60 VDD1.n59 10.4732
R1806 VDD1.n35 VDD1.n18 10.4732
R1807 VDD1.n108 VDD1.n91 10.4732
R1808 VDD1.n133 VDD1.n132 10.4732
R1809 VDD1.n56 VDD1.n6 9.69747
R1810 VDD1.n36 VDD1.n16 9.69747
R1811 VDD1.n109 VDD1.n89 9.69747
R1812 VDD1.n129 VDD1.n79 9.69747
R1813 VDD1.n70 VDD1.n69 9.45567
R1814 VDD1.n143 VDD1.n142 9.45567
R1815 VDD1.n10 VDD1.n9 9.3005
R1816 VDD1.n53 VDD1.n52 9.3005
R1817 VDD1.n55 VDD1.n54 9.3005
R1818 VDD1.n6 VDD1.n5 9.3005
R1819 VDD1.n61 VDD1.n60 9.3005
R1820 VDD1.n63 VDD1.n62 9.3005
R1821 VDD1.n2 VDD1.n1 9.3005
R1822 VDD1.n69 VDD1.n68 9.3005
R1823 VDD1.n47 VDD1.n46 9.3005
R1824 VDD1.n45 VDD1.n44 9.3005
R1825 VDD1.n14 VDD1.n13 9.3005
R1826 VDD1.n39 VDD1.n38 9.3005
R1827 VDD1.n37 VDD1.n36 9.3005
R1828 VDD1.n18 VDD1.n17 9.3005
R1829 VDD1.n31 VDD1.n30 9.3005
R1830 VDD1.n29 VDD1.n28 9.3005
R1831 VDD1.n22 VDD1.n21 9.3005
R1832 VDD1.n118 VDD1.n117 9.3005
R1833 VDD1.n87 VDD1.n86 9.3005
R1834 VDD1.n112 VDD1.n111 9.3005
R1835 VDD1.n110 VDD1.n109 9.3005
R1836 VDD1.n91 VDD1.n90 9.3005
R1837 VDD1.n104 VDD1.n103 9.3005
R1838 VDD1.n102 VDD1.n101 9.3005
R1839 VDD1.n95 VDD1.n94 9.3005
R1840 VDD1.n120 VDD1.n119 9.3005
R1841 VDD1.n83 VDD1.n82 9.3005
R1842 VDD1.n126 VDD1.n125 9.3005
R1843 VDD1.n128 VDD1.n127 9.3005
R1844 VDD1.n79 VDD1.n78 9.3005
R1845 VDD1.n134 VDD1.n133 9.3005
R1846 VDD1.n136 VDD1.n135 9.3005
R1847 VDD1.n75 VDD1.n74 9.3005
R1848 VDD1.n142 VDD1.n141 9.3005
R1849 VDD1.n55 VDD1.n8 8.92171
R1850 VDD1.n40 VDD1.n39 8.92171
R1851 VDD1.n113 VDD1.n112 8.92171
R1852 VDD1.n128 VDD1.n81 8.92171
R1853 VDD1.n70 VDD1.n0 8.2187
R1854 VDD1.n143 VDD1.n73 8.2187
R1855 VDD1.n52 VDD1.n51 8.14595
R1856 VDD1.n43 VDD1.n14 8.14595
R1857 VDD1.n116 VDD1.n87 8.14595
R1858 VDD1.n125 VDD1.n124 8.14595
R1859 VDD1.n48 VDD1.n10 7.3702
R1860 VDD1.n44 VDD1.n12 7.3702
R1861 VDD1.n117 VDD1.n85 7.3702
R1862 VDD1.n121 VDD1.n83 7.3702
R1863 VDD1.n48 VDD1.n47 6.59444
R1864 VDD1.n47 VDD1.n12 6.59444
R1865 VDD1.n120 VDD1.n85 6.59444
R1866 VDD1.n121 VDD1.n120 6.59444
R1867 VDD1.n51 VDD1.n10 5.81868
R1868 VDD1.n44 VDD1.n43 5.81868
R1869 VDD1.n117 VDD1.n116 5.81868
R1870 VDD1.n124 VDD1.n83 5.81868
R1871 VDD1.n68 VDD1.n0 5.3904
R1872 VDD1.n141 VDD1.n73 5.3904
R1873 VDD1.n52 VDD1.n8 5.04292
R1874 VDD1.n40 VDD1.n14 5.04292
R1875 VDD1.n113 VDD1.n87 5.04292
R1876 VDD1.n125 VDD1.n81 5.04292
R1877 VDD1.n96 VDD1.n94 4.38563
R1878 VDD1.n23 VDD1.n21 4.38563
R1879 VDD1.n56 VDD1.n55 4.26717
R1880 VDD1.n39 VDD1.n16 4.26717
R1881 VDD1.n112 VDD1.n89 4.26717
R1882 VDD1.n129 VDD1.n128 4.26717
R1883 VDD1.n59 VDD1.n6 3.49141
R1884 VDD1.n36 VDD1.n35 3.49141
R1885 VDD1.n109 VDD1.n108 3.49141
R1886 VDD1.n132 VDD1.n79 3.49141
R1887 VDD1.n60 VDD1.n4 2.71565
R1888 VDD1.n32 VDD1.n18 2.71565
R1889 VDD1.n105 VDD1.n91 2.71565
R1890 VDD1.n133 VDD1.n77 2.71565
R1891 VDD1.n64 VDD1.n63 1.93989
R1892 VDD1.n31 VDD1.n20 1.93989
R1893 VDD1.n104 VDD1.n93 1.93989
R1894 VDD1.n137 VDD1.n136 1.93989
R1895 VDD1.n148 VDD1.t6 1.49259
R1896 VDD1.n148 VDD1.t9 1.49259
R1897 VDD1.n71 VDD1.t2 1.49259
R1898 VDD1.n71 VDD1.t7 1.49259
R1899 VDD1.n146 VDD1.t3 1.49259
R1900 VDD1.n146 VDD1.t4 1.49259
R1901 VDD1.n144 VDD1.t5 1.49259
R1902 VDD1.n144 VDD1.t1 1.49259
R1903 VDD1 VDD1.n149 1.17722
R1904 VDD1.n67 VDD1.n2 1.16414
R1905 VDD1.n28 VDD1.n27 1.16414
R1906 VDD1.n101 VDD1.n100 1.16414
R1907 VDD1.n140 VDD1.n75 1.16414
R1908 VDD1 VDD1.n72 0.470328
R1909 VDD1.n24 VDD1.n22 0.388379
R1910 VDD1.n97 VDD1.n95 0.388379
R1911 VDD1.n147 VDD1.n145 0.356792
R1912 VDD1.n69 VDD1.n1 0.155672
R1913 VDD1.n62 VDD1.n1 0.155672
R1914 VDD1.n62 VDD1.n61 0.155672
R1915 VDD1.n61 VDD1.n5 0.155672
R1916 VDD1.n54 VDD1.n5 0.155672
R1917 VDD1.n54 VDD1.n53 0.155672
R1918 VDD1.n53 VDD1.n9 0.155672
R1919 VDD1.n46 VDD1.n9 0.155672
R1920 VDD1.n46 VDD1.n45 0.155672
R1921 VDD1.n45 VDD1.n13 0.155672
R1922 VDD1.n38 VDD1.n13 0.155672
R1923 VDD1.n38 VDD1.n37 0.155672
R1924 VDD1.n37 VDD1.n17 0.155672
R1925 VDD1.n30 VDD1.n17 0.155672
R1926 VDD1.n30 VDD1.n29 0.155672
R1927 VDD1.n29 VDD1.n21 0.155672
R1928 VDD1.n102 VDD1.n94 0.155672
R1929 VDD1.n103 VDD1.n102 0.155672
R1930 VDD1.n103 VDD1.n90 0.155672
R1931 VDD1.n110 VDD1.n90 0.155672
R1932 VDD1.n111 VDD1.n110 0.155672
R1933 VDD1.n111 VDD1.n86 0.155672
R1934 VDD1.n118 VDD1.n86 0.155672
R1935 VDD1.n119 VDD1.n118 0.155672
R1936 VDD1.n119 VDD1.n82 0.155672
R1937 VDD1.n126 VDD1.n82 0.155672
R1938 VDD1.n127 VDD1.n126 0.155672
R1939 VDD1.n127 VDD1.n78 0.155672
R1940 VDD1.n134 VDD1.n78 0.155672
R1941 VDD1.n135 VDD1.n134 0.155672
R1942 VDD1.n135 VDD1.n74 0.155672
R1943 VDD1.n142 VDD1.n74 0.155672
R1944 VTAIL.n296 VTAIL.n230 214.453
R1945 VTAIL.n68 VTAIL.n2 214.453
R1946 VTAIL.n224 VTAIL.n158 214.453
R1947 VTAIL.n148 VTAIL.n82 214.453
R1948 VTAIL.n255 VTAIL.n254 185
R1949 VTAIL.n257 VTAIL.n256 185
R1950 VTAIL.n250 VTAIL.n249 185
R1951 VTAIL.n263 VTAIL.n262 185
R1952 VTAIL.n265 VTAIL.n264 185
R1953 VTAIL.n246 VTAIL.n245 185
R1954 VTAIL.n271 VTAIL.n270 185
R1955 VTAIL.n273 VTAIL.n272 185
R1956 VTAIL.n242 VTAIL.n241 185
R1957 VTAIL.n279 VTAIL.n278 185
R1958 VTAIL.n281 VTAIL.n280 185
R1959 VTAIL.n238 VTAIL.n237 185
R1960 VTAIL.n287 VTAIL.n286 185
R1961 VTAIL.n289 VTAIL.n288 185
R1962 VTAIL.n234 VTAIL.n233 185
R1963 VTAIL.n295 VTAIL.n294 185
R1964 VTAIL.n297 VTAIL.n296 185
R1965 VTAIL.n27 VTAIL.n26 185
R1966 VTAIL.n29 VTAIL.n28 185
R1967 VTAIL.n22 VTAIL.n21 185
R1968 VTAIL.n35 VTAIL.n34 185
R1969 VTAIL.n37 VTAIL.n36 185
R1970 VTAIL.n18 VTAIL.n17 185
R1971 VTAIL.n43 VTAIL.n42 185
R1972 VTAIL.n45 VTAIL.n44 185
R1973 VTAIL.n14 VTAIL.n13 185
R1974 VTAIL.n51 VTAIL.n50 185
R1975 VTAIL.n53 VTAIL.n52 185
R1976 VTAIL.n10 VTAIL.n9 185
R1977 VTAIL.n59 VTAIL.n58 185
R1978 VTAIL.n61 VTAIL.n60 185
R1979 VTAIL.n6 VTAIL.n5 185
R1980 VTAIL.n67 VTAIL.n66 185
R1981 VTAIL.n69 VTAIL.n68 185
R1982 VTAIL.n225 VTAIL.n224 185
R1983 VTAIL.n223 VTAIL.n222 185
R1984 VTAIL.n162 VTAIL.n161 185
R1985 VTAIL.n217 VTAIL.n216 185
R1986 VTAIL.n215 VTAIL.n214 185
R1987 VTAIL.n166 VTAIL.n165 185
R1988 VTAIL.n209 VTAIL.n208 185
R1989 VTAIL.n207 VTAIL.n206 185
R1990 VTAIL.n170 VTAIL.n169 185
R1991 VTAIL.n201 VTAIL.n200 185
R1992 VTAIL.n199 VTAIL.n198 185
R1993 VTAIL.n174 VTAIL.n173 185
R1994 VTAIL.n193 VTAIL.n192 185
R1995 VTAIL.n191 VTAIL.n190 185
R1996 VTAIL.n178 VTAIL.n177 185
R1997 VTAIL.n185 VTAIL.n184 185
R1998 VTAIL.n183 VTAIL.n182 185
R1999 VTAIL.n149 VTAIL.n148 185
R2000 VTAIL.n147 VTAIL.n146 185
R2001 VTAIL.n86 VTAIL.n85 185
R2002 VTAIL.n141 VTAIL.n140 185
R2003 VTAIL.n139 VTAIL.n138 185
R2004 VTAIL.n90 VTAIL.n89 185
R2005 VTAIL.n133 VTAIL.n132 185
R2006 VTAIL.n131 VTAIL.n130 185
R2007 VTAIL.n94 VTAIL.n93 185
R2008 VTAIL.n125 VTAIL.n124 185
R2009 VTAIL.n123 VTAIL.n122 185
R2010 VTAIL.n98 VTAIL.n97 185
R2011 VTAIL.n117 VTAIL.n116 185
R2012 VTAIL.n115 VTAIL.n114 185
R2013 VTAIL.n102 VTAIL.n101 185
R2014 VTAIL.n109 VTAIL.n108 185
R2015 VTAIL.n107 VTAIL.n106 185
R2016 VTAIL.n253 VTAIL.t4 147.659
R2017 VTAIL.n25 VTAIL.t18 147.659
R2018 VTAIL.n181 VTAIL.t10 147.659
R2019 VTAIL.n105 VTAIL.t2 147.659
R2020 VTAIL.n256 VTAIL.n255 104.615
R2021 VTAIL.n256 VTAIL.n249 104.615
R2022 VTAIL.n263 VTAIL.n249 104.615
R2023 VTAIL.n264 VTAIL.n263 104.615
R2024 VTAIL.n264 VTAIL.n245 104.615
R2025 VTAIL.n271 VTAIL.n245 104.615
R2026 VTAIL.n272 VTAIL.n271 104.615
R2027 VTAIL.n272 VTAIL.n241 104.615
R2028 VTAIL.n279 VTAIL.n241 104.615
R2029 VTAIL.n280 VTAIL.n279 104.615
R2030 VTAIL.n280 VTAIL.n237 104.615
R2031 VTAIL.n287 VTAIL.n237 104.615
R2032 VTAIL.n288 VTAIL.n287 104.615
R2033 VTAIL.n288 VTAIL.n233 104.615
R2034 VTAIL.n295 VTAIL.n233 104.615
R2035 VTAIL.n296 VTAIL.n295 104.615
R2036 VTAIL.n28 VTAIL.n27 104.615
R2037 VTAIL.n28 VTAIL.n21 104.615
R2038 VTAIL.n35 VTAIL.n21 104.615
R2039 VTAIL.n36 VTAIL.n35 104.615
R2040 VTAIL.n36 VTAIL.n17 104.615
R2041 VTAIL.n43 VTAIL.n17 104.615
R2042 VTAIL.n44 VTAIL.n43 104.615
R2043 VTAIL.n44 VTAIL.n13 104.615
R2044 VTAIL.n51 VTAIL.n13 104.615
R2045 VTAIL.n52 VTAIL.n51 104.615
R2046 VTAIL.n52 VTAIL.n9 104.615
R2047 VTAIL.n59 VTAIL.n9 104.615
R2048 VTAIL.n60 VTAIL.n59 104.615
R2049 VTAIL.n60 VTAIL.n5 104.615
R2050 VTAIL.n67 VTAIL.n5 104.615
R2051 VTAIL.n68 VTAIL.n67 104.615
R2052 VTAIL.n224 VTAIL.n223 104.615
R2053 VTAIL.n223 VTAIL.n161 104.615
R2054 VTAIL.n216 VTAIL.n161 104.615
R2055 VTAIL.n216 VTAIL.n215 104.615
R2056 VTAIL.n215 VTAIL.n165 104.615
R2057 VTAIL.n208 VTAIL.n165 104.615
R2058 VTAIL.n208 VTAIL.n207 104.615
R2059 VTAIL.n207 VTAIL.n169 104.615
R2060 VTAIL.n200 VTAIL.n169 104.615
R2061 VTAIL.n200 VTAIL.n199 104.615
R2062 VTAIL.n199 VTAIL.n173 104.615
R2063 VTAIL.n192 VTAIL.n173 104.615
R2064 VTAIL.n192 VTAIL.n191 104.615
R2065 VTAIL.n191 VTAIL.n177 104.615
R2066 VTAIL.n184 VTAIL.n177 104.615
R2067 VTAIL.n184 VTAIL.n183 104.615
R2068 VTAIL.n148 VTAIL.n147 104.615
R2069 VTAIL.n147 VTAIL.n85 104.615
R2070 VTAIL.n140 VTAIL.n85 104.615
R2071 VTAIL.n140 VTAIL.n139 104.615
R2072 VTAIL.n139 VTAIL.n89 104.615
R2073 VTAIL.n132 VTAIL.n89 104.615
R2074 VTAIL.n132 VTAIL.n131 104.615
R2075 VTAIL.n131 VTAIL.n93 104.615
R2076 VTAIL.n124 VTAIL.n93 104.615
R2077 VTAIL.n124 VTAIL.n123 104.615
R2078 VTAIL.n123 VTAIL.n97 104.615
R2079 VTAIL.n116 VTAIL.n97 104.615
R2080 VTAIL.n116 VTAIL.n115 104.615
R2081 VTAIL.n115 VTAIL.n101 104.615
R2082 VTAIL.n108 VTAIL.n101 104.615
R2083 VTAIL.n108 VTAIL.n107 104.615
R2084 VTAIL.n255 VTAIL.t4 52.3082
R2085 VTAIL.n27 VTAIL.t18 52.3082
R2086 VTAIL.n183 VTAIL.t10 52.3082
R2087 VTAIL.n107 VTAIL.t2 52.3082
R2088 VTAIL.n157 VTAIL.n156 45.7984
R2089 VTAIL.n155 VTAIL.n154 45.7984
R2090 VTAIL.n81 VTAIL.n80 45.7984
R2091 VTAIL.n79 VTAIL.n78 45.7984
R2092 VTAIL.n303 VTAIL.n302 45.7983
R2093 VTAIL.n1 VTAIL.n0 45.7983
R2094 VTAIL.n75 VTAIL.n74 45.7983
R2095 VTAIL.n77 VTAIL.n76 45.7983
R2096 VTAIL.n301 VTAIL.n300 33.5429
R2097 VTAIL.n73 VTAIL.n72 33.5429
R2098 VTAIL.n229 VTAIL.n228 33.5429
R2099 VTAIL.n153 VTAIL.n152 33.5429
R2100 VTAIL.n79 VTAIL.n77 27.0996
R2101 VTAIL.n301 VTAIL.n229 25.4531
R2102 VTAIL.n254 VTAIL.n253 15.6677
R2103 VTAIL.n26 VTAIL.n25 15.6677
R2104 VTAIL.n182 VTAIL.n181 15.6677
R2105 VTAIL.n106 VTAIL.n105 15.6677
R2106 VTAIL.n257 VTAIL.n252 12.8005
R2107 VTAIL.n298 VTAIL.n297 12.8005
R2108 VTAIL.n29 VTAIL.n24 12.8005
R2109 VTAIL.n70 VTAIL.n69 12.8005
R2110 VTAIL.n226 VTAIL.n225 12.8005
R2111 VTAIL.n185 VTAIL.n180 12.8005
R2112 VTAIL.n150 VTAIL.n149 12.8005
R2113 VTAIL.n109 VTAIL.n104 12.8005
R2114 VTAIL.n258 VTAIL.n250 12.0247
R2115 VTAIL.n294 VTAIL.n232 12.0247
R2116 VTAIL.n30 VTAIL.n22 12.0247
R2117 VTAIL.n66 VTAIL.n4 12.0247
R2118 VTAIL.n222 VTAIL.n160 12.0247
R2119 VTAIL.n186 VTAIL.n178 12.0247
R2120 VTAIL.n146 VTAIL.n84 12.0247
R2121 VTAIL.n110 VTAIL.n102 12.0247
R2122 VTAIL.n262 VTAIL.n261 11.249
R2123 VTAIL.n293 VTAIL.n234 11.249
R2124 VTAIL.n34 VTAIL.n33 11.249
R2125 VTAIL.n65 VTAIL.n6 11.249
R2126 VTAIL.n221 VTAIL.n162 11.249
R2127 VTAIL.n190 VTAIL.n189 11.249
R2128 VTAIL.n145 VTAIL.n86 11.249
R2129 VTAIL.n114 VTAIL.n113 11.249
R2130 VTAIL.n265 VTAIL.n248 10.4732
R2131 VTAIL.n290 VTAIL.n289 10.4732
R2132 VTAIL.n37 VTAIL.n20 10.4732
R2133 VTAIL.n62 VTAIL.n61 10.4732
R2134 VTAIL.n218 VTAIL.n217 10.4732
R2135 VTAIL.n193 VTAIL.n176 10.4732
R2136 VTAIL.n142 VTAIL.n141 10.4732
R2137 VTAIL.n117 VTAIL.n100 10.4732
R2138 VTAIL.n266 VTAIL.n246 9.69747
R2139 VTAIL.n286 VTAIL.n236 9.69747
R2140 VTAIL.n38 VTAIL.n18 9.69747
R2141 VTAIL.n58 VTAIL.n8 9.69747
R2142 VTAIL.n214 VTAIL.n164 9.69747
R2143 VTAIL.n194 VTAIL.n174 9.69747
R2144 VTAIL.n138 VTAIL.n88 9.69747
R2145 VTAIL.n118 VTAIL.n98 9.69747
R2146 VTAIL.n300 VTAIL.n299 9.45567
R2147 VTAIL.n72 VTAIL.n71 9.45567
R2148 VTAIL.n228 VTAIL.n227 9.45567
R2149 VTAIL.n152 VTAIL.n151 9.45567
R2150 VTAIL.n275 VTAIL.n274 9.3005
R2151 VTAIL.n244 VTAIL.n243 9.3005
R2152 VTAIL.n269 VTAIL.n268 9.3005
R2153 VTAIL.n267 VTAIL.n266 9.3005
R2154 VTAIL.n248 VTAIL.n247 9.3005
R2155 VTAIL.n261 VTAIL.n260 9.3005
R2156 VTAIL.n259 VTAIL.n258 9.3005
R2157 VTAIL.n252 VTAIL.n251 9.3005
R2158 VTAIL.n277 VTAIL.n276 9.3005
R2159 VTAIL.n240 VTAIL.n239 9.3005
R2160 VTAIL.n283 VTAIL.n282 9.3005
R2161 VTAIL.n285 VTAIL.n284 9.3005
R2162 VTAIL.n236 VTAIL.n235 9.3005
R2163 VTAIL.n291 VTAIL.n290 9.3005
R2164 VTAIL.n293 VTAIL.n292 9.3005
R2165 VTAIL.n232 VTAIL.n231 9.3005
R2166 VTAIL.n299 VTAIL.n298 9.3005
R2167 VTAIL.n47 VTAIL.n46 9.3005
R2168 VTAIL.n16 VTAIL.n15 9.3005
R2169 VTAIL.n41 VTAIL.n40 9.3005
R2170 VTAIL.n39 VTAIL.n38 9.3005
R2171 VTAIL.n20 VTAIL.n19 9.3005
R2172 VTAIL.n33 VTAIL.n32 9.3005
R2173 VTAIL.n31 VTAIL.n30 9.3005
R2174 VTAIL.n24 VTAIL.n23 9.3005
R2175 VTAIL.n49 VTAIL.n48 9.3005
R2176 VTAIL.n12 VTAIL.n11 9.3005
R2177 VTAIL.n55 VTAIL.n54 9.3005
R2178 VTAIL.n57 VTAIL.n56 9.3005
R2179 VTAIL.n8 VTAIL.n7 9.3005
R2180 VTAIL.n63 VTAIL.n62 9.3005
R2181 VTAIL.n65 VTAIL.n64 9.3005
R2182 VTAIL.n4 VTAIL.n3 9.3005
R2183 VTAIL.n71 VTAIL.n70 9.3005
R2184 VTAIL.n168 VTAIL.n167 9.3005
R2185 VTAIL.n211 VTAIL.n210 9.3005
R2186 VTAIL.n213 VTAIL.n212 9.3005
R2187 VTAIL.n164 VTAIL.n163 9.3005
R2188 VTAIL.n219 VTAIL.n218 9.3005
R2189 VTAIL.n221 VTAIL.n220 9.3005
R2190 VTAIL.n160 VTAIL.n159 9.3005
R2191 VTAIL.n227 VTAIL.n226 9.3005
R2192 VTAIL.n205 VTAIL.n204 9.3005
R2193 VTAIL.n203 VTAIL.n202 9.3005
R2194 VTAIL.n172 VTAIL.n171 9.3005
R2195 VTAIL.n197 VTAIL.n196 9.3005
R2196 VTAIL.n195 VTAIL.n194 9.3005
R2197 VTAIL.n176 VTAIL.n175 9.3005
R2198 VTAIL.n189 VTAIL.n188 9.3005
R2199 VTAIL.n187 VTAIL.n186 9.3005
R2200 VTAIL.n180 VTAIL.n179 9.3005
R2201 VTAIL.n92 VTAIL.n91 9.3005
R2202 VTAIL.n135 VTAIL.n134 9.3005
R2203 VTAIL.n137 VTAIL.n136 9.3005
R2204 VTAIL.n88 VTAIL.n87 9.3005
R2205 VTAIL.n143 VTAIL.n142 9.3005
R2206 VTAIL.n145 VTAIL.n144 9.3005
R2207 VTAIL.n84 VTAIL.n83 9.3005
R2208 VTAIL.n151 VTAIL.n150 9.3005
R2209 VTAIL.n129 VTAIL.n128 9.3005
R2210 VTAIL.n127 VTAIL.n126 9.3005
R2211 VTAIL.n96 VTAIL.n95 9.3005
R2212 VTAIL.n121 VTAIL.n120 9.3005
R2213 VTAIL.n119 VTAIL.n118 9.3005
R2214 VTAIL.n100 VTAIL.n99 9.3005
R2215 VTAIL.n113 VTAIL.n112 9.3005
R2216 VTAIL.n111 VTAIL.n110 9.3005
R2217 VTAIL.n104 VTAIL.n103 9.3005
R2218 VTAIL.n270 VTAIL.n269 8.92171
R2219 VTAIL.n285 VTAIL.n238 8.92171
R2220 VTAIL.n42 VTAIL.n41 8.92171
R2221 VTAIL.n57 VTAIL.n10 8.92171
R2222 VTAIL.n213 VTAIL.n166 8.92171
R2223 VTAIL.n198 VTAIL.n197 8.92171
R2224 VTAIL.n137 VTAIL.n90 8.92171
R2225 VTAIL.n122 VTAIL.n121 8.92171
R2226 VTAIL.n300 VTAIL.n230 8.2187
R2227 VTAIL.n72 VTAIL.n2 8.2187
R2228 VTAIL.n228 VTAIL.n158 8.2187
R2229 VTAIL.n152 VTAIL.n82 8.2187
R2230 VTAIL.n273 VTAIL.n244 8.14595
R2231 VTAIL.n282 VTAIL.n281 8.14595
R2232 VTAIL.n45 VTAIL.n16 8.14595
R2233 VTAIL.n54 VTAIL.n53 8.14595
R2234 VTAIL.n210 VTAIL.n209 8.14595
R2235 VTAIL.n201 VTAIL.n172 8.14595
R2236 VTAIL.n134 VTAIL.n133 8.14595
R2237 VTAIL.n125 VTAIL.n96 8.14595
R2238 VTAIL.n274 VTAIL.n242 7.3702
R2239 VTAIL.n278 VTAIL.n240 7.3702
R2240 VTAIL.n46 VTAIL.n14 7.3702
R2241 VTAIL.n50 VTAIL.n12 7.3702
R2242 VTAIL.n206 VTAIL.n168 7.3702
R2243 VTAIL.n202 VTAIL.n170 7.3702
R2244 VTAIL.n130 VTAIL.n92 7.3702
R2245 VTAIL.n126 VTAIL.n94 7.3702
R2246 VTAIL.n277 VTAIL.n242 6.59444
R2247 VTAIL.n278 VTAIL.n277 6.59444
R2248 VTAIL.n49 VTAIL.n14 6.59444
R2249 VTAIL.n50 VTAIL.n49 6.59444
R2250 VTAIL.n206 VTAIL.n205 6.59444
R2251 VTAIL.n205 VTAIL.n170 6.59444
R2252 VTAIL.n130 VTAIL.n129 6.59444
R2253 VTAIL.n129 VTAIL.n94 6.59444
R2254 VTAIL.n274 VTAIL.n273 5.81868
R2255 VTAIL.n281 VTAIL.n240 5.81868
R2256 VTAIL.n46 VTAIL.n45 5.81868
R2257 VTAIL.n53 VTAIL.n12 5.81868
R2258 VTAIL.n209 VTAIL.n168 5.81868
R2259 VTAIL.n202 VTAIL.n201 5.81868
R2260 VTAIL.n133 VTAIL.n92 5.81868
R2261 VTAIL.n126 VTAIL.n125 5.81868
R2262 VTAIL.n298 VTAIL.n230 5.3904
R2263 VTAIL.n70 VTAIL.n2 5.3904
R2264 VTAIL.n226 VTAIL.n158 5.3904
R2265 VTAIL.n150 VTAIL.n82 5.3904
R2266 VTAIL.n270 VTAIL.n244 5.04292
R2267 VTAIL.n282 VTAIL.n238 5.04292
R2268 VTAIL.n42 VTAIL.n16 5.04292
R2269 VTAIL.n54 VTAIL.n10 5.04292
R2270 VTAIL.n210 VTAIL.n166 5.04292
R2271 VTAIL.n198 VTAIL.n172 5.04292
R2272 VTAIL.n134 VTAIL.n90 5.04292
R2273 VTAIL.n122 VTAIL.n96 5.04292
R2274 VTAIL.n253 VTAIL.n251 4.38563
R2275 VTAIL.n25 VTAIL.n23 4.38563
R2276 VTAIL.n181 VTAIL.n179 4.38563
R2277 VTAIL.n105 VTAIL.n103 4.38563
R2278 VTAIL.n269 VTAIL.n246 4.26717
R2279 VTAIL.n286 VTAIL.n285 4.26717
R2280 VTAIL.n41 VTAIL.n18 4.26717
R2281 VTAIL.n58 VTAIL.n57 4.26717
R2282 VTAIL.n214 VTAIL.n213 4.26717
R2283 VTAIL.n197 VTAIL.n174 4.26717
R2284 VTAIL.n138 VTAIL.n137 4.26717
R2285 VTAIL.n121 VTAIL.n98 4.26717
R2286 VTAIL.n266 VTAIL.n265 3.49141
R2287 VTAIL.n289 VTAIL.n236 3.49141
R2288 VTAIL.n38 VTAIL.n37 3.49141
R2289 VTAIL.n61 VTAIL.n8 3.49141
R2290 VTAIL.n217 VTAIL.n164 3.49141
R2291 VTAIL.n194 VTAIL.n193 3.49141
R2292 VTAIL.n141 VTAIL.n88 3.49141
R2293 VTAIL.n118 VTAIL.n117 3.49141
R2294 VTAIL.n262 VTAIL.n248 2.71565
R2295 VTAIL.n290 VTAIL.n234 2.71565
R2296 VTAIL.n34 VTAIL.n20 2.71565
R2297 VTAIL.n62 VTAIL.n6 2.71565
R2298 VTAIL.n218 VTAIL.n162 2.71565
R2299 VTAIL.n190 VTAIL.n176 2.71565
R2300 VTAIL.n142 VTAIL.n86 2.71565
R2301 VTAIL.n114 VTAIL.n100 2.71565
R2302 VTAIL.n261 VTAIL.n250 1.93989
R2303 VTAIL.n294 VTAIL.n293 1.93989
R2304 VTAIL.n33 VTAIL.n22 1.93989
R2305 VTAIL.n66 VTAIL.n65 1.93989
R2306 VTAIL.n222 VTAIL.n221 1.93989
R2307 VTAIL.n189 VTAIL.n178 1.93989
R2308 VTAIL.n146 VTAIL.n145 1.93989
R2309 VTAIL.n113 VTAIL.n102 1.93989
R2310 VTAIL.n81 VTAIL.n79 1.64705
R2311 VTAIL.n153 VTAIL.n81 1.64705
R2312 VTAIL.n157 VTAIL.n155 1.64705
R2313 VTAIL.n229 VTAIL.n157 1.64705
R2314 VTAIL.n77 VTAIL.n75 1.64705
R2315 VTAIL.n75 VTAIL.n73 1.64705
R2316 VTAIL.n303 VTAIL.n301 1.64705
R2317 VTAIL.n302 VTAIL.t1 1.49259
R2318 VTAIL.n302 VTAIL.t7 1.49259
R2319 VTAIL.n0 VTAIL.t8 1.49259
R2320 VTAIL.n0 VTAIL.t3 1.49259
R2321 VTAIL.n74 VTAIL.t17 1.49259
R2322 VTAIL.n74 VTAIL.t11 1.49259
R2323 VTAIL.n76 VTAIL.t13 1.49259
R2324 VTAIL.n76 VTAIL.t16 1.49259
R2325 VTAIL.n156 VTAIL.t12 1.49259
R2326 VTAIL.n156 VTAIL.t15 1.49259
R2327 VTAIL.n154 VTAIL.t14 1.49259
R2328 VTAIL.n154 VTAIL.t19 1.49259
R2329 VTAIL.n80 VTAIL.t5 1.49259
R2330 VTAIL.n80 VTAIL.t9 1.49259
R2331 VTAIL.n78 VTAIL.t0 1.49259
R2332 VTAIL.n78 VTAIL.t6 1.49259
R2333 VTAIL.n155 VTAIL.n153 1.2936
R2334 VTAIL.n73 VTAIL.n1 1.2936
R2335 VTAIL VTAIL.n1 1.2936
R2336 VTAIL.n258 VTAIL.n257 1.16414
R2337 VTAIL.n297 VTAIL.n232 1.16414
R2338 VTAIL.n30 VTAIL.n29 1.16414
R2339 VTAIL.n69 VTAIL.n4 1.16414
R2340 VTAIL.n225 VTAIL.n160 1.16414
R2341 VTAIL.n186 VTAIL.n185 1.16414
R2342 VTAIL.n149 VTAIL.n84 1.16414
R2343 VTAIL.n110 VTAIL.n109 1.16414
R2344 VTAIL.n254 VTAIL.n252 0.388379
R2345 VTAIL.n26 VTAIL.n24 0.388379
R2346 VTAIL.n182 VTAIL.n180 0.388379
R2347 VTAIL.n106 VTAIL.n104 0.388379
R2348 VTAIL VTAIL.n303 0.353948
R2349 VTAIL.n259 VTAIL.n251 0.155672
R2350 VTAIL.n260 VTAIL.n259 0.155672
R2351 VTAIL.n260 VTAIL.n247 0.155672
R2352 VTAIL.n267 VTAIL.n247 0.155672
R2353 VTAIL.n268 VTAIL.n267 0.155672
R2354 VTAIL.n268 VTAIL.n243 0.155672
R2355 VTAIL.n275 VTAIL.n243 0.155672
R2356 VTAIL.n276 VTAIL.n275 0.155672
R2357 VTAIL.n276 VTAIL.n239 0.155672
R2358 VTAIL.n283 VTAIL.n239 0.155672
R2359 VTAIL.n284 VTAIL.n283 0.155672
R2360 VTAIL.n284 VTAIL.n235 0.155672
R2361 VTAIL.n291 VTAIL.n235 0.155672
R2362 VTAIL.n292 VTAIL.n291 0.155672
R2363 VTAIL.n292 VTAIL.n231 0.155672
R2364 VTAIL.n299 VTAIL.n231 0.155672
R2365 VTAIL.n31 VTAIL.n23 0.155672
R2366 VTAIL.n32 VTAIL.n31 0.155672
R2367 VTAIL.n32 VTAIL.n19 0.155672
R2368 VTAIL.n39 VTAIL.n19 0.155672
R2369 VTAIL.n40 VTAIL.n39 0.155672
R2370 VTAIL.n40 VTAIL.n15 0.155672
R2371 VTAIL.n47 VTAIL.n15 0.155672
R2372 VTAIL.n48 VTAIL.n47 0.155672
R2373 VTAIL.n48 VTAIL.n11 0.155672
R2374 VTAIL.n55 VTAIL.n11 0.155672
R2375 VTAIL.n56 VTAIL.n55 0.155672
R2376 VTAIL.n56 VTAIL.n7 0.155672
R2377 VTAIL.n63 VTAIL.n7 0.155672
R2378 VTAIL.n64 VTAIL.n63 0.155672
R2379 VTAIL.n64 VTAIL.n3 0.155672
R2380 VTAIL.n71 VTAIL.n3 0.155672
R2381 VTAIL.n227 VTAIL.n159 0.155672
R2382 VTAIL.n220 VTAIL.n159 0.155672
R2383 VTAIL.n220 VTAIL.n219 0.155672
R2384 VTAIL.n219 VTAIL.n163 0.155672
R2385 VTAIL.n212 VTAIL.n163 0.155672
R2386 VTAIL.n212 VTAIL.n211 0.155672
R2387 VTAIL.n211 VTAIL.n167 0.155672
R2388 VTAIL.n204 VTAIL.n167 0.155672
R2389 VTAIL.n204 VTAIL.n203 0.155672
R2390 VTAIL.n203 VTAIL.n171 0.155672
R2391 VTAIL.n196 VTAIL.n171 0.155672
R2392 VTAIL.n196 VTAIL.n195 0.155672
R2393 VTAIL.n195 VTAIL.n175 0.155672
R2394 VTAIL.n188 VTAIL.n175 0.155672
R2395 VTAIL.n188 VTAIL.n187 0.155672
R2396 VTAIL.n187 VTAIL.n179 0.155672
R2397 VTAIL.n151 VTAIL.n83 0.155672
R2398 VTAIL.n144 VTAIL.n83 0.155672
R2399 VTAIL.n144 VTAIL.n143 0.155672
R2400 VTAIL.n143 VTAIL.n87 0.155672
R2401 VTAIL.n136 VTAIL.n87 0.155672
R2402 VTAIL.n136 VTAIL.n135 0.155672
R2403 VTAIL.n135 VTAIL.n91 0.155672
R2404 VTAIL.n128 VTAIL.n91 0.155672
R2405 VTAIL.n128 VTAIL.n127 0.155672
R2406 VTAIL.n127 VTAIL.n95 0.155672
R2407 VTAIL.n120 VTAIL.n95 0.155672
R2408 VTAIL.n120 VTAIL.n119 0.155672
R2409 VTAIL.n119 VTAIL.n99 0.155672
R2410 VTAIL.n112 VTAIL.n99 0.155672
R2411 VTAIL.n112 VTAIL.n111 0.155672
R2412 VTAIL.n111 VTAIL.n103 0.155672
R2413 VN.n6 VN.t1 232.237
R2414 VN.n36 VN.t5 232.237
R2415 VN.n7 VN.t7 202.411
R2416 VN.n14 VN.t8 202.411
R2417 VN.n21 VN.t3 202.411
R2418 VN.n28 VN.t6 202.411
R2419 VN.n37 VN.t2 202.411
R2420 VN.n44 VN.t9 202.411
R2421 VN.n51 VN.t4 202.411
R2422 VN.n58 VN.t0 202.411
R2423 VN.n29 VN.n28 182.343
R2424 VN.n59 VN.n58 182.343
R2425 VN.n57 VN.n30 161.3
R2426 VN.n56 VN.n55 161.3
R2427 VN.n54 VN.n31 161.3
R2428 VN.n53 VN.n52 161.3
R2429 VN.n50 VN.n32 161.3
R2430 VN.n49 VN.n48 161.3
R2431 VN.n47 VN.n33 161.3
R2432 VN.n46 VN.n45 161.3
R2433 VN.n43 VN.n34 161.3
R2434 VN.n42 VN.n41 161.3
R2435 VN.n40 VN.n35 161.3
R2436 VN.n39 VN.n38 161.3
R2437 VN.n27 VN.n0 161.3
R2438 VN.n26 VN.n25 161.3
R2439 VN.n24 VN.n1 161.3
R2440 VN.n23 VN.n22 161.3
R2441 VN.n20 VN.n2 161.3
R2442 VN.n19 VN.n18 161.3
R2443 VN.n17 VN.n3 161.3
R2444 VN.n16 VN.n15 161.3
R2445 VN.n13 VN.n4 161.3
R2446 VN.n12 VN.n11 161.3
R2447 VN.n10 VN.n5 161.3
R2448 VN.n9 VN.n8 161.3
R2449 VN.n7 VN.n6 59.0939
R2450 VN.n37 VN.n36 59.0939
R2451 VN.n12 VN.n5 56.5193
R2452 VN.n19 VN.n3 56.5193
R2453 VN.n42 VN.n35 56.5193
R2454 VN.n49 VN.n33 56.5193
R2455 VN.n26 VN.n1 51.663
R2456 VN.n56 VN.n31 51.663
R2457 VN VN.n59 48.7562
R2458 VN.n22 VN.n1 29.3238
R2459 VN.n52 VN.n31 29.3238
R2460 VN.n8 VN.n5 24.4675
R2461 VN.n13 VN.n12 24.4675
R2462 VN.n15 VN.n3 24.4675
R2463 VN.n20 VN.n19 24.4675
R2464 VN.n27 VN.n26 24.4675
R2465 VN.n38 VN.n35 24.4675
R2466 VN.n45 VN.n33 24.4675
R2467 VN.n43 VN.n42 24.4675
R2468 VN.n50 VN.n49 24.4675
R2469 VN.n57 VN.n56 24.4675
R2470 VN.n39 VN.n36 18.5156
R2471 VN.n9 VN.n6 18.5156
R2472 VN.n22 VN.n21 16.6381
R2473 VN.n52 VN.n51 16.6381
R2474 VN.n14 VN.n13 12.234
R2475 VN.n15 VN.n14 12.234
R2476 VN.n45 VN.n44 12.234
R2477 VN.n44 VN.n43 12.234
R2478 VN.n8 VN.n7 7.82994
R2479 VN.n21 VN.n20 7.82994
R2480 VN.n38 VN.n37 7.82994
R2481 VN.n51 VN.n50 7.82994
R2482 VN.n28 VN.n27 3.42588
R2483 VN.n58 VN.n57 3.42588
R2484 VN.n59 VN.n30 0.189894
R2485 VN.n55 VN.n30 0.189894
R2486 VN.n55 VN.n54 0.189894
R2487 VN.n54 VN.n53 0.189894
R2488 VN.n53 VN.n32 0.189894
R2489 VN.n48 VN.n32 0.189894
R2490 VN.n48 VN.n47 0.189894
R2491 VN.n47 VN.n46 0.189894
R2492 VN.n46 VN.n34 0.189894
R2493 VN.n41 VN.n34 0.189894
R2494 VN.n41 VN.n40 0.189894
R2495 VN.n40 VN.n39 0.189894
R2496 VN.n10 VN.n9 0.189894
R2497 VN.n11 VN.n10 0.189894
R2498 VN.n11 VN.n4 0.189894
R2499 VN.n16 VN.n4 0.189894
R2500 VN.n17 VN.n16 0.189894
R2501 VN.n18 VN.n17 0.189894
R2502 VN.n18 VN.n2 0.189894
R2503 VN.n23 VN.n2 0.189894
R2504 VN.n24 VN.n23 0.189894
R2505 VN.n25 VN.n24 0.189894
R2506 VN.n25 VN.n0 0.189894
R2507 VN.n29 VN.n0 0.189894
R2508 VN VN.n29 0.0516364
R2509 VDD2.n141 VDD2.n75 214.453
R2510 VDD2.n66 VDD2.n0 214.453
R2511 VDD2.n142 VDD2.n141 185
R2512 VDD2.n140 VDD2.n139 185
R2513 VDD2.n79 VDD2.n78 185
R2514 VDD2.n134 VDD2.n133 185
R2515 VDD2.n132 VDD2.n131 185
R2516 VDD2.n83 VDD2.n82 185
R2517 VDD2.n126 VDD2.n125 185
R2518 VDD2.n124 VDD2.n123 185
R2519 VDD2.n87 VDD2.n86 185
R2520 VDD2.n118 VDD2.n117 185
R2521 VDD2.n116 VDD2.n115 185
R2522 VDD2.n91 VDD2.n90 185
R2523 VDD2.n110 VDD2.n109 185
R2524 VDD2.n108 VDD2.n107 185
R2525 VDD2.n95 VDD2.n94 185
R2526 VDD2.n102 VDD2.n101 185
R2527 VDD2.n100 VDD2.n99 185
R2528 VDD2.n25 VDD2.n24 185
R2529 VDD2.n27 VDD2.n26 185
R2530 VDD2.n20 VDD2.n19 185
R2531 VDD2.n33 VDD2.n32 185
R2532 VDD2.n35 VDD2.n34 185
R2533 VDD2.n16 VDD2.n15 185
R2534 VDD2.n41 VDD2.n40 185
R2535 VDD2.n43 VDD2.n42 185
R2536 VDD2.n12 VDD2.n11 185
R2537 VDD2.n49 VDD2.n48 185
R2538 VDD2.n51 VDD2.n50 185
R2539 VDD2.n8 VDD2.n7 185
R2540 VDD2.n57 VDD2.n56 185
R2541 VDD2.n59 VDD2.n58 185
R2542 VDD2.n4 VDD2.n3 185
R2543 VDD2.n65 VDD2.n64 185
R2544 VDD2.n67 VDD2.n66 185
R2545 VDD2.n23 VDD2.t8 147.659
R2546 VDD2.n98 VDD2.t9 147.659
R2547 VDD2.n141 VDD2.n140 104.615
R2548 VDD2.n140 VDD2.n78 104.615
R2549 VDD2.n133 VDD2.n78 104.615
R2550 VDD2.n133 VDD2.n132 104.615
R2551 VDD2.n132 VDD2.n82 104.615
R2552 VDD2.n125 VDD2.n82 104.615
R2553 VDD2.n125 VDD2.n124 104.615
R2554 VDD2.n124 VDD2.n86 104.615
R2555 VDD2.n117 VDD2.n86 104.615
R2556 VDD2.n117 VDD2.n116 104.615
R2557 VDD2.n116 VDD2.n90 104.615
R2558 VDD2.n109 VDD2.n90 104.615
R2559 VDD2.n109 VDD2.n108 104.615
R2560 VDD2.n108 VDD2.n94 104.615
R2561 VDD2.n101 VDD2.n94 104.615
R2562 VDD2.n101 VDD2.n100 104.615
R2563 VDD2.n26 VDD2.n25 104.615
R2564 VDD2.n26 VDD2.n19 104.615
R2565 VDD2.n33 VDD2.n19 104.615
R2566 VDD2.n34 VDD2.n33 104.615
R2567 VDD2.n34 VDD2.n15 104.615
R2568 VDD2.n41 VDD2.n15 104.615
R2569 VDD2.n42 VDD2.n41 104.615
R2570 VDD2.n42 VDD2.n11 104.615
R2571 VDD2.n49 VDD2.n11 104.615
R2572 VDD2.n50 VDD2.n49 104.615
R2573 VDD2.n50 VDD2.n7 104.615
R2574 VDD2.n57 VDD2.n7 104.615
R2575 VDD2.n58 VDD2.n57 104.615
R2576 VDD2.n58 VDD2.n3 104.615
R2577 VDD2.n65 VDD2.n3 104.615
R2578 VDD2.n66 VDD2.n65 104.615
R2579 VDD2.n74 VDD2.n73 63.6566
R2580 VDD2 VDD2.n149 63.6538
R2581 VDD2.n148 VDD2.n147 62.4772
R2582 VDD2.n72 VDD2.n71 62.477
R2583 VDD2.n100 VDD2.t9 52.3082
R2584 VDD2.n25 VDD2.t8 52.3082
R2585 VDD2.n72 VDD2.n70 51.8683
R2586 VDD2.n146 VDD2.n145 50.2217
R2587 VDD2.n146 VDD2.n74 42.9761
R2588 VDD2.n99 VDD2.n98 15.6677
R2589 VDD2.n24 VDD2.n23 15.6677
R2590 VDD2.n143 VDD2.n142 12.8005
R2591 VDD2.n102 VDD2.n97 12.8005
R2592 VDD2.n27 VDD2.n22 12.8005
R2593 VDD2.n68 VDD2.n67 12.8005
R2594 VDD2.n139 VDD2.n77 12.0247
R2595 VDD2.n103 VDD2.n95 12.0247
R2596 VDD2.n28 VDD2.n20 12.0247
R2597 VDD2.n64 VDD2.n2 12.0247
R2598 VDD2.n138 VDD2.n79 11.249
R2599 VDD2.n107 VDD2.n106 11.249
R2600 VDD2.n32 VDD2.n31 11.249
R2601 VDD2.n63 VDD2.n4 11.249
R2602 VDD2.n135 VDD2.n134 10.4732
R2603 VDD2.n110 VDD2.n93 10.4732
R2604 VDD2.n35 VDD2.n18 10.4732
R2605 VDD2.n60 VDD2.n59 10.4732
R2606 VDD2.n131 VDD2.n81 9.69747
R2607 VDD2.n111 VDD2.n91 9.69747
R2608 VDD2.n36 VDD2.n16 9.69747
R2609 VDD2.n56 VDD2.n6 9.69747
R2610 VDD2.n145 VDD2.n144 9.45567
R2611 VDD2.n70 VDD2.n69 9.45567
R2612 VDD2.n85 VDD2.n84 9.3005
R2613 VDD2.n128 VDD2.n127 9.3005
R2614 VDD2.n130 VDD2.n129 9.3005
R2615 VDD2.n81 VDD2.n80 9.3005
R2616 VDD2.n136 VDD2.n135 9.3005
R2617 VDD2.n138 VDD2.n137 9.3005
R2618 VDD2.n77 VDD2.n76 9.3005
R2619 VDD2.n144 VDD2.n143 9.3005
R2620 VDD2.n122 VDD2.n121 9.3005
R2621 VDD2.n120 VDD2.n119 9.3005
R2622 VDD2.n89 VDD2.n88 9.3005
R2623 VDD2.n114 VDD2.n113 9.3005
R2624 VDD2.n112 VDD2.n111 9.3005
R2625 VDD2.n93 VDD2.n92 9.3005
R2626 VDD2.n106 VDD2.n105 9.3005
R2627 VDD2.n104 VDD2.n103 9.3005
R2628 VDD2.n97 VDD2.n96 9.3005
R2629 VDD2.n45 VDD2.n44 9.3005
R2630 VDD2.n14 VDD2.n13 9.3005
R2631 VDD2.n39 VDD2.n38 9.3005
R2632 VDD2.n37 VDD2.n36 9.3005
R2633 VDD2.n18 VDD2.n17 9.3005
R2634 VDD2.n31 VDD2.n30 9.3005
R2635 VDD2.n29 VDD2.n28 9.3005
R2636 VDD2.n22 VDD2.n21 9.3005
R2637 VDD2.n47 VDD2.n46 9.3005
R2638 VDD2.n10 VDD2.n9 9.3005
R2639 VDD2.n53 VDD2.n52 9.3005
R2640 VDD2.n55 VDD2.n54 9.3005
R2641 VDD2.n6 VDD2.n5 9.3005
R2642 VDD2.n61 VDD2.n60 9.3005
R2643 VDD2.n63 VDD2.n62 9.3005
R2644 VDD2.n2 VDD2.n1 9.3005
R2645 VDD2.n69 VDD2.n68 9.3005
R2646 VDD2.n130 VDD2.n83 8.92171
R2647 VDD2.n115 VDD2.n114 8.92171
R2648 VDD2.n40 VDD2.n39 8.92171
R2649 VDD2.n55 VDD2.n8 8.92171
R2650 VDD2.n145 VDD2.n75 8.2187
R2651 VDD2.n70 VDD2.n0 8.2187
R2652 VDD2.n127 VDD2.n126 8.14595
R2653 VDD2.n118 VDD2.n89 8.14595
R2654 VDD2.n43 VDD2.n14 8.14595
R2655 VDD2.n52 VDD2.n51 8.14595
R2656 VDD2.n123 VDD2.n85 7.3702
R2657 VDD2.n119 VDD2.n87 7.3702
R2658 VDD2.n44 VDD2.n12 7.3702
R2659 VDD2.n48 VDD2.n10 7.3702
R2660 VDD2.n123 VDD2.n122 6.59444
R2661 VDD2.n122 VDD2.n87 6.59444
R2662 VDD2.n47 VDD2.n12 6.59444
R2663 VDD2.n48 VDD2.n47 6.59444
R2664 VDD2.n126 VDD2.n85 5.81868
R2665 VDD2.n119 VDD2.n118 5.81868
R2666 VDD2.n44 VDD2.n43 5.81868
R2667 VDD2.n51 VDD2.n10 5.81868
R2668 VDD2.n143 VDD2.n75 5.3904
R2669 VDD2.n68 VDD2.n0 5.3904
R2670 VDD2.n127 VDD2.n83 5.04292
R2671 VDD2.n115 VDD2.n89 5.04292
R2672 VDD2.n40 VDD2.n14 5.04292
R2673 VDD2.n52 VDD2.n8 5.04292
R2674 VDD2.n23 VDD2.n21 4.38563
R2675 VDD2.n98 VDD2.n96 4.38563
R2676 VDD2.n131 VDD2.n130 4.26717
R2677 VDD2.n114 VDD2.n91 4.26717
R2678 VDD2.n39 VDD2.n16 4.26717
R2679 VDD2.n56 VDD2.n55 4.26717
R2680 VDD2.n134 VDD2.n81 3.49141
R2681 VDD2.n111 VDD2.n110 3.49141
R2682 VDD2.n36 VDD2.n35 3.49141
R2683 VDD2.n59 VDD2.n6 3.49141
R2684 VDD2.n135 VDD2.n79 2.71565
R2685 VDD2.n107 VDD2.n93 2.71565
R2686 VDD2.n32 VDD2.n18 2.71565
R2687 VDD2.n60 VDD2.n4 2.71565
R2688 VDD2.n139 VDD2.n138 1.93989
R2689 VDD2.n106 VDD2.n95 1.93989
R2690 VDD2.n31 VDD2.n20 1.93989
R2691 VDD2.n64 VDD2.n63 1.93989
R2692 VDD2.n148 VDD2.n146 1.64705
R2693 VDD2.n149 VDD2.t7 1.49259
R2694 VDD2.n149 VDD2.t4 1.49259
R2695 VDD2.n147 VDD2.t5 1.49259
R2696 VDD2.n147 VDD2.t0 1.49259
R2697 VDD2.n73 VDD2.t6 1.49259
R2698 VDD2.n73 VDD2.t3 1.49259
R2699 VDD2.n71 VDD2.t2 1.49259
R2700 VDD2.n71 VDD2.t1 1.49259
R2701 VDD2.n142 VDD2.n77 1.16414
R2702 VDD2.n103 VDD2.n102 1.16414
R2703 VDD2.n28 VDD2.n27 1.16414
R2704 VDD2.n67 VDD2.n2 1.16414
R2705 VDD2 VDD2.n148 0.470328
R2706 VDD2.n99 VDD2.n97 0.388379
R2707 VDD2.n24 VDD2.n22 0.388379
R2708 VDD2.n74 VDD2.n72 0.356792
R2709 VDD2.n144 VDD2.n76 0.155672
R2710 VDD2.n137 VDD2.n76 0.155672
R2711 VDD2.n137 VDD2.n136 0.155672
R2712 VDD2.n136 VDD2.n80 0.155672
R2713 VDD2.n129 VDD2.n80 0.155672
R2714 VDD2.n129 VDD2.n128 0.155672
R2715 VDD2.n128 VDD2.n84 0.155672
R2716 VDD2.n121 VDD2.n84 0.155672
R2717 VDD2.n121 VDD2.n120 0.155672
R2718 VDD2.n120 VDD2.n88 0.155672
R2719 VDD2.n113 VDD2.n88 0.155672
R2720 VDD2.n113 VDD2.n112 0.155672
R2721 VDD2.n112 VDD2.n92 0.155672
R2722 VDD2.n105 VDD2.n92 0.155672
R2723 VDD2.n105 VDD2.n104 0.155672
R2724 VDD2.n104 VDD2.n96 0.155672
R2725 VDD2.n29 VDD2.n21 0.155672
R2726 VDD2.n30 VDD2.n29 0.155672
R2727 VDD2.n30 VDD2.n17 0.155672
R2728 VDD2.n37 VDD2.n17 0.155672
R2729 VDD2.n38 VDD2.n37 0.155672
R2730 VDD2.n38 VDD2.n13 0.155672
R2731 VDD2.n45 VDD2.n13 0.155672
R2732 VDD2.n46 VDD2.n45 0.155672
R2733 VDD2.n46 VDD2.n9 0.155672
R2734 VDD2.n53 VDD2.n9 0.155672
R2735 VDD2.n54 VDD2.n53 0.155672
R2736 VDD2.n54 VDD2.n5 0.155672
R2737 VDD2.n61 VDD2.n5 0.155672
R2738 VDD2.n62 VDD2.n61 0.155672
R2739 VDD2.n62 VDD2.n1 0.155672
R2740 VDD2.n69 VDD2.n1 0.155672
C0 VN VDD2 10.3531f
C1 VTAIL VDD2 11.6123f
C2 VN VDD1 0.151073f
C3 VP VN 7.13281f
C4 VTAIL VDD1 11.5702f
C5 VP VTAIL 10.5313f
C6 VN VTAIL 10.5169f
C7 VDD1 VDD2 1.51171f
C8 VP VDD2 0.453743f
C9 VP VDD1 10.651401f
C10 VDD2 B 6.233635f
C11 VDD1 B 6.211672f
C12 VTAIL B 7.859111f
C13 VN B 13.48592f
C14 VP B 11.82733f
C15 VDD2.n0 B 0.02955f
C16 VDD2.n1 B 0.022424f
C17 VDD2.n2 B 0.01205f
C18 VDD2.n3 B 0.028481f
C19 VDD2.n4 B 0.012758f
C20 VDD2.n5 B 0.022424f
C21 VDD2.n6 B 0.01205f
C22 VDD2.n7 B 0.028481f
C23 VDD2.n8 B 0.012758f
C24 VDD2.n9 B 0.022424f
C25 VDD2.n10 B 0.01205f
C26 VDD2.n11 B 0.028481f
C27 VDD2.n12 B 0.012758f
C28 VDD2.n13 B 0.022424f
C29 VDD2.n14 B 0.01205f
C30 VDD2.n15 B 0.028481f
C31 VDD2.n16 B 0.012758f
C32 VDD2.n17 B 0.022424f
C33 VDD2.n18 B 0.01205f
C34 VDD2.n19 B 0.028481f
C35 VDD2.n20 B 0.012758f
C36 VDD2.n21 B 1.28115f
C37 VDD2.n22 B 0.01205f
C38 VDD2.t8 B 0.046829f
C39 VDD2.n23 B 0.136528f
C40 VDD2.n24 B 0.016825f
C41 VDD2.n25 B 0.021361f
C42 VDD2.n26 B 0.028481f
C43 VDD2.n27 B 0.012758f
C44 VDD2.n28 B 0.01205f
C45 VDD2.n29 B 0.022424f
C46 VDD2.n30 B 0.022424f
C47 VDD2.n31 B 0.01205f
C48 VDD2.n32 B 0.012758f
C49 VDD2.n33 B 0.028481f
C50 VDD2.n34 B 0.028481f
C51 VDD2.n35 B 0.012758f
C52 VDD2.n36 B 0.01205f
C53 VDD2.n37 B 0.022424f
C54 VDD2.n38 B 0.022424f
C55 VDD2.n39 B 0.01205f
C56 VDD2.n40 B 0.012758f
C57 VDD2.n41 B 0.028481f
C58 VDD2.n42 B 0.028481f
C59 VDD2.n43 B 0.012758f
C60 VDD2.n44 B 0.01205f
C61 VDD2.n45 B 0.022424f
C62 VDD2.n46 B 0.022424f
C63 VDD2.n47 B 0.01205f
C64 VDD2.n48 B 0.012758f
C65 VDD2.n49 B 0.028481f
C66 VDD2.n50 B 0.028481f
C67 VDD2.n51 B 0.012758f
C68 VDD2.n52 B 0.01205f
C69 VDD2.n53 B 0.022424f
C70 VDD2.n54 B 0.022424f
C71 VDD2.n55 B 0.01205f
C72 VDD2.n56 B 0.012758f
C73 VDD2.n57 B 0.028481f
C74 VDD2.n58 B 0.028481f
C75 VDD2.n59 B 0.012758f
C76 VDD2.n60 B 0.01205f
C77 VDD2.n61 B 0.022424f
C78 VDD2.n62 B 0.022424f
C79 VDD2.n63 B 0.01205f
C80 VDD2.n64 B 0.012758f
C81 VDD2.n65 B 0.028481f
C82 VDD2.n66 B 0.057182f
C83 VDD2.n67 B 0.012758f
C84 VDD2.n68 B 0.023561f
C85 VDD2.n69 B 0.053976f
C86 VDD2.n70 B 0.078163f
C87 VDD2.t2 B 0.235146f
C88 VDD2.t1 B 0.235146f
C89 VDD2.n71 B 2.11415f
C90 VDD2.n72 B 0.484725f
C91 VDD2.t6 B 0.235146f
C92 VDD2.t3 B 0.235146f
C93 VDD2.n73 B 2.12145f
C94 VDD2.n74 B 2.19193f
C95 VDD2.n75 B 0.02955f
C96 VDD2.n76 B 0.022424f
C97 VDD2.n77 B 0.01205f
C98 VDD2.n78 B 0.028481f
C99 VDD2.n79 B 0.012758f
C100 VDD2.n80 B 0.022424f
C101 VDD2.n81 B 0.01205f
C102 VDD2.n82 B 0.028481f
C103 VDD2.n83 B 0.012758f
C104 VDD2.n84 B 0.022424f
C105 VDD2.n85 B 0.01205f
C106 VDD2.n86 B 0.028481f
C107 VDD2.n87 B 0.012758f
C108 VDD2.n88 B 0.022424f
C109 VDD2.n89 B 0.01205f
C110 VDD2.n90 B 0.028481f
C111 VDD2.n91 B 0.012758f
C112 VDD2.n92 B 0.022424f
C113 VDD2.n93 B 0.01205f
C114 VDD2.n94 B 0.028481f
C115 VDD2.n95 B 0.012758f
C116 VDD2.n96 B 1.28115f
C117 VDD2.n97 B 0.01205f
C118 VDD2.t9 B 0.046829f
C119 VDD2.n98 B 0.136528f
C120 VDD2.n99 B 0.016825f
C121 VDD2.n100 B 0.021361f
C122 VDD2.n101 B 0.028481f
C123 VDD2.n102 B 0.012758f
C124 VDD2.n103 B 0.01205f
C125 VDD2.n104 B 0.022424f
C126 VDD2.n105 B 0.022424f
C127 VDD2.n106 B 0.01205f
C128 VDD2.n107 B 0.012758f
C129 VDD2.n108 B 0.028481f
C130 VDD2.n109 B 0.028481f
C131 VDD2.n110 B 0.012758f
C132 VDD2.n111 B 0.01205f
C133 VDD2.n112 B 0.022424f
C134 VDD2.n113 B 0.022424f
C135 VDD2.n114 B 0.01205f
C136 VDD2.n115 B 0.012758f
C137 VDD2.n116 B 0.028481f
C138 VDD2.n117 B 0.028481f
C139 VDD2.n118 B 0.012758f
C140 VDD2.n119 B 0.01205f
C141 VDD2.n120 B 0.022424f
C142 VDD2.n121 B 0.022424f
C143 VDD2.n122 B 0.01205f
C144 VDD2.n123 B 0.012758f
C145 VDD2.n124 B 0.028481f
C146 VDD2.n125 B 0.028481f
C147 VDD2.n126 B 0.012758f
C148 VDD2.n127 B 0.01205f
C149 VDD2.n128 B 0.022424f
C150 VDD2.n129 B 0.022424f
C151 VDD2.n130 B 0.01205f
C152 VDD2.n131 B 0.012758f
C153 VDD2.n132 B 0.028481f
C154 VDD2.n133 B 0.028481f
C155 VDD2.n134 B 0.012758f
C156 VDD2.n135 B 0.01205f
C157 VDD2.n136 B 0.022424f
C158 VDD2.n137 B 0.022424f
C159 VDD2.n138 B 0.01205f
C160 VDD2.n139 B 0.012758f
C161 VDD2.n140 B 0.028481f
C162 VDD2.n141 B 0.057182f
C163 VDD2.n142 B 0.012758f
C164 VDD2.n143 B 0.023561f
C165 VDD2.n144 B 0.053976f
C166 VDD2.n145 B 0.072976f
C167 VDD2.n146 B 2.32657f
C168 VDD2.t5 B 0.235146f
C169 VDD2.t0 B 0.235146f
C170 VDD2.n147 B 2.11416f
C171 VDD2.n148 B 0.333269f
C172 VDD2.t7 B 0.235146f
C173 VDD2.t4 B 0.235146f
C174 VDD2.n149 B 2.12142f
C175 VN.n0 B 0.028843f
C176 VN.t6 B 1.65218f
C177 VN.n1 B 0.028621f
C178 VN.n2 B 0.028843f
C179 VN.t3 B 1.65218f
C180 VN.n3 B 0.038491f
C181 VN.n4 B 0.028843f
C182 VN.t8 B 1.65218f
C183 VN.n5 B 0.045725f
C184 VN.t1 B 1.74289f
C185 VN.n6 B 0.666862f
C186 VN.t7 B 1.65218f
C187 VN.n7 B 0.643296f
C188 VN.n8 B 0.035709f
C189 VN.n9 B 0.181147f
C190 VN.n10 B 0.028843f
C191 VN.n11 B 0.028843f
C192 VN.n12 B 0.038491f
C193 VN.n13 B 0.040486f
C194 VN.n14 B 0.591458f
C195 VN.n15 B 0.040486f
C196 VN.n16 B 0.028843f
C197 VN.n17 B 0.028843f
C198 VN.n18 B 0.028843f
C199 VN.n19 B 0.045725f
C200 VN.n20 B 0.035709f
C201 VN.n21 B 0.591458f
C202 VN.n22 B 0.048779f
C203 VN.n23 B 0.028843f
C204 VN.n24 B 0.028843f
C205 VN.n25 B 0.028843f
C206 VN.n26 B 0.052079f
C207 VN.n27 B 0.030932f
C208 VN.n28 B 0.646054f
C209 VN.n29 B 0.029474f
C210 VN.n30 B 0.028843f
C211 VN.t0 B 1.65218f
C212 VN.n31 B 0.028621f
C213 VN.n32 B 0.028843f
C214 VN.t4 B 1.65218f
C215 VN.n33 B 0.038491f
C216 VN.n34 B 0.028843f
C217 VN.t9 B 1.65218f
C218 VN.n35 B 0.045725f
C219 VN.t5 B 1.74289f
C220 VN.n36 B 0.666862f
C221 VN.t2 B 1.65218f
C222 VN.n37 B 0.643296f
C223 VN.n38 B 0.035709f
C224 VN.n39 B 0.181147f
C225 VN.n40 B 0.028843f
C226 VN.n41 B 0.028843f
C227 VN.n42 B 0.038491f
C228 VN.n43 B 0.040486f
C229 VN.n44 B 0.591458f
C230 VN.n45 B 0.040486f
C231 VN.n46 B 0.028843f
C232 VN.n47 B 0.028843f
C233 VN.n48 B 0.028843f
C234 VN.n49 B 0.045725f
C235 VN.n50 B 0.035709f
C236 VN.n51 B 0.591458f
C237 VN.n52 B 0.048779f
C238 VN.n53 B 0.028843f
C239 VN.n54 B 0.028843f
C240 VN.n55 B 0.028843f
C241 VN.n56 B 0.052079f
C242 VN.n57 B 0.030932f
C243 VN.n58 B 0.646054f
C244 VN.n59 B 1.51738f
C245 VTAIL.t8 B 0.253426f
C246 VTAIL.t3 B 0.253426f
C247 VTAIL.n0 B 2.20939f
C248 VTAIL.n1 B 0.432039f
C249 VTAIL.n2 B 0.031848f
C250 VTAIL.n3 B 0.024167f
C251 VTAIL.n4 B 0.012986f
C252 VTAIL.n5 B 0.030695f
C253 VTAIL.n6 B 0.01375f
C254 VTAIL.n7 B 0.024167f
C255 VTAIL.n8 B 0.012986f
C256 VTAIL.n9 B 0.030695f
C257 VTAIL.n10 B 0.01375f
C258 VTAIL.n11 B 0.024167f
C259 VTAIL.n12 B 0.012986f
C260 VTAIL.n13 B 0.030695f
C261 VTAIL.n14 B 0.01375f
C262 VTAIL.n15 B 0.024167f
C263 VTAIL.n16 B 0.012986f
C264 VTAIL.n17 B 0.030695f
C265 VTAIL.n18 B 0.01375f
C266 VTAIL.n19 B 0.024167f
C267 VTAIL.n20 B 0.012986f
C268 VTAIL.n21 B 0.030695f
C269 VTAIL.n22 B 0.01375f
C270 VTAIL.n23 B 1.38074f
C271 VTAIL.n24 B 0.012986f
C272 VTAIL.t18 B 0.050469f
C273 VTAIL.n25 B 0.147141f
C274 VTAIL.n26 B 0.018133f
C275 VTAIL.n27 B 0.023021f
C276 VTAIL.n28 B 0.030695f
C277 VTAIL.n29 B 0.01375f
C278 VTAIL.n30 B 0.012986f
C279 VTAIL.n31 B 0.024167f
C280 VTAIL.n32 B 0.024167f
C281 VTAIL.n33 B 0.012986f
C282 VTAIL.n34 B 0.01375f
C283 VTAIL.n35 B 0.030695f
C284 VTAIL.n36 B 0.030695f
C285 VTAIL.n37 B 0.01375f
C286 VTAIL.n38 B 0.012986f
C287 VTAIL.n39 B 0.024167f
C288 VTAIL.n40 B 0.024167f
C289 VTAIL.n41 B 0.012986f
C290 VTAIL.n42 B 0.01375f
C291 VTAIL.n43 B 0.030695f
C292 VTAIL.n44 B 0.030695f
C293 VTAIL.n45 B 0.01375f
C294 VTAIL.n46 B 0.012986f
C295 VTAIL.n47 B 0.024167f
C296 VTAIL.n48 B 0.024167f
C297 VTAIL.n49 B 0.012986f
C298 VTAIL.n50 B 0.01375f
C299 VTAIL.n51 B 0.030695f
C300 VTAIL.n52 B 0.030695f
C301 VTAIL.n53 B 0.01375f
C302 VTAIL.n54 B 0.012986f
C303 VTAIL.n55 B 0.024167f
C304 VTAIL.n56 B 0.024167f
C305 VTAIL.n57 B 0.012986f
C306 VTAIL.n58 B 0.01375f
C307 VTAIL.n59 B 0.030695f
C308 VTAIL.n60 B 0.030695f
C309 VTAIL.n61 B 0.01375f
C310 VTAIL.n62 B 0.012986f
C311 VTAIL.n63 B 0.024167f
C312 VTAIL.n64 B 0.024167f
C313 VTAIL.n65 B 0.012986f
C314 VTAIL.n66 B 0.01375f
C315 VTAIL.n67 B 0.030695f
C316 VTAIL.n68 B 0.061628f
C317 VTAIL.n69 B 0.01375f
C318 VTAIL.n70 B 0.025393f
C319 VTAIL.n71 B 0.058173f
C320 VTAIL.n72 B 0.06198f
C321 VTAIL.n73 B 0.250864f
C322 VTAIL.t17 B 0.253426f
C323 VTAIL.t11 B 0.253426f
C324 VTAIL.n74 B 2.20939f
C325 VTAIL.n75 B 0.487087f
C326 VTAIL.t13 B 0.253426f
C327 VTAIL.t16 B 0.253426f
C328 VTAIL.n76 B 2.20939f
C329 VTAIL.n77 B 1.83442f
C330 VTAIL.t0 B 0.253426f
C331 VTAIL.t6 B 0.253426f
C332 VTAIL.n78 B 2.2094f
C333 VTAIL.n79 B 1.83441f
C334 VTAIL.t5 B 0.253426f
C335 VTAIL.t9 B 0.253426f
C336 VTAIL.n80 B 2.2094f
C337 VTAIL.n81 B 0.487074f
C338 VTAIL.n82 B 0.031848f
C339 VTAIL.n83 B 0.024167f
C340 VTAIL.n84 B 0.012986f
C341 VTAIL.n85 B 0.030695f
C342 VTAIL.n86 B 0.01375f
C343 VTAIL.n87 B 0.024167f
C344 VTAIL.n88 B 0.012986f
C345 VTAIL.n89 B 0.030695f
C346 VTAIL.n90 B 0.01375f
C347 VTAIL.n91 B 0.024167f
C348 VTAIL.n92 B 0.012986f
C349 VTAIL.n93 B 0.030695f
C350 VTAIL.n94 B 0.01375f
C351 VTAIL.n95 B 0.024167f
C352 VTAIL.n96 B 0.012986f
C353 VTAIL.n97 B 0.030695f
C354 VTAIL.n98 B 0.01375f
C355 VTAIL.n99 B 0.024167f
C356 VTAIL.n100 B 0.012986f
C357 VTAIL.n101 B 0.030695f
C358 VTAIL.n102 B 0.01375f
C359 VTAIL.n103 B 1.38074f
C360 VTAIL.n104 B 0.012986f
C361 VTAIL.t2 B 0.050469f
C362 VTAIL.n105 B 0.147141f
C363 VTAIL.n106 B 0.018133f
C364 VTAIL.n107 B 0.023021f
C365 VTAIL.n108 B 0.030695f
C366 VTAIL.n109 B 0.01375f
C367 VTAIL.n110 B 0.012986f
C368 VTAIL.n111 B 0.024167f
C369 VTAIL.n112 B 0.024167f
C370 VTAIL.n113 B 0.012986f
C371 VTAIL.n114 B 0.01375f
C372 VTAIL.n115 B 0.030695f
C373 VTAIL.n116 B 0.030695f
C374 VTAIL.n117 B 0.01375f
C375 VTAIL.n118 B 0.012986f
C376 VTAIL.n119 B 0.024167f
C377 VTAIL.n120 B 0.024167f
C378 VTAIL.n121 B 0.012986f
C379 VTAIL.n122 B 0.01375f
C380 VTAIL.n123 B 0.030695f
C381 VTAIL.n124 B 0.030695f
C382 VTAIL.n125 B 0.01375f
C383 VTAIL.n126 B 0.012986f
C384 VTAIL.n127 B 0.024167f
C385 VTAIL.n128 B 0.024167f
C386 VTAIL.n129 B 0.012986f
C387 VTAIL.n130 B 0.01375f
C388 VTAIL.n131 B 0.030695f
C389 VTAIL.n132 B 0.030695f
C390 VTAIL.n133 B 0.01375f
C391 VTAIL.n134 B 0.012986f
C392 VTAIL.n135 B 0.024167f
C393 VTAIL.n136 B 0.024167f
C394 VTAIL.n137 B 0.012986f
C395 VTAIL.n138 B 0.01375f
C396 VTAIL.n139 B 0.030695f
C397 VTAIL.n140 B 0.030695f
C398 VTAIL.n141 B 0.01375f
C399 VTAIL.n142 B 0.012986f
C400 VTAIL.n143 B 0.024167f
C401 VTAIL.n144 B 0.024167f
C402 VTAIL.n145 B 0.012986f
C403 VTAIL.n146 B 0.01375f
C404 VTAIL.n147 B 0.030695f
C405 VTAIL.n148 B 0.061628f
C406 VTAIL.n149 B 0.01375f
C407 VTAIL.n150 B 0.025393f
C408 VTAIL.n151 B 0.058173f
C409 VTAIL.n152 B 0.06198f
C410 VTAIL.n153 B 0.250864f
C411 VTAIL.t14 B 0.253426f
C412 VTAIL.t19 B 0.253426f
C413 VTAIL.n154 B 2.2094f
C414 VTAIL.n155 B 0.45955f
C415 VTAIL.t12 B 0.253426f
C416 VTAIL.t15 B 0.253426f
C417 VTAIL.n156 B 2.2094f
C418 VTAIL.n157 B 0.487074f
C419 VTAIL.n158 B 0.031848f
C420 VTAIL.n159 B 0.024167f
C421 VTAIL.n160 B 0.012986f
C422 VTAIL.n161 B 0.030695f
C423 VTAIL.n162 B 0.01375f
C424 VTAIL.n163 B 0.024167f
C425 VTAIL.n164 B 0.012986f
C426 VTAIL.n165 B 0.030695f
C427 VTAIL.n166 B 0.01375f
C428 VTAIL.n167 B 0.024167f
C429 VTAIL.n168 B 0.012986f
C430 VTAIL.n169 B 0.030695f
C431 VTAIL.n170 B 0.01375f
C432 VTAIL.n171 B 0.024167f
C433 VTAIL.n172 B 0.012986f
C434 VTAIL.n173 B 0.030695f
C435 VTAIL.n174 B 0.01375f
C436 VTAIL.n175 B 0.024167f
C437 VTAIL.n176 B 0.012986f
C438 VTAIL.n177 B 0.030695f
C439 VTAIL.n178 B 0.01375f
C440 VTAIL.n179 B 1.38074f
C441 VTAIL.n180 B 0.012986f
C442 VTAIL.t10 B 0.050469f
C443 VTAIL.n181 B 0.147141f
C444 VTAIL.n182 B 0.018133f
C445 VTAIL.n183 B 0.023021f
C446 VTAIL.n184 B 0.030695f
C447 VTAIL.n185 B 0.01375f
C448 VTAIL.n186 B 0.012986f
C449 VTAIL.n187 B 0.024167f
C450 VTAIL.n188 B 0.024167f
C451 VTAIL.n189 B 0.012986f
C452 VTAIL.n190 B 0.01375f
C453 VTAIL.n191 B 0.030695f
C454 VTAIL.n192 B 0.030695f
C455 VTAIL.n193 B 0.01375f
C456 VTAIL.n194 B 0.012986f
C457 VTAIL.n195 B 0.024167f
C458 VTAIL.n196 B 0.024167f
C459 VTAIL.n197 B 0.012986f
C460 VTAIL.n198 B 0.01375f
C461 VTAIL.n199 B 0.030695f
C462 VTAIL.n200 B 0.030695f
C463 VTAIL.n201 B 0.01375f
C464 VTAIL.n202 B 0.012986f
C465 VTAIL.n203 B 0.024167f
C466 VTAIL.n204 B 0.024167f
C467 VTAIL.n205 B 0.012986f
C468 VTAIL.n206 B 0.01375f
C469 VTAIL.n207 B 0.030695f
C470 VTAIL.n208 B 0.030695f
C471 VTAIL.n209 B 0.01375f
C472 VTAIL.n210 B 0.012986f
C473 VTAIL.n211 B 0.024167f
C474 VTAIL.n212 B 0.024167f
C475 VTAIL.n213 B 0.012986f
C476 VTAIL.n214 B 0.01375f
C477 VTAIL.n215 B 0.030695f
C478 VTAIL.n216 B 0.030695f
C479 VTAIL.n217 B 0.01375f
C480 VTAIL.n218 B 0.012986f
C481 VTAIL.n219 B 0.024167f
C482 VTAIL.n220 B 0.024167f
C483 VTAIL.n221 B 0.012986f
C484 VTAIL.n222 B 0.01375f
C485 VTAIL.n223 B 0.030695f
C486 VTAIL.n224 B 0.061628f
C487 VTAIL.n225 B 0.01375f
C488 VTAIL.n226 B 0.025393f
C489 VTAIL.n227 B 0.058173f
C490 VTAIL.n228 B 0.06198f
C491 VTAIL.n229 B 1.4975f
C492 VTAIL.n230 B 0.031848f
C493 VTAIL.n231 B 0.024167f
C494 VTAIL.n232 B 0.012986f
C495 VTAIL.n233 B 0.030695f
C496 VTAIL.n234 B 0.01375f
C497 VTAIL.n235 B 0.024167f
C498 VTAIL.n236 B 0.012986f
C499 VTAIL.n237 B 0.030695f
C500 VTAIL.n238 B 0.01375f
C501 VTAIL.n239 B 0.024167f
C502 VTAIL.n240 B 0.012986f
C503 VTAIL.n241 B 0.030695f
C504 VTAIL.n242 B 0.01375f
C505 VTAIL.n243 B 0.024167f
C506 VTAIL.n244 B 0.012986f
C507 VTAIL.n245 B 0.030695f
C508 VTAIL.n246 B 0.01375f
C509 VTAIL.n247 B 0.024167f
C510 VTAIL.n248 B 0.012986f
C511 VTAIL.n249 B 0.030695f
C512 VTAIL.n250 B 0.01375f
C513 VTAIL.n251 B 1.38074f
C514 VTAIL.n252 B 0.012986f
C515 VTAIL.t4 B 0.050469f
C516 VTAIL.n253 B 0.147141f
C517 VTAIL.n254 B 0.018133f
C518 VTAIL.n255 B 0.023021f
C519 VTAIL.n256 B 0.030695f
C520 VTAIL.n257 B 0.01375f
C521 VTAIL.n258 B 0.012986f
C522 VTAIL.n259 B 0.024167f
C523 VTAIL.n260 B 0.024167f
C524 VTAIL.n261 B 0.012986f
C525 VTAIL.n262 B 0.01375f
C526 VTAIL.n263 B 0.030695f
C527 VTAIL.n264 B 0.030695f
C528 VTAIL.n265 B 0.01375f
C529 VTAIL.n266 B 0.012986f
C530 VTAIL.n267 B 0.024167f
C531 VTAIL.n268 B 0.024167f
C532 VTAIL.n269 B 0.012986f
C533 VTAIL.n270 B 0.01375f
C534 VTAIL.n271 B 0.030695f
C535 VTAIL.n272 B 0.030695f
C536 VTAIL.n273 B 0.01375f
C537 VTAIL.n274 B 0.012986f
C538 VTAIL.n275 B 0.024167f
C539 VTAIL.n276 B 0.024167f
C540 VTAIL.n277 B 0.012986f
C541 VTAIL.n278 B 0.01375f
C542 VTAIL.n279 B 0.030695f
C543 VTAIL.n280 B 0.030695f
C544 VTAIL.n281 B 0.01375f
C545 VTAIL.n282 B 0.012986f
C546 VTAIL.n283 B 0.024167f
C547 VTAIL.n284 B 0.024167f
C548 VTAIL.n285 B 0.012986f
C549 VTAIL.n286 B 0.01375f
C550 VTAIL.n287 B 0.030695f
C551 VTAIL.n288 B 0.030695f
C552 VTAIL.n289 B 0.01375f
C553 VTAIL.n290 B 0.012986f
C554 VTAIL.n291 B 0.024167f
C555 VTAIL.n292 B 0.024167f
C556 VTAIL.n293 B 0.012986f
C557 VTAIL.n294 B 0.01375f
C558 VTAIL.n295 B 0.030695f
C559 VTAIL.n296 B 0.061628f
C560 VTAIL.n297 B 0.01375f
C561 VTAIL.n298 B 0.025393f
C562 VTAIL.n299 B 0.058173f
C563 VTAIL.n300 B 0.06198f
C564 VTAIL.n301 B 1.4975f
C565 VTAIL.t1 B 0.253426f
C566 VTAIL.t7 B 0.253426f
C567 VTAIL.n302 B 2.20939f
C568 VTAIL.n303 B 0.38639f
C569 VDD1.n0 B 0.029841f
C570 VDD1.n1 B 0.022645f
C571 VDD1.n2 B 0.012168f
C572 VDD1.n3 B 0.028761f
C573 VDD1.n4 B 0.012884f
C574 VDD1.n5 B 0.022645f
C575 VDD1.n6 B 0.012168f
C576 VDD1.n7 B 0.028761f
C577 VDD1.n8 B 0.012884f
C578 VDD1.n9 B 0.022645f
C579 VDD1.n10 B 0.012168f
C580 VDD1.n11 B 0.028761f
C581 VDD1.n12 B 0.012884f
C582 VDD1.n13 B 0.022645f
C583 VDD1.n14 B 0.012168f
C584 VDD1.n15 B 0.028761f
C585 VDD1.n16 B 0.012884f
C586 VDD1.n17 B 0.022645f
C587 VDD1.n18 B 0.012168f
C588 VDD1.n19 B 0.028761f
C589 VDD1.n20 B 0.012884f
C590 VDD1.n21 B 1.29375f
C591 VDD1.n22 B 0.012168f
C592 VDD1.t8 B 0.047289f
C593 VDD1.n23 B 0.13787f
C594 VDD1.n24 B 0.01699f
C595 VDD1.n25 B 0.021571f
C596 VDD1.n26 B 0.028761f
C597 VDD1.n27 B 0.012884f
C598 VDD1.n28 B 0.012168f
C599 VDD1.n29 B 0.022645f
C600 VDD1.n30 B 0.022645f
C601 VDD1.n31 B 0.012168f
C602 VDD1.n32 B 0.012884f
C603 VDD1.n33 B 0.028761f
C604 VDD1.n34 B 0.028761f
C605 VDD1.n35 B 0.012884f
C606 VDD1.n36 B 0.012168f
C607 VDD1.n37 B 0.022645f
C608 VDD1.n38 B 0.022645f
C609 VDD1.n39 B 0.012168f
C610 VDD1.n40 B 0.012884f
C611 VDD1.n41 B 0.028761f
C612 VDD1.n42 B 0.028761f
C613 VDD1.n43 B 0.012884f
C614 VDD1.n44 B 0.012168f
C615 VDD1.n45 B 0.022645f
C616 VDD1.n46 B 0.022645f
C617 VDD1.n47 B 0.012168f
C618 VDD1.n48 B 0.012884f
C619 VDD1.n49 B 0.028761f
C620 VDD1.n50 B 0.028761f
C621 VDD1.n51 B 0.012884f
C622 VDD1.n52 B 0.012168f
C623 VDD1.n53 B 0.022645f
C624 VDD1.n54 B 0.022645f
C625 VDD1.n55 B 0.012168f
C626 VDD1.n56 B 0.012884f
C627 VDD1.n57 B 0.028761f
C628 VDD1.n58 B 0.028761f
C629 VDD1.n59 B 0.012884f
C630 VDD1.n60 B 0.012168f
C631 VDD1.n61 B 0.022645f
C632 VDD1.n62 B 0.022645f
C633 VDD1.n63 B 0.012168f
C634 VDD1.n64 B 0.012884f
C635 VDD1.n65 B 0.028761f
C636 VDD1.n66 B 0.057745f
C637 VDD1.n67 B 0.012884f
C638 VDD1.n68 B 0.023793f
C639 VDD1.n69 B 0.054507f
C640 VDD1.n70 B 0.078931f
C641 VDD1.t2 B 0.237459f
C642 VDD1.t7 B 0.237459f
C643 VDD1.n71 B 2.13495f
C644 VDD1.n72 B 0.496294f
C645 VDD1.n73 B 0.029841f
C646 VDD1.n74 B 0.022645f
C647 VDD1.n75 B 0.012168f
C648 VDD1.n76 B 0.028761f
C649 VDD1.n77 B 0.012884f
C650 VDD1.n78 B 0.022645f
C651 VDD1.n79 B 0.012168f
C652 VDD1.n80 B 0.028761f
C653 VDD1.n81 B 0.012884f
C654 VDD1.n82 B 0.022645f
C655 VDD1.n83 B 0.012168f
C656 VDD1.n84 B 0.028761f
C657 VDD1.n85 B 0.012884f
C658 VDD1.n86 B 0.022645f
C659 VDD1.n87 B 0.012168f
C660 VDD1.n88 B 0.028761f
C661 VDD1.n89 B 0.012884f
C662 VDD1.n90 B 0.022645f
C663 VDD1.n91 B 0.012168f
C664 VDD1.n92 B 0.028761f
C665 VDD1.n93 B 0.012884f
C666 VDD1.n94 B 1.29375f
C667 VDD1.n95 B 0.012168f
C668 VDD1.t0 B 0.047289f
C669 VDD1.n96 B 0.13787f
C670 VDD1.n97 B 0.01699f
C671 VDD1.n98 B 0.021571f
C672 VDD1.n99 B 0.028761f
C673 VDD1.n100 B 0.012884f
C674 VDD1.n101 B 0.012168f
C675 VDD1.n102 B 0.022645f
C676 VDD1.n103 B 0.022645f
C677 VDD1.n104 B 0.012168f
C678 VDD1.n105 B 0.012884f
C679 VDD1.n106 B 0.028761f
C680 VDD1.n107 B 0.028761f
C681 VDD1.n108 B 0.012884f
C682 VDD1.n109 B 0.012168f
C683 VDD1.n110 B 0.022645f
C684 VDD1.n111 B 0.022645f
C685 VDD1.n112 B 0.012168f
C686 VDD1.n113 B 0.012884f
C687 VDD1.n114 B 0.028761f
C688 VDD1.n115 B 0.028761f
C689 VDD1.n116 B 0.012884f
C690 VDD1.n117 B 0.012168f
C691 VDD1.n118 B 0.022645f
C692 VDD1.n119 B 0.022645f
C693 VDD1.n120 B 0.012168f
C694 VDD1.n121 B 0.012884f
C695 VDD1.n122 B 0.028761f
C696 VDD1.n123 B 0.028761f
C697 VDD1.n124 B 0.012884f
C698 VDD1.n125 B 0.012168f
C699 VDD1.n126 B 0.022645f
C700 VDD1.n127 B 0.022645f
C701 VDD1.n128 B 0.012168f
C702 VDD1.n129 B 0.012884f
C703 VDD1.n130 B 0.028761f
C704 VDD1.n131 B 0.028761f
C705 VDD1.n132 B 0.012884f
C706 VDD1.n133 B 0.012168f
C707 VDD1.n134 B 0.022645f
C708 VDD1.n135 B 0.022645f
C709 VDD1.n136 B 0.012168f
C710 VDD1.n137 B 0.012884f
C711 VDD1.n138 B 0.028761f
C712 VDD1.n139 B 0.057745f
C713 VDD1.n140 B 0.012884f
C714 VDD1.n141 B 0.023793f
C715 VDD1.n142 B 0.054507f
C716 VDD1.n143 B 0.078931f
C717 VDD1.t5 B 0.237459f
C718 VDD1.t1 B 0.237459f
C719 VDD1.n144 B 2.13494f
C720 VDD1.n145 B 0.489492f
C721 VDD1.t3 B 0.237459f
C722 VDD1.t4 B 0.237459f
C723 VDD1.n146 B 2.14232f
C724 VDD1.n147 B 2.30325f
C725 VDD1.t6 B 0.237459f
C726 VDD1.t9 B 0.237459f
C727 VDD1.n148 B 2.13494f
C728 VDD1.n149 B 2.5756f
C729 VP.n0 B 0.029194f
C730 VP.t1 B 1.67231f
C731 VP.n1 B 0.028969f
C732 VP.n2 B 0.029194f
C733 VP.t8 B 1.67231f
C734 VP.n3 B 0.03896f
C735 VP.n4 B 0.029194f
C736 VP.t2 B 1.67231f
C737 VP.n5 B 0.046282f
C738 VP.n6 B 0.029194f
C739 VP.t3 B 1.67231f
C740 VP.n7 B 0.052714f
C741 VP.n8 B 0.029194f
C742 VP.t9 B 1.67231f
C743 VP.n9 B 0.028969f
C744 VP.n10 B 0.029194f
C745 VP.t4 B 1.67231f
C746 VP.n11 B 0.03896f
C747 VP.n12 B 0.029194f
C748 VP.t7 B 1.67231f
C749 VP.n13 B 0.046282f
C750 VP.t5 B 1.76412f
C751 VP.n14 B 0.674984f
C752 VP.t0 B 1.67231f
C753 VP.n15 B 0.651131f
C754 VP.n16 B 0.036144f
C755 VP.n17 B 0.183354f
C756 VP.n18 B 0.029194f
C757 VP.n19 B 0.029194f
C758 VP.n20 B 0.03896f
C759 VP.n21 B 0.040979f
C760 VP.n22 B 0.598662f
C761 VP.n23 B 0.040979f
C762 VP.n24 B 0.029194f
C763 VP.n25 B 0.029194f
C764 VP.n26 B 0.029194f
C765 VP.n27 B 0.046282f
C766 VP.n28 B 0.036144f
C767 VP.n29 B 0.598662f
C768 VP.n30 B 0.049374f
C769 VP.n31 B 0.029194f
C770 VP.n32 B 0.029194f
C771 VP.n33 B 0.029194f
C772 VP.n34 B 0.052714f
C773 VP.n35 B 0.031309f
C774 VP.n36 B 0.653922f
C775 VP.n37 B 1.51685f
C776 VP.n38 B 1.53855f
C777 VP.t6 B 1.67231f
C778 VP.n39 B 0.653922f
C779 VP.n40 B 0.031309f
C780 VP.n41 B 0.029194f
C781 VP.n42 B 0.029194f
C782 VP.n43 B 0.029194f
C783 VP.n44 B 0.028969f
C784 VP.n45 B 0.049374f
C785 VP.n46 B 0.598662f
C786 VP.n47 B 0.036144f
C787 VP.n48 B 0.029194f
C788 VP.n49 B 0.029194f
C789 VP.n50 B 0.029194f
C790 VP.n51 B 0.03896f
C791 VP.n52 B 0.040979f
C792 VP.n53 B 0.598662f
C793 VP.n54 B 0.040979f
C794 VP.n55 B 0.029194f
C795 VP.n56 B 0.029194f
C796 VP.n57 B 0.029194f
C797 VP.n58 B 0.046282f
C798 VP.n59 B 0.036144f
C799 VP.n60 B 0.598662f
C800 VP.n61 B 0.049374f
C801 VP.n62 B 0.029194f
C802 VP.n63 B 0.029194f
C803 VP.n64 B 0.029194f
C804 VP.n65 B 0.052714f
C805 VP.n66 B 0.031309f
C806 VP.n67 B 0.653922f
C807 VP.n68 B 0.029833f
.ends

