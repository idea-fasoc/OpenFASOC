* NGSPICE file created from diff_pair_sample_0915.ext - technology: sky130A

.subckt diff_pair_sample_0915 VTAIL VN VP B VDD2 VDD1
X0 B.t11 B.t9 B.t10 w_n2470_n2220# sky130_fd_pr__pfet_01v8 ad=2.4414 pd=13.3 as=0 ps=0 w=6.26 l=2.17
X1 B.t8 B.t6 B.t7 w_n2470_n2220# sky130_fd_pr__pfet_01v8 ad=2.4414 pd=13.3 as=0 ps=0 w=6.26 l=2.17
X2 VTAIL.t7 VP.t0 VDD1.t1 w_n2470_n2220# sky130_fd_pr__pfet_01v8 ad=2.4414 pd=13.3 as=1.0329 ps=6.59 w=6.26 l=2.17
X3 B.t5 B.t3 B.t4 w_n2470_n2220# sky130_fd_pr__pfet_01v8 ad=2.4414 pd=13.3 as=0 ps=0 w=6.26 l=2.17
X4 VTAIL.t3 VN.t0 VDD2.t3 w_n2470_n2220# sky130_fd_pr__pfet_01v8 ad=2.4414 pd=13.3 as=1.0329 ps=6.59 w=6.26 l=2.17
X5 VDD1.t3 VP.t1 VTAIL.t6 w_n2470_n2220# sky130_fd_pr__pfet_01v8 ad=1.0329 pd=6.59 as=2.4414 ps=13.3 w=6.26 l=2.17
X6 VDD2.t2 VN.t1 VTAIL.t1 w_n2470_n2220# sky130_fd_pr__pfet_01v8 ad=1.0329 pd=6.59 as=2.4414 ps=13.3 w=6.26 l=2.17
X7 VDD1.t0 VP.t2 VTAIL.t5 w_n2470_n2220# sky130_fd_pr__pfet_01v8 ad=1.0329 pd=6.59 as=2.4414 ps=13.3 w=6.26 l=2.17
X8 B.t2 B.t0 B.t1 w_n2470_n2220# sky130_fd_pr__pfet_01v8 ad=2.4414 pd=13.3 as=0 ps=0 w=6.26 l=2.17
X9 VDD2.t1 VN.t2 VTAIL.t2 w_n2470_n2220# sky130_fd_pr__pfet_01v8 ad=1.0329 pd=6.59 as=2.4414 ps=13.3 w=6.26 l=2.17
X10 VTAIL.t4 VP.t3 VDD1.t2 w_n2470_n2220# sky130_fd_pr__pfet_01v8 ad=2.4414 pd=13.3 as=1.0329 ps=6.59 w=6.26 l=2.17
X11 VTAIL.t0 VN.t3 VDD2.t0 w_n2470_n2220# sky130_fd_pr__pfet_01v8 ad=2.4414 pd=13.3 as=1.0329 ps=6.59 w=6.26 l=2.17
R0 B.n356 B.n355 585
R1 B.n357 B.n50 585
R2 B.n359 B.n358 585
R3 B.n360 B.n49 585
R4 B.n362 B.n361 585
R5 B.n363 B.n48 585
R6 B.n365 B.n364 585
R7 B.n366 B.n47 585
R8 B.n368 B.n367 585
R9 B.n369 B.n46 585
R10 B.n371 B.n370 585
R11 B.n372 B.n45 585
R12 B.n374 B.n373 585
R13 B.n375 B.n44 585
R14 B.n377 B.n376 585
R15 B.n378 B.n43 585
R16 B.n380 B.n379 585
R17 B.n381 B.n42 585
R18 B.n383 B.n382 585
R19 B.n384 B.n41 585
R20 B.n386 B.n385 585
R21 B.n387 B.n40 585
R22 B.n389 B.n388 585
R23 B.n390 B.n39 585
R24 B.n392 B.n391 585
R25 B.n394 B.n393 585
R26 B.n395 B.n35 585
R27 B.n397 B.n396 585
R28 B.n398 B.n34 585
R29 B.n400 B.n399 585
R30 B.n401 B.n33 585
R31 B.n403 B.n402 585
R32 B.n404 B.n32 585
R33 B.n406 B.n405 585
R34 B.n408 B.n29 585
R35 B.n410 B.n409 585
R36 B.n411 B.n28 585
R37 B.n413 B.n412 585
R38 B.n414 B.n27 585
R39 B.n416 B.n415 585
R40 B.n417 B.n26 585
R41 B.n419 B.n418 585
R42 B.n420 B.n25 585
R43 B.n422 B.n421 585
R44 B.n423 B.n24 585
R45 B.n425 B.n424 585
R46 B.n426 B.n23 585
R47 B.n428 B.n427 585
R48 B.n429 B.n22 585
R49 B.n431 B.n430 585
R50 B.n432 B.n21 585
R51 B.n434 B.n433 585
R52 B.n435 B.n20 585
R53 B.n437 B.n436 585
R54 B.n438 B.n19 585
R55 B.n440 B.n439 585
R56 B.n441 B.n18 585
R57 B.n443 B.n442 585
R58 B.n444 B.n17 585
R59 B.n354 B.n51 585
R60 B.n353 B.n352 585
R61 B.n351 B.n52 585
R62 B.n350 B.n349 585
R63 B.n348 B.n53 585
R64 B.n347 B.n346 585
R65 B.n345 B.n54 585
R66 B.n344 B.n343 585
R67 B.n342 B.n55 585
R68 B.n341 B.n340 585
R69 B.n339 B.n56 585
R70 B.n338 B.n337 585
R71 B.n336 B.n57 585
R72 B.n335 B.n334 585
R73 B.n333 B.n58 585
R74 B.n332 B.n331 585
R75 B.n330 B.n59 585
R76 B.n329 B.n328 585
R77 B.n327 B.n60 585
R78 B.n326 B.n325 585
R79 B.n324 B.n61 585
R80 B.n323 B.n322 585
R81 B.n321 B.n62 585
R82 B.n320 B.n319 585
R83 B.n318 B.n63 585
R84 B.n317 B.n316 585
R85 B.n315 B.n64 585
R86 B.n314 B.n313 585
R87 B.n312 B.n65 585
R88 B.n311 B.n310 585
R89 B.n309 B.n66 585
R90 B.n308 B.n307 585
R91 B.n306 B.n67 585
R92 B.n305 B.n304 585
R93 B.n303 B.n68 585
R94 B.n302 B.n301 585
R95 B.n300 B.n69 585
R96 B.n299 B.n298 585
R97 B.n297 B.n70 585
R98 B.n296 B.n295 585
R99 B.n294 B.n71 585
R100 B.n293 B.n292 585
R101 B.n291 B.n72 585
R102 B.n290 B.n289 585
R103 B.n288 B.n73 585
R104 B.n287 B.n286 585
R105 B.n285 B.n74 585
R106 B.n284 B.n283 585
R107 B.n282 B.n75 585
R108 B.n281 B.n280 585
R109 B.n279 B.n76 585
R110 B.n278 B.n277 585
R111 B.n276 B.n77 585
R112 B.n275 B.n274 585
R113 B.n273 B.n78 585
R114 B.n272 B.n271 585
R115 B.n270 B.n79 585
R116 B.n269 B.n268 585
R117 B.n267 B.n80 585
R118 B.n266 B.n265 585
R119 B.n264 B.n81 585
R120 B.n174 B.n115 585
R121 B.n176 B.n175 585
R122 B.n177 B.n114 585
R123 B.n179 B.n178 585
R124 B.n180 B.n113 585
R125 B.n182 B.n181 585
R126 B.n183 B.n112 585
R127 B.n185 B.n184 585
R128 B.n186 B.n111 585
R129 B.n188 B.n187 585
R130 B.n189 B.n110 585
R131 B.n191 B.n190 585
R132 B.n192 B.n109 585
R133 B.n194 B.n193 585
R134 B.n195 B.n108 585
R135 B.n197 B.n196 585
R136 B.n198 B.n107 585
R137 B.n200 B.n199 585
R138 B.n201 B.n106 585
R139 B.n203 B.n202 585
R140 B.n204 B.n105 585
R141 B.n206 B.n205 585
R142 B.n207 B.n104 585
R143 B.n209 B.n208 585
R144 B.n210 B.n101 585
R145 B.n213 B.n212 585
R146 B.n214 B.n100 585
R147 B.n216 B.n215 585
R148 B.n217 B.n99 585
R149 B.n219 B.n218 585
R150 B.n220 B.n98 585
R151 B.n222 B.n221 585
R152 B.n223 B.n97 585
R153 B.n225 B.n224 585
R154 B.n227 B.n226 585
R155 B.n228 B.n93 585
R156 B.n230 B.n229 585
R157 B.n231 B.n92 585
R158 B.n233 B.n232 585
R159 B.n234 B.n91 585
R160 B.n236 B.n235 585
R161 B.n237 B.n90 585
R162 B.n239 B.n238 585
R163 B.n240 B.n89 585
R164 B.n242 B.n241 585
R165 B.n243 B.n88 585
R166 B.n245 B.n244 585
R167 B.n246 B.n87 585
R168 B.n248 B.n247 585
R169 B.n249 B.n86 585
R170 B.n251 B.n250 585
R171 B.n252 B.n85 585
R172 B.n254 B.n253 585
R173 B.n255 B.n84 585
R174 B.n257 B.n256 585
R175 B.n258 B.n83 585
R176 B.n260 B.n259 585
R177 B.n261 B.n82 585
R178 B.n263 B.n262 585
R179 B.n173 B.n172 585
R180 B.n171 B.n116 585
R181 B.n170 B.n169 585
R182 B.n168 B.n117 585
R183 B.n167 B.n166 585
R184 B.n165 B.n118 585
R185 B.n164 B.n163 585
R186 B.n162 B.n119 585
R187 B.n161 B.n160 585
R188 B.n159 B.n120 585
R189 B.n158 B.n157 585
R190 B.n156 B.n121 585
R191 B.n155 B.n154 585
R192 B.n153 B.n122 585
R193 B.n152 B.n151 585
R194 B.n150 B.n123 585
R195 B.n149 B.n148 585
R196 B.n147 B.n124 585
R197 B.n146 B.n145 585
R198 B.n144 B.n125 585
R199 B.n143 B.n142 585
R200 B.n141 B.n126 585
R201 B.n140 B.n139 585
R202 B.n138 B.n127 585
R203 B.n137 B.n136 585
R204 B.n135 B.n128 585
R205 B.n134 B.n133 585
R206 B.n132 B.n129 585
R207 B.n131 B.n130 585
R208 B.n2 B.n0 585
R209 B.n489 B.n1 585
R210 B.n488 B.n487 585
R211 B.n486 B.n3 585
R212 B.n485 B.n484 585
R213 B.n483 B.n4 585
R214 B.n482 B.n481 585
R215 B.n480 B.n5 585
R216 B.n479 B.n478 585
R217 B.n477 B.n6 585
R218 B.n476 B.n475 585
R219 B.n474 B.n7 585
R220 B.n473 B.n472 585
R221 B.n471 B.n8 585
R222 B.n470 B.n469 585
R223 B.n468 B.n9 585
R224 B.n467 B.n466 585
R225 B.n465 B.n10 585
R226 B.n464 B.n463 585
R227 B.n462 B.n11 585
R228 B.n461 B.n460 585
R229 B.n459 B.n12 585
R230 B.n458 B.n457 585
R231 B.n456 B.n13 585
R232 B.n455 B.n454 585
R233 B.n453 B.n14 585
R234 B.n452 B.n451 585
R235 B.n450 B.n15 585
R236 B.n449 B.n448 585
R237 B.n447 B.n16 585
R238 B.n446 B.n445 585
R239 B.n491 B.n490 585
R240 B.n172 B.n115 530.939
R241 B.n446 B.n17 530.939
R242 B.n262 B.n81 530.939
R243 B.n356 B.n51 530.939
R244 B.n94 B.t6 276.815
R245 B.n102 B.t9 276.815
R246 B.n30 B.t0 276.815
R247 B.n36 B.t3 276.815
R248 B.n172 B.n171 163.367
R249 B.n171 B.n170 163.367
R250 B.n170 B.n117 163.367
R251 B.n166 B.n117 163.367
R252 B.n166 B.n165 163.367
R253 B.n165 B.n164 163.367
R254 B.n164 B.n119 163.367
R255 B.n160 B.n119 163.367
R256 B.n160 B.n159 163.367
R257 B.n159 B.n158 163.367
R258 B.n158 B.n121 163.367
R259 B.n154 B.n121 163.367
R260 B.n154 B.n153 163.367
R261 B.n153 B.n152 163.367
R262 B.n152 B.n123 163.367
R263 B.n148 B.n123 163.367
R264 B.n148 B.n147 163.367
R265 B.n147 B.n146 163.367
R266 B.n146 B.n125 163.367
R267 B.n142 B.n125 163.367
R268 B.n142 B.n141 163.367
R269 B.n141 B.n140 163.367
R270 B.n140 B.n127 163.367
R271 B.n136 B.n127 163.367
R272 B.n136 B.n135 163.367
R273 B.n135 B.n134 163.367
R274 B.n134 B.n129 163.367
R275 B.n130 B.n129 163.367
R276 B.n130 B.n2 163.367
R277 B.n490 B.n2 163.367
R278 B.n490 B.n489 163.367
R279 B.n489 B.n488 163.367
R280 B.n488 B.n3 163.367
R281 B.n484 B.n3 163.367
R282 B.n484 B.n483 163.367
R283 B.n483 B.n482 163.367
R284 B.n482 B.n5 163.367
R285 B.n478 B.n5 163.367
R286 B.n478 B.n477 163.367
R287 B.n477 B.n476 163.367
R288 B.n476 B.n7 163.367
R289 B.n472 B.n7 163.367
R290 B.n472 B.n471 163.367
R291 B.n471 B.n470 163.367
R292 B.n470 B.n9 163.367
R293 B.n466 B.n9 163.367
R294 B.n466 B.n465 163.367
R295 B.n465 B.n464 163.367
R296 B.n464 B.n11 163.367
R297 B.n460 B.n11 163.367
R298 B.n460 B.n459 163.367
R299 B.n459 B.n458 163.367
R300 B.n458 B.n13 163.367
R301 B.n454 B.n13 163.367
R302 B.n454 B.n453 163.367
R303 B.n453 B.n452 163.367
R304 B.n452 B.n15 163.367
R305 B.n448 B.n15 163.367
R306 B.n448 B.n447 163.367
R307 B.n447 B.n446 163.367
R308 B.n176 B.n115 163.367
R309 B.n177 B.n176 163.367
R310 B.n178 B.n177 163.367
R311 B.n178 B.n113 163.367
R312 B.n182 B.n113 163.367
R313 B.n183 B.n182 163.367
R314 B.n184 B.n183 163.367
R315 B.n184 B.n111 163.367
R316 B.n188 B.n111 163.367
R317 B.n189 B.n188 163.367
R318 B.n190 B.n189 163.367
R319 B.n190 B.n109 163.367
R320 B.n194 B.n109 163.367
R321 B.n195 B.n194 163.367
R322 B.n196 B.n195 163.367
R323 B.n196 B.n107 163.367
R324 B.n200 B.n107 163.367
R325 B.n201 B.n200 163.367
R326 B.n202 B.n201 163.367
R327 B.n202 B.n105 163.367
R328 B.n206 B.n105 163.367
R329 B.n207 B.n206 163.367
R330 B.n208 B.n207 163.367
R331 B.n208 B.n101 163.367
R332 B.n213 B.n101 163.367
R333 B.n214 B.n213 163.367
R334 B.n215 B.n214 163.367
R335 B.n215 B.n99 163.367
R336 B.n219 B.n99 163.367
R337 B.n220 B.n219 163.367
R338 B.n221 B.n220 163.367
R339 B.n221 B.n97 163.367
R340 B.n225 B.n97 163.367
R341 B.n226 B.n225 163.367
R342 B.n226 B.n93 163.367
R343 B.n230 B.n93 163.367
R344 B.n231 B.n230 163.367
R345 B.n232 B.n231 163.367
R346 B.n232 B.n91 163.367
R347 B.n236 B.n91 163.367
R348 B.n237 B.n236 163.367
R349 B.n238 B.n237 163.367
R350 B.n238 B.n89 163.367
R351 B.n242 B.n89 163.367
R352 B.n243 B.n242 163.367
R353 B.n244 B.n243 163.367
R354 B.n244 B.n87 163.367
R355 B.n248 B.n87 163.367
R356 B.n249 B.n248 163.367
R357 B.n250 B.n249 163.367
R358 B.n250 B.n85 163.367
R359 B.n254 B.n85 163.367
R360 B.n255 B.n254 163.367
R361 B.n256 B.n255 163.367
R362 B.n256 B.n83 163.367
R363 B.n260 B.n83 163.367
R364 B.n261 B.n260 163.367
R365 B.n262 B.n261 163.367
R366 B.n266 B.n81 163.367
R367 B.n267 B.n266 163.367
R368 B.n268 B.n267 163.367
R369 B.n268 B.n79 163.367
R370 B.n272 B.n79 163.367
R371 B.n273 B.n272 163.367
R372 B.n274 B.n273 163.367
R373 B.n274 B.n77 163.367
R374 B.n278 B.n77 163.367
R375 B.n279 B.n278 163.367
R376 B.n280 B.n279 163.367
R377 B.n280 B.n75 163.367
R378 B.n284 B.n75 163.367
R379 B.n285 B.n284 163.367
R380 B.n286 B.n285 163.367
R381 B.n286 B.n73 163.367
R382 B.n290 B.n73 163.367
R383 B.n291 B.n290 163.367
R384 B.n292 B.n291 163.367
R385 B.n292 B.n71 163.367
R386 B.n296 B.n71 163.367
R387 B.n297 B.n296 163.367
R388 B.n298 B.n297 163.367
R389 B.n298 B.n69 163.367
R390 B.n302 B.n69 163.367
R391 B.n303 B.n302 163.367
R392 B.n304 B.n303 163.367
R393 B.n304 B.n67 163.367
R394 B.n308 B.n67 163.367
R395 B.n309 B.n308 163.367
R396 B.n310 B.n309 163.367
R397 B.n310 B.n65 163.367
R398 B.n314 B.n65 163.367
R399 B.n315 B.n314 163.367
R400 B.n316 B.n315 163.367
R401 B.n316 B.n63 163.367
R402 B.n320 B.n63 163.367
R403 B.n321 B.n320 163.367
R404 B.n322 B.n321 163.367
R405 B.n322 B.n61 163.367
R406 B.n326 B.n61 163.367
R407 B.n327 B.n326 163.367
R408 B.n328 B.n327 163.367
R409 B.n328 B.n59 163.367
R410 B.n332 B.n59 163.367
R411 B.n333 B.n332 163.367
R412 B.n334 B.n333 163.367
R413 B.n334 B.n57 163.367
R414 B.n338 B.n57 163.367
R415 B.n339 B.n338 163.367
R416 B.n340 B.n339 163.367
R417 B.n340 B.n55 163.367
R418 B.n344 B.n55 163.367
R419 B.n345 B.n344 163.367
R420 B.n346 B.n345 163.367
R421 B.n346 B.n53 163.367
R422 B.n350 B.n53 163.367
R423 B.n351 B.n350 163.367
R424 B.n352 B.n351 163.367
R425 B.n352 B.n51 163.367
R426 B.n442 B.n17 163.367
R427 B.n442 B.n441 163.367
R428 B.n441 B.n440 163.367
R429 B.n440 B.n19 163.367
R430 B.n436 B.n19 163.367
R431 B.n436 B.n435 163.367
R432 B.n435 B.n434 163.367
R433 B.n434 B.n21 163.367
R434 B.n430 B.n21 163.367
R435 B.n430 B.n429 163.367
R436 B.n429 B.n428 163.367
R437 B.n428 B.n23 163.367
R438 B.n424 B.n23 163.367
R439 B.n424 B.n423 163.367
R440 B.n423 B.n422 163.367
R441 B.n422 B.n25 163.367
R442 B.n418 B.n25 163.367
R443 B.n418 B.n417 163.367
R444 B.n417 B.n416 163.367
R445 B.n416 B.n27 163.367
R446 B.n412 B.n27 163.367
R447 B.n412 B.n411 163.367
R448 B.n411 B.n410 163.367
R449 B.n410 B.n29 163.367
R450 B.n405 B.n29 163.367
R451 B.n405 B.n404 163.367
R452 B.n404 B.n403 163.367
R453 B.n403 B.n33 163.367
R454 B.n399 B.n33 163.367
R455 B.n399 B.n398 163.367
R456 B.n398 B.n397 163.367
R457 B.n397 B.n35 163.367
R458 B.n393 B.n35 163.367
R459 B.n393 B.n392 163.367
R460 B.n392 B.n39 163.367
R461 B.n388 B.n39 163.367
R462 B.n388 B.n387 163.367
R463 B.n387 B.n386 163.367
R464 B.n386 B.n41 163.367
R465 B.n382 B.n41 163.367
R466 B.n382 B.n381 163.367
R467 B.n381 B.n380 163.367
R468 B.n380 B.n43 163.367
R469 B.n376 B.n43 163.367
R470 B.n376 B.n375 163.367
R471 B.n375 B.n374 163.367
R472 B.n374 B.n45 163.367
R473 B.n370 B.n45 163.367
R474 B.n370 B.n369 163.367
R475 B.n369 B.n368 163.367
R476 B.n368 B.n47 163.367
R477 B.n364 B.n47 163.367
R478 B.n364 B.n363 163.367
R479 B.n363 B.n362 163.367
R480 B.n362 B.n49 163.367
R481 B.n358 B.n49 163.367
R482 B.n358 B.n357 163.367
R483 B.n357 B.n356 163.367
R484 B.n94 B.t8 161.855
R485 B.n36 B.t4 161.855
R486 B.n102 B.t11 161.847
R487 B.n30 B.t1 161.847
R488 B.n95 B.t7 113.37
R489 B.n37 B.t5 113.37
R490 B.n103 B.t10 113.362
R491 B.n31 B.t2 113.362
R492 B.n96 B.n95 59.5399
R493 B.n211 B.n103 59.5399
R494 B.n407 B.n31 59.5399
R495 B.n38 B.n37 59.5399
R496 B.n95 B.n94 48.4853
R497 B.n103 B.n102 48.4853
R498 B.n31 B.n30 48.4853
R499 B.n37 B.n36 48.4853
R500 B.n445 B.n444 34.4981
R501 B.n355 B.n354 34.4981
R502 B.n264 B.n263 34.4981
R503 B.n174 B.n173 34.4981
R504 B B.n491 18.0485
R505 B.n444 B.n443 10.6151
R506 B.n443 B.n18 10.6151
R507 B.n439 B.n18 10.6151
R508 B.n439 B.n438 10.6151
R509 B.n438 B.n437 10.6151
R510 B.n437 B.n20 10.6151
R511 B.n433 B.n20 10.6151
R512 B.n433 B.n432 10.6151
R513 B.n432 B.n431 10.6151
R514 B.n431 B.n22 10.6151
R515 B.n427 B.n22 10.6151
R516 B.n427 B.n426 10.6151
R517 B.n426 B.n425 10.6151
R518 B.n425 B.n24 10.6151
R519 B.n421 B.n24 10.6151
R520 B.n421 B.n420 10.6151
R521 B.n420 B.n419 10.6151
R522 B.n419 B.n26 10.6151
R523 B.n415 B.n26 10.6151
R524 B.n415 B.n414 10.6151
R525 B.n414 B.n413 10.6151
R526 B.n413 B.n28 10.6151
R527 B.n409 B.n28 10.6151
R528 B.n409 B.n408 10.6151
R529 B.n406 B.n32 10.6151
R530 B.n402 B.n32 10.6151
R531 B.n402 B.n401 10.6151
R532 B.n401 B.n400 10.6151
R533 B.n400 B.n34 10.6151
R534 B.n396 B.n34 10.6151
R535 B.n396 B.n395 10.6151
R536 B.n395 B.n394 10.6151
R537 B.n391 B.n390 10.6151
R538 B.n390 B.n389 10.6151
R539 B.n389 B.n40 10.6151
R540 B.n385 B.n40 10.6151
R541 B.n385 B.n384 10.6151
R542 B.n384 B.n383 10.6151
R543 B.n383 B.n42 10.6151
R544 B.n379 B.n42 10.6151
R545 B.n379 B.n378 10.6151
R546 B.n378 B.n377 10.6151
R547 B.n377 B.n44 10.6151
R548 B.n373 B.n44 10.6151
R549 B.n373 B.n372 10.6151
R550 B.n372 B.n371 10.6151
R551 B.n371 B.n46 10.6151
R552 B.n367 B.n46 10.6151
R553 B.n367 B.n366 10.6151
R554 B.n366 B.n365 10.6151
R555 B.n365 B.n48 10.6151
R556 B.n361 B.n48 10.6151
R557 B.n361 B.n360 10.6151
R558 B.n360 B.n359 10.6151
R559 B.n359 B.n50 10.6151
R560 B.n355 B.n50 10.6151
R561 B.n265 B.n264 10.6151
R562 B.n265 B.n80 10.6151
R563 B.n269 B.n80 10.6151
R564 B.n270 B.n269 10.6151
R565 B.n271 B.n270 10.6151
R566 B.n271 B.n78 10.6151
R567 B.n275 B.n78 10.6151
R568 B.n276 B.n275 10.6151
R569 B.n277 B.n276 10.6151
R570 B.n277 B.n76 10.6151
R571 B.n281 B.n76 10.6151
R572 B.n282 B.n281 10.6151
R573 B.n283 B.n282 10.6151
R574 B.n283 B.n74 10.6151
R575 B.n287 B.n74 10.6151
R576 B.n288 B.n287 10.6151
R577 B.n289 B.n288 10.6151
R578 B.n289 B.n72 10.6151
R579 B.n293 B.n72 10.6151
R580 B.n294 B.n293 10.6151
R581 B.n295 B.n294 10.6151
R582 B.n295 B.n70 10.6151
R583 B.n299 B.n70 10.6151
R584 B.n300 B.n299 10.6151
R585 B.n301 B.n300 10.6151
R586 B.n301 B.n68 10.6151
R587 B.n305 B.n68 10.6151
R588 B.n306 B.n305 10.6151
R589 B.n307 B.n306 10.6151
R590 B.n307 B.n66 10.6151
R591 B.n311 B.n66 10.6151
R592 B.n312 B.n311 10.6151
R593 B.n313 B.n312 10.6151
R594 B.n313 B.n64 10.6151
R595 B.n317 B.n64 10.6151
R596 B.n318 B.n317 10.6151
R597 B.n319 B.n318 10.6151
R598 B.n319 B.n62 10.6151
R599 B.n323 B.n62 10.6151
R600 B.n324 B.n323 10.6151
R601 B.n325 B.n324 10.6151
R602 B.n325 B.n60 10.6151
R603 B.n329 B.n60 10.6151
R604 B.n330 B.n329 10.6151
R605 B.n331 B.n330 10.6151
R606 B.n331 B.n58 10.6151
R607 B.n335 B.n58 10.6151
R608 B.n336 B.n335 10.6151
R609 B.n337 B.n336 10.6151
R610 B.n337 B.n56 10.6151
R611 B.n341 B.n56 10.6151
R612 B.n342 B.n341 10.6151
R613 B.n343 B.n342 10.6151
R614 B.n343 B.n54 10.6151
R615 B.n347 B.n54 10.6151
R616 B.n348 B.n347 10.6151
R617 B.n349 B.n348 10.6151
R618 B.n349 B.n52 10.6151
R619 B.n353 B.n52 10.6151
R620 B.n354 B.n353 10.6151
R621 B.n175 B.n174 10.6151
R622 B.n175 B.n114 10.6151
R623 B.n179 B.n114 10.6151
R624 B.n180 B.n179 10.6151
R625 B.n181 B.n180 10.6151
R626 B.n181 B.n112 10.6151
R627 B.n185 B.n112 10.6151
R628 B.n186 B.n185 10.6151
R629 B.n187 B.n186 10.6151
R630 B.n187 B.n110 10.6151
R631 B.n191 B.n110 10.6151
R632 B.n192 B.n191 10.6151
R633 B.n193 B.n192 10.6151
R634 B.n193 B.n108 10.6151
R635 B.n197 B.n108 10.6151
R636 B.n198 B.n197 10.6151
R637 B.n199 B.n198 10.6151
R638 B.n199 B.n106 10.6151
R639 B.n203 B.n106 10.6151
R640 B.n204 B.n203 10.6151
R641 B.n205 B.n204 10.6151
R642 B.n205 B.n104 10.6151
R643 B.n209 B.n104 10.6151
R644 B.n210 B.n209 10.6151
R645 B.n212 B.n100 10.6151
R646 B.n216 B.n100 10.6151
R647 B.n217 B.n216 10.6151
R648 B.n218 B.n217 10.6151
R649 B.n218 B.n98 10.6151
R650 B.n222 B.n98 10.6151
R651 B.n223 B.n222 10.6151
R652 B.n224 B.n223 10.6151
R653 B.n228 B.n227 10.6151
R654 B.n229 B.n228 10.6151
R655 B.n229 B.n92 10.6151
R656 B.n233 B.n92 10.6151
R657 B.n234 B.n233 10.6151
R658 B.n235 B.n234 10.6151
R659 B.n235 B.n90 10.6151
R660 B.n239 B.n90 10.6151
R661 B.n240 B.n239 10.6151
R662 B.n241 B.n240 10.6151
R663 B.n241 B.n88 10.6151
R664 B.n245 B.n88 10.6151
R665 B.n246 B.n245 10.6151
R666 B.n247 B.n246 10.6151
R667 B.n247 B.n86 10.6151
R668 B.n251 B.n86 10.6151
R669 B.n252 B.n251 10.6151
R670 B.n253 B.n252 10.6151
R671 B.n253 B.n84 10.6151
R672 B.n257 B.n84 10.6151
R673 B.n258 B.n257 10.6151
R674 B.n259 B.n258 10.6151
R675 B.n259 B.n82 10.6151
R676 B.n263 B.n82 10.6151
R677 B.n173 B.n116 10.6151
R678 B.n169 B.n116 10.6151
R679 B.n169 B.n168 10.6151
R680 B.n168 B.n167 10.6151
R681 B.n167 B.n118 10.6151
R682 B.n163 B.n118 10.6151
R683 B.n163 B.n162 10.6151
R684 B.n162 B.n161 10.6151
R685 B.n161 B.n120 10.6151
R686 B.n157 B.n120 10.6151
R687 B.n157 B.n156 10.6151
R688 B.n156 B.n155 10.6151
R689 B.n155 B.n122 10.6151
R690 B.n151 B.n122 10.6151
R691 B.n151 B.n150 10.6151
R692 B.n150 B.n149 10.6151
R693 B.n149 B.n124 10.6151
R694 B.n145 B.n124 10.6151
R695 B.n145 B.n144 10.6151
R696 B.n144 B.n143 10.6151
R697 B.n143 B.n126 10.6151
R698 B.n139 B.n126 10.6151
R699 B.n139 B.n138 10.6151
R700 B.n138 B.n137 10.6151
R701 B.n137 B.n128 10.6151
R702 B.n133 B.n128 10.6151
R703 B.n133 B.n132 10.6151
R704 B.n132 B.n131 10.6151
R705 B.n131 B.n0 10.6151
R706 B.n487 B.n1 10.6151
R707 B.n487 B.n486 10.6151
R708 B.n486 B.n485 10.6151
R709 B.n485 B.n4 10.6151
R710 B.n481 B.n4 10.6151
R711 B.n481 B.n480 10.6151
R712 B.n480 B.n479 10.6151
R713 B.n479 B.n6 10.6151
R714 B.n475 B.n6 10.6151
R715 B.n475 B.n474 10.6151
R716 B.n474 B.n473 10.6151
R717 B.n473 B.n8 10.6151
R718 B.n469 B.n8 10.6151
R719 B.n469 B.n468 10.6151
R720 B.n468 B.n467 10.6151
R721 B.n467 B.n10 10.6151
R722 B.n463 B.n10 10.6151
R723 B.n463 B.n462 10.6151
R724 B.n462 B.n461 10.6151
R725 B.n461 B.n12 10.6151
R726 B.n457 B.n12 10.6151
R727 B.n457 B.n456 10.6151
R728 B.n456 B.n455 10.6151
R729 B.n455 B.n14 10.6151
R730 B.n451 B.n14 10.6151
R731 B.n451 B.n450 10.6151
R732 B.n450 B.n449 10.6151
R733 B.n449 B.n16 10.6151
R734 B.n445 B.n16 10.6151
R735 B.n407 B.n406 6.5566
R736 B.n394 B.n38 6.5566
R737 B.n212 B.n211 6.5566
R738 B.n224 B.n96 6.5566
R739 B.n408 B.n407 4.05904
R740 B.n391 B.n38 4.05904
R741 B.n211 B.n210 4.05904
R742 B.n227 B.n96 4.05904
R743 B.n491 B.n0 2.81026
R744 B.n491 B.n1 2.81026
R745 VP.n12 VP.n0 161.3
R746 VP.n11 VP.n10 161.3
R747 VP.n9 VP.n1 161.3
R748 VP.n8 VP.n7 161.3
R749 VP.n6 VP.n2 161.3
R750 VP.n3 VP.t0 105.07
R751 VP.n3 VP.t2 104.438
R752 VP.n5 VP.n4 98.6123
R753 VP.n14 VP.n13 98.6123
R754 VP.n5 VP.t3 69.524
R755 VP.n13 VP.t1 69.524
R756 VP.n4 VP.n3 46.452
R757 VP.n7 VP.n1 40.577
R758 VP.n11 VP.n1 40.577
R759 VP.n7 VP.n6 24.5923
R760 VP.n12 VP.n11 24.5923
R761 VP.n6 VP.n5 12.2964
R762 VP.n13 VP.n12 12.2964
R763 VP.n4 VP.n2 0.278335
R764 VP.n14 VP.n0 0.278335
R765 VP.n8 VP.n2 0.189894
R766 VP.n9 VP.n8 0.189894
R767 VP.n10 VP.n9 0.189894
R768 VP.n10 VP.n0 0.189894
R769 VP VP.n14 0.153485
R770 VDD1 VDD1.n1 124.391
R771 VDD1 VDD1.n0 88.3471
R772 VDD1.n0 VDD1.t1 5.19299
R773 VDD1.n0 VDD1.t0 5.19299
R774 VDD1.n1 VDD1.t2 5.19299
R775 VDD1.n1 VDD1.t3 5.19299
R776 VTAIL.n5 VTAIL.t7 76.8027
R777 VTAIL.n4 VTAIL.t1 76.8027
R778 VTAIL.n3 VTAIL.t0 76.8027
R779 VTAIL.n7 VTAIL.t2 76.8026
R780 VTAIL.n0 VTAIL.t3 76.8026
R781 VTAIL.n1 VTAIL.t6 76.8026
R782 VTAIL.n2 VTAIL.t4 76.8026
R783 VTAIL.n6 VTAIL.t5 76.8026
R784 VTAIL.n7 VTAIL.n6 19.9186
R785 VTAIL.n3 VTAIL.n2 19.9186
R786 VTAIL.n4 VTAIL.n3 2.15567
R787 VTAIL.n6 VTAIL.n5 2.15567
R788 VTAIL.n2 VTAIL.n1 2.15567
R789 VTAIL VTAIL.n0 1.13628
R790 VTAIL VTAIL.n7 1.0199
R791 VTAIL.n5 VTAIL.n4 0.470328
R792 VTAIL.n1 VTAIL.n0 0.470328
R793 VN.n0 VN.t0 105.07
R794 VN.n1 VN.t1 105.07
R795 VN.n0 VN.t2 104.438
R796 VN.n1 VN.t3 104.438
R797 VN VN.n1 46.7309
R798 VN VN.n0 5.90891
R799 VDD2.n2 VDD2.n0 123.865
R800 VDD2.n2 VDD2.n1 88.2889
R801 VDD2.n1 VDD2.t0 5.19299
R802 VDD2.n1 VDD2.t2 5.19299
R803 VDD2.n0 VDD2.t3 5.19299
R804 VDD2.n0 VDD2.t1 5.19299
R805 VDD2 VDD2.n2 0.0586897
C0 VDD1 VP 2.76581f
C1 VN VTAIL 2.73744f
C2 VN B 0.960127f
C3 B VTAIL 2.90449f
C4 VN VDD2 2.54811f
C5 VP w_n2470_n2220# 4.32154f
C6 VTAIL VDD2 3.95598f
C7 B VDD2 1.07774f
C8 VDD1 w_n2470_n2220# 1.21277f
C9 VN VP 4.81845f
C10 VTAIL VP 2.75155f
C11 VN VDD1 0.148773f
C12 B VP 1.48325f
C13 VTAIL VDD1 3.90465f
C14 VP VDD2 0.367105f
C15 B VDD1 1.03265f
C16 VN w_n2470_n2220# 4.0051f
C17 VDD1 VDD2 0.924313f
C18 VTAIL w_n2470_n2220# 2.65715f
C19 B w_n2470_n2220# 7.11486f
C20 w_n2470_n2220# VDD2 1.25927f
C21 VDD2 VSUBS 0.731528f
C22 VDD1 VSUBS 4.737888f
C23 VTAIL VSUBS 0.679472f
C24 VN VSUBS 5.05586f
C25 VP VSUBS 1.740282f
C26 B VSUBS 3.41641f
C27 w_n2470_n2220# VSUBS 68.3795f
C28 VDD2.t3 VSUBS 0.135004f
C29 VDD2.t1 VSUBS 0.135004f
C30 VDD2.n0 VSUBS 1.33716f
C31 VDD2.t0 VSUBS 0.135004f
C32 VDD2.t2 VSUBS 0.135004f
C33 VDD2.n1 VSUBS 0.901432f
C34 VDD2.n2 VSUBS 3.52599f
C35 VN.t0 VSUBS 1.83666f
C36 VN.t2 VSUBS 1.83168f
C37 VN.n0 VSUBS 1.22299f
C38 VN.t1 VSUBS 1.83666f
C39 VN.t3 VSUBS 1.83168f
C40 VN.n1 VSUBS 3.04839f
C41 VTAIL.t3 VSUBS 1.07863f
C42 VTAIL.n0 VSUBS 0.71915f
C43 VTAIL.t6 VSUBS 1.07863f
C44 VTAIL.n1 VSUBS 0.807392f
C45 VTAIL.t4 VSUBS 1.07863f
C46 VTAIL.n2 VSUBS 1.78535f
C47 VTAIL.t0 VSUBS 1.07864f
C48 VTAIL.n3 VSUBS 1.78534f
C49 VTAIL.t1 VSUBS 1.07864f
C50 VTAIL.n4 VSUBS 0.807386f
C51 VTAIL.t7 VSUBS 1.07864f
C52 VTAIL.n5 VSUBS 0.807386f
C53 VTAIL.t5 VSUBS 1.07863f
C54 VTAIL.n6 VSUBS 1.78535f
C55 VTAIL.t2 VSUBS 1.07863f
C56 VTAIL.n7 VSUBS 1.68703f
C57 VDD1.t1 VSUBS 0.137033f
C58 VDD1.t0 VSUBS 0.137033f
C59 VDD1.n0 VSUBS 0.91542f
C60 VDD1.t2 VSUBS 0.137033f
C61 VDD1.t3 VSUBS 0.137033f
C62 VDD1.n1 VSUBS 1.37813f
C63 VP.n0 VSUBS 0.060061f
C64 VP.t1 VSUBS 1.64203f
C65 VP.n1 VSUBS 0.036796f
C66 VP.n2 VSUBS 0.060061f
C67 VP.t3 VSUBS 1.64203f
C68 VP.t2 VSUBS 1.93164f
C69 VP.t0 VSUBS 1.93689f
C70 VP.n3 VSUBS 3.19089f
C71 VP.n4 VSUBS 2.14155f
C72 VP.n5 VSUBS 0.750467f
C73 VP.n6 VSUBS 0.06363f
C74 VP.n7 VSUBS 0.09007f
C75 VP.n8 VSUBS 0.045558f
C76 VP.n9 VSUBS 0.045558f
C77 VP.n10 VSUBS 0.045558f
C78 VP.n11 VSUBS 0.09007f
C79 VP.n12 VSUBS 0.06363f
C80 VP.n13 VSUBS 0.750467f
C81 VP.n14 VSUBS 0.065829f
C82 B.n0 VSUBS 0.005267f
C83 B.n1 VSUBS 0.005267f
C84 B.n2 VSUBS 0.008328f
C85 B.n3 VSUBS 0.008328f
C86 B.n4 VSUBS 0.008328f
C87 B.n5 VSUBS 0.008328f
C88 B.n6 VSUBS 0.008328f
C89 B.n7 VSUBS 0.008328f
C90 B.n8 VSUBS 0.008328f
C91 B.n9 VSUBS 0.008328f
C92 B.n10 VSUBS 0.008328f
C93 B.n11 VSUBS 0.008328f
C94 B.n12 VSUBS 0.008328f
C95 B.n13 VSUBS 0.008328f
C96 B.n14 VSUBS 0.008328f
C97 B.n15 VSUBS 0.008328f
C98 B.n16 VSUBS 0.008328f
C99 B.n17 VSUBS 0.020765f
C100 B.n18 VSUBS 0.008328f
C101 B.n19 VSUBS 0.008328f
C102 B.n20 VSUBS 0.008328f
C103 B.n21 VSUBS 0.008328f
C104 B.n22 VSUBS 0.008328f
C105 B.n23 VSUBS 0.008328f
C106 B.n24 VSUBS 0.008328f
C107 B.n25 VSUBS 0.008328f
C108 B.n26 VSUBS 0.008328f
C109 B.n27 VSUBS 0.008328f
C110 B.n28 VSUBS 0.008328f
C111 B.n29 VSUBS 0.008328f
C112 B.t2 VSUBS 0.219389f
C113 B.t1 VSUBS 0.240479f
C114 B.t0 VSUBS 0.75563f
C115 B.n30 VSUBS 0.13642f
C116 B.n31 VSUBS 0.082277f
C117 B.n32 VSUBS 0.008328f
C118 B.n33 VSUBS 0.008328f
C119 B.n34 VSUBS 0.008328f
C120 B.n35 VSUBS 0.008328f
C121 B.t5 VSUBS 0.219389f
C122 B.t4 VSUBS 0.240477f
C123 B.t3 VSUBS 0.75563f
C124 B.n36 VSUBS 0.136422f
C125 B.n37 VSUBS 0.082278f
C126 B.n38 VSUBS 0.019296f
C127 B.n39 VSUBS 0.008328f
C128 B.n40 VSUBS 0.008328f
C129 B.n41 VSUBS 0.008328f
C130 B.n42 VSUBS 0.008328f
C131 B.n43 VSUBS 0.008328f
C132 B.n44 VSUBS 0.008328f
C133 B.n45 VSUBS 0.008328f
C134 B.n46 VSUBS 0.008328f
C135 B.n47 VSUBS 0.008328f
C136 B.n48 VSUBS 0.008328f
C137 B.n49 VSUBS 0.008328f
C138 B.n50 VSUBS 0.008328f
C139 B.n51 VSUBS 0.019652f
C140 B.n52 VSUBS 0.008328f
C141 B.n53 VSUBS 0.008328f
C142 B.n54 VSUBS 0.008328f
C143 B.n55 VSUBS 0.008328f
C144 B.n56 VSUBS 0.008328f
C145 B.n57 VSUBS 0.008328f
C146 B.n58 VSUBS 0.008328f
C147 B.n59 VSUBS 0.008328f
C148 B.n60 VSUBS 0.008328f
C149 B.n61 VSUBS 0.008328f
C150 B.n62 VSUBS 0.008328f
C151 B.n63 VSUBS 0.008328f
C152 B.n64 VSUBS 0.008328f
C153 B.n65 VSUBS 0.008328f
C154 B.n66 VSUBS 0.008328f
C155 B.n67 VSUBS 0.008328f
C156 B.n68 VSUBS 0.008328f
C157 B.n69 VSUBS 0.008328f
C158 B.n70 VSUBS 0.008328f
C159 B.n71 VSUBS 0.008328f
C160 B.n72 VSUBS 0.008328f
C161 B.n73 VSUBS 0.008328f
C162 B.n74 VSUBS 0.008328f
C163 B.n75 VSUBS 0.008328f
C164 B.n76 VSUBS 0.008328f
C165 B.n77 VSUBS 0.008328f
C166 B.n78 VSUBS 0.008328f
C167 B.n79 VSUBS 0.008328f
C168 B.n80 VSUBS 0.008328f
C169 B.n81 VSUBS 0.019652f
C170 B.n82 VSUBS 0.008328f
C171 B.n83 VSUBS 0.008328f
C172 B.n84 VSUBS 0.008328f
C173 B.n85 VSUBS 0.008328f
C174 B.n86 VSUBS 0.008328f
C175 B.n87 VSUBS 0.008328f
C176 B.n88 VSUBS 0.008328f
C177 B.n89 VSUBS 0.008328f
C178 B.n90 VSUBS 0.008328f
C179 B.n91 VSUBS 0.008328f
C180 B.n92 VSUBS 0.008328f
C181 B.n93 VSUBS 0.008328f
C182 B.t7 VSUBS 0.219389f
C183 B.t8 VSUBS 0.240477f
C184 B.t6 VSUBS 0.75563f
C185 B.n94 VSUBS 0.136422f
C186 B.n95 VSUBS 0.082278f
C187 B.n96 VSUBS 0.019296f
C188 B.n97 VSUBS 0.008328f
C189 B.n98 VSUBS 0.008328f
C190 B.n99 VSUBS 0.008328f
C191 B.n100 VSUBS 0.008328f
C192 B.n101 VSUBS 0.008328f
C193 B.t10 VSUBS 0.219389f
C194 B.t11 VSUBS 0.240479f
C195 B.t9 VSUBS 0.75563f
C196 B.n102 VSUBS 0.13642f
C197 B.n103 VSUBS 0.082277f
C198 B.n104 VSUBS 0.008328f
C199 B.n105 VSUBS 0.008328f
C200 B.n106 VSUBS 0.008328f
C201 B.n107 VSUBS 0.008328f
C202 B.n108 VSUBS 0.008328f
C203 B.n109 VSUBS 0.008328f
C204 B.n110 VSUBS 0.008328f
C205 B.n111 VSUBS 0.008328f
C206 B.n112 VSUBS 0.008328f
C207 B.n113 VSUBS 0.008328f
C208 B.n114 VSUBS 0.008328f
C209 B.n115 VSUBS 0.020765f
C210 B.n116 VSUBS 0.008328f
C211 B.n117 VSUBS 0.008328f
C212 B.n118 VSUBS 0.008328f
C213 B.n119 VSUBS 0.008328f
C214 B.n120 VSUBS 0.008328f
C215 B.n121 VSUBS 0.008328f
C216 B.n122 VSUBS 0.008328f
C217 B.n123 VSUBS 0.008328f
C218 B.n124 VSUBS 0.008328f
C219 B.n125 VSUBS 0.008328f
C220 B.n126 VSUBS 0.008328f
C221 B.n127 VSUBS 0.008328f
C222 B.n128 VSUBS 0.008328f
C223 B.n129 VSUBS 0.008328f
C224 B.n130 VSUBS 0.008328f
C225 B.n131 VSUBS 0.008328f
C226 B.n132 VSUBS 0.008328f
C227 B.n133 VSUBS 0.008328f
C228 B.n134 VSUBS 0.008328f
C229 B.n135 VSUBS 0.008328f
C230 B.n136 VSUBS 0.008328f
C231 B.n137 VSUBS 0.008328f
C232 B.n138 VSUBS 0.008328f
C233 B.n139 VSUBS 0.008328f
C234 B.n140 VSUBS 0.008328f
C235 B.n141 VSUBS 0.008328f
C236 B.n142 VSUBS 0.008328f
C237 B.n143 VSUBS 0.008328f
C238 B.n144 VSUBS 0.008328f
C239 B.n145 VSUBS 0.008328f
C240 B.n146 VSUBS 0.008328f
C241 B.n147 VSUBS 0.008328f
C242 B.n148 VSUBS 0.008328f
C243 B.n149 VSUBS 0.008328f
C244 B.n150 VSUBS 0.008328f
C245 B.n151 VSUBS 0.008328f
C246 B.n152 VSUBS 0.008328f
C247 B.n153 VSUBS 0.008328f
C248 B.n154 VSUBS 0.008328f
C249 B.n155 VSUBS 0.008328f
C250 B.n156 VSUBS 0.008328f
C251 B.n157 VSUBS 0.008328f
C252 B.n158 VSUBS 0.008328f
C253 B.n159 VSUBS 0.008328f
C254 B.n160 VSUBS 0.008328f
C255 B.n161 VSUBS 0.008328f
C256 B.n162 VSUBS 0.008328f
C257 B.n163 VSUBS 0.008328f
C258 B.n164 VSUBS 0.008328f
C259 B.n165 VSUBS 0.008328f
C260 B.n166 VSUBS 0.008328f
C261 B.n167 VSUBS 0.008328f
C262 B.n168 VSUBS 0.008328f
C263 B.n169 VSUBS 0.008328f
C264 B.n170 VSUBS 0.008328f
C265 B.n171 VSUBS 0.008328f
C266 B.n172 VSUBS 0.019652f
C267 B.n173 VSUBS 0.019652f
C268 B.n174 VSUBS 0.020765f
C269 B.n175 VSUBS 0.008328f
C270 B.n176 VSUBS 0.008328f
C271 B.n177 VSUBS 0.008328f
C272 B.n178 VSUBS 0.008328f
C273 B.n179 VSUBS 0.008328f
C274 B.n180 VSUBS 0.008328f
C275 B.n181 VSUBS 0.008328f
C276 B.n182 VSUBS 0.008328f
C277 B.n183 VSUBS 0.008328f
C278 B.n184 VSUBS 0.008328f
C279 B.n185 VSUBS 0.008328f
C280 B.n186 VSUBS 0.008328f
C281 B.n187 VSUBS 0.008328f
C282 B.n188 VSUBS 0.008328f
C283 B.n189 VSUBS 0.008328f
C284 B.n190 VSUBS 0.008328f
C285 B.n191 VSUBS 0.008328f
C286 B.n192 VSUBS 0.008328f
C287 B.n193 VSUBS 0.008328f
C288 B.n194 VSUBS 0.008328f
C289 B.n195 VSUBS 0.008328f
C290 B.n196 VSUBS 0.008328f
C291 B.n197 VSUBS 0.008328f
C292 B.n198 VSUBS 0.008328f
C293 B.n199 VSUBS 0.008328f
C294 B.n200 VSUBS 0.008328f
C295 B.n201 VSUBS 0.008328f
C296 B.n202 VSUBS 0.008328f
C297 B.n203 VSUBS 0.008328f
C298 B.n204 VSUBS 0.008328f
C299 B.n205 VSUBS 0.008328f
C300 B.n206 VSUBS 0.008328f
C301 B.n207 VSUBS 0.008328f
C302 B.n208 VSUBS 0.008328f
C303 B.n209 VSUBS 0.008328f
C304 B.n210 VSUBS 0.005756f
C305 B.n211 VSUBS 0.019296f
C306 B.n212 VSUBS 0.006736f
C307 B.n213 VSUBS 0.008328f
C308 B.n214 VSUBS 0.008328f
C309 B.n215 VSUBS 0.008328f
C310 B.n216 VSUBS 0.008328f
C311 B.n217 VSUBS 0.008328f
C312 B.n218 VSUBS 0.008328f
C313 B.n219 VSUBS 0.008328f
C314 B.n220 VSUBS 0.008328f
C315 B.n221 VSUBS 0.008328f
C316 B.n222 VSUBS 0.008328f
C317 B.n223 VSUBS 0.008328f
C318 B.n224 VSUBS 0.006736f
C319 B.n225 VSUBS 0.008328f
C320 B.n226 VSUBS 0.008328f
C321 B.n227 VSUBS 0.005756f
C322 B.n228 VSUBS 0.008328f
C323 B.n229 VSUBS 0.008328f
C324 B.n230 VSUBS 0.008328f
C325 B.n231 VSUBS 0.008328f
C326 B.n232 VSUBS 0.008328f
C327 B.n233 VSUBS 0.008328f
C328 B.n234 VSUBS 0.008328f
C329 B.n235 VSUBS 0.008328f
C330 B.n236 VSUBS 0.008328f
C331 B.n237 VSUBS 0.008328f
C332 B.n238 VSUBS 0.008328f
C333 B.n239 VSUBS 0.008328f
C334 B.n240 VSUBS 0.008328f
C335 B.n241 VSUBS 0.008328f
C336 B.n242 VSUBS 0.008328f
C337 B.n243 VSUBS 0.008328f
C338 B.n244 VSUBS 0.008328f
C339 B.n245 VSUBS 0.008328f
C340 B.n246 VSUBS 0.008328f
C341 B.n247 VSUBS 0.008328f
C342 B.n248 VSUBS 0.008328f
C343 B.n249 VSUBS 0.008328f
C344 B.n250 VSUBS 0.008328f
C345 B.n251 VSUBS 0.008328f
C346 B.n252 VSUBS 0.008328f
C347 B.n253 VSUBS 0.008328f
C348 B.n254 VSUBS 0.008328f
C349 B.n255 VSUBS 0.008328f
C350 B.n256 VSUBS 0.008328f
C351 B.n257 VSUBS 0.008328f
C352 B.n258 VSUBS 0.008328f
C353 B.n259 VSUBS 0.008328f
C354 B.n260 VSUBS 0.008328f
C355 B.n261 VSUBS 0.008328f
C356 B.n262 VSUBS 0.020765f
C357 B.n263 VSUBS 0.020765f
C358 B.n264 VSUBS 0.019652f
C359 B.n265 VSUBS 0.008328f
C360 B.n266 VSUBS 0.008328f
C361 B.n267 VSUBS 0.008328f
C362 B.n268 VSUBS 0.008328f
C363 B.n269 VSUBS 0.008328f
C364 B.n270 VSUBS 0.008328f
C365 B.n271 VSUBS 0.008328f
C366 B.n272 VSUBS 0.008328f
C367 B.n273 VSUBS 0.008328f
C368 B.n274 VSUBS 0.008328f
C369 B.n275 VSUBS 0.008328f
C370 B.n276 VSUBS 0.008328f
C371 B.n277 VSUBS 0.008328f
C372 B.n278 VSUBS 0.008328f
C373 B.n279 VSUBS 0.008328f
C374 B.n280 VSUBS 0.008328f
C375 B.n281 VSUBS 0.008328f
C376 B.n282 VSUBS 0.008328f
C377 B.n283 VSUBS 0.008328f
C378 B.n284 VSUBS 0.008328f
C379 B.n285 VSUBS 0.008328f
C380 B.n286 VSUBS 0.008328f
C381 B.n287 VSUBS 0.008328f
C382 B.n288 VSUBS 0.008328f
C383 B.n289 VSUBS 0.008328f
C384 B.n290 VSUBS 0.008328f
C385 B.n291 VSUBS 0.008328f
C386 B.n292 VSUBS 0.008328f
C387 B.n293 VSUBS 0.008328f
C388 B.n294 VSUBS 0.008328f
C389 B.n295 VSUBS 0.008328f
C390 B.n296 VSUBS 0.008328f
C391 B.n297 VSUBS 0.008328f
C392 B.n298 VSUBS 0.008328f
C393 B.n299 VSUBS 0.008328f
C394 B.n300 VSUBS 0.008328f
C395 B.n301 VSUBS 0.008328f
C396 B.n302 VSUBS 0.008328f
C397 B.n303 VSUBS 0.008328f
C398 B.n304 VSUBS 0.008328f
C399 B.n305 VSUBS 0.008328f
C400 B.n306 VSUBS 0.008328f
C401 B.n307 VSUBS 0.008328f
C402 B.n308 VSUBS 0.008328f
C403 B.n309 VSUBS 0.008328f
C404 B.n310 VSUBS 0.008328f
C405 B.n311 VSUBS 0.008328f
C406 B.n312 VSUBS 0.008328f
C407 B.n313 VSUBS 0.008328f
C408 B.n314 VSUBS 0.008328f
C409 B.n315 VSUBS 0.008328f
C410 B.n316 VSUBS 0.008328f
C411 B.n317 VSUBS 0.008328f
C412 B.n318 VSUBS 0.008328f
C413 B.n319 VSUBS 0.008328f
C414 B.n320 VSUBS 0.008328f
C415 B.n321 VSUBS 0.008328f
C416 B.n322 VSUBS 0.008328f
C417 B.n323 VSUBS 0.008328f
C418 B.n324 VSUBS 0.008328f
C419 B.n325 VSUBS 0.008328f
C420 B.n326 VSUBS 0.008328f
C421 B.n327 VSUBS 0.008328f
C422 B.n328 VSUBS 0.008328f
C423 B.n329 VSUBS 0.008328f
C424 B.n330 VSUBS 0.008328f
C425 B.n331 VSUBS 0.008328f
C426 B.n332 VSUBS 0.008328f
C427 B.n333 VSUBS 0.008328f
C428 B.n334 VSUBS 0.008328f
C429 B.n335 VSUBS 0.008328f
C430 B.n336 VSUBS 0.008328f
C431 B.n337 VSUBS 0.008328f
C432 B.n338 VSUBS 0.008328f
C433 B.n339 VSUBS 0.008328f
C434 B.n340 VSUBS 0.008328f
C435 B.n341 VSUBS 0.008328f
C436 B.n342 VSUBS 0.008328f
C437 B.n343 VSUBS 0.008328f
C438 B.n344 VSUBS 0.008328f
C439 B.n345 VSUBS 0.008328f
C440 B.n346 VSUBS 0.008328f
C441 B.n347 VSUBS 0.008328f
C442 B.n348 VSUBS 0.008328f
C443 B.n349 VSUBS 0.008328f
C444 B.n350 VSUBS 0.008328f
C445 B.n351 VSUBS 0.008328f
C446 B.n352 VSUBS 0.008328f
C447 B.n353 VSUBS 0.008328f
C448 B.n354 VSUBS 0.020584f
C449 B.n355 VSUBS 0.019834f
C450 B.n356 VSUBS 0.020765f
C451 B.n357 VSUBS 0.008328f
C452 B.n358 VSUBS 0.008328f
C453 B.n359 VSUBS 0.008328f
C454 B.n360 VSUBS 0.008328f
C455 B.n361 VSUBS 0.008328f
C456 B.n362 VSUBS 0.008328f
C457 B.n363 VSUBS 0.008328f
C458 B.n364 VSUBS 0.008328f
C459 B.n365 VSUBS 0.008328f
C460 B.n366 VSUBS 0.008328f
C461 B.n367 VSUBS 0.008328f
C462 B.n368 VSUBS 0.008328f
C463 B.n369 VSUBS 0.008328f
C464 B.n370 VSUBS 0.008328f
C465 B.n371 VSUBS 0.008328f
C466 B.n372 VSUBS 0.008328f
C467 B.n373 VSUBS 0.008328f
C468 B.n374 VSUBS 0.008328f
C469 B.n375 VSUBS 0.008328f
C470 B.n376 VSUBS 0.008328f
C471 B.n377 VSUBS 0.008328f
C472 B.n378 VSUBS 0.008328f
C473 B.n379 VSUBS 0.008328f
C474 B.n380 VSUBS 0.008328f
C475 B.n381 VSUBS 0.008328f
C476 B.n382 VSUBS 0.008328f
C477 B.n383 VSUBS 0.008328f
C478 B.n384 VSUBS 0.008328f
C479 B.n385 VSUBS 0.008328f
C480 B.n386 VSUBS 0.008328f
C481 B.n387 VSUBS 0.008328f
C482 B.n388 VSUBS 0.008328f
C483 B.n389 VSUBS 0.008328f
C484 B.n390 VSUBS 0.008328f
C485 B.n391 VSUBS 0.005756f
C486 B.n392 VSUBS 0.008328f
C487 B.n393 VSUBS 0.008328f
C488 B.n394 VSUBS 0.006736f
C489 B.n395 VSUBS 0.008328f
C490 B.n396 VSUBS 0.008328f
C491 B.n397 VSUBS 0.008328f
C492 B.n398 VSUBS 0.008328f
C493 B.n399 VSUBS 0.008328f
C494 B.n400 VSUBS 0.008328f
C495 B.n401 VSUBS 0.008328f
C496 B.n402 VSUBS 0.008328f
C497 B.n403 VSUBS 0.008328f
C498 B.n404 VSUBS 0.008328f
C499 B.n405 VSUBS 0.008328f
C500 B.n406 VSUBS 0.006736f
C501 B.n407 VSUBS 0.019296f
C502 B.n408 VSUBS 0.005756f
C503 B.n409 VSUBS 0.008328f
C504 B.n410 VSUBS 0.008328f
C505 B.n411 VSUBS 0.008328f
C506 B.n412 VSUBS 0.008328f
C507 B.n413 VSUBS 0.008328f
C508 B.n414 VSUBS 0.008328f
C509 B.n415 VSUBS 0.008328f
C510 B.n416 VSUBS 0.008328f
C511 B.n417 VSUBS 0.008328f
C512 B.n418 VSUBS 0.008328f
C513 B.n419 VSUBS 0.008328f
C514 B.n420 VSUBS 0.008328f
C515 B.n421 VSUBS 0.008328f
C516 B.n422 VSUBS 0.008328f
C517 B.n423 VSUBS 0.008328f
C518 B.n424 VSUBS 0.008328f
C519 B.n425 VSUBS 0.008328f
C520 B.n426 VSUBS 0.008328f
C521 B.n427 VSUBS 0.008328f
C522 B.n428 VSUBS 0.008328f
C523 B.n429 VSUBS 0.008328f
C524 B.n430 VSUBS 0.008328f
C525 B.n431 VSUBS 0.008328f
C526 B.n432 VSUBS 0.008328f
C527 B.n433 VSUBS 0.008328f
C528 B.n434 VSUBS 0.008328f
C529 B.n435 VSUBS 0.008328f
C530 B.n436 VSUBS 0.008328f
C531 B.n437 VSUBS 0.008328f
C532 B.n438 VSUBS 0.008328f
C533 B.n439 VSUBS 0.008328f
C534 B.n440 VSUBS 0.008328f
C535 B.n441 VSUBS 0.008328f
C536 B.n442 VSUBS 0.008328f
C537 B.n443 VSUBS 0.008328f
C538 B.n444 VSUBS 0.020765f
C539 B.n445 VSUBS 0.019652f
C540 B.n446 VSUBS 0.019652f
C541 B.n447 VSUBS 0.008328f
C542 B.n448 VSUBS 0.008328f
C543 B.n449 VSUBS 0.008328f
C544 B.n450 VSUBS 0.008328f
C545 B.n451 VSUBS 0.008328f
C546 B.n452 VSUBS 0.008328f
C547 B.n453 VSUBS 0.008328f
C548 B.n454 VSUBS 0.008328f
C549 B.n455 VSUBS 0.008328f
C550 B.n456 VSUBS 0.008328f
C551 B.n457 VSUBS 0.008328f
C552 B.n458 VSUBS 0.008328f
C553 B.n459 VSUBS 0.008328f
C554 B.n460 VSUBS 0.008328f
C555 B.n461 VSUBS 0.008328f
C556 B.n462 VSUBS 0.008328f
C557 B.n463 VSUBS 0.008328f
C558 B.n464 VSUBS 0.008328f
C559 B.n465 VSUBS 0.008328f
C560 B.n466 VSUBS 0.008328f
C561 B.n467 VSUBS 0.008328f
C562 B.n468 VSUBS 0.008328f
C563 B.n469 VSUBS 0.008328f
C564 B.n470 VSUBS 0.008328f
C565 B.n471 VSUBS 0.008328f
C566 B.n472 VSUBS 0.008328f
C567 B.n473 VSUBS 0.008328f
C568 B.n474 VSUBS 0.008328f
C569 B.n475 VSUBS 0.008328f
C570 B.n476 VSUBS 0.008328f
C571 B.n477 VSUBS 0.008328f
C572 B.n478 VSUBS 0.008328f
C573 B.n479 VSUBS 0.008328f
C574 B.n480 VSUBS 0.008328f
C575 B.n481 VSUBS 0.008328f
C576 B.n482 VSUBS 0.008328f
C577 B.n483 VSUBS 0.008328f
C578 B.n484 VSUBS 0.008328f
C579 B.n485 VSUBS 0.008328f
C580 B.n486 VSUBS 0.008328f
C581 B.n487 VSUBS 0.008328f
C582 B.n488 VSUBS 0.008328f
C583 B.n489 VSUBS 0.008328f
C584 B.n490 VSUBS 0.008328f
C585 B.n491 VSUBS 0.018859f
.ends

