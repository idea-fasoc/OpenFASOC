* NGSPICE file created from diff_pair_sample_1415.ext - technology: sky130A

.subckt diff_pair_sample_1415 VTAIL VN VP B VDD2 VDD1
X0 B.t19 B.t17 B.t18 B.t7 sky130_fd_pr__nfet_01v8 ad=4.5318 pd=24.02 as=0 ps=0 w=11.62 l=1.46
X1 VTAIL.t11 VN.t0 VDD2.t0 B.t3 sky130_fd_pr__nfet_01v8 ad=1.9173 pd=11.95 as=1.9173 ps=11.95 w=11.62 l=1.46
X2 VTAIL.t1 VP.t0 VDD1.t5 B.t3 sky130_fd_pr__nfet_01v8 ad=1.9173 pd=11.95 as=1.9173 ps=11.95 w=11.62 l=1.46
X3 VDD1.t4 VP.t1 VTAIL.t5 B.t0 sky130_fd_pr__nfet_01v8 ad=4.5318 pd=24.02 as=1.9173 ps=11.95 w=11.62 l=1.46
X4 B.t16 B.t14 B.t15 B.t11 sky130_fd_pr__nfet_01v8 ad=4.5318 pd=24.02 as=0 ps=0 w=11.62 l=1.46
X5 VDD1.t3 VP.t2 VTAIL.t4 B.t1 sky130_fd_pr__nfet_01v8 ad=4.5318 pd=24.02 as=1.9173 ps=11.95 w=11.62 l=1.46
X6 VDD2.t5 VN.t1 VTAIL.t10 B.t1 sky130_fd_pr__nfet_01v8 ad=4.5318 pd=24.02 as=1.9173 ps=11.95 w=11.62 l=1.46
X7 VTAIL.t2 VP.t3 VDD1.t2 B.t4 sky130_fd_pr__nfet_01v8 ad=1.9173 pd=11.95 as=1.9173 ps=11.95 w=11.62 l=1.46
X8 B.t13 B.t10 B.t12 B.t11 sky130_fd_pr__nfet_01v8 ad=4.5318 pd=24.02 as=0 ps=0 w=11.62 l=1.46
X9 VTAIL.t9 VN.t2 VDD2.t1 B.t4 sky130_fd_pr__nfet_01v8 ad=1.9173 pd=11.95 as=1.9173 ps=11.95 w=11.62 l=1.46
X10 VDD2.t3 VN.t3 VTAIL.t8 B.t2 sky130_fd_pr__nfet_01v8 ad=1.9173 pd=11.95 as=4.5318 ps=24.02 w=11.62 l=1.46
X11 VDD2.t2 VN.t4 VTAIL.t7 B.t0 sky130_fd_pr__nfet_01v8 ad=4.5318 pd=24.02 as=1.9173 ps=11.95 w=11.62 l=1.46
X12 B.t9 B.t6 B.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=4.5318 pd=24.02 as=0 ps=0 w=11.62 l=1.46
X13 VDD1.t1 VP.t4 VTAIL.t3 B.t5 sky130_fd_pr__nfet_01v8 ad=1.9173 pd=11.95 as=4.5318 ps=24.02 w=11.62 l=1.46
X14 VDD2.t4 VN.t5 VTAIL.t6 B.t5 sky130_fd_pr__nfet_01v8 ad=1.9173 pd=11.95 as=4.5318 ps=24.02 w=11.62 l=1.46
X15 VDD1.t0 VP.t5 VTAIL.t0 B.t2 sky130_fd_pr__nfet_01v8 ad=1.9173 pd=11.95 as=4.5318 ps=24.02 w=11.62 l=1.46
R0 B.n701 B.n700 585
R1 B.n702 B.n701 585
R2 B.n286 B.n101 585
R3 B.n285 B.n284 585
R4 B.n283 B.n282 585
R5 B.n281 B.n280 585
R6 B.n279 B.n278 585
R7 B.n277 B.n276 585
R8 B.n275 B.n274 585
R9 B.n273 B.n272 585
R10 B.n271 B.n270 585
R11 B.n269 B.n268 585
R12 B.n267 B.n266 585
R13 B.n265 B.n264 585
R14 B.n263 B.n262 585
R15 B.n261 B.n260 585
R16 B.n259 B.n258 585
R17 B.n257 B.n256 585
R18 B.n255 B.n254 585
R19 B.n253 B.n252 585
R20 B.n251 B.n250 585
R21 B.n249 B.n248 585
R22 B.n247 B.n246 585
R23 B.n245 B.n244 585
R24 B.n243 B.n242 585
R25 B.n241 B.n240 585
R26 B.n239 B.n238 585
R27 B.n237 B.n236 585
R28 B.n235 B.n234 585
R29 B.n233 B.n232 585
R30 B.n231 B.n230 585
R31 B.n229 B.n228 585
R32 B.n227 B.n226 585
R33 B.n225 B.n224 585
R34 B.n223 B.n222 585
R35 B.n221 B.n220 585
R36 B.n219 B.n218 585
R37 B.n217 B.n216 585
R38 B.n215 B.n214 585
R39 B.n213 B.n212 585
R40 B.n211 B.n210 585
R41 B.n209 B.n208 585
R42 B.n207 B.n206 585
R43 B.n205 B.n204 585
R44 B.n203 B.n202 585
R45 B.n201 B.n200 585
R46 B.n199 B.n198 585
R47 B.n197 B.n196 585
R48 B.n195 B.n194 585
R49 B.n193 B.n192 585
R50 B.n191 B.n190 585
R51 B.n188 B.n187 585
R52 B.n186 B.n185 585
R53 B.n184 B.n183 585
R54 B.n182 B.n181 585
R55 B.n180 B.n179 585
R56 B.n178 B.n177 585
R57 B.n176 B.n175 585
R58 B.n174 B.n173 585
R59 B.n172 B.n171 585
R60 B.n170 B.n169 585
R61 B.n168 B.n167 585
R62 B.n166 B.n165 585
R63 B.n164 B.n163 585
R64 B.n162 B.n161 585
R65 B.n160 B.n159 585
R66 B.n158 B.n157 585
R67 B.n156 B.n155 585
R68 B.n154 B.n153 585
R69 B.n152 B.n151 585
R70 B.n150 B.n149 585
R71 B.n148 B.n147 585
R72 B.n146 B.n145 585
R73 B.n144 B.n143 585
R74 B.n142 B.n141 585
R75 B.n140 B.n139 585
R76 B.n138 B.n137 585
R77 B.n136 B.n135 585
R78 B.n134 B.n133 585
R79 B.n132 B.n131 585
R80 B.n130 B.n129 585
R81 B.n128 B.n127 585
R82 B.n126 B.n125 585
R83 B.n124 B.n123 585
R84 B.n122 B.n121 585
R85 B.n120 B.n119 585
R86 B.n118 B.n117 585
R87 B.n116 B.n115 585
R88 B.n114 B.n113 585
R89 B.n112 B.n111 585
R90 B.n110 B.n109 585
R91 B.n108 B.n107 585
R92 B.n699 B.n55 585
R93 B.n703 B.n55 585
R94 B.n698 B.n54 585
R95 B.n704 B.n54 585
R96 B.n697 B.n696 585
R97 B.n696 B.n50 585
R98 B.n695 B.n49 585
R99 B.n710 B.n49 585
R100 B.n694 B.n48 585
R101 B.n711 B.n48 585
R102 B.n693 B.n47 585
R103 B.n712 B.n47 585
R104 B.n692 B.n691 585
R105 B.n691 B.n43 585
R106 B.n690 B.n42 585
R107 B.n718 B.n42 585
R108 B.n689 B.n41 585
R109 B.n719 B.n41 585
R110 B.n688 B.n40 585
R111 B.n720 B.n40 585
R112 B.n687 B.n686 585
R113 B.n686 B.n36 585
R114 B.n685 B.n35 585
R115 B.n726 B.n35 585
R116 B.n684 B.n34 585
R117 B.n727 B.n34 585
R118 B.n683 B.n33 585
R119 B.n728 B.n33 585
R120 B.n682 B.n681 585
R121 B.n681 B.n32 585
R122 B.n680 B.n28 585
R123 B.n734 B.n28 585
R124 B.n679 B.n27 585
R125 B.n735 B.n27 585
R126 B.n678 B.n26 585
R127 B.n736 B.n26 585
R128 B.n677 B.n676 585
R129 B.n676 B.n22 585
R130 B.n675 B.n21 585
R131 B.n742 B.n21 585
R132 B.n674 B.n20 585
R133 B.n743 B.n20 585
R134 B.n673 B.n19 585
R135 B.n744 B.n19 585
R136 B.n672 B.n671 585
R137 B.n671 B.n15 585
R138 B.n670 B.n14 585
R139 B.n750 B.n14 585
R140 B.n669 B.n13 585
R141 B.n751 B.n13 585
R142 B.n668 B.n12 585
R143 B.n752 B.n12 585
R144 B.n667 B.n666 585
R145 B.n666 B.n8 585
R146 B.n665 B.n7 585
R147 B.n758 B.n7 585
R148 B.n664 B.n6 585
R149 B.n759 B.n6 585
R150 B.n663 B.n5 585
R151 B.n760 B.n5 585
R152 B.n662 B.n661 585
R153 B.n661 B.n4 585
R154 B.n660 B.n287 585
R155 B.n660 B.n659 585
R156 B.n650 B.n288 585
R157 B.n289 B.n288 585
R158 B.n652 B.n651 585
R159 B.n653 B.n652 585
R160 B.n649 B.n293 585
R161 B.n297 B.n293 585
R162 B.n648 B.n647 585
R163 B.n647 B.n646 585
R164 B.n295 B.n294 585
R165 B.n296 B.n295 585
R166 B.n639 B.n638 585
R167 B.n640 B.n639 585
R168 B.n637 B.n302 585
R169 B.n302 B.n301 585
R170 B.n636 B.n635 585
R171 B.n635 B.n634 585
R172 B.n304 B.n303 585
R173 B.n305 B.n304 585
R174 B.n627 B.n626 585
R175 B.n628 B.n627 585
R176 B.n625 B.n310 585
R177 B.n310 B.n309 585
R178 B.n624 B.n623 585
R179 B.n623 B.n622 585
R180 B.n312 B.n311 585
R181 B.n615 B.n312 585
R182 B.n614 B.n613 585
R183 B.n616 B.n614 585
R184 B.n612 B.n317 585
R185 B.n317 B.n316 585
R186 B.n611 B.n610 585
R187 B.n610 B.n609 585
R188 B.n319 B.n318 585
R189 B.n320 B.n319 585
R190 B.n602 B.n601 585
R191 B.n603 B.n602 585
R192 B.n600 B.n325 585
R193 B.n325 B.n324 585
R194 B.n599 B.n598 585
R195 B.n598 B.n597 585
R196 B.n327 B.n326 585
R197 B.n328 B.n327 585
R198 B.n590 B.n589 585
R199 B.n591 B.n590 585
R200 B.n588 B.n333 585
R201 B.n333 B.n332 585
R202 B.n587 B.n586 585
R203 B.n586 B.n585 585
R204 B.n335 B.n334 585
R205 B.n336 B.n335 585
R206 B.n578 B.n577 585
R207 B.n579 B.n578 585
R208 B.n576 B.n341 585
R209 B.n341 B.n340 585
R210 B.n570 B.n569 585
R211 B.n568 B.n388 585
R212 B.n567 B.n387 585
R213 B.n572 B.n387 585
R214 B.n566 B.n565 585
R215 B.n564 B.n563 585
R216 B.n562 B.n561 585
R217 B.n560 B.n559 585
R218 B.n558 B.n557 585
R219 B.n556 B.n555 585
R220 B.n554 B.n553 585
R221 B.n552 B.n551 585
R222 B.n550 B.n549 585
R223 B.n548 B.n547 585
R224 B.n546 B.n545 585
R225 B.n544 B.n543 585
R226 B.n542 B.n541 585
R227 B.n540 B.n539 585
R228 B.n538 B.n537 585
R229 B.n536 B.n535 585
R230 B.n534 B.n533 585
R231 B.n532 B.n531 585
R232 B.n530 B.n529 585
R233 B.n528 B.n527 585
R234 B.n526 B.n525 585
R235 B.n524 B.n523 585
R236 B.n522 B.n521 585
R237 B.n520 B.n519 585
R238 B.n518 B.n517 585
R239 B.n516 B.n515 585
R240 B.n514 B.n513 585
R241 B.n512 B.n511 585
R242 B.n510 B.n509 585
R243 B.n508 B.n507 585
R244 B.n506 B.n505 585
R245 B.n504 B.n503 585
R246 B.n502 B.n501 585
R247 B.n500 B.n499 585
R248 B.n498 B.n497 585
R249 B.n496 B.n495 585
R250 B.n494 B.n493 585
R251 B.n492 B.n491 585
R252 B.n490 B.n489 585
R253 B.n488 B.n487 585
R254 B.n486 B.n485 585
R255 B.n484 B.n483 585
R256 B.n482 B.n481 585
R257 B.n480 B.n479 585
R258 B.n478 B.n477 585
R259 B.n476 B.n475 585
R260 B.n474 B.n473 585
R261 B.n471 B.n470 585
R262 B.n469 B.n468 585
R263 B.n467 B.n466 585
R264 B.n465 B.n464 585
R265 B.n463 B.n462 585
R266 B.n461 B.n460 585
R267 B.n459 B.n458 585
R268 B.n457 B.n456 585
R269 B.n455 B.n454 585
R270 B.n453 B.n452 585
R271 B.n451 B.n450 585
R272 B.n449 B.n448 585
R273 B.n447 B.n446 585
R274 B.n445 B.n444 585
R275 B.n443 B.n442 585
R276 B.n441 B.n440 585
R277 B.n439 B.n438 585
R278 B.n437 B.n436 585
R279 B.n435 B.n434 585
R280 B.n433 B.n432 585
R281 B.n431 B.n430 585
R282 B.n429 B.n428 585
R283 B.n427 B.n426 585
R284 B.n425 B.n424 585
R285 B.n423 B.n422 585
R286 B.n421 B.n420 585
R287 B.n419 B.n418 585
R288 B.n417 B.n416 585
R289 B.n415 B.n414 585
R290 B.n413 B.n412 585
R291 B.n411 B.n410 585
R292 B.n409 B.n408 585
R293 B.n407 B.n406 585
R294 B.n405 B.n404 585
R295 B.n403 B.n402 585
R296 B.n401 B.n400 585
R297 B.n399 B.n398 585
R298 B.n397 B.n396 585
R299 B.n395 B.n394 585
R300 B.n343 B.n342 585
R301 B.n575 B.n574 585
R302 B.n339 B.n338 585
R303 B.n340 B.n339 585
R304 B.n581 B.n580 585
R305 B.n580 B.n579 585
R306 B.n582 B.n337 585
R307 B.n337 B.n336 585
R308 B.n584 B.n583 585
R309 B.n585 B.n584 585
R310 B.n331 B.n330 585
R311 B.n332 B.n331 585
R312 B.n593 B.n592 585
R313 B.n592 B.n591 585
R314 B.n594 B.n329 585
R315 B.n329 B.n328 585
R316 B.n596 B.n595 585
R317 B.n597 B.n596 585
R318 B.n323 B.n322 585
R319 B.n324 B.n323 585
R320 B.n605 B.n604 585
R321 B.n604 B.n603 585
R322 B.n606 B.n321 585
R323 B.n321 B.n320 585
R324 B.n608 B.n607 585
R325 B.n609 B.n608 585
R326 B.n315 B.n314 585
R327 B.n316 B.n315 585
R328 B.n618 B.n617 585
R329 B.n617 B.n616 585
R330 B.n619 B.n313 585
R331 B.n615 B.n313 585
R332 B.n621 B.n620 585
R333 B.n622 B.n621 585
R334 B.n308 B.n307 585
R335 B.n309 B.n308 585
R336 B.n630 B.n629 585
R337 B.n629 B.n628 585
R338 B.n631 B.n306 585
R339 B.n306 B.n305 585
R340 B.n633 B.n632 585
R341 B.n634 B.n633 585
R342 B.n300 B.n299 585
R343 B.n301 B.n300 585
R344 B.n642 B.n641 585
R345 B.n641 B.n640 585
R346 B.n643 B.n298 585
R347 B.n298 B.n296 585
R348 B.n645 B.n644 585
R349 B.n646 B.n645 585
R350 B.n292 B.n291 585
R351 B.n297 B.n292 585
R352 B.n655 B.n654 585
R353 B.n654 B.n653 585
R354 B.n656 B.n290 585
R355 B.n290 B.n289 585
R356 B.n658 B.n657 585
R357 B.n659 B.n658 585
R358 B.n2 B.n0 585
R359 B.n4 B.n2 585
R360 B.n3 B.n1 585
R361 B.n759 B.n3 585
R362 B.n757 B.n756 585
R363 B.n758 B.n757 585
R364 B.n755 B.n9 585
R365 B.n9 B.n8 585
R366 B.n754 B.n753 585
R367 B.n753 B.n752 585
R368 B.n11 B.n10 585
R369 B.n751 B.n11 585
R370 B.n749 B.n748 585
R371 B.n750 B.n749 585
R372 B.n747 B.n16 585
R373 B.n16 B.n15 585
R374 B.n746 B.n745 585
R375 B.n745 B.n744 585
R376 B.n18 B.n17 585
R377 B.n743 B.n18 585
R378 B.n741 B.n740 585
R379 B.n742 B.n741 585
R380 B.n739 B.n23 585
R381 B.n23 B.n22 585
R382 B.n738 B.n737 585
R383 B.n737 B.n736 585
R384 B.n25 B.n24 585
R385 B.n735 B.n25 585
R386 B.n733 B.n732 585
R387 B.n734 B.n733 585
R388 B.n731 B.n29 585
R389 B.n32 B.n29 585
R390 B.n730 B.n729 585
R391 B.n729 B.n728 585
R392 B.n31 B.n30 585
R393 B.n727 B.n31 585
R394 B.n725 B.n724 585
R395 B.n726 B.n725 585
R396 B.n723 B.n37 585
R397 B.n37 B.n36 585
R398 B.n722 B.n721 585
R399 B.n721 B.n720 585
R400 B.n39 B.n38 585
R401 B.n719 B.n39 585
R402 B.n717 B.n716 585
R403 B.n718 B.n717 585
R404 B.n715 B.n44 585
R405 B.n44 B.n43 585
R406 B.n714 B.n713 585
R407 B.n713 B.n712 585
R408 B.n46 B.n45 585
R409 B.n711 B.n46 585
R410 B.n709 B.n708 585
R411 B.n710 B.n709 585
R412 B.n707 B.n51 585
R413 B.n51 B.n50 585
R414 B.n706 B.n705 585
R415 B.n705 B.n704 585
R416 B.n53 B.n52 585
R417 B.n703 B.n53 585
R418 B.n762 B.n761 585
R419 B.n761 B.n760 585
R420 B.n570 B.n339 492.5
R421 B.n107 B.n53 492.5
R422 B.n574 B.n341 492.5
R423 B.n701 B.n55 492.5
R424 B.n392 B.t14 397.098
R425 B.n389 B.t10 397.098
R426 B.n105 B.t6 397.098
R427 B.n102 B.t17 397.098
R428 B.n702 B.n100 256.663
R429 B.n702 B.n99 256.663
R430 B.n702 B.n98 256.663
R431 B.n702 B.n97 256.663
R432 B.n702 B.n96 256.663
R433 B.n702 B.n95 256.663
R434 B.n702 B.n94 256.663
R435 B.n702 B.n93 256.663
R436 B.n702 B.n92 256.663
R437 B.n702 B.n91 256.663
R438 B.n702 B.n90 256.663
R439 B.n702 B.n89 256.663
R440 B.n702 B.n88 256.663
R441 B.n702 B.n87 256.663
R442 B.n702 B.n86 256.663
R443 B.n702 B.n85 256.663
R444 B.n702 B.n84 256.663
R445 B.n702 B.n83 256.663
R446 B.n702 B.n82 256.663
R447 B.n702 B.n81 256.663
R448 B.n702 B.n80 256.663
R449 B.n702 B.n79 256.663
R450 B.n702 B.n78 256.663
R451 B.n702 B.n77 256.663
R452 B.n702 B.n76 256.663
R453 B.n702 B.n75 256.663
R454 B.n702 B.n74 256.663
R455 B.n702 B.n73 256.663
R456 B.n702 B.n72 256.663
R457 B.n702 B.n71 256.663
R458 B.n702 B.n70 256.663
R459 B.n702 B.n69 256.663
R460 B.n702 B.n68 256.663
R461 B.n702 B.n67 256.663
R462 B.n702 B.n66 256.663
R463 B.n702 B.n65 256.663
R464 B.n702 B.n64 256.663
R465 B.n702 B.n63 256.663
R466 B.n702 B.n62 256.663
R467 B.n702 B.n61 256.663
R468 B.n702 B.n60 256.663
R469 B.n702 B.n59 256.663
R470 B.n702 B.n58 256.663
R471 B.n702 B.n57 256.663
R472 B.n702 B.n56 256.663
R473 B.n572 B.n571 256.663
R474 B.n572 B.n344 256.663
R475 B.n572 B.n345 256.663
R476 B.n572 B.n346 256.663
R477 B.n572 B.n347 256.663
R478 B.n572 B.n348 256.663
R479 B.n572 B.n349 256.663
R480 B.n572 B.n350 256.663
R481 B.n572 B.n351 256.663
R482 B.n572 B.n352 256.663
R483 B.n572 B.n353 256.663
R484 B.n572 B.n354 256.663
R485 B.n572 B.n355 256.663
R486 B.n572 B.n356 256.663
R487 B.n572 B.n357 256.663
R488 B.n572 B.n358 256.663
R489 B.n572 B.n359 256.663
R490 B.n572 B.n360 256.663
R491 B.n572 B.n361 256.663
R492 B.n572 B.n362 256.663
R493 B.n572 B.n363 256.663
R494 B.n572 B.n364 256.663
R495 B.n572 B.n365 256.663
R496 B.n572 B.n366 256.663
R497 B.n572 B.n367 256.663
R498 B.n572 B.n368 256.663
R499 B.n572 B.n369 256.663
R500 B.n572 B.n370 256.663
R501 B.n572 B.n371 256.663
R502 B.n572 B.n372 256.663
R503 B.n572 B.n373 256.663
R504 B.n572 B.n374 256.663
R505 B.n572 B.n375 256.663
R506 B.n572 B.n376 256.663
R507 B.n572 B.n377 256.663
R508 B.n572 B.n378 256.663
R509 B.n572 B.n379 256.663
R510 B.n572 B.n380 256.663
R511 B.n572 B.n381 256.663
R512 B.n572 B.n382 256.663
R513 B.n572 B.n383 256.663
R514 B.n572 B.n384 256.663
R515 B.n572 B.n385 256.663
R516 B.n572 B.n386 256.663
R517 B.n573 B.n572 256.663
R518 B.n580 B.n339 163.367
R519 B.n580 B.n337 163.367
R520 B.n584 B.n337 163.367
R521 B.n584 B.n331 163.367
R522 B.n592 B.n331 163.367
R523 B.n592 B.n329 163.367
R524 B.n596 B.n329 163.367
R525 B.n596 B.n323 163.367
R526 B.n604 B.n323 163.367
R527 B.n604 B.n321 163.367
R528 B.n608 B.n321 163.367
R529 B.n608 B.n315 163.367
R530 B.n617 B.n315 163.367
R531 B.n617 B.n313 163.367
R532 B.n621 B.n313 163.367
R533 B.n621 B.n308 163.367
R534 B.n629 B.n308 163.367
R535 B.n629 B.n306 163.367
R536 B.n633 B.n306 163.367
R537 B.n633 B.n300 163.367
R538 B.n641 B.n300 163.367
R539 B.n641 B.n298 163.367
R540 B.n645 B.n298 163.367
R541 B.n645 B.n292 163.367
R542 B.n654 B.n292 163.367
R543 B.n654 B.n290 163.367
R544 B.n658 B.n290 163.367
R545 B.n658 B.n2 163.367
R546 B.n761 B.n2 163.367
R547 B.n761 B.n3 163.367
R548 B.n757 B.n3 163.367
R549 B.n757 B.n9 163.367
R550 B.n753 B.n9 163.367
R551 B.n753 B.n11 163.367
R552 B.n749 B.n11 163.367
R553 B.n749 B.n16 163.367
R554 B.n745 B.n16 163.367
R555 B.n745 B.n18 163.367
R556 B.n741 B.n18 163.367
R557 B.n741 B.n23 163.367
R558 B.n737 B.n23 163.367
R559 B.n737 B.n25 163.367
R560 B.n733 B.n25 163.367
R561 B.n733 B.n29 163.367
R562 B.n729 B.n29 163.367
R563 B.n729 B.n31 163.367
R564 B.n725 B.n31 163.367
R565 B.n725 B.n37 163.367
R566 B.n721 B.n37 163.367
R567 B.n721 B.n39 163.367
R568 B.n717 B.n39 163.367
R569 B.n717 B.n44 163.367
R570 B.n713 B.n44 163.367
R571 B.n713 B.n46 163.367
R572 B.n709 B.n46 163.367
R573 B.n709 B.n51 163.367
R574 B.n705 B.n51 163.367
R575 B.n705 B.n53 163.367
R576 B.n388 B.n387 163.367
R577 B.n565 B.n387 163.367
R578 B.n563 B.n562 163.367
R579 B.n559 B.n558 163.367
R580 B.n555 B.n554 163.367
R581 B.n551 B.n550 163.367
R582 B.n547 B.n546 163.367
R583 B.n543 B.n542 163.367
R584 B.n539 B.n538 163.367
R585 B.n535 B.n534 163.367
R586 B.n531 B.n530 163.367
R587 B.n527 B.n526 163.367
R588 B.n523 B.n522 163.367
R589 B.n519 B.n518 163.367
R590 B.n515 B.n514 163.367
R591 B.n511 B.n510 163.367
R592 B.n507 B.n506 163.367
R593 B.n503 B.n502 163.367
R594 B.n499 B.n498 163.367
R595 B.n495 B.n494 163.367
R596 B.n491 B.n490 163.367
R597 B.n487 B.n486 163.367
R598 B.n483 B.n482 163.367
R599 B.n479 B.n478 163.367
R600 B.n475 B.n474 163.367
R601 B.n470 B.n469 163.367
R602 B.n466 B.n465 163.367
R603 B.n462 B.n461 163.367
R604 B.n458 B.n457 163.367
R605 B.n454 B.n453 163.367
R606 B.n450 B.n449 163.367
R607 B.n446 B.n445 163.367
R608 B.n442 B.n441 163.367
R609 B.n438 B.n437 163.367
R610 B.n434 B.n433 163.367
R611 B.n430 B.n429 163.367
R612 B.n426 B.n425 163.367
R613 B.n422 B.n421 163.367
R614 B.n418 B.n417 163.367
R615 B.n414 B.n413 163.367
R616 B.n410 B.n409 163.367
R617 B.n406 B.n405 163.367
R618 B.n402 B.n401 163.367
R619 B.n398 B.n397 163.367
R620 B.n394 B.n343 163.367
R621 B.n578 B.n341 163.367
R622 B.n578 B.n335 163.367
R623 B.n586 B.n335 163.367
R624 B.n586 B.n333 163.367
R625 B.n590 B.n333 163.367
R626 B.n590 B.n327 163.367
R627 B.n598 B.n327 163.367
R628 B.n598 B.n325 163.367
R629 B.n602 B.n325 163.367
R630 B.n602 B.n319 163.367
R631 B.n610 B.n319 163.367
R632 B.n610 B.n317 163.367
R633 B.n614 B.n317 163.367
R634 B.n614 B.n312 163.367
R635 B.n623 B.n312 163.367
R636 B.n623 B.n310 163.367
R637 B.n627 B.n310 163.367
R638 B.n627 B.n304 163.367
R639 B.n635 B.n304 163.367
R640 B.n635 B.n302 163.367
R641 B.n639 B.n302 163.367
R642 B.n639 B.n295 163.367
R643 B.n647 B.n295 163.367
R644 B.n647 B.n293 163.367
R645 B.n652 B.n293 163.367
R646 B.n652 B.n288 163.367
R647 B.n660 B.n288 163.367
R648 B.n661 B.n660 163.367
R649 B.n661 B.n5 163.367
R650 B.n6 B.n5 163.367
R651 B.n7 B.n6 163.367
R652 B.n666 B.n7 163.367
R653 B.n666 B.n12 163.367
R654 B.n13 B.n12 163.367
R655 B.n14 B.n13 163.367
R656 B.n671 B.n14 163.367
R657 B.n671 B.n19 163.367
R658 B.n20 B.n19 163.367
R659 B.n21 B.n20 163.367
R660 B.n676 B.n21 163.367
R661 B.n676 B.n26 163.367
R662 B.n27 B.n26 163.367
R663 B.n28 B.n27 163.367
R664 B.n681 B.n28 163.367
R665 B.n681 B.n33 163.367
R666 B.n34 B.n33 163.367
R667 B.n35 B.n34 163.367
R668 B.n686 B.n35 163.367
R669 B.n686 B.n40 163.367
R670 B.n41 B.n40 163.367
R671 B.n42 B.n41 163.367
R672 B.n691 B.n42 163.367
R673 B.n691 B.n47 163.367
R674 B.n48 B.n47 163.367
R675 B.n49 B.n48 163.367
R676 B.n696 B.n49 163.367
R677 B.n696 B.n54 163.367
R678 B.n55 B.n54 163.367
R679 B.n111 B.n110 163.367
R680 B.n115 B.n114 163.367
R681 B.n119 B.n118 163.367
R682 B.n123 B.n122 163.367
R683 B.n127 B.n126 163.367
R684 B.n131 B.n130 163.367
R685 B.n135 B.n134 163.367
R686 B.n139 B.n138 163.367
R687 B.n143 B.n142 163.367
R688 B.n147 B.n146 163.367
R689 B.n151 B.n150 163.367
R690 B.n155 B.n154 163.367
R691 B.n159 B.n158 163.367
R692 B.n163 B.n162 163.367
R693 B.n167 B.n166 163.367
R694 B.n171 B.n170 163.367
R695 B.n175 B.n174 163.367
R696 B.n179 B.n178 163.367
R697 B.n183 B.n182 163.367
R698 B.n187 B.n186 163.367
R699 B.n192 B.n191 163.367
R700 B.n196 B.n195 163.367
R701 B.n200 B.n199 163.367
R702 B.n204 B.n203 163.367
R703 B.n208 B.n207 163.367
R704 B.n212 B.n211 163.367
R705 B.n216 B.n215 163.367
R706 B.n220 B.n219 163.367
R707 B.n224 B.n223 163.367
R708 B.n228 B.n227 163.367
R709 B.n232 B.n231 163.367
R710 B.n236 B.n235 163.367
R711 B.n240 B.n239 163.367
R712 B.n244 B.n243 163.367
R713 B.n248 B.n247 163.367
R714 B.n252 B.n251 163.367
R715 B.n256 B.n255 163.367
R716 B.n260 B.n259 163.367
R717 B.n264 B.n263 163.367
R718 B.n268 B.n267 163.367
R719 B.n272 B.n271 163.367
R720 B.n276 B.n275 163.367
R721 B.n280 B.n279 163.367
R722 B.n284 B.n283 163.367
R723 B.n701 B.n101 163.367
R724 B.n392 B.t16 103.722
R725 B.n102 B.t18 103.722
R726 B.n389 B.t13 103.707
R727 B.n105 B.t8 103.707
R728 B.n572 B.n340 87.8963
R729 B.n703 B.n702 87.8963
R730 B.n571 B.n570 71.676
R731 B.n565 B.n344 71.676
R732 B.n562 B.n345 71.676
R733 B.n558 B.n346 71.676
R734 B.n554 B.n347 71.676
R735 B.n550 B.n348 71.676
R736 B.n546 B.n349 71.676
R737 B.n542 B.n350 71.676
R738 B.n538 B.n351 71.676
R739 B.n534 B.n352 71.676
R740 B.n530 B.n353 71.676
R741 B.n526 B.n354 71.676
R742 B.n522 B.n355 71.676
R743 B.n518 B.n356 71.676
R744 B.n514 B.n357 71.676
R745 B.n510 B.n358 71.676
R746 B.n506 B.n359 71.676
R747 B.n502 B.n360 71.676
R748 B.n498 B.n361 71.676
R749 B.n494 B.n362 71.676
R750 B.n490 B.n363 71.676
R751 B.n486 B.n364 71.676
R752 B.n482 B.n365 71.676
R753 B.n478 B.n366 71.676
R754 B.n474 B.n367 71.676
R755 B.n469 B.n368 71.676
R756 B.n465 B.n369 71.676
R757 B.n461 B.n370 71.676
R758 B.n457 B.n371 71.676
R759 B.n453 B.n372 71.676
R760 B.n449 B.n373 71.676
R761 B.n445 B.n374 71.676
R762 B.n441 B.n375 71.676
R763 B.n437 B.n376 71.676
R764 B.n433 B.n377 71.676
R765 B.n429 B.n378 71.676
R766 B.n425 B.n379 71.676
R767 B.n421 B.n380 71.676
R768 B.n417 B.n381 71.676
R769 B.n413 B.n382 71.676
R770 B.n409 B.n383 71.676
R771 B.n405 B.n384 71.676
R772 B.n401 B.n385 71.676
R773 B.n397 B.n386 71.676
R774 B.n573 B.n343 71.676
R775 B.n107 B.n56 71.676
R776 B.n111 B.n57 71.676
R777 B.n115 B.n58 71.676
R778 B.n119 B.n59 71.676
R779 B.n123 B.n60 71.676
R780 B.n127 B.n61 71.676
R781 B.n131 B.n62 71.676
R782 B.n135 B.n63 71.676
R783 B.n139 B.n64 71.676
R784 B.n143 B.n65 71.676
R785 B.n147 B.n66 71.676
R786 B.n151 B.n67 71.676
R787 B.n155 B.n68 71.676
R788 B.n159 B.n69 71.676
R789 B.n163 B.n70 71.676
R790 B.n167 B.n71 71.676
R791 B.n171 B.n72 71.676
R792 B.n175 B.n73 71.676
R793 B.n179 B.n74 71.676
R794 B.n183 B.n75 71.676
R795 B.n187 B.n76 71.676
R796 B.n192 B.n77 71.676
R797 B.n196 B.n78 71.676
R798 B.n200 B.n79 71.676
R799 B.n204 B.n80 71.676
R800 B.n208 B.n81 71.676
R801 B.n212 B.n82 71.676
R802 B.n216 B.n83 71.676
R803 B.n220 B.n84 71.676
R804 B.n224 B.n85 71.676
R805 B.n228 B.n86 71.676
R806 B.n232 B.n87 71.676
R807 B.n236 B.n88 71.676
R808 B.n240 B.n89 71.676
R809 B.n244 B.n90 71.676
R810 B.n248 B.n91 71.676
R811 B.n252 B.n92 71.676
R812 B.n256 B.n93 71.676
R813 B.n260 B.n94 71.676
R814 B.n264 B.n95 71.676
R815 B.n268 B.n96 71.676
R816 B.n272 B.n97 71.676
R817 B.n276 B.n98 71.676
R818 B.n280 B.n99 71.676
R819 B.n284 B.n100 71.676
R820 B.n101 B.n100 71.676
R821 B.n283 B.n99 71.676
R822 B.n279 B.n98 71.676
R823 B.n275 B.n97 71.676
R824 B.n271 B.n96 71.676
R825 B.n267 B.n95 71.676
R826 B.n263 B.n94 71.676
R827 B.n259 B.n93 71.676
R828 B.n255 B.n92 71.676
R829 B.n251 B.n91 71.676
R830 B.n247 B.n90 71.676
R831 B.n243 B.n89 71.676
R832 B.n239 B.n88 71.676
R833 B.n235 B.n87 71.676
R834 B.n231 B.n86 71.676
R835 B.n227 B.n85 71.676
R836 B.n223 B.n84 71.676
R837 B.n219 B.n83 71.676
R838 B.n215 B.n82 71.676
R839 B.n211 B.n81 71.676
R840 B.n207 B.n80 71.676
R841 B.n203 B.n79 71.676
R842 B.n199 B.n78 71.676
R843 B.n195 B.n77 71.676
R844 B.n191 B.n76 71.676
R845 B.n186 B.n75 71.676
R846 B.n182 B.n74 71.676
R847 B.n178 B.n73 71.676
R848 B.n174 B.n72 71.676
R849 B.n170 B.n71 71.676
R850 B.n166 B.n70 71.676
R851 B.n162 B.n69 71.676
R852 B.n158 B.n68 71.676
R853 B.n154 B.n67 71.676
R854 B.n150 B.n66 71.676
R855 B.n146 B.n65 71.676
R856 B.n142 B.n64 71.676
R857 B.n138 B.n63 71.676
R858 B.n134 B.n62 71.676
R859 B.n130 B.n61 71.676
R860 B.n126 B.n60 71.676
R861 B.n122 B.n59 71.676
R862 B.n118 B.n58 71.676
R863 B.n114 B.n57 71.676
R864 B.n110 B.n56 71.676
R865 B.n571 B.n388 71.676
R866 B.n563 B.n344 71.676
R867 B.n559 B.n345 71.676
R868 B.n555 B.n346 71.676
R869 B.n551 B.n347 71.676
R870 B.n547 B.n348 71.676
R871 B.n543 B.n349 71.676
R872 B.n539 B.n350 71.676
R873 B.n535 B.n351 71.676
R874 B.n531 B.n352 71.676
R875 B.n527 B.n353 71.676
R876 B.n523 B.n354 71.676
R877 B.n519 B.n355 71.676
R878 B.n515 B.n356 71.676
R879 B.n511 B.n357 71.676
R880 B.n507 B.n358 71.676
R881 B.n503 B.n359 71.676
R882 B.n499 B.n360 71.676
R883 B.n495 B.n361 71.676
R884 B.n491 B.n362 71.676
R885 B.n487 B.n363 71.676
R886 B.n483 B.n364 71.676
R887 B.n479 B.n365 71.676
R888 B.n475 B.n366 71.676
R889 B.n470 B.n367 71.676
R890 B.n466 B.n368 71.676
R891 B.n462 B.n369 71.676
R892 B.n458 B.n370 71.676
R893 B.n454 B.n371 71.676
R894 B.n450 B.n372 71.676
R895 B.n446 B.n373 71.676
R896 B.n442 B.n374 71.676
R897 B.n438 B.n375 71.676
R898 B.n434 B.n376 71.676
R899 B.n430 B.n377 71.676
R900 B.n426 B.n378 71.676
R901 B.n422 B.n379 71.676
R902 B.n418 B.n380 71.676
R903 B.n414 B.n381 71.676
R904 B.n410 B.n382 71.676
R905 B.n406 B.n383 71.676
R906 B.n402 B.n384 71.676
R907 B.n398 B.n385 71.676
R908 B.n394 B.n386 71.676
R909 B.n574 B.n573 71.676
R910 B.n393 B.t15 69.007
R911 B.n103 B.t19 69.007
R912 B.n390 B.t12 68.9923
R913 B.n106 B.t9 68.9923
R914 B.n472 B.n393 59.5399
R915 B.n391 B.n390 59.5399
R916 B.n189 B.n106 59.5399
R917 B.n104 B.n103 59.5399
R918 B.n579 B.n340 44.274
R919 B.n579 B.n336 44.274
R920 B.n585 B.n336 44.274
R921 B.n585 B.n332 44.274
R922 B.n591 B.n332 44.274
R923 B.n597 B.n328 44.274
R924 B.n597 B.n324 44.274
R925 B.n603 B.n324 44.274
R926 B.n603 B.n320 44.274
R927 B.n609 B.n320 44.274
R928 B.n609 B.n316 44.274
R929 B.n616 B.n316 44.274
R930 B.n616 B.n615 44.274
R931 B.n622 B.n309 44.274
R932 B.n628 B.n309 44.274
R933 B.n628 B.n305 44.274
R934 B.n634 B.n305 44.274
R935 B.n640 B.n301 44.274
R936 B.n640 B.n296 44.274
R937 B.n646 B.n296 44.274
R938 B.n646 B.n297 44.274
R939 B.n653 B.n289 44.274
R940 B.n659 B.n289 44.274
R941 B.n659 B.n4 44.274
R942 B.n760 B.n4 44.274
R943 B.n760 B.n759 44.274
R944 B.n759 B.n758 44.274
R945 B.n758 B.n8 44.274
R946 B.n752 B.n8 44.274
R947 B.n751 B.n750 44.274
R948 B.n750 B.n15 44.274
R949 B.n744 B.n15 44.274
R950 B.n744 B.n743 44.274
R951 B.n742 B.n22 44.274
R952 B.n736 B.n22 44.274
R953 B.n736 B.n735 44.274
R954 B.n735 B.n734 44.274
R955 B.n728 B.n32 44.274
R956 B.n728 B.n727 44.274
R957 B.n727 B.n726 44.274
R958 B.n726 B.n36 44.274
R959 B.n720 B.n36 44.274
R960 B.n720 B.n719 44.274
R961 B.n719 B.n718 44.274
R962 B.n718 B.n43 44.274
R963 B.n712 B.n711 44.274
R964 B.n711 B.n710 44.274
R965 B.n710 B.n50 44.274
R966 B.n704 B.n50 44.274
R967 B.n704 B.n703 44.274
R968 B.n393 B.n392 34.7157
R969 B.n390 B.n389 34.7157
R970 B.n106 B.n105 34.7157
R971 B.n103 B.n102 34.7157
R972 B.n591 B.t11 33.8567
R973 B.n622 B.t1 33.8567
R974 B.n297 B.t2 33.8567
R975 B.t0 B.n751 33.8567
R976 B.n734 B.t5 33.8567
R977 B.n712 B.t7 33.8567
R978 B.n108 B.n52 32.0005
R979 B.n700 B.n699 32.0005
R980 B.n576 B.n575 32.0005
R981 B.n569 B.n338 32.0005
R982 B.n634 B.t3 22.1372
R983 B.t3 B.n301 22.1372
R984 B.n743 B.t4 22.1372
R985 B.t4 B.n742 22.1372
R986 B B.n762 18.0485
R987 B.n109 B.n108 10.6151
R988 B.n112 B.n109 10.6151
R989 B.n113 B.n112 10.6151
R990 B.n116 B.n113 10.6151
R991 B.n117 B.n116 10.6151
R992 B.n120 B.n117 10.6151
R993 B.n121 B.n120 10.6151
R994 B.n124 B.n121 10.6151
R995 B.n125 B.n124 10.6151
R996 B.n128 B.n125 10.6151
R997 B.n129 B.n128 10.6151
R998 B.n132 B.n129 10.6151
R999 B.n133 B.n132 10.6151
R1000 B.n136 B.n133 10.6151
R1001 B.n137 B.n136 10.6151
R1002 B.n140 B.n137 10.6151
R1003 B.n141 B.n140 10.6151
R1004 B.n144 B.n141 10.6151
R1005 B.n145 B.n144 10.6151
R1006 B.n148 B.n145 10.6151
R1007 B.n149 B.n148 10.6151
R1008 B.n152 B.n149 10.6151
R1009 B.n153 B.n152 10.6151
R1010 B.n156 B.n153 10.6151
R1011 B.n157 B.n156 10.6151
R1012 B.n160 B.n157 10.6151
R1013 B.n161 B.n160 10.6151
R1014 B.n164 B.n161 10.6151
R1015 B.n165 B.n164 10.6151
R1016 B.n168 B.n165 10.6151
R1017 B.n169 B.n168 10.6151
R1018 B.n172 B.n169 10.6151
R1019 B.n173 B.n172 10.6151
R1020 B.n176 B.n173 10.6151
R1021 B.n177 B.n176 10.6151
R1022 B.n180 B.n177 10.6151
R1023 B.n181 B.n180 10.6151
R1024 B.n184 B.n181 10.6151
R1025 B.n185 B.n184 10.6151
R1026 B.n188 B.n185 10.6151
R1027 B.n193 B.n190 10.6151
R1028 B.n194 B.n193 10.6151
R1029 B.n197 B.n194 10.6151
R1030 B.n198 B.n197 10.6151
R1031 B.n201 B.n198 10.6151
R1032 B.n202 B.n201 10.6151
R1033 B.n205 B.n202 10.6151
R1034 B.n206 B.n205 10.6151
R1035 B.n210 B.n209 10.6151
R1036 B.n213 B.n210 10.6151
R1037 B.n214 B.n213 10.6151
R1038 B.n217 B.n214 10.6151
R1039 B.n218 B.n217 10.6151
R1040 B.n221 B.n218 10.6151
R1041 B.n222 B.n221 10.6151
R1042 B.n225 B.n222 10.6151
R1043 B.n226 B.n225 10.6151
R1044 B.n229 B.n226 10.6151
R1045 B.n230 B.n229 10.6151
R1046 B.n233 B.n230 10.6151
R1047 B.n234 B.n233 10.6151
R1048 B.n237 B.n234 10.6151
R1049 B.n238 B.n237 10.6151
R1050 B.n241 B.n238 10.6151
R1051 B.n242 B.n241 10.6151
R1052 B.n245 B.n242 10.6151
R1053 B.n246 B.n245 10.6151
R1054 B.n249 B.n246 10.6151
R1055 B.n250 B.n249 10.6151
R1056 B.n253 B.n250 10.6151
R1057 B.n254 B.n253 10.6151
R1058 B.n257 B.n254 10.6151
R1059 B.n258 B.n257 10.6151
R1060 B.n261 B.n258 10.6151
R1061 B.n262 B.n261 10.6151
R1062 B.n265 B.n262 10.6151
R1063 B.n266 B.n265 10.6151
R1064 B.n269 B.n266 10.6151
R1065 B.n270 B.n269 10.6151
R1066 B.n273 B.n270 10.6151
R1067 B.n274 B.n273 10.6151
R1068 B.n277 B.n274 10.6151
R1069 B.n278 B.n277 10.6151
R1070 B.n281 B.n278 10.6151
R1071 B.n282 B.n281 10.6151
R1072 B.n285 B.n282 10.6151
R1073 B.n286 B.n285 10.6151
R1074 B.n700 B.n286 10.6151
R1075 B.n577 B.n576 10.6151
R1076 B.n577 B.n334 10.6151
R1077 B.n587 B.n334 10.6151
R1078 B.n588 B.n587 10.6151
R1079 B.n589 B.n588 10.6151
R1080 B.n589 B.n326 10.6151
R1081 B.n599 B.n326 10.6151
R1082 B.n600 B.n599 10.6151
R1083 B.n601 B.n600 10.6151
R1084 B.n601 B.n318 10.6151
R1085 B.n611 B.n318 10.6151
R1086 B.n612 B.n611 10.6151
R1087 B.n613 B.n612 10.6151
R1088 B.n613 B.n311 10.6151
R1089 B.n624 B.n311 10.6151
R1090 B.n625 B.n624 10.6151
R1091 B.n626 B.n625 10.6151
R1092 B.n626 B.n303 10.6151
R1093 B.n636 B.n303 10.6151
R1094 B.n637 B.n636 10.6151
R1095 B.n638 B.n637 10.6151
R1096 B.n638 B.n294 10.6151
R1097 B.n648 B.n294 10.6151
R1098 B.n649 B.n648 10.6151
R1099 B.n651 B.n649 10.6151
R1100 B.n651 B.n650 10.6151
R1101 B.n650 B.n287 10.6151
R1102 B.n662 B.n287 10.6151
R1103 B.n663 B.n662 10.6151
R1104 B.n664 B.n663 10.6151
R1105 B.n665 B.n664 10.6151
R1106 B.n667 B.n665 10.6151
R1107 B.n668 B.n667 10.6151
R1108 B.n669 B.n668 10.6151
R1109 B.n670 B.n669 10.6151
R1110 B.n672 B.n670 10.6151
R1111 B.n673 B.n672 10.6151
R1112 B.n674 B.n673 10.6151
R1113 B.n675 B.n674 10.6151
R1114 B.n677 B.n675 10.6151
R1115 B.n678 B.n677 10.6151
R1116 B.n679 B.n678 10.6151
R1117 B.n680 B.n679 10.6151
R1118 B.n682 B.n680 10.6151
R1119 B.n683 B.n682 10.6151
R1120 B.n684 B.n683 10.6151
R1121 B.n685 B.n684 10.6151
R1122 B.n687 B.n685 10.6151
R1123 B.n688 B.n687 10.6151
R1124 B.n689 B.n688 10.6151
R1125 B.n690 B.n689 10.6151
R1126 B.n692 B.n690 10.6151
R1127 B.n693 B.n692 10.6151
R1128 B.n694 B.n693 10.6151
R1129 B.n695 B.n694 10.6151
R1130 B.n697 B.n695 10.6151
R1131 B.n698 B.n697 10.6151
R1132 B.n699 B.n698 10.6151
R1133 B.n569 B.n568 10.6151
R1134 B.n568 B.n567 10.6151
R1135 B.n567 B.n566 10.6151
R1136 B.n566 B.n564 10.6151
R1137 B.n564 B.n561 10.6151
R1138 B.n561 B.n560 10.6151
R1139 B.n560 B.n557 10.6151
R1140 B.n557 B.n556 10.6151
R1141 B.n556 B.n553 10.6151
R1142 B.n553 B.n552 10.6151
R1143 B.n552 B.n549 10.6151
R1144 B.n549 B.n548 10.6151
R1145 B.n548 B.n545 10.6151
R1146 B.n545 B.n544 10.6151
R1147 B.n544 B.n541 10.6151
R1148 B.n541 B.n540 10.6151
R1149 B.n540 B.n537 10.6151
R1150 B.n537 B.n536 10.6151
R1151 B.n536 B.n533 10.6151
R1152 B.n533 B.n532 10.6151
R1153 B.n532 B.n529 10.6151
R1154 B.n529 B.n528 10.6151
R1155 B.n528 B.n525 10.6151
R1156 B.n525 B.n524 10.6151
R1157 B.n524 B.n521 10.6151
R1158 B.n521 B.n520 10.6151
R1159 B.n520 B.n517 10.6151
R1160 B.n517 B.n516 10.6151
R1161 B.n516 B.n513 10.6151
R1162 B.n513 B.n512 10.6151
R1163 B.n512 B.n509 10.6151
R1164 B.n509 B.n508 10.6151
R1165 B.n508 B.n505 10.6151
R1166 B.n505 B.n504 10.6151
R1167 B.n504 B.n501 10.6151
R1168 B.n501 B.n500 10.6151
R1169 B.n500 B.n497 10.6151
R1170 B.n497 B.n496 10.6151
R1171 B.n496 B.n493 10.6151
R1172 B.n493 B.n492 10.6151
R1173 B.n489 B.n488 10.6151
R1174 B.n488 B.n485 10.6151
R1175 B.n485 B.n484 10.6151
R1176 B.n484 B.n481 10.6151
R1177 B.n481 B.n480 10.6151
R1178 B.n480 B.n477 10.6151
R1179 B.n477 B.n476 10.6151
R1180 B.n476 B.n473 10.6151
R1181 B.n471 B.n468 10.6151
R1182 B.n468 B.n467 10.6151
R1183 B.n467 B.n464 10.6151
R1184 B.n464 B.n463 10.6151
R1185 B.n463 B.n460 10.6151
R1186 B.n460 B.n459 10.6151
R1187 B.n459 B.n456 10.6151
R1188 B.n456 B.n455 10.6151
R1189 B.n455 B.n452 10.6151
R1190 B.n452 B.n451 10.6151
R1191 B.n451 B.n448 10.6151
R1192 B.n448 B.n447 10.6151
R1193 B.n447 B.n444 10.6151
R1194 B.n444 B.n443 10.6151
R1195 B.n443 B.n440 10.6151
R1196 B.n440 B.n439 10.6151
R1197 B.n439 B.n436 10.6151
R1198 B.n436 B.n435 10.6151
R1199 B.n435 B.n432 10.6151
R1200 B.n432 B.n431 10.6151
R1201 B.n431 B.n428 10.6151
R1202 B.n428 B.n427 10.6151
R1203 B.n427 B.n424 10.6151
R1204 B.n424 B.n423 10.6151
R1205 B.n423 B.n420 10.6151
R1206 B.n420 B.n419 10.6151
R1207 B.n419 B.n416 10.6151
R1208 B.n416 B.n415 10.6151
R1209 B.n415 B.n412 10.6151
R1210 B.n412 B.n411 10.6151
R1211 B.n411 B.n408 10.6151
R1212 B.n408 B.n407 10.6151
R1213 B.n407 B.n404 10.6151
R1214 B.n404 B.n403 10.6151
R1215 B.n403 B.n400 10.6151
R1216 B.n400 B.n399 10.6151
R1217 B.n399 B.n396 10.6151
R1218 B.n396 B.n395 10.6151
R1219 B.n395 B.n342 10.6151
R1220 B.n575 B.n342 10.6151
R1221 B.n581 B.n338 10.6151
R1222 B.n582 B.n581 10.6151
R1223 B.n583 B.n582 10.6151
R1224 B.n583 B.n330 10.6151
R1225 B.n593 B.n330 10.6151
R1226 B.n594 B.n593 10.6151
R1227 B.n595 B.n594 10.6151
R1228 B.n595 B.n322 10.6151
R1229 B.n605 B.n322 10.6151
R1230 B.n606 B.n605 10.6151
R1231 B.n607 B.n606 10.6151
R1232 B.n607 B.n314 10.6151
R1233 B.n618 B.n314 10.6151
R1234 B.n619 B.n618 10.6151
R1235 B.n620 B.n619 10.6151
R1236 B.n620 B.n307 10.6151
R1237 B.n630 B.n307 10.6151
R1238 B.n631 B.n630 10.6151
R1239 B.n632 B.n631 10.6151
R1240 B.n632 B.n299 10.6151
R1241 B.n642 B.n299 10.6151
R1242 B.n643 B.n642 10.6151
R1243 B.n644 B.n643 10.6151
R1244 B.n644 B.n291 10.6151
R1245 B.n655 B.n291 10.6151
R1246 B.n656 B.n655 10.6151
R1247 B.n657 B.n656 10.6151
R1248 B.n657 B.n0 10.6151
R1249 B.n756 B.n1 10.6151
R1250 B.n756 B.n755 10.6151
R1251 B.n755 B.n754 10.6151
R1252 B.n754 B.n10 10.6151
R1253 B.n748 B.n10 10.6151
R1254 B.n748 B.n747 10.6151
R1255 B.n747 B.n746 10.6151
R1256 B.n746 B.n17 10.6151
R1257 B.n740 B.n17 10.6151
R1258 B.n740 B.n739 10.6151
R1259 B.n739 B.n738 10.6151
R1260 B.n738 B.n24 10.6151
R1261 B.n732 B.n24 10.6151
R1262 B.n732 B.n731 10.6151
R1263 B.n731 B.n730 10.6151
R1264 B.n730 B.n30 10.6151
R1265 B.n724 B.n30 10.6151
R1266 B.n724 B.n723 10.6151
R1267 B.n723 B.n722 10.6151
R1268 B.n722 B.n38 10.6151
R1269 B.n716 B.n38 10.6151
R1270 B.n716 B.n715 10.6151
R1271 B.n715 B.n714 10.6151
R1272 B.n714 B.n45 10.6151
R1273 B.n708 B.n45 10.6151
R1274 B.n708 B.n707 10.6151
R1275 B.n707 B.n706 10.6151
R1276 B.n706 B.n52 10.6151
R1277 B.t11 B.n328 10.4178
R1278 B.n615 B.t1 10.4178
R1279 B.n653 B.t2 10.4178
R1280 B.n752 B.t0 10.4178
R1281 B.n32 B.t5 10.4178
R1282 B.t7 B.n43 10.4178
R1283 B.n190 B.n189 6.5566
R1284 B.n206 B.n104 6.5566
R1285 B.n489 B.n391 6.5566
R1286 B.n473 B.n472 6.5566
R1287 B.n189 B.n188 4.05904
R1288 B.n209 B.n104 4.05904
R1289 B.n492 B.n391 4.05904
R1290 B.n472 B.n471 4.05904
R1291 B.n762 B.n0 2.81026
R1292 B.n762 B.n1 2.81026
R1293 VN.n3 VN.t4 228.529
R1294 VN.n13 VN.t3 228.529
R1295 VN.n2 VN.t2 191.81
R1296 VN.n8 VN.t5 191.81
R1297 VN.n12 VN.t0 191.81
R1298 VN.n18 VN.t1 191.81
R1299 VN.n9 VN.n8 171.63
R1300 VN.n19 VN.n18 171.63
R1301 VN.n17 VN.n10 161.3
R1302 VN.n16 VN.n15 161.3
R1303 VN.n14 VN.n11 161.3
R1304 VN.n7 VN.n0 161.3
R1305 VN.n6 VN.n5 161.3
R1306 VN.n4 VN.n1 161.3
R1307 VN.n6 VN.n1 50.7491
R1308 VN.n16 VN.n11 50.7491
R1309 VN VN.n19 44.2789
R1310 VN.n3 VN.n2 41.9508
R1311 VN.n13 VN.n12 41.9508
R1312 VN.n7 VN.n6 30.405
R1313 VN.n17 VN.n16 30.405
R1314 VN.n2 VN.n1 24.5923
R1315 VN.n12 VN.n11 24.5923
R1316 VN.n14 VN.n13 17.3014
R1317 VN.n4 VN.n3 17.3014
R1318 VN.n8 VN.n7 14.2638
R1319 VN.n18 VN.n17 14.2638
R1320 VN.n19 VN.n10 0.189894
R1321 VN.n15 VN.n10 0.189894
R1322 VN.n15 VN.n14 0.189894
R1323 VN.n5 VN.n4 0.189894
R1324 VN.n5 VN.n0 0.189894
R1325 VN.n9 VN.n0 0.189894
R1326 VN VN.n9 0.0516364
R1327 VDD2.n1 VDD2.t2 68.4027
R1328 VDD2.n2 VDD2.t5 67.3017
R1329 VDD2.n1 VDD2.n0 65.9271
R1330 VDD2 VDD2.n3 65.9242
R1331 VDD2.n2 VDD2.n1 38.7476
R1332 VDD2.n3 VDD2.t0 1.70446
R1333 VDD2.n3 VDD2.t3 1.70446
R1334 VDD2.n0 VDD2.t1 1.70446
R1335 VDD2.n0 VDD2.t4 1.70446
R1336 VDD2 VDD2.n2 1.21602
R1337 VTAIL.n7 VTAIL.t8 50.6229
R1338 VTAIL.n11 VTAIL.t6 50.6219
R1339 VTAIL.n2 VTAIL.t0 50.6219
R1340 VTAIL.n10 VTAIL.t3 50.6218
R1341 VTAIL.n9 VTAIL.n8 48.9189
R1342 VTAIL.n6 VTAIL.n5 48.9189
R1343 VTAIL.n1 VTAIL.n0 48.9179
R1344 VTAIL.n4 VTAIL.n3 48.9179
R1345 VTAIL.n6 VTAIL.n4 25.4703
R1346 VTAIL.n11 VTAIL.n10 23.9272
R1347 VTAIL.n0 VTAIL.t7 1.70446
R1348 VTAIL.n0 VTAIL.t9 1.70446
R1349 VTAIL.n3 VTAIL.t4 1.70446
R1350 VTAIL.n3 VTAIL.t1 1.70446
R1351 VTAIL.n8 VTAIL.t5 1.70446
R1352 VTAIL.n8 VTAIL.t2 1.70446
R1353 VTAIL.n5 VTAIL.t10 1.70446
R1354 VTAIL.n5 VTAIL.t11 1.70446
R1355 VTAIL.n7 VTAIL.n6 1.5436
R1356 VTAIL.n10 VTAIL.n9 1.5436
R1357 VTAIL.n4 VTAIL.n2 1.5436
R1358 VTAIL.n9 VTAIL.n7 1.24188
R1359 VTAIL.n2 VTAIL.n1 1.24188
R1360 VTAIL VTAIL.n11 1.09964
R1361 VTAIL VTAIL.n1 0.444466
R1362 VP.n7 VP.t1 228.529
R1363 VP.n20 VP.t0 191.81
R1364 VP.n14 VP.t2 191.81
R1365 VP.n26 VP.t5 191.81
R1366 VP.n6 VP.t3 191.81
R1367 VP.n12 VP.t4 191.81
R1368 VP.n15 VP.n14 171.63
R1369 VP.n27 VP.n26 171.63
R1370 VP.n13 VP.n12 171.63
R1371 VP.n8 VP.n5 161.3
R1372 VP.n10 VP.n9 161.3
R1373 VP.n11 VP.n4 161.3
R1374 VP.n25 VP.n0 161.3
R1375 VP.n24 VP.n23 161.3
R1376 VP.n22 VP.n1 161.3
R1377 VP.n21 VP.n20 161.3
R1378 VP.n19 VP.n2 161.3
R1379 VP.n18 VP.n17 161.3
R1380 VP.n16 VP.n3 161.3
R1381 VP.n19 VP.n18 50.7491
R1382 VP.n24 VP.n1 50.7491
R1383 VP.n10 VP.n5 50.7491
R1384 VP.n15 VP.n13 43.8982
R1385 VP.n7 VP.n6 41.9508
R1386 VP.n18 VP.n3 30.405
R1387 VP.n25 VP.n24 30.405
R1388 VP.n11 VP.n10 30.405
R1389 VP.n20 VP.n19 24.5923
R1390 VP.n20 VP.n1 24.5923
R1391 VP.n6 VP.n5 24.5923
R1392 VP.n8 VP.n7 17.3014
R1393 VP.n14 VP.n3 14.2638
R1394 VP.n26 VP.n25 14.2638
R1395 VP.n12 VP.n11 14.2638
R1396 VP.n9 VP.n8 0.189894
R1397 VP.n9 VP.n4 0.189894
R1398 VP.n13 VP.n4 0.189894
R1399 VP.n16 VP.n15 0.189894
R1400 VP.n17 VP.n16 0.189894
R1401 VP.n17 VP.n2 0.189894
R1402 VP.n21 VP.n2 0.189894
R1403 VP.n22 VP.n21 0.189894
R1404 VP.n23 VP.n22 0.189894
R1405 VP.n23 VP.n0 0.189894
R1406 VP.n27 VP.n0 0.189894
R1407 VP VP.n27 0.0516364
R1408 VDD1 VDD1.t4 68.5172
R1409 VDD1.n1 VDD1.t3 68.4027
R1410 VDD1.n1 VDD1.n0 65.9271
R1411 VDD1.n3 VDD1.n2 65.5966
R1412 VDD1.n3 VDD1.n1 40.1022
R1413 VDD1.n2 VDD1.t2 1.70446
R1414 VDD1.n2 VDD1.t1 1.70446
R1415 VDD1.n0 VDD1.t5 1.70446
R1416 VDD1.n0 VDD1.t0 1.70446
R1417 VDD1 VDD1.n3 0.328086
C0 VP VN 5.7424f
C1 VP VDD1 5.86494f
C2 VDD2 VN 5.656f
C3 VP VTAIL 5.58079f
C4 VDD2 VDD1 0.991663f
C5 VDD1 VN 0.149465f
C6 VDD2 VTAIL 7.89695f
C7 VTAIL VN 5.56637f
C8 VDD1 VTAIL 7.855391f
C9 VDD2 VP 0.362042f
C10 VDD2 B 5.007337f
C11 VDD1 B 5.273879f
C12 VTAIL B 6.859082f
C13 VN B 9.62757f
C14 VP B 8.022514f
C15 VDD1.t4 B 2.31367f
C16 VDD1.t3 B 2.31302f
C17 VDD1.t5 B 0.202501f
C18 VDD1.t0 B 0.202501f
C19 VDD1.n0 B 1.81195f
C20 VDD1.n1 B 2.17215f
C21 VDD1.t2 B 0.202501f
C22 VDD1.t1 B 0.202501f
C23 VDD1.n2 B 1.81036f
C24 VDD1.n3 B 2.1424f
C25 VP.n0 B 0.033557f
C26 VP.t5 B 1.5497f
C27 VP.n1 B 0.060962f
C28 VP.n2 B 0.033557f
C29 VP.t0 B 1.5497f
C30 VP.n3 B 0.05379f
C31 VP.n4 B 0.033557f
C32 VP.t4 B 1.5497f
C33 VP.n5 B 0.060962f
C34 VP.t1 B 1.66092f
C35 VP.t3 B 1.5497f
C36 VP.n6 B 0.64016f
C37 VP.n7 B 0.628783f
C38 VP.n8 B 0.213423f
C39 VP.n9 B 0.033557f
C40 VP.n10 B 0.032136f
C41 VP.n11 B 0.05379f
C42 VP.n12 B 0.635463f
C43 VP.n13 B 1.49408f
C44 VP.t2 B 1.5497f
C45 VP.n14 B 0.635463f
C46 VP.n15 B 1.52163f
C47 VP.n16 B 0.033557f
C48 VP.n17 B 0.033557f
C49 VP.n18 B 0.032136f
C50 VP.n19 B 0.060962f
C51 VP.n20 B 0.594051f
C52 VP.n21 B 0.033557f
C53 VP.n22 B 0.033557f
C54 VP.n23 B 0.033557f
C55 VP.n24 B 0.032136f
C56 VP.n25 B 0.05379f
C57 VP.n26 B 0.635463f
C58 VP.n27 B 0.030675f
C59 VTAIL.t7 B 0.215372f
C60 VTAIL.t9 B 0.215372f
C61 VTAIL.n0 B 1.86438f
C62 VTAIL.n1 B 0.340097f
C63 VTAIL.t0 B 2.37648f
C64 VTAIL.n2 B 0.498447f
C65 VTAIL.t4 B 0.215372f
C66 VTAIL.t1 B 0.215372f
C67 VTAIL.n3 B 1.86438f
C68 VTAIL.n4 B 1.63826f
C69 VTAIL.t10 B 0.215372f
C70 VTAIL.t11 B 0.215372f
C71 VTAIL.n5 B 1.86437f
C72 VTAIL.n6 B 1.63827f
C73 VTAIL.t8 B 2.37648f
C74 VTAIL.n7 B 0.498449f
C75 VTAIL.t5 B 0.215372f
C76 VTAIL.t2 B 0.215372f
C77 VTAIL.n8 B 1.86437f
C78 VTAIL.n9 B 0.423173f
C79 VTAIL.t3 B 2.37647f
C80 VTAIL.n10 B 1.59693f
C81 VTAIL.t6 B 2.37648f
C82 VTAIL.n11 B 1.56337f
C83 VDD2.t2 B 2.29303f
C84 VDD2.t1 B 0.200751f
C85 VDD2.t4 B 0.200751f
C86 VDD2.n0 B 1.79629f
C87 VDD2.n1 B 2.07025f
C88 VDD2.t5 B 2.288f
C89 VDD2.n2 B 2.13432f
C90 VDD2.t0 B 0.200751f
C91 VDD2.t3 B 0.200751f
C92 VDD2.n3 B 1.79626f
C93 VN.n0 B 0.033076f
C94 VN.t5 B 1.52749f
C95 VN.n1 B 0.060089f
C96 VN.t4 B 1.63711f
C97 VN.t2 B 1.52749f
C98 VN.n2 B 0.630986f
C99 VN.n3 B 0.619772f
C100 VN.n4 B 0.210365f
C101 VN.n5 B 0.033076f
C102 VN.n6 B 0.031675f
C103 VN.n7 B 0.053019f
C104 VN.n8 B 0.626356f
C105 VN.n9 B 0.030235f
C106 VN.n10 B 0.033076f
C107 VN.t1 B 1.52749f
C108 VN.n11 B 0.060089f
C109 VN.t3 B 1.63711f
C110 VN.t0 B 1.52749f
C111 VN.n12 B 0.630986f
C112 VN.n13 B 0.619772f
C113 VN.n14 B 0.210365f
C114 VN.n15 B 0.033076f
C115 VN.n16 B 0.031675f
C116 VN.n17 B 0.053019f
C117 VN.n18 B 0.626356f
C118 VN.n19 B 1.49432f
.ends

