* NGSPICE file created from diff_pair_sample_1729.ext - technology: sky130A

.subckt diff_pair_sample_1729 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t10 VN.t0 VDD2.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=2.1021 pd=13.07 as=2.1021 ps=13.07 w=12.74 l=3.07
X1 VDD1.t5 VP.t0 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=2.1021 pd=13.07 as=4.9686 ps=26.26 w=12.74 l=3.07
X2 VDD1.t4 VP.t1 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=4.9686 pd=26.26 as=2.1021 ps=13.07 w=12.74 l=3.07
X3 B.t19 B.t17 B.t18 B.t14 sky130_fd_pr__nfet_01v8 ad=4.9686 pd=26.26 as=0 ps=0 w=12.74 l=3.07
X4 VTAIL.t9 VN.t1 VDD2.t1 B.t5 sky130_fd_pr__nfet_01v8 ad=2.1021 pd=13.07 as=2.1021 ps=13.07 w=12.74 l=3.07
X5 B.t16 B.t13 B.t15 B.t14 sky130_fd_pr__nfet_01v8 ad=4.9686 pd=26.26 as=0 ps=0 w=12.74 l=3.07
X6 B.t12 B.t10 B.t11 B.t7 sky130_fd_pr__nfet_01v8 ad=4.9686 pd=26.26 as=0 ps=0 w=12.74 l=3.07
X7 VDD2.t3 VN.t2 VTAIL.t8 B.t2 sky130_fd_pr__nfet_01v8 ad=4.9686 pd=26.26 as=2.1021 ps=13.07 w=12.74 l=3.07
X8 VTAIL.t11 VP.t2 VDD1.t3 B.t5 sky130_fd_pr__nfet_01v8 ad=2.1021 pd=13.07 as=2.1021 ps=13.07 w=12.74 l=3.07
X9 VDD2.t5 VN.t3 VTAIL.t7 B.t1 sky130_fd_pr__nfet_01v8 ad=4.9686 pd=26.26 as=2.1021 ps=13.07 w=12.74 l=3.07
X10 VDD1.t2 VP.t3 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=4.9686 pd=26.26 as=2.1021 ps=13.07 w=12.74 l=3.07
X11 VDD2.t4 VN.t4 VTAIL.t6 B.t3 sky130_fd_pr__nfet_01v8 ad=2.1021 pd=13.07 as=4.9686 ps=26.26 w=12.74 l=3.07
X12 B.t9 B.t6 B.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=4.9686 pd=26.26 as=0 ps=0 w=12.74 l=3.07
X13 VDD1.t1 VP.t4 VTAIL.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=2.1021 pd=13.07 as=4.9686 ps=26.26 w=12.74 l=3.07
X14 VTAIL.t0 VP.t5 VDD1.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=2.1021 pd=13.07 as=2.1021 ps=13.07 w=12.74 l=3.07
X15 VDD2.t2 VN.t5 VTAIL.t5 B.t4 sky130_fd_pr__nfet_01v8 ad=2.1021 pd=13.07 as=4.9686 ps=26.26 w=12.74 l=3.07
R0 VN.n30 VN.n29 161.3
R1 VN.n28 VN.n17 161.3
R2 VN.n27 VN.n26 161.3
R3 VN.n25 VN.n18 161.3
R4 VN.n24 VN.n23 161.3
R5 VN.n22 VN.n19 161.3
R6 VN.n14 VN.n13 161.3
R7 VN.n12 VN.n1 161.3
R8 VN.n11 VN.n10 161.3
R9 VN.n9 VN.n2 161.3
R10 VN.n8 VN.n7 161.3
R11 VN.n6 VN.n3 161.3
R12 VN.n20 VN.t4 133.322
R13 VN.n4 VN.t2 133.322
R14 VN.n5 VN.t1 100.011
R15 VN.n0 VN.t5 100.011
R16 VN.n21 VN.t0 100.011
R17 VN.n16 VN.t3 100.011
R18 VN.n15 VN.n0 70.4162
R19 VN.n31 VN.n16 70.4162
R20 VN.n11 VN.n2 56.4773
R21 VN.n27 VN.n18 56.4773
R22 VN VN.n31 51.3767
R23 VN.n5 VN.n4 49.2698
R24 VN.n21 VN.n20 49.2698
R25 VN.n6 VN.n5 24.3439
R26 VN.n7 VN.n6 24.3439
R27 VN.n7 VN.n2 24.3439
R28 VN.n12 VN.n11 24.3439
R29 VN.n13 VN.n12 24.3439
R30 VN.n23 VN.n18 24.3439
R31 VN.n23 VN.n22 24.3439
R32 VN.n22 VN.n21 24.3439
R33 VN.n29 VN.n28 24.3439
R34 VN.n28 VN.n27 24.3439
R35 VN.n13 VN.n0 19.4752
R36 VN.n29 VN.n16 19.4752
R37 VN.n20 VN.n19 3.94998
R38 VN.n4 VN.n3 3.94998
R39 VN.n31 VN.n30 0.355081
R40 VN.n15 VN.n14 0.355081
R41 VN VN.n15 0.26685
R42 VN.n30 VN.n17 0.189894
R43 VN.n26 VN.n17 0.189894
R44 VN.n26 VN.n25 0.189894
R45 VN.n25 VN.n24 0.189894
R46 VN.n24 VN.n19 0.189894
R47 VN.n8 VN.n3 0.189894
R48 VN.n9 VN.n8 0.189894
R49 VN.n10 VN.n9 0.189894
R50 VN.n10 VN.n1 0.189894
R51 VN.n14 VN.n1 0.189894
R52 VDD2.n135 VDD2.n71 289.615
R53 VDD2.n64 VDD2.n0 289.615
R54 VDD2.n136 VDD2.n135 185
R55 VDD2.n134 VDD2.n133 185
R56 VDD2.n75 VDD2.n74 185
R57 VDD2.n128 VDD2.n127 185
R58 VDD2.n126 VDD2.n125 185
R59 VDD2.n79 VDD2.n78 185
R60 VDD2.n120 VDD2.n119 185
R61 VDD2.n118 VDD2.n117 185
R62 VDD2.n116 VDD2.n82 185
R63 VDD2.n86 VDD2.n83 185
R64 VDD2.n111 VDD2.n110 185
R65 VDD2.n109 VDD2.n108 185
R66 VDD2.n88 VDD2.n87 185
R67 VDD2.n103 VDD2.n102 185
R68 VDD2.n101 VDD2.n100 185
R69 VDD2.n92 VDD2.n91 185
R70 VDD2.n95 VDD2.n94 185
R71 VDD2.n23 VDD2.n22 185
R72 VDD2.n20 VDD2.n19 185
R73 VDD2.n29 VDD2.n28 185
R74 VDD2.n31 VDD2.n30 185
R75 VDD2.n16 VDD2.n15 185
R76 VDD2.n37 VDD2.n36 185
R77 VDD2.n40 VDD2.n39 185
R78 VDD2.n38 VDD2.n12 185
R79 VDD2.n45 VDD2.n11 185
R80 VDD2.n47 VDD2.n46 185
R81 VDD2.n49 VDD2.n48 185
R82 VDD2.n8 VDD2.n7 185
R83 VDD2.n55 VDD2.n54 185
R84 VDD2.n57 VDD2.n56 185
R85 VDD2.n4 VDD2.n3 185
R86 VDD2.n63 VDD2.n62 185
R87 VDD2.n65 VDD2.n64 185
R88 VDD2.t5 VDD2.n93 149.524
R89 VDD2.t3 VDD2.n21 149.524
R90 VDD2.n135 VDD2.n134 104.615
R91 VDD2.n134 VDD2.n74 104.615
R92 VDD2.n127 VDD2.n74 104.615
R93 VDD2.n127 VDD2.n126 104.615
R94 VDD2.n126 VDD2.n78 104.615
R95 VDD2.n119 VDD2.n78 104.615
R96 VDD2.n119 VDD2.n118 104.615
R97 VDD2.n118 VDD2.n82 104.615
R98 VDD2.n86 VDD2.n82 104.615
R99 VDD2.n110 VDD2.n86 104.615
R100 VDD2.n110 VDD2.n109 104.615
R101 VDD2.n109 VDD2.n87 104.615
R102 VDD2.n102 VDD2.n87 104.615
R103 VDD2.n102 VDD2.n101 104.615
R104 VDD2.n101 VDD2.n91 104.615
R105 VDD2.n94 VDD2.n91 104.615
R106 VDD2.n22 VDD2.n19 104.615
R107 VDD2.n29 VDD2.n19 104.615
R108 VDD2.n30 VDD2.n29 104.615
R109 VDD2.n30 VDD2.n15 104.615
R110 VDD2.n37 VDD2.n15 104.615
R111 VDD2.n39 VDD2.n37 104.615
R112 VDD2.n39 VDD2.n38 104.615
R113 VDD2.n38 VDD2.n11 104.615
R114 VDD2.n47 VDD2.n11 104.615
R115 VDD2.n48 VDD2.n47 104.615
R116 VDD2.n48 VDD2.n7 104.615
R117 VDD2.n55 VDD2.n7 104.615
R118 VDD2.n56 VDD2.n55 104.615
R119 VDD2.n56 VDD2.n3 104.615
R120 VDD2.n63 VDD2.n3 104.615
R121 VDD2.n64 VDD2.n63 104.615
R122 VDD2.n70 VDD2.n69 60.4413
R123 VDD2 VDD2.n141 60.4383
R124 VDD2.n94 VDD2.t5 52.3082
R125 VDD2.n22 VDD2.t3 52.3082
R126 VDD2.n70 VDD2.n68 49.0677
R127 VDD2.n140 VDD2.n139 46.9247
R128 VDD2.n140 VDD2.n70 44.2239
R129 VDD2.n117 VDD2.n116 13.1884
R130 VDD2.n46 VDD2.n45 13.1884
R131 VDD2.n120 VDD2.n81 12.8005
R132 VDD2.n115 VDD2.n83 12.8005
R133 VDD2.n44 VDD2.n12 12.8005
R134 VDD2.n49 VDD2.n10 12.8005
R135 VDD2.n121 VDD2.n79 12.0247
R136 VDD2.n112 VDD2.n111 12.0247
R137 VDD2.n41 VDD2.n40 12.0247
R138 VDD2.n50 VDD2.n8 12.0247
R139 VDD2.n125 VDD2.n124 11.249
R140 VDD2.n108 VDD2.n85 11.249
R141 VDD2.n36 VDD2.n14 11.249
R142 VDD2.n54 VDD2.n53 11.249
R143 VDD2.n128 VDD2.n77 10.4732
R144 VDD2.n107 VDD2.n88 10.4732
R145 VDD2.n35 VDD2.n16 10.4732
R146 VDD2.n57 VDD2.n6 10.4732
R147 VDD2.n95 VDD2.n93 10.2747
R148 VDD2.n23 VDD2.n21 10.2747
R149 VDD2.n129 VDD2.n75 9.69747
R150 VDD2.n104 VDD2.n103 9.69747
R151 VDD2.n32 VDD2.n31 9.69747
R152 VDD2.n58 VDD2.n4 9.69747
R153 VDD2.n139 VDD2.n138 9.45567
R154 VDD2.n68 VDD2.n67 9.45567
R155 VDD2.n97 VDD2.n96 9.3005
R156 VDD2.n99 VDD2.n98 9.3005
R157 VDD2.n90 VDD2.n89 9.3005
R158 VDD2.n105 VDD2.n104 9.3005
R159 VDD2.n107 VDD2.n106 9.3005
R160 VDD2.n85 VDD2.n84 9.3005
R161 VDD2.n113 VDD2.n112 9.3005
R162 VDD2.n115 VDD2.n114 9.3005
R163 VDD2.n138 VDD2.n137 9.3005
R164 VDD2.n73 VDD2.n72 9.3005
R165 VDD2.n132 VDD2.n131 9.3005
R166 VDD2.n130 VDD2.n129 9.3005
R167 VDD2.n77 VDD2.n76 9.3005
R168 VDD2.n124 VDD2.n123 9.3005
R169 VDD2.n122 VDD2.n121 9.3005
R170 VDD2.n81 VDD2.n80 9.3005
R171 VDD2.n2 VDD2.n1 9.3005
R172 VDD2.n61 VDD2.n60 9.3005
R173 VDD2.n59 VDD2.n58 9.3005
R174 VDD2.n6 VDD2.n5 9.3005
R175 VDD2.n53 VDD2.n52 9.3005
R176 VDD2.n51 VDD2.n50 9.3005
R177 VDD2.n10 VDD2.n9 9.3005
R178 VDD2.n25 VDD2.n24 9.3005
R179 VDD2.n27 VDD2.n26 9.3005
R180 VDD2.n18 VDD2.n17 9.3005
R181 VDD2.n33 VDD2.n32 9.3005
R182 VDD2.n35 VDD2.n34 9.3005
R183 VDD2.n14 VDD2.n13 9.3005
R184 VDD2.n42 VDD2.n41 9.3005
R185 VDD2.n44 VDD2.n43 9.3005
R186 VDD2.n67 VDD2.n66 9.3005
R187 VDD2.n133 VDD2.n132 8.92171
R188 VDD2.n100 VDD2.n90 8.92171
R189 VDD2.n28 VDD2.n18 8.92171
R190 VDD2.n62 VDD2.n61 8.92171
R191 VDD2.n136 VDD2.n73 8.14595
R192 VDD2.n99 VDD2.n92 8.14595
R193 VDD2.n27 VDD2.n20 8.14595
R194 VDD2.n65 VDD2.n2 8.14595
R195 VDD2.n137 VDD2.n71 7.3702
R196 VDD2.n96 VDD2.n95 7.3702
R197 VDD2.n24 VDD2.n23 7.3702
R198 VDD2.n66 VDD2.n0 7.3702
R199 VDD2.n139 VDD2.n71 6.59444
R200 VDD2.n68 VDD2.n0 6.59444
R201 VDD2.n137 VDD2.n136 5.81868
R202 VDD2.n96 VDD2.n92 5.81868
R203 VDD2.n24 VDD2.n20 5.81868
R204 VDD2.n66 VDD2.n65 5.81868
R205 VDD2.n133 VDD2.n73 5.04292
R206 VDD2.n100 VDD2.n99 5.04292
R207 VDD2.n28 VDD2.n27 5.04292
R208 VDD2.n62 VDD2.n2 5.04292
R209 VDD2.n132 VDD2.n75 4.26717
R210 VDD2.n103 VDD2.n90 4.26717
R211 VDD2.n31 VDD2.n18 4.26717
R212 VDD2.n61 VDD2.n4 4.26717
R213 VDD2.n129 VDD2.n128 3.49141
R214 VDD2.n104 VDD2.n88 3.49141
R215 VDD2.n32 VDD2.n16 3.49141
R216 VDD2.n58 VDD2.n57 3.49141
R217 VDD2.n97 VDD2.n93 2.84303
R218 VDD2.n25 VDD2.n21 2.84303
R219 VDD2.n125 VDD2.n77 2.71565
R220 VDD2.n108 VDD2.n107 2.71565
R221 VDD2.n36 VDD2.n35 2.71565
R222 VDD2.n54 VDD2.n6 2.71565
R223 VDD2 VDD2.n140 2.25697
R224 VDD2.n124 VDD2.n79 1.93989
R225 VDD2.n111 VDD2.n85 1.93989
R226 VDD2.n40 VDD2.n14 1.93989
R227 VDD2.n53 VDD2.n8 1.93989
R228 VDD2.n141 VDD2.t0 1.55466
R229 VDD2.n141 VDD2.t4 1.55466
R230 VDD2.n69 VDD2.t1 1.55466
R231 VDD2.n69 VDD2.t2 1.55466
R232 VDD2.n121 VDD2.n120 1.16414
R233 VDD2.n112 VDD2.n83 1.16414
R234 VDD2.n41 VDD2.n12 1.16414
R235 VDD2.n50 VDD2.n49 1.16414
R236 VDD2.n117 VDD2.n81 0.388379
R237 VDD2.n116 VDD2.n115 0.388379
R238 VDD2.n45 VDD2.n44 0.388379
R239 VDD2.n46 VDD2.n10 0.388379
R240 VDD2.n138 VDD2.n72 0.155672
R241 VDD2.n131 VDD2.n72 0.155672
R242 VDD2.n131 VDD2.n130 0.155672
R243 VDD2.n130 VDD2.n76 0.155672
R244 VDD2.n123 VDD2.n76 0.155672
R245 VDD2.n123 VDD2.n122 0.155672
R246 VDD2.n122 VDD2.n80 0.155672
R247 VDD2.n114 VDD2.n80 0.155672
R248 VDD2.n114 VDD2.n113 0.155672
R249 VDD2.n113 VDD2.n84 0.155672
R250 VDD2.n106 VDD2.n84 0.155672
R251 VDD2.n106 VDD2.n105 0.155672
R252 VDD2.n105 VDD2.n89 0.155672
R253 VDD2.n98 VDD2.n89 0.155672
R254 VDD2.n98 VDD2.n97 0.155672
R255 VDD2.n26 VDD2.n25 0.155672
R256 VDD2.n26 VDD2.n17 0.155672
R257 VDD2.n33 VDD2.n17 0.155672
R258 VDD2.n34 VDD2.n33 0.155672
R259 VDD2.n34 VDD2.n13 0.155672
R260 VDD2.n42 VDD2.n13 0.155672
R261 VDD2.n43 VDD2.n42 0.155672
R262 VDD2.n43 VDD2.n9 0.155672
R263 VDD2.n51 VDD2.n9 0.155672
R264 VDD2.n52 VDD2.n51 0.155672
R265 VDD2.n52 VDD2.n5 0.155672
R266 VDD2.n59 VDD2.n5 0.155672
R267 VDD2.n60 VDD2.n59 0.155672
R268 VDD2.n60 VDD2.n1 0.155672
R269 VDD2.n67 VDD2.n1 0.155672
R270 VTAIL.n282 VTAIL.n218 289.615
R271 VTAIL.n66 VTAIL.n2 289.615
R272 VTAIL.n212 VTAIL.n148 289.615
R273 VTAIL.n140 VTAIL.n76 289.615
R274 VTAIL.n241 VTAIL.n240 185
R275 VTAIL.n238 VTAIL.n237 185
R276 VTAIL.n247 VTAIL.n246 185
R277 VTAIL.n249 VTAIL.n248 185
R278 VTAIL.n234 VTAIL.n233 185
R279 VTAIL.n255 VTAIL.n254 185
R280 VTAIL.n258 VTAIL.n257 185
R281 VTAIL.n256 VTAIL.n230 185
R282 VTAIL.n263 VTAIL.n229 185
R283 VTAIL.n265 VTAIL.n264 185
R284 VTAIL.n267 VTAIL.n266 185
R285 VTAIL.n226 VTAIL.n225 185
R286 VTAIL.n273 VTAIL.n272 185
R287 VTAIL.n275 VTAIL.n274 185
R288 VTAIL.n222 VTAIL.n221 185
R289 VTAIL.n281 VTAIL.n280 185
R290 VTAIL.n283 VTAIL.n282 185
R291 VTAIL.n25 VTAIL.n24 185
R292 VTAIL.n22 VTAIL.n21 185
R293 VTAIL.n31 VTAIL.n30 185
R294 VTAIL.n33 VTAIL.n32 185
R295 VTAIL.n18 VTAIL.n17 185
R296 VTAIL.n39 VTAIL.n38 185
R297 VTAIL.n42 VTAIL.n41 185
R298 VTAIL.n40 VTAIL.n14 185
R299 VTAIL.n47 VTAIL.n13 185
R300 VTAIL.n49 VTAIL.n48 185
R301 VTAIL.n51 VTAIL.n50 185
R302 VTAIL.n10 VTAIL.n9 185
R303 VTAIL.n57 VTAIL.n56 185
R304 VTAIL.n59 VTAIL.n58 185
R305 VTAIL.n6 VTAIL.n5 185
R306 VTAIL.n65 VTAIL.n64 185
R307 VTAIL.n67 VTAIL.n66 185
R308 VTAIL.n213 VTAIL.n212 185
R309 VTAIL.n211 VTAIL.n210 185
R310 VTAIL.n152 VTAIL.n151 185
R311 VTAIL.n205 VTAIL.n204 185
R312 VTAIL.n203 VTAIL.n202 185
R313 VTAIL.n156 VTAIL.n155 185
R314 VTAIL.n197 VTAIL.n196 185
R315 VTAIL.n195 VTAIL.n194 185
R316 VTAIL.n193 VTAIL.n159 185
R317 VTAIL.n163 VTAIL.n160 185
R318 VTAIL.n188 VTAIL.n187 185
R319 VTAIL.n186 VTAIL.n185 185
R320 VTAIL.n165 VTAIL.n164 185
R321 VTAIL.n180 VTAIL.n179 185
R322 VTAIL.n178 VTAIL.n177 185
R323 VTAIL.n169 VTAIL.n168 185
R324 VTAIL.n172 VTAIL.n171 185
R325 VTAIL.n141 VTAIL.n140 185
R326 VTAIL.n139 VTAIL.n138 185
R327 VTAIL.n80 VTAIL.n79 185
R328 VTAIL.n133 VTAIL.n132 185
R329 VTAIL.n131 VTAIL.n130 185
R330 VTAIL.n84 VTAIL.n83 185
R331 VTAIL.n125 VTAIL.n124 185
R332 VTAIL.n123 VTAIL.n122 185
R333 VTAIL.n121 VTAIL.n87 185
R334 VTAIL.n91 VTAIL.n88 185
R335 VTAIL.n116 VTAIL.n115 185
R336 VTAIL.n114 VTAIL.n113 185
R337 VTAIL.n93 VTAIL.n92 185
R338 VTAIL.n108 VTAIL.n107 185
R339 VTAIL.n106 VTAIL.n105 185
R340 VTAIL.n97 VTAIL.n96 185
R341 VTAIL.n100 VTAIL.n99 185
R342 VTAIL.t5 VTAIL.n239 149.524
R343 VTAIL.t3 VTAIL.n23 149.524
R344 VTAIL.t4 VTAIL.n170 149.524
R345 VTAIL.t6 VTAIL.n98 149.524
R346 VTAIL.n240 VTAIL.n237 104.615
R347 VTAIL.n247 VTAIL.n237 104.615
R348 VTAIL.n248 VTAIL.n247 104.615
R349 VTAIL.n248 VTAIL.n233 104.615
R350 VTAIL.n255 VTAIL.n233 104.615
R351 VTAIL.n257 VTAIL.n255 104.615
R352 VTAIL.n257 VTAIL.n256 104.615
R353 VTAIL.n256 VTAIL.n229 104.615
R354 VTAIL.n265 VTAIL.n229 104.615
R355 VTAIL.n266 VTAIL.n265 104.615
R356 VTAIL.n266 VTAIL.n225 104.615
R357 VTAIL.n273 VTAIL.n225 104.615
R358 VTAIL.n274 VTAIL.n273 104.615
R359 VTAIL.n274 VTAIL.n221 104.615
R360 VTAIL.n281 VTAIL.n221 104.615
R361 VTAIL.n282 VTAIL.n281 104.615
R362 VTAIL.n24 VTAIL.n21 104.615
R363 VTAIL.n31 VTAIL.n21 104.615
R364 VTAIL.n32 VTAIL.n31 104.615
R365 VTAIL.n32 VTAIL.n17 104.615
R366 VTAIL.n39 VTAIL.n17 104.615
R367 VTAIL.n41 VTAIL.n39 104.615
R368 VTAIL.n41 VTAIL.n40 104.615
R369 VTAIL.n40 VTAIL.n13 104.615
R370 VTAIL.n49 VTAIL.n13 104.615
R371 VTAIL.n50 VTAIL.n49 104.615
R372 VTAIL.n50 VTAIL.n9 104.615
R373 VTAIL.n57 VTAIL.n9 104.615
R374 VTAIL.n58 VTAIL.n57 104.615
R375 VTAIL.n58 VTAIL.n5 104.615
R376 VTAIL.n65 VTAIL.n5 104.615
R377 VTAIL.n66 VTAIL.n65 104.615
R378 VTAIL.n212 VTAIL.n211 104.615
R379 VTAIL.n211 VTAIL.n151 104.615
R380 VTAIL.n204 VTAIL.n151 104.615
R381 VTAIL.n204 VTAIL.n203 104.615
R382 VTAIL.n203 VTAIL.n155 104.615
R383 VTAIL.n196 VTAIL.n155 104.615
R384 VTAIL.n196 VTAIL.n195 104.615
R385 VTAIL.n195 VTAIL.n159 104.615
R386 VTAIL.n163 VTAIL.n159 104.615
R387 VTAIL.n187 VTAIL.n163 104.615
R388 VTAIL.n187 VTAIL.n186 104.615
R389 VTAIL.n186 VTAIL.n164 104.615
R390 VTAIL.n179 VTAIL.n164 104.615
R391 VTAIL.n179 VTAIL.n178 104.615
R392 VTAIL.n178 VTAIL.n168 104.615
R393 VTAIL.n171 VTAIL.n168 104.615
R394 VTAIL.n140 VTAIL.n139 104.615
R395 VTAIL.n139 VTAIL.n79 104.615
R396 VTAIL.n132 VTAIL.n79 104.615
R397 VTAIL.n132 VTAIL.n131 104.615
R398 VTAIL.n131 VTAIL.n83 104.615
R399 VTAIL.n124 VTAIL.n83 104.615
R400 VTAIL.n124 VTAIL.n123 104.615
R401 VTAIL.n123 VTAIL.n87 104.615
R402 VTAIL.n91 VTAIL.n87 104.615
R403 VTAIL.n115 VTAIL.n91 104.615
R404 VTAIL.n115 VTAIL.n114 104.615
R405 VTAIL.n114 VTAIL.n92 104.615
R406 VTAIL.n107 VTAIL.n92 104.615
R407 VTAIL.n107 VTAIL.n106 104.615
R408 VTAIL.n106 VTAIL.n96 104.615
R409 VTAIL.n99 VTAIL.n96 104.615
R410 VTAIL.n240 VTAIL.t5 52.3082
R411 VTAIL.n24 VTAIL.t3 52.3082
R412 VTAIL.n171 VTAIL.t4 52.3082
R413 VTAIL.n99 VTAIL.t6 52.3082
R414 VTAIL.n1 VTAIL.n0 43.0851
R415 VTAIL.n73 VTAIL.n72 43.0851
R416 VTAIL.n147 VTAIL.n146 43.0851
R417 VTAIL.n75 VTAIL.n74 43.0851
R418 VTAIL.n287 VTAIL.n286 30.246
R419 VTAIL.n71 VTAIL.n70 30.246
R420 VTAIL.n217 VTAIL.n216 30.246
R421 VTAIL.n145 VTAIL.n144 30.246
R422 VTAIL.n75 VTAIL.n73 29.2117
R423 VTAIL.n287 VTAIL.n217 26.2807
R424 VTAIL.n264 VTAIL.n263 13.1884
R425 VTAIL.n48 VTAIL.n47 13.1884
R426 VTAIL.n194 VTAIL.n193 13.1884
R427 VTAIL.n122 VTAIL.n121 13.1884
R428 VTAIL.n262 VTAIL.n230 12.8005
R429 VTAIL.n267 VTAIL.n228 12.8005
R430 VTAIL.n46 VTAIL.n14 12.8005
R431 VTAIL.n51 VTAIL.n12 12.8005
R432 VTAIL.n197 VTAIL.n158 12.8005
R433 VTAIL.n192 VTAIL.n160 12.8005
R434 VTAIL.n125 VTAIL.n86 12.8005
R435 VTAIL.n120 VTAIL.n88 12.8005
R436 VTAIL.n259 VTAIL.n258 12.0247
R437 VTAIL.n268 VTAIL.n226 12.0247
R438 VTAIL.n43 VTAIL.n42 12.0247
R439 VTAIL.n52 VTAIL.n10 12.0247
R440 VTAIL.n198 VTAIL.n156 12.0247
R441 VTAIL.n189 VTAIL.n188 12.0247
R442 VTAIL.n126 VTAIL.n84 12.0247
R443 VTAIL.n117 VTAIL.n116 12.0247
R444 VTAIL.n254 VTAIL.n232 11.249
R445 VTAIL.n272 VTAIL.n271 11.249
R446 VTAIL.n38 VTAIL.n16 11.249
R447 VTAIL.n56 VTAIL.n55 11.249
R448 VTAIL.n202 VTAIL.n201 11.249
R449 VTAIL.n185 VTAIL.n162 11.249
R450 VTAIL.n130 VTAIL.n129 11.249
R451 VTAIL.n113 VTAIL.n90 11.249
R452 VTAIL.n253 VTAIL.n234 10.4732
R453 VTAIL.n275 VTAIL.n224 10.4732
R454 VTAIL.n37 VTAIL.n18 10.4732
R455 VTAIL.n59 VTAIL.n8 10.4732
R456 VTAIL.n205 VTAIL.n154 10.4732
R457 VTAIL.n184 VTAIL.n165 10.4732
R458 VTAIL.n133 VTAIL.n82 10.4732
R459 VTAIL.n112 VTAIL.n93 10.4732
R460 VTAIL.n241 VTAIL.n239 10.2747
R461 VTAIL.n25 VTAIL.n23 10.2747
R462 VTAIL.n172 VTAIL.n170 10.2747
R463 VTAIL.n100 VTAIL.n98 10.2747
R464 VTAIL.n250 VTAIL.n249 9.69747
R465 VTAIL.n276 VTAIL.n222 9.69747
R466 VTAIL.n34 VTAIL.n33 9.69747
R467 VTAIL.n60 VTAIL.n6 9.69747
R468 VTAIL.n206 VTAIL.n152 9.69747
R469 VTAIL.n181 VTAIL.n180 9.69747
R470 VTAIL.n134 VTAIL.n80 9.69747
R471 VTAIL.n109 VTAIL.n108 9.69747
R472 VTAIL.n286 VTAIL.n285 9.45567
R473 VTAIL.n70 VTAIL.n69 9.45567
R474 VTAIL.n216 VTAIL.n215 9.45567
R475 VTAIL.n144 VTAIL.n143 9.45567
R476 VTAIL.n220 VTAIL.n219 9.3005
R477 VTAIL.n279 VTAIL.n278 9.3005
R478 VTAIL.n277 VTAIL.n276 9.3005
R479 VTAIL.n224 VTAIL.n223 9.3005
R480 VTAIL.n271 VTAIL.n270 9.3005
R481 VTAIL.n269 VTAIL.n268 9.3005
R482 VTAIL.n228 VTAIL.n227 9.3005
R483 VTAIL.n243 VTAIL.n242 9.3005
R484 VTAIL.n245 VTAIL.n244 9.3005
R485 VTAIL.n236 VTAIL.n235 9.3005
R486 VTAIL.n251 VTAIL.n250 9.3005
R487 VTAIL.n253 VTAIL.n252 9.3005
R488 VTAIL.n232 VTAIL.n231 9.3005
R489 VTAIL.n260 VTAIL.n259 9.3005
R490 VTAIL.n262 VTAIL.n261 9.3005
R491 VTAIL.n285 VTAIL.n284 9.3005
R492 VTAIL.n4 VTAIL.n3 9.3005
R493 VTAIL.n63 VTAIL.n62 9.3005
R494 VTAIL.n61 VTAIL.n60 9.3005
R495 VTAIL.n8 VTAIL.n7 9.3005
R496 VTAIL.n55 VTAIL.n54 9.3005
R497 VTAIL.n53 VTAIL.n52 9.3005
R498 VTAIL.n12 VTAIL.n11 9.3005
R499 VTAIL.n27 VTAIL.n26 9.3005
R500 VTAIL.n29 VTAIL.n28 9.3005
R501 VTAIL.n20 VTAIL.n19 9.3005
R502 VTAIL.n35 VTAIL.n34 9.3005
R503 VTAIL.n37 VTAIL.n36 9.3005
R504 VTAIL.n16 VTAIL.n15 9.3005
R505 VTAIL.n44 VTAIL.n43 9.3005
R506 VTAIL.n46 VTAIL.n45 9.3005
R507 VTAIL.n69 VTAIL.n68 9.3005
R508 VTAIL.n174 VTAIL.n173 9.3005
R509 VTAIL.n176 VTAIL.n175 9.3005
R510 VTAIL.n167 VTAIL.n166 9.3005
R511 VTAIL.n182 VTAIL.n181 9.3005
R512 VTAIL.n184 VTAIL.n183 9.3005
R513 VTAIL.n162 VTAIL.n161 9.3005
R514 VTAIL.n190 VTAIL.n189 9.3005
R515 VTAIL.n192 VTAIL.n191 9.3005
R516 VTAIL.n215 VTAIL.n214 9.3005
R517 VTAIL.n150 VTAIL.n149 9.3005
R518 VTAIL.n209 VTAIL.n208 9.3005
R519 VTAIL.n207 VTAIL.n206 9.3005
R520 VTAIL.n154 VTAIL.n153 9.3005
R521 VTAIL.n201 VTAIL.n200 9.3005
R522 VTAIL.n199 VTAIL.n198 9.3005
R523 VTAIL.n158 VTAIL.n157 9.3005
R524 VTAIL.n102 VTAIL.n101 9.3005
R525 VTAIL.n104 VTAIL.n103 9.3005
R526 VTAIL.n95 VTAIL.n94 9.3005
R527 VTAIL.n110 VTAIL.n109 9.3005
R528 VTAIL.n112 VTAIL.n111 9.3005
R529 VTAIL.n90 VTAIL.n89 9.3005
R530 VTAIL.n118 VTAIL.n117 9.3005
R531 VTAIL.n120 VTAIL.n119 9.3005
R532 VTAIL.n143 VTAIL.n142 9.3005
R533 VTAIL.n78 VTAIL.n77 9.3005
R534 VTAIL.n137 VTAIL.n136 9.3005
R535 VTAIL.n135 VTAIL.n134 9.3005
R536 VTAIL.n82 VTAIL.n81 9.3005
R537 VTAIL.n129 VTAIL.n128 9.3005
R538 VTAIL.n127 VTAIL.n126 9.3005
R539 VTAIL.n86 VTAIL.n85 9.3005
R540 VTAIL.n246 VTAIL.n236 8.92171
R541 VTAIL.n280 VTAIL.n279 8.92171
R542 VTAIL.n30 VTAIL.n20 8.92171
R543 VTAIL.n64 VTAIL.n63 8.92171
R544 VTAIL.n210 VTAIL.n209 8.92171
R545 VTAIL.n177 VTAIL.n167 8.92171
R546 VTAIL.n138 VTAIL.n137 8.92171
R547 VTAIL.n105 VTAIL.n95 8.92171
R548 VTAIL.n245 VTAIL.n238 8.14595
R549 VTAIL.n283 VTAIL.n220 8.14595
R550 VTAIL.n29 VTAIL.n22 8.14595
R551 VTAIL.n67 VTAIL.n4 8.14595
R552 VTAIL.n213 VTAIL.n150 8.14595
R553 VTAIL.n176 VTAIL.n169 8.14595
R554 VTAIL.n141 VTAIL.n78 8.14595
R555 VTAIL.n104 VTAIL.n97 8.14595
R556 VTAIL.n242 VTAIL.n241 7.3702
R557 VTAIL.n284 VTAIL.n218 7.3702
R558 VTAIL.n26 VTAIL.n25 7.3702
R559 VTAIL.n68 VTAIL.n2 7.3702
R560 VTAIL.n214 VTAIL.n148 7.3702
R561 VTAIL.n173 VTAIL.n172 7.3702
R562 VTAIL.n142 VTAIL.n76 7.3702
R563 VTAIL.n101 VTAIL.n100 7.3702
R564 VTAIL.n286 VTAIL.n218 6.59444
R565 VTAIL.n70 VTAIL.n2 6.59444
R566 VTAIL.n216 VTAIL.n148 6.59444
R567 VTAIL.n144 VTAIL.n76 6.59444
R568 VTAIL.n242 VTAIL.n238 5.81868
R569 VTAIL.n284 VTAIL.n283 5.81868
R570 VTAIL.n26 VTAIL.n22 5.81868
R571 VTAIL.n68 VTAIL.n67 5.81868
R572 VTAIL.n214 VTAIL.n213 5.81868
R573 VTAIL.n173 VTAIL.n169 5.81868
R574 VTAIL.n142 VTAIL.n141 5.81868
R575 VTAIL.n101 VTAIL.n97 5.81868
R576 VTAIL.n246 VTAIL.n245 5.04292
R577 VTAIL.n280 VTAIL.n220 5.04292
R578 VTAIL.n30 VTAIL.n29 5.04292
R579 VTAIL.n64 VTAIL.n4 5.04292
R580 VTAIL.n210 VTAIL.n150 5.04292
R581 VTAIL.n177 VTAIL.n176 5.04292
R582 VTAIL.n138 VTAIL.n78 5.04292
R583 VTAIL.n105 VTAIL.n104 5.04292
R584 VTAIL.n249 VTAIL.n236 4.26717
R585 VTAIL.n279 VTAIL.n222 4.26717
R586 VTAIL.n33 VTAIL.n20 4.26717
R587 VTAIL.n63 VTAIL.n6 4.26717
R588 VTAIL.n209 VTAIL.n152 4.26717
R589 VTAIL.n180 VTAIL.n167 4.26717
R590 VTAIL.n137 VTAIL.n80 4.26717
R591 VTAIL.n108 VTAIL.n95 4.26717
R592 VTAIL.n250 VTAIL.n234 3.49141
R593 VTAIL.n276 VTAIL.n275 3.49141
R594 VTAIL.n34 VTAIL.n18 3.49141
R595 VTAIL.n60 VTAIL.n59 3.49141
R596 VTAIL.n206 VTAIL.n205 3.49141
R597 VTAIL.n181 VTAIL.n165 3.49141
R598 VTAIL.n134 VTAIL.n133 3.49141
R599 VTAIL.n109 VTAIL.n93 3.49141
R600 VTAIL.n145 VTAIL.n75 2.93153
R601 VTAIL.n217 VTAIL.n147 2.93153
R602 VTAIL.n73 VTAIL.n71 2.93153
R603 VTAIL.n243 VTAIL.n239 2.84303
R604 VTAIL.n27 VTAIL.n23 2.84303
R605 VTAIL.n174 VTAIL.n170 2.84303
R606 VTAIL.n102 VTAIL.n98 2.84303
R607 VTAIL.n254 VTAIL.n253 2.71565
R608 VTAIL.n272 VTAIL.n224 2.71565
R609 VTAIL.n38 VTAIL.n37 2.71565
R610 VTAIL.n56 VTAIL.n8 2.71565
R611 VTAIL.n202 VTAIL.n154 2.71565
R612 VTAIL.n185 VTAIL.n184 2.71565
R613 VTAIL.n130 VTAIL.n82 2.71565
R614 VTAIL.n113 VTAIL.n112 2.71565
R615 VTAIL VTAIL.n287 2.14059
R616 VTAIL.n258 VTAIL.n232 1.93989
R617 VTAIL.n271 VTAIL.n226 1.93989
R618 VTAIL.n42 VTAIL.n16 1.93989
R619 VTAIL.n55 VTAIL.n10 1.93989
R620 VTAIL.n201 VTAIL.n156 1.93989
R621 VTAIL.n188 VTAIL.n162 1.93989
R622 VTAIL.n129 VTAIL.n84 1.93989
R623 VTAIL.n116 VTAIL.n90 1.93989
R624 VTAIL.n147 VTAIL.n145 1.93584
R625 VTAIL.n71 VTAIL.n1 1.93584
R626 VTAIL.n0 VTAIL.t8 1.55466
R627 VTAIL.n0 VTAIL.t9 1.55466
R628 VTAIL.n72 VTAIL.t1 1.55466
R629 VTAIL.n72 VTAIL.t0 1.55466
R630 VTAIL.n146 VTAIL.t2 1.55466
R631 VTAIL.n146 VTAIL.t11 1.55466
R632 VTAIL.n74 VTAIL.t7 1.55466
R633 VTAIL.n74 VTAIL.t10 1.55466
R634 VTAIL.n259 VTAIL.n230 1.16414
R635 VTAIL.n268 VTAIL.n267 1.16414
R636 VTAIL.n43 VTAIL.n14 1.16414
R637 VTAIL.n52 VTAIL.n51 1.16414
R638 VTAIL.n198 VTAIL.n197 1.16414
R639 VTAIL.n189 VTAIL.n160 1.16414
R640 VTAIL.n126 VTAIL.n125 1.16414
R641 VTAIL.n117 VTAIL.n88 1.16414
R642 VTAIL VTAIL.n1 0.791448
R643 VTAIL.n263 VTAIL.n262 0.388379
R644 VTAIL.n264 VTAIL.n228 0.388379
R645 VTAIL.n47 VTAIL.n46 0.388379
R646 VTAIL.n48 VTAIL.n12 0.388379
R647 VTAIL.n194 VTAIL.n158 0.388379
R648 VTAIL.n193 VTAIL.n192 0.388379
R649 VTAIL.n122 VTAIL.n86 0.388379
R650 VTAIL.n121 VTAIL.n120 0.388379
R651 VTAIL.n244 VTAIL.n243 0.155672
R652 VTAIL.n244 VTAIL.n235 0.155672
R653 VTAIL.n251 VTAIL.n235 0.155672
R654 VTAIL.n252 VTAIL.n251 0.155672
R655 VTAIL.n252 VTAIL.n231 0.155672
R656 VTAIL.n260 VTAIL.n231 0.155672
R657 VTAIL.n261 VTAIL.n260 0.155672
R658 VTAIL.n261 VTAIL.n227 0.155672
R659 VTAIL.n269 VTAIL.n227 0.155672
R660 VTAIL.n270 VTAIL.n269 0.155672
R661 VTAIL.n270 VTAIL.n223 0.155672
R662 VTAIL.n277 VTAIL.n223 0.155672
R663 VTAIL.n278 VTAIL.n277 0.155672
R664 VTAIL.n278 VTAIL.n219 0.155672
R665 VTAIL.n285 VTAIL.n219 0.155672
R666 VTAIL.n28 VTAIL.n27 0.155672
R667 VTAIL.n28 VTAIL.n19 0.155672
R668 VTAIL.n35 VTAIL.n19 0.155672
R669 VTAIL.n36 VTAIL.n35 0.155672
R670 VTAIL.n36 VTAIL.n15 0.155672
R671 VTAIL.n44 VTAIL.n15 0.155672
R672 VTAIL.n45 VTAIL.n44 0.155672
R673 VTAIL.n45 VTAIL.n11 0.155672
R674 VTAIL.n53 VTAIL.n11 0.155672
R675 VTAIL.n54 VTAIL.n53 0.155672
R676 VTAIL.n54 VTAIL.n7 0.155672
R677 VTAIL.n61 VTAIL.n7 0.155672
R678 VTAIL.n62 VTAIL.n61 0.155672
R679 VTAIL.n62 VTAIL.n3 0.155672
R680 VTAIL.n69 VTAIL.n3 0.155672
R681 VTAIL.n215 VTAIL.n149 0.155672
R682 VTAIL.n208 VTAIL.n149 0.155672
R683 VTAIL.n208 VTAIL.n207 0.155672
R684 VTAIL.n207 VTAIL.n153 0.155672
R685 VTAIL.n200 VTAIL.n153 0.155672
R686 VTAIL.n200 VTAIL.n199 0.155672
R687 VTAIL.n199 VTAIL.n157 0.155672
R688 VTAIL.n191 VTAIL.n157 0.155672
R689 VTAIL.n191 VTAIL.n190 0.155672
R690 VTAIL.n190 VTAIL.n161 0.155672
R691 VTAIL.n183 VTAIL.n161 0.155672
R692 VTAIL.n183 VTAIL.n182 0.155672
R693 VTAIL.n182 VTAIL.n166 0.155672
R694 VTAIL.n175 VTAIL.n166 0.155672
R695 VTAIL.n175 VTAIL.n174 0.155672
R696 VTAIL.n143 VTAIL.n77 0.155672
R697 VTAIL.n136 VTAIL.n77 0.155672
R698 VTAIL.n136 VTAIL.n135 0.155672
R699 VTAIL.n135 VTAIL.n81 0.155672
R700 VTAIL.n128 VTAIL.n81 0.155672
R701 VTAIL.n128 VTAIL.n127 0.155672
R702 VTAIL.n127 VTAIL.n85 0.155672
R703 VTAIL.n119 VTAIL.n85 0.155672
R704 VTAIL.n119 VTAIL.n118 0.155672
R705 VTAIL.n118 VTAIL.n89 0.155672
R706 VTAIL.n111 VTAIL.n89 0.155672
R707 VTAIL.n111 VTAIL.n110 0.155672
R708 VTAIL.n110 VTAIL.n94 0.155672
R709 VTAIL.n103 VTAIL.n94 0.155672
R710 VTAIL.n103 VTAIL.n102 0.155672
R711 B.n882 B.n881 585
R712 B.n883 B.n882 585
R713 B.n333 B.n138 585
R714 B.n332 B.n331 585
R715 B.n330 B.n329 585
R716 B.n328 B.n327 585
R717 B.n326 B.n325 585
R718 B.n324 B.n323 585
R719 B.n322 B.n321 585
R720 B.n320 B.n319 585
R721 B.n318 B.n317 585
R722 B.n316 B.n315 585
R723 B.n314 B.n313 585
R724 B.n312 B.n311 585
R725 B.n310 B.n309 585
R726 B.n308 B.n307 585
R727 B.n306 B.n305 585
R728 B.n304 B.n303 585
R729 B.n302 B.n301 585
R730 B.n300 B.n299 585
R731 B.n298 B.n297 585
R732 B.n296 B.n295 585
R733 B.n294 B.n293 585
R734 B.n292 B.n291 585
R735 B.n290 B.n289 585
R736 B.n288 B.n287 585
R737 B.n286 B.n285 585
R738 B.n284 B.n283 585
R739 B.n282 B.n281 585
R740 B.n280 B.n279 585
R741 B.n278 B.n277 585
R742 B.n276 B.n275 585
R743 B.n274 B.n273 585
R744 B.n272 B.n271 585
R745 B.n270 B.n269 585
R746 B.n268 B.n267 585
R747 B.n266 B.n265 585
R748 B.n264 B.n263 585
R749 B.n262 B.n261 585
R750 B.n260 B.n259 585
R751 B.n258 B.n257 585
R752 B.n256 B.n255 585
R753 B.n254 B.n253 585
R754 B.n252 B.n251 585
R755 B.n250 B.n249 585
R756 B.n247 B.n246 585
R757 B.n245 B.n244 585
R758 B.n243 B.n242 585
R759 B.n241 B.n240 585
R760 B.n239 B.n238 585
R761 B.n237 B.n236 585
R762 B.n235 B.n234 585
R763 B.n233 B.n232 585
R764 B.n231 B.n230 585
R765 B.n229 B.n228 585
R766 B.n227 B.n226 585
R767 B.n225 B.n224 585
R768 B.n223 B.n222 585
R769 B.n221 B.n220 585
R770 B.n219 B.n218 585
R771 B.n217 B.n216 585
R772 B.n215 B.n214 585
R773 B.n213 B.n212 585
R774 B.n211 B.n210 585
R775 B.n209 B.n208 585
R776 B.n207 B.n206 585
R777 B.n205 B.n204 585
R778 B.n203 B.n202 585
R779 B.n201 B.n200 585
R780 B.n199 B.n198 585
R781 B.n197 B.n196 585
R782 B.n195 B.n194 585
R783 B.n193 B.n192 585
R784 B.n191 B.n190 585
R785 B.n189 B.n188 585
R786 B.n187 B.n186 585
R787 B.n185 B.n184 585
R788 B.n183 B.n182 585
R789 B.n181 B.n180 585
R790 B.n179 B.n178 585
R791 B.n177 B.n176 585
R792 B.n175 B.n174 585
R793 B.n173 B.n172 585
R794 B.n171 B.n170 585
R795 B.n169 B.n168 585
R796 B.n167 B.n166 585
R797 B.n165 B.n164 585
R798 B.n163 B.n162 585
R799 B.n161 B.n160 585
R800 B.n159 B.n158 585
R801 B.n157 B.n156 585
R802 B.n155 B.n154 585
R803 B.n153 B.n152 585
R804 B.n151 B.n150 585
R805 B.n149 B.n148 585
R806 B.n147 B.n146 585
R807 B.n145 B.n144 585
R808 B.n88 B.n87 585
R809 B.n880 B.n89 585
R810 B.n884 B.n89 585
R811 B.n879 B.n878 585
R812 B.n878 B.n85 585
R813 B.n877 B.n84 585
R814 B.n890 B.n84 585
R815 B.n876 B.n83 585
R816 B.n891 B.n83 585
R817 B.n875 B.n82 585
R818 B.n892 B.n82 585
R819 B.n874 B.n873 585
R820 B.n873 B.n78 585
R821 B.n872 B.n77 585
R822 B.n898 B.n77 585
R823 B.n871 B.n76 585
R824 B.n899 B.n76 585
R825 B.n870 B.n75 585
R826 B.n900 B.n75 585
R827 B.n869 B.n868 585
R828 B.n868 B.n71 585
R829 B.n867 B.n70 585
R830 B.n906 B.n70 585
R831 B.n866 B.n69 585
R832 B.n907 B.n69 585
R833 B.n865 B.n68 585
R834 B.n908 B.n68 585
R835 B.n864 B.n863 585
R836 B.n863 B.n64 585
R837 B.n862 B.n63 585
R838 B.n914 B.n63 585
R839 B.n861 B.n62 585
R840 B.n915 B.n62 585
R841 B.n860 B.n61 585
R842 B.n916 B.n61 585
R843 B.n859 B.n858 585
R844 B.n858 B.n57 585
R845 B.n857 B.n56 585
R846 B.n922 B.n56 585
R847 B.n856 B.n55 585
R848 B.n923 B.n55 585
R849 B.n855 B.n54 585
R850 B.n924 B.n54 585
R851 B.n854 B.n853 585
R852 B.n853 B.n53 585
R853 B.n852 B.n49 585
R854 B.n930 B.n49 585
R855 B.n851 B.n48 585
R856 B.n931 B.n48 585
R857 B.n850 B.n47 585
R858 B.n932 B.n47 585
R859 B.n849 B.n848 585
R860 B.n848 B.n43 585
R861 B.n847 B.n42 585
R862 B.n938 B.n42 585
R863 B.n846 B.n41 585
R864 B.n939 B.n41 585
R865 B.n845 B.n40 585
R866 B.n940 B.n40 585
R867 B.n844 B.n843 585
R868 B.n843 B.n36 585
R869 B.n842 B.n35 585
R870 B.n946 B.n35 585
R871 B.n841 B.n34 585
R872 B.n947 B.n34 585
R873 B.n840 B.n33 585
R874 B.n948 B.n33 585
R875 B.n839 B.n838 585
R876 B.n838 B.n29 585
R877 B.n837 B.n28 585
R878 B.n954 B.n28 585
R879 B.n836 B.n27 585
R880 B.n955 B.n27 585
R881 B.n835 B.n26 585
R882 B.n956 B.n26 585
R883 B.n834 B.n833 585
R884 B.n833 B.n22 585
R885 B.n832 B.n21 585
R886 B.n962 B.n21 585
R887 B.n831 B.n20 585
R888 B.n963 B.n20 585
R889 B.n830 B.n19 585
R890 B.n964 B.n19 585
R891 B.n829 B.n828 585
R892 B.n828 B.n18 585
R893 B.n827 B.n14 585
R894 B.n970 B.n14 585
R895 B.n826 B.n13 585
R896 B.n971 B.n13 585
R897 B.n825 B.n12 585
R898 B.n972 B.n12 585
R899 B.n824 B.n823 585
R900 B.n823 B.n8 585
R901 B.n822 B.n7 585
R902 B.n978 B.n7 585
R903 B.n821 B.n6 585
R904 B.n979 B.n6 585
R905 B.n820 B.n5 585
R906 B.n980 B.n5 585
R907 B.n819 B.n818 585
R908 B.n818 B.n4 585
R909 B.n817 B.n334 585
R910 B.n817 B.n816 585
R911 B.n807 B.n335 585
R912 B.n336 B.n335 585
R913 B.n809 B.n808 585
R914 B.n810 B.n809 585
R915 B.n806 B.n341 585
R916 B.n341 B.n340 585
R917 B.n805 B.n804 585
R918 B.n804 B.n803 585
R919 B.n343 B.n342 585
R920 B.n796 B.n343 585
R921 B.n795 B.n794 585
R922 B.n797 B.n795 585
R923 B.n793 B.n348 585
R924 B.n348 B.n347 585
R925 B.n792 B.n791 585
R926 B.n791 B.n790 585
R927 B.n350 B.n349 585
R928 B.n351 B.n350 585
R929 B.n783 B.n782 585
R930 B.n784 B.n783 585
R931 B.n781 B.n356 585
R932 B.n356 B.n355 585
R933 B.n780 B.n779 585
R934 B.n779 B.n778 585
R935 B.n358 B.n357 585
R936 B.n359 B.n358 585
R937 B.n771 B.n770 585
R938 B.n772 B.n771 585
R939 B.n769 B.n363 585
R940 B.n367 B.n363 585
R941 B.n768 B.n767 585
R942 B.n767 B.n766 585
R943 B.n365 B.n364 585
R944 B.n366 B.n365 585
R945 B.n759 B.n758 585
R946 B.n760 B.n759 585
R947 B.n757 B.n372 585
R948 B.n372 B.n371 585
R949 B.n756 B.n755 585
R950 B.n755 B.n754 585
R951 B.n374 B.n373 585
R952 B.n375 B.n374 585
R953 B.n747 B.n746 585
R954 B.n748 B.n747 585
R955 B.n745 B.n380 585
R956 B.n380 B.n379 585
R957 B.n744 B.n743 585
R958 B.n743 B.n742 585
R959 B.n382 B.n381 585
R960 B.n735 B.n382 585
R961 B.n734 B.n733 585
R962 B.n736 B.n734 585
R963 B.n732 B.n387 585
R964 B.n387 B.n386 585
R965 B.n731 B.n730 585
R966 B.n730 B.n729 585
R967 B.n389 B.n388 585
R968 B.n390 B.n389 585
R969 B.n722 B.n721 585
R970 B.n723 B.n722 585
R971 B.n720 B.n395 585
R972 B.n395 B.n394 585
R973 B.n719 B.n718 585
R974 B.n718 B.n717 585
R975 B.n397 B.n396 585
R976 B.n398 B.n397 585
R977 B.n710 B.n709 585
R978 B.n711 B.n710 585
R979 B.n708 B.n403 585
R980 B.n403 B.n402 585
R981 B.n707 B.n706 585
R982 B.n706 B.n705 585
R983 B.n405 B.n404 585
R984 B.n406 B.n405 585
R985 B.n698 B.n697 585
R986 B.n699 B.n698 585
R987 B.n696 B.n411 585
R988 B.n411 B.n410 585
R989 B.n695 B.n694 585
R990 B.n694 B.n693 585
R991 B.n413 B.n412 585
R992 B.n414 B.n413 585
R993 B.n686 B.n685 585
R994 B.n687 B.n686 585
R995 B.n684 B.n419 585
R996 B.n419 B.n418 585
R997 B.n683 B.n682 585
R998 B.n682 B.n681 585
R999 B.n421 B.n420 585
R1000 B.n422 B.n421 585
R1001 B.n674 B.n673 585
R1002 B.n675 B.n674 585
R1003 B.n425 B.n424 585
R1004 B.n481 B.n479 585
R1005 B.n482 B.n478 585
R1006 B.n482 B.n426 585
R1007 B.n485 B.n484 585
R1008 B.n486 B.n477 585
R1009 B.n488 B.n487 585
R1010 B.n490 B.n476 585
R1011 B.n493 B.n492 585
R1012 B.n494 B.n475 585
R1013 B.n496 B.n495 585
R1014 B.n498 B.n474 585
R1015 B.n501 B.n500 585
R1016 B.n502 B.n473 585
R1017 B.n504 B.n503 585
R1018 B.n506 B.n472 585
R1019 B.n509 B.n508 585
R1020 B.n510 B.n471 585
R1021 B.n512 B.n511 585
R1022 B.n514 B.n470 585
R1023 B.n517 B.n516 585
R1024 B.n518 B.n469 585
R1025 B.n520 B.n519 585
R1026 B.n522 B.n468 585
R1027 B.n525 B.n524 585
R1028 B.n526 B.n467 585
R1029 B.n528 B.n527 585
R1030 B.n530 B.n466 585
R1031 B.n533 B.n532 585
R1032 B.n534 B.n465 585
R1033 B.n536 B.n535 585
R1034 B.n538 B.n464 585
R1035 B.n541 B.n540 585
R1036 B.n542 B.n463 585
R1037 B.n544 B.n543 585
R1038 B.n546 B.n462 585
R1039 B.n549 B.n548 585
R1040 B.n550 B.n461 585
R1041 B.n552 B.n551 585
R1042 B.n554 B.n460 585
R1043 B.n557 B.n556 585
R1044 B.n558 B.n459 585
R1045 B.n560 B.n559 585
R1046 B.n562 B.n458 585
R1047 B.n565 B.n564 585
R1048 B.n567 B.n455 585
R1049 B.n569 B.n568 585
R1050 B.n571 B.n454 585
R1051 B.n574 B.n573 585
R1052 B.n575 B.n453 585
R1053 B.n577 B.n576 585
R1054 B.n579 B.n452 585
R1055 B.n582 B.n581 585
R1056 B.n583 B.n449 585
R1057 B.n586 B.n585 585
R1058 B.n588 B.n448 585
R1059 B.n591 B.n590 585
R1060 B.n592 B.n447 585
R1061 B.n594 B.n593 585
R1062 B.n596 B.n446 585
R1063 B.n599 B.n598 585
R1064 B.n600 B.n445 585
R1065 B.n602 B.n601 585
R1066 B.n604 B.n444 585
R1067 B.n607 B.n606 585
R1068 B.n608 B.n443 585
R1069 B.n610 B.n609 585
R1070 B.n612 B.n442 585
R1071 B.n615 B.n614 585
R1072 B.n616 B.n441 585
R1073 B.n618 B.n617 585
R1074 B.n620 B.n440 585
R1075 B.n623 B.n622 585
R1076 B.n624 B.n439 585
R1077 B.n626 B.n625 585
R1078 B.n628 B.n438 585
R1079 B.n631 B.n630 585
R1080 B.n632 B.n437 585
R1081 B.n634 B.n633 585
R1082 B.n636 B.n436 585
R1083 B.n639 B.n638 585
R1084 B.n640 B.n435 585
R1085 B.n642 B.n641 585
R1086 B.n644 B.n434 585
R1087 B.n647 B.n646 585
R1088 B.n648 B.n433 585
R1089 B.n650 B.n649 585
R1090 B.n652 B.n432 585
R1091 B.n655 B.n654 585
R1092 B.n656 B.n431 585
R1093 B.n658 B.n657 585
R1094 B.n660 B.n430 585
R1095 B.n663 B.n662 585
R1096 B.n664 B.n429 585
R1097 B.n666 B.n665 585
R1098 B.n668 B.n428 585
R1099 B.n671 B.n670 585
R1100 B.n672 B.n427 585
R1101 B.n677 B.n676 585
R1102 B.n676 B.n675 585
R1103 B.n678 B.n423 585
R1104 B.n423 B.n422 585
R1105 B.n680 B.n679 585
R1106 B.n681 B.n680 585
R1107 B.n417 B.n416 585
R1108 B.n418 B.n417 585
R1109 B.n689 B.n688 585
R1110 B.n688 B.n687 585
R1111 B.n690 B.n415 585
R1112 B.n415 B.n414 585
R1113 B.n692 B.n691 585
R1114 B.n693 B.n692 585
R1115 B.n409 B.n408 585
R1116 B.n410 B.n409 585
R1117 B.n701 B.n700 585
R1118 B.n700 B.n699 585
R1119 B.n702 B.n407 585
R1120 B.n407 B.n406 585
R1121 B.n704 B.n703 585
R1122 B.n705 B.n704 585
R1123 B.n401 B.n400 585
R1124 B.n402 B.n401 585
R1125 B.n713 B.n712 585
R1126 B.n712 B.n711 585
R1127 B.n714 B.n399 585
R1128 B.n399 B.n398 585
R1129 B.n716 B.n715 585
R1130 B.n717 B.n716 585
R1131 B.n393 B.n392 585
R1132 B.n394 B.n393 585
R1133 B.n725 B.n724 585
R1134 B.n724 B.n723 585
R1135 B.n726 B.n391 585
R1136 B.n391 B.n390 585
R1137 B.n728 B.n727 585
R1138 B.n729 B.n728 585
R1139 B.n385 B.n384 585
R1140 B.n386 B.n385 585
R1141 B.n738 B.n737 585
R1142 B.n737 B.n736 585
R1143 B.n739 B.n383 585
R1144 B.n735 B.n383 585
R1145 B.n741 B.n740 585
R1146 B.n742 B.n741 585
R1147 B.n378 B.n377 585
R1148 B.n379 B.n378 585
R1149 B.n750 B.n749 585
R1150 B.n749 B.n748 585
R1151 B.n751 B.n376 585
R1152 B.n376 B.n375 585
R1153 B.n753 B.n752 585
R1154 B.n754 B.n753 585
R1155 B.n370 B.n369 585
R1156 B.n371 B.n370 585
R1157 B.n762 B.n761 585
R1158 B.n761 B.n760 585
R1159 B.n763 B.n368 585
R1160 B.n368 B.n366 585
R1161 B.n765 B.n764 585
R1162 B.n766 B.n765 585
R1163 B.n362 B.n361 585
R1164 B.n367 B.n362 585
R1165 B.n774 B.n773 585
R1166 B.n773 B.n772 585
R1167 B.n775 B.n360 585
R1168 B.n360 B.n359 585
R1169 B.n777 B.n776 585
R1170 B.n778 B.n777 585
R1171 B.n354 B.n353 585
R1172 B.n355 B.n354 585
R1173 B.n786 B.n785 585
R1174 B.n785 B.n784 585
R1175 B.n787 B.n352 585
R1176 B.n352 B.n351 585
R1177 B.n789 B.n788 585
R1178 B.n790 B.n789 585
R1179 B.n346 B.n345 585
R1180 B.n347 B.n346 585
R1181 B.n799 B.n798 585
R1182 B.n798 B.n797 585
R1183 B.n800 B.n344 585
R1184 B.n796 B.n344 585
R1185 B.n802 B.n801 585
R1186 B.n803 B.n802 585
R1187 B.n339 B.n338 585
R1188 B.n340 B.n339 585
R1189 B.n812 B.n811 585
R1190 B.n811 B.n810 585
R1191 B.n813 B.n337 585
R1192 B.n337 B.n336 585
R1193 B.n815 B.n814 585
R1194 B.n816 B.n815 585
R1195 B.n2 B.n0 585
R1196 B.n4 B.n2 585
R1197 B.n3 B.n1 585
R1198 B.n979 B.n3 585
R1199 B.n977 B.n976 585
R1200 B.n978 B.n977 585
R1201 B.n975 B.n9 585
R1202 B.n9 B.n8 585
R1203 B.n974 B.n973 585
R1204 B.n973 B.n972 585
R1205 B.n11 B.n10 585
R1206 B.n971 B.n11 585
R1207 B.n969 B.n968 585
R1208 B.n970 B.n969 585
R1209 B.n967 B.n15 585
R1210 B.n18 B.n15 585
R1211 B.n966 B.n965 585
R1212 B.n965 B.n964 585
R1213 B.n17 B.n16 585
R1214 B.n963 B.n17 585
R1215 B.n961 B.n960 585
R1216 B.n962 B.n961 585
R1217 B.n959 B.n23 585
R1218 B.n23 B.n22 585
R1219 B.n958 B.n957 585
R1220 B.n957 B.n956 585
R1221 B.n25 B.n24 585
R1222 B.n955 B.n25 585
R1223 B.n953 B.n952 585
R1224 B.n954 B.n953 585
R1225 B.n951 B.n30 585
R1226 B.n30 B.n29 585
R1227 B.n950 B.n949 585
R1228 B.n949 B.n948 585
R1229 B.n32 B.n31 585
R1230 B.n947 B.n32 585
R1231 B.n945 B.n944 585
R1232 B.n946 B.n945 585
R1233 B.n943 B.n37 585
R1234 B.n37 B.n36 585
R1235 B.n942 B.n941 585
R1236 B.n941 B.n940 585
R1237 B.n39 B.n38 585
R1238 B.n939 B.n39 585
R1239 B.n937 B.n936 585
R1240 B.n938 B.n937 585
R1241 B.n935 B.n44 585
R1242 B.n44 B.n43 585
R1243 B.n934 B.n933 585
R1244 B.n933 B.n932 585
R1245 B.n46 B.n45 585
R1246 B.n931 B.n46 585
R1247 B.n929 B.n928 585
R1248 B.n930 B.n929 585
R1249 B.n927 B.n50 585
R1250 B.n53 B.n50 585
R1251 B.n926 B.n925 585
R1252 B.n925 B.n924 585
R1253 B.n52 B.n51 585
R1254 B.n923 B.n52 585
R1255 B.n921 B.n920 585
R1256 B.n922 B.n921 585
R1257 B.n919 B.n58 585
R1258 B.n58 B.n57 585
R1259 B.n918 B.n917 585
R1260 B.n917 B.n916 585
R1261 B.n60 B.n59 585
R1262 B.n915 B.n60 585
R1263 B.n913 B.n912 585
R1264 B.n914 B.n913 585
R1265 B.n911 B.n65 585
R1266 B.n65 B.n64 585
R1267 B.n910 B.n909 585
R1268 B.n909 B.n908 585
R1269 B.n67 B.n66 585
R1270 B.n907 B.n67 585
R1271 B.n905 B.n904 585
R1272 B.n906 B.n905 585
R1273 B.n903 B.n72 585
R1274 B.n72 B.n71 585
R1275 B.n902 B.n901 585
R1276 B.n901 B.n900 585
R1277 B.n74 B.n73 585
R1278 B.n899 B.n74 585
R1279 B.n897 B.n896 585
R1280 B.n898 B.n897 585
R1281 B.n895 B.n79 585
R1282 B.n79 B.n78 585
R1283 B.n894 B.n893 585
R1284 B.n893 B.n892 585
R1285 B.n81 B.n80 585
R1286 B.n891 B.n81 585
R1287 B.n889 B.n888 585
R1288 B.n890 B.n889 585
R1289 B.n887 B.n86 585
R1290 B.n86 B.n85 585
R1291 B.n886 B.n885 585
R1292 B.n885 B.n884 585
R1293 B.n982 B.n981 585
R1294 B.n981 B.n980 585
R1295 B.n676 B.n425 530.939
R1296 B.n885 B.n88 530.939
R1297 B.n674 B.n427 530.939
R1298 B.n882 B.n89 530.939
R1299 B.n450 B.t16 360.824
R1300 B.n139 B.t8 360.824
R1301 B.n456 B.t19 360.824
R1302 B.n141 B.t11 360.824
R1303 B.n450 B.t13 308.673
R1304 B.n456 B.t17 308.673
R1305 B.n141 B.t10 308.673
R1306 B.n139 B.t6 308.673
R1307 B.n451 B.t15 294.885
R1308 B.n140 B.t9 294.885
R1309 B.n457 B.t18 294.885
R1310 B.n142 B.t12 294.885
R1311 B.n883 B.n137 256.663
R1312 B.n883 B.n136 256.663
R1313 B.n883 B.n135 256.663
R1314 B.n883 B.n134 256.663
R1315 B.n883 B.n133 256.663
R1316 B.n883 B.n132 256.663
R1317 B.n883 B.n131 256.663
R1318 B.n883 B.n130 256.663
R1319 B.n883 B.n129 256.663
R1320 B.n883 B.n128 256.663
R1321 B.n883 B.n127 256.663
R1322 B.n883 B.n126 256.663
R1323 B.n883 B.n125 256.663
R1324 B.n883 B.n124 256.663
R1325 B.n883 B.n123 256.663
R1326 B.n883 B.n122 256.663
R1327 B.n883 B.n121 256.663
R1328 B.n883 B.n120 256.663
R1329 B.n883 B.n119 256.663
R1330 B.n883 B.n118 256.663
R1331 B.n883 B.n117 256.663
R1332 B.n883 B.n116 256.663
R1333 B.n883 B.n115 256.663
R1334 B.n883 B.n114 256.663
R1335 B.n883 B.n113 256.663
R1336 B.n883 B.n112 256.663
R1337 B.n883 B.n111 256.663
R1338 B.n883 B.n110 256.663
R1339 B.n883 B.n109 256.663
R1340 B.n883 B.n108 256.663
R1341 B.n883 B.n107 256.663
R1342 B.n883 B.n106 256.663
R1343 B.n883 B.n105 256.663
R1344 B.n883 B.n104 256.663
R1345 B.n883 B.n103 256.663
R1346 B.n883 B.n102 256.663
R1347 B.n883 B.n101 256.663
R1348 B.n883 B.n100 256.663
R1349 B.n883 B.n99 256.663
R1350 B.n883 B.n98 256.663
R1351 B.n883 B.n97 256.663
R1352 B.n883 B.n96 256.663
R1353 B.n883 B.n95 256.663
R1354 B.n883 B.n94 256.663
R1355 B.n883 B.n93 256.663
R1356 B.n883 B.n92 256.663
R1357 B.n883 B.n91 256.663
R1358 B.n883 B.n90 256.663
R1359 B.n480 B.n426 256.663
R1360 B.n483 B.n426 256.663
R1361 B.n489 B.n426 256.663
R1362 B.n491 B.n426 256.663
R1363 B.n497 B.n426 256.663
R1364 B.n499 B.n426 256.663
R1365 B.n505 B.n426 256.663
R1366 B.n507 B.n426 256.663
R1367 B.n513 B.n426 256.663
R1368 B.n515 B.n426 256.663
R1369 B.n521 B.n426 256.663
R1370 B.n523 B.n426 256.663
R1371 B.n529 B.n426 256.663
R1372 B.n531 B.n426 256.663
R1373 B.n537 B.n426 256.663
R1374 B.n539 B.n426 256.663
R1375 B.n545 B.n426 256.663
R1376 B.n547 B.n426 256.663
R1377 B.n553 B.n426 256.663
R1378 B.n555 B.n426 256.663
R1379 B.n561 B.n426 256.663
R1380 B.n563 B.n426 256.663
R1381 B.n570 B.n426 256.663
R1382 B.n572 B.n426 256.663
R1383 B.n578 B.n426 256.663
R1384 B.n580 B.n426 256.663
R1385 B.n587 B.n426 256.663
R1386 B.n589 B.n426 256.663
R1387 B.n595 B.n426 256.663
R1388 B.n597 B.n426 256.663
R1389 B.n603 B.n426 256.663
R1390 B.n605 B.n426 256.663
R1391 B.n611 B.n426 256.663
R1392 B.n613 B.n426 256.663
R1393 B.n619 B.n426 256.663
R1394 B.n621 B.n426 256.663
R1395 B.n627 B.n426 256.663
R1396 B.n629 B.n426 256.663
R1397 B.n635 B.n426 256.663
R1398 B.n637 B.n426 256.663
R1399 B.n643 B.n426 256.663
R1400 B.n645 B.n426 256.663
R1401 B.n651 B.n426 256.663
R1402 B.n653 B.n426 256.663
R1403 B.n659 B.n426 256.663
R1404 B.n661 B.n426 256.663
R1405 B.n667 B.n426 256.663
R1406 B.n669 B.n426 256.663
R1407 B.n676 B.n423 163.367
R1408 B.n680 B.n423 163.367
R1409 B.n680 B.n417 163.367
R1410 B.n688 B.n417 163.367
R1411 B.n688 B.n415 163.367
R1412 B.n692 B.n415 163.367
R1413 B.n692 B.n409 163.367
R1414 B.n700 B.n409 163.367
R1415 B.n700 B.n407 163.367
R1416 B.n704 B.n407 163.367
R1417 B.n704 B.n401 163.367
R1418 B.n712 B.n401 163.367
R1419 B.n712 B.n399 163.367
R1420 B.n716 B.n399 163.367
R1421 B.n716 B.n393 163.367
R1422 B.n724 B.n393 163.367
R1423 B.n724 B.n391 163.367
R1424 B.n728 B.n391 163.367
R1425 B.n728 B.n385 163.367
R1426 B.n737 B.n385 163.367
R1427 B.n737 B.n383 163.367
R1428 B.n741 B.n383 163.367
R1429 B.n741 B.n378 163.367
R1430 B.n749 B.n378 163.367
R1431 B.n749 B.n376 163.367
R1432 B.n753 B.n376 163.367
R1433 B.n753 B.n370 163.367
R1434 B.n761 B.n370 163.367
R1435 B.n761 B.n368 163.367
R1436 B.n765 B.n368 163.367
R1437 B.n765 B.n362 163.367
R1438 B.n773 B.n362 163.367
R1439 B.n773 B.n360 163.367
R1440 B.n777 B.n360 163.367
R1441 B.n777 B.n354 163.367
R1442 B.n785 B.n354 163.367
R1443 B.n785 B.n352 163.367
R1444 B.n789 B.n352 163.367
R1445 B.n789 B.n346 163.367
R1446 B.n798 B.n346 163.367
R1447 B.n798 B.n344 163.367
R1448 B.n802 B.n344 163.367
R1449 B.n802 B.n339 163.367
R1450 B.n811 B.n339 163.367
R1451 B.n811 B.n337 163.367
R1452 B.n815 B.n337 163.367
R1453 B.n815 B.n2 163.367
R1454 B.n981 B.n2 163.367
R1455 B.n981 B.n3 163.367
R1456 B.n977 B.n3 163.367
R1457 B.n977 B.n9 163.367
R1458 B.n973 B.n9 163.367
R1459 B.n973 B.n11 163.367
R1460 B.n969 B.n11 163.367
R1461 B.n969 B.n15 163.367
R1462 B.n965 B.n15 163.367
R1463 B.n965 B.n17 163.367
R1464 B.n961 B.n17 163.367
R1465 B.n961 B.n23 163.367
R1466 B.n957 B.n23 163.367
R1467 B.n957 B.n25 163.367
R1468 B.n953 B.n25 163.367
R1469 B.n953 B.n30 163.367
R1470 B.n949 B.n30 163.367
R1471 B.n949 B.n32 163.367
R1472 B.n945 B.n32 163.367
R1473 B.n945 B.n37 163.367
R1474 B.n941 B.n37 163.367
R1475 B.n941 B.n39 163.367
R1476 B.n937 B.n39 163.367
R1477 B.n937 B.n44 163.367
R1478 B.n933 B.n44 163.367
R1479 B.n933 B.n46 163.367
R1480 B.n929 B.n46 163.367
R1481 B.n929 B.n50 163.367
R1482 B.n925 B.n50 163.367
R1483 B.n925 B.n52 163.367
R1484 B.n921 B.n52 163.367
R1485 B.n921 B.n58 163.367
R1486 B.n917 B.n58 163.367
R1487 B.n917 B.n60 163.367
R1488 B.n913 B.n60 163.367
R1489 B.n913 B.n65 163.367
R1490 B.n909 B.n65 163.367
R1491 B.n909 B.n67 163.367
R1492 B.n905 B.n67 163.367
R1493 B.n905 B.n72 163.367
R1494 B.n901 B.n72 163.367
R1495 B.n901 B.n74 163.367
R1496 B.n897 B.n74 163.367
R1497 B.n897 B.n79 163.367
R1498 B.n893 B.n79 163.367
R1499 B.n893 B.n81 163.367
R1500 B.n889 B.n81 163.367
R1501 B.n889 B.n86 163.367
R1502 B.n885 B.n86 163.367
R1503 B.n482 B.n481 163.367
R1504 B.n484 B.n482 163.367
R1505 B.n488 B.n477 163.367
R1506 B.n492 B.n490 163.367
R1507 B.n496 B.n475 163.367
R1508 B.n500 B.n498 163.367
R1509 B.n504 B.n473 163.367
R1510 B.n508 B.n506 163.367
R1511 B.n512 B.n471 163.367
R1512 B.n516 B.n514 163.367
R1513 B.n520 B.n469 163.367
R1514 B.n524 B.n522 163.367
R1515 B.n528 B.n467 163.367
R1516 B.n532 B.n530 163.367
R1517 B.n536 B.n465 163.367
R1518 B.n540 B.n538 163.367
R1519 B.n544 B.n463 163.367
R1520 B.n548 B.n546 163.367
R1521 B.n552 B.n461 163.367
R1522 B.n556 B.n554 163.367
R1523 B.n560 B.n459 163.367
R1524 B.n564 B.n562 163.367
R1525 B.n569 B.n455 163.367
R1526 B.n573 B.n571 163.367
R1527 B.n577 B.n453 163.367
R1528 B.n581 B.n579 163.367
R1529 B.n586 B.n449 163.367
R1530 B.n590 B.n588 163.367
R1531 B.n594 B.n447 163.367
R1532 B.n598 B.n596 163.367
R1533 B.n602 B.n445 163.367
R1534 B.n606 B.n604 163.367
R1535 B.n610 B.n443 163.367
R1536 B.n614 B.n612 163.367
R1537 B.n618 B.n441 163.367
R1538 B.n622 B.n620 163.367
R1539 B.n626 B.n439 163.367
R1540 B.n630 B.n628 163.367
R1541 B.n634 B.n437 163.367
R1542 B.n638 B.n636 163.367
R1543 B.n642 B.n435 163.367
R1544 B.n646 B.n644 163.367
R1545 B.n650 B.n433 163.367
R1546 B.n654 B.n652 163.367
R1547 B.n658 B.n431 163.367
R1548 B.n662 B.n660 163.367
R1549 B.n666 B.n429 163.367
R1550 B.n670 B.n668 163.367
R1551 B.n674 B.n421 163.367
R1552 B.n682 B.n421 163.367
R1553 B.n682 B.n419 163.367
R1554 B.n686 B.n419 163.367
R1555 B.n686 B.n413 163.367
R1556 B.n694 B.n413 163.367
R1557 B.n694 B.n411 163.367
R1558 B.n698 B.n411 163.367
R1559 B.n698 B.n405 163.367
R1560 B.n706 B.n405 163.367
R1561 B.n706 B.n403 163.367
R1562 B.n710 B.n403 163.367
R1563 B.n710 B.n397 163.367
R1564 B.n718 B.n397 163.367
R1565 B.n718 B.n395 163.367
R1566 B.n722 B.n395 163.367
R1567 B.n722 B.n389 163.367
R1568 B.n730 B.n389 163.367
R1569 B.n730 B.n387 163.367
R1570 B.n734 B.n387 163.367
R1571 B.n734 B.n382 163.367
R1572 B.n743 B.n382 163.367
R1573 B.n743 B.n380 163.367
R1574 B.n747 B.n380 163.367
R1575 B.n747 B.n374 163.367
R1576 B.n755 B.n374 163.367
R1577 B.n755 B.n372 163.367
R1578 B.n759 B.n372 163.367
R1579 B.n759 B.n365 163.367
R1580 B.n767 B.n365 163.367
R1581 B.n767 B.n363 163.367
R1582 B.n771 B.n363 163.367
R1583 B.n771 B.n358 163.367
R1584 B.n779 B.n358 163.367
R1585 B.n779 B.n356 163.367
R1586 B.n783 B.n356 163.367
R1587 B.n783 B.n350 163.367
R1588 B.n791 B.n350 163.367
R1589 B.n791 B.n348 163.367
R1590 B.n795 B.n348 163.367
R1591 B.n795 B.n343 163.367
R1592 B.n804 B.n343 163.367
R1593 B.n804 B.n341 163.367
R1594 B.n809 B.n341 163.367
R1595 B.n809 B.n335 163.367
R1596 B.n817 B.n335 163.367
R1597 B.n818 B.n817 163.367
R1598 B.n818 B.n5 163.367
R1599 B.n6 B.n5 163.367
R1600 B.n7 B.n6 163.367
R1601 B.n823 B.n7 163.367
R1602 B.n823 B.n12 163.367
R1603 B.n13 B.n12 163.367
R1604 B.n14 B.n13 163.367
R1605 B.n828 B.n14 163.367
R1606 B.n828 B.n19 163.367
R1607 B.n20 B.n19 163.367
R1608 B.n21 B.n20 163.367
R1609 B.n833 B.n21 163.367
R1610 B.n833 B.n26 163.367
R1611 B.n27 B.n26 163.367
R1612 B.n28 B.n27 163.367
R1613 B.n838 B.n28 163.367
R1614 B.n838 B.n33 163.367
R1615 B.n34 B.n33 163.367
R1616 B.n35 B.n34 163.367
R1617 B.n843 B.n35 163.367
R1618 B.n843 B.n40 163.367
R1619 B.n41 B.n40 163.367
R1620 B.n42 B.n41 163.367
R1621 B.n848 B.n42 163.367
R1622 B.n848 B.n47 163.367
R1623 B.n48 B.n47 163.367
R1624 B.n49 B.n48 163.367
R1625 B.n853 B.n49 163.367
R1626 B.n853 B.n54 163.367
R1627 B.n55 B.n54 163.367
R1628 B.n56 B.n55 163.367
R1629 B.n858 B.n56 163.367
R1630 B.n858 B.n61 163.367
R1631 B.n62 B.n61 163.367
R1632 B.n63 B.n62 163.367
R1633 B.n863 B.n63 163.367
R1634 B.n863 B.n68 163.367
R1635 B.n69 B.n68 163.367
R1636 B.n70 B.n69 163.367
R1637 B.n868 B.n70 163.367
R1638 B.n868 B.n75 163.367
R1639 B.n76 B.n75 163.367
R1640 B.n77 B.n76 163.367
R1641 B.n873 B.n77 163.367
R1642 B.n873 B.n82 163.367
R1643 B.n83 B.n82 163.367
R1644 B.n84 B.n83 163.367
R1645 B.n878 B.n84 163.367
R1646 B.n878 B.n89 163.367
R1647 B.n146 B.n145 163.367
R1648 B.n150 B.n149 163.367
R1649 B.n154 B.n153 163.367
R1650 B.n158 B.n157 163.367
R1651 B.n162 B.n161 163.367
R1652 B.n166 B.n165 163.367
R1653 B.n170 B.n169 163.367
R1654 B.n174 B.n173 163.367
R1655 B.n178 B.n177 163.367
R1656 B.n182 B.n181 163.367
R1657 B.n186 B.n185 163.367
R1658 B.n190 B.n189 163.367
R1659 B.n194 B.n193 163.367
R1660 B.n198 B.n197 163.367
R1661 B.n202 B.n201 163.367
R1662 B.n206 B.n205 163.367
R1663 B.n210 B.n209 163.367
R1664 B.n214 B.n213 163.367
R1665 B.n218 B.n217 163.367
R1666 B.n222 B.n221 163.367
R1667 B.n226 B.n225 163.367
R1668 B.n230 B.n229 163.367
R1669 B.n234 B.n233 163.367
R1670 B.n238 B.n237 163.367
R1671 B.n242 B.n241 163.367
R1672 B.n246 B.n245 163.367
R1673 B.n251 B.n250 163.367
R1674 B.n255 B.n254 163.367
R1675 B.n259 B.n258 163.367
R1676 B.n263 B.n262 163.367
R1677 B.n267 B.n266 163.367
R1678 B.n271 B.n270 163.367
R1679 B.n275 B.n274 163.367
R1680 B.n279 B.n278 163.367
R1681 B.n283 B.n282 163.367
R1682 B.n287 B.n286 163.367
R1683 B.n291 B.n290 163.367
R1684 B.n295 B.n294 163.367
R1685 B.n299 B.n298 163.367
R1686 B.n303 B.n302 163.367
R1687 B.n307 B.n306 163.367
R1688 B.n311 B.n310 163.367
R1689 B.n315 B.n314 163.367
R1690 B.n319 B.n318 163.367
R1691 B.n323 B.n322 163.367
R1692 B.n327 B.n326 163.367
R1693 B.n331 B.n330 163.367
R1694 B.n882 B.n138 163.367
R1695 B.n675 B.n426 79.9894
R1696 B.n884 B.n883 79.9894
R1697 B.n480 B.n425 71.676
R1698 B.n484 B.n483 71.676
R1699 B.n489 B.n488 71.676
R1700 B.n492 B.n491 71.676
R1701 B.n497 B.n496 71.676
R1702 B.n500 B.n499 71.676
R1703 B.n505 B.n504 71.676
R1704 B.n508 B.n507 71.676
R1705 B.n513 B.n512 71.676
R1706 B.n516 B.n515 71.676
R1707 B.n521 B.n520 71.676
R1708 B.n524 B.n523 71.676
R1709 B.n529 B.n528 71.676
R1710 B.n532 B.n531 71.676
R1711 B.n537 B.n536 71.676
R1712 B.n540 B.n539 71.676
R1713 B.n545 B.n544 71.676
R1714 B.n548 B.n547 71.676
R1715 B.n553 B.n552 71.676
R1716 B.n556 B.n555 71.676
R1717 B.n561 B.n560 71.676
R1718 B.n564 B.n563 71.676
R1719 B.n570 B.n569 71.676
R1720 B.n573 B.n572 71.676
R1721 B.n578 B.n577 71.676
R1722 B.n581 B.n580 71.676
R1723 B.n587 B.n586 71.676
R1724 B.n590 B.n589 71.676
R1725 B.n595 B.n594 71.676
R1726 B.n598 B.n597 71.676
R1727 B.n603 B.n602 71.676
R1728 B.n606 B.n605 71.676
R1729 B.n611 B.n610 71.676
R1730 B.n614 B.n613 71.676
R1731 B.n619 B.n618 71.676
R1732 B.n622 B.n621 71.676
R1733 B.n627 B.n626 71.676
R1734 B.n630 B.n629 71.676
R1735 B.n635 B.n634 71.676
R1736 B.n638 B.n637 71.676
R1737 B.n643 B.n642 71.676
R1738 B.n646 B.n645 71.676
R1739 B.n651 B.n650 71.676
R1740 B.n654 B.n653 71.676
R1741 B.n659 B.n658 71.676
R1742 B.n662 B.n661 71.676
R1743 B.n667 B.n666 71.676
R1744 B.n670 B.n669 71.676
R1745 B.n90 B.n88 71.676
R1746 B.n146 B.n91 71.676
R1747 B.n150 B.n92 71.676
R1748 B.n154 B.n93 71.676
R1749 B.n158 B.n94 71.676
R1750 B.n162 B.n95 71.676
R1751 B.n166 B.n96 71.676
R1752 B.n170 B.n97 71.676
R1753 B.n174 B.n98 71.676
R1754 B.n178 B.n99 71.676
R1755 B.n182 B.n100 71.676
R1756 B.n186 B.n101 71.676
R1757 B.n190 B.n102 71.676
R1758 B.n194 B.n103 71.676
R1759 B.n198 B.n104 71.676
R1760 B.n202 B.n105 71.676
R1761 B.n206 B.n106 71.676
R1762 B.n210 B.n107 71.676
R1763 B.n214 B.n108 71.676
R1764 B.n218 B.n109 71.676
R1765 B.n222 B.n110 71.676
R1766 B.n226 B.n111 71.676
R1767 B.n230 B.n112 71.676
R1768 B.n234 B.n113 71.676
R1769 B.n238 B.n114 71.676
R1770 B.n242 B.n115 71.676
R1771 B.n246 B.n116 71.676
R1772 B.n251 B.n117 71.676
R1773 B.n255 B.n118 71.676
R1774 B.n259 B.n119 71.676
R1775 B.n263 B.n120 71.676
R1776 B.n267 B.n121 71.676
R1777 B.n271 B.n122 71.676
R1778 B.n275 B.n123 71.676
R1779 B.n279 B.n124 71.676
R1780 B.n283 B.n125 71.676
R1781 B.n287 B.n126 71.676
R1782 B.n291 B.n127 71.676
R1783 B.n295 B.n128 71.676
R1784 B.n299 B.n129 71.676
R1785 B.n303 B.n130 71.676
R1786 B.n307 B.n131 71.676
R1787 B.n311 B.n132 71.676
R1788 B.n315 B.n133 71.676
R1789 B.n319 B.n134 71.676
R1790 B.n323 B.n135 71.676
R1791 B.n327 B.n136 71.676
R1792 B.n331 B.n137 71.676
R1793 B.n138 B.n137 71.676
R1794 B.n330 B.n136 71.676
R1795 B.n326 B.n135 71.676
R1796 B.n322 B.n134 71.676
R1797 B.n318 B.n133 71.676
R1798 B.n314 B.n132 71.676
R1799 B.n310 B.n131 71.676
R1800 B.n306 B.n130 71.676
R1801 B.n302 B.n129 71.676
R1802 B.n298 B.n128 71.676
R1803 B.n294 B.n127 71.676
R1804 B.n290 B.n126 71.676
R1805 B.n286 B.n125 71.676
R1806 B.n282 B.n124 71.676
R1807 B.n278 B.n123 71.676
R1808 B.n274 B.n122 71.676
R1809 B.n270 B.n121 71.676
R1810 B.n266 B.n120 71.676
R1811 B.n262 B.n119 71.676
R1812 B.n258 B.n118 71.676
R1813 B.n254 B.n117 71.676
R1814 B.n250 B.n116 71.676
R1815 B.n245 B.n115 71.676
R1816 B.n241 B.n114 71.676
R1817 B.n237 B.n113 71.676
R1818 B.n233 B.n112 71.676
R1819 B.n229 B.n111 71.676
R1820 B.n225 B.n110 71.676
R1821 B.n221 B.n109 71.676
R1822 B.n217 B.n108 71.676
R1823 B.n213 B.n107 71.676
R1824 B.n209 B.n106 71.676
R1825 B.n205 B.n105 71.676
R1826 B.n201 B.n104 71.676
R1827 B.n197 B.n103 71.676
R1828 B.n193 B.n102 71.676
R1829 B.n189 B.n101 71.676
R1830 B.n185 B.n100 71.676
R1831 B.n181 B.n99 71.676
R1832 B.n177 B.n98 71.676
R1833 B.n173 B.n97 71.676
R1834 B.n169 B.n96 71.676
R1835 B.n165 B.n95 71.676
R1836 B.n161 B.n94 71.676
R1837 B.n157 B.n93 71.676
R1838 B.n153 B.n92 71.676
R1839 B.n149 B.n91 71.676
R1840 B.n145 B.n90 71.676
R1841 B.n481 B.n480 71.676
R1842 B.n483 B.n477 71.676
R1843 B.n490 B.n489 71.676
R1844 B.n491 B.n475 71.676
R1845 B.n498 B.n497 71.676
R1846 B.n499 B.n473 71.676
R1847 B.n506 B.n505 71.676
R1848 B.n507 B.n471 71.676
R1849 B.n514 B.n513 71.676
R1850 B.n515 B.n469 71.676
R1851 B.n522 B.n521 71.676
R1852 B.n523 B.n467 71.676
R1853 B.n530 B.n529 71.676
R1854 B.n531 B.n465 71.676
R1855 B.n538 B.n537 71.676
R1856 B.n539 B.n463 71.676
R1857 B.n546 B.n545 71.676
R1858 B.n547 B.n461 71.676
R1859 B.n554 B.n553 71.676
R1860 B.n555 B.n459 71.676
R1861 B.n562 B.n561 71.676
R1862 B.n563 B.n455 71.676
R1863 B.n571 B.n570 71.676
R1864 B.n572 B.n453 71.676
R1865 B.n579 B.n578 71.676
R1866 B.n580 B.n449 71.676
R1867 B.n588 B.n587 71.676
R1868 B.n589 B.n447 71.676
R1869 B.n596 B.n595 71.676
R1870 B.n597 B.n445 71.676
R1871 B.n604 B.n603 71.676
R1872 B.n605 B.n443 71.676
R1873 B.n612 B.n611 71.676
R1874 B.n613 B.n441 71.676
R1875 B.n620 B.n619 71.676
R1876 B.n621 B.n439 71.676
R1877 B.n628 B.n627 71.676
R1878 B.n629 B.n437 71.676
R1879 B.n636 B.n635 71.676
R1880 B.n637 B.n435 71.676
R1881 B.n644 B.n643 71.676
R1882 B.n645 B.n433 71.676
R1883 B.n652 B.n651 71.676
R1884 B.n653 B.n431 71.676
R1885 B.n660 B.n659 71.676
R1886 B.n661 B.n429 71.676
R1887 B.n668 B.n667 71.676
R1888 B.n669 B.n427 71.676
R1889 B.n451 B.n450 65.9399
R1890 B.n457 B.n456 65.9399
R1891 B.n142 B.n141 65.9399
R1892 B.n140 B.n139 65.9399
R1893 B.n584 B.n451 59.5399
R1894 B.n566 B.n457 59.5399
R1895 B.n143 B.n142 59.5399
R1896 B.n248 B.n140 59.5399
R1897 B.n675 B.n422 41.5215
R1898 B.n681 B.n422 41.5215
R1899 B.n681 B.n418 41.5215
R1900 B.n687 B.n418 41.5215
R1901 B.n687 B.n414 41.5215
R1902 B.n693 B.n414 41.5215
R1903 B.n693 B.n410 41.5215
R1904 B.n699 B.n410 41.5215
R1905 B.n705 B.n406 41.5215
R1906 B.n705 B.n402 41.5215
R1907 B.n711 B.n402 41.5215
R1908 B.n711 B.n398 41.5215
R1909 B.n717 B.n398 41.5215
R1910 B.n717 B.n394 41.5215
R1911 B.n723 B.n394 41.5215
R1912 B.n723 B.n390 41.5215
R1913 B.n729 B.n390 41.5215
R1914 B.n729 B.n386 41.5215
R1915 B.n736 B.n386 41.5215
R1916 B.n736 B.n735 41.5215
R1917 B.n742 B.n379 41.5215
R1918 B.n748 B.n379 41.5215
R1919 B.n748 B.n375 41.5215
R1920 B.n754 B.n375 41.5215
R1921 B.n754 B.n371 41.5215
R1922 B.n760 B.n371 41.5215
R1923 B.n760 B.n366 41.5215
R1924 B.n766 B.n366 41.5215
R1925 B.n766 B.n367 41.5215
R1926 B.n772 B.n359 41.5215
R1927 B.n778 B.n359 41.5215
R1928 B.n778 B.n355 41.5215
R1929 B.n784 B.n355 41.5215
R1930 B.n784 B.n351 41.5215
R1931 B.n790 B.n351 41.5215
R1932 B.n790 B.n347 41.5215
R1933 B.n797 B.n347 41.5215
R1934 B.n797 B.n796 41.5215
R1935 B.n803 B.n340 41.5215
R1936 B.n810 B.n340 41.5215
R1937 B.n810 B.n336 41.5215
R1938 B.n816 B.n336 41.5215
R1939 B.n816 B.n4 41.5215
R1940 B.n980 B.n4 41.5215
R1941 B.n980 B.n979 41.5215
R1942 B.n979 B.n978 41.5215
R1943 B.n978 B.n8 41.5215
R1944 B.n972 B.n8 41.5215
R1945 B.n972 B.n971 41.5215
R1946 B.n971 B.n970 41.5215
R1947 B.n964 B.n18 41.5215
R1948 B.n964 B.n963 41.5215
R1949 B.n963 B.n962 41.5215
R1950 B.n962 B.n22 41.5215
R1951 B.n956 B.n22 41.5215
R1952 B.n956 B.n955 41.5215
R1953 B.n955 B.n954 41.5215
R1954 B.n954 B.n29 41.5215
R1955 B.n948 B.n29 41.5215
R1956 B.n947 B.n946 41.5215
R1957 B.n946 B.n36 41.5215
R1958 B.n940 B.n36 41.5215
R1959 B.n940 B.n939 41.5215
R1960 B.n939 B.n938 41.5215
R1961 B.n938 B.n43 41.5215
R1962 B.n932 B.n43 41.5215
R1963 B.n932 B.n931 41.5215
R1964 B.n931 B.n930 41.5215
R1965 B.n924 B.n53 41.5215
R1966 B.n924 B.n923 41.5215
R1967 B.n923 B.n922 41.5215
R1968 B.n922 B.n57 41.5215
R1969 B.n916 B.n57 41.5215
R1970 B.n916 B.n915 41.5215
R1971 B.n915 B.n914 41.5215
R1972 B.n914 B.n64 41.5215
R1973 B.n908 B.n64 41.5215
R1974 B.n908 B.n907 41.5215
R1975 B.n907 B.n906 41.5215
R1976 B.n906 B.n71 41.5215
R1977 B.n900 B.n899 41.5215
R1978 B.n899 B.n898 41.5215
R1979 B.n898 B.n78 41.5215
R1980 B.n892 B.n78 41.5215
R1981 B.n892 B.n891 41.5215
R1982 B.n891 B.n890 41.5215
R1983 B.n890 B.n85 41.5215
R1984 B.n884 B.n85 41.5215
R1985 B.n886 B.n87 34.4981
R1986 B.n881 B.n880 34.4981
R1987 B.n673 B.n672 34.4981
R1988 B.n677 B.n424 34.4981
R1989 B.t14 B.n406 33.5836
R1990 B.t7 B.n71 33.5836
R1991 B.n742 B.t1 25.0352
R1992 B.n772 B.t0 25.0352
R1993 B.n803 B.t3 25.0352
R1994 B.n970 B.t2 25.0352
R1995 B.n948 B.t5 25.0352
R1996 B.n930 B.t4 25.0352
R1997 B B.n982 18.0485
R1998 B.n735 B.t1 16.4868
R1999 B.n367 B.t0 16.4868
R2000 B.n796 B.t3 16.4868
R2001 B.n18 B.t2 16.4868
R2002 B.t5 B.n947 16.4868
R2003 B.n53 B.t4 16.4868
R2004 B.n144 B.n87 10.6151
R2005 B.n147 B.n144 10.6151
R2006 B.n148 B.n147 10.6151
R2007 B.n151 B.n148 10.6151
R2008 B.n152 B.n151 10.6151
R2009 B.n155 B.n152 10.6151
R2010 B.n156 B.n155 10.6151
R2011 B.n159 B.n156 10.6151
R2012 B.n160 B.n159 10.6151
R2013 B.n163 B.n160 10.6151
R2014 B.n164 B.n163 10.6151
R2015 B.n167 B.n164 10.6151
R2016 B.n168 B.n167 10.6151
R2017 B.n171 B.n168 10.6151
R2018 B.n172 B.n171 10.6151
R2019 B.n175 B.n172 10.6151
R2020 B.n176 B.n175 10.6151
R2021 B.n179 B.n176 10.6151
R2022 B.n180 B.n179 10.6151
R2023 B.n183 B.n180 10.6151
R2024 B.n184 B.n183 10.6151
R2025 B.n187 B.n184 10.6151
R2026 B.n188 B.n187 10.6151
R2027 B.n191 B.n188 10.6151
R2028 B.n192 B.n191 10.6151
R2029 B.n195 B.n192 10.6151
R2030 B.n196 B.n195 10.6151
R2031 B.n199 B.n196 10.6151
R2032 B.n200 B.n199 10.6151
R2033 B.n203 B.n200 10.6151
R2034 B.n204 B.n203 10.6151
R2035 B.n207 B.n204 10.6151
R2036 B.n208 B.n207 10.6151
R2037 B.n211 B.n208 10.6151
R2038 B.n212 B.n211 10.6151
R2039 B.n215 B.n212 10.6151
R2040 B.n216 B.n215 10.6151
R2041 B.n219 B.n216 10.6151
R2042 B.n220 B.n219 10.6151
R2043 B.n223 B.n220 10.6151
R2044 B.n224 B.n223 10.6151
R2045 B.n227 B.n224 10.6151
R2046 B.n228 B.n227 10.6151
R2047 B.n232 B.n231 10.6151
R2048 B.n235 B.n232 10.6151
R2049 B.n236 B.n235 10.6151
R2050 B.n239 B.n236 10.6151
R2051 B.n240 B.n239 10.6151
R2052 B.n243 B.n240 10.6151
R2053 B.n244 B.n243 10.6151
R2054 B.n247 B.n244 10.6151
R2055 B.n252 B.n249 10.6151
R2056 B.n253 B.n252 10.6151
R2057 B.n256 B.n253 10.6151
R2058 B.n257 B.n256 10.6151
R2059 B.n260 B.n257 10.6151
R2060 B.n261 B.n260 10.6151
R2061 B.n264 B.n261 10.6151
R2062 B.n265 B.n264 10.6151
R2063 B.n268 B.n265 10.6151
R2064 B.n269 B.n268 10.6151
R2065 B.n272 B.n269 10.6151
R2066 B.n273 B.n272 10.6151
R2067 B.n276 B.n273 10.6151
R2068 B.n277 B.n276 10.6151
R2069 B.n280 B.n277 10.6151
R2070 B.n281 B.n280 10.6151
R2071 B.n284 B.n281 10.6151
R2072 B.n285 B.n284 10.6151
R2073 B.n288 B.n285 10.6151
R2074 B.n289 B.n288 10.6151
R2075 B.n292 B.n289 10.6151
R2076 B.n293 B.n292 10.6151
R2077 B.n296 B.n293 10.6151
R2078 B.n297 B.n296 10.6151
R2079 B.n300 B.n297 10.6151
R2080 B.n301 B.n300 10.6151
R2081 B.n304 B.n301 10.6151
R2082 B.n305 B.n304 10.6151
R2083 B.n308 B.n305 10.6151
R2084 B.n309 B.n308 10.6151
R2085 B.n312 B.n309 10.6151
R2086 B.n313 B.n312 10.6151
R2087 B.n316 B.n313 10.6151
R2088 B.n317 B.n316 10.6151
R2089 B.n320 B.n317 10.6151
R2090 B.n321 B.n320 10.6151
R2091 B.n324 B.n321 10.6151
R2092 B.n325 B.n324 10.6151
R2093 B.n328 B.n325 10.6151
R2094 B.n329 B.n328 10.6151
R2095 B.n332 B.n329 10.6151
R2096 B.n333 B.n332 10.6151
R2097 B.n881 B.n333 10.6151
R2098 B.n673 B.n420 10.6151
R2099 B.n683 B.n420 10.6151
R2100 B.n684 B.n683 10.6151
R2101 B.n685 B.n684 10.6151
R2102 B.n685 B.n412 10.6151
R2103 B.n695 B.n412 10.6151
R2104 B.n696 B.n695 10.6151
R2105 B.n697 B.n696 10.6151
R2106 B.n697 B.n404 10.6151
R2107 B.n707 B.n404 10.6151
R2108 B.n708 B.n707 10.6151
R2109 B.n709 B.n708 10.6151
R2110 B.n709 B.n396 10.6151
R2111 B.n719 B.n396 10.6151
R2112 B.n720 B.n719 10.6151
R2113 B.n721 B.n720 10.6151
R2114 B.n721 B.n388 10.6151
R2115 B.n731 B.n388 10.6151
R2116 B.n732 B.n731 10.6151
R2117 B.n733 B.n732 10.6151
R2118 B.n733 B.n381 10.6151
R2119 B.n744 B.n381 10.6151
R2120 B.n745 B.n744 10.6151
R2121 B.n746 B.n745 10.6151
R2122 B.n746 B.n373 10.6151
R2123 B.n756 B.n373 10.6151
R2124 B.n757 B.n756 10.6151
R2125 B.n758 B.n757 10.6151
R2126 B.n758 B.n364 10.6151
R2127 B.n768 B.n364 10.6151
R2128 B.n769 B.n768 10.6151
R2129 B.n770 B.n769 10.6151
R2130 B.n770 B.n357 10.6151
R2131 B.n780 B.n357 10.6151
R2132 B.n781 B.n780 10.6151
R2133 B.n782 B.n781 10.6151
R2134 B.n782 B.n349 10.6151
R2135 B.n792 B.n349 10.6151
R2136 B.n793 B.n792 10.6151
R2137 B.n794 B.n793 10.6151
R2138 B.n794 B.n342 10.6151
R2139 B.n805 B.n342 10.6151
R2140 B.n806 B.n805 10.6151
R2141 B.n808 B.n806 10.6151
R2142 B.n808 B.n807 10.6151
R2143 B.n807 B.n334 10.6151
R2144 B.n819 B.n334 10.6151
R2145 B.n820 B.n819 10.6151
R2146 B.n821 B.n820 10.6151
R2147 B.n822 B.n821 10.6151
R2148 B.n824 B.n822 10.6151
R2149 B.n825 B.n824 10.6151
R2150 B.n826 B.n825 10.6151
R2151 B.n827 B.n826 10.6151
R2152 B.n829 B.n827 10.6151
R2153 B.n830 B.n829 10.6151
R2154 B.n831 B.n830 10.6151
R2155 B.n832 B.n831 10.6151
R2156 B.n834 B.n832 10.6151
R2157 B.n835 B.n834 10.6151
R2158 B.n836 B.n835 10.6151
R2159 B.n837 B.n836 10.6151
R2160 B.n839 B.n837 10.6151
R2161 B.n840 B.n839 10.6151
R2162 B.n841 B.n840 10.6151
R2163 B.n842 B.n841 10.6151
R2164 B.n844 B.n842 10.6151
R2165 B.n845 B.n844 10.6151
R2166 B.n846 B.n845 10.6151
R2167 B.n847 B.n846 10.6151
R2168 B.n849 B.n847 10.6151
R2169 B.n850 B.n849 10.6151
R2170 B.n851 B.n850 10.6151
R2171 B.n852 B.n851 10.6151
R2172 B.n854 B.n852 10.6151
R2173 B.n855 B.n854 10.6151
R2174 B.n856 B.n855 10.6151
R2175 B.n857 B.n856 10.6151
R2176 B.n859 B.n857 10.6151
R2177 B.n860 B.n859 10.6151
R2178 B.n861 B.n860 10.6151
R2179 B.n862 B.n861 10.6151
R2180 B.n864 B.n862 10.6151
R2181 B.n865 B.n864 10.6151
R2182 B.n866 B.n865 10.6151
R2183 B.n867 B.n866 10.6151
R2184 B.n869 B.n867 10.6151
R2185 B.n870 B.n869 10.6151
R2186 B.n871 B.n870 10.6151
R2187 B.n872 B.n871 10.6151
R2188 B.n874 B.n872 10.6151
R2189 B.n875 B.n874 10.6151
R2190 B.n876 B.n875 10.6151
R2191 B.n877 B.n876 10.6151
R2192 B.n879 B.n877 10.6151
R2193 B.n880 B.n879 10.6151
R2194 B.n479 B.n424 10.6151
R2195 B.n479 B.n478 10.6151
R2196 B.n485 B.n478 10.6151
R2197 B.n486 B.n485 10.6151
R2198 B.n487 B.n486 10.6151
R2199 B.n487 B.n476 10.6151
R2200 B.n493 B.n476 10.6151
R2201 B.n494 B.n493 10.6151
R2202 B.n495 B.n494 10.6151
R2203 B.n495 B.n474 10.6151
R2204 B.n501 B.n474 10.6151
R2205 B.n502 B.n501 10.6151
R2206 B.n503 B.n502 10.6151
R2207 B.n503 B.n472 10.6151
R2208 B.n509 B.n472 10.6151
R2209 B.n510 B.n509 10.6151
R2210 B.n511 B.n510 10.6151
R2211 B.n511 B.n470 10.6151
R2212 B.n517 B.n470 10.6151
R2213 B.n518 B.n517 10.6151
R2214 B.n519 B.n518 10.6151
R2215 B.n519 B.n468 10.6151
R2216 B.n525 B.n468 10.6151
R2217 B.n526 B.n525 10.6151
R2218 B.n527 B.n526 10.6151
R2219 B.n527 B.n466 10.6151
R2220 B.n533 B.n466 10.6151
R2221 B.n534 B.n533 10.6151
R2222 B.n535 B.n534 10.6151
R2223 B.n535 B.n464 10.6151
R2224 B.n541 B.n464 10.6151
R2225 B.n542 B.n541 10.6151
R2226 B.n543 B.n542 10.6151
R2227 B.n543 B.n462 10.6151
R2228 B.n549 B.n462 10.6151
R2229 B.n550 B.n549 10.6151
R2230 B.n551 B.n550 10.6151
R2231 B.n551 B.n460 10.6151
R2232 B.n557 B.n460 10.6151
R2233 B.n558 B.n557 10.6151
R2234 B.n559 B.n558 10.6151
R2235 B.n559 B.n458 10.6151
R2236 B.n565 B.n458 10.6151
R2237 B.n568 B.n567 10.6151
R2238 B.n568 B.n454 10.6151
R2239 B.n574 B.n454 10.6151
R2240 B.n575 B.n574 10.6151
R2241 B.n576 B.n575 10.6151
R2242 B.n576 B.n452 10.6151
R2243 B.n582 B.n452 10.6151
R2244 B.n583 B.n582 10.6151
R2245 B.n585 B.n448 10.6151
R2246 B.n591 B.n448 10.6151
R2247 B.n592 B.n591 10.6151
R2248 B.n593 B.n592 10.6151
R2249 B.n593 B.n446 10.6151
R2250 B.n599 B.n446 10.6151
R2251 B.n600 B.n599 10.6151
R2252 B.n601 B.n600 10.6151
R2253 B.n601 B.n444 10.6151
R2254 B.n607 B.n444 10.6151
R2255 B.n608 B.n607 10.6151
R2256 B.n609 B.n608 10.6151
R2257 B.n609 B.n442 10.6151
R2258 B.n615 B.n442 10.6151
R2259 B.n616 B.n615 10.6151
R2260 B.n617 B.n616 10.6151
R2261 B.n617 B.n440 10.6151
R2262 B.n623 B.n440 10.6151
R2263 B.n624 B.n623 10.6151
R2264 B.n625 B.n624 10.6151
R2265 B.n625 B.n438 10.6151
R2266 B.n631 B.n438 10.6151
R2267 B.n632 B.n631 10.6151
R2268 B.n633 B.n632 10.6151
R2269 B.n633 B.n436 10.6151
R2270 B.n639 B.n436 10.6151
R2271 B.n640 B.n639 10.6151
R2272 B.n641 B.n640 10.6151
R2273 B.n641 B.n434 10.6151
R2274 B.n647 B.n434 10.6151
R2275 B.n648 B.n647 10.6151
R2276 B.n649 B.n648 10.6151
R2277 B.n649 B.n432 10.6151
R2278 B.n655 B.n432 10.6151
R2279 B.n656 B.n655 10.6151
R2280 B.n657 B.n656 10.6151
R2281 B.n657 B.n430 10.6151
R2282 B.n663 B.n430 10.6151
R2283 B.n664 B.n663 10.6151
R2284 B.n665 B.n664 10.6151
R2285 B.n665 B.n428 10.6151
R2286 B.n671 B.n428 10.6151
R2287 B.n672 B.n671 10.6151
R2288 B.n678 B.n677 10.6151
R2289 B.n679 B.n678 10.6151
R2290 B.n679 B.n416 10.6151
R2291 B.n689 B.n416 10.6151
R2292 B.n690 B.n689 10.6151
R2293 B.n691 B.n690 10.6151
R2294 B.n691 B.n408 10.6151
R2295 B.n701 B.n408 10.6151
R2296 B.n702 B.n701 10.6151
R2297 B.n703 B.n702 10.6151
R2298 B.n703 B.n400 10.6151
R2299 B.n713 B.n400 10.6151
R2300 B.n714 B.n713 10.6151
R2301 B.n715 B.n714 10.6151
R2302 B.n715 B.n392 10.6151
R2303 B.n725 B.n392 10.6151
R2304 B.n726 B.n725 10.6151
R2305 B.n727 B.n726 10.6151
R2306 B.n727 B.n384 10.6151
R2307 B.n738 B.n384 10.6151
R2308 B.n739 B.n738 10.6151
R2309 B.n740 B.n739 10.6151
R2310 B.n740 B.n377 10.6151
R2311 B.n750 B.n377 10.6151
R2312 B.n751 B.n750 10.6151
R2313 B.n752 B.n751 10.6151
R2314 B.n752 B.n369 10.6151
R2315 B.n762 B.n369 10.6151
R2316 B.n763 B.n762 10.6151
R2317 B.n764 B.n763 10.6151
R2318 B.n764 B.n361 10.6151
R2319 B.n774 B.n361 10.6151
R2320 B.n775 B.n774 10.6151
R2321 B.n776 B.n775 10.6151
R2322 B.n776 B.n353 10.6151
R2323 B.n786 B.n353 10.6151
R2324 B.n787 B.n786 10.6151
R2325 B.n788 B.n787 10.6151
R2326 B.n788 B.n345 10.6151
R2327 B.n799 B.n345 10.6151
R2328 B.n800 B.n799 10.6151
R2329 B.n801 B.n800 10.6151
R2330 B.n801 B.n338 10.6151
R2331 B.n812 B.n338 10.6151
R2332 B.n813 B.n812 10.6151
R2333 B.n814 B.n813 10.6151
R2334 B.n814 B.n0 10.6151
R2335 B.n976 B.n1 10.6151
R2336 B.n976 B.n975 10.6151
R2337 B.n975 B.n974 10.6151
R2338 B.n974 B.n10 10.6151
R2339 B.n968 B.n10 10.6151
R2340 B.n968 B.n967 10.6151
R2341 B.n967 B.n966 10.6151
R2342 B.n966 B.n16 10.6151
R2343 B.n960 B.n16 10.6151
R2344 B.n960 B.n959 10.6151
R2345 B.n959 B.n958 10.6151
R2346 B.n958 B.n24 10.6151
R2347 B.n952 B.n24 10.6151
R2348 B.n952 B.n951 10.6151
R2349 B.n951 B.n950 10.6151
R2350 B.n950 B.n31 10.6151
R2351 B.n944 B.n31 10.6151
R2352 B.n944 B.n943 10.6151
R2353 B.n943 B.n942 10.6151
R2354 B.n942 B.n38 10.6151
R2355 B.n936 B.n38 10.6151
R2356 B.n936 B.n935 10.6151
R2357 B.n935 B.n934 10.6151
R2358 B.n934 B.n45 10.6151
R2359 B.n928 B.n45 10.6151
R2360 B.n928 B.n927 10.6151
R2361 B.n927 B.n926 10.6151
R2362 B.n926 B.n51 10.6151
R2363 B.n920 B.n51 10.6151
R2364 B.n920 B.n919 10.6151
R2365 B.n919 B.n918 10.6151
R2366 B.n918 B.n59 10.6151
R2367 B.n912 B.n59 10.6151
R2368 B.n912 B.n911 10.6151
R2369 B.n911 B.n910 10.6151
R2370 B.n910 B.n66 10.6151
R2371 B.n904 B.n66 10.6151
R2372 B.n904 B.n903 10.6151
R2373 B.n903 B.n902 10.6151
R2374 B.n902 B.n73 10.6151
R2375 B.n896 B.n73 10.6151
R2376 B.n896 B.n895 10.6151
R2377 B.n895 B.n894 10.6151
R2378 B.n894 B.n80 10.6151
R2379 B.n888 B.n80 10.6151
R2380 B.n888 B.n887 10.6151
R2381 B.n887 B.n886 10.6151
R2382 B.n699 B.t14 7.93833
R2383 B.n900 B.t7 7.93833
R2384 B.n231 B.n143 6.5566
R2385 B.n248 B.n247 6.5566
R2386 B.n567 B.n566 6.5566
R2387 B.n584 B.n583 6.5566
R2388 B.n228 B.n143 4.05904
R2389 B.n249 B.n248 4.05904
R2390 B.n566 B.n565 4.05904
R2391 B.n585 B.n584 4.05904
R2392 B.n982 B.n0 2.81026
R2393 B.n982 B.n1 2.81026
R2394 VP.n13 VP.n10 161.3
R2395 VP.n15 VP.n14 161.3
R2396 VP.n16 VP.n9 161.3
R2397 VP.n18 VP.n17 161.3
R2398 VP.n19 VP.n8 161.3
R2399 VP.n21 VP.n20 161.3
R2400 VP.n44 VP.n43 161.3
R2401 VP.n42 VP.n1 161.3
R2402 VP.n41 VP.n40 161.3
R2403 VP.n39 VP.n2 161.3
R2404 VP.n38 VP.n37 161.3
R2405 VP.n36 VP.n3 161.3
R2406 VP.n35 VP.n34 161.3
R2407 VP.n33 VP.n4 161.3
R2408 VP.n32 VP.n31 161.3
R2409 VP.n30 VP.n5 161.3
R2410 VP.n29 VP.n28 161.3
R2411 VP.n27 VP.n6 161.3
R2412 VP.n26 VP.n25 161.3
R2413 VP.n11 VP.t1 133.321
R2414 VP.n35 VP.t5 100.011
R2415 VP.n24 VP.t3 100.011
R2416 VP.n0 VP.t0 100.011
R2417 VP.n12 VP.t2 100.011
R2418 VP.n7 VP.t4 100.011
R2419 VP.n24 VP.n23 70.4162
R2420 VP.n45 VP.n0 70.4162
R2421 VP.n22 VP.n7 70.4162
R2422 VP.n30 VP.n29 56.4773
R2423 VP.n41 VP.n2 56.4773
R2424 VP.n18 VP.n9 56.4773
R2425 VP.n23 VP.n22 51.2112
R2426 VP.n12 VP.n11 49.2698
R2427 VP.n25 VP.n6 24.3439
R2428 VP.n29 VP.n6 24.3439
R2429 VP.n31 VP.n30 24.3439
R2430 VP.n31 VP.n4 24.3439
R2431 VP.n35 VP.n4 24.3439
R2432 VP.n36 VP.n35 24.3439
R2433 VP.n37 VP.n36 24.3439
R2434 VP.n37 VP.n2 24.3439
R2435 VP.n42 VP.n41 24.3439
R2436 VP.n43 VP.n42 24.3439
R2437 VP.n19 VP.n18 24.3439
R2438 VP.n20 VP.n19 24.3439
R2439 VP.n13 VP.n12 24.3439
R2440 VP.n14 VP.n13 24.3439
R2441 VP.n14 VP.n9 24.3439
R2442 VP.n25 VP.n24 19.4752
R2443 VP.n43 VP.n0 19.4752
R2444 VP.n20 VP.n7 19.4752
R2445 VP.n11 VP.n10 3.94995
R2446 VP.n22 VP.n21 0.355081
R2447 VP.n26 VP.n23 0.355081
R2448 VP.n45 VP.n44 0.355081
R2449 VP VP.n45 0.26685
R2450 VP.n15 VP.n10 0.189894
R2451 VP.n16 VP.n15 0.189894
R2452 VP.n17 VP.n16 0.189894
R2453 VP.n17 VP.n8 0.189894
R2454 VP.n21 VP.n8 0.189894
R2455 VP.n27 VP.n26 0.189894
R2456 VP.n28 VP.n27 0.189894
R2457 VP.n28 VP.n5 0.189894
R2458 VP.n32 VP.n5 0.189894
R2459 VP.n33 VP.n32 0.189894
R2460 VP.n34 VP.n33 0.189894
R2461 VP.n34 VP.n3 0.189894
R2462 VP.n38 VP.n3 0.189894
R2463 VP.n39 VP.n38 0.189894
R2464 VP.n40 VP.n39 0.189894
R2465 VP.n40 VP.n1 0.189894
R2466 VP.n44 VP.n1 0.189894
R2467 VDD1.n64 VDD1.n0 289.615
R2468 VDD1.n133 VDD1.n69 289.615
R2469 VDD1.n65 VDD1.n64 185
R2470 VDD1.n63 VDD1.n62 185
R2471 VDD1.n4 VDD1.n3 185
R2472 VDD1.n57 VDD1.n56 185
R2473 VDD1.n55 VDD1.n54 185
R2474 VDD1.n8 VDD1.n7 185
R2475 VDD1.n49 VDD1.n48 185
R2476 VDD1.n47 VDD1.n46 185
R2477 VDD1.n45 VDD1.n11 185
R2478 VDD1.n15 VDD1.n12 185
R2479 VDD1.n40 VDD1.n39 185
R2480 VDD1.n38 VDD1.n37 185
R2481 VDD1.n17 VDD1.n16 185
R2482 VDD1.n32 VDD1.n31 185
R2483 VDD1.n30 VDD1.n29 185
R2484 VDD1.n21 VDD1.n20 185
R2485 VDD1.n24 VDD1.n23 185
R2486 VDD1.n92 VDD1.n91 185
R2487 VDD1.n89 VDD1.n88 185
R2488 VDD1.n98 VDD1.n97 185
R2489 VDD1.n100 VDD1.n99 185
R2490 VDD1.n85 VDD1.n84 185
R2491 VDD1.n106 VDD1.n105 185
R2492 VDD1.n109 VDD1.n108 185
R2493 VDD1.n107 VDD1.n81 185
R2494 VDD1.n114 VDD1.n80 185
R2495 VDD1.n116 VDD1.n115 185
R2496 VDD1.n118 VDD1.n117 185
R2497 VDD1.n77 VDD1.n76 185
R2498 VDD1.n124 VDD1.n123 185
R2499 VDD1.n126 VDD1.n125 185
R2500 VDD1.n73 VDD1.n72 185
R2501 VDD1.n132 VDD1.n131 185
R2502 VDD1.n134 VDD1.n133 185
R2503 VDD1.t4 VDD1.n22 149.524
R2504 VDD1.t2 VDD1.n90 149.524
R2505 VDD1.n64 VDD1.n63 104.615
R2506 VDD1.n63 VDD1.n3 104.615
R2507 VDD1.n56 VDD1.n3 104.615
R2508 VDD1.n56 VDD1.n55 104.615
R2509 VDD1.n55 VDD1.n7 104.615
R2510 VDD1.n48 VDD1.n7 104.615
R2511 VDD1.n48 VDD1.n47 104.615
R2512 VDD1.n47 VDD1.n11 104.615
R2513 VDD1.n15 VDD1.n11 104.615
R2514 VDD1.n39 VDD1.n15 104.615
R2515 VDD1.n39 VDD1.n38 104.615
R2516 VDD1.n38 VDD1.n16 104.615
R2517 VDD1.n31 VDD1.n16 104.615
R2518 VDD1.n31 VDD1.n30 104.615
R2519 VDD1.n30 VDD1.n20 104.615
R2520 VDD1.n23 VDD1.n20 104.615
R2521 VDD1.n91 VDD1.n88 104.615
R2522 VDD1.n98 VDD1.n88 104.615
R2523 VDD1.n99 VDD1.n98 104.615
R2524 VDD1.n99 VDD1.n84 104.615
R2525 VDD1.n106 VDD1.n84 104.615
R2526 VDD1.n108 VDD1.n106 104.615
R2527 VDD1.n108 VDD1.n107 104.615
R2528 VDD1.n107 VDD1.n80 104.615
R2529 VDD1.n116 VDD1.n80 104.615
R2530 VDD1.n117 VDD1.n116 104.615
R2531 VDD1.n117 VDD1.n76 104.615
R2532 VDD1.n124 VDD1.n76 104.615
R2533 VDD1.n125 VDD1.n124 104.615
R2534 VDD1.n125 VDD1.n72 104.615
R2535 VDD1.n132 VDD1.n72 104.615
R2536 VDD1.n133 VDD1.n132 104.615
R2537 VDD1.n139 VDD1.n138 60.4413
R2538 VDD1.n141 VDD1.n140 59.7637
R2539 VDD1.n23 VDD1.t4 52.3082
R2540 VDD1.n91 VDD1.t2 52.3082
R2541 VDD1 VDD1.n68 49.1812
R2542 VDD1.n139 VDD1.n137 49.0677
R2543 VDD1.n141 VDD1.n139 46.2724
R2544 VDD1.n46 VDD1.n45 13.1884
R2545 VDD1.n115 VDD1.n114 13.1884
R2546 VDD1.n49 VDD1.n10 12.8005
R2547 VDD1.n44 VDD1.n12 12.8005
R2548 VDD1.n113 VDD1.n81 12.8005
R2549 VDD1.n118 VDD1.n79 12.8005
R2550 VDD1.n50 VDD1.n8 12.0247
R2551 VDD1.n41 VDD1.n40 12.0247
R2552 VDD1.n110 VDD1.n109 12.0247
R2553 VDD1.n119 VDD1.n77 12.0247
R2554 VDD1.n54 VDD1.n53 11.249
R2555 VDD1.n37 VDD1.n14 11.249
R2556 VDD1.n105 VDD1.n83 11.249
R2557 VDD1.n123 VDD1.n122 11.249
R2558 VDD1.n57 VDD1.n6 10.4732
R2559 VDD1.n36 VDD1.n17 10.4732
R2560 VDD1.n104 VDD1.n85 10.4732
R2561 VDD1.n126 VDD1.n75 10.4732
R2562 VDD1.n24 VDD1.n22 10.2747
R2563 VDD1.n92 VDD1.n90 10.2747
R2564 VDD1.n58 VDD1.n4 9.69747
R2565 VDD1.n33 VDD1.n32 9.69747
R2566 VDD1.n101 VDD1.n100 9.69747
R2567 VDD1.n127 VDD1.n73 9.69747
R2568 VDD1.n68 VDD1.n67 9.45567
R2569 VDD1.n137 VDD1.n136 9.45567
R2570 VDD1.n26 VDD1.n25 9.3005
R2571 VDD1.n28 VDD1.n27 9.3005
R2572 VDD1.n19 VDD1.n18 9.3005
R2573 VDD1.n34 VDD1.n33 9.3005
R2574 VDD1.n36 VDD1.n35 9.3005
R2575 VDD1.n14 VDD1.n13 9.3005
R2576 VDD1.n42 VDD1.n41 9.3005
R2577 VDD1.n44 VDD1.n43 9.3005
R2578 VDD1.n67 VDD1.n66 9.3005
R2579 VDD1.n2 VDD1.n1 9.3005
R2580 VDD1.n61 VDD1.n60 9.3005
R2581 VDD1.n59 VDD1.n58 9.3005
R2582 VDD1.n6 VDD1.n5 9.3005
R2583 VDD1.n53 VDD1.n52 9.3005
R2584 VDD1.n51 VDD1.n50 9.3005
R2585 VDD1.n10 VDD1.n9 9.3005
R2586 VDD1.n71 VDD1.n70 9.3005
R2587 VDD1.n130 VDD1.n129 9.3005
R2588 VDD1.n128 VDD1.n127 9.3005
R2589 VDD1.n75 VDD1.n74 9.3005
R2590 VDD1.n122 VDD1.n121 9.3005
R2591 VDD1.n120 VDD1.n119 9.3005
R2592 VDD1.n79 VDD1.n78 9.3005
R2593 VDD1.n94 VDD1.n93 9.3005
R2594 VDD1.n96 VDD1.n95 9.3005
R2595 VDD1.n87 VDD1.n86 9.3005
R2596 VDD1.n102 VDD1.n101 9.3005
R2597 VDD1.n104 VDD1.n103 9.3005
R2598 VDD1.n83 VDD1.n82 9.3005
R2599 VDD1.n111 VDD1.n110 9.3005
R2600 VDD1.n113 VDD1.n112 9.3005
R2601 VDD1.n136 VDD1.n135 9.3005
R2602 VDD1.n62 VDD1.n61 8.92171
R2603 VDD1.n29 VDD1.n19 8.92171
R2604 VDD1.n97 VDD1.n87 8.92171
R2605 VDD1.n131 VDD1.n130 8.92171
R2606 VDD1.n65 VDD1.n2 8.14595
R2607 VDD1.n28 VDD1.n21 8.14595
R2608 VDD1.n96 VDD1.n89 8.14595
R2609 VDD1.n134 VDD1.n71 8.14595
R2610 VDD1.n66 VDD1.n0 7.3702
R2611 VDD1.n25 VDD1.n24 7.3702
R2612 VDD1.n93 VDD1.n92 7.3702
R2613 VDD1.n135 VDD1.n69 7.3702
R2614 VDD1.n68 VDD1.n0 6.59444
R2615 VDD1.n137 VDD1.n69 6.59444
R2616 VDD1.n66 VDD1.n65 5.81868
R2617 VDD1.n25 VDD1.n21 5.81868
R2618 VDD1.n93 VDD1.n89 5.81868
R2619 VDD1.n135 VDD1.n134 5.81868
R2620 VDD1.n62 VDD1.n2 5.04292
R2621 VDD1.n29 VDD1.n28 5.04292
R2622 VDD1.n97 VDD1.n96 5.04292
R2623 VDD1.n131 VDD1.n71 5.04292
R2624 VDD1.n61 VDD1.n4 4.26717
R2625 VDD1.n32 VDD1.n19 4.26717
R2626 VDD1.n100 VDD1.n87 4.26717
R2627 VDD1.n130 VDD1.n73 4.26717
R2628 VDD1.n58 VDD1.n57 3.49141
R2629 VDD1.n33 VDD1.n17 3.49141
R2630 VDD1.n101 VDD1.n85 3.49141
R2631 VDD1.n127 VDD1.n126 3.49141
R2632 VDD1.n26 VDD1.n22 2.84303
R2633 VDD1.n94 VDD1.n90 2.84303
R2634 VDD1.n54 VDD1.n6 2.71565
R2635 VDD1.n37 VDD1.n36 2.71565
R2636 VDD1.n105 VDD1.n104 2.71565
R2637 VDD1.n123 VDD1.n75 2.71565
R2638 VDD1.n53 VDD1.n8 1.93989
R2639 VDD1.n40 VDD1.n14 1.93989
R2640 VDD1.n109 VDD1.n83 1.93989
R2641 VDD1.n122 VDD1.n77 1.93989
R2642 VDD1.n140 VDD1.t3 1.55466
R2643 VDD1.n140 VDD1.t1 1.55466
R2644 VDD1.n138 VDD1.t0 1.55466
R2645 VDD1.n138 VDD1.t5 1.55466
R2646 VDD1.n50 VDD1.n49 1.16414
R2647 VDD1.n41 VDD1.n12 1.16414
R2648 VDD1.n110 VDD1.n81 1.16414
R2649 VDD1.n119 VDD1.n118 1.16414
R2650 VDD1 VDD1.n141 0.675069
R2651 VDD1.n46 VDD1.n10 0.388379
R2652 VDD1.n45 VDD1.n44 0.388379
R2653 VDD1.n114 VDD1.n113 0.388379
R2654 VDD1.n115 VDD1.n79 0.388379
R2655 VDD1.n67 VDD1.n1 0.155672
R2656 VDD1.n60 VDD1.n1 0.155672
R2657 VDD1.n60 VDD1.n59 0.155672
R2658 VDD1.n59 VDD1.n5 0.155672
R2659 VDD1.n52 VDD1.n5 0.155672
R2660 VDD1.n52 VDD1.n51 0.155672
R2661 VDD1.n51 VDD1.n9 0.155672
R2662 VDD1.n43 VDD1.n9 0.155672
R2663 VDD1.n43 VDD1.n42 0.155672
R2664 VDD1.n42 VDD1.n13 0.155672
R2665 VDD1.n35 VDD1.n13 0.155672
R2666 VDD1.n35 VDD1.n34 0.155672
R2667 VDD1.n34 VDD1.n18 0.155672
R2668 VDD1.n27 VDD1.n18 0.155672
R2669 VDD1.n27 VDD1.n26 0.155672
R2670 VDD1.n95 VDD1.n94 0.155672
R2671 VDD1.n95 VDD1.n86 0.155672
R2672 VDD1.n102 VDD1.n86 0.155672
R2673 VDD1.n103 VDD1.n102 0.155672
R2674 VDD1.n103 VDD1.n82 0.155672
R2675 VDD1.n111 VDD1.n82 0.155672
R2676 VDD1.n112 VDD1.n111 0.155672
R2677 VDD1.n112 VDD1.n78 0.155672
R2678 VDD1.n120 VDD1.n78 0.155672
R2679 VDD1.n121 VDD1.n120 0.155672
R2680 VDD1.n121 VDD1.n74 0.155672
R2681 VDD1.n128 VDD1.n74 0.155672
R2682 VDD1.n129 VDD1.n128 0.155672
R2683 VDD1.n129 VDD1.n70 0.155672
R2684 VDD1.n136 VDD1.n70 0.155672
C0 VDD1 VDD2 1.59096f
C1 VTAIL VDD1 8.10421f
C2 VP VN 7.527441f
C3 VP VDD2 0.497975f
C4 VP VTAIL 7.57766f
C5 VN VDD2 7.32442f
C6 VN VTAIL 7.5634f
C7 VP VDD1 7.668049f
C8 VTAIL VDD2 8.158501f
C9 VN VDD1 0.151137f
C10 VDD2 B 6.481663f
C11 VDD1 B 6.626123f
C12 VTAIL B 8.428585f
C13 VN B 14.331632f
C14 VP B 12.998486f
C15 VDD1.n0 B 0.029548f
C16 VDD1.n1 B 0.021645f
C17 VDD1.n2 B 0.011631f
C18 VDD1.n3 B 0.027492f
C19 VDD1.n4 B 0.012315f
C20 VDD1.n5 B 0.021645f
C21 VDD1.n6 B 0.011631f
C22 VDD1.n7 B 0.027492f
C23 VDD1.n8 B 0.012315f
C24 VDD1.n9 B 0.021645f
C25 VDD1.n10 B 0.011631f
C26 VDD1.n11 B 0.027492f
C27 VDD1.n12 B 0.012315f
C28 VDD1.n13 B 0.021645f
C29 VDD1.n14 B 0.011631f
C30 VDD1.n15 B 0.027492f
C31 VDD1.n16 B 0.027492f
C32 VDD1.n17 B 0.012315f
C33 VDD1.n18 B 0.021645f
C34 VDD1.n19 B 0.011631f
C35 VDD1.n20 B 0.027492f
C36 VDD1.n21 B 0.012315f
C37 VDD1.n22 B 0.162211f
C38 VDD1.t4 B 0.046519f
C39 VDD1.n23 B 0.020619f
C40 VDD1.n24 B 0.019435f
C41 VDD1.n25 B 0.011631f
C42 VDD1.n26 B 1.16322f
C43 VDD1.n27 B 0.021645f
C44 VDD1.n28 B 0.011631f
C45 VDD1.n29 B 0.012315f
C46 VDD1.n30 B 0.027492f
C47 VDD1.n31 B 0.027492f
C48 VDD1.n32 B 0.012315f
C49 VDD1.n33 B 0.011631f
C50 VDD1.n34 B 0.021645f
C51 VDD1.n35 B 0.021645f
C52 VDD1.n36 B 0.011631f
C53 VDD1.n37 B 0.012315f
C54 VDD1.n38 B 0.027492f
C55 VDD1.n39 B 0.027492f
C56 VDD1.n40 B 0.012315f
C57 VDD1.n41 B 0.011631f
C58 VDD1.n42 B 0.021645f
C59 VDD1.n43 B 0.021645f
C60 VDD1.n44 B 0.011631f
C61 VDD1.n45 B 0.011973f
C62 VDD1.n46 B 0.011973f
C63 VDD1.n47 B 0.027492f
C64 VDD1.n48 B 0.027492f
C65 VDD1.n49 B 0.012315f
C66 VDD1.n50 B 0.011631f
C67 VDD1.n51 B 0.021645f
C68 VDD1.n52 B 0.021645f
C69 VDD1.n53 B 0.011631f
C70 VDD1.n54 B 0.012315f
C71 VDD1.n55 B 0.027492f
C72 VDD1.n56 B 0.027492f
C73 VDD1.n57 B 0.012315f
C74 VDD1.n58 B 0.011631f
C75 VDD1.n59 B 0.021645f
C76 VDD1.n60 B 0.021645f
C77 VDD1.n61 B 0.011631f
C78 VDD1.n62 B 0.012315f
C79 VDD1.n63 B 0.027492f
C80 VDD1.n64 B 0.057967f
C81 VDD1.n65 B 0.012315f
C82 VDD1.n66 B 0.011631f
C83 VDD1.n67 B 0.047075f
C84 VDD1.n68 B 0.056208f
C85 VDD1.n69 B 0.029548f
C86 VDD1.n70 B 0.021645f
C87 VDD1.n71 B 0.011631f
C88 VDD1.n72 B 0.027492f
C89 VDD1.n73 B 0.012315f
C90 VDD1.n74 B 0.021645f
C91 VDD1.n75 B 0.011631f
C92 VDD1.n76 B 0.027492f
C93 VDD1.n77 B 0.012315f
C94 VDD1.n78 B 0.021645f
C95 VDD1.n79 B 0.011631f
C96 VDD1.n80 B 0.027492f
C97 VDD1.n81 B 0.012315f
C98 VDD1.n82 B 0.021645f
C99 VDD1.n83 B 0.011631f
C100 VDD1.n84 B 0.027492f
C101 VDD1.n85 B 0.012315f
C102 VDD1.n86 B 0.021645f
C103 VDD1.n87 B 0.011631f
C104 VDD1.n88 B 0.027492f
C105 VDD1.n89 B 0.012315f
C106 VDD1.n90 B 0.162211f
C107 VDD1.t2 B 0.046519f
C108 VDD1.n91 B 0.020619f
C109 VDD1.n92 B 0.019435f
C110 VDD1.n93 B 0.011631f
C111 VDD1.n94 B 1.16322f
C112 VDD1.n95 B 0.021645f
C113 VDD1.n96 B 0.011631f
C114 VDD1.n97 B 0.012315f
C115 VDD1.n98 B 0.027492f
C116 VDD1.n99 B 0.027492f
C117 VDD1.n100 B 0.012315f
C118 VDD1.n101 B 0.011631f
C119 VDD1.n102 B 0.021645f
C120 VDD1.n103 B 0.021645f
C121 VDD1.n104 B 0.011631f
C122 VDD1.n105 B 0.012315f
C123 VDD1.n106 B 0.027492f
C124 VDD1.n107 B 0.027492f
C125 VDD1.n108 B 0.027492f
C126 VDD1.n109 B 0.012315f
C127 VDD1.n110 B 0.011631f
C128 VDD1.n111 B 0.021645f
C129 VDD1.n112 B 0.021645f
C130 VDD1.n113 B 0.011631f
C131 VDD1.n114 B 0.011973f
C132 VDD1.n115 B 0.011973f
C133 VDD1.n116 B 0.027492f
C134 VDD1.n117 B 0.027492f
C135 VDD1.n118 B 0.012315f
C136 VDD1.n119 B 0.011631f
C137 VDD1.n120 B 0.021645f
C138 VDD1.n121 B 0.021645f
C139 VDD1.n122 B 0.011631f
C140 VDD1.n123 B 0.012315f
C141 VDD1.n124 B 0.027492f
C142 VDD1.n125 B 0.027492f
C143 VDD1.n126 B 0.012315f
C144 VDD1.n127 B 0.011631f
C145 VDD1.n128 B 0.021645f
C146 VDD1.n129 B 0.021645f
C147 VDD1.n130 B 0.011631f
C148 VDD1.n131 B 0.012315f
C149 VDD1.n132 B 0.027492f
C150 VDD1.n133 B 0.057967f
C151 VDD1.n134 B 0.012315f
C152 VDD1.n135 B 0.011631f
C153 VDD1.n136 B 0.047075f
C154 VDD1.n137 B 0.055437f
C155 VDD1.t0 B 0.217917f
C156 VDD1.t5 B 0.217917f
C157 VDD1.n138 B 1.95136f
C158 VDD1.n139 B 2.65452f
C159 VDD1.t3 B 0.217917f
C160 VDD1.t1 B 0.217917f
C161 VDD1.n140 B 1.94639f
C162 VDD1.n141 B 2.58272f
C163 VP.t0 B 2.25599f
C164 VP.n0 B 0.876875f
C165 VP.n1 B 0.021135f
C166 VP.n2 B 0.028022f
C167 VP.n3 B 0.021135f
C168 VP.t5 B 2.25599f
C169 VP.n4 B 0.039588f
C170 VP.n5 B 0.021135f
C171 VP.n6 B 0.039588f
C172 VP.t4 B 2.25599f
C173 VP.n7 B 0.876875f
C174 VP.n8 B 0.021135f
C175 VP.n9 B 0.028022f
C176 VP.n10 B 0.240641f
C177 VP.t2 B 2.25599f
C178 VP.t1 B 2.49127f
C179 VP.n11 B 0.827548f
C180 VP.n12 B 0.871372f
C181 VP.n13 B 0.039588f
C182 VP.n14 B 0.039588f
C183 VP.n15 B 0.021135f
C184 VP.n16 B 0.021135f
C185 VP.n17 B 0.021135f
C186 VP.n18 B 0.033953f
C187 VP.n19 B 0.039588f
C188 VP.n20 B 0.035679f
C189 VP.n21 B 0.034117f
C190 VP.n22 B 1.23785f
C191 VP.n23 B 1.25264f
C192 VP.t3 B 2.25599f
C193 VP.n24 B 0.876875f
C194 VP.n25 B 0.035679f
C195 VP.n26 B 0.034117f
C196 VP.n27 B 0.021135f
C197 VP.n28 B 0.021135f
C198 VP.n29 B 0.033953f
C199 VP.n30 B 0.028022f
C200 VP.n31 B 0.039588f
C201 VP.n32 B 0.021135f
C202 VP.n33 B 0.021135f
C203 VP.n34 B 0.021135f
C204 VP.n35 B 0.811787f
C205 VP.n36 B 0.039588f
C206 VP.n37 B 0.039588f
C207 VP.n38 B 0.021135f
C208 VP.n39 B 0.021135f
C209 VP.n40 B 0.021135f
C210 VP.n41 B 0.033953f
C211 VP.n42 B 0.039588f
C212 VP.n43 B 0.035679f
C213 VP.n44 B 0.034117f
C214 VP.n45 B 0.04492f
C215 VTAIL.t8 B 0.240383f
C216 VTAIL.t9 B 0.240383f
C217 VTAIL.n0 B 2.07101f
C218 VTAIL.n1 B 0.454319f
C219 VTAIL.n2 B 0.032595f
C220 VTAIL.n3 B 0.023877f
C221 VTAIL.n4 B 0.01283f
C222 VTAIL.n5 B 0.030326f
C223 VTAIL.n6 B 0.013585f
C224 VTAIL.n7 B 0.023877f
C225 VTAIL.n8 B 0.01283f
C226 VTAIL.n9 B 0.030326f
C227 VTAIL.n10 B 0.013585f
C228 VTAIL.n11 B 0.023877f
C229 VTAIL.n12 B 0.01283f
C230 VTAIL.n13 B 0.030326f
C231 VTAIL.n14 B 0.013585f
C232 VTAIL.n15 B 0.023877f
C233 VTAIL.n16 B 0.01283f
C234 VTAIL.n17 B 0.030326f
C235 VTAIL.n18 B 0.013585f
C236 VTAIL.n19 B 0.023877f
C237 VTAIL.n20 B 0.01283f
C238 VTAIL.n21 B 0.030326f
C239 VTAIL.n22 B 0.013585f
C240 VTAIL.n23 B 0.178934f
C241 VTAIL.t3 B 0.051315f
C242 VTAIL.n24 B 0.022745f
C243 VTAIL.n25 B 0.021438f
C244 VTAIL.n26 B 0.01283f
C245 VTAIL.n27 B 1.28314f
C246 VTAIL.n28 B 0.023877f
C247 VTAIL.n29 B 0.01283f
C248 VTAIL.n30 B 0.013585f
C249 VTAIL.n31 B 0.030326f
C250 VTAIL.n32 B 0.030326f
C251 VTAIL.n33 B 0.013585f
C252 VTAIL.n34 B 0.01283f
C253 VTAIL.n35 B 0.023877f
C254 VTAIL.n36 B 0.023877f
C255 VTAIL.n37 B 0.01283f
C256 VTAIL.n38 B 0.013585f
C257 VTAIL.n39 B 0.030326f
C258 VTAIL.n40 B 0.030326f
C259 VTAIL.n41 B 0.030326f
C260 VTAIL.n42 B 0.013585f
C261 VTAIL.n43 B 0.01283f
C262 VTAIL.n44 B 0.023877f
C263 VTAIL.n45 B 0.023877f
C264 VTAIL.n46 B 0.01283f
C265 VTAIL.n47 B 0.013208f
C266 VTAIL.n48 B 0.013208f
C267 VTAIL.n49 B 0.030326f
C268 VTAIL.n50 B 0.030326f
C269 VTAIL.n51 B 0.013585f
C270 VTAIL.n52 B 0.01283f
C271 VTAIL.n53 B 0.023877f
C272 VTAIL.n54 B 0.023877f
C273 VTAIL.n55 B 0.01283f
C274 VTAIL.n56 B 0.013585f
C275 VTAIL.n57 B 0.030326f
C276 VTAIL.n58 B 0.030326f
C277 VTAIL.n59 B 0.013585f
C278 VTAIL.n60 B 0.01283f
C279 VTAIL.n61 B 0.023877f
C280 VTAIL.n62 B 0.023877f
C281 VTAIL.n63 B 0.01283f
C282 VTAIL.n64 B 0.013585f
C283 VTAIL.n65 B 0.030326f
C284 VTAIL.n66 B 0.063943f
C285 VTAIL.n67 B 0.013585f
C286 VTAIL.n68 B 0.01283f
C287 VTAIL.n69 B 0.051929f
C288 VTAIL.n70 B 0.0355f
C289 VTAIL.n71 B 0.392959f
C290 VTAIL.t1 B 0.240383f
C291 VTAIL.t0 B 0.240383f
C292 VTAIL.n72 B 2.07101f
C293 VTAIL.n73 B 2.0904f
C294 VTAIL.t7 B 0.240383f
C295 VTAIL.t10 B 0.240383f
C296 VTAIL.n74 B 2.07102f
C297 VTAIL.n75 B 2.0904f
C298 VTAIL.n76 B 0.032595f
C299 VTAIL.n77 B 0.023877f
C300 VTAIL.n78 B 0.01283f
C301 VTAIL.n79 B 0.030326f
C302 VTAIL.n80 B 0.013585f
C303 VTAIL.n81 B 0.023877f
C304 VTAIL.n82 B 0.01283f
C305 VTAIL.n83 B 0.030326f
C306 VTAIL.n84 B 0.013585f
C307 VTAIL.n85 B 0.023877f
C308 VTAIL.n86 B 0.01283f
C309 VTAIL.n87 B 0.030326f
C310 VTAIL.n88 B 0.013585f
C311 VTAIL.n89 B 0.023877f
C312 VTAIL.n90 B 0.01283f
C313 VTAIL.n91 B 0.030326f
C314 VTAIL.n92 B 0.030326f
C315 VTAIL.n93 B 0.013585f
C316 VTAIL.n94 B 0.023877f
C317 VTAIL.n95 B 0.01283f
C318 VTAIL.n96 B 0.030326f
C319 VTAIL.n97 B 0.013585f
C320 VTAIL.n98 B 0.178934f
C321 VTAIL.t6 B 0.051315f
C322 VTAIL.n99 B 0.022745f
C323 VTAIL.n100 B 0.021438f
C324 VTAIL.n101 B 0.01283f
C325 VTAIL.n102 B 1.28314f
C326 VTAIL.n103 B 0.023877f
C327 VTAIL.n104 B 0.01283f
C328 VTAIL.n105 B 0.013585f
C329 VTAIL.n106 B 0.030326f
C330 VTAIL.n107 B 0.030326f
C331 VTAIL.n108 B 0.013585f
C332 VTAIL.n109 B 0.01283f
C333 VTAIL.n110 B 0.023877f
C334 VTAIL.n111 B 0.023877f
C335 VTAIL.n112 B 0.01283f
C336 VTAIL.n113 B 0.013585f
C337 VTAIL.n114 B 0.030326f
C338 VTAIL.n115 B 0.030326f
C339 VTAIL.n116 B 0.013585f
C340 VTAIL.n117 B 0.01283f
C341 VTAIL.n118 B 0.023877f
C342 VTAIL.n119 B 0.023877f
C343 VTAIL.n120 B 0.01283f
C344 VTAIL.n121 B 0.013208f
C345 VTAIL.n122 B 0.013208f
C346 VTAIL.n123 B 0.030326f
C347 VTAIL.n124 B 0.030326f
C348 VTAIL.n125 B 0.013585f
C349 VTAIL.n126 B 0.01283f
C350 VTAIL.n127 B 0.023877f
C351 VTAIL.n128 B 0.023877f
C352 VTAIL.n129 B 0.01283f
C353 VTAIL.n130 B 0.013585f
C354 VTAIL.n131 B 0.030326f
C355 VTAIL.n132 B 0.030326f
C356 VTAIL.n133 B 0.013585f
C357 VTAIL.n134 B 0.01283f
C358 VTAIL.n135 B 0.023877f
C359 VTAIL.n136 B 0.023877f
C360 VTAIL.n137 B 0.01283f
C361 VTAIL.n138 B 0.013585f
C362 VTAIL.n139 B 0.030326f
C363 VTAIL.n140 B 0.063943f
C364 VTAIL.n141 B 0.013585f
C365 VTAIL.n142 B 0.01283f
C366 VTAIL.n143 B 0.051929f
C367 VTAIL.n144 B 0.0355f
C368 VTAIL.n145 B 0.392959f
C369 VTAIL.t2 B 0.240383f
C370 VTAIL.t11 B 0.240383f
C371 VTAIL.n146 B 2.07102f
C372 VTAIL.n147 B 0.618968f
C373 VTAIL.n148 B 0.032595f
C374 VTAIL.n149 B 0.023877f
C375 VTAIL.n150 B 0.01283f
C376 VTAIL.n151 B 0.030326f
C377 VTAIL.n152 B 0.013585f
C378 VTAIL.n153 B 0.023877f
C379 VTAIL.n154 B 0.01283f
C380 VTAIL.n155 B 0.030326f
C381 VTAIL.n156 B 0.013585f
C382 VTAIL.n157 B 0.023877f
C383 VTAIL.n158 B 0.01283f
C384 VTAIL.n159 B 0.030326f
C385 VTAIL.n160 B 0.013585f
C386 VTAIL.n161 B 0.023877f
C387 VTAIL.n162 B 0.01283f
C388 VTAIL.n163 B 0.030326f
C389 VTAIL.n164 B 0.030326f
C390 VTAIL.n165 B 0.013585f
C391 VTAIL.n166 B 0.023877f
C392 VTAIL.n167 B 0.01283f
C393 VTAIL.n168 B 0.030326f
C394 VTAIL.n169 B 0.013585f
C395 VTAIL.n170 B 0.178934f
C396 VTAIL.t4 B 0.051315f
C397 VTAIL.n171 B 0.022745f
C398 VTAIL.n172 B 0.021438f
C399 VTAIL.n173 B 0.01283f
C400 VTAIL.n174 B 1.28314f
C401 VTAIL.n175 B 0.023877f
C402 VTAIL.n176 B 0.01283f
C403 VTAIL.n177 B 0.013585f
C404 VTAIL.n178 B 0.030326f
C405 VTAIL.n179 B 0.030326f
C406 VTAIL.n180 B 0.013585f
C407 VTAIL.n181 B 0.01283f
C408 VTAIL.n182 B 0.023877f
C409 VTAIL.n183 B 0.023877f
C410 VTAIL.n184 B 0.01283f
C411 VTAIL.n185 B 0.013585f
C412 VTAIL.n186 B 0.030326f
C413 VTAIL.n187 B 0.030326f
C414 VTAIL.n188 B 0.013585f
C415 VTAIL.n189 B 0.01283f
C416 VTAIL.n190 B 0.023877f
C417 VTAIL.n191 B 0.023877f
C418 VTAIL.n192 B 0.01283f
C419 VTAIL.n193 B 0.013208f
C420 VTAIL.n194 B 0.013208f
C421 VTAIL.n195 B 0.030326f
C422 VTAIL.n196 B 0.030326f
C423 VTAIL.n197 B 0.013585f
C424 VTAIL.n198 B 0.01283f
C425 VTAIL.n199 B 0.023877f
C426 VTAIL.n200 B 0.023877f
C427 VTAIL.n201 B 0.01283f
C428 VTAIL.n202 B 0.013585f
C429 VTAIL.n203 B 0.030326f
C430 VTAIL.n204 B 0.030326f
C431 VTAIL.n205 B 0.013585f
C432 VTAIL.n206 B 0.01283f
C433 VTAIL.n207 B 0.023877f
C434 VTAIL.n208 B 0.023877f
C435 VTAIL.n209 B 0.01283f
C436 VTAIL.n210 B 0.013585f
C437 VTAIL.n211 B 0.030326f
C438 VTAIL.n212 B 0.063943f
C439 VTAIL.n213 B 0.013585f
C440 VTAIL.n214 B 0.01283f
C441 VTAIL.n215 B 0.051929f
C442 VTAIL.n216 B 0.0355f
C443 VTAIL.n217 B 1.63889f
C444 VTAIL.n218 B 0.032595f
C445 VTAIL.n219 B 0.023877f
C446 VTAIL.n220 B 0.01283f
C447 VTAIL.n221 B 0.030326f
C448 VTAIL.n222 B 0.013585f
C449 VTAIL.n223 B 0.023877f
C450 VTAIL.n224 B 0.01283f
C451 VTAIL.n225 B 0.030326f
C452 VTAIL.n226 B 0.013585f
C453 VTAIL.n227 B 0.023877f
C454 VTAIL.n228 B 0.01283f
C455 VTAIL.n229 B 0.030326f
C456 VTAIL.n230 B 0.013585f
C457 VTAIL.n231 B 0.023877f
C458 VTAIL.n232 B 0.01283f
C459 VTAIL.n233 B 0.030326f
C460 VTAIL.n234 B 0.013585f
C461 VTAIL.n235 B 0.023877f
C462 VTAIL.n236 B 0.01283f
C463 VTAIL.n237 B 0.030326f
C464 VTAIL.n238 B 0.013585f
C465 VTAIL.n239 B 0.178934f
C466 VTAIL.t5 B 0.051315f
C467 VTAIL.n240 B 0.022745f
C468 VTAIL.n241 B 0.021438f
C469 VTAIL.n242 B 0.01283f
C470 VTAIL.n243 B 1.28314f
C471 VTAIL.n244 B 0.023877f
C472 VTAIL.n245 B 0.01283f
C473 VTAIL.n246 B 0.013585f
C474 VTAIL.n247 B 0.030326f
C475 VTAIL.n248 B 0.030326f
C476 VTAIL.n249 B 0.013585f
C477 VTAIL.n250 B 0.01283f
C478 VTAIL.n251 B 0.023877f
C479 VTAIL.n252 B 0.023877f
C480 VTAIL.n253 B 0.01283f
C481 VTAIL.n254 B 0.013585f
C482 VTAIL.n255 B 0.030326f
C483 VTAIL.n256 B 0.030326f
C484 VTAIL.n257 B 0.030326f
C485 VTAIL.n258 B 0.013585f
C486 VTAIL.n259 B 0.01283f
C487 VTAIL.n260 B 0.023877f
C488 VTAIL.n261 B 0.023877f
C489 VTAIL.n262 B 0.01283f
C490 VTAIL.n263 B 0.013208f
C491 VTAIL.n264 B 0.013208f
C492 VTAIL.n265 B 0.030326f
C493 VTAIL.n266 B 0.030326f
C494 VTAIL.n267 B 0.013585f
C495 VTAIL.n268 B 0.01283f
C496 VTAIL.n269 B 0.023877f
C497 VTAIL.n270 B 0.023877f
C498 VTAIL.n271 B 0.01283f
C499 VTAIL.n272 B 0.013585f
C500 VTAIL.n273 B 0.030326f
C501 VTAIL.n274 B 0.030326f
C502 VTAIL.n275 B 0.013585f
C503 VTAIL.n276 B 0.01283f
C504 VTAIL.n277 B 0.023877f
C505 VTAIL.n278 B 0.023877f
C506 VTAIL.n279 B 0.01283f
C507 VTAIL.n280 B 0.013585f
C508 VTAIL.n281 B 0.030326f
C509 VTAIL.n282 B 0.063943f
C510 VTAIL.n283 B 0.013585f
C511 VTAIL.n284 B 0.01283f
C512 VTAIL.n285 B 0.051929f
C513 VTAIL.n286 B 0.0355f
C514 VTAIL.n287 B 1.57803f
C515 VDD2.n0 B 0.029135f
C516 VDD2.n1 B 0.021343f
C517 VDD2.n2 B 0.011468f
C518 VDD2.n3 B 0.027107f
C519 VDD2.n4 B 0.012143f
C520 VDD2.n5 B 0.021343f
C521 VDD2.n6 B 0.011468f
C522 VDD2.n7 B 0.027107f
C523 VDD2.n8 B 0.012143f
C524 VDD2.n9 B 0.021343f
C525 VDD2.n10 B 0.011468f
C526 VDD2.n11 B 0.027107f
C527 VDD2.n12 B 0.012143f
C528 VDD2.n13 B 0.021343f
C529 VDD2.n14 B 0.011468f
C530 VDD2.n15 B 0.027107f
C531 VDD2.n16 B 0.012143f
C532 VDD2.n17 B 0.021343f
C533 VDD2.n18 B 0.011468f
C534 VDD2.n19 B 0.027107f
C535 VDD2.n20 B 0.012143f
C536 VDD2.n21 B 0.15994f
C537 VDD2.t3 B 0.045868f
C538 VDD2.n22 B 0.020331f
C539 VDD2.n23 B 0.019163f
C540 VDD2.n24 B 0.011468f
C541 VDD2.n25 B 1.14694f
C542 VDD2.n26 B 0.021343f
C543 VDD2.n27 B 0.011468f
C544 VDD2.n28 B 0.012143f
C545 VDD2.n29 B 0.027107f
C546 VDD2.n30 B 0.027107f
C547 VDD2.n31 B 0.012143f
C548 VDD2.n32 B 0.011468f
C549 VDD2.n33 B 0.021343f
C550 VDD2.n34 B 0.021343f
C551 VDD2.n35 B 0.011468f
C552 VDD2.n36 B 0.012143f
C553 VDD2.n37 B 0.027107f
C554 VDD2.n38 B 0.027107f
C555 VDD2.n39 B 0.027107f
C556 VDD2.n40 B 0.012143f
C557 VDD2.n41 B 0.011468f
C558 VDD2.n42 B 0.021343f
C559 VDD2.n43 B 0.021343f
C560 VDD2.n44 B 0.011468f
C561 VDD2.n45 B 0.011806f
C562 VDD2.n46 B 0.011806f
C563 VDD2.n47 B 0.027107f
C564 VDD2.n48 B 0.027107f
C565 VDD2.n49 B 0.012143f
C566 VDD2.n50 B 0.011468f
C567 VDD2.n51 B 0.021343f
C568 VDD2.n52 B 0.021343f
C569 VDD2.n53 B 0.011468f
C570 VDD2.n54 B 0.012143f
C571 VDD2.n55 B 0.027107f
C572 VDD2.n56 B 0.027107f
C573 VDD2.n57 B 0.012143f
C574 VDD2.n58 B 0.011468f
C575 VDD2.n59 B 0.021343f
C576 VDD2.n60 B 0.021343f
C577 VDD2.n61 B 0.011468f
C578 VDD2.n62 B 0.012143f
C579 VDD2.n63 B 0.027107f
C580 VDD2.n64 B 0.057155f
C581 VDD2.n65 B 0.012143f
C582 VDD2.n66 B 0.011468f
C583 VDD2.n67 B 0.046416f
C584 VDD2.n68 B 0.054661f
C585 VDD2.t1 B 0.214866f
C586 VDD2.t2 B 0.214866f
C587 VDD2.n69 B 1.92405f
C588 VDD2.n70 B 2.5003f
C589 VDD2.n71 B 0.029135f
C590 VDD2.n72 B 0.021343f
C591 VDD2.n73 B 0.011468f
C592 VDD2.n74 B 0.027107f
C593 VDD2.n75 B 0.012143f
C594 VDD2.n76 B 0.021343f
C595 VDD2.n77 B 0.011468f
C596 VDD2.n78 B 0.027107f
C597 VDD2.n79 B 0.012143f
C598 VDD2.n80 B 0.021343f
C599 VDD2.n81 B 0.011468f
C600 VDD2.n82 B 0.027107f
C601 VDD2.n83 B 0.012143f
C602 VDD2.n84 B 0.021343f
C603 VDD2.n85 B 0.011468f
C604 VDD2.n86 B 0.027107f
C605 VDD2.n87 B 0.027107f
C606 VDD2.n88 B 0.012143f
C607 VDD2.n89 B 0.021343f
C608 VDD2.n90 B 0.011468f
C609 VDD2.n91 B 0.027107f
C610 VDD2.n92 B 0.012143f
C611 VDD2.n93 B 0.15994f
C612 VDD2.t5 B 0.045868f
C613 VDD2.n94 B 0.020331f
C614 VDD2.n95 B 0.019163f
C615 VDD2.n96 B 0.011468f
C616 VDD2.n97 B 1.14694f
C617 VDD2.n98 B 0.021343f
C618 VDD2.n99 B 0.011468f
C619 VDD2.n100 B 0.012143f
C620 VDD2.n101 B 0.027107f
C621 VDD2.n102 B 0.027107f
C622 VDD2.n103 B 0.012143f
C623 VDD2.n104 B 0.011468f
C624 VDD2.n105 B 0.021343f
C625 VDD2.n106 B 0.021343f
C626 VDD2.n107 B 0.011468f
C627 VDD2.n108 B 0.012143f
C628 VDD2.n109 B 0.027107f
C629 VDD2.n110 B 0.027107f
C630 VDD2.n111 B 0.012143f
C631 VDD2.n112 B 0.011468f
C632 VDD2.n113 B 0.021343f
C633 VDD2.n114 B 0.021343f
C634 VDD2.n115 B 0.011468f
C635 VDD2.n116 B 0.011806f
C636 VDD2.n117 B 0.011806f
C637 VDD2.n118 B 0.027107f
C638 VDD2.n119 B 0.027107f
C639 VDD2.n120 B 0.012143f
C640 VDD2.n121 B 0.011468f
C641 VDD2.n122 B 0.021343f
C642 VDD2.n123 B 0.021343f
C643 VDD2.n124 B 0.011468f
C644 VDD2.n125 B 0.012143f
C645 VDD2.n126 B 0.027107f
C646 VDD2.n127 B 0.027107f
C647 VDD2.n128 B 0.012143f
C648 VDD2.n129 B 0.011468f
C649 VDD2.n130 B 0.021343f
C650 VDD2.n131 B 0.021343f
C651 VDD2.n132 B 0.011468f
C652 VDD2.n133 B 0.012143f
C653 VDD2.n134 B 0.027107f
C654 VDD2.n135 B 0.057155f
C655 VDD2.n136 B 0.012143f
C656 VDD2.n137 B 0.011468f
C657 VDD2.n138 B 0.046416f
C658 VDD2.n139 B 0.046493f
C659 VDD2.n140 B 2.34319f
C660 VDD2.t0 B 0.214866f
C661 VDD2.t4 B 0.214866f
C662 VDD2.n141 B 1.92401f
C663 VN.t5 B 2.21352f
C664 VN.n0 B 0.86037f
C665 VN.n1 B 0.020737f
C666 VN.n2 B 0.027494f
C667 VN.n3 B 0.236111f
C668 VN.t1 B 2.21352f
C669 VN.t2 B 2.44438f
C670 VN.n4 B 0.811971f
C671 VN.n5 B 0.854971f
C672 VN.n6 B 0.038843f
C673 VN.n7 B 0.038843f
C674 VN.n8 B 0.020737f
C675 VN.n9 B 0.020737f
C676 VN.n10 B 0.020737f
C677 VN.n11 B 0.033314f
C678 VN.n12 B 0.038843f
C679 VN.n13 B 0.035007f
C680 VN.n14 B 0.033475f
C681 VN.n15 B 0.044074f
C682 VN.t3 B 2.21352f
C683 VN.n16 B 0.86037f
C684 VN.n17 B 0.020737f
C685 VN.n18 B 0.027494f
C686 VN.n19 B 0.236111f
C687 VN.t0 B 2.21352f
C688 VN.t4 B 2.44438f
C689 VN.n20 B 0.811971f
C690 VN.n21 B 0.854971f
C691 VN.n22 B 0.038843f
C692 VN.n23 B 0.038843f
C693 VN.n24 B 0.020737f
C694 VN.n25 B 0.020737f
C695 VN.n26 B 0.020737f
C696 VN.n27 B 0.033314f
C697 VN.n28 B 0.038843f
C698 VN.n29 B 0.035007f
C699 VN.n30 B 0.033475f
C700 VN.n31 B 1.22297f
.ends

