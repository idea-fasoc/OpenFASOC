* NGSPICE file created from diff_pair_sample_0401.ext - technology: sky130A

.subckt diff_pair_sample_0401 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t7 VN.t0 VDD2.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=6.4155 pd=33.68 as=2.71425 ps=16.78 w=16.45 l=2.31
X1 VDD2.t1 VN.t1 VTAIL.t6 B.t1 sky130_fd_pr__nfet_01v8 ad=2.71425 pd=16.78 as=6.4155 ps=33.68 w=16.45 l=2.31
X2 B.t17 B.t15 B.t16 B.t12 sky130_fd_pr__nfet_01v8 ad=6.4155 pd=33.68 as=0 ps=0 w=16.45 l=2.31
X3 VTAIL.t0 VP.t0 VDD1.t3 B.t0 sky130_fd_pr__nfet_01v8 ad=6.4155 pd=33.68 as=2.71425 ps=16.78 w=16.45 l=2.31
X4 VDD1.t2 VP.t1 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=2.71425 pd=16.78 as=6.4155 ps=33.68 w=16.45 l=2.31
X5 B.t14 B.t11 B.t13 B.t12 sky130_fd_pr__nfet_01v8 ad=6.4155 pd=33.68 as=0 ps=0 w=16.45 l=2.31
X6 VDD2.t3 VN.t2 VTAIL.t5 B.t3 sky130_fd_pr__nfet_01v8 ad=2.71425 pd=16.78 as=6.4155 ps=33.68 w=16.45 l=2.31
X7 B.t10 B.t8 B.t9 B.t5 sky130_fd_pr__nfet_01v8 ad=6.4155 pd=33.68 as=0 ps=0 w=16.45 l=2.31
X8 VTAIL.t4 VN.t3 VDD2.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=6.4155 pd=33.68 as=2.71425 ps=16.78 w=16.45 l=2.31
X9 B.t7 B.t4 B.t6 B.t5 sky130_fd_pr__nfet_01v8 ad=6.4155 pd=33.68 as=0 ps=0 w=16.45 l=2.31
X10 VDD1.t1 VP.t2 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=2.71425 pd=16.78 as=6.4155 ps=33.68 w=16.45 l=2.31
X11 VTAIL.t2 VP.t3 VDD1.t0 B.t2 sky130_fd_pr__nfet_01v8 ad=6.4155 pd=33.68 as=2.71425 ps=16.78 w=16.45 l=2.31
R0 VN.n0 VN.t3 208.026
R1 VN.n1 VN.t2 208.026
R2 VN.n0 VN.t1 207.371
R3 VN.n1 VN.t0 207.371
R4 VN VN.n1 54.613
R5 VN VN.n0 5.54102
R6 VDD2.n2 VDD2.n0 105.666
R7 VDD2.n2 VDD2.n1 60.9434
R8 VDD2.n1 VDD2.t2 1.20415
R9 VDD2.n1 VDD2.t3 1.20415
R10 VDD2.n0 VDD2.t0 1.20415
R11 VDD2.n0 VDD2.t1 1.20415
R12 VDD2 VDD2.n2 0.0586897
R13 VTAIL.n5 VTAIL.t0 45.4684
R14 VTAIL.n4 VTAIL.t5 45.4684
R15 VTAIL.n3 VTAIL.t7 45.4684
R16 VTAIL.n6 VTAIL.t1 45.4682
R17 VTAIL.n7 VTAIL.t6 45.4682
R18 VTAIL.n0 VTAIL.t4 45.4682
R19 VTAIL.n1 VTAIL.t3 45.4682
R20 VTAIL.n2 VTAIL.t2 45.4682
R21 VTAIL.n7 VTAIL.n6 28.8238
R22 VTAIL.n3 VTAIL.n2 28.8238
R23 VTAIL.n4 VTAIL.n3 2.27636
R24 VTAIL.n6 VTAIL.n5 2.27636
R25 VTAIL.n2 VTAIL.n1 2.27636
R26 VTAIL VTAIL.n0 1.19662
R27 VTAIL VTAIL.n7 1.08024
R28 VTAIL.n5 VTAIL.n4 0.470328
R29 VTAIL.n1 VTAIL.n0 0.470328
R30 B.n857 B.n856 585
R31 B.n858 B.n857 585
R32 B.n358 B.n120 585
R33 B.n357 B.n356 585
R34 B.n355 B.n354 585
R35 B.n353 B.n352 585
R36 B.n351 B.n350 585
R37 B.n349 B.n348 585
R38 B.n347 B.n346 585
R39 B.n345 B.n344 585
R40 B.n343 B.n342 585
R41 B.n341 B.n340 585
R42 B.n339 B.n338 585
R43 B.n337 B.n336 585
R44 B.n335 B.n334 585
R45 B.n333 B.n332 585
R46 B.n331 B.n330 585
R47 B.n329 B.n328 585
R48 B.n327 B.n326 585
R49 B.n325 B.n324 585
R50 B.n323 B.n322 585
R51 B.n321 B.n320 585
R52 B.n319 B.n318 585
R53 B.n317 B.n316 585
R54 B.n315 B.n314 585
R55 B.n313 B.n312 585
R56 B.n311 B.n310 585
R57 B.n309 B.n308 585
R58 B.n307 B.n306 585
R59 B.n305 B.n304 585
R60 B.n303 B.n302 585
R61 B.n301 B.n300 585
R62 B.n299 B.n298 585
R63 B.n297 B.n296 585
R64 B.n295 B.n294 585
R65 B.n293 B.n292 585
R66 B.n291 B.n290 585
R67 B.n289 B.n288 585
R68 B.n287 B.n286 585
R69 B.n285 B.n284 585
R70 B.n283 B.n282 585
R71 B.n281 B.n280 585
R72 B.n279 B.n278 585
R73 B.n277 B.n276 585
R74 B.n275 B.n274 585
R75 B.n273 B.n272 585
R76 B.n271 B.n270 585
R77 B.n269 B.n268 585
R78 B.n267 B.n266 585
R79 B.n265 B.n264 585
R80 B.n263 B.n262 585
R81 B.n261 B.n260 585
R82 B.n259 B.n258 585
R83 B.n257 B.n256 585
R84 B.n255 B.n254 585
R85 B.n253 B.n252 585
R86 B.n251 B.n250 585
R87 B.n249 B.n248 585
R88 B.n247 B.n246 585
R89 B.n245 B.n244 585
R90 B.n243 B.n242 585
R91 B.n241 B.n240 585
R92 B.n239 B.n238 585
R93 B.n237 B.n236 585
R94 B.n235 B.n234 585
R95 B.n232 B.n231 585
R96 B.n230 B.n229 585
R97 B.n228 B.n227 585
R98 B.n226 B.n225 585
R99 B.n224 B.n223 585
R100 B.n222 B.n221 585
R101 B.n220 B.n219 585
R102 B.n218 B.n217 585
R103 B.n216 B.n215 585
R104 B.n214 B.n213 585
R105 B.n212 B.n211 585
R106 B.n210 B.n209 585
R107 B.n208 B.n207 585
R108 B.n206 B.n205 585
R109 B.n204 B.n203 585
R110 B.n202 B.n201 585
R111 B.n200 B.n199 585
R112 B.n198 B.n197 585
R113 B.n196 B.n195 585
R114 B.n194 B.n193 585
R115 B.n192 B.n191 585
R116 B.n190 B.n189 585
R117 B.n188 B.n187 585
R118 B.n186 B.n185 585
R119 B.n184 B.n183 585
R120 B.n182 B.n181 585
R121 B.n180 B.n179 585
R122 B.n178 B.n177 585
R123 B.n176 B.n175 585
R124 B.n174 B.n173 585
R125 B.n172 B.n171 585
R126 B.n170 B.n169 585
R127 B.n168 B.n167 585
R128 B.n166 B.n165 585
R129 B.n164 B.n163 585
R130 B.n162 B.n161 585
R131 B.n160 B.n159 585
R132 B.n158 B.n157 585
R133 B.n156 B.n155 585
R134 B.n154 B.n153 585
R135 B.n152 B.n151 585
R136 B.n150 B.n149 585
R137 B.n148 B.n147 585
R138 B.n146 B.n145 585
R139 B.n144 B.n143 585
R140 B.n142 B.n141 585
R141 B.n140 B.n139 585
R142 B.n138 B.n137 585
R143 B.n136 B.n135 585
R144 B.n134 B.n133 585
R145 B.n132 B.n131 585
R146 B.n130 B.n129 585
R147 B.n128 B.n127 585
R148 B.n61 B.n60 585
R149 B.n861 B.n860 585
R150 B.n855 B.n121 585
R151 B.n121 B.n58 585
R152 B.n854 B.n57 585
R153 B.n865 B.n57 585
R154 B.n853 B.n56 585
R155 B.n866 B.n56 585
R156 B.n852 B.n55 585
R157 B.n867 B.n55 585
R158 B.n851 B.n850 585
R159 B.n850 B.n51 585
R160 B.n849 B.n50 585
R161 B.n873 B.n50 585
R162 B.n848 B.n49 585
R163 B.n874 B.n49 585
R164 B.n847 B.n48 585
R165 B.n875 B.n48 585
R166 B.n846 B.n845 585
R167 B.n845 B.n44 585
R168 B.n844 B.n43 585
R169 B.n881 B.n43 585
R170 B.n843 B.n42 585
R171 B.n882 B.n42 585
R172 B.n842 B.n41 585
R173 B.n883 B.n41 585
R174 B.n841 B.n840 585
R175 B.n840 B.n37 585
R176 B.n839 B.n36 585
R177 B.n889 B.n36 585
R178 B.n838 B.n35 585
R179 B.n890 B.n35 585
R180 B.n837 B.n34 585
R181 B.n891 B.n34 585
R182 B.n836 B.n835 585
R183 B.n835 B.n30 585
R184 B.n834 B.n29 585
R185 B.n897 B.n29 585
R186 B.n833 B.n28 585
R187 B.n898 B.n28 585
R188 B.n832 B.n27 585
R189 B.n899 B.n27 585
R190 B.n831 B.n830 585
R191 B.n830 B.n23 585
R192 B.n829 B.n22 585
R193 B.n905 B.n22 585
R194 B.n828 B.n21 585
R195 B.n906 B.n21 585
R196 B.n827 B.n20 585
R197 B.n907 B.n20 585
R198 B.n826 B.n825 585
R199 B.n825 B.n16 585
R200 B.n824 B.n15 585
R201 B.n913 B.n15 585
R202 B.n823 B.n14 585
R203 B.n914 B.n14 585
R204 B.n822 B.n13 585
R205 B.n915 B.n13 585
R206 B.n821 B.n820 585
R207 B.n820 B.n12 585
R208 B.n819 B.n818 585
R209 B.n819 B.n8 585
R210 B.n817 B.n7 585
R211 B.n922 B.n7 585
R212 B.n816 B.n6 585
R213 B.n923 B.n6 585
R214 B.n815 B.n5 585
R215 B.n924 B.n5 585
R216 B.n814 B.n813 585
R217 B.n813 B.n4 585
R218 B.n812 B.n359 585
R219 B.n812 B.n811 585
R220 B.n802 B.n360 585
R221 B.n361 B.n360 585
R222 B.n804 B.n803 585
R223 B.n805 B.n804 585
R224 B.n801 B.n365 585
R225 B.n369 B.n365 585
R226 B.n800 B.n799 585
R227 B.n799 B.n798 585
R228 B.n367 B.n366 585
R229 B.n368 B.n367 585
R230 B.n791 B.n790 585
R231 B.n792 B.n791 585
R232 B.n789 B.n374 585
R233 B.n374 B.n373 585
R234 B.n788 B.n787 585
R235 B.n787 B.n786 585
R236 B.n376 B.n375 585
R237 B.n377 B.n376 585
R238 B.n779 B.n778 585
R239 B.n780 B.n779 585
R240 B.n777 B.n381 585
R241 B.n385 B.n381 585
R242 B.n776 B.n775 585
R243 B.n775 B.n774 585
R244 B.n383 B.n382 585
R245 B.n384 B.n383 585
R246 B.n767 B.n766 585
R247 B.n768 B.n767 585
R248 B.n765 B.n390 585
R249 B.n390 B.n389 585
R250 B.n764 B.n763 585
R251 B.n763 B.n762 585
R252 B.n392 B.n391 585
R253 B.n393 B.n392 585
R254 B.n755 B.n754 585
R255 B.n756 B.n755 585
R256 B.n753 B.n398 585
R257 B.n398 B.n397 585
R258 B.n752 B.n751 585
R259 B.n751 B.n750 585
R260 B.n400 B.n399 585
R261 B.n401 B.n400 585
R262 B.n743 B.n742 585
R263 B.n744 B.n743 585
R264 B.n741 B.n406 585
R265 B.n406 B.n405 585
R266 B.n740 B.n739 585
R267 B.n739 B.n738 585
R268 B.n408 B.n407 585
R269 B.n409 B.n408 585
R270 B.n731 B.n730 585
R271 B.n732 B.n731 585
R272 B.n729 B.n414 585
R273 B.n414 B.n413 585
R274 B.n728 B.n727 585
R275 B.n727 B.n726 585
R276 B.n416 B.n415 585
R277 B.n417 B.n416 585
R278 B.n722 B.n721 585
R279 B.n420 B.n419 585
R280 B.n718 B.n717 585
R281 B.n719 B.n718 585
R282 B.n716 B.n479 585
R283 B.n715 B.n714 585
R284 B.n713 B.n712 585
R285 B.n711 B.n710 585
R286 B.n709 B.n708 585
R287 B.n707 B.n706 585
R288 B.n705 B.n704 585
R289 B.n703 B.n702 585
R290 B.n701 B.n700 585
R291 B.n699 B.n698 585
R292 B.n697 B.n696 585
R293 B.n695 B.n694 585
R294 B.n693 B.n692 585
R295 B.n691 B.n690 585
R296 B.n689 B.n688 585
R297 B.n687 B.n686 585
R298 B.n685 B.n684 585
R299 B.n683 B.n682 585
R300 B.n681 B.n680 585
R301 B.n679 B.n678 585
R302 B.n677 B.n676 585
R303 B.n675 B.n674 585
R304 B.n673 B.n672 585
R305 B.n671 B.n670 585
R306 B.n669 B.n668 585
R307 B.n667 B.n666 585
R308 B.n665 B.n664 585
R309 B.n663 B.n662 585
R310 B.n661 B.n660 585
R311 B.n659 B.n658 585
R312 B.n657 B.n656 585
R313 B.n655 B.n654 585
R314 B.n653 B.n652 585
R315 B.n651 B.n650 585
R316 B.n649 B.n648 585
R317 B.n647 B.n646 585
R318 B.n645 B.n644 585
R319 B.n643 B.n642 585
R320 B.n641 B.n640 585
R321 B.n639 B.n638 585
R322 B.n637 B.n636 585
R323 B.n635 B.n634 585
R324 B.n633 B.n632 585
R325 B.n631 B.n630 585
R326 B.n629 B.n628 585
R327 B.n627 B.n626 585
R328 B.n625 B.n624 585
R329 B.n623 B.n622 585
R330 B.n621 B.n620 585
R331 B.n619 B.n618 585
R332 B.n617 B.n616 585
R333 B.n615 B.n614 585
R334 B.n613 B.n612 585
R335 B.n611 B.n610 585
R336 B.n609 B.n608 585
R337 B.n607 B.n606 585
R338 B.n605 B.n604 585
R339 B.n603 B.n602 585
R340 B.n601 B.n600 585
R341 B.n599 B.n598 585
R342 B.n597 B.n596 585
R343 B.n594 B.n593 585
R344 B.n592 B.n591 585
R345 B.n590 B.n589 585
R346 B.n588 B.n587 585
R347 B.n586 B.n585 585
R348 B.n584 B.n583 585
R349 B.n582 B.n581 585
R350 B.n580 B.n579 585
R351 B.n578 B.n577 585
R352 B.n576 B.n575 585
R353 B.n574 B.n573 585
R354 B.n572 B.n571 585
R355 B.n570 B.n569 585
R356 B.n568 B.n567 585
R357 B.n566 B.n565 585
R358 B.n564 B.n563 585
R359 B.n562 B.n561 585
R360 B.n560 B.n559 585
R361 B.n558 B.n557 585
R362 B.n556 B.n555 585
R363 B.n554 B.n553 585
R364 B.n552 B.n551 585
R365 B.n550 B.n549 585
R366 B.n548 B.n547 585
R367 B.n546 B.n545 585
R368 B.n544 B.n543 585
R369 B.n542 B.n541 585
R370 B.n540 B.n539 585
R371 B.n538 B.n537 585
R372 B.n536 B.n535 585
R373 B.n534 B.n533 585
R374 B.n532 B.n531 585
R375 B.n530 B.n529 585
R376 B.n528 B.n527 585
R377 B.n526 B.n525 585
R378 B.n524 B.n523 585
R379 B.n522 B.n521 585
R380 B.n520 B.n519 585
R381 B.n518 B.n517 585
R382 B.n516 B.n515 585
R383 B.n514 B.n513 585
R384 B.n512 B.n511 585
R385 B.n510 B.n509 585
R386 B.n508 B.n507 585
R387 B.n506 B.n505 585
R388 B.n504 B.n503 585
R389 B.n502 B.n501 585
R390 B.n500 B.n499 585
R391 B.n498 B.n497 585
R392 B.n496 B.n495 585
R393 B.n494 B.n493 585
R394 B.n492 B.n491 585
R395 B.n490 B.n489 585
R396 B.n488 B.n487 585
R397 B.n486 B.n485 585
R398 B.n723 B.n418 585
R399 B.n418 B.n417 585
R400 B.n725 B.n724 585
R401 B.n726 B.n725 585
R402 B.n412 B.n411 585
R403 B.n413 B.n412 585
R404 B.n734 B.n733 585
R405 B.n733 B.n732 585
R406 B.n735 B.n410 585
R407 B.n410 B.n409 585
R408 B.n737 B.n736 585
R409 B.n738 B.n737 585
R410 B.n404 B.n403 585
R411 B.n405 B.n404 585
R412 B.n746 B.n745 585
R413 B.n745 B.n744 585
R414 B.n747 B.n402 585
R415 B.n402 B.n401 585
R416 B.n749 B.n748 585
R417 B.n750 B.n749 585
R418 B.n396 B.n395 585
R419 B.n397 B.n396 585
R420 B.n758 B.n757 585
R421 B.n757 B.n756 585
R422 B.n759 B.n394 585
R423 B.n394 B.n393 585
R424 B.n761 B.n760 585
R425 B.n762 B.n761 585
R426 B.n388 B.n387 585
R427 B.n389 B.n388 585
R428 B.n770 B.n769 585
R429 B.n769 B.n768 585
R430 B.n771 B.n386 585
R431 B.n386 B.n384 585
R432 B.n773 B.n772 585
R433 B.n774 B.n773 585
R434 B.n380 B.n379 585
R435 B.n385 B.n380 585
R436 B.n782 B.n781 585
R437 B.n781 B.n780 585
R438 B.n783 B.n378 585
R439 B.n378 B.n377 585
R440 B.n785 B.n784 585
R441 B.n786 B.n785 585
R442 B.n372 B.n371 585
R443 B.n373 B.n372 585
R444 B.n794 B.n793 585
R445 B.n793 B.n792 585
R446 B.n795 B.n370 585
R447 B.n370 B.n368 585
R448 B.n797 B.n796 585
R449 B.n798 B.n797 585
R450 B.n364 B.n363 585
R451 B.n369 B.n364 585
R452 B.n807 B.n806 585
R453 B.n806 B.n805 585
R454 B.n808 B.n362 585
R455 B.n362 B.n361 585
R456 B.n810 B.n809 585
R457 B.n811 B.n810 585
R458 B.n3 B.n0 585
R459 B.n4 B.n3 585
R460 B.n921 B.n1 585
R461 B.n922 B.n921 585
R462 B.n920 B.n919 585
R463 B.n920 B.n8 585
R464 B.n918 B.n9 585
R465 B.n12 B.n9 585
R466 B.n917 B.n916 585
R467 B.n916 B.n915 585
R468 B.n11 B.n10 585
R469 B.n914 B.n11 585
R470 B.n912 B.n911 585
R471 B.n913 B.n912 585
R472 B.n910 B.n17 585
R473 B.n17 B.n16 585
R474 B.n909 B.n908 585
R475 B.n908 B.n907 585
R476 B.n19 B.n18 585
R477 B.n906 B.n19 585
R478 B.n904 B.n903 585
R479 B.n905 B.n904 585
R480 B.n902 B.n24 585
R481 B.n24 B.n23 585
R482 B.n901 B.n900 585
R483 B.n900 B.n899 585
R484 B.n26 B.n25 585
R485 B.n898 B.n26 585
R486 B.n896 B.n895 585
R487 B.n897 B.n896 585
R488 B.n894 B.n31 585
R489 B.n31 B.n30 585
R490 B.n893 B.n892 585
R491 B.n892 B.n891 585
R492 B.n33 B.n32 585
R493 B.n890 B.n33 585
R494 B.n888 B.n887 585
R495 B.n889 B.n888 585
R496 B.n886 B.n38 585
R497 B.n38 B.n37 585
R498 B.n885 B.n884 585
R499 B.n884 B.n883 585
R500 B.n40 B.n39 585
R501 B.n882 B.n40 585
R502 B.n880 B.n879 585
R503 B.n881 B.n880 585
R504 B.n878 B.n45 585
R505 B.n45 B.n44 585
R506 B.n877 B.n876 585
R507 B.n876 B.n875 585
R508 B.n47 B.n46 585
R509 B.n874 B.n47 585
R510 B.n872 B.n871 585
R511 B.n873 B.n872 585
R512 B.n870 B.n52 585
R513 B.n52 B.n51 585
R514 B.n869 B.n868 585
R515 B.n868 B.n867 585
R516 B.n54 B.n53 585
R517 B.n866 B.n54 585
R518 B.n864 B.n863 585
R519 B.n865 B.n864 585
R520 B.n862 B.n59 585
R521 B.n59 B.n58 585
R522 B.n925 B.n924 585
R523 B.n923 B.n2 585
R524 B.n860 B.n59 482.89
R525 B.n857 B.n121 482.89
R526 B.n485 B.n416 482.89
R527 B.n721 B.n418 482.89
R528 B.n125 B.t4 379.185
R529 B.n122 B.t8 379.185
R530 B.n483 B.t11 379.185
R531 B.n480 B.t15 379.185
R532 B.n858 B.n119 256.663
R533 B.n858 B.n118 256.663
R534 B.n858 B.n117 256.663
R535 B.n858 B.n116 256.663
R536 B.n858 B.n115 256.663
R537 B.n858 B.n114 256.663
R538 B.n858 B.n113 256.663
R539 B.n858 B.n112 256.663
R540 B.n858 B.n111 256.663
R541 B.n858 B.n110 256.663
R542 B.n858 B.n109 256.663
R543 B.n858 B.n108 256.663
R544 B.n858 B.n107 256.663
R545 B.n858 B.n106 256.663
R546 B.n858 B.n105 256.663
R547 B.n858 B.n104 256.663
R548 B.n858 B.n103 256.663
R549 B.n858 B.n102 256.663
R550 B.n858 B.n101 256.663
R551 B.n858 B.n100 256.663
R552 B.n858 B.n99 256.663
R553 B.n858 B.n98 256.663
R554 B.n858 B.n97 256.663
R555 B.n858 B.n96 256.663
R556 B.n858 B.n95 256.663
R557 B.n858 B.n94 256.663
R558 B.n858 B.n93 256.663
R559 B.n858 B.n92 256.663
R560 B.n858 B.n91 256.663
R561 B.n858 B.n90 256.663
R562 B.n858 B.n89 256.663
R563 B.n858 B.n88 256.663
R564 B.n858 B.n87 256.663
R565 B.n858 B.n86 256.663
R566 B.n858 B.n85 256.663
R567 B.n858 B.n84 256.663
R568 B.n858 B.n83 256.663
R569 B.n858 B.n82 256.663
R570 B.n858 B.n81 256.663
R571 B.n858 B.n80 256.663
R572 B.n858 B.n79 256.663
R573 B.n858 B.n78 256.663
R574 B.n858 B.n77 256.663
R575 B.n858 B.n76 256.663
R576 B.n858 B.n75 256.663
R577 B.n858 B.n74 256.663
R578 B.n858 B.n73 256.663
R579 B.n858 B.n72 256.663
R580 B.n858 B.n71 256.663
R581 B.n858 B.n70 256.663
R582 B.n858 B.n69 256.663
R583 B.n858 B.n68 256.663
R584 B.n858 B.n67 256.663
R585 B.n858 B.n66 256.663
R586 B.n858 B.n65 256.663
R587 B.n858 B.n64 256.663
R588 B.n858 B.n63 256.663
R589 B.n858 B.n62 256.663
R590 B.n859 B.n858 256.663
R591 B.n720 B.n719 256.663
R592 B.n719 B.n421 256.663
R593 B.n719 B.n422 256.663
R594 B.n719 B.n423 256.663
R595 B.n719 B.n424 256.663
R596 B.n719 B.n425 256.663
R597 B.n719 B.n426 256.663
R598 B.n719 B.n427 256.663
R599 B.n719 B.n428 256.663
R600 B.n719 B.n429 256.663
R601 B.n719 B.n430 256.663
R602 B.n719 B.n431 256.663
R603 B.n719 B.n432 256.663
R604 B.n719 B.n433 256.663
R605 B.n719 B.n434 256.663
R606 B.n719 B.n435 256.663
R607 B.n719 B.n436 256.663
R608 B.n719 B.n437 256.663
R609 B.n719 B.n438 256.663
R610 B.n719 B.n439 256.663
R611 B.n719 B.n440 256.663
R612 B.n719 B.n441 256.663
R613 B.n719 B.n442 256.663
R614 B.n719 B.n443 256.663
R615 B.n719 B.n444 256.663
R616 B.n719 B.n445 256.663
R617 B.n719 B.n446 256.663
R618 B.n719 B.n447 256.663
R619 B.n719 B.n448 256.663
R620 B.n719 B.n449 256.663
R621 B.n719 B.n450 256.663
R622 B.n719 B.n451 256.663
R623 B.n719 B.n452 256.663
R624 B.n719 B.n453 256.663
R625 B.n719 B.n454 256.663
R626 B.n719 B.n455 256.663
R627 B.n719 B.n456 256.663
R628 B.n719 B.n457 256.663
R629 B.n719 B.n458 256.663
R630 B.n719 B.n459 256.663
R631 B.n719 B.n460 256.663
R632 B.n719 B.n461 256.663
R633 B.n719 B.n462 256.663
R634 B.n719 B.n463 256.663
R635 B.n719 B.n464 256.663
R636 B.n719 B.n465 256.663
R637 B.n719 B.n466 256.663
R638 B.n719 B.n467 256.663
R639 B.n719 B.n468 256.663
R640 B.n719 B.n469 256.663
R641 B.n719 B.n470 256.663
R642 B.n719 B.n471 256.663
R643 B.n719 B.n472 256.663
R644 B.n719 B.n473 256.663
R645 B.n719 B.n474 256.663
R646 B.n719 B.n475 256.663
R647 B.n719 B.n476 256.663
R648 B.n719 B.n477 256.663
R649 B.n719 B.n478 256.663
R650 B.n927 B.n926 256.663
R651 B.n127 B.n61 163.367
R652 B.n131 B.n130 163.367
R653 B.n135 B.n134 163.367
R654 B.n139 B.n138 163.367
R655 B.n143 B.n142 163.367
R656 B.n147 B.n146 163.367
R657 B.n151 B.n150 163.367
R658 B.n155 B.n154 163.367
R659 B.n159 B.n158 163.367
R660 B.n163 B.n162 163.367
R661 B.n167 B.n166 163.367
R662 B.n171 B.n170 163.367
R663 B.n175 B.n174 163.367
R664 B.n179 B.n178 163.367
R665 B.n183 B.n182 163.367
R666 B.n187 B.n186 163.367
R667 B.n191 B.n190 163.367
R668 B.n195 B.n194 163.367
R669 B.n199 B.n198 163.367
R670 B.n203 B.n202 163.367
R671 B.n207 B.n206 163.367
R672 B.n211 B.n210 163.367
R673 B.n215 B.n214 163.367
R674 B.n219 B.n218 163.367
R675 B.n223 B.n222 163.367
R676 B.n227 B.n226 163.367
R677 B.n231 B.n230 163.367
R678 B.n236 B.n235 163.367
R679 B.n240 B.n239 163.367
R680 B.n244 B.n243 163.367
R681 B.n248 B.n247 163.367
R682 B.n252 B.n251 163.367
R683 B.n256 B.n255 163.367
R684 B.n260 B.n259 163.367
R685 B.n264 B.n263 163.367
R686 B.n268 B.n267 163.367
R687 B.n272 B.n271 163.367
R688 B.n276 B.n275 163.367
R689 B.n280 B.n279 163.367
R690 B.n284 B.n283 163.367
R691 B.n288 B.n287 163.367
R692 B.n292 B.n291 163.367
R693 B.n296 B.n295 163.367
R694 B.n300 B.n299 163.367
R695 B.n304 B.n303 163.367
R696 B.n308 B.n307 163.367
R697 B.n312 B.n311 163.367
R698 B.n316 B.n315 163.367
R699 B.n320 B.n319 163.367
R700 B.n324 B.n323 163.367
R701 B.n328 B.n327 163.367
R702 B.n332 B.n331 163.367
R703 B.n336 B.n335 163.367
R704 B.n340 B.n339 163.367
R705 B.n344 B.n343 163.367
R706 B.n348 B.n347 163.367
R707 B.n352 B.n351 163.367
R708 B.n356 B.n355 163.367
R709 B.n857 B.n120 163.367
R710 B.n727 B.n416 163.367
R711 B.n727 B.n414 163.367
R712 B.n731 B.n414 163.367
R713 B.n731 B.n408 163.367
R714 B.n739 B.n408 163.367
R715 B.n739 B.n406 163.367
R716 B.n743 B.n406 163.367
R717 B.n743 B.n400 163.367
R718 B.n751 B.n400 163.367
R719 B.n751 B.n398 163.367
R720 B.n755 B.n398 163.367
R721 B.n755 B.n392 163.367
R722 B.n763 B.n392 163.367
R723 B.n763 B.n390 163.367
R724 B.n767 B.n390 163.367
R725 B.n767 B.n383 163.367
R726 B.n775 B.n383 163.367
R727 B.n775 B.n381 163.367
R728 B.n779 B.n381 163.367
R729 B.n779 B.n376 163.367
R730 B.n787 B.n376 163.367
R731 B.n787 B.n374 163.367
R732 B.n791 B.n374 163.367
R733 B.n791 B.n367 163.367
R734 B.n799 B.n367 163.367
R735 B.n799 B.n365 163.367
R736 B.n804 B.n365 163.367
R737 B.n804 B.n360 163.367
R738 B.n812 B.n360 163.367
R739 B.n813 B.n812 163.367
R740 B.n813 B.n5 163.367
R741 B.n6 B.n5 163.367
R742 B.n7 B.n6 163.367
R743 B.n819 B.n7 163.367
R744 B.n820 B.n819 163.367
R745 B.n820 B.n13 163.367
R746 B.n14 B.n13 163.367
R747 B.n15 B.n14 163.367
R748 B.n825 B.n15 163.367
R749 B.n825 B.n20 163.367
R750 B.n21 B.n20 163.367
R751 B.n22 B.n21 163.367
R752 B.n830 B.n22 163.367
R753 B.n830 B.n27 163.367
R754 B.n28 B.n27 163.367
R755 B.n29 B.n28 163.367
R756 B.n835 B.n29 163.367
R757 B.n835 B.n34 163.367
R758 B.n35 B.n34 163.367
R759 B.n36 B.n35 163.367
R760 B.n840 B.n36 163.367
R761 B.n840 B.n41 163.367
R762 B.n42 B.n41 163.367
R763 B.n43 B.n42 163.367
R764 B.n845 B.n43 163.367
R765 B.n845 B.n48 163.367
R766 B.n49 B.n48 163.367
R767 B.n50 B.n49 163.367
R768 B.n850 B.n50 163.367
R769 B.n850 B.n55 163.367
R770 B.n56 B.n55 163.367
R771 B.n57 B.n56 163.367
R772 B.n121 B.n57 163.367
R773 B.n718 B.n420 163.367
R774 B.n718 B.n479 163.367
R775 B.n714 B.n713 163.367
R776 B.n710 B.n709 163.367
R777 B.n706 B.n705 163.367
R778 B.n702 B.n701 163.367
R779 B.n698 B.n697 163.367
R780 B.n694 B.n693 163.367
R781 B.n690 B.n689 163.367
R782 B.n686 B.n685 163.367
R783 B.n682 B.n681 163.367
R784 B.n678 B.n677 163.367
R785 B.n674 B.n673 163.367
R786 B.n670 B.n669 163.367
R787 B.n666 B.n665 163.367
R788 B.n662 B.n661 163.367
R789 B.n658 B.n657 163.367
R790 B.n654 B.n653 163.367
R791 B.n650 B.n649 163.367
R792 B.n646 B.n645 163.367
R793 B.n642 B.n641 163.367
R794 B.n638 B.n637 163.367
R795 B.n634 B.n633 163.367
R796 B.n630 B.n629 163.367
R797 B.n626 B.n625 163.367
R798 B.n622 B.n621 163.367
R799 B.n618 B.n617 163.367
R800 B.n614 B.n613 163.367
R801 B.n610 B.n609 163.367
R802 B.n606 B.n605 163.367
R803 B.n602 B.n601 163.367
R804 B.n598 B.n597 163.367
R805 B.n593 B.n592 163.367
R806 B.n589 B.n588 163.367
R807 B.n585 B.n584 163.367
R808 B.n581 B.n580 163.367
R809 B.n577 B.n576 163.367
R810 B.n573 B.n572 163.367
R811 B.n569 B.n568 163.367
R812 B.n565 B.n564 163.367
R813 B.n561 B.n560 163.367
R814 B.n557 B.n556 163.367
R815 B.n553 B.n552 163.367
R816 B.n549 B.n548 163.367
R817 B.n545 B.n544 163.367
R818 B.n541 B.n540 163.367
R819 B.n537 B.n536 163.367
R820 B.n533 B.n532 163.367
R821 B.n529 B.n528 163.367
R822 B.n525 B.n524 163.367
R823 B.n521 B.n520 163.367
R824 B.n517 B.n516 163.367
R825 B.n513 B.n512 163.367
R826 B.n509 B.n508 163.367
R827 B.n505 B.n504 163.367
R828 B.n501 B.n500 163.367
R829 B.n497 B.n496 163.367
R830 B.n493 B.n492 163.367
R831 B.n489 B.n488 163.367
R832 B.n725 B.n418 163.367
R833 B.n725 B.n412 163.367
R834 B.n733 B.n412 163.367
R835 B.n733 B.n410 163.367
R836 B.n737 B.n410 163.367
R837 B.n737 B.n404 163.367
R838 B.n745 B.n404 163.367
R839 B.n745 B.n402 163.367
R840 B.n749 B.n402 163.367
R841 B.n749 B.n396 163.367
R842 B.n757 B.n396 163.367
R843 B.n757 B.n394 163.367
R844 B.n761 B.n394 163.367
R845 B.n761 B.n388 163.367
R846 B.n769 B.n388 163.367
R847 B.n769 B.n386 163.367
R848 B.n773 B.n386 163.367
R849 B.n773 B.n380 163.367
R850 B.n781 B.n380 163.367
R851 B.n781 B.n378 163.367
R852 B.n785 B.n378 163.367
R853 B.n785 B.n372 163.367
R854 B.n793 B.n372 163.367
R855 B.n793 B.n370 163.367
R856 B.n797 B.n370 163.367
R857 B.n797 B.n364 163.367
R858 B.n806 B.n364 163.367
R859 B.n806 B.n362 163.367
R860 B.n810 B.n362 163.367
R861 B.n810 B.n3 163.367
R862 B.n925 B.n3 163.367
R863 B.n921 B.n2 163.367
R864 B.n921 B.n920 163.367
R865 B.n920 B.n9 163.367
R866 B.n916 B.n9 163.367
R867 B.n916 B.n11 163.367
R868 B.n912 B.n11 163.367
R869 B.n912 B.n17 163.367
R870 B.n908 B.n17 163.367
R871 B.n908 B.n19 163.367
R872 B.n904 B.n19 163.367
R873 B.n904 B.n24 163.367
R874 B.n900 B.n24 163.367
R875 B.n900 B.n26 163.367
R876 B.n896 B.n26 163.367
R877 B.n896 B.n31 163.367
R878 B.n892 B.n31 163.367
R879 B.n892 B.n33 163.367
R880 B.n888 B.n33 163.367
R881 B.n888 B.n38 163.367
R882 B.n884 B.n38 163.367
R883 B.n884 B.n40 163.367
R884 B.n880 B.n40 163.367
R885 B.n880 B.n45 163.367
R886 B.n876 B.n45 163.367
R887 B.n876 B.n47 163.367
R888 B.n872 B.n47 163.367
R889 B.n872 B.n52 163.367
R890 B.n868 B.n52 163.367
R891 B.n868 B.n54 163.367
R892 B.n864 B.n54 163.367
R893 B.n864 B.n59 163.367
R894 B.n122 B.t9 121.072
R895 B.n483 B.t14 121.072
R896 B.n125 B.t6 121.049
R897 B.n480 B.t17 121.049
R898 B.n860 B.n859 71.676
R899 B.n127 B.n62 71.676
R900 B.n131 B.n63 71.676
R901 B.n135 B.n64 71.676
R902 B.n139 B.n65 71.676
R903 B.n143 B.n66 71.676
R904 B.n147 B.n67 71.676
R905 B.n151 B.n68 71.676
R906 B.n155 B.n69 71.676
R907 B.n159 B.n70 71.676
R908 B.n163 B.n71 71.676
R909 B.n167 B.n72 71.676
R910 B.n171 B.n73 71.676
R911 B.n175 B.n74 71.676
R912 B.n179 B.n75 71.676
R913 B.n183 B.n76 71.676
R914 B.n187 B.n77 71.676
R915 B.n191 B.n78 71.676
R916 B.n195 B.n79 71.676
R917 B.n199 B.n80 71.676
R918 B.n203 B.n81 71.676
R919 B.n207 B.n82 71.676
R920 B.n211 B.n83 71.676
R921 B.n215 B.n84 71.676
R922 B.n219 B.n85 71.676
R923 B.n223 B.n86 71.676
R924 B.n227 B.n87 71.676
R925 B.n231 B.n88 71.676
R926 B.n236 B.n89 71.676
R927 B.n240 B.n90 71.676
R928 B.n244 B.n91 71.676
R929 B.n248 B.n92 71.676
R930 B.n252 B.n93 71.676
R931 B.n256 B.n94 71.676
R932 B.n260 B.n95 71.676
R933 B.n264 B.n96 71.676
R934 B.n268 B.n97 71.676
R935 B.n272 B.n98 71.676
R936 B.n276 B.n99 71.676
R937 B.n280 B.n100 71.676
R938 B.n284 B.n101 71.676
R939 B.n288 B.n102 71.676
R940 B.n292 B.n103 71.676
R941 B.n296 B.n104 71.676
R942 B.n300 B.n105 71.676
R943 B.n304 B.n106 71.676
R944 B.n308 B.n107 71.676
R945 B.n312 B.n108 71.676
R946 B.n316 B.n109 71.676
R947 B.n320 B.n110 71.676
R948 B.n324 B.n111 71.676
R949 B.n328 B.n112 71.676
R950 B.n332 B.n113 71.676
R951 B.n336 B.n114 71.676
R952 B.n340 B.n115 71.676
R953 B.n344 B.n116 71.676
R954 B.n348 B.n117 71.676
R955 B.n352 B.n118 71.676
R956 B.n356 B.n119 71.676
R957 B.n120 B.n119 71.676
R958 B.n355 B.n118 71.676
R959 B.n351 B.n117 71.676
R960 B.n347 B.n116 71.676
R961 B.n343 B.n115 71.676
R962 B.n339 B.n114 71.676
R963 B.n335 B.n113 71.676
R964 B.n331 B.n112 71.676
R965 B.n327 B.n111 71.676
R966 B.n323 B.n110 71.676
R967 B.n319 B.n109 71.676
R968 B.n315 B.n108 71.676
R969 B.n311 B.n107 71.676
R970 B.n307 B.n106 71.676
R971 B.n303 B.n105 71.676
R972 B.n299 B.n104 71.676
R973 B.n295 B.n103 71.676
R974 B.n291 B.n102 71.676
R975 B.n287 B.n101 71.676
R976 B.n283 B.n100 71.676
R977 B.n279 B.n99 71.676
R978 B.n275 B.n98 71.676
R979 B.n271 B.n97 71.676
R980 B.n267 B.n96 71.676
R981 B.n263 B.n95 71.676
R982 B.n259 B.n94 71.676
R983 B.n255 B.n93 71.676
R984 B.n251 B.n92 71.676
R985 B.n247 B.n91 71.676
R986 B.n243 B.n90 71.676
R987 B.n239 B.n89 71.676
R988 B.n235 B.n88 71.676
R989 B.n230 B.n87 71.676
R990 B.n226 B.n86 71.676
R991 B.n222 B.n85 71.676
R992 B.n218 B.n84 71.676
R993 B.n214 B.n83 71.676
R994 B.n210 B.n82 71.676
R995 B.n206 B.n81 71.676
R996 B.n202 B.n80 71.676
R997 B.n198 B.n79 71.676
R998 B.n194 B.n78 71.676
R999 B.n190 B.n77 71.676
R1000 B.n186 B.n76 71.676
R1001 B.n182 B.n75 71.676
R1002 B.n178 B.n74 71.676
R1003 B.n174 B.n73 71.676
R1004 B.n170 B.n72 71.676
R1005 B.n166 B.n71 71.676
R1006 B.n162 B.n70 71.676
R1007 B.n158 B.n69 71.676
R1008 B.n154 B.n68 71.676
R1009 B.n150 B.n67 71.676
R1010 B.n146 B.n66 71.676
R1011 B.n142 B.n65 71.676
R1012 B.n138 B.n64 71.676
R1013 B.n134 B.n63 71.676
R1014 B.n130 B.n62 71.676
R1015 B.n859 B.n61 71.676
R1016 B.n721 B.n720 71.676
R1017 B.n479 B.n421 71.676
R1018 B.n713 B.n422 71.676
R1019 B.n709 B.n423 71.676
R1020 B.n705 B.n424 71.676
R1021 B.n701 B.n425 71.676
R1022 B.n697 B.n426 71.676
R1023 B.n693 B.n427 71.676
R1024 B.n689 B.n428 71.676
R1025 B.n685 B.n429 71.676
R1026 B.n681 B.n430 71.676
R1027 B.n677 B.n431 71.676
R1028 B.n673 B.n432 71.676
R1029 B.n669 B.n433 71.676
R1030 B.n665 B.n434 71.676
R1031 B.n661 B.n435 71.676
R1032 B.n657 B.n436 71.676
R1033 B.n653 B.n437 71.676
R1034 B.n649 B.n438 71.676
R1035 B.n645 B.n439 71.676
R1036 B.n641 B.n440 71.676
R1037 B.n637 B.n441 71.676
R1038 B.n633 B.n442 71.676
R1039 B.n629 B.n443 71.676
R1040 B.n625 B.n444 71.676
R1041 B.n621 B.n445 71.676
R1042 B.n617 B.n446 71.676
R1043 B.n613 B.n447 71.676
R1044 B.n609 B.n448 71.676
R1045 B.n605 B.n449 71.676
R1046 B.n601 B.n450 71.676
R1047 B.n597 B.n451 71.676
R1048 B.n592 B.n452 71.676
R1049 B.n588 B.n453 71.676
R1050 B.n584 B.n454 71.676
R1051 B.n580 B.n455 71.676
R1052 B.n576 B.n456 71.676
R1053 B.n572 B.n457 71.676
R1054 B.n568 B.n458 71.676
R1055 B.n564 B.n459 71.676
R1056 B.n560 B.n460 71.676
R1057 B.n556 B.n461 71.676
R1058 B.n552 B.n462 71.676
R1059 B.n548 B.n463 71.676
R1060 B.n544 B.n464 71.676
R1061 B.n540 B.n465 71.676
R1062 B.n536 B.n466 71.676
R1063 B.n532 B.n467 71.676
R1064 B.n528 B.n468 71.676
R1065 B.n524 B.n469 71.676
R1066 B.n520 B.n470 71.676
R1067 B.n516 B.n471 71.676
R1068 B.n512 B.n472 71.676
R1069 B.n508 B.n473 71.676
R1070 B.n504 B.n474 71.676
R1071 B.n500 B.n475 71.676
R1072 B.n496 B.n476 71.676
R1073 B.n492 B.n477 71.676
R1074 B.n488 B.n478 71.676
R1075 B.n720 B.n420 71.676
R1076 B.n714 B.n421 71.676
R1077 B.n710 B.n422 71.676
R1078 B.n706 B.n423 71.676
R1079 B.n702 B.n424 71.676
R1080 B.n698 B.n425 71.676
R1081 B.n694 B.n426 71.676
R1082 B.n690 B.n427 71.676
R1083 B.n686 B.n428 71.676
R1084 B.n682 B.n429 71.676
R1085 B.n678 B.n430 71.676
R1086 B.n674 B.n431 71.676
R1087 B.n670 B.n432 71.676
R1088 B.n666 B.n433 71.676
R1089 B.n662 B.n434 71.676
R1090 B.n658 B.n435 71.676
R1091 B.n654 B.n436 71.676
R1092 B.n650 B.n437 71.676
R1093 B.n646 B.n438 71.676
R1094 B.n642 B.n439 71.676
R1095 B.n638 B.n440 71.676
R1096 B.n634 B.n441 71.676
R1097 B.n630 B.n442 71.676
R1098 B.n626 B.n443 71.676
R1099 B.n622 B.n444 71.676
R1100 B.n618 B.n445 71.676
R1101 B.n614 B.n446 71.676
R1102 B.n610 B.n447 71.676
R1103 B.n606 B.n448 71.676
R1104 B.n602 B.n449 71.676
R1105 B.n598 B.n450 71.676
R1106 B.n593 B.n451 71.676
R1107 B.n589 B.n452 71.676
R1108 B.n585 B.n453 71.676
R1109 B.n581 B.n454 71.676
R1110 B.n577 B.n455 71.676
R1111 B.n573 B.n456 71.676
R1112 B.n569 B.n457 71.676
R1113 B.n565 B.n458 71.676
R1114 B.n561 B.n459 71.676
R1115 B.n557 B.n460 71.676
R1116 B.n553 B.n461 71.676
R1117 B.n549 B.n462 71.676
R1118 B.n545 B.n463 71.676
R1119 B.n541 B.n464 71.676
R1120 B.n537 B.n465 71.676
R1121 B.n533 B.n466 71.676
R1122 B.n529 B.n467 71.676
R1123 B.n525 B.n468 71.676
R1124 B.n521 B.n469 71.676
R1125 B.n517 B.n470 71.676
R1126 B.n513 B.n471 71.676
R1127 B.n509 B.n472 71.676
R1128 B.n505 B.n473 71.676
R1129 B.n501 B.n474 71.676
R1130 B.n497 B.n475 71.676
R1131 B.n493 B.n476 71.676
R1132 B.n489 B.n477 71.676
R1133 B.n485 B.n478 71.676
R1134 B.n926 B.n925 71.676
R1135 B.n926 B.n2 71.676
R1136 B.n123 B.t10 69.8713
R1137 B.n484 B.t13 69.8713
R1138 B.n126 B.t7 69.8495
R1139 B.n481 B.t16 69.8495
R1140 B.n233 B.n126 59.5399
R1141 B.n124 B.n123 59.5399
R1142 B.n595 B.n484 59.5399
R1143 B.n482 B.n481 59.5399
R1144 B.n719 B.n417 59.241
R1145 B.n858 B.n58 59.241
R1146 B.n126 B.n125 51.2005
R1147 B.n123 B.n122 51.2005
R1148 B.n484 B.n483 51.2005
R1149 B.n481 B.n480 51.2005
R1150 B.n726 B.n417 34.4309
R1151 B.n726 B.n413 34.4309
R1152 B.n732 B.n413 34.4309
R1153 B.n732 B.n409 34.4309
R1154 B.n738 B.n409 34.4309
R1155 B.n738 B.n405 34.4309
R1156 B.n744 B.n405 34.4309
R1157 B.n750 B.n401 34.4309
R1158 B.n750 B.n397 34.4309
R1159 B.n756 B.n397 34.4309
R1160 B.n756 B.n393 34.4309
R1161 B.n762 B.n393 34.4309
R1162 B.n762 B.n389 34.4309
R1163 B.n768 B.n389 34.4309
R1164 B.n768 B.n384 34.4309
R1165 B.n774 B.n384 34.4309
R1166 B.n774 B.n385 34.4309
R1167 B.n780 B.n377 34.4309
R1168 B.n786 B.n377 34.4309
R1169 B.n786 B.n373 34.4309
R1170 B.n792 B.n373 34.4309
R1171 B.n792 B.n368 34.4309
R1172 B.n798 B.n368 34.4309
R1173 B.n798 B.n369 34.4309
R1174 B.n805 B.n361 34.4309
R1175 B.n811 B.n361 34.4309
R1176 B.n811 B.n4 34.4309
R1177 B.n924 B.n4 34.4309
R1178 B.n924 B.n923 34.4309
R1179 B.n923 B.n922 34.4309
R1180 B.n922 B.n8 34.4309
R1181 B.n12 B.n8 34.4309
R1182 B.n915 B.n12 34.4309
R1183 B.n914 B.n913 34.4309
R1184 B.n913 B.n16 34.4309
R1185 B.n907 B.n16 34.4309
R1186 B.n907 B.n906 34.4309
R1187 B.n906 B.n905 34.4309
R1188 B.n905 B.n23 34.4309
R1189 B.n899 B.n23 34.4309
R1190 B.n898 B.n897 34.4309
R1191 B.n897 B.n30 34.4309
R1192 B.n891 B.n30 34.4309
R1193 B.n891 B.n890 34.4309
R1194 B.n890 B.n889 34.4309
R1195 B.n889 B.n37 34.4309
R1196 B.n883 B.n37 34.4309
R1197 B.n883 B.n882 34.4309
R1198 B.n882 B.n881 34.4309
R1199 B.n881 B.n44 34.4309
R1200 B.n875 B.n874 34.4309
R1201 B.n874 B.n873 34.4309
R1202 B.n873 B.n51 34.4309
R1203 B.n867 B.n51 34.4309
R1204 B.n867 B.n866 34.4309
R1205 B.n866 B.n865 34.4309
R1206 B.n865 B.n58 34.4309
R1207 B.n805 B.t3 33.9245
R1208 B.n915 B.t0 33.9245
R1209 B.n723 B.n722 31.3761
R1210 B.n486 B.n415 31.3761
R1211 B.n856 B.n855 31.3761
R1212 B.n862 B.n861 31.3761
R1213 B.n780 B.t2 25.8233
R1214 B.n899 B.t1 25.8233
R1215 B.t12 B.n401 24.8106
R1216 B.t5 B.n44 24.8106
R1217 B B.n927 18.0485
R1218 B.n724 B.n723 10.6151
R1219 B.n724 B.n411 10.6151
R1220 B.n734 B.n411 10.6151
R1221 B.n735 B.n734 10.6151
R1222 B.n736 B.n735 10.6151
R1223 B.n736 B.n403 10.6151
R1224 B.n746 B.n403 10.6151
R1225 B.n747 B.n746 10.6151
R1226 B.n748 B.n747 10.6151
R1227 B.n748 B.n395 10.6151
R1228 B.n758 B.n395 10.6151
R1229 B.n759 B.n758 10.6151
R1230 B.n760 B.n759 10.6151
R1231 B.n760 B.n387 10.6151
R1232 B.n770 B.n387 10.6151
R1233 B.n771 B.n770 10.6151
R1234 B.n772 B.n771 10.6151
R1235 B.n772 B.n379 10.6151
R1236 B.n782 B.n379 10.6151
R1237 B.n783 B.n782 10.6151
R1238 B.n784 B.n783 10.6151
R1239 B.n784 B.n371 10.6151
R1240 B.n794 B.n371 10.6151
R1241 B.n795 B.n794 10.6151
R1242 B.n796 B.n795 10.6151
R1243 B.n796 B.n363 10.6151
R1244 B.n807 B.n363 10.6151
R1245 B.n808 B.n807 10.6151
R1246 B.n809 B.n808 10.6151
R1247 B.n809 B.n0 10.6151
R1248 B.n722 B.n419 10.6151
R1249 B.n717 B.n419 10.6151
R1250 B.n717 B.n716 10.6151
R1251 B.n716 B.n715 10.6151
R1252 B.n715 B.n712 10.6151
R1253 B.n712 B.n711 10.6151
R1254 B.n711 B.n708 10.6151
R1255 B.n708 B.n707 10.6151
R1256 B.n707 B.n704 10.6151
R1257 B.n704 B.n703 10.6151
R1258 B.n703 B.n700 10.6151
R1259 B.n700 B.n699 10.6151
R1260 B.n699 B.n696 10.6151
R1261 B.n696 B.n695 10.6151
R1262 B.n695 B.n692 10.6151
R1263 B.n692 B.n691 10.6151
R1264 B.n691 B.n688 10.6151
R1265 B.n688 B.n687 10.6151
R1266 B.n687 B.n684 10.6151
R1267 B.n684 B.n683 10.6151
R1268 B.n683 B.n680 10.6151
R1269 B.n680 B.n679 10.6151
R1270 B.n679 B.n676 10.6151
R1271 B.n676 B.n675 10.6151
R1272 B.n675 B.n672 10.6151
R1273 B.n672 B.n671 10.6151
R1274 B.n671 B.n668 10.6151
R1275 B.n668 B.n667 10.6151
R1276 B.n667 B.n664 10.6151
R1277 B.n664 B.n663 10.6151
R1278 B.n663 B.n660 10.6151
R1279 B.n660 B.n659 10.6151
R1280 B.n659 B.n656 10.6151
R1281 B.n656 B.n655 10.6151
R1282 B.n655 B.n652 10.6151
R1283 B.n652 B.n651 10.6151
R1284 B.n651 B.n648 10.6151
R1285 B.n648 B.n647 10.6151
R1286 B.n647 B.n644 10.6151
R1287 B.n644 B.n643 10.6151
R1288 B.n643 B.n640 10.6151
R1289 B.n640 B.n639 10.6151
R1290 B.n639 B.n636 10.6151
R1291 B.n636 B.n635 10.6151
R1292 B.n635 B.n632 10.6151
R1293 B.n632 B.n631 10.6151
R1294 B.n631 B.n628 10.6151
R1295 B.n628 B.n627 10.6151
R1296 B.n627 B.n624 10.6151
R1297 B.n624 B.n623 10.6151
R1298 B.n623 B.n620 10.6151
R1299 B.n620 B.n619 10.6151
R1300 B.n619 B.n616 10.6151
R1301 B.n616 B.n615 10.6151
R1302 B.n612 B.n611 10.6151
R1303 B.n611 B.n608 10.6151
R1304 B.n608 B.n607 10.6151
R1305 B.n607 B.n604 10.6151
R1306 B.n604 B.n603 10.6151
R1307 B.n603 B.n600 10.6151
R1308 B.n600 B.n599 10.6151
R1309 B.n599 B.n596 10.6151
R1310 B.n594 B.n591 10.6151
R1311 B.n591 B.n590 10.6151
R1312 B.n590 B.n587 10.6151
R1313 B.n587 B.n586 10.6151
R1314 B.n586 B.n583 10.6151
R1315 B.n583 B.n582 10.6151
R1316 B.n582 B.n579 10.6151
R1317 B.n579 B.n578 10.6151
R1318 B.n578 B.n575 10.6151
R1319 B.n575 B.n574 10.6151
R1320 B.n574 B.n571 10.6151
R1321 B.n571 B.n570 10.6151
R1322 B.n570 B.n567 10.6151
R1323 B.n567 B.n566 10.6151
R1324 B.n566 B.n563 10.6151
R1325 B.n563 B.n562 10.6151
R1326 B.n562 B.n559 10.6151
R1327 B.n559 B.n558 10.6151
R1328 B.n558 B.n555 10.6151
R1329 B.n555 B.n554 10.6151
R1330 B.n554 B.n551 10.6151
R1331 B.n551 B.n550 10.6151
R1332 B.n550 B.n547 10.6151
R1333 B.n547 B.n546 10.6151
R1334 B.n546 B.n543 10.6151
R1335 B.n543 B.n542 10.6151
R1336 B.n542 B.n539 10.6151
R1337 B.n539 B.n538 10.6151
R1338 B.n538 B.n535 10.6151
R1339 B.n535 B.n534 10.6151
R1340 B.n534 B.n531 10.6151
R1341 B.n531 B.n530 10.6151
R1342 B.n530 B.n527 10.6151
R1343 B.n527 B.n526 10.6151
R1344 B.n526 B.n523 10.6151
R1345 B.n523 B.n522 10.6151
R1346 B.n522 B.n519 10.6151
R1347 B.n519 B.n518 10.6151
R1348 B.n518 B.n515 10.6151
R1349 B.n515 B.n514 10.6151
R1350 B.n514 B.n511 10.6151
R1351 B.n511 B.n510 10.6151
R1352 B.n510 B.n507 10.6151
R1353 B.n507 B.n506 10.6151
R1354 B.n506 B.n503 10.6151
R1355 B.n503 B.n502 10.6151
R1356 B.n502 B.n499 10.6151
R1357 B.n499 B.n498 10.6151
R1358 B.n498 B.n495 10.6151
R1359 B.n495 B.n494 10.6151
R1360 B.n494 B.n491 10.6151
R1361 B.n491 B.n490 10.6151
R1362 B.n490 B.n487 10.6151
R1363 B.n487 B.n486 10.6151
R1364 B.n728 B.n415 10.6151
R1365 B.n729 B.n728 10.6151
R1366 B.n730 B.n729 10.6151
R1367 B.n730 B.n407 10.6151
R1368 B.n740 B.n407 10.6151
R1369 B.n741 B.n740 10.6151
R1370 B.n742 B.n741 10.6151
R1371 B.n742 B.n399 10.6151
R1372 B.n752 B.n399 10.6151
R1373 B.n753 B.n752 10.6151
R1374 B.n754 B.n753 10.6151
R1375 B.n754 B.n391 10.6151
R1376 B.n764 B.n391 10.6151
R1377 B.n765 B.n764 10.6151
R1378 B.n766 B.n765 10.6151
R1379 B.n766 B.n382 10.6151
R1380 B.n776 B.n382 10.6151
R1381 B.n777 B.n776 10.6151
R1382 B.n778 B.n777 10.6151
R1383 B.n778 B.n375 10.6151
R1384 B.n788 B.n375 10.6151
R1385 B.n789 B.n788 10.6151
R1386 B.n790 B.n789 10.6151
R1387 B.n790 B.n366 10.6151
R1388 B.n800 B.n366 10.6151
R1389 B.n801 B.n800 10.6151
R1390 B.n803 B.n801 10.6151
R1391 B.n803 B.n802 10.6151
R1392 B.n802 B.n359 10.6151
R1393 B.n814 B.n359 10.6151
R1394 B.n815 B.n814 10.6151
R1395 B.n816 B.n815 10.6151
R1396 B.n817 B.n816 10.6151
R1397 B.n818 B.n817 10.6151
R1398 B.n821 B.n818 10.6151
R1399 B.n822 B.n821 10.6151
R1400 B.n823 B.n822 10.6151
R1401 B.n824 B.n823 10.6151
R1402 B.n826 B.n824 10.6151
R1403 B.n827 B.n826 10.6151
R1404 B.n828 B.n827 10.6151
R1405 B.n829 B.n828 10.6151
R1406 B.n831 B.n829 10.6151
R1407 B.n832 B.n831 10.6151
R1408 B.n833 B.n832 10.6151
R1409 B.n834 B.n833 10.6151
R1410 B.n836 B.n834 10.6151
R1411 B.n837 B.n836 10.6151
R1412 B.n838 B.n837 10.6151
R1413 B.n839 B.n838 10.6151
R1414 B.n841 B.n839 10.6151
R1415 B.n842 B.n841 10.6151
R1416 B.n843 B.n842 10.6151
R1417 B.n844 B.n843 10.6151
R1418 B.n846 B.n844 10.6151
R1419 B.n847 B.n846 10.6151
R1420 B.n848 B.n847 10.6151
R1421 B.n849 B.n848 10.6151
R1422 B.n851 B.n849 10.6151
R1423 B.n852 B.n851 10.6151
R1424 B.n853 B.n852 10.6151
R1425 B.n854 B.n853 10.6151
R1426 B.n855 B.n854 10.6151
R1427 B.n919 B.n1 10.6151
R1428 B.n919 B.n918 10.6151
R1429 B.n918 B.n917 10.6151
R1430 B.n917 B.n10 10.6151
R1431 B.n911 B.n10 10.6151
R1432 B.n911 B.n910 10.6151
R1433 B.n910 B.n909 10.6151
R1434 B.n909 B.n18 10.6151
R1435 B.n903 B.n18 10.6151
R1436 B.n903 B.n902 10.6151
R1437 B.n902 B.n901 10.6151
R1438 B.n901 B.n25 10.6151
R1439 B.n895 B.n25 10.6151
R1440 B.n895 B.n894 10.6151
R1441 B.n894 B.n893 10.6151
R1442 B.n893 B.n32 10.6151
R1443 B.n887 B.n32 10.6151
R1444 B.n887 B.n886 10.6151
R1445 B.n886 B.n885 10.6151
R1446 B.n885 B.n39 10.6151
R1447 B.n879 B.n39 10.6151
R1448 B.n879 B.n878 10.6151
R1449 B.n878 B.n877 10.6151
R1450 B.n877 B.n46 10.6151
R1451 B.n871 B.n46 10.6151
R1452 B.n871 B.n870 10.6151
R1453 B.n870 B.n869 10.6151
R1454 B.n869 B.n53 10.6151
R1455 B.n863 B.n53 10.6151
R1456 B.n863 B.n862 10.6151
R1457 B.n861 B.n60 10.6151
R1458 B.n128 B.n60 10.6151
R1459 B.n129 B.n128 10.6151
R1460 B.n132 B.n129 10.6151
R1461 B.n133 B.n132 10.6151
R1462 B.n136 B.n133 10.6151
R1463 B.n137 B.n136 10.6151
R1464 B.n140 B.n137 10.6151
R1465 B.n141 B.n140 10.6151
R1466 B.n144 B.n141 10.6151
R1467 B.n145 B.n144 10.6151
R1468 B.n148 B.n145 10.6151
R1469 B.n149 B.n148 10.6151
R1470 B.n152 B.n149 10.6151
R1471 B.n153 B.n152 10.6151
R1472 B.n156 B.n153 10.6151
R1473 B.n157 B.n156 10.6151
R1474 B.n160 B.n157 10.6151
R1475 B.n161 B.n160 10.6151
R1476 B.n164 B.n161 10.6151
R1477 B.n165 B.n164 10.6151
R1478 B.n168 B.n165 10.6151
R1479 B.n169 B.n168 10.6151
R1480 B.n172 B.n169 10.6151
R1481 B.n173 B.n172 10.6151
R1482 B.n176 B.n173 10.6151
R1483 B.n177 B.n176 10.6151
R1484 B.n180 B.n177 10.6151
R1485 B.n181 B.n180 10.6151
R1486 B.n184 B.n181 10.6151
R1487 B.n185 B.n184 10.6151
R1488 B.n188 B.n185 10.6151
R1489 B.n189 B.n188 10.6151
R1490 B.n192 B.n189 10.6151
R1491 B.n193 B.n192 10.6151
R1492 B.n196 B.n193 10.6151
R1493 B.n197 B.n196 10.6151
R1494 B.n200 B.n197 10.6151
R1495 B.n201 B.n200 10.6151
R1496 B.n204 B.n201 10.6151
R1497 B.n205 B.n204 10.6151
R1498 B.n208 B.n205 10.6151
R1499 B.n209 B.n208 10.6151
R1500 B.n212 B.n209 10.6151
R1501 B.n213 B.n212 10.6151
R1502 B.n216 B.n213 10.6151
R1503 B.n217 B.n216 10.6151
R1504 B.n220 B.n217 10.6151
R1505 B.n221 B.n220 10.6151
R1506 B.n224 B.n221 10.6151
R1507 B.n225 B.n224 10.6151
R1508 B.n228 B.n225 10.6151
R1509 B.n229 B.n228 10.6151
R1510 B.n232 B.n229 10.6151
R1511 B.n237 B.n234 10.6151
R1512 B.n238 B.n237 10.6151
R1513 B.n241 B.n238 10.6151
R1514 B.n242 B.n241 10.6151
R1515 B.n245 B.n242 10.6151
R1516 B.n246 B.n245 10.6151
R1517 B.n249 B.n246 10.6151
R1518 B.n250 B.n249 10.6151
R1519 B.n254 B.n253 10.6151
R1520 B.n257 B.n254 10.6151
R1521 B.n258 B.n257 10.6151
R1522 B.n261 B.n258 10.6151
R1523 B.n262 B.n261 10.6151
R1524 B.n265 B.n262 10.6151
R1525 B.n266 B.n265 10.6151
R1526 B.n269 B.n266 10.6151
R1527 B.n270 B.n269 10.6151
R1528 B.n273 B.n270 10.6151
R1529 B.n274 B.n273 10.6151
R1530 B.n277 B.n274 10.6151
R1531 B.n278 B.n277 10.6151
R1532 B.n281 B.n278 10.6151
R1533 B.n282 B.n281 10.6151
R1534 B.n285 B.n282 10.6151
R1535 B.n286 B.n285 10.6151
R1536 B.n289 B.n286 10.6151
R1537 B.n290 B.n289 10.6151
R1538 B.n293 B.n290 10.6151
R1539 B.n294 B.n293 10.6151
R1540 B.n297 B.n294 10.6151
R1541 B.n298 B.n297 10.6151
R1542 B.n301 B.n298 10.6151
R1543 B.n302 B.n301 10.6151
R1544 B.n305 B.n302 10.6151
R1545 B.n306 B.n305 10.6151
R1546 B.n309 B.n306 10.6151
R1547 B.n310 B.n309 10.6151
R1548 B.n313 B.n310 10.6151
R1549 B.n314 B.n313 10.6151
R1550 B.n317 B.n314 10.6151
R1551 B.n318 B.n317 10.6151
R1552 B.n321 B.n318 10.6151
R1553 B.n322 B.n321 10.6151
R1554 B.n325 B.n322 10.6151
R1555 B.n326 B.n325 10.6151
R1556 B.n329 B.n326 10.6151
R1557 B.n330 B.n329 10.6151
R1558 B.n333 B.n330 10.6151
R1559 B.n334 B.n333 10.6151
R1560 B.n337 B.n334 10.6151
R1561 B.n338 B.n337 10.6151
R1562 B.n341 B.n338 10.6151
R1563 B.n342 B.n341 10.6151
R1564 B.n345 B.n342 10.6151
R1565 B.n346 B.n345 10.6151
R1566 B.n349 B.n346 10.6151
R1567 B.n350 B.n349 10.6151
R1568 B.n353 B.n350 10.6151
R1569 B.n354 B.n353 10.6151
R1570 B.n357 B.n354 10.6151
R1571 B.n358 B.n357 10.6151
R1572 B.n856 B.n358 10.6151
R1573 B.n744 B.t12 9.62075
R1574 B.n875 B.t5 9.62075
R1575 B.n385 B.t2 8.60809
R1576 B.t1 B.n898 8.60809
R1577 B.n927 B.n0 8.11757
R1578 B.n927 B.n1 8.11757
R1579 B.n612 B.n482 6.5566
R1580 B.n596 B.n595 6.5566
R1581 B.n234 B.n233 6.5566
R1582 B.n250 B.n124 6.5566
R1583 B.n615 B.n482 4.05904
R1584 B.n595 B.n594 4.05904
R1585 B.n233 B.n232 4.05904
R1586 B.n253 B.n124 4.05904
R1587 B.n369 B.t3 0.506829
R1588 B.t0 B.n914 0.506829
R1589 VP.n3 VP.t0 208.026
R1590 VP.n3 VP.t2 207.371
R1591 VP.n5 VP.t3 171.621
R1592 VP.n13 VP.t1 171.621
R1593 VP.n12 VP.n0 161.3
R1594 VP.n11 VP.n10 161.3
R1595 VP.n9 VP.n1 161.3
R1596 VP.n8 VP.n7 161.3
R1597 VP.n6 VP.n2 161.3
R1598 VP.n5 VP.n4 95.0976
R1599 VP.n14 VP.n13 95.0976
R1600 VP.n4 VP.n3 54.3341
R1601 VP.n7 VP.n1 40.4934
R1602 VP.n11 VP.n1 40.4934
R1603 VP.n7 VP.n6 24.4675
R1604 VP.n12 VP.n11 24.4675
R1605 VP.n6 VP.n5 15.6594
R1606 VP.n13 VP.n12 15.6594
R1607 VP.n4 VP.n2 0.278367
R1608 VP.n14 VP.n0 0.278367
R1609 VP.n8 VP.n2 0.189894
R1610 VP.n9 VP.n8 0.189894
R1611 VP.n10 VP.n9 0.189894
R1612 VP.n10 VP.n0 0.189894
R1613 VP VP.n14 0.153454
R1614 VDD1 VDD1.n1 106.192
R1615 VDD1 VDD1.n0 61.0016
R1616 VDD1.n0 VDD1.t3 1.20415
R1617 VDD1.n0 VDD1.t1 1.20415
R1618 VDD1.n1 VDD1.t0 1.20415
R1619 VDD1.n1 VDD1.t2 1.20415
C0 VP VN 6.80552f
C1 VN VDD1 0.148568f
C2 VN VTAIL 5.92904f
C3 VP VDD1 6.48315f
C4 VP VTAIL 5.94315f
C5 VN VDD2 6.256701f
C6 VP VDD2 0.375682f
C7 VTAIL VDD1 6.48449f
C8 VDD2 VDD1 0.959552f
C9 VTAIL VDD2 6.53675f
C10 VDD2 B 3.940197f
C11 VDD1 B 8.440801f
C12 VTAIL B 12.569495f
C13 VN B 10.54827f
C14 VP B 8.621383f
C15 VDD1.t3 B 0.347809f
C16 VDD1.t1 B 0.347809f
C17 VDD1.n0 B 3.1573f
C18 VDD1.t0 B 0.347809f
C19 VDD1.t2 B 0.347809f
C20 VDD1.n1 B 4.00977f
C21 VP.n0 B 0.03533f
C22 VP.t1 B 2.79589f
C23 VP.n1 B 0.021663f
C24 VP.n2 B 0.03533f
C25 VP.t3 B 2.79589f
C26 VP.t2 B 2.99103f
C27 VP.t0 B 2.99456f
C28 VP.n3 B 3.44104f
C29 VP.n4 B 1.62179f
C30 VP.n5 B 1.06373f
C31 VP.n6 B 0.041067f
C32 VP.n7 B 0.05326f
C33 VP.n8 B 0.026797f
C34 VP.n9 B 0.026797f
C35 VP.n10 B 0.026797f
C36 VP.n11 B 0.05326f
C37 VP.n12 B 0.041067f
C38 VP.n13 B 1.06373f
C39 VP.n14 B 0.03735f
C40 VTAIL.t4 B 2.25546f
C41 VTAIL.n0 B 0.290877f
C42 VTAIL.t3 B 2.25546f
C43 VTAIL.n1 B 0.344343f
C44 VTAIL.t2 B 2.25546f
C45 VTAIL.n2 B 1.34473f
C46 VTAIL.t7 B 2.25546f
C47 VTAIL.n3 B 1.34473f
C48 VTAIL.t5 B 2.25546f
C49 VTAIL.n4 B 0.34434f
C50 VTAIL.t0 B 2.25546f
C51 VTAIL.n5 B 0.34434f
C52 VTAIL.t1 B 2.25546f
C53 VTAIL.n6 B 1.34473f
C54 VTAIL.t6 B 2.25546f
C55 VTAIL.n7 B 1.2855f
C56 VDD2.t0 B 0.345081f
C57 VDD2.t1 B 0.345081f
C58 VDD2.n0 B 3.95045f
C59 VDD2.t2 B 0.345081f
C60 VDD2.t3 B 0.345081f
C61 VDD2.n1 B 3.13213f
C62 VDD2.n2 B 4.13671f
C63 VN.t3 B 2.95756f
C64 VN.t1 B 2.95408f
C65 VN.n0 B 1.93795f
C66 VN.t2 B 2.95756f
C67 VN.t0 B 2.95408f
C68 VN.n1 B 3.41221f
.ends

