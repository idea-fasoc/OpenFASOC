* NGSPICE file created from diff_pair_sample_1138.ext - technology: sky130A

.subckt diff_pair_sample_1138 VTAIL VN VP B VDD2 VDD1
X0 B.t15 B.t13 B.t14 B.t3 sky130_fd_pr__nfet_01v8 ad=3.4827 pd=18.64 as=0 ps=0 w=8.93 l=1.86
X1 B.t12 B.t10 B.t11 B.t7 sky130_fd_pr__nfet_01v8 ad=3.4827 pd=18.64 as=0 ps=0 w=8.93 l=1.86
X2 B.t9 B.t6 B.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=3.4827 pd=18.64 as=0 ps=0 w=8.93 l=1.86
X3 VDD1.t1 VP.t0 VTAIL.t2 B.t0 sky130_fd_pr__nfet_01v8 ad=3.4827 pd=18.64 as=3.4827 ps=18.64 w=8.93 l=1.86
X4 VDD2.t1 VN.t0 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=3.4827 pd=18.64 as=3.4827 ps=18.64 w=8.93 l=1.86
X5 B.t5 B.t2 B.t4 B.t3 sky130_fd_pr__nfet_01v8 ad=3.4827 pd=18.64 as=0 ps=0 w=8.93 l=1.86
X6 VDD1.t0 VP.t1 VTAIL.t3 B.t1 sky130_fd_pr__nfet_01v8 ad=3.4827 pd=18.64 as=3.4827 ps=18.64 w=8.93 l=1.86
X7 VDD2.t0 VN.t1 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=3.4827 pd=18.64 as=3.4827 ps=18.64 w=8.93 l=1.86
R0 B.n557 B.n556 585
R1 B.n558 B.n557 585
R2 B.n232 B.n79 585
R3 B.n231 B.n230 585
R4 B.n229 B.n228 585
R5 B.n227 B.n226 585
R6 B.n225 B.n224 585
R7 B.n223 B.n222 585
R8 B.n221 B.n220 585
R9 B.n219 B.n218 585
R10 B.n217 B.n216 585
R11 B.n215 B.n214 585
R12 B.n213 B.n212 585
R13 B.n211 B.n210 585
R14 B.n209 B.n208 585
R15 B.n207 B.n206 585
R16 B.n205 B.n204 585
R17 B.n203 B.n202 585
R18 B.n201 B.n200 585
R19 B.n199 B.n198 585
R20 B.n197 B.n196 585
R21 B.n195 B.n194 585
R22 B.n193 B.n192 585
R23 B.n191 B.n190 585
R24 B.n189 B.n188 585
R25 B.n187 B.n186 585
R26 B.n185 B.n184 585
R27 B.n183 B.n182 585
R28 B.n181 B.n180 585
R29 B.n179 B.n178 585
R30 B.n177 B.n176 585
R31 B.n175 B.n174 585
R32 B.n173 B.n172 585
R33 B.n171 B.n170 585
R34 B.n169 B.n168 585
R35 B.n167 B.n166 585
R36 B.n165 B.n164 585
R37 B.n163 B.n162 585
R38 B.n161 B.n160 585
R39 B.n159 B.n158 585
R40 B.n157 B.n156 585
R41 B.n155 B.n154 585
R42 B.n153 B.n152 585
R43 B.n150 B.n149 585
R44 B.n148 B.n147 585
R45 B.n146 B.n145 585
R46 B.n144 B.n143 585
R47 B.n142 B.n141 585
R48 B.n140 B.n139 585
R49 B.n138 B.n137 585
R50 B.n136 B.n135 585
R51 B.n134 B.n133 585
R52 B.n132 B.n131 585
R53 B.n130 B.n129 585
R54 B.n128 B.n127 585
R55 B.n126 B.n125 585
R56 B.n124 B.n123 585
R57 B.n122 B.n121 585
R58 B.n120 B.n119 585
R59 B.n118 B.n117 585
R60 B.n116 B.n115 585
R61 B.n114 B.n113 585
R62 B.n112 B.n111 585
R63 B.n110 B.n109 585
R64 B.n108 B.n107 585
R65 B.n106 B.n105 585
R66 B.n104 B.n103 585
R67 B.n102 B.n101 585
R68 B.n100 B.n99 585
R69 B.n98 B.n97 585
R70 B.n96 B.n95 585
R71 B.n94 B.n93 585
R72 B.n92 B.n91 585
R73 B.n90 B.n89 585
R74 B.n88 B.n87 585
R75 B.n86 B.n85 585
R76 B.n555 B.n41 585
R77 B.n559 B.n41 585
R78 B.n554 B.n40 585
R79 B.n560 B.n40 585
R80 B.n553 B.n552 585
R81 B.n552 B.n36 585
R82 B.n551 B.n35 585
R83 B.n566 B.n35 585
R84 B.n550 B.n34 585
R85 B.n567 B.n34 585
R86 B.n549 B.n33 585
R87 B.n568 B.n33 585
R88 B.n548 B.n547 585
R89 B.n547 B.n32 585
R90 B.n546 B.n28 585
R91 B.n574 B.n28 585
R92 B.n545 B.n27 585
R93 B.n575 B.n27 585
R94 B.n544 B.n26 585
R95 B.n576 B.n26 585
R96 B.n543 B.n542 585
R97 B.n542 B.n22 585
R98 B.n541 B.n21 585
R99 B.n582 B.n21 585
R100 B.n540 B.n20 585
R101 B.n583 B.n20 585
R102 B.n539 B.n19 585
R103 B.n584 B.n19 585
R104 B.n538 B.n537 585
R105 B.n537 B.n15 585
R106 B.n536 B.n14 585
R107 B.n590 B.n14 585
R108 B.n535 B.n13 585
R109 B.n591 B.n13 585
R110 B.n534 B.n12 585
R111 B.n592 B.n12 585
R112 B.n533 B.n532 585
R113 B.n532 B.n8 585
R114 B.n531 B.n7 585
R115 B.n598 B.n7 585
R116 B.n530 B.n6 585
R117 B.n599 B.n6 585
R118 B.n529 B.n5 585
R119 B.n600 B.n5 585
R120 B.n528 B.n527 585
R121 B.n527 B.n4 585
R122 B.n526 B.n233 585
R123 B.n526 B.n525 585
R124 B.n516 B.n234 585
R125 B.n235 B.n234 585
R126 B.n518 B.n517 585
R127 B.n519 B.n518 585
R128 B.n515 B.n239 585
R129 B.n243 B.n239 585
R130 B.n514 B.n513 585
R131 B.n513 B.n512 585
R132 B.n241 B.n240 585
R133 B.n242 B.n241 585
R134 B.n505 B.n504 585
R135 B.n506 B.n505 585
R136 B.n503 B.n248 585
R137 B.n248 B.n247 585
R138 B.n502 B.n501 585
R139 B.n501 B.n500 585
R140 B.n250 B.n249 585
R141 B.n251 B.n250 585
R142 B.n493 B.n492 585
R143 B.n494 B.n493 585
R144 B.n491 B.n256 585
R145 B.n256 B.n255 585
R146 B.n490 B.n489 585
R147 B.n489 B.n488 585
R148 B.n258 B.n257 585
R149 B.n481 B.n258 585
R150 B.n480 B.n479 585
R151 B.n482 B.n480 585
R152 B.n478 B.n263 585
R153 B.n263 B.n262 585
R154 B.n477 B.n476 585
R155 B.n476 B.n475 585
R156 B.n265 B.n264 585
R157 B.n266 B.n265 585
R158 B.n468 B.n467 585
R159 B.n469 B.n468 585
R160 B.n466 B.n271 585
R161 B.n271 B.n270 585
R162 B.n460 B.n459 585
R163 B.n458 B.n310 585
R164 B.n457 B.n309 585
R165 B.n462 B.n309 585
R166 B.n456 B.n455 585
R167 B.n454 B.n453 585
R168 B.n452 B.n451 585
R169 B.n450 B.n449 585
R170 B.n448 B.n447 585
R171 B.n446 B.n445 585
R172 B.n444 B.n443 585
R173 B.n442 B.n441 585
R174 B.n440 B.n439 585
R175 B.n438 B.n437 585
R176 B.n436 B.n435 585
R177 B.n434 B.n433 585
R178 B.n432 B.n431 585
R179 B.n430 B.n429 585
R180 B.n428 B.n427 585
R181 B.n426 B.n425 585
R182 B.n424 B.n423 585
R183 B.n422 B.n421 585
R184 B.n420 B.n419 585
R185 B.n418 B.n417 585
R186 B.n416 B.n415 585
R187 B.n414 B.n413 585
R188 B.n412 B.n411 585
R189 B.n410 B.n409 585
R190 B.n408 B.n407 585
R191 B.n406 B.n405 585
R192 B.n404 B.n403 585
R193 B.n402 B.n401 585
R194 B.n400 B.n399 585
R195 B.n398 B.n397 585
R196 B.n396 B.n395 585
R197 B.n394 B.n393 585
R198 B.n392 B.n391 585
R199 B.n390 B.n389 585
R200 B.n388 B.n387 585
R201 B.n386 B.n385 585
R202 B.n384 B.n383 585
R203 B.n382 B.n381 585
R204 B.n380 B.n379 585
R205 B.n377 B.n376 585
R206 B.n375 B.n374 585
R207 B.n373 B.n372 585
R208 B.n371 B.n370 585
R209 B.n369 B.n368 585
R210 B.n367 B.n366 585
R211 B.n365 B.n364 585
R212 B.n363 B.n362 585
R213 B.n361 B.n360 585
R214 B.n359 B.n358 585
R215 B.n357 B.n356 585
R216 B.n355 B.n354 585
R217 B.n353 B.n352 585
R218 B.n351 B.n350 585
R219 B.n349 B.n348 585
R220 B.n347 B.n346 585
R221 B.n345 B.n344 585
R222 B.n343 B.n342 585
R223 B.n341 B.n340 585
R224 B.n339 B.n338 585
R225 B.n337 B.n336 585
R226 B.n335 B.n334 585
R227 B.n333 B.n332 585
R228 B.n331 B.n330 585
R229 B.n329 B.n328 585
R230 B.n327 B.n326 585
R231 B.n325 B.n324 585
R232 B.n323 B.n322 585
R233 B.n321 B.n320 585
R234 B.n319 B.n318 585
R235 B.n317 B.n316 585
R236 B.n273 B.n272 585
R237 B.n465 B.n464 585
R238 B.n269 B.n268 585
R239 B.n270 B.n269 585
R240 B.n471 B.n470 585
R241 B.n470 B.n469 585
R242 B.n472 B.n267 585
R243 B.n267 B.n266 585
R244 B.n474 B.n473 585
R245 B.n475 B.n474 585
R246 B.n261 B.n260 585
R247 B.n262 B.n261 585
R248 B.n484 B.n483 585
R249 B.n483 B.n482 585
R250 B.n485 B.n259 585
R251 B.n481 B.n259 585
R252 B.n487 B.n486 585
R253 B.n488 B.n487 585
R254 B.n254 B.n253 585
R255 B.n255 B.n254 585
R256 B.n496 B.n495 585
R257 B.n495 B.n494 585
R258 B.n497 B.n252 585
R259 B.n252 B.n251 585
R260 B.n499 B.n498 585
R261 B.n500 B.n499 585
R262 B.n246 B.n245 585
R263 B.n247 B.n246 585
R264 B.n508 B.n507 585
R265 B.n507 B.n506 585
R266 B.n509 B.n244 585
R267 B.n244 B.n242 585
R268 B.n511 B.n510 585
R269 B.n512 B.n511 585
R270 B.n238 B.n237 585
R271 B.n243 B.n238 585
R272 B.n521 B.n520 585
R273 B.n520 B.n519 585
R274 B.n522 B.n236 585
R275 B.n236 B.n235 585
R276 B.n524 B.n523 585
R277 B.n525 B.n524 585
R278 B.n2 B.n0 585
R279 B.n4 B.n2 585
R280 B.n3 B.n1 585
R281 B.n599 B.n3 585
R282 B.n597 B.n596 585
R283 B.n598 B.n597 585
R284 B.n595 B.n9 585
R285 B.n9 B.n8 585
R286 B.n594 B.n593 585
R287 B.n593 B.n592 585
R288 B.n11 B.n10 585
R289 B.n591 B.n11 585
R290 B.n589 B.n588 585
R291 B.n590 B.n589 585
R292 B.n587 B.n16 585
R293 B.n16 B.n15 585
R294 B.n586 B.n585 585
R295 B.n585 B.n584 585
R296 B.n18 B.n17 585
R297 B.n583 B.n18 585
R298 B.n581 B.n580 585
R299 B.n582 B.n581 585
R300 B.n579 B.n23 585
R301 B.n23 B.n22 585
R302 B.n578 B.n577 585
R303 B.n577 B.n576 585
R304 B.n25 B.n24 585
R305 B.n575 B.n25 585
R306 B.n573 B.n572 585
R307 B.n574 B.n573 585
R308 B.n571 B.n29 585
R309 B.n32 B.n29 585
R310 B.n570 B.n569 585
R311 B.n569 B.n568 585
R312 B.n31 B.n30 585
R313 B.n567 B.n31 585
R314 B.n565 B.n564 585
R315 B.n566 B.n565 585
R316 B.n563 B.n37 585
R317 B.n37 B.n36 585
R318 B.n562 B.n561 585
R319 B.n561 B.n560 585
R320 B.n39 B.n38 585
R321 B.n559 B.n39 585
R322 B.n602 B.n601 585
R323 B.n601 B.n600 585
R324 B.n460 B.n269 478.086
R325 B.n85 B.n39 478.086
R326 B.n464 B.n271 478.086
R327 B.n557 B.n41 478.086
R328 B.n314 B.t13 322.276
R329 B.n311 B.t2 322.276
R330 B.n83 B.t6 322.276
R331 B.n80 B.t10 322.276
R332 B.n558 B.n78 256.663
R333 B.n558 B.n77 256.663
R334 B.n558 B.n76 256.663
R335 B.n558 B.n75 256.663
R336 B.n558 B.n74 256.663
R337 B.n558 B.n73 256.663
R338 B.n558 B.n72 256.663
R339 B.n558 B.n71 256.663
R340 B.n558 B.n70 256.663
R341 B.n558 B.n69 256.663
R342 B.n558 B.n68 256.663
R343 B.n558 B.n67 256.663
R344 B.n558 B.n66 256.663
R345 B.n558 B.n65 256.663
R346 B.n558 B.n64 256.663
R347 B.n558 B.n63 256.663
R348 B.n558 B.n62 256.663
R349 B.n558 B.n61 256.663
R350 B.n558 B.n60 256.663
R351 B.n558 B.n59 256.663
R352 B.n558 B.n58 256.663
R353 B.n558 B.n57 256.663
R354 B.n558 B.n56 256.663
R355 B.n558 B.n55 256.663
R356 B.n558 B.n54 256.663
R357 B.n558 B.n53 256.663
R358 B.n558 B.n52 256.663
R359 B.n558 B.n51 256.663
R360 B.n558 B.n50 256.663
R361 B.n558 B.n49 256.663
R362 B.n558 B.n48 256.663
R363 B.n558 B.n47 256.663
R364 B.n558 B.n46 256.663
R365 B.n558 B.n45 256.663
R366 B.n558 B.n44 256.663
R367 B.n558 B.n43 256.663
R368 B.n558 B.n42 256.663
R369 B.n462 B.n461 256.663
R370 B.n462 B.n274 256.663
R371 B.n462 B.n275 256.663
R372 B.n462 B.n276 256.663
R373 B.n462 B.n277 256.663
R374 B.n462 B.n278 256.663
R375 B.n462 B.n279 256.663
R376 B.n462 B.n280 256.663
R377 B.n462 B.n281 256.663
R378 B.n462 B.n282 256.663
R379 B.n462 B.n283 256.663
R380 B.n462 B.n284 256.663
R381 B.n462 B.n285 256.663
R382 B.n462 B.n286 256.663
R383 B.n462 B.n287 256.663
R384 B.n462 B.n288 256.663
R385 B.n462 B.n289 256.663
R386 B.n462 B.n290 256.663
R387 B.n462 B.n291 256.663
R388 B.n462 B.n292 256.663
R389 B.n462 B.n293 256.663
R390 B.n462 B.n294 256.663
R391 B.n462 B.n295 256.663
R392 B.n462 B.n296 256.663
R393 B.n462 B.n297 256.663
R394 B.n462 B.n298 256.663
R395 B.n462 B.n299 256.663
R396 B.n462 B.n300 256.663
R397 B.n462 B.n301 256.663
R398 B.n462 B.n302 256.663
R399 B.n462 B.n303 256.663
R400 B.n462 B.n304 256.663
R401 B.n462 B.n305 256.663
R402 B.n462 B.n306 256.663
R403 B.n462 B.n307 256.663
R404 B.n462 B.n308 256.663
R405 B.n463 B.n462 256.663
R406 B.n470 B.n269 163.367
R407 B.n470 B.n267 163.367
R408 B.n474 B.n267 163.367
R409 B.n474 B.n261 163.367
R410 B.n483 B.n261 163.367
R411 B.n483 B.n259 163.367
R412 B.n487 B.n259 163.367
R413 B.n487 B.n254 163.367
R414 B.n495 B.n254 163.367
R415 B.n495 B.n252 163.367
R416 B.n499 B.n252 163.367
R417 B.n499 B.n246 163.367
R418 B.n507 B.n246 163.367
R419 B.n507 B.n244 163.367
R420 B.n511 B.n244 163.367
R421 B.n511 B.n238 163.367
R422 B.n520 B.n238 163.367
R423 B.n520 B.n236 163.367
R424 B.n524 B.n236 163.367
R425 B.n524 B.n2 163.367
R426 B.n601 B.n2 163.367
R427 B.n601 B.n3 163.367
R428 B.n597 B.n3 163.367
R429 B.n597 B.n9 163.367
R430 B.n593 B.n9 163.367
R431 B.n593 B.n11 163.367
R432 B.n589 B.n11 163.367
R433 B.n589 B.n16 163.367
R434 B.n585 B.n16 163.367
R435 B.n585 B.n18 163.367
R436 B.n581 B.n18 163.367
R437 B.n581 B.n23 163.367
R438 B.n577 B.n23 163.367
R439 B.n577 B.n25 163.367
R440 B.n573 B.n25 163.367
R441 B.n573 B.n29 163.367
R442 B.n569 B.n29 163.367
R443 B.n569 B.n31 163.367
R444 B.n565 B.n31 163.367
R445 B.n565 B.n37 163.367
R446 B.n561 B.n37 163.367
R447 B.n561 B.n39 163.367
R448 B.n310 B.n309 163.367
R449 B.n455 B.n309 163.367
R450 B.n453 B.n452 163.367
R451 B.n449 B.n448 163.367
R452 B.n445 B.n444 163.367
R453 B.n441 B.n440 163.367
R454 B.n437 B.n436 163.367
R455 B.n433 B.n432 163.367
R456 B.n429 B.n428 163.367
R457 B.n425 B.n424 163.367
R458 B.n421 B.n420 163.367
R459 B.n417 B.n416 163.367
R460 B.n413 B.n412 163.367
R461 B.n409 B.n408 163.367
R462 B.n405 B.n404 163.367
R463 B.n401 B.n400 163.367
R464 B.n397 B.n396 163.367
R465 B.n393 B.n392 163.367
R466 B.n389 B.n388 163.367
R467 B.n385 B.n384 163.367
R468 B.n381 B.n380 163.367
R469 B.n376 B.n375 163.367
R470 B.n372 B.n371 163.367
R471 B.n368 B.n367 163.367
R472 B.n364 B.n363 163.367
R473 B.n360 B.n359 163.367
R474 B.n356 B.n355 163.367
R475 B.n352 B.n351 163.367
R476 B.n348 B.n347 163.367
R477 B.n344 B.n343 163.367
R478 B.n340 B.n339 163.367
R479 B.n336 B.n335 163.367
R480 B.n332 B.n331 163.367
R481 B.n328 B.n327 163.367
R482 B.n324 B.n323 163.367
R483 B.n320 B.n319 163.367
R484 B.n316 B.n273 163.367
R485 B.n468 B.n271 163.367
R486 B.n468 B.n265 163.367
R487 B.n476 B.n265 163.367
R488 B.n476 B.n263 163.367
R489 B.n480 B.n263 163.367
R490 B.n480 B.n258 163.367
R491 B.n489 B.n258 163.367
R492 B.n489 B.n256 163.367
R493 B.n493 B.n256 163.367
R494 B.n493 B.n250 163.367
R495 B.n501 B.n250 163.367
R496 B.n501 B.n248 163.367
R497 B.n505 B.n248 163.367
R498 B.n505 B.n241 163.367
R499 B.n513 B.n241 163.367
R500 B.n513 B.n239 163.367
R501 B.n518 B.n239 163.367
R502 B.n518 B.n234 163.367
R503 B.n526 B.n234 163.367
R504 B.n527 B.n526 163.367
R505 B.n527 B.n5 163.367
R506 B.n6 B.n5 163.367
R507 B.n7 B.n6 163.367
R508 B.n532 B.n7 163.367
R509 B.n532 B.n12 163.367
R510 B.n13 B.n12 163.367
R511 B.n14 B.n13 163.367
R512 B.n537 B.n14 163.367
R513 B.n537 B.n19 163.367
R514 B.n20 B.n19 163.367
R515 B.n21 B.n20 163.367
R516 B.n542 B.n21 163.367
R517 B.n542 B.n26 163.367
R518 B.n27 B.n26 163.367
R519 B.n28 B.n27 163.367
R520 B.n547 B.n28 163.367
R521 B.n547 B.n33 163.367
R522 B.n34 B.n33 163.367
R523 B.n35 B.n34 163.367
R524 B.n552 B.n35 163.367
R525 B.n552 B.n40 163.367
R526 B.n41 B.n40 163.367
R527 B.n89 B.n88 163.367
R528 B.n93 B.n92 163.367
R529 B.n97 B.n96 163.367
R530 B.n101 B.n100 163.367
R531 B.n105 B.n104 163.367
R532 B.n109 B.n108 163.367
R533 B.n113 B.n112 163.367
R534 B.n117 B.n116 163.367
R535 B.n121 B.n120 163.367
R536 B.n125 B.n124 163.367
R537 B.n129 B.n128 163.367
R538 B.n133 B.n132 163.367
R539 B.n137 B.n136 163.367
R540 B.n141 B.n140 163.367
R541 B.n145 B.n144 163.367
R542 B.n149 B.n148 163.367
R543 B.n154 B.n153 163.367
R544 B.n158 B.n157 163.367
R545 B.n162 B.n161 163.367
R546 B.n166 B.n165 163.367
R547 B.n170 B.n169 163.367
R548 B.n174 B.n173 163.367
R549 B.n178 B.n177 163.367
R550 B.n182 B.n181 163.367
R551 B.n186 B.n185 163.367
R552 B.n190 B.n189 163.367
R553 B.n194 B.n193 163.367
R554 B.n198 B.n197 163.367
R555 B.n202 B.n201 163.367
R556 B.n206 B.n205 163.367
R557 B.n210 B.n209 163.367
R558 B.n214 B.n213 163.367
R559 B.n218 B.n217 163.367
R560 B.n222 B.n221 163.367
R561 B.n226 B.n225 163.367
R562 B.n230 B.n229 163.367
R563 B.n557 B.n79 163.367
R564 B.n314 B.t15 112.572
R565 B.n80 B.t11 112.572
R566 B.n311 B.t5 112.561
R567 B.n83 B.t8 112.561
R568 B.n462 B.n270 95.2486
R569 B.n559 B.n558 95.2486
R570 B.n461 B.n460 71.676
R571 B.n455 B.n274 71.676
R572 B.n452 B.n275 71.676
R573 B.n448 B.n276 71.676
R574 B.n444 B.n277 71.676
R575 B.n440 B.n278 71.676
R576 B.n436 B.n279 71.676
R577 B.n432 B.n280 71.676
R578 B.n428 B.n281 71.676
R579 B.n424 B.n282 71.676
R580 B.n420 B.n283 71.676
R581 B.n416 B.n284 71.676
R582 B.n412 B.n285 71.676
R583 B.n408 B.n286 71.676
R584 B.n404 B.n287 71.676
R585 B.n400 B.n288 71.676
R586 B.n396 B.n289 71.676
R587 B.n392 B.n290 71.676
R588 B.n388 B.n291 71.676
R589 B.n384 B.n292 71.676
R590 B.n380 B.n293 71.676
R591 B.n375 B.n294 71.676
R592 B.n371 B.n295 71.676
R593 B.n367 B.n296 71.676
R594 B.n363 B.n297 71.676
R595 B.n359 B.n298 71.676
R596 B.n355 B.n299 71.676
R597 B.n351 B.n300 71.676
R598 B.n347 B.n301 71.676
R599 B.n343 B.n302 71.676
R600 B.n339 B.n303 71.676
R601 B.n335 B.n304 71.676
R602 B.n331 B.n305 71.676
R603 B.n327 B.n306 71.676
R604 B.n323 B.n307 71.676
R605 B.n319 B.n308 71.676
R606 B.n463 B.n273 71.676
R607 B.n85 B.n42 71.676
R608 B.n89 B.n43 71.676
R609 B.n93 B.n44 71.676
R610 B.n97 B.n45 71.676
R611 B.n101 B.n46 71.676
R612 B.n105 B.n47 71.676
R613 B.n109 B.n48 71.676
R614 B.n113 B.n49 71.676
R615 B.n117 B.n50 71.676
R616 B.n121 B.n51 71.676
R617 B.n125 B.n52 71.676
R618 B.n129 B.n53 71.676
R619 B.n133 B.n54 71.676
R620 B.n137 B.n55 71.676
R621 B.n141 B.n56 71.676
R622 B.n145 B.n57 71.676
R623 B.n149 B.n58 71.676
R624 B.n154 B.n59 71.676
R625 B.n158 B.n60 71.676
R626 B.n162 B.n61 71.676
R627 B.n166 B.n62 71.676
R628 B.n170 B.n63 71.676
R629 B.n174 B.n64 71.676
R630 B.n178 B.n65 71.676
R631 B.n182 B.n66 71.676
R632 B.n186 B.n67 71.676
R633 B.n190 B.n68 71.676
R634 B.n194 B.n69 71.676
R635 B.n198 B.n70 71.676
R636 B.n202 B.n71 71.676
R637 B.n206 B.n72 71.676
R638 B.n210 B.n73 71.676
R639 B.n214 B.n74 71.676
R640 B.n218 B.n75 71.676
R641 B.n222 B.n76 71.676
R642 B.n226 B.n77 71.676
R643 B.n230 B.n78 71.676
R644 B.n79 B.n78 71.676
R645 B.n229 B.n77 71.676
R646 B.n225 B.n76 71.676
R647 B.n221 B.n75 71.676
R648 B.n217 B.n74 71.676
R649 B.n213 B.n73 71.676
R650 B.n209 B.n72 71.676
R651 B.n205 B.n71 71.676
R652 B.n201 B.n70 71.676
R653 B.n197 B.n69 71.676
R654 B.n193 B.n68 71.676
R655 B.n189 B.n67 71.676
R656 B.n185 B.n66 71.676
R657 B.n181 B.n65 71.676
R658 B.n177 B.n64 71.676
R659 B.n173 B.n63 71.676
R660 B.n169 B.n62 71.676
R661 B.n165 B.n61 71.676
R662 B.n161 B.n60 71.676
R663 B.n157 B.n59 71.676
R664 B.n153 B.n58 71.676
R665 B.n148 B.n57 71.676
R666 B.n144 B.n56 71.676
R667 B.n140 B.n55 71.676
R668 B.n136 B.n54 71.676
R669 B.n132 B.n53 71.676
R670 B.n128 B.n52 71.676
R671 B.n124 B.n51 71.676
R672 B.n120 B.n50 71.676
R673 B.n116 B.n49 71.676
R674 B.n112 B.n48 71.676
R675 B.n108 B.n47 71.676
R676 B.n104 B.n46 71.676
R677 B.n100 B.n45 71.676
R678 B.n96 B.n44 71.676
R679 B.n92 B.n43 71.676
R680 B.n88 B.n42 71.676
R681 B.n461 B.n310 71.676
R682 B.n453 B.n274 71.676
R683 B.n449 B.n275 71.676
R684 B.n445 B.n276 71.676
R685 B.n441 B.n277 71.676
R686 B.n437 B.n278 71.676
R687 B.n433 B.n279 71.676
R688 B.n429 B.n280 71.676
R689 B.n425 B.n281 71.676
R690 B.n421 B.n282 71.676
R691 B.n417 B.n283 71.676
R692 B.n413 B.n284 71.676
R693 B.n409 B.n285 71.676
R694 B.n405 B.n286 71.676
R695 B.n401 B.n287 71.676
R696 B.n397 B.n288 71.676
R697 B.n393 B.n289 71.676
R698 B.n389 B.n290 71.676
R699 B.n385 B.n291 71.676
R700 B.n381 B.n292 71.676
R701 B.n376 B.n293 71.676
R702 B.n372 B.n294 71.676
R703 B.n368 B.n295 71.676
R704 B.n364 B.n296 71.676
R705 B.n360 B.n297 71.676
R706 B.n356 B.n298 71.676
R707 B.n352 B.n299 71.676
R708 B.n348 B.n300 71.676
R709 B.n344 B.n301 71.676
R710 B.n340 B.n302 71.676
R711 B.n336 B.n303 71.676
R712 B.n332 B.n304 71.676
R713 B.n328 B.n305 71.676
R714 B.n324 B.n306 71.676
R715 B.n320 B.n307 71.676
R716 B.n316 B.n308 71.676
R717 B.n464 B.n463 71.676
R718 B.n315 B.t14 70.0983
R719 B.n81 B.t12 70.0983
R720 B.n312 B.t4 70.0875
R721 B.n84 B.t9 70.0875
R722 B.n378 B.n315 59.5399
R723 B.n313 B.n312 59.5399
R724 B.n151 B.n84 59.5399
R725 B.n82 B.n81 59.5399
R726 B.n469 B.n270 52.658
R727 B.n469 B.n266 52.658
R728 B.n475 B.n266 52.658
R729 B.n475 B.n262 52.658
R730 B.n482 B.n262 52.658
R731 B.n482 B.n481 52.658
R732 B.n488 B.n255 52.658
R733 B.n494 B.n255 52.658
R734 B.n494 B.n251 52.658
R735 B.n500 B.n251 52.658
R736 B.n500 B.n247 52.658
R737 B.n506 B.n247 52.658
R738 B.n506 B.n242 52.658
R739 B.n512 B.n242 52.658
R740 B.n512 B.n243 52.658
R741 B.n519 B.n235 52.658
R742 B.n525 B.n235 52.658
R743 B.n525 B.n4 52.658
R744 B.n600 B.n4 52.658
R745 B.n600 B.n599 52.658
R746 B.n599 B.n598 52.658
R747 B.n598 B.n8 52.658
R748 B.n592 B.n8 52.658
R749 B.n591 B.n590 52.658
R750 B.n590 B.n15 52.658
R751 B.n584 B.n15 52.658
R752 B.n584 B.n583 52.658
R753 B.n583 B.n582 52.658
R754 B.n582 B.n22 52.658
R755 B.n576 B.n22 52.658
R756 B.n576 B.n575 52.658
R757 B.n575 B.n574 52.658
R758 B.n568 B.n32 52.658
R759 B.n568 B.n567 52.658
R760 B.n567 B.n566 52.658
R761 B.n566 B.n36 52.658
R762 B.n560 B.n36 52.658
R763 B.n560 B.n559 52.658
R764 B.n519 B.t1 43.3655
R765 B.n592 B.t0 43.3655
R766 B.n315 B.n314 42.4732
R767 B.n312 B.n311 42.4732
R768 B.n84 B.n83 42.4732
R769 B.n81 B.n80 42.4732
R770 B.n86 B.n38 31.0639
R771 B.n556 B.n555 31.0639
R772 B.n466 B.n465 31.0639
R773 B.n459 B.n268 31.0639
R774 B.n481 B.t3 27.878
R775 B.n32 B.t7 27.878
R776 B.n488 B.t3 24.7805
R777 B.n574 B.t7 24.7805
R778 B B.n602 18.0485
R779 B.n87 B.n86 10.6151
R780 B.n90 B.n87 10.6151
R781 B.n91 B.n90 10.6151
R782 B.n94 B.n91 10.6151
R783 B.n95 B.n94 10.6151
R784 B.n98 B.n95 10.6151
R785 B.n99 B.n98 10.6151
R786 B.n102 B.n99 10.6151
R787 B.n103 B.n102 10.6151
R788 B.n106 B.n103 10.6151
R789 B.n107 B.n106 10.6151
R790 B.n110 B.n107 10.6151
R791 B.n111 B.n110 10.6151
R792 B.n114 B.n111 10.6151
R793 B.n115 B.n114 10.6151
R794 B.n118 B.n115 10.6151
R795 B.n119 B.n118 10.6151
R796 B.n122 B.n119 10.6151
R797 B.n123 B.n122 10.6151
R798 B.n126 B.n123 10.6151
R799 B.n127 B.n126 10.6151
R800 B.n130 B.n127 10.6151
R801 B.n131 B.n130 10.6151
R802 B.n134 B.n131 10.6151
R803 B.n135 B.n134 10.6151
R804 B.n138 B.n135 10.6151
R805 B.n139 B.n138 10.6151
R806 B.n142 B.n139 10.6151
R807 B.n143 B.n142 10.6151
R808 B.n146 B.n143 10.6151
R809 B.n147 B.n146 10.6151
R810 B.n150 B.n147 10.6151
R811 B.n155 B.n152 10.6151
R812 B.n156 B.n155 10.6151
R813 B.n159 B.n156 10.6151
R814 B.n160 B.n159 10.6151
R815 B.n163 B.n160 10.6151
R816 B.n164 B.n163 10.6151
R817 B.n167 B.n164 10.6151
R818 B.n168 B.n167 10.6151
R819 B.n172 B.n171 10.6151
R820 B.n175 B.n172 10.6151
R821 B.n176 B.n175 10.6151
R822 B.n179 B.n176 10.6151
R823 B.n180 B.n179 10.6151
R824 B.n183 B.n180 10.6151
R825 B.n184 B.n183 10.6151
R826 B.n187 B.n184 10.6151
R827 B.n188 B.n187 10.6151
R828 B.n191 B.n188 10.6151
R829 B.n192 B.n191 10.6151
R830 B.n195 B.n192 10.6151
R831 B.n196 B.n195 10.6151
R832 B.n199 B.n196 10.6151
R833 B.n200 B.n199 10.6151
R834 B.n203 B.n200 10.6151
R835 B.n204 B.n203 10.6151
R836 B.n207 B.n204 10.6151
R837 B.n208 B.n207 10.6151
R838 B.n211 B.n208 10.6151
R839 B.n212 B.n211 10.6151
R840 B.n215 B.n212 10.6151
R841 B.n216 B.n215 10.6151
R842 B.n219 B.n216 10.6151
R843 B.n220 B.n219 10.6151
R844 B.n223 B.n220 10.6151
R845 B.n224 B.n223 10.6151
R846 B.n227 B.n224 10.6151
R847 B.n228 B.n227 10.6151
R848 B.n231 B.n228 10.6151
R849 B.n232 B.n231 10.6151
R850 B.n556 B.n232 10.6151
R851 B.n467 B.n466 10.6151
R852 B.n467 B.n264 10.6151
R853 B.n477 B.n264 10.6151
R854 B.n478 B.n477 10.6151
R855 B.n479 B.n478 10.6151
R856 B.n479 B.n257 10.6151
R857 B.n490 B.n257 10.6151
R858 B.n491 B.n490 10.6151
R859 B.n492 B.n491 10.6151
R860 B.n492 B.n249 10.6151
R861 B.n502 B.n249 10.6151
R862 B.n503 B.n502 10.6151
R863 B.n504 B.n503 10.6151
R864 B.n504 B.n240 10.6151
R865 B.n514 B.n240 10.6151
R866 B.n515 B.n514 10.6151
R867 B.n517 B.n515 10.6151
R868 B.n517 B.n516 10.6151
R869 B.n516 B.n233 10.6151
R870 B.n528 B.n233 10.6151
R871 B.n529 B.n528 10.6151
R872 B.n530 B.n529 10.6151
R873 B.n531 B.n530 10.6151
R874 B.n533 B.n531 10.6151
R875 B.n534 B.n533 10.6151
R876 B.n535 B.n534 10.6151
R877 B.n536 B.n535 10.6151
R878 B.n538 B.n536 10.6151
R879 B.n539 B.n538 10.6151
R880 B.n540 B.n539 10.6151
R881 B.n541 B.n540 10.6151
R882 B.n543 B.n541 10.6151
R883 B.n544 B.n543 10.6151
R884 B.n545 B.n544 10.6151
R885 B.n546 B.n545 10.6151
R886 B.n548 B.n546 10.6151
R887 B.n549 B.n548 10.6151
R888 B.n550 B.n549 10.6151
R889 B.n551 B.n550 10.6151
R890 B.n553 B.n551 10.6151
R891 B.n554 B.n553 10.6151
R892 B.n555 B.n554 10.6151
R893 B.n459 B.n458 10.6151
R894 B.n458 B.n457 10.6151
R895 B.n457 B.n456 10.6151
R896 B.n456 B.n454 10.6151
R897 B.n454 B.n451 10.6151
R898 B.n451 B.n450 10.6151
R899 B.n450 B.n447 10.6151
R900 B.n447 B.n446 10.6151
R901 B.n446 B.n443 10.6151
R902 B.n443 B.n442 10.6151
R903 B.n442 B.n439 10.6151
R904 B.n439 B.n438 10.6151
R905 B.n438 B.n435 10.6151
R906 B.n435 B.n434 10.6151
R907 B.n434 B.n431 10.6151
R908 B.n431 B.n430 10.6151
R909 B.n430 B.n427 10.6151
R910 B.n427 B.n426 10.6151
R911 B.n426 B.n423 10.6151
R912 B.n423 B.n422 10.6151
R913 B.n422 B.n419 10.6151
R914 B.n419 B.n418 10.6151
R915 B.n418 B.n415 10.6151
R916 B.n415 B.n414 10.6151
R917 B.n414 B.n411 10.6151
R918 B.n411 B.n410 10.6151
R919 B.n410 B.n407 10.6151
R920 B.n407 B.n406 10.6151
R921 B.n406 B.n403 10.6151
R922 B.n403 B.n402 10.6151
R923 B.n402 B.n399 10.6151
R924 B.n399 B.n398 10.6151
R925 B.n395 B.n394 10.6151
R926 B.n394 B.n391 10.6151
R927 B.n391 B.n390 10.6151
R928 B.n390 B.n387 10.6151
R929 B.n387 B.n386 10.6151
R930 B.n386 B.n383 10.6151
R931 B.n383 B.n382 10.6151
R932 B.n382 B.n379 10.6151
R933 B.n377 B.n374 10.6151
R934 B.n374 B.n373 10.6151
R935 B.n373 B.n370 10.6151
R936 B.n370 B.n369 10.6151
R937 B.n369 B.n366 10.6151
R938 B.n366 B.n365 10.6151
R939 B.n365 B.n362 10.6151
R940 B.n362 B.n361 10.6151
R941 B.n361 B.n358 10.6151
R942 B.n358 B.n357 10.6151
R943 B.n357 B.n354 10.6151
R944 B.n354 B.n353 10.6151
R945 B.n353 B.n350 10.6151
R946 B.n350 B.n349 10.6151
R947 B.n349 B.n346 10.6151
R948 B.n346 B.n345 10.6151
R949 B.n345 B.n342 10.6151
R950 B.n342 B.n341 10.6151
R951 B.n341 B.n338 10.6151
R952 B.n338 B.n337 10.6151
R953 B.n337 B.n334 10.6151
R954 B.n334 B.n333 10.6151
R955 B.n333 B.n330 10.6151
R956 B.n330 B.n329 10.6151
R957 B.n329 B.n326 10.6151
R958 B.n326 B.n325 10.6151
R959 B.n325 B.n322 10.6151
R960 B.n322 B.n321 10.6151
R961 B.n321 B.n318 10.6151
R962 B.n318 B.n317 10.6151
R963 B.n317 B.n272 10.6151
R964 B.n465 B.n272 10.6151
R965 B.n471 B.n268 10.6151
R966 B.n472 B.n471 10.6151
R967 B.n473 B.n472 10.6151
R968 B.n473 B.n260 10.6151
R969 B.n484 B.n260 10.6151
R970 B.n485 B.n484 10.6151
R971 B.n486 B.n485 10.6151
R972 B.n486 B.n253 10.6151
R973 B.n496 B.n253 10.6151
R974 B.n497 B.n496 10.6151
R975 B.n498 B.n497 10.6151
R976 B.n498 B.n245 10.6151
R977 B.n508 B.n245 10.6151
R978 B.n509 B.n508 10.6151
R979 B.n510 B.n509 10.6151
R980 B.n510 B.n237 10.6151
R981 B.n521 B.n237 10.6151
R982 B.n522 B.n521 10.6151
R983 B.n523 B.n522 10.6151
R984 B.n523 B.n0 10.6151
R985 B.n596 B.n1 10.6151
R986 B.n596 B.n595 10.6151
R987 B.n595 B.n594 10.6151
R988 B.n594 B.n10 10.6151
R989 B.n588 B.n10 10.6151
R990 B.n588 B.n587 10.6151
R991 B.n587 B.n586 10.6151
R992 B.n586 B.n17 10.6151
R993 B.n580 B.n17 10.6151
R994 B.n580 B.n579 10.6151
R995 B.n579 B.n578 10.6151
R996 B.n578 B.n24 10.6151
R997 B.n572 B.n24 10.6151
R998 B.n572 B.n571 10.6151
R999 B.n571 B.n570 10.6151
R1000 B.n570 B.n30 10.6151
R1001 B.n564 B.n30 10.6151
R1002 B.n564 B.n563 10.6151
R1003 B.n563 B.n562 10.6151
R1004 B.n562 B.n38 10.6151
R1005 B.n243 B.t1 9.293
R1006 B.t0 B.n591 9.293
R1007 B.n152 B.n151 6.5566
R1008 B.n168 B.n82 6.5566
R1009 B.n395 B.n313 6.5566
R1010 B.n379 B.n378 6.5566
R1011 B.n151 B.n150 4.05904
R1012 B.n171 B.n82 4.05904
R1013 B.n398 B.n313 4.05904
R1014 B.n378 B.n377 4.05904
R1015 B.n602 B.n0 2.81026
R1016 B.n602 B.n1 2.81026
R1017 VP.n0 VP.t0 214.935
R1018 VP.n0 VP.t1 174.567
R1019 VP VP.n0 0.241678
R1020 VTAIL.n1 VTAIL.t1 49.7185
R1021 VTAIL.n3 VTAIL.t0 49.7182
R1022 VTAIL.n0 VTAIL.t3 49.7182
R1023 VTAIL.n2 VTAIL.t2 49.7182
R1024 VTAIL.n1 VTAIL.n0 23.841
R1025 VTAIL.n3 VTAIL.n2 21.9531
R1026 VTAIL.n2 VTAIL.n1 1.41429
R1027 VTAIL VTAIL.n0 1.0005
R1028 VTAIL VTAIL.n3 0.414293
R1029 VDD1 VDD1.t0 102.528
R1030 VDD1 VDD1.t1 66.9272
R1031 VN VN.t0 215.126
R1032 VN VN.t1 174.809
R1033 VDD2.n0 VDD2.t0 101.531
R1034 VDD2.n0 VDD2.t1 66.397
R1035 VDD2 VDD2.n0 0.530672
C0 VN VDD1 0.147783f
C1 VP VDD2 0.301739f
C2 VDD2 VTAIL 4.20006f
C3 VDD1 VDD2 0.586639f
C4 VN VDD2 2.01163f
C5 VP VTAIL 1.77271f
C6 VP VDD1 2.16326f
C7 VDD1 VTAIL 4.15444f
C8 VN VP 4.53993f
C9 VN VTAIL 1.75841f
C10 VDD2 B 3.619661f
C11 VDD1 B 6.38337f
C12 VTAIL B 5.749966f
C13 VN B 8.38649f
C14 VP B 5.260527f
C15 VDD2.t0 B 2.01859f
C16 VDD2.t1 B 1.59884f
C17 VDD2.n0 B 2.48516f
C18 VN.t1 B 1.56137f
C19 VN.t0 B 1.87535f
C20 VDD1.t1 B 1.63269f
C21 VDD1.t0 B 2.0884f
C22 VTAIL.t3 B 1.12733f
C23 VTAIL.n0 B 0.998356f
C24 VTAIL.t1 B 1.12734f
C25 VTAIL.n1 B 1.0184f
C26 VTAIL.t2 B 1.12733f
C27 VTAIL.n2 B 0.926925f
C28 VTAIL.t0 B 1.12733f
C29 VTAIL.n3 B 0.87847f
C30 VP.t0 B 1.94166f
C31 VP.t1 B 1.61917f
C32 VP.n0 B 3.09041f
.ends

