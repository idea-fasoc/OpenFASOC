* NGSPICE file created from diff_pair_sample_0186.ext - technology: sky130A

.subckt diff_pair_sample_0186 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t11 VN.t0 VDD2.t1 B.t4 sky130_fd_pr__nfet_01v8 ad=1.48005 pd=9.3 as=1.48005 ps=9.3 w=8.97 l=2.2
X1 VDD1.t5 VP.t0 VTAIL.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=3.4983 pd=18.72 as=1.48005 ps=9.3 w=8.97 l=2.2
X2 VDD1.t4 VP.t1 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=1.48005 pd=9.3 as=3.4983 ps=18.72 w=8.97 l=2.2
X3 VTAIL.t10 VN.t1 VDD2.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=1.48005 pd=9.3 as=1.48005 ps=9.3 w=8.97 l=2.2
X4 VTAIL.t4 VP.t2 VDD1.t3 B.t4 sky130_fd_pr__nfet_01v8 ad=1.48005 pd=9.3 as=1.48005 ps=9.3 w=8.97 l=2.2
X5 B.t19 B.t17 B.t18 B.t7 sky130_fd_pr__nfet_01v8 ad=3.4983 pd=18.72 as=0 ps=0 w=8.97 l=2.2
X6 B.t16 B.t14 B.t15 B.t11 sky130_fd_pr__nfet_01v8 ad=3.4983 pd=18.72 as=0 ps=0 w=8.97 l=2.2
X7 VDD2.t5 VN.t2 VTAIL.t9 B.t1 sky130_fd_pr__nfet_01v8 ad=1.48005 pd=9.3 as=3.4983 ps=18.72 w=8.97 l=2.2
X8 VDD2.t4 VN.t3 VTAIL.t8 B.t5 sky130_fd_pr__nfet_01v8 ad=3.4983 pd=18.72 as=1.48005 ps=9.3 w=8.97 l=2.2
X9 VDD1.t2 VP.t3 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=1.48005 pd=9.3 as=3.4983 ps=18.72 w=8.97 l=2.2
X10 VDD1.t1 VP.t4 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=3.4983 pd=18.72 as=1.48005 ps=9.3 w=8.97 l=2.2
X11 B.t13 B.t10 B.t12 B.t11 sky130_fd_pr__nfet_01v8 ad=3.4983 pd=18.72 as=0 ps=0 w=8.97 l=2.2
X12 VTAIL.t3 VP.t5 VDD1.t0 B.t3 sky130_fd_pr__nfet_01v8 ad=1.48005 pd=9.3 as=1.48005 ps=9.3 w=8.97 l=2.2
X13 VDD2.t2 VN.t4 VTAIL.t7 B.t2 sky130_fd_pr__nfet_01v8 ad=3.4983 pd=18.72 as=1.48005 ps=9.3 w=8.97 l=2.2
X14 VDD2.t0 VN.t5 VTAIL.t6 B.t0 sky130_fd_pr__nfet_01v8 ad=1.48005 pd=9.3 as=3.4983 ps=18.72 w=8.97 l=2.2
X15 B.t9 B.t6 B.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=3.4983 pd=18.72 as=0 ps=0 w=8.97 l=2.2
R0 VN.n25 VN.n14 161.3
R1 VN.n24 VN.n23 161.3
R2 VN.n22 VN.n15 161.3
R3 VN.n21 VN.n20 161.3
R4 VN.n19 VN.n16 161.3
R5 VN.n11 VN.n0 161.3
R6 VN.n10 VN.n9 161.3
R7 VN.n8 VN.n1 161.3
R8 VN.n7 VN.n6 161.3
R9 VN.n5 VN.n2 161.3
R10 VN.n3 VN.t3 130.69
R11 VN.n17 VN.t2 130.69
R12 VN.n4 VN.t1 98.2628
R13 VN.n12 VN.t5 98.2628
R14 VN.n18 VN.t0 98.2628
R15 VN.n26 VN.t4 98.2628
R16 VN.n13 VN.n12 97.0549
R17 VN.n27 VN.n26 97.0549
R18 VN.n4 VN.n3 59.2585
R19 VN.n18 VN.n17 59.2585
R20 VN VN.n27 45.0701
R21 VN.n10 VN.n1 41.9503
R22 VN.n24 VN.n15 41.9503
R23 VN.n6 VN.n1 39.0365
R24 VN.n20 VN.n15 39.0365
R25 VN.n6 VN.n5 24.4675
R26 VN.n11 VN.n10 24.4675
R27 VN.n20 VN.n19 24.4675
R28 VN.n25 VN.n24 24.4675
R29 VN.n12 VN.n11 13.702
R30 VN.n26 VN.n25 13.702
R31 VN.n5 VN.n4 12.234
R32 VN.n19 VN.n18 12.234
R33 VN.n17 VN.n16 9.58252
R34 VN.n3 VN.n2 9.58252
R35 VN.n27 VN.n14 0.278367
R36 VN.n13 VN.n0 0.278367
R37 VN.n23 VN.n14 0.189894
R38 VN.n23 VN.n22 0.189894
R39 VN.n22 VN.n21 0.189894
R40 VN.n21 VN.n16 0.189894
R41 VN.n7 VN.n2 0.189894
R42 VN.n8 VN.n7 0.189894
R43 VN.n9 VN.n8 0.189894
R44 VN.n9 VN.n0 0.189894
R45 VN VN.n13 0.153454
R46 VDD2.n1 VDD2.t4 68.7433
R47 VDD2.n2 VDD2.t2 67.1631
R48 VDD2.n1 VDD2.n0 65.4454
R49 VDD2 VDD2.n3 65.4427
R50 VDD2.n2 VDD2.n1 38.5364
R51 VDD2.n3 VDD2.t1 2.20786
R52 VDD2.n3 VDD2.t5 2.20786
R53 VDD2.n0 VDD2.t3 2.20786
R54 VDD2.n0 VDD2.t0 2.20786
R55 VDD2 VDD2.n2 1.69447
R56 VTAIL.n7 VTAIL.t9 50.4843
R57 VTAIL.n11 VTAIL.t6 50.4841
R58 VTAIL.n2 VTAIL.t1 50.4841
R59 VTAIL.n10 VTAIL.t0 50.4841
R60 VTAIL.n9 VTAIL.n8 48.277
R61 VTAIL.n6 VTAIL.n5 48.277
R62 VTAIL.n1 VTAIL.n0 48.2767
R63 VTAIL.n4 VTAIL.n3 48.2767
R64 VTAIL.n6 VTAIL.n4 24.4617
R65 VTAIL.n11 VTAIL.n10 22.2807
R66 VTAIL.n0 VTAIL.t8 2.20786
R67 VTAIL.n0 VTAIL.t10 2.20786
R68 VTAIL.n3 VTAIL.t2 2.20786
R69 VTAIL.n3 VTAIL.t4 2.20786
R70 VTAIL.n8 VTAIL.t5 2.20786
R71 VTAIL.n8 VTAIL.t3 2.20786
R72 VTAIL.n5 VTAIL.t7 2.20786
R73 VTAIL.n5 VTAIL.t11 2.20786
R74 VTAIL.n7 VTAIL.n6 2.18153
R75 VTAIL.n10 VTAIL.n9 2.18153
R76 VTAIL.n4 VTAIL.n2 2.18153
R77 VTAIL VTAIL.n11 1.57809
R78 VTAIL.n9 VTAIL.n7 1.56084
R79 VTAIL.n2 VTAIL.n1 1.56084
R80 VTAIL VTAIL.n1 0.603948
R81 B.n544 B.n114 585
R82 B.n114 B.n71 585
R83 B.n546 B.n545 585
R84 B.n548 B.n113 585
R85 B.n551 B.n550 585
R86 B.n552 B.n112 585
R87 B.n554 B.n553 585
R88 B.n556 B.n111 585
R89 B.n559 B.n558 585
R90 B.n560 B.n110 585
R91 B.n562 B.n561 585
R92 B.n564 B.n109 585
R93 B.n567 B.n566 585
R94 B.n568 B.n108 585
R95 B.n570 B.n569 585
R96 B.n572 B.n107 585
R97 B.n575 B.n574 585
R98 B.n576 B.n106 585
R99 B.n578 B.n577 585
R100 B.n580 B.n105 585
R101 B.n583 B.n582 585
R102 B.n584 B.n104 585
R103 B.n586 B.n585 585
R104 B.n588 B.n103 585
R105 B.n591 B.n590 585
R106 B.n592 B.n102 585
R107 B.n594 B.n593 585
R108 B.n596 B.n101 585
R109 B.n599 B.n598 585
R110 B.n600 B.n100 585
R111 B.n602 B.n601 585
R112 B.n604 B.n99 585
R113 B.n606 B.n605 585
R114 B.n608 B.n607 585
R115 B.n611 B.n610 585
R116 B.n612 B.n94 585
R117 B.n614 B.n613 585
R118 B.n616 B.n93 585
R119 B.n619 B.n618 585
R120 B.n620 B.n92 585
R121 B.n622 B.n621 585
R122 B.n624 B.n91 585
R123 B.n627 B.n626 585
R124 B.n629 B.n88 585
R125 B.n631 B.n630 585
R126 B.n633 B.n87 585
R127 B.n636 B.n635 585
R128 B.n637 B.n86 585
R129 B.n639 B.n638 585
R130 B.n641 B.n85 585
R131 B.n644 B.n643 585
R132 B.n645 B.n84 585
R133 B.n647 B.n646 585
R134 B.n649 B.n83 585
R135 B.n652 B.n651 585
R136 B.n653 B.n82 585
R137 B.n655 B.n654 585
R138 B.n657 B.n81 585
R139 B.n660 B.n659 585
R140 B.n661 B.n80 585
R141 B.n663 B.n662 585
R142 B.n665 B.n79 585
R143 B.n668 B.n667 585
R144 B.n669 B.n78 585
R145 B.n671 B.n670 585
R146 B.n673 B.n77 585
R147 B.n676 B.n675 585
R148 B.n677 B.n76 585
R149 B.n679 B.n678 585
R150 B.n681 B.n75 585
R151 B.n684 B.n683 585
R152 B.n685 B.n74 585
R153 B.n687 B.n686 585
R154 B.n689 B.n73 585
R155 B.n692 B.n691 585
R156 B.n693 B.n72 585
R157 B.n543 B.n70 585
R158 B.n696 B.n70 585
R159 B.n542 B.n69 585
R160 B.n697 B.n69 585
R161 B.n541 B.n68 585
R162 B.n698 B.n68 585
R163 B.n540 B.n539 585
R164 B.n539 B.n64 585
R165 B.n538 B.n63 585
R166 B.n704 B.n63 585
R167 B.n537 B.n62 585
R168 B.n705 B.n62 585
R169 B.n536 B.n61 585
R170 B.n706 B.n61 585
R171 B.n535 B.n534 585
R172 B.n534 B.n60 585
R173 B.n533 B.n56 585
R174 B.n712 B.n56 585
R175 B.n532 B.n55 585
R176 B.n713 B.n55 585
R177 B.n531 B.n54 585
R178 B.n714 B.n54 585
R179 B.n530 B.n529 585
R180 B.n529 B.n50 585
R181 B.n528 B.n49 585
R182 B.n720 B.n49 585
R183 B.n527 B.n48 585
R184 B.n721 B.n48 585
R185 B.n526 B.n47 585
R186 B.n722 B.n47 585
R187 B.n525 B.n524 585
R188 B.n524 B.n43 585
R189 B.n523 B.n42 585
R190 B.n728 B.n42 585
R191 B.n522 B.n41 585
R192 B.n729 B.n41 585
R193 B.n521 B.n40 585
R194 B.n730 B.n40 585
R195 B.n520 B.n519 585
R196 B.n519 B.n36 585
R197 B.n518 B.n35 585
R198 B.n736 B.n35 585
R199 B.n517 B.n34 585
R200 B.n737 B.n34 585
R201 B.n516 B.n33 585
R202 B.n738 B.n33 585
R203 B.n515 B.n514 585
R204 B.n514 B.n29 585
R205 B.n513 B.n28 585
R206 B.n744 B.n28 585
R207 B.n512 B.n27 585
R208 B.n745 B.n27 585
R209 B.n511 B.n26 585
R210 B.n746 B.n26 585
R211 B.n510 B.n509 585
R212 B.n509 B.n22 585
R213 B.n508 B.n21 585
R214 B.n752 B.n21 585
R215 B.n507 B.n20 585
R216 B.n753 B.n20 585
R217 B.n506 B.n19 585
R218 B.n754 B.n19 585
R219 B.n505 B.n504 585
R220 B.n504 B.n15 585
R221 B.n503 B.n14 585
R222 B.n760 B.n14 585
R223 B.n502 B.n13 585
R224 B.n761 B.n13 585
R225 B.n501 B.n12 585
R226 B.n762 B.n12 585
R227 B.n500 B.n499 585
R228 B.n499 B.n8 585
R229 B.n498 B.n7 585
R230 B.n768 B.n7 585
R231 B.n497 B.n6 585
R232 B.n769 B.n6 585
R233 B.n496 B.n5 585
R234 B.n770 B.n5 585
R235 B.n495 B.n494 585
R236 B.n494 B.n4 585
R237 B.n493 B.n115 585
R238 B.n493 B.n492 585
R239 B.n483 B.n116 585
R240 B.n117 B.n116 585
R241 B.n485 B.n484 585
R242 B.n486 B.n485 585
R243 B.n482 B.n122 585
R244 B.n122 B.n121 585
R245 B.n481 B.n480 585
R246 B.n480 B.n479 585
R247 B.n124 B.n123 585
R248 B.n125 B.n124 585
R249 B.n472 B.n471 585
R250 B.n473 B.n472 585
R251 B.n470 B.n130 585
R252 B.n130 B.n129 585
R253 B.n469 B.n468 585
R254 B.n468 B.n467 585
R255 B.n132 B.n131 585
R256 B.n133 B.n132 585
R257 B.n460 B.n459 585
R258 B.n461 B.n460 585
R259 B.n458 B.n137 585
R260 B.n141 B.n137 585
R261 B.n457 B.n456 585
R262 B.n456 B.n455 585
R263 B.n139 B.n138 585
R264 B.n140 B.n139 585
R265 B.n448 B.n447 585
R266 B.n449 B.n448 585
R267 B.n446 B.n146 585
R268 B.n146 B.n145 585
R269 B.n445 B.n444 585
R270 B.n444 B.n443 585
R271 B.n148 B.n147 585
R272 B.n149 B.n148 585
R273 B.n436 B.n435 585
R274 B.n437 B.n436 585
R275 B.n434 B.n153 585
R276 B.n157 B.n153 585
R277 B.n433 B.n432 585
R278 B.n432 B.n431 585
R279 B.n155 B.n154 585
R280 B.n156 B.n155 585
R281 B.n424 B.n423 585
R282 B.n425 B.n424 585
R283 B.n422 B.n162 585
R284 B.n162 B.n161 585
R285 B.n421 B.n420 585
R286 B.n420 B.n419 585
R287 B.n164 B.n163 585
R288 B.n165 B.n164 585
R289 B.n412 B.n411 585
R290 B.n413 B.n412 585
R291 B.n410 B.n170 585
R292 B.n170 B.n169 585
R293 B.n409 B.n408 585
R294 B.n408 B.n407 585
R295 B.n172 B.n171 585
R296 B.n400 B.n172 585
R297 B.n399 B.n398 585
R298 B.n401 B.n399 585
R299 B.n397 B.n177 585
R300 B.n177 B.n176 585
R301 B.n396 B.n395 585
R302 B.n395 B.n394 585
R303 B.n179 B.n178 585
R304 B.n180 B.n179 585
R305 B.n387 B.n386 585
R306 B.n388 B.n387 585
R307 B.n385 B.n185 585
R308 B.n185 B.n184 585
R309 B.n384 B.n383 585
R310 B.n383 B.n382 585
R311 B.n379 B.n189 585
R312 B.n378 B.n377 585
R313 B.n375 B.n190 585
R314 B.n375 B.n188 585
R315 B.n374 B.n373 585
R316 B.n372 B.n371 585
R317 B.n370 B.n192 585
R318 B.n368 B.n367 585
R319 B.n366 B.n193 585
R320 B.n365 B.n364 585
R321 B.n362 B.n194 585
R322 B.n360 B.n359 585
R323 B.n358 B.n195 585
R324 B.n357 B.n356 585
R325 B.n354 B.n196 585
R326 B.n352 B.n351 585
R327 B.n350 B.n197 585
R328 B.n349 B.n348 585
R329 B.n346 B.n198 585
R330 B.n344 B.n343 585
R331 B.n342 B.n199 585
R332 B.n341 B.n340 585
R333 B.n338 B.n200 585
R334 B.n336 B.n335 585
R335 B.n334 B.n201 585
R336 B.n333 B.n332 585
R337 B.n330 B.n202 585
R338 B.n328 B.n327 585
R339 B.n326 B.n203 585
R340 B.n325 B.n324 585
R341 B.n322 B.n204 585
R342 B.n320 B.n319 585
R343 B.n318 B.n205 585
R344 B.n317 B.n316 585
R345 B.n314 B.n313 585
R346 B.n312 B.n311 585
R347 B.n310 B.n210 585
R348 B.n308 B.n307 585
R349 B.n306 B.n211 585
R350 B.n305 B.n304 585
R351 B.n302 B.n212 585
R352 B.n300 B.n299 585
R353 B.n298 B.n213 585
R354 B.n296 B.n295 585
R355 B.n293 B.n216 585
R356 B.n291 B.n290 585
R357 B.n289 B.n217 585
R358 B.n288 B.n287 585
R359 B.n285 B.n218 585
R360 B.n283 B.n282 585
R361 B.n281 B.n219 585
R362 B.n280 B.n279 585
R363 B.n277 B.n220 585
R364 B.n275 B.n274 585
R365 B.n273 B.n221 585
R366 B.n272 B.n271 585
R367 B.n269 B.n222 585
R368 B.n267 B.n266 585
R369 B.n265 B.n223 585
R370 B.n264 B.n263 585
R371 B.n261 B.n224 585
R372 B.n259 B.n258 585
R373 B.n257 B.n225 585
R374 B.n256 B.n255 585
R375 B.n253 B.n226 585
R376 B.n251 B.n250 585
R377 B.n249 B.n227 585
R378 B.n248 B.n247 585
R379 B.n245 B.n228 585
R380 B.n243 B.n242 585
R381 B.n241 B.n229 585
R382 B.n240 B.n239 585
R383 B.n237 B.n230 585
R384 B.n235 B.n234 585
R385 B.n233 B.n232 585
R386 B.n187 B.n186 585
R387 B.n381 B.n380 585
R388 B.n382 B.n381 585
R389 B.n183 B.n182 585
R390 B.n184 B.n183 585
R391 B.n390 B.n389 585
R392 B.n389 B.n388 585
R393 B.n391 B.n181 585
R394 B.n181 B.n180 585
R395 B.n393 B.n392 585
R396 B.n394 B.n393 585
R397 B.n175 B.n174 585
R398 B.n176 B.n175 585
R399 B.n403 B.n402 585
R400 B.n402 B.n401 585
R401 B.n404 B.n173 585
R402 B.n400 B.n173 585
R403 B.n406 B.n405 585
R404 B.n407 B.n406 585
R405 B.n168 B.n167 585
R406 B.n169 B.n168 585
R407 B.n415 B.n414 585
R408 B.n414 B.n413 585
R409 B.n416 B.n166 585
R410 B.n166 B.n165 585
R411 B.n418 B.n417 585
R412 B.n419 B.n418 585
R413 B.n160 B.n159 585
R414 B.n161 B.n160 585
R415 B.n427 B.n426 585
R416 B.n426 B.n425 585
R417 B.n428 B.n158 585
R418 B.n158 B.n156 585
R419 B.n430 B.n429 585
R420 B.n431 B.n430 585
R421 B.n152 B.n151 585
R422 B.n157 B.n152 585
R423 B.n439 B.n438 585
R424 B.n438 B.n437 585
R425 B.n440 B.n150 585
R426 B.n150 B.n149 585
R427 B.n442 B.n441 585
R428 B.n443 B.n442 585
R429 B.n144 B.n143 585
R430 B.n145 B.n144 585
R431 B.n451 B.n450 585
R432 B.n450 B.n449 585
R433 B.n452 B.n142 585
R434 B.n142 B.n140 585
R435 B.n454 B.n453 585
R436 B.n455 B.n454 585
R437 B.n136 B.n135 585
R438 B.n141 B.n136 585
R439 B.n463 B.n462 585
R440 B.n462 B.n461 585
R441 B.n464 B.n134 585
R442 B.n134 B.n133 585
R443 B.n466 B.n465 585
R444 B.n467 B.n466 585
R445 B.n128 B.n127 585
R446 B.n129 B.n128 585
R447 B.n475 B.n474 585
R448 B.n474 B.n473 585
R449 B.n476 B.n126 585
R450 B.n126 B.n125 585
R451 B.n478 B.n477 585
R452 B.n479 B.n478 585
R453 B.n120 B.n119 585
R454 B.n121 B.n120 585
R455 B.n488 B.n487 585
R456 B.n487 B.n486 585
R457 B.n489 B.n118 585
R458 B.n118 B.n117 585
R459 B.n491 B.n490 585
R460 B.n492 B.n491 585
R461 B.n2 B.n0 585
R462 B.n4 B.n2 585
R463 B.n3 B.n1 585
R464 B.n769 B.n3 585
R465 B.n767 B.n766 585
R466 B.n768 B.n767 585
R467 B.n765 B.n9 585
R468 B.n9 B.n8 585
R469 B.n764 B.n763 585
R470 B.n763 B.n762 585
R471 B.n11 B.n10 585
R472 B.n761 B.n11 585
R473 B.n759 B.n758 585
R474 B.n760 B.n759 585
R475 B.n757 B.n16 585
R476 B.n16 B.n15 585
R477 B.n756 B.n755 585
R478 B.n755 B.n754 585
R479 B.n18 B.n17 585
R480 B.n753 B.n18 585
R481 B.n751 B.n750 585
R482 B.n752 B.n751 585
R483 B.n749 B.n23 585
R484 B.n23 B.n22 585
R485 B.n748 B.n747 585
R486 B.n747 B.n746 585
R487 B.n25 B.n24 585
R488 B.n745 B.n25 585
R489 B.n743 B.n742 585
R490 B.n744 B.n743 585
R491 B.n741 B.n30 585
R492 B.n30 B.n29 585
R493 B.n740 B.n739 585
R494 B.n739 B.n738 585
R495 B.n32 B.n31 585
R496 B.n737 B.n32 585
R497 B.n735 B.n734 585
R498 B.n736 B.n735 585
R499 B.n733 B.n37 585
R500 B.n37 B.n36 585
R501 B.n732 B.n731 585
R502 B.n731 B.n730 585
R503 B.n39 B.n38 585
R504 B.n729 B.n39 585
R505 B.n727 B.n726 585
R506 B.n728 B.n727 585
R507 B.n725 B.n44 585
R508 B.n44 B.n43 585
R509 B.n724 B.n723 585
R510 B.n723 B.n722 585
R511 B.n46 B.n45 585
R512 B.n721 B.n46 585
R513 B.n719 B.n718 585
R514 B.n720 B.n719 585
R515 B.n717 B.n51 585
R516 B.n51 B.n50 585
R517 B.n716 B.n715 585
R518 B.n715 B.n714 585
R519 B.n53 B.n52 585
R520 B.n713 B.n53 585
R521 B.n711 B.n710 585
R522 B.n712 B.n711 585
R523 B.n709 B.n57 585
R524 B.n60 B.n57 585
R525 B.n708 B.n707 585
R526 B.n707 B.n706 585
R527 B.n59 B.n58 585
R528 B.n705 B.n59 585
R529 B.n703 B.n702 585
R530 B.n704 B.n703 585
R531 B.n701 B.n65 585
R532 B.n65 B.n64 585
R533 B.n700 B.n699 585
R534 B.n699 B.n698 585
R535 B.n67 B.n66 585
R536 B.n697 B.n67 585
R537 B.n695 B.n694 585
R538 B.n696 B.n695 585
R539 B.n772 B.n771 585
R540 B.n771 B.n770 585
R541 B.n381 B.n189 478.086
R542 B.n695 B.n72 478.086
R543 B.n383 B.n187 478.086
R544 B.n114 B.n70 478.086
R545 B.n214 B.t17 305.613
R546 B.n206 B.t6 305.613
R547 B.n89 B.t14 305.613
R548 B.n95 B.t10 305.613
R549 B.n547 B.n71 256.663
R550 B.n549 B.n71 256.663
R551 B.n555 B.n71 256.663
R552 B.n557 B.n71 256.663
R553 B.n563 B.n71 256.663
R554 B.n565 B.n71 256.663
R555 B.n571 B.n71 256.663
R556 B.n573 B.n71 256.663
R557 B.n579 B.n71 256.663
R558 B.n581 B.n71 256.663
R559 B.n587 B.n71 256.663
R560 B.n589 B.n71 256.663
R561 B.n595 B.n71 256.663
R562 B.n597 B.n71 256.663
R563 B.n603 B.n71 256.663
R564 B.n98 B.n71 256.663
R565 B.n609 B.n71 256.663
R566 B.n615 B.n71 256.663
R567 B.n617 B.n71 256.663
R568 B.n623 B.n71 256.663
R569 B.n625 B.n71 256.663
R570 B.n632 B.n71 256.663
R571 B.n634 B.n71 256.663
R572 B.n640 B.n71 256.663
R573 B.n642 B.n71 256.663
R574 B.n648 B.n71 256.663
R575 B.n650 B.n71 256.663
R576 B.n656 B.n71 256.663
R577 B.n658 B.n71 256.663
R578 B.n664 B.n71 256.663
R579 B.n666 B.n71 256.663
R580 B.n672 B.n71 256.663
R581 B.n674 B.n71 256.663
R582 B.n680 B.n71 256.663
R583 B.n682 B.n71 256.663
R584 B.n688 B.n71 256.663
R585 B.n690 B.n71 256.663
R586 B.n376 B.n188 256.663
R587 B.n191 B.n188 256.663
R588 B.n369 B.n188 256.663
R589 B.n363 B.n188 256.663
R590 B.n361 B.n188 256.663
R591 B.n355 B.n188 256.663
R592 B.n353 B.n188 256.663
R593 B.n347 B.n188 256.663
R594 B.n345 B.n188 256.663
R595 B.n339 B.n188 256.663
R596 B.n337 B.n188 256.663
R597 B.n331 B.n188 256.663
R598 B.n329 B.n188 256.663
R599 B.n323 B.n188 256.663
R600 B.n321 B.n188 256.663
R601 B.n315 B.n188 256.663
R602 B.n209 B.n188 256.663
R603 B.n309 B.n188 256.663
R604 B.n303 B.n188 256.663
R605 B.n301 B.n188 256.663
R606 B.n294 B.n188 256.663
R607 B.n292 B.n188 256.663
R608 B.n286 B.n188 256.663
R609 B.n284 B.n188 256.663
R610 B.n278 B.n188 256.663
R611 B.n276 B.n188 256.663
R612 B.n270 B.n188 256.663
R613 B.n268 B.n188 256.663
R614 B.n262 B.n188 256.663
R615 B.n260 B.n188 256.663
R616 B.n254 B.n188 256.663
R617 B.n252 B.n188 256.663
R618 B.n246 B.n188 256.663
R619 B.n244 B.n188 256.663
R620 B.n238 B.n188 256.663
R621 B.n236 B.n188 256.663
R622 B.n231 B.n188 256.663
R623 B.n381 B.n183 163.367
R624 B.n389 B.n183 163.367
R625 B.n389 B.n181 163.367
R626 B.n393 B.n181 163.367
R627 B.n393 B.n175 163.367
R628 B.n402 B.n175 163.367
R629 B.n402 B.n173 163.367
R630 B.n406 B.n173 163.367
R631 B.n406 B.n168 163.367
R632 B.n414 B.n168 163.367
R633 B.n414 B.n166 163.367
R634 B.n418 B.n166 163.367
R635 B.n418 B.n160 163.367
R636 B.n426 B.n160 163.367
R637 B.n426 B.n158 163.367
R638 B.n430 B.n158 163.367
R639 B.n430 B.n152 163.367
R640 B.n438 B.n152 163.367
R641 B.n438 B.n150 163.367
R642 B.n442 B.n150 163.367
R643 B.n442 B.n144 163.367
R644 B.n450 B.n144 163.367
R645 B.n450 B.n142 163.367
R646 B.n454 B.n142 163.367
R647 B.n454 B.n136 163.367
R648 B.n462 B.n136 163.367
R649 B.n462 B.n134 163.367
R650 B.n466 B.n134 163.367
R651 B.n466 B.n128 163.367
R652 B.n474 B.n128 163.367
R653 B.n474 B.n126 163.367
R654 B.n478 B.n126 163.367
R655 B.n478 B.n120 163.367
R656 B.n487 B.n120 163.367
R657 B.n487 B.n118 163.367
R658 B.n491 B.n118 163.367
R659 B.n491 B.n2 163.367
R660 B.n771 B.n2 163.367
R661 B.n771 B.n3 163.367
R662 B.n767 B.n3 163.367
R663 B.n767 B.n9 163.367
R664 B.n763 B.n9 163.367
R665 B.n763 B.n11 163.367
R666 B.n759 B.n11 163.367
R667 B.n759 B.n16 163.367
R668 B.n755 B.n16 163.367
R669 B.n755 B.n18 163.367
R670 B.n751 B.n18 163.367
R671 B.n751 B.n23 163.367
R672 B.n747 B.n23 163.367
R673 B.n747 B.n25 163.367
R674 B.n743 B.n25 163.367
R675 B.n743 B.n30 163.367
R676 B.n739 B.n30 163.367
R677 B.n739 B.n32 163.367
R678 B.n735 B.n32 163.367
R679 B.n735 B.n37 163.367
R680 B.n731 B.n37 163.367
R681 B.n731 B.n39 163.367
R682 B.n727 B.n39 163.367
R683 B.n727 B.n44 163.367
R684 B.n723 B.n44 163.367
R685 B.n723 B.n46 163.367
R686 B.n719 B.n46 163.367
R687 B.n719 B.n51 163.367
R688 B.n715 B.n51 163.367
R689 B.n715 B.n53 163.367
R690 B.n711 B.n53 163.367
R691 B.n711 B.n57 163.367
R692 B.n707 B.n57 163.367
R693 B.n707 B.n59 163.367
R694 B.n703 B.n59 163.367
R695 B.n703 B.n65 163.367
R696 B.n699 B.n65 163.367
R697 B.n699 B.n67 163.367
R698 B.n695 B.n67 163.367
R699 B.n377 B.n375 163.367
R700 B.n375 B.n374 163.367
R701 B.n371 B.n370 163.367
R702 B.n368 B.n193 163.367
R703 B.n364 B.n362 163.367
R704 B.n360 B.n195 163.367
R705 B.n356 B.n354 163.367
R706 B.n352 B.n197 163.367
R707 B.n348 B.n346 163.367
R708 B.n344 B.n199 163.367
R709 B.n340 B.n338 163.367
R710 B.n336 B.n201 163.367
R711 B.n332 B.n330 163.367
R712 B.n328 B.n203 163.367
R713 B.n324 B.n322 163.367
R714 B.n320 B.n205 163.367
R715 B.n316 B.n314 163.367
R716 B.n311 B.n310 163.367
R717 B.n308 B.n211 163.367
R718 B.n304 B.n302 163.367
R719 B.n300 B.n213 163.367
R720 B.n295 B.n293 163.367
R721 B.n291 B.n217 163.367
R722 B.n287 B.n285 163.367
R723 B.n283 B.n219 163.367
R724 B.n279 B.n277 163.367
R725 B.n275 B.n221 163.367
R726 B.n271 B.n269 163.367
R727 B.n267 B.n223 163.367
R728 B.n263 B.n261 163.367
R729 B.n259 B.n225 163.367
R730 B.n255 B.n253 163.367
R731 B.n251 B.n227 163.367
R732 B.n247 B.n245 163.367
R733 B.n243 B.n229 163.367
R734 B.n239 B.n237 163.367
R735 B.n235 B.n232 163.367
R736 B.n383 B.n185 163.367
R737 B.n387 B.n185 163.367
R738 B.n387 B.n179 163.367
R739 B.n395 B.n179 163.367
R740 B.n395 B.n177 163.367
R741 B.n399 B.n177 163.367
R742 B.n399 B.n172 163.367
R743 B.n408 B.n172 163.367
R744 B.n408 B.n170 163.367
R745 B.n412 B.n170 163.367
R746 B.n412 B.n164 163.367
R747 B.n420 B.n164 163.367
R748 B.n420 B.n162 163.367
R749 B.n424 B.n162 163.367
R750 B.n424 B.n155 163.367
R751 B.n432 B.n155 163.367
R752 B.n432 B.n153 163.367
R753 B.n436 B.n153 163.367
R754 B.n436 B.n148 163.367
R755 B.n444 B.n148 163.367
R756 B.n444 B.n146 163.367
R757 B.n448 B.n146 163.367
R758 B.n448 B.n139 163.367
R759 B.n456 B.n139 163.367
R760 B.n456 B.n137 163.367
R761 B.n460 B.n137 163.367
R762 B.n460 B.n132 163.367
R763 B.n468 B.n132 163.367
R764 B.n468 B.n130 163.367
R765 B.n472 B.n130 163.367
R766 B.n472 B.n124 163.367
R767 B.n480 B.n124 163.367
R768 B.n480 B.n122 163.367
R769 B.n485 B.n122 163.367
R770 B.n485 B.n116 163.367
R771 B.n493 B.n116 163.367
R772 B.n494 B.n493 163.367
R773 B.n494 B.n5 163.367
R774 B.n6 B.n5 163.367
R775 B.n7 B.n6 163.367
R776 B.n499 B.n7 163.367
R777 B.n499 B.n12 163.367
R778 B.n13 B.n12 163.367
R779 B.n14 B.n13 163.367
R780 B.n504 B.n14 163.367
R781 B.n504 B.n19 163.367
R782 B.n20 B.n19 163.367
R783 B.n21 B.n20 163.367
R784 B.n509 B.n21 163.367
R785 B.n509 B.n26 163.367
R786 B.n27 B.n26 163.367
R787 B.n28 B.n27 163.367
R788 B.n514 B.n28 163.367
R789 B.n514 B.n33 163.367
R790 B.n34 B.n33 163.367
R791 B.n35 B.n34 163.367
R792 B.n519 B.n35 163.367
R793 B.n519 B.n40 163.367
R794 B.n41 B.n40 163.367
R795 B.n42 B.n41 163.367
R796 B.n524 B.n42 163.367
R797 B.n524 B.n47 163.367
R798 B.n48 B.n47 163.367
R799 B.n49 B.n48 163.367
R800 B.n529 B.n49 163.367
R801 B.n529 B.n54 163.367
R802 B.n55 B.n54 163.367
R803 B.n56 B.n55 163.367
R804 B.n534 B.n56 163.367
R805 B.n534 B.n61 163.367
R806 B.n62 B.n61 163.367
R807 B.n63 B.n62 163.367
R808 B.n539 B.n63 163.367
R809 B.n539 B.n68 163.367
R810 B.n69 B.n68 163.367
R811 B.n70 B.n69 163.367
R812 B.n691 B.n689 163.367
R813 B.n687 B.n74 163.367
R814 B.n683 B.n681 163.367
R815 B.n679 B.n76 163.367
R816 B.n675 B.n673 163.367
R817 B.n671 B.n78 163.367
R818 B.n667 B.n665 163.367
R819 B.n663 B.n80 163.367
R820 B.n659 B.n657 163.367
R821 B.n655 B.n82 163.367
R822 B.n651 B.n649 163.367
R823 B.n647 B.n84 163.367
R824 B.n643 B.n641 163.367
R825 B.n639 B.n86 163.367
R826 B.n635 B.n633 163.367
R827 B.n631 B.n88 163.367
R828 B.n626 B.n624 163.367
R829 B.n622 B.n92 163.367
R830 B.n618 B.n616 163.367
R831 B.n614 B.n94 163.367
R832 B.n610 B.n608 163.367
R833 B.n605 B.n604 163.367
R834 B.n602 B.n100 163.367
R835 B.n598 B.n596 163.367
R836 B.n594 B.n102 163.367
R837 B.n590 B.n588 163.367
R838 B.n586 B.n104 163.367
R839 B.n582 B.n580 163.367
R840 B.n578 B.n106 163.367
R841 B.n574 B.n572 163.367
R842 B.n570 B.n108 163.367
R843 B.n566 B.n564 163.367
R844 B.n562 B.n110 163.367
R845 B.n558 B.n556 163.367
R846 B.n554 B.n112 163.367
R847 B.n550 B.n548 163.367
R848 B.n546 B.n114 163.367
R849 B.n214 B.t19 119.93
R850 B.n95 B.t12 119.93
R851 B.n206 B.t9 119.921
R852 B.n89 B.t15 119.921
R853 B.n382 B.n188 88.8036
R854 B.n696 B.n71 88.8036
R855 B.n376 B.n189 71.676
R856 B.n374 B.n191 71.676
R857 B.n370 B.n369 71.676
R858 B.n363 B.n193 71.676
R859 B.n362 B.n361 71.676
R860 B.n355 B.n195 71.676
R861 B.n354 B.n353 71.676
R862 B.n347 B.n197 71.676
R863 B.n346 B.n345 71.676
R864 B.n339 B.n199 71.676
R865 B.n338 B.n337 71.676
R866 B.n331 B.n201 71.676
R867 B.n330 B.n329 71.676
R868 B.n323 B.n203 71.676
R869 B.n322 B.n321 71.676
R870 B.n315 B.n205 71.676
R871 B.n314 B.n209 71.676
R872 B.n310 B.n309 71.676
R873 B.n303 B.n211 71.676
R874 B.n302 B.n301 71.676
R875 B.n294 B.n213 71.676
R876 B.n293 B.n292 71.676
R877 B.n286 B.n217 71.676
R878 B.n285 B.n284 71.676
R879 B.n278 B.n219 71.676
R880 B.n277 B.n276 71.676
R881 B.n270 B.n221 71.676
R882 B.n269 B.n268 71.676
R883 B.n262 B.n223 71.676
R884 B.n261 B.n260 71.676
R885 B.n254 B.n225 71.676
R886 B.n253 B.n252 71.676
R887 B.n246 B.n227 71.676
R888 B.n245 B.n244 71.676
R889 B.n238 B.n229 71.676
R890 B.n237 B.n236 71.676
R891 B.n232 B.n231 71.676
R892 B.n690 B.n72 71.676
R893 B.n689 B.n688 71.676
R894 B.n682 B.n74 71.676
R895 B.n681 B.n680 71.676
R896 B.n674 B.n76 71.676
R897 B.n673 B.n672 71.676
R898 B.n666 B.n78 71.676
R899 B.n665 B.n664 71.676
R900 B.n658 B.n80 71.676
R901 B.n657 B.n656 71.676
R902 B.n650 B.n82 71.676
R903 B.n649 B.n648 71.676
R904 B.n642 B.n84 71.676
R905 B.n641 B.n640 71.676
R906 B.n634 B.n86 71.676
R907 B.n633 B.n632 71.676
R908 B.n625 B.n88 71.676
R909 B.n624 B.n623 71.676
R910 B.n617 B.n92 71.676
R911 B.n616 B.n615 71.676
R912 B.n609 B.n94 71.676
R913 B.n608 B.n98 71.676
R914 B.n604 B.n603 71.676
R915 B.n597 B.n100 71.676
R916 B.n596 B.n595 71.676
R917 B.n589 B.n102 71.676
R918 B.n588 B.n587 71.676
R919 B.n581 B.n104 71.676
R920 B.n580 B.n579 71.676
R921 B.n573 B.n106 71.676
R922 B.n572 B.n571 71.676
R923 B.n565 B.n108 71.676
R924 B.n564 B.n563 71.676
R925 B.n557 B.n110 71.676
R926 B.n556 B.n555 71.676
R927 B.n549 B.n112 71.676
R928 B.n548 B.n547 71.676
R929 B.n547 B.n546 71.676
R930 B.n550 B.n549 71.676
R931 B.n555 B.n554 71.676
R932 B.n558 B.n557 71.676
R933 B.n563 B.n562 71.676
R934 B.n566 B.n565 71.676
R935 B.n571 B.n570 71.676
R936 B.n574 B.n573 71.676
R937 B.n579 B.n578 71.676
R938 B.n582 B.n581 71.676
R939 B.n587 B.n586 71.676
R940 B.n590 B.n589 71.676
R941 B.n595 B.n594 71.676
R942 B.n598 B.n597 71.676
R943 B.n603 B.n602 71.676
R944 B.n605 B.n98 71.676
R945 B.n610 B.n609 71.676
R946 B.n615 B.n614 71.676
R947 B.n618 B.n617 71.676
R948 B.n623 B.n622 71.676
R949 B.n626 B.n625 71.676
R950 B.n632 B.n631 71.676
R951 B.n635 B.n634 71.676
R952 B.n640 B.n639 71.676
R953 B.n643 B.n642 71.676
R954 B.n648 B.n647 71.676
R955 B.n651 B.n650 71.676
R956 B.n656 B.n655 71.676
R957 B.n659 B.n658 71.676
R958 B.n664 B.n663 71.676
R959 B.n667 B.n666 71.676
R960 B.n672 B.n671 71.676
R961 B.n675 B.n674 71.676
R962 B.n680 B.n679 71.676
R963 B.n683 B.n682 71.676
R964 B.n688 B.n687 71.676
R965 B.n691 B.n690 71.676
R966 B.n377 B.n376 71.676
R967 B.n371 B.n191 71.676
R968 B.n369 B.n368 71.676
R969 B.n364 B.n363 71.676
R970 B.n361 B.n360 71.676
R971 B.n356 B.n355 71.676
R972 B.n353 B.n352 71.676
R973 B.n348 B.n347 71.676
R974 B.n345 B.n344 71.676
R975 B.n340 B.n339 71.676
R976 B.n337 B.n336 71.676
R977 B.n332 B.n331 71.676
R978 B.n329 B.n328 71.676
R979 B.n324 B.n323 71.676
R980 B.n321 B.n320 71.676
R981 B.n316 B.n315 71.676
R982 B.n311 B.n209 71.676
R983 B.n309 B.n308 71.676
R984 B.n304 B.n303 71.676
R985 B.n301 B.n300 71.676
R986 B.n295 B.n294 71.676
R987 B.n292 B.n291 71.676
R988 B.n287 B.n286 71.676
R989 B.n284 B.n283 71.676
R990 B.n279 B.n278 71.676
R991 B.n276 B.n275 71.676
R992 B.n271 B.n270 71.676
R993 B.n268 B.n267 71.676
R994 B.n263 B.n262 71.676
R995 B.n260 B.n259 71.676
R996 B.n255 B.n254 71.676
R997 B.n252 B.n251 71.676
R998 B.n247 B.n246 71.676
R999 B.n244 B.n243 71.676
R1000 B.n239 B.n238 71.676
R1001 B.n236 B.n235 71.676
R1002 B.n231 B.n187 71.676
R1003 B.n215 B.t18 70.8641
R1004 B.n96 B.t13 70.8641
R1005 B.n207 B.t8 70.8534
R1006 B.n90 B.t16 70.8534
R1007 B.n297 B.n215 59.5399
R1008 B.n208 B.n207 59.5399
R1009 B.n628 B.n90 59.5399
R1010 B.n97 B.n96 59.5399
R1011 B.n382 B.n184 52.5102
R1012 B.n388 B.n184 52.5102
R1013 B.n388 B.n180 52.5102
R1014 B.n394 B.n180 52.5102
R1015 B.n394 B.n176 52.5102
R1016 B.n401 B.n176 52.5102
R1017 B.n401 B.n400 52.5102
R1018 B.n407 B.n169 52.5102
R1019 B.n413 B.n169 52.5102
R1020 B.n413 B.n165 52.5102
R1021 B.n419 B.n165 52.5102
R1022 B.n419 B.n161 52.5102
R1023 B.n425 B.n161 52.5102
R1024 B.n425 B.n156 52.5102
R1025 B.n431 B.n156 52.5102
R1026 B.n431 B.n157 52.5102
R1027 B.n437 B.n149 52.5102
R1028 B.n443 B.n149 52.5102
R1029 B.n443 B.n145 52.5102
R1030 B.n449 B.n145 52.5102
R1031 B.n449 B.n140 52.5102
R1032 B.n455 B.n140 52.5102
R1033 B.n455 B.n141 52.5102
R1034 B.n461 B.n133 52.5102
R1035 B.n467 B.n133 52.5102
R1036 B.n467 B.n129 52.5102
R1037 B.n473 B.n129 52.5102
R1038 B.n473 B.n125 52.5102
R1039 B.n479 B.n125 52.5102
R1040 B.n486 B.n121 52.5102
R1041 B.n486 B.n117 52.5102
R1042 B.n492 B.n117 52.5102
R1043 B.n492 B.n4 52.5102
R1044 B.n770 B.n4 52.5102
R1045 B.n770 B.n769 52.5102
R1046 B.n769 B.n768 52.5102
R1047 B.n768 B.n8 52.5102
R1048 B.n762 B.n8 52.5102
R1049 B.n762 B.n761 52.5102
R1050 B.n760 B.n15 52.5102
R1051 B.n754 B.n15 52.5102
R1052 B.n754 B.n753 52.5102
R1053 B.n753 B.n752 52.5102
R1054 B.n752 B.n22 52.5102
R1055 B.n746 B.n22 52.5102
R1056 B.n745 B.n744 52.5102
R1057 B.n744 B.n29 52.5102
R1058 B.n738 B.n29 52.5102
R1059 B.n738 B.n737 52.5102
R1060 B.n737 B.n736 52.5102
R1061 B.n736 B.n36 52.5102
R1062 B.n730 B.n36 52.5102
R1063 B.n729 B.n728 52.5102
R1064 B.n728 B.n43 52.5102
R1065 B.n722 B.n43 52.5102
R1066 B.n722 B.n721 52.5102
R1067 B.n721 B.n720 52.5102
R1068 B.n720 B.n50 52.5102
R1069 B.n714 B.n50 52.5102
R1070 B.n714 B.n713 52.5102
R1071 B.n713 B.n712 52.5102
R1072 B.n706 B.n60 52.5102
R1073 B.n706 B.n705 52.5102
R1074 B.n705 B.n704 52.5102
R1075 B.n704 B.n64 52.5102
R1076 B.n698 B.n64 52.5102
R1077 B.n698 B.n697 52.5102
R1078 B.n697 B.n696 52.5102
R1079 B.n215 B.n214 49.0672
R1080 B.n207 B.n206 49.0672
R1081 B.n90 B.n89 49.0672
R1082 B.n96 B.n95 49.0672
R1083 B.n407 B.t7 44.7881
R1084 B.n712 B.t11 44.7881
R1085 B.n157 B.t2 41.6993
R1086 B.t0 B.n729 41.6993
R1087 B.n461 B.t4 40.1549
R1088 B.n746 B.t3 40.1549
R1089 B.n479 B.t1 35.5217
R1090 B.t5 B.n760 35.5217
R1091 B.n694 B.n693 31.0639
R1092 B.n544 B.n543 31.0639
R1093 B.n384 B.n186 31.0639
R1094 B.n380 B.n379 31.0639
R1095 B B.n772 18.0485
R1096 B.t1 B.n121 16.9889
R1097 B.n761 B.t5 16.9889
R1098 B.n141 B.t4 12.3557
R1099 B.t3 B.n745 12.3557
R1100 B.n437 B.t2 10.8113
R1101 B.n730 B.t0 10.8113
R1102 B.n693 B.n692 10.6151
R1103 B.n692 B.n73 10.6151
R1104 B.n686 B.n73 10.6151
R1105 B.n686 B.n685 10.6151
R1106 B.n685 B.n684 10.6151
R1107 B.n684 B.n75 10.6151
R1108 B.n678 B.n75 10.6151
R1109 B.n678 B.n677 10.6151
R1110 B.n677 B.n676 10.6151
R1111 B.n676 B.n77 10.6151
R1112 B.n670 B.n77 10.6151
R1113 B.n670 B.n669 10.6151
R1114 B.n669 B.n668 10.6151
R1115 B.n668 B.n79 10.6151
R1116 B.n662 B.n79 10.6151
R1117 B.n662 B.n661 10.6151
R1118 B.n661 B.n660 10.6151
R1119 B.n660 B.n81 10.6151
R1120 B.n654 B.n81 10.6151
R1121 B.n654 B.n653 10.6151
R1122 B.n653 B.n652 10.6151
R1123 B.n652 B.n83 10.6151
R1124 B.n646 B.n83 10.6151
R1125 B.n646 B.n645 10.6151
R1126 B.n645 B.n644 10.6151
R1127 B.n644 B.n85 10.6151
R1128 B.n638 B.n85 10.6151
R1129 B.n638 B.n637 10.6151
R1130 B.n637 B.n636 10.6151
R1131 B.n636 B.n87 10.6151
R1132 B.n630 B.n87 10.6151
R1133 B.n630 B.n629 10.6151
R1134 B.n627 B.n91 10.6151
R1135 B.n621 B.n91 10.6151
R1136 B.n621 B.n620 10.6151
R1137 B.n620 B.n619 10.6151
R1138 B.n619 B.n93 10.6151
R1139 B.n613 B.n93 10.6151
R1140 B.n613 B.n612 10.6151
R1141 B.n612 B.n611 10.6151
R1142 B.n607 B.n606 10.6151
R1143 B.n606 B.n99 10.6151
R1144 B.n601 B.n99 10.6151
R1145 B.n601 B.n600 10.6151
R1146 B.n600 B.n599 10.6151
R1147 B.n599 B.n101 10.6151
R1148 B.n593 B.n101 10.6151
R1149 B.n593 B.n592 10.6151
R1150 B.n592 B.n591 10.6151
R1151 B.n591 B.n103 10.6151
R1152 B.n585 B.n103 10.6151
R1153 B.n585 B.n584 10.6151
R1154 B.n584 B.n583 10.6151
R1155 B.n583 B.n105 10.6151
R1156 B.n577 B.n105 10.6151
R1157 B.n577 B.n576 10.6151
R1158 B.n576 B.n575 10.6151
R1159 B.n575 B.n107 10.6151
R1160 B.n569 B.n107 10.6151
R1161 B.n569 B.n568 10.6151
R1162 B.n568 B.n567 10.6151
R1163 B.n567 B.n109 10.6151
R1164 B.n561 B.n109 10.6151
R1165 B.n561 B.n560 10.6151
R1166 B.n560 B.n559 10.6151
R1167 B.n559 B.n111 10.6151
R1168 B.n553 B.n111 10.6151
R1169 B.n553 B.n552 10.6151
R1170 B.n552 B.n551 10.6151
R1171 B.n551 B.n113 10.6151
R1172 B.n545 B.n113 10.6151
R1173 B.n545 B.n544 10.6151
R1174 B.n385 B.n384 10.6151
R1175 B.n386 B.n385 10.6151
R1176 B.n386 B.n178 10.6151
R1177 B.n396 B.n178 10.6151
R1178 B.n397 B.n396 10.6151
R1179 B.n398 B.n397 10.6151
R1180 B.n398 B.n171 10.6151
R1181 B.n409 B.n171 10.6151
R1182 B.n410 B.n409 10.6151
R1183 B.n411 B.n410 10.6151
R1184 B.n411 B.n163 10.6151
R1185 B.n421 B.n163 10.6151
R1186 B.n422 B.n421 10.6151
R1187 B.n423 B.n422 10.6151
R1188 B.n423 B.n154 10.6151
R1189 B.n433 B.n154 10.6151
R1190 B.n434 B.n433 10.6151
R1191 B.n435 B.n434 10.6151
R1192 B.n435 B.n147 10.6151
R1193 B.n445 B.n147 10.6151
R1194 B.n446 B.n445 10.6151
R1195 B.n447 B.n446 10.6151
R1196 B.n447 B.n138 10.6151
R1197 B.n457 B.n138 10.6151
R1198 B.n458 B.n457 10.6151
R1199 B.n459 B.n458 10.6151
R1200 B.n459 B.n131 10.6151
R1201 B.n469 B.n131 10.6151
R1202 B.n470 B.n469 10.6151
R1203 B.n471 B.n470 10.6151
R1204 B.n471 B.n123 10.6151
R1205 B.n481 B.n123 10.6151
R1206 B.n482 B.n481 10.6151
R1207 B.n484 B.n482 10.6151
R1208 B.n484 B.n483 10.6151
R1209 B.n483 B.n115 10.6151
R1210 B.n495 B.n115 10.6151
R1211 B.n496 B.n495 10.6151
R1212 B.n497 B.n496 10.6151
R1213 B.n498 B.n497 10.6151
R1214 B.n500 B.n498 10.6151
R1215 B.n501 B.n500 10.6151
R1216 B.n502 B.n501 10.6151
R1217 B.n503 B.n502 10.6151
R1218 B.n505 B.n503 10.6151
R1219 B.n506 B.n505 10.6151
R1220 B.n507 B.n506 10.6151
R1221 B.n508 B.n507 10.6151
R1222 B.n510 B.n508 10.6151
R1223 B.n511 B.n510 10.6151
R1224 B.n512 B.n511 10.6151
R1225 B.n513 B.n512 10.6151
R1226 B.n515 B.n513 10.6151
R1227 B.n516 B.n515 10.6151
R1228 B.n517 B.n516 10.6151
R1229 B.n518 B.n517 10.6151
R1230 B.n520 B.n518 10.6151
R1231 B.n521 B.n520 10.6151
R1232 B.n522 B.n521 10.6151
R1233 B.n523 B.n522 10.6151
R1234 B.n525 B.n523 10.6151
R1235 B.n526 B.n525 10.6151
R1236 B.n527 B.n526 10.6151
R1237 B.n528 B.n527 10.6151
R1238 B.n530 B.n528 10.6151
R1239 B.n531 B.n530 10.6151
R1240 B.n532 B.n531 10.6151
R1241 B.n533 B.n532 10.6151
R1242 B.n535 B.n533 10.6151
R1243 B.n536 B.n535 10.6151
R1244 B.n537 B.n536 10.6151
R1245 B.n538 B.n537 10.6151
R1246 B.n540 B.n538 10.6151
R1247 B.n541 B.n540 10.6151
R1248 B.n542 B.n541 10.6151
R1249 B.n543 B.n542 10.6151
R1250 B.n379 B.n378 10.6151
R1251 B.n378 B.n190 10.6151
R1252 B.n373 B.n190 10.6151
R1253 B.n373 B.n372 10.6151
R1254 B.n372 B.n192 10.6151
R1255 B.n367 B.n192 10.6151
R1256 B.n367 B.n366 10.6151
R1257 B.n366 B.n365 10.6151
R1258 B.n365 B.n194 10.6151
R1259 B.n359 B.n194 10.6151
R1260 B.n359 B.n358 10.6151
R1261 B.n358 B.n357 10.6151
R1262 B.n357 B.n196 10.6151
R1263 B.n351 B.n196 10.6151
R1264 B.n351 B.n350 10.6151
R1265 B.n350 B.n349 10.6151
R1266 B.n349 B.n198 10.6151
R1267 B.n343 B.n198 10.6151
R1268 B.n343 B.n342 10.6151
R1269 B.n342 B.n341 10.6151
R1270 B.n341 B.n200 10.6151
R1271 B.n335 B.n200 10.6151
R1272 B.n335 B.n334 10.6151
R1273 B.n334 B.n333 10.6151
R1274 B.n333 B.n202 10.6151
R1275 B.n327 B.n202 10.6151
R1276 B.n327 B.n326 10.6151
R1277 B.n326 B.n325 10.6151
R1278 B.n325 B.n204 10.6151
R1279 B.n319 B.n204 10.6151
R1280 B.n319 B.n318 10.6151
R1281 B.n318 B.n317 10.6151
R1282 B.n313 B.n312 10.6151
R1283 B.n312 B.n210 10.6151
R1284 B.n307 B.n210 10.6151
R1285 B.n307 B.n306 10.6151
R1286 B.n306 B.n305 10.6151
R1287 B.n305 B.n212 10.6151
R1288 B.n299 B.n212 10.6151
R1289 B.n299 B.n298 10.6151
R1290 B.n296 B.n216 10.6151
R1291 B.n290 B.n216 10.6151
R1292 B.n290 B.n289 10.6151
R1293 B.n289 B.n288 10.6151
R1294 B.n288 B.n218 10.6151
R1295 B.n282 B.n218 10.6151
R1296 B.n282 B.n281 10.6151
R1297 B.n281 B.n280 10.6151
R1298 B.n280 B.n220 10.6151
R1299 B.n274 B.n220 10.6151
R1300 B.n274 B.n273 10.6151
R1301 B.n273 B.n272 10.6151
R1302 B.n272 B.n222 10.6151
R1303 B.n266 B.n222 10.6151
R1304 B.n266 B.n265 10.6151
R1305 B.n265 B.n264 10.6151
R1306 B.n264 B.n224 10.6151
R1307 B.n258 B.n224 10.6151
R1308 B.n258 B.n257 10.6151
R1309 B.n257 B.n256 10.6151
R1310 B.n256 B.n226 10.6151
R1311 B.n250 B.n226 10.6151
R1312 B.n250 B.n249 10.6151
R1313 B.n249 B.n248 10.6151
R1314 B.n248 B.n228 10.6151
R1315 B.n242 B.n228 10.6151
R1316 B.n242 B.n241 10.6151
R1317 B.n241 B.n240 10.6151
R1318 B.n240 B.n230 10.6151
R1319 B.n234 B.n230 10.6151
R1320 B.n234 B.n233 10.6151
R1321 B.n233 B.n186 10.6151
R1322 B.n380 B.n182 10.6151
R1323 B.n390 B.n182 10.6151
R1324 B.n391 B.n390 10.6151
R1325 B.n392 B.n391 10.6151
R1326 B.n392 B.n174 10.6151
R1327 B.n403 B.n174 10.6151
R1328 B.n404 B.n403 10.6151
R1329 B.n405 B.n404 10.6151
R1330 B.n405 B.n167 10.6151
R1331 B.n415 B.n167 10.6151
R1332 B.n416 B.n415 10.6151
R1333 B.n417 B.n416 10.6151
R1334 B.n417 B.n159 10.6151
R1335 B.n427 B.n159 10.6151
R1336 B.n428 B.n427 10.6151
R1337 B.n429 B.n428 10.6151
R1338 B.n429 B.n151 10.6151
R1339 B.n439 B.n151 10.6151
R1340 B.n440 B.n439 10.6151
R1341 B.n441 B.n440 10.6151
R1342 B.n441 B.n143 10.6151
R1343 B.n451 B.n143 10.6151
R1344 B.n452 B.n451 10.6151
R1345 B.n453 B.n452 10.6151
R1346 B.n453 B.n135 10.6151
R1347 B.n463 B.n135 10.6151
R1348 B.n464 B.n463 10.6151
R1349 B.n465 B.n464 10.6151
R1350 B.n465 B.n127 10.6151
R1351 B.n475 B.n127 10.6151
R1352 B.n476 B.n475 10.6151
R1353 B.n477 B.n476 10.6151
R1354 B.n477 B.n119 10.6151
R1355 B.n488 B.n119 10.6151
R1356 B.n489 B.n488 10.6151
R1357 B.n490 B.n489 10.6151
R1358 B.n490 B.n0 10.6151
R1359 B.n766 B.n1 10.6151
R1360 B.n766 B.n765 10.6151
R1361 B.n765 B.n764 10.6151
R1362 B.n764 B.n10 10.6151
R1363 B.n758 B.n10 10.6151
R1364 B.n758 B.n757 10.6151
R1365 B.n757 B.n756 10.6151
R1366 B.n756 B.n17 10.6151
R1367 B.n750 B.n17 10.6151
R1368 B.n750 B.n749 10.6151
R1369 B.n749 B.n748 10.6151
R1370 B.n748 B.n24 10.6151
R1371 B.n742 B.n24 10.6151
R1372 B.n742 B.n741 10.6151
R1373 B.n741 B.n740 10.6151
R1374 B.n740 B.n31 10.6151
R1375 B.n734 B.n31 10.6151
R1376 B.n734 B.n733 10.6151
R1377 B.n733 B.n732 10.6151
R1378 B.n732 B.n38 10.6151
R1379 B.n726 B.n38 10.6151
R1380 B.n726 B.n725 10.6151
R1381 B.n725 B.n724 10.6151
R1382 B.n724 B.n45 10.6151
R1383 B.n718 B.n45 10.6151
R1384 B.n718 B.n717 10.6151
R1385 B.n717 B.n716 10.6151
R1386 B.n716 B.n52 10.6151
R1387 B.n710 B.n52 10.6151
R1388 B.n710 B.n709 10.6151
R1389 B.n709 B.n708 10.6151
R1390 B.n708 B.n58 10.6151
R1391 B.n702 B.n58 10.6151
R1392 B.n702 B.n701 10.6151
R1393 B.n701 B.n700 10.6151
R1394 B.n700 B.n66 10.6151
R1395 B.n694 B.n66 10.6151
R1396 B.n400 B.t7 7.72251
R1397 B.n60 B.t11 7.72251
R1398 B.n628 B.n627 6.5566
R1399 B.n611 B.n97 6.5566
R1400 B.n313 B.n208 6.5566
R1401 B.n298 B.n297 6.5566
R1402 B.n629 B.n628 4.05904
R1403 B.n607 B.n97 4.05904
R1404 B.n317 B.n208 4.05904
R1405 B.n297 B.n296 4.05904
R1406 B.n772 B.n0 2.81026
R1407 B.n772 B.n1 2.81026
R1408 VP.n11 VP.n8 161.3
R1409 VP.n13 VP.n12 161.3
R1410 VP.n14 VP.n7 161.3
R1411 VP.n16 VP.n15 161.3
R1412 VP.n17 VP.n6 161.3
R1413 VP.n36 VP.n0 161.3
R1414 VP.n35 VP.n34 161.3
R1415 VP.n33 VP.n1 161.3
R1416 VP.n32 VP.n31 161.3
R1417 VP.n30 VP.n2 161.3
R1418 VP.n28 VP.n27 161.3
R1419 VP.n26 VP.n3 161.3
R1420 VP.n25 VP.n24 161.3
R1421 VP.n23 VP.n4 161.3
R1422 VP.n22 VP.n21 161.3
R1423 VP.n9 VP.t0 130.69
R1424 VP.n5 VP.t4 98.2628
R1425 VP.n29 VP.t2 98.2628
R1426 VP.n37 VP.t3 98.2628
R1427 VP.n18 VP.t1 98.2628
R1428 VP.n10 VP.t5 98.2628
R1429 VP.n20 VP.n5 97.0549
R1430 VP.n38 VP.n37 97.0549
R1431 VP.n19 VP.n18 97.0549
R1432 VP.n10 VP.n9 59.2585
R1433 VP.n20 VP.n19 44.7913
R1434 VP.n24 VP.n23 41.9503
R1435 VP.n35 VP.n1 41.9503
R1436 VP.n16 VP.n7 41.9503
R1437 VP.n24 VP.n3 39.0365
R1438 VP.n31 VP.n1 39.0365
R1439 VP.n12 VP.n7 39.0365
R1440 VP.n23 VP.n22 24.4675
R1441 VP.n28 VP.n3 24.4675
R1442 VP.n31 VP.n30 24.4675
R1443 VP.n36 VP.n35 24.4675
R1444 VP.n17 VP.n16 24.4675
R1445 VP.n12 VP.n11 24.4675
R1446 VP.n22 VP.n5 13.702
R1447 VP.n37 VP.n36 13.702
R1448 VP.n18 VP.n17 13.702
R1449 VP.n29 VP.n28 12.234
R1450 VP.n30 VP.n29 12.234
R1451 VP.n11 VP.n10 12.234
R1452 VP.n9 VP.n8 9.58252
R1453 VP.n19 VP.n6 0.278367
R1454 VP.n21 VP.n20 0.278367
R1455 VP.n38 VP.n0 0.278367
R1456 VP.n13 VP.n8 0.189894
R1457 VP.n14 VP.n13 0.189894
R1458 VP.n15 VP.n14 0.189894
R1459 VP.n15 VP.n6 0.189894
R1460 VP.n21 VP.n4 0.189894
R1461 VP.n25 VP.n4 0.189894
R1462 VP.n26 VP.n25 0.189894
R1463 VP.n27 VP.n26 0.189894
R1464 VP.n27 VP.n2 0.189894
R1465 VP.n32 VP.n2 0.189894
R1466 VP.n33 VP.n32 0.189894
R1467 VP.n34 VP.n33 0.189894
R1468 VP.n34 VP.n0 0.189894
R1469 VP VP.n38 0.153454
R1470 VDD1 VDD1.t5 68.8571
R1471 VDD1.n1 VDD1.t1 68.7433
R1472 VDD1.n1 VDD1.n0 65.4454
R1473 VDD1.n3 VDD1.n2 64.9556
R1474 VDD1.n3 VDD1.n1 40.2099
R1475 VDD1.n2 VDD1.t0 2.20786
R1476 VDD1.n2 VDD1.t4 2.20786
R1477 VDD1.n0 VDD1.t3 2.20786
R1478 VDD1.n0 VDD1.t2 2.20786
R1479 VDD1 VDD1.n3 0.487569
C0 VN VDD1 0.149994f
C1 VDD2 VP 0.423959f
C2 VTAIL VDD1 6.53037f
C3 VDD2 VDD1 1.24944f
C4 VDD1 VP 5.22626f
C5 VTAIL VN 5.1501f
C6 VDD2 VN 4.95502f
C7 VN VP 5.97954f
C8 VTAIL VDD2 6.57886f
C9 VTAIL VP 5.16437f
C10 VDD2 B 5.141494f
C11 VDD1 B 5.437647f
C12 VTAIL B 6.343787f
C13 VN B 11.49759f
C14 VP B 10.108589f
C15 VDD1.t5 B 1.72618f
C16 VDD1.t1 B 1.72543f
C17 VDD1.t3 B 0.154371f
C18 VDD1.t2 B 0.154371f
C19 VDD1.n0 B 1.35232f
C20 VDD1.n1 B 2.3055f
C21 VDD1.t0 B 0.154371f
C22 VDD1.t4 B 0.154371f
C23 VDD1.n2 B 1.34954f
C24 VDD1.n3 B 2.12374f
C25 VP.n0 B 0.036089f
C26 VP.t3 B 1.4576f
C27 VP.n1 B 0.022209f
C28 VP.n2 B 0.027373f
C29 VP.t2 B 1.4576f
C30 VP.n3 B 0.054777f
C31 VP.n4 B 0.027373f
C32 VP.t4 B 1.4576f
C33 VP.n5 B 0.612118f
C34 VP.n6 B 0.036089f
C35 VP.t1 B 1.4576f
C36 VP.n7 B 0.022209f
C37 VP.n8 B 0.233009f
C38 VP.t5 B 1.4576f
C39 VP.t0 B 1.62544f
C40 VP.n9 B 0.592041f
C41 VP.n10 B 0.600426f
C42 VP.n11 B 0.038423f
C43 VP.n12 B 0.054777f
C44 VP.n13 B 0.027373f
C45 VP.n14 B 0.027373f
C46 VP.n15 B 0.027373f
C47 VP.n16 B 0.053956f
C48 VP.n17 B 0.039935f
C49 VP.n18 B 0.612118f
C50 VP.n19 B 1.28328f
C51 VP.n20 B 1.30525f
C52 VP.n21 B 0.036089f
C53 VP.n22 B 0.039935f
C54 VP.n23 B 0.053956f
C55 VP.n24 B 0.022209f
C56 VP.n25 B 0.027373f
C57 VP.n26 B 0.027373f
C58 VP.n27 B 0.027373f
C59 VP.n28 B 0.038423f
C60 VP.n29 B 0.529805f
C61 VP.n30 B 0.038423f
C62 VP.n31 B 0.054777f
C63 VP.n32 B 0.027373f
C64 VP.n33 B 0.027373f
C65 VP.n34 B 0.027373f
C66 VP.n35 B 0.053956f
C67 VP.n36 B 0.039935f
C68 VP.n37 B 0.612118f
C69 VP.n38 B 0.038842f
C70 VTAIL.t8 B 0.174317f
C71 VTAIL.t10 B 0.174317f
C72 VTAIL.n0 B 1.45736f
C73 VTAIL.n1 B 0.40191f
C74 VTAIL.t1 B 1.85588f
C75 VTAIL.n2 B 0.603806f
C76 VTAIL.t2 B 0.174317f
C77 VTAIL.t4 B 0.174317f
C78 VTAIL.n3 B 1.45736f
C79 VTAIL.n4 B 1.69574f
C80 VTAIL.t7 B 0.174317f
C81 VTAIL.t11 B 0.174317f
C82 VTAIL.n5 B 1.45736f
C83 VTAIL.n6 B 1.69573f
C84 VTAIL.t9 B 1.85588f
C85 VTAIL.n7 B 0.603802f
C86 VTAIL.t5 B 0.174317f
C87 VTAIL.t3 B 0.174317f
C88 VTAIL.n8 B 1.45736f
C89 VTAIL.n9 B 0.526915f
C90 VTAIL.t0 B 1.85588f
C91 VTAIL.n10 B 1.5998f
C92 VTAIL.t6 B 1.85588f
C93 VTAIL.n11 B 1.55198f
C94 VDD2.t4 B 1.72253f
C95 VDD2.t3 B 0.154111f
C96 VDD2.t0 B 0.154111f
C97 VDD2.n0 B 1.35005f
C98 VDD2.n1 B 2.20468f
C99 VDD2.t2 B 1.71455f
C100 VDD2.n2 B 2.12157f
C101 VDD2.t1 B 0.154111f
C102 VDD2.t5 B 0.154111f
C103 VDD2.n3 B 1.35002f
C104 VN.n0 B 0.035565f
C105 VN.t5 B 1.43645f
C106 VN.n1 B 0.021887f
C107 VN.n2 B 0.229629f
C108 VN.t1 B 1.43645f
C109 VN.t3 B 1.60185f
C110 VN.n3 B 0.583452f
C111 VN.n4 B 0.591716f
C112 VN.n5 B 0.037866f
C113 VN.n6 B 0.053983f
C114 VN.n7 B 0.026976f
C115 VN.n8 B 0.026976f
C116 VN.n9 B 0.026976f
C117 VN.n10 B 0.053173f
C118 VN.n11 B 0.039355f
C119 VN.n12 B 0.603238f
C120 VN.n13 B 0.038279f
C121 VN.n14 B 0.035565f
C122 VN.t4 B 1.43645f
C123 VN.n15 B 0.021887f
C124 VN.n16 B 0.229629f
C125 VN.t0 B 1.43645f
C126 VN.t2 B 1.60185f
C127 VN.n17 B 0.583452f
C128 VN.n18 B 0.591716f
C129 VN.n19 B 0.037866f
C130 VN.n20 B 0.053983f
C131 VN.n21 B 0.026976f
C132 VN.n22 B 0.026976f
C133 VN.n23 B 0.026976f
C134 VN.n24 B 0.053173f
C135 VN.n25 B 0.039355f
C136 VN.n26 B 0.603238f
C137 VN.n27 B 1.27943f
.ends

