* NGSPICE file created from diff_pair_sample_0549.ext - technology: sky130A

.subckt diff_pair_sample_0549 VTAIL VN VP B VDD2 VDD1
X0 B.t11 B.t9 B.t10 w_n5506_n4706# sky130_fd_pr__pfet_01v8 ad=7.2891 pd=38.16 as=0 ps=0 w=18.69 l=3.45
X1 VTAIL.t19 VP.t0 VDD1.t7 w_n5506_n4706# sky130_fd_pr__pfet_01v8 ad=3.08385 pd=19.02 as=3.08385 ps=19.02 w=18.69 l=3.45
X2 VDD1.t6 VP.t1 VTAIL.t18 w_n5506_n4706# sky130_fd_pr__pfet_01v8 ad=3.08385 pd=19.02 as=7.2891 ps=38.16 w=18.69 l=3.45
X3 VTAIL.t9 VN.t0 VDD2.t9 w_n5506_n4706# sky130_fd_pr__pfet_01v8 ad=3.08385 pd=19.02 as=3.08385 ps=19.02 w=18.69 l=3.45
X4 VDD2.t8 VN.t1 VTAIL.t8 w_n5506_n4706# sky130_fd_pr__pfet_01v8 ad=3.08385 pd=19.02 as=3.08385 ps=19.02 w=18.69 l=3.45
X5 VDD2.t7 VN.t2 VTAIL.t7 w_n5506_n4706# sky130_fd_pr__pfet_01v8 ad=3.08385 pd=19.02 as=3.08385 ps=19.02 w=18.69 l=3.45
X6 VTAIL.t17 VP.t2 VDD1.t9 w_n5506_n4706# sky130_fd_pr__pfet_01v8 ad=3.08385 pd=19.02 as=3.08385 ps=19.02 w=18.69 l=3.45
X7 VDD2.t6 VN.t3 VTAIL.t6 w_n5506_n4706# sky130_fd_pr__pfet_01v8 ad=7.2891 pd=38.16 as=3.08385 ps=19.02 w=18.69 l=3.45
X8 VDD1.t3 VP.t3 VTAIL.t16 w_n5506_n4706# sky130_fd_pr__pfet_01v8 ad=3.08385 pd=19.02 as=3.08385 ps=19.02 w=18.69 l=3.45
X9 B.t8 B.t6 B.t7 w_n5506_n4706# sky130_fd_pr__pfet_01v8 ad=7.2891 pd=38.16 as=0 ps=0 w=18.69 l=3.45
X10 B.t5 B.t3 B.t4 w_n5506_n4706# sky130_fd_pr__pfet_01v8 ad=7.2891 pd=38.16 as=0 ps=0 w=18.69 l=3.45
X11 VDD2.t5 VN.t4 VTAIL.t5 w_n5506_n4706# sky130_fd_pr__pfet_01v8 ad=3.08385 pd=19.02 as=7.2891 ps=38.16 w=18.69 l=3.45
X12 VTAIL.t4 VN.t5 VDD2.t4 w_n5506_n4706# sky130_fd_pr__pfet_01v8 ad=3.08385 pd=19.02 as=3.08385 ps=19.02 w=18.69 l=3.45
X13 B.t2 B.t0 B.t1 w_n5506_n4706# sky130_fd_pr__pfet_01v8 ad=7.2891 pd=38.16 as=0 ps=0 w=18.69 l=3.45
X14 VDD1.t8 VP.t4 VTAIL.t15 w_n5506_n4706# sky130_fd_pr__pfet_01v8 ad=7.2891 pd=38.16 as=3.08385 ps=19.02 w=18.69 l=3.45
X15 VDD2.t3 VN.t6 VTAIL.t3 w_n5506_n4706# sky130_fd_pr__pfet_01v8 ad=7.2891 pd=38.16 as=3.08385 ps=19.02 w=18.69 l=3.45
X16 VTAIL.t14 VP.t5 VDD1.t5 w_n5506_n4706# sky130_fd_pr__pfet_01v8 ad=3.08385 pd=19.02 as=3.08385 ps=19.02 w=18.69 l=3.45
X17 VDD1.t4 VP.t6 VTAIL.t13 w_n5506_n4706# sky130_fd_pr__pfet_01v8 ad=3.08385 pd=19.02 as=7.2891 ps=38.16 w=18.69 l=3.45
X18 VDD1.t1 VP.t7 VTAIL.t12 w_n5506_n4706# sky130_fd_pr__pfet_01v8 ad=3.08385 pd=19.02 as=3.08385 ps=19.02 w=18.69 l=3.45
X19 VTAIL.t2 VN.t7 VDD2.t2 w_n5506_n4706# sky130_fd_pr__pfet_01v8 ad=3.08385 pd=19.02 as=3.08385 ps=19.02 w=18.69 l=3.45
X20 VDD1.t2 VP.t8 VTAIL.t11 w_n5506_n4706# sky130_fd_pr__pfet_01v8 ad=7.2891 pd=38.16 as=3.08385 ps=19.02 w=18.69 l=3.45
X21 VTAIL.t1 VN.t8 VDD2.t1 w_n5506_n4706# sky130_fd_pr__pfet_01v8 ad=3.08385 pd=19.02 as=3.08385 ps=19.02 w=18.69 l=3.45
X22 VDD2.t0 VN.t9 VTAIL.t0 w_n5506_n4706# sky130_fd_pr__pfet_01v8 ad=3.08385 pd=19.02 as=7.2891 ps=38.16 w=18.69 l=3.45
X23 VTAIL.t10 VP.t9 VDD1.t0 w_n5506_n4706# sky130_fd_pr__pfet_01v8 ad=3.08385 pd=19.02 as=3.08385 ps=19.02 w=18.69 l=3.45
R0 B.n831 B.n830 585
R1 B.n832 B.n109 585
R2 B.n834 B.n833 585
R3 B.n835 B.n108 585
R4 B.n837 B.n836 585
R5 B.n838 B.n107 585
R6 B.n840 B.n839 585
R7 B.n841 B.n106 585
R8 B.n843 B.n842 585
R9 B.n844 B.n105 585
R10 B.n846 B.n845 585
R11 B.n847 B.n104 585
R12 B.n849 B.n848 585
R13 B.n850 B.n103 585
R14 B.n852 B.n851 585
R15 B.n853 B.n102 585
R16 B.n855 B.n854 585
R17 B.n856 B.n101 585
R18 B.n858 B.n857 585
R19 B.n859 B.n100 585
R20 B.n861 B.n860 585
R21 B.n862 B.n99 585
R22 B.n864 B.n863 585
R23 B.n865 B.n98 585
R24 B.n867 B.n866 585
R25 B.n868 B.n97 585
R26 B.n870 B.n869 585
R27 B.n871 B.n96 585
R28 B.n873 B.n872 585
R29 B.n874 B.n95 585
R30 B.n876 B.n875 585
R31 B.n877 B.n94 585
R32 B.n879 B.n878 585
R33 B.n880 B.n93 585
R34 B.n882 B.n881 585
R35 B.n883 B.n92 585
R36 B.n885 B.n884 585
R37 B.n886 B.n91 585
R38 B.n888 B.n887 585
R39 B.n889 B.n90 585
R40 B.n891 B.n890 585
R41 B.n892 B.n89 585
R42 B.n894 B.n893 585
R43 B.n895 B.n88 585
R44 B.n897 B.n896 585
R45 B.n898 B.n87 585
R46 B.n900 B.n899 585
R47 B.n901 B.n86 585
R48 B.n903 B.n902 585
R49 B.n904 B.n85 585
R50 B.n906 B.n905 585
R51 B.n907 B.n84 585
R52 B.n909 B.n908 585
R53 B.n910 B.n83 585
R54 B.n912 B.n911 585
R55 B.n913 B.n82 585
R56 B.n915 B.n914 585
R57 B.n916 B.n81 585
R58 B.n918 B.n917 585
R59 B.n919 B.n80 585
R60 B.n921 B.n920 585
R61 B.n923 B.n77 585
R62 B.n925 B.n924 585
R63 B.n926 B.n76 585
R64 B.n928 B.n927 585
R65 B.n929 B.n75 585
R66 B.n931 B.n930 585
R67 B.n932 B.n74 585
R68 B.n934 B.n933 585
R69 B.n935 B.n73 585
R70 B.n937 B.n936 585
R71 B.n939 B.n938 585
R72 B.n940 B.n69 585
R73 B.n942 B.n941 585
R74 B.n943 B.n68 585
R75 B.n945 B.n944 585
R76 B.n946 B.n67 585
R77 B.n948 B.n947 585
R78 B.n949 B.n66 585
R79 B.n951 B.n950 585
R80 B.n952 B.n65 585
R81 B.n954 B.n953 585
R82 B.n955 B.n64 585
R83 B.n957 B.n956 585
R84 B.n958 B.n63 585
R85 B.n960 B.n959 585
R86 B.n961 B.n62 585
R87 B.n963 B.n962 585
R88 B.n964 B.n61 585
R89 B.n966 B.n965 585
R90 B.n967 B.n60 585
R91 B.n969 B.n968 585
R92 B.n970 B.n59 585
R93 B.n972 B.n971 585
R94 B.n973 B.n58 585
R95 B.n975 B.n974 585
R96 B.n976 B.n57 585
R97 B.n978 B.n977 585
R98 B.n979 B.n56 585
R99 B.n981 B.n980 585
R100 B.n982 B.n55 585
R101 B.n984 B.n983 585
R102 B.n985 B.n54 585
R103 B.n987 B.n986 585
R104 B.n988 B.n53 585
R105 B.n990 B.n989 585
R106 B.n991 B.n52 585
R107 B.n993 B.n992 585
R108 B.n994 B.n51 585
R109 B.n996 B.n995 585
R110 B.n997 B.n50 585
R111 B.n999 B.n998 585
R112 B.n1000 B.n49 585
R113 B.n1002 B.n1001 585
R114 B.n1003 B.n48 585
R115 B.n1005 B.n1004 585
R116 B.n1006 B.n47 585
R117 B.n1008 B.n1007 585
R118 B.n1009 B.n46 585
R119 B.n1011 B.n1010 585
R120 B.n1012 B.n45 585
R121 B.n1014 B.n1013 585
R122 B.n1015 B.n44 585
R123 B.n1017 B.n1016 585
R124 B.n1018 B.n43 585
R125 B.n1020 B.n1019 585
R126 B.n1021 B.n42 585
R127 B.n1023 B.n1022 585
R128 B.n1024 B.n41 585
R129 B.n1026 B.n1025 585
R130 B.n1027 B.n40 585
R131 B.n1029 B.n1028 585
R132 B.n829 B.n110 585
R133 B.n828 B.n827 585
R134 B.n826 B.n111 585
R135 B.n825 B.n824 585
R136 B.n823 B.n112 585
R137 B.n822 B.n821 585
R138 B.n820 B.n113 585
R139 B.n819 B.n818 585
R140 B.n817 B.n114 585
R141 B.n816 B.n815 585
R142 B.n814 B.n115 585
R143 B.n813 B.n812 585
R144 B.n811 B.n116 585
R145 B.n810 B.n809 585
R146 B.n808 B.n117 585
R147 B.n807 B.n806 585
R148 B.n805 B.n118 585
R149 B.n804 B.n803 585
R150 B.n802 B.n119 585
R151 B.n801 B.n800 585
R152 B.n799 B.n120 585
R153 B.n798 B.n797 585
R154 B.n796 B.n121 585
R155 B.n795 B.n794 585
R156 B.n793 B.n122 585
R157 B.n792 B.n791 585
R158 B.n790 B.n123 585
R159 B.n789 B.n788 585
R160 B.n787 B.n124 585
R161 B.n786 B.n785 585
R162 B.n784 B.n125 585
R163 B.n783 B.n782 585
R164 B.n781 B.n126 585
R165 B.n780 B.n779 585
R166 B.n778 B.n127 585
R167 B.n777 B.n776 585
R168 B.n775 B.n128 585
R169 B.n774 B.n773 585
R170 B.n772 B.n129 585
R171 B.n771 B.n770 585
R172 B.n769 B.n130 585
R173 B.n768 B.n767 585
R174 B.n766 B.n131 585
R175 B.n765 B.n764 585
R176 B.n763 B.n132 585
R177 B.n762 B.n761 585
R178 B.n760 B.n133 585
R179 B.n759 B.n758 585
R180 B.n757 B.n134 585
R181 B.n756 B.n755 585
R182 B.n754 B.n135 585
R183 B.n753 B.n752 585
R184 B.n751 B.n136 585
R185 B.n750 B.n749 585
R186 B.n748 B.n137 585
R187 B.n747 B.n746 585
R188 B.n745 B.n138 585
R189 B.n744 B.n743 585
R190 B.n742 B.n139 585
R191 B.n741 B.n740 585
R192 B.n739 B.n140 585
R193 B.n738 B.n737 585
R194 B.n736 B.n141 585
R195 B.n735 B.n734 585
R196 B.n733 B.n142 585
R197 B.n732 B.n731 585
R198 B.n730 B.n143 585
R199 B.n729 B.n728 585
R200 B.n727 B.n144 585
R201 B.n726 B.n725 585
R202 B.n724 B.n145 585
R203 B.n723 B.n722 585
R204 B.n721 B.n146 585
R205 B.n720 B.n719 585
R206 B.n718 B.n147 585
R207 B.n717 B.n716 585
R208 B.n715 B.n148 585
R209 B.n714 B.n713 585
R210 B.n712 B.n149 585
R211 B.n711 B.n710 585
R212 B.n709 B.n150 585
R213 B.n708 B.n707 585
R214 B.n706 B.n151 585
R215 B.n705 B.n704 585
R216 B.n703 B.n152 585
R217 B.n702 B.n701 585
R218 B.n700 B.n153 585
R219 B.n699 B.n698 585
R220 B.n697 B.n154 585
R221 B.n696 B.n695 585
R222 B.n694 B.n155 585
R223 B.n693 B.n692 585
R224 B.n691 B.n156 585
R225 B.n690 B.n689 585
R226 B.n688 B.n157 585
R227 B.n687 B.n686 585
R228 B.n685 B.n158 585
R229 B.n684 B.n683 585
R230 B.n682 B.n159 585
R231 B.n681 B.n680 585
R232 B.n679 B.n160 585
R233 B.n678 B.n677 585
R234 B.n676 B.n161 585
R235 B.n675 B.n674 585
R236 B.n673 B.n162 585
R237 B.n672 B.n671 585
R238 B.n670 B.n163 585
R239 B.n669 B.n668 585
R240 B.n667 B.n164 585
R241 B.n666 B.n665 585
R242 B.n664 B.n165 585
R243 B.n663 B.n662 585
R244 B.n661 B.n166 585
R245 B.n660 B.n659 585
R246 B.n658 B.n167 585
R247 B.n657 B.n656 585
R248 B.n655 B.n168 585
R249 B.n654 B.n653 585
R250 B.n652 B.n169 585
R251 B.n651 B.n650 585
R252 B.n649 B.n170 585
R253 B.n648 B.n647 585
R254 B.n646 B.n171 585
R255 B.n645 B.n644 585
R256 B.n643 B.n172 585
R257 B.n642 B.n641 585
R258 B.n640 B.n173 585
R259 B.n639 B.n638 585
R260 B.n637 B.n174 585
R261 B.n636 B.n635 585
R262 B.n634 B.n175 585
R263 B.n633 B.n632 585
R264 B.n631 B.n176 585
R265 B.n630 B.n629 585
R266 B.n628 B.n177 585
R267 B.n627 B.n626 585
R268 B.n625 B.n178 585
R269 B.n624 B.n623 585
R270 B.n622 B.n179 585
R271 B.n621 B.n620 585
R272 B.n619 B.n180 585
R273 B.n618 B.n617 585
R274 B.n616 B.n181 585
R275 B.n615 B.n614 585
R276 B.n613 B.n182 585
R277 B.n612 B.n611 585
R278 B.n610 B.n183 585
R279 B.n609 B.n608 585
R280 B.n607 B.n184 585
R281 B.n606 B.n605 585
R282 B.n604 B.n185 585
R283 B.n405 B.n404 585
R284 B.n406 B.n255 585
R285 B.n408 B.n407 585
R286 B.n409 B.n254 585
R287 B.n411 B.n410 585
R288 B.n412 B.n253 585
R289 B.n414 B.n413 585
R290 B.n415 B.n252 585
R291 B.n417 B.n416 585
R292 B.n418 B.n251 585
R293 B.n420 B.n419 585
R294 B.n421 B.n250 585
R295 B.n423 B.n422 585
R296 B.n424 B.n249 585
R297 B.n426 B.n425 585
R298 B.n427 B.n248 585
R299 B.n429 B.n428 585
R300 B.n430 B.n247 585
R301 B.n432 B.n431 585
R302 B.n433 B.n246 585
R303 B.n435 B.n434 585
R304 B.n436 B.n245 585
R305 B.n438 B.n437 585
R306 B.n439 B.n244 585
R307 B.n441 B.n440 585
R308 B.n442 B.n243 585
R309 B.n444 B.n443 585
R310 B.n445 B.n242 585
R311 B.n447 B.n446 585
R312 B.n448 B.n241 585
R313 B.n450 B.n449 585
R314 B.n451 B.n240 585
R315 B.n453 B.n452 585
R316 B.n454 B.n239 585
R317 B.n456 B.n455 585
R318 B.n457 B.n238 585
R319 B.n459 B.n458 585
R320 B.n460 B.n237 585
R321 B.n462 B.n461 585
R322 B.n463 B.n236 585
R323 B.n465 B.n464 585
R324 B.n466 B.n235 585
R325 B.n468 B.n467 585
R326 B.n469 B.n234 585
R327 B.n471 B.n470 585
R328 B.n472 B.n233 585
R329 B.n474 B.n473 585
R330 B.n475 B.n232 585
R331 B.n477 B.n476 585
R332 B.n478 B.n231 585
R333 B.n480 B.n479 585
R334 B.n481 B.n230 585
R335 B.n483 B.n482 585
R336 B.n484 B.n229 585
R337 B.n486 B.n485 585
R338 B.n487 B.n228 585
R339 B.n489 B.n488 585
R340 B.n490 B.n227 585
R341 B.n492 B.n491 585
R342 B.n493 B.n226 585
R343 B.n495 B.n494 585
R344 B.n497 B.n223 585
R345 B.n499 B.n498 585
R346 B.n500 B.n222 585
R347 B.n502 B.n501 585
R348 B.n503 B.n221 585
R349 B.n505 B.n504 585
R350 B.n506 B.n220 585
R351 B.n508 B.n507 585
R352 B.n509 B.n219 585
R353 B.n511 B.n510 585
R354 B.n513 B.n512 585
R355 B.n514 B.n215 585
R356 B.n516 B.n515 585
R357 B.n517 B.n214 585
R358 B.n519 B.n518 585
R359 B.n520 B.n213 585
R360 B.n522 B.n521 585
R361 B.n523 B.n212 585
R362 B.n525 B.n524 585
R363 B.n526 B.n211 585
R364 B.n528 B.n527 585
R365 B.n529 B.n210 585
R366 B.n531 B.n530 585
R367 B.n532 B.n209 585
R368 B.n534 B.n533 585
R369 B.n535 B.n208 585
R370 B.n537 B.n536 585
R371 B.n538 B.n207 585
R372 B.n540 B.n539 585
R373 B.n541 B.n206 585
R374 B.n543 B.n542 585
R375 B.n544 B.n205 585
R376 B.n546 B.n545 585
R377 B.n547 B.n204 585
R378 B.n549 B.n548 585
R379 B.n550 B.n203 585
R380 B.n552 B.n551 585
R381 B.n553 B.n202 585
R382 B.n555 B.n554 585
R383 B.n556 B.n201 585
R384 B.n558 B.n557 585
R385 B.n559 B.n200 585
R386 B.n561 B.n560 585
R387 B.n562 B.n199 585
R388 B.n564 B.n563 585
R389 B.n565 B.n198 585
R390 B.n567 B.n566 585
R391 B.n568 B.n197 585
R392 B.n570 B.n569 585
R393 B.n571 B.n196 585
R394 B.n573 B.n572 585
R395 B.n574 B.n195 585
R396 B.n576 B.n575 585
R397 B.n577 B.n194 585
R398 B.n579 B.n578 585
R399 B.n580 B.n193 585
R400 B.n582 B.n581 585
R401 B.n583 B.n192 585
R402 B.n585 B.n584 585
R403 B.n586 B.n191 585
R404 B.n588 B.n587 585
R405 B.n589 B.n190 585
R406 B.n591 B.n590 585
R407 B.n592 B.n189 585
R408 B.n594 B.n593 585
R409 B.n595 B.n188 585
R410 B.n597 B.n596 585
R411 B.n598 B.n187 585
R412 B.n600 B.n599 585
R413 B.n601 B.n186 585
R414 B.n603 B.n602 585
R415 B.n403 B.n256 585
R416 B.n402 B.n401 585
R417 B.n400 B.n257 585
R418 B.n399 B.n398 585
R419 B.n397 B.n258 585
R420 B.n396 B.n395 585
R421 B.n394 B.n259 585
R422 B.n393 B.n392 585
R423 B.n391 B.n260 585
R424 B.n390 B.n389 585
R425 B.n388 B.n261 585
R426 B.n387 B.n386 585
R427 B.n385 B.n262 585
R428 B.n384 B.n383 585
R429 B.n382 B.n263 585
R430 B.n381 B.n380 585
R431 B.n379 B.n264 585
R432 B.n378 B.n377 585
R433 B.n376 B.n265 585
R434 B.n375 B.n374 585
R435 B.n373 B.n266 585
R436 B.n372 B.n371 585
R437 B.n370 B.n267 585
R438 B.n369 B.n368 585
R439 B.n367 B.n268 585
R440 B.n366 B.n365 585
R441 B.n364 B.n269 585
R442 B.n363 B.n362 585
R443 B.n361 B.n270 585
R444 B.n360 B.n359 585
R445 B.n358 B.n271 585
R446 B.n357 B.n356 585
R447 B.n355 B.n272 585
R448 B.n354 B.n353 585
R449 B.n352 B.n273 585
R450 B.n351 B.n350 585
R451 B.n349 B.n274 585
R452 B.n348 B.n347 585
R453 B.n346 B.n275 585
R454 B.n345 B.n344 585
R455 B.n343 B.n276 585
R456 B.n342 B.n341 585
R457 B.n340 B.n277 585
R458 B.n339 B.n338 585
R459 B.n337 B.n278 585
R460 B.n336 B.n335 585
R461 B.n334 B.n279 585
R462 B.n333 B.n332 585
R463 B.n331 B.n280 585
R464 B.n330 B.n329 585
R465 B.n328 B.n281 585
R466 B.n327 B.n326 585
R467 B.n325 B.n282 585
R468 B.n324 B.n323 585
R469 B.n322 B.n283 585
R470 B.n321 B.n320 585
R471 B.n319 B.n284 585
R472 B.n318 B.n317 585
R473 B.n316 B.n285 585
R474 B.n315 B.n314 585
R475 B.n313 B.n286 585
R476 B.n312 B.n311 585
R477 B.n310 B.n287 585
R478 B.n309 B.n308 585
R479 B.n307 B.n288 585
R480 B.n306 B.n305 585
R481 B.n304 B.n289 585
R482 B.n303 B.n302 585
R483 B.n301 B.n290 585
R484 B.n300 B.n299 585
R485 B.n298 B.n291 585
R486 B.n297 B.n296 585
R487 B.n295 B.n292 585
R488 B.n294 B.n293 585
R489 B.n2 B.n0 585
R490 B.n1141 B.n1 585
R491 B.n1140 B.n1139 585
R492 B.n1138 B.n3 585
R493 B.n1137 B.n1136 585
R494 B.n1135 B.n4 585
R495 B.n1134 B.n1133 585
R496 B.n1132 B.n5 585
R497 B.n1131 B.n1130 585
R498 B.n1129 B.n6 585
R499 B.n1128 B.n1127 585
R500 B.n1126 B.n7 585
R501 B.n1125 B.n1124 585
R502 B.n1123 B.n8 585
R503 B.n1122 B.n1121 585
R504 B.n1120 B.n9 585
R505 B.n1119 B.n1118 585
R506 B.n1117 B.n10 585
R507 B.n1116 B.n1115 585
R508 B.n1114 B.n11 585
R509 B.n1113 B.n1112 585
R510 B.n1111 B.n12 585
R511 B.n1110 B.n1109 585
R512 B.n1108 B.n13 585
R513 B.n1107 B.n1106 585
R514 B.n1105 B.n14 585
R515 B.n1104 B.n1103 585
R516 B.n1102 B.n15 585
R517 B.n1101 B.n1100 585
R518 B.n1099 B.n16 585
R519 B.n1098 B.n1097 585
R520 B.n1096 B.n17 585
R521 B.n1095 B.n1094 585
R522 B.n1093 B.n18 585
R523 B.n1092 B.n1091 585
R524 B.n1090 B.n19 585
R525 B.n1089 B.n1088 585
R526 B.n1087 B.n20 585
R527 B.n1086 B.n1085 585
R528 B.n1084 B.n21 585
R529 B.n1083 B.n1082 585
R530 B.n1081 B.n22 585
R531 B.n1080 B.n1079 585
R532 B.n1078 B.n23 585
R533 B.n1077 B.n1076 585
R534 B.n1075 B.n24 585
R535 B.n1074 B.n1073 585
R536 B.n1072 B.n25 585
R537 B.n1071 B.n1070 585
R538 B.n1069 B.n26 585
R539 B.n1068 B.n1067 585
R540 B.n1066 B.n27 585
R541 B.n1065 B.n1064 585
R542 B.n1063 B.n28 585
R543 B.n1062 B.n1061 585
R544 B.n1060 B.n29 585
R545 B.n1059 B.n1058 585
R546 B.n1057 B.n30 585
R547 B.n1056 B.n1055 585
R548 B.n1054 B.n31 585
R549 B.n1053 B.n1052 585
R550 B.n1051 B.n32 585
R551 B.n1050 B.n1049 585
R552 B.n1048 B.n33 585
R553 B.n1047 B.n1046 585
R554 B.n1045 B.n34 585
R555 B.n1044 B.n1043 585
R556 B.n1042 B.n35 585
R557 B.n1041 B.n1040 585
R558 B.n1039 B.n36 585
R559 B.n1038 B.n1037 585
R560 B.n1036 B.n37 585
R561 B.n1035 B.n1034 585
R562 B.n1033 B.n38 585
R563 B.n1032 B.n1031 585
R564 B.n1030 B.n39 585
R565 B.n1143 B.n1142 585
R566 B.n404 B.n403 482.89
R567 B.n1028 B.n39 482.89
R568 B.n602 B.n185 482.89
R569 B.n830 B.n829 482.89
R570 B.n216 B.t9 339.608
R571 B.n224 B.t0 339.608
R572 B.n70 B.t6 339.608
R573 B.n78 B.t3 339.608
R574 B.n216 B.t11 185.847
R575 B.n78 B.t4 185.847
R576 B.n224 B.t2 185.823
R577 B.n70 B.t7 185.823
R578 B.n403 B.n402 163.367
R579 B.n402 B.n257 163.367
R580 B.n398 B.n257 163.367
R581 B.n398 B.n397 163.367
R582 B.n397 B.n396 163.367
R583 B.n396 B.n259 163.367
R584 B.n392 B.n259 163.367
R585 B.n392 B.n391 163.367
R586 B.n391 B.n390 163.367
R587 B.n390 B.n261 163.367
R588 B.n386 B.n261 163.367
R589 B.n386 B.n385 163.367
R590 B.n385 B.n384 163.367
R591 B.n384 B.n263 163.367
R592 B.n380 B.n263 163.367
R593 B.n380 B.n379 163.367
R594 B.n379 B.n378 163.367
R595 B.n378 B.n265 163.367
R596 B.n374 B.n265 163.367
R597 B.n374 B.n373 163.367
R598 B.n373 B.n372 163.367
R599 B.n372 B.n267 163.367
R600 B.n368 B.n267 163.367
R601 B.n368 B.n367 163.367
R602 B.n367 B.n366 163.367
R603 B.n366 B.n269 163.367
R604 B.n362 B.n269 163.367
R605 B.n362 B.n361 163.367
R606 B.n361 B.n360 163.367
R607 B.n360 B.n271 163.367
R608 B.n356 B.n271 163.367
R609 B.n356 B.n355 163.367
R610 B.n355 B.n354 163.367
R611 B.n354 B.n273 163.367
R612 B.n350 B.n273 163.367
R613 B.n350 B.n349 163.367
R614 B.n349 B.n348 163.367
R615 B.n348 B.n275 163.367
R616 B.n344 B.n275 163.367
R617 B.n344 B.n343 163.367
R618 B.n343 B.n342 163.367
R619 B.n342 B.n277 163.367
R620 B.n338 B.n277 163.367
R621 B.n338 B.n337 163.367
R622 B.n337 B.n336 163.367
R623 B.n336 B.n279 163.367
R624 B.n332 B.n279 163.367
R625 B.n332 B.n331 163.367
R626 B.n331 B.n330 163.367
R627 B.n330 B.n281 163.367
R628 B.n326 B.n281 163.367
R629 B.n326 B.n325 163.367
R630 B.n325 B.n324 163.367
R631 B.n324 B.n283 163.367
R632 B.n320 B.n283 163.367
R633 B.n320 B.n319 163.367
R634 B.n319 B.n318 163.367
R635 B.n318 B.n285 163.367
R636 B.n314 B.n285 163.367
R637 B.n314 B.n313 163.367
R638 B.n313 B.n312 163.367
R639 B.n312 B.n287 163.367
R640 B.n308 B.n287 163.367
R641 B.n308 B.n307 163.367
R642 B.n307 B.n306 163.367
R643 B.n306 B.n289 163.367
R644 B.n302 B.n289 163.367
R645 B.n302 B.n301 163.367
R646 B.n301 B.n300 163.367
R647 B.n300 B.n291 163.367
R648 B.n296 B.n291 163.367
R649 B.n296 B.n295 163.367
R650 B.n295 B.n294 163.367
R651 B.n294 B.n2 163.367
R652 B.n1142 B.n2 163.367
R653 B.n1142 B.n1141 163.367
R654 B.n1141 B.n1140 163.367
R655 B.n1140 B.n3 163.367
R656 B.n1136 B.n3 163.367
R657 B.n1136 B.n1135 163.367
R658 B.n1135 B.n1134 163.367
R659 B.n1134 B.n5 163.367
R660 B.n1130 B.n5 163.367
R661 B.n1130 B.n1129 163.367
R662 B.n1129 B.n1128 163.367
R663 B.n1128 B.n7 163.367
R664 B.n1124 B.n7 163.367
R665 B.n1124 B.n1123 163.367
R666 B.n1123 B.n1122 163.367
R667 B.n1122 B.n9 163.367
R668 B.n1118 B.n9 163.367
R669 B.n1118 B.n1117 163.367
R670 B.n1117 B.n1116 163.367
R671 B.n1116 B.n11 163.367
R672 B.n1112 B.n11 163.367
R673 B.n1112 B.n1111 163.367
R674 B.n1111 B.n1110 163.367
R675 B.n1110 B.n13 163.367
R676 B.n1106 B.n13 163.367
R677 B.n1106 B.n1105 163.367
R678 B.n1105 B.n1104 163.367
R679 B.n1104 B.n15 163.367
R680 B.n1100 B.n15 163.367
R681 B.n1100 B.n1099 163.367
R682 B.n1099 B.n1098 163.367
R683 B.n1098 B.n17 163.367
R684 B.n1094 B.n17 163.367
R685 B.n1094 B.n1093 163.367
R686 B.n1093 B.n1092 163.367
R687 B.n1092 B.n19 163.367
R688 B.n1088 B.n19 163.367
R689 B.n1088 B.n1087 163.367
R690 B.n1087 B.n1086 163.367
R691 B.n1086 B.n21 163.367
R692 B.n1082 B.n21 163.367
R693 B.n1082 B.n1081 163.367
R694 B.n1081 B.n1080 163.367
R695 B.n1080 B.n23 163.367
R696 B.n1076 B.n23 163.367
R697 B.n1076 B.n1075 163.367
R698 B.n1075 B.n1074 163.367
R699 B.n1074 B.n25 163.367
R700 B.n1070 B.n25 163.367
R701 B.n1070 B.n1069 163.367
R702 B.n1069 B.n1068 163.367
R703 B.n1068 B.n27 163.367
R704 B.n1064 B.n27 163.367
R705 B.n1064 B.n1063 163.367
R706 B.n1063 B.n1062 163.367
R707 B.n1062 B.n29 163.367
R708 B.n1058 B.n29 163.367
R709 B.n1058 B.n1057 163.367
R710 B.n1057 B.n1056 163.367
R711 B.n1056 B.n31 163.367
R712 B.n1052 B.n31 163.367
R713 B.n1052 B.n1051 163.367
R714 B.n1051 B.n1050 163.367
R715 B.n1050 B.n33 163.367
R716 B.n1046 B.n33 163.367
R717 B.n1046 B.n1045 163.367
R718 B.n1045 B.n1044 163.367
R719 B.n1044 B.n35 163.367
R720 B.n1040 B.n35 163.367
R721 B.n1040 B.n1039 163.367
R722 B.n1039 B.n1038 163.367
R723 B.n1038 B.n37 163.367
R724 B.n1034 B.n37 163.367
R725 B.n1034 B.n1033 163.367
R726 B.n1033 B.n1032 163.367
R727 B.n1032 B.n39 163.367
R728 B.n404 B.n255 163.367
R729 B.n408 B.n255 163.367
R730 B.n409 B.n408 163.367
R731 B.n410 B.n409 163.367
R732 B.n410 B.n253 163.367
R733 B.n414 B.n253 163.367
R734 B.n415 B.n414 163.367
R735 B.n416 B.n415 163.367
R736 B.n416 B.n251 163.367
R737 B.n420 B.n251 163.367
R738 B.n421 B.n420 163.367
R739 B.n422 B.n421 163.367
R740 B.n422 B.n249 163.367
R741 B.n426 B.n249 163.367
R742 B.n427 B.n426 163.367
R743 B.n428 B.n427 163.367
R744 B.n428 B.n247 163.367
R745 B.n432 B.n247 163.367
R746 B.n433 B.n432 163.367
R747 B.n434 B.n433 163.367
R748 B.n434 B.n245 163.367
R749 B.n438 B.n245 163.367
R750 B.n439 B.n438 163.367
R751 B.n440 B.n439 163.367
R752 B.n440 B.n243 163.367
R753 B.n444 B.n243 163.367
R754 B.n445 B.n444 163.367
R755 B.n446 B.n445 163.367
R756 B.n446 B.n241 163.367
R757 B.n450 B.n241 163.367
R758 B.n451 B.n450 163.367
R759 B.n452 B.n451 163.367
R760 B.n452 B.n239 163.367
R761 B.n456 B.n239 163.367
R762 B.n457 B.n456 163.367
R763 B.n458 B.n457 163.367
R764 B.n458 B.n237 163.367
R765 B.n462 B.n237 163.367
R766 B.n463 B.n462 163.367
R767 B.n464 B.n463 163.367
R768 B.n464 B.n235 163.367
R769 B.n468 B.n235 163.367
R770 B.n469 B.n468 163.367
R771 B.n470 B.n469 163.367
R772 B.n470 B.n233 163.367
R773 B.n474 B.n233 163.367
R774 B.n475 B.n474 163.367
R775 B.n476 B.n475 163.367
R776 B.n476 B.n231 163.367
R777 B.n480 B.n231 163.367
R778 B.n481 B.n480 163.367
R779 B.n482 B.n481 163.367
R780 B.n482 B.n229 163.367
R781 B.n486 B.n229 163.367
R782 B.n487 B.n486 163.367
R783 B.n488 B.n487 163.367
R784 B.n488 B.n227 163.367
R785 B.n492 B.n227 163.367
R786 B.n493 B.n492 163.367
R787 B.n494 B.n493 163.367
R788 B.n494 B.n223 163.367
R789 B.n499 B.n223 163.367
R790 B.n500 B.n499 163.367
R791 B.n501 B.n500 163.367
R792 B.n501 B.n221 163.367
R793 B.n505 B.n221 163.367
R794 B.n506 B.n505 163.367
R795 B.n507 B.n506 163.367
R796 B.n507 B.n219 163.367
R797 B.n511 B.n219 163.367
R798 B.n512 B.n511 163.367
R799 B.n512 B.n215 163.367
R800 B.n516 B.n215 163.367
R801 B.n517 B.n516 163.367
R802 B.n518 B.n517 163.367
R803 B.n518 B.n213 163.367
R804 B.n522 B.n213 163.367
R805 B.n523 B.n522 163.367
R806 B.n524 B.n523 163.367
R807 B.n524 B.n211 163.367
R808 B.n528 B.n211 163.367
R809 B.n529 B.n528 163.367
R810 B.n530 B.n529 163.367
R811 B.n530 B.n209 163.367
R812 B.n534 B.n209 163.367
R813 B.n535 B.n534 163.367
R814 B.n536 B.n535 163.367
R815 B.n536 B.n207 163.367
R816 B.n540 B.n207 163.367
R817 B.n541 B.n540 163.367
R818 B.n542 B.n541 163.367
R819 B.n542 B.n205 163.367
R820 B.n546 B.n205 163.367
R821 B.n547 B.n546 163.367
R822 B.n548 B.n547 163.367
R823 B.n548 B.n203 163.367
R824 B.n552 B.n203 163.367
R825 B.n553 B.n552 163.367
R826 B.n554 B.n553 163.367
R827 B.n554 B.n201 163.367
R828 B.n558 B.n201 163.367
R829 B.n559 B.n558 163.367
R830 B.n560 B.n559 163.367
R831 B.n560 B.n199 163.367
R832 B.n564 B.n199 163.367
R833 B.n565 B.n564 163.367
R834 B.n566 B.n565 163.367
R835 B.n566 B.n197 163.367
R836 B.n570 B.n197 163.367
R837 B.n571 B.n570 163.367
R838 B.n572 B.n571 163.367
R839 B.n572 B.n195 163.367
R840 B.n576 B.n195 163.367
R841 B.n577 B.n576 163.367
R842 B.n578 B.n577 163.367
R843 B.n578 B.n193 163.367
R844 B.n582 B.n193 163.367
R845 B.n583 B.n582 163.367
R846 B.n584 B.n583 163.367
R847 B.n584 B.n191 163.367
R848 B.n588 B.n191 163.367
R849 B.n589 B.n588 163.367
R850 B.n590 B.n589 163.367
R851 B.n590 B.n189 163.367
R852 B.n594 B.n189 163.367
R853 B.n595 B.n594 163.367
R854 B.n596 B.n595 163.367
R855 B.n596 B.n187 163.367
R856 B.n600 B.n187 163.367
R857 B.n601 B.n600 163.367
R858 B.n602 B.n601 163.367
R859 B.n606 B.n185 163.367
R860 B.n607 B.n606 163.367
R861 B.n608 B.n607 163.367
R862 B.n608 B.n183 163.367
R863 B.n612 B.n183 163.367
R864 B.n613 B.n612 163.367
R865 B.n614 B.n613 163.367
R866 B.n614 B.n181 163.367
R867 B.n618 B.n181 163.367
R868 B.n619 B.n618 163.367
R869 B.n620 B.n619 163.367
R870 B.n620 B.n179 163.367
R871 B.n624 B.n179 163.367
R872 B.n625 B.n624 163.367
R873 B.n626 B.n625 163.367
R874 B.n626 B.n177 163.367
R875 B.n630 B.n177 163.367
R876 B.n631 B.n630 163.367
R877 B.n632 B.n631 163.367
R878 B.n632 B.n175 163.367
R879 B.n636 B.n175 163.367
R880 B.n637 B.n636 163.367
R881 B.n638 B.n637 163.367
R882 B.n638 B.n173 163.367
R883 B.n642 B.n173 163.367
R884 B.n643 B.n642 163.367
R885 B.n644 B.n643 163.367
R886 B.n644 B.n171 163.367
R887 B.n648 B.n171 163.367
R888 B.n649 B.n648 163.367
R889 B.n650 B.n649 163.367
R890 B.n650 B.n169 163.367
R891 B.n654 B.n169 163.367
R892 B.n655 B.n654 163.367
R893 B.n656 B.n655 163.367
R894 B.n656 B.n167 163.367
R895 B.n660 B.n167 163.367
R896 B.n661 B.n660 163.367
R897 B.n662 B.n661 163.367
R898 B.n662 B.n165 163.367
R899 B.n666 B.n165 163.367
R900 B.n667 B.n666 163.367
R901 B.n668 B.n667 163.367
R902 B.n668 B.n163 163.367
R903 B.n672 B.n163 163.367
R904 B.n673 B.n672 163.367
R905 B.n674 B.n673 163.367
R906 B.n674 B.n161 163.367
R907 B.n678 B.n161 163.367
R908 B.n679 B.n678 163.367
R909 B.n680 B.n679 163.367
R910 B.n680 B.n159 163.367
R911 B.n684 B.n159 163.367
R912 B.n685 B.n684 163.367
R913 B.n686 B.n685 163.367
R914 B.n686 B.n157 163.367
R915 B.n690 B.n157 163.367
R916 B.n691 B.n690 163.367
R917 B.n692 B.n691 163.367
R918 B.n692 B.n155 163.367
R919 B.n696 B.n155 163.367
R920 B.n697 B.n696 163.367
R921 B.n698 B.n697 163.367
R922 B.n698 B.n153 163.367
R923 B.n702 B.n153 163.367
R924 B.n703 B.n702 163.367
R925 B.n704 B.n703 163.367
R926 B.n704 B.n151 163.367
R927 B.n708 B.n151 163.367
R928 B.n709 B.n708 163.367
R929 B.n710 B.n709 163.367
R930 B.n710 B.n149 163.367
R931 B.n714 B.n149 163.367
R932 B.n715 B.n714 163.367
R933 B.n716 B.n715 163.367
R934 B.n716 B.n147 163.367
R935 B.n720 B.n147 163.367
R936 B.n721 B.n720 163.367
R937 B.n722 B.n721 163.367
R938 B.n722 B.n145 163.367
R939 B.n726 B.n145 163.367
R940 B.n727 B.n726 163.367
R941 B.n728 B.n727 163.367
R942 B.n728 B.n143 163.367
R943 B.n732 B.n143 163.367
R944 B.n733 B.n732 163.367
R945 B.n734 B.n733 163.367
R946 B.n734 B.n141 163.367
R947 B.n738 B.n141 163.367
R948 B.n739 B.n738 163.367
R949 B.n740 B.n739 163.367
R950 B.n740 B.n139 163.367
R951 B.n744 B.n139 163.367
R952 B.n745 B.n744 163.367
R953 B.n746 B.n745 163.367
R954 B.n746 B.n137 163.367
R955 B.n750 B.n137 163.367
R956 B.n751 B.n750 163.367
R957 B.n752 B.n751 163.367
R958 B.n752 B.n135 163.367
R959 B.n756 B.n135 163.367
R960 B.n757 B.n756 163.367
R961 B.n758 B.n757 163.367
R962 B.n758 B.n133 163.367
R963 B.n762 B.n133 163.367
R964 B.n763 B.n762 163.367
R965 B.n764 B.n763 163.367
R966 B.n764 B.n131 163.367
R967 B.n768 B.n131 163.367
R968 B.n769 B.n768 163.367
R969 B.n770 B.n769 163.367
R970 B.n770 B.n129 163.367
R971 B.n774 B.n129 163.367
R972 B.n775 B.n774 163.367
R973 B.n776 B.n775 163.367
R974 B.n776 B.n127 163.367
R975 B.n780 B.n127 163.367
R976 B.n781 B.n780 163.367
R977 B.n782 B.n781 163.367
R978 B.n782 B.n125 163.367
R979 B.n786 B.n125 163.367
R980 B.n787 B.n786 163.367
R981 B.n788 B.n787 163.367
R982 B.n788 B.n123 163.367
R983 B.n792 B.n123 163.367
R984 B.n793 B.n792 163.367
R985 B.n794 B.n793 163.367
R986 B.n794 B.n121 163.367
R987 B.n798 B.n121 163.367
R988 B.n799 B.n798 163.367
R989 B.n800 B.n799 163.367
R990 B.n800 B.n119 163.367
R991 B.n804 B.n119 163.367
R992 B.n805 B.n804 163.367
R993 B.n806 B.n805 163.367
R994 B.n806 B.n117 163.367
R995 B.n810 B.n117 163.367
R996 B.n811 B.n810 163.367
R997 B.n812 B.n811 163.367
R998 B.n812 B.n115 163.367
R999 B.n816 B.n115 163.367
R1000 B.n817 B.n816 163.367
R1001 B.n818 B.n817 163.367
R1002 B.n818 B.n113 163.367
R1003 B.n822 B.n113 163.367
R1004 B.n823 B.n822 163.367
R1005 B.n824 B.n823 163.367
R1006 B.n824 B.n111 163.367
R1007 B.n828 B.n111 163.367
R1008 B.n829 B.n828 163.367
R1009 B.n1028 B.n1027 163.367
R1010 B.n1027 B.n1026 163.367
R1011 B.n1026 B.n41 163.367
R1012 B.n1022 B.n41 163.367
R1013 B.n1022 B.n1021 163.367
R1014 B.n1021 B.n1020 163.367
R1015 B.n1020 B.n43 163.367
R1016 B.n1016 B.n43 163.367
R1017 B.n1016 B.n1015 163.367
R1018 B.n1015 B.n1014 163.367
R1019 B.n1014 B.n45 163.367
R1020 B.n1010 B.n45 163.367
R1021 B.n1010 B.n1009 163.367
R1022 B.n1009 B.n1008 163.367
R1023 B.n1008 B.n47 163.367
R1024 B.n1004 B.n47 163.367
R1025 B.n1004 B.n1003 163.367
R1026 B.n1003 B.n1002 163.367
R1027 B.n1002 B.n49 163.367
R1028 B.n998 B.n49 163.367
R1029 B.n998 B.n997 163.367
R1030 B.n997 B.n996 163.367
R1031 B.n996 B.n51 163.367
R1032 B.n992 B.n51 163.367
R1033 B.n992 B.n991 163.367
R1034 B.n991 B.n990 163.367
R1035 B.n990 B.n53 163.367
R1036 B.n986 B.n53 163.367
R1037 B.n986 B.n985 163.367
R1038 B.n985 B.n984 163.367
R1039 B.n984 B.n55 163.367
R1040 B.n980 B.n55 163.367
R1041 B.n980 B.n979 163.367
R1042 B.n979 B.n978 163.367
R1043 B.n978 B.n57 163.367
R1044 B.n974 B.n57 163.367
R1045 B.n974 B.n973 163.367
R1046 B.n973 B.n972 163.367
R1047 B.n972 B.n59 163.367
R1048 B.n968 B.n59 163.367
R1049 B.n968 B.n967 163.367
R1050 B.n967 B.n966 163.367
R1051 B.n966 B.n61 163.367
R1052 B.n962 B.n61 163.367
R1053 B.n962 B.n961 163.367
R1054 B.n961 B.n960 163.367
R1055 B.n960 B.n63 163.367
R1056 B.n956 B.n63 163.367
R1057 B.n956 B.n955 163.367
R1058 B.n955 B.n954 163.367
R1059 B.n954 B.n65 163.367
R1060 B.n950 B.n65 163.367
R1061 B.n950 B.n949 163.367
R1062 B.n949 B.n948 163.367
R1063 B.n948 B.n67 163.367
R1064 B.n944 B.n67 163.367
R1065 B.n944 B.n943 163.367
R1066 B.n943 B.n942 163.367
R1067 B.n942 B.n69 163.367
R1068 B.n938 B.n69 163.367
R1069 B.n938 B.n937 163.367
R1070 B.n937 B.n73 163.367
R1071 B.n933 B.n73 163.367
R1072 B.n933 B.n932 163.367
R1073 B.n932 B.n931 163.367
R1074 B.n931 B.n75 163.367
R1075 B.n927 B.n75 163.367
R1076 B.n927 B.n926 163.367
R1077 B.n926 B.n925 163.367
R1078 B.n925 B.n77 163.367
R1079 B.n920 B.n77 163.367
R1080 B.n920 B.n919 163.367
R1081 B.n919 B.n918 163.367
R1082 B.n918 B.n81 163.367
R1083 B.n914 B.n81 163.367
R1084 B.n914 B.n913 163.367
R1085 B.n913 B.n912 163.367
R1086 B.n912 B.n83 163.367
R1087 B.n908 B.n83 163.367
R1088 B.n908 B.n907 163.367
R1089 B.n907 B.n906 163.367
R1090 B.n906 B.n85 163.367
R1091 B.n902 B.n85 163.367
R1092 B.n902 B.n901 163.367
R1093 B.n901 B.n900 163.367
R1094 B.n900 B.n87 163.367
R1095 B.n896 B.n87 163.367
R1096 B.n896 B.n895 163.367
R1097 B.n895 B.n894 163.367
R1098 B.n894 B.n89 163.367
R1099 B.n890 B.n89 163.367
R1100 B.n890 B.n889 163.367
R1101 B.n889 B.n888 163.367
R1102 B.n888 B.n91 163.367
R1103 B.n884 B.n91 163.367
R1104 B.n884 B.n883 163.367
R1105 B.n883 B.n882 163.367
R1106 B.n882 B.n93 163.367
R1107 B.n878 B.n93 163.367
R1108 B.n878 B.n877 163.367
R1109 B.n877 B.n876 163.367
R1110 B.n876 B.n95 163.367
R1111 B.n872 B.n95 163.367
R1112 B.n872 B.n871 163.367
R1113 B.n871 B.n870 163.367
R1114 B.n870 B.n97 163.367
R1115 B.n866 B.n97 163.367
R1116 B.n866 B.n865 163.367
R1117 B.n865 B.n864 163.367
R1118 B.n864 B.n99 163.367
R1119 B.n860 B.n99 163.367
R1120 B.n860 B.n859 163.367
R1121 B.n859 B.n858 163.367
R1122 B.n858 B.n101 163.367
R1123 B.n854 B.n101 163.367
R1124 B.n854 B.n853 163.367
R1125 B.n853 B.n852 163.367
R1126 B.n852 B.n103 163.367
R1127 B.n848 B.n103 163.367
R1128 B.n848 B.n847 163.367
R1129 B.n847 B.n846 163.367
R1130 B.n846 B.n105 163.367
R1131 B.n842 B.n105 163.367
R1132 B.n842 B.n841 163.367
R1133 B.n841 B.n840 163.367
R1134 B.n840 B.n107 163.367
R1135 B.n836 B.n107 163.367
R1136 B.n836 B.n835 163.367
R1137 B.n835 B.n834 163.367
R1138 B.n834 B.n109 163.367
R1139 B.n830 B.n109 163.367
R1140 B.n217 B.t10 112.538
R1141 B.n79 B.t5 112.538
R1142 B.n225 B.t1 112.514
R1143 B.n71 B.t8 112.514
R1144 B.n217 B.n216 73.3096
R1145 B.n225 B.n224 73.3096
R1146 B.n71 B.n70 73.3096
R1147 B.n79 B.n78 73.3096
R1148 B.n218 B.n217 59.5399
R1149 B.n496 B.n225 59.5399
R1150 B.n72 B.n71 59.5399
R1151 B.n922 B.n79 59.5399
R1152 B.n1030 B.n1029 31.3761
R1153 B.n831 B.n110 31.3761
R1154 B.n604 B.n603 31.3761
R1155 B.n405 B.n256 31.3761
R1156 B B.n1143 18.0485
R1157 B.n1029 B.n40 10.6151
R1158 B.n1025 B.n40 10.6151
R1159 B.n1025 B.n1024 10.6151
R1160 B.n1024 B.n1023 10.6151
R1161 B.n1023 B.n42 10.6151
R1162 B.n1019 B.n42 10.6151
R1163 B.n1019 B.n1018 10.6151
R1164 B.n1018 B.n1017 10.6151
R1165 B.n1017 B.n44 10.6151
R1166 B.n1013 B.n44 10.6151
R1167 B.n1013 B.n1012 10.6151
R1168 B.n1012 B.n1011 10.6151
R1169 B.n1011 B.n46 10.6151
R1170 B.n1007 B.n46 10.6151
R1171 B.n1007 B.n1006 10.6151
R1172 B.n1006 B.n1005 10.6151
R1173 B.n1005 B.n48 10.6151
R1174 B.n1001 B.n48 10.6151
R1175 B.n1001 B.n1000 10.6151
R1176 B.n1000 B.n999 10.6151
R1177 B.n999 B.n50 10.6151
R1178 B.n995 B.n50 10.6151
R1179 B.n995 B.n994 10.6151
R1180 B.n994 B.n993 10.6151
R1181 B.n993 B.n52 10.6151
R1182 B.n989 B.n52 10.6151
R1183 B.n989 B.n988 10.6151
R1184 B.n988 B.n987 10.6151
R1185 B.n987 B.n54 10.6151
R1186 B.n983 B.n54 10.6151
R1187 B.n983 B.n982 10.6151
R1188 B.n982 B.n981 10.6151
R1189 B.n981 B.n56 10.6151
R1190 B.n977 B.n56 10.6151
R1191 B.n977 B.n976 10.6151
R1192 B.n976 B.n975 10.6151
R1193 B.n975 B.n58 10.6151
R1194 B.n971 B.n58 10.6151
R1195 B.n971 B.n970 10.6151
R1196 B.n970 B.n969 10.6151
R1197 B.n969 B.n60 10.6151
R1198 B.n965 B.n60 10.6151
R1199 B.n965 B.n964 10.6151
R1200 B.n964 B.n963 10.6151
R1201 B.n963 B.n62 10.6151
R1202 B.n959 B.n62 10.6151
R1203 B.n959 B.n958 10.6151
R1204 B.n958 B.n957 10.6151
R1205 B.n957 B.n64 10.6151
R1206 B.n953 B.n64 10.6151
R1207 B.n953 B.n952 10.6151
R1208 B.n952 B.n951 10.6151
R1209 B.n951 B.n66 10.6151
R1210 B.n947 B.n66 10.6151
R1211 B.n947 B.n946 10.6151
R1212 B.n946 B.n945 10.6151
R1213 B.n945 B.n68 10.6151
R1214 B.n941 B.n68 10.6151
R1215 B.n941 B.n940 10.6151
R1216 B.n940 B.n939 10.6151
R1217 B.n936 B.n935 10.6151
R1218 B.n935 B.n934 10.6151
R1219 B.n934 B.n74 10.6151
R1220 B.n930 B.n74 10.6151
R1221 B.n930 B.n929 10.6151
R1222 B.n929 B.n928 10.6151
R1223 B.n928 B.n76 10.6151
R1224 B.n924 B.n76 10.6151
R1225 B.n924 B.n923 10.6151
R1226 B.n921 B.n80 10.6151
R1227 B.n917 B.n80 10.6151
R1228 B.n917 B.n916 10.6151
R1229 B.n916 B.n915 10.6151
R1230 B.n915 B.n82 10.6151
R1231 B.n911 B.n82 10.6151
R1232 B.n911 B.n910 10.6151
R1233 B.n910 B.n909 10.6151
R1234 B.n909 B.n84 10.6151
R1235 B.n905 B.n84 10.6151
R1236 B.n905 B.n904 10.6151
R1237 B.n904 B.n903 10.6151
R1238 B.n903 B.n86 10.6151
R1239 B.n899 B.n86 10.6151
R1240 B.n899 B.n898 10.6151
R1241 B.n898 B.n897 10.6151
R1242 B.n897 B.n88 10.6151
R1243 B.n893 B.n88 10.6151
R1244 B.n893 B.n892 10.6151
R1245 B.n892 B.n891 10.6151
R1246 B.n891 B.n90 10.6151
R1247 B.n887 B.n90 10.6151
R1248 B.n887 B.n886 10.6151
R1249 B.n886 B.n885 10.6151
R1250 B.n885 B.n92 10.6151
R1251 B.n881 B.n92 10.6151
R1252 B.n881 B.n880 10.6151
R1253 B.n880 B.n879 10.6151
R1254 B.n879 B.n94 10.6151
R1255 B.n875 B.n94 10.6151
R1256 B.n875 B.n874 10.6151
R1257 B.n874 B.n873 10.6151
R1258 B.n873 B.n96 10.6151
R1259 B.n869 B.n96 10.6151
R1260 B.n869 B.n868 10.6151
R1261 B.n868 B.n867 10.6151
R1262 B.n867 B.n98 10.6151
R1263 B.n863 B.n98 10.6151
R1264 B.n863 B.n862 10.6151
R1265 B.n862 B.n861 10.6151
R1266 B.n861 B.n100 10.6151
R1267 B.n857 B.n100 10.6151
R1268 B.n857 B.n856 10.6151
R1269 B.n856 B.n855 10.6151
R1270 B.n855 B.n102 10.6151
R1271 B.n851 B.n102 10.6151
R1272 B.n851 B.n850 10.6151
R1273 B.n850 B.n849 10.6151
R1274 B.n849 B.n104 10.6151
R1275 B.n845 B.n104 10.6151
R1276 B.n845 B.n844 10.6151
R1277 B.n844 B.n843 10.6151
R1278 B.n843 B.n106 10.6151
R1279 B.n839 B.n106 10.6151
R1280 B.n839 B.n838 10.6151
R1281 B.n838 B.n837 10.6151
R1282 B.n837 B.n108 10.6151
R1283 B.n833 B.n108 10.6151
R1284 B.n833 B.n832 10.6151
R1285 B.n832 B.n831 10.6151
R1286 B.n605 B.n604 10.6151
R1287 B.n605 B.n184 10.6151
R1288 B.n609 B.n184 10.6151
R1289 B.n610 B.n609 10.6151
R1290 B.n611 B.n610 10.6151
R1291 B.n611 B.n182 10.6151
R1292 B.n615 B.n182 10.6151
R1293 B.n616 B.n615 10.6151
R1294 B.n617 B.n616 10.6151
R1295 B.n617 B.n180 10.6151
R1296 B.n621 B.n180 10.6151
R1297 B.n622 B.n621 10.6151
R1298 B.n623 B.n622 10.6151
R1299 B.n623 B.n178 10.6151
R1300 B.n627 B.n178 10.6151
R1301 B.n628 B.n627 10.6151
R1302 B.n629 B.n628 10.6151
R1303 B.n629 B.n176 10.6151
R1304 B.n633 B.n176 10.6151
R1305 B.n634 B.n633 10.6151
R1306 B.n635 B.n634 10.6151
R1307 B.n635 B.n174 10.6151
R1308 B.n639 B.n174 10.6151
R1309 B.n640 B.n639 10.6151
R1310 B.n641 B.n640 10.6151
R1311 B.n641 B.n172 10.6151
R1312 B.n645 B.n172 10.6151
R1313 B.n646 B.n645 10.6151
R1314 B.n647 B.n646 10.6151
R1315 B.n647 B.n170 10.6151
R1316 B.n651 B.n170 10.6151
R1317 B.n652 B.n651 10.6151
R1318 B.n653 B.n652 10.6151
R1319 B.n653 B.n168 10.6151
R1320 B.n657 B.n168 10.6151
R1321 B.n658 B.n657 10.6151
R1322 B.n659 B.n658 10.6151
R1323 B.n659 B.n166 10.6151
R1324 B.n663 B.n166 10.6151
R1325 B.n664 B.n663 10.6151
R1326 B.n665 B.n664 10.6151
R1327 B.n665 B.n164 10.6151
R1328 B.n669 B.n164 10.6151
R1329 B.n670 B.n669 10.6151
R1330 B.n671 B.n670 10.6151
R1331 B.n671 B.n162 10.6151
R1332 B.n675 B.n162 10.6151
R1333 B.n676 B.n675 10.6151
R1334 B.n677 B.n676 10.6151
R1335 B.n677 B.n160 10.6151
R1336 B.n681 B.n160 10.6151
R1337 B.n682 B.n681 10.6151
R1338 B.n683 B.n682 10.6151
R1339 B.n683 B.n158 10.6151
R1340 B.n687 B.n158 10.6151
R1341 B.n688 B.n687 10.6151
R1342 B.n689 B.n688 10.6151
R1343 B.n689 B.n156 10.6151
R1344 B.n693 B.n156 10.6151
R1345 B.n694 B.n693 10.6151
R1346 B.n695 B.n694 10.6151
R1347 B.n695 B.n154 10.6151
R1348 B.n699 B.n154 10.6151
R1349 B.n700 B.n699 10.6151
R1350 B.n701 B.n700 10.6151
R1351 B.n701 B.n152 10.6151
R1352 B.n705 B.n152 10.6151
R1353 B.n706 B.n705 10.6151
R1354 B.n707 B.n706 10.6151
R1355 B.n707 B.n150 10.6151
R1356 B.n711 B.n150 10.6151
R1357 B.n712 B.n711 10.6151
R1358 B.n713 B.n712 10.6151
R1359 B.n713 B.n148 10.6151
R1360 B.n717 B.n148 10.6151
R1361 B.n718 B.n717 10.6151
R1362 B.n719 B.n718 10.6151
R1363 B.n719 B.n146 10.6151
R1364 B.n723 B.n146 10.6151
R1365 B.n724 B.n723 10.6151
R1366 B.n725 B.n724 10.6151
R1367 B.n725 B.n144 10.6151
R1368 B.n729 B.n144 10.6151
R1369 B.n730 B.n729 10.6151
R1370 B.n731 B.n730 10.6151
R1371 B.n731 B.n142 10.6151
R1372 B.n735 B.n142 10.6151
R1373 B.n736 B.n735 10.6151
R1374 B.n737 B.n736 10.6151
R1375 B.n737 B.n140 10.6151
R1376 B.n741 B.n140 10.6151
R1377 B.n742 B.n741 10.6151
R1378 B.n743 B.n742 10.6151
R1379 B.n743 B.n138 10.6151
R1380 B.n747 B.n138 10.6151
R1381 B.n748 B.n747 10.6151
R1382 B.n749 B.n748 10.6151
R1383 B.n749 B.n136 10.6151
R1384 B.n753 B.n136 10.6151
R1385 B.n754 B.n753 10.6151
R1386 B.n755 B.n754 10.6151
R1387 B.n755 B.n134 10.6151
R1388 B.n759 B.n134 10.6151
R1389 B.n760 B.n759 10.6151
R1390 B.n761 B.n760 10.6151
R1391 B.n761 B.n132 10.6151
R1392 B.n765 B.n132 10.6151
R1393 B.n766 B.n765 10.6151
R1394 B.n767 B.n766 10.6151
R1395 B.n767 B.n130 10.6151
R1396 B.n771 B.n130 10.6151
R1397 B.n772 B.n771 10.6151
R1398 B.n773 B.n772 10.6151
R1399 B.n773 B.n128 10.6151
R1400 B.n777 B.n128 10.6151
R1401 B.n778 B.n777 10.6151
R1402 B.n779 B.n778 10.6151
R1403 B.n779 B.n126 10.6151
R1404 B.n783 B.n126 10.6151
R1405 B.n784 B.n783 10.6151
R1406 B.n785 B.n784 10.6151
R1407 B.n785 B.n124 10.6151
R1408 B.n789 B.n124 10.6151
R1409 B.n790 B.n789 10.6151
R1410 B.n791 B.n790 10.6151
R1411 B.n791 B.n122 10.6151
R1412 B.n795 B.n122 10.6151
R1413 B.n796 B.n795 10.6151
R1414 B.n797 B.n796 10.6151
R1415 B.n797 B.n120 10.6151
R1416 B.n801 B.n120 10.6151
R1417 B.n802 B.n801 10.6151
R1418 B.n803 B.n802 10.6151
R1419 B.n803 B.n118 10.6151
R1420 B.n807 B.n118 10.6151
R1421 B.n808 B.n807 10.6151
R1422 B.n809 B.n808 10.6151
R1423 B.n809 B.n116 10.6151
R1424 B.n813 B.n116 10.6151
R1425 B.n814 B.n813 10.6151
R1426 B.n815 B.n814 10.6151
R1427 B.n815 B.n114 10.6151
R1428 B.n819 B.n114 10.6151
R1429 B.n820 B.n819 10.6151
R1430 B.n821 B.n820 10.6151
R1431 B.n821 B.n112 10.6151
R1432 B.n825 B.n112 10.6151
R1433 B.n826 B.n825 10.6151
R1434 B.n827 B.n826 10.6151
R1435 B.n827 B.n110 10.6151
R1436 B.n406 B.n405 10.6151
R1437 B.n407 B.n406 10.6151
R1438 B.n407 B.n254 10.6151
R1439 B.n411 B.n254 10.6151
R1440 B.n412 B.n411 10.6151
R1441 B.n413 B.n412 10.6151
R1442 B.n413 B.n252 10.6151
R1443 B.n417 B.n252 10.6151
R1444 B.n418 B.n417 10.6151
R1445 B.n419 B.n418 10.6151
R1446 B.n419 B.n250 10.6151
R1447 B.n423 B.n250 10.6151
R1448 B.n424 B.n423 10.6151
R1449 B.n425 B.n424 10.6151
R1450 B.n425 B.n248 10.6151
R1451 B.n429 B.n248 10.6151
R1452 B.n430 B.n429 10.6151
R1453 B.n431 B.n430 10.6151
R1454 B.n431 B.n246 10.6151
R1455 B.n435 B.n246 10.6151
R1456 B.n436 B.n435 10.6151
R1457 B.n437 B.n436 10.6151
R1458 B.n437 B.n244 10.6151
R1459 B.n441 B.n244 10.6151
R1460 B.n442 B.n441 10.6151
R1461 B.n443 B.n442 10.6151
R1462 B.n443 B.n242 10.6151
R1463 B.n447 B.n242 10.6151
R1464 B.n448 B.n447 10.6151
R1465 B.n449 B.n448 10.6151
R1466 B.n449 B.n240 10.6151
R1467 B.n453 B.n240 10.6151
R1468 B.n454 B.n453 10.6151
R1469 B.n455 B.n454 10.6151
R1470 B.n455 B.n238 10.6151
R1471 B.n459 B.n238 10.6151
R1472 B.n460 B.n459 10.6151
R1473 B.n461 B.n460 10.6151
R1474 B.n461 B.n236 10.6151
R1475 B.n465 B.n236 10.6151
R1476 B.n466 B.n465 10.6151
R1477 B.n467 B.n466 10.6151
R1478 B.n467 B.n234 10.6151
R1479 B.n471 B.n234 10.6151
R1480 B.n472 B.n471 10.6151
R1481 B.n473 B.n472 10.6151
R1482 B.n473 B.n232 10.6151
R1483 B.n477 B.n232 10.6151
R1484 B.n478 B.n477 10.6151
R1485 B.n479 B.n478 10.6151
R1486 B.n479 B.n230 10.6151
R1487 B.n483 B.n230 10.6151
R1488 B.n484 B.n483 10.6151
R1489 B.n485 B.n484 10.6151
R1490 B.n485 B.n228 10.6151
R1491 B.n489 B.n228 10.6151
R1492 B.n490 B.n489 10.6151
R1493 B.n491 B.n490 10.6151
R1494 B.n491 B.n226 10.6151
R1495 B.n495 B.n226 10.6151
R1496 B.n498 B.n497 10.6151
R1497 B.n498 B.n222 10.6151
R1498 B.n502 B.n222 10.6151
R1499 B.n503 B.n502 10.6151
R1500 B.n504 B.n503 10.6151
R1501 B.n504 B.n220 10.6151
R1502 B.n508 B.n220 10.6151
R1503 B.n509 B.n508 10.6151
R1504 B.n510 B.n509 10.6151
R1505 B.n514 B.n513 10.6151
R1506 B.n515 B.n514 10.6151
R1507 B.n515 B.n214 10.6151
R1508 B.n519 B.n214 10.6151
R1509 B.n520 B.n519 10.6151
R1510 B.n521 B.n520 10.6151
R1511 B.n521 B.n212 10.6151
R1512 B.n525 B.n212 10.6151
R1513 B.n526 B.n525 10.6151
R1514 B.n527 B.n526 10.6151
R1515 B.n527 B.n210 10.6151
R1516 B.n531 B.n210 10.6151
R1517 B.n532 B.n531 10.6151
R1518 B.n533 B.n532 10.6151
R1519 B.n533 B.n208 10.6151
R1520 B.n537 B.n208 10.6151
R1521 B.n538 B.n537 10.6151
R1522 B.n539 B.n538 10.6151
R1523 B.n539 B.n206 10.6151
R1524 B.n543 B.n206 10.6151
R1525 B.n544 B.n543 10.6151
R1526 B.n545 B.n544 10.6151
R1527 B.n545 B.n204 10.6151
R1528 B.n549 B.n204 10.6151
R1529 B.n550 B.n549 10.6151
R1530 B.n551 B.n550 10.6151
R1531 B.n551 B.n202 10.6151
R1532 B.n555 B.n202 10.6151
R1533 B.n556 B.n555 10.6151
R1534 B.n557 B.n556 10.6151
R1535 B.n557 B.n200 10.6151
R1536 B.n561 B.n200 10.6151
R1537 B.n562 B.n561 10.6151
R1538 B.n563 B.n562 10.6151
R1539 B.n563 B.n198 10.6151
R1540 B.n567 B.n198 10.6151
R1541 B.n568 B.n567 10.6151
R1542 B.n569 B.n568 10.6151
R1543 B.n569 B.n196 10.6151
R1544 B.n573 B.n196 10.6151
R1545 B.n574 B.n573 10.6151
R1546 B.n575 B.n574 10.6151
R1547 B.n575 B.n194 10.6151
R1548 B.n579 B.n194 10.6151
R1549 B.n580 B.n579 10.6151
R1550 B.n581 B.n580 10.6151
R1551 B.n581 B.n192 10.6151
R1552 B.n585 B.n192 10.6151
R1553 B.n586 B.n585 10.6151
R1554 B.n587 B.n586 10.6151
R1555 B.n587 B.n190 10.6151
R1556 B.n591 B.n190 10.6151
R1557 B.n592 B.n591 10.6151
R1558 B.n593 B.n592 10.6151
R1559 B.n593 B.n188 10.6151
R1560 B.n597 B.n188 10.6151
R1561 B.n598 B.n597 10.6151
R1562 B.n599 B.n598 10.6151
R1563 B.n599 B.n186 10.6151
R1564 B.n603 B.n186 10.6151
R1565 B.n401 B.n256 10.6151
R1566 B.n401 B.n400 10.6151
R1567 B.n400 B.n399 10.6151
R1568 B.n399 B.n258 10.6151
R1569 B.n395 B.n258 10.6151
R1570 B.n395 B.n394 10.6151
R1571 B.n394 B.n393 10.6151
R1572 B.n393 B.n260 10.6151
R1573 B.n389 B.n260 10.6151
R1574 B.n389 B.n388 10.6151
R1575 B.n388 B.n387 10.6151
R1576 B.n387 B.n262 10.6151
R1577 B.n383 B.n262 10.6151
R1578 B.n383 B.n382 10.6151
R1579 B.n382 B.n381 10.6151
R1580 B.n381 B.n264 10.6151
R1581 B.n377 B.n264 10.6151
R1582 B.n377 B.n376 10.6151
R1583 B.n376 B.n375 10.6151
R1584 B.n375 B.n266 10.6151
R1585 B.n371 B.n266 10.6151
R1586 B.n371 B.n370 10.6151
R1587 B.n370 B.n369 10.6151
R1588 B.n369 B.n268 10.6151
R1589 B.n365 B.n268 10.6151
R1590 B.n365 B.n364 10.6151
R1591 B.n364 B.n363 10.6151
R1592 B.n363 B.n270 10.6151
R1593 B.n359 B.n270 10.6151
R1594 B.n359 B.n358 10.6151
R1595 B.n358 B.n357 10.6151
R1596 B.n357 B.n272 10.6151
R1597 B.n353 B.n272 10.6151
R1598 B.n353 B.n352 10.6151
R1599 B.n352 B.n351 10.6151
R1600 B.n351 B.n274 10.6151
R1601 B.n347 B.n274 10.6151
R1602 B.n347 B.n346 10.6151
R1603 B.n346 B.n345 10.6151
R1604 B.n345 B.n276 10.6151
R1605 B.n341 B.n276 10.6151
R1606 B.n341 B.n340 10.6151
R1607 B.n340 B.n339 10.6151
R1608 B.n339 B.n278 10.6151
R1609 B.n335 B.n278 10.6151
R1610 B.n335 B.n334 10.6151
R1611 B.n334 B.n333 10.6151
R1612 B.n333 B.n280 10.6151
R1613 B.n329 B.n280 10.6151
R1614 B.n329 B.n328 10.6151
R1615 B.n328 B.n327 10.6151
R1616 B.n327 B.n282 10.6151
R1617 B.n323 B.n282 10.6151
R1618 B.n323 B.n322 10.6151
R1619 B.n322 B.n321 10.6151
R1620 B.n321 B.n284 10.6151
R1621 B.n317 B.n284 10.6151
R1622 B.n317 B.n316 10.6151
R1623 B.n316 B.n315 10.6151
R1624 B.n315 B.n286 10.6151
R1625 B.n311 B.n286 10.6151
R1626 B.n311 B.n310 10.6151
R1627 B.n310 B.n309 10.6151
R1628 B.n309 B.n288 10.6151
R1629 B.n305 B.n288 10.6151
R1630 B.n305 B.n304 10.6151
R1631 B.n304 B.n303 10.6151
R1632 B.n303 B.n290 10.6151
R1633 B.n299 B.n290 10.6151
R1634 B.n299 B.n298 10.6151
R1635 B.n298 B.n297 10.6151
R1636 B.n297 B.n292 10.6151
R1637 B.n293 B.n292 10.6151
R1638 B.n293 B.n0 10.6151
R1639 B.n1139 B.n1 10.6151
R1640 B.n1139 B.n1138 10.6151
R1641 B.n1138 B.n1137 10.6151
R1642 B.n1137 B.n4 10.6151
R1643 B.n1133 B.n4 10.6151
R1644 B.n1133 B.n1132 10.6151
R1645 B.n1132 B.n1131 10.6151
R1646 B.n1131 B.n6 10.6151
R1647 B.n1127 B.n6 10.6151
R1648 B.n1127 B.n1126 10.6151
R1649 B.n1126 B.n1125 10.6151
R1650 B.n1125 B.n8 10.6151
R1651 B.n1121 B.n8 10.6151
R1652 B.n1121 B.n1120 10.6151
R1653 B.n1120 B.n1119 10.6151
R1654 B.n1119 B.n10 10.6151
R1655 B.n1115 B.n10 10.6151
R1656 B.n1115 B.n1114 10.6151
R1657 B.n1114 B.n1113 10.6151
R1658 B.n1113 B.n12 10.6151
R1659 B.n1109 B.n12 10.6151
R1660 B.n1109 B.n1108 10.6151
R1661 B.n1108 B.n1107 10.6151
R1662 B.n1107 B.n14 10.6151
R1663 B.n1103 B.n14 10.6151
R1664 B.n1103 B.n1102 10.6151
R1665 B.n1102 B.n1101 10.6151
R1666 B.n1101 B.n16 10.6151
R1667 B.n1097 B.n16 10.6151
R1668 B.n1097 B.n1096 10.6151
R1669 B.n1096 B.n1095 10.6151
R1670 B.n1095 B.n18 10.6151
R1671 B.n1091 B.n18 10.6151
R1672 B.n1091 B.n1090 10.6151
R1673 B.n1090 B.n1089 10.6151
R1674 B.n1089 B.n20 10.6151
R1675 B.n1085 B.n20 10.6151
R1676 B.n1085 B.n1084 10.6151
R1677 B.n1084 B.n1083 10.6151
R1678 B.n1083 B.n22 10.6151
R1679 B.n1079 B.n22 10.6151
R1680 B.n1079 B.n1078 10.6151
R1681 B.n1078 B.n1077 10.6151
R1682 B.n1077 B.n24 10.6151
R1683 B.n1073 B.n24 10.6151
R1684 B.n1073 B.n1072 10.6151
R1685 B.n1072 B.n1071 10.6151
R1686 B.n1071 B.n26 10.6151
R1687 B.n1067 B.n26 10.6151
R1688 B.n1067 B.n1066 10.6151
R1689 B.n1066 B.n1065 10.6151
R1690 B.n1065 B.n28 10.6151
R1691 B.n1061 B.n28 10.6151
R1692 B.n1061 B.n1060 10.6151
R1693 B.n1060 B.n1059 10.6151
R1694 B.n1059 B.n30 10.6151
R1695 B.n1055 B.n30 10.6151
R1696 B.n1055 B.n1054 10.6151
R1697 B.n1054 B.n1053 10.6151
R1698 B.n1053 B.n32 10.6151
R1699 B.n1049 B.n32 10.6151
R1700 B.n1049 B.n1048 10.6151
R1701 B.n1048 B.n1047 10.6151
R1702 B.n1047 B.n34 10.6151
R1703 B.n1043 B.n34 10.6151
R1704 B.n1043 B.n1042 10.6151
R1705 B.n1042 B.n1041 10.6151
R1706 B.n1041 B.n36 10.6151
R1707 B.n1037 B.n36 10.6151
R1708 B.n1037 B.n1036 10.6151
R1709 B.n1036 B.n1035 10.6151
R1710 B.n1035 B.n38 10.6151
R1711 B.n1031 B.n38 10.6151
R1712 B.n1031 B.n1030 10.6151
R1713 B.n939 B.n72 9.36635
R1714 B.n922 B.n921 9.36635
R1715 B.n496 B.n495 9.36635
R1716 B.n513 B.n218 9.36635
R1717 B.n1143 B.n0 2.81026
R1718 B.n1143 B.n1 2.81026
R1719 B.n936 B.n72 1.24928
R1720 B.n923 B.n922 1.24928
R1721 B.n497 B.n496 1.24928
R1722 B.n510 B.n218 1.24928
R1723 VP.n31 VP.t4 163.417
R1724 VP.n32 VP.n29 161.3
R1725 VP.n34 VP.n33 161.3
R1726 VP.n35 VP.n28 161.3
R1727 VP.n37 VP.n36 161.3
R1728 VP.n38 VP.n27 161.3
R1729 VP.n40 VP.n39 161.3
R1730 VP.n41 VP.n26 161.3
R1731 VP.n44 VP.n43 161.3
R1732 VP.n45 VP.n25 161.3
R1733 VP.n47 VP.n46 161.3
R1734 VP.n48 VP.n24 161.3
R1735 VP.n50 VP.n49 161.3
R1736 VP.n51 VP.n23 161.3
R1737 VP.n53 VP.n52 161.3
R1738 VP.n54 VP.n22 161.3
R1739 VP.n56 VP.n55 161.3
R1740 VP.n58 VP.n57 161.3
R1741 VP.n59 VP.n20 161.3
R1742 VP.n61 VP.n60 161.3
R1743 VP.n62 VP.n19 161.3
R1744 VP.n64 VP.n63 161.3
R1745 VP.n65 VP.n18 161.3
R1746 VP.n67 VP.n66 161.3
R1747 VP.n117 VP.n116 161.3
R1748 VP.n115 VP.n1 161.3
R1749 VP.n114 VP.n113 161.3
R1750 VP.n112 VP.n2 161.3
R1751 VP.n111 VP.n110 161.3
R1752 VP.n109 VP.n3 161.3
R1753 VP.n108 VP.n107 161.3
R1754 VP.n106 VP.n105 161.3
R1755 VP.n104 VP.n5 161.3
R1756 VP.n103 VP.n102 161.3
R1757 VP.n101 VP.n6 161.3
R1758 VP.n100 VP.n99 161.3
R1759 VP.n98 VP.n7 161.3
R1760 VP.n97 VP.n96 161.3
R1761 VP.n95 VP.n8 161.3
R1762 VP.n94 VP.n93 161.3
R1763 VP.n91 VP.n9 161.3
R1764 VP.n90 VP.n89 161.3
R1765 VP.n88 VP.n10 161.3
R1766 VP.n87 VP.n86 161.3
R1767 VP.n85 VP.n11 161.3
R1768 VP.n84 VP.n83 161.3
R1769 VP.n82 VP.n12 161.3
R1770 VP.n81 VP.n80 161.3
R1771 VP.n78 VP.n13 161.3
R1772 VP.n77 VP.n76 161.3
R1773 VP.n75 VP.n14 161.3
R1774 VP.n74 VP.n73 161.3
R1775 VP.n72 VP.n15 161.3
R1776 VP.n71 VP.n70 161.3
R1777 VP.n16 VP.t8 130.56
R1778 VP.n79 VP.t5 130.56
R1779 VP.n92 VP.t3 130.56
R1780 VP.n4 VP.t9 130.56
R1781 VP.n0 VP.t6 130.56
R1782 VP.n17 VP.t1 130.56
R1783 VP.n21 VP.t2 130.56
R1784 VP.n42 VP.t7 130.56
R1785 VP.n30 VP.t0 130.56
R1786 VP.n69 VP.n16 74.8979
R1787 VP.n118 VP.n0 74.8979
R1788 VP.n68 VP.n17 74.8979
R1789 VP.n31 VP.n30 73.2461
R1790 VP.n69 VP.n68 62.9615
R1791 VP.n86 VP.n10 54.0911
R1792 VP.n99 VP.n6 54.0911
R1793 VP.n49 VP.n23 54.0911
R1794 VP.n36 VP.n27 54.0911
R1795 VP.n77 VP.n14 48.2635
R1796 VP.n110 VP.n2 48.2635
R1797 VP.n60 VP.n19 48.2635
R1798 VP.n73 VP.n14 32.7233
R1799 VP.n114 VP.n2 32.7233
R1800 VP.n64 VP.n19 32.7233
R1801 VP.n90 VP.n10 26.8957
R1802 VP.n99 VP.n98 26.8957
R1803 VP.n49 VP.n48 26.8957
R1804 VP.n40 VP.n27 26.8957
R1805 VP.n72 VP.n71 24.4675
R1806 VP.n73 VP.n72 24.4675
R1807 VP.n78 VP.n77 24.4675
R1808 VP.n80 VP.n78 24.4675
R1809 VP.n84 VP.n12 24.4675
R1810 VP.n85 VP.n84 24.4675
R1811 VP.n86 VP.n85 24.4675
R1812 VP.n91 VP.n90 24.4675
R1813 VP.n93 VP.n91 24.4675
R1814 VP.n97 VP.n8 24.4675
R1815 VP.n98 VP.n97 24.4675
R1816 VP.n103 VP.n6 24.4675
R1817 VP.n104 VP.n103 24.4675
R1818 VP.n105 VP.n104 24.4675
R1819 VP.n109 VP.n108 24.4675
R1820 VP.n110 VP.n109 24.4675
R1821 VP.n115 VP.n114 24.4675
R1822 VP.n116 VP.n115 24.4675
R1823 VP.n65 VP.n64 24.4675
R1824 VP.n66 VP.n65 24.4675
R1825 VP.n53 VP.n23 24.4675
R1826 VP.n54 VP.n53 24.4675
R1827 VP.n55 VP.n54 24.4675
R1828 VP.n59 VP.n58 24.4675
R1829 VP.n60 VP.n59 24.4675
R1830 VP.n41 VP.n40 24.4675
R1831 VP.n43 VP.n41 24.4675
R1832 VP.n47 VP.n25 24.4675
R1833 VP.n48 VP.n47 24.4675
R1834 VP.n34 VP.n29 24.4675
R1835 VP.n35 VP.n34 24.4675
R1836 VP.n36 VP.n35 24.4675
R1837 VP.n80 VP.n79 22.9995
R1838 VP.n108 VP.n4 22.9995
R1839 VP.n58 VP.n21 22.9995
R1840 VP.n71 VP.n16 15.17
R1841 VP.n116 VP.n0 15.17
R1842 VP.n66 VP.n17 15.17
R1843 VP.n93 VP.n92 12.234
R1844 VP.n92 VP.n8 12.234
R1845 VP.n43 VP.n42 12.234
R1846 VP.n42 VP.n25 12.234
R1847 VP.n32 VP.n31 4.14768
R1848 VP.n79 VP.n12 1.46852
R1849 VP.n105 VP.n4 1.46852
R1850 VP.n55 VP.n21 1.46852
R1851 VP.n30 VP.n29 1.46852
R1852 VP.n68 VP.n67 0.354971
R1853 VP.n70 VP.n69 0.354971
R1854 VP.n118 VP.n117 0.354971
R1855 VP VP.n118 0.26696
R1856 VP.n33 VP.n32 0.189894
R1857 VP.n33 VP.n28 0.189894
R1858 VP.n37 VP.n28 0.189894
R1859 VP.n38 VP.n37 0.189894
R1860 VP.n39 VP.n38 0.189894
R1861 VP.n39 VP.n26 0.189894
R1862 VP.n44 VP.n26 0.189894
R1863 VP.n45 VP.n44 0.189894
R1864 VP.n46 VP.n45 0.189894
R1865 VP.n46 VP.n24 0.189894
R1866 VP.n50 VP.n24 0.189894
R1867 VP.n51 VP.n50 0.189894
R1868 VP.n52 VP.n51 0.189894
R1869 VP.n52 VP.n22 0.189894
R1870 VP.n56 VP.n22 0.189894
R1871 VP.n57 VP.n56 0.189894
R1872 VP.n57 VP.n20 0.189894
R1873 VP.n61 VP.n20 0.189894
R1874 VP.n62 VP.n61 0.189894
R1875 VP.n63 VP.n62 0.189894
R1876 VP.n63 VP.n18 0.189894
R1877 VP.n67 VP.n18 0.189894
R1878 VP.n70 VP.n15 0.189894
R1879 VP.n74 VP.n15 0.189894
R1880 VP.n75 VP.n74 0.189894
R1881 VP.n76 VP.n75 0.189894
R1882 VP.n76 VP.n13 0.189894
R1883 VP.n81 VP.n13 0.189894
R1884 VP.n82 VP.n81 0.189894
R1885 VP.n83 VP.n82 0.189894
R1886 VP.n83 VP.n11 0.189894
R1887 VP.n87 VP.n11 0.189894
R1888 VP.n88 VP.n87 0.189894
R1889 VP.n89 VP.n88 0.189894
R1890 VP.n89 VP.n9 0.189894
R1891 VP.n94 VP.n9 0.189894
R1892 VP.n95 VP.n94 0.189894
R1893 VP.n96 VP.n95 0.189894
R1894 VP.n96 VP.n7 0.189894
R1895 VP.n100 VP.n7 0.189894
R1896 VP.n101 VP.n100 0.189894
R1897 VP.n102 VP.n101 0.189894
R1898 VP.n102 VP.n5 0.189894
R1899 VP.n106 VP.n5 0.189894
R1900 VP.n107 VP.n106 0.189894
R1901 VP.n107 VP.n3 0.189894
R1902 VP.n111 VP.n3 0.189894
R1903 VP.n112 VP.n111 0.189894
R1904 VP.n113 VP.n112 0.189894
R1905 VP.n113 VP.n1 0.189894
R1906 VP.n117 VP.n1 0.189894
R1907 VDD1.n1 VDD1.t8 75.2757
R1908 VDD1.n3 VDD1.t2 75.2756
R1909 VDD1.n5 VDD1.n4 72.6664
R1910 VDD1.n1 VDD1.n0 70.278
R1911 VDD1.n7 VDD1.n6 70.2778
R1912 VDD1.n3 VDD1.n2 70.2777
R1913 VDD1.n7 VDD1.n5 57.5181
R1914 VDD1 VDD1.n7 2.38628
R1915 VDD1.n6 VDD1.t9 1.73967
R1916 VDD1.n6 VDD1.t6 1.73967
R1917 VDD1.n0 VDD1.t7 1.73967
R1918 VDD1.n0 VDD1.t1 1.73967
R1919 VDD1.n4 VDD1.t0 1.73967
R1920 VDD1.n4 VDD1.t4 1.73967
R1921 VDD1.n2 VDD1.t5 1.73967
R1922 VDD1.n2 VDD1.t3 1.73967
R1923 VDD1 VDD1.n1 0.873345
R1924 VDD1.n5 VDD1.n3 0.759809
R1925 VTAIL.n11 VTAIL.t5 55.3383
R1926 VTAIL.n17 VTAIL.t0 55.3382
R1927 VTAIL.n2 VTAIL.t13 55.3382
R1928 VTAIL.n16 VTAIL.t18 55.3382
R1929 VTAIL.n15 VTAIL.n14 53.5992
R1930 VTAIL.n13 VTAIL.n12 53.5992
R1931 VTAIL.n10 VTAIL.n9 53.5992
R1932 VTAIL.n8 VTAIL.n7 53.5992
R1933 VTAIL.n19 VTAIL.n18 53.599
R1934 VTAIL.n1 VTAIL.n0 53.599
R1935 VTAIL.n4 VTAIL.n3 53.599
R1936 VTAIL.n6 VTAIL.n5 53.599
R1937 VTAIL.n8 VTAIL.n6 34.9962
R1938 VTAIL.n17 VTAIL.n16 31.7376
R1939 VTAIL.n10 VTAIL.n8 3.25912
R1940 VTAIL.n11 VTAIL.n10 3.25912
R1941 VTAIL.n15 VTAIL.n13 3.25912
R1942 VTAIL.n16 VTAIL.n15 3.25912
R1943 VTAIL.n6 VTAIL.n4 3.25912
R1944 VTAIL.n4 VTAIL.n2 3.25912
R1945 VTAIL.n19 VTAIL.n17 3.25912
R1946 VTAIL VTAIL.n1 2.50266
R1947 VTAIL.n13 VTAIL.n11 2.09964
R1948 VTAIL.n2 VTAIL.n1 2.09964
R1949 VTAIL.n18 VTAIL.t7 1.73967
R1950 VTAIL.n18 VTAIL.t4 1.73967
R1951 VTAIL.n0 VTAIL.t3 1.73967
R1952 VTAIL.n0 VTAIL.t1 1.73967
R1953 VTAIL.n3 VTAIL.t16 1.73967
R1954 VTAIL.n3 VTAIL.t10 1.73967
R1955 VTAIL.n5 VTAIL.t11 1.73967
R1956 VTAIL.n5 VTAIL.t14 1.73967
R1957 VTAIL.n14 VTAIL.t12 1.73967
R1958 VTAIL.n14 VTAIL.t17 1.73967
R1959 VTAIL.n12 VTAIL.t15 1.73967
R1960 VTAIL.n12 VTAIL.t19 1.73967
R1961 VTAIL.n9 VTAIL.t8 1.73967
R1962 VTAIL.n9 VTAIL.t9 1.73967
R1963 VTAIL.n7 VTAIL.t6 1.73967
R1964 VTAIL.n7 VTAIL.t2 1.73967
R1965 VTAIL VTAIL.n19 0.756965
R1966 VN.n67 VN.t4 163.417
R1967 VN.n14 VN.t6 163.417
R1968 VN.n102 VN.n101 161.3
R1969 VN.n100 VN.n53 161.3
R1970 VN.n99 VN.n98 161.3
R1971 VN.n97 VN.n54 161.3
R1972 VN.n96 VN.n95 161.3
R1973 VN.n94 VN.n55 161.3
R1974 VN.n93 VN.n92 161.3
R1975 VN.n91 VN.n90 161.3
R1976 VN.n89 VN.n57 161.3
R1977 VN.n88 VN.n87 161.3
R1978 VN.n86 VN.n58 161.3
R1979 VN.n85 VN.n84 161.3
R1980 VN.n83 VN.n59 161.3
R1981 VN.n82 VN.n81 161.3
R1982 VN.n80 VN.n60 161.3
R1983 VN.n79 VN.n78 161.3
R1984 VN.n77 VN.n61 161.3
R1985 VN.n76 VN.n75 161.3
R1986 VN.n74 VN.n63 161.3
R1987 VN.n73 VN.n72 161.3
R1988 VN.n71 VN.n64 161.3
R1989 VN.n70 VN.n69 161.3
R1990 VN.n68 VN.n65 161.3
R1991 VN.n50 VN.n49 161.3
R1992 VN.n48 VN.n1 161.3
R1993 VN.n47 VN.n46 161.3
R1994 VN.n45 VN.n2 161.3
R1995 VN.n44 VN.n43 161.3
R1996 VN.n42 VN.n3 161.3
R1997 VN.n41 VN.n40 161.3
R1998 VN.n39 VN.n38 161.3
R1999 VN.n37 VN.n5 161.3
R2000 VN.n36 VN.n35 161.3
R2001 VN.n34 VN.n6 161.3
R2002 VN.n33 VN.n32 161.3
R2003 VN.n31 VN.n7 161.3
R2004 VN.n30 VN.n29 161.3
R2005 VN.n28 VN.n8 161.3
R2006 VN.n27 VN.n26 161.3
R2007 VN.n24 VN.n9 161.3
R2008 VN.n23 VN.n22 161.3
R2009 VN.n21 VN.n10 161.3
R2010 VN.n20 VN.n19 161.3
R2011 VN.n18 VN.n11 161.3
R2012 VN.n17 VN.n16 161.3
R2013 VN.n15 VN.n12 161.3
R2014 VN.n13 VN.t8 130.56
R2015 VN.n25 VN.t2 130.56
R2016 VN.n4 VN.t5 130.56
R2017 VN.n0 VN.t9 130.56
R2018 VN.n66 VN.t0 130.56
R2019 VN.n62 VN.t1 130.56
R2020 VN.n56 VN.t7 130.56
R2021 VN.n52 VN.t3 130.56
R2022 VN.n51 VN.n0 74.8979
R2023 VN.n103 VN.n52 74.8979
R2024 VN.n14 VN.n13 73.246
R2025 VN.n67 VN.n66 73.246
R2026 VN VN.n103 63.1268
R2027 VN.n19 VN.n10 54.0911
R2028 VN.n32 VN.n6 54.0911
R2029 VN.n72 VN.n63 54.0911
R2030 VN.n84 VN.n58 54.0911
R2031 VN.n43 VN.n2 48.2635
R2032 VN.n95 VN.n54 48.2635
R2033 VN.n47 VN.n2 32.7233
R2034 VN.n99 VN.n54 32.7233
R2035 VN.n23 VN.n10 26.8957
R2036 VN.n32 VN.n31 26.8957
R2037 VN.n76 VN.n63 26.8957
R2038 VN.n84 VN.n83 26.8957
R2039 VN.n17 VN.n12 24.4675
R2040 VN.n18 VN.n17 24.4675
R2041 VN.n19 VN.n18 24.4675
R2042 VN.n24 VN.n23 24.4675
R2043 VN.n26 VN.n24 24.4675
R2044 VN.n30 VN.n8 24.4675
R2045 VN.n31 VN.n30 24.4675
R2046 VN.n36 VN.n6 24.4675
R2047 VN.n37 VN.n36 24.4675
R2048 VN.n38 VN.n37 24.4675
R2049 VN.n42 VN.n41 24.4675
R2050 VN.n43 VN.n42 24.4675
R2051 VN.n48 VN.n47 24.4675
R2052 VN.n49 VN.n48 24.4675
R2053 VN.n72 VN.n71 24.4675
R2054 VN.n71 VN.n70 24.4675
R2055 VN.n70 VN.n65 24.4675
R2056 VN.n83 VN.n82 24.4675
R2057 VN.n82 VN.n60 24.4675
R2058 VN.n78 VN.n77 24.4675
R2059 VN.n77 VN.n76 24.4675
R2060 VN.n95 VN.n94 24.4675
R2061 VN.n94 VN.n93 24.4675
R2062 VN.n90 VN.n89 24.4675
R2063 VN.n89 VN.n88 24.4675
R2064 VN.n88 VN.n58 24.4675
R2065 VN.n101 VN.n100 24.4675
R2066 VN.n100 VN.n99 24.4675
R2067 VN.n41 VN.n4 22.9995
R2068 VN.n93 VN.n56 22.9995
R2069 VN.n49 VN.n0 15.17
R2070 VN.n101 VN.n52 15.17
R2071 VN.n26 VN.n25 12.234
R2072 VN.n25 VN.n8 12.234
R2073 VN.n62 VN.n60 12.234
R2074 VN.n78 VN.n62 12.234
R2075 VN.n15 VN.n14 4.14771
R2076 VN.n68 VN.n67 4.14771
R2077 VN.n13 VN.n12 1.46852
R2078 VN.n38 VN.n4 1.46852
R2079 VN.n66 VN.n65 1.46852
R2080 VN.n90 VN.n56 1.46852
R2081 VN.n103 VN.n102 0.354971
R2082 VN.n51 VN.n50 0.354971
R2083 VN VN.n51 0.26696
R2084 VN.n102 VN.n53 0.189894
R2085 VN.n98 VN.n53 0.189894
R2086 VN.n98 VN.n97 0.189894
R2087 VN.n97 VN.n96 0.189894
R2088 VN.n96 VN.n55 0.189894
R2089 VN.n92 VN.n55 0.189894
R2090 VN.n92 VN.n91 0.189894
R2091 VN.n91 VN.n57 0.189894
R2092 VN.n87 VN.n57 0.189894
R2093 VN.n87 VN.n86 0.189894
R2094 VN.n86 VN.n85 0.189894
R2095 VN.n85 VN.n59 0.189894
R2096 VN.n81 VN.n59 0.189894
R2097 VN.n81 VN.n80 0.189894
R2098 VN.n80 VN.n79 0.189894
R2099 VN.n79 VN.n61 0.189894
R2100 VN.n75 VN.n61 0.189894
R2101 VN.n75 VN.n74 0.189894
R2102 VN.n74 VN.n73 0.189894
R2103 VN.n73 VN.n64 0.189894
R2104 VN.n69 VN.n64 0.189894
R2105 VN.n69 VN.n68 0.189894
R2106 VN.n16 VN.n15 0.189894
R2107 VN.n16 VN.n11 0.189894
R2108 VN.n20 VN.n11 0.189894
R2109 VN.n21 VN.n20 0.189894
R2110 VN.n22 VN.n21 0.189894
R2111 VN.n22 VN.n9 0.189894
R2112 VN.n27 VN.n9 0.189894
R2113 VN.n28 VN.n27 0.189894
R2114 VN.n29 VN.n28 0.189894
R2115 VN.n29 VN.n7 0.189894
R2116 VN.n33 VN.n7 0.189894
R2117 VN.n34 VN.n33 0.189894
R2118 VN.n35 VN.n34 0.189894
R2119 VN.n35 VN.n5 0.189894
R2120 VN.n39 VN.n5 0.189894
R2121 VN.n40 VN.n39 0.189894
R2122 VN.n40 VN.n3 0.189894
R2123 VN.n44 VN.n3 0.189894
R2124 VN.n45 VN.n44 0.189894
R2125 VN.n46 VN.n45 0.189894
R2126 VN.n46 VN.n1 0.189894
R2127 VN.n50 VN.n1 0.189894
R2128 VDD2.n1 VDD2.t3 75.2756
R2129 VDD2.n3 VDD2.n2 72.6664
R2130 VDD2 VDD2.n7 72.6636
R2131 VDD2.n4 VDD2.t6 72.0171
R2132 VDD2.n6 VDD2.n5 70.278
R2133 VDD2.n1 VDD2.n0 70.2777
R2134 VDD2.n4 VDD2.n3 55.3058
R2135 VDD2.n6 VDD2.n4 3.25912
R2136 VDD2.n7 VDD2.t9 1.73967
R2137 VDD2.n7 VDD2.t5 1.73967
R2138 VDD2.n5 VDD2.t2 1.73967
R2139 VDD2.n5 VDD2.t8 1.73967
R2140 VDD2.n2 VDD2.t4 1.73967
R2141 VDD2.n2 VDD2.t0 1.73967
R2142 VDD2.n0 VDD2.t1 1.73967
R2143 VDD2.n0 VDD2.t7 1.73967
R2144 VDD2 VDD2.n6 0.873345
R2145 VDD2.n3 VDD2.n1 0.759809
C0 VDD1 B 3.34883f
C1 VP w_n5506_n4706# 12.8741f
C2 VN w_n5506_n4706# 12.154599f
C3 VTAIL w_n5506_n4706# 4.24138f
C4 VN VP 10.8888f
C5 VTAIL VP 17.870302f
C6 VDD2 w_n5506_n4706# 3.75705f
C7 VDD2 VP 0.692418f
C8 VTAIL VN 17.856f
C9 VDD2 VN 17.1637f
C10 VDD2 VTAIL 13.527901f
C11 B w_n5506_n4706# 13.8514f
C12 B VP 2.79269f
C13 VDD1 w_n5506_n4706# 3.56932f
C14 B VN 1.57816f
C15 VDD1 VP 17.696098f
C16 B VTAIL 5.63255f
C17 VDD1 VN 0.155265f
C18 B VDD2 3.49984f
C19 VDD1 VTAIL 13.4717f
C20 VDD1 VDD2 2.72841f
C21 VDD2 VSUBS 2.59914f
C22 VDD1 VSUBS 2.478714f
C23 VTAIL VSUBS 1.730414f
C24 VN VSUBS 9.327741f
C25 VP VSUBS 5.569039f
C26 B VSUBS 6.98488f
C27 w_n5506_n4706# VSUBS 0.316683p
C28 VDD2.t3 VSUBS 4.651721f
C29 VDD2.t1 VSUBS 0.424923f
C30 VDD2.t7 VSUBS 0.424923f
C31 VDD2.n0 VSUBS 3.55399f
C32 VDD2.n1 VSUBS 1.87304f
C33 VDD2.t4 VSUBS 0.424923f
C34 VDD2.t0 VSUBS 0.424923f
C35 VDD2.n2 VSUBS 3.59007f
C36 VDD2.n3 VSUBS 4.65578f
C37 VDD2.t6 VSUBS 4.60933f
C38 VDD2.n4 VSUBS 4.91391f
C39 VDD2.t2 VSUBS 0.424923f
C40 VDD2.t8 VSUBS 0.424923f
C41 VDD2.n5 VSUBS 3.55399f
C42 VDD2.n6 VSUBS 0.945428f
C43 VDD2.t9 VSUBS 0.424923f
C44 VDD2.t5 VSUBS 0.424923f
C45 VDD2.n7 VSUBS 3.59001f
C46 VN.t9 VSUBS 3.78168f
C47 VN.n0 VSUBS 1.39106f
C48 VN.n1 VSUBS 0.021307f
C49 VN.n2 VSUBS 0.019043f
C50 VN.n3 VSUBS 0.021307f
C51 VN.t5 VSUBS 3.78168f
C52 VN.n4 VSUBS 1.30306f
C53 VN.n5 VSUBS 0.021307f
C54 VN.n6 VSUBS 0.037348f
C55 VN.n7 VSUBS 0.021307f
C56 VN.n8 VSUBS 0.029909f
C57 VN.n9 VSUBS 0.021307f
C58 VN.n10 VSUBS 0.02327f
C59 VN.n11 VSUBS 0.021307f
C60 VN.n12 VSUBS 0.021282f
C61 VN.t8 VSUBS 3.78168f
C62 VN.n13 VSUBS 1.36843f
C63 VN.t6 VSUBS 4.07519f
C64 VN.n14 VSUBS 1.31329f
C65 VN.n15 VSUBS 0.25423f
C66 VN.n16 VSUBS 0.021307f
C67 VN.n17 VSUBS 0.039712f
C68 VN.n18 VSUBS 0.039712f
C69 VN.n19 VSUBS 0.037348f
C70 VN.n20 VSUBS 0.021307f
C71 VN.n21 VSUBS 0.021307f
C72 VN.n22 VSUBS 0.021307f
C73 VN.n23 VSUBS 0.041304f
C74 VN.n24 VSUBS 0.039712f
C75 VN.t2 VSUBS 3.78168f
C76 VN.n25 VSUBS 1.30306f
C77 VN.n26 VSUBS 0.029909f
C78 VN.n27 VSUBS 0.021307f
C79 VN.n28 VSUBS 0.021307f
C80 VN.n29 VSUBS 0.021307f
C81 VN.n30 VSUBS 0.039712f
C82 VN.n31 VSUBS 0.041304f
C83 VN.n32 VSUBS 0.02327f
C84 VN.n33 VSUBS 0.021307f
C85 VN.n34 VSUBS 0.021307f
C86 VN.n35 VSUBS 0.021307f
C87 VN.n36 VSUBS 0.039712f
C88 VN.n37 VSUBS 0.039712f
C89 VN.n38 VSUBS 0.021282f
C90 VN.n39 VSUBS 0.021307f
C91 VN.n40 VSUBS 0.021307f
C92 VN.n41 VSUBS 0.038535f
C93 VN.n42 VSUBS 0.039712f
C94 VN.n43 VSUBS 0.039903f
C95 VN.n44 VSUBS 0.021307f
C96 VN.n45 VSUBS 0.021307f
C97 VN.n46 VSUBS 0.021307f
C98 VN.n47 VSUBS 0.042975f
C99 VN.n48 VSUBS 0.039712f
C100 VN.n49 VSUBS 0.032261f
C101 VN.n50 VSUBS 0.03439f
C102 VN.n51 VSUBS 0.052426f
C103 VN.t3 VSUBS 3.78168f
C104 VN.n52 VSUBS 1.39106f
C105 VN.n53 VSUBS 0.021307f
C106 VN.n54 VSUBS 0.019043f
C107 VN.n55 VSUBS 0.021307f
C108 VN.t7 VSUBS 3.78168f
C109 VN.n56 VSUBS 1.30306f
C110 VN.n57 VSUBS 0.021307f
C111 VN.n58 VSUBS 0.037348f
C112 VN.n59 VSUBS 0.021307f
C113 VN.n60 VSUBS 0.029909f
C114 VN.n61 VSUBS 0.021307f
C115 VN.t1 VSUBS 3.78168f
C116 VN.n62 VSUBS 1.30306f
C117 VN.n63 VSUBS 0.02327f
C118 VN.n64 VSUBS 0.021307f
C119 VN.n65 VSUBS 0.021282f
C120 VN.t4 VSUBS 4.07519f
C121 VN.t0 VSUBS 3.78168f
C122 VN.n66 VSUBS 1.36843f
C123 VN.n67 VSUBS 1.31329f
C124 VN.n68 VSUBS 0.25423f
C125 VN.n69 VSUBS 0.021307f
C126 VN.n70 VSUBS 0.039712f
C127 VN.n71 VSUBS 0.039712f
C128 VN.n72 VSUBS 0.037348f
C129 VN.n73 VSUBS 0.021307f
C130 VN.n74 VSUBS 0.021307f
C131 VN.n75 VSUBS 0.021307f
C132 VN.n76 VSUBS 0.041304f
C133 VN.n77 VSUBS 0.039712f
C134 VN.n78 VSUBS 0.029909f
C135 VN.n79 VSUBS 0.021307f
C136 VN.n80 VSUBS 0.021307f
C137 VN.n81 VSUBS 0.021307f
C138 VN.n82 VSUBS 0.039712f
C139 VN.n83 VSUBS 0.041304f
C140 VN.n84 VSUBS 0.02327f
C141 VN.n85 VSUBS 0.021307f
C142 VN.n86 VSUBS 0.021307f
C143 VN.n87 VSUBS 0.021307f
C144 VN.n88 VSUBS 0.039712f
C145 VN.n89 VSUBS 0.039712f
C146 VN.n90 VSUBS 0.021282f
C147 VN.n91 VSUBS 0.021307f
C148 VN.n92 VSUBS 0.021307f
C149 VN.n93 VSUBS 0.038535f
C150 VN.n94 VSUBS 0.039712f
C151 VN.n95 VSUBS 0.039903f
C152 VN.n96 VSUBS 0.021307f
C153 VN.n97 VSUBS 0.021307f
C154 VN.n98 VSUBS 0.021307f
C155 VN.n99 VSUBS 0.042975f
C156 VN.n100 VSUBS 0.039712f
C157 VN.n101 VSUBS 0.032261f
C158 VN.n102 VSUBS 0.03439f
C159 VN.n103 VSUBS 1.67353f
C160 VTAIL.t3 VSUBS 0.409554f
C161 VTAIL.t1 VSUBS 0.409554f
C162 VTAIL.n0 VSUBS 3.25841f
C163 VTAIL.n1 VSUBS 1.08257f
C164 VTAIL.t13 VSUBS 4.25072f
C165 VTAIL.n2 VSUBS 1.27481f
C166 VTAIL.t16 VSUBS 0.409554f
C167 VTAIL.t10 VSUBS 0.409554f
C168 VTAIL.n3 VSUBS 3.25841f
C169 VTAIL.n4 VSUBS 1.25376f
C170 VTAIL.t11 VSUBS 0.409554f
C171 VTAIL.t14 VSUBS 0.409554f
C172 VTAIL.n5 VSUBS 3.25841f
C173 VTAIL.n6 VSUBS 3.36125f
C174 VTAIL.t6 VSUBS 0.409554f
C175 VTAIL.t2 VSUBS 0.409554f
C176 VTAIL.n7 VSUBS 3.25841f
C177 VTAIL.n8 VSUBS 3.36125f
C178 VTAIL.t8 VSUBS 0.409554f
C179 VTAIL.t9 VSUBS 0.409554f
C180 VTAIL.n9 VSUBS 3.25841f
C181 VTAIL.n10 VSUBS 1.25376f
C182 VTAIL.t5 VSUBS 4.25075f
C183 VTAIL.n11 VSUBS 1.27478f
C184 VTAIL.t15 VSUBS 0.409554f
C185 VTAIL.t19 VSUBS 0.409554f
C186 VTAIL.n12 VSUBS 3.25841f
C187 VTAIL.n13 VSUBS 1.15016f
C188 VTAIL.t12 VSUBS 0.409554f
C189 VTAIL.t17 VSUBS 0.409554f
C190 VTAIL.n14 VSUBS 3.25841f
C191 VTAIL.n15 VSUBS 1.25376f
C192 VTAIL.t18 VSUBS 4.25072f
C193 VTAIL.n16 VSUBS 3.19474f
C194 VTAIL.t0 VSUBS 4.25072f
C195 VTAIL.n17 VSUBS 3.19474f
C196 VTAIL.t7 VSUBS 0.409554f
C197 VTAIL.t4 VSUBS 0.409554f
C198 VTAIL.n18 VSUBS 3.25841f
C199 VTAIL.n19 VSUBS 1.03019f
C200 VDD1.t8 VSUBS 4.65102f
C201 VDD1.t7 VSUBS 0.424858f
C202 VDD1.t1 VSUBS 0.424858f
C203 VDD1.n0 VSUBS 3.55345f
C204 VDD1.n1 VSUBS 1.88237f
C205 VDD1.t2 VSUBS 4.651f
C206 VDD1.t5 VSUBS 0.424858f
C207 VDD1.t3 VSUBS 0.424858f
C208 VDD1.n2 VSUBS 3.55344f
C209 VDD1.n3 VSUBS 1.87275f
C210 VDD1.t0 VSUBS 0.424858f
C211 VDD1.t4 VSUBS 0.424858f
C212 VDD1.n4 VSUBS 3.58952f
C213 VDD1.n5 VSUBS 4.83095f
C214 VDD1.t9 VSUBS 0.424858f
C215 VDD1.t6 VSUBS 0.424858f
C216 VDD1.n6 VSUBS 3.55343f
C217 VDD1.n7 VSUBS 4.96115f
C218 VP.t6 VSUBS 4.04367f
C219 VP.n0 VSUBS 1.48743f
C220 VP.n1 VSUBS 0.022784f
C221 VP.n2 VSUBS 0.020363f
C222 VP.n3 VSUBS 0.022784f
C223 VP.t9 VSUBS 4.04367f
C224 VP.n4 VSUBS 1.39333f
C225 VP.n5 VSUBS 0.022784f
C226 VP.n6 VSUBS 0.039935f
C227 VP.n7 VSUBS 0.022784f
C228 VP.n8 VSUBS 0.031981f
C229 VP.n9 VSUBS 0.022784f
C230 VP.n10 VSUBS 0.024883f
C231 VP.n11 VSUBS 0.022784f
C232 VP.n12 VSUBS 0.022757f
C233 VP.n13 VSUBS 0.022784f
C234 VP.n14 VSUBS 0.020363f
C235 VP.n15 VSUBS 0.022784f
C236 VP.t8 VSUBS 4.04367f
C237 VP.n16 VSUBS 1.48743f
C238 VP.t1 VSUBS 4.04367f
C239 VP.n17 VSUBS 1.48743f
C240 VP.n18 VSUBS 0.022784f
C241 VP.n19 VSUBS 0.020363f
C242 VP.n20 VSUBS 0.022784f
C243 VP.t2 VSUBS 4.04367f
C244 VP.n21 VSUBS 1.39333f
C245 VP.n22 VSUBS 0.022784f
C246 VP.n23 VSUBS 0.039935f
C247 VP.n24 VSUBS 0.022784f
C248 VP.n25 VSUBS 0.031981f
C249 VP.n26 VSUBS 0.022784f
C250 VP.n27 VSUBS 0.024883f
C251 VP.n28 VSUBS 0.022784f
C252 VP.n29 VSUBS 0.022757f
C253 VP.t4 VSUBS 4.35751f
C254 VP.t0 VSUBS 4.04367f
C255 VP.n30 VSUBS 1.46323f
C256 VP.n31 VSUBS 1.40427f
C257 VP.n32 VSUBS 0.271843f
C258 VP.n33 VSUBS 0.022784f
C259 VP.n34 VSUBS 0.042463f
C260 VP.n35 VSUBS 0.042463f
C261 VP.n36 VSUBS 0.039935f
C262 VP.n37 VSUBS 0.022784f
C263 VP.n38 VSUBS 0.022784f
C264 VP.n39 VSUBS 0.022784f
C265 VP.n40 VSUBS 0.044165f
C266 VP.n41 VSUBS 0.042463f
C267 VP.t7 VSUBS 4.04367f
C268 VP.n42 VSUBS 1.39333f
C269 VP.n43 VSUBS 0.031981f
C270 VP.n44 VSUBS 0.022784f
C271 VP.n45 VSUBS 0.022784f
C272 VP.n46 VSUBS 0.022784f
C273 VP.n47 VSUBS 0.042463f
C274 VP.n48 VSUBS 0.044165f
C275 VP.n49 VSUBS 0.024883f
C276 VP.n50 VSUBS 0.022784f
C277 VP.n51 VSUBS 0.022784f
C278 VP.n52 VSUBS 0.022784f
C279 VP.n53 VSUBS 0.042463f
C280 VP.n54 VSUBS 0.042463f
C281 VP.n55 VSUBS 0.022757f
C282 VP.n56 VSUBS 0.022784f
C283 VP.n57 VSUBS 0.022784f
C284 VP.n58 VSUBS 0.041205f
C285 VP.n59 VSUBS 0.042463f
C286 VP.n60 VSUBS 0.042668f
C287 VP.n61 VSUBS 0.022784f
C288 VP.n62 VSUBS 0.022784f
C289 VP.n63 VSUBS 0.022784f
C290 VP.n64 VSUBS 0.045952f
C291 VP.n65 VSUBS 0.042463f
C292 VP.n66 VSUBS 0.034496f
C293 VP.n67 VSUBS 0.036772f
C294 VP.n68 VSUBS 1.78082f
C295 VP.n69 VSUBS 1.79382f
C296 VP.n70 VSUBS 0.036772f
C297 VP.n71 VSUBS 0.034496f
C298 VP.n72 VSUBS 0.042463f
C299 VP.n73 VSUBS 0.045952f
C300 VP.n74 VSUBS 0.022784f
C301 VP.n75 VSUBS 0.022784f
C302 VP.n76 VSUBS 0.022784f
C303 VP.n77 VSUBS 0.042668f
C304 VP.n78 VSUBS 0.042463f
C305 VP.t5 VSUBS 4.04367f
C306 VP.n79 VSUBS 1.39333f
C307 VP.n80 VSUBS 0.041205f
C308 VP.n81 VSUBS 0.022784f
C309 VP.n82 VSUBS 0.022784f
C310 VP.n83 VSUBS 0.022784f
C311 VP.n84 VSUBS 0.042463f
C312 VP.n85 VSUBS 0.042463f
C313 VP.n86 VSUBS 0.039935f
C314 VP.n87 VSUBS 0.022784f
C315 VP.n88 VSUBS 0.022784f
C316 VP.n89 VSUBS 0.022784f
C317 VP.n90 VSUBS 0.044165f
C318 VP.n91 VSUBS 0.042463f
C319 VP.t3 VSUBS 4.04367f
C320 VP.n92 VSUBS 1.39333f
C321 VP.n93 VSUBS 0.031981f
C322 VP.n94 VSUBS 0.022784f
C323 VP.n95 VSUBS 0.022784f
C324 VP.n96 VSUBS 0.022784f
C325 VP.n97 VSUBS 0.042463f
C326 VP.n98 VSUBS 0.044165f
C327 VP.n99 VSUBS 0.024883f
C328 VP.n100 VSUBS 0.022784f
C329 VP.n101 VSUBS 0.022784f
C330 VP.n102 VSUBS 0.022784f
C331 VP.n103 VSUBS 0.042463f
C332 VP.n104 VSUBS 0.042463f
C333 VP.n105 VSUBS 0.022757f
C334 VP.n106 VSUBS 0.022784f
C335 VP.n107 VSUBS 0.022784f
C336 VP.n108 VSUBS 0.041205f
C337 VP.n109 VSUBS 0.042463f
C338 VP.n110 VSUBS 0.042668f
C339 VP.n111 VSUBS 0.022784f
C340 VP.n112 VSUBS 0.022784f
C341 VP.n113 VSUBS 0.022784f
C342 VP.n114 VSUBS 0.045952f
C343 VP.n115 VSUBS 0.042463f
C344 VP.n116 VSUBS 0.034496f
C345 VP.n117 VSUBS 0.036772f
C346 VP.n118 VSUBS 0.056058f
C347 B.n0 VSUBS 0.004796f
C348 B.n1 VSUBS 0.004796f
C349 B.n2 VSUBS 0.007585f
C350 B.n3 VSUBS 0.007585f
C351 B.n4 VSUBS 0.007585f
C352 B.n5 VSUBS 0.007585f
C353 B.n6 VSUBS 0.007585f
C354 B.n7 VSUBS 0.007585f
C355 B.n8 VSUBS 0.007585f
C356 B.n9 VSUBS 0.007585f
C357 B.n10 VSUBS 0.007585f
C358 B.n11 VSUBS 0.007585f
C359 B.n12 VSUBS 0.007585f
C360 B.n13 VSUBS 0.007585f
C361 B.n14 VSUBS 0.007585f
C362 B.n15 VSUBS 0.007585f
C363 B.n16 VSUBS 0.007585f
C364 B.n17 VSUBS 0.007585f
C365 B.n18 VSUBS 0.007585f
C366 B.n19 VSUBS 0.007585f
C367 B.n20 VSUBS 0.007585f
C368 B.n21 VSUBS 0.007585f
C369 B.n22 VSUBS 0.007585f
C370 B.n23 VSUBS 0.007585f
C371 B.n24 VSUBS 0.007585f
C372 B.n25 VSUBS 0.007585f
C373 B.n26 VSUBS 0.007585f
C374 B.n27 VSUBS 0.007585f
C375 B.n28 VSUBS 0.007585f
C376 B.n29 VSUBS 0.007585f
C377 B.n30 VSUBS 0.007585f
C378 B.n31 VSUBS 0.007585f
C379 B.n32 VSUBS 0.007585f
C380 B.n33 VSUBS 0.007585f
C381 B.n34 VSUBS 0.007585f
C382 B.n35 VSUBS 0.007585f
C383 B.n36 VSUBS 0.007585f
C384 B.n37 VSUBS 0.007585f
C385 B.n38 VSUBS 0.007585f
C386 B.n39 VSUBS 0.017051f
C387 B.n40 VSUBS 0.007585f
C388 B.n41 VSUBS 0.007585f
C389 B.n42 VSUBS 0.007585f
C390 B.n43 VSUBS 0.007585f
C391 B.n44 VSUBS 0.007585f
C392 B.n45 VSUBS 0.007585f
C393 B.n46 VSUBS 0.007585f
C394 B.n47 VSUBS 0.007585f
C395 B.n48 VSUBS 0.007585f
C396 B.n49 VSUBS 0.007585f
C397 B.n50 VSUBS 0.007585f
C398 B.n51 VSUBS 0.007585f
C399 B.n52 VSUBS 0.007585f
C400 B.n53 VSUBS 0.007585f
C401 B.n54 VSUBS 0.007585f
C402 B.n55 VSUBS 0.007585f
C403 B.n56 VSUBS 0.007585f
C404 B.n57 VSUBS 0.007585f
C405 B.n58 VSUBS 0.007585f
C406 B.n59 VSUBS 0.007585f
C407 B.n60 VSUBS 0.007585f
C408 B.n61 VSUBS 0.007585f
C409 B.n62 VSUBS 0.007585f
C410 B.n63 VSUBS 0.007585f
C411 B.n64 VSUBS 0.007585f
C412 B.n65 VSUBS 0.007585f
C413 B.n66 VSUBS 0.007585f
C414 B.n67 VSUBS 0.007585f
C415 B.n68 VSUBS 0.007585f
C416 B.n69 VSUBS 0.007585f
C417 B.t8 VSUBS 0.68549f
C418 B.t7 VSUBS 0.713556f
C419 B.t6 VSUBS 3.15535f
C420 B.n70 VSUBS 0.436089f
C421 B.n71 VSUBS 0.081958f
C422 B.n72 VSUBS 0.017574f
C423 B.n73 VSUBS 0.007585f
C424 B.n74 VSUBS 0.007585f
C425 B.n75 VSUBS 0.007585f
C426 B.n76 VSUBS 0.007585f
C427 B.n77 VSUBS 0.007585f
C428 B.t5 VSUBS 0.685464f
C429 B.t4 VSUBS 0.713536f
C430 B.t3 VSUBS 3.15535f
C431 B.n78 VSUBS 0.436109f
C432 B.n79 VSUBS 0.081984f
C433 B.n80 VSUBS 0.007585f
C434 B.n81 VSUBS 0.007585f
C435 B.n82 VSUBS 0.007585f
C436 B.n83 VSUBS 0.007585f
C437 B.n84 VSUBS 0.007585f
C438 B.n85 VSUBS 0.007585f
C439 B.n86 VSUBS 0.007585f
C440 B.n87 VSUBS 0.007585f
C441 B.n88 VSUBS 0.007585f
C442 B.n89 VSUBS 0.007585f
C443 B.n90 VSUBS 0.007585f
C444 B.n91 VSUBS 0.007585f
C445 B.n92 VSUBS 0.007585f
C446 B.n93 VSUBS 0.007585f
C447 B.n94 VSUBS 0.007585f
C448 B.n95 VSUBS 0.007585f
C449 B.n96 VSUBS 0.007585f
C450 B.n97 VSUBS 0.007585f
C451 B.n98 VSUBS 0.007585f
C452 B.n99 VSUBS 0.007585f
C453 B.n100 VSUBS 0.007585f
C454 B.n101 VSUBS 0.007585f
C455 B.n102 VSUBS 0.007585f
C456 B.n103 VSUBS 0.007585f
C457 B.n104 VSUBS 0.007585f
C458 B.n105 VSUBS 0.007585f
C459 B.n106 VSUBS 0.007585f
C460 B.n107 VSUBS 0.007585f
C461 B.n108 VSUBS 0.007585f
C462 B.n109 VSUBS 0.007585f
C463 B.n110 VSUBS 0.017983f
C464 B.n111 VSUBS 0.007585f
C465 B.n112 VSUBS 0.007585f
C466 B.n113 VSUBS 0.007585f
C467 B.n114 VSUBS 0.007585f
C468 B.n115 VSUBS 0.007585f
C469 B.n116 VSUBS 0.007585f
C470 B.n117 VSUBS 0.007585f
C471 B.n118 VSUBS 0.007585f
C472 B.n119 VSUBS 0.007585f
C473 B.n120 VSUBS 0.007585f
C474 B.n121 VSUBS 0.007585f
C475 B.n122 VSUBS 0.007585f
C476 B.n123 VSUBS 0.007585f
C477 B.n124 VSUBS 0.007585f
C478 B.n125 VSUBS 0.007585f
C479 B.n126 VSUBS 0.007585f
C480 B.n127 VSUBS 0.007585f
C481 B.n128 VSUBS 0.007585f
C482 B.n129 VSUBS 0.007585f
C483 B.n130 VSUBS 0.007585f
C484 B.n131 VSUBS 0.007585f
C485 B.n132 VSUBS 0.007585f
C486 B.n133 VSUBS 0.007585f
C487 B.n134 VSUBS 0.007585f
C488 B.n135 VSUBS 0.007585f
C489 B.n136 VSUBS 0.007585f
C490 B.n137 VSUBS 0.007585f
C491 B.n138 VSUBS 0.007585f
C492 B.n139 VSUBS 0.007585f
C493 B.n140 VSUBS 0.007585f
C494 B.n141 VSUBS 0.007585f
C495 B.n142 VSUBS 0.007585f
C496 B.n143 VSUBS 0.007585f
C497 B.n144 VSUBS 0.007585f
C498 B.n145 VSUBS 0.007585f
C499 B.n146 VSUBS 0.007585f
C500 B.n147 VSUBS 0.007585f
C501 B.n148 VSUBS 0.007585f
C502 B.n149 VSUBS 0.007585f
C503 B.n150 VSUBS 0.007585f
C504 B.n151 VSUBS 0.007585f
C505 B.n152 VSUBS 0.007585f
C506 B.n153 VSUBS 0.007585f
C507 B.n154 VSUBS 0.007585f
C508 B.n155 VSUBS 0.007585f
C509 B.n156 VSUBS 0.007585f
C510 B.n157 VSUBS 0.007585f
C511 B.n158 VSUBS 0.007585f
C512 B.n159 VSUBS 0.007585f
C513 B.n160 VSUBS 0.007585f
C514 B.n161 VSUBS 0.007585f
C515 B.n162 VSUBS 0.007585f
C516 B.n163 VSUBS 0.007585f
C517 B.n164 VSUBS 0.007585f
C518 B.n165 VSUBS 0.007585f
C519 B.n166 VSUBS 0.007585f
C520 B.n167 VSUBS 0.007585f
C521 B.n168 VSUBS 0.007585f
C522 B.n169 VSUBS 0.007585f
C523 B.n170 VSUBS 0.007585f
C524 B.n171 VSUBS 0.007585f
C525 B.n172 VSUBS 0.007585f
C526 B.n173 VSUBS 0.007585f
C527 B.n174 VSUBS 0.007585f
C528 B.n175 VSUBS 0.007585f
C529 B.n176 VSUBS 0.007585f
C530 B.n177 VSUBS 0.007585f
C531 B.n178 VSUBS 0.007585f
C532 B.n179 VSUBS 0.007585f
C533 B.n180 VSUBS 0.007585f
C534 B.n181 VSUBS 0.007585f
C535 B.n182 VSUBS 0.007585f
C536 B.n183 VSUBS 0.007585f
C537 B.n184 VSUBS 0.007585f
C538 B.n185 VSUBS 0.017051f
C539 B.n186 VSUBS 0.007585f
C540 B.n187 VSUBS 0.007585f
C541 B.n188 VSUBS 0.007585f
C542 B.n189 VSUBS 0.007585f
C543 B.n190 VSUBS 0.007585f
C544 B.n191 VSUBS 0.007585f
C545 B.n192 VSUBS 0.007585f
C546 B.n193 VSUBS 0.007585f
C547 B.n194 VSUBS 0.007585f
C548 B.n195 VSUBS 0.007585f
C549 B.n196 VSUBS 0.007585f
C550 B.n197 VSUBS 0.007585f
C551 B.n198 VSUBS 0.007585f
C552 B.n199 VSUBS 0.007585f
C553 B.n200 VSUBS 0.007585f
C554 B.n201 VSUBS 0.007585f
C555 B.n202 VSUBS 0.007585f
C556 B.n203 VSUBS 0.007585f
C557 B.n204 VSUBS 0.007585f
C558 B.n205 VSUBS 0.007585f
C559 B.n206 VSUBS 0.007585f
C560 B.n207 VSUBS 0.007585f
C561 B.n208 VSUBS 0.007585f
C562 B.n209 VSUBS 0.007585f
C563 B.n210 VSUBS 0.007585f
C564 B.n211 VSUBS 0.007585f
C565 B.n212 VSUBS 0.007585f
C566 B.n213 VSUBS 0.007585f
C567 B.n214 VSUBS 0.007585f
C568 B.n215 VSUBS 0.007585f
C569 B.t10 VSUBS 0.685464f
C570 B.t11 VSUBS 0.713536f
C571 B.t9 VSUBS 3.15535f
C572 B.n216 VSUBS 0.436109f
C573 B.n217 VSUBS 0.081984f
C574 B.n218 VSUBS 0.017574f
C575 B.n219 VSUBS 0.007585f
C576 B.n220 VSUBS 0.007585f
C577 B.n221 VSUBS 0.007585f
C578 B.n222 VSUBS 0.007585f
C579 B.n223 VSUBS 0.007585f
C580 B.t1 VSUBS 0.68549f
C581 B.t2 VSUBS 0.713556f
C582 B.t0 VSUBS 3.15535f
C583 B.n224 VSUBS 0.436089f
C584 B.n225 VSUBS 0.081958f
C585 B.n226 VSUBS 0.007585f
C586 B.n227 VSUBS 0.007585f
C587 B.n228 VSUBS 0.007585f
C588 B.n229 VSUBS 0.007585f
C589 B.n230 VSUBS 0.007585f
C590 B.n231 VSUBS 0.007585f
C591 B.n232 VSUBS 0.007585f
C592 B.n233 VSUBS 0.007585f
C593 B.n234 VSUBS 0.007585f
C594 B.n235 VSUBS 0.007585f
C595 B.n236 VSUBS 0.007585f
C596 B.n237 VSUBS 0.007585f
C597 B.n238 VSUBS 0.007585f
C598 B.n239 VSUBS 0.007585f
C599 B.n240 VSUBS 0.007585f
C600 B.n241 VSUBS 0.007585f
C601 B.n242 VSUBS 0.007585f
C602 B.n243 VSUBS 0.007585f
C603 B.n244 VSUBS 0.007585f
C604 B.n245 VSUBS 0.007585f
C605 B.n246 VSUBS 0.007585f
C606 B.n247 VSUBS 0.007585f
C607 B.n248 VSUBS 0.007585f
C608 B.n249 VSUBS 0.007585f
C609 B.n250 VSUBS 0.007585f
C610 B.n251 VSUBS 0.007585f
C611 B.n252 VSUBS 0.007585f
C612 B.n253 VSUBS 0.007585f
C613 B.n254 VSUBS 0.007585f
C614 B.n255 VSUBS 0.007585f
C615 B.n256 VSUBS 0.017051f
C616 B.n257 VSUBS 0.007585f
C617 B.n258 VSUBS 0.007585f
C618 B.n259 VSUBS 0.007585f
C619 B.n260 VSUBS 0.007585f
C620 B.n261 VSUBS 0.007585f
C621 B.n262 VSUBS 0.007585f
C622 B.n263 VSUBS 0.007585f
C623 B.n264 VSUBS 0.007585f
C624 B.n265 VSUBS 0.007585f
C625 B.n266 VSUBS 0.007585f
C626 B.n267 VSUBS 0.007585f
C627 B.n268 VSUBS 0.007585f
C628 B.n269 VSUBS 0.007585f
C629 B.n270 VSUBS 0.007585f
C630 B.n271 VSUBS 0.007585f
C631 B.n272 VSUBS 0.007585f
C632 B.n273 VSUBS 0.007585f
C633 B.n274 VSUBS 0.007585f
C634 B.n275 VSUBS 0.007585f
C635 B.n276 VSUBS 0.007585f
C636 B.n277 VSUBS 0.007585f
C637 B.n278 VSUBS 0.007585f
C638 B.n279 VSUBS 0.007585f
C639 B.n280 VSUBS 0.007585f
C640 B.n281 VSUBS 0.007585f
C641 B.n282 VSUBS 0.007585f
C642 B.n283 VSUBS 0.007585f
C643 B.n284 VSUBS 0.007585f
C644 B.n285 VSUBS 0.007585f
C645 B.n286 VSUBS 0.007585f
C646 B.n287 VSUBS 0.007585f
C647 B.n288 VSUBS 0.007585f
C648 B.n289 VSUBS 0.007585f
C649 B.n290 VSUBS 0.007585f
C650 B.n291 VSUBS 0.007585f
C651 B.n292 VSUBS 0.007585f
C652 B.n293 VSUBS 0.007585f
C653 B.n294 VSUBS 0.007585f
C654 B.n295 VSUBS 0.007585f
C655 B.n296 VSUBS 0.007585f
C656 B.n297 VSUBS 0.007585f
C657 B.n298 VSUBS 0.007585f
C658 B.n299 VSUBS 0.007585f
C659 B.n300 VSUBS 0.007585f
C660 B.n301 VSUBS 0.007585f
C661 B.n302 VSUBS 0.007585f
C662 B.n303 VSUBS 0.007585f
C663 B.n304 VSUBS 0.007585f
C664 B.n305 VSUBS 0.007585f
C665 B.n306 VSUBS 0.007585f
C666 B.n307 VSUBS 0.007585f
C667 B.n308 VSUBS 0.007585f
C668 B.n309 VSUBS 0.007585f
C669 B.n310 VSUBS 0.007585f
C670 B.n311 VSUBS 0.007585f
C671 B.n312 VSUBS 0.007585f
C672 B.n313 VSUBS 0.007585f
C673 B.n314 VSUBS 0.007585f
C674 B.n315 VSUBS 0.007585f
C675 B.n316 VSUBS 0.007585f
C676 B.n317 VSUBS 0.007585f
C677 B.n318 VSUBS 0.007585f
C678 B.n319 VSUBS 0.007585f
C679 B.n320 VSUBS 0.007585f
C680 B.n321 VSUBS 0.007585f
C681 B.n322 VSUBS 0.007585f
C682 B.n323 VSUBS 0.007585f
C683 B.n324 VSUBS 0.007585f
C684 B.n325 VSUBS 0.007585f
C685 B.n326 VSUBS 0.007585f
C686 B.n327 VSUBS 0.007585f
C687 B.n328 VSUBS 0.007585f
C688 B.n329 VSUBS 0.007585f
C689 B.n330 VSUBS 0.007585f
C690 B.n331 VSUBS 0.007585f
C691 B.n332 VSUBS 0.007585f
C692 B.n333 VSUBS 0.007585f
C693 B.n334 VSUBS 0.007585f
C694 B.n335 VSUBS 0.007585f
C695 B.n336 VSUBS 0.007585f
C696 B.n337 VSUBS 0.007585f
C697 B.n338 VSUBS 0.007585f
C698 B.n339 VSUBS 0.007585f
C699 B.n340 VSUBS 0.007585f
C700 B.n341 VSUBS 0.007585f
C701 B.n342 VSUBS 0.007585f
C702 B.n343 VSUBS 0.007585f
C703 B.n344 VSUBS 0.007585f
C704 B.n345 VSUBS 0.007585f
C705 B.n346 VSUBS 0.007585f
C706 B.n347 VSUBS 0.007585f
C707 B.n348 VSUBS 0.007585f
C708 B.n349 VSUBS 0.007585f
C709 B.n350 VSUBS 0.007585f
C710 B.n351 VSUBS 0.007585f
C711 B.n352 VSUBS 0.007585f
C712 B.n353 VSUBS 0.007585f
C713 B.n354 VSUBS 0.007585f
C714 B.n355 VSUBS 0.007585f
C715 B.n356 VSUBS 0.007585f
C716 B.n357 VSUBS 0.007585f
C717 B.n358 VSUBS 0.007585f
C718 B.n359 VSUBS 0.007585f
C719 B.n360 VSUBS 0.007585f
C720 B.n361 VSUBS 0.007585f
C721 B.n362 VSUBS 0.007585f
C722 B.n363 VSUBS 0.007585f
C723 B.n364 VSUBS 0.007585f
C724 B.n365 VSUBS 0.007585f
C725 B.n366 VSUBS 0.007585f
C726 B.n367 VSUBS 0.007585f
C727 B.n368 VSUBS 0.007585f
C728 B.n369 VSUBS 0.007585f
C729 B.n370 VSUBS 0.007585f
C730 B.n371 VSUBS 0.007585f
C731 B.n372 VSUBS 0.007585f
C732 B.n373 VSUBS 0.007585f
C733 B.n374 VSUBS 0.007585f
C734 B.n375 VSUBS 0.007585f
C735 B.n376 VSUBS 0.007585f
C736 B.n377 VSUBS 0.007585f
C737 B.n378 VSUBS 0.007585f
C738 B.n379 VSUBS 0.007585f
C739 B.n380 VSUBS 0.007585f
C740 B.n381 VSUBS 0.007585f
C741 B.n382 VSUBS 0.007585f
C742 B.n383 VSUBS 0.007585f
C743 B.n384 VSUBS 0.007585f
C744 B.n385 VSUBS 0.007585f
C745 B.n386 VSUBS 0.007585f
C746 B.n387 VSUBS 0.007585f
C747 B.n388 VSUBS 0.007585f
C748 B.n389 VSUBS 0.007585f
C749 B.n390 VSUBS 0.007585f
C750 B.n391 VSUBS 0.007585f
C751 B.n392 VSUBS 0.007585f
C752 B.n393 VSUBS 0.007585f
C753 B.n394 VSUBS 0.007585f
C754 B.n395 VSUBS 0.007585f
C755 B.n396 VSUBS 0.007585f
C756 B.n397 VSUBS 0.007585f
C757 B.n398 VSUBS 0.007585f
C758 B.n399 VSUBS 0.007585f
C759 B.n400 VSUBS 0.007585f
C760 B.n401 VSUBS 0.007585f
C761 B.n402 VSUBS 0.007585f
C762 B.n403 VSUBS 0.017051f
C763 B.n404 VSUBS 0.017528f
C764 B.n405 VSUBS 0.017528f
C765 B.n406 VSUBS 0.007585f
C766 B.n407 VSUBS 0.007585f
C767 B.n408 VSUBS 0.007585f
C768 B.n409 VSUBS 0.007585f
C769 B.n410 VSUBS 0.007585f
C770 B.n411 VSUBS 0.007585f
C771 B.n412 VSUBS 0.007585f
C772 B.n413 VSUBS 0.007585f
C773 B.n414 VSUBS 0.007585f
C774 B.n415 VSUBS 0.007585f
C775 B.n416 VSUBS 0.007585f
C776 B.n417 VSUBS 0.007585f
C777 B.n418 VSUBS 0.007585f
C778 B.n419 VSUBS 0.007585f
C779 B.n420 VSUBS 0.007585f
C780 B.n421 VSUBS 0.007585f
C781 B.n422 VSUBS 0.007585f
C782 B.n423 VSUBS 0.007585f
C783 B.n424 VSUBS 0.007585f
C784 B.n425 VSUBS 0.007585f
C785 B.n426 VSUBS 0.007585f
C786 B.n427 VSUBS 0.007585f
C787 B.n428 VSUBS 0.007585f
C788 B.n429 VSUBS 0.007585f
C789 B.n430 VSUBS 0.007585f
C790 B.n431 VSUBS 0.007585f
C791 B.n432 VSUBS 0.007585f
C792 B.n433 VSUBS 0.007585f
C793 B.n434 VSUBS 0.007585f
C794 B.n435 VSUBS 0.007585f
C795 B.n436 VSUBS 0.007585f
C796 B.n437 VSUBS 0.007585f
C797 B.n438 VSUBS 0.007585f
C798 B.n439 VSUBS 0.007585f
C799 B.n440 VSUBS 0.007585f
C800 B.n441 VSUBS 0.007585f
C801 B.n442 VSUBS 0.007585f
C802 B.n443 VSUBS 0.007585f
C803 B.n444 VSUBS 0.007585f
C804 B.n445 VSUBS 0.007585f
C805 B.n446 VSUBS 0.007585f
C806 B.n447 VSUBS 0.007585f
C807 B.n448 VSUBS 0.007585f
C808 B.n449 VSUBS 0.007585f
C809 B.n450 VSUBS 0.007585f
C810 B.n451 VSUBS 0.007585f
C811 B.n452 VSUBS 0.007585f
C812 B.n453 VSUBS 0.007585f
C813 B.n454 VSUBS 0.007585f
C814 B.n455 VSUBS 0.007585f
C815 B.n456 VSUBS 0.007585f
C816 B.n457 VSUBS 0.007585f
C817 B.n458 VSUBS 0.007585f
C818 B.n459 VSUBS 0.007585f
C819 B.n460 VSUBS 0.007585f
C820 B.n461 VSUBS 0.007585f
C821 B.n462 VSUBS 0.007585f
C822 B.n463 VSUBS 0.007585f
C823 B.n464 VSUBS 0.007585f
C824 B.n465 VSUBS 0.007585f
C825 B.n466 VSUBS 0.007585f
C826 B.n467 VSUBS 0.007585f
C827 B.n468 VSUBS 0.007585f
C828 B.n469 VSUBS 0.007585f
C829 B.n470 VSUBS 0.007585f
C830 B.n471 VSUBS 0.007585f
C831 B.n472 VSUBS 0.007585f
C832 B.n473 VSUBS 0.007585f
C833 B.n474 VSUBS 0.007585f
C834 B.n475 VSUBS 0.007585f
C835 B.n476 VSUBS 0.007585f
C836 B.n477 VSUBS 0.007585f
C837 B.n478 VSUBS 0.007585f
C838 B.n479 VSUBS 0.007585f
C839 B.n480 VSUBS 0.007585f
C840 B.n481 VSUBS 0.007585f
C841 B.n482 VSUBS 0.007585f
C842 B.n483 VSUBS 0.007585f
C843 B.n484 VSUBS 0.007585f
C844 B.n485 VSUBS 0.007585f
C845 B.n486 VSUBS 0.007585f
C846 B.n487 VSUBS 0.007585f
C847 B.n488 VSUBS 0.007585f
C848 B.n489 VSUBS 0.007585f
C849 B.n490 VSUBS 0.007585f
C850 B.n491 VSUBS 0.007585f
C851 B.n492 VSUBS 0.007585f
C852 B.n493 VSUBS 0.007585f
C853 B.n494 VSUBS 0.007585f
C854 B.n495 VSUBS 0.007139f
C855 B.n496 VSUBS 0.017574f
C856 B.n497 VSUBS 0.004239f
C857 B.n498 VSUBS 0.007585f
C858 B.n499 VSUBS 0.007585f
C859 B.n500 VSUBS 0.007585f
C860 B.n501 VSUBS 0.007585f
C861 B.n502 VSUBS 0.007585f
C862 B.n503 VSUBS 0.007585f
C863 B.n504 VSUBS 0.007585f
C864 B.n505 VSUBS 0.007585f
C865 B.n506 VSUBS 0.007585f
C866 B.n507 VSUBS 0.007585f
C867 B.n508 VSUBS 0.007585f
C868 B.n509 VSUBS 0.007585f
C869 B.n510 VSUBS 0.004239f
C870 B.n511 VSUBS 0.007585f
C871 B.n512 VSUBS 0.007585f
C872 B.n513 VSUBS 0.007139f
C873 B.n514 VSUBS 0.007585f
C874 B.n515 VSUBS 0.007585f
C875 B.n516 VSUBS 0.007585f
C876 B.n517 VSUBS 0.007585f
C877 B.n518 VSUBS 0.007585f
C878 B.n519 VSUBS 0.007585f
C879 B.n520 VSUBS 0.007585f
C880 B.n521 VSUBS 0.007585f
C881 B.n522 VSUBS 0.007585f
C882 B.n523 VSUBS 0.007585f
C883 B.n524 VSUBS 0.007585f
C884 B.n525 VSUBS 0.007585f
C885 B.n526 VSUBS 0.007585f
C886 B.n527 VSUBS 0.007585f
C887 B.n528 VSUBS 0.007585f
C888 B.n529 VSUBS 0.007585f
C889 B.n530 VSUBS 0.007585f
C890 B.n531 VSUBS 0.007585f
C891 B.n532 VSUBS 0.007585f
C892 B.n533 VSUBS 0.007585f
C893 B.n534 VSUBS 0.007585f
C894 B.n535 VSUBS 0.007585f
C895 B.n536 VSUBS 0.007585f
C896 B.n537 VSUBS 0.007585f
C897 B.n538 VSUBS 0.007585f
C898 B.n539 VSUBS 0.007585f
C899 B.n540 VSUBS 0.007585f
C900 B.n541 VSUBS 0.007585f
C901 B.n542 VSUBS 0.007585f
C902 B.n543 VSUBS 0.007585f
C903 B.n544 VSUBS 0.007585f
C904 B.n545 VSUBS 0.007585f
C905 B.n546 VSUBS 0.007585f
C906 B.n547 VSUBS 0.007585f
C907 B.n548 VSUBS 0.007585f
C908 B.n549 VSUBS 0.007585f
C909 B.n550 VSUBS 0.007585f
C910 B.n551 VSUBS 0.007585f
C911 B.n552 VSUBS 0.007585f
C912 B.n553 VSUBS 0.007585f
C913 B.n554 VSUBS 0.007585f
C914 B.n555 VSUBS 0.007585f
C915 B.n556 VSUBS 0.007585f
C916 B.n557 VSUBS 0.007585f
C917 B.n558 VSUBS 0.007585f
C918 B.n559 VSUBS 0.007585f
C919 B.n560 VSUBS 0.007585f
C920 B.n561 VSUBS 0.007585f
C921 B.n562 VSUBS 0.007585f
C922 B.n563 VSUBS 0.007585f
C923 B.n564 VSUBS 0.007585f
C924 B.n565 VSUBS 0.007585f
C925 B.n566 VSUBS 0.007585f
C926 B.n567 VSUBS 0.007585f
C927 B.n568 VSUBS 0.007585f
C928 B.n569 VSUBS 0.007585f
C929 B.n570 VSUBS 0.007585f
C930 B.n571 VSUBS 0.007585f
C931 B.n572 VSUBS 0.007585f
C932 B.n573 VSUBS 0.007585f
C933 B.n574 VSUBS 0.007585f
C934 B.n575 VSUBS 0.007585f
C935 B.n576 VSUBS 0.007585f
C936 B.n577 VSUBS 0.007585f
C937 B.n578 VSUBS 0.007585f
C938 B.n579 VSUBS 0.007585f
C939 B.n580 VSUBS 0.007585f
C940 B.n581 VSUBS 0.007585f
C941 B.n582 VSUBS 0.007585f
C942 B.n583 VSUBS 0.007585f
C943 B.n584 VSUBS 0.007585f
C944 B.n585 VSUBS 0.007585f
C945 B.n586 VSUBS 0.007585f
C946 B.n587 VSUBS 0.007585f
C947 B.n588 VSUBS 0.007585f
C948 B.n589 VSUBS 0.007585f
C949 B.n590 VSUBS 0.007585f
C950 B.n591 VSUBS 0.007585f
C951 B.n592 VSUBS 0.007585f
C952 B.n593 VSUBS 0.007585f
C953 B.n594 VSUBS 0.007585f
C954 B.n595 VSUBS 0.007585f
C955 B.n596 VSUBS 0.007585f
C956 B.n597 VSUBS 0.007585f
C957 B.n598 VSUBS 0.007585f
C958 B.n599 VSUBS 0.007585f
C959 B.n600 VSUBS 0.007585f
C960 B.n601 VSUBS 0.007585f
C961 B.n602 VSUBS 0.017528f
C962 B.n603 VSUBS 0.017528f
C963 B.n604 VSUBS 0.017051f
C964 B.n605 VSUBS 0.007585f
C965 B.n606 VSUBS 0.007585f
C966 B.n607 VSUBS 0.007585f
C967 B.n608 VSUBS 0.007585f
C968 B.n609 VSUBS 0.007585f
C969 B.n610 VSUBS 0.007585f
C970 B.n611 VSUBS 0.007585f
C971 B.n612 VSUBS 0.007585f
C972 B.n613 VSUBS 0.007585f
C973 B.n614 VSUBS 0.007585f
C974 B.n615 VSUBS 0.007585f
C975 B.n616 VSUBS 0.007585f
C976 B.n617 VSUBS 0.007585f
C977 B.n618 VSUBS 0.007585f
C978 B.n619 VSUBS 0.007585f
C979 B.n620 VSUBS 0.007585f
C980 B.n621 VSUBS 0.007585f
C981 B.n622 VSUBS 0.007585f
C982 B.n623 VSUBS 0.007585f
C983 B.n624 VSUBS 0.007585f
C984 B.n625 VSUBS 0.007585f
C985 B.n626 VSUBS 0.007585f
C986 B.n627 VSUBS 0.007585f
C987 B.n628 VSUBS 0.007585f
C988 B.n629 VSUBS 0.007585f
C989 B.n630 VSUBS 0.007585f
C990 B.n631 VSUBS 0.007585f
C991 B.n632 VSUBS 0.007585f
C992 B.n633 VSUBS 0.007585f
C993 B.n634 VSUBS 0.007585f
C994 B.n635 VSUBS 0.007585f
C995 B.n636 VSUBS 0.007585f
C996 B.n637 VSUBS 0.007585f
C997 B.n638 VSUBS 0.007585f
C998 B.n639 VSUBS 0.007585f
C999 B.n640 VSUBS 0.007585f
C1000 B.n641 VSUBS 0.007585f
C1001 B.n642 VSUBS 0.007585f
C1002 B.n643 VSUBS 0.007585f
C1003 B.n644 VSUBS 0.007585f
C1004 B.n645 VSUBS 0.007585f
C1005 B.n646 VSUBS 0.007585f
C1006 B.n647 VSUBS 0.007585f
C1007 B.n648 VSUBS 0.007585f
C1008 B.n649 VSUBS 0.007585f
C1009 B.n650 VSUBS 0.007585f
C1010 B.n651 VSUBS 0.007585f
C1011 B.n652 VSUBS 0.007585f
C1012 B.n653 VSUBS 0.007585f
C1013 B.n654 VSUBS 0.007585f
C1014 B.n655 VSUBS 0.007585f
C1015 B.n656 VSUBS 0.007585f
C1016 B.n657 VSUBS 0.007585f
C1017 B.n658 VSUBS 0.007585f
C1018 B.n659 VSUBS 0.007585f
C1019 B.n660 VSUBS 0.007585f
C1020 B.n661 VSUBS 0.007585f
C1021 B.n662 VSUBS 0.007585f
C1022 B.n663 VSUBS 0.007585f
C1023 B.n664 VSUBS 0.007585f
C1024 B.n665 VSUBS 0.007585f
C1025 B.n666 VSUBS 0.007585f
C1026 B.n667 VSUBS 0.007585f
C1027 B.n668 VSUBS 0.007585f
C1028 B.n669 VSUBS 0.007585f
C1029 B.n670 VSUBS 0.007585f
C1030 B.n671 VSUBS 0.007585f
C1031 B.n672 VSUBS 0.007585f
C1032 B.n673 VSUBS 0.007585f
C1033 B.n674 VSUBS 0.007585f
C1034 B.n675 VSUBS 0.007585f
C1035 B.n676 VSUBS 0.007585f
C1036 B.n677 VSUBS 0.007585f
C1037 B.n678 VSUBS 0.007585f
C1038 B.n679 VSUBS 0.007585f
C1039 B.n680 VSUBS 0.007585f
C1040 B.n681 VSUBS 0.007585f
C1041 B.n682 VSUBS 0.007585f
C1042 B.n683 VSUBS 0.007585f
C1043 B.n684 VSUBS 0.007585f
C1044 B.n685 VSUBS 0.007585f
C1045 B.n686 VSUBS 0.007585f
C1046 B.n687 VSUBS 0.007585f
C1047 B.n688 VSUBS 0.007585f
C1048 B.n689 VSUBS 0.007585f
C1049 B.n690 VSUBS 0.007585f
C1050 B.n691 VSUBS 0.007585f
C1051 B.n692 VSUBS 0.007585f
C1052 B.n693 VSUBS 0.007585f
C1053 B.n694 VSUBS 0.007585f
C1054 B.n695 VSUBS 0.007585f
C1055 B.n696 VSUBS 0.007585f
C1056 B.n697 VSUBS 0.007585f
C1057 B.n698 VSUBS 0.007585f
C1058 B.n699 VSUBS 0.007585f
C1059 B.n700 VSUBS 0.007585f
C1060 B.n701 VSUBS 0.007585f
C1061 B.n702 VSUBS 0.007585f
C1062 B.n703 VSUBS 0.007585f
C1063 B.n704 VSUBS 0.007585f
C1064 B.n705 VSUBS 0.007585f
C1065 B.n706 VSUBS 0.007585f
C1066 B.n707 VSUBS 0.007585f
C1067 B.n708 VSUBS 0.007585f
C1068 B.n709 VSUBS 0.007585f
C1069 B.n710 VSUBS 0.007585f
C1070 B.n711 VSUBS 0.007585f
C1071 B.n712 VSUBS 0.007585f
C1072 B.n713 VSUBS 0.007585f
C1073 B.n714 VSUBS 0.007585f
C1074 B.n715 VSUBS 0.007585f
C1075 B.n716 VSUBS 0.007585f
C1076 B.n717 VSUBS 0.007585f
C1077 B.n718 VSUBS 0.007585f
C1078 B.n719 VSUBS 0.007585f
C1079 B.n720 VSUBS 0.007585f
C1080 B.n721 VSUBS 0.007585f
C1081 B.n722 VSUBS 0.007585f
C1082 B.n723 VSUBS 0.007585f
C1083 B.n724 VSUBS 0.007585f
C1084 B.n725 VSUBS 0.007585f
C1085 B.n726 VSUBS 0.007585f
C1086 B.n727 VSUBS 0.007585f
C1087 B.n728 VSUBS 0.007585f
C1088 B.n729 VSUBS 0.007585f
C1089 B.n730 VSUBS 0.007585f
C1090 B.n731 VSUBS 0.007585f
C1091 B.n732 VSUBS 0.007585f
C1092 B.n733 VSUBS 0.007585f
C1093 B.n734 VSUBS 0.007585f
C1094 B.n735 VSUBS 0.007585f
C1095 B.n736 VSUBS 0.007585f
C1096 B.n737 VSUBS 0.007585f
C1097 B.n738 VSUBS 0.007585f
C1098 B.n739 VSUBS 0.007585f
C1099 B.n740 VSUBS 0.007585f
C1100 B.n741 VSUBS 0.007585f
C1101 B.n742 VSUBS 0.007585f
C1102 B.n743 VSUBS 0.007585f
C1103 B.n744 VSUBS 0.007585f
C1104 B.n745 VSUBS 0.007585f
C1105 B.n746 VSUBS 0.007585f
C1106 B.n747 VSUBS 0.007585f
C1107 B.n748 VSUBS 0.007585f
C1108 B.n749 VSUBS 0.007585f
C1109 B.n750 VSUBS 0.007585f
C1110 B.n751 VSUBS 0.007585f
C1111 B.n752 VSUBS 0.007585f
C1112 B.n753 VSUBS 0.007585f
C1113 B.n754 VSUBS 0.007585f
C1114 B.n755 VSUBS 0.007585f
C1115 B.n756 VSUBS 0.007585f
C1116 B.n757 VSUBS 0.007585f
C1117 B.n758 VSUBS 0.007585f
C1118 B.n759 VSUBS 0.007585f
C1119 B.n760 VSUBS 0.007585f
C1120 B.n761 VSUBS 0.007585f
C1121 B.n762 VSUBS 0.007585f
C1122 B.n763 VSUBS 0.007585f
C1123 B.n764 VSUBS 0.007585f
C1124 B.n765 VSUBS 0.007585f
C1125 B.n766 VSUBS 0.007585f
C1126 B.n767 VSUBS 0.007585f
C1127 B.n768 VSUBS 0.007585f
C1128 B.n769 VSUBS 0.007585f
C1129 B.n770 VSUBS 0.007585f
C1130 B.n771 VSUBS 0.007585f
C1131 B.n772 VSUBS 0.007585f
C1132 B.n773 VSUBS 0.007585f
C1133 B.n774 VSUBS 0.007585f
C1134 B.n775 VSUBS 0.007585f
C1135 B.n776 VSUBS 0.007585f
C1136 B.n777 VSUBS 0.007585f
C1137 B.n778 VSUBS 0.007585f
C1138 B.n779 VSUBS 0.007585f
C1139 B.n780 VSUBS 0.007585f
C1140 B.n781 VSUBS 0.007585f
C1141 B.n782 VSUBS 0.007585f
C1142 B.n783 VSUBS 0.007585f
C1143 B.n784 VSUBS 0.007585f
C1144 B.n785 VSUBS 0.007585f
C1145 B.n786 VSUBS 0.007585f
C1146 B.n787 VSUBS 0.007585f
C1147 B.n788 VSUBS 0.007585f
C1148 B.n789 VSUBS 0.007585f
C1149 B.n790 VSUBS 0.007585f
C1150 B.n791 VSUBS 0.007585f
C1151 B.n792 VSUBS 0.007585f
C1152 B.n793 VSUBS 0.007585f
C1153 B.n794 VSUBS 0.007585f
C1154 B.n795 VSUBS 0.007585f
C1155 B.n796 VSUBS 0.007585f
C1156 B.n797 VSUBS 0.007585f
C1157 B.n798 VSUBS 0.007585f
C1158 B.n799 VSUBS 0.007585f
C1159 B.n800 VSUBS 0.007585f
C1160 B.n801 VSUBS 0.007585f
C1161 B.n802 VSUBS 0.007585f
C1162 B.n803 VSUBS 0.007585f
C1163 B.n804 VSUBS 0.007585f
C1164 B.n805 VSUBS 0.007585f
C1165 B.n806 VSUBS 0.007585f
C1166 B.n807 VSUBS 0.007585f
C1167 B.n808 VSUBS 0.007585f
C1168 B.n809 VSUBS 0.007585f
C1169 B.n810 VSUBS 0.007585f
C1170 B.n811 VSUBS 0.007585f
C1171 B.n812 VSUBS 0.007585f
C1172 B.n813 VSUBS 0.007585f
C1173 B.n814 VSUBS 0.007585f
C1174 B.n815 VSUBS 0.007585f
C1175 B.n816 VSUBS 0.007585f
C1176 B.n817 VSUBS 0.007585f
C1177 B.n818 VSUBS 0.007585f
C1178 B.n819 VSUBS 0.007585f
C1179 B.n820 VSUBS 0.007585f
C1180 B.n821 VSUBS 0.007585f
C1181 B.n822 VSUBS 0.007585f
C1182 B.n823 VSUBS 0.007585f
C1183 B.n824 VSUBS 0.007585f
C1184 B.n825 VSUBS 0.007585f
C1185 B.n826 VSUBS 0.007585f
C1186 B.n827 VSUBS 0.007585f
C1187 B.n828 VSUBS 0.007585f
C1188 B.n829 VSUBS 0.017051f
C1189 B.n830 VSUBS 0.017528f
C1190 B.n831 VSUBS 0.016595f
C1191 B.n832 VSUBS 0.007585f
C1192 B.n833 VSUBS 0.007585f
C1193 B.n834 VSUBS 0.007585f
C1194 B.n835 VSUBS 0.007585f
C1195 B.n836 VSUBS 0.007585f
C1196 B.n837 VSUBS 0.007585f
C1197 B.n838 VSUBS 0.007585f
C1198 B.n839 VSUBS 0.007585f
C1199 B.n840 VSUBS 0.007585f
C1200 B.n841 VSUBS 0.007585f
C1201 B.n842 VSUBS 0.007585f
C1202 B.n843 VSUBS 0.007585f
C1203 B.n844 VSUBS 0.007585f
C1204 B.n845 VSUBS 0.007585f
C1205 B.n846 VSUBS 0.007585f
C1206 B.n847 VSUBS 0.007585f
C1207 B.n848 VSUBS 0.007585f
C1208 B.n849 VSUBS 0.007585f
C1209 B.n850 VSUBS 0.007585f
C1210 B.n851 VSUBS 0.007585f
C1211 B.n852 VSUBS 0.007585f
C1212 B.n853 VSUBS 0.007585f
C1213 B.n854 VSUBS 0.007585f
C1214 B.n855 VSUBS 0.007585f
C1215 B.n856 VSUBS 0.007585f
C1216 B.n857 VSUBS 0.007585f
C1217 B.n858 VSUBS 0.007585f
C1218 B.n859 VSUBS 0.007585f
C1219 B.n860 VSUBS 0.007585f
C1220 B.n861 VSUBS 0.007585f
C1221 B.n862 VSUBS 0.007585f
C1222 B.n863 VSUBS 0.007585f
C1223 B.n864 VSUBS 0.007585f
C1224 B.n865 VSUBS 0.007585f
C1225 B.n866 VSUBS 0.007585f
C1226 B.n867 VSUBS 0.007585f
C1227 B.n868 VSUBS 0.007585f
C1228 B.n869 VSUBS 0.007585f
C1229 B.n870 VSUBS 0.007585f
C1230 B.n871 VSUBS 0.007585f
C1231 B.n872 VSUBS 0.007585f
C1232 B.n873 VSUBS 0.007585f
C1233 B.n874 VSUBS 0.007585f
C1234 B.n875 VSUBS 0.007585f
C1235 B.n876 VSUBS 0.007585f
C1236 B.n877 VSUBS 0.007585f
C1237 B.n878 VSUBS 0.007585f
C1238 B.n879 VSUBS 0.007585f
C1239 B.n880 VSUBS 0.007585f
C1240 B.n881 VSUBS 0.007585f
C1241 B.n882 VSUBS 0.007585f
C1242 B.n883 VSUBS 0.007585f
C1243 B.n884 VSUBS 0.007585f
C1244 B.n885 VSUBS 0.007585f
C1245 B.n886 VSUBS 0.007585f
C1246 B.n887 VSUBS 0.007585f
C1247 B.n888 VSUBS 0.007585f
C1248 B.n889 VSUBS 0.007585f
C1249 B.n890 VSUBS 0.007585f
C1250 B.n891 VSUBS 0.007585f
C1251 B.n892 VSUBS 0.007585f
C1252 B.n893 VSUBS 0.007585f
C1253 B.n894 VSUBS 0.007585f
C1254 B.n895 VSUBS 0.007585f
C1255 B.n896 VSUBS 0.007585f
C1256 B.n897 VSUBS 0.007585f
C1257 B.n898 VSUBS 0.007585f
C1258 B.n899 VSUBS 0.007585f
C1259 B.n900 VSUBS 0.007585f
C1260 B.n901 VSUBS 0.007585f
C1261 B.n902 VSUBS 0.007585f
C1262 B.n903 VSUBS 0.007585f
C1263 B.n904 VSUBS 0.007585f
C1264 B.n905 VSUBS 0.007585f
C1265 B.n906 VSUBS 0.007585f
C1266 B.n907 VSUBS 0.007585f
C1267 B.n908 VSUBS 0.007585f
C1268 B.n909 VSUBS 0.007585f
C1269 B.n910 VSUBS 0.007585f
C1270 B.n911 VSUBS 0.007585f
C1271 B.n912 VSUBS 0.007585f
C1272 B.n913 VSUBS 0.007585f
C1273 B.n914 VSUBS 0.007585f
C1274 B.n915 VSUBS 0.007585f
C1275 B.n916 VSUBS 0.007585f
C1276 B.n917 VSUBS 0.007585f
C1277 B.n918 VSUBS 0.007585f
C1278 B.n919 VSUBS 0.007585f
C1279 B.n920 VSUBS 0.007585f
C1280 B.n921 VSUBS 0.007139f
C1281 B.n922 VSUBS 0.017574f
C1282 B.n923 VSUBS 0.004239f
C1283 B.n924 VSUBS 0.007585f
C1284 B.n925 VSUBS 0.007585f
C1285 B.n926 VSUBS 0.007585f
C1286 B.n927 VSUBS 0.007585f
C1287 B.n928 VSUBS 0.007585f
C1288 B.n929 VSUBS 0.007585f
C1289 B.n930 VSUBS 0.007585f
C1290 B.n931 VSUBS 0.007585f
C1291 B.n932 VSUBS 0.007585f
C1292 B.n933 VSUBS 0.007585f
C1293 B.n934 VSUBS 0.007585f
C1294 B.n935 VSUBS 0.007585f
C1295 B.n936 VSUBS 0.004239f
C1296 B.n937 VSUBS 0.007585f
C1297 B.n938 VSUBS 0.007585f
C1298 B.n939 VSUBS 0.007139f
C1299 B.n940 VSUBS 0.007585f
C1300 B.n941 VSUBS 0.007585f
C1301 B.n942 VSUBS 0.007585f
C1302 B.n943 VSUBS 0.007585f
C1303 B.n944 VSUBS 0.007585f
C1304 B.n945 VSUBS 0.007585f
C1305 B.n946 VSUBS 0.007585f
C1306 B.n947 VSUBS 0.007585f
C1307 B.n948 VSUBS 0.007585f
C1308 B.n949 VSUBS 0.007585f
C1309 B.n950 VSUBS 0.007585f
C1310 B.n951 VSUBS 0.007585f
C1311 B.n952 VSUBS 0.007585f
C1312 B.n953 VSUBS 0.007585f
C1313 B.n954 VSUBS 0.007585f
C1314 B.n955 VSUBS 0.007585f
C1315 B.n956 VSUBS 0.007585f
C1316 B.n957 VSUBS 0.007585f
C1317 B.n958 VSUBS 0.007585f
C1318 B.n959 VSUBS 0.007585f
C1319 B.n960 VSUBS 0.007585f
C1320 B.n961 VSUBS 0.007585f
C1321 B.n962 VSUBS 0.007585f
C1322 B.n963 VSUBS 0.007585f
C1323 B.n964 VSUBS 0.007585f
C1324 B.n965 VSUBS 0.007585f
C1325 B.n966 VSUBS 0.007585f
C1326 B.n967 VSUBS 0.007585f
C1327 B.n968 VSUBS 0.007585f
C1328 B.n969 VSUBS 0.007585f
C1329 B.n970 VSUBS 0.007585f
C1330 B.n971 VSUBS 0.007585f
C1331 B.n972 VSUBS 0.007585f
C1332 B.n973 VSUBS 0.007585f
C1333 B.n974 VSUBS 0.007585f
C1334 B.n975 VSUBS 0.007585f
C1335 B.n976 VSUBS 0.007585f
C1336 B.n977 VSUBS 0.007585f
C1337 B.n978 VSUBS 0.007585f
C1338 B.n979 VSUBS 0.007585f
C1339 B.n980 VSUBS 0.007585f
C1340 B.n981 VSUBS 0.007585f
C1341 B.n982 VSUBS 0.007585f
C1342 B.n983 VSUBS 0.007585f
C1343 B.n984 VSUBS 0.007585f
C1344 B.n985 VSUBS 0.007585f
C1345 B.n986 VSUBS 0.007585f
C1346 B.n987 VSUBS 0.007585f
C1347 B.n988 VSUBS 0.007585f
C1348 B.n989 VSUBS 0.007585f
C1349 B.n990 VSUBS 0.007585f
C1350 B.n991 VSUBS 0.007585f
C1351 B.n992 VSUBS 0.007585f
C1352 B.n993 VSUBS 0.007585f
C1353 B.n994 VSUBS 0.007585f
C1354 B.n995 VSUBS 0.007585f
C1355 B.n996 VSUBS 0.007585f
C1356 B.n997 VSUBS 0.007585f
C1357 B.n998 VSUBS 0.007585f
C1358 B.n999 VSUBS 0.007585f
C1359 B.n1000 VSUBS 0.007585f
C1360 B.n1001 VSUBS 0.007585f
C1361 B.n1002 VSUBS 0.007585f
C1362 B.n1003 VSUBS 0.007585f
C1363 B.n1004 VSUBS 0.007585f
C1364 B.n1005 VSUBS 0.007585f
C1365 B.n1006 VSUBS 0.007585f
C1366 B.n1007 VSUBS 0.007585f
C1367 B.n1008 VSUBS 0.007585f
C1368 B.n1009 VSUBS 0.007585f
C1369 B.n1010 VSUBS 0.007585f
C1370 B.n1011 VSUBS 0.007585f
C1371 B.n1012 VSUBS 0.007585f
C1372 B.n1013 VSUBS 0.007585f
C1373 B.n1014 VSUBS 0.007585f
C1374 B.n1015 VSUBS 0.007585f
C1375 B.n1016 VSUBS 0.007585f
C1376 B.n1017 VSUBS 0.007585f
C1377 B.n1018 VSUBS 0.007585f
C1378 B.n1019 VSUBS 0.007585f
C1379 B.n1020 VSUBS 0.007585f
C1380 B.n1021 VSUBS 0.007585f
C1381 B.n1022 VSUBS 0.007585f
C1382 B.n1023 VSUBS 0.007585f
C1383 B.n1024 VSUBS 0.007585f
C1384 B.n1025 VSUBS 0.007585f
C1385 B.n1026 VSUBS 0.007585f
C1386 B.n1027 VSUBS 0.007585f
C1387 B.n1028 VSUBS 0.017528f
C1388 B.n1029 VSUBS 0.017528f
C1389 B.n1030 VSUBS 0.017051f
C1390 B.n1031 VSUBS 0.007585f
C1391 B.n1032 VSUBS 0.007585f
C1392 B.n1033 VSUBS 0.007585f
C1393 B.n1034 VSUBS 0.007585f
C1394 B.n1035 VSUBS 0.007585f
C1395 B.n1036 VSUBS 0.007585f
C1396 B.n1037 VSUBS 0.007585f
C1397 B.n1038 VSUBS 0.007585f
C1398 B.n1039 VSUBS 0.007585f
C1399 B.n1040 VSUBS 0.007585f
C1400 B.n1041 VSUBS 0.007585f
C1401 B.n1042 VSUBS 0.007585f
C1402 B.n1043 VSUBS 0.007585f
C1403 B.n1044 VSUBS 0.007585f
C1404 B.n1045 VSUBS 0.007585f
C1405 B.n1046 VSUBS 0.007585f
C1406 B.n1047 VSUBS 0.007585f
C1407 B.n1048 VSUBS 0.007585f
C1408 B.n1049 VSUBS 0.007585f
C1409 B.n1050 VSUBS 0.007585f
C1410 B.n1051 VSUBS 0.007585f
C1411 B.n1052 VSUBS 0.007585f
C1412 B.n1053 VSUBS 0.007585f
C1413 B.n1054 VSUBS 0.007585f
C1414 B.n1055 VSUBS 0.007585f
C1415 B.n1056 VSUBS 0.007585f
C1416 B.n1057 VSUBS 0.007585f
C1417 B.n1058 VSUBS 0.007585f
C1418 B.n1059 VSUBS 0.007585f
C1419 B.n1060 VSUBS 0.007585f
C1420 B.n1061 VSUBS 0.007585f
C1421 B.n1062 VSUBS 0.007585f
C1422 B.n1063 VSUBS 0.007585f
C1423 B.n1064 VSUBS 0.007585f
C1424 B.n1065 VSUBS 0.007585f
C1425 B.n1066 VSUBS 0.007585f
C1426 B.n1067 VSUBS 0.007585f
C1427 B.n1068 VSUBS 0.007585f
C1428 B.n1069 VSUBS 0.007585f
C1429 B.n1070 VSUBS 0.007585f
C1430 B.n1071 VSUBS 0.007585f
C1431 B.n1072 VSUBS 0.007585f
C1432 B.n1073 VSUBS 0.007585f
C1433 B.n1074 VSUBS 0.007585f
C1434 B.n1075 VSUBS 0.007585f
C1435 B.n1076 VSUBS 0.007585f
C1436 B.n1077 VSUBS 0.007585f
C1437 B.n1078 VSUBS 0.007585f
C1438 B.n1079 VSUBS 0.007585f
C1439 B.n1080 VSUBS 0.007585f
C1440 B.n1081 VSUBS 0.007585f
C1441 B.n1082 VSUBS 0.007585f
C1442 B.n1083 VSUBS 0.007585f
C1443 B.n1084 VSUBS 0.007585f
C1444 B.n1085 VSUBS 0.007585f
C1445 B.n1086 VSUBS 0.007585f
C1446 B.n1087 VSUBS 0.007585f
C1447 B.n1088 VSUBS 0.007585f
C1448 B.n1089 VSUBS 0.007585f
C1449 B.n1090 VSUBS 0.007585f
C1450 B.n1091 VSUBS 0.007585f
C1451 B.n1092 VSUBS 0.007585f
C1452 B.n1093 VSUBS 0.007585f
C1453 B.n1094 VSUBS 0.007585f
C1454 B.n1095 VSUBS 0.007585f
C1455 B.n1096 VSUBS 0.007585f
C1456 B.n1097 VSUBS 0.007585f
C1457 B.n1098 VSUBS 0.007585f
C1458 B.n1099 VSUBS 0.007585f
C1459 B.n1100 VSUBS 0.007585f
C1460 B.n1101 VSUBS 0.007585f
C1461 B.n1102 VSUBS 0.007585f
C1462 B.n1103 VSUBS 0.007585f
C1463 B.n1104 VSUBS 0.007585f
C1464 B.n1105 VSUBS 0.007585f
C1465 B.n1106 VSUBS 0.007585f
C1466 B.n1107 VSUBS 0.007585f
C1467 B.n1108 VSUBS 0.007585f
C1468 B.n1109 VSUBS 0.007585f
C1469 B.n1110 VSUBS 0.007585f
C1470 B.n1111 VSUBS 0.007585f
C1471 B.n1112 VSUBS 0.007585f
C1472 B.n1113 VSUBS 0.007585f
C1473 B.n1114 VSUBS 0.007585f
C1474 B.n1115 VSUBS 0.007585f
C1475 B.n1116 VSUBS 0.007585f
C1476 B.n1117 VSUBS 0.007585f
C1477 B.n1118 VSUBS 0.007585f
C1478 B.n1119 VSUBS 0.007585f
C1479 B.n1120 VSUBS 0.007585f
C1480 B.n1121 VSUBS 0.007585f
C1481 B.n1122 VSUBS 0.007585f
C1482 B.n1123 VSUBS 0.007585f
C1483 B.n1124 VSUBS 0.007585f
C1484 B.n1125 VSUBS 0.007585f
C1485 B.n1126 VSUBS 0.007585f
C1486 B.n1127 VSUBS 0.007585f
C1487 B.n1128 VSUBS 0.007585f
C1488 B.n1129 VSUBS 0.007585f
C1489 B.n1130 VSUBS 0.007585f
C1490 B.n1131 VSUBS 0.007585f
C1491 B.n1132 VSUBS 0.007585f
C1492 B.n1133 VSUBS 0.007585f
C1493 B.n1134 VSUBS 0.007585f
C1494 B.n1135 VSUBS 0.007585f
C1495 B.n1136 VSUBS 0.007585f
C1496 B.n1137 VSUBS 0.007585f
C1497 B.n1138 VSUBS 0.007585f
C1498 B.n1139 VSUBS 0.007585f
C1499 B.n1140 VSUBS 0.007585f
C1500 B.n1141 VSUBS 0.007585f
C1501 B.n1142 VSUBS 0.007585f
C1502 B.n1143 VSUBS 0.017175f
.ends

