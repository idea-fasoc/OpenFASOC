* NGSPICE file created from diff_pair_sample_0328.ext - technology: sky130A

.subckt diff_pair_sample_0328 VTAIL VN VP B VDD2 VDD1
X0 B.t17 B.t15 B.t16 B.t5 sky130_fd_pr__nfet_01v8 ad=6.6066 pd=34.66 as=0 ps=0 w=16.94 l=1.49
X1 VTAIL.t7 VN.t0 VDD2.t2 B.t0 sky130_fd_pr__nfet_01v8 ad=6.6066 pd=34.66 as=2.7951 ps=17.27 w=16.94 l=1.49
X2 VTAIL.t1 VP.t0 VDD1.t3 B.t1 sky130_fd_pr__nfet_01v8 ad=6.6066 pd=34.66 as=2.7951 ps=17.27 w=16.94 l=1.49
X3 VTAIL.t6 VN.t1 VDD2.t3 B.t1 sky130_fd_pr__nfet_01v8 ad=6.6066 pd=34.66 as=2.7951 ps=17.27 w=16.94 l=1.49
X4 B.t14 B.t12 B.t13 B.t9 sky130_fd_pr__nfet_01v8 ad=6.6066 pd=34.66 as=0 ps=0 w=16.94 l=1.49
X5 VDD1.t2 VP.t1 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=2.7951 pd=17.27 as=6.6066 ps=34.66 w=16.94 l=1.49
X6 VDD2.t1 VN.t2 VTAIL.t5 B.t3 sky130_fd_pr__nfet_01v8 ad=2.7951 pd=17.27 as=6.6066 ps=34.66 w=16.94 l=1.49
X7 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=6.6066 pd=34.66 as=0 ps=0 w=16.94 l=1.49
X8 VDD2.t0 VN.t3 VTAIL.t4 B.t2 sky130_fd_pr__nfet_01v8 ad=2.7951 pd=17.27 as=6.6066 ps=34.66 w=16.94 l=1.49
X9 B.t7 B.t4 B.t6 B.t5 sky130_fd_pr__nfet_01v8 ad=6.6066 pd=34.66 as=0 ps=0 w=16.94 l=1.49
X10 VDD1.t1 VP.t2 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=2.7951 pd=17.27 as=6.6066 ps=34.66 w=16.94 l=1.49
X11 VTAIL.t0 VP.t3 VDD1.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=6.6066 pd=34.66 as=2.7951 ps=17.27 w=16.94 l=1.49
R0 B.n814 B.n813 585
R1 B.n353 B.n108 585
R2 B.n352 B.n351 585
R3 B.n350 B.n349 585
R4 B.n348 B.n347 585
R5 B.n346 B.n345 585
R6 B.n344 B.n343 585
R7 B.n342 B.n341 585
R8 B.n340 B.n339 585
R9 B.n338 B.n337 585
R10 B.n336 B.n335 585
R11 B.n334 B.n333 585
R12 B.n332 B.n331 585
R13 B.n330 B.n329 585
R14 B.n328 B.n327 585
R15 B.n326 B.n325 585
R16 B.n324 B.n323 585
R17 B.n322 B.n321 585
R18 B.n320 B.n319 585
R19 B.n318 B.n317 585
R20 B.n316 B.n315 585
R21 B.n314 B.n313 585
R22 B.n312 B.n311 585
R23 B.n310 B.n309 585
R24 B.n308 B.n307 585
R25 B.n306 B.n305 585
R26 B.n304 B.n303 585
R27 B.n302 B.n301 585
R28 B.n300 B.n299 585
R29 B.n298 B.n297 585
R30 B.n296 B.n295 585
R31 B.n294 B.n293 585
R32 B.n292 B.n291 585
R33 B.n290 B.n289 585
R34 B.n288 B.n287 585
R35 B.n286 B.n285 585
R36 B.n284 B.n283 585
R37 B.n282 B.n281 585
R38 B.n280 B.n279 585
R39 B.n278 B.n277 585
R40 B.n276 B.n275 585
R41 B.n274 B.n273 585
R42 B.n272 B.n271 585
R43 B.n270 B.n269 585
R44 B.n268 B.n267 585
R45 B.n266 B.n265 585
R46 B.n264 B.n263 585
R47 B.n262 B.n261 585
R48 B.n260 B.n259 585
R49 B.n258 B.n257 585
R50 B.n256 B.n255 585
R51 B.n254 B.n253 585
R52 B.n252 B.n251 585
R53 B.n250 B.n249 585
R54 B.n248 B.n247 585
R55 B.n246 B.n245 585
R56 B.n244 B.n243 585
R57 B.n242 B.n241 585
R58 B.n240 B.n239 585
R59 B.n238 B.n237 585
R60 B.n236 B.n235 585
R61 B.n234 B.n233 585
R62 B.n232 B.n231 585
R63 B.n230 B.n229 585
R64 B.n228 B.n227 585
R65 B.n226 B.n225 585
R66 B.n224 B.n223 585
R67 B.n222 B.n221 585
R68 B.n220 B.n219 585
R69 B.n218 B.n217 585
R70 B.n216 B.n215 585
R71 B.n214 B.n213 585
R72 B.n212 B.n211 585
R73 B.n210 B.n209 585
R74 B.n208 B.n207 585
R75 B.n206 B.n205 585
R76 B.n204 B.n203 585
R77 B.n202 B.n201 585
R78 B.n200 B.n199 585
R79 B.n198 B.n197 585
R80 B.n196 B.n195 585
R81 B.n194 B.n193 585
R82 B.n192 B.n191 585
R83 B.n190 B.n189 585
R84 B.n188 B.n187 585
R85 B.n186 B.n185 585
R86 B.n184 B.n183 585
R87 B.n182 B.n181 585
R88 B.n180 B.n179 585
R89 B.n178 B.n177 585
R90 B.n176 B.n175 585
R91 B.n174 B.n173 585
R92 B.n172 B.n171 585
R93 B.n170 B.n169 585
R94 B.n168 B.n167 585
R95 B.n166 B.n165 585
R96 B.n164 B.n163 585
R97 B.n162 B.n161 585
R98 B.n160 B.n159 585
R99 B.n158 B.n157 585
R100 B.n156 B.n155 585
R101 B.n154 B.n153 585
R102 B.n152 B.n151 585
R103 B.n150 B.n149 585
R104 B.n148 B.n147 585
R105 B.n146 B.n145 585
R106 B.n144 B.n143 585
R107 B.n142 B.n141 585
R108 B.n140 B.n139 585
R109 B.n138 B.n137 585
R110 B.n136 B.n135 585
R111 B.n134 B.n133 585
R112 B.n132 B.n131 585
R113 B.n130 B.n129 585
R114 B.n128 B.n127 585
R115 B.n126 B.n125 585
R116 B.n124 B.n123 585
R117 B.n122 B.n121 585
R118 B.n120 B.n119 585
R119 B.n118 B.n117 585
R120 B.n116 B.n115 585
R121 B.n46 B.n45 585
R122 B.n812 B.n47 585
R123 B.n817 B.n47 585
R124 B.n811 B.n810 585
R125 B.n810 B.n43 585
R126 B.n809 B.n42 585
R127 B.n823 B.n42 585
R128 B.n808 B.n41 585
R129 B.n824 B.n41 585
R130 B.n807 B.n40 585
R131 B.n825 B.n40 585
R132 B.n806 B.n805 585
R133 B.n805 B.n39 585
R134 B.n804 B.n35 585
R135 B.n831 B.n35 585
R136 B.n803 B.n34 585
R137 B.n832 B.n34 585
R138 B.n802 B.n33 585
R139 B.n833 B.n33 585
R140 B.n801 B.n800 585
R141 B.n800 B.n29 585
R142 B.n799 B.n28 585
R143 B.n839 B.n28 585
R144 B.n798 B.n27 585
R145 B.n840 B.n27 585
R146 B.n797 B.n26 585
R147 B.n841 B.n26 585
R148 B.n796 B.n795 585
R149 B.n795 B.n22 585
R150 B.n794 B.n21 585
R151 B.n847 B.n21 585
R152 B.n793 B.n20 585
R153 B.n848 B.n20 585
R154 B.n792 B.n19 585
R155 B.n849 B.n19 585
R156 B.n791 B.n790 585
R157 B.n790 B.n15 585
R158 B.n789 B.n14 585
R159 B.n855 B.n14 585
R160 B.n788 B.n13 585
R161 B.n856 B.n13 585
R162 B.n787 B.n12 585
R163 B.n857 B.n12 585
R164 B.n786 B.n785 585
R165 B.n785 B.n8 585
R166 B.n784 B.n7 585
R167 B.n863 B.n7 585
R168 B.n783 B.n6 585
R169 B.n864 B.n6 585
R170 B.n782 B.n5 585
R171 B.n865 B.n5 585
R172 B.n781 B.n780 585
R173 B.n780 B.n4 585
R174 B.n779 B.n354 585
R175 B.n779 B.n778 585
R176 B.n769 B.n355 585
R177 B.n356 B.n355 585
R178 B.n771 B.n770 585
R179 B.n772 B.n771 585
R180 B.n768 B.n360 585
R181 B.n364 B.n360 585
R182 B.n767 B.n766 585
R183 B.n766 B.n765 585
R184 B.n362 B.n361 585
R185 B.n363 B.n362 585
R186 B.n758 B.n757 585
R187 B.n759 B.n758 585
R188 B.n756 B.n369 585
R189 B.n369 B.n368 585
R190 B.n755 B.n754 585
R191 B.n754 B.n753 585
R192 B.n371 B.n370 585
R193 B.n372 B.n371 585
R194 B.n746 B.n745 585
R195 B.n747 B.n746 585
R196 B.n744 B.n377 585
R197 B.n377 B.n376 585
R198 B.n743 B.n742 585
R199 B.n742 B.n741 585
R200 B.n379 B.n378 585
R201 B.n380 B.n379 585
R202 B.n734 B.n733 585
R203 B.n735 B.n734 585
R204 B.n732 B.n385 585
R205 B.n385 B.n384 585
R206 B.n731 B.n730 585
R207 B.n730 B.n729 585
R208 B.n387 B.n386 585
R209 B.n722 B.n387 585
R210 B.n721 B.n720 585
R211 B.n723 B.n721 585
R212 B.n719 B.n392 585
R213 B.n392 B.n391 585
R214 B.n718 B.n717 585
R215 B.n717 B.n716 585
R216 B.n394 B.n393 585
R217 B.n395 B.n394 585
R218 B.n709 B.n708 585
R219 B.n710 B.n709 585
R220 B.n398 B.n397 585
R221 B.n465 B.n463 585
R222 B.n466 B.n462 585
R223 B.n466 B.n399 585
R224 B.n469 B.n468 585
R225 B.n470 B.n461 585
R226 B.n472 B.n471 585
R227 B.n474 B.n460 585
R228 B.n477 B.n476 585
R229 B.n478 B.n459 585
R230 B.n480 B.n479 585
R231 B.n482 B.n458 585
R232 B.n485 B.n484 585
R233 B.n486 B.n457 585
R234 B.n488 B.n487 585
R235 B.n490 B.n456 585
R236 B.n493 B.n492 585
R237 B.n494 B.n455 585
R238 B.n496 B.n495 585
R239 B.n498 B.n454 585
R240 B.n501 B.n500 585
R241 B.n502 B.n453 585
R242 B.n504 B.n503 585
R243 B.n506 B.n452 585
R244 B.n509 B.n508 585
R245 B.n510 B.n451 585
R246 B.n512 B.n511 585
R247 B.n514 B.n450 585
R248 B.n517 B.n516 585
R249 B.n518 B.n449 585
R250 B.n520 B.n519 585
R251 B.n522 B.n448 585
R252 B.n525 B.n524 585
R253 B.n526 B.n447 585
R254 B.n528 B.n527 585
R255 B.n530 B.n446 585
R256 B.n533 B.n532 585
R257 B.n534 B.n445 585
R258 B.n536 B.n535 585
R259 B.n538 B.n444 585
R260 B.n541 B.n540 585
R261 B.n542 B.n443 585
R262 B.n544 B.n543 585
R263 B.n546 B.n442 585
R264 B.n549 B.n548 585
R265 B.n550 B.n441 585
R266 B.n552 B.n551 585
R267 B.n554 B.n440 585
R268 B.n557 B.n556 585
R269 B.n558 B.n439 585
R270 B.n560 B.n559 585
R271 B.n562 B.n438 585
R272 B.n565 B.n564 585
R273 B.n566 B.n437 585
R274 B.n568 B.n567 585
R275 B.n570 B.n436 585
R276 B.n573 B.n572 585
R277 B.n575 B.n433 585
R278 B.n577 B.n576 585
R279 B.n579 B.n432 585
R280 B.n582 B.n581 585
R281 B.n583 B.n431 585
R282 B.n585 B.n584 585
R283 B.n587 B.n430 585
R284 B.n590 B.n589 585
R285 B.n591 B.n429 585
R286 B.n596 B.n595 585
R287 B.n598 B.n428 585
R288 B.n601 B.n600 585
R289 B.n602 B.n427 585
R290 B.n604 B.n603 585
R291 B.n606 B.n426 585
R292 B.n609 B.n608 585
R293 B.n610 B.n425 585
R294 B.n612 B.n611 585
R295 B.n614 B.n424 585
R296 B.n617 B.n616 585
R297 B.n618 B.n423 585
R298 B.n620 B.n619 585
R299 B.n622 B.n422 585
R300 B.n625 B.n624 585
R301 B.n626 B.n421 585
R302 B.n628 B.n627 585
R303 B.n630 B.n420 585
R304 B.n633 B.n632 585
R305 B.n634 B.n419 585
R306 B.n636 B.n635 585
R307 B.n638 B.n418 585
R308 B.n641 B.n640 585
R309 B.n642 B.n417 585
R310 B.n644 B.n643 585
R311 B.n646 B.n416 585
R312 B.n649 B.n648 585
R313 B.n650 B.n415 585
R314 B.n652 B.n651 585
R315 B.n654 B.n414 585
R316 B.n657 B.n656 585
R317 B.n658 B.n413 585
R318 B.n660 B.n659 585
R319 B.n662 B.n412 585
R320 B.n665 B.n664 585
R321 B.n666 B.n411 585
R322 B.n668 B.n667 585
R323 B.n670 B.n410 585
R324 B.n673 B.n672 585
R325 B.n674 B.n409 585
R326 B.n676 B.n675 585
R327 B.n678 B.n408 585
R328 B.n681 B.n680 585
R329 B.n682 B.n407 585
R330 B.n684 B.n683 585
R331 B.n686 B.n406 585
R332 B.n689 B.n688 585
R333 B.n690 B.n405 585
R334 B.n692 B.n691 585
R335 B.n694 B.n404 585
R336 B.n697 B.n696 585
R337 B.n698 B.n403 585
R338 B.n700 B.n699 585
R339 B.n702 B.n402 585
R340 B.n703 B.n401 585
R341 B.n706 B.n705 585
R342 B.n707 B.n400 585
R343 B.n400 B.n399 585
R344 B.n712 B.n711 585
R345 B.n711 B.n710 585
R346 B.n713 B.n396 585
R347 B.n396 B.n395 585
R348 B.n715 B.n714 585
R349 B.n716 B.n715 585
R350 B.n390 B.n389 585
R351 B.n391 B.n390 585
R352 B.n725 B.n724 585
R353 B.n724 B.n723 585
R354 B.n726 B.n388 585
R355 B.n722 B.n388 585
R356 B.n728 B.n727 585
R357 B.n729 B.n728 585
R358 B.n383 B.n382 585
R359 B.n384 B.n383 585
R360 B.n737 B.n736 585
R361 B.n736 B.n735 585
R362 B.n738 B.n381 585
R363 B.n381 B.n380 585
R364 B.n740 B.n739 585
R365 B.n741 B.n740 585
R366 B.n375 B.n374 585
R367 B.n376 B.n375 585
R368 B.n749 B.n748 585
R369 B.n748 B.n747 585
R370 B.n750 B.n373 585
R371 B.n373 B.n372 585
R372 B.n752 B.n751 585
R373 B.n753 B.n752 585
R374 B.n367 B.n366 585
R375 B.n368 B.n367 585
R376 B.n761 B.n760 585
R377 B.n760 B.n759 585
R378 B.n762 B.n365 585
R379 B.n365 B.n363 585
R380 B.n764 B.n763 585
R381 B.n765 B.n764 585
R382 B.n359 B.n358 585
R383 B.n364 B.n359 585
R384 B.n774 B.n773 585
R385 B.n773 B.n772 585
R386 B.n775 B.n357 585
R387 B.n357 B.n356 585
R388 B.n777 B.n776 585
R389 B.n778 B.n777 585
R390 B.n2 B.n0 585
R391 B.n4 B.n2 585
R392 B.n3 B.n1 585
R393 B.n864 B.n3 585
R394 B.n862 B.n861 585
R395 B.n863 B.n862 585
R396 B.n860 B.n9 585
R397 B.n9 B.n8 585
R398 B.n859 B.n858 585
R399 B.n858 B.n857 585
R400 B.n11 B.n10 585
R401 B.n856 B.n11 585
R402 B.n854 B.n853 585
R403 B.n855 B.n854 585
R404 B.n852 B.n16 585
R405 B.n16 B.n15 585
R406 B.n851 B.n850 585
R407 B.n850 B.n849 585
R408 B.n18 B.n17 585
R409 B.n848 B.n18 585
R410 B.n846 B.n845 585
R411 B.n847 B.n846 585
R412 B.n844 B.n23 585
R413 B.n23 B.n22 585
R414 B.n843 B.n842 585
R415 B.n842 B.n841 585
R416 B.n25 B.n24 585
R417 B.n840 B.n25 585
R418 B.n838 B.n837 585
R419 B.n839 B.n838 585
R420 B.n836 B.n30 585
R421 B.n30 B.n29 585
R422 B.n835 B.n834 585
R423 B.n834 B.n833 585
R424 B.n32 B.n31 585
R425 B.n832 B.n32 585
R426 B.n830 B.n829 585
R427 B.n831 B.n830 585
R428 B.n828 B.n36 585
R429 B.n39 B.n36 585
R430 B.n827 B.n826 585
R431 B.n826 B.n825 585
R432 B.n38 B.n37 585
R433 B.n824 B.n38 585
R434 B.n822 B.n821 585
R435 B.n823 B.n822 585
R436 B.n820 B.n44 585
R437 B.n44 B.n43 585
R438 B.n819 B.n818 585
R439 B.n818 B.n817 585
R440 B.n867 B.n866 585
R441 B.n866 B.n865 585
R442 B.n711 B.n398 516.524
R443 B.n818 B.n46 516.524
R444 B.n709 B.n400 516.524
R445 B.n814 B.n47 516.524
R446 B.n592 B.t4 479.399
R447 B.n434 B.t15 479.399
R448 B.n112 B.t8 479.399
R449 B.n109 B.t12 479.399
R450 B.n592 B.t7 402.783
R451 B.n109 B.t13 402.783
R452 B.n434 B.t17 402.783
R453 B.n112 B.t10 402.783
R454 B.n593 B.t6 367.486
R455 B.n110 B.t14 367.486
R456 B.n435 B.t16 367.486
R457 B.n113 B.t11 367.486
R458 B.n816 B.n815 256.663
R459 B.n816 B.n107 256.663
R460 B.n816 B.n106 256.663
R461 B.n816 B.n105 256.663
R462 B.n816 B.n104 256.663
R463 B.n816 B.n103 256.663
R464 B.n816 B.n102 256.663
R465 B.n816 B.n101 256.663
R466 B.n816 B.n100 256.663
R467 B.n816 B.n99 256.663
R468 B.n816 B.n98 256.663
R469 B.n816 B.n97 256.663
R470 B.n816 B.n96 256.663
R471 B.n816 B.n95 256.663
R472 B.n816 B.n94 256.663
R473 B.n816 B.n93 256.663
R474 B.n816 B.n92 256.663
R475 B.n816 B.n91 256.663
R476 B.n816 B.n90 256.663
R477 B.n816 B.n89 256.663
R478 B.n816 B.n88 256.663
R479 B.n816 B.n87 256.663
R480 B.n816 B.n86 256.663
R481 B.n816 B.n85 256.663
R482 B.n816 B.n84 256.663
R483 B.n816 B.n83 256.663
R484 B.n816 B.n82 256.663
R485 B.n816 B.n81 256.663
R486 B.n816 B.n80 256.663
R487 B.n816 B.n79 256.663
R488 B.n816 B.n78 256.663
R489 B.n816 B.n77 256.663
R490 B.n816 B.n76 256.663
R491 B.n816 B.n75 256.663
R492 B.n816 B.n74 256.663
R493 B.n816 B.n73 256.663
R494 B.n816 B.n72 256.663
R495 B.n816 B.n71 256.663
R496 B.n816 B.n70 256.663
R497 B.n816 B.n69 256.663
R498 B.n816 B.n68 256.663
R499 B.n816 B.n67 256.663
R500 B.n816 B.n66 256.663
R501 B.n816 B.n65 256.663
R502 B.n816 B.n64 256.663
R503 B.n816 B.n63 256.663
R504 B.n816 B.n62 256.663
R505 B.n816 B.n61 256.663
R506 B.n816 B.n60 256.663
R507 B.n816 B.n59 256.663
R508 B.n816 B.n58 256.663
R509 B.n816 B.n57 256.663
R510 B.n816 B.n56 256.663
R511 B.n816 B.n55 256.663
R512 B.n816 B.n54 256.663
R513 B.n816 B.n53 256.663
R514 B.n816 B.n52 256.663
R515 B.n816 B.n51 256.663
R516 B.n816 B.n50 256.663
R517 B.n816 B.n49 256.663
R518 B.n816 B.n48 256.663
R519 B.n464 B.n399 256.663
R520 B.n467 B.n399 256.663
R521 B.n473 B.n399 256.663
R522 B.n475 B.n399 256.663
R523 B.n481 B.n399 256.663
R524 B.n483 B.n399 256.663
R525 B.n489 B.n399 256.663
R526 B.n491 B.n399 256.663
R527 B.n497 B.n399 256.663
R528 B.n499 B.n399 256.663
R529 B.n505 B.n399 256.663
R530 B.n507 B.n399 256.663
R531 B.n513 B.n399 256.663
R532 B.n515 B.n399 256.663
R533 B.n521 B.n399 256.663
R534 B.n523 B.n399 256.663
R535 B.n529 B.n399 256.663
R536 B.n531 B.n399 256.663
R537 B.n537 B.n399 256.663
R538 B.n539 B.n399 256.663
R539 B.n545 B.n399 256.663
R540 B.n547 B.n399 256.663
R541 B.n553 B.n399 256.663
R542 B.n555 B.n399 256.663
R543 B.n561 B.n399 256.663
R544 B.n563 B.n399 256.663
R545 B.n569 B.n399 256.663
R546 B.n571 B.n399 256.663
R547 B.n578 B.n399 256.663
R548 B.n580 B.n399 256.663
R549 B.n586 B.n399 256.663
R550 B.n588 B.n399 256.663
R551 B.n597 B.n399 256.663
R552 B.n599 B.n399 256.663
R553 B.n605 B.n399 256.663
R554 B.n607 B.n399 256.663
R555 B.n613 B.n399 256.663
R556 B.n615 B.n399 256.663
R557 B.n621 B.n399 256.663
R558 B.n623 B.n399 256.663
R559 B.n629 B.n399 256.663
R560 B.n631 B.n399 256.663
R561 B.n637 B.n399 256.663
R562 B.n639 B.n399 256.663
R563 B.n645 B.n399 256.663
R564 B.n647 B.n399 256.663
R565 B.n653 B.n399 256.663
R566 B.n655 B.n399 256.663
R567 B.n661 B.n399 256.663
R568 B.n663 B.n399 256.663
R569 B.n669 B.n399 256.663
R570 B.n671 B.n399 256.663
R571 B.n677 B.n399 256.663
R572 B.n679 B.n399 256.663
R573 B.n685 B.n399 256.663
R574 B.n687 B.n399 256.663
R575 B.n693 B.n399 256.663
R576 B.n695 B.n399 256.663
R577 B.n701 B.n399 256.663
R578 B.n704 B.n399 256.663
R579 B.n711 B.n396 163.367
R580 B.n715 B.n396 163.367
R581 B.n715 B.n390 163.367
R582 B.n724 B.n390 163.367
R583 B.n724 B.n388 163.367
R584 B.n728 B.n388 163.367
R585 B.n728 B.n383 163.367
R586 B.n736 B.n383 163.367
R587 B.n736 B.n381 163.367
R588 B.n740 B.n381 163.367
R589 B.n740 B.n375 163.367
R590 B.n748 B.n375 163.367
R591 B.n748 B.n373 163.367
R592 B.n752 B.n373 163.367
R593 B.n752 B.n367 163.367
R594 B.n760 B.n367 163.367
R595 B.n760 B.n365 163.367
R596 B.n764 B.n365 163.367
R597 B.n764 B.n359 163.367
R598 B.n773 B.n359 163.367
R599 B.n773 B.n357 163.367
R600 B.n777 B.n357 163.367
R601 B.n777 B.n2 163.367
R602 B.n866 B.n2 163.367
R603 B.n866 B.n3 163.367
R604 B.n862 B.n3 163.367
R605 B.n862 B.n9 163.367
R606 B.n858 B.n9 163.367
R607 B.n858 B.n11 163.367
R608 B.n854 B.n11 163.367
R609 B.n854 B.n16 163.367
R610 B.n850 B.n16 163.367
R611 B.n850 B.n18 163.367
R612 B.n846 B.n18 163.367
R613 B.n846 B.n23 163.367
R614 B.n842 B.n23 163.367
R615 B.n842 B.n25 163.367
R616 B.n838 B.n25 163.367
R617 B.n838 B.n30 163.367
R618 B.n834 B.n30 163.367
R619 B.n834 B.n32 163.367
R620 B.n830 B.n32 163.367
R621 B.n830 B.n36 163.367
R622 B.n826 B.n36 163.367
R623 B.n826 B.n38 163.367
R624 B.n822 B.n38 163.367
R625 B.n822 B.n44 163.367
R626 B.n818 B.n44 163.367
R627 B.n466 B.n465 163.367
R628 B.n468 B.n466 163.367
R629 B.n472 B.n461 163.367
R630 B.n476 B.n474 163.367
R631 B.n480 B.n459 163.367
R632 B.n484 B.n482 163.367
R633 B.n488 B.n457 163.367
R634 B.n492 B.n490 163.367
R635 B.n496 B.n455 163.367
R636 B.n500 B.n498 163.367
R637 B.n504 B.n453 163.367
R638 B.n508 B.n506 163.367
R639 B.n512 B.n451 163.367
R640 B.n516 B.n514 163.367
R641 B.n520 B.n449 163.367
R642 B.n524 B.n522 163.367
R643 B.n528 B.n447 163.367
R644 B.n532 B.n530 163.367
R645 B.n536 B.n445 163.367
R646 B.n540 B.n538 163.367
R647 B.n544 B.n443 163.367
R648 B.n548 B.n546 163.367
R649 B.n552 B.n441 163.367
R650 B.n556 B.n554 163.367
R651 B.n560 B.n439 163.367
R652 B.n564 B.n562 163.367
R653 B.n568 B.n437 163.367
R654 B.n572 B.n570 163.367
R655 B.n577 B.n433 163.367
R656 B.n581 B.n579 163.367
R657 B.n585 B.n431 163.367
R658 B.n589 B.n587 163.367
R659 B.n596 B.n429 163.367
R660 B.n600 B.n598 163.367
R661 B.n604 B.n427 163.367
R662 B.n608 B.n606 163.367
R663 B.n612 B.n425 163.367
R664 B.n616 B.n614 163.367
R665 B.n620 B.n423 163.367
R666 B.n624 B.n622 163.367
R667 B.n628 B.n421 163.367
R668 B.n632 B.n630 163.367
R669 B.n636 B.n419 163.367
R670 B.n640 B.n638 163.367
R671 B.n644 B.n417 163.367
R672 B.n648 B.n646 163.367
R673 B.n652 B.n415 163.367
R674 B.n656 B.n654 163.367
R675 B.n660 B.n413 163.367
R676 B.n664 B.n662 163.367
R677 B.n668 B.n411 163.367
R678 B.n672 B.n670 163.367
R679 B.n676 B.n409 163.367
R680 B.n680 B.n678 163.367
R681 B.n684 B.n407 163.367
R682 B.n688 B.n686 163.367
R683 B.n692 B.n405 163.367
R684 B.n696 B.n694 163.367
R685 B.n700 B.n403 163.367
R686 B.n703 B.n702 163.367
R687 B.n705 B.n400 163.367
R688 B.n709 B.n394 163.367
R689 B.n717 B.n394 163.367
R690 B.n717 B.n392 163.367
R691 B.n721 B.n392 163.367
R692 B.n721 B.n387 163.367
R693 B.n730 B.n387 163.367
R694 B.n730 B.n385 163.367
R695 B.n734 B.n385 163.367
R696 B.n734 B.n379 163.367
R697 B.n742 B.n379 163.367
R698 B.n742 B.n377 163.367
R699 B.n746 B.n377 163.367
R700 B.n746 B.n371 163.367
R701 B.n754 B.n371 163.367
R702 B.n754 B.n369 163.367
R703 B.n758 B.n369 163.367
R704 B.n758 B.n362 163.367
R705 B.n766 B.n362 163.367
R706 B.n766 B.n360 163.367
R707 B.n771 B.n360 163.367
R708 B.n771 B.n355 163.367
R709 B.n779 B.n355 163.367
R710 B.n780 B.n779 163.367
R711 B.n780 B.n5 163.367
R712 B.n6 B.n5 163.367
R713 B.n7 B.n6 163.367
R714 B.n785 B.n7 163.367
R715 B.n785 B.n12 163.367
R716 B.n13 B.n12 163.367
R717 B.n14 B.n13 163.367
R718 B.n790 B.n14 163.367
R719 B.n790 B.n19 163.367
R720 B.n20 B.n19 163.367
R721 B.n21 B.n20 163.367
R722 B.n795 B.n21 163.367
R723 B.n795 B.n26 163.367
R724 B.n27 B.n26 163.367
R725 B.n28 B.n27 163.367
R726 B.n800 B.n28 163.367
R727 B.n800 B.n33 163.367
R728 B.n34 B.n33 163.367
R729 B.n35 B.n34 163.367
R730 B.n805 B.n35 163.367
R731 B.n805 B.n40 163.367
R732 B.n41 B.n40 163.367
R733 B.n42 B.n41 163.367
R734 B.n810 B.n42 163.367
R735 B.n810 B.n47 163.367
R736 B.n117 B.n116 163.367
R737 B.n121 B.n120 163.367
R738 B.n125 B.n124 163.367
R739 B.n129 B.n128 163.367
R740 B.n133 B.n132 163.367
R741 B.n137 B.n136 163.367
R742 B.n141 B.n140 163.367
R743 B.n145 B.n144 163.367
R744 B.n149 B.n148 163.367
R745 B.n153 B.n152 163.367
R746 B.n157 B.n156 163.367
R747 B.n161 B.n160 163.367
R748 B.n165 B.n164 163.367
R749 B.n169 B.n168 163.367
R750 B.n173 B.n172 163.367
R751 B.n177 B.n176 163.367
R752 B.n181 B.n180 163.367
R753 B.n185 B.n184 163.367
R754 B.n189 B.n188 163.367
R755 B.n193 B.n192 163.367
R756 B.n197 B.n196 163.367
R757 B.n201 B.n200 163.367
R758 B.n205 B.n204 163.367
R759 B.n209 B.n208 163.367
R760 B.n213 B.n212 163.367
R761 B.n217 B.n216 163.367
R762 B.n221 B.n220 163.367
R763 B.n225 B.n224 163.367
R764 B.n229 B.n228 163.367
R765 B.n233 B.n232 163.367
R766 B.n237 B.n236 163.367
R767 B.n241 B.n240 163.367
R768 B.n245 B.n244 163.367
R769 B.n249 B.n248 163.367
R770 B.n253 B.n252 163.367
R771 B.n257 B.n256 163.367
R772 B.n261 B.n260 163.367
R773 B.n265 B.n264 163.367
R774 B.n269 B.n268 163.367
R775 B.n273 B.n272 163.367
R776 B.n277 B.n276 163.367
R777 B.n281 B.n280 163.367
R778 B.n285 B.n284 163.367
R779 B.n289 B.n288 163.367
R780 B.n293 B.n292 163.367
R781 B.n297 B.n296 163.367
R782 B.n301 B.n300 163.367
R783 B.n305 B.n304 163.367
R784 B.n309 B.n308 163.367
R785 B.n313 B.n312 163.367
R786 B.n317 B.n316 163.367
R787 B.n321 B.n320 163.367
R788 B.n325 B.n324 163.367
R789 B.n329 B.n328 163.367
R790 B.n333 B.n332 163.367
R791 B.n337 B.n336 163.367
R792 B.n341 B.n340 163.367
R793 B.n345 B.n344 163.367
R794 B.n349 B.n348 163.367
R795 B.n351 B.n108 163.367
R796 B.n464 B.n398 71.676
R797 B.n468 B.n467 71.676
R798 B.n473 B.n472 71.676
R799 B.n476 B.n475 71.676
R800 B.n481 B.n480 71.676
R801 B.n484 B.n483 71.676
R802 B.n489 B.n488 71.676
R803 B.n492 B.n491 71.676
R804 B.n497 B.n496 71.676
R805 B.n500 B.n499 71.676
R806 B.n505 B.n504 71.676
R807 B.n508 B.n507 71.676
R808 B.n513 B.n512 71.676
R809 B.n516 B.n515 71.676
R810 B.n521 B.n520 71.676
R811 B.n524 B.n523 71.676
R812 B.n529 B.n528 71.676
R813 B.n532 B.n531 71.676
R814 B.n537 B.n536 71.676
R815 B.n540 B.n539 71.676
R816 B.n545 B.n544 71.676
R817 B.n548 B.n547 71.676
R818 B.n553 B.n552 71.676
R819 B.n556 B.n555 71.676
R820 B.n561 B.n560 71.676
R821 B.n564 B.n563 71.676
R822 B.n569 B.n568 71.676
R823 B.n572 B.n571 71.676
R824 B.n578 B.n577 71.676
R825 B.n581 B.n580 71.676
R826 B.n586 B.n585 71.676
R827 B.n589 B.n588 71.676
R828 B.n597 B.n596 71.676
R829 B.n600 B.n599 71.676
R830 B.n605 B.n604 71.676
R831 B.n608 B.n607 71.676
R832 B.n613 B.n612 71.676
R833 B.n616 B.n615 71.676
R834 B.n621 B.n620 71.676
R835 B.n624 B.n623 71.676
R836 B.n629 B.n628 71.676
R837 B.n632 B.n631 71.676
R838 B.n637 B.n636 71.676
R839 B.n640 B.n639 71.676
R840 B.n645 B.n644 71.676
R841 B.n648 B.n647 71.676
R842 B.n653 B.n652 71.676
R843 B.n656 B.n655 71.676
R844 B.n661 B.n660 71.676
R845 B.n664 B.n663 71.676
R846 B.n669 B.n668 71.676
R847 B.n672 B.n671 71.676
R848 B.n677 B.n676 71.676
R849 B.n680 B.n679 71.676
R850 B.n685 B.n684 71.676
R851 B.n688 B.n687 71.676
R852 B.n693 B.n692 71.676
R853 B.n696 B.n695 71.676
R854 B.n701 B.n700 71.676
R855 B.n704 B.n703 71.676
R856 B.n48 B.n46 71.676
R857 B.n117 B.n49 71.676
R858 B.n121 B.n50 71.676
R859 B.n125 B.n51 71.676
R860 B.n129 B.n52 71.676
R861 B.n133 B.n53 71.676
R862 B.n137 B.n54 71.676
R863 B.n141 B.n55 71.676
R864 B.n145 B.n56 71.676
R865 B.n149 B.n57 71.676
R866 B.n153 B.n58 71.676
R867 B.n157 B.n59 71.676
R868 B.n161 B.n60 71.676
R869 B.n165 B.n61 71.676
R870 B.n169 B.n62 71.676
R871 B.n173 B.n63 71.676
R872 B.n177 B.n64 71.676
R873 B.n181 B.n65 71.676
R874 B.n185 B.n66 71.676
R875 B.n189 B.n67 71.676
R876 B.n193 B.n68 71.676
R877 B.n197 B.n69 71.676
R878 B.n201 B.n70 71.676
R879 B.n205 B.n71 71.676
R880 B.n209 B.n72 71.676
R881 B.n213 B.n73 71.676
R882 B.n217 B.n74 71.676
R883 B.n221 B.n75 71.676
R884 B.n225 B.n76 71.676
R885 B.n229 B.n77 71.676
R886 B.n233 B.n78 71.676
R887 B.n237 B.n79 71.676
R888 B.n241 B.n80 71.676
R889 B.n245 B.n81 71.676
R890 B.n249 B.n82 71.676
R891 B.n253 B.n83 71.676
R892 B.n257 B.n84 71.676
R893 B.n261 B.n85 71.676
R894 B.n265 B.n86 71.676
R895 B.n269 B.n87 71.676
R896 B.n273 B.n88 71.676
R897 B.n277 B.n89 71.676
R898 B.n281 B.n90 71.676
R899 B.n285 B.n91 71.676
R900 B.n289 B.n92 71.676
R901 B.n293 B.n93 71.676
R902 B.n297 B.n94 71.676
R903 B.n301 B.n95 71.676
R904 B.n305 B.n96 71.676
R905 B.n309 B.n97 71.676
R906 B.n313 B.n98 71.676
R907 B.n317 B.n99 71.676
R908 B.n321 B.n100 71.676
R909 B.n325 B.n101 71.676
R910 B.n329 B.n102 71.676
R911 B.n333 B.n103 71.676
R912 B.n337 B.n104 71.676
R913 B.n341 B.n105 71.676
R914 B.n345 B.n106 71.676
R915 B.n349 B.n107 71.676
R916 B.n815 B.n108 71.676
R917 B.n815 B.n814 71.676
R918 B.n351 B.n107 71.676
R919 B.n348 B.n106 71.676
R920 B.n344 B.n105 71.676
R921 B.n340 B.n104 71.676
R922 B.n336 B.n103 71.676
R923 B.n332 B.n102 71.676
R924 B.n328 B.n101 71.676
R925 B.n324 B.n100 71.676
R926 B.n320 B.n99 71.676
R927 B.n316 B.n98 71.676
R928 B.n312 B.n97 71.676
R929 B.n308 B.n96 71.676
R930 B.n304 B.n95 71.676
R931 B.n300 B.n94 71.676
R932 B.n296 B.n93 71.676
R933 B.n292 B.n92 71.676
R934 B.n288 B.n91 71.676
R935 B.n284 B.n90 71.676
R936 B.n280 B.n89 71.676
R937 B.n276 B.n88 71.676
R938 B.n272 B.n87 71.676
R939 B.n268 B.n86 71.676
R940 B.n264 B.n85 71.676
R941 B.n260 B.n84 71.676
R942 B.n256 B.n83 71.676
R943 B.n252 B.n82 71.676
R944 B.n248 B.n81 71.676
R945 B.n244 B.n80 71.676
R946 B.n240 B.n79 71.676
R947 B.n236 B.n78 71.676
R948 B.n232 B.n77 71.676
R949 B.n228 B.n76 71.676
R950 B.n224 B.n75 71.676
R951 B.n220 B.n74 71.676
R952 B.n216 B.n73 71.676
R953 B.n212 B.n72 71.676
R954 B.n208 B.n71 71.676
R955 B.n204 B.n70 71.676
R956 B.n200 B.n69 71.676
R957 B.n196 B.n68 71.676
R958 B.n192 B.n67 71.676
R959 B.n188 B.n66 71.676
R960 B.n184 B.n65 71.676
R961 B.n180 B.n64 71.676
R962 B.n176 B.n63 71.676
R963 B.n172 B.n62 71.676
R964 B.n168 B.n61 71.676
R965 B.n164 B.n60 71.676
R966 B.n160 B.n59 71.676
R967 B.n156 B.n58 71.676
R968 B.n152 B.n57 71.676
R969 B.n148 B.n56 71.676
R970 B.n144 B.n55 71.676
R971 B.n140 B.n54 71.676
R972 B.n136 B.n53 71.676
R973 B.n132 B.n52 71.676
R974 B.n128 B.n51 71.676
R975 B.n124 B.n50 71.676
R976 B.n120 B.n49 71.676
R977 B.n116 B.n48 71.676
R978 B.n465 B.n464 71.676
R979 B.n467 B.n461 71.676
R980 B.n474 B.n473 71.676
R981 B.n475 B.n459 71.676
R982 B.n482 B.n481 71.676
R983 B.n483 B.n457 71.676
R984 B.n490 B.n489 71.676
R985 B.n491 B.n455 71.676
R986 B.n498 B.n497 71.676
R987 B.n499 B.n453 71.676
R988 B.n506 B.n505 71.676
R989 B.n507 B.n451 71.676
R990 B.n514 B.n513 71.676
R991 B.n515 B.n449 71.676
R992 B.n522 B.n521 71.676
R993 B.n523 B.n447 71.676
R994 B.n530 B.n529 71.676
R995 B.n531 B.n445 71.676
R996 B.n538 B.n537 71.676
R997 B.n539 B.n443 71.676
R998 B.n546 B.n545 71.676
R999 B.n547 B.n441 71.676
R1000 B.n554 B.n553 71.676
R1001 B.n555 B.n439 71.676
R1002 B.n562 B.n561 71.676
R1003 B.n563 B.n437 71.676
R1004 B.n570 B.n569 71.676
R1005 B.n571 B.n433 71.676
R1006 B.n579 B.n578 71.676
R1007 B.n580 B.n431 71.676
R1008 B.n587 B.n586 71.676
R1009 B.n588 B.n429 71.676
R1010 B.n598 B.n597 71.676
R1011 B.n599 B.n427 71.676
R1012 B.n606 B.n605 71.676
R1013 B.n607 B.n425 71.676
R1014 B.n614 B.n613 71.676
R1015 B.n615 B.n423 71.676
R1016 B.n622 B.n621 71.676
R1017 B.n623 B.n421 71.676
R1018 B.n630 B.n629 71.676
R1019 B.n631 B.n419 71.676
R1020 B.n638 B.n637 71.676
R1021 B.n639 B.n417 71.676
R1022 B.n646 B.n645 71.676
R1023 B.n647 B.n415 71.676
R1024 B.n654 B.n653 71.676
R1025 B.n655 B.n413 71.676
R1026 B.n662 B.n661 71.676
R1027 B.n663 B.n411 71.676
R1028 B.n670 B.n669 71.676
R1029 B.n671 B.n409 71.676
R1030 B.n678 B.n677 71.676
R1031 B.n679 B.n407 71.676
R1032 B.n686 B.n685 71.676
R1033 B.n687 B.n405 71.676
R1034 B.n694 B.n693 71.676
R1035 B.n695 B.n403 71.676
R1036 B.n702 B.n701 71.676
R1037 B.n705 B.n704 71.676
R1038 B.n710 B.n399 66.8472
R1039 B.n817 B.n816 66.8472
R1040 B.n594 B.n593 59.5399
R1041 B.n574 B.n435 59.5399
R1042 B.n114 B.n113 59.5399
R1043 B.n111 B.n110 59.5399
R1044 B.n593 B.n592 35.2975
R1045 B.n435 B.n434 35.2975
R1046 B.n113 B.n112 35.2975
R1047 B.n110 B.n109 35.2975
R1048 B.n710 B.n395 33.6714
R1049 B.n716 B.n395 33.6714
R1050 B.n716 B.n391 33.6714
R1051 B.n723 B.n391 33.6714
R1052 B.n723 B.n722 33.6714
R1053 B.n729 B.n384 33.6714
R1054 B.n735 B.n384 33.6714
R1055 B.n735 B.n380 33.6714
R1056 B.n741 B.n380 33.6714
R1057 B.n741 B.n376 33.6714
R1058 B.n747 B.n376 33.6714
R1059 B.n747 B.n372 33.6714
R1060 B.n753 B.n372 33.6714
R1061 B.n759 B.n368 33.6714
R1062 B.n759 B.n363 33.6714
R1063 B.n765 B.n363 33.6714
R1064 B.n765 B.n364 33.6714
R1065 B.n772 B.n356 33.6714
R1066 B.n778 B.n356 33.6714
R1067 B.n778 B.n4 33.6714
R1068 B.n865 B.n4 33.6714
R1069 B.n865 B.n864 33.6714
R1070 B.n864 B.n863 33.6714
R1071 B.n863 B.n8 33.6714
R1072 B.n857 B.n8 33.6714
R1073 B.n856 B.n855 33.6714
R1074 B.n855 B.n15 33.6714
R1075 B.n849 B.n15 33.6714
R1076 B.n849 B.n848 33.6714
R1077 B.n847 B.n22 33.6714
R1078 B.n841 B.n22 33.6714
R1079 B.n841 B.n840 33.6714
R1080 B.n840 B.n839 33.6714
R1081 B.n839 B.n29 33.6714
R1082 B.n833 B.n29 33.6714
R1083 B.n833 B.n832 33.6714
R1084 B.n832 B.n831 33.6714
R1085 B.n825 B.n39 33.6714
R1086 B.n825 B.n824 33.6714
R1087 B.n824 B.n823 33.6714
R1088 B.n823 B.n43 33.6714
R1089 B.n817 B.n43 33.6714
R1090 B.n819 B.n45 33.5615
R1091 B.n813 B.n812 33.5615
R1092 B.n708 B.n707 33.5615
R1093 B.n712 B.n397 33.5615
R1094 B.n722 B.t5 27.2344
R1095 B.n39 B.t9 27.2344
R1096 B.n364 B.t2 24.2634
R1097 B.t1 B.n856 24.2634
R1098 B.t0 B.n368 21.2924
R1099 B.n848 B.t3 21.2924
R1100 B B.n867 18.0485
R1101 B.n753 B.t0 12.3795
R1102 B.t3 B.n847 12.3795
R1103 B.n115 B.n45 10.6151
R1104 B.n118 B.n115 10.6151
R1105 B.n119 B.n118 10.6151
R1106 B.n122 B.n119 10.6151
R1107 B.n123 B.n122 10.6151
R1108 B.n126 B.n123 10.6151
R1109 B.n127 B.n126 10.6151
R1110 B.n130 B.n127 10.6151
R1111 B.n131 B.n130 10.6151
R1112 B.n134 B.n131 10.6151
R1113 B.n135 B.n134 10.6151
R1114 B.n138 B.n135 10.6151
R1115 B.n139 B.n138 10.6151
R1116 B.n142 B.n139 10.6151
R1117 B.n143 B.n142 10.6151
R1118 B.n146 B.n143 10.6151
R1119 B.n147 B.n146 10.6151
R1120 B.n150 B.n147 10.6151
R1121 B.n151 B.n150 10.6151
R1122 B.n154 B.n151 10.6151
R1123 B.n155 B.n154 10.6151
R1124 B.n158 B.n155 10.6151
R1125 B.n159 B.n158 10.6151
R1126 B.n162 B.n159 10.6151
R1127 B.n163 B.n162 10.6151
R1128 B.n166 B.n163 10.6151
R1129 B.n167 B.n166 10.6151
R1130 B.n170 B.n167 10.6151
R1131 B.n171 B.n170 10.6151
R1132 B.n174 B.n171 10.6151
R1133 B.n175 B.n174 10.6151
R1134 B.n178 B.n175 10.6151
R1135 B.n179 B.n178 10.6151
R1136 B.n182 B.n179 10.6151
R1137 B.n183 B.n182 10.6151
R1138 B.n186 B.n183 10.6151
R1139 B.n187 B.n186 10.6151
R1140 B.n190 B.n187 10.6151
R1141 B.n191 B.n190 10.6151
R1142 B.n194 B.n191 10.6151
R1143 B.n195 B.n194 10.6151
R1144 B.n198 B.n195 10.6151
R1145 B.n199 B.n198 10.6151
R1146 B.n202 B.n199 10.6151
R1147 B.n203 B.n202 10.6151
R1148 B.n206 B.n203 10.6151
R1149 B.n207 B.n206 10.6151
R1150 B.n210 B.n207 10.6151
R1151 B.n211 B.n210 10.6151
R1152 B.n214 B.n211 10.6151
R1153 B.n215 B.n214 10.6151
R1154 B.n218 B.n215 10.6151
R1155 B.n219 B.n218 10.6151
R1156 B.n222 B.n219 10.6151
R1157 B.n223 B.n222 10.6151
R1158 B.n227 B.n226 10.6151
R1159 B.n230 B.n227 10.6151
R1160 B.n231 B.n230 10.6151
R1161 B.n234 B.n231 10.6151
R1162 B.n235 B.n234 10.6151
R1163 B.n238 B.n235 10.6151
R1164 B.n239 B.n238 10.6151
R1165 B.n242 B.n239 10.6151
R1166 B.n243 B.n242 10.6151
R1167 B.n247 B.n246 10.6151
R1168 B.n250 B.n247 10.6151
R1169 B.n251 B.n250 10.6151
R1170 B.n254 B.n251 10.6151
R1171 B.n255 B.n254 10.6151
R1172 B.n258 B.n255 10.6151
R1173 B.n259 B.n258 10.6151
R1174 B.n262 B.n259 10.6151
R1175 B.n263 B.n262 10.6151
R1176 B.n266 B.n263 10.6151
R1177 B.n267 B.n266 10.6151
R1178 B.n270 B.n267 10.6151
R1179 B.n271 B.n270 10.6151
R1180 B.n274 B.n271 10.6151
R1181 B.n275 B.n274 10.6151
R1182 B.n278 B.n275 10.6151
R1183 B.n279 B.n278 10.6151
R1184 B.n282 B.n279 10.6151
R1185 B.n283 B.n282 10.6151
R1186 B.n286 B.n283 10.6151
R1187 B.n287 B.n286 10.6151
R1188 B.n290 B.n287 10.6151
R1189 B.n291 B.n290 10.6151
R1190 B.n294 B.n291 10.6151
R1191 B.n295 B.n294 10.6151
R1192 B.n298 B.n295 10.6151
R1193 B.n299 B.n298 10.6151
R1194 B.n302 B.n299 10.6151
R1195 B.n303 B.n302 10.6151
R1196 B.n306 B.n303 10.6151
R1197 B.n307 B.n306 10.6151
R1198 B.n310 B.n307 10.6151
R1199 B.n311 B.n310 10.6151
R1200 B.n314 B.n311 10.6151
R1201 B.n315 B.n314 10.6151
R1202 B.n318 B.n315 10.6151
R1203 B.n319 B.n318 10.6151
R1204 B.n322 B.n319 10.6151
R1205 B.n323 B.n322 10.6151
R1206 B.n326 B.n323 10.6151
R1207 B.n327 B.n326 10.6151
R1208 B.n330 B.n327 10.6151
R1209 B.n331 B.n330 10.6151
R1210 B.n334 B.n331 10.6151
R1211 B.n335 B.n334 10.6151
R1212 B.n338 B.n335 10.6151
R1213 B.n339 B.n338 10.6151
R1214 B.n342 B.n339 10.6151
R1215 B.n343 B.n342 10.6151
R1216 B.n346 B.n343 10.6151
R1217 B.n347 B.n346 10.6151
R1218 B.n350 B.n347 10.6151
R1219 B.n352 B.n350 10.6151
R1220 B.n353 B.n352 10.6151
R1221 B.n813 B.n353 10.6151
R1222 B.n708 B.n393 10.6151
R1223 B.n718 B.n393 10.6151
R1224 B.n719 B.n718 10.6151
R1225 B.n720 B.n719 10.6151
R1226 B.n720 B.n386 10.6151
R1227 B.n731 B.n386 10.6151
R1228 B.n732 B.n731 10.6151
R1229 B.n733 B.n732 10.6151
R1230 B.n733 B.n378 10.6151
R1231 B.n743 B.n378 10.6151
R1232 B.n744 B.n743 10.6151
R1233 B.n745 B.n744 10.6151
R1234 B.n745 B.n370 10.6151
R1235 B.n755 B.n370 10.6151
R1236 B.n756 B.n755 10.6151
R1237 B.n757 B.n756 10.6151
R1238 B.n757 B.n361 10.6151
R1239 B.n767 B.n361 10.6151
R1240 B.n768 B.n767 10.6151
R1241 B.n770 B.n768 10.6151
R1242 B.n770 B.n769 10.6151
R1243 B.n769 B.n354 10.6151
R1244 B.n781 B.n354 10.6151
R1245 B.n782 B.n781 10.6151
R1246 B.n783 B.n782 10.6151
R1247 B.n784 B.n783 10.6151
R1248 B.n786 B.n784 10.6151
R1249 B.n787 B.n786 10.6151
R1250 B.n788 B.n787 10.6151
R1251 B.n789 B.n788 10.6151
R1252 B.n791 B.n789 10.6151
R1253 B.n792 B.n791 10.6151
R1254 B.n793 B.n792 10.6151
R1255 B.n794 B.n793 10.6151
R1256 B.n796 B.n794 10.6151
R1257 B.n797 B.n796 10.6151
R1258 B.n798 B.n797 10.6151
R1259 B.n799 B.n798 10.6151
R1260 B.n801 B.n799 10.6151
R1261 B.n802 B.n801 10.6151
R1262 B.n803 B.n802 10.6151
R1263 B.n804 B.n803 10.6151
R1264 B.n806 B.n804 10.6151
R1265 B.n807 B.n806 10.6151
R1266 B.n808 B.n807 10.6151
R1267 B.n809 B.n808 10.6151
R1268 B.n811 B.n809 10.6151
R1269 B.n812 B.n811 10.6151
R1270 B.n463 B.n397 10.6151
R1271 B.n463 B.n462 10.6151
R1272 B.n469 B.n462 10.6151
R1273 B.n470 B.n469 10.6151
R1274 B.n471 B.n470 10.6151
R1275 B.n471 B.n460 10.6151
R1276 B.n477 B.n460 10.6151
R1277 B.n478 B.n477 10.6151
R1278 B.n479 B.n478 10.6151
R1279 B.n479 B.n458 10.6151
R1280 B.n485 B.n458 10.6151
R1281 B.n486 B.n485 10.6151
R1282 B.n487 B.n486 10.6151
R1283 B.n487 B.n456 10.6151
R1284 B.n493 B.n456 10.6151
R1285 B.n494 B.n493 10.6151
R1286 B.n495 B.n494 10.6151
R1287 B.n495 B.n454 10.6151
R1288 B.n501 B.n454 10.6151
R1289 B.n502 B.n501 10.6151
R1290 B.n503 B.n502 10.6151
R1291 B.n503 B.n452 10.6151
R1292 B.n509 B.n452 10.6151
R1293 B.n510 B.n509 10.6151
R1294 B.n511 B.n510 10.6151
R1295 B.n511 B.n450 10.6151
R1296 B.n517 B.n450 10.6151
R1297 B.n518 B.n517 10.6151
R1298 B.n519 B.n518 10.6151
R1299 B.n519 B.n448 10.6151
R1300 B.n525 B.n448 10.6151
R1301 B.n526 B.n525 10.6151
R1302 B.n527 B.n526 10.6151
R1303 B.n527 B.n446 10.6151
R1304 B.n533 B.n446 10.6151
R1305 B.n534 B.n533 10.6151
R1306 B.n535 B.n534 10.6151
R1307 B.n535 B.n444 10.6151
R1308 B.n541 B.n444 10.6151
R1309 B.n542 B.n541 10.6151
R1310 B.n543 B.n542 10.6151
R1311 B.n543 B.n442 10.6151
R1312 B.n549 B.n442 10.6151
R1313 B.n550 B.n549 10.6151
R1314 B.n551 B.n550 10.6151
R1315 B.n551 B.n440 10.6151
R1316 B.n557 B.n440 10.6151
R1317 B.n558 B.n557 10.6151
R1318 B.n559 B.n558 10.6151
R1319 B.n559 B.n438 10.6151
R1320 B.n565 B.n438 10.6151
R1321 B.n566 B.n565 10.6151
R1322 B.n567 B.n566 10.6151
R1323 B.n567 B.n436 10.6151
R1324 B.n573 B.n436 10.6151
R1325 B.n576 B.n575 10.6151
R1326 B.n576 B.n432 10.6151
R1327 B.n582 B.n432 10.6151
R1328 B.n583 B.n582 10.6151
R1329 B.n584 B.n583 10.6151
R1330 B.n584 B.n430 10.6151
R1331 B.n590 B.n430 10.6151
R1332 B.n591 B.n590 10.6151
R1333 B.n595 B.n591 10.6151
R1334 B.n601 B.n428 10.6151
R1335 B.n602 B.n601 10.6151
R1336 B.n603 B.n602 10.6151
R1337 B.n603 B.n426 10.6151
R1338 B.n609 B.n426 10.6151
R1339 B.n610 B.n609 10.6151
R1340 B.n611 B.n610 10.6151
R1341 B.n611 B.n424 10.6151
R1342 B.n617 B.n424 10.6151
R1343 B.n618 B.n617 10.6151
R1344 B.n619 B.n618 10.6151
R1345 B.n619 B.n422 10.6151
R1346 B.n625 B.n422 10.6151
R1347 B.n626 B.n625 10.6151
R1348 B.n627 B.n626 10.6151
R1349 B.n627 B.n420 10.6151
R1350 B.n633 B.n420 10.6151
R1351 B.n634 B.n633 10.6151
R1352 B.n635 B.n634 10.6151
R1353 B.n635 B.n418 10.6151
R1354 B.n641 B.n418 10.6151
R1355 B.n642 B.n641 10.6151
R1356 B.n643 B.n642 10.6151
R1357 B.n643 B.n416 10.6151
R1358 B.n649 B.n416 10.6151
R1359 B.n650 B.n649 10.6151
R1360 B.n651 B.n650 10.6151
R1361 B.n651 B.n414 10.6151
R1362 B.n657 B.n414 10.6151
R1363 B.n658 B.n657 10.6151
R1364 B.n659 B.n658 10.6151
R1365 B.n659 B.n412 10.6151
R1366 B.n665 B.n412 10.6151
R1367 B.n666 B.n665 10.6151
R1368 B.n667 B.n666 10.6151
R1369 B.n667 B.n410 10.6151
R1370 B.n673 B.n410 10.6151
R1371 B.n674 B.n673 10.6151
R1372 B.n675 B.n674 10.6151
R1373 B.n675 B.n408 10.6151
R1374 B.n681 B.n408 10.6151
R1375 B.n682 B.n681 10.6151
R1376 B.n683 B.n682 10.6151
R1377 B.n683 B.n406 10.6151
R1378 B.n689 B.n406 10.6151
R1379 B.n690 B.n689 10.6151
R1380 B.n691 B.n690 10.6151
R1381 B.n691 B.n404 10.6151
R1382 B.n697 B.n404 10.6151
R1383 B.n698 B.n697 10.6151
R1384 B.n699 B.n698 10.6151
R1385 B.n699 B.n402 10.6151
R1386 B.n402 B.n401 10.6151
R1387 B.n706 B.n401 10.6151
R1388 B.n707 B.n706 10.6151
R1389 B.n713 B.n712 10.6151
R1390 B.n714 B.n713 10.6151
R1391 B.n714 B.n389 10.6151
R1392 B.n725 B.n389 10.6151
R1393 B.n726 B.n725 10.6151
R1394 B.n727 B.n726 10.6151
R1395 B.n727 B.n382 10.6151
R1396 B.n737 B.n382 10.6151
R1397 B.n738 B.n737 10.6151
R1398 B.n739 B.n738 10.6151
R1399 B.n739 B.n374 10.6151
R1400 B.n749 B.n374 10.6151
R1401 B.n750 B.n749 10.6151
R1402 B.n751 B.n750 10.6151
R1403 B.n751 B.n366 10.6151
R1404 B.n761 B.n366 10.6151
R1405 B.n762 B.n761 10.6151
R1406 B.n763 B.n762 10.6151
R1407 B.n763 B.n358 10.6151
R1408 B.n774 B.n358 10.6151
R1409 B.n775 B.n774 10.6151
R1410 B.n776 B.n775 10.6151
R1411 B.n776 B.n0 10.6151
R1412 B.n861 B.n1 10.6151
R1413 B.n861 B.n860 10.6151
R1414 B.n860 B.n859 10.6151
R1415 B.n859 B.n10 10.6151
R1416 B.n853 B.n10 10.6151
R1417 B.n853 B.n852 10.6151
R1418 B.n852 B.n851 10.6151
R1419 B.n851 B.n17 10.6151
R1420 B.n845 B.n17 10.6151
R1421 B.n845 B.n844 10.6151
R1422 B.n844 B.n843 10.6151
R1423 B.n843 B.n24 10.6151
R1424 B.n837 B.n24 10.6151
R1425 B.n837 B.n836 10.6151
R1426 B.n836 B.n835 10.6151
R1427 B.n835 B.n31 10.6151
R1428 B.n829 B.n31 10.6151
R1429 B.n829 B.n828 10.6151
R1430 B.n828 B.n827 10.6151
R1431 B.n827 B.n37 10.6151
R1432 B.n821 B.n37 10.6151
R1433 B.n821 B.n820 10.6151
R1434 B.n820 B.n819 10.6151
R1435 B.n772 B.t2 9.40856
R1436 B.n857 B.t1 9.40856
R1437 B.n223 B.n114 9.36635
R1438 B.n246 B.n111 9.36635
R1439 B.n574 B.n573 9.36635
R1440 B.n594 B.n428 9.36635
R1441 B.n729 B.t5 6.43759
R1442 B.n831 B.t9 6.43759
R1443 B.n867 B.n0 2.81026
R1444 B.n867 B.n1 2.81026
R1445 B.n226 B.n114 1.24928
R1446 B.n243 B.n111 1.24928
R1447 B.n575 B.n574 1.24928
R1448 B.n595 B.n594 1.24928
R1449 VN.n0 VN.t1 310.13
R1450 VN.n1 VN.t3 310.13
R1451 VN.n0 VN.t2 309.815
R1452 VN.n1 VN.t0 309.815
R1453 VN VN.n1 60.0265
R1454 VN VN.n0 13.1212
R1455 VDD2.n2 VDD2.n0 106.465
R1456 VDD2.n2 VDD2.n1 63.4398
R1457 VDD2.n1 VDD2.t2 1.16933
R1458 VDD2.n1 VDD2.t0 1.16933
R1459 VDD2.n0 VDD2.t3 1.16933
R1460 VDD2.n0 VDD2.t1 1.16933
R1461 VDD2 VDD2.n2 0.0586897
R1462 VTAIL.n746 VTAIL.n658 289.615
R1463 VTAIL.n88 VTAIL.n0 289.615
R1464 VTAIL.n182 VTAIL.n94 289.615
R1465 VTAIL.n276 VTAIL.n188 289.615
R1466 VTAIL.n652 VTAIL.n564 289.615
R1467 VTAIL.n558 VTAIL.n470 289.615
R1468 VTAIL.n464 VTAIL.n376 289.615
R1469 VTAIL.n370 VTAIL.n282 289.615
R1470 VTAIL.n689 VTAIL.n688 185
R1471 VTAIL.n686 VTAIL.n685 185
R1472 VTAIL.n695 VTAIL.n694 185
R1473 VTAIL.n697 VTAIL.n696 185
R1474 VTAIL.n682 VTAIL.n681 185
R1475 VTAIL.n703 VTAIL.n702 185
R1476 VTAIL.n705 VTAIL.n704 185
R1477 VTAIL.n678 VTAIL.n677 185
R1478 VTAIL.n711 VTAIL.n710 185
R1479 VTAIL.n713 VTAIL.n712 185
R1480 VTAIL.n674 VTAIL.n673 185
R1481 VTAIL.n719 VTAIL.n718 185
R1482 VTAIL.n721 VTAIL.n720 185
R1483 VTAIL.n670 VTAIL.n669 185
R1484 VTAIL.n727 VTAIL.n726 185
R1485 VTAIL.n730 VTAIL.n729 185
R1486 VTAIL.n728 VTAIL.n666 185
R1487 VTAIL.n735 VTAIL.n665 185
R1488 VTAIL.n737 VTAIL.n736 185
R1489 VTAIL.n739 VTAIL.n738 185
R1490 VTAIL.n662 VTAIL.n661 185
R1491 VTAIL.n745 VTAIL.n744 185
R1492 VTAIL.n747 VTAIL.n746 185
R1493 VTAIL.n31 VTAIL.n30 185
R1494 VTAIL.n28 VTAIL.n27 185
R1495 VTAIL.n37 VTAIL.n36 185
R1496 VTAIL.n39 VTAIL.n38 185
R1497 VTAIL.n24 VTAIL.n23 185
R1498 VTAIL.n45 VTAIL.n44 185
R1499 VTAIL.n47 VTAIL.n46 185
R1500 VTAIL.n20 VTAIL.n19 185
R1501 VTAIL.n53 VTAIL.n52 185
R1502 VTAIL.n55 VTAIL.n54 185
R1503 VTAIL.n16 VTAIL.n15 185
R1504 VTAIL.n61 VTAIL.n60 185
R1505 VTAIL.n63 VTAIL.n62 185
R1506 VTAIL.n12 VTAIL.n11 185
R1507 VTAIL.n69 VTAIL.n68 185
R1508 VTAIL.n72 VTAIL.n71 185
R1509 VTAIL.n70 VTAIL.n8 185
R1510 VTAIL.n77 VTAIL.n7 185
R1511 VTAIL.n79 VTAIL.n78 185
R1512 VTAIL.n81 VTAIL.n80 185
R1513 VTAIL.n4 VTAIL.n3 185
R1514 VTAIL.n87 VTAIL.n86 185
R1515 VTAIL.n89 VTAIL.n88 185
R1516 VTAIL.n125 VTAIL.n124 185
R1517 VTAIL.n122 VTAIL.n121 185
R1518 VTAIL.n131 VTAIL.n130 185
R1519 VTAIL.n133 VTAIL.n132 185
R1520 VTAIL.n118 VTAIL.n117 185
R1521 VTAIL.n139 VTAIL.n138 185
R1522 VTAIL.n141 VTAIL.n140 185
R1523 VTAIL.n114 VTAIL.n113 185
R1524 VTAIL.n147 VTAIL.n146 185
R1525 VTAIL.n149 VTAIL.n148 185
R1526 VTAIL.n110 VTAIL.n109 185
R1527 VTAIL.n155 VTAIL.n154 185
R1528 VTAIL.n157 VTAIL.n156 185
R1529 VTAIL.n106 VTAIL.n105 185
R1530 VTAIL.n163 VTAIL.n162 185
R1531 VTAIL.n166 VTAIL.n165 185
R1532 VTAIL.n164 VTAIL.n102 185
R1533 VTAIL.n171 VTAIL.n101 185
R1534 VTAIL.n173 VTAIL.n172 185
R1535 VTAIL.n175 VTAIL.n174 185
R1536 VTAIL.n98 VTAIL.n97 185
R1537 VTAIL.n181 VTAIL.n180 185
R1538 VTAIL.n183 VTAIL.n182 185
R1539 VTAIL.n219 VTAIL.n218 185
R1540 VTAIL.n216 VTAIL.n215 185
R1541 VTAIL.n225 VTAIL.n224 185
R1542 VTAIL.n227 VTAIL.n226 185
R1543 VTAIL.n212 VTAIL.n211 185
R1544 VTAIL.n233 VTAIL.n232 185
R1545 VTAIL.n235 VTAIL.n234 185
R1546 VTAIL.n208 VTAIL.n207 185
R1547 VTAIL.n241 VTAIL.n240 185
R1548 VTAIL.n243 VTAIL.n242 185
R1549 VTAIL.n204 VTAIL.n203 185
R1550 VTAIL.n249 VTAIL.n248 185
R1551 VTAIL.n251 VTAIL.n250 185
R1552 VTAIL.n200 VTAIL.n199 185
R1553 VTAIL.n257 VTAIL.n256 185
R1554 VTAIL.n260 VTAIL.n259 185
R1555 VTAIL.n258 VTAIL.n196 185
R1556 VTAIL.n265 VTAIL.n195 185
R1557 VTAIL.n267 VTAIL.n266 185
R1558 VTAIL.n269 VTAIL.n268 185
R1559 VTAIL.n192 VTAIL.n191 185
R1560 VTAIL.n275 VTAIL.n274 185
R1561 VTAIL.n277 VTAIL.n276 185
R1562 VTAIL.n653 VTAIL.n652 185
R1563 VTAIL.n651 VTAIL.n650 185
R1564 VTAIL.n568 VTAIL.n567 185
R1565 VTAIL.n645 VTAIL.n644 185
R1566 VTAIL.n643 VTAIL.n642 185
R1567 VTAIL.n641 VTAIL.n571 185
R1568 VTAIL.n575 VTAIL.n572 185
R1569 VTAIL.n636 VTAIL.n635 185
R1570 VTAIL.n634 VTAIL.n633 185
R1571 VTAIL.n577 VTAIL.n576 185
R1572 VTAIL.n628 VTAIL.n627 185
R1573 VTAIL.n626 VTAIL.n625 185
R1574 VTAIL.n581 VTAIL.n580 185
R1575 VTAIL.n620 VTAIL.n619 185
R1576 VTAIL.n618 VTAIL.n617 185
R1577 VTAIL.n585 VTAIL.n584 185
R1578 VTAIL.n612 VTAIL.n611 185
R1579 VTAIL.n610 VTAIL.n609 185
R1580 VTAIL.n589 VTAIL.n588 185
R1581 VTAIL.n604 VTAIL.n603 185
R1582 VTAIL.n602 VTAIL.n601 185
R1583 VTAIL.n593 VTAIL.n592 185
R1584 VTAIL.n596 VTAIL.n595 185
R1585 VTAIL.n559 VTAIL.n558 185
R1586 VTAIL.n557 VTAIL.n556 185
R1587 VTAIL.n474 VTAIL.n473 185
R1588 VTAIL.n551 VTAIL.n550 185
R1589 VTAIL.n549 VTAIL.n548 185
R1590 VTAIL.n547 VTAIL.n477 185
R1591 VTAIL.n481 VTAIL.n478 185
R1592 VTAIL.n542 VTAIL.n541 185
R1593 VTAIL.n540 VTAIL.n539 185
R1594 VTAIL.n483 VTAIL.n482 185
R1595 VTAIL.n534 VTAIL.n533 185
R1596 VTAIL.n532 VTAIL.n531 185
R1597 VTAIL.n487 VTAIL.n486 185
R1598 VTAIL.n526 VTAIL.n525 185
R1599 VTAIL.n524 VTAIL.n523 185
R1600 VTAIL.n491 VTAIL.n490 185
R1601 VTAIL.n518 VTAIL.n517 185
R1602 VTAIL.n516 VTAIL.n515 185
R1603 VTAIL.n495 VTAIL.n494 185
R1604 VTAIL.n510 VTAIL.n509 185
R1605 VTAIL.n508 VTAIL.n507 185
R1606 VTAIL.n499 VTAIL.n498 185
R1607 VTAIL.n502 VTAIL.n501 185
R1608 VTAIL.n465 VTAIL.n464 185
R1609 VTAIL.n463 VTAIL.n462 185
R1610 VTAIL.n380 VTAIL.n379 185
R1611 VTAIL.n457 VTAIL.n456 185
R1612 VTAIL.n455 VTAIL.n454 185
R1613 VTAIL.n453 VTAIL.n383 185
R1614 VTAIL.n387 VTAIL.n384 185
R1615 VTAIL.n448 VTAIL.n447 185
R1616 VTAIL.n446 VTAIL.n445 185
R1617 VTAIL.n389 VTAIL.n388 185
R1618 VTAIL.n440 VTAIL.n439 185
R1619 VTAIL.n438 VTAIL.n437 185
R1620 VTAIL.n393 VTAIL.n392 185
R1621 VTAIL.n432 VTAIL.n431 185
R1622 VTAIL.n430 VTAIL.n429 185
R1623 VTAIL.n397 VTAIL.n396 185
R1624 VTAIL.n424 VTAIL.n423 185
R1625 VTAIL.n422 VTAIL.n421 185
R1626 VTAIL.n401 VTAIL.n400 185
R1627 VTAIL.n416 VTAIL.n415 185
R1628 VTAIL.n414 VTAIL.n413 185
R1629 VTAIL.n405 VTAIL.n404 185
R1630 VTAIL.n408 VTAIL.n407 185
R1631 VTAIL.n371 VTAIL.n370 185
R1632 VTAIL.n369 VTAIL.n368 185
R1633 VTAIL.n286 VTAIL.n285 185
R1634 VTAIL.n363 VTAIL.n362 185
R1635 VTAIL.n361 VTAIL.n360 185
R1636 VTAIL.n359 VTAIL.n289 185
R1637 VTAIL.n293 VTAIL.n290 185
R1638 VTAIL.n354 VTAIL.n353 185
R1639 VTAIL.n352 VTAIL.n351 185
R1640 VTAIL.n295 VTAIL.n294 185
R1641 VTAIL.n346 VTAIL.n345 185
R1642 VTAIL.n344 VTAIL.n343 185
R1643 VTAIL.n299 VTAIL.n298 185
R1644 VTAIL.n338 VTAIL.n337 185
R1645 VTAIL.n336 VTAIL.n335 185
R1646 VTAIL.n303 VTAIL.n302 185
R1647 VTAIL.n330 VTAIL.n329 185
R1648 VTAIL.n328 VTAIL.n327 185
R1649 VTAIL.n307 VTAIL.n306 185
R1650 VTAIL.n322 VTAIL.n321 185
R1651 VTAIL.n320 VTAIL.n319 185
R1652 VTAIL.n311 VTAIL.n310 185
R1653 VTAIL.n314 VTAIL.n313 185
R1654 VTAIL.t3 VTAIL.n594 147.659
R1655 VTAIL.t1 VTAIL.n500 147.659
R1656 VTAIL.t4 VTAIL.n406 147.659
R1657 VTAIL.t7 VTAIL.n312 147.659
R1658 VTAIL.t5 VTAIL.n687 147.659
R1659 VTAIL.t6 VTAIL.n29 147.659
R1660 VTAIL.t2 VTAIL.n123 147.659
R1661 VTAIL.t0 VTAIL.n217 147.659
R1662 VTAIL.n688 VTAIL.n685 104.615
R1663 VTAIL.n695 VTAIL.n685 104.615
R1664 VTAIL.n696 VTAIL.n695 104.615
R1665 VTAIL.n696 VTAIL.n681 104.615
R1666 VTAIL.n703 VTAIL.n681 104.615
R1667 VTAIL.n704 VTAIL.n703 104.615
R1668 VTAIL.n704 VTAIL.n677 104.615
R1669 VTAIL.n711 VTAIL.n677 104.615
R1670 VTAIL.n712 VTAIL.n711 104.615
R1671 VTAIL.n712 VTAIL.n673 104.615
R1672 VTAIL.n719 VTAIL.n673 104.615
R1673 VTAIL.n720 VTAIL.n719 104.615
R1674 VTAIL.n720 VTAIL.n669 104.615
R1675 VTAIL.n727 VTAIL.n669 104.615
R1676 VTAIL.n729 VTAIL.n727 104.615
R1677 VTAIL.n729 VTAIL.n728 104.615
R1678 VTAIL.n728 VTAIL.n665 104.615
R1679 VTAIL.n737 VTAIL.n665 104.615
R1680 VTAIL.n738 VTAIL.n737 104.615
R1681 VTAIL.n738 VTAIL.n661 104.615
R1682 VTAIL.n745 VTAIL.n661 104.615
R1683 VTAIL.n746 VTAIL.n745 104.615
R1684 VTAIL.n30 VTAIL.n27 104.615
R1685 VTAIL.n37 VTAIL.n27 104.615
R1686 VTAIL.n38 VTAIL.n37 104.615
R1687 VTAIL.n38 VTAIL.n23 104.615
R1688 VTAIL.n45 VTAIL.n23 104.615
R1689 VTAIL.n46 VTAIL.n45 104.615
R1690 VTAIL.n46 VTAIL.n19 104.615
R1691 VTAIL.n53 VTAIL.n19 104.615
R1692 VTAIL.n54 VTAIL.n53 104.615
R1693 VTAIL.n54 VTAIL.n15 104.615
R1694 VTAIL.n61 VTAIL.n15 104.615
R1695 VTAIL.n62 VTAIL.n61 104.615
R1696 VTAIL.n62 VTAIL.n11 104.615
R1697 VTAIL.n69 VTAIL.n11 104.615
R1698 VTAIL.n71 VTAIL.n69 104.615
R1699 VTAIL.n71 VTAIL.n70 104.615
R1700 VTAIL.n70 VTAIL.n7 104.615
R1701 VTAIL.n79 VTAIL.n7 104.615
R1702 VTAIL.n80 VTAIL.n79 104.615
R1703 VTAIL.n80 VTAIL.n3 104.615
R1704 VTAIL.n87 VTAIL.n3 104.615
R1705 VTAIL.n88 VTAIL.n87 104.615
R1706 VTAIL.n124 VTAIL.n121 104.615
R1707 VTAIL.n131 VTAIL.n121 104.615
R1708 VTAIL.n132 VTAIL.n131 104.615
R1709 VTAIL.n132 VTAIL.n117 104.615
R1710 VTAIL.n139 VTAIL.n117 104.615
R1711 VTAIL.n140 VTAIL.n139 104.615
R1712 VTAIL.n140 VTAIL.n113 104.615
R1713 VTAIL.n147 VTAIL.n113 104.615
R1714 VTAIL.n148 VTAIL.n147 104.615
R1715 VTAIL.n148 VTAIL.n109 104.615
R1716 VTAIL.n155 VTAIL.n109 104.615
R1717 VTAIL.n156 VTAIL.n155 104.615
R1718 VTAIL.n156 VTAIL.n105 104.615
R1719 VTAIL.n163 VTAIL.n105 104.615
R1720 VTAIL.n165 VTAIL.n163 104.615
R1721 VTAIL.n165 VTAIL.n164 104.615
R1722 VTAIL.n164 VTAIL.n101 104.615
R1723 VTAIL.n173 VTAIL.n101 104.615
R1724 VTAIL.n174 VTAIL.n173 104.615
R1725 VTAIL.n174 VTAIL.n97 104.615
R1726 VTAIL.n181 VTAIL.n97 104.615
R1727 VTAIL.n182 VTAIL.n181 104.615
R1728 VTAIL.n218 VTAIL.n215 104.615
R1729 VTAIL.n225 VTAIL.n215 104.615
R1730 VTAIL.n226 VTAIL.n225 104.615
R1731 VTAIL.n226 VTAIL.n211 104.615
R1732 VTAIL.n233 VTAIL.n211 104.615
R1733 VTAIL.n234 VTAIL.n233 104.615
R1734 VTAIL.n234 VTAIL.n207 104.615
R1735 VTAIL.n241 VTAIL.n207 104.615
R1736 VTAIL.n242 VTAIL.n241 104.615
R1737 VTAIL.n242 VTAIL.n203 104.615
R1738 VTAIL.n249 VTAIL.n203 104.615
R1739 VTAIL.n250 VTAIL.n249 104.615
R1740 VTAIL.n250 VTAIL.n199 104.615
R1741 VTAIL.n257 VTAIL.n199 104.615
R1742 VTAIL.n259 VTAIL.n257 104.615
R1743 VTAIL.n259 VTAIL.n258 104.615
R1744 VTAIL.n258 VTAIL.n195 104.615
R1745 VTAIL.n267 VTAIL.n195 104.615
R1746 VTAIL.n268 VTAIL.n267 104.615
R1747 VTAIL.n268 VTAIL.n191 104.615
R1748 VTAIL.n275 VTAIL.n191 104.615
R1749 VTAIL.n276 VTAIL.n275 104.615
R1750 VTAIL.n652 VTAIL.n651 104.615
R1751 VTAIL.n651 VTAIL.n567 104.615
R1752 VTAIL.n644 VTAIL.n567 104.615
R1753 VTAIL.n644 VTAIL.n643 104.615
R1754 VTAIL.n643 VTAIL.n571 104.615
R1755 VTAIL.n575 VTAIL.n571 104.615
R1756 VTAIL.n635 VTAIL.n575 104.615
R1757 VTAIL.n635 VTAIL.n634 104.615
R1758 VTAIL.n634 VTAIL.n576 104.615
R1759 VTAIL.n627 VTAIL.n576 104.615
R1760 VTAIL.n627 VTAIL.n626 104.615
R1761 VTAIL.n626 VTAIL.n580 104.615
R1762 VTAIL.n619 VTAIL.n580 104.615
R1763 VTAIL.n619 VTAIL.n618 104.615
R1764 VTAIL.n618 VTAIL.n584 104.615
R1765 VTAIL.n611 VTAIL.n584 104.615
R1766 VTAIL.n611 VTAIL.n610 104.615
R1767 VTAIL.n610 VTAIL.n588 104.615
R1768 VTAIL.n603 VTAIL.n588 104.615
R1769 VTAIL.n603 VTAIL.n602 104.615
R1770 VTAIL.n602 VTAIL.n592 104.615
R1771 VTAIL.n595 VTAIL.n592 104.615
R1772 VTAIL.n558 VTAIL.n557 104.615
R1773 VTAIL.n557 VTAIL.n473 104.615
R1774 VTAIL.n550 VTAIL.n473 104.615
R1775 VTAIL.n550 VTAIL.n549 104.615
R1776 VTAIL.n549 VTAIL.n477 104.615
R1777 VTAIL.n481 VTAIL.n477 104.615
R1778 VTAIL.n541 VTAIL.n481 104.615
R1779 VTAIL.n541 VTAIL.n540 104.615
R1780 VTAIL.n540 VTAIL.n482 104.615
R1781 VTAIL.n533 VTAIL.n482 104.615
R1782 VTAIL.n533 VTAIL.n532 104.615
R1783 VTAIL.n532 VTAIL.n486 104.615
R1784 VTAIL.n525 VTAIL.n486 104.615
R1785 VTAIL.n525 VTAIL.n524 104.615
R1786 VTAIL.n524 VTAIL.n490 104.615
R1787 VTAIL.n517 VTAIL.n490 104.615
R1788 VTAIL.n517 VTAIL.n516 104.615
R1789 VTAIL.n516 VTAIL.n494 104.615
R1790 VTAIL.n509 VTAIL.n494 104.615
R1791 VTAIL.n509 VTAIL.n508 104.615
R1792 VTAIL.n508 VTAIL.n498 104.615
R1793 VTAIL.n501 VTAIL.n498 104.615
R1794 VTAIL.n464 VTAIL.n463 104.615
R1795 VTAIL.n463 VTAIL.n379 104.615
R1796 VTAIL.n456 VTAIL.n379 104.615
R1797 VTAIL.n456 VTAIL.n455 104.615
R1798 VTAIL.n455 VTAIL.n383 104.615
R1799 VTAIL.n387 VTAIL.n383 104.615
R1800 VTAIL.n447 VTAIL.n387 104.615
R1801 VTAIL.n447 VTAIL.n446 104.615
R1802 VTAIL.n446 VTAIL.n388 104.615
R1803 VTAIL.n439 VTAIL.n388 104.615
R1804 VTAIL.n439 VTAIL.n438 104.615
R1805 VTAIL.n438 VTAIL.n392 104.615
R1806 VTAIL.n431 VTAIL.n392 104.615
R1807 VTAIL.n431 VTAIL.n430 104.615
R1808 VTAIL.n430 VTAIL.n396 104.615
R1809 VTAIL.n423 VTAIL.n396 104.615
R1810 VTAIL.n423 VTAIL.n422 104.615
R1811 VTAIL.n422 VTAIL.n400 104.615
R1812 VTAIL.n415 VTAIL.n400 104.615
R1813 VTAIL.n415 VTAIL.n414 104.615
R1814 VTAIL.n414 VTAIL.n404 104.615
R1815 VTAIL.n407 VTAIL.n404 104.615
R1816 VTAIL.n370 VTAIL.n369 104.615
R1817 VTAIL.n369 VTAIL.n285 104.615
R1818 VTAIL.n362 VTAIL.n285 104.615
R1819 VTAIL.n362 VTAIL.n361 104.615
R1820 VTAIL.n361 VTAIL.n289 104.615
R1821 VTAIL.n293 VTAIL.n289 104.615
R1822 VTAIL.n353 VTAIL.n293 104.615
R1823 VTAIL.n353 VTAIL.n352 104.615
R1824 VTAIL.n352 VTAIL.n294 104.615
R1825 VTAIL.n345 VTAIL.n294 104.615
R1826 VTAIL.n345 VTAIL.n344 104.615
R1827 VTAIL.n344 VTAIL.n298 104.615
R1828 VTAIL.n337 VTAIL.n298 104.615
R1829 VTAIL.n337 VTAIL.n336 104.615
R1830 VTAIL.n336 VTAIL.n302 104.615
R1831 VTAIL.n329 VTAIL.n302 104.615
R1832 VTAIL.n329 VTAIL.n328 104.615
R1833 VTAIL.n328 VTAIL.n306 104.615
R1834 VTAIL.n321 VTAIL.n306 104.615
R1835 VTAIL.n321 VTAIL.n320 104.615
R1836 VTAIL.n320 VTAIL.n310 104.615
R1837 VTAIL.n313 VTAIL.n310 104.615
R1838 VTAIL.n688 VTAIL.t5 52.3082
R1839 VTAIL.n30 VTAIL.t6 52.3082
R1840 VTAIL.n124 VTAIL.t2 52.3082
R1841 VTAIL.n218 VTAIL.t0 52.3082
R1842 VTAIL.n595 VTAIL.t3 52.3082
R1843 VTAIL.n501 VTAIL.t1 52.3082
R1844 VTAIL.n407 VTAIL.t4 52.3082
R1845 VTAIL.n313 VTAIL.t7 52.3082
R1846 VTAIL.n751 VTAIL.n750 34.9005
R1847 VTAIL.n93 VTAIL.n92 34.9005
R1848 VTAIL.n187 VTAIL.n186 34.9005
R1849 VTAIL.n281 VTAIL.n280 34.9005
R1850 VTAIL.n657 VTAIL.n656 34.9005
R1851 VTAIL.n563 VTAIL.n562 34.9005
R1852 VTAIL.n469 VTAIL.n468 34.9005
R1853 VTAIL.n375 VTAIL.n374 34.9005
R1854 VTAIL.n751 VTAIL.n657 28.5393
R1855 VTAIL.n375 VTAIL.n281 28.5393
R1856 VTAIL.n689 VTAIL.n687 15.6677
R1857 VTAIL.n31 VTAIL.n29 15.6677
R1858 VTAIL.n125 VTAIL.n123 15.6677
R1859 VTAIL.n219 VTAIL.n217 15.6677
R1860 VTAIL.n596 VTAIL.n594 15.6677
R1861 VTAIL.n502 VTAIL.n500 15.6677
R1862 VTAIL.n408 VTAIL.n406 15.6677
R1863 VTAIL.n314 VTAIL.n312 15.6677
R1864 VTAIL.n736 VTAIL.n735 13.1884
R1865 VTAIL.n78 VTAIL.n77 13.1884
R1866 VTAIL.n172 VTAIL.n171 13.1884
R1867 VTAIL.n266 VTAIL.n265 13.1884
R1868 VTAIL.n642 VTAIL.n641 13.1884
R1869 VTAIL.n548 VTAIL.n547 13.1884
R1870 VTAIL.n454 VTAIL.n453 13.1884
R1871 VTAIL.n360 VTAIL.n359 13.1884
R1872 VTAIL.n690 VTAIL.n686 12.8005
R1873 VTAIL.n734 VTAIL.n666 12.8005
R1874 VTAIL.n739 VTAIL.n664 12.8005
R1875 VTAIL.n32 VTAIL.n28 12.8005
R1876 VTAIL.n76 VTAIL.n8 12.8005
R1877 VTAIL.n81 VTAIL.n6 12.8005
R1878 VTAIL.n126 VTAIL.n122 12.8005
R1879 VTAIL.n170 VTAIL.n102 12.8005
R1880 VTAIL.n175 VTAIL.n100 12.8005
R1881 VTAIL.n220 VTAIL.n216 12.8005
R1882 VTAIL.n264 VTAIL.n196 12.8005
R1883 VTAIL.n269 VTAIL.n194 12.8005
R1884 VTAIL.n645 VTAIL.n570 12.8005
R1885 VTAIL.n640 VTAIL.n572 12.8005
R1886 VTAIL.n597 VTAIL.n593 12.8005
R1887 VTAIL.n551 VTAIL.n476 12.8005
R1888 VTAIL.n546 VTAIL.n478 12.8005
R1889 VTAIL.n503 VTAIL.n499 12.8005
R1890 VTAIL.n457 VTAIL.n382 12.8005
R1891 VTAIL.n452 VTAIL.n384 12.8005
R1892 VTAIL.n409 VTAIL.n405 12.8005
R1893 VTAIL.n363 VTAIL.n288 12.8005
R1894 VTAIL.n358 VTAIL.n290 12.8005
R1895 VTAIL.n315 VTAIL.n311 12.8005
R1896 VTAIL.n694 VTAIL.n693 12.0247
R1897 VTAIL.n731 VTAIL.n730 12.0247
R1898 VTAIL.n740 VTAIL.n662 12.0247
R1899 VTAIL.n36 VTAIL.n35 12.0247
R1900 VTAIL.n73 VTAIL.n72 12.0247
R1901 VTAIL.n82 VTAIL.n4 12.0247
R1902 VTAIL.n130 VTAIL.n129 12.0247
R1903 VTAIL.n167 VTAIL.n166 12.0247
R1904 VTAIL.n176 VTAIL.n98 12.0247
R1905 VTAIL.n224 VTAIL.n223 12.0247
R1906 VTAIL.n261 VTAIL.n260 12.0247
R1907 VTAIL.n270 VTAIL.n192 12.0247
R1908 VTAIL.n646 VTAIL.n568 12.0247
R1909 VTAIL.n637 VTAIL.n636 12.0247
R1910 VTAIL.n601 VTAIL.n600 12.0247
R1911 VTAIL.n552 VTAIL.n474 12.0247
R1912 VTAIL.n543 VTAIL.n542 12.0247
R1913 VTAIL.n507 VTAIL.n506 12.0247
R1914 VTAIL.n458 VTAIL.n380 12.0247
R1915 VTAIL.n449 VTAIL.n448 12.0247
R1916 VTAIL.n413 VTAIL.n412 12.0247
R1917 VTAIL.n364 VTAIL.n286 12.0247
R1918 VTAIL.n355 VTAIL.n354 12.0247
R1919 VTAIL.n319 VTAIL.n318 12.0247
R1920 VTAIL.n697 VTAIL.n684 11.249
R1921 VTAIL.n726 VTAIL.n668 11.249
R1922 VTAIL.n744 VTAIL.n743 11.249
R1923 VTAIL.n39 VTAIL.n26 11.249
R1924 VTAIL.n68 VTAIL.n10 11.249
R1925 VTAIL.n86 VTAIL.n85 11.249
R1926 VTAIL.n133 VTAIL.n120 11.249
R1927 VTAIL.n162 VTAIL.n104 11.249
R1928 VTAIL.n180 VTAIL.n179 11.249
R1929 VTAIL.n227 VTAIL.n214 11.249
R1930 VTAIL.n256 VTAIL.n198 11.249
R1931 VTAIL.n274 VTAIL.n273 11.249
R1932 VTAIL.n650 VTAIL.n649 11.249
R1933 VTAIL.n633 VTAIL.n574 11.249
R1934 VTAIL.n604 VTAIL.n591 11.249
R1935 VTAIL.n556 VTAIL.n555 11.249
R1936 VTAIL.n539 VTAIL.n480 11.249
R1937 VTAIL.n510 VTAIL.n497 11.249
R1938 VTAIL.n462 VTAIL.n461 11.249
R1939 VTAIL.n445 VTAIL.n386 11.249
R1940 VTAIL.n416 VTAIL.n403 11.249
R1941 VTAIL.n368 VTAIL.n367 11.249
R1942 VTAIL.n351 VTAIL.n292 11.249
R1943 VTAIL.n322 VTAIL.n309 11.249
R1944 VTAIL.n698 VTAIL.n682 10.4732
R1945 VTAIL.n725 VTAIL.n670 10.4732
R1946 VTAIL.n747 VTAIL.n660 10.4732
R1947 VTAIL.n40 VTAIL.n24 10.4732
R1948 VTAIL.n67 VTAIL.n12 10.4732
R1949 VTAIL.n89 VTAIL.n2 10.4732
R1950 VTAIL.n134 VTAIL.n118 10.4732
R1951 VTAIL.n161 VTAIL.n106 10.4732
R1952 VTAIL.n183 VTAIL.n96 10.4732
R1953 VTAIL.n228 VTAIL.n212 10.4732
R1954 VTAIL.n255 VTAIL.n200 10.4732
R1955 VTAIL.n277 VTAIL.n190 10.4732
R1956 VTAIL.n653 VTAIL.n566 10.4732
R1957 VTAIL.n632 VTAIL.n577 10.4732
R1958 VTAIL.n605 VTAIL.n589 10.4732
R1959 VTAIL.n559 VTAIL.n472 10.4732
R1960 VTAIL.n538 VTAIL.n483 10.4732
R1961 VTAIL.n511 VTAIL.n495 10.4732
R1962 VTAIL.n465 VTAIL.n378 10.4732
R1963 VTAIL.n444 VTAIL.n389 10.4732
R1964 VTAIL.n417 VTAIL.n401 10.4732
R1965 VTAIL.n371 VTAIL.n284 10.4732
R1966 VTAIL.n350 VTAIL.n295 10.4732
R1967 VTAIL.n323 VTAIL.n307 10.4732
R1968 VTAIL.n702 VTAIL.n701 9.69747
R1969 VTAIL.n722 VTAIL.n721 9.69747
R1970 VTAIL.n748 VTAIL.n658 9.69747
R1971 VTAIL.n44 VTAIL.n43 9.69747
R1972 VTAIL.n64 VTAIL.n63 9.69747
R1973 VTAIL.n90 VTAIL.n0 9.69747
R1974 VTAIL.n138 VTAIL.n137 9.69747
R1975 VTAIL.n158 VTAIL.n157 9.69747
R1976 VTAIL.n184 VTAIL.n94 9.69747
R1977 VTAIL.n232 VTAIL.n231 9.69747
R1978 VTAIL.n252 VTAIL.n251 9.69747
R1979 VTAIL.n278 VTAIL.n188 9.69747
R1980 VTAIL.n654 VTAIL.n564 9.69747
R1981 VTAIL.n629 VTAIL.n628 9.69747
R1982 VTAIL.n609 VTAIL.n608 9.69747
R1983 VTAIL.n560 VTAIL.n470 9.69747
R1984 VTAIL.n535 VTAIL.n534 9.69747
R1985 VTAIL.n515 VTAIL.n514 9.69747
R1986 VTAIL.n466 VTAIL.n376 9.69747
R1987 VTAIL.n441 VTAIL.n440 9.69747
R1988 VTAIL.n421 VTAIL.n420 9.69747
R1989 VTAIL.n372 VTAIL.n282 9.69747
R1990 VTAIL.n347 VTAIL.n346 9.69747
R1991 VTAIL.n327 VTAIL.n326 9.69747
R1992 VTAIL.n750 VTAIL.n749 9.45567
R1993 VTAIL.n92 VTAIL.n91 9.45567
R1994 VTAIL.n186 VTAIL.n185 9.45567
R1995 VTAIL.n280 VTAIL.n279 9.45567
R1996 VTAIL.n656 VTAIL.n655 9.45567
R1997 VTAIL.n562 VTAIL.n561 9.45567
R1998 VTAIL.n468 VTAIL.n467 9.45567
R1999 VTAIL.n374 VTAIL.n373 9.45567
R2000 VTAIL.n749 VTAIL.n748 9.3005
R2001 VTAIL.n660 VTAIL.n659 9.3005
R2002 VTAIL.n743 VTAIL.n742 9.3005
R2003 VTAIL.n741 VTAIL.n740 9.3005
R2004 VTAIL.n664 VTAIL.n663 9.3005
R2005 VTAIL.n709 VTAIL.n708 9.3005
R2006 VTAIL.n707 VTAIL.n706 9.3005
R2007 VTAIL.n680 VTAIL.n679 9.3005
R2008 VTAIL.n701 VTAIL.n700 9.3005
R2009 VTAIL.n699 VTAIL.n698 9.3005
R2010 VTAIL.n684 VTAIL.n683 9.3005
R2011 VTAIL.n693 VTAIL.n692 9.3005
R2012 VTAIL.n691 VTAIL.n690 9.3005
R2013 VTAIL.n676 VTAIL.n675 9.3005
R2014 VTAIL.n715 VTAIL.n714 9.3005
R2015 VTAIL.n717 VTAIL.n716 9.3005
R2016 VTAIL.n672 VTAIL.n671 9.3005
R2017 VTAIL.n723 VTAIL.n722 9.3005
R2018 VTAIL.n725 VTAIL.n724 9.3005
R2019 VTAIL.n668 VTAIL.n667 9.3005
R2020 VTAIL.n732 VTAIL.n731 9.3005
R2021 VTAIL.n734 VTAIL.n733 9.3005
R2022 VTAIL.n91 VTAIL.n90 9.3005
R2023 VTAIL.n2 VTAIL.n1 9.3005
R2024 VTAIL.n85 VTAIL.n84 9.3005
R2025 VTAIL.n83 VTAIL.n82 9.3005
R2026 VTAIL.n6 VTAIL.n5 9.3005
R2027 VTAIL.n51 VTAIL.n50 9.3005
R2028 VTAIL.n49 VTAIL.n48 9.3005
R2029 VTAIL.n22 VTAIL.n21 9.3005
R2030 VTAIL.n43 VTAIL.n42 9.3005
R2031 VTAIL.n41 VTAIL.n40 9.3005
R2032 VTAIL.n26 VTAIL.n25 9.3005
R2033 VTAIL.n35 VTAIL.n34 9.3005
R2034 VTAIL.n33 VTAIL.n32 9.3005
R2035 VTAIL.n18 VTAIL.n17 9.3005
R2036 VTAIL.n57 VTAIL.n56 9.3005
R2037 VTAIL.n59 VTAIL.n58 9.3005
R2038 VTAIL.n14 VTAIL.n13 9.3005
R2039 VTAIL.n65 VTAIL.n64 9.3005
R2040 VTAIL.n67 VTAIL.n66 9.3005
R2041 VTAIL.n10 VTAIL.n9 9.3005
R2042 VTAIL.n74 VTAIL.n73 9.3005
R2043 VTAIL.n76 VTAIL.n75 9.3005
R2044 VTAIL.n185 VTAIL.n184 9.3005
R2045 VTAIL.n96 VTAIL.n95 9.3005
R2046 VTAIL.n179 VTAIL.n178 9.3005
R2047 VTAIL.n177 VTAIL.n176 9.3005
R2048 VTAIL.n100 VTAIL.n99 9.3005
R2049 VTAIL.n145 VTAIL.n144 9.3005
R2050 VTAIL.n143 VTAIL.n142 9.3005
R2051 VTAIL.n116 VTAIL.n115 9.3005
R2052 VTAIL.n137 VTAIL.n136 9.3005
R2053 VTAIL.n135 VTAIL.n134 9.3005
R2054 VTAIL.n120 VTAIL.n119 9.3005
R2055 VTAIL.n129 VTAIL.n128 9.3005
R2056 VTAIL.n127 VTAIL.n126 9.3005
R2057 VTAIL.n112 VTAIL.n111 9.3005
R2058 VTAIL.n151 VTAIL.n150 9.3005
R2059 VTAIL.n153 VTAIL.n152 9.3005
R2060 VTAIL.n108 VTAIL.n107 9.3005
R2061 VTAIL.n159 VTAIL.n158 9.3005
R2062 VTAIL.n161 VTAIL.n160 9.3005
R2063 VTAIL.n104 VTAIL.n103 9.3005
R2064 VTAIL.n168 VTAIL.n167 9.3005
R2065 VTAIL.n170 VTAIL.n169 9.3005
R2066 VTAIL.n279 VTAIL.n278 9.3005
R2067 VTAIL.n190 VTAIL.n189 9.3005
R2068 VTAIL.n273 VTAIL.n272 9.3005
R2069 VTAIL.n271 VTAIL.n270 9.3005
R2070 VTAIL.n194 VTAIL.n193 9.3005
R2071 VTAIL.n239 VTAIL.n238 9.3005
R2072 VTAIL.n237 VTAIL.n236 9.3005
R2073 VTAIL.n210 VTAIL.n209 9.3005
R2074 VTAIL.n231 VTAIL.n230 9.3005
R2075 VTAIL.n229 VTAIL.n228 9.3005
R2076 VTAIL.n214 VTAIL.n213 9.3005
R2077 VTAIL.n223 VTAIL.n222 9.3005
R2078 VTAIL.n221 VTAIL.n220 9.3005
R2079 VTAIL.n206 VTAIL.n205 9.3005
R2080 VTAIL.n245 VTAIL.n244 9.3005
R2081 VTAIL.n247 VTAIL.n246 9.3005
R2082 VTAIL.n202 VTAIL.n201 9.3005
R2083 VTAIL.n253 VTAIL.n252 9.3005
R2084 VTAIL.n255 VTAIL.n254 9.3005
R2085 VTAIL.n198 VTAIL.n197 9.3005
R2086 VTAIL.n262 VTAIL.n261 9.3005
R2087 VTAIL.n264 VTAIL.n263 9.3005
R2088 VTAIL.n622 VTAIL.n621 9.3005
R2089 VTAIL.n624 VTAIL.n623 9.3005
R2090 VTAIL.n579 VTAIL.n578 9.3005
R2091 VTAIL.n630 VTAIL.n629 9.3005
R2092 VTAIL.n632 VTAIL.n631 9.3005
R2093 VTAIL.n574 VTAIL.n573 9.3005
R2094 VTAIL.n638 VTAIL.n637 9.3005
R2095 VTAIL.n640 VTAIL.n639 9.3005
R2096 VTAIL.n655 VTAIL.n654 9.3005
R2097 VTAIL.n566 VTAIL.n565 9.3005
R2098 VTAIL.n649 VTAIL.n648 9.3005
R2099 VTAIL.n647 VTAIL.n646 9.3005
R2100 VTAIL.n570 VTAIL.n569 9.3005
R2101 VTAIL.n583 VTAIL.n582 9.3005
R2102 VTAIL.n616 VTAIL.n615 9.3005
R2103 VTAIL.n614 VTAIL.n613 9.3005
R2104 VTAIL.n587 VTAIL.n586 9.3005
R2105 VTAIL.n608 VTAIL.n607 9.3005
R2106 VTAIL.n606 VTAIL.n605 9.3005
R2107 VTAIL.n591 VTAIL.n590 9.3005
R2108 VTAIL.n600 VTAIL.n599 9.3005
R2109 VTAIL.n598 VTAIL.n597 9.3005
R2110 VTAIL.n528 VTAIL.n527 9.3005
R2111 VTAIL.n530 VTAIL.n529 9.3005
R2112 VTAIL.n485 VTAIL.n484 9.3005
R2113 VTAIL.n536 VTAIL.n535 9.3005
R2114 VTAIL.n538 VTAIL.n537 9.3005
R2115 VTAIL.n480 VTAIL.n479 9.3005
R2116 VTAIL.n544 VTAIL.n543 9.3005
R2117 VTAIL.n546 VTAIL.n545 9.3005
R2118 VTAIL.n561 VTAIL.n560 9.3005
R2119 VTAIL.n472 VTAIL.n471 9.3005
R2120 VTAIL.n555 VTAIL.n554 9.3005
R2121 VTAIL.n553 VTAIL.n552 9.3005
R2122 VTAIL.n476 VTAIL.n475 9.3005
R2123 VTAIL.n489 VTAIL.n488 9.3005
R2124 VTAIL.n522 VTAIL.n521 9.3005
R2125 VTAIL.n520 VTAIL.n519 9.3005
R2126 VTAIL.n493 VTAIL.n492 9.3005
R2127 VTAIL.n514 VTAIL.n513 9.3005
R2128 VTAIL.n512 VTAIL.n511 9.3005
R2129 VTAIL.n497 VTAIL.n496 9.3005
R2130 VTAIL.n506 VTAIL.n505 9.3005
R2131 VTAIL.n504 VTAIL.n503 9.3005
R2132 VTAIL.n434 VTAIL.n433 9.3005
R2133 VTAIL.n436 VTAIL.n435 9.3005
R2134 VTAIL.n391 VTAIL.n390 9.3005
R2135 VTAIL.n442 VTAIL.n441 9.3005
R2136 VTAIL.n444 VTAIL.n443 9.3005
R2137 VTAIL.n386 VTAIL.n385 9.3005
R2138 VTAIL.n450 VTAIL.n449 9.3005
R2139 VTAIL.n452 VTAIL.n451 9.3005
R2140 VTAIL.n467 VTAIL.n466 9.3005
R2141 VTAIL.n378 VTAIL.n377 9.3005
R2142 VTAIL.n461 VTAIL.n460 9.3005
R2143 VTAIL.n459 VTAIL.n458 9.3005
R2144 VTAIL.n382 VTAIL.n381 9.3005
R2145 VTAIL.n395 VTAIL.n394 9.3005
R2146 VTAIL.n428 VTAIL.n427 9.3005
R2147 VTAIL.n426 VTAIL.n425 9.3005
R2148 VTAIL.n399 VTAIL.n398 9.3005
R2149 VTAIL.n420 VTAIL.n419 9.3005
R2150 VTAIL.n418 VTAIL.n417 9.3005
R2151 VTAIL.n403 VTAIL.n402 9.3005
R2152 VTAIL.n412 VTAIL.n411 9.3005
R2153 VTAIL.n410 VTAIL.n409 9.3005
R2154 VTAIL.n340 VTAIL.n339 9.3005
R2155 VTAIL.n342 VTAIL.n341 9.3005
R2156 VTAIL.n297 VTAIL.n296 9.3005
R2157 VTAIL.n348 VTAIL.n347 9.3005
R2158 VTAIL.n350 VTAIL.n349 9.3005
R2159 VTAIL.n292 VTAIL.n291 9.3005
R2160 VTAIL.n356 VTAIL.n355 9.3005
R2161 VTAIL.n358 VTAIL.n357 9.3005
R2162 VTAIL.n373 VTAIL.n372 9.3005
R2163 VTAIL.n284 VTAIL.n283 9.3005
R2164 VTAIL.n367 VTAIL.n366 9.3005
R2165 VTAIL.n365 VTAIL.n364 9.3005
R2166 VTAIL.n288 VTAIL.n287 9.3005
R2167 VTAIL.n301 VTAIL.n300 9.3005
R2168 VTAIL.n334 VTAIL.n333 9.3005
R2169 VTAIL.n332 VTAIL.n331 9.3005
R2170 VTAIL.n305 VTAIL.n304 9.3005
R2171 VTAIL.n326 VTAIL.n325 9.3005
R2172 VTAIL.n324 VTAIL.n323 9.3005
R2173 VTAIL.n309 VTAIL.n308 9.3005
R2174 VTAIL.n318 VTAIL.n317 9.3005
R2175 VTAIL.n316 VTAIL.n315 9.3005
R2176 VTAIL.n705 VTAIL.n680 8.92171
R2177 VTAIL.n718 VTAIL.n672 8.92171
R2178 VTAIL.n47 VTAIL.n22 8.92171
R2179 VTAIL.n60 VTAIL.n14 8.92171
R2180 VTAIL.n141 VTAIL.n116 8.92171
R2181 VTAIL.n154 VTAIL.n108 8.92171
R2182 VTAIL.n235 VTAIL.n210 8.92171
R2183 VTAIL.n248 VTAIL.n202 8.92171
R2184 VTAIL.n625 VTAIL.n579 8.92171
R2185 VTAIL.n612 VTAIL.n587 8.92171
R2186 VTAIL.n531 VTAIL.n485 8.92171
R2187 VTAIL.n518 VTAIL.n493 8.92171
R2188 VTAIL.n437 VTAIL.n391 8.92171
R2189 VTAIL.n424 VTAIL.n399 8.92171
R2190 VTAIL.n343 VTAIL.n297 8.92171
R2191 VTAIL.n330 VTAIL.n305 8.92171
R2192 VTAIL.n706 VTAIL.n678 8.14595
R2193 VTAIL.n717 VTAIL.n674 8.14595
R2194 VTAIL.n48 VTAIL.n20 8.14595
R2195 VTAIL.n59 VTAIL.n16 8.14595
R2196 VTAIL.n142 VTAIL.n114 8.14595
R2197 VTAIL.n153 VTAIL.n110 8.14595
R2198 VTAIL.n236 VTAIL.n208 8.14595
R2199 VTAIL.n247 VTAIL.n204 8.14595
R2200 VTAIL.n624 VTAIL.n581 8.14595
R2201 VTAIL.n613 VTAIL.n585 8.14595
R2202 VTAIL.n530 VTAIL.n487 8.14595
R2203 VTAIL.n519 VTAIL.n491 8.14595
R2204 VTAIL.n436 VTAIL.n393 8.14595
R2205 VTAIL.n425 VTAIL.n397 8.14595
R2206 VTAIL.n342 VTAIL.n299 8.14595
R2207 VTAIL.n331 VTAIL.n303 8.14595
R2208 VTAIL.n710 VTAIL.n709 7.3702
R2209 VTAIL.n714 VTAIL.n713 7.3702
R2210 VTAIL.n52 VTAIL.n51 7.3702
R2211 VTAIL.n56 VTAIL.n55 7.3702
R2212 VTAIL.n146 VTAIL.n145 7.3702
R2213 VTAIL.n150 VTAIL.n149 7.3702
R2214 VTAIL.n240 VTAIL.n239 7.3702
R2215 VTAIL.n244 VTAIL.n243 7.3702
R2216 VTAIL.n621 VTAIL.n620 7.3702
R2217 VTAIL.n617 VTAIL.n616 7.3702
R2218 VTAIL.n527 VTAIL.n526 7.3702
R2219 VTAIL.n523 VTAIL.n522 7.3702
R2220 VTAIL.n433 VTAIL.n432 7.3702
R2221 VTAIL.n429 VTAIL.n428 7.3702
R2222 VTAIL.n339 VTAIL.n338 7.3702
R2223 VTAIL.n335 VTAIL.n334 7.3702
R2224 VTAIL.n710 VTAIL.n676 6.59444
R2225 VTAIL.n713 VTAIL.n676 6.59444
R2226 VTAIL.n52 VTAIL.n18 6.59444
R2227 VTAIL.n55 VTAIL.n18 6.59444
R2228 VTAIL.n146 VTAIL.n112 6.59444
R2229 VTAIL.n149 VTAIL.n112 6.59444
R2230 VTAIL.n240 VTAIL.n206 6.59444
R2231 VTAIL.n243 VTAIL.n206 6.59444
R2232 VTAIL.n620 VTAIL.n583 6.59444
R2233 VTAIL.n617 VTAIL.n583 6.59444
R2234 VTAIL.n526 VTAIL.n489 6.59444
R2235 VTAIL.n523 VTAIL.n489 6.59444
R2236 VTAIL.n432 VTAIL.n395 6.59444
R2237 VTAIL.n429 VTAIL.n395 6.59444
R2238 VTAIL.n338 VTAIL.n301 6.59444
R2239 VTAIL.n335 VTAIL.n301 6.59444
R2240 VTAIL.n709 VTAIL.n678 5.81868
R2241 VTAIL.n714 VTAIL.n674 5.81868
R2242 VTAIL.n51 VTAIL.n20 5.81868
R2243 VTAIL.n56 VTAIL.n16 5.81868
R2244 VTAIL.n145 VTAIL.n114 5.81868
R2245 VTAIL.n150 VTAIL.n110 5.81868
R2246 VTAIL.n239 VTAIL.n208 5.81868
R2247 VTAIL.n244 VTAIL.n204 5.81868
R2248 VTAIL.n621 VTAIL.n581 5.81868
R2249 VTAIL.n616 VTAIL.n585 5.81868
R2250 VTAIL.n527 VTAIL.n487 5.81868
R2251 VTAIL.n522 VTAIL.n491 5.81868
R2252 VTAIL.n433 VTAIL.n393 5.81868
R2253 VTAIL.n428 VTAIL.n397 5.81868
R2254 VTAIL.n339 VTAIL.n299 5.81868
R2255 VTAIL.n334 VTAIL.n303 5.81868
R2256 VTAIL.n706 VTAIL.n705 5.04292
R2257 VTAIL.n718 VTAIL.n717 5.04292
R2258 VTAIL.n48 VTAIL.n47 5.04292
R2259 VTAIL.n60 VTAIL.n59 5.04292
R2260 VTAIL.n142 VTAIL.n141 5.04292
R2261 VTAIL.n154 VTAIL.n153 5.04292
R2262 VTAIL.n236 VTAIL.n235 5.04292
R2263 VTAIL.n248 VTAIL.n247 5.04292
R2264 VTAIL.n625 VTAIL.n624 5.04292
R2265 VTAIL.n613 VTAIL.n612 5.04292
R2266 VTAIL.n531 VTAIL.n530 5.04292
R2267 VTAIL.n519 VTAIL.n518 5.04292
R2268 VTAIL.n437 VTAIL.n436 5.04292
R2269 VTAIL.n425 VTAIL.n424 5.04292
R2270 VTAIL.n343 VTAIL.n342 5.04292
R2271 VTAIL.n331 VTAIL.n330 5.04292
R2272 VTAIL.n598 VTAIL.n594 4.38563
R2273 VTAIL.n504 VTAIL.n500 4.38563
R2274 VTAIL.n410 VTAIL.n406 4.38563
R2275 VTAIL.n316 VTAIL.n312 4.38563
R2276 VTAIL.n691 VTAIL.n687 4.38563
R2277 VTAIL.n33 VTAIL.n29 4.38563
R2278 VTAIL.n127 VTAIL.n123 4.38563
R2279 VTAIL.n221 VTAIL.n217 4.38563
R2280 VTAIL.n702 VTAIL.n680 4.26717
R2281 VTAIL.n721 VTAIL.n672 4.26717
R2282 VTAIL.n750 VTAIL.n658 4.26717
R2283 VTAIL.n44 VTAIL.n22 4.26717
R2284 VTAIL.n63 VTAIL.n14 4.26717
R2285 VTAIL.n92 VTAIL.n0 4.26717
R2286 VTAIL.n138 VTAIL.n116 4.26717
R2287 VTAIL.n157 VTAIL.n108 4.26717
R2288 VTAIL.n186 VTAIL.n94 4.26717
R2289 VTAIL.n232 VTAIL.n210 4.26717
R2290 VTAIL.n251 VTAIL.n202 4.26717
R2291 VTAIL.n280 VTAIL.n188 4.26717
R2292 VTAIL.n656 VTAIL.n564 4.26717
R2293 VTAIL.n628 VTAIL.n579 4.26717
R2294 VTAIL.n609 VTAIL.n587 4.26717
R2295 VTAIL.n562 VTAIL.n470 4.26717
R2296 VTAIL.n534 VTAIL.n485 4.26717
R2297 VTAIL.n515 VTAIL.n493 4.26717
R2298 VTAIL.n468 VTAIL.n376 4.26717
R2299 VTAIL.n440 VTAIL.n391 4.26717
R2300 VTAIL.n421 VTAIL.n399 4.26717
R2301 VTAIL.n374 VTAIL.n282 4.26717
R2302 VTAIL.n346 VTAIL.n297 4.26717
R2303 VTAIL.n327 VTAIL.n305 4.26717
R2304 VTAIL.n701 VTAIL.n682 3.49141
R2305 VTAIL.n722 VTAIL.n670 3.49141
R2306 VTAIL.n748 VTAIL.n747 3.49141
R2307 VTAIL.n43 VTAIL.n24 3.49141
R2308 VTAIL.n64 VTAIL.n12 3.49141
R2309 VTAIL.n90 VTAIL.n89 3.49141
R2310 VTAIL.n137 VTAIL.n118 3.49141
R2311 VTAIL.n158 VTAIL.n106 3.49141
R2312 VTAIL.n184 VTAIL.n183 3.49141
R2313 VTAIL.n231 VTAIL.n212 3.49141
R2314 VTAIL.n252 VTAIL.n200 3.49141
R2315 VTAIL.n278 VTAIL.n277 3.49141
R2316 VTAIL.n654 VTAIL.n653 3.49141
R2317 VTAIL.n629 VTAIL.n577 3.49141
R2318 VTAIL.n608 VTAIL.n589 3.49141
R2319 VTAIL.n560 VTAIL.n559 3.49141
R2320 VTAIL.n535 VTAIL.n483 3.49141
R2321 VTAIL.n514 VTAIL.n495 3.49141
R2322 VTAIL.n466 VTAIL.n465 3.49141
R2323 VTAIL.n441 VTAIL.n389 3.49141
R2324 VTAIL.n420 VTAIL.n401 3.49141
R2325 VTAIL.n372 VTAIL.n371 3.49141
R2326 VTAIL.n347 VTAIL.n295 3.49141
R2327 VTAIL.n326 VTAIL.n307 3.49141
R2328 VTAIL.n698 VTAIL.n697 2.71565
R2329 VTAIL.n726 VTAIL.n725 2.71565
R2330 VTAIL.n744 VTAIL.n660 2.71565
R2331 VTAIL.n40 VTAIL.n39 2.71565
R2332 VTAIL.n68 VTAIL.n67 2.71565
R2333 VTAIL.n86 VTAIL.n2 2.71565
R2334 VTAIL.n134 VTAIL.n133 2.71565
R2335 VTAIL.n162 VTAIL.n161 2.71565
R2336 VTAIL.n180 VTAIL.n96 2.71565
R2337 VTAIL.n228 VTAIL.n227 2.71565
R2338 VTAIL.n256 VTAIL.n255 2.71565
R2339 VTAIL.n274 VTAIL.n190 2.71565
R2340 VTAIL.n650 VTAIL.n566 2.71565
R2341 VTAIL.n633 VTAIL.n632 2.71565
R2342 VTAIL.n605 VTAIL.n604 2.71565
R2343 VTAIL.n556 VTAIL.n472 2.71565
R2344 VTAIL.n539 VTAIL.n538 2.71565
R2345 VTAIL.n511 VTAIL.n510 2.71565
R2346 VTAIL.n462 VTAIL.n378 2.71565
R2347 VTAIL.n445 VTAIL.n444 2.71565
R2348 VTAIL.n417 VTAIL.n416 2.71565
R2349 VTAIL.n368 VTAIL.n284 2.71565
R2350 VTAIL.n351 VTAIL.n350 2.71565
R2351 VTAIL.n323 VTAIL.n322 2.71565
R2352 VTAIL.n694 VTAIL.n684 1.93989
R2353 VTAIL.n730 VTAIL.n668 1.93989
R2354 VTAIL.n743 VTAIL.n662 1.93989
R2355 VTAIL.n36 VTAIL.n26 1.93989
R2356 VTAIL.n72 VTAIL.n10 1.93989
R2357 VTAIL.n85 VTAIL.n4 1.93989
R2358 VTAIL.n130 VTAIL.n120 1.93989
R2359 VTAIL.n166 VTAIL.n104 1.93989
R2360 VTAIL.n179 VTAIL.n98 1.93989
R2361 VTAIL.n224 VTAIL.n214 1.93989
R2362 VTAIL.n260 VTAIL.n198 1.93989
R2363 VTAIL.n273 VTAIL.n192 1.93989
R2364 VTAIL.n649 VTAIL.n568 1.93989
R2365 VTAIL.n636 VTAIL.n574 1.93989
R2366 VTAIL.n601 VTAIL.n591 1.93989
R2367 VTAIL.n555 VTAIL.n474 1.93989
R2368 VTAIL.n542 VTAIL.n480 1.93989
R2369 VTAIL.n507 VTAIL.n497 1.93989
R2370 VTAIL.n461 VTAIL.n380 1.93989
R2371 VTAIL.n448 VTAIL.n386 1.93989
R2372 VTAIL.n413 VTAIL.n403 1.93989
R2373 VTAIL.n367 VTAIL.n286 1.93989
R2374 VTAIL.n354 VTAIL.n292 1.93989
R2375 VTAIL.n319 VTAIL.n309 1.93989
R2376 VTAIL.n469 VTAIL.n375 1.56947
R2377 VTAIL.n657 VTAIL.n563 1.56947
R2378 VTAIL.n281 VTAIL.n187 1.56947
R2379 VTAIL.n693 VTAIL.n686 1.16414
R2380 VTAIL.n731 VTAIL.n666 1.16414
R2381 VTAIL.n740 VTAIL.n739 1.16414
R2382 VTAIL.n35 VTAIL.n28 1.16414
R2383 VTAIL.n73 VTAIL.n8 1.16414
R2384 VTAIL.n82 VTAIL.n81 1.16414
R2385 VTAIL.n129 VTAIL.n122 1.16414
R2386 VTAIL.n167 VTAIL.n102 1.16414
R2387 VTAIL.n176 VTAIL.n175 1.16414
R2388 VTAIL.n223 VTAIL.n216 1.16414
R2389 VTAIL.n261 VTAIL.n196 1.16414
R2390 VTAIL.n270 VTAIL.n269 1.16414
R2391 VTAIL.n646 VTAIL.n645 1.16414
R2392 VTAIL.n637 VTAIL.n572 1.16414
R2393 VTAIL.n600 VTAIL.n593 1.16414
R2394 VTAIL.n552 VTAIL.n551 1.16414
R2395 VTAIL.n543 VTAIL.n478 1.16414
R2396 VTAIL.n506 VTAIL.n499 1.16414
R2397 VTAIL.n458 VTAIL.n457 1.16414
R2398 VTAIL.n449 VTAIL.n384 1.16414
R2399 VTAIL.n412 VTAIL.n405 1.16414
R2400 VTAIL.n364 VTAIL.n363 1.16414
R2401 VTAIL.n355 VTAIL.n290 1.16414
R2402 VTAIL.n318 VTAIL.n311 1.16414
R2403 VTAIL VTAIL.n93 0.843172
R2404 VTAIL VTAIL.n751 0.726793
R2405 VTAIL.n563 VTAIL.n469 0.470328
R2406 VTAIL.n187 VTAIL.n93 0.470328
R2407 VTAIL.n690 VTAIL.n689 0.388379
R2408 VTAIL.n735 VTAIL.n734 0.388379
R2409 VTAIL.n736 VTAIL.n664 0.388379
R2410 VTAIL.n32 VTAIL.n31 0.388379
R2411 VTAIL.n77 VTAIL.n76 0.388379
R2412 VTAIL.n78 VTAIL.n6 0.388379
R2413 VTAIL.n126 VTAIL.n125 0.388379
R2414 VTAIL.n171 VTAIL.n170 0.388379
R2415 VTAIL.n172 VTAIL.n100 0.388379
R2416 VTAIL.n220 VTAIL.n219 0.388379
R2417 VTAIL.n265 VTAIL.n264 0.388379
R2418 VTAIL.n266 VTAIL.n194 0.388379
R2419 VTAIL.n642 VTAIL.n570 0.388379
R2420 VTAIL.n641 VTAIL.n640 0.388379
R2421 VTAIL.n597 VTAIL.n596 0.388379
R2422 VTAIL.n548 VTAIL.n476 0.388379
R2423 VTAIL.n547 VTAIL.n546 0.388379
R2424 VTAIL.n503 VTAIL.n502 0.388379
R2425 VTAIL.n454 VTAIL.n382 0.388379
R2426 VTAIL.n453 VTAIL.n452 0.388379
R2427 VTAIL.n409 VTAIL.n408 0.388379
R2428 VTAIL.n360 VTAIL.n288 0.388379
R2429 VTAIL.n359 VTAIL.n358 0.388379
R2430 VTAIL.n315 VTAIL.n314 0.388379
R2431 VTAIL.n692 VTAIL.n691 0.155672
R2432 VTAIL.n692 VTAIL.n683 0.155672
R2433 VTAIL.n699 VTAIL.n683 0.155672
R2434 VTAIL.n700 VTAIL.n699 0.155672
R2435 VTAIL.n700 VTAIL.n679 0.155672
R2436 VTAIL.n707 VTAIL.n679 0.155672
R2437 VTAIL.n708 VTAIL.n707 0.155672
R2438 VTAIL.n708 VTAIL.n675 0.155672
R2439 VTAIL.n715 VTAIL.n675 0.155672
R2440 VTAIL.n716 VTAIL.n715 0.155672
R2441 VTAIL.n716 VTAIL.n671 0.155672
R2442 VTAIL.n723 VTAIL.n671 0.155672
R2443 VTAIL.n724 VTAIL.n723 0.155672
R2444 VTAIL.n724 VTAIL.n667 0.155672
R2445 VTAIL.n732 VTAIL.n667 0.155672
R2446 VTAIL.n733 VTAIL.n732 0.155672
R2447 VTAIL.n733 VTAIL.n663 0.155672
R2448 VTAIL.n741 VTAIL.n663 0.155672
R2449 VTAIL.n742 VTAIL.n741 0.155672
R2450 VTAIL.n742 VTAIL.n659 0.155672
R2451 VTAIL.n749 VTAIL.n659 0.155672
R2452 VTAIL.n34 VTAIL.n33 0.155672
R2453 VTAIL.n34 VTAIL.n25 0.155672
R2454 VTAIL.n41 VTAIL.n25 0.155672
R2455 VTAIL.n42 VTAIL.n41 0.155672
R2456 VTAIL.n42 VTAIL.n21 0.155672
R2457 VTAIL.n49 VTAIL.n21 0.155672
R2458 VTAIL.n50 VTAIL.n49 0.155672
R2459 VTAIL.n50 VTAIL.n17 0.155672
R2460 VTAIL.n57 VTAIL.n17 0.155672
R2461 VTAIL.n58 VTAIL.n57 0.155672
R2462 VTAIL.n58 VTAIL.n13 0.155672
R2463 VTAIL.n65 VTAIL.n13 0.155672
R2464 VTAIL.n66 VTAIL.n65 0.155672
R2465 VTAIL.n66 VTAIL.n9 0.155672
R2466 VTAIL.n74 VTAIL.n9 0.155672
R2467 VTAIL.n75 VTAIL.n74 0.155672
R2468 VTAIL.n75 VTAIL.n5 0.155672
R2469 VTAIL.n83 VTAIL.n5 0.155672
R2470 VTAIL.n84 VTAIL.n83 0.155672
R2471 VTAIL.n84 VTAIL.n1 0.155672
R2472 VTAIL.n91 VTAIL.n1 0.155672
R2473 VTAIL.n128 VTAIL.n127 0.155672
R2474 VTAIL.n128 VTAIL.n119 0.155672
R2475 VTAIL.n135 VTAIL.n119 0.155672
R2476 VTAIL.n136 VTAIL.n135 0.155672
R2477 VTAIL.n136 VTAIL.n115 0.155672
R2478 VTAIL.n143 VTAIL.n115 0.155672
R2479 VTAIL.n144 VTAIL.n143 0.155672
R2480 VTAIL.n144 VTAIL.n111 0.155672
R2481 VTAIL.n151 VTAIL.n111 0.155672
R2482 VTAIL.n152 VTAIL.n151 0.155672
R2483 VTAIL.n152 VTAIL.n107 0.155672
R2484 VTAIL.n159 VTAIL.n107 0.155672
R2485 VTAIL.n160 VTAIL.n159 0.155672
R2486 VTAIL.n160 VTAIL.n103 0.155672
R2487 VTAIL.n168 VTAIL.n103 0.155672
R2488 VTAIL.n169 VTAIL.n168 0.155672
R2489 VTAIL.n169 VTAIL.n99 0.155672
R2490 VTAIL.n177 VTAIL.n99 0.155672
R2491 VTAIL.n178 VTAIL.n177 0.155672
R2492 VTAIL.n178 VTAIL.n95 0.155672
R2493 VTAIL.n185 VTAIL.n95 0.155672
R2494 VTAIL.n222 VTAIL.n221 0.155672
R2495 VTAIL.n222 VTAIL.n213 0.155672
R2496 VTAIL.n229 VTAIL.n213 0.155672
R2497 VTAIL.n230 VTAIL.n229 0.155672
R2498 VTAIL.n230 VTAIL.n209 0.155672
R2499 VTAIL.n237 VTAIL.n209 0.155672
R2500 VTAIL.n238 VTAIL.n237 0.155672
R2501 VTAIL.n238 VTAIL.n205 0.155672
R2502 VTAIL.n245 VTAIL.n205 0.155672
R2503 VTAIL.n246 VTAIL.n245 0.155672
R2504 VTAIL.n246 VTAIL.n201 0.155672
R2505 VTAIL.n253 VTAIL.n201 0.155672
R2506 VTAIL.n254 VTAIL.n253 0.155672
R2507 VTAIL.n254 VTAIL.n197 0.155672
R2508 VTAIL.n262 VTAIL.n197 0.155672
R2509 VTAIL.n263 VTAIL.n262 0.155672
R2510 VTAIL.n263 VTAIL.n193 0.155672
R2511 VTAIL.n271 VTAIL.n193 0.155672
R2512 VTAIL.n272 VTAIL.n271 0.155672
R2513 VTAIL.n272 VTAIL.n189 0.155672
R2514 VTAIL.n279 VTAIL.n189 0.155672
R2515 VTAIL.n655 VTAIL.n565 0.155672
R2516 VTAIL.n648 VTAIL.n565 0.155672
R2517 VTAIL.n648 VTAIL.n647 0.155672
R2518 VTAIL.n647 VTAIL.n569 0.155672
R2519 VTAIL.n639 VTAIL.n569 0.155672
R2520 VTAIL.n639 VTAIL.n638 0.155672
R2521 VTAIL.n638 VTAIL.n573 0.155672
R2522 VTAIL.n631 VTAIL.n573 0.155672
R2523 VTAIL.n631 VTAIL.n630 0.155672
R2524 VTAIL.n630 VTAIL.n578 0.155672
R2525 VTAIL.n623 VTAIL.n578 0.155672
R2526 VTAIL.n623 VTAIL.n622 0.155672
R2527 VTAIL.n622 VTAIL.n582 0.155672
R2528 VTAIL.n615 VTAIL.n582 0.155672
R2529 VTAIL.n615 VTAIL.n614 0.155672
R2530 VTAIL.n614 VTAIL.n586 0.155672
R2531 VTAIL.n607 VTAIL.n586 0.155672
R2532 VTAIL.n607 VTAIL.n606 0.155672
R2533 VTAIL.n606 VTAIL.n590 0.155672
R2534 VTAIL.n599 VTAIL.n590 0.155672
R2535 VTAIL.n599 VTAIL.n598 0.155672
R2536 VTAIL.n561 VTAIL.n471 0.155672
R2537 VTAIL.n554 VTAIL.n471 0.155672
R2538 VTAIL.n554 VTAIL.n553 0.155672
R2539 VTAIL.n553 VTAIL.n475 0.155672
R2540 VTAIL.n545 VTAIL.n475 0.155672
R2541 VTAIL.n545 VTAIL.n544 0.155672
R2542 VTAIL.n544 VTAIL.n479 0.155672
R2543 VTAIL.n537 VTAIL.n479 0.155672
R2544 VTAIL.n537 VTAIL.n536 0.155672
R2545 VTAIL.n536 VTAIL.n484 0.155672
R2546 VTAIL.n529 VTAIL.n484 0.155672
R2547 VTAIL.n529 VTAIL.n528 0.155672
R2548 VTAIL.n528 VTAIL.n488 0.155672
R2549 VTAIL.n521 VTAIL.n488 0.155672
R2550 VTAIL.n521 VTAIL.n520 0.155672
R2551 VTAIL.n520 VTAIL.n492 0.155672
R2552 VTAIL.n513 VTAIL.n492 0.155672
R2553 VTAIL.n513 VTAIL.n512 0.155672
R2554 VTAIL.n512 VTAIL.n496 0.155672
R2555 VTAIL.n505 VTAIL.n496 0.155672
R2556 VTAIL.n505 VTAIL.n504 0.155672
R2557 VTAIL.n467 VTAIL.n377 0.155672
R2558 VTAIL.n460 VTAIL.n377 0.155672
R2559 VTAIL.n460 VTAIL.n459 0.155672
R2560 VTAIL.n459 VTAIL.n381 0.155672
R2561 VTAIL.n451 VTAIL.n381 0.155672
R2562 VTAIL.n451 VTAIL.n450 0.155672
R2563 VTAIL.n450 VTAIL.n385 0.155672
R2564 VTAIL.n443 VTAIL.n385 0.155672
R2565 VTAIL.n443 VTAIL.n442 0.155672
R2566 VTAIL.n442 VTAIL.n390 0.155672
R2567 VTAIL.n435 VTAIL.n390 0.155672
R2568 VTAIL.n435 VTAIL.n434 0.155672
R2569 VTAIL.n434 VTAIL.n394 0.155672
R2570 VTAIL.n427 VTAIL.n394 0.155672
R2571 VTAIL.n427 VTAIL.n426 0.155672
R2572 VTAIL.n426 VTAIL.n398 0.155672
R2573 VTAIL.n419 VTAIL.n398 0.155672
R2574 VTAIL.n419 VTAIL.n418 0.155672
R2575 VTAIL.n418 VTAIL.n402 0.155672
R2576 VTAIL.n411 VTAIL.n402 0.155672
R2577 VTAIL.n411 VTAIL.n410 0.155672
R2578 VTAIL.n373 VTAIL.n283 0.155672
R2579 VTAIL.n366 VTAIL.n283 0.155672
R2580 VTAIL.n366 VTAIL.n365 0.155672
R2581 VTAIL.n365 VTAIL.n287 0.155672
R2582 VTAIL.n357 VTAIL.n287 0.155672
R2583 VTAIL.n357 VTAIL.n356 0.155672
R2584 VTAIL.n356 VTAIL.n291 0.155672
R2585 VTAIL.n349 VTAIL.n291 0.155672
R2586 VTAIL.n349 VTAIL.n348 0.155672
R2587 VTAIL.n348 VTAIL.n296 0.155672
R2588 VTAIL.n341 VTAIL.n296 0.155672
R2589 VTAIL.n341 VTAIL.n340 0.155672
R2590 VTAIL.n340 VTAIL.n300 0.155672
R2591 VTAIL.n333 VTAIL.n300 0.155672
R2592 VTAIL.n333 VTAIL.n332 0.155672
R2593 VTAIL.n332 VTAIL.n304 0.155672
R2594 VTAIL.n325 VTAIL.n304 0.155672
R2595 VTAIL.n325 VTAIL.n324 0.155672
R2596 VTAIL.n324 VTAIL.n308 0.155672
R2597 VTAIL.n317 VTAIL.n308 0.155672
R2598 VTAIL.n317 VTAIL.n316 0.155672
R2599 VP.n2 VP.t0 310.13
R2600 VP.n2 VP.t2 309.815
R2601 VP.n4 VP.t3 273.997
R2602 VP.n11 VP.t1 273.997
R2603 VP.n4 VP.n3 177.855
R2604 VP.n12 VP.n11 177.855
R2605 VP.n10 VP.n0 161.3
R2606 VP.n9 VP.n8 161.3
R2607 VP.n7 VP.n1 161.3
R2608 VP.n6 VP.n5 161.3
R2609 VP.n3 VP.n2 59.6458
R2610 VP.n9 VP.n1 56.4773
R2611 VP.n5 VP.n1 24.3439
R2612 VP.n10 VP.n9 24.3439
R2613 VP.n5 VP.n4 7.7904
R2614 VP.n11 VP.n10 7.7904
R2615 VP.n6 VP.n3 0.189894
R2616 VP.n7 VP.n6 0.189894
R2617 VP.n8 VP.n7 0.189894
R2618 VP.n8 VP.n0 0.189894
R2619 VP.n12 VP.n0 0.189894
R2620 VP VP.n12 0.0516364
R2621 VDD1 VDD1.n1 106.99
R2622 VDD1 VDD1.n0 63.498
R2623 VDD1.n0 VDD1.t3 1.16933
R2624 VDD1.n0 VDD1.t1 1.16933
R2625 VDD1.n1 VDD1.t0 1.16933
R2626 VDD1.n1 VDD1.t2 1.16933
C0 VP VN 6.31034f
C1 VDD1 VTAIL 7.0317f
C2 VDD2 VTAIL 7.07846f
C3 VP VTAIL 5.32807f
C4 VN VTAIL 5.31397f
C5 VDD1 VDD2 0.757267f
C6 VDD1 VP 5.9466f
C7 VDD2 VP 0.323459f
C8 VDD1 VN 0.147781f
C9 VDD2 VN 5.771379f
C10 VDD2 B 3.53176f
C11 VDD1 B 7.82473f
C12 VTAIL B 12.301917f
C13 VN B 9.33837f
C14 VP B 6.901174f
C15 VDD1.t3 B 0.35523f
C16 VDD1.t1 B 0.35523f
C17 VDD1.n0 B 3.23165f
C18 VDD1.t0 B 0.35523f
C19 VDD1.t2 B 0.35523f
C20 VDD1.n1 B 4.02922f
C21 VP.n0 B 0.034755f
C22 VP.t1 B 2.41006f
C23 VP.n1 B 0.050957f
C24 VP.t0 B 2.52551f
C25 VP.t2 B 2.52448f
C26 VP.n2 B 3.27345f
C27 VP.n3 B 2.14185f
C28 VP.t3 B 2.41006f
C29 VP.n4 B 0.919406f
C30 VP.n5 B 0.043243f
C31 VP.n6 B 0.034755f
C32 VP.n7 B 0.034755f
C33 VP.n8 B 0.034755f
C34 VP.n9 B 0.050957f
C35 VP.n10 B 0.043243f
C36 VP.n11 B 0.919406f
C37 VP.n12 B 0.03389f
C38 VTAIL.n0 B 0.021915f
C39 VTAIL.n1 B 0.015155f
C40 VTAIL.n2 B 0.008144f
C41 VTAIL.n3 B 0.019249f
C42 VTAIL.n4 B 0.008623f
C43 VTAIL.n5 B 0.015155f
C44 VTAIL.n6 B 0.008144f
C45 VTAIL.n7 B 0.019249f
C46 VTAIL.n8 B 0.008623f
C47 VTAIL.n9 B 0.015155f
C48 VTAIL.n10 B 0.008144f
C49 VTAIL.n11 B 0.019249f
C50 VTAIL.n12 B 0.008623f
C51 VTAIL.n13 B 0.015155f
C52 VTAIL.n14 B 0.008144f
C53 VTAIL.n15 B 0.019249f
C54 VTAIL.n16 B 0.008623f
C55 VTAIL.n17 B 0.015155f
C56 VTAIL.n18 B 0.008144f
C57 VTAIL.n19 B 0.019249f
C58 VTAIL.n20 B 0.008623f
C59 VTAIL.n21 B 0.015155f
C60 VTAIL.n22 B 0.008144f
C61 VTAIL.n23 B 0.019249f
C62 VTAIL.n24 B 0.008623f
C63 VTAIL.n25 B 0.015155f
C64 VTAIL.n26 B 0.008144f
C65 VTAIL.n27 B 0.019249f
C66 VTAIL.n28 B 0.008623f
C67 VTAIL.n29 B 0.106215f
C68 VTAIL.t6 B 0.031839f
C69 VTAIL.n30 B 0.014436f
C70 VTAIL.n31 B 0.011371f
C71 VTAIL.n32 B 0.008144f
C72 VTAIL.n33 B 1.12075f
C73 VTAIL.n34 B 0.015155f
C74 VTAIL.n35 B 0.008144f
C75 VTAIL.n36 B 0.008623f
C76 VTAIL.n37 B 0.019249f
C77 VTAIL.n38 B 0.019249f
C78 VTAIL.n39 B 0.008623f
C79 VTAIL.n40 B 0.008144f
C80 VTAIL.n41 B 0.015155f
C81 VTAIL.n42 B 0.015155f
C82 VTAIL.n43 B 0.008144f
C83 VTAIL.n44 B 0.008623f
C84 VTAIL.n45 B 0.019249f
C85 VTAIL.n46 B 0.019249f
C86 VTAIL.n47 B 0.008623f
C87 VTAIL.n48 B 0.008144f
C88 VTAIL.n49 B 0.015155f
C89 VTAIL.n50 B 0.015155f
C90 VTAIL.n51 B 0.008144f
C91 VTAIL.n52 B 0.008623f
C92 VTAIL.n53 B 0.019249f
C93 VTAIL.n54 B 0.019249f
C94 VTAIL.n55 B 0.008623f
C95 VTAIL.n56 B 0.008144f
C96 VTAIL.n57 B 0.015155f
C97 VTAIL.n58 B 0.015155f
C98 VTAIL.n59 B 0.008144f
C99 VTAIL.n60 B 0.008623f
C100 VTAIL.n61 B 0.019249f
C101 VTAIL.n62 B 0.019249f
C102 VTAIL.n63 B 0.008623f
C103 VTAIL.n64 B 0.008144f
C104 VTAIL.n65 B 0.015155f
C105 VTAIL.n66 B 0.015155f
C106 VTAIL.n67 B 0.008144f
C107 VTAIL.n68 B 0.008623f
C108 VTAIL.n69 B 0.019249f
C109 VTAIL.n70 B 0.019249f
C110 VTAIL.n71 B 0.019249f
C111 VTAIL.n72 B 0.008623f
C112 VTAIL.n73 B 0.008144f
C113 VTAIL.n74 B 0.015155f
C114 VTAIL.n75 B 0.015155f
C115 VTAIL.n76 B 0.008144f
C116 VTAIL.n77 B 0.008383f
C117 VTAIL.n78 B 0.008383f
C118 VTAIL.n79 B 0.019249f
C119 VTAIL.n80 B 0.019249f
C120 VTAIL.n81 B 0.008623f
C121 VTAIL.n82 B 0.008144f
C122 VTAIL.n83 B 0.015155f
C123 VTAIL.n84 B 0.015155f
C124 VTAIL.n85 B 0.008144f
C125 VTAIL.n86 B 0.008623f
C126 VTAIL.n87 B 0.019249f
C127 VTAIL.n88 B 0.042755f
C128 VTAIL.n89 B 0.008623f
C129 VTAIL.n90 B 0.008144f
C130 VTAIL.n91 B 0.037928f
C131 VTAIL.n92 B 0.02412f
C132 VTAIL.n93 B 0.078675f
C133 VTAIL.n94 B 0.021915f
C134 VTAIL.n95 B 0.015155f
C135 VTAIL.n96 B 0.008144f
C136 VTAIL.n97 B 0.019249f
C137 VTAIL.n98 B 0.008623f
C138 VTAIL.n99 B 0.015155f
C139 VTAIL.n100 B 0.008144f
C140 VTAIL.n101 B 0.019249f
C141 VTAIL.n102 B 0.008623f
C142 VTAIL.n103 B 0.015155f
C143 VTAIL.n104 B 0.008144f
C144 VTAIL.n105 B 0.019249f
C145 VTAIL.n106 B 0.008623f
C146 VTAIL.n107 B 0.015155f
C147 VTAIL.n108 B 0.008144f
C148 VTAIL.n109 B 0.019249f
C149 VTAIL.n110 B 0.008623f
C150 VTAIL.n111 B 0.015155f
C151 VTAIL.n112 B 0.008144f
C152 VTAIL.n113 B 0.019249f
C153 VTAIL.n114 B 0.008623f
C154 VTAIL.n115 B 0.015155f
C155 VTAIL.n116 B 0.008144f
C156 VTAIL.n117 B 0.019249f
C157 VTAIL.n118 B 0.008623f
C158 VTAIL.n119 B 0.015155f
C159 VTAIL.n120 B 0.008144f
C160 VTAIL.n121 B 0.019249f
C161 VTAIL.n122 B 0.008623f
C162 VTAIL.n123 B 0.106215f
C163 VTAIL.t2 B 0.031839f
C164 VTAIL.n124 B 0.014436f
C165 VTAIL.n125 B 0.011371f
C166 VTAIL.n126 B 0.008144f
C167 VTAIL.n127 B 1.12075f
C168 VTAIL.n128 B 0.015155f
C169 VTAIL.n129 B 0.008144f
C170 VTAIL.n130 B 0.008623f
C171 VTAIL.n131 B 0.019249f
C172 VTAIL.n132 B 0.019249f
C173 VTAIL.n133 B 0.008623f
C174 VTAIL.n134 B 0.008144f
C175 VTAIL.n135 B 0.015155f
C176 VTAIL.n136 B 0.015155f
C177 VTAIL.n137 B 0.008144f
C178 VTAIL.n138 B 0.008623f
C179 VTAIL.n139 B 0.019249f
C180 VTAIL.n140 B 0.019249f
C181 VTAIL.n141 B 0.008623f
C182 VTAIL.n142 B 0.008144f
C183 VTAIL.n143 B 0.015155f
C184 VTAIL.n144 B 0.015155f
C185 VTAIL.n145 B 0.008144f
C186 VTAIL.n146 B 0.008623f
C187 VTAIL.n147 B 0.019249f
C188 VTAIL.n148 B 0.019249f
C189 VTAIL.n149 B 0.008623f
C190 VTAIL.n150 B 0.008144f
C191 VTAIL.n151 B 0.015155f
C192 VTAIL.n152 B 0.015155f
C193 VTAIL.n153 B 0.008144f
C194 VTAIL.n154 B 0.008623f
C195 VTAIL.n155 B 0.019249f
C196 VTAIL.n156 B 0.019249f
C197 VTAIL.n157 B 0.008623f
C198 VTAIL.n158 B 0.008144f
C199 VTAIL.n159 B 0.015155f
C200 VTAIL.n160 B 0.015155f
C201 VTAIL.n161 B 0.008144f
C202 VTAIL.n162 B 0.008623f
C203 VTAIL.n163 B 0.019249f
C204 VTAIL.n164 B 0.019249f
C205 VTAIL.n165 B 0.019249f
C206 VTAIL.n166 B 0.008623f
C207 VTAIL.n167 B 0.008144f
C208 VTAIL.n168 B 0.015155f
C209 VTAIL.n169 B 0.015155f
C210 VTAIL.n170 B 0.008144f
C211 VTAIL.n171 B 0.008383f
C212 VTAIL.n172 B 0.008383f
C213 VTAIL.n173 B 0.019249f
C214 VTAIL.n174 B 0.019249f
C215 VTAIL.n175 B 0.008623f
C216 VTAIL.n176 B 0.008144f
C217 VTAIL.n177 B 0.015155f
C218 VTAIL.n178 B 0.015155f
C219 VTAIL.n179 B 0.008144f
C220 VTAIL.n180 B 0.008623f
C221 VTAIL.n181 B 0.019249f
C222 VTAIL.n182 B 0.042755f
C223 VTAIL.n183 B 0.008623f
C224 VTAIL.n184 B 0.008144f
C225 VTAIL.n185 B 0.037928f
C226 VTAIL.n186 B 0.02412f
C227 VTAIL.n187 B 0.114142f
C228 VTAIL.n188 B 0.021915f
C229 VTAIL.n189 B 0.015155f
C230 VTAIL.n190 B 0.008144f
C231 VTAIL.n191 B 0.019249f
C232 VTAIL.n192 B 0.008623f
C233 VTAIL.n193 B 0.015155f
C234 VTAIL.n194 B 0.008144f
C235 VTAIL.n195 B 0.019249f
C236 VTAIL.n196 B 0.008623f
C237 VTAIL.n197 B 0.015155f
C238 VTAIL.n198 B 0.008144f
C239 VTAIL.n199 B 0.019249f
C240 VTAIL.n200 B 0.008623f
C241 VTAIL.n201 B 0.015155f
C242 VTAIL.n202 B 0.008144f
C243 VTAIL.n203 B 0.019249f
C244 VTAIL.n204 B 0.008623f
C245 VTAIL.n205 B 0.015155f
C246 VTAIL.n206 B 0.008144f
C247 VTAIL.n207 B 0.019249f
C248 VTAIL.n208 B 0.008623f
C249 VTAIL.n209 B 0.015155f
C250 VTAIL.n210 B 0.008144f
C251 VTAIL.n211 B 0.019249f
C252 VTAIL.n212 B 0.008623f
C253 VTAIL.n213 B 0.015155f
C254 VTAIL.n214 B 0.008144f
C255 VTAIL.n215 B 0.019249f
C256 VTAIL.n216 B 0.008623f
C257 VTAIL.n217 B 0.106215f
C258 VTAIL.t0 B 0.031839f
C259 VTAIL.n218 B 0.014436f
C260 VTAIL.n219 B 0.011371f
C261 VTAIL.n220 B 0.008144f
C262 VTAIL.n221 B 1.12075f
C263 VTAIL.n222 B 0.015155f
C264 VTAIL.n223 B 0.008144f
C265 VTAIL.n224 B 0.008623f
C266 VTAIL.n225 B 0.019249f
C267 VTAIL.n226 B 0.019249f
C268 VTAIL.n227 B 0.008623f
C269 VTAIL.n228 B 0.008144f
C270 VTAIL.n229 B 0.015155f
C271 VTAIL.n230 B 0.015155f
C272 VTAIL.n231 B 0.008144f
C273 VTAIL.n232 B 0.008623f
C274 VTAIL.n233 B 0.019249f
C275 VTAIL.n234 B 0.019249f
C276 VTAIL.n235 B 0.008623f
C277 VTAIL.n236 B 0.008144f
C278 VTAIL.n237 B 0.015155f
C279 VTAIL.n238 B 0.015155f
C280 VTAIL.n239 B 0.008144f
C281 VTAIL.n240 B 0.008623f
C282 VTAIL.n241 B 0.019249f
C283 VTAIL.n242 B 0.019249f
C284 VTAIL.n243 B 0.008623f
C285 VTAIL.n244 B 0.008144f
C286 VTAIL.n245 B 0.015155f
C287 VTAIL.n246 B 0.015155f
C288 VTAIL.n247 B 0.008144f
C289 VTAIL.n248 B 0.008623f
C290 VTAIL.n249 B 0.019249f
C291 VTAIL.n250 B 0.019249f
C292 VTAIL.n251 B 0.008623f
C293 VTAIL.n252 B 0.008144f
C294 VTAIL.n253 B 0.015155f
C295 VTAIL.n254 B 0.015155f
C296 VTAIL.n255 B 0.008144f
C297 VTAIL.n256 B 0.008623f
C298 VTAIL.n257 B 0.019249f
C299 VTAIL.n258 B 0.019249f
C300 VTAIL.n259 B 0.019249f
C301 VTAIL.n260 B 0.008623f
C302 VTAIL.n261 B 0.008144f
C303 VTAIL.n262 B 0.015155f
C304 VTAIL.n263 B 0.015155f
C305 VTAIL.n264 B 0.008144f
C306 VTAIL.n265 B 0.008383f
C307 VTAIL.n266 B 0.008383f
C308 VTAIL.n267 B 0.019249f
C309 VTAIL.n268 B 0.019249f
C310 VTAIL.n269 B 0.008623f
C311 VTAIL.n270 B 0.008144f
C312 VTAIL.n271 B 0.015155f
C313 VTAIL.n272 B 0.015155f
C314 VTAIL.n273 B 0.008144f
C315 VTAIL.n274 B 0.008623f
C316 VTAIL.n275 B 0.019249f
C317 VTAIL.n276 B 0.042755f
C318 VTAIL.n277 B 0.008623f
C319 VTAIL.n278 B 0.008144f
C320 VTAIL.n279 B 0.037928f
C321 VTAIL.n280 B 0.02412f
C322 VTAIL.n281 B 1.0868f
C323 VTAIL.n282 B 0.021915f
C324 VTAIL.n283 B 0.015155f
C325 VTAIL.n284 B 0.008144f
C326 VTAIL.n285 B 0.019249f
C327 VTAIL.n286 B 0.008623f
C328 VTAIL.n287 B 0.015155f
C329 VTAIL.n288 B 0.008144f
C330 VTAIL.n289 B 0.019249f
C331 VTAIL.n290 B 0.008623f
C332 VTAIL.n291 B 0.015155f
C333 VTAIL.n292 B 0.008144f
C334 VTAIL.n293 B 0.019249f
C335 VTAIL.n294 B 0.019249f
C336 VTAIL.n295 B 0.008623f
C337 VTAIL.n296 B 0.015155f
C338 VTAIL.n297 B 0.008144f
C339 VTAIL.n298 B 0.019249f
C340 VTAIL.n299 B 0.008623f
C341 VTAIL.n300 B 0.015155f
C342 VTAIL.n301 B 0.008144f
C343 VTAIL.n302 B 0.019249f
C344 VTAIL.n303 B 0.008623f
C345 VTAIL.n304 B 0.015155f
C346 VTAIL.n305 B 0.008144f
C347 VTAIL.n306 B 0.019249f
C348 VTAIL.n307 B 0.008623f
C349 VTAIL.n308 B 0.015155f
C350 VTAIL.n309 B 0.008144f
C351 VTAIL.n310 B 0.019249f
C352 VTAIL.n311 B 0.008623f
C353 VTAIL.n312 B 0.106215f
C354 VTAIL.t7 B 0.031839f
C355 VTAIL.n313 B 0.014436f
C356 VTAIL.n314 B 0.011371f
C357 VTAIL.n315 B 0.008144f
C358 VTAIL.n316 B 1.12075f
C359 VTAIL.n317 B 0.015155f
C360 VTAIL.n318 B 0.008144f
C361 VTAIL.n319 B 0.008623f
C362 VTAIL.n320 B 0.019249f
C363 VTAIL.n321 B 0.019249f
C364 VTAIL.n322 B 0.008623f
C365 VTAIL.n323 B 0.008144f
C366 VTAIL.n324 B 0.015155f
C367 VTAIL.n325 B 0.015155f
C368 VTAIL.n326 B 0.008144f
C369 VTAIL.n327 B 0.008623f
C370 VTAIL.n328 B 0.019249f
C371 VTAIL.n329 B 0.019249f
C372 VTAIL.n330 B 0.008623f
C373 VTAIL.n331 B 0.008144f
C374 VTAIL.n332 B 0.015155f
C375 VTAIL.n333 B 0.015155f
C376 VTAIL.n334 B 0.008144f
C377 VTAIL.n335 B 0.008623f
C378 VTAIL.n336 B 0.019249f
C379 VTAIL.n337 B 0.019249f
C380 VTAIL.n338 B 0.008623f
C381 VTAIL.n339 B 0.008144f
C382 VTAIL.n340 B 0.015155f
C383 VTAIL.n341 B 0.015155f
C384 VTAIL.n342 B 0.008144f
C385 VTAIL.n343 B 0.008623f
C386 VTAIL.n344 B 0.019249f
C387 VTAIL.n345 B 0.019249f
C388 VTAIL.n346 B 0.008623f
C389 VTAIL.n347 B 0.008144f
C390 VTAIL.n348 B 0.015155f
C391 VTAIL.n349 B 0.015155f
C392 VTAIL.n350 B 0.008144f
C393 VTAIL.n351 B 0.008623f
C394 VTAIL.n352 B 0.019249f
C395 VTAIL.n353 B 0.019249f
C396 VTAIL.n354 B 0.008623f
C397 VTAIL.n355 B 0.008144f
C398 VTAIL.n356 B 0.015155f
C399 VTAIL.n357 B 0.015155f
C400 VTAIL.n358 B 0.008144f
C401 VTAIL.n359 B 0.008383f
C402 VTAIL.n360 B 0.008383f
C403 VTAIL.n361 B 0.019249f
C404 VTAIL.n362 B 0.019249f
C405 VTAIL.n363 B 0.008623f
C406 VTAIL.n364 B 0.008144f
C407 VTAIL.n365 B 0.015155f
C408 VTAIL.n366 B 0.015155f
C409 VTAIL.n367 B 0.008144f
C410 VTAIL.n368 B 0.008623f
C411 VTAIL.n369 B 0.019249f
C412 VTAIL.n370 B 0.042755f
C413 VTAIL.n371 B 0.008623f
C414 VTAIL.n372 B 0.008144f
C415 VTAIL.n373 B 0.037928f
C416 VTAIL.n374 B 0.02412f
C417 VTAIL.n375 B 1.0868f
C418 VTAIL.n376 B 0.021915f
C419 VTAIL.n377 B 0.015155f
C420 VTAIL.n378 B 0.008144f
C421 VTAIL.n379 B 0.019249f
C422 VTAIL.n380 B 0.008623f
C423 VTAIL.n381 B 0.015155f
C424 VTAIL.n382 B 0.008144f
C425 VTAIL.n383 B 0.019249f
C426 VTAIL.n384 B 0.008623f
C427 VTAIL.n385 B 0.015155f
C428 VTAIL.n386 B 0.008144f
C429 VTAIL.n387 B 0.019249f
C430 VTAIL.n388 B 0.019249f
C431 VTAIL.n389 B 0.008623f
C432 VTAIL.n390 B 0.015155f
C433 VTAIL.n391 B 0.008144f
C434 VTAIL.n392 B 0.019249f
C435 VTAIL.n393 B 0.008623f
C436 VTAIL.n394 B 0.015155f
C437 VTAIL.n395 B 0.008144f
C438 VTAIL.n396 B 0.019249f
C439 VTAIL.n397 B 0.008623f
C440 VTAIL.n398 B 0.015155f
C441 VTAIL.n399 B 0.008144f
C442 VTAIL.n400 B 0.019249f
C443 VTAIL.n401 B 0.008623f
C444 VTAIL.n402 B 0.015155f
C445 VTAIL.n403 B 0.008144f
C446 VTAIL.n404 B 0.019249f
C447 VTAIL.n405 B 0.008623f
C448 VTAIL.n406 B 0.106215f
C449 VTAIL.t4 B 0.031839f
C450 VTAIL.n407 B 0.014436f
C451 VTAIL.n408 B 0.011371f
C452 VTAIL.n409 B 0.008144f
C453 VTAIL.n410 B 1.12075f
C454 VTAIL.n411 B 0.015155f
C455 VTAIL.n412 B 0.008144f
C456 VTAIL.n413 B 0.008623f
C457 VTAIL.n414 B 0.019249f
C458 VTAIL.n415 B 0.019249f
C459 VTAIL.n416 B 0.008623f
C460 VTAIL.n417 B 0.008144f
C461 VTAIL.n418 B 0.015155f
C462 VTAIL.n419 B 0.015155f
C463 VTAIL.n420 B 0.008144f
C464 VTAIL.n421 B 0.008623f
C465 VTAIL.n422 B 0.019249f
C466 VTAIL.n423 B 0.019249f
C467 VTAIL.n424 B 0.008623f
C468 VTAIL.n425 B 0.008144f
C469 VTAIL.n426 B 0.015155f
C470 VTAIL.n427 B 0.015155f
C471 VTAIL.n428 B 0.008144f
C472 VTAIL.n429 B 0.008623f
C473 VTAIL.n430 B 0.019249f
C474 VTAIL.n431 B 0.019249f
C475 VTAIL.n432 B 0.008623f
C476 VTAIL.n433 B 0.008144f
C477 VTAIL.n434 B 0.015155f
C478 VTAIL.n435 B 0.015155f
C479 VTAIL.n436 B 0.008144f
C480 VTAIL.n437 B 0.008623f
C481 VTAIL.n438 B 0.019249f
C482 VTAIL.n439 B 0.019249f
C483 VTAIL.n440 B 0.008623f
C484 VTAIL.n441 B 0.008144f
C485 VTAIL.n442 B 0.015155f
C486 VTAIL.n443 B 0.015155f
C487 VTAIL.n444 B 0.008144f
C488 VTAIL.n445 B 0.008623f
C489 VTAIL.n446 B 0.019249f
C490 VTAIL.n447 B 0.019249f
C491 VTAIL.n448 B 0.008623f
C492 VTAIL.n449 B 0.008144f
C493 VTAIL.n450 B 0.015155f
C494 VTAIL.n451 B 0.015155f
C495 VTAIL.n452 B 0.008144f
C496 VTAIL.n453 B 0.008383f
C497 VTAIL.n454 B 0.008383f
C498 VTAIL.n455 B 0.019249f
C499 VTAIL.n456 B 0.019249f
C500 VTAIL.n457 B 0.008623f
C501 VTAIL.n458 B 0.008144f
C502 VTAIL.n459 B 0.015155f
C503 VTAIL.n460 B 0.015155f
C504 VTAIL.n461 B 0.008144f
C505 VTAIL.n462 B 0.008623f
C506 VTAIL.n463 B 0.019249f
C507 VTAIL.n464 B 0.042755f
C508 VTAIL.n465 B 0.008623f
C509 VTAIL.n466 B 0.008144f
C510 VTAIL.n467 B 0.037928f
C511 VTAIL.n468 B 0.02412f
C512 VTAIL.n469 B 0.114142f
C513 VTAIL.n470 B 0.021915f
C514 VTAIL.n471 B 0.015155f
C515 VTAIL.n472 B 0.008144f
C516 VTAIL.n473 B 0.019249f
C517 VTAIL.n474 B 0.008623f
C518 VTAIL.n475 B 0.015155f
C519 VTAIL.n476 B 0.008144f
C520 VTAIL.n477 B 0.019249f
C521 VTAIL.n478 B 0.008623f
C522 VTAIL.n479 B 0.015155f
C523 VTAIL.n480 B 0.008144f
C524 VTAIL.n481 B 0.019249f
C525 VTAIL.n482 B 0.019249f
C526 VTAIL.n483 B 0.008623f
C527 VTAIL.n484 B 0.015155f
C528 VTAIL.n485 B 0.008144f
C529 VTAIL.n486 B 0.019249f
C530 VTAIL.n487 B 0.008623f
C531 VTAIL.n488 B 0.015155f
C532 VTAIL.n489 B 0.008144f
C533 VTAIL.n490 B 0.019249f
C534 VTAIL.n491 B 0.008623f
C535 VTAIL.n492 B 0.015155f
C536 VTAIL.n493 B 0.008144f
C537 VTAIL.n494 B 0.019249f
C538 VTAIL.n495 B 0.008623f
C539 VTAIL.n496 B 0.015155f
C540 VTAIL.n497 B 0.008144f
C541 VTAIL.n498 B 0.019249f
C542 VTAIL.n499 B 0.008623f
C543 VTAIL.n500 B 0.106215f
C544 VTAIL.t1 B 0.031839f
C545 VTAIL.n501 B 0.014436f
C546 VTAIL.n502 B 0.011371f
C547 VTAIL.n503 B 0.008144f
C548 VTAIL.n504 B 1.12075f
C549 VTAIL.n505 B 0.015155f
C550 VTAIL.n506 B 0.008144f
C551 VTAIL.n507 B 0.008623f
C552 VTAIL.n508 B 0.019249f
C553 VTAIL.n509 B 0.019249f
C554 VTAIL.n510 B 0.008623f
C555 VTAIL.n511 B 0.008144f
C556 VTAIL.n512 B 0.015155f
C557 VTAIL.n513 B 0.015155f
C558 VTAIL.n514 B 0.008144f
C559 VTAIL.n515 B 0.008623f
C560 VTAIL.n516 B 0.019249f
C561 VTAIL.n517 B 0.019249f
C562 VTAIL.n518 B 0.008623f
C563 VTAIL.n519 B 0.008144f
C564 VTAIL.n520 B 0.015155f
C565 VTAIL.n521 B 0.015155f
C566 VTAIL.n522 B 0.008144f
C567 VTAIL.n523 B 0.008623f
C568 VTAIL.n524 B 0.019249f
C569 VTAIL.n525 B 0.019249f
C570 VTAIL.n526 B 0.008623f
C571 VTAIL.n527 B 0.008144f
C572 VTAIL.n528 B 0.015155f
C573 VTAIL.n529 B 0.015155f
C574 VTAIL.n530 B 0.008144f
C575 VTAIL.n531 B 0.008623f
C576 VTAIL.n532 B 0.019249f
C577 VTAIL.n533 B 0.019249f
C578 VTAIL.n534 B 0.008623f
C579 VTAIL.n535 B 0.008144f
C580 VTAIL.n536 B 0.015155f
C581 VTAIL.n537 B 0.015155f
C582 VTAIL.n538 B 0.008144f
C583 VTAIL.n539 B 0.008623f
C584 VTAIL.n540 B 0.019249f
C585 VTAIL.n541 B 0.019249f
C586 VTAIL.n542 B 0.008623f
C587 VTAIL.n543 B 0.008144f
C588 VTAIL.n544 B 0.015155f
C589 VTAIL.n545 B 0.015155f
C590 VTAIL.n546 B 0.008144f
C591 VTAIL.n547 B 0.008383f
C592 VTAIL.n548 B 0.008383f
C593 VTAIL.n549 B 0.019249f
C594 VTAIL.n550 B 0.019249f
C595 VTAIL.n551 B 0.008623f
C596 VTAIL.n552 B 0.008144f
C597 VTAIL.n553 B 0.015155f
C598 VTAIL.n554 B 0.015155f
C599 VTAIL.n555 B 0.008144f
C600 VTAIL.n556 B 0.008623f
C601 VTAIL.n557 B 0.019249f
C602 VTAIL.n558 B 0.042755f
C603 VTAIL.n559 B 0.008623f
C604 VTAIL.n560 B 0.008144f
C605 VTAIL.n561 B 0.037928f
C606 VTAIL.n562 B 0.02412f
C607 VTAIL.n563 B 0.114142f
C608 VTAIL.n564 B 0.021915f
C609 VTAIL.n565 B 0.015155f
C610 VTAIL.n566 B 0.008144f
C611 VTAIL.n567 B 0.019249f
C612 VTAIL.n568 B 0.008623f
C613 VTAIL.n569 B 0.015155f
C614 VTAIL.n570 B 0.008144f
C615 VTAIL.n571 B 0.019249f
C616 VTAIL.n572 B 0.008623f
C617 VTAIL.n573 B 0.015155f
C618 VTAIL.n574 B 0.008144f
C619 VTAIL.n575 B 0.019249f
C620 VTAIL.n576 B 0.019249f
C621 VTAIL.n577 B 0.008623f
C622 VTAIL.n578 B 0.015155f
C623 VTAIL.n579 B 0.008144f
C624 VTAIL.n580 B 0.019249f
C625 VTAIL.n581 B 0.008623f
C626 VTAIL.n582 B 0.015155f
C627 VTAIL.n583 B 0.008144f
C628 VTAIL.n584 B 0.019249f
C629 VTAIL.n585 B 0.008623f
C630 VTAIL.n586 B 0.015155f
C631 VTAIL.n587 B 0.008144f
C632 VTAIL.n588 B 0.019249f
C633 VTAIL.n589 B 0.008623f
C634 VTAIL.n590 B 0.015155f
C635 VTAIL.n591 B 0.008144f
C636 VTAIL.n592 B 0.019249f
C637 VTAIL.n593 B 0.008623f
C638 VTAIL.n594 B 0.106215f
C639 VTAIL.t3 B 0.031839f
C640 VTAIL.n595 B 0.014436f
C641 VTAIL.n596 B 0.011371f
C642 VTAIL.n597 B 0.008144f
C643 VTAIL.n598 B 1.12075f
C644 VTAIL.n599 B 0.015155f
C645 VTAIL.n600 B 0.008144f
C646 VTAIL.n601 B 0.008623f
C647 VTAIL.n602 B 0.019249f
C648 VTAIL.n603 B 0.019249f
C649 VTAIL.n604 B 0.008623f
C650 VTAIL.n605 B 0.008144f
C651 VTAIL.n606 B 0.015155f
C652 VTAIL.n607 B 0.015155f
C653 VTAIL.n608 B 0.008144f
C654 VTAIL.n609 B 0.008623f
C655 VTAIL.n610 B 0.019249f
C656 VTAIL.n611 B 0.019249f
C657 VTAIL.n612 B 0.008623f
C658 VTAIL.n613 B 0.008144f
C659 VTAIL.n614 B 0.015155f
C660 VTAIL.n615 B 0.015155f
C661 VTAIL.n616 B 0.008144f
C662 VTAIL.n617 B 0.008623f
C663 VTAIL.n618 B 0.019249f
C664 VTAIL.n619 B 0.019249f
C665 VTAIL.n620 B 0.008623f
C666 VTAIL.n621 B 0.008144f
C667 VTAIL.n622 B 0.015155f
C668 VTAIL.n623 B 0.015155f
C669 VTAIL.n624 B 0.008144f
C670 VTAIL.n625 B 0.008623f
C671 VTAIL.n626 B 0.019249f
C672 VTAIL.n627 B 0.019249f
C673 VTAIL.n628 B 0.008623f
C674 VTAIL.n629 B 0.008144f
C675 VTAIL.n630 B 0.015155f
C676 VTAIL.n631 B 0.015155f
C677 VTAIL.n632 B 0.008144f
C678 VTAIL.n633 B 0.008623f
C679 VTAIL.n634 B 0.019249f
C680 VTAIL.n635 B 0.019249f
C681 VTAIL.n636 B 0.008623f
C682 VTAIL.n637 B 0.008144f
C683 VTAIL.n638 B 0.015155f
C684 VTAIL.n639 B 0.015155f
C685 VTAIL.n640 B 0.008144f
C686 VTAIL.n641 B 0.008383f
C687 VTAIL.n642 B 0.008383f
C688 VTAIL.n643 B 0.019249f
C689 VTAIL.n644 B 0.019249f
C690 VTAIL.n645 B 0.008623f
C691 VTAIL.n646 B 0.008144f
C692 VTAIL.n647 B 0.015155f
C693 VTAIL.n648 B 0.015155f
C694 VTAIL.n649 B 0.008144f
C695 VTAIL.n650 B 0.008623f
C696 VTAIL.n651 B 0.019249f
C697 VTAIL.n652 B 0.042755f
C698 VTAIL.n653 B 0.008623f
C699 VTAIL.n654 B 0.008144f
C700 VTAIL.n655 B 0.037928f
C701 VTAIL.n656 B 0.02412f
C702 VTAIL.n657 B 1.0868f
C703 VTAIL.n658 B 0.021915f
C704 VTAIL.n659 B 0.015155f
C705 VTAIL.n660 B 0.008144f
C706 VTAIL.n661 B 0.019249f
C707 VTAIL.n662 B 0.008623f
C708 VTAIL.n663 B 0.015155f
C709 VTAIL.n664 B 0.008144f
C710 VTAIL.n665 B 0.019249f
C711 VTAIL.n666 B 0.008623f
C712 VTAIL.n667 B 0.015155f
C713 VTAIL.n668 B 0.008144f
C714 VTAIL.n669 B 0.019249f
C715 VTAIL.n670 B 0.008623f
C716 VTAIL.n671 B 0.015155f
C717 VTAIL.n672 B 0.008144f
C718 VTAIL.n673 B 0.019249f
C719 VTAIL.n674 B 0.008623f
C720 VTAIL.n675 B 0.015155f
C721 VTAIL.n676 B 0.008144f
C722 VTAIL.n677 B 0.019249f
C723 VTAIL.n678 B 0.008623f
C724 VTAIL.n679 B 0.015155f
C725 VTAIL.n680 B 0.008144f
C726 VTAIL.n681 B 0.019249f
C727 VTAIL.n682 B 0.008623f
C728 VTAIL.n683 B 0.015155f
C729 VTAIL.n684 B 0.008144f
C730 VTAIL.n685 B 0.019249f
C731 VTAIL.n686 B 0.008623f
C732 VTAIL.n687 B 0.106215f
C733 VTAIL.t5 B 0.031839f
C734 VTAIL.n688 B 0.014436f
C735 VTAIL.n689 B 0.011371f
C736 VTAIL.n690 B 0.008144f
C737 VTAIL.n691 B 1.12075f
C738 VTAIL.n692 B 0.015155f
C739 VTAIL.n693 B 0.008144f
C740 VTAIL.n694 B 0.008623f
C741 VTAIL.n695 B 0.019249f
C742 VTAIL.n696 B 0.019249f
C743 VTAIL.n697 B 0.008623f
C744 VTAIL.n698 B 0.008144f
C745 VTAIL.n699 B 0.015155f
C746 VTAIL.n700 B 0.015155f
C747 VTAIL.n701 B 0.008144f
C748 VTAIL.n702 B 0.008623f
C749 VTAIL.n703 B 0.019249f
C750 VTAIL.n704 B 0.019249f
C751 VTAIL.n705 B 0.008623f
C752 VTAIL.n706 B 0.008144f
C753 VTAIL.n707 B 0.015155f
C754 VTAIL.n708 B 0.015155f
C755 VTAIL.n709 B 0.008144f
C756 VTAIL.n710 B 0.008623f
C757 VTAIL.n711 B 0.019249f
C758 VTAIL.n712 B 0.019249f
C759 VTAIL.n713 B 0.008623f
C760 VTAIL.n714 B 0.008144f
C761 VTAIL.n715 B 0.015155f
C762 VTAIL.n716 B 0.015155f
C763 VTAIL.n717 B 0.008144f
C764 VTAIL.n718 B 0.008623f
C765 VTAIL.n719 B 0.019249f
C766 VTAIL.n720 B 0.019249f
C767 VTAIL.n721 B 0.008623f
C768 VTAIL.n722 B 0.008144f
C769 VTAIL.n723 B 0.015155f
C770 VTAIL.n724 B 0.015155f
C771 VTAIL.n725 B 0.008144f
C772 VTAIL.n726 B 0.008623f
C773 VTAIL.n727 B 0.019249f
C774 VTAIL.n728 B 0.019249f
C775 VTAIL.n729 B 0.019249f
C776 VTAIL.n730 B 0.008623f
C777 VTAIL.n731 B 0.008144f
C778 VTAIL.n732 B 0.015155f
C779 VTAIL.n733 B 0.015155f
C780 VTAIL.n734 B 0.008144f
C781 VTAIL.n735 B 0.008383f
C782 VTAIL.n736 B 0.008383f
C783 VTAIL.n737 B 0.019249f
C784 VTAIL.n738 B 0.019249f
C785 VTAIL.n739 B 0.008623f
C786 VTAIL.n740 B 0.008144f
C787 VTAIL.n741 B 0.015155f
C788 VTAIL.n742 B 0.015155f
C789 VTAIL.n743 B 0.008144f
C790 VTAIL.n744 B 0.008623f
C791 VTAIL.n745 B 0.019249f
C792 VTAIL.n746 B 0.042755f
C793 VTAIL.n747 B 0.008623f
C794 VTAIL.n748 B 0.008144f
C795 VTAIL.n749 B 0.037928f
C796 VTAIL.n750 B 0.02412f
C797 VTAIL.n751 B 1.04565f
C798 VDD2.t3 B 0.35795f
C799 VDD2.t1 B 0.35795f
C800 VDD2.n0 B 4.03279f
C801 VDD2.t2 B 0.35795f
C802 VDD2.t0 B 0.35795f
C803 VDD2.n1 B 3.25605f
C804 VDD2.n2 B 4.03842f
C805 VN.t1 B 2.50409f
C806 VN.t2 B 2.50307f
C807 VN.n0 B 1.78657f
C808 VN.t3 B 2.50409f
C809 VN.t0 B 2.50307f
C810 VN.n1 B 3.26587f
.ends

