* NGSPICE file created from diff_pair_sample_0494.ext - technology: sky130A

.subckt diff_pair_sample_0494 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t10 VN.t0 VDD2.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=2.77695 pd=17.16 as=2.77695 ps=17.16 w=16.83 l=0.87
X1 B.t19 B.t17 B.t18 B.t11 sky130_fd_pr__nfet_01v8 ad=6.5637 pd=34.44 as=0 ps=0 w=16.83 l=0.87
X2 VDD2.t4 VN.t1 VTAIL.t9 B.t1 sky130_fd_pr__nfet_01v8 ad=6.5637 pd=34.44 as=2.77695 ps=17.16 w=16.83 l=0.87
X3 VDD1.t5 VP.t0 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=2.77695 pd=17.16 as=6.5637 ps=34.44 w=16.83 l=0.87
X4 VTAIL.t3 VP.t1 VDD1.t4 B.t3 sky130_fd_pr__nfet_01v8 ad=2.77695 pd=17.16 as=2.77695 ps=17.16 w=16.83 l=0.87
X5 B.t16 B.t14 B.t15 B.t7 sky130_fd_pr__nfet_01v8 ad=6.5637 pd=34.44 as=0 ps=0 w=16.83 l=0.87
X6 VDD1.t3 VP.t2 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=6.5637 pd=34.44 as=2.77695 ps=17.16 w=16.83 l=0.87
X7 VDD1.t2 VP.t3 VTAIL.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=2.77695 pd=17.16 as=6.5637 ps=34.44 w=16.83 l=0.87
X8 VDD1.t1 VP.t4 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=6.5637 pd=34.44 as=2.77695 ps=17.16 w=16.83 l=0.87
X9 VDD2.t5 VN.t2 VTAIL.t8 B.t4 sky130_fd_pr__nfet_01v8 ad=2.77695 pd=17.16 as=6.5637 ps=34.44 w=16.83 l=0.87
X10 VDD2.t2 VN.t3 VTAIL.t7 B.t2 sky130_fd_pr__nfet_01v8 ad=6.5637 pd=34.44 as=2.77695 ps=17.16 w=16.83 l=0.87
X11 B.t13 B.t10 B.t12 B.t11 sky130_fd_pr__nfet_01v8 ad=6.5637 pd=34.44 as=0 ps=0 w=16.83 l=0.87
X12 VDD2.t0 VN.t4 VTAIL.t6 B.t0 sky130_fd_pr__nfet_01v8 ad=2.77695 pd=17.16 as=6.5637 ps=34.44 w=16.83 l=0.87
X13 VTAIL.t11 VP.t5 VDD1.t0 B.t5 sky130_fd_pr__nfet_01v8 ad=2.77695 pd=17.16 as=2.77695 ps=17.16 w=16.83 l=0.87
X14 B.t9 B.t6 B.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=6.5637 pd=34.44 as=0 ps=0 w=16.83 l=0.87
X15 VTAIL.t5 VN.t5 VDD2.t1 B.t5 sky130_fd_pr__nfet_01v8 ad=2.77695 pd=17.16 as=2.77695 ps=17.16 w=16.83 l=0.87
R0 VN.n2 VN.t1 527.88
R1 VN.n10 VN.t2 527.88
R2 VN.n6 VN.t4 511.64
R3 VN.n14 VN.t3 511.64
R4 VN.n1 VN.t5 466.211
R5 VN.n9 VN.t0 466.211
R6 VN.n7 VN.n6 161.3
R7 VN.n15 VN.n14 161.3
R8 VN.n13 VN.n8 161.3
R9 VN.n12 VN.n11 161.3
R10 VN.n5 VN.n0 161.3
R11 VN.n4 VN.n3 161.3
R12 VN.n5 VN.n4 55.0624
R13 VN.n13 VN.n12 55.0624
R14 VN VN.n15 45.8888
R15 VN.n11 VN.n10 43.7084
R16 VN.n3 VN.n2 43.7084
R17 VN.n2 VN.n1 42.6481
R18 VN.n10 VN.n9 42.6481
R19 VN.n4 VN.n1 12.234
R20 VN.n12 VN.n9 12.234
R21 VN.n6 VN.n5 2.19141
R22 VN.n14 VN.n13 2.19141
R23 VN.n15 VN.n8 0.189894
R24 VN.n11 VN.n8 0.189894
R25 VN.n3 VN.n0 0.189894
R26 VN.n7 VN.n0 0.189894
R27 VN VN.n7 0.0516364
R28 VDD2.n183 VDD2.n95 289.615
R29 VDD2.n88 VDD2.n0 289.615
R30 VDD2.n184 VDD2.n183 185
R31 VDD2.n182 VDD2.n181 185
R32 VDD2.n99 VDD2.n98 185
R33 VDD2.n176 VDD2.n175 185
R34 VDD2.n174 VDD2.n173 185
R35 VDD2.n172 VDD2.n102 185
R36 VDD2.n106 VDD2.n103 185
R37 VDD2.n167 VDD2.n166 185
R38 VDD2.n165 VDD2.n164 185
R39 VDD2.n108 VDD2.n107 185
R40 VDD2.n159 VDD2.n158 185
R41 VDD2.n157 VDD2.n156 185
R42 VDD2.n112 VDD2.n111 185
R43 VDD2.n151 VDD2.n150 185
R44 VDD2.n149 VDD2.n148 185
R45 VDD2.n116 VDD2.n115 185
R46 VDD2.n143 VDD2.n142 185
R47 VDD2.n141 VDD2.n140 185
R48 VDD2.n120 VDD2.n119 185
R49 VDD2.n135 VDD2.n134 185
R50 VDD2.n133 VDD2.n132 185
R51 VDD2.n124 VDD2.n123 185
R52 VDD2.n127 VDD2.n126 185
R53 VDD2.n31 VDD2.n30 185
R54 VDD2.n28 VDD2.n27 185
R55 VDD2.n37 VDD2.n36 185
R56 VDD2.n39 VDD2.n38 185
R57 VDD2.n24 VDD2.n23 185
R58 VDD2.n45 VDD2.n44 185
R59 VDD2.n47 VDD2.n46 185
R60 VDD2.n20 VDD2.n19 185
R61 VDD2.n53 VDD2.n52 185
R62 VDD2.n55 VDD2.n54 185
R63 VDD2.n16 VDD2.n15 185
R64 VDD2.n61 VDD2.n60 185
R65 VDD2.n63 VDD2.n62 185
R66 VDD2.n12 VDD2.n11 185
R67 VDD2.n69 VDD2.n68 185
R68 VDD2.n72 VDD2.n71 185
R69 VDD2.n70 VDD2.n8 185
R70 VDD2.n77 VDD2.n7 185
R71 VDD2.n79 VDD2.n78 185
R72 VDD2.n81 VDD2.n80 185
R73 VDD2.n4 VDD2.n3 185
R74 VDD2.n87 VDD2.n86 185
R75 VDD2.n89 VDD2.n88 185
R76 VDD2.t2 VDD2.n125 147.659
R77 VDD2.t4 VDD2.n29 147.659
R78 VDD2.n183 VDD2.n182 104.615
R79 VDD2.n182 VDD2.n98 104.615
R80 VDD2.n175 VDD2.n98 104.615
R81 VDD2.n175 VDD2.n174 104.615
R82 VDD2.n174 VDD2.n102 104.615
R83 VDD2.n106 VDD2.n102 104.615
R84 VDD2.n166 VDD2.n106 104.615
R85 VDD2.n166 VDD2.n165 104.615
R86 VDD2.n165 VDD2.n107 104.615
R87 VDD2.n158 VDD2.n107 104.615
R88 VDD2.n158 VDD2.n157 104.615
R89 VDD2.n157 VDD2.n111 104.615
R90 VDD2.n150 VDD2.n111 104.615
R91 VDD2.n150 VDD2.n149 104.615
R92 VDD2.n149 VDD2.n115 104.615
R93 VDD2.n142 VDD2.n115 104.615
R94 VDD2.n142 VDD2.n141 104.615
R95 VDD2.n141 VDD2.n119 104.615
R96 VDD2.n134 VDD2.n119 104.615
R97 VDD2.n134 VDD2.n133 104.615
R98 VDD2.n133 VDD2.n123 104.615
R99 VDD2.n126 VDD2.n123 104.615
R100 VDD2.n30 VDD2.n27 104.615
R101 VDD2.n37 VDD2.n27 104.615
R102 VDD2.n38 VDD2.n37 104.615
R103 VDD2.n38 VDD2.n23 104.615
R104 VDD2.n45 VDD2.n23 104.615
R105 VDD2.n46 VDD2.n45 104.615
R106 VDD2.n46 VDD2.n19 104.615
R107 VDD2.n53 VDD2.n19 104.615
R108 VDD2.n54 VDD2.n53 104.615
R109 VDD2.n54 VDD2.n15 104.615
R110 VDD2.n61 VDD2.n15 104.615
R111 VDD2.n62 VDD2.n61 104.615
R112 VDD2.n62 VDD2.n11 104.615
R113 VDD2.n69 VDD2.n11 104.615
R114 VDD2.n71 VDD2.n69 104.615
R115 VDD2.n71 VDD2.n70 104.615
R116 VDD2.n70 VDD2.n7 104.615
R117 VDD2.n79 VDD2.n7 104.615
R118 VDD2.n80 VDD2.n79 104.615
R119 VDD2.n80 VDD2.n3 104.615
R120 VDD2.n87 VDD2.n3 104.615
R121 VDD2.n88 VDD2.n87 104.615
R122 VDD2.n94 VDD2.n93 61.5097
R123 VDD2 VDD2.n189 61.5069
R124 VDD2.n126 VDD2.t2 52.3082
R125 VDD2.n30 VDD2.t4 52.3082
R126 VDD2.n94 VDD2.n92 50.1665
R127 VDD2.n188 VDD2.n187 49.446
R128 VDD2.n188 VDD2.n94 41.586
R129 VDD2.n127 VDD2.n125 15.6677
R130 VDD2.n31 VDD2.n29 15.6677
R131 VDD2.n173 VDD2.n172 13.1884
R132 VDD2.n78 VDD2.n77 13.1884
R133 VDD2.n176 VDD2.n101 12.8005
R134 VDD2.n171 VDD2.n103 12.8005
R135 VDD2.n128 VDD2.n124 12.8005
R136 VDD2.n32 VDD2.n28 12.8005
R137 VDD2.n76 VDD2.n8 12.8005
R138 VDD2.n81 VDD2.n6 12.8005
R139 VDD2.n177 VDD2.n99 12.0247
R140 VDD2.n168 VDD2.n167 12.0247
R141 VDD2.n132 VDD2.n131 12.0247
R142 VDD2.n36 VDD2.n35 12.0247
R143 VDD2.n73 VDD2.n72 12.0247
R144 VDD2.n82 VDD2.n4 12.0247
R145 VDD2.n181 VDD2.n180 11.249
R146 VDD2.n164 VDD2.n105 11.249
R147 VDD2.n135 VDD2.n122 11.249
R148 VDD2.n39 VDD2.n26 11.249
R149 VDD2.n68 VDD2.n10 11.249
R150 VDD2.n86 VDD2.n85 11.249
R151 VDD2.n184 VDD2.n97 10.4732
R152 VDD2.n163 VDD2.n108 10.4732
R153 VDD2.n136 VDD2.n120 10.4732
R154 VDD2.n40 VDD2.n24 10.4732
R155 VDD2.n67 VDD2.n12 10.4732
R156 VDD2.n89 VDD2.n2 10.4732
R157 VDD2.n185 VDD2.n95 9.69747
R158 VDD2.n160 VDD2.n159 9.69747
R159 VDD2.n140 VDD2.n139 9.69747
R160 VDD2.n44 VDD2.n43 9.69747
R161 VDD2.n64 VDD2.n63 9.69747
R162 VDD2.n90 VDD2.n0 9.69747
R163 VDD2.n187 VDD2.n186 9.45567
R164 VDD2.n92 VDD2.n91 9.45567
R165 VDD2.n153 VDD2.n152 9.3005
R166 VDD2.n155 VDD2.n154 9.3005
R167 VDD2.n110 VDD2.n109 9.3005
R168 VDD2.n161 VDD2.n160 9.3005
R169 VDD2.n163 VDD2.n162 9.3005
R170 VDD2.n105 VDD2.n104 9.3005
R171 VDD2.n169 VDD2.n168 9.3005
R172 VDD2.n171 VDD2.n170 9.3005
R173 VDD2.n186 VDD2.n185 9.3005
R174 VDD2.n97 VDD2.n96 9.3005
R175 VDD2.n180 VDD2.n179 9.3005
R176 VDD2.n178 VDD2.n177 9.3005
R177 VDD2.n101 VDD2.n100 9.3005
R178 VDD2.n114 VDD2.n113 9.3005
R179 VDD2.n147 VDD2.n146 9.3005
R180 VDD2.n145 VDD2.n144 9.3005
R181 VDD2.n118 VDD2.n117 9.3005
R182 VDD2.n139 VDD2.n138 9.3005
R183 VDD2.n137 VDD2.n136 9.3005
R184 VDD2.n122 VDD2.n121 9.3005
R185 VDD2.n131 VDD2.n130 9.3005
R186 VDD2.n129 VDD2.n128 9.3005
R187 VDD2.n91 VDD2.n90 9.3005
R188 VDD2.n2 VDD2.n1 9.3005
R189 VDD2.n85 VDD2.n84 9.3005
R190 VDD2.n83 VDD2.n82 9.3005
R191 VDD2.n6 VDD2.n5 9.3005
R192 VDD2.n51 VDD2.n50 9.3005
R193 VDD2.n49 VDD2.n48 9.3005
R194 VDD2.n22 VDD2.n21 9.3005
R195 VDD2.n43 VDD2.n42 9.3005
R196 VDD2.n41 VDD2.n40 9.3005
R197 VDD2.n26 VDD2.n25 9.3005
R198 VDD2.n35 VDD2.n34 9.3005
R199 VDD2.n33 VDD2.n32 9.3005
R200 VDD2.n18 VDD2.n17 9.3005
R201 VDD2.n57 VDD2.n56 9.3005
R202 VDD2.n59 VDD2.n58 9.3005
R203 VDD2.n14 VDD2.n13 9.3005
R204 VDD2.n65 VDD2.n64 9.3005
R205 VDD2.n67 VDD2.n66 9.3005
R206 VDD2.n10 VDD2.n9 9.3005
R207 VDD2.n74 VDD2.n73 9.3005
R208 VDD2.n76 VDD2.n75 9.3005
R209 VDD2.n156 VDD2.n110 8.92171
R210 VDD2.n143 VDD2.n118 8.92171
R211 VDD2.n47 VDD2.n22 8.92171
R212 VDD2.n60 VDD2.n14 8.92171
R213 VDD2.n155 VDD2.n112 8.14595
R214 VDD2.n144 VDD2.n116 8.14595
R215 VDD2.n48 VDD2.n20 8.14595
R216 VDD2.n59 VDD2.n16 8.14595
R217 VDD2.n152 VDD2.n151 7.3702
R218 VDD2.n148 VDD2.n147 7.3702
R219 VDD2.n52 VDD2.n51 7.3702
R220 VDD2.n56 VDD2.n55 7.3702
R221 VDD2.n151 VDD2.n114 6.59444
R222 VDD2.n148 VDD2.n114 6.59444
R223 VDD2.n52 VDD2.n18 6.59444
R224 VDD2.n55 VDD2.n18 6.59444
R225 VDD2.n152 VDD2.n112 5.81868
R226 VDD2.n147 VDD2.n116 5.81868
R227 VDD2.n51 VDD2.n20 5.81868
R228 VDD2.n56 VDD2.n16 5.81868
R229 VDD2.n156 VDD2.n155 5.04292
R230 VDD2.n144 VDD2.n143 5.04292
R231 VDD2.n48 VDD2.n47 5.04292
R232 VDD2.n60 VDD2.n59 5.04292
R233 VDD2.n129 VDD2.n125 4.38563
R234 VDD2.n33 VDD2.n29 4.38563
R235 VDD2.n187 VDD2.n95 4.26717
R236 VDD2.n159 VDD2.n110 4.26717
R237 VDD2.n140 VDD2.n118 4.26717
R238 VDD2.n44 VDD2.n22 4.26717
R239 VDD2.n63 VDD2.n14 4.26717
R240 VDD2.n92 VDD2.n0 4.26717
R241 VDD2.n185 VDD2.n184 3.49141
R242 VDD2.n160 VDD2.n108 3.49141
R243 VDD2.n139 VDD2.n120 3.49141
R244 VDD2.n43 VDD2.n24 3.49141
R245 VDD2.n64 VDD2.n12 3.49141
R246 VDD2.n90 VDD2.n89 3.49141
R247 VDD2.n181 VDD2.n97 2.71565
R248 VDD2.n164 VDD2.n163 2.71565
R249 VDD2.n136 VDD2.n135 2.71565
R250 VDD2.n40 VDD2.n39 2.71565
R251 VDD2.n68 VDD2.n67 2.71565
R252 VDD2.n86 VDD2.n2 2.71565
R253 VDD2.n180 VDD2.n99 1.93989
R254 VDD2.n167 VDD2.n105 1.93989
R255 VDD2.n132 VDD2.n122 1.93989
R256 VDD2.n36 VDD2.n26 1.93989
R257 VDD2.n72 VDD2.n10 1.93989
R258 VDD2.n85 VDD2.n4 1.93989
R259 VDD2.n189 VDD2.t3 1.17697
R260 VDD2.n189 VDD2.t5 1.17697
R261 VDD2.n93 VDD2.t1 1.17697
R262 VDD2.n93 VDD2.t0 1.17697
R263 VDD2.n177 VDD2.n176 1.16414
R264 VDD2.n168 VDD2.n103 1.16414
R265 VDD2.n131 VDD2.n124 1.16414
R266 VDD2.n35 VDD2.n28 1.16414
R267 VDD2.n73 VDD2.n8 1.16414
R268 VDD2.n82 VDD2.n81 1.16414
R269 VDD2 VDD2.n188 0.834552
R270 VDD2.n173 VDD2.n101 0.388379
R271 VDD2.n172 VDD2.n171 0.388379
R272 VDD2.n128 VDD2.n127 0.388379
R273 VDD2.n32 VDD2.n31 0.388379
R274 VDD2.n77 VDD2.n76 0.388379
R275 VDD2.n78 VDD2.n6 0.388379
R276 VDD2.n186 VDD2.n96 0.155672
R277 VDD2.n179 VDD2.n96 0.155672
R278 VDD2.n179 VDD2.n178 0.155672
R279 VDD2.n178 VDD2.n100 0.155672
R280 VDD2.n170 VDD2.n100 0.155672
R281 VDD2.n170 VDD2.n169 0.155672
R282 VDD2.n169 VDD2.n104 0.155672
R283 VDD2.n162 VDD2.n104 0.155672
R284 VDD2.n162 VDD2.n161 0.155672
R285 VDD2.n161 VDD2.n109 0.155672
R286 VDD2.n154 VDD2.n109 0.155672
R287 VDD2.n154 VDD2.n153 0.155672
R288 VDD2.n153 VDD2.n113 0.155672
R289 VDD2.n146 VDD2.n113 0.155672
R290 VDD2.n146 VDD2.n145 0.155672
R291 VDD2.n145 VDD2.n117 0.155672
R292 VDD2.n138 VDD2.n117 0.155672
R293 VDD2.n138 VDD2.n137 0.155672
R294 VDD2.n137 VDD2.n121 0.155672
R295 VDD2.n130 VDD2.n121 0.155672
R296 VDD2.n130 VDD2.n129 0.155672
R297 VDD2.n34 VDD2.n33 0.155672
R298 VDD2.n34 VDD2.n25 0.155672
R299 VDD2.n41 VDD2.n25 0.155672
R300 VDD2.n42 VDD2.n41 0.155672
R301 VDD2.n42 VDD2.n21 0.155672
R302 VDD2.n49 VDD2.n21 0.155672
R303 VDD2.n50 VDD2.n49 0.155672
R304 VDD2.n50 VDD2.n17 0.155672
R305 VDD2.n57 VDD2.n17 0.155672
R306 VDD2.n58 VDD2.n57 0.155672
R307 VDD2.n58 VDD2.n13 0.155672
R308 VDD2.n65 VDD2.n13 0.155672
R309 VDD2.n66 VDD2.n65 0.155672
R310 VDD2.n66 VDD2.n9 0.155672
R311 VDD2.n74 VDD2.n9 0.155672
R312 VDD2.n75 VDD2.n74 0.155672
R313 VDD2.n75 VDD2.n5 0.155672
R314 VDD2.n83 VDD2.n5 0.155672
R315 VDD2.n84 VDD2.n83 0.155672
R316 VDD2.n84 VDD2.n1 0.155672
R317 VDD2.n91 VDD2.n1 0.155672
R318 VTAIL.n378 VTAIL.n290 289.615
R319 VTAIL.n90 VTAIL.n2 289.615
R320 VTAIL.n284 VTAIL.n196 289.615
R321 VTAIL.n188 VTAIL.n100 289.615
R322 VTAIL.n321 VTAIL.n320 185
R323 VTAIL.n318 VTAIL.n317 185
R324 VTAIL.n327 VTAIL.n326 185
R325 VTAIL.n329 VTAIL.n328 185
R326 VTAIL.n314 VTAIL.n313 185
R327 VTAIL.n335 VTAIL.n334 185
R328 VTAIL.n337 VTAIL.n336 185
R329 VTAIL.n310 VTAIL.n309 185
R330 VTAIL.n343 VTAIL.n342 185
R331 VTAIL.n345 VTAIL.n344 185
R332 VTAIL.n306 VTAIL.n305 185
R333 VTAIL.n351 VTAIL.n350 185
R334 VTAIL.n353 VTAIL.n352 185
R335 VTAIL.n302 VTAIL.n301 185
R336 VTAIL.n359 VTAIL.n358 185
R337 VTAIL.n362 VTAIL.n361 185
R338 VTAIL.n360 VTAIL.n298 185
R339 VTAIL.n367 VTAIL.n297 185
R340 VTAIL.n369 VTAIL.n368 185
R341 VTAIL.n371 VTAIL.n370 185
R342 VTAIL.n294 VTAIL.n293 185
R343 VTAIL.n377 VTAIL.n376 185
R344 VTAIL.n379 VTAIL.n378 185
R345 VTAIL.n33 VTAIL.n32 185
R346 VTAIL.n30 VTAIL.n29 185
R347 VTAIL.n39 VTAIL.n38 185
R348 VTAIL.n41 VTAIL.n40 185
R349 VTAIL.n26 VTAIL.n25 185
R350 VTAIL.n47 VTAIL.n46 185
R351 VTAIL.n49 VTAIL.n48 185
R352 VTAIL.n22 VTAIL.n21 185
R353 VTAIL.n55 VTAIL.n54 185
R354 VTAIL.n57 VTAIL.n56 185
R355 VTAIL.n18 VTAIL.n17 185
R356 VTAIL.n63 VTAIL.n62 185
R357 VTAIL.n65 VTAIL.n64 185
R358 VTAIL.n14 VTAIL.n13 185
R359 VTAIL.n71 VTAIL.n70 185
R360 VTAIL.n74 VTAIL.n73 185
R361 VTAIL.n72 VTAIL.n10 185
R362 VTAIL.n79 VTAIL.n9 185
R363 VTAIL.n81 VTAIL.n80 185
R364 VTAIL.n83 VTAIL.n82 185
R365 VTAIL.n6 VTAIL.n5 185
R366 VTAIL.n89 VTAIL.n88 185
R367 VTAIL.n91 VTAIL.n90 185
R368 VTAIL.n285 VTAIL.n284 185
R369 VTAIL.n283 VTAIL.n282 185
R370 VTAIL.n200 VTAIL.n199 185
R371 VTAIL.n277 VTAIL.n276 185
R372 VTAIL.n275 VTAIL.n274 185
R373 VTAIL.n273 VTAIL.n203 185
R374 VTAIL.n207 VTAIL.n204 185
R375 VTAIL.n268 VTAIL.n267 185
R376 VTAIL.n266 VTAIL.n265 185
R377 VTAIL.n209 VTAIL.n208 185
R378 VTAIL.n260 VTAIL.n259 185
R379 VTAIL.n258 VTAIL.n257 185
R380 VTAIL.n213 VTAIL.n212 185
R381 VTAIL.n252 VTAIL.n251 185
R382 VTAIL.n250 VTAIL.n249 185
R383 VTAIL.n217 VTAIL.n216 185
R384 VTAIL.n244 VTAIL.n243 185
R385 VTAIL.n242 VTAIL.n241 185
R386 VTAIL.n221 VTAIL.n220 185
R387 VTAIL.n236 VTAIL.n235 185
R388 VTAIL.n234 VTAIL.n233 185
R389 VTAIL.n225 VTAIL.n224 185
R390 VTAIL.n228 VTAIL.n227 185
R391 VTAIL.n189 VTAIL.n188 185
R392 VTAIL.n187 VTAIL.n186 185
R393 VTAIL.n104 VTAIL.n103 185
R394 VTAIL.n181 VTAIL.n180 185
R395 VTAIL.n179 VTAIL.n178 185
R396 VTAIL.n177 VTAIL.n107 185
R397 VTAIL.n111 VTAIL.n108 185
R398 VTAIL.n172 VTAIL.n171 185
R399 VTAIL.n170 VTAIL.n169 185
R400 VTAIL.n113 VTAIL.n112 185
R401 VTAIL.n164 VTAIL.n163 185
R402 VTAIL.n162 VTAIL.n161 185
R403 VTAIL.n117 VTAIL.n116 185
R404 VTAIL.n156 VTAIL.n155 185
R405 VTAIL.n154 VTAIL.n153 185
R406 VTAIL.n121 VTAIL.n120 185
R407 VTAIL.n148 VTAIL.n147 185
R408 VTAIL.n146 VTAIL.n145 185
R409 VTAIL.n125 VTAIL.n124 185
R410 VTAIL.n140 VTAIL.n139 185
R411 VTAIL.n138 VTAIL.n137 185
R412 VTAIL.n129 VTAIL.n128 185
R413 VTAIL.n132 VTAIL.n131 185
R414 VTAIL.t0 VTAIL.n226 147.659
R415 VTAIL.t8 VTAIL.n130 147.659
R416 VTAIL.t6 VTAIL.n319 147.659
R417 VTAIL.t4 VTAIL.n31 147.659
R418 VTAIL.n320 VTAIL.n317 104.615
R419 VTAIL.n327 VTAIL.n317 104.615
R420 VTAIL.n328 VTAIL.n327 104.615
R421 VTAIL.n328 VTAIL.n313 104.615
R422 VTAIL.n335 VTAIL.n313 104.615
R423 VTAIL.n336 VTAIL.n335 104.615
R424 VTAIL.n336 VTAIL.n309 104.615
R425 VTAIL.n343 VTAIL.n309 104.615
R426 VTAIL.n344 VTAIL.n343 104.615
R427 VTAIL.n344 VTAIL.n305 104.615
R428 VTAIL.n351 VTAIL.n305 104.615
R429 VTAIL.n352 VTAIL.n351 104.615
R430 VTAIL.n352 VTAIL.n301 104.615
R431 VTAIL.n359 VTAIL.n301 104.615
R432 VTAIL.n361 VTAIL.n359 104.615
R433 VTAIL.n361 VTAIL.n360 104.615
R434 VTAIL.n360 VTAIL.n297 104.615
R435 VTAIL.n369 VTAIL.n297 104.615
R436 VTAIL.n370 VTAIL.n369 104.615
R437 VTAIL.n370 VTAIL.n293 104.615
R438 VTAIL.n377 VTAIL.n293 104.615
R439 VTAIL.n378 VTAIL.n377 104.615
R440 VTAIL.n32 VTAIL.n29 104.615
R441 VTAIL.n39 VTAIL.n29 104.615
R442 VTAIL.n40 VTAIL.n39 104.615
R443 VTAIL.n40 VTAIL.n25 104.615
R444 VTAIL.n47 VTAIL.n25 104.615
R445 VTAIL.n48 VTAIL.n47 104.615
R446 VTAIL.n48 VTAIL.n21 104.615
R447 VTAIL.n55 VTAIL.n21 104.615
R448 VTAIL.n56 VTAIL.n55 104.615
R449 VTAIL.n56 VTAIL.n17 104.615
R450 VTAIL.n63 VTAIL.n17 104.615
R451 VTAIL.n64 VTAIL.n63 104.615
R452 VTAIL.n64 VTAIL.n13 104.615
R453 VTAIL.n71 VTAIL.n13 104.615
R454 VTAIL.n73 VTAIL.n71 104.615
R455 VTAIL.n73 VTAIL.n72 104.615
R456 VTAIL.n72 VTAIL.n9 104.615
R457 VTAIL.n81 VTAIL.n9 104.615
R458 VTAIL.n82 VTAIL.n81 104.615
R459 VTAIL.n82 VTAIL.n5 104.615
R460 VTAIL.n89 VTAIL.n5 104.615
R461 VTAIL.n90 VTAIL.n89 104.615
R462 VTAIL.n284 VTAIL.n283 104.615
R463 VTAIL.n283 VTAIL.n199 104.615
R464 VTAIL.n276 VTAIL.n199 104.615
R465 VTAIL.n276 VTAIL.n275 104.615
R466 VTAIL.n275 VTAIL.n203 104.615
R467 VTAIL.n207 VTAIL.n203 104.615
R468 VTAIL.n267 VTAIL.n207 104.615
R469 VTAIL.n267 VTAIL.n266 104.615
R470 VTAIL.n266 VTAIL.n208 104.615
R471 VTAIL.n259 VTAIL.n208 104.615
R472 VTAIL.n259 VTAIL.n258 104.615
R473 VTAIL.n258 VTAIL.n212 104.615
R474 VTAIL.n251 VTAIL.n212 104.615
R475 VTAIL.n251 VTAIL.n250 104.615
R476 VTAIL.n250 VTAIL.n216 104.615
R477 VTAIL.n243 VTAIL.n216 104.615
R478 VTAIL.n243 VTAIL.n242 104.615
R479 VTAIL.n242 VTAIL.n220 104.615
R480 VTAIL.n235 VTAIL.n220 104.615
R481 VTAIL.n235 VTAIL.n234 104.615
R482 VTAIL.n234 VTAIL.n224 104.615
R483 VTAIL.n227 VTAIL.n224 104.615
R484 VTAIL.n188 VTAIL.n187 104.615
R485 VTAIL.n187 VTAIL.n103 104.615
R486 VTAIL.n180 VTAIL.n103 104.615
R487 VTAIL.n180 VTAIL.n179 104.615
R488 VTAIL.n179 VTAIL.n107 104.615
R489 VTAIL.n111 VTAIL.n107 104.615
R490 VTAIL.n171 VTAIL.n111 104.615
R491 VTAIL.n171 VTAIL.n170 104.615
R492 VTAIL.n170 VTAIL.n112 104.615
R493 VTAIL.n163 VTAIL.n112 104.615
R494 VTAIL.n163 VTAIL.n162 104.615
R495 VTAIL.n162 VTAIL.n116 104.615
R496 VTAIL.n155 VTAIL.n116 104.615
R497 VTAIL.n155 VTAIL.n154 104.615
R498 VTAIL.n154 VTAIL.n120 104.615
R499 VTAIL.n147 VTAIL.n120 104.615
R500 VTAIL.n147 VTAIL.n146 104.615
R501 VTAIL.n146 VTAIL.n124 104.615
R502 VTAIL.n139 VTAIL.n124 104.615
R503 VTAIL.n139 VTAIL.n138 104.615
R504 VTAIL.n138 VTAIL.n128 104.615
R505 VTAIL.n131 VTAIL.n128 104.615
R506 VTAIL.n320 VTAIL.t6 52.3082
R507 VTAIL.n32 VTAIL.t4 52.3082
R508 VTAIL.n227 VTAIL.t0 52.3082
R509 VTAIL.n131 VTAIL.t8 52.3082
R510 VTAIL.n195 VTAIL.n194 44.6278
R511 VTAIL.n99 VTAIL.n98 44.6278
R512 VTAIL.n1 VTAIL.n0 44.6277
R513 VTAIL.n97 VTAIL.n96 44.6277
R514 VTAIL.n383 VTAIL.n382 32.7672
R515 VTAIL.n95 VTAIL.n94 32.7672
R516 VTAIL.n289 VTAIL.n288 32.7672
R517 VTAIL.n193 VTAIL.n192 32.7672
R518 VTAIL.n99 VTAIL.n97 28.9445
R519 VTAIL.n383 VTAIL.n289 27.91
R520 VTAIL.n321 VTAIL.n319 15.6677
R521 VTAIL.n33 VTAIL.n31 15.6677
R522 VTAIL.n228 VTAIL.n226 15.6677
R523 VTAIL.n132 VTAIL.n130 15.6677
R524 VTAIL.n368 VTAIL.n367 13.1884
R525 VTAIL.n80 VTAIL.n79 13.1884
R526 VTAIL.n274 VTAIL.n273 13.1884
R527 VTAIL.n178 VTAIL.n177 13.1884
R528 VTAIL.n322 VTAIL.n318 12.8005
R529 VTAIL.n366 VTAIL.n298 12.8005
R530 VTAIL.n371 VTAIL.n296 12.8005
R531 VTAIL.n34 VTAIL.n30 12.8005
R532 VTAIL.n78 VTAIL.n10 12.8005
R533 VTAIL.n83 VTAIL.n8 12.8005
R534 VTAIL.n277 VTAIL.n202 12.8005
R535 VTAIL.n272 VTAIL.n204 12.8005
R536 VTAIL.n229 VTAIL.n225 12.8005
R537 VTAIL.n181 VTAIL.n106 12.8005
R538 VTAIL.n176 VTAIL.n108 12.8005
R539 VTAIL.n133 VTAIL.n129 12.8005
R540 VTAIL.n326 VTAIL.n325 12.0247
R541 VTAIL.n363 VTAIL.n362 12.0247
R542 VTAIL.n372 VTAIL.n294 12.0247
R543 VTAIL.n38 VTAIL.n37 12.0247
R544 VTAIL.n75 VTAIL.n74 12.0247
R545 VTAIL.n84 VTAIL.n6 12.0247
R546 VTAIL.n278 VTAIL.n200 12.0247
R547 VTAIL.n269 VTAIL.n268 12.0247
R548 VTAIL.n233 VTAIL.n232 12.0247
R549 VTAIL.n182 VTAIL.n104 12.0247
R550 VTAIL.n173 VTAIL.n172 12.0247
R551 VTAIL.n137 VTAIL.n136 12.0247
R552 VTAIL.n329 VTAIL.n316 11.249
R553 VTAIL.n358 VTAIL.n300 11.249
R554 VTAIL.n376 VTAIL.n375 11.249
R555 VTAIL.n41 VTAIL.n28 11.249
R556 VTAIL.n70 VTAIL.n12 11.249
R557 VTAIL.n88 VTAIL.n87 11.249
R558 VTAIL.n282 VTAIL.n281 11.249
R559 VTAIL.n265 VTAIL.n206 11.249
R560 VTAIL.n236 VTAIL.n223 11.249
R561 VTAIL.n186 VTAIL.n185 11.249
R562 VTAIL.n169 VTAIL.n110 11.249
R563 VTAIL.n140 VTAIL.n127 11.249
R564 VTAIL.n330 VTAIL.n314 10.4732
R565 VTAIL.n357 VTAIL.n302 10.4732
R566 VTAIL.n379 VTAIL.n292 10.4732
R567 VTAIL.n42 VTAIL.n26 10.4732
R568 VTAIL.n69 VTAIL.n14 10.4732
R569 VTAIL.n91 VTAIL.n4 10.4732
R570 VTAIL.n285 VTAIL.n198 10.4732
R571 VTAIL.n264 VTAIL.n209 10.4732
R572 VTAIL.n237 VTAIL.n221 10.4732
R573 VTAIL.n189 VTAIL.n102 10.4732
R574 VTAIL.n168 VTAIL.n113 10.4732
R575 VTAIL.n141 VTAIL.n125 10.4732
R576 VTAIL.n334 VTAIL.n333 9.69747
R577 VTAIL.n354 VTAIL.n353 9.69747
R578 VTAIL.n380 VTAIL.n290 9.69747
R579 VTAIL.n46 VTAIL.n45 9.69747
R580 VTAIL.n66 VTAIL.n65 9.69747
R581 VTAIL.n92 VTAIL.n2 9.69747
R582 VTAIL.n286 VTAIL.n196 9.69747
R583 VTAIL.n261 VTAIL.n260 9.69747
R584 VTAIL.n241 VTAIL.n240 9.69747
R585 VTAIL.n190 VTAIL.n100 9.69747
R586 VTAIL.n165 VTAIL.n164 9.69747
R587 VTAIL.n145 VTAIL.n144 9.69747
R588 VTAIL.n382 VTAIL.n381 9.45567
R589 VTAIL.n94 VTAIL.n93 9.45567
R590 VTAIL.n288 VTAIL.n287 9.45567
R591 VTAIL.n192 VTAIL.n191 9.45567
R592 VTAIL.n381 VTAIL.n380 9.3005
R593 VTAIL.n292 VTAIL.n291 9.3005
R594 VTAIL.n375 VTAIL.n374 9.3005
R595 VTAIL.n373 VTAIL.n372 9.3005
R596 VTAIL.n296 VTAIL.n295 9.3005
R597 VTAIL.n341 VTAIL.n340 9.3005
R598 VTAIL.n339 VTAIL.n338 9.3005
R599 VTAIL.n312 VTAIL.n311 9.3005
R600 VTAIL.n333 VTAIL.n332 9.3005
R601 VTAIL.n331 VTAIL.n330 9.3005
R602 VTAIL.n316 VTAIL.n315 9.3005
R603 VTAIL.n325 VTAIL.n324 9.3005
R604 VTAIL.n323 VTAIL.n322 9.3005
R605 VTAIL.n308 VTAIL.n307 9.3005
R606 VTAIL.n347 VTAIL.n346 9.3005
R607 VTAIL.n349 VTAIL.n348 9.3005
R608 VTAIL.n304 VTAIL.n303 9.3005
R609 VTAIL.n355 VTAIL.n354 9.3005
R610 VTAIL.n357 VTAIL.n356 9.3005
R611 VTAIL.n300 VTAIL.n299 9.3005
R612 VTAIL.n364 VTAIL.n363 9.3005
R613 VTAIL.n366 VTAIL.n365 9.3005
R614 VTAIL.n93 VTAIL.n92 9.3005
R615 VTAIL.n4 VTAIL.n3 9.3005
R616 VTAIL.n87 VTAIL.n86 9.3005
R617 VTAIL.n85 VTAIL.n84 9.3005
R618 VTAIL.n8 VTAIL.n7 9.3005
R619 VTAIL.n53 VTAIL.n52 9.3005
R620 VTAIL.n51 VTAIL.n50 9.3005
R621 VTAIL.n24 VTAIL.n23 9.3005
R622 VTAIL.n45 VTAIL.n44 9.3005
R623 VTAIL.n43 VTAIL.n42 9.3005
R624 VTAIL.n28 VTAIL.n27 9.3005
R625 VTAIL.n37 VTAIL.n36 9.3005
R626 VTAIL.n35 VTAIL.n34 9.3005
R627 VTAIL.n20 VTAIL.n19 9.3005
R628 VTAIL.n59 VTAIL.n58 9.3005
R629 VTAIL.n61 VTAIL.n60 9.3005
R630 VTAIL.n16 VTAIL.n15 9.3005
R631 VTAIL.n67 VTAIL.n66 9.3005
R632 VTAIL.n69 VTAIL.n68 9.3005
R633 VTAIL.n12 VTAIL.n11 9.3005
R634 VTAIL.n76 VTAIL.n75 9.3005
R635 VTAIL.n78 VTAIL.n77 9.3005
R636 VTAIL.n254 VTAIL.n253 9.3005
R637 VTAIL.n256 VTAIL.n255 9.3005
R638 VTAIL.n211 VTAIL.n210 9.3005
R639 VTAIL.n262 VTAIL.n261 9.3005
R640 VTAIL.n264 VTAIL.n263 9.3005
R641 VTAIL.n206 VTAIL.n205 9.3005
R642 VTAIL.n270 VTAIL.n269 9.3005
R643 VTAIL.n272 VTAIL.n271 9.3005
R644 VTAIL.n287 VTAIL.n286 9.3005
R645 VTAIL.n198 VTAIL.n197 9.3005
R646 VTAIL.n281 VTAIL.n280 9.3005
R647 VTAIL.n279 VTAIL.n278 9.3005
R648 VTAIL.n202 VTAIL.n201 9.3005
R649 VTAIL.n215 VTAIL.n214 9.3005
R650 VTAIL.n248 VTAIL.n247 9.3005
R651 VTAIL.n246 VTAIL.n245 9.3005
R652 VTAIL.n219 VTAIL.n218 9.3005
R653 VTAIL.n240 VTAIL.n239 9.3005
R654 VTAIL.n238 VTAIL.n237 9.3005
R655 VTAIL.n223 VTAIL.n222 9.3005
R656 VTAIL.n232 VTAIL.n231 9.3005
R657 VTAIL.n230 VTAIL.n229 9.3005
R658 VTAIL.n158 VTAIL.n157 9.3005
R659 VTAIL.n160 VTAIL.n159 9.3005
R660 VTAIL.n115 VTAIL.n114 9.3005
R661 VTAIL.n166 VTAIL.n165 9.3005
R662 VTAIL.n168 VTAIL.n167 9.3005
R663 VTAIL.n110 VTAIL.n109 9.3005
R664 VTAIL.n174 VTAIL.n173 9.3005
R665 VTAIL.n176 VTAIL.n175 9.3005
R666 VTAIL.n191 VTAIL.n190 9.3005
R667 VTAIL.n102 VTAIL.n101 9.3005
R668 VTAIL.n185 VTAIL.n184 9.3005
R669 VTAIL.n183 VTAIL.n182 9.3005
R670 VTAIL.n106 VTAIL.n105 9.3005
R671 VTAIL.n119 VTAIL.n118 9.3005
R672 VTAIL.n152 VTAIL.n151 9.3005
R673 VTAIL.n150 VTAIL.n149 9.3005
R674 VTAIL.n123 VTAIL.n122 9.3005
R675 VTAIL.n144 VTAIL.n143 9.3005
R676 VTAIL.n142 VTAIL.n141 9.3005
R677 VTAIL.n127 VTAIL.n126 9.3005
R678 VTAIL.n136 VTAIL.n135 9.3005
R679 VTAIL.n134 VTAIL.n133 9.3005
R680 VTAIL.n337 VTAIL.n312 8.92171
R681 VTAIL.n350 VTAIL.n304 8.92171
R682 VTAIL.n49 VTAIL.n24 8.92171
R683 VTAIL.n62 VTAIL.n16 8.92171
R684 VTAIL.n257 VTAIL.n211 8.92171
R685 VTAIL.n244 VTAIL.n219 8.92171
R686 VTAIL.n161 VTAIL.n115 8.92171
R687 VTAIL.n148 VTAIL.n123 8.92171
R688 VTAIL.n338 VTAIL.n310 8.14595
R689 VTAIL.n349 VTAIL.n306 8.14595
R690 VTAIL.n50 VTAIL.n22 8.14595
R691 VTAIL.n61 VTAIL.n18 8.14595
R692 VTAIL.n256 VTAIL.n213 8.14595
R693 VTAIL.n245 VTAIL.n217 8.14595
R694 VTAIL.n160 VTAIL.n117 8.14595
R695 VTAIL.n149 VTAIL.n121 8.14595
R696 VTAIL.n342 VTAIL.n341 7.3702
R697 VTAIL.n346 VTAIL.n345 7.3702
R698 VTAIL.n54 VTAIL.n53 7.3702
R699 VTAIL.n58 VTAIL.n57 7.3702
R700 VTAIL.n253 VTAIL.n252 7.3702
R701 VTAIL.n249 VTAIL.n248 7.3702
R702 VTAIL.n157 VTAIL.n156 7.3702
R703 VTAIL.n153 VTAIL.n152 7.3702
R704 VTAIL.n342 VTAIL.n308 6.59444
R705 VTAIL.n345 VTAIL.n308 6.59444
R706 VTAIL.n54 VTAIL.n20 6.59444
R707 VTAIL.n57 VTAIL.n20 6.59444
R708 VTAIL.n252 VTAIL.n215 6.59444
R709 VTAIL.n249 VTAIL.n215 6.59444
R710 VTAIL.n156 VTAIL.n119 6.59444
R711 VTAIL.n153 VTAIL.n119 6.59444
R712 VTAIL.n341 VTAIL.n310 5.81868
R713 VTAIL.n346 VTAIL.n306 5.81868
R714 VTAIL.n53 VTAIL.n22 5.81868
R715 VTAIL.n58 VTAIL.n18 5.81868
R716 VTAIL.n253 VTAIL.n213 5.81868
R717 VTAIL.n248 VTAIL.n217 5.81868
R718 VTAIL.n157 VTAIL.n117 5.81868
R719 VTAIL.n152 VTAIL.n121 5.81868
R720 VTAIL.n338 VTAIL.n337 5.04292
R721 VTAIL.n350 VTAIL.n349 5.04292
R722 VTAIL.n50 VTAIL.n49 5.04292
R723 VTAIL.n62 VTAIL.n61 5.04292
R724 VTAIL.n257 VTAIL.n256 5.04292
R725 VTAIL.n245 VTAIL.n244 5.04292
R726 VTAIL.n161 VTAIL.n160 5.04292
R727 VTAIL.n149 VTAIL.n148 5.04292
R728 VTAIL.n230 VTAIL.n226 4.38563
R729 VTAIL.n134 VTAIL.n130 4.38563
R730 VTAIL.n323 VTAIL.n319 4.38563
R731 VTAIL.n35 VTAIL.n31 4.38563
R732 VTAIL.n334 VTAIL.n312 4.26717
R733 VTAIL.n353 VTAIL.n304 4.26717
R734 VTAIL.n382 VTAIL.n290 4.26717
R735 VTAIL.n46 VTAIL.n24 4.26717
R736 VTAIL.n65 VTAIL.n16 4.26717
R737 VTAIL.n94 VTAIL.n2 4.26717
R738 VTAIL.n288 VTAIL.n196 4.26717
R739 VTAIL.n260 VTAIL.n211 4.26717
R740 VTAIL.n241 VTAIL.n219 4.26717
R741 VTAIL.n192 VTAIL.n100 4.26717
R742 VTAIL.n164 VTAIL.n115 4.26717
R743 VTAIL.n145 VTAIL.n123 4.26717
R744 VTAIL.n333 VTAIL.n314 3.49141
R745 VTAIL.n354 VTAIL.n302 3.49141
R746 VTAIL.n380 VTAIL.n379 3.49141
R747 VTAIL.n45 VTAIL.n26 3.49141
R748 VTAIL.n66 VTAIL.n14 3.49141
R749 VTAIL.n92 VTAIL.n91 3.49141
R750 VTAIL.n286 VTAIL.n285 3.49141
R751 VTAIL.n261 VTAIL.n209 3.49141
R752 VTAIL.n240 VTAIL.n221 3.49141
R753 VTAIL.n190 VTAIL.n189 3.49141
R754 VTAIL.n165 VTAIL.n113 3.49141
R755 VTAIL.n144 VTAIL.n125 3.49141
R756 VTAIL.n330 VTAIL.n329 2.71565
R757 VTAIL.n358 VTAIL.n357 2.71565
R758 VTAIL.n376 VTAIL.n292 2.71565
R759 VTAIL.n42 VTAIL.n41 2.71565
R760 VTAIL.n70 VTAIL.n69 2.71565
R761 VTAIL.n88 VTAIL.n4 2.71565
R762 VTAIL.n282 VTAIL.n198 2.71565
R763 VTAIL.n265 VTAIL.n264 2.71565
R764 VTAIL.n237 VTAIL.n236 2.71565
R765 VTAIL.n186 VTAIL.n102 2.71565
R766 VTAIL.n169 VTAIL.n168 2.71565
R767 VTAIL.n141 VTAIL.n140 2.71565
R768 VTAIL.n326 VTAIL.n316 1.93989
R769 VTAIL.n362 VTAIL.n300 1.93989
R770 VTAIL.n375 VTAIL.n294 1.93989
R771 VTAIL.n38 VTAIL.n28 1.93989
R772 VTAIL.n74 VTAIL.n12 1.93989
R773 VTAIL.n87 VTAIL.n6 1.93989
R774 VTAIL.n281 VTAIL.n200 1.93989
R775 VTAIL.n268 VTAIL.n206 1.93989
R776 VTAIL.n233 VTAIL.n223 1.93989
R777 VTAIL.n185 VTAIL.n104 1.93989
R778 VTAIL.n172 VTAIL.n110 1.93989
R779 VTAIL.n137 VTAIL.n127 1.93989
R780 VTAIL.n0 VTAIL.t9 1.17697
R781 VTAIL.n0 VTAIL.t5 1.17697
R782 VTAIL.n96 VTAIL.t2 1.17697
R783 VTAIL.n96 VTAIL.t3 1.17697
R784 VTAIL.n194 VTAIL.t1 1.17697
R785 VTAIL.n194 VTAIL.t11 1.17697
R786 VTAIL.n98 VTAIL.t7 1.17697
R787 VTAIL.n98 VTAIL.t10 1.17697
R788 VTAIL.n325 VTAIL.n318 1.16414
R789 VTAIL.n363 VTAIL.n298 1.16414
R790 VTAIL.n372 VTAIL.n371 1.16414
R791 VTAIL.n37 VTAIL.n30 1.16414
R792 VTAIL.n75 VTAIL.n10 1.16414
R793 VTAIL.n84 VTAIL.n83 1.16414
R794 VTAIL.n278 VTAIL.n277 1.16414
R795 VTAIL.n269 VTAIL.n204 1.16414
R796 VTAIL.n232 VTAIL.n225 1.16414
R797 VTAIL.n182 VTAIL.n181 1.16414
R798 VTAIL.n173 VTAIL.n108 1.16414
R799 VTAIL.n136 VTAIL.n129 1.16414
R800 VTAIL.n193 VTAIL.n99 1.03498
R801 VTAIL.n289 VTAIL.n195 1.03498
R802 VTAIL.n97 VTAIL.n95 1.03498
R803 VTAIL.n195 VTAIL.n193 0.987569
R804 VTAIL.n95 VTAIL.n1 0.987569
R805 VTAIL VTAIL.n383 0.718172
R806 VTAIL.n322 VTAIL.n321 0.388379
R807 VTAIL.n367 VTAIL.n366 0.388379
R808 VTAIL.n368 VTAIL.n296 0.388379
R809 VTAIL.n34 VTAIL.n33 0.388379
R810 VTAIL.n79 VTAIL.n78 0.388379
R811 VTAIL.n80 VTAIL.n8 0.388379
R812 VTAIL.n274 VTAIL.n202 0.388379
R813 VTAIL.n273 VTAIL.n272 0.388379
R814 VTAIL.n229 VTAIL.n228 0.388379
R815 VTAIL.n178 VTAIL.n106 0.388379
R816 VTAIL.n177 VTAIL.n176 0.388379
R817 VTAIL.n133 VTAIL.n132 0.388379
R818 VTAIL VTAIL.n1 0.31731
R819 VTAIL.n324 VTAIL.n323 0.155672
R820 VTAIL.n324 VTAIL.n315 0.155672
R821 VTAIL.n331 VTAIL.n315 0.155672
R822 VTAIL.n332 VTAIL.n331 0.155672
R823 VTAIL.n332 VTAIL.n311 0.155672
R824 VTAIL.n339 VTAIL.n311 0.155672
R825 VTAIL.n340 VTAIL.n339 0.155672
R826 VTAIL.n340 VTAIL.n307 0.155672
R827 VTAIL.n347 VTAIL.n307 0.155672
R828 VTAIL.n348 VTAIL.n347 0.155672
R829 VTAIL.n348 VTAIL.n303 0.155672
R830 VTAIL.n355 VTAIL.n303 0.155672
R831 VTAIL.n356 VTAIL.n355 0.155672
R832 VTAIL.n356 VTAIL.n299 0.155672
R833 VTAIL.n364 VTAIL.n299 0.155672
R834 VTAIL.n365 VTAIL.n364 0.155672
R835 VTAIL.n365 VTAIL.n295 0.155672
R836 VTAIL.n373 VTAIL.n295 0.155672
R837 VTAIL.n374 VTAIL.n373 0.155672
R838 VTAIL.n374 VTAIL.n291 0.155672
R839 VTAIL.n381 VTAIL.n291 0.155672
R840 VTAIL.n36 VTAIL.n35 0.155672
R841 VTAIL.n36 VTAIL.n27 0.155672
R842 VTAIL.n43 VTAIL.n27 0.155672
R843 VTAIL.n44 VTAIL.n43 0.155672
R844 VTAIL.n44 VTAIL.n23 0.155672
R845 VTAIL.n51 VTAIL.n23 0.155672
R846 VTAIL.n52 VTAIL.n51 0.155672
R847 VTAIL.n52 VTAIL.n19 0.155672
R848 VTAIL.n59 VTAIL.n19 0.155672
R849 VTAIL.n60 VTAIL.n59 0.155672
R850 VTAIL.n60 VTAIL.n15 0.155672
R851 VTAIL.n67 VTAIL.n15 0.155672
R852 VTAIL.n68 VTAIL.n67 0.155672
R853 VTAIL.n68 VTAIL.n11 0.155672
R854 VTAIL.n76 VTAIL.n11 0.155672
R855 VTAIL.n77 VTAIL.n76 0.155672
R856 VTAIL.n77 VTAIL.n7 0.155672
R857 VTAIL.n85 VTAIL.n7 0.155672
R858 VTAIL.n86 VTAIL.n85 0.155672
R859 VTAIL.n86 VTAIL.n3 0.155672
R860 VTAIL.n93 VTAIL.n3 0.155672
R861 VTAIL.n287 VTAIL.n197 0.155672
R862 VTAIL.n280 VTAIL.n197 0.155672
R863 VTAIL.n280 VTAIL.n279 0.155672
R864 VTAIL.n279 VTAIL.n201 0.155672
R865 VTAIL.n271 VTAIL.n201 0.155672
R866 VTAIL.n271 VTAIL.n270 0.155672
R867 VTAIL.n270 VTAIL.n205 0.155672
R868 VTAIL.n263 VTAIL.n205 0.155672
R869 VTAIL.n263 VTAIL.n262 0.155672
R870 VTAIL.n262 VTAIL.n210 0.155672
R871 VTAIL.n255 VTAIL.n210 0.155672
R872 VTAIL.n255 VTAIL.n254 0.155672
R873 VTAIL.n254 VTAIL.n214 0.155672
R874 VTAIL.n247 VTAIL.n214 0.155672
R875 VTAIL.n247 VTAIL.n246 0.155672
R876 VTAIL.n246 VTAIL.n218 0.155672
R877 VTAIL.n239 VTAIL.n218 0.155672
R878 VTAIL.n239 VTAIL.n238 0.155672
R879 VTAIL.n238 VTAIL.n222 0.155672
R880 VTAIL.n231 VTAIL.n222 0.155672
R881 VTAIL.n231 VTAIL.n230 0.155672
R882 VTAIL.n191 VTAIL.n101 0.155672
R883 VTAIL.n184 VTAIL.n101 0.155672
R884 VTAIL.n184 VTAIL.n183 0.155672
R885 VTAIL.n183 VTAIL.n105 0.155672
R886 VTAIL.n175 VTAIL.n105 0.155672
R887 VTAIL.n175 VTAIL.n174 0.155672
R888 VTAIL.n174 VTAIL.n109 0.155672
R889 VTAIL.n167 VTAIL.n109 0.155672
R890 VTAIL.n167 VTAIL.n166 0.155672
R891 VTAIL.n166 VTAIL.n114 0.155672
R892 VTAIL.n159 VTAIL.n114 0.155672
R893 VTAIL.n159 VTAIL.n158 0.155672
R894 VTAIL.n158 VTAIL.n118 0.155672
R895 VTAIL.n151 VTAIL.n118 0.155672
R896 VTAIL.n151 VTAIL.n150 0.155672
R897 VTAIL.n150 VTAIL.n122 0.155672
R898 VTAIL.n143 VTAIL.n122 0.155672
R899 VTAIL.n143 VTAIL.n142 0.155672
R900 VTAIL.n142 VTAIL.n126 0.155672
R901 VTAIL.n135 VTAIL.n126 0.155672
R902 VTAIL.n135 VTAIL.n134 0.155672
R903 B.n185 B.t17 668.167
R904 B.n179 B.t10 668.167
R905 B.n73 B.t14 668.167
R906 B.n79 B.t6 668.167
R907 B.n553 B.n108 585
R908 B.n108 B.n43 585
R909 B.n555 B.n554 585
R910 B.n557 B.n107 585
R911 B.n560 B.n559 585
R912 B.n561 B.n106 585
R913 B.n563 B.n562 585
R914 B.n565 B.n105 585
R915 B.n568 B.n567 585
R916 B.n569 B.n104 585
R917 B.n571 B.n570 585
R918 B.n573 B.n103 585
R919 B.n576 B.n575 585
R920 B.n577 B.n102 585
R921 B.n579 B.n578 585
R922 B.n581 B.n101 585
R923 B.n584 B.n583 585
R924 B.n585 B.n100 585
R925 B.n587 B.n586 585
R926 B.n589 B.n99 585
R927 B.n592 B.n591 585
R928 B.n593 B.n98 585
R929 B.n595 B.n594 585
R930 B.n597 B.n97 585
R931 B.n600 B.n599 585
R932 B.n601 B.n96 585
R933 B.n603 B.n602 585
R934 B.n605 B.n95 585
R935 B.n608 B.n607 585
R936 B.n609 B.n94 585
R937 B.n611 B.n610 585
R938 B.n613 B.n93 585
R939 B.n616 B.n615 585
R940 B.n617 B.n92 585
R941 B.n619 B.n618 585
R942 B.n621 B.n91 585
R943 B.n624 B.n623 585
R944 B.n625 B.n90 585
R945 B.n627 B.n626 585
R946 B.n629 B.n89 585
R947 B.n632 B.n631 585
R948 B.n633 B.n88 585
R949 B.n635 B.n634 585
R950 B.n637 B.n87 585
R951 B.n640 B.n639 585
R952 B.n641 B.n86 585
R953 B.n643 B.n642 585
R954 B.n645 B.n85 585
R955 B.n648 B.n647 585
R956 B.n649 B.n84 585
R957 B.n651 B.n650 585
R958 B.n653 B.n83 585
R959 B.n656 B.n655 585
R960 B.n657 B.n82 585
R961 B.n659 B.n658 585
R962 B.n661 B.n81 585
R963 B.n664 B.n663 585
R964 B.n666 B.n78 585
R965 B.n668 B.n667 585
R966 B.n670 B.n77 585
R967 B.n673 B.n672 585
R968 B.n674 B.n76 585
R969 B.n676 B.n675 585
R970 B.n678 B.n75 585
R971 B.n681 B.n680 585
R972 B.n682 B.n72 585
R973 B.n685 B.n684 585
R974 B.n687 B.n71 585
R975 B.n690 B.n689 585
R976 B.n691 B.n70 585
R977 B.n693 B.n692 585
R978 B.n695 B.n69 585
R979 B.n698 B.n697 585
R980 B.n699 B.n68 585
R981 B.n701 B.n700 585
R982 B.n703 B.n67 585
R983 B.n706 B.n705 585
R984 B.n707 B.n66 585
R985 B.n709 B.n708 585
R986 B.n711 B.n65 585
R987 B.n714 B.n713 585
R988 B.n715 B.n64 585
R989 B.n717 B.n716 585
R990 B.n719 B.n63 585
R991 B.n722 B.n721 585
R992 B.n723 B.n62 585
R993 B.n725 B.n724 585
R994 B.n727 B.n61 585
R995 B.n730 B.n729 585
R996 B.n731 B.n60 585
R997 B.n733 B.n732 585
R998 B.n735 B.n59 585
R999 B.n738 B.n737 585
R1000 B.n739 B.n58 585
R1001 B.n741 B.n740 585
R1002 B.n743 B.n57 585
R1003 B.n746 B.n745 585
R1004 B.n747 B.n56 585
R1005 B.n749 B.n748 585
R1006 B.n751 B.n55 585
R1007 B.n754 B.n753 585
R1008 B.n755 B.n54 585
R1009 B.n757 B.n756 585
R1010 B.n759 B.n53 585
R1011 B.n762 B.n761 585
R1012 B.n763 B.n52 585
R1013 B.n765 B.n764 585
R1014 B.n767 B.n51 585
R1015 B.n770 B.n769 585
R1016 B.n771 B.n50 585
R1017 B.n773 B.n772 585
R1018 B.n775 B.n49 585
R1019 B.n778 B.n777 585
R1020 B.n779 B.n48 585
R1021 B.n781 B.n780 585
R1022 B.n783 B.n47 585
R1023 B.n786 B.n785 585
R1024 B.n787 B.n46 585
R1025 B.n789 B.n788 585
R1026 B.n791 B.n45 585
R1027 B.n794 B.n793 585
R1028 B.n795 B.n44 585
R1029 B.n552 B.n42 585
R1030 B.n798 B.n42 585
R1031 B.n551 B.n41 585
R1032 B.n799 B.n41 585
R1033 B.n550 B.n40 585
R1034 B.n800 B.n40 585
R1035 B.n549 B.n548 585
R1036 B.n548 B.n36 585
R1037 B.n547 B.n35 585
R1038 B.n806 B.n35 585
R1039 B.n546 B.n34 585
R1040 B.n807 B.n34 585
R1041 B.n545 B.n33 585
R1042 B.n808 B.n33 585
R1043 B.n544 B.n543 585
R1044 B.n543 B.n29 585
R1045 B.n542 B.n28 585
R1046 B.n814 B.n28 585
R1047 B.n541 B.n27 585
R1048 B.n815 B.n27 585
R1049 B.n540 B.n26 585
R1050 B.n816 B.n26 585
R1051 B.n539 B.n538 585
R1052 B.n538 B.n25 585
R1053 B.n537 B.n21 585
R1054 B.n822 B.n21 585
R1055 B.n536 B.n20 585
R1056 B.n823 B.n20 585
R1057 B.n535 B.n19 585
R1058 B.n824 B.n19 585
R1059 B.n534 B.n533 585
R1060 B.n533 B.n18 585
R1061 B.n532 B.n14 585
R1062 B.n830 B.n14 585
R1063 B.n531 B.n13 585
R1064 B.n831 B.n13 585
R1065 B.n530 B.n12 585
R1066 B.n832 B.n12 585
R1067 B.n529 B.n528 585
R1068 B.n528 B.n8 585
R1069 B.n527 B.n7 585
R1070 B.n838 B.n7 585
R1071 B.n526 B.n6 585
R1072 B.n839 B.n6 585
R1073 B.n525 B.n5 585
R1074 B.n840 B.n5 585
R1075 B.n524 B.n523 585
R1076 B.n523 B.n4 585
R1077 B.n522 B.n109 585
R1078 B.n522 B.n521 585
R1079 B.n512 B.n110 585
R1080 B.n111 B.n110 585
R1081 B.n514 B.n513 585
R1082 B.n515 B.n514 585
R1083 B.n511 B.n116 585
R1084 B.n116 B.n115 585
R1085 B.n510 B.n509 585
R1086 B.n509 B.n508 585
R1087 B.n118 B.n117 585
R1088 B.n501 B.n118 585
R1089 B.n500 B.n499 585
R1090 B.n502 B.n500 585
R1091 B.n498 B.n123 585
R1092 B.n123 B.n122 585
R1093 B.n497 B.n496 585
R1094 B.n496 B.n495 585
R1095 B.n125 B.n124 585
R1096 B.n488 B.n125 585
R1097 B.n487 B.n486 585
R1098 B.n489 B.n487 585
R1099 B.n485 B.n130 585
R1100 B.n130 B.n129 585
R1101 B.n484 B.n483 585
R1102 B.n483 B.n482 585
R1103 B.n132 B.n131 585
R1104 B.n133 B.n132 585
R1105 B.n475 B.n474 585
R1106 B.n476 B.n475 585
R1107 B.n473 B.n138 585
R1108 B.n138 B.n137 585
R1109 B.n472 B.n471 585
R1110 B.n471 B.n470 585
R1111 B.n140 B.n139 585
R1112 B.n141 B.n140 585
R1113 B.n463 B.n462 585
R1114 B.n464 B.n463 585
R1115 B.n461 B.n146 585
R1116 B.n146 B.n145 585
R1117 B.n460 B.n459 585
R1118 B.n459 B.n458 585
R1119 B.n455 B.n150 585
R1120 B.n454 B.n453 585
R1121 B.n451 B.n151 585
R1122 B.n451 B.n149 585
R1123 B.n450 B.n449 585
R1124 B.n448 B.n447 585
R1125 B.n446 B.n153 585
R1126 B.n444 B.n443 585
R1127 B.n442 B.n154 585
R1128 B.n441 B.n440 585
R1129 B.n438 B.n155 585
R1130 B.n436 B.n435 585
R1131 B.n434 B.n156 585
R1132 B.n433 B.n432 585
R1133 B.n430 B.n157 585
R1134 B.n428 B.n427 585
R1135 B.n426 B.n158 585
R1136 B.n425 B.n424 585
R1137 B.n422 B.n159 585
R1138 B.n420 B.n419 585
R1139 B.n418 B.n160 585
R1140 B.n417 B.n416 585
R1141 B.n414 B.n161 585
R1142 B.n412 B.n411 585
R1143 B.n410 B.n162 585
R1144 B.n409 B.n408 585
R1145 B.n406 B.n163 585
R1146 B.n404 B.n403 585
R1147 B.n402 B.n164 585
R1148 B.n401 B.n400 585
R1149 B.n398 B.n165 585
R1150 B.n396 B.n395 585
R1151 B.n394 B.n166 585
R1152 B.n393 B.n392 585
R1153 B.n390 B.n167 585
R1154 B.n388 B.n387 585
R1155 B.n386 B.n168 585
R1156 B.n385 B.n384 585
R1157 B.n382 B.n169 585
R1158 B.n380 B.n379 585
R1159 B.n378 B.n170 585
R1160 B.n377 B.n376 585
R1161 B.n374 B.n171 585
R1162 B.n372 B.n371 585
R1163 B.n370 B.n172 585
R1164 B.n369 B.n368 585
R1165 B.n366 B.n173 585
R1166 B.n364 B.n363 585
R1167 B.n362 B.n174 585
R1168 B.n361 B.n360 585
R1169 B.n358 B.n175 585
R1170 B.n356 B.n355 585
R1171 B.n354 B.n176 585
R1172 B.n353 B.n352 585
R1173 B.n350 B.n177 585
R1174 B.n348 B.n347 585
R1175 B.n346 B.n178 585
R1176 B.n344 B.n343 585
R1177 B.n341 B.n181 585
R1178 B.n339 B.n338 585
R1179 B.n337 B.n182 585
R1180 B.n336 B.n335 585
R1181 B.n333 B.n183 585
R1182 B.n331 B.n330 585
R1183 B.n329 B.n184 585
R1184 B.n328 B.n327 585
R1185 B.n325 B.n324 585
R1186 B.n323 B.n322 585
R1187 B.n321 B.n189 585
R1188 B.n319 B.n318 585
R1189 B.n317 B.n190 585
R1190 B.n316 B.n315 585
R1191 B.n313 B.n191 585
R1192 B.n311 B.n310 585
R1193 B.n309 B.n192 585
R1194 B.n308 B.n307 585
R1195 B.n305 B.n193 585
R1196 B.n303 B.n302 585
R1197 B.n301 B.n194 585
R1198 B.n300 B.n299 585
R1199 B.n297 B.n195 585
R1200 B.n295 B.n294 585
R1201 B.n293 B.n196 585
R1202 B.n292 B.n291 585
R1203 B.n289 B.n197 585
R1204 B.n287 B.n286 585
R1205 B.n285 B.n198 585
R1206 B.n284 B.n283 585
R1207 B.n281 B.n199 585
R1208 B.n279 B.n278 585
R1209 B.n277 B.n200 585
R1210 B.n276 B.n275 585
R1211 B.n273 B.n201 585
R1212 B.n271 B.n270 585
R1213 B.n269 B.n202 585
R1214 B.n268 B.n267 585
R1215 B.n265 B.n203 585
R1216 B.n263 B.n262 585
R1217 B.n261 B.n204 585
R1218 B.n260 B.n259 585
R1219 B.n257 B.n205 585
R1220 B.n255 B.n254 585
R1221 B.n253 B.n206 585
R1222 B.n252 B.n251 585
R1223 B.n249 B.n207 585
R1224 B.n247 B.n246 585
R1225 B.n245 B.n208 585
R1226 B.n244 B.n243 585
R1227 B.n241 B.n209 585
R1228 B.n239 B.n238 585
R1229 B.n237 B.n210 585
R1230 B.n236 B.n235 585
R1231 B.n233 B.n211 585
R1232 B.n231 B.n230 585
R1233 B.n229 B.n212 585
R1234 B.n228 B.n227 585
R1235 B.n225 B.n213 585
R1236 B.n223 B.n222 585
R1237 B.n221 B.n214 585
R1238 B.n220 B.n219 585
R1239 B.n217 B.n215 585
R1240 B.n148 B.n147 585
R1241 B.n457 B.n456 585
R1242 B.n458 B.n457 585
R1243 B.n144 B.n143 585
R1244 B.n145 B.n144 585
R1245 B.n466 B.n465 585
R1246 B.n465 B.n464 585
R1247 B.n467 B.n142 585
R1248 B.n142 B.n141 585
R1249 B.n469 B.n468 585
R1250 B.n470 B.n469 585
R1251 B.n136 B.n135 585
R1252 B.n137 B.n136 585
R1253 B.n478 B.n477 585
R1254 B.n477 B.n476 585
R1255 B.n479 B.n134 585
R1256 B.n134 B.n133 585
R1257 B.n481 B.n480 585
R1258 B.n482 B.n481 585
R1259 B.n128 B.n127 585
R1260 B.n129 B.n128 585
R1261 B.n491 B.n490 585
R1262 B.n490 B.n489 585
R1263 B.n492 B.n126 585
R1264 B.n488 B.n126 585
R1265 B.n494 B.n493 585
R1266 B.n495 B.n494 585
R1267 B.n121 B.n120 585
R1268 B.n122 B.n121 585
R1269 B.n504 B.n503 585
R1270 B.n503 B.n502 585
R1271 B.n505 B.n119 585
R1272 B.n501 B.n119 585
R1273 B.n507 B.n506 585
R1274 B.n508 B.n507 585
R1275 B.n114 B.n113 585
R1276 B.n115 B.n114 585
R1277 B.n517 B.n516 585
R1278 B.n516 B.n515 585
R1279 B.n518 B.n112 585
R1280 B.n112 B.n111 585
R1281 B.n520 B.n519 585
R1282 B.n521 B.n520 585
R1283 B.n2 B.n0 585
R1284 B.n4 B.n2 585
R1285 B.n3 B.n1 585
R1286 B.n839 B.n3 585
R1287 B.n837 B.n836 585
R1288 B.n838 B.n837 585
R1289 B.n835 B.n9 585
R1290 B.n9 B.n8 585
R1291 B.n834 B.n833 585
R1292 B.n833 B.n832 585
R1293 B.n11 B.n10 585
R1294 B.n831 B.n11 585
R1295 B.n829 B.n828 585
R1296 B.n830 B.n829 585
R1297 B.n827 B.n15 585
R1298 B.n18 B.n15 585
R1299 B.n826 B.n825 585
R1300 B.n825 B.n824 585
R1301 B.n17 B.n16 585
R1302 B.n823 B.n17 585
R1303 B.n821 B.n820 585
R1304 B.n822 B.n821 585
R1305 B.n819 B.n22 585
R1306 B.n25 B.n22 585
R1307 B.n818 B.n817 585
R1308 B.n817 B.n816 585
R1309 B.n24 B.n23 585
R1310 B.n815 B.n24 585
R1311 B.n813 B.n812 585
R1312 B.n814 B.n813 585
R1313 B.n811 B.n30 585
R1314 B.n30 B.n29 585
R1315 B.n810 B.n809 585
R1316 B.n809 B.n808 585
R1317 B.n32 B.n31 585
R1318 B.n807 B.n32 585
R1319 B.n805 B.n804 585
R1320 B.n806 B.n805 585
R1321 B.n803 B.n37 585
R1322 B.n37 B.n36 585
R1323 B.n802 B.n801 585
R1324 B.n801 B.n800 585
R1325 B.n39 B.n38 585
R1326 B.n799 B.n39 585
R1327 B.n797 B.n796 585
R1328 B.n798 B.n797 585
R1329 B.n842 B.n841 585
R1330 B.n841 B.n840 585
R1331 B.n457 B.n150 554.963
R1332 B.n797 B.n44 554.963
R1333 B.n459 B.n148 554.963
R1334 B.n108 B.n42 554.963
R1335 B.n185 B.t19 388.625
R1336 B.n79 B.t8 388.625
R1337 B.n179 B.t13 388.625
R1338 B.n73 B.t15 388.625
R1339 B.n186 B.t18 365.353
R1340 B.n80 B.t9 365.353
R1341 B.n180 B.t12 365.353
R1342 B.n74 B.t16 365.353
R1343 B.n556 B.n43 256.663
R1344 B.n558 B.n43 256.663
R1345 B.n564 B.n43 256.663
R1346 B.n566 B.n43 256.663
R1347 B.n572 B.n43 256.663
R1348 B.n574 B.n43 256.663
R1349 B.n580 B.n43 256.663
R1350 B.n582 B.n43 256.663
R1351 B.n588 B.n43 256.663
R1352 B.n590 B.n43 256.663
R1353 B.n596 B.n43 256.663
R1354 B.n598 B.n43 256.663
R1355 B.n604 B.n43 256.663
R1356 B.n606 B.n43 256.663
R1357 B.n612 B.n43 256.663
R1358 B.n614 B.n43 256.663
R1359 B.n620 B.n43 256.663
R1360 B.n622 B.n43 256.663
R1361 B.n628 B.n43 256.663
R1362 B.n630 B.n43 256.663
R1363 B.n636 B.n43 256.663
R1364 B.n638 B.n43 256.663
R1365 B.n644 B.n43 256.663
R1366 B.n646 B.n43 256.663
R1367 B.n652 B.n43 256.663
R1368 B.n654 B.n43 256.663
R1369 B.n660 B.n43 256.663
R1370 B.n662 B.n43 256.663
R1371 B.n669 B.n43 256.663
R1372 B.n671 B.n43 256.663
R1373 B.n677 B.n43 256.663
R1374 B.n679 B.n43 256.663
R1375 B.n686 B.n43 256.663
R1376 B.n688 B.n43 256.663
R1377 B.n694 B.n43 256.663
R1378 B.n696 B.n43 256.663
R1379 B.n702 B.n43 256.663
R1380 B.n704 B.n43 256.663
R1381 B.n710 B.n43 256.663
R1382 B.n712 B.n43 256.663
R1383 B.n718 B.n43 256.663
R1384 B.n720 B.n43 256.663
R1385 B.n726 B.n43 256.663
R1386 B.n728 B.n43 256.663
R1387 B.n734 B.n43 256.663
R1388 B.n736 B.n43 256.663
R1389 B.n742 B.n43 256.663
R1390 B.n744 B.n43 256.663
R1391 B.n750 B.n43 256.663
R1392 B.n752 B.n43 256.663
R1393 B.n758 B.n43 256.663
R1394 B.n760 B.n43 256.663
R1395 B.n766 B.n43 256.663
R1396 B.n768 B.n43 256.663
R1397 B.n774 B.n43 256.663
R1398 B.n776 B.n43 256.663
R1399 B.n782 B.n43 256.663
R1400 B.n784 B.n43 256.663
R1401 B.n790 B.n43 256.663
R1402 B.n792 B.n43 256.663
R1403 B.n452 B.n149 256.663
R1404 B.n152 B.n149 256.663
R1405 B.n445 B.n149 256.663
R1406 B.n439 B.n149 256.663
R1407 B.n437 B.n149 256.663
R1408 B.n431 B.n149 256.663
R1409 B.n429 B.n149 256.663
R1410 B.n423 B.n149 256.663
R1411 B.n421 B.n149 256.663
R1412 B.n415 B.n149 256.663
R1413 B.n413 B.n149 256.663
R1414 B.n407 B.n149 256.663
R1415 B.n405 B.n149 256.663
R1416 B.n399 B.n149 256.663
R1417 B.n397 B.n149 256.663
R1418 B.n391 B.n149 256.663
R1419 B.n389 B.n149 256.663
R1420 B.n383 B.n149 256.663
R1421 B.n381 B.n149 256.663
R1422 B.n375 B.n149 256.663
R1423 B.n373 B.n149 256.663
R1424 B.n367 B.n149 256.663
R1425 B.n365 B.n149 256.663
R1426 B.n359 B.n149 256.663
R1427 B.n357 B.n149 256.663
R1428 B.n351 B.n149 256.663
R1429 B.n349 B.n149 256.663
R1430 B.n342 B.n149 256.663
R1431 B.n340 B.n149 256.663
R1432 B.n334 B.n149 256.663
R1433 B.n332 B.n149 256.663
R1434 B.n326 B.n149 256.663
R1435 B.n188 B.n149 256.663
R1436 B.n320 B.n149 256.663
R1437 B.n314 B.n149 256.663
R1438 B.n312 B.n149 256.663
R1439 B.n306 B.n149 256.663
R1440 B.n304 B.n149 256.663
R1441 B.n298 B.n149 256.663
R1442 B.n296 B.n149 256.663
R1443 B.n290 B.n149 256.663
R1444 B.n288 B.n149 256.663
R1445 B.n282 B.n149 256.663
R1446 B.n280 B.n149 256.663
R1447 B.n274 B.n149 256.663
R1448 B.n272 B.n149 256.663
R1449 B.n266 B.n149 256.663
R1450 B.n264 B.n149 256.663
R1451 B.n258 B.n149 256.663
R1452 B.n256 B.n149 256.663
R1453 B.n250 B.n149 256.663
R1454 B.n248 B.n149 256.663
R1455 B.n242 B.n149 256.663
R1456 B.n240 B.n149 256.663
R1457 B.n234 B.n149 256.663
R1458 B.n232 B.n149 256.663
R1459 B.n226 B.n149 256.663
R1460 B.n224 B.n149 256.663
R1461 B.n218 B.n149 256.663
R1462 B.n216 B.n149 256.663
R1463 B.n457 B.n144 163.367
R1464 B.n465 B.n144 163.367
R1465 B.n465 B.n142 163.367
R1466 B.n469 B.n142 163.367
R1467 B.n469 B.n136 163.367
R1468 B.n477 B.n136 163.367
R1469 B.n477 B.n134 163.367
R1470 B.n481 B.n134 163.367
R1471 B.n481 B.n128 163.367
R1472 B.n490 B.n128 163.367
R1473 B.n490 B.n126 163.367
R1474 B.n494 B.n126 163.367
R1475 B.n494 B.n121 163.367
R1476 B.n503 B.n121 163.367
R1477 B.n503 B.n119 163.367
R1478 B.n507 B.n119 163.367
R1479 B.n507 B.n114 163.367
R1480 B.n516 B.n114 163.367
R1481 B.n516 B.n112 163.367
R1482 B.n520 B.n112 163.367
R1483 B.n520 B.n2 163.367
R1484 B.n841 B.n2 163.367
R1485 B.n841 B.n3 163.367
R1486 B.n837 B.n3 163.367
R1487 B.n837 B.n9 163.367
R1488 B.n833 B.n9 163.367
R1489 B.n833 B.n11 163.367
R1490 B.n829 B.n11 163.367
R1491 B.n829 B.n15 163.367
R1492 B.n825 B.n15 163.367
R1493 B.n825 B.n17 163.367
R1494 B.n821 B.n17 163.367
R1495 B.n821 B.n22 163.367
R1496 B.n817 B.n22 163.367
R1497 B.n817 B.n24 163.367
R1498 B.n813 B.n24 163.367
R1499 B.n813 B.n30 163.367
R1500 B.n809 B.n30 163.367
R1501 B.n809 B.n32 163.367
R1502 B.n805 B.n32 163.367
R1503 B.n805 B.n37 163.367
R1504 B.n801 B.n37 163.367
R1505 B.n801 B.n39 163.367
R1506 B.n797 B.n39 163.367
R1507 B.n453 B.n451 163.367
R1508 B.n451 B.n450 163.367
R1509 B.n447 B.n446 163.367
R1510 B.n444 B.n154 163.367
R1511 B.n440 B.n438 163.367
R1512 B.n436 B.n156 163.367
R1513 B.n432 B.n430 163.367
R1514 B.n428 B.n158 163.367
R1515 B.n424 B.n422 163.367
R1516 B.n420 B.n160 163.367
R1517 B.n416 B.n414 163.367
R1518 B.n412 B.n162 163.367
R1519 B.n408 B.n406 163.367
R1520 B.n404 B.n164 163.367
R1521 B.n400 B.n398 163.367
R1522 B.n396 B.n166 163.367
R1523 B.n392 B.n390 163.367
R1524 B.n388 B.n168 163.367
R1525 B.n384 B.n382 163.367
R1526 B.n380 B.n170 163.367
R1527 B.n376 B.n374 163.367
R1528 B.n372 B.n172 163.367
R1529 B.n368 B.n366 163.367
R1530 B.n364 B.n174 163.367
R1531 B.n360 B.n358 163.367
R1532 B.n356 B.n176 163.367
R1533 B.n352 B.n350 163.367
R1534 B.n348 B.n178 163.367
R1535 B.n343 B.n341 163.367
R1536 B.n339 B.n182 163.367
R1537 B.n335 B.n333 163.367
R1538 B.n331 B.n184 163.367
R1539 B.n327 B.n325 163.367
R1540 B.n322 B.n321 163.367
R1541 B.n319 B.n190 163.367
R1542 B.n315 B.n313 163.367
R1543 B.n311 B.n192 163.367
R1544 B.n307 B.n305 163.367
R1545 B.n303 B.n194 163.367
R1546 B.n299 B.n297 163.367
R1547 B.n295 B.n196 163.367
R1548 B.n291 B.n289 163.367
R1549 B.n287 B.n198 163.367
R1550 B.n283 B.n281 163.367
R1551 B.n279 B.n200 163.367
R1552 B.n275 B.n273 163.367
R1553 B.n271 B.n202 163.367
R1554 B.n267 B.n265 163.367
R1555 B.n263 B.n204 163.367
R1556 B.n259 B.n257 163.367
R1557 B.n255 B.n206 163.367
R1558 B.n251 B.n249 163.367
R1559 B.n247 B.n208 163.367
R1560 B.n243 B.n241 163.367
R1561 B.n239 B.n210 163.367
R1562 B.n235 B.n233 163.367
R1563 B.n231 B.n212 163.367
R1564 B.n227 B.n225 163.367
R1565 B.n223 B.n214 163.367
R1566 B.n219 B.n217 163.367
R1567 B.n459 B.n146 163.367
R1568 B.n463 B.n146 163.367
R1569 B.n463 B.n140 163.367
R1570 B.n471 B.n140 163.367
R1571 B.n471 B.n138 163.367
R1572 B.n475 B.n138 163.367
R1573 B.n475 B.n132 163.367
R1574 B.n483 B.n132 163.367
R1575 B.n483 B.n130 163.367
R1576 B.n487 B.n130 163.367
R1577 B.n487 B.n125 163.367
R1578 B.n496 B.n125 163.367
R1579 B.n496 B.n123 163.367
R1580 B.n500 B.n123 163.367
R1581 B.n500 B.n118 163.367
R1582 B.n509 B.n118 163.367
R1583 B.n509 B.n116 163.367
R1584 B.n514 B.n116 163.367
R1585 B.n514 B.n110 163.367
R1586 B.n522 B.n110 163.367
R1587 B.n523 B.n522 163.367
R1588 B.n523 B.n5 163.367
R1589 B.n6 B.n5 163.367
R1590 B.n7 B.n6 163.367
R1591 B.n528 B.n7 163.367
R1592 B.n528 B.n12 163.367
R1593 B.n13 B.n12 163.367
R1594 B.n14 B.n13 163.367
R1595 B.n533 B.n14 163.367
R1596 B.n533 B.n19 163.367
R1597 B.n20 B.n19 163.367
R1598 B.n21 B.n20 163.367
R1599 B.n538 B.n21 163.367
R1600 B.n538 B.n26 163.367
R1601 B.n27 B.n26 163.367
R1602 B.n28 B.n27 163.367
R1603 B.n543 B.n28 163.367
R1604 B.n543 B.n33 163.367
R1605 B.n34 B.n33 163.367
R1606 B.n35 B.n34 163.367
R1607 B.n548 B.n35 163.367
R1608 B.n548 B.n40 163.367
R1609 B.n41 B.n40 163.367
R1610 B.n42 B.n41 163.367
R1611 B.n793 B.n791 163.367
R1612 B.n789 B.n46 163.367
R1613 B.n785 B.n783 163.367
R1614 B.n781 B.n48 163.367
R1615 B.n777 B.n775 163.367
R1616 B.n773 B.n50 163.367
R1617 B.n769 B.n767 163.367
R1618 B.n765 B.n52 163.367
R1619 B.n761 B.n759 163.367
R1620 B.n757 B.n54 163.367
R1621 B.n753 B.n751 163.367
R1622 B.n749 B.n56 163.367
R1623 B.n745 B.n743 163.367
R1624 B.n741 B.n58 163.367
R1625 B.n737 B.n735 163.367
R1626 B.n733 B.n60 163.367
R1627 B.n729 B.n727 163.367
R1628 B.n725 B.n62 163.367
R1629 B.n721 B.n719 163.367
R1630 B.n717 B.n64 163.367
R1631 B.n713 B.n711 163.367
R1632 B.n709 B.n66 163.367
R1633 B.n705 B.n703 163.367
R1634 B.n701 B.n68 163.367
R1635 B.n697 B.n695 163.367
R1636 B.n693 B.n70 163.367
R1637 B.n689 B.n687 163.367
R1638 B.n685 B.n72 163.367
R1639 B.n680 B.n678 163.367
R1640 B.n676 B.n76 163.367
R1641 B.n672 B.n670 163.367
R1642 B.n668 B.n78 163.367
R1643 B.n663 B.n661 163.367
R1644 B.n659 B.n82 163.367
R1645 B.n655 B.n653 163.367
R1646 B.n651 B.n84 163.367
R1647 B.n647 B.n645 163.367
R1648 B.n643 B.n86 163.367
R1649 B.n639 B.n637 163.367
R1650 B.n635 B.n88 163.367
R1651 B.n631 B.n629 163.367
R1652 B.n627 B.n90 163.367
R1653 B.n623 B.n621 163.367
R1654 B.n619 B.n92 163.367
R1655 B.n615 B.n613 163.367
R1656 B.n611 B.n94 163.367
R1657 B.n607 B.n605 163.367
R1658 B.n603 B.n96 163.367
R1659 B.n599 B.n597 163.367
R1660 B.n595 B.n98 163.367
R1661 B.n591 B.n589 163.367
R1662 B.n587 B.n100 163.367
R1663 B.n583 B.n581 163.367
R1664 B.n579 B.n102 163.367
R1665 B.n575 B.n573 163.367
R1666 B.n571 B.n104 163.367
R1667 B.n567 B.n565 163.367
R1668 B.n563 B.n106 163.367
R1669 B.n559 B.n557 163.367
R1670 B.n555 B.n108 163.367
R1671 B.n452 B.n150 71.676
R1672 B.n450 B.n152 71.676
R1673 B.n446 B.n445 71.676
R1674 B.n439 B.n154 71.676
R1675 B.n438 B.n437 71.676
R1676 B.n431 B.n156 71.676
R1677 B.n430 B.n429 71.676
R1678 B.n423 B.n158 71.676
R1679 B.n422 B.n421 71.676
R1680 B.n415 B.n160 71.676
R1681 B.n414 B.n413 71.676
R1682 B.n407 B.n162 71.676
R1683 B.n406 B.n405 71.676
R1684 B.n399 B.n164 71.676
R1685 B.n398 B.n397 71.676
R1686 B.n391 B.n166 71.676
R1687 B.n390 B.n389 71.676
R1688 B.n383 B.n168 71.676
R1689 B.n382 B.n381 71.676
R1690 B.n375 B.n170 71.676
R1691 B.n374 B.n373 71.676
R1692 B.n367 B.n172 71.676
R1693 B.n366 B.n365 71.676
R1694 B.n359 B.n174 71.676
R1695 B.n358 B.n357 71.676
R1696 B.n351 B.n176 71.676
R1697 B.n350 B.n349 71.676
R1698 B.n342 B.n178 71.676
R1699 B.n341 B.n340 71.676
R1700 B.n334 B.n182 71.676
R1701 B.n333 B.n332 71.676
R1702 B.n326 B.n184 71.676
R1703 B.n325 B.n188 71.676
R1704 B.n321 B.n320 71.676
R1705 B.n314 B.n190 71.676
R1706 B.n313 B.n312 71.676
R1707 B.n306 B.n192 71.676
R1708 B.n305 B.n304 71.676
R1709 B.n298 B.n194 71.676
R1710 B.n297 B.n296 71.676
R1711 B.n290 B.n196 71.676
R1712 B.n289 B.n288 71.676
R1713 B.n282 B.n198 71.676
R1714 B.n281 B.n280 71.676
R1715 B.n274 B.n200 71.676
R1716 B.n273 B.n272 71.676
R1717 B.n266 B.n202 71.676
R1718 B.n265 B.n264 71.676
R1719 B.n258 B.n204 71.676
R1720 B.n257 B.n256 71.676
R1721 B.n250 B.n206 71.676
R1722 B.n249 B.n248 71.676
R1723 B.n242 B.n208 71.676
R1724 B.n241 B.n240 71.676
R1725 B.n234 B.n210 71.676
R1726 B.n233 B.n232 71.676
R1727 B.n226 B.n212 71.676
R1728 B.n225 B.n224 71.676
R1729 B.n218 B.n214 71.676
R1730 B.n217 B.n216 71.676
R1731 B.n792 B.n44 71.676
R1732 B.n791 B.n790 71.676
R1733 B.n784 B.n46 71.676
R1734 B.n783 B.n782 71.676
R1735 B.n776 B.n48 71.676
R1736 B.n775 B.n774 71.676
R1737 B.n768 B.n50 71.676
R1738 B.n767 B.n766 71.676
R1739 B.n760 B.n52 71.676
R1740 B.n759 B.n758 71.676
R1741 B.n752 B.n54 71.676
R1742 B.n751 B.n750 71.676
R1743 B.n744 B.n56 71.676
R1744 B.n743 B.n742 71.676
R1745 B.n736 B.n58 71.676
R1746 B.n735 B.n734 71.676
R1747 B.n728 B.n60 71.676
R1748 B.n727 B.n726 71.676
R1749 B.n720 B.n62 71.676
R1750 B.n719 B.n718 71.676
R1751 B.n712 B.n64 71.676
R1752 B.n711 B.n710 71.676
R1753 B.n704 B.n66 71.676
R1754 B.n703 B.n702 71.676
R1755 B.n696 B.n68 71.676
R1756 B.n695 B.n694 71.676
R1757 B.n688 B.n70 71.676
R1758 B.n687 B.n686 71.676
R1759 B.n679 B.n72 71.676
R1760 B.n678 B.n677 71.676
R1761 B.n671 B.n76 71.676
R1762 B.n670 B.n669 71.676
R1763 B.n662 B.n78 71.676
R1764 B.n661 B.n660 71.676
R1765 B.n654 B.n82 71.676
R1766 B.n653 B.n652 71.676
R1767 B.n646 B.n84 71.676
R1768 B.n645 B.n644 71.676
R1769 B.n638 B.n86 71.676
R1770 B.n637 B.n636 71.676
R1771 B.n630 B.n88 71.676
R1772 B.n629 B.n628 71.676
R1773 B.n622 B.n90 71.676
R1774 B.n621 B.n620 71.676
R1775 B.n614 B.n92 71.676
R1776 B.n613 B.n612 71.676
R1777 B.n606 B.n94 71.676
R1778 B.n605 B.n604 71.676
R1779 B.n598 B.n96 71.676
R1780 B.n597 B.n596 71.676
R1781 B.n590 B.n98 71.676
R1782 B.n589 B.n588 71.676
R1783 B.n582 B.n100 71.676
R1784 B.n581 B.n580 71.676
R1785 B.n574 B.n102 71.676
R1786 B.n573 B.n572 71.676
R1787 B.n566 B.n104 71.676
R1788 B.n565 B.n564 71.676
R1789 B.n558 B.n106 71.676
R1790 B.n557 B.n556 71.676
R1791 B.n556 B.n555 71.676
R1792 B.n559 B.n558 71.676
R1793 B.n564 B.n563 71.676
R1794 B.n567 B.n566 71.676
R1795 B.n572 B.n571 71.676
R1796 B.n575 B.n574 71.676
R1797 B.n580 B.n579 71.676
R1798 B.n583 B.n582 71.676
R1799 B.n588 B.n587 71.676
R1800 B.n591 B.n590 71.676
R1801 B.n596 B.n595 71.676
R1802 B.n599 B.n598 71.676
R1803 B.n604 B.n603 71.676
R1804 B.n607 B.n606 71.676
R1805 B.n612 B.n611 71.676
R1806 B.n615 B.n614 71.676
R1807 B.n620 B.n619 71.676
R1808 B.n623 B.n622 71.676
R1809 B.n628 B.n627 71.676
R1810 B.n631 B.n630 71.676
R1811 B.n636 B.n635 71.676
R1812 B.n639 B.n638 71.676
R1813 B.n644 B.n643 71.676
R1814 B.n647 B.n646 71.676
R1815 B.n652 B.n651 71.676
R1816 B.n655 B.n654 71.676
R1817 B.n660 B.n659 71.676
R1818 B.n663 B.n662 71.676
R1819 B.n669 B.n668 71.676
R1820 B.n672 B.n671 71.676
R1821 B.n677 B.n676 71.676
R1822 B.n680 B.n679 71.676
R1823 B.n686 B.n685 71.676
R1824 B.n689 B.n688 71.676
R1825 B.n694 B.n693 71.676
R1826 B.n697 B.n696 71.676
R1827 B.n702 B.n701 71.676
R1828 B.n705 B.n704 71.676
R1829 B.n710 B.n709 71.676
R1830 B.n713 B.n712 71.676
R1831 B.n718 B.n717 71.676
R1832 B.n721 B.n720 71.676
R1833 B.n726 B.n725 71.676
R1834 B.n729 B.n728 71.676
R1835 B.n734 B.n733 71.676
R1836 B.n737 B.n736 71.676
R1837 B.n742 B.n741 71.676
R1838 B.n745 B.n744 71.676
R1839 B.n750 B.n749 71.676
R1840 B.n753 B.n752 71.676
R1841 B.n758 B.n757 71.676
R1842 B.n761 B.n760 71.676
R1843 B.n766 B.n765 71.676
R1844 B.n769 B.n768 71.676
R1845 B.n774 B.n773 71.676
R1846 B.n777 B.n776 71.676
R1847 B.n782 B.n781 71.676
R1848 B.n785 B.n784 71.676
R1849 B.n790 B.n789 71.676
R1850 B.n793 B.n792 71.676
R1851 B.n453 B.n452 71.676
R1852 B.n447 B.n152 71.676
R1853 B.n445 B.n444 71.676
R1854 B.n440 B.n439 71.676
R1855 B.n437 B.n436 71.676
R1856 B.n432 B.n431 71.676
R1857 B.n429 B.n428 71.676
R1858 B.n424 B.n423 71.676
R1859 B.n421 B.n420 71.676
R1860 B.n416 B.n415 71.676
R1861 B.n413 B.n412 71.676
R1862 B.n408 B.n407 71.676
R1863 B.n405 B.n404 71.676
R1864 B.n400 B.n399 71.676
R1865 B.n397 B.n396 71.676
R1866 B.n392 B.n391 71.676
R1867 B.n389 B.n388 71.676
R1868 B.n384 B.n383 71.676
R1869 B.n381 B.n380 71.676
R1870 B.n376 B.n375 71.676
R1871 B.n373 B.n372 71.676
R1872 B.n368 B.n367 71.676
R1873 B.n365 B.n364 71.676
R1874 B.n360 B.n359 71.676
R1875 B.n357 B.n356 71.676
R1876 B.n352 B.n351 71.676
R1877 B.n349 B.n348 71.676
R1878 B.n343 B.n342 71.676
R1879 B.n340 B.n339 71.676
R1880 B.n335 B.n334 71.676
R1881 B.n332 B.n331 71.676
R1882 B.n327 B.n326 71.676
R1883 B.n322 B.n188 71.676
R1884 B.n320 B.n319 71.676
R1885 B.n315 B.n314 71.676
R1886 B.n312 B.n311 71.676
R1887 B.n307 B.n306 71.676
R1888 B.n304 B.n303 71.676
R1889 B.n299 B.n298 71.676
R1890 B.n296 B.n295 71.676
R1891 B.n291 B.n290 71.676
R1892 B.n288 B.n287 71.676
R1893 B.n283 B.n282 71.676
R1894 B.n280 B.n279 71.676
R1895 B.n275 B.n274 71.676
R1896 B.n272 B.n271 71.676
R1897 B.n267 B.n266 71.676
R1898 B.n264 B.n263 71.676
R1899 B.n259 B.n258 71.676
R1900 B.n256 B.n255 71.676
R1901 B.n251 B.n250 71.676
R1902 B.n248 B.n247 71.676
R1903 B.n243 B.n242 71.676
R1904 B.n240 B.n239 71.676
R1905 B.n235 B.n234 71.676
R1906 B.n232 B.n231 71.676
R1907 B.n227 B.n226 71.676
R1908 B.n224 B.n223 71.676
R1909 B.n219 B.n218 71.676
R1910 B.n216 B.n148 71.676
R1911 B.n458 B.n149 69.1704
R1912 B.n798 B.n43 69.1704
R1913 B.n187 B.n186 59.5399
R1914 B.n345 B.n180 59.5399
R1915 B.n683 B.n74 59.5399
R1916 B.n665 B.n80 59.5399
R1917 B.n553 B.n552 36.059
R1918 B.n796 B.n795 36.059
R1919 B.n460 B.n147 36.059
R1920 B.n456 B.n455 36.059
R1921 B.n458 B.n145 33.839
R1922 B.n464 B.n145 33.839
R1923 B.n464 B.n141 33.839
R1924 B.n470 B.n141 33.839
R1925 B.n476 B.n137 33.839
R1926 B.n476 B.n133 33.839
R1927 B.n482 B.n133 33.839
R1928 B.n482 B.n129 33.839
R1929 B.n489 B.n129 33.839
R1930 B.n489 B.n488 33.839
R1931 B.n495 B.n122 33.839
R1932 B.n502 B.n122 33.839
R1933 B.n502 B.n501 33.839
R1934 B.n508 B.n115 33.839
R1935 B.n515 B.n115 33.839
R1936 B.n521 B.n111 33.839
R1937 B.n521 B.n4 33.839
R1938 B.n840 B.n4 33.839
R1939 B.n840 B.n839 33.839
R1940 B.n839 B.n838 33.839
R1941 B.n838 B.n8 33.839
R1942 B.n832 B.n831 33.839
R1943 B.n831 B.n830 33.839
R1944 B.n824 B.n18 33.839
R1945 B.n824 B.n823 33.839
R1946 B.n823 B.n822 33.839
R1947 B.n816 B.n25 33.839
R1948 B.n816 B.n815 33.839
R1949 B.n815 B.n814 33.839
R1950 B.n814 B.n29 33.839
R1951 B.n808 B.n29 33.839
R1952 B.n808 B.n807 33.839
R1953 B.n806 B.n36 33.839
R1954 B.n800 B.n36 33.839
R1955 B.n800 B.n799 33.839
R1956 B.n799 B.n798 33.839
R1957 B.n508 B.t3 30.3556
R1958 B.n830 B.t5 30.3556
R1959 B.n470 B.t11 28.3651
R1960 B.t7 B.n806 28.3651
R1961 B.n186 B.n185 23.2732
R1962 B.n180 B.n179 23.2732
R1963 B.n74 B.n73 23.2732
R1964 B.n80 B.n79 23.2732
R1965 B.n515 B.t4 21.3984
R1966 B.n832 B.t1 21.3984
R1967 B.n488 B.t2 19.4079
R1968 B.n25 B.t0 19.4079
R1969 B B.n842 18.0485
R1970 B.n495 B.t2 14.4316
R1971 B.n822 B.t0 14.4316
R1972 B.t4 B.n111 12.4411
R1973 B.t1 B.n8 12.4411
R1974 B.n795 B.n794 10.6151
R1975 B.n794 B.n45 10.6151
R1976 B.n788 B.n45 10.6151
R1977 B.n788 B.n787 10.6151
R1978 B.n787 B.n786 10.6151
R1979 B.n786 B.n47 10.6151
R1980 B.n780 B.n47 10.6151
R1981 B.n780 B.n779 10.6151
R1982 B.n779 B.n778 10.6151
R1983 B.n778 B.n49 10.6151
R1984 B.n772 B.n49 10.6151
R1985 B.n772 B.n771 10.6151
R1986 B.n771 B.n770 10.6151
R1987 B.n770 B.n51 10.6151
R1988 B.n764 B.n51 10.6151
R1989 B.n764 B.n763 10.6151
R1990 B.n763 B.n762 10.6151
R1991 B.n762 B.n53 10.6151
R1992 B.n756 B.n53 10.6151
R1993 B.n756 B.n755 10.6151
R1994 B.n755 B.n754 10.6151
R1995 B.n754 B.n55 10.6151
R1996 B.n748 B.n55 10.6151
R1997 B.n748 B.n747 10.6151
R1998 B.n747 B.n746 10.6151
R1999 B.n746 B.n57 10.6151
R2000 B.n740 B.n57 10.6151
R2001 B.n740 B.n739 10.6151
R2002 B.n739 B.n738 10.6151
R2003 B.n738 B.n59 10.6151
R2004 B.n732 B.n59 10.6151
R2005 B.n732 B.n731 10.6151
R2006 B.n731 B.n730 10.6151
R2007 B.n730 B.n61 10.6151
R2008 B.n724 B.n61 10.6151
R2009 B.n724 B.n723 10.6151
R2010 B.n723 B.n722 10.6151
R2011 B.n722 B.n63 10.6151
R2012 B.n716 B.n63 10.6151
R2013 B.n716 B.n715 10.6151
R2014 B.n715 B.n714 10.6151
R2015 B.n714 B.n65 10.6151
R2016 B.n708 B.n65 10.6151
R2017 B.n708 B.n707 10.6151
R2018 B.n707 B.n706 10.6151
R2019 B.n706 B.n67 10.6151
R2020 B.n700 B.n67 10.6151
R2021 B.n700 B.n699 10.6151
R2022 B.n699 B.n698 10.6151
R2023 B.n698 B.n69 10.6151
R2024 B.n692 B.n69 10.6151
R2025 B.n692 B.n691 10.6151
R2026 B.n691 B.n690 10.6151
R2027 B.n690 B.n71 10.6151
R2028 B.n684 B.n71 10.6151
R2029 B.n682 B.n681 10.6151
R2030 B.n681 B.n75 10.6151
R2031 B.n675 B.n75 10.6151
R2032 B.n675 B.n674 10.6151
R2033 B.n674 B.n673 10.6151
R2034 B.n673 B.n77 10.6151
R2035 B.n667 B.n77 10.6151
R2036 B.n667 B.n666 10.6151
R2037 B.n664 B.n81 10.6151
R2038 B.n658 B.n81 10.6151
R2039 B.n658 B.n657 10.6151
R2040 B.n657 B.n656 10.6151
R2041 B.n656 B.n83 10.6151
R2042 B.n650 B.n83 10.6151
R2043 B.n650 B.n649 10.6151
R2044 B.n649 B.n648 10.6151
R2045 B.n648 B.n85 10.6151
R2046 B.n642 B.n85 10.6151
R2047 B.n642 B.n641 10.6151
R2048 B.n641 B.n640 10.6151
R2049 B.n640 B.n87 10.6151
R2050 B.n634 B.n87 10.6151
R2051 B.n634 B.n633 10.6151
R2052 B.n633 B.n632 10.6151
R2053 B.n632 B.n89 10.6151
R2054 B.n626 B.n89 10.6151
R2055 B.n626 B.n625 10.6151
R2056 B.n625 B.n624 10.6151
R2057 B.n624 B.n91 10.6151
R2058 B.n618 B.n91 10.6151
R2059 B.n618 B.n617 10.6151
R2060 B.n617 B.n616 10.6151
R2061 B.n616 B.n93 10.6151
R2062 B.n610 B.n93 10.6151
R2063 B.n610 B.n609 10.6151
R2064 B.n609 B.n608 10.6151
R2065 B.n608 B.n95 10.6151
R2066 B.n602 B.n95 10.6151
R2067 B.n602 B.n601 10.6151
R2068 B.n601 B.n600 10.6151
R2069 B.n600 B.n97 10.6151
R2070 B.n594 B.n97 10.6151
R2071 B.n594 B.n593 10.6151
R2072 B.n593 B.n592 10.6151
R2073 B.n592 B.n99 10.6151
R2074 B.n586 B.n99 10.6151
R2075 B.n586 B.n585 10.6151
R2076 B.n585 B.n584 10.6151
R2077 B.n584 B.n101 10.6151
R2078 B.n578 B.n101 10.6151
R2079 B.n578 B.n577 10.6151
R2080 B.n577 B.n576 10.6151
R2081 B.n576 B.n103 10.6151
R2082 B.n570 B.n103 10.6151
R2083 B.n570 B.n569 10.6151
R2084 B.n569 B.n568 10.6151
R2085 B.n568 B.n105 10.6151
R2086 B.n562 B.n105 10.6151
R2087 B.n562 B.n561 10.6151
R2088 B.n561 B.n560 10.6151
R2089 B.n560 B.n107 10.6151
R2090 B.n554 B.n107 10.6151
R2091 B.n554 B.n553 10.6151
R2092 B.n461 B.n460 10.6151
R2093 B.n462 B.n461 10.6151
R2094 B.n462 B.n139 10.6151
R2095 B.n472 B.n139 10.6151
R2096 B.n473 B.n472 10.6151
R2097 B.n474 B.n473 10.6151
R2098 B.n474 B.n131 10.6151
R2099 B.n484 B.n131 10.6151
R2100 B.n485 B.n484 10.6151
R2101 B.n486 B.n485 10.6151
R2102 B.n486 B.n124 10.6151
R2103 B.n497 B.n124 10.6151
R2104 B.n498 B.n497 10.6151
R2105 B.n499 B.n498 10.6151
R2106 B.n499 B.n117 10.6151
R2107 B.n510 B.n117 10.6151
R2108 B.n511 B.n510 10.6151
R2109 B.n513 B.n511 10.6151
R2110 B.n513 B.n512 10.6151
R2111 B.n512 B.n109 10.6151
R2112 B.n524 B.n109 10.6151
R2113 B.n525 B.n524 10.6151
R2114 B.n526 B.n525 10.6151
R2115 B.n527 B.n526 10.6151
R2116 B.n529 B.n527 10.6151
R2117 B.n530 B.n529 10.6151
R2118 B.n531 B.n530 10.6151
R2119 B.n532 B.n531 10.6151
R2120 B.n534 B.n532 10.6151
R2121 B.n535 B.n534 10.6151
R2122 B.n536 B.n535 10.6151
R2123 B.n537 B.n536 10.6151
R2124 B.n539 B.n537 10.6151
R2125 B.n540 B.n539 10.6151
R2126 B.n541 B.n540 10.6151
R2127 B.n542 B.n541 10.6151
R2128 B.n544 B.n542 10.6151
R2129 B.n545 B.n544 10.6151
R2130 B.n546 B.n545 10.6151
R2131 B.n547 B.n546 10.6151
R2132 B.n549 B.n547 10.6151
R2133 B.n550 B.n549 10.6151
R2134 B.n551 B.n550 10.6151
R2135 B.n552 B.n551 10.6151
R2136 B.n455 B.n454 10.6151
R2137 B.n454 B.n151 10.6151
R2138 B.n449 B.n151 10.6151
R2139 B.n449 B.n448 10.6151
R2140 B.n448 B.n153 10.6151
R2141 B.n443 B.n153 10.6151
R2142 B.n443 B.n442 10.6151
R2143 B.n442 B.n441 10.6151
R2144 B.n441 B.n155 10.6151
R2145 B.n435 B.n155 10.6151
R2146 B.n435 B.n434 10.6151
R2147 B.n434 B.n433 10.6151
R2148 B.n433 B.n157 10.6151
R2149 B.n427 B.n157 10.6151
R2150 B.n427 B.n426 10.6151
R2151 B.n426 B.n425 10.6151
R2152 B.n425 B.n159 10.6151
R2153 B.n419 B.n159 10.6151
R2154 B.n419 B.n418 10.6151
R2155 B.n418 B.n417 10.6151
R2156 B.n417 B.n161 10.6151
R2157 B.n411 B.n161 10.6151
R2158 B.n411 B.n410 10.6151
R2159 B.n410 B.n409 10.6151
R2160 B.n409 B.n163 10.6151
R2161 B.n403 B.n163 10.6151
R2162 B.n403 B.n402 10.6151
R2163 B.n402 B.n401 10.6151
R2164 B.n401 B.n165 10.6151
R2165 B.n395 B.n165 10.6151
R2166 B.n395 B.n394 10.6151
R2167 B.n394 B.n393 10.6151
R2168 B.n393 B.n167 10.6151
R2169 B.n387 B.n167 10.6151
R2170 B.n387 B.n386 10.6151
R2171 B.n386 B.n385 10.6151
R2172 B.n385 B.n169 10.6151
R2173 B.n379 B.n169 10.6151
R2174 B.n379 B.n378 10.6151
R2175 B.n378 B.n377 10.6151
R2176 B.n377 B.n171 10.6151
R2177 B.n371 B.n171 10.6151
R2178 B.n371 B.n370 10.6151
R2179 B.n370 B.n369 10.6151
R2180 B.n369 B.n173 10.6151
R2181 B.n363 B.n173 10.6151
R2182 B.n363 B.n362 10.6151
R2183 B.n362 B.n361 10.6151
R2184 B.n361 B.n175 10.6151
R2185 B.n355 B.n175 10.6151
R2186 B.n355 B.n354 10.6151
R2187 B.n354 B.n353 10.6151
R2188 B.n353 B.n177 10.6151
R2189 B.n347 B.n177 10.6151
R2190 B.n347 B.n346 10.6151
R2191 B.n344 B.n181 10.6151
R2192 B.n338 B.n181 10.6151
R2193 B.n338 B.n337 10.6151
R2194 B.n337 B.n336 10.6151
R2195 B.n336 B.n183 10.6151
R2196 B.n330 B.n183 10.6151
R2197 B.n330 B.n329 10.6151
R2198 B.n329 B.n328 10.6151
R2199 B.n324 B.n323 10.6151
R2200 B.n323 B.n189 10.6151
R2201 B.n318 B.n189 10.6151
R2202 B.n318 B.n317 10.6151
R2203 B.n317 B.n316 10.6151
R2204 B.n316 B.n191 10.6151
R2205 B.n310 B.n191 10.6151
R2206 B.n310 B.n309 10.6151
R2207 B.n309 B.n308 10.6151
R2208 B.n308 B.n193 10.6151
R2209 B.n302 B.n193 10.6151
R2210 B.n302 B.n301 10.6151
R2211 B.n301 B.n300 10.6151
R2212 B.n300 B.n195 10.6151
R2213 B.n294 B.n195 10.6151
R2214 B.n294 B.n293 10.6151
R2215 B.n293 B.n292 10.6151
R2216 B.n292 B.n197 10.6151
R2217 B.n286 B.n197 10.6151
R2218 B.n286 B.n285 10.6151
R2219 B.n285 B.n284 10.6151
R2220 B.n284 B.n199 10.6151
R2221 B.n278 B.n199 10.6151
R2222 B.n278 B.n277 10.6151
R2223 B.n277 B.n276 10.6151
R2224 B.n276 B.n201 10.6151
R2225 B.n270 B.n201 10.6151
R2226 B.n270 B.n269 10.6151
R2227 B.n269 B.n268 10.6151
R2228 B.n268 B.n203 10.6151
R2229 B.n262 B.n203 10.6151
R2230 B.n262 B.n261 10.6151
R2231 B.n261 B.n260 10.6151
R2232 B.n260 B.n205 10.6151
R2233 B.n254 B.n205 10.6151
R2234 B.n254 B.n253 10.6151
R2235 B.n253 B.n252 10.6151
R2236 B.n252 B.n207 10.6151
R2237 B.n246 B.n207 10.6151
R2238 B.n246 B.n245 10.6151
R2239 B.n245 B.n244 10.6151
R2240 B.n244 B.n209 10.6151
R2241 B.n238 B.n209 10.6151
R2242 B.n238 B.n237 10.6151
R2243 B.n237 B.n236 10.6151
R2244 B.n236 B.n211 10.6151
R2245 B.n230 B.n211 10.6151
R2246 B.n230 B.n229 10.6151
R2247 B.n229 B.n228 10.6151
R2248 B.n228 B.n213 10.6151
R2249 B.n222 B.n213 10.6151
R2250 B.n222 B.n221 10.6151
R2251 B.n221 B.n220 10.6151
R2252 B.n220 B.n215 10.6151
R2253 B.n215 B.n147 10.6151
R2254 B.n456 B.n143 10.6151
R2255 B.n466 B.n143 10.6151
R2256 B.n467 B.n466 10.6151
R2257 B.n468 B.n467 10.6151
R2258 B.n468 B.n135 10.6151
R2259 B.n478 B.n135 10.6151
R2260 B.n479 B.n478 10.6151
R2261 B.n480 B.n479 10.6151
R2262 B.n480 B.n127 10.6151
R2263 B.n491 B.n127 10.6151
R2264 B.n492 B.n491 10.6151
R2265 B.n493 B.n492 10.6151
R2266 B.n493 B.n120 10.6151
R2267 B.n504 B.n120 10.6151
R2268 B.n505 B.n504 10.6151
R2269 B.n506 B.n505 10.6151
R2270 B.n506 B.n113 10.6151
R2271 B.n517 B.n113 10.6151
R2272 B.n518 B.n517 10.6151
R2273 B.n519 B.n518 10.6151
R2274 B.n519 B.n0 10.6151
R2275 B.n836 B.n1 10.6151
R2276 B.n836 B.n835 10.6151
R2277 B.n835 B.n834 10.6151
R2278 B.n834 B.n10 10.6151
R2279 B.n828 B.n10 10.6151
R2280 B.n828 B.n827 10.6151
R2281 B.n827 B.n826 10.6151
R2282 B.n826 B.n16 10.6151
R2283 B.n820 B.n16 10.6151
R2284 B.n820 B.n819 10.6151
R2285 B.n819 B.n818 10.6151
R2286 B.n818 B.n23 10.6151
R2287 B.n812 B.n23 10.6151
R2288 B.n812 B.n811 10.6151
R2289 B.n811 B.n810 10.6151
R2290 B.n810 B.n31 10.6151
R2291 B.n804 B.n31 10.6151
R2292 B.n804 B.n803 10.6151
R2293 B.n803 B.n802 10.6151
R2294 B.n802 B.n38 10.6151
R2295 B.n796 B.n38 10.6151
R2296 B.n683 B.n682 6.5566
R2297 B.n666 B.n665 6.5566
R2298 B.n345 B.n344 6.5566
R2299 B.n328 B.n187 6.5566
R2300 B.t11 B.n137 5.47437
R2301 B.n807 B.t7 5.47437
R2302 B.n684 B.n683 4.05904
R2303 B.n665 B.n664 4.05904
R2304 B.n346 B.n345 4.05904
R2305 B.n324 B.n187 4.05904
R2306 B.n501 B.t3 3.48387
R2307 B.n18 B.t5 3.48387
R2308 B.n842 B.n0 2.81026
R2309 B.n842 B.n1 2.81026
R2310 VP.n5 VP.t2 527.88
R2311 VP.n12 VP.t4 511.64
R2312 VP.n19 VP.t3 511.64
R2313 VP.n9 VP.t0 511.64
R2314 VP.n1 VP.t1 466.211
R2315 VP.n4 VP.t5 466.211
R2316 VP.n20 VP.n19 161.3
R2317 VP.n7 VP.n6 161.3
R2318 VP.n8 VP.n3 161.3
R2319 VP.n10 VP.n9 161.3
R2320 VP.n18 VP.n0 161.3
R2321 VP.n17 VP.n16 161.3
R2322 VP.n15 VP.n14 161.3
R2323 VP.n13 VP.n2 161.3
R2324 VP.n12 VP.n11 161.3
R2325 VP.n14 VP.n13 55.0624
R2326 VP.n18 VP.n17 55.0624
R2327 VP.n8 VP.n7 55.0624
R2328 VP.n11 VP.n10 45.5081
R2329 VP.n6 VP.n5 43.7084
R2330 VP.n5 VP.n4 42.6481
R2331 VP.n14 VP.n1 12.234
R2332 VP.n17 VP.n1 12.234
R2333 VP.n7 VP.n4 12.234
R2334 VP.n13 VP.n12 2.19141
R2335 VP.n19 VP.n18 2.19141
R2336 VP.n9 VP.n8 2.19141
R2337 VP.n6 VP.n3 0.189894
R2338 VP.n10 VP.n3 0.189894
R2339 VP.n11 VP.n2 0.189894
R2340 VP.n15 VP.n2 0.189894
R2341 VP.n16 VP.n15 0.189894
R2342 VP.n16 VP.n0 0.189894
R2343 VP.n20 VP.n0 0.189894
R2344 VP VP.n20 0.0516364
R2345 VDD1.n88 VDD1.n0 289.615
R2346 VDD1.n181 VDD1.n93 289.615
R2347 VDD1.n89 VDD1.n88 185
R2348 VDD1.n87 VDD1.n86 185
R2349 VDD1.n4 VDD1.n3 185
R2350 VDD1.n81 VDD1.n80 185
R2351 VDD1.n79 VDD1.n78 185
R2352 VDD1.n77 VDD1.n7 185
R2353 VDD1.n11 VDD1.n8 185
R2354 VDD1.n72 VDD1.n71 185
R2355 VDD1.n70 VDD1.n69 185
R2356 VDD1.n13 VDD1.n12 185
R2357 VDD1.n64 VDD1.n63 185
R2358 VDD1.n62 VDD1.n61 185
R2359 VDD1.n17 VDD1.n16 185
R2360 VDD1.n56 VDD1.n55 185
R2361 VDD1.n54 VDD1.n53 185
R2362 VDD1.n21 VDD1.n20 185
R2363 VDD1.n48 VDD1.n47 185
R2364 VDD1.n46 VDD1.n45 185
R2365 VDD1.n25 VDD1.n24 185
R2366 VDD1.n40 VDD1.n39 185
R2367 VDD1.n38 VDD1.n37 185
R2368 VDD1.n29 VDD1.n28 185
R2369 VDD1.n32 VDD1.n31 185
R2370 VDD1.n124 VDD1.n123 185
R2371 VDD1.n121 VDD1.n120 185
R2372 VDD1.n130 VDD1.n129 185
R2373 VDD1.n132 VDD1.n131 185
R2374 VDD1.n117 VDD1.n116 185
R2375 VDD1.n138 VDD1.n137 185
R2376 VDD1.n140 VDD1.n139 185
R2377 VDD1.n113 VDD1.n112 185
R2378 VDD1.n146 VDD1.n145 185
R2379 VDD1.n148 VDD1.n147 185
R2380 VDD1.n109 VDD1.n108 185
R2381 VDD1.n154 VDD1.n153 185
R2382 VDD1.n156 VDD1.n155 185
R2383 VDD1.n105 VDD1.n104 185
R2384 VDD1.n162 VDD1.n161 185
R2385 VDD1.n165 VDD1.n164 185
R2386 VDD1.n163 VDD1.n101 185
R2387 VDD1.n170 VDD1.n100 185
R2388 VDD1.n172 VDD1.n171 185
R2389 VDD1.n174 VDD1.n173 185
R2390 VDD1.n97 VDD1.n96 185
R2391 VDD1.n180 VDD1.n179 185
R2392 VDD1.n182 VDD1.n181 185
R2393 VDD1.t3 VDD1.n30 147.659
R2394 VDD1.t1 VDD1.n122 147.659
R2395 VDD1.n88 VDD1.n87 104.615
R2396 VDD1.n87 VDD1.n3 104.615
R2397 VDD1.n80 VDD1.n3 104.615
R2398 VDD1.n80 VDD1.n79 104.615
R2399 VDD1.n79 VDD1.n7 104.615
R2400 VDD1.n11 VDD1.n7 104.615
R2401 VDD1.n71 VDD1.n11 104.615
R2402 VDD1.n71 VDD1.n70 104.615
R2403 VDD1.n70 VDD1.n12 104.615
R2404 VDD1.n63 VDD1.n12 104.615
R2405 VDD1.n63 VDD1.n62 104.615
R2406 VDD1.n62 VDD1.n16 104.615
R2407 VDD1.n55 VDD1.n16 104.615
R2408 VDD1.n55 VDD1.n54 104.615
R2409 VDD1.n54 VDD1.n20 104.615
R2410 VDD1.n47 VDD1.n20 104.615
R2411 VDD1.n47 VDD1.n46 104.615
R2412 VDD1.n46 VDD1.n24 104.615
R2413 VDD1.n39 VDD1.n24 104.615
R2414 VDD1.n39 VDD1.n38 104.615
R2415 VDD1.n38 VDD1.n28 104.615
R2416 VDD1.n31 VDD1.n28 104.615
R2417 VDD1.n123 VDD1.n120 104.615
R2418 VDD1.n130 VDD1.n120 104.615
R2419 VDD1.n131 VDD1.n130 104.615
R2420 VDD1.n131 VDD1.n116 104.615
R2421 VDD1.n138 VDD1.n116 104.615
R2422 VDD1.n139 VDD1.n138 104.615
R2423 VDD1.n139 VDD1.n112 104.615
R2424 VDD1.n146 VDD1.n112 104.615
R2425 VDD1.n147 VDD1.n146 104.615
R2426 VDD1.n147 VDD1.n108 104.615
R2427 VDD1.n154 VDD1.n108 104.615
R2428 VDD1.n155 VDD1.n154 104.615
R2429 VDD1.n155 VDD1.n104 104.615
R2430 VDD1.n162 VDD1.n104 104.615
R2431 VDD1.n164 VDD1.n162 104.615
R2432 VDD1.n164 VDD1.n163 104.615
R2433 VDD1.n163 VDD1.n100 104.615
R2434 VDD1.n172 VDD1.n100 104.615
R2435 VDD1.n173 VDD1.n172 104.615
R2436 VDD1.n173 VDD1.n96 104.615
R2437 VDD1.n180 VDD1.n96 104.615
R2438 VDD1.n181 VDD1.n180 104.615
R2439 VDD1.n187 VDD1.n186 61.5097
R2440 VDD1.n189 VDD1.n188 61.3065
R2441 VDD1.n31 VDD1.t3 52.3082
R2442 VDD1.n123 VDD1.t1 52.3082
R2443 VDD1 VDD1.n92 50.28
R2444 VDD1.n187 VDD1.n185 50.1665
R2445 VDD1.n189 VDD1.n187 42.6862
R2446 VDD1.n32 VDD1.n30 15.6677
R2447 VDD1.n124 VDD1.n122 15.6677
R2448 VDD1.n78 VDD1.n77 13.1884
R2449 VDD1.n171 VDD1.n170 13.1884
R2450 VDD1.n81 VDD1.n6 12.8005
R2451 VDD1.n76 VDD1.n8 12.8005
R2452 VDD1.n33 VDD1.n29 12.8005
R2453 VDD1.n125 VDD1.n121 12.8005
R2454 VDD1.n169 VDD1.n101 12.8005
R2455 VDD1.n174 VDD1.n99 12.8005
R2456 VDD1.n82 VDD1.n4 12.0247
R2457 VDD1.n73 VDD1.n72 12.0247
R2458 VDD1.n37 VDD1.n36 12.0247
R2459 VDD1.n129 VDD1.n128 12.0247
R2460 VDD1.n166 VDD1.n165 12.0247
R2461 VDD1.n175 VDD1.n97 12.0247
R2462 VDD1.n86 VDD1.n85 11.249
R2463 VDD1.n69 VDD1.n10 11.249
R2464 VDD1.n40 VDD1.n27 11.249
R2465 VDD1.n132 VDD1.n119 11.249
R2466 VDD1.n161 VDD1.n103 11.249
R2467 VDD1.n179 VDD1.n178 11.249
R2468 VDD1.n89 VDD1.n2 10.4732
R2469 VDD1.n68 VDD1.n13 10.4732
R2470 VDD1.n41 VDD1.n25 10.4732
R2471 VDD1.n133 VDD1.n117 10.4732
R2472 VDD1.n160 VDD1.n105 10.4732
R2473 VDD1.n182 VDD1.n95 10.4732
R2474 VDD1.n90 VDD1.n0 9.69747
R2475 VDD1.n65 VDD1.n64 9.69747
R2476 VDD1.n45 VDD1.n44 9.69747
R2477 VDD1.n137 VDD1.n136 9.69747
R2478 VDD1.n157 VDD1.n156 9.69747
R2479 VDD1.n183 VDD1.n93 9.69747
R2480 VDD1.n92 VDD1.n91 9.45567
R2481 VDD1.n185 VDD1.n184 9.45567
R2482 VDD1.n58 VDD1.n57 9.3005
R2483 VDD1.n60 VDD1.n59 9.3005
R2484 VDD1.n15 VDD1.n14 9.3005
R2485 VDD1.n66 VDD1.n65 9.3005
R2486 VDD1.n68 VDD1.n67 9.3005
R2487 VDD1.n10 VDD1.n9 9.3005
R2488 VDD1.n74 VDD1.n73 9.3005
R2489 VDD1.n76 VDD1.n75 9.3005
R2490 VDD1.n91 VDD1.n90 9.3005
R2491 VDD1.n2 VDD1.n1 9.3005
R2492 VDD1.n85 VDD1.n84 9.3005
R2493 VDD1.n83 VDD1.n82 9.3005
R2494 VDD1.n6 VDD1.n5 9.3005
R2495 VDD1.n19 VDD1.n18 9.3005
R2496 VDD1.n52 VDD1.n51 9.3005
R2497 VDD1.n50 VDD1.n49 9.3005
R2498 VDD1.n23 VDD1.n22 9.3005
R2499 VDD1.n44 VDD1.n43 9.3005
R2500 VDD1.n42 VDD1.n41 9.3005
R2501 VDD1.n27 VDD1.n26 9.3005
R2502 VDD1.n36 VDD1.n35 9.3005
R2503 VDD1.n34 VDD1.n33 9.3005
R2504 VDD1.n184 VDD1.n183 9.3005
R2505 VDD1.n95 VDD1.n94 9.3005
R2506 VDD1.n178 VDD1.n177 9.3005
R2507 VDD1.n176 VDD1.n175 9.3005
R2508 VDD1.n99 VDD1.n98 9.3005
R2509 VDD1.n144 VDD1.n143 9.3005
R2510 VDD1.n142 VDD1.n141 9.3005
R2511 VDD1.n115 VDD1.n114 9.3005
R2512 VDD1.n136 VDD1.n135 9.3005
R2513 VDD1.n134 VDD1.n133 9.3005
R2514 VDD1.n119 VDD1.n118 9.3005
R2515 VDD1.n128 VDD1.n127 9.3005
R2516 VDD1.n126 VDD1.n125 9.3005
R2517 VDD1.n111 VDD1.n110 9.3005
R2518 VDD1.n150 VDD1.n149 9.3005
R2519 VDD1.n152 VDD1.n151 9.3005
R2520 VDD1.n107 VDD1.n106 9.3005
R2521 VDD1.n158 VDD1.n157 9.3005
R2522 VDD1.n160 VDD1.n159 9.3005
R2523 VDD1.n103 VDD1.n102 9.3005
R2524 VDD1.n167 VDD1.n166 9.3005
R2525 VDD1.n169 VDD1.n168 9.3005
R2526 VDD1.n61 VDD1.n15 8.92171
R2527 VDD1.n48 VDD1.n23 8.92171
R2528 VDD1.n140 VDD1.n115 8.92171
R2529 VDD1.n153 VDD1.n107 8.92171
R2530 VDD1.n60 VDD1.n17 8.14595
R2531 VDD1.n49 VDD1.n21 8.14595
R2532 VDD1.n141 VDD1.n113 8.14595
R2533 VDD1.n152 VDD1.n109 8.14595
R2534 VDD1.n57 VDD1.n56 7.3702
R2535 VDD1.n53 VDD1.n52 7.3702
R2536 VDD1.n145 VDD1.n144 7.3702
R2537 VDD1.n149 VDD1.n148 7.3702
R2538 VDD1.n56 VDD1.n19 6.59444
R2539 VDD1.n53 VDD1.n19 6.59444
R2540 VDD1.n145 VDD1.n111 6.59444
R2541 VDD1.n148 VDD1.n111 6.59444
R2542 VDD1.n57 VDD1.n17 5.81868
R2543 VDD1.n52 VDD1.n21 5.81868
R2544 VDD1.n144 VDD1.n113 5.81868
R2545 VDD1.n149 VDD1.n109 5.81868
R2546 VDD1.n61 VDD1.n60 5.04292
R2547 VDD1.n49 VDD1.n48 5.04292
R2548 VDD1.n141 VDD1.n140 5.04292
R2549 VDD1.n153 VDD1.n152 5.04292
R2550 VDD1.n34 VDD1.n30 4.38563
R2551 VDD1.n126 VDD1.n122 4.38563
R2552 VDD1.n92 VDD1.n0 4.26717
R2553 VDD1.n64 VDD1.n15 4.26717
R2554 VDD1.n45 VDD1.n23 4.26717
R2555 VDD1.n137 VDD1.n115 4.26717
R2556 VDD1.n156 VDD1.n107 4.26717
R2557 VDD1.n185 VDD1.n93 4.26717
R2558 VDD1.n90 VDD1.n89 3.49141
R2559 VDD1.n65 VDD1.n13 3.49141
R2560 VDD1.n44 VDD1.n25 3.49141
R2561 VDD1.n136 VDD1.n117 3.49141
R2562 VDD1.n157 VDD1.n105 3.49141
R2563 VDD1.n183 VDD1.n182 3.49141
R2564 VDD1.n86 VDD1.n2 2.71565
R2565 VDD1.n69 VDD1.n68 2.71565
R2566 VDD1.n41 VDD1.n40 2.71565
R2567 VDD1.n133 VDD1.n132 2.71565
R2568 VDD1.n161 VDD1.n160 2.71565
R2569 VDD1.n179 VDD1.n95 2.71565
R2570 VDD1.n85 VDD1.n4 1.93989
R2571 VDD1.n72 VDD1.n10 1.93989
R2572 VDD1.n37 VDD1.n27 1.93989
R2573 VDD1.n129 VDD1.n119 1.93989
R2574 VDD1.n165 VDD1.n103 1.93989
R2575 VDD1.n178 VDD1.n97 1.93989
R2576 VDD1.n188 VDD1.t0 1.17697
R2577 VDD1.n188 VDD1.t5 1.17697
R2578 VDD1.n186 VDD1.t4 1.17697
R2579 VDD1.n186 VDD1.t2 1.17697
R2580 VDD1.n82 VDD1.n81 1.16414
R2581 VDD1.n73 VDD1.n8 1.16414
R2582 VDD1.n36 VDD1.n29 1.16414
R2583 VDD1.n128 VDD1.n121 1.16414
R2584 VDD1.n166 VDD1.n101 1.16414
R2585 VDD1.n175 VDD1.n174 1.16414
R2586 VDD1.n78 VDD1.n6 0.388379
R2587 VDD1.n77 VDD1.n76 0.388379
R2588 VDD1.n33 VDD1.n32 0.388379
R2589 VDD1.n125 VDD1.n124 0.388379
R2590 VDD1.n170 VDD1.n169 0.388379
R2591 VDD1.n171 VDD1.n99 0.388379
R2592 VDD1 VDD1.n189 0.200931
R2593 VDD1.n91 VDD1.n1 0.155672
R2594 VDD1.n84 VDD1.n1 0.155672
R2595 VDD1.n84 VDD1.n83 0.155672
R2596 VDD1.n83 VDD1.n5 0.155672
R2597 VDD1.n75 VDD1.n5 0.155672
R2598 VDD1.n75 VDD1.n74 0.155672
R2599 VDD1.n74 VDD1.n9 0.155672
R2600 VDD1.n67 VDD1.n9 0.155672
R2601 VDD1.n67 VDD1.n66 0.155672
R2602 VDD1.n66 VDD1.n14 0.155672
R2603 VDD1.n59 VDD1.n14 0.155672
R2604 VDD1.n59 VDD1.n58 0.155672
R2605 VDD1.n58 VDD1.n18 0.155672
R2606 VDD1.n51 VDD1.n18 0.155672
R2607 VDD1.n51 VDD1.n50 0.155672
R2608 VDD1.n50 VDD1.n22 0.155672
R2609 VDD1.n43 VDD1.n22 0.155672
R2610 VDD1.n43 VDD1.n42 0.155672
R2611 VDD1.n42 VDD1.n26 0.155672
R2612 VDD1.n35 VDD1.n26 0.155672
R2613 VDD1.n35 VDD1.n34 0.155672
R2614 VDD1.n127 VDD1.n126 0.155672
R2615 VDD1.n127 VDD1.n118 0.155672
R2616 VDD1.n134 VDD1.n118 0.155672
R2617 VDD1.n135 VDD1.n134 0.155672
R2618 VDD1.n135 VDD1.n114 0.155672
R2619 VDD1.n142 VDD1.n114 0.155672
R2620 VDD1.n143 VDD1.n142 0.155672
R2621 VDD1.n143 VDD1.n110 0.155672
R2622 VDD1.n150 VDD1.n110 0.155672
R2623 VDD1.n151 VDD1.n150 0.155672
R2624 VDD1.n151 VDD1.n106 0.155672
R2625 VDD1.n158 VDD1.n106 0.155672
R2626 VDD1.n159 VDD1.n158 0.155672
R2627 VDD1.n159 VDD1.n102 0.155672
R2628 VDD1.n167 VDD1.n102 0.155672
R2629 VDD1.n168 VDD1.n167 0.155672
R2630 VDD1.n168 VDD1.n98 0.155672
R2631 VDD1.n176 VDD1.n98 0.155672
R2632 VDD1.n177 VDD1.n176 0.155672
R2633 VDD1.n177 VDD1.n94 0.155672
R2634 VDD1.n184 VDD1.n94 0.155672
C0 VP VN 6.14161f
C1 VDD2 VN 6.59276f
C2 VN VTAIL 6.13224f
C3 VDD2 VP 0.312675f
C4 VN VDD1 0.148398f
C5 VP VTAIL 6.14697f
C6 VDD2 VTAIL 12.132599f
C7 VP VDD1 6.75118f
C8 VDD2 VDD1 0.773981f
C9 VTAIL VDD1 12.0992f
C10 VDD2 B 5.489718f
C11 VDD1 B 5.521994f
C12 VTAIL B 8.341793f
C13 VN B 8.69303f
C14 VP B 6.603522f
C15 VDD1.n0 B 0.031244f
C16 VDD1.n1 B 0.022775f
C17 VDD1.n2 B 0.012238f
C18 VDD1.n3 B 0.028927f
C19 VDD1.n4 B 0.012958f
C20 VDD1.n5 B 0.022775f
C21 VDD1.n6 B 0.012238f
C22 VDD1.n7 B 0.028927f
C23 VDD1.n8 B 0.012958f
C24 VDD1.n9 B 0.022775f
C25 VDD1.n10 B 0.012238f
C26 VDD1.n11 B 0.028927f
C27 VDD1.n12 B 0.028927f
C28 VDD1.n13 B 0.012958f
C29 VDD1.n14 B 0.022775f
C30 VDD1.n15 B 0.012238f
C31 VDD1.n16 B 0.028927f
C32 VDD1.n17 B 0.012958f
C33 VDD1.n18 B 0.022775f
C34 VDD1.n19 B 0.012238f
C35 VDD1.n20 B 0.028927f
C36 VDD1.n21 B 0.012958f
C37 VDD1.n22 B 0.022775f
C38 VDD1.n23 B 0.012238f
C39 VDD1.n24 B 0.028927f
C40 VDD1.n25 B 0.012958f
C41 VDD1.n26 B 0.022775f
C42 VDD1.n27 B 0.012238f
C43 VDD1.n28 B 0.028927f
C44 VDD1.n29 B 0.012958f
C45 VDD1.n30 B 0.158995f
C46 VDD1.t3 B 0.04784f
C47 VDD1.n31 B 0.021695f
C48 VDD1.n32 B 0.017088f
C49 VDD1.n33 B 0.012238f
C50 VDD1.n34 B 1.6728f
C51 VDD1.n35 B 0.022775f
C52 VDD1.n36 B 0.012238f
C53 VDD1.n37 B 0.012958f
C54 VDD1.n38 B 0.028927f
C55 VDD1.n39 B 0.028927f
C56 VDD1.n40 B 0.012958f
C57 VDD1.n41 B 0.012238f
C58 VDD1.n42 B 0.022775f
C59 VDD1.n43 B 0.022775f
C60 VDD1.n44 B 0.012238f
C61 VDD1.n45 B 0.012958f
C62 VDD1.n46 B 0.028927f
C63 VDD1.n47 B 0.028927f
C64 VDD1.n48 B 0.012958f
C65 VDD1.n49 B 0.012238f
C66 VDD1.n50 B 0.022775f
C67 VDD1.n51 B 0.022775f
C68 VDD1.n52 B 0.012238f
C69 VDD1.n53 B 0.012958f
C70 VDD1.n54 B 0.028927f
C71 VDD1.n55 B 0.028927f
C72 VDD1.n56 B 0.012958f
C73 VDD1.n57 B 0.012238f
C74 VDD1.n58 B 0.022775f
C75 VDD1.n59 B 0.022775f
C76 VDD1.n60 B 0.012238f
C77 VDD1.n61 B 0.012958f
C78 VDD1.n62 B 0.028927f
C79 VDD1.n63 B 0.028927f
C80 VDD1.n64 B 0.012958f
C81 VDD1.n65 B 0.012238f
C82 VDD1.n66 B 0.022775f
C83 VDD1.n67 B 0.022775f
C84 VDD1.n68 B 0.012238f
C85 VDD1.n69 B 0.012958f
C86 VDD1.n70 B 0.028927f
C87 VDD1.n71 B 0.028927f
C88 VDD1.n72 B 0.012958f
C89 VDD1.n73 B 0.012238f
C90 VDD1.n74 B 0.022775f
C91 VDD1.n75 B 0.022775f
C92 VDD1.n76 B 0.012238f
C93 VDD1.n77 B 0.012598f
C94 VDD1.n78 B 0.012598f
C95 VDD1.n79 B 0.028927f
C96 VDD1.n80 B 0.028927f
C97 VDD1.n81 B 0.012958f
C98 VDD1.n82 B 0.012238f
C99 VDD1.n83 B 0.022775f
C100 VDD1.n84 B 0.022775f
C101 VDD1.n85 B 0.012238f
C102 VDD1.n86 B 0.012958f
C103 VDD1.n87 B 0.028927f
C104 VDD1.n88 B 0.061264f
C105 VDD1.n89 B 0.012958f
C106 VDD1.n90 B 0.012238f
C107 VDD1.n91 B 0.053577f
C108 VDD1.n92 B 0.051638f
C109 VDD1.n93 B 0.031244f
C110 VDD1.n94 B 0.022775f
C111 VDD1.n95 B 0.012238f
C112 VDD1.n96 B 0.028927f
C113 VDD1.n97 B 0.012958f
C114 VDD1.n98 B 0.022775f
C115 VDD1.n99 B 0.012238f
C116 VDD1.n100 B 0.028927f
C117 VDD1.n101 B 0.012958f
C118 VDD1.n102 B 0.022775f
C119 VDD1.n103 B 0.012238f
C120 VDD1.n104 B 0.028927f
C121 VDD1.n105 B 0.012958f
C122 VDD1.n106 B 0.022775f
C123 VDD1.n107 B 0.012238f
C124 VDD1.n108 B 0.028927f
C125 VDD1.n109 B 0.012958f
C126 VDD1.n110 B 0.022775f
C127 VDD1.n111 B 0.012238f
C128 VDD1.n112 B 0.028927f
C129 VDD1.n113 B 0.012958f
C130 VDD1.n114 B 0.022775f
C131 VDD1.n115 B 0.012238f
C132 VDD1.n116 B 0.028927f
C133 VDD1.n117 B 0.012958f
C134 VDD1.n118 B 0.022775f
C135 VDD1.n119 B 0.012238f
C136 VDD1.n120 B 0.028927f
C137 VDD1.n121 B 0.012958f
C138 VDD1.n122 B 0.158995f
C139 VDD1.t1 B 0.04784f
C140 VDD1.n123 B 0.021695f
C141 VDD1.n124 B 0.017088f
C142 VDD1.n125 B 0.012238f
C143 VDD1.n126 B 1.6728f
C144 VDD1.n127 B 0.022775f
C145 VDD1.n128 B 0.012238f
C146 VDD1.n129 B 0.012958f
C147 VDD1.n130 B 0.028927f
C148 VDD1.n131 B 0.028927f
C149 VDD1.n132 B 0.012958f
C150 VDD1.n133 B 0.012238f
C151 VDD1.n134 B 0.022775f
C152 VDD1.n135 B 0.022775f
C153 VDD1.n136 B 0.012238f
C154 VDD1.n137 B 0.012958f
C155 VDD1.n138 B 0.028927f
C156 VDD1.n139 B 0.028927f
C157 VDD1.n140 B 0.012958f
C158 VDD1.n141 B 0.012238f
C159 VDD1.n142 B 0.022775f
C160 VDD1.n143 B 0.022775f
C161 VDD1.n144 B 0.012238f
C162 VDD1.n145 B 0.012958f
C163 VDD1.n146 B 0.028927f
C164 VDD1.n147 B 0.028927f
C165 VDD1.n148 B 0.012958f
C166 VDD1.n149 B 0.012238f
C167 VDD1.n150 B 0.022775f
C168 VDD1.n151 B 0.022775f
C169 VDD1.n152 B 0.012238f
C170 VDD1.n153 B 0.012958f
C171 VDD1.n154 B 0.028927f
C172 VDD1.n155 B 0.028927f
C173 VDD1.n156 B 0.012958f
C174 VDD1.n157 B 0.012238f
C175 VDD1.n158 B 0.022775f
C176 VDD1.n159 B 0.022775f
C177 VDD1.n160 B 0.012238f
C178 VDD1.n161 B 0.012958f
C179 VDD1.n162 B 0.028927f
C180 VDD1.n163 B 0.028927f
C181 VDD1.n164 B 0.028927f
C182 VDD1.n165 B 0.012958f
C183 VDD1.n166 B 0.012238f
C184 VDD1.n167 B 0.022775f
C185 VDD1.n168 B 0.022775f
C186 VDD1.n169 B 0.012238f
C187 VDD1.n170 B 0.012598f
C188 VDD1.n171 B 0.012598f
C189 VDD1.n172 B 0.028927f
C190 VDD1.n173 B 0.028927f
C191 VDD1.n174 B 0.012958f
C192 VDD1.n175 B 0.012238f
C193 VDD1.n176 B 0.022775f
C194 VDD1.n177 B 0.022775f
C195 VDD1.n178 B 0.012238f
C196 VDD1.n179 B 0.012958f
C197 VDD1.n180 B 0.028927f
C198 VDD1.n181 B 0.061264f
C199 VDD1.n182 B 0.012958f
C200 VDD1.n183 B 0.012238f
C201 VDD1.n184 B 0.053577f
C202 VDD1.n185 B 0.051294f
C203 VDD1.t4 B 0.302901f
C204 VDD1.t2 B 0.302901f
C205 VDD1.n186 B 2.75331f
C206 VDD1.n187 B 2.10276f
C207 VDD1.t0 B 0.302901f
C208 VDD1.t5 B 0.302901f
C209 VDD1.n188 B 2.75235f
C210 VDD1.n189 B 2.4351f
C211 VP.n0 B 0.042252f
C212 VP.t1 B 1.69944f
C213 VP.n1 B 0.616805f
C214 VP.n2 B 0.042252f
C215 VP.n3 B 0.042252f
C216 VP.t0 B 1.75576f
C217 VP.t5 B 1.69944f
C218 VP.n4 B 0.655277f
C219 VP.t2 B 1.77639f
C220 VP.n5 B 0.667027f
C221 VP.n6 B 0.175191f
C222 VP.n7 B 0.053688f
C223 VP.n8 B 0.013302f
C224 VP.n9 B 0.658289f
C225 VP.n10 B 1.9867f
C226 VP.n11 B 2.02007f
C227 VP.t4 B 1.75576f
C228 VP.n12 B 0.658289f
C229 VP.n13 B 0.013302f
C230 VP.n14 B 0.053688f
C231 VP.n15 B 0.042252f
C232 VP.n16 B 0.042252f
C233 VP.n17 B 0.053688f
C234 VP.n18 B 0.013302f
C235 VP.t3 B 1.75576f
C236 VP.n19 B 0.658289f
C237 VP.n20 B 0.032744f
C238 VTAIL.t9 B 0.30755f
C239 VTAIL.t5 B 0.30755f
C240 VTAIL.n0 B 2.72499f
C241 VTAIL.n1 B 0.325958f
C242 VTAIL.n2 B 0.031724f
C243 VTAIL.n3 B 0.023125f
C244 VTAIL.n4 B 0.012426f
C245 VTAIL.n5 B 0.029371f
C246 VTAIL.n6 B 0.013157f
C247 VTAIL.n7 B 0.023125f
C248 VTAIL.n8 B 0.012426f
C249 VTAIL.n9 B 0.029371f
C250 VTAIL.n10 B 0.013157f
C251 VTAIL.n11 B 0.023125f
C252 VTAIL.n12 B 0.012426f
C253 VTAIL.n13 B 0.029371f
C254 VTAIL.n14 B 0.013157f
C255 VTAIL.n15 B 0.023125f
C256 VTAIL.n16 B 0.012426f
C257 VTAIL.n17 B 0.029371f
C258 VTAIL.n18 B 0.013157f
C259 VTAIL.n19 B 0.023125f
C260 VTAIL.n20 B 0.012426f
C261 VTAIL.n21 B 0.029371f
C262 VTAIL.n22 B 0.013157f
C263 VTAIL.n23 B 0.023125f
C264 VTAIL.n24 B 0.012426f
C265 VTAIL.n25 B 0.029371f
C266 VTAIL.n26 B 0.013157f
C267 VTAIL.n27 B 0.023125f
C268 VTAIL.n28 B 0.012426f
C269 VTAIL.n29 B 0.029371f
C270 VTAIL.n30 B 0.013157f
C271 VTAIL.n31 B 0.161435f
C272 VTAIL.t4 B 0.048575f
C273 VTAIL.n32 B 0.022028f
C274 VTAIL.n33 B 0.01735f
C275 VTAIL.n34 B 0.012426f
C276 VTAIL.n35 B 1.69848f
C277 VTAIL.n36 B 0.023125f
C278 VTAIL.n37 B 0.012426f
C279 VTAIL.n38 B 0.013157f
C280 VTAIL.n39 B 0.029371f
C281 VTAIL.n40 B 0.029371f
C282 VTAIL.n41 B 0.013157f
C283 VTAIL.n42 B 0.012426f
C284 VTAIL.n43 B 0.023125f
C285 VTAIL.n44 B 0.023125f
C286 VTAIL.n45 B 0.012426f
C287 VTAIL.n46 B 0.013157f
C288 VTAIL.n47 B 0.029371f
C289 VTAIL.n48 B 0.029371f
C290 VTAIL.n49 B 0.013157f
C291 VTAIL.n50 B 0.012426f
C292 VTAIL.n51 B 0.023125f
C293 VTAIL.n52 B 0.023125f
C294 VTAIL.n53 B 0.012426f
C295 VTAIL.n54 B 0.013157f
C296 VTAIL.n55 B 0.029371f
C297 VTAIL.n56 B 0.029371f
C298 VTAIL.n57 B 0.013157f
C299 VTAIL.n58 B 0.012426f
C300 VTAIL.n59 B 0.023125f
C301 VTAIL.n60 B 0.023125f
C302 VTAIL.n61 B 0.012426f
C303 VTAIL.n62 B 0.013157f
C304 VTAIL.n63 B 0.029371f
C305 VTAIL.n64 B 0.029371f
C306 VTAIL.n65 B 0.013157f
C307 VTAIL.n66 B 0.012426f
C308 VTAIL.n67 B 0.023125f
C309 VTAIL.n68 B 0.023125f
C310 VTAIL.n69 B 0.012426f
C311 VTAIL.n70 B 0.013157f
C312 VTAIL.n71 B 0.029371f
C313 VTAIL.n72 B 0.029371f
C314 VTAIL.n73 B 0.029371f
C315 VTAIL.n74 B 0.013157f
C316 VTAIL.n75 B 0.012426f
C317 VTAIL.n76 B 0.023125f
C318 VTAIL.n77 B 0.023125f
C319 VTAIL.n78 B 0.012426f
C320 VTAIL.n79 B 0.012792f
C321 VTAIL.n80 B 0.012792f
C322 VTAIL.n81 B 0.029371f
C323 VTAIL.n82 B 0.029371f
C324 VTAIL.n83 B 0.013157f
C325 VTAIL.n84 B 0.012426f
C326 VTAIL.n85 B 0.023125f
C327 VTAIL.n86 B 0.023125f
C328 VTAIL.n87 B 0.012426f
C329 VTAIL.n88 B 0.013157f
C330 VTAIL.n89 B 0.029371f
C331 VTAIL.n90 B 0.062204f
C332 VTAIL.n91 B 0.013157f
C333 VTAIL.n92 B 0.012426f
C334 VTAIL.n93 B 0.0544f
C335 VTAIL.n94 B 0.034693f
C336 VTAIL.n95 B 0.170918f
C337 VTAIL.t2 B 0.30755f
C338 VTAIL.t3 B 0.30755f
C339 VTAIL.n96 B 2.72499f
C340 VTAIL.n97 B 1.85526f
C341 VTAIL.t7 B 0.30755f
C342 VTAIL.t10 B 0.30755f
C343 VTAIL.n98 B 2.725f
C344 VTAIL.n99 B 1.85524f
C345 VTAIL.n100 B 0.031724f
C346 VTAIL.n101 B 0.023125f
C347 VTAIL.n102 B 0.012426f
C348 VTAIL.n103 B 0.029371f
C349 VTAIL.n104 B 0.013157f
C350 VTAIL.n105 B 0.023125f
C351 VTAIL.n106 B 0.012426f
C352 VTAIL.n107 B 0.029371f
C353 VTAIL.n108 B 0.013157f
C354 VTAIL.n109 B 0.023125f
C355 VTAIL.n110 B 0.012426f
C356 VTAIL.n111 B 0.029371f
C357 VTAIL.n112 B 0.029371f
C358 VTAIL.n113 B 0.013157f
C359 VTAIL.n114 B 0.023125f
C360 VTAIL.n115 B 0.012426f
C361 VTAIL.n116 B 0.029371f
C362 VTAIL.n117 B 0.013157f
C363 VTAIL.n118 B 0.023125f
C364 VTAIL.n119 B 0.012426f
C365 VTAIL.n120 B 0.029371f
C366 VTAIL.n121 B 0.013157f
C367 VTAIL.n122 B 0.023125f
C368 VTAIL.n123 B 0.012426f
C369 VTAIL.n124 B 0.029371f
C370 VTAIL.n125 B 0.013157f
C371 VTAIL.n126 B 0.023125f
C372 VTAIL.n127 B 0.012426f
C373 VTAIL.n128 B 0.029371f
C374 VTAIL.n129 B 0.013157f
C375 VTAIL.n130 B 0.161435f
C376 VTAIL.t8 B 0.048575f
C377 VTAIL.n131 B 0.022028f
C378 VTAIL.n132 B 0.01735f
C379 VTAIL.n133 B 0.012426f
C380 VTAIL.n134 B 1.69848f
C381 VTAIL.n135 B 0.023125f
C382 VTAIL.n136 B 0.012426f
C383 VTAIL.n137 B 0.013157f
C384 VTAIL.n138 B 0.029371f
C385 VTAIL.n139 B 0.029371f
C386 VTAIL.n140 B 0.013157f
C387 VTAIL.n141 B 0.012426f
C388 VTAIL.n142 B 0.023125f
C389 VTAIL.n143 B 0.023125f
C390 VTAIL.n144 B 0.012426f
C391 VTAIL.n145 B 0.013157f
C392 VTAIL.n146 B 0.029371f
C393 VTAIL.n147 B 0.029371f
C394 VTAIL.n148 B 0.013157f
C395 VTAIL.n149 B 0.012426f
C396 VTAIL.n150 B 0.023125f
C397 VTAIL.n151 B 0.023125f
C398 VTAIL.n152 B 0.012426f
C399 VTAIL.n153 B 0.013157f
C400 VTAIL.n154 B 0.029371f
C401 VTAIL.n155 B 0.029371f
C402 VTAIL.n156 B 0.013157f
C403 VTAIL.n157 B 0.012426f
C404 VTAIL.n158 B 0.023125f
C405 VTAIL.n159 B 0.023125f
C406 VTAIL.n160 B 0.012426f
C407 VTAIL.n161 B 0.013157f
C408 VTAIL.n162 B 0.029371f
C409 VTAIL.n163 B 0.029371f
C410 VTAIL.n164 B 0.013157f
C411 VTAIL.n165 B 0.012426f
C412 VTAIL.n166 B 0.023125f
C413 VTAIL.n167 B 0.023125f
C414 VTAIL.n168 B 0.012426f
C415 VTAIL.n169 B 0.013157f
C416 VTAIL.n170 B 0.029371f
C417 VTAIL.n171 B 0.029371f
C418 VTAIL.n172 B 0.013157f
C419 VTAIL.n173 B 0.012426f
C420 VTAIL.n174 B 0.023125f
C421 VTAIL.n175 B 0.023125f
C422 VTAIL.n176 B 0.012426f
C423 VTAIL.n177 B 0.012792f
C424 VTAIL.n178 B 0.012792f
C425 VTAIL.n179 B 0.029371f
C426 VTAIL.n180 B 0.029371f
C427 VTAIL.n181 B 0.013157f
C428 VTAIL.n182 B 0.012426f
C429 VTAIL.n183 B 0.023125f
C430 VTAIL.n184 B 0.023125f
C431 VTAIL.n185 B 0.012426f
C432 VTAIL.n186 B 0.013157f
C433 VTAIL.n187 B 0.029371f
C434 VTAIL.n188 B 0.062204f
C435 VTAIL.n189 B 0.013157f
C436 VTAIL.n190 B 0.012426f
C437 VTAIL.n191 B 0.0544f
C438 VTAIL.n192 B 0.034693f
C439 VTAIL.n193 B 0.170918f
C440 VTAIL.t1 B 0.30755f
C441 VTAIL.t11 B 0.30755f
C442 VTAIL.n194 B 2.725f
C443 VTAIL.n195 B 0.379421f
C444 VTAIL.n196 B 0.031724f
C445 VTAIL.n197 B 0.023125f
C446 VTAIL.n198 B 0.012426f
C447 VTAIL.n199 B 0.029371f
C448 VTAIL.n200 B 0.013157f
C449 VTAIL.n201 B 0.023125f
C450 VTAIL.n202 B 0.012426f
C451 VTAIL.n203 B 0.029371f
C452 VTAIL.n204 B 0.013157f
C453 VTAIL.n205 B 0.023125f
C454 VTAIL.n206 B 0.012426f
C455 VTAIL.n207 B 0.029371f
C456 VTAIL.n208 B 0.029371f
C457 VTAIL.n209 B 0.013157f
C458 VTAIL.n210 B 0.023125f
C459 VTAIL.n211 B 0.012426f
C460 VTAIL.n212 B 0.029371f
C461 VTAIL.n213 B 0.013157f
C462 VTAIL.n214 B 0.023125f
C463 VTAIL.n215 B 0.012426f
C464 VTAIL.n216 B 0.029371f
C465 VTAIL.n217 B 0.013157f
C466 VTAIL.n218 B 0.023125f
C467 VTAIL.n219 B 0.012426f
C468 VTAIL.n220 B 0.029371f
C469 VTAIL.n221 B 0.013157f
C470 VTAIL.n222 B 0.023125f
C471 VTAIL.n223 B 0.012426f
C472 VTAIL.n224 B 0.029371f
C473 VTAIL.n225 B 0.013157f
C474 VTAIL.n226 B 0.161435f
C475 VTAIL.t0 B 0.048575f
C476 VTAIL.n227 B 0.022028f
C477 VTAIL.n228 B 0.01735f
C478 VTAIL.n229 B 0.012426f
C479 VTAIL.n230 B 1.69848f
C480 VTAIL.n231 B 0.023125f
C481 VTAIL.n232 B 0.012426f
C482 VTAIL.n233 B 0.013157f
C483 VTAIL.n234 B 0.029371f
C484 VTAIL.n235 B 0.029371f
C485 VTAIL.n236 B 0.013157f
C486 VTAIL.n237 B 0.012426f
C487 VTAIL.n238 B 0.023125f
C488 VTAIL.n239 B 0.023125f
C489 VTAIL.n240 B 0.012426f
C490 VTAIL.n241 B 0.013157f
C491 VTAIL.n242 B 0.029371f
C492 VTAIL.n243 B 0.029371f
C493 VTAIL.n244 B 0.013157f
C494 VTAIL.n245 B 0.012426f
C495 VTAIL.n246 B 0.023125f
C496 VTAIL.n247 B 0.023125f
C497 VTAIL.n248 B 0.012426f
C498 VTAIL.n249 B 0.013157f
C499 VTAIL.n250 B 0.029371f
C500 VTAIL.n251 B 0.029371f
C501 VTAIL.n252 B 0.013157f
C502 VTAIL.n253 B 0.012426f
C503 VTAIL.n254 B 0.023125f
C504 VTAIL.n255 B 0.023125f
C505 VTAIL.n256 B 0.012426f
C506 VTAIL.n257 B 0.013157f
C507 VTAIL.n258 B 0.029371f
C508 VTAIL.n259 B 0.029371f
C509 VTAIL.n260 B 0.013157f
C510 VTAIL.n261 B 0.012426f
C511 VTAIL.n262 B 0.023125f
C512 VTAIL.n263 B 0.023125f
C513 VTAIL.n264 B 0.012426f
C514 VTAIL.n265 B 0.013157f
C515 VTAIL.n266 B 0.029371f
C516 VTAIL.n267 B 0.029371f
C517 VTAIL.n268 B 0.013157f
C518 VTAIL.n269 B 0.012426f
C519 VTAIL.n270 B 0.023125f
C520 VTAIL.n271 B 0.023125f
C521 VTAIL.n272 B 0.012426f
C522 VTAIL.n273 B 0.012792f
C523 VTAIL.n274 B 0.012792f
C524 VTAIL.n275 B 0.029371f
C525 VTAIL.n276 B 0.029371f
C526 VTAIL.n277 B 0.013157f
C527 VTAIL.n278 B 0.012426f
C528 VTAIL.n279 B 0.023125f
C529 VTAIL.n280 B 0.023125f
C530 VTAIL.n281 B 0.012426f
C531 VTAIL.n282 B 0.013157f
C532 VTAIL.n283 B 0.029371f
C533 VTAIL.n284 B 0.062204f
C534 VTAIL.n285 B 0.013157f
C535 VTAIL.n286 B 0.012426f
C536 VTAIL.n287 B 0.0544f
C537 VTAIL.n288 B 0.034693f
C538 VTAIL.n289 B 1.56966f
C539 VTAIL.n290 B 0.031724f
C540 VTAIL.n291 B 0.023125f
C541 VTAIL.n292 B 0.012426f
C542 VTAIL.n293 B 0.029371f
C543 VTAIL.n294 B 0.013157f
C544 VTAIL.n295 B 0.023125f
C545 VTAIL.n296 B 0.012426f
C546 VTAIL.n297 B 0.029371f
C547 VTAIL.n298 B 0.013157f
C548 VTAIL.n299 B 0.023125f
C549 VTAIL.n300 B 0.012426f
C550 VTAIL.n301 B 0.029371f
C551 VTAIL.n302 B 0.013157f
C552 VTAIL.n303 B 0.023125f
C553 VTAIL.n304 B 0.012426f
C554 VTAIL.n305 B 0.029371f
C555 VTAIL.n306 B 0.013157f
C556 VTAIL.n307 B 0.023125f
C557 VTAIL.n308 B 0.012426f
C558 VTAIL.n309 B 0.029371f
C559 VTAIL.n310 B 0.013157f
C560 VTAIL.n311 B 0.023125f
C561 VTAIL.n312 B 0.012426f
C562 VTAIL.n313 B 0.029371f
C563 VTAIL.n314 B 0.013157f
C564 VTAIL.n315 B 0.023125f
C565 VTAIL.n316 B 0.012426f
C566 VTAIL.n317 B 0.029371f
C567 VTAIL.n318 B 0.013157f
C568 VTAIL.n319 B 0.161435f
C569 VTAIL.t6 B 0.048575f
C570 VTAIL.n320 B 0.022028f
C571 VTAIL.n321 B 0.01735f
C572 VTAIL.n322 B 0.012426f
C573 VTAIL.n323 B 1.69848f
C574 VTAIL.n324 B 0.023125f
C575 VTAIL.n325 B 0.012426f
C576 VTAIL.n326 B 0.013157f
C577 VTAIL.n327 B 0.029371f
C578 VTAIL.n328 B 0.029371f
C579 VTAIL.n329 B 0.013157f
C580 VTAIL.n330 B 0.012426f
C581 VTAIL.n331 B 0.023125f
C582 VTAIL.n332 B 0.023125f
C583 VTAIL.n333 B 0.012426f
C584 VTAIL.n334 B 0.013157f
C585 VTAIL.n335 B 0.029371f
C586 VTAIL.n336 B 0.029371f
C587 VTAIL.n337 B 0.013157f
C588 VTAIL.n338 B 0.012426f
C589 VTAIL.n339 B 0.023125f
C590 VTAIL.n340 B 0.023125f
C591 VTAIL.n341 B 0.012426f
C592 VTAIL.n342 B 0.013157f
C593 VTAIL.n343 B 0.029371f
C594 VTAIL.n344 B 0.029371f
C595 VTAIL.n345 B 0.013157f
C596 VTAIL.n346 B 0.012426f
C597 VTAIL.n347 B 0.023125f
C598 VTAIL.n348 B 0.023125f
C599 VTAIL.n349 B 0.012426f
C600 VTAIL.n350 B 0.013157f
C601 VTAIL.n351 B 0.029371f
C602 VTAIL.n352 B 0.029371f
C603 VTAIL.n353 B 0.013157f
C604 VTAIL.n354 B 0.012426f
C605 VTAIL.n355 B 0.023125f
C606 VTAIL.n356 B 0.023125f
C607 VTAIL.n357 B 0.012426f
C608 VTAIL.n358 B 0.013157f
C609 VTAIL.n359 B 0.029371f
C610 VTAIL.n360 B 0.029371f
C611 VTAIL.n361 B 0.029371f
C612 VTAIL.n362 B 0.013157f
C613 VTAIL.n363 B 0.012426f
C614 VTAIL.n364 B 0.023125f
C615 VTAIL.n365 B 0.023125f
C616 VTAIL.n366 B 0.012426f
C617 VTAIL.n367 B 0.012792f
C618 VTAIL.n368 B 0.012792f
C619 VTAIL.n369 B 0.029371f
C620 VTAIL.n370 B 0.029371f
C621 VTAIL.n371 B 0.013157f
C622 VTAIL.n372 B 0.012426f
C623 VTAIL.n373 B 0.023125f
C624 VTAIL.n374 B 0.023125f
C625 VTAIL.n375 B 0.012426f
C626 VTAIL.n376 B 0.013157f
C627 VTAIL.n377 B 0.029371f
C628 VTAIL.n378 B 0.062204f
C629 VTAIL.n379 B 0.013157f
C630 VTAIL.n380 B 0.012426f
C631 VTAIL.n381 B 0.0544f
C632 VTAIL.n382 B 0.034693f
C633 VTAIL.n383 B 1.54605f
C634 VDD2.n0 B 0.031052f
C635 VDD2.n1 B 0.022635f
C636 VDD2.n2 B 0.012163f
C637 VDD2.n3 B 0.028749f
C638 VDD2.n4 B 0.012878f
C639 VDD2.n5 B 0.022635f
C640 VDD2.n6 B 0.012163f
C641 VDD2.n7 B 0.028749f
C642 VDD2.n8 B 0.012878f
C643 VDD2.n9 B 0.022635f
C644 VDD2.n10 B 0.012163f
C645 VDD2.n11 B 0.028749f
C646 VDD2.n12 B 0.012878f
C647 VDD2.n13 B 0.022635f
C648 VDD2.n14 B 0.012163f
C649 VDD2.n15 B 0.028749f
C650 VDD2.n16 B 0.012878f
C651 VDD2.n17 B 0.022635f
C652 VDD2.n18 B 0.012163f
C653 VDD2.n19 B 0.028749f
C654 VDD2.n20 B 0.012878f
C655 VDD2.n21 B 0.022635f
C656 VDD2.n22 B 0.012163f
C657 VDD2.n23 B 0.028749f
C658 VDD2.n24 B 0.012878f
C659 VDD2.n25 B 0.022635f
C660 VDD2.n26 B 0.012163f
C661 VDD2.n27 B 0.028749f
C662 VDD2.n28 B 0.012878f
C663 VDD2.n29 B 0.158016f
C664 VDD2.t4 B 0.047546f
C665 VDD2.n30 B 0.021562f
C666 VDD2.n31 B 0.016983f
C667 VDD2.n32 B 0.012163f
C668 VDD2.n33 B 1.6625f
C669 VDD2.n34 B 0.022635f
C670 VDD2.n35 B 0.012163f
C671 VDD2.n36 B 0.012878f
C672 VDD2.n37 B 0.028749f
C673 VDD2.n38 B 0.028749f
C674 VDD2.n39 B 0.012878f
C675 VDD2.n40 B 0.012163f
C676 VDD2.n41 B 0.022635f
C677 VDD2.n42 B 0.022635f
C678 VDD2.n43 B 0.012163f
C679 VDD2.n44 B 0.012878f
C680 VDD2.n45 B 0.028749f
C681 VDD2.n46 B 0.028749f
C682 VDD2.n47 B 0.012878f
C683 VDD2.n48 B 0.012163f
C684 VDD2.n49 B 0.022635f
C685 VDD2.n50 B 0.022635f
C686 VDD2.n51 B 0.012163f
C687 VDD2.n52 B 0.012878f
C688 VDD2.n53 B 0.028749f
C689 VDD2.n54 B 0.028749f
C690 VDD2.n55 B 0.012878f
C691 VDD2.n56 B 0.012163f
C692 VDD2.n57 B 0.022635f
C693 VDD2.n58 B 0.022635f
C694 VDD2.n59 B 0.012163f
C695 VDD2.n60 B 0.012878f
C696 VDD2.n61 B 0.028749f
C697 VDD2.n62 B 0.028749f
C698 VDD2.n63 B 0.012878f
C699 VDD2.n64 B 0.012163f
C700 VDD2.n65 B 0.022635f
C701 VDD2.n66 B 0.022635f
C702 VDD2.n67 B 0.012163f
C703 VDD2.n68 B 0.012878f
C704 VDD2.n69 B 0.028749f
C705 VDD2.n70 B 0.028749f
C706 VDD2.n71 B 0.028749f
C707 VDD2.n72 B 0.012878f
C708 VDD2.n73 B 0.012163f
C709 VDD2.n74 B 0.022635f
C710 VDD2.n75 B 0.022635f
C711 VDD2.n76 B 0.012163f
C712 VDD2.n77 B 0.012521f
C713 VDD2.n78 B 0.012521f
C714 VDD2.n79 B 0.028749f
C715 VDD2.n80 B 0.028749f
C716 VDD2.n81 B 0.012878f
C717 VDD2.n82 B 0.012163f
C718 VDD2.n83 B 0.022635f
C719 VDD2.n84 B 0.022635f
C720 VDD2.n85 B 0.012163f
C721 VDD2.n86 B 0.012878f
C722 VDD2.n87 B 0.028749f
C723 VDD2.n88 B 0.060887f
C724 VDD2.n89 B 0.012878f
C725 VDD2.n90 B 0.012163f
C726 VDD2.n91 B 0.053247f
C727 VDD2.n92 B 0.050978f
C728 VDD2.t1 B 0.301035f
C729 VDD2.t0 B 0.301035f
C730 VDD2.n93 B 2.73635f
C731 VDD2.n94 B 2.01499f
C732 VDD2.n95 B 0.031052f
C733 VDD2.n96 B 0.022635f
C734 VDD2.n97 B 0.012163f
C735 VDD2.n98 B 0.028749f
C736 VDD2.n99 B 0.012878f
C737 VDD2.n100 B 0.022635f
C738 VDD2.n101 B 0.012163f
C739 VDD2.n102 B 0.028749f
C740 VDD2.n103 B 0.012878f
C741 VDD2.n104 B 0.022635f
C742 VDD2.n105 B 0.012163f
C743 VDD2.n106 B 0.028749f
C744 VDD2.n107 B 0.028749f
C745 VDD2.n108 B 0.012878f
C746 VDD2.n109 B 0.022635f
C747 VDD2.n110 B 0.012163f
C748 VDD2.n111 B 0.028749f
C749 VDD2.n112 B 0.012878f
C750 VDD2.n113 B 0.022635f
C751 VDD2.n114 B 0.012163f
C752 VDD2.n115 B 0.028749f
C753 VDD2.n116 B 0.012878f
C754 VDD2.n117 B 0.022635f
C755 VDD2.n118 B 0.012163f
C756 VDD2.n119 B 0.028749f
C757 VDD2.n120 B 0.012878f
C758 VDD2.n121 B 0.022635f
C759 VDD2.n122 B 0.012163f
C760 VDD2.n123 B 0.028749f
C761 VDD2.n124 B 0.012878f
C762 VDD2.n125 B 0.158016f
C763 VDD2.t2 B 0.047546f
C764 VDD2.n126 B 0.021562f
C765 VDD2.n127 B 0.016983f
C766 VDD2.n128 B 0.012163f
C767 VDD2.n129 B 1.6625f
C768 VDD2.n130 B 0.022635f
C769 VDD2.n131 B 0.012163f
C770 VDD2.n132 B 0.012878f
C771 VDD2.n133 B 0.028749f
C772 VDD2.n134 B 0.028749f
C773 VDD2.n135 B 0.012878f
C774 VDD2.n136 B 0.012163f
C775 VDD2.n137 B 0.022635f
C776 VDD2.n138 B 0.022635f
C777 VDD2.n139 B 0.012163f
C778 VDD2.n140 B 0.012878f
C779 VDD2.n141 B 0.028749f
C780 VDD2.n142 B 0.028749f
C781 VDD2.n143 B 0.012878f
C782 VDD2.n144 B 0.012163f
C783 VDD2.n145 B 0.022635f
C784 VDD2.n146 B 0.022635f
C785 VDD2.n147 B 0.012163f
C786 VDD2.n148 B 0.012878f
C787 VDD2.n149 B 0.028749f
C788 VDD2.n150 B 0.028749f
C789 VDD2.n151 B 0.012878f
C790 VDD2.n152 B 0.012163f
C791 VDD2.n153 B 0.022635f
C792 VDD2.n154 B 0.022635f
C793 VDD2.n155 B 0.012163f
C794 VDD2.n156 B 0.012878f
C795 VDD2.n157 B 0.028749f
C796 VDD2.n158 B 0.028749f
C797 VDD2.n159 B 0.012878f
C798 VDD2.n160 B 0.012163f
C799 VDD2.n161 B 0.022635f
C800 VDD2.n162 B 0.022635f
C801 VDD2.n163 B 0.012163f
C802 VDD2.n164 B 0.012878f
C803 VDD2.n165 B 0.028749f
C804 VDD2.n166 B 0.028749f
C805 VDD2.n167 B 0.012878f
C806 VDD2.n168 B 0.012163f
C807 VDD2.n169 B 0.022635f
C808 VDD2.n170 B 0.022635f
C809 VDD2.n171 B 0.012163f
C810 VDD2.n172 B 0.012521f
C811 VDD2.n173 B 0.012521f
C812 VDD2.n174 B 0.028749f
C813 VDD2.n175 B 0.028749f
C814 VDD2.n176 B 0.012878f
C815 VDD2.n177 B 0.012163f
C816 VDD2.n178 B 0.022635f
C817 VDD2.n179 B 0.022635f
C818 VDD2.n180 B 0.012163f
C819 VDD2.n181 B 0.012878f
C820 VDD2.n182 B 0.028749f
C821 VDD2.n183 B 0.060887f
C822 VDD2.n184 B 0.012878f
C823 VDD2.n185 B 0.012163f
C824 VDD2.n186 B 0.053247f
C825 VDD2.n187 B 0.049579f
C826 VDD2.n188 B 2.23049f
C827 VDD2.t3 B 0.301035f
C828 VDD2.t5 B 0.301035f
C829 VDD2.n189 B 2.73633f
C830 VN.n0 B 0.041677f
C831 VN.t5 B 1.67631f
C832 VN.n1 B 0.646358f
C833 VN.t1 B 1.75221f
C834 VN.n2 B 0.657949f
C835 VN.n3 B 0.172806f
C836 VN.n4 B 0.052958f
C837 VN.n5 B 0.013121f
C838 VN.t4 B 1.73186f
C839 VN.n6 B 0.64933f
C840 VN.n7 B 0.032298f
C841 VN.n8 B 0.041677f
C842 VN.t0 B 1.67631f
C843 VN.n9 B 0.646358f
C844 VN.t2 B 1.75221f
C845 VN.n10 B 0.657949f
C846 VN.n11 B 0.172806f
C847 VN.n12 B 0.052958f
C848 VN.n13 B 0.013121f
C849 VN.t3 B 1.73186f
C850 VN.n14 B 0.64933f
C851 VN.n15 B 1.98689f
.ends

