* NGSPICE file created from diff_pair_sample_0677.ext - technology: sky130A

.subckt diff_pair_sample_0677 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t1 VP.t0 VTAIL.t1 B.t0 sky130_fd_pr__nfet_01v8 ad=7.3242 pd=38.34 as=7.3242 ps=38.34 w=18.78 l=2.3
X1 B.t15 B.t13 B.t14 B.t3 sky130_fd_pr__nfet_01v8 ad=7.3242 pd=38.34 as=0 ps=0 w=18.78 l=2.3
X2 VDD2.t1 VN.t0 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=7.3242 pd=38.34 as=7.3242 ps=38.34 w=18.78 l=2.3
X3 B.t12 B.t10 B.t11 B.t7 sky130_fd_pr__nfet_01v8 ad=7.3242 pd=38.34 as=0 ps=0 w=18.78 l=2.3
X4 VDD1.t0 VP.t1 VTAIL.t2 B.t1 sky130_fd_pr__nfet_01v8 ad=7.3242 pd=38.34 as=7.3242 ps=38.34 w=18.78 l=2.3
X5 B.t9 B.t6 B.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=7.3242 pd=38.34 as=0 ps=0 w=18.78 l=2.3
X6 VDD2.t0 VN.t1 VTAIL.t3 B.t1 sky130_fd_pr__nfet_01v8 ad=7.3242 pd=38.34 as=7.3242 ps=38.34 w=18.78 l=2.3
X7 B.t5 B.t2 B.t4 B.t3 sky130_fd_pr__nfet_01v8 ad=7.3242 pd=38.34 as=0 ps=0 w=18.78 l=2.3
R0 VP.n0 VP.t0 294.906
R1 VP.n0 VP.t1 245.909
R2 VP VP.n0 0.336784
R3 VTAIL.n414 VTAIL.n413 289.615
R4 VTAIL.n102 VTAIL.n101 289.615
R5 VTAIL.n310 VTAIL.n309 289.615
R6 VTAIL.n206 VTAIL.n205 289.615
R7 VTAIL.n347 VTAIL.n346 185
R8 VTAIL.n349 VTAIL.n348 185
R9 VTAIL.n342 VTAIL.n341 185
R10 VTAIL.n355 VTAIL.n354 185
R11 VTAIL.n357 VTAIL.n356 185
R12 VTAIL.n338 VTAIL.n337 185
R13 VTAIL.n364 VTAIL.n363 185
R14 VTAIL.n365 VTAIL.n336 185
R15 VTAIL.n367 VTAIL.n366 185
R16 VTAIL.n334 VTAIL.n333 185
R17 VTAIL.n373 VTAIL.n372 185
R18 VTAIL.n375 VTAIL.n374 185
R19 VTAIL.n330 VTAIL.n329 185
R20 VTAIL.n381 VTAIL.n380 185
R21 VTAIL.n383 VTAIL.n382 185
R22 VTAIL.n326 VTAIL.n325 185
R23 VTAIL.n389 VTAIL.n388 185
R24 VTAIL.n391 VTAIL.n390 185
R25 VTAIL.n322 VTAIL.n321 185
R26 VTAIL.n397 VTAIL.n396 185
R27 VTAIL.n399 VTAIL.n398 185
R28 VTAIL.n318 VTAIL.n317 185
R29 VTAIL.n405 VTAIL.n404 185
R30 VTAIL.n407 VTAIL.n406 185
R31 VTAIL.n314 VTAIL.n313 185
R32 VTAIL.n413 VTAIL.n412 185
R33 VTAIL.n35 VTAIL.n34 185
R34 VTAIL.n37 VTAIL.n36 185
R35 VTAIL.n30 VTAIL.n29 185
R36 VTAIL.n43 VTAIL.n42 185
R37 VTAIL.n45 VTAIL.n44 185
R38 VTAIL.n26 VTAIL.n25 185
R39 VTAIL.n52 VTAIL.n51 185
R40 VTAIL.n53 VTAIL.n24 185
R41 VTAIL.n55 VTAIL.n54 185
R42 VTAIL.n22 VTAIL.n21 185
R43 VTAIL.n61 VTAIL.n60 185
R44 VTAIL.n63 VTAIL.n62 185
R45 VTAIL.n18 VTAIL.n17 185
R46 VTAIL.n69 VTAIL.n68 185
R47 VTAIL.n71 VTAIL.n70 185
R48 VTAIL.n14 VTAIL.n13 185
R49 VTAIL.n77 VTAIL.n76 185
R50 VTAIL.n79 VTAIL.n78 185
R51 VTAIL.n10 VTAIL.n9 185
R52 VTAIL.n85 VTAIL.n84 185
R53 VTAIL.n87 VTAIL.n86 185
R54 VTAIL.n6 VTAIL.n5 185
R55 VTAIL.n93 VTAIL.n92 185
R56 VTAIL.n95 VTAIL.n94 185
R57 VTAIL.n2 VTAIL.n1 185
R58 VTAIL.n101 VTAIL.n100 185
R59 VTAIL.n309 VTAIL.n308 185
R60 VTAIL.n210 VTAIL.n209 185
R61 VTAIL.n303 VTAIL.n302 185
R62 VTAIL.n301 VTAIL.n300 185
R63 VTAIL.n214 VTAIL.n213 185
R64 VTAIL.n295 VTAIL.n294 185
R65 VTAIL.n293 VTAIL.n292 185
R66 VTAIL.n218 VTAIL.n217 185
R67 VTAIL.n287 VTAIL.n286 185
R68 VTAIL.n285 VTAIL.n284 185
R69 VTAIL.n222 VTAIL.n221 185
R70 VTAIL.n279 VTAIL.n278 185
R71 VTAIL.n277 VTAIL.n276 185
R72 VTAIL.n226 VTAIL.n225 185
R73 VTAIL.n271 VTAIL.n270 185
R74 VTAIL.n269 VTAIL.n268 185
R75 VTAIL.n230 VTAIL.n229 185
R76 VTAIL.n234 VTAIL.n232 185
R77 VTAIL.n263 VTAIL.n262 185
R78 VTAIL.n261 VTAIL.n260 185
R79 VTAIL.n236 VTAIL.n235 185
R80 VTAIL.n255 VTAIL.n254 185
R81 VTAIL.n253 VTAIL.n252 185
R82 VTAIL.n240 VTAIL.n239 185
R83 VTAIL.n247 VTAIL.n246 185
R84 VTAIL.n245 VTAIL.n244 185
R85 VTAIL.n205 VTAIL.n204 185
R86 VTAIL.n106 VTAIL.n105 185
R87 VTAIL.n199 VTAIL.n198 185
R88 VTAIL.n197 VTAIL.n196 185
R89 VTAIL.n110 VTAIL.n109 185
R90 VTAIL.n191 VTAIL.n190 185
R91 VTAIL.n189 VTAIL.n188 185
R92 VTAIL.n114 VTAIL.n113 185
R93 VTAIL.n183 VTAIL.n182 185
R94 VTAIL.n181 VTAIL.n180 185
R95 VTAIL.n118 VTAIL.n117 185
R96 VTAIL.n175 VTAIL.n174 185
R97 VTAIL.n173 VTAIL.n172 185
R98 VTAIL.n122 VTAIL.n121 185
R99 VTAIL.n167 VTAIL.n166 185
R100 VTAIL.n165 VTAIL.n164 185
R101 VTAIL.n126 VTAIL.n125 185
R102 VTAIL.n130 VTAIL.n128 185
R103 VTAIL.n159 VTAIL.n158 185
R104 VTAIL.n157 VTAIL.n156 185
R105 VTAIL.n132 VTAIL.n131 185
R106 VTAIL.n151 VTAIL.n150 185
R107 VTAIL.n149 VTAIL.n148 185
R108 VTAIL.n136 VTAIL.n135 185
R109 VTAIL.n143 VTAIL.n142 185
R110 VTAIL.n141 VTAIL.n140 185
R111 VTAIL.n345 VTAIL.t0 149.524
R112 VTAIL.n33 VTAIL.t2 149.524
R113 VTAIL.n243 VTAIL.t1 149.524
R114 VTAIL.n139 VTAIL.t3 149.524
R115 VTAIL.n348 VTAIL.n347 104.615
R116 VTAIL.n348 VTAIL.n341 104.615
R117 VTAIL.n355 VTAIL.n341 104.615
R118 VTAIL.n356 VTAIL.n355 104.615
R119 VTAIL.n356 VTAIL.n337 104.615
R120 VTAIL.n364 VTAIL.n337 104.615
R121 VTAIL.n365 VTAIL.n364 104.615
R122 VTAIL.n366 VTAIL.n365 104.615
R123 VTAIL.n366 VTAIL.n333 104.615
R124 VTAIL.n373 VTAIL.n333 104.615
R125 VTAIL.n374 VTAIL.n373 104.615
R126 VTAIL.n374 VTAIL.n329 104.615
R127 VTAIL.n381 VTAIL.n329 104.615
R128 VTAIL.n382 VTAIL.n381 104.615
R129 VTAIL.n382 VTAIL.n325 104.615
R130 VTAIL.n389 VTAIL.n325 104.615
R131 VTAIL.n390 VTAIL.n389 104.615
R132 VTAIL.n390 VTAIL.n321 104.615
R133 VTAIL.n397 VTAIL.n321 104.615
R134 VTAIL.n398 VTAIL.n397 104.615
R135 VTAIL.n398 VTAIL.n317 104.615
R136 VTAIL.n405 VTAIL.n317 104.615
R137 VTAIL.n406 VTAIL.n405 104.615
R138 VTAIL.n406 VTAIL.n313 104.615
R139 VTAIL.n413 VTAIL.n313 104.615
R140 VTAIL.n36 VTAIL.n35 104.615
R141 VTAIL.n36 VTAIL.n29 104.615
R142 VTAIL.n43 VTAIL.n29 104.615
R143 VTAIL.n44 VTAIL.n43 104.615
R144 VTAIL.n44 VTAIL.n25 104.615
R145 VTAIL.n52 VTAIL.n25 104.615
R146 VTAIL.n53 VTAIL.n52 104.615
R147 VTAIL.n54 VTAIL.n53 104.615
R148 VTAIL.n54 VTAIL.n21 104.615
R149 VTAIL.n61 VTAIL.n21 104.615
R150 VTAIL.n62 VTAIL.n61 104.615
R151 VTAIL.n62 VTAIL.n17 104.615
R152 VTAIL.n69 VTAIL.n17 104.615
R153 VTAIL.n70 VTAIL.n69 104.615
R154 VTAIL.n70 VTAIL.n13 104.615
R155 VTAIL.n77 VTAIL.n13 104.615
R156 VTAIL.n78 VTAIL.n77 104.615
R157 VTAIL.n78 VTAIL.n9 104.615
R158 VTAIL.n85 VTAIL.n9 104.615
R159 VTAIL.n86 VTAIL.n85 104.615
R160 VTAIL.n86 VTAIL.n5 104.615
R161 VTAIL.n93 VTAIL.n5 104.615
R162 VTAIL.n94 VTAIL.n93 104.615
R163 VTAIL.n94 VTAIL.n1 104.615
R164 VTAIL.n101 VTAIL.n1 104.615
R165 VTAIL.n309 VTAIL.n209 104.615
R166 VTAIL.n302 VTAIL.n209 104.615
R167 VTAIL.n302 VTAIL.n301 104.615
R168 VTAIL.n301 VTAIL.n213 104.615
R169 VTAIL.n294 VTAIL.n213 104.615
R170 VTAIL.n294 VTAIL.n293 104.615
R171 VTAIL.n293 VTAIL.n217 104.615
R172 VTAIL.n286 VTAIL.n217 104.615
R173 VTAIL.n286 VTAIL.n285 104.615
R174 VTAIL.n285 VTAIL.n221 104.615
R175 VTAIL.n278 VTAIL.n221 104.615
R176 VTAIL.n278 VTAIL.n277 104.615
R177 VTAIL.n277 VTAIL.n225 104.615
R178 VTAIL.n270 VTAIL.n225 104.615
R179 VTAIL.n270 VTAIL.n269 104.615
R180 VTAIL.n269 VTAIL.n229 104.615
R181 VTAIL.n234 VTAIL.n229 104.615
R182 VTAIL.n262 VTAIL.n234 104.615
R183 VTAIL.n262 VTAIL.n261 104.615
R184 VTAIL.n261 VTAIL.n235 104.615
R185 VTAIL.n254 VTAIL.n235 104.615
R186 VTAIL.n254 VTAIL.n253 104.615
R187 VTAIL.n253 VTAIL.n239 104.615
R188 VTAIL.n246 VTAIL.n239 104.615
R189 VTAIL.n246 VTAIL.n245 104.615
R190 VTAIL.n205 VTAIL.n105 104.615
R191 VTAIL.n198 VTAIL.n105 104.615
R192 VTAIL.n198 VTAIL.n197 104.615
R193 VTAIL.n197 VTAIL.n109 104.615
R194 VTAIL.n190 VTAIL.n109 104.615
R195 VTAIL.n190 VTAIL.n189 104.615
R196 VTAIL.n189 VTAIL.n113 104.615
R197 VTAIL.n182 VTAIL.n113 104.615
R198 VTAIL.n182 VTAIL.n181 104.615
R199 VTAIL.n181 VTAIL.n117 104.615
R200 VTAIL.n174 VTAIL.n117 104.615
R201 VTAIL.n174 VTAIL.n173 104.615
R202 VTAIL.n173 VTAIL.n121 104.615
R203 VTAIL.n166 VTAIL.n121 104.615
R204 VTAIL.n166 VTAIL.n165 104.615
R205 VTAIL.n165 VTAIL.n125 104.615
R206 VTAIL.n130 VTAIL.n125 104.615
R207 VTAIL.n158 VTAIL.n130 104.615
R208 VTAIL.n158 VTAIL.n157 104.615
R209 VTAIL.n157 VTAIL.n131 104.615
R210 VTAIL.n150 VTAIL.n131 104.615
R211 VTAIL.n150 VTAIL.n149 104.615
R212 VTAIL.n149 VTAIL.n135 104.615
R213 VTAIL.n142 VTAIL.n135 104.615
R214 VTAIL.n142 VTAIL.n141 104.615
R215 VTAIL.n347 VTAIL.t0 52.3082
R216 VTAIL.n35 VTAIL.t2 52.3082
R217 VTAIL.n245 VTAIL.t1 52.3082
R218 VTAIL.n141 VTAIL.t3 52.3082
R219 VTAIL.n415 VTAIL.n414 35.2884
R220 VTAIL.n103 VTAIL.n102 35.2884
R221 VTAIL.n311 VTAIL.n310 35.2884
R222 VTAIL.n207 VTAIL.n206 35.2884
R223 VTAIL.n207 VTAIL.n103 33.091
R224 VTAIL.n415 VTAIL.n311 30.8238
R225 VTAIL.n367 VTAIL.n334 13.1884
R226 VTAIL.n55 VTAIL.n22 13.1884
R227 VTAIL.n232 VTAIL.n230 13.1884
R228 VTAIL.n128 VTAIL.n126 13.1884
R229 VTAIL.n368 VTAIL.n336 12.8005
R230 VTAIL.n372 VTAIL.n371 12.8005
R231 VTAIL.n412 VTAIL.n312 12.8005
R232 VTAIL.n56 VTAIL.n24 12.8005
R233 VTAIL.n60 VTAIL.n59 12.8005
R234 VTAIL.n100 VTAIL.n0 12.8005
R235 VTAIL.n308 VTAIL.n208 12.8005
R236 VTAIL.n268 VTAIL.n267 12.8005
R237 VTAIL.n264 VTAIL.n263 12.8005
R238 VTAIL.n204 VTAIL.n104 12.8005
R239 VTAIL.n164 VTAIL.n163 12.8005
R240 VTAIL.n160 VTAIL.n159 12.8005
R241 VTAIL.n363 VTAIL.n362 12.0247
R242 VTAIL.n375 VTAIL.n332 12.0247
R243 VTAIL.n411 VTAIL.n314 12.0247
R244 VTAIL.n51 VTAIL.n50 12.0247
R245 VTAIL.n63 VTAIL.n20 12.0247
R246 VTAIL.n99 VTAIL.n2 12.0247
R247 VTAIL.n307 VTAIL.n210 12.0247
R248 VTAIL.n271 VTAIL.n228 12.0247
R249 VTAIL.n260 VTAIL.n233 12.0247
R250 VTAIL.n203 VTAIL.n106 12.0247
R251 VTAIL.n167 VTAIL.n124 12.0247
R252 VTAIL.n156 VTAIL.n129 12.0247
R253 VTAIL.n361 VTAIL.n338 11.249
R254 VTAIL.n376 VTAIL.n330 11.249
R255 VTAIL.n408 VTAIL.n407 11.249
R256 VTAIL.n49 VTAIL.n26 11.249
R257 VTAIL.n64 VTAIL.n18 11.249
R258 VTAIL.n96 VTAIL.n95 11.249
R259 VTAIL.n304 VTAIL.n303 11.249
R260 VTAIL.n272 VTAIL.n226 11.249
R261 VTAIL.n259 VTAIL.n236 11.249
R262 VTAIL.n200 VTAIL.n199 11.249
R263 VTAIL.n168 VTAIL.n122 11.249
R264 VTAIL.n155 VTAIL.n132 11.249
R265 VTAIL.n358 VTAIL.n357 10.4732
R266 VTAIL.n380 VTAIL.n379 10.4732
R267 VTAIL.n404 VTAIL.n316 10.4732
R268 VTAIL.n46 VTAIL.n45 10.4732
R269 VTAIL.n68 VTAIL.n67 10.4732
R270 VTAIL.n92 VTAIL.n4 10.4732
R271 VTAIL.n300 VTAIL.n212 10.4732
R272 VTAIL.n276 VTAIL.n275 10.4732
R273 VTAIL.n256 VTAIL.n255 10.4732
R274 VTAIL.n196 VTAIL.n108 10.4732
R275 VTAIL.n172 VTAIL.n171 10.4732
R276 VTAIL.n152 VTAIL.n151 10.4732
R277 VTAIL.n346 VTAIL.n345 10.2747
R278 VTAIL.n34 VTAIL.n33 10.2747
R279 VTAIL.n244 VTAIL.n243 10.2747
R280 VTAIL.n140 VTAIL.n139 10.2747
R281 VTAIL.n354 VTAIL.n340 9.69747
R282 VTAIL.n383 VTAIL.n328 9.69747
R283 VTAIL.n403 VTAIL.n318 9.69747
R284 VTAIL.n42 VTAIL.n28 9.69747
R285 VTAIL.n71 VTAIL.n16 9.69747
R286 VTAIL.n91 VTAIL.n6 9.69747
R287 VTAIL.n299 VTAIL.n214 9.69747
R288 VTAIL.n279 VTAIL.n224 9.69747
R289 VTAIL.n252 VTAIL.n238 9.69747
R290 VTAIL.n195 VTAIL.n110 9.69747
R291 VTAIL.n175 VTAIL.n120 9.69747
R292 VTAIL.n148 VTAIL.n134 9.69747
R293 VTAIL.n410 VTAIL.n312 9.45567
R294 VTAIL.n98 VTAIL.n0 9.45567
R295 VTAIL.n306 VTAIL.n208 9.45567
R296 VTAIL.n202 VTAIL.n104 9.45567
R297 VTAIL.n393 VTAIL.n392 9.3005
R298 VTAIL.n395 VTAIL.n394 9.3005
R299 VTAIL.n320 VTAIL.n319 9.3005
R300 VTAIL.n401 VTAIL.n400 9.3005
R301 VTAIL.n403 VTAIL.n402 9.3005
R302 VTAIL.n316 VTAIL.n315 9.3005
R303 VTAIL.n409 VTAIL.n408 9.3005
R304 VTAIL.n411 VTAIL.n410 9.3005
R305 VTAIL.n387 VTAIL.n386 9.3005
R306 VTAIL.n385 VTAIL.n384 9.3005
R307 VTAIL.n328 VTAIL.n327 9.3005
R308 VTAIL.n379 VTAIL.n378 9.3005
R309 VTAIL.n377 VTAIL.n376 9.3005
R310 VTAIL.n332 VTAIL.n331 9.3005
R311 VTAIL.n371 VTAIL.n370 9.3005
R312 VTAIL.n344 VTAIL.n343 9.3005
R313 VTAIL.n351 VTAIL.n350 9.3005
R314 VTAIL.n353 VTAIL.n352 9.3005
R315 VTAIL.n340 VTAIL.n339 9.3005
R316 VTAIL.n359 VTAIL.n358 9.3005
R317 VTAIL.n361 VTAIL.n360 9.3005
R318 VTAIL.n362 VTAIL.n335 9.3005
R319 VTAIL.n369 VTAIL.n368 9.3005
R320 VTAIL.n324 VTAIL.n323 9.3005
R321 VTAIL.n81 VTAIL.n80 9.3005
R322 VTAIL.n83 VTAIL.n82 9.3005
R323 VTAIL.n8 VTAIL.n7 9.3005
R324 VTAIL.n89 VTAIL.n88 9.3005
R325 VTAIL.n91 VTAIL.n90 9.3005
R326 VTAIL.n4 VTAIL.n3 9.3005
R327 VTAIL.n97 VTAIL.n96 9.3005
R328 VTAIL.n99 VTAIL.n98 9.3005
R329 VTAIL.n75 VTAIL.n74 9.3005
R330 VTAIL.n73 VTAIL.n72 9.3005
R331 VTAIL.n16 VTAIL.n15 9.3005
R332 VTAIL.n67 VTAIL.n66 9.3005
R333 VTAIL.n65 VTAIL.n64 9.3005
R334 VTAIL.n20 VTAIL.n19 9.3005
R335 VTAIL.n59 VTAIL.n58 9.3005
R336 VTAIL.n32 VTAIL.n31 9.3005
R337 VTAIL.n39 VTAIL.n38 9.3005
R338 VTAIL.n41 VTAIL.n40 9.3005
R339 VTAIL.n28 VTAIL.n27 9.3005
R340 VTAIL.n47 VTAIL.n46 9.3005
R341 VTAIL.n49 VTAIL.n48 9.3005
R342 VTAIL.n50 VTAIL.n23 9.3005
R343 VTAIL.n57 VTAIL.n56 9.3005
R344 VTAIL.n12 VTAIL.n11 9.3005
R345 VTAIL.n307 VTAIL.n306 9.3005
R346 VTAIL.n305 VTAIL.n304 9.3005
R347 VTAIL.n212 VTAIL.n211 9.3005
R348 VTAIL.n299 VTAIL.n298 9.3005
R349 VTAIL.n297 VTAIL.n296 9.3005
R350 VTAIL.n216 VTAIL.n215 9.3005
R351 VTAIL.n291 VTAIL.n290 9.3005
R352 VTAIL.n289 VTAIL.n288 9.3005
R353 VTAIL.n220 VTAIL.n219 9.3005
R354 VTAIL.n283 VTAIL.n282 9.3005
R355 VTAIL.n281 VTAIL.n280 9.3005
R356 VTAIL.n224 VTAIL.n223 9.3005
R357 VTAIL.n275 VTAIL.n274 9.3005
R358 VTAIL.n273 VTAIL.n272 9.3005
R359 VTAIL.n228 VTAIL.n227 9.3005
R360 VTAIL.n267 VTAIL.n266 9.3005
R361 VTAIL.n265 VTAIL.n264 9.3005
R362 VTAIL.n233 VTAIL.n231 9.3005
R363 VTAIL.n259 VTAIL.n258 9.3005
R364 VTAIL.n257 VTAIL.n256 9.3005
R365 VTAIL.n238 VTAIL.n237 9.3005
R366 VTAIL.n251 VTAIL.n250 9.3005
R367 VTAIL.n249 VTAIL.n248 9.3005
R368 VTAIL.n242 VTAIL.n241 9.3005
R369 VTAIL.n138 VTAIL.n137 9.3005
R370 VTAIL.n145 VTAIL.n144 9.3005
R371 VTAIL.n147 VTAIL.n146 9.3005
R372 VTAIL.n134 VTAIL.n133 9.3005
R373 VTAIL.n153 VTAIL.n152 9.3005
R374 VTAIL.n155 VTAIL.n154 9.3005
R375 VTAIL.n129 VTAIL.n127 9.3005
R376 VTAIL.n161 VTAIL.n160 9.3005
R377 VTAIL.n187 VTAIL.n186 9.3005
R378 VTAIL.n112 VTAIL.n111 9.3005
R379 VTAIL.n193 VTAIL.n192 9.3005
R380 VTAIL.n195 VTAIL.n194 9.3005
R381 VTAIL.n108 VTAIL.n107 9.3005
R382 VTAIL.n201 VTAIL.n200 9.3005
R383 VTAIL.n203 VTAIL.n202 9.3005
R384 VTAIL.n185 VTAIL.n184 9.3005
R385 VTAIL.n116 VTAIL.n115 9.3005
R386 VTAIL.n179 VTAIL.n178 9.3005
R387 VTAIL.n177 VTAIL.n176 9.3005
R388 VTAIL.n120 VTAIL.n119 9.3005
R389 VTAIL.n171 VTAIL.n170 9.3005
R390 VTAIL.n169 VTAIL.n168 9.3005
R391 VTAIL.n124 VTAIL.n123 9.3005
R392 VTAIL.n163 VTAIL.n162 9.3005
R393 VTAIL.n353 VTAIL.n342 8.92171
R394 VTAIL.n384 VTAIL.n326 8.92171
R395 VTAIL.n400 VTAIL.n399 8.92171
R396 VTAIL.n41 VTAIL.n30 8.92171
R397 VTAIL.n72 VTAIL.n14 8.92171
R398 VTAIL.n88 VTAIL.n87 8.92171
R399 VTAIL.n296 VTAIL.n295 8.92171
R400 VTAIL.n280 VTAIL.n222 8.92171
R401 VTAIL.n251 VTAIL.n240 8.92171
R402 VTAIL.n192 VTAIL.n191 8.92171
R403 VTAIL.n176 VTAIL.n118 8.92171
R404 VTAIL.n147 VTAIL.n136 8.92171
R405 VTAIL.n350 VTAIL.n349 8.14595
R406 VTAIL.n388 VTAIL.n387 8.14595
R407 VTAIL.n396 VTAIL.n320 8.14595
R408 VTAIL.n38 VTAIL.n37 8.14595
R409 VTAIL.n76 VTAIL.n75 8.14595
R410 VTAIL.n84 VTAIL.n8 8.14595
R411 VTAIL.n292 VTAIL.n216 8.14595
R412 VTAIL.n284 VTAIL.n283 8.14595
R413 VTAIL.n248 VTAIL.n247 8.14595
R414 VTAIL.n188 VTAIL.n112 8.14595
R415 VTAIL.n180 VTAIL.n179 8.14595
R416 VTAIL.n144 VTAIL.n143 8.14595
R417 VTAIL.n346 VTAIL.n344 7.3702
R418 VTAIL.n391 VTAIL.n324 7.3702
R419 VTAIL.n395 VTAIL.n322 7.3702
R420 VTAIL.n34 VTAIL.n32 7.3702
R421 VTAIL.n79 VTAIL.n12 7.3702
R422 VTAIL.n83 VTAIL.n10 7.3702
R423 VTAIL.n291 VTAIL.n218 7.3702
R424 VTAIL.n287 VTAIL.n220 7.3702
R425 VTAIL.n244 VTAIL.n242 7.3702
R426 VTAIL.n187 VTAIL.n114 7.3702
R427 VTAIL.n183 VTAIL.n116 7.3702
R428 VTAIL.n140 VTAIL.n138 7.3702
R429 VTAIL.n392 VTAIL.n391 6.59444
R430 VTAIL.n392 VTAIL.n322 6.59444
R431 VTAIL.n80 VTAIL.n79 6.59444
R432 VTAIL.n80 VTAIL.n10 6.59444
R433 VTAIL.n288 VTAIL.n218 6.59444
R434 VTAIL.n288 VTAIL.n287 6.59444
R435 VTAIL.n184 VTAIL.n114 6.59444
R436 VTAIL.n184 VTAIL.n183 6.59444
R437 VTAIL.n349 VTAIL.n344 5.81868
R438 VTAIL.n388 VTAIL.n324 5.81868
R439 VTAIL.n396 VTAIL.n395 5.81868
R440 VTAIL.n37 VTAIL.n32 5.81868
R441 VTAIL.n76 VTAIL.n12 5.81868
R442 VTAIL.n84 VTAIL.n83 5.81868
R443 VTAIL.n292 VTAIL.n291 5.81868
R444 VTAIL.n284 VTAIL.n220 5.81868
R445 VTAIL.n247 VTAIL.n242 5.81868
R446 VTAIL.n188 VTAIL.n187 5.81868
R447 VTAIL.n180 VTAIL.n116 5.81868
R448 VTAIL.n143 VTAIL.n138 5.81868
R449 VTAIL.n350 VTAIL.n342 5.04292
R450 VTAIL.n387 VTAIL.n326 5.04292
R451 VTAIL.n399 VTAIL.n320 5.04292
R452 VTAIL.n38 VTAIL.n30 5.04292
R453 VTAIL.n75 VTAIL.n14 5.04292
R454 VTAIL.n87 VTAIL.n8 5.04292
R455 VTAIL.n295 VTAIL.n216 5.04292
R456 VTAIL.n283 VTAIL.n222 5.04292
R457 VTAIL.n248 VTAIL.n240 5.04292
R458 VTAIL.n191 VTAIL.n112 5.04292
R459 VTAIL.n179 VTAIL.n118 5.04292
R460 VTAIL.n144 VTAIL.n136 5.04292
R461 VTAIL.n354 VTAIL.n353 4.26717
R462 VTAIL.n384 VTAIL.n383 4.26717
R463 VTAIL.n400 VTAIL.n318 4.26717
R464 VTAIL.n42 VTAIL.n41 4.26717
R465 VTAIL.n72 VTAIL.n71 4.26717
R466 VTAIL.n88 VTAIL.n6 4.26717
R467 VTAIL.n296 VTAIL.n214 4.26717
R468 VTAIL.n280 VTAIL.n279 4.26717
R469 VTAIL.n252 VTAIL.n251 4.26717
R470 VTAIL.n192 VTAIL.n110 4.26717
R471 VTAIL.n176 VTAIL.n175 4.26717
R472 VTAIL.n148 VTAIL.n147 4.26717
R473 VTAIL.n357 VTAIL.n340 3.49141
R474 VTAIL.n380 VTAIL.n328 3.49141
R475 VTAIL.n404 VTAIL.n403 3.49141
R476 VTAIL.n45 VTAIL.n28 3.49141
R477 VTAIL.n68 VTAIL.n16 3.49141
R478 VTAIL.n92 VTAIL.n91 3.49141
R479 VTAIL.n300 VTAIL.n299 3.49141
R480 VTAIL.n276 VTAIL.n224 3.49141
R481 VTAIL.n255 VTAIL.n238 3.49141
R482 VTAIL.n196 VTAIL.n195 3.49141
R483 VTAIL.n172 VTAIL.n120 3.49141
R484 VTAIL.n151 VTAIL.n134 3.49141
R485 VTAIL.n345 VTAIL.n343 2.84303
R486 VTAIL.n33 VTAIL.n31 2.84303
R487 VTAIL.n243 VTAIL.n241 2.84303
R488 VTAIL.n139 VTAIL.n137 2.84303
R489 VTAIL.n358 VTAIL.n338 2.71565
R490 VTAIL.n379 VTAIL.n330 2.71565
R491 VTAIL.n407 VTAIL.n316 2.71565
R492 VTAIL.n46 VTAIL.n26 2.71565
R493 VTAIL.n67 VTAIL.n18 2.71565
R494 VTAIL.n95 VTAIL.n4 2.71565
R495 VTAIL.n303 VTAIL.n212 2.71565
R496 VTAIL.n275 VTAIL.n226 2.71565
R497 VTAIL.n256 VTAIL.n236 2.71565
R498 VTAIL.n199 VTAIL.n108 2.71565
R499 VTAIL.n171 VTAIL.n122 2.71565
R500 VTAIL.n152 VTAIL.n132 2.71565
R501 VTAIL.n363 VTAIL.n361 1.93989
R502 VTAIL.n376 VTAIL.n375 1.93989
R503 VTAIL.n408 VTAIL.n314 1.93989
R504 VTAIL.n51 VTAIL.n49 1.93989
R505 VTAIL.n64 VTAIL.n63 1.93989
R506 VTAIL.n96 VTAIL.n2 1.93989
R507 VTAIL.n304 VTAIL.n210 1.93989
R508 VTAIL.n272 VTAIL.n271 1.93989
R509 VTAIL.n260 VTAIL.n259 1.93989
R510 VTAIL.n200 VTAIL.n106 1.93989
R511 VTAIL.n168 VTAIL.n167 1.93989
R512 VTAIL.n156 VTAIL.n155 1.93989
R513 VTAIL.n311 VTAIL.n207 1.60395
R514 VTAIL.n362 VTAIL.n336 1.16414
R515 VTAIL.n372 VTAIL.n332 1.16414
R516 VTAIL.n412 VTAIL.n411 1.16414
R517 VTAIL.n50 VTAIL.n24 1.16414
R518 VTAIL.n60 VTAIL.n20 1.16414
R519 VTAIL.n100 VTAIL.n99 1.16414
R520 VTAIL.n308 VTAIL.n307 1.16414
R521 VTAIL.n268 VTAIL.n228 1.16414
R522 VTAIL.n263 VTAIL.n233 1.16414
R523 VTAIL.n204 VTAIL.n203 1.16414
R524 VTAIL.n164 VTAIL.n124 1.16414
R525 VTAIL.n159 VTAIL.n129 1.16414
R526 VTAIL VTAIL.n103 1.09533
R527 VTAIL VTAIL.n415 0.509121
R528 VTAIL.n368 VTAIL.n367 0.388379
R529 VTAIL.n371 VTAIL.n334 0.388379
R530 VTAIL.n414 VTAIL.n312 0.388379
R531 VTAIL.n56 VTAIL.n55 0.388379
R532 VTAIL.n59 VTAIL.n22 0.388379
R533 VTAIL.n102 VTAIL.n0 0.388379
R534 VTAIL.n310 VTAIL.n208 0.388379
R535 VTAIL.n267 VTAIL.n230 0.388379
R536 VTAIL.n264 VTAIL.n232 0.388379
R537 VTAIL.n206 VTAIL.n104 0.388379
R538 VTAIL.n163 VTAIL.n126 0.388379
R539 VTAIL.n160 VTAIL.n128 0.388379
R540 VTAIL.n351 VTAIL.n343 0.155672
R541 VTAIL.n352 VTAIL.n351 0.155672
R542 VTAIL.n352 VTAIL.n339 0.155672
R543 VTAIL.n359 VTAIL.n339 0.155672
R544 VTAIL.n360 VTAIL.n359 0.155672
R545 VTAIL.n360 VTAIL.n335 0.155672
R546 VTAIL.n369 VTAIL.n335 0.155672
R547 VTAIL.n370 VTAIL.n369 0.155672
R548 VTAIL.n370 VTAIL.n331 0.155672
R549 VTAIL.n377 VTAIL.n331 0.155672
R550 VTAIL.n378 VTAIL.n377 0.155672
R551 VTAIL.n378 VTAIL.n327 0.155672
R552 VTAIL.n385 VTAIL.n327 0.155672
R553 VTAIL.n386 VTAIL.n385 0.155672
R554 VTAIL.n386 VTAIL.n323 0.155672
R555 VTAIL.n393 VTAIL.n323 0.155672
R556 VTAIL.n394 VTAIL.n393 0.155672
R557 VTAIL.n394 VTAIL.n319 0.155672
R558 VTAIL.n401 VTAIL.n319 0.155672
R559 VTAIL.n402 VTAIL.n401 0.155672
R560 VTAIL.n402 VTAIL.n315 0.155672
R561 VTAIL.n409 VTAIL.n315 0.155672
R562 VTAIL.n410 VTAIL.n409 0.155672
R563 VTAIL.n39 VTAIL.n31 0.155672
R564 VTAIL.n40 VTAIL.n39 0.155672
R565 VTAIL.n40 VTAIL.n27 0.155672
R566 VTAIL.n47 VTAIL.n27 0.155672
R567 VTAIL.n48 VTAIL.n47 0.155672
R568 VTAIL.n48 VTAIL.n23 0.155672
R569 VTAIL.n57 VTAIL.n23 0.155672
R570 VTAIL.n58 VTAIL.n57 0.155672
R571 VTAIL.n58 VTAIL.n19 0.155672
R572 VTAIL.n65 VTAIL.n19 0.155672
R573 VTAIL.n66 VTAIL.n65 0.155672
R574 VTAIL.n66 VTAIL.n15 0.155672
R575 VTAIL.n73 VTAIL.n15 0.155672
R576 VTAIL.n74 VTAIL.n73 0.155672
R577 VTAIL.n74 VTAIL.n11 0.155672
R578 VTAIL.n81 VTAIL.n11 0.155672
R579 VTAIL.n82 VTAIL.n81 0.155672
R580 VTAIL.n82 VTAIL.n7 0.155672
R581 VTAIL.n89 VTAIL.n7 0.155672
R582 VTAIL.n90 VTAIL.n89 0.155672
R583 VTAIL.n90 VTAIL.n3 0.155672
R584 VTAIL.n97 VTAIL.n3 0.155672
R585 VTAIL.n98 VTAIL.n97 0.155672
R586 VTAIL.n306 VTAIL.n305 0.155672
R587 VTAIL.n305 VTAIL.n211 0.155672
R588 VTAIL.n298 VTAIL.n211 0.155672
R589 VTAIL.n298 VTAIL.n297 0.155672
R590 VTAIL.n297 VTAIL.n215 0.155672
R591 VTAIL.n290 VTAIL.n215 0.155672
R592 VTAIL.n290 VTAIL.n289 0.155672
R593 VTAIL.n289 VTAIL.n219 0.155672
R594 VTAIL.n282 VTAIL.n219 0.155672
R595 VTAIL.n282 VTAIL.n281 0.155672
R596 VTAIL.n281 VTAIL.n223 0.155672
R597 VTAIL.n274 VTAIL.n223 0.155672
R598 VTAIL.n274 VTAIL.n273 0.155672
R599 VTAIL.n273 VTAIL.n227 0.155672
R600 VTAIL.n266 VTAIL.n227 0.155672
R601 VTAIL.n266 VTAIL.n265 0.155672
R602 VTAIL.n265 VTAIL.n231 0.155672
R603 VTAIL.n258 VTAIL.n231 0.155672
R604 VTAIL.n258 VTAIL.n257 0.155672
R605 VTAIL.n257 VTAIL.n237 0.155672
R606 VTAIL.n250 VTAIL.n237 0.155672
R607 VTAIL.n250 VTAIL.n249 0.155672
R608 VTAIL.n249 VTAIL.n241 0.155672
R609 VTAIL.n202 VTAIL.n201 0.155672
R610 VTAIL.n201 VTAIL.n107 0.155672
R611 VTAIL.n194 VTAIL.n107 0.155672
R612 VTAIL.n194 VTAIL.n193 0.155672
R613 VTAIL.n193 VTAIL.n111 0.155672
R614 VTAIL.n186 VTAIL.n111 0.155672
R615 VTAIL.n186 VTAIL.n185 0.155672
R616 VTAIL.n185 VTAIL.n115 0.155672
R617 VTAIL.n178 VTAIL.n115 0.155672
R618 VTAIL.n178 VTAIL.n177 0.155672
R619 VTAIL.n177 VTAIL.n119 0.155672
R620 VTAIL.n170 VTAIL.n119 0.155672
R621 VTAIL.n170 VTAIL.n169 0.155672
R622 VTAIL.n169 VTAIL.n123 0.155672
R623 VTAIL.n162 VTAIL.n123 0.155672
R624 VTAIL.n162 VTAIL.n161 0.155672
R625 VTAIL.n161 VTAIL.n127 0.155672
R626 VTAIL.n154 VTAIL.n127 0.155672
R627 VTAIL.n154 VTAIL.n153 0.155672
R628 VTAIL.n153 VTAIL.n133 0.155672
R629 VTAIL.n146 VTAIL.n133 0.155672
R630 VTAIL.n146 VTAIL.n145 0.155672
R631 VTAIL.n145 VTAIL.n137 0.155672
R632 VDD1.n102 VDD1.n101 289.615
R633 VDD1.n205 VDD1.n204 289.615
R634 VDD1.n101 VDD1.n100 185
R635 VDD1.n2 VDD1.n1 185
R636 VDD1.n95 VDD1.n94 185
R637 VDD1.n93 VDD1.n92 185
R638 VDD1.n6 VDD1.n5 185
R639 VDD1.n87 VDD1.n86 185
R640 VDD1.n85 VDD1.n84 185
R641 VDD1.n10 VDD1.n9 185
R642 VDD1.n79 VDD1.n78 185
R643 VDD1.n77 VDD1.n76 185
R644 VDD1.n14 VDD1.n13 185
R645 VDD1.n71 VDD1.n70 185
R646 VDD1.n69 VDD1.n68 185
R647 VDD1.n18 VDD1.n17 185
R648 VDD1.n63 VDD1.n62 185
R649 VDD1.n61 VDD1.n60 185
R650 VDD1.n22 VDD1.n21 185
R651 VDD1.n26 VDD1.n24 185
R652 VDD1.n55 VDD1.n54 185
R653 VDD1.n53 VDD1.n52 185
R654 VDD1.n28 VDD1.n27 185
R655 VDD1.n47 VDD1.n46 185
R656 VDD1.n45 VDD1.n44 185
R657 VDD1.n32 VDD1.n31 185
R658 VDD1.n39 VDD1.n38 185
R659 VDD1.n37 VDD1.n36 185
R660 VDD1.n138 VDD1.n137 185
R661 VDD1.n140 VDD1.n139 185
R662 VDD1.n133 VDD1.n132 185
R663 VDD1.n146 VDD1.n145 185
R664 VDD1.n148 VDD1.n147 185
R665 VDD1.n129 VDD1.n128 185
R666 VDD1.n155 VDD1.n154 185
R667 VDD1.n156 VDD1.n127 185
R668 VDD1.n158 VDD1.n157 185
R669 VDD1.n125 VDD1.n124 185
R670 VDD1.n164 VDD1.n163 185
R671 VDD1.n166 VDD1.n165 185
R672 VDD1.n121 VDD1.n120 185
R673 VDD1.n172 VDD1.n171 185
R674 VDD1.n174 VDD1.n173 185
R675 VDD1.n117 VDD1.n116 185
R676 VDD1.n180 VDD1.n179 185
R677 VDD1.n182 VDD1.n181 185
R678 VDD1.n113 VDD1.n112 185
R679 VDD1.n188 VDD1.n187 185
R680 VDD1.n190 VDD1.n189 185
R681 VDD1.n109 VDD1.n108 185
R682 VDD1.n196 VDD1.n195 185
R683 VDD1.n198 VDD1.n197 185
R684 VDD1.n105 VDD1.n104 185
R685 VDD1.n204 VDD1.n203 185
R686 VDD1.n35 VDD1.t1 149.524
R687 VDD1.n136 VDD1.t0 149.524
R688 VDD1.n101 VDD1.n1 104.615
R689 VDD1.n94 VDD1.n1 104.615
R690 VDD1.n94 VDD1.n93 104.615
R691 VDD1.n93 VDD1.n5 104.615
R692 VDD1.n86 VDD1.n5 104.615
R693 VDD1.n86 VDD1.n85 104.615
R694 VDD1.n85 VDD1.n9 104.615
R695 VDD1.n78 VDD1.n9 104.615
R696 VDD1.n78 VDD1.n77 104.615
R697 VDD1.n77 VDD1.n13 104.615
R698 VDD1.n70 VDD1.n13 104.615
R699 VDD1.n70 VDD1.n69 104.615
R700 VDD1.n69 VDD1.n17 104.615
R701 VDD1.n62 VDD1.n17 104.615
R702 VDD1.n62 VDD1.n61 104.615
R703 VDD1.n61 VDD1.n21 104.615
R704 VDD1.n26 VDD1.n21 104.615
R705 VDD1.n54 VDD1.n26 104.615
R706 VDD1.n54 VDD1.n53 104.615
R707 VDD1.n53 VDD1.n27 104.615
R708 VDD1.n46 VDD1.n27 104.615
R709 VDD1.n46 VDD1.n45 104.615
R710 VDD1.n45 VDD1.n31 104.615
R711 VDD1.n38 VDD1.n31 104.615
R712 VDD1.n38 VDD1.n37 104.615
R713 VDD1.n139 VDD1.n138 104.615
R714 VDD1.n139 VDD1.n132 104.615
R715 VDD1.n146 VDD1.n132 104.615
R716 VDD1.n147 VDD1.n146 104.615
R717 VDD1.n147 VDD1.n128 104.615
R718 VDD1.n155 VDD1.n128 104.615
R719 VDD1.n156 VDD1.n155 104.615
R720 VDD1.n157 VDD1.n156 104.615
R721 VDD1.n157 VDD1.n124 104.615
R722 VDD1.n164 VDD1.n124 104.615
R723 VDD1.n165 VDD1.n164 104.615
R724 VDD1.n165 VDD1.n120 104.615
R725 VDD1.n172 VDD1.n120 104.615
R726 VDD1.n173 VDD1.n172 104.615
R727 VDD1.n173 VDD1.n116 104.615
R728 VDD1.n180 VDD1.n116 104.615
R729 VDD1.n181 VDD1.n180 104.615
R730 VDD1.n181 VDD1.n112 104.615
R731 VDD1.n188 VDD1.n112 104.615
R732 VDD1.n189 VDD1.n188 104.615
R733 VDD1.n189 VDD1.n108 104.615
R734 VDD1.n196 VDD1.n108 104.615
R735 VDD1.n197 VDD1.n196 104.615
R736 VDD1.n197 VDD1.n104 104.615
R737 VDD1.n204 VDD1.n104 104.615
R738 VDD1 VDD1.n205 97.4424
R739 VDD1 VDD1.n102 52.5922
R740 VDD1.n37 VDD1.t1 52.3082
R741 VDD1.n138 VDD1.t0 52.3082
R742 VDD1.n24 VDD1.n22 13.1884
R743 VDD1.n158 VDD1.n125 13.1884
R744 VDD1.n100 VDD1.n0 12.8005
R745 VDD1.n60 VDD1.n59 12.8005
R746 VDD1.n56 VDD1.n55 12.8005
R747 VDD1.n159 VDD1.n127 12.8005
R748 VDD1.n163 VDD1.n162 12.8005
R749 VDD1.n203 VDD1.n103 12.8005
R750 VDD1.n99 VDD1.n2 12.0247
R751 VDD1.n63 VDD1.n20 12.0247
R752 VDD1.n52 VDD1.n25 12.0247
R753 VDD1.n154 VDD1.n153 12.0247
R754 VDD1.n166 VDD1.n123 12.0247
R755 VDD1.n202 VDD1.n105 12.0247
R756 VDD1.n96 VDD1.n95 11.249
R757 VDD1.n64 VDD1.n18 11.249
R758 VDD1.n51 VDD1.n28 11.249
R759 VDD1.n152 VDD1.n129 11.249
R760 VDD1.n167 VDD1.n121 11.249
R761 VDD1.n199 VDD1.n198 11.249
R762 VDD1.n92 VDD1.n4 10.4732
R763 VDD1.n68 VDD1.n67 10.4732
R764 VDD1.n48 VDD1.n47 10.4732
R765 VDD1.n149 VDD1.n148 10.4732
R766 VDD1.n171 VDD1.n170 10.4732
R767 VDD1.n195 VDD1.n107 10.4732
R768 VDD1.n36 VDD1.n35 10.2747
R769 VDD1.n137 VDD1.n136 10.2747
R770 VDD1.n91 VDD1.n6 9.69747
R771 VDD1.n71 VDD1.n16 9.69747
R772 VDD1.n44 VDD1.n30 9.69747
R773 VDD1.n145 VDD1.n131 9.69747
R774 VDD1.n174 VDD1.n119 9.69747
R775 VDD1.n194 VDD1.n109 9.69747
R776 VDD1.n98 VDD1.n0 9.45567
R777 VDD1.n201 VDD1.n103 9.45567
R778 VDD1.n99 VDD1.n98 9.3005
R779 VDD1.n97 VDD1.n96 9.3005
R780 VDD1.n4 VDD1.n3 9.3005
R781 VDD1.n91 VDD1.n90 9.3005
R782 VDD1.n89 VDD1.n88 9.3005
R783 VDD1.n8 VDD1.n7 9.3005
R784 VDD1.n83 VDD1.n82 9.3005
R785 VDD1.n81 VDD1.n80 9.3005
R786 VDD1.n12 VDD1.n11 9.3005
R787 VDD1.n75 VDD1.n74 9.3005
R788 VDD1.n73 VDD1.n72 9.3005
R789 VDD1.n16 VDD1.n15 9.3005
R790 VDD1.n67 VDD1.n66 9.3005
R791 VDD1.n65 VDD1.n64 9.3005
R792 VDD1.n20 VDD1.n19 9.3005
R793 VDD1.n59 VDD1.n58 9.3005
R794 VDD1.n57 VDD1.n56 9.3005
R795 VDD1.n25 VDD1.n23 9.3005
R796 VDD1.n51 VDD1.n50 9.3005
R797 VDD1.n49 VDD1.n48 9.3005
R798 VDD1.n30 VDD1.n29 9.3005
R799 VDD1.n43 VDD1.n42 9.3005
R800 VDD1.n41 VDD1.n40 9.3005
R801 VDD1.n34 VDD1.n33 9.3005
R802 VDD1.n184 VDD1.n183 9.3005
R803 VDD1.n186 VDD1.n185 9.3005
R804 VDD1.n111 VDD1.n110 9.3005
R805 VDD1.n192 VDD1.n191 9.3005
R806 VDD1.n194 VDD1.n193 9.3005
R807 VDD1.n107 VDD1.n106 9.3005
R808 VDD1.n200 VDD1.n199 9.3005
R809 VDD1.n202 VDD1.n201 9.3005
R810 VDD1.n178 VDD1.n177 9.3005
R811 VDD1.n176 VDD1.n175 9.3005
R812 VDD1.n119 VDD1.n118 9.3005
R813 VDD1.n170 VDD1.n169 9.3005
R814 VDD1.n168 VDD1.n167 9.3005
R815 VDD1.n123 VDD1.n122 9.3005
R816 VDD1.n162 VDD1.n161 9.3005
R817 VDD1.n135 VDD1.n134 9.3005
R818 VDD1.n142 VDD1.n141 9.3005
R819 VDD1.n144 VDD1.n143 9.3005
R820 VDD1.n131 VDD1.n130 9.3005
R821 VDD1.n150 VDD1.n149 9.3005
R822 VDD1.n152 VDD1.n151 9.3005
R823 VDD1.n153 VDD1.n126 9.3005
R824 VDD1.n160 VDD1.n159 9.3005
R825 VDD1.n115 VDD1.n114 9.3005
R826 VDD1.n88 VDD1.n87 8.92171
R827 VDD1.n72 VDD1.n14 8.92171
R828 VDD1.n43 VDD1.n32 8.92171
R829 VDD1.n144 VDD1.n133 8.92171
R830 VDD1.n175 VDD1.n117 8.92171
R831 VDD1.n191 VDD1.n190 8.92171
R832 VDD1.n84 VDD1.n8 8.14595
R833 VDD1.n76 VDD1.n75 8.14595
R834 VDD1.n40 VDD1.n39 8.14595
R835 VDD1.n141 VDD1.n140 8.14595
R836 VDD1.n179 VDD1.n178 8.14595
R837 VDD1.n187 VDD1.n111 8.14595
R838 VDD1.n83 VDD1.n10 7.3702
R839 VDD1.n79 VDD1.n12 7.3702
R840 VDD1.n36 VDD1.n34 7.3702
R841 VDD1.n137 VDD1.n135 7.3702
R842 VDD1.n182 VDD1.n115 7.3702
R843 VDD1.n186 VDD1.n113 7.3702
R844 VDD1.n80 VDD1.n10 6.59444
R845 VDD1.n80 VDD1.n79 6.59444
R846 VDD1.n183 VDD1.n182 6.59444
R847 VDD1.n183 VDD1.n113 6.59444
R848 VDD1.n84 VDD1.n83 5.81868
R849 VDD1.n76 VDD1.n12 5.81868
R850 VDD1.n39 VDD1.n34 5.81868
R851 VDD1.n140 VDD1.n135 5.81868
R852 VDD1.n179 VDD1.n115 5.81868
R853 VDD1.n187 VDD1.n186 5.81868
R854 VDD1.n87 VDD1.n8 5.04292
R855 VDD1.n75 VDD1.n14 5.04292
R856 VDD1.n40 VDD1.n32 5.04292
R857 VDD1.n141 VDD1.n133 5.04292
R858 VDD1.n178 VDD1.n117 5.04292
R859 VDD1.n190 VDD1.n111 5.04292
R860 VDD1.n88 VDD1.n6 4.26717
R861 VDD1.n72 VDD1.n71 4.26717
R862 VDD1.n44 VDD1.n43 4.26717
R863 VDD1.n145 VDD1.n144 4.26717
R864 VDD1.n175 VDD1.n174 4.26717
R865 VDD1.n191 VDD1.n109 4.26717
R866 VDD1.n92 VDD1.n91 3.49141
R867 VDD1.n68 VDD1.n16 3.49141
R868 VDD1.n47 VDD1.n30 3.49141
R869 VDD1.n148 VDD1.n131 3.49141
R870 VDD1.n171 VDD1.n119 3.49141
R871 VDD1.n195 VDD1.n194 3.49141
R872 VDD1.n136 VDD1.n134 2.84303
R873 VDD1.n35 VDD1.n33 2.84303
R874 VDD1.n95 VDD1.n4 2.71565
R875 VDD1.n67 VDD1.n18 2.71565
R876 VDD1.n48 VDD1.n28 2.71565
R877 VDD1.n149 VDD1.n129 2.71565
R878 VDD1.n170 VDD1.n121 2.71565
R879 VDD1.n198 VDD1.n107 2.71565
R880 VDD1.n96 VDD1.n2 1.93989
R881 VDD1.n64 VDD1.n63 1.93989
R882 VDD1.n52 VDD1.n51 1.93989
R883 VDD1.n154 VDD1.n152 1.93989
R884 VDD1.n167 VDD1.n166 1.93989
R885 VDD1.n199 VDD1.n105 1.93989
R886 VDD1.n100 VDD1.n99 1.16414
R887 VDD1.n60 VDD1.n20 1.16414
R888 VDD1.n55 VDD1.n25 1.16414
R889 VDD1.n153 VDD1.n127 1.16414
R890 VDD1.n163 VDD1.n123 1.16414
R891 VDD1.n203 VDD1.n202 1.16414
R892 VDD1.n102 VDD1.n0 0.388379
R893 VDD1.n59 VDD1.n22 0.388379
R894 VDD1.n56 VDD1.n24 0.388379
R895 VDD1.n159 VDD1.n158 0.388379
R896 VDD1.n162 VDD1.n125 0.388379
R897 VDD1.n205 VDD1.n103 0.388379
R898 VDD1.n98 VDD1.n97 0.155672
R899 VDD1.n97 VDD1.n3 0.155672
R900 VDD1.n90 VDD1.n3 0.155672
R901 VDD1.n90 VDD1.n89 0.155672
R902 VDD1.n89 VDD1.n7 0.155672
R903 VDD1.n82 VDD1.n7 0.155672
R904 VDD1.n82 VDD1.n81 0.155672
R905 VDD1.n81 VDD1.n11 0.155672
R906 VDD1.n74 VDD1.n11 0.155672
R907 VDD1.n74 VDD1.n73 0.155672
R908 VDD1.n73 VDD1.n15 0.155672
R909 VDD1.n66 VDD1.n15 0.155672
R910 VDD1.n66 VDD1.n65 0.155672
R911 VDD1.n65 VDD1.n19 0.155672
R912 VDD1.n58 VDD1.n19 0.155672
R913 VDD1.n58 VDD1.n57 0.155672
R914 VDD1.n57 VDD1.n23 0.155672
R915 VDD1.n50 VDD1.n23 0.155672
R916 VDD1.n50 VDD1.n49 0.155672
R917 VDD1.n49 VDD1.n29 0.155672
R918 VDD1.n42 VDD1.n29 0.155672
R919 VDD1.n42 VDD1.n41 0.155672
R920 VDD1.n41 VDD1.n33 0.155672
R921 VDD1.n142 VDD1.n134 0.155672
R922 VDD1.n143 VDD1.n142 0.155672
R923 VDD1.n143 VDD1.n130 0.155672
R924 VDD1.n150 VDD1.n130 0.155672
R925 VDD1.n151 VDD1.n150 0.155672
R926 VDD1.n151 VDD1.n126 0.155672
R927 VDD1.n160 VDD1.n126 0.155672
R928 VDD1.n161 VDD1.n160 0.155672
R929 VDD1.n161 VDD1.n122 0.155672
R930 VDD1.n168 VDD1.n122 0.155672
R931 VDD1.n169 VDD1.n168 0.155672
R932 VDD1.n169 VDD1.n118 0.155672
R933 VDD1.n176 VDD1.n118 0.155672
R934 VDD1.n177 VDD1.n176 0.155672
R935 VDD1.n177 VDD1.n114 0.155672
R936 VDD1.n184 VDD1.n114 0.155672
R937 VDD1.n185 VDD1.n184 0.155672
R938 VDD1.n185 VDD1.n110 0.155672
R939 VDD1.n192 VDD1.n110 0.155672
R940 VDD1.n193 VDD1.n192 0.155672
R941 VDD1.n193 VDD1.n106 0.155672
R942 VDD1.n200 VDD1.n106 0.155672
R943 VDD1.n201 VDD1.n200 0.155672
R944 B.n863 B.n862 585
R945 B.n864 B.n863 585
R946 B.n379 B.n113 585
R947 B.n378 B.n377 585
R948 B.n376 B.n375 585
R949 B.n374 B.n373 585
R950 B.n372 B.n371 585
R951 B.n370 B.n369 585
R952 B.n368 B.n367 585
R953 B.n366 B.n365 585
R954 B.n364 B.n363 585
R955 B.n362 B.n361 585
R956 B.n360 B.n359 585
R957 B.n358 B.n357 585
R958 B.n356 B.n355 585
R959 B.n354 B.n353 585
R960 B.n352 B.n351 585
R961 B.n350 B.n349 585
R962 B.n348 B.n347 585
R963 B.n346 B.n345 585
R964 B.n344 B.n343 585
R965 B.n342 B.n341 585
R966 B.n340 B.n339 585
R967 B.n338 B.n337 585
R968 B.n336 B.n335 585
R969 B.n334 B.n333 585
R970 B.n332 B.n331 585
R971 B.n330 B.n329 585
R972 B.n328 B.n327 585
R973 B.n326 B.n325 585
R974 B.n324 B.n323 585
R975 B.n322 B.n321 585
R976 B.n320 B.n319 585
R977 B.n318 B.n317 585
R978 B.n316 B.n315 585
R979 B.n314 B.n313 585
R980 B.n312 B.n311 585
R981 B.n310 B.n309 585
R982 B.n308 B.n307 585
R983 B.n306 B.n305 585
R984 B.n304 B.n303 585
R985 B.n302 B.n301 585
R986 B.n300 B.n299 585
R987 B.n298 B.n297 585
R988 B.n296 B.n295 585
R989 B.n294 B.n293 585
R990 B.n292 B.n291 585
R991 B.n290 B.n289 585
R992 B.n288 B.n287 585
R993 B.n286 B.n285 585
R994 B.n284 B.n283 585
R995 B.n282 B.n281 585
R996 B.n280 B.n279 585
R997 B.n278 B.n277 585
R998 B.n276 B.n275 585
R999 B.n274 B.n273 585
R1000 B.n272 B.n271 585
R1001 B.n270 B.n269 585
R1002 B.n268 B.n267 585
R1003 B.n266 B.n265 585
R1004 B.n264 B.n263 585
R1005 B.n262 B.n261 585
R1006 B.n260 B.n259 585
R1007 B.n257 B.n256 585
R1008 B.n255 B.n254 585
R1009 B.n253 B.n252 585
R1010 B.n251 B.n250 585
R1011 B.n249 B.n248 585
R1012 B.n247 B.n246 585
R1013 B.n245 B.n244 585
R1014 B.n243 B.n242 585
R1015 B.n241 B.n240 585
R1016 B.n239 B.n238 585
R1017 B.n237 B.n236 585
R1018 B.n235 B.n234 585
R1019 B.n233 B.n232 585
R1020 B.n231 B.n230 585
R1021 B.n229 B.n228 585
R1022 B.n227 B.n226 585
R1023 B.n225 B.n224 585
R1024 B.n223 B.n222 585
R1025 B.n221 B.n220 585
R1026 B.n219 B.n218 585
R1027 B.n217 B.n216 585
R1028 B.n215 B.n214 585
R1029 B.n213 B.n212 585
R1030 B.n211 B.n210 585
R1031 B.n209 B.n208 585
R1032 B.n207 B.n206 585
R1033 B.n205 B.n204 585
R1034 B.n203 B.n202 585
R1035 B.n201 B.n200 585
R1036 B.n199 B.n198 585
R1037 B.n197 B.n196 585
R1038 B.n195 B.n194 585
R1039 B.n193 B.n192 585
R1040 B.n191 B.n190 585
R1041 B.n189 B.n188 585
R1042 B.n187 B.n186 585
R1043 B.n185 B.n184 585
R1044 B.n183 B.n182 585
R1045 B.n181 B.n180 585
R1046 B.n179 B.n178 585
R1047 B.n177 B.n176 585
R1048 B.n175 B.n174 585
R1049 B.n173 B.n172 585
R1050 B.n171 B.n170 585
R1051 B.n169 B.n168 585
R1052 B.n167 B.n166 585
R1053 B.n165 B.n164 585
R1054 B.n163 B.n162 585
R1055 B.n161 B.n160 585
R1056 B.n159 B.n158 585
R1057 B.n157 B.n156 585
R1058 B.n155 B.n154 585
R1059 B.n153 B.n152 585
R1060 B.n151 B.n150 585
R1061 B.n149 B.n148 585
R1062 B.n147 B.n146 585
R1063 B.n145 B.n144 585
R1064 B.n143 B.n142 585
R1065 B.n141 B.n140 585
R1066 B.n139 B.n138 585
R1067 B.n137 B.n136 585
R1068 B.n135 B.n134 585
R1069 B.n133 B.n132 585
R1070 B.n131 B.n130 585
R1071 B.n129 B.n128 585
R1072 B.n127 B.n126 585
R1073 B.n125 B.n124 585
R1074 B.n123 B.n122 585
R1075 B.n121 B.n120 585
R1076 B.n47 B.n46 585
R1077 B.n867 B.n866 585
R1078 B.n861 B.n114 585
R1079 B.n114 B.n44 585
R1080 B.n860 B.n43 585
R1081 B.n871 B.n43 585
R1082 B.n859 B.n42 585
R1083 B.n872 B.n42 585
R1084 B.n858 B.n41 585
R1085 B.n873 B.n41 585
R1086 B.n857 B.n856 585
R1087 B.n856 B.n37 585
R1088 B.n855 B.n36 585
R1089 B.n879 B.n36 585
R1090 B.n854 B.n35 585
R1091 B.n880 B.n35 585
R1092 B.n853 B.n34 585
R1093 B.n881 B.n34 585
R1094 B.n852 B.n851 585
R1095 B.n851 B.n30 585
R1096 B.n850 B.n29 585
R1097 B.n887 B.n29 585
R1098 B.n849 B.n28 585
R1099 B.n888 B.n28 585
R1100 B.n848 B.n27 585
R1101 B.n889 B.n27 585
R1102 B.n847 B.n846 585
R1103 B.n846 B.n23 585
R1104 B.n845 B.n22 585
R1105 B.n895 B.n22 585
R1106 B.n844 B.n21 585
R1107 B.n896 B.n21 585
R1108 B.n843 B.n20 585
R1109 B.n897 B.n20 585
R1110 B.n842 B.n841 585
R1111 B.n841 B.n16 585
R1112 B.n840 B.n15 585
R1113 B.n903 B.n15 585
R1114 B.n839 B.n14 585
R1115 B.n904 B.n14 585
R1116 B.n838 B.n13 585
R1117 B.n905 B.n13 585
R1118 B.n837 B.n836 585
R1119 B.n836 B.n12 585
R1120 B.n835 B.n834 585
R1121 B.n835 B.n8 585
R1122 B.n833 B.n7 585
R1123 B.n912 B.n7 585
R1124 B.n832 B.n6 585
R1125 B.n913 B.n6 585
R1126 B.n831 B.n5 585
R1127 B.n914 B.n5 585
R1128 B.n830 B.n829 585
R1129 B.n829 B.n4 585
R1130 B.n828 B.n380 585
R1131 B.n828 B.n827 585
R1132 B.n818 B.n381 585
R1133 B.n382 B.n381 585
R1134 B.n820 B.n819 585
R1135 B.n821 B.n820 585
R1136 B.n817 B.n386 585
R1137 B.n390 B.n386 585
R1138 B.n816 B.n815 585
R1139 B.n815 B.n814 585
R1140 B.n388 B.n387 585
R1141 B.n389 B.n388 585
R1142 B.n807 B.n806 585
R1143 B.n808 B.n807 585
R1144 B.n805 B.n395 585
R1145 B.n395 B.n394 585
R1146 B.n804 B.n803 585
R1147 B.n803 B.n802 585
R1148 B.n397 B.n396 585
R1149 B.n398 B.n397 585
R1150 B.n795 B.n794 585
R1151 B.n796 B.n795 585
R1152 B.n793 B.n403 585
R1153 B.n403 B.n402 585
R1154 B.n792 B.n791 585
R1155 B.n791 B.n790 585
R1156 B.n405 B.n404 585
R1157 B.n406 B.n405 585
R1158 B.n783 B.n782 585
R1159 B.n784 B.n783 585
R1160 B.n781 B.n411 585
R1161 B.n411 B.n410 585
R1162 B.n780 B.n779 585
R1163 B.n779 B.n778 585
R1164 B.n413 B.n412 585
R1165 B.n414 B.n413 585
R1166 B.n771 B.n770 585
R1167 B.n772 B.n771 585
R1168 B.n769 B.n419 585
R1169 B.n419 B.n418 585
R1170 B.n768 B.n767 585
R1171 B.n767 B.n766 585
R1172 B.n421 B.n420 585
R1173 B.n422 B.n421 585
R1174 B.n762 B.n761 585
R1175 B.n425 B.n424 585
R1176 B.n758 B.n757 585
R1177 B.n759 B.n758 585
R1178 B.n756 B.n491 585
R1179 B.n755 B.n754 585
R1180 B.n753 B.n752 585
R1181 B.n751 B.n750 585
R1182 B.n749 B.n748 585
R1183 B.n747 B.n746 585
R1184 B.n745 B.n744 585
R1185 B.n743 B.n742 585
R1186 B.n741 B.n740 585
R1187 B.n739 B.n738 585
R1188 B.n737 B.n736 585
R1189 B.n735 B.n734 585
R1190 B.n733 B.n732 585
R1191 B.n731 B.n730 585
R1192 B.n729 B.n728 585
R1193 B.n727 B.n726 585
R1194 B.n725 B.n724 585
R1195 B.n723 B.n722 585
R1196 B.n721 B.n720 585
R1197 B.n719 B.n718 585
R1198 B.n717 B.n716 585
R1199 B.n715 B.n714 585
R1200 B.n713 B.n712 585
R1201 B.n711 B.n710 585
R1202 B.n709 B.n708 585
R1203 B.n707 B.n706 585
R1204 B.n705 B.n704 585
R1205 B.n703 B.n702 585
R1206 B.n701 B.n700 585
R1207 B.n699 B.n698 585
R1208 B.n697 B.n696 585
R1209 B.n695 B.n694 585
R1210 B.n693 B.n692 585
R1211 B.n691 B.n690 585
R1212 B.n689 B.n688 585
R1213 B.n687 B.n686 585
R1214 B.n685 B.n684 585
R1215 B.n683 B.n682 585
R1216 B.n681 B.n680 585
R1217 B.n679 B.n678 585
R1218 B.n677 B.n676 585
R1219 B.n675 B.n674 585
R1220 B.n673 B.n672 585
R1221 B.n671 B.n670 585
R1222 B.n669 B.n668 585
R1223 B.n667 B.n666 585
R1224 B.n665 B.n664 585
R1225 B.n663 B.n662 585
R1226 B.n661 B.n660 585
R1227 B.n659 B.n658 585
R1228 B.n657 B.n656 585
R1229 B.n655 B.n654 585
R1230 B.n653 B.n652 585
R1231 B.n651 B.n650 585
R1232 B.n649 B.n648 585
R1233 B.n647 B.n646 585
R1234 B.n645 B.n644 585
R1235 B.n643 B.n642 585
R1236 B.n641 B.n640 585
R1237 B.n638 B.n637 585
R1238 B.n636 B.n635 585
R1239 B.n634 B.n633 585
R1240 B.n632 B.n631 585
R1241 B.n630 B.n629 585
R1242 B.n628 B.n627 585
R1243 B.n626 B.n625 585
R1244 B.n624 B.n623 585
R1245 B.n622 B.n621 585
R1246 B.n620 B.n619 585
R1247 B.n618 B.n617 585
R1248 B.n616 B.n615 585
R1249 B.n614 B.n613 585
R1250 B.n612 B.n611 585
R1251 B.n610 B.n609 585
R1252 B.n608 B.n607 585
R1253 B.n606 B.n605 585
R1254 B.n604 B.n603 585
R1255 B.n602 B.n601 585
R1256 B.n600 B.n599 585
R1257 B.n598 B.n597 585
R1258 B.n596 B.n595 585
R1259 B.n594 B.n593 585
R1260 B.n592 B.n591 585
R1261 B.n590 B.n589 585
R1262 B.n588 B.n587 585
R1263 B.n586 B.n585 585
R1264 B.n584 B.n583 585
R1265 B.n582 B.n581 585
R1266 B.n580 B.n579 585
R1267 B.n578 B.n577 585
R1268 B.n576 B.n575 585
R1269 B.n574 B.n573 585
R1270 B.n572 B.n571 585
R1271 B.n570 B.n569 585
R1272 B.n568 B.n567 585
R1273 B.n566 B.n565 585
R1274 B.n564 B.n563 585
R1275 B.n562 B.n561 585
R1276 B.n560 B.n559 585
R1277 B.n558 B.n557 585
R1278 B.n556 B.n555 585
R1279 B.n554 B.n553 585
R1280 B.n552 B.n551 585
R1281 B.n550 B.n549 585
R1282 B.n548 B.n547 585
R1283 B.n546 B.n545 585
R1284 B.n544 B.n543 585
R1285 B.n542 B.n541 585
R1286 B.n540 B.n539 585
R1287 B.n538 B.n537 585
R1288 B.n536 B.n535 585
R1289 B.n534 B.n533 585
R1290 B.n532 B.n531 585
R1291 B.n530 B.n529 585
R1292 B.n528 B.n527 585
R1293 B.n526 B.n525 585
R1294 B.n524 B.n523 585
R1295 B.n522 B.n521 585
R1296 B.n520 B.n519 585
R1297 B.n518 B.n517 585
R1298 B.n516 B.n515 585
R1299 B.n514 B.n513 585
R1300 B.n512 B.n511 585
R1301 B.n510 B.n509 585
R1302 B.n508 B.n507 585
R1303 B.n506 B.n505 585
R1304 B.n504 B.n503 585
R1305 B.n502 B.n501 585
R1306 B.n500 B.n499 585
R1307 B.n498 B.n497 585
R1308 B.n763 B.n423 585
R1309 B.n423 B.n422 585
R1310 B.n765 B.n764 585
R1311 B.n766 B.n765 585
R1312 B.n417 B.n416 585
R1313 B.n418 B.n417 585
R1314 B.n774 B.n773 585
R1315 B.n773 B.n772 585
R1316 B.n775 B.n415 585
R1317 B.n415 B.n414 585
R1318 B.n777 B.n776 585
R1319 B.n778 B.n777 585
R1320 B.n409 B.n408 585
R1321 B.n410 B.n409 585
R1322 B.n786 B.n785 585
R1323 B.n785 B.n784 585
R1324 B.n787 B.n407 585
R1325 B.n407 B.n406 585
R1326 B.n789 B.n788 585
R1327 B.n790 B.n789 585
R1328 B.n401 B.n400 585
R1329 B.n402 B.n401 585
R1330 B.n798 B.n797 585
R1331 B.n797 B.n796 585
R1332 B.n799 B.n399 585
R1333 B.n399 B.n398 585
R1334 B.n801 B.n800 585
R1335 B.n802 B.n801 585
R1336 B.n393 B.n392 585
R1337 B.n394 B.n393 585
R1338 B.n810 B.n809 585
R1339 B.n809 B.n808 585
R1340 B.n811 B.n391 585
R1341 B.n391 B.n389 585
R1342 B.n813 B.n812 585
R1343 B.n814 B.n813 585
R1344 B.n385 B.n384 585
R1345 B.n390 B.n385 585
R1346 B.n823 B.n822 585
R1347 B.n822 B.n821 585
R1348 B.n824 B.n383 585
R1349 B.n383 B.n382 585
R1350 B.n826 B.n825 585
R1351 B.n827 B.n826 585
R1352 B.n3 B.n0 585
R1353 B.n4 B.n3 585
R1354 B.n911 B.n1 585
R1355 B.n912 B.n911 585
R1356 B.n910 B.n909 585
R1357 B.n910 B.n8 585
R1358 B.n908 B.n9 585
R1359 B.n12 B.n9 585
R1360 B.n907 B.n906 585
R1361 B.n906 B.n905 585
R1362 B.n11 B.n10 585
R1363 B.n904 B.n11 585
R1364 B.n902 B.n901 585
R1365 B.n903 B.n902 585
R1366 B.n900 B.n17 585
R1367 B.n17 B.n16 585
R1368 B.n899 B.n898 585
R1369 B.n898 B.n897 585
R1370 B.n19 B.n18 585
R1371 B.n896 B.n19 585
R1372 B.n894 B.n893 585
R1373 B.n895 B.n894 585
R1374 B.n892 B.n24 585
R1375 B.n24 B.n23 585
R1376 B.n891 B.n890 585
R1377 B.n890 B.n889 585
R1378 B.n26 B.n25 585
R1379 B.n888 B.n26 585
R1380 B.n886 B.n885 585
R1381 B.n887 B.n886 585
R1382 B.n884 B.n31 585
R1383 B.n31 B.n30 585
R1384 B.n883 B.n882 585
R1385 B.n882 B.n881 585
R1386 B.n33 B.n32 585
R1387 B.n880 B.n33 585
R1388 B.n878 B.n877 585
R1389 B.n879 B.n878 585
R1390 B.n876 B.n38 585
R1391 B.n38 B.n37 585
R1392 B.n875 B.n874 585
R1393 B.n874 B.n873 585
R1394 B.n40 B.n39 585
R1395 B.n872 B.n40 585
R1396 B.n870 B.n869 585
R1397 B.n871 B.n870 585
R1398 B.n868 B.n45 585
R1399 B.n45 B.n44 585
R1400 B.n915 B.n914 585
R1401 B.n913 B.n2 585
R1402 B.n866 B.n45 487.695
R1403 B.n863 B.n114 487.695
R1404 B.n497 B.n421 487.695
R1405 B.n761 B.n423 487.695
R1406 B.n117 B.t8 449.75
R1407 B.n115 B.t11 449.75
R1408 B.n494 B.t5 449.75
R1409 B.n492 B.t15 449.75
R1410 B.n117 B.t6 404.327
R1411 B.n115 B.t10 404.327
R1412 B.n494 B.t2 404.327
R1413 B.n492 B.t13 404.327
R1414 B.n116 B.t12 398.745
R1415 B.n495 B.t4 398.745
R1416 B.n118 B.t9 398.745
R1417 B.n493 B.t14 398.745
R1418 B.n864 B.n112 256.663
R1419 B.n864 B.n111 256.663
R1420 B.n864 B.n110 256.663
R1421 B.n864 B.n109 256.663
R1422 B.n864 B.n108 256.663
R1423 B.n864 B.n107 256.663
R1424 B.n864 B.n106 256.663
R1425 B.n864 B.n105 256.663
R1426 B.n864 B.n104 256.663
R1427 B.n864 B.n103 256.663
R1428 B.n864 B.n102 256.663
R1429 B.n864 B.n101 256.663
R1430 B.n864 B.n100 256.663
R1431 B.n864 B.n99 256.663
R1432 B.n864 B.n98 256.663
R1433 B.n864 B.n97 256.663
R1434 B.n864 B.n96 256.663
R1435 B.n864 B.n95 256.663
R1436 B.n864 B.n94 256.663
R1437 B.n864 B.n93 256.663
R1438 B.n864 B.n92 256.663
R1439 B.n864 B.n91 256.663
R1440 B.n864 B.n90 256.663
R1441 B.n864 B.n89 256.663
R1442 B.n864 B.n88 256.663
R1443 B.n864 B.n87 256.663
R1444 B.n864 B.n86 256.663
R1445 B.n864 B.n85 256.663
R1446 B.n864 B.n84 256.663
R1447 B.n864 B.n83 256.663
R1448 B.n864 B.n82 256.663
R1449 B.n864 B.n81 256.663
R1450 B.n864 B.n80 256.663
R1451 B.n864 B.n79 256.663
R1452 B.n864 B.n78 256.663
R1453 B.n864 B.n77 256.663
R1454 B.n864 B.n76 256.663
R1455 B.n864 B.n75 256.663
R1456 B.n864 B.n74 256.663
R1457 B.n864 B.n73 256.663
R1458 B.n864 B.n72 256.663
R1459 B.n864 B.n71 256.663
R1460 B.n864 B.n70 256.663
R1461 B.n864 B.n69 256.663
R1462 B.n864 B.n68 256.663
R1463 B.n864 B.n67 256.663
R1464 B.n864 B.n66 256.663
R1465 B.n864 B.n65 256.663
R1466 B.n864 B.n64 256.663
R1467 B.n864 B.n63 256.663
R1468 B.n864 B.n62 256.663
R1469 B.n864 B.n61 256.663
R1470 B.n864 B.n60 256.663
R1471 B.n864 B.n59 256.663
R1472 B.n864 B.n58 256.663
R1473 B.n864 B.n57 256.663
R1474 B.n864 B.n56 256.663
R1475 B.n864 B.n55 256.663
R1476 B.n864 B.n54 256.663
R1477 B.n864 B.n53 256.663
R1478 B.n864 B.n52 256.663
R1479 B.n864 B.n51 256.663
R1480 B.n864 B.n50 256.663
R1481 B.n864 B.n49 256.663
R1482 B.n864 B.n48 256.663
R1483 B.n865 B.n864 256.663
R1484 B.n760 B.n759 256.663
R1485 B.n759 B.n426 256.663
R1486 B.n759 B.n427 256.663
R1487 B.n759 B.n428 256.663
R1488 B.n759 B.n429 256.663
R1489 B.n759 B.n430 256.663
R1490 B.n759 B.n431 256.663
R1491 B.n759 B.n432 256.663
R1492 B.n759 B.n433 256.663
R1493 B.n759 B.n434 256.663
R1494 B.n759 B.n435 256.663
R1495 B.n759 B.n436 256.663
R1496 B.n759 B.n437 256.663
R1497 B.n759 B.n438 256.663
R1498 B.n759 B.n439 256.663
R1499 B.n759 B.n440 256.663
R1500 B.n759 B.n441 256.663
R1501 B.n759 B.n442 256.663
R1502 B.n759 B.n443 256.663
R1503 B.n759 B.n444 256.663
R1504 B.n759 B.n445 256.663
R1505 B.n759 B.n446 256.663
R1506 B.n759 B.n447 256.663
R1507 B.n759 B.n448 256.663
R1508 B.n759 B.n449 256.663
R1509 B.n759 B.n450 256.663
R1510 B.n759 B.n451 256.663
R1511 B.n759 B.n452 256.663
R1512 B.n759 B.n453 256.663
R1513 B.n759 B.n454 256.663
R1514 B.n759 B.n455 256.663
R1515 B.n759 B.n456 256.663
R1516 B.n759 B.n457 256.663
R1517 B.n759 B.n458 256.663
R1518 B.n759 B.n459 256.663
R1519 B.n759 B.n460 256.663
R1520 B.n759 B.n461 256.663
R1521 B.n759 B.n462 256.663
R1522 B.n759 B.n463 256.663
R1523 B.n759 B.n464 256.663
R1524 B.n759 B.n465 256.663
R1525 B.n759 B.n466 256.663
R1526 B.n759 B.n467 256.663
R1527 B.n759 B.n468 256.663
R1528 B.n759 B.n469 256.663
R1529 B.n759 B.n470 256.663
R1530 B.n759 B.n471 256.663
R1531 B.n759 B.n472 256.663
R1532 B.n759 B.n473 256.663
R1533 B.n759 B.n474 256.663
R1534 B.n759 B.n475 256.663
R1535 B.n759 B.n476 256.663
R1536 B.n759 B.n477 256.663
R1537 B.n759 B.n478 256.663
R1538 B.n759 B.n479 256.663
R1539 B.n759 B.n480 256.663
R1540 B.n759 B.n481 256.663
R1541 B.n759 B.n482 256.663
R1542 B.n759 B.n483 256.663
R1543 B.n759 B.n484 256.663
R1544 B.n759 B.n485 256.663
R1545 B.n759 B.n486 256.663
R1546 B.n759 B.n487 256.663
R1547 B.n759 B.n488 256.663
R1548 B.n759 B.n489 256.663
R1549 B.n759 B.n490 256.663
R1550 B.n917 B.n916 256.663
R1551 B.n120 B.n47 163.367
R1552 B.n124 B.n123 163.367
R1553 B.n128 B.n127 163.367
R1554 B.n132 B.n131 163.367
R1555 B.n136 B.n135 163.367
R1556 B.n140 B.n139 163.367
R1557 B.n144 B.n143 163.367
R1558 B.n148 B.n147 163.367
R1559 B.n152 B.n151 163.367
R1560 B.n156 B.n155 163.367
R1561 B.n160 B.n159 163.367
R1562 B.n164 B.n163 163.367
R1563 B.n168 B.n167 163.367
R1564 B.n172 B.n171 163.367
R1565 B.n176 B.n175 163.367
R1566 B.n180 B.n179 163.367
R1567 B.n184 B.n183 163.367
R1568 B.n188 B.n187 163.367
R1569 B.n192 B.n191 163.367
R1570 B.n196 B.n195 163.367
R1571 B.n200 B.n199 163.367
R1572 B.n204 B.n203 163.367
R1573 B.n208 B.n207 163.367
R1574 B.n212 B.n211 163.367
R1575 B.n216 B.n215 163.367
R1576 B.n220 B.n219 163.367
R1577 B.n224 B.n223 163.367
R1578 B.n228 B.n227 163.367
R1579 B.n232 B.n231 163.367
R1580 B.n236 B.n235 163.367
R1581 B.n240 B.n239 163.367
R1582 B.n244 B.n243 163.367
R1583 B.n248 B.n247 163.367
R1584 B.n252 B.n251 163.367
R1585 B.n256 B.n255 163.367
R1586 B.n261 B.n260 163.367
R1587 B.n265 B.n264 163.367
R1588 B.n269 B.n268 163.367
R1589 B.n273 B.n272 163.367
R1590 B.n277 B.n276 163.367
R1591 B.n281 B.n280 163.367
R1592 B.n285 B.n284 163.367
R1593 B.n289 B.n288 163.367
R1594 B.n293 B.n292 163.367
R1595 B.n297 B.n296 163.367
R1596 B.n301 B.n300 163.367
R1597 B.n305 B.n304 163.367
R1598 B.n309 B.n308 163.367
R1599 B.n313 B.n312 163.367
R1600 B.n317 B.n316 163.367
R1601 B.n321 B.n320 163.367
R1602 B.n325 B.n324 163.367
R1603 B.n329 B.n328 163.367
R1604 B.n333 B.n332 163.367
R1605 B.n337 B.n336 163.367
R1606 B.n341 B.n340 163.367
R1607 B.n345 B.n344 163.367
R1608 B.n349 B.n348 163.367
R1609 B.n353 B.n352 163.367
R1610 B.n357 B.n356 163.367
R1611 B.n361 B.n360 163.367
R1612 B.n365 B.n364 163.367
R1613 B.n369 B.n368 163.367
R1614 B.n373 B.n372 163.367
R1615 B.n377 B.n376 163.367
R1616 B.n863 B.n113 163.367
R1617 B.n767 B.n421 163.367
R1618 B.n767 B.n419 163.367
R1619 B.n771 B.n419 163.367
R1620 B.n771 B.n413 163.367
R1621 B.n779 B.n413 163.367
R1622 B.n779 B.n411 163.367
R1623 B.n783 B.n411 163.367
R1624 B.n783 B.n405 163.367
R1625 B.n791 B.n405 163.367
R1626 B.n791 B.n403 163.367
R1627 B.n795 B.n403 163.367
R1628 B.n795 B.n397 163.367
R1629 B.n803 B.n397 163.367
R1630 B.n803 B.n395 163.367
R1631 B.n807 B.n395 163.367
R1632 B.n807 B.n388 163.367
R1633 B.n815 B.n388 163.367
R1634 B.n815 B.n386 163.367
R1635 B.n820 B.n386 163.367
R1636 B.n820 B.n381 163.367
R1637 B.n828 B.n381 163.367
R1638 B.n829 B.n828 163.367
R1639 B.n829 B.n5 163.367
R1640 B.n6 B.n5 163.367
R1641 B.n7 B.n6 163.367
R1642 B.n835 B.n7 163.367
R1643 B.n836 B.n835 163.367
R1644 B.n836 B.n13 163.367
R1645 B.n14 B.n13 163.367
R1646 B.n15 B.n14 163.367
R1647 B.n841 B.n15 163.367
R1648 B.n841 B.n20 163.367
R1649 B.n21 B.n20 163.367
R1650 B.n22 B.n21 163.367
R1651 B.n846 B.n22 163.367
R1652 B.n846 B.n27 163.367
R1653 B.n28 B.n27 163.367
R1654 B.n29 B.n28 163.367
R1655 B.n851 B.n29 163.367
R1656 B.n851 B.n34 163.367
R1657 B.n35 B.n34 163.367
R1658 B.n36 B.n35 163.367
R1659 B.n856 B.n36 163.367
R1660 B.n856 B.n41 163.367
R1661 B.n42 B.n41 163.367
R1662 B.n43 B.n42 163.367
R1663 B.n114 B.n43 163.367
R1664 B.n758 B.n425 163.367
R1665 B.n758 B.n491 163.367
R1666 B.n754 B.n753 163.367
R1667 B.n750 B.n749 163.367
R1668 B.n746 B.n745 163.367
R1669 B.n742 B.n741 163.367
R1670 B.n738 B.n737 163.367
R1671 B.n734 B.n733 163.367
R1672 B.n730 B.n729 163.367
R1673 B.n726 B.n725 163.367
R1674 B.n722 B.n721 163.367
R1675 B.n718 B.n717 163.367
R1676 B.n714 B.n713 163.367
R1677 B.n710 B.n709 163.367
R1678 B.n706 B.n705 163.367
R1679 B.n702 B.n701 163.367
R1680 B.n698 B.n697 163.367
R1681 B.n694 B.n693 163.367
R1682 B.n690 B.n689 163.367
R1683 B.n686 B.n685 163.367
R1684 B.n682 B.n681 163.367
R1685 B.n678 B.n677 163.367
R1686 B.n674 B.n673 163.367
R1687 B.n670 B.n669 163.367
R1688 B.n666 B.n665 163.367
R1689 B.n662 B.n661 163.367
R1690 B.n658 B.n657 163.367
R1691 B.n654 B.n653 163.367
R1692 B.n650 B.n649 163.367
R1693 B.n646 B.n645 163.367
R1694 B.n642 B.n641 163.367
R1695 B.n637 B.n636 163.367
R1696 B.n633 B.n632 163.367
R1697 B.n629 B.n628 163.367
R1698 B.n625 B.n624 163.367
R1699 B.n621 B.n620 163.367
R1700 B.n617 B.n616 163.367
R1701 B.n613 B.n612 163.367
R1702 B.n609 B.n608 163.367
R1703 B.n605 B.n604 163.367
R1704 B.n601 B.n600 163.367
R1705 B.n597 B.n596 163.367
R1706 B.n593 B.n592 163.367
R1707 B.n589 B.n588 163.367
R1708 B.n585 B.n584 163.367
R1709 B.n581 B.n580 163.367
R1710 B.n577 B.n576 163.367
R1711 B.n573 B.n572 163.367
R1712 B.n569 B.n568 163.367
R1713 B.n565 B.n564 163.367
R1714 B.n561 B.n560 163.367
R1715 B.n557 B.n556 163.367
R1716 B.n553 B.n552 163.367
R1717 B.n549 B.n548 163.367
R1718 B.n545 B.n544 163.367
R1719 B.n541 B.n540 163.367
R1720 B.n537 B.n536 163.367
R1721 B.n533 B.n532 163.367
R1722 B.n529 B.n528 163.367
R1723 B.n525 B.n524 163.367
R1724 B.n521 B.n520 163.367
R1725 B.n517 B.n516 163.367
R1726 B.n513 B.n512 163.367
R1727 B.n509 B.n508 163.367
R1728 B.n505 B.n504 163.367
R1729 B.n501 B.n500 163.367
R1730 B.n765 B.n423 163.367
R1731 B.n765 B.n417 163.367
R1732 B.n773 B.n417 163.367
R1733 B.n773 B.n415 163.367
R1734 B.n777 B.n415 163.367
R1735 B.n777 B.n409 163.367
R1736 B.n785 B.n409 163.367
R1737 B.n785 B.n407 163.367
R1738 B.n789 B.n407 163.367
R1739 B.n789 B.n401 163.367
R1740 B.n797 B.n401 163.367
R1741 B.n797 B.n399 163.367
R1742 B.n801 B.n399 163.367
R1743 B.n801 B.n393 163.367
R1744 B.n809 B.n393 163.367
R1745 B.n809 B.n391 163.367
R1746 B.n813 B.n391 163.367
R1747 B.n813 B.n385 163.367
R1748 B.n822 B.n385 163.367
R1749 B.n822 B.n383 163.367
R1750 B.n826 B.n383 163.367
R1751 B.n826 B.n3 163.367
R1752 B.n915 B.n3 163.367
R1753 B.n911 B.n2 163.367
R1754 B.n911 B.n910 163.367
R1755 B.n910 B.n9 163.367
R1756 B.n906 B.n9 163.367
R1757 B.n906 B.n11 163.367
R1758 B.n902 B.n11 163.367
R1759 B.n902 B.n17 163.367
R1760 B.n898 B.n17 163.367
R1761 B.n898 B.n19 163.367
R1762 B.n894 B.n19 163.367
R1763 B.n894 B.n24 163.367
R1764 B.n890 B.n24 163.367
R1765 B.n890 B.n26 163.367
R1766 B.n886 B.n26 163.367
R1767 B.n886 B.n31 163.367
R1768 B.n882 B.n31 163.367
R1769 B.n882 B.n33 163.367
R1770 B.n878 B.n33 163.367
R1771 B.n878 B.n38 163.367
R1772 B.n874 B.n38 163.367
R1773 B.n874 B.n40 163.367
R1774 B.n870 B.n40 163.367
R1775 B.n870 B.n45 163.367
R1776 B.n866 B.n865 71.676
R1777 B.n120 B.n48 71.676
R1778 B.n124 B.n49 71.676
R1779 B.n128 B.n50 71.676
R1780 B.n132 B.n51 71.676
R1781 B.n136 B.n52 71.676
R1782 B.n140 B.n53 71.676
R1783 B.n144 B.n54 71.676
R1784 B.n148 B.n55 71.676
R1785 B.n152 B.n56 71.676
R1786 B.n156 B.n57 71.676
R1787 B.n160 B.n58 71.676
R1788 B.n164 B.n59 71.676
R1789 B.n168 B.n60 71.676
R1790 B.n172 B.n61 71.676
R1791 B.n176 B.n62 71.676
R1792 B.n180 B.n63 71.676
R1793 B.n184 B.n64 71.676
R1794 B.n188 B.n65 71.676
R1795 B.n192 B.n66 71.676
R1796 B.n196 B.n67 71.676
R1797 B.n200 B.n68 71.676
R1798 B.n204 B.n69 71.676
R1799 B.n208 B.n70 71.676
R1800 B.n212 B.n71 71.676
R1801 B.n216 B.n72 71.676
R1802 B.n220 B.n73 71.676
R1803 B.n224 B.n74 71.676
R1804 B.n228 B.n75 71.676
R1805 B.n232 B.n76 71.676
R1806 B.n236 B.n77 71.676
R1807 B.n240 B.n78 71.676
R1808 B.n244 B.n79 71.676
R1809 B.n248 B.n80 71.676
R1810 B.n252 B.n81 71.676
R1811 B.n256 B.n82 71.676
R1812 B.n261 B.n83 71.676
R1813 B.n265 B.n84 71.676
R1814 B.n269 B.n85 71.676
R1815 B.n273 B.n86 71.676
R1816 B.n277 B.n87 71.676
R1817 B.n281 B.n88 71.676
R1818 B.n285 B.n89 71.676
R1819 B.n289 B.n90 71.676
R1820 B.n293 B.n91 71.676
R1821 B.n297 B.n92 71.676
R1822 B.n301 B.n93 71.676
R1823 B.n305 B.n94 71.676
R1824 B.n309 B.n95 71.676
R1825 B.n313 B.n96 71.676
R1826 B.n317 B.n97 71.676
R1827 B.n321 B.n98 71.676
R1828 B.n325 B.n99 71.676
R1829 B.n329 B.n100 71.676
R1830 B.n333 B.n101 71.676
R1831 B.n337 B.n102 71.676
R1832 B.n341 B.n103 71.676
R1833 B.n345 B.n104 71.676
R1834 B.n349 B.n105 71.676
R1835 B.n353 B.n106 71.676
R1836 B.n357 B.n107 71.676
R1837 B.n361 B.n108 71.676
R1838 B.n365 B.n109 71.676
R1839 B.n369 B.n110 71.676
R1840 B.n373 B.n111 71.676
R1841 B.n377 B.n112 71.676
R1842 B.n113 B.n112 71.676
R1843 B.n376 B.n111 71.676
R1844 B.n372 B.n110 71.676
R1845 B.n368 B.n109 71.676
R1846 B.n364 B.n108 71.676
R1847 B.n360 B.n107 71.676
R1848 B.n356 B.n106 71.676
R1849 B.n352 B.n105 71.676
R1850 B.n348 B.n104 71.676
R1851 B.n344 B.n103 71.676
R1852 B.n340 B.n102 71.676
R1853 B.n336 B.n101 71.676
R1854 B.n332 B.n100 71.676
R1855 B.n328 B.n99 71.676
R1856 B.n324 B.n98 71.676
R1857 B.n320 B.n97 71.676
R1858 B.n316 B.n96 71.676
R1859 B.n312 B.n95 71.676
R1860 B.n308 B.n94 71.676
R1861 B.n304 B.n93 71.676
R1862 B.n300 B.n92 71.676
R1863 B.n296 B.n91 71.676
R1864 B.n292 B.n90 71.676
R1865 B.n288 B.n89 71.676
R1866 B.n284 B.n88 71.676
R1867 B.n280 B.n87 71.676
R1868 B.n276 B.n86 71.676
R1869 B.n272 B.n85 71.676
R1870 B.n268 B.n84 71.676
R1871 B.n264 B.n83 71.676
R1872 B.n260 B.n82 71.676
R1873 B.n255 B.n81 71.676
R1874 B.n251 B.n80 71.676
R1875 B.n247 B.n79 71.676
R1876 B.n243 B.n78 71.676
R1877 B.n239 B.n77 71.676
R1878 B.n235 B.n76 71.676
R1879 B.n231 B.n75 71.676
R1880 B.n227 B.n74 71.676
R1881 B.n223 B.n73 71.676
R1882 B.n219 B.n72 71.676
R1883 B.n215 B.n71 71.676
R1884 B.n211 B.n70 71.676
R1885 B.n207 B.n69 71.676
R1886 B.n203 B.n68 71.676
R1887 B.n199 B.n67 71.676
R1888 B.n195 B.n66 71.676
R1889 B.n191 B.n65 71.676
R1890 B.n187 B.n64 71.676
R1891 B.n183 B.n63 71.676
R1892 B.n179 B.n62 71.676
R1893 B.n175 B.n61 71.676
R1894 B.n171 B.n60 71.676
R1895 B.n167 B.n59 71.676
R1896 B.n163 B.n58 71.676
R1897 B.n159 B.n57 71.676
R1898 B.n155 B.n56 71.676
R1899 B.n151 B.n55 71.676
R1900 B.n147 B.n54 71.676
R1901 B.n143 B.n53 71.676
R1902 B.n139 B.n52 71.676
R1903 B.n135 B.n51 71.676
R1904 B.n131 B.n50 71.676
R1905 B.n127 B.n49 71.676
R1906 B.n123 B.n48 71.676
R1907 B.n865 B.n47 71.676
R1908 B.n761 B.n760 71.676
R1909 B.n491 B.n426 71.676
R1910 B.n753 B.n427 71.676
R1911 B.n749 B.n428 71.676
R1912 B.n745 B.n429 71.676
R1913 B.n741 B.n430 71.676
R1914 B.n737 B.n431 71.676
R1915 B.n733 B.n432 71.676
R1916 B.n729 B.n433 71.676
R1917 B.n725 B.n434 71.676
R1918 B.n721 B.n435 71.676
R1919 B.n717 B.n436 71.676
R1920 B.n713 B.n437 71.676
R1921 B.n709 B.n438 71.676
R1922 B.n705 B.n439 71.676
R1923 B.n701 B.n440 71.676
R1924 B.n697 B.n441 71.676
R1925 B.n693 B.n442 71.676
R1926 B.n689 B.n443 71.676
R1927 B.n685 B.n444 71.676
R1928 B.n681 B.n445 71.676
R1929 B.n677 B.n446 71.676
R1930 B.n673 B.n447 71.676
R1931 B.n669 B.n448 71.676
R1932 B.n665 B.n449 71.676
R1933 B.n661 B.n450 71.676
R1934 B.n657 B.n451 71.676
R1935 B.n653 B.n452 71.676
R1936 B.n649 B.n453 71.676
R1937 B.n645 B.n454 71.676
R1938 B.n641 B.n455 71.676
R1939 B.n636 B.n456 71.676
R1940 B.n632 B.n457 71.676
R1941 B.n628 B.n458 71.676
R1942 B.n624 B.n459 71.676
R1943 B.n620 B.n460 71.676
R1944 B.n616 B.n461 71.676
R1945 B.n612 B.n462 71.676
R1946 B.n608 B.n463 71.676
R1947 B.n604 B.n464 71.676
R1948 B.n600 B.n465 71.676
R1949 B.n596 B.n466 71.676
R1950 B.n592 B.n467 71.676
R1951 B.n588 B.n468 71.676
R1952 B.n584 B.n469 71.676
R1953 B.n580 B.n470 71.676
R1954 B.n576 B.n471 71.676
R1955 B.n572 B.n472 71.676
R1956 B.n568 B.n473 71.676
R1957 B.n564 B.n474 71.676
R1958 B.n560 B.n475 71.676
R1959 B.n556 B.n476 71.676
R1960 B.n552 B.n477 71.676
R1961 B.n548 B.n478 71.676
R1962 B.n544 B.n479 71.676
R1963 B.n540 B.n480 71.676
R1964 B.n536 B.n481 71.676
R1965 B.n532 B.n482 71.676
R1966 B.n528 B.n483 71.676
R1967 B.n524 B.n484 71.676
R1968 B.n520 B.n485 71.676
R1969 B.n516 B.n486 71.676
R1970 B.n512 B.n487 71.676
R1971 B.n508 B.n488 71.676
R1972 B.n504 B.n489 71.676
R1973 B.n500 B.n490 71.676
R1974 B.n760 B.n425 71.676
R1975 B.n754 B.n426 71.676
R1976 B.n750 B.n427 71.676
R1977 B.n746 B.n428 71.676
R1978 B.n742 B.n429 71.676
R1979 B.n738 B.n430 71.676
R1980 B.n734 B.n431 71.676
R1981 B.n730 B.n432 71.676
R1982 B.n726 B.n433 71.676
R1983 B.n722 B.n434 71.676
R1984 B.n718 B.n435 71.676
R1985 B.n714 B.n436 71.676
R1986 B.n710 B.n437 71.676
R1987 B.n706 B.n438 71.676
R1988 B.n702 B.n439 71.676
R1989 B.n698 B.n440 71.676
R1990 B.n694 B.n441 71.676
R1991 B.n690 B.n442 71.676
R1992 B.n686 B.n443 71.676
R1993 B.n682 B.n444 71.676
R1994 B.n678 B.n445 71.676
R1995 B.n674 B.n446 71.676
R1996 B.n670 B.n447 71.676
R1997 B.n666 B.n448 71.676
R1998 B.n662 B.n449 71.676
R1999 B.n658 B.n450 71.676
R2000 B.n654 B.n451 71.676
R2001 B.n650 B.n452 71.676
R2002 B.n646 B.n453 71.676
R2003 B.n642 B.n454 71.676
R2004 B.n637 B.n455 71.676
R2005 B.n633 B.n456 71.676
R2006 B.n629 B.n457 71.676
R2007 B.n625 B.n458 71.676
R2008 B.n621 B.n459 71.676
R2009 B.n617 B.n460 71.676
R2010 B.n613 B.n461 71.676
R2011 B.n609 B.n462 71.676
R2012 B.n605 B.n463 71.676
R2013 B.n601 B.n464 71.676
R2014 B.n597 B.n465 71.676
R2015 B.n593 B.n466 71.676
R2016 B.n589 B.n467 71.676
R2017 B.n585 B.n468 71.676
R2018 B.n581 B.n469 71.676
R2019 B.n577 B.n470 71.676
R2020 B.n573 B.n471 71.676
R2021 B.n569 B.n472 71.676
R2022 B.n565 B.n473 71.676
R2023 B.n561 B.n474 71.676
R2024 B.n557 B.n475 71.676
R2025 B.n553 B.n476 71.676
R2026 B.n549 B.n477 71.676
R2027 B.n545 B.n478 71.676
R2028 B.n541 B.n479 71.676
R2029 B.n537 B.n480 71.676
R2030 B.n533 B.n481 71.676
R2031 B.n529 B.n482 71.676
R2032 B.n525 B.n483 71.676
R2033 B.n521 B.n484 71.676
R2034 B.n517 B.n485 71.676
R2035 B.n513 B.n486 71.676
R2036 B.n509 B.n487 71.676
R2037 B.n505 B.n488 71.676
R2038 B.n501 B.n489 71.676
R2039 B.n497 B.n490 71.676
R2040 B.n916 B.n915 71.676
R2041 B.n916 B.n2 71.676
R2042 B.n119 B.n118 59.5399
R2043 B.n258 B.n116 59.5399
R2044 B.n496 B.n495 59.5399
R2045 B.n639 B.n493 59.5399
R2046 B.n759 B.n422 58.9903
R2047 B.n864 B.n44 58.9903
R2048 B.n118 B.n117 51.0066
R2049 B.n116 B.n115 51.0066
R2050 B.n495 B.n494 51.0066
R2051 B.n493 B.n492 51.0066
R2052 B.n763 B.n762 31.6883
R2053 B.n498 B.n420 31.6883
R2054 B.n862 B.n861 31.6883
R2055 B.n868 B.n867 31.6883
R2056 B.n766 B.n422 31.0959
R2057 B.n766 B.n418 31.0959
R2058 B.n772 B.n418 31.0959
R2059 B.n772 B.n414 31.0959
R2060 B.n778 B.n414 31.0959
R2061 B.n778 B.n410 31.0959
R2062 B.n784 B.n410 31.0959
R2063 B.n790 B.n406 31.0959
R2064 B.n790 B.n402 31.0959
R2065 B.n796 B.n402 31.0959
R2066 B.n796 B.n398 31.0959
R2067 B.n802 B.n398 31.0959
R2068 B.n802 B.n394 31.0959
R2069 B.n808 B.n394 31.0959
R2070 B.n808 B.n389 31.0959
R2071 B.n814 B.n389 31.0959
R2072 B.n814 B.n390 31.0959
R2073 B.n821 B.n382 31.0959
R2074 B.n827 B.n382 31.0959
R2075 B.n827 B.n4 31.0959
R2076 B.n914 B.n4 31.0959
R2077 B.n914 B.n913 31.0959
R2078 B.n913 B.n912 31.0959
R2079 B.n912 B.n8 31.0959
R2080 B.n12 B.n8 31.0959
R2081 B.n905 B.n12 31.0959
R2082 B.n904 B.n903 31.0959
R2083 B.n903 B.n16 31.0959
R2084 B.n897 B.n16 31.0959
R2085 B.n897 B.n896 31.0959
R2086 B.n896 B.n895 31.0959
R2087 B.n895 B.n23 31.0959
R2088 B.n889 B.n23 31.0959
R2089 B.n889 B.n888 31.0959
R2090 B.n888 B.n887 31.0959
R2091 B.n887 B.n30 31.0959
R2092 B.n881 B.n880 31.0959
R2093 B.n880 B.n879 31.0959
R2094 B.n879 B.n37 31.0959
R2095 B.n873 B.n37 31.0959
R2096 B.n873 B.n872 31.0959
R2097 B.n872 B.n871 31.0959
R2098 B.n871 B.n44 31.0959
R2099 B.n821 B.t1 30.1813
R2100 B.n905 B.t0 30.1813
R2101 B.t3 B.n406 28.3522
R2102 B.t7 B.n30 28.3522
R2103 B B.n917 18.0485
R2104 B.n764 B.n763 10.6151
R2105 B.n764 B.n416 10.6151
R2106 B.n774 B.n416 10.6151
R2107 B.n775 B.n774 10.6151
R2108 B.n776 B.n775 10.6151
R2109 B.n776 B.n408 10.6151
R2110 B.n786 B.n408 10.6151
R2111 B.n787 B.n786 10.6151
R2112 B.n788 B.n787 10.6151
R2113 B.n788 B.n400 10.6151
R2114 B.n798 B.n400 10.6151
R2115 B.n799 B.n798 10.6151
R2116 B.n800 B.n799 10.6151
R2117 B.n800 B.n392 10.6151
R2118 B.n810 B.n392 10.6151
R2119 B.n811 B.n810 10.6151
R2120 B.n812 B.n811 10.6151
R2121 B.n812 B.n384 10.6151
R2122 B.n823 B.n384 10.6151
R2123 B.n824 B.n823 10.6151
R2124 B.n825 B.n824 10.6151
R2125 B.n825 B.n0 10.6151
R2126 B.n762 B.n424 10.6151
R2127 B.n757 B.n424 10.6151
R2128 B.n757 B.n756 10.6151
R2129 B.n756 B.n755 10.6151
R2130 B.n755 B.n752 10.6151
R2131 B.n752 B.n751 10.6151
R2132 B.n751 B.n748 10.6151
R2133 B.n748 B.n747 10.6151
R2134 B.n747 B.n744 10.6151
R2135 B.n744 B.n743 10.6151
R2136 B.n743 B.n740 10.6151
R2137 B.n740 B.n739 10.6151
R2138 B.n739 B.n736 10.6151
R2139 B.n736 B.n735 10.6151
R2140 B.n735 B.n732 10.6151
R2141 B.n732 B.n731 10.6151
R2142 B.n731 B.n728 10.6151
R2143 B.n728 B.n727 10.6151
R2144 B.n727 B.n724 10.6151
R2145 B.n724 B.n723 10.6151
R2146 B.n723 B.n720 10.6151
R2147 B.n720 B.n719 10.6151
R2148 B.n719 B.n716 10.6151
R2149 B.n716 B.n715 10.6151
R2150 B.n715 B.n712 10.6151
R2151 B.n712 B.n711 10.6151
R2152 B.n711 B.n708 10.6151
R2153 B.n708 B.n707 10.6151
R2154 B.n707 B.n704 10.6151
R2155 B.n704 B.n703 10.6151
R2156 B.n703 B.n700 10.6151
R2157 B.n700 B.n699 10.6151
R2158 B.n699 B.n696 10.6151
R2159 B.n696 B.n695 10.6151
R2160 B.n695 B.n692 10.6151
R2161 B.n692 B.n691 10.6151
R2162 B.n691 B.n688 10.6151
R2163 B.n688 B.n687 10.6151
R2164 B.n687 B.n684 10.6151
R2165 B.n684 B.n683 10.6151
R2166 B.n683 B.n680 10.6151
R2167 B.n680 B.n679 10.6151
R2168 B.n679 B.n676 10.6151
R2169 B.n676 B.n675 10.6151
R2170 B.n675 B.n672 10.6151
R2171 B.n672 B.n671 10.6151
R2172 B.n671 B.n668 10.6151
R2173 B.n668 B.n667 10.6151
R2174 B.n667 B.n664 10.6151
R2175 B.n664 B.n663 10.6151
R2176 B.n663 B.n660 10.6151
R2177 B.n660 B.n659 10.6151
R2178 B.n659 B.n656 10.6151
R2179 B.n656 B.n655 10.6151
R2180 B.n655 B.n652 10.6151
R2181 B.n652 B.n651 10.6151
R2182 B.n651 B.n648 10.6151
R2183 B.n648 B.n647 10.6151
R2184 B.n647 B.n644 10.6151
R2185 B.n644 B.n643 10.6151
R2186 B.n643 B.n640 10.6151
R2187 B.n638 B.n635 10.6151
R2188 B.n635 B.n634 10.6151
R2189 B.n634 B.n631 10.6151
R2190 B.n631 B.n630 10.6151
R2191 B.n630 B.n627 10.6151
R2192 B.n627 B.n626 10.6151
R2193 B.n626 B.n623 10.6151
R2194 B.n623 B.n622 10.6151
R2195 B.n619 B.n618 10.6151
R2196 B.n618 B.n615 10.6151
R2197 B.n615 B.n614 10.6151
R2198 B.n614 B.n611 10.6151
R2199 B.n611 B.n610 10.6151
R2200 B.n610 B.n607 10.6151
R2201 B.n607 B.n606 10.6151
R2202 B.n606 B.n603 10.6151
R2203 B.n603 B.n602 10.6151
R2204 B.n602 B.n599 10.6151
R2205 B.n599 B.n598 10.6151
R2206 B.n598 B.n595 10.6151
R2207 B.n595 B.n594 10.6151
R2208 B.n594 B.n591 10.6151
R2209 B.n591 B.n590 10.6151
R2210 B.n590 B.n587 10.6151
R2211 B.n587 B.n586 10.6151
R2212 B.n586 B.n583 10.6151
R2213 B.n583 B.n582 10.6151
R2214 B.n582 B.n579 10.6151
R2215 B.n579 B.n578 10.6151
R2216 B.n578 B.n575 10.6151
R2217 B.n575 B.n574 10.6151
R2218 B.n574 B.n571 10.6151
R2219 B.n571 B.n570 10.6151
R2220 B.n570 B.n567 10.6151
R2221 B.n567 B.n566 10.6151
R2222 B.n566 B.n563 10.6151
R2223 B.n563 B.n562 10.6151
R2224 B.n562 B.n559 10.6151
R2225 B.n559 B.n558 10.6151
R2226 B.n558 B.n555 10.6151
R2227 B.n555 B.n554 10.6151
R2228 B.n554 B.n551 10.6151
R2229 B.n551 B.n550 10.6151
R2230 B.n550 B.n547 10.6151
R2231 B.n547 B.n546 10.6151
R2232 B.n546 B.n543 10.6151
R2233 B.n543 B.n542 10.6151
R2234 B.n542 B.n539 10.6151
R2235 B.n539 B.n538 10.6151
R2236 B.n538 B.n535 10.6151
R2237 B.n535 B.n534 10.6151
R2238 B.n534 B.n531 10.6151
R2239 B.n531 B.n530 10.6151
R2240 B.n530 B.n527 10.6151
R2241 B.n527 B.n526 10.6151
R2242 B.n526 B.n523 10.6151
R2243 B.n523 B.n522 10.6151
R2244 B.n522 B.n519 10.6151
R2245 B.n519 B.n518 10.6151
R2246 B.n518 B.n515 10.6151
R2247 B.n515 B.n514 10.6151
R2248 B.n514 B.n511 10.6151
R2249 B.n511 B.n510 10.6151
R2250 B.n510 B.n507 10.6151
R2251 B.n507 B.n506 10.6151
R2252 B.n506 B.n503 10.6151
R2253 B.n503 B.n502 10.6151
R2254 B.n502 B.n499 10.6151
R2255 B.n499 B.n498 10.6151
R2256 B.n768 B.n420 10.6151
R2257 B.n769 B.n768 10.6151
R2258 B.n770 B.n769 10.6151
R2259 B.n770 B.n412 10.6151
R2260 B.n780 B.n412 10.6151
R2261 B.n781 B.n780 10.6151
R2262 B.n782 B.n781 10.6151
R2263 B.n782 B.n404 10.6151
R2264 B.n792 B.n404 10.6151
R2265 B.n793 B.n792 10.6151
R2266 B.n794 B.n793 10.6151
R2267 B.n794 B.n396 10.6151
R2268 B.n804 B.n396 10.6151
R2269 B.n805 B.n804 10.6151
R2270 B.n806 B.n805 10.6151
R2271 B.n806 B.n387 10.6151
R2272 B.n816 B.n387 10.6151
R2273 B.n817 B.n816 10.6151
R2274 B.n819 B.n817 10.6151
R2275 B.n819 B.n818 10.6151
R2276 B.n818 B.n380 10.6151
R2277 B.n830 B.n380 10.6151
R2278 B.n831 B.n830 10.6151
R2279 B.n832 B.n831 10.6151
R2280 B.n833 B.n832 10.6151
R2281 B.n834 B.n833 10.6151
R2282 B.n837 B.n834 10.6151
R2283 B.n838 B.n837 10.6151
R2284 B.n839 B.n838 10.6151
R2285 B.n840 B.n839 10.6151
R2286 B.n842 B.n840 10.6151
R2287 B.n843 B.n842 10.6151
R2288 B.n844 B.n843 10.6151
R2289 B.n845 B.n844 10.6151
R2290 B.n847 B.n845 10.6151
R2291 B.n848 B.n847 10.6151
R2292 B.n849 B.n848 10.6151
R2293 B.n850 B.n849 10.6151
R2294 B.n852 B.n850 10.6151
R2295 B.n853 B.n852 10.6151
R2296 B.n854 B.n853 10.6151
R2297 B.n855 B.n854 10.6151
R2298 B.n857 B.n855 10.6151
R2299 B.n858 B.n857 10.6151
R2300 B.n859 B.n858 10.6151
R2301 B.n860 B.n859 10.6151
R2302 B.n861 B.n860 10.6151
R2303 B.n909 B.n1 10.6151
R2304 B.n909 B.n908 10.6151
R2305 B.n908 B.n907 10.6151
R2306 B.n907 B.n10 10.6151
R2307 B.n901 B.n10 10.6151
R2308 B.n901 B.n900 10.6151
R2309 B.n900 B.n899 10.6151
R2310 B.n899 B.n18 10.6151
R2311 B.n893 B.n18 10.6151
R2312 B.n893 B.n892 10.6151
R2313 B.n892 B.n891 10.6151
R2314 B.n891 B.n25 10.6151
R2315 B.n885 B.n25 10.6151
R2316 B.n885 B.n884 10.6151
R2317 B.n884 B.n883 10.6151
R2318 B.n883 B.n32 10.6151
R2319 B.n877 B.n32 10.6151
R2320 B.n877 B.n876 10.6151
R2321 B.n876 B.n875 10.6151
R2322 B.n875 B.n39 10.6151
R2323 B.n869 B.n39 10.6151
R2324 B.n869 B.n868 10.6151
R2325 B.n867 B.n46 10.6151
R2326 B.n121 B.n46 10.6151
R2327 B.n122 B.n121 10.6151
R2328 B.n125 B.n122 10.6151
R2329 B.n126 B.n125 10.6151
R2330 B.n129 B.n126 10.6151
R2331 B.n130 B.n129 10.6151
R2332 B.n133 B.n130 10.6151
R2333 B.n134 B.n133 10.6151
R2334 B.n137 B.n134 10.6151
R2335 B.n138 B.n137 10.6151
R2336 B.n141 B.n138 10.6151
R2337 B.n142 B.n141 10.6151
R2338 B.n145 B.n142 10.6151
R2339 B.n146 B.n145 10.6151
R2340 B.n149 B.n146 10.6151
R2341 B.n150 B.n149 10.6151
R2342 B.n153 B.n150 10.6151
R2343 B.n154 B.n153 10.6151
R2344 B.n157 B.n154 10.6151
R2345 B.n158 B.n157 10.6151
R2346 B.n161 B.n158 10.6151
R2347 B.n162 B.n161 10.6151
R2348 B.n165 B.n162 10.6151
R2349 B.n166 B.n165 10.6151
R2350 B.n169 B.n166 10.6151
R2351 B.n170 B.n169 10.6151
R2352 B.n173 B.n170 10.6151
R2353 B.n174 B.n173 10.6151
R2354 B.n177 B.n174 10.6151
R2355 B.n178 B.n177 10.6151
R2356 B.n181 B.n178 10.6151
R2357 B.n182 B.n181 10.6151
R2358 B.n185 B.n182 10.6151
R2359 B.n186 B.n185 10.6151
R2360 B.n189 B.n186 10.6151
R2361 B.n190 B.n189 10.6151
R2362 B.n193 B.n190 10.6151
R2363 B.n194 B.n193 10.6151
R2364 B.n197 B.n194 10.6151
R2365 B.n198 B.n197 10.6151
R2366 B.n201 B.n198 10.6151
R2367 B.n202 B.n201 10.6151
R2368 B.n205 B.n202 10.6151
R2369 B.n206 B.n205 10.6151
R2370 B.n209 B.n206 10.6151
R2371 B.n210 B.n209 10.6151
R2372 B.n213 B.n210 10.6151
R2373 B.n214 B.n213 10.6151
R2374 B.n217 B.n214 10.6151
R2375 B.n218 B.n217 10.6151
R2376 B.n221 B.n218 10.6151
R2377 B.n222 B.n221 10.6151
R2378 B.n225 B.n222 10.6151
R2379 B.n226 B.n225 10.6151
R2380 B.n229 B.n226 10.6151
R2381 B.n230 B.n229 10.6151
R2382 B.n233 B.n230 10.6151
R2383 B.n234 B.n233 10.6151
R2384 B.n237 B.n234 10.6151
R2385 B.n238 B.n237 10.6151
R2386 B.n242 B.n241 10.6151
R2387 B.n245 B.n242 10.6151
R2388 B.n246 B.n245 10.6151
R2389 B.n249 B.n246 10.6151
R2390 B.n250 B.n249 10.6151
R2391 B.n253 B.n250 10.6151
R2392 B.n254 B.n253 10.6151
R2393 B.n257 B.n254 10.6151
R2394 B.n262 B.n259 10.6151
R2395 B.n263 B.n262 10.6151
R2396 B.n266 B.n263 10.6151
R2397 B.n267 B.n266 10.6151
R2398 B.n270 B.n267 10.6151
R2399 B.n271 B.n270 10.6151
R2400 B.n274 B.n271 10.6151
R2401 B.n275 B.n274 10.6151
R2402 B.n278 B.n275 10.6151
R2403 B.n279 B.n278 10.6151
R2404 B.n282 B.n279 10.6151
R2405 B.n283 B.n282 10.6151
R2406 B.n286 B.n283 10.6151
R2407 B.n287 B.n286 10.6151
R2408 B.n290 B.n287 10.6151
R2409 B.n291 B.n290 10.6151
R2410 B.n294 B.n291 10.6151
R2411 B.n295 B.n294 10.6151
R2412 B.n298 B.n295 10.6151
R2413 B.n299 B.n298 10.6151
R2414 B.n302 B.n299 10.6151
R2415 B.n303 B.n302 10.6151
R2416 B.n306 B.n303 10.6151
R2417 B.n307 B.n306 10.6151
R2418 B.n310 B.n307 10.6151
R2419 B.n311 B.n310 10.6151
R2420 B.n314 B.n311 10.6151
R2421 B.n315 B.n314 10.6151
R2422 B.n318 B.n315 10.6151
R2423 B.n319 B.n318 10.6151
R2424 B.n322 B.n319 10.6151
R2425 B.n323 B.n322 10.6151
R2426 B.n326 B.n323 10.6151
R2427 B.n327 B.n326 10.6151
R2428 B.n330 B.n327 10.6151
R2429 B.n331 B.n330 10.6151
R2430 B.n334 B.n331 10.6151
R2431 B.n335 B.n334 10.6151
R2432 B.n338 B.n335 10.6151
R2433 B.n339 B.n338 10.6151
R2434 B.n342 B.n339 10.6151
R2435 B.n343 B.n342 10.6151
R2436 B.n346 B.n343 10.6151
R2437 B.n347 B.n346 10.6151
R2438 B.n350 B.n347 10.6151
R2439 B.n351 B.n350 10.6151
R2440 B.n354 B.n351 10.6151
R2441 B.n355 B.n354 10.6151
R2442 B.n358 B.n355 10.6151
R2443 B.n359 B.n358 10.6151
R2444 B.n362 B.n359 10.6151
R2445 B.n363 B.n362 10.6151
R2446 B.n366 B.n363 10.6151
R2447 B.n367 B.n366 10.6151
R2448 B.n370 B.n367 10.6151
R2449 B.n371 B.n370 10.6151
R2450 B.n374 B.n371 10.6151
R2451 B.n375 B.n374 10.6151
R2452 B.n378 B.n375 10.6151
R2453 B.n379 B.n378 10.6151
R2454 B.n862 B.n379 10.6151
R2455 B.n917 B.n0 8.11757
R2456 B.n917 B.n1 8.11757
R2457 B.n639 B.n638 6.5566
R2458 B.n622 B.n496 6.5566
R2459 B.n241 B.n119 6.5566
R2460 B.n258 B.n257 6.5566
R2461 B.n640 B.n639 4.05904
R2462 B.n619 B.n496 4.05904
R2463 B.n238 B.n119 4.05904
R2464 B.n259 B.n258 4.05904
R2465 B.n784 B.t3 2.74421
R2466 B.n881 B.t7 2.74421
R2467 B.n390 B.t1 0.915071
R2468 B.t0 B.n904 0.915071
R2469 VN VN.t1 295.002
R2470 VN VN.t0 246.244
R2471 VDD2.n205 VDD2.n204 289.615
R2472 VDD2.n102 VDD2.n101 289.615
R2473 VDD2.n204 VDD2.n203 185
R2474 VDD2.n105 VDD2.n104 185
R2475 VDD2.n198 VDD2.n197 185
R2476 VDD2.n196 VDD2.n195 185
R2477 VDD2.n109 VDD2.n108 185
R2478 VDD2.n190 VDD2.n189 185
R2479 VDD2.n188 VDD2.n187 185
R2480 VDD2.n113 VDD2.n112 185
R2481 VDD2.n182 VDD2.n181 185
R2482 VDD2.n180 VDD2.n179 185
R2483 VDD2.n117 VDD2.n116 185
R2484 VDD2.n174 VDD2.n173 185
R2485 VDD2.n172 VDD2.n171 185
R2486 VDD2.n121 VDD2.n120 185
R2487 VDD2.n166 VDD2.n165 185
R2488 VDD2.n164 VDD2.n163 185
R2489 VDD2.n125 VDD2.n124 185
R2490 VDD2.n129 VDD2.n127 185
R2491 VDD2.n158 VDD2.n157 185
R2492 VDD2.n156 VDD2.n155 185
R2493 VDD2.n131 VDD2.n130 185
R2494 VDD2.n150 VDD2.n149 185
R2495 VDD2.n148 VDD2.n147 185
R2496 VDD2.n135 VDD2.n134 185
R2497 VDD2.n142 VDD2.n141 185
R2498 VDD2.n140 VDD2.n139 185
R2499 VDD2.n35 VDD2.n34 185
R2500 VDD2.n37 VDD2.n36 185
R2501 VDD2.n30 VDD2.n29 185
R2502 VDD2.n43 VDD2.n42 185
R2503 VDD2.n45 VDD2.n44 185
R2504 VDD2.n26 VDD2.n25 185
R2505 VDD2.n52 VDD2.n51 185
R2506 VDD2.n53 VDD2.n24 185
R2507 VDD2.n55 VDD2.n54 185
R2508 VDD2.n22 VDD2.n21 185
R2509 VDD2.n61 VDD2.n60 185
R2510 VDD2.n63 VDD2.n62 185
R2511 VDD2.n18 VDD2.n17 185
R2512 VDD2.n69 VDD2.n68 185
R2513 VDD2.n71 VDD2.n70 185
R2514 VDD2.n14 VDD2.n13 185
R2515 VDD2.n77 VDD2.n76 185
R2516 VDD2.n79 VDD2.n78 185
R2517 VDD2.n10 VDD2.n9 185
R2518 VDD2.n85 VDD2.n84 185
R2519 VDD2.n87 VDD2.n86 185
R2520 VDD2.n6 VDD2.n5 185
R2521 VDD2.n93 VDD2.n92 185
R2522 VDD2.n95 VDD2.n94 185
R2523 VDD2.n2 VDD2.n1 185
R2524 VDD2.n101 VDD2.n100 185
R2525 VDD2.n138 VDD2.t0 149.524
R2526 VDD2.n33 VDD2.t1 149.524
R2527 VDD2.n204 VDD2.n104 104.615
R2528 VDD2.n197 VDD2.n104 104.615
R2529 VDD2.n197 VDD2.n196 104.615
R2530 VDD2.n196 VDD2.n108 104.615
R2531 VDD2.n189 VDD2.n108 104.615
R2532 VDD2.n189 VDD2.n188 104.615
R2533 VDD2.n188 VDD2.n112 104.615
R2534 VDD2.n181 VDD2.n112 104.615
R2535 VDD2.n181 VDD2.n180 104.615
R2536 VDD2.n180 VDD2.n116 104.615
R2537 VDD2.n173 VDD2.n116 104.615
R2538 VDD2.n173 VDD2.n172 104.615
R2539 VDD2.n172 VDD2.n120 104.615
R2540 VDD2.n165 VDD2.n120 104.615
R2541 VDD2.n165 VDD2.n164 104.615
R2542 VDD2.n164 VDD2.n124 104.615
R2543 VDD2.n129 VDD2.n124 104.615
R2544 VDD2.n157 VDD2.n129 104.615
R2545 VDD2.n157 VDD2.n156 104.615
R2546 VDD2.n156 VDD2.n130 104.615
R2547 VDD2.n149 VDD2.n130 104.615
R2548 VDD2.n149 VDD2.n148 104.615
R2549 VDD2.n148 VDD2.n134 104.615
R2550 VDD2.n141 VDD2.n134 104.615
R2551 VDD2.n141 VDD2.n140 104.615
R2552 VDD2.n36 VDD2.n35 104.615
R2553 VDD2.n36 VDD2.n29 104.615
R2554 VDD2.n43 VDD2.n29 104.615
R2555 VDD2.n44 VDD2.n43 104.615
R2556 VDD2.n44 VDD2.n25 104.615
R2557 VDD2.n52 VDD2.n25 104.615
R2558 VDD2.n53 VDD2.n52 104.615
R2559 VDD2.n54 VDD2.n53 104.615
R2560 VDD2.n54 VDD2.n21 104.615
R2561 VDD2.n61 VDD2.n21 104.615
R2562 VDD2.n62 VDD2.n61 104.615
R2563 VDD2.n62 VDD2.n17 104.615
R2564 VDD2.n69 VDD2.n17 104.615
R2565 VDD2.n70 VDD2.n69 104.615
R2566 VDD2.n70 VDD2.n13 104.615
R2567 VDD2.n77 VDD2.n13 104.615
R2568 VDD2.n78 VDD2.n77 104.615
R2569 VDD2.n78 VDD2.n9 104.615
R2570 VDD2.n85 VDD2.n9 104.615
R2571 VDD2.n86 VDD2.n85 104.615
R2572 VDD2.n86 VDD2.n5 104.615
R2573 VDD2.n93 VDD2.n5 104.615
R2574 VDD2.n94 VDD2.n93 104.615
R2575 VDD2.n94 VDD2.n1 104.615
R2576 VDD2.n101 VDD2.n1 104.615
R2577 VDD2.n206 VDD2.n102 96.3508
R2578 VDD2.n140 VDD2.t0 52.3082
R2579 VDD2.n35 VDD2.t1 52.3082
R2580 VDD2.n206 VDD2.n205 51.9672
R2581 VDD2.n127 VDD2.n125 13.1884
R2582 VDD2.n55 VDD2.n22 13.1884
R2583 VDD2.n203 VDD2.n103 12.8005
R2584 VDD2.n163 VDD2.n162 12.8005
R2585 VDD2.n159 VDD2.n158 12.8005
R2586 VDD2.n56 VDD2.n24 12.8005
R2587 VDD2.n60 VDD2.n59 12.8005
R2588 VDD2.n100 VDD2.n0 12.8005
R2589 VDD2.n202 VDD2.n105 12.0247
R2590 VDD2.n166 VDD2.n123 12.0247
R2591 VDD2.n155 VDD2.n128 12.0247
R2592 VDD2.n51 VDD2.n50 12.0247
R2593 VDD2.n63 VDD2.n20 12.0247
R2594 VDD2.n99 VDD2.n2 12.0247
R2595 VDD2.n199 VDD2.n198 11.249
R2596 VDD2.n167 VDD2.n121 11.249
R2597 VDD2.n154 VDD2.n131 11.249
R2598 VDD2.n49 VDD2.n26 11.249
R2599 VDD2.n64 VDD2.n18 11.249
R2600 VDD2.n96 VDD2.n95 11.249
R2601 VDD2.n195 VDD2.n107 10.4732
R2602 VDD2.n171 VDD2.n170 10.4732
R2603 VDD2.n151 VDD2.n150 10.4732
R2604 VDD2.n46 VDD2.n45 10.4732
R2605 VDD2.n68 VDD2.n67 10.4732
R2606 VDD2.n92 VDD2.n4 10.4732
R2607 VDD2.n139 VDD2.n138 10.2747
R2608 VDD2.n34 VDD2.n33 10.2747
R2609 VDD2.n194 VDD2.n109 9.69747
R2610 VDD2.n174 VDD2.n119 9.69747
R2611 VDD2.n147 VDD2.n133 9.69747
R2612 VDD2.n42 VDD2.n28 9.69747
R2613 VDD2.n71 VDD2.n16 9.69747
R2614 VDD2.n91 VDD2.n6 9.69747
R2615 VDD2.n201 VDD2.n103 9.45567
R2616 VDD2.n98 VDD2.n0 9.45567
R2617 VDD2.n202 VDD2.n201 9.3005
R2618 VDD2.n200 VDD2.n199 9.3005
R2619 VDD2.n107 VDD2.n106 9.3005
R2620 VDD2.n194 VDD2.n193 9.3005
R2621 VDD2.n192 VDD2.n191 9.3005
R2622 VDD2.n111 VDD2.n110 9.3005
R2623 VDD2.n186 VDD2.n185 9.3005
R2624 VDD2.n184 VDD2.n183 9.3005
R2625 VDD2.n115 VDD2.n114 9.3005
R2626 VDD2.n178 VDD2.n177 9.3005
R2627 VDD2.n176 VDD2.n175 9.3005
R2628 VDD2.n119 VDD2.n118 9.3005
R2629 VDD2.n170 VDD2.n169 9.3005
R2630 VDD2.n168 VDD2.n167 9.3005
R2631 VDD2.n123 VDD2.n122 9.3005
R2632 VDD2.n162 VDD2.n161 9.3005
R2633 VDD2.n160 VDD2.n159 9.3005
R2634 VDD2.n128 VDD2.n126 9.3005
R2635 VDD2.n154 VDD2.n153 9.3005
R2636 VDD2.n152 VDD2.n151 9.3005
R2637 VDD2.n133 VDD2.n132 9.3005
R2638 VDD2.n146 VDD2.n145 9.3005
R2639 VDD2.n144 VDD2.n143 9.3005
R2640 VDD2.n137 VDD2.n136 9.3005
R2641 VDD2.n81 VDD2.n80 9.3005
R2642 VDD2.n83 VDD2.n82 9.3005
R2643 VDD2.n8 VDD2.n7 9.3005
R2644 VDD2.n89 VDD2.n88 9.3005
R2645 VDD2.n91 VDD2.n90 9.3005
R2646 VDD2.n4 VDD2.n3 9.3005
R2647 VDD2.n97 VDD2.n96 9.3005
R2648 VDD2.n99 VDD2.n98 9.3005
R2649 VDD2.n75 VDD2.n74 9.3005
R2650 VDD2.n73 VDD2.n72 9.3005
R2651 VDD2.n16 VDD2.n15 9.3005
R2652 VDD2.n67 VDD2.n66 9.3005
R2653 VDD2.n65 VDD2.n64 9.3005
R2654 VDD2.n20 VDD2.n19 9.3005
R2655 VDD2.n59 VDD2.n58 9.3005
R2656 VDD2.n32 VDD2.n31 9.3005
R2657 VDD2.n39 VDD2.n38 9.3005
R2658 VDD2.n41 VDD2.n40 9.3005
R2659 VDD2.n28 VDD2.n27 9.3005
R2660 VDD2.n47 VDD2.n46 9.3005
R2661 VDD2.n49 VDD2.n48 9.3005
R2662 VDD2.n50 VDD2.n23 9.3005
R2663 VDD2.n57 VDD2.n56 9.3005
R2664 VDD2.n12 VDD2.n11 9.3005
R2665 VDD2.n191 VDD2.n190 8.92171
R2666 VDD2.n175 VDD2.n117 8.92171
R2667 VDD2.n146 VDD2.n135 8.92171
R2668 VDD2.n41 VDD2.n30 8.92171
R2669 VDD2.n72 VDD2.n14 8.92171
R2670 VDD2.n88 VDD2.n87 8.92171
R2671 VDD2.n187 VDD2.n111 8.14595
R2672 VDD2.n179 VDD2.n178 8.14595
R2673 VDD2.n143 VDD2.n142 8.14595
R2674 VDD2.n38 VDD2.n37 8.14595
R2675 VDD2.n76 VDD2.n75 8.14595
R2676 VDD2.n84 VDD2.n8 8.14595
R2677 VDD2.n186 VDD2.n113 7.3702
R2678 VDD2.n182 VDD2.n115 7.3702
R2679 VDD2.n139 VDD2.n137 7.3702
R2680 VDD2.n34 VDD2.n32 7.3702
R2681 VDD2.n79 VDD2.n12 7.3702
R2682 VDD2.n83 VDD2.n10 7.3702
R2683 VDD2.n183 VDD2.n113 6.59444
R2684 VDD2.n183 VDD2.n182 6.59444
R2685 VDD2.n80 VDD2.n79 6.59444
R2686 VDD2.n80 VDD2.n10 6.59444
R2687 VDD2.n187 VDD2.n186 5.81868
R2688 VDD2.n179 VDD2.n115 5.81868
R2689 VDD2.n142 VDD2.n137 5.81868
R2690 VDD2.n37 VDD2.n32 5.81868
R2691 VDD2.n76 VDD2.n12 5.81868
R2692 VDD2.n84 VDD2.n83 5.81868
R2693 VDD2.n190 VDD2.n111 5.04292
R2694 VDD2.n178 VDD2.n117 5.04292
R2695 VDD2.n143 VDD2.n135 5.04292
R2696 VDD2.n38 VDD2.n30 5.04292
R2697 VDD2.n75 VDD2.n14 5.04292
R2698 VDD2.n87 VDD2.n8 5.04292
R2699 VDD2.n191 VDD2.n109 4.26717
R2700 VDD2.n175 VDD2.n174 4.26717
R2701 VDD2.n147 VDD2.n146 4.26717
R2702 VDD2.n42 VDD2.n41 4.26717
R2703 VDD2.n72 VDD2.n71 4.26717
R2704 VDD2.n88 VDD2.n6 4.26717
R2705 VDD2.n195 VDD2.n194 3.49141
R2706 VDD2.n171 VDD2.n119 3.49141
R2707 VDD2.n150 VDD2.n133 3.49141
R2708 VDD2.n45 VDD2.n28 3.49141
R2709 VDD2.n68 VDD2.n16 3.49141
R2710 VDD2.n92 VDD2.n91 3.49141
R2711 VDD2.n33 VDD2.n31 2.84303
R2712 VDD2.n138 VDD2.n136 2.84303
R2713 VDD2.n198 VDD2.n107 2.71565
R2714 VDD2.n170 VDD2.n121 2.71565
R2715 VDD2.n151 VDD2.n131 2.71565
R2716 VDD2.n46 VDD2.n26 2.71565
R2717 VDD2.n67 VDD2.n18 2.71565
R2718 VDD2.n95 VDD2.n4 2.71565
R2719 VDD2.n199 VDD2.n105 1.93989
R2720 VDD2.n167 VDD2.n166 1.93989
R2721 VDD2.n155 VDD2.n154 1.93989
R2722 VDD2.n51 VDD2.n49 1.93989
R2723 VDD2.n64 VDD2.n63 1.93989
R2724 VDD2.n96 VDD2.n2 1.93989
R2725 VDD2.n203 VDD2.n202 1.16414
R2726 VDD2.n163 VDD2.n123 1.16414
R2727 VDD2.n158 VDD2.n128 1.16414
R2728 VDD2.n50 VDD2.n24 1.16414
R2729 VDD2.n60 VDD2.n20 1.16414
R2730 VDD2.n100 VDD2.n99 1.16414
R2731 VDD2 VDD2.n206 0.6255
R2732 VDD2.n205 VDD2.n103 0.388379
R2733 VDD2.n162 VDD2.n125 0.388379
R2734 VDD2.n159 VDD2.n127 0.388379
R2735 VDD2.n56 VDD2.n55 0.388379
R2736 VDD2.n59 VDD2.n22 0.388379
R2737 VDD2.n102 VDD2.n0 0.388379
R2738 VDD2.n201 VDD2.n200 0.155672
R2739 VDD2.n200 VDD2.n106 0.155672
R2740 VDD2.n193 VDD2.n106 0.155672
R2741 VDD2.n193 VDD2.n192 0.155672
R2742 VDD2.n192 VDD2.n110 0.155672
R2743 VDD2.n185 VDD2.n110 0.155672
R2744 VDD2.n185 VDD2.n184 0.155672
R2745 VDD2.n184 VDD2.n114 0.155672
R2746 VDD2.n177 VDD2.n114 0.155672
R2747 VDD2.n177 VDD2.n176 0.155672
R2748 VDD2.n176 VDD2.n118 0.155672
R2749 VDD2.n169 VDD2.n118 0.155672
R2750 VDD2.n169 VDD2.n168 0.155672
R2751 VDD2.n168 VDD2.n122 0.155672
R2752 VDD2.n161 VDD2.n122 0.155672
R2753 VDD2.n161 VDD2.n160 0.155672
R2754 VDD2.n160 VDD2.n126 0.155672
R2755 VDD2.n153 VDD2.n126 0.155672
R2756 VDD2.n153 VDD2.n152 0.155672
R2757 VDD2.n152 VDD2.n132 0.155672
R2758 VDD2.n145 VDD2.n132 0.155672
R2759 VDD2.n145 VDD2.n144 0.155672
R2760 VDD2.n144 VDD2.n136 0.155672
R2761 VDD2.n39 VDD2.n31 0.155672
R2762 VDD2.n40 VDD2.n39 0.155672
R2763 VDD2.n40 VDD2.n27 0.155672
R2764 VDD2.n47 VDD2.n27 0.155672
R2765 VDD2.n48 VDD2.n47 0.155672
R2766 VDD2.n48 VDD2.n23 0.155672
R2767 VDD2.n57 VDD2.n23 0.155672
R2768 VDD2.n58 VDD2.n57 0.155672
R2769 VDD2.n58 VDD2.n19 0.155672
R2770 VDD2.n65 VDD2.n19 0.155672
R2771 VDD2.n66 VDD2.n65 0.155672
R2772 VDD2.n66 VDD2.n15 0.155672
R2773 VDD2.n73 VDD2.n15 0.155672
R2774 VDD2.n74 VDD2.n73 0.155672
R2775 VDD2.n74 VDD2.n11 0.155672
R2776 VDD2.n81 VDD2.n11 0.155672
R2777 VDD2.n82 VDD2.n81 0.155672
R2778 VDD2.n82 VDD2.n7 0.155672
R2779 VDD2.n89 VDD2.n7 0.155672
R2780 VDD2.n90 VDD2.n89 0.155672
R2781 VDD2.n90 VDD2.n3 0.155672
R2782 VDD2.n97 VDD2.n3 0.155672
R2783 VDD2.n98 VDD2.n97 0.155672
C0 VDD1 VTAIL 6.86575f
C1 VDD1 VDD2 0.639638f
C2 VDD2 VTAIL 6.91223f
C3 VDD1 VN 0.14765f
C4 VN VTAIL 3.45935f
C5 VDD2 VN 4.126339f
C6 VDD1 VP 4.29543f
C7 VTAIL VP 3.47378f
C8 VDD2 VP 0.320738f
C9 VN VP 6.57469f
C10 VDD2 B 5.542786f
C11 VDD1 B 8.752629f
C12 VTAIL B 9.957382f
C13 VN B 12.0914f
C14 VP B 6.486495f
C15 VDD2.n0 B 0.011167f
C16 VDD2.n1 B 0.025177f
C17 VDD2.n2 B 0.011278f
C18 VDD2.n3 B 0.019822f
C19 VDD2.n4 B 0.010652f
C20 VDD2.n5 B 0.025177f
C21 VDD2.n6 B 0.011278f
C22 VDD2.n7 B 0.019822f
C23 VDD2.n8 B 0.010652f
C24 VDD2.n9 B 0.025177f
C25 VDD2.n10 B 0.011278f
C26 VDD2.n11 B 0.019822f
C27 VDD2.n12 B 0.010652f
C28 VDD2.n13 B 0.025177f
C29 VDD2.n14 B 0.011278f
C30 VDD2.n15 B 0.019822f
C31 VDD2.n16 B 0.010652f
C32 VDD2.n17 B 0.025177f
C33 VDD2.n18 B 0.011278f
C34 VDD2.n19 B 0.019822f
C35 VDD2.n20 B 0.010652f
C36 VDD2.n21 B 0.025177f
C37 VDD2.n22 B 0.010965f
C38 VDD2.n23 B 0.019822f
C39 VDD2.n24 B 0.011278f
C40 VDD2.n25 B 0.025177f
C41 VDD2.n26 B 0.011278f
C42 VDD2.n27 B 0.019822f
C43 VDD2.n28 B 0.010652f
C44 VDD2.n29 B 0.025177f
C45 VDD2.n30 B 0.011278f
C46 VDD2.n31 B 1.59776f
C47 VDD2.n32 B 0.010652f
C48 VDD2.t1 B 0.043245f
C49 VDD2.n33 B 0.194512f
C50 VDD2.n34 B 0.017798f
C51 VDD2.n35 B 0.018882f
C52 VDD2.n36 B 0.025177f
C53 VDD2.n37 B 0.011278f
C54 VDD2.n38 B 0.010652f
C55 VDD2.n39 B 0.019822f
C56 VDD2.n40 B 0.019822f
C57 VDD2.n41 B 0.010652f
C58 VDD2.n42 B 0.011278f
C59 VDD2.n43 B 0.025177f
C60 VDD2.n44 B 0.025177f
C61 VDD2.n45 B 0.011278f
C62 VDD2.n46 B 0.010652f
C63 VDD2.n47 B 0.019822f
C64 VDD2.n48 B 0.019822f
C65 VDD2.n49 B 0.010652f
C66 VDD2.n50 B 0.010652f
C67 VDD2.n51 B 0.011278f
C68 VDD2.n52 B 0.025177f
C69 VDD2.n53 B 0.025177f
C70 VDD2.n54 B 0.025177f
C71 VDD2.n55 B 0.010965f
C72 VDD2.n56 B 0.010652f
C73 VDD2.n57 B 0.019822f
C74 VDD2.n58 B 0.019822f
C75 VDD2.n59 B 0.010652f
C76 VDD2.n60 B 0.011278f
C77 VDD2.n61 B 0.025177f
C78 VDD2.n62 B 0.025177f
C79 VDD2.n63 B 0.011278f
C80 VDD2.n64 B 0.010652f
C81 VDD2.n65 B 0.019822f
C82 VDD2.n66 B 0.019822f
C83 VDD2.n67 B 0.010652f
C84 VDD2.n68 B 0.011278f
C85 VDD2.n69 B 0.025177f
C86 VDD2.n70 B 0.025177f
C87 VDD2.n71 B 0.011278f
C88 VDD2.n72 B 0.010652f
C89 VDD2.n73 B 0.019822f
C90 VDD2.n74 B 0.019822f
C91 VDD2.n75 B 0.010652f
C92 VDD2.n76 B 0.011278f
C93 VDD2.n77 B 0.025177f
C94 VDD2.n78 B 0.025177f
C95 VDD2.n79 B 0.011278f
C96 VDD2.n80 B 0.010652f
C97 VDD2.n81 B 0.019822f
C98 VDD2.n82 B 0.019822f
C99 VDD2.n83 B 0.010652f
C100 VDD2.n84 B 0.011278f
C101 VDD2.n85 B 0.025177f
C102 VDD2.n86 B 0.025177f
C103 VDD2.n87 B 0.011278f
C104 VDD2.n88 B 0.010652f
C105 VDD2.n89 B 0.019822f
C106 VDD2.n90 B 0.019822f
C107 VDD2.n91 B 0.010652f
C108 VDD2.n92 B 0.011278f
C109 VDD2.n93 B 0.025177f
C110 VDD2.n94 B 0.025177f
C111 VDD2.n95 B 0.011278f
C112 VDD2.n96 B 0.010652f
C113 VDD2.n97 B 0.019822f
C114 VDD2.n98 B 0.050692f
C115 VDD2.n99 B 0.010652f
C116 VDD2.n100 B 0.011278f
C117 VDD2.n101 B 0.051192f
C118 VDD2.n102 B 0.757991f
C119 VDD2.n103 B 0.011167f
C120 VDD2.n104 B 0.025177f
C121 VDD2.n105 B 0.011278f
C122 VDD2.n106 B 0.019822f
C123 VDD2.n107 B 0.010652f
C124 VDD2.n108 B 0.025177f
C125 VDD2.n109 B 0.011278f
C126 VDD2.n110 B 0.019822f
C127 VDD2.n111 B 0.010652f
C128 VDD2.n112 B 0.025177f
C129 VDD2.n113 B 0.011278f
C130 VDD2.n114 B 0.019822f
C131 VDD2.n115 B 0.010652f
C132 VDD2.n116 B 0.025177f
C133 VDD2.n117 B 0.011278f
C134 VDD2.n118 B 0.019822f
C135 VDD2.n119 B 0.010652f
C136 VDD2.n120 B 0.025177f
C137 VDD2.n121 B 0.011278f
C138 VDD2.n122 B 0.019822f
C139 VDD2.n123 B 0.010652f
C140 VDD2.n124 B 0.025177f
C141 VDD2.n125 B 0.010965f
C142 VDD2.n126 B 0.019822f
C143 VDD2.n127 B 0.010965f
C144 VDD2.n128 B 0.010652f
C145 VDD2.n129 B 0.025177f
C146 VDD2.n130 B 0.025177f
C147 VDD2.n131 B 0.011278f
C148 VDD2.n132 B 0.019822f
C149 VDD2.n133 B 0.010652f
C150 VDD2.n134 B 0.025177f
C151 VDD2.n135 B 0.011278f
C152 VDD2.n136 B 1.59776f
C153 VDD2.n137 B 0.010652f
C154 VDD2.t0 B 0.043245f
C155 VDD2.n138 B 0.194512f
C156 VDD2.n139 B 0.017798f
C157 VDD2.n140 B 0.018882f
C158 VDD2.n141 B 0.025177f
C159 VDD2.n142 B 0.011278f
C160 VDD2.n143 B 0.010652f
C161 VDD2.n144 B 0.019822f
C162 VDD2.n145 B 0.019822f
C163 VDD2.n146 B 0.010652f
C164 VDD2.n147 B 0.011278f
C165 VDD2.n148 B 0.025177f
C166 VDD2.n149 B 0.025177f
C167 VDD2.n150 B 0.011278f
C168 VDD2.n151 B 0.010652f
C169 VDD2.n152 B 0.019822f
C170 VDD2.n153 B 0.019822f
C171 VDD2.n154 B 0.010652f
C172 VDD2.n155 B 0.011278f
C173 VDD2.n156 B 0.025177f
C174 VDD2.n157 B 0.025177f
C175 VDD2.n158 B 0.011278f
C176 VDD2.n159 B 0.010652f
C177 VDD2.n160 B 0.019822f
C178 VDD2.n161 B 0.019822f
C179 VDD2.n162 B 0.010652f
C180 VDD2.n163 B 0.011278f
C181 VDD2.n164 B 0.025177f
C182 VDD2.n165 B 0.025177f
C183 VDD2.n166 B 0.011278f
C184 VDD2.n167 B 0.010652f
C185 VDD2.n168 B 0.019822f
C186 VDD2.n169 B 0.019822f
C187 VDD2.n170 B 0.010652f
C188 VDD2.n171 B 0.011278f
C189 VDD2.n172 B 0.025177f
C190 VDD2.n173 B 0.025177f
C191 VDD2.n174 B 0.011278f
C192 VDD2.n175 B 0.010652f
C193 VDD2.n176 B 0.019822f
C194 VDD2.n177 B 0.019822f
C195 VDD2.n178 B 0.010652f
C196 VDD2.n179 B 0.011278f
C197 VDD2.n180 B 0.025177f
C198 VDD2.n181 B 0.025177f
C199 VDD2.n182 B 0.011278f
C200 VDD2.n183 B 0.010652f
C201 VDD2.n184 B 0.019822f
C202 VDD2.n185 B 0.019822f
C203 VDD2.n186 B 0.010652f
C204 VDD2.n187 B 0.011278f
C205 VDD2.n188 B 0.025177f
C206 VDD2.n189 B 0.025177f
C207 VDD2.n190 B 0.011278f
C208 VDD2.n191 B 0.010652f
C209 VDD2.n192 B 0.019822f
C210 VDD2.n193 B 0.019822f
C211 VDD2.n194 B 0.010652f
C212 VDD2.n195 B 0.011278f
C213 VDD2.n196 B 0.025177f
C214 VDD2.n197 B 0.025177f
C215 VDD2.n198 B 0.011278f
C216 VDD2.n199 B 0.010652f
C217 VDD2.n200 B 0.019822f
C218 VDD2.n201 B 0.050692f
C219 VDD2.n202 B 0.010652f
C220 VDD2.n203 B 0.011278f
C221 VDD2.n204 B 0.051192f
C222 VDD2.n205 B 0.056606f
C223 VDD2.n206 B 2.94745f
C224 VN.t0 B 4.07262f
C225 VN.t1 B 4.57106f
C226 VDD1.n0 B 0.011294f
C227 VDD1.n1 B 0.025465f
C228 VDD1.n2 B 0.011407f
C229 VDD1.n3 B 0.020049f
C230 VDD1.n4 B 0.010774f
C231 VDD1.n5 B 0.025465f
C232 VDD1.n6 B 0.011407f
C233 VDD1.n7 B 0.020049f
C234 VDD1.n8 B 0.010774f
C235 VDD1.n9 B 0.025465f
C236 VDD1.n10 B 0.011407f
C237 VDD1.n11 B 0.020049f
C238 VDD1.n12 B 0.010774f
C239 VDD1.n13 B 0.025465f
C240 VDD1.n14 B 0.011407f
C241 VDD1.n15 B 0.020049f
C242 VDD1.n16 B 0.010774f
C243 VDD1.n17 B 0.025465f
C244 VDD1.n18 B 0.011407f
C245 VDD1.n19 B 0.020049f
C246 VDD1.n20 B 0.010774f
C247 VDD1.n21 B 0.025465f
C248 VDD1.n22 B 0.01109f
C249 VDD1.n23 B 0.020049f
C250 VDD1.n24 B 0.01109f
C251 VDD1.n25 B 0.010774f
C252 VDD1.n26 B 0.025465f
C253 VDD1.n27 B 0.025465f
C254 VDD1.n28 B 0.011407f
C255 VDD1.n29 B 0.020049f
C256 VDD1.n30 B 0.010774f
C257 VDD1.n31 B 0.025465f
C258 VDD1.n32 B 0.011407f
C259 VDD1.n33 B 1.61606f
C260 VDD1.n34 B 0.010774f
C261 VDD1.t1 B 0.04374f
C262 VDD1.n35 B 0.196739f
C263 VDD1.n36 B 0.018002f
C264 VDD1.n37 B 0.019099f
C265 VDD1.n38 B 0.025465f
C266 VDD1.n39 B 0.011407f
C267 VDD1.n40 B 0.010774f
C268 VDD1.n41 B 0.020049f
C269 VDD1.n42 B 0.020049f
C270 VDD1.n43 B 0.010774f
C271 VDD1.n44 B 0.011407f
C272 VDD1.n45 B 0.025465f
C273 VDD1.n46 B 0.025465f
C274 VDD1.n47 B 0.011407f
C275 VDD1.n48 B 0.010774f
C276 VDD1.n49 B 0.020049f
C277 VDD1.n50 B 0.020049f
C278 VDD1.n51 B 0.010774f
C279 VDD1.n52 B 0.011407f
C280 VDD1.n53 B 0.025465f
C281 VDD1.n54 B 0.025465f
C282 VDD1.n55 B 0.011407f
C283 VDD1.n56 B 0.010774f
C284 VDD1.n57 B 0.020049f
C285 VDD1.n58 B 0.020049f
C286 VDD1.n59 B 0.010774f
C287 VDD1.n60 B 0.011407f
C288 VDD1.n61 B 0.025465f
C289 VDD1.n62 B 0.025465f
C290 VDD1.n63 B 0.011407f
C291 VDD1.n64 B 0.010774f
C292 VDD1.n65 B 0.020049f
C293 VDD1.n66 B 0.020049f
C294 VDD1.n67 B 0.010774f
C295 VDD1.n68 B 0.011407f
C296 VDD1.n69 B 0.025465f
C297 VDD1.n70 B 0.025465f
C298 VDD1.n71 B 0.011407f
C299 VDD1.n72 B 0.010774f
C300 VDD1.n73 B 0.020049f
C301 VDD1.n74 B 0.020049f
C302 VDD1.n75 B 0.010774f
C303 VDD1.n76 B 0.011407f
C304 VDD1.n77 B 0.025465f
C305 VDD1.n78 B 0.025465f
C306 VDD1.n79 B 0.011407f
C307 VDD1.n80 B 0.010774f
C308 VDD1.n81 B 0.020049f
C309 VDD1.n82 B 0.020049f
C310 VDD1.n83 B 0.010774f
C311 VDD1.n84 B 0.011407f
C312 VDD1.n85 B 0.025465f
C313 VDD1.n86 B 0.025465f
C314 VDD1.n87 B 0.011407f
C315 VDD1.n88 B 0.010774f
C316 VDD1.n89 B 0.020049f
C317 VDD1.n90 B 0.020049f
C318 VDD1.n91 B 0.010774f
C319 VDD1.n92 B 0.011407f
C320 VDD1.n93 B 0.025465f
C321 VDD1.n94 B 0.025465f
C322 VDD1.n95 B 0.011407f
C323 VDD1.n96 B 0.010774f
C324 VDD1.n97 B 0.020049f
C325 VDD1.n98 B 0.051273f
C326 VDD1.n99 B 0.010774f
C327 VDD1.n100 B 0.011407f
C328 VDD1.n101 B 0.051778f
C329 VDD1.n102 B 0.058222f
C330 VDD1.n103 B 0.011294f
C331 VDD1.n104 B 0.025465f
C332 VDD1.n105 B 0.011407f
C333 VDD1.n106 B 0.020049f
C334 VDD1.n107 B 0.010774f
C335 VDD1.n108 B 0.025465f
C336 VDD1.n109 B 0.011407f
C337 VDD1.n110 B 0.020049f
C338 VDD1.n111 B 0.010774f
C339 VDD1.n112 B 0.025465f
C340 VDD1.n113 B 0.011407f
C341 VDD1.n114 B 0.020049f
C342 VDD1.n115 B 0.010774f
C343 VDD1.n116 B 0.025465f
C344 VDD1.n117 B 0.011407f
C345 VDD1.n118 B 0.020049f
C346 VDD1.n119 B 0.010774f
C347 VDD1.n120 B 0.025465f
C348 VDD1.n121 B 0.011407f
C349 VDD1.n122 B 0.020049f
C350 VDD1.n123 B 0.010774f
C351 VDD1.n124 B 0.025465f
C352 VDD1.n125 B 0.01109f
C353 VDD1.n126 B 0.020049f
C354 VDD1.n127 B 0.011407f
C355 VDD1.n128 B 0.025465f
C356 VDD1.n129 B 0.011407f
C357 VDD1.n130 B 0.020049f
C358 VDD1.n131 B 0.010774f
C359 VDD1.n132 B 0.025465f
C360 VDD1.n133 B 0.011407f
C361 VDD1.n134 B 1.61606f
C362 VDD1.n135 B 0.010774f
C363 VDD1.t0 B 0.04374f
C364 VDD1.n136 B 0.196739f
C365 VDD1.n137 B 0.018002f
C366 VDD1.n138 B 0.019099f
C367 VDD1.n139 B 0.025465f
C368 VDD1.n140 B 0.011407f
C369 VDD1.n141 B 0.010774f
C370 VDD1.n142 B 0.020049f
C371 VDD1.n143 B 0.020049f
C372 VDD1.n144 B 0.010774f
C373 VDD1.n145 B 0.011407f
C374 VDD1.n146 B 0.025465f
C375 VDD1.n147 B 0.025465f
C376 VDD1.n148 B 0.011407f
C377 VDD1.n149 B 0.010774f
C378 VDD1.n150 B 0.020049f
C379 VDD1.n151 B 0.020049f
C380 VDD1.n152 B 0.010774f
C381 VDD1.n153 B 0.010774f
C382 VDD1.n154 B 0.011407f
C383 VDD1.n155 B 0.025465f
C384 VDD1.n156 B 0.025465f
C385 VDD1.n157 B 0.025465f
C386 VDD1.n158 B 0.01109f
C387 VDD1.n159 B 0.010774f
C388 VDD1.n160 B 0.020049f
C389 VDD1.n161 B 0.020049f
C390 VDD1.n162 B 0.010774f
C391 VDD1.n163 B 0.011407f
C392 VDD1.n164 B 0.025465f
C393 VDD1.n165 B 0.025465f
C394 VDD1.n166 B 0.011407f
C395 VDD1.n167 B 0.010774f
C396 VDD1.n168 B 0.020049f
C397 VDD1.n169 B 0.020049f
C398 VDD1.n170 B 0.010774f
C399 VDD1.n171 B 0.011407f
C400 VDD1.n172 B 0.025465f
C401 VDD1.n173 B 0.025465f
C402 VDD1.n174 B 0.011407f
C403 VDD1.n175 B 0.010774f
C404 VDD1.n176 B 0.020049f
C405 VDD1.n177 B 0.020049f
C406 VDD1.n178 B 0.010774f
C407 VDD1.n179 B 0.011407f
C408 VDD1.n180 B 0.025465f
C409 VDD1.n181 B 0.025465f
C410 VDD1.n182 B 0.011407f
C411 VDD1.n183 B 0.010774f
C412 VDD1.n184 B 0.020049f
C413 VDD1.n185 B 0.020049f
C414 VDD1.n186 B 0.010774f
C415 VDD1.n187 B 0.011407f
C416 VDD1.n188 B 0.025465f
C417 VDD1.n189 B 0.025465f
C418 VDD1.n190 B 0.011407f
C419 VDD1.n191 B 0.010774f
C420 VDD1.n192 B 0.020049f
C421 VDD1.n193 B 0.020049f
C422 VDD1.n194 B 0.010774f
C423 VDD1.n195 B 0.011407f
C424 VDD1.n196 B 0.025465f
C425 VDD1.n197 B 0.025465f
C426 VDD1.n198 B 0.011407f
C427 VDD1.n199 B 0.010774f
C428 VDD1.n200 B 0.020049f
C429 VDD1.n201 B 0.051273f
C430 VDD1.n202 B 0.010774f
C431 VDD1.n203 B 0.011407f
C432 VDD1.n204 B 0.051778f
C433 VDD1.n205 B 0.806885f
C434 VTAIL.n0 B 0.011065f
C435 VTAIL.n1 B 0.024947f
C436 VTAIL.n2 B 0.011175f
C437 VTAIL.n3 B 0.019642f
C438 VTAIL.n4 B 0.010554f
C439 VTAIL.n5 B 0.024947f
C440 VTAIL.n6 B 0.011175f
C441 VTAIL.n7 B 0.019642f
C442 VTAIL.n8 B 0.010554f
C443 VTAIL.n9 B 0.024947f
C444 VTAIL.n10 B 0.011175f
C445 VTAIL.n11 B 0.019642f
C446 VTAIL.n12 B 0.010554f
C447 VTAIL.n13 B 0.024947f
C448 VTAIL.n14 B 0.011175f
C449 VTAIL.n15 B 0.019642f
C450 VTAIL.n16 B 0.010554f
C451 VTAIL.n17 B 0.024947f
C452 VTAIL.n18 B 0.011175f
C453 VTAIL.n19 B 0.019642f
C454 VTAIL.n20 B 0.010554f
C455 VTAIL.n21 B 0.024947f
C456 VTAIL.n22 B 0.010865f
C457 VTAIL.n23 B 0.019642f
C458 VTAIL.n24 B 0.011175f
C459 VTAIL.n25 B 0.024947f
C460 VTAIL.n26 B 0.011175f
C461 VTAIL.n27 B 0.019642f
C462 VTAIL.n28 B 0.010554f
C463 VTAIL.n29 B 0.024947f
C464 VTAIL.n30 B 0.011175f
C465 VTAIL.n31 B 1.5832f
C466 VTAIL.n32 B 0.010554f
C467 VTAIL.t2 B 0.042851f
C468 VTAIL.n33 B 0.19274f
C469 VTAIL.n34 B 0.017636f
C470 VTAIL.n35 B 0.01871f
C471 VTAIL.n36 B 0.024947f
C472 VTAIL.n37 B 0.011175f
C473 VTAIL.n38 B 0.010554f
C474 VTAIL.n39 B 0.019642f
C475 VTAIL.n40 B 0.019642f
C476 VTAIL.n41 B 0.010554f
C477 VTAIL.n42 B 0.011175f
C478 VTAIL.n43 B 0.024947f
C479 VTAIL.n44 B 0.024947f
C480 VTAIL.n45 B 0.011175f
C481 VTAIL.n46 B 0.010554f
C482 VTAIL.n47 B 0.019642f
C483 VTAIL.n48 B 0.019642f
C484 VTAIL.n49 B 0.010554f
C485 VTAIL.n50 B 0.010554f
C486 VTAIL.n51 B 0.011175f
C487 VTAIL.n52 B 0.024947f
C488 VTAIL.n53 B 0.024947f
C489 VTAIL.n54 B 0.024947f
C490 VTAIL.n55 B 0.010865f
C491 VTAIL.n56 B 0.010554f
C492 VTAIL.n57 B 0.019642f
C493 VTAIL.n58 B 0.019642f
C494 VTAIL.n59 B 0.010554f
C495 VTAIL.n60 B 0.011175f
C496 VTAIL.n61 B 0.024947f
C497 VTAIL.n62 B 0.024947f
C498 VTAIL.n63 B 0.011175f
C499 VTAIL.n64 B 0.010554f
C500 VTAIL.n65 B 0.019642f
C501 VTAIL.n66 B 0.019642f
C502 VTAIL.n67 B 0.010554f
C503 VTAIL.n68 B 0.011175f
C504 VTAIL.n69 B 0.024947f
C505 VTAIL.n70 B 0.024947f
C506 VTAIL.n71 B 0.011175f
C507 VTAIL.n72 B 0.010554f
C508 VTAIL.n73 B 0.019642f
C509 VTAIL.n74 B 0.019642f
C510 VTAIL.n75 B 0.010554f
C511 VTAIL.n76 B 0.011175f
C512 VTAIL.n77 B 0.024947f
C513 VTAIL.n78 B 0.024947f
C514 VTAIL.n79 B 0.011175f
C515 VTAIL.n80 B 0.010554f
C516 VTAIL.n81 B 0.019642f
C517 VTAIL.n82 B 0.019642f
C518 VTAIL.n83 B 0.010554f
C519 VTAIL.n84 B 0.011175f
C520 VTAIL.n85 B 0.024947f
C521 VTAIL.n86 B 0.024947f
C522 VTAIL.n87 B 0.011175f
C523 VTAIL.n88 B 0.010554f
C524 VTAIL.n89 B 0.019642f
C525 VTAIL.n90 B 0.019642f
C526 VTAIL.n91 B 0.010554f
C527 VTAIL.n92 B 0.011175f
C528 VTAIL.n93 B 0.024947f
C529 VTAIL.n94 B 0.024947f
C530 VTAIL.n95 B 0.011175f
C531 VTAIL.n96 B 0.010554f
C532 VTAIL.n97 B 0.019642f
C533 VTAIL.n98 B 0.05023f
C534 VTAIL.n99 B 0.010554f
C535 VTAIL.n100 B 0.011175f
C536 VTAIL.n101 B 0.050725f
C537 VTAIL.n102 B 0.042558f
C538 VTAIL.n103 B 1.66692f
C539 VTAIL.n104 B 0.011065f
C540 VTAIL.n105 B 0.024947f
C541 VTAIL.n106 B 0.011175f
C542 VTAIL.n107 B 0.019642f
C543 VTAIL.n108 B 0.010554f
C544 VTAIL.n109 B 0.024947f
C545 VTAIL.n110 B 0.011175f
C546 VTAIL.n111 B 0.019642f
C547 VTAIL.n112 B 0.010554f
C548 VTAIL.n113 B 0.024947f
C549 VTAIL.n114 B 0.011175f
C550 VTAIL.n115 B 0.019642f
C551 VTAIL.n116 B 0.010554f
C552 VTAIL.n117 B 0.024947f
C553 VTAIL.n118 B 0.011175f
C554 VTAIL.n119 B 0.019642f
C555 VTAIL.n120 B 0.010554f
C556 VTAIL.n121 B 0.024947f
C557 VTAIL.n122 B 0.011175f
C558 VTAIL.n123 B 0.019642f
C559 VTAIL.n124 B 0.010554f
C560 VTAIL.n125 B 0.024947f
C561 VTAIL.n126 B 0.010865f
C562 VTAIL.n127 B 0.019642f
C563 VTAIL.n128 B 0.010865f
C564 VTAIL.n129 B 0.010554f
C565 VTAIL.n130 B 0.024947f
C566 VTAIL.n131 B 0.024947f
C567 VTAIL.n132 B 0.011175f
C568 VTAIL.n133 B 0.019642f
C569 VTAIL.n134 B 0.010554f
C570 VTAIL.n135 B 0.024947f
C571 VTAIL.n136 B 0.011175f
C572 VTAIL.n137 B 1.5832f
C573 VTAIL.n138 B 0.010554f
C574 VTAIL.t3 B 0.042851f
C575 VTAIL.n139 B 0.19274f
C576 VTAIL.n140 B 0.017636f
C577 VTAIL.n141 B 0.01871f
C578 VTAIL.n142 B 0.024947f
C579 VTAIL.n143 B 0.011175f
C580 VTAIL.n144 B 0.010554f
C581 VTAIL.n145 B 0.019642f
C582 VTAIL.n146 B 0.019642f
C583 VTAIL.n147 B 0.010554f
C584 VTAIL.n148 B 0.011175f
C585 VTAIL.n149 B 0.024947f
C586 VTAIL.n150 B 0.024947f
C587 VTAIL.n151 B 0.011175f
C588 VTAIL.n152 B 0.010554f
C589 VTAIL.n153 B 0.019642f
C590 VTAIL.n154 B 0.019642f
C591 VTAIL.n155 B 0.010554f
C592 VTAIL.n156 B 0.011175f
C593 VTAIL.n157 B 0.024947f
C594 VTAIL.n158 B 0.024947f
C595 VTAIL.n159 B 0.011175f
C596 VTAIL.n160 B 0.010554f
C597 VTAIL.n161 B 0.019642f
C598 VTAIL.n162 B 0.019642f
C599 VTAIL.n163 B 0.010554f
C600 VTAIL.n164 B 0.011175f
C601 VTAIL.n165 B 0.024947f
C602 VTAIL.n166 B 0.024947f
C603 VTAIL.n167 B 0.011175f
C604 VTAIL.n168 B 0.010554f
C605 VTAIL.n169 B 0.019642f
C606 VTAIL.n170 B 0.019642f
C607 VTAIL.n171 B 0.010554f
C608 VTAIL.n172 B 0.011175f
C609 VTAIL.n173 B 0.024947f
C610 VTAIL.n174 B 0.024947f
C611 VTAIL.n175 B 0.011175f
C612 VTAIL.n176 B 0.010554f
C613 VTAIL.n177 B 0.019642f
C614 VTAIL.n178 B 0.019642f
C615 VTAIL.n179 B 0.010554f
C616 VTAIL.n180 B 0.011175f
C617 VTAIL.n181 B 0.024947f
C618 VTAIL.n182 B 0.024947f
C619 VTAIL.n183 B 0.011175f
C620 VTAIL.n184 B 0.010554f
C621 VTAIL.n185 B 0.019642f
C622 VTAIL.n186 B 0.019642f
C623 VTAIL.n187 B 0.010554f
C624 VTAIL.n188 B 0.011175f
C625 VTAIL.n189 B 0.024947f
C626 VTAIL.n190 B 0.024947f
C627 VTAIL.n191 B 0.011175f
C628 VTAIL.n192 B 0.010554f
C629 VTAIL.n193 B 0.019642f
C630 VTAIL.n194 B 0.019642f
C631 VTAIL.n195 B 0.010554f
C632 VTAIL.n196 B 0.011175f
C633 VTAIL.n197 B 0.024947f
C634 VTAIL.n198 B 0.024947f
C635 VTAIL.n199 B 0.011175f
C636 VTAIL.n200 B 0.010554f
C637 VTAIL.n201 B 0.019642f
C638 VTAIL.n202 B 0.05023f
C639 VTAIL.n203 B 0.010554f
C640 VTAIL.n204 B 0.011175f
C641 VTAIL.n205 B 0.050725f
C642 VTAIL.n206 B 0.042558f
C643 VTAIL.n207 B 1.69911f
C644 VTAIL.n208 B 0.011065f
C645 VTAIL.n209 B 0.024947f
C646 VTAIL.n210 B 0.011175f
C647 VTAIL.n211 B 0.019642f
C648 VTAIL.n212 B 0.010554f
C649 VTAIL.n213 B 0.024947f
C650 VTAIL.n214 B 0.011175f
C651 VTAIL.n215 B 0.019642f
C652 VTAIL.n216 B 0.010554f
C653 VTAIL.n217 B 0.024947f
C654 VTAIL.n218 B 0.011175f
C655 VTAIL.n219 B 0.019642f
C656 VTAIL.n220 B 0.010554f
C657 VTAIL.n221 B 0.024947f
C658 VTAIL.n222 B 0.011175f
C659 VTAIL.n223 B 0.019642f
C660 VTAIL.n224 B 0.010554f
C661 VTAIL.n225 B 0.024947f
C662 VTAIL.n226 B 0.011175f
C663 VTAIL.n227 B 0.019642f
C664 VTAIL.n228 B 0.010554f
C665 VTAIL.n229 B 0.024947f
C666 VTAIL.n230 B 0.010865f
C667 VTAIL.n231 B 0.019642f
C668 VTAIL.n232 B 0.010865f
C669 VTAIL.n233 B 0.010554f
C670 VTAIL.n234 B 0.024947f
C671 VTAIL.n235 B 0.024947f
C672 VTAIL.n236 B 0.011175f
C673 VTAIL.n237 B 0.019642f
C674 VTAIL.n238 B 0.010554f
C675 VTAIL.n239 B 0.024947f
C676 VTAIL.n240 B 0.011175f
C677 VTAIL.n241 B 1.5832f
C678 VTAIL.n242 B 0.010554f
C679 VTAIL.t1 B 0.042851f
C680 VTAIL.n243 B 0.19274f
C681 VTAIL.n244 B 0.017636f
C682 VTAIL.n245 B 0.01871f
C683 VTAIL.n246 B 0.024947f
C684 VTAIL.n247 B 0.011175f
C685 VTAIL.n248 B 0.010554f
C686 VTAIL.n249 B 0.019642f
C687 VTAIL.n250 B 0.019642f
C688 VTAIL.n251 B 0.010554f
C689 VTAIL.n252 B 0.011175f
C690 VTAIL.n253 B 0.024947f
C691 VTAIL.n254 B 0.024947f
C692 VTAIL.n255 B 0.011175f
C693 VTAIL.n256 B 0.010554f
C694 VTAIL.n257 B 0.019642f
C695 VTAIL.n258 B 0.019642f
C696 VTAIL.n259 B 0.010554f
C697 VTAIL.n260 B 0.011175f
C698 VTAIL.n261 B 0.024947f
C699 VTAIL.n262 B 0.024947f
C700 VTAIL.n263 B 0.011175f
C701 VTAIL.n264 B 0.010554f
C702 VTAIL.n265 B 0.019642f
C703 VTAIL.n266 B 0.019642f
C704 VTAIL.n267 B 0.010554f
C705 VTAIL.n268 B 0.011175f
C706 VTAIL.n269 B 0.024947f
C707 VTAIL.n270 B 0.024947f
C708 VTAIL.n271 B 0.011175f
C709 VTAIL.n272 B 0.010554f
C710 VTAIL.n273 B 0.019642f
C711 VTAIL.n274 B 0.019642f
C712 VTAIL.n275 B 0.010554f
C713 VTAIL.n276 B 0.011175f
C714 VTAIL.n277 B 0.024947f
C715 VTAIL.n278 B 0.024947f
C716 VTAIL.n279 B 0.011175f
C717 VTAIL.n280 B 0.010554f
C718 VTAIL.n281 B 0.019642f
C719 VTAIL.n282 B 0.019642f
C720 VTAIL.n283 B 0.010554f
C721 VTAIL.n284 B 0.011175f
C722 VTAIL.n285 B 0.024947f
C723 VTAIL.n286 B 0.024947f
C724 VTAIL.n287 B 0.011175f
C725 VTAIL.n288 B 0.010554f
C726 VTAIL.n289 B 0.019642f
C727 VTAIL.n290 B 0.019642f
C728 VTAIL.n291 B 0.010554f
C729 VTAIL.n292 B 0.011175f
C730 VTAIL.n293 B 0.024947f
C731 VTAIL.n294 B 0.024947f
C732 VTAIL.n295 B 0.011175f
C733 VTAIL.n296 B 0.010554f
C734 VTAIL.n297 B 0.019642f
C735 VTAIL.n298 B 0.019642f
C736 VTAIL.n299 B 0.010554f
C737 VTAIL.n300 B 0.011175f
C738 VTAIL.n301 B 0.024947f
C739 VTAIL.n302 B 0.024947f
C740 VTAIL.n303 B 0.011175f
C741 VTAIL.n304 B 0.010554f
C742 VTAIL.n305 B 0.019642f
C743 VTAIL.n306 B 0.05023f
C744 VTAIL.n307 B 0.010554f
C745 VTAIL.n308 B 0.011175f
C746 VTAIL.n309 B 0.050725f
C747 VTAIL.n310 B 0.042558f
C748 VTAIL.n311 B 1.55562f
C749 VTAIL.n312 B 0.011065f
C750 VTAIL.n313 B 0.024947f
C751 VTAIL.n314 B 0.011175f
C752 VTAIL.n315 B 0.019642f
C753 VTAIL.n316 B 0.010554f
C754 VTAIL.n317 B 0.024947f
C755 VTAIL.n318 B 0.011175f
C756 VTAIL.n319 B 0.019642f
C757 VTAIL.n320 B 0.010554f
C758 VTAIL.n321 B 0.024947f
C759 VTAIL.n322 B 0.011175f
C760 VTAIL.n323 B 0.019642f
C761 VTAIL.n324 B 0.010554f
C762 VTAIL.n325 B 0.024947f
C763 VTAIL.n326 B 0.011175f
C764 VTAIL.n327 B 0.019642f
C765 VTAIL.n328 B 0.010554f
C766 VTAIL.n329 B 0.024947f
C767 VTAIL.n330 B 0.011175f
C768 VTAIL.n331 B 0.019642f
C769 VTAIL.n332 B 0.010554f
C770 VTAIL.n333 B 0.024947f
C771 VTAIL.n334 B 0.010865f
C772 VTAIL.n335 B 0.019642f
C773 VTAIL.n336 B 0.011175f
C774 VTAIL.n337 B 0.024947f
C775 VTAIL.n338 B 0.011175f
C776 VTAIL.n339 B 0.019642f
C777 VTAIL.n340 B 0.010554f
C778 VTAIL.n341 B 0.024947f
C779 VTAIL.n342 B 0.011175f
C780 VTAIL.n343 B 1.5832f
C781 VTAIL.n344 B 0.010554f
C782 VTAIL.t0 B 0.042851f
C783 VTAIL.n345 B 0.19274f
C784 VTAIL.n346 B 0.017636f
C785 VTAIL.n347 B 0.01871f
C786 VTAIL.n348 B 0.024947f
C787 VTAIL.n349 B 0.011175f
C788 VTAIL.n350 B 0.010554f
C789 VTAIL.n351 B 0.019642f
C790 VTAIL.n352 B 0.019642f
C791 VTAIL.n353 B 0.010554f
C792 VTAIL.n354 B 0.011175f
C793 VTAIL.n355 B 0.024947f
C794 VTAIL.n356 B 0.024947f
C795 VTAIL.n357 B 0.011175f
C796 VTAIL.n358 B 0.010554f
C797 VTAIL.n359 B 0.019642f
C798 VTAIL.n360 B 0.019642f
C799 VTAIL.n361 B 0.010554f
C800 VTAIL.n362 B 0.010554f
C801 VTAIL.n363 B 0.011175f
C802 VTAIL.n364 B 0.024947f
C803 VTAIL.n365 B 0.024947f
C804 VTAIL.n366 B 0.024947f
C805 VTAIL.n367 B 0.010865f
C806 VTAIL.n368 B 0.010554f
C807 VTAIL.n369 B 0.019642f
C808 VTAIL.n370 B 0.019642f
C809 VTAIL.n371 B 0.010554f
C810 VTAIL.n372 B 0.011175f
C811 VTAIL.n373 B 0.024947f
C812 VTAIL.n374 B 0.024947f
C813 VTAIL.n375 B 0.011175f
C814 VTAIL.n376 B 0.010554f
C815 VTAIL.n377 B 0.019642f
C816 VTAIL.n378 B 0.019642f
C817 VTAIL.n379 B 0.010554f
C818 VTAIL.n380 B 0.011175f
C819 VTAIL.n381 B 0.024947f
C820 VTAIL.n382 B 0.024947f
C821 VTAIL.n383 B 0.011175f
C822 VTAIL.n384 B 0.010554f
C823 VTAIL.n385 B 0.019642f
C824 VTAIL.n386 B 0.019642f
C825 VTAIL.n387 B 0.010554f
C826 VTAIL.n388 B 0.011175f
C827 VTAIL.n389 B 0.024947f
C828 VTAIL.n390 B 0.024947f
C829 VTAIL.n391 B 0.011175f
C830 VTAIL.n392 B 0.010554f
C831 VTAIL.n393 B 0.019642f
C832 VTAIL.n394 B 0.019642f
C833 VTAIL.n395 B 0.010554f
C834 VTAIL.n396 B 0.011175f
C835 VTAIL.n397 B 0.024947f
C836 VTAIL.n398 B 0.024947f
C837 VTAIL.n399 B 0.011175f
C838 VTAIL.n400 B 0.010554f
C839 VTAIL.n401 B 0.019642f
C840 VTAIL.n402 B 0.019642f
C841 VTAIL.n403 B 0.010554f
C842 VTAIL.n404 B 0.011175f
C843 VTAIL.n405 B 0.024947f
C844 VTAIL.n406 B 0.024947f
C845 VTAIL.n407 B 0.011175f
C846 VTAIL.n408 B 0.010554f
C847 VTAIL.n409 B 0.019642f
C848 VTAIL.n410 B 0.05023f
C849 VTAIL.n411 B 0.010554f
C850 VTAIL.n412 B 0.011175f
C851 VTAIL.n413 B 0.050725f
C852 VTAIL.n414 B 0.042558f
C853 VTAIL.n415 B 1.48633f
C854 VP.t0 B 4.64741f
C855 VP.t1 B 4.14115f
C856 VP.n0 B 5.54306f
.ends

