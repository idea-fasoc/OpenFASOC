* NGSPICE file created from diff_pair_sample_1337.ext - technology: sky130A

.subckt diff_pair_sample_1337 VTAIL VN VP B VDD2 VDD1
X0 B.t11 B.t9 B.t10 w_n1924_n1682# sky130_fd_pr__pfet_01v8 ad=1.3923 pd=7.92 as=0 ps=0 w=3.57 l=1.26
X1 VTAIL.t7 VN.t0 VDD2.t2 w_n1924_n1682# sky130_fd_pr__pfet_01v8 ad=1.3923 pd=7.92 as=0.58905 ps=3.9 w=3.57 l=1.26
X2 VDD1.t3 VP.t0 VTAIL.t3 w_n1924_n1682# sky130_fd_pr__pfet_01v8 ad=0.58905 pd=3.9 as=1.3923 ps=7.92 w=3.57 l=1.26
X3 VDD2.t1 VN.t1 VTAIL.t6 w_n1924_n1682# sky130_fd_pr__pfet_01v8 ad=0.58905 pd=3.9 as=1.3923 ps=7.92 w=3.57 l=1.26
X4 B.t8 B.t6 B.t7 w_n1924_n1682# sky130_fd_pr__pfet_01v8 ad=1.3923 pd=7.92 as=0 ps=0 w=3.57 l=1.26
X5 VDD2.t0 VN.t2 VTAIL.t5 w_n1924_n1682# sky130_fd_pr__pfet_01v8 ad=0.58905 pd=3.9 as=1.3923 ps=7.92 w=3.57 l=1.26
X6 B.t5 B.t3 B.t4 w_n1924_n1682# sky130_fd_pr__pfet_01v8 ad=1.3923 pd=7.92 as=0 ps=0 w=3.57 l=1.26
X7 VTAIL.t4 VN.t3 VDD2.t3 w_n1924_n1682# sky130_fd_pr__pfet_01v8 ad=1.3923 pd=7.92 as=0.58905 ps=3.9 w=3.57 l=1.26
X8 VTAIL.t2 VP.t1 VDD1.t2 w_n1924_n1682# sky130_fd_pr__pfet_01v8 ad=1.3923 pd=7.92 as=0.58905 ps=3.9 w=3.57 l=1.26
X9 VTAIL.t0 VP.t2 VDD1.t1 w_n1924_n1682# sky130_fd_pr__pfet_01v8 ad=1.3923 pd=7.92 as=0.58905 ps=3.9 w=3.57 l=1.26
X10 B.t2 B.t0 B.t1 w_n1924_n1682# sky130_fd_pr__pfet_01v8 ad=1.3923 pd=7.92 as=0 ps=0 w=3.57 l=1.26
X11 VDD1.t0 VP.t3 VTAIL.t1 w_n1924_n1682# sky130_fd_pr__pfet_01v8 ad=0.58905 pd=3.9 as=1.3923 ps=7.92 w=3.57 l=1.26
R0 B.n264 B.n263 585
R1 B.n265 B.n38 585
R2 B.n267 B.n266 585
R3 B.n268 B.n37 585
R4 B.n270 B.n269 585
R5 B.n271 B.n36 585
R6 B.n273 B.n272 585
R7 B.n274 B.n35 585
R8 B.n276 B.n275 585
R9 B.n277 B.n34 585
R10 B.n279 B.n278 585
R11 B.n280 B.n33 585
R12 B.n282 B.n281 585
R13 B.n283 B.n32 585
R14 B.n285 B.n284 585
R15 B.n286 B.n31 585
R16 B.n288 B.n287 585
R17 B.n290 B.n289 585
R18 B.n291 B.n27 585
R19 B.n293 B.n292 585
R20 B.n294 B.n26 585
R21 B.n296 B.n295 585
R22 B.n297 B.n25 585
R23 B.n299 B.n298 585
R24 B.n300 B.n24 585
R25 B.n302 B.n301 585
R26 B.n304 B.n21 585
R27 B.n306 B.n305 585
R28 B.n307 B.n20 585
R29 B.n309 B.n308 585
R30 B.n310 B.n19 585
R31 B.n312 B.n311 585
R32 B.n313 B.n18 585
R33 B.n315 B.n314 585
R34 B.n316 B.n17 585
R35 B.n318 B.n317 585
R36 B.n319 B.n16 585
R37 B.n321 B.n320 585
R38 B.n322 B.n15 585
R39 B.n324 B.n323 585
R40 B.n325 B.n14 585
R41 B.n327 B.n326 585
R42 B.n328 B.n13 585
R43 B.n262 B.n39 585
R44 B.n261 B.n260 585
R45 B.n259 B.n40 585
R46 B.n258 B.n257 585
R47 B.n256 B.n41 585
R48 B.n255 B.n254 585
R49 B.n253 B.n42 585
R50 B.n252 B.n251 585
R51 B.n250 B.n43 585
R52 B.n249 B.n248 585
R53 B.n247 B.n44 585
R54 B.n246 B.n245 585
R55 B.n244 B.n45 585
R56 B.n243 B.n242 585
R57 B.n241 B.n46 585
R58 B.n240 B.n239 585
R59 B.n238 B.n47 585
R60 B.n237 B.n236 585
R61 B.n235 B.n48 585
R62 B.n234 B.n233 585
R63 B.n232 B.n49 585
R64 B.n231 B.n230 585
R65 B.n229 B.n50 585
R66 B.n228 B.n227 585
R67 B.n226 B.n51 585
R68 B.n225 B.n224 585
R69 B.n223 B.n52 585
R70 B.n222 B.n221 585
R71 B.n220 B.n53 585
R72 B.n219 B.n218 585
R73 B.n217 B.n54 585
R74 B.n216 B.n215 585
R75 B.n214 B.n55 585
R76 B.n213 B.n212 585
R77 B.n211 B.n56 585
R78 B.n210 B.n209 585
R79 B.n208 B.n57 585
R80 B.n207 B.n206 585
R81 B.n205 B.n58 585
R82 B.n204 B.n203 585
R83 B.n202 B.n59 585
R84 B.n201 B.n200 585
R85 B.n199 B.n60 585
R86 B.n198 B.n197 585
R87 B.n196 B.n61 585
R88 B.n130 B.n87 585
R89 B.n132 B.n131 585
R90 B.n133 B.n86 585
R91 B.n135 B.n134 585
R92 B.n136 B.n85 585
R93 B.n138 B.n137 585
R94 B.n139 B.n84 585
R95 B.n141 B.n140 585
R96 B.n142 B.n83 585
R97 B.n144 B.n143 585
R98 B.n145 B.n82 585
R99 B.n147 B.n146 585
R100 B.n148 B.n81 585
R101 B.n150 B.n149 585
R102 B.n151 B.n80 585
R103 B.n153 B.n152 585
R104 B.n154 B.n77 585
R105 B.n157 B.n156 585
R106 B.n158 B.n76 585
R107 B.n160 B.n159 585
R108 B.n161 B.n75 585
R109 B.n163 B.n162 585
R110 B.n164 B.n74 585
R111 B.n166 B.n165 585
R112 B.n167 B.n73 585
R113 B.n169 B.n168 585
R114 B.n171 B.n170 585
R115 B.n172 B.n69 585
R116 B.n174 B.n173 585
R117 B.n175 B.n68 585
R118 B.n177 B.n176 585
R119 B.n178 B.n67 585
R120 B.n180 B.n179 585
R121 B.n181 B.n66 585
R122 B.n183 B.n182 585
R123 B.n184 B.n65 585
R124 B.n186 B.n185 585
R125 B.n187 B.n64 585
R126 B.n189 B.n188 585
R127 B.n190 B.n63 585
R128 B.n192 B.n191 585
R129 B.n193 B.n62 585
R130 B.n195 B.n194 585
R131 B.n129 B.n128 585
R132 B.n127 B.n88 585
R133 B.n126 B.n125 585
R134 B.n124 B.n89 585
R135 B.n123 B.n122 585
R136 B.n121 B.n90 585
R137 B.n120 B.n119 585
R138 B.n118 B.n91 585
R139 B.n117 B.n116 585
R140 B.n115 B.n92 585
R141 B.n114 B.n113 585
R142 B.n112 B.n93 585
R143 B.n111 B.n110 585
R144 B.n109 B.n94 585
R145 B.n108 B.n107 585
R146 B.n106 B.n95 585
R147 B.n105 B.n104 585
R148 B.n103 B.n96 585
R149 B.n102 B.n101 585
R150 B.n100 B.n97 585
R151 B.n99 B.n98 585
R152 B.n2 B.n0 585
R153 B.n361 B.n1 585
R154 B.n360 B.n359 585
R155 B.n358 B.n3 585
R156 B.n357 B.n356 585
R157 B.n355 B.n4 585
R158 B.n354 B.n353 585
R159 B.n352 B.n5 585
R160 B.n351 B.n350 585
R161 B.n349 B.n6 585
R162 B.n348 B.n347 585
R163 B.n346 B.n7 585
R164 B.n345 B.n344 585
R165 B.n343 B.n8 585
R166 B.n342 B.n341 585
R167 B.n340 B.n9 585
R168 B.n339 B.n338 585
R169 B.n337 B.n10 585
R170 B.n336 B.n335 585
R171 B.n334 B.n11 585
R172 B.n333 B.n332 585
R173 B.n331 B.n12 585
R174 B.n330 B.n329 585
R175 B.n363 B.n362 585
R176 B.n128 B.n87 540.549
R177 B.n330 B.n13 540.549
R178 B.n194 B.n61 540.549
R179 B.n264 B.n39 540.549
R180 B.n70 B.t0 272.702
R181 B.n78 B.t3 272.702
R182 B.n22 B.t9 272.702
R183 B.n28 B.t6 272.702
R184 B.n128 B.n127 163.367
R185 B.n127 B.n126 163.367
R186 B.n126 B.n89 163.367
R187 B.n122 B.n89 163.367
R188 B.n122 B.n121 163.367
R189 B.n121 B.n120 163.367
R190 B.n120 B.n91 163.367
R191 B.n116 B.n91 163.367
R192 B.n116 B.n115 163.367
R193 B.n115 B.n114 163.367
R194 B.n114 B.n93 163.367
R195 B.n110 B.n93 163.367
R196 B.n110 B.n109 163.367
R197 B.n109 B.n108 163.367
R198 B.n108 B.n95 163.367
R199 B.n104 B.n95 163.367
R200 B.n104 B.n103 163.367
R201 B.n103 B.n102 163.367
R202 B.n102 B.n97 163.367
R203 B.n98 B.n97 163.367
R204 B.n98 B.n2 163.367
R205 B.n362 B.n2 163.367
R206 B.n362 B.n361 163.367
R207 B.n361 B.n360 163.367
R208 B.n360 B.n3 163.367
R209 B.n356 B.n3 163.367
R210 B.n356 B.n355 163.367
R211 B.n355 B.n354 163.367
R212 B.n354 B.n5 163.367
R213 B.n350 B.n5 163.367
R214 B.n350 B.n349 163.367
R215 B.n349 B.n348 163.367
R216 B.n348 B.n7 163.367
R217 B.n344 B.n7 163.367
R218 B.n344 B.n343 163.367
R219 B.n343 B.n342 163.367
R220 B.n342 B.n9 163.367
R221 B.n338 B.n9 163.367
R222 B.n338 B.n337 163.367
R223 B.n337 B.n336 163.367
R224 B.n336 B.n11 163.367
R225 B.n332 B.n11 163.367
R226 B.n332 B.n331 163.367
R227 B.n331 B.n330 163.367
R228 B.n132 B.n87 163.367
R229 B.n133 B.n132 163.367
R230 B.n134 B.n133 163.367
R231 B.n134 B.n85 163.367
R232 B.n138 B.n85 163.367
R233 B.n139 B.n138 163.367
R234 B.n140 B.n139 163.367
R235 B.n140 B.n83 163.367
R236 B.n144 B.n83 163.367
R237 B.n145 B.n144 163.367
R238 B.n146 B.n145 163.367
R239 B.n146 B.n81 163.367
R240 B.n150 B.n81 163.367
R241 B.n151 B.n150 163.367
R242 B.n152 B.n151 163.367
R243 B.n152 B.n77 163.367
R244 B.n157 B.n77 163.367
R245 B.n158 B.n157 163.367
R246 B.n159 B.n158 163.367
R247 B.n159 B.n75 163.367
R248 B.n163 B.n75 163.367
R249 B.n164 B.n163 163.367
R250 B.n165 B.n164 163.367
R251 B.n165 B.n73 163.367
R252 B.n169 B.n73 163.367
R253 B.n170 B.n169 163.367
R254 B.n170 B.n69 163.367
R255 B.n174 B.n69 163.367
R256 B.n175 B.n174 163.367
R257 B.n176 B.n175 163.367
R258 B.n176 B.n67 163.367
R259 B.n180 B.n67 163.367
R260 B.n181 B.n180 163.367
R261 B.n182 B.n181 163.367
R262 B.n182 B.n65 163.367
R263 B.n186 B.n65 163.367
R264 B.n187 B.n186 163.367
R265 B.n188 B.n187 163.367
R266 B.n188 B.n63 163.367
R267 B.n192 B.n63 163.367
R268 B.n193 B.n192 163.367
R269 B.n194 B.n193 163.367
R270 B.n198 B.n61 163.367
R271 B.n199 B.n198 163.367
R272 B.n200 B.n199 163.367
R273 B.n200 B.n59 163.367
R274 B.n204 B.n59 163.367
R275 B.n205 B.n204 163.367
R276 B.n206 B.n205 163.367
R277 B.n206 B.n57 163.367
R278 B.n210 B.n57 163.367
R279 B.n211 B.n210 163.367
R280 B.n212 B.n211 163.367
R281 B.n212 B.n55 163.367
R282 B.n216 B.n55 163.367
R283 B.n217 B.n216 163.367
R284 B.n218 B.n217 163.367
R285 B.n218 B.n53 163.367
R286 B.n222 B.n53 163.367
R287 B.n223 B.n222 163.367
R288 B.n224 B.n223 163.367
R289 B.n224 B.n51 163.367
R290 B.n228 B.n51 163.367
R291 B.n229 B.n228 163.367
R292 B.n230 B.n229 163.367
R293 B.n230 B.n49 163.367
R294 B.n234 B.n49 163.367
R295 B.n235 B.n234 163.367
R296 B.n236 B.n235 163.367
R297 B.n236 B.n47 163.367
R298 B.n240 B.n47 163.367
R299 B.n241 B.n240 163.367
R300 B.n242 B.n241 163.367
R301 B.n242 B.n45 163.367
R302 B.n246 B.n45 163.367
R303 B.n247 B.n246 163.367
R304 B.n248 B.n247 163.367
R305 B.n248 B.n43 163.367
R306 B.n252 B.n43 163.367
R307 B.n253 B.n252 163.367
R308 B.n254 B.n253 163.367
R309 B.n254 B.n41 163.367
R310 B.n258 B.n41 163.367
R311 B.n259 B.n258 163.367
R312 B.n260 B.n259 163.367
R313 B.n260 B.n39 163.367
R314 B.n326 B.n13 163.367
R315 B.n326 B.n325 163.367
R316 B.n325 B.n324 163.367
R317 B.n324 B.n15 163.367
R318 B.n320 B.n15 163.367
R319 B.n320 B.n319 163.367
R320 B.n319 B.n318 163.367
R321 B.n318 B.n17 163.367
R322 B.n314 B.n17 163.367
R323 B.n314 B.n313 163.367
R324 B.n313 B.n312 163.367
R325 B.n312 B.n19 163.367
R326 B.n308 B.n19 163.367
R327 B.n308 B.n307 163.367
R328 B.n307 B.n306 163.367
R329 B.n306 B.n21 163.367
R330 B.n301 B.n21 163.367
R331 B.n301 B.n300 163.367
R332 B.n300 B.n299 163.367
R333 B.n299 B.n25 163.367
R334 B.n295 B.n25 163.367
R335 B.n295 B.n294 163.367
R336 B.n294 B.n293 163.367
R337 B.n293 B.n27 163.367
R338 B.n289 B.n27 163.367
R339 B.n289 B.n288 163.367
R340 B.n288 B.n31 163.367
R341 B.n284 B.n31 163.367
R342 B.n284 B.n283 163.367
R343 B.n283 B.n282 163.367
R344 B.n282 B.n33 163.367
R345 B.n278 B.n33 163.367
R346 B.n278 B.n277 163.367
R347 B.n277 B.n276 163.367
R348 B.n276 B.n35 163.367
R349 B.n272 B.n35 163.367
R350 B.n272 B.n271 163.367
R351 B.n271 B.n270 163.367
R352 B.n270 B.n37 163.367
R353 B.n266 B.n37 163.367
R354 B.n266 B.n265 163.367
R355 B.n265 B.n264 163.367
R356 B.n70 B.t2 160.308
R357 B.n28 B.t7 160.308
R358 B.n78 B.t5 160.304
R359 B.n22 B.t10 160.304
R360 B.n71 B.t1 129.47
R361 B.n29 B.t8 129.47
R362 B.n79 B.t4 129.468
R363 B.n23 B.t11 129.468
R364 B.n72 B.n71 59.5399
R365 B.n155 B.n79 59.5399
R366 B.n303 B.n23 59.5399
R367 B.n30 B.n29 59.5399
R368 B.n329 B.n328 35.1225
R369 B.n263 B.n262 35.1225
R370 B.n196 B.n195 35.1225
R371 B.n130 B.n129 35.1225
R372 B.n71 B.n70 30.8369
R373 B.n79 B.n78 30.8369
R374 B.n23 B.n22 30.8369
R375 B.n29 B.n28 30.8369
R376 B B.n363 18.0485
R377 B.n328 B.n327 10.6151
R378 B.n327 B.n14 10.6151
R379 B.n323 B.n14 10.6151
R380 B.n323 B.n322 10.6151
R381 B.n322 B.n321 10.6151
R382 B.n321 B.n16 10.6151
R383 B.n317 B.n16 10.6151
R384 B.n317 B.n316 10.6151
R385 B.n316 B.n315 10.6151
R386 B.n315 B.n18 10.6151
R387 B.n311 B.n18 10.6151
R388 B.n311 B.n310 10.6151
R389 B.n310 B.n309 10.6151
R390 B.n309 B.n20 10.6151
R391 B.n305 B.n20 10.6151
R392 B.n305 B.n304 10.6151
R393 B.n302 B.n24 10.6151
R394 B.n298 B.n24 10.6151
R395 B.n298 B.n297 10.6151
R396 B.n297 B.n296 10.6151
R397 B.n296 B.n26 10.6151
R398 B.n292 B.n26 10.6151
R399 B.n292 B.n291 10.6151
R400 B.n291 B.n290 10.6151
R401 B.n287 B.n286 10.6151
R402 B.n286 B.n285 10.6151
R403 B.n285 B.n32 10.6151
R404 B.n281 B.n32 10.6151
R405 B.n281 B.n280 10.6151
R406 B.n280 B.n279 10.6151
R407 B.n279 B.n34 10.6151
R408 B.n275 B.n34 10.6151
R409 B.n275 B.n274 10.6151
R410 B.n274 B.n273 10.6151
R411 B.n273 B.n36 10.6151
R412 B.n269 B.n36 10.6151
R413 B.n269 B.n268 10.6151
R414 B.n268 B.n267 10.6151
R415 B.n267 B.n38 10.6151
R416 B.n263 B.n38 10.6151
R417 B.n197 B.n196 10.6151
R418 B.n197 B.n60 10.6151
R419 B.n201 B.n60 10.6151
R420 B.n202 B.n201 10.6151
R421 B.n203 B.n202 10.6151
R422 B.n203 B.n58 10.6151
R423 B.n207 B.n58 10.6151
R424 B.n208 B.n207 10.6151
R425 B.n209 B.n208 10.6151
R426 B.n209 B.n56 10.6151
R427 B.n213 B.n56 10.6151
R428 B.n214 B.n213 10.6151
R429 B.n215 B.n214 10.6151
R430 B.n215 B.n54 10.6151
R431 B.n219 B.n54 10.6151
R432 B.n220 B.n219 10.6151
R433 B.n221 B.n220 10.6151
R434 B.n221 B.n52 10.6151
R435 B.n225 B.n52 10.6151
R436 B.n226 B.n225 10.6151
R437 B.n227 B.n226 10.6151
R438 B.n227 B.n50 10.6151
R439 B.n231 B.n50 10.6151
R440 B.n232 B.n231 10.6151
R441 B.n233 B.n232 10.6151
R442 B.n233 B.n48 10.6151
R443 B.n237 B.n48 10.6151
R444 B.n238 B.n237 10.6151
R445 B.n239 B.n238 10.6151
R446 B.n239 B.n46 10.6151
R447 B.n243 B.n46 10.6151
R448 B.n244 B.n243 10.6151
R449 B.n245 B.n244 10.6151
R450 B.n245 B.n44 10.6151
R451 B.n249 B.n44 10.6151
R452 B.n250 B.n249 10.6151
R453 B.n251 B.n250 10.6151
R454 B.n251 B.n42 10.6151
R455 B.n255 B.n42 10.6151
R456 B.n256 B.n255 10.6151
R457 B.n257 B.n256 10.6151
R458 B.n257 B.n40 10.6151
R459 B.n261 B.n40 10.6151
R460 B.n262 B.n261 10.6151
R461 B.n131 B.n130 10.6151
R462 B.n131 B.n86 10.6151
R463 B.n135 B.n86 10.6151
R464 B.n136 B.n135 10.6151
R465 B.n137 B.n136 10.6151
R466 B.n137 B.n84 10.6151
R467 B.n141 B.n84 10.6151
R468 B.n142 B.n141 10.6151
R469 B.n143 B.n142 10.6151
R470 B.n143 B.n82 10.6151
R471 B.n147 B.n82 10.6151
R472 B.n148 B.n147 10.6151
R473 B.n149 B.n148 10.6151
R474 B.n149 B.n80 10.6151
R475 B.n153 B.n80 10.6151
R476 B.n154 B.n153 10.6151
R477 B.n156 B.n76 10.6151
R478 B.n160 B.n76 10.6151
R479 B.n161 B.n160 10.6151
R480 B.n162 B.n161 10.6151
R481 B.n162 B.n74 10.6151
R482 B.n166 B.n74 10.6151
R483 B.n167 B.n166 10.6151
R484 B.n168 B.n167 10.6151
R485 B.n172 B.n171 10.6151
R486 B.n173 B.n172 10.6151
R487 B.n173 B.n68 10.6151
R488 B.n177 B.n68 10.6151
R489 B.n178 B.n177 10.6151
R490 B.n179 B.n178 10.6151
R491 B.n179 B.n66 10.6151
R492 B.n183 B.n66 10.6151
R493 B.n184 B.n183 10.6151
R494 B.n185 B.n184 10.6151
R495 B.n185 B.n64 10.6151
R496 B.n189 B.n64 10.6151
R497 B.n190 B.n189 10.6151
R498 B.n191 B.n190 10.6151
R499 B.n191 B.n62 10.6151
R500 B.n195 B.n62 10.6151
R501 B.n129 B.n88 10.6151
R502 B.n125 B.n88 10.6151
R503 B.n125 B.n124 10.6151
R504 B.n124 B.n123 10.6151
R505 B.n123 B.n90 10.6151
R506 B.n119 B.n90 10.6151
R507 B.n119 B.n118 10.6151
R508 B.n118 B.n117 10.6151
R509 B.n117 B.n92 10.6151
R510 B.n113 B.n92 10.6151
R511 B.n113 B.n112 10.6151
R512 B.n112 B.n111 10.6151
R513 B.n111 B.n94 10.6151
R514 B.n107 B.n94 10.6151
R515 B.n107 B.n106 10.6151
R516 B.n106 B.n105 10.6151
R517 B.n105 B.n96 10.6151
R518 B.n101 B.n96 10.6151
R519 B.n101 B.n100 10.6151
R520 B.n100 B.n99 10.6151
R521 B.n99 B.n0 10.6151
R522 B.n359 B.n1 10.6151
R523 B.n359 B.n358 10.6151
R524 B.n358 B.n357 10.6151
R525 B.n357 B.n4 10.6151
R526 B.n353 B.n4 10.6151
R527 B.n353 B.n352 10.6151
R528 B.n352 B.n351 10.6151
R529 B.n351 B.n6 10.6151
R530 B.n347 B.n6 10.6151
R531 B.n347 B.n346 10.6151
R532 B.n346 B.n345 10.6151
R533 B.n345 B.n8 10.6151
R534 B.n341 B.n8 10.6151
R535 B.n341 B.n340 10.6151
R536 B.n340 B.n339 10.6151
R537 B.n339 B.n10 10.6151
R538 B.n335 B.n10 10.6151
R539 B.n335 B.n334 10.6151
R540 B.n334 B.n333 10.6151
R541 B.n333 B.n12 10.6151
R542 B.n329 B.n12 10.6151
R543 B.n303 B.n302 6.5566
R544 B.n290 B.n30 6.5566
R545 B.n156 B.n155 6.5566
R546 B.n168 B.n72 6.5566
R547 B.n304 B.n303 4.05904
R548 B.n287 B.n30 4.05904
R549 B.n155 B.n154 4.05904
R550 B.n171 B.n72 4.05904
R551 B.n363 B.n0 2.81026
R552 B.n363 B.n1 2.81026
R553 VN.n0 VN.t0 105.194
R554 VN.n1 VN.t1 105.194
R555 VN.n0 VN.t2 104.969
R556 VN.n1 VN.t3 104.969
R557 VN VN.n1 54.2953
R558 VN VN.n0 18.2006
R559 VDD2.n2 VDD2.n0 152.558
R560 VDD2.n2 VDD2.n1 121.653
R561 VDD2.n1 VDD2.t3 9.10554
R562 VDD2.n1 VDD2.t1 9.10554
R563 VDD2.n0 VDD2.t2 9.10554
R564 VDD2.n0 VDD2.t0 9.10554
R565 VDD2 VDD2.n2 0.0586897
R566 VTAIL.n5 VTAIL.t2 114.079
R567 VTAIL.n4 VTAIL.t6 114.079
R568 VTAIL.n3 VTAIL.t4 114.079
R569 VTAIL.n7 VTAIL.t5 114.079
R570 VTAIL.n0 VTAIL.t7 114.079
R571 VTAIL.n1 VTAIL.t1 114.079
R572 VTAIL.n2 VTAIL.t0 114.079
R573 VTAIL.n6 VTAIL.t3 114.079
R574 VTAIL.n7 VTAIL.n6 16.8152
R575 VTAIL.n3 VTAIL.n2 16.8152
R576 VTAIL.n4 VTAIL.n3 1.37119
R577 VTAIL.n6 VTAIL.n5 1.37119
R578 VTAIL.n2 VTAIL.n1 1.37119
R579 VTAIL VTAIL.n0 0.744035
R580 VTAIL VTAIL.n7 0.627655
R581 VTAIL.n5 VTAIL.n4 0.470328
R582 VTAIL.n1 VTAIL.n0 0.470328
R583 VP.n4 VP.n3 171.332
R584 VP.n10 VP.n9 171.332
R585 VP.n8 VP.n0 161.3
R586 VP.n7 VP.n6 161.3
R587 VP.n5 VP.n1 161.3
R588 VP.n2 VP.t1 105.194
R589 VP.n2 VP.t0 104.969
R590 VP.n3 VP.t2 68.2838
R591 VP.n9 VP.t3 68.2838
R592 VP.n4 VP.n2 53.9146
R593 VP.n7 VP.n1 40.4934
R594 VP.n8 VP.n7 40.4934
R595 VP.n3 VP.n1 14.436
R596 VP.n9 VP.n8 14.436
R597 VP.n5 VP.n4 0.189894
R598 VP.n6 VP.n5 0.189894
R599 VP.n6 VP.n0 0.189894
R600 VP.n10 VP.n0 0.189894
R601 VP VP.n10 0.0516364
R602 VDD1 VDD1.n1 153.083
R603 VDD1 VDD1.n0 121.712
R604 VDD1.n0 VDD1.t2 9.10554
R605 VDD1.n0 VDD1.t3 9.10554
R606 VDD1.n1 VDD1.t1 9.10554
R607 VDD1.n1 VDD1.t0 9.10554
C0 VTAIL VDD1 2.95055f
C1 VDD2 VDD1 0.698925f
C2 VTAIL VN 1.53451f
C3 VDD2 VN 1.39728f
C4 w_n1924_n1682# VTAIL 1.97801f
C5 w_n1924_n1682# VDD2 0.980639f
C6 VP VDD1 1.55811f
C7 B VTAIL 1.72715f
C8 B VDD2 0.828198f
C9 VP VN 3.67068f
C10 w_n1924_n1682# VP 3.08758f
C11 VDD1 VN 0.152127f
C12 B VP 1.14946f
C13 w_n1924_n1682# VDD1 0.954685f
C14 w_n1924_n1682# VN 2.84509f
C15 B VDD1 0.79778f
C16 B VN 0.751165f
C17 B w_n1924_n1682# 5.2356f
C18 VDD2 VTAIL 2.99578f
C19 VP VTAIL 1.54862f
C20 VP VDD2 0.313802f
C21 VDD2 VSUBS 0.498657f
C22 VDD1 VSUBS 2.720535f
C23 VTAIL VSUBS 0.403463f
C24 VN VSUBS 3.95825f
C25 VP VSUBS 1.144767f
C26 B VSUBS 2.282791f
C27 w_n1924_n1682# VSUBS 40.842697f
C28 VDD1.t2 VSUBS 0.051192f
C29 VDD1.t3 VSUBS 0.051192f
C30 VDD1.n0 VSUBS 0.287638f
C31 VDD1.t1 VSUBS 0.051192f
C32 VDD1.t0 VSUBS 0.051192f
C33 VDD1.n1 VSUBS 0.459917f
C34 VP.n0 VSUBS 0.044251f
C35 VP.t3 VSUBS 0.505749f
C36 VP.n1 VSUBS 0.071253f
C37 VP.t1 VSUBS 0.63728f
C38 VP.t0 VSUBS 0.636449f
C39 VP.n2 VSUBS 1.57598f
C40 VP.t2 VSUBS 0.505749f
C41 VP.n3 VSUBS 0.308517f
C42 VP.n4 VSUBS 1.95184f
C43 VP.n5 VSUBS 0.044251f
C44 VP.n6 VSUBS 0.044251f
C45 VP.n7 VSUBS 0.035773f
C46 VP.n8 VSUBS 0.071253f
C47 VP.n9 VSUBS 0.308517f
C48 VP.n10 VSUBS 0.039384f
C49 VTAIL.t7 VSUBS 0.272501f
C50 VTAIL.n0 VSUBS 0.269371f
C51 VTAIL.t1 VSUBS 0.272501f
C52 VTAIL.n1 VSUBS 0.297001f
C53 VTAIL.t0 VSUBS 0.272501f
C54 VTAIL.n2 VSUBS 0.657997f
C55 VTAIL.t4 VSUBS 0.272502f
C56 VTAIL.n3 VSUBS 0.657996f
C57 VTAIL.t6 VSUBS 0.272502f
C58 VTAIL.n4 VSUBS 0.296999f
C59 VTAIL.t2 VSUBS 0.272502f
C60 VTAIL.n5 VSUBS 0.296999f
C61 VTAIL.t3 VSUBS 0.272501f
C62 VTAIL.n6 VSUBS 0.657998f
C63 VTAIL.t5 VSUBS 0.272501f
C64 VTAIL.n7 VSUBS 0.625241f
C65 VDD2.t2 VSUBS 0.052361f
C66 VDD2.t0 VSUBS 0.052361f
C67 VDD2.n0 VSUBS 0.460367f
C68 VDD2.t3 VSUBS 0.052361f
C69 VDD2.t1 VSUBS 0.052361f
C70 VDD2.n1 VSUBS 0.294046f
C71 VDD2.n2 VSUBS 1.95017f
C72 VN.t0 VSUBS 0.603643f
C73 VN.t2 VSUBS 0.602855f
C74 VN.n0 VSUBS 0.507717f
C75 VN.t1 VSUBS 0.603643f
C76 VN.t3 VSUBS 0.602855f
C77 VN.n1 VSUBS 1.51482f
C78 B.n0 VSUBS 0.004747f
C79 B.n1 VSUBS 0.004747f
C80 B.n2 VSUBS 0.007507f
C81 B.n3 VSUBS 0.007507f
C82 B.n4 VSUBS 0.007507f
C83 B.n5 VSUBS 0.007507f
C84 B.n6 VSUBS 0.007507f
C85 B.n7 VSUBS 0.007507f
C86 B.n8 VSUBS 0.007507f
C87 B.n9 VSUBS 0.007507f
C88 B.n10 VSUBS 0.007507f
C89 B.n11 VSUBS 0.007507f
C90 B.n12 VSUBS 0.007507f
C91 B.n13 VSUBS 0.018849f
C92 B.n14 VSUBS 0.007507f
C93 B.n15 VSUBS 0.007507f
C94 B.n16 VSUBS 0.007507f
C95 B.n17 VSUBS 0.007507f
C96 B.n18 VSUBS 0.007507f
C97 B.n19 VSUBS 0.007507f
C98 B.n20 VSUBS 0.007507f
C99 B.n21 VSUBS 0.007507f
C100 B.t11 VSUBS 0.097176f
C101 B.t10 VSUBS 0.107888f
C102 B.t9 VSUBS 0.225913f
C103 B.n22 VSUBS 0.081292f
C104 B.n23 VSUBS 0.066392f
C105 B.n24 VSUBS 0.007507f
C106 B.n25 VSUBS 0.007507f
C107 B.n26 VSUBS 0.007507f
C108 B.n27 VSUBS 0.007507f
C109 B.t8 VSUBS 0.097176f
C110 B.t7 VSUBS 0.107888f
C111 B.t6 VSUBS 0.225913f
C112 B.n28 VSUBS 0.081292f
C113 B.n29 VSUBS 0.066392f
C114 B.n30 VSUBS 0.017393f
C115 B.n31 VSUBS 0.007507f
C116 B.n32 VSUBS 0.007507f
C117 B.n33 VSUBS 0.007507f
C118 B.n34 VSUBS 0.007507f
C119 B.n35 VSUBS 0.007507f
C120 B.n36 VSUBS 0.007507f
C121 B.n37 VSUBS 0.007507f
C122 B.n38 VSUBS 0.007507f
C123 B.n39 VSUBS 0.018024f
C124 B.n40 VSUBS 0.007507f
C125 B.n41 VSUBS 0.007507f
C126 B.n42 VSUBS 0.007507f
C127 B.n43 VSUBS 0.007507f
C128 B.n44 VSUBS 0.007507f
C129 B.n45 VSUBS 0.007507f
C130 B.n46 VSUBS 0.007507f
C131 B.n47 VSUBS 0.007507f
C132 B.n48 VSUBS 0.007507f
C133 B.n49 VSUBS 0.007507f
C134 B.n50 VSUBS 0.007507f
C135 B.n51 VSUBS 0.007507f
C136 B.n52 VSUBS 0.007507f
C137 B.n53 VSUBS 0.007507f
C138 B.n54 VSUBS 0.007507f
C139 B.n55 VSUBS 0.007507f
C140 B.n56 VSUBS 0.007507f
C141 B.n57 VSUBS 0.007507f
C142 B.n58 VSUBS 0.007507f
C143 B.n59 VSUBS 0.007507f
C144 B.n60 VSUBS 0.007507f
C145 B.n61 VSUBS 0.018024f
C146 B.n62 VSUBS 0.007507f
C147 B.n63 VSUBS 0.007507f
C148 B.n64 VSUBS 0.007507f
C149 B.n65 VSUBS 0.007507f
C150 B.n66 VSUBS 0.007507f
C151 B.n67 VSUBS 0.007507f
C152 B.n68 VSUBS 0.007507f
C153 B.n69 VSUBS 0.007507f
C154 B.t1 VSUBS 0.097176f
C155 B.t2 VSUBS 0.107888f
C156 B.t0 VSUBS 0.225913f
C157 B.n70 VSUBS 0.081292f
C158 B.n71 VSUBS 0.066392f
C159 B.n72 VSUBS 0.017393f
C160 B.n73 VSUBS 0.007507f
C161 B.n74 VSUBS 0.007507f
C162 B.n75 VSUBS 0.007507f
C163 B.n76 VSUBS 0.007507f
C164 B.n77 VSUBS 0.007507f
C165 B.t4 VSUBS 0.097176f
C166 B.t5 VSUBS 0.107888f
C167 B.t3 VSUBS 0.225913f
C168 B.n78 VSUBS 0.081292f
C169 B.n79 VSUBS 0.066392f
C170 B.n80 VSUBS 0.007507f
C171 B.n81 VSUBS 0.007507f
C172 B.n82 VSUBS 0.007507f
C173 B.n83 VSUBS 0.007507f
C174 B.n84 VSUBS 0.007507f
C175 B.n85 VSUBS 0.007507f
C176 B.n86 VSUBS 0.007507f
C177 B.n87 VSUBS 0.018849f
C178 B.n88 VSUBS 0.007507f
C179 B.n89 VSUBS 0.007507f
C180 B.n90 VSUBS 0.007507f
C181 B.n91 VSUBS 0.007507f
C182 B.n92 VSUBS 0.007507f
C183 B.n93 VSUBS 0.007507f
C184 B.n94 VSUBS 0.007507f
C185 B.n95 VSUBS 0.007507f
C186 B.n96 VSUBS 0.007507f
C187 B.n97 VSUBS 0.007507f
C188 B.n98 VSUBS 0.007507f
C189 B.n99 VSUBS 0.007507f
C190 B.n100 VSUBS 0.007507f
C191 B.n101 VSUBS 0.007507f
C192 B.n102 VSUBS 0.007507f
C193 B.n103 VSUBS 0.007507f
C194 B.n104 VSUBS 0.007507f
C195 B.n105 VSUBS 0.007507f
C196 B.n106 VSUBS 0.007507f
C197 B.n107 VSUBS 0.007507f
C198 B.n108 VSUBS 0.007507f
C199 B.n109 VSUBS 0.007507f
C200 B.n110 VSUBS 0.007507f
C201 B.n111 VSUBS 0.007507f
C202 B.n112 VSUBS 0.007507f
C203 B.n113 VSUBS 0.007507f
C204 B.n114 VSUBS 0.007507f
C205 B.n115 VSUBS 0.007507f
C206 B.n116 VSUBS 0.007507f
C207 B.n117 VSUBS 0.007507f
C208 B.n118 VSUBS 0.007507f
C209 B.n119 VSUBS 0.007507f
C210 B.n120 VSUBS 0.007507f
C211 B.n121 VSUBS 0.007507f
C212 B.n122 VSUBS 0.007507f
C213 B.n123 VSUBS 0.007507f
C214 B.n124 VSUBS 0.007507f
C215 B.n125 VSUBS 0.007507f
C216 B.n126 VSUBS 0.007507f
C217 B.n127 VSUBS 0.007507f
C218 B.n128 VSUBS 0.018024f
C219 B.n129 VSUBS 0.018024f
C220 B.n130 VSUBS 0.018849f
C221 B.n131 VSUBS 0.007507f
C222 B.n132 VSUBS 0.007507f
C223 B.n133 VSUBS 0.007507f
C224 B.n134 VSUBS 0.007507f
C225 B.n135 VSUBS 0.007507f
C226 B.n136 VSUBS 0.007507f
C227 B.n137 VSUBS 0.007507f
C228 B.n138 VSUBS 0.007507f
C229 B.n139 VSUBS 0.007507f
C230 B.n140 VSUBS 0.007507f
C231 B.n141 VSUBS 0.007507f
C232 B.n142 VSUBS 0.007507f
C233 B.n143 VSUBS 0.007507f
C234 B.n144 VSUBS 0.007507f
C235 B.n145 VSUBS 0.007507f
C236 B.n146 VSUBS 0.007507f
C237 B.n147 VSUBS 0.007507f
C238 B.n148 VSUBS 0.007507f
C239 B.n149 VSUBS 0.007507f
C240 B.n150 VSUBS 0.007507f
C241 B.n151 VSUBS 0.007507f
C242 B.n152 VSUBS 0.007507f
C243 B.n153 VSUBS 0.007507f
C244 B.n154 VSUBS 0.005189f
C245 B.n155 VSUBS 0.017393f
C246 B.n156 VSUBS 0.006072f
C247 B.n157 VSUBS 0.007507f
C248 B.n158 VSUBS 0.007507f
C249 B.n159 VSUBS 0.007507f
C250 B.n160 VSUBS 0.007507f
C251 B.n161 VSUBS 0.007507f
C252 B.n162 VSUBS 0.007507f
C253 B.n163 VSUBS 0.007507f
C254 B.n164 VSUBS 0.007507f
C255 B.n165 VSUBS 0.007507f
C256 B.n166 VSUBS 0.007507f
C257 B.n167 VSUBS 0.007507f
C258 B.n168 VSUBS 0.006072f
C259 B.n169 VSUBS 0.007507f
C260 B.n170 VSUBS 0.007507f
C261 B.n171 VSUBS 0.005189f
C262 B.n172 VSUBS 0.007507f
C263 B.n173 VSUBS 0.007507f
C264 B.n174 VSUBS 0.007507f
C265 B.n175 VSUBS 0.007507f
C266 B.n176 VSUBS 0.007507f
C267 B.n177 VSUBS 0.007507f
C268 B.n178 VSUBS 0.007507f
C269 B.n179 VSUBS 0.007507f
C270 B.n180 VSUBS 0.007507f
C271 B.n181 VSUBS 0.007507f
C272 B.n182 VSUBS 0.007507f
C273 B.n183 VSUBS 0.007507f
C274 B.n184 VSUBS 0.007507f
C275 B.n185 VSUBS 0.007507f
C276 B.n186 VSUBS 0.007507f
C277 B.n187 VSUBS 0.007507f
C278 B.n188 VSUBS 0.007507f
C279 B.n189 VSUBS 0.007507f
C280 B.n190 VSUBS 0.007507f
C281 B.n191 VSUBS 0.007507f
C282 B.n192 VSUBS 0.007507f
C283 B.n193 VSUBS 0.007507f
C284 B.n194 VSUBS 0.018849f
C285 B.n195 VSUBS 0.018849f
C286 B.n196 VSUBS 0.018024f
C287 B.n197 VSUBS 0.007507f
C288 B.n198 VSUBS 0.007507f
C289 B.n199 VSUBS 0.007507f
C290 B.n200 VSUBS 0.007507f
C291 B.n201 VSUBS 0.007507f
C292 B.n202 VSUBS 0.007507f
C293 B.n203 VSUBS 0.007507f
C294 B.n204 VSUBS 0.007507f
C295 B.n205 VSUBS 0.007507f
C296 B.n206 VSUBS 0.007507f
C297 B.n207 VSUBS 0.007507f
C298 B.n208 VSUBS 0.007507f
C299 B.n209 VSUBS 0.007507f
C300 B.n210 VSUBS 0.007507f
C301 B.n211 VSUBS 0.007507f
C302 B.n212 VSUBS 0.007507f
C303 B.n213 VSUBS 0.007507f
C304 B.n214 VSUBS 0.007507f
C305 B.n215 VSUBS 0.007507f
C306 B.n216 VSUBS 0.007507f
C307 B.n217 VSUBS 0.007507f
C308 B.n218 VSUBS 0.007507f
C309 B.n219 VSUBS 0.007507f
C310 B.n220 VSUBS 0.007507f
C311 B.n221 VSUBS 0.007507f
C312 B.n222 VSUBS 0.007507f
C313 B.n223 VSUBS 0.007507f
C314 B.n224 VSUBS 0.007507f
C315 B.n225 VSUBS 0.007507f
C316 B.n226 VSUBS 0.007507f
C317 B.n227 VSUBS 0.007507f
C318 B.n228 VSUBS 0.007507f
C319 B.n229 VSUBS 0.007507f
C320 B.n230 VSUBS 0.007507f
C321 B.n231 VSUBS 0.007507f
C322 B.n232 VSUBS 0.007507f
C323 B.n233 VSUBS 0.007507f
C324 B.n234 VSUBS 0.007507f
C325 B.n235 VSUBS 0.007507f
C326 B.n236 VSUBS 0.007507f
C327 B.n237 VSUBS 0.007507f
C328 B.n238 VSUBS 0.007507f
C329 B.n239 VSUBS 0.007507f
C330 B.n240 VSUBS 0.007507f
C331 B.n241 VSUBS 0.007507f
C332 B.n242 VSUBS 0.007507f
C333 B.n243 VSUBS 0.007507f
C334 B.n244 VSUBS 0.007507f
C335 B.n245 VSUBS 0.007507f
C336 B.n246 VSUBS 0.007507f
C337 B.n247 VSUBS 0.007507f
C338 B.n248 VSUBS 0.007507f
C339 B.n249 VSUBS 0.007507f
C340 B.n250 VSUBS 0.007507f
C341 B.n251 VSUBS 0.007507f
C342 B.n252 VSUBS 0.007507f
C343 B.n253 VSUBS 0.007507f
C344 B.n254 VSUBS 0.007507f
C345 B.n255 VSUBS 0.007507f
C346 B.n256 VSUBS 0.007507f
C347 B.n257 VSUBS 0.007507f
C348 B.n258 VSUBS 0.007507f
C349 B.n259 VSUBS 0.007507f
C350 B.n260 VSUBS 0.007507f
C351 B.n261 VSUBS 0.007507f
C352 B.n262 VSUBS 0.018849f
C353 B.n263 VSUBS 0.018024f
C354 B.n264 VSUBS 0.018849f
C355 B.n265 VSUBS 0.007507f
C356 B.n266 VSUBS 0.007507f
C357 B.n267 VSUBS 0.007507f
C358 B.n268 VSUBS 0.007507f
C359 B.n269 VSUBS 0.007507f
C360 B.n270 VSUBS 0.007507f
C361 B.n271 VSUBS 0.007507f
C362 B.n272 VSUBS 0.007507f
C363 B.n273 VSUBS 0.007507f
C364 B.n274 VSUBS 0.007507f
C365 B.n275 VSUBS 0.007507f
C366 B.n276 VSUBS 0.007507f
C367 B.n277 VSUBS 0.007507f
C368 B.n278 VSUBS 0.007507f
C369 B.n279 VSUBS 0.007507f
C370 B.n280 VSUBS 0.007507f
C371 B.n281 VSUBS 0.007507f
C372 B.n282 VSUBS 0.007507f
C373 B.n283 VSUBS 0.007507f
C374 B.n284 VSUBS 0.007507f
C375 B.n285 VSUBS 0.007507f
C376 B.n286 VSUBS 0.007507f
C377 B.n287 VSUBS 0.005189f
C378 B.n288 VSUBS 0.007507f
C379 B.n289 VSUBS 0.007507f
C380 B.n290 VSUBS 0.006072f
C381 B.n291 VSUBS 0.007507f
C382 B.n292 VSUBS 0.007507f
C383 B.n293 VSUBS 0.007507f
C384 B.n294 VSUBS 0.007507f
C385 B.n295 VSUBS 0.007507f
C386 B.n296 VSUBS 0.007507f
C387 B.n297 VSUBS 0.007507f
C388 B.n298 VSUBS 0.007507f
C389 B.n299 VSUBS 0.007507f
C390 B.n300 VSUBS 0.007507f
C391 B.n301 VSUBS 0.007507f
C392 B.n302 VSUBS 0.006072f
C393 B.n303 VSUBS 0.017393f
C394 B.n304 VSUBS 0.005189f
C395 B.n305 VSUBS 0.007507f
C396 B.n306 VSUBS 0.007507f
C397 B.n307 VSUBS 0.007507f
C398 B.n308 VSUBS 0.007507f
C399 B.n309 VSUBS 0.007507f
C400 B.n310 VSUBS 0.007507f
C401 B.n311 VSUBS 0.007507f
C402 B.n312 VSUBS 0.007507f
C403 B.n313 VSUBS 0.007507f
C404 B.n314 VSUBS 0.007507f
C405 B.n315 VSUBS 0.007507f
C406 B.n316 VSUBS 0.007507f
C407 B.n317 VSUBS 0.007507f
C408 B.n318 VSUBS 0.007507f
C409 B.n319 VSUBS 0.007507f
C410 B.n320 VSUBS 0.007507f
C411 B.n321 VSUBS 0.007507f
C412 B.n322 VSUBS 0.007507f
C413 B.n323 VSUBS 0.007507f
C414 B.n324 VSUBS 0.007507f
C415 B.n325 VSUBS 0.007507f
C416 B.n326 VSUBS 0.007507f
C417 B.n327 VSUBS 0.007507f
C418 B.n328 VSUBS 0.018849f
C419 B.n329 VSUBS 0.018024f
C420 B.n330 VSUBS 0.018024f
C421 B.n331 VSUBS 0.007507f
C422 B.n332 VSUBS 0.007507f
C423 B.n333 VSUBS 0.007507f
C424 B.n334 VSUBS 0.007507f
C425 B.n335 VSUBS 0.007507f
C426 B.n336 VSUBS 0.007507f
C427 B.n337 VSUBS 0.007507f
C428 B.n338 VSUBS 0.007507f
C429 B.n339 VSUBS 0.007507f
C430 B.n340 VSUBS 0.007507f
C431 B.n341 VSUBS 0.007507f
C432 B.n342 VSUBS 0.007507f
C433 B.n343 VSUBS 0.007507f
C434 B.n344 VSUBS 0.007507f
C435 B.n345 VSUBS 0.007507f
C436 B.n346 VSUBS 0.007507f
C437 B.n347 VSUBS 0.007507f
C438 B.n348 VSUBS 0.007507f
C439 B.n349 VSUBS 0.007507f
C440 B.n350 VSUBS 0.007507f
C441 B.n351 VSUBS 0.007507f
C442 B.n352 VSUBS 0.007507f
C443 B.n353 VSUBS 0.007507f
C444 B.n354 VSUBS 0.007507f
C445 B.n355 VSUBS 0.007507f
C446 B.n356 VSUBS 0.007507f
C447 B.n357 VSUBS 0.007507f
C448 B.n358 VSUBS 0.007507f
C449 B.n359 VSUBS 0.007507f
C450 B.n360 VSUBS 0.007507f
C451 B.n361 VSUBS 0.007507f
C452 B.n362 VSUBS 0.007507f
C453 B.n363 VSUBS 0.016998f
.ends

