* NGSPICE file created from diff_pair_sample_1215.ext - technology: sky130A

.subckt diff_pair_sample_1215 VTAIL VN VP B VDD2 VDD1
X0 B.t11 B.t9 B.t10 w_n1750_n1582# sky130_fd_pr__pfet_01v8 ad=1.1973 pd=6.92 as=0 ps=0 w=3.07 l=1.62
X1 B.t8 B.t6 B.t7 w_n1750_n1582# sky130_fd_pr__pfet_01v8 ad=1.1973 pd=6.92 as=0 ps=0 w=3.07 l=1.62
X2 B.t5 B.t3 B.t4 w_n1750_n1582# sky130_fd_pr__pfet_01v8 ad=1.1973 pd=6.92 as=0 ps=0 w=3.07 l=1.62
X3 VDD1.t1 VP.t0 VTAIL.t2 w_n1750_n1582# sky130_fd_pr__pfet_01v8 ad=1.1973 pd=6.92 as=1.1973 ps=6.92 w=3.07 l=1.62
X4 VDD2.t1 VN.t0 VTAIL.t1 w_n1750_n1582# sky130_fd_pr__pfet_01v8 ad=1.1973 pd=6.92 as=1.1973 ps=6.92 w=3.07 l=1.62
X5 B.t2 B.t0 B.t1 w_n1750_n1582# sky130_fd_pr__pfet_01v8 ad=1.1973 pd=6.92 as=0 ps=0 w=3.07 l=1.62
X6 VDD2.t0 VN.t1 VTAIL.t0 w_n1750_n1582# sky130_fd_pr__pfet_01v8 ad=1.1973 pd=6.92 as=1.1973 ps=6.92 w=3.07 l=1.62
X7 VDD1.t0 VP.t1 VTAIL.t3 w_n1750_n1582# sky130_fd_pr__pfet_01v8 ad=1.1973 pd=6.92 as=1.1973 ps=6.92 w=3.07 l=1.62
R0 B.n177 B.n56 585
R1 B.n176 B.n175 585
R2 B.n174 B.n57 585
R3 B.n173 B.n172 585
R4 B.n171 B.n58 585
R5 B.n170 B.n169 585
R6 B.n168 B.n59 585
R7 B.n167 B.n166 585
R8 B.n165 B.n60 585
R9 B.n164 B.n163 585
R10 B.n162 B.n61 585
R11 B.n161 B.n160 585
R12 B.n159 B.n62 585
R13 B.n158 B.n157 585
R14 B.n156 B.n63 585
R15 B.n154 B.n153 585
R16 B.n152 B.n66 585
R17 B.n151 B.n150 585
R18 B.n149 B.n67 585
R19 B.n148 B.n147 585
R20 B.n146 B.n68 585
R21 B.n145 B.n144 585
R22 B.n143 B.n69 585
R23 B.n142 B.n141 585
R24 B.n140 B.n70 585
R25 B.n139 B.n138 585
R26 B.n134 B.n71 585
R27 B.n133 B.n132 585
R28 B.n131 B.n72 585
R29 B.n130 B.n129 585
R30 B.n128 B.n73 585
R31 B.n127 B.n126 585
R32 B.n125 B.n74 585
R33 B.n124 B.n123 585
R34 B.n122 B.n75 585
R35 B.n121 B.n120 585
R36 B.n119 B.n76 585
R37 B.n118 B.n117 585
R38 B.n116 B.n77 585
R39 B.n115 B.n114 585
R40 B.n179 B.n178 585
R41 B.n180 B.n55 585
R42 B.n182 B.n181 585
R43 B.n183 B.n54 585
R44 B.n185 B.n184 585
R45 B.n186 B.n53 585
R46 B.n188 B.n187 585
R47 B.n189 B.n52 585
R48 B.n191 B.n190 585
R49 B.n192 B.n51 585
R50 B.n194 B.n193 585
R51 B.n195 B.n50 585
R52 B.n197 B.n196 585
R53 B.n198 B.n49 585
R54 B.n200 B.n199 585
R55 B.n201 B.n48 585
R56 B.n203 B.n202 585
R57 B.n204 B.n47 585
R58 B.n206 B.n205 585
R59 B.n207 B.n46 585
R60 B.n209 B.n208 585
R61 B.n210 B.n45 585
R62 B.n212 B.n211 585
R63 B.n213 B.n44 585
R64 B.n215 B.n214 585
R65 B.n216 B.n43 585
R66 B.n218 B.n217 585
R67 B.n219 B.n42 585
R68 B.n221 B.n220 585
R69 B.n222 B.n41 585
R70 B.n224 B.n223 585
R71 B.n225 B.n40 585
R72 B.n227 B.n226 585
R73 B.n228 B.n39 585
R74 B.n230 B.n229 585
R75 B.n231 B.n38 585
R76 B.n233 B.n232 585
R77 B.n234 B.n37 585
R78 B.n236 B.n235 585
R79 B.n237 B.n36 585
R80 B.n299 B.n298 585
R81 B.n297 B.n12 585
R82 B.n296 B.n295 585
R83 B.n294 B.n13 585
R84 B.n293 B.n292 585
R85 B.n291 B.n14 585
R86 B.n290 B.n289 585
R87 B.n288 B.n15 585
R88 B.n287 B.n286 585
R89 B.n285 B.n16 585
R90 B.n284 B.n283 585
R91 B.n282 B.n17 585
R92 B.n281 B.n280 585
R93 B.n279 B.n18 585
R94 B.n278 B.n277 585
R95 B.n275 B.n19 585
R96 B.n274 B.n273 585
R97 B.n272 B.n22 585
R98 B.n271 B.n270 585
R99 B.n269 B.n23 585
R100 B.n268 B.n267 585
R101 B.n266 B.n24 585
R102 B.n265 B.n264 585
R103 B.n263 B.n25 585
R104 B.n262 B.n261 585
R105 B.n260 B.n259 585
R106 B.n258 B.n29 585
R107 B.n257 B.n256 585
R108 B.n255 B.n30 585
R109 B.n254 B.n253 585
R110 B.n252 B.n31 585
R111 B.n251 B.n250 585
R112 B.n249 B.n32 585
R113 B.n248 B.n247 585
R114 B.n246 B.n33 585
R115 B.n245 B.n244 585
R116 B.n243 B.n34 585
R117 B.n242 B.n241 585
R118 B.n240 B.n35 585
R119 B.n239 B.n238 585
R120 B.n300 B.n11 585
R121 B.n302 B.n301 585
R122 B.n303 B.n10 585
R123 B.n305 B.n304 585
R124 B.n306 B.n9 585
R125 B.n308 B.n307 585
R126 B.n309 B.n8 585
R127 B.n311 B.n310 585
R128 B.n312 B.n7 585
R129 B.n314 B.n313 585
R130 B.n315 B.n6 585
R131 B.n317 B.n316 585
R132 B.n318 B.n5 585
R133 B.n320 B.n319 585
R134 B.n321 B.n4 585
R135 B.n323 B.n322 585
R136 B.n324 B.n3 585
R137 B.n326 B.n325 585
R138 B.n327 B.n0 585
R139 B.n2 B.n1 585
R140 B.n88 B.n87 585
R141 B.n89 B.n86 585
R142 B.n91 B.n90 585
R143 B.n92 B.n85 585
R144 B.n94 B.n93 585
R145 B.n95 B.n84 585
R146 B.n97 B.n96 585
R147 B.n98 B.n83 585
R148 B.n100 B.n99 585
R149 B.n101 B.n82 585
R150 B.n103 B.n102 585
R151 B.n104 B.n81 585
R152 B.n106 B.n105 585
R153 B.n107 B.n80 585
R154 B.n109 B.n108 585
R155 B.n110 B.n79 585
R156 B.n112 B.n111 585
R157 B.n113 B.n78 585
R158 B.n114 B.n113 535.745
R159 B.n178 B.n177 535.745
R160 B.n238 B.n237 535.745
R161 B.n298 B.n11 535.745
R162 B.n64 B.t1 260.858
R163 B.n26 B.t8 260.858
R164 B.n135 B.t4 260.858
R165 B.n20 B.t11 260.858
R166 B.n329 B.n328 256.663
R167 B.n135 B.t3 251.531
R168 B.n64 B.t0 251.531
R169 B.n26 B.t6 251.531
R170 B.n20 B.t9 251.531
R171 B.n328 B.n327 235.042
R172 B.n328 B.n2 235.042
R173 B.n65 B.t2 223.04
R174 B.n27 B.t7 223.04
R175 B.n136 B.t5 223.04
R176 B.n21 B.t10 223.04
R177 B.n114 B.n77 163.367
R178 B.n118 B.n77 163.367
R179 B.n119 B.n118 163.367
R180 B.n120 B.n119 163.367
R181 B.n120 B.n75 163.367
R182 B.n124 B.n75 163.367
R183 B.n125 B.n124 163.367
R184 B.n126 B.n125 163.367
R185 B.n126 B.n73 163.367
R186 B.n130 B.n73 163.367
R187 B.n131 B.n130 163.367
R188 B.n132 B.n131 163.367
R189 B.n132 B.n71 163.367
R190 B.n139 B.n71 163.367
R191 B.n140 B.n139 163.367
R192 B.n141 B.n140 163.367
R193 B.n141 B.n69 163.367
R194 B.n145 B.n69 163.367
R195 B.n146 B.n145 163.367
R196 B.n147 B.n146 163.367
R197 B.n147 B.n67 163.367
R198 B.n151 B.n67 163.367
R199 B.n152 B.n151 163.367
R200 B.n153 B.n152 163.367
R201 B.n153 B.n63 163.367
R202 B.n158 B.n63 163.367
R203 B.n159 B.n158 163.367
R204 B.n160 B.n159 163.367
R205 B.n160 B.n61 163.367
R206 B.n164 B.n61 163.367
R207 B.n165 B.n164 163.367
R208 B.n166 B.n165 163.367
R209 B.n166 B.n59 163.367
R210 B.n170 B.n59 163.367
R211 B.n171 B.n170 163.367
R212 B.n172 B.n171 163.367
R213 B.n172 B.n57 163.367
R214 B.n176 B.n57 163.367
R215 B.n177 B.n176 163.367
R216 B.n237 B.n236 163.367
R217 B.n236 B.n37 163.367
R218 B.n232 B.n37 163.367
R219 B.n232 B.n231 163.367
R220 B.n231 B.n230 163.367
R221 B.n230 B.n39 163.367
R222 B.n226 B.n39 163.367
R223 B.n226 B.n225 163.367
R224 B.n225 B.n224 163.367
R225 B.n224 B.n41 163.367
R226 B.n220 B.n41 163.367
R227 B.n220 B.n219 163.367
R228 B.n219 B.n218 163.367
R229 B.n218 B.n43 163.367
R230 B.n214 B.n43 163.367
R231 B.n214 B.n213 163.367
R232 B.n213 B.n212 163.367
R233 B.n212 B.n45 163.367
R234 B.n208 B.n45 163.367
R235 B.n208 B.n207 163.367
R236 B.n207 B.n206 163.367
R237 B.n206 B.n47 163.367
R238 B.n202 B.n47 163.367
R239 B.n202 B.n201 163.367
R240 B.n201 B.n200 163.367
R241 B.n200 B.n49 163.367
R242 B.n196 B.n49 163.367
R243 B.n196 B.n195 163.367
R244 B.n195 B.n194 163.367
R245 B.n194 B.n51 163.367
R246 B.n190 B.n51 163.367
R247 B.n190 B.n189 163.367
R248 B.n189 B.n188 163.367
R249 B.n188 B.n53 163.367
R250 B.n184 B.n53 163.367
R251 B.n184 B.n183 163.367
R252 B.n183 B.n182 163.367
R253 B.n182 B.n55 163.367
R254 B.n178 B.n55 163.367
R255 B.n298 B.n297 163.367
R256 B.n297 B.n296 163.367
R257 B.n296 B.n13 163.367
R258 B.n292 B.n13 163.367
R259 B.n292 B.n291 163.367
R260 B.n291 B.n290 163.367
R261 B.n290 B.n15 163.367
R262 B.n286 B.n15 163.367
R263 B.n286 B.n285 163.367
R264 B.n285 B.n284 163.367
R265 B.n284 B.n17 163.367
R266 B.n280 B.n17 163.367
R267 B.n280 B.n279 163.367
R268 B.n279 B.n278 163.367
R269 B.n278 B.n19 163.367
R270 B.n273 B.n19 163.367
R271 B.n273 B.n272 163.367
R272 B.n272 B.n271 163.367
R273 B.n271 B.n23 163.367
R274 B.n267 B.n23 163.367
R275 B.n267 B.n266 163.367
R276 B.n266 B.n265 163.367
R277 B.n265 B.n25 163.367
R278 B.n261 B.n25 163.367
R279 B.n261 B.n260 163.367
R280 B.n260 B.n29 163.367
R281 B.n256 B.n29 163.367
R282 B.n256 B.n255 163.367
R283 B.n255 B.n254 163.367
R284 B.n254 B.n31 163.367
R285 B.n250 B.n31 163.367
R286 B.n250 B.n249 163.367
R287 B.n249 B.n248 163.367
R288 B.n248 B.n33 163.367
R289 B.n244 B.n33 163.367
R290 B.n244 B.n243 163.367
R291 B.n243 B.n242 163.367
R292 B.n242 B.n35 163.367
R293 B.n238 B.n35 163.367
R294 B.n302 B.n11 163.367
R295 B.n303 B.n302 163.367
R296 B.n304 B.n303 163.367
R297 B.n304 B.n9 163.367
R298 B.n308 B.n9 163.367
R299 B.n309 B.n308 163.367
R300 B.n310 B.n309 163.367
R301 B.n310 B.n7 163.367
R302 B.n314 B.n7 163.367
R303 B.n315 B.n314 163.367
R304 B.n316 B.n315 163.367
R305 B.n316 B.n5 163.367
R306 B.n320 B.n5 163.367
R307 B.n321 B.n320 163.367
R308 B.n322 B.n321 163.367
R309 B.n322 B.n3 163.367
R310 B.n326 B.n3 163.367
R311 B.n327 B.n326 163.367
R312 B.n88 B.n2 163.367
R313 B.n89 B.n88 163.367
R314 B.n90 B.n89 163.367
R315 B.n90 B.n85 163.367
R316 B.n94 B.n85 163.367
R317 B.n95 B.n94 163.367
R318 B.n96 B.n95 163.367
R319 B.n96 B.n83 163.367
R320 B.n100 B.n83 163.367
R321 B.n101 B.n100 163.367
R322 B.n102 B.n101 163.367
R323 B.n102 B.n81 163.367
R324 B.n106 B.n81 163.367
R325 B.n107 B.n106 163.367
R326 B.n108 B.n107 163.367
R327 B.n108 B.n79 163.367
R328 B.n112 B.n79 163.367
R329 B.n113 B.n112 163.367
R330 B.n137 B.n136 59.5399
R331 B.n155 B.n65 59.5399
R332 B.n28 B.n27 59.5399
R333 B.n276 B.n21 59.5399
R334 B.n136 B.n135 37.8187
R335 B.n65 B.n64 37.8187
R336 B.n27 B.n26 37.8187
R337 B.n21 B.n20 37.8187
R338 B.n300 B.n299 34.8103
R339 B.n239 B.n36 34.8103
R340 B.n115 B.n78 34.8103
R341 B.n179 B.n56 34.8103
R342 B B.n329 18.0485
R343 B.n301 B.n300 10.6151
R344 B.n301 B.n10 10.6151
R345 B.n305 B.n10 10.6151
R346 B.n306 B.n305 10.6151
R347 B.n307 B.n306 10.6151
R348 B.n307 B.n8 10.6151
R349 B.n311 B.n8 10.6151
R350 B.n312 B.n311 10.6151
R351 B.n313 B.n312 10.6151
R352 B.n313 B.n6 10.6151
R353 B.n317 B.n6 10.6151
R354 B.n318 B.n317 10.6151
R355 B.n319 B.n318 10.6151
R356 B.n319 B.n4 10.6151
R357 B.n323 B.n4 10.6151
R358 B.n324 B.n323 10.6151
R359 B.n325 B.n324 10.6151
R360 B.n325 B.n0 10.6151
R361 B.n299 B.n12 10.6151
R362 B.n295 B.n12 10.6151
R363 B.n295 B.n294 10.6151
R364 B.n294 B.n293 10.6151
R365 B.n293 B.n14 10.6151
R366 B.n289 B.n14 10.6151
R367 B.n289 B.n288 10.6151
R368 B.n288 B.n287 10.6151
R369 B.n287 B.n16 10.6151
R370 B.n283 B.n16 10.6151
R371 B.n283 B.n282 10.6151
R372 B.n282 B.n281 10.6151
R373 B.n281 B.n18 10.6151
R374 B.n277 B.n18 10.6151
R375 B.n275 B.n274 10.6151
R376 B.n274 B.n22 10.6151
R377 B.n270 B.n22 10.6151
R378 B.n270 B.n269 10.6151
R379 B.n269 B.n268 10.6151
R380 B.n268 B.n24 10.6151
R381 B.n264 B.n24 10.6151
R382 B.n264 B.n263 10.6151
R383 B.n263 B.n262 10.6151
R384 B.n259 B.n258 10.6151
R385 B.n258 B.n257 10.6151
R386 B.n257 B.n30 10.6151
R387 B.n253 B.n30 10.6151
R388 B.n253 B.n252 10.6151
R389 B.n252 B.n251 10.6151
R390 B.n251 B.n32 10.6151
R391 B.n247 B.n32 10.6151
R392 B.n247 B.n246 10.6151
R393 B.n246 B.n245 10.6151
R394 B.n245 B.n34 10.6151
R395 B.n241 B.n34 10.6151
R396 B.n241 B.n240 10.6151
R397 B.n240 B.n239 10.6151
R398 B.n235 B.n36 10.6151
R399 B.n235 B.n234 10.6151
R400 B.n234 B.n233 10.6151
R401 B.n233 B.n38 10.6151
R402 B.n229 B.n38 10.6151
R403 B.n229 B.n228 10.6151
R404 B.n228 B.n227 10.6151
R405 B.n227 B.n40 10.6151
R406 B.n223 B.n40 10.6151
R407 B.n223 B.n222 10.6151
R408 B.n222 B.n221 10.6151
R409 B.n221 B.n42 10.6151
R410 B.n217 B.n42 10.6151
R411 B.n217 B.n216 10.6151
R412 B.n216 B.n215 10.6151
R413 B.n215 B.n44 10.6151
R414 B.n211 B.n44 10.6151
R415 B.n211 B.n210 10.6151
R416 B.n210 B.n209 10.6151
R417 B.n209 B.n46 10.6151
R418 B.n205 B.n46 10.6151
R419 B.n205 B.n204 10.6151
R420 B.n204 B.n203 10.6151
R421 B.n203 B.n48 10.6151
R422 B.n199 B.n48 10.6151
R423 B.n199 B.n198 10.6151
R424 B.n198 B.n197 10.6151
R425 B.n197 B.n50 10.6151
R426 B.n193 B.n50 10.6151
R427 B.n193 B.n192 10.6151
R428 B.n192 B.n191 10.6151
R429 B.n191 B.n52 10.6151
R430 B.n187 B.n52 10.6151
R431 B.n187 B.n186 10.6151
R432 B.n186 B.n185 10.6151
R433 B.n185 B.n54 10.6151
R434 B.n181 B.n54 10.6151
R435 B.n181 B.n180 10.6151
R436 B.n180 B.n179 10.6151
R437 B.n87 B.n1 10.6151
R438 B.n87 B.n86 10.6151
R439 B.n91 B.n86 10.6151
R440 B.n92 B.n91 10.6151
R441 B.n93 B.n92 10.6151
R442 B.n93 B.n84 10.6151
R443 B.n97 B.n84 10.6151
R444 B.n98 B.n97 10.6151
R445 B.n99 B.n98 10.6151
R446 B.n99 B.n82 10.6151
R447 B.n103 B.n82 10.6151
R448 B.n104 B.n103 10.6151
R449 B.n105 B.n104 10.6151
R450 B.n105 B.n80 10.6151
R451 B.n109 B.n80 10.6151
R452 B.n110 B.n109 10.6151
R453 B.n111 B.n110 10.6151
R454 B.n111 B.n78 10.6151
R455 B.n116 B.n115 10.6151
R456 B.n117 B.n116 10.6151
R457 B.n117 B.n76 10.6151
R458 B.n121 B.n76 10.6151
R459 B.n122 B.n121 10.6151
R460 B.n123 B.n122 10.6151
R461 B.n123 B.n74 10.6151
R462 B.n127 B.n74 10.6151
R463 B.n128 B.n127 10.6151
R464 B.n129 B.n128 10.6151
R465 B.n129 B.n72 10.6151
R466 B.n133 B.n72 10.6151
R467 B.n134 B.n133 10.6151
R468 B.n138 B.n134 10.6151
R469 B.n142 B.n70 10.6151
R470 B.n143 B.n142 10.6151
R471 B.n144 B.n143 10.6151
R472 B.n144 B.n68 10.6151
R473 B.n148 B.n68 10.6151
R474 B.n149 B.n148 10.6151
R475 B.n150 B.n149 10.6151
R476 B.n150 B.n66 10.6151
R477 B.n154 B.n66 10.6151
R478 B.n157 B.n156 10.6151
R479 B.n157 B.n62 10.6151
R480 B.n161 B.n62 10.6151
R481 B.n162 B.n161 10.6151
R482 B.n163 B.n162 10.6151
R483 B.n163 B.n60 10.6151
R484 B.n167 B.n60 10.6151
R485 B.n168 B.n167 10.6151
R486 B.n169 B.n168 10.6151
R487 B.n169 B.n58 10.6151
R488 B.n173 B.n58 10.6151
R489 B.n174 B.n173 10.6151
R490 B.n175 B.n174 10.6151
R491 B.n175 B.n56 10.6151
R492 B.n277 B.n276 9.36635
R493 B.n259 B.n28 9.36635
R494 B.n138 B.n137 9.36635
R495 B.n156 B.n155 9.36635
R496 B.n329 B.n0 8.11757
R497 B.n329 B.n1 8.11757
R498 B.n276 B.n275 1.24928
R499 B.n262 B.n28 1.24928
R500 B.n137 B.n70 1.24928
R501 B.n155 B.n154 1.24928
R502 VP.n0 VP.t1 139.825
R503 VP.n0 VP.t0 104.532
R504 VP VP.n0 0.241678
R505 VTAIL.n58 VTAIL.n48 756.745
R506 VTAIL.n10 VTAIL.n0 756.745
R507 VTAIL.n42 VTAIL.n32 756.745
R508 VTAIL.n26 VTAIL.n16 756.745
R509 VTAIL.n52 VTAIL.n51 585
R510 VTAIL.n57 VTAIL.n56 585
R511 VTAIL.n59 VTAIL.n58 585
R512 VTAIL.n4 VTAIL.n3 585
R513 VTAIL.n9 VTAIL.n8 585
R514 VTAIL.n11 VTAIL.n10 585
R515 VTAIL.n43 VTAIL.n42 585
R516 VTAIL.n41 VTAIL.n40 585
R517 VTAIL.n36 VTAIL.n35 585
R518 VTAIL.n27 VTAIL.n26 585
R519 VTAIL.n25 VTAIL.n24 585
R520 VTAIL.n20 VTAIL.n19 585
R521 VTAIL.n53 VTAIL.t0 336.901
R522 VTAIL.n5 VTAIL.t2 336.901
R523 VTAIL.n37 VTAIL.t3 336.901
R524 VTAIL.n21 VTAIL.t1 336.901
R525 VTAIL.n57 VTAIL.n51 171.744
R526 VTAIL.n58 VTAIL.n57 171.744
R527 VTAIL.n9 VTAIL.n3 171.744
R528 VTAIL.n10 VTAIL.n9 171.744
R529 VTAIL.n42 VTAIL.n41 171.744
R530 VTAIL.n41 VTAIL.n35 171.744
R531 VTAIL.n26 VTAIL.n25 171.744
R532 VTAIL.n25 VTAIL.n19 171.744
R533 VTAIL.t0 VTAIL.n51 85.8723
R534 VTAIL.t2 VTAIL.n3 85.8723
R535 VTAIL.t3 VTAIL.n35 85.8723
R536 VTAIL.t1 VTAIL.n19 85.8723
R537 VTAIL.n63 VTAIL.n62 31.2157
R538 VTAIL.n15 VTAIL.n14 31.2157
R539 VTAIL.n47 VTAIL.n46 31.2157
R540 VTAIL.n31 VTAIL.n30 31.2157
R541 VTAIL.n31 VTAIL.n15 18.3755
R542 VTAIL.n63 VTAIL.n47 16.6945
R543 VTAIL.n53 VTAIL.n52 16.193
R544 VTAIL.n5 VTAIL.n4 16.193
R545 VTAIL.n37 VTAIL.n36 16.193
R546 VTAIL.n21 VTAIL.n20 16.193
R547 VTAIL.n56 VTAIL.n55 12.8005
R548 VTAIL.n8 VTAIL.n7 12.8005
R549 VTAIL.n40 VTAIL.n39 12.8005
R550 VTAIL.n24 VTAIL.n23 12.8005
R551 VTAIL.n59 VTAIL.n50 12.0247
R552 VTAIL.n11 VTAIL.n2 12.0247
R553 VTAIL.n43 VTAIL.n34 12.0247
R554 VTAIL.n27 VTAIL.n18 12.0247
R555 VTAIL.n60 VTAIL.n48 11.249
R556 VTAIL.n12 VTAIL.n0 11.249
R557 VTAIL.n44 VTAIL.n32 11.249
R558 VTAIL.n28 VTAIL.n16 11.249
R559 VTAIL.n62 VTAIL.n61 9.45567
R560 VTAIL.n14 VTAIL.n13 9.45567
R561 VTAIL.n46 VTAIL.n45 9.45567
R562 VTAIL.n30 VTAIL.n29 9.45567
R563 VTAIL.n61 VTAIL.n60 9.3005
R564 VTAIL.n50 VTAIL.n49 9.3005
R565 VTAIL.n55 VTAIL.n54 9.3005
R566 VTAIL.n13 VTAIL.n12 9.3005
R567 VTAIL.n2 VTAIL.n1 9.3005
R568 VTAIL.n7 VTAIL.n6 9.3005
R569 VTAIL.n45 VTAIL.n44 9.3005
R570 VTAIL.n34 VTAIL.n33 9.3005
R571 VTAIL.n39 VTAIL.n38 9.3005
R572 VTAIL.n29 VTAIL.n28 9.3005
R573 VTAIL.n18 VTAIL.n17 9.3005
R574 VTAIL.n23 VTAIL.n22 9.3005
R575 VTAIL.n38 VTAIL.n37 3.91276
R576 VTAIL.n22 VTAIL.n21 3.91276
R577 VTAIL.n54 VTAIL.n53 3.91276
R578 VTAIL.n6 VTAIL.n5 3.91276
R579 VTAIL.n62 VTAIL.n48 2.71565
R580 VTAIL.n14 VTAIL.n0 2.71565
R581 VTAIL.n46 VTAIL.n32 2.71565
R582 VTAIL.n30 VTAIL.n16 2.71565
R583 VTAIL.n60 VTAIL.n59 1.93989
R584 VTAIL.n12 VTAIL.n11 1.93989
R585 VTAIL.n44 VTAIL.n43 1.93989
R586 VTAIL.n28 VTAIL.n27 1.93989
R587 VTAIL.n47 VTAIL.n31 1.31084
R588 VTAIL.n56 VTAIL.n50 1.16414
R589 VTAIL.n8 VTAIL.n2 1.16414
R590 VTAIL.n40 VTAIL.n34 1.16414
R591 VTAIL.n24 VTAIL.n18 1.16414
R592 VTAIL VTAIL.n15 0.948776
R593 VTAIL.n55 VTAIL.n52 0.388379
R594 VTAIL.n7 VTAIL.n4 0.388379
R595 VTAIL.n39 VTAIL.n36 0.388379
R596 VTAIL.n23 VTAIL.n20 0.388379
R597 VTAIL VTAIL.n63 0.362569
R598 VTAIL.n54 VTAIL.n49 0.155672
R599 VTAIL.n61 VTAIL.n49 0.155672
R600 VTAIL.n6 VTAIL.n1 0.155672
R601 VTAIL.n13 VTAIL.n1 0.155672
R602 VTAIL.n45 VTAIL.n33 0.155672
R603 VTAIL.n38 VTAIL.n33 0.155672
R604 VTAIL.n29 VTAIL.n17 0.155672
R605 VTAIL.n22 VTAIL.n17 0.155672
R606 VDD1.n10 VDD1.n0 756.745
R607 VDD1.n25 VDD1.n15 756.745
R608 VDD1.n11 VDD1.n10 585
R609 VDD1.n9 VDD1.n8 585
R610 VDD1.n4 VDD1.n3 585
R611 VDD1.n19 VDD1.n18 585
R612 VDD1.n24 VDD1.n23 585
R613 VDD1.n26 VDD1.n25 585
R614 VDD1.n5 VDD1.t0 336.901
R615 VDD1.n20 VDD1.t1 336.901
R616 VDD1.n10 VDD1.n9 171.744
R617 VDD1.n9 VDD1.n3 171.744
R618 VDD1.n24 VDD1.n18 171.744
R619 VDD1.n25 VDD1.n24 171.744
R620 VDD1.t0 VDD1.n3 85.8723
R621 VDD1.t1 VDD1.n18 85.8723
R622 VDD1 VDD1.n29 78.5076
R623 VDD1 VDD1.n14 48.3729
R624 VDD1.n5 VDD1.n4 16.193
R625 VDD1.n20 VDD1.n19 16.193
R626 VDD1.n8 VDD1.n7 12.8005
R627 VDD1.n23 VDD1.n22 12.8005
R628 VDD1.n11 VDD1.n2 12.0247
R629 VDD1.n26 VDD1.n17 12.0247
R630 VDD1.n12 VDD1.n0 11.249
R631 VDD1.n27 VDD1.n15 11.249
R632 VDD1.n14 VDD1.n13 9.45567
R633 VDD1.n29 VDD1.n28 9.45567
R634 VDD1.n13 VDD1.n12 9.3005
R635 VDD1.n2 VDD1.n1 9.3005
R636 VDD1.n7 VDD1.n6 9.3005
R637 VDD1.n28 VDD1.n27 9.3005
R638 VDD1.n17 VDD1.n16 9.3005
R639 VDD1.n22 VDD1.n21 9.3005
R640 VDD1.n6 VDD1.n5 3.91276
R641 VDD1.n21 VDD1.n20 3.91276
R642 VDD1.n14 VDD1.n0 2.71565
R643 VDD1.n29 VDD1.n15 2.71565
R644 VDD1.n12 VDD1.n11 1.93989
R645 VDD1.n27 VDD1.n26 1.93989
R646 VDD1.n8 VDD1.n2 1.16414
R647 VDD1.n23 VDD1.n17 1.16414
R648 VDD1.n7 VDD1.n4 0.388379
R649 VDD1.n22 VDD1.n19 0.388379
R650 VDD1.n13 VDD1.n1 0.155672
R651 VDD1.n6 VDD1.n1 0.155672
R652 VDD1.n21 VDD1.n16 0.155672
R653 VDD1.n28 VDD1.n16 0.155672
R654 VN VN.t0 140.016
R655 VN VN.t1 104.773
R656 VDD2.n25 VDD2.n15 756.745
R657 VDD2.n10 VDD2.n0 756.745
R658 VDD2.n26 VDD2.n25 585
R659 VDD2.n24 VDD2.n23 585
R660 VDD2.n19 VDD2.n18 585
R661 VDD2.n4 VDD2.n3 585
R662 VDD2.n9 VDD2.n8 585
R663 VDD2.n11 VDD2.n10 585
R664 VDD2.n20 VDD2.t1 336.901
R665 VDD2.n5 VDD2.t0 336.901
R666 VDD2.n25 VDD2.n24 171.744
R667 VDD2.n24 VDD2.n18 171.744
R668 VDD2.n9 VDD2.n3 171.744
R669 VDD2.n10 VDD2.n9 171.744
R670 VDD2.t1 VDD2.n18 85.8723
R671 VDD2.t0 VDD2.n3 85.8723
R672 VDD2.n30 VDD2.n14 77.5625
R673 VDD2.n30 VDD2.n29 47.8944
R674 VDD2.n20 VDD2.n19 16.193
R675 VDD2.n5 VDD2.n4 16.193
R676 VDD2.n23 VDD2.n22 12.8005
R677 VDD2.n8 VDD2.n7 12.8005
R678 VDD2.n26 VDD2.n17 12.0247
R679 VDD2.n11 VDD2.n2 12.0247
R680 VDD2.n27 VDD2.n15 11.249
R681 VDD2.n12 VDD2.n0 11.249
R682 VDD2.n29 VDD2.n28 9.45567
R683 VDD2.n14 VDD2.n13 9.45567
R684 VDD2.n28 VDD2.n27 9.3005
R685 VDD2.n17 VDD2.n16 9.3005
R686 VDD2.n22 VDD2.n21 9.3005
R687 VDD2.n13 VDD2.n12 9.3005
R688 VDD2.n2 VDD2.n1 9.3005
R689 VDD2.n7 VDD2.n6 9.3005
R690 VDD2.n21 VDD2.n20 3.91276
R691 VDD2.n6 VDD2.n5 3.91276
R692 VDD2.n29 VDD2.n15 2.71565
R693 VDD2.n14 VDD2.n0 2.71565
R694 VDD2.n27 VDD2.n26 1.93989
R695 VDD2.n12 VDD2.n11 1.93989
R696 VDD2.n23 VDD2.n17 1.16414
R697 VDD2.n8 VDD2.n2 1.16414
R698 VDD2 VDD2.n30 0.478948
R699 VDD2.n22 VDD2.n19 0.388379
R700 VDD2.n7 VDD2.n4 0.388379
R701 VDD2.n28 VDD2.n16 0.155672
R702 VDD2.n21 VDD2.n16 0.155672
R703 VDD2.n6 VDD2.n1 0.155672
R704 VDD2.n13 VDD2.n1 0.155672
C0 B w_n1750_n1582# 5.24977f
C1 VDD1 VN 0.152695f
C2 VN B 0.767019f
C3 VDD2 VP 0.296543f
C4 VP VTAIL 0.93259f
C5 VDD2 VTAIL 2.48726f
C6 VDD1 B 0.881553f
C7 VP w_n1750_n1582# 2.37528f
C8 VDD2 w_n1750_n1582# 1.04676f
C9 w_n1750_n1582# VTAIL 1.42129f
C10 VN VP 3.35214f
C11 VDD2 VN 0.835387f
C12 VN VTAIL 0.918408f
C13 VDD1 VP 0.977682f
C14 VDD1 VDD2 0.558125f
C15 VDD1 VTAIL 2.44155f
C16 VP B 1.12569f
C17 VN w_n1750_n1582# 2.15669f
C18 VDD2 B 0.903124f
C19 B VTAIL 1.34427f
C20 VDD1 w_n1750_n1582# 1.03312f
C21 VDD2 VSUBS 0.497459f
C22 VDD1 VSUBS 1.881966f
C23 VTAIL VSUBS 0.369016f
C24 VN VSUBS 4.91441f
C25 VP VSUBS 0.969294f
C26 B VSUBS 2.29325f
C27 w_n1750_n1582# VSUBS 35.049f
C28 VDD2.n0 VSUBS 0.016199f
C29 VDD2.n1 VSUBS 0.01611f
C30 VDD2.n2 VSUBS 0.008657f
C31 VDD2.n3 VSUBS 0.015346f
C32 VDD2.n4 VSUBS 0.012632f
C33 VDD2.t0 VSUBS 0.044684f
C34 VDD2.n5 VSUBS 0.056992f
C35 VDD2.n6 VSUBS 0.155055f
C36 VDD2.n7 VSUBS 0.008657f
C37 VDD2.n8 VSUBS 0.009166f
C38 VDD2.n9 VSUBS 0.020461f
C39 VDD2.n10 VSUBS 0.044419f
C40 VDD2.n11 VSUBS 0.009166f
C41 VDD2.n12 VSUBS 0.008657f
C42 VDD2.n13 VSUBS 0.036136f
C43 VDD2.n14 VSUBS 0.254393f
C44 VDD2.n15 VSUBS 0.016199f
C45 VDD2.n16 VSUBS 0.01611f
C46 VDD2.n17 VSUBS 0.008657f
C47 VDD2.n18 VSUBS 0.015346f
C48 VDD2.n19 VSUBS 0.012632f
C49 VDD2.t1 VSUBS 0.044684f
C50 VDD2.n20 VSUBS 0.056992f
C51 VDD2.n21 VSUBS 0.155055f
C52 VDD2.n22 VSUBS 0.008657f
C53 VDD2.n23 VSUBS 0.009166f
C54 VDD2.n24 VSUBS 0.020461f
C55 VDD2.n25 VSUBS 0.044419f
C56 VDD2.n26 VSUBS 0.009166f
C57 VDD2.n27 VSUBS 0.008657f
C58 VDD2.n28 VSUBS 0.036136f
C59 VDD2.n29 VSUBS 0.033209f
C60 VDD2.n30 VSUBS 1.21882f
C61 VN.t1 VSUBS 0.906383f
C62 VN.t0 VSUBS 1.3766f
C63 VDD1.n0 VSUBS 0.01519f
C64 VDD1.n1 VSUBS 0.015106f
C65 VDD1.n2 VSUBS 0.008117f
C66 VDD1.n3 VSUBS 0.014389f
C67 VDD1.n4 VSUBS 0.011845f
C68 VDD1.t0 VSUBS 0.0419f
C69 VDD1.n5 VSUBS 0.05344f
C70 VDD1.n6 VSUBS 0.145392f
C71 VDD1.n7 VSUBS 0.008117f
C72 VDD1.n8 VSUBS 0.008595f
C73 VDD1.n9 VSUBS 0.019186f
C74 VDD1.n10 VSUBS 0.041651f
C75 VDD1.n11 VSUBS 0.008595f
C76 VDD1.n12 VSUBS 0.008117f
C77 VDD1.n13 VSUBS 0.033884f
C78 VDD1.n14 VSUBS 0.031652f
C79 VDD1.n15 VSUBS 0.01519f
C80 VDD1.n16 VSUBS 0.015106f
C81 VDD1.n17 VSUBS 0.008117f
C82 VDD1.n18 VSUBS 0.014389f
C83 VDD1.n19 VSUBS 0.011845f
C84 VDD1.t1 VSUBS 0.0419f
C85 VDD1.n20 VSUBS 0.05344f
C86 VDD1.n21 VSUBS 0.145392f
C87 VDD1.n22 VSUBS 0.008117f
C88 VDD1.n23 VSUBS 0.008595f
C89 VDD1.n24 VSUBS 0.019186f
C90 VDD1.n25 VSUBS 0.041651f
C91 VDD1.n26 VSUBS 0.008595f
C92 VDD1.n27 VSUBS 0.008117f
C93 VDD1.n28 VSUBS 0.033884f
C94 VDD1.n29 VSUBS 0.258886f
C95 VTAIL.n0 VSUBS 0.018852f
C96 VTAIL.n1 VSUBS 0.018747f
C97 VTAIL.n2 VSUBS 0.010074f
C98 VTAIL.n3 VSUBS 0.017858f
C99 VTAIL.n4 VSUBS 0.0147f
C100 VTAIL.t2 VSUBS 0.052f
C101 VTAIL.n5 VSUBS 0.066322f
C102 VTAIL.n6 VSUBS 0.18044f
C103 VTAIL.n7 VSUBS 0.010074f
C104 VTAIL.n8 VSUBS 0.010666f
C105 VTAIL.n9 VSUBS 0.023811f
C106 VTAIL.n10 VSUBS 0.051692f
C107 VTAIL.n11 VSUBS 0.010666f
C108 VTAIL.n12 VSUBS 0.010074f
C109 VTAIL.n13 VSUBS 0.042052f
C110 VTAIL.n14 VSUBS 0.025691f
C111 VTAIL.n15 VSUBS 0.690184f
C112 VTAIL.n16 VSUBS 0.018852f
C113 VTAIL.n17 VSUBS 0.018747f
C114 VTAIL.n18 VSUBS 0.010074f
C115 VTAIL.n19 VSUBS 0.017858f
C116 VTAIL.n20 VSUBS 0.0147f
C117 VTAIL.t1 VSUBS 0.052f
C118 VTAIL.n21 VSUBS 0.066322f
C119 VTAIL.n22 VSUBS 0.18044f
C120 VTAIL.n23 VSUBS 0.010074f
C121 VTAIL.n24 VSUBS 0.010666f
C122 VTAIL.n25 VSUBS 0.023811f
C123 VTAIL.n26 VSUBS 0.051692f
C124 VTAIL.n27 VSUBS 0.010666f
C125 VTAIL.n28 VSUBS 0.010074f
C126 VTAIL.n29 VSUBS 0.042052f
C127 VTAIL.n30 VSUBS 0.025691f
C128 VTAIL.n31 VSUBS 0.712055f
C129 VTAIL.n32 VSUBS 0.018852f
C130 VTAIL.n33 VSUBS 0.018747f
C131 VTAIL.n34 VSUBS 0.010074f
C132 VTAIL.n35 VSUBS 0.017858f
C133 VTAIL.n36 VSUBS 0.0147f
C134 VTAIL.t3 VSUBS 0.052f
C135 VTAIL.n37 VSUBS 0.066322f
C136 VTAIL.n38 VSUBS 0.18044f
C137 VTAIL.n39 VSUBS 0.010074f
C138 VTAIL.n40 VSUBS 0.010666f
C139 VTAIL.n41 VSUBS 0.023811f
C140 VTAIL.n42 VSUBS 0.051692f
C141 VTAIL.n43 VSUBS 0.010666f
C142 VTAIL.n44 VSUBS 0.010074f
C143 VTAIL.n45 VSUBS 0.042052f
C144 VTAIL.n46 VSUBS 0.025691f
C145 VTAIL.n47 VSUBS 0.61051f
C146 VTAIL.n48 VSUBS 0.018852f
C147 VTAIL.n49 VSUBS 0.018747f
C148 VTAIL.n50 VSUBS 0.010074f
C149 VTAIL.n51 VSUBS 0.017858f
C150 VTAIL.n52 VSUBS 0.0147f
C151 VTAIL.t0 VSUBS 0.052f
C152 VTAIL.n53 VSUBS 0.066322f
C153 VTAIL.n54 VSUBS 0.18044f
C154 VTAIL.n55 VSUBS 0.010074f
C155 VTAIL.n56 VSUBS 0.010666f
C156 VTAIL.n57 VSUBS 0.023811f
C157 VTAIL.n58 VSUBS 0.051692f
C158 VTAIL.n59 VSUBS 0.010666f
C159 VTAIL.n60 VSUBS 0.010074f
C160 VTAIL.n61 VSUBS 0.042052f
C161 VTAIL.n62 VSUBS 0.025691f
C162 VTAIL.n63 VSUBS 0.553228f
C163 VP.t1 VSUBS 1.43537f
C164 VP.t0 VSUBS 0.949862f
C165 VP.n0 VSUBS 3.34263f
C166 B.n0 VSUBS 0.006985f
C167 B.n1 VSUBS 0.006985f
C168 B.n2 VSUBS 0.010331f
C169 B.n3 VSUBS 0.007917f
C170 B.n4 VSUBS 0.007917f
C171 B.n5 VSUBS 0.007917f
C172 B.n6 VSUBS 0.007917f
C173 B.n7 VSUBS 0.007917f
C174 B.n8 VSUBS 0.007917f
C175 B.n9 VSUBS 0.007917f
C176 B.n10 VSUBS 0.007917f
C177 B.n11 VSUBS 0.018952f
C178 B.n12 VSUBS 0.007917f
C179 B.n13 VSUBS 0.007917f
C180 B.n14 VSUBS 0.007917f
C181 B.n15 VSUBS 0.007917f
C182 B.n16 VSUBS 0.007917f
C183 B.n17 VSUBS 0.007917f
C184 B.n18 VSUBS 0.007917f
C185 B.n19 VSUBS 0.007917f
C186 B.t10 VSUBS 0.050859f
C187 B.t11 VSUBS 0.064137f
C188 B.t9 VSUBS 0.268881f
C189 B.n20 VSUBS 0.116333f
C190 B.n21 VSUBS 0.102879f
C191 B.n22 VSUBS 0.007917f
C192 B.n23 VSUBS 0.007917f
C193 B.n24 VSUBS 0.007917f
C194 B.n25 VSUBS 0.007917f
C195 B.t7 VSUBS 0.05086f
C196 B.t8 VSUBS 0.064138f
C197 B.t6 VSUBS 0.268881f
C198 B.n26 VSUBS 0.116333f
C199 B.n27 VSUBS 0.102878f
C200 B.n28 VSUBS 0.018342f
C201 B.n29 VSUBS 0.007917f
C202 B.n30 VSUBS 0.007917f
C203 B.n31 VSUBS 0.007917f
C204 B.n32 VSUBS 0.007917f
C205 B.n33 VSUBS 0.007917f
C206 B.n34 VSUBS 0.007917f
C207 B.n35 VSUBS 0.007917f
C208 B.n36 VSUBS 0.018952f
C209 B.n37 VSUBS 0.007917f
C210 B.n38 VSUBS 0.007917f
C211 B.n39 VSUBS 0.007917f
C212 B.n40 VSUBS 0.007917f
C213 B.n41 VSUBS 0.007917f
C214 B.n42 VSUBS 0.007917f
C215 B.n43 VSUBS 0.007917f
C216 B.n44 VSUBS 0.007917f
C217 B.n45 VSUBS 0.007917f
C218 B.n46 VSUBS 0.007917f
C219 B.n47 VSUBS 0.007917f
C220 B.n48 VSUBS 0.007917f
C221 B.n49 VSUBS 0.007917f
C222 B.n50 VSUBS 0.007917f
C223 B.n51 VSUBS 0.007917f
C224 B.n52 VSUBS 0.007917f
C225 B.n53 VSUBS 0.007917f
C226 B.n54 VSUBS 0.007917f
C227 B.n55 VSUBS 0.007917f
C228 B.n56 VSUBS 0.018823f
C229 B.n57 VSUBS 0.007917f
C230 B.n58 VSUBS 0.007917f
C231 B.n59 VSUBS 0.007917f
C232 B.n60 VSUBS 0.007917f
C233 B.n61 VSUBS 0.007917f
C234 B.n62 VSUBS 0.007917f
C235 B.n63 VSUBS 0.007917f
C236 B.t2 VSUBS 0.05086f
C237 B.t1 VSUBS 0.064138f
C238 B.t0 VSUBS 0.268881f
C239 B.n64 VSUBS 0.116333f
C240 B.n65 VSUBS 0.102878f
C241 B.n66 VSUBS 0.007917f
C242 B.n67 VSUBS 0.007917f
C243 B.n68 VSUBS 0.007917f
C244 B.n69 VSUBS 0.007917f
C245 B.n70 VSUBS 0.004424f
C246 B.n71 VSUBS 0.007917f
C247 B.n72 VSUBS 0.007917f
C248 B.n73 VSUBS 0.007917f
C249 B.n74 VSUBS 0.007917f
C250 B.n75 VSUBS 0.007917f
C251 B.n76 VSUBS 0.007917f
C252 B.n77 VSUBS 0.007917f
C253 B.n78 VSUBS 0.018952f
C254 B.n79 VSUBS 0.007917f
C255 B.n80 VSUBS 0.007917f
C256 B.n81 VSUBS 0.007917f
C257 B.n82 VSUBS 0.007917f
C258 B.n83 VSUBS 0.007917f
C259 B.n84 VSUBS 0.007917f
C260 B.n85 VSUBS 0.007917f
C261 B.n86 VSUBS 0.007917f
C262 B.n87 VSUBS 0.007917f
C263 B.n88 VSUBS 0.007917f
C264 B.n89 VSUBS 0.007917f
C265 B.n90 VSUBS 0.007917f
C266 B.n91 VSUBS 0.007917f
C267 B.n92 VSUBS 0.007917f
C268 B.n93 VSUBS 0.007917f
C269 B.n94 VSUBS 0.007917f
C270 B.n95 VSUBS 0.007917f
C271 B.n96 VSUBS 0.007917f
C272 B.n97 VSUBS 0.007917f
C273 B.n98 VSUBS 0.007917f
C274 B.n99 VSUBS 0.007917f
C275 B.n100 VSUBS 0.007917f
C276 B.n101 VSUBS 0.007917f
C277 B.n102 VSUBS 0.007917f
C278 B.n103 VSUBS 0.007917f
C279 B.n104 VSUBS 0.007917f
C280 B.n105 VSUBS 0.007917f
C281 B.n106 VSUBS 0.007917f
C282 B.n107 VSUBS 0.007917f
C283 B.n108 VSUBS 0.007917f
C284 B.n109 VSUBS 0.007917f
C285 B.n110 VSUBS 0.007917f
C286 B.n111 VSUBS 0.007917f
C287 B.n112 VSUBS 0.007917f
C288 B.n113 VSUBS 0.018952f
C289 B.n114 VSUBS 0.019701f
C290 B.n115 VSUBS 0.019701f
C291 B.n116 VSUBS 0.007917f
C292 B.n117 VSUBS 0.007917f
C293 B.n118 VSUBS 0.007917f
C294 B.n119 VSUBS 0.007917f
C295 B.n120 VSUBS 0.007917f
C296 B.n121 VSUBS 0.007917f
C297 B.n122 VSUBS 0.007917f
C298 B.n123 VSUBS 0.007917f
C299 B.n124 VSUBS 0.007917f
C300 B.n125 VSUBS 0.007917f
C301 B.n126 VSUBS 0.007917f
C302 B.n127 VSUBS 0.007917f
C303 B.n128 VSUBS 0.007917f
C304 B.n129 VSUBS 0.007917f
C305 B.n130 VSUBS 0.007917f
C306 B.n131 VSUBS 0.007917f
C307 B.n132 VSUBS 0.007917f
C308 B.n133 VSUBS 0.007917f
C309 B.n134 VSUBS 0.007917f
C310 B.t5 VSUBS 0.050859f
C311 B.t4 VSUBS 0.064137f
C312 B.t3 VSUBS 0.268881f
C313 B.n135 VSUBS 0.116333f
C314 B.n136 VSUBS 0.102879f
C315 B.n137 VSUBS 0.018342f
C316 B.n138 VSUBS 0.007451f
C317 B.n139 VSUBS 0.007917f
C318 B.n140 VSUBS 0.007917f
C319 B.n141 VSUBS 0.007917f
C320 B.n142 VSUBS 0.007917f
C321 B.n143 VSUBS 0.007917f
C322 B.n144 VSUBS 0.007917f
C323 B.n145 VSUBS 0.007917f
C324 B.n146 VSUBS 0.007917f
C325 B.n147 VSUBS 0.007917f
C326 B.n148 VSUBS 0.007917f
C327 B.n149 VSUBS 0.007917f
C328 B.n150 VSUBS 0.007917f
C329 B.n151 VSUBS 0.007917f
C330 B.n152 VSUBS 0.007917f
C331 B.n153 VSUBS 0.007917f
C332 B.n154 VSUBS 0.004424f
C333 B.n155 VSUBS 0.018342f
C334 B.n156 VSUBS 0.007451f
C335 B.n157 VSUBS 0.007917f
C336 B.n158 VSUBS 0.007917f
C337 B.n159 VSUBS 0.007917f
C338 B.n160 VSUBS 0.007917f
C339 B.n161 VSUBS 0.007917f
C340 B.n162 VSUBS 0.007917f
C341 B.n163 VSUBS 0.007917f
C342 B.n164 VSUBS 0.007917f
C343 B.n165 VSUBS 0.007917f
C344 B.n166 VSUBS 0.007917f
C345 B.n167 VSUBS 0.007917f
C346 B.n168 VSUBS 0.007917f
C347 B.n169 VSUBS 0.007917f
C348 B.n170 VSUBS 0.007917f
C349 B.n171 VSUBS 0.007917f
C350 B.n172 VSUBS 0.007917f
C351 B.n173 VSUBS 0.007917f
C352 B.n174 VSUBS 0.007917f
C353 B.n175 VSUBS 0.007917f
C354 B.n176 VSUBS 0.007917f
C355 B.n177 VSUBS 0.019701f
C356 B.n178 VSUBS 0.018952f
C357 B.n179 VSUBS 0.019829f
C358 B.n180 VSUBS 0.007917f
C359 B.n181 VSUBS 0.007917f
C360 B.n182 VSUBS 0.007917f
C361 B.n183 VSUBS 0.007917f
C362 B.n184 VSUBS 0.007917f
C363 B.n185 VSUBS 0.007917f
C364 B.n186 VSUBS 0.007917f
C365 B.n187 VSUBS 0.007917f
C366 B.n188 VSUBS 0.007917f
C367 B.n189 VSUBS 0.007917f
C368 B.n190 VSUBS 0.007917f
C369 B.n191 VSUBS 0.007917f
C370 B.n192 VSUBS 0.007917f
C371 B.n193 VSUBS 0.007917f
C372 B.n194 VSUBS 0.007917f
C373 B.n195 VSUBS 0.007917f
C374 B.n196 VSUBS 0.007917f
C375 B.n197 VSUBS 0.007917f
C376 B.n198 VSUBS 0.007917f
C377 B.n199 VSUBS 0.007917f
C378 B.n200 VSUBS 0.007917f
C379 B.n201 VSUBS 0.007917f
C380 B.n202 VSUBS 0.007917f
C381 B.n203 VSUBS 0.007917f
C382 B.n204 VSUBS 0.007917f
C383 B.n205 VSUBS 0.007917f
C384 B.n206 VSUBS 0.007917f
C385 B.n207 VSUBS 0.007917f
C386 B.n208 VSUBS 0.007917f
C387 B.n209 VSUBS 0.007917f
C388 B.n210 VSUBS 0.007917f
C389 B.n211 VSUBS 0.007917f
C390 B.n212 VSUBS 0.007917f
C391 B.n213 VSUBS 0.007917f
C392 B.n214 VSUBS 0.007917f
C393 B.n215 VSUBS 0.007917f
C394 B.n216 VSUBS 0.007917f
C395 B.n217 VSUBS 0.007917f
C396 B.n218 VSUBS 0.007917f
C397 B.n219 VSUBS 0.007917f
C398 B.n220 VSUBS 0.007917f
C399 B.n221 VSUBS 0.007917f
C400 B.n222 VSUBS 0.007917f
C401 B.n223 VSUBS 0.007917f
C402 B.n224 VSUBS 0.007917f
C403 B.n225 VSUBS 0.007917f
C404 B.n226 VSUBS 0.007917f
C405 B.n227 VSUBS 0.007917f
C406 B.n228 VSUBS 0.007917f
C407 B.n229 VSUBS 0.007917f
C408 B.n230 VSUBS 0.007917f
C409 B.n231 VSUBS 0.007917f
C410 B.n232 VSUBS 0.007917f
C411 B.n233 VSUBS 0.007917f
C412 B.n234 VSUBS 0.007917f
C413 B.n235 VSUBS 0.007917f
C414 B.n236 VSUBS 0.007917f
C415 B.n237 VSUBS 0.018952f
C416 B.n238 VSUBS 0.019701f
C417 B.n239 VSUBS 0.019701f
C418 B.n240 VSUBS 0.007917f
C419 B.n241 VSUBS 0.007917f
C420 B.n242 VSUBS 0.007917f
C421 B.n243 VSUBS 0.007917f
C422 B.n244 VSUBS 0.007917f
C423 B.n245 VSUBS 0.007917f
C424 B.n246 VSUBS 0.007917f
C425 B.n247 VSUBS 0.007917f
C426 B.n248 VSUBS 0.007917f
C427 B.n249 VSUBS 0.007917f
C428 B.n250 VSUBS 0.007917f
C429 B.n251 VSUBS 0.007917f
C430 B.n252 VSUBS 0.007917f
C431 B.n253 VSUBS 0.007917f
C432 B.n254 VSUBS 0.007917f
C433 B.n255 VSUBS 0.007917f
C434 B.n256 VSUBS 0.007917f
C435 B.n257 VSUBS 0.007917f
C436 B.n258 VSUBS 0.007917f
C437 B.n259 VSUBS 0.007451f
C438 B.n260 VSUBS 0.007917f
C439 B.n261 VSUBS 0.007917f
C440 B.n262 VSUBS 0.004424f
C441 B.n263 VSUBS 0.007917f
C442 B.n264 VSUBS 0.007917f
C443 B.n265 VSUBS 0.007917f
C444 B.n266 VSUBS 0.007917f
C445 B.n267 VSUBS 0.007917f
C446 B.n268 VSUBS 0.007917f
C447 B.n269 VSUBS 0.007917f
C448 B.n270 VSUBS 0.007917f
C449 B.n271 VSUBS 0.007917f
C450 B.n272 VSUBS 0.007917f
C451 B.n273 VSUBS 0.007917f
C452 B.n274 VSUBS 0.007917f
C453 B.n275 VSUBS 0.004424f
C454 B.n276 VSUBS 0.018342f
C455 B.n277 VSUBS 0.007451f
C456 B.n278 VSUBS 0.007917f
C457 B.n279 VSUBS 0.007917f
C458 B.n280 VSUBS 0.007917f
C459 B.n281 VSUBS 0.007917f
C460 B.n282 VSUBS 0.007917f
C461 B.n283 VSUBS 0.007917f
C462 B.n284 VSUBS 0.007917f
C463 B.n285 VSUBS 0.007917f
C464 B.n286 VSUBS 0.007917f
C465 B.n287 VSUBS 0.007917f
C466 B.n288 VSUBS 0.007917f
C467 B.n289 VSUBS 0.007917f
C468 B.n290 VSUBS 0.007917f
C469 B.n291 VSUBS 0.007917f
C470 B.n292 VSUBS 0.007917f
C471 B.n293 VSUBS 0.007917f
C472 B.n294 VSUBS 0.007917f
C473 B.n295 VSUBS 0.007917f
C474 B.n296 VSUBS 0.007917f
C475 B.n297 VSUBS 0.007917f
C476 B.n298 VSUBS 0.019701f
C477 B.n299 VSUBS 0.019701f
C478 B.n300 VSUBS 0.018952f
C479 B.n301 VSUBS 0.007917f
C480 B.n302 VSUBS 0.007917f
C481 B.n303 VSUBS 0.007917f
C482 B.n304 VSUBS 0.007917f
C483 B.n305 VSUBS 0.007917f
C484 B.n306 VSUBS 0.007917f
C485 B.n307 VSUBS 0.007917f
C486 B.n308 VSUBS 0.007917f
C487 B.n309 VSUBS 0.007917f
C488 B.n310 VSUBS 0.007917f
C489 B.n311 VSUBS 0.007917f
C490 B.n312 VSUBS 0.007917f
C491 B.n313 VSUBS 0.007917f
C492 B.n314 VSUBS 0.007917f
C493 B.n315 VSUBS 0.007917f
C494 B.n316 VSUBS 0.007917f
C495 B.n317 VSUBS 0.007917f
C496 B.n318 VSUBS 0.007917f
C497 B.n319 VSUBS 0.007917f
C498 B.n320 VSUBS 0.007917f
C499 B.n321 VSUBS 0.007917f
C500 B.n322 VSUBS 0.007917f
C501 B.n323 VSUBS 0.007917f
C502 B.n324 VSUBS 0.007917f
C503 B.n325 VSUBS 0.007917f
C504 B.n326 VSUBS 0.007917f
C505 B.n327 VSUBS 0.010331f
C506 B.n328 VSUBS 0.011005f
C507 B.n329 VSUBS 0.021885f
.ends

