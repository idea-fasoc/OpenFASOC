* NGSPICE file created from diff_pair_sample_1373.ext - technology: sky130A

.subckt diff_pair_sample_1373 VTAIL VN VP B VDD2 VDD1
X0 B.t11 B.t9 B.t10 w_n2486_n3820# sky130_fd_pr__pfet_01v8 ad=5.5614 pd=29.3 as=0 ps=0 w=14.26 l=3.46
X1 B.t8 B.t6 B.t7 w_n2486_n3820# sky130_fd_pr__pfet_01v8 ad=5.5614 pd=29.3 as=0 ps=0 w=14.26 l=3.46
X2 VDD1.t1 VP.t0 VTAIL.t2 w_n2486_n3820# sky130_fd_pr__pfet_01v8 ad=5.5614 pd=29.3 as=5.5614 ps=29.3 w=14.26 l=3.46
X3 VDD2.t1 VN.t0 VTAIL.t0 w_n2486_n3820# sky130_fd_pr__pfet_01v8 ad=5.5614 pd=29.3 as=5.5614 ps=29.3 w=14.26 l=3.46
X4 B.t5 B.t3 B.t4 w_n2486_n3820# sky130_fd_pr__pfet_01v8 ad=5.5614 pd=29.3 as=0 ps=0 w=14.26 l=3.46
X5 B.t2 B.t0 B.t1 w_n2486_n3820# sky130_fd_pr__pfet_01v8 ad=5.5614 pd=29.3 as=0 ps=0 w=14.26 l=3.46
X6 VDD2.t0 VN.t1 VTAIL.t1 w_n2486_n3820# sky130_fd_pr__pfet_01v8 ad=5.5614 pd=29.3 as=5.5614 ps=29.3 w=14.26 l=3.46
X7 VDD1.t0 VP.t1 VTAIL.t3 w_n2486_n3820# sky130_fd_pr__pfet_01v8 ad=5.5614 pd=29.3 as=5.5614 ps=29.3 w=14.26 l=3.46
R0 B.n381 B.n380 585
R1 B.n379 B.n106 585
R2 B.n378 B.n377 585
R3 B.n376 B.n107 585
R4 B.n375 B.n374 585
R5 B.n373 B.n108 585
R6 B.n372 B.n371 585
R7 B.n370 B.n109 585
R8 B.n369 B.n368 585
R9 B.n367 B.n110 585
R10 B.n366 B.n365 585
R11 B.n364 B.n111 585
R12 B.n363 B.n362 585
R13 B.n361 B.n112 585
R14 B.n360 B.n359 585
R15 B.n358 B.n113 585
R16 B.n357 B.n356 585
R17 B.n355 B.n114 585
R18 B.n354 B.n353 585
R19 B.n352 B.n115 585
R20 B.n351 B.n350 585
R21 B.n349 B.n116 585
R22 B.n348 B.n347 585
R23 B.n346 B.n117 585
R24 B.n345 B.n344 585
R25 B.n343 B.n118 585
R26 B.n342 B.n341 585
R27 B.n340 B.n119 585
R28 B.n339 B.n338 585
R29 B.n337 B.n120 585
R30 B.n336 B.n335 585
R31 B.n334 B.n121 585
R32 B.n333 B.n332 585
R33 B.n331 B.n122 585
R34 B.n330 B.n329 585
R35 B.n328 B.n123 585
R36 B.n327 B.n326 585
R37 B.n325 B.n124 585
R38 B.n324 B.n323 585
R39 B.n322 B.n125 585
R40 B.n321 B.n320 585
R41 B.n319 B.n126 585
R42 B.n318 B.n317 585
R43 B.n316 B.n127 585
R44 B.n315 B.n314 585
R45 B.n313 B.n128 585
R46 B.n312 B.n311 585
R47 B.n310 B.n129 585
R48 B.n308 B.n307 585
R49 B.n306 B.n132 585
R50 B.n305 B.n304 585
R51 B.n303 B.n133 585
R52 B.n302 B.n301 585
R53 B.n300 B.n134 585
R54 B.n299 B.n298 585
R55 B.n297 B.n135 585
R56 B.n296 B.n295 585
R57 B.n294 B.n136 585
R58 B.n293 B.n292 585
R59 B.n288 B.n137 585
R60 B.n287 B.n286 585
R61 B.n285 B.n138 585
R62 B.n284 B.n283 585
R63 B.n282 B.n139 585
R64 B.n281 B.n280 585
R65 B.n279 B.n140 585
R66 B.n278 B.n277 585
R67 B.n276 B.n141 585
R68 B.n275 B.n274 585
R69 B.n273 B.n142 585
R70 B.n272 B.n271 585
R71 B.n270 B.n143 585
R72 B.n269 B.n268 585
R73 B.n267 B.n144 585
R74 B.n266 B.n265 585
R75 B.n264 B.n145 585
R76 B.n263 B.n262 585
R77 B.n261 B.n146 585
R78 B.n260 B.n259 585
R79 B.n258 B.n147 585
R80 B.n257 B.n256 585
R81 B.n255 B.n148 585
R82 B.n254 B.n253 585
R83 B.n252 B.n149 585
R84 B.n251 B.n250 585
R85 B.n249 B.n150 585
R86 B.n248 B.n247 585
R87 B.n246 B.n151 585
R88 B.n245 B.n244 585
R89 B.n243 B.n152 585
R90 B.n242 B.n241 585
R91 B.n240 B.n153 585
R92 B.n239 B.n238 585
R93 B.n237 B.n154 585
R94 B.n236 B.n235 585
R95 B.n234 B.n155 585
R96 B.n233 B.n232 585
R97 B.n231 B.n156 585
R98 B.n230 B.n229 585
R99 B.n228 B.n157 585
R100 B.n227 B.n226 585
R101 B.n225 B.n158 585
R102 B.n224 B.n223 585
R103 B.n222 B.n159 585
R104 B.n221 B.n220 585
R105 B.n219 B.n160 585
R106 B.n382 B.n105 585
R107 B.n384 B.n383 585
R108 B.n385 B.n104 585
R109 B.n387 B.n386 585
R110 B.n388 B.n103 585
R111 B.n390 B.n389 585
R112 B.n391 B.n102 585
R113 B.n393 B.n392 585
R114 B.n394 B.n101 585
R115 B.n396 B.n395 585
R116 B.n397 B.n100 585
R117 B.n399 B.n398 585
R118 B.n400 B.n99 585
R119 B.n402 B.n401 585
R120 B.n403 B.n98 585
R121 B.n405 B.n404 585
R122 B.n406 B.n97 585
R123 B.n408 B.n407 585
R124 B.n409 B.n96 585
R125 B.n411 B.n410 585
R126 B.n412 B.n95 585
R127 B.n414 B.n413 585
R128 B.n415 B.n94 585
R129 B.n417 B.n416 585
R130 B.n418 B.n93 585
R131 B.n420 B.n419 585
R132 B.n421 B.n92 585
R133 B.n423 B.n422 585
R134 B.n424 B.n91 585
R135 B.n426 B.n425 585
R136 B.n427 B.n90 585
R137 B.n429 B.n428 585
R138 B.n430 B.n89 585
R139 B.n432 B.n431 585
R140 B.n433 B.n88 585
R141 B.n435 B.n434 585
R142 B.n436 B.n87 585
R143 B.n438 B.n437 585
R144 B.n439 B.n86 585
R145 B.n441 B.n440 585
R146 B.n442 B.n85 585
R147 B.n444 B.n443 585
R148 B.n445 B.n84 585
R149 B.n447 B.n446 585
R150 B.n448 B.n83 585
R151 B.n450 B.n449 585
R152 B.n451 B.n82 585
R153 B.n453 B.n452 585
R154 B.n454 B.n81 585
R155 B.n456 B.n455 585
R156 B.n457 B.n80 585
R157 B.n459 B.n458 585
R158 B.n460 B.n79 585
R159 B.n462 B.n461 585
R160 B.n463 B.n78 585
R161 B.n465 B.n464 585
R162 B.n466 B.n77 585
R163 B.n468 B.n467 585
R164 B.n469 B.n76 585
R165 B.n471 B.n470 585
R166 B.n472 B.n75 585
R167 B.n474 B.n473 585
R168 B.n634 B.n17 585
R169 B.n633 B.n632 585
R170 B.n631 B.n18 585
R171 B.n630 B.n629 585
R172 B.n628 B.n19 585
R173 B.n627 B.n626 585
R174 B.n625 B.n20 585
R175 B.n624 B.n623 585
R176 B.n622 B.n21 585
R177 B.n621 B.n620 585
R178 B.n619 B.n22 585
R179 B.n618 B.n617 585
R180 B.n616 B.n23 585
R181 B.n615 B.n614 585
R182 B.n613 B.n24 585
R183 B.n612 B.n611 585
R184 B.n610 B.n25 585
R185 B.n609 B.n608 585
R186 B.n607 B.n26 585
R187 B.n606 B.n605 585
R188 B.n604 B.n27 585
R189 B.n603 B.n602 585
R190 B.n601 B.n28 585
R191 B.n600 B.n599 585
R192 B.n598 B.n29 585
R193 B.n597 B.n596 585
R194 B.n595 B.n30 585
R195 B.n594 B.n593 585
R196 B.n592 B.n31 585
R197 B.n591 B.n590 585
R198 B.n589 B.n32 585
R199 B.n588 B.n587 585
R200 B.n586 B.n33 585
R201 B.n585 B.n584 585
R202 B.n583 B.n34 585
R203 B.n582 B.n581 585
R204 B.n580 B.n35 585
R205 B.n579 B.n578 585
R206 B.n577 B.n36 585
R207 B.n576 B.n575 585
R208 B.n574 B.n37 585
R209 B.n573 B.n572 585
R210 B.n571 B.n38 585
R211 B.n570 B.n569 585
R212 B.n568 B.n39 585
R213 B.n567 B.n566 585
R214 B.n565 B.n40 585
R215 B.n564 B.n563 585
R216 B.n561 B.n41 585
R217 B.n560 B.n559 585
R218 B.n558 B.n44 585
R219 B.n557 B.n556 585
R220 B.n555 B.n45 585
R221 B.n554 B.n553 585
R222 B.n552 B.n46 585
R223 B.n551 B.n550 585
R224 B.n549 B.n47 585
R225 B.n548 B.n547 585
R226 B.n546 B.n545 585
R227 B.n544 B.n51 585
R228 B.n543 B.n542 585
R229 B.n541 B.n52 585
R230 B.n540 B.n539 585
R231 B.n538 B.n53 585
R232 B.n537 B.n536 585
R233 B.n535 B.n54 585
R234 B.n534 B.n533 585
R235 B.n532 B.n55 585
R236 B.n531 B.n530 585
R237 B.n529 B.n56 585
R238 B.n528 B.n527 585
R239 B.n526 B.n57 585
R240 B.n525 B.n524 585
R241 B.n523 B.n58 585
R242 B.n522 B.n521 585
R243 B.n520 B.n59 585
R244 B.n519 B.n518 585
R245 B.n517 B.n60 585
R246 B.n516 B.n515 585
R247 B.n514 B.n61 585
R248 B.n513 B.n512 585
R249 B.n511 B.n62 585
R250 B.n510 B.n509 585
R251 B.n508 B.n63 585
R252 B.n507 B.n506 585
R253 B.n505 B.n64 585
R254 B.n504 B.n503 585
R255 B.n502 B.n65 585
R256 B.n501 B.n500 585
R257 B.n499 B.n66 585
R258 B.n498 B.n497 585
R259 B.n496 B.n67 585
R260 B.n495 B.n494 585
R261 B.n493 B.n68 585
R262 B.n492 B.n491 585
R263 B.n490 B.n69 585
R264 B.n489 B.n488 585
R265 B.n487 B.n70 585
R266 B.n486 B.n485 585
R267 B.n484 B.n71 585
R268 B.n483 B.n482 585
R269 B.n481 B.n72 585
R270 B.n480 B.n479 585
R271 B.n478 B.n73 585
R272 B.n477 B.n476 585
R273 B.n475 B.n74 585
R274 B.n636 B.n635 585
R275 B.n637 B.n16 585
R276 B.n639 B.n638 585
R277 B.n640 B.n15 585
R278 B.n642 B.n641 585
R279 B.n643 B.n14 585
R280 B.n645 B.n644 585
R281 B.n646 B.n13 585
R282 B.n648 B.n647 585
R283 B.n649 B.n12 585
R284 B.n651 B.n650 585
R285 B.n652 B.n11 585
R286 B.n654 B.n653 585
R287 B.n655 B.n10 585
R288 B.n657 B.n656 585
R289 B.n658 B.n9 585
R290 B.n660 B.n659 585
R291 B.n661 B.n8 585
R292 B.n663 B.n662 585
R293 B.n664 B.n7 585
R294 B.n666 B.n665 585
R295 B.n667 B.n6 585
R296 B.n669 B.n668 585
R297 B.n670 B.n5 585
R298 B.n672 B.n671 585
R299 B.n673 B.n4 585
R300 B.n675 B.n674 585
R301 B.n676 B.n3 585
R302 B.n678 B.n677 585
R303 B.n679 B.n0 585
R304 B.n2 B.n1 585
R305 B.n176 B.n175 585
R306 B.n177 B.n174 585
R307 B.n179 B.n178 585
R308 B.n180 B.n173 585
R309 B.n182 B.n181 585
R310 B.n183 B.n172 585
R311 B.n185 B.n184 585
R312 B.n186 B.n171 585
R313 B.n188 B.n187 585
R314 B.n189 B.n170 585
R315 B.n191 B.n190 585
R316 B.n192 B.n169 585
R317 B.n194 B.n193 585
R318 B.n195 B.n168 585
R319 B.n197 B.n196 585
R320 B.n198 B.n167 585
R321 B.n200 B.n199 585
R322 B.n201 B.n166 585
R323 B.n203 B.n202 585
R324 B.n204 B.n165 585
R325 B.n206 B.n205 585
R326 B.n207 B.n164 585
R327 B.n209 B.n208 585
R328 B.n210 B.n163 585
R329 B.n212 B.n211 585
R330 B.n213 B.n162 585
R331 B.n215 B.n214 585
R332 B.n216 B.n161 585
R333 B.n218 B.n217 585
R334 B.n219 B.n218 492.5
R335 B.n380 B.n105 492.5
R336 B.n475 B.n474 492.5
R337 B.n636 B.n17 492.5
R338 B.n130 B.t1 490.041
R339 B.n48 B.t11 490.041
R340 B.n289 B.t4 490.041
R341 B.n42 B.t8 490.041
R342 B.n131 B.t2 416.538
R343 B.n49 B.t10 416.538
R344 B.n290 B.t5 416.538
R345 B.n43 B.t7 416.538
R346 B.n289 B.t3 308.384
R347 B.n130 B.t0 308.384
R348 B.n48 B.t9 308.384
R349 B.n42 B.t6 308.384
R350 B.n681 B.n680 256.663
R351 B.n680 B.n679 235.042
R352 B.n680 B.n2 235.042
R353 B.n220 B.n219 163.367
R354 B.n220 B.n159 163.367
R355 B.n224 B.n159 163.367
R356 B.n225 B.n224 163.367
R357 B.n226 B.n225 163.367
R358 B.n226 B.n157 163.367
R359 B.n230 B.n157 163.367
R360 B.n231 B.n230 163.367
R361 B.n232 B.n231 163.367
R362 B.n232 B.n155 163.367
R363 B.n236 B.n155 163.367
R364 B.n237 B.n236 163.367
R365 B.n238 B.n237 163.367
R366 B.n238 B.n153 163.367
R367 B.n242 B.n153 163.367
R368 B.n243 B.n242 163.367
R369 B.n244 B.n243 163.367
R370 B.n244 B.n151 163.367
R371 B.n248 B.n151 163.367
R372 B.n249 B.n248 163.367
R373 B.n250 B.n249 163.367
R374 B.n250 B.n149 163.367
R375 B.n254 B.n149 163.367
R376 B.n255 B.n254 163.367
R377 B.n256 B.n255 163.367
R378 B.n256 B.n147 163.367
R379 B.n260 B.n147 163.367
R380 B.n261 B.n260 163.367
R381 B.n262 B.n261 163.367
R382 B.n262 B.n145 163.367
R383 B.n266 B.n145 163.367
R384 B.n267 B.n266 163.367
R385 B.n268 B.n267 163.367
R386 B.n268 B.n143 163.367
R387 B.n272 B.n143 163.367
R388 B.n273 B.n272 163.367
R389 B.n274 B.n273 163.367
R390 B.n274 B.n141 163.367
R391 B.n278 B.n141 163.367
R392 B.n279 B.n278 163.367
R393 B.n280 B.n279 163.367
R394 B.n280 B.n139 163.367
R395 B.n284 B.n139 163.367
R396 B.n285 B.n284 163.367
R397 B.n286 B.n285 163.367
R398 B.n286 B.n137 163.367
R399 B.n293 B.n137 163.367
R400 B.n294 B.n293 163.367
R401 B.n295 B.n294 163.367
R402 B.n295 B.n135 163.367
R403 B.n299 B.n135 163.367
R404 B.n300 B.n299 163.367
R405 B.n301 B.n300 163.367
R406 B.n301 B.n133 163.367
R407 B.n305 B.n133 163.367
R408 B.n306 B.n305 163.367
R409 B.n307 B.n306 163.367
R410 B.n307 B.n129 163.367
R411 B.n312 B.n129 163.367
R412 B.n313 B.n312 163.367
R413 B.n314 B.n313 163.367
R414 B.n314 B.n127 163.367
R415 B.n318 B.n127 163.367
R416 B.n319 B.n318 163.367
R417 B.n320 B.n319 163.367
R418 B.n320 B.n125 163.367
R419 B.n324 B.n125 163.367
R420 B.n325 B.n324 163.367
R421 B.n326 B.n325 163.367
R422 B.n326 B.n123 163.367
R423 B.n330 B.n123 163.367
R424 B.n331 B.n330 163.367
R425 B.n332 B.n331 163.367
R426 B.n332 B.n121 163.367
R427 B.n336 B.n121 163.367
R428 B.n337 B.n336 163.367
R429 B.n338 B.n337 163.367
R430 B.n338 B.n119 163.367
R431 B.n342 B.n119 163.367
R432 B.n343 B.n342 163.367
R433 B.n344 B.n343 163.367
R434 B.n344 B.n117 163.367
R435 B.n348 B.n117 163.367
R436 B.n349 B.n348 163.367
R437 B.n350 B.n349 163.367
R438 B.n350 B.n115 163.367
R439 B.n354 B.n115 163.367
R440 B.n355 B.n354 163.367
R441 B.n356 B.n355 163.367
R442 B.n356 B.n113 163.367
R443 B.n360 B.n113 163.367
R444 B.n361 B.n360 163.367
R445 B.n362 B.n361 163.367
R446 B.n362 B.n111 163.367
R447 B.n366 B.n111 163.367
R448 B.n367 B.n366 163.367
R449 B.n368 B.n367 163.367
R450 B.n368 B.n109 163.367
R451 B.n372 B.n109 163.367
R452 B.n373 B.n372 163.367
R453 B.n374 B.n373 163.367
R454 B.n374 B.n107 163.367
R455 B.n378 B.n107 163.367
R456 B.n379 B.n378 163.367
R457 B.n380 B.n379 163.367
R458 B.n474 B.n75 163.367
R459 B.n470 B.n75 163.367
R460 B.n470 B.n469 163.367
R461 B.n469 B.n468 163.367
R462 B.n468 B.n77 163.367
R463 B.n464 B.n77 163.367
R464 B.n464 B.n463 163.367
R465 B.n463 B.n462 163.367
R466 B.n462 B.n79 163.367
R467 B.n458 B.n79 163.367
R468 B.n458 B.n457 163.367
R469 B.n457 B.n456 163.367
R470 B.n456 B.n81 163.367
R471 B.n452 B.n81 163.367
R472 B.n452 B.n451 163.367
R473 B.n451 B.n450 163.367
R474 B.n450 B.n83 163.367
R475 B.n446 B.n83 163.367
R476 B.n446 B.n445 163.367
R477 B.n445 B.n444 163.367
R478 B.n444 B.n85 163.367
R479 B.n440 B.n85 163.367
R480 B.n440 B.n439 163.367
R481 B.n439 B.n438 163.367
R482 B.n438 B.n87 163.367
R483 B.n434 B.n87 163.367
R484 B.n434 B.n433 163.367
R485 B.n433 B.n432 163.367
R486 B.n432 B.n89 163.367
R487 B.n428 B.n89 163.367
R488 B.n428 B.n427 163.367
R489 B.n427 B.n426 163.367
R490 B.n426 B.n91 163.367
R491 B.n422 B.n91 163.367
R492 B.n422 B.n421 163.367
R493 B.n421 B.n420 163.367
R494 B.n420 B.n93 163.367
R495 B.n416 B.n93 163.367
R496 B.n416 B.n415 163.367
R497 B.n415 B.n414 163.367
R498 B.n414 B.n95 163.367
R499 B.n410 B.n95 163.367
R500 B.n410 B.n409 163.367
R501 B.n409 B.n408 163.367
R502 B.n408 B.n97 163.367
R503 B.n404 B.n97 163.367
R504 B.n404 B.n403 163.367
R505 B.n403 B.n402 163.367
R506 B.n402 B.n99 163.367
R507 B.n398 B.n99 163.367
R508 B.n398 B.n397 163.367
R509 B.n397 B.n396 163.367
R510 B.n396 B.n101 163.367
R511 B.n392 B.n101 163.367
R512 B.n392 B.n391 163.367
R513 B.n391 B.n390 163.367
R514 B.n390 B.n103 163.367
R515 B.n386 B.n103 163.367
R516 B.n386 B.n385 163.367
R517 B.n385 B.n384 163.367
R518 B.n384 B.n105 163.367
R519 B.n632 B.n17 163.367
R520 B.n632 B.n631 163.367
R521 B.n631 B.n630 163.367
R522 B.n630 B.n19 163.367
R523 B.n626 B.n19 163.367
R524 B.n626 B.n625 163.367
R525 B.n625 B.n624 163.367
R526 B.n624 B.n21 163.367
R527 B.n620 B.n21 163.367
R528 B.n620 B.n619 163.367
R529 B.n619 B.n618 163.367
R530 B.n618 B.n23 163.367
R531 B.n614 B.n23 163.367
R532 B.n614 B.n613 163.367
R533 B.n613 B.n612 163.367
R534 B.n612 B.n25 163.367
R535 B.n608 B.n25 163.367
R536 B.n608 B.n607 163.367
R537 B.n607 B.n606 163.367
R538 B.n606 B.n27 163.367
R539 B.n602 B.n27 163.367
R540 B.n602 B.n601 163.367
R541 B.n601 B.n600 163.367
R542 B.n600 B.n29 163.367
R543 B.n596 B.n29 163.367
R544 B.n596 B.n595 163.367
R545 B.n595 B.n594 163.367
R546 B.n594 B.n31 163.367
R547 B.n590 B.n31 163.367
R548 B.n590 B.n589 163.367
R549 B.n589 B.n588 163.367
R550 B.n588 B.n33 163.367
R551 B.n584 B.n33 163.367
R552 B.n584 B.n583 163.367
R553 B.n583 B.n582 163.367
R554 B.n582 B.n35 163.367
R555 B.n578 B.n35 163.367
R556 B.n578 B.n577 163.367
R557 B.n577 B.n576 163.367
R558 B.n576 B.n37 163.367
R559 B.n572 B.n37 163.367
R560 B.n572 B.n571 163.367
R561 B.n571 B.n570 163.367
R562 B.n570 B.n39 163.367
R563 B.n566 B.n39 163.367
R564 B.n566 B.n565 163.367
R565 B.n565 B.n564 163.367
R566 B.n564 B.n41 163.367
R567 B.n559 B.n41 163.367
R568 B.n559 B.n558 163.367
R569 B.n558 B.n557 163.367
R570 B.n557 B.n45 163.367
R571 B.n553 B.n45 163.367
R572 B.n553 B.n552 163.367
R573 B.n552 B.n551 163.367
R574 B.n551 B.n47 163.367
R575 B.n547 B.n47 163.367
R576 B.n547 B.n546 163.367
R577 B.n546 B.n51 163.367
R578 B.n542 B.n51 163.367
R579 B.n542 B.n541 163.367
R580 B.n541 B.n540 163.367
R581 B.n540 B.n53 163.367
R582 B.n536 B.n53 163.367
R583 B.n536 B.n535 163.367
R584 B.n535 B.n534 163.367
R585 B.n534 B.n55 163.367
R586 B.n530 B.n55 163.367
R587 B.n530 B.n529 163.367
R588 B.n529 B.n528 163.367
R589 B.n528 B.n57 163.367
R590 B.n524 B.n57 163.367
R591 B.n524 B.n523 163.367
R592 B.n523 B.n522 163.367
R593 B.n522 B.n59 163.367
R594 B.n518 B.n59 163.367
R595 B.n518 B.n517 163.367
R596 B.n517 B.n516 163.367
R597 B.n516 B.n61 163.367
R598 B.n512 B.n61 163.367
R599 B.n512 B.n511 163.367
R600 B.n511 B.n510 163.367
R601 B.n510 B.n63 163.367
R602 B.n506 B.n63 163.367
R603 B.n506 B.n505 163.367
R604 B.n505 B.n504 163.367
R605 B.n504 B.n65 163.367
R606 B.n500 B.n65 163.367
R607 B.n500 B.n499 163.367
R608 B.n499 B.n498 163.367
R609 B.n498 B.n67 163.367
R610 B.n494 B.n67 163.367
R611 B.n494 B.n493 163.367
R612 B.n493 B.n492 163.367
R613 B.n492 B.n69 163.367
R614 B.n488 B.n69 163.367
R615 B.n488 B.n487 163.367
R616 B.n487 B.n486 163.367
R617 B.n486 B.n71 163.367
R618 B.n482 B.n71 163.367
R619 B.n482 B.n481 163.367
R620 B.n481 B.n480 163.367
R621 B.n480 B.n73 163.367
R622 B.n476 B.n73 163.367
R623 B.n476 B.n475 163.367
R624 B.n637 B.n636 163.367
R625 B.n638 B.n637 163.367
R626 B.n638 B.n15 163.367
R627 B.n642 B.n15 163.367
R628 B.n643 B.n642 163.367
R629 B.n644 B.n643 163.367
R630 B.n644 B.n13 163.367
R631 B.n648 B.n13 163.367
R632 B.n649 B.n648 163.367
R633 B.n650 B.n649 163.367
R634 B.n650 B.n11 163.367
R635 B.n654 B.n11 163.367
R636 B.n655 B.n654 163.367
R637 B.n656 B.n655 163.367
R638 B.n656 B.n9 163.367
R639 B.n660 B.n9 163.367
R640 B.n661 B.n660 163.367
R641 B.n662 B.n661 163.367
R642 B.n662 B.n7 163.367
R643 B.n666 B.n7 163.367
R644 B.n667 B.n666 163.367
R645 B.n668 B.n667 163.367
R646 B.n668 B.n5 163.367
R647 B.n672 B.n5 163.367
R648 B.n673 B.n672 163.367
R649 B.n674 B.n673 163.367
R650 B.n674 B.n3 163.367
R651 B.n678 B.n3 163.367
R652 B.n679 B.n678 163.367
R653 B.n176 B.n2 163.367
R654 B.n177 B.n176 163.367
R655 B.n178 B.n177 163.367
R656 B.n178 B.n173 163.367
R657 B.n182 B.n173 163.367
R658 B.n183 B.n182 163.367
R659 B.n184 B.n183 163.367
R660 B.n184 B.n171 163.367
R661 B.n188 B.n171 163.367
R662 B.n189 B.n188 163.367
R663 B.n190 B.n189 163.367
R664 B.n190 B.n169 163.367
R665 B.n194 B.n169 163.367
R666 B.n195 B.n194 163.367
R667 B.n196 B.n195 163.367
R668 B.n196 B.n167 163.367
R669 B.n200 B.n167 163.367
R670 B.n201 B.n200 163.367
R671 B.n202 B.n201 163.367
R672 B.n202 B.n165 163.367
R673 B.n206 B.n165 163.367
R674 B.n207 B.n206 163.367
R675 B.n208 B.n207 163.367
R676 B.n208 B.n163 163.367
R677 B.n212 B.n163 163.367
R678 B.n213 B.n212 163.367
R679 B.n214 B.n213 163.367
R680 B.n214 B.n161 163.367
R681 B.n218 B.n161 163.367
R682 B.n290 B.n289 73.5035
R683 B.n131 B.n130 73.5035
R684 B.n49 B.n48 73.5035
R685 B.n43 B.n42 73.5035
R686 B.n291 B.n290 59.5399
R687 B.n309 B.n131 59.5399
R688 B.n50 B.n49 59.5399
R689 B.n562 B.n43 59.5399
R690 B.n635 B.n634 32.0005
R691 B.n473 B.n74 32.0005
R692 B.n382 B.n381 32.0005
R693 B.n217 B.n160 32.0005
R694 B B.n681 18.0485
R695 B.n635 B.n16 10.6151
R696 B.n639 B.n16 10.6151
R697 B.n640 B.n639 10.6151
R698 B.n641 B.n640 10.6151
R699 B.n641 B.n14 10.6151
R700 B.n645 B.n14 10.6151
R701 B.n646 B.n645 10.6151
R702 B.n647 B.n646 10.6151
R703 B.n647 B.n12 10.6151
R704 B.n651 B.n12 10.6151
R705 B.n652 B.n651 10.6151
R706 B.n653 B.n652 10.6151
R707 B.n653 B.n10 10.6151
R708 B.n657 B.n10 10.6151
R709 B.n658 B.n657 10.6151
R710 B.n659 B.n658 10.6151
R711 B.n659 B.n8 10.6151
R712 B.n663 B.n8 10.6151
R713 B.n664 B.n663 10.6151
R714 B.n665 B.n664 10.6151
R715 B.n665 B.n6 10.6151
R716 B.n669 B.n6 10.6151
R717 B.n670 B.n669 10.6151
R718 B.n671 B.n670 10.6151
R719 B.n671 B.n4 10.6151
R720 B.n675 B.n4 10.6151
R721 B.n676 B.n675 10.6151
R722 B.n677 B.n676 10.6151
R723 B.n677 B.n0 10.6151
R724 B.n634 B.n633 10.6151
R725 B.n633 B.n18 10.6151
R726 B.n629 B.n18 10.6151
R727 B.n629 B.n628 10.6151
R728 B.n628 B.n627 10.6151
R729 B.n627 B.n20 10.6151
R730 B.n623 B.n20 10.6151
R731 B.n623 B.n622 10.6151
R732 B.n622 B.n621 10.6151
R733 B.n621 B.n22 10.6151
R734 B.n617 B.n22 10.6151
R735 B.n617 B.n616 10.6151
R736 B.n616 B.n615 10.6151
R737 B.n615 B.n24 10.6151
R738 B.n611 B.n24 10.6151
R739 B.n611 B.n610 10.6151
R740 B.n610 B.n609 10.6151
R741 B.n609 B.n26 10.6151
R742 B.n605 B.n26 10.6151
R743 B.n605 B.n604 10.6151
R744 B.n604 B.n603 10.6151
R745 B.n603 B.n28 10.6151
R746 B.n599 B.n28 10.6151
R747 B.n599 B.n598 10.6151
R748 B.n598 B.n597 10.6151
R749 B.n597 B.n30 10.6151
R750 B.n593 B.n30 10.6151
R751 B.n593 B.n592 10.6151
R752 B.n592 B.n591 10.6151
R753 B.n591 B.n32 10.6151
R754 B.n587 B.n32 10.6151
R755 B.n587 B.n586 10.6151
R756 B.n586 B.n585 10.6151
R757 B.n585 B.n34 10.6151
R758 B.n581 B.n34 10.6151
R759 B.n581 B.n580 10.6151
R760 B.n580 B.n579 10.6151
R761 B.n579 B.n36 10.6151
R762 B.n575 B.n36 10.6151
R763 B.n575 B.n574 10.6151
R764 B.n574 B.n573 10.6151
R765 B.n573 B.n38 10.6151
R766 B.n569 B.n38 10.6151
R767 B.n569 B.n568 10.6151
R768 B.n568 B.n567 10.6151
R769 B.n567 B.n40 10.6151
R770 B.n563 B.n40 10.6151
R771 B.n561 B.n560 10.6151
R772 B.n560 B.n44 10.6151
R773 B.n556 B.n44 10.6151
R774 B.n556 B.n555 10.6151
R775 B.n555 B.n554 10.6151
R776 B.n554 B.n46 10.6151
R777 B.n550 B.n46 10.6151
R778 B.n550 B.n549 10.6151
R779 B.n549 B.n548 10.6151
R780 B.n545 B.n544 10.6151
R781 B.n544 B.n543 10.6151
R782 B.n543 B.n52 10.6151
R783 B.n539 B.n52 10.6151
R784 B.n539 B.n538 10.6151
R785 B.n538 B.n537 10.6151
R786 B.n537 B.n54 10.6151
R787 B.n533 B.n54 10.6151
R788 B.n533 B.n532 10.6151
R789 B.n532 B.n531 10.6151
R790 B.n531 B.n56 10.6151
R791 B.n527 B.n56 10.6151
R792 B.n527 B.n526 10.6151
R793 B.n526 B.n525 10.6151
R794 B.n525 B.n58 10.6151
R795 B.n521 B.n58 10.6151
R796 B.n521 B.n520 10.6151
R797 B.n520 B.n519 10.6151
R798 B.n519 B.n60 10.6151
R799 B.n515 B.n60 10.6151
R800 B.n515 B.n514 10.6151
R801 B.n514 B.n513 10.6151
R802 B.n513 B.n62 10.6151
R803 B.n509 B.n62 10.6151
R804 B.n509 B.n508 10.6151
R805 B.n508 B.n507 10.6151
R806 B.n507 B.n64 10.6151
R807 B.n503 B.n64 10.6151
R808 B.n503 B.n502 10.6151
R809 B.n502 B.n501 10.6151
R810 B.n501 B.n66 10.6151
R811 B.n497 B.n66 10.6151
R812 B.n497 B.n496 10.6151
R813 B.n496 B.n495 10.6151
R814 B.n495 B.n68 10.6151
R815 B.n491 B.n68 10.6151
R816 B.n491 B.n490 10.6151
R817 B.n490 B.n489 10.6151
R818 B.n489 B.n70 10.6151
R819 B.n485 B.n70 10.6151
R820 B.n485 B.n484 10.6151
R821 B.n484 B.n483 10.6151
R822 B.n483 B.n72 10.6151
R823 B.n479 B.n72 10.6151
R824 B.n479 B.n478 10.6151
R825 B.n478 B.n477 10.6151
R826 B.n477 B.n74 10.6151
R827 B.n473 B.n472 10.6151
R828 B.n472 B.n471 10.6151
R829 B.n471 B.n76 10.6151
R830 B.n467 B.n76 10.6151
R831 B.n467 B.n466 10.6151
R832 B.n466 B.n465 10.6151
R833 B.n465 B.n78 10.6151
R834 B.n461 B.n78 10.6151
R835 B.n461 B.n460 10.6151
R836 B.n460 B.n459 10.6151
R837 B.n459 B.n80 10.6151
R838 B.n455 B.n80 10.6151
R839 B.n455 B.n454 10.6151
R840 B.n454 B.n453 10.6151
R841 B.n453 B.n82 10.6151
R842 B.n449 B.n82 10.6151
R843 B.n449 B.n448 10.6151
R844 B.n448 B.n447 10.6151
R845 B.n447 B.n84 10.6151
R846 B.n443 B.n84 10.6151
R847 B.n443 B.n442 10.6151
R848 B.n442 B.n441 10.6151
R849 B.n441 B.n86 10.6151
R850 B.n437 B.n86 10.6151
R851 B.n437 B.n436 10.6151
R852 B.n436 B.n435 10.6151
R853 B.n435 B.n88 10.6151
R854 B.n431 B.n88 10.6151
R855 B.n431 B.n430 10.6151
R856 B.n430 B.n429 10.6151
R857 B.n429 B.n90 10.6151
R858 B.n425 B.n90 10.6151
R859 B.n425 B.n424 10.6151
R860 B.n424 B.n423 10.6151
R861 B.n423 B.n92 10.6151
R862 B.n419 B.n92 10.6151
R863 B.n419 B.n418 10.6151
R864 B.n418 B.n417 10.6151
R865 B.n417 B.n94 10.6151
R866 B.n413 B.n94 10.6151
R867 B.n413 B.n412 10.6151
R868 B.n412 B.n411 10.6151
R869 B.n411 B.n96 10.6151
R870 B.n407 B.n96 10.6151
R871 B.n407 B.n406 10.6151
R872 B.n406 B.n405 10.6151
R873 B.n405 B.n98 10.6151
R874 B.n401 B.n98 10.6151
R875 B.n401 B.n400 10.6151
R876 B.n400 B.n399 10.6151
R877 B.n399 B.n100 10.6151
R878 B.n395 B.n100 10.6151
R879 B.n395 B.n394 10.6151
R880 B.n394 B.n393 10.6151
R881 B.n393 B.n102 10.6151
R882 B.n389 B.n102 10.6151
R883 B.n389 B.n388 10.6151
R884 B.n388 B.n387 10.6151
R885 B.n387 B.n104 10.6151
R886 B.n383 B.n104 10.6151
R887 B.n383 B.n382 10.6151
R888 B.n175 B.n1 10.6151
R889 B.n175 B.n174 10.6151
R890 B.n179 B.n174 10.6151
R891 B.n180 B.n179 10.6151
R892 B.n181 B.n180 10.6151
R893 B.n181 B.n172 10.6151
R894 B.n185 B.n172 10.6151
R895 B.n186 B.n185 10.6151
R896 B.n187 B.n186 10.6151
R897 B.n187 B.n170 10.6151
R898 B.n191 B.n170 10.6151
R899 B.n192 B.n191 10.6151
R900 B.n193 B.n192 10.6151
R901 B.n193 B.n168 10.6151
R902 B.n197 B.n168 10.6151
R903 B.n198 B.n197 10.6151
R904 B.n199 B.n198 10.6151
R905 B.n199 B.n166 10.6151
R906 B.n203 B.n166 10.6151
R907 B.n204 B.n203 10.6151
R908 B.n205 B.n204 10.6151
R909 B.n205 B.n164 10.6151
R910 B.n209 B.n164 10.6151
R911 B.n210 B.n209 10.6151
R912 B.n211 B.n210 10.6151
R913 B.n211 B.n162 10.6151
R914 B.n215 B.n162 10.6151
R915 B.n216 B.n215 10.6151
R916 B.n217 B.n216 10.6151
R917 B.n221 B.n160 10.6151
R918 B.n222 B.n221 10.6151
R919 B.n223 B.n222 10.6151
R920 B.n223 B.n158 10.6151
R921 B.n227 B.n158 10.6151
R922 B.n228 B.n227 10.6151
R923 B.n229 B.n228 10.6151
R924 B.n229 B.n156 10.6151
R925 B.n233 B.n156 10.6151
R926 B.n234 B.n233 10.6151
R927 B.n235 B.n234 10.6151
R928 B.n235 B.n154 10.6151
R929 B.n239 B.n154 10.6151
R930 B.n240 B.n239 10.6151
R931 B.n241 B.n240 10.6151
R932 B.n241 B.n152 10.6151
R933 B.n245 B.n152 10.6151
R934 B.n246 B.n245 10.6151
R935 B.n247 B.n246 10.6151
R936 B.n247 B.n150 10.6151
R937 B.n251 B.n150 10.6151
R938 B.n252 B.n251 10.6151
R939 B.n253 B.n252 10.6151
R940 B.n253 B.n148 10.6151
R941 B.n257 B.n148 10.6151
R942 B.n258 B.n257 10.6151
R943 B.n259 B.n258 10.6151
R944 B.n259 B.n146 10.6151
R945 B.n263 B.n146 10.6151
R946 B.n264 B.n263 10.6151
R947 B.n265 B.n264 10.6151
R948 B.n265 B.n144 10.6151
R949 B.n269 B.n144 10.6151
R950 B.n270 B.n269 10.6151
R951 B.n271 B.n270 10.6151
R952 B.n271 B.n142 10.6151
R953 B.n275 B.n142 10.6151
R954 B.n276 B.n275 10.6151
R955 B.n277 B.n276 10.6151
R956 B.n277 B.n140 10.6151
R957 B.n281 B.n140 10.6151
R958 B.n282 B.n281 10.6151
R959 B.n283 B.n282 10.6151
R960 B.n283 B.n138 10.6151
R961 B.n287 B.n138 10.6151
R962 B.n288 B.n287 10.6151
R963 B.n292 B.n288 10.6151
R964 B.n296 B.n136 10.6151
R965 B.n297 B.n296 10.6151
R966 B.n298 B.n297 10.6151
R967 B.n298 B.n134 10.6151
R968 B.n302 B.n134 10.6151
R969 B.n303 B.n302 10.6151
R970 B.n304 B.n303 10.6151
R971 B.n304 B.n132 10.6151
R972 B.n308 B.n132 10.6151
R973 B.n311 B.n310 10.6151
R974 B.n311 B.n128 10.6151
R975 B.n315 B.n128 10.6151
R976 B.n316 B.n315 10.6151
R977 B.n317 B.n316 10.6151
R978 B.n317 B.n126 10.6151
R979 B.n321 B.n126 10.6151
R980 B.n322 B.n321 10.6151
R981 B.n323 B.n322 10.6151
R982 B.n323 B.n124 10.6151
R983 B.n327 B.n124 10.6151
R984 B.n328 B.n327 10.6151
R985 B.n329 B.n328 10.6151
R986 B.n329 B.n122 10.6151
R987 B.n333 B.n122 10.6151
R988 B.n334 B.n333 10.6151
R989 B.n335 B.n334 10.6151
R990 B.n335 B.n120 10.6151
R991 B.n339 B.n120 10.6151
R992 B.n340 B.n339 10.6151
R993 B.n341 B.n340 10.6151
R994 B.n341 B.n118 10.6151
R995 B.n345 B.n118 10.6151
R996 B.n346 B.n345 10.6151
R997 B.n347 B.n346 10.6151
R998 B.n347 B.n116 10.6151
R999 B.n351 B.n116 10.6151
R1000 B.n352 B.n351 10.6151
R1001 B.n353 B.n352 10.6151
R1002 B.n353 B.n114 10.6151
R1003 B.n357 B.n114 10.6151
R1004 B.n358 B.n357 10.6151
R1005 B.n359 B.n358 10.6151
R1006 B.n359 B.n112 10.6151
R1007 B.n363 B.n112 10.6151
R1008 B.n364 B.n363 10.6151
R1009 B.n365 B.n364 10.6151
R1010 B.n365 B.n110 10.6151
R1011 B.n369 B.n110 10.6151
R1012 B.n370 B.n369 10.6151
R1013 B.n371 B.n370 10.6151
R1014 B.n371 B.n108 10.6151
R1015 B.n375 B.n108 10.6151
R1016 B.n376 B.n375 10.6151
R1017 B.n377 B.n376 10.6151
R1018 B.n377 B.n106 10.6151
R1019 B.n381 B.n106 10.6151
R1020 B.n563 B.n562 9.36635
R1021 B.n545 B.n50 9.36635
R1022 B.n292 B.n291 9.36635
R1023 B.n310 B.n309 9.36635
R1024 B.n681 B.n0 8.11757
R1025 B.n681 B.n1 8.11757
R1026 B.n562 B.n561 1.24928
R1027 B.n548 B.n50 1.24928
R1028 B.n291 B.n136 1.24928
R1029 B.n309 B.n308 1.24928
R1030 VP.n0 VP.t1 186.821
R1031 VP.n0 VP.t0 138.172
R1032 VP VP.n0 0.526373
R1033 VTAIL.n306 VTAIL.n234 756.745
R1034 VTAIL.n72 VTAIL.n0 756.745
R1035 VTAIL.n228 VTAIL.n156 756.745
R1036 VTAIL.n150 VTAIL.n78 756.745
R1037 VTAIL.n258 VTAIL.n257 585
R1038 VTAIL.n263 VTAIL.n262 585
R1039 VTAIL.n265 VTAIL.n264 585
R1040 VTAIL.n254 VTAIL.n253 585
R1041 VTAIL.n271 VTAIL.n270 585
R1042 VTAIL.n273 VTAIL.n272 585
R1043 VTAIL.n250 VTAIL.n249 585
R1044 VTAIL.n280 VTAIL.n279 585
R1045 VTAIL.n281 VTAIL.n248 585
R1046 VTAIL.n283 VTAIL.n282 585
R1047 VTAIL.n246 VTAIL.n245 585
R1048 VTAIL.n289 VTAIL.n288 585
R1049 VTAIL.n291 VTAIL.n290 585
R1050 VTAIL.n242 VTAIL.n241 585
R1051 VTAIL.n297 VTAIL.n296 585
R1052 VTAIL.n299 VTAIL.n298 585
R1053 VTAIL.n238 VTAIL.n237 585
R1054 VTAIL.n305 VTAIL.n304 585
R1055 VTAIL.n307 VTAIL.n306 585
R1056 VTAIL.n24 VTAIL.n23 585
R1057 VTAIL.n29 VTAIL.n28 585
R1058 VTAIL.n31 VTAIL.n30 585
R1059 VTAIL.n20 VTAIL.n19 585
R1060 VTAIL.n37 VTAIL.n36 585
R1061 VTAIL.n39 VTAIL.n38 585
R1062 VTAIL.n16 VTAIL.n15 585
R1063 VTAIL.n46 VTAIL.n45 585
R1064 VTAIL.n47 VTAIL.n14 585
R1065 VTAIL.n49 VTAIL.n48 585
R1066 VTAIL.n12 VTAIL.n11 585
R1067 VTAIL.n55 VTAIL.n54 585
R1068 VTAIL.n57 VTAIL.n56 585
R1069 VTAIL.n8 VTAIL.n7 585
R1070 VTAIL.n63 VTAIL.n62 585
R1071 VTAIL.n65 VTAIL.n64 585
R1072 VTAIL.n4 VTAIL.n3 585
R1073 VTAIL.n71 VTAIL.n70 585
R1074 VTAIL.n73 VTAIL.n72 585
R1075 VTAIL.n229 VTAIL.n228 585
R1076 VTAIL.n227 VTAIL.n226 585
R1077 VTAIL.n160 VTAIL.n159 585
R1078 VTAIL.n221 VTAIL.n220 585
R1079 VTAIL.n219 VTAIL.n218 585
R1080 VTAIL.n164 VTAIL.n163 585
R1081 VTAIL.n213 VTAIL.n212 585
R1082 VTAIL.n211 VTAIL.n210 585
R1083 VTAIL.n168 VTAIL.n167 585
R1084 VTAIL.n205 VTAIL.n204 585
R1085 VTAIL.n203 VTAIL.n170 585
R1086 VTAIL.n202 VTAIL.n201 585
R1087 VTAIL.n173 VTAIL.n171 585
R1088 VTAIL.n196 VTAIL.n195 585
R1089 VTAIL.n194 VTAIL.n193 585
R1090 VTAIL.n177 VTAIL.n176 585
R1091 VTAIL.n188 VTAIL.n187 585
R1092 VTAIL.n186 VTAIL.n185 585
R1093 VTAIL.n181 VTAIL.n180 585
R1094 VTAIL.n151 VTAIL.n150 585
R1095 VTAIL.n149 VTAIL.n148 585
R1096 VTAIL.n82 VTAIL.n81 585
R1097 VTAIL.n143 VTAIL.n142 585
R1098 VTAIL.n141 VTAIL.n140 585
R1099 VTAIL.n86 VTAIL.n85 585
R1100 VTAIL.n135 VTAIL.n134 585
R1101 VTAIL.n133 VTAIL.n132 585
R1102 VTAIL.n90 VTAIL.n89 585
R1103 VTAIL.n127 VTAIL.n126 585
R1104 VTAIL.n125 VTAIL.n92 585
R1105 VTAIL.n124 VTAIL.n123 585
R1106 VTAIL.n95 VTAIL.n93 585
R1107 VTAIL.n118 VTAIL.n117 585
R1108 VTAIL.n116 VTAIL.n115 585
R1109 VTAIL.n99 VTAIL.n98 585
R1110 VTAIL.n110 VTAIL.n109 585
R1111 VTAIL.n108 VTAIL.n107 585
R1112 VTAIL.n103 VTAIL.n102 585
R1113 VTAIL.n259 VTAIL.t1 329.036
R1114 VTAIL.n25 VTAIL.t2 329.036
R1115 VTAIL.n104 VTAIL.t0 329.036
R1116 VTAIL.n182 VTAIL.t3 329.036
R1117 VTAIL.n263 VTAIL.n257 171.744
R1118 VTAIL.n264 VTAIL.n263 171.744
R1119 VTAIL.n264 VTAIL.n253 171.744
R1120 VTAIL.n271 VTAIL.n253 171.744
R1121 VTAIL.n272 VTAIL.n271 171.744
R1122 VTAIL.n272 VTAIL.n249 171.744
R1123 VTAIL.n280 VTAIL.n249 171.744
R1124 VTAIL.n281 VTAIL.n280 171.744
R1125 VTAIL.n282 VTAIL.n281 171.744
R1126 VTAIL.n282 VTAIL.n245 171.744
R1127 VTAIL.n289 VTAIL.n245 171.744
R1128 VTAIL.n290 VTAIL.n289 171.744
R1129 VTAIL.n290 VTAIL.n241 171.744
R1130 VTAIL.n297 VTAIL.n241 171.744
R1131 VTAIL.n298 VTAIL.n297 171.744
R1132 VTAIL.n298 VTAIL.n237 171.744
R1133 VTAIL.n305 VTAIL.n237 171.744
R1134 VTAIL.n306 VTAIL.n305 171.744
R1135 VTAIL.n29 VTAIL.n23 171.744
R1136 VTAIL.n30 VTAIL.n29 171.744
R1137 VTAIL.n30 VTAIL.n19 171.744
R1138 VTAIL.n37 VTAIL.n19 171.744
R1139 VTAIL.n38 VTAIL.n37 171.744
R1140 VTAIL.n38 VTAIL.n15 171.744
R1141 VTAIL.n46 VTAIL.n15 171.744
R1142 VTAIL.n47 VTAIL.n46 171.744
R1143 VTAIL.n48 VTAIL.n47 171.744
R1144 VTAIL.n48 VTAIL.n11 171.744
R1145 VTAIL.n55 VTAIL.n11 171.744
R1146 VTAIL.n56 VTAIL.n55 171.744
R1147 VTAIL.n56 VTAIL.n7 171.744
R1148 VTAIL.n63 VTAIL.n7 171.744
R1149 VTAIL.n64 VTAIL.n63 171.744
R1150 VTAIL.n64 VTAIL.n3 171.744
R1151 VTAIL.n71 VTAIL.n3 171.744
R1152 VTAIL.n72 VTAIL.n71 171.744
R1153 VTAIL.n228 VTAIL.n227 171.744
R1154 VTAIL.n227 VTAIL.n159 171.744
R1155 VTAIL.n220 VTAIL.n159 171.744
R1156 VTAIL.n220 VTAIL.n219 171.744
R1157 VTAIL.n219 VTAIL.n163 171.744
R1158 VTAIL.n212 VTAIL.n163 171.744
R1159 VTAIL.n212 VTAIL.n211 171.744
R1160 VTAIL.n211 VTAIL.n167 171.744
R1161 VTAIL.n204 VTAIL.n167 171.744
R1162 VTAIL.n204 VTAIL.n203 171.744
R1163 VTAIL.n203 VTAIL.n202 171.744
R1164 VTAIL.n202 VTAIL.n171 171.744
R1165 VTAIL.n195 VTAIL.n171 171.744
R1166 VTAIL.n195 VTAIL.n194 171.744
R1167 VTAIL.n194 VTAIL.n176 171.744
R1168 VTAIL.n187 VTAIL.n176 171.744
R1169 VTAIL.n187 VTAIL.n186 171.744
R1170 VTAIL.n186 VTAIL.n180 171.744
R1171 VTAIL.n150 VTAIL.n149 171.744
R1172 VTAIL.n149 VTAIL.n81 171.744
R1173 VTAIL.n142 VTAIL.n81 171.744
R1174 VTAIL.n142 VTAIL.n141 171.744
R1175 VTAIL.n141 VTAIL.n85 171.744
R1176 VTAIL.n134 VTAIL.n85 171.744
R1177 VTAIL.n134 VTAIL.n133 171.744
R1178 VTAIL.n133 VTAIL.n89 171.744
R1179 VTAIL.n126 VTAIL.n89 171.744
R1180 VTAIL.n126 VTAIL.n125 171.744
R1181 VTAIL.n125 VTAIL.n124 171.744
R1182 VTAIL.n124 VTAIL.n93 171.744
R1183 VTAIL.n117 VTAIL.n93 171.744
R1184 VTAIL.n117 VTAIL.n116 171.744
R1185 VTAIL.n116 VTAIL.n98 171.744
R1186 VTAIL.n109 VTAIL.n98 171.744
R1187 VTAIL.n109 VTAIL.n108 171.744
R1188 VTAIL.n108 VTAIL.n102 171.744
R1189 VTAIL.t1 VTAIL.n257 85.8723
R1190 VTAIL.t2 VTAIL.n23 85.8723
R1191 VTAIL.t3 VTAIL.n180 85.8723
R1192 VTAIL.t0 VTAIL.n102 85.8723
R1193 VTAIL.n311 VTAIL.n310 31.7975
R1194 VTAIL.n77 VTAIL.n76 31.7975
R1195 VTAIL.n233 VTAIL.n232 31.7975
R1196 VTAIL.n155 VTAIL.n154 31.7975
R1197 VTAIL.n155 VTAIL.n77 31.1945
R1198 VTAIL.n311 VTAIL.n233 27.9272
R1199 VTAIL.n283 VTAIL.n248 13.1884
R1200 VTAIL.n49 VTAIL.n14 13.1884
R1201 VTAIL.n205 VTAIL.n170 13.1884
R1202 VTAIL.n127 VTAIL.n92 13.1884
R1203 VTAIL.n279 VTAIL.n278 12.8005
R1204 VTAIL.n284 VTAIL.n246 12.8005
R1205 VTAIL.n45 VTAIL.n44 12.8005
R1206 VTAIL.n50 VTAIL.n12 12.8005
R1207 VTAIL.n206 VTAIL.n168 12.8005
R1208 VTAIL.n201 VTAIL.n172 12.8005
R1209 VTAIL.n128 VTAIL.n90 12.8005
R1210 VTAIL.n123 VTAIL.n94 12.8005
R1211 VTAIL.n277 VTAIL.n250 12.0247
R1212 VTAIL.n288 VTAIL.n287 12.0247
R1213 VTAIL.n43 VTAIL.n16 12.0247
R1214 VTAIL.n54 VTAIL.n53 12.0247
R1215 VTAIL.n210 VTAIL.n209 12.0247
R1216 VTAIL.n200 VTAIL.n173 12.0247
R1217 VTAIL.n132 VTAIL.n131 12.0247
R1218 VTAIL.n122 VTAIL.n95 12.0247
R1219 VTAIL.n274 VTAIL.n273 11.249
R1220 VTAIL.n291 VTAIL.n244 11.249
R1221 VTAIL.n40 VTAIL.n39 11.249
R1222 VTAIL.n57 VTAIL.n10 11.249
R1223 VTAIL.n213 VTAIL.n166 11.249
R1224 VTAIL.n197 VTAIL.n196 11.249
R1225 VTAIL.n135 VTAIL.n88 11.249
R1226 VTAIL.n119 VTAIL.n118 11.249
R1227 VTAIL.n259 VTAIL.n258 10.7239
R1228 VTAIL.n25 VTAIL.n24 10.7239
R1229 VTAIL.n182 VTAIL.n181 10.7239
R1230 VTAIL.n104 VTAIL.n103 10.7239
R1231 VTAIL.n270 VTAIL.n252 10.4732
R1232 VTAIL.n292 VTAIL.n242 10.4732
R1233 VTAIL.n36 VTAIL.n18 10.4732
R1234 VTAIL.n58 VTAIL.n8 10.4732
R1235 VTAIL.n214 VTAIL.n164 10.4732
R1236 VTAIL.n193 VTAIL.n175 10.4732
R1237 VTAIL.n136 VTAIL.n86 10.4732
R1238 VTAIL.n115 VTAIL.n97 10.4732
R1239 VTAIL.n269 VTAIL.n254 9.69747
R1240 VTAIL.n296 VTAIL.n295 9.69747
R1241 VTAIL.n35 VTAIL.n20 9.69747
R1242 VTAIL.n62 VTAIL.n61 9.69747
R1243 VTAIL.n218 VTAIL.n217 9.69747
R1244 VTAIL.n192 VTAIL.n177 9.69747
R1245 VTAIL.n140 VTAIL.n139 9.69747
R1246 VTAIL.n114 VTAIL.n99 9.69747
R1247 VTAIL.n310 VTAIL.n309 9.45567
R1248 VTAIL.n76 VTAIL.n75 9.45567
R1249 VTAIL.n232 VTAIL.n231 9.45567
R1250 VTAIL.n154 VTAIL.n153 9.45567
R1251 VTAIL.n236 VTAIL.n235 9.3005
R1252 VTAIL.n309 VTAIL.n308 9.3005
R1253 VTAIL.n301 VTAIL.n300 9.3005
R1254 VTAIL.n240 VTAIL.n239 9.3005
R1255 VTAIL.n295 VTAIL.n294 9.3005
R1256 VTAIL.n293 VTAIL.n292 9.3005
R1257 VTAIL.n244 VTAIL.n243 9.3005
R1258 VTAIL.n287 VTAIL.n286 9.3005
R1259 VTAIL.n285 VTAIL.n284 9.3005
R1260 VTAIL.n261 VTAIL.n260 9.3005
R1261 VTAIL.n256 VTAIL.n255 9.3005
R1262 VTAIL.n267 VTAIL.n266 9.3005
R1263 VTAIL.n269 VTAIL.n268 9.3005
R1264 VTAIL.n252 VTAIL.n251 9.3005
R1265 VTAIL.n275 VTAIL.n274 9.3005
R1266 VTAIL.n277 VTAIL.n276 9.3005
R1267 VTAIL.n278 VTAIL.n247 9.3005
R1268 VTAIL.n303 VTAIL.n302 9.3005
R1269 VTAIL.n2 VTAIL.n1 9.3005
R1270 VTAIL.n75 VTAIL.n74 9.3005
R1271 VTAIL.n67 VTAIL.n66 9.3005
R1272 VTAIL.n6 VTAIL.n5 9.3005
R1273 VTAIL.n61 VTAIL.n60 9.3005
R1274 VTAIL.n59 VTAIL.n58 9.3005
R1275 VTAIL.n10 VTAIL.n9 9.3005
R1276 VTAIL.n53 VTAIL.n52 9.3005
R1277 VTAIL.n51 VTAIL.n50 9.3005
R1278 VTAIL.n27 VTAIL.n26 9.3005
R1279 VTAIL.n22 VTAIL.n21 9.3005
R1280 VTAIL.n33 VTAIL.n32 9.3005
R1281 VTAIL.n35 VTAIL.n34 9.3005
R1282 VTAIL.n18 VTAIL.n17 9.3005
R1283 VTAIL.n41 VTAIL.n40 9.3005
R1284 VTAIL.n43 VTAIL.n42 9.3005
R1285 VTAIL.n44 VTAIL.n13 9.3005
R1286 VTAIL.n69 VTAIL.n68 9.3005
R1287 VTAIL.n158 VTAIL.n157 9.3005
R1288 VTAIL.n225 VTAIL.n224 9.3005
R1289 VTAIL.n223 VTAIL.n222 9.3005
R1290 VTAIL.n162 VTAIL.n161 9.3005
R1291 VTAIL.n217 VTAIL.n216 9.3005
R1292 VTAIL.n215 VTAIL.n214 9.3005
R1293 VTAIL.n166 VTAIL.n165 9.3005
R1294 VTAIL.n209 VTAIL.n208 9.3005
R1295 VTAIL.n207 VTAIL.n206 9.3005
R1296 VTAIL.n172 VTAIL.n169 9.3005
R1297 VTAIL.n200 VTAIL.n199 9.3005
R1298 VTAIL.n198 VTAIL.n197 9.3005
R1299 VTAIL.n175 VTAIL.n174 9.3005
R1300 VTAIL.n192 VTAIL.n191 9.3005
R1301 VTAIL.n190 VTAIL.n189 9.3005
R1302 VTAIL.n179 VTAIL.n178 9.3005
R1303 VTAIL.n184 VTAIL.n183 9.3005
R1304 VTAIL.n231 VTAIL.n230 9.3005
R1305 VTAIL.n106 VTAIL.n105 9.3005
R1306 VTAIL.n101 VTAIL.n100 9.3005
R1307 VTAIL.n112 VTAIL.n111 9.3005
R1308 VTAIL.n114 VTAIL.n113 9.3005
R1309 VTAIL.n97 VTAIL.n96 9.3005
R1310 VTAIL.n120 VTAIL.n119 9.3005
R1311 VTAIL.n122 VTAIL.n121 9.3005
R1312 VTAIL.n94 VTAIL.n91 9.3005
R1313 VTAIL.n153 VTAIL.n152 9.3005
R1314 VTAIL.n80 VTAIL.n79 9.3005
R1315 VTAIL.n147 VTAIL.n146 9.3005
R1316 VTAIL.n145 VTAIL.n144 9.3005
R1317 VTAIL.n84 VTAIL.n83 9.3005
R1318 VTAIL.n139 VTAIL.n138 9.3005
R1319 VTAIL.n137 VTAIL.n136 9.3005
R1320 VTAIL.n88 VTAIL.n87 9.3005
R1321 VTAIL.n131 VTAIL.n130 9.3005
R1322 VTAIL.n129 VTAIL.n128 9.3005
R1323 VTAIL.n266 VTAIL.n265 8.92171
R1324 VTAIL.n299 VTAIL.n240 8.92171
R1325 VTAIL.n32 VTAIL.n31 8.92171
R1326 VTAIL.n65 VTAIL.n6 8.92171
R1327 VTAIL.n221 VTAIL.n162 8.92171
R1328 VTAIL.n189 VTAIL.n188 8.92171
R1329 VTAIL.n143 VTAIL.n84 8.92171
R1330 VTAIL.n111 VTAIL.n110 8.92171
R1331 VTAIL.n262 VTAIL.n256 8.14595
R1332 VTAIL.n300 VTAIL.n238 8.14595
R1333 VTAIL.n310 VTAIL.n234 8.14595
R1334 VTAIL.n28 VTAIL.n22 8.14595
R1335 VTAIL.n66 VTAIL.n4 8.14595
R1336 VTAIL.n76 VTAIL.n0 8.14595
R1337 VTAIL.n232 VTAIL.n156 8.14595
R1338 VTAIL.n222 VTAIL.n160 8.14595
R1339 VTAIL.n185 VTAIL.n179 8.14595
R1340 VTAIL.n154 VTAIL.n78 8.14595
R1341 VTAIL.n144 VTAIL.n82 8.14595
R1342 VTAIL.n107 VTAIL.n101 8.14595
R1343 VTAIL.n261 VTAIL.n258 7.3702
R1344 VTAIL.n304 VTAIL.n303 7.3702
R1345 VTAIL.n308 VTAIL.n307 7.3702
R1346 VTAIL.n27 VTAIL.n24 7.3702
R1347 VTAIL.n70 VTAIL.n69 7.3702
R1348 VTAIL.n74 VTAIL.n73 7.3702
R1349 VTAIL.n230 VTAIL.n229 7.3702
R1350 VTAIL.n226 VTAIL.n225 7.3702
R1351 VTAIL.n184 VTAIL.n181 7.3702
R1352 VTAIL.n152 VTAIL.n151 7.3702
R1353 VTAIL.n148 VTAIL.n147 7.3702
R1354 VTAIL.n106 VTAIL.n103 7.3702
R1355 VTAIL.n304 VTAIL.n236 6.59444
R1356 VTAIL.n307 VTAIL.n236 6.59444
R1357 VTAIL.n70 VTAIL.n2 6.59444
R1358 VTAIL.n73 VTAIL.n2 6.59444
R1359 VTAIL.n229 VTAIL.n158 6.59444
R1360 VTAIL.n226 VTAIL.n158 6.59444
R1361 VTAIL.n151 VTAIL.n80 6.59444
R1362 VTAIL.n148 VTAIL.n80 6.59444
R1363 VTAIL.n262 VTAIL.n261 5.81868
R1364 VTAIL.n303 VTAIL.n238 5.81868
R1365 VTAIL.n308 VTAIL.n234 5.81868
R1366 VTAIL.n28 VTAIL.n27 5.81868
R1367 VTAIL.n69 VTAIL.n4 5.81868
R1368 VTAIL.n74 VTAIL.n0 5.81868
R1369 VTAIL.n230 VTAIL.n156 5.81868
R1370 VTAIL.n225 VTAIL.n160 5.81868
R1371 VTAIL.n185 VTAIL.n184 5.81868
R1372 VTAIL.n152 VTAIL.n78 5.81868
R1373 VTAIL.n147 VTAIL.n82 5.81868
R1374 VTAIL.n107 VTAIL.n106 5.81868
R1375 VTAIL.n265 VTAIL.n256 5.04292
R1376 VTAIL.n300 VTAIL.n299 5.04292
R1377 VTAIL.n31 VTAIL.n22 5.04292
R1378 VTAIL.n66 VTAIL.n65 5.04292
R1379 VTAIL.n222 VTAIL.n221 5.04292
R1380 VTAIL.n188 VTAIL.n179 5.04292
R1381 VTAIL.n144 VTAIL.n143 5.04292
R1382 VTAIL.n110 VTAIL.n101 5.04292
R1383 VTAIL.n266 VTAIL.n254 4.26717
R1384 VTAIL.n296 VTAIL.n240 4.26717
R1385 VTAIL.n32 VTAIL.n20 4.26717
R1386 VTAIL.n62 VTAIL.n6 4.26717
R1387 VTAIL.n218 VTAIL.n162 4.26717
R1388 VTAIL.n189 VTAIL.n177 4.26717
R1389 VTAIL.n140 VTAIL.n84 4.26717
R1390 VTAIL.n111 VTAIL.n99 4.26717
R1391 VTAIL.n270 VTAIL.n269 3.49141
R1392 VTAIL.n295 VTAIL.n242 3.49141
R1393 VTAIL.n36 VTAIL.n35 3.49141
R1394 VTAIL.n61 VTAIL.n8 3.49141
R1395 VTAIL.n217 VTAIL.n164 3.49141
R1396 VTAIL.n193 VTAIL.n192 3.49141
R1397 VTAIL.n139 VTAIL.n86 3.49141
R1398 VTAIL.n115 VTAIL.n114 3.49141
R1399 VTAIL.n273 VTAIL.n252 2.71565
R1400 VTAIL.n292 VTAIL.n291 2.71565
R1401 VTAIL.n39 VTAIL.n18 2.71565
R1402 VTAIL.n58 VTAIL.n57 2.71565
R1403 VTAIL.n214 VTAIL.n213 2.71565
R1404 VTAIL.n196 VTAIL.n175 2.71565
R1405 VTAIL.n136 VTAIL.n135 2.71565
R1406 VTAIL.n118 VTAIL.n97 2.71565
R1407 VTAIL.n183 VTAIL.n182 2.41282
R1408 VTAIL.n105 VTAIL.n104 2.41282
R1409 VTAIL.n260 VTAIL.n259 2.41282
R1410 VTAIL.n26 VTAIL.n25 2.41282
R1411 VTAIL.n233 VTAIL.n155 2.10395
R1412 VTAIL.n274 VTAIL.n250 1.93989
R1413 VTAIL.n288 VTAIL.n244 1.93989
R1414 VTAIL.n40 VTAIL.n16 1.93989
R1415 VTAIL.n54 VTAIL.n10 1.93989
R1416 VTAIL.n210 VTAIL.n166 1.93989
R1417 VTAIL.n197 VTAIL.n173 1.93989
R1418 VTAIL.n132 VTAIL.n88 1.93989
R1419 VTAIL.n119 VTAIL.n95 1.93989
R1420 VTAIL VTAIL.n77 1.34533
R1421 VTAIL.n279 VTAIL.n277 1.16414
R1422 VTAIL.n287 VTAIL.n246 1.16414
R1423 VTAIL.n45 VTAIL.n43 1.16414
R1424 VTAIL.n53 VTAIL.n12 1.16414
R1425 VTAIL.n209 VTAIL.n168 1.16414
R1426 VTAIL.n201 VTAIL.n200 1.16414
R1427 VTAIL.n131 VTAIL.n90 1.16414
R1428 VTAIL.n123 VTAIL.n122 1.16414
R1429 VTAIL VTAIL.n311 0.759121
R1430 VTAIL.n278 VTAIL.n248 0.388379
R1431 VTAIL.n284 VTAIL.n283 0.388379
R1432 VTAIL.n44 VTAIL.n14 0.388379
R1433 VTAIL.n50 VTAIL.n49 0.388379
R1434 VTAIL.n206 VTAIL.n205 0.388379
R1435 VTAIL.n172 VTAIL.n170 0.388379
R1436 VTAIL.n128 VTAIL.n127 0.388379
R1437 VTAIL.n94 VTAIL.n92 0.388379
R1438 VTAIL.n260 VTAIL.n255 0.155672
R1439 VTAIL.n267 VTAIL.n255 0.155672
R1440 VTAIL.n268 VTAIL.n267 0.155672
R1441 VTAIL.n268 VTAIL.n251 0.155672
R1442 VTAIL.n275 VTAIL.n251 0.155672
R1443 VTAIL.n276 VTAIL.n275 0.155672
R1444 VTAIL.n276 VTAIL.n247 0.155672
R1445 VTAIL.n285 VTAIL.n247 0.155672
R1446 VTAIL.n286 VTAIL.n285 0.155672
R1447 VTAIL.n286 VTAIL.n243 0.155672
R1448 VTAIL.n293 VTAIL.n243 0.155672
R1449 VTAIL.n294 VTAIL.n293 0.155672
R1450 VTAIL.n294 VTAIL.n239 0.155672
R1451 VTAIL.n301 VTAIL.n239 0.155672
R1452 VTAIL.n302 VTAIL.n301 0.155672
R1453 VTAIL.n302 VTAIL.n235 0.155672
R1454 VTAIL.n309 VTAIL.n235 0.155672
R1455 VTAIL.n26 VTAIL.n21 0.155672
R1456 VTAIL.n33 VTAIL.n21 0.155672
R1457 VTAIL.n34 VTAIL.n33 0.155672
R1458 VTAIL.n34 VTAIL.n17 0.155672
R1459 VTAIL.n41 VTAIL.n17 0.155672
R1460 VTAIL.n42 VTAIL.n41 0.155672
R1461 VTAIL.n42 VTAIL.n13 0.155672
R1462 VTAIL.n51 VTAIL.n13 0.155672
R1463 VTAIL.n52 VTAIL.n51 0.155672
R1464 VTAIL.n52 VTAIL.n9 0.155672
R1465 VTAIL.n59 VTAIL.n9 0.155672
R1466 VTAIL.n60 VTAIL.n59 0.155672
R1467 VTAIL.n60 VTAIL.n5 0.155672
R1468 VTAIL.n67 VTAIL.n5 0.155672
R1469 VTAIL.n68 VTAIL.n67 0.155672
R1470 VTAIL.n68 VTAIL.n1 0.155672
R1471 VTAIL.n75 VTAIL.n1 0.155672
R1472 VTAIL.n231 VTAIL.n157 0.155672
R1473 VTAIL.n224 VTAIL.n157 0.155672
R1474 VTAIL.n224 VTAIL.n223 0.155672
R1475 VTAIL.n223 VTAIL.n161 0.155672
R1476 VTAIL.n216 VTAIL.n161 0.155672
R1477 VTAIL.n216 VTAIL.n215 0.155672
R1478 VTAIL.n215 VTAIL.n165 0.155672
R1479 VTAIL.n208 VTAIL.n165 0.155672
R1480 VTAIL.n208 VTAIL.n207 0.155672
R1481 VTAIL.n207 VTAIL.n169 0.155672
R1482 VTAIL.n199 VTAIL.n169 0.155672
R1483 VTAIL.n199 VTAIL.n198 0.155672
R1484 VTAIL.n198 VTAIL.n174 0.155672
R1485 VTAIL.n191 VTAIL.n174 0.155672
R1486 VTAIL.n191 VTAIL.n190 0.155672
R1487 VTAIL.n190 VTAIL.n178 0.155672
R1488 VTAIL.n183 VTAIL.n178 0.155672
R1489 VTAIL.n153 VTAIL.n79 0.155672
R1490 VTAIL.n146 VTAIL.n79 0.155672
R1491 VTAIL.n146 VTAIL.n145 0.155672
R1492 VTAIL.n145 VTAIL.n83 0.155672
R1493 VTAIL.n138 VTAIL.n83 0.155672
R1494 VTAIL.n138 VTAIL.n137 0.155672
R1495 VTAIL.n137 VTAIL.n87 0.155672
R1496 VTAIL.n130 VTAIL.n87 0.155672
R1497 VTAIL.n130 VTAIL.n129 0.155672
R1498 VTAIL.n129 VTAIL.n91 0.155672
R1499 VTAIL.n121 VTAIL.n91 0.155672
R1500 VTAIL.n121 VTAIL.n120 0.155672
R1501 VTAIL.n120 VTAIL.n96 0.155672
R1502 VTAIL.n113 VTAIL.n96 0.155672
R1503 VTAIL.n113 VTAIL.n112 0.155672
R1504 VTAIL.n112 VTAIL.n100 0.155672
R1505 VTAIL.n105 VTAIL.n100 0.155672
R1506 VDD1.n72 VDD1.n0 756.745
R1507 VDD1.n149 VDD1.n77 756.745
R1508 VDD1.n73 VDD1.n72 585
R1509 VDD1.n71 VDD1.n70 585
R1510 VDD1.n4 VDD1.n3 585
R1511 VDD1.n65 VDD1.n64 585
R1512 VDD1.n63 VDD1.n62 585
R1513 VDD1.n8 VDD1.n7 585
R1514 VDD1.n57 VDD1.n56 585
R1515 VDD1.n55 VDD1.n54 585
R1516 VDD1.n12 VDD1.n11 585
R1517 VDD1.n49 VDD1.n48 585
R1518 VDD1.n47 VDD1.n14 585
R1519 VDD1.n46 VDD1.n45 585
R1520 VDD1.n17 VDD1.n15 585
R1521 VDD1.n40 VDD1.n39 585
R1522 VDD1.n38 VDD1.n37 585
R1523 VDD1.n21 VDD1.n20 585
R1524 VDD1.n32 VDD1.n31 585
R1525 VDD1.n30 VDD1.n29 585
R1526 VDD1.n25 VDD1.n24 585
R1527 VDD1.n101 VDD1.n100 585
R1528 VDD1.n106 VDD1.n105 585
R1529 VDD1.n108 VDD1.n107 585
R1530 VDD1.n97 VDD1.n96 585
R1531 VDD1.n114 VDD1.n113 585
R1532 VDD1.n116 VDD1.n115 585
R1533 VDD1.n93 VDD1.n92 585
R1534 VDD1.n123 VDD1.n122 585
R1535 VDD1.n124 VDD1.n91 585
R1536 VDD1.n126 VDD1.n125 585
R1537 VDD1.n89 VDD1.n88 585
R1538 VDD1.n132 VDD1.n131 585
R1539 VDD1.n134 VDD1.n133 585
R1540 VDD1.n85 VDD1.n84 585
R1541 VDD1.n140 VDD1.n139 585
R1542 VDD1.n142 VDD1.n141 585
R1543 VDD1.n81 VDD1.n80 585
R1544 VDD1.n148 VDD1.n147 585
R1545 VDD1.n150 VDD1.n149 585
R1546 VDD1.n102 VDD1.t1 329.036
R1547 VDD1.n26 VDD1.t0 329.036
R1548 VDD1.n72 VDD1.n71 171.744
R1549 VDD1.n71 VDD1.n3 171.744
R1550 VDD1.n64 VDD1.n3 171.744
R1551 VDD1.n64 VDD1.n63 171.744
R1552 VDD1.n63 VDD1.n7 171.744
R1553 VDD1.n56 VDD1.n7 171.744
R1554 VDD1.n56 VDD1.n55 171.744
R1555 VDD1.n55 VDD1.n11 171.744
R1556 VDD1.n48 VDD1.n11 171.744
R1557 VDD1.n48 VDD1.n47 171.744
R1558 VDD1.n47 VDD1.n46 171.744
R1559 VDD1.n46 VDD1.n15 171.744
R1560 VDD1.n39 VDD1.n15 171.744
R1561 VDD1.n39 VDD1.n38 171.744
R1562 VDD1.n38 VDD1.n20 171.744
R1563 VDD1.n31 VDD1.n20 171.744
R1564 VDD1.n31 VDD1.n30 171.744
R1565 VDD1.n30 VDD1.n24 171.744
R1566 VDD1.n106 VDD1.n100 171.744
R1567 VDD1.n107 VDD1.n106 171.744
R1568 VDD1.n107 VDD1.n96 171.744
R1569 VDD1.n114 VDD1.n96 171.744
R1570 VDD1.n115 VDD1.n114 171.744
R1571 VDD1.n115 VDD1.n92 171.744
R1572 VDD1.n123 VDD1.n92 171.744
R1573 VDD1.n124 VDD1.n123 171.744
R1574 VDD1.n125 VDD1.n124 171.744
R1575 VDD1.n125 VDD1.n88 171.744
R1576 VDD1.n132 VDD1.n88 171.744
R1577 VDD1.n133 VDD1.n132 171.744
R1578 VDD1.n133 VDD1.n84 171.744
R1579 VDD1.n140 VDD1.n84 171.744
R1580 VDD1.n141 VDD1.n140 171.744
R1581 VDD1.n141 VDD1.n80 171.744
R1582 VDD1.n148 VDD1.n80 171.744
R1583 VDD1.n149 VDD1.n148 171.744
R1584 VDD1 VDD1.n153 92.3049
R1585 VDD1.t0 VDD1.n24 85.8723
R1586 VDD1.t1 VDD1.n100 85.8723
R1587 VDD1 VDD1.n76 49.3513
R1588 VDD1.n49 VDD1.n14 13.1884
R1589 VDD1.n126 VDD1.n91 13.1884
R1590 VDD1.n50 VDD1.n12 12.8005
R1591 VDD1.n45 VDD1.n16 12.8005
R1592 VDD1.n122 VDD1.n121 12.8005
R1593 VDD1.n127 VDD1.n89 12.8005
R1594 VDD1.n54 VDD1.n53 12.0247
R1595 VDD1.n44 VDD1.n17 12.0247
R1596 VDD1.n120 VDD1.n93 12.0247
R1597 VDD1.n131 VDD1.n130 12.0247
R1598 VDD1.n57 VDD1.n10 11.249
R1599 VDD1.n41 VDD1.n40 11.249
R1600 VDD1.n117 VDD1.n116 11.249
R1601 VDD1.n134 VDD1.n87 11.249
R1602 VDD1.n26 VDD1.n25 10.7239
R1603 VDD1.n102 VDD1.n101 10.7239
R1604 VDD1.n58 VDD1.n8 10.4732
R1605 VDD1.n37 VDD1.n19 10.4732
R1606 VDD1.n113 VDD1.n95 10.4732
R1607 VDD1.n135 VDD1.n85 10.4732
R1608 VDD1.n62 VDD1.n61 9.69747
R1609 VDD1.n36 VDD1.n21 9.69747
R1610 VDD1.n112 VDD1.n97 9.69747
R1611 VDD1.n139 VDD1.n138 9.69747
R1612 VDD1.n76 VDD1.n75 9.45567
R1613 VDD1.n153 VDD1.n152 9.45567
R1614 VDD1.n2 VDD1.n1 9.3005
R1615 VDD1.n69 VDD1.n68 9.3005
R1616 VDD1.n67 VDD1.n66 9.3005
R1617 VDD1.n6 VDD1.n5 9.3005
R1618 VDD1.n61 VDD1.n60 9.3005
R1619 VDD1.n59 VDD1.n58 9.3005
R1620 VDD1.n10 VDD1.n9 9.3005
R1621 VDD1.n53 VDD1.n52 9.3005
R1622 VDD1.n51 VDD1.n50 9.3005
R1623 VDD1.n16 VDD1.n13 9.3005
R1624 VDD1.n44 VDD1.n43 9.3005
R1625 VDD1.n42 VDD1.n41 9.3005
R1626 VDD1.n19 VDD1.n18 9.3005
R1627 VDD1.n36 VDD1.n35 9.3005
R1628 VDD1.n34 VDD1.n33 9.3005
R1629 VDD1.n23 VDD1.n22 9.3005
R1630 VDD1.n28 VDD1.n27 9.3005
R1631 VDD1.n75 VDD1.n74 9.3005
R1632 VDD1.n79 VDD1.n78 9.3005
R1633 VDD1.n152 VDD1.n151 9.3005
R1634 VDD1.n144 VDD1.n143 9.3005
R1635 VDD1.n83 VDD1.n82 9.3005
R1636 VDD1.n138 VDD1.n137 9.3005
R1637 VDD1.n136 VDD1.n135 9.3005
R1638 VDD1.n87 VDD1.n86 9.3005
R1639 VDD1.n130 VDD1.n129 9.3005
R1640 VDD1.n128 VDD1.n127 9.3005
R1641 VDD1.n104 VDD1.n103 9.3005
R1642 VDD1.n99 VDD1.n98 9.3005
R1643 VDD1.n110 VDD1.n109 9.3005
R1644 VDD1.n112 VDD1.n111 9.3005
R1645 VDD1.n95 VDD1.n94 9.3005
R1646 VDD1.n118 VDD1.n117 9.3005
R1647 VDD1.n120 VDD1.n119 9.3005
R1648 VDD1.n121 VDD1.n90 9.3005
R1649 VDD1.n146 VDD1.n145 9.3005
R1650 VDD1.n65 VDD1.n6 8.92171
R1651 VDD1.n33 VDD1.n32 8.92171
R1652 VDD1.n109 VDD1.n108 8.92171
R1653 VDD1.n142 VDD1.n83 8.92171
R1654 VDD1.n76 VDD1.n0 8.14595
R1655 VDD1.n66 VDD1.n4 8.14595
R1656 VDD1.n29 VDD1.n23 8.14595
R1657 VDD1.n105 VDD1.n99 8.14595
R1658 VDD1.n143 VDD1.n81 8.14595
R1659 VDD1.n153 VDD1.n77 8.14595
R1660 VDD1.n74 VDD1.n73 7.3702
R1661 VDD1.n70 VDD1.n69 7.3702
R1662 VDD1.n28 VDD1.n25 7.3702
R1663 VDD1.n104 VDD1.n101 7.3702
R1664 VDD1.n147 VDD1.n146 7.3702
R1665 VDD1.n151 VDD1.n150 7.3702
R1666 VDD1.n73 VDD1.n2 6.59444
R1667 VDD1.n70 VDD1.n2 6.59444
R1668 VDD1.n147 VDD1.n79 6.59444
R1669 VDD1.n150 VDD1.n79 6.59444
R1670 VDD1.n74 VDD1.n0 5.81868
R1671 VDD1.n69 VDD1.n4 5.81868
R1672 VDD1.n29 VDD1.n28 5.81868
R1673 VDD1.n105 VDD1.n104 5.81868
R1674 VDD1.n146 VDD1.n81 5.81868
R1675 VDD1.n151 VDD1.n77 5.81868
R1676 VDD1.n66 VDD1.n65 5.04292
R1677 VDD1.n32 VDD1.n23 5.04292
R1678 VDD1.n108 VDD1.n99 5.04292
R1679 VDD1.n143 VDD1.n142 5.04292
R1680 VDD1.n62 VDD1.n6 4.26717
R1681 VDD1.n33 VDD1.n21 4.26717
R1682 VDD1.n109 VDD1.n97 4.26717
R1683 VDD1.n139 VDD1.n83 4.26717
R1684 VDD1.n61 VDD1.n8 3.49141
R1685 VDD1.n37 VDD1.n36 3.49141
R1686 VDD1.n113 VDD1.n112 3.49141
R1687 VDD1.n138 VDD1.n85 3.49141
R1688 VDD1.n58 VDD1.n57 2.71565
R1689 VDD1.n40 VDD1.n19 2.71565
R1690 VDD1.n116 VDD1.n95 2.71565
R1691 VDD1.n135 VDD1.n134 2.71565
R1692 VDD1.n27 VDD1.n26 2.41282
R1693 VDD1.n103 VDD1.n102 2.41282
R1694 VDD1.n54 VDD1.n10 1.93989
R1695 VDD1.n41 VDD1.n17 1.93989
R1696 VDD1.n117 VDD1.n93 1.93989
R1697 VDD1.n131 VDD1.n87 1.93989
R1698 VDD1.n53 VDD1.n12 1.16414
R1699 VDD1.n45 VDD1.n44 1.16414
R1700 VDD1.n122 VDD1.n120 1.16414
R1701 VDD1.n130 VDD1.n89 1.16414
R1702 VDD1.n50 VDD1.n49 0.388379
R1703 VDD1.n16 VDD1.n14 0.388379
R1704 VDD1.n121 VDD1.n91 0.388379
R1705 VDD1.n127 VDD1.n126 0.388379
R1706 VDD1.n75 VDD1.n1 0.155672
R1707 VDD1.n68 VDD1.n1 0.155672
R1708 VDD1.n68 VDD1.n67 0.155672
R1709 VDD1.n67 VDD1.n5 0.155672
R1710 VDD1.n60 VDD1.n5 0.155672
R1711 VDD1.n60 VDD1.n59 0.155672
R1712 VDD1.n59 VDD1.n9 0.155672
R1713 VDD1.n52 VDD1.n9 0.155672
R1714 VDD1.n52 VDD1.n51 0.155672
R1715 VDD1.n51 VDD1.n13 0.155672
R1716 VDD1.n43 VDD1.n13 0.155672
R1717 VDD1.n43 VDD1.n42 0.155672
R1718 VDD1.n42 VDD1.n18 0.155672
R1719 VDD1.n35 VDD1.n18 0.155672
R1720 VDD1.n35 VDD1.n34 0.155672
R1721 VDD1.n34 VDD1.n22 0.155672
R1722 VDD1.n27 VDD1.n22 0.155672
R1723 VDD1.n103 VDD1.n98 0.155672
R1724 VDD1.n110 VDD1.n98 0.155672
R1725 VDD1.n111 VDD1.n110 0.155672
R1726 VDD1.n111 VDD1.n94 0.155672
R1727 VDD1.n118 VDD1.n94 0.155672
R1728 VDD1.n119 VDD1.n118 0.155672
R1729 VDD1.n119 VDD1.n90 0.155672
R1730 VDD1.n128 VDD1.n90 0.155672
R1731 VDD1.n129 VDD1.n128 0.155672
R1732 VDD1.n129 VDD1.n86 0.155672
R1733 VDD1.n136 VDD1.n86 0.155672
R1734 VDD1.n137 VDD1.n136 0.155672
R1735 VDD1.n137 VDD1.n82 0.155672
R1736 VDD1.n144 VDD1.n82 0.155672
R1737 VDD1.n145 VDD1.n144 0.155672
R1738 VDD1.n145 VDD1.n78 0.155672
R1739 VDD1.n152 VDD1.n78 0.155672
R1740 VN VN.t0 186.727
R1741 VN VN.t1 138.697
R1742 VDD2.n149 VDD2.n77 756.745
R1743 VDD2.n72 VDD2.n0 756.745
R1744 VDD2.n150 VDD2.n149 585
R1745 VDD2.n148 VDD2.n147 585
R1746 VDD2.n81 VDD2.n80 585
R1747 VDD2.n142 VDD2.n141 585
R1748 VDD2.n140 VDD2.n139 585
R1749 VDD2.n85 VDD2.n84 585
R1750 VDD2.n134 VDD2.n133 585
R1751 VDD2.n132 VDD2.n131 585
R1752 VDD2.n89 VDD2.n88 585
R1753 VDD2.n126 VDD2.n125 585
R1754 VDD2.n124 VDD2.n91 585
R1755 VDD2.n123 VDD2.n122 585
R1756 VDD2.n94 VDD2.n92 585
R1757 VDD2.n117 VDD2.n116 585
R1758 VDD2.n115 VDD2.n114 585
R1759 VDD2.n98 VDD2.n97 585
R1760 VDD2.n109 VDD2.n108 585
R1761 VDD2.n107 VDD2.n106 585
R1762 VDD2.n102 VDD2.n101 585
R1763 VDD2.n24 VDD2.n23 585
R1764 VDD2.n29 VDD2.n28 585
R1765 VDD2.n31 VDD2.n30 585
R1766 VDD2.n20 VDD2.n19 585
R1767 VDD2.n37 VDD2.n36 585
R1768 VDD2.n39 VDD2.n38 585
R1769 VDD2.n16 VDD2.n15 585
R1770 VDD2.n46 VDD2.n45 585
R1771 VDD2.n47 VDD2.n14 585
R1772 VDD2.n49 VDD2.n48 585
R1773 VDD2.n12 VDD2.n11 585
R1774 VDD2.n55 VDD2.n54 585
R1775 VDD2.n57 VDD2.n56 585
R1776 VDD2.n8 VDD2.n7 585
R1777 VDD2.n63 VDD2.n62 585
R1778 VDD2.n65 VDD2.n64 585
R1779 VDD2.n4 VDD2.n3 585
R1780 VDD2.n71 VDD2.n70 585
R1781 VDD2.n73 VDD2.n72 585
R1782 VDD2.n25 VDD2.t0 329.036
R1783 VDD2.n103 VDD2.t1 329.036
R1784 VDD2.n149 VDD2.n148 171.744
R1785 VDD2.n148 VDD2.n80 171.744
R1786 VDD2.n141 VDD2.n80 171.744
R1787 VDD2.n141 VDD2.n140 171.744
R1788 VDD2.n140 VDD2.n84 171.744
R1789 VDD2.n133 VDD2.n84 171.744
R1790 VDD2.n133 VDD2.n132 171.744
R1791 VDD2.n132 VDD2.n88 171.744
R1792 VDD2.n125 VDD2.n88 171.744
R1793 VDD2.n125 VDD2.n124 171.744
R1794 VDD2.n124 VDD2.n123 171.744
R1795 VDD2.n123 VDD2.n92 171.744
R1796 VDD2.n116 VDD2.n92 171.744
R1797 VDD2.n116 VDD2.n115 171.744
R1798 VDD2.n115 VDD2.n97 171.744
R1799 VDD2.n108 VDD2.n97 171.744
R1800 VDD2.n108 VDD2.n107 171.744
R1801 VDD2.n107 VDD2.n101 171.744
R1802 VDD2.n29 VDD2.n23 171.744
R1803 VDD2.n30 VDD2.n29 171.744
R1804 VDD2.n30 VDD2.n19 171.744
R1805 VDD2.n37 VDD2.n19 171.744
R1806 VDD2.n38 VDD2.n37 171.744
R1807 VDD2.n38 VDD2.n15 171.744
R1808 VDD2.n46 VDD2.n15 171.744
R1809 VDD2.n47 VDD2.n46 171.744
R1810 VDD2.n48 VDD2.n47 171.744
R1811 VDD2.n48 VDD2.n11 171.744
R1812 VDD2.n55 VDD2.n11 171.744
R1813 VDD2.n56 VDD2.n55 171.744
R1814 VDD2.n56 VDD2.n7 171.744
R1815 VDD2.n63 VDD2.n7 171.744
R1816 VDD2.n64 VDD2.n63 171.744
R1817 VDD2.n64 VDD2.n3 171.744
R1818 VDD2.n71 VDD2.n3 171.744
R1819 VDD2.n72 VDD2.n71 171.744
R1820 VDD2.n154 VDD2.n76 90.9633
R1821 VDD2.t1 VDD2.n101 85.8723
R1822 VDD2.t0 VDD2.n23 85.8723
R1823 VDD2.n154 VDD2.n153 48.4763
R1824 VDD2.n126 VDD2.n91 13.1884
R1825 VDD2.n49 VDD2.n14 13.1884
R1826 VDD2.n127 VDD2.n89 12.8005
R1827 VDD2.n122 VDD2.n93 12.8005
R1828 VDD2.n45 VDD2.n44 12.8005
R1829 VDD2.n50 VDD2.n12 12.8005
R1830 VDD2.n131 VDD2.n130 12.0247
R1831 VDD2.n121 VDD2.n94 12.0247
R1832 VDD2.n43 VDD2.n16 12.0247
R1833 VDD2.n54 VDD2.n53 12.0247
R1834 VDD2.n134 VDD2.n87 11.249
R1835 VDD2.n118 VDD2.n117 11.249
R1836 VDD2.n40 VDD2.n39 11.249
R1837 VDD2.n57 VDD2.n10 11.249
R1838 VDD2.n103 VDD2.n102 10.7239
R1839 VDD2.n25 VDD2.n24 10.7239
R1840 VDD2.n135 VDD2.n85 10.4732
R1841 VDD2.n114 VDD2.n96 10.4732
R1842 VDD2.n36 VDD2.n18 10.4732
R1843 VDD2.n58 VDD2.n8 10.4732
R1844 VDD2.n139 VDD2.n138 9.69747
R1845 VDD2.n113 VDD2.n98 9.69747
R1846 VDD2.n35 VDD2.n20 9.69747
R1847 VDD2.n62 VDD2.n61 9.69747
R1848 VDD2.n153 VDD2.n152 9.45567
R1849 VDD2.n76 VDD2.n75 9.45567
R1850 VDD2.n79 VDD2.n78 9.3005
R1851 VDD2.n146 VDD2.n145 9.3005
R1852 VDD2.n144 VDD2.n143 9.3005
R1853 VDD2.n83 VDD2.n82 9.3005
R1854 VDD2.n138 VDD2.n137 9.3005
R1855 VDD2.n136 VDD2.n135 9.3005
R1856 VDD2.n87 VDD2.n86 9.3005
R1857 VDD2.n130 VDD2.n129 9.3005
R1858 VDD2.n128 VDD2.n127 9.3005
R1859 VDD2.n93 VDD2.n90 9.3005
R1860 VDD2.n121 VDD2.n120 9.3005
R1861 VDD2.n119 VDD2.n118 9.3005
R1862 VDD2.n96 VDD2.n95 9.3005
R1863 VDD2.n113 VDD2.n112 9.3005
R1864 VDD2.n111 VDD2.n110 9.3005
R1865 VDD2.n100 VDD2.n99 9.3005
R1866 VDD2.n105 VDD2.n104 9.3005
R1867 VDD2.n152 VDD2.n151 9.3005
R1868 VDD2.n2 VDD2.n1 9.3005
R1869 VDD2.n75 VDD2.n74 9.3005
R1870 VDD2.n67 VDD2.n66 9.3005
R1871 VDD2.n6 VDD2.n5 9.3005
R1872 VDD2.n61 VDD2.n60 9.3005
R1873 VDD2.n59 VDD2.n58 9.3005
R1874 VDD2.n10 VDD2.n9 9.3005
R1875 VDD2.n53 VDD2.n52 9.3005
R1876 VDD2.n51 VDD2.n50 9.3005
R1877 VDD2.n27 VDD2.n26 9.3005
R1878 VDD2.n22 VDD2.n21 9.3005
R1879 VDD2.n33 VDD2.n32 9.3005
R1880 VDD2.n35 VDD2.n34 9.3005
R1881 VDD2.n18 VDD2.n17 9.3005
R1882 VDD2.n41 VDD2.n40 9.3005
R1883 VDD2.n43 VDD2.n42 9.3005
R1884 VDD2.n44 VDD2.n13 9.3005
R1885 VDD2.n69 VDD2.n68 9.3005
R1886 VDD2.n142 VDD2.n83 8.92171
R1887 VDD2.n110 VDD2.n109 8.92171
R1888 VDD2.n32 VDD2.n31 8.92171
R1889 VDD2.n65 VDD2.n6 8.92171
R1890 VDD2.n153 VDD2.n77 8.14595
R1891 VDD2.n143 VDD2.n81 8.14595
R1892 VDD2.n106 VDD2.n100 8.14595
R1893 VDD2.n28 VDD2.n22 8.14595
R1894 VDD2.n66 VDD2.n4 8.14595
R1895 VDD2.n76 VDD2.n0 8.14595
R1896 VDD2.n151 VDD2.n150 7.3702
R1897 VDD2.n147 VDD2.n146 7.3702
R1898 VDD2.n105 VDD2.n102 7.3702
R1899 VDD2.n27 VDD2.n24 7.3702
R1900 VDD2.n70 VDD2.n69 7.3702
R1901 VDD2.n74 VDD2.n73 7.3702
R1902 VDD2.n150 VDD2.n79 6.59444
R1903 VDD2.n147 VDD2.n79 6.59444
R1904 VDD2.n70 VDD2.n2 6.59444
R1905 VDD2.n73 VDD2.n2 6.59444
R1906 VDD2.n151 VDD2.n77 5.81868
R1907 VDD2.n146 VDD2.n81 5.81868
R1908 VDD2.n106 VDD2.n105 5.81868
R1909 VDD2.n28 VDD2.n27 5.81868
R1910 VDD2.n69 VDD2.n4 5.81868
R1911 VDD2.n74 VDD2.n0 5.81868
R1912 VDD2.n143 VDD2.n142 5.04292
R1913 VDD2.n109 VDD2.n100 5.04292
R1914 VDD2.n31 VDD2.n22 5.04292
R1915 VDD2.n66 VDD2.n65 5.04292
R1916 VDD2.n139 VDD2.n83 4.26717
R1917 VDD2.n110 VDD2.n98 4.26717
R1918 VDD2.n32 VDD2.n20 4.26717
R1919 VDD2.n62 VDD2.n6 4.26717
R1920 VDD2.n138 VDD2.n85 3.49141
R1921 VDD2.n114 VDD2.n113 3.49141
R1922 VDD2.n36 VDD2.n35 3.49141
R1923 VDD2.n61 VDD2.n8 3.49141
R1924 VDD2.n135 VDD2.n134 2.71565
R1925 VDD2.n117 VDD2.n96 2.71565
R1926 VDD2.n39 VDD2.n18 2.71565
R1927 VDD2.n58 VDD2.n57 2.71565
R1928 VDD2.n104 VDD2.n103 2.41282
R1929 VDD2.n26 VDD2.n25 2.41282
R1930 VDD2.n131 VDD2.n87 1.93989
R1931 VDD2.n118 VDD2.n94 1.93989
R1932 VDD2.n40 VDD2.n16 1.93989
R1933 VDD2.n54 VDD2.n10 1.93989
R1934 VDD2.n130 VDD2.n89 1.16414
R1935 VDD2.n122 VDD2.n121 1.16414
R1936 VDD2.n45 VDD2.n43 1.16414
R1937 VDD2.n53 VDD2.n12 1.16414
R1938 VDD2 VDD2.n154 0.8755
R1939 VDD2.n127 VDD2.n126 0.388379
R1940 VDD2.n93 VDD2.n91 0.388379
R1941 VDD2.n44 VDD2.n14 0.388379
R1942 VDD2.n50 VDD2.n49 0.388379
R1943 VDD2.n152 VDD2.n78 0.155672
R1944 VDD2.n145 VDD2.n78 0.155672
R1945 VDD2.n145 VDD2.n144 0.155672
R1946 VDD2.n144 VDD2.n82 0.155672
R1947 VDD2.n137 VDD2.n82 0.155672
R1948 VDD2.n137 VDD2.n136 0.155672
R1949 VDD2.n136 VDD2.n86 0.155672
R1950 VDD2.n129 VDD2.n86 0.155672
R1951 VDD2.n129 VDD2.n128 0.155672
R1952 VDD2.n128 VDD2.n90 0.155672
R1953 VDD2.n120 VDD2.n90 0.155672
R1954 VDD2.n120 VDD2.n119 0.155672
R1955 VDD2.n119 VDD2.n95 0.155672
R1956 VDD2.n112 VDD2.n95 0.155672
R1957 VDD2.n112 VDD2.n111 0.155672
R1958 VDD2.n111 VDD2.n99 0.155672
R1959 VDD2.n104 VDD2.n99 0.155672
R1960 VDD2.n26 VDD2.n21 0.155672
R1961 VDD2.n33 VDD2.n21 0.155672
R1962 VDD2.n34 VDD2.n33 0.155672
R1963 VDD2.n34 VDD2.n17 0.155672
R1964 VDD2.n41 VDD2.n17 0.155672
R1965 VDD2.n42 VDD2.n41 0.155672
R1966 VDD2.n42 VDD2.n13 0.155672
R1967 VDD2.n51 VDD2.n13 0.155672
R1968 VDD2.n52 VDD2.n51 0.155672
R1969 VDD2.n52 VDD2.n9 0.155672
R1970 VDD2.n59 VDD2.n9 0.155672
R1971 VDD2.n60 VDD2.n59 0.155672
R1972 VDD2.n60 VDD2.n5 0.155672
R1973 VDD2.n67 VDD2.n5 0.155672
R1974 VDD2.n68 VDD2.n67 0.155672
R1975 VDD2.n68 VDD2.n1 0.155672
R1976 VDD2.n75 VDD2.n1 0.155672
C0 VDD1 VN 0.148851f
C1 VDD2 VN 3.386f
C2 w_n2486_n3820# VDD1 2.03331f
C3 w_n2486_n3820# VDD2 2.06985f
C4 VDD1 VP 3.60434f
C5 VP VDD2 0.369677f
C6 VN B 1.2255f
C7 VDD1 VTAIL 5.80119f
C8 VTAIL VDD2 5.85792f
C9 w_n2486_n3820# B 10.3716f
C10 VP B 1.75261f
C11 VTAIL B 4.50879f
C12 VDD1 VDD2 0.779832f
C13 VDD1 B 2.0012f
C14 w_n2486_n3820# VN 3.5528f
C15 VDD2 B 2.03894f
C16 VP VN 6.27369f
C17 w_n2486_n3820# VP 3.87132f
C18 VTAIL VN 3.00135f
C19 w_n2486_n3820# VTAIL 3.07315f
C20 VTAIL VP 3.01561f
C21 VDD2 VSUBS 1.09905f
C22 VDD1 VSUBS 5.44533f
C23 VTAIL VSUBS 1.179271f
C24 VN VSUBS 8.55391f
C25 VP VSUBS 2.021076f
C26 B VSUBS 4.731739f
C27 w_n2486_n3820# VSUBS 0.116554p
C28 VDD2.n0 VSUBS 0.033348f
C29 VDD2.n1 VSUBS 0.02933f
C30 VDD2.n2 VSUBS 0.015761f
C31 VDD2.n3 VSUBS 0.037253f
C32 VDD2.n4 VSUBS 0.016688f
C33 VDD2.n5 VSUBS 0.02933f
C34 VDD2.n6 VSUBS 0.015761f
C35 VDD2.n7 VSUBS 0.037253f
C36 VDD2.n8 VSUBS 0.016688f
C37 VDD2.n9 VSUBS 0.02933f
C38 VDD2.n10 VSUBS 0.015761f
C39 VDD2.n11 VSUBS 0.037253f
C40 VDD2.n12 VSUBS 0.016688f
C41 VDD2.n13 VSUBS 0.02933f
C42 VDD2.n14 VSUBS 0.016224f
C43 VDD2.n15 VSUBS 0.037253f
C44 VDD2.n16 VSUBS 0.016688f
C45 VDD2.n17 VSUBS 0.02933f
C46 VDD2.n18 VSUBS 0.015761f
C47 VDD2.n19 VSUBS 0.037253f
C48 VDD2.n20 VSUBS 0.016688f
C49 VDD2.n21 VSUBS 0.02933f
C50 VDD2.n22 VSUBS 0.015761f
C51 VDD2.n23 VSUBS 0.02794f
C52 VDD2.n24 VSUBS 0.028023f
C53 VDD2.t0 VSUBS 0.080496f
C54 VDD2.n25 VSUBS 0.260962f
C55 VDD2.n26 VSUBS 1.73154f
C56 VDD2.n27 VSUBS 0.015761f
C57 VDD2.n28 VSUBS 0.016688f
C58 VDD2.n29 VSUBS 0.037253f
C59 VDD2.n30 VSUBS 0.037253f
C60 VDD2.n31 VSUBS 0.016688f
C61 VDD2.n32 VSUBS 0.015761f
C62 VDD2.n33 VSUBS 0.02933f
C63 VDD2.n34 VSUBS 0.02933f
C64 VDD2.n35 VSUBS 0.015761f
C65 VDD2.n36 VSUBS 0.016688f
C66 VDD2.n37 VSUBS 0.037253f
C67 VDD2.n38 VSUBS 0.037253f
C68 VDD2.n39 VSUBS 0.016688f
C69 VDD2.n40 VSUBS 0.015761f
C70 VDD2.n41 VSUBS 0.02933f
C71 VDD2.n42 VSUBS 0.02933f
C72 VDD2.n43 VSUBS 0.015761f
C73 VDD2.n44 VSUBS 0.015761f
C74 VDD2.n45 VSUBS 0.016688f
C75 VDD2.n46 VSUBS 0.037253f
C76 VDD2.n47 VSUBS 0.037253f
C77 VDD2.n48 VSUBS 0.037253f
C78 VDD2.n49 VSUBS 0.016224f
C79 VDD2.n50 VSUBS 0.015761f
C80 VDD2.n51 VSUBS 0.02933f
C81 VDD2.n52 VSUBS 0.02933f
C82 VDD2.n53 VSUBS 0.015761f
C83 VDD2.n54 VSUBS 0.016688f
C84 VDD2.n55 VSUBS 0.037253f
C85 VDD2.n56 VSUBS 0.037253f
C86 VDD2.n57 VSUBS 0.016688f
C87 VDD2.n58 VSUBS 0.015761f
C88 VDD2.n59 VSUBS 0.02933f
C89 VDD2.n60 VSUBS 0.02933f
C90 VDD2.n61 VSUBS 0.015761f
C91 VDD2.n62 VSUBS 0.016688f
C92 VDD2.n63 VSUBS 0.037253f
C93 VDD2.n64 VSUBS 0.037253f
C94 VDD2.n65 VSUBS 0.016688f
C95 VDD2.n66 VSUBS 0.015761f
C96 VDD2.n67 VSUBS 0.02933f
C97 VDD2.n68 VSUBS 0.02933f
C98 VDD2.n69 VSUBS 0.015761f
C99 VDD2.n70 VSUBS 0.016688f
C100 VDD2.n71 VSUBS 0.037253f
C101 VDD2.n72 VSUBS 0.094002f
C102 VDD2.n73 VSUBS 0.016688f
C103 VDD2.n74 VSUBS 0.015761f
C104 VDD2.n75 VSUBS 0.066994f
C105 VDD2.n76 VSUBS 1.03361f
C106 VDD2.n77 VSUBS 0.033348f
C107 VDD2.n78 VSUBS 0.02933f
C108 VDD2.n79 VSUBS 0.015761f
C109 VDD2.n80 VSUBS 0.037253f
C110 VDD2.n81 VSUBS 0.016688f
C111 VDD2.n82 VSUBS 0.02933f
C112 VDD2.n83 VSUBS 0.015761f
C113 VDD2.n84 VSUBS 0.037253f
C114 VDD2.n85 VSUBS 0.016688f
C115 VDD2.n86 VSUBS 0.02933f
C116 VDD2.n87 VSUBS 0.015761f
C117 VDD2.n88 VSUBS 0.037253f
C118 VDD2.n89 VSUBS 0.016688f
C119 VDD2.n90 VSUBS 0.02933f
C120 VDD2.n91 VSUBS 0.016224f
C121 VDD2.n92 VSUBS 0.037253f
C122 VDD2.n93 VSUBS 0.015761f
C123 VDD2.n94 VSUBS 0.016688f
C124 VDD2.n95 VSUBS 0.02933f
C125 VDD2.n96 VSUBS 0.015761f
C126 VDD2.n97 VSUBS 0.037253f
C127 VDD2.n98 VSUBS 0.016688f
C128 VDD2.n99 VSUBS 0.02933f
C129 VDD2.n100 VSUBS 0.015761f
C130 VDD2.n101 VSUBS 0.02794f
C131 VDD2.n102 VSUBS 0.028023f
C132 VDD2.t1 VSUBS 0.080496f
C133 VDD2.n103 VSUBS 0.260962f
C134 VDD2.n104 VSUBS 1.73154f
C135 VDD2.n105 VSUBS 0.015761f
C136 VDD2.n106 VSUBS 0.016688f
C137 VDD2.n107 VSUBS 0.037253f
C138 VDD2.n108 VSUBS 0.037253f
C139 VDD2.n109 VSUBS 0.016688f
C140 VDD2.n110 VSUBS 0.015761f
C141 VDD2.n111 VSUBS 0.02933f
C142 VDD2.n112 VSUBS 0.02933f
C143 VDD2.n113 VSUBS 0.015761f
C144 VDD2.n114 VSUBS 0.016688f
C145 VDD2.n115 VSUBS 0.037253f
C146 VDD2.n116 VSUBS 0.037253f
C147 VDD2.n117 VSUBS 0.016688f
C148 VDD2.n118 VSUBS 0.015761f
C149 VDD2.n119 VSUBS 0.02933f
C150 VDD2.n120 VSUBS 0.02933f
C151 VDD2.n121 VSUBS 0.015761f
C152 VDD2.n122 VSUBS 0.016688f
C153 VDD2.n123 VSUBS 0.037253f
C154 VDD2.n124 VSUBS 0.037253f
C155 VDD2.n125 VSUBS 0.037253f
C156 VDD2.n126 VSUBS 0.016224f
C157 VDD2.n127 VSUBS 0.015761f
C158 VDD2.n128 VSUBS 0.02933f
C159 VDD2.n129 VSUBS 0.02933f
C160 VDD2.n130 VSUBS 0.015761f
C161 VDD2.n131 VSUBS 0.016688f
C162 VDD2.n132 VSUBS 0.037253f
C163 VDD2.n133 VSUBS 0.037253f
C164 VDD2.n134 VSUBS 0.016688f
C165 VDD2.n135 VSUBS 0.015761f
C166 VDD2.n136 VSUBS 0.02933f
C167 VDD2.n137 VSUBS 0.02933f
C168 VDD2.n138 VSUBS 0.015761f
C169 VDD2.n139 VSUBS 0.016688f
C170 VDD2.n140 VSUBS 0.037253f
C171 VDD2.n141 VSUBS 0.037253f
C172 VDD2.n142 VSUBS 0.016688f
C173 VDD2.n143 VSUBS 0.015761f
C174 VDD2.n144 VSUBS 0.02933f
C175 VDD2.n145 VSUBS 0.02933f
C176 VDD2.n146 VSUBS 0.015761f
C177 VDD2.n147 VSUBS 0.016688f
C178 VDD2.n148 VSUBS 0.037253f
C179 VDD2.n149 VSUBS 0.094002f
C180 VDD2.n150 VSUBS 0.016688f
C181 VDD2.n151 VSUBS 0.015761f
C182 VDD2.n152 VSUBS 0.066994f
C183 VDD2.n153 VSUBS 0.067676f
C184 VDD2.n154 VSUBS 4.04275f
C185 VN.t1 VSUBS 4.89296f
C186 VN.t0 VSUBS 5.7276f
C187 VDD1.n0 VSUBS 0.033081f
C188 VDD1.n1 VSUBS 0.029095f
C189 VDD1.n2 VSUBS 0.015634f
C190 VDD1.n3 VSUBS 0.036954f
C191 VDD1.n4 VSUBS 0.016554f
C192 VDD1.n5 VSUBS 0.029095f
C193 VDD1.n6 VSUBS 0.015634f
C194 VDD1.n7 VSUBS 0.036954f
C195 VDD1.n8 VSUBS 0.016554f
C196 VDD1.n9 VSUBS 0.029095f
C197 VDD1.n10 VSUBS 0.015634f
C198 VDD1.n11 VSUBS 0.036954f
C199 VDD1.n12 VSUBS 0.016554f
C200 VDD1.n13 VSUBS 0.029095f
C201 VDD1.n14 VSUBS 0.016094f
C202 VDD1.n15 VSUBS 0.036954f
C203 VDD1.n16 VSUBS 0.015634f
C204 VDD1.n17 VSUBS 0.016554f
C205 VDD1.n18 VSUBS 0.029095f
C206 VDD1.n19 VSUBS 0.015634f
C207 VDD1.n20 VSUBS 0.036954f
C208 VDD1.n21 VSUBS 0.016554f
C209 VDD1.n22 VSUBS 0.029095f
C210 VDD1.n23 VSUBS 0.015634f
C211 VDD1.n24 VSUBS 0.027716f
C212 VDD1.n25 VSUBS 0.027799f
C213 VDD1.t0 VSUBS 0.079851f
C214 VDD1.n26 VSUBS 0.258869f
C215 VDD1.n27 VSUBS 1.71765f
C216 VDD1.n28 VSUBS 0.015634f
C217 VDD1.n29 VSUBS 0.016554f
C218 VDD1.n30 VSUBS 0.036954f
C219 VDD1.n31 VSUBS 0.036954f
C220 VDD1.n32 VSUBS 0.016554f
C221 VDD1.n33 VSUBS 0.015634f
C222 VDD1.n34 VSUBS 0.029095f
C223 VDD1.n35 VSUBS 0.029095f
C224 VDD1.n36 VSUBS 0.015634f
C225 VDD1.n37 VSUBS 0.016554f
C226 VDD1.n38 VSUBS 0.036954f
C227 VDD1.n39 VSUBS 0.036954f
C228 VDD1.n40 VSUBS 0.016554f
C229 VDD1.n41 VSUBS 0.015634f
C230 VDD1.n42 VSUBS 0.029095f
C231 VDD1.n43 VSUBS 0.029095f
C232 VDD1.n44 VSUBS 0.015634f
C233 VDD1.n45 VSUBS 0.016554f
C234 VDD1.n46 VSUBS 0.036954f
C235 VDD1.n47 VSUBS 0.036954f
C236 VDD1.n48 VSUBS 0.036954f
C237 VDD1.n49 VSUBS 0.016094f
C238 VDD1.n50 VSUBS 0.015634f
C239 VDD1.n51 VSUBS 0.029095f
C240 VDD1.n52 VSUBS 0.029095f
C241 VDD1.n53 VSUBS 0.015634f
C242 VDD1.n54 VSUBS 0.016554f
C243 VDD1.n55 VSUBS 0.036954f
C244 VDD1.n56 VSUBS 0.036954f
C245 VDD1.n57 VSUBS 0.016554f
C246 VDD1.n58 VSUBS 0.015634f
C247 VDD1.n59 VSUBS 0.029095f
C248 VDD1.n60 VSUBS 0.029095f
C249 VDD1.n61 VSUBS 0.015634f
C250 VDD1.n62 VSUBS 0.016554f
C251 VDD1.n63 VSUBS 0.036954f
C252 VDD1.n64 VSUBS 0.036954f
C253 VDD1.n65 VSUBS 0.016554f
C254 VDD1.n66 VSUBS 0.015634f
C255 VDD1.n67 VSUBS 0.029095f
C256 VDD1.n68 VSUBS 0.029095f
C257 VDD1.n69 VSUBS 0.015634f
C258 VDD1.n70 VSUBS 0.016554f
C259 VDD1.n71 VSUBS 0.036954f
C260 VDD1.n72 VSUBS 0.093248f
C261 VDD1.n73 VSUBS 0.016554f
C262 VDD1.n74 VSUBS 0.015634f
C263 VDD1.n75 VSUBS 0.066457f
C264 VDD1.n76 VSUBS 0.069573f
C265 VDD1.n77 VSUBS 0.033081f
C266 VDD1.n78 VSUBS 0.029095f
C267 VDD1.n79 VSUBS 0.015634f
C268 VDD1.n80 VSUBS 0.036954f
C269 VDD1.n81 VSUBS 0.016554f
C270 VDD1.n82 VSUBS 0.029095f
C271 VDD1.n83 VSUBS 0.015634f
C272 VDD1.n84 VSUBS 0.036954f
C273 VDD1.n85 VSUBS 0.016554f
C274 VDD1.n86 VSUBS 0.029095f
C275 VDD1.n87 VSUBS 0.015634f
C276 VDD1.n88 VSUBS 0.036954f
C277 VDD1.n89 VSUBS 0.016554f
C278 VDD1.n90 VSUBS 0.029095f
C279 VDD1.n91 VSUBS 0.016094f
C280 VDD1.n92 VSUBS 0.036954f
C281 VDD1.n93 VSUBS 0.016554f
C282 VDD1.n94 VSUBS 0.029095f
C283 VDD1.n95 VSUBS 0.015634f
C284 VDD1.n96 VSUBS 0.036954f
C285 VDD1.n97 VSUBS 0.016554f
C286 VDD1.n98 VSUBS 0.029095f
C287 VDD1.n99 VSUBS 0.015634f
C288 VDD1.n100 VSUBS 0.027716f
C289 VDD1.n101 VSUBS 0.027799f
C290 VDD1.t1 VSUBS 0.079851f
C291 VDD1.n102 VSUBS 0.258869f
C292 VDD1.n103 VSUBS 1.71765f
C293 VDD1.n104 VSUBS 0.015634f
C294 VDD1.n105 VSUBS 0.016554f
C295 VDD1.n106 VSUBS 0.036954f
C296 VDD1.n107 VSUBS 0.036954f
C297 VDD1.n108 VSUBS 0.016554f
C298 VDD1.n109 VSUBS 0.015634f
C299 VDD1.n110 VSUBS 0.029095f
C300 VDD1.n111 VSUBS 0.029095f
C301 VDD1.n112 VSUBS 0.015634f
C302 VDD1.n113 VSUBS 0.016554f
C303 VDD1.n114 VSUBS 0.036954f
C304 VDD1.n115 VSUBS 0.036954f
C305 VDD1.n116 VSUBS 0.016554f
C306 VDD1.n117 VSUBS 0.015634f
C307 VDD1.n118 VSUBS 0.029095f
C308 VDD1.n119 VSUBS 0.029095f
C309 VDD1.n120 VSUBS 0.015634f
C310 VDD1.n121 VSUBS 0.015634f
C311 VDD1.n122 VSUBS 0.016554f
C312 VDD1.n123 VSUBS 0.036954f
C313 VDD1.n124 VSUBS 0.036954f
C314 VDD1.n125 VSUBS 0.036954f
C315 VDD1.n126 VSUBS 0.016094f
C316 VDD1.n127 VSUBS 0.015634f
C317 VDD1.n128 VSUBS 0.029095f
C318 VDD1.n129 VSUBS 0.029095f
C319 VDD1.n130 VSUBS 0.015634f
C320 VDD1.n131 VSUBS 0.016554f
C321 VDD1.n132 VSUBS 0.036954f
C322 VDD1.n133 VSUBS 0.036954f
C323 VDD1.n134 VSUBS 0.016554f
C324 VDD1.n135 VSUBS 0.015634f
C325 VDD1.n136 VSUBS 0.029095f
C326 VDD1.n137 VSUBS 0.029095f
C327 VDD1.n138 VSUBS 0.015634f
C328 VDD1.n139 VSUBS 0.016554f
C329 VDD1.n140 VSUBS 0.036954f
C330 VDD1.n141 VSUBS 0.036954f
C331 VDD1.n142 VSUBS 0.016554f
C332 VDD1.n143 VSUBS 0.015634f
C333 VDD1.n144 VSUBS 0.029095f
C334 VDD1.n145 VSUBS 0.029095f
C335 VDD1.n146 VSUBS 0.015634f
C336 VDD1.n147 VSUBS 0.016554f
C337 VDD1.n148 VSUBS 0.036954f
C338 VDD1.n149 VSUBS 0.093248f
C339 VDD1.n150 VSUBS 0.016554f
C340 VDD1.n151 VSUBS 0.015634f
C341 VDD1.n152 VSUBS 0.066457f
C342 VDD1.n153 VSUBS 1.09414f
C343 VTAIL.n0 VSUBS 0.033464f
C344 VTAIL.n1 VSUBS 0.029431f
C345 VTAIL.n2 VSUBS 0.015815f
C346 VTAIL.n3 VSUBS 0.037381f
C347 VTAIL.n4 VSUBS 0.016746f
C348 VTAIL.n5 VSUBS 0.029431f
C349 VTAIL.n6 VSUBS 0.015815f
C350 VTAIL.n7 VSUBS 0.037381f
C351 VTAIL.n8 VSUBS 0.016746f
C352 VTAIL.n9 VSUBS 0.029431f
C353 VTAIL.n10 VSUBS 0.015815f
C354 VTAIL.n11 VSUBS 0.037381f
C355 VTAIL.n12 VSUBS 0.016746f
C356 VTAIL.n13 VSUBS 0.029431f
C357 VTAIL.n14 VSUBS 0.01628f
C358 VTAIL.n15 VSUBS 0.037381f
C359 VTAIL.n16 VSUBS 0.016746f
C360 VTAIL.n17 VSUBS 0.029431f
C361 VTAIL.n18 VSUBS 0.015815f
C362 VTAIL.n19 VSUBS 0.037381f
C363 VTAIL.n20 VSUBS 0.016746f
C364 VTAIL.n21 VSUBS 0.029431f
C365 VTAIL.n22 VSUBS 0.015815f
C366 VTAIL.n23 VSUBS 0.028036f
C367 VTAIL.n24 VSUBS 0.02812f
C368 VTAIL.t2 VSUBS 0.080774f
C369 VTAIL.n25 VSUBS 0.261863f
C370 VTAIL.n26 VSUBS 1.73751f
C371 VTAIL.n27 VSUBS 0.015815f
C372 VTAIL.n28 VSUBS 0.016746f
C373 VTAIL.n29 VSUBS 0.037381f
C374 VTAIL.n30 VSUBS 0.037381f
C375 VTAIL.n31 VSUBS 0.016746f
C376 VTAIL.n32 VSUBS 0.015815f
C377 VTAIL.n33 VSUBS 0.029431f
C378 VTAIL.n34 VSUBS 0.029431f
C379 VTAIL.n35 VSUBS 0.015815f
C380 VTAIL.n36 VSUBS 0.016746f
C381 VTAIL.n37 VSUBS 0.037381f
C382 VTAIL.n38 VSUBS 0.037381f
C383 VTAIL.n39 VSUBS 0.016746f
C384 VTAIL.n40 VSUBS 0.015815f
C385 VTAIL.n41 VSUBS 0.029431f
C386 VTAIL.n42 VSUBS 0.029431f
C387 VTAIL.n43 VSUBS 0.015815f
C388 VTAIL.n44 VSUBS 0.015815f
C389 VTAIL.n45 VSUBS 0.016746f
C390 VTAIL.n46 VSUBS 0.037381f
C391 VTAIL.n47 VSUBS 0.037381f
C392 VTAIL.n48 VSUBS 0.037381f
C393 VTAIL.n49 VSUBS 0.01628f
C394 VTAIL.n50 VSUBS 0.015815f
C395 VTAIL.n51 VSUBS 0.029431f
C396 VTAIL.n52 VSUBS 0.029431f
C397 VTAIL.n53 VSUBS 0.015815f
C398 VTAIL.n54 VSUBS 0.016746f
C399 VTAIL.n55 VSUBS 0.037381f
C400 VTAIL.n56 VSUBS 0.037381f
C401 VTAIL.n57 VSUBS 0.016746f
C402 VTAIL.n58 VSUBS 0.015815f
C403 VTAIL.n59 VSUBS 0.029431f
C404 VTAIL.n60 VSUBS 0.029431f
C405 VTAIL.n61 VSUBS 0.015815f
C406 VTAIL.n62 VSUBS 0.016746f
C407 VTAIL.n63 VSUBS 0.037381f
C408 VTAIL.n64 VSUBS 0.037381f
C409 VTAIL.n65 VSUBS 0.016746f
C410 VTAIL.n66 VSUBS 0.015815f
C411 VTAIL.n67 VSUBS 0.029431f
C412 VTAIL.n68 VSUBS 0.029431f
C413 VTAIL.n69 VSUBS 0.015815f
C414 VTAIL.n70 VSUBS 0.016746f
C415 VTAIL.n71 VSUBS 0.037381f
C416 VTAIL.n72 VSUBS 0.094327f
C417 VTAIL.n73 VSUBS 0.016746f
C418 VTAIL.n74 VSUBS 0.015815f
C419 VTAIL.n75 VSUBS 0.067225f
C420 VTAIL.n76 VSUBS 0.047581f
C421 VTAIL.n77 VSUBS 2.33752f
C422 VTAIL.n78 VSUBS 0.033464f
C423 VTAIL.n79 VSUBS 0.029431f
C424 VTAIL.n80 VSUBS 0.015815f
C425 VTAIL.n81 VSUBS 0.037381f
C426 VTAIL.n82 VSUBS 0.016746f
C427 VTAIL.n83 VSUBS 0.029431f
C428 VTAIL.n84 VSUBS 0.015815f
C429 VTAIL.n85 VSUBS 0.037381f
C430 VTAIL.n86 VSUBS 0.016746f
C431 VTAIL.n87 VSUBS 0.029431f
C432 VTAIL.n88 VSUBS 0.015815f
C433 VTAIL.n89 VSUBS 0.037381f
C434 VTAIL.n90 VSUBS 0.016746f
C435 VTAIL.n91 VSUBS 0.029431f
C436 VTAIL.n92 VSUBS 0.01628f
C437 VTAIL.n93 VSUBS 0.037381f
C438 VTAIL.n94 VSUBS 0.015815f
C439 VTAIL.n95 VSUBS 0.016746f
C440 VTAIL.n96 VSUBS 0.029431f
C441 VTAIL.n97 VSUBS 0.015815f
C442 VTAIL.n98 VSUBS 0.037381f
C443 VTAIL.n99 VSUBS 0.016746f
C444 VTAIL.n100 VSUBS 0.029431f
C445 VTAIL.n101 VSUBS 0.015815f
C446 VTAIL.n102 VSUBS 0.028036f
C447 VTAIL.n103 VSUBS 0.02812f
C448 VTAIL.t0 VSUBS 0.080774f
C449 VTAIL.n104 VSUBS 0.261863f
C450 VTAIL.n105 VSUBS 1.73751f
C451 VTAIL.n106 VSUBS 0.015815f
C452 VTAIL.n107 VSUBS 0.016746f
C453 VTAIL.n108 VSUBS 0.037381f
C454 VTAIL.n109 VSUBS 0.037381f
C455 VTAIL.n110 VSUBS 0.016746f
C456 VTAIL.n111 VSUBS 0.015815f
C457 VTAIL.n112 VSUBS 0.029431f
C458 VTAIL.n113 VSUBS 0.029431f
C459 VTAIL.n114 VSUBS 0.015815f
C460 VTAIL.n115 VSUBS 0.016746f
C461 VTAIL.n116 VSUBS 0.037381f
C462 VTAIL.n117 VSUBS 0.037381f
C463 VTAIL.n118 VSUBS 0.016746f
C464 VTAIL.n119 VSUBS 0.015815f
C465 VTAIL.n120 VSUBS 0.029431f
C466 VTAIL.n121 VSUBS 0.029431f
C467 VTAIL.n122 VSUBS 0.015815f
C468 VTAIL.n123 VSUBS 0.016746f
C469 VTAIL.n124 VSUBS 0.037381f
C470 VTAIL.n125 VSUBS 0.037381f
C471 VTAIL.n126 VSUBS 0.037381f
C472 VTAIL.n127 VSUBS 0.01628f
C473 VTAIL.n128 VSUBS 0.015815f
C474 VTAIL.n129 VSUBS 0.029431f
C475 VTAIL.n130 VSUBS 0.029431f
C476 VTAIL.n131 VSUBS 0.015815f
C477 VTAIL.n132 VSUBS 0.016746f
C478 VTAIL.n133 VSUBS 0.037381f
C479 VTAIL.n134 VSUBS 0.037381f
C480 VTAIL.n135 VSUBS 0.016746f
C481 VTAIL.n136 VSUBS 0.015815f
C482 VTAIL.n137 VSUBS 0.029431f
C483 VTAIL.n138 VSUBS 0.029431f
C484 VTAIL.n139 VSUBS 0.015815f
C485 VTAIL.n140 VSUBS 0.016746f
C486 VTAIL.n141 VSUBS 0.037381f
C487 VTAIL.n142 VSUBS 0.037381f
C488 VTAIL.n143 VSUBS 0.016746f
C489 VTAIL.n144 VSUBS 0.015815f
C490 VTAIL.n145 VSUBS 0.029431f
C491 VTAIL.n146 VSUBS 0.029431f
C492 VTAIL.n147 VSUBS 0.015815f
C493 VTAIL.n148 VSUBS 0.016746f
C494 VTAIL.n149 VSUBS 0.037381f
C495 VTAIL.n150 VSUBS 0.094327f
C496 VTAIL.n151 VSUBS 0.016746f
C497 VTAIL.n152 VSUBS 0.015815f
C498 VTAIL.n153 VSUBS 0.067225f
C499 VTAIL.n154 VSUBS 0.047581f
C500 VTAIL.n155 VSUBS 2.40947f
C501 VTAIL.n156 VSUBS 0.033464f
C502 VTAIL.n157 VSUBS 0.029431f
C503 VTAIL.n158 VSUBS 0.015815f
C504 VTAIL.n159 VSUBS 0.037381f
C505 VTAIL.n160 VSUBS 0.016746f
C506 VTAIL.n161 VSUBS 0.029431f
C507 VTAIL.n162 VSUBS 0.015815f
C508 VTAIL.n163 VSUBS 0.037381f
C509 VTAIL.n164 VSUBS 0.016746f
C510 VTAIL.n165 VSUBS 0.029431f
C511 VTAIL.n166 VSUBS 0.015815f
C512 VTAIL.n167 VSUBS 0.037381f
C513 VTAIL.n168 VSUBS 0.016746f
C514 VTAIL.n169 VSUBS 0.029431f
C515 VTAIL.n170 VSUBS 0.01628f
C516 VTAIL.n171 VSUBS 0.037381f
C517 VTAIL.n172 VSUBS 0.015815f
C518 VTAIL.n173 VSUBS 0.016746f
C519 VTAIL.n174 VSUBS 0.029431f
C520 VTAIL.n175 VSUBS 0.015815f
C521 VTAIL.n176 VSUBS 0.037381f
C522 VTAIL.n177 VSUBS 0.016746f
C523 VTAIL.n178 VSUBS 0.029431f
C524 VTAIL.n179 VSUBS 0.015815f
C525 VTAIL.n180 VSUBS 0.028036f
C526 VTAIL.n181 VSUBS 0.02812f
C527 VTAIL.t3 VSUBS 0.080774f
C528 VTAIL.n182 VSUBS 0.261863f
C529 VTAIL.n183 VSUBS 1.73751f
C530 VTAIL.n184 VSUBS 0.015815f
C531 VTAIL.n185 VSUBS 0.016746f
C532 VTAIL.n186 VSUBS 0.037381f
C533 VTAIL.n187 VSUBS 0.037381f
C534 VTAIL.n188 VSUBS 0.016746f
C535 VTAIL.n189 VSUBS 0.015815f
C536 VTAIL.n190 VSUBS 0.029431f
C537 VTAIL.n191 VSUBS 0.029431f
C538 VTAIL.n192 VSUBS 0.015815f
C539 VTAIL.n193 VSUBS 0.016746f
C540 VTAIL.n194 VSUBS 0.037381f
C541 VTAIL.n195 VSUBS 0.037381f
C542 VTAIL.n196 VSUBS 0.016746f
C543 VTAIL.n197 VSUBS 0.015815f
C544 VTAIL.n198 VSUBS 0.029431f
C545 VTAIL.n199 VSUBS 0.029431f
C546 VTAIL.n200 VSUBS 0.015815f
C547 VTAIL.n201 VSUBS 0.016746f
C548 VTAIL.n202 VSUBS 0.037381f
C549 VTAIL.n203 VSUBS 0.037381f
C550 VTAIL.n204 VSUBS 0.037381f
C551 VTAIL.n205 VSUBS 0.01628f
C552 VTAIL.n206 VSUBS 0.015815f
C553 VTAIL.n207 VSUBS 0.029431f
C554 VTAIL.n208 VSUBS 0.029431f
C555 VTAIL.n209 VSUBS 0.015815f
C556 VTAIL.n210 VSUBS 0.016746f
C557 VTAIL.n211 VSUBS 0.037381f
C558 VTAIL.n212 VSUBS 0.037381f
C559 VTAIL.n213 VSUBS 0.016746f
C560 VTAIL.n214 VSUBS 0.015815f
C561 VTAIL.n215 VSUBS 0.029431f
C562 VTAIL.n216 VSUBS 0.029431f
C563 VTAIL.n217 VSUBS 0.015815f
C564 VTAIL.n218 VSUBS 0.016746f
C565 VTAIL.n219 VSUBS 0.037381f
C566 VTAIL.n220 VSUBS 0.037381f
C567 VTAIL.n221 VSUBS 0.016746f
C568 VTAIL.n222 VSUBS 0.015815f
C569 VTAIL.n223 VSUBS 0.029431f
C570 VTAIL.n224 VSUBS 0.029431f
C571 VTAIL.n225 VSUBS 0.015815f
C572 VTAIL.n226 VSUBS 0.016746f
C573 VTAIL.n227 VSUBS 0.037381f
C574 VTAIL.n228 VSUBS 0.094327f
C575 VTAIL.n229 VSUBS 0.016746f
C576 VTAIL.n230 VSUBS 0.015815f
C577 VTAIL.n231 VSUBS 0.067225f
C578 VTAIL.n232 VSUBS 0.047581f
C579 VTAIL.n233 VSUBS 2.09962f
C580 VTAIL.n234 VSUBS 0.033464f
C581 VTAIL.n235 VSUBS 0.029431f
C582 VTAIL.n236 VSUBS 0.015815f
C583 VTAIL.n237 VSUBS 0.037381f
C584 VTAIL.n238 VSUBS 0.016746f
C585 VTAIL.n239 VSUBS 0.029431f
C586 VTAIL.n240 VSUBS 0.015815f
C587 VTAIL.n241 VSUBS 0.037381f
C588 VTAIL.n242 VSUBS 0.016746f
C589 VTAIL.n243 VSUBS 0.029431f
C590 VTAIL.n244 VSUBS 0.015815f
C591 VTAIL.n245 VSUBS 0.037381f
C592 VTAIL.n246 VSUBS 0.016746f
C593 VTAIL.n247 VSUBS 0.029431f
C594 VTAIL.n248 VSUBS 0.01628f
C595 VTAIL.n249 VSUBS 0.037381f
C596 VTAIL.n250 VSUBS 0.016746f
C597 VTAIL.n251 VSUBS 0.029431f
C598 VTAIL.n252 VSUBS 0.015815f
C599 VTAIL.n253 VSUBS 0.037381f
C600 VTAIL.n254 VSUBS 0.016746f
C601 VTAIL.n255 VSUBS 0.029431f
C602 VTAIL.n256 VSUBS 0.015815f
C603 VTAIL.n257 VSUBS 0.028036f
C604 VTAIL.n258 VSUBS 0.02812f
C605 VTAIL.t1 VSUBS 0.080774f
C606 VTAIL.n259 VSUBS 0.261863f
C607 VTAIL.n260 VSUBS 1.73751f
C608 VTAIL.n261 VSUBS 0.015815f
C609 VTAIL.n262 VSUBS 0.016746f
C610 VTAIL.n263 VSUBS 0.037381f
C611 VTAIL.n264 VSUBS 0.037381f
C612 VTAIL.n265 VSUBS 0.016746f
C613 VTAIL.n266 VSUBS 0.015815f
C614 VTAIL.n267 VSUBS 0.029431f
C615 VTAIL.n268 VSUBS 0.029431f
C616 VTAIL.n269 VSUBS 0.015815f
C617 VTAIL.n270 VSUBS 0.016746f
C618 VTAIL.n271 VSUBS 0.037381f
C619 VTAIL.n272 VSUBS 0.037381f
C620 VTAIL.n273 VSUBS 0.016746f
C621 VTAIL.n274 VSUBS 0.015815f
C622 VTAIL.n275 VSUBS 0.029431f
C623 VTAIL.n276 VSUBS 0.029431f
C624 VTAIL.n277 VSUBS 0.015815f
C625 VTAIL.n278 VSUBS 0.015815f
C626 VTAIL.n279 VSUBS 0.016746f
C627 VTAIL.n280 VSUBS 0.037381f
C628 VTAIL.n281 VSUBS 0.037381f
C629 VTAIL.n282 VSUBS 0.037381f
C630 VTAIL.n283 VSUBS 0.01628f
C631 VTAIL.n284 VSUBS 0.015815f
C632 VTAIL.n285 VSUBS 0.029431f
C633 VTAIL.n286 VSUBS 0.029431f
C634 VTAIL.n287 VSUBS 0.015815f
C635 VTAIL.n288 VSUBS 0.016746f
C636 VTAIL.n289 VSUBS 0.037381f
C637 VTAIL.n290 VSUBS 0.037381f
C638 VTAIL.n291 VSUBS 0.016746f
C639 VTAIL.n292 VSUBS 0.015815f
C640 VTAIL.n293 VSUBS 0.029431f
C641 VTAIL.n294 VSUBS 0.029431f
C642 VTAIL.n295 VSUBS 0.015815f
C643 VTAIL.n296 VSUBS 0.016746f
C644 VTAIL.n297 VSUBS 0.037381f
C645 VTAIL.n298 VSUBS 0.037381f
C646 VTAIL.n299 VSUBS 0.016746f
C647 VTAIL.n300 VSUBS 0.015815f
C648 VTAIL.n301 VSUBS 0.029431f
C649 VTAIL.n302 VSUBS 0.029431f
C650 VTAIL.n303 VSUBS 0.015815f
C651 VTAIL.n304 VSUBS 0.016746f
C652 VTAIL.n305 VSUBS 0.037381f
C653 VTAIL.n306 VSUBS 0.094327f
C654 VTAIL.n307 VSUBS 0.016746f
C655 VTAIL.n308 VSUBS 0.015815f
C656 VTAIL.n309 VSUBS 0.067225f
C657 VTAIL.n310 VSUBS 0.047581f
C658 VTAIL.n311 VSUBS 1.97208f
C659 VP.t1 VSUBS 5.9201f
C660 VP.t0 VSUBS 5.05131f
C661 VP.n0 VSUBS 5.70485f
C662 B.n0 VSUBS 0.006043f
C663 B.n1 VSUBS 0.006043f
C664 B.n2 VSUBS 0.008937f
C665 B.n3 VSUBS 0.006849f
C666 B.n4 VSUBS 0.006849f
C667 B.n5 VSUBS 0.006849f
C668 B.n6 VSUBS 0.006849f
C669 B.n7 VSUBS 0.006849f
C670 B.n8 VSUBS 0.006849f
C671 B.n9 VSUBS 0.006849f
C672 B.n10 VSUBS 0.006849f
C673 B.n11 VSUBS 0.006849f
C674 B.n12 VSUBS 0.006849f
C675 B.n13 VSUBS 0.006849f
C676 B.n14 VSUBS 0.006849f
C677 B.n15 VSUBS 0.006849f
C678 B.n16 VSUBS 0.006849f
C679 B.n17 VSUBS 0.016105f
C680 B.n18 VSUBS 0.006849f
C681 B.n19 VSUBS 0.006849f
C682 B.n20 VSUBS 0.006849f
C683 B.n21 VSUBS 0.006849f
C684 B.n22 VSUBS 0.006849f
C685 B.n23 VSUBS 0.006849f
C686 B.n24 VSUBS 0.006849f
C687 B.n25 VSUBS 0.006849f
C688 B.n26 VSUBS 0.006849f
C689 B.n27 VSUBS 0.006849f
C690 B.n28 VSUBS 0.006849f
C691 B.n29 VSUBS 0.006849f
C692 B.n30 VSUBS 0.006849f
C693 B.n31 VSUBS 0.006849f
C694 B.n32 VSUBS 0.006849f
C695 B.n33 VSUBS 0.006849f
C696 B.n34 VSUBS 0.006849f
C697 B.n35 VSUBS 0.006849f
C698 B.n36 VSUBS 0.006849f
C699 B.n37 VSUBS 0.006849f
C700 B.n38 VSUBS 0.006849f
C701 B.n39 VSUBS 0.006849f
C702 B.n40 VSUBS 0.006849f
C703 B.n41 VSUBS 0.006849f
C704 B.t7 VSUBS 0.256955f
C705 B.t8 VSUBS 0.297389f
C706 B.t6 VSUBS 2.21731f
C707 B.n42 VSUBS 0.472017f
C708 B.n43 VSUBS 0.279344f
C709 B.n44 VSUBS 0.006849f
C710 B.n45 VSUBS 0.006849f
C711 B.n46 VSUBS 0.006849f
C712 B.n47 VSUBS 0.006849f
C713 B.t10 VSUBS 0.256958f
C714 B.t11 VSUBS 0.297392f
C715 B.t9 VSUBS 2.21731f
C716 B.n48 VSUBS 0.472015f
C717 B.n49 VSUBS 0.279341f
C718 B.n50 VSUBS 0.015868f
C719 B.n51 VSUBS 0.006849f
C720 B.n52 VSUBS 0.006849f
C721 B.n53 VSUBS 0.006849f
C722 B.n54 VSUBS 0.006849f
C723 B.n55 VSUBS 0.006849f
C724 B.n56 VSUBS 0.006849f
C725 B.n57 VSUBS 0.006849f
C726 B.n58 VSUBS 0.006849f
C727 B.n59 VSUBS 0.006849f
C728 B.n60 VSUBS 0.006849f
C729 B.n61 VSUBS 0.006849f
C730 B.n62 VSUBS 0.006849f
C731 B.n63 VSUBS 0.006849f
C732 B.n64 VSUBS 0.006849f
C733 B.n65 VSUBS 0.006849f
C734 B.n66 VSUBS 0.006849f
C735 B.n67 VSUBS 0.006849f
C736 B.n68 VSUBS 0.006849f
C737 B.n69 VSUBS 0.006849f
C738 B.n70 VSUBS 0.006849f
C739 B.n71 VSUBS 0.006849f
C740 B.n72 VSUBS 0.006849f
C741 B.n73 VSUBS 0.006849f
C742 B.n74 VSUBS 0.016105f
C743 B.n75 VSUBS 0.006849f
C744 B.n76 VSUBS 0.006849f
C745 B.n77 VSUBS 0.006849f
C746 B.n78 VSUBS 0.006849f
C747 B.n79 VSUBS 0.006849f
C748 B.n80 VSUBS 0.006849f
C749 B.n81 VSUBS 0.006849f
C750 B.n82 VSUBS 0.006849f
C751 B.n83 VSUBS 0.006849f
C752 B.n84 VSUBS 0.006849f
C753 B.n85 VSUBS 0.006849f
C754 B.n86 VSUBS 0.006849f
C755 B.n87 VSUBS 0.006849f
C756 B.n88 VSUBS 0.006849f
C757 B.n89 VSUBS 0.006849f
C758 B.n90 VSUBS 0.006849f
C759 B.n91 VSUBS 0.006849f
C760 B.n92 VSUBS 0.006849f
C761 B.n93 VSUBS 0.006849f
C762 B.n94 VSUBS 0.006849f
C763 B.n95 VSUBS 0.006849f
C764 B.n96 VSUBS 0.006849f
C765 B.n97 VSUBS 0.006849f
C766 B.n98 VSUBS 0.006849f
C767 B.n99 VSUBS 0.006849f
C768 B.n100 VSUBS 0.006849f
C769 B.n101 VSUBS 0.006849f
C770 B.n102 VSUBS 0.006849f
C771 B.n103 VSUBS 0.006849f
C772 B.n104 VSUBS 0.006849f
C773 B.n105 VSUBS 0.015521f
C774 B.n106 VSUBS 0.006849f
C775 B.n107 VSUBS 0.006849f
C776 B.n108 VSUBS 0.006849f
C777 B.n109 VSUBS 0.006849f
C778 B.n110 VSUBS 0.006849f
C779 B.n111 VSUBS 0.006849f
C780 B.n112 VSUBS 0.006849f
C781 B.n113 VSUBS 0.006849f
C782 B.n114 VSUBS 0.006849f
C783 B.n115 VSUBS 0.006849f
C784 B.n116 VSUBS 0.006849f
C785 B.n117 VSUBS 0.006849f
C786 B.n118 VSUBS 0.006849f
C787 B.n119 VSUBS 0.006849f
C788 B.n120 VSUBS 0.006849f
C789 B.n121 VSUBS 0.006849f
C790 B.n122 VSUBS 0.006849f
C791 B.n123 VSUBS 0.006849f
C792 B.n124 VSUBS 0.006849f
C793 B.n125 VSUBS 0.006849f
C794 B.n126 VSUBS 0.006849f
C795 B.n127 VSUBS 0.006849f
C796 B.n128 VSUBS 0.006849f
C797 B.n129 VSUBS 0.006849f
C798 B.t2 VSUBS 0.256958f
C799 B.t1 VSUBS 0.297392f
C800 B.t0 VSUBS 2.21731f
C801 B.n130 VSUBS 0.472015f
C802 B.n131 VSUBS 0.279341f
C803 B.n132 VSUBS 0.006849f
C804 B.n133 VSUBS 0.006849f
C805 B.n134 VSUBS 0.006849f
C806 B.n135 VSUBS 0.006849f
C807 B.n136 VSUBS 0.003827f
C808 B.n137 VSUBS 0.006849f
C809 B.n138 VSUBS 0.006849f
C810 B.n139 VSUBS 0.006849f
C811 B.n140 VSUBS 0.006849f
C812 B.n141 VSUBS 0.006849f
C813 B.n142 VSUBS 0.006849f
C814 B.n143 VSUBS 0.006849f
C815 B.n144 VSUBS 0.006849f
C816 B.n145 VSUBS 0.006849f
C817 B.n146 VSUBS 0.006849f
C818 B.n147 VSUBS 0.006849f
C819 B.n148 VSUBS 0.006849f
C820 B.n149 VSUBS 0.006849f
C821 B.n150 VSUBS 0.006849f
C822 B.n151 VSUBS 0.006849f
C823 B.n152 VSUBS 0.006849f
C824 B.n153 VSUBS 0.006849f
C825 B.n154 VSUBS 0.006849f
C826 B.n155 VSUBS 0.006849f
C827 B.n156 VSUBS 0.006849f
C828 B.n157 VSUBS 0.006849f
C829 B.n158 VSUBS 0.006849f
C830 B.n159 VSUBS 0.006849f
C831 B.n160 VSUBS 0.016105f
C832 B.n161 VSUBS 0.006849f
C833 B.n162 VSUBS 0.006849f
C834 B.n163 VSUBS 0.006849f
C835 B.n164 VSUBS 0.006849f
C836 B.n165 VSUBS 0.006849f
C837 B.n166 VSUBS 0.006849f
C838 B.n167 VSUBS 0.006849f
C839 B.n168 VSUBS 0.006849f
C840 B.n169 VSUBS 0.006849f
C841 B.n170 VSUBS 0.006849f
C842 B.n171 VSUBS 0.006849f
C843 B.n172 VSUBS 0.006849f
C844 B.n173 VSUBS 0.006849f
C845 B.n174 VSUBS 0.006849f
C846 B.n175 VSUBS 0.006849f
C847 B.n176 VSUBS 0.006849f
C848 B.n177 VSUBS 0.006849f
C849 B.n178 VSUBS 0.006849f
C850 B.n179 VSUBS 0.006849f
C851 B.n180 VSUBS 0.006849f
C852 B.n181 VSUBS 0.006849f
C853 B.n182 VSUBS 0.006849f
C854 B.n183 VSUBS 0.006849f
C855 B.n184 VSUBS 0.006849f
C856 B.n185 VSUBS 0.006849f
C857 B.n186 VSUBS 0.006849f
C858 B.n187 VSUBS 0.006849f
C859 B.n188 VSUBS 0.006849f
C860 B.n189 VSUBS 0.006849f
C861 B.n190 VSUBS 0.006849f
C862 B.n191 VSUBS 0.006849f
C863 B.n192 VSUBS 0.006849f
C864 B.n193 VSUBS 0.006849f
C865 B.n194 VSUBS 0.006849f
C866 B.n195 VSUBS 0.006849f
C867 B.n196 VSUBS 0.006849f
C868 B.n197 VSUBS 0.006849f
C869 B.n198 VSUBS 0.006849f
C870 B.n199 VSUBS 0.006849f
C871 B.n200 VSUBS 0.006849f
C872 B.n201 VSUBS 0.006849f
C873 B.n202 VSUBS 0.006849f
C874 B.n203 VSUBS 0.006849f
C875 B.n204 VSUBS 0.006849f
C876 B.n205 VSUBS 0.006849f
C877 B.n206 VSUBS 0.006849f
C878 B.n207 VSUBS 0.006849f
C879 B.n208 VSUBS 0.006849f
C880 B.n209 VSUBS 0.006849f
C881 B.n210 VSUBS 0.006849f
C882 B.n211 VSUBS 0.006849f
C883 B.n212 VSUBS 0.006849f
C884 B.n213 VSUBS 0.006849f
C885 B.n214 VSUBS 0.006849f
C886 B.n215 VSUBS 0.006849f
C887 B.n216 VSUBS 0.006849f
C888 B.n217 VSUBS 0.015521f
C889 B.n218 VSUBS 0.015521f
C890 B.n219 VSUBS 0.016105f
C891 B.n220 VSUBS 0.006849f
C892 B.n221 VSUBS 0.006849f
C893 B.n222 VSUBS 0.006849f
C894 B.n223 VSUBS 0.006849f
C895 B.n224 VSUBS 0.006849f
C896 B.n225 VSUBS 0.006849f
C897 B.n226 VSUBS 0.006849f
C898 B.n227 VSUBS 0.006849f
C899 B.n228 VSUBS 0.006849f
C900 B.n229 VSUBS 0.006849f
C901 B.n230 VSUBS 0.006849f
C902 B.n231 VSUBS 0.006849f
C903 B.n232 VSUBS 0.006849f
C904 B.n233 VSUBS 0.006849f
C905 B.n234 VSUBS 0.006849f
C906 B.n235 VSUBS 0.006849f
C907 B.n236 VSUBS 0.006849f
C908 B.n237 VSUBS 0.006849f
C909 B.n238 VSUBS 0.006849f
C910 B.n239 VSUBS 0.006849f
C911 B.n240 VSUBS 0.006849f
C912 B.n241 VSUBS 0.006849f
C913 B.n242 VSUBS 0.006849f
C914 B.n243 VSUBS 0.006849f
C915 B.n244 VSUBS 0.006849f
C916 B.n245 VSUBS 0.006849f
C917 B.n246 VSUBS 0.006849f
C918 B.n247 VSUBS 0.006849f
C919 B.n248 VSUBS 0.006849f
C920 B.n249 VSUBS 0.006849f
C921 B.n250 VSUBS 0.006849f
C922 B.n251 VSUBS 0.006849f
C923 B.n252 VSUBS 0.006849f
C924 B.n253 VSUBS 0.006849f
C925 B.n254 VSUBS 0.006849f
C926 B.n255 VSUBS 0.006849f
C927 B.n256 VSUBS 0.006849f
C928 B.n257 VSUBS 0.006849f
C929 B.n258 VSUBS 0.006849f
C930 B.n259 VSUBS 0.006849f
C931 B.n260 VSUBS 0.006849f
C932 B.n261 VSUBS 0.006849f
C933 B.n262 VSUBS 0.006849f
C934 B.n263 VSUBS 0.006849f
C935 B.n264 VSUBS 0.006849f
C936 B.n265 VSUBS 0.006849f
C937 B.n266 VSUBS 0.006849f
C938 B.n267 VSUBS 0.006849f
C939 B.n268 VSUBS 0.006849f
C940 B.n269 VSUBS 0.006849f
C941 B.n270 VSUBS 0.006849f
C942 B.n271 VSUBS 0.006849f
C943 B.n272 VSUBS 0.006849f
C944 B.n273 VSUBS 0.006849f
C945 B.n274 VSUBS 0.006849f
C946 B.n275 VSUBS 0.006849f
C947 B.n276 VSUBS 0.006849f
C948 B.n277 VSUBS 0.006849f
C949 B.n278 VSUBS 0.006849f
C950 B.n279 VSUBS 0.006849f
C951 B.n280 VSUBS 0.006849f
C952 B.n281 VSUBS 0.006849f
C953 B.n282 VSUBS 0.006849f
C954 B.n283 VSUBS 0.006849f
C955 B.n284 VSUBS 0.006849f
C956 B.n285 VSUBS 0.006849f
C957 B.n286 VSUBS 0.006849f
C958 B.n287 VSUBS 0.006849f
C959 B.n288 VSUBS 0.006849f
C960 B.t5 VSUBS 0.256955f
C961 B.t4 VSUBS 0.297389f
C962 B.t3 VSUBS 2.21731f
C963 B.n289 VSUBS 0.472017f
C964 B.n290 VSUBS 0.279344f
C965 B.n291 VSUBS 0.015868f
C966 B.n292 VSUBS 0.006446f
C967 B.n293 VSUBS 0.006849f
C968 B.n294 VSUBS 0.006849f
C969 B.n295 VSUBS 0.006849f
C970 B.n296 VSUBS 0.006849f
C971 B.n297 VSUBS 0.006849f
C972 B.n298 VSUBS 0.006849f
C973 B.n299 VSUBS 0.006849f
C974 B.n300 VSUBS 0.006849f
C975 B.n301 VSUBS 0.006849f
C976 B.n302 VSUBS 0.006849f
C977 B.n303 VSUBS 0.006849f
C978 B.n304 VSUBS 0.006849f
C979 B.n305 VSUBS 0.006849f
C980 B.n306 VSUBS 0.006849f
C981 B.n307 VSUBS 0.006849f
C982 B.n308 VSUBS 0.003827f
C983 B.n309 VSUBS 0.015868f
C984 B.n310 VSUBS 0.006446f
C985 B.n311 VSUBS 0.006849f
C986 B.n312 VSUBS 0.006849f
C987 B.n313 VSUBS 0.006849f
C988 B.n314 VSUBS 0.006849f
C989 B.n315 VSUBS 0.006849f
C990 B.n316 VSUBS 0.006849f
C991 B.n317 VSUBS 0.006849f
C992 B.n318 VSUBS 0.006849f
C993 B.n319 VSUBS 0.006849f
C994 B.n320 VSUBS 0.006849f
C995 B.n321 VSUBS 0.006849f
C996 B.n322 VSUBS 0.006849f
C997 B.n323 VSUBS 0.006849f
C998 B.n324 VSUBS 0.006849f
C999 B.n325 VSUBS 0.006849f
C1000 B.n326 VSUBS 0.006849f
C1001 B.n327 VSUBS 0.006849f
C1002 B.n328 VSUBS 0.006849f
C1003 B.n329 VSUBS 0.006849f
C1004 B.n330 VSUBS 0.006849f
C1005 B.n331 VSUBS 0.006849f
C1006 B.n332 VSUBS 0.006849f
C1007 B.n333 VSUBS 0.006849f
C1008 B.n334 VSUBS 0.006849f
C1009 B.n335 VSUBS 0.006849f
C1010 B.n336 VSUBS 0.006849f
C1011 B.n337 VSUBS 0.006849f
C1012 B.n338 VSUBS 0.006849f
C1013 B.n339 VSUBS 0.006849f
C1014 B.n340 VSUBS 0.006849f
C1015 B.n341 VSUBS 0.006849f
C1016 B.n342 VSUBS 0.006849f
C1017 B.n343 VSUBS 0.006849f
C1018 B.n344 VSUBS 0.006849f
C1019 B.n345 VSUBS 0.006849f
C1020 B.n346 VSUBS 0.006849f
C1021 B.n347 VSUBS 0.006849f
C1022 B.n348 VSUBS 0.006849f
C1023 B.n349 VSUBS 0.006849f
C1024 B.n350 VSUBS 0.006849f
C1025 B.n351 VSUBS 0.006849f
C1026 B.n352 VSUBS 0.006849f
C1027 B.n353 VSUBS 0.006849f
C1028 B.n354 VSUBS 0.006849f
C1029 B.n355 VSUBS 0.006849f
C1030 B.n356 VSUBS 0.006849f
C1031 B.n357 VSUBS 0.006849f
C1032 B.n358 VSUBS 0.006849f
C1033 B.n359 VSUBS 0.006849f
C1034 B.n360 VSUBS 0.006849f
C1035 B.n361 VSUBS 0.006849f
C1036 B.n362 VSUBS 0.006849f
C1037 B.n363 VSUBS 0.006849f
C1038 B.n364 VSUBS 0.006849f
C1039 B.n365 VSUBS 0.006849f
C1040 B.n366 VSUBS 0.006849f
C1041 B.n367 VSUBS 0.006849f
C1042 B.n368 VSUBS 0.006849f
C1043 B.n369 VSUBS 0.006849f
C1044 B.n370 VSUBS 0.006849f
C1045 B.n371 VSUBS 0.006849f
C1046 B.n372 VSUBS 0.006849f
C1047 B.n373 VSUBS 0.006849f
C1048 B.n374 VSUBS 0.006849f
C1049 B.n375 VSUBS 0.006849f
C1050 B.n376 VSUBS 0.006849f
C1051 B.n377 VSUBS 0.006849f
C1052 B.n378 VSUBS 0.006849f
C1053 B.n379 VSUBS 0.006849f
C1054 B.n380 VSUBS 0.016105f
C1055 B.n381 VSUBS 0.015279f
C1056 B.n382 VSUBS 0.016347f
C1057 B.n383 VSUBS 0.006849f
C1058 B.n384 VSUBS 0.006849f
C1059 B.n385 VSUBS 0.006849f
C1060 B.n386 VSUBS 0.006849f
C1061 B.n387 VSUBS 0.006849f
C1062 B.n388 VSUBS 0.006849f
C1063 B.n389 VSUBS 0.006849f
C1064 B.n390 VSUBS 0.006849f
C1065 B.n391 VSUBS 0.006849f
C1066 B.n392 VSUBS 0.006849f
C1067 B.n393 VSUBS 0.006849f
C1068 B.n394 VSUBS 0.006849f
C1069 B.n395 VSUBS 0.006849f
C1070 B.n396 VSUBS 0.006849f
C1071 B.n397 VSUBS 0.006849f
C1072 B.n398 VSUBS 0.006849f
C1073 B.n399 VSUBS 0.006849f
C1074 B.n400 VSUBS 0.006849f
C1075 B.n401 VSUBS 0.006849f
C1076 B.n402 VSUBS 0.006849f
C1077 B.n403 VSUBS 0.006849f
C1078 B.n404 VSUBS 0.006849f
C1079 B.n405 VSUBS 0.006849f
C1080 B.n406 VSUBS 0.006849f
C1081 B.n407 VSUBS 0.006849f
C1082 B.n408 VSUBS 0.006849f
C1083 B.n409 VSUBS 0.006849f
C1084 B.n410 VSUBS 0.006849f
C1085 B.n411 VSUBS 0.006849f
C1086 B.n412 VSUBS 0.006849f
C1087 B.n413 VSUBS 0.006849f
C1088 B.n414 VSUBS 0.006849f
C1089 B.n415 VSUBS 0.006849f
C1090 B.n416 VSUBS 0.006849f
C1091 B.n417 VSUBS 0.006849f
C1092 B.n418 VSUBS 0.006849f
C1093 B.n419 VSUBS 0.006849f
C1094 B.n420 VSUBS 0.006849f
C1095 B.n421 VSUBS 0.006849f
C1096 B.n422 VSUBS 0.006849f
C1097 B.n423 VSUBS 0.006849f
C1098 B.n424 VSUBS 0.006849f
C1099 B.n425 VSUBS 0.006849f
C1100 B.n426 VSUBS 0.006849f
C1101 B.n427 VSUBS 0.006849f
C1102 B.n428 VSUBS 0.006849f
C1103 B.n429 VSUBS 0.006849f
C1104 B.n430 VSUBS 0.006849f
C1105 B.n431 VSUBS 0.006849f
C1106 B.n432 VSUBS 0.006849f
C1107 B.n433 VSUBS 0.006849f
C1108 B.n434 VSUBS 0.006849f
C1109 B.n435 VSUBS 0.006849f
C1110 B.n436 VSUBS 0.006849f
C1111 B.n437 VSUBS 0.006849f
C1112 B.n438 VSUBS 0.006849f
C1113 B.n439 VSUBS 0.006849f
C1114 B.n440 VSUBS 0.006849f
C1115 B.n441 VSUBS 0.006849f
C1116 B.n442 VSUBS 0.006849f
C1117 B.n443 VSUBS 0.006849f
C1118 B.n444 VSUBS 0.006849f
C1119 B.n445 VSUBS 0.006849f
C1120 B.n446 VSUBS 0.006849f
C1121 B.n447 VSUBS 0.006849f
C1122 B.n448 VSUBS 0.006849f
C1123 B.n449 VSUBS 0.006849f
C1124 B.n450 VSUBS 0.006849f
C1125 B.n451 VSUBS 0.006849f
C1126 B.n452 VSUBS 0.006849f
C1127 B.n453 VSUBS 0.006849f
C1128 B.n454 VSUBS 0.006849f
C1129 B.n455 VSUBS 0.006849f
C1130 B.n456 VSUBS 0.006849f
C1131 B.n457 VSUBS 0.006849f
C1132 B.n458 VSUBS 0.006849f
C1133 B.n459 VSUBS 0.006849f
C1134 B.n460 VSUBS 0.006849f
C1135 B.n461 VSUBS 0.006849f
C1136 B.n462 VSUBS 0.006849f
C1137 B.n463 VSUBS 0.006849f
C1138 B.n464 VSUBS 0.006849f
C1139 B.n465 VSUBS 0.006849f
C1140 B.n466 VSUBS 0.006849f
C1141 B.n467 VSUBS 0.006849f
C1142 B.n468 VSUBS 0.006849f
C1143 B.n469 VSUBS 0.006849f
C1144 B.n470 VSUBS 0.006849f
C1145 B.n471 VSUBS 0.006849f
C1146 B.n472 VSUBS 0.006849f
C1147 B.n473 VSUBS 0.015521f
C1148 B.n474 VSUBS 0.015521f
C1149 B.n475 VSUBS 0.016105f
C1150 B.n476 VSUBS 0.006849f
C1151 B.n477 VSUBS 0.006849f
C1152 B.n478 VSUBS 0.006849f
C1153 B.n479 VSUBS 0.006849f
C1154 B.n480 VSUBS 0.006849f
C1155 B.n481 VSUBS 0.006849f
C1156 B.n482 VSUBS 0.006849f
C1157 B.n483 VSUBS 0.006849f
C1158 B.n484 VSUBS 0.006849f
C1159 B.n485 VSUBS 0.006849f
C1160 B.n486 VSUBS 0.006849f
C1161 B.n487 VSUBS 0.006849f
C1162 B.n488 VSUBS 0.006849f
C1163 B.n489 VSUBS 0.006849f
C1164 B.n490 VSUBS 0.006849f
C1165 B.n491 VSUBS 0.006849f
C1166 B.n492 VSUBS 0.006849f
C1167 B.n493 VSUBS 0.006849f
C1168 B.n494 VSUBS 0.006849f
C1169 B.n495 VSUBS 0.006849f
C1170 B.n496 VSUBS 0.006849f
C1171 B.n497 VSUBS 0.006849f
C1172 B.n498 VSUBS 0.006849f
C1173 B.n499 VSUBS 0.006849f
C1174 B.n500 VSUBS 0.006849f
C1175 B.n501 VSUBS 0.006849f
C1176 B.n502 VSUBS 0.006849f
C1177 B.n503 VSUBS 0.006849f
C1178 B.n504 VSUBS 0.006849f
C1179 B.n505 VSUBS 0.006849f
C1180 B.n506 VSUBS 0.006849f
C1181 B.n507 VSUBS 0.006849f
C1182 B.n508 VSUBS 0.006849f
C1183 B.n509 VSUBS 0.006849f
C1184 B.n510 VSUBS 0.006849f
C1185 B.n511 VSUBS 0.006849f
C1186 B.n512 VSUBS 0.006849f
C1187 B.n513 VSUBS 0.006849f
C1188 B.n514 VSUBS 0.006849f
C1189 B.n515 VSUBS 0.006849f
C1190 B.n516 VSUBS 0.006849f
C1191 B.n517 VSUBS 0.006849f
C1192 B.n518 VSUBS 0.006849f
C1193 B.n519 VSUBS 0.006849f
C1194 B.n520 VSUBS 0.006849f
C1195 B.n521 VSUBS 0.006849f
C1196 B.n522 VSUBS 0.006849f
C1197 B.n523 VSUBS 0.006849f
C1198 B.n524 VSUBS 0.006849f
C1199 B.n525 VSUBS 0.006849f
C1200 B.n526 VSUBS 0.006849f
C1201 B.n527 VSUBS 0.006849f
C1202 B.n528 VSUBS 0.006849f
C1203 B.n529 VSUBS 0.006849f
C1204 B.n530 VSUBS 0.006849f
C1205 B.n531 VSUBS 0.006849f
C1206 B.n532 VSUBS 0.006849f
C1207 B.n533 VSUBS 0.006849f
C1208 B.n534 VSUBS 0.006849f
C1209 B.n535 VSUBS 0.006849f
C1210 B.n536 VSUBS 0.006849f
C1211 B.n537 VSUBS 0.006849f
C1212 B.n538 VSUBS 0.006849f
C1213 B.n539 VSUBS 0.006849f
C1214 B.n540 VSUBS 0.006849f
C1215 B.n541 VSUBS 0.006849f
C1216 B.n542 VSUBS 0.006849f
C1217 B.n543 VSUBS 0.006849f
C1218 B.n544 VSUBS 0.006849f
C1219 B.n545 VSUBS 0.006446f
C1220 B.n546 VSUBS 0.006849f
C1221 B.n547 VSUBS 0.006849f
C1222 B.n548 VSUBS 0.003827f
C1223 B.n549 VSUBS 0.006849f
C1224 B.n550 VSUBS 0.006849f
C1225 B.n551 VSUBS 0.006849f
C1226 B.n552 VSUBS 0.006849f
C1227 B.n553 VSUBS 0.006849f
C1228 B.n554 VSUBS 0.006849f
C1229 B.n555 VSUBS 0.006849f
C1230 B.n556 VSUBS 0.006849f
C1231 B.n557 VSUBS 0.006849f
C1232 B.n558 VSUBS 0.006849f
C1233 B.n559 VSUBS 0.006849f
C1234 B.n560 VSUBS 0.006849f
C1235 B.n561 VSUBS 0.003827f
C1236 B.n562 VSUBS 0.015868f
C1237 B.n563 VSUBS 0.006446f
C1238 B.n564 VSUBS 0.006849f
C1239 B.n565 VSUBS 0.006849f
C1240 B.n566 VSUBS 0.006849f
C1241 B.n567 VSUBS 0.006849f
C1242 B.n568 VSUBS 0.006849f
C1243 B.n569 VSUBS 0.006849f
C1244 B.n570 VSUBS 0.006849f
C1245 B.n571 VSUBS 0.006849f
C1246 B.n572 VSUBS 0.006849f
C1247 B.n573 VSUBS 0.006849f
C1248 B.n574 VSUBS 0.006849f
C1249 B.n575 VSUBS 0.006849f
C1250 B.n576 VSUBS 0.006849f
C1251 B.n577 VSUBS 0.006849f
C1252 B.n578 VSUBS 0.006849f
C1253 B.n579 VSUBS 0.006849f
C1254 B.n580 VSUBS 0.006849f
C1255 B.n581 VSUBS 0.006849f
C1256 B.n582 VSUBS 0.006849f
C1257 B.n583 VSUBS 0.006849f
C1258 B.n584 VSUBS 0.006849f
C1259 B.n585 VSUBS 0.006849f
C1260 B.n586 VSUBS 0.006849f
C1261 B.n587 VSUBS 0.006849f
C1262 B.n588 VSUBS 0.006849f
C1263 B.n589 VSUBS 0.006849f
C1264 B.n590 VSUBS 0.006849f
C1265 B.n591 VSUBS 0.006849f
C1266 B.n592 VSUBS 0.006849f
C1267 B.n593 VSUBS 0.006849f
C1268 B.n594 VSUBS 0.006849f
C1269 B.n595 VSUBS 0.006849f
C1270 B.n596 VSUBS 0.006849f
C1271 B.n597 VSUBS 0.006849f
C1272 B.n598 VSUBS 0.006849f
C1273 B.n599 VSUBS 0.006849f
C1274 B.n600 VSUBS 0.006849f
C1275 B.n601 VSUBS 0.006849f
C1276 B.n602 VSUBS 0.006849f
C1277 B.n603 VSUBS 0.006849f
C1278 B.n604 VSUBS 0.006849f
C1279 B.n605 VSUBS 0.006849f
C1280 B.n606 VSUBS 0.006849f
C1281 B.n607 VSUBS 0.006849f
C1282 B.n608 VSUBS 0.006849f
C1283 B.n609 VSUBS 0.006849f
C1284 B.n610 VSUBS 0.006849f
C1285 B.n611 VSUBS 0.006849f
C1286 B.n612 VSUBS 0.006849f
C1287 B.n613 VSUBS 0.006849f
C1288 B.n614 VSUBS 0.006849f
C1289 B.n615 VSUBS 0.006849f
C1290 B.n616 VSUBS 0.006849f
C1291 B.n617 VSUBS 0.006849f
C1292 B.n618 VSUBS 0.006849f
C1293 B.n619 VSUBS 0.006849f
C1294 B.n620 VSUBS 0.006849f
C1295 B.n621 VSUBS 0.006849f
C1296 B.n622 VSUBS 0.006849f
C1297 B.n623 VSUBS 0.006849f
C1298 B.n624 VSUBS 0.006849f
C1299 B.n625 VSUBS 0.006849f
C1300 B.n626 VSUBS 0.006849f
C1301 B.n627 VSUBS 0.006849f
C1302 B.n628 VSUBS 0.006849f
C1303 B.n629 VSUBS 0.006849f
C1304 B.n630 VSUBS 0.006849f
C1305 B.n631 VSUBS 0.006849f
C1306 B.n632 VSUBS 0.006849f
C1307 B.n633 VSUBS 0.006849f
C1308 B.n634 VSUBS 0.016105f
C1309 B.n635 VSUBS 0.015521f
C1310 B.n636 VSUBS 0.015521f
C1311 B.n637 VSUBS 0.006849f
C1312 B.n638 VSUBS 0.006849f
C1313 B.n639 VSUBS 0.006849f
C1314 B.n640 VSUBS 0.006849f
C1315 B.n641 VSUBS 0.006849f
C1316 B.n642 VSUBS 0.006849f
C1317 B.n643 VSUBS 0.006849f
C1318 B.n644 VSUBS 0.006849f
C1319 B.n645 VSUBS 0.006849f
C1320 B.n646 VSUBS 0.006849f
C1321 B.n647 VSUBS 0.006849f
C1322 B.n648 VSUBS 0.006849f
C1323 B.n649 VSUBS 0.006849f
C1324 B.n650 VSUBS 0.006849f
C1325 B.n651 VSUBS 0.006849f
C1326 B.n652 VSUBS 0.006849f
C1327 B.n653 VSUBS 0.006849f
C1328 B.n654 VSUBS 0.006849f
C1329 B.n655 VSUBS 0.006849f
C1330 B.n656 VSUBS 0.006849f
C1331 B.n657 VSUBS 0.006849f
C1332 B.n658 VSUBS 0.006849f
C1333 B.n659 VSUBS 0.006849f
C1334 B.n660 VSUBS 0.006849f
C1335 B.n661 VSUBS 0.006849f
C1336 B.n662 VSUBS 0.006849f
C1337 B.n663 VSUBS 0.006849f
C1338 B.n664 VSUBS 0.006849f
C1339 B.n665 VSUBS 0.006849f
C1340 B.n666 VSUBS 0.006849f
C1341 B.n667 VSUBS 0.006849f
C1342 B.n668 VSUBS 0.006849f
C1343 B.n669 VSUBS 0.006849f
C1344 B.n670 VSUBS 0.006849f
C1345 B.n671 VSUBS 0.006849f
C1346 B.n672 VSUBS 0.006849f
C1347 B.n673 VSUBS 0.006849f
C1348 B.n674 VSUBS 0.006849f
C1349 B.n675 VSUBS 0.006849f
C1350 B.n676 VSUBS 0.006849f
C1351 B.n677 VSUBS 0.006849f
C1352 B.n678 VSUBS 0.006849f
C1353 B.n679 VSUBS 0.008937f
C1354 B.n680 VSUBS 0.009521f
C1355 B.n681 VSUBS 0.018933f
.ends

