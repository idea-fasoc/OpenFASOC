* NGSPICE file created from diff_pair_sample_1290.ext - technology: sky130A

.subckt diff_pair_sample_1290 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t15 VN.t0 VDD2.t7 B.t7 sky130_fd_pr__nfet_01v8 ad=7.2969 pd=38.2 as=3.08715 ps=19.04 w=18.71 l=3.13
X1 B.t21 B.t19 B.t20 B.t16 sky130_fd_pr__nfet_01v8 ad=7.2969 pd=38.2 as=0 ps=0 w=18.71 l=3.13
X2 VTAIL.t14 VN.t1 VDD2.t6 B.t0 sky130_fd_pr__nfet_01v8 ad=3.08715 pd=19.04 as=3.08715 ps=19.04 w=18.71 l=3.13
X3 VDD1.t7 VP.t0 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=3.08715 pd=19.04 as=7.2969 ps=38.2 w=18.71 l=3.13
X4 VTAIL.t0 VP.t1 VDD1.t6 B.t0 sky130_fd_pr__nfet_01v8 ad=3.08715 pd=19.04 as=3.08715 ps=19.04 w=18.71 l=3.13
X5 B.t18 B.t15 B.t17 B.t16 sky130_fd_pr__nfet_01v8 ad=7.2969 pd=38.2 as=0 ps=0 w=18.71 l=3.13
X6 VTAIL.t1 VP.t2 VDD1.t5 B.t1 sky130_fd_pr__nfet_01v8 ad=7.2969 pd=38.2 as=3.08715 ps=19.04 w=18.71 l=3.13
X7 VDD2.t5 VN.t2 VTAIL.t13 B.t6 sky130_fd_pr__nfet_01v8 ad=3.08715 pd=19.04 as=7.2969 ps=38.2 w=18.71 l=3.13
X8 VTAIL.t12 VN.t3 VDD2.t4 B.t3 sky130_fd_pr__nfet_01v8 ad=3.08715 pd=19.04 as=3.08715 ps=19.04 w=18.71 l=3.13
X9 VDD1.t4 VP.t3 VTAIL.t6 B.t6 sky130_fd_pr__nfet_01v8 ad=3.08715 pd=19.04 as=7.2969 ps=38.2 w=18.71 l=3.13
X10 VDD2.t1 VN.t4 VTAIL.t11 B.t4 sky130_fd_pr__nfet_01v8 ad=3.08715 pd=19.04 as=3.08715 ps=19.04 w=18.71 l=3.13
X11 VDD2.t0 VN.t5 VTAIL.t10 B.t2 sky130_fd_pr__nfet_01v8 ad=3.08715 pd=19.04 as=7.2969 ps=38.2 w=18.71 l=3.13
X12 VTAIL.t9 VN.t6 VDD2.t3 B.t1 sky130_fd_pr__nfet_01v8 ad=7.2969 pd=38.2 as=3.08715 ps=19.04 w=18.71 l=3.13
X13 B.t14 B.t12 B.t13 B.t9 sky130_fd_pr__nfet_01v8 ad=7.2969 pd=38.2 as=0 ps=0 w=18.71 l=3.13
X14 VDD1.t3 VP.t4 VTAIL.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=3.08715 pd=19.04 as=3.08715 ps=19.04 w=18.71 l=3.13
X15 VDD2.t2 VN.t7 VTAIL.t8 B.t5 sky130_fd_pr__nfet_01v8 ad=3.08715 pd=19.04 as=3.08715 ps=19.04 w=18.71 l=3.13
X16 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=7.2969 pd=38.2 as=0 ps=0 w=18.71 l=3.13
X17 VTAIL.t7 VP.t5 VDD1.t2 B.t7 sky130_fd_pr__nfet_01v8 ad=7.2969 pd=38.2 as=3.08715 ps=19.04 w=18.71 l=3.13
X18 VTAIL.t3 VP.t6 VDD1.t1 B.t3 sky130_fd_pr__nfet_01v8 ad=3.08715 pd=19.04 as=3.08715 ps=19.04 w=18.71 l=3.13
X19 VDD1.t0 VP.t7 VTAIL.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=3.08715 pd=19.04 as=3.08715 ps=19.04 w=18.71 l=3.13
R0 VN.n39 VN.t5 177.48
R1 VN.n8 VN.t6 177.48
R2 VN.n60 VN.n59 161.3
R3 VN.n58 VN.n32 161.3
R4 VN.n57 VN.n56 161.3
R5 VN.n55 VN.n33 161.3
R6 VN.n54 VN.n53 161.3
R7 VN.n52 VN.n34 161.3
R8 VN.n51 VN.n50 161.3
R9 VN.n49 VN.n48 161.3
R10 VN.n47 VN.n36 161.3
R11 VN.n46 VN.n45 161.3
R12 VN.n44 VN.n37 161.3
R13 VN.n43 VN.n42 161.3
R14 VN.n41 VN.n38 161.3
R15 VN.n29 VN.n28 161.3
R16 VN.n27 VN.n1 161.3
R17 VN.n26 VN.n25 161.3
R18 VN.n24 VN.n2 161.3
R19 VN.n23 VN.n22 161.3
R20 VN.n21 VN.n3 161.3
R21 VN.n20 VN.n19 161.3
R22 VN.n18 VN.n17 161.3
R23 VN.n16 VN.n5 161.3
R24 VN.n15 VN.n14 161.3
R25 VN.n13 VN.n6 161.3
R26 VN.n12 VN.n11 161.3
R27 VN.n10 VN.n7 161.3
R28 VN.n9 VN.t4 144.061
R29 VN.n4 VN.t3 144.061
R30 VN.n0 VN.t2 144.061
R31 VN.n40 VN.t1 144.061
R32 VN.n35 VN.t7 144.061
R33 VN.n31 VN.t0 144.061
R34 VN.n30 VN.n0 68.5364
R35 VN.n61 VN.n31 68.5364
R36 VN VN.n61 58.8011
R37 VN.n15 VN.n6 56.5193
R38 VN.n26 VN.n2 56.5193
R39 VN.n46 VN.n37 56.5193
R40 VN.n57 VN.n33 56.5193
R41 VN.n9 VN.n8 50.4514
R42 VN.n40 VN.n39 50.4514
R43 VN.n11 VN.n10 24.4675
R44 VN.n11 VN.n6 24.4675
R45 VN.n16 VN.n15 24.4675
R46 VN.n17 VN.n16 24.4675
R47 VN.n21 VN.n20 24.4675
R48 VN.n22 VN.n21 24.4675
R49 VN.n22 VN.n2 24.4675
R50 VN.n27 VN.n26 24.4675
R51 VN.n28 VN.n27 24.4675
R52 VN.n42 VN.n37 24.4675
R53 VN.n42 VN.n41 24.4675
R54 VN.n53 VN.n33 24.4675
R55 VN.n53 VN.n52 24.4675
R56 VN.n52 VN.n51 24.4675
R57 VN.n48 VN.n47 24.4675
R58 VN.n47 VN.n46 24.4675
R59 VN.n59 VN.n58 24.4675
R60 VN.n58 VN.n57 24.4675
R61 VN.n10 VN.n9 23.4888
R62 VN.n17 VN.n4 23.4888
R63 VN.n41 VN.n40 23.4888
R64 VN.n48 VN.n35 23.4888
R65 VN.n28 VN.n0 21.5315
R66 VN.n59 VN.n31 21.5315
R67 VN.n39 VN.n38 3.84099
R68 VN.n8 VN.n7 3.84099
R69 VN.n20 VN.n4 0.97918
R70 VN.n51 VN.n35 0.97918
R71 VN.n61 VN.n60 0.354971
R72 VN.n30 VN.n29 0.354971
R73 VN VN.n30 0.26696
R74 VN.n60 VN.n32 0.189894
R75 VN.n56 VN.n32 0.189894
R76 VN.n56 VN.n55 0.189894
R77 VN.n55 VN.n54 0.189894
R78 VN.n54 VN.n34 0.189894
R79 VN.n50 VN.n34 0.189894
R80 VN.n50 VN.n49 0.189894
R81 VN.n49 VN.n36 0.189894
R82 VN.n45 VN.n36 0.189894
R83 VN.n45 VN.n44 0.189894
R84 VN.n44 VN.n43 0.189894
R85 VN.n43 VN.n38 0.189894
R86 VN.n12 VN.n7 0.189894
R87 VN.n13 VN.n12 0.189894
R88 VN.n14 VN.n13 0.189894
R89 VN.n14 VN.n5 0.189894
R90 VN.n18 VN.n5 0.189894
R91 VN.n19 VN.n18 0.189894
R92 VN.n19 VN.n3 0.189894
R93 VN.n23 VN.n3 0.189894
R94 VN.n24 VN.n23 0.189894
R95 VN.n25 VN.n24 0.189894
R96 VN.n25 VN.n1 0.189894
R97 VN.n29 VN.n1 0.189894
R98 VDD2.n2 VDD2.n1 63.7374
R99 VDD2.n2 VDD2.n0 63.7374
R100 VDD2 VDD2.n5 63.7344
R101 VDD2.n4 VDD2.n3 62.3024
R102 VDD2.n4 VDD2.n2 53.267
R103 VDD2 VDD2.n4 1.55007
R104 VDD2.n5 VDD2.t6 1.05876
R105 VDD2.n5 VDD2.t0 1.05876
R106 VDD2.n3 VDD2.t7 1.05876
R107 VDD2.n3 VDD2.t2 1.05876
R108 VDD2.n1 VDD2.t4 1.05876
R109 VDD2.n1 VDD2.t5 1.05876
R110 VDD2.n0 VDD2.t3 1.05876
R111 VDD2.n0 VDD2.t1 1.05876
R112 VTAIL.n838 VTAIL.n837 289.615
R113 VTAIL.n104 VTAIL.n103 289.615
R114 VTAIL.n208 VTAIL.n207 289.615
R115 VTAIL.n314 VTAIL.n313 289.615
R116 VTAIL.n734 VTAIL.n733 289.615
R117 VTAIL.n628 VTAIL.n627 289.615
R118 VTAIL.n524 VTAIL.n523 289.615
R119 VTAIL.n418 VTAIL.n417 289.615
R120 VTAIL.n771 VTAIL.n770 185
R121 VTAIL.n773 VTAIL.n772 185
R122 VTAIL.n766 VTAIL.n765 185
R123 VTAIL.n779 VTAIL.n778 185
R124 VTAIL.n781 VTAIL.n780 185
R125 VTAIL.n762 VTAIL.n761 185
R126 VTAIL.n788 VTAIL.n787 185
R127 VTAIL.n789 VTAIL.n760 185
R128 VTAIL.n791 VTAIL.n790 185
R129 VTAIL.n758 VTAIL.n757 185
R130 VTAIL.n797 VTAIL.n796 185
R131 VTAIL.n799 VTAIL.n798 185
R132 VTAIL.n754 VTAIL.n753 185
R133 VTAIL.n805 VTAIL.n804 185
R134 VTAIL.n807 VTAIL.n806 185
R135 VTAIL.n750 VTAIL.n749 185
R136 VTAIL.n813 VTAIL.n812 185
R137 VTAIL.n815 VTAIL.n814 185
R138 VTAIL.n746 VTAIL.n745 185
R139 VTAIL.n821 VTAIL.n820 185
R140 VTAIL.n823 VTAIL.n822 185
R141 VTAIL.n742 VTAIL.n741 185
R142 VTAIL.n829 VTAIL.n828 185
R143 VTAIL.n831 VTAIL.n830 185
R144 VTAIL.n738 VTAIL.n737 185
R145 VTAIL.n837 VTAIL.n836 185
R146 VTAIL.n37 VTAIL.n36 185
R147 VTAIL.n39 VTAIL.n38 185
R148 VTAIL.n32 VTAIL.n31 185
R149 VTAIL.n45 VTAIL.n44 185
R150 VTAIL.n47 VTAIL.n46 185
R151 VTAIL.n28 VTAIL.n27 185
R152 VTAIL.n54 VTAIL.n53 185
R153 VTAIL.n55 VTAIL.n26 185
R154 VTAIL.n57 VTAIL.n56 185
R155 VTAIL.n24 VTAIL.n23 185
R156 VTAIL.n63 VTAIL.n62 185
R157 VTAIL.n65 VTAIL.n64 185
R158 VTAIL.n20 VTAIL.n19 185
R159 VTAIL.n71 VTAIL.n70 185
R160 VTAIL.n73 VTAIL.n72 185
R161 VTAIL.n16 VTAIL.n15 185
R162 VTAIL.n79 VTAIL.n78 185
R163 VTAIL.n81 VTAIL.n80 185
R164 VTAIL.n12 VTAIL.n11 185
R165 VTAIL.n87 VTAIL.n86 185
R166 VTAIL.n89 VTAIL.n88 185
R167 VTAIL.n8 VTAIL.n7 185
R168 VTAIL.n95 VTAIL.n94 185
R169 VTAIL.n97 VTAIL.n96 185
R170 VTAIL.n4 VTAIL.n3 185
R171 VTAIL.n103 VTAIL.n102 185
R172 VTAIL.n141 VTAIL.n140 185
R173 VTAIL.n143 VTAIL.n142 185
R174 VTAIL.n136 VTAIL.n135 185
R175 VTAIL.n149 VTAIL.n148 185
R176 VTAIL.n151 VTAIL.n150 185
R177 VTAIL.n132 VTAIL.n131 185
R178 VTAIL.n158 VTAIL.n157 185
R179 VTAIL.n159 VTAIL.n130 185
R180 VTAIL.n161 VTAIL.n160 185
R181 VTAIL.n128 VTAIL.n127 185
R182 VTAIL.n167 VTAIL.n166 185
R183 VTAIL.n169 VTAIL.n168 185
R184 VTAIL.n124 VTAIL.n123 185
R185 VTAIL.n175 VTAIL.n174 185
R186 VTAIL.n177 VTAIL.n176 185
R187 VTAIL.n120 VTAIL.n119 185
R188 VTAIL.n183 VTAIL.n182 185
R189 VTAIL.n185 VTAIL.n184 185
R190 VTAIL.n116 VTAIL.n115 185
R191 VTAIL.n191 VTAIL.n190 185
R192 VTAIL.n193 VTAIL.n192 185
R193 VTAIL.n112 VTAIL.n111 185
R194 VTAIL.n199 VTAIL.n198 185
R195 VTAIL.n201 VTAIL.n200 185
R196 VTAIL.n108 VTAIL.n107 185
R197 VTAIL.n207 VTAIL.n206 185
R198 VTAIL.n247 VTAIL.n246 185
R199 VTAIL.n249 VTAIL.n248 185
R200 VTAIL.n242 VTAIL.n241 185
R201 VTAIL.n255 VTAIL.n254 185
R202 VTAIL.n257 VTAIL.n256 185
R203 VTAIL.n238 VTAIL.n237 185
R204 VTAIL.n264 VTAIL.n263 185
R205 VTAIL.n265 VTAIL.n236 185
R206 VTAIL.n267 VTAIL.n266 185
R207 VTAIL.n234 VTAIL.n233 185
R208 VTAIL.n273 VTAIL.n272 185
R209 VTAIL.n275 VTAIL.n274 185
R210 VTAIL.n230 VTAIL.n229 185
R211 VTAIL.n281 VTAIL.n280 185
R212 VTAIL.n283 VTAIL.n282 185
R213 VTAIL.n226 VTAIL.n225 185
R214 VTAIL.n289 VTAIL.n288 185
R215 VTAIL.n291 VTAIL.n290 185
R216 VTAIL.n222 VTAIL.n221 185
R217 VTAIL.n297 VTAIL.n296 185
R218 VTAIL.n299 VTAIL.n298 185
R219 VTAIL.n218 VTAIL.n217 185
R220 VTAIL.n305 VTAIL.n304 185
R221 VTAIL.n307 VTAIL.n306 185
R222 VTAIL.n214 VTAIL.n213 185
R223 VTAIL.n313 VTAIL.n312 185
R224 VTAIL.n733 VTAIL.n732 185
R225 VTAIL.n634 VTAIL.n633 185
R226 VTAIL.n727 VTAIL.n726 185
R227 VTAIL.n725 VTAIL.n724 185
R228 VTAIL.n638 VTAIL.n637 185
R229 VTAIL.n719 VTAIL.n718 185
R230 VTAIL.n717 VTAIL.n716 185
R231 VTAIL.n642 VTAIL.n641 185
R232 VTAIL.n711 VTAIL.n710 185
R233 VTAIL.n709 VTAIL.n708 185
R234 VTAIL.n646 VTAIL.n645 185
R235 VTAIL.n703 VTAIL.n702 185
R236 VTAIL.n701 VTAIL.n700 185
R237 VTAIL.n650 VTAIL.n649 185
R238 VTAIL.n695 VTAIL.n694 185
R239 VTAIL.n693 VTAIL.n692 185
R240 VTAIL.n654 VTAIL.n653 185
R241 VTAIL.n658 VTAIL.n656 185
R242 VTAIL.n687 VTAIL.n686 185
R243 VTAIL.n685 VTAIL.n684 185
R244 VTAIL.n660 VTAIL.n659 185
R245 VTAIL.n679 VTAIL.n678 185
R246 VTAIL.n677 VTAIL.n676 185
R247 VTAIL.n664 VTAIL.n663 185
R248 VTAIL.n671 VTAIL.n670 185
R249 VTAIL.n669 VTAIL.n668 185
R250 VTAIL.n627 VTAIL.n626 185
R251 VTAIL.n528 VTAIL.n527 185
R252 VTAIL.n621 VTAIL.n620 185
R253 VTAIL.n619 VTAIL.n618 185
R254 VTAIL.n532 VTAIL.n531 185
R255 VTAIL.n613 VTAIL.n612 185
R256 VTAIL.n611 VTAIL.n610 185
R257 VTAIL.n536 VTAIL.n535 185
R258 VTAIL.n605 VTAIL.n604 185
R259 VTAIL.n603 VTAIL.n602 185
R260 VTAIL.n540 VTAIL.n539 185
R261 VTAIL.n597 VTAIL.n596 185
R262 VTAIL.n595 VTAIL.n594 185
R263 VTAIL.n544 VTAIL.n543 185
R264 VTAIL.n589 VTAIL.n588 185
R265 VTAIL.n587 VTAIL.n586 185
R266 VTAIL.n548 VTAIL.n547 185
R267 VTAIL.n552 VTAIL.n550 185
R268 VTAIL.n581 VTAIL.n580 185
R269 VTAIL.n579 VTAIL.n578 185
R270 VTAIL.n554 VTAIL.n553 185
R271 VTAIL.n573 VTAIL.n572 185
R272 VTAIL.n571 VTAIL.n570 185
R273 VTAIL.n558 VTAIL.n557 185
R274 VTAIL.n565 VTAIL.n564 185
R275 VTAIL.n563 VTAIL.n562 185
R276 VTAIL.n523 VTAIL.n522 185
R277 VTAIL.n424 VTAIL.n423 185
R278 VTAIL.n517 VTAIL.n516 185
R279 VTAIL.n515 VTAIL.n514 185
R280 VTAIL.n428 VTAIL.n427 185
R281 VTAIL.n509 VTAIL.n508 185
R282 VTAIL.n507 VTAIL.n506 185
R283 VTAIL.n432 VTAIL.n431 185
R284 VTAIL.n501 VTAIL.n500 185
R285 VTAIL.n499 VTAIL.n498 185
R286 VTAIL.n436 VTAIL.n435 185
R287 VTAIL.n493 VTAIL.n492 185
R288 VTAIL.n491 VTAIL.n490 185
R289 VTAIL.n440 VTAIL.n439 185
R290 VTAIL.n485 VTAIL.n484 185
R291 VTAIL.n483 VTAIL.n482 185
R292 VTAIL.n444 VTAIL.n443 185
R293 VTAIL.n448 VTAIL.n446 185
R294 VTAIL.n477 VTAIL.n476 185
R295 VTAIL.n475 VTAIL.n474 185
R296 VTAIL.n450 VTAIL.n449 185
R297 VTAIL.n469 VTAIL.n468 185
R298 VTAIL.n467 VTAIL.n466 185
R299 VTAIL.n454 VTAIL.n453 185
R300 VTAIL.n461 VTAIL.n460 185
R301 VTAIL.n459 VTAIL.n458 185
R302 VTAIL.n417 VTAIL.n416 185
R303 VTAIL.n318 VTAIL.n317 185
R304 VTAIL.n411 VTAIL.n410 185
R305 VTAIL.n409 VTAIL.n408 185
R306 VTAIL.n322 VTAIL.n321 185
R307 VTAIL.n403 VTAIL.n402 185
R308 VTAIL.n401 VTAIL.n400 185
R309 VTAIL.n326 VTAIL.n325 185
R310 VTAIL.n395 VTAIL.n394 185
R311 VTAIL.n393 VTAIL.n392 185
R312 VTAIL.n330 VTAIL.n329 185
R313 VTAIL.n387 VTAIL.n386 185
R314 VTAIL.n385 VTAIL.n384 185
R315 VTAIL.n334 VTAIL.n333 185
R316 VTAIL.n379 VTAIL.n378 185
R317 VTAIL.n377 VTAIL.n376 185
R318 VTAIL.n338 VTAIL.n337 185
R319 VTAIL.n342 VTAIL.n340 185
R320 VTAIL.n371 VTAIL.n370 185
R321 VTAIL.n369 VTAIL.n368 185
R322 VTAIL.n344 VTAIL.n343 185
R323 VTAIL.n363 VTAIL.n362 185
R324 VTAIL.n361 VTAIL.n360 185
R325 VTAIL.n348 VTAIL.n347 185
R326 VTAIL.n355 VTAIL.n354 185
R327 VTAIL.n353 VTAIL.n352 185
R328 VTAIL.n769 VTAIL.t13 149.524
R329 VTAIL.n35 VTAIL.t9 149.524
R330 VTAIL.n139 VTAIL.t2 149.524
R331 VTAIL.n245 VTAIL.t7 149.524
R332 VTAIL.n667 VTAIL.t6 149.524
R333 VTAIL.n561 VTAIL.t1 149.524
R334 VTAIL.n457 VTAIL.t10 149.524
R335 VTAIL.n351 VTAIL.t15 149.524
R336 VTAIL.n772 VTAIL.n771 104.615
R337 VTAIL.n772 VTAIL.n765 104.615
R338 VTAIL.n779 VTAIL.n765 104.615
R339 VTAIL.n780 VTAIL.n779 104.615
R340 VTAIL.n780 VTAIL.n761 104.615
R341 VTAIL.n788 VTAIL.n761 104.615
R342 VTAIL.n789 VTAIL.n788 104.615
R343 VTAIL.n790 VTAIL.n789 104.615
R344 VTAIL.n790 VTAIL.n757 104.615
R345 VTAIL.n797 VTAIL.n757 104.615
R346 VTAIL.n798 VTAIL.n797 104.615
R347 VTAIL.n798 VTAIL.n753 104.615
R348 VTAIL.n805 VTAIL.n753 104.615
R349 VTAIL.n806 VTAIL.n805 104.615
R350 VTAIL.n806 VTAIL.n749 104.615
R351 VTAIL.n813 VTAIL.n749 104.615
R352 VTAIL.n814 VTAIL.n813 104.615
R353 VTAIL.n814 VTAIL.n745 104.615
R354 VTAIL.n821 VTAIL.n745 104.615
R355 VTAIL.n822 VTAIL.n821 104.615
R356 VTAIL.n822 VTAIL.n741 104.615
R357 VTAIL.n829 VTAIL.n741 104.615
R358 VTAIL.n830 VTAIL.n829 104.615
R359 VTAIL.n830 VTAIL.n737 104.615
R360 VTAIL.n837 VTAIL.n737 104.615
R361 VTAIL.n38 VTAIL.n37 104.615
R362 VTAIL.n38 VTAIL.n31 104.615
R363 VTAIL.n45 VTAIL.n31 104.615
R364 VTAIL.n46 VTAIL.n45 104.615
R365 VTAIL.n46 VTAIL.n27 104.615
R366 VTAIL.n54 VTAIL.n27 104.615
R367 VTAIL.n55 VTAIL.n54 104.615
R368 VTAIL.n56 VTAIL.n55 104.615
R369 VTAIL.n56 VTAIL.n23 104.615
R370 VTAIL.n63 VTAIL.n23 104.615
R371 VTAIL.n64 VTAIL.n63 104.615
R372 VTAIL.n64 VTAIL.n19 104.615
R373 VTAIL.n71 VTAIL.n19 104.615
R374 VTAIL.n72 VTAIL.n71 104.615
R375 VTAIL.n72 VTAIL.n15 104.615
R376 VTAIL.n79 VTAIL.n15 104.615
R377 VTAIL.n80 VTAIL.n79 104.615
R378 VTAIL.n80 VTAIL.n11 104.615
R379 VTAIL.n87 VTAIL.n11 104.615
R380 VTAIL.n88 VTAIL.n87 104.615
R381 VTAIL.n88 VTAIL.n7 104.615
R382 VTAIL.n95 VTAIL.n7 104.615
R383 VTAIL.n96 VTAIL.n95 104.615
R384 VTAIL.n96 VTAIL.n3 104.615
R385 VTAIL.n103 VTAIL.n3 104.615
R386 VTAIL.n142 VTAIL.n141 104.615
R387 VTAIL.n142 VTAIL.n135 104.615
R388 VTAIL.n149 VTAIL.n135 104.615
R389 VTAIL.n150 VTAIL.n149 104.615
R390 VTAIL.n150 VTAIL.n131 104.615
R391 VTAIL.n158 VTAIL.n131 104.615
R392 VTAIL.n159 VTAIL.n158 104.615
R393 VTAIL.n160 VTAIL.n159 104.615
R394 VTAIL.n160 VTAIL.n127 104.615
R395 VTAIL.n167 VTAIL.n127 104.615
R396 VTAIL.n168 VTAIL.n167 104.615
R397 VTAIL.n168 VTAIL.n123 104.615
R398 VTAIL.n175 VTAIL.n123 104.615
R399 VTAIL.n176 VTAIL.n175 104.615
R400 VTAIL.n176 VTAIL.n119 104.615
R401 VTAIL.n183 VTAIL.n119 104.615
R402 VTAIL.n184 VTAIL.n183 104.615
R403 VTAIL.n184 VTAIL.n115 104.615
R404 VTAIL.n191 VTAIL.n115 104.615
R405 VTAIL.n192 VTAIL.n191 104.615
R406 VTAIL.n192 VTAIL.n111 104.615
R407 VTAIL.n199 VTAIL.n111 104.615
R408 VTAIL.n200 VTAIL.n199 104.615
R409 VTAIL.n200 VTAIL.n107 104.615
R410 VTAIL.n207 VTAIL.n107 104.615
R411 VTAIL.n248 VTAIL.n247 104.615
R412 VTAIL.n248 VTAIL.n241 104.615
R413 VTAIL.n255 VTAIL.n241 104.615
R414 VTAIL.n256 VTAIL.n255 104.615
R415 VTAIL.n256 VTAIL.n237 104.615
R416 VTAIL.n264 VTAIL.n237 104.615
R417 VTAIL.n265 VTAIL.n264 104.615
R418 VTAIL.n266 VTAIL.n265 104.615
R419 VTAIL.n266 VTAIL.n233 104.615
R420 VTAIL.n273 VTAIL.n233 104.615
R421 VTAIL.n274 VTAIL.n273 104.615
R422 VTAIL.n274 VTAIL.n229 104.615
R423 VTAIL.n281 VTAIL.n229 104.615
R424 VTAIL.n282 VTAIL.n281 104.615
R425 VTAIL.n282 VTAIL.n225 104.615
R426 VTAIL.n289 VTAIL.n225 104.615
R427 VTAIL.n290 VTAIL.n289 104.615
R428 VTAIL.n290 VTAIL.n221 104.615
R429 VTAIL.n297 VTAIL.n221 104.615
R430 VTAIL.n298 VTAIL.n297 104.615
R431 VTAIL.n298 VTAIL.n217 104.615
R432 VTAIL.n305 VTAIL.n217 104.615
R433 VTAIL.n306 VTAIL.n305 104.615
R434 VTAIL.n306 VTAIL.n213 104.615
R435 VTAIL.n313 VTAIL.n213 104.615
R436 VTAIL.n733 VTAIL.n633 104.615
R437 VTAIL.n726 VTAIL.n633 104.615
R438 VTAIL.n726 VTAIL.n725 104.615
R439 VTAIL.n725 VTAIL.n637 104.615
R440 VTAIL.n718 VTAIL.n637 104.615
R441 VTAIL.n718 VTAIL.n717 104.615
R442 VTAIL.n717 VTAIL.n641 104.615
R443 VTAIL.n710 VTAIL.n641 104.615
R444 VTAIL.n710 VTAIL.n709 104.615
R445 VTAIL.n709 VTAIL.n645 104.615
R446 VTAIL.n702 VTAIL.n645 104.615
R447 VTAIL.n702 VTAIL.n701 104.615
R448 VTAIL.n701 VTAIL.n649 104.615
R449 VTAIL.n694 VTAIL.n649 104.615
R450 VTAIL.n694 VTAIL.n693 104.615
R451 VTAIL.n693 VTAIL.n653 104.615
R452 VTAIL.n658 VTAIL.n653 104.615
R453 VTAIL.n686 VTAIL.n658 104.615
R454 VTAIL.n686 VTAIL.n685 104.615
R455 VTAIL.n685 VTAIL.n659 104.615
R456 VTAIL.n678 VTAIL.n659 104.615
R457 VTAIL.n678 VTAIL.n677 104.615
R458 VTAIL.n677 VTAIL.n663 104.615
R459 VTAIL.n670 VTAIL.n663 104.615
R460 VTAIL.n670 VTAIL.n669 104.615
R461 VTAIL.n627 VTAIL.n527 104.615
R462 VTAIL.n620 VTAIL.n527 104.615
R463 VTAIL.n620 VTAIL.n619 104.615
R464 VTAIL.n619 VTAIL.n531 104.615
R465 VTAIL.n612 VTAIL.n531 104.615
R466 VTAIL.n612 VTAIL.n611 104.615
R467 VTAIL.n611 VTAIL.n535 104.615
R468 VTAIL.n604 VTAIL.n535 104.615
R469 VTAIL.n604 VTAIL.n603 104.615
R470 VTAIL.n603 VTAIL.n539 104.615
R471 VTAIL.n596 VTAIL.n539 104.615
R472 VTAIL.n596 VTAIL.n595 104.615
R473 VTAIL.n595 VTAIL.n543 104.615
R474 VTAIL.n588 VTAIL.n543 104.615
R475 VTAIL.n588 VTAIL.n587 104.615
R476 VTAIL.n587 VTAIL.n547 104.615
R477 VTAIL.n552 VTAIL.n547 104.615
R478 VTAIL.n580 VTAIL.n552 104.615
R479 VTAIL.n580 VTAIL.n579 104.615
R480 VTAIL.n579 VTAIL.n553 104.615
R481 VTAIL.n572 VTAIL.n553 104.615
R482 VTAIL.n572 VTAIL.n571 104.615
R483 VTAIL.n571 VTAIL.n557 104.615
R484 VTAIL.n564 VTAIL.n557 104.615
R485 VTAIL.n564 VTAIL.n563 104.615
R486 VTAIL.n523 VTAIL.n423 104.615
R487 VTAIL.n516 VTAIL.n423 104.615
R488 VTAIL.n516 VTAIL.n515 104.615
R489 VTAIL.n515 VTAIL.n427 104.615
R490 VTAIL.n508 VTAIL.n427 104.615
R491 VTAIL.n508 VTAIL.n507 104.615
R492 VTAIL.n507 VTAIL.n431 104.615
R493 VTAIL.n500 VTAIL.n431 104.615
R494 VTAIL.n500 VTAIL.n499 104.615
R495 VTAIL.n499 VTAIL.n435 104.615
R496 VTAIL.n492 VTAIL.n435 104.615
R497 VTAIL.n492 VTAIL.n491 104.615
R498 VTAIL.n491 VTAIL.n439 104.615
R499 VTAIL.n484 VTAIL.n439 104.615
R500 VTAIL.n484 VTAIL.n483 104.615
R501 VTAIL.n483 VTAIL.n443 104.615
R502 VTAIL.n448 VTAIL.n443 104.615
R503 VTAIL.n476 VTAIL.n448 104.615
R504 VTAIL.n476 VTAIL.n475 104.615
R505 VTAIL.n475 VTAIL.n449 104.615
R506 VTAIL.n468 VTAIL.n449 104.615
R507 VTAIL.n468 VTAIL.n467 104.615
R508 VTAIL.n467 VTAIL.n453 104.615
R509 VTAIL.n460 VTAIL.n453 104.615
R510 VTAIL.n460 VTAIL.n459 104.615
R511 VTAIL.n417 VTAIL.n317 104.615
R512 VTAIL.n410 VTAIL.n317 104.615
R513 VTAIL.n410 VTAIL.n409 104.615
R514 VTAIL.n409 VTAIL.n321 104.615
R515 VTAIL.n402 VTAIL.n321 104.615
R516 VTAIL.n402 VTAIL.n401 104.615
R517 VTAIL.n401 VTAIL.n325 104.615
R518 VTAIL.n394 VTAIL.n325 104.615
R519 VTAIL.n394 VTAIL.n393 104.615
R520 VTAIL.n393 VTAIL.n329 104.615
R521 VTAIL.n386 VTAIL.n329 104.615
R522 VTAIL.n386 VTAIL.n385 104.615
R523 VTAIL.n385 VTAIL.n333 104.615
R524 VTAIL.n378 VTAIL.n333 104.615
R525 VTAIL.n378 VTAIL.n377 104.615
R526 VTAIL.n377 VTAIL.n337 104.615
R527 VTAIL.n342 VTAIL.n337 104.615
R528 VTAIL.n370 VTAIL.n342 104.615
R529 VTAIL.n370 VTAIL.n369 104.615
R530 VTAIL.n369 VTAIL.n343 104.615
R531 VTAIL.n362 VTAIL.n343 104.615
R532 VTAIL.n362 VTAIL.n361 104.615
R533 VTAIL.n361 VTAIL.n347 104.615
R534 VTAIL.n354 VTAIL.n347 104.615
R535 VTAIL.n354 VTAIL.n353 104.615
R536 VTAIL.n771 VTAIL.t13 52.3082
R537 VTAIL.n37 VTAIL.t9 52.3082
R538 VTAIL.n141 VTAIL.t2 52.3082
R539 VTAIL.n247 VTAIL.t7 52.3082
R540 VTAIL.n669 VTAIL.t6 52.3082
R541 VTAIL.n563 VTAIL.t1 52.3082
R542 VTAIL.n459 VTAIL.t10 52.3082
R543 VTAIL.n353 VTAIL.t15 52.3082
R544 VTAIL.n631 VTAIL.n630 45.6236
R545 VTAIL.n421 VTAIL.n420 45.6236
R546 VTAIL.n1 VTAIL.n0 45.6226
R547 VTAIL.n211 VTAIL.n210 45.6226
R548 VTAIL.n839 VTAIL.n838 33.9308
R549 VTAIL.n105 VTAIL.n104 33.9308
R550 VTAIL.n209 VTAIL.n208 33.9308
R551 VTAIL.n315 VTAIL.n314 33.9308
R552 VTAIL.n735 VTAIL.n734 33.9308
R553 VTAIL.n629 VTAIL.n628 33.9308
R554 VTAIL.n525 VTAIL.n524 33.9308
R555 VTAIL.n419 VTAIL.n418 33.9308
R556 VTAIL.n839 VTAIL.n735 31.4789
R557 VTAIL.n419 VTAIL.n315 31.4789
R558 VTAIL.n791 VTAIL.n758 13.1884
R559 VTAIL.n57 VTAIL.n24 13.1884
R560 VTAIL.n161 VTAIL.n128 13.1884
R561 VTAIL.n267 VTAIL.n234 13.1884
R562 VTAIL.n656 VTAIL.n654 13.1884
R563 VTAIL.n550 VTAIL.n548 13.1884
R564 VTAIL.n446 VTAIL.n444 13.1884
R565 VTAIL.n340 VTAIL.n338 13.1884
R566 VTAIL.n792 VTAIL.n760 12.8005
R567 VTAIL.n796 VTAIL.n795 12.8005
R568 VTAIL.n836 VTAIL.n736 12.8005
R569 VTAIL.n58 VTAIL.n26 12.8005
R570 VTAIL.n62 VTAIL.n61 12.8005
R571 VTAIL.n102 VTAIL.n2 12.8005
R572 VTAIL.n162 VTAIL.n130 12.8005
R573 VTAIL.n166 VTAIL.n165 12.8005
R574 VTAIL.n206 VTAIL.n106 12.8005
R575 VTAIL.n268 VTAIL.n236 12.8005
R576 VTAIL.n272 VTAIL.n271 12.8005
R577 VTAIL.n312 VTAIL.n212 12.8005
R578 VTAIL.n732 VTAIL.n632 12.8005
R579 VTAIL.n692 VTAIL.n691 12.8005
R580 VTAIL.n688 VTAIL.n687 12.8005
R581 VTAIL.n626 VTAIL.n526 12.8005
R582 VTAIL.n586 VTAIL.n585 12.8005
R583 VTAIL.n582 VTAIL.n581 12.8005
R584 VTAIL.n522 VTAIL.n422 12.8005
R585 VTAIL.n482 VTAIL.n481 12.8005
R586 VTAIL.n478 VTAIL.n477 12.8005
R587 VTAIL.n416 VTAIL.n316 12.8005
R588 VTAIL.n376 VTAIL.n375 12.8005
R589 VTAIL.n372 VTAIL.n371 12.8005
R590 VTAIL.n787 VTAIL.n786 12.0247
R591 VTAIL.n799 VTAIL.n756 12.0247
R592 VTAIL.n835 VTAIL.n738 12.0247
R593 VTAIL.n53 VTAIL.n52 12.0247
R594 VTAIL.n65 VTAIL.n22 12.0247
R595 VTAIL.n101 VTAIL.n4 12.0247
R596 VTAIL.n157 VTAIL.n156 12.0247
R597 VTAIL.n169 VTAIL.n126 12.0247
R598 VTAIL.n205 VTAIL.n108 12.0247
R599 VTAIL.n263 VTAIL.n262 12.0247
R600 VTAIL.n275 VTAIL.n232 12.0247
R601 VTAIL.n311 VTAIL.n214 12.0247
R602 VTAIL.n731 VTAIL.n634 12.0247
R603 VTAIL.n695 VTAIL.n652 12.0247
R604 VTAIL.n684 VTAIL.n657 12.0247
R605 VTAIL.n625 VTAIL.n528 12.0247
R606 VTAIL.n589 VTAIL.n546 12.0247
R607 VTAIL.n578 VTAIL.n551 12.0247
R608 VTAIL.n521 VTAIL.n424 12.0247
R609 VTAIL.n485 VTAIL.n442 12.0247
R610 VTAIL.n474 VTAIL.n447 12.0247
R611 VTAIL.n415 VTAIL.n318 12.0247
R612 VTAIL.n379 VTAIL.n336 12.0247
R613 VTAIL.n368 VTAIL.n341 12.0247
R614 VTAIL.n785 VTAIL.n762 11.249
R615 VTAIL.n800 VTAIL.n754 11.249
R616 VTAIL.n832 VTAIL.n831 11.249
R617 VTAIL.n51 VTAIL.n28 11.249
R618 VTAIL.n66 VTAIL.n20 11.249
R619 VTAIL.n98 VTAIL.n97 11.249
R620 VTAIL.n155 VTAIL.n132 11.249
R621 VTAIL.n170 VTAIL.n124 11.249
R622 VTAIL.n202 VTAIL.n201 11.249
R623 VTAIL.n261 VTAIL.n238 11.249
R624 VTAIL.n276 VTAIL.n230 11.249
R625 VTAIL.n308 VTAIL.n307 11.249
R626 VTAIL.n728 VTAIL.n727 11.249
R627 VTAIL.n696 VTAIL.n650 11.249
R628 VTAIL.n683 VTAIL.n660 11.249
R629 VTAIL.n622 VTAIL.n621 11.249
R630 VTAIL.n590 VTAIL.n544 11.249
R631 VTAIL.n577 VTAIL.n554 11.249
R632 VTAIL.n518 VTAIL.n517 11.249
R633 VTAIL.n486 VTAIL.n440 11.249
R634 VTAIL.n473 VTAIL.n450 11.249
R635 VTAIL.n412 VTAIL.n411 11.249
R636 VTAIL.n380 VTAIL.n334 11.249
R637 VTAIL.n367 VTAIL.n344 11.249
R638 VTAIL.n782 VTAIL.n781 10.4732
R639 VTAIL.n804 VTAIL.n803 10.4732
R640 VTAIL.n828 VTAIL.n740 10.4732
R641 VTAIL.n48 VTAIL.n47 10.4732
R642 VTAIL.n70 VTAIL.n69 10.4732
R643 VTAIL.n94 VTAIL.n6 10.4732
R644 VTAIL.n152 VTAIL.n151 10.4732
R645 VTAIL.n174 VTAIL.n173 10.4732
R646 VTAIL.n198 VTAIL.n110 10.4732
R647 VTAIL.n258 VTAIL.n257 10.4732
R648 VTAIL.n280 VTAIL.n279 10.4732
R649 VTAIL.n304 VTAIL.n216 10.4732
R650 VTAIL.n724 VTAIL.n636 10.4732
R651 VTAIL.n700 VTAIL.n699 10.4732
R652 VTAIL.n680 VTAIL.n679 10.4732
R653 VTAIL.n618 VTAIL.n530 10.4732
R654 VTAIL.n594 VTAIL.n593 10.4732
R655 VTAIL.n574 VTAIL.n573 10.4732
R656 VTAIL.n514 VTAIL.n426 10.4732
R657 VTAIL.n490 VTAIL.n489 10.4732
R658 VTAIL.n470 VTAIL.n469 10.4732
R659 VTAIL.n408 VTAIL.n320 10.4732
R660 VTAIL.n384 VTAIL.n383 10.4732
R661 VTAIL.n364 VTAIL.n363 10.4732
R662 VTAIL.n770 VTAIL.n769 10.2747
R663 VTAIL.n36 VTAIL.n35 10.2747
R664 VTAIL.n140 VTAIL.n139 10.2747
R665 VTAIL.n246 VTAIL.n245 10.2747
R666 VTAIL.n668 VTAIL.n667 10.2747
R667 VTAIL.n562 VTAIL.n561 10.2747
R668 VTAIL.n458 VTAIL.n457 10.2747
R669 VTAIL.n352 VTAIL.n351 10.2747
R670 VTAIL.n778 VTAIL.n764 9.69747
R671 VTAIL.n807 VTAIL.n752 9.69747
R672 VTAIL.n827 VTAIL.n742 9.69747
R673 VTAIL.n44 VTAIL.n30 9.69747
R674 VTAIL.n73 VTAIL.n18 9.69747
R675 VTAIL.n93 VTAIL.n8 9.69747
R676 VTAIL.n148 VTAIL.n134 9.69747
R677 VTAIL.n177 VTAIL.n122 9.69747
R678 VTAIL.n197 VTAIL.n112 9.69747
R679 VTAIL.n254 VTAIL.n240 9.69747
R680 VTAIL.n283 VTAIL.n228 9.69747
R681 VTAIL.n303 VTAIL.n218 9.69747
R682 VTAIL.n723 VTAIL.n638 9.69747
R683 VTAIL.n703 VTAIL.n648 9.69747
R684 VTAIL.n676 VTAIL.n662 9.69747
R685 VTAIL.n617 VTAIL.n532 9.69747
R686 VTAIL.n597 VTAIL.n542 9.69747
R687 VTAIL.n570 VTAIL.n556 9.69747
R688 VTAIL.n513 VTAIL.n428 9.69747
R689 VTAIL.n493 VTAIL.n438 9.69747
R690 VTAIL.n466 VTAIL.n452 9.69747
R691 VTAIL.n407 VTAIL.n322 9.69747
R692 VTAIL.n387 VTAIL.n332 9.69747
R693 VTAIL.n360 VTAIL.n346 9.69747
R694 VTAIL.n834 VTAIL.n736 9.45567
R695 VTAIL.n100 VTAIL.n2 9.45567
R696 VTAIL.n204 VTAIL.n106 9.45567
R697 VTAIL.n310 VTAIL.n212 9.45567
R698 VTAIL.n730 VTAIL.n632 9.45567
R699 VTAIL.n624 VTAIL.n526 9.45567
R700 VTAIL.n520 VTAIL.n422 9.45567
R701 VTAIL.n414 VTAIL.n316 9.45567
R702 VTAIL.n817 VTAIL.n816 9.3005
R703 VTAIL.n819 VTAIL.n818 9.3005
R704 VTAIL.n744 VTAIL.n743 9.3005
R705 VTAIL.n825 VTAIL.n824 9.3005
R706 VTAIL.n827 VTAIL.n826 9.3005
R707 VTAIL.n740 VTAIL.n739 9.3005
R708 VTAIL.n833 VTAIL.n832 9.3005
R709 VTAIL.n835 VTAIL.n834 9.3005
R710 VTAIL.n811 VTAIL.n810 9.3005
R711 VTAIL.n809 VTAIL.n808 9.3005
R712 VTAIL.n752 VTAIL.n751 9.3005
R713 VTAIL.n803 VTAIL.n802 9.3005
R714 VTAIL.n801 VTAIL.n800 9.3005
R715 VTAIL.n756 VTAIL.n755 9.3005
R716 VTAIL.n795 VTAIL.n794 9.3005
R717 VTAIL.n768 VTAIL.n767 9.3005
R718 VTAIL.n775 VTAIL.n774 9.3005
R719 VTAIL.n777 VTAIL.n776 9.3005
R720 VTAIL.n764 VTAIL.n763 9.3005
R721 VTAIL.n783 VTAIL.n782 9.3005
R722 VTAIL.n785 VTAIL.n784 9.3005
R723 VTAIL.n786 VTAIL.n759 9.3005
R724 VTAIL.n793 VTAIL.n792 9.3005
R725 VTAIL.n748 VTAIL.n747 9.3005
R726 VTAIL.n83 VTAIL.n82 9.3005
R727 VTAIL.n85 VTAIL.n84 9.3005
R728 VTAIL.n10 VTAIL.n9 9.3005
R729 VTAIL.n91 VTAIL.n90 9.3005
R730 VTAIL.n93 VTAIL.n92 9.3005
R731 VTAIL.n6 VTAIL.n5 9.3005
R732 VTAIL.n99 VTAIL.n98 9.3005
R733 VTAIL.n101 VTAIL.n100 9.3005
R734 VTAIL.n77 VTAIL.n76 9.3005
R735 VTAIL.n75 VTAIL.n74 9.3005
R736 VTAIL.n18 VTAIL.n17 9.3005
R737 VTAIL.n69 VTAIL.n68 9.3005
R738 VTAIL.n67 VTAIL.n66 9.3005
R739 VTAIL.n22 VTAIL.n21 9.3005
R740 VTAIL.n61 VTAIL.n60 9.3005
R741 VTAIL.n34 VTAIL.n33 9.3005
R742 VTAIL.n41 VTAIL.n40 9.3005
R743 VTAIL.n43 VTAIL.n42 9.3005
R744 VTAIL.n30 VTAIL.n29 9.3005
R745 VTAIL.n49 VTAIL.n48 9.3005
R746 VTAIL.n51 VTAIL.n50 9.3005
R747 VTAIL.n52 VTAIL.n25 9.3005
R748 VTAIL.n59 VTAIL.n58 9.3005
R749 VTAIL.n14 VTAIL.n13 9.3005
R750 VTAIL.n187 VTAIL.n186 9.3005
R751 VTAIL.n189 VTAIL.n188 9.3005
R752 VTAIL.n114 VTAIL.n113 9.3005
R753 VTAIL.n195 VTAIL.n194 9.3005
R754 VTAIL.n197 VTAIL.n196 9.3005
R755 VTAIL.n110 VTAIL.n109 9.3005
R756 VTAIL.n203 VTAIL.n202 9.3005
R757 VTAIL.n205 VTAIL.n204 9.3005
R758 VTAIL.n181 VTAIL.n180 9.3005
R759 VTAIL.n179 VTAIL.n178 9.3005
R760 VTAIL.n122 VTAIL.n121 9.3005
R761 VTAIL.n173 VTAIL.n172 9.3005
R762 VTAIL.n171 VTAIL.n170 9.3005
R763 VTAIL.n126 VTAIL.n125 9.3005
R764 VTAIL.n165 VTAIL.n164 9.3005
R765 VTAIL.n138 VTAIL.n137 9.3005
R766 VTAIL.n145 VTAIL.n144 9.3005
R767 VTAIL.n147 VTAIL.n146 9.3005
R768 VTAIL.n134 VTAIL.n133 9.3005
R769 VTAIL.n153 VTAIL.n152 9.3005
R770 VTAIL.n155 VTAIL.n154 9.3005
R771 VTAIL.n156 VTAIL.n129 9.3005
R772 VTAIL.n163 VTAIL.n162 9.3005
R773 VTAIL.n118 VTAIL.n117 9.3005
R774 VTAIL.n293 VTAIL.n292 9.3005
R775 VTAIL.n295 VTAIL.n294 9.3005
R776 VTAIL.n220 VTAIL.n219 9.3005
R777 VTAIL.n301 VTAIL.n300 9.3005
R778 VTAIL.n303 VTAIL.n302 9.3005
R779 VTAIL.n216 VTAIL.n215 9.3005
R780 VTAIL.n309 VTAIL.n308 9.3005
R781 VTAIL.n311 VTAIL.n310 9.3005
R782 VTAIL.n287 VTAIL.n286 9.3005
R783 VTAIL.n285 VTAIL.n284 9.3005
R784 VTAIL.n228 VTAIL.n227 9.3005
R785 VTAIL.n279 VTAIL.n278 9.3005
R786 VTAIL.n277 VTAIL.n276 9.3005
R787 VTAIL.n232 VTAIL.n231 9.3005
R788 VTAIL.n271 VTAIL.n270 9.3005
R789 VTAIL.n244 VTAIL.n243 9.3005
R790 VTAIL.n251 VTAIL.n250 9.3005
R791 VTAIL.n253 VTAIL.n252 9.3005
R792 VTAIL.n240 VTAIL.n239 9.3005
R793 VTAIL.n259 VTAIL.n258 9.3005
R794 VTAIL.n261 VTAIL.n260 9.3005
R795 VTAIL.n262 VTAIL.n235 9.3005
R796 VTAIL.n269 VTAIL.n268 9.3005
R797 VTAIL.n224 VTAIL.n223 9.3005
R798 VTAIL.n731 VTAIL.n730 9.3005
R799 VTAIL.n729 VTAIL.n728 9.3005
R800 VTAIL.n636 VTAIL.n635 9.3005
R801 VTAIL.n723 VTAIL.n722 9.3005
R802 VTAIL.n721 VTAIL.n720 9.3005
R803 VTAIL.n640 VTAIL.n639 9.3005
R804 VTAIL.n715 VTAIL.n714 9.3005
R805 VTAIL.n713 VTAIL.n712 9.3005
R806 VTAIL.n644 VTAIL.n643 9.3005
R807 VTAIL.n707 VTAIL.n706 9.3005
R808 VTAIL.n705 VTAIL.n704 9.3005
R809 VTAIL.n648 VTAIL.n647 9.3005
R810 VTAIL.n699 VTAIL.n698 9.3005
R811 VTAIL.n697 VTAIL.n696 9.3005
R812 VTAIL.n652 VTAIL.n651 9.3005
R813 VTAIL.n691 VTAIL.n690 9.3005
R814 VTAIL.n689 VTAIL.n688 9.3005
R815 VTAIL.n657 VTAIL.n655 9.3005
R816 VTAIL.n683 VTAIL.n682 9.3005
R817 VTAIL.n681 VTAIL.n680 9.3005
R818 VTAIL.n662 VTAIL.n661 9.3005
R819 VTAIL.n675 VTAIL.n674 9.3005
R820 VTAIL.n673 VTAIL.n672 9.3005
R821 VTAIL.n666 VTAIL.n665 9.3005
R822 VTAIL.n560 VTAIL.n559 9.3005
R823 VTAIL.n567 VTAIL.n566 9.3005
R824 VTAIL.n569 VTAIL.n568 9.3005
R825 VTAIL.n556 VTAIL.n555 9.3005
R826 VTAIL.n575 VTAIL.n574 9.3005
R827 VTAIL.n577 VTAIL.n576 9.3005
R828 VTAIL.n551 VTAIL.n549 9.3005
R829 VTAIL.n583 VTAIL.n582 9.3005
R830 VTAIL.n609 VTAIL.n608 9.3005
R831 VTAIL.n534 VTAIL.n533 9.3005
R832 VTAIL.n615 VTAIL.n614 9.3005
R833 VTAIL.n617 VTAIL.n616 9.3005
R834 VTAIL.n530 VTAIL.n529 9.3005
R835 VTAIL.n623 VTAIL.n622 9.3005
R836 VTAIL.n625 VTAIL.n624 9.3005
R837 VTAIL.n607 VTAIL.n606 9.3005
R838 VTAIL.n538 VTAIL.n537 9.3005
R839 VTAIL.n601 VTAIL.n600 9.3005
R840 VTAIL.n599 VTAIL.n598 9.3005
R841 VTAIL.n542 VTAIL.n541 9.3005
R842 VTAIL.n593 VTAIL.n592 9.3005
R843 VTAIL.n591 VTAIL.n590 9.3005
R844 VTAIL.n546 VTAIL.n545 9.3005
R845 VTAIL.n585 VTAIL.n584 9.3005
R846 VTAIL.n456 VTAIL.n455 9.3005
R847 VTAIL.n463 VTAIL.n462 9.3005
R848 VTAIL.n465 VTAIL.n464 9.3005
R849 VTAIL.n452 VTAIL.n451 9.3005
R850 VTAIL.n471 VTAIL.n470 9.3005
R851 VTAIL.n473 VTAIL.n472 9.3005
R852 VTAIL.n447 VTAIL.n445 9.3005
R853 VTAIL.n479 VTAIL.n478 9.3005
R854 VTAIL.n505 VTAIL.n504 9.3005
R855 VTAIL.n430 VTAIL.n429 9.3005
R856 VTAIL.n511 VTAIL.n510 9.3005
R857 VTAIL.n513 VTAIL.n512 9.3005
R858 VTAIL.n426 VTAIL.n425 9.3005
R859 VTAIL.n519 VTAIL.n518 9.3005
R860 VTAIL.n521 VTAIL.n520 9.3005
R861 VTAIL.n503 VTAIL.n502 9.3005
R862 VTAIL.n434 VTAIL.n433 9.3005
R863 VTAIL.n497 VTAIL.n496 9.3005
R864 VTAIL.n495 VTAIL.n494 9.3005
R865 VTAIL.n438 VTAIL.n437 9.3005
R866 VTAIL.n489 VTAIL.n488 9.3005
R867 VTAIL.n487 VTAIL.n486 9.3005
R868 VTAIL.n442 VTAIL.n441 9.3005
R869 VTAIL.n481 VTAIL.n480 9.3005
R870 VTAIL.n350 VTAIL.n349 9.3005
R871 VTAIL.n357 VTAIL.n356 9.3005
R872 VTAIL.n359 VTAIL.n358 9.3005
R873 VTAIL.n346 VTAIL.n345 9.3005
R874 VTAIL.n365 VTAIL.n364 9.3005
R875 VTAIL.n367 VTAIL.n366 9.3005
R876 VTAIL.n341 VTAIL.n339 9.3005
R877 VTAIL.n373 VTAIL.n372 9.3005
R878 VTAIL.n399 VTAIL.n398 9.3005
R879 VTAIL.n324 VTAIL.n323 9.3005
R880 VTAIL.n405 VTAIL.n404 9.3005
R881 VTAIL.n407 VTAIL.n406 9.3005
R882 VTAIL.n320 VTAIL.n319 9.3005
R883 VTAIL.n413 VTAIL.n412 9.3005
R884 VTAIL.n415 VTAIL.n414 9.3005
R885 VTAIL.n397 VTAIL.n396 9.3005
R886 VTAIL.n328 VTAIL.n327 9.3005
R887 VTAIL.n391 VTAIL.n390 9.3005
R888 VTAIL.n389 VTAIL.n388 9.3005
R889 VTAIL.n332 VTAIL.n331 9.3005
R890 VTAIL.n383 VTAIL.n382 9.3005
R891 VTAIL.n381 VTAIL.n380 9.3005
R892 VTAIL.n336 VTAIL.n335 9.3005
R893 VTAIL.n375 VTAIL.n374 9.3005
R894 VTAIL.n777 VTAIL.n766 8.92171
R895 VTAIL.n808 VTAIL.n750 8.92171
R896 VTAIL.n824 VTAIL.n823 8.92171
R897 VTAIL.n43 VTAIL.n32 8.92171
R898 VTAIL.n74 VTAIL.n16 8.92171
R899 VTAIL.n90 VTAIL.n89 8.92171
R900 VTAIL.n147 VTAIL.n136 8.92171
R901 VTAIL.n178 VTAIL.n120 8.92171
R902 VTAIL.n194 VTAIL.n193 8.92171
R903 VTAIL.n253 VTAIL.n242 8.92171
R904 VTAIL.n284 VTAIL.n226 8.92171
R905 VTAIL.n300 VTAIL.n299 8.92171
R906 VTAIL.n720 VTAIL.n719 8.92171
R907 VTAIL.n704 VTAIL.n646 8.92171
R908 VTAIL.n675 VTAIL.n664 8.92171
R909 VTAIL.n614 VTAIL.n613 8.92171
R910 VTAIL.n598 VTAIL.n540 8.92171
R911 VTAIL.n569 VTAIL.n558 8.92171
R912 VTAIL.n510 VTAIL.n509 8.92171
R913 VTAIL.n494 VTAIL.n436 8.92171
R914 VTAIL.n465 VTAIL.n454 8.92171
R915 VTAIL.n404 VTAIL.n403 8.92171
R916 VTAIL.n388 VTAIL.n330 8.92171
R917 VTAIL.n359 VTAIL.n348 8.92171
R918 VTAIL.n774 VTAIL.n773 8.14595
R919 VTAIL.n812 VTAIL.n811 8.14595
R920 VTAIL.n820 VTAIL.n744 8.14595
R921 VTAIL.n40 VTAIL.n39 8.14595
R922 VTAIL.n78 VTAIL.n77 8.14595
R923 VTAIL.n86 VTAIL.n10 8.14595
R924 VTAIL.n144 VTAIL.n143 8.14595
R925 VTAIL.n182 VTAIL.n181 8.14595
R926 VTAIL.n190 VTAIL.n114 8.14595
R927 VTAIL.n250 VTAIL.n249 8.14595
R928 VTAIL.n288 VTAIL.n287 8.14595
R929 VTAIL.n296 VTAIL.n220 8.14595
R930 VTAIL.n716 VTAIL.n640 8.14595
R931 VTAIL.n708 VTAIL.n707 8.14595
R932 VTAIL.n672 VTAIL.n671 8.14595
R933 VTAIL.n610 VTAIL.n534 8.14595
R934 VTAIL.n602 VTAIL.n601 8.14595
R935 VTAIL.n566 VTAIL.n565 8.14595
R936 VTAIL.n506 VTAIL.n430 8.14595
R937 VTAIL.n498 VTAIL.n497 8.14595
R938 VTAIL.n462 VTAIL.n461 8.14595
R939 VTAIL.n400 VTAIL.n324 8.14595
R940 VTAIL.n392 VTAIL.n391 8.14595
R941 VTAIL.n356 VTAIL.n355 8.14595
R942 VTAIL.n770 VTAIL.n768 7.3702
R943 VTAIL.n815 VTAIL.n748 7.3702
R944 VTAIL.n819 VTAIL.n746 7.3702
R945 VTAIL.n36 VTAIL.n34 7.3702
R946 VTAIL.n81 VTAIL.n14 7.3702
R947 VTAIL.n85 VTAIL.n12 7.3702
R948 VTAIL.n140 VTAIL.n138 7.3702
R949 VTAIL.n185 VTAIL.n118 7.3702
R950 VTAIL.n189 VTAIL.n116 7.3702
R951 VTAIL.n246 VTAIL.n244 7.3702
R952 VTAIL.n291 VTAIL.n224 7.3702
R953 VTAIL.n295 VTAIL.n222 7.3702
R954 VTAIL.n715 VTAIL.n642 7.3702
R955 VTAIL.n711 VTAIL.n644 7.3702
R956 VTAIL.n668 VTAIL.n666 7.3702
R957 VTAIL.n609 VTAIL.n536 7.3702
R958 VTAIL.n605 VTAIL.n538 7.3702
R959 VTAIL.n562 VTAIL.n560 7.3702
R960 VTAIL.n505 VTAIL.n432 7.3702
R961 VTAIL.n501 VTAIL.n434 7.3702
R962 VTAIL.n458 VTAIL.n456 7.3702
R963 VTAIL.n399 VTAIL.n326 7.3702
R964 VTAIL.n395 VTAIL.n328 7.3702
R965 VTAIL.n352 VTAIL.n350 7.3702
R966 VTAIL.n816 VTAIL.n815 6.59444
R967 VTAIL.n816 VTAIL.n746 6.59444
R968 VTAIL.n82 VTAIL.n81 6.59444
R969 VTAIL.n82 VTAIL.n12 6.59444
R970 VTAIL.n186 VTAIL.n185 6.59444
R971 VTAIL.n186 VTAIL.n116 6.59444
R972 VTAIL.n292 VTAIL.n291 6.59444
R973 VTAIL.n292 VTAIL.n222 6.59444
R974 VTAIL.n712 VTAIL.n642 6.59444
R975 VTAIL.n712 VTAIL.n711 6.59444
R976 VTAIL.n606 VTAIL.n536 6.59444
R977 VTAIL.n606 VTAIL.n605 6.59444
R978 VTAIL.n502 VTAIL.n432 6.59444
R979 VTAIL.n502 VTAIL.n501 6.59444
R980 VTAIL.n396 VTAIL.n326 6.59444
R981 VTAIL.n396 VTAIL.n395 6.59444
R982 VTAIL.n773 VTAIL.n768 5.81868
R983 VTAIL.n812 VTAIL.n748 5.81868
R984 VTAIL.n820 VTAIL.n819 5.81868
R985 VTAIL.n39 VTAIL.n34 5.81868
R986 VTAIL.n78 VTAIL.n14 5.81868
R987 VTAIL.n86 VTAIL.n85 5.81868
R988 VTAIL.n143 VTAIL.n138 5.81868
R989 VTAIL.n182 VTAIL.n118 5.81868
R990 VTAIL.n190 VTAIL.n189 5.81868
R991 VTAIL.n249 VTAIL.n244 5.81868
R992 VTAIL.n288 VTAIL.n224 5.81868
R993 VTAIL.n296 VTAIL.n295 5.81868
R994 VTAIL.n716 VTAIL.n715 5.81868
R995 VTAIL.n708 VTAIL.n644 5.81868
R996 VTAIL.n671 VTAIL.n666 5.81868
R997 VTAIL.n610 VTAIL.n609 5.81868
R998 VTAIL.n602 VTAIL.n538 5.81868
R999 VTAIL.n565 VTAIL.n560 5.81868
R1000 VTAIL.n506 VTAIL.n505 5.81868
R1001 VTAIL.n498 VTAIL.n434 5.81868
R1002 VTAIL.n461 VTAIL.n456 5.81868
R1003 VTAIL.n400 VTAIL.n399 5.81868
R1004 VTAIL.n392 VTAIL.n328 5.81868
R1005 VTAIL.n355 VTAIL.n350 5.81868
R1006 VTAIL.n774 VTAIL.n766 5.04292
R1007 VTAIL.n811 VTAIL.n750 5.04292
R1008 VTAIL.n823 VTAIL.n744 5.04292
R1009 VTAIL.n40 VTAIL.n32 5.04292
R1010 VTAIL.n77 VTAIL.n16 5.04292
R1011 VTAIL.n89 VTAIL.n10 5.04292
R1012 VTAIL.n144 VTAIL.n136 5.04292
R1013 VTAIL.n181 VTAIL.n120 5.04292
R1014 VTAIL.n193 VTAIL.n114 5.04292
R1015 VTAIL.n250 VTAIL.n242 5.04292
R1016 VTAIL.n287 VTAIL.n226 5.04292
R1017 VTAIL.n299 VTAIL.n220 5.04292
R1018 VTAIL.n719 VTAIL.n640 5.04292
R1019 VTAIL.n707 VTAIL.n646 5.04292
R1020 VTAIL.n672 VTAIL.n664 5.04292
R1021 VTAIL.n613 VTAIL.n534 5.04292
R1022 VTAIL.n601 VTAIL.n540 5.04292
R1023 VTAIL.n566 VTAIL.n558 5.04292
R1024 VTAIL.n509 VTAIL.n430 5.04292
R1025 VTAIL.n497 VTAIL.n436 5.04292
R1026 VTAIL.n462 VTAIL.n454 5.04292
R1027 VTAIL.n403 VTAIL.n324 5.04292
R1028 VTAIL.n391 VTAIL.n330 5.04292
R1029 VTAIL.n356 VTAIL.n348 5.04292
R1030 VTAIL.n778 VTAIL.n777 4.26717
R1031 VTAIL.n808 VTAIL.n807 4.26717
R1032 VTAIL.n824 VTAIL.n742 4.26717
R1033 VTAIL.n44 VTAIL.n43 4.26717
R1034 VTAIL.n74 VTAIL.n73 4.26717
R1035 VTAIL.n90 VTAIL.n8 4.26717
R1036 VTAIL.n148 VTAIL.n147 4.26717
R1037 VTAIL.n178 VTAIL.n177 4.26717
R1038 VTAIL.n194 VTAIL.n112 4.26717
R1039 VTAIL.n254 VTAIL.n253 4.26717
R1040 VTAIL.n284 VTAIL.n283 4.26717
R1041 VTAIL.n300 VTAIL.n218 4.26717
R1042 VTAIL.n720 VTAIL.n638 4.26717
R1043 VTAIL.n704 VTAIL.n703 4.26717
R1044 VTAIL.n676 VTAIL.n675 4.26717
R1045 VTAIL.n614 VTAIL.n532 4.26717
R1046 VTAIL.n598 VTAIL.n597 4.26717
R1047 VTAIL.n570 VTAIL.n569 4.26717
R1048 VTAIL.n510 VTAIL.n428 4.26717
R1049 VTAIL.n494 VTAIL.n493 4.26717
R1050 VTAIL.n466 VTAIL.n465 4.26717
R1051 VTAIL.n404 VTAIL.n322 4.26717
R1052 VTAIL.n388 VTAIL.n387 4.26717
R1053 VTAIL.n360 VTAIL.n359 4.26717
R1054 VTAIL.n781 VTAIL.n764 3.49141
R1055 VTAIL.n804 VTAIL.n752 3.49141
R1056 VTAIL.n828 VTAIL.n827 3.49141
R1057 VTAIL.n47 VTAIL.n30 3.49141
R1058 VTAIL.n70 VTAIL.n18 3.49141
R1059 VTAIL.n94 VTAIL.n93 3.49141
R1060 VTAIL.n151 VTAIL.n134 3.49141
R1061 VTAIL.n174 VTAIL.n122 3.49141
R1062 VTAIL.n198 VTAIL.n197 3.49141
R1063 VTAIL.n257 VTAIL.n240 3.49141
R1064 VTAIL.n280 VTAIL.n228 3.49141
R1065 VTAIL.n304 VTAIL.n303 3.49141
R1066 VTAIL.n724 VTAIL.n723 3.49141
R1067 VTAIL.n700 VTAIL.n648 3.49141
R1068 VTAIL.n679 VTAIL.n662 3.49141
R1069 VTAIL.n618 VTAIL.n617 3.49141
R1070 VTAIL.n594 VTAIL.n542 3.49141
R1071 VTAIL.n573 VTAIL.n556 3.49141
R1072 VTAIL.n514 VTAIL.n513 3.49141
R1073 VTAIL.n490 VTAIL.n438 3.49141
R1074 VTAIL.n469 VTAIL.n452 3.49141
R1075 VTAIL.n408 VTAIL.n407 3.49141
R1076 VTAIL.n384 VTAIL.n332 3.49141
R1077 VTAIL.n363 VTAIL.n346 3.49141
R1078 VTAIL.n421 VTAIL.n419 2.98326
R1079 VTAIL.n525 VTAIL.n421 2.98326
R1080 VTAIL.n631 VTAIL.n629 2.98326
R1081 VTAIL.n735 VTAIL.n631 2.98326
R1082 VTAIL.n315 VTAIL.n211 2.98326
R1083 VTAIL.n211 VTAIL.n209 2.98326
R1084 VTAIL.n105 VTAIL.n1 2.98326
R1085 VTAIL VTAIL.n839 2.92507
R1086 VTAIL.n769 VTAIL.n767 2.84303
R1087 VTAIL.n35 VTAIL.n33 2.84303
R1088 VTAIL.n139 VTAIL.n137 2.84303
R1089 VTAIL.n245 VTAIL.n243 2.84303
R1090 VTAIL.n667 VTAIL.n665 2.84303
R1091 VTAIL.n561 VTAIL.n559 2.84303
R1092 VTAIL.n457 VTAIL.n455 2.84303
R1093 VTAIL.n351 VTAIL.n349 2.84303
R1094 VTAIL.n782 VTAIL.n762 2.71565
R1095 VTAIL.n803 VTAIL.n754 2.71565
R1096 VTAIL.n831 VTAIL.n740 2.71565
R1097 VTAIL.n48 VTAIL.n28 2.71565
R1098 VTAIL.n69 VTAIL.n20 2.71565
R1099 VTAIL.n97 VTAIL.n6 2.71565
R1100 VTAIL.n152 VTAIL.n132 2.71565
R1101 VTAIL.n173 VTAIL.n124 2.71565
R1102 VTAIL.n201 VTAIL.n110 2.71565
R1103 VTAIL.n258 VTAIL.n238 2.71565
R1104 VTAIL.n279 VTAIL.n230 2.71565
R1105 VTAIL.n307 VTAIL.n216 2.71565
R1106 VTAIL.n727 VTAIL.n636 2.71565
R1107 VTAIL.n699 VTAIL.n650 2.71565
R1108 VTAIL.n680 VTAIL.n660 2.71565
R1109 VTAIL.n621 VTAIL.n530 2.71565
R1110 VTAIL.n593 VTAIL.n544 2.71565
R1111 VTAIL.n574 VTAIL.n554 2.71565
R1112 VTAIL.n517 VTAIL.n426 2.71565
R1113 VTAIL.n489 VTAIL.n440 2.71565
R1114 VTAIL.n470 VTAIL.n450 2.71565
R1115 VTAIL.n411 VTAIL.n320 2.71565
R1116 VTAIL.n383 VTAIL.n334 2.71565
R1117 VTAIL.n364 VTAIL.n344 2.71565
R1118 VTAIL.n787 VTAIL.n785 1.93989
R1119 VTAIL.n800 VTAIL.n799 1.93989
R1120 VTAIL.n832 VTAIL.n738 1.93989
R1121 VTAIL.n53 VTAIL.n51 1.93989
R1122 VTAIL.n66 VTAIL.n65 1.93989
R1123 VTAIL.n98 VTAIL.n4 1.93989
R1124 VTAIL.n157 VTAIL.n155 1.93989
R1125 VTAIL.n170 VTAIL.n169 1.93989
R1126 VTAIL.n202 VTAIL.n108 1.93989
R1127 VTAIL.n263 VTAIL.n261 1.93989
R1128 VTAIL.n276 VTAIL.n275 1.93989
R1129 VTAIL.n308 VTAIL.n214 1.93989
R1130 VTAIL.n728 VTAIL.n634 1.93989
R1131 VTAIL.n696 VTAIL.n695 1.93989
R1132 VTAIL.n684 VTAIL.n683 1.93989
R1133 VTAIL.n622 VTAIL.n528 1.93989
R1134 VTAIL.n590 VTAIL.n589 1.93989
R1135 VTAIL.n578 VTAIL.n577 1.93989
R1136 VTAIL.n518 VTAIL.n424 1.93989
R1137 VTAIL.n486 VTAIL.n485 1.93989
R1138 VTAIL.n474 VTAIL.n473 1.93989
R1139 VTAIL.n412 VTAIL.n318 1.93989
R1140 VTAIL.n380 VTAIL.n379 1.93989
R1141 VTAIL.n368 VTAIL.n367 1.93989
R1142 VTAIL.n786 VTAIL.n760 1.16414
R1143 VTAIL.n796 VTAIL.n756 1.16414
R1144 VTAIL.n836 VTAIL.n835 1.16414
R1145 VTAIL.n52 VTAIL.n26 1.16414
R1146 VTAIL.n62 VTAIL.n22 1.16414
R1147 VTAIL.n102 VTAIL.n101 1.16414
R1148 VTAIL.n156 VTAIL.n130 1.16414
R1149 VTAIL.n166 VTAIL.n126 1.16414
R1150 VTAIL.n206 VTAIL.n205 1.16414
R1151 VTAIL.n262 VTAIL.n236 1.16414
R1152 VTAIL.n272 VTAIL.n232 1.16414
R1153 VTAIL.n312 VTAIL.n311 1.16414
R1154 VTAIL.n732 VTAIL.n731 1.16414
R1155 VTAIL.n692 VTAIL.n652 1.16414
R1156 VTAIL.n687 VTAIL.n657 1.16414
R1157 VTAIL.n626 VTAIL.n625 1.16414
R1158 VTAIL.n586 VTAIL.n546 1.16414
R1159 VTAIL.n581 VTAIL.n551 1.16414
R1160 VTAIL.n522 VTAIL.n521 1.16414
R1161 VTAIL.n482 VTAIL.n442 1.16414
R1162 VTAIL.n477 VTAIL.n447 1.16414
R1163 VTAIL.n416 VTAIL.n415 1.16414
R1164 VTAIL.n376 VTAIL.n336 1.16414
R1165 VTAIL.n371 VTAIL.n341 1.16414
R1166 VTAIL.n0 VTAIL.t11 1.05876
R1167 VTAIL.n0 VTAIL.t12 1.05876
R1168 VTAIL.n210 VTAIL.t5 1.05876
R1169 VTAIL.n210 VTAIL.t0 1.05876
R1170 VTAIL.n630 VTAIL.t4 1.05876
R1171 VTAIL.n630 VTAIL.t3 1.05876
R1172 VTAIL.n420 VTAIL.t8 1.05876
R1173 VTAIL.n420 VTAIL.t14 1.05876
R1174 VTAIL.n629 VTAIL.n525 0.470328
R1175 VTAIL.n209 VTAIL.n105 0.470328
R1176 VTAIL.n792 VTAIL.n791 0.388379
R1177 VTAIL.n795 VTAIL.n758 0.388379
R1178 VTAIL.n838 VTAIL.n736 0.388379
R1179 VTAIL.n58 VTAIL.n57 0.388379
R1180 VTAIL.n61 VTAIL.n24 0.388379
R1181 VTAIL.n104 VTAIL.n2 0.388379
R1182 VTAIL.n162 VTAIL.n161 0.388379
R1183 VTAIL.n165 VTAIL.n128 0.388379
R1184 VTAIL.n208 VTAIL.n106 0.388379
R1185 VTAIL.n268 VTAIL.n267 0.388379
R1186 VTAIL.n271 VTAIL.n234 0.388379
R1187 VTAIL.n314 VTAIL.n212 0.388379
R1188 VTAIL.n734 VTAIL.n632 0.388379
R1189 VTAIL.n691 VTAIL.n654 0.388379
R1190 VTAIL.n688 VTAIL.n656 0.388379
R1191 VTAIL.n628 VTAIL.n526 0.388379
R1192 VTAIL.n585 VTAIL.n548 0.388379
R1193 VTAIL.n582 VTAIL.n550 0.388379
R1194 VTAIL.n524 VTAIL.n422 0.388379
R1195 VTAIL.n481 VTAIL.n444 0.388379
R1196 VTAIL.n478 VTAIL.n446 0.388379
R1197 VTAIL.n418 VTAIL.n316 0.388379
R1198 VTAIL.n375 VTAIL.n338 0.388379
R1199 VTAIL.n372 VTAIL.n340 0.388379
R1200 VTAIL.n775 VTAIL.n767 0.155672
R1201 VTAIL.n776 VTAIL.n775 0.155672
R1202 VTAIL.n776 VTAIL.n763 0.155672
R1203 VTAIL.n783 VTAIL.n763 0.155672
R1204 VTAIL.n784 VTAIL.n783 0.155672
R1205 VTAIL.n784 VTAIL.n759 0.155672
R1206 VTAIL.n793 VTAIL.n759 0.155672
R1207 VTAIL.n794 VTAIL.n793 0.155672
R1208 VTAIL.n794 VTAIL.n755 0.155672
R1209 VTAIL.n801 VTAIL.n755 0.155672
R1210 VTAIL.n802 VTAIL.n801 0.155672
R1211 VTAIL.n802 VTAIL.n751 0.155672
R1212 VTAIL.n809 VTAIL.n751 0.155672
R1213 VTAIL.n810 VTAIL.n809 0.155672
R1214 VTAIL.n810 VTAIL.n747 0.155672
R1215 VTAIL.n817 VTAIL.n747 0.155672
R1216 VTAIL.n818 VTAIL.n817 0.155672
R1217 VTAIL.n818 VTAIL.n743 0.155672
R1218 VTAIL.n825 VTAIL.n743 0.155672
R1219 VTAIL.n826 VTAIL.n825 0.155672
R1220 VTAIL.n826 VTAIL.n739 0.155672
R1221 VTAIL.n833 VTAIL.n739 0.155672
R1222 VTAIL.n834 VTAIL.n833 0.155672
R1223 VTAIL.n41 VTAIL.n33 0.155672
R1224 VTAIL.n42 VTAIL.n41 0.155672
R1225 VTAIL.n42 VTAIL.n29 0.155672
R1226 VTAIL.n49 VTAIL.n29 0.155672
R1227 VTAIL.n50 VTAIL.n49 0.155672
R1228 VTAIL.n50 VTAIL.n25 0.155672
R1229 VTAIL.n59 VTAIL.n25 0.155672
R1230 VTAIL.n60 VTAIL.n59 0.155672
R1231 VTAIL.n60 VTAIL.n21 0.155672
R1232 VTAIL.n67 VTAIL.n21 0.155672
R1233 VTAIL.n68 VTAIL.n67 0.155672
R1234 VTAIL.n68 VTAIL.n17 0.155672
R1235 VTAIL.n75 VTAIL.n17 0.155672
R1236 VTAIL.n76 VTAIL.n75 0.155672
R1237 VTAIL.n76 VTAIL.n13 0.155672
R1238 VTAIL.n83 VTAIL.n13 0.155672
R1239 VTAIL.n84 VTAIL.n83 0.155672
R1240 VTAIL.n84 VTAIL.n9 0.155672
R1241 VTAIL.n91 VTAIL.n9 0.155672
R1242 VTAIL.n92 VTAIL.n91 0.155672
R1243 VTAIL.n92 VTAIL.n5 0.155672
R1244 VTAIL.n99 VTAIL.n5 0.155672
R1245 VTAIL.n100 VTAIL.n99 0.155672
R1246 VTAIL.n145 VTAIL.n137 0.155672
R1247 VTAIL.n146 VTAIL.n145 0.155672
R1248 VTAIL.n146 VTAIL.n133 0.155672
R1249 VTAIL.n153 VTAIL.n133 0.155672
R1250 VTAIL.n154 VTAIL.n153 0.155672
R1251 VTAIL.n154 VTAIL.n129 0.155672
R1252 VTAIL.n163 VTAIL.n129 0.155672
R1253 VTAIL.n164 VTAIL.n163 0.155672
R1254 VTAIL.n164 VTAIL.n125 0.155672
R1255 VTAIL.n171 VTAIL.n125 0.155672
R1256 VTAIL.n172 VTAIL.n171 0.155672
R1257 VTAIL.n172 VTAIL.n121 0.155672
R1258 VTAIL.n179 VTAIL.n121 0.155672
R1259 VTAIL.n180 VTAIL.n179 0.155672
R1260 VTAIL.n180 VTAIL.n117 0.155672
R1261 VTAIL.n187 VTAIL.n117 0.155672
R1262 VTAIL.n188 VTAIL.n187 0.155672
R1263 VTAIL.n188 VTAIL.n113 0.155672
R1264 VTAIL.n195 VTAIL.n113 0.155672
R1265 VTAIL.n196 VTAIL.n195 0.155672
R1266 VTAIL.n196 VTAIL.n109 0.155672
R1267 VTAIL.n203 VTAIL.n109 0.155672
R1268 VTAIL.n204 VTAIL.n203 0.155672
R1269 VTAIL.n251 VTAIL.n243 0.155672
R1270 VTAIL.n252 VTAIL.n251 0.155672
R1271 VTAIL.n252 VTAIL.n239 0.155672
R1272 VTAIL.n259 VTAIL.n239 0.155672
R1273 VTAIL.n260 VTAIL.n259 0.155672
R1274 VTAIL.n260 VTAIL.n235 0.155672
R1275 VTAIL.n269 VTAIL.n235 0.155672
R1276 VTAIL.n270 VTAIL.n269 0.155672
R1277 VTAIL.n270 VTAIL.n231 0.155672
R1278 VTAIL.n277 VTAIL.n231 0.155672
R1279 VTAIL.n278 VTAIL.n277 0.155672
R1280 VTAIL.n278 VTAIL.n227 0.155672
R1281 VTAIL.n285 VTAIL.n227 0.155672
R1282 VTAIL.n286 VTAIL.n285 0.155672
R1283 VTAIL.n286 VTAIL.n223 0.155672
R1284 VTAIL.n293 VTAIL.n223 0.155672
R1285 VTAIL.n294 VTAIL.n293 0.155672
R1286 VTAIL.n294 VTAIL.n219 0.155672
R1287 VTAIL.n301 VTAIL.n219 0.155672
R1288 VTAIL.n302 VTAIL.n301 0.155672
R1289 VTAIL.n302 VTAIL.n215 0.155672
R1290 VTAIL.n309 VTAIL.n215 0.155672
R1291 VTAIL.n310 VTAIL.n309 0.155672
R1292 VTAIL.n730 VTAIL.n729 0.155672
R1293 VTAIL.n729 VTAIL.n635 0.155672
R1294 VTAIL.n722 VTAIL.n635 0.155672
R1295 VTAIL.n722 VTAIL.n721 0.155672
R1296 VTAIL.n721 VTAIL.n639 0.155672
R1297 VTAIL.n714 VTAIL.n639 0.155672
R1298 VTAIL.n714 VTAIL.n713 0.155672
R1299 VTAIL.n713 VTAIL.n643 0.155672
R1300 VTAIL.n706 VTAIL.n643 0.155672
R1301 VTAIL.n706 VTAIL.n705 0.155672
R1302 VTAIL.n705 VTAIL.n647 0.155672
R1303 VTAIL.n698 VTAIL.n647 0.155672
R1304 VTAIL.n698 VTAIL.n697 0.155672
R1305 VTAIL.n697 VTAIL.n651 0.155672
R1306 VTAIL.n690 VTAIL.n651 0.155672
R1307 VTAIL.n690 VTAIL.n689 0.155672
R1308 VTAIL.n689 VTAIL.n655 0.155672
R1309 VTAIL.n682 VTAIL.n655 0.155672
R1310 VTAIL.n682 VTAIL.n681 0.155672
R1311 VTAIL.n681 VTAIL.n661 0.155672
R1312 VTAIL.n674 VTAIL.n661 0.155672
R1313 VTAIL.n674 VTAIL.n673 0.155672
R1314 VTAIL.n673 VTAIL.n665 0.155672
R1315 VTAIL.n624 VTAIL.n623 0.155672
R1316 VTAIL.n623 VTAIL.n529 0.155672
R1317 VTAIL.n616 VTAIL.n529 0.155672
R1318 VTAIL.n616 VTAIL.n615 0.155672
R1319 VTAIL.n615 VTAIL.n533 0.155672
R1320 VTAIL.n608 VTAIL.n533 0.155672
R1321 VTAIL.n608 VTAIL.n607 0.155672
R1322 VTAIL.n607 VTAIL.n537 0.155672
R1323 VTAIL.n600 VTAIL.n537 0.155672
R1324 VTAIL.n600 VTAIL.n599 0.155672
R1325 VTAIL.n599 VTAIL.n541 0.155672
R1326 VTAIL.n592 VTAIL.n541 0.155672
R1327 VTAIL.n592 VTAIL.n591 0.155672
R1328 VTAIL.n591 VTAIL.n545 0.155672
R1329 VTAIL.n584 VTAIL.n545 0.155672
R1330 VTAIL.n584 VTAIL.n583 0.155672
R1331 VTAIL.n583 VTAIL.n549 0.155672
R1332 VTAIL.n576 VTAIL.n549 0.155672
R1333 VTAIL.n576 VTAIL.n575 0.155672
R1334 VTAIL.n575 VTAIL.n555 0.155672
R1335 VTAIL.n568 VTAIL.n555 0.155672
R1336 VTAIL.n568 VTAIL.n567 0.155672
R1337 VTAIL.n567 VTAIL.n559 0.155672
R1338 VTAIL.n520 VTAIL.n519 0.155672
R1339 VTAIL.n519 VTAIL.n425 0.155672
R1340 VTAIL.n512 VTAIL.n425 0.155672
R1341 VTAIL.n512 VTAIL.n511 0.155672
R1342 VTAIL.n511 VTAIL.n429 0.155672
R1343 VTAIL.n504 VTAIL.n429 0.155672
R1344 VTAIL.n504 VTAIL.n503 0.155672
R1345 VTAIL.n503 VTAIL.n433 0.155672
R1346 VTAIL.n496 VTAIL.n433 0.155672
R1347 VTAIL.n496 VTAIL.n495 0.155672
R1348 VTAIL.n495 VTAIL.n437 0.155672
R1349 VTAIL.n488 VTAIL.n437 0.155672
R1350 VTAIL.n488 VTAIL.n487 0.155672
R1351 VTAIL.n487 VTAIL.n441 0.155672
R1352 VTAIL.n480 VTAIL.n441 0.155672
R1353 VTAIL.n480 VTAIL.n479 0.155672
R1354 VTAIL.n479 VTAIL.n445 0.155672
R1355 VTAIL.n472 VTAIL.n445 0.155672
R1356 VTAIL.n472 VTAIL.n471 0.155672
R1357 VTAIL.n471 VTAIL.n451 0.155672
R1358 VTAIL.n464 VTAIL.n451 0.155672
R1359 VTAIL.n464 VTAIL.n463 0.155672
R1360 VTAIL.n463 VTAIL.n455 0.155672
R1361 VTAIL.n414 VTAIL.n413 0.155672
R1362 VTAIL.n413 VTAIL.n319 0.155672
R1363 VTAIL.n406 VTAIL.n319 0.155672
R1364 VTAIL.n406 VTAIL.n405 0.155672
R1365 VTAIL.n405 VTAIL.n323 0.155672
R1366 VTAIL.n398 VTAIL.n323 0.155672
R1367 VTAIL.n398 VTAIL.n397 0.155672
R1368 VTAIL.n397 VTAIL.n327 0.155672
R1369 VTAIL.n390 VTAIL.n327 0.155672
R1370 VTAIL.n390 VTAIL.n389 0.155672
R1371 VTAIL.n389 VTAIL.n331 0.155672
R1372 VTAIL.n382 VTAIL.n331 0.155672
R1373 VTAIL.n382 VTAIL.n381 0.155672
R1374 VTAIL.n381 VTAIL.n335 0.155672
R1375 VTAIL.n374 VTAIL.n335 0.155672
R1376 VTAIL.n374 VTAIL.n373 0.155672
R1377 VTAIL.n373 VTAIL.n339 0.155672
R1378 VTAIL.n366 VTAIL.n339 0.155672
R1379 VTAIL.n366 VTAIL.n365 0.155672
R1380 VTAIL.n365 VTAIL.n345 0.155672
R1381 VTAIL.n358 VTAIL.n345 0.155672
R1382 VTAIL.n358 VTAIL.n357 0.155672
R1383 VTAIL.n357 VTAIL.n349 0.155672
R1384 VTAIL VTAIL.n1 0.0586897
R1385 B.n1142 B.n1141 585
R1386 B.n438 B.n174 585
R1387 B.n437 B.n436 585
R1388 B.n435 B.n434 585
R1389 B.n433 B.n432 585
R1390 B.n431 B.n430 585
R1391 B.n429 B.n428 585
R1392 B.n427 B.n426 585
R1393 B.n425 B.n424 585
R1394 B.n423 B.n422 585
R1395 B.n421 B.n420 585
R1396 B.n419 B.n418 585
R1397 B.n417 B.n416 585
R1398 B.n415 B.n414 585
R1399 B.n413 B.n412 585
R1400 B.n411 B.n410 585
R1401 B.n409 B.n408 585
R1402 B.n407 B.n406 585
R1403 B.n405 B.n404 585
R1404 B.n403 B.n402 585
R1405 B.n401 B.n400 585
R1406 B.n399 B.n398 585
R1407 B.n397 B.n396 585
R1408 B.n395 B.n394 585
R1409 B.n393 B.n392 585
R1410 B.n391 B.n390 585
R1411 B.n389 B.n388 585
R1412 B.n387 B.n386 585
R1413 B.n385 B.n384 585
R1414 B.n383 B.n382 585
R1415 B.n381 B.n380 585
R1416 B.n379 B.n378 585
R1417 B.n377 B.n376 585
R1418 B.n375 B.n374 585
R1419 B.n373 B.n372 585
R1420 B.n371 B.n370 585
R1421 B.n369 B.n368 585
R1422 B.n367 B.n366 585
R1423 B.n365 B.n364 585
R1424 B.n363 B.n362 585
R1425 B.n361 B.n360 585
R1426 B.n359 B.n358 585
R1427 B.n357 B.n356 585
R1428 B.n355 B.n354 585
R1429 B.n353 B.n352 585
R1430 B.n351 B.n350 585
R1431 B.n349 B.n348 585
R1432 B.n347 B.n346 585
R1433 B.n345 B.n344 585
R1434 B.n343 B.n342 585
R1435 B.n341 B.n340 585
R1436 B.n339 B.n338 585
R1437 B.n337 B.n336 585
R1438 B.n335 B.n334 585
R1439 B.n333 B.n332 585
R1440 B.n331 B.n330 585
R1441 B.n329 B.n328 585
R1442 B.n327 B.n326 585
R1443 B.n325 B.n324 585
R1444 B.n323 B.n322 585
R1445 B.n321 B.n320 585
R1446 B.n318 B.n317 585
R1447 B.n316 B.n315 585
R1448 B.n314 B.n313 585
R1449 B.n312 B.n311 585
R1450 B.n310 B.n309 585
R1451 B.n308 B.n307 585
R1452 B.n306 B.n305 585
R1453 B.n304 B.n303 585
R1454 B.n302 B.n301 585
R1455 B.n300 B.n299 585
R1456 B.n297 B.n296 585
R1457 B.n295 B.n294 585
R1458 B.n293 B.n292 585
R1459 B.n291 B.n290 585
R1460 B.n289 B.n288 585
R1461 B.n287 B.n286 585
R1462 B.n285 B.n284 585
R1463 B.n283 B.n282 585
R1464 B.n281 B.n280 585
R1465 B.n279 B.n278 585
R1466 B.n277 B.n276 585
R1467 B.n275 B.n274 585
R1468 B.n273 B.n272 585
R1469 B.n271 B.n270 585
R1470 B.n269 B.n268 585
R1471 B.n267 B.n266 585
R1472 B.n265 B.n264 585
R1473 B.n263 B.n262 585
R1474 B.n261 B.n260 585
R1475 B.n259 B.n258 585
R1476 B.n257 B.n256 585
R1477 B.n255 B.n254 585
R1478 B.n253 B.n252 585
R1479 B.n251 B.n250 585
R1480 B.n249 B.n248 585
R1481 B.n247 B.n246 585
R1482 B.n245 B.n244 585
R1483 B.n243 B.n242 585
R1484 B.n241 B.n240 585
R1485 B.n239 B.n238 585
R1486 B.n237 B.n236 585
R1487 B.n235 B.n234 585
R1488 B.n233 B.n232 585
R1489 B.n231 B.n230 585
R1490 B.n229 B.n228 585
R1491 B.n227 B.n226 585
R1492 B.n225 B.n224 585
R1493 B.n223 B.n222 585
R1494 B.n221 B.n220 585
R1495 B.n219 B.n218 585
R1496 B.n217 B.n216 585
R1497 B.n215 B.n214 585
R1498 B.n213 B.n212 585
R1499 B.n211 B.n210 585
R1500 B.n209 B.n208 585
R1501 B.n207 B.n206 585
R1502 B.n205 B.n204 585
R1503 B.n203 B.n202 585
R1504 B.n201 B.n200 585
R1505 B.n199 B.n198 585
R1506 B.n197 B.n196 585
R1507 B.n195 B.n194 585
R1508 B.n193 B.n192 585
R1509 B.n191 B.n190 585
R1510 B.n189 B.n188 585
R1511 B.n187 B.n186 585
R1512 B.n185 B.n184 585
R1513 B.n183 B.n182 585
R1514 B.n181 B.n180 585
R1515 B.n109 B.n108 585
R1516 B.n1147 B.n1146 585
R1517 B.n1140 B.n175 585
R1518 B.n175 B.n106 585
R1519 B.n1139 B.n105 585
R1520 B.n1151 B.n105 585
R1521 B.n1138 B.n104 585
R1522 B.n1152 B.n104 585
R1523 B.n1137 B.n103 585
R1524 B.n1153 B.n103 585
R1525 B.n1136 B.n1135 585
R1526 B.n1135 B.n99 585
R1527 B.n1134 B.n98 585
R1528 B.n1159 B.n98 585
R1529 B.n1133 B.n97 585
R1530 B.n1160 B.n97 585
R1531 B.n1132 B.n96 585
R1532 B.n1161 B.n96 585
R1533 B.n1131 B.n1130 585
R1534 B.n1130 B.n95 585
R1535 B.n1129 B.n91 585
R1536 B.n1167 B.n91 585
R1537 B.n1128 B.n90 585
R1538 B.n1168 B.n90 585
R1539 B.n1127 B.n89 585
R1540 B.n1169 B.n89 585
R1541 B.n1126 B.n1125 585
R1542 B.n1125 B.n85 585
R1543 B.n1124 B.n84 585
R1544 B.n1175 B.n84 585
R1545 B.n1123 B.n83 585
R1546 B.n1176 B.n83 585
R1547 B.n1122 B.n82 585
R1548 B.n1177 B.n82 585
R1549 B.n1121 B.n1120 585
R1550 B.n1120 B.n78 585
R1551 B.n1119 B.n77 585
R1552 B.n1183 B.n77 585
R1553 B.n1118 B.n76 585
R1554 B.n1184 B.n76 585
R1555 B.n1117 B.n75 585
R1556 B.n1185 B.n75 585
R1557 B.n1116 B.n1115 585
R1558 B.n1115 B.n71 585
R1559 B.n1114 B.n70 585
R1560 B.n1191 B.n70 585
R1561 B.n1113 B.n69 585
R1562 B.n1192 B.n69 585
R1563 B.n1112 B.n68 585
R1564 B.n1193 B.n68 585
R1565 B.n1111 B.n1110 585
R1566 B.n1110 B.n64 585
R1567 B.n1109 B.n63 585
R1568 B.n1199 B.n63 585
R1569 B.n1108 B.n62 585
R1570 B.n1200 B.n62 585
R1571 B.n1107 B.n61 585
R1572 B.n1201 B.n61 585
R1573 B.n1106 B.n1105 585
R1574 B.n1105 B.n57 585
R1575 B.n1104 B.n56 585
R1576 B.n1207 B.n56 585
R1577 B.n1103 B.n55 585
R1578 B.n1208 B.n55 585
R1579 B.n1102 B.n54 585
R1580 B.n1209 B.n54 585
R1581 B.n1101 B.n1100 585
R1582 B.n1100 B.n50 585
R1583 B.n1099 B.n49 585
R1584 B.n1215 B.n49 585
R1585 B.n1098 B.n48 585
R1586 B.n1216 B.n48 585
R1587 B.n1097 B.n47 585
R1588 B.n1217 B.n47 585
R1589 B.n1096 B.n1095 585
R1590 B.n1095 B.n43 585
R1591 B.n1094 B.n42 585
R1592 B.n1223 B.n42 585
R1593 B.n1093 B.n41 585
R1594 B.n1224 B.n41 585
R1595 B.n1092 B.n40 585
R1596 B.n1225 B.n40 585
R1597 B.n1091 B.n1090 585
R1598 B.n1090 B.n36 585
R1599 B.n1089 B.n35 585
R1600 B.n1231 B.n35 585
R1601 B.n1088 B.n34 585
R1602 B.n1232 B.n34 585
R1603 B.n1087 B.n33 585
R1604 B.n1233 B.n33 585
R1605 B.n1086 B.n1085 585
R1606 B.n1085 B.n29 585
R1607 B.n1084 B.n28 585
R1608 B.n1239 B.n28 585
R1609 B.n1083 B.n27 585
R1610 B.n1240 B.n27 585
R1611 B.n1082 B.n26 585
R1612 B.n1241 B.n26 585
R1613 B.n1081 B.n1080 585
R1614 B.n1080 B.n22 585
R1615 B.n1079 B.n21 585
R1616 B.n1247 B.n21 585
R1617 B.n1078 B.n20 585
R1618 B.n1248 B.n20 585
R1619 B.n1077 B.n19 585
R1620 B.n1249 B.n19 585
R1621 B.n1076 B.n1075 585
R1622 B.n1075 B.n18 585
R1623 B.n1074 B.n14 585
R1624 B.n1255 B.n14 585
R1625 B.n1073 B.n13 585
R1626 B.n1256 B.n13 585
R1627 B.n1072 B.n12 585
R1628 B.n1257 B.n12 585
R1629 B.n1071 B.n1070 585
R1630 B.n1070 B.n8 585
R1631 B.n1069 B.n7 585
R1632 B.n1263 B.n7 585
R1633 B.n1068 B.n6 585
R1634 B.n1264 B.n6 585
R1635 B.n1067 B.n5 585
R1636 B.n1265 B.n5 585
R1637 B.n1066 B.n1065 585
R1638 B.n1065 B.n4 585
R1639 B.n1064 B.n439 585
R1640 B.n1064 B.n1063 585
R1641 B.n1054 B.n440 585
R1642 B.n441 B.n440 585
R1643 B.n1056 B.n1055 585
R1644 B.n1057 B.n1056 585
R1645 B.n1053 B.n446 585
R1646 B.n446 B.n445 585
R1647 B.n1052 B.n1051 585
R1648 B.n1051 B.n1050 585
R1649 B.n448 B.n447 585
R1650 B.n1043 B.n448 585
R1651 B.n1042 B.n1041 585
R1652 B.n1044 B.n1042 585
R1653 B.n1040 B.n453 585
R1654 B.n453 B.n452 585
R1655 B.n1039 B.n1038 585
R1656 B.n1038 B.n1037 585
R1657 B.n455 B.n454 585
R1658 B.n456 B.n455 585
R1659 B.n1030 B.n1029 585
R1660 B.n1031 B.n1030 585
R1661 B.n1028 B.n461 585
R1662 B.n461 B.n460 585
R1663 B.n1027 B.n1026 585
R1664 B.n1026 B.n1025 585
R1665 B.n463 B.n462 585
R1666 B.n464 B.n463 585
R1667 B.n1018 B.n1017 585
R1668 B.n1019 B.n1018 585
R1669 B.n1016 B.n468 585
R1670 B.n472 B.n468 585
R1671 B.n1015 B.n1014 585
R1672 B.n1014 B.n1013 585
R1673 B.n470 B.n469 585
R1674 B.n471 B.n470 585
R1675 B.n1006 B.n1005 585
R1676 B.n1007 B.n1006 585
R1677 B.n1004 B.n477 585
R1678 B.n477 B.n476 585
R1679 B.n1003 B.n1002 585
R1680 B.n1002 B.n1001 585
R1681 B.n479 B.n478 585
R1682 B.n480 B.n479 585
R1683 B.n994 B.n993 585
R1684 B.n995 B.n994 585
R1685 B.n992 B.n485 585
R1686 B.n485 B.n484 585
R1687 B.n991 B.n990 585
R1688 B.n990 B.n989 585
R1689 B.n487 B.n486 585
R1690 B.n488 B.n487 585
R1691 B.n982 B.n981 585
R1692 B.n983 B.n982 585
R1693 B.n980 B.n493 585
R1694 B.n493 B.n492 585
R1695 B.n979 B.n978 585
R1696 B.n978 B.n977 585
R1697 B.n495 B.n494 585
R1698 B.n496 B.n495 585
R1699 B.n970 B.n969 585
R1700 B.n971 B.n970 585
R1701 B.n968 B.n501 585
R1702 B.n501 B.n500 585
R1703 B.n967 B.n966 585
R1704 B.n966 B.n965 585
R1705 B.n503 B.n502 585
R1706 B.n504 B.n503 585
R1707 B.n958 B.n957 585
R1708 B.n959 B.n958 585
R1709 B.n956 B.n509 585
R1710 B.n509 B.n508 585
R1711 B.n955 B.n954 585
R1712 B.n954 B.n953 585
R1713 B.n511 B.n510 585
R1714 B.n512 B.n511 585
R1715 B.n946 B.n945 585
R1716 B.n947 B.n946 585
R1717 B.n944 B.n517 585
R1718 B.n517 B.n516 585
R1719 B.n943 B.n942 585
R1720 B.n942 B.n941 585
R1721 B.n519 B.n518 585
R1722 B.n520 B.n519 585
R1723 B.n934 B.n933 585
R1724 B.n935 B.n934 585
R1725 B.n932 B.n525 585
R1726 B.n525 B.n524 585
R1727 B.n931 B.n930 585
R1728 B.n930 B.n929 585
R1729 B.n527 B.n526 585
R1730 B.n528 B.n527 585
R1731 B.n922 B.n921 585
R1732 B.n923 B.n922 585
R1733 B.n920 B.n533 585
R1734 B.n533 B.n532 585
R1735 B.n919 B.n918 585
R1736 B.n918 B.n917 585
R1737 B.n535 B.n534 585
R1738 B.n910 B.n535 585
R1739 B.n909 B.n908 585
R1740 B.n911 B.n909 585
R1741 B.n907 B.n540 585
R1742 B.n540 B.n539 585
R1743 B.n906 B.n905 585
R1744 B.n905 B.n904 585
R1745 B.n542 B.n541 585
R1746 B.n543 B.n542 585
R1747 B.n897 B.n896 585
R1748 B.n898 B.n897 585
R1749 B.n895 B.n548 585
R1750 B.n548 B.n547 585
R1751 B.n894 B.n893 585
R1752 B.n893 B.n892 585
R1753 B.n550 B.n549 585
R1754 B.n551 B.n550 585
R1755 B.n888 B.n887 585
R1756 B.n554 B.n553 585
R1757 B.n884 B.n883 585
R1758 B.n885 B.n884 585
R1759 B.n882 B.n620 585
R1760 B.n881 B.n880 585
R1761 B.n879 B.n878 585
R1762 B.n877 B.n876 585
R1763 B.n875 B.n874 585
R1764 B.n873 B.n872 585
R1765 B.n871 B.n870 585
R1766 B.n869 B.n868 585
R1767 B.n867 B.n866 585
R1768 B.n865 B.n864 585
R1769 B.n863 B.n862 585
R1770 B.n861 B.n860 585
R1771 B.n859 B.n858 585
R1772 B.n857 B.n856 585
R1773 B.n855 B.n854 585
R1774 B.n853 B.n852 585
R1775 B.n851 B.n850 585
R1776 B.n849 B.n848 585
R1777 B.n847 B.n846 585
R1778 B.n845 B.n844 585
R1779 B.n843 B.n842 585
R1780 B.n841 B.n840 585
R1781 B.n839 B.n838 585
R1782 B.n837 B.n836 585
R1783 B.n835 B.n834 585
R1784 B.n833 B.n832 585
R1785 B.n831 B.n830 585
R1786 B.n829 B.n828 585
R1787 B.n827 B.n826 585
R1788 B.n825 B.n824 585
R1789 B.n823 B.n822 585
R1790 B.n821 B.n820 585
R1791 B.n819 B.n818 585
R1792 B.n817 B.n816 585
R1793 B.n815 B.n814 585
R1794 B.n813 B.n812 585
R1795 B.n811 B.n810 585
R1796 B.n809 B.n808 585
R1797 B.n807 B.n806 585
R1798 B.n805 B.n804 585
R1799 B.n803 B.n802 585
R1800 B.n801 B.n800 585
R1801 B.n799 B.n798 585
R1802 B.n797 B.n796 585
R1803 B.n795 B.n794 585
R1804 B.n793 B.n792 585
R1805 B.n791 B.n790 585
R1806 B.n789 B.n788 585
R1807 B.n787 B.n786 585
R1808 B.n785 B.n784 585
R1809 B.n783 B.n782 585
R1810 B.n781 B.n780 585
R1811 B.n779 B.n778 585
R1812 B.n777 B.n776 585
R1813 B.n775 B.n774 585
R1814 B.n773 B.n772 585
R1815 B.n771 B.n770 585
R1816 B.n769 B.n768 585
R1817 B.n767 B.n766 585
R1818 B.n765 B.n764 585
R1819 B.n763 B.n762 585
R1820 B.n761 B.n760 585
R1821 B.n759 B.n758 585
R1822 B.n757 B.n756 585
R1823 B.n755 B.n754 585
R1824 B.n753 B.n752 585
R1825 B.n751 B.n750 585
R1826 B.n749 B.n748 585
R1827 B.n747 B.n746 585
R1828 B.n745 B.n744 585
R1829 B.n743 B.n742 585
R1830 B.n741 B.n740 585
R1831 B.n739 B.n738 585
R1832 B.n737 B.n736 585
R1833 B.n735 B.n734 585
R1834 B.n733 B.n732 585
R1835 B.n731 B.n730 585
R1836 B.n729 B.n728 585
R1837 B.n727 B.n726 585
R1838 B.n725 B.n724 585
R1839 B.n723 B.n722 585
R1840 B.n721 B.n720 585
R1841 B.n719 B.n718 585
R1842 B.n717 B.n716 585
R1843 B.n715 B.n714 585
R1844 B.n713 B.n712 585
R1845 B.n711 B.n710 585
R1846 B.n709 B.n708 585
R1847 B.n707 B.n706 585
R1848 B.n705 B.n704 585
R1849 B.n703 B.n702 585
R1850 B.n701 B.n700 585
R1851 B.n699 B.n698 585
R1852 B.n697 B.n696 585
R1853 B.n695 B.n694 585
R1854 B.n693 B.n692 585
R1855 B.n691 B.n690 585
R1856 B.n689 B.n688 585
R1857 B.n687 B.n686 585
R1858 B.n685 B.n684 585
R1859 B.n683 B.n682 585
R1860 B.n681 B.n680 585
R1861 B.n679 B.n678 585
R1862 B.n677 B.n676 585
R1863 B.n675 B.n674 585
R1864 B.n673 B.n672 585
R1865 B.n671 B.n670 585
R1866 B.n669 B.n668 585
R1867 B.n667 B.n666 585
R1868 B.n665 B.n664 585
R1869 B.n663 B.n662 585
R1870 B.n661 B.n660 585
R1871 B.n659 B.n658 585
R1872 B.n657 B.n656 585
R1873 B.n655 B.n654 585
R1874 B.n653 B.n652 585
R1875 B.n651 B.n650 585
R1876 B.n649 B.n648 585
R1877 B.n647 B.n646 585
R1878 B.n645 B.n644 585
R1879 B.n643 B.n642 585
R1880 B.n641 B.n640 585
R1881 B.n639 B.n638 585
R1882 B.n637 B.n636 585
R1883 B.n635 B.n634 585
R1884 B.n633 B.n632 585
R1885 B.n631 B.n630 585
R1886 B.n629 B.n628 585
R1887 B.n627 B.n619 585
R1888 B.n885 B.n619 585
R1889 B.n889 B.n552 585
R1890 B.n552 B.n551 585
R1891 B.n891 B.n890 585
R1892 B.n892 B.n891 585
R1893 B.n546 B.n545 585
R1894 B.n547 B.n546 585
R1895 B.n900 B.n899 585
R1896 B.n899 B.n898 585
R1897 B.n901 B.n544 585
R1898 B.n544 B.n543 585
R1899 B.n903 B.n902 585
R1900 B.n904 B.n903 585
R1901 B.n538 B.n537 585
R1902 B.n539 B.n538 585
R1903 B.n913 B.n912 585
R1904 B.n912 B.n911 585
R1905 B.n914 B.n536 585
R1906 B.n910 B.n536 585
R1907 B.n916 B.n915 585
R1908 B.n917 B.n916 585
R1909 B.n531 B.n530 585
R1910 B.n532 B.n531 585
R1911 B.n925 B.n924 585
R1912 B.n924 B.n923 585
R1913 B.n926 B.n529 585
R1914 B.n529 B.n528 585
R1915 B.n928 B.n927 585
R1916 B.n929 B.n928 585
R1917 B.n523 B.n522 585
R1918 B.n524 B.n523 585
R1919 B.n937 B.n936 585
R1920 B.n936 B.n935 585
R1921 B.n938 B.n521 585
R1922 B.n521 B.n520 585
R1923 B.n940 B.n939 585
R1924 B.n941 B.n940 585
R1925 B.n515 B.n514 585
R1926 B.n516 B.n515 585
R1927 B.n949 B.n948 585
R1928 B.n948 B.n947 585
R1929 B.n950 B.n513 585
R1930 B.n513 B.n512 585
R1931 B.n952 B.n951 585
R1932 B.n953 B.n952 585
R1933 B.n507 B.n506 585
R1934 B.n508 B.n507 585
R1935 B.n961 B.n960 585
R1936 B.n960 B.n959 585
R1937 B.n962 B.n505 585
R1938 B.n505 B.n504 585
R1939 B.n964 B.n963 585
R1940 B.n965 B.n964 585
R1941 B.n499 B.n498 585
R1942 B.n500 B.n499 585
R1943 B.n973 B.n972 585
R1944 B.n972 B.n971 585
R1945 B.n974 B.n497 585
R1946 B.n497 B.n496 585
R1947 B.n976 B.n975 585
R1948 B.n977 B.n976 585
R1949 B.n491 B.n490 585
R1950 B.n492 B.n491 585
R1951 B.n985 B.n984 585
R1952 B.n984 B.n983 585
R1953 B.n986 B.n489 585
R1954 B.n489 B.n488 585
R1955 B.n988 B.n987 585
R1956 B.n989 B.n988 585
R1957 B.n483 B.n482 585
R1958 B.n484 B.n483 585
R1959 B.n997 B.n996 585
R1960 B.n996 B.n995 585
R1961 B.n998 B.n481 585
R1962 B.n481 B.n480 585
R1963 B.n1000 B.n999 585
R1964 B.n1001 B.n1000 585
R1965 B.n475 B.n474 585
R1966 B.n476 B.n475 585
R1967 B.n1009 B.n1008 585
R1968 B.n1008 B.n1007 585
R1969 B.n1010 B.n473 585
R1970 B.n473 B.n471 585
R1971 B.n1012 B.n1011 585
R1972 B.n1013 B.n1012 585
R1973 B.n467 B.n466 585
R1974 B.n472 B.n467 585
R1975 B.n1021 B.n1020 585
R1976 B.n1020 B.n1019 585
R1977 B.n1022 B.n465 585
R1978 B.n465 B.n464 585
R1979 B.n1024 B.n1023 585
R1980 B.n1025 B.n1024 585
R1981 B.n459 B.n458 585
R1982 B.n460 B.n459 585
R1983 B.n1033 B.n1032 585
R1984 B.n1032 B.n1031 585
R1985 B.n1034 B.n457 585
R1986 B.n457 B.n456 585
R1987 B.n1036 B.n1035 585
R1988 B.n1037 B.n1036 585
R1989 B.n451 B.n450 585
R1990 B.n452 B.n451 585
R1991 B.n1046 B.n1045 585
R1992 B.n1045 B.n1044 585
R1993 B.n1047 B.n449 585
R1994 B.n1043 B.n449 585
R1995 B.n1049 B.n1048 585
R1996 B.n1050 B.n1049 585
R1997 B.n444 B.n443 585
R1998 B.n445 B.n444 585
R1999 B.n1059 B.n1058 585
R2000 B.n1058 B.n1057 585
R2001 B.n1060 B.n442 585
R2002 B.n442 B.n441 585
R2003 B.n1062 B.n1061 585
R2004 B.n1063 B.n1062 585
R2005 B.n2 B.n0 585
R2006 B.n4 B.n2 585
R2007 B.n3 B.n1 585
R2008 B.n1264 B.n3 585
R2009 B.n1262 B.n1261 585
R2010 B.n1263 B.n1262 585
R2011 B.n1260 B.n9 585
R2012 B.n9 B.n8 585
R2013 B.n1259 B.n1258 585
R2014 B.n1258 B.n1257 585
R2015 B.n11 B.n10 585
R2016 B.n1256 B.n11 585
R2017 B.n1254 B.n1253 585
R2018 B.n1255 B.n1254 585
R2019 B.n1252 B.n15 585
R2020 B.n18 B.n15 585
R2021 B.n1251 B.n1250 585
R2022 B.n1250 B.n1249 585
R2023 B.n17 B.n16 585
R2024 B.n1248 B.n17 585
R2025 B.n1246 B.n1245 585
R2026 B.n1247 B.n1246 585
R2027 B.n1244 B.n23 585
R2028 B.n23 B.n22 585
R2029 B.n1243 B.n1242 585
R2030 B.n1242 B.n1241 585
R2031 B.n25 B.n24 585
R2032 B.n1240 B.n25 585
R2033 B.n1238 B.n1237 585
R2034 B.n1239 B.n1238 585
R2035 B.n1236 B.n30 585
R2036 B.n30 B.n29 585
R2037 B.n1235 B.n1234 585
R2038 B.n1234 B.n1233 585
R2039 B.n32 B.n31 585
R2040 B.n1232 B.n32 585
R2041 B.n1230 B.n1229 585
R2042 B.n1231 B.n1230 585
R2043 B.n1228 B.n37 585
R2044 B.n37 B.n36 585
R2045 B.n1227 B.n1226 585
R2046 B.n1226 B.n1225 585
R2047 B.n39 B.n38 585
R2048 B.n1224 B.n39 585
R2049 B.n1222 B.n1221 585
R2050 B.n1223 B.n1222 585
R2051 B.n1220 B.n44 585
R2052 B.n44 B.n43 585
R2053 B.n1219 B.n1218 585
R2054 B.n1218 B.n1217 585
R2055 B.n46 B.n45 585
R2056 B.n1216 B.n46 585
R2057 B.n1214 B.n1213 585
R2058 B.n1215 B.n1214 585
R2059 B.n1212 B.n51 585
R2060 B.n51 B.n50 585
R2061 B.n1211 B.n1210 585
R2062 B.n1210 B.n1209 585
R2063 B.n53 B.n52 585
R2064 B.n1208 B.n53 585
R2065 B.n1206 B.n1205 585
R2066 B.n1207 B.n1206 585
R2067 B.n1204 B.n58 585
R2068 B.n58 B.n57 585
R2069 B.n1203 B.n1202 585
R2070 B.n1202 B.n1201 585
R2071 B.n60 B.n59 585
R2072 B.n1200 B.n60 585
R2073 B.n1198 B.n1197 585
R2074 B.n1199 B.n1198 585
R2075 B.n1196 B.n65 585
R2076 B.n65 B.n64 585
R2077 B.n1195 B.n1194 585
R2078 B.n1194 B.n1193 585
R2079 B.n67 B.n66 585
R2080 B.n1192 B.n67 585
R2081 B.n1190 B.n1189 585
R2082 B.n1191 B.n1190 585
R2083 B.n1188 B.n72 585
R2084 B.n72 B.n71 585
R2085 B.n1187 B.n1186 585
R2086 B.n1186 B.n1185 585
R2087 B.n74 B.n73 585
R2088 B.n1184 B.n74 585
R2089 B.n1182 B.n1181 585
R2090 B.n1183 B.n1182 585
R2091 B.n1180 B.n79 585
R2092 B.n79 B.n78 585
R2093 B.n1179 B.n1178 585
R2094 B.n1178 B.n1177 585
R2095 B.n81 B.n80 585
R2096 B.n1176 B.n81 585
R2097 B.n1174 B.n1173 585
R2098 B.n1175 B.n1174 585
R2099 B.n1172 B.n86 585
R2100 B.n86 B.n85 585
R2101 B.n1171 B.n1170 585
R2102 B.n1170 B.n1169 585
R2103 B.n88 B.n87 585
R2104 B.n1168 B.n88 585
R2105 B.n1166 B.n1165 585
R2106 B.n1167 B.n1166 585
R2107 B.n1164 B.n92 585
R2108 B.n95 B.n92 585
R2109 B.n1163 B.n1162 585
R2110 B.n1162 B.n1161 585
R2111 B.n94 B.n93 585
R2112 B.n1160 B.n94 585
R2113 B.n1158 B.n1157 585
R2114 B.n1159 B.n1158 585
R2115 B.n1156 B.n100 585
R2116 B.n100 B.n99 585
R2117 B.n1155 B.n1154 585
R2118 B.n1154 B.n1153 585
R2119 B.n102 B.n101 585
R2120 B.n1152 B.n102 585
R2121 B.n1150 B.n1149 585
R2122 B.n1151 B.n1150 585
R2123 B.n1148 B.n107 585
R2124 B.n107 B.n106 585
R2125 B.n1267 B.n1266 585
R2126 B.n1266 B.n1265 585
R2127 B.n887 B.n552 521.33
R2128 B.n1146 B.n107 521.33
R2129 B.n619 B.n550 521.33
R2130 B.n1142 B.n175 521.33
R2131 B.n624 B.t14 464.49
R2132 B.n176 B.t20 464.49
R2133 B.n621 B.t11 464.49
R2134 B.n178 B.t17 464.49
R2135 B.n625 B.t13 397.387
R2136 B.n177 B.t21 397.387
R2137 B.n622 B.t10 397.387
R2138 B.n179 B.t18 397.387
R2139 B.n624 B.t12 352.788
R2140 B.n621 B.t8 352.788
R2141 B.n178 B.t15 352.788
R2142 B.n176 B.t19 352.788
R2143 B.n1144 B.n1143 256.663
R2144 B.n1144 B.n173 256.663
R2145 B.n1144 B.n172 256.663
R2146 B.n1144 B.n171 256.663
R2147 B.n1144 B.n170 256.663
R2148 B.n1144 B.n169 256.663
R2149 B.n1144 B.n168 256.663
R2150 B.n1144 B.n167 256.663
R2151 B.n1144 B.n166 256.663
R2152 B.n1144 B.n165 256.663
R2153 B.n1144 B.n164 256.663
R2154 B.n1144 B.n163 256.663
R2155 B.n1144 B.n162 256.663
R2156 B.n1144 B.n161 256.663
R2157 B.n1144 B.n160 256.663
R2158 B.n1144 B.n159 256.663
R2159 B.n1144 B.n158 256.663
R2160 B.n1144 B.n157 256.663
R2161 B.n1144 B.n156 256.663
R2162 B.n1144 B.n155 256.663
R2163 B.n1144 B.n154 256.663
R2164 B.n1144 B.n153 256.663
R2165 B.n1144 B.n152 256.663
R2166 B.n1144 B.n151 256.663
R2167 B.n1144 B.n150 256.663
R2168 B.n1144 B.n149 256.663
R2169 B.n1144 B.n148 256.663
R2170 B.n1144 B.n147 256.663
R2171 B.n1144 B.n146 256.663
R2172 B.n1144 B.n145 256.663
R2173 B.n1144 B.n144 256.663
R2174 B.n1144 B.n143 256.663
R2175 B.n1144 B.n142 256.663
R2176 B.n1144 B.n141 256.663
R2177 B.n1144 B.n140 256.663
R2178 B.n1144 B.n139 256.663
R2179 B.n1144 B.n138 256.663
R2180 B.n1144 B.n137 256.663
R2181 B.n1144 B.n136 256.663
R2182 B.n1144 B.n135 256.663
R2183 B.n1144 B.n134 256.663
R2184 B.n1144 B.n133 256.663
R2185 B.n1144 B.n132 256.663
R2186 B.n1144 B.n131 256.663
R2187 B.n1144 B.n130 256.663
R2188 B.n1144 B.n129 256.663
R2189 B.n1144 B.n128 256.663
R2190 B.n1144 B.n127 256.663
R2191 B.n1144 B.n126 256.663
R2192 B.n1144 B.n125 256.663
R2193 B.n1144 B.n124 256.663
R2194 B.n1144 B.n123 256.663
R2195 B.n1144 B.n122 256.663
R2196 B.n1144 B.n121 256.663
R2197 B.n1144 B.n120 256.663
R2198 B.n1144 B.n119 256.663
R2199 B.n1144 B.n118 256.663
R2200 B.n1144 B.n117 256.663
R2201 B.n1144 B.n116 256.663
R2202 B.n1144 B.n115 256.663
R2203 B.n1144 B.n114 256.663
R2204 B.n1144 B.n113 256.663
R2205 B.n1144 B.n112 256.663
R2206 B.n1144 B.n111 256.663
R2207 B.n1144 B.n110 256.663
R2208 B.n1145 B.n1144 256.663
R2209 B.n886 B.n885 256.663
R2210 B.n885 B.n555 256.663
R2211 B.n885 B.n556 256.663
R2212 B.n885 B.n557 256.663
R2213 B.n885 B.n558 256.663
R2214 B.n885 B.n559 256.663
R2215 B.n885 B.n560 256.663
R2216 B.n885 B.n561 256.663
R2217 B.n885 B.n562 256.663
R2218 B.n885 B.n563 256.663
R2219 B.n885 B.n564 256.663
R2220 B.n885 B.n565 256.663
R2221 B.n885 B.n566 256.663
R2222 B.n885 B.n567 256.663
R2223 B.n885 B.n568 256.663
R2224 B.n885 B.n569 256.663
R2225 B.n885 B.n570 256.663
R2226 B.n885 B.n571 256.663
R2227 B.n885 B.n572 256.663
R2228 B.n885 B.n573 256.663
R2229 B.n885 B.n574 256.663
R2230 B.n885 B.n575 256.663
R2231 B.n885 B.n576 256.663
R2232 B.n885 B.n577 256.663
R2233 B.n885 B.n578 256.663
R2234 B.n885 B.n579 256.663
R2235 B.n885 B.n580 256.663
R2236 B.n885 B.n581 256.663
R2237 B.n885 B.n582 256.663
R2238 B.n885 B.n583 256.663
R2239 B.n885 B.n584 256.663
R2240 B.n885 B.n585 256.663
R2241 B.n885 B.n586 256.663
R2242 B.n885 B.n587 256.663
R2243 B.n885 B.n588 256.663
R2244 B.n885 B.n589 256.663
R2245 B.n885 B.n590 256.663
R2246 B.n885 B.n591 256.663
R2247 B.n885 B.n592 256.663
R2248 B.n885 B.n593 256.663
R2249 B.n885 B.n594 256.663
R2250 B.n885 B.n595 256.663
R2251 B.n885 B.n596 256.663
R2252 B.n885 B.n597 256.663
R2253 B.n885 B.n598 256.663
R2254 B.n885 B.n599 256.663
R2255 B.n885 B.n600 256.663
R2256 B.n885 B.n601 256.663
R2257 B.n885 B.n602 256.663
R2258 B.n885 B.n603 256.663
R2259 B.n885 B.n604 256.663
R2260 B.n885 B.n605 256.663
R2261 B.n885 B.n606 256.663
R2262 B.n885 B.n607 256.663
R2263 B.n885 B.n608 256.663
R2264 B.n885 B.n609 256.663
R2265 B.n885 B.n610 256.663
R2266 B.n885 B.n611 256.663
R2267 B.n885 B.n612 256.663
R2268 B.n885 B.n613 256.663
R2269 B.n885 B.n614 256.663
R2270 B.n885 B.n615 256.663
R2271 B.n885 B.n616 256.663
R2272 B.n885 B.n617 256.663
R2273 B.n885 B.n618 256.663
R2274 B.n891 B.n552 163.367
R2275 B.n891 B.n546 163.367
R2276 B.n899 B.n546 163.367
R2277 B.n899 B.n544 163.367
R2278 B.n903 B.n544 163.367
R2279 B.n903 B.n538 163.367
R2280 B.n912 B.n538 163.367
R2281 B.n912 B.n536 163.367
R2282 B.n916 B.n536 163.367
R2283 B.n916 B.n531 163.367
R2284 B.n924 B.n531 163.367
R2285 B.n924 B.n529 163.367
R2286 B.n928 B.n529 163.367
R2287 B.n928 B.n523 163.367
R2288 B.n936 B.n523 163.367
R2289 B.n936 B.n521 163.367
R2290 B.n940 B.n521 163.367
R2291 B.n940 B.n515 163.367
R2292 B.n948 B.n515 163.367
R2293 B.n948 B.n513 163.367
R2294 B.n952 B.n513 163.367
R2295 B.n952 B.n507 163.367
R2296 B.n960 B.n507 163.367
R2297 B.n960 B.n505 163.367
R2298 B.n964 B.n505 163.367
R2299 B.n964 B.n499 163.367
R2300 B.n972 B.n499 163.367
R2301 B.n972 B.n497 163.367
R2302 B.n976 B.n497 163.367
R2303 B.n976 B.n491 163.367
R2304 B.n984 B.n491 163.367
R2305 B.n984 B.n489 163.367
R2306 B.n988 B.n489 163.367
R2307 B.n988 B.n483 163.367
R2308 B.n996 B.n483 163.367
R2309 B.n996 B.n481 163.367
R2310 B.n1000 B.n481 163.367
R2311 B.n1000 B.n475 163.367
R2312 B.n1008 B.n475 163.367
R2313 B.n1008 B.n473 163.367
R2314 B.n1012 B.n473 163.367
R2315 B.n1012 B.n467 163.367
R2316 B.n1020 B.n467 163.367
R2317 B.n1020 B.n465 163.367
R2318 B.n1024 B.n465 163.367
R2319 B.n1024 B.n459 163.367
R2320 B.n1032 B.n459 163.367
R2321 B.n1032 B.n457 163.367
R2322 B.n1036 B.n457 163.367
R2323 B.n1036 B.n451 163.367
R2324 B.n1045 B.n451 163.367
R2325 B.n1045 B.n449 163.367
R2326 B.n1049 B.n449 163.367
R2327 B.n1049 B.n444 163.367
R2328 B.n1058 B.n444 163.367
R2329 B.n1058 B.n442 163.367
R2330 B.n1062 B.n442 163.367
R2331 B.n1062 B.n2 163.367
R2332 B.n1266 B.n2 163.367
R2333 B.n1266 B.n3 163.367
R2334 B.n1262 B.n3 163.367
R2335 B.n1262 B.n9 163.367
R2336 B.n1258 B.n9 163.367
R2337 B.n1258 B.n11 163.367
R2338 B.n1254 B.n11 163.367
R2339 B.n1254 B.n15 163.367
R2340 B.n1250 B.n15 163.367
R2341 B.n1250 B.n17 163.367
R2342 B.n1246 B.n17 163.367
R2343 B.n1246 B.n23 163.367
R2344 B.n1242 B.n23 163.367
R2345 B.n1242 B.n25 163.367
R2346 B.n1238 B.n25 163.367
R2347 B.n1238 B.n30 163.367
R2348 B.n1234 B.n30 163.367
R2349 B.n1234 B.n32 163.367
R2350 B.n1230 B.n32 163.367
R2351 B.n1230 B.n37 163.367
R2352 B.n1226 B.n37 163.367
R2353 B.n1226 B.n39 163.367
R2354 B.n1222 B.n39 163.367
R2355 B.n1222 B.n44 163.367
R2356 B.n1218 B.n44 163.367
R2357 B.n1218 B.n46 163.367
R2358 B.n1214 B.n46 163.367
R2359 B.n1214 B.n51 163.367
R2360 B.n1210 B.n51 163.367
R2361 B.n1210 B.n53 163.367
R2362 B.n1206 B.n53 163.367
R2363 B.n1206 B.n58 163.367
R2364 B.n1202 B.n58 163.367
R2365 B.n1202 B.n60 163.367
R2366 B.n1198 B.n60 163.367
R2367 B.n1198 B.n65 163.367
R2368 B.n1194 B.n65 163.367
R2369 B.n1194 B.n67 163.367
R2370 B.n1190 B.n67 163.367
R2371 B.n1190 B.n72 163.367
R2372 B.n1186 B.n72 163.367
R2373 B.n1186 B.n74 163.367
R2374 B.n1182 B.n74 163.367
R2375 B.n1182 B.n79 163.367
R2376 B.n1178 B.n79 163.367
R2377 B.n1178 B.n81 163.367
R2378 B.n1174 B.n81 163.367
R2379 B.n1174 B.n86 163.367
R2380 B.n1170 B.n86 163.367
R2381 B.n1170 B.n88 163.367
R2382 B.n1166 B.n88 163.367
R2383 B.n1166 B.n92 163.367
R2384 B.n1162 B.n92 163.367
R2385 B.n1162 B.n94 163.367
R2386 B.n1158 B.n94 163.367
R2387 B.n1158 B.n100 163.367
R2388 B.n1154 B.n100 163.367
R2389 B.n1154 B.n102 163.367
R2390 B.n1150 B.n102 163.367
R2391 B.n1150 B.n107 163.367
R2392 B.n884 B.n554 163.367
R2393 B.n884 B.n620 163.367
R2394 B.n880 B.n879 163.367
R2395 B.n876 B.n875 163.367
R2396 B.n872 B.n871 163.367
R2397 B.n868 B.n867 163.367
R2398 B.n864 B.n863 163.367
R2399 B.n860 B.n859 163.367
R2400 B.n856 B.n855 163.367
R2401 B.n852 B.n851 163.367
R2402 B.n848 B.n847 163.367
R2403 B.n844 B.n843 163.367
R2404 B.n840 B.n839 163.367
R2405 B.n836 B.n835 163.367
R2406 B.n832 B.n831 163.367
R2407 B.n828 B.n827 163.367
R2408 B.n824 B.n823 163.367
R2409 B.n820 B.n819 163.367
R2410 B.n816 B.n815 163.367
R2411 B.n812 B.n811 163.367
R2412 B.n808 B.n807 163.367
R2413 B.n804 B.n803 163.367
R2414 B.n800 B.n799 163.367
R2415 B.n796 B.n795 163.367
R2416 B.n792 B.n791 163.367
R2417 B.n788 B.n787 163.367
R2418 B.n784 B.n783 163.367
R2419 B.n780 B.n779 163.367
R2420 B.n776 B.n775 163.367
R2421 B.n772 B.n771 163.367
R2422 B.n768 B.n767 163.367
R2423 B.n764 B.n763 163.367
R2424 B.n760 B.n759 163.367
R2425 B.n756 B.n755 163.367
R2426 B.n752 B.n751 163.367
R2427 B.n748 B.n747 163.367
R2428 B.n744 B.n743 163.367
R2429 B.n740 B.n739 163.367
R2430 B.n736 B.n735 163.367
R2431 B.n732 B.n731 163.367
R2432 B.n728 B.n727 163.367
R2433 B.n724 B.n723 163.367
R2434 B.n720 B.n719 163.367
R2435 B.n716 B.n715 163.367
R2436 B.n712 B.n711 163.367
R2437 B.n708 B.n707 163.367
R2438 B.n704 B.n703 163.367
R2439 B.n700 B.n699 163.367
R2440 B.n696 B.n695 163.367
R2441 B.n692 B.n691 163.367
R2442 B.n688 B.n687 163.367
R2443 B.n684 B.n683 163.367
R2444 B.n680 B.n679 163.367
R2445 B.n676 B.n675 163.367
R2446 B.n672 B.n671 163.367
R2447 B.n668 B.n667 163.367
R2448 B.n664 B.n663 163.367
R2449 B.n660 B.n659 163.367
R2450 B.n656 B.n655 163.367
R2451 B.n652 B.n651 163.367
R2452 B.n648 B.n647 163.367
R2453 B.n644 B.n643 163.367
R2454 B.n640 B.n639 163.367
R2455 B.n636 B.n635 163.367
R2456 B.n632 B.n631 163.367
R2457 B.n628 B.n619 163.367
R2458 B.n893 B.n550 163.367
R2459 B.n893 B.n548 163.367
R2460 B.n897 B.n548 163.367
R2461 B.n897 B.n542 163.367
R2462 B.n905 B.n542 163.367
R2463 B.n905 B.n540 163.367
R2464 B.n909 B.n540 163.367
R2465 B.n909 B.n535 163.367
R2466 B.n918 B.n535 163.367
R2467 B.n918 B.n533 163.367
R2468 B.n922 B.n533 163.367
R2469 B.n922 B.n527 163.367
R2470 B.n930 B.n527 163.367
R2471 B.n930 B.n525 163.367
R2472 B.n934 B.n525 163.367
R2473 B.n934 B.n519 163.367
R2474 B.n942 B.n519 163.367
R2475 B.n942 B.n517 163.367
R2476 B.n946 B.n517 163.367
R2477 B.n946 B.n511 163.367
R2478 B.n954 B.n511 163.367
R2479 B.n954 B.n509 163.367
R2480 B.n958 B.n509 163.367
R2481 B.n958 B.n503 163.367
R2482 B.n966 B.n503 163.367
R2483 B.n966 B.n501 163.367
R2484 B.n970 B.n501 163.367
R2485 B.n970 B.n495 163.367
R2486 B.n978 B.n495 163.367
R2487 B.n978 B.n493 163.367
R2488 B.n982 B.n493 163.367
R2489 B.n982 B.n487 163.367
R2490 B.n990 B.n487 163.367
R2491 B.n990 B.n485 163.367
R2492 B.n994 B.n485 163.367
R2493 B.n994 B.n479 163.367
R2494 B.n1002 B.n479 163.367
R2495 B.n1002 B.n477 163.367
R2496 B.n1006 B.n477 163.367
R2497 B.n1006 B.n470 163.367
R2498 B.n1014 B.n470 163.367
R2499 B.n1014 B.n468 163.367
R2500 B.n1018 B.n468 163.367
R2501 B.n1018 B.n463 163.367
R2502 B.n1026 B.n463 163.367
R2503 B.n1026 B.n461 163.367
R2504 B.n1030 B.n461 163.367
R2505 B.n1030 B.n455 163.367
R2506 B.n1038 B.n455 163.367
R2507 B.n1038 B.n453 163.367
R2508 B.n1042 B.n453 163.367
R2509 B.n1042 B.n448 163.367
R2510 B.n1051 B.n448 163.367
R2511 B.n1051 B.n446 163.367
R2512 B.n1056 B.n446 163.367
R2513 B.n1056 B.n440 163.367
R2514 B.n1064 B.n440 163.367
R2515 B.n1065 B.n1064 163.367
R2516 B.n1065 B.n5 163.367
R2517 B.n6 B.n5 163.367
R2518 B.n7 B.n6 163.367
R2519 B.n1070 B.n7 163.367
R2520 B.n1070 B.n12 163.367
R2521 B.n13 B.n12 163.367
R2522 B.n14 B.n13 163.367
R2523 B.n1075 B.n14 163.367
R2524 B.n1075 B.n19 163.367
R2525 B.n20 B.n19 163.367
R2526 B.n21 B.n20 163.367
R2527 B.n1080 B.n21 163.367
R2528 B.n1080 B.n26 163.367
R2529 B.n27 B.n26 163.367
R2530 B.n28 B.n27 163.367
R2531 B.n1085 B.n28 163.367
R2532 B.n1085 B.n33 163.367
R2533 B.n34 B.n33 163.367
R2534 B.n35 B.n34 163.367
R2535 B.n1090 B.n35 163.367
R2536 B.n1090 B.n40 163.367
R2537 B.n41 B.n40 163.367
R2538 B.n42 B.n41 163.367
R2539 B.n1095 B.n42 163.367
R2540 B.n1095 B.n47 163.367
R2541 B.n48 B.n47 163.367
R2542 B.n49 B.n48 163.367
R2543 B.n1100 B.n49 163.367
R2544 B.n1100 B.n54 163.367
R2545 B.n55 B.n54 163.367
R2546 B.n56 B.n55 163.367
R2547 B.n1105 B.n56 163.367
R2548 B.n1105 B.n61 163.367
R2549 B.n62 B.n61 163.367
R2550 B.n63 B.n62 163.367
R2551 B.n1110 B.n63 163.367
R2552 B.n1110 B.n68 163.367
R2553 B.n69 B.n68 163.367
R2554 B.n70 B.n69 163.367
R2555 B.n1115 B.n70 163.367
R2556 B.n1115 B.n75 163.367
R2557 B.n76 B.n75 163.367
R2558 B.n77 B.n76 163.367
R2559 B.n1120 B.n77 163.367
R2560 B.n1120 B.n82 163.367
R2561 B.n83 B.n82 163.367
R2562 B.n84 B.n83 163.367
R2563 B.n1125 B.n84 163.367
R2564 B.n1125 B.n89 163.367
R2565 B.n90 B.n89 163.367
R2566 B.n91 B.n90 163.367
R2567 B.n1130 B.n91 163.367
R2568 B.n1130 B.n96 163.367
R2569 B.n97 B.n96 163.367
R2570 B.n98 B.n97 163.367
R2571 B.n1135 B.n98 163.367
R2572 B.n1135 B.n103 163.367
R2573 B.n104 B.n103 163.367
R2574 B.n105 B.n104 163.367
R2575 B.n175 B.n105 163.367
R2576 B.n180 B.n109 163.367
R2577 B.n184 B.n183 163.367
R2578 B.n188 B.n187 163.367
R2579 B.n192 B.n191 163.367
R2580 B.n196 B.n195 163.367
R2581 B.n200 B.n199 163.367
R2582 B.n204 B.n203 163.367
R2583 B.n208 B.n207 163.367
R2584 B.n212 B.n211 163.367
R2585 B.n216 B.n215 163.367
R2586 B.n220 B.n219 163.367
R2587 B.n224 B.n223 163.367
R2588 B.n228 B.n227 163.367
R2589 B.n232 B.n231 163.367
R2590 B.n236 B.n235 163.367
R2591 B.n240 B.n239 163.367
R2592 B.n244 B.n243 163.367
R2593 B.n248 B.n247 163.367
R2594 B.n252 B.n251 163.367
R2595 B.n256 B.n255 163.367
R2596 B.n260 B.n259 163.367
R2597 B.n264 B.n263 163.367
R2598 B.n268 B.n267 163.367
R2599 B.n272 B.n271 163.367
R2600 B.n276 B.n275 163.367
R2601 B.n280 B.n279 163.367
R2602 B.n284 B.n283 163.367
R2603 B.n288 B.n287 163.367
R2604 B.n292 B.n291 163.367
R2605 B.n296 B.n295 163.367
R2606 B.n301 B.n300 163.367
R2607 B.n305 B.n304 163.367
R2608 B.n309 B.n308 163.367
R2609 B.n313 B.n312 163.367
R2610 B.n317 B.n316 163.367
R2611 B.n322 B.n321 163.367
R2612 B.n326 B.n325 163.367
R2613 B.n330 B.n329 163.367
R2614 B.n334 B.n333 163.367
R2615 B.n338 B.n337 163.367
R2616 B.n342 B.n341 163.367
R2617 B.n346 B.n345 163.367
R2618 B.n350 B.n349 163.367
R2619 B.n354 B.n353 163.367
R2620 B.n358 B.n357 163.367
R2621 B.n362 B.n361 163.367
R2622 B.n366 B.n365 163.367
R2623 B.n370 B.n369 163.367
R2624 B.n374 B.n373 163.367
R2625 B.n378 B.n377 163.367
R2626 B.n382 B.n381 163.367
R2627 B.n386 B.n385 163.367
R2628 B.n390 B.n389 163.367
R2629 B.n394 B.n393 163.367
R2630 B.n398 B.n397 163.367
R2631 B.n402 B.n401 163.367
R2632 B.n406 B.n405 163.367
R2633 B.n410 B.n409 163.367
R2634 B.n414 B.n413 163.367
R2635 B.n418 B.n417 163.367
R2636 B.n422 B.n421 163.367
R2637 B.n426 B.n425 163.367
R2638 B.n430 B.n429 163.367
R2639 B.n434 B.n433 163.367
R2640 B.n436 B.n174 163.367
R2641 B.n887 B.n886 71.676
R2642 B.n620 B.n555 71.676
R2643 B.n879 B.n556 71.676
R2644 B.n875 B.n557 71.676
R2645 B.n871 B.n558 71.676
R2646 B.n867 B.n559 71.676
R2647 B.n863 B.n560 71.676
R2648 B.n859 B.n561 71.676
R2649 B.n855 B.n562 71.676
R2650 B.n851 B.n563 71.676
R2651 B.n847 B.n564 71.676
R2652 B.n843 B.n565 71.676
R2653 B.n839 B.n566 71.676
R2654 B.n835 B.n567 71.676
R2655 B.n831 B.n568 71.676
R2656 B.n827 B.n569 71.676
R2657 B.n823 B.n570 71.676
R2658 B.n819 B.n571 71.676
R2659 B.n815 B.n572 71.676
R2660 B.n811 B.n573 71.676
R2661 B.n807 B.n574 71.676
R2662 B.n803 B.n575 71.676
R2663 B.n799 B.n576 71.676
R2664 B.n795 B.n577 71.676
R2665 B.n791 B.n578 71.676
R2666 B.n787 B.n579 71.676
R2667 B.n783 B.n580 71.676
R2668 B.n779 B.n581 71.676
R2669 B.n775 B.n582 71.676
R2670 B.n771 B.n583 71.676
R2671 B.n767 B.n584 71.676
R2672 B.n763 B.n585 71.676
R2673 B.n759 B.n586 71.676
R2674 B.n755 B.n587 71.676
R2675 B.n751 B.n588 71.676
R2676 B.n747 B.n589 71.676
R2677 B.n743 B.n590 71.676
R2678 B.n739 B.n591 71.676
R2679 B.n735 B.n592 71.676
R2680 B.n731 B.n593 71.676
R2681 B.n727 B.n594 71.676
R2682 B.n723 B.n595 71.676
R2683 B.n719 B.n596 71.676
R2684 B.n715 B.n597 71.676
R2685 B.n711 B.n598 71.676
R2686 B.n707 B.n599 71.676
R2687 B.n703 B.n600 71.676
R2688 B.n699 B.n601 71.676
R2689 B.n695 B.n602 71.676
R2690 B.n691 B.n603 71.676
R2691 B.n687 B.n604 71.676
R2692 B.n683 B.n605 71.676
R2693 B.n679 B.n606 71.676
R2694 B.n675 B.n607 71.676
R2695 B.n671 B.n608 71.676
R2696 B.n667 B.n609 71.676
R2697 B.n663 B.n610 71.676
R2698 B.n659 B.n611 71.676
R2699 B.n655 B.n612 71.676
R2700 B.n651 B.n613 71.676
R2701 B.n647 B.n614 71.676
R2702 B.n643 B.n615 71.676
R2703 B.n639 B.n616 71.676
R2704 B.n635 B.n617 71.676
R2705 B.n631 B.n618 71.676
R2706 B.n1146 B.n1145 71.676
R2707 B.n180 B.n110 71.676
R2708 B.n184 B.n111 71.676
R2709 B.n188 B.n112 71.676
R2710 B.n192 B.n113 71.676
R2711 B.n196 B.n114 71.676
R2712 B.n200 B.n115 71.676
R2713 B.n204 B.n116 71.676
R2714 B.n208 B.n117 71.676
R2715 B.n212 B.n118 71.676
R2716 B.n216 B.n119 71.676
R2717 B.n220 B.n120 71.676
R2718 B.n224 B.n121 71.676
R2719 B.n228 B.n122 71.676
R2720 B.n232 B.n123 71.676
R2721 B.n236 B.n124 71.676
R2722 B.n240 B.n125 71.676
R2723 B.n244 B.n126 71.676
R2724 B.n248 B.n127 71.676
R2725 B.n252 B.n128 71.676
R2726 B.n256 B.n129 71.676
R2727 B.n260 B.n130 71.676
R2728 B.n264 B.n131 71.676
R2729 B.n268 B.n132 71.676
R2730 B.n272 B.n133 71.676
R2731 B.n276 B.n134 71.676
R2732 B.n280 B.n135 71.676
R2733 B.n284 B.n136 71.676
R2734 B.n288 B.n137 71.676
R2735 B.n292 B.n138 71.676
R2736 B.n296 B.n139 71.676
R2737 B.n301 B.n140 71.676
R2738 B.n305 B.n141 71.676
R2739 B.n309 B.n142 71.676
R2740 B.n313 B.n143 71.676
R2741 B.n317 B.n144 71.676
R2742 B.n322 B.n145 71.676
R2743 B.n326 B.n146 71.676
R2744 B.n330 B.n147 71.676
R2745 B.n334 B.n148 71.676
R2746 B.n338 B.n149 71.676
R2747 B.n342 B.n150 71.676
R2748 B.n346 B.n151 71.676
R2749 B.n350 B.n152 71.676
R2750 B.n354 B.n153 71.676
R2751 B.n358 B.n154 71.676
R2752 B.n362 B.n155 71.676
R2753 B.n366 B.n156 71.676
R2754 B.n370 B.n157 71.676
R2755 B.n374 B.n158 71.676
R2756 B.n378 B.n159 71.676
R2757 B.n382 B.n160 71.676
R2758 B.n386 B.n161 71.676
R2759 B.n390 B.n162 71.676
R2760 B.n394 B.n163 71.676
R2761 B.n398 B.n164 71.676
R2762 B.n402 B.n165 71.676
R2763 B.n406 B.n166 71.676
R2764 B.n410 B.n167 71.676
R2765 B.n414 B.n168 71.676
R2766 B.n418 B.n169 71.676
R2767 B.n422 B.n170 71.676
R2768 B.n426 B.n171 71.676
R2769 B.n430 B.n172 71.676
R2770 B.n434 B.n173 71.676
R2771 B.n1143 B.n174 71.676
R2772 B.n1143 B.n1142 71.676
R2773 B.n436 B.n173 71.676
R2774 B.n433 B.n172 71.676
R2775 B.n429 B.n171 71.676
R2776 B.n425 B.n170 71.676
R2777 B.n421 B.n169 71.676
R2778 B.n417 B.n168 71.676
R2779 B.n413 B.n167 71.676
R2780 B.n409 B.n166 71.676
R2781 B.n405 B.n165 71.676
R2782 B.n401 B.n164 71.676
R2783 B.n397 B.n163 71.676
R2784 B.n393 B.n162 71.676
R2785 B.n389 B.n161 71.676
R2786 B.n385 B.n160 71.676
R2787 B.n381 B.n159 71.676
R2788 B.n377 B.n158 71.676
R2789 B.n373 B.n157 71.676
R2790 B.n369 B.n156 71.676
R2791 B.n365 B.n155 71.676
R2792 B.n361 B.n154 71.676
R2793 B.n357 B.n153 71.676
R2794 B.n353 B.n152 71.676
R2795 B.n349 B.n151 71.676
R2796 B.n345 B.n150 71.676
R2797 B.n341 B.n149 71.676
R2798 B.n337 B.n148 71.676
R2799 B.n333 B.n147 71.676
R2800 B.n329 B.n146 71.676
R2801 B.n325 B.n145 71.676
R2802 B.n321 B.n144 71.676
R2803 B.n316 B.n143 71.676
R2804 B.n312 B.n142 71.676
R2805 B.n308 B.n141 71.676
R2806 B.n304 B.n140 71.676
R2807 B.n300 B.n139 71.676
R2808 B.n295 B.n138 71.676
R2809 B.n291 B.n137 71.676
R2810 B.n287 B.n136 71.676
R2811 B.n283 B.n135 71.676
R2812 B.n279 B.n134 71.676
R2813 B.n275 B.n133 71.676
R2814 B.n271 B.n132 71.676
R2815 B.n267 B.n131 71.676
R2816 B.n263 B.n130 71.676
R2817 B.n259 B.n129 71.676
R2818 B.n255 B.n128 71.676
R2819 B.n251 B.n127 71.676
R2820 B.n247 B.n126 71.676
R2821 B.n243 B.n125 71.676
R2822 B.n239 B.n124 71.676
R2823 B.n235 B.n123 71.676
R2824 B.n231 B.n122 71.676
R2825 B.n227 B.n121 71.676
R2826 B.n223 B.n120 71.676
R2827 B.n219 B.n119 71.676
R2828 B.n215 B.n118 71.676
R2829 B.n211 B.n117 71.676
R2830 B.n207 B.n116 71.676
R2831 B.n203 B.n115 71.676
R2832 B.n199 B.n114 71.676
R2833 B.n195 B.n113 71.676
R2834 B.n191 B.n112 71.676
R2835 B.n187 B.n111 71.676
R2836 B.n183 B.n110 71.676
R2837 B.n1145 B.n109 71.676
R2838 B.n886 B.n554 71.676
R2839 B.n880 B.n555 71.676
R2840 B.n876 B.n556 71.676
R2841 B.n872 B.n557 71.676
R2842 B.n868 B.n558 71.676
R2843 B.n864 B.n559 71.676
R2844 B.n860 B.n560 71.676
R2845 B.n856 B.n561 71.676
R2846 B.n852 B.n562 71.676
R2847 B.n848 B.n563 71.676
R2848 B.n844 B.n564 71.676
R2849 B.n840 B.n565 71.676
R2850 B.n836 B.n566 71.676
R2851 B.n832 B.n567 71.676
R2852 B.n828 B.n568 71.676
R2853 B.n824 B.n569 71.676
R2854 B.n820 B.n570 71.676
R2855 B.n816 B.n571 71.676
R2856 B.n812 B.n572 71.676
R2857 B.n808 B.n573 71.676
R2858 B.n804 B.n574 71.676
R2859 B.n800 B.n575 71.676
R2860 B.n796 B.n576 71.676
R2861 B.n792 B.n577 71.676
R2862 B.n788 B.n578 71.676
R2863 B.n784 B.n579 71.676
R2864 B.n780 B.n580 71.676
R2865 B.n776 B.n581 71.676
R2866 B.n772 B.n582 71.676
R2867 B.n768 B.n583 71.676
R2868 B.n764 B.n584 71.676
R2869 B.n760 B.n585 71.676
R2870 B.n756 B.n586 71.676
R2871 B.n752 B.n587 71.676
R2872 B.n748 B.n588 71.676
R2873 B.n744 B.n589 71.676
R2874 B.n740 B.n590 71.676
R2875 B.n736 B.n591 71.676
R2876 B.n732 B.n592 71.676
R2877 B.n728 B.n593 71.676
R2878 B.n724 B.n594 71.676
R2879 B.n720 B.n595 71.676
R2880 B.n716 B.n596 71.676
R2881 B.n712 B.n597 71.676
R2882 B.n708 B.n598 71.676
R2883 B.n704 B.n599 71.676
R2884 B.n700 B.n600 71.676
R2885 B.n696 B.n601 71.676
R2886 B.n692 B.n602 71.676
R2887 B.n688 B.n603 71.676
R2888 B.n684 B.n604 71.676
R2889 B.n680 B.n605 71.676
R2890 B.n676 B.n606 71.676
R2891 B.n672 B.n607 71.676
R2892 B.n668 B.n608 71.676
R2893 B.n664 B.n609 71.676
R2894 B.n660 B.n610 71.676
R2895 B.n656 B.n611 71.676
R2896 B.n652 B.n612 71.676
R2897 B.n648 B.n613 71.676
R2898 B.n644 B.n614 71.676
R2899 B.n640 B.n615 71.676
R2900 B.n636 B.n616 71.676
R2901 B.n632 B.n617 71.676
R2902 B.n628 B.n618 71.676
R2903 B.n625 B.n624 67.1035
R2904 B.n622 B.n621 67.1035
R2905 B.n179 B.n178 67.1035
R2906 B.n177 B.n176 67.1035
R2907 B.n626 B.n625 59.5399
R2908 B.n623 B.n622 59.5399
R2909 B.n298 B.n179 59.5399
R2910 B.n319 B.n177 59.5399
R2911 B.n885 B.n551 56.4108
R2912 B.n1144 B.n106 56.4108
R2913 B.n1148 B.n1147 33.8737
R2914 B.n1141 B.n1140 33.8737
R2915 B.n627 B.n549 33.8737
R2916 B.n889 B.n888 33.8737
R2917 B.n892 B.n551 31.1867
R2918 B.n892 B.n547 31.1867
R2919 B.n898 B.n547 31.1867
R2920 B.n898 B.n543 31.1867
R2921 B.n904 B.n543 31.1867
R2922 B.n904 B.n539 31.1867
R2923 B.n911 B.n539 31.1867
R2924 B.n911 B.n910 31.1867
R2925 B.n917 B.n532 31.1867
R2926 B.n923 B.n532 31.1867
R2927 B.n923 B.n528 31.1867
R2928 B.n929 B.n528 31.1867
R2929 B.n929 B.n524 31.1867
R2930 B.n935 B.n524 31.1867
R2931 B.n935 B.n520 31.1867
R2932 B.n941 B.n520 31.1867
R2933 B.n941 B.n516 31.1867
R2934 B.n947 B.n516 31.1867
R2935 B.n947 B.n512 31.1867
R2936 B.n953 B.n512 31.1867
R2937 B.n959 B.n508 31.1867
R2938 B.n959 B.n504 31.1867
R2939 B.n965 B.n504 31.1867
R2940 B.n965 B.n500 31.1867
R2941 B.n971 B.n500 31.1867
R2942 B.n971 B.n496 31.1867
R2943 B.n977 B.n496 31.1867
R2944 B.n977 B.n492 31.1867
R2945 B.n983 B.n492 31.1867
R2946 B.n989 B.n488 31.1867
R2947 B.n989 B.n484 31.1867
R2948 B.n995 B.n484 31.1867
R2949 B.n995 B.n480 31.1867
R2950 B.n1001 B.n480 31.1867
R2951 B.n1001 B.n476 31.1867
R2952 B.n1007 B.n476 31.1867
R2953 B.n1007 B.n471 31.1867
R2954 B.n1013 B.n471 31.1867
R2955 B.n1013 B.n472 31.1867
R2956 B.n1019 B.n464 31.1867
R2957 B.n1025 B.n464 31.1867
R2958 B.n1025 B.n460 31.1867
R2959 B.n1031 B.n460 31.1867
R2960 B.n1031 B.n456 31.1867
R2961 B.n1037 B.n456 31.1867
R2962 B.n1037 B.n452 31.1867
R2963 B.n1044 B.n452 31.1867
R2964 B.n1044 B.n1043 31.1867
R2965 B.n1050 B.n445 31.1867
R2966 B.n1057 B.n445 31.1867
R2967 B.n1057 B.n441 31.1867
R2968 B.n1063 B.n441 31.1867
R2969 B.n1063 B.n4 31.1867
R2970 B.n1265 B.n4 31.1867
R2971 B.n1265 B.n1264 31.1867
R2972 B.n1264 B.n1263 31.1867
R2973 B.n1263 B.n8 31.1867
R2974 B.n1257 B.n8 31.1867
R2975 B.n1257 B.n1256 31.1867
R2976 B.n1256 B.n1255 31.1867
R2977 B.n1249 B.n18 31.1867
R2978 B.n1249 B.n1248 31.1867
R2979 B.n1248 B.n1247 31.1867
R2980 B.n1247 B.n22 31.1867
R2981 B.n1241 B.n22 31.1867
R2982 B.n1241 B.n1240 31.1867
R2983 B.n1240 B.n1239 31.1867
R2984 B.n1239 B.n29 31.1867
R2985 B.n1233 B.n29 31.1867
R2986 B.n1232 B.n1231 31.1867
R2987 B.n1231 B.n36 31.1867
R2988 B.n1225 B.n36 31.1867
R2989 B.n1225 B.n1224 31.1867
R2990 B.n1224 B.n1223 31.1867
R2991 B.n1223 B.n43 31.1867
R2992 B.n1217 B.n43 31.1867
R2993 B.n1217 B.n1216 31.1867
R2994 B.n1216 B.n1215 31.1867
R2995 B.n1215 B.n50 31.1867
R2996 B.n1209 B.n1208 31.1867
R2997 B.n1208 B.n1207 31.1867
R2998 B.n1207 B.n57 31.1867
R2999 B.n1201 B.n57 31.1867
R3000 B.n1201 B.n1200 31.1867
R3001 B.n1200 B.n1199 31.1867
R3002 B.n1199 B.n64 31.1867
R3003 B.n1193 B.n64 31.1867
R3004 B.n1193 B.n1192 31.1867
R3005 B.n1191 B.n71 31.1867
R3006 B.n1185 B.n71 31.1867
R3007 B.n1185 B.n1184 31.1867
R3008 B.n1184 B.n1183 31.1867
R3009 B.n1183 B.n78 31.1867
R3010 B.n1177 B.n78 31.1867
R3011 B.n1177 B.n1176 31.1867
R3012 B.n1176 B.n1175 31.1867
R3013 B.n1175 B.n85 31.1867
R3014 B.n1169 B.n85 31.1867
R3015 B.n1169 B.n1168 31.1867
R3016 B.n1168 B.n1167 31.1867
R3017 B.n1161 B.n95 31.1867
R3018 B.n1161 B.n1160 31.1867
R3019 B.n1160 B.n1159 31.1867
R3020 B.n1159 B.n99 31.1867
R3021 B.n1153 B.n99 31.1867
R3022 B.n1153 B.n1152 31.1867
R3023 B.n1152 B.n1151 31.1867
R3024 B.n1151 B.n106 31.1867
R3025 B.n983 B.t5 29.8108
R3026 B.n1209 B.t3 29.8108
R3027 B.n1019 B.t0 27.0591
R3028 B.n1233 B.t4 27.0591
R3029 B.n953 B.t7 24.3074
R3030 B.t6 B.n1191 24.3074
R3031 B.n1050 B.t2 21.5556
R3032 B.n1255 B.t1 21.5556
R3033 B.n917 B.t9 18.8039
R3034 B.n1167 B.t16 18.8039
R3035 B B.n1267 18.0485
R3036 B.n910 B.t9 12.3832
R3037 B.n95 B.t16 12.3832
R3038 B.n1147 B.n108 10.6151
R3039 B.n181 B.n108 10.6151
R3040 B.n182 B.n181 10.6151
R3041 B.n185 B.n182 10.6151
R3042 B.n186 B.n185 10.6151
R3043 B.n189 B.n186 10.6151
R3044 B.n190 B.n189 10.6151
R3045 B.n193 B.n190 10.6151
R3046 B.n194 B.n193 10.6151
R3047 B.n197 B.n194 10.6151
R3048 B.n198 B.n197 10.6151
R3049 B.n201 B.n198 10.6151
R3050 B.n202 B.n201 10.6151
R3051 B.n205 B.n202 10.6151
R3052 B.n206 B.n205 10.6151
R3053 B.n209 B.n206 10.6151
R3054 B.n210 B.n209 10.6151
R3055 B.n213 B.n210 10.6151
R3056 B.n214 B.n213 10.6151
R3057 B.n217 B.n214 10.6151
R3058 B.n218 B.n217 10.6151
R3059 B.n221 B.n218 10.6151
R3060 B.n222 B.n221 10.6151
R3061 B.n225 B.n222 10.6151
R3062 B.n226 B.n225 10.6151
R3063 B.n229 B.n226 10.6151
R3064 B.n230 B.n229 10.6151
R3065 B.n233 B.n230 10.6151
R3066 B.n234 B.n233 10.6151
R3067 B.n237 B.n234 10.6151
R3068 B.n238 B.n237 10.6151
R3069 B.n241 B.n238 10.6151
R3070 B.n242 B.n241 10.6151
R3071 B.n245 B.n242 10.6151
R3072 B.n246 B.n245 10.6151
R3073 B.n249 B.n246 10.6151
R3074 B.n250 B.n249 10.6151
R3075 B.n253 B.n250 10.6151
R3076 B.n254 B.n253 10.6151
R3077 B.n257 B.n254 10.6151
R3078 B.n258 B.n257 10.6151
R3079 B.n261 B.n258 10.6151
R3080 B.n262 B.n261 10.6151
R3081 B.n265 B.n262 10.6151
R3082 B.n266 B.n265 10.6151
R3083 B.n269 B.n266 10.6151
R3084 B.n270 B.n269 10.6151
R3085 B.n273 B.n270 10.6151
R3086 B.n274 B.n273 10.6151
R3087 B.n277 B.n274 10.6151
R3088 B.n278 B.n277 10.6151
R3089 B.n281 B.n278 10.6151
R3090 B.n282 B.n281 10.6151
R3091 B.n285 B.n282 10.6151
R3092 B.n286 B.n285 10.6151
R3093 B.n289 B.n286 10.6151
R3094 B.n290 B.n289 10.6151
R3095 B.n293 B.n290 10.6151
R3096 B.n294 B.n293 10.6151
R3097 B.n297 B.n294 10.6151
R3098 B.n302 B.n299 10.6151
R3099 B.n303 B.n302 10.6151
R3100 B.n306 B.n303 10.6151
R3101 B.n307 B.n306 10.6151
R3102 B.n310 B.n307 10.6151
R3103 B.n311 B.n310 10.6151
R3104 B.n314 B.n311 10.6151
R3105 B.n315 B.n314 10.6151
R3106 B.n318 B.n315 10.6151
R3107 B.n323 B.n320 10.6151
R3108 B.n324 B.n323 10.6151
R3109 B.n327 B.n324 10.6151
R3110 B.n328 B.n327 10.6151
R3111 B.n331 B.n328 10.6151
R3112 B.n332 B.n331 10.6151
R3113 B.n335 B.n332 10.6151
R3114 B.n336 B.n335 10.6151
R3115 B.n339 B.n336 10.6151
R3116 B.n340 B.n339 10.6151
R3117 B.n343 B.n340 10.6151
R3118 B.n344 B.n343 10.6151
R3119 B.n347 B.n344 10.6151
R3120 B.n348 B.n347 10.6151
R3121 B.n351 B.n348 10.6151
R3122 B.n352 B.n351 10.6151
R3123 B.n355 B.n352 10.6151
R3124 B.n356 B.n355 10.6151
R3125 B.n359 B.n356 10.6151
R3126 B.n360 B.n359 10.6151
R3127 B.n363 B.n360 10.6151
R3128 B.n364 B.n363 10.6151
R3129 B.n367 B.n364 10.6151
R3130 B.n368 B.n367 10.6151
R3131 B.n371 B.n368 10.6151
R3132 B.n372 B.n371 10.6151
R3133 B.n375 B.n372 10.6151
R3134 B.n376 B.n375 10.6151
R3135 B.n379 B.n376 10.6151
R3136 B.n380 B.n379 10.6151
R3137 B.n383 B.n380 10.6151
R3138 B.n384 B.n383 10.6151
R3139 B.n387 B.n384 10.6151
R3140 B.n388 B.n387 10.6151
R3141 B.n391 B.n388 10.6151
R3142 B.n392 B.n391 10.6151
R3143 B.n395 B.n392 10.6151
R3144 B.n396 B.n395 10.6151
R3145 B.n399 B.n396 10.6151
R3146 B.n400 B.n399 10.6151
R3147 B.n403 B.n400 10.6151
R3148 B.n404 B.n403 10.6151
R3149 B.n407 B.n404 10.6151
R3150 B.n408 B.n407 10.6151
R3151 B.n411 B.n408 10.6151
R3152 B.n412 B.n411 10.6151
R3153 B.n415 B.n412 10.6151
R3154 B.n416 B.n415 10.6151
R3155 B.n419 B.n416 10.6151
R3156 B.n420 B.n419 10.6151
R3157 B.n423 B.n420 10.6151
R3158 B.n424 B.n423 10.6151
R3159 B.n427 B.n424 10.6151
R3160 B.n428 B.n427 10.6151
R3161 B.n431 B.n428 10.6151
R3162 B.n432 B.n431 10.6151
R3163 B.n435 B.n432 10.6151
R3164 B.n437 B.n435 10.6151
R3165 B.n438 B.n437 10.6151
R3166 B.n1141 B.n438 10.6151
R3167 B.n894 B.n549 10.6151
R3168 B.n895 B.n894 10.6151
R3169 B.n896 B.n895 10.6151
R3170 B.n896 B.n541 10.6151
R3171 B.n906 B.n541 10.6151
R3172 B.n907 B.n906 10.6151
R3173 B.n908 B.n907 10.6151
R3174 B.n908 B.n534 10.6151
R3175 B.n919 B.n534 10.6151
R3176 B.n920 B.n919 10.6151
R3177 B.n921 B.n920 10.6151
R3178 B.n921 B.n526 10.6151
R3179 B.n931 B.n526 10.6151
R3180 B.n932 B.n931 10.6151
R3181 B.n933 B.n932 10.6151
R3182 B.n933 B.n518 10.6151
R3183 B.n943 B.n518 10.6151
R3184 B.n944 B.n943 10.6151
R3185 B.n945 B.n944 10.6151
R3186 B.n945 B.n510 10.6151
R3187 B.n955 B.n510 10.6151
R3188 B.n956 B.n955 10.6151
R3189 B.n957 B.n956 10.6151
R3190 B.n957 B.n502 10.6151
R3191 B.n967 B.n502 10.6151
R3192 B.n968 B.n967 10.6151
R3193 B.n969 B.n968 10.6151
R3194 B.n969 B.n494 10.6151
R3195 B.n979 B.n494 10.6151
R3196 B.n980 B.n979 10.6151
R3197 B.n981 B.n980 10.6151
R3198 B.n981 B.n486 10.6151
R3199 B.n991 B.n486 10.6151
R3200 B.n992 B.n991 10.6151
R3201 B.n993 B.n992 10.6151
R3202 B.n993 B.n478 10.6151
R3203 B.n1003 B.n478 10.6151
R3204 B.n1004 B.n1003 10.6151
R3205 B.n1005 B.n1004 10.6151
R3206 B.n1005 B.n469 10.6151
R3207 B.n1015 B.n469 10.6151
R3208 B.n1016 B.n1015 10.6151
R3209 B.n1017 B.n1016 10.6151
R3210 B.n1017 B.n462 10.6151
R3211 B.n1027 B.n462 10.6151
R3212 B.n1028 B.n1027 10.6151
R3213 B.n1029 B.n1028 10.6151
R3214 B.n1029 B.n454 10.6151
R3215 B.n1039 B.n454 10.6151
R3216 B.n1040 B.n1039 10.6151
R3217 B.n1041 B.n1040 10.6151
R3218 B.n1041 B.n447 10.6151
R3219 B.n1052 B.n447 10.6151
R3220 B.n1053 B.n1052 10.6151
R3221 B.n1055 B.n1053 10.6151
R3222 B.n1055 B.n1054 10.6151
R3223 B.n1054 B.n439 10.6151
R3224 B.n1066 B.n439 10.6151
R3225 B.n1067 B.n1066 10.6151
R3226 B.n1068 B.n1067 10.6151
R3227 B.n1069 B.n1068 10.6151
R3228 B.n1071 B.n1069 10.6151
R3229 B.n1072 B.n1071 10.6151
R3230 B.n1073 B.n1072 10.6151
R3231 B.n1074 B.n1073 10.6151
R3232 B.n1076 B.n1074 10.6151
R3233 B.n1077 B.n1076 10.6151
R3234 B.n1078 B.n1077 10.6151
R3235 B.n1079 B.n1078 10.6151
R3236 B.n1081 B.n1079 10.6151
R3237 B.n1082 B.n1081 10.6151
R3238 B.n1083 B.n1082 10.6151
R3239 B.n1084 B.n1083 10.6151
R3240 B.n1086 B.n1084 10.6151
R3241 B.n1087 B.n1086 10.6151
R3242 B.n1088 B.n1087 10.6151
R3243 B.n1089 B.n1088 10.6151
R3244 B.n1091 B.n1089 10.6151
R3245 B.n1092 B.n1091 10.6151
R3246 B.n1093 B.n1092 10.6151
R3247 B.n1094 B.n1093 10.6151
R3248 B.n1096 B.n1094 10.6151
R3249 B.n1097 B.n1096 10.6151
R3250 B.n1098 B.n1097 10.6151
R3251 B.n1099 B.n1098 10.6151
R3252 B.n1101 B.n1099 10.6151
R3253 B.n1102 B.n1101 10.6151
R3254 B.n1103 B.n1102 10.6151
R3255 B.n1104 B.n1103 10.6151
R3256 B.n1106 B.n1104 10.6151
R3257 B.n1107 B.n1106 10.6151
R3258 B.n1108 B.n1107 10.6151
R3259 B.n1109 B.n1108 10.6151
R3260 B.n1111 B.n1109 10.6151
R3261 B.n1112 B.n1111 10.6151
R3262 B.n1113 B.n1112 10.6151
R3263 B.n1114 B.n1113 10.6151
R3264 B.n1116 B.n1114 10.6151
R3265 B.n1117 B.n1116 10.6151
R3266 B.n1118 B.n1117 10.6151
R3267 B.n1119 B.n1118 10.6151
R3268 B.n1121 B.n1119 10.6151
R3269 B.n1122 B.n1121 10.6151
R3270 B.n1123 B.n1122 10.6151
R3271 B.n1124 B.n1123 10.6151
R3272 B.n1126 B.n1124 10.6151
R3273 B.n1127 B.n1126 10.6151
R3274 B.n1128 B.n1127 10.6151
R3275 B.n1129 B.n1128 10.6151
R3276 B.n1131 B.n1129 10.6151
R3277 B.n1132 B.n1131 10.6151
R3278 B.n1133 B.n1132 10.6151
R3279 B.n1134 B.n1133 10.6151
R3280 B.n1136 B.n1134 10.6151
R3281 B.n1137 B.n1136 10.6151
R3282 B.n1138 B.n1137 10.6151
R3283 B.n1139 B.n1138 10.6151
R3284 B.n1140 B.n1139 10.6151
R3285 B.n888 B.n553 10.6151
R3286 B.n883 B.n553 10.6151
R3287 B.n883 B.n882 10.6151
R3288 B.n882 B.n881 10.6151
R3289 B.n881 B.n878 10.6151
R3290 B.n878 B.n877 10.6151
R3291 B.n877 B.n874 10.6151
R3292 B.n874 B.n873 10.6151
R3293 B.n873 B.n870 10.6151
R3294 B.n870 B.n869 10.6151
R3295 B.n869 B.n866 10.6151
R3296 B.n866 B.n865 10.6151
R3297 B.n865 B.n862 10.6151
R3298 B.n862 B.n861 10.6151
R3299 B.n861 B.n858 10.6151
R3300 B.n858 B.n857 10.6151
R3301 B.n857 B.n854 10.6151
R3302 B.n854 B.n853 10.6151
R3303 B.n853 B.n850 10.6151
R3304 B.n850 B.n849 10.6151
R3305 B.n849 B.n846 10.6151
R3306 B.n846 B.n845 10.6151
R3307 B.n845 B.n842 10.6151
R3308 B.n842 B.n841 10.6151
R3309 B.n841 B.n838 10.6151
R3310 B.n838 B.n837 10.6151
R3311 B.n837 B.n834 10.6151
R3312 B.n834 B.n833 10.6151
R3313 B.n833 B.n830 10.6151
R3314 B.n830 B.n829 10.6151
R3315 B.n829 B.n826 10.6151
R3316 B.n826 B.n825 10.6151
R3317 B.n825 B.n822 10.6151
R3318 B.n822 B.n821 10.6151
R3319 B.n821 B.n818 10.6151
R3320 B.n818 B.n817 10.6151
R3321 B.n817 B.n814 10.6151
R3322 B.n814 B.n813 10.6151
R3323 B.n813 B.n810 10.6151
R3324 B.n810 B.n809 10.6151
R3325 B.n809 B.n806 10.6151
R3326 B.n806 B.n805 10.6151
R3327 B.n805 B.n802 10.6151
R3328 B.n802 B.n801 10.6151
R3329 B.n801 B.n798 10.6151
R3330 B.n798 B.n797 10.6151
R3331 B.n797 B.n794 10.6151
R3332 B.n794 B.n793 10.6151
R3333 B.n793 B.n790 10.6151
R3334 B.n790 B.n789 10.6151
R3335 B.n789 B.n786 10.6151
R3336 B.n786 B.n785 10.6151
R3337 B.n785 B.n782 10.6151
R3338 B.n782 B.n781 10.6151
R3339 B.n781 B.n778 10.6151
R3340 B.n778 B.n777 10.6151
R3341 B.n777 B.n774 10.6151
R3342 B.n774 B.n773 10.6151
R3343 B.n773 B.n770 10.6151
R3344 B.n770 B.n769 10.6151
R3345 B.n766 B.n765 10.6151
R3346 B.n765 B.n762 10.6151
R3347 B.n762 B.n761 10.6151
R3348 B.n761 B.n758 10.6151
R3349 B.n758 B.n757 10.6151
R3350 B.n757 B.n754 10.6151
R3351 B.n754 B.n753 10.6151
R3352 B.n753 B.n750 10.6151
R3353 B.n750 B.n749 10.6151
R3354 B.n746 B.n745 10.6151
R3355 B.n745 B.n742 10.6151
R3356 B.n742 B.n741 10.6151
R3357 B.n741 B.n738 10.6151
R3358 B.n738 B.n737 10.6151
R3359 B.n737 B.n734 10.6151
R3360 B.n734 B.n733 10.6151
R3361 B.n733 B.n730 10.6151
R3362 B.n730 B.n729 10.6151
R3363 B.n729 B.n726 10.6151
R3364 B.n726 B.n725 10.6151
R3365 B.n725 B.n722 10.6151
R3366 B.n722 B.n721 10.6151
R3367 B.n721 B.n718 10.6151
R3368 B.n718 B.n717 10.6151
R3369 B.n717 B.n714 10.6151
R3370 B.n714 B.n713 10.6151
R3371 B.n713 B.n710 10.6151
R3372 B.n710 B.n709 10.6151
R3373 B.n709 B.n706 10.6151
R3374 B.n706 B.n705 10.6151
R3375 B.n705 B.n702 10.6151
R3376 B.n702 B.n701 10.6151
R3377 B.n701 B.n698 10.6151
R3378 B.n698 B.n697 10.6151
R3379 B.n697 B.n694 10.6151
R3380 B.n694 B.n693 10.6151
R3381 B.n693 B.n690 10.6151
R3382 B.n690 B.n689 10.6151
R3383 B.n689 B.n686 10.6151
R3384 B.n686 B.n685 10.6151
R3385 B.n685 B.n682 10.6151
R3386 B.n682 B.n681 10.6151
R3387 B.n681 B.n678 10.6151
R3388 B.n678 B.n677 10.6151
R3389 B.n677 B.n674 10.6151
R3390 B.n674 B.n673 10.6151
R3391 B.n673 B.n670 10.6151
R3392 B.n670 B.n669 10.6151
R3393 B.n669 B.n666 10.6151
R3394 B.n666 B.n665 10.6151
R3395 B.n665 B.n662 10.6151
R3396 B.n662 B.n661 10.6151
R3397 B.n661 B.n658 10.6151
R3398 B.n658 B.n657 10.6151
R3399 B.n657 B.n654 10.6151
R3400 B.n654 B.n653 10.6151
R3401 B.n653 B.n650 10.6151
R3402 B.n650 B.n649 10.6151
R3403 B.n649 B.n646 10.6151
R3404 B.n646 B.n645 10.6151
R3405 B.n645 B.n642 10.6151
R3406 B.n642 B.n641 10.6151
R3407 B.n641 B.n638 10.6151
R3408 B.n638 B.n637 10.6151
R3409 B.n637 B.n634 10.6151
R3410 B.n634 B.n633 10.6151
R3411 B.n633 B.n630 10.6151
R3412 B.n630 B.n629 10.6151
R3413 B.n629 B.n627 10.6151
R3414 B.n890 B.n889 10.6151
R3415 B.n890 B.n545 10.6151
R3416 B.n900 B.n545 10.6151
R3417 B.n901 B.n900 10.6151
R3418 B.n902 B.n901 10.6151
R3419 B.n902 B.n537 10.6151
R3420 B.n913 B.n537 10.6151
R3421 B.n914 B.n913 10.6151
R3422 B.n915 B.n914 10.6151
R3423 B.n915 B.n530 10.6151
R3424 B.n925 B.n530 10.6151
R3425 B.n926 B.n925 10.6151
R3426 B.n927 B.n926 10.6151
R3427 B.n927 B.n522 10.6151
R3428 B.n937 B.n522 10.6151
R3429 B.n938 B.n937 10.6151
R3430 B.n939 B.n938 10.6151
R3431 B.n939 B.n514 10.6151
R3432 B.n949 B.n514 10.6151
R3433 B.n950 B.n949 10.6151
R3434 B.n951 B.n950 10.6151
R3435 B.n951 B.n506 10.6151
R3436 B.n961 B.n506 10.6151
R3437 B.n962 B.n961 10.6151
R3438 B.n963 B.n962 10.6151
R3439 B.n963 B.n498 10.6151
R3440 B.n973 B.n498 10.6151
R3441 B.n974 B.n973 10.6151
R3442 B.n975 B.n974 10.6151
R3443 B.n975 B.n490 10.6151
R3444 B.n985 B.n490 10.6151
R3445 B.n986 B.n985 10.6151
R3446 B.n987 B.n986 10.6151
R3447 B.n987 B.n482 10.6151
R3448 B.n997 B.n482 10.6151
R3449 B.n998 B.n997 10.6151
R3450 B.n999 B.n998 10.6151
R3451 B.n999 B.n474 10.6151
R3452 B.n1009 B.n474 10.6151
R3453 B.n1010 B.n1009 10.6151
R3454 B.n1011 B.n1010 10.6151
R3455 B.n1011 B.n466 10.6151
R3456 B.n1021 B.n466 10.6151
R3457 B.n1022 B.n1021 10.6151
R3458 B.n1023 B.n1022 10.6151
R3459 B.n1023 B.n458 10.6151
R3460 B.n1033 B.n458 10.6151
R3461 B.n1034 B.n1033 10.6151
R3462 B.n1035 B.n1034 10.6151
R3463 B.n1035 B.n450 10.6151
R3464 B.n1046 B.n450 10.6151
R3465 B.n1047 B.n1046 10.6151
R3466 B.n1048 B.n1047 10.6151
R3467 B.n1048 B.n443 10.6151
R3468 B.n1059 B.n443 10.6151
R3469 B.n1060 B.n1059 10.6151
R3470 B.n1061 B.n1060 10.6151
R3471 B.n1061 B.n0 10.6151
R3472 B.n1261 B.n1 10.6151
R3473 B.n1261 B.n1260 10.6151
R3474 B.n1260 B.n1259 10.6151
R3475 B.n1259 B.n10 10.6151
R3476 B.n1253 B.n10 10.6151
R3477 B.n1253 B.n1252 10.6151
R3478 B.n1252 B.n1251 10.6151
R3479 B.n1251 B.n16 10.6151
R3480 B.n1245 B.n16 10.6151
R3481 B.n1245 B.n1244 10.6151
R3482 B.n1244 B.n1243 10.6151
R3483 B.n1243 B.n24 10.6151
R3484 B.n1237 B.n24 10.6151
R3485 B.n1237 B.n1236 10.6151
R3486 B.n1236 B.n1235 10.6151
R3487 B.n1235 B.n31 10.6151
R3488 B.n1229 B.n31 10.6151
R3489 B.n1229 B.n1228 10.6151
R3490 B.n1228 B.n1227 10.6151
R3491 B.n1227 B.n38 10.6151
R3492 B.n1221 B.n38 10.6151
R3493 B.n1221 B.n1220 10.6151
R3494 B.n1220 B.n1219 10.6151
R3495 B.n1219 B.n45 10.6151
R3496 B.n1213 B.n45 10.6151
R3497 B.n1213 B.n1212 10.6151
R3498 B.n1212 B.n1211 10.6151
R3499 B.n1211 B.n52 10.6151
R3500 B.n1205 B.n52 10.6151
R3501 B.n1205 B.n1204 10.6151
R3502 B.n1204 B.n1203 10.6151
R3503 B.n1203 B.n59 10.6151
R3504 B.n1197 B.n59 10.6151
R3505 B.n1197 B.n1196 10.6151
R3506 B.n1196 B.n1195 10.6151
R3507 B.n1195 B.n66 10.6151
R3508 B.n1189 B.n66 10.6151
R3509 B.n1189 B.n1188 10.6151
R3510 B.n1188 B.n1187 10.6151
R3511 B.n1187 B.n73 10.6151
R3512 B.n1181 B.n73 10.6151
R3513 B.n1181 B.n1180 10.6151
R3514 B.n1180 B.n1179 10.6151
R3515 B.n1179 B.n80 10.6151
R3516 B.n1173 B.n80 10.6151
R3517 B.n1173 B.n1172 10.6151
R3518 B.n1172 B.n1171 10.6151
R3519 B.n1171 B.n87 10.6151
R3520 B.n1165 B.n87 10.6151
R3521 B.n1165 B.n1164 10.6151
R3522 B.n1164 B.n1163 10.6151
R3523 B.n1163 B.n93 10.6151
R3524 B.n1157 B.n93 10.6151
R3525 B.n1157 B.n1156 10.6151
R3526 B.n1156 B.n1155 10.6151
R3527 B.n1155 B.n101 10.6151
R3528 B.n1149 B.n101 10.6151
R3529 B.n1149 B.n1148 10.6151
R3530 B.n1043 B.t2 9.63152
R3531 B.n18 B.t1 9.63152
R3532 B.n298 B.n297 9.36635
R3533 B.n320 B.n319 9.36635
R3534 B.n769 B.n623 9.36635
R3535 B.n746 B.n626 9.36635
R3536 B.t7 B.n508 6.8798
R3537 B.n1192 B.t6 6.8798
R3538 B.n472 B.t0 4.12808
R3539 B.t4 B.n1232 4.12808
R3540 B.n1267 B.n0 2.81026
R3541 B.n1267 B.n1 2.81026
R3542 B.t5 B.n488 1.37636
R3543 B.t3 B.n50 1.37636
R3544 B.n299 B.n298 1.24928
R3545 B.n319 B.n318 1.24928
R3546 B.n766 B.n623 1.24928
R3547 B.n749 B.n626 1.24928
R3548 VP.n19 VP.t2 177.478
R3549 VP.n21 VP.n18 161.3
R3550 VP.n23 VP.n22 161.3
R3551 VP.n24 VP.n17 161.3
R3552 VP.n26 VP.n25 161.3
R3553 VP.n27 VP.n16 161.3
R3554 VP.n29 VP.n28 161.3
R3555 VP.n31 VP.n30 161.3
R3556 VP.n32 VP.n14 161.3
R3557 VP.n34 VP.n33 161.3
R3558 VP.n35 VP.n13 161.3
R3559 VP.n37 VP.n36 161.3
R3560 VP.n38 VP.n12 161.3
R3561 VP.n40 VP.n39 161.3
R3562 VP.n75 VP.n74 161.3
R3563 VP.n73 VP.n1 161.3
R3564 VP.n72 VP.n71 161.3
R3565 VP.n70 VP.n2 161.3
R3566 VP.n69 VP.n68 161.3
R3567 VP.n67 VP.n3 161.3
R3568 VP.n66 VP.n65 161.3
R3569 VP.n64 VP.n63 161.3
R3570 VP.n62 VP.n5 161.3
R3571 VP.n61 VP.n60 161.3
R3572 VP.n59 VP.n6 161.3
R3573 VP.n58 VP.n57 161.3
R3574 VP.n56 VP.n7 161.3
R3575 VP.n54 VP.n53 161.3
R3576 VP.n52 VP.n8 161.3
R3577 VP.n51 VP.n50 161.3
R3578 VP.n49 VP.n9 161.3
R3579 VP.n48 VP.n47 161.3
R3580 VP.n46 VP.n10 161.3
R3581 VP.n45 VP.n44 161.3
R3582 VP.n43 VP.t5 144.061
R3583 VP.n55 VP.t7 144.061
R3584 VP.n4 VP.t1 144.061
R3585 VP.n0 VP.t0 144.061
R3586 VP.n11 VP.t3 144.061
R3587 VP.n15 VP.t6 144.061
R3588 VP.n20 VP.t4 144.061
R3589 VP.n43 VP.n42 68.5364
R3590 VP.n76 VP.n0 68.5364
R3591 VP.n41 VP.n11 68.5364
R3592 VP.n42 VP.n41 58.6357
R3593 VP.n49 VP.n48 56.5193
R3594 VP.n61 VP.n6 56.5193
R3595 VP.n72 VP.n2 56.5193
R3596 VP.n37 VP.n13 56.5193
R3597 VP.n26 VP.n17 56.5193
R3598 VP.n20 VP.n19 50.4515
R3599 VP.n44 VP.n10 24.4675
R3600 VP.n48 VP.n10 24.4675
R3601 VP.n50 VP.n49 24.4675
R3602 VP.n50 VP.n8 24.4675
R3603 VP.n54 VP.n8 24.4675
R3604 VP.n57 VP.n56 24.4675
R3605 VP.n57 VP.n6 24.4675
R3606 VP.n62 VP.n61 24.4675
R3607 VP.n63 VP.n62 24.4675
R3608 VP.n67 VP.n66 24.4675
R3609 VP.n68 VP.n67 24.4675
R3610 VP.n68 VP.n2 24.4675
R3611 VP.n73 VP.n72 24.4675
R3612 VP.n74 VP.n73 24.4675
R3613 VP.n38 VP.n37 24.4675
R3614 VP.n39 VP.n38 24.4675
R3615 VP.n27 VP.n26 24.4675
R3616 VP.n28 VP.n27 24.4675
R3617 VP.n32 VP.n31 24.4675
R3618 VP.n33 VP.n32 24.4675
R3619 VP.n33 VP.n13 24.4675
R3620 VP.n22 VP.n21 24.4675
R3621 VP.n22 VP.n17 24.4675
R3622 VP.n56 VP.n55 23.4888
R3623 VP.n63 VP.n4 23.4888
R3624 VP.n28 VP.n15 23.4888
R3625 VP.n21 VP.n20 23.4888
R3626 VP.n44 VP.n43 21.5315
R3627 VP.n74 VP.n0 21.5315
R3628 VP.n39 VP.n11 21.5315
R3629 VP.n19 VP.n18 3.84097
R3630 VP.n55 VP.n54 0.97918
R3631 VP.n66 VP.n4 0.97918
R3632 VP.n31 VP.n15 0.97918
R3633 VP.n41 VP.n40 0.354971
R3634 VP.n45 VP.n42 0.354971
R3635 VP.n76 VP.n75 0.354971
R3636 VP VP.n76 0.26696
R3637 VP.n23 VP.n18 0.189894
R3638 VP.n24 VP.n23 0.189894
R3639 VP.n25 VP.n24 0.189894
R3640 VP.n25 VP.n16 0.189894
R3641 VP.n29 VP.n16 0.189894
R3642 VP.n30 VP.n29 0.189894
R3643 VP.n30 VP.n14 0.189894
R3644 VP.n34 VP.n14 0.189894
R3645 VP.n35 VP.n34 0.189894
R3646 VP.n36 VP.n35 0.189894
R3647 VP.n36 VP.n12 0.189894
R3648 VP.n40 VP.n12 0.189894
R3649 VP.n46 VP.n45 0.189894
R3650 VP.n47 VP.n46 0.189894
R3651 VP.n47 VP.n9 0.189894
R3652 VP.n51 VP.n9 0.189894
R3653 VP.n52 VP.n51 0.189894
R3654 VP.n53 VP.n52 0.189894
R3655 VP.n53 VP.n7 0.189894
R3656 VP.n58 VP.n7 0.189894
R3657 VP.n59 VP.n58 0.189894
R3658 VP.n60 VP.n59 0.189894
R3659 VP.n60 VP.n5 0.189894
R3660 VP.n64 VP.n5 0.189894
R3661 VP.n65 VP.n64 0.189894
R3662 VP.n65 VP.n3 0.189894
R3663 VP.n69 VP.n3 0.189894
R3664 VP.n70 VP.n69 0.189894
R3665 VP.n71 VP.n70 0.189894
R3666 VP.n71 VP.n1 0.189894
R3667 VP.n75 VP.n1 0.189894
R3668 VDD1 VDD1.n0 63.852
R3669 VDD1.n3 VDD1.n2 63.7374
R3670 VDD1.n3 VDD1.n1 63.7374
R3671 VDD1.n5 VDD1.n4 62.3013
R3672 VDD1.n5 VDD1.n3 53.85
R3673 VDD1 VDD1.n5 1.43369
R3674 VDD1.n4 VDD1.t1 1.05876
R3675 VDD1.n4 VDD1.t4 1.05876
R3676 VDD1.n0 VDD1.t5 1.05876
R3677 VDD1.n0 VDD1.t3 1.05876
R3678 VDD1.n2 VDD1.t6 1.05876
R3679 VDD1.n2 VDD1.t7 1.05876
R3680 VDD1.n1 VDD1.t2 1.05876
R3681 VDD1.n1 VDD1.t0 1.05876
C0 VP VTAIL 14.038401f
C1 VDD1 VDD2 2.05437f
C2 VDD1 VP 14.176901f
C3 VDD2 VP 0.576193f
C4 VN VTAIL 14.0243f
C5 VDD1 VN 0.15281f
C6 VDD2 VN 13.755099f
C7 VDD1 VTAIL 10.2922f
C8 VP VN 9.552509f
C9 VDD2 VTAIL 10.350201f
C10 VDD2 B 6.434165f
C11 VDD1 B 6.923973f
C12 VTAIL B 14.89656f
C13 VN B 18.08693f
C14 VP B 16.6275f
C15 VDD1.t5 B 0.392702f
C16 VDD1.t3 B 0.392702f
C17 VDD1.n0 B 3.60596f
C18 VDD1.t2 B 0.392702f
C19 VDD1.t0 B 0.392702f
C20 VDD1.n1 B 3.6047f
C21 VDD1.t6 B 0.392702f
C22 VDD1.t7 B 0.392702f
C23 VDD1.n2 B 3.6047f
C24 VDD1.n3 B 4.3051f
C25 VDD1.t1 B 0.392702f
C26 VDD1.t4 B 0.392702f
C27 VDD1.n4 B 3.59112f
C28 VDD1.n5 B 3.8947f
C29 VP.t0 B 3.03169f
C30 VP.n0 B 1.12544f
C31 VP.n1 B 0.018808f
C32 VP.n2 B 0.025359f
C33 VP.n3 B 0.018808f
C34 VP.t1 B 3.03169f
C35 VP.n4 B 1.0462f
C36 VP.n5 B 0.018808f
C37 VP.n6 B 0.027456f
C38 VP.n7 B 0.018808f
C39 VP.t7 B 3.03169f
C40 VP.n8 B 0.035053f
C41 VP.n9 B 0.018808f
C42 VP.n10 B 0.035053f
C43 VP.t3 B 3.03169f
C44 VP.n11 B 1.12544f
C45 VP.n12 B 0.018808f
C46 VP.n13 B 0.025359f
C47 VP.n14 B 0.018808f
C48 VP.t6 B 3.03169f
C49 VP.n15 B 1.0462f
C50 VP.n16 B 0.018808f
C51 VP.n17 B 0.027456f
C52 VP.n18 B 0.21436f
C53 VP.t4 B 3.03169f
C54 VP.t2 B 3.25429f
C55 VP.n19 B 1.07098f
C56 VP.n20 B 1.11633f
C57 VP.n21 B 0.03436f
C58 VP.n22 B 0.035053f
C59 VP.n23 B 0.018808f
C60 VP.n24 B 0.018808f
C61 VP.n25 B 0.018808f
C62 VP.n26 B 0.027456f
C63 VP.n27 B 0.035053f
C64 VP.n28 B 0.03436f
C65 VP.n29 B 0.018808f
C66 VP.n30 B 0.018808f
C67 VP.n31 B 0.018439f
C68 VP.n32 B 0.035053f
C69 VP.n33 B 0.035053f
C70 VP.n34 B 0.018808f
C71 VP.n35 B 0.018808f
C72 VP.n36 B 0.018808f
C73 VP.n37 B 0.029552f
C74 VP.n38 B 0.035053f
C75 VP.n39 B 0.032976f
C76 VP.n40 B 0.030355f
C77 VP.n41 B 1.32909f
C78 VP.n42 B 1.34062f
C79 VP.t5 B 3.03169f
C80 VP.n43 B 1.12544f
C81 VP.n44 B 0.032976f
C82 VP.n45 B 0.030355f
C83 VP.n46 B 0.018808f
C84 VP.n47 B 0.018808f
C85 VP.n48 B 0.029552f
C86 VP.n49 B 0.025359f
C87 VP.n50 B 0.035053f
C88 VP.n51 B 0.018808f
C89 VP.n52 B 0.018808f
C90 VP.n53 B 0.018808f
C91 VP.n54 B 0.018439f
C92 VP.n55 B 1.0462f
C93 VP.n56 B 0.03436f
C94 VP.n57 B 0.035053f
C95 VP.n58 B 0.018808f
C96 VP.n59 B 0.018808f
C97 VP.n60 B 0.018808f
C98 VP.n61 B 0.027456f
C99 VP.n62 B 0.035053f
C100 VP.n63 B 0.03436f
C101 VP.n64 B 0.018808f
C102 VP.n65 B 0.018808f
C103 VP.n66 B 0.018439f
C104 VP.n67 B 0.035053f
C105 VP.n68 B 0.035053f
C106 VP.n69 B 0.018808f
C107 VP.n70 B 0.018808f
C108 VP.n71 B 0.018808f
C109 VP.n72 B 0.029552f
C110 VP.n73 B 0.035053f
C111 VP.n74 B 0.032976f
C112 VP.n75 B 0.030355f
C113 VP.n76 B 0.038531f
C114 VTAIL.t11 B 0.276535f
C115 VTAIL.t12 B 0.276535f
C116 VTAIL.n0 B 2.47527f
C117 VTAIL.n1 B 0.36144f
C118 VTAIL.n2 B 0.010507f
C119 VTAIL.n3 B 0.023756f
C120 VTAIL.n4 B 0.010642f
C121 VTAIL.n5 B 0.018703f
C122 VTAIL.n6 B 0.01005f
C123 VTAIL.n7 B 0.023756f
C124 VTAIL.n8 B 0.010642f
C125 VTAIL.n9 B 0.018703f
C126 VTAIL.n10 B 0.01005f
C127 VTAIL.n11 B 0.023756f
C128 VTAIL.n12 B 0.010642f
C129 VTAIL.n13 B 0.018703f
C130 VTAIL.n14 B 0.01005f
C131 VTAIL.n15 B 0.023756f
C132 VTAIL.n16 B 0.010642f
C133 VTAIL.n17 B 0.018703f
C134 VTAIL.n18 B 0.01005f
C135 VTAIL.n19 B 0.023756f
C136 VTAIL.n20 B 0.010642f
C137 VTAIL.n21 B 0.018703f
C138 VTAIL.n22 B 0.01005f
C139 VTAIL.n23 B 0.023756f
C140 VTAIL.n24 B 0.010346f
C141 VTAIL.n25 B 0.018703f
C142 VTAIL.n26 B 0.010642f
C143 VTAIL.n27 B 0.023756f
C144 VTAIL.n28 B 0.010642f
C145 VTAIL.n29 B 0.018703f
C146 VTAIL.n30 B 0.01005f
C147 VTAIL.n31 B 0.023756f
C148 VTAIL.n32 B 0.010642f
C149 VTAIL.n33 B 1.50177f
C150 VTAIL.n34 B 0.01005f
C151 VTAIL.t9 B 0.040797f
C152 VTAIL.n35 B 0.183032f
C153 VTAIL.n36 B 0.016793f
C154 VTAIL.n37 B 0.017817f
C155 VTAIL.n38 B 0.023756f
C156 VTAIL.n39 B 0.010642f
C157 VTAIL.n40 B 0.01005f
C158 VTAIL.n41 B 0.018703f
C159 VTAIL.n42 B 0.018703f
C160 VTAIL.n43 B 0.01005f
C161 VTAIL.n44 B 0.010642f
C162 VTAIL.n45 B 0.023756f
C163 VTAIL.n46 B 0.023756f
C164 VTAIL.n47 B 0.010642f
C165 VTAIL.n48 B 0.01005f
C166 VTAIL.n49 B 0.018703f
C167 VTAIL.n50 B 0.018703f
C168 VTAIL.n51 B 0.01005f
C169 VTAIL.n52 B 0.01005f
C170 VTAIL.n53 B 0.010642f
C171 VTAIL.n54 B 0.023756f
C172 VTAIL.n55 B 0.023756f
C173 VTAIL.n56 B 0.023756f
C174 VTAIL.n57 B 0.010346f
C175 VTAIL.n58 B 0.01005f
C176 VTAIL.n59 B 0.018703f
C177 VTAIL.n60 B 0.018703f
C178 VTAIL.n61 B 0.01005f
C179 VTAIL.n62 B 0.010642f
C180 VTAIL.n63 B 0.023756f
C181 VTAIL.n64 B 0.023756f
C182 VTAIL.n65 B 0.010642f
C183 VTAIL.n66 B 0.01005f
C184 VTAIL.n67 B 0.018703f
C185 VTAIL.n68 B 0.018703f
C186 VTAIL.n69 B 0.01005f
C187 VTAIL.n70 B 0.010642f
C188 VTAIL.n71 B 0.023756f
C189 VTAIL.n72 B 0.023756f
C190 VTAIL.n73 B 0.010642f
C191 VTAIL.n74 B 0.01005f
C192 VTAIL.n75 B 0.018703f
C193 VTAIL.n76 B 0.018703f
C194 VTAIL.n77 B 0.01005f
C195 VTAIL.n78 B 0.010642f
C196 VTAIL.n79 B 0.023756f
C197 VTAIL.n80 B 0.023756f
C198 VTAIL.n81 B 0.010642f
C199 VTAIL.n82 B 0.01005f
C200 VTAIL.n83 B 0.018703f
C201 VTAIL.n84 B 0.018703f
C202 VTAIL.n85 B 0.01005f
C203 VTAIL.n86 B 0.010642f
C204 VTAIL.n87 B 0.023756f
C205 VTAIL.n88 B 0.023756f
C206 VTAIL.n89 B 0.010642f
C207 VTAIL.n90 B 0.01005f
C208 VTAIL.n91 B 0.018703f
C209 VTAIL.n92 B 0.018703f
C210 VTAIL.n93 B 0.01005f
C211 VTAIL.n94 B 0.010642f
C212 VTAIL.n95 B 0.023756f
C213 VTAIL.n96 B 0.023756f
C214 VTAIL.n97 B 0.010642f
C215 VTAIL.n98 B 0.01005f
C216 VTAIL.n99 B 0.018703f
C217 VTAIL.n100 B 0.046043f
C218 VTAIL.n101 B 0.01005f
C219 VTAIL.n102 B 0.010642f
C220 VTAIL.n103 B 0.046741f
C221 VTAIL.n104 B 0.038586f
C222 VTAIL.n105 B 0.22535f
C223 VTAIL.n106 B 0.010507f
C224 VTAIL.n107 B 0.023756f
C225 VTAIL.n108 B 0.010642f
C226 VTAIL.n109 B 0.018703f
C227 VTAIL.n110 B 0.01005f
C228 VTAIL.n111 B 0.023756f
C229 VTAIL.n112 B 0.010642f
C230 VTAIL.n113 B 0.018703f
C231 VTAIL.n114 B 0.01005f
C232 VTAIL.n115 B 0.023756f
C233 VTAIL.n116 B 0.010642f
C234 VTAIL.n117 B 0.018703f
C235 VTAIL.n118 B 0.01005f
C236 VTAIL.n119 B 0.023756f
C237 VTAIL.n120 B 0.010642f
C238 VTAIL.n121 B 0.018703f
C239 VTAIL.n122 B 0.01005f
C240 VTAIL.n123 B 0.023756f
C241 VTAIL.n124 B 0.010642f
C242 VTAIL.n125 B 0.018703f
C243 VTAIL.n126 B 0.01005f
C244 VTAIL.n127 B 0.023756f
C245 VTAIL.n128 B 0.010346f
C246 VTAIL.n129 B 0.018703f
C247 VTAIL.n130 B 0.010642f
C248 VTAIL.n131 B 0.023756f
C249 VTAIL.n132 B 0.010642f
C250 VTAIL.n133 B 0.018703f
C251 VTAIL.n134 B 0.01005f
C252 VTAIL.n135 B 0.023756f
C253 VTAIL.n136 B 0.010642f
C254 VTAIL.n137 B 1.50177f
C255 VTAIL.n138 B 0.01005f
C256 VTAIL.t2 B 0.040797f
C257 VTAIL.n139 B 0.183032f
C258 VTAIL.n140 B 0.016793f
C259 VTAIL.n141 B 0.017817f
C260 VTAIL.n142 B 0.023756f
C261 VTAIL.n143 B 0.010642f
C262 VTAIL.n144 B 0.01005f
C263 VTAIL.n145 B 0.018703f
C264 VTAIL.n146 B 0.018703f
C265 VTAIL.n147 B 0.01005f
C266 VTAIL.n148 B 0.010642f
C267 VTAIL.n149 B 0.023756f
C268 VTAIL.n150 B 0.023756f
C269 VTAIL.n151 B 0.010642f
C270 VTAIL.n152 B 0.01005f
C271 VTAIL.n153 B 0.018703f
C272 VTAIL.n154 B 0.018703f
C273 VTAIL.n155 B 0.01005f
C274 VTAIL.n156 B 0.01005f
C275 VTAIL.n157 B 0.010642f
C276 VTAIL.n158 B 0.023756f
C277 VTAIL.n159 B 0.023756f
C278 VTAIL.n160 B 0.023756f
C279 VTAIL.n161 B 0.010346f
C280 VTAIL.n162 B 0.01005f
C281 VTAIL.n163 B 0.018703f
C282 VTAIL.n164 B 0.018703f
C283 VTAIL.n165 B 0.01005f
C284 VTAIL.n166 B 0.010642f
C285 VTAIL.n167 B 0.023756f
C286 VTAIL.n168 B 0.023756f
C287 VTAIL.n169 B 0.010642f
C288 VTAIL.n170 B 0.01005f
C289 VTAIL.n171 B 0.018703f
C290 VTAIL.n172 B 0.018703f
C291 VTAIL.n173 B 0.01005f
C292 VTAIL.n174 B 0.010642f
C293 VTAIL.n175 B 0.023756f
C294 VTAIL.n176 B 0.023756f
C295 VTAIL.n177 B 0.010642f
C296 VTAIL.n178 B 0.01005f
C297 VTAIL.n179 B 0.018703f
C298 VTAIL.n180 B 0.018703f
C299 VTAIL.n181 B 0.01005f
C300 VTAIL.n182 B 0.010642f
C301 VTAIL.n183 B 0.023756f
C302 VTAIL.n184 B 0.023756f
C303 VTAIL.n185 B 0.010642f
C304 VTAIL.n186 B 0.01005f
C305 VTAIL.n187 B 0.018703f
C306 VTAIL.n188 B 0.018703f
C307 VTAIL.n189 B 0.01005f
C308 VTAIL.n190 B 0.010642f
C309 VTAIL.n191 B 0.023756f
C310 VTAIL.n192 B 0.023756f
C311 VTAIL.n193 B 0.010642f
C312 VTAIL.n194 B 0.01005f
C313 VTAIL.n195 B 0.018703f
C314 VTAIL.n196 B 0.018703f
C315 VTAIL.n197 B 0.01005f
C316 VTAIL.n198 B 0.010642f
C317 VTAIL.n199 B 0.023756f
C318 VTAIL.n200 B 0.023756f
C319 VTAIL.n201 B 0.010642f
C320 VTAIL.n202 B 0.01005f
C321 VTAIL.n203 B 0.018703f
C322 VTAIL.n204 B 0.046043f
C323 VTAIL.n205 B 0.01005f
C324 VTAIL.n206 B 0.010642f
C325 VTAIL.n207 B 0.046741f
C326 VTAIL.n208 B 0.038586f
C327 VTAIL.n209 B 0.22535f
C328 VTAIL.t5 B 0.276535f
C329 VTAIL.t0 B 0.276535f
C330 VTAIL.n210 B 2.47527f
C331 VTAIL.n211 B 0.537695f
C332 VTAIL.n212 B 0.010507f
C333 VTAIL.n213 B 0.023756f
C334 VTAIL.n214 B 0.010642f
C335 VTAIL.n215 B 0.018703f
C336 VTAIL.n216 B 0.01005f
C337 VTAIL.n217 B 0.023756f
C338 VTAIL.n218 B 0.010642f
C339 VTAIL.n219 B 0.018703f
C340 VTAIL.n220 B 0.01005f
C341 VTAIL.n221 B 0.023756f
C342 VTAIL.n222 B 0.010642f
C343 VTAIL.n223 B 0.018703f
C344 VTAIL.n224 B 0.01005f
C345 VTAIL.n225 B 0.023756f
C346 VTAIL.n226 B 0.010642f
C347 VTAIL.n227 B 0.018703f
C348 VTAIL.n228 B 0.01005f
C349 VTAIL.n229 B 0.023756f
C350 VTAIL.n230 B 0.010642f
C351 VTAIL.n231 B 0.018703f
C352 VTAIL.n232 B 0.01005f
C353 VTAIL.n233 B 0.023756f
C354 VTAIL.n234 B 0.010346f
C355 VTAIL.n235 B 0.018703f
C356 VTAIL.n236 B 0.010642f
C357 VTAIL.n237 B 0.023756f
C358 VTAIL.n238 B 0.010642f
C359 VTAIL.n239 B 0.018703f
C360 VTAIL.n240 B 0.01005f
C361 VTAIL.n241 B 0.023756f
C362 VTAIL.n242 B 0.010642f
C363 VTAIL.n243 B 1.50177f
C364 VTAIL.n244 B 0.01005f
C365 VTAIL.t7 B 0.040797f
C366 VTAIL.n245 B 0.183032f
C367 VTAIL.n246 B 0.016793f
C368 VTAIL.n247 B 0.017817f
C369 VTAIL.n248 B 0.023756f
C370 VTAIL.n249 B 0.010642f
C371 VTAIL.n250 B 0.01005f
C372 VTAIL.n251 B 0.018703f
C373 VTAIL.n252 B 0.018703f
C374 VTAIL.n253 B 0.01005f
C375 VTAIL.n254 B 0.010642f
C376 VTAIL.n255 B 0.023756f
C377 VTAIL.n256 B 0.023756f
C378 VTAIL.n257 B 0.010642f
C379 VTAIL.n258 B 0.01005f
C380 VTAIL.n259 B 0.018703f
C381 VTAIL.n260 B 0.018703f
C382 VTAIL.n261 B 0.01005f
C383 VTAIL.n262 B 0.01005f
C384 VTAIL.n263 B 0.010642f
C385 VTAIL.n264 B 0.023756f
C386 VTAIL.n265 B 0.023756f
C387 VTAIL.n266 B 0.023756f
C388 VTAIL.n267 B 0.010346f
C389 VTAIL.n268 B 0.01005f
C390 VTAIL.n269 B 0.018703f
C391 VTAIL.n270 B 0.018703f
C392 VTAIL.n271 B 0.01005f
C393 VTAIL.n272 B 0.010642f
C394 VTAIL.n273 B 0.023756f
C395 VTAIL.n274 B 0.023756f
C396 VTAIL.n275 B 0.010642f
C397 VTAIL.n276 B 0.01005f
C398 VTAIL.n277 B 0.018703f
C399 VTAIL.n278 B 0.018703f
C400 VTAIL.n279 B 0.01005f
C401 VTAIL.n280 B 0.010642f
C402 VTAIL.n281 B 0.023756f
C403 VTAIL.n282 B 0.023756f
C404 VTAIL.n283 B 0.010642f
C405 VTAIL.n284 B 0.01005f
C406 VTAIL.n285 B 0.018703f
C407 VTAIL.n286 B 0.018703f
C408 VTAIL.n287 B 0.01005f
C409 VTAIL.n288 B 0.010642f
C410 VTAIL.n289 B 0.023756f
C411 VTAIL.n290 B 0.023756f
C412 VTAIL.n291 B 0.010642f
C413 VTAIL.n292 B 0.01005f
C414 VTAIL.n293 B 0.018703f
C415 VTAIL.n294 B 0.018703f
C416 VTAIL.n295 B 0.01005f
C417 VTAIL.n296 B 0.010642f
C418 VTAIL.n297 B 0.023756f
C419 VTAIL.n298 B 0.023756f
C420 VTAIL.n299 B 0.010642f
C421 VTAIL.n300 B 0.01005f
C422 VTAIL.n301 B 0.018703f
C423 VTAIL.n302 B 0.018703f
C424 VTAIL.n303 B 0.01005f
C425 VTAIL.n304 B 0.010642f
C426 VTAIL.n305 B 0.023756f
C427 VTAIL.n306 B 0.023756f
C428 VTAIL.n307 B 0.010642f
C429 VTAIL.n308 B 0.01005f
C430 VTAIL.n309 B 0.018703f
C431 VTAIL.n310 B 0.046043f
C432 VTAIL.n311 B 0.01005f
C433 VTAIL.n312 B 0.010642f
C434 VTAIL.n313 B 0.046741f
C435 VTAIL.n314 B 0.038586f
C436 VTAIL.n315 B 1.60292f
C437 VTAIL.n316 B 0.010507f
C438 VTAIL.n317 B 0.023756f
C439 VTAIL.n318 B 0.010642f
C440 VTAIL.n319 B 0.018703f
C441 VTAIL.n320 B 0.01005f
C442 VTAIL.n321 B 0.023756f
C443 VTAIL.n322 B 0.010642f
C444 VTAIL.n323 B 0.018703f
C445 VTAIL.n324 B 0.01005f
C446 VTAIL.n325 B 0.023756f
C447 VTAIL.n326 B 0.010642f
C448 VTAIL.n327 B 0.018703f
C449 VTAIL.n328 B 0.01005f
C450 VTAIL.n329 B 0.023756f
C451 VTAIL.n330 B 0.010642f
C452 VTAIL.n331 B 0.018703f
C453 VTAIL.n332 B 0.01005f
C454 VTAIL.n333 B 0.023756f
C455 VTAIL.n334 B 0.010642f
C456 VTAIL.n335 B 0.018703f
C457 VTAIL.n336 B 0.01005f
C458 VTAIL.n337 B 0.023756f
C459 VTAIL.n338 B 0.010346f
C460 VTAIL.n339 B 0.018703f
C461 VTAIL.n340 B 0.010346f
C462 VTAIL.n341 B 0.01005f
C463 VTAIL.n342 B 0.023756f
C464 VTAIL.n343 B 0.023756f
C465 VTAIL.n344 B 0.010642f
C466 VTAIL.n345 B 0.018703f
C467 VTAIL.n346 B 0.01005f
C468 VTAIL.n347 B 0.023756f
C469 VTAIL.n348 B 0.010642f
C470 VTAIL.n349 B 1.50177f
C471 VTAIL.n350 B 0.01005f
C472 VTAIL.t15 B 0.040797f
C473 VTAIL.n351 B 0.183032f
C474 VTAIL.n352 B 0.016793f
C475 VTAIL.n353 B 0.017817f
C476 VTAIL.n354 B 0.023756f
C477 VTAIL.n355 B 0.010642f
C478 VTAIL.n356 B 0.01005f
C479 VTAIL.n357 B 0.018703f
C480 VTAIL.n358 B 0.018703f
C481 VTAIL.n359 B 0.01005f
C482 VTAIL.n360 B 0.010642f
C483 VTAIL.n361 B 0.023756f
C484 VTAIL.n362 B 0.023756f
C485 VTAIL.n363 B 0.010642f
C486 VTAIL.n364 B 0.01005f
C487 VTAIL.n365 B 0.018703f
C488 VTAIL.n366 B 0.018703f
C489 VTAIL.n367 B 0.01005f
C490 VTAIL.n368 B 0.010642f
C491 VTAIL.n369 B 0.023756f
C492 VTAIL.n370 B 0.023756f
C493 VTAIL.n371 B 0.010642f
C494 VTAIL.n372 B 0.01005f
C495 VTAIL.n373 B 0.018703f
C496 VTAIL.n374 B 0.018703f
C497 VTAIL.n375 B 0.01005f
C498 VTAIL.n376 B 0.010642f
C499 VTAIL.n377 B 0.023756f
C500 VTAIL.n378 B 0.023756f
C501 VTAIL.n379 B 0.010642f
C502 VTAIL.n380 B 0.01005f
C503 VTAIL.n381 B 0.018703f
C504 VTAIL.n382 B 0.018703f
C505 VTAIL.n383 B 0.01005f
C506 VTAIL.n384 B 0.010642f
C507 VTAIL.n385 B 0.023756f
C508 VTAIL.n386 B 0.023756f
C509 VTAIL.n387 B 0.010642f
C510 VTAIL.n388 B 0.01005f
C511 VTAIL.n389 B 0.018703f
C512 VTAIL.n390 B 0.018703f
C513 VTAIL.n391 B 0.01005f
C514 VTAIL.n392 B 0.010642f
C515 VTAIL.n393 B 0.023756f
C516 VTAIL.n394 B 0.023756f
C517 VTAIL.n395 B 0.010642f
C518 VTAIL.n396 B 0.01005f
C519 VTAIL.n397 B 0.018703f
C520 VTAIL.n398 B 0.018703f
C521 VTAIL.n399 B 0.01005f
C522 VTAIL.n400 B 0.010642f
C523 VTAIL.n401 B 0.023756f
C524 VTAIL.n402 B 0.023756f
C525 VTAIL.n403 B 0.010642f
C526 VTAIL.n404 B 0.01005f
C527 VTAIL.n405 B 0.018703f
C528 VTAIL.n406 B 0.018703f
C529 VTAIL.n407 B 0.01005f
C530 VTAIL.n408 B 0.010642f
C531 VTAIL.n409 B 0.023756f
C532 VTAIL.n410 B 0.023756f
C533 VTAIL.n411 B 0.010642f
C534 VTAIL.n412 B 0.01005f
C535 VTAIL.n413 B 0.018703f
C536 VTAIL.n414 B 0.046043f
C537 VTAIL.n415 B 0.01005f
C538 VTAIL.n416 B 0.010642f
C539 VTAIL.n417 B 0.046741f
C540 VTAIL.n418 B 0.038586f
C541 VTAIL.n419 B 1.60292f
C542 VTAIL.t8 B 0.276535f
C543 VTAIL.t14 B 0.276535f
C544 VTAIL.n420 B 2.47526f
C545 VTAIL.n421 B 0.537701f
C546 VTAIL.n422 B 0.010507f
C547 VTAIL.n423 B 0.023756f
C548 VTAIL.n424 B 0.010642f
C549 VTAIL.n425 B 0.018703f
C550 VTAIL.n426 B 0.01005f
C551 VTAIL.n427 B 0.023756f
C552 VTAIL.n428 B 0.010642f
C553 VTAIL.n429 B 0.018703f
C554 VTAIL.n430 B 0.01005f
C555 VTAIL.n431 B 0.023756f
C556 VTAIL.n432 B 0.010642f
C557 VTAIL.n433 B 0.018703f
C558 VTAIL.n434 B 0.01005f
C559 VTAIL.n435 B 0.023756f
C560 VTAIL.n436 B 0.010642f
C561 VTAIL.n437 B 0.018703f
C562 VTAIL.n438 B 0.01005f
C563 VTAIL.n439 B 0.023756f
C564 VTAIL.n440 B 0.010642f
C565 VTAIL.n441 B 0.018703f
C566 VTAIL.n442 B 0.01005f
C567 VTAIL.n443 B 0.023756f
C568 VTAIL.n444 B 0.010346f
C569 VTAIL.n445 B 0.018703f
C570 VTAIL.n446 B 0.010346f
C571 VTAIL.n447 B 0.01005f
C572 VTAIL.n448 B 0.023756f
C573 VTAIL.n449 B 0.023756f
C574 VTAIL.n450 B 0.010642f
C575 VTAIL.n451 B 0.018703f
C576 VTAIL.n452 B 0.01005f
C577 VTAIL.n453 B 0.023756f
C578 VTAIL.n454 B 0.010642f
C579 VTAIL.n455 B 1.50177f
C580 VTAIL.n456 B 0.01005f
C581 VTAIL.t10 B 0.040797f
C582 VTAIL.n457 B 0.183032f
C583 VTAIL.n458 B 0.016793f
C584 VTAIL.n459 B 0.017817f
C585 VTAIL.n460 B 0.023756f
C586 VTAIL.n461 B 0.010642f
C587 VTAIL.n462 B 0.01005f
C588 VTAIL.n463 B 0.018703f
C589 VTAIL.n464 B 0.018703f
C590 VTAIL.n465 B 0.01005f
C591 VTAIL.n466 B 0.010642f
C592 VTAIL.n467 B 0.023756f
C593 VTAIL.n468 B 0.023756f
C594 VTAIL.n469 B 0.010642f
C595 VTAIL.n470 B 0.01005f
C596 VTAIL.n471 B 0.018703f
C597 VTAIL.n472 B 0.018703f
C598 VTAIL.n473 B 0.01005f
C599 VTAIL.n474 B 0.010642f
C600 VTAIL.n475 B 0.023756f
C601 VTAIL.n476 B 0.023756f
C602 VTAIL.n477 B 0.010642f
C603 VTAIL.n478 B 0.01005f
C604 VTAIL.n479 B 0.018703f
C605 VTAIL.n480 B 0.018703f
C606 VTAIL.n481 B 0.01005f
C607 VTAIL.n482 B 0.010642f
C608 VTAIL.n483 B 0.023756f
C609 VTAIL.n484 B 0.023756f
C610 VTAIL.n485 B 0.010642f
C611 VTAIL.n486 B 0.01005f
C612 VTAIL.n487 B 0.018703f
C613 VTAIL.n488 B 0.018703f
C614 VTAIL.n489 B 0.01005f
C615 VTAIL.n490 B 0.010642f
C616 VTAIL.n491 B 0.023756f
C617 VTAIL.n492 B 0.023756f
C618 VTAIL.n493 B 0.010642f
C619 VTAIL.n494 B 0.01005f
C620 VTAIL.n495 B 0.018703f
C621 VTAIL.n496 B 0.018703f
C622 VTAIL.n497 B 0.01005f
C623 VTAIL.n498 B 0.010642f
C624 VTAIL.n499 B 0.023756f
C625 VTAIL.n500 B 0.023756f
C626 VTAIL.n501 B 0.010642f
C627 VTAIL.n502 B 0.01005f
C628 VTAIL.n503 B 0.018703f
C629 VTAIL.n504 B 0.018703f
C630 VTAIL.n505 B 0.01005f
C631 VTAIL.n506 B 0.010642f
C632 VTAIL.n507 B 0.023756f
C633 VTAIL.n508 B 0.023756f
C634 VTAIL.n509 B 0.010642f
C635 VTAIL.n510 B 0.01005f
C636 VTAIL.n511 B 0.018703f
C637 VTAIL.n512 B 0.018703f
C638 VTAIL.n513 B 0.01005f
C639 VTAIL.n514 B 0.010642f
C640 VTAIL.n515 B 0.023756f
C641 VTAIL.n516 B 0.023756f
C642 VTAIL.n517 B 0.010642f
C643 VTAIL.n518 B 0.01005f
C644 VTAIL.n519 B 0.018703f
C645 VTAIL.n520 B 0.046043f
C646 VTAIL.n521 B 0.01005f
C647 VTAIL.n522 B 0.010642f
C648 VTAIL.n523 B 0.046741f
C649 VTAIL.n524 B 0.038586f
C650 VTAIL.n525 B 0.22535f
C651 VTAIL.n526 B 0.010507f
C652 VTAIL.n527 B 0.023756f
C653 VTAIL.n528 B 0.010642f
C654 VTAIL.n529 B 0.018703f
C655 VTAIL.n530 B 0.01005f
C656 VTAIL.n531 B 0.023756f
C657 VTAIL.n532 B 0.010642f
C658 VTAIL.n533 B 0.018703f
C659 VTAIL.n534 B 0.01005f
C660 VTAIL.n535 B 0.023756f
C661 VTAIL.n536 B 0.010642f
C662 VTAIL.n537 B 0.018703f
C663 VTAIL.n538 B 0.01005f
C664 VTAIL.n539 B 0.023756f
C665 VTAIL.n540 B 0.010642f
C666 VTAIL.n541 B 0.018703f
C667 VTAIL.n542 B 0.01005f
C668 VTAIL.n543 B 0.023756f
C669 VTAIL.n544 B 0.010642f
C670 VTAIL.n545 B 0.018703f
C671 VTAIL.n546 B 0.01005f
C672 VTAIL.n547 B 0.023756f
C673 VTAIL.n548 B 0.010346f
C674 VTAIL.n549 B 0.018703f
C675 VTAIL.n550 B 0.010346f
C676 VTAIL.n551 B 0.01005f
C677 VTAIL.n552 B 0.023756f
C678 VTAIL.n553 B 0.023756f
C679 VTAIL.n554 B 0.010642f
C680 VTAIL.n555 B 0.018703f
C681 VTAIL.n556 B 0.01005f
C682 VTAIL.n557 B 0.023756f
C683 VTAIL.n558 B 0.010642f
C684 VTAIL.n559 B 1.50177f
C685 VTAIL.n560 B 0.01005f
C686 VTAIL.t1 B 0.040797f
C687 VTAIL.n561 B 0.183032f
C688 VTAIL.n562 B 0.016793f
C689 VTAIL.n563 B 0.017817f
C690 VTAIL.n564 B 0.023756f
C691 VTAIL.n565 B 0.010642f
C692 VTAIL.n566 B 0.01005f
C693 VTAIL.n567 B 0.018703f
C694 VTAIL.n568 B 0.018703f
C695 VTAIL.n569 B 0.01005f
C696 VTAIL.n570 B 0.010642f
C697 VTAIL.n571 B 0.023756f
C698 VTAIL.n572 B 0.023756f
C699 VTAIL.n573 B 0.010642f
C700 VTAIL.n574 B 0.01005f
C701 VTAIL.n575 B 0.018703f
C702 VTAIL.n576 B 0.018703f
C703 VTAIL.n577 B 0.01005f
C704 VTAIL.n578 B 0.010642f
C705 VTAIL.n579 B 0.023756f
C706 VTAIL.n580 B 0.023756f
C707 VTAIL.n581 B 0.010642f
C708 VTAIL.n582 B 0.01005f
C709 VTAIL.n583 B 0.018703f
C710 VTAIL.n584 B 0.018703f
C711 VTAIL.n585 B 0.01005f
C712 VTAIL.n586 B 0.010642f
C713 VTAIL.n587 B 0.023756f
C714 VTAIL.n588 B 0.023756f
C715 VTAIL.n589 B 0.010642f
C716 VTAIL.n590 B 0.01005f
C717 VTAIL.n591 B 0.018703f
C718 VTAIL.n592 B 0.018703f
C719 VTAIL.n593 B 0.01005f
C720 VTAIL.n594 B 0.010642f
C721 VTAIL.n595 B 0.023756f
C722 VTAIL.n596 B 0.023756f
C723 VTAIL.n597 B 0.010642f
C724 VTAIL.n598 B 0.01005f
C725 VTAIL.n599 B 0.018703f
C726 VTAIL.n600 B 0.018703f
C727 VTAIL.n601 B 0.01005f
C728 VTAIL.n602 B 0.010642f
C729 VTAIL.n603 B 0.023756f
C730 VTAIL.n604 B 0.023756f
C731 VTAIL.n605 B 0.010642f
C732 VTAIL.n606 B 0.01005f
C733 VTAIL.n607 B 0.018703f
C734 VTAIL.n608 B 0.018703f
C735 VTAIL.n609 B 0.01005f
C736 VTAIL.n610 B 0.010642f
C737 VTAIL.n611 B 0.023756f
C738 VTAIL.n612 B 0.023756f
C739 VTAIL.n613 B 0.010642f
C740 VTAIL.n614 B 0.01005f
C741 VTAIL.n615 B 0.018703f
C742 VTAIL.n616 B 0.018703f
C743 VTAIL.n617 B 0.01005f
C744 VTAIL.n618 B 0.010642f
C745 VTAIL.n619 B 0.023756f
C746 VTAIL.n620 B 0.023756f
C747 VTAIL.n621 B 0.010642f
C748 VTAIL.n622 B 0.01005f
C749 VTAIL.n623 B 0.018703f
C750 VTAIL.n624 B 0.046043f
C751 VTAIL.n625 B 0.01005f
C752 VTAIL.n626 B 0.010642f
C753 VTAIL.n627 B 0.046741f
C754 VTAIL.n628 B 0.038586f
C755 VTAIL.n629 B 0.22535f
C756 VTAIL.t4 B 0.276535f
C757 VTAIL.t3 B 0.276535f
C758 VTAIL.n630 B 2.47526f
C759 VTAIL.n631 B 0.537701f
C760 VTAIL.n632 B 0.010507f
C761 VTAIL.n633 B 0.023756f
C762 VTAIL.n634 B 0.010642f
C763 VTAIL.n635 B 0.018703f
C764 VTAIL.n636 B 0.01005f
C765 VTAIL.n637 B 0.023756f
C766 VTAIL.n638 B 0.010642f
C767 VTAIL.n639 B 0.018703f
C768 VTAIL.n640 B 0.01005f
C769 VTAIL.n641 B 0.023756f
C770 VTAIL.n642 B 0.010642f
C771 VTAIL.n643 B 0.018703f
C772 VTAIL.n644 B 0.01005f
C773 VTAIL.n645 B 0.023756f
C774 VTAIL.n646 B 0.010642f
C775 VTAIL.n647 B 0.018703f
C776 VTAIL.n648 B 0.01005f
C777 VTAIL.n649 B 0.023756f
C778 VTAIL.n650 B 0.010642f
C779 VTAIL.n651 B 0.018703f
C780 VTAIL.n652 B 0.01005f
C781 VTAIL.n653 B 0.023756f
C782 VTAIL.n654 B 0.010346f
C783 VTAIL.n655 B 0.018703f
C784 VTAIL.n656 B 0.010346f
C785 VTAIL.n657 B 0.01005f
C786 VTAIL.n658 B 0.023756f
C787 VTAIL.n659 B 0.023756f
C788 VTAIL.n660 B 0.010642f
C789 VTAIL.n661 B 0.018703f
C790 VTAIL.n662 B 0.01005f
C791 VTAIL.n663 B 0.023756f
C792 VTAIL.n664 B 0.010642f
C793 VTAIL.n665 B 1.50177f
C794 VTAIL.n666 B 0.01005f
C795 VTAIL.t6 B 0.040797f
C796 VTAIL.n667 B 0.183032f
C797 VTAIL.n668 B 0.016793f
C798 VTAIL.n669 B 0.017817f
C799 VTAIL.n670 B 0.023756f
C800 VTAIL.n671 B 0.010642f
C801 VTAIL.n672 B 0.01005f
C802 VTAIL.n673 B 0.018703f
C803 VTAIL.n674 B 0.018703f
C804 VTAIL.n675 B 0.01005f
C805 VTAIL.n676 B 0.010642f
C806 VTAIL.n677 B 0.023756f
C807 VTAIL.n678 B 0.023756f
C808 VTAIL.n679 B 0.010642f
C809 VTAIL.n680 B 0.01005f
C810 VTAIL.n681 B 0.018703f
C811 VTAIL.n682 B 0.018703f
C812 VTAIL.n683 B 0.01005f
C813 VTAIL.n684 B 0.010642f
C814 VTAIL.n685 B 0.023756f
C815 VTAIL.n686 B 0.023756f
C816 VTAIL.n687 B 0.010642f
C817 VTAIL.n688 B 0.01005f
C818 VTAIL.n689 B 0.018703f
C819 VTAIL.n690 B 0.018703f
C820 VTAIL.n691 B 0.01005f
C821 VTAIL.n692 B 0.010642f
C822 VTAIL.n693 B 0.023756f
C823 VTAIL.n694 B 0.023756f
C824 VTAIL.n695 B 0.010642f
C825 VTAIL.n696 B 0.01005f
C826 VTAIL.n697 B 0.018703f
C827 VTAIL.n698 B 0.018703f
C828 VTAIL.n699 B 0.01005f
C829 VTAIL.n700 B 0.010642f
C830 VTAIL.n701 B 0.023756f
C831 VTAIL.n702 B 0.023756f
C832 VTAIL.n703 B 0.010642f
C833 VTAIL.n704 B 0.01005f
C834 VTAIL.n705 B 0.018703f
C835 VTAIL.n706 B 0.018703f
C836 VTAIL.n707 B 0.01005f
C837 VTAIL.n708 B 0.010642f
C838 VTAIL.n709 B 0.023756f
C839 VTAIL.n710 B 0.023756f
C840 VTAIL.n711 B 0.010642f
C841 VTAIL.n712 B 0.01005f
C842 VTAIL.n713 B 0.018703f
C843 VTAIL.n714 B 0.018703f
C844 VTAIL.n715 B 0.01005f
C845 VTAIL.n716 B 0.010642f
C846 VTAIL.n717 B 0.023756f
C847 VTAIL.n718 B 0.023756f
C848 VTAIL.n719 B 0.010642f
C849 VTAIL.n720 B 0.01005f
C850 VTAIL.n721 B 0.018703f
C851 VTAIL.n722 B 0.018703f
C852 VTAIL.n723 B 0.01005f
C853 VTAIL.n724 B 0.010642f
C854 VTAIL.n725 B 0.023756f
C855 VTAIL.n726 B 0.023756f
C856 VTAIL.n727 B 0.010642f
C857 VTAIL.n728 B 0.01005f
C858 VTAIL.n729 B 0.018703f
C859 VTAIL.n730 B 0.046043f
C860 VTAIL.n731 B 0.01005f
C861 VTAIL.n732 B 0.010642f
C862 VTAIL.n733 B 0.046741f
C863 VTAIL.n734 B 0.038586f
C864 VTAIL.n735 B 1.60292f
C865 VTAIL.n736 B 0.010507f
C866 VTAIL.n737 B 0.023756f
C867 VTAIL.n738 B 0.010642f
C868 VTAIL.n739 B 0.018703f
C869 VTAIL.n740 B 0.01005f
C870 VTAIL.n741 B 0.023756f
C871 VTAIL.n742 B 0.010642f
C872 VTAIL.n743 B 0.018703f
C873 VTAIL.n744 B 0.01005f
C874 VTAIL.n745 B 0.023756f
C875 VTAIL.n746 B 0.010642f
C876 VTAIL.n747 B 0.018703f
C877 VTAIL.n748 B 0.01005f
C878 VTAIL.n749 B 0.023756f
C879 VTAIL.n750 B 0.010642f
C880 VTAIL.n751 B 0.018703f
C881 VTAIL.n752 B 0.01005f
C882 VTAIL.n753 B 0.023756f
C883 VTAIL.n754 B 0.010642f
C884 VTAIL.n755 B 0.018703f
C885 VTAIL.n756 B 0.01005f
C886 VTAIL.n757 B 0.023756f
C887 VTAIL.n758 B 0.010346f
C888 VTAIL.n759 B 0.018703f
C889 VTAIL.n760 B 0.010642f
C890 VTAIL.n761 B 0.023756f
C891 VTAIL.n762 B 0.010642f
C892 VTAIL.n763 B 0.018703f
C893 VTAIL.n764 B 0.01005f
C894 VTAIL.n765 B 0.023756f
C895 VTAIL.n766 B 0.010642f
C896 VTAIL.n767 B 1.50177f
C897 VTAIL.n768 B 0.01005f
C898 VTAIL.t13 B 0.040797f
C899 VTAIL.n769 B 0.183032f
C900 VTAIL.n770 B 0.016793f
C901 VTAIL.n771 B 0.017817f
C902 VTAIL.n772 B 0.023756f
C903 VTAIL.n773 B 0.010642f
C904 VTAIL.n774 B 0.01005f
C905 VTAIL.n775 B 0.018703f
C906 VTAIL.n776 B 0.018703f
C907 VTAIL.n777 B 0.01005f
C908 VTAIL.n778 B 0.010642f
C909 VTAIL.n779 B 0.023756f
C910 VTAIL.n780 B 0.023756f
C911 VTAIL.n781 B 0.010642f
C912 VTAIL.n782 B 0.01005f
C913 VTAIL.n783 B 0.018703f
C914 VTAIL.n784 B 0.018703f
C915 VTAIL.n785 B 0.01005f
C916 VTAIL.n786 B 0.01005f
C917 VTAIL.n787 B 0.010642f
C918 VTAIL.n788 B 0.023756f
C919 VTAIL.n789 B 0.023756f
C920 VTAIL.n790 B 0.023756f
C921 VTAIL.n791 B 0.010346f
C922 VTAIL.n792 B 0.01005f
C923 VTAIL.n793 B 0.018703f
C924 VTAIL.n794 B 0.018703f
C925 VTAIL.n795 B 0.01005f
C926 VTAIL.n796 B 0.010642f
C927 VTAIL.n797 B 0.023756f
C928 VTAIL.n798 B 0.023756f
C929 VTAIL.n799 B 0.010642f
C930 VTAIL.n800 B 0.01005f
C931 VTAIL.n801 B 0.018703f
C932 VTAIL.n802 B 0.018703f
C933 VTAIL.n803 B 0.01005f
C934 VTAIL.n804 B 0.010642f
C935 VTAIL.n805 B 0.023756f
C936 VTAIL.n806 B 0.023756f
C937 VTAIL.n807 B 0.010642f
C938 VTAIL.n808 B 0.01005f
C939 VTAIL.n809 B 0.018703f
C940 VTAIL.n810 B 0.018703f
C941 VTAIL.n811 B 0.01005f
C942 VTAIL.n812 B 0.010642f
C943 VTAIL.n813 B 0.023756f
C944 VTAIL.n814 B 0.023756f
C945 VTAIL.n815 B 0.010642f
C946 VTAIL.n816 B 0.01005f
C947 VTAIL.n817 B 0.018703f
C948 VTAIL.n818 B 0.018703f
C949 VTAIL.n819 B 0.01005f
C950 VTAIL.n820 B 0.010642f
C951 VTAIL.n821 B 0.023756f
C952 VTAIL.n822 B 0.023756f
C953 VTAIL.n823 B 0.010642f
C954 VTAIL.n824 B 0.01005f
C955 VTAIL.n825 B 0.018703f
C956 VTAIL.n826 B 0.018703f
C957 VTAIL.n827 B 0.01005f
C958 VTAIL.n828 B 0.010642f
C959 VTAIL.n829 B 0.023756f
C960 VTAIL.n830 B 0.023756f
C961 VTAIL.n831 B 0.010642f
C962 VTAIL.n832 B 0.01005f
C963 VTAIL.n833 B 0.018703f
C964 VTAIL.n834 B 0.046043f
C965 VTAIL.n835 B 0.01005f
C966 VTAIL.n836 B 0.010642f
C967 VTAIL.n837 B 0.046741f
C968 VTAIL.n838 B 0.038586f
C969 VTAIL.n839 B 1.59941f
C970 VDD2.t3 B 0.38971f
C971 VDD2.t1 B 0.38971f
C972 VDD2.n0 B 3.57724f
C973 VDD2.t4 B 0.38971f
C974 VDD2.t5 B 0.38971f
C975 VDD2.n1 B 3.57724f
C976 VDD2.n2 B 4.21798f
C977 VDD2.t7 B 0.38971f
C978 VDD2.t2 B 0.38971f
C979 VDD2.n3 B 3.56376f
C980 VDD2.n4 B 3.83188f
C981 VDD2.t6 B 0.38971f
C982 VDD2.t0 B 0.38971f
C983 VDD2.n5 B 3.57719f
C984 VN.t2 B 2.99752f
C985 VN.n0 B 1.11275f
C986 VN.n1 B 0.018596f
C987 VN.n2 B 0.025074f
C988 VN.n3 B 0.018596f
C989 VN.t3 B 2.99752f
C990 VN.n4 B 1.03441f
C991 VN.n5 B 0.018596f
C992 VN.n6 B 0.027146f
C993 VN.n7 B 0.211944f
C994 VN.t4 B 2.99752f
C995 VN.t6 B 3.2176f
C996 VN.n8 B 1.05891f
C997 VN.n9 B 1.10374f
C998 VN.n10 B 0.033973f
C999 VN.n11 B 0.034658f
C1000 VN.n12 B 0.018596f
C1001 VN.n13 B 0.018596f
C1002 VN.n14 B 0.018596f
C1003 VN.n15 B 0.027146f
C1004 VN.n16 B 0.034658f
C1005 VN.n17 B 0.033973f
C1006 VN.n18 B 0.018596f
C1007 VN.n19 B 0.018596f
C1008 VN.n20 B 0.018231f
C1009 VN.n21 B 0.034658f
C1010 VN.n22 B 0.034658f
C1011 VN.n23 B 0.018596f
C1012 VN.n24 B 0.018596f
C1013 VN.n25 B 0.018596f
C1014 VN.n26 B 0.029219f
C1015 VN.n27 B 0.034658f
C1016 VN.n28 B 0.032604f
C1017 VN.n29 B 0.030013f
C1018 VN.n30 B 0.038096f
C1019 VN.t0 B 2.99752f
C1020 VN.n31 B 1.11275f
C1021 VN.n32 B 0.018596f
C1022 VN.n33 B 0.025074f
C1023 VN.n34 B 0.018596f
C1024 VN.t7 B 2.99752f
C1025 VN.n35 B 1.03441f
C1026 VN.n36 B 0.018596f
C1027 VN.n37 B 0.027146f
C1028 VN.n38 B 0.211944f
C1029 VN.t1 B 2.99752f
C1030 VN.t5 B 3.2176f
C1031 VN.n39 B 1.05891f
C1032 VN.n40 B 1.10374f
C1033 VN.n41 B 0.033973f
C1034 VN.n42 B 0.034658f
C1035 VN.n43 B 0.018596f
C1036 VN.n44 B 0.018596f
C1037 VN.n45 B 0.018596f
C1038 VN.n46 B 0.027146f
C1039 VN.n47 B 0.034658f
C1040 VN.n48 B 0.033973f
C1041 VN.n49 B 0.018596f
C1042 VN.n50 B 0.018596f
C1043 VN.n51 B 0.018231f
C1044 VN.n52 B 0.034658f
C1045 VN.n53 B 0.034658f
C1046 VN.n54 B 0.018596f
C1047 VN.n55 B 0.018596f
C1048 VN.n56 B 0.018596f
C1049 VN.n57 B 0.029219f
C1050 VN.n58 B 0.034658f
C1051 VN.n59 B 0.032604f
C1052 VN.n60 B 0.030013f
C1053 VN.n61 B 1.32133f
.ends

