* NGSPICE file created from diff_pair_sample_1631.ext - technology: sky130A

.subckt diff_pair_sample_1631 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t7 VN.t0 VDD2.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=6.6456 pd=34.86 as=2.8116 ps=17.37 w=17.04 l=2.85
X1 VTAIL.t6 VN.t1 VDD2.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=6.6456 pd=34.86 as=2.8116 ps=17.37 w=17.04 l=2.85
X2 B.t17 B.t15 B.t16 B.t12 sky130_fd_pr__nfet_01v8 ad=6.6456 pd=34.86 as=0 ps=0 w=17.04 l=2.85
X3 VTAIL.t3 VP.t0 VDD1.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=6.6456 pd=34.86 as=2.8116 ps=17.37 w=17.04 l=2.85
X4 B.t14 B.t11 B.t13 B.t12 sky130_fd_pr__nfet_01v8 ad=6.6456 pd=34.86 as=0 ps=0 w=17.04 l=2.85
X5 VTAIL.t2 VP.t1 VDD1.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=6.6456 pd=34.86 as=2.8116 ps=17.37 w=17.04 l=2.85
X6 VDD1.t1 VP.t2 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=2.8116 pd=17.37 as=6.6456 ps=34.86 w=17.04 l=2.85
X7 VDD2.t1 VN.t2 VTAIL.t5 B.t0 sky130_fd_pr__nfet_01v8 ad=2.8116 pd=17.37 as=6.6456 ps=34.86 w=17.04 l=2.85
X8 B.t10 B.t8 B.t9 B.t5 sky130_fd_pr__nfet_01v8 ad=6.6456 pd=34.86 as=0 ps=0 w=17.04 l=2.85
X9 B.t7 B.t4 B.t6 B.t5 sky130_fd_pr__nfet_01v8 ad=6.6456 pd=34.86 as=0 ps=0 w=17.04 l=2.85
X10 VDD1.t0 VP.t3 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=2.8116 pd=17.37 as=6.6456 ps=34.86 w=17.04 l=2.85
X11 VDD2.t0 VN.t3 VTAIL.t4 B.t1 sky130_fd_pr__nfet_01v8 ad=2.8116 pd=17.37 as=6.6456 ps=34.86 w=17.04 l=2.85
R0 VN.n0 VN.t0 179.571
R1 VN.n1 VN.t2 179.571
R2 VN.n0 VN.t3 178.672
R3 VN.n1 VN.t1 178.672
R4 VN VN.n1 54.6105
R5 VN VN.n0 3.4249
R6 VDD2.n2 VDD2.n0 105.004
R7 VDD2.n2 VDD2.n1 58.3746
R8 VDD2.n1 VDD2.t2 1.16247
R9 VDD2.n1 VDD2.t1 1.16247
R10 VDD2.n0 VDD2.t3 1.16247
R11 VDD2.n0 VDD2.t0 1.16247
R12 VDD2 VDD2.n2 0.0586897
R13 VTAIL.n5 VTAIL.t3 42.8579
R14 VTAIL.n4 VTAIL.t5 42.8579
R15 VTAIL.n3 VTAIL.t6 42.8579
R16 VTAIL.n7 VTAIL.t4 42.8578
R17 VTAIL.n0 VTAIL.t7 42.8578
R18 VTAIL.n1 VTAIL.t0 42.8578
R19 VTAIL.n2 VTAIL.t2 42.8578
R20 VTAIL.n6 VTAIL.t1 42.8578
R21 VTAIL.n7 VTAIL.n6 29.7979
R22 VTAIL.n3 VTAIL.n2 29.7979
R23 VTAIL.n4 VTAIL.n3 2.74188
R24 VTAIL.n6 VTAIL.n5 2.74188
R25 VTAIL.n2 VTAIL.n1 2.74188
R26 VTAIL VTAIL.n0 1.42938
R27 VTAIL VTAIL.n7 1.313
R28 VTAIL.n5 VTAIL.n4 0.470328
R29 VTAIL.n1 VTAIL.n0 0.470328
R30 B.n910 B.n909 585
R31 B.n374 B.n129 585
R32 B.n373 B.n372 585
R33 B.n371 B.n370 585
R34 B.n369 B.n368 585
R35 B.n367 B.n366 585
R36 B.n365 B.n364 585
R37 B.n363 B.n362 585
R38 B.n361 B.n360 585
R39 B.n359 B.n358 585
R40 B.n357 B.n356 585
R41 B.n355 B.n354 585
R42 B.n353 B.n352 585
R43 B.n351 B.n350 585
R44 B.n349 B.n348 585
R45 B.n347 B.n346 585
R46 B.n345 B.n344 585
R47 B.n343 B.n342 585
R48 B.n341 B.n340 585
R49 B.n339 B.n338 585
R50 B.n337 B.n336 585
R51 B.n335 B.n334 585
R52 B.n333 B.n332 585
R53 B.n331 B.n330 585
R54 B.n329 B.n328 585
R55 B.n327 B.n326 585
R56 B.n325 B.n324 585
R57 B.n323 B.n322 585
R58 B.n321 B.n320 585
R59 B.n319 B.n318 585
R60 B.n317 B.n316 585
R61 B.n315 B.n314 585
R62 B.n313 B.n312 585
R63 B.n311 B.n310 585
R64 B.n309 B.n308 585
R65 B.n307 B.n306 585
R66 B.n305 B.n304 585
R67 B.n303 B.n302 585
R68 B.n301 B.n300 585
R69 B.n299 B.n298 585
R70 B.n297 B.n296 585
R71 B.n295 B.n294 585
R72 B.n293 B.n292 585
R73 B.n291 B.n290 585
R74 B.n289 B.n288 585
R75 B.n287 B.n286 585
R76 B.n285 B.n284 585
R77 B.n283 B.n282 585
R78 B.n281 B.n280 585
R79 B.n279 B.n278 585
R80 B.n277 B.n276 585
R81 B.n275 B.n274 585
R82 B.n273 B.n272 585
R83 B.n271 B.n270 585
R84 B.n269 B.n268 585
R85 B.n267 B.n266 585
R86 B.n265 B.n264 585
R87 B.n263 B.n262 585
R88 B.n261 B.n260 585
R89 B.n259 B.n258 585
R90 B.n257 B.n256 585
R91 B.n255 B.n254 585
R92 B.n253 B.n252 585
R93 B.n251 B.n250 585
R94 B.n249 B.n248 585
R95 B.n247 B.n246 585
R96 B.n245 B.n244 585
R97 B.n243 B.n242 585
R98 B.n241 B.n240 585
R99 B.n239 B.n238 585
R100 B.n237 B.n236 585
R101 B.n235 B.n234 585
R102 B.n233 B.n232 585
R103 B.n231 B.n230 585
R104 B.n229 B.n228 585
R105 B.n227 B.n226 585
R106 B.n225 B.n224 585
R107 B.n223 B.n222 585
R108 B.n221 B.n220 585
R109 B.n219 B.n218 585
R110 B.n217 B.n216 585
R111 B.n215 B.n214 585
R112 B.n213 B.n212 585
R113 B.n211 B.n210 585
R114 B.n209 B.n208 585
R115 B.n207 B.n206 585
R116 B.n205 B.n204 585
R117 B.n203 B.n202 585
R118 B.n201 B.n200 585
R119 B.n199 B.n198 585
R120 B.n197 B.n196 585
R121 B.n195 B.n194 585
R122 B.n193 B.n192 585
R123 B.n191 B.n190 585
R124 B.n189 B.n188 585
R125 B.n187 B.n186 585
R126 B.n185 B.n184 585
R127 B.n183 B.n182 585
R128 B.n181 B.n180 585
R129 B.n179 B.n178 585
R130 B.n177 B.n176 585
R131 B.n175 B.n174 585
R132 B.n173 B.n172 585
R133 B.n171 B.n170 585
R134 B.n169 B.n168 585
R135 B.n167 B.n166 585
R136 B.n165 B.n164 585
R137 B.n163 B.n162 585
R138 B.n161 B.n160 585
R139 B.n159 B.n158 585
R140 B.n157 B.n156 585
R141 B.n155 B.n154 585
R142 B.n153 B.n152 585
R143 B.n151 B.n150 585
R144 B.n149 B.n148 585
R145 B.n147 B.n146 585
R146 B.n145 B.n144 585
R147 B.n143 B.n142 585
R148 B.n141 B.n140 585
R149 B.n139 B.n138 585
R150 B.n137 B.n136 585
R151 B.n67 B.n66 585
R152 B.n908 B.n68 585
R153 B.n913 B.n68 585
R154 B.n907 B.n906 585
R155 B.n906 B.n64 585
R156 B.n905 B.n63 585
R157 B.n919 B.n63 585
R158 B.n904 B.n62 585
R159 B.n920 B.n62 585
R160 B.n903 B.n61 585
R161 B.n921 B.n61 585
R162 B.n902 B.n901 585
R163 B.n901 B.n57 585
R164 B.n900 B.n56 585
R165 B.n927 B.n56 585
R166 B.n899 B.n55 585
R167 B.n928 B.n55 585
R168 B.n898 B.n54 585
R169 B.n929 B.n54 585
R170 B.n897 B.n896 585
R171 B.n896 B.n50 585
R172 B.n895 B.n49 585
R173 B.n935 B.n49 585
R174 B.n894 B.n48 585
R175 B.n936 B.n48 585
R176 B.n893 B.n47 585
R177 B.n937 B.n47 585
R178 B.n892 B.n891 585
R179 B.n891 B.n43 585
R180 B.n890 B.n42 585
R181 B.n943 B.n42 585
R182 B.n889 B.n41 585
R183 B.n944 B.n41 585
R184 B.n888 B.n40 585
R185 B.n945 B.n40 585
R186 B.n887 B.n886 585
R187 B.n886 B.n36 585
R188 B.n885 B.n35 585
R189 B.n951 B.n35 585
R190 B.n884 B.n34 585
R191 B.n952 B.n34 585
R192 B.n883 B.n33 585
R193 B.n953 B.n33 585
R194 B.n882 B.n881 585
R195 B.n881 B.n29 585
R196 B.n880 B.n28 585
R197 B.n959 B.n28 585
R198 B.n879 B.n27 585
R199 B.n960 B.n27 585
R200 B.n878 B.n26 585
R201 B.n961 B.n26 585
R202 B.n877 B.n876 585
R203 B.n876 B.n22 585
R204 B.n875 B.n21 585
R205 B.n967 B.n21 585
R206 B.n874 B.n20 585
R207 B.n968 B.n20 585
R208 B.n873 B.n19 585
R209 B.n969 B.n19 585
R210 B.n872 B.n871 585
R211 B.n871 B.n18 585
R212 B.n870 B.n14 585
R213 B.n975 B.n14 585
R214 B.n869 B.n13 585
R215 B.n976 B.n13 585
R216 B.n868 B.n12 585
R217 B.n977 B.n12 585
R218 B.n867 B.n866 585
R219 B.n866 B.n8 585
R220 B.n865 B.n7 585
R221 B.n983 B.n7 585
R222 B.n864 B.n6 585
R223 B.n984 B.n6 585
R224 B.n863 B.n5 585
R225 B.n985 B.n5 585
R226 B.n862 B.n861 585
R227 B.n861 B.n4 585
R228 B.n860 B.n375 585
R229 B.n860 B.n859 585
R230 B.n850 B.n376 585
R231 B.n377 B.n376 585
R232 B.n852 B.n851 585
R233 B.n853 B.n852 585
R234 B.n849 B.n382 585
R235 B.n382 B.n381 585
R236 B.n848 B.n847 585
R237 B.n847 B.n846 585
R238 B.n384 B.n383 585
R239 B.n839 B.n384 585
R240 B.n838 B.n837 585
R241 B.n840 B.n838 585
R242 B.n836 B.n389 585
R243 B.n389 B.n388 585
R244 B.n835 B.n834 585
R245 B.n834 B.n833 585
R246 B.n391 B.n390 585
R247 B.n392 B.n391 585
R248 B.n826 B.n825 585
R249 B.n827 B.n826 585
R250 B.n824 B.n397 585
R251 B.n397 B.n396 585
R252 B.n823 B.n822 585
R253 B.n822 B.n821 585
R254 B.n399 B.n398 585
R255 B.n400 B.n399 585
R256 B.n814 B.n813 585
R257 B.n815 B.n814 585
R258 B.n812 B.n405 585
R259 B.n405 B.n404 585
R260 B.n811 B.n810 585
R261 B.n810 B.n809 585
R262 B.n407 B.n406 585
R263 B.n408 B.n407 585
R264 B.n802 B.n801 585
R265 B.n803 B.n802 585
R266 B.n800 B.n413 585
R267 B.n413 B.n412 585
R268 B.n799 B.n798 585
R269 B.n798 B.n797 585
R270 B.n415 B.n414 585
R271 B.n416 B.n415 585
R272 B.n790 B.n789 585
R273 B.n791 B.n790 585
R274 B.n788 B.n421 585
R275 B.n421 B.n420 585
R276 B.n787 B.n786 585
R277 B.n786 B.n785 585
R278 B.n423 B.n422 585
R279 B.n424 B.n423 585
R280 B.n778 B.n777 585
R281 B.n779 B.n778 585
R282 B.n776 B.n428 585
R283 B.n432 B.n428 585
R284 B.n775 B.n774 585
R285 B.n774 B.n773 585
R286 B.n430 B.n429 585
R287 B.n431 B.n430 585
R288 B.n766 B.n765 585
R289 B.n767 B.n766 585
R290 B.n764 B.n437 585
R291 B.n437 B.n436 585
R292 B.n763 B.n762 585
R293 B.n762 B.n761 585
R294 B.n439 B.n438 585
R295 B.n440 B.n439 585
R296 B.n754 B.n753 585
R297 B.n755 B.n754 585
R298 B.n443 B.n442 585
R299 B.n510 B.n508 585
R300 B.n511 B.n507 585
R301 B.n511 B.n444 585
R302 B.n514 B.n513 585
R303 B.n515 B.n506 585
R304 B.n517 B.n516 585
R305 B.n519 B.n505 585
R306 B.n522 B.n521 585
R307 B.n523 B.n504 585
R308 B.n525 B.n524 585
R309 B.n527 B.n503 585
R310 B.n530 B.n529 585
R311 B.n531 B.n502 585
R312 B.n533 B.n532 585
R313 B.n535 B.n501 585
R314 B.n538 B.n537 585
R315 B.n539 B.n500 585
R316 B.n541 B.n540 585
R317 B.n543 B.n499 585
R318 B.n546 B.n545 585
R319 B.n547 B.n498 585
R320 B.n549 B.n548 585
R321 B.n551 B.n497 585
R322 B.n554 B.n553 585
R323 B.n555 B.n496 585
R324 B.n557 B.n556 585
R325 B.n559 B.n495 585
R326 B.n562 B.n561 585
R327 B.n563 B.n494 585
R328 B.n565 B.n564 585
R329 B.n567 B.n493 585
R330 B.n570 B.n569 585
R331 B.n571 B.n492 585
R332 B.n573 B.n572 585
R333 B.n575 B.n491 585
R334 B.n578 B.n577 585
R335 B.n579 B.n490 585
R336 B.n581 B.n580 585
R337 B.n583 B.n489 585
R338 B.n586 B.n585 585
R339 B.n587 B.n488 585
R340 B.n589 B.n588 585
R341 B.n591 B.n487 585
R342 B.n594 B.n593 585
R343 B.n595 B.n486 585
R344 B.n597 B.n596 585
R345 B.n599 B.n485 585
R346 B.n602 B.n601 585
R347 B.n603 B.n484 585
R348 B.n605 B.n604 585
R349 B.n607 B.n483 585
R350 B.n610 B.n609 585
R351 B.n611 B.n482 585
R352 B.n613 B.n612 585
R353 B.n615 B.n481 585
R354 B.n618 B.n617 585
R355 B.n620 B.n478 585
R356 B.n622 B.n621 585
R357 B.n624 B.n477 585
R358 B.n627 B.n626 585
R359 B.n628 B.n476 585
R360 B.n630 B.n629 585
R361 B.n632 B.n475 585
R362 B.n635 B.n634 585
R363 B.n636 B.n474 585
R364 B.n641 B.n640 585
R365 B.n643 B.n473 585
R366 B.n646 B.n645 585
R367 B.n647 B.n472 585
R368 B.n649 B.n648 585
R369 B.n651 B.n471 585
R370 B.n654 B.n653 585
R371 B.n655 B.n470 585
R372 B.n657 B.n656 585
R373 B.n659 B.n469 585
R374 B.n662 B.n661 585
R375 B.n663 B.n468 585
R376 B.n665 B.n664 585
R377 B.n667 B.n467 585
R378 B.n670 B.n669 585
R379 B.n671 B.n466 585
R380 B.n673 B.n672 585
R381 B.n675 B.n465 585
R382 B.n678 B.n677 585
R383 B.n679 B.n464 585
R384 B.n681 B.n680 585
R385 B.n683 B.n463 585
R386 B.n686 B.n685 585
R387 B.n687 B.n462 585
R388 B.n689 B.n688 585
R389 B.n691 B.n461 585
R390 B.n694 B.n693 585
R391 B.n695 B.n460 585
R392 B.n697 B.n696 585
R393 B.n699 B.n459 585
R394 B.n702 B.n701 585
R395 B.n703 B.n458 585
R396 B.n705 B.n704 585
R397 B.n707 B.n457 585
R398 B.n710 B.n709 585
R399 B.n711 B.n456 585
R400 B.n713 B.n712 585
R401 B.n715 B.n455 585
R402 B.n718 B.n717 585
R403 B.n719 B.n454 585
R404 B.n721 B.n720 585
R405 B.n723 B.n453 585
R406 B.n726 B.n725 585
R407 B.n727 B.n452 585
R408 B.n729 B.n728 585
R409 B.n731 B.n451 585
R410 B.n734 B.n733 585
R411 B.n735 B.n450 585
R412 B.n737 B.n736 585
R413 B.n739 B.n449 585
R414 B.n742 B.n741 585
R415 B.n743 B.n448 585
R416 B.n745 B.n744 585
R417 B.n747 B.n447 585
R418 B.n748 B.n446 585
R419 B.n751 B.n750 585
R420 B.n752 B.n445 585
R421 B.n445 B.n444 585
R422 B.n757 B.n756 585
R423 B.n756 B.n755 585
R424 B.n758 B.n441 585
R425 B.n441 B.n440 585
R426 B.n760 B.n759 585
R427 B.n761 B.n760 585
R428 B.n435 B.n434 585
R429 B.n436 B.n435 585
R430 B.n769 B.n768 585
R431 B.n768 B.n767 585
R432 B.n770 B.n433 585
R433 B.n433 B.n431 585
R434 B.n772 B.n771 585
R435 B.n773 B.n772 585
R436 B.n427 B.n426 585
R437 B.n432 B.n427 585
R438 B.n781 B.n780 585
R439 B.n780 B.n779 585
R440 B.n782 B.n425 585
R441 B.n425 B.n424 585
R442 B.n784 B.n783 585
R443 B.n785 B.n784 585
R444 B.n419 B.n418 585
R445 B.n420 B.n419 585
R446 B.n793 B.n792 585
R447 B.n792 B.n791 585
R448 B.n794 B.n417 585
R449 B.n417 B.n416 585
R450 B.n796 B.n795 585
R451 B.n797 B.n796 585
R452 B.n411 B.n410 585
R453 B.n412 B.n411 585
R454 B.n805 B.n804 585
R455 B.n804 B.n803 585
R456 B.n806 B.n409 585
R457 B.n409 B.n408 585
R458 B.n808 B.n807 585
R459 B.n809 B.n808 585
R460 B.n403 B.n402 585
R461 B.n404 B.n403 585
R462 B.n817 B.n816 585
R463 B.n816 B.n815 585
R464 B.n818 B.n401 585
R465 B.n401 B.n400 585
R466 B.n820 B.n819 585
R467 B.n821 B.n820 585
R468 B.n395 B.n394 585
R469 B.n396 B.n395 585
R470 B.n829 B.n828 585
R471 B.n828 B.n827 585
R472 B.n830 B.n393 585
R473 B.n393 B.n392 585
R474 B.n832 B.n831 585
R475 B.n833 B.n832 585
R476 B.n387 B.n386 585
R477 B.n388 B.n387 585
R478 B.n842 B.n841 585
R479 B.n841 B.n840 585
R480 B.n843 B.n385 585
R481 B.n839 B.n385 585
R482 B.n845 B.n844 585
R483 B.n846 B.n845 585
R484 B.n380 B.n379 585
R485 B.n381 B.n380 585
R486 B.n855 B.n854 585
R487 B.n854 B.n853 585
R488 B.n856 B.n378 585
R489 B.n378 B.n377 585
R490 B.n858 B.n857 585
R491 B.n859 B.n858 585
R492 B.n2 B.n0 585
R493 B.n4 B.n2 585
R494 B.n3 B.n1 585
R495 B.n984 B.n3 585
R496 B.n982 B.n981 585
R497 B.n983 B.n982 585
R498 B.n980 B.n9 585
R499 B.n9 B.n8 585
R500 B.n979 B.n978 585
R501 B.n978 B.n977 585
R502 B.n11 B.n10 585
R503 B.n976 B.n11 585
R504 B.n974 B.n973 585
R505 B.n975 B.n974 585
R506 B.n972 B.n15 585
R507 B.n18 B.n15 585
R508 B.n971 B.n970 585
R509 B.n970 B.n969 585
R510 B.n17 B.n16 585
R511 B.n968 B.n17 585
R512 B.n966 B.n965 585
R513 B.n967 B.n966 585
R514 B.n964 B.n23 585
R515 B.n23 B.n22 585
R516 B.n963 B.n962 585
R517 B.n962 B.n961 585
R518 B.n25 B.n24 585
R519 B.n960 B.n25 585
R520 B.n958 B.n957 585
R521 B.n959 B.n958 585
R522 B.n956 B.n30 585
R523 B.n30 B.n29 585
R524 B.n955 B.n954 585
R525 B.n954 B.n953 585
R526 B.n32 B.n31 585
R527 B.n952 B.n32 585
R528 B.n950 B.n949 585
R529 B.n951 B.n950 585
R530 B.n948 B.n37 585
R531 B.n37 B.n36 585
R532 B.n947 B.n946 585
R533 B.n946 B.n945 585
R534 B.n39 B.n38 585
R535 B.n944 B.n39 585
R536 B.n942 B.n941 585
R537 B.n943 B.n942 585
R538 B.n940 B.n44 585
R539 B.n44 B.n43 585
R540 B.n939 B.n938 585
R541 B.n938 B.n937 585
R542 B.n46 B.n45 585
R543 B.n936 B.n46 585
R544 B.n934 B.n933 585
R545 B.n935 B.n934 585
R546 B.n932 B.n51 585
R547 B.n51 B.n50 585
R548 B.n931 B.n930 585
R549 B.n930 B.n929 585
R550 B.n53 B.n52 585
R551 B.n928 B.n53 585
R552 B.n926 B.n925 585
R553 B.n927 B.n926 585
R554 B.n924 B.n58 585
R555 B.n58 B.n57 585
R556 B.n923 B.n922 585
R557 B.n922 B.n921 585
R558 B.n60 B.n59 585
R559 B.n920 B.n60 585
R560 B.n918 B.n917 585
R561 B.n919 B.n918 585
R562 B.n916 B.n65 585
R563 B.n65 B.n64 585
R564 B.n915 B.n914 585
R565 B.n914 B.n913 585
R566 B.n987 B.n986 585
R567 B.n986 B.n985 585
R568 B.n756 B.n443 564.573
R569 B.n914 B.n67 564.573
R570 B.n754 B.n445 564.573
R571 B.n910 B.n68 564.573
R572 B.n637 B.t15 352.488
R573 B.n479 B.t11 352.488
R574 B.n133 B.t4 352.488
R575 B.n130 B.t8 352.488
R576 B.n912 B.n911 256.663
R577 B.n912 B.n128 256.663
R578 B.n912 B.n127 256.663
R579 B.n912 B.n126 256.663
R580 B.n912 B.n125 256.663
R581 B.n912 B.n124 256.663
R582 B.n912 B.n123 256.663
R583 B.n912 B.n122 256.663
R584 B.n912 B.n121 256.663
R585 B.n912 B.n120 256.663
R586 B.n912 B.n119 256.663
R587 B.n912 B.n118 256.663
R588 B.n912 B.n117 256.663
R589 B.n912 B.n116 256.663
R590 B.n912 B.n115 256.663
R591 B.n912 B.n114 256.663
R592 B.n912 B.n113 256.663
R593 B.n912 B.n112 256.663
R594 B.n912 B.n111 256.663
R595 B.n912 B.n110 256.663
R596 B.n912 B.n109 256.663
R597 B.n912 B.n108 256.663
R598 B.n912 B.n107 256.663
R599 B.n912 B.n106 256.663
R600 B.n912 B.n105 256.663
R601 B.n912 B.n104 256.663
R602 B.n912 B.n103 256.663
R603 B.n912 B.n102 256.663
R604 B.n912 B.n101 256.663
R605 B.n912 B.n100 256.663
R606 B.n912 B.n99 256.663
R607 B.n912 B.n98 256.663
R608 B.n912 B.n97 256.663
R609 B.n912 B.n96 256.663
R610 B.n912 B.n95 256.663
R611 B.n912 B.n94 256.663
R612 B.n912 B.n93 256.663
R613 B.n912 B.n92 256.663
R614 B.n912 B.n91 256.663
R615 B.n912 B.n90 256.663
R616 B.n912 B.n89 256.663
R617 B.n912 B.n88 256.663
R618 B.n912 B.n87 256.663
R619 B.n912 B.n86 256.663
R620 B.n912 B.n85 256.663
R621 B.n912 B.n84 256.663
R622 B.n912 B.n83 256.663
R623 B.n912 B.n82 256.663
R624 B.n912 B.n81 256.663
R625 B.n912 B.n80 256.663
R626 B.n912 B.n79 256.663
R627 B.n912 B.n78 256.663
R628 B.n912 B.n77 256.663
R629 B.n912 B.n76 256.663
R630 B.n912 B.n75 256.663
R631 B.n912 B.n74 256.663
R632 B.n912 B.n73 256.663
R633 B.n912 B.n72 256.663
R634 B.n912 B.n71 256.663
R635 B.n912 B.n70 256.663
R636 B.n912 B.n69 256.663
R637 B.n509 B.n444 256.663
R638 B.n512 B.n444 256.663
R639 B.n518 B.n444 256.663
R640 B.n520 B.n444 256.663
R641 B.n526 B.n444 256.663
R642 B.n528 B.n444 256.663
R643 B.n534 B.n444 256.663
R644 B.n536 B.n444 256.663
R645 B.n542 B.n444 256.663
R646 B.n544 B.n444 256.663
R647 B.n550 B.n444 256.663
R648 B.n552 B.n444 256.663
R649 B.n558 B.n444 256.663
R650 B.n560 B.n444 256.663
R651 B.n566 B.n444 256.663
R652 B.n568 B.n444 256.663
R653 B.n574 B.n444 256.663
R654 B.n576 B.n444 256.663
R655 B.n582 B.n444 256.663
R656 B.n584 B.n444 256.663
R657 B.n590 B.n444 256.663
R658 B.n592 B.n444 256.663
R659 B.n598 B.n444 256.663
R660 B.n600 B.n444 256.663
R661 B.n606 B.n444 256.663
R662 B.n608 B.n444 256.663
R663 B.n614 B.n444 256.663
R664 B.n616 B.n444 256.663
R665 B.n623 B.n444 256.663
R666 B.n625 B.n444 256.663
R667 B.n631 B.n444 256.663
R668 B.n633 B.n444 256.663
R669 B.n642 B.n444 256.663
R670 B.n644 B.n444 256.663
R671 B.n650 B.n444 256.663
R672 B.n652 B.n444 256.663
R673 B.n658 B.n444 256.663
R674 B.n660 B.n444 256.663
R675 B.n666 B.n444 256.663
R676 B.n668 B.n444 256.663
R677 B.n674 B.n444 256.663
R678 B.n676 B.n444 256.663
R679 B.n682 B.n444 256.663
R680 B.n684 B.n444 256.663
R681 B.n690 B.n444 256.663
R682 B.n692 B.n444 256.663
R683 B.n698 B.n444 256.663
R684 B.n700 B.n444 256.663
R685 B.n706 B.n444 256.663
R686 B.n708 B.n444 256.663
R687 B.n714 B.n444 256.663
R688 B.n716 B.n444 256.663
R689 B.n722 B.n444 256.663
R690 B.n724 B.n444 256.663
R691 B.n730 B.n444 256.663
R692 B.n732 B.n444 256.663
R693 B.n738 B.n444 256.663
R694 B.n740 B.n444 256.663
R695 B.n746 B.n444 256.663
R696 B.n749 B.n444 256.663
R697 B.n756 B.n441 163.367
R698 B.n760 B.n441 163.367
R699 B.n760 B.n435 163.367
R700 B.n768 B.n435 163.367
R701 B.n768 B.n433 163.367
R702 B.n772 B.n433 163.367
R703 B.n772 B.n427 163.367
R704 B.n780 B.n427 163.367
R705 B.n780 B.n425 163.367
R706 B.n784 B.n425 163.367
R707 B.n784 B.n419 163.367
R708 B.n792 B.n419 163.367
R709 B.n792 B.n417 163.367
R710 B.n796 B.n417 163.367
R711 B.n796 B.n411 163.367
R712 B.n804 B.n411 163.367
R713 B.n804 B.n409 163.367
R714 B.n808 B.n409 163.367
R715 B.n808 B.n403 163.367
R716 B.n816 B.n403 163.367
R717 B.n816 B.n401 163.367
R718 B.n820 B.n401 163.367
R719 B.n820 B.n395 163.367
R720 B.n828 B.n395 163.367
R721 B.n828 B.n393 163.367
R722 B.n832 B.n393 163.367
R723 B.n832 B.n387 163.367
R724 B.n841 B.n387 163.367
R725 B.n841 B.n385 163.367
R726 B.n845 B.n385 163.367
R727 B.n845 B.n380 163.367
R728 B.n854 B.n380 163.367
R729 B.n854 B.n378 163.367
R730 B.n858 B.n378 163.367
R731 B.n858 B.n2 163.367
R732 B.n986 B.n2 163.367
R733 B.n986 B.n3 163.367
R734 B.n982 B.n3 163.367
R735 B.n982 B.n9 163.367
R736 B.n978 B.n9 163.367
R737 B.n978 B.n11 163.367
R738 B.n974 B.n11 163.367
R739 B.n974 B.n15 163.367
R740 B.n970 B.n15 163.367
R741 B.n970 B.n17 163.367
R742 B.n966 B.n17 163.367
R743 B.n966 B.n23 163.367
R744 B.n962 B.n23 163.367
R745 B.n962 B.n25 163.367
R746 B.n958 B.n25 163.367
R747 B.n958 B.n30 163.367
R748 B.n954 B.n30 163.367
R749 B.n954 B.n32 163.367
R750 B.n950 B.n32 163.367
R751 B.n950 B.n37 163.367
R752 B.n946 B.n37 163.367
R753 B.n946 B.n39 163.367
R754 B.n942 B.n39 163.367
R755 B.n942 B.n44 163.367
R756 B.n938 B.n44 163.367
R757 B.n938 B.n46 163.367
R758 B.n934 B.n46 163.367
R759 B.n934 B.n51 163.367
R760 B.n930 B.n51 163.367
R761 B.n930 B.n53 163.367
R762 B.n926 B.n53 163.367
R763 B.n926 B.n58 163.367
R764 B.n922 B.n58 163.367
R765 B.n922 B.n60 163.367
R766 B.n918 B.n60 163.367
R767 B.n918 B.n65 163.367
R768 B.n914 B.n65 163.367
R769 B.n511 B.n510 163.367
R770 B.n513 B.n511 163.367
R771 B.n517 B.n506 163.367
R772 B.n521 B.n519 163.367
R773 B.n525 B.n504 163.367
R774 B.n529 B.n527 163.367
R775 B.n533 B.n502 163.367
R776 B.n537 B.n535 163.367
R777 B.n541 B.n500 163.367
R778 B.n545 B.n543 163.367
R779 B.n549 B.n498 163.367
R780 B.n553 B.n551 163.367
R781 B.n557 B.n496 163.367
R782 B.n561 B.n559 163.367
R783 B.n565 B.n494 163.367
R784 B.n569 B.n567 163.367
R785 B.n573 B.n492 163.367
R786 B.n577 B.n575 163.367
R787 B.n581 B.n490 163.367
R788 B.n585 B.n583 163.367
R789 B.n589 B.n488 163.367
R790 B.n593 B.n591 163.367
R791 B.n597 B.n486 163.367
R792 B.n601 B.n599 163.367
R793 B.n605 B.n484 163.367
R794 B.n609 B.n607 163.367
R795 B.n613 B.n482 163.367
R796 B.n617 B.n615 163.367
R797 B.n622 B.n478 163.367
R798 B.n626 B.n624 163.367
R799 B.n630 B.n476 163.367
R800 B.n634 B.n632 163.367
R801 B.n641 B.n474 163.367
R802 B.n645 B.n643 163.367
R803 B.n649 B.n472 163.367
R804 B.n653 B.n651 163.367
R805 B.n657 B.n470 163.367
R806 B.n661 B.n659 163.367
R807 B.n665 B.n468 163.367
R808 B.n669 B.n667 163.367
R809 B.n673 B.n466 163.367
R810 B.n677 B.n675 163.367
R811 B.n681 B.n464 163.367
R812 B.n685 B.n683 163.367
R813 B.n689 B.n462 163.367
R814 B.n693 B.n691 163.367
R815 B.n697 B.n460 163.367
R816 B.n701 B.n699 163.367
R817 B.n705 B.n458 163.367
R818 B.n709 B.n707 163.367
R819 B.n713 B.n456 163.367
R820 B.n717 B.n715 163.367
R821 B.n721 B.n454 163.367
R822 B.n725 B.n723 163.367
R823 B.n729 B.n452 163.367
R824 B.n733 B.n731 163.367
R825 B.n737 B.n450 163.367
R826 B.n741 B.n739 163.367
R827 B.n745 B.n448 163.367
R828 B.n748 B.n747 163.367
R829 B.n750 B.n445 163.367
R830 B.n754 B.n439 163.367
R831 B.n762 B.n439 163.367
R832 B.n762 B.n437 163.367
R833 B.n766 B.n437 163.367
R834 B.n766 B.n430 163.367
R835 B.n774 B.n430 163.367
R836 B.n774 B.n428 163.367
R837 B.n778 B.n428 163.367
R838 B.n778 B.n423 163.367
R839 B.n786 B.n423 163.367
R840 B.n786 B.n421 163.367
R841 B.n790 B.n421 163.367
R842 B.n790 B.n415 163.367
R843 B.n798 B.n415 163.367
R844 B.n798 B.n413 163.367
R845 B.n802 B.n413 163.367
R846 B.n802 B.n407 163.367
R847 B.n810 B.n407 163.367
R848 B.n810 B.n405 163.367
R849 B.n814 B.n405 163.367
R850 B.n814 B.n399 163.367
R851 B.n822 B.n399 163.367
R852 B.n822 B.n397 163.367
R853 B.n826 B.n397 163.367
R854 B.n826 B.n391 163.367
R855 B.n834 B.n391 163.367
R856 B.n834 B.n389 163.367
R857 B.n838 B.n389 163.367
R858 B.n838 B.n384 163.367
R859 B.n847 B.n384 163.367
R860 B.n847 B.n382 163.367
R861 B.n852 B.n382 163.367
R862 B.n852 B.n376 163.367
R863 B.n860 B.n376 163.367
R864 B.n861 B.n860 163.367
R865 B.n861 B.n5 163.367
R866 B.n6 B.n5 163.367
R867 B.n7 B.n6 163.367
R868 B.n866 B.n7 163.367
R869 B.n866 B.n12 163.367
R870 B.n13 B.n12 163.367
R871 B.n14 B.n13 163.367
R872 B.n871 B.n14 163.367
R873 B.n871 B.n19 163.367
R874 B.n20 B.n19 163.367
R875 B.n21 B.n20 163.367
R876 B.n876 B.n21 163.367
R877 B.n876 B.n26 163.367
R878 B.n27 B.n26 163.367
R879 B.n28 B.n27 163.367
R880 B.n881 B.n28 163.367
R881 B.n881 B.n33 163.367
R882 B.n34 B.n33 163.367
R883 B.n35 B.n34 163.367
R884 B.n886 B.n35 163.367
R885 B.n886 B.n40 163.367
R886 B.n41 B.n40 163.367
R887 B.n42 B.n41 163.367
R888 B.n891 B.n42 163.367
R889 B.n891 B.n47 163.367
R890 B.n48 B.n47 163.367
R891 B.n49 B.n48 163.367
R892 B.n896 B.n49 163.367
R893 B.n896 B.n54 163.367
R894 B.n55 B.n54 163.367
R895 B.n56 B.n55 163.367
R896 B.n901 B.n56 163.367
R897 B.n901 B.n61 163.367
R898 B.n62 B.n61 163.367
R899 B.n63 B.n62 163.367
R900 B.n906 B.n63 163.367
R901 B.n906 B.n68 163.367
R902 B.n138 B.n137 163.367
R903 B.n142 B.n141 163.367
R904 B.n146 B.n145 163.367
R905 B.n150 B.n149 163.367
R906 B.n154 B.n153 163.367
R907 B.n158 B.n157 163.367
R908 B.n162 B.n161 163.367
R909 B.n166 B.n165 163.367
R910 B.n170 B.n169 163.367
R911 B.n174 B.n173 163.367
R912 B.n178 B.n177 163.367
R913 B.n182 B.n181 163.367
R914 B.n186 B.n185 163.367
R915 B.n190 B.n189 163.367
R916 B.n194 B.n193 163.367
R917 B.n198 B.n197 163.367
R918 B.n202 B.n201 163.367
R919 B.n206 B.n205 163.367
R920 B.n210 B.n209 163.367
R921 B.n214 B.n213 163.367
R922 B.n218 B.n217 163.367
R923 B.n222 B.n221 163.367
R924 B.n226 B.n225 163.367
R925 B.n230 B.n229 163.367
R926 B.n234 B.n233 163.367
R927 B.n238 B.n237 163.367
R928 B.n242 B.n241 163.367
R929 B.n246 B.n245 163.367
R930 B.n250 B.n249 163.367
R931 B.n254 B.n253 163.367
R932 B.n258 B.n257 163.367
R933 B.n262 B.n261 163.367
R934 B.n266 B.n265 163.367
R935 B.n270 B.n269 163.367
R936 B.n274 B.n273 163.367
R937 B.n278 B.n277 163.367
R938 B.n282 B.n281 163.367
R939 B.n286 B.n285 163.367
R940 B.n290 B.n289 163.367
R941 B.n294 B.n293 163.367
R942 B.n298 B.n297 163.367
R943 B.n302 B.n301 163.367
R944 B.n306 B.n305 163.367
R945 B.n310 B.n309 163.367
R946 B.n314 B.n313 163.367
R947 B.n318 B.n317 163.367
R948 B.n322 B.n321 163.367
R949 B.n326 B.n325 163.367
R950 B.n330 B.n329 163.367
R951 B.n334 B.n333 163.367
R952 B.n338 B.n337 163.367
R953 B.n342 B.n341 163.367
R954 B.n346 B.n345 163.367
R955 B.n350 B.n349 163.367
R956 B.n354 B.n353 163.367
R957 B.n358 B.n357 163.367
R958 B.n362 B.n361 163.367
R959 B.n366 B.n365 163.367
R960 B.n370 B.n369 163.367
R961 B.n372 B.n129 163.367
R962 B.n637 B.t17 129.757
R963 B.n130 B.t9 129.757
R964 B.n479 B.t14 129.736
R965 B.n133 B.t6 129.736
R966 B.n509 B.n443 71.676
R967 B.n513 B.n512 71.676
R968 B.n518 B.n517 71.676
R969 B.n521 B.n520 71.676
R970 B.n526 B.n525 71.676
R971 B.n529 B.n528 71.676
R972 B.n534 B.n533 71.676
R973 B.n537 B.n536 71.676
R974 B.n542 B.n541 71.676
R975 B.n545 B.n544 71.676
R976 B.n550 B.n549 71.676
R977 B.n553 B.n552 71.676
R978 B.n558 B.n557 71.676
R979 B.n561 B.n560 71.676
R980 B.n566 B.n565 71.676
R981 B.n569 B.n568 71.676
R982 B.n574 B.n573 71.676
R983 B.n577 B.n576 71.676
R984 B.n582 B.n581 71.676
R985 B.n585 B.n584 71.676
R986 B.n590 B.n589 71.676
R987 B.n593 B.n592 71.676
R988 B.n598 B.n597 71.676
R989 B.n601 B.n600 71.676
R990 B.n606 B.n605 71.676
R991 B.n609 B.n608 71.676
R992 B.n614 B.n613 71.676
R993 B.n617 B.n616 71.676
R994 B.n623 B.n622 71.676
R995 B.n626 B.n625 71.676
R996 B.n631 B.n630 71.676
R997 B.n634 B.n633 71.676
R998 B.n642 B.n641 71.676
R999 B.n645 B.n644 71.676
R1000 B.n650 B.n649 71.676
R1001 B.n653 B.n652 71.676
R1002 B.n658 B.n657 71.676
R1003 B.n661 B.n660 71.676
R1004 B.n666 B.n665 71.676
R1005 B.n669 B.n668 71.676
R1006 B.n674 B.n673 71.676
R1007 B.n677 B.n676 71.676
R1008 B.n682 B.n681 71.676
R1009 B.n685 B.n684 71.676
R1010 B.n690 B.n689 71.676
R1011 B.n693 B.n692 71.676
R1012 B.n698 B.n697 71.676
R1013 B.n701 B.n700 71.676
R1014 B.n706 B.n705 71.676
R1015 B.n709 B.n708 71.676
R1016 B.n714 B.n713 71.676
R1017 B.n717 B.n716 71.676
R1018 B.n722 B.n721 71.676
R1019 B.n725 B.n724 71.676
R1020 B.n730 B.n729 71.676
R1021 B.n733 B.n732 71.676
R1022 B.n738 B.n737 71.676
R1023 B.n741 B.n740 71.676
R1024 B.n746 B.n745 71.676
R1025 B.n749 B.n748 71.676
R1026 B.n69 B.n67 71.676
R1027 B.n138 B.n70 71.676
R1028 B.n142 B.n71 71.676
R1029 B.n146 B.n72 71.676
R1030 B.n150 B.n73 71.676
R1031 B.n154 B.n74 71.676
R1032 B.n158 B.n75 71.676
R1033 B.n162 B.n76 71.676
R1034 B.n166 B.n77 71.676
R1035 B.n170 B.n78 71.676
R1036 B.n174 B.n79 71.676
R1037 B.n178 B.n80 71.676
R1038 B.n182 B.n81 71.676
R1039 B.n186 B.n82 71.676
R1040 B.n190 B.n83 71.676
R1041 B.n194 B.n84 71.676
R1042 B.n198 B.n85 71.676
R1043 B.n202 B.n86 71.676
R1044 B.n206 B.n87 71.676
R1045 B.n210 B.n88 71.676
R1046 B.n214 B.n89 71.676
R1047 B.n218 B.n90 71.676
R1048 B.n222 B.n91 71.676
R1049 B.n226 B.n92 71.676
R1050 B.n230 B.n93 71.676
R1051 B.n234 B.n94 71.676
R1052 B.n238 B.n95 71.676
R1053 B.n242 B.n96 71.676
R1054 B.n246 B.n97 71.676
R1055 B.n250 B.n98 71.676
R1056 B.n254 B.n99 71.676
R1057 B.n258 B.n100 71.676
R1058 B.n262 B.n101 71.676
R1059 B.n266 B.n102 71.676
R1060 B.n270 B.n103 71.676
R1061 B.n274 B.n104 71.676
R1062 B.n278 B.n105 71.676
R1063 B.n282 B.n106 71.676
R1064 B.n286 B.n107 71.676
R1065 B.n290 B.n108 71.676
R1066 B.n294 B.n109 71.676
R1067 B.n298 B.n110 71.676
R1068 B.n302 B.n111 71.676
R1069 B.n306 B.n112 71.676
R1070 B.n310 B.n113 71.676
R1071 B.n314 B.n114 71.676
R1072 B.n318 B.n115 71.676
R1073 B.n322 B.n116 71.676
R1074 B.n326 B.n117 71.676
R1075 B.n330 B.n118 71.676
R1076 B.n334 B.n119 71.676
R1077 B.n338 B.n120 71.676
R1078 B.n342 B.n121 71.676
R1079 B.n346 B.n122 71.676
R1080 B.n350 B.n123 71.676
R1081 B.n354 B.n124 71.676
R1082 B.n358 B.n125 71.676
R1083 B.n362 B.n126 71.676
R1084 B.n366 B.n127 71.676
R1085 B.n370 B.n128 71.676
R1086 B.n911 B.n129 71.676
R1087 B.n911 B.n910 71.676
R1088 B.n372 B.n128 71.676
R1089 B.n369 B.n127 71.676
R1090 B.n365 B.n126 71.676
R1091 B.n361 B.n125 71.676
R1092 B.n357 B.n124 71.676
R1093 B.n353 B.n123 71.676
R1094 B.n349 B.n122 71.676
R1095 B.n345 B.n121 71.676
R1096 B.n341 B.n120 71.676
R1097 B.n337 B.n119 71.676
R1098 B.n333 B.n118 71.676
R1099 B.n329 B.n117 71.676
R1100 B.n325 B.n116 71.676
R1101 B.n321 B.n115 71.676
R1102 B.n317 B.n114 71.676
R1103 B.n313 B.n113 71.676
R1104 B.n309 B.n112 71.676
R1105 B.n305 B.n111 71.676
R1106 B.n301 B.n110 71.676
R1107 B.n297 B.n109 71.676
R1108 B.n293 B.n108 71.676
R1109 B.n289 B.n107 71.676
R1110 B.n285 B.n106 71.676
R1111 B.n281 B.n105 71.676
R1112 B.n277 B.n104 71.676
R1113 B.n273 B.n103 71.676
R1114 B.n269 B.n102 71.676
R1115 B.n265 B.n101 71.676
R1116 B.n261 B.n100 71.676
R1117 B.n257 B.n99 71.676
R1118 B.n253 B.n98 71.676
R1119 B.n249 B.n97 71.676
R1120 B.n245 B.n96 71.676
R1121 B.n241 B.n95 71.676
R1122 B.n237 B.n94 71.676
R1123 B.n233 B.n93 71.676
R1124 B.n229 B.n92 71.676
R1125 B.n225 B.n91 71.676
R1126 B.n221 B.n90 71.676
R1127 B.n217 B.n89 71.676
R1128 B.n213 B.n88 71.676
R1129 B.n209 B.n87 71.676
R1130 B.n205 B.n86 71.676
R1131 B.n201 B.n85 71.676
R1132 B.n197 B.n84 71.676
R1133 B.n193 B.n83 71.676
R1134 B.n189 B.n82 71.676
R1135 B.n185 B.n81 71.676
R1136 B.n181 B.n80 71.676
R1137 B.n177 B.n79 71.676
R1138 B.n173 B.n78 71.676
R1139 B.n169 B.n77 71.676
R1140 B.n165 B.n76 71.676
R1141 B.n161 B.n75 71.676
R1142 B.n157 B.n74 71.676
R1143 B.n153 B.n73 71.676
R1144 B.n149 B.n72 71.676
R1145 B.n145 B.n71 71.676
R1146 B.n141 B.n70 71.676
R1147 B.n137 B.n69 71.676
R1148 B.n510 B.n509 71.676
R1149 B.n512 B.n506 71.676
R1150 B.n519 B.n518 71.676
R1151 B.n520 B.n504 71.676
R1152 B.n527 B.n526 71.676
R1153 B.n528 B.n502 71.676
R1154 B.n535 B.n534 71.676
R1155 B.n536 B.n500 71.676
R1156 B.n543 B.n542 71.676
R1157 B.n544 B.n498 71.676
R1158 B.n551 B.n550 71.676
R1159 B.n552 B.n496 71.676
R1160 B.n559 B.n558 71.676
R1161 B.n560 B.n494 71.676
R1162 B.n567 B.n566 71.676
R1163 B.n568 B.n492 71.676
R1164 B.n575 B.n574 71.676
R1165 B.n576 B.n490 71.676
R1166 B.n583 B.n582 71.676
R1167 B.n584 B.n488 71.676
R1168 B.n591 B.n590 71.676
R1169 B.n592 B.n486 71.676
R1170 B.n599 B.n598 71.676
R1171 B.n600 B.n484 71.676
R1172 B.n607 B.n606 71.676
R1173 B.n608 B.n482 71.676
R1174 B.n615 B.n614 71.676
R1175 B.n616 B.n478 71.676
R1176 B.n624 B.n623 71.676
R1177 B.n625 B.n476 71.676
R1178 B.n632 B.n631 71.676
R1179 B.n633 B.n474 71.676
R1180 B.n643 B.n642 71.676
R1181 B.n644 B.n472 71.676
R1182 B.n651 B.n650 71.676
R1183 B.n652 B.n470 71.676
R1184 B.n659 B.n658 71.676
R1185 B.n660 B.n468 71.676
R1186 B.n667 B.n666 71.676
R1187 B.n668 B.n466 71.676
R1188 B.n675 B.n674 71.676
R1189 B.n676 B.n464 71.676
R1190 B.n683 B.n682 71.676
R1191 B.n684 B.n462 71.676
R1192 B.n691 B.n690 71.676
R1193 B.n692 B.n460 71.676
R1194 B.n699 B.n698 71.676
R1195 B.n700 B.n458 71.676
R1196 B.n707 B.n706 71.676
R1197 B.n708 B.n456 71.676
R1198 B.n715 B.n714 71.676
R1199 B.n716 B.n454 71.676
R1200 B.n723 B.n722 71.676
R1201 B.n724 B.n452 71.676
R1202 B.n731 B.n730 71.676
R1203 B.n732 B.n450 71.676
R1204 B.n739 B.n738 71.676
R1205 B.n740 B.n448 71.676
R1206 B.n747 B.n746 71.676
R1207 B.n750 B.n749 71.676
R1208 B.n638 B.t16 68.0851
R1209 B.n131 B.t10 68.0851
R1210 B.n480 B.t13 68.0624
R1211 B.n134 B.t7 68.0624
R1212 B.n755 B.n444 66.5477
R1213 B.n913 B.n912 66.5477
R1214 B.n638 B.n637 61.6732
R1215 B.n480 B.n479 61.6732
R1216 B.n134 B.n133 61.6732
R1217 B.n131 B.n130 61.6732
R1218 B.n639 B.n638 59.5399
R1219 B.n619 B.n480 59.5399
R1220 B.n135 B.n134 59.5399
R1221 B.n132 B.n131 59.5399
R1222 B.n915 B.n66 36.6834
R1223 B.n909 B.n908 36.6834
R1224 B.n753 B.n752 36.6834
R1225 B.n757 B.n442 36.6834
R1226 B.n755 B.n440 33.5206
R1227 B.n761 B.n440 33.5206
R1228 B.n761 B.n436 33.5206
R1229 B.n767 B.n436 33.5206
R1230 B.n767 B.n431 33.5206
R1231 B.n773 B.n431 33.5206
R1232 B.n773 B.n432 33.5206
R1233 B.n779 B.n424 33.5206
R1234 B.n785 B.n424 33.5206
R1235 B.n785 B.n420 33.5206
R1236 B.n791 B.n420 33.5206
R1237 B.n791 B.n416 33.5206
R1238 B.n797 B.n416 33.5206
R1239 B.n797 B.n412 33.5206
R1240 B.n803 B.n412 33.5206
R1241 B.n803 B.n408 33.5206
R1242 B.n809 B.n408 33.5206
R1243 B.n809 B.n404 33.5206
R1244 B.n815 B.n404 33.5206
R1245 B.n821 B.n400 33.5206
R1246 B.n821 B.n396 33.5206
R1247 B.n827 B.n396 33.5206
R1248 B.n827 B.n392 33.5206
R1249 B.n833 B.n392 33.5206
R1250 B.n833 B.n388 33.5206
R1251 B.n840 B.n388 33.5206
R1252 B.n840 B.n839 33.5206
R1253 B.n846 B.n381 33.5206
R1254 B.n853 B.n381 33.5206
R1255 B.n853 B.n377 33.5206
R1256 B.n859 B.n377 33.5206
R1257 B.n859 B.n4 33.5206
R1258 B.n985 B.n4 33.5206
R1259 B.n985 B.n984 33.5206
R1260 B.n984 B.n983 33.5206
R1261 B.n983 B.n8 33.5206
R1262 B.n977 B.n8 33.5206
R1263 B.n977 B.n976 33.5206
R1264 B.n976 B.n975 33.5206
R1265 B.n969 B.n18 33.5206
R1266 B.n969 B.n968 33.5206
R1267 B.n968 B.n967 33.5206
R1268 B.n967 B.n22 33.5206
R1269 B.n961 B.n22 33.5206
R1270 B.n961 B.n960 33.5206
R1271 B.n960 B.n959 33.5206
R1272 B.n959 B.n29 33.5206
R1273 B.n953 B.n952 33.5206
R1274 B.n952 B.n951 33.5206
R1275 B.n951 B.n36 33.5206
R1276 B.n945 B.n36 33.5206
R1277 B.n945 B.n944 33.5206
R1278 B.n944 B.n943 33.5206
R1279 B.n943 B.n43 33.5206
R1280 B.n937 B.n43 33.5206
R1281 B.n937 B.n936 33.5206
R1282 B.n936 B.n935 33.5206
R1283 B.n935 B.n50 33.5206
R1284 B.n929 B.n50 33.5206
R1285 B.n928 B.n927 33.5206
R1286 B.n927 B.n57 33.5206
R1287 B.n921 B.n57 33.5206
R1288 B.n921 B.n920 33.5206
R1289 B.n920 B.n919 33.5206
R1290 B.n919 B.n64 33.5206
R1291 B.n913 B.n64 33.5206
R1292 B.n432 B.t12 27.1123
R1293 B.t5 B.n928 27.1123
R1294 B.n839 B.t0 24.1547
R1295 B.n18 B.t3 24.1547
R1296 B.t2 B.n400 21.197
R1297 B.t1 B.n29 21.197
R1298 B B.n987 18.0485
R1299 B.n815 B.t2 12.324
R1300 B.n953 B.t1 12.324
R1301 B.n136 B.n66 10.6151
R1302 B.n139 B.n136 10.6151
R1303 B.n140 B.n139 10.6151
R1304 B.n143 B.n140 10.6151
R1305 B.n144 B.n143 10.6151
R1306 B.n147 B.n144 10.6151
R1307 B.n148 B.n147 10.6151
R1308 B.n151 B.n148 10.6151
R1309 B.n152 B.n151 10.6151
R1310 B.n155 B.n152 10.6151
R1311 B.n156 B.n155 10.6151
R1312 B.n159 B.n156 10.6151
R1313 B.n160 B.n159 10.6151
R1314 B.n163 B.n160 10.6151
R1315 B.n164 B.n163 10.6151
R1316 B.n167 B.n164 10.6151
R1317 B.n168 B.n167 10.6151
R1318 B.n171 B.n168 10.6151
R1319 B.n172 B.n171 10.6151
R1320 B.n175 B.n172 10.6151
R1321 B.n176 B.n175 10.6151
R1322 B.n179 B.n176 10.6151
R1323 B.n180 B.n179 10.6151
R1324 B.n183 B.n180 10.6151
R1325 B.n184 B.n183 10.6151
R1326 B.n187 B.n184 10.6151
R1327 B.n188 B.n187 10.6151
R1328 B.n191 B.n188 10.6151
R1329 B.n192 B.n191 10.6151
R1330 B.n195 B.n192 10.6151
R1331 B.n196 B.n195 10.6151
R1332 B.n199 B.n196 10.6151
R1333 B.n200 B.n199 10.6151
R1334 B.n203 B.n200 10.6151
R1335 B.n204 B.n203 10.6151
R1336 B.n207 B.n204 10.6151
R1337 B.n208 B.n207 10.6151
R1338 B.n211 B.n208 10.6151
R1339 B.n212 B.n211 10.6151
R1340 B.n215 B.n212 10.6151
R1341 B.n216 B.n215 10.6151
R1342 B.n219 B.n216 10.6151
R1343 B.n220 B.n219 10.6151
R1344 B.n223 B.n220 10.6151
R1345 B.n224 B.n223 10.6151
R1346 B.n227 B.n224 10.6151
R1347 B.n228 B.n227 10.6151
R1348 B.n231 B.n228 10.6151
R1349 B.n232 B.n231 10.6151
R1350 B.n235 B.n232 10.6151
R1351 B.n236 B.n235 10.6151
R1352 B.n239 B.n236 10.6151
R1353 B.n240 B.n239 10.6151
R1354 B.n243 B.n240 10.6151
R1355 B.n244 B.n243 10.6151
R1356 B.n248 B.n247 10.6151
R1357 B.n251 B.n248 10.6151
R1358 B.n252 B.n251 10.6151
R1359 B.n255 B.n252 10.6151
R1360 B.n256 B.n255 10.6151
R1361 B.n259 B.n256 10.6151
R1362 B.n260 B.n259 10.6151
R1363 B.n263 B.n260 10.6151
R1364 B.n264 B.n263 10.6151
R1365 B.n268 B.n267 10.6151
R1366 B.n271 B.n268 10.6151
R1367 B.n272 B.n271 10.6151
R1368 B.n275 B.n272 10.6151
R1369 B.n276 B.n275 10.6151
R1370 B.n279 B.n276 10.6151
R1371 B.n280 B.n279 10.6151
R1372 B.n283 B.n280 10.6151
R1373 B.n284 B.n283 10.6151
R1374 B.n287 B.n284 10.6151
R1375 B.n288 B.n287 10.6151
R1376 B.n291 B.n288 10.6151
R1377 B.n292 B.n291 10.6151
R1378 B.n295 B.n292 10.6151
R1379 B.n296 B.n295 10.6151
R1380 B.n299 B.n296 10.6151
R1381 B.n300 B.n299 10.6151
R1382 B.n303 B.n300 10.6151
R1383 B.n304 B.n303 10.6151
R1384 B.n307 B.n304 10.6151
R1385 B.n308 B.n307 10.6151
R1386 B.n311 B.n308 10.6151
R1387 B.n312 B.n311 10.6151
R1388 B.n315 B.n312 10.6151
R1389 B.n316 B.n315 10.6151
R1390 B.n319 B.n316 10.6151
R1391 B.n320 B.n319 10.6151
R1392 B.n323 B.n320 10.6151
R1393 B.n324 B.n323 10.6151
R1394 B.n327 B.n324 10.6151
R1395 B.n328 B.n327 10.6151
R1396 B.n331 B.n328 10.6151
R1397 B.n332 B.n331 10.6151
R1398 B.n335 B.n332 10.6151
R1399 B.n336 B.n335 10.6151
R1400 B.n339 B.n336 10.6151
R1401 B.n340 B.n339 10.6151
R1402 B.n343 B.n340 10.6151
R1403 B.n344 B.n343 10.6151
R1404 B.n347 B.n344 10.6151
R1405 B.n348 B.n347 10.6151
R1406 B.n351 B.n348 10.6151
R1407 B.n352 B.n351 10.6151
R1408 B.n355 B.n352 10.6151
R1409 B.n356 B.n355 10.6151
R1410 B.n359 B.n356 10.6151
R1411 B.n360 B.n359 10.6151
R1412 B.n363 B.n360 10.6151
R1413 B.n364 B.n363 10.6151
R1414 B.n367 B.n364 10.6151
R1415 B.n368 B.n367 10.6151
R1416 B.n371 B.n368 10.6151
R1417 B.n373 B.n371 10.6151
R1418 B.n374 B.n373 10.6151
R1419 B.n909 B.n374 10.6151
R1420 B.n753 B.n438 10.6151
R1421 B.n763 B.n438 10.6151
R1422 B.n764 B.n763 10.6151
R1423 B.n765 B.n764 10.6151
R1424 B.n765 B.n429 10.6151
R1425 B.n775 B.n429 10.6151
R1426 B.n776 B.n775 10.6151
R1427 B.n777 B.n776 10.6151
R1428 B.n777 B.n422 10.6151
R1429 B.n787 B.n422 10.6151
R1430 B.n788 B.n787 10.6151
R1431 B.n789 B.n788 10.6151
R1432 B.n789 B.n414 10.6151
R1433 B.n799 B.n414 10.6151
R1434 B.n800 B.n799 10.6151
R1435 B.n801 B.n800 10.6151
R1436 B.n801 B.n406 10.6151
R1437 B.n811 B.n406 10.6151
R1438 B.n812 B.n811 10.6151
R1439 B.n813 B.n812 10.6151
R1440 B.n813 B.n398 10.6151
R1441 B.n823 B.n398 10.6151
R1442 B.n824 B.n823 10.6151
R1443 B.n825 B.n824 10.6151
R1444 B.n825 B.n390 10.6151
R1445 B.n835 B.n390 10.6151
R1446 B.n836 B.n835 10.6151
R1447 B.n837 B.n836 10.6151
R1448 B.n837 B.n383 10.6151
R1449 B.n848 B.n383 10.6151
R1450 B.n849 B.n848 10.6151
R1451 B.n851 B.n849 10.6151
R1452 B.n851 B.n850 10.6151
R1453 B.n850 B.n375 10.6151
R1454 B.n862 B.n375 10.6151
R1455 B.n863 B.n862 10.6151
R1456 B.n864 B.n863 10.6151
R1457 B.n865 B.n864 10.6151
R1458 B.n867 B.n865 10.6151
R1459 B.n868 B.n867 10.6151
R1460 B.n869 B.n868 10.6151
R1461 B.n870 B.n869 10.6151
R1462 B.n872 B.n870 10.6151
R1463 B.n873 B.n872 10.6151
R1464 B.n874 B.n873 10.6151
R1465 B.n875 B.n874 10.6151
R1466 B.n877 B.n875 10.6151
R1467 B.n878 B.n877 10.6151
R1468 B.n879 B.n878 10.6151
R1469 B.n880 B.n879 10.6151
R1470 B.n882 B.n880 10.6151
R1471 B.n883 B.n882 10.6151
R1472 B.n884 B.n883 10.6151
R1473 B.n885 B.n884 10.6151
R1474 B.n887 B.n885 10.6151
R1475 B.n888 B.n887 10.6151
R1476 B.n889 B.n888 10.6151
R1477 B.n890 B.n889 10.6151
R1478 B.n892 B.n890 10.6151
R1479 B.n893 B.n892 10.6151
R1480 B.n894 B.n893 10.6151
R1481 B.n895 B.n894 10.6151
R1482 B.n897 B.n895 10.6151
R1483 B.n898 B.n897 10.6151
R1484 B.n899 B.n898 10.6151
R1485 B.n900 B.n899 10.6151
R1486 B.n902 B.n900 10.6151
R1487 B.n903 B.n902 10.6151
R1488 B.n904 B.n903 10.6151
R1489 B.n905 B.n904 10.6151
R1490 B.n907 B.n905 10.6151
R1491 B.n908 B.n907 10.6151
R1492 B.n508 B.n442 10.6151
R1493 B.n508 B.n507 10.6151
R1494 B.n514 B.n507 10.6151
R1495 B.n515 B.n514 10.6151
R1496 B.n516 B.n515 10.6151
R1497 B.n516 B.n505 10.6151
R1498 B.n522 B.n505 10.6151
R1499 B.n523 B.n522 10.6151
R1500 B.n524 B.n523 10.6151
R1501 B.n524 B.n503 10.6151
R1502 B.n530 B.n503 10.6151
R1503 B.n531 B.n530 10.6151
R1504 B.n532 B.n531 10.6151
R1505 B.n532 B.n501 10.6151
R1506 B.n538 B.n501 10.6151
R1507 B.n539 B.n538 10.6151
R1508 B.n540 B.n539 10.6151
R1509 B.n540 B.n499 10.6151
R1510 B.n546 B.n499 10.6151
R1511 B.n547 B.n546 10.6151
R1512 B.n548 B.n547 10.6151
R1513 B.n548 B.n497 10.6151
R1514 B.n554 B.n497 10.6151
R1515 B.n555 B.n554 10.6151
R1516 B.n556 B.n555 10.6151
R1517 B.n556 B.n495 10.6151
R1518 B.n562 B.n495 10.6151
R1519 B.n563 B.n562 10.6151
R1520 B.n564 B.n563 10.6151
R1521 B.n564 B.n493 10.6151
R1522 B.n570 B.n493 10.6151
R1523 B.n571 B.n570 10.6151
R1524 B.n572 B.n571 10.6151
R1525 B.n572 B.n491 10.6151
R1526 B.n578 B.n491 10.6151
R1527 B.n579 B.n578 10.6151
R1528 B.n580 B.n579 10.6151
R1529 B.n580 B.n489 10.6151
R1530 B.n586 B.n489 10.6151
R1531 B.n587 B.n586 10.6151
R1532 B.n588 B.n587 10.6151
R1533 B.n588 B.n487 10.6151
R1534 B.n594 B.n487 10.6151
R1535 B.n595 B.n594 10.6151
R1536 B.n596 B.n595 10.6151
R1537 B.n596 B.n485 10.6151
R1538 B.n602 B.n485 10.6151
R1539 B.n603 B.n602 10.6151
R1540 B.n604 B.n603 10.6151
R1541 B.n604 B.n483 10.6151
R1542 B.n610 B.n483 10.6151
R1543 B.n611 B.n610 10.6151
R1544 B.n612 B.n611 10.6151
R1545 B.n612 B.n481 10.6151
R1546 B.n618 B.n481 10.6151
R1547 B.n621 B.n620 10.6151
R1548 B.n621 B.n477 10.6151
R1549 B.n627 B.n477 10.6151
R1550 B.n628 B.n627 10.6151
R1551 B.n629 B.n628 10.6151
R1552 B.n629 B.n475 10.6151
R1553 B.n635 B.n475 10.6151
R1554 B.n636 B.n635 10.6151
R1555 B.n640 B.n636 10.6151
R1556 B.n646 B.n473 10.6151
R1557 B.n647 B.n646 10.6151
R1558 B.n648 B.n647 10.6151
R1559 B.n648 B.n471 10.6151
R1560 B.n654 B.n471 10.6151
R1561 B.n655 B.n654 10.6151
R1562 B.n656 B.n655 10.6151
R1563 B.n656 B.n469 10.6151
R1564 B.n662 B.n469 10.6151
R1565 B.n663 B.n662 10.6151
R1566 B.n664 B.n663 10.6151
R1567 B.n664 B.n467 10.6151
R1568 B.n670 B.n467 10.6151
R1569 B.n671 B.n670 10.6151
R1570 B.n672 B.n671 10.6151
R1571 B.n672 B.n465 10.6151
R1572 B.n678 B.n465 10.6151
R1573 B.n679 B.n678 10.6151
R1574 B.n680 B.n679 10.6151
R1575 B.n680 B.n463 10.6151
R1576 B.n686 B.n463 10.6151
R1577 B.n687 B.n686 10.6151
R1578 B.n688 B.n687 10.6151
R1579 B.n688 B.n461 10.6151
R1580 B.n694 B.n461 10.6151
R1581 B.n695 B.n694 10.6151
R1582 B.n696 B.n695 10.6151
R1583 B.n696 B.n459 10.6151
R1584 B.n702 B.n459 10.6151
R1585 B.n703 B.n702 10.6151
R1586 B.n704 B.n703 10.6151
R1587 B.n704 B.n457 10.6151
R1588 B.n710 B.n457 10.6151
R1589 B.n711 B.n710 10.6151
R1590 B.n712 B.n711 10.6151
R1591 B.n712 B.n455 10.6151
R1592 B.n718 B.n455 10.6151
R1593 B.n719 B.n718 10.6151
R1594 B.n720 B.n719 10.6151
R1595 B.n720 B.n453 10.6151
R1596 B.n726 B.n453 10.6151
R1597 B.n727 B.n726 10.6151
R1598 B.n728 B.n727 10.6151
R1599 B.n728 B.n451 10.6151
R1600 B.n734 B.n451 10.6151
R1601 B.n735 B.n734 10.6151
R1602 B.n736 B.n735 10.6151
R1603 B.n736 B.n449 10.6151
R1604 B.n742 B.n449 10.6151
R1605 B.n743 B.n742 10.6151
R1606 B.n744 B.n743 10.6151
R1607 B.n744 B.n447 10.6151
R1608 B.n447 B.n446 10.6151
R1609 B.n751 B.n446 10.6151
R1610 B.n752 B.n751 10.6151
R1611 B.n758 B.n757 10.6151
R1612 B.n759 B.n758 10.6151
R1613 B.n759 B.n434 10.6151
R1614 B.n769 B.n434 10.6151
R1615 B.n770 B.n769 10.6151
R1616 B.n771 B.n770 10.6151
R1617 B.n771 B.n426 10.6151
R1618 B.n781 B.n426 10.6151
R1619 B.n782 B.n781 10.6151
R1620 B.n783 B.n782 10.6151
R1621 B.n783 B.n418 10.6151
R1622 B.n793 B.n418 10.6151
R1623 B.n794 B.n793 10.6151
R1624 B.n795 B.n794 10.6151
R1625 B.n795 B.n410 10.6151
R1626 B.n805 B.n410 10.6151
R1627 B.n806 B.n805 10.6151
R1628 B.n807 B.n806 10.6151
R1629 B.n807 B.n402 10.6151
R1630 B.n817 B.n402 10.6151
R1631 B.n818 B.n817 10.6151
R1632 B.n819 B.n818 10.6151
R1633 B.n819 B.n394 10.6151
R1634 B.n829 B.n394 10.6151
R1635 B.n830 B.n829 10.6151
R1636 B.n831 B.n830 10.6151
R1637 B.n831 B.n386 10.6151
R1638 B.n842 B.n386 10.6151
R1639 B.n843 B.n842 10.6151
R1640 B.n844 B.n843 10.6151
R1641 B.n844 B.n379 10.6151
R1642 B.n855 B.n379 10.6151
R1643 B.n856 B.n855 10.6151
R1644 B.n857 B.n856 10.6151
R1645 B.n857 B.n0 10.6151
R1646 B.n981 B.n1 10.6151
R1647 B.n981 B.n980 10.6151
R1648 B.n980 B.n979 10.6151
R1649 B.n979 B.n10 10.6151
R1650 B.n973 B.n10 10.6151
R1651 B.n973 B.n972 10.6151
R1652 B.n972 B.n971 10.6151
R1653 B.n971 B.n16 10.6151
R1654 B.n965 B.n16 10.6151
R1655 B.n965 B.n964 10.6151
R1656 B.n964 B.n963 10.6151
R1657 B.n963 B.n24 10.6151
R1658 B.n957 B.n24 10.6151
R1659 B.n957 B.n956 10.6151
R1660 B.n956 B.n955 10.6151
R1661 B.n955 B.n31 10.6151
R1662 B.n949 B.n31 10.6151
R1663 B.n949 B.n948 10.6151
R1664 B.n948 B.n947 10.6151
R1665 B.n947 B.n38 10.6151
R1666 B.n941 B.n38 10.6151
R1667 B.n941 B.n940 10.6151
R1668 B.n940 B.n939 10.6151
R1669 B.n939 B.n45 10.6151
R1670 B.n933 B.n45 10.6151
R1671 B.n933 B.n932 10.6151
R1672 B.n932 B.n931 10.6151
R1673 B.n931 B.n52 10.6151
R1674 B.n925 B.n52 10.6151
R1675 B.n925 B.n924 10.6151
R1676 B.n924 B.n923 10.6151
R1677 B.n923 B.n59 10.6151
R1678 B.n917 B.n59 10.6151
R1679 B.n917 B.n916 10.6151
R1680 B.n916 B.n915 10.6151
R1681 B.n846 B.t0 9.3664
R1682 B.n975 B.t3 9.3664
R1683 B.n244 B.n135 9.36635
R1684 B.n267 B.n132 9.36635
R1685 B.n619 B.n618 9.36635
R1686 B.n639 B.n473 9.36635
R1687 B.n779 B.t12 6.40875
R1688 B.n929 B.t5 6.40875
R1689 B.n987 B.n0 2.81026
R1690 B.n987 B.n1 2.81026
R1691 B.n247 B.n135 1.24928
R1692 B.n264 B.n132 1.24928
R1693 B.n620 B.n619 1.24928
R1694 B.n640 B.n639 1.24928
R1695 VP.n4 VP.t0 179.571
R1696 VP.n4 VP.t3 178.672
R1697 VP.n16 VP.n0 161.3
R1698 VP.n15 VP.n14 161.3
R1699 VP.n13 VP.n1 161.3
R1700 VP.n12 VP.n11 161.3
R1701 VP.n10 VP.n2 161.3
R1702 VP.n9 VP.n8 161.3
R1703 VP.n7 VP.n3 161.3
R1704 VP.n5 VP.t1 144.094
R1705 VP.n17 VP.t2 144.094
R1706 VP.n6 VP.n5 106.481
R1707 VP.n18 VP.n17 106.481
R1708 VP.n6 VP.n4 54.3317
R1709 VP.n11 VP.n10 40.577
R1710 VP.n11 VP.n1 40.577
R1711 VP.n9 VP.n3 24.5923
R1712 VP.n10 VP.n9 24.5923
R1713 VP.n15 VP.n1 24.5923
R1714 VP.n16 VP.n15 24.5923
R1715 VP.n5 VP.n3 4.42703
R1716 VP.n17 VP.n16 4.42703
R1717 VP.n7 VP.n6 0.278335
R1718 VP.n18 VP.n0 0.278335
R1719 VP.n8 VP.n7 0.189894
R1720 VP.n8 VP.n2 0.189894
R1721 VP.n12 VP.n2 0.189894
R1722 VP.n13 VP.n12 0.189894
R1723 VP.n14 VP.n13 0.189894
R1724 VP.n14 VP.n0 0.189894
R1725 VP VP.n18 0.153485
R1726 VDD1 VDD1.n1 105.528
R1727 VDD1 VDD1.n0 58.4328
R1728 VDD1.n0 VDD1.t3 1.16247
R1729 VDD1.n0 VDD1.t0 1.16247
R1730 VDD1.n1 VDD1.t2 1.16247
R1731 VDD1.n1 VDD1.t1 1.16247
C0 VDD2 VTAIL 6.66741f
C1 VN VTAIL 6.44143f
C2 VDD1 VTAIL 6.61153f
C3 VP VTAIL 6.45554f
C4 VDD2 VN 6.724259f
C5 VDD2 VDD1 1.0826f
C6 VP VDD2 0.410386f
C7 VN VDD1 0.149399f
C8 VP VN 7.29868f
C9 VP VDD1 6.98445f
C10 VDD2 B 4.301904f
C11 VDD1 B 9.01824f
C12 VTAIL B 13.256029f
C13 VN B 11.56651f
C14 VP B 9.798078f
C15 VDD1.t3 B 0.360929f
C16 VDD1.t0 B 0.360929f
C17 VDD1.n0 B 3.2776f
C18 VDD1.t2 B 0.360929f
C19 VDD1.t1 B 0.360929f
C20 VDD1.n1 B 4.209549f
C21 VP.n0 B 0.030769f
C22 VP.t2 B 3.11438f
C23 VP.n1 B 0.046143f
C24 VP.n2 B 0.02334f
C25 VP.n3 B 0.025761f
C26 VP.t3 B 3.35387f
C27 VP.t0 B 3.35991f
C28 VP.n4 B 3.58342f
C29 VP.t1 B 3.11438f
C30 VP.n5 B 1.15855f
C31 VP.n6 B 1.45558f
C32 VP.n7 B 0.030769f
C33 VP.n8 B 0.02334f
C34 VP.n9 B 0.043281f
C35 VP.n10 B 0.046143f
C36 VP.n11 B 0.018851f
C37 VP.n12 B 0.02334f
C38 VP.n13 B 0.02334f
C39 VP.n14 B 0.02334f
C40 VP.n15 B 0.043281f
C41 VP.n16 B 0.025761f
C42 VP.n17 B 1.15855f
C43 VP.n18 B 0.043174f
C44 VTAIL.t7 B 2.36239f
C45 VTAIL.n0 B 0.315996f
C46 VTAIL.t0 B 2.36239f
C47 VTAIL.n1 B 0.381794f
C48 VTAIL.t2 B 2.36239f
C49 VTAIL.n2 B 1.44343f
C50 VTAIL.t6 B 2.36241f
C51 VTAIL.n3 B 1.44341f
C52 VTAIL.t5 B 2.36241f
C53 VTAIL.n4 B 0.381779f
C54 VTAIL.t3 B 2.36241f
C55 VTAIL.n5 B 0.381779f
C56 VTAIL.t1 B 2.36239f
C57 VTAIL.n6 B 1.44342f
C58 VTAIL.t4 B 2.36239f
C59 VTAIL.n7 B 1.37179f
C60 VDD2.t3 B 0.358229f
C61 VDD2.t0 B 0.358229f
C62 VDD2.n0 B 4.14911f
C63 VDD2.t2 B 0.358229f
C64 VDD2.t1 B 0.358229f
C65 VDD2.n1 B 3.25261f
C66 VDD2.n2 B 4.32464f
C67 VN.t0 B 3.2901f
C68 VN.t3 B 3.2842f
C69 VN.n0 B 2.07545f
C70 VN.t2 B 3.2901f
C71 VN.t1 B 3.2842f
C72 VN.n1 B 3.52095f
.ends

