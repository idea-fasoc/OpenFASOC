* NGSPICE file created from diff_pair_sample_1615.ext - technology: sky130A

.subckt diff_pair_sample_1615 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t7 VN.t0 VTAIL.t11 B.t6 sky130_fd_pr__nfet_01v8 ad=3.17955 pd=19.6 as=7.5153 ps=39.32 w=19.27 l=1.89
X1 VDD2.t6 VN.t1 VTAIL.t12 B.t2 sky130_fd_pr__nfet_01v8 ad=3.17955 pd=19.6 as=3.17955 ps=19.6 w=19.27 l=1.89
X2 VDD1.t7 VP.t0 VTAIL.t6 B.t6 sky130_fd_pr__nfet_01v8 ad=3.17955 pd=19.6 as=7.5153 ps=39.32 w=19.27 l=1.89
X3 VTAIL.t10 VN.t2 VDD2.t5 B.t4 sky130_fd_pr__nfet_01v8 ad=3.17955 pd=19.6 as=3.17955 ps=19.6 w=19.27 l=1.89
X4 B.t21 B.t19 B.t20 B.t9 sky130_fd_pr__nfet_01v8 ad=7.5153 pd=39.32 as=0 ps=0 w=19.27 l=1.89
X5 VDD1.t6 VP.t1 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=3.17955 pd=19.6 as=3.17955 ps=19.6 w=19.27 l=1.89
X6 VTAIL.t9 VN.t3 VDD2.t4 B.t0 sky130_fd_pr__nfet_01v8 ad=7.5153 pd=39.32 as=3.17955 ps=19.6 w=19.27 l=1.89
X7 B.t18 B.t16 B.t17 B.t13 sky130_fd_pr__nfet_01v8 ad=7.5153 pd=39.32 as=0 ps=0 w=19.27 l=1.89
X8 B.t15 B.t12 B.t14 B.t13 sky130_fd_pr__nfet_01v8 ad=7.5153 pd=39.32 as=0 ps=0 w=19.27 l=1.89
X9 VTAIL.t5 VP.t2 VDD1.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=7.5153 pd=39.32 as=3.17955 ps=19.6 w=19.27 l=1.89
X10 VDD1.t4 VP.t3 VTAIL.t7 B.t7 sky130_fd_pr__nfet_01v8 ad=3.17955 pd=19.6 as=7.5153 ps=39.32 w=19.27 l=1.89
X11 VTAIL.t3 VP.t4 VDD1.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=3.17955 pd=19.6 as=3.17955 ps=19.6 w=19.27 l=1.89
X12 VDD2.t3 VN.t4 VTAIL.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=3.17955 pd=19.6 as=7.5153 ps=39.32 w=19.27 l=1.89
X13 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=7.5153 pd=39.32 as=0 ps=0 w=19.27 l=1.89
X14 VTAIL.t14 VN.t5 VDD2.t2 B.t3 sky130_fd_pr__nfet_01v8 ad=3.17955 pd=19.6 as=3.17955 ps=19.6 w=19.27 l=1.89
X15 VTAIL.t15 VN.t6 VDD2.t1 B.t5 sky130_fd_pr__nfet_01v8 ad=7.5153 pd=39.32 as=3.17955 ps=19.6 w=19.27 l=1.89
X16 VTAIL.t0 VP.t5 VDD1.t2 B.t0 sky130_fd_pr__nfet_01v8 ad=7.5153 pd=39.32 as=3.17955 ps=19.6 w=19.27 l=1.89
X17 VDD2.t0 VN.t7 VTAIL.t13 B.t1 sky130_fd_pr__nfet_01v8 ad=3.17955 pd=19.6 as=3.17955 ps=19.6 w=19.27 l=1.89
X18 VDD1.t1 VP.t6 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=3.17955 pd=19.6 as=3.17955 ps=19.6 w=19.27 l=1.89
X19 VTAIL.t4 VP.t7 VDD1.t0 B.t4 sky130_fd_pr__nfet_01v8 ad=3.17955 pd=19.6 as=3.17955 ps=19.6 w=19.27 l=1.89
R0 VN.n5 VN.t6 280.058
R1 VN.n28 VN.t4 280.058
R2 VN.n6 VN.t1 245.719
R3 VN.n13 VN.t5 245.719
R4 VN.n21 VN.t0 245.719
R5 VN.n29 VN.t2 245.719
R6 VN.n36 VN.t7 245.719
R7 VN.n44 VN.t3 245.719
R8 VN.n22 VN.n21 181.852
R9 VN.n45 VN.n44 181.852
R10 VN.n43 VN.n23 161.3
R11 VN.n42 VN.n41 161.3
R12 VN.n40 VN.n24 161.3
R13 VN.n39 VN.n38 161.3
R14 VN.n37 VN.n25 161.3
R15 VN.n35 VN.n34 161.3
R16 VN.n33 VN.n26 161.3
R17 VN.n32 VN.n31 161.3
R18 VN.n30 VN.n27 161.3
R19 VN.n20 VN.n0 161.3
R20 VN.n19 VN.n18 161.3
R21 VN.n17 VN.n1 161.3
R22 VN.n16 VN.n15 161.3
R23 VN.n14 VN.n2 161.3
R24 VN.n12 VN.n11 161.3
R25 VN.n10 VN.n3 161.3
R26 VN.n9 VN.n8 161.3
R27 VN.n7 VN.n4 161.3
R28 VN.n8 VN.n3 56.5193
R29 VN.n31 VN.n26 56.5193
R30 VN VN.n45 53.3888
R31 VN.n6 VN.n5 52.0405
R32 VN.n29 VN.n28 52.0405
R33 VN.n15 VN.n1 43.4072
R34 VN.n38 VN.n24 43.4072
R35 VN.n19 VN.n1 37.5796
R36 VN.n42 VN.n24 37.5796
R37 VN.n8 VN.n7 24.4675
R38 VN.n12 VN.n3 24.4675
R39 VN.n15 VN.n14 24.4675
R40 VN.n20 VN.n19 24.4675
R41 VN.n31 VN.n30 24.4675
R42 VN.n38 VN.n37 24.4675
R43 VN.n35 VN.n26 24.4675
R44 VN.n43 VN.n42 24.4675
R45 VN.n7 VN.n6 17.6167
R46 VN.n13 VN.n12 17.6167
R47 VN.n30 VN.n29 17.6167
R48 VN.n36 VN.n35 17.6167
R49 VN.n28 VN.n27 12.2976
R50 VN.n5 VN.n4 12.2976
R51 VN.n14 VN.n13 6.85126
R52 VN.n37 VN.n36 6.85126
R53 VN.n21 VN.n20 3.91522
R54 VN.n44 VN.n43 3.91522
R55 VN.n45 VN.n23 0.189894
R56 VN.n41 VN.n23 0.189894
R57 VN.n41 VN.n40 0.189894
R58 VN.n40 VN.n39 0.189894
R59 VN.n39 VN.n25 0.189894
R60 VN.n34 VN.n25 0.189894
R61 VN.n34 VN.n33 0.189894
R62 VN.n33 VN.n32 0.189894
R63 VN.n32 VN.n27 0.189894
R64 VN.n9 VN.n4 0.189894
R65 VN.n10 VN.n9 0.189894
R66 VN.n11 VN.n10 0.189894
R67 VN.n11 VN.n2 0.189894
R68 VN.n16 VN.n2 0.189894
R69 VN.n17 VN.n16 0.189894
R70 VN.n18 VN.n17 0.189894
R71 VN.n18 VN.n0 0.189894
R72 VN.n22 VN.n0 0.189894
R73 VN VN.n22 0.0516364
R74 VTAIL.n11 VTAIL.t5 43.9902
R75 VTAIL.n10 VTAIL.t8 43.9902
R76 VTAIL.n7 VTAIL.t9 43.9902
R77 VTAIL.n15 VTAIL.t11 43.9899
R78 VTAIL.n2 VTAIL.t15 43.9899
R79 VTAIL.n3 VTAIL.t7 43.9899
R80 VTAIL.n6 VTAIL.t0 43.9899
R81 VTAIL.n14 VTAIL.t6 43.9899
R82 VTAIL.n13 VTAIL.n12 42.9627
R83 VTAIL.n9 VTAIL.n8 42.9627
R84 VTAIL.n1 VTAIL.n0 42.9626
R85 VTAIL.n5 VTAIL.n4 42.9626
R86 VTAIL.n15 VTAIL.n14 30.8927
R87 VTAIL.n7 VTAIL.n6 30.8927
R88 VTAIL.n9 VTAIL.n7 1.91429
R89 VTAIL.n10 VTAIL.n9 1.91429
R90 VTAIL.n13 VTAIL.n11 1.91429
R91 VTAIL.n14 VTAIL.n13 1.91429
R92 VTAIL.n6 VTAIL.n5 1.91429
R93 VTAIL.n5 VTAIL.n3 1.91429
R94 VTAIL.n2 VTAIL.n1 1.91429
R95 VTAIL VTAIL.n15 1.8561
R96 VTAIL.n0 VTAIL.t12 1.028
R97 VTAIL.n0 VTAIL.t14 1.028
R98 VTAIL.n4 VTAIL.t1 1.028
R99 VTAIL.n4 VTAIL.t4 1.028
R100 VTAIL.n12 VTAIL.t2 1.028
R101 VTAIL.n12 VTAIL.t3 1.028
R102 VTAIL.n8 VTAIL.t13 1.028
R103 VTAIL.n8 VTAIL.t10 1.028
R104 VTAIL.n11 VTAIL.n10 0.470328
R105 VTAIL.n3 VTAIL.n2 0.470328
R106 VTAIL VTAIL.n1 0.0586897
R107 VDD2.n2 VDD2.n1 60.5429
R108 VDD2.n2 VDD2.n0 60.5429
R109 VDD2 VDD2.n5 60.54
R110 VDD2.n4 VDD2.n3 59.6414
R111 VDD2.n4 VDD2.n2 48.9394
R112 VDD2.n5 VDD2.t5 1.028
R113 VDD2.n5 VDD2.t3 1.028
R114 VDD2.n3 VDD2.t4 1.028
R115 VDD2.n3 VDD2.t0 1.028
R116 VDD2.n1 VDD2.t2 1.028
R117 VDD2.n1 VDD2.t7 1.028
R118 VDD2.n0 VDD2.t1 1.028
R119 VDD2.n0 VDD2.t6 1.028
R120 VDD2 VDD2.n4 1.01559
R121 B.n1015 B.n1014 585
R122 B.n417 B.n144 585
R123 B.n416 B.n415 585
R124 B.n414 B.n413 585
R125 B.n412 B.n411 585
R126 B.n410 B.n409 585
R127 B.n408 B.n407 585
R128 B.n406 B.n405 585
R129 B.n404 B.n403 585
R130 B.n402 B.n401 585
R131 B.n400 B.n399 585
R132 B.n398 B.n397 585
R133 B.n396 B.n395 585
R134 B.n394 B.n393 585
R135 B.n392 B.n391 585
R136 B.n390 B.n389 585
R137 B.n388 B.n387 585
R138 B.n386 B.n385 585
R139 B.n384 B.n383 585
R140 B.n382 B.n381 585
R141 B.n380 B.n379 585
R142 B.n378 B.n377 585
R143 B.n376 B.n375 585
R144 B.n374 B.n373 585
R145 B.n372 B.n371 585
R146 B.n370 B.n369 585
R147 B.n368 B.n367 585
R148 B.n366 B.n365 585
R149 B.n364 B.n363 585
R150 B.n362 B.n361 585
R151 B.n360 B.n359 585
R152 B.n358 B.n357 585
R153 B.n356 B.n355 585
R154 B.n354 B.n353 585
R155 B.n352 B.n351 585
R156 B.n350 B.n349 585
R157 B.n348 B.n347 585
R158 B.n346 B.n345 585
R159 B.n344 B.n343 585
R160 B.n342 B.n341 585
R161 B.n340 B.n339 585
R162 B.n338 B.n337 585
R163 B.n336 B.n335 585
R164 B.n334 B.n333 585
R165 B.n332 B.n331 585
R166 B.n330 B.n329 585
R167 B.n328 B.n327 585
R168 B.n326 B.n325 585
R169 B.n324 B.n323 585
R170 B.n322 B.n321 585
R171 B.n320 B.n319 585
R172 B.n318 B.n317 585
R173 B.n316 B.n315 585
R174 B.n314 B.n313 585
R175 B.n312 B.n311 585
R176 B.n310 B.n309 585
R177 B.n308 B.n307 585
R178 B.n306 B.n305 585
R179 B.n304 B.n303 585
R180 B.n302 B.n301 585
R181 B.n300 B.n299 585
R182 B.n298 B.n297 585
R183 B.n296 B.n295 585
R184 B.n293 B.n292 585
R185 B.n291 B.n290 585
R186 B.n289 B.n288 585
R187 B.n287 B.n286 585
R188 B.n285 B.n284 585
R189 B.n283 B.n282 585
R190 B.n281 B.n280 585
R191 B.n279 B.n278 585
R192 B.n277 B.n276 585
R193 B.n275 B.n274 585
R194 B.n272 B.n271 585
R195 B.n270 B.n269 585
R196 B.n268 B.n267 585
R197 B.n266 B.n265 585
R198 B.n264 B.n263 585
R199 B.n262 B.n261 585
R200 B.n260 B.n259 585
R201 B.n258 B.n257 585
R202 B.n256 B.n255 585
R203 B.n254 B.n253 585
R204 B.n252 B.n251 585
R205 B.n250 B.n249 585
R206 B.n248 B.n247 585
R207 B.n246 B.n245 585
R208 B.n244 B.n243 585
R209 B.n242 B.n241 585
R210 B.n240 B.n239 585
R211 B.n238 B.n237 585
R212 B.n236 B.n235 585
R213 B.n234 B.n233 585
R214 B.n232 B.n231 585
R215 B.n230 B.n229 585
R216 B.n228 B.n227 585
R217 B.n226 B.n225 585
R218 B.n224 B.n223 585
R219 B.n222 B.n221 585
R220 B.n220 B.n219 585
R221 B.n218 B.n217 585
R222 B.n216 B.n215 585
R223 B.n214 B.n213 585
R224 B.n212 B.n211 585
R225 B.n210 B.n209 585
R226 B.n208 B.n207 585
R227 B.n206 B.n205 585
R228 B.n204 B.n203 585
R229 B.n202 B.n201 585
R230 B.n200 B.n199 585
R231 B.n198 B.n197 585
R232 B.n196 B.n195 585
R233 B.n194 B.n193 585
R234 B.n192 B.n191 585
R235 B.n190 B.n189 585
R236 B.n188 B.n187 585
R237 B.n186 B.n185 585
R238 B.n184 B.n183 585
R239 B.n182 B.n181 585
R240 B.n180 B.n179 585
R241 B.n178 B.n177 585
R242 B.n176 B.n175 585
R243 B.n174 B.n173 585
R244 B.n172 B.n171 585
R245 B.n170 B.n169 585
R246 B.n168 B.n167 585
R247 B.n166 B.n165 585
R248 B.n164 B.n163 585
R249 B.n162 B.n161 585
R250 B.n160 B.n159 585
R251 B.n158 B.n157 585
R252 B.n156 B.n155 585
R253 B.n154 B.n153 585
R254 B.n152 B.n151 585
R255 B.n150 B.n149 585
R256 B.n75 B.n74 585
R257 B.n1013 B.n76 585
R258 B.n1018 B.n76 585
R259 B.n1012 B.n1011 585
R260 B.n1011 B.n72 585
R261 B.n1010 B.n71 585
R262 B.n1024 B.n71 585
R263 B.n1009 B.n70 585
R264 B.n1025 B.n70 585
R265 B.n1008 B.n69 585
R266 B.n1026 B.n69 585
R267 B.n1007 B.n1006 585
R268 B.n1006 B.n65 585
R269 B.n1005 B.n64 585
R270 B.n1032 B.n64 585
R271 B.n1004 B.n63 585
R272 B.n1033 B.n63 585
R273 B.n1003 B.n62 585
R274 B.n1034 B.n62 585
R275 B.n1002 B.n1001 585
R276 B.n1001 B.n58 585
R277 B.n1000 B.n57 585
R278 B.n1040 B.n57 585
R279 B.n999 B.n56 585
R280 B.n1041 B.n56 585
R281 B.n998 B.n55 585
R282 B.n1042 B.n55 585
R283 B.n997 B.n996 585
R284 B.n996 B.n51 585
R285 B.n995 B.n50 585
R286 B.n1048 B.n50 585
R287 B.n994 B.n49 585
R288 B.n1049 B.n49 585
R289 B.n993 B.n48 585
R290 B.n1050 B.n48 585
R291 B.n992 B.n991 585
R292 B.n991 B.n44 585
R293 B.n990 B.n43 585
R294 B.n1056 B.n43 585
R295 B.n989 B.n42 585
R296 B.n1057 B.n42 585
R297 B.n988 B.n41 585
R298 B.n1058 B.n41 585
R299 B.n987 B.n986 585
R300 B.n986 B.n37 585
R301 B.n985 B.n36 585
R302 B.n1064 B.n36 585
R303 B.n984 B.n35 585
R304 B.n1065 B.n35 585
R305 B.n983 B.n34 585
R306 B.n1066 B.n34 585
R307 B.n982 B.n981 585
R308 B.n981 B.n30 585
R309 B.n980 B.n29 585
R310 B.n1072 B.n29 585
R311 B.n979 B.n28 585
R312 B.n1073 B.n28 585
R313 B.n978 B.n27 585
R314 B.n1074 B.n27 585
R315 B.n977 B.n976 585
R316 B.n976 B.n26 585
R317 B.n975 B.n22 585
R318 B.n1080 B.n22 585
R319 B.n974 B.n21 585
R320 B.n1081 B.n21 585
R321 B.n973 B.n20 585
R322 B.n1082 B.n20 585
R323 B.n972 B.n971 585
R324 B.n971 B.n16 585
R325 B.n970 B.n15 585
R326 B.n1088 B.n15 585
R327 B.n969 B.n14 585
R328 B.n1089 B.n14 585
R329 B.n968 B.n13 585
R330 B.n1090 B.n13 585
R331 B.n967 B.n966 585
R332 B.n966 B.n12 585
R333 B.n965 B.n964 585
R334 B.n965 B.n8 585
R335 B.n963 B.n7 585
R336 B.n1097 B.n7 585
R337 B.n962 B.n6 585
R338 B.n1098 B.n6 585
R339 B.n961 B.n5 585
R340 B.n1099 B.n5 585
R341 B.n960 B.n959 585
R342 B.n959 B.n4 585
R343 B.n958 B.n418 585
R344 B.n958 B.n957 585
R345 B.n948 B.n419 585
R346 B.n420 B.n419 585
R347 B.n950 B.n949 585
R348 B.n951 B.n950 585
R349 B.n947 B.n424 585
R350 B.n428 B.n424 585
R351 B.n946 B.n945 585
R352 B.n945 B.n944 585
R353 B.n426 B.n425 585
R354 B.n427 B.n426 585
R355 B.n937 B.n936 585
R356 B.n938 B.n937 585
R357 B.n935 B.n433 585
R358 B.n433 B.n432 585
R359 B.n934 B.n933 585
R360 B.n933 B.n932 585
R361 B.n435 B.n434 585
R362 B.n925 B.n435 585
R363 B.n924 B.n923 585
R364 B.n926 B.n924 585
R365 B.n922 B.n440 585
R366 B.n440 B.n439 585
R367 B.n921 B.n920 585
R368 B.n920 B.n919 585
R369 B.n442 B.n441 585
R370 B.n443 B.n442 585
R371 B.n912 B.n911 585
R372 B.n913 B.n912 585
R373 B.n910 B.n448 585
R374 B.n448 B.n447 585
R375 B.n909 B.n908 585
R376 B.n908 B.n907 585
R377 B.n450 B.n449 585
R378 B.n451 B.n450 585
R379 B.n900 B.n899 585
R380 B.n901 B.n900 585
R381 B.n898 B.n456 585
R382 B.n456 B.n455 585
R383 B.n897 B.n896 585
R384 B.n896 B.n895 585
R385 B.n458 B.n457 585
R386 B.n459 B.n458 585
R387 B.n888 B.n887 585
R388 B.n889 B.n888 585
R389 B.n886 B.n464 585
R390 B.n464 B.n463 585
R391 B.n885 B.n884 585
R392 B.n884 B.n883 585
R393 B.n466 B.n465 585
R394 B.n467 B.n466 585
R395 B.n876 B.n875 585
R396 B.n877 B.n876 585
R397 B.n874 B.n472 585
R398 B.n472 B.n471 585
R399 B.n873 B.n872 585
R400 B.n872 B.n871 585
R401 B.n474 B.n473 585
R402 B.n475 B.n474 585
R403 B.n864 B.n863 585
R404 B.n865 B.n864 585
R405 B.n862 B.n480 585
R406 B.n480 B.n479 585
R407 B.n861 B.n860 585
R408 B.n860 B.n859 585
R409 B.n482 B.n481 585
R410 B.n483 B.n482 585
R411 B.n852 B.n851 585
R412 B.n853 B.n852 585
R413 B.n850 B.n488 585
R414 B.n488 B.n487 585
R415 B.n849 B.n848 585
R416 B.n848 B.n847 585
R417 B.n490 B.n489 585
R418 B.n491 B.n490 585
R419 B.n840 B.n839 585
R420 B.n841 B.n840 585
R421 B.n494 B.n493 585
R422 B.n571 B.n570 585
R423 B.n572 B.n568 585
R424 B.n568 B.n495 585
R425 B.n574 B.n573 585
R426 B.n576 B.n567 585
R427 B.n579 B.n578 585
R428 B.n580 B.n566 585
R429 B.n582 B.n581 585
R430 B.n584 B.n565 585
R431 B.n587 B.n586 585
R432 B.n588 B.n564 585
R433 B.n590 B.n589 585
R434 B.n592 B.n563 585
R435 B.n595 B.n594 585
R436 B.n596 B.n562 585
R437 B.n598 B.n597 585
R438 B.n600 B.n561 585
R439 B.n603 B.n602 585
R440 B.n604 B.n560 585
R441 B.n606 B.n605 585
R442 B.n608 B.n559 585
R443 B.n611 B.n610 585
R444 B.n612 B.n558 585
R445 B.n614 B.n613 585
R446 B.n616 B.n557 585
R447 B.n619 B.n618 585
R448 B.n620 B.n556 585
R449 B.n622 B.n621 585
R450 B.n624 B.n555 585
R451 B.n627 B.n626 585
R452 B.n628 B.n554 585
R453 B.n630 B.n629 585
R454 B.n632 B.n553 585
R455 B.n635 B.n634 585
R456 B.n636 B.n552 585
R457 B.n638 B.n637 585
R458 B.n640 B.n551 585
R459 B.n643 B.n642 585
R460 B.n644 B.n550 585
R461 B.n646 B.n645 585
R462 B.n648 B.n549 585
R463 B.n651 B.n650 585
R464 B.n652 B.n548 585
R465 B.n654 B.n653 585
R466 B.n656 B.n547 585
R467 B.n659 B.n658 585
R468 B.n660 B.n546 585
R469 B.n662 B.n661 585
R470 B.n664 B.n545 585
R471 B.n667 B.n666 585
R472 B.n668 B.n544 585
R473 B.n670 B.n669 585
R474 B.n672 B.n543 585
R475 B.n675 B.n674 585
R476 B.n676 B.n542 585
R477 B.n678 B.n677 585
R478 B.n680 B.n541 585
R479 B.n683 B.n682 585
R480 B.n684 B.n540 585
R481 B.n686 B.n685 585
R482 B.n688 B.n539 585
R483 B.n691 B.n690 585
R484 B.n692 B.n536 585
R485 B.n695 B.n694 585
R486 B.n697 B.n535 585
R487 B.n700 B.n699 585
R488 B.n701 B.n534 585
R489 B.n703 B.n702 585
R490 B.n705 B.n533 585
R491 B.n708 B.n707 585
R492 B.n709 B.n532 585
R493 B.n711 B.n710 585
R494 B.n713 B.n531 585
R495 B.n716 B.n715 585
R496 B.n717 B.n527 585
R497 B.n719 B.n718 585
R498 B.n721 B.n526 585
R499 B.n724 B.n723 585
R500 B.n725 B.n525 585
R501 B.n727 B.n726 585
R502 B.n729 B.n524 585
R503 B.n732 B.n731 585
R504 B.n733 B.n523 585
R505 B.n735 B.n734 585
R506 B.n737 B.n522 585
R507 B.n740 B.n739 585
R508 B.n741 B.n521 585
R509 B.n743 B.n742 585
R510 B.n745 B.n520 585
R511 B.n748 B.n747 585
R512 B.n749 B.n519 585
R513 B.n751 B.n750 585
R514 B.n753 B.n518 585
R515 B.n756 B.n755 585
R516 B.n757 B.n517 585
R517 B.n759 B.n758 585
R518 B.n761 B.n516 585
R519 B.n764 B.n763 585
R520 B.n765 B.n515 585
R521 B.n767 B.n766 585
R522 B.n769 B.n514 585
R523 B.n772 B.n771 585
R524 B.n773 B.n513 585
R525 B.n775 B.n774 585
R526 B.n777 B.n512 585
R527 B.n780 B.n779 585
R528 B.n781 B.n511 585
R529 B.n783 B.n782 585
R530 B.n785 B.n510 585
R531 B.n788 B.n787 585
R532 B.n789 B.n509 585
R533 B.n791 B.n790 585
R534 B.n793 B.n508 585
R535 B.n796 B.n795 585
R536 B.n797 B.n507 585
R537 B.n799 B.n798 585
R538 B.n801 B.n506 585
R539 B.n804 B.n803 585
R540 B.n805 B.n505 585
R541 B.n807 B.n806 585
R542 B.n809 B.n504 585
R543 B.n812 B.n811 585
R544 B.n813 B.n503 585
R545 B.n815 B.n814 585
R546 B.n817 B.n502 585
R547 B.n820 B.n819 585
R548 B.n821 B.n501 585
R549 B.n823 B.n822 585
R550 B.n825 B.n500 585
R551 B.n828 B.n827 585
R552 B.n829 B.n499 585
R553 B.n831 B.n830 585
R554 B.n833 B.n498 585
R555 B.n834 B.n497 585
R556 B.n837 B.n836 585
R557 B.n838 B.n496 585
R558 B.n496 B.n495 585
R559 B.n843 B.n842 585
R560 B.n842 B.n841 585
R561 B.n844 B.n492 585
R562 B.n492 B.n491 585
R563 B.n846 B.n845 585
R564 B.n847 B.n846 585
R565 B.n486 B.n485 585
R566 B.n487 B.n486 585
R567 B.n855 B.n854 585
R568 B.n854 B.n853 585
R569 B.n856 B.n484 585
R570 B.n484 B.n483 585
R571 B.n858 B.n857 585
R572 B.n859 B.n858 585
R573 B.n478 B.n477 585
R574 B.n479 B.n478 585
R575 B.n867 B.n866 585
R576 B.n866 B.n865 585
R577 B.n868 B.n476 585
R578 B.n476 B.n475 585
R579 B.n870 B.n869 585
R580 B.n871 B.n870 585
R581 B.n470 B.n469 585
R582 B.n471 B.n470 585
R583 B.n879 B.n878 585
R584 B.n878 B.n877 585
R585 B.n880 B.n468 585
R586 B.n468 B.n467 585
R587 B.n882 B.n881 585
R588 B.n883 B.n882 585
R589 B.n462 B.n461 585
R590 B.n463 B.n462 585
R591 B.n891 B.n890 585
R592 B.n890 B.n889 585
R593 B.n892 B.n460 585
R594 B.n460 B.n459 585
R595 B.n894 B.n893 585
R596 B.n895 B.n894 585
R597 B.n454 B.n453 585
R598 B.n455 B.n454 585
R599 B.n903 B.n902 585
R600 B.n902 B.n901 585
R601 B.n904 B.n452 585
R602 B.n452 B.n451 585
R603 B.n906 B.n905 585
R604 B.n907 B.n906 585
R605 B.n446 B.n445 585
R606 B.n447 B.n446 585
R607 B.n915 B.n914 585
R608 B.n914 B.n913 585
R609 B.n916 B.n444 585
R610 B.n444 B.n443 585
R611 B.n918 B.n917 585
R612 B.n919 B.n918 585
R613 B.n438 B.n437 585
R614 B.n439 B.n438 585
R615 B.n928 B.n927 585
R616 B.n927 B.n926 585
R617 B.n929 B.n436 585
R618 B.n925 B.n436 585
R619 B.n931 B.n930 585
R620 B.n932 B.n931 585
R621 B.n431 B.n430 585
R622 B.n432 B.n431 585
R623 B.n940 B.n939 585
R624 B.n939 B.n938 585
R625 B.n941 B.n429 585
R626 B.n429 B.n427 585
R627 B.n943 B.n942 585
R628 B.n944 B.n943 585
R629 B.n423 B.n422 585
R630 B.n428 B.n423 585
R631 B.n953 B.n952 585
R632 B.n952 B.n951 585
R633 B.n954 B.n421 585
R634 B.n421 B.n420 585
R635 B.n956 B.n955 585
R636 B.n957 B.n956 585
R637 B.n3 B.n0 585
R638 B.n4 B.n3 585
R639 B.n1096 B.n1 585
R640 B.n1097 B.n1096 585
R641 B.n1095 B.n1094 585
R642 B.n1095 B.n8 585
R643 B.n1093 B.n9 585
R644 B.n12 B.n9 585
R645 B.n1092 B.n1091 585
R646 B.n1091 B.n1090 585
R647 B.n11 B.n10 585
R648 B.n1089 B.n11 585
R649 B.n1087 B.n1086 585
R650 B.n1088 B.n1087 585
R651 B.n1085 B.n17 585
R652 B.n17 B.n16 585
R653 B.n1084 B.n1083 585
R654 B.n1083 B.n1082 585
R655 B.n19 B.n18 585
R656 B.n1081 B.n19 585
R657 B.n1079 B.n1078 585
R658 B.n1080 B.n1079 585
R659 B.n1077 B.n23 585
R660 B.n26 B.n23 585
R661 B.n1076 B.n1075 585
R662 B.n1075 B.n1074 585
R663 B.n25 B.n24 585
R664 B.n1073 B.n25 585
R665 B.n1071 B.n1070 585
R666 B.n1072 B.n1071 585
R667 B.n1069 B.n31 585
R668 B.n31 B.n30 585
R669 B.n1068 B.n1067 585
R670 B.n1067 B.n1066 585
R671 B.n33 B.n32 585
R672 B.n1065 B.n33 585
R673 B.n1063 B.n1062 585
R674 B.n1064 B.n1063 585
R675 B.n1061 B.n38 585
R676 B.n38 B.n37 585
R677 B.n1060 B.n1059 585
R678 B.n1059 B.n1058 585
R679 B.n40 B.n39 585
R680 B.n1057 B.n40 585
R681 B.n1055 B.n1054 585
R682 B.n1056 B.n1055 585
R683 B.n1053 B.n45 585
R684 B.n45 B.n44 585
R685 B.n1052 B.n1051 585
R686 B.n1051 B.n1050 585
R687 B.n47 B.n46 585
R688 B.n1049 B.n47 585
R689 B.n1047 B.n1046 585
R690 B.n1048 B.n1047 585
R691 B.n1045 B.n52 585
R692 B.n52 B.n51 585
R693 B.n1044 B.n1043 585
R694 B.n1043 B.n1042 585
R695 B.n54 B.n53 585
R696 B.n1041 B.n54 585
R697 B.n1039 B.n1038 585
R698 B.n1040 B.n1039 585
R699 B.n1037 B.n59 585
R700 B.n59 B.n58 585
R701 B.n1036 B.n1035 585
R702 B.n1035 B.n1034 585
R703 B.n61 B.n60 585
R704 B.n1033 B.n61 585
R705 B.n1031 B.n1030 585
R706 B.n1032 B.n1031 585
R707 B.n1029 B.n66 585
R708 B.n66 B.n65 585
R709 B.n1028 B.n1027 585
R710 B.n1027 B.n1026 585
R711 B.n68 B.n67 585
R712 B.n1025 B.n68 585
R713 B.n1023 B.n1022 585
R714 B.n1024 B.n1023 585
R715 B.n1021 B.n73 585
R716 B.n73 B.n72 585
R717 B.n1020 B.n1019 585
R718 B.n1019 B.n1018 585
R719 B.n1100 B.n1099 585
R720 B.n1098 B.n2 585
R721 B.n1019 B.n75 506.916
R722 B.n1015 B.n76 506.916
R723 B.n840 B.n496 506.916
R724 B.n842 B.n494 506.916
R725 B.n147 B.t19 452.365
R726 B.n145 B.t8 452.365
R727 B.n528 B.t12 452.365
R728 B.n537 B.t16 452.365
R729 B.n1017 B.n1016 256.663
R730 B.n1017 B.n143 256.663
R731 B.n1017 B.n142 256.663
R732 B.n1017 B.n141 256.663
R733 B.n1017 B.n140 256.663
R734 B.n1017 B.n139 256.663
R735 B.n1017 B.n138 256.663
R736 B.n1017 B.n137 256.663
R737 B.n1017 B.n136 256.663
R738 B.n1017 B.n135 256.663
R739 B.n1017 B.n134 256.663
R740 B.n1017 B.n133 256.663
R741 B.n1017 B.n132 256.663
R742 B.n1017 B.n131 256.663
R743 B.n1017 B.n130 256.663
R744 B.n1017 B.n129 256.663
R745 B.n1017 B.n128 256.663
R746 B.n1017 B.n127 256.663
R747 B.n1017 B.n126 256.663
R748 B.n1017 B.n125 256.663
R749 B.n1017 B.n124 256.663
R750 B.n1017 B.n123 256.663
R751 B.n1017 B.n122 256.663
R752 B.n1017 B.n121 256.663
R753 B.n1017 B.n120 256.663
R754 B.n1017 B.n119 256.663
R755 B.n1017 B.n118 256.663
R756 B.n1017 B.n117 256.663
R757 B.n1017 B.n116 256.663
R758 B.n1017 B.n115 256.663
R759 B.n1017 B.n114 256.663
R760 B.n1017 B.n113 256.663
R761 B.n1017 B.n112 256.663
R762 B.n1017 B.n111 256.663
R763 B.n1017 B.n110 256.663
R764 B.n1017 B.n109 256.663
R765 B.n1017 B.n108 256.663
R766 B.n1017 B.n107 256.663
R767 B.n1017 B.n106 256.663
R768 B.n1017 B.n105 256.663
R769 B.n1017 B.n104 256.663
R770 B.n1017 B.n103 256.663
R771 B.n1017 B.n102 256.663
R772 B.n1017 B.n101 256.663
R773 B.n1017 B.n100 256.663
R774 B.n1017 B.n99 256.663
R775 B.n1017 B.n98 256.663
R776 B.n1017 B.n97 256.663
R777 B.n1017 B.n96 256.663
R778 B.n1017 B.n95 256.663
R779 B.n1017 B.n94 256.663
R780 B.n1017 B.n93 256.663
R781 B.n1017 B.n92 256.663
R782 B.n1017 B.n91 256.663
R783 B.n1017 B.n90 256.663
R784 B.n1017 B.n89 256.663
R785 B.n1017 B.n88 256.663
R786 B.n1017 B.n87 256.663
R787 B.n1017 B.n86 256.663
R788 B.n1017 B.n85 256.663
R789 B.n1017 B.n84 256.663
R790 B.n1017 B.n83 256.663
R791 B.n1017 B.n82 256.663
R792 B.n1017 B.n81 256.663
R793 B.n1017 B.n80 256.663
R794 B.n1017 B.n79 256.663
R795 B.n1017 B.n78 256.663
R796 B.n1017 B.n77 256.663
R797 B.n569 B.n495 256.663
R798 B.n575 B.n495 256.663
R799 B.n577 B.n495 256.663
R800 B.n583 B.n495 256.663
R801 B.n585 B.n495 256.663
R802 B.n591 B.n495 256.663
R803 B.n593 B.n495 256.663
R804 B.n599 B.n495 256.663
R805 B.n601 B.n495 256.663
R806 B.n607 B.n495 256.663
R807 B.n609 B.n495 256.663
R808 B.n615 B.n495 256.663
R809 B.n617 B.n495 256.663
R810 B.n623 B.n495 256.663
R811 B.n625 B.n495 256.663
R812 B.n631 B.n495 256.663
R813 B.n633 B.n495 256.663
R814 B.n639 B.n495 256.663
R815 B.n641 B.n495 256.663
R816 B.n647 B.n495 256.663
R817 B.n649 B.n495 256.663
R818 B.n655 B.n495 256.663
R819 B.n657 B.n495 256.663
R820 B.n663 B.n495 256.663
R821 B.n665 B.n495 256.663
R822 B.n671 B.n495 256.663
R823 B.n673 B.n495 256.663
R824 B.n679 B.n495 256.663
R825 B.n681 B.n495 256.663
R826 B.n687 B.n495 256.663
R827 B.n689 B.n495 256.663
R828 B.n696 B.n495 256.663
R829 B.n698 B.n495 256.663
R830 B.n704 B.n495 256.663
R831 B.n706 B.n495 256.663
R832 B.n712 B.n495 256.663
R833 B.n714 B.n495 256.663
R834 B.n720 B.n495 256.663
R835 B.n722 B.n495 256.663
R836 B.n728 B.n495 256.663
R837 B.n730 B.n495 256.663
R838 B.n736 B.n495 256.663
R839 B.n738 B.n495 256.663
R840 B.n744 B.n495 256.663
R841 B.n746 B.n495 256.663
R842 B.n752 B.n495 256.663
R843 B.n754 B.n495 256.663
R844 B.n760 B.n495 256.663
R845 B.n762 B.n495 256.663
R846 B.n768 B.n495 256.663
R847 B.n770 B.n495 256.663
R848 B.n776 B.n495 256.663
R849 B.n778 B.n495 256.663
R850 B.n784 B.n495 256.663
R851 B.n786 B.n495 256.663
R852 B.n792 B.n495 256.663
R853 B.n794 B.n495 256.663
R854 B.n800 B.n495 256.663
R855 B.n802 B.n495 256.663
R856 B.n808 B.n495 256.663
R857 B.n810 B.n495 256.663
R858 B.n816 B.n495 256.663
R859 B.n818 B.n495 256.663
R860 B.n824 B.n495 256.663
R861 B.n826 B.n495 256.663
R862 B.n832 B.n495 256.663
R863 B.n835 B.n495 256.663
R864 B.n1102 B.n1101 256.663
R865 B.n151 B.n150 163.367
R866 B.n155 B.n154 163.367
R867 B.n159 B.n158 163.367
R868 B.n163 B.n162 163.367
R869 B.n167 B.n166 163.367
R870 B.n171 B.n170 163.367
R871 B.n175 B.n174 163.367
R872 B.n179 B.n178 163.367
R873 B.n183 B.n182 163.367
R874 B.n187 B.n186 163.367
R875 B.n191 B.n190 163.367
R876 B.n195 B.n194 163.367
R877 B.n199 B.n198 163.367
R878 B.n203 B.n202 163.367
R879 B.n207 B.n206 163.367
R880 B.n211 B.n210 163.367
R881 B.n215 B.n214 163.367
R882 B.n219 B.n218 163.367
R883 B.n223 B.n222 163.367
R884 B.n227 B.n226 163.367
R885 B.n231 B.n230 163.367
R886 B.n235 B.n234 163.367
R887 B.n239 B.n238 163.367
R888 B.n243 B.n242 163.367
R889 B.n247 B.n246 163.367
R890 B.n251 B.n250 163.367
R891 B.n255 B.n254 163.367
R892 B.n259 B.n258 163.367
R893 B.n263 B.n262 163.367
R894 B.n267 B.n266 163.367
R895 B.n271 B.n270 163.367
R896 B.n276 B.n275 163.367
R897 B.n280 B.n279 163.367
R898 B.n284 B.n283 163.367
R899 B.n288 B.n287 163.367
R900 B.n292 B.n291 163.367
R901 B.n297 B.n296 163.367
R902 B.n301 B.n300 163.367
R903 B.n305 B.n304 163.367
R904 B.n309 B.n308 163.367
R905 B.n313 B.n312 163.367
R906 B.n317 B.n316 163.367
R907 B.n321 B.n320 163.367
R908 B.n325 B.n324 163.367
R909 B.n329 B.n328 163.367
R910 B.n333 B.n332 163.367
R911 B.n337 B.n336 163.367
R912 B.n341 B.n340 163.367
R913 B.n345 B.n344 163.367
R914 B.n349 B.n348 163.367
R915 B.n353 B.n352 163.367
R916 B.n357 B.n356 163.367
R917 B.n361 B.n360 163.367
R918 B.n365 B.n364 163.367
R919 B.n369 B.n368 163.367
R920 B.n373 B.n372 163.367
R921 B.n377 B.n376 163.367
R922 B.n381 B.n380 163.367
R923 B.n385 B.n384 163.367
R924 B.n389 B.n388 163.367
R925 B.n393 B.n392 163.367
R926 B.n397 B.n396 163.367
R927 B.n401 B.n400 163.367
R928 B.n405 B.n404 163.367
R929 B.n409 B.n408 163.367
R930 B.n413 B.n412 163.367
R931 B.n415 B.n144 163.367
R932 B.n840 B.n490 163.367
R933 B.n848 B.n490 163.367
R934 B.n848 B.n488 163.367
R935 B.n852 B.n488 163.367
R936 B.n852 B.n482 163.367
R937 B.n860 B.n482 163.367
R938 B.n860 B.n480 163.367
R939 B.n864 B.n480 163.367
R940 B.n864 B.n474 163.367
R941 B.n872 B.n474 163.367
R942 B.n872 B.n472 163.367
R943 B.n876 B.n472 163.367
R944 B.n876 B.n466 163.367
R945 B.n884 B.n466 163.367
R946 B.n884 B.n464 163.367
R947 B.n888 B.n464 163.367
R948 B.n888 B.n458 163.367
R949 B.n896 B.n458 163.367
R950 B.n896 B.n456 163.367
R951 B.n900 B.n456 163.367
R952 B.n900 B.n450 163.367
R953 B.n908 B.n450 163.367
R954 B.n908 B.n448 163.367
R955 B.n912 B.n448 163.367
R956 B.n912 B.n442 163.367
R957 B.n920 B.n442 163.367
R958 B.n920 B.n440 163.367
R959 B.n924 B.n440 163.367
R960 B.n924 B.n435 163.367
R961 B.n933 B.n435 163.367
R962 B.n933 B.n433 163.367
R963 B.n937 B.n433 163.367
R964 B.n937 B.n426 163.367
R965 B.n945 B.n426 163.367
R966 B.n945 B.n424 163.367
R967 B.n950 B.n424 163.367
R968 B.n950 B.n419 163.367
R969 B.n958 B.n419 163.367
R970 B.n959 B.n958 163.367
R971 B.n959 B.n5 163.367
R972 B.n6 B.n5 163.367
R973 B.n7 B.n6 163.367
R974 B.n965 B.n7 163.367
R975 B.n966 B.n965 163.367
R976 B.n966 B.n13 163.367
R977 B.n14 B.n13 163.367
R978 B.n15 B.n14 163.367
R979 B.n971 B.n15 163.367
R980 B.n971 B.n20 163.367
R981 B.n21 B.n20 163.367
R982 B.n22 B.n21 163.367
R983 B.n976 B.n22 163.367
R984 B.n976 B.n27 163.367
R985 B.n28 B.n27 163.367
R986 B.n29 B.n28 163.367
R987 B.n981 B.n29 163.367
R988 B.n981 B.n34 163.367
R989 B.n35 B.n34 163.367
R990 B.n36 B.n35 163.367
R991 B.n986 B.n36 163.367
R992 B.n986 B.n41 163.367
R993 B.n42 B.n41 163.367
R994 B.n43 B.n42 163.367
R995 B.n991 B.n43 163.367
R996 B.n991 B.n48 163.367
R997 B.n49 B.n48 163.367
R998 B.n50 B.n49 163.367
R999 B.n996 B.n50 163.367
R1000 B.n996 B.n55 163.367
R1001 B.n56 B.n55 163.367
R1002 B.n57 B.n56 163.367
R1003 B.n1001 B.n57 163.367
R1004 B.n1001 B.n62 163.367
R1005 B.n63 B.n62 163.367
R1006 B.n64 B.n63 163.367
R1007 B.n1006 B.n64 163.367
R1008 B.n1006 B.n69 163.367
R1009 B.n70 B.n69 163.367
R1010 B.n71 B.n70 163.367
R1011 B.n1011 B.n71 163.367
R1012 B.n1011 B.n76 163.367
R1013 B.n570 B.n568 163.367
R1014 B.n574 B.n568 163.367
R1015 B.n578 B.n576 163.367
R1016 B.n582 B.n566 163.367
R1017 B.n586 B.n584 163.367
R1018 B.n590 B.n564 163.367
R1019 B.n594 B.n592 163.367
R1020 B.n598 B.n562 163.367
R1021 B.n602 B.n600 163.367
R1022 B.n606 B.n560 163.367
R1023 B.n610 B.n608 163.367
R1024 B.n614 B.n558 163.367
R1025 B.n618 B.n616 163.367
R1026 B.n622 B.n556 163.367
R1027 B.n626 B.n624 163.367
R1028 B.n630 B.n554 163.367
R1029 B.n634 B.n632 163.367
R1030 B.n638 B.n552 163.367
R1031 B.n642 B.n640 163.367
R1032 B.n646 B.n550 163.367
R1033 B.n650 B.n648 163.367
R1034 B.n654 B.n548 163.367
R1035 B.n658 B.n656 163.367
R1036 B.n662 B.n546 163.367
R1037 B.n666 B.n664 163.367
R1038 B.n670 B.n544 163.367
R1039 B.n674 B.n672 163.367
R1040 B.n678 B.n542 163.367
R1041 B.n682 B.n680 163.367
R1042 B.n686 B.n540 163.367
R1043 B.n690 B.n688 163.367
R1044 B.n695 B.n536 163.367
R1045 B.n699 B.n697 163.367
R1046 B.n703 B.n534 163.367
R1047 B.n707 B.n705 163.367
R1048 B.n711 B.n532 163.367
R1049 B.n715 B.n713 163.367
R1050 B.n719 B.n527 163.367
R1051 B.n723 B.n721 163.367
R1052 B.n727 B.n525 163.367
R1053 B.n731 B.n729 163.367
R1054 B.n735 B.n523 163.367
R1055 B.n739 B.n737 163.367
R1056 B.n743 B.n521 163.367
R1057 B.n747 B.n745 163.367
R1058 B.n751 B.n519 163.367
R1059 B.n755 B.n753 163.367
R1060 B.n759 B.n517 163.367
R1061 B.n763 B.n761 163.367
R1062 B.n767 B.n515 163.367
R1063 B.n771 B.n769 163.367
R1064 B.n775 B.n513 163.367
R1065 B.n779 B.n777 163.367
R1066 B.n783 B.n511 163.367
R1067 B.n787 B.n785 163.367
R1068 B.n791 B.n509 163.367
R1069 B.n795 B.n793 163.367
R1070 B.n799 B.n507 163.367
R1071 B.n803 B.n801 163.367
R1072 B.n807 B.n505 163.367
R1073 B.n811 B.n809 163.367
R1074 B.n815 B.n503 163.367
R1075 B.n819 B.n817 163.367
R1076 B.n823 B.n501 163.367
R1077 B.n827 B.n825 163.367
R1078 B.n831 B.n499 163.367
R1079 B.n834 B.n833 163.367
R1080 B.n836 B.n496 163.367
R1081 B.n842 B.n492 163.367
R1082 B.n846 B.n492 163.367
R1083 B.n846 B.n486 163.367
R1084 B.n854 B.n486 163.367
R1085 B.n854 B.n484 163.367
R1086 B.n858 B.n484 163.367
R1087 B.n858 B.n478 163.367
R1088 B.n866 B.n478 163.367
R1089 B.n866 B.n476 163.367
R1090 B.n870 B.n476 163.367
R1091 B.n870 B.n470 163.367
R1092 B.n878 B.n470 163.367
R1093 B.n878 B.n468 163.367
R1094 B.n882 B.n468 163.367
R1095 B.n882 B.n462 163.367
R1096 B.n890 B.n462 163.367
R1097 B.n890 B.n460 163.367
R1098 B.n894 B.n460 163.367
R1099 B.n894 B.n454 163.367
R1100 B.n902 B.n454 163.367
R1101 B.n902 B.n452 163.367
R1102 B.n906 B.n452 163.367
R1103 B.n906 B.n446 163.367
R1104 B.n914 B.n446 163.367
R1105 B.n914 B.n444 163.367
R1106 B.n918 B.n444 163.367
R1107 B.n918 B.n438 163.367
R1108 B.n927 B.n438 163.367
R1109 B.n927 B.n436 163.367
R1110 B.n931 B.n436 163.367
R1111 B.n931 B.n431 163.367
R1112 B.n939 B.n431 163.367
R1113 B.n939 B.n429 163.367
R1114 B.n943 B.n429 163.367
R1115 B.n943 B.n423 163.367
R1116 B.n952 B.n423 163.367
R1117 B.n952 B.n421 163.367
R1118 B.n956 B.n421 163.367
R1119 B.n956 B.n3 163.367
R1120 B.n1100 B.n3 163.367
R1121 B.n1096 B.n2 163.367
R1122 B.n1096 B.n1095 163.367
R1123 B.n1095 B.n9 163.367
R1124 B.n1091 B.n9 163.367
R1125 B.n1091 B.n11 163.367
R1126 B.n1087 B.n11 163.367
R1127 B.n1087 B.n17 163.367
R1128 B.n1083 B.n17 163.367
R1129 B.n1083 B.n19 163.367
R1130 B.n1079 B.n19 163.367
R1131 B.n1079 B.n23 163.367
R1132 B.n1075 B.n23 163.367
R1133 B.n1075 B.n25 163.367
R1134 B.n1071 B.n25 163.367
R1135 B.n1071 B.n31 163.367
R1136 B.n1067 B.n31 163.367
R1137 B.n1067 B.n33 163.367
R1138 B.n1063 B.n33 163.367
R1139 B.n1063 B.n38 163.367
R1140 B.n1059 B.n38 163.367
R1141 B.n1059 B.n40 163.367
R1142 B.n1055 B.n40 163.367
R1143 B.n1055 B.n45 163.367
R1144 B.n1051 B.n45 163.367
R1145 B.n1051 B.n47 163.367
R1146 B.n1047 B.n47 163.367
R1147 B.n1047 B.n52 163.367
R1148 B.n1043 B.n52 163.367
R1149 B.n1043 B.n54 163.367
R1150 B.n1039 B.n54 163.367
R1151 B.n1039 B.n59 163.367
R1152 B.n1035 B.n59 163.367
R1153 B.n1035 B.n61 163.367
R1154 B.n1031 B.n61 163.367
R1155 B.n1031 B.n66 163.367
R1156 B.n1027 B.n66 163.367
R1157 B.n1027 B.n68 163.367
R1158 B.n1023 B.n68 163.367
R1159 B.n1023 B.n73 163.367
R1160 B.n1019 B.n73 163.367
R1161 B.n145 B.t10 114.694
R1162 B.n528 B.t15 114.694
R1163 B.n147 B.t20 114.668
R1164 B.n537 B.t18 114.668
R1165 B.n77 B.n75 71.676
R1166 B.n151 B.n78 71.676
R1167 B.n155 B.n79 71.676
R1168 B.n159 B.n80 71.676
R1169 B.n163 B.n81 71.676
R1170 B.n167 B.n82 71.676
R1171 B.n171 B.n83 71.676
R1172 B.n175 B.n84 71.676
R1173 B.n179 B.n85 71.676
R1174 B.n183 B.n86 71.676
R1175 B.n187 B.n87 71.676
R1176 B.n191 B.n88 71.676
R1177 B.n195 B.n89 71.676
R1178 B.n199 B.n90 71.676
R1179 B.n203 B.n91 71.676
R1180 B.n207 B.n92 71.676
R1181 B.n211 B.n93 71.676
R1182 B.n215 B.n94 71.676
R1183 B.n219 B.n95 71.676
R1184 B.n223 B.n96 71.676
R1185 B.n227 B.n97 71.676
R1186 B.n231 B.n98 71.676
R1187 B.n235 B.n99 71.676
R1188 B.n239 B.n100 71.676
R1189 B.n243 B.n101 71.676
R1190 B.n247 B.n102 71.676
R1191 B.n251 B.n103 71.676
R1192 B.n255 B.n104 71.676
R1193 B.n259 B.n105 71.676
R1194 B.n263 B.n106 71.676
R1195 B.n267 B.n107 71.676
R1196 B.n271 B.n108 71.676
R1197 B.n276 B.n109 71.676
R1198 B.n280 B.n110 71.676
R1199 B.n284 B.n111 71.676
R1200 B.n288 B.n112 71.676
R1201 B.n292 B.n113 71.676
R1202 B.n297 B.n114 71.676
R1203 B.n301 B.n115 71.676
R1204 B.n305 B.n116 71.676
R1205 B.n309 B.n117 71.676
R1206 B.n313 B.n118 71.676
R1207 B.n317 B.n119 71.676
R1208 B.n321 B.n120 71.676
R1209 B.n325 B.n121 71.676
R1210 B.n329 B.n122 71.676
R1211 B.n333 B.n123 71.676
R1212 B.n337 B.n124 71.676
R1213 B.n341 B.n125 71.676
R1214 B.n345 B.n126 71.676
R1215 B.n349 B.n127 71.676
R1216 B.n353 B.n128 71.676
R1217 B.n357 B.n129 71.676
R1218 B.n361 B.n130 71.676
R1219 B.n365 B.n131 71.676
R1220 B.n369 B.n132 71.676
R1221 B.n373 B.n133 71.676
R1222 B.n377 B.n134 71.676
R1223 B.n381 B.n135 71.676
R1224 B.n385 B.n136 71.676
R1225 B.n389 B.n137 71.676
R1226 B.n393 B.n138 71.676
R1227 B.n397 B.n139 71.676
R1228 B.n401 B.n140 71.676
R1229 B.n405 B.n141 71.676
R1230 B.n409 B.n142 71.676
R1231 B.n413 B.n143 71.676
R1232 B.n1016 B.n144 71.676
R1233 B.n1016 B.n1015 71.676
R1234 B.n415 B.n143 71.676
R1235 B.n412 B.n142 71.676
R1236 B.n408 B.n141 71.676
R1237 B.n404 B.n140 71.676
R1238 B.n400 B.n139 71.676
R1239 B.n396 B.n138 71.676
R1240 B.n392 B.n137 71.676
R1241 B.n388 B.n136 71.676
R1242 B.n384 B.n135 71.676
R1243 B.n380 B.n134 71.676
R1244 B.n376 B.n133 71.676
R1245 B.n372 B.n132 71.676
R1246 B.n368 B.n131 71.676
R1247 B.n364 B.n130 71.676
R1248 B.n360 B.n129 71.676
R1249 B.n356 B.n128 71.676
R1250 B.n352 B.n127 71.676
R1251 B.n348 B.n126 71.676
R1252 B.n344 B.n125 71.676
R1253 B.n340 B.n124 71.676
R1254 B.n336 B.n123 71.676
R1255 B.n332 B.n122 71.676
R1256 B.n328 B.n121 71.676
R1257 B.n324 B.n120 71.676
R1258 B.n320 B.n119 71.676
R1259 B.n316 B.n118 71.676
R1260 B.n312 B.n117 71.676
R1261 B.n308 B.n116 71.676
R1262 B.n304 B.n115 71.676
R1263 B.n300 B.n114 71.676
R1264 B.n296 B.n113 71.676
R1265 B.n291 B.n112 71.676
R1266 B.n287 B.n111 71.676
R1267 B.n283 B.n110 71.676
R1268 B.n279 B.n109 71.676
R1269 B.n275 B.n108 71.676
R1270 B.n270 B.n107 71.676
R1271 B.n266 B.n106 71.676
R1272 B.n262 B.n105 71.676
R1273 B.n258 B.n104 71.676
R1274 B.n254 B.n103 71.676
R1275 B.n250 B.n102 71.676
R1276 B.n246 B.n101 71.676
R1277 B.n242 B.n100 71.676
R1278 B.n238 B.n99 71.676
R1279 B.n234 B.n98 71.676
R1280 B.n230 B.n97 71.676
R1281 B.n226 B.n96 71.676
R1282 B.n222 B.n95 71.676
R1283 B.n218 B.n94 71.676
R1284 B.n214 B.n93 71.676
R1285 B.n210 B.n92 71.676
R1286 B.n206 B.n91 71.676
R1287 B.n202 B.n90 71.676
R1288 B.n198 B.n89 71.676
R1289 B.n194 B.n88 71.676
R1290 B.n190 B.n87 71.676
R1291 B.n186 B.n86 71.676
R1292 B.n182 B.n85 71.676
R1293 B.n178 B.n84 71.676
R1294 B.n174 B.n83 71.676
R1295 B.n170 B.n82 71.676
R1296 B.n166 B.n81 71.676
R1297 B.n162 B.n80 71.676
R1298 B.n158 B.n79 71.676
R1299 B.n154 B.n78 71.676
R1300 B.n150 B.n77 71.676
R1301 B.n569 B.n494 71.676
R1302 B.n575 B.n574 71.676
R1303 B.n578 B.n577 71.676
R1304 B.n583 B.n582 71.676
R1305 B.n586 B.n585 71.676
R1306 B.n591 B.n590 71.676
R1307 B.n594 B.n593 71.676
R1308 B.n599 B.n598 71.676
R1309 B.n602 B.n601 71.676
R1310 B.n607 B.n606 71.676
R1311 B.n610 B.n609 71.676
R1312 B.n615 B.n614 71.676
R1313 B.n618 B.n617 71.676
R1314 B.n623 B.n622 71.676
R1315 B.n626 B.n625 71.676
R1316 B.n631 B.n630 71.676
R1317 B.n634 B.n633 71.676
R1318 B.n639 B.n638 71.676
R1319 B.n642 B.n641 71.676
R1320 B.n647 B.n646 71.676
R1321 B.n650 B.n649 71.676
R1322 B.n655 B.n654 71.676
R1323 B.n658 B.n657 71.676
R1324 B.n663 B.n662 71.676
R1325 B.n666 B.n665 71.676
R1326 B.n671 B.n670 71.676
R1327 B.n674 B.n673 71.676
R1328 B.n679 B.n678 71.676
R1329 B.n682 B.n681 71.676
R1330 B.n687 B.n686 71.676
R1331 B.n690 B.n689 71.676
R1332 B.n696 B.n695 71.676
R1333 B.n699 B.n698 71.676
R1334 B.n704 B.n703 71.676
R1335 B.n707 B.n706 71.676
R1336 B.n712 B.n711 71.676
R1337 B.n715 B.n714 71.676
R1338 B.n720 B.n719 71.676
R1339 B.n723 B.n722 71.676
R1340 B.n728 B.n727 71.676
R1341 B.n731 B.n730 71.676
R1342 B.n736 B.n735 71.676
R1343 B.n739 B.n738 71.676
R1344 B.n744 B.n743 71.676
R1345 B.n747 B.n746 71.676
R1346 B.n752 B.n751 71.676
R1347 B.n755 B.n754 71.676
R1348 B.n760 B.n759 71.676
R1349 B.n763 B.n762 71.676
R1350 B.n768 B.n767 71.676
R1351 B.n771 B.n770 71.676
R1352 B.n776 B.n775 71.676
R1353 B.n779 B.n778 71.676
R1354 B.n784 B.n783 71.676
R1355 B.n787 B.n786 71.676
R1356 B.n792 B.n791 71.676
R1357 B.n795 B.n794 71.676
R1358 B.n800 B.n799 71.676
R1359 B.n803 B.n802 71.676
R1360 B.n808 B.n807 71.676
R1361 B.n811 B.n810 71.676
R1362 B.n816 B.n815 71.676
R1363 B.n819 B.n818 71.676
R1364 B.n824 B.n823 71.676
R1365 B.n827 B.n826 71.676
R1366 B.n832 B.n831 71.676
R1367 B.n835 B.n834 71.676
R1368 B.n570 B.n569 71.676
R1369 B.n576 B.n575 71.676
R1370 B.n577 B.n566 71.676
R1371 B.n584 B.n583 71.676
R1372 B.n585 B.n564 71.676
R1373 B.n592 B.n591 71.676
R1374 B.n593 B.n562 71.676
R1375 B.n600 B.n599 71.676
R1376 B.n601 B.n560 71.676
R1377 B.n608 B.n607 71.676
R1378 B.n609 B.n558 71.676
R1379 B.n616 B.n615 71.676
R1380 B.n617 B.n556 71.676
R1381 B.n624 B.n623 71.676
R1382 B.n625 B.n554 71.676
R1383 B.n632 B.n631 71.676
R1384 B.n633 B.n552 71.676
R1385 B.n640 B.n639 71.676
R1386 B.n641 B.n550 71.676
R1387 B.n648 B.n647 71.676
R1388 B.n649 B.n548 71.676
R1389 B.n656 B.n655 71.676
R1390 B.n657 B.n546 71.676
R1391 B.n664 B.n663 71.676
R1392 B.n665 B.n544 71.676
R1393 B.n672 B.n671 71.676
R1394 B.n673 B.n542 71.676
R1395 B.n680 B.n679 71.676
R1396 B.n681 B.n540 71.676
R1397 B.n688 B.n687 71.676
R1398 B.n689 B.n536 71.676
R1399 B.n697 B.n696 71.676
R1400 B.n698 B.n534 71.676
R1401 B.n705 B.n704 71.676
R1402 B.n706 B.n532 71.676
R1403 B.n713 B.n712 71.676
R1404 B.n714 B.n527 71.676
R1405 B.n721 B.n720 71.676
R1406 B.n722 B.n525 71.676
R1407 B.n729 B.n728 71.676
R1408 B.n730 B.n523 71.676
R1409 B.n737 B.n736 71.676
R1410 B.n738 B.n521 71.676
R1411 B.n745 B.n744 71.676
R1412 B.n746 B.n519 71.676
R1413 B.n753 B.n752 71.676
R1414 B.n754 B.n517 71.676
R1415 B.n761 B.n760 71.676
R1416 B.n762 B.n515 71.676
R1417 B.n769 B.n768 71.676
R1418 B.n770 B.n513 71.676
R1419 B.n777 B.n776 71.676
R1420 B.n778 B.n511 71.676
R1421 B.n785 B.n784 71.676
R1422 B.n786 B.n509 71.676
R1423 B.n793 B.n792 71.676
R1424 B.n794 B.n507 71.676
R1425 B.n801 B.n800 71.676
R1426 B.n802 B.n505 71.676
R1427 B.n809 B.n808 71.676
R1428 B.n810 B.n503 71.676
R1429 B.n817 B.n816 71.676
R1430 B.n818 B.n501 71.676
R1431 B.n825 B.n824 71.676
R1432 B.n826 B.n499 71.676
R1433 B.n833 B.n832 71.676
R1434 B.n836 B.n835 71.676
R1435 B.n1101 B.n1100 71.676
R1436 B.n1101 B.n2 71.676
R1437 B.n146 B.t11 71.6385
R1438 B.n529 B.t14 71.6385
R1439 B.n148 B.t21 71.6128
R1440 B.n538 B.t17 71.6128
R1441 B.n841 B.n495 63.1906
R1442 B.n1018 B.n1017 63.1906
R1443 B.n273 B.n148 59.5399
R1444 B.n294 B.n146 59.5399
R1445 B.n530 B.n529 59.5399
R1446 B.n693 B.n538 59.5399
R1447 B.n148 B.n147 43.055
R1448 B.n146 B.n145 43.055
R1449 B.n529 B.n528 43.055
R1450 B.n538 B.n537 43.055
R1451 B.n843 B.n493 32.9371
R1452 B.n839 B.n838 32.9371
R1453 B.n1014 B.n1013 32.9371
R1454 B.n1020 B.n74 32.9371
R1455 B.n841 B.n491 30.4751
R1456 B.n847 B.n491 30.4751
R1457 B.n847 B.n487 30.4751
R1458 B.n853 B.n487 30.4751
R1459 B.n853 B.n483 30.4751
R1460 B.n859 B.n483 30.4751
R1461 B.n865 B.n479 30.4751
R1462 B.n865 B.n475 30.4751
R1463 B.n871 B.n475 30.4751
R1464 B.n871 B.n471 30.4751
R1465 B.n877 B.n471 30.4751
R1466 B.n877 B.n467 30.4751
R1467 B.n883 B.n467 30.4751
R1468 B.n883 B.n463 30.4751
R1469 B.n889 B.n463 30.4751
R1470 B.n895 B.n459 30.4751
R1471 B.n895 B.n455 30.4751
R1472 B.n901 B.n455 30.4751
R1473 B.n901 B.n451 30.4751
R1474 B.n907 B.n451 30.4751
R1475 B.n913 B.n447 30.4751
R1476 B.n913 B.n443 30.4751
R1477 B.n919 B.n443 30.4751
R1478 B.n919 B.n439 30.4751
R1479 B.n926 B.n439 30.4751
R1480 B.n926 B.n925 30.4751
R1481 B.n932 B.n432 30.4751
R1482 B.n938 B.n432 30.4751
R1483 B.n938 B.n427 30.4751
R1484 B.n944 B.n427 30.4751
R1485 B.n944 B.n428 30.4751
R1486 B.n951 B.n420 30.4751
R1487 B.n957 B.n420 30.4751
R1488 B.n957 B.n4 30.4751
R1489 B.n1099 B.n4 30.4751
R1490 B.n1099 B.n1098 30.4751
R1491 B.n1098 B.n1097 30.4751
R1492 B.n1097 B.n8 30.4751
R1493 B.n12 B.n8 30.4751
R1494 B.n1090 B.n12 30.4751
R1495 B.n1089 B.n1088 30.4751
R1496 B.n1088 B.n16 30.4751
R1497 B.n1082 B.n16 30.4751
R1498 B.n1082 B.n1081 30.4751
R1499 B.n1081 B.n1080 30.4751
R1500 B.n1074 B.n26 30.4751
R1501 B.n1074 B.n1073 30.4751
R1502 B.n1073 B.n1072 30.4751
R1503 B.n1072 B.n30 30.4751
R1504 B.n1066 B.n30 30.4751
R1505 B.n1066 B.n1065 30.4751
R1506 B.n1064 B.n37 30.4751
R1507 B.n1058 B.n37 30.4751
R1508 B.n1058 B.n1057 30.4751
R1509 B.n1057 B.n1056 30.4751
R1510 B.n1056 B.n44 30.4751
R1511 B.n1050 B.n1049 30.4751
R1512 B.n1049 B.n1048 30.4751
R1513 B.n1048 B.n51 30.4751
R1514 B.n1042 B.n51 30.4751
R1515 B.n1042 B.n1041 30.4751
R1516 B.n1041 B.n1040 30.4751
R1517 B.n1040 B.n58 30.4751
R1518 B.n1034 B.n58 30.4751
R1519 B.n1034 B.n1033 30.4751
R1520 B.n1032 B.n65 30.4751
R1521 B.n1026 B.n65 30.4751
R1522 B.n1026 B.n1025 30.4751
R1523 B.n1025 B.n1024 30.4751
R1524 B.n1024 B.n72 30.4751
R1525 B.n1018 B.n72 30.4751
R1526 B.t0 B.n459 29.1307
R1527 B.t6 B.n44 29.1307
R1528 B.n932 B.t4 27.338
R1529 B.n1080 B.t2 27.338
R1530 B.t13 B.n479 21.0639
R1531 B.n1033 B.t9 21.0639
R1532 B.n428 B.t7 19.2712
R1533 B.t5 B.n1089 19.2712
R1534 B B.n1102 18.0485
R1535 B.n907 B.t1 17.4786
R1536 B.t3 B.n1064 17.4786
R1537 B.t1 B.n447 12.997
R1538 B.n1065 B.t3 12.997
R1539 B.n951 B.t7 11.2044
R1540 B.n1090 B.t5 11.2044
R1541 B.n844 B.n843 10.6151
R1542 B.n845 B.n844 10.6151
R1543 B.n845 B.n485 10.6151
R1544 B.n855 B.n485 10.6151
R1545 B.n856 B.n855 10.6151
R1546 B.n857 B.n856 10.6151
R1547 B.n857 B.n477 10.6151
R1548 B.n867 B.n477 10.6151
R1549 B.n868 B.n867 10.6151
R1550 B.n869 B.n868 10.6151
R1551 B.n869 B.n469 10.6151
R1552 B.n879 B.n469 10.6151
R1553 B.n880 B.n879 10.6151
R1554 B.n881 B.n880 10.6151
R1555 B.n881 B.n461 10.6151
R1556 B.n891 B.n461 10.6151
R1557 B.n892 B.n891 10.6151
R1558 B.n893 B.n892 10.6151
R1559 B.n893 B.n453 10.6151
R1560 B.n903 B.n453 10.6151
R1561 B.n904 B.n903 10.6151
R1562 B.n905 B.n904 10.6151
R1563 B.n905 B.n445 10.6151
R1564 B.n915 B.n445 10.6151
R1565 B.n916 B.n915 10.6151
R1566 B.n917 B.n916 10.6151
R1567 B.n917 B.n437 10.6151
R1568 B.n928 B.n437 10.6151
R1569 B.n929 B.n928 10.6151
R1570 B.n930 B.n929 10.6151
R1571 B.n930 B.n430 10.6151
R1572 B.n940 B.n430 10.6151
R1573 B.n941 B.n940 10.6151
R1574 B.n942 B.n941 10.6151
R1575 B.n942 B.n422 10.6151
R1576 B.n953 B.n422 10.6151
R1577 B.n954 B.n953 10.6151
R1578 B.n955 B.n954 10.6151
R1579 B.n955 B.n0 10.6151
R1580 B.n571 B.n493 10.6151
R1581 B.n572 B.n571 10.6151
R1582 B.n573 B.n572 10.6151
R1583 B.n573 B.n567 10.6151
R1584 B.n579 B.n567 10.6151
R1585 B.n580 B.n579 10.6151
R1586 B.n581 B.n580 10.6151
R1587 B.n581 B.n565 10.6151
R1588 B.n587 B.n565 10.6151
R1589 B.n588 B.n587 10.6151
R1590 B.n589 B.n588 10.6151
R1591 B.n589 B.n563 10.6151
R1592 B.n595 B.n563 10.6151
R1593 B.n596 B.n595 10.6151
R1594 B.n597 B.n596 10.6151
R1595 B.n597 B.n561 10.6151
R1596 B.n603 B.n561 10.6151
R1597 B.n604 B.n603 10.6151
R1598 B.n605 B.n604 10.6151
R1599 B.n605 B.n559 10.6151
R1600 B.n611 B.n559 10.6151
R1601 B.n612 B.n611 10.6151
R1602 B.n613 B.n612 10.6151
R1603 B.n613 B.n557 10.6151
R1604 B.n619 B.n557 10.6151
R1605 B.n620 B.n619 10.6151
R1606 B.n621 B.n620 10.6151
R1607 B.n621 B.n555 10.6151
R1608 B.n627 B.n555 10.6151
R1609 B.n628 B.n627 10.6151
R1610 B.n629 B.n628 10.6151
R1611 B.n629 B.n553 10.6151
R1612 B.n635 B.n553 10.6151
R1613 B.n636 B.n635 10.6151
R1614 B.n637 B.n636 10.6151
R1615 B.n637 B.n551 10.6151
R1616 B.n643 B.n551 10.6151
R1617 B.n644 B.n643 10.6151
R1618 B.n645 B.n644 10.6151
R1619 B.n645 B.n549 10.6151
R1620 B.n651 B.n549 10.6151
R1621 B.n652 B.n651 10.6151
R1622 B.n653 B.n652 10.6151
R1623 B.n653 B.n547 10.6151
R1624 B.n659 B.n547 10.6151
R1625 B.n660 B.n659 10.6151
R1626 B.n661 B.n660 10.6151
R1627 B.n661 B.n545 10.6151
R1628 B.n667 B.n545 10.6151
R1629 B.n668 B.n667 10.6151
R1630 B.n669 B.n668 10.6151
R1631 B.n669 B.n543 10.6151
R1632 B.n675 B.n543 10.6151
R1633 B.n676 B.n675 10.6151
R1634 B.n677 B.n676 10.6151
R1635 B.n677 B.n541 10.6151
R1636 B.n683 B.n541 10.6151
R1637 B.n684 B.n683 10.6151
R1638 B.n685 B.n684 10.6151
R1639 B.n685 B.n539 10.6151
R1640 B.n691 B.n539 10.6151
R1641 B.n692 B.n691 10.6151
R1642 B.n694 B.n535 10.6151
R1643 B.n700 B.n535 10.6151
R1644 B.n701 B.n700 10.6151
R1645 B.n702 B.n701 10.6151
R1646 B.n702 B.n533 10.6151
R1647 B.n708 B.n533 10.6151
R1648 B.n709 B.n708 10.6151
R1649 B.n710 B.n709 10.6151
R1650 B.n710 B.n531 10.6151
R1651 B.n717 B.n716 10.6151
R1652 B.n718 B.n717 10.6151
R1653 B.n718 B.n526 10.6151
R1654 B.n724 B.n526 10.6151
R1655 B.n725 B.n724 10.6151
R1656 B.n726 B.n725 10.6151
R1657 B.n726 B.n524 10.6151
R1658 B.n732 B.n524 10.6151
R1659 B.n733 B.n732 10.6151
R1660 B.n734 B.n733 10.6151
R1661 B.n734 B.n522 10.6151
R1662 B.n740 B.n522 10.6151
R1663 B.n741 B.n740 10.6151
R1664 B.n742 B.n741 10.6151
R1665 B.n742 B.n520 10.6151
R1666 B.n748 B.n520 10.6151
R1667 B.n749 B.n748 10.6151
R1668 B.n750 B.n749 10.6151
R1669 B.n750 B.n518 10.6151
R1670 B.n756 B.n518 10.6151
R1671 B.n757 B.n756 10.6151
R1672 B.n758 B.n757 10.6151
R1673 B.n758 B.n516 10.6151
R1674 B.n764 B.n516 10.6151
R1675 B.n765 B.n764 10.6151
R1676 B.n766 B.n765 10.6151
R1677 B.n766 B.n514 10.6151
R1678 B.n772 B.n514 10.6151
R1679 B.n773 B.n772 10.6151
R1680 B.n774 B.n773 10.6151
R1681 B.n774 B.n512 10.6151
R1682 B.n780 B.n512 10.6151
R1683 B.n781 B.n780 10.6151
R1684 B.n782 B.n781 10.6151
R1685 B.n782 B.n510 10.6151
R1686 B.n788 B.n510 10.6151
R1687 B.n789 B.n788 10.6151
R1688 B.n790 B.n789 10.6151
R1689 B.n790 B.n508 10.6151
R1690 B.n796 B.n508 10.6151
R1691 B.n797 B.n796 10.6151
R1692 B.n798 B.n797 10.6151
R1693 B.n798 B.n506 10.6151
R1694 B.n804 B.n506 10.6151
R1695 B.n805 B.n804 10.6151
R1696 B.n806 B.n805 10.6151
R1697 B.n806 B.n504 10.6151
R1698 B.n812 B.n504 10.6151
R1699 B.n813 B.n812 10.6151
R1700 B.n814 B.n813 10.6151
R1701 B.n814 B.n502 10.6151
R1702 B.n820 B.n502 10.6151
R1703 B.n821 B.n820 10.6151
R1704 B.n822 B.n821 10.6151
R1705 B.n822 B.n500 10.6151
R1706 B.n828 B.n500 10.6151
R1707 B.n829 B.n828 10.6151
R1708 B.n830 B.n829 10.6151
R1709 B.n830 B.n498 10.6151
R1710 B.n498 B.n497 10.6151
R1711 B.n837 B.n497 10.6151
R1712 B.n838 B.n837 10.6151
R1713 B.n839 B.n489 10.6151
R1714 B.n849 B.n489 10.6151
R1715 B.n850 B.n849 10.6151
R1716 B.n851 B.n850 10.6151
R1717 B.n851 B.n481 10.6151
R1718 B.n861 B.n481 10.6151
R1719 B.n862 B.n861 10.6151
R1720 B.n863 B.n862 10.6151
R1721 B.n863 B.n473 10.6151
R1722 B.n873 B.n473 10.6151
R1723 B.n874 B.n873 10.6151
R1724 B.n875 B.n874 10.6151
R1725 B.n875 B.n465 10.6151
R1726 B.n885 B.n465 10.6151
R1727 B.n886 B.n885 10.6151
R1728 B.n887 B.n886 10.6151
R1729 B.n887 B.n457 10.6151
R1730 B.n897 B.n457 10.6151
R1731 B.n898 B.n897 10.6151
R1732 B.n899 B.n898 10.6151
R1733 B.n899 B.n449 10.6151
R1734 B.n909 B.n449 10.6151
R1735 B.n910 B.n909 10.6151
R1736 B.n911 B.n910 10.6151
R1737 B.n911 B.n441 10.6151
R1738 B.n921 B.n441 10.6151
R1739 B.n922 B.n921 10.6151
R1740 B.n923 B.n922 10.6151
R1741 B.n923 B.n434 10.6151
R1742 B.n934 B.n434 10.6151
R1743 B.n935 B.n934 10.6151
R1744 B.n936 B.n935 10.6151
R1745 B.n936 B.n425 10.6151
R1746 B.n946 B.n425 10.6151
R1747 B.n947 B.n946 10.6151
R1748 B.n949 B.n947 10.6151
R1749 B.n949 B.n948 10.6151
R1750 B.n948 B.n418 10.6151
R1751 B.n960 B.n418 10.6151
R1752 B.n961 B.n960 10.6151
R1753 B.n962 B.n961 10.6151
R1754 B.n963 B.n962 10.6151
R1755 B.n964 B.n963 10.6151
R1756 B.n967 B.n964 10.6151
R1757 B.n968 B.n967 10.6151
R1758 B.n969 B.n968 10.6151
R1759 B.n970 B.n969 10.6151
R1760 B.n972 B.n970 10.6151
R1761 B.n973 B.n972 10.6151
R1762 B.n974 B.n973 10.6151
R1763 B.n975 B.n974 10.6151
R1764 B.n977 B.n975 10.6151
R1765 B.n978 B.n977 10.6151
R1766 B.n979 B.n978 10.6151
R1767 B.n980 B.n979 10.6151
R1768 B.n982 B.n980 10.6151
R1769 B.n983 B.n982 10.6151
R1770 B.n984 B.n983 10.6151
R1771 B.n985 B.n984 10.6151
R1772 B.n987 B.n985 10.6151
R1773 B.n988 B.n987 10.6151
R1774 B.n989 B.n988 10.6151
R1775 B.n990 B.n989 10.6151
R1776 B.n992 B.n990 10.6151
R1777 B.n993 B.n992 10.6151
R1778 B.n994 B.n993 10.6151
R1779 B.n995 B.n994 10.6151
R1780 B.n997 B.n995 10.6151
R1781 B.n998 B.n997 10.6151
R1782 B.n999 B.n998 10.6151
R1783 B.n1000 B.n999 10.6151
R1784 B.n1002 B.n1000 10.6151
R1785 B.n1003 B.n1002 10.6151
R1786 B.n1004 B.n1003 10.6151
R1787 B.n1005 B.n1004 10.6151
R1788 B.n1007 B.n1005 10.6151
R1789 B.n1008 B.n1007 10.6151
R1790 B.n1009 B.n1008 10.6151
R1791 B.n1010 B.n1009 10.6151
R1792 B.n1012 B.n1010 10.6151
R1793 B.n1013 B.n1012 10.6151
R1794 B.n1094 B.n1 10.6151
R1795 B.n1094 B.n1093 10.6151
R1796 B.n1093 B.n1092 10.6151
R1797 B.n1092 B.n10 10.6151
R1798 B.n1086 B.n10 10.6151
R1799 B.n1086 B.n1085 10.6151
R1800 B.n1085 B.n1084 10.6151
R1801 B.n1084 B.n18 10.6151
R1802 B.n1078 B.n18 10.6151
R1803 B.n1078 B.n1077 10.6151
R1804 B.n1077 B.n1076 10.6151
R1805 B.n1076 B.n24 10.6151
R1806 B.n1070 B.n24 10.6151
R1807 B.n1070 B.n1069 10.6151
R1808 B.n1069 B.n1068 10.6151
R1809 B.n1068 B.n32 10.6151
R1810 B.n1062 B.n32 10.6151
R1811 B.n1062 B.n1061 10.6151
R1812 B.n1061 B.n1060 10.6151
R1813 B.n1060 B.n39 10.6151
R1814 B.n1054 B.n39 10.6151
R1815 B.n1054 B.n1053 10.6151
R1816 B.n1053 B.n1052 10.6151
R1817 B.n1052 B.n46 10.6151
R1818 B.n1046 B.n46 10.6151
R1819 B.n1046 B.n1045 10.6151
R1820 B.n1045 B.n1044 10.6151
R1821 B.n1044 B.n53 10.6151
R1822 B.n1038 B.n53 10.6151
R1823 B.n1038 B.n1037 10.6151
R1824 B.n1037 B.n1036 10.6151
R1825 B.n1036 B.n60 10.6151
R1826 B.n1030 B.n60 10.6151
R1827 B.n1030 B.n1029 10.6151
R1828 B.n1029 B.n1028 10.6151
R1829 B.n1028 B.n67 10.6151
R1830 B.n1022 B.n67 10.6151
R1831 B.n1022 B.n1021 10.6151
R1832 B.n1021 B.n1020 10.6151
R1833 B.n149 B.n74 10.6151
R1834 B.n152 B.n149 10.6151
R1835 B.n153 B.n152 10.6151
R1836 B.n156 B.n153 10.6151
R1837 B.n157 B.n156 10.6151
R1838 B.n160 B.n157 10.6151
R1839 B.n161 B.n160 10.6151
R1840 B.n164 B.n161 10.6151
R1841 B.n165 B.n164 10.6151
R1842 B.n168 B.n165 10.6151
R1843 B.n169 B.n168 10.6151
R1844 B.n172 B.n169 10.6151
R1845 B.n173 B.n172 10.6151
R1846 B.n176 B.n173 10.6151
R1847 B.n177 B.n176 10.6151
R1848 B.n180 B.n177 10.6151
R1849 B.n181 B.n180 10.6151
R1850 B.n184 B.n181 10.6151
R1851 B.n185 B.n184 10.6151
R1852 B.n188 B.n185 10.6151
R1853 B.n189 B.n188 10.6151
R1854 B.n192 B.n189 10.6151
R1855 B.n193 B.n192 10.6151
R1856 B.n196 B.n193 10.6151
R1857 B.n197 B.n196 10.6151
R1858 B.n200 B.n197 10.6151
R1859 B.n201 B.n200 10.6151
R1860 B.n204 B.n201 10.6151
R1861 B.n205 B.n204 10.6151
R1862 B.n208 B.n205 10.6151
R1863 B.n209 B.n208 10.6151
R1864 B.n212 B.n209 10.6151
R1865 B.n213 B.n212 10.6151
R1866 B.n216 B.n213 10.6151
R1867 B.n217 B.n216 10.6151
R1868 B.n220 B.n217 10.6151
R1869 B.n221 B.n220 10.6151
R1870 B.n224 B.n221 10.6151
R1871 B.n225 B.n224 10.6151
R1872 B.n228 B.n225 10.6151
R1873 B.n229 B.n228 10.6151
R1874 B.n232 B.n229 10.6151
R1875 B.n233 B.n232 10.6151
R1876 B.n236 B.n233 10.6151
R1877 B.n237 B.n236 10.6151
R1878 B.n240 B.n237 10.6151
R1879 B.n241 B.n240 10.6151
R1880 B.n244 B.n241 10.6151
R1881 B.n245 B.n244 10.6151
R1882 B.n248 B.n245 10.6151
R1883 B.n249 B.n248 10.6151
R1884 B.n252 B.n249 10.6151
R1885 B.n253 B.n252 10.6151
R1886 B.n256 B.n253 10.6151
R1887 B.n257 B.n256 10.6151
R1888 B.n260 B.n257 10.6151
R1889 B.n261 B.n260 10.6151
R1890 B.n264 B.n261 10.6151
R1891 B.n265 B.n264 10.6151
R1892 B.n268 B.n265 10.6151
R1893 B.n269 B.n268 10.6151
R1894 B.n272 B.n269 10.6151
R1895 B.n277 B.n274 10.6151
R1896 B.n278 B.n277 10.6151
R1897 B.n281 B.n278 10.6151
R1898 B.n282 B.n281 10.6151
R1899 B.n285 B.n282 10.6151
R1900 B.n286 B.n285 10.6151
R1901 B.n289 B.n286 10.6151
R1902 B.n290 B.n289 10.6151
R1903 B.n293 B.n290 10.6151
R1904 B.n298 B.n295 10.6151
R1905 B.n299 B.n298 10.6151
R1906 B.n302 B.n299 10.6151
R1907 B.n303 B.n302 10.6151
R1908 B.n306 B.n303 10.6151
R1909 B.n307 B.n306 10.6151
R1910 B.n310 B.n307 10.6151
R1911 B.n311 B.n310 10.6151
R1912 B.n314 B.n311 10.6151
R1913 B.n315 B.n314 10.6151
R1914 B.n318 B.n315 10.6151
R1915 B.n319 B.n318 10.6151
R1916 B.n322 B.n319 10.6151
R1917 B.n323 B.n322 10.6151
R1918 B.n326 B.n323 10.6151
R1919 B.n327 B.n326 10.6151
R1920 B.n330 B.n327 10.6151
R1921 B.n331 B.n330 10.6151
R1922 B.n334 B.n331 10.6151
R1923 B.n335 B.n334 10.6151
R1924 B.n338 B.n335 10.6151
R1925 B.n339 B.n338 10.6151
R1926 B.n342 B.n339 10.6151
R1927 B.n343 B.n342 10.6151
R1928 B.n346 B.n343 10.6151
R1929 B.n347 B.n346 10.6151
R1930 B.n350 B.n347 10.6151
R1931 B.n351 B.n350 10.6151
R1932 B.n354 B.n351 10.6151
R1933 B.n355 B.n354 10.6151
R1934 B.n358 B.n355 10.6151
R1935 B.n359 B.n358 10.6151
R1936 B.n362 B.n359 10.6151
R1937 B.n363 B.n362 10.6151
R1938 B.n366 B.n363 10.6151
R1939 B.n367 B.n366 10.6151
R1940 B.n370 B.n367 10.6151
R1941 B.n371 B.n370 10.6151
R1942 B.n374 B.n371 10.6151
R1943 B.n375 B.n374 10.6151
R1944 B.n378 B.n375 10.6151
R1945 B.n379 B.n378 10.6151
R1946 B.n382 B.n379 10.6151
R1947 B.n383 B.n382 10.6151
R1948 B.n386 B.n383 10.6151
R1949 B.n387 B.n386 10.6151
R1950 B.n390 B.n387 10.6151
R1951 B.n391 B.n390 10.6151
R1952 B.n394 B.n391 10.6151
R1953 B.n395 B.n394 10.6151
R1954 B.n398 B.n395 10.6151
R1955 B.n399 B.n398 10.6151
R1956 B.n402 B.n399 10.6151
R1957 B.n403 B.n402 10.6151
R1958 B.n406 B.n403 10.6151
R1959 B.n407 B.n406 10.6151
R1960 B.n410 B.n407 10.6151
R1961 B.n411 B.n410 10.6151
R1962 B.n414 B.n411 10.6151
R1963 B.n416 B.n414 10.6151
R1964 B.n417 B.n416 10.6151
R1965 B.n1014 B.n417 10.6151
R1966 B.n859 B.t13 9.41179
R1967 B.t9 B.n1032 9.41179
R1968 B.n693 B.n692 9.36635
R1969 B.n716 B.n530 9.36635
R1970 B.n273 B.n272 9.36635
R1971 B.n295 B.n294 9.36635
R1972 B.n1102 B.n0 8.11757
R1973 B.n1102 B.n1 8.11757
R1974 B.n925 B.t4 3.1376
R1975 B.n26 B.t2 3.1376
R1976 B.n889 B.t0 1.34497
R1977 B.n1050 B.t6 1.34497
R1978 B.n694 B.n693 1.24928
R1979 B.n531 B.n530 1.24928
R1980 B.n274 B.n273 1.24928
R1981 B.n294 B.n293 1.24928
R1982 VP.n13 VP.t2 280.058
R1983 VP.n7 VP.t5 245.719
R1984 VP.n40 VP.t1 245.719
R1985 VP.n47 VP.t7 245.719
R1986 VP.n55 VP.t3 245.719
R1987 VP.n29 VP.t0 245.719
R1988 VP.n21 VP.t4 245.719
R1989 VP.n14 VP.t6 245.719
R1990 VP.n31 VP.n7 181.852
R1991 VP.n56 VP.n55 181.852
R1992 VP.n30 VP.n29 181.852
R1993 VP.n15 VP.n12 161.3
R1994 VP.n17 VP.n16 161.3
R1995 VP.n18 VP.n11 161.3
R1996 VP.n20 VP.n19 161.3
R1997 VP.n22 VP.n10 161.3
R1998 VP.n24 VP.n23 161.3
R1999 VP.n25 VP.n9 161.3
R2000 VP.n27 VP.n26 161.3
R2001 VP.n28 VP.n8 161.3
R2002 VP.n54 VP.n0 161.3
R2003 VP.n53 VP.n52 161.3
R2004 VP.n51 VP.n1 161.3
R2005 VP.n50 VP.n49 161.3
R2006 VP.n48 VP.n2 161.3
R2007 VP.n46 VP.n45 161.3
R2008 VP.n44 VP.n3 161.3
R2009 VP.n43 VP.n42 161.3
R2010 VP.n41 VP.n4 161.3
R2011 VP.n39 VP.n38 161.3
R2012 VP.n37 VP.n5 161.3
R2013 VP.n36 VP.n35 161.3
R2014 VP.n34 VP.n6 161.3
R2015 VP.n33 VP.n32 161.3
R2016 VP.n42 VP.n3 56.5193
R2017 VP.n16 VP.n11 56.5193
R2018 VP.n31 VP.n30 53.0081
R2019 VP.n14 VP.n13 52.0405
R2020 VP.n35 VP.n5 43.4072
R2021 VP.n49 VP.n1 43.4072
R2022 VP.n23 VP.n9 43.4072
R2023 VP.n35 VP.n34 37.5796
R2024 VP.n53 VP.n1 37.5796
R2025 VP.n27 VP.n9 37.5796
R2026 VP.n34 VP.n33 24.4675
R2027 VP.n39 VP.n5 24.4675
R2028 VP.n42 VP.n41 24.4675
R2029 VP.n46 VP.n3 24.4675
R2030 VP.n49 VP.n48 24.4675
R2031 VP.n54 VP.n53 24.4675
R2032 VP.n28 VP.n27 24.4675
R2033 VP.n20 VP.n11 24.4675
R2034 VP.n23 VP.n22 24.4675
R2035 VP.n16 VP.n15 24.4675
R2036 VP.n41 VP.n40 17.6167
R2037 VP.n47 VP.n46 17.6167
R2038 VP.n21 VP.n20 17.6167
R2039 VP.n15 VP.n14 17.6167
R2040 VP.n13 VP.n12 12.2976
R2041 VP.n40 VP.n39 6.85126
R2042 VP.n48 VP.n47 6.85126
R2043 VP.n22 VP.n21 6.85126
R2044 VP.n33 VP.n7 3.91522
R2045 VP.n55 VP.n54 3.91522
R2046 VP.n29 VP.n28 3.91522
R2047 VP.n17 VP.n12 0.189894
R2048 VP.n18 VP.n17 0.189894
R2049 VP.n19 VP.n18 0.189894
R2050 VP.n19 VP.n10 0.189894
R2051 VP.n24 VP.n10 0.189894
R2052 VP.n25 VP.n24 0.189894
R2053 VP.n26 VP.n25 0.189894
R2054 VP.n26 VP.n8 0.189894
R2055 VP.n30 VP.n8 0.189894
R2056 VP.n32 VP.n31 0.189894
R2057 VP.n32 VP.n6 0.189894
R2058 VP.n36 VP.n6 0.189894
R2059 VP.n37 VP.n36 0.189894
R2060 VP.n38 VP.n37 0.189894
R2061 VP.n38 VP.n4 0.189894
R2062 VP.n43 VP.n4 0.189894
R2063 VP.n44 VP.n43 0.189894
R2064 VP.n45 VP.n44 0.189894
R2065 VP.n45 VP.n2 0.189894
R2066 VP.n50 VP.n2 0.189894
R2067 VP.n51 VP.n50 0.189894
R2068 VP.n52 VP.n51 0.189894
R2069 VP.n52 VP.n0 0.189894
R2070 VP.n56 VP.n0 0.189894
R2071 VP VP.n56 0.0516364
R2072 VDD1 VDD1.n0 60.6565
R2073 VDD1.n3 VDD1.n2 60.5429
R2074 VDD1.n3 VDD1.n1 60.5429
R2075 VDD1.n5 VDD1.n4 59.6413
R2076 VDD1.n5 VDD1.n3 49.5224
R2077 VDD1.n4 VDD1.t3 1.028
R2078 VDD1.n4 VDD1.t7 1.028
R2079 VDD1.n0 VDD1.t5 1.028
R2080 VDD1.n0 VDD1.t1 1.028
R2081 VDD1.n2 VDD1.t0 1.028
R2082 VDD1.n2 VDD1.t4 1.028
R2083 VDD1.n1 VDD1.t2 1.028
R2084 VDD1.n1 VDD1.t6 1.028
R2085 VDD1 VDD1.n5 0.899207
C0 VDD1 VN 0.150031f
C1 VDD1 VTAIL 11.0774f
C2 VTAIL VN 12.588901f
C3 VDD2 VDD1 1.40507f
C4 VDD2 VN 12.732201f
C5 VDD2 VTAIL 11.127f
C6 VDD1 VP 13.0249f
C7 VN VP 8.13818f
C8 VTAIL VP 12.603f
C9 VDD2 VP 0.443706f
C10 VDD2 B 5.225632f
C11 VDD1 B 5.58605f
C12 VTAIL B 14.280013f
C13 VN B 13.477871f
C14 VP B 11.779814f
C15 VDD1.t5 B 0.378389f
C16 VDD1.t1 B 0.378389f
C17 VDD1.n0 B 3.46196f
C18 VDD1.t2 B 0.378389f
C19 VDD1.t6 B 0.378389f
C20 VDD1.n1 B 3.46101f
C21 VDD1.t0 B 0.378389f
C22 VDD1.t4 B 0.378389f
C23 VDD1.n2 B 3.46101f
C24 VDD1.n3 B 3.36435f
C25 VDD1.t3 B 0.378389f
C26 VDD1.t7 B 0.378389f
C27 VDD1.n4 B 3.45436f
C28 VDD1.n5 B 3.27077f
C29 VP.n0 B 0.026259f
C30 VP.t3 B 2.63384f
C31 VP.n1 B 0.021533f
C32 VP.n2 B 0.026259f
C33 VP.t7 B 2.63384f
C34 VP.n3 B 0.038334f
C35 VP.n4 B 0.026259f
C36 VP.t1 B 2.63384f
C37 VP.n5 B 0.051258f
C38 VP.n6 B 0.026259f
C39 VP.t5 B 2.63384f
C40 VP.n7 B 0.98112f
C41 VP.n8 B 0.026259f
C42 VP.t0 B 2.63384f
C43 VP.n9 B 0.021533f
C44 VP.n10 B 0.026259f
C45 VP.t4 B 2.63384f
C46 VP.n11 B 0.038334f
C47 VP.n12 B 0.195385f
C48 VP.t6 B 2.63384f
C49 VP.t2 B 2.76219f
C50 VP.n13 B 0.978568f
C51 VP.n14 B 0.983002f
C52 VP.n15 B 0.042175f
C53 VP.n16 B 0.038334f
C54 VP.n17 B 0.026259f
C55 VP.n18 B 0.026259f
C56 VP.n19 B 0.026259f
C57 VP.n20 B 0.042175f
C58 VP.n21 B 0.917565f
C59 VP.n22 B 0.031544f
C60 VP.n23 B 0.051258f
C61 VP.n24 B 0.026259f
C62 VP.n25 B 0.026259f
C63 VP.n26 B 0.026259f
C64 VP.n27 B 0.052817f
C65 VP.n28 B 0.028644f
C66 VP.n29 B 0.98112f
C67 VP.n30 B 1.56484f
C68 VP.n31 B 1.58265f
C69 VP.n32 B 0.026259f
C70 VP.n33 B 0.028644f
C71 VP.n34 B 0.052817f
C72 VP.n35 B 0.021533f
C73 VP.n36 B 0.026259f
C74 VP.n37 B 0.026259f
C75 VP.n38 B 0.026259f
C76 VP.n39 B 0.031544f
C77 VP.n40 B 0.917565f
C78 VP.n41 B 0.042175f
C79 VP.n42 B 0.038334f
C80 VP.n43 B 0.026259f
C81 VP.n44 B 0.026259f
C82 VP.n45 B 0.026259f
C83 VP.n46 B 0.042175f
C84 VP.n47 B 0.917565f
C85 VP.n48 B 0.031544f
C86 VP.n49 B 0.051258f
C87 VP.n50 B 0.026259f
C88 VP.n51 B 0.026259f
C89 VP.n52 B 0.026259f
C90 VP.n53 B 0.052817f
C91 VP.n54 B 0.028644f
C92 VP.n55 B 0.98112f
C93 VP.n56 B 0.028448f
C94 VDD2.t1 B 0.375107f
C95 VDD2.t6 B 0.375107f
C96 VDD2.n0 B 3.43099f
C97 VDD2.t2 B 0.375107f
C98 VDD2.t7 B 0.375107f
C99 VDD2.n1 B 3.43099f
C100 VDD2.n2 B 3.28379f
C101 VDD2.t4 B 0.375107f
C102 VDD2.t0 B 0.375107f
C103 VDD2.n3 B 3.42441f
C104 VDD2.n4 B 3.21203f
C105 VDD2.t5 B 0.375107f
C106 VDD2.t3 B 0.375107f
C107 VDD2.n5 B 3.43094f
C108 VTAIL.t12 B 0.277096f
C109 VTAIL.t14 B 0.277096f
C110 VTAIL.n0 B 2.47151f
C111 VTAIL.n1 B 0.3023f
C112 VTAIL.t15 B 3.1583f
C113 VTAIL.n2 B 0.395354f
C114 VTAIL.t7 B 3.1583f
C115 VTAIL.n3 B 0.395354f
C116 VTAIL.t1 B 0.277096f
C117 VTAIL.t4 B 0.277096f
C118 VTAIL.n4 B 2.47151f
C119 VTAIL.n5 B 0.411102f
C120 VTAIL.t0 B 3.1583f
C121 VTAIL.n6 B 1.70124f
C122 VTAIL.t9 B 3.15831f
C123 VTAIL.n7 B 1.70123f
C124 VTAIL.t13 B 0.277096f
C125 VTAIL.t10 B 0.277096f
C126 VTAIL.n8 B 2.4715f
C127 VTAIL.n9 B 0.411107f
C128 VTAIL.t8 B 3.15831f
C129 VTAIL.n10 B 0.39535f
C130 VTAIL.t5 B 3.15831f
C131 VTAIL.n11 B 0.39535f
C132 VTAIL.t2 B 0.277096f
C133 VTAIL.t3 B 0.277096f
C134 VTAIL.n12 B 2.4715f
C135 VTAIL.n13 B 0.411107f
C136 VTAIL.t6 B 3.1583f
C137 VTAIL.n14 B 1.70124f
C138 VTAIL.t11 B 3.1583f
C139 VTAIL.n15 B 1.69782f
C140 VN.n0 B 0.025997f
C141 VN.t0 B 2.60754f
C142 VN.n1 B 0.021318f
C143 VN.n2 B 0.025997f
C144 VN.t5 B 2.60754f
C145 VN.n3 B 0.037951f
C146 VN.n4 B 0.193434f
C147 VN.t1 B 2.60754f
C148 VN.t6 B 2.7346f
C149 VN.n5 B 0.968796f
C150 VN.n6 B 0.973186f
C151 VN.n7 B 0.041754f
C152 VN.n8 B 0.037951f
C153 VN.n9 B 0.025997f
C154 VN.n10 B 0.025997f
C155 VN.n11 B 0.025997f
C156 VN.n12 B 0.041754f
C157 VN.n13 B 0.908401f
C158 VN.n14 B 0.031229f
C159 VN.n15 B 0.050746f
C160 VN.n16 B 0.025997f
C161 VN.n17 B 0.025997f
C162 VN.n18 B 0.025997f
C163 VN.n19 B 0.05229f
C164 VN.n20 B 0.028358f
C165 VN.n21 B 0.971322f
C166 VN.n22 B 0.028164f
C167 VN.n23 B 0.025997f
C168 VN.t3 B 2.60754f
C169 VN.n24 B 0.021318f
C170 VN.n25 B 0.025997f
C171 VN.t7 B 2.60754f
C172 VN.n26 B 0.037951f
C173 VN.n27 B 0.193434f
C174 VN.t2 B 2.60754f
C175 VN.t4 B 2.7346f
C176 VN.n28 B 0.968796f
C177 VN.n29 B 0.973186f
C178 VN.n30 B 0.041754f
C179 VN.n31 B 0.037951f
C180 VN.n32 B 0.025997f
C181 VN.n33 B 0.025997f
C182 VN.n34 B 0.025997f
C183 VN.n35 B 0.041754f
C184 VN.n36 B 0.908401f
C185 VN.n37 B 0.031229f
C186 VN.n38 B 0.050746f
C187 VN.n39 B 0.025997f
C188 VN.n40 B 0.025997f
C189 VN.n41 B 0.025997f
C190 VN.n42 B 0.05229f
C191 VN.n43 B 0.028358f
C192 VN.n44 B 0.971322f
C193 VN.n45 B 1.56607f
.ends

