* NGSPICE file created from diff_pair_sample_0575.ext - technology: sky130A

.subckt diff_pair_sample_0575 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t9 VP.t0 VDD1.t2 B.t5 sky130_fd_pr__nfet_01v8 ad=1.4553 pd=9.15 as=1.4553 ps=9.15 w=8.82 l=3.08
X1 VDD2.t5 VN.t0 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=3.4398 pd=18.42 as=1.4553 ps=9.15 w=8.82 l=3.08
X2 VDD2.t4 VN.t1 VTAIL.t10 B.t4 sky130_fd_pr__nfet_01v8 ad=3.4398 pd=18.42 as=1.4553 ps=9.15 w=8.82 l=3.08
X3 B.t19 B.t17 B.t18 B.t7 sky130_fd_pr__nfet_01v8 ad=3.4398 pd=18.42 as=0 ps=0 w=8.82 l=3.08
X4 VTAIL.t0 VN.t2 VDD2.t3 B.t0 sky130_fd_pr__nfet_01v8 ad=1.4553 pd=9.15 as=1.4553 ps=9.15 w=8.82 l=3.08
X5 VDD2.t2 VN.t3 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=1.4553 pd=9.15 as=3.4398 ps=18.42 w=8.82 l=3.08
X6 B.t16 B.t14 B.t15 B.t11 sky130_fd_pr__nfet_01v8 ad=3.4398 pd=18.42 as=0 ps=0 w=8.82 l=3.08
X7 VDD1.t1 VP.t1 VTAIL.t8 B.t4 sky130_fd_pr__nfet_01v8 ad=3.4398 pd=18.42 as=1.4553 ps=9.15 w=8.82 l=3.08
X8 VTAIL.t11 VN.t4 VDD2.t1 B.t5 sky130_fd_pr__nfet_01v8 ad=1.4553 pd=9.15 as=1.4553 ps=9.15 w=8.82 l=3.08
X9 VDD1.t0 VP.t2 VTAIL.t7 B.t1 sky130_fd_pr__nfet_01v8 ad=1.4553 pd=9.15 as=3.4398 ps=18.42 w=8.82 l=3.08
X10 VDD2.t0 VN.t5 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=1.4553 pd=9.15 as=3.4398 ps=18.42 w=8.82 l=3.08
X11 VDD1.t5 VP.t3 VTAIL.t6 B.t3 sky130_fd_pr__nfet_01v8 ad=1.4553 pd=9.15 as=3.4398 ps=18.42 w=8.82 l=3.08
X12 B.t13 B.t10 B.t12 B.t11 sky130_fd_pr__nfet_01v8 ad=3.4398 pd=18.42 as=0 ps=0 w=8.82 l=3.08
X13 VTAIL.t5 VP.t4 VDD1.t3 B.t0 sky130_fd_pr__nfet_01v8 ad=1.4553 pd=9.15 as=1.4553 ps=9.15 w=8.82 l=3.08
X14 VDD1.t4 VP.t5 VTAIL.t4 B.t2 sky130_fd_pr__nfet_01v8 ad=3.4398 pd=18.42 as=1.4553 ps=9.15 w=8.82 l=3.08
X15 B.t9 B.t6 B.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=3.4398 pd=18.42 as=0 ps=0 w=8.82 l=3.08
R0 VP.n13 VP.n10 161.3
R1 VP.n15 VP.n14 161.3
R2 VP.n16 VP.n9 161.3
R3 VP.n18 VP.n17 161.3
R4 VP.n19 VP.n8 161.3
R5 VP.n21 VP.n20 161.3
R6 VP.n44 VP.n43 161.3
R7 VP.n42 VP.n1 161.3
R8 VP.n41 VP.n40 161.3
R9 VP.n39 VP.n2 161.3
R10 VP.n38 VP.n37 161.3
R11 VP.n36 VP.n3 161.3
R12 VP.n35 VP.n34 161.3
R13 VP.n33 VP.n4 161.3
R14 VP.n32 VP.n31 161.3
R15 VP.n30 VP.n5 161.3
R16 VP.n29 VP.n28 161.3
R17 VP.n27 VP.n6 161.3
R18 VP.n26 VP.n25 161.3
R19 VP.n11 VP.t1 102.337
R20 VP.n24 VP.n23 69.9294
R21 VP.n45 VP.n0 69.9294
R22 VP.n22 VP.n7 69.9294
R23 VP.n35 VP.t4 69.0141
R24 VP.n24 VP.t5 69.0141
R25 VP.n0 VP.t2 69.0141
R26 VP.n12 VP.t0 69.0141
R27 VP.n7 VP.t3 69.0141
R28 VP.n30 VP.n29 56.4773
R29 VP.n41 VP.n2 56.4773
R30 VP.n18 VP.n9 56.4773
R31 VP.n12 VP.n11 49.2934
R32 VP.n23 VP.n22 48.2908
R33 VP.n25 VP.n6 24.3439
R34 VP.n29 VP.n6 24.3439
R35 VP.n31 VP.n30 24.3439
R36 VP.n31 VP.n4 24.3439
R37 VP.n35 VP.n4 24.3439
R38 VP.n36 VP.n35 24.3439
R39 VP.n37 VP.n36 24.3439
R40 VP.n37 VP.n2 24.3439
R41 VP.n42 VP.n41 24.3439
R42 VP.n43 VP.n42 24.3439
R43 VP.n19 VP.n18 24.3439
R44 VP.n20 VP.n19 24.3439
R45 VP.n13 VP.n12 24.3439
R46 VP.n14 VP.n13 24.3439
R47 VP.n14 VP.n9 24.3439
R48 VP.n25 VP.n24 19.9621
R49 VP.n43 VP.n0 19.9621
R50 VP.n20 VP.n7 19.9621
R51 VP.n11 VP.n10 3.92639
R52 VP.n22 VP.n21 0.355081
R53 VP.n26 VP.n23 0.355081
R54 VP.n45 VP.n44 0.355081
R55 VP VP.n45 0.26685
R56 VP.n15 VP.n10 0.189894
R57 VP.n16 VP.n15 0.189894
R58 VP.n17 VP.n16 0.189894
R59 VP.n17 VP.n8 0.189894
R60 VP.n21 VP.n8 0.189894
R61 VP.n27 VP.n26 0.189894
R62 VP.n28 VP.n27 0.189894
R63 VP.n28 VP.n5 0.189894
R64 VP.n32 VP.n5 0.189894
R65 VP.n33 VP.n32 0.189894
R66 VP.n34 VP.n33 0.189894
R67 VP.n34 VP.n3 0.189894
R68 VP.n38 VP.n3 0.189894
R69 VP.n39 VP.n38 0.189894
R70 VP.n40 VP.n39 0.189894
R71 VP.n40 VP.n1 0.189894
R72 VP.n44 VP.n1 0.189894
R73 VDD1.n42 VDD1.n0 289.615
R74 VDD1.n89 VDD1.n47 289.615
R75 VDD1.n43 VDD1.n42 185
R76 VDD1.n41 VDD1.n40 185
R77 VDD1.n4 VDD1.n3 185
R78 VDD1.n35 VDD1.n34 185
R79 VDD1.n33 VDD1.n32 185
R80 VDD1.n8 VDD1.n7 185
R81 VDD1.n27 VDD1.n26 185
R82 VDD1.n25 VDD1.n24 185
R83 VDD1.n12 VDD1.n11 185
R84 VDD1.n19 VDD1.n18 185
R85 VDD1.n17 VDD1.n16 185
R86 VDD1.n64 VDD1.n63 185
R87 VDD1.n66 VDD1.n65 185
R88 VDD1.n59 VDD1.n58 185
R89 VDD1.n72 VDD1.n71 185
R90 VDD1.n74 VDD1.n73 185
R91 VDD1.n55 VDD1.n54 185
R92 VDD1.n80 VDD1.n79 185
R93 VDD1.n82 VDD1.n81 185
R94 VDD1.n51 VDD1.n50 185
R95 VDD1.n88 VDD1.n87 185
R96 VDD1.n90 VDD1.n89 185
R97 VDD1.n15 VDD1.t1 147.659
R98 VDD1.n62 VDD1.t4 147.659
R99 VDD1.n42 VDD1.n41 104.615
R100 VDD1.n41 VDD1.n3 104.615
R101 VDD1.n34 VDD1.n3 104.615
R102 VDD1.n34 VDD1.n33 104.615
R103 VDD1.n33 VDD1.n7 104.615
R104 VDD1.n26 VDD1.n7 104.615
R105 VDD1.n26 VDD1.n25 104.615
R106 VDD1.n25 VDD1.n11 104.615
R107 VDD1.n18 VDD1.n11 104.615
R108 VDD1.n18 VDD1.n17 104.615
R109 VDD1.n65 VDD1.n64 104.615
R110 VDD1.n65 VDD1.n58 104.615
R111 VDD1.n72 VDD1.n58 104.615
R112 VDD1.n73 VDD1.n72 104.615
R113 VDD1.n73 VDD1.n54 104.615
R114 VDD1.n80 VDD1.n54 104.615
R115 VDD1.n81 VDD1.n80 104.615
R116 VDD1.n81 VDD1.n50 104.615
R117 VDD1.n88 VDD1.n50 104.615
R118 VDD1.n89 VDD1.n88 104.615
R119 VDD1.n95 VDD1.n94 63.4539
R120 VDD1.n97 VDD1.n96 62.7745
R121 VDD1.n17 VDD1.t1 52.3082
R122 VDD1.n64 VDD1.t4 52.3082
R123 VDD1 VDD1.n46 49.9634
R124 VDD1.n95 VDD1.n93 49.8499
R125 VDD1.n97 VDD1.n95 42.9255
R126 VDD1.n16 VDD1.n15 15.6677
R127 VDD1.n63 VDD1.n62 15.6677
R128 VDD1.n19 VDD1.n14 12.8005
R129 VDD1.n66 VDD1.n61 12.8005
R130 VDD1.n20 VDD1.n12 12.0247
R131 VDD1.n67 VDD1.n59 12.0247
R132 VDD1.n24 VDD1.n23 11.249
R133 VDD1.n71 VDD1.n70 11.249
R134 VDD1.n27 VDD1.n10 10.4732
R135 VDD1.n74 VDD1.n57 10.4732
R136 VDD1.n28 VDD1.n8 9.69747
R137 VDD1.n75 VDD1.n55 9.69747
R138 VDD1.n46 VDD1.n45 9.45567
R139 VDD1.n93 VDD1.n92 9.45567
R140 VDD1.n2 VDD1.n1 9.3005
R141 VDD1.n45 VDD1.n44 9.3005
R142 VDD1.n39 VDD1.n38 9.3005
R143 VDD1.n37 VDD1.n36 9.3005
R144 VDD1.n6 VDD1.n5 9.3005
R145 VDD1.n31 VDD1.n30 9.3005
R146 VDD1.n29 VDD1.n28 9.3005
R147 VDD1.n10 VDD1.n9 9.3005
R148 VDD1.n23 VDD1.n22 9.3005
R149 VDD1.n21 VDD1.n20 9.3005
R150 VDD1.n14 VDD1.n13 9.3005
R151 VDD1.n86 VDD1.n85 9.3005
R152 VDD1.n49 VDD1.n48 9.3005
R153 VDD1.n92 VDD1.n91 9.3005
R154 VDD1.n53 VDD1.n52 9.3005
R155 VDD1.n78 VDD1.n77 9.3005
R156 VDD1.n76 VDD1.n75 9.3005
R157 VDD1.n57 VDD1.n56 9.3005
R158 VDD1.n70 VDD1.n69 9.3005
R159 VDD1.n68 VDD1.n67 9.3005
R160 VDD1.n61 VDD1.n60 9.3005
R161 VDD1.n84 VDD1.n83 9.3005
R162 VDD1.n46 VDD1.n0 8.92171
R163 VDD1.n32 VDD1.n31 8.92171
R164 VDD1.n79 VDD1.n78 8.92171
R165 VDD1.n93 VDD1.n47 8.92171
R166 VDD1.n44 VDD1.n43 8.14595
R167 VDD1.n35 VDD1.n6 8.14595
R168 VDD1.n82 VDD1.n53 8.14595
R169 VDD1.n91 VDD1.n90 8.14595
R170 VDD1.n40 VDD1.n2 7.3702
R171 VDD1.n36 VDD1.n4 7.3702
R172 VDD1.n83 VDD1.n51 7.3702
R173 VDD1.n87 VDD1.n49 7.3702
R174 VDD1.n40 VDD1.n39 6.59444
R175 VDD1.n39 VDD1.n4 6.59444
R176 VDD1.n86 VDD1.n51 6.59444
R177 VDD1.n87 VDD1.n86 6.59444
R178 VDD1.n43 VDD1.n2 5.81868
R179 VDD1.n36 VDD1.n35 5.81868
R180 VDD1.n83 VDD1.n82 5.81868
R181 VDD1.n90 VDD1.n49 5.81868
R182 VDD1.n44 VDD1.n0 5.04292
R183 VDD1.n32 VDD1.n6 5.04292
R184 VDD1.n79 VDD1.n53 5.04292
R185 VDD1.n91 VDD1.n47 5.04292
R186 VDD1.n15 VDD1.n13 4.38563
R187 VDD1.n62 VDD1.n60 4.38563
R188 VDD1.n31 VDD1.n8 4.26717
R189 VDD1.n78 VDD1.n55 4.26717
R190 VDD1.n28 VDD1.n27 3.49141
R191 VDD1.n75 VDD1.n74 3.49141
R192 VDD1.n24 VDD1.n10 2.71565
R193 VDD1.n71 VDD1.n57 2.71565
R194 VDD1.n96 VDD1.t2 2.2454
R195 VDD1.n96 VDD1.t5 2.2454
R196 VDD1.n94 VDD1.t3 2.2454
R197 VDD1.n94 VDD1.t0 2.2454
R198 VDD1.n23 VDD1.n12 1.93989
R199 VDD1.n70 VDD1.n59 1.93989
R200 VDD1.n20 VDD1.n19 1.16414
R201 VDD1.n67 VDD1.n66 1.16414
R202 VDD1 VDD1.n97 0.677224
R203 VDD1.n16 VDD1.n14 0.388379
R204 VDD1.n63 VDD1.n61 0.388379
R205 VDD1.n45 VDD1.n1 0.155672
R206 VDD1.n38 VDD1.n1 0.155672
R207 VDD1.n38 VDD1.n37 0.155672
R208 VDD1.n37 VDD1.n5 0.155672
R209 VDD1.n30 VDD1.n5 0.155672
R210 VDD1.n30 VDD1.n29 0.155672
R211 VDD1.n29 VDD1.n9 0.155672
R212 VDD1.n22 VDD1.n9 0.155672
R213 VDD1.n22 VDD1.n21 0.155672
R214 VDD1.n21 VDD1.n13 0.155672
R215 VDD1.n68 VDD1.n60 0.155672
R216 VDD1.n69 VDD1.n68 0.155672
R217 VDD1.n69 VDD1.n56 0.155672
R218 VDD1.n76 VDD1.n56 0.155672
R219 VDD1.n77 VDD1.n76 0.155672
R220 VDD1.n77 VDD1.n52 0.155672
R221 VDD1.n84 VDD1.n52 0.155672
R222 VDD1.n85 VDD1.n84 0.155672
R223 VDD1.n85 VDD1.n48 0.155672
R224 VDD1.n92 VDD1.n48 0.155672
R225 VTAIL.n194 VTAIL.n152 289.615
R226 VTAIL.n44 VTAIL.n2 289.615
R227 VTAIL.n146 VTAIL.n104 289.615
R228 VTAIL.n96 VTAIL.n54 289.615
R229 VTAIL.n169 VTAIL.n168 185
R230 VTAIL.n171 VTAIL.n170 185
R231 VTAIL.n164 VTAIL.n163 185
R232 VTAIL.n177 VTAIL.n176 185
R233 VTAIL.n179 VTAIL.n178 185
R234 VTAIL.n160 VTAIL.n159 185
R235 VTAIL.n185 VTAIL.n184 185
R236 VTAIL.n187 VTAIL.n186 185
R237 VTAIL.n156 VTAIL.n155 185
R238 VTAIL.n193 VTAIL.n192 185
R239 VTAIL.n195 VTAIL.n194 185
R240 VTAIL.n19 VTAIL.n18 185
R241 VTAIL.n21 VTAIL.n20 185
R242 VTAIL.n14 VTAIL.n13 185
R243 VTAIL.n27 VTAIL.n26 185
R244 VTAIL.n29 VTAIL.n28 185
R245 VTAIL.n10 VTAIL.n9 185
R246 VTAIL.n35 VTAIL.n34 185
R247 VTAIL.n37 VTAIL.n36 185
R248 VTAIL.n6 VTAIL.n5 185
R249 VTAIL.n43 VTAIL.n42 185
R250 VTAIL.n45 VTAIL.n44 185
R251 VTAIL.n147 VTAIL.n146 185
R252 VTAIL.n145 VTAIL.n144 185
R253 VTAIL.n108 VTAIL.n107 185
R254 VTAIL.n139 VTAIL.n138 185
R255 VTAIL.n137 VTAIL.n136 185
R256 VTAIL.n112 VTAIL.n111 185
R257 VTAIL.n131 VTAIL.n130 185
R258 VTAIL.n129 VTAIL.n128 185
R259 VTAIL.n116 VTAIL.n115 185
R260 VTAIL.n123 VTAIL.n122 185
R261 VTAIL.n121 VTAIL.n120 185
R262 VTAIL.n97 VTAIL.n96 185
R263 VTAIL.n95 VTAIL.n94 185
R264 VTAIL.n58 VTAIL.n57 185
R265 VTAIL.n89 VTAIL.n88 185
R266 VTAIL.n87 VTAIL.n86 185
R267 VTAIL.n62 VTAIL.n61 185
R268 VTAIL.n81 VTAIL.n80 185
R269 VTAIL.n79 VTAIL.n78 185
R270 VTAIL.n66 VTAIL.n65 185
R271 VTAIL.n73 VTAIL.n72 185
R272 VTAIL.n71 VTAIL.n70 185
R273 VTAIL.n69 VTAIL.t1 147.659
R274 VTAIL.n167 VTAIL.t3 147.659
R275 VTAIL.n17 VTAIL.t7 147.659
R276 VTAIL.n119 VTAIL.t6 147.659
R277 VTAIL.n170 VTAIL.n169 104.615
R278 VTAIL.n170 VTAIL.n163 104.615
R279 VTAIL.n177 VTAIL.n163 104.615
R280 VTAIL.n178 VTAIL.n177 104.615
R281 VTAIL.n178 VTAIL.n159 104.615
R282 VTAIL.n185 VTAIL.n159 104.615
R283 VTAIL.n186 VTAIL.n185 104.615
R284 VTAIL.n186 VTAIL.n155 104.615
R285 VTAIL.n193 VTAIL.n155 104.615
R286 VTAIL.n194 VTAIL.n193 104.615
R287 VTAIL.n20 VTAIL.n19 104.615
R288 VTAIL.n20 VTAIL.n13 104.615
R289 VTAIL.n27 VTAIL.n13 104.615
R290 VTAIL.n28 VTAIL.n27 104.615
R291 VTAIL.n28 VTAIL.n9 104.615
R292 VTAIL.n35 VTAIL.n9 104.615
R293 VTAIL.n36 VTAIL.n35 104.615
R294 VTAIL.n36 VTAIL.n5 104.615
R295 VTAIL.n43 VTAIL.n5 104.615
R296 VTAIL.n44 VTAIL.n43 104.615
R297 VTAIL.n146 VTAIL.n145 104.615
R298 VTAIL.n145 VTAIL.n107 104.615
R299 VTAIL.n138 VTAIL.n107 104.615
R300 VTAIL.n138 VTAIL.n137 104.615
R301 VTAIL.n137 VTAIL.n111 104.615
R302 VTAIL.n130 VTAIL.n111 104.615
R303 VTAIL.n130 VTAIL.n129 104.615
R304 VTAIL.n129 VTAIL.n115 104.615
R305 VTAIL.n122 VTAIL.n115 104.615
R306 VTAIL.n122 VTAIL.n121 104.615
R307 VTAIL.n96 VTAIL.n95 104.615
R308 VTAIL.n95 VTAIL.n57 104.615
R309 VTAIL.n88 VTAIL.n57 104.615
R310 VTAIL.n88 VTAIL.n87 104.615
R311 VTAIL.n87 VTAIL.n61 104.615
R312 VTAIL.n80 VTAIL.n61 104.615
R313 VTAIL.n80 VTAIL.n79 104.615
R314 VTAIL.n79 VTAIL.n65 104.615
R315 VTAIL.n72 VTAIL.n65 104.615
R316 VTAIL.n72 VTAIL.n71 104.615
R317 VTAIL.n169 VTAIL.t3 52.3082
R318 VTAIL.n19 VTAIL.t7 52.3082
R319 VTAIL.n121 VTAIL.t6 52.3082
R320 VTAIL.n71 VTAIL.t1 52.3082
R321 VTAIL.n103 VTAIL.n102 46.0957
R322 VTAIL.n53 VTAIL.n52 46.0957
R323 VTAIL.n1 VTAIL.n0 46.0956
R324 VTAIL.n51 VTAIL.n50 46.0956
R325 VTAIL.n199 VTAIL.n198 31.0217
R326 VTAIL.n49 VTAIL.n48 31.0217
R327 VTAIL.n151 VTAIL.n150 31.0217
R328 VTAIL.n101 VTAIL.n100 31.0217
R329 VTAIL.n53 VTAIL.n51 25.8496
R330 VTAIL.n199 VTAIL.n151 22.91
R331 VTAIL.n168 VTAIL.n167 15.6677
R332 VTAIL.n18 VTAIL.n17 15.6677
R333 VTAIL.n120 VTAIL.n119 15.6677
R334 VTAIL.n70 VTAIL.n69 15.6677
R335 VTAIL.n171 VTAIL.n166 12.8005
R336 VTAIL.n21 VTAIL.n16 12.8005
R337 VTAIL.n123 VTAIL.n118 12.8005
R338 VTAIL.n73 VTAIL.n68 12.8005
R339 VTAIL.n172 VTAIL.n164 12.0247
R340 VTAIL.n22 VTAIL.n14 12.0247
R341 VTAIL.n124 VTAIL.n116 12.0247
R342 VTAIL.n74 VTAIL.n66 12.0247
R343 VTAIL.n176 VTAIL.n175 11.249
R344 VTAIL.n26 VTAIL.n25 11.249
R345 VTAIL.n128 VTAIL.n127 11.249
R346 VTAIL.n78 VTAIL.n77 11.249
R347 VTAIL.n179 VTAIL.n162 10.4732
R348 VTAIL.n29 VTAIL.n12 10.4732
R349 VTAIL.n131 VTAIL.n114 10.4732
R350 VTAIL.n81 VTAIL.n64 10.4732
R351 VTAIL.n180 VTAIL.n160 9.69747
R352 VTAIL.n30 VTAIL.n10 9.69747
R353 VTAIL.n132 VTAIL.n112 9.69747
R354 VTAIL.n82 VTAIL.n62 9.69747
R355 VTAIL.n198 VTAIL.n197 9.45567
R356 VTAIL.n48 VTAIL.n47 9.45567
R357 VTAIL.n150 VTAIL.n149 9.45567
R358 VTAIL.n100 VTAIL.n99 9.45567
R359 VTAIL.n191 VTAIL.n190 9.3005
R360 VTAIL.n154 VTAIL.n153 9.3005
R361 VTAIL.n197 VTAIL.n196 9.3005
R362 VTAIL.n158 VTAIL.n157 9.3005
R363 VTAIL.n183 VTAIL.n182 9.3005
R364 VTAIL.n181 VTAIL.n180 9.3005
R365 VTAIL.n162 VTAIL.n161 9.3005
R366 VTAIL.n175 VTAIL.n174 9.3005
R367 VTAIL.n173 VTAIL.n172 9.3005
R368 VTAIL.n166 VTAIL.n165 9.3005
R369 VTAIL.n189 VTAIL.n188 9.3005
R370 VTAIL.n41 VTAIL.n40 9.3005
R371 VTAIL.n4 VTAIL.n3 9.3005
R372 VTAIL.n47 VTAIL.n46 9.3005
R373 VTAIL.n8 VTAIL.n7 9.3005
R374 VTAIL.n33 VTAIL.n32 9.3005
R375 VTAIL.n31 VTAIL.n30 9.3005
R376 VTAIL.n12 VTAIL.n11 9.3005
R377 VTAIL.n25 VTAIL.n24 9.3005
R378 VTAIL.n23 VTAIL.n22 9.3005
R379 VTAIL.n16 VTAIL.n15 9.3005
R380 VTAIL.n39 VTAIL.n38 9.3005
R381 VTAIL.n106 VTAIL.n105 9.3005
R382 VTAIL.n143 VTAIL.n142 9.3005
R383 VTAIL.n141 VTAIL.n140 9.3005
R384 VTAIL.n110 VTAIL.n109 9.3005
R385 VTAIL.n135 VTAIL.n134 9.3005
R386 VTAIL.n133 VTAIL.n132 9.3005
R387 VTAIL.n114 VTAIL.n113 9.3005
R388 VTAIL.n127 VTAIL.n126 9.3005
R389 VTAIL.n125 VTAIL.n124 9.3005
R390 VTAIL.n118 VTAIL.n117 9.3005
R391 VTAIL.n149 VTAIL.n148 9.3005
R392 VTAIL.n56 VTAIL.n55 9.3005
R393 VTAIL.n99 VTAIL.n98 9.3005
R394 VTAIL.n93 VTAIL.n92 9.3005
R395 VTAIL.n91 VTAIL.n90 9.3005
R396 VTAIL.n60 VTAIL.n59 9.3005
R397 VTAIL.n85 VTAIL.n84 9.3005
R398 VTAIL.n83 VTAIL.n82 9.3005
R399 VTAIL.n64 VTAIL.n63 9.3005
R400 VTAIL.n77 VTAIL.n76 9.3005
R401 VTAIL.n75 VTAIL.n74 9.3005
R402 VTAIL.n68 VTAIL.n67 9.3005
R403 VTAIL.n184 VTAIL.n183 8.92171
R404 VTAIL.n198 VTAIL.n152 8.92171
R405 VTAIL.n34 VTAIL.n33 8.92171
R406 VTAIL.n48 VTAIL.n2 8.92171
R407 VTAIL.n150 VTAIL.n104 8.92171
R408 VTAIL.n136 VTAIL.n135 8.92171
R409 VTAIL.n100 VTAIL.n54 8.92171
R410 VTAIL.n86 VTAIL.n85 8.92171
R411 VTAIL.n187 VTAIL.n158 8.14595
R412 VTAIL.n196 VTAIL.n195 8.14595
R413 VTAIL.n37 VTAIL.n8 8.14595
R414 VTAIL.n46 VTAIL.n45 8.14595
R415 VTAIL.n148 VTAIL.n147 8.14595
R416 VTAIL.n139 VTAIL.n110 8.14595
R417 VTAIL.n98 VTAIL.n97 8.14595
R418 VTAIL.n89 VTAIL.n60 8.14595
R419 VTAIL.n188 VTAIL.n156 7.3702
R420 VTAIL.n192 VTAIL.n154 7.3702
R421 VTAIL.n38 VTAIL.n6 7.3702
R422 VTAIL.n42 VTAIL.n4 7.3702
R423 VTAIL.n144 VTAIL.n106 7.3702
R424 VTAIL.n140 VTAIL.n108 7.3702
R425 VTAIL.n94 VTAIL.n56 7.3702
R426 VTAIL.n90 VTAIL.n58 7.3702
R427 VTAIL.n191 VTAIL.n156 6.59444
R428 VTAIL.n192 VTAIL.n191 6.59444
R429 VTAIL.n41 VTAIL.n6 6.59444
R430 VTAIL.n42 VTAIL.n41 6.59444
R431 VTAIL.n144 VTAIL.n143 6.59444
R432 VTAIL.n143 VTAIL.n108 6.59444
R433 VTAIL.n94 VTAIL.n93 6.59444
R434 VTAIL.n93 VTAIL.n58 6.59444
R435 VTAIL.n188 VTAIL.n187 5.81868
R436 VTAIL.n195 VTAIL.n154 5.81868
R437 VTAIL.n38 VTAIL.n37 5.81868
R438 VTAIL.n45 VTAIL.n4 5.81868
R439 VTAIL.n147 VTAIL.n106 5.81868
R440 VTAIL.n140 VTAIL.n139 5.81868
R441 VTAIL.n97 VTAIL.n56 5.81868
R442 VTAIL.n90 VTAIL.n89 5.81868
R443 VTAIL.n184 VTAIL.n158 5.04292
R444 VTAIL.n196 VTAIL.n152 5.04292
R445 VTAIL.n34 VTAIL.n8 5.04292
R446 VTAIL.n46 VTAIL.n2 5.04292
R447 VTAIL.n148 VTAIL.n104 5.04292
R448 VTAIL.n136 VTAIL.n110 5.04292
R449 VTAIL.n98 VTAIL.n54 5.04292
R450 VTAIL.n86 VTAIL.n60 5.04292
R451 VTAIL.n167 VTAIL.n165 4.38563
R452 VTAIL.n17 VTAIL.n15 4.38563
R453 VTAIL.n119 VTAIL.n117 4.38563
R454 VTAIL.n69 VTAIL.n67 4.38563
R455 VTAIL.n183 VTAIL.n160 4.26717
R456 VTAIL.n33 VTAIL.n10 4.26717
R457 VTAIL.n135 VTAIL.n112 4.26717
R458 VTAIL.n85 VTAIL.n62 4.26717
R459 VTAIL.n180 VTAIL.n179 3.49141
R460 VTAIL.n30 VTAIL.n29 3.49141
R461 VTAIL.n132 VTAIL.n131 3.49141
R462 VTAIL.n82 VTAIL.n81 3.49141
R463 VTAIL.n101 VTAIL.n53 2.94016
R464 VTAIL.n151 VTAIL.n103 2.94016
R465 VTAIL.n51 VTAIL.n49 2.94016
R466 VTAIL.n176 VTAIL.n162 2.71565
R467 VTAIL.n26 VTAIL.n12 2.71565
R468 VTAIL.n128 VTAIL.n114 2.71565
R469 VTAIL.n78 VTAIL.n64 2.71565
R470 VTAIL.n0 VTAIL.t10 2.2454
R471 VTAIL.n0 VTAIL.t11 2.2454
R472 VTAIL.n50 VTAIL.t4 2.2454
R473 VTAIL.n50 VTAIL.t5 2.2454
R474 VTAIL.n102 VTAIL.t8 2.2454
R475 VTAIL.n102 VTAIL.t9 2.2454
R476 VTAIL.n52 VTAIL.t2 2.2454
R477 VTAIL.n52 VTAIL.t0 2.2454
R478 VTAIL VTAIL.n199 2.14705
R479 VTAIL.n103 VTAIL.n101 1.94016
R480 VTAIL.n49 VTAIL.n1 1.94016
R481 VTAIL.n175 VTAIL.n164 1.93989
R482 VTAIL.n25 VTAIL.n14 1.93989
R483 VTAIL.n127 VTAIL.n116 1.93989
R484 VTAIL.n77 VTAIL.n66 1.93989
R485 VTAIL.n172 VTAIL.n171 1.16414
R486 VTAIL.n22 VTAIL.n21 1.16414
R487 VTAIL.n124 VTAIL.n123 1.16414
R488 VTAIL.n74 VTAIL.n73 1.16414
R489 VTAIL VTAIL.n1 0.793603
R490 VTAIL.n168 VTAIL.n166 0.388379
R491 VTAIL.n18 VTAIL.n16 0.388379
R492 VTAIL.n120 VTAIL.n118 0.388379
R493 VTAIL.n70 VTAIL.n68 0.388379
R494 VTAIL.n173 VTAIL.n165 0.155672
R495 VTAIL.n174 VTAIL.n173 0.155672
R496 VTAIL.n174 VTAIL.n161 0.155672
R497 VTAIL.n181 VTAIL.n161 0.155672
R498 VTAIL.n182 VTAIL.n181 0.155672
R499 VTAIL.n182 VTAIL.n157 0.155672
R500 VTAIL.n189 VTAIL.n157 0.155672
R501 VTAIL.n190 VTAIL.n189 0.155672
R502 VTAIL.n190 VTAIL.n153 0.155672
R503 VTAIL.n197 VTAIL.n153 0.155672
R504 VTAIL.n23 VTAIL.n15 0.155672
R505 VTAIL.n24 VTAIL.n23 0.155672
R506 VTAIL.n24 VTAIL.n11 0.155672
R507 VTAIL.n31 VTAIL.n11 0.155672
R508 VTAIL.n32 VTAIL.n31 0.155672
R509 VTAIL.n32 VTAIL.n7 0.155672
R510 VTAIL.n39 VTAIL.n7 0.155672
R511 VTAIL.n40 VTAIL.n39 0.155672
R512 VTAIL.n40 VTAIL.n3 0.155672
R513 VTAIL.n47 VTAIL.n3 0.155672
R514 VTAIL.n149 VTAIL.n105 0.155672
R515 VTAIL.n142 VTAIL.n105 0.155672
R516 VTAIL.n142 VTAIL.n141 0.155672
R517 VTAIL.n141 VTAIL.n109 0.155672
R518 VTAIL.n134 VTAIL.n109 0.155672
R519 VTAIL.n134 VTAIL.n133 0.155672
R520 VTAIL.n133 VTAIL.n113 0.155672
R521 VTAIL.n126 VTAIL.n113 0.155672
R522 VTAIL.n126 VTAIL.n125 0.155672
R523 VTAIL.n125 VTAIL.n117 0.155672
R524 VTAIL.n99 VTAIL.n55 0.155672
R525 VTAIL.n92 VTAIL.n55 0.155672
R526 VTAIL.n92 VTAIL.n91 0.155672
R527 VTAIL.n91 VTAIL.n59 0.155672
R528 VTAIL.n84 VTAIL.n59 0.155672
R529 VTAIL.n84 VTAIL.n83 0.155672
R530 VTAIL.n83 VTAIL.n63 0.155672
R531 VTAIL.n76 VTAIL.n63 0.155672
R532 VTAIL.n76 VTAIL.n75 0.155672
R533 VTAIL.n75 VTAIL.n67 0.155672
R534 B.n766 B.n765 585
R535 B.n275 B.n126 585
R536 B.n274 B.n273 585
R537 B.n272 B.n271 585
R538 B.n270 B.n269 585
R539 B.n268 B.n267 585
R540 B.n266 B.n265 585
R541 B.n264 B.n263 585
R542 B.n262 B.n261 585
R543 B.n260 B.n259 585
R544 B.n258 B.n257 585
R545 B.n256 B.n255 585
R546 B.n254 B.n253 585
R547 B.n252 B.n251 585
R548 B.n250 B.n249 585
R549 B.n248 B.n247 585
R550 B.n246 B.n245 585
R551 B.n244 B.n243 585
R552 B.n242 B.n241 585
R553 B.n240 B.n239 585
R554 B.n238 B.n237 585
R555 B.n236 B.n235 585
R556 B.n234 B.n233 585
R557 B.n232 B.n231 585
R558 B.n230 B.n229 585
R559 B.n228 B.n227 585
R560 B.n226 B.n225 585
R561 B.n224 B.n223 585
R562 B.n222 B.n221 585
R563 B.n220 B.n219 585
R564 B.n218 B.n217 585
R565 B.n216 B.n215 585
R566 B.n214 B.n213 585
R567 B.n212 B.n211 585
R568 B.n210 B.n209 585
R569 B.n208 B.n207 585
R570 B.n206 B.n205 585
R571 B.n204 B.n203 585
R572 B.n202 B.n201 585
R573 B.n200 B.n199 585
R574 B.n198 B.n197 585
R575 B.n196 B.n195 585
R576 B.n194 B.n193 585
R577 B.n192 B.n191 585
R578 B.n190 B.n189 585
R579 B.n188 B.n187 585
R580 B.n186 B.n185 585
R581 B.n184 B.n183 585
R582 B.n182 B.n181 585
R583 B.n180 B.n179 585
R584 B.n178 B.n177 585
R585 B.n176 B.n175 585
R586 B.n174 B.n173 585
R587 B.n172 B.n171 585
R588 B.n170 B.n169 585
R589 B.n168 B.n167 585
R590 B.n166 B.n165 585
R591 B.n164 B.n163 585
R592 B.n162 B.n161 585
R593 B.n160 B.n159 585
R594 B.n158 B.n157 585
R595 B.n156 B.n155 585
R596 B.n154 B.n153 585
R597 B.n152 B.n151 585
R598 B.n150 B.n149 585
R599 B.n148 B.n147 585
R600 B.n146 B.n145 585
R601 B.n144 B.n143 585
R602 B.n142 B.n141 585
R603 B.n140 B.n139 585
R604 B.n138 B.n137 585
R605 B.n136 B.n135 585
R606 B.n134 B.n133 585
R607 B.n88 B.n87 585
R608 B.n764 B.n89 585
R609 B.n769 B.n89 585
R610 B.n763 B.n762 585
R611 B.n762 B.n85 585
R612 B.n761 B.n84 585
R613 B.n775 B.n84 585
R614 B.n760 B.n83 585
R615 B.n776 B.n83 585
R616 B.n759 B.n82 585
R617 B.n777 B.n82 585
R618 B.n758 B.n757 585
R619 B.n757 B.n78 585
R620 B.n756 B.n77 585
R621 B.n783 B.n77 585
R622 B.n755 B.n76 585
R623 B.n784 B.n76 585
R624 B.n754 B.n75 585
R625 B.n785 B.n75 585
R626 B.n753 B.n752 585
R627 B.n752 B.n71 585
R628 B.n751 B.n70 585
R629 B.n791 B.n70 585
R630 B.n750 B.n69 585
R631 B.n792 B.n69 585
R632 B.n749 B.n68 585
R633 B.n793 B.n68 585
R634 B.n748 B.n747 585
R635 B.n747 B.n64 585
R636 B.n746 B.n63 585
R637 B.n799 B.n63 585
R638 B.n745 B.n62 585
R639 B.n800 B.n62 585
R640 B.n744 B.n61 585
R641 B.n801 B.n61 585
R642 B.n743 B.n742 585
R643 B.n742 B.n57 585
R644 B.n741 B.n56 585
R645 B.n807 B.n56 585
R646 B.n740 B.n55 585
R647 B.n808 B.n55 585
R648 B.n739 B.n54 585
R649 B.n809 B.n54 585
R650 B.n738 B.n737 585
R651 B.n737 B.n53 585
R652 B.n736 B.n49 585
R653 B.n815 B.n49 585
R654 B.n735 B.n48 585
R655 B.n816 B.n48 585
R656 B.n734 B.n47 585
R657 B.n817 B.n47 585
R658 B.n733 B.n732 585
R659 B.n732 B.n43 585
R660 B.n731 B.n42 585
R661 B.n823 B.n42 585
R662 B.n730 B.n41 585
R663 B.n824 B.n41 585
R664 B.n729 B.n40 585
R665 B.n825 B.n40 585
R666 B.n728 B.n727 585
R667 B.n727 B.n36 585
R668 B.n726 B.n35 585
R669 B.n831 B.n35 585
R670 B.n725 B.n34 585
R671 B.n832 B.n34 585
R672 B.n724 B.n33 585
R673 B.n833 B.n33 585
R674 B.n723 B.n722 585
R675 B.n722 B.n29 585
R676 B.n721 B.n28 585
R677 B.n839 B.n28 585
R678 B.n720 B.n27 585
R679 B.n840 B.n27 585
R680 B.n719 B.n26 585
R681 B.n841 B.n26 585
R682 B.n718 B.n717 585
R683 B.n717 B.n22 585
R684 B.n716 B.n21 585
R685 B.n847 B.n21 585
R686 B.n715 B.n20 585
R687 B.n848 B.n20 585
R688 B.n714 B.n19 585
R689 B.n849 B.n19 585
R690 B.n713 B.n712 585
R691 B.n712 B.n18 585
R692 B.n711 B.n14 585
R693 B.n855 B.n14 585
R694 B.n710 B.n13 585
R695 B.n856 B.n13 585
R696 B.n709 B.n12 585
R697 B.n857 B.n12 585
R698 B.n708 B.n707 585
R699 B.n707 B.n8 585
R700 B.n706 B.n7 585
R701 B.n863 B.n7 585
R702 B.n705 B.n6 585
R703 B.n864 B.n6 585
R704 B.n704 B.n5 585
R705 B.n865 B.n5 585
R706 B.n703 B.n702 585
R707 B.n702 B.n4 585
R708 B.n701 B.n276 585
R709 B.n701 B.n700 585
R710 B.n691 B.n277 585
R711 B.n278 B.n277 585
R712 B.n693 B.n692 585
R713 B.n694 B.n693 585
R714 B.n690 B.n283 585
R715 B.n283 B.n282 585
R716 B.n689 B.n688 585
R717 B.n688 B.n687 585
R718 B.n285 B.n284 585
R719 B.n680 B.n285 585
R720 B.n679 B.n678 585
R721 B.n681 B.n679 585
R722 B.n677 B.n290 585
R723 B.n290 B.n289 585
R724 B.n676 B.n675 585
R725 B.n675 B.n674 585
R726 B.n292 B.n291 585
R727 B.n293 B.n292 585
R728 B.n667 B.n666 585
R729 B.n668 B.n667 585
R730 B.n665 B.n298 585
R731 B.n298 B.n297 585
R732 B.n664 B.n663 585
R733 B.n663 B.n662 585
R734 B.n300 B.n299 585
R735 B.n301 B.n300 585
R736 B.n655 B.n654 585
R737 B.n656 B.n655 585
R738 B.n653 B.n305 585
R739 B.n309 B.n305 585
R740 B.n652 B.n651 585
R741 B.n651 B.n650 585
R742 B.n307 B.n306 585
R743 B.n308 B.n307 585
R744 B.n643 B.n642 585
R745 B.n644 B.n643 585
R746 B.n641 B.n314 585
R747 B.n314 B.n313 585
R748 B.n640 B.n639 585
R749 B.n639 B.n638 585
R750 B.n316 B.n315 585
R751 B.n317 B.n316 585
R752 B.n631 B.n630 585
R753 B.n632 B.n631 585
R754 B.n629 B.n322 585
R755 B.n322 B.n321 585
R756 B.n628 B.n627 585
R757 B.n627 B.n626 585
R758 B.n324 B.n323 585
R759 B.n619 B.n324 585
R760 B.n618 B.n617 585
R761 B.n620 B.n618 585
R762 B.n616 B.n329 585
R763 B.n329 B.n328 585
R764 B.n615 B.n614 585
R765 B.n614 B.n613 585
R766 B.n331 B.n330 585
R767 B.n332 B.n331 585
R768 B.n606 B.n605 585
R769 B.n607 B.n606 585
R770 B.n604 B.n337 585
R771 B.n337 B.n336 585
R772 B.n603 B.n602 585
R773 B.n602 B.n601 585
R774 B.n339 B.n338 585
R775 B.n340 B.n339 585
R776 B.n594 B.n593 585
R777 B.n595 B.n594 585
R778 B.n592 B.n345 585
R779 B.n345 B.n344 585
R780 B.n591 B.n590 585
R781 B.n590 B.n589 585
R782 B.n347 B.n346 585
R783 B.n348 B.n347 585
R784 B.n582 B.n581 585
R785 B.n583 B.n582 585
R786 B.n580 B.n353 585
R787 B.n353 B.n352 585
R788 B.n579 B.n578 585
R789 B.n578 B.n577 585
R790 B.n355 B.n354 585
R791 B.n356 B.n355 585
R792 B.n570 B.n569 585
R793 B.n571 B.n570 585
R794 B.n568 B.n361 585
R795 B.n361 B.n360 585
R796 B.n567 B.n566 585
R797 B.n566 B.n565 585
R798 B.n363 B.n362 585
R799 B.n364 B.n363 585
R800 B.n558 B.n557 585
R801 B.n559 B.n558 585
R802 B.n367 B.n366 585
R803 B.n410 B.n408 585
R804 B.n411 B.n407 585
R805 B.n411 B.n368 585
R806 B.n414 B.n413 585
R807 B.n415 B.n406 585
R808 B.n417 B.n416 585
R809 B.n419 B.n405 585
R810 B.n422 B.n421 585
R811 B.n423 B.n404 585
R812 B.n425 B.n424 585
R813 B.n427 B.n403 585
R814 B.n430 B.n429 585
R815 B.n431 B.n402 585
R816 B.n433 B.n432 585
R817 B.n435 B.n401 585
R818 B.n438 B.n437 585
R819 B.n439 B.n400 585
R820 B.n441 B.n440 585
R821 B.n443 B.n399 585
R822 B.n446 B.n445 585
R823 B.n447 B.n398 585
R824 B.n449 B.n448 585
R825 B.n451 B.n397 585
R826 B.n454 B.n453 585
R827 B.n455 B.n396 585
R828 B.n457 B.n456 585
R829 B.n459 B.n395 585
R830 B.n462 B.n461 585
R831 B.n463 B.n394 585
R832 B.n465 B.n464 585
R833 B.n467 B.n393 585
R834 B.n470 B.n469 585
R835 B.n472 B.n390 585
R836 B.n474 B.n473 585
R837 B.n476 B.n389 585
R838 B.n479 B.n478 585
R839 B.n480 B.n388 585
R840 B.n482 B.n481 585
R841 B.n484 B.n387 585
R842 B.n487 B.n486 585
R843 B.n488 B.n386 585
R844 B.n493 B.n492 585
R845 B.n495 B.n385 585
R846 B.n498 B.n497 585
R847 B.n499 B.n384 585
R848 B.n501 B.n500 585
R849 B.n503 B.n383 585
R850 B.n506 B.n505 585
R851 B.n507 B.n382 585
R852 B.n509 B.n508 585
R853 B.n511 B.n381 585
R854 B.n514 B.n513 585
R855 B.n515 B.n380 585
R856 B.n517 B.n516 585
R857 B.n519 B.n379 585
R858 B.n522 B.n521 585
R859 B.n523 B.n378 585
R860 B.n525 B.n524 585
R861 B.n527 B.n377 585
R862 B.n530 B.n529 585
R863 B.n531 B.n376 585
R864 B.n533 B.n532 585
R865 B.n535 B.n375 585
R866 B.n538 B.n537 585
R867 B.n539 B.n374 585
R868 B.n541 B.n540 585
R869 B.n543 B.n373 585
R870 B.n546 B.n545 585
R871 B.n547 B.n372 585
R872 B.n549 B.n548 585
R873 B.n551 B.n371 585
R874 B.n552 B.n370 585
R875 B.n555 B.n554 585
R876 B.n556 B.n369 585
R877 B.n369 B.n368 585
R878 B.n561 B.n560 585
R879 B.n560 B.n559 585
R880 B.n562 B.n365 585
R881 B.n365 B.n364 585
R882 B.n564 B.n563 585
R883 B.n565 B.n564 585
R884 B.n359 B.n358 585
R885 B.n360 B.n359 585
R886 B.n573 B.n572 585
R887 B.n572 B.n571 585
R888 B.n574 B.n357 585
R889 B.n357 B.n356 585
R890 B.n576 B.n575 585
R891 B.n577 B.n576 585
R892 B.n351 B.n350 585
R893 B.n352 B.n351 585
R894 B.n585 B.n584 585
R895 B.n584 B.n583 585
R896 B.n586 B.n349 585
R897 B.n349 B.n348 585
R898 B.n588 B.n587 585
R899 B.n589 B.n588 585
R900 B.n343 B.n342 585
R901 B.n344 B.n343 585
R902 B.n597 B.n596 585
R903 B.n596 B.n595 585
R904 B.n598 B.n341 585
R905 B.n341 B.n340 585
R906 B.n600 B.n599 585
R907 B.n601 B.n600 585
R908 B.n335 B.n334 585
R909 B.n336 B.n335 585
R910 B.n609 B.n608 585
R911 B.n608 B.n607 585
R912 B.n610 B.n333 585
R913 B.n333 B.n332 585
R914 B.n612 B.n611 585
R915 B.n613 B.n612 585
R916 B.n327 B.n326 585
R917 B.n328 B.n327 585
R918 B.n622 B.n621 585
R919 B.n621 B.n620 585
R920 B.n623 B.n325 585
R921 B.n619 B.n325 585
R922 B.n625 B.n624 585
R923 B.n626 B.n625 585
R924 B.n320 B.n319 585
R925 B.n321 B.n320 585
R926 B.n634 B.n633 585
R927 B.n633 B.n632 585
R928 B.n635 B.n318 585
R929 B.n318 B.n317 585
R930 B.n637 B.n636 585
R931 B.n638 B.n637 585
R932 B.n312 B.n311 585
R933 B.n313 B.n312 585
R934 B.n646 B.n645 585
R935 B.n645 B.n644 585
R936 B.n647 B.n310 585
R937 B.n310 B.n308 585
R938 B.n649 B.n648 585
R939 B.n650 B.n649 585
R940 B.n304 B.n303 585
R941 B.n309 B.n304 585
R942 B.n658 B.n657 585
R943 B.n657 B.n656 585
R944 B.n659 B.n302 585
R945 B.n302 B.n301 585
R946 B.n661 B.n660 585
R947 B.n662 B.n661 585
R948 B.n296 B.n295 585
R949 B.n297 B.n296 585
R950 B.n670 B.n669 585
R951 B.n669 B.n668 585
R952 B.n671 B.n294 585
R953 B.n294 B.n293 585
R954 B.n673 B.n672 585
R955 B.n674 B.n673 585
R956 B.n288 B.n287 585
R957 B.n289 B.n288 585
R958 B.n683 B.n682 585
R959 B.n682 B.n681 585
R960 B.n684 B.n286 585
R961 B.n680 B.n286 585
R962 B.n686 B.n685 585
R963 B.n687 B.n686 585
R964 B.n281 B.n280 585
R965 B.n282 B.n281 585
R966 B.n696 B.n695 585
R967 B.n695 B.n694 585
R968 B.n697 B.n279 585
R969 B.n279 B.n278 585
R970 B.n699 B.n698 585
R971 B.n700 B.n699 585
R972 B.n2 B.n0 585
R973 B.n4 B.n2 585
R974 B.n3 B.n1 585
R975 B.n864 B.n3 585
R976 B.n862 B.n861 585
R977 B.n863 B.n862 585
R978 B.n860 B.n9 585
R979 B.n9 B.n8 585
R980 B.n859 B.n858 585
R981 B.n858 B.n857 585
R982 B.n11 B.n10 585
R983 B.n856 B.n11 585
R984 B.n854 B.n853 585
R985 B.n855 B.n854 585
R986 B.n852 B.n15 585
R987 B.n18 B.n15 585
R988 B.n851 B.n850 585
R989 B.n850 B.n849 585
R990 B.n17 B.n16 585
R991 B.n848 B.n17 585
R992 B.n846 B.n845 585
R993 B.n847 B.n846 585
R994 B.n844 B.n23 585
R995 B.n23 B.n22 585
R996 B.n843 B.n842 585
R997 B.n842 B.n841 585
R998 B.n25 B.n24 585
R999 B.n840 B.n25 585
R1000 B.n838 B.n837 585
R1001 B.n839 B.n838 585
R1002 B.n836 B.n30 585
R1003 B.n30 B.n29 585
R1004 B.n835 B.n834 585
R1005 B.n834 B.n833 585
R1006 B.n32 B.n31 585
R1007 B.n832 B.n32 585
R1008 B.n830 B.n829 585
R1009 B.n831 B.n830 585
R1010 B.n828 B.n37 585
R1011 B.n37 B.n36 585
R1012 B.n827 B.n826 585
R1013 B.n826 B.n825 585
R1014 B.n39 B.n38 585
R1015 B.n824 B.n39 585
R1016 B.n822 B.n821 585
R1017 B.n823 B.n822 585
R1018 B.n820 B.n44 585
R1019 B.n44 B.n43 585
R1020 B.n819 B.n818 585
R1021 B.n818 B.n817 585
R1022 B.n46 B.n45 585
R1023 B.n816 B.n46 585
R1024 B.n814 B.n813 585
R1025 B.n815 B.n814 585
R1026 B.n812 B.n50 585
R1027 B.n53 B.n50 585
R1028 B.n811 B.n810 585
R1029 B.n810 B.n809 585
R1030 B.n52 B.n51 585
R1031 B.n808 B.n52 585
R1032 B.n806 B.n805 585
R1033 B.n807 B.n806 585
R1034 B.n804 B.n58 585
R1035 B.n58 B.n57 585
R1036 B.n803 B.n802 585
R1037 B.n802 B.n801 585
R1038 B.n60 B.n59 585
R1039 B.n800 B.n60 585
R1040 B.n798 B.n797 585
R1041 B.n799 B.n798 585
R1042 B.n796 B.n65 585
R1043 B.n65 B.n64 585
R1044 B.n795 B.n794 585
R1045 B.n794 B.n793 585
R1046 B.n67 B.n66 585
R1047 B.n792 B.n67 585
R1048 B.n790 B.n789 585
R1049 B.n791 B.n790 585
R1050 B.n788 B.n72 585
R1051 B.n72 B.n71 585
R1052 B.n787 B.n786 585
R1053 B.n786 B.n785 585
R1054 B.n74 B.n73 585
R1055 B.n784 B.n74 585
R1056 B.n782 B.n781 585
R1057 B.n783 B.n782 585
R1058 B.n780 B.n79 585
R1059 B.n79 B.n78 585
R1060 B.n779 B.n778 585
R1061 B.n778 B.n777 585
R1062 B.n81 B.n80 585
R1063 B.n776 B.n81 585
R1064 B.n774 B.n773 585
R1065 B.n775 B.n774 585
R1066 B.n772 B.n86 585
R1067 B.n86 B.n85 585
R1068 B.n771 B.n770 585
R1069 B.n770 B.n769 585
R1070 B.n867 B.n866 585
R1071 B.n866 B.n865 585
R1072 B.n560 B.n367 545.355
R1073 B.n770 B.n88 545.355
R1074 B.n558 B.n369 545.355
R1075 B.n766 B.n89 545.355
R1076 B.n489 B.t9 293.849
R1077 B.n127 B.t15 293.849
R1078 B.n391 B.t19 293.849
R1079 B.n130 B.t12 293.849
R1080 B.n489 B.t6 277.685
R1081 B.n391 B.t17 277.685
R1082 B.n130 B.t10 277.685
R1083 B.n127 B.t14 277.685
R1084 B.n768 B.n767 256.663
R1085 B.n768 B.n125 256.663
R1086 B.n768 B.n124 256.663
R1087 B.n768 B.n123 256.663
R1088 B.n768 B.n122 256.663
R1089 B.n768 B.n121 256.663
R1090 B.n768 B.n120 256.663
R1091 B.n768 B.n119 256.663
R1092 B.n768 B.n118 256.663
R1093 B.n768 B.n117 256.663
R1094 B.n768 B.n116 256.663
R1095 B.n768 B.n115 256.663
R1096 B.n768 B.n114 256.663
R1097 B.n768 B.n113 256.663
R1098 B.n768 B.n112 256.663
R1099 B.n768 B.n111 256.663
R1100 B.n768 B.n110 256.663
R1101 B.n768 B.n109 256.663
R1102 B.n768 B.n108 256.663
R1103 B.n768 B.n107 256.663
R1104 B.n768 B.n106 256.663
R1105 B.n768 B.n105 256.663
R1106 B.n768 B.n104 256.663
R1107 B.n768 B.n103 256.663
R1108 B.n768 B.n102 256.663
R1109 B.n768 B.n101 256.663
R1110 B.n768 B.n100 256.663
R1111 B.n768 B.n99 256.663
R1112 B.n768 B.n98 256.663
R1113 B.n768 B.n97 256.663
R1114 B.n768 B.n96 256.663
R1115 B.n768 B.n95 256.663
R1116 B.n768 B.n94 256.663
R1117 B.n768 B.n93 256.663
R1118 B.n768 B.n92 256.663
R1119 B.n768 B.n91 256.663
R1120 B.n768 B.n90 256.663
R1121 B.n409 B.n368 256.663
R1122 B.n412 B.n368 256.663
R1123 B.n418 B.n368 256.663
R1124 B.n420 B.n368 256.663
R1125 B.n426 B.n368 256.663
R1126 B.n428 B.n368 256.663
R1127 B.n434 B.n368 256.663
R1128 B.n436 B.n368 256.663
R1129 B.n442 B.n368 256.663
R1130 B.n444 B.n368 256.663
R1131 B.n450 B.n368 256.663
R1132 B.n452 B.n368 256.663
R1133 B.n458 B.n368 256.663
R1134 B.n460 B.n368 256.663
R1135 B.n466 B.n368 256.663
R1136 B.n468 B.n368 256.663
R1137 B.n475 B.n368 256.663
R1138 B.n477 B.n368 256.663
R1139 B.n483 B.n368 256.663
R1140 B.n485 B.n368 256.663
R1141 B.n494 B.n368 256.663
R1142 B.n496 B.n368 256.663
R1143 B.n502 B.n368 256.663
R1144 B.n504 B.n368 256.663
R1145 B.n510 B.n368 256.663
R1146 B.n512 B.n368 256.663
R1147 B.n518 B.n368 256.663
R1148 B.n520 B.n368 256.663
R1149 B.n526 B.n368 256.663
R1150 B.n528 B.n368 256.663
R1151 B.n534 B.n368 256.663
R1152 B.n536 B.n368 256.663
R1153 B.n542 B.n368 256.663
R1154 B.n544 B.n368 256.663
R1155 B.n550 B.n368 256.663
R1156 B.n553 B.n368 256.663
R1157 B.n490 B.t8 227.715
R1158 B.n128 B.t16 227.715
R1159 B.n392 B.t18 227.715
R1160 B.n131 B.t13 227.715
R1161 B.n560 B.n365 163.367
R1162 B.n564 B.n365 163.367
R1163 B.n564 B.n359 163.367
R1164 B.n572 B.n359 163.367
R1165 B.n572 B.n357 163.367
R1166 B.n576 B.n357 163.367
R1167 B.n576 B.n351 163.367
R1168 B.n584 B.n351 163.367
R1169 B.n584 B.n349 163.367
R1170 B.n588 B.n349 163.367
R1171 B.n588 B.n343 163.367
R1172 B.n596 B.n343 163.367
R1173 B.n596 B.n341 163.367
R1174 B.n600 B.n341 163.367
R1175 B.n600 B.n335 163.367
R1176 B.n608 B.n335 163.367
R1177 B.n608 B.n333 163.367
R1178 B.n612 B.n333 163.367
R1179 B.n612 B.n327 163.367
R1180 B.n621 B.n327 163.367
R1181 B.n621 B.n325 163.367
R1182 B.n625 B.n325 163.367
R1183 B.n625 B.n320 163.367
R1184 B.n633 B.n320 163.367
R1185 B.n633 B.n318 163.367
R1186 B.n637 B.n318 163.367
R1187 B.n637 B.n312 163.367
R1188 B.n645 B.n312 163.367
R1189 B.n645 B.n310 163.367
R1190 B.n649 B.n310 163.367
R1191 B.n649 B.n304 163.367
R1192 B.n657 B.n304 163.367
R1193 B.n657 B.n302 163.367
R1194 B.n661 B.n302 163.367
R1195 B.n661 B.n296 163.367
R1196 B.n669 B.n296 163.367
R1197 B.n669 B.n294 163.367
R1198 B.n673 B.n294 163.367
R1199 B.n673 B.n288 163.367
R1200 B.n682 B.n288 163.367
R1201 B.n682 B.n286 163.367
R1202 B.n686 B.n286 163.367
R1203 B.n686 B.n281 163.367
R1204 B.n695 B.n281 163.367
R1205 B.n695 B.n279 163.367
R1206 B.n699 B.n279 163.367
R1207 B.n699 B.n2 163.367
R1208 B.n866 B.n2 163.367
R1209 B.n866 B.n3 163.367
R1210 B.n862 B.n3 163.367
R1211 B.n862 B.n9 163.367
R1212 B.n858 B.n9 163.367
R1213 B.n858 B.n11 163.367
R1214 B.n854 B.n11 163.367
R1215 B.n854 B.n15 163.367
R1216 B.n850 B.n15 163.367
R1217 B.n850 B.n17 163.367
R1218 B.n846 B.n17 163.367
R1219 B.n846 B.n23 163.367
R1220 B.n842 B.n23 163.367
R1221 B.n842 B.n25 163.367
R1222 B.n838 B.n25 163.367
R1223 B.n838 B.n30 163.367
R1224 B.n834 B.n30 163.367
R1225 B.n834 B.n32 163.367
R1226 B.n830 B.n32 163.367
R1227 B.n830 B.n37 163.367
R1228 B.n826 B.n37 163.367
R1229 B.n826 B.n39 163.367
R1230 B.n822 B.n39 163.367
R1231 B.n822 B.n44 163.367
R1232 B.n818 B.n44 163.367
R1233 B.n818 B.n46 163.367
R1234 B.n814 B.n46 163.367
R1235 B.n814 B.n50 163.367
R1236 B.n810 B.n50 163.367
R1237 B.n810 B.n52 163.367
R1238 B.n806 B.n52 163.367
R1239 B.n806 B.n58 163.367
R1240 B.n802 B.n58 163.367
R1241 B.n802 B.n60 163.367
R1242 B.n798 B.n60 163.367
R1243 B.n798 B.n65 163.367
R1244 B.n794 B.n65 163.367
R1245 B.n794 B.n67 163.367
R1246 B.n790 B.n67 163.367
R1247 B.n790 B.n72 163.367
R1248 B.n786 B.n72 163.367
R1249 B.n786 B.n74 163.367
R1250 B.n782 B.n74 163.367
R1251 B.n782 B.n79 163.367
R1252 B.n778 B.n79 163.367
R1253 B.n778 B.n81 163.367
R1254 B.n774 B.n81 163.367
R1255 B.n774 B.n86 163.367
R1256 B.n770 B.n86 163.367
R1257 B.n411 B.n410 163.367
R1258 B.n413 B.n411 163.367
R1259 B.n417 B.n406 163.367
R1260 B.n421 B.n419 163.367
R1261 B.n425 B.n404 163.367
R1262 B.n429 B.n427 163.367
R1263 B.n433 B.n402 163.367
R1264 B.n437 B.n435 163.367
R1265 B.n441 B.n400 163.367
R1266 B.n445 B.n443 163.367
R1267 B.n449 B.n398 163.367
R1268 B.n453 B.n451 163.367
R1269 B.n457 B.n396 163.367
R1270 B.n461 B.n459 163.367
R1271 B.n465 B.n394 163.367
R1272 B.n469 B.n467 163.367
R1273 B.n474 B.n390 163.367
R1274 B.n478 B.n476 163.367
R1275 B.n482 B.n388 163.367
R1276 B.n486 B.n484 163.367
R1277 B.n493 B.n386 163.367
R1278 B.n497 B.n495 163.367
R1279 B.n501 B.n384 163.367
R1280 B.n505 B.n503 163.367
R1281 B.n509 B.n382 163.367
R1282 B.n513 B.n511 163.367
R1283 B.n517 B.n380 163.367
R1284 B.n521 B.n519 163.367
R1285 B.n525 B.n378 163.367
R1286 B.n529 B.n527 163.367
R1287 B.n533 B.n376 163.367
R1288 B.n537 B.n535 163.367
R1289 B.n541 B.n374 163.367
R1290 B.n545 B.n543 163.367
R1291 B.n549 B.n372 163.367
R1292 B.n552 B.n551 163.367
R1293 B.n554 B.n369 163.367
R1294 B.n558 B.n363 163.367
R1295 B.n566 B.n363 163.367
R1296 B.n566 B.n361 163.367
R1297 B.n570 B.n361 163.367
R1298 B.n570 B.n355 163.367
R1299 B.n578 B.n355 163.367
R1300 B.n578 B.n353 163.367
R1301 B.n582 B.n353 163.367
R1302 B.n582 B.n347 163.367
R1303 B.n590 B.n347 163.367
R1304 B.n590 B.n345 163.367
R1305 B.n594 B.n345 163.367
R1306 B.n594 B.n339 163.367
R1307 B.n602 B.n339 163.367
R1308 B.n602 B.n337 163.367
R1309 B.n606 B.n337 163.367
R1310 B.n606 B.n331 163.367
R1311 B.n614 B.n331 163.367
R1312 B.n614 B.n329 163.367
R1313 B.n618 B.n329 163.367
R1314 B.n618 B.n324 163.367
R1315 B.n627 B.n324 163.367
R1316 B.n627 B.n322 163.367
R1317 B.n631 B.n322 163.367
R1318 B.n631 B.n316 163.367
R1319 B.n639 B.n316 163.367
R1320 B.n639 B.n314 163.367
R1321 B.n643 B.n314 163.367
R1322 B.n643 B.n307 163.367
R1323 B.n651 B.n307 163.367
R1324 B.n651 B.n305 163.367
R1325 B.n655 B.n305 163.367
R1326 B.n655 B.n300 163.367
R1327 B.n663 B.n300 163.367
R1328 B.n663 B.n298 163.367
R1329 B.n667 B.n298 163.367
R1330 B.n667 B.n292 163.367
R1331 B.n675 B.n292 163.367
R1332 B.n675 B.n290 163.367
R1333 B.n679 B.n290 163.367
R1334 B.n679 B.n285 163.367
R1335 B.n688 B.n285 163.367
R1336 B.n688 B.n283 163.367
R1337 B.n693 B.n283 163.367
R1338 B.n693 B.n277 163.367
R1339 B.n701 B.n277 163.367
R1340 B.n702 B.n701 163.367
R1341 B.n702 B.n5 163.367
R1342 B.n6 B.n5 163.367
R1343 B.n7 B.n6 163.367
R1344 B.n707 B.n7 163.367
R1345 B.n707 B.n12 163.367
R1346 B.n13 B.n12 163.367
R1347 B.n14 B.n13 163.367
R1348 B.n712 B.n14 163.367
R1349 B.n712 B.n19 163.367
R1350 B.n20 B.n19 163.367
R1351 B.n21 B.n20 163.367
R1352 B.n717 B.n21 163.367
R1353 B.n717 B.n26 163.367
R1354 B.n27 B.n26 163.367
R1355 B.n28 B.n27 163.367
R1356 B.n722 B.n28 163.367
R1357 B.n722 B.n33 163.367
R1358 B.n34 B.n33 163.367
R1359 B.n35 B.n34 163.367
R1360 B.n727 B.n35 163.367
R1361 B.n727 B.n40 163.367
R1362 B.n41 B.n40 163.367
R1363 B.n42 B.n41 163.367
R1364 B.n732 B.n42 163.367
R1365 B.n732 B.n47 163.367
R1366 B.n48 B.n47 163.367
R1367 B.n49 B.n48 163.367
R1368 B.n737 B.n49 163.367
R1369 B.n737 B.n54 163.367
R1370 B.n55 B.n54 163.367
R1371 B.n56 B.n55 163.367
R1372 B.n742 B.n56 163.367
R1373 B.n742 B.n61 163.367
R1374 B.n62 B.n61 163.367
R1375 B.n63 B.n62 163.367
R1376 B.n747 B.n63 163.367
R1377 B.n747 B.n68 163.367
R1378 B.n69 B.n68 163.367
R1379 B.n70 B.n69 163.367
R1380 B.n752 B.n70 163.367
R1381 B.n752 B.n75 163.367
R1382 B.n76 B.n75 163.367
R1383 B.n77 B.n76 163.367
R1384 B.n757 B.n77 163.367
R1385 B.n757 B.n82 163.367
R1386 B.n83 B.n82 163.367
R1387 B.n84 B.n83 163.367
R1388 B.n762 B.n84 163.367
R1389 B.n762 B.n89 163.367
R1390 B.n135 B.n134 163.367
R1391 B.n139 B.n138 163.367
R1392 B.n143 B.n142 163.367
R1393 B.n147 B.n146 163.367
R1394 B.n151 B.n150 163.367
R1395 B.n155 B.n154 163.367
R1396 B.n159 B.n158 163.367
R1397 B.n163 B.n162 163.367
R1398 B.n167 B.n166 163.367
R1399 B.n171 B.n170 163.367
R1400 B.n175 B.n174 163.367
R1401 B.n179 B.n178 163.367
R1402 B.n183 B.n182 163.367
R1403 B.n187 B.n186 163.367
R1404 B.n191 B.n190 163.367
R1405 B.n195 B.n194 163.367
R1406 B.n199 B.n198 163.367
R1407 B.n203 B.n202 163.367
R1408 B.n207 B.n206 163.367
R1409 B.n211 B.n210 163.367
R1410 B.n215 B.n214 163.367
R1411 B.n219 B.n218 163.367
R1412 B.n223 B.n222 163.367
R1413 B.n227 B.n226 163.367
R1414 B.n231 B.n230 163.367
R1415 B.n235 B.n234 163.367
R1416 B.n239 B.n238 163.367
R1417 B.n243 B.n242 163.367
R1418 B.n247 B.n246 163.367
R1419 B.n251 B.n250 163.367
R1420 B.n255 B.n254 163.367
R1421 B.n259 B.n258 163.367
R1422 B.n263 B.n262 163.367
R1423 B.n267 B.n266 163.367
R1424 B.n271 B.n270 163.367
R1425 B.n273 B.n126 163.367
R1426 B.n559 B.n368 108.478
R1427 B.n769 B.n768 108.478
R1428 B.n409 B.n367 71.676
R1429 B.n413 B.n412 71.676
R1430 B.n418 B.n417 71.676
R1431 B.n421 B.n420 71.676
R1432 B.n426 B.n425 71.676
R1433 B.n429 B.n428 71.676
R1434 B.n434 B.n433 71.676
R1435 B.n437 B.n436 71.676
R1436 B.n442 B.n441 71.676
R1437 B.n445 B.n444 71.676
R1438 B.n450 B.n449 71.676
R1439 B.n453 B.n452 71.676
R1440 B.n458 B.n457 71.676
R1441 B.n461 B.n460 71.676
R1442 B.n466 B.n465 71.676
R1443 B.n469 B.n468 71.676
R1444 B.n475 B.n474 71.676
R1445 B.n478 B.n477 71.676
R1446 B.n483 B.n482 71.676
R1447 B.n486 B.n485 71.676
R1448 B.n494 B.n493 71.676
R1449 B.n497 B.n496 71.676
R1450 B.n502 B.n501 71.676
R1451 B.n505 B.n504 71.676
R1452 B.n510 B.n509 71.676
R1453 B.n513 B.n512 71.676
R1454 B.n518 B.n517 71.676
R1455 B.n521 B.n520 71.676
R1456 B.n526 B.n525 71.676
R1457 B.n529 B.n528 71.676
R1458 B.n534 B.n533 71.676
R1459 B.n537 B.n536 71.676
R1460 B.n542 B.n541 71.676
R1461 B.n545 B.n544 71.676
R1462 B.n550 B.n549 71.676
R1463 B.n553 B.n552 71.676
R1464 B.n90 B.n88 71.676
R1465 B.n135 B.n91 71.676
R1466 B.n139 B.n92 71.676
R1467 B.n143 B.n93 71.676
R1468 B.n147 B.n94 71.676
R1469 B.n151 B.n95 71.676
R1470 B.n155 B.n96 71.676
R1471 B.n159 B.n97 71.676
R1472 B.n163 B.n98 71.676
R1473 B.n167 B.n99 71.676
R1474 B.n171 B.n100 71.676
R1475 B.n175 B.n101 71.676
R1476 B.n179 B.n102 71.676
R1477 B.n183 B.n103 71.676
R1478 B.n187 B.n104 71.676
R1479 B.n191 B.n105 71.676
R1480 B.n195 B.n106 71.676
R1481 B.n199 B.n107 71.676
R1482 B.n203 B.n108 71.676
R1483 B.n207 B.n109 71.676
R1484 B.n211 B.n110 71.676
R1485 B.n215 B.n111 71.676
R1486 B.n219 B.n112 71.676
R1487 B.n223 B.n113 71.676
R1488 B.n227 B.n114 71.676
R1489 B.n231 B.n115 71.676
R1490 B.n235 B.n116 71.676
R1491 B.n239 B.n117 71.676
R1492 B.n243 B.n118 71.676
R1493 B.n247 B.n119 71.676
R1494 B.n251 B.n120 71.676
R1495 B.n255 B.n121 71.676
R1496 B.n259 B.n122 71.676
R1497 B.n263 B.n123 71.676
R1498 B.n267 B.n124 71.676
R1499 B.n271 B.n125 71.676
R1500 B.n767 B.n126 71.676
R1501 B.n767 B.n766 71.676
R1502 B.n273 B.n125 71.676
R1503 B.n270 B.n124 71.676
R1504 B.n266 B.n123 71.676
R1505 B.n262 B.n122 71.676
R1506 B.n258 B.n121 71.676
R1507 B.n254 B.n120 71.676
R1508 B.n250 B.n119 71.676
R1509 B.n246 B.n118 71.676
R1510 B.n242 B.n117 71.676
R1511 B.n238 B.n116 71.676
R1512 B.n234 B.n115 71.676
R1513 B.n230 B.n114 71.676
R1514 B.n226 B.n113 71.676
R1515 B.n222 B.n112 71.676
R1516 B.n218 B.n111 71.676
R1517 B.n214 B.n110 71.676
R1518 B.n210 B.n109 71.676
R1519 B.n206 B.n108 71.676
R1520 B.n202 B.n107 71.676
R1521 B.n198 B.n106 71.676
R1522 B.n194 B.n105 71.676
R1523 B.n190 B.n104 71.676
R1524 B.n186 B.n103 71.676
R1525 B.n182 B.n102 71.676
R1526 B.n178 B.n101 71.676
R1527 B.n174 B.n100 71.676
R1528 B.n170 B.n99 71.676
R1529 B.n166 B.n98 71.676
R1530 B.n162 B.n97 71.676
R1531 B.n158 B.n96 71.676
R1532 B.n154 B.n95 71.676
R1533 B.n150 B.n94 71.676
R1534 B.n146 B.n93 71.676
R1535 B.n142 B.n92 71.676
R1536 B.n138 B.n91 71.676
R1537 B.n134 B.n90 71.676
R1538 B.n410 B.n409 71.676
R1539 B.n412 B.n406 71.676
R1540 B.n419 B.n418 71.676
R1541 B.n420 B.n404 71.676
R1542 B.n427 B.n426 71.676
R1543 B.n428 B.n402 71.676
R1544 B.n435 B.n434 71.676
R1545 B.n436 B.n400 71.676
R1546 B.n443 B.n442 71.676
R1547 B.n444 B.n398 71.676
R1548 B.n451 B.n450 71.676
R1549 B.n452 B.n396 71.676
R1550 B.n459 B.n458 71.676
R1551 B.n460 B.n394 71.676
R1552 B.n467 B.n466 71.676
R1553 B.n468 B.n390 71.676
R1554 B.n476 B.n475 71.676
R1555 B.n477 B.n388 71.676
R1556 B.n484 B.n483 71.676
R1557 B.n485 B.n386 71.676
R1558 B.n495 B.n494 71.676
R1559 B.n496 B.n384 71.676
R1560 B.n503 B.n502 71.676
R1561 B.n504 B.n382 71.676
R1562 B.n511 B.n510 71.676
R1563 B.n512 B.n380 71.676
R1564 B.n519 B.n518 71.676
R1565 B.n520 B.n378 71.676
R1566 B.n527 B.n526 71.676
R1567 B.n528 B.n376 71.676
R1568 B.n535 B.n534 71.676
R1569 B.n536 B.n374 71.676
R1570 B.n543 B.n542 71.676
R1571 B.n544 B.n372 71.676
R1572 B.n551 B.n550 71.676
R1573 B.n554 B.n553 71.676
R1574 B.n490 B.n489 66.1338
R1575 B.n392 B.n391 66.1338
R1576 B.n131 B.n130 66.1338
R1577 B.n128 B.n127 66.1338
R1578 B.n491 B.n490 59.5399
R1579 B.n471 B.n392 59.5399
R1580 B.n132 B.n131 59.5399
R1581 B.n129 B.n128 59.5399
R1582 B.n559 B.n364 53.069
R1583 B.n565 B.n364 53.069
R1584 B.n565 B.n360 53.069
R1585 B.n571 B.n360 53.069
R1586 B.n571 B.n356 53.069
R1587 B.n577 B.n356 53.069
R1588 B.n577 B.n352 53.069
R1589 B.n583 B.n352 53.069
R1590 B.n589 B.n348 53.069
R1591 B.n589 B.n344 53.069
R1592 B.n595 B.n344 53.069
R1593 B.n595 B.n340 53.069
R1594 B.n601 B.n340 53.069
R1595 B.n601 B.n336 53.069
R1596 B.n607 B.n336 53.069
R1597 B.n607 B.n332 53.069
R1598 B.n613 B.n332 53.069
R1599 B.n613 B.n328 53.069
R1600 B.n620 B.n328 53.069
R1601 B.n620 B.n619 53.069
R1602 B.n626 B.n321 53.069
R1603 B.n632 B.n321 53.069
R1604 B.n632 B.n317 53.069
R1605 B.n638 B.n317 53.069
R1606 B.n638 B.n313 53.069
R1607 B.n644 B.n313 53.069
R1608 B.n644 B.n308 53.069
R1609 B.n650 B.n308 53.069
R1610 B.n650 B.n309 53.069
R1611 B.n656 B.n301 53.069
R1612 B.n662 B.n301 53.069
R1613 B.n662 B.n297 53.069
R1614 B.n668 B.n297 53.069
R1615 B.n668 B.n293 53.069
R1616 B.n674 B.n293 53.069
R1617 B.n674 B.n289 53.069
R1618 B.n681 B.n289 53.069
R1619 B.n681 B.n680 53.069
R1620 B.n687 B.n282 53.069
R1621 B.n694 B.n282 53.069
R1622 B.n694 B.n278 53.069
R1623 B.n700 B.n278 53.069
R1624 B.n700 B.n4 53.069
R1625 B.n865 B.n4 53.069
R1626 B.n865 B.n864 53.069
R1627 B.n864 B.n863 53.069
R1628 B.n863 B.n8 53.069
R1629 B.n857 B.n8 53.069
R1630 B.n857 B.n856 53.069
R1631 B.n856 B.n855 53.069
R1632 B.n849 B.n18 53.069
R1633 B.n849 B.n848 53.069
R1634 B.n848 B.n847 53.069
R1635 B.n847 B.n22 53.069
R1636 B.n841 B.n22 53.069
R1637 B.n841 B.n840 53.069
R1638 B.n840 B.n839 53.069
R1639 B.n839 B.n29 53.069
R1640 B.n833 B.n29 53.069
R1641 B.n832 B.n831 53.069
R1642 B.n831 B.n36 53.069
R1643 B.n825 B.n36 53.069
R1644 B.n825 B.n824 53.069
R1645 B.n824 B.n823 53.069
R1646 B.n823 B.n43 53.069
R1647 B.n817 B.n43 53.069
R1648 B.n817 B.n816 53.069
R1649 B.n816 B.n815 53.069
R1650 B.n809 B.n53 53.069
R1651 B.n809 B.n808 53.069
R1652 B.n808 B.n807 53.069
R1653 B.n807 B.n57 53.069
R1654 B.n801 B.n57 53.069
R1655 B.n801 B.n800 53.069
R1656 B.n800 B.n799 53.069
R1657 B.n799 B.n64 53.069
R1658 B.n793 B.n64 53.069
R1659 B.n793 B.n792 53.069
R1660 B.n792 B.n791 53.069
R1661 B.n791 B.n71 53.069
R1662 B.n785 B.n784 53.069
R1663 B.n784 B.n783 53.069
R1664 B.n783 B.n78 53.069
R1665 B.n777 B.n78 53.069
R1666 B.n777 B.n776 53.069
R1667 B.n776 B.n775 53.069
R1668 B.n775 B.n85 53.069
R1669 B.n769 B.n85 53.069
R1670 B.t7 B.n348 48.3865
R1671 B.t11 B.n71 48.3865
R1672 B.n626 B.t2 35.8998
R1673 B.n815 B.t3 35.8998
R1674 B.n765 B.n764 35.4346
R1675 B.n771 B.n87 35.4346
R1676 B.n557 B.n556 35.4346
R1677 B.n561 B.n366 35.4346
R1678 B.n656 B.t0 34.3389
R1679 B.n833 B.t5 34.3389
R1680 B.n687 B.t1 32.7781
R1681 B.n855 B.t4 32.7781
R1682 B.n680 B.t1 20.2914
R1683 B.n18 B.t4 20.2914
R1684 B.n309 B.t0 18.7305
R1685 B.t5 B.n832 18.7305
R1686 B B.n867 18.0485
R1687 B.n619 B.t2 17.1697
R1688 B.n53 B.t3 17.1697
R1689 B.n133 B.n87 10.6151
R1690 B.n136 B.n133 10.6151
R1691 B.n137 B.n136 10.6151
R1692 B.n140 B.n137 10.6151
R1693 B.n141 B.n140 10.6151
R1694 B.n144 B.n141 10.6151
R1695 B.n145 B.n144 10.6151
R1696 B.n148 B.n145 10.6151
R1697 B.n149 B.n148 10.6151
R1698 B.n152 B.n149 10.6151
R1699 B.n153 B.n152 10.6151
R1700 B.n156 B.n153 10.6151
R1701 B.n157 B.n156 10.6151
R1702 B.n160 B.n157 10.6151
R1703 B.n161 B.n160 10.6151
R1704 B.n164 B.n161 10.6151
R1705 B.n165 B.n164 10.6151
R1706 B.n168 B.n165 10.6151
R1707 B.n169 B.n168 10.6151
R1708 B.n172 B.n169 10.6151
R1709 B.n173 B.n172 10.6151
R1710 B.n176 B.n173 10.6151
R1711 B.n177 B.n176 10.6151
R1712 B.n180 B.n177 10.6151
R1713 B.n181 B.n180 10.6151
R1714 B.n184 B.n181 10.6151
R1715 B.n185 B.n184 10.6151
R1716 B.n188 B.n185 10.6151
R1717 B.n189 B.n188 10.6151
R1718 B.n192 B.n189 10.6151
R1719 B.n193 B.n192 10.6151
R1720 B.n197 B.n196 10.6151
R1721 B.n200 B.n197 10.6151
R1722 B.n201 B.n200 10.6151
R1723 B.n204 B.n201 10.6151
R1724 B.n205 B.n204 10.6151
R1725 B.n208 B.n205 10.6151
R1726 B.n209 B.n208 10.6151
R1727 B.n212 B.n209 10.6151
R1728 B.n213 B.n212 10.6151
R1729 B.n217 B.n216 10.6151
R1730 B.n220 B.n217 10.6151
R1731 B.n221 B.n220 10.6151
R1732 B.n224 B.n221 10.6151
R1733 B.n225 B.n224 10.6151
R1734 B.n228 B.n225 10.6151
R1735 B.n229 B.n228 10.6151
R1736 B.n232 B.n229 10.6151
R1737 B.n233 B.n232 10.6151
R1738 B.n236 B.n233 10.6151
R1739 B.n237 B.n236 10.6151
R1740 B.n240 B.n237 10.6151
R1741 B.n241 B.n240 10.6151
R1742 B.n244 B.n241 10.6151
R1743 B.n245 B.n244 10.6151
R1744 B.n248 B.n245 10.6151
R1745 B.n249 B.n248 10.6151
R1746 B.n252 B.n249 10.6151
R1747 B.n253 B.n252 10.6151
R1748 B.n256 B.n253 10.6151
R1749 B.n257 B.n256 10.6151
R1750 B.n260 B.n257 10.6151
R1751 B.n261 B.n260 10.6151
R1752 B.n264 B.n261 10.6151
R1753 B.n265 B.n264 10.6151
R1754 B.n268 B.n265 10.6151
R1755 B.n269 B.n268 10.6151
R1756 B.n272 B.n269 10.6151
R1757 B.n274 B.n272 10.6151
R1758 B.n275 B.n274 10.6151
R1759 B.n765 B.n275 10.6151
R1760 B.n557 B.n362 10.6151
R1761 B.n567 B.n362 10.6151
R1762 B.n568 B.n567 10.6151
R1763 B.n569 B.n568 10.6151
R1764 B.n569 B.n354 10.6151
R1765 B.n579 B.n354 10.6151
R1766 B.n580 B.n579 10.6151
R1767 B.n581 B.n580 10.6151
R1768 B.n581 B.n346 10.6151
R1769 B.n591 B.n346 10.6151
R1770 B.n592 B.n591 10.6151
R1771 B.n593 B.n592 10.6151
R1772 B.n593 B.n338 10.6151
R1773 B.n603 B.n338 10.6151
R1774 B.n604 B.n603 10.6151
R1775 B.n605 B.n604 10.6151
R1776 B.n605 B.n330 10.6151
R1777 B.n615 B.n330 10.6151
R1778 B.n616 B.n615 10.6151
R1779 B.n617 B.n616 10.6151
R1780 B.n617 B.n323 10.6151
R1781 B.n628 B.n323 10.6151
R1782 B.n629 B.n628 10.6151
R1783 B.n630 B.n629 10.6151
R1784 B.n630 B.n315 10.6151
R1785 B.n640 B.n315 10.6151
R1786 B.n641 B.n640 10.6151
R1787 B.n642 B.n641 10.6151
R1788 B.n642 B.n306 10.6151
R1789 B.n652 B.n306 10.6151
R1790 B.n653 B.n652 10.6151
R1791 B.n654 B.n653 10.6151
R1792 B.n654 B.n299 10.6151
R1793 B.n664 B.n299 10.6151
R1794 B.n665 B.n664 10.6151
R1795 B.n666 B.n665 10.6151
R1796 B.n666 B.n291 10.6151
R1797 B.n676 B.n291 10.6151
R1798 B.n677 B.n676 10.6151
R1799 B.n678 B.n677 10.6151
R1800 B.n678 B.n284 10.6151
R1801 B.n689 B.n284 10.6151
R1802 B.n690 B.n689 10.6151
R1803 B.n692 B.n690 10.6151
R1804 B.n692 B.n691 10.6151
R1805 B.n691 B.n276 10.6151
R1806 B.n703 B.n276 10.6151
R1807 B.n704 B.n703 10.6151
R1808 B.n705 B.n704 10.6151
R1809 B.n706 B.n705 10.6151
R1810 B.n708 B.n706 10.6151
R1811 B.n709 B.n708 10.6151
R1812 B.n710 B.n709 10.6151
R1813 B.n711 B.n710 10.6151
R1814 B.n713 B.n711 10.6151
R1815 B.n714 B.n713 10.6151
R1816 B.n715 B.n714 10.6151
R1817 B.n716 B.n715 10.6151
R1818 B.n718 B.n716 10.6151
R1819 B.n719 B.n718 10.6151
R1820 B.n720 B.n719 10.6151
R1821 B.n721 B.n720 10.6151
R1822 B.n723 B.n721 10.6151
R1823 B.n724 B.n723 10.6151
R1824 B.n725 B.n724 10.6151
R1825 B.n726 B.n725 10.6151
R1826 B.n728 B.n726 10.6151
R1827 B.n729 B.n728 10.6151
R1828 B.n730 B.n729 10.6151
R1829 B.n731 B.n730 10.6151
R1830 B.n733 B.n731 10.6151
R1831 B.n734 B.n733 10.6151
R1832 B.n735 B.n734 10.6151
R1833 B.n736 B.n735 10.6151
R1834 B.n738 B.n736 10.6151
R1835 B.n739 B.n738 10.6151
R1836 B.n740 B.n739 10.6151
R1837 B.n741 B.n740 10.6151
R1838 B.n743 B.n741 10.6151
R1839 B.n744 B.n743 10.6151
R1840 B.n745 B.n744 10.6151
R1841 B.n746 B.n745 10.6151
R1842 B.n748 B.n746 10.6151
R1843 B.n749 B.n748 10.6151
R1844 B.n750 B.n749 10.6151
R1845 B.n751 B.n750 10.6151
R1846 B.n753 B.n751 10.6151
R1847 B.n754 B.n753 10.6151
R1848 B.n755 B.n754 10.6151
R1849 B.n756 B.n755 10.6151
R1850 B.n758 B.n756 10.6151
R1851 B.n759 B.n758 10.6151
R1852 B.n760 B.n759 10.6151
R1853 B.n761 B.n760 10.6151
R1854 B.n763 B.n761 10.6151
R1855 B.n764 B.n763 10.6151
R1856 B.n408 B.n366 10.6151
R1857 B.n408 B.n407 10.6151
R1858 B.n414 B.n407 10.6151
R1859 B.n415 B.n414 10.6151
R1860 B.n416 B.n415 10.6151
R1861 B.n416 B.n405 10.6151
R1862 B.n422 B.n405 10.6151
R1863 B.n423 B.n422 10.6151
R1864 B.n424 B.n423 10.6151
R1865 B.n424 B.n403 10.6151
R1866 B.n430 B.n403 10.6151
R1867 B.n431 B.n430 10.6151
R1868 B.n432 B.n431 10.6151
R1869 B.n432 B.n401 10.6151
R1870 B.n438 B.n401 10.6151
R1871 B.n439 B.n438 10.6151
R1872 B.n440 B.n439 10.6151
R1873 B.n440 B.n399 10.6151
R1874 B.n446 B.n399 10.6151
R1875 B.n447 B.n446 10.6151
R1876 B.n448 B.n447 10.6151
R1877 B.n448 B.n397 10.6151
R1878 B.n454 B.n397 10.6151
R1879 B.n455 B.n454 10.6151
R1880 B.n456 B.n455 10.6151
R1881 B.n456 B.n395 10.6151
R1882 B.n462 B.n395 10.6151
R1883 B.n463 B.n462 10.6151
R1884 B.n464 B.n463 10.6151
R1885 B.n464 B.n393 10.6151
R1886 B.n470 B.n393 10.6151
R1887 B.n473 B.n472 10.6151
R1888 B.n473 B.n389 10.6151
R1889 B.n479 B.n389 10.6151
R1890 B.n480 B.n479 10.6151
R1891 B.n481 B.n480 10.6151
R1892 B.n481 B.n387 10.6151
R1893 B.n487 B.n387 10.6151
R1894 B.n488 B.n487 10.6151
R1895 B.n492 B.n488 10.6151
R1896 B.n498 B.n385 10.6151
R1897 B.n499 B.n498 10.6151
R1898 B.n500 B.n499 10.6151
R1899 B.n500 B.n383 10.6151
R1900 B.n506 B.n383 10.6151
R1901 B.n507 B.n506 10.6151
R1902 B.n508 B.n507 10.6151
R1903 B.n508 B.n381 10.6151
R1904 B.n514 B.n381 10.6151
R1905 B.n515 B.n514 10.6151
R1906 B.n516 B.n515 10.6151
R1907 B.n516 B.n379 10.6151
R1908 B.n522 B.n379 10.6151
R1909 B.n523 B.n522 10.6151
R1910 B.n524 B.n523 10.6151
R1911 B.n524 B.n377 10.6151
R1912 B.n530 B.n377 10.6151
R1913 B.n531 B.n530 10.6151
R1914 B.n532 B.n531 10.6151
R1915 B.n532 B.n375 10.6151
R1916 B.n538 B.n375 10.6151
R1917 B.n539 B.n538 10.6151
R1918 B.n540 B.n539 10.6151
R1919 B.n540 B.n373 10.6151
R1920 B.n546 B.n373 10.6151
R1921 B.n547 B.n546 10.6151
R1922 B.n548 B.n547 10.6151
R1923 B.n548 B.n371 10.6151
R1924 B.n371 B.n370 10.6151
R1925 B.n555 B.n370 10.6151
R1926 B.n556 B.n555 10.6151
R1927 B.n562 B.n561 10.6151
R1928 B.n563 B.n562 10.6151
R1929 B.n563 B.n358 10.6151
R1930 B.n573 B.n358 10.6151
R1931 B.n574 B.n573 10.6151
R1932 B.n575 B.n574 10.6151
R1933 B.n575 B.n350 10.6151
R1934 B.n585 B.n350 10.6151
R1935 B.n586 B.n585 10.6151
R1936 B.n587 B.n586 10.6151
R1937 B.n587 B.n342 10.6151
R1938 B.n597 B.n342 10.6151
R1939 B.n598 B.n597 10.6151
R1940 B.n599 B.n598 10.6151
R1941 B.n599 B.n334 10.6151
R1942 B.n609 B.n334 10.6151
R1943 B.n610 B.n609 10.6151
R1944 B.n611 B.n610 10.6151
R1945 B.n611 B.n326 10.6151
R1946 B.n622 B.n326 10.6151
R1947 B.n623 B.n622 10.6151
R1948 B.n624 B.n623 10.6151
R1949 B.n624 B.n319 10.6151
R1950 B.n634 B.n319 10.6151
R1951 B.n635 B.n634 10.6151
R1952 B.n636 B.n635 10.6151
R1953 B.n636 B.n311 10.6151
R1954 B.n646 B.n311 10.6151
R1955 B.n647 B.n646 10.6151
R1956 B.n648 B.n647 10.6151
R1957 B.n648 B.n303 10.6151
R1958 B.n658 B.n303 10.6151
R1959 B.n659 B.n658 10.6151
R1960 B.n660 B.n659 10.6151
R1961 B.n660 B.n295 10.6151
R1962 B.n670 B.n295 10.6151
R1963 B.n671 B.n670 10.6151
R1964 B.n672 B.n671 10.6151
R1965 B.n672 B.n287 10.6151
R1966 B.n683 B.n287 10.6151
R1967 B.n684 B.n683 10.6151
R1968 B.n685 B.n684 10.6151
R1969 B.n685 B.n280 10.6151
R1970 B.n696 B.n280 10.6151
R1971 B.n697 B.n696 10.6151
R1972 B.n698 B.n697 10.6151
R1973 B.n698 B.n0 10.6151
R1974 B.n861 B.n1 10.6151
R1975 B.n861 B.n860 10.6151
R1976 B.n860 B.n859 10.6151
R1977 B.n859 B.n10 10.6151
R1978 B.n853 B.n10 10.6151
R1979 B.n853 B.n852 10.6151
R1980 B.n852 B.n851 10.6151
R1981 B.n851 B.n16 10.6151
R1982 B.n845 B.n16 10.6151
R1983 B.n845 B.n844 10.6151
R1984 B.n844 B.n843 10.6151
R1985 B.n843 B.n24 10.6151
R1986 B.n837 B.n24 10.6151
R1987 B.n837 B.n836 10.6151
R1988 B.n836 B.n835 10.6151
R1989 B.n835 B.n31 10.6151
R1990 B.n829 B.n31 10.6151
R1991 B.n829 B.n828 10.6151
R1992 B.n828 B.n827 10.6151
R1993 B.n827 B.n38 10.6151
R1994 B.n821 B.n38 10.6151
R1995 B.n821 B.n820 10.6151
R1996 B.n820 B.n819 10.6151
R1997 B.n819 B.n45 10.6151
R1998 B.n813 B.n45 10.6151
R1999 B.n813 B.n812 10.6151
R2000 B.n812 B.n811 10.6151
R2001 B.n811 B.n51 10.6151
R2002 B.n805 B.n51 10.6151
R2003 B.n805 B.n804 10.6151
R2004 B.n804 B.n803 10.6151
R2005 B.n803 B.n59 10.6151
R2006 B.n797 B.n59 10.6151
R2007 B.n797 B.n796 10.6151
R2008 B.n796 B.n795 10.6151
R2009 B.n795 B.n66 10.6151
R2010 B.n789 B.n66 10.6151
R2011 B.n789 B.n788 10.6151
R2012 B.n788 B.n787 10.6151
R2013 B.n787 B.n73 10.6151
R2014 B.n781 B.n73 10.6151
R2015 B.n781 B.n780 10.6151
R2016 B.n780 B.n779 10.6151
R2017 B.n779 B.n80 10.6151
R2018 B.n773 B.n80 10.6151
R2019 B.n773 B.n772 10.6151
R2020 B.n772 B.n771 10.6151
R2021 B.n193 B.n132 9.36635
R2022 B.n216 B.n129 9.36635
R2023 B.n471 B.n470 9.36635
R2024 B.n491 B.n385 9.36635
R2025 B.n583 B.t7 4.68301
R2026 B.n785 B.t11 4.68301
R2027 B.n867 B.n0 2.81026
R2028 B.n867 B.n1 2.81026
R2029 B.n196 B.n132 1.24928
R2030 B.n213 B.n129 1.24928
R2031 B.n472 B.n471 1.24928
R2032 B.n492 B.n491 1.24928
R2033 VN.n30 VN.n29 161.3
R2034 VN.n28 VN.n17 161.3
R2035 VN.n27 VN.n26 161.3
R2036 VN.n25 VN.n18 161.3
R2037 VN.n24 VN.n23 161.3
R2038 VN.n22 VN.n19 161.3
R2039 VN.n14 VN.n13 161.3
R2040 VN.n12 VN.n1 161.3
R2041 VN.n11 VN.n10 161.3
R2042 VN.n9 VN.n2 161.3
R2043 VN.n8 VN.n7 161.3
R2044 VN.n6 VN.n3 161.3
R2045 VN.n20 VN.t5 102.338
R2046 VN.n4 VN.t1 102.338
R2047 VN.n15 VN.n0 69.9294
R2048 VN.n31 VN.n16 69.9294
R2049 VN.n5 VN.t4 69.0141
R2050 VN.n0 VN.t3 69.0141
R2051 VN.n21 VN.t2 69.0141
R2052 VN.n16 VN.t0 69.0141
R2053 VN.n11 VN.n2 56.4773
R2054 VN.n27 VN.n18 56.4773
R2055 VN.n21 VN.n20 49.2933
R2056 VN.n5 VN.n4 49.2933
R2057 VN VN.n31 48.4562
R2058 VN.n6 VN.n5 24.3439
R2059 VN.n7 VN.n6 24.3439
R2060 VN.n7 VN.n2 24.3439
R2061 VN.n12 VN.n11 24.3439
R2062 VN.n13 VN.n12 24.3439
R2063 VN.n23 VN.n18 24.3439
R2064 VN.n23 VN.n22 24.3439
R2065 VN.n22 VN.n21 24.3439
R2066 VN.n29 VN.n28 24.3439
R2067 VN.n28 VN.n27 24.3439
R2068 VN.n13 VN.n0 19.9621
R2069 VN.n29 VN.n16 19.9621
R2070 VN.n20 VN.n19 3.92641
R2071 VN.n4 VN.n3 3.92641
R2072 VN.n31 VN.n30 0.355081
R2073 VN.n15 VN.n14 0.355081
R2074 VN VN.n15 0.26685
R2075 VN.n30 VN.n17 0.189894
R2076 VN.n26 VN.n17 0.189894
R2077 VN.n26 VN.n25 0.189894
R2078 VN.n25 VN.n24 0.189894
R2079 VN.n24 VN.n19 0.189894
R2080 VN.n8 VN.n3 0.189894
R2081 VN.n9 VN.n8 0.189894
R2082 VN.n10 VN.n9 0.189894
R2083 VN.n10 VN.n1 0.189894
R2084 VN.n14 VN.n1 0.189894
R2085 VDD2.n91 VDD2.n49 289.615
R2086 VDD2.n42 VDD2.n0 289.615
R2087 VDD2.n92 VDD2.n91 185
R2088 VDD2.n90 VDD2.n89 185
R2089 VDD2.n53 VDD2.n52 185
R2090 VDD2.n84 VDD2.n83 185
R2091 VDD2.n82 VDD2.n81 185
R2092 VDD2.n57 VDD2.n56 185
R2093 VDD2.n76 VDD2.n75 185
R2094 VDD2.n74 VDD2.n73 185
R2095 VDD2.n61 VDD2.n60 185
R2096 VDD2.n68 VDD2.n67 185
R2097 VDD2.n66 VDD2.n65 185
R2098 VDD2.n17 VDD2.n16 185
R2099 VDD2.n19 VDD2.n18 185
R2100 VDD2.n12 VDD2.n11 185
R2101 VDD2.n25 VDD2.n24 185
R2102 VDD2.n27 VDD2.n26 185
R2103 VDD2.n8 VDD2.n7 185
R2104 VDD2.n33 VDD2.n32 185
R2105 VDD2.n35 VDD2.n34 185
R2106 VDD2.n4 VDD2.n3 185
R2107 VDD2.n41 VDD2.n40 185
R2108 VDD2.n43 VDD2.n42 185
R2109 VDD2.n64 VDD2.t5 147.659
R2110 VDD2.n15 VDD2.t4 147.659
R2111 VDD2.n91 VDD2.n90 104.615
R2112 VDD2.n90 VDD2.n52 104.615
R2113 VDD2.n83 VDD2.n52 104.615
R2114 VDD2.n83 VDD2.n82 104.615
R2115 VDD2.n82 VDD2.n56 104.615
R2116 VDD2.n75 VDD2.n56 104.615
R2117 VDD2.n75 VDD2.n74 104.615
R2118 VDD2.n74 VDD2.n60 104.615
R2119 VDD2.n67 VDD2.n60 104.615
R2120 VDD2.n67 VDD2.n66 104.615
R2121 VDD2.n18 VDD2.n17 104.615
R2122 VDD2.n18 VDD2.n11 104.615
R2123 VDD2.n25 VDD2.n11 104.615
R2124 VDD2.n26 VDD2.n25 104.615
R2125 VDD2.n26 VDD2.n7 104.615
R2126 VDD2.n33 VDD2.n7 104.615
R2127 VDD2.n34 VDD2.n33 104.615
R2128 VDD2.n34 VDD2.n3 104.615
R2129 VDD2.n41 VDD2.n3 104.615
R2130 VDD2.n42 VDD2.n41 104.615
R2131 VDD2.n48 VDD2.n47 63.4539
R2132 VDD2 VDD2.n97 63.4512
R2133 VDD2.n66 VDD2.t5 52.3082
R2134 VDD2.n17 VDD2.t4 52.3082
R2135 VDD2.n48 VDD2.n46 49.8499
R2136 VDD2.n96 VDD2.n95 47.7005
R2137 VDD2.n96 VDD2.n48 40.8726
R2138 VDD2.n65 VDD2.n64 15.6677
R2139 VDD2.n16 VDD2.n15 15.6677
R2140 VDD2.n68 VDD2.n63 12.8005
R2141 VDD2.n19 VDD2.n14 12.8005
R2142 VDD2.n69 VDD2.n61 12.0247
R2143 VDD2.n20 VDD2.n12 12.0247
R2144 VDD2.n73 VDD2.n72 11.249
R2145 VDD2.n24 VDD2.n23 11.249
R2146 VDD2.n76 VDD2.n59 10.4732
R2147 VDD2.n27 VDD2.n10 10.4732
R2148 VDD2.n77 VDD2.n57 9.69747
R2149 VDD2.n28 VDD2.n8 9.69747
R2150 VDD2.n95 VDD2.n94 9.45567
R2151 VDD2.n46 VDD2.n45 9.45567
R2152 VDD2.n51 VDD2.n50 9.3005
R2153 VDD2.n94 VDD2.n93 9.3005
R2154 VDD2.n88 VDD2.n87 9.3005
R2155 VDD2.n86 VDD2.n85 9.3005
R2156 VDD2.n55 VDD2.n54 9.3005
R2157 VDD2.n80 VDD2.n79 9.3005
R2158 VDD2.n78 VDD2.n77 9.3005
R2159 VDD2.n59 VDD2.n58 9.3005
R2160 VDD2.n72 VDD2.n71 9.3005
R2161 VDD2.n70 VDD2.n69 9.3005
R2162 VDD2.n63 VDD2.n62 9.3005
R2163 VDD2.n39 VDD2.n38 9.3005
R2164 VDD2.n2 VDD2.n1 9.3005
R2165 VDD2.n45 VDD2.n44 9.3005
R2166 VDD2.n6 VDD2.n5 9.3005
R2167 VDD2.n31 VDD2.n30 9.3005
R2168 VDD2.n29 VDD2.n28 9.3005
R2169 VDD2.n10 VDD2.n9 9.3005
R2170 VDD2.n23 VDD2.n22 9.3005
R2171 VDD2.n21 VDD2.n20 9.3005
R2172 VDD2.n14 VDD2.n13 9.3005
R2173 VDD2.n37 VDD2.n36 9.3005
R2174 VDD2.n95 VDD2.n49 8.92171
R2175 VDD2.n81 VDD2.n80 8.92171
R2176 VDD2.n32 VDD2.n31 8.92171
R2177 VDD2.n46 VDD2.n0 8.92171
R2178 VDD2.n93 VDD2.n92 8.14595
R2179 VDD2.n84 VDD2.n55 8.14595
R2180 VDD2.n35 VDD2.n6 8.14595
R2181 VDD2.n44 VDD2.n43 8.14595
R2182 VDD2.n89 VDD2.n51 7.3702
R2183 VDD2.n85 VDD2.n53 7.3702
R2184 VDD2.n36 VDD2.n4 7.3702
R2185 VDD2.n40 VDD2.n2 7.3702
R2186 VDD2.n89 VDD2.n88 6.59444
R2187 VDD2.n88 VDD2.n53 6.59444
R2188 VDD2.n39 VDD2.n4 6.59444
R2189 VDD2.n40 VDD2.n39 6.59444
R2190 VDD2.n92 VDD2.n51 5.81868
R2191 VDD2.n85 VDD2.n84 5.81868
R2192 VDD2.n36 VDD2.n35 5.81868
R2193 VDD2.n43 VDD2.n2 5.81868
R2194 VDD2.n93 VDD2.n49 5.04292
R2195 VDD2.n81 VDD2.n55 5.04292
R2196 VDD2.n32 VDD2.n6 5.04292
R2197 VDD2.n44 VDD2.n0 5.04292
R2198 VDD2.n64 VDD2.n62 4.38563
R2199 VDD2.n15 VDD2.n13 4.38563
R2200 VDD2.n80 VDD2.n57 4.26717
R2201 VDD2.n31 VDD2.n8 4.26717
R2202 VDD2.n77 VDD2.n76 3.49141
R2203 VDD2.n28 VDD2.n27 3.49141
R2204 VDD2.n73 VDD2.n59 2.71565
R2205 VDD2.n24 VDD2.n10 2.71565
R2206 VDD2 VDD2.n96 2.26343
R2207 VDD2.n97 VDD2.t3 2.2454
R2208 VDD2.n97 VDD2.t0 2.2454
R2209 VDD2.n47 VDD2.t1 2.2454
R2210 VDD2.n47 VDD2.t2 2.2454
R2211 VDD2.n72 VDD2.n61 1.93989
R2212 VDD2.n23 VDD2.n12 1.93989
R2213 VDD2.n69 VDD2.n68 1.16414
R2214 VDD2.n20 VDD2.n19 1.16414
R2215 VDD2.n65 VDD2.n63 0.388379
R2216 VDD2.n16 VDD2.n14 0.388379
R2217 VDD2.n94 VDD2.n50 0.155672
R2218 VDD2.n87 VDD2.n50 0.155672
R2219 VDD2.n87 VDD2.n86 0.155672
R2220 VDD2.n86 VDD2.n54 0.155672
R2221 VDD2.n79 VDD2.n54 0.155672
R2222 VDD2.n79 VDD2.n78 0.155672
R2223 VDD2.n78 VDD2.n58 0.155672
R2224 VDD2.n71 VDD2.n58 0.155672
R2225 VDD2.n71 VDD2.n70 0.155672
R2226 VDD2.n70 VDD2.n62 0.155672
R2227 VDD2.n21 VDD2.n13 0.155672
R2228 VDD2.n22 VDD2.n21 0.155672
R2229 VDD2.n22 VDD2.n9 0.155672
R2230 VDD2.n29 VDD2.n9 0.155672
R2231 VDD2.n30 VDD2.n29 0.155672
R2232 VDD2.n30 VDD2.n5 0.155672
R2233 VDD2.n37 VDD2.n5 0.155672
R2234 VDD2.n38 VDD2.n37 0.155672
R2235 VDD2.n38 VDD2.n1 0.155672
R2236 VDD2.n45 VDD2.n1 0.155672
C0 VN VP 6.81075f
C1 VTAIL VDD1 6.77101f
C2 VDD2 VTAIL 6.82614f
C3 VTAIL VP 5.62742f
C4 VTAIL VN 5.61321f
C5 VDD2 VDD1 1.59448f
C6 VP VDD1 5.53709f
C7 VDD2 VP 0.498549f
C8 VN VDD1 0.15115f
C9 VDD2 VN 5.1923f
C10 VDD2 B 5.795253f
C11 VDD1 B 5.940182f
C12 VTAIL B 6.851472f
C13 VN B 14.05992f
C14 VP B 12.764749f
C15 VDD2.n0 B 0.0317f
C16 VDD2.n1 B 0.02152f
C17 VDD2.n2 B 0.011564f
C18 VDD2.n3 B 0.027332f
C19 VDD2.n4 B 0.012244f
C20 VDD2.n5 B 0.02152f
C21 VDD2.n6 B 0.011564f
C22 VDD2.n7 B 0.027332f
C23 VDD2.n8 B 0.012244f
C24 VDD2.n9 B 0.02152f
C25 VDD2.n10 B 0.011564f
C26 VDD2.n11 B 0.027332f
C27 VDD2.n12 B 0.012244f
C28 VDD2.n13 B 0.790561f
C29 VDD2.n14 B 0.011564f
C30 VDD2.t4 B 0.044622f
C31 VDD2.n15 B 0.107033f
C32 VDD2.n16 B 0.016146f
C33 VDD2.n17 B 0.020499f
C34 VDD2.n18 B 0.027332f
C35 VDD2.n19 B 0.012244f
C36 VDD2.n20 B 0.011564f
C37 VDD2.n21 B 0.02152f
C38 VDD2.n22 B 0.02152f
C39 VDD2.n23 B 0.011564f
C40 VDD2.n24 B 0.012244f
C41 VDD2.n25 B 0.027332f
C42 VDD2.n26 B 0.027332f
C43 VDD2.n27 B 0.012244f
C44 VDD2.n28 B 0.011564f
C45 VDD2.n29 B 0.02152f
C46 VDD2.n30 B 0.02152f
C47 VDD2.n31 B 0.011564f
C48 VDD2.n32 B 0.012244f
C49 VDD2.n33 B 0.027332f
C50 VDD2.n34 B 0.027332f
C51 VDD2.n35 B 0.012244f
C52 VDD2.n36 B 0.011564f
C53 VDD2.n37 B 0.02152f
C54 VDD2.n38 B 0.02152f
C55 VDD2.n39 B 0.011564f
C56 VDD2.n40 B 0.012244f
C57 VDD2.n41 B 0.027332f
C58 VDD2.n42 B 0.061737f
C59 VDD2.n43 B 0.012244f
C60 VDD2.n44 B 0.011564f
C61 VDD2.n45 B 0.047977f
C62 VDD2.n46 B 0.057806f
C63 VDD2.t1 B 0.149988f
C64 VDD2.t2 B 0.149988f
C65 VDD2.n47 B 1.30533f
C66 VDD2.n48 B 2.31859f
C67 VDD2.n49 B 0.0317f
C68 VDD2.n50 B 0.02152f
C69 VDD2.n51 B 0.011564f
C70 VDD2.n52 B 0.027332f
C71 VDD2.n53 B 0.012244f
C72 VDD2.n54 B 0.02152f
C73 VDD2.n55 B 0.011564f
C74 VDD2.n56 B 0.027332f
C75 VDD2.n57 B 0.012244f
C76 VDD2.n58 B 0.02152f
C77 VDD2.n59 B 0.011564f
C78 VDD2.n60 B 0.027332f
C79 VDD2.n61 B 0.012244f
C80 VDD2.n62 B 0.790561f
C81 VDD2.n63 B 0.011564f
C82 VDD2.t5 B 0.044622f
C83 VDD2.n64 B 0.107033f
C84 VDD2.n65 B 0.016146f
C85 VDD2.n66 B 0.020499f
C86 VDD2.n67 B 0.027332f
C87 VDD2.n68 B 0.012244f
C88 VDD2.n69 B 0.011564f
C89 VDD2.n70 B 0.02152f
C90 VDD2.n71 B 0.02152f
C91 VDD2.n72 B 0.011564f
C92 VDD2.n73 B 0.012244f
C93 VDD2.n74 B 0.027332f
C94 VDD2.n75 B 0.027332f
C95 VDD2.n76 B 0.012244f
C96 VDD2.n77 B 0.011564f
C97 VDD2.n78 B 0.02152f
C98 VDD2.n79 B 0.02152f
C99 VDD2.n80 B 0.011564f
C100 VDD2.n81 B 0.012244f
C101 VDD2.n82 B 0.027332f
C102 VDD2.n83 B 0.027332f
C103 VDD2.n84 B 0.012244f
C104 VDD2.n85 B 0.011564f
C105 VDD2.n86 B 0.02152f
C106 VDD2.n87 B 0.02152f
C107 VDD2.n88 B 0.011564f
C108 VDD2.n89 B 0.012244f
C109 VDD2.n90 B 0.027332f
C110 VDD2.n91 B 0.061737f
C111 VDD2.n92 B 0.012244f
C112 VDD2.n93 B 0.011564f
C113 VDD2.n94 B 0.047977f
C114 VDD2.n95 B 0.049627f
C115 VDD2.n96 B 2.10435f
C116 VDD2.t3 B 0.149988f
C117 VDD2.t0 B 0.149988f
C118 VDD2.n97 B 1.30531f
C119 VN.t3 B 1.60546f
C120 VN.n0 B 0.665725f
C121 VN.n1 B 0.021916f
C122 VN.n2 B 0.029366f
C123 VN.n3 B 0.249536f
C124 VN.t4 B 1.60546f
C125 VN.t1 B 1.84405f
C126 VN.n4 B 0.620432f
C127 VN.n5 B 0.659156f
C128 VN.n6 B 0.041051f
C129 VN.n7 B 0.041051f
C130 VN.n8 B 0.021916f
C131 VN.n9 B 0.021916f
C132 VN.n10 B 0.021916f
C133 VN.n11 B 0.034901f
C134 VN.n12 B 0.041051f
C135 VN.n13 B 0.037403f
C136 VN.n14 B 0.035378f
C137 VN.n15 B 0.046156f
C138 VN.t0 B 1.60546f
C139 VN.n16 B 0.665725f
C140 VN.n17 B 0.021916f
C141 VN.n18 B 0.029366f
C142 VN.n19 B 0.249537f
C143 VN.t2 B 1.60546f
C144 VN.t5 B 1.84405f
C145 VN.n20 B 0.620432f
C146 VN.n21 B 0.659156f
C147 VN.n22 B 0.041051f
C148 VN.n23 B 0.041051f
C149 VN.n24 B 0.021916f
C150 VN.n25 B 0.021916f
C151 VN.n26 B 0.021916f
C152 VN.n27 B 0.034901f
C153 VN.n28 B 0.041051f
C154 VN.n29 B 0.037403f
C155 VN.n30 B 0.035378f
C156 VN.n31 B 1.18786f
C157 VTAIL.t10 B 0.176061f
C158 VTAIL.t11 B 0.176061f
C159 VTAIL.n0 B 1.45142f
C160 VTAIL.n1 B 0.476196f
C161 VTAIL.n2 B 0.03721f
C162 VTAIL.n3 B 0.02526f
C163 VTAIL.n4 B 0.013574f
C164 VTAIL.n5 B 0.032084f
C165 VTAIL.n6 B 0.014372f
C166 VTAIL.n7 B 0.02526f
C167 VTAIL.n8 B 0.013574f
C168 VTAIL.n9 B 0.032084f
C169 VTAIL.n10 B 0.014372f
C170 VTAIL.n11 B 0.02526f
C171 VTAIL.n12 B 0.013574f
C172 VTAIL.n13 B 0.032084f
C173 VTAIL.n14 B 0.014372f
C174 VTAIL.n15 B 0.927989f
C175 VTAIL.n16 B 0.013574f
C176 VTAIL.t7 B 0.052379f
C177 VTAIL.n17 B 0.125639f
C178 VTAIL.n18 B 0.018953f
C179 VTAIL.n19 B 0.024063f
C180 VTAIL.n20 B 0.032084f
C181 VTAIL.n21 B 0.014372f
C182 VTAIL.n22 B 0.013574f
C183 VTAIL.n23 B 0.02526f
C184 VTAIL.n24 B 0.02526f
C185 VTAIL.n25 B 0.013574f
C186 VTAIL.n26 B 0.014372f
C187 VTAIL.n27 B 0.032084f
C188 VTAIL.n28 B 0.032084f
C189 VTAIL.n29 B 0.014372f
C190 VTAIL.n30 B 0.013574f
C191 VTAIL.n31 B 0.02526f
C192 VTAIL.n32 B 0.02526f
C193 VTAIL.n33 B 0.013574f
C194 VTAIL.n34 B 0.014372f
C195 VTAIL.n35 B 0.032084f
C196 VTAIL.n36 B 0.032084f
C197 VTAIL.n37 B 0.014372f
C198 VTAIL.n38 B 0.013574f
C199 VTAIL.n39 B 0.02526f
C200 VTAIL.n40 B 0.02526f
C201 VTAIL.n41 B 0.013574f
C202 VTAIL.n42 B 0.014372f
C203 VTAIL.n43 B 0.032084f
C204 VTAIL.n44 B 0.072469f
C205 VTAIL.n45 B 0.014372f
C206 VTAIL.n46 B 0.013574f
C207 VTAIL.n47 B 0.056318f
C208 VTAIL.n48 B 0.040795f
C209 VTAIL.n49 B 0.417556f
C210 VTAIL.t4 B 0.176061f
C211 VTAIL.t5 B 0.176061f
C212 VTAIL.n50 B 1.45142f
C213 VTAIL.n51 B 1.93359f
C214 VTAIL.t2 B 0.176061f
C215 VTAIL.t0 B 0.176061f
C216 VTAIL.n52 B 1.45143f
C217 VTAIL.n53 B 1.93358f
C218 VTAIL.n54 B 0.03721f
C219 VTAIL.n55 B 0.02526f
C220 VTAIL.n56 B 0.013574f
C221 VTAIL.n57 B 0.032084f
C222 VTAIL.n58 B 0.014372f
C223 VTAIL.n59 B 0.02526f
C224 VTAIL.n60 B 0.013574f
C225 VTAIL.n61 B 0.032084f
C226 VTAIL.n62 B 0.014372f
C227 VTAIL.n63 B 0.02526f
C228 VTAIL.n64 B 0.013574f
C229 VTAIL.n65 B 0.032084f
C230 VTAIL.n66 B 0.014372f
C231 VTAIL.n67 B 0.927989f
C232 VTAIL.n68 B 0.013574f
C233 VTAIL.t1 B 0.052379f
C234 VTAIL.n69 B 0.125639f
C235 VTAIL.n70 B 0.018953f
C236 VTAIL.n71 B 0.024063f
C237 VTAIL.n72 B 0.032084f
C238 VTAIL.n73 B 0.014372f
C239 VTAIL.n74 B 0.013574f
C240 VTAIL.n75 B 0.02526f
C241 VTAIL.n76 B 0.02526f
C242 VTAIL.n77 B 0.013574f
C243 VTAIL.n78 B 0.014372f
C244 VTAIL.n79 B 0.032084f
C245 VTAIL.n80 B 0.032084f
C246 VTAIL.n81 B 0.014372f
C247 VTAIL.n82 B 0.013574f
C248 VTAIL.n83 B 0.02526f
C249 VTAIL.n84 B 0.02526f
C250 VTAIL.n85 B 0.013574f
C251 VTAIL.n86 B 0.014372f
C252 VTAIL.n87 B 0.032084f
C253 VTAIL.n88 B 0.032084f
C254 VTAIL.n89 B 0.014372f
C255 VTAIL.n90 B 0.013574f
C256 VTAIL.n91 B 0.02526f
C257 VTAIL.n92 B 0.02526f
C258 VTAIL.n93 B 0.013574f
C259 VTAIL.n94 B 0.014372f
C260 VTAIL.n95 B 0.032084f
C261 VTAIL.n96 B 0.072469f
C262 VTAIL.n97 B 0.014372f
C263 VTAIL.n98 B 0.013574f
C264 VTAIL.n99 B 0.056318f
C265 VTAIL.n100 B 0.040795f
C266 VTAIL.n101 B 0.417556f
C267 VTAIL.t8 B 0.176061f
C268 VTAIL.t9 B 0.176061f
C269 VTAIL.n102 B 1.45143f
C270 VTAIL.n103 B 0.650905f
C271 VTAIL.n104 B 0.03721f
C272 VTAIL.n105 B 0.02526f
C273 VTAIL.n106 B 0.013574f
C274 VTAIL.n107 B 0.032084f
C275 VTAIL.n108 B 0.014372f
C276 VTAIL.n109 B 0.02526f
C277 VTAIL.n110 B 0.013574f
C278 VTAIL.n111 B 0.032084f
C279 VTAIL.n112 B 0.014372f
C280 VTAIL.n113 B 0.02526f
C281 VTAIL.n114 B 0.013574f
C282 VTAIL.n115 B 0.032084f
C283 VTAIL.n116 B 0.014372f
C284 VTAIL.n117 B 0.927989f
C285 VTAIL.n118 B 0.013574f
C286 VTAIL.t6 B 0.052379f
C287 VTAIL.n119 B 0.125639f
C288 VTAIL.n120 B 0.018953f
C289 VTAIL.n121 B 0.024063f
C290 VTAIL.n122 B 0.032084f
C291 VTAIL.n123 B 0.014372f
C292 VTAIL.n124 B 0.013574f
C293 VTAIL.n125 B 0.02526f
C294 VTAIL.n126 B 0.02526f
C295 VTAIL.n127 B 0.013574f
C296 VTAIL.n128 B 0.014372f
C297 VTAIL.n129 B 0.032084f
C298 VTAIL.n130 B 0.032084f
C299 VTAIL.n131 B 0.014372f
C300 VTAIL.n132 B 0.013574f
C301 VTAIL.n133 B 0.02526f
C302 VTAIL.n134 B 0.02526f
C303 VTAIL.n135 B 0.013574f
C304 VTAIL.n136 B 0.014372f
C305 VTAIL.n137 B 0.032084f
C306 VTAIL.n138 B 0.032084f
C307 VTAIL.n139 B 0.014372f
C308 VTAIL.n140 B 0.013574f
C309 VTAIL.n141 B 0.02526f
C310 VTAIL.n142 B 0.02526f
C311 VTAIL.n143 B 0.013574f
C312 VTAIL.n144 B 0.014372f
C313 VTAIL.n145 B 0.032084f
C314 VTAIL.n146 B 0.072469f
C315 VTAIL.n147 B 0.014372f
C316 VTAIL.n148 B 0.013574f
C317 VTAIL.n149 B 0.056318f
C318 VTAIL.n150 B 0.040795f
C319 VTAIL.n151 B 1.46096f
C320 VTAIL.n152 B 0.03721f
C321 VTAIL.n153 B 0.02526f
C322 VTAIL.n154 B 0.013574f
C323 VTAIL.n155 B 0.032084f
C324 VTAIL.n156 B 0.014372f
C325 VTAIL.n157 B 0.02526f
C326 VTAIL.n158 B 0.013574f
C327 VTAIL.n159 B 0.032084f
C328 VTAIL.n160 B 0.014372f
C329 VTAIL.n161 B 0.02526f
C330 VTAIL.n162 B 0.013574f
C331 VTAIL.n163 B 0.032084f
C332 VTAIL.n164 B 0.014372f
C333 VTAIL.n165 B 0.927989f
C334 VTAIL.n166 B 0.013574f
C335 VTAIL.t3 B 0.052379f
C336 VTAIL.n167 B 0.125639f
C337 VTAIL.n168 B 0.018953f
C338 VTAIL.n169 B 0.024063f
C339 VTAIL.n170 B 0.032084f
C340 VTAIL.n171 B 0.014372f
C341 VTAIL.n172 B 0.013574f
C342 VTAIL.n173 B 0.02526f
C343 VTAIL.n174 B 0.02526f
C344 VTAIL.n175 B 0.013574f
C345 VTAIL.n176 B 0.014372f
C346 VTAIL.n177 B 0.032084f
C347 VTAIL.n178 B 0.032084f
C348 VTAIL.n179 B 0.014372f
C349 VTAIL.n180 B 0.013574f
C350 VTAIL.n181 B 0.02526f
C351 VTAIL.n182 B 0.02526f
C352 VTAIL.n183 B 0.013574f
C353 VTAIL.n184 B 0.014372f
C354 VTAIL.n185 B 0.032084f
C355 VTAIL.n186 B 0.032084f
C356 VTAIL.n187 B 0.014372f
C357 VTAIL.n188 B 0.013574f
C358 VTAIL.n189 B 0.02526f
C359 VTAIL.n190 B 0.02526f
C360 VTAIL.n191 B 0.013574f
C361 VTAIL.n192 B 0.014372f
C362 VTAIL.n193 B 0.032084f
C363 VTAIL.n194 B 0.072469f
C364 VTAIL.n195 B 0.014372f
C365 VTAIL.n196 B 0.013574f
C366 VTAIL.n197 B 0.056318f
C367 VTAIL.n198 B 0.040795f
C368 VTAIL.n199 B 1.39641f
C369 VDD1.n0 B 0.032278f
C370 VDD1.n1 B 0.021912f
C371 VDD1.n2 B 0.011775f
C372 VDD1.n3 B 0.027831f
C373 VDD1.n4 B 0.012467f
C374 VDD1.n5 B 0.021912f
C375 VDD1.n6 B 0.011775f
C376 VDD1.n7 B 0.027831f
C377 VDD1.n8 B 0.012467f
C378 VDD1.n9 B 0.021912f
C379 VDD1.n10 B 0.011775f
C380 VDD1.n11 B 0.027831f
C381 VDD1.n12 B 0.012467f
C382 VDD1.n13 B 0.804993f
C383 VDD1.n14 B 0.011775f
C384 VDD1.t1 B 0.045436f
C385 VDD1.n15 B 0.108987f
C386 VDD1.n16 B 0.016441f
C387 VDD1.n17 B 0.020873f
C388 VDD1.n18 B 0.027831f
C389 VDD1.n19 B 0.012467f
C390 VDD1.n20 B 0.011775f
C391 VDD1.n21 B 0.021912f
C392 VDD1.n22 B 0.021912f
C393 VDD1.n23 B 0.011775f
C394 VDD1.n24 B 0.012467f
C395 VDD1.n25 B 0.027831f
C396 VDD1.n26 B 0.027831f
C397 VDD1.n27 B 0.012467f
C398 VDD1.n28 B 0.011775f
C399 VDD1.n29 B 0.021912f
C400 VDD1.n30 B 0.021912f
C401 VDD1.n31 B 0.011775f
C402 VDD1.n32 B 0.012467f
C403 VDD1.n33 B 0.027831f
C404 VDD1.n34 B 0.027831f
C405 VDD1.n35 B 0.012467f
C406 VDD1.n36 B 0.011775f
C407 VDD1.n37 B 0.021912f
C408 VDD1.n38 B 0.021912f
C409 VDD1.n39 B 0.011775f
C410 VDD1.n40 B 0.012467f
C411 VDD1.n41 B 0.027831f
C412 VDD1.n42 B 0.062864f
C413 VDD1.n43 B 0.012467f
C414 VDD1.n44 B 0.011775f
C415 VDD1.n45 B 0.048853f
C416 VDD1.n46 B 0.059634f
C417 VDD1.n47 B 0.032278f
C418 VDD1.n48 B 0.021912f
C419 VDD1.n49 B 0.011775f
C420 VDD1.n50 B 0.027831f
C421 VDD1.n51 B 0.012467f
C422 VDD1.n52 B 0.021912f
C423 VDD1.n53 B 0.011775f
C424 VDD1.n54 B 0.027831f
C425 VDD1.n55 B 0.012467f
C426 VDD1.n56 B 0.021912f
C427 VDD1.n57 B 0.011775f
C428 VDD1.n58 B 0.027831f
C429 VDD1.n59 B 0.012467f
C430 VDD1.n60 B 0.804993f
C431 VDD1.n61 B 0.011775f
C432 VDD1.t4 B 0.045436f
C433 VDD1.n62 B 0.108987f
C434 VDD1.n63 B 0.016441f
C435 VDD1.n64 B 0.020873f
C436 VDD1.n65 B 0.027831f
C437 VDD1.n66 B 0.012467f
C438 VDD1.n67 B 0.011775f
C439 VDD1.n68 B 0.021912f
C440 VDD1.n69 B 0.021912f
C441 VDD1.n70 B 0.011775f
C442 VDD1.n71 B 0.012467f
C443 VDD1.n72 B 0.027831f
C444 VDD1.n73 B 0.027831f
C445 VDD1.n74 B 0.012467f
C446 VDD1.n75 B 0.011775f
C447 VDD1.n76 B 0.021912f
C448 VDD1.n77 B 0.021912f
C449 VDD1.n78 B 0.011775f
C450 VDD1.n79 B 0.012467f
C451 VDD1.n80 B 0.027831f
C452 VDD1.n81 B 0.027831f
C453 VDD1.n82 B 0.012467f
C454 VDD1.n83 B 0.011775f
C455 VDD1.n84 B 0.021912f
C456 VDD1.n85 B 0.021912f
C457 VDD1.n86 B 0.011775f
C458 VDD1.n87 B 0.012467f
C459 VDD1.n88 B 0.027831f
C460 VDD1.n89 B 0.062864f
C461 VDD1.n90 B 0.012467f
C462 VDD1.n91 B 0.011775f
C463 VDD1.n92 B 0.048853f
C464 VDD1.n93 B 0.058861f
C465 VDD1.t3 B 0.152726f
C466 VDD1.t0 B 0.152726f
C467 VDD1.n94 B 1.32916f
C468 VDD1.n95 B 2.4782f
C469 VDD1.t2 B 0.152726f
C470 VDD1.t5 B 0.152726f
C471 VDD1.n96 B 1.32435f
C472 VDD1.n97 B 2.35426f
C473 VP.t2 B 1.63569f
C474 VP.n0 B 0.67826f
C475 VP.n1 B 0.022329f
C476 VP.n2 B 0.029919f
C477 VP.n3 B 0.022329f
C478 VP.t4 B 1.63569f
C479 VP.n4 B 0.041824f
C480 VP.n5 B 0.022329f
C481 VP.n6 B 0.041824f
C482 VP.t3 B 1.63569f
C483 VP.n7 B 0.67826f
C484 VP.n8 B 0.022329f
C485 VP.n9 B 0.029919f
C486 VP.n10 B 0.254235f
C487 VP.t0 B 1.63569f
C488 VP.t1 B 1.87877f
C489 VP.n11 B 0.632115f
C490 VP.n12 B 0.671568f
C491 VP.n13 B 0.041824f
C492 VP.n14 B 0.041824f
C493 VP.n15 B 0.022329f
C494 VP.n16 B 0.022329f
C495 VP.n17 B 0.022329f
C496 VP.n18 B 0.035558f
C497 VP.n19 B 0.041824f
C498 VP.n20 B 0.038107f
C499 VP.n21 B 0.036044f
C500 VP.n22 B 1.20097f
C501 VP.n23 B 1.21755f
C502 VP.t5 B 1.63569f
C503 VP.n24 B 0.67826f
C504 VP.n25 B 0.038107f
C505 VP.n26 B 0.036044f
C506 VP.n27 B 0.022329f
C507 VP.n28 B 0.022329f
C508 VP.n29 B 0.035558f
C509 VP.n30 B 0.029919f
C510 VP.n31 B 0.041824f
C511 VP.n32 B 0.022329f
C512 VP.n33 B 0.022329f
C513 VP.n34 B 0.022329f
C514 VP.n35 B 0.608468f
C515 VP.n36 B 0.041824f
C516 VP.n37 B 0.041824f
C517 VP.n38 B 0.022329f
C518 VP.n39 B 0.022329f
C519 VP.n40 B 0.022329f
C520 VP.n41 B 0.035558f
C521 VP.n42 B 0.041824f
C522 VP.n43 B 0.038107f
C523 VP.n44 B 0.036044f
C524 VP.n45 B 0.047025f
.ends

