* NGSPICE file created from diff_pair_sample_1151.ext - technology: sky130A

.subckt diff_pair_sample_1151 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t1 VN.t0 VTAIL.t3 w_n1734_n4250# sky130_fd_pr__pfet_01v8 ad=6.3999 pd=33.6 as=6.3999 ps=33.6 w=16.41 l=1.58
X1 VDD1.t1 VP.t0 VTAIL.t1 w_n1734_n4250# sky130_fd_pr__pfet_01v8 ad=6.3999 pd=33.6 as=6.3999 ps=33.6 w=16.41 l=1.58
X2 VDD1.t0 VP.t1 VTAIL.t0 w_n1734_n4250# sky130_fd_pr__pfet_01v8 ad=6.3999 pd=33.6 as=6.3999 ps=33.6 w=16.41 l=1.58
X3 B.t11 B.t9 B.t10 w_n1734_n4250# sky130_fd_pr__pfet_01v8 ad=6.3999 pd=33.6 as=0 ps=0 w=16.41 l=1.58
X4 VDD2.t0 VN.t1 VTAIL.t2 w_n1734_n4250# sky130_fd_pr__pfet_01v8 ad=6.3999 pd=33.6 as=6.3999 ps=33.6 w=16.41 l=1.58
X5 B.t8 B.t6 B.t7 w_n1734_n4250# sky130_fd_pr__pfet_01v8 ad=6.3999 pd=33.6 as=0 ps=0 w=16.41 l=1.58
X6 B.t5 B.t3 B.t4 w_n1734_n4250# sky130_fd_pr__pfet_01v8 ad=6.3999 pd=33.6 as=0 ps=0 w=16.41 l=1.58
X7 B.t2 B.t0 B.t1 w_n1734_n4250# sky130_fd_pr__pfet_01v8 ad=6.3999 pd=33.6 as=0 ps=0 w=16.41 l=1.58
R0 VN VN.t1 401.502
R1 VN VN.t0 356.07
R2 VTAIL.n1 VTAIL.t2 54.3117
R3 VTAIL.n3 VTAIL.t3 54.3114
R4 VTAIL.n0 VTAIL.t0 54.3114
R5 VTAIL.n2 VTAIL.t1 54.3114
R6 VTAIL.n1 VTAIL.n0 29.8065
R7 VTAIL.n3 VTAIL.n2 28.16
R8 VTAIL.n2 VTAIL.n1 1.2936
R9 VTAIL VTAIL.n0 0.940155
R10 VTAIL VTAIL.n3 0.353948
R11 VDD2.n0 VDD2.t1 112.09
R12 VDD2.n0 VDD2.t0 70.9902
R13 VDD2 VDD2.n0 0.470328
R14 VP.n0 VP.t0 401.216
R15 VP.n0 VP.t1 355.923
R16 VP VP.n0 0.146778
R17 VDD1 VDD1.t0 113.025
R18 VDD1 VDD1.t1 71.46
R19 B.n374 B.n95 585
R20 B.n373 B.n372 585
R21 B.n371 B.n96 585
R22 B.n370 B.n369 585
R23 B.n368 B.n97 585
R24 B.n367 B.n366 585
R25 B.n365 B.n98 585
R26 B.n364 B.n363 585
R27 B.n362 B.n99 585
R28 B.n361 B.n360 585
R29 B.n359 B.n100 585
R30 B.n358 B.n357 585
R31 B.n356 B.n101 585
R32 B.n355 B.n354 585
R33 B.n353 B.n102 585
R34 B.n352 B.n351 585
R35 B.n350 B.n103 585
R36 B.n349 B.n348 585
R37 B.n347 B.n104 585
R38 B.n346 B.n345 585
R39 B.n344 B.n105 585
R40 B.n343 B.n342 585
R41 B.n341 B.n106 585
R42 B.n340 B.n339 585
R43 B.n338 B.n107 585
R44 B.n337 B.n336 585
R45 B.n335 B.n108 585
R46 B.n334 B.n333 585
R47 B.n332 B.n109 585
R48 B.n331 B.n330 585
R49 B.n329 B.n110 585
R50 B.n328 B.n327 585
R51 B.n326 B.n111 585
R52 B.n325 B.n324 585
R53 B.n323 B.n112 585
R54 B.n322 B.n321 585
R55 B.n320 B.n113 585
R56 B.n319 B.n318 585
R57 B.n317 B.n114 585
R58 B.n316 B.n315 585
R59 B.n314 B.n115 585
R60 B.n313 B.n312 585
R61 B.n311 B.n116 585
R62 B.n310 B.n309 585
R63 B.n308 B.n117 585
R64 B.n307 B.n306 585
R65 B.n305 B.n118 585
R66 B.n304 B.n303 585
R67 B.n302 B.n119 585
R68 B.n301 B.n300 585
R69 B.n299 B.n120 585
R70 B.n298 B.n297 585
R71 B.n296 B.n121 585
R72 B.n295 B.n294 585
R73 B.n293 B.n122 585
R74 B.n292 B.n291 585
R75 B.n287 B.n123 585
R76 B.n286 B.n285 585
R77 B.n284 B.n124 585
R78 B.n283 B.n282 585
R79 B.n281 B.n125 585
R80 B.n280 B.n279 585
R81 B.n278 B.n126 585
R82 B.n277 B.n276 585
R83 B.n274 B.n127 585
R84 B.n273 B.n272 585
R85 B.n271 B.n130 585
R86 B.n270 B.n269 585
R87 B.n268 B.n131 585
R88 B.n267 B.n266 585
R89 B.n265 B.n132 585
R90 B.n264 B.n263 585
R91 B.n262 B.n133 585
R92 B.n261 B.n260 585
R93 B.n259 B.n134 585
R94 B.n258 B.n257 585
R95 B.n256 B.n135 585
R96 B.n255 B.n254 585
R97 B.n253 B.n136 585
R98 B.n252 B.n251 585
R99 B.n250 B.n137 585
R100 B.n249 B.n248 585
R101 B.n247 B.n138 585
R102 B.n246 B.n245 585
R103 B.n244 B.n139 585
R104 B.n243 B.n242 585
R105 B.n241 B.n140 585
R106 B.n240 B.n239 585
R107 B.n238 B.n141 585
R108 B.n237 B.n236 585
R109 B.n235 B.n142 585
R110 B.n234 B.n233 585
R111 B.n232 B.n143 585
R112 B.n231 B.n230 585
R113 B.n229 B.n144 585
R114 B.n228 B.n227 585
R115 B.n226 B.n145 585
R116 B.n225 B.n224 585
R117 B.n223 B.n146 585
R118 B.n222 B.n221 585
R119 B.n220 B.n147 585
R120 B.n219 B.n218 585
R121 B.n217 B.n148 585
R122 B.n216 B.n215 585
R123 B.n214 B.n149 585
R124 B.n213 B.n212 585
R125 B.n211 B.n150 585
R126 B.n210 B.n209 585
R127 B.n208 B.n151 585
R128 B.n207 B.n206 585
R129 B.n205 B.n152 585
R130 B.n204 B.n203 585
R131 B.n202 B.n153 585
R132 B.n201 B.n200 585
R133 B.n199 B.n154 585
R134 B.n198 B.n197 585
R135 B.n196 B.n155 585
R136 B.n195 B.n194 585
R137 B.n193 B.n156 585
R138 B.n376 B.n375 585
R139 B.n377 B.n94 585
R140 B.n379 B.n378 585
R141 B.n380 B.n93 585
R142 B.n382 B.n381 585
R143 B.n383 B.n92 585
R144 B.n385 B.n384 585
R145 B.n386 B.n91 585
R146 B.n388 B.n387 585
R147 B.n389 B.n90 585
R148 B.n391 B.n390 585
R149 B.n392 B.n89 585
R150 B.n394 B.n393 585
R151 B.n395 B.n88 585
R152 B.n397 B.n396 585
R153 B.n398 B.n87 585
R154 B.n400 B.n399 585
R155 B.n401 B.n86 585
R156 B.n403 B.n402 585
R157 B.n404 B.n85 585
R158 B.n406 B.n405 585
R159 B.n407 B.n84 585
R160 B.n409 B.n408 585
R161 B.n410 B.n83 585
R162 B.n412 B.n411 585
R163 B.n413 B.n82 585
R164 B.n415 B.n414 585
R165 B.n416 B.n81 585
R166 B.n418 B.n417 585
R167 B.n419 B.n80 585
R168 B.n421 B.n420 585
R169 B.n422 B.n79 585
R170 B.n424 B.n423 585
R171 B.n425 B.n78 585
R172 B.n427 B.n426 585
R173 B.n428 B.n77 585
R174 B.n430 B.n429 585
R175 B.n431 B.n76 585
R176 B.n433 B.n432 585
R177 B.n434 B.n75 585
R178 B.n615 B.n614 585
R179 B.n613 B.n12 585
R180 B.n612 B.n611 585
R181 B.n610 B.n13 585
R182 B.n609 B.n608 585
R183 B.n607 B.n14 585
R184 B.n606 B.n605 585
R185 B.n604 B.n15 585
R186 B.n603 B.n602 585
R187 B.n601 B.n16 585
R188 B.n600 B.n599 585
R189 B.n598 B.n17 585
R190 B.n597 B.n596 585
R191 B.n595 B.n18 585
R192 B.n594 B.n593 585
R193 B.n592 B.n19 585
R194 B.n591 B.n590 585
R195 B.n589 B.n20 585
R196 B.n588 B.n587 585
R197 B.n586 B.n21 585
R198 B.n585 B.n584 585
R199 B.n583 B.n22 585
R200 B.n582 B.n581 585
R201 B.n580 B.n23 585
R202 B.n579 B.n578 585
R203 B.n577 B.n24 585
R204 B.n576 B.n575 585
R205 B.n574 B.n25 585
R206 B.n573 B.n572 585
R207 B.n571 B.n26 585
R208 B.n570 B.n569 585
R209 B.n568 B.n27 585
R210 B.n567 B.n566 585
R211 B.n565 B.n28 585
R212 B.n564 B.n563 585
R213 B.n562 B.n29 585
R214 B.n561 B.n560 585
R215 B.n559 B.n30 585
R216 B.n558 B.n557 585
R217 B.n556 B.n31 585
R218 B.n555 B.n554 585
R219 B.n553 B.n32 585
R220 B.n552 B.n551 585
R221 B.n550 B.n33 585
R222 B.n549 B.n548 585
R223 B.n547 B.n34 585
R224 B.n546 B.n545 585
R225 B.n544 B.n35 585
R226 B.n543 B.n542 585
R227 B.n541 B.n36 585
R228 B.n540 B.n539 585
R229 B.n538 B.n37 585
R230 B.n537 B.n536 585
R231 B.n535 B.n38 585
R232 B.n534 B.n533 585
R233 B.n531 B.n39 585
R234 B.n530 B.n529 585
R235 B.n528 B.n42 585
R236 B.n527 B.n526 585
R237 B.n525 B.n43 585
R238 B.n524 B.n523 585
R239 B.n522 B.n44 585
R240 B.n521 B.n520 585
R241 B.n519 B.n45 585
R242 B.n517 B.n516 585
R243 B.n515 B.n48 585
R244 B.n514 B.n513 585
R245 B.n512 B.n49 585
R246 B.n511 B.n510 585
R247 B.n509 B.n50 585
R248 B.n508 B.n507 585
R249 B.n506 B.n51 585
R250 B.n505 B.n504 585
R251 B.n503 B.n52 585
R252 B.n502 B.n501 585
R253 B.n500 B.n53 585
R254 B.n499 B.n498 585
R255 B.n497 B.n54 585
R256 B.n496 B.n495 585
R257 B.n494 B.n55 585
R258 B.n493 B.n492 585
R259 B.n491 B.n56 585
R260 B.n490 B.n489 585
R261 B.n488 B.n57 585
R262 B.n487 B.n486 585
R263 B.n485 B.n58 585
R264 B.n484 B.n483 585
R265 B.n482 B.n59 585
R266 B.n481 B.n480 585
R267 B.n479 B.n60 585
R268 B.n478 B.n477 585
R269 B.n476 B.n61 585
R270 B.n475 B.n474 585
R271 B.n473 B.n62 585
R272 B.n472 B.n471 585
R273 B.n470 B.n63 585
R274 B.n469 B.n468 585
R275 B.n467 B.n64 585
R276 B.n466 B.n465 585
R277 B.n464 B.n65 585
R278 B.n463 B.n462 585
R279 B.n461 B.n66 585
R280 B.n460 B.n459 585
R281 B.n458 B.n67 585
R282 B.n457 B.n456 585
R283 B.n455 B.n68 585
R284 B.n454 B.n453 585
R285 B.n452 B.n69 585
R286 B.n451 B.n450 585
R287 B.n449 B.n70 585
R288 B.n448 B.n447 585
R289 B.n446 B.n71 585
R290 B.n445 B.n444 585
R291 B.n443 B.n72 585
R292 B.n442 B.n441 585
R293 B.n440 B.n73 585
R294 B.n439 B.n438 585
R295 B.n437 B.n74 585
R296 B.n436 B.n435 585
R297 B.n616 B.n11 585
R298 B.n618 B.n617 585
R299 B.n619 B.n10 585
R300 B.n621 B.n620 585
R301 B.n622 B.n9 585
R302 B.n624 B.n623 585
R303 B.n625 B.n8 585
R304 B.n627 B.n626 585
R305 B.n628 B.n7 585
R306 B.n630 B.n629 585
R307 B.n631 B.n6 585
R308 B.n633 B.n632 585
R309 B.n634 B.n5 585
R310 B.n636 B.n635 585
R311 B.n637 B.n4 585
R312 B.n639 B.n638 585
R313 B.n640 B.n3 585
R314 B.n642 B.n641 585
R315 B.n643 B.n0 585
R316 B.n2 B.n1 585
R317 B.n166 B.n165 585
R318 B.n168 B.n167 585
R319 B.n169 B.n164 585
R320 B.n171 B.n170 585
R321 B.n172 B.n163 585
R322 B.n174 B.n173 585
R323 B.n175 B.n162 585
R324 B.n177 B.n176 585
R325 B.n178 B.n161 585
R326 B.n180 B.n179 585
R327 B.n181 B.n160 585
R328 B.n183 B.n182 585
R329 B.n184 B.n159 585
R330 B.n186 B.n185 585
R331 B.n187 B.n158 585
R332 B.n189 B.n188 585
R333 B.n190 B.n157 585
R334 B.n192 B.n191 585
R335 B.n128 B.t9 456.031
R336 B.n288 B.t3 456.031
R337 B.n46 B.t0 456.031
R338 B.n40 B.t6 456.031
R339 B.n193 B.n192 454.062
R340 B.n376 B.n95 454.062
R341 B.n436 B.n75 454.062
R342 B.n614 B.n11 454.062
R343 B.n645 B.n644 256.663
R344 B.n644 B.n643 235.042
R345 B.n644 B.n2 235.042
R346 B.n194 B.n193 163.367
R347 B.n194 B.n155 163.367
R348 B.n198 B.n155 163.367
R349 B.n199 B.n198 163.367
R350 B.n200 B.n199 163.367
R351 B.n200 B.n153 163.367
R352 B.n204 B.n153 163.367
R353 B.n205 B.n204 163.367
R354 B.n206 B.n205 163.367
R355 B.n206 B.n151 163.367
R356 B.n210 B.n151 163.367
R357 B.n211 B.n210 163.367
R358 B.n212 B.n211 163.367
R359 B.n212 B.n149 163.367
R360 B.n216 B.n149 163.367
R361 B.n217 B.n216 163.367
R362 B.n218 B.n217 163.367
R363 B.n218 B.n147 163.367
R364 B.n222 B.n147 163.367
R365 B.n223 B.n222 163.367
R366 B.n224 B.n223 163.367
R367 B.n224 B.n145 163.367
R368 B.n228 B.n145 163.367
R369 B.n229 B.n228 163.367
R370 B.n230 B.n229 163.367
R371 B.n230 B.n143 163.367
R372 B.n234 B.n143 163.367
R373 B.n235 B.n234 163.367
R374 B.n236 B.n235 163.367
R375 B.n236 B.n141 163.367
R376 B.n240 B.n141 163.367
R377 B.n241 B.n240 163.367
R378 B.n242 B.n241 163.367
R379 B.n242 B.n139 163.367
R380 B.n246 B.n139 163.367
R381 B.n247 B.n246 163.367
R382 B.n248 B.n247 163.367
R383 B.n248 B.n137 163.367
R384 B.n252 B.n137 163.367
R385 B.n253 B.n252 163.367
R386 B.n254 B.n253 163.367
R387 B.n254 B.n135 163.367
R388 B.n258 B.n135 163.367
R389 B.n259 B.n258 163.367
R390 B.n260 B.n259 163.367
R391 B.n260 B.n133 163.367
R392 B.n264 B.n133 163.367
R393 B.n265 B.n264 163.367
R394 B.n266 B.n265 163.367
R395 B.n266 B.n131 163.367
R396 B.n270 B.n131 163.367
R397 B.n271 B.n270 163.367
R398 B.n272 B.n271 163.367
R399 B.n272 B.n127 163.367
R400 B.n277 B.n127 163.367
R401 B.n278 B.n277 163.367
R402 B.n279 B.n278 163.367
R403 B.n279 B.n125 163.367
R404 B.n283 B.n125 163.367
R405 B.n284 B.n283 163.367
R406 B.n285 B.n284 163.367
R407 B.n285 B.n123 163.367
R408 B.n292 B.n123 163.367
R409 B.n293 B.n292 163.367
R410 B.n294 B.n293 163.367
R411 B.n294 B.n121 163.367
R412 B.n298 B.n121 163.367
R413 B.n299 B.n298 163.367
R414 B.n300 B.n299 163.367
R415 B.n300 B.n119 163.367
R416 B.n304 B.n119 163.367
R417 B.n305 B.n304 163.367
R418 B.n306 B.n305 163.367
R419 B.n306 B.n117 163.367
R420 B.n310 B.n117 163.367
R421 B.n311 B.n310 163.367
R422 B.n312 B.n311 163.367
R423 B.n312 B.n115 163.367
R424 B.n316 B.n115 163.367
R425 B.n317 B.n316 163.367
R426 B.n318 B.n317 163.367
R427 B.n318 B.n113 163.367
R428 B.n322 B.n113 163.367
R429 B.n323 B.n322 163.367
R430 B.n324 B.n323 163.367
R431 B.n324 B.n111 163.367
R432 B.n328 B.n111 163.367
R433 B.n329 B.n328 163.367
R434 B.n330 B.n329 163.367
R435 B.n330 B.n109 163.367
R436 B.n334 B.n109 163.367
R437 B.n335 B.n334 163.367
R438 B.n336 B.n335 163.367
R439 B.n336 B.n107 163.367
R440 B.n340 B.n107 163.367
R441 B.n341 B.n340 163.367
R442 B.n342 B.n341 163.367
R443 B.n342 B.n105 163.367
R444 B.n346 B.n105 163.367
R445 B.n347 B.n346 163.367
R446 B.n348 B.n347 163.367
R447 B.n348 B.n103 163.367
R448 B.n352 B.n103 163.367
R449 B.n353 B.n352 163.367
R450 B.n354 B.n353 163.367
R451 B.n354 B.n101 163.367
R452 B.n358 B.n101 163.367
R453 B.n359 B.n358 163.367
R454 B.n360 B.n359 163.367
R455 B.n360 B.n99 163.367
R456 B.n364 B.n99 163.367
R457 B.n365 B.n364 163.367
R458 B.n366 B.n365 163.367
R459 B.n366 B.n97 163.367
R460 B.n370 B.n97 163.367
R461 B.n371 B.n370 163.367
R462 B.n372 B.n371 163.367
R463 B.n372 B.n95 163.367
R464 B.n432 B.n75 163.367
R465 B.n432 B.n431 163.367
R466 B.n431 B.n430 163.367
R467 B.n430 B.n77 163.367
R468 B.n426 B.n77 163.367
R469 B.n426 B.n425 163.367
R470 B.n425 B.n424 163.367
R471 B.n424 B.n79 163.367
R472 B.n420 B.n79 163.367
R473 B.n420 B.n419 163.367
R474 B.n419 B.n418 163.367
R475 B.n418 B.n81 163.367
R476 B.n414 B.n81 163.367
R477 B.n414 B.n413 163.367
R478 B.n413 B.n412 163.367
R479 B.n412 B.n83 163.367
R480 B.n408 B.n83 163.367
R481 B.n408 B.n407 163.367
R482 B.n407 B.n406 163.367
R483 B.n406 B.n85 163.367
R484 B.n402 B.n85 163.367
R485 B.n402 B.n401 163.367
R486 B.n401 B.n400 163.367
R487 B.n400 B.n87 163.367
R488 B.n396 B.n87 163.367
R489 B.n396 B.n395 163.367
R490 B.n395 B.n394 163.367
R491 B.n394 B.n89 163.367
R492 B.n390 B.n89 163.367
R493 B.n390 B.n389 163.367
R494 B.n389 B.n388 163.367
R495 B.n388 B.n91 163.367
R496 B.n384 B.n91 163.367
R497 B.n384 B.n383 163.367
R498 B.n383 B.n382 163.367
R499 B.n382 B.n93 163.367
R500 B.n378 B.n93 163.367
R501 B.n378 B.n377 163.367
R502 B.n377 B.n376 163.367
R503 B.n614 B.n613 163.367
R504 B.n613 B.n612 163.367
R505 B.n612 B.n13 163.367
R506 B.n608 B.n13 163.367
R507 B.n608 B.n607 163.367
R508 B.n607 B.n606 163.367
R509 B.n606 B.n15 163.367
R510 B.n602 B.n15 163.367
R511 B.n602 B.n601 163.367
R512 B.n601 B.n600 163.367
R513 B.n600 B.n17 163.367
R514 B.n596 B.n17 163.367
R515 B.n596 B.n595 163.367
R516 B.n595 B.n594 163.367
R517 B.n594 B.n19 163.367
R518 B.n590 B.n19 163.367
R519 B.n590 B.n589 163.367
R520 B.n589 B.n588 163.367
R521 B.n588 B.n21 163.367
R522 B.n584 B.n21 163.367
R523 B.n584 B.n583 163.367
R524 B.n583 B.n582 163.367
R525 B.n582 B.n23 163.367
R526 B.n578 B.n23 163.367
R527 B.n578 B.n577 163.367
R528 B.n577 B.n576 163.367
R529 B.n576 B.n25 163.367
R530 B.n572 B.n25 163.367
R531 B.n572 B.n571 163.367
R532 B.n571 B.n570 163.367
R533 B.n570 B.n27 163.367
R534 B.n566 B.n27 163.367
R535 B.n566 B.n565 163.367
R536 B.n565 B.n564 163.367
R537 B.n564 B.n29 163.367
R538 B.n560 B.n29 163.367
R539 B.n560 B.n559 163.367
R540 B.n559 B.n558 163.367
R541 B.n558 B.n31 163.367
R542 B.n554 B.n31 163.367
R543 B.n554 B.n553 163.367
R544 B.n553 B.n552 163.367
R545 B.n552 B.n33 163.367
R546 B.n548 B.n33 163.367
R547 B.n548 B.n547 163.367
R548 B.n547 B.n546 163.367
R549 B.n546 B.n35 163.367
R550 B.n542 B.n35 163.367
R551 B.n542 B.n541 163.367
R552 B.n541 B.n540 163.367
R553 B.n540 B.n37 163.367
R554 B.n536 B.n37 163.367
R555 B.n536 B.n535 163.367
R556 B.n535 B.n534 163.367
R557 B.n534 B.n39 163.367
R558 B.n529 B.n39 163.367
R559 B.n529 B.n528 163.367
R560 B.n528 B.n527 163.367
R561 B.n527 B.n43 163.367
R562 B.n523 B.n43 163.367
R563 B.n523 B.n522 163.367
R564 B.n522 B.n521 163.367
R565 B.n521 B.n45 163.367
R566 B.n516 B.n45 163.367
R567 B.n516 B.n515 163.367
R568 B.n515 B.n514 163.367
R569 B.n514 B.n49 163.367
R570 B.n510 B.n49 163.367
R571 B.n510 B.n509 163.367
R572 B.n509 B.n508 163.367
R573 B.n508 B.n51 163.367
R574 B.n504 B.n51 163.367
R575 B.n504 B.n503 163.367
R576 B.n503 B.n502 163.367
R577 B.n502 B.n53 163.367
R578 B.n498 B.n53 163.367
R579 B.n498 B.n497 163.367
R580 B.n497 B.n496 163.367
R581 B.n496 B.n55 163.367
R582 B.n492 B.n55 163.367
R583 B.n492 B.n491 163.367
R584 B.n491 B.n490 163.367
R585 B.n490 B.n57 163.367
R586 B.n486 B.n57 163.367
R587 B.n486 B.n485 163.367
R588 B.n485 B.n484 163.367
R589 B.n484 B.n59 163.367
R590 B.n480 B.n59 163.367
R591 B.n480 B.n479 163.367
R592 B.n479 B.n478 163.367
R593 B.n478 B.n61 163.367
R594 B.n474 B.n61 163.367
R595 B.n474 B.n473 163.367
R596 B.n473 B.n472 163.367
R597 B.n472 B.n63 163.367
R598 B.n468 B.n63 163.367
R599 B.n468 B.n467 163.367
R600 B.n467 B.n466 163.367
R601 B.n466 B.n65 163.367
R602 B.n462 B.n65 163.367
R603 B.n462 B.n461 163.367
R604 B.n461 B.n460 163.367
R605 B.n460 B.n67 163.367
R606 B.n456 B.n67 163.367
R607 B.n456 B.n455 163.367
R608 B.n455 B.n454 163.367
R609 B.n454 B.n69 163.367
R610 B.n450 B.n69 163.367
R611 B.n450 B.n449 163.367
R612 B.n449 B.n448 163.367
R613 B.n448 B.n71 163.367
R614 B.n444 B.n71 163.367
R615 B.n444 B.n443 163.367
R616 B.n443 B.n442 163.367
R617 B.n442 B.n73 163.367
R618 B.n438 B.n73 163.367
R619 B.n438 B.n437 163.367
R620 B.n437 B.n436 163.367
R621 B.n618 B.n11 163.367
R622 B.n619 B.n618 163.367
R623 B.n620 B.n619 163.367
R624 B.n620 B.n9 163.367
R625 B.n624 B.n9 163.367
R626 B.n625 B.n624 163.367
R627 B.n626 B.n625 163.367
R628 B.n626 B.n7 163.367
R629 B.n630 B.n7 163.367
R630 B.n631 B.n630 163.367
R631 B.n632 B.n631 163.367
R632 B.n632 B.n5 163.367
R633 B.n636 B.n5 163.367
R634 B.n637 B.n636 163.367
R635 B.n638 B.n637 163.367
R636 B.n638 B.n3 163.367
R637 B.n642 B.n3 163.367
R638 B.n643 B.n642 163.367
R639 B.n165 B.n2 163.367
R640 B.n168 B.n165 163.367
R641 B.n169 B.n168 163.367
R642 B.n170 B.n169 163.367
R643 B.n170 B.n163 163.367
R644 B.n174 B.n163 163.367
R645 B.n175 B.n174 163.367
R646 B.n176 B.n175 163.367
R647 B.n176 B.n161 163.367
R648 B.n180 B.n161 163.367
R649 B.n181 B.n180 163.367
R650 B.n182 B.n181 163.367
R651 B.n182 B.n159 163.367
R652 B.n186 B.n159 163.367
R653 B.n187 B.n186 163.367
R654 B.n188 B.n187 163.367
R655 B.n188 B.n157 163.367
R656 B.n192 B.n157 163.367
R657 B.n288 B.t4 145.165
R658 B.n46 B.t2 145.165
R659 B.n128 B.t10 145.143
R660 B.n40 B.t8 145.143
R661 B.n289 B.t5 108.123
R662 B.n47 B.t1 108.123
R663 B.n129 B.t11 108.102
R664 B.n41 B.t7 108.102
R665 B.n275 B.n129 59.5399
R666 B.n290 B.n289 59.5399
R667 B.n518 B.n47 59.5399
R668 B.n532 B.n41 59.5399
R669 B.n129 B.n128 37.0429
R670 B.n289 B.n288 37.0429
R671 B.n47 B.n46 37.0429
R672 B.n41 B.n40 37.0429
R673 B.n616 B.n615 29.5029
R674 B.n435 B.n434 29.5029
R675 B.n375 B.n374 29.5029
R676 B.n191 B.n156 29.5029
R677 B B.n645 18.0485
R678 B.n617 B.n616 10.6151
R679 B.n617 B.n10 10.6151
R680 B.n621 B.n10 10.6151
R681 B.n622 B.n621 10.6151
R682 B.n623 B.n622 10.6151
R683 B.n623 B.n8 10.6151
R684 B.n627 B.n8 10.6151
R685 B.n628 B.n627 10.6151
R686 B.n629 B.n628 10.6151
R687 B.n629 B.n6 10.6151
R688 B.n633 B.n6 10.6151
R689 B.n634 B.n633 10.6151
R690 B.n635 B.n634 10.6151
R691 B.n635 B.n4 10.6151
R692 B.n639 B.n4 10.6151
R693 B.n640 B.n639 10.6151
R694 B.n641 B.n640 10.6151
R695 B.n641 B.n0 10.6151
R696 B.n615 B.n12 10.6151
R697 B.n611 B.n12 10.6151
R698 B.n611 B.n610 10.6151
R699 B.n610 B.n609 10.6151
R700 B.n609 B.n14 10.6151
R701 B.n605 B.n14 10.6151
R702 B.n605 B.n604 10.6151
R703 B.n604 B.n603 10.6151
R704 B.n603 B.n16 10.6151
R705 B.n599 B.n16 10.6151
R706 B.n599 B.n598 10.6151
R707 B.n598 B.n597 10.6151
R708 B.n597 B.n18 10.6151
R709 B.n593 B.n18 10.6151
R710 B.n593 B.n592 10.6151
R711 B.n592 B.n591 10.6151
R712 B.n591 B.n20 10.6151
R713 B.n587 B.n20 10.6151
R714 B.n587 B.n586 10.6151
R715 B.n586 B.n585 10.6151
R716 B.n585 B.n22 10.6151
R717 B.n581 B.n22 10.6151
R718 B.n581 B.n580 10.6151
R719 B.n580 B.n579 10.6151
R720 B.n579 B.n24 10.6151
R721 B.n575 B.n24 10.6151
R722 B.n575 B.n574 10.6151
R723 B.n574 B.n573 10.6151
R724 B.n573 B.n26 10.6151
R725 B.n569 B.n26 10.6151
R726 B.n569 B.n568 10.6151
R727 B.n568 B.n567 10.6151
R728 B.n567 B.n28 10.6151
R729 B.n563 B.n28 10.6151
R730 B.n563 B.n562 10.6151
R731 B.n562 B.n561 10.6151
R732 B.n561 B.n30 10.6151
R733 B.n557 B.n30 10.6151
R734 B.n557 B.n556 10.6151
R735 B.n556 B.n555 10.6151
R736 B.n555 B.n32 10.6151
R737 B.n551 B.n32 10.6151
R738 B.n551 B.n550 10.6151
R739 B.n550 B.n549 10.6151
R740 B.n549 B.n34 10.6151
R741 B.n545 B.n34 10.6151
R742 B.n545 B.n544 10.6151
R743 B.n544 B.n543 10.6151
R744 B.n543 B.n36 10.6151
R745 B.n539 B.n36 10.6151
R746 B.n539 B.n538 10.6151
R747 B.n538 B.n537 10.6151
R748 B.n537 B.n38 10.6151
R749 B.n533 B.n38 10.6151
R750 B.n531 B.n530 10.6151
R751 B.n530 B.n42 10.6151
R752 B.n526 B.n42 10.6151
R753 B.n526 B.n525 10.6151
R754 B.n525 B.n524 10.6151
R755 B.n524 B.n44 10.6151
R756 B.n520 B.n44 10.6151
R757 B.n520 B.n519 10.6151
R758 B.n517 B.n48 10.6151
R759 B.n513 B.n48 10.6151
R760 B.n513 B.n512 10.6151
R761 B.n512 B.n511 10.6151
R762 B.n511 B.n50 10.6151
R763 B.n507 B.n50 10.6151
R764 B.n507 B.n506 10.6151
R765 B.n506 B.n505 10.6151
R766 B.n505 B.n52 10.6151
R767 B.n501 B.n52 10.6151
R768 B.n501 B.n500 10.6151
R769 B.n500 B.n499 10.6151
R770 B.n499 B.n54 10.6151
R771 B.n495 B.n54 10.6151
R772 B.n495 B.n494 10.6151
R773 B.n494 B.n493 10.6151
R774 B.n493 B.n56 10.6151
R775 B.n489 B.n56 10.6151
R776 B.n489 B.n488 10.6151
R777 B.n488 B.n487 10.6151
R778 B.n487 B.n58 10.6151
R779 B.n483 B.n58 10.6151
R780 B.n483 B.n482 10.6151
R781 B.n482 B.n481 10.6151
R782 B.n481 B.n60 10.6151
R783 B.n477 B.n60 10.6151
R784 B.n477 B.n476 10.6151
R785 B.n476 B.n475 10.6151
R786 B.n475 B.n62 10.6151
R787 B.n471 B.n62 10.6151
R788 B.n471 B.n470 10.6151
R789 B.n470 B.n469 10.6151
R790 B.n469 B.n64 10.6151
R791 B.n465 B.n64 10.6151
R792 B.n465 B.n464 10.6151
R793 B.n464 B.n463 10.6151
R794 B.n463 B.n66 10.6151
R795 B.n459 B.n66 10.6151
R796 B.n459 B.n458 10.6151
R797 B.n458 B.n457 10.6151
R798 B.n457 B.n68 10.6151
R799 B.n453 B.n68 10.6151
R800 B.n453 B.n452 10.6151
R801 B.n452 B.n451 10.6151
R802 B.n451 B.n70 10.6151
R803 B.n447 B.n70 10.6151
R804 B.n447 B.n446 10.6151
R805 B.n446 B.n445 10.6151
R806 B.n445 B.n72 10.6151
R807 B.n441 B.n72 10.6151
R808 B.n441 B.n440 10.6151
R809 B.n440 B.n439 10.6151
R810 B.n439 B.n74 10.6151
R811 B.n435 B.n74 10.6151
R812 B.n434 B.n433 10.6151
R813 B.n433 B.n76 10.6151
R814 B.n429 B.n76 10.6151
R815 B.n429 B.n428 10.6151
R816 B.n428 B.n427 10.6151
R817 B.n427 B.n78 10.6151
R818 B.n423 B.n78 10.6151
R819 B.n423 B.n422 10.6151
R820 B.n422 B.n421 10.6151
R821 B.n421 B.n80 10.6151
R822 B.n417 B.n80 10.6151
R823 B.n417 B.n416 10.6151
R824 B.n416 B.n415 10.6151
R825 B.n415 B.n82 10.6151
R826 B.n411 B.n82 10.6151
R827 B.n411 B.n410 10.6151
R828 B.n410 B.n409 10.6151
R829 B.n409 B.n84 10.6151
R830 B.n405 B.n84 10.6151
R831 B.n405 B.n404 10.6151
R832 B.n404 B.n403 10.6151
R833 B.n403 B.n86 10.6151
R834 B.n399 B.n86 10.6151
R835 B.n399 B.n398 10.6151
R836 B.n398 B.n397 10.6151
R837 B.n397 B.n88 10.6151
R838 B.n393 B.n88 10.6151
R839 B.n393 B.n392 10.6151
R840 B.n392 B.n391 10.6151
R841 B.n391 B.n90 10.6151
R842 B.n387 B.n90 10.6151
R843 B.n387 B.n386 10.6151
R844 B.n386 B.n385 10.6151
R845 B.n385 B.n92 10.6151
R846 B.n381 B.n92 10.6151
R847 B.n381 B.n380 10.6151
R848 B.n380 B.n379 10.6151
R849 B.n379 B.n94 10.6151
R850 B.n375 B.n94 10.6151
R851 B.n166 B.n1 10.6151
R852 B.n167 B.n166 10.6151
R853 B.n167 B.n164 10.6151
R854 B.n171 B.n164 10.6151
R855 B.n172 B.n171 10.6151
R856 B.n173 B.n172 10.6151
R857 B.n173 B.n162 10.6151
R858 B.n177 B.n162 10.6151
R859 B.n178 B.n177 10.6151
R860 B.n179 B.n178 10.6151
R861 B.n179 B.n160 10.6151
R862 B.n183 B.n160 10.6151
R863 B.n184 B.n183 10.6151
R864 B.n185 B.n184 10.6151
R865 B.n185 B.n158 10.6151
R866 B.n189 B.n158 10.6151
R867 B.n190 B.n189 10.6151
R868 B.n191 B.n190 10.6151
R869 B.n195 B.n156 10.6151
R870 B.n196 B.n195 10.6151
R871 B.n197 B.n196 10.6151
R872 B.n197 B.n154 10.6151
R873 B.n201 B.n154 10.6151
R874 B.n202 B.n201 10.6151
R875 B.n203 B.n202 10.6151
R876 B.n203 B.n152 10.6151
R877 B.n207 B.n152 10.6151
R878 B.n208 B.n207 10.6151
R879 B.n209 B.n208 10.6151
R880 B.n209 B.n150 10.6151
R881 B.n213 B.n150 10.6151
R882 B.n214 B.n213 10.6151
R883 B.n215 B.n214 10.6151
R884 B.n215 B.n148 10.6151
R885 B.n219 B.n148 10.6151
R886 B.n220 B.n219 10.6151
R887 B.n221 B.n220 10.6151
R888 B.n221 B.n146 10.6151
R889 B.n225 B.n146 10.6151
R890 B.n226 B.n225 10.6151
R891 B.n227 B.n226 10.6151
R892 B.n227 B.n144 10.6151
R893 B.n231 B.n144 10.6151
R894 B.n232 B.n231 10.6151
R895 B.n233 B.n232 10.6151
R896 B.n233 B.n142 10.6151
R897 B.n237 B.n142 10.6151
R898 B.n238 B.n237 10.6151
R899 B.n239 B.n238 10.6151
R900 B.n239 B.n140 10.6151
R901 B.n243 B.n140 10.6151
R902 B.n244 B.n243 10.6151
R903 B.n245 B.n244 10.6151
R904 B.n245 B.n138 10.6151
R905 B.n249 B.n138 10.6151
R906 B.n250 B.n249 10.6151
R907 B.n251 B.n250 10.6151
R908 B.n251 B.n136 10.6151
R909 B.n255 B.n136 10.6151
R910 B.n256 B.n255 10.6151
R911 B.n257 B.n256 10.6151
R912 B.n257 B.n134 10.6151
R913 B.n261 B.n134 10.6151
R914 B.n262 B.n261 10.6151
R915 B.n263 B.n262 10.6151
R916 B.n263 B.n132 10.6151
R917 B.n267 B.n132 10.6151
R918 B.n268 B.n267 10.6151
R919 B.n269 B.n268 10.6151
R920 B.n269 B.n130 10.6151
R921 B.n273 B.n130 10.6151
R922 B.n274 B.n273 10.6151
R923 B.n276 B.n126 10.6151
R924 B.n280 B.n126 10.6151
R925 B.n281 B.n280 10.6151
R926 B.n282 B.n281 10.6151
R927 B.n282 B.n124 10.6151
R928 B.n286 B.n124 10.6151
R929 B.n287 B.n286 10.6151
R930 B.n291 B.n287 10.6151
R931 B.n295 B.n122 10.6151
R932 B.n296 B.n295 10.6151
R933 B.n297 B.n296 10.6151
R934 B.n297 B.n120 10.6151
R935 B.n301 B.n120 10.6151
R936 B.n302 B.n301 10.6151
R937 B.n303 B.n302 10.6151
R938 B.n303 B.n118 10.6151
R939 B.n307 B.n118 10.6151
R940 B.n308 B.n307 10.6151
R941 B.n309 B.n308 10.6151
R942 B.n309 B.n116 10.6151
R943 B.n313 B.n116 10.6151
R944 B.n314 B.n313 10.6151
R945 B.n315 B.n314 10.6151
R946 B.n315 B.n114 10.6151
R947 B.n319 B.n114 10.6151
R948 B.n320 B.n319 10.6151
R949 B.n321 B.n320 10.6151
R950 B.n321 B.n112 10.6151
R951 B.n325 B.n112 10.6151
R952 B.n326 B.n325 10.6151
R953 B.n327 B.n326 10.6151
R954 B.n327 B.n110 10.6151
R955 B.n331 B.n110 10.6151
R956 B.n332 B.n331 10.6151
R957 B.n333 B.n332 10.6151
R958 B.n333 B.n108 10.6151
R959 B.n337 B.n108 10.6151
R960 B.n338 B.n337 10.6151
R961 B.n339 B.n338 10.6151
R962 B.n339 B.n106 10.6151
R963 B.n343 B.n106 10.6151
R964 B.n344 B.n343 10.6151
R965 B.n345 B.n344 10.6151
R966 B.n345 B.n104 10.6151
R967 B.n349 B.n104 10.6151
R968 B.n350 B.n349 10.6151
R969 B.n351 B.n350 10.6151
R970 B.n351 B.n102 10.6151
R971 B.n355 B.n102 10.6151
R972 B.n356 B.n355 10.6151
R973 B.n357 B.n356 10.6151
R974 B.n357 B.n100 10.6151
R975 B.n361 B.n100 10.6151
R976 B.n362 B.n361 10.6151
R977 B.n363 B.n362 10.6151
R978 B.n363 B.n98 10.6151
R979 B.n367 B.n98 10.6151
R980 B.n368 B.n367 10.6151
R981 B.n369 B.n368 10.6151
R982 B.n369 B.n96 10.6151
R983 B.n373 B.n96 10.6151
R984 B.n374 B.n373 10.6151
R985 B.n645 B.n0 8.11757
R986 B.n645 B.n1 8.11757
R987 B.n532 B.n531 6.5566
R988 B.n519 B.n518 6.5566
R989 B.n276 B.n275 6.5566
R990 B.n291 B.n290 6.5566
R991 B.n533 B.n532 4.05904
R992 B.n518 B.n517 4.05904
R993 B.n275 B.n274 4.05904
R994 B.n290 B.n122 4.05904
C0 VDD2 VN 3.36958f
C1 VDD2 VDD1 0.555947f
C2 VN VTAIL 2.77868f
C3 VTAIL VDD1 6.34158f
C4 VP B 1.28473f
C5 VN VDD1 0.147654f
C6 w_n1734_n4250# B 8.94277f
C7 VDD2 B 1.91913f
C8 w_n1734_n4250# VP 2.59735f
C9 VDD2 VP 0.290819f
C10 VTAIL B 4.09787f
C11 VDD2 w_n1734_n4250# 1.99513f
C12 VN B 0.929306f
C13 B VDD1 1.89806f
C14 VTAIL VP 2.7932f
C15 w_n1734_n4250# VTAIL 3.44932f
C16 VN VP 5.78986f
C17 VP VDD1 3.50842f
C18 VDD2 VTAIL 6.38228f
C19 VN w_n1734_n4250# 2.37867f
C20 w_n1734_n4250# VDD1 1.98146f
C21 VDD2 VSUBS 0.951546f
C22 VDD1 VSUBS 4.668389f
C23 VTAIL VSUBS 1.057585f
C24 VN VSUBS 8.52273f
C25 VP VSUBS 1.537298f
C26 B VSUBS 3.51159f
C27 w_n1734_n4250# VSUBS 90.2443f
C28 B.n0 VSUBS 0.005408f
C29 B.n1 VSUBS 0.005408f
C30 B.n2 VSUBS 0.007999f
C31 B.n3 VSUBS 0.006129f
C32 B.n4 VSUBS 0.006129f
C33 B.n5 VSUBS 0.006129f
C34 B.n6 VSUBS 0.006129f
C35 B.n7 VSUBS 0.006129f
C36 B.n8 VSUBS 0.006129f
C37 B.n9 VSUBS 0.006129f
C38 B.n10 VSUBS 0.006129f
C39 B.n11 VSUBS 0.013069f
C40 B.n12 VSUBS 0.006129f
C41 B.n13 VSUBS 0.006129f
C42 B.n14 VSUBS 0.006129f
C43 B.n15 VSUBS 0.006129f
C44 B.n16 VSUBS 0.006129f
C45 B.n17 VSUBS 0.006129f
C46 B.n18 VSUBS 0.006129f
C47 B.n19 VSUBS 0.006129f
C48 B.n20 VSUBS 0.006129f
C49 B.n21 VSUBS 0.006129f
C50 B.n22 VSUBS 0.006129f
C51 B.n23 VSUBS 0.006129f
C52 B.n24 VSUBS 0.006129f
C53 B.n25 VSUBS 0.006129f
C54 B.n26 VSUBS 0.006129f
C55 B.n27 VSUBS 0.006129f
C56 B.n28 VSUBS 0.006129f
C57 B.n29 VSUBS 0.006129f
C58 B.n30 VSUBS 0.006129f
C59 B.n31 VSUBS 0.006129f
C60 B.n32 VSUBS 0.006129f
C61 B.n33 VSUBS 0.006129f
C62 B.n34 VSUBS 0.006129f
C63 B.n35 VSUBS 0.006129f
C64 B.n36 VSUBS 0.006129f
C65 B.n37 VSUBS 0.006129f
C66 B.n38 VSUBS 0.006129f
C67 B.n39 VSUBS 0.006129f
C68 B.t7 VSUBS 0.481804f
C69 B.t8 VSUBS 0.494732f
C70 B.t6 VSUBS 0.975537f
C71 B.n40 VSUBS 0.220871f
C72 B.n41 VSUBS 0.059398f
C73 B.n42 VSUBS 0.006129f
C74 B.n43 VSUBS 0.006129f
C75 B.n44 VSUBS 0.006129f
C76 B.n45 VSUBS 0.006129f
C77 B.t1 VSUBS 0.481788f
C78 B.t2 VSUBS 0.494718f
C79 B.t0 VSUBS 0.975537f
C80 B.n46 VSUBS 0.220885f
C81 B.n47 VSUBS 0.059414f
C82 B.n48 VSUBS 0.006129f
C83 B.n49 VSUBS 0.006129f
C84 B.n50 VSUBS 0.006129f
C85 B.n51 VSUBS 0.006129f
C86 B.n52 VSUBS 0.006129f
C87 B.n53 VSUBS 0.006129f
C88 B.n54 VSUBS 0.006129f
C89 B.n55 VSUBS 0.006129f
C90 B.n56 VSUBS 0.006129f
C91 B.n57 VSUBS 0.006129f
C92 B.n58 VSUBS 0.006129f
C93 B.n59 VSUBS 0.006129f
C94 B.n60 VSUBS 0.006129f
C95 B.n61 VSUBS 0.006129f
C96 B.n62 VSUBS 0.006129f
C97 B.n63 VSUBS 0.006129f
C98 B.n64 VSUBS 0.006129f
C99 B.n65 VSUBS 0.006129f
C100 B.n66 VSUBS 0.006129f
C101 B.n67 VSUBS 0.006129f
C102 B.n68 VSUBS 0.006129f
C103 B.n69 VSUBS 0.006129f
C104 B.n70 VSUBS 0.006129f
C105 B.n71 VSUBS 0.006129f
C106 B.n72 VSUBS 0.006129f
C107 B.n73 VSUBS 0.006129f
C108 B.n74 VSUBS 0.006129f
C109 B.n75 VSUBS 0.013069f
C110 B.n76 VSUBS 0.006129f
C111 B.n77 VSUBS 0.006129f
C112 B.n78 VSUBS 0.006129f
C113 B.n79 VSUBS 0.006129f
C114 B.n80 VSUBS 0.006129f
C115 B.n81 VSUBS 0.006129f
C116 B.n82 VSUBS 0.006129f
C117 B.n83 VSUBS 0.006129f
C118 B.n84 VSUBS 0.006129f
C119 B.n85 VSUBS 0.006129f
C120 B.n86 VSUBS 0.006129f
C121 B.n87 VSUBS 0.006129f
C122 B.n88 VSUBS 0.006129f
C123 B.n89 VSUBS 0.006129f
C124 B.n90 VSUBS 0.006129f
C125 B.n91 VSUBS 0.006129f
C126 B.n92 VSUBS 0.006129f
C127 B.n93 VSUBS 0.006129f
C128 B.n94 VSUBS 0.006129f
C129 B.n95 VSUBS 0.013792f
C130 B.n96 VSUBS 0.006129f
C131 B.n97 VSUBS 0.006129f
C132 B.n98 VSUBS 0.006129f
C133 B.n99 VSUBS 0.006129f
C134 B.n100 VSUBS 0.006129f
C135 B.n101 VSUBS 0.006129f
C136 B.n102 VSUBS 0.006129f
C137 B.n103 VSUBS 0.006129f
C138 B.n104 VSUBS 0.006129f
C139 B.n105 VSUBS 0.006129f
C140 B.n106 VSUBS 0.006129f
C141 B.n107 VSUBS 0.006129f
C142 B.n108 VSUBS 0.006129f
C143 B.n109 VSUBS 0.006129f
C144 B.n110 VSUBS 0.006129f
C145 B.n111 VSUBS 0.006129f
C146 B.n112 VSUBS 0.006129f
C147 B.n113 VSUBS 0.006129f
C148 B.n114 VSUBS 0.006129f
C149 B.n115 VSUBS 0.006129f
C150 B.n116 VSUBS 0.006129f
C151 B.n117 VSUBS 0.006129f
C152 B.n118 VSUBS 0.006129f
C153 B.n119 VSUBS 0.006129f
C154 B.n120 VSUBS 0.006129f
C155 B.n121 VSUBS 0.006129f
C156 B.n122 VSUBS 0.004236f
C157 B.n123 VSUBS 0.006129f
C158 B.n124 VSUBS 0.006129f
C159 B.n125 VSUBS 0.006129f
C160 B.n126 VSUBS 0.006129f
C161 B.n127 VSUBS 0.006129f
C162 B.t11 VSUBS 0.481804f
C163 B.t10 VSUBS 0.494732f
C164 B.t9 VSUBS 0.975537f
C165 B.n128 VSUBS 0.220871f
C166 B.n129 VSUBS 0.059398f
C167 B.n130 VSUBS 0.006129f
C168 B.n131 VSUBS 0.006129f
C169 B.n132 VSUBS 0.006129f
C170 B.n133 VSUBS 0.006129f
C171 B.n134 VSUBS 0.006129f
C172 B.n135 VSUBS 0.006129f
C173 B.n136 VSUBS 0.006129f
C174 B.n137 VSUBS 0.006129f
C175 B.n138 VSUBS 0.006129f
C176 B.n139 VSUBS 0.006129f
C177 B.n140 VSUBS 0.006129f
C178 B.n141 VSUBS 0.006129f
C179 B.n142 VSUBS 0.006129f
C180 B.n143 VSUBS 0.006129f
C181 B.n144 VSUBS 0.006129f
C182 B.n145 VSUBS 0.006129f
C183 B.n146 VSUBS 0.006129f
C184 B.n147 VSUBS 0.006129f
C185 B.n148 VSUBS 0.006129f
C186 B.n149 VSUBS 0.006129f
C187 B.n150 VSUBS 0.006129f
C188 B.n151 VSUBS 0.006129f
C189 B.n152 VSUBS 0.006129f
C190 B.n153 VSUBS 0.006129f
C191 B.n154 VSUBS 0.006129f
C192 B.n155 VSUBS 0.006129f
C193 B.n156 VSUBS 0.013792f
C194 B.n157 VSUBS 0.006129f
C195 B.n158 VSUBS 0.006129f
C196 B.n159 VSUBS 0.006129f
C197 B.n160 VSUBS 0.006129f
C198 B.n161 VSUBS 0.006129f
C199 B.n162 VSUBS 0.006129f
C200 B.n163 VSUBS 0.006129f
C201 B.n164 VSUBS 0.006129f
C202 B.n165 VSUBS 0.006129f
C203 B.n166 VSUBS 0.006129f
C204 B.n167 VSUBS 0.006129f
C205 B.n168 VSUBS 0.006129f
C206 B.n169 VSUBS 0.006129f
C207 B.n170 VSUBS 0.006129f
C208 B.n171 VSUBS 0.006129f
C209 B.n172 VSUBS 0.006129f
C210 B.n173 VSUBS 0.006129f
C211 B.n174 VSUBS 0.006129f
C212 B.n175 VSUBS 0.006129f
C213 B.n176 VSUBS 0.006129f
C214 B.n177 VSUBS 0.006129f
C215 B.n178 VSUBS 0.006129f
C216 B.n179 VSUBS 0.006129f
C217 B.n180 VSUBS 0.006129f
C218 B.n181 VSUBS 0.006129f
C219 B.n182 VSUBS 0.006129f
C220 B.n183 VSUBS 0.006129f
C221 B.n184 VSUBS 0.006129f
C222 B.n185 VSUBS 0.006129f
C223 B.n186 VSUBS 0.006129f
C224 B.n187 VSUBS 0.006129f
C225 B.n188 VSUBS 0.006129f
C226 B.n189 VSUBS 0.006129f
C227 B.n190 VSUBS 0.006129f
C228 B.n191 VSUBS 0.013069f
C229 B.n192 VSUBS 0.013069f
C230 B.n193 VSUBS 0.013792f
C231 B.n194 VSUBS 0.006129f
C232 B.n195 VSUBS 0.006129f
C233 B.n196 VSUBS 0.006129f
C234 B.n197 VSUBS 0.006129f
C235 B.n198 VSUBS 0.006129f
C236 B.n199 VSUBS 0.006129f
C237 B.n200 VSUBS 0.006129f
C238 B.n201 VSUBS 0.006129f
C239 B.n202 VSUBS 0.006129f
C240 B.n203 VSUBS 0.006129f
C241 B.n204 VSUBS 0.006129f
C242 B.n205 VSUBS 0.006129f
C243 B.n206 VSUBS 0.006129f
C244 B.n207 VSUBS 0.006129f
C245 B.n208 VSUBS 0.006129f
C246 B.n209 VSUBS 0.006129f
C247 B.n210 VSUBS 0.006129f
C248 B.n211 VSUBS 0.006129f
C249 B.n212 VSUBS 0.006129f
C250 B.n213 VSUBS 0.006129f
C251 B.n214 VSUBS 0.006129f
C252 B.n215 VSUBS 0.006129f
C253 B.n216 VSUBS 0.006129f
C254 B.n217 VSUBS 0.006129f
C255 B.n218 VSUBS 0.006129f
C256 B.n219 VSUBS 0.006129f
C257 B.n220 VSUBS 0.006129f
C258 B.n221 VSUBS 0.006129f
C259 B.n222 VSUBS 0.006129f
C260 B.n223 VSUBS 0.006129f
C261 B.n224 VSUBS 0.006129f
C262 B.n225 VSUBS 0.006129f
C263 B.n226 VSUBS 0.006129f
C264 B.n227 VSUBS 0.006129f
C265 B.n228 VSUBS 0.006129f
C266 B.n229 VSUBS 0.006129f
C267 B.n230 VSUBS 0.006129f
C268 B.n231 VSUBS 0.006129f
C269 B.n232 VSUBS 0.006129f
C270 B.n233 VSUBS 0.006129f
C271 B.n234 VSUBS 0.006129f
C272 B.n235 VSUBS 0.006129f
C273 B.n236 VSUBS 0.006129f
C274 B.n237 VSUBS 0.006129f
C275 B.n238 VSUBS 0.006129f
C276 B.n239 VSUBS 0.006129f
C277 B.n240 VSUBS 0.006129f
C278 B.n241 VSUBS 0.006129f
C279 B.n242 VSUBS 0.006129f
C280 B.n243 VSUBS 0.006129f
C281 B.n244 VSUBS 0.006129f
C282 B.n245 VSUBS 0.006129f
C283 B.n246 VSUBS 0.006129f
C284 B.n247 VSUBS 0.006129f
C285 B.n248 VSUBS 0.006129f
C286 B.n249 VSUBS 0.006129f
C287 B.n250 VSUBS 0.006129f
C288 B.n251 VSUBS 0.006129f
C289 B.n252 VSUBS 0.006129f
C290 B.n253 VSUBS 0.006129f
C291 B.n254 VSUBS 0.006129f
C292 B.n255 VSUBS 0.006129f
C293 B.n256 VSUBS 0.006129f
C294 B.n257 VSUBS 0.006129f
C295 B.n258 VSUBS 0.006129f
C296 B.n259 VSUBS 0.006129f
C297 B.n260 VSUBS 0.006129f
C298 B.n261 VSUBS 0.006129f
C299 B.n262 VSUBS 0.006129f
C300 B.n263 VSUBS 0.006129f
C301 B.n264 VSUBS 0.006129f
C302 B.n265 VSUBS 0.006129f
C303 B.n266 VSUBS 0.006129f
C304 B.n267 VSUBS 0.006129f
C305 B.n268 VSUBS 0.006129f
C306 B.n269 VSUBS 0.006129f
C307 B.n270 VSUBS 0.006129f
C308 B.n271 VSUBS 0.006129f
C309 B.n272 VSUBS 0.006129f
C310 B.n273 VSUBS 0.006129f
C311 B.n274 VSUBS 0.004236f
C312 B.n275 VSUBS 0.014201f
C313 B.n276 VSUBS 0.004958f
C314 B.n277 VSUBS 0.006129f
C315 B.n278 VSUBS 0.006129f
C316 B.n279 VSUBS 0.006129f
C317 B.n280 VSUBS 0.006129f
C318 B.n281 VSUBS 0.006129f
C319 B.n282 VSUBS 0.006129f
C320 B.n283 VSUBS 0.006129f
C321 B.n284 VSUBS 0.006129f
C322 B.n285 VSUBS 0.006129f
C323 B.n286 VSUBS 0.006129f
C324 B.n287 VSUBS 0.006129f
C325 B.t5 VSUBS 0.481788f
C326 B.t4 VSUBS 0.494718f
C327 B.t3 VSUBS 0.975537f
C328 B.n288 VSUBS 0.220885f
C329 B.n289 VSUBS 0.059414f
C330 B.n290 VSUBS 0.014201f
C331 B.n291 VSUBS 0.004958f
C332 B.n292 VSUBS 0.006129f
C333 B.n293 VSUBS 0.006129f
C334 B.n294 VSUBS 0.006129f
C335 B.n295 VSUBS 0.006129f
C336 B.n296 VSUBS 0.006129f
C337 B.n297 VSUBS 0.006129f
C338 B.n298 VSUBS 0.006129f
C339 B.n299 VSUBS 0.006129f
C340 B.n300 VSUBS 0.006129f
C341 B.n301 VSUBS 0.006129f
C342 B.n302 VSUBS 0.006129f
C343 B.n303 VSUBS 0.006129f
C344 B.n304 VSUBS 0.006129f
C345 B.n305 VSUBS 0.006129f
C346 B.n306 VSUBS 0.006129f
C347 B.n307 VSUBS 0.006129f
C348 B.n308 VSUBS 0.006129f
C349 B.n309 VSUBS 0.006129f
C350 B.n310 VSUBS 0.006129f
C351 B.n311 VSUBS 0.006129f
C352 B.n312 VSUBS 0.006129f
C353 B.n313 VSUBS 0.006129f
C354 B.n314 VSUBS 0.006129f
C355 B.n315 VSUBS 0.006129f
C356 B.n316 VSUBS 0.006129f
C357 B.n317 VSUBS 0.006129f
C358 B.n318 VSUBS 0.006129f
C359 B.n319 VSUBS 0.006129f
C360 B.n320 VSUBS 0.006129f
C361 B.n321 VSUBS 0.006129f
C362 B.n322 VSUBS 0.006129f
C363 B.n323 VSUBS 0.006129f
C364 B.n324 VSUBS 0.006129f
C365 B.n325 VSUBS 0.006129f
C366 B.n326 VSUBS 0.006129f
C367 B.n327 VSUBS 0.006129f
C368 B.n328 VSUBS 0.006129f
C369 B.n329 VSUBS 0.006129f
C370 B.n330 VSUBS 0.006129f
C371 B.n331 VSUBS 0.006129f
C372 B.n332 VSUBS 0.006129f
C373 B.n333 VSUBS 0.006129f
C374 B.n334 VSUBS 0.006129f
C375 B.n335 VSUBS 0.006129f
C376 B.n336 VSUBS 0.006129f
C377 B.n337 VSUBS 0.006129f
C378 B.n338 VSUBS 0.006129f
C379 B.n339 VSUBS 0.006129f
C380 B.n340 VSUBS 0.006129f
C381 B.n341 VSUBS 0.006129f
C382 B.n342 VSUBS 0.006129f
C383 B.n343 VSUBS 0.006129f
C384 B.n344 VSUBS 0.006129f
C385 B.n345 VSUBS 0.006129f
C386 B.n346 VSUBS 0.006129f
C387 B.n347 VSUBS 0.006129f
C388 B.n348 VSUBS 0.006129f
C389 B.n349 VSUBS 0.006129f
C390 B.n350 VSUBS 0.006129f
C391 B.n351 VSUBS 0.006129f
C392 B.n352 VSUBS 0.006129f
C393 B.n353 VSUBS 0.006129f
C394 B.n354 VSUBS 0.006129f
C395 B.n355 VSUBS 0.006129f
C396 B.n356 VSUBS 0.006129f
C397 B.n357 VSUBS 0.006129f
C398 B.n358 VSUBS 0.006129f
C399 B.n359 VSUBS 0.006129f
C400 B.n360 VSUBS 0.006129f
C401 B.n361 VSUBS 0.006129f
C402 B.n362 VSUBS 0.006129f
C403 B.n363 VSUBS 0.006129f
C404 B.n364 VSUBS 0.006129f
C405 B.n365 VSUBS 0.006129f
C406 B.n366 VSUBS 0.006129f
C407 B.n367 VSUBS 0.006129f
C408 B.n368 VSUBS 0.006129f
C409 B.n369 VSUBS 0.006129f
C410 B.n370 VSUBS 0.006129f
C411 B.n371 VSUBS 0.006129f
C412 B.n372 VSUBS 0.006129f
C413 B.n373 VSUBS 0.006129f
C414 B.n374 VSUBS 0.012991f
C415 B.n375 VSUBS 0.01387f
C416 B.n376 VSUBS 0.013069f
C417 B.n377 VSUBS 0.006129f
C418 B.n378 VSUBS 0.006129f
C419 B.n379 VSUBS 0.006129f
C420 B.n380 VSUBS 0.006129f
C421 B.n381 VSUBS 0.006129f
C422 B.n382 VSUBS 0.006129f
C423 B.n383 VSUBS 0.006129f
C424 B.n384 VSUBS 0.006129f
C425 B.n385 VSUBS 0.006129f
C426 B.n386 VSUBS 0.006129f
C427 B.n387 VSUBS 0.006129f
C428 B.n388 VSUBS 0.006129f
C429 B.n389 VSUBS 0.006129f
C430 B.n390 VSUBS 0.006129f
C431 B.n391 VSUBS 0.006129f
C432 B.n392 VSUBS 0.006129f
C433 B.n393 VSUBS 0.006129f
C434 B.n394 VSUBS 0.006129f
C435 B.n395 VSUBS 0.006129f
C436 B.n396 VSUBS 0.006129f
C437 B.n397 VSUBS 0.006129f
C438 B.n398 VSUBS 0.006129f
C439 B.n399 VSUBS 0.006129f
C440 B.n400 VSUBS 0.006129f
C441 B.n401 VSUBS 0.006129f
C442 B.n402 VSUBS 0.006129f
C443 B.n403 VSUBS 0.006129f
C444 B.n404 VSUBS 0.006129f
C445 B.n405 VSUBS 0.006129f
C446 B.n406 VSUBS 0.006129f
C447 B.n407 VSUBS 0.006129f
C448 B.n408 VSUBS 0.006129f
C449 B.n409 VSUBS 0.006129f
C450 B.n410 VSUBS 0.006129f
C451 B.n411 VSUBS 0.006129f
C452 B.n412 VSUBS 0.006129f
C453 B.n413 VSUBS 0.006129f
C454 B.n414 VSUBS 0.006129f
C455 B.n415 VSUBS 0.006129f
C456 B.n416 VSUBS 0.006129f
C457 B.n417 VSUBS 0.006129f
C458 B.n418 VSUBS 0.006129f
C459 B.n419 VSUBS 0.006129f
C460 B.n420 VSUBS 0.006129f
C461 B.n421 VSUBS 0.006129f
C462 B.n422 VSUBS 0.006129f
C463 B.n423 VSUBS 0.006129f
C464 B.n424 VSUBS 0.006129f
C465 B.n425 VSUBS 0.006129f
C466 B.n426 VSUBS 0.006129f
C467 B.n427 VSUBS 0.006129f
C468 B.n428 VSUBS 0.006129f
C469 B.n429 VSUBS 0.006129f
C470 B.n430 VSUBS 0.006129f
C471 B.n431 VSUBS 0.006129f
C472 B.n432 VSUBS 0.006129f
C473 B.n433 VSUBS 0.006129f
C474 B.n434 VSUBS 0.013069f
C475 B.n435 VSUBS 0.013792f
C476 B.n436 VSUBS 0.013792f
C477 B.n437 VSUBS 0.006129f
C478 B.n438 VSUBS 0.006129f
C479 B.n439 VSUBS 0.006129f
C480 B.n440 VSUBS 0.006129f
C481 B.n441 VSUBS 0.006129f
C482 B.n442 VSUBS 0.006129f
C483 B.n443 VSUBS 0.006129f
C484 B.n444 VSUBS 0.006129f
C485 B.n445 VSUBS 0.006129f
C486 B.n446 VSUBS 0.006129f
C487 B.n447 VSUBS 0.006129f
C488 B.n448 VSUBS 0.006129f
C489 B.n449 VSUBS 0.006129f
C490 B.n450 VSUBS 0.006129f
C491 B.n451 VSUBS 0.006129f
C492 B.n452 VSUBS 0.006129f
C493 B.n453 VSUBS 0.006129f
C494 B.n454 VSUBS 0.006129f
C495 B.n455 VSUBS 0.006129f
C496 B.n456 VSUBS 0.006129f
C497 B.n457 VSUBS 0.006129f
C498 B.n458 VSUBS 0.006129f
C499 B.n459 VSUBS 0.006129f
C500 B.n460 VSUBS 0.006129f
C501 B.n461 VSUBS 0.006129f
C502 B.n462 VSUBS 0.006129f
C503 B.n463 VSUBS 0.006129f
C504 B.n464 VSUBS 0.006129f
C505 B.n465 VSUBS 0.006129f
C506 B.n466 VSUBS 0.006129f
C507 B.n467 VSUBS 0.006129f
C508 B.n468 VSUBS 0.006129f
C509 B.n469 VSUBS 0.006129f
C510 B.n470 VSUBS 0.006129f
C511 B.n471 VSUBS 0.006129f
C512 B.n472 VSUBS 0.006129f
C513 B.n473 VSUBS 0.006129f
C514 B.n474 VSUBS 0.006129f
C515 B.n475 VSUBS 0.006129f
C516 B.n476 VSUBS 0.006129f
C517 B.n477 VSUBS 0.006129f
C518 B.n478 VSUBS 0.006129f
C519 B.n479 VSUBS 0.006129f
C520 B.n480 VSUBS 0.006129f
C521 B.n481 VSUBS 0.006129f
C522 B.n482 VSUBS 0.006129f
C523 B.n483 VSUBS 0.006129f
C524 B.n484 VSUBS 0.006129f
C525 B.n485 VSUBS 0.006129f
C526 B.n486 VSUBS 0.006129f
C527 B.n487 VSUBS 0.006129f
C528 B.n488 VSUBS 0.006129f
C529 B.n489 VSUBS 0.006129f
C530 B.n490 VSUBS 0.006129f
C531 B.n491 VSUBS 0.006129f
C532 B.n492 VSUBS 0.006129f
C533 B.n493 VSUBS 0.006129f
C534 B.n494 VSUBS 0.006129f
C535 B.n495 VSUBS 0.006129f
C536 B.n496 VSUBS 0.006129f
C537 B.n497 VSUBS 0.006129f
C538 B.n498 VSUBS 0.006129f
C539 B.n499 VSUBS 0.006129f
C540 B.n500 VSUBS 0.006129f
C541 B.n501 VSUBS 0.006129f
C542 B.n502 VSUBS 0.006129f
C543 B.n503 VSUBS 0.006129f
C544 B.n504 VSUBS 0.006129f
C545 B.n505 VSUBS 0.006129f
C546 B.n506 VSUBS 0.006129f
C547 B.n507 VSUBS 0.006129f
C548 B.n508 VSUBS 0.006129f
C549 B.n509 VSUBS 0.006129f
C550 B.n510 VSUBS 0.006129f
C551 B.n511 VSUBS 0.006129f
C552 B.n512 VSUBS 0.006129f
C553 B.n513 VSUBS 0.006129f
C554 B.n514 VSUBS 0.006129f
C555 B.n515 VSUBS 0.006129f
C556 B.n516 VSUBS 0.006129f
C557 B.n517 VSUBS 0.004236f
C558 B.n518 VSUBS 0.014201f
C559 B.n519 VSUBS 0.004958f
C560 B.n520 VSUBS 0.006129f
C561 B.n521 VSUBS 0.006129f
C562 B.n522 VSUBS 0.006129f
C563 B.n523 VSUBS 0.006129f
C564 B.n524 VSUBS 0.006129f
C565 B.n525 VSUBS 0.006129f
C566 B.n526 VSUBS 0.006129f
C567 B.n527 VSUBS 0.006129f
C568 B.n528 VSUBS 0.006129f
C569 B.n529 VSUBS 0.006129f
C570 B.n530 VSUBS 0.006129f
C571 B.n531 VSUBS 0.004958f
C572 B.n532 VSUBS 0.014201f
C573 B.n533 VSUBS 0.004236f
C574 B.n534 VSUBS 0.006129f
C575 B.n535 VSUBS 0.006129f
C576 B.n536 VSUBS 0.006129f
C577 B.n537 VSUBS 0.006129f
C578 B.n538 VSUBS 0.006129f
C579 B.n539 VSUBS 0.006129f
C580 B.n540 VSUBS 0.006129f
C581 B.n541 VSUBS 0.006129f
C582 B.n542 VSUBS 0.006129f
C583 B.n543 VSUBS 0.006129f
C584 B.n544 VSUBS 0.006129f
C585 B.n545 VSUBS 0.006129f
C586 B.n546 VSUBS 0.006129f
C587 B.n547 VSUBS 0.006129f
C588 B.n548 VSUBS 0.006129f
C589 B.n549 VSUBS 0.006129f
C590 B.n550 VSUBS 0.006129f
C591 B.n551 VSUBS 0.006129f
C592 B.n552 VSUBS 0.006129f
C593 B.n553 VSUBS 0.006129f
C594 B.n554 VSUBS 0.006129f
C595 B.n555 VSUBS 0.006129f
C596 B.n556 VSUBS 0.006129f
C597 B.n557 VSUBS 0.006129f
C598 B.n558 VSUBS 0.006129f
C599 B.n559 VSUBS 0.006129f
C600 B.n560 VSUBS 0.006129f
C601 B.n561 VSUBS 0.006129f
C602 B.n562 VSUBS 0.006129f
C603 B.n563 VSUBS 0.006129f
C604 B.n564 VSUBS 0.006129f
C605 B.n565 VSUBS 0.006129f
C606 B.n566 VSUBS 0.006129f
C607 B.n567 VSUBS 0.006129f
C608 B.n568 VSUBS 0.006129f
C609 B.n569 VSUBS 0.006129f
C610 B.n570 VSUBS 0.006129f
C611 B.n571 VSUBS 0.006129f
C612 B.n572 VSUBS 0.006129f
C613 B.n573 VSUBS 0.006129f
C614 B.n574 VSUBS 0.006129f
C615 B.n575 VSUBS 0.006129f
C616 B.n576 VSUBS 0.006129f
C617 B.n577 VSUBS 0.006129f
C618 B.n578 VSUBS 0.006129f
C619 B.n579 VSUBS 0.006129f
C620 B.n580 VSUBS 0.006129f
C621 B.n581 VSUBS 0.006129f
C622 B.n582 VSUBS 0.006129f
C623 B.n583 VSUBS 0.006129f
C624 B.n584 VSUBS 0.006129f
C625 B.n585 VSUBS 0.006129f
C626 B.n586 VSUBS 0.006129f
C627 B.n587 VSUBS 0.006129f
C628 B.n588 VSUBS 0.006129f
C629 B.n589 VSUBS 0.006129f
C630 B.n590 VSUBS 0.006129f
C631 B.n591 VSUBS 0.006129f
C632 B.n592 VSUBS 0.006129f
C633 B.n593 VSUBS 0.006129f
C634 B.n594 VSUBS 0.006129f
C635 B.n595 VSUBS 0.006129f
C636 B.n596 VSUBS 0.006129f
C637 B.n597 VSUBS 0.006129f
C638 B.n598 VSUBS 0.006129f
C639 B.n599 VSUBS 0.006129f
C640 B.n600 VSUBS 0.006129f
C641 B.n601 VSUBS 0.006129f
C642 B.n602 VSUBS 0.006129f
C643 B.n603 VSUBS 0.006129f
C644 B.n604 VSUBS 0.006129f
C645 B.n605 VSUBS 0.006129f
C646 B.n606 VSUBS 0.006129f
C647 B.n607 VSUBS 0.006129f
C648 B.n608 VSUBS 0.006129f
C649 B.n609 VSUBS 0.006129f
C650 B.n610 VSUBS 0.006129f
C651 B.n611 VSUBS 0.006129f
C652 B.n612 VSUBS 0.006129f
C653 B.n613 VSUBS 0.006129f
C654 B.n614 VSUBS 0.013792f
C655 B.n615 VSUBS 0.013792f
C656 B.n616 VSUBS 0.013069f
C657 B.n617 VSUBS 0.006129f
C658 B.n618 VSUBS 0.006129f
C659 B.n619 VSUBS 0.006129f
C660 B.n620 VSUBS 0.006129f
C661 B.n621 VSUBS 0.006129f
C662 B.n622 VSUBS 0.006129f
C663 B.n623 VSUBS 0.006129f
C664 B.n624 VSUBS 0.006129f
C665 B.n625 VSUBS 0.006129f
C666 B.n626 VSUBS 0.006129f
C667 B.n627 VSUBS 0.006129f
C668 B.n628 VSUBS 0.006129f
C669 B.n629 VSUBS 0.006129f
C670 B.n630 VSUBS 0.006129f
C671 B.n631 VSUBS 0.006129f
C672 B.n632 VSUBS 0.006129f
C673 B.n633 VSUBS 0.006129f
C674 B.n634 VSUBS 0.006129f
C675 B.n635 VSUBS 0.006129f
C676 B.n636 VSUBS 0.006129f
C677 B.n637 VSUBS 0.006129f
C678 B.n638 VSUBS 0.006129f
C679 B.n639 VSUBS 0.006129f
C680 B.n640 VSUBS 0.006129f
C681 B.n641 VSUBS 0.006129f
C682 B.n642 VSUBS 0.006129f
C683 B.n643 VSUBS 0.007999f
C684 B.n644 VSUBS 0.00852f
C685 B.n645 VSUBS 0.016944f
C686 VDD1.t1 VSUBS 2.76252f
C687 VDD1.t0 VSUBS 3.44356f
C688 VP.t0 VSUBS 4.31377f
C689 VP.t1 VSUBS 3.92988f
C690 VP.n0 VSUBS 6.40288f
C691 VDD2.t1 VSUBS 3.43835f
C692 VDD2.t0 VSUBS 2.78016f
C693 VDD2.n0 VSUBS 3.49707f
C694 VTAIL.t0 VSUBS 3.65619f
C695 VTAIL.n0 VSUBS 2.83603f
C696 VTAIL.t2 VSUBS 3.6562f
C697 VTAIL.n1 VSUBS 2.8678f
C698 VTAIL.t1 VSUBS 3.65619f
C699 VTAIL.n2 VSUBS 2.71981f
C700 VTAIL.t3 VSUBS 3.65619f
C701 VTAIL.n3 VSUBS 2.63535f
C702 VN.t0 VSUBS 3.8321f
C703 VN.t1 VSUBS 4.21105f
.ends

