* NGSPICE file created from diff_pair_sample_1630.ext - technology: sky130A

.subckt diff_pair_sample_1630 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t15 VP.t0 VDD1.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=5.0154 pd=26.5 as=2.1219 ps=13.19 w=12.86 l=1.57
X1 VDD1.t3 VP.t1 VTAIL.t14 B.t1 sky130_fd_pr__nfet_01v8 ad=2.1219 pd=13.19 as=2.1219 ps=13.19 w=12.86 l=1.57
X2 B.t21 B.t19 B.t20 B.t9 sky130_fd_pr__nfet_01v8 ad=5.0154 pd=26.5 as=0 ps=0 w=12.86 l=1.57
X3 VDD2.t7 VN.t0 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=2.1219 pd=13.19 as=2.1219 ps=13.19 w=12.86 l=1.57
X4 B.t18 B.t16 B.t17 B.t13 sky130_fd_pr__nfet_01v8 ad=5.0154 pd=26.5 as=0 ps=0 w=12.86 l=1.57
X5 B.t15 B.t12 B.t14 B.t13 sky130_fd_pr__nfet_01v8 ad=5.0154 pd=26.5 as=0 ps=0 w=12.86 l=1.57
X6 VDD1.t5 VP.t2 VTAIL.t13 B.t0 sky130_fd_pr__nfet_01v8 ad=2.1219 pd=13.19 as=2.1219 ps=13.19 w=12.86 l=1.57
X7 VTAIL.t2 VN.t1 VDD2.t6 B.t2 sky130_fd_pr__nfet_01v8 ad=5.0154 pd=26.5 as=2.1219 ps=13.19 w=12.86 l=1.57
X8 VDD2.t5 VN.t2 VTAIL.t6 B.t6 sky130_fd_pr__nfet_01v8 ad=2.1219 pd=13.19 as=5.0154 ps=26.5 w=12.86 l=1.57
X9 VTAIL.t4 VN.t3 VDD2.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=5.0154 pd=26.5 as=2.1219 ps=13.19 w=12.86 l=1.57
X10 VDD2.t3 VN.t4 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=2.1219 pd=13.19 as=2.1219 ps=13.19 w=12.86 l=1.57
X11 VTAIL.t12 VP.t3 VDD1.t7 B.t7 sky130_fd_pr__nfet_01v8 ad=2.1219 pd=13.19 as=2.1219 ps=13.19 w=12.86 l=1.57
X12 VDD2.t2 VN.t5 VTAIL.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=2.1219 pd=13.19 as=5.0154 ps=26.5 w=12.86 l=1.57
X13 VTAIL.t7 VN.t6 VDD2.t1 B.t7 sky130_fd_pr__nfet_01v8 ad=2.1219 pd=13.19 as=2.1219 ps=13.19 w=12.86 l=1.57
X14 VTAIL.t11 VP.t4 VDD1.t6 B.t2 sky130_fd_pr__nfet_01v8 ad=5.0154 pd=26.5 as=2.1219 ps=13.19 w=12.86 l=1.57
X15 VDD1.t2 VP.t5 VTAIL.t10 B.t6 sky130_fd_pr__nfet_01v8 ad=2.1219 pd=13.19 as=5.0154 ps=26.5 w=12.86 l=1.57
X16 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=5.0154 pd=26.5 as=0 ps=0 w=12.86 l=1.57
X17 VDD1.t0 VP.t6 VTAIL.t9 B.t5 sky130_fd_pr__nfet_01v8 ad=2.1219 pd=13.19 as=5.0154 ps=26.5 w=12.86 l=1.57
X18 VTAIL.t3 VN.t7 VDD2.t0 B.t3 sky130_fd_pr__nfet_01v8 ad=2.1219 pd=13.19 as=2.1219 ps=13.19 w=12.86 l=1.57
X19 VTAIL.t8 VP.t7 VDD1.t1 B.t3 sky130_fd_pr__nfet_01v8 ad=2.1219 pd=13.19 as=2.1219 ps=13.19 w=12.86 l=1.57
R0 VP.n10 VP.t0 228.359
R1 VP.n28 VP.t4 197.405
R2 VP.n35 VP.t1 197.405
R3 VP.n42 VP.t7 197.405
R4 VP.n49 VP.t6 197.405
R5 VP.n25 VP.t5 197.405
R6 VP.n18 VP.t3 197.405
R7 VP.n11 VP.t2 197.405
R8 VP.n28 VP.n27 180.974
R9 VP.n50 VP.n49 180.974
R10 VP.n26 VP.n25 180.974
R11 VP.n13 VP.n12 161.3
R12 VP.n14 VP.n9 161.3
R13 VP.n16 VP.n15 161.3
R14 VP.n17 VP.n8 161.3
R15 VP.n20 VP.n19 161.3
R16 VP.n21 VP.n7 161.3
R17 VP.n23 VP.n22 161.3
R18 VP.n24 VP.n6 161.3
R19 VP.n48 VP.n0 161.3
R20 VP.n47 VP.n46 161.3
R21 VP.n45 VP.n1 161.3
R22 VP.n44 VP.n43 161.3
R23 VP.n41 VP.n2 161.3
R24 VP.n40 VP.n39 161.3
R25 VP.n38 VP.n3 161.3
R26 VP.n37 VP.n36 161.3
R27 VP.n34 VP.n4 161.3
R28 VP.n33 VP.n32 161.3
R29 VP.n31 VP.n5 161.3
R30 VP.n30 VP.n29 161.3
R31 VP.n11 VP.n10 56.6077
R32 VP.n40 VP.n3 56.5617
R33 VP.n16 VP.n9 56.5617
R34 VP.n33 VP.n5 55.1086
R35 VP.n47 VP.n1 55.1086
R36 VP.n23 VP.n7 55.1086
R37 VP.n27 VP.n26 46.5914
R38 VP.n34 VP.n33 26.0455
R39 VP.n43 VP.n1 26.0455
R40 VP.n19 VP.n7 26.0455
R41 VP.n29 VP.n5 24.5923
R42 VP.n36 VP.n3 24.5923
R43 VP.n41 VP.n40 24.5923
R44 VP.n48 VP.n47 24.5923
R45 VP.n24 VP.n23 24.5923
R46 VP.n17 VP.n16 24.5923
R47 VP.n12 VP.n9 24.5923
R48 VP.n13 VP.n10 18.2882
R49 VP.n35 VP.n34 14.7556
R50 VP.n43 VP.n42 14.7556
R51 VP.n19 VP.n18 14.7556
R52 VP.n36 VP.n35 9.83723
R53 VP.n42 VP.n41 9.83723
R54 VP.n18 VP.n17 9.83723
R55 VP.n12 VP.n11 9.83723
R56 VP.n29 VP.n28 4.91887
R57 VP.n49 VP.n48 4.91887
R58 VP.n25 VP.n24 4.91887
R59 VP.n14 VP.n13 0.189894
R60 VP.n15 VP.n14 0.189894
R61 VP.n15 VP.n8 0.189894
R62 VP.n20 VP.n8 0.189894
R63 VP.n21 VP.n20 0.189894
R64 VP.n22 VP.n21 0.189894
R65 VP.n22 VP.n6 0.189894
R66 VP.n26 VP.n6 0.189894
R67 VP.n30 VP.n27 0.189894
R68 VP.n31 VP.n30 0.189894
R69 VP.n32 VP.n31 0.189894
R70 VP.n32 VP.n4 0.189894
R71 VP.n37 VP.n4 0.189894
R72 VP.n38 VP.n37 0.189894
R73 VP.n39 VP.n38 0.189894
R74 VP.n39 VP.n2 0.189894
R75 VP.n44 VP.n2 0.189894
R76 VP.n45 VP.n44 0.189894
R77 VP.n46 VP.n45 0.189894
R78 VP.n46 VP.n0 0.189894
R79 VP.n50 VP.n0 0.189894
R80 VP VP.n50 0.0516364
R81 VDD1 VDD1.n0 62.9683
R82 VDD1.n3 VDD1.n2 62.8548
R83 VDD1.n3 VDD1.n1 62.8548
R84 VDD1.n5 VDD1.n4 62.091
R85 VDD1.n5 VDD1.n3 42.7552
R86 VDD1.n4 VDD1.t7 1.54016
R87 VDD1.n4 VDD1.t2 1.54016
R88 VDD1.n0 VDD1.t4 1.54016
R89 VDD1.n0 VDD1.t5 1.54016
R90 VDD1.n2 VDD1.t1 1.54016
R91 VDD1.n2 VDD1.t0 1.54016
R92 VDD1.n1 VDD1.t6 1.54016
R93 VDD1.n1 VDD1.t3 1.54016
R94 VDD1 VDD1.n5 0.761276
R95 VTAIL.n562 VTAIL.n498 289.615
R96 VTAIL.n66 VTAIL.n2 289.615
R97 VTAIL.n136 VTAIL.n72 289.615
R98 VTAIL.n208 VTAIL.n144 289.615
R99 VTAIL.n492 VTAIL.n428 289.615
R100 VTAIL.n420 VTAIL.n356 289.615
R101 VTAIL.n350 VTAIL.n286 289.615
R102 VTAIL.n278 VTAIL.n214 289.615
R103 VTAIL.n521 VTAIL.n520 185
R104 VTAIL.n518 VTAIL.n517 185
R105 VTAIL.n527 VTAIL.n526 185
R106 VTAIL.n529 VTAIL.n528 185
R107 VTAIL.n514 VTAIL.n513 185
R108 VTAIL.n535 VTAIL.n534 185
R109 VTAIL.n538 VTAIL.n537 185
R110 VTAIL.n536 VTAIL.n510 185
R111 VTAIL.n543 VTAIL.n509 185
R112 VTAIL.n545 VTAIL.n544 185
R113 VTAIL.n547 VTAIL.n546 185
R114 VTAIL.n506 VTAIL.n505 185
R115 VTAIL.n553 VTAIL.n552 185
R116 VTAIL.n555 VTAIL.n554 185
R117 VTAIL.n502 VTAIL.n501 185
R118 VTAIL.n561 VTAIL.n560 185
R119 VTAIL.n563 VTAIL.n562 185
R120 VTAIL.n25 VTAIL.n24 185
R121 VTAIL.n22 VTAIL.n21 185
R122 VTAIL.n31 VTAIL.n30 185
R123 VTAIL.n33 VTAIL.n32 185
R124 VTAIL.n18 VTAIL.n17 185
R125 VTAIL.n39 VTAIL.n38 185
R126 VTAIL.n42 VTAIL.n41 185
R127 VTAIL.n40 VTAIL.n14 185
R128 VTAIL.n47 VTAIL.n13 185
R129 VTAIL.n49 VTAIL.n48 185
R130 VTAIL.n51 VTAIL.n50 185
R131 VTAIL.n10 VTAIL.n9 185
R132 VTAIL.n57 VTAIL.n56 185
R133 VTAIL.n59 VTAIL.n58 185
R134 VTAIL.n6 VTAIL.n5 185
R135 VTAIL.n65 VTAIL.n64 185
R136 VTAIL.n67 VTAIL.n66 185
R137 VTAIL.n95 VTAIL.n94 185
R138 VTAIL.n92 VTAIL.n91 185
R139 VTAIL.n101 VTAIL.n100 185
R140 VTAIL.n103 VTAIL.n102 185
R141 VTAIL.n88 VTAIL.n87 185
R142 VTAIL.n109 VTAIL.n108 185
R143 VTAIL.n112 VTAIL.n111 185
R144 VTAIL.n110 VTAIL.n84 185
R145 VTAIL.n117 VTAIL.n83 185
R146 VTAIL.n119 VTAIL.n118 185
R147 VTAIL.n121 VTAIL.n120 185
R148 VTAIL.n80 VTAIL.n79 185
R149 VTAIL.n127 VTAIL.n126 185
R150 VTAIL.n129 VTAIL.n128 185
R151 VTAIL.n76 VTAIL.n75 185
R152 VTAIL.n135 VTAIL.n134 185
R153 VTAIL.n137 VTAIL.n136 185
R154 VTAIL.n167 VTAIL.n166 185
R155 VTAIL.n164 VTAIL.n163 185
R156 VTAIL.n173 VTAIL.n172 185
R157 VTAIL.n175 VTAIL.n174 185
R158 VTAIL.n160 VTAIL.n159 185
R159 VTAIL.n181 VTAIL.n180 185
R160 VTAIL.n184 VTAIL.n183 185
R161 VTAIL.n182 VTAIL.n156 185
R162 VTAIL.n189 VTAIL.n155 185
R163 VTAIL.n191 VTAIL.n190 185
R164 VTAIL.n193 VTAIL.n192 185
R165 VTAIL.n152 VTAIL.n151 185
R166 VTAIL.n199 VTAIL.n198 185
R167 VTAIL.n201 VTAIL.n200 185
R168 VTAIL.n148 VTAIL.n147 185
R169 VTAIL.n207 VTAIL.n206 185
R170 VTAIL.n209 VTAIL.n208 185
R171 VTAIL.n493 VTAIL.n492 185
R172 VTAIL.n491 VTAIL.n490 185
R173 VTAIL.n432 VTAIL.n431 185
R174 VTAIL.n485 VTAIL.n484 185
R175 VTAIL.n483 VTAIL.n482 185
R176 VTAIL.n436 VTAIL.n435 185
R177 VTAIL.n477 VTAIL.n476 185
R178 VTAIL.n475 VTAIL.n474 185
R179 VTAIL.n473 VTAIL.n439 185
R180 VTAIL.n443 VTAIL.n440 185
R181 VTAIL.n468 VTAIL.n467 185
R182 VTAIL.n466 VTAIL.n465 185
R183 VTAIL.n445 VTAIL.n444 185
R184 VTAIL.n460 VTAIL.n459 185
R185 VTAIL.n458 VTAIL.n457 185
R186 VTAIL.n449 VTAIL.n448 185
R187 VTAIL.n452 VTAIL.n451 185
R188 VTAIL.n421 VTAIL.n420 185
R189 VTAIL.n419 VTAIL.n418 185
R190 VTAIL.n360 VTAIL.n359 185
R191 VTAIL.n413 VTAIL.n412 185
R192 VTAIL.n411 VTAIL.n410 185
R193 VTAIL.n364 VTAIL.n363 185
R194 VTAIL.n405 VTAIL.n404 185
R195 VTAIL.n403 VTAIL.n402 185
R196 VTAIL.n401 VTAIL.n367 185
R197 VTAIL.n371 VTAIL.n368 185
R198 VTAIL.n396 VTAIL.n395 185
R199 VTAIL.n394 VTAIL.n393 185
R200 VTAIL.n373 VTAIL.n372 185
R201 VTAIL.n388 VTAIL.n387 185
R202 VTAIL.n386 VTAIL.n385 185
R203 VTAIL.n377 VTAIL.n376 185
R204 VTAIL.n380 VTAIL.n379 185
R205 VTAIL.n351 VTAIL.n350 185
R206 VTAIL.n349 VTAIL.n348 185
R207 VTAIL.n290 VTAIL.n289 185
R208 VTAIL.n343 VTAIL.n342 185
R209 VTAIL.n341 VTAIL.n340 185
R210 VTAIL.n294 VTAIL.n293 185
R211 VTAIL.n335 VTAIL.n334 185
R212 VTAIL.n333 VTAIL.n332 185
R213 VTAIL.n331 VTAIL.n297 185
R214 VTAIL.n301 VTAIL.n298 185
R215 VTAIL.n326 VTAIL.n325 185
R216 VTAIL.n324 VTAIL.n323 185
R217 VTAIL.n303 VTAIL.n302 185
R218 VTAIL.n318 VTAIL.n317 185
R219 VTAIL.n316 VTAIL.n315 185
R220 VTAIL.n307 VTAIL.n306 185
R221 VTAIL.n310 VTAIL.n309 185
R222 VTAIL.n279 VTAIL.n278 185
R223 VTAIL.n277 VTAIL.n276 185
R224 VTAIL.n218 VTAIL.n217 185
R225 VTAIL.n271 VTAIL.n270 185
R226 VTAIL.n269 VTAIL.n268 185
R227 VTAIL.n222 VTAIL.n221 185
R228 VTAIL.n263 VTAIL.n262 185
R229 VTAIL.n261 VTAIL.n260 185
R230 VTAIL.n259 VTAIL.n225 185
R231 VTAIL.n229 VTAIL.n226 185
R232 VTAIL.n254 VTAIL.n253 185
R233 VTAIL.n252 VTAIL.n251 185
R234 VTAIL.n231 VTAIL.n230 185
R235 VTAIL.n246 VTAIL.n245 185
R236 VTAIL.n244 VTAIL.n243 185
R237 VTAIL.n235 VTAIL.n234 185
R238 VTAIL.n238 VTAIL.n237 185
R239 VTAIL.t6 VTAIL.n519 149.524
R240 VTAIL.t4 VTAIL.n23 149.524
R241 VTAIL.t9 VTAIL.n93 149.524
R242 VTAIL.t11 VTAIL.n165 149.524
R243 VTAIL.t10 VTAIL.n450 149.524
R244 VTAIL.t15 VTAIL.n378 149.524
R245 VTAIL.t5 VTAIL.n308 149.524
R246 VTAIL.t2 VTAIL.n236 149.524
R247 VTAIL.n520 VTAIL.n517 104.615
R248 VTAIL.n527 VTAIL.n517 104.615
R249 VTAIL.n528 VTAIL.n527 104.615
R250 VTAIL.n528 VTAIL.n513 104.615
R251 VTAIL.n535 VTAIL.n513 104.615
R252 VTAIL.n537 VTAIL.n535 104.615
R253 VTAIL.n537 VTAIL.n536 104.615
R254 VTAIL.n536 VTAIL.n509 104.615
R255 VTAIL.n545 VTAIL.n509 104.615
R256 VTAIL.n546 VTAIL.n545 104.615
R257 VTAIL.n546 VTAIL.n505 104.615
R258 VTAIL.n553 VTAIL.n505 104.615
R259 VTAIL.n554 VTAIL.n553 104.615
R260 VTAIL.n554 VTAIL.n501 104.615
R261 VTAIL.n561 VTAIL.n501 104.615
R262 VTAIL.n562 VTAIL.n561 104.615
R263 VTAIL.n24 VTAIL.n21 104.615
R264 VTAIL.n31 VTAIL.n21 104.615
R265 VTAIL.n32 VTAIL.n31 104.615
R266 VTAIL.n32 VTAIL.n17 104.615
R267 VTAIL.n39 VTAIL.n17 104.615
R268 VTAIL.n41 VTAIL.n39 104.615
R269 VTAIL.n41 VTAIL.n40 104.615
R270 VTAIL.n40 VTAIL.n13 104.615
R271 VTAIL.n49 VTAIL.n13 104.615
R272 VTAIL.n50 VTAIL.n49 104.615
R273 VTAIL.n50 VTAIL.n9 104.615
R274 VTAIL.n57 VTAIL.n9 104.615
R275 VTAIL.n58 VTAIL.n57 104.615
R276 VTAIL.n58 VTAIL.n5 104.615
R277 VTAIL.n65 VTAIL.n5 104.615
R278 VTAIL.n66 VTAIL.n65 104.615
R279 VTAIL.n94 VTAIL.n91 104.615
R280 VTAIL.n101 VTAIL.n91 104.615
R281 VTAIL.n102 VTAIL.n101 104.615
R282 VTAIL.n102 VTAIL.n87 104.615
R283 VTAIL.n109 VTAIL.n87 104.615
R284 VTAIL.n111 VTAIL.n109 104.615
R285 VTAIL.n111 VTAIL.n110 104.615
R286 VTAIL.n110 VTAIL.n83 104.615
R287 VTAIL.n119 VTAIL.n83 104.615
R288 VTAIL.n120 VTAIL.n119 104.615
R289 VTAIL.n120 VTAIL.n79 104.615
R290 VTAIL.n127 VTAIL.n79 104.615
R291 VTAIL.n128 VTAIL.n127 104.615
R292 VTAIL.n128 VTAIL.n75 104.615
R293 VTAIL.n135 VTAIL.n75 104.615
R294 VTAIL.n136 VTAIL.n135 104.615
R295 VTAIL.n166 VTAIL.n163 104.615
R296 VTAIL.n173 VTAIL.n163 104.615
R297 VTAIL.n174 VTAIL.n173 104.615
R298 VTAIL.n174 VTAIL.n159 104.615
R299 VTAIL.n181 VTAIL.n159 104.615
R300 VTAIL.n183 VTAIL.n181 104.615
R301 VTAIL.n183 VTAIL.n182 104.615
R302 VTAIL.n182 VTAIL.n155 104.615
R303 VTAIL.n191 VTAIL.n155 104.615
R304 VTAIL.n192 VTAIL.n191 104.615
R305 VTAIL.n192 VTAIL.n151 104.615
R306 VTAIL.n199 VTAIL.n151 104.615
R307 VTAIL.n200 VTAIL.n199 104.615
R308 VTAIL.n200 VTAIL.n147 104.615
R309 VTAIL.n207 VTAIL.n147 104.615
R310 VTAIL.n208 VTAIL.n207 104.615
R311 VTAIL.n492 VTAIL.n491 104.615
R312 VTAIL.n491 VTAIL.n431 104.615
R313 VTAIL.n484 VTAIL.n431 104.615
R314 VTAIL.n484 VTAIL.n483 104.615
R315 VTAIL.n483 VTAIL.n435 104.615
R316 VTAIL.n476 VTAIL.n435 104.615
R317 VTAIL.n476 VTAIL.n475 104.615
R318 VTAIL.n475 VTAIL.n439 104.615
R319 VTAIL.n443 VTAIL.n439 104.615
R320 VTAIL.n467 VTAIL.n443 104.615
R321 VTAIL.n467 VTAIL.n466 104.615
R322 VTAIL.n466 VTAIL.n444 104.615
R323 VTAIL.n459 VTAIL.n444 104.615
R324 VTAIL.n459 VTAIL.n458 104.615
R325 VTAIL.n458 VTAIL.n448 104.615
R326 VTAIL.n451 VTAIL.n448 104.615
R327 VTAIL.n420 VTAIL.n419 104.615
R328 VTAIL.n419 VTAIL.n359 104.615
R329 VTAIL.n412 VTAIL.n359 104.615
R330 VTAIL.n412 VTAIL.n411 104.615
R331 VTAIL.n411 VTAIL.n363 104.615
R332 VTAIL.n404 VTAIL.n363 104.615
R333 VTAIL.n404 VTAIL.n403 104.615
R334 VTAIL.n403 VTAIL.n367 104.615
R335 VTAIL.n371 VTAIL.n367 104.615
R336 VTAIL.n395 VTAIL.n371 104.615
R337 VTAIL.n395 VTAIL.n394 104.615
R338 VTAIL.n394 VTAIL.n372 104.615
R339 VTAIL.n387 VTAIL.n372 104.615
R340 VTAIL.n387 VTAIL.n386 104.615
R341 VTAIL.n386 VTAIL.n376 104.615
R342 VTAIL.n379 VTAIL.n376 104.615
R343 VTAIL.n350 VTAIL.n349 104.615
R344 VTAIL.n349 VTAIL.n289 104.615
R345 VTAIL.n342 VTAIL.n289 104.615
R346 VTAIL.n342 VTAIL.n341 104.615
R347 VTAIL.n341 VTAIL.n293 104.615
R348 VTAIL.n334 VTAIL.n293 104.615
R349 VTAIL.n334 VTAIL.n333 104.615
R350 VTAIL.n333 VTAIL.n297 104.615
R351 VTAIL.n301 VTAIL.n297 104.615
R352 VTAIL.n325 VTAIL.n301 104.615
R353 VTAIL.n325 VTAIL.n324 104.615
R354 VTAIL.n324 VTAIL.n302 104.615
R355 VTAIL.n317 VTAIL.n302 104.615
R356 VTAIL.n317 VTAIL.n316 104.615
R357 VTAIL.n316 VTAIL.n306 104.615
R358 VTAIL.n309 VTAIL.n306 104.615
R359 VTAIL.n278 VTAIL.n277 104.615
R360 VTAIL.n277 VTAIL.n217 104.615
R361 VTAIL.n270 VTAIL.n217 104.615
R362 VTAIL.n270 VTAIL.n269 104.615
R363 VTAIL.n269 VTAIL.n221 104.615
R364 VTAIL.n262 VTAIL.n221 104.615
R365 VTAIL.n262 VTAIL.n261 104.615
R366 VTAIL.n261 VTAIL.n225 104.615
R367 VTAIL.n229 VTAIL.n225 104.615
R368 VTAIL.n253 VTAIL.n229 104.615
R369 VTAIL.n253 VTAIL.n252 104.615
R370 VTAIL.n252 VTAIL.n230 104.615
R371 VTAIL.n245 VTAIL.n230 104.615
R372 VTAIL.n245 VTAIL.n244 104.615
R373 VTAIL.n244 VTAIL.n234 104.615
R374 VTAIL.n237 VTAIL.n234 104.615
R375 VTAIL.n520 VTAIL.t6 52.3082
R376 VTAIL.n24 VTAIL.t4 52.3082
R377 VTAIL.n94 VTAIL.t9 52.3082
R378 VTAIL.n166 VTAIL.t11 52.3082
R379 VTAIL.n451 VTAIL.t10 52.3082
R380 VTAIL.n379 VTAIL.t15 52.3082
R381 VTAIL.n309 VTAIL.t5 52.3082
R382 VTAIL.n237 VTAIL.t2 52.3082
R383 VTAIL.n1 VTAIL.n0 45.4123
R384 VTAIL.n143 VTAIL.n142 45.4123
R385 VTAIL.n427 VTAIL.n426 45.4123
R386 VTAIL.n285 VTAIL.n284 45.4123
R387 VTAIL.n567 VTAIL.n566 32.5732
R388 VTAIL.n71 VTAIL.n70 32.5732
R389 VTAIL.n141 VTAIL.n140 32.5732
R390 VTAIL.n213 VTAIL.n212 32.5732
R391 VTAIL.n497 VTAIL.n496 32.5732
R392 VTAIL.n425 VTAIL.n424 32.5732
R393 VTAIL.n355 VTAIL.n354 32.5732
R394 VTAIL.n283 VTAIL.n282 32.5732
R395 VTAIL.n567 VTAIL.n497 25.091
R396 VTAIL.n283 VTAIL.n213 25.091
R397 VTAIL.n544 VTAIL.n543 13.1884
R398 VTAIL.n48 VTAIL.n47 13.1884
R399 VTAIL.n118 VTAIL.n117 13.1884
R400 VTAIL.n190 VTAIL.n189 13.1884
R401 VTAIL.n474 VTAIL.n473 13.1884
R402 VTAIL.n402 VTAIL.n401 13.1884
R403 VTAIL.n332 VTAIL.n331 13.1884
R404 VTAIL.n260 VTAIL.n259 13.1884
R405 VTAIL.n542 VTAIL.n510 12.8005
R406 VTAIL.n547 VTAIL.n508 12.8005
R407 VTAIL.n46 VTAIL.n14 12.8005
R408 VTAIL.n51 VTAIL.n12 12.8005
R409 VTAIL.n116 VTAIL.n84 12.8005
R410 VTAIL.n121 VTAIL.n82 12.8005
R411 VTAIL.n188 VTAIL.n156 12.8005
R412 VTAIL.n193 VTAIL.n154 12.8005
R413 VTAIL.n477 VTAIL.n438 12.8005
R414 VTAIL.n472 VTAIL.n440 12.8005
R415 VTAIL.n405 VTAIL.n366 12.8005
R416 VTAIL.n400 VTAIL.n368 12.8005
R417 VTAIL.n335 VTAIL.n296 12.8005
R418 VTAIL.n330 VTAIL.n298 12.8005
R419 VTAIL.n263 VTAIL.n224 12.8005
R420 VTAIL.n258 VTAIL.n226 12.8005
R421 VTAIL.n539 VTAIL.n538 12.0247
R422 VTAIL.n548 VTAIL.n506 12.0247
R423 VTAIL.n43 VTAIL.n42 12.0247
R424 VTAIL.n52 VTAIL.n10 12.0247
R425 VTAIL.n113 VTAIL.n112 12.0247
R426 VTAIL.n122 VTAIL.n80 12.0247
R427 VTAIL.n185 VTAIL.n184 12.0247
R428 VTAIL.n194 VTAIL.n152 12.0247
R429 VTAIL.n478 VTAIL.n436 12.0247
R430 VTAIL.n469 VTAIL.n468 12.0247
R431 VTAIL.n406 VTAIL.n364 12.0247
R432 VTAIL.n397 VTAIL.n396 12.0247
R433 VTAIL.n336 VTAIL.n294 12.0247
R434 VTAIL.n327 VTAIL.n326 12.0247
R435 VTAIL.n264 VTAIL.n222 12.0247
R436 VTAIL.n255 VTAIL.n254 12.0247
R437 VTAIL.n534 VTAIL.n512 11.249
R438 VTAIL.n552 VTAIL.n551 11.249
R439 VTAIL.n38 VTAIL.n16 11.249
R440 VTAIL.n56 VTAIL.n55 11.249
R441 VTAIL.n108 VTAIL.n86 11.249
R442 VTAIL.n126 VTAIL.n125 11.249
R443 VTAIL.n180 VTAIL.n158 11.249
R444 VTAIL.n198 VTAIL.n197 11.249
R445 VTAIL.n482 VTAIL.n481 11.249
R446 VTAIL.n465 VTAIL.n442 11.249
R447 VTAIL.n410 VTAIL.n409 11.249
R448 VTAIL.n393 VTAIL.n370 11.249
R449 VTAIL.n340 VTAIL.n339 11.249
R450 VTAIL.n323 VTAIL.n300 11.249
R451 VTAIL.n268 VTAIL.n267 11.249
R452 VTAIL.n251 VTAIL.n228 11.249
R453 VTAIL.n533 VTAIL.n514 10.4732
R454 VTAIL.n555 VTAIL.n504 10.4732
R455 VTAIL.n37 VTAIL.n18 10.4732
R456 VTAIL.n59 VTAIL.n8 10.4732
R457 VTAIL.n107 VTAIL.n88 10.4732
R458 VTAIL.n129 VTAIL.n78 10.4732
R459 VTAIL.n179 VTAIL.n160 10.4732
R460 VTAIL.n201 VTAIL.n150 10.4732
R461 VTAIL.n485 VTAIL.n434 10.4732
R462 VTAIL.n464 VTAIL.n445 10.4732
R463 VTAIL.n413 VTAIL.n362 10.4732
R464 VTAIL.n392 VTAIL.n373 10.4732
R465 VTAIL.n343 VTAIL.n292 10.4732
R466 VTAIL.n322 VTAIL.n303 10.4732
R467 VTAIL.n271 VTAIL.n220 10.4732
R468 VTAIL.n250 VTAIL.n231 10.4732
R469 VTAIL.n521 VTAIL.n519 10.2747
R470 VTAIL.n25 VTAIL.n23 10.2747
R471 VTAIL.n95 VTAIL.n93 10.2747
R472 VTAIL.n167 VTAIL.n165 10.2747
R473 VTAIL.n452 VTAIL.n450 10.2747
R474 VTAIL.n380 VTAIL.n378 10.2747
R475 VTAIL.n310 VTAIL.n308 10.2747
R476 VTAIL.n238 VTAIL.n236 10.2747
R477 VTAIL.n530 VTAIL.n529 9.69747
R478 VTAIL.n556 VTAIL.n502 9.69747
R479 VTAIL.n34 VTAIL.n33 9.69747
R480 VTAIL.n60 VTAIL.n6 9.69747
R481 VTAIL.n104 VTAIL.n103 9.69747
R482 VTAIL.n130 VTAIL.n76 9.69747
R483 VTAIL.n176 VTAIL.n175 9.69747
R484 VTAIL.n202 VTAIL.n148 9.69747
R485 VTAIL.n486 VTAIL.n432 9.69747
R486 VTAIL.n461 VTAIL.n460 9.69747
R487 VTAIL.n414 VTAIL.n360 9.69747
R488 VTAIL.n389 VTAIL.n388 9.69747
R489 VTAIL.n344 VTAIL.n290 9.69747
R490 VTAIL.n319 VTAIL.n318 9.69747
R491 VTAIL.n272 VTAIL.n218 9.69747
R492 VTAIL.n247 VTAIL.n246 9.69747
R493 VTAIL.n566 VTAIL.n565 9.45567
R494 VTAIL.n70 VTAIL.n69 9.45567
R495 VTAIL.n140 VTAIL.n139 9.45567
R496 VTAIL.n212 VTAIL.n211 9.45567
R497 VTAIL.n496 VTAIL.n495 9.45567
R498 VTAIL.n424 VTAIL.n423 9.45567
R499 VTAIL.n354 VTAIL.n353 9.45567
R500 VTAIL.n282 VTAIL.n281 9.45567
R501 VTAIL.n500 VTAIL.n499 9.3005
R502 VTAIL.n559 VTAIL.n558 9.3005
R503 VTAIL.n557 VTAIL.n556 9.3005
R504 VTAIL.n504 VTAIL.n503 9.3005
R505 VTAIL.n551 VTAIL.n550 9.3005
R506 VTAIL.n549 VTAIL.n548 9.3005
R507 VTAIL.n508 VTAIL.n507 9.3005
R508 VTAIL.n523 VTAIL.n522 9.3005
R509 VTAIL.n525 VTAIL.n524 9.3005
R510 VTAIL.n516 VTAIL.n515 9.3005
R511 VTAIL.n531 VTAIL.n530 9.3005
R512 VTAIL.n533 VTAIL.n532 9.3005
R513 VTAIL.n512 VTAIL.n511 9.3005
R514 VTAIL.n540 VTAIL.n539 9.3005
R515 VTAIL.n542 VTAIL.n541 9.3005
R516 VTAIL.n565 VTAIL.n564 9.3005
R517 VTAIL.n4 VTAIL.n3 9.3005
R518 VTAIL.n63 VTAIL.n62 9.3005
R519 VTAIL.n61 VTAIL.n60 9.3005
R520 VTAIL.n8 VTAIL.n7 9.3005
R521 VTAIL.n55 VTAIL.n54 9.3005
R522 VTAIL.n53 VTAIL.n52 9.3005
R523 VTAIL.n12 VTAIL.n11 9.3005
R524 VTAIL.n27 VTAIL.n26 9.3005
R525 VTAIL.n29 VTAIL.n28 9.3005
R526 VTAIL.n20 VTAIL.n19 9.3005
R527 VTAIL.n35 VTAIL.n34 9.3005
R528 VTAIL.n37 VTAIL.n36 9.3005
R529 VTAIL.n16 VTAIL.n15 9.3005
R530 VTAIL.n44 VTAIL.n43 9.3005
R531 VTAIL.n46 VTAIL.n45 9.3005
R532 VTAIL.n69 VTAIL.n68 9.3005
R533 VTAIL.n74 VTAIL.n73 9.3005
R534 VTAIL.n133 VTAIL.n132 9.3005
R535 VTAIL.n131 VTAIL.n130 9.3005
R536 VTAIL.n78 VTAIL.n77 9.3005
R537 VTAIL.n125 VTAIL.n124 9.3005
R538 VTAIL.n123 VTAIL.n122 9.3005
R539 VTAIL.n82 VTAIL.n81 9.3005
R540 VTAIL.n97 VTAIL.n96 9.3005
R541 VTAIL.n99 VTAIL.n98 9.3005
R542 VTAIL.n90 VTAIL.n89 9.3005
R543 VTAIL.n105 VTAIL.n104 9.3005
R544 VTAIL.n107 VTAIL.n106 9.3005
R545 VTAIL.n86 VTAIL.n85 9.3005
R546 VTAIL.n114 VTAIL.n113 9.3005
R547 VTAIL.n116 VTAIL.n115 9.3005
R548 VTAIL.n139 VTAIL.n138 9.3005
R549 VTAIL.n146 VTAIL.n145 9.3005
R550 VTAIL.n205 VTAIL.n204 9.3005
R551 VTAIL.n203 VTAIL.n202 9.3005
R552 VTAIL.n150 VTAIL.n149 9.3005
R553 VTAIL.n197 VTAIL.n196 9.3005
R554 VTAIL.n195 VTAIL.n194 9.3005
R555 VTAIL.n154 VTAIL.n153 9.3005
R556 VTAIL.n169 VTAIL.n168 9.3005
R557 VTAIL.n171 VTAIL.n170 9.3005
R558 VTAIL.n162 VTAIL.n161 9.3005
R559 VTAIL.n177 VTAIL.n176 9.3005
R560 VTAIL.n179 VTAIL.n178 9.3005
R561 VTAIL.n158 VTAIL.n157 9.3005
R562 VTAIL.n186 VTAIL.n185 9.3005
R563 VTAIL.n188 VTAIL.n187 9.3005
R564 VTAIL.n211 VTAIL.n210 9.3005
R565 VTAIL.n454 VTAIL.n453 9.3005
R566 VTAIL.n456 VTAIL.n455 9.3005
R567 VTAIL.n447 VTAIL.n446 9.3005
R568 VTAIL.n462 VTAIL.n461 9.3005
R569 VTAIL.n464 VTAIL.n463 9.3005
R570 VTAIL.n442 VTAIL.n441 9.3005
R571 VTAIL.n470 VTAIL.n469 9.3005
R572 VTAIL.n472 VTAIL.n471 9.3005
R573 VTAIL.n495 VTAIL.n494 9.3005
R574 VTAIL.n430 VTAIL.n429 9.3005
R575 VTAIL.n489 VTAIL.n488 9.3005
R576 VTAIL.n487 VTAIL.n486 9.3005
R577 VTAIL.n434 VTAIL.n433 9.3005
R578 VTAIL.n481 VTAIL.n480 9.3005
R579 VTAIL.n479 VTAIL.n478 9.3005
R580 VTAIL.n438 VTAIL.n437 9.3005
R581 VTAIL.n382 VTAIL.n381 9.3005
R582 VTAIL.n384 VTAIL.n383 9.3005
R583 VTAIL.n375 VTAIL.n374 9.3005
R584 VTAIL.n390 VTAIL.n389 9.3005
R585 VTAIL.n392 VTAIL.n391 9.3005
R586 VTAIL.n370 VTAIL.n369 9.3005
R587 VTAIL.n398 VTAIL.n397 9.3005
R588 VTAIL.n400 VTAIL.n399 9.3005
R589 VTAIL.n423 VTAIL.n422 9.3005
R590 VTAIL.n358 VTAIL.n357 9.3005
R591 VTAIL.n417 VTAIL.n416 9.3005
R592 VTAIL.n415 VTAIL.n414 9.3005
R593 VTAIL.n362 VTAIL.n361 9.3005
R594 VTAIL.n409 VTAIL.n408 9.3005
R595 VTAIL.n407 VTAIL.n406 9.3005
R596 VTAIL.n366 VTAIL.n365 9.3005
R597 VTAIL.n312 VTAIL.n311 9.3005
R598 VTAIL.n314 VTAIL.n313 9.3005
R599 VTAIL.n305 VTAIL.n304 9.3005
R600 VTAIL.n320 VTAIL.n319 9.3005
R601 VTAIL.n322 VTAIL.n321 9.3005
R602 VTAIL.n300 VTAIL.n299 9.3005
R603 VTAIL.n328 VTAIL.n327 9.3005
R604 VTAIL.n330 VTAIL.n329 9.3005
R605 VTAIL.n353 VTAIL.n352 9.3005
R606 VTAIL.n288 VTAIL.n287 9.3005
R607 VTAIL.n347 VTAIL.n346 9.3005
R608 VTAIL.n345 VTAIL.n344 9.3005
R609 VTAIL.n292 VTAIL.n291 9.3005
R610 VTAIL.n339 VTAIL.n338 9.3005
R611 VTAIL.n337 VTAIL.n336 9.3005
R612 VTAIL.n296 VTAIL.n295 9.3005
R613 VTAIL.n240 VTAIL.n239 9.3005
R614 VTAIL.n242 VTAIL.n241 9.3005
R615 VTAIL.n233 VTAIL.n232 9.3005
R616 VTAIL.n248 VTAIL.n247 9.3005
R617 VTAIL.n250 VTAIL.n249 9.3005
R618 VTAIL.n228 VTAIL.n227 9.3005
R619 VTAIL.n256 VTAIL.n255 9.3005
R620 VTAIL.n258 VTAIL.n257 9.3005
R621 VTAIL.n281 VTAIL.n280 9.3005
R622 VTAIL.n216 VTAIL.n215 9.3005
R623 VTAIL.n275 VTAIL.n274 9.3005
R624 VTAIL.n273 VTAIL.n272 9.3005
R625 VTAIL.n220 VTAIL.n219 9.3005
R626 VTAIL.n267 VTAIL.n266 9.3005
R627 VTAIL.n265 VTAIL.n264 9.3005
R628 VTAIL.n224 VTAIL.n223 9.3005
R629 VTAIL.n526 VTAIL.n516 8.92171
R630 VTAIL.n560 VTAIL.n559 8.92171
R631 VTAIL.n30 VTAIL.n20 8.92171
R632 VTAIL.n64 VTAIL.n63 8.92171
R633 VTAIL.n100 VTAIL.n90 8.92171
R634 VTAIL.n134 VTAIL.n133 8.92171
R635 VTAIL.n172 VTAIL.n162 8.92171
R636 VTAIL.n206 VTAIL.n205 8.92171
R637 VTAIL.n490 VTAIL.n489 8.92171
R638 VTAIL.n457 VTAIL.n447 8.92171
R639 VTAIL.n418 VTAIL.n417 8.92171
R640 VTAIL.n385 VTAIL.n375 8.92171
R641 VTAIL.n348 VTAIL.n347 8.92171
R642 VTAIL.n315 VTAIL.n305 8.92171
R643 VTAIL.n276 VTAIL.n275 8.92171
R644 VTAIL.n243 VTAIL.n233 8.92171
R645 VTAIL.n525 VTAIL.n518 8.14595
R646 VTAIL.n563 VTAIL.n500 8.14595
R647 VTAIL.n29 VTAIL.n22 8.14595
R648 VTAIL.n67 VTAIL.n4 8.14595
R649 VTAIL.n99 VTAIL.n92 8.14595
R650 VTAIL.n137 VTAIL.n74 8.14595
R651 VTAIL.n171 VTAIL.n164 8.14595
R652 VTAIL.n209 VTAIL.n146 8.14595
R653 VTAIL.n493 VTAIL.n430 8.14595
R654 VTAIL.n456 VTAIL.n449 8.14595
R655 VTAIL.n421 VTAIL.n358 8.14595
R656 VTAIL.n384 VTAIL.n377 8.14595
R657 VTAIL.n351 VTAIL.n288 8.14595
R658 VTAIL.n314 VTAIL.n307 8.14595
R659 VTAIL.n279 VTAIL.n216 8.14595
R660 VTAIL.n242 VTAIL.n235 8.14595
R661 VTAIL.n522 VTAIL.n521 7.3702
R662 VTAIL.n564 VTAIL.n498 7.3702
R663 VTAIL.n26 VTAIL.n25 7.3702
R664 VTAIL.n68 VTAIL.n2 7.3702
R665 VTAIL.n96 VTAIL.n95 7.3702
R666 VTAIL.n138 VTAIL.n72 7.3702
R667 VTAIL.n168 VTAIL.n167 7.3702
R668 VTAIL.n210 VTAIL.n144 7.3702
R669 VTAIL.n494 VTAIL.n428 7.3702
R670 VTAIL.n453 VTAIL.n452 7.3702
R671 VTAIL.n422 VTAIL.n356 7.3702
R672 VTAIL.n381 VTAIL.n380 7.3702
R673 VTAIL.n352 VTAIL.n286 7.3702
R674 VTAIL.n311 VTAIL.n310 7.3702
R675 VTAIL.n280 VTAIL.n214 7.3702
R676 VTAIL.n239 VTAIL.n238 7.3702
R677 VTAIL.n566 VTAIL.n498 6.59444
R678 VTAIL.n70 VTAIL.n2 6.59444
R679 VTAIL.n140 VTAIL.n72 6.59444
R680 VTAIL.n212 VTAIL.n144 6.59444
R681 VTAIL.n496 VTAIL.n428 6.59444
R682 VTAIL.n424 VTAIL.n356 6.59444
R683 VTAIL.n354 VTAIL.n286 6.59444
R684 VTAIL.n282 VTAIL.n214 6.59444
R685 VTAIL.n522 VTAIL.n518 5.81868
R686 VTAIL.n564 VTAIL.n563 5.81868
R687 VTAIL.n26 VTAIL.n22 5.81868
R688 VTAIL.n68 VTAIL.n67 5.81868
R689 VTAIL.n96 VTAIL.n92 5.81868
R690 VTAIL.n138 VTAIL.n137 5.81868
R691 VTAIL.n168 VTAIL.n164 5.81868
R692 VTAIL.n210 VTAIL.n209 5.81868
R693 VTAIL.n494 VTAIL.n493 5.81868
R694 VTAIL.n453 VTAIL.n449 5.81868
R695 VTAIL.n422 VTAIL.n421 5.81868
R696 VTAIL.n381 VTAIL.n377 5.81868
R697 VTAIL.n352 VTAIL.n351 5.81868
R698 VTAIL.n311 VTAIL.n307 5.81868
R699 VTAIL.n280 VTAIL.n279 5.81868
R700 VTAIL.n239 VTAIL.n235 5.81868
R701 VTAIL.n526 VTAIL.n525 5.04292
R702 VTAIL.n560 VTAIL.n500 5.04292
R703 VTAIL.n30 VTAIL.n29 5.04292
R704 VTAIL.n64 VTAIL.n4 5.04292
R705 VTAIL.n100 VTAIL.n99 5.04292
R706 VTAIL.n134 VTAIL.n74 5.04292
R707 VTAIL.n172 VTAIL.n171 5.04292
R708 VTAIL.n206 VTAIL.n146 5.04292
R709 VTAIL.n490 VTAIL.n430 5.04292
R710 VTAIL.n457 VTAIL.n456 5.04292
R711 VTAIL.n418 VTAIL.n358 5.04292
R712 VTAIL.n385 VTAIL.n384 5.04292
R713 VTAIL.n348 VTAIL.n288 5.04292
R714 VTAIL.n315 VTAIL.n314 5.04292
R715 VTAIL.n276 VTAIL.n216 5.04292
R716 VTAIL.n243 VTAIL.n242 5.04292
R717 VTAIL.n529 VTAIL.n516 4.26717
R718 VTAIL.n559 VTAIL.n502 4.26717
R719 VTAIL.n33 VTAIL.n20 4.26717
R720 VTAIL.n63 VTAIL.n6 4.26717
R721 VTAIL.n103 VTAIL.n90 4.26717
R722 VTAIL.n133 VTAIL.n76 4.26717
R723 VTAIL.n175 VTAIL.n162 4.26717
R724 VTAIL.n205 VTAIL.n148 4.26717
R725 VTAIL.n489 VTAIL.n432 4.26717
R726 VTAIL.n460 VTAIL.n447 4.26717
R727 VTAIL.n417 VTAIL.n360 4.26717
R728 VTAIL.n388 VTAIL.n375 4.26717
R729 VTAIL.n347 VTAIL.n290 4.26717
R730 VTAIL.n318 VTAIL.n305 4.26717
R731 VTAIL.n275 VTAIL.n218 4.26717
R732 VTAIL.n246 VTAIL.n233 4.26717
R733 VTAIL.n530 VTAIL.n514 3.49141
R734 VTAIL.n556 VTAIL.n555 3.49141
R735 VTAIL.n34 VTAIL.n18 3.49141
R736 VTAIL.n60 VTAIL.n59 3.49141
R737 VTAIL.n104 VTAIL.n88 3.49141
R738 VTAIL.n130 VTAIL.n129 3.49141
R739 VTAIL.n176 VTAIL.n160 3.49141
R740 VTAIL.n202 VTAIL.n201 3.49141
R741 VTAIL.n486 VTAIL.n485 3.49141
R742 VTAIL.n461 VTAIL.n445 3.49141
R743 VTAIL.n414 VTAIL.n413 3.49141
R744 VTAIL.n389 VTAIL.n373 3.49141
R745 VTAIL.n344 VTAIL.n343 3.49141
R746 VTAIL.n319 VTAIL.n303 3.49141
R747 VTAIL.n272 VTAIL.n271 3.49141
R748 VTAIL.n247 VTAIL.n231 3.49141
R749 VTAIL.n523 VTAIL.n519 2.84303
R750 VTAIL.n27 VTAIL.n23 2.84303
R751 VTAIL.n97 VTAIL.n93 2.84303
R752 VTAIL.n169 VTAIL.n165 2.84303
R753 VTAIL.n454 VTAIL.n450 2.84303
R754 VTAIL.n382 VTAIL.n378 2.84303
R755 VTAIL.n312 VTAIL.n308 2.84303
R756 VTAIL.n240 VTAIL.n236 2.84303
R757 VTAIL.n534 VTAIL.n533 2.71565
R758 VTAIL.n552 VTAIL.n504 2.71565
R759 VTAIL.n38 VTAIL.n37 2.71565
R760 VTAIL.n56 VTAIL.n8 2.71565
R761 VTAIL.n108 VTAIL.n107 2.71565
R762 VTAIL.n126 VTAIL.n78 2.71565
R763 VTAIL.n180 VTAIL.n179 2.71565
R764 VTAIL.n198 VTAIL.n150 2.71565
R765 VTAIL.n482 VTAIL.n434 2.71565
R766 VTAIL.n465 VTAIL.n464 2.71565
R767 VTAIL.n410 VTAIL.n362 2.71565
R768 VTAIL.n393 VTAIL.n392 2.71565
R769 VTAIL.n340 VTAIL.n292 2.71565
R770 VTAIL.n323 VTAIL.n322 2.71565
R771 VTAIL.n268 VTAIL.n220 2.71565
R772 VTAIL.n251 VTAIL.n250 2.71565
R773 VTAIL.n538 VTAIL.n512 1.93989
R774 VTAIL.n551 VTAIL.n506 1.93989
R775 VTAIL.n42 VTAIL.n16 1.93989
R776 VTAIL.n55 VTAIL.n10 1.93989
R777 VTAIL.n112 VTAIL.n86 1.93989
R778 VTAIL.n125 VTAIL.n80 1.93989
R779 VTAIL.n184 VTAIL.n158 1.93989
R780 VTAIL.n197 VTAIL.n152 1.93989
R781 VTAIL.n481 VTAIL.n436 1.93989
R782 VTAIL.n468 VTAIL.n442 1.93989
R783 VTAIL.n409 VTAIL.n364 1.93989
R784 VTAIL.n396 VTAIL.n370 1.93989
R785 VTAIL.n339 VTAIL.n294 1.93989
R786 VTAIL.n326 VTAIL.n300 1.93989
R787 VTAIL.n267 VTAIL.n222 1.93989
R788 VTAIL.n254 VTAIL.n228 1.93989
R789 VTAIL.n285 VTAIL.n283 1.63843
R790 VTAIL.n355 VTAIL.n285 1.63843
R791 VTAIL.n427 VTAIL.n425 1.63843
R792 VTAIL.n497 VTAIL.n427 1.63843
R793 VTAIL.n213 VTAIL.n143 1.63843
R794 VTAIL.n143 VTAIL.n141 1.63843
R795 VTAIL.n71 VTAIL.n1 1.63843
R796 VTAIL VTAIL.n567 1.58024
R797 VTAIL.n0 VTAIL.t0 1.54016
R798 VTAIL.n0 VTAIL.t7 1.54016
R799 VTAIL.n142 VTAIL.t14 1.54016
R800 VTAIL.n142 VTAIL.t8 1.54016
R801 VTAIL.n426 VTAIL.t13 1.54016
R802 VTAIL.n426 VTAIL.t12 1.54016
R803 VTAIL.n284 VTAIL.t1 1.54016
R804 VTAIL.n284 VTAIL.t3 1.54016
R805 VTAIL.n539 VTAIL.n510 1.16414
R806 VTAIL.n548 VTAIL.n547 1.16414
R807 VTAIL.n43 VTAIL.n14 1.16414
R808 VTAIL.n52 VTAIL.n51 1.16414
R809 VTAIL.n113 VTAIL.n84 1.16414
R810 VTAIL.n122 VTAIL.n121 1.16414
R811 VTAIL.n185 VTAIL.n156 1.16414
R812 VTAIL.n194 VTAIL.n193 1.16414
R813 VTAIL.n478 VTAIL.n477 1.16414
R814 VTAIL.n469 VTAIL.n440 1.16414
R815 VTAIL.n406 VTAIL.n405 1.16414
R816 VTAIL.n397 VTAIL.n368 1.16414
R817 VTAIL.n336 VTAIL.n335 1.16414
R818 VTAIL.n327 VTAIL.n298 1.16414
R819 VTAIL.n264 VTAIL.n263 1.16414
R820 VTAIL.n255 VTAIL.n226 1.16414
R821 VTAIL.n425 VTAIL.n355 0.470328
R822 VTAIL.n141 VTAIL.n71 0.470328
R823 VTAIL.n543 VTAIL.n542 0.388379
R824 VTAIL.n544 VTAIL.n508 0.388379
R825 VTAIL.n47 VTAIL.n46 0.388379
R826 VTAIL.n48 VTAIL.n12 0.388379
R827 VTAIL.n117 VTAIL.n116 0.388379
R828 VTAIL.n118 VTAIL.n82 0.388379
R829 VTAIL.n189 VTAIL.n188 0.388379
R830 VTAIL.n190 VTAIL.n154 0.388379
R831 VTAIL.n474 VTAIL.n438 0.388379
R832 VTAIL.n473 VTAIL.n472 0.388379
R833 VTAIL.n402 VTAIL.n366 0.388379
R834 VTAIL.n401 VTAIL.n400 0.388379
R835 VTAIL.n332 VTAIL.n296 0.388379
R836 VTAIL.n331 VTAIL.n330 0.388379
R837 VTAIL.n260 VTAIL.n224 0.388379
R838 VTAIL.n259 VTAIL.n258 0.388379
R839 VTAIL.n524 VTAIL.n523 0.155672
R840 VTAIL.n524 VTAIL.n515 0.155672
R841 VTAIL.n531 VTAIL.n515 0.155672
R842 VTAIL.n532 VTAIL.n531 0.155672
R843 VTAIL.n532 VTAIL.n511 0.155672
R844 VTAIL.n540 VTAIL.n511 0.155672
R845 VTAIL.n541 VTAIL.n540 0.155672
R846 VTAIL.n541 VTAIL.n507 0.155672
R847 VTAIL.n549 VTAIL.n507 0.155672
R848 VTAIL.n550 VTAIL.n549 0.155672
R849 VTAIL.n550 VTAIL.n503 0.155672
R850 VTAIL.n557 VTAIL.n503 0.155672
R851 VTAIL.n558 VTAIL.n557 0.155672
R852 VTAIL.n558 VTAIL.n499 0.155672
R853 VTAIL.n565 VTAIL.n499 0.155672
R854 VTAIL.n28 VTAIL.n27 0.155672
R855 VTAIL.n28 VTAIL.n19 0.155672
R856 VTAIL.n35 VTAIL.n19 0.155672
R857 VTAIL.n36 VTAIL.n35 0.155672
R858 VTAIL.n36 VTAIL.n15 0.155672
R859 VTAIL.n44 VTAIL.n15 0.155672
R860 VTAIL.n45 VTAIL.n44 0.155672
R861 VTAIL.n45 VTAIL.n11 0.155672
R862 VTAIL.n53 VTAIL.n11 0.155672
R863 VTAIL.n54 VTAIL.n53 0.155672
R864 VTAIL.n54 VTAIL.n7 0.155672
R865 VTAIL.n61 VTAIL.n7 0.155672
R866 VTAIL.n62 VTAIL.n61 0.155672
R867 VTAIL.n62 VTAIL.n3 0.155672
R868 VTAIL.n69 VTAIL.n3 0.155672
R869 VTAIL.n98 VTAIL.n97 0.155672
R870 VTAIL.n98 VTAIL.n89 0.155672
R871 VTAIL.n105 VTAIL.n89 0.155672
R872 VTAIL.n106 VTAIL.n105 0.155672
R873 VTAIL.n106 VTAIL.n85 0.155672
R874 VTAIL.n114 VTAIL.n85 0.155672
R875 VTAIL.n115 VTAIL.n114 0.155672
R876 VTAIL.n115 VTAIL.n81 0.155672
R877 VTAIL.n123 VTAIL.n81 0.155672
R878 VTAIL.n124 VTAIL.n123 0.155672
R879 VTAIL.n124 VTAIL.n77 0.155672
R880 VTAIL.n131 VTAIL.n77 0.155672
R881 VTAIL.n132 VTAIL.n131 0.155672
R882 VTAIL.n132 VTAIL.n73 0.155672
R883 VTAIL.n139 VTAIL.n73 0.155672
R884 VTAIL.n170 VTAIL.n169 0.155672
R885 VTAIL.n170 VTAIL.n161 0.155672
R886 VTAIL.n177 VTAIL.n161 0.155672
R887 VTAIL.n178 VTAIL.n177 0.155672
R888 VTAIL.n178 VTAIL.n157 0.155672
R889 VTAIL.n186 VTAIL.n157 0.155672
R890 VTAIL.n187 VTAIL.n186 0.155672
R891 VTAIL.n187 VTAIL.n153 0.155672
R892 VTAIL.n195 VTAIL.n153 0.155672
R893 VTAIL.n196 VTAIL.n195 0.155672
R894 VTAIL.n196 VTAIL.n149 0.155672
R895 VTAIL.n203 VTAIL.n149 0.155672
R896 VTAIL.n204 VTAIL.n203 0.155672
R897 VTAIL.n204 VTAIL.n145 0.155672
R898 VTAIL.n211 VTAIL.n145 0.155672
R899 VTAIL.n495 VTAIL.n429 0.155672
R900 VTAIL.n488 VTAIL.n429 0.155672
R901 VTAIL.n488 VTAIL.n487 0.155672
R902 VTAIL.n487 VTAIL.n433 0.155672
R903 VTAIL.n480 VTAIL.n433 0.155672
R904 VTAIL.n480 VTAIL.n479 0.155672
R905 VTAIL.n479 VTAIL.n437 0.155672
R906 VTAIL.n471 VTAIL.n437 0.155672
R907 VTAIL.n471 VTAIL.n470 0.155672
R908 VTAIL.n470 VTAIL.n441 0.155672
R909 VTAIL.n463 VTAIL.n441 0.155672
R910 VTAIL.n463 VTAIL.n462 0.155672
R911 VTAIL.n462 VTAIL.n446 0.155672
R912 VTAIL.n455 VTAIL.n446 0.155672
R913 VTAIL.n455 VTAIL.n454 0.155672
R914 VTAIL.n423 VTAIL.n357 0.155672
R915 VTAIL.n416 VTAIL.n357 0.155672
R916 VTAIL.n416 VTAIL.n415 0.155672
R917 VTAIL.n415 VTAIL.n361 0.155672
R918 VTAIL.n408 VTAIL.n361 0.155672
R919 VTAIL.n408 VTAIL.n407 0.155672
R920 VTAIL.n407 VTAIL.n365 0.155672
R921 VTAIL.n399 VTAIL.n365 0.155672
R922 VTAIL.n399 VTAIL.n398 0.155672
R923 VTAIL.n398 VTAIL.n369 0.155672
R924 VTAIL.n391 VTAIL.n369 0.155672
R925 VTAIL.n391 VTAIL.n390 0.155672
R926 VTAIL.n390 VTAIL.n374 0.155672
R927 VTAIL.n383 VTAIL.n374 0.155672
R928 VTAIL.n383 VTAIL.n382 0.155672
R929 VTAIL.n353 VTAIL.n287 0.155672
R930 VTAIL.n346 VTAIL.n287 0.155672
R931 VTAIL.n346 VTAIL.n345 0.155672
R932 VTAIL.n345 VTAIL.n291 0.155672
R933 VTAIL.n338 VTAIL.n291 0.155672
R934 VTAIL.n338 VTAIL.n337 0.155672
R935 VTAIL.n337 VTAIL.n295 0.155672
R936 VTAIL.n329 VTAIL.n295 0.155672
R937 VTAIL.n329 VTAIL.n328 0.155672
R938 VTAIL.n328 VTAIL.n299 0.155672
R939 VTAIL.n321 VTAIL.n299 0.155672
R940 VTAIL.n321 VTAIL.n320 0.155672
R941 VTAIL.n320 VTAIL.n304 0.155672
R942 VTAIL.n313 VTAIL.n304 0.155672
R943 VTAIL.n313 VTAIL.n312 0.155672
R944 VTAIL.n281 VTAIL.n215 0.155672
R945 VTAIL.n274 VTAIL.n215 0.155672
R946 VTAIL.n274 VTAIL.n273 0.155672
R947 VTAIL.n273 VTAIL.n219 0.155672
R948 VTAIL.n266 VTAIL.n219 0.155672
R949 VTAIL.n266 VTAIL.n265 0.155672
R950 VTAIL.n265 VTAIL.n223 0.155672
R951 VTAIL.n257 VTAIL.n223 0.155672
R952 VTAIL.n257 VTAIL.n256 0.155672
R953 VTAIL.n256 VTAIL.n227 0.155672
R954 VTAIL.n249 VTAIL.n227 0.155672
R955 VTAIL.n249 VTAIL.n248 0.155672
R956 VTAIL.n248 VTAIL.n232 0.155672
R957 VTAIL.n241 VTAIL.n232 0.155672
R958 VTAIL.n241 VTAIL.n240 0.155672
R959 VTAIL VTAIL.n1 0.0586897
R960 B.n790 B.n789 585
R961 B.n314 B.n117 585
R962 B.n313 B.n312 585
R963 B.n311 B.n310 585
R964 B.n309 B.n308 585
R965 B.n307 B.n306 585
R966 B.n305 B.n304 585
R967 B.n303 B.n302 585
R968 B.n301 B.n300 585
R969 B.n299 B.n298 585
R970 B.n297 B.n296 585
R971 B.n295 B.n294 585
R972 B.n293 B.n292 585
R973 B.n291 B.n290 585
R974 B.n289 B.n288 585
R975 B.n287 B.n286 585
R976 B.n285 B.n284 585
R977 B.n283 B.n282 585
R978 B.n281 B.n280 585
R979 B.n279 B.n278 585
R980 B.n277 B.n276 585
R981 B.n275 B.n274 585
R982 B.n273 B.n272 585
R983 B.n271 B.n270 585
R984 B.n269 B.n268 585
R985 B.n267 B.n266 585
R986 B.n265 B.n264 585
R987 B.n263 B.n262 585
R988 B.n261 B.n260 585
R989 B.n259 B.n258 585
R990 B.n257 B.n256 585
R991 B.n255 B.n254 585
R992 B.n253 B.n252 585
R993 B.n251 B.n250 585
R994 B.n249 B.n248 585
R995 B.n247 B.n246 585
R996 B.n245 B.n244 585
R997 B.n243 B.n242 585
R998 B.n241 B.n240 585
R999 B.n239 B.n238 585
R1000 B.n237 B.n236 585
R1001 B.n235 B.n234 585
R1002 B.n233 B.n232 585
R1003 B.n231 B.n230 585
R1004 B.n229 B.n228 585
R1005 B.n227 B.n226 585
R1006 B.n225 B.n224 585
R1007 B.n223 B.n222 585
R1008 B.n221 B.n220 585
R1009 B.n219 B.n218 585
R1010 B.n217 B.n216 585
R1011 B.n215 B.n214 585
R1012 B.n213 B.n212 585
R1013 B.n211 B.n210 585
R1014 B.n209 B.n208 585
R1015 B.n207 B.n206 585
R1016 B.n205 B.n204 585
R1017 B.n203 B.n202 585
R1018 B.n201 B.n200 585
R1019 B.n199 B.n198 585
R1020 B.n197 B.n196 585
R1021 B.n195 B.n194 585
R1022 B.n193 B.n192 585
R1023 B.n191 B.n190 585
R1024 B.n189 B.n188 585
R1025 B.n187 B.n186 585
R1026 B.n185 B.n184 585
R1027 B.n183 B.n182 585
R1028 B.n181 B.n180 585
R1029 B.n179 B.n178 585
R1030 B.n177 B.n176 585
R1031 B.n175 B.n174 585
R1032 B.n173 B.n172 585
R1033 B.n171 B.n170 585
R1034 B.n169 B.n168 585
R1035 B.n167 B.n166 585
R1036 B.n165 B.n164 585
R1037 B.n163 B.n162 585
R1038 B.n161 B.n160 585
R1039 B.n159 B.n158 585
R1040 B.n157 B.n156 585
R1041 B.n155 B.n154 585
R1042 B.n153 B.n152 585
R1043 B.n151 B.n150 585
R1044 B.n149 B.n148 585
R1045 B.n147 B.n146 585
R1046 B.n145 B.n144 585
R1047 B.n143 B.n142 585
R1048 B.n141 B.n140 585
R1049 B.n139 B.n138 585
R1050 B.n137 B.n136 585
R1051 B.n135 B.n134 585
R1052 B.n133 B.n132 585
R1053 B.n131 B.n130 585
R1054 B.n129 B.n128 585
R1055 B.n127 B.n126 585
R1056 B.n125 B.n124 585
R1057 B.n67 B.n66 585
R1058 B.n788 B.n68 585
R1059 B.n793 B.n68 585
R1060 B.n787 B.n786 585
R1061 B.n786 B.n64 585
R1062 B.n785 B.n63 585
R1063 B.n799 B.n63 585
R1064 B.n784 B.n62 585
R1065 B.n800 B.n62 585
R1066 B.n783 B.n61 585
R1067 B.n801 B.n61 585
R1068 B.n782 B.n781 585
R1069 B.n781 B.n57 585
R1070 B.n780 B.n56 585
R1071 B.n807 B.n56 585
R1072 B.n779 B.n55 585
R1073 B.n808 B.n55 585
R1074 B.n778 B.n54 585
R1075 B.n809 B.n54 585
R1076 B.n777 B.n776 585
R1077 B.n776 B.n50 585
R1078 B.n775 B.n49 585
R1079 B.n815 B.n49 585
R1080 B.n774 B.n48 585
R1081 B.n816 B.n48 585
R1082 B.n773 B.n47 585
R1083 B.n817 B.n47 585
R1084 B.n772 B.n771 585
R1085 B.n771 B.n43 585
R1086 B.n770 B.n42 585
R1087 B.n823 B.n42 585
R1088 B.n769 B.n41 585
R1089 B.n824 B.n41 585
R1090 B.n768 B.n40 585
R1091 B.n825 B.n40 585
R1092 B.n767 B.n766 585
R1093 B.n766 B.n36 585
R1094 B.n765 B.n35 585
R1095 B.n831 B.n35 585
R1096 B.n764 B.n34 585
R1097 B.n832 B.n34 585
R1098 B.n763 B.n33 585
R1099 B.n833 B.n33 585
R1100 B.n762 B.n761 585
R1101 B.n761 B.n29 585
R1102 B.n760 B.n28 585
R1103 B.n839 B.n28 585
R1104 B.n759 B.n27 585
R1105 B.n840 B.n27 585
R1106 B.n758 B.n26 585
R1107 B.n841 B.n26 585
R1108 B.n757 B.n756 585
R1109 B.n756 B.n22 585
R1110 B.n755 B.n21 585
R1111 B.n847 B.n21 585
R1112 B.n754 B.n20 585
R1113 B.n848 B.n20 585
R1114 B.n753 B.n19 585
R1115 B.n849 B.n19 585
R1116 B.n752 B.n751 585
R1117 B.n751 B.n15 585
R1118 B.n750 B.n14 585
R1119 B.n855 B.n14 585
R1120 B.n749 B.n13 585
R1121 B.n856 B.n13 585
R1122 B.n748 B.n12 585
R1123 B.n857 B.n12 585
R1124 B.n747 B.n746 585
R1125 B.n746 B.n8 585
R1126 B.n745 B.n7 585
R1127 B.n863 B.n7 585
R1128 B.n744 B.n6 585
R1129 B.n864 B.n6 585
R1130 B.n743 B.n5 585
R1131 B.n865 B.n5 585
R1132 B.n742 B.n741 585
R1133 B.n741 B.n4 585
R1134 B.n740 B.n315 585
R1135 B.n740 B.n739 585
R1136 B.n730 B.n316 585
R1137 B.n317 B.n316 585
R1138 B.n732 B.n731 585
R1139 B.n733 B.n732 585
R1140 B.n729 B.n321 585
R1141 B.n325 B.n321 585
R1142 B.n728 B.n727 585
R1143 B.n727 B.n726 585
R1144 B.n323 B.n322 585
R1145 B.n324 B.n323 585
R1146 B.n719 B.n718 585
R1147 B.n720 B.n719 585
R1148 B.n717 B.n330 585
R1149 B.n330 B.n329 585
R1150 B.n716 B.n715 585
R1151 B.n715 B.n714 585
R1152 B.n332 B.n331 585
R1153 B.n333 B.n332 585
R1154 B.n707 B.n706 585
R1155 B.n708 B.n707 585
R1156 B.n705 B.n338 585
R1157 B.n338 B.n337 585
R1158 B.n704 B.n703 585
R1159 B.n703 B.n702 585
R1160 B.n340 B.n339 585
R1161 B.n341 B.n340 585
R1162 B.n695 B.n694 585
R1163 B.n696 B.n695 585
R1164 B.n693 B.n346 585
R1165 B.n346 B.n345 585
R1166 B.n692 B.n691 585
R1167 B.n691 B.n690 585
R1168 B.n348 B.n347 585
R1169 B.n349 B.n348 585
R1170 B.n683 B.n682 585
R1171 B.n684 B.n683 585
R1172 B.n681 B.n354 585
R1173 B.n354 B.n353 585
R1174 B.n680 B.n679 585
R1175 B.n679 B.n678 585
R1176 B.n356 B.n355 585
R1177 B.n357 B.n356 585
R1178 B.n671 B.n670 585
R1179 B.n672 B.n671 585
R1180 B.n669 B.n362 585
R1181 B.n362 B.n361 585
R1182 B.n668 B.n667 585
R1183 B.n667 B.n666 585
R1184 B.n364 B.n363 585
R1185 B.n365 B.n364 585
R1186 B.n659 B.n658 585
R1187 B.n660 B.n659 585
R1188 B.n657 B.n370 585
R1189 B.n370 B.n369 585
R1190 B.n656 B.n655 585
R1191 B.n655 B.n654 585
R1192 B.n372 B.n371 585
R1193 B.n373 B.n372 585
R1194 B.n647 B.n646 585
R1195 B.n648 B.n647 585
R1196 B.n645 B.n378 585
R1197 B.n378 B.n377 585
R1198 B.n644 B.n643 585
R1199 B.n643 B.n642 585
R1200 B.n380 B.n379 585
R1201 B.n381 B.n380 585
R1202 B.n635 B.n634 585
R1203 B.n636 B.n635 585
R1204 B.n384 B.n383 585
R1205 B.n439 B.n437 585
R1206 B.n440 B.n436 585
R1207 B.n440 B.n385 585
R1208 B.n443 B.n442 585
R1209 B.n444 B.n435 585
R1210 B.n446 B.n445 585
R1211 B.n448 B.n434 585
R1212 B.n451 B.n450 585
R1213 B.n452 B.n433 585
R1214 B.n454 B.n453 585
R1215 B.n456 B.n432 585
R1216 B.n459 B.n458 585
R1217 B.n460 B.n431 585
R1218 B.n462 B.n461 585
R1219 B.n464 B.n430 585
R1220 B.n467 B.n466 585
R1221 B.n468 B.n429 585
R1222 B.n470 B.n469 585
R1223 B.n472 B.n428 585
R1224 B.n475 B.n474 585
R1225 B.n476 B.n427 585
R1226 B.n478 B.n477 585
R1227 B.n480 B.n426 585
R1228 B.n483 B.n482 585
R1229 B.n484 B.n425 585
R1230 B.n486 B.n485 585
R1231 B.n488 B.n424 585
R1232 B.n491 B.n490 585
R1233 B.n492 B.n423 585
R1234 B.n494 B.n493 585
R1235 B.n496 B.n422 585
R1236 B.n499 B.n498 585
R1237 B.n500 B.n421 585
R1238 B.n502 B.n501 585
R1239 B.n504 B.n420 585
R1240 B.n507 B.n506 585
R1241 B.n508 B.n419 585
R1242 B.n510 B.n509 585
R1243 B.n512 B.n418 585
R1244 B.n515 B.n514 585
R1245 B.n516 B.n417 585
R1246 B.n518 B.n517 585
R1247 B.n520 B.n416 585
R1248 B.n523 B.n522 585
R1249 B.n525 B.n413 585
R1250 B.n527 B.n526 585
R1251 B.n529 B.n412 585
R1252 B.n532 B.n531 585
R1253 B.n533 B.n411 585
R1254 B.n535 B.n534 585
R1255 B.n537 B.n410 585
R1256 B.n540 B.n539 585
R1257 B.n541 B.n409 585
R1258 B.n546 B.n545 585
R1259 B.n548 B.n408 585
R1260 B.n551 B.n550 585
R1261 B.n552 B.n407 585
R1262 B.n554 B.n553 585
R1263 B.n556 B.n406 585
R1264 B.n559 B.n558 585
R1265 B.n560 B.n405 585
R1266 B.n562 B.n561 585
R1267 B.n564 B.n404 585
R1268 B.n567 B.n566 585
R1269 B.n568 B.n403 585
R1270 B.n570 B.n569 585
R1271 B.n572 B.n402 585
R1272 B.n575 B.n574 585
R1273 B.n576 B.n401 585
R1274 B.n578 B.n577 585
R1275 B.n580 B.n400 585
R1276 B.n583 B.n582 585
R1277 B.n584 B.n399 585
R1278 B.n586 B.n585 585
R1279 B.n588 B.n398 585
R1280 B.n591 B.n590 585
R1281 B.n592 B.n397 585
R1282 B.n594 B.n593 585
R1283 B.n596 B.n396 585
R1284 B.n599 B.n598 585
R1285 B.n600 B.n395 585
R1286 B.n602 B.n601 585
R1287 B.n604 B.n394 585
R1288 B.n607 B.n606 585
R1289 B.n608 B.n393 585
R1290 B.n610 B.n609 585
R1291 B.n612 B.n392 585
R1292 B.n615 B.n614 585
R1293 B.n616 B.n391 585
R1294 B.n618 B.n617 585
R1295 B.n620 B.n390 585
R1296 B.n623 B.n622 585
R1297 B.n624 B.n389 585
R1298 B.n626 B.n625 585
R1299 B.n628 B.n388 585
R1300 B.n629 B.n387 585
R1301 B.n632 B.n631 585
R1302 B.n633 B.n386 585
R1303 B.n386 B.n385 585
R1304 B.n638 B.n637 585
R1305 B.n637 B.n636 585
R1306 B.n639 B.n382 585
R1307 B.n382 B.n381 585
R1308 B.n641 B.n640 585
R1309 B.n642 B.n641 585
R1310 B.n376 B.n375 585
R1311 B.n377 B.n376 585
R1312 B.n650 B.n649 585
R1313 B.n649 B.n648 585
R1314 B.n651 B.n374 585
R1315 B.n374 B.n373 585
R1316 B.n653 B.n652 585
R1317 B.n654 B.n653 585
R1318 B.n368 B.n367 585
R1319 B.n369 B.n368 585
R1320 B.n662 B.n661 585
R1321 B.n661 B.n660 585
R1322 B.n663 B.n366 585
R1323 B.n366 B.n365 585
R1324 B.n665 B.n664 585
R1325 B.n666 B.n665 585
R1326 B.n360 B.n359 585
R1327 B.n361 B.n360 585
R1328 B.n674 B.n673 585
R1329 B.n673 B.n672 585
R1330 B.n675 B.n358 585
R1331 B.n358 B.n357 585
R1332 B.n677 B.n676 585
R1333 B.n678 B.n677 585
R1334 B.n352 B.n351 585
R1335 B.n353 B.n352 585
R1336 B.n686 B.n685 585
R1337 B.n685 B.n684 585
R1338 B.n687 B.n350 585
R1339 B.n350 B.n349 585
R1340 B.n689 B.n688 585
R1341 B.n690 B.n689 585
R1342 B.n344 B.n343 585
R1343 B.n345 B.n344 585
R1344 B.n698 B.n697 585
R1345 B.n697 B.n696 585
R1346 B.n699 B.n342 585
R1347 B.n342 B.n341 585
R1348 B.n701 B.n700 585
R1349 B.n702 B.n701 585
R1350 B.n336 B.n335 585
R1351 B.n337 B.n336 585
R1352 B.n710 B.n709 585
R1353 B.n709 B.n708 585
R1354 B.n711 B.n334 585
R1355 B.n334 B.n333 585
R1356 B.n713 B.n712 585
R1357 B.n714 B.n713 585
R1358 B.n328 B.n327 585
R1359 B.n329 B.n328 585
R1360 B.n722 B.n721 585
R1361 B.n721 B.n720 585
R1362 B.n723 B.n326 585
R1363 B.n326 B.n324 585
R1364 B.n725 B.n724 585
R1365 B.n726 B.n725 585
R1366 B.n320 B.n319 585
R1367 B.n325 B.n320 585
R1368 B.n735 B.n734 585
R1369 B.n734 B.n733 585
R1370 B.n736 B.n318 585
R1371 B.n318 B.n317 585
R1372 B.n738 B.n737 585
R1373 B.n739 B.n738 585
R1374 B.n2 B.n0 585
R1375 B.n4 B.n2 585
R1376 B.n3 B.n1 585
R1377 B.n864 B.n3 585
R1378 B.n862 B.n861 585
R1379 B.n863 B.n862 585
R1380 B.n860 B.n9 585
R1381 B.n9 B.n8 585
R1382 B.n859 B.n858 585
R1383 B.n858 B.n857 585
R1384 B.n11 B.n10 585
R1385 B.n856 B.n11 585
R1386 B.n854 B.n853 585
R1387 B.n855 B.n854 585
R1388 B.n852 B.n16 585
R1389 B.n16 B.n15 585
R1390 B.n851 B.n850 585
R1391 B.n850 B.n849 585
R1392 B.n18 B.n17 585
R1393 B.n848 B.n18 585
R1394 B.n846 B.n845 585
R1395 B.n847 B.n846 585
R1396 B.n844 B.n23 585
R1397 B.n23 B.n22 585
R1398 B.n843 B.n842 585
R1399 B.n842 B.n841 585
R1400 B.n25 B.n24 585
R1401 B.n840 B.n25 585
R1402 B.n838 B.n837 585
R1403 B.n839 B.n838 585
R1404 B.n836 B.n30 585
R1405 B.n30 B.n29 585
R1406 B.n835 B.n834 585
R1407 B.n834 B.n833 585
R1408 B.n32 B.n31 585
R1409 B.n832 B.n32 585
R1410 B.n830 B.n829 585
R1411 B.n831 B.n830 585
R1412 B.n828 B.n37 585
R1413 B.n37 B.n36 585
R1414 B.n827 B.n826 585
R1415 B.n826 B.n825 585
R1416 B.n39 B.n38 585
R1417 B.n824 B.n39 585
R1418 B.n822 B.n821 585
R1419 B.n823 B.n822 585
R1420 B.n820 B.n44 585
R1421 B.n44 B.n43 585
R1422 B.n819 B.n818 585
R1423 B.n818 B.n817 585
R1424 B.n46 B.n45 585
R1425 B.n816 B.n46 585
R1426 B.n814 B.n813 585
R1427 B.n815 B.n814 585
R1428 B.n812 B.n51 585
R1429 B.n51 B.n50 585
R1430 B.n811 B.n810 585
R1431 B.n810 B.n809 585
R1432 B.n53 B.n52 585
R1433 B.n808 B.n53 585
R1434 B.n806 B.n805 585
R1435 B.n807 B.n806 585
R1436 B.n804 B.n58 585
R1437 B.n58 B.n57 585
R1438 B.n803 B.n802 585
R1439 B.n802 B.n801 585
R1440 B.n60 B.n59 585
R1441 B.n800 B.n60 585
R1442 B.n798 B.n797 585
R1443 B.n799 B.n798 585
R1444 B.n796 B.n65 585
R1445 B.n65 B.n64 585
R1446 B.n795 B.n794 585
R1447 B.n794 B.n793 585
R1448 B.n867 B.n866 585
R1449 B.n866 B.n865 585
R1450 B.n637 B.n384 497.305
R1451 B.n794 B.n67 497.305
R1452 B.n635 B.n386 497.305
R1453 B.n790 B.n68 497.305
R1454 B.n542 B.t8 403.096
R1455 B.n414 B.t19 403.096
R1456 B.n121 B.t16 403.096
R1457 B.n118 B.t12 403.096
R1458 B.n542 B.t11 334.06
R1459 B.n118 B.t14 334.06
R1460 B.n414 B.t21 334.06
R1461 B.n121 B.t17 334.06
R1462 B.n543 B.t10 297.212
R1463 B.n119 B.t15 297.212
R1464 B.n415 B.t20 297.212
R1465 B.n122 B.t18 297.212
R1466 B.n792 B.n791 256.663
R1467 B.n792 B.n116 256.663
R1468 B.n792 B.n115 256.663
R1469 B.n792 B.n114 256.663
R1470 B.n792 B.n113 256.663
R1471 B.n792 B.n112 256.663
R1472 B.n792 B.n111 256.663
R1473 B.n792 B.n110 256.663
R1474 B.n792 B.n109 256.663
R1475 B.n792 B.n108 256.663
R1476 B.n792 B.n107 256.663
R1477 B.n792 B.n106 256.663
R1478 B.n792 B.n105 256.663
R1479 B.n792 B.n104 256.663
R1480 B.n792 B.n103 256.663
R1481 B.n792 B.n102 256.663
R1482 B.n792 B.n101 256.663
R1483 B.n792 B.n100 256.663
R1484 B.n792 B.n99 256.663
R1485 B.n792 B.n98 256.663
R1486 B.n792 B.n97 256.663
R1487 B.n792 B.n96 256.663
R1488 B.n792 B.n95 256.663
R1489 B.n792 B.n94 256.663
R1490 B.n792 B.n93 256.663
R1491 B.n792 B.n92 256.663
R1492 B.n792 B.n91 256.663
R1493 B.n792 B.n90 256.663
R1494 B.n792 B.n89 256.663
R1495 B.n792 B.n88 256.663
R1496 B.n792 B.n87 256.663
R1497 B.n792 B.n86 256.663
R1498 B.n792 B.n85 256.663
R1499 B.n792 B.n84 256.663
R1500 B.n792 B.n83 256.663
R1501 B.n792 B.n82 256.663
R1502 B.n792 B.n81 256.663
R1503 B.n792 B.n80 256.663
R1504 B.n792 B.n79 256.663
R1505 B.n792 B.n78 256.663
R1506 B.n792 B.n77 256.663
R1507 B.n792 B.n76 256.663
R1508 B.n792 B.n75 256.663
R1509 B.n792 B.n74 256.663
R1510 B.n792 B.n73 256.663
R1511 B.n792 B.n72 256.663
R1512 B.n792 B.n71 256.663
R1513 B.n792 B.n70 256.663
R1514 B.n792 B.n69 256.663
R1515 B.n438 B.n385 256.663
R1516 B.n441 B.n385 256.663
R1517 B.n447 B.n385 256.663
R1518 B.n449 B.n385 256.663
R1519 B.n455 B.n385 256.663
R1520 B.n457 B.n385 256.663
R1521 B.n463 B.n385 256.663
R1522 B.n465 B.n385 256.663
R1523 B.n471 B.n385 256.663
R1524 B.n473 B.n385 256.663
R1525 B.n479 B.n385 256.663
R1526 B.n481 B.n385 256.663
R1527 B.n487 B.n385 256.663
R1528 B.n489 B.n385 256.663
R1529 B.n495 B.n385 256.663
R1530 B.n497 B.n385 256.663
R1531 B.n503 B.n385 256.663
R1532 B.n505 B.n385 256.663
R1533 B.n511 B.n385 256.663
R1534 B.n513 B.n385 256.663
R1535 B.n519 B.n385 256.663
R1536 B.n521 B.n385 256.663
R1537 B.n528 B.n385 256.663
R1538 B.n530 B.n385 256.663
R1539 B.n536 B.n385 256.663
R1540 B.n538 B.n385 256.663
R1541 B.n547 B.n385 256.663
R1542 B.n549 B.n385 256.663
R1543 B.n555 B.n385 256.663
R1544 B.n557 B.n385 256.663
R1545 B.n563 B.n385 256.663
R1546 B.n565 B.n385 256.663
R1547 B.n571 B.n385 256.663
R1548 B.n573 B.n385 256.663
R1549 B.n579 B.n385 256.663
R1550 B.n581 B.n385 256.663
R1551 B.n587 B.n385 256.663
R1552 B.n589 B.n385 256.663
R1553 B.n595 B.n385 256.663
R1554 B.n597 B.n385 256.663
R1555 B.n603 B.n385 256.663
R1556 B.n605 B.n385 256.663
R1557 B.n611 B.n385 256.663
R1558 B.n613 B.n385 256.663
R1559 B.n619 B.n385 256.663
R1560 B.n621 B.n385 256.663
R1561 B.n627 B.n385 256.663
R1562 B.n630 B.n385 256.663
R1563 B.n637 B.n382 163.367
R1564 B.n641 B.n382 163.367
R1565 B.n641 B.n376 163.367
R1566 B.n649 B.n376 163.367
R1567 B.n649 B.n374 163.367
R1568 B.n653 B.n374 163.367
R1569 B.n653 B.n368 163.367
R1570 B.n661 B.n368 163.367
R1571 B.n661 B.n366 163.367
R1572 B.n665 B.n366 163.367
R1573 B.n665 B.n360 163.367
R1574 B.n673 B.n360 163.367
R1575 B.n673 B.n358 163.367
R1576 B.n677 B.n358 163.367
R1577 B.n677 B.n352 163.367
R1578 B.n685 B.n352 163.367
R1579 B.n685 B.n350 163.367
R1580 B.n689 B.n350 163.367
R1581 B.n689 B.n344 163.367
R1582 B.n697 B.n344 163.367
R1583 B.n697 B.n342 163.367
R1584 B.n701 B.n342 163.367
R1585 B.n701 B.n336 163.367
R1586 B.n709 B.n336 163.367
R1587 B.n709 B.n334 163.367
R1588 B.n713 B.n334 163.367
R1589 B.n713 B.n328 163.367
R1590 B.n721 B.n328 163.367
R1591 B.n721 B.n326 163.367
R1592 B.n725 B.n326 163.367
R1593 B.n725 B.n320 163.367
R1594 B.n734 B.n320 163.367
R1595 B.n734 B.n318 163.367
R1596 B.n738 B.n318 163.367
R1597 B.n738 B.n2 163.367
R1598 B.n866 B.n2 163.367
R1599 B.n866 B.n3 163.367
R1600 B.n862 B.n3 163.367
R1601 B.n862 B.n9 163.367
R1602 B.n858 B.n9 163.367
R1603 B.n858 B.n11 163.367
R1604 B.n854 B.n11 163.367
R1605 B.n854 B.n16 163.367
R1606 B.n850 B.n16 163.367
R1607 B.n850 B.n18 163.367
R1608 B.n846 B.n18 163.367
R1609 B.n846 B.n23 163.367
R1610 B.n842 B.n23 163.367
R1611 B.n842 B.n25 163.367
R1612 B.n838 B.n25 163.367
R1613 B.n838 B.n30 163.367
R1614 B.n834 B.n30 163.367
R1615 B.n834 B.n32 163.367
R1616 B.n830 B.n32 163.367
R1617 B.n830 B.n37 163.367
R1618 B.n826 B.n37 163.367
R1619 B.n826 B.n39 163.367
R1620 B.n822 B.n39 163.367
R1621 B.n822 B.n44 163.367
R1622 B.n818 B.n44 163.367
R1623 B.n818 B.n46 163.367
R1624 B.n814 B.n46 163.367
R1625 B.n814 B.n51 163.367
R1626 B.n810 B.n51 163.367
R1627 B.n810 B.n53 163.367
R1628 B.n806 B.n53 163.367
R1629 B.n806 B.n58 163.367
R1630 B.n802 B.n58 163.367
R1631 B.n802 B.n60 163.367
R1632 B.n798 B.n60 163.367
R1633 B.n798 B.n65 163.367
R1634 B.n794 B.n65 163.367
R1635 B.n440 B.n439 163.367
R1636 B.n442 B.n440 163.367
R1637 B.n446 B.n435 163.367
R1638 B.n450 B.n448 163.367
R1639 B.n454 B.n433 163.367
R1640 B.n458 B.n456 163.367
R1641 B.n462 B.n431 163.367
R1642 B.n466 B.n464 163.367
R1643 B.n470 B.n429 163.367
R1644 B.n474 B.n472 163.367
R1645 B.n478 B.n427 163.367
R1646 B.n482 B.n480 163.367
R1647 B.n486 B.n425 163.367
R1648 B.n490 B.n488 163.367
R1649 B.n494 B.n423 163.367
R1650 B.n498 B.n496 163.367
R1651 B.n502 B.n421 163.367
R1652 B.n506 B.n504 163.367
R1653 B.n510 B.n419 163.367
R1654 B.n514 B.n512 163.367
R1655 B.n518 B.n417 163.367
R1656 B.n522 B.n520 163.367
R1657 B.n527 B.n413 163.367
R1658 B.n531 B.n529 163.367
R1659 B.n535 B.n411 163.367
R1660 B.n539 B.n537 163.367
R1661 B.n546 B.n409 163.367
R1662 B.n550 B.n548 163.367
R1663 B.n554 B.n407 163.367
R1664 B.n558 B.n556 163.367
R1665 B.n562 B.n405 163.367
R1666 B.n566 B.n564 163.367
R1667 B.n570 B.n403 163.367
R1668 B.n574 B.n572 163.367
R1669 B.n578 B.n401 163.367
R1670 B.n582 B.n580 163.367
R1671 B.n586 B.n399 163.367
R1672 B.n590 B.n588 163.367
R1673 B.n594 B.n397 163.367
R1674 B.n598 B.n596 163.367
R1675 B.n602 B.n395 163.367
R1676 B.n606 B.n604 163.367
R1677 B.n610 B.n393 163.367
R1678 B.n614 B.n612 163.367
R1679 B.n618 B.n391 163.367
R1680 B.n622 B.n620 163.367
R1681 B.n626 B.n389 163.367
R1682 B.n629 B.n628 163.367
R1683 B.n631 B.n386 163.367
R1684 B.n635 B.n380 163.367
R1685 B.n643 B.n380 163.367
R1686 B.n643 B.n378 163.367
R1687 B.n647 B.n378 163.367
R1688 B.n647 B.n372 163.367
R1689 B.n655 B.n372 163.367
R1690 B.n655 B.n370 163.367
R1691 B.n659 B.n370 163.367
R1692 B.n659 B.n364 163.367
R1693 B.n667 B.n364 163.367
R1694 B.n667 B.n362 163.367
R1695 B.n671 B.n362 163.367
R1696 B.n671 B.n356 163.367
R1697 B.n679 B.n356 163.367
R1698 B.n679 B.n354 163.367
R1699 B.n683 B.n354 163.367
R1700 B.n683 B.n348 163.367
R1701 B.n691 B.n348 163.367
R1702 B.n691 B.n346 163.367
R1703 B.n695 B.n346 163.367
R1704 B.n695 B.n340 163.367
R1705 B.n703 B.n340 163.367
R1706 B.n703 B.n338 163.367
R1707 B.n707 B.n338 163.367
R1708 B.n707 B.n332 163.367
R1709 B.n715 B.n332 163.367
R1710 B.n715 B.n330 163.367
R1711 B.n719 B.n330 163.367
R1712 B.n719 B.n323 163.367
R1713 B.n727 B.n323 163.367
R1714 B.n727 B.n321 163.367
R1715 B.n732 B.n321 163.367
R1716 B.n732 B.n316 163.367
R1717 B.n740 B.n316 163.367
R1718 B.n741 B.n740 163.367
R1719 B.n741 B.n5 163.367
R1720 B.n6 B.n5 163.367
R1721 B.n7 B.n6 163.367
R1722 B.n746 B.n7 163.367
R1723 B.n746 B.n12 163.367
R1724 B.n13 B.n12 163.367
R1725 B.n14 B.n13 163.367
R1726 B.n751 B.n14 163.367
R1727 B.n751 B.n19 163.367
R1728 B.n20 B.n19 163.367
R1729 B.n21 B.n20 163.367
R1730 B.n756 B.n21 163.367
R1731 B.n756 B.n26 163.367
R1732 B.n27 B.n26 163.367
R1733 B.n28 B.n27 163.367
R1734 B.n761 B.n28 163.367
R1735 B.n761 B.n33 163.367
R1736 B.n34 B.n33 163.367
R1737 B.n35 B.n34 163.367
R1738 B.n766 B.n35 163.367
R1739 B.n766 B.n40 163.367
R1740 B.n41 B.n40 163.367
R1741 B.n42 B.n41 163.367
R1742 B.n771 B.n42 163.367
R1743 B.n771 B.n47 163.367
R1744 B.n48 B.n47 163.367
R1745 B.n49 B.n48 163.367
R1746 B.n776 B.n49 163.367
R1747 B.n776 B.n54 163.367
R1748 B.n55 B.n54 163.367
R1749 B.n56 B.n55 163.367
R1750 B.n781 B.n56 163.367
R1751 B.n781 B.n61 163.367
R1752 B.n62 B.n61 163.367
R1753 B.n63 B.n62 163.367
R1754 B.n786 B.n63 163.367
R1755 B.n786 B.n68 163.367
R1756 B.n126 B.n125 163.367
R1757 B.n130 B.n129 163.367
R1758 B.n134 B.n133 163.367
R1759 B.n138 B.n137 163.367
R1760 B.n142 B.n141 163.367
R1761 B.n146 B.n145 163.367
R1762 B.n150 B.n149 163.367
R1763 B.n154 B.n153 163.367
R1764 B.n158 B.n157 163.367
R1765 B.n162 B.n161 163.367
R1766 B.n166 B.n165 163.367
R1767 B.n170 B.n169 163.367
R1768 B.n174 B.n173 163.367
R1769 B.n178 B.n177 163.367
R1770 B.n182 B.n181 163.367
R1771 B.n186 B.n185 163.367
R1772 B.n190 B.n189 163.367
R1773 B.n194 B.n193 163.367
R1774 B.n198 B.n197 163.367
R1775 B.n202 B.n201 163.367
R1776 B.n206 B.n205 163.367
R1777 B.n210 B.n209 163.367
R1778 B.n214 B.n213 163.367
R1779 B.n218 B.n217 163.367
R1780 B.n222 B.n221 163.367
R1781 B.n226 B.n225 163.367
R1782 B.n230 B.n229 163.367
R1783 B.n234 B.n233 163.367
R1784 B.n238 B.n237 163.367
R1785 B.n242 B.n241 163.367
R1786 B.n246 B.n245 163.367
R1787 B.n250 B.n249 163.367
R1788 B.n254 B.n253 163.367
R1789 B.n258 B.n257 163.367
R1790 B.n262 B.n261 163.367
R1791 B.n266 B.n265 163.367
R1792 B.n270 B.n269 163.367
R1793 B.n274 B.n273 163.367
R1794 B.n278 B.n277 163.367
R1795 B.n282 B.n281 163.367
R1796 B.n286 B.n285 163.367
R1797 B.n290 B.n289 163.367
R1798 B.n294 B.n293 163.367
R1799 B.n298 B.n297 163.367
R1800 B.n302 B.n301 163.367
R1801 B.n306 B.n305 163.367
R1802 B.n310 B.n309 163.367
R1803 B.n312 B.n117 163.367
R1804 B.n636 B.n385 77.0339
R1805 B.n793 B.n792 77.0339
R1806 B.n438 B.n384 71.676
R1807 B.n442 B.n441 71.676
R1808 B.n447 B.n446 71.676
R1809 B.n450 B.n449 71.676
R1810 B.n455 B.n454 71.676
R1811 B.n458 B.n457 71.676
R1812 B.n463 B.n462 71.676
R1813 B.n466 B.n465 71.676
R1814 B.n471 B.n470 71.676
R1815 B.n474 B.n473 71.676
R1816 B.n479 B.n478 71.676
R1817 B.n482 B.n481 71.676
R1818 B.n487 B.n486 71.676
R1819 B.n490 B.n489 71.676
R1820 B.n495 B.n494 71.676
R1821 B.n498 B.n497 71.676
R1822 B.n503 B.n502 71.676
R1823 B.n506 B.n505 71.676
R1824 B.n511 B.n510 71.676
R1825 B.n514 B.n513 71.676
R1826 B.n519 B.n518 71.676
R1827 B.n522 B.n521 71.676
R1828 B.n528 B.n527 71.676
R1829 B.n531 B.n530 71.676
R1830 B.n536 B.n535 71.676
R1831 B.n539 B.n538 71.676
R1832 B.n547 B.n546 71.676
R1833 B.n550 B.n549 71.676
R1834 B.n555 B.n554 71.676
R1835 B.n558 B.n557 71.676
R1836 B.n563 B.n562 71.676
R1837 B.n566 B.n565 71.676
R1838 B.n571 B.n570 71.676
R1839 B.n574 B.n573 71.676
R1840 B.n579 B.n578 71.676
R1841 B.n582 B.n581 71.676
R1842 B.n587 B.n586 71.676
R1843 B.n590 B.n589 71.676
R1844 B.n595 B.n594 71.676
R1845 B.n598 B.n597 71.676
R1846 B.n603 B.n602 71.676
R1847 B.n606 B.n605 71.676
R1848 B.n611 B.n610 71.676
R1849 B.n614 B.n613 71.676
R1850 B.n619 B.n618 71.676
R1851 B.n622 B.n621 71.676
R1852 B.n627 B.n626 71.676
R1853 B.n630 B.n629 71.676
R1854 B.n69 B.n67 71.676
R1855 B.n126 B.n70 71.676
R1856 B.n130 B.n71 71.676
R1857 B.n134 B.n72 71.676
R1858 B.n138 B.n73 71.676
R1859 B.n142 B.n74 71.676
R1860 B.n146 B.n75 71.676
R1861 B.n150 B.n76 71.676
R1862 B.n154 B.n77 71.676
R1863 B.n158 B.n78 71.676
R1864 B.n162 B.n79 71.676
R1865 B.n166 B.n80 71.676
R1866 B.n170 B.n81 71.676
R1867 B.n174 B.n82 71.676
R1868 B.n178 B.n83 71.676
R1869 B.n182 B.n84 71.676
R1870 B.n186 B.n85 71.676
R1871 B.n190 B.n86 71.676
R1872 B.n194 B.n87 71.676
R1873 B.n198 B.n88 71.676
R1874 B.n202 B.n89 71.676
R1875 B.n206 B.n90 71.676
R1876 B.n210 B.n91 71.676
R1877 B.n214 B.n92 71.676
R1878 B.n218 B.n93 71.676
R1879 B.n222 B.n94 71.676
R1880 B.n226 B.n95 71.676
R1881 B.n230 B.n96 71.676
R1882 B.n234 B.n97 71.676
R1883 B.n238 B.n98 71.676
R1884 B.n242 B.n99 71.676
R1885 B.n246 B.n100 71.676
R1886 B.n250 B.n101 71.676
R1887 B.n254 B.n102 71.676
R1888 B.n258 B.n103 71.676
R1889 B.n262 B.n104 71.676
R1890 B.n266 B.n105 71.676
R1891 B.n270 B.n106 71.676
R1892 B.n274 B.n107 71.676
R1893 B.n278 B.n108 71.676
R1894 B.n282 B.n109 71.676
R1895 B.n286 B.n110 71.676
R1896 B.n290 B.n111 71.676
R1897 B.n294 B.n112 71.676
R1898 B.n298 B.n113 71.676
R1899 B.n302 B.n114 71.676
R1900 B.n306 B.n115 71.676
R1901 B.n310 B.n116 71.676
R1902 B.n791 B.n117 71.676
R1903 B.n791 B.n790 71.676
R1904 B.n312 B.n116 71.676
R1905 B.n309 B.n115 71.676
R1906 B.n305 B.n114 71.676
R1907 B.n301 B.n113 71.676
R1908 B.n297 B.n112 71.676
R1909 B.n293 B.n111 71.676
R1910 B.n289 B.n110 71.676
R1911 B.n285 B.n109 71.676
R1912 B.n281 B.n108 71.676
R1913 B.n277 B.n107 71.676
R1914 B.n273 B.n106 71.676
R1915 B.n269 B.n105 71.676
R1916 B.n265 B.n104 71.676
R1917 B.n261 B.n103 71.676
R1918 B.n257 B.n102 71.676
R1919 B.n253 B.n101 71.676
R1920 B.n249 B.n100 71.676
R1921 B.n245 B.n99 71.676
R1922 B.n241 B.n98 71.676
R1923 B.n237 B.n97 71.676
R1924 B.n233 B.n96 71.676
R1925 B.n229 B.n95 71.676
R1926 B.n225 B.n94 71.676
R1927 B.n221 B.n93 71.676
R1928 B.n217 B.n92 71.676
R1929 B.n213 B.n91 71.676
R1930 B.n209 B.n90 71.676
R1931 B.n205 B.n89 71.676
R1932 B.n201 B.n88 71.676
R1933 B.n197 B.n87 71.676
R1934 B.n193 B.n86 71.676
R1935 B.n189 B.n85 71.676
R1936 B.n185 B.n84 71.676
R1937 B.n181 B.n83 71.676
R1938 B.n177 B.n82 71.676
R1939 B.n173 B.n81 71.676
R1940 B.n169 B.n80 71.676
R1941 B.n165 B.n79 71.676
R1942 B.n161 B.n78 71.676
R1943 B.n157 B.n77 71.676
R1944 B.n153 B.n76 71.676
R1945 B.n149 B.n75 71.676
R1946 B.n145 B.n74 71.676
R1947 B.n141 B.n73 71.676
R1948 B.n137 B.n72 71.676
R1949 B.n133 B.n71 71.676
R1950 B.n129 B.n70 71.676
R1951 B.n125 B.n69 71.676
R1952 B.n439 B.n438 71.676
R1953 B.n441 B.n435 71.676
R1954 B.n448 B.n447 71.676
R1955 B.n449 B.n433 71.676
R1956 B.n456 B.n455 71.676
R1957 B.n457 B.n431 71.676
R1958 B.n464 B.n463 71.676
R1959 B.n465 B.n429 71.676
R1960 B.n472 B.n471 71.676
R1961 B.n473 B.n427 71.676
R1962 B.n480 B.n479 71.676
R1963 B.n481 B.n425 71.676
R1964 B.n488 B.n487 71.676
R1965 B.n489 B.n423 71.676
R1966 B.n496 B.n495 71.676
R1967 B.n497 B.n421 71.676
R1968 B.n504 B.n503 71.676
R1969 B.n505 B.n419 71.676
R1970 B.n512 B.n511 71.676
R1971 B.n513 B.n417 71.676
R1972 B.n520 B.n519 71.676
R1973 B.n521 B.n413 71.676
R1974 B.n529 B.n528 71.676
R1975 B.n530 B.n411 71.676
R1976 B.n537 B.n536 71.676
R1977 B.n538 B.n409 71.676
R1978 B.n548 B.n547 71.676
R1979 B.n549 B.n407 71.676
R1980 B.n556 B.n555 71.676
R1981 B.n557 B.n405 71.676
R1982 B.n564 B.n563 71.676
R1983 B.n565 B.n403 71.676
R1984 B.n572 B.n571 71.676
R1985 B.n573 B.n401 71.676
R1986 B.n580 B.n579 71.676
R1987 B.n581 B.n399 71.676
R1988 B.n588 B.n587 71.676
R1989 B.n589 B.n397 71.676
R1990 B.n596 B.n595 71.676
R1991 B.n597 B.n395 71.676
R1992 B.n604 B.n603 71.676
R1993 B.n605 B.n393 71.676
R1994 B.n612 B.n611 71.676
R1995 B.n613 B.n391 71.676
R1996 B.n620 B.n619 71.676
R1997 B.n621 B.n389 71.676
R1998 B.n628 B.n627 71.676
R1999 B.n631 B.n630 71.676
R2000 B.n544 B.n543 59.5399
R2001 B.n524 B.n415 59.5399
R2002 B.n123 B.n122 59.5399
R2003 B.n120 B.n119 59.5399
R2004 B.n636 B.n381 41.2467
R2005 B.n642 B.n381 41.2467
R2006 B.n642 B.n377 41.2467
R2007 B.n648 B.n377 41.2467
R2008 B.n648 B.n373 41.2467
R2009 B.n654 B.n373 41.2467
R2010 B.n660 B.n369 41.2467
R2011 B.n660 B.n365 41.2467
R2012 B.n666 B.n365 41.2467
R2013 B.n666 B.n361 41.2467
R2014 B.n672 B.n361 41.2467
R2015 B.n672 B.n357 41.2467
R2016 B.n678 B.n357 41.2467
R2017 B.n684 B.n353 41.2467
R2018 B.n684 B.n349 41.2467
R2019 B.n690 B.n349 41.2467
R2020 B.n690 B.n345 41.2467
R2021 B.n696 B.n345 41.2467
R2022 B.n702 B.n341 41.2467
R2023 B.n702 B.n337 41.2467
R2024 B.n708 B.n337 41.2467
R2025 B.n708 B.n333 41.2467
R2026 B.n714 B.n333 41.2467
R2027 B.n720 B.n329 41.2467
R2028 B.n720 B.n324 41.2467
R2029 B.n726 B.n324 41.2467
R2030 B.n726 B.n325 41.2467
R2031 B.n733 B.n317 41.2467
R2032 B.n739 B.n317 41.2467
R2033 B.n739 B.n4 41.2467
R2034 B.n865 B.n4 41.2467
R2035 B.n865 B.n864 41.2467
R2036 B.n864 B.n863 41.2467
R2037 B.n863 B.n8 41.2467
R2038 B.n857 B.n8 41.2467
R2039 B.n856 B.n855 41.2467
R2040 B.n855 B.n15 41.2467
R2041 B.n849 B.n15 41.2467
R2042 B.n849 B.n848 41.2467
R2043 B.n847 B.n22 41.2467
R2044 B.n841 B.n22 41.2467
R2045 B.n841 B.n840 41.2467
R2046 B.n840 B.n839 41.2467
R2047 B.n839 B.n29 41.2467
R2048 B.n833 B.n832 41.2467
R2049 B.n832 B.n831 41.2467
R2050 B.n831 B.n36 41.2467
R2051 B.n825 B.n36 41.2467
R2052 B.n825 B.n824 41.2467
R2053 B.n823 B.n43 41.2467
R2054 B.n817 B.n43 41.2467
R2055 B.n817 B.n816 41.2467
R2056 B.n816 B.n815 41.2467
R2057 B.n815 B.n50 41.2467
R2058 B.n809 B.n50 41.2467
R2059 B.n809 B.n808 41.2467
R2060 B.n807 B.n57 41.2467
R2061 B.n801 B.n57 41.2467
R2062 B.n801 B.n800 41.2467
R2063 B.n800 B.n799 41.2467
R2064 B.n799 B.n64 41.2467
R2065 B.n793 B.n64 41.2467
R2066 B.t3 B.n329 40.6401
R2067 B.n848 B.t0 40.6401
R2068 B.t9 B.n369 39.427
R2069 B.n808 B.t13 39.427
R2070 B.n543 B.n542 36.849
R2071 B.n415 B.n414 36.849
R2072 B.n122 B.n121 36.849
R2073 B.n119 B.n118 36.849
R2074 B.n678 B.t2 34.5745
R2075 B.t6 B.n823 34.5745
R2076 B.n795 B.n66 32.3127
R2077 B.n789 B.n788 32.3127
R2078 B.n634 B.n633 32.3127
R2079 B.n638 B.n383 32.3127
R2080 B.n325 B.t5 24.8695
R2081 B.t4 B.n856 24.8695
R2082 B.t1 B.n341 23.6564
R2083 B.t7 B.n29 23.6564
R2084 B B.n867 18.0485
R2085 B.n696 B.t1 17.5908
R2086 B.n833 B.t7 17.5908
R2087 B.n733 B.t5 16.3777
R2088 B.n857 B.t4 16.3777
R2089 B.n124 B.n66 10.6151
R2090 B.n127 B.n124 10.6151
R2091 B.n128 B.n127 10.6151
R2092 B.n131 B.n128 10.6151
R2093 B.n132 B.n131 10.6151
R2094 B.n135 B.n132 10.6151
R2095 B.n136 B.n135 10.6151
R2096 B.n139 B.n136 10.6151
R2097 B.n140 B.n139 10.6151
R2098 B.n143 B.n140 10.6151
R2099 B.n144 B.n143 10.6151
R2100 B.n147 B.n144 10.6151
R2101 B.n148 B.n147 10.6151
R2102 B.n151 B.n148 10.6151
R2103 B.n152 B.n151 10.6151
R2104 B.n155 B.n152 10.6151
R2105 B.n156 B.n155 10.6151
R2106 B.n159 B.n156 10.6151
R2107 B.n160 B.n159 10.6151
R2108 B.n163 B.n160 10.6151
R2109 B.n164 B.n163 10.6151
R2110 B.n167 B.n164 10.6151
R2111 B.n168 B.n167 10.6151
R2112 B.n171 B.n168 10.6151
R2113 B.n172 B.n171 10.6151
R2114 B.n175 B.n172 10.6151
R2115 B.n176 B.n175 10.6151
R2116 B.n179 B.n176 10.6151
R2117 B.n180 B.n179 10.6151
R2118 B.n183 B.n180 10.6151
R2119 B.n184 B.n183 10.6151
R2120 B.n187 B.n184 10.6151
R2121 B.n188 B.n187 10.6151
R2122 B.n191 B.n188 10.6151
R2123 B.n192 B.n191 10.6151
R2124 B.n195 B.n192 10.6151
R2125 B.n196 B.n195 10.6151
R2126 B.n199 B.n196 10.6151
R2127 B.n200 B.n199 10.6151
R2128 B.n203 B.n200 10.6151
R2129 B.n204 B.n203 10.6151
R2130 B.n207 B.n204 10.6151
R2131 B.n208 B.n207 10.6151
R2132 B.n212 B.n211 10.6151
R2133 B.n215 B.n212 10.6151
R2134 B.n216 B.n215 10.6151
R2135 B.n219 B.n216 10.6151
R2136 B.n220 B.n219 10.6151
R2137 B.n223 B.n220 10.6151
R2138 B.n224 B.n223 10.6151
R2139 B.n227 B.n224 10.6151
R2140 B.n228 B.n227 10.6151
R2141 B.n232 B.n231 10.6151
R2142 B.n235 B.n232 10.6151
R2143 B.n236 B.n235 10.6151
R2144 B.n239 B.n236 10.6151
R2145 B.n240 B.n239 10.6151
R2146 B.n243 B.n240 10.6151
R2147 B.n244 B.n243 10.6151
R2148 B.n247 B.n244 10.6151
R2149 B.n248 B.n247 10.6151
R2150 B.n251 B.n248 10.6151
R2151 B.n252 B.n251 10.6151
R2152 B.n255 B.n252 10.6151
R2153 B.n256 B.n255 10.6151
R2154 B.n259 B.n256 10.6151
R2155 B.n260 B.n259 10.6151
R2156 B.n263 B.n260 10.6151
R2157 B.n264 B.n263 10.6151
R2158 B.n267 B.n264 10.6151
R2159 B.n268 B.n267 10.6151
R2160 B.n271 B.n268 10.6151
R2161 B.n272 B.n271 10.6151
R2162 B.n275 B.n272 10.6151
R2163 B.n276 B.n275 10.6151
R2164 B.n279 B.n276 10.6151
R2165 B.n280 B.n279 10.6151
R2166 B.n283 B.n280 10.6151
R2167 B.n284 B.n283 10.6151
R2168 B.n287 B.n284 10.6151
R2169 B.n288 B.n287 10.6151
R2170 B.n291 B.n288 10.6151
R2171 B.n292 B.n291 10.6151
R2172 B.n295 B.n292 10.6151
R2173 B.n296 B.n295 10.6151
R2174 B.n299 B.n296 10.6151
R2175 B.n300 B.n299 10.6151
R2176 B.n303 B.n300 10.6151
R2177 B.n304 B.n303 10.6151
R2178 B.n307 B.n304 10.6151
R2179 B.n308 B.n307 10.6151
R2180 B.n311 B.n308 10.6151
R2181 B.n313 B.n311 10.6151
R2182 B.n314 B.n313 10.6151
R2183 B.n789 B.n314 10.6151
R2184 B.n634 B.n379 10.6151
R2185 B.n644 B.n379 10.6151
R2186 B.n645 B.n644 10.6151
R2187 B.n646 B.n645 10.6151
R2188 B.n646 B.n371 10.6151
R2189 B.n656 B.n371 10.6151
R2190 B.n657 B.n656 10.6151
R2191 B.n658 B.n657 10.6151
R2192 B.n658 B.n363 10.6151
R2193 B.n668 B.n363 10.6151
R2194 B.n669 B.n668 10.6151
R2195 B.n670 B.n669 10.6151
R2196 B.n670 B.n355 10.6151
R2197 B.n680 B.n355 10.6151
R2198 B.n681 B.n680 10.6151
R2199 B.n682 B.n681 10.6151
R2200 B.n682 B.n347 10.6151
R2201 B.n692 B.n347 10.6151
R2202 B.n693 B.n692 10.6151
R2203 B.n694 B.n693 10.6151
R2204 B.n694 B.n339 10.6151
R2205 B.n704 B.n339 10.6151
R2206 B.n705 B.n704 10.6151
R2207 B.n706 B.n705 10.6151
R2208 B.n706 B.n331 10.6151
R2209 B.n716 B.n331 10.6151
R2210 B.n717 B.n716 10.6151
R2211 B.n718 B.n717 10.6151
R2212 B.n718 B.n322 10.6151
R2213 B.n728 B.n322 10.6151
R2214 B.n729 B.n728 10.6151
R2215 B.n731 B.n729 10.6151
R2216 B.n731 B.n730 10.6151
R2217 B.n730 B.n315 10.6151
R2218 B.n742 B.n315 10.6151
R2219 B.n743 B.n742 10.6151
R2220 B.n744 B.n743 10.6151
R2221 B.n745 B.n744 10.6151
R2222 B.n747 B.n745 10.6151
R2223 B.n748 B.n747 10.6151
R2224 B.n749 B.n748 10.6151
R2225 B.n750 B.n749 10.6151
R2226 B.n752 B.n750 10.6151
R2227 B.n753 B.n752 10.6151
R2228 B.n754 B.n753 10.6151
R2229 B.n755 B.n754 10.6151
R2230 B.n757 B.n755 10.6151
R2231 B.n758 B.n757 10.6151
R2232 B.n759 B.n758 10.6151
R2233 B.n760 B.n759 10.6151
R2234 B.n762 B.n760 10.6151
R2235 B.n763 B.n762 10.6151
R2236 B.n764 B.n763 10.6151
R2237 B.n765 B.n764 10.6151
R2238 B.n767 B.n765 10.6151
R2239 B.n768 B.n767 10.6151
R2240 B.n769 B.n768 10.6151
R2241 B.n770 B.n769 10.6151
R2242 B.n772 B.n770 10.6151
R2243 B.n773 B.n772 10.6151
R2244 B.n774 B.n773 10.6151
R2245 B.n775 B.n774 10.6151
R2246 B.n777 B.n775 10.6151
R2247 B.n778 B.n777 10.6151
R2248 B.n779 B.n778 10.6151
R2249 B.n780 B.n779 10.6151
R2250 B.n782 B.n780 10.6151
R2251 B.n783 B.n782 10.6151
R2252 B.n784 B.n783 10.6151
R2253 B.n785 B.n784 10.6151
R2254 B.n787 B.n785 10.6151
R2255 B.n788 B.n787 10.6151
R2256 B.n437 B.n383 10.6151
R2257 B.n437 B.n436 10.6151
R2258 B.n443 B.n436 10.6151
R2259 B.n444 B.n443 10.6151
R2260 B.n445 B.n444 10.6151
R2261 B.n445 B.n434 10.6151
R2262 B.n451 B.n434 10.6151
R2263 B.n452 B.n451 10.6151
R2264 B.n453 B.n452 10.6151
R2265 B.n453 B.n432 10.6151
R2266 B.n459 B.n432 10.6151
R2267 B.n460 B.n459 10.6151
R2268 B.n461 B.n460 10.6151
R2269 B.n461 B.n430 10.6151
R2270 B.n467 B.n430 10.6151
R2271 B.n468 B.n467 10.6151
R2272 B.n469 B.n468 10.6151
R2273 B.n469 B.n428 10.6151
R2274 B.n475 B.n428 10.6151
R2275 B.n476 B.n475 10.6151
R2276 B.n477 B.n476 10.6151
R2277 B.n477 B.n426 10.6151
R2278 B.n483 B.n426 10.6151
R2279 B.n484 B.n483 10.6151
R2280 B.n485 B.n484 10.6151
R2281 B.n485 B.n424 10.6151
R2282 B.n491 B.n424 10.6151
R2283 B.n492 B.n491 10.6151
R2284 B.n493 B.n492 10.6151
R2285 B.n493 B.n422 10.6151
R2286 B.n499 B.n422 10.6151
R2287 B.n500 B.n499 10.6151
R2288 B.n501 B.n500 10.6151
R2289 B.n501 B.n420 10.6151
R2290 B.n507 B.n420 10.6151
R2291 B.n508 B.n507 10.6151
R2292 B.n509 B.n508 10.6151
R2293 B.n509 B.n418 10.6151
R2294 B.n515 B.n418 10.6151
R2295 B.n516 B.n515 10.6151
R2296 B.n517 B.n516 10.6151
R2297 B.n517 B.n416 10.6151
R2298 B.n523 B.n416 10.6151
R2299 B.n526 B.n525 10.6151
R2300 B.n526 B.n412 10.6151
R2301 B.n532 B.n412 10.6151
R2302 B.n533 B.n532 10.6151
R2303 B.n534 B.n533 10.6151
R2304 B.n534 B.n410 10.6151
R2305 B.n540 B.n410 10.6151
R2306 B.n541 B.n540 10.6151
R2307 B.n545 B.n541 10.6151
R2308 B.n551 B.n408 10.6151
R2309 B.n552 B.n551 10.6151
R2310 B.n553 B.n552 10.6151
R2311 B.n553 B.n406 10.6151
R2312 B.n559 B.n406 10.6151
R2313 B.n560 B.n559 10.6151
R2314 B.n561 B.n560 10.6151
R2315 B.n561 B.n404 10.6151
R2316 B.n567 B.n404 10.6151
R2317 B.n568 B.n567 10.6151
R2318 B.n569 B.n568 10.6151
R2319 B.n569 B.n402 10.6151
R2320 B.n575 B.n402 10.6151
R2321 B.n576 B.n575 10.6151
R2322 B.n577 B.n576 10.6151
R2323 B.n577 B.n400 10.6151
R2324 B.n583 B.n400 10.6151
R2325 B.n584 B.n583 10.6151
R2326 B.n585 B.n584 10.6151
R2327 B.n585 B.n398 10.6151
R2328 B.n591 B.n398 10.6151
R2329 B.n592 B.n591 10.6151
R2330 B.n593 B.n592 10.6151
R2331 B.n593 B.n396 10.6151
R2332 B.n599 B.n396 10.6151
R2333 B.n600 B.n599 10.6151
R2334 B.n601 B.n600 10.6151
R2335 B.n601 B.n394 10.6151
R2336 B.n607 B.n394 10.6151
R2337 B.n608 B.n607 10.6151
R2338 B.n609 B.n608 10.6151
R2339 B.n609 B.n392 10.6151
R2340 B.n615 B.n392 10.6151
R2341 B.n616 B.n615 10.6151
R2342 B.n617 B.n616 10.6151
R2343 B.n617 B.n390 10.6151
R2344 B.n623 B.n390 10.6151
R2345 B.n624 B.n623 10.6151
R2346 B.n625 B.n624 10.6151
R2347 B.n625 B.n388 10.6151
R2348 B.n388 B.n387 10.6151
R2349 B.n632 B.n387 10.6151
R2350 B.n633 B.n632 10.6151
R2351 B.n639 B.n638 10.6151
R2352 B.n640 B.n639 10.6151
R2353 B.n640 B.n375 10.6151
R2354 B.n650 B.n375 10.6151
R2355 B.n651 B.n650 10.6151
R2356 B.n652 B.n651 10.6151
R2357 B.n652 B.n367 10.6151
R2358 B.n662 B.n367 10.6151
R2359 B.n663 B.n662 10.6151
R2360 B.n664 B.n663 10.6151
R2361 B.n664 B.n359 10.6151
R2362 B.n674 B.n359 10.6151
R2363 B.n675 B.n674 10.6151
R2364 B.n676 B.n675 10.6151
R2365 B.n676 B.n351 10.6151
R2366 B.n686 B.n351 10.6151
R2367 B.n687 B.n686 10.6151
R2368 B.n688 B.n687 10.6151
R2369 B.n688 B.n343 10.6151
R2370 B.n698 B.n343 10.6151
R2371 B.n699 B.n698 10.6151
R2372 B.n700 B.n699 10.6151
R2373 B.n700 B.n335 10.6151
R2374 B.n710 B.n335 10.6151
R2375 B.n711 B.n710 10.6151
R2376 B.n712 B.n711 10.6151
R2377 B.n712 B.n327 10.6151
R2378 B.n722 B.n327 10.6151
R2379 B.n723 B.n722 10.6151
R2380 B.n724 B.n723 10.6151
R2381 B.n724 B.n319 10.6151
R2382 B.n735 B.n319 10.6151
R2383 B.n736 B.n735 10.6151
R2384 B.n737 B.n736 10.6151
R2385 B.n737 B.n0 10.6151
R2386 B.n861 B.n1 10.6151
R2387 B.n861 B.n860 10.6151
R2388 B.n860 B.n859 10.6151
R2389 B.n859 B.n10 10.6151
R2390 B.n853 B.n10 10.6151
R2391 B.n853 B.n852 10.6151
R2392 B.n852 B.n851 10.6151
R2393 B.n851 B.n17 10.6151
R2394 B.n845 B.n17 10.6151
R2395 B.n845 B.n844 10.6151
R2396 B.n844 B.n843 10.6151
R2397 B.n843 B.n24 10.6151
R2398 B.n837 B.n24 10.6151
R2399 B.n837 B.n836 10.6151
R2400 B.n836 B.n835 10.6151
R2401 B.n835 B.n31 10.6151
R2402 B.n829 B.n31 10.6151
R2403 B.n829 B.n828 10.6151
R2404 B.n828 B.n827 10.6151
R2405 B.n827 B.n38 10.6151
R2406 B.n821 B.n38 10.6151
R2407 B.n821 B.n820 10.6151
R2408 B.n820 B.n819 10.6151
R2409 B.n819 B.n45 10.6151
R2410 B.n813 B.n45 10.6151
R2411 B.n813 B.n812 10.6151
R2412 B.n812 B.n811 10.6151
R2413 B.n811 B.n52 10.6151
R2414 B.n805 B.n52 10.6151
R2415 B.n805 B.n804 10.6151
R2416 B.n804 B.n803 10.6151
R2417 B.n803 B.n59 10.6151
R2418 B.n797 B.n59 10.6151
R2419 B.n797 B.n796 10.6151
R2420 B.n796 B.n795 10.6151
R2421 B.n208 B.n123 9.36635
R2422 B.n231 B.n120 9.36635
R2423 B.n524 B.n523 9.36635
R2424 B.n544 B.n408 9.36635
R2425 B.t2 B.n353 6.67268
R2426 B.n824 B.t6 6.67268
R2427 B.n867 B.n0 2.81026
R2428 B.n867 B.n1 2.81026
R2429 B.n654 B.t9 1.82019
R2430 B.t13 B.n807 1.82019
R2431 B.n211 B.n123 1.24928
R2432 B.n228 B.n120 1.24928
R2433 B.n525 B.n524 1.24928
R2434 B.n545 B.n544 1.24928
R2435 B.n714 B.t3 0.607062
R2436 B.t0 B.n847 0.607062
R2437 VN.n4 VN.t3 228.359
R2438 VN.n25 VN.t5 228.359
R2439 VN.n5 VN.t4 197.405
R2440 VN.n12 VN.t6 197.405
R2441 VN.n19 VN.t2 197.405
R2442 VN.n26 VN.t7 197.405
R2443 VN.n33 VN.t0 197.405
R2444 VN.n40 VN.t1 197.405
R2445 VN.n20 VN.n19 180.974
R2446 VN.n41 VN.n40 180.974
R2447 VN.n39 VN.n21 161.3
R2448 VN.n38 VN.n37 161.3
R2449 VN.n36 VN.n22 161.3
R2450 VN.n35 VN.n34 161.3
R2451 VN.n32 VN.n23 161.3
R2452 VN.n31 VN.n30 161.3
R2453 VN.n29 VN.n24 161.3
R2454 VN.n28 VN.n27 161.3
R2455 VN.n18 VN.n0 161.3
R2456 VN.n17 VN.n16 161.3
R2457 VN.n15 VN.n1 161.3
R2458 VN.n14 VN.n13 161.3
R2459 VN.n11 VN.n2 161.3
R2460 VN.n10 VN.n9 161.3
R2461 VN.n8 VN.n3 161.3
R2462 VN.n7 VN.n6 161.3
R2463 VN.n5 VN.n4 56.6077
R2464 VN.n26 VN.n25 56.6077
R2465 VN.n10 VN.n3 56.5617
R2466 VN.n31 VN.n24 56.5617
R2467 VN.n17 VN.n1 55.1086
R2468 VN.n38 VN.n22 55.1086
R2469 VN VN.n41 46.9721
R2470 VN.n13 VN.n1 26.0455
R2471 VN.n34 VN.n22 26.0455
R2472 VN.n6 VN.n3 24.5923
R2473 VN.n11 VN.n10 24.5923
R2474 VN.n18 VN.n17 24.5923
R2475 VN.n27 VN.n24 24.5923
R2476 VN.n32 VN.n31 24.5923
R2477 VN.n39 VN.n38 24.5923
R2478 VN.n28 VN.n25 18.2882
R2479 VN.n7 VN.n4 18.2882
R2480 VN.n13 VN.n12 14.7556
R2481 VN.n34 VN.n33 14.7556
R2482 VN.n6 VN.n5 9.83723
R2483 VN.n12 VN.n11 9.83723
R2484 VN.n27 VN.n26 9.83723
R2485 VN.n33 VN.n32 9.83723
R2486 VN.n19 VN.n18 4.91887
R2487 VN.n40 VN.n39 4.91887
R2488 VN.n41 VN.n21 0.189894
R2489 VN.n37 VN.n21 0.189894
R2490 VN.n37 VN.n36 0.189894
R2491 VN.n36 VN.n35 0.189894
R2492 VN.n35 VN.n23 0.189894
R2493 VN.n30 VN.n23 0.189894
R2494 VN.n30 VN.n29 0.189894
R2495 VN.n29 VN.n28 0.189894
R2496 VN.n8 VN.n7 0.189894
R2497 VN.n9 VN.n8 0.189894
R2498 VN.n9 VN.n2 0.189894
R2499 VN.n14 VN.n2 0.189894
R2500 VN.n15 VN.n14 0.189894
R2501 VN.n16 VN.n15 0.189894
R2502 VN.n16 VN.n0 0.189894
R2503 VN.n20 VN.n0 0.189894
R2504 VN VN.n20 0.0516364
R2505 VDD2.n2 VDD2.n1 62.8548
R2506 VDD2.n2 VDD2.n0 62.8548
R2507 VDD2 VDD2.n5 62.8517
R2508 VDD2.n4 VDD2.n3 62.0911
R2509 VDD2.n4 VDD2.n2 42.1722
R2510 VDD2.n5 VDD2.t0 1.54016
R2511 VDD2.n5 VDD2.t2 1.54016
R2512 VDD2.n3 VDD2.t6 1.54016
R2513 VDD2.n3 VDD2.t7 1.54016
R2514 VDD2.n1 VDD2.t1 1.54016
R2515 VDD2.n1 VDD2.t5 1.54016
R2516 VDD2.n0 VDD2.t4 1.54016
R2517 VDD2.n0 VDD2.t3 1.54016
R2518 VDD2 VDD2.n4 0.877655
C0 VP VN 6.55981f
C1 VP VDD2 0.410401f
C2 VP VTAIL 8.231071f
C3 VP VDD1 8.44849f
C4 VN VTAIL 8.21696f
C5 VN VDD2 8.18916f
C6 VTAIL VDD2 8.824459f
C7 VN VDD1 0.150199f
C8 VTAIL VDD1 8.77695f
C9 VDD1 VDD2 1.25637f
C10 VDD2 B 4.410112f
C11 VDD1 B 4.73597f
C12 VTAIL B 10.209249f
C13 VN B 11.71205f
C14 VP B 10.093964f
C15 VDD2.t4 B 0.252932f
C16 VDD2.t3 B 0.252932f
C17 VDD2.n0 B 2.26808f
C18 VDD2.t1 B 0.252932f
C19 VDD2.t5 B 0.252932f
C20 VDD2.n1 B 2.26808f
C21 VDD2.n2 B 2.72475f
C22 VDD2.t6 B 0.252932f
C23 VDD2.t7 B 0.252932f
C24 VDD2.n3 B 2.2631f
C25 VDD2.n4 B 2.64876f
C26 VDD2.t0 B 0.252932f
C27 VDD2.t2 B 0.252932f
C28 VDD2.n5 B 2.26805f
C29 VN.n0 B 0.029987f
C30 VN.t2 B 1.65276f
C31 VN.n1 B 0.034086f
C32 VN.n2 B 0.029987f
C33 VN.t6 B 1.65276f
C34 VN.n3 B 0.043591f
C35 VN.t3 B 1.74921f
C36 VN.n4 B 0.668123f
C37 VN.t4 B 1.65276f
C38 VN.n5 B 0.647936f
C39 VN.n6 B 0.039137f
C40 VN.n7 B 0.188856f
C41 VN.n8 B 0.029987f
C42 VN.n9 B 0.029987f
C43 VN.n10 B 0.043591f
C44 VN.n11 B 0.039137f
C45 VN.n12 B 0.593031f
C46 VN.n13 B 0.046067f
C47 VN.n14 B 0.029987f
C48 VN.n15 B 0.029987f
C49 VN.n16 B 0.029987f
C50 VN.n17 B 0.051656f
C51 VN.n18 B 0.033646f
C52 VN.n19 B 0.650913f
C53 VN.n20 B 0.030299f
C54 VN.n21 B 0.029987f
C55 VN.t1 B 1.65276f
C56 VN.n22 B 0.034086f
C57 VN.n23 B 0.029987f
C58 VN.t0 B 1.65276f
C59 VN.n24 B 0.043591f
C60 VN.t5 B 1.74921f
C61 VN.n25 B 0.668123f
C62 VN.t7 B 1.65276f
C63 VN.n26 B 0.647936f
C64 VN.n27 B 0.039137f
C65 VN.n28 B 0.188856f
C66 VN.n29 B 0.029987f
C67 VN.n30 B 0.029987f
C68 VN.n31 B 0.043591f
C69 VN.n32 B 0.039137f
C70 VN.n33 B 0.593031f
C71 VN.n34 B 0.046067f
C72 VN.n35 B 0.029987f
C73 VN.n36 B 0.029987f
C74 VN.n37 B 0.029987f
C75 VN.n38 B 0.051656f
C76 VN.n39 B 0.033646f
C77 VN.n40 B 0.650913f
C78 VN.n41 B 1.48973f
C79 VTAIL.t0 B 0.193413f
C80 VTAIL.t7 B 0.193413f
C81 VTAIL.n0 B 1.67378f
C82 VTAIL.n1 B 0.293154f
C83 VTAIL.n2 B 0.027522f
C84 VTAIL.n3 B 0.019032f
C85 VTAIL.n4 B 0.010227f
C86 VTAIL.n5 B 0.024173f
C87 VTAIL.n6 B 0.010829f
C88 VTAIL.n7 B 0.019032f
C89 VTAIL.n8 B 0.010227f
C90 VTAIL.n9 B 0.024173f
C91 VTAIL.n10 B 0.010829f
C92 VTAIL.n11 B 0.019032f
C93 VTAIL.n12 B 0.010227f
C94 VTAIL.n13 B 0.024173f
C95 VTAIL.n14 B 0.010829f
C96 VTAIL.n15 B 0.019032f
C97 VTAIL.n16 B 0.010227f
C98 VTAIL.n17 B 0.024173f
C99 VTAIL.n18 B 0.010829f
C100 VTAIL.n19 B 0.019032f
C101 VTAIL.n20 B 0.010227f
C102 VTAIL.n21 B 0.024173f
C103 VTAIL.n22 B 0.010829f
C104 VTAIL.n23 B 0.143504f
C105 VTAIL.t4 B 0.040915f
C106 VTAIL.n24 B 0.01813f
C107 VTAIL.n25 B 0.017089f
C108 VTAIL.n26 B 0.010227f
C109 VTAIL.n27 B 1.03295f
C110 VTAIL.n28 B 0.019032f
C111 VTAIL.n29 B 0.010227f
C112 VTAIL.n30 B 0.010829f
C113 VTAIL.n31 B 0.024173f
C114 VTAIL.n32 B 0.024173f
C115 VTAIL.n33 B 0.010829f
C116 VTAIL.n34 B 0.010227f
C117 VTAIL.n35 B 0.019032f
C118 VTAIL.n36 B 0.019032f
C119 VTAIL.n37 B 0.010227f
C120 VTAIL.n38 B 0.010829f
C121 VTAIL.n39 B 0.024173f
C122 VTAIL.n40 B 0.024173f
C123 VTAIL.n41 B 0.024173f
C124 VTAIL.n42 B 0.010829f
C125 VTAIL.n43 B 0.010227f
C126 VTAIL.n44 B 0.019032f
C127 VTAIL.n45 B 0.019032f
C128 VTAIL.n46 B 0.010227f
C129 VTAIL.n47 B 0.010528f
C130 VTAIL.n48 B 0.010528f
C131 VTAIL.n49 B 0.024173f
C132 VTAIL.n50 B 0.024173f
C133 VTAIL.n51 B 0.010829f
C134 VTAIL.n52 B 0.010227f
C135 VTAIL.n53 B 0.019032f
C136 VTAIL.n54 B 0.019032f
C137 VTAIL.n55 B 0.010227f
C138 VTAIL.n56 B 0.010829f
C139 VTAIL.n57 B 0.024173f
C140 VTAIL.n58 B 0.024173f
C141 VTAIL.n59 B 0.010829f
C142 VTAIL.n60 B 0.010227f
C143 VTAIL.n61 B 0.019032f
C144 VTAIL.n62 B 0.019032f
C145 VTAIL.n63 B 0.010227f
C146 VTAIL.n64 B 0.010829f
C147 VTAIL.n65 B 0.024173f
C148 VTAIL.n66 B 0.053693f
C149 VTAIL.n67 B 0.010829f
C150 VTAIL.n68 B 0.010227f
C151 VTAIL.n69 B 0.044512f
C152 VTAIL.n70 B 0.030199f
C153 VTAIL.n71 B 0.145809f
C154 VTAIL.n72 B 0.027522f
C155 VTAIL.n73 B 0.019032f
C156 VTAIL.n74 B 0.010227f
C157 VTAIL.n75 B 0.024173f
C158 VTAIL.n76 B 0.010829f
C159 VTAIL.n77 B 0.019032f
C160 VTAIL.n78 B 0.010227f
C161 VTAIL.n79 B 0.024173f
C162 VTAIL.n80 B 0.010829f
C163 VTAIL.n81 B 0.019032f
C164 VTAIL.n82 B 0.010227f
C165 VTAIL.n83 B 0.024173f
C166 VTAIL.n84 B 0.010829f
C167 VTAIL.n85 B 0.019032f
C168 VTAIL.n86 B 0.010227f
C169 VTAIL.n87 B 0.024173f
C170 VTAIL.n88 B 0.010829f
C171 VTAIL.n89 B 0.019032f
C172 VTAIL.n90 B 0.010227f
C173 VTAIL.n91 B 0.024173f
C174 VTAIL.n92 B 0.010829f
C175 VTAIL.n93 B 0.143504f
C176 VTAIL.t9 B 0.040915f
C177 VTAIL.n94 B 0.01813f
C178 VTAIL.n95 B 0.017089f
C179 VTAIL.n96 B 0.010227f
C180 VTAIL.n97 B 1.03295f
C181 VTAIL.n98 B 0.019032f
C182 VTAIL.n99 B 0.010227f
C183 VTAIL.n100 B 0.010829f
C184 VTAIL.n101 B 0.024173f
C185 VTAIL.n102 B 0.024173f
C186 VTAIL.n103 B 0.010829f
C187 VTAIL.n104 B 0.010227f
C188 VTAIL.n105 B 0.019032f
C189 VTAIL.n106 B 0.019032f
C190 VTAIL.n107 B 0.010227f
C191 VTAIL.n108 B 0.010829f
C192 VTAIL.n109 B 0.024173f
C193 VTAIL.n110 B 0.024173f
C194 VTAIL.n111 B 0.024173f
C195 VTAIL.n112 B 0.010829f
C196 VTAIL.n113 B 0.010227f
C197 VTAIL.n114 B 0.019032f
C198 VTAIL.n115 B 0.019032f
C199 VTAIL.n116 B 0.010227f
C200 VTAIL.n117 B 0.010528f
C201 VTAIL.n118 B 0.010528f
C202 VTAIL.n119 B 0.024173f
C203 VTAIL.n120 B 0.024173f
C204 VTAIL.n121 B 0.010829f
C205 VTAIL.n122 B 0.010227f
C206 VTAIL.n123 B 0.019032f
C207 VTAIL.n124 B 0.019032f
C208 VTAIL.n125 B 0.010227f
C209 VTAIL.n126 B 0.010829f
C210 VTAIL.n127 B 0.024173f
C211 VTAIL.n128 B 0.024173f
C212 VTAIL.n129 B 0.010829f
C213 VTAIL.n130 B 0.010227f
C214 VTAIL.n131 B 0.019032f
C215 VTAIL.n132 B 0.019032f
C216 VTAIL.n133 B 0.010227f
C217 VTAIL.n134 B 0.010829f
C218 VTAIL.n135 B 0.024173f
C219 VTAIL.n136 B 0.053693f
C220 VTAIL.n137 B 0.010829f
C221 VTAIL.n138 B 0.010227f
C222 VTAIL.n139 B 0.044512f
C223 VTAIL.n140 B 0.030199f
C224 VTAIL.n141 B 0.145809f
C225 VTAIL.t14 B 0.193413f
C226 VTAIL.t8 B 0.193413f
C227 VTAIL.n142 B 1.67378f
C228 VTAIL.n143 B 0.390033f
C229 VTAIL.n144 B 0.027522f
C230 VTAIL.n145 B 0.019032f
C231 VTAIL.n146 B 0.010227f
C232 VTAIL.n147 B 0.024173f
C233 VTAIL.n148 B 0.010829f
C234 VTAIL.n149 B 0.019032f
C235 VTAIL.n150 B 0.010227f
C236 VTAIL.n151 B 0.024173f
C237 VTAIL.n152 B 0.010829f
C238 VTAIL.n153 B 0.019032f
C239 VTAIL.n154 B 0.010227f
C240 VTAIL.n155 B 0.024173f
C241 VTAIL.n156 B 0.010829f
C242 VTAIL.n157 B 0.019032f
C243 VTAIL.n158 B 0.010227f
C244 VTAIL.n159 B 0.024173f
C245 VTAIL.n160 B 0.010829f
C246 VTAIL.n161 B 0.019032f
C247 VTAIL.n162 B 0.010227f
C248 VTAIL.n163 B 0.024173f
C249 VTAIL.n164 B 0.010829f
C250 VTAIL.n165 B 0.143504f
C251 VTAIL.t11 B 0.040915f
C252 VTAIL.n166 B 0.01813f
C253 VTAIL.n167 B 0.017089f
C254 VTAIL.n168 B 0.010227f
C255 VTAIL.n169 B 1.03295f
C256 VTAIL.n170 B 0.019032f
C257 VTAIL.n171 B 0.010227f
C258 VTAIL.n172 B 0.010829f
C259 VTAIL.n173 B 0.024173f
C260 VTAIL.n174 B 0.024173f
C261 VTAIL.n175 B 0.010829f
C262 VTAIL.n176 B 0.010227f
C263 VTAIL.n177 B 0.019032f
C264 VTAIL.n178 B 0.019032f
C265 VTAIL.n179 B 0.010227f
C266 VTAIL.n180 B 0.010829f
C267 VTAIL.n181 B 0.024173f
C268 VTAIL.n182 B 0.024173f
C269 VTAIL.n183 B 0.024173f
C270 VTAIL.n184 B 0.010829f
C271 VTAIL.n185 B 0.010227f
C272 VTAIL.n186 B 0.019032f
C273 VTAIL.n187 B 0.019032f
C274 VTAIL.n188 B 0.010227f
C275 VTAIL.n189 B 0.010528f
C276 VTAIL.n190 B 0.010528f
C277 VTAIL.n191 B 0.024173f
C278 VTAIL.n192 B 0.024173f
C279 VTAIL.n193 B 0.010829f
C280 VTAIL.n194 B 0.010227f
C281 VTAIL.n195 B 0.019032f
C282 VTAIL.n196 B 0.019032f
C283 VTAIL.n197 B 0.010227f
C284 VTAIL.n198 B 0.010829f
C285 VTAIL.n199 B 0.024173f
C286 VTAIL.n200 B 0.024173f
C287 VTAIL.n201 B 0.010829f
C288 VTAIL.n202 B 0.010227f
C289 VTAIL.n203 B 0.019032f
C290 VTAIL.n204 B 0.019032f
C291 VTAIL.n205 B 0.010227f
C292 VTAIL.n206 B 0.010829f
C293 VTAIL.n207 B 0.024173f
C294 VTAIL.n208 B 0.053693f
C295 VTAIL.n209 B 0.010829f
C296 VTAIL.n210 B 0.010227f
C297 VTAIL.n211 B 0.044512f
C298 VTAIL.n212 B 0.030199f
C299 VTAIL.n213 B 1.15585f
C300 VTAIL.n214 B 0.027522f
C301 VTAIL.n215 B 0.019032f
C302 VTAIL.n216 B 0.010227f
C303 VTAIL.n217 B 0.024173f
C304 VTAIL.n218 B 0.010829f
C305 VTAIL.n219 B 0.019032f
C306 VTAIL.n220 B 0.010227f
C307 VTAIL.n221 B 0.024173f
C308 VTAIL.n222 B 0.010829f
C309 VTAIL.n223 B 0.019032f
C310 VTAIL.n224 B 0.010227f
C311 VTAIL.n225 B 0.024173f
C312 VTAIL.n226 B 0.010829f
C313 VTAIL.n227 B 0.019032f
C314 VTAIL.n228 B 0.010227f
C315 VTAIL.n229 B 0.024173f
C316 VTAIL.n230 B 0.024173f
C317 VTAIL.n231 B 0.010829f
C318 VTAIL.n232 B 0.019032f
C319 VTAIL.n233 B 0.010227f
C320 VTAIL.n234 B 0.024173f
C321 VTAIL.n235 B 0.010829f
C322 VTAIL.n236 B 0.143504f
C323 VTAIL.t2 B 0.040915f
C324 VTAIL.n237 B 0.01813f
C325 VTAIL.n238 B 0.017089f
C326 VTAIL.n239 B 0.010227f
C327 VTAIL.n240 B 1.03295f
C328 VTAIL.n241 B 0.019032f
C329 VTAIL.n242 B 0.010227f
C330 VTAIL.n243 B 0.010829f
C331 VTAIL.n244 B 0.024173f
C332 VTAIL.n245 B 0.024173f
C333 VTAIL.n246 B 0.010829f
C334 VTAIL.n247 B 0.010227f
C335 VTAIL.n248 B 0.019032f
C336 VTAIL.n249 B 0.019032f
C337 VTAIL.n250 B 0.010227f
C338 VTAIL.n251 B 0.010829f
C339 VTAIL.n252 B 0.024173f
C340 VTAIL.n253 B 0.024173f
C341 VTAIL.n254 B 0.010829f
C342 VTAIL.n255 B 0.010227f
C343 VTAIL.n256 B 0.019032f
C344 VTAIL.n257 B 0.019032f
C345 VTAIL.n258 B 0.010227f
C346 VTAIL.n259 B 0.010528f
C347 VTAIL.n260 B 0.010528f
C348 VTAIL.n261 B 0.024173f
C349 VTAIL.n262 B 0.024173f
C350 VTAIL.n263 B 0.010829f
C351 VTAIL.n264 B 0.010227f
C352 VTAIL.n265 B 0.019032f
C353 VTAIL.n266 B 0.019032f
C354 VTAIL.n267 B 0.010227f
C355 VTAIL.n268 B 0.010829f
C356 VTAIL.n269 B 0.024173f
C357 VTAIL.n270 B 0.024173f
C358 VTAIL.n271 B 0.010829f
C359 VTAIL.n272 B 0.010227f
C360 VTAIL.n273 B 0.019032f
C361 VTAIL.n274 B 0.019032f
C362 VTAIL.n275 B 0.010227f
C363 VTAIL.n276 B 0.010829f
C364 VTAIL.n277 B 0.024173f
C365 VTAIL.n278 B 0.053693f
C366 VTAIL.n279 B 0.010829f
C367 VTAIL.n280 B 0.010227f
C368 VTAIL.n281 B 0.044512f
C369 VTAIL.n282 B 0.030199f
C370 VTAIL.n283 B 1.15585f
C371 VTAIL.t1 B 0.193413f
C372 VTAIL.t3 B 0.193413f
C373 VTAIL.n284 B 1.67378f
C374 VTAIL.n285 B 0.390031f
C375 VTAIL.n286 B 0.027522f
C376 VTAIL.n287 B 0.019032f
C377 VTAIL.n288 B 0.010227f
C378 VTAIL.n289 B 0.024173f
C379 VTAIL.n290 B 0.010829f
C380 VTAIL.n291 B 0.019032f
C381 VTAIL.n292 B 0.010227f
C382 VTAIL.n293 B 0.024173f
C383 VTAIL.n294 B 0.010829f
C384 VTAIL.n295 B 0.019032f
C385 VTAIL.n296 B 0.010227f
C386 VTAIL.n297 B 0.024173f
C387 VTAIL.n298 B 0.010829f
C388 VTAIL.n299 B 0.019032f
C389 VTAIL.n300 B 0.010227f
C390 VTAIL.n301 B 0.024173f
C391 VTAIL.n302 B 0.024173f
C392 VTAIL.n303 B 0.010829f
C393 VTAIL.n304 B 0.019032f
C394 VTAIL.n305 B 0.010227f
C395 VTAIL.n306 B 0.024173f
C396 VTAIL.n307 B 0.010829f
C397 VTAIL.n308 B 0.143504f
C398 VTAIL.t5 B 0.040915f
C399 VTAIL.n309 B 0.01813f
C400 VTAIL.n310 B 0.017089f
C401 VTAIL.n311 B 0.010227f
C402 VTAIL.n312 B 1.03295f
C403 VTAIL.n313 B 0.019032f
C404 VTAIL.n314 B 0.010227f
C405 VTAIL.n315 B 0.010829f
C406 VTAIL.n316 B 0.024173f
C407 VTAIL.n317 B 0.024173f
C408 VTAIL.n318 B 0.010829f
C409 VTAIL.n319 B 0.010227f
C410 VTAIL.n320 B 0.019032f
C411 VTAIL.n321 B 0.019032f
C412 VTAIL.n322 B 0.010227f
C413 VTAIL.n323 B 0.010829f
C414 VTAIL.n324 B 0.024173f
C415 VTAIL.n325 B 0.024173f
C416 VTAIL.n326 B 0.010829f
C417 VTAIL.n327 B 0.010227f
C418 VTAIL.n328 B 0.019032f
C419 VTAIL.n329 B 0.019032f
C420 VTAIL.n330 B 0.010227f
C421 VTAIL.n331 B 0.010528f
C422 VTAIL.n332 B 0.010528f
C423 VTAIL.n333 B 0.024173f
C424 VTAIL.n334 B 0.024173f
C425 VTAIL.n335 B 0.010829f
C426 VTAIL.n336 B 0.010227f
C427 VTAIL.n337 B 0.019032f
C428 VTAIL.n338 B 0.019032f
C429 VTAIL.n339 B 0.010227f
C430 VTAIL.n340 B 0.010829f
C431 VTAIL.n341 B 0.024173f
C432 VTAIL.n342 B 0.024173f
C433 VTAIL.n343 B 0.010829f
C434 VTAIL.n344 B 0.010227f
C435 VTAIL.n345 B 0.019032f
C436 VTAIL.n346 B 0.019032f
C437 VTAIL.n347 B 0.010227f
C438 VTAIL.n348 B 0.010829f
C439 VTAIL.n349 B 0.024173f
C440 VTAIL.n350 B 0.053693f
C441 VTAIL.n351 B 0.010829f
C442 VTAIL.n352 B 0.010227f
C443 VTAIL.n353 B 0.044512f
C444 VTAIL.n354 B 0.030199f
C445 VTAIL.n355 B 0.145809f
C446 VTAIL.n356 B 0.027522f
C447 VTAIL.n357 B 0.019032f
C448 VTAIL.n358 B 0.010227f
C449 VTAIL.n359 B 0.024173f
C450 VTAIL.n360 B 0.010829f
C451 VTAIL.n361 B 0.019032f
C452 VTAIL.n362 B 0.010227f
C453 VTAIL.n363 B 0.024173f
C454 VTAIL.n364 B 0.010829f
C455 VTAIL.n365 B 0.019032f
C456 VTAIL.n366 B 0.010227f
C457 VTAIL.n367 B 0.024173f
C458 VTAIL.n368 B 0.010829f
C459 VTAIL.n369 B 0.019032f
C460 VTAIL.n370 B 0.010227f
C461 VTAIL.n371 B 0.024173f
C462 VTAIL.n372 B 0.024173f
C463 VTAIL.n373 B 0.010829f
C464 VTAIL.n374 B 0.019032f
C465 VTAIL.n375 B 0.010227f
C466 VTAIL.n376 B 0.024173f
C467 VTAIL.n377 B 0.010829f
C468 VTAIL.n378 B 0.143504f
C469 VTAIL.t15 B 0.040915f
C470 VTAIL.n379 B 0.01813f
C471 VTAIL.n380 B 0.017089f
C472 VTAIL.n381 B 0.010227f
C473 VTAIL.n382 B 1.03295f
C474 VTAIL.n383 B 0.019032f
C475 VTAIL.n384 B 0.010227f
C476 VTAIL.n385 B 0.010829f
C477 VTAIL.n386 B 0.024173f
C478 VTAIL.n387 B 0.024173f
C479 VTAIL.n388 B 0.010829f
C480 VTAIL.n389 B 0.010227f
C481 VTAIL.n390 B 0.019032f
C482 VTAIL.n391 B 0.019032f
C483 VTAIL.n392 B 0.010227f
C484 VTAIL.n393 B 0.010829f
C485 VTAIL.n394 B 0.024173f
C486 VTAIL.n395 B 0.024173f
C487 VTAIL.n396 B 0.010829f
C488 VTAIL.n397 B 0.010227f
C489 VTAIL.n398 B 0.019032f
C490 VTAIL.n399 B 0.019032f
C491 VTAIL.n400 B 0.010227f
C492 VTAIL.n401 B 0.010528f
C493 VTAIL.n402 B 0.010528f
C494 VTAIL.n403 B 0.024173f
C495 VTAIL.n404 B 0.024173f
C496 VTAIL.n405 B 0.010829f
C497 VTAIL.n406 B 0.010227f
C498 VTAIL.n407 B 0.019032f
C499 VTAIL.n408 B 0.019032f
C500 VTAIL.n409 B 0.010227f
C501 VTAIL.n410 B 0.010829f
C502 VTAIL.n411 B 0.024173f
C503 VTAIL.n412 B 0.024173f
C504 VTAIL.n413 B 0.010829f
C505 VTAIL.n414 B 0.010227f
C506 VTAIL.n415 B 0.019032f
C507 VTAIL.n416 B 0.019032f
C508 VTAIL.n417 B 0.010227f
C509 VTAIL.n418 B 0.010829f
C510 VTAIL.n419 B 0.024173f
C511 VTAIL.n420 B 0.053693f
C512 VTAIL.n421 B 0.010829f
C513 VTAIL.n422 B 0.010227f
C514 VTAIL.n423 B 0.044512f
C515 VTAIL.n424 B 0.030199f
C516 VTAIL.n425 B 0.145809f
C517 VTAIL.t13 B 0.193413f
C518 VTAIL.t12 B 0.193413f
C519 VTAIL.n426 B 1.67378f
C520 VTAIL.n427 B 0.390031f
C521 VTAIL.n428 B 0.027522f
C522 VTAIL.n429 B 0.019032f
C523 VTAIL.n430 B 0.010227f
C524 VTAIL.n431 B 0.024173f
C525 VTAIL.n432 B 0.010829f
C526 VTAIL.n433 B 0.019032f
C527 VTAIL.n434 B 0.010227f
C528 VTAIL.n435 B 0.024173f
C529 VTAIL.n436 B 0.010829f
C530 VTAIL.n437 B 0.019032f
C531 VTAIL.n438 B 0.010227f
C532 VTAIL.n439 B 0.024173f
C533 VTAIL.n440 B 0.010829f
C534 VTAIL.n441 B 0.019032f
C535 VTAIL.n442 B 0.010227f
C536 VTAIL.n443 B 0.024173f
C537 VTAIL.n444 B 0.024173f
C538 VTAIL.n445 B 0.010829f
C539 VTAIL.n446 B 0.019032f
C540 VTAIL.n447 B 0.010227f
C541 VTAIL.n448 B 0.024173f
C542 VTAIL.n449 B 0.010829f
C543 VTAIL.n450 B 0.143504f
C544 VTAIL.t10 B 0.040915f
C545 VTAIL.n451 B 0.01813f
C546 VTAIL.n452 B 0.017089f
C547 VTAIL.n453 B 0.010227f
C548 VTAIL.n454 B 1.03295f
C549 VTAIL.n455 B 0.019032f
C550 VTAIL.n456 B 0.010227f
C551 VTAIL.n457 B 0.010829f
C552 VTAIL.n458 B 0.024173f
C553 VTAIL.n459 B 0.024173f
C554 VTAIL.n460 B 0.010829f
C555 VTAIL.n461 B 0.010227f
C556 VTAIL.n462 B 0.019032f
C557 VTAIL.n463 B 0.019032f
C558 VTAIL.n464 B 0.010227f
C559 VTAIL.n465 B 0.010829f
C560 VTAIL.n466 B 0.024173f
C561 VTAIL.n467 B 0.024173f
C562 VTAIL.n468 B 0.010829f
C563 VTAIL.n469 B 0.010227f
C564 VTAIL.n470 B 0.019032f
C565 VTAIL.n471 B 0.019032f
C566 VTAIL.n472 B 0.010227f
C567 VTAIL.n473 B 0.010528f
C568 VTAIL.n474 B 0.010528f
C569 VTAIL.n475 B 0.024173f
C570 VTAIL.n476 B 0.024173f
C571 VTAIL.n477 B 0.010829f
C572 VTAIL.n478 B 0.010227f
C573 VTAIL.n479 B 0.019032f
C574 VTAIL.n480 B 0.019032f
C575 VTAIL.n481 B 0.010227f
C576 VTAIL.n482 B 0.010829f
C577 VTAIL.n483 B 0.024173f
C578 VTAIL.n484 B 0.024173f
C579 VTAIL.n485 B 0.010829f
C580 VTAIL.n486 B 0.010227f
C581 VTAIL.n487 B 0.019032f
C582 VTAIL.n488 B 0.019032f
C583 VTAIL.n489 B 0.010227f
C584 VTAIL.n490 B 0.010829f
C585 VTAIL.n491 B 0.024173f
C586 VTAIL.n492 B 0.053693f
C587 VTAIL.n493 B 0.010829f
C588 VTAIL.n494 B 0.010227f
C589 VTAIL.n495 B 0.044512f
C590 VTAIL.n496 B 0.030199f
C591 VTAIL.n497 B 1.15585f
C592 VTAIL.n498 B 0.027522f
C593 VTAIL.n499 B 0.019032f
C594 VTAIL.n500 B 0.010227f
C595 VTAIL.n501 B 0.024173f
C596 VTAIL.n502 B 0.010829f
C597 VTAIL.n503 B 0.019032f
C598 VTAIL.n504 B 0.010227f
C599 VTAIL.n505 B 0.024173f
C600 VTAIL.n506 B 0.010829f
C601 VTAIL.n507 B 0.019032f
C602 VTAIL.n508 B 0.010227f
C603 VTAIL.n509 B 0.024173f
C604 VTAIL.n510 B 0.010829f
C605 VTAIL.n511 B 0.019032f
C606 VTAIL.n512 B 0.010227f
C607 VTAIL.n513 B 0.024173f
C608 VTAIL.n514 B 0.010829f
C609 VTAIL.n515 B 0.019032f
C610 VTAIL.n516 B 0.010227f
C611 VTAIL.n517 B 0.024173f
C612 VTAIL.n518 B 0.010829f
C613 VTAIL.n519 B 0.143504f
C614 VTAIL.t6 B 0.040915f
C615 VTAIL.n520 B 0.01813f
C616 VTAIL.n521 B 0.017089f
C617 VTAIL.n522 B 0.010227f
C618 VTAIL.n523 B 1.03295f
C619 VTAIL.n524 B 0.019032f
C620 VTAIL.n525 B 0.010227f
C621 VTAIL.n526 B 0.010829f
C622 VTAIL.n527 B 0.024173f
C623 VTAIL.n528 B 0.024173f
C624 VTAIL.n529 B 0.010829f
C625 VTAIL.n530 B 0.010227f
C626 VTAIL.n531 B 0.019032f
C627 VTAIL.n532 B 0.019032f
C628 VTAIL.n533 B 0.010227f
C629 VTAIL.n534 B 0.010829f
C630 VTAIL.n535 B 0.024173f
C631 VTAIL.n536 B 0.024173f
C632 VTAIL.n537 B 0.024173f
C633 VTAIL.n538 B 0.010829f
C634 VTAIL.n539 B 0.010227f
C635 VTAIL.n540 B 0.019032f
C636 VTAIL.n541 B 0.019032f
C637 VTAIL.n542 B 0.010227f
C638 VTAIL.n543 B 0.010528f
C639 VTAIL.n544 B 0.010528f
C640 VTAIL.n545 B 0.024173f
C641 VTAIL.n546 B 0.024173f
C642 VTAIL.n547 B 0.010829f
C643 VTAIL.n548 B 0.010227f
C644 VTAIL.n549 B 0.019032f
C645 VTAIL.n550 B 0.019032f
C646 VTAIL.n551 B 0.010227f
C647 VTAIL.n552 B 0.010829f
C648 VTAIL.n553 B 0.024173f
C649 VTAIL.n554 B 0.024173f
C650 VTAIL.n555 B 0.010829f
C651 VTAIL.n556 B 0.010227f
C652 VTAIL.n557 B 0.019032f
C653 VTAIL.n558 B 0.019032f
C654 VTAIL.n559 B 0.010227f
C655 VTAIL.n560 B 0.010829f
C656 VTAIL.n561 B 0.024173f
C657 VTAIL.n562 B 0.053693f
C658 VTAIL.n563 B 0.010829f
C659 VTAIL.n564 B 0.010227f
C660 VTAIL.n565 B 0.044512f
C661 VTAIL.n566 B 0.030199f
C662 VTAIL.n567 B 1.15228f
C663 VDD1.t4 B 0.254531f
C664 VDD1.t5 B 0.254531f
C665 VDD1.n0 B 2.28328f
C666 VDD1.t6 B 0.254531f
C667 VDD1.t3 B 0.254531f
C668 VDD1.n1 B 2.28243f
C669 VDD1.t1 B 0.254531f
C670 VDD1.t0 B 0.254531f
C671 VDD1.n2 B 2.28243f
C672 VDD1.n3 B 2.79474f
C673 VDD1.t7 B 0.254531f
C674 VDD1.t2 B 0.254531f
C675 VDD1.n4 B 2.2774f
C676 VDD1.n5 B 2.69587f
C677 VP.n0 B 0.030303f
C678 VP.t6 B 1.67019f
C679 VP.n1 B 0.034446f
C680 VP.n2 B 0.030303f
C681 VP.t7 B 1.67019f
C682 VP.n3 B 0.04405f
C683 VP.n4 B 0.030303f
C684 VP.t1 B 1.67019f
C685 VP.n5 B 0.0522f
C686 VP.n6 B 0.030303f
C687 VP.t5 B 1.67019f
C688 VP.n7 B 0.034446f
C689 VP.n8 B 0.030303f
C690 VP.t3 B 1.67019f
C691 VP.n9 B 0.04405f
C692 VP.t0 B 1.76766f
C693 VP.n10 B 0.67517f
C694 VP.t2 B 1.67019f
C695 VP.n11 B 0.65477f
C696 VP.n12 B 0.039549f
C697 VP.n13 B 0.190848f
C698 VP.n14 B 0.030303f
C699 VP.n15 B 0.030303f
C700 VP.n16 B 0.04405f
C701 VP.n17 B 0.039549f
C702 VP.n18 B 0.599286f
C703 VP.n19 B 0.046553f
C704 VP.n20 B 0.030303f
C705 VP.n21 B 0.030303f
C706 VP.n22 B 0.030303f
C707 VP.n23 B 0.0522f
C708 VP.n24 B 0.034001f
C709 VP.n25 B 0.657779f
C710 VP.n26 B 1.48567f
C711 VP.n27 B 1.50912f
C712 VP.t4 B 1.67019f
C713 VP.n28 B 0.657779f
C714 VP.n29 B 0.034001f
C715 VP.n30 B 0.030303f
C716 VP.n31 B 0.030303f
C717 VP.n32 B 0.030303f
C718 VP.n33 B 0.034446f
C719 VP.n34 B 0.046553f
C720 VP.n35 B 0.599286f
C721 VP.n36 B 0.039549f
C722 VP.n37 B 0.030303f
C723 VP.n38 B 0.030303f
C724 VP.n39 B 0.030303f
C725 VP.n40 B 0.04405f
C726 VP.n41 B 0.039549f
C727 VP.n42 B 0.599286f
C728 VP.n43 B 0.046553f
C729 VP.n44 B 0.030303f
C730 VP.n45 B 0.030303f
C731 VP.n46 B 0.030303f
C732 VP.n47 B 0.0522f
C733 VP.n48 B 0.034001f
C734 VP.n49 B 0.657779f
C735 VP.n50 B 0.030618f
.ends

