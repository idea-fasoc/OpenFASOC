* NGSPICE file created from diff_pair_sample_0780.ext - technology: sky130A

.subckt diff_pair_sample_0780 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t11 VP.t0 VDD1.t1 w_n2514_n4224# sky130_fd_pr__pfet_01v8 ad=2.6862 pd=16.61 as=2.6862 ps=16.61 w=16.28 l=1.6
X1 VDD2.t5 VN.t0 VTAIL.t3 w_n2514_n4224# sky130_fd_pr__pfet_01v8 ad=6.3492 pd=33.34 as=2.6862 ps=16.61 w=16.28 l=1.6
X2 B.t11 B.t9 B.t10 w_n2514_n4224# sky130_fd_pr__pfet_01v8 ad=6.3492 pd=33.34 as=0 ps=0 w=16.28 l=1.6
X3 VDD1.t0 VP.t1 VTAIL.t10 w_n2514_n4224# sky130_fd_pr__pfet_01v8 ad=6.3492 pd=33.34 as=2.6862 ps=16.61 w=16.28 l=1.6
X4 VTAIL.t9 VP.t2 VDD1.t4 w_n2514_n4224# sky130_fd_pr__pfet_01v8 ad=2.6862 pd=16.61 as=2.6862 ps=16.61 w=16.28 l=1.6
X5 B.t8 B.t6 B.t7 w_n2514_n4224# sky130_fd_pr__pfet_01v8 ad=6.3492 pd=33.34 as=0 ps=0 w=16.28 l=1.6
X6 VDD2.t4 VN.t1 VTAIL.t1 w_n2514_n4224# sky130_fd_pr__pfet_01v8 ad=6.3492 pd=33.34 as=2.6862 ps=16.61 w=16.28 l=1.6
X7 VDD2.t3 VN.t2 VTAIL.t5 w_n2514_n4224# sky130_fd_pr__pfet_01v8 ad=2.6862 pd=16.61 as=6.3492 ps=33.34 w=16.28 l=1.6
X8 B.t5 B.t3 B.t4 w_n2514_n4224# sky130_fd_pr__pfet_01v8 ad=6.3492 pd=33.34 as=0 ps=0 w=16.28 l=1.6
X9 VDD1.t2 VP.t3 VTAIL.t8 w_n2514_n4224# sky130_fd_pr__pfet_01v8 ad=2.6862 pd=16.61 as=6.3492 ps=33.34 w=16.28 l=1.6
X10 VTAIL.t0 VN.t3 VDD2.t2 w_n2514_n4224# sky130_fd_pr__pfet_01v8 ad=2.6862 pd=16.61 as=2.6862 ps=16.61 w=16.28 l=1.6
X11 VDD2.t1 VN.t4 VTAIL.t2 w_n2514_n4224# sky130_fd_pr__pfet_01v8 ad=2.6862 pd=16.61 as=6.3492 ps=33.34 w=16.28 l=1.6
X12 VTAIL.t4 VN.t5 VDD2.t0 w_n2514_n4224# sky130_fd_pr__pfet_01v8 ad=2.6862 pd=16.61 as=2.6862 ps=16.61 w=16.28 l=1.6
X13 VDD1.t5 VP.t4 VTAIL.t7 w_n2514_n4224# sky130_fd_pr__pfet_01v8 ad=2.6862 pd=16.61 as=6.3492 ps=33.34 w=16.28 l=1.6
X14 VDD1.t3 VP.t5 VTAIL.t6 w_n2514_n4224# sky130_fd_pr__pfet_01v8 ad=6.3492 pd=33.34 as=2.6862 ps=16.61 w=16.28 l=1.6
X15 B.t2 B.t0 B.t1 w_n2514_n4224# sky130_fd_pr__pfet_01v8 ad=6.3492 pd=33.34 as=0 ps=0 w=16.28 l=1.6
R0 VP.n6 VP.t5 278.24
R1 VP.n17 VP.t1 245.218
R2 VP.n24 VP.t0 245.218
R3 VP.n31 VP.t4 245.218
R4 VP.n14 VP.t3 245.218
R5 VP.n7 VP.t2 245.218
R6 VP.n17 VP.n16 176.881
R7 VP.n32 VP.n31 176.881
R8 VP.n15 VP.n14 176.881
R9 VP.n9 VP.n8 161.3
R10 VP.n10 VP.n5 161.3
R11 VP.n12 VP.n11 161.3
R12 VP.n13 VP.n4 161.3
R13 VP.n30 VP.n0 161.3
R14 VP.n29 VP.n28 161.3
R15 VP.n27 VP.n1 161.3
R16 VP.n26 VP.n25 161.3
R17 VP.n23 VP.n2 161.3
R18 VP.n22 VP.n21 161.3
R19 VP.n20 VP.n3 161.3
R20 VP.n19 VP.n18 161.3
R21 VP.n22 VP.n3 56.4773
R22 VP.n29 VP.n1 56.4773
R23 VP.n12 VP.n5 56.4773
R24 VP.n7 VP.n6 53.8729
R25 VP.n16 VP.n15 47.9285
R26 VP.n18 VP.n3 24.3439
R27 VP.n23 VP.n22 24.3439
R28 VP.n25 VP.n1 24.3439
R29 VP.n30 VP.n29 24.3439
R30 VP.n13 VP.n12 24.3439
R31 VP.n8 VP.n5 24.3439
R32 VP.n9 VP.n6 17.9272
R33 VP.n24 VP.n23 12.1722
R34 VP.n25 VP.n24 12.1722
R35 VP.n8 VP.n7 12.1722
R36 VP.n18 VP.n17 8.76414
R37 VP.n31 VP.n30 8.76414
R38 VP.n14 VP.n13 8.76414
R39 VP.n10 VP.n9 0.189894
R40 VP.n11 VP.n10 0.189894
R41 VP.n11 VP.n4 0.189894
R42 VP.n15 VP.n4 0.189894
R43 VP.n19 VP.n16 0.189894
R44 VP.n20 VP.n19 0.189894
R45 VP.n21 VP.n20 0.189894
R46 VP.n21 VP.n2 0.189894
R47 VP.n26 VP.n2 0.189894
R48 VP.n27 VP.n26 0.189894
R49 VP.n28 VP.n27 0.189894
R50 VP.n28 VP.n0 0.189894
R51 VP.n32 VP.n0 0.189894
R52 VP VP.n32 0.0516364
R53 VDD1.n84 VDD1.n0 756.745
R54 VDD1.n173 VDD1.n89 756.745
R55 VDD1.n85 VDD1.n84 585
R56 VDD1.n83 VDD1.n82 585
R57 VDD1.n4 VDD1.n3 585
R58 VDD1.n77 VDD1.n76 585
R59 VDD1.n75 VDD1.n6 585
R60 VDD1.n74 VDD1.n73 585
R61 VDD1.n9 VDD1.n7 585
R62 VDD1.n68 VDD1.n67 585
R63 VDD1.n66 VDD1.n65 585
R64 VDD1.n13 VDD1.n12 585
R65 VDD1.n60 VDD1.n59 585
R66 VDD1.n58 VDD1.n57 585
R67 VDD1.n17 VDD1.n16 585
R68 VDD1.n52 VDD1.n51 585
R69 VDD1.n50 VDD1.n49 585
R70 VDD1.n21 VDD1.n20 585
R71 VDD1.n44 VDD1.n43 585
R72 VDD1.n42 VDD1.n41 585
R73 VDD1.n25 VDD1.n24 585
R74 VDD1.n36 VDD1.n35 585
R75 VDD1.n34 VDD1.n33 585
R76 VDD1.n29 VDD1.n28 585
R77 VDD1.n117 VDD1.n116 585
R78 VDD1.n122 VDD1.n121 585
R79 VDD1.n124 VDD1.n123 585
R80 VDD1.n113 VDD1.n112 585
R81 VDD1.n130 VDD1.n129 585
R82 VDD1.n132 VDD1.n131 585
R83 VDD1.n109 VDD1.n108 585
R84 VDD1.n138 VDD1.n137 585
R85 VDD1.n140 VDD1.n139 585
R86 VDD1.n105 VDD1.n104 585
R87 VDD1.n146 VDD1.n145 585
R88 VDD1.n148 VDD1.n147 585
R89 VDD1.n101 VDD1.n100 585
R90 VDD1.n154 VDD1.n153 585
R91 VDD1.n156 VDD1.n155 585
R92 VDD1.n97 VDD1.n96 585
R93 VDD1.n163 VDD1.n162 585
R94 VDD1.n164 VDD1.n95 585
R95 VDD1.n166 VDD1.n165 585
R96 VDD1.n93 VDD1.n92 585
R97 VDD1.n172 VDD1.n171 585
R98 VDD1.n174 VDD1.n173 585
R99 VDD1.n30 VDD1.t3 327.466
R100 VDD1.n118 VDD1.t0 327.466
R101 VDD1.n84 VDD1.n83 171.744
R102 VDD1.n83 VDD1.n3 171.744
R103 VDD1.n76 VDD1.n3 171.744
R104 VDD1.n76 VDD1.n75 171.744
R105 VDD1.n75 VDD1.n74 171.744
R106 VDD1.n74 VDD1.n7 171.744
R107 VDD1.n67 VDD1.n7 171.744
R108 VDD1.n67 VDD1.n66 171.744
R109 VDD1.n66 VDD1.n12 171.744
R110 VDD1.n59 VDD1.n12 171.744
R111 VDD1.n59 VDD1.n58 171.744
R112 VDD1.n58 VDD1.n16 171.744
R113 VDD1.n51 VDD1.n16 171.744
R114 VDD1.n51 VDD1.n50 171.744
R115 VDD1.n50 VDD1.n20 171.744
R116 VDD1.n43 VDD1.n20 171.744
R117 VDD1.n43 VDD1.n42 171.744
R118 VDD1.n42 VDD1.n24 171.744
R119 VDD1.n35 VDD1.n24 171.744
R120 VDD1.n35 VDD1.n34 171.744
R121 VDD1.n34 VDD1.n28 171.744
R122 VDD1.n122 VDD1.n116 171.744
R123 VDD1.n123 VDD1.n122 171.744
R124 VDD1.n123 VDD1.n112 171.744
R125 VDD1.n130 VDD1.n112 171.744
R126 VDD1.n131 VDD1.n130 171.744
R127 VDD1.n131 VDD1.n108 171.744
R128 VDD1.n138 VDD1.n108 171.744
R129 VDD1.n139 VDD1.n138 171.744
R130 VDD1.n139 VDD1.n104 171.744
R131 VDD1.n146 VDD1.n104 171.744
R132 VDD1.n147 VDD1.n146 171.744
R133 VDD1.n147 VDD1.n100 171.744
R134 VDD1.n154 VDD1.n100 171.744
R135 VDD1.n155 VDD1.n154 171.744
R136 VDD1.n155 VDD1.n96 171.744
R137 VDD1.n163 VDD1.n96 171.744
R138 VDD1.n164 VDD1.n163 171.744
R139 VDD1.n165 VDD1.n164 171.744
R140 VDD1.n165 VDD1.n92 171.744
R141 VDD1.n172 VDD1.n92 171.744
R142 VDD1.n173 VDD1.n172 171.744
R143 VDD1.t3 VDD1.n28 85.8723
R144 VDD1.t0 VDD1.n116 85.8723
R145 VDD1.n179 VDD1.n178 74.0413
R146 VDD1.n181 VDD1.n180 73.6807
R147 VDD1 VDD1.n88 54.049
R148 VDD1.n179 VDD1.n177 53.9354
R149 VDD1.n181 VDD1.n179 44.572
R150 VDD1.n30 VDD1.n29 16.3895
R151 VDD1.n118 VDD1.n117 16.3895
R152 VDD1.n77 VDD1.n6 13.1884
R153 VDD1.n166 VDD1.n95 13.1884
R154 VDD1.n78 VDD1.n4 12.8005
R155 VDD1.n73 VDD1.n8 12.8005
R156 VDD1.n33 VDD1.n32 12.8005
R157 VDD1.n121 VDD1.n120 12.8005
R158 VDD1.n162 VDD1.n161 12.8005
R159 VDD1.n167 VDD1.n93 12.8005
R160 VDD1.n82 VDD1.n81 12.0247
R161 VDD1.n72 VDD1.n9 12.0247
R162 VDD1.n36 VDD1.n27 12.0247
R163 VDD1.n124 VDD1.n115 12.0247
R164 VDD1.n160 VDD1.n97 12.0247
R165 VDD1.n171 VDD1.n170 12.0247
R166 VDD1.n85 VDD1.n2 11.249
R167 VDD1.n69 VDD1.n68 11.249
R168 VDD1.n37 VDD1.n25 11.249
R169 VDD1.n125 VDD1.n113 11.249
R170 VDD1.n157 VDD1.n156 11.249
R171 VDD1.n174 VDD1.n91 11.249
R172 VDD1.n86 VDD1.n0 10.4732
R173 VDD1.n65 VDD1.n11 10.4732
R174 VDD1.n41 VDD1.n40 10.4732
R175 VDD1.n129 VDD1.n128 10.4732
R176 VDD1.n153 VDD1.n99 10.4732
R177 VDD1.n175 VDD1.n89 10.4732
R178 VDD1.n64 VDD1.n13 9.69747
R179 VDD1.n44 VDD1.n23 9.69747
R180 VDD1.n132 VDD1.n111 9.69747
R181 VDD1.n152 VDD1.n101 9.69747
R182 VDD1.n88 VDD1.n87 9.45567
R183 VDD1.n177 VDD1.n176 9.45567
R184 VDD1.n56 VDD1.n55 9.3005
R185 VDD1.n15 VDD1.n14 9.3005
R186 VDD1.n62 VDD1.n61 9.3005
R187 VDD1.n64 VDD1.n63 9.3005
R188 VDD1.n11 VDD1.n10 9.3005
R189 VDD1.n70 VDD1.n69 9.3005
R190 VDD1.n72 VDD1.n71 9.3005
R191 VDD1.n8 VDD1.n5 9.3005
R192 VDD1.n87 VDD1.n86 9.3005
R193 VDD1.n2 VDD1.n1 9.3005
R194 VDD1.n81 VDD1.n80 9.3005
R195 VDD1.n79 VDD1.n78 9.3005
R196 VDD1.n54 VDD1.n53 9.3005
R197 VDD1.n19 VDD1.n18 9.3005
R198 VDD1.n48 VDD1.n47 9.3005
R199 VDD1.n46 VDD1.n45 9.3005
R200 VDD1.n23 VDD1.n22 9.3005
R201 VDD1.n40 VDD1.n39 9.3005
R202 VDD1.n38 VDD1.n37 9.3005
R203 VDD1.n27 VDD1.n26 9.3005
R204 VDD1.n32 VDD1.n31 9.3005
R205 VDD1.n176 VDD1.n175 9.3005
R206 VDD1.n91 VDD1.n90 9.3005
R207 VDD1.n170 VDD1.n169 9.3005
R208 VDD1.n168 VDD1.n167 9.3005
R209 VDD1.n107 VDD1.n106 9.3005
R210 VDD1.n136 VDD1.n135 9.3005
R211 VDD1.n134 VDD1.n133 9.3005
R212 VDD1.n111 VDD1.n110 9.3005
R213 VDD1.n128 VDD1.n127 9.3005
R214 VDD1.n126 VDD1.n125 9.3005
R215 VDD1.n115 VDD1.n114 9.3005
R216 VDD1.n120 VDD1.n119 9.3005
R217 VDD1.n142 VDD1.n141 9.3005
R218 VDD1.n144 VDD1.n143 9.3005
R219 VDD1.n103 VDD1.n102 9.3005
R220 VDD1.n150 VDD1.n149 9.3005
R221 VDD1.n152 VDD1.n151 9.3005
R222 VDD1.n99 VDD1.n98 9.3005
R223 VDD1.n158 VDD1.n157 9.3005
R224 VDD1.n160 VDD1.n159 9.3005
R225 VDD1.n161 VDD1.n94 9.3005
R226 VDD1.n61 VDD1.n60 8.92171
R227 VDD1.n45 VDD1.n21 8.92171
R228 VDD1.n133 VDD1.n109 8.92171
R229 VDD1.n149 VDD1.n148 8.92171
R230 VDD1.n57 VDD1.n15 8.14595
R231 VDD1.n49 VDD1.n48 8.14595
R232 VDD1.n137 VDD1.n136 8.14595
R233 VDD1.n145 VDD1.n103 8.14595
R234 VDD1.n56 VDD1.n17 7.3702
R235 VDD1.n52 VDD1.n19 7.3702
R236 VDD1.n140 VDD1.n107 7.3702
R237 VDD1.n144 VDD1.n105 7.3702
R238 VDD1.n53 VDD1.n17 6.59444
R239 VDD1.n53 VDD1.n52 6.59444
R240 VDD1.n141 VDD1.n140 6.59444
R241 VDD1.n141 VDD1.n105 6.59444
R242 VDD1.n57 VDD1.n56 5.81868
R243 VDD1.n49 VDD1.n19 5.81868
R244 VDD1.n137 VDD1.n107 5.81868
R245 VDD1.n145 VDD1.n144 5.81868
R246 VDD1.n60 VDD1.n15 5.04292
R247 VDD1.n48 VDD1.n21 5.04292
R248 VDD1.n136 VDD1.n109 5.04292
R249 VDD1.n148 VDD1.n103 5.04292
R250 VDD1.n61 VDD1.n13 4.26717
R251 VDD1.n45 VDD1.n44 4.26717
R252 VDD1.n133 VDD1.n132 4.26717
R253 VDD1.n149 VDD1.n101 4.26717
R254 VDD1.n31 VDD1.n30 3.70982
R255 VDD1.n119 VDD1.n118 3.70982
R256 VDD1.n88 VDD1.n0 3.49141
R257 VDD1.n65 VDD1.n64 3.49141
R258 VDD1.n41 VDD1.n23 3.49141
R259 VDD1.n129 VDD1.n111 3.49141
R260 VDD1.n153 VDD1.n152 3.49141
R261 VDD1.n177 VDD1.n89 3.49141
R262 VDD1.n86 VDD1.n85 2.71565
R263 VDD1.n68 VDD1.n11 2.71565
R264 VDD1.n40 VDD1.n25 2.71565
R265 VDD1.n128 VDD1.n113 2.71565
R266 VDD1.n156 VDD1.n99 2.71565
R267 VDD1.n175 VDD1.n174 2.71565
R268 VDD1.n180 VDD1.t4 1.99712
R269 VDD1.n180 VDD1.t2 1.99712
R270 VDD1.n178 VDD1.t1 1.99712
R271 VDD1.n178 VDD1.t5 1.99712
R272 VDD1.n82 VDD1.n2 1.93989
R273 VDD1.n69 VDD1.n9 1.93989
R274 VDD1.n37 VDD1.n36 1.93989
R275 VDD1.n125 VDD1.n124 1.93989
R276 VDD1.n157 VDD1.n97 1.93989
R277 VDD1.n171 VDD1.n91 1.93989
R278 VDD1.n81 VDD1.n4 1.16414
R279 VDD1.n73 VDD1.n72 1.16414
R280 VDD1.n33 VDD1.n27 1.16414
R281 VDD1.n121 VDD1.n115 1.16414
R282 VDD1.n162 VDD1.n160 1.16414
R283 VDD1.n170 VDD1.n93 1.16414
R284 VDD1.n78 VDD1.n77 0.388379
R285 VDD1.n8 VDD1.n6 0.388379
R286 VDD1.n32 VDD1.n29 0.388379
R287 VDD1.n120 VDD1.n117 0.388379
R288 VDD1.n161 VDD1.n95 0.388379
R289 VDD1.n167 VDD1.n166 0.388379
R290 VDD1 VDD1.n181 0.358259
R291 VDD1.n87 VDD1.n1 0.155672
R292 VDD1.n80 VDD1.n1 0.155672
R293 VDD1.n80 VDD1.n79 0.155672
R294 VDD1.n79 VDD1.n5 0.155672
R295 VDD1.n71 VDD1.n5 0.155672
R296 VDD1.n71 VDD1.n70 0.155672
R297 VDD1.n70 VDD1.n10 0.155672
R298 VDD1.n63 VDD1.n10 0.155672
R299 VDD1.n63 VDD1.n62 0.155672
R300 VDD1.n62 VDD1.n14 0.155672
R301 VDD1.n55 VDD1.n14 0.155672
R302 VDD1.n55 VDD1.n54 0.155672
R303 VDD1.n54 VDD1.n18 0.155672
R304 VDD1.n47 VDD1.n18 0.155672
R305 VDD1.n47 VDD1.n46 0.155672
R306 VDD1.n46 VDD1.n22 0.155672
R307 VDD1.n39 VDD1.n22 0.155672
R308 VDD1.n39 VDD1.n38 0.155672
R309 VDD1.n38 VDD1.n26 0.155672
R310 VDD1.n31 VDD1.n26 0.155672
R311 VDD1.n119 VDD1.n114 0.155672
R312 VDD1.n126 VDD1.n114 0.155672
R313 VDD1.n127 VDD1.n126 0.155672
R314 VDD1.n127 VDD1.n110 0.155672
R315 VDD1.n134 VDD1.n110 0.155672
R316 VDD1.n135 VDD1.n134 0.155672
R317 VDD1.n135 VDD1.n106 0.155672
R318 VDD1.n142 VDD1.n106 0.155672
R319 VDD1.n143 VDD1.n142 0.155672
R320 VDD1.n143 VDD1.n102 0.155672
R321 VDD1.n150 VDD1.n102 0.155672
R322 VDD1.n151 VDD1.n150 0.155672
R323 VDD1.n151 VDD1.n98 0.155672
R324 VDD1.n158 VDD1.n98 0.155672
R325 VDD1.n159 VDD1.n158 0.155672
R326 VDD1.n159 VDD1.n94 0.155672
R327 VDD1.n168 VDD1.n94 0.155672
R328 VDD1.n169 VDD1.n168 0.155672
R329 VDD1.n169 VDD1.n90 0.155672
R330 VDD1.n176 VDD1.n90 0.155672
R331 VTAIL.n362 VTAIL.n278 756.745
R332 VTAIL.n86 VTAIL.n2 756.745
R333 VTAIL.n272 VTAIL.n188 756.745
R334 VTAIL.n180 VTAIL.n96 756.745
R335 VTAIL.n306 VTAIL.n305 585
R336 VTAIL.n311 VTAIL.n310 585
R337 VTAIL.n313 VTAIL.n312 585
R338 VTAIL.n302 VTAIL.n301 585
R339 VTAIL.n319 VTAIL.n318 585
R340 VTAIL.n321 VTAIL.n320 585
R341 VTAIL.n298 VTAIL.n297 585
R342 VTAIL.n327 VTAIL.n326 585
R343 VTAIL.n329 VTAIL.n328 585
R344 VTAIL.n294 VTAIL.n293 585
R345 VTAIL.n335 VTAIL.n334 585
R346 VTAIL.n337 VTAIL.n336 585
R347 VTAIL.n290 VTAIL.n289 585
R348 VTAIL.n343 VTAIL.n342 585
R349 VTAIL.n345 VTAIL.n344 585
R350 VTAIL.n286 VTAIL.n285 585
R351 VTAIL.n352 VTAIL.n351 585
R352 VTAIL.n353 VTAIL.n284 585
R353 VTAIL.n355 VTAIL.n354 585
R354 VTAIL.n282 VTAIL.n281 585
R355 VTAIL.n361 VTAIL.n360 585
R356 VTAIL.n363 VTAIL.n362 585
R357 VTAIL.n30 VTAIL.n29 585
R358 VTAIL.n35 VTAIL.n34 585
R359 VTAIL.n37 VTAIL.n36 585
R360 VTAIL.n26 VTAIL.n25 585
R361 VTAIL.n43 VTAIL.n42 585
R362 VTAIL.n45 VTAIL.n44 585
R363 VTAIL.n22 VTAIL.n21 585
R364 VTAIL.n51 VTAIL.n50 585
R365 VTAIL.n53 VTAIL.n52 585
R366 VTAIL.n18 VTAIL.n17 585
R367 VTAIL.n59 VTAIL.n58 585
R368 VTAIL.n61 VTAIL.n60 585
R369 VTAIL.n14 VTAIL.n13 585
R370 VTAIL.n67 VTAIL.n66 585
R371 VTAIL.n69 VTAIL.n68 585
R372 VTAIL.n10 VTAIL.n9 585
R373 VTAIL.n76 VTAIL.n75 585
R374 VTAIL.n77 VTAIL.n8 585
R375 VTAIL.n79 VTAIL.n78 585
R376 VTAIL.n6 VTAIL.n5 585
R377 VTAIL.n85 VTAIL.n84 585
R378 VTAIL.n87 VTAIL.n86 585
R379 VTAIL.n273 VTAIL.n272 585
R380 VTAIL.n271 VTAIL.n270 585
R381 VTAIL.n192 VTAIL.n191 585
R382 VTAIL.n265 VTAIL.n264 585
R383 VTAIL.n263 VTAIL.n194 585
R384 VTAIL.n262 VTAIL.n261 585
R385 VTAIL.n197 VTAIL.n195 585
R386 VTAIL.n256 VTAIL.n255 585
R387 VTAIL.n254 VTAIL.n253 585
R388 VTAIL.n201 VTAIL.n200 585
R389 VTAIL.n248 VTAIL.n247 585
R390 VTAIL.n246 VTAIL.n245 585
R391 VTAIL.n205 VTAIL.n204 585
R392 VTAIL.n240 VTAIL.n239 585
R393 VTAIL.n238 VTAIL.n237 585
R394 VTAIL.n209 VTAIL.n208 585
R395 VTAIL.n232 VTAIL.n231 585
R396 VTAIL.n230 VTAIL.n229 585
R397 VTAIL.n213 VTAIL.n212 585
R398 VTAIL.n224 VTAIL.n223 585
R399 VTAIL.n222 VTAIL.n221 585
R400 VTAIL.n217 VTAIL.n216 585
R401 VTAIL.n181 VTAIL.n180 585
R402 VTAIL.n179 VTAIL.n178 585
R403 VTAIL.n100 VTAIL.n99 585
R404 VTAIL.n173 VTAIL.n172 585
R405 VTAIL.n171 VTAIL.n102 585
R406 VTAIL.n170 VTAIL.n169 585
R407 VTAIL.n105 VTAIL.n103 585
R408 VTAIL.n164 VTAIL.n163 585
R409 VTAIL.n162 VTAIL.n161 585
R410 VTAIL.n109 VTAIL.n108 585
R411 VTAIL.n156 VTAIL.n155 585
R412 VTAIL.n154 VTAIL.n153 585
R413 VTAIL.n113 VTAIL.n112 585
R414 VTAIL.n148 VTAIL.n147 585
R415 VTAIL.n146 VTAIL.n145 585
R416 VTAIL.n117 VTAIL.n116 585
R417 VTAIL.n140 VTAIL.n139 585
R418 VTAIL.n138 VTAIL.n137 585
R419 VTAIL.n121 VTAIL.n120 585
R420 VTAIL.n132 VTAIL.n131 585
R421 VTAIL.n130 VTAIL.n129 585
R422 VTAIL.n125 VTAIL.n124 585
R423 VTAIL.n307 VTAIL.t2 327.466
R424 VTAIL.n31 VTAIL.t7 327.466
R425 VTAIL.n218 VTAIL.t8 327.466
R426 VTAIL.n126 VTAIL.t5 327.466
R427 VTAIL.n311 VTAIL.n305 171.744
R428 VTAIL.n312 VTAIL.n311 171.744
R429 VTAIL.n312 VTAIL.n301 171.744
R430 VTAIL.n319 VTAIL.n301 171.744
R431 VTAIL.n320 VTAIL.n319 171.744
R432 VTAIL.n320 VTAIL.n297 171.744
R433 VTAIL.n327 VTAIL.n297 171.744
R434 VTAIL.n328 VTAIL.n327 171.744
R435 VTAIL.n328 VTAIL.n293 171.744
R436 VTAIL.n335 VTAIL.n293 171.744
R437 VTAIL.n336 VTAIL.n335 171.744
R438 VTAIL.n336 VTAIL.n289 171.744
R439 VTAIL.n343 VTAIL.n289 171.744
R440 VTAIL.n344 VTAIL.n343 171.744
R441 VTAIL.n344 VTAIL.n285 171.744
R442 VTAIL.n352 VTAIL.n285 171.744
R443 VTAIL.n353 VTAIL.n352 171.744
R444 VTAIL.n354 VTAIL.n353 171.744
R445 VTAIL.n354 VTAIL.n281 171.744
R446 VTAIL.n361 VTAIL.n281 171.744
R447 VTAIL.n362 VTAIL.n361 171.744
R448 VTAIL.n35 VTAIL.n29 171.744
R449 VTAIL.n36 VTAIL.n35 171.744
R450 VTAIL.n36 VTAIL.n25 171.744
R451 VTAIL.n43 VTAIL.n25 171.744
R452 VTAIL.n44 VTAIL.n43 171.744
R453 VTAIL.n44 VTAIL.n21 171.744
R454 VTAIL.n51 VTAIL.n21 171.744
R455 VTAIL.n52 VTAIL.n51 171.744
R456 VTAIL.n52 VTAIL.n17 171.744
R457 VTAIL.n59 VTAIL.n17 171.744
R458 VTAIL.n60 VTAIL.n59 171.744
R459 VTAIL.n60 VTAIL.n13 171.744
R460 VTAIL.n67 VTAIL.n13 171.744
R461 VTAIL.n68 VTAIL.n67 171.744
R462 VTAIL.n68 VTAIL.n9 171.744
R463 VTAIL.n76 VTAIL.n9 171.744
R464 VTAIL.n77 VTAIL.n76 171.744
R465 VTAIL.n78 VTAIL.n77 171.744
R466 VTAIL.n78 VTAIL.n5 171.744
R467 VTAIL.n85 VTAIL.n5 171.744
R468 VTAIL.n86 VTAIL.n85 171.744
R469 VTAIL.n272 VTAIL.n271 171.744
R470 VTAIL.n271 VTAIL.n191 171.744
R471 VTAIL.n264 VTAIL.n191 171.744
R472 VTAIL.n264 VTAIL.n263 171.744
R473 VTAIL.n263 VTAIL.n262 171.744
R474 VTAIL.n262 VTAIL.n195 171.744
R475 VTAIL.n255 VTAIL.n195 171.744
R476 VTAIL.n255 VTAIL.n254 171.744
R477 VTAIL.n254 VTAIL.n200 171.744
R478 VTAIL.n247 VTAIL.n200 171.744
R479 VTAIL.n247 VTAIL.n246 171.744
R480 VTAIL.n246 VTAIL.n204 171.744
R481 VTAIL.n239 VTAIL.n204 171.744
R482 VTAIL.n239 VTAIL.n238 171.744
R483 VTAIL.n238 VTAIL.n208 171.744
R484 VTAIL.n231 VTAIL.n208 171.744
R485 VTAIL.n231 VTAIL.n230 171.744
R486 VTAIL.n230 VTAIL.n212 171.744
R487 VTAIL.n223 VTAIL.n212 171.744
R488 VTAIL.n223 VTAIL.n222 171.744
R489 VTAIL.n222 VTAIL.n216 171.744
R490 VTAIL.n180 VTAIL.n179 171.744
R491 VTAIL.n179 VTAIL.n99 171.744
R492 VTAIL.n172 VTAIL.n99 171.744
R493 VTAIL.n172 VTAIL.n171 171.744
R494 VTAIL.n171 VTAIL.n170 171.744
R495 VTAIL.n170 VTAIL.n103 171.744
R496 VTAIL.n163 VTAIL.n103 171.744
R497 VTAIL.n163 VTAIL.n162 171.744
R498 VTAIL.n162 VTAIL.n108 171.744
R499 VTAIL.n155 VTAIL.n108 171.744
R500 VTAIL.n155 VTAIL.n154 171.744
R501 VTAIL.n154 VTAIL.n112 171.744
R502 VTAIL.n147 VTAIL.n112 171.744
R503 VTAIL.n147 VTAIL.n146 171.744
R504 VTAIL.n146 VTAIL.n116 171.744
R505 VTAIL.n139 VTAIL.n116 171.744
R506 VTAIL.n139 VTAIL.n138 171.744
R507 VTAIL.n138 VTAIL.n120 171.744
R508 VTAIL.n131 VTAIL.n120 171.744
R509 VTAIL.n131 VTAIL.n130 171.744
R510 VTAIL.n130 VTAIL.n124 171.744
R511 VTAIL.t2 VTAIL.n305 85.8723
R512 VTAIL.t7 VTAIL.n29 85.8723
R513 VTAIL.t8 VTAIL.n216 85.8723
R514 VTAIL.t5 VTAIL.n124 85.8723
R515 VTAIL.n187 VTAIL.n186 57.0021
R516 VTAIL.n95 VTAIL.n94 57.0021
R517 VTAIL.n1 VTAIL.n0 57.0019
R518 VTAIL.n93 VTAIL.n92 57.0019
R519 VTAIL.n367 VTAIL.n366 36.0641
R520 VTAIL.n91 VTAIL.n90 36.0641
R521 VTAIL.n277 VTAIL.n276 36.0641
R522 VTAIL.n185 VTAIL.n184 36.0641
R523 VTAIL.n95 VTAIL.n93 29.7289
R524 VTAIL.n367 VTAIL.n277 28.0652
R525 VTAIL.n307 VTAIL.n306 16.3895
R526 VTAIL.n31 VTAIL.n30 16.3895
R527 VTAIL.n218 VTAIL.n217 16.3895
R528 VTAIL.n126 VTAIL.n125 16.3895
R529 VTAIL.n355 VTAIL.n284 13.1884
R530 VTAIL.n79 VTAIL.n8 13.1884
R531 VTAIL.n265 VTAIL.n194 13.1884
R532 VTAIL.n173 VTAIL.n102 13.1884
R533 VTAIL.n310 VTAIL.n309 12.8005
R534 VTAIL.n351 VTAIL.n350 12.8005
R535 VTAIL.n356 VTAIL.n282 12.8005
R536 VTAIL.n34 VTAIL.n33 12.8005
R537 VTAIL.n75 VTAIL.n74 12.8005
R538 VTAIL.n80 VTAIL.n6 12.8005
R539 VTAIL.n266 VTAIL.n192 12.8005
R540 VTAIL.n261 VTAIL.n196 12.8005
R541 VTAIL.n221 VTAIL.n220 12.8005
R542 VTAIL.n174 VTAIL.n100 12.8005
R543 VTAIL.n169 VTAIL.n104 12.8005
R544 VTAIL.n129 VTAIL.n128 12.8005
R545 VTAIL.n313 VTAIL.n304 12.0247
R546 VTAIL.n349 VTAIL.n286 12.0247
R547 VTAIL.n360 VTAIL.n359 12.0247
R548 VTAIL.n37 VTAIL.n28 12.0247
R549 VTAIL.n73 VTAIL.n10 12.0247
R550 VTAIL.n84 VTAIL.n83 12.0247
R551 VTAIL.n270 VTAIL.n269 12.0247
R552 VTAIL.n260 VTAIL.n197 12.0247
R553 VTAIL.n224 VTAIL.n215 12.0247
R554 VTAIL.n178 VTAIL.n177 12.0247
R555 VTAIL.n168 VTAIL.n105 12.0247
R556 VTAIL.n132 VTAIL.n123 12.0247
R557 VTAIL.n314 VTAIL.n302 11.249
R558 VTAIL.n346 VTAIL.n345 11.249
R559 VTAIL.n363 VTAIL.n280 11.249
R560 VTAIL.n38 VTAIL.n26 11.249
R561 VTAIL.n70 VTAIL.n69 11.249
R562 VTAIL.n87 VTAIL.n4 11.249
R563 VTAIL.n273 VTAIL.n190 11.249
R564 VTAIL.n257 VTAIL.n256 11.249
R565 VTAIL.n225 VTAIL.n213 11.249
R566 VTAIL.n181 VTAIL.n98 11.249
R567 VTAIL.n165 VTAIL.n164 11.249
R568 VTAIL.n133 VTAIL.n121 11.249
R569 VTAIL.n318 VTAIL.n317 10.4732
R570 VTAIL.n342 VTAIL.n288 10.4732
R571 VTAIL.n364 VTAIL.n278 10.4732
R572 VTAIL.n42 VTAIL.n41 10.4732
R573 VTAIL.n66 VTAIL.n12 10.4732
R574 VTAIL.n88 VTAIL.n2 10.4732
R575 VTAIL.n274 VTAIL.n188 10.4732
R576 VTAIL.n253 VTAIL.n199 10.4732
R577 VTAIL.n229 VTAIL.n228 10.4732
R578 VTAIL.n182 VTAIL.n96 10.4732
R579 VTAIL.n161 VTAIL.n107 10.4732
R580 VTAIL.n137 VTAIL.n136 10.4732
R581 VTAIL.n321 VTAIL.n300 9.69747
R582 VTAIL.n341 VTAIL.n290 9.69747
R583 VTAIL.n45 VTAIL.n24 9.69747
R584 VTAIL.n65 VTAIL.n14 9.69747
R585 VTAIL.n252 VTAIL.n201 9.69747
R586 VTAIL.n232 VTAIL.n211 9.69747
R587 VTAIL.n160 VTAIL.n109 9.69747
R588 VTAIL.n140 VTAIL.n119 9.69747
R589 VTAIL.n366 VTAIL.n365 9.45567
R590 VTAIL.n90 VTAIL.n89 9.45567
R591 VTAIL.n276 VTAIL.n275 9.45567
R592 VTAIL.n184 VTAIL.n183 9.45567
R593 VTAIL.n365 VTAIL.n364 9.3005
R594 VTAIL.n280 VTAIL.n279 9.3005
R595 VTAIL.n359 VTAIL.n358 9.3005
R596 VTAIL.n357 VTAIL.n356 9.3005
R597 VTAIL.n296 VTAIL.n295 9.3005
R598 VTAIL.n325 VTAIL.n324 9.3005
R599 VTAIL.n323 VTAIL.n322 9.3005
R600 VTAIL.n300 VTAIL.n299 9.3005
R601 VTAIL.n317 VTAIL.n316 9.3005
R602 VTAIL.n315 VTAIL.n314 9.3005
R603 VTAIL.n304 VTAIL.n303 9.3005
R604 VTAIL.n309 VTAIL.n308 9.3005
R605 VTAIL.n331 VTAIL.n330 9.3005
R606 VTAIL.n333 VTAIL.n332 9.3005
R607 VTAIL.n292 VTAIL.n291 9.3005
R608 VTAIL.n339 VTAIL.n338 9.3005
R609 VTAIL.n341 VTAIL.n340 9.3005
R610 VTAIL.n288 VTAIL.n287 9.3005
R611 VTAIL.n347 VTAIL.n346 9.3005
R612 VTAIL.n349 VTAIL.n348 9.3005
R613 VTAIL.n350 VTAIL.n283 9.3005
R614 VTAIL.n89 VTAIL.n88 9.3005
R615 VTAIL.n4 VTAIL.n3 9.3005
R616 VTAIL.n83 VTAIL.n82 9.3005
R617 VTAIL.n81 VTAIL.n80 9.3005
R618 VTAIL.n20 VTAIL.n19 9.3005
R619 VTAIL.n49 VTAIL.n48 9.3005
R620 VTAIL.n47 VTAIL.n46 9.3005
R621 VTAIL.n24 VTAIL.n23 9.3005
R622 VTAIL.n41 VTAIL.n40 9.3005
R623 VTAIL.n39 VTAIL.n38 9.3005
R624 VTAIL.n28 VTAIL.n27 9.3005
R625 VTAIL.n33 VTAIL.n32 9.3005
R626 VTAIL.n55 VTAIL.n54 9.3005
R627 VTAIL.n57 VTAIL.n56 9.3005
R628 VTAIL.n16 VTAIL.n15 9.3005
R629 VTAIL.n63 VTAIL.n62 9.3005
R630 VTAIL.n65 VTAIL.n64 9.3005
R631 VTAIL.n12 VTAIL.n11 9.3005
R632 VTAIL.n71 VTAIL.n70 9.3005
R633 VTAIL.n73 VTAIL.n72 9.3005
R634 VTAIL.n74 VTAIL.n7 9.3005
R635 VTAIL.n244 VTAIL.n243 9.3005
R636 VTAIL.n203 VTAIL.n202 9.3005
R637 VTAIL.n250 VTAIL.n249 9.3005
R638 VTAIL.n252 VTAIL.n251 9.3005
R639 VTAIL.n199 VTAIL.n198 9.3005
R640 VTAIL.n258 VTAIL.n257 9.3005
R641 VTAIL.n260 VTAIL.n259 9.3005
R642 VTAIL.n196 VTAIL.n193 9.3005
R643 VTAIL.n275 VTAIL.n274 9.3005
R644 VTAIL.n190 VTAIL.n189 9.3005
R645 VTAIL.n269 VTAIL.n268 9.3005
R646 VTAIL.n267 VTAIL.n266 9.3005
R647 VTAIL.n242 VTAIL.n241 9.3005
R648 VTAIL.n207 VTAIL.n206 9.3005
R649 VTAIL.n236 VTAIL.n235 9.3005
R650 VTAIL.n234 VTAIL.n233 9.3005
R651 VTAIL.n211 VTAIL.n210 9.3005
R652 VTAIL.n228 VTAIL.n227 9.3005
R653 VTAIL.n226 VTAIL.n225 9.3005
R654 VTAIL.n215 VTAIL.n214 9.3005
R655 VTAIL.n220 VTAIL.n219 9.3005
R656 VTAIL.n152 VTAIL.n151 9.3005
R657 VTAIL.n111 VTAIL.n110 9.3005
R658 VTAIL.n158 VTAIL.n157 9.3005
R659 VTAIL.n160 VTAIL.n159 9.3005
R660 VTAIL.n107 VTAIL.n106 9.3005
R661 VTAIL.n166 VTAIL.n165 9.3005
R662 VTAIL.n168 VTAIL.n167 9.3005
R663 VTAIL.n104 VTAIL.n101 9.3005
R664 VTAIL.n183 VTAIL.n182 9.3005
R665 VTAIL.n98 VTAIL.n97 9.3005
R666 VTAIL.n177 VTAIL.n176 9.3005
R667 VTAIL.n175 VTAIL.n174 9.3005
R668 VTAIL.n150 VTAIL.n149 9.3005
R669 VTAIL.n115 VTAIL.n114 9.3005
R670 VTAIL.n144 VTAIL.n143 9.3005
R671 VTAIL.n142 VTAIL.n141 9.3005
R672 VTAIL.n119 VTAIL.n118 9.3005
R673 VTAIL.n136 VTAIL.n135 9.3005
R674 VTAIL.n134 VTAIL.n133 9.3005
R675 VTAIL.n123 VTAIL.n122 9.3005
R676 VTAIL.n128 VTAIL.n127 9.3005
R677 VTAIL.n322 VTAIL.n298 8.92171
R678 VTAIL.n338 VTAIL.n337 8.92171
R679 VTAIL.n46 VTAIL.n22 8.92171
R680 VTAIL.n62 VTAIL.n61 8.92171
R681 VTAIL.n249 VTAIL.n248 8.92171
R682 VTAIL.n233 VTAIL.n209 8.92171
R683 VTAIL.n157 VTAIL.n156 8.92171
R684 VTAIL.n141 VTAIL.n117 8.92171
R685 VTAIL.n326 VTAIL.n325 8.14595
R686 VTAIL.n334 VTAIL.n292 8.14595
R687 VTAIL.n50 VTAIL.n49 8.14595
R688 VTAIL.n58 VTAIL.n16 8.14595
R689 VTAIL.n245 VTAIL.n203 8.14595
R690 VTAIL.n237 VTAIL.n236 8.14595
R691 VTAIL.n153 VTAIL.n111 8.14595
R692 VTAIL.n145 VTAIL.n144 8.14595
R693 VTAIL.n329 VTAIL.n296 7.3702
R694 VTAIL.n333 VTAIL.n294 7.3702
R695 VTAIL.n53 VTAIL.n20 7.3702
R696 VTAIL.n57 VTAIL.n18 7.3702
R697 VTAIL.n244 VTAIL.n205 7.3702
R698 VTAIL.n240 VTAIL.n207 7.3702
R699 VTAIL.n152 VTAIL.n113 7.3702
R700 VTAIL.n148 VTAIL.n115 7.3702
R701 VTAIL.n330 VTAIL.n329 6.59444
R702 VTAIL.n330 VTAIL.n294 6.59444
R703 VTAIL.n54 VTAIL.n53 6.59444
R704 VTAIL.n54 VTAIL.n18 6.59444
R705 VTAIL.n241 VTAIL.n205 6.59444
R706 VTAIL.n241 VTAIL.n240 6.59444
R707 VTAIL.n149 VTAIL.n113 6.59444
R708 VTAIL.n149 VTAIL.n148 6.59444
R709 VTAIL.n326 VTAIL.n296 5.81868
R710 VTAIL.n334 VTAIL.n333 5.81868
R711 VTAIL.n50 VTAIL.n20 5.81868
R712 VTAIL.n58 VTAIL.n57 5.81868
R713 VTAIL.n245 VTAIL.n244 5.81868
R714 VTAIL.n237 VTAIL.n207 5.81868
R715 VTAIL.n153 VTAIL.n152 5.81868
R716 VTAIL.n145 VTAIL.n115 5.81868
R717 VTAIL.n325 VTAIL.n298 5.04292
R718 VTAIL.n337 VTAIL.n292 5.04292
R719 VTAIL.n49 VTAIL.n22 5.04292
R720 VTAIL.n61 VTAIL.n16 5.04292
R721 VTAIL.n248 VTAIL.n203 5.04292
R722 VTAIL.n236 VTAIL.n209 5.04292
R723 VTAIL.n156 VTAIL.n111 5.04292
R724 VTAIL.n144 VTAIL.n117 5.04292
R725 VTAIL.n322 VTAIL.n321 4.26717
R726 VTAIL.n338 VTAIL.n290 4.26717
R727 VTAIL.n46 VTAIL.n45 4.26717
R728 VTAIL.n62 VTAIL.n14 4.26717
R729 VTAIL.n249 VTAIL.n201 4.26717
R730 VTAIL.n233 VTAIL.n232 4.26717
R731 VTAIL.n157 VTAIL.n109 4.26717
R732 VTAIL.n141 VTAIL.n140 4.26717
R733 VTAIL.n308 VTAIL.n307 3.70982
R734 VTAIL.n32 VTAIL.n31 3.70982
R735 VTAIL.n219 VTAIL.n218 3.70982
R736 VTAIL.n127 VTAIL.n126 3.70982
R737 VTAIL.n318 VTAIL.n300 3.49141
R738 VTAIL.n342 VTAIL.n341 3.49141
R739 VTAIL.n366 VTAIL.n278 3.49141
R740 VTAIL.n42 VTAIL.n24 3.49141
R741 VTAIL.n66 VTAIL.n65 3.49141
R742 VTAIL.n90 VTAIL.n2 3.49141
R743 VTAIL.n276 VTAIL.n188 3.49141
R744 VTAIL.n253 VTAIL.n252 3.49141
R745 VTAIL.n229 VTAIL.n211 3.49141
R746 VTAIL.n184 VTAIL.n96 3.49141
R747 VTAIL.n161 VTAIL.n160 3.49141
R748 VTAIL.n137 VTAIL.n119 3.49141
R749 VTAIL.n317 VTAIL.n302 2.71565
R750 VTAIL.n345 VTAIL.n288 2.71565
R751 VTAIL.n364 VTAIL.n363 2.71565
R752 VTAIL.n41 VTAIL.n26 2.71565
R753 VTAIL.n69 VTAIL.n12 2.71565
R754 VTAIL.n88 VTAIL.n87 2.71565
R755 VTAIL.n274 VTAIL.n273 2.71565
R756 VTAIL.n256 VTAIL.n199 2.71565
R757 VTAIL.n228 VTAIL.n213 2.71565
R758 VTAIL.n182 VTAIL.n181 2.71565
R759 VTAIL.n164 VTAIL.n107 2.71565
R760 VTAIL.n136 VTAIL.n121 2.71565
R761 VTAIL.n0 VTAIL.t1 1.99712
R762 VTAIL.n0 VTAIL.t0 1.99712
R763 VTAIL.n92 VTAIL.t10 1.99712
R764 VTAIL.n92 VTAIL.t11 1.99712
R765 VTAIL.n186 VTAIL.t6 1.99712
R766 VTAIL.n186 VTAIL.t9 1.99712
R767 VTAIL.n94 VTAIL.t3 1.99712
R768 VTAIL.n94 VTAIL.t4 1.99712
R769 VTAIL.n314 VTAIL.n313 1.93989
R770 VTAIL.n346 VTAIL.n286 1.93989
R771 VTAIL.n360 VTAIL.n280 1.93989
R772 VTAIL.n38 VTAIL.n37 1.93989
R773 VTAIL.n70 VTAIL.n10 1.93989
R774 VTAIL.n84 VTAIL.n4 1.93989
R775 VTAIL.n270 VTAIL.n190 1.93989
R776 VTAIL.n257 VTAIL.n197 1.93989
R777 VTAIL.n225 VTAIL.n224 1.93989
R778 VTAIL.n178 VTAIL.n98 1.93989
R779 VTAIL.n165 VTAIL.n105 1.93989
R780 VTAIL.n133 VTAIL.n132 1.93989
R781 VTAIL.n185 VTAIL.n95 1.66429
R782 VTAIL.n277 VTAIL.n187 1.66429
R783 VTAIL.n93 VTAIL.n91 1.66429
R784 VTAIL.n187 VTAIL.n185 1.30222
R785 VTAIL.n91 VTAIL.n1 1.30222
R786 VTAIL VTAIL.n367 1.19016
R787 VTAIL.n310 VTAIL.n304 1.16414
R788 VTAIL.n351 VTAIL.n349 1.16414
R789 VTAIL.n359 VTAIL.n282 1.16414
R790 VTAIL.n34 VTAIL.n28 1.16414
R791 VTAIL.n75 VTAIL.n73 1.16414
R792 VTAIL.n83 VTAIL.n6 1.16414
R793 VTAIL.n269 VTAIL.n192 1.16414
R794 VTAIL.n261 VTAIL.n260 1.16414
R795 VTAIL.n221 VTAIL.n215 1.16414
R796 VTAIL.n177 VTAIL.n100 1.16414
R797 VTAIL.n169 VTAIL.n168 1.16414
R798 VTAIL.n129 VTAIL.n123 1.16414
R799 VTAIL VTAIL.n1 0.474638
R800 VTAIL.n309 VTAIL.n306 0.388379
R801 VTAIL.n350 VTAIL.n284 0.388379
R802 VTAIL.n356 VTAIL.n355 0.388379
R803 VTAIL.n33 VTAIL.n30 0.388379
R804 VTAIL.n74 VTAIL.n8 0.388379
R805 VTAIL.n80 VTAIL.n79 0.388379
R806 VTAIL.n266 VTAIL.n265 0.388379
R807 VTAIL.n196 VTAIL.n194 0.388379
R808 VTAIL.n220 VTAIL.n217 0.388379
R809 VTAIL.n174 VTAIL.n173 0.388379
R810 VTAIL.n104 VTAIL.n102 0.388379
R811 VTAIL.n128 VTAIL.n125 0.388379
R812 VTAIL.n308 VTAIL.n303 0.155672
R813 VTAIL.n315 VTAIL.n303 0.155672
R814 VTAIL.n316 VTAIL.n315 0.155672
R815 VTAIL.n316 VTAIL.n299 0.155672
R816 VTAIL.n323 VTAIL.n299 0.155672
R817 VTAIL.n324 VTAIL.n323 0.155672
R818 VTAIL.n324 VTAIL.n295 0.155672
R819 VTAIL.n331 VTAIL.n295 0.155672
R820 VTAIL.n332 VTAIL.n331 0.155672
R821 VTAIL.n332 VTAIL.n291 0.155672
R822 VTAIL.n339 VTAIL.n291 0.155672
R823 VTAIL.n340 VTAIL.n339 0.155672
R824 VTAIL.n340 VTAIL.n287 0.155672
R825 VTAIL.n347 VTAIL.n287 0.155672
R826 VTAIL.n348 VTAIL.n347 0.155672
R827 VTAIL.n348 VTAIL.n283 0.155672
R828 VTAIL.n357 VTAIL.n283 0.155672
R829 VTAIL.n358 VTAIL.n357 0.155672
R830 VTAIL.n358 VTAIL.n279 0.155672
R831 VTAIL.n365 VTAIL.n279 0.155672
R832 VTAIL.n32 VTAIL.n27 0.155672
R833 VTAIL.n39 VTAIL.n27 0.155672
R834 VTAIL.n40 VTAIL.n39 0.155672
R835 VTAIL.n40 VTAIL.n23 0.155672
R836 VTAIL.n47 VTAIL.n23 0.155672
R837 VTAIL.n48 VTAIL.n47 0.155672
R838 VTAIL.n48 VTAIL.n19 0.155672
R839 VTAIL.n55 VTAIL.n19 0.155672
R840 VTAIL.n56 VTAIL.n55 0.155672
R841 VTAIL.n56 VTAIL.n15 0.155672
R842 VTAIL.n63 VTAIL.n15 0.155672
R843 VTAIL.n64 VTAIL.n63 0.155672
R844 VTAIL.n64 VTAIL.n11 0.155672
R845 VTAIL.n71 VTAIL.n11 0.155672
R846 VTAIL.n72 VTAIL.n71 0.155672
R847 VTAIL.n72 VTAIL.n7 0.155672
R848 VTAIL.n81 VTAIL.n7 0.155672
R849 VTAIL.n82 VTAIL.n81 0.155672
R850 VTAIL.n82 VTAIL.n3 0.155672
R851 VTAIL.n89 VTAIL.n3 0.155672
R852 VTAIL.n275 VTAIL.n189 0.155672
R853 VTAIL.n268 VTAIL.n189 0.155672
R854 VTAIL.n268 VTAIL.n267 0.155672
R855 VTAIL.n267 VTAIL.n193 0.155672
R856 VTAIL.n259 VTAIL.n193 0.155672
R857 VTAIL.n259 VTAIL.n258 0.155672
R858 VTAIL.n258 VTAIL.n198 0.155672
R859 VTAIL.n251 VTAIL.n198 0.155672
R860 VTAIL.n251 VTAIL.n250 0.155672
R861 VTAIL.n250 VTAIL.n202 0.155672
R862 VTAIL.n243 VTAIL.n202 0.155672
R863 VTAIL.n243 VTAIL.n242 0.155672
R864 VTAIL.n242 VTAIL.n206 0.155672
R865 VTAIL.n235 VTAIL.n206 0.155672
R866 VTAIL.n235 VTAIL.n234 0.155672
R867 VTAIL.n234 VTAIL.n210 0.155672
R868 VTAIL.n227 VTAIL.n210 0.155672
R869 VTAIL.n227 VTAIL.n226 0.155672
R870 VTAIL.n226 VTAIL.n214 0.155672
R871 VTAIL.n219 VTAIL.n214 0.155672
R872 VTAIL.n183 VTAIL.n97 0.155672
R873 VTAIL.n176 VTAIL.n97 0.155672
R874 VTAIL.n176 VTAIL.n175 0.155672
R875 VTAIL.n175 VTAIL.n101 0.155672
R876 VTAIL.n167 VTAIL.n101 0.155672
R877 VTAIL.n167 VTAIL.n166 0.155672
R878 VTAIL.n166 VTAIL.n106 0.155672
R879 VTAIL.n159 VTAIL.n106 0.155672
R880 VTAIL.n159 VTAIL.n158 0.155672
R881 VTAIL.n158 VTAIL.n110 0.155672
R882 VTAIL.n151 VTAIL.n110 0.155672
R883 VTAIL.n151 VTAIL.n150 0.155672
R884 VTAIL.n150 VTAIL.n114 0.155672
R885 VTAIL.n143 VTAIL.n114 0.155672
R886 VTAIL.n143 VTAIL.n142 0.155672
R887 VTAIL.n142 VTAIL.n118 0.155672
R888 VTAIL.n135 VTAIL.n118 0.155672
R889 VTAIL.n135 VTAIL.n134 0.155672
R890 VTAIL.n134 VTAIL.n122 0.155672
R891 VTAIL.n127 VTAIL.n122 0.155672
R892 VN.n2 VN.t1 278.24
R893 VN.n14 VN.t2 278.24
R894 VN.n3 VN.t3 245.218
R895 VN.n10 VN.t4 245.218
R896 VN.n15 VN.t5 245.218
R897 VN.n22 VN.t0 245.218
R898 VN.n11 VN.n10 176.881
R899 VN.n23 VN.n22 176.881
R900 VN.n21 VN.n12 161.3
R901 VN.n20 VN.n19 161.3
R902 VN.n18 VN.n13 161.3
R903 VN.n17 VN.n16 161.3
R904 VN.n9 VN.n0 161.3
R905 VN.n8 VN.n7 161.3
R906 VN.n6 VN.n1 161.3
R907 VN.n5 VN.n4 161.3
R908 VN.n8 VN.n1 56.4773
R909 VN.n20 VN.n13 56.4773
R910 VN.n3 VN.n2 53.8729
R911 VN.n15 VN.n14 53.8729
R912 VN VN.n23 48.3092
R913 VN.n4 VN.n1 24.3439
R914 VN.n9 VN.n8 24.3439
R915 VN.n16 VN.n13 24.3439
R916 VN.n21 VN.n20 24.3439
R917 VN.n17 VN.n14 17.9272
R918 VN.n5 VN.n2 17.9272
R919 VN.n4 VN.n3 12.1722
R920 VN.n16 VN.n15 12.1722
R921 VN.n10 VN.n9 8.76414
R922 VN.n22 VN.n21 8.76414
R923 VN.n23 VN.n12 0.189894
R924 VN.n19 VN.n12 0.189894
R925 VN.n19 VN.n18 0.189894
R926 VN.n18 VN.n17 0.189894
R927 VN.n6 VN.n5 0.189894
R928 VN.n7 VN.n6 0.189894
R929 VN.n7 VN.n0 0.189894
R930 VN.n11 VN.n0 0.189894
R931 VN VN.n11 0.0516364
R932 VDD2.n175 VDD2.n91 756.745
R933 VDD2.n84 VDD2.n0 756.745
R934 VDD2.n176 VDD2.n175 585
R935 VDD2.n174 VDD2.n173 585
R936 VDD2.n95 VDD2.n94 585
R937 VDD2.n168 VDD2.n167 585
R938 VDD2.n166 VDD2.n97 585
R939 VDD2.n165 VDD2.n164 585
R940 VDD2.n100 VDD2.n98 585
R941 VDD2.n159 VDD2.n158 585
R942 VDD2.n157 VDD2.n156 585
R943 VDD2.n104 VDD2.n103 585
R944 VDD2.n151 VDD2.n150 585
R945 VDD2.n149 VDD2.n148 585
R946 VDD2.n108 VDD2.n107 585
R947 VDD2.n143 VDD2.n142 585
R948 VDD2.n141 VDD2.n140 585
R949 VDD2.n112 VDD2.n111 585
R950 VDD2.n135 VDD2.n134 585
R951 VDD2.n133 VDD2.n132 585
R952 VDD2.n116 VDD2.n115 585
R953 VDD2.n127 VDD2.n126 585
R954 VDD2.n125 VDD2.n124 585
R955 VDD2.n120 VDD2.n119 585
R956 VDD2.n28 VDD2.n27 585
R957 VDD2.n33 VDD2.n32 585
R958 VDD2.n35 VDD2.n34 585
R959 VDD2.n24 VDD2.n23 585
R960 VDD2.n41 VDD2.n40 585
R961 VDD2.n43 VDD2.n42 585
R962 VDD2.n20 VDD2.n19 585
R963 VDD2.n49 VDD2.n48 585
R964 VDD2.n51 VDD2.n50 585
R965 VDD2.n16 VDD2.n15 585
R966 VDD2.n57 VDD2.n56 585
R967 VDD2.n59 VDD2.n58 585
R968 VDD2.n12 VDD2.n11 585
R969 VDD2.n65 VDD2.n64 585
R970 VDD2.n67 VDD2.n66 585
R971 VDD2.n8 VDD2.n7 585
R972 VDD2.n74 VDD2.n73 585
R973 VDD2.n75 VDD2.n6 585
R974 VDD2.n77 VDD2.n76 585
R975 VDD2.n4 VDD2.n3 585
R976 VDD2.n83 VDD2.n82 585
R977 VDD2.n85 VDD2.n84 585
R978 VDD2.n121 VDD2.t5 327.466
R979 VDD2.n29 VDD2.t4 327.466
R980 VDD2.n175 VDD2.n174 171.744
R981 VDD2.n174 VDD2.n94 171.744
R982 VDD2.n167 VDD2.n94 171.744
R983 VDD2.n167 VDD2.n166 171.744
R984 VDD2.n166 VDD2.n165 171.744
R985 VDD2.n165 VDD2.n98 171.744
R986 VDD2.n158 VDD2.n98 171.744
R987 VDD2.n158 VDD2.n157 171.744
R988 VDD2.n157 VDD2.n103 171.744
R989 VDD2.n150 VDD2.n103 171.744
R990 VDD2.n150 VDD2.n149 171.744
R991 VDD2.n149 VDD2.n107 171.744
R992 VDD2.n142 VDD2.n107 171.744
R993 VDD2.n142 VDD2.n141 171.744
R994 VDD2.n141 VDD2.n111 171.744
R995 VDD2.n134 VDD2.n111 171.744
R996 VDD2.n134 VDD2.n133 171.744
R997 VDD2.n133 VDD2.n115 171.744
R998 VDD2.n126 VDD2.n115 171.744
R999 VDD2.n126 VDD2.n125 171.744
R1000 VDD2.n125 VDD2.n119 171.744
R1001 VDD2.n33 VDD2.n27 171.744
R1002 VDD2.n34 VDD2.n33 171.744
R1003 VDD2.n34 VDD2.n23 171.744
R1004 VDD2.n41 VDD2.n23 171.744
R1005 VDD2.n42 VDD2.n41 171.744
R1006 VDD2.n42 VDD2.n19 171.744
R1007 VDD2.n49 VDD2.n19 171.744
R1008 VDD2.n50 VDD2.n49 171.744
R1009 VDD2.n50 VDD2.n15 171.744
R1010 VDD2.n57 VDD2.n15 171.744
R1011 VDD2.n58 VDD2.n57 171.744
R1012 VDD2.n58 VDD2.n11 171.744
R1013 VDD2.n65 VDD2.n11 171.744
R1014 VDD2.n66 VDD2.n65 171.744
R1015 VDD2.n66 VDD2.n7 171.744
R1016 VDD2.n74 VDD2.n7 171.744
R1017 VDD2.n75 VDD2.n74 171.744
R1018 VDD2.n76 VDD2.n75 171.744
R1019 VDD2.n76 VDD2.n3 171.744
R1020 VDD2.n83 VDD2.n3 171.744
R1021 VDD2.n84 VDD2.n83 171.744
R1022 VDD2.t5 VDD2.n119 85.8723
R1023 VDD2.t4 VDD2.n27 85.8723
R1024 VDD2.n90 VDD2.n89 74.0413
R1025 VDD2 VDD2.n181 74.0385
R1026 VDD2.n90 VDD2.n88 53.9354
R1027 VDD2.n180 VDD2.n179 52.7429
R1028 VDD2.n180 VDD2.n90 43.1571
R1029 VDD2.n121 VDD2.n120 16.3895
R1030 VDD2.n29 VDD2.n28 16.3895
R1031 VDD2.n168 VDD2.n97 13.1884
R1032 VDD2.n77 VDD2.n6 13.1884
R1033 VDD2.n169 VDD2.n95 12.8005
R1034 VDD2.n164 VDD2.n99 12.8005
R1035 VDD2.n124 VDD2.n123 12.8005
R1036 VDD2.n32 VDD2.n31 12.8005
R1037 VDD2.n73 VDD2.n72 12.8005
R1038 VDD2.n78 VDD2.n4 12.8005
R1039 VDD2.n173 VDD2.n172 12.0247
R1040 VDD2.n163 VDD2.n100 12.0247
R1041 VDD2.n127 VDD2.n118 12.0247
R1042 VDD2.n35 VDD2.n26 12.0247
R1043 VDD2.n71 VDD2.n8 12.0247
R1044 VDD2.n82 VDD2.n81 12.0247
R1045 VDD2.n176 VDD2.n93 11.249
R1046 VDD2.n160 VDD2.n159 11.249
R1047 VDD2.n128 VDD2.n116 11.249
R1048 VDD2.n36 VDD2.n24 11.249
R1049 VDD2.n68 VDD2.n67 11.249
R1050 VDD2.n85 VDD2.n2 11.249
R1051 VDD2.n177 VDD2.n91 10.4732
R1052 VDD2.n156 VDD2.n102 10.4732
R1053 VDD2.n132 VDD2.n131 10.4732
R1054 VDD2.n40 VDD2.n39 10.4732
R1055 VDD2.n64 VDD2.n10 10.4732
R1056 VDD2.n86 VDD2.n0 10.4732
R1057 VDD2.n155 VDD2.n104 9.69747
R1058 VDD2.n135 VDD2.n114 9.69747
R1059 VDD2.n43 VDD2.n22 9.69747
R1060 VDD2.n63 VDD2.n12 9.69747
R1061 VDD2.n179 VDD2.n178 9.45567
R1062 VDD2.n88 VDD2.n87 9.45567
R1063 VDD2.n147 VDD2.n146 9.3005
R1064 VDD2.n106 VDD2.n105 9.3005
R1065 VDD2.n153 VDD2.n152 9.3005
R1066 VDD2.n155 VDD2.n154 9.3005
R1067 VDD2.n102 VDD2.n101 9.3005
R1068 VDD2.n161 VDD2.n160 9.3005
R1069 VDD2.n163 VDD2.n162 9.3005
R1070 VDD2.n99 VDD2.n96 9.3005
R1071 VDD2.n178 VDD2.n177 9.3005
R1072 VDD2.n93 VDD2.n92 9.3005
R1073 VDD2.n172 VDD2.n171 9.3005
R1074 VDD2.n170 VDD2.n169 9.3005
R1075 VDD2.n145 VDD2.n144 9.3005
R1076 VDD2.n110 VDD2.n109 9.3005
R1077 VDD2.n139 VDD2.n138 9.3005
R1078 VDD2.n137 VDD2.n136 9.3005
R1079 VDD2.n114 VDD2.n113 9.3005
R1080 VDD2.n131 VDD2.n130 9.3005
R1081 VDD2.n129 VDD2.n128 9.3005
R1082 VDD2.n118 VDD2.n117 9.3005
R1083 VDD2.n123 VDD2.n122 9.3005
R1084 VDD2.n87 VDD2.n86 9.3005
R1085 VDD2.n2 VDD2.n1 9.3005
R1086 VDD2.n81 VDD2.n80 9.3005
R1087 VDD2.n79 VDD2.n78 9.3005
R1088 VDD2.n18 VDD2.n17 9.3005
R1089 VDD2.n47 VDD2.n46 9.3005
R1090 VDD2.n45 VDD2.n44 9.3005
R1091 VDD2.n22 VDD2.n21 9.3005
R1092 VDD2.n39 VDD2.n38 9.3005
R1093 VDD2.n37 VDD2.n36 9.3005
R1094 VDD2.n26 VDD2.n25 9.3005
R1095 VDD2.n31 VDD2.n30 9.3005
R1096 VDD2.n53 VDD2.n52 9.3005
R1097 VDD2.n55 VDD2.n54 9.3005
R1098 VDD2.n14 VDD2.n13 9.3005
R1099 VDD2.n61 VDD2.n60 9.3005
R1100 VDD2.n63 VDD2.n62 9.3005
R1101 VDD2.n10 VDD2.n9 9.3005
R1102 VDD2.n69 VDD2.n68 9.3005
R1103 VDD2.n71 VDD2.n70 9.3005
R1104 VDD2.n72 VDD2.n5 9.3005
R1105 VDD2.n152 VDD2.n151 8.92171
R1106 VDD2.n136 VDD2.n112 8.92171
R1107 VDD2.n44 VDD2.n20 8.92171
R1108 VDD2.n60 VDD2.n59 8.92171
R1109 VDD2.n148 VDD2.n106 8.14595
R1110 VDD2.n140 VDD2.n139 8.14595
R1111 VDD2.n48 VDD2.n47 8.14595
R1112 VDD2.n56 VDD2.n14 8.14595
R1113 VDD2.n147 VDD2.n108 7.3702
R1114 VDD2.n143 VDD2.n110 7.3702
R1115 VDD2.n51 VDD2.n18 7.3702
R1116 VDD2.n55 VDD2.n16 7.3702
R1117 VDD2.n144 VDD2.n108 6.59444
R1118 VDD2.n144 VDD2.n143 6.59444
R1119 VDD2.n52 VDD2.n51 6.59444
R1120 VDD2.n52 VDD2.n16 6.59444
R1121 VDD2.n148 VDD2.n147 5.81868
R1122 VDD2.n140 VDD2.n110 5.81868
R1123 VDD2.n48 VDD2.n18 5.81868
R1124 VDD2.n56 VDD2.n55 5.81868
R1125 VDD2.n151 VDD2.n106 5.04292
R1126 VDD2.n139 VDD2.n112 5.04292
R1127 VDD2.n47 VDD2.n20 5.04292
R1128 VDD2.n59 VDD2.n14 5.04292
R1129 VDD2.n152 VDD2.n104 4.26717
R1130 VDD2.n136 VDD2.n135 4.26717
R1131 VDD2.n44 VDD2.n43 4.26717
R1132 VDD2.n60 VDD2.n12 4.26717
R1133 VDD2.n122 VDD2.n121 3.70982
R1134 VDD2.n30 VDD2.n29 3.70982
R1135 VDD2.n179 VDD2.n91 3.49141
R1136 VDD2.n156 VDD2.n155 3.49141
R1137 VDD2.n132 VDD2.n114 3.49141
R1138 VDD2.n40 VDD2.n22 3.49141
R1139 VDD2.n64 VDD2.n63 3.49141
R1140 VDD2.n88 VDD2.n0 3.49141
R1141 VDD2.n177 VDD2.n176 2.71565
R1142 VDD2.n159 VDD2.n102 2.71565
R1143 VDD2.n131 VDD2.n116 2.71565
R1144 VDD2.n39 VDD2.n24 2.71565
R1145 VDD2.n67 VDD2.n10 2.71565
R1146 VDD2.n86 VDD2.n85 2.71565
R1147 VDD2.n181 VDD2.t0 1.99712
R1148 VDD2.n181 VDD2.t3 1.99712
R1149 VDD2.n89 VDD2.t2 1.99712
R1150 VDD2.n89 VDD2.t1 1.99712
R1151 VDD2.n173 VDD2.n93 1.93989
R1152 VDD2.n160 VDD2.n100 1.93989
R1153 VDD2.n128 VDD2.n127 1.93989
R1154 VDD2.n36 VDD2.n35 1.93989
R1155 VDD2.n68 VDD2.n8 1.93989
R1156 VDD2.n82 VDD2.n2 1.93989
R1157 VDD2 VDD2.n180 1.30653
R1158 VDD2.n172 VDD2.n95 1.16414
R1159 VDD2.n164 VDD2.n163 1.16414
R1160 VDD2.n124 VDD2.n118 1.16414
R1161 VDD2.n32 VDD2.n26 1.16414
R1162 VDD2.n73 VDD2.n71 1.16414
R1163 VDD2.n81 VDD2.n4 1.16414
R1164 VDD2.n169 VDD2.n168 0.388379
R1165 VDD2.n99 VDD2.n97 0.388379
R1166 VDD2.n123 VDD2.n120 0.388379
R1167 VDD2.n31 VDD2.n28 0.388379
R1168 VDD2.n72 VDD2.n6 0.388379
R1169 VDD2.n78 VDD2.n77 0.388379
R1170 VDD2.n178 VDD2.n92 0.155672
R1171 VDD2.n171 VDD2.n92 0.155672
R1172 VDD2.n171 VDD2.n170 0.155672
R1173 VDD2.n170 VDD2.n96 0.155672
R1174 VDD2.n162 VDD2.n96 0.155672
R1175 VDD2.n162 VDD2.n161 0.155672
R1176 VDD2.n161 VDD2.n101 0.155672
R1177 VDD2.n154 VDD2.n101 0.155672
R1178 VDD2.n154 VDD2.n153 0.155672
R1179 VDD2.n153 VDD2.n105 0.155672
R1180 VDD2.n146 VDD2.n105 0.155672
R1181 VDD2.n146 VDD2.n145 0.155672
R1182 VDD2.n145 VDD2.n109 0.155672
R1183 VDD2.n138 VDD2.n109 0.155672
R1184 VDD2.n138 VDD2.n137 0.155672
R1185 VDD2.n137 VDD2.n113 0.155672
R1186 VDD2.n130 VDD2.n113 0.155672
R1187 VDD2.n130 VDD2.n129 0.155672
R1188 VDD2.n129 VDD2.n117 0.155672
R1189 VDD2.n122 VDD2.n117 0.155672
R1190 VDD2.n30 VDD2.n25 0.155672
R1191 VDD2.n37 VDD2.n25 0.155672
R1192 VDD2.n38 VDD2.n37 0.155672
R1193 VDD2.n38 VDD2.n21 0.155672
R1194 VDD2.n45 VDD2.n21 0.155672
R1195 VDD2.n46 VDD2.n45 0.155672
R1196 VDD2.n46 VDD2.n17 0.155672
R1197 VDD2.n53 VDD2.n17 0.155672
R1198 VDD2.n54 VDD2.n53 0.155672
R1199 VDD2.n54 VDD2.n13 0.155672
R1200 VDD2.n61 VDD2.n13 0.155672
R1201 VDD2.n62 VDD2.n61 0.155672
R1202 VDD2.n62 VDD2.n9 0.155672
R1203 VDD2.n69 VDD2.n9 0.155672
R1204 VDD2.n70 VDD2.n69 0.155672
R1205 VDD2.n70 VDD2.n5 0.155672
R1206 VDD2.n79 VDD2.n5 0.155672
R1207 VDD2.n80 VDD2.n79 0.155672
R1208 VDD2.n80 VDD2.n1 0.155672
R1209 VDD2.n87 VDD2.n1 0.155672
R1210 B.n510 B.n81 585
R1211 B.n512 B.n511 585
R1212 B.n513 B.n80 585
R1213 B.n515 B.n514 585
R1214 B.n516 B.n79 585
R1215 B.n518 B.n517 585
R1216 B.n519 B.n78 585
R1217 B.n521 B.n520 585
R1218 B.n522 B.n77 585
R1219 B.n524 B.n523 585
R1220 B.n525 B.n76 585
R1221 B.n527 B.n526 585
R1222 B.n528 B.n75 585
R1223 B.n530 B.n529 585
R1224 B.n531 B.n74 585
R1225 B.n533 B.n532 585
R1226 B.n534 B.n73 585
R1227 B.n536 B.n535 585
R1228 B.n537 B.n72 585
R1229 B.n539 B.n538 585
R1230 B.n540 B.n71 585
R1231 B.n542 B.n541 585
R1232 B.n543 B.n70 585
R1233 B.n545 B.n544 585
R1234 B.n546 B.n69 585
R1235 B.n548 B.n547 585
R1236 B.n549 B.n68 585
R1237 B.n551 B.n550 585
R1238 B.n552 B.n67 585
R1239 B.n554 B.n553 585
R1240 B.n555 B.n66 585
R1241 B.n557 B.n556 585
R1242 B.n558 B.n65 585
R1243 B.n560 B.n559 585
R1244 B.n561 B.n64 585
R1245 B.n563 B.n562 585
R1246 B.n564 B.n63 585
R1247 B.n566 B.n565 585
R1248 B.n567 B.n62 585
R1249 B.n569 B.n568 585
R1250 B.n570 B.n61 585
R1251 B.n572 B.n571 585
R1252 B.n573 B.n60 585
R1253 B.n575 B.n574 585
R1254 B.n576 B.n59 585
R1255 B.n578 B.n577 585
R1256 B.n579 B.n58 585
R1257 B.n581 B.n580 585
R1258 B.n582 B.n57 585
R1259 B.n584 B.n583 585
R1260 B.n585 B.n56 585
R1261 B.n587 B.n586 585
R1262 B.n588 B.n55 585
R1263 B.n590 B.n589 585
R1264 B.n592 B.n52 585
R1265 B.n594 B.n593 585
R1266 B.n595 B.n51 585
R1267 B.n597 B.n596 585
R1268 B.n598 B.n50 585
R1269 B.n600 B.n599 585
R1270 B.n601 B.n49 585
R1271 B.n603 B.n602 585
R1272 B.n604 B.n45 585
R1273 B.n606 B.n605 585
R1274 B.n607 B.n44 585
R1275 B.n609 B.n608 585
R1276 B.n610 B.n43 585
R1277 B.n612 B.n611 585
R1278 B.n613 B.n42 585
R1279 B.n615 B.n614 585
R1280 B.n616 B.n41 585
R1281 B.n618 B.n617 585
R1282 B.n619 B.n40 585
R1283 B.n621 B.n620 585
R1284 B.n622 B.n39 585
R1285 B.n624 B.n623 585
R1286 B.n625 B.n38 585
R1287 B.n627 B.n626 585
R1288 B.n628 B.n37 585
R1289 B.n630 B.n629 585
R1290 B.n631 B.n36 585
R1291 B.n633 B.n632 585
R1292 B.n634 B.n35 585
R1293 B.n636 B.n635 585
R1294 B.n637 B.n34 585
R1295 B.n639 B.n638 585
R1296 B.n640 B.n33 585
R1297 B.n642 B.n641 585
R1298 B.n643 B.n32 585
R1299 B.n645 B.n644 585
R1300 B.n646 B.n31 585
R1301 B.n648 B.n647 585
R1302 B.n649 B.n30 585
R1303 B.n651 B.n650 585
R1304 B.n652 B.n29 585
R1305 B.n654 B.n653 585
R1306 B.n655 B.n28 585
R1307 B.n657 B.n656 585
R1308 B.n658 B.n27 585
R1309 B.n660 B.n659 585
R1310 B.n661 B.n26 585
R1311 B.n663 B.n662 585
R1312 B.n664 B.n25 585
R1313 B.n666 B.n665 585
R1314 B.n667 B.n24 585
R1315 B.n669 B.n668 585
R1316 B.n670 B.n23 585
R1317 B.n672 B.n671 585
R1318 B.n673 B.n22 585
R1319 B.n675 B.n674 585
R1320 B.n676 B.n21 585
R1321 B.n678 B.n677 585
R1322 B.n679 B.n20 585
R1323 B.n681 B.n680 585
R1324 B.n682 B.n19 585
R1325 B.n684 B.n683 585
R1326 B.n685 B.n18 585
R1327 B.n687 B.n686 585
R1328 B.n509 B.n508 585
R1329 B.n507 B.n82 585
R1330 B.n506 B.n505 585
R1331 B.n504 B.n83 585
R1332 B.n503 B.n502 585
R1333 B.n501 B.n84 585
R1334 B.n500 B.n499 585
R1335 B.n498 B.n85 585
R1336 B.n497 B.n496 585
R1337 B.n495 B.n86 585
R1338 B.n494 B.n493 585
R1339 B.n492 B.n87 585
R1340 B.n491 B.n490 585
R1341 B.n489 B.n88 585
R1342 B.n488 B.n487 585
R1343 B.n486 B.n89 585
R1344 B.n485 B.n484 585
R1345 B.n483 B.n90 585
R1346 B.n482 B.n481 585
R1347 B.n480 B.n91 585
R1348 B.n479 B.n478 585
R1349 B.n477 B.n92 585
R1350 B.n476 B.n475 585
R1351 B.n474 B.n93 585
R1352 B.n473 B.n472 585
R1353 B.n471 B.n94 585
R1354 B.n470 B.n469 585
R1355 B.n468 B.n95 585
R1356 B.n467 B.n466 585
R1357 B.n465 B.n96 585
R1358 B.n464 B.n463 585
R1359 B.n462 B.n97 585
R1360 B.n461 B.n460 585
R1361 B.n459 B.n98 585
R1362 B.n458 B.n457 585
R1363 B.n456 B.n99 585
R1364 B.n455 B.n454 585
R1365 B.n453 B.n100 585
R1366 B.n452 B.n451 585
R1367 B.n450 B.n101 585
R1368 B.n449 B.n448 585
R1369 B.n447 B.n102 585
R1370 B.n446 B.n445 585
R1371 B.n444 B.n103 585
R1372 B.n443 B.n442 585
R1373 B.n441 B.n104 585
R1374 B.n440 B.n439 585
R1375 B.n438 B.n105 585
R1376 B.n437 B.n436 585
R1377 B.n435 B.n106 585
R1378 B.n434 B.n433 585
R1379 B.n432 B.n107 585
R1380 B.n431 B.n430 585
R1381 B.n429 B.n108 585
R1382 B.n428 B.n427 585
R1383 B.n426 B.n109 585
R1384 B.n425 B.n424 585
R1385 B.n423 B.n110 585
R1386 B.n422 B.n421 585
R1387 B.n420 B.n111 585
R1388 B.n419 B.n418 585
R1389 B.n417 B.n112 585
R1390 B.n416 B.n415 585
R1391 B.n237 B.n176 585
R1392 B.n239 B.n238 585
R1393 B.n240 B.n175 585
R1394 B.n242 B.n241 585
R1395 B.n243 B.n174 585
R1396 B.n245 B.n244 585
R1397 B.n246 B.n173 585
R1398 B.n248 B.n247 585
R1399 B.n249 B.n172 585
R1400 B.n251 B.n250 585
R1401 B.n252 B.n171 585
R1402 B.n254 B.n253 585
R1403 B.n255 B.n170 585
R1404 B.n257 B.n256 585
R1405 B.n258 B.n169 585
R1406 B.n260 B.n259 585
R1407 B.n261 B.n168 585
R1408 B.n263 B.n262 585
R1409 B.n264 B.n167 585
R1410 B.n266 B.n265 585
R1411 B.n267 B.n166 585
R1412 B.n269 B.n268 585
R1413 B.n270 B.n165 585
R1414 B.n272 B.n271 585
R1415 B.n273 B.n164 585
R1416 B.n275 B.n274 585
R1417 B.n276 B.n163 585
R1418 B.n278 B.n277 585
R1419 B.n279 B.n162 585
R1420 B.n281 B.n280 585
R1421 B.n282 B.n161 585
R1422 B.n284 B.n283 585
R1423 B.n285 B.n160 585
R1424 B.n287 B.n286 585
R1425 B.n288 B.n159 585
R1426 B.n290 B.n289 585
R1427 B.n291 B.n158 585
R1428 B.n293 B.n292 585
R1429 B.n294 B.n157 585
R1430 B.n296 B.n295 585
R1431 B.n297 B.n156 585
R1432 B.n299 B.n298 585
R1433 B.n300 B.n155 585
R1434 B.n302 B.n301 585
R1435 B.n303 B.n154 585
R1436 B.n305 B.n304 585
R1437 B.n306 B.n153 585
R1438 B.n308 B.n307 585
R1439 B.n309 B.n152 585
R1440 B.n311 B.n310 585
R1441 B.n312 B.n151 585
R1442 B.n314 B.n313 585
R1443 B.n315 B.n150 585
R1444 B.n317 B.n316 585
R1445 B.n319 B.n318 585
R1446 B.n320 B.n146 585
R1447 B.n322 B.n321 585
R1448 B.n323 B.n145 585
R1449 B.n325 B.n324 585
R1450 B.n326 B.n144 585
R1451 B.n328 B.n327 585
R1452 B.n329 B.n143 585
R1453 B.n331 B.n330 585
R1454 B.n332 B.n140 585
R1455 B.n335 B.n334 585
R1456 B.n336 B.n139 585
R1457 B.n338 B.n337 585
R1458 B.n339 B.n138 585
R1459 B.n341 B.n340 585
R1460 B.n342 B.n137 585
R1461 B.n344 B.n343 585
R1462 B.n345 B.n136 585
R1463 B.n347 B.n346 585
R1464 B.n348 B.n135 585
R1465 B.n350 B.n349 585
R1466 B.n351 B.n134 585
R1467 B.n353 B.n352 585
R1468 B.n354 B.n133 585
R1469 B.n356 B.n355 585
R1470 B.n357 B.n132 585
R1471 B.n359 B.n358 585
R1472 B.n360 B.n131 585
R1473 B.n362 B.n361 585
R1474 B.n363 B.n130 585
R1475 B.n365 B.n364 585
R1476 B.n366 B.n129 585
R1477 B.n368 B.n367 585
R1478 B.n369 B.n128 585
R1479 B.n371 B.n370 585
R1480 B.n372 B.n127 585
R1481 B.n374 B.n373 585
R1482 B.n375 B.n126 585
R1483 B.n377 B.n376 585
R1484 B.n378 B.n125 585
R1485 B.n380 B.n379 585
R1486 B.n381 B.n124 585
R1487 B.n383 B.n382 585
R1488 B.n384 B.n123 585
R1489 B.n386 B.n385 585
R1490 B.n387 B.n122 585
R1491 B.n389 B.n388 585
R1492 B.n390 B.n121 585
R1493 B.n392 B.n391 585
R1494 B.n393 B.n120 585
R1495 B.n395 B.n394 585
R1496 B.n396 B.n119 585
R1497 B.n398 B.n397 585
R1498 B.n399 B.n118 585
R1499 B.n401 B.n400 585
R1500 B.n402 B.n117 585
R1501 B.n404 B.n403 585
R1502 B.n405 B.n116 585
R1503 B.n407 B.n406 585
R1504 B.n408 B.n115 585
R1505 B.n410 B.n409 585
R1506 B.n411 B.n114 585
R1507 B.n413 B.n412 585
R1508 B.n414 B.n113 585
R1509 B.n236 B.n235 585
R1510 B.n234 B.n177 585
R1511 B.n233 B.n232 585
R1512 B.n231 B.n178 585
R1513 B.n230 B.n229 585
R1514 B.n228 B.n179 585
R1515 B.n227 B.n226 585
R1516 B.n225 B.n180 585
R1517 B.n224 B.n223 585
R1518 B.n222 B.n181 585
R1519 B.n221 B.n220 585
R1520 B.n219 B.n182 585
R1521 B.n218 B.n217 585
R1522 B.n216 B.n183 585
R1523 B.n215 B.n214 585
R1524 B.n213 B.n184 585
R1525 B.n212 B.n211 585
R1526 B.n210 B.n185 585
R1527 B.n209 B.n208 585
R1528 B.n207 B.n186 585
R1529 B.n206 B.n205 585
R1530 B.n204 B.n187 585
R1531 B.n203 B.n202 585
R1532 B.n201 B.n188 585
R1533 B.n200 B.n199 585
R1534 B.n198 B.n189 585
R1535 B.n197 B.n196 585
R1536 B.n195 B.n190 585
R1537 B.n194 B.n193 585
R1538 B.n192 B.n191 585
R1539 B.n2 B.n0 585
R1540 B.n733 B.n1 585
R1541 B.n732 B.n731 585
R1542 B.n730 B.n3 585
R1543 B.n729 B.n728 585
R1544 B.n727 B.n4 585
R1545 B.n726 B.n725 585
R1546 B.n724 B.n5 585
R1547 B.n723 B.n722 585
R1548 B.n721 B.n6 585
R1549 B.n720 B.n719 585
R1550 B.n718 B.n7 585
R1551 B.n717 B.n716 585
R1552 B.n715 B.n8 585
R1553 B.n714 B.n713 585
R1554 B.n712 B.n9 585
R1555 B.n711 B.n710 585
R1556 B.n709 B.n10 585
R1557 B.n708 B.n707 585
R1558 B.n706 B.n11 585
R1559 B.n705 B.n704 585
R1560 B.n703 B.n12 585
R1561 B.n702 B.n701 585
R1562 B.n700 B.n13 585
R1563 B.n699 B.n698 585
R1564 B.n697 B.n14 585
R1565 B.n696 B.n695 585
R1566 B.n694 B.n15 585
R1567 B.n693 B.n692 585
R1568 B.n691 B.n16 585
R1569 B.n690 B.n689 585
R1570 B.n688 B.n17 585
R1571 B.n735 B.n734 585
R1572 B.n141 B.t8 490.325
R1573 B.n53 B.t1 490.325
R1574 B.n147 B.t11 490.325
R1575 B.n46 B.t4 490.325
R1576 B.n235 B.n176 468.476
R1577 B.n686 B.n17 468.476
R1578 B.n415 B.n414 468.476
R1579 B.n510 B.n509 468.476
R1580 B.n142 B.t7 452.896
R1581 B.n54 B.t2 452.896
R1582 B.n148 B.t10 452.896
R1583 B.n47 B.t5 452.896
R1584 B.n141 B.t6 451.012
R1585 B.n147 B.t9 451.012
R1586 B.n46 B.t3 451.012
R1587 B.n53 B.t0 451.012
R1588 B.n235 B.n234 163.367
R1589 B.n234 B.n233 163.367
R1590 B.n233 B.n178 163.367
R1591 B.n229 B.n178 163.367
R1592 B.n229 B.n228 163.367
R1593 B.n228 B.n227 163.367
R1594 B.n227 B.n180 163.367
R1595 B.n223 B.n180 163.367
R1596 B.n223 B.n222 163.367
R1597 B.n222 B.n221 163.367
R1598 B.n221 B.n182 163.367
R1599 B.n217 B.n182 163.367
R1600 B.n217 B.n216 163.367
R1601 B.n216 B.n215 163.367
R1602 B.n215 B.n184 163.367
R1603 B.n211 B.n184 163.367
R1604 B.n211 B.n210 163.367
R1605 B.n210 B.n209 163.367
R1606 B.n209 B.n186 163.367
R1607 B.n205 B.n186 163.367
R1608 B.n205 B.n204 163.367
R1609 B.n204 B.n203 163.367
R1610 B.n203 B.n188 163.367
R1611 B.n199 B.n188 163.367
R1612 B.n199 B.n198 163.367
R1613 B.n198 B.n197 163.367
R1614 B.n197 B.n190 163.367
R1615 B.n193 B.n190 163.367
R1616 B.n193 B.n192 163.367
R1617 B.n192 B.n2 163.367
R1618 B.n734 B.n2 163.367
R1619 B.n734 B.n733 163.367
R1620 B.n733 B.n732 163.367
R1621 B.n732 B.n3 163.367
R1622 B.n728 B.n3 163.367
R1623 B.n728 B.n727 163.367
R1624 B.n727 B.n726 163.367
R1625 B.n726 B.n5 163.367
R1626 B.n722 B.n5 163.367
R1627 B.n722 B.n721 163.367
R1628 B.n721 B.n720 163.367
R1629 B.n720 B.n7 163.367
R1630 B.n716 B.n7 163.367
R1631 B.n716 B.n715 163.367
R1632 B.n715 B.n714 163.367
R1633 B.n714 B.n9 163.367
R1634 B.n710 B.n9 163.367
R1635 B.n710 B.n709 163.367
R1636 B.n709 B.n708 163.367
R1637 B.n708 B.n11 163.367
R1638 B.n704 B.n11 163.367
R1639 B.n704 B.n703 163.367
R1640 B.n703 B.n702 163.367
R1641 B.n702 B.n13 163.367
R1642 B.n698 B.n13 163.367
R1643 B.n698 B.n697 163.367
R1644 B.n697 B.n696 163.367
R1645 B.n696 B.n15 163.367
R1646 B.n692 B.n15 163.367
R1647 B.n692 B.n691 163.367
R1648 B.n691 B.n690 163.367
R1649 B.n690 B.n17 163.367
R1650 B.n239 B.n176 163.367
R1651 B.n240 B.n239 163.367
R1652 B.n241 B.n240 163.367
R1653 B.n241 B.n174 163.367
R1654 B.n245 B.n174 163.367
R1655 B.n246 B.n245 163.367
R1656 B.n247 B.n246 163.367
R1657 B.n247 B.n172 163.367
R1658 B.n251 B.n172 163.367
R1659 B.n252 B.n251 163.367
R1660 B.n253 B.n252 163.367
R1661 B.n253 B.n170 163.367
R1662 B.n257 B.n170 163.367
R1663 B.n258 B.n257 163.367
R1664 B.n259 B.n258 163.367
R1665 B.n259 B.n168 163.367
R1666 B.n263 B.n168 163.367
R1667 B.n264 B.n263 163.367
R1668 B.n265 B.n264 163.367
R1669 B.n265 B.n166 163.367
R1670 B.n269 B.n166 163.367
R1671 B.n270 B.n269 163.367
R1672 B.n271 B.n270 163.367
R1673 B.n271 B.n164 163.367
R1674 B.n275 B.n164 163.367
R1675 B.n276 B.n275 163.367
R1676 B.n277 B.n276 163.367
R1677 B.n277 B.n162 163.367
R1678 B.n281 B.n162 163.367
R1679 B.n282 B.n281 163.367
R1680 B.n283 B.n282 163.367
R1681 B.n283 B.n160 163.367
R1682 B.n287 B.n160 163.367
R1683 B.n288 B.n287 163.367
R1684 B.n289 B.n288 163.367
R1685 B.n289 B.n158 163.367
R1686 B.n293 B.n158 163.367
R1687 B.n294 B.n293 163.367
R1688 B.n295 B.n294 163.367
R1689 B.n295 B.n156 163.367
R1690 B.n299 B.n156 163.367
R1691 B.n300 B.n299 163.367
R1692 B.n301 B.n300 163.367
R1693 B.n301 B.n154 163.367
R1694 B.n305 B.n154 163.367
R1695 B.n306 B.n305 163.367
R1696 B.n307 B.n306 163.367
R1697 B.n307 B.n152 163.367
R1698 B.n311 B.n152 163.367
R1699 B.n312 B.n311 163.367
R1700 B.n313 B.n312 163.367
R1701 B.n313 B.n150 163.367
R1702 B.n317 B.n150 163.367
R1703 B.n318 B.n317 163.367
R1704 B.n318 B.n146 163.367
R1705 B.n322 B.n146 163.367
R1706 B.n323 B.n322 163.367
R1707 B.n324 B.n323 163.367
R1708 B.n324 B.n144 163.367
R1709 B.n328 B.n144 163.367
R1710 B.n329 B.n328 163.367
R1711 B.n330 B.n329 163.367
R1712 B.n330 B.n140 163.367
R1713 B.n335 B.n140 163.367
R1714 B.n336 B.n335 163.367
R1715 B.n337 B.n336 163.367
R1716 B.n337 B.n138 163.367
R1717 B.n341 B.n138 163.367
R1718 B.n342 B.n341 163.367
R1719 B.n343 B.n342 163.367
R1720 B.n343 B.n136 163.367
R1721 B.n347 B.n136 163.367
R1722 B.n348 B.n347 163.367
R1723 B.n349 B.n348 163.367
R1724 B.n349 B.n134 163.367
R1725 B.n353 B.n134 163.367
R1726 B.n354 B.n353 163.367
R1727 B.n355 B.n354 163.367
R1728 B.n355 B.n132 163.367
R1729 B.n359 B.n132 163.367
R1730 B.n360 B.n359 163.367
R1731 B.n361 B.n360 163.367
R1732 B.n361 B.n130 163.367
R1733 B.n365 B.n130 163.367
R1734 B.n366 B.n365 163.367
R1735 B.n367 B.n366 163.367
R1736 B.n367 B.n128 163.367
R1737 B.n371 B.n128 163.367
R1738 B.n372 B.n371 163.367
R1739 B.n373 B.n372 163.367
R1740 B.n373 B.n126 163.367
R1741 B.n377 B.n126 163.367
R1742 B.n378 B.n377 163.367
R1743 B.n379 B.n378 163.367
R1744 B.n379 B.n124 163.367
R1745 B.n383 B.n124 163.367
R1746 B.n384 B.n383 163.367
R1747 B.n385 B.n384 163.367
R1748 B.n385 B.n122 163.367
R1749 B.n389 B.n122 163.367
R1750 B.n390 B.n389 163.367
R1751 B.n391 B.n390 163.367
R1752 B.n391 B.n120 163.367
R1753 B.n395 B.n120 163.367
R1754 B.n396 B.n395 163.367
R1755 B.n397 B.n396 163.367
R1756 B.n397 B.n118 163.367
R1757 B.n401 B.n118 163.367
R1758 B.n402 B.n401 163.367
R1759 B.n403 B.n402 163.367
R1760 B.n403 B.n116 163.367
R1761 B.n407 B.n116 163.367
R1762 B.n408 B.n407 163.367
R1763 B.n409 B.n408 163.367
R1764 B.n409 B.n114 163.367
R1765 B.n413 B.n114 163.367
R1766 B.n414 B.n413 163.367
R1767 B.n415 B.n112 163.367
R1768 B.n419 B.n112 163.367
R1769 B.n420 B.n419 163.367
R1770 B.n421 B.n420 163.367
R1771 B.n421 B.n110 163.367
R1772 B.n425 B.n110 163.367
R1773 B.n426 B.n425 163.367
R1774 B.n427 B.n426 163.367
R1775 B.n427 B.n108 163.367
R1776 B.n431 B.n108 163.367
R1777 B.n432 B.n431 163.367
R1778 B.n433 B.n432 163.367
R1779 B.n433 B.n106 163.367
R1780 B.n437 B.n106 163.367
R1781 B.n438 B.n437 163.367
R1782 B.n439 B.n438 163.367
R1783 B.n439 B.n104 163.367
R1784 B.n443 B.n104 163.367
R1785 B.n444 B.n443 163.367
R1786 B.n445 B.n444 163.367
R1787 B.n445 B.n102 163.367
R1788 B.n449 B.n102 163.367
R1789 B.n450 B.n449 163.367
R1790 B.n451 B.n450 163.367
R1791 B.n451 B.n100 163.367
R1792 B.n455 B.n100 163.367
R1793 B.n456 B.n455 163.367
R1794 B.n457 B.n456 163.367
R1795 B.n457 B.n98 163.367
R1796 B.n461 B.n98 163.367
R1797 B.n462 B.n461 163.367
R1798 B.n463 B.n462 163.367
R1799 B.n463 B.n96 163.367
R1800 B.n467 B.n96 163.367
R1801 B.n468 B.n467 163.367
R1802 B.n469 B.n468 163.367
R1803 B.n469 B.n94 163.367
R1804 B.n473 B.n94 163.367
R1805 B.n474 B.n473 163.367
R1806 B.n475 B.n474 163.367
R1807 B.n475 B.n92 163.367
R1808 B.n479 B.n92 163.367
R1809 B.n480 B.n479 163.367
R1810 B.n481 B.n480 163.367
R1811 B.n481 B.n90 163.367
R1812 B.n485 B.n90 163.367
R1813 B.n486 B.n485 163.367
R1814 B.n487 B.n486 163.367
R1815 B.n487 B.n88 163.367
R1816 B.n491 B.n88 163.367
R1817 B.n492 B.n491 163.367
R1818 B.n493 B.n492 163.367
R1819 B.n493 B.n86 163.367
R1820 B.n497 B.n86 163.367
R1821 B.n498 B.n497 163.367
R1822 B.n499 B.n498 163.367
R1823 B.n499 B.n84 163.367
R1824 B.n503 B.n84 163.367
R1825 B.n504 B.n503 163.367
R1826 B.n505 B.n504 163.367
R1827 B.n505 B.n82 163.367
R1828 B.n509 B.n82 163.367
R1829 B.n686 B.n685 163.367
R1830 B.n685 B.n684 163.367
R1831 B.n684 B.n19 163.367
R1832 B.n680 B.n19 163.367
R1833 B.n680 B.n679 163.367
R1834 B.n679 B.n678 163.367
R1835 B.n678 B.n21 163.367
R1836 B.n674 B.n21 163.367
R1837 B.n674 B.n673 163.367
R1838 B.n673 B.n672 163.367
R1839 B.n672 B.n23 163.367
R1840 B.n668 B.n23 163.367
R1841 B.n668 B.n667 163.367
R1842 B.n667 B.n666 163.367
R1843 B.n666 B.n25 163.367
R1844 B.n662 B.n25 163.367
R1845 B.n662 B.n661 163.367
R1846 B.n661 B.n660 163.367
R1847 B.n660 B.n27 163.367
R1848 B.n656 B.n27 163.367
R1849 B.n656 B.n655 163.367
R1850 B.n655 B.n654 163.367
R1851 B.n654 B.n29 163.367
R1852 B.n650 B.n29 163.367
R1853 B.n650 B.n649 163.367
R1854 B.n649 B.n648 163.367
R1855 B.n648 B.n31 163.367
R1856 B.n644 B.n31 163.367
R1857 B.n644 B.n643 163.367
R1858 B.n643 B.n642 163.367
R1859 B.n642 B.n33 163.367
R1860 B.n638 B.n33 163.367
R1861 B.n638 B.n637 163.367
R1862 B.n637 B.n636 163.367
R1863 B.n636 B.n35 163.367
R1864 B.n632 B.n35 163.367
R1865 B.n632 B.n631 163.367
R1866 B.n631 B.n630 163.367
R1867 B.n630 B.n37 163.367
R1868 B.n626 B.n37 163.367
R1869 B.n626 B.n625 163.367
R1870 B.n625 B.n624 163.367
R1871 B.n624 B.n39 163.367
R1872 B.n620 B.n39 163.367
R1873 B.n620 B.n619 163.367
R1874 B.n619 B.n618 163.367
R1875 B.n618 B.n41 163.367
R1876 B.n614 B.n41 163.367
R1877 B.n614 B.n613 163.367
R1878 B.n613 B.n612 163.367
R1879 B.n612 B.n43 163.367
R1880 B.n608 B.n43 163.367
R1881 B.n608 B.n607 163.367
R1882 B.n607 B.n606 163.367
R1883 B.n606 B.n45 163.367
R1884 B.n602 B.n45 163.367
R1885 B.n602 B.n601 163.367
R1886 B.n601 B.n600 163.367
R1887 B.n600 B.n50 163.367
R1888 B.n596 B.n50 163.367
R1889 B.n596 B.n595 163.367
R1890 B.n595 B.n594 163.367
R1891 B.n594 B.n52 163.367
R1892 B.n589 B.n52 163.367
R1893 B.n589 B.n588 163.367
R1894 B.n588 B.n587 163.367
R1895 B.n587 B.n56 163.367
R1896 B.n583 B.n56 163.367
R1897 B.n583 B.n582 163.367
R1898 B.n582 B.n581 163.367
R1899 B.n581 B.n58 163.367
R1900 B.n577 B.n58 163.367
R1901 B.n577 B.n576 163.367
R1902 B.n576 B.n575 163.367
R1903 B.n575 B.n60 163.367
R1904 B.n571 B.n60 163.367
R1905 B.n571 B.n570 163.367
R1906 B.n570 B.n569 163.367
R1907 B.n569 B.n62 163.367
R1908 B.n565 B.n62 163.367
R1909 B.n565 B.n564 163.367
R1910 B.n564 B.n563 163.367
R1911 B.n563 B.n64 163.367
R1912 B.n559 B.n64 163.367
R1913 B.n559 B.n558 163.367
R1914 B.n558 B.n557 163.367
R1915 B.n557 B.n66 163.367
R1916 B.n553 B.n66 163.367
R1917 B.n553 B.n552 163.367
R1918 B.n552 B.n551 163.367
R1919 B.n551 B.n68 163.367
R1920 B.n547 B.n68 163.367
R1921 B.n547 B.n546 163.367
R1922 B.n546 B.n545 163.367
R1923 B.n545 B.n70 163.367
R1924 B.n541 B.n70 163.367
R1925 B.n541 B.n540 163.367
R1926 B.n540 B.n539 163.367
R1927 B.n539 B.n72 163.367
R1928 B.n535 B.n72 163.367
R1929 B.n535 B.n534 163.367
R1930 B.n534 B.n533 163.367
R1931 B.n533 B.n74 163.367
R1932 B.n529 B.n74 163.367
R1933 B.n529 B.n528 163.367
R1934 B.n528 B.n527 163.367
R1935 B.n527 B.n76 163.367
R1936 B.n523 B.n76 163.367
R1937 B.n523 B.n522 163.367
R1938 B.n522 B.n521 163.367
R1939 B.n521 B.n78 163.367
R1940 B.n517 B.n78 163.367
R1941 B.n517 B.n516 163.367
R1942 B.n516 B.n515 163.367
R1943 B.n515 B.n80 163.367
R1944 B.n511 B.n80 163.367
R1945 B.n511 B.n510 163.367
R1946 B.n333 B.n142 59.5399
R1947 B.n149 B.n148 59.5399
R1948 B.n48 B.n47 59.5399
R1949 B.n591 B.n54 59.5399
R1950 B.n142 B.n141 37.4308
R1951 B.n148 B.n147 37.4308
R1952 B.n47 B.n46 37.4308
R1953 B.n54 B.n53 37.4308
R1954 B.n688 B.n687 30.4395
R1955 B.n416 B.n113 30.4395
R1956 B.n237 B.n236 30.4395
R1957 B.n508 B.n81 30.4395
R1958 B B.n735 18.0485
R1959 B.n687 B.n18 10.6151
R1960 B.n683 B.n18 10.6151
R1961 B.n683 B.n682 10.6151
R1962 B.n682 B.n681 10.6151
R1963 B.n681 B.n20 10.6151
R1964 B.n677 B.n20 10.6151
R1965 B.n677 B.n676 10.6151
R1966 B.n676 B.n675 10.6151
R1967 B.n675 B.n22 10.6151
R1968 B.n671 B.n22 10.6151
R1969 B.n671 B.n670 10.6151
R1970 B.n670 B.n669 10.6151
R1971 B.n669 B.n24 10.6151
R1972 B.n665 B.n24 10.6151
R1973 B.n665 B.n664 10.6151
R1974 B.n664 B.n663 10.6151
R1975 B.n663 B.n26 10.6151
R1976 B.n659 B.n26 10.6151
R1977 B.n659 B.n658 10.6151
R1978 B.n658 B.n657 10.6151
R1979 B.n657 B.n28 10.6151
R1980 B.n653 B.n28 10.6151
R1981 B.n653 B.n652 10.6151
R1982 B.n652 B.n651 10.6151
R1983 B.n651 B.n30 10.6151
R1984 B.n647 B.n30 10.6151
R1985 B.n647 B.n646 10.6151
R1986 B.n646 B.n645 10.6151
R1987 B.n645 B.n32 10.6151
R1988 B.n641 B.n32 10.6151
R1989 B.n641 B.n640 10.6151
R1990 B.n640 B.n639 10.6151
R1991 B.n639 B.n34 10.6151
R1992 B.n635 B.n34 10.6151
R1993 B.n635 B.n634 10.6151
R1994 B.n634 B.n633 10.6151
R1995 B.n633 B.n36 10.6151
R1996 B.n629 B.n36 10.6151
R1997 B.n629 B.n628 10.6151
R1998 B.n628 B.n627 10.6151
R1999 B.n627 B.n38 10.6151
R2000 B.n623 B.n38 10.6151
R2001 B.n623 B.n622 10.6151
R2002 B.n622 B.n621 10.6151
R2003 B.n621 B.n40 10.6151
R2004 B.n617 B.n40 10.6151
R2005 B.n617 B.n616 10.6151
R2006 B.n616 B.n615 10.6151
R2007 B.n615 B.n42 10.6151
R2008 B.n611 B.n42 10.6151
R2009 B.n611 B.n610 10.6151
R2010 B.n610 B.n609 10.6151
R2011 B.n609 B.n44 10.6151
R2012 B.n605 B.n604 10.6151
R2013 B.n604 B.n603 10.6151
R2014 B.n603 B.n49 10.6151
R2015 B.n599 B.n49 10.6151
R2016 B.n599 B.n598 10.6151
R2017 B.n598 B.n597 10.6151
R2018 B.n597 B.n51 10.6151
R2019 B.n593 B.n51 10.6151
R2020 B.n593 B.n592 10.6151
R2021 B.n590 B.n55 10.6151
R2022 B.n586 B.n55 10.6151
R2023 B.n586 B.n585 10.6151
R2024 B.n585 B.n584 10.6151
R2025 B.n584 B.n57 10.6151
R2026 B.n580 B.n57 10.6151
R2027 B.n580 B.n579 10.6151
R2028 B.n579 B.n578 10.6151
R2029 B.n578 B.n59 10.6151
R2030 B.n574 B.n59 10.6151
R2031 B.n574 B.n573 10.6151
R2032 B.n573 B.n572 10.6151
R2033 B.n572 B.n61 10.6151
R2034 B.n568 B.n61 10.6151
R2035 B.n568 B.n567 10.6151
R2036 B.n567 B.n566 10.6151
R2037 B.n566 B.n63 10.6151
R2038 B.n562 B.n63 10.6151
R2039 B.n562 B.n561 10.6151
R2040 B.n561 B.n560 10.6151
R2041 B.n560 B.n65 10.6151
R2042 B.n556 B.n65 10.6151
R2043 B.n556 B.n555 10.6151
R2044 B.n555 B.n554 10.6151
R2045 B.n554 B.n67 10.6151
R2046 B.n550 B.n67 10.6151
R2047 B.n550 B.n549 10.6151
R2048 B.n549 B.n548 10.6151
R2049 B.n548 B.n69 10.6151
R2050 B.n544 B.n69 10.6151
R2051 B.n544 B.n543 10.6151
R2052 B.n543 B.n542 10.6151
R2053 B.n542 B.n71 10.6151
R2054 B.n538 B.n71 10.6151
R2055 B.n538 B.n537 10.6151
R2056 B.n537 B.n536 10.6151
R2057 B.n536 B.n73 10.6151
R2058 B.n532 B.n73 10.6151
R2059 B.n532 B.n531 10.6151
R2060 B.n531 B.n530 10.6151
R2061 B.n530 B.n75 10.6151
R2062 B.n526 B.n75 10.6151
R2063 B.n526 B.n525 10.6151
R2064 B.n525 B.n524 10.6151
R2065 B.n524 B.n77 10.6151
R2066 B.n520 B.n77 10.6151
R2067 B.n520 B.n519 10.6151
R2068 B.n519 B.n518 10.6151
R2069 B.n518 B.n79 10.6151
R2070 B.n514 B.n79 10.6151
R2071 B.n514 B.n513 10.6151
R2072 B.n513 B.n512 10.6151
R2073 B.n512 B.n81 10.6151
R2074 B.n417 B.n416 10.6151
R2075 B.n418 B.n417 10.6151
R2076 B.n418 B.n111 10.6151
R2077 B.n422 B.n111 10.6151
R2078 B.n423 B.n422 10.6151
R2079 B.n424 B.n423 10.6151
R2080 B.n424 B.n109 10.6151
R2081 B.n428 B.n109 10.6151
R2082 B.n429 B.n428 10.6151
R2083 B.n430 B.n429 10.6151
R2084 B.n430 B.n107 10.6151
R2085 B.n434 B.n107 10.6151
R2086 B.n435 B.n434 10.6151
R2087 B.n436 B.n435 10.6151
R2088 B.n436 B.n105 10.6151
R2089 B.n440 B.n105 10.6151
R2090 B.n441 B.n440 10.6151
R2091 B.n442 B.n441 10.6151
R2092 B.n442 B.n103 10.6151
R2093 B.n446 B.n103 10.6151
R2094 B.n447 B.n446 10.6151
R2095 B.n448 B.n447 10.6151
R2096 B.n448 B.n101 10.6151
R2097 B.n452 B.n101 10.6151
R2098 B.n453 B.n452 10.6151
R2099 B.n454 B.n453 10.6151
R2100 B.n454 B.n99 10.6151
R2101 B.n458 B.n99 10.6151
R2102 B.n459 B.n458 10.6151
R2103 B.n460 B.n459 10.6151
R2104 B.n460 B.n97 10.6151
R2105 B.n464 B.n97 10.6151
R2106 B.n465 B.n464 10.6151
R2107 B.n466 B.n465 10.6151
R2108 B.n466 B.n95 10.6151
R2109 B.n470 B.n95 10.6151
R2110 B.n471 B.n470 10.6151
R2111 B.n472 B.n471 10.6151
R2112 B.n472 B.n93 10.6151
R2113 B.n476 B.n93 10.6151
R2114 B.n477 B.n476 10.6151
R2115 B.n478 B.n477 10.6151
R2116 B.n478 B.n91 10.6151
R2117 B.n482 B.n91 10.6151
R2118 B.n483 B.n482 10.6151
R2119 B.n484 B.n483 10.6151
R2120 B.n484 B.n89 10.6151
R2121 B.n488 B.n89 10.6151
R2122 B.n489 B.n488 10.6151
R2123 B.n490 B.n489 10.6151
R2124 B.n490 B.n87 10.6151
R2125 B.n494 B.n87 10.6151
R2126 B.n495 B.n494 10.6151
R2127 B.n496 B.n495 10.6151
R2128 B.n496 B.n85 10.6151
R2129 B.n500 B.n85 10.6151
R2130 B.n501 B.n500 10.6151
R2131 B.n502 B.n501 10.6151
R2132 B.n502 B.n83 10.6151
R2133 B.n506 B.n83 10.6151
R2134 B.n507 B.n506 10.6151
R2135 B.n508 B.n507 10.6151
R2136 B.n238 B.n237 10.6151
R2137 B.n238 B.n175 10.6151
R2138 B.n242 B.n175 10.6151
R2139 B.n243 B.n242 10.6151
R2140 B.n244 B.n243 10.6151
R2141 B.n244 B.n173 10.6151
R2142 B.n248 B.n173 10.6151
R2143 B.n249 B.n248 10.6151
R2144 B.n250 B.n249 10.6151
R2145 B.n250 B.n171 10.6151
R2146 B.n254 B.n171 10.6151
R2147 B.n255 B.n254 10.6151
R2148 B.n256 B.n255 10.6151
R2149 B.n256 B.n169 10.6151
R2150 B.n260 B.n169 10.6151
R2151 B.n261 B.n260 10.6151
R2152 B.n262 B.n261 10.6151
R2153 B.n262 B.n167 10.6151
R2154 B.n266 B.n167 10.6151
R2155 B.n267 B.n266 10.6151
R2156 B.n268 B.n267 10.6151
R2157 B.n268 B.n165 10.6151
R2158 B.n272 B.n165 10.6151
R2159 B.n273 B.n272 10.6151
R2160 B.n274 B.n273 10.6151
R2161 B.n274 B.n163 10.6151
R2162 B.n278 B.n163 10.6151
R2163 B.n279 B.n278 10.6151
R2164 B.n280 B.n279 10.6151
R2165 B.n280 B.n161 10.6151
R2166 B.n284 B.n161 10.6151
R2167 B.n285 B.n284 10.6151
R2168 B.n286 B.n285 10.6151
R2169 B.n286 B.n159 10.6151
R2170 B.n290 B.n159 10.6151
R2171 B.n291 B.n290 10.6151
R2172 B.n292 B.n291 10.6151
R2173 B.n292 B.n157 10.6151
R2174 B.n296 B.n157 10.6151
R2175 B.n297 B.n296 10.6151
R2176 B.n298 B.n297 10.6151
R2177 B.n298 B.n155 10.6151
R2178 B.n302 B.n155 10.6151
R2179 B.n303 B.n302 10.6151
R2180 B.n304 B.n303 10.6151
R2181 B.n304 B.n153 10.6151
R2182 B.n308 B.n153 10.6151
R2183 B.n309 B.n308 10.6151
R2184 B.n310 B.n309 10.6151
R2185 B.n310 B.n151 10.6151
R2186 B.n314 B.n151 10.6151
R2187 B.n315 B.n314 10.6151
R2188 B.n316 B.n315 10.6151
R2189 B.n320 B.n319 10.6151
R2190 B.n321 B.n320 10.6151
R2191 B.n321 B.n145 10.6151
R2192 B.n325 B.n145 10.6151
R2193 B.n326 B.n325 10.6151
R2194 B.n327 B.n326 10.6151
R2195 B.n327 B.n143 10.6151
R2196 B.n331 B.n143 10.6151
R2197 B.n332 B.n331 10.6151
R2198 B.n334 B.n139 10.6151
R2199 B.n338 B.n139 10.6151
R2200 B.n339 B.n338 10.6151
R2201 B.n340 B.n339 10.6151
R2202 B.n340 B.n137 10.6151
R2203 B.n344 B.n137 10.6151
R2204 B.n345 B.n344 10.6151
R2205 B.n346 B.n345 10.6151
R2206 B.n346 B.n135 10.6151
R2207 B.n350 B.n135 10.6151
R2208 B.n351 B.n350 10.6151
R2209 B.n352 B.n351 10.6151
R2210 B.n352 B.n133 10.6151
R2211 B.n356 B.n133 10.6151
R2212 B.n357 B.n356 10.6151
R2213 B.n358 B.n357 10.6151
R2214 B.n358 B.n131 10.6151
R2215 B.n362 B.n131 10.6151
R2216 B.n363 B.n362 10.6151
R2217 B.n364 B.n363 10.6151
R2218 B.n364 B.n129 10.6151
R2219 B.n368 B.n129 10.6151
R2220 B.n369 B.n368 10.6151
R2221 B.n370 B.n369 10.6151
R2222 B.n370 B.n127 10.6151
R2223 B.n374 B.n127 10.6151
R2224 B.n375 B.n374 10.6151
R2225 B.n376 B.n375 10.6151
R2226 B.n376 B.n125 10.6151
R2227 B.n380 B.n125 10.6151
R2228 B.n381 B.n380 10.6151
R2229 B.n382 B.n381 10.6151
R2230 B.n382 B.n123 10.6151
R2231 B.n386 B.n123 10.6151
R2232 B.n387 B.n386 10.6151
R2233 B.n388 B.n387 10.6151
R2234 B.n388 B.n121 10.6151
R2235 B.n392 B.n121 10.6151
R2236 B.n393 B.n392 10.6151
R2237 B.n394 B.n393 10.6151
R2238 B.n394 B.n119 10.6151
R2239 B.n398 B.n119 10.6151
R2240 B.n399 B.n398 10.6151
R2241 B.n400 B.n399 10.6151
R2242 B.n400 B.n117 10.6151
R2243 B.n404 B.n117 10.6151
R2244 B.n405 B.n404 10.6151
R2245 B.n406 B.n405 10.6151
R2246 B.n406 B.n115 10.6151
R2247 B.n410 B.n115 10.6151
R2248 B.n411 B.n410 10.6151
R2249 B.n412 B.n411 10.6151
R2250 B.n412 B.n113 10.6151
R2251 B.n236 B.n177 10.6151
R2252 B.n232 B.n177 10.6151
R2253 B.n232 B.n231 10.6151
R2254 B.n231 B.n230 10.6151
R2255 B.n230 B.n179 10.6151
R2256 B.n226 B.n179 10.6151
R2257 B.n226 B.n225 10.6151
R2258 B.n225 B.n224 10.6151
R2259 B.n224 B.n181 10.6151
R2260 B.n220 B.n181 10.6151
R2261 B.n220 B.n219 10.6151
R2262 B.n219 B.n218 10.6151
R2263 B.n218 B.n183 10.6151
R2264 B.n214 B.n183 10.6151
R2265 B.n214 B.n213 10.6151
R2266 B.n213 B.n212 10.6151
R2267 B.n212 B.n185 10.6151
R2268 B.n208 B.n185 10.6151
R2269 B.n208 B.n207 10.6151
R2270 B.n207 B.n206 10.6151
R2271 B.n206 B.n187 10.6151
R2272 B.n202 B.n187 10.6151
R2273 B.n202 B.n201 10.6151
R2274 B.n201 B.n200 10.6151
R2275 B.n200 B.n189 10.6151
R2276 B.n196 B.n189 10.6151
R2277 B.n196 B.n195 10.6151
R2278 B.n195 B.n194 10.6151
R2279 B.n194 B.n191 10.6151
R2280 B.n191 B.n0 10.6151
R2281 B.n731 B.n1 10.6151
R2282 B.n731 B.n730 10.6151
R2283 B.n730 B.n729 10.6151
R2284 B.n729 B.n4 10.6151
R2285 B.n725 B.n4 10.6151
R2286 B.n725 B.n724 10.6151
R2287 B.n724 B.n723 10.6151
R2288 B.n723 B.n6 10.6151
R2289 B.n719 B.n6 10.6151
R2290 B.n719 B.n718 10.6151
R2291 B.n718 B.n717 10.6151
R2292 B.n717 B.n8 10.6151
R2293 B.n713 B.n8 10.6151
R2294 B.n713 B.n712 10.6151
R2295 B.n712 B.n711 10.6151
R2296 B.n711 B.n10 10.6151
R2297 B.n707 B.n10 10.6151
R2298 B.n707 B.n706 10.6151
R2299 B.n706 B.n705 10.6151
R2300 B.n705 B.n12 10.6151
R2301 B.n701 B.n12 10.6151
R2302 B.n701 B.n700 10.6151
R2303 B.n700 B.n699 10.6151
R2304 B.n699 B.n14 10.6151
R2305 B.n695 B.n14 10.6151
R2306 B.n695 B.n694 10.6151
R2307 B.n694 B.n693 10.6151
R2308 B.n693 B.n16 10.6151
R2309 B.n689 B.n16 10.6151
R2310 B.n689 B.n688 10.6151
R2311 B.n48 B.n44 9.36635
R2312 B.n591 B.n590 9.36635
R2313 B.n316 B.n149 9.36635
R2314 B.n334 B.n333 9.36635
R2315 B.n735 B.n0 2.81026
R2316 B.n735 B.n1 2.81026
R2317 B.n605 B.n48 1.24928
R2318 B.n592 B.n591 1.24928
R2319 B.n319 B.n149 1.24928
R2320 B.n333 B.n332 1.24928
C0 VDD1 VN 0.149107f
C1 VN VTAIL 7.747721f
C2 VDD1 B 2.15064f
C3 VDD2 VN 7.99746f
C4 VTAIL B 4.11347f
C5 VDD2 B 2.20084f
C6 VDD1 VP 8.21753f
C7 w_n2514_n4224# VDD1 2.35154f
C8 VTAIL VP 7.76223f
C9 w_n2514_n4224# VTAIL 3.53792f
C10 VN B 1.00293f
C11 VDD2 VP 0.373844f
C12 w_n2514_n4224# VDD2 2.40451f
C13 VN VP 6.75032f
C14 w_n2514_n4224# VN 4.60055f
C15 B VP 1.53591f
C16 w_n2514_n4224# B 9.49522f
C17 w_n2514_n4224# VP 4.92279f
C18 VDD1 VTAIL 9.814569f
C19 VDD1 VDD2 1.04611f
C20 VDD2 VTAIL 9.85572f
C21 VDD2 VSUBS 1.753146f
C22 VDD1 VSUBS 1.596699f
C23 VTAIL VSUBS 1.143023f
C24 VN VSUBS 5.1837f
C25 VP VSUBS 2.309098f
C26 B VSUBS 4.012077f
C27 w_n2514_n4224# VSUBS 0.130054p
C28 B.n0 VSUBS 0.005155f
C29 B.n1 VSUBS 0.005155f
C30 B.n2 VSUBS 0.008152f
C31 B.n3 VSUBS 0.008152f
C32 B.n4 VSUBS 0.008152f
C33 B.n5 VSUBS 0.008152f
C34 B.n6 VSUBS 0.008152f
C35 B.n7 VSUBS 0.008152f
C36 B.n8 VSUBS 0.008152f
C37 B.n9 VSUBS 0.008152f
C38 B.n10 VSUBS 0.008152f
C39 B.n11 VSUBS 0.008152f
C40 B.n12 VSUBS 0.008152f
C41 B.n13 VSUBS 0.008152f
C42 B.n14 VSUBS 0.008152f
C43 B.n15 VSUBS 0.008152f
C44 B.n16 VSUBS 0.008152f
C45 B.n17 VSUBS 0.017883f
C46 B.n18 VSUBS 0.008152f
C47 B.n19 VSUBS 0.008152f
C48 B.n20 VSUBS 0.008152f
C49 B.n21 VSUBS 0.008152f
C50 B.n22 VSUBS 0.008152f
C51 B.n23 VSUBS 0.008152f
C52 B.n24 VSUBS 0.008152f
C53 B.n25 VSUBS 0.008152f
C54 B.n26 VSUBS 0.008152f
C55 B.n27 VSUBS 0.008152f
C56 B.n28 VSUBS 0.008152f
C57 B.n29 VSUBS 0.008152f
C58 B.n30 VSUBS 0.008152f
C59 B.n31 VSUBS 0.008152f
C60 B.n32 VSUBS 0.008152f
C61 B.n33 VSUBS 0.008152f
C62 B.n34 VSUBS 0.008152f
C63 B.n35 VSUBS 0.008152f
C64 B.n36 VSUBS 0.008152f
C65 B.n37 VSUBS 0.008152f
C66 B.n38 VSUBS 0.008152f
C67 B.n39 VSUBS 0.008152f
C68 B.n40 VSUBS 0.008152f
C69 B.n41 VSUBS 0.008152f
C70 B.n42 VSUBS 0.008152f
C71 B.n43 VSUBS 0.008152f
C72 B.n44 VSUBS 0.007673f
C73 B.n45 VSUBS 0.008152f
C74 B.t5 VSUBS 0.361054f
C75 B.t4 VSUBS 0.387145f
C76 B.t3 VSUBS 1.30555f
C77 B.n46 VSUBS 0.558492f
C78 B.n47 VSUBS 0.353407f
C79 B.n48 VSUBS 0.018889f
C80 B.n49 VSUBS 0.008152f
C81 B.n50 VSUBS 0.008152f
C82 B.n51 VSUBS 0.008152f
C83 B.n52 VSUBS 0.008152f
C84 B.t2 VSUBS 0.361058f
C85 B.t1 VSUBS 0.387148f
C86 B.t0 VSUBS 1.30555f
C87 B.n53 VSUBS 0.558488f
C88 B.n54 VSUBS 0.353403f
C89 B.n55 VSUBS 0.008152f
C90 B.n56 VSUBS 0.008152f
C91 B.n57 VSUBS 0.008152f
C92 B.n58 VSUBS 0.008152f
C93 B.n59 VSUBS 0.008152f
C94 B.n60 VSUBS 0.008152f
C95 B.n61 VSUBS 0.008152f
C96 B.n62 VSUBS 0.008152f
C97 B.n63 VSUBS 0.008152f
C98 B.n64 VSUBS 0.008152f
C99 B.n65 VSUBS 0.008152f
C100 B.n66 VSUBS 0.008152f
C101 B.n67 VSUBS 0.008152f
C102 B.n68 VSUBS 0.008152f
C103 B.n69 VSUBS 0.008152f
C104 B.n70 VSUBS 0.008152f
C105 B.n71 VSUBS 0.008152f
C106 B.n72 VSUBS 0.008152f
C107 B.n73 VSUBS 0.008152f
C108 B.n74 VSUBS 0.008152f
C109 B.n75 VSUBS 0.008152f
C110 B.n76 VSUBS 0.008152f
C111 B.n77 VSUBS 0.008152f
C112 B.n78 VSUBS 0.008152f
C113 B.n79 VSUBS 0.008152f
C114 B.n80 VSUBS 0.008152f
C115 B.n81 VSUBS 0.01753f
C116 B.n82 VSUBS 0.008152f
C117 B.n83 VSUBS 0.008152f
C118 B.n84 VSUBS 0.008152f
C119 B.n85 VSUBS 0.008152f
C120 B.n86 VSUBS 0.008152f
C121 B.n87 VSUBS 0.008152f
C122 B.n88 VSUBS 0.008152f
C123 B.n89 VSUBS 0.008152f
C124 B.n90 VSUBS 0.008152f
C125 B.n91 VSUBS 0.008152f
C126 B.n92 VSUBS 0.008152f
C127 B.n93 VSUBS 0.008152f
C128 B.n94 VSUBS 0.008152f
C129 B.n95 VSUBS 0.008152f
C130 B.n96 VSUBS 0.008152f
C131 B.n97 VSUBS 0.008152f
C132 B.n98 VSUBS 0.008152f
C133 B.n99 VSUBS 0.008152f
C134 B.n100 VSUBS 0.008152f
C135 B.n101 VSUBS 0.008152f
C136 B.n102 VSUBS 0.008152f
C137 B.n103 VSUBS 0.008152f
C138 B.n104 VSUBS 0.008152f
C139 B.n105 VSUBS 0.008152f
C140 B.n106 VSUBS 0.008152f
C141 B.n107 VSUBS 0.008152f
C142 B.n108 VSUBS 0.008152f
C143 B.n109 VSUBS 0.008152f
C144 B.n110 VSUBS 0.008152f
C145 B.n111 VSUBS 0.008152f
C146 B.n112 VSUBS 0.008152f
C147 B.n113 VSUBS 0.018563f
C148 B.n114 VSUBS 0.008152f
C149 B.n115 VSUBS 0.008152f
C150 B.n116 VSUBS 0.008152f
C151 B.n117 VSUBS 0.008152f
C152 B.n118 VSUBS 0.008152f
C153 B.n119 VSUBS 0.008152f
C154 B.n120 VSUBS 0.008152f
C155 B.n121 VSUBS 0.008152f
C156 B.n122 VSUBS 0.008152f
C157 B.n123 VSUBS 0.008152f
C158 B.n124 VSUBS 0.008152f
C159 B.n125 VSUBS 0.008152f
C160 B.n126 VSUBS 0.008152f
C161 B.n127 VSUBS 0.008152f
C162 B.n128 VSUBS 0.008152f
C163 B.n129 VSUBS 0.008152f
C164 B.n130 VSUBS 0.008152f
C165 B.n131 VSUBS 0.008152f
C166 B.n132 VSUBS 0.008152f
C167 B.n133 VSUBS 0.008152f
C168 B.n134 VSUBS 0.008152f
C169 B.n135 VSUBS 0.008152f
C170 B.n136 VSUBS 0.008152f
C171 B.n137 VSUBS 0.008152f
C172 B.n138 VSUBS 0.008152f
C173 B.n139 VSUBS 0.008152f
C174 B.n140 VSUBS 0.008152f
C175 B.t7 VSUBS 0.361058f
C176 B.t8 VSUBS 0.387148f
C177 B.t6 VSUBS 1.30555f
C178 B.n141 VSUBS 0.558488f
C179 B.n142 VSUBS 0.353403f
C180 B.n143 VSUBS 0.008152f
C181 B.n144 VSUBS 0.008152f
C182 B.n145 VSUBS 0.008152f
C183 B.n146 VSUBS 0.008152f
C184 B.t10 VSUBS 0.361054f
C185 B.t11 VSUBS 0.387145f
C186 B.t9 VSUBS 1.30555f
C187 B.n147 VSUBS 0.558492f
C188 B.n148 VSUBS 0.353407f
C189 B.n149 VSUBS 0.018889f
C190 B.n150 VSUBS 0.008152f
C191 B.n151 VSUBS 0.008152f
C192 B.n152 VSUBS 0.008152f
C193 B.n153 VSUBS 0.008152f
C194 B.n154 VSUBS 0.008152f
C195 B.n155 VSUBS 0.008152f
C196 B.n156 VSUBS 0.008152f
C197 B.n157 VSUBS 0.008152f
C198 B.n158 VSUBS 0.008152f
C199 B.n159 VSUBS 0.008152f
C200 B.n160 VSUBS 0.008152f
C201 B.n161 VSUBS 0.008152f
C202 B.n162 VSUBS 0.008152f
C203 B.n163 VSUBS 0.008152f
C204 B.n164 VSUBS 0.008152f
C205 B.n165 VSUBS 0.008152f
C206 B.n166 VSUBS 0.008152f
C207 B.n167 VSUBS 0.008152f
C208 B.n168 VSUBS 0.008152f
C209 B.n169 VSUBS 0.008152f
C210 B.n170 VSUBS 0.008152f
C211 B.n171 VSUBS 0.008152f
C212 B.n172 VSUBS 0.008152f
C213 B.n173 VSUBS 0.008152f
C214 B.n174 VSUBS 0.008152f
C215 B.n175 VSUBS 0.008152f
C216 B.n176 VSUBS 0.018563f
C217 B.n177 VSUBS 0.008152f
C218 B.n178 VSUBS 0.008152f
C219 B.n179 VSUBS 0.008152f
C220 B.n180 VSUBS 0.008152f
C221 B.n181 VSUBS 0.008152f
C222 B.n182 VSUBS 0.008152f
C223 B.n183 VSUBS 0.008152f
C224 B.n184 VSUBS 0.008152f
C225 B.n185 VSUBS 0.008152f
C226 B.n186 VSUBS 0.008152f
C227 B.n187 VSUBS 0.008152f
C228 B.n188 VSUBS 0.008152f
C229 B.n189 VSUBS 0.008152f
C230 B.n190 VSUBS 0.008152f
C231 B.n191 VSUBS 0.008152f
C232 B.n192 VSUBS 0.008152f
C233 B.n193 VSUBS 0.008152f
C234 B.n194 VSUBS 0.008152f
C235 B.n195 VSUBS 0.008152f
C236 B.n196 VSUBS 0.008152f
C237 B.n197 VSUBS 0.008152f
C238 B.n198 VSUBS 0.008152f
C239 B.n199 VSUBS 0.008152f
C240 B.n200 VSUBS 0.008152f
C241 B.n201 VSUBS 0.008152f
C242 B.n202 VSUBS 0.008152f
C243 B.n203 VSUBS 0.008152f
C244 B.n204 VSUBS 0.008152f
C245 B.n205 VSUBS 0.008152f
C246 B.n206 VSUBS 0.008152f
C247 B.n207 VSUBS 0.008152f
C248 B.n208 VSUBS 0.008152f
C249 B.n209 VSUBS 0.008152f
C250 B.n210 VSUBS 0.008152f
C251 B.n211 VSUBS 0.008152f
C252 B.n212 VSUBS 0.008152f
C253 B.n213 VSUBS 0.008152f
C254 B.n214 VSUBS 0.008152f
C255 B.n215 VSUBS 0.008152f
C256 B.n216 VSUBS 0.008152f
C257 B.n217 VSUBS 0.008152f
C258 B.n218 VSUBS 0.008152f
C259 B.n219 VSUBS 0.008152f
C260 B.n220 VSUBS 0.008152f
C261 B.n221 VSUBS 0.008152f
C262 B.n222 VSUBS 0.008152f
C263 B.n223 VSUBS 0.008152f
C264 B.n224 VSUBS 0.008152f
C265 B.n225 VSUBS 0.008152f
C266 B.n226 VSUBS 0.008152f
C267 B.n227 VSUBS 0.008152f
C268 B.n228 VSUBS 0.008152f
C269 B.n229 VSUBS 0.008152f
C270 B.n230 VSUBS 0.008152f
C271 B.n231 VSUBS 0.008152f
C272 B.n232 VSUBS 0.008152f
C273 B.n233 VSUBS 0.008152f
C274 B.n234 VSUBS 0.008152f
C275 B.n235 VSUBS 0.017883f
C276 B.n236 VSUBS 0.017883f
C277 B.n237 VSUBS 0.018563f
C278 B.n238 VSUBS 0.008152f
C279 B.n239 VSUBS 0.008152f
C280 B.n240 VSUBS 0.008152f
C281 B.n241 VSUBS 0.008152f
C282 B.n242 VSUBS 0.008152f
C283 B.n243 VSUBS 0.008152f
C284 B.n244 VSUBS 0.008152f
C285 B.n245 VSUBS 0.008152f
C286 B.n246 VSUBS 0.008152f
C287 B.n247 VSUBS 0.008152f
C288 B.n248 VSUBS 0.008152f
C289 B.n249 VSUBS 0.008152f
C290 B.n250 VSUBS 0.008152f
C291 B.n251 VSUBS 0.008152f
C292 B.n252 VSUBS 0.008152f
C293 B.n253 VSUBS 0.008152f
C294 B.n254 VSUBS 0.008152f
C295 B.n255 VSUBS 0.008152f
C296 B.n256 VSUBS 0.008152f
C297 B.n257 VSUBS 0.008152f
C298 B.n258 VSUBS 0.008152f
C299 B.n259 VSUBS 0.008152f
C300 B.n260 VSUBS 0.008152f
C301 B.n261 VSUBS 0.008152f
C302 B.n262 VSUBS 0.008152f
C303 B.n263 VSUBS 0.008152f
C304 B.n264 VSUBS 0.008152f
C305 B.n265 VSUBS 0.008152f
C306 B.n266 VSUBS 0.008152f
C307 B.n267 VSUBS 0.008152f
C308 B.n268 VSUBS 0.008152f
C309 B.n269 VSUBS 0.008152f
C310 B.n270 VSUBS 0.008152f
C311 B.n271 VSUBS 0.008152f
C312 B.n272 VSUBS 0.008152f
C313 B.n273 VSUBS 0.008152f
C314 B.n274 VSUBS 0.008152f
C315 B.n275 VSUBS 0.008152f
C316 B.n276 VSUBS 0.008152f
C317 B.n277 VSUBS 0.008152f
C318 B.n278 VSUBS 0.008152f
C319 B.n279 VSUBS 0.008152f
C320 B.n280 VSUBS 0.008152f
C321 B.n281 VSUBS 0.008152f
C322 B.n282 VSUBS 0.008152f
C323 B.n283 VSUBS 0.008152f
C324 B.n284 VSUBS 0.008152f
C325 B.n285 VSUBS 0.008152f
C326 B.n286 VSUBS 0.008152f
C327 B.n287 VSUBS 0.008152f
C328 B.n288 VSUBS 0.008152f
C329 B.n289 VSUBS 0.008152f
C330 B.n290 VSUBS 0.008152f
C331 B.n291 VSUBS 0.008152f
C332 B.n292 VSUBS 0.008152f
C333 B.n293 VSUBS 0.008152f
C334 B.n294 VSUBS 0.008152f
C335 B.n295 VSUBS 0.008152f
C336 B.n296 VSUBS 0.008152f
C337 B.n297 VSUBS 0.008152f
C338 B.n298 VSUBS 0.008152f
C339 B.n299 VSUBS 0.008152f
C340 B.n300 VSUBS 0.008152f
C341 B.n301 VSUBS 0.008152f
C342 B.n302 VSUBS 0.008152f
C343 B.n303 VSUBS 0.008152f
C344 B.n304 VSUBS 0.008152f
C345 B.n305 VSUBS 0.008152f
C346 B.n306 VSUBS 0.008152f
C347 B.n307 VSUBS 0.008152f
C348 B.n308 VSUBS 0.008152f
C349 B.n309 VSUBS 0.008152f
C350 B.n310 VSUBS 0.008152f
C351 B.n311 VSUBS 0.008152f
C352 B.n312 VSUBS 0.008152f
C353 B.n313 VSUBS 0.008152f
C354 B.n314 VSUBS 0.008152f
C355 B.n315 VSUBS 0.008152f
C356 B.n316 VSUBS 0.007673f
C357 B.n317 VSUBS 0.008152f
C358 B.n318 VSUBS 0.008152f
C359 B.n319 VSUBS 0.004556f
C360 B.n320 VSUBS 0.008152f
C361 B.n321 VSUBS 0.008152f
C362 B.n322 VSUBS 0.008152f
C363 B.n323 VSUBS 0.008152f
C364 B.n324 VSUBS 0.008152f
C365 B.n325 VSUBS 0.008152f
C366 B.n326 VSUBS 0.008152f
C367 B.n327 VSUBS 0.008152f
C368 B.n328 VSUBS 0.008152f
C369 B.n329 VSUBS 0.008152f
C370 B.n330 VSUBS 0.008152f
C371 B.n331 VSUBS 0.008152f
C372 B.n332 VSUBS 0.004556f
C373 B.n333 VSUBS 0.018889f
C374 B.n334 VSUBS 0.007673f
C375 B.n335 VSUBS 0.008152f
C376 B.n336 VSUBS 0.008152f
C377 B.n337 VSUBS 0.008152f
C378 B.n338 VSUBS 0.008152f
C379 B.n339 VSUBS 0.008152f
C380 B.n340 VSUBS 0.008152f
C381 B.n341 VSUBS 0.008152f
C382 B.n342 VSUBS 0.008152f
C383 B.n343 VSUBS 0.008152f
C384 B.n344 VSUBS 0.008152f
C385 B.n345 VSUBS 0.008152f
C386 B.n346 VSUBS 0.008152f
C387 B.n347 VSUBS 0.008152f
C388 B.n348 VSUBS 0.008152f
C389 B.n349 VSUBS 0.008152f
C390 B.n350 VSUBS 0.008152f
C391 B.n351 VSUBS 0.008152f
C392 B.n352 VSUBS 0.008152f
C393 B.n353 VSUBS 0.008152f
C394 B.n354 VSUBS 0.008152f
C395 B.n355 VSUBS 0.008152f
C396 B.n356 VSUBS 0.008152f
C397 B.n357 VSUBS 0.008152f
C398 B.n358 VSUBS 0.008152f
C399 B.n359 VSUBS 0.008152f
C400 B.n360 VSUBS 0.008152f
C401 B.n361 VSUBS 0.008152f
C402 B.n362 VSUBS 0.008152f
C403 B.n363 VSUBS 0.008152f
C404 B.n364 VSUBS 0.008152f
C405 B.n365 VSUBS 0.008152f
C406 B.n366 VSUBS 0.008152f
C407 B.n367 VSUBS 0.008152f
C408 B.n368 VSUBS 0.008152f
C409 B.n369 VSUBS 0.008152f
C410 B.n370 VSUBS 0.008152f
C411 B.n371 VSUBS 0.008152f
C412 B.n372 VSUBS 0.008152f
C413 B.n373 VSUBS 0.008152f
C414 B.n374 VSUBS 0.008152f
C415 B.n375 VSUBS 0.008152f
C416 B.n376 VSUBS 0.008152f
C417 B.n377 VSUBS 0.008152f
C418 B.n378 VSUBS 0.008152f
C419 B.n379 VSUBS 0.008152f
C420 B.n380 VSUBS 0.008152f
C421 B.n381 VSUBS 0.008152f
C422 B.n382 VSUBS 0.008152f
C423 B.n383 VSUBS 0.008152f
C424 B.n384 VSUBS 0.008152f
C425 B.n385 VSUBS 0.008152f
C426 B.n386 VSUBS 0.008152f
C427 B.n387 VSUBS 0.008152f
C428 B.n388 VSUBS 0.008152f
C429 B.n389 VSUBS 0.008152f
C430 B.n390 VSUBS 0.008152f
C431 B.n391 VSUBS 0.008152f
C432 B.n392 VSUBS 0.008152f
C433 B.n393 VSUBS 0.008152f
C434 B.n394 VSUBS 0.008152f
C435 B.n395 VSUBS 0.008152f
C436 B.n396 VSUBS 0.008152f
C437 B.n397 VSUBS 0.008152f
C438 B.n398 VSUBS 0.008152f
C439 B.n399 VSUBS 0.008152f
C440 B.n400 VSUBS 0.008152f
C441 B.n401 VSUBS 0.008152f
C442 B.n402 VSUBS 0.008152f
C443 B.n403 VSUBS 0.008152f
C444 B.n404 VSUBS 0.008152f
C445 B.n405 VSUBS 0.008152f
C446 B.n406 VSUBS 0.008152f
C447 B.n407 VSUBS 0.008152f
C448 B.n408 VSUBS 0.008152f
C449 B.n409 VSUBS 0.008152f
C450 B.n410 VSUBS 0.008152f
C451 B.n411 VSUBS 0.008152f
C452 B.n412 VSUBS 0.008152f
C453 B.n413 VSUBS 0.008152f
C454 B.n414 VSUBS 0.018563f
C455 B.n415 VSUBS 0.017883f
C456 B.n416 VSUBS 0.017883f
C457 B.n417 VSUBS 0.008152f
C458 B.n418 VSUBS 0.008152f
C459 B.n419 VSUBS 0.008152f
C460 B.n420 VSUBS 0.008152f
C461 B.n421 VSUBS 0.008152f
C462 B.n422 VSUBS 0.008152f
C463 B.n423 VSUBS 0.008152f
C464 B.n424 VSUBS 0.008152f
C465 B.n425 VSUBS 0.008152f
C466 B.n426 VSUBS 0.008152f
C467 B.n427 VSUBS 0.008152f
C468 B.n428 VSUBS 0.008152f
C469 B.n429 VSUBS 0.008152f
C470 B.n430 VSUBS 0.008152f
C471 B.n431 VSUBS 0.008152f
C472 B.n432 VSUBS 0.008152f
C473 B.n433 VSUBS 0.008152f
C474 B.n434 VSUBS 0.008152f
C475 B.n435 VSUBS 0.008152f
C476 B.n436 VSUBS 0.008152f
C477 B.n437 VSUBS 0.008152f
C478 B.n438 VSUBS 0.008152f
C479 B.n439 VSUBS 0.008152f
C480 B.n440 VSUBS 0.008152f
C481 B.n441 VSUBS 0.008152f
C482 B.n442 VSUBS 0.008152f
C483 B.n443 VSUBS 0.008152f
C484 B.n444 VSUBS 0.008152f
C485 B.n445 VSUBS 0.008152f
C486 B.n446 VSUBS 0.008152f
C487 B.n447 VSUBS 0.008152f
C488 B.n448 VSUBS 0.008152f
C489 B.n449 VSUBS 0.008152f
C490 B.n450 VSUBS 0.008152f
C491 B.n451 VSUBS 0.008152f
C492 B.n452 VSUBS 0.008152f
C493 B.n453 VSUBS 0.008152f
C494 B.n454 VSUBS 0.008152f
C495 B.n455 VSUBS 0.008152f
C496 B.n456 VSUBS 0.008152f
C497 B.n457 VSUBS 0.008152f
C498 B.n458 VSUBS 0.008152f
C499 B.n459 VSUBS 0.008152f
C500 B.n460 VSUBS 0.008152f
C501 B.n461 VSUBS 0.008152f
C502 B.n462 VSUBS 0.008152f
C503 B.n463 VSUBS 0.008152f
C504 B.n464 VSUBS 0.008152f
C505 B.n465 VSUBS 0.008152f
C506 B.n466 VSUBS 0.008152f
C507 B.n467 VSUBS 0.008152f
C508 B.n468 VSUBS 0.008152f
C509 B.n469 VSUBS 0.008152f
C510 B.n470 VSUBS 0.008152f
C511 B.n471 VSUBS 0.008152f
C512 B.n472 VSUBS 0.008152f
C513 B.n473 VSUBS 0.008152f
C514 B.n474 VSUBS 0.008152f
C515 B.n475 VSUBS 0.008152f
C516 B.n476 VSUBS 0.008152f
C517 B.n477 VSUBS 0.008152f
C518 B.n478 VSUBS 0.008152f
C519 B.n479 VSUBS 0.008152f
C520 B.n480 VSUBS 0.008152f
C521 B.n481 VSUBS 0.008152f
C522 B.n482 VSUBS 0.008152f
C523 B.n483 VSUBS 0.008152f
C524 B.n484 VSUBS 0.008152f
C525 B.n485 VSUBS 0.008152f
C526 B.n486 VSUBS 0.008152f
C527 B.n487 VSUBS 0.008152f
C528 B.n488 VSUBS 0.008152f
C529 B.n489 VSUBS 0.008152f
C530 B.n490 VSUBS 0.008152f
C531 B.n491 VSUBS 0.008152f
C532 B.n492 VSUBS 0.008152f
C533 B.n493 VSUBS 0.008152f
C534 B.n494 VSUBS 0.008152f
C535 B.n495 VSUBS 0.008152f
C536 B.n496 VSUBS 0.008152f
C537 B.n497 VSUBS 0.008152f
C538 B.n498 VSUBS 0.008152f
C539 B.n499 VSUBS 0.008152f
C540 B.n500 VSUBS 0.008152f
C541 B.n501 VSUBS 0.008152f
C542 B.n502 VSUBS 0.008152f
C543 B.n503 VSUBS 0.008152f
C544 B.n504 VSUBS 0.008152f
C545 B.n505 VSUBS 0.008152f
C546 B.n506 VSUBS 0.008152f
C547 B.n507 VSUBS 0.008152f
C548 B.n508 VSUBS 0.018916f
C549 B.n509 VSUBS 0.017883f
C550 B.n510 VSUBS 0.018563f
C551 B.n511 VSUBS 0.008152f
C552 B.n512 VSUBS 0.008152f
C553 B.n513 VSUBS 0.008152f
C554 B.n514 VSUBS 0.008152f
C555 B.n515 VSUBS 0.008152f
C556 B.n516 VSUBS 0.008152f
C557 B.n517 VSUBS 0.008152f
C558 B.n518 VSUBS 0.008152f
C559 B.n519 VSUBS 0.008152f
C560 B.n520 VSUBS 0.008152f
C561 B.n521 VSUBS 0.008152f
C562 B.n522 VSUBS 0.008152f
C563 B.n523 VSUBS 0.008152f
C564 B.n524 VSUBS 0.008152f
C565 B.n525 VSUBS 0.008152f
C566 B.n526 VSUBS 0.008152f
C567 B.n527 VSUBS 0.008152f
C568 B.n528 VSUBS 0.008152f
C569 B.n529 VSUBS 0.008152f
C570 B.n530 VSUBS 0.008152f
C571 B.n531 VSUBS 0.008152f
C572 B.n532 VSUBS 0.008152f
C573 B.n533 VSUBS 0.008152f
C574 B.n534 VSUBS 0.008152f
C575 B.n535 VSUBS 0.008152f
C576 B.n536 VSUBS 0.008152f
C577 B.n537 VSUBS 0.008152f
C578 B.n538 VSUBS 0.008152f
C579 B.n539 VSUBS 0.008152f
C580 B.n540 VSUBS 0.008152f
C581 B.n541 VSUBS 0.008152f
C582 B.n542 VSUBS 0.008152f
C583 B.n543 VSUBS 0.008152f
C584 B.n544 VSUBS 0.008152f
C585 B.n545 VSUBS 0.008152f
C586 B.n546 VSUBS 0.008152f
C587 B.n547 VSUBS 0.008152f
C588 B.n548 VSUBS 0.008152f
C589 B.n549 VSUBS 0.008152f
C590 B.n550 VSUBS 0.008152f
C591 B.n551 VSUBS 0.008152f
C592 B.n552 VSUBS 0.008152f
C593 B.n553 VSUBS 0.008152f
C594 B.n554 VSUBS 0.008152f
C595 B.n555 VSUBS 0.008152f
C596 B.n556 VSUBS 0.008152f
C597 B.n557 VSUBS 0.008152f
C598 B.n558 VSUBS 0.008152f
C599 B.n559 VSUBS 0.008152f
C600 B.n560 VSUBS 0.008152f
C601 B.n561 VSUBS 0.008152f
C602 B.n562 VSUBS 0.008152f
C603 B.n563 VSUBS 0.008152f
C604 B.n564 VSUBS 0.008152f
C605 B.n565 VSUBS 0.008152f
C606 B.n566 VSUBS 0.008152f
C607 B.n567 VSUBS 0.008152f
C608 B.n568 VSUBS 0.008152f
C609 B.n569 VSUBS 0.008152f
C610 B.n570 VSUBS 0.008152f
C611 B.n571 VSUBS 0.008152f
C612 B.n572 VSUBS 0.008152f
C613 B.n573 VSUBS 0.008152f
C614 B.n574 VSUBS 0.008152f
C615 B.n575 VSUBS 0.008152f
C616 B.n576 VSUBS 0.008152f
C617 B.n577 VSUBS 0.008152f
C618 B.n578 VSUBS 0.008152f
C619 B.n579 VSUBS 0.008152f
C620 B.n580 VSUBS 0.008152f
C621 B.n581 VSUBS 0.008152f
C622 B.n582 VSUBS 0.008152f
C623 B.n583 VSUBS 0.008152f
C624 B.n584 VSUBS 0.008152f
C625 B.n585 VSUBS 0.008152f
C626 B.n586 VSUBS 0.008152f
C627 B.n587 VSUBS 0.008152f
C628 B.n588 VSUBS 0.008152f
C629 B.n589 VSUBS 0.008152f
C630 B.n590 VSUBS 0.007673f
C631 B.n591 VSUBS 0.018889f
C632 B.n592 VSUBS 0.004556f
C633 B.n593 VSUBS 0.008152f
C634 B.n594 VSUBS 0.008152f
C635 B.n595 VSUBS 0.008152f
C636 B.n596 VSUBS 0.008152f
C637 B.n597 VSUBS 0.008152f
C638 B.n598 VSUBS 0.008152f
C639 B.n599 VSUBS 0.008152f
C640 B.n600 VSUBS 0.008152f
C641 B.n601 VSUBS 0.008152f
C642 B.n602 VSUBS 0.008152f
C643 B.n603 VSUBS 0.008152f
C644 B.n604 VSUBS 0.008152f
C645 B.n605 VSUBS 0.004556f
C646 B.n606 VSUBS 0.008152f
C647 B.n607 VSUBS 0.008152f
C648 B.n608 VSUBS 0.008152f
C649 B.n609 VSUBS 0.008152f
C650 B.n610 VSUBS 0.008152f
C651 B.n611 VSUBS 0.008152f
C652 B.n612 VSUBS 0.008152f
C653 B.n613 VSUBS 0.008152f
C654 B.n614 VSUBS 0.008152f
C655 B.n615 VSUBS 0.008152f
C656 B.n616 VSUBS 0.008152f
C657 B.n617 VSUBS 0.008152f
C658 B.n618 VSUBS 0.008152f
C659 B.n619 VSUBS 0.008152f
C660 B.n620 VSUBS 0.008152f
C661 B.n621 VSUBS 0.008152f
C662 B.n622 VSUBS 0.008152f
C663 B.n623 VSUBS 0.008152f
C664 B.n624 VSUBS 0.008152f
C665 B.n625 VSUBS 0.008152f
C666 B.n626 VSUBS 0.008152f
C667 B.n627 VSUBS 0.008152f
C668 B.n628 VSUBS 0.008152f
C669 B.n629 VSUBS 0.008152f
C670 B.n630 VSUBS 0.008152f
C671 B.n631 VSUBS 0.008152f
C672 B.n632 VSUBS 0.008152f
C673 B.n633 VSUBS 0.008152f
C674 B.n634 VSUBS 0.008152f
C675 B.n635 VSUBS 0.008152f
C676 B.n636 VSUBS 0.008152f
C677 B.n637 VSUBS 0.008152f
C678 B.n638 VSUBS 0.008152f
C679 B.n639 VSUBS 0.008152f
C680 B.n640 VSUBS 0.008152f
C681 B.n641 VSUBS 0.008152f
C682 B.n642 VSUBS 0.008152f
C683 B.n643 VSUBS 0.008152f
C684 B.n644 VSUBS 0.008152f
C685 B.n645 VSUBS 0.008152f
C686 B.n646 VSUBS 0.008152f
C687 B.n647 VSUBS 0.008152f
C688 B.n648 VSUBS 0.008152f
C689 B.n649 VSUBS 0.008152f
C690 B.n650 VSUBS 0.008152f
C691 B.n651 VSUBS 0.008152f
C692 B.n652 VSUBS 0.008152f
C693 B.n653 VSUBS 0.008152f
C694 B.n654 VSUBS 0.008152f
C695 B.n655 VSUBS 0.008152f
C696 B.n656 VSUBS 0.008152f
C697 B.n657 VSUBS 0.008152f
C698 B.n658 VSUBS 0.008152f
C699 B.n659 VSUBS 0.008152f
C700 B.n660 VSUBS 0.008152f
C701 B.n661 VSUBS 0.008152f
C702 B.n662 VSUBS 0.008152f
C703 B.n663 VSUBS 0.008152f
C704 B.n664 VSUBS 0.008152f
C705 B.n665 VSUBS 0.008152f
C706 B.n666 VSUBS 0.008152f
C707 B.n667 VSUBS 0.008152f
C708 B.n668 VSUBS 0.008152f
C709 B.n669 VSUBS 0.008152f
C710 B.n670 VSUBS 0.008152f
C711 B.n671 VSUBS 0.008152f
C712 B.n672 VSUBS 0.008152f
C713 B.n673 VSUBS 0.008152f
C714 B.n674 VSUBS 0.008152f
C715 B.n675 VSUBS 0.008152f
C716 B.n676 VSUBS 0.008152f
C717 B.n677 VSUBS 0.008152f
C718 B.n678 VSUBS 0.008152f
C719 B.n679 VSUBS 0.008152f
C720 B.n680 VSUBS 0.008152f
C721 B.n681 VSUBS 0.008152f
C722 B.n682 VSUBS 0.008152f
C723 B.n683 VSUBS 0.008152f
C724 B.n684 VSUBS 0.008152f
C725 B.n685 VSUBS 0.008152f
C726 B.n686 VSUBS 0.018563f
C727 B.n687 VSUBS 0.018563f
C728 B.n688 VSUBS 0.017883f
C729 B.n689 VSUBS 0.008152f
C730 B.n690 VSUBS 0.008152f
C731 B.n691 VSUBS 0.008152f
C732 B.n692 VSUBS 0.008152f
C733 B.n693 VSUBS 0.008152f
C734 B.n694 VSUBS 0.008152f
C735 B.n695 VSUBS 0.008152f
C736 B.n696 VSUBS 0.008152f
C737 B.n697 VSUBS 0.008152f
C738 B.n698 VSUBS 0.008152f
C739 B.n699 VSUBS 0.008152f
C740 B.n700 VSUBS 0.008152f
C741 B.n701 VSUBS 0.008152f
C742 B.n702 VSUBS 0.008152f
C743 B.n703 VSUBS 0.008152f
C744 B.n704 VSUBS 0.008152f
C745 B.n705 VSUBS 0.008152f
C746 B.n706 VSUBS 0.008152f
C747 B.n707 VSUBS 0.008152f
C748 B.n708 VSUBS 0.008152f
C749 B.n709 VSUBS 0.008152f
C750 B.n710 VSUBS 0.008152f
C751 B.n711 VSUBS 0.008152f
C752 B.n712 VSUBS 0.008152f
C753 B.n713 VSUBS 0.008152f
C754 B.n714 VSUBS 0.008152f
C755 B.n715 VSUBS 0.008152f
C756 B.n716 VSUBS 0.008152f
C757 B.n717 VSUBS 0.008152f
C758 B.n718 VSUBS 0.008152f
C759 B.n719 VSUBS 0.008152f
C760 B.n720 VSUBS 0.008152f
C761 B.n721 VSUBS 0.008152f
C762 B.n722 VSUBS 0.008152f
C763 B.n723 VSUBS 0.008152f
C764 B.n724 VSUBS 0.008152f
C765 B.n725 VSUBS 0.008152f
C766 B.n726 VSUBS 0.008152f
C767 B.n727 VSUBS 0.008152f
C768 B.n728 VSUBS 0.008152f
C769 B.n729 VSUBS 0.008152f
C770 B.n730 VSUBS 0.008152f
C771 B.n731 VSUBS 0.008152f
C772 B.n732 VSUBS 0.008152f
C773 B.n733 VSUBS 0.008152f
C774 B.n734 VSUBS 0.008152f
C775 B.n735 VSUBS 0.01846f
C776 VDD2.n0 VSUBS 0.030674f
C777 VDD2.n1 VSUBS 0.027181f
C778 VDD2.n2 VSUBS 0.014606f
C779 VDD2.n3 VSUBS 0.034522f
C780 VDD2.n4 VSUBS 0.015465f
C781 VDD2.n5 VSUBS 0.027181f
C782 VDD2.n6 VSUBS 0.015035f
C783 VDD2.n7 VSUBS 0.034522f
C784 VDD2.n8 VSUBS 0.015465f
C785 VDD2.n9 VSUBS 0.027181f
C786 VDD2.n10 VSUBS 0.014606f
C787 VDD2.n11 VSUBS 0.034522f
C788 VDD2.n12 VSUBS 0.015465f
C789 VDD2.n13 VSUBS 0.027181f
C790 VDD2.n14 VSUBS 0.014606f
C791 VDD2.n15 VSUBS 0.034522f
C792 VDD2.n16 VSUBS 0.015465f
C793 VDD2.n17 VSUBS 0.027181f
C794 VDD2.n18 VSUBS 0.014606f
C795 VDD2.n19 VSUBS 0.034522f
C796 VDD2.n20 VSUBS 0.015465f
C797 VDD2.n21 VSUBS 0.027181f
C798 VDD2.n22 VSUBS 0.014606f
C799 VDD2.n23 VSUBS 0.034522f
C800 VDD2.n24 VSUBS 0.015465f
C801 VDD2.n25 VSUBS 0.027181f
C802 VDD2.n26 VSUBS 0.014606f
C803 VDD2.n27 VSUBS 0.025892f
C804 VDD2.n28 VSUBS 0.021962f
C805 VDD2.t4 VSUBS 0.073992f
C806 VDD2.n29 VSUBS 0.201862f
C807 VDD2.n30 VSUBS 1.89348f
C808 VDD2.n31 VSUBS 0.014606f
C809 VDD2.n32 VSUBS 0.015465f
C810 VDD2.n33 VSUBS 0.034522f
C811 VDD2.n34 VSUBS 0.034522f
C812 VDD2.n35 VSUBS 0.015465f
C813 VDD2.n36 VSUBS 0.014606f
C814 VDD2.n37 VSUBS 0.027181f
C815 VDD2.n38 VSUBS 0.027181f
C816 VDD2.n39 VSUBS 0.014606f
C817 VDD2.n40 VSUBS 0.015465f
C818 VDD2.n41 VSUBS 0.034522f
C819 VDD2.n42 VSUBS 0.034522f
C820 VDD2.n43 VSUBS 0.015465f
C821 VDD2.n44 VSUBS 0.014606f
C822 VDD2.n45 VSUBS 0.027181f
C823 VDD2.n46 VSUBS 0.027181f
C824 VDD2.n47 VSUBS 0.014606f
C825 VDD2.n48 VSUBS 0.015465f
C826 VDD2.n49 VSUBS 0.034522f
C827 VDD2.n50 VSUBS 0.034522f
C828 VDD2.n51 VSUBS 0.015465f
C829 VDD2.n52 VSUBS 0.014606f
C830 VDD2.n53 VSUBS 0.027181f
C831 VDD2.n54 VSUBS 0.027181f
C832 VDD2.n55 VSUBS 0.014606f
C833 VDD2.n56 VSUBS 0.015465f
C834 VDD2.n57 VSUBS 0.034522f
C835 VDD2.n58 VSUBS 0.034522f
C836 VDD2.n59 VSUBS 0.015465f
C837 VDD2.n60 VSUBS 0.014606f
C838 VDD2.n61 VSUBS 0.027181f
C839 VDD2.n62 VSUBS 0.027181f
C840 VDD2.n63 VSUBS 0.014606f
C841 VDD2.n64 VSUBS 0.015465f
C842 VDD2.n65 VSUBS 0.034522f
C843 VDD2.n66 VSUBS 0.034522f
C844 VDD2.n67 VSUBS 0.015465f
C845 VDD2.n68 VSUBS 0.014606f
C846 VDD2.n69 VSUBS 0.027181f
C847 VDD2.n70 VSUBS 0.027181f
C848 VDD2.n71 VSUBS 0.014606f
C849 VDD2.n72 VSUBS 0.014606f
C850 VDD2.n73 VSUBS 0.015465f
C851 VDD2.n74 VSUBS 0.034522f
C852 VDD2.n75 VSUBS 0.034522f
C853 VDD2.n76 VSUBS 0.034522f
C854 VDD2.n77 VSUBS 0.015035f
C855 VDD2.n78 VSUBS 0.014606f
C856 VDD2.n79 VSUBS 0.027181f
C857 VDD2.n80 VSUBS 0.027181f
C858 VDD2.n81 VSUBS 0.014606f
C859 VDD2.n82 VSUBS 0.015465f
C860 VDD2.n83 VSUBS 0.034522f
C861 VDD2.n84 VSUBS 0.086328f
C862 VDD2.n85 VSUBS 0.015465f
C863 VDD2.n86 VSUBS 0.014606f
C864 VDD2.n87 VSUBS 0.070253f
C865 VDD2.n88 VSUBS 0.066041f
C866 VDD2.t2 VSUBS 0.349677f
C867 VDD2.t1 VSUBS 0.349677f
C868 VDD2.n89 VSUBS 2.88828f
C869 VDD2.n90 VSUBS 3.01965f
C870 VDD2.n91 VSUBS 0.030674f
C871 VDD2.n92 VSUBS 0.027181f
C872 VDD2.n93 VSUBS 0.014606f
C873 VDD2.n94 VSUBS 0.034522f
C874 VDD2.n95 VSUBS 0.015465f
C875 VDD2.n96 VSUBS 0.027181f
C876 VDD2.n97 VSUBS 0.015035f
C877 VDD2.n98 VSUBS 0.034522f
C878 VDD2.n99 VSUBS 0.014606f
C879 VDD2.n100 VSUBS 0.015465f
C880 VDD2.n101 VSUBS 0.027181f
C881 VDD2.n102 VSUBS 0.014606f
C882 VDD2.n103 VSUBS 0.034522f
C883 VDD2.n104 VSUBS 0.015465f
C884 VDD2.n105 VSUBS 0.027181f
C885 VDD2.n106 VSUBS 0.014606f
C886 VDD2.n107 VSUBS 0.034522f
C887 VDD2.n108 VSUBS 0.015465f
C888 VDD2.n109 VSUBS 0.027181f
C889 VDD2.n110 VSUBS 0.014606f
C890 VDD2.n111 VSUBS 0.034522f
C891 VDD2.n112 VSUBS 0.015465f
C892 VDD2.n113 VSUBS 0.027181f
C893 VDD2.n114 VSUBS 0.014606f
C894 VDD2.n115 VSUBS 0.034522f
C895 VDD2.n116 VSUBS 0.015465f
C896 VDD2.n117 VSUBS 0.027181f
C897 VDD2.n118 VSUBS 0.014606f
C898 VDD2.n119 VSUBS 0.025892f
C899 VDD2.n120 VSUBS 0.021962f
C900 VDD2.t5 VSUBS 0.073992f
C901 VDD2.n121 VSUBS 0.201862f
C902 VDD2.n122 VSUBS 1.89348f
C903 VDD2.n123 VSUBS 0.014606f
C904 VDD2.n124 VSUBS 0.015465f
C905 VDD2.n125 VSUBS 0.034522f
C906 VDD2.n126 VSUBS 0.034522f
C907 VDD2.n127 VSUBS 0.015465f
C908 VDD2.n128 VSUBS 0.014606f
C909 VDD2.n129 VSUBS 0.027181f
C910 VDD2.n130 VSUBS 0.027181f
C911 VDD2.n131 VSUBS 0.014606f
C912 VDD2.n132 VSUBS 0.015465f
C913 VDD2.n133 VSUBS 0.034522f
C914 VDD2.n134 VSUBS 0.034522f
C915 VDD2.n135 VSUBS 0.015465f
C916 VDD2.n136 VSUBS 0.014606f
C917 VDD2.n137 VSUBS 0.027181f
C918 VDD2.n138 VSUBS 0.027181f
C919 VDD2.n139 VSUBS 0.014606f
C920 VDD2.n140 VSUBS 0.015465f
C921 VDD2.n141 VSUBS 0.034522f
C922 VDD2.n142 VSUBS 0.034522f
C923 VDD2.n143 VSUBS 0.015465f
C924 VDD2.n144 VSUBS 0.014606f
C925 VDD2.n145 VSUBS 0.027181f
C926 VDD2.n146 VSUBS 0.027181f
C927 VDD2.n147 VSUBS 0.014606f
C928 VDD2.n148 VSUBS 0.015465f
C929 VDD2.n149 VSUBS 0.034522f
C930 VDD2.n150 VSUBS 0.034522f
C931 VDD2.n151 VSUBS 0.015465f
C932 VDD2.n152 VSUBS 0.014606f
C933 VDD2.n153 VSUBS 0.027181f
C934 VDD2.n154 VSUBS 0.027181f
C935 VDD2.n155 VSUBS 0.014606f
C936 VDD2.n156 VSUBS 0.015465f
C937 VDD2.n157 VSUBS 0.034522f
C938 VDD2.n158 VSUBS 0.034522f
C939 VDD2.n159 VSUBS 0.015465f
C940 VDD2.n160 VSUBS 0.014606f
C941 VDD2.n161 VSUBS 0.027181f
C942 VDD2.n162 VSUBS 0.027181f
C943 VDD2.n163 VSUBS 0.014606f
C944 VDD2.n164 VSUBS 0.015465f
C945 VDD2.n165 VSUBS 0.034522f
C946 VDD2.n166 VSUBS 0.034522f
C947 VDD2.n167 VSUBS 0.034522f
C948 VDD2.n168 VSUBS 0.015035f
C949 VDD2.n169 VSUBS 0.014606f
C950 VDD2.n170 VSUBS 0.027181f
C951 VDD2.n171 VSUBS 0.027181f
C952 VDD2.n172 VSUBS 0.014606f
C953 VDD2.n173 VSUBS 0.015465f
C954 VDD2.n174 VSUBS 0.034522f
C955 VDD2.n175 VSUBS 0.086328f
C956 VDD2.n176 VSUBS 0.015465f
C957 VDD2.n177 VSUBS 0.014606f
C958 VDD2.n178 VSUBS 0.070253f
C959 VDD2.n179 VSUBS 0.062469f
C960 VDD2.n180 VSUBS 2.85085f
C961 VDD2.t0 VSUBS 0.349677f
C962 VDD2.t3 VSUBS 0.349677f
C963 VDD2.n181 VSUBS 2.88825f
C964 VN.n0 VSUBS 0.036855f
C965 VN.t4 VSUBS 2.63528f
C966 VN.n1 VSUBS 0.050416f
C967 VN.t1 VSUBS 2.76373f
C968 VN.n2 VSUBS 1.02195f
C969 VN.t3 VSUBS 2.63528f
C970 VN.n3 VSUBS 1.00299f
C971 VN.n4 VSUBS 0.051991f
C972 VN.n5 VSUBS 0.235347f
C973 VN.n6 VSUBS 0.036855f
C974 VN.n7 VSUBS 0.036855f
C975 VN.n8 VSUBS 0.057656f
C976 VN.n9 VSUBS 0.047219f
C977 VN.n10 VSUBS 1.01123f
C978 VN.n11 VSUBS 0.036323f
C979 VN.n12 VSUBS 0.036855f
C980 VN.t0 VSUBS 2.63528f
C981 VN.n13 VSUBS 0.050416f
C982 VN.t2 VSUBS 2.76373f
C983 VN.n14 VSUBS 1.02195f
C984 VN.t5 VSUBS 2.63528f
C985 VN.n15 VSUBS 1.00299f
C986 VN.n16 VSUBS 0.051991f
C987 VN.n17 VSUBS 0.235347f
C988 VN.n18 VSUBS 0.036855f
C989 VN.n19 VSUBS 0.036855f
C990 VN.n20 VSUBS 0.057656f
C991 VN.n21 VSUBS 0.047219f
C992 VN.n22 VSUBS 1.01123f
C993 VN.n23 VSUBS 1.91067f
C994 VTAIL.t1 VSUBS 0.353165f
C995 VTAIL.t0 VSUBS 0.353165f
C996 VTAIL.n0 VSUBS 2.764f
C997 VTAIL.n1 VSUBS 0.786042f
C998 VTAIL.n2 VSUBS 0.03098f
C999 VTAIL.n3 VSUBS 0.027452f
C1000 VTAIL.n4 VSUBS 0.014751f
C1001 VTAIL.n5 VSUBS 0.034867f
C1002 VTAIL.n6 VSUBS 0.015619f
C1003 VTAIL.n7 VSUBS 0.027452f
C1004 VTAIL.n8 VSUBS 0.015185f
C1005 VTAIL.n9 VSUBS 0.034867f
C1006 VTAIL.n10 VSUBS 0.015619f
C1007 VTAIL.n11 VSUBS 0.027452f
C1008 VTAIL.n12 VSUBS 0.014751f
C1009 VTAIL.n13 VSUBS 0.034867f
C1010 VTAIL.n14 VSUBS 0.015619f
C1011 VTAIL.n15 VSUBS 0.027452f
C1012 VTAIL.n16 VSUBS 0.014751f
C1013 VTAIL.n17 VSUBS 0.034867f
C1014 VTAIL.n18 VSUBS 0.015619f
C1015 VTAIL.n19 VSUBS 0.027452f
C1016 VTAIL.n20 VSUBS 0.014751f
C1017 VTAIL.n21 VSUBS 0.034867f
C1018 VTAIL.n22 VSUBS 0.015619f
C1019 VTAIL.n23 VSUBS 0.027452f
C1020 VTAIL.n24 VSUBS 0.014751f
C1021 VTAIL.n25 VSUBS 0.034867f
C1022 VTAIL.n26 VSUBS 0.015619f
C1023 VTAIL.n27 VSUBS 0.027452f
C1024 VTAIL.n28 VSUBS 0.014751f
C1025 VTAIL.n29 VSUBS 0.02615f
C1026 VTAIL.n30 VSUBS 0.022181f
C1027 VTAIL.t7 VSUBS 0.07473f
C1028 VTAIL.n31 VSUBS 0.203875f
C1029 VTAIL.n32 VSUBS 1.91237f
C1030 VTAIL.n33 VSUBS 0.014751f
C1031 VTAIL.n34 VSUBS 0.015619f
C1032 VTAIL.n35 VSUBS 0.034867f
C1033 VTAIL.n36 VSUBS 0.034867f
C1034 VTAIL.n37 VSUBS 0.015619f
C1035 VTAIL.n38 VSUBS 0.014751f
C1036 VTAIL.n39 VSUBS 0.027452f
C1037 VTAIL.n40 VSUBS 0.027452f
C1038 VTAIL.n41 VSUBS 0.014751f
C1039 VTAIL.n42 VSUBS 0.015619f
C1040 VTAIL.n43 VSUBS 0.034867f
C1041 VTAIL.n44 VSUBS 0.034867f
C1042 VTAIL.n45 VSUBS 0.015619f
C1043 VTAIL.n46 VSUBS 0.014751f
C1044 VTAIL.n47 VSUBS 0.027452f
C1045 VTAIL.n48 VSUBS 0.027452f
C1046 VTAIL.n49 VSUBS 0.014751f
C1047 VTAIL.n50 VSUBS 0.015619f
C1048 VTAIL.n51 VSUBS 0.034867f
C1049 VTAIL.n52 VSUBS 0.034867f
C1050 VTAIL.n53 VSUBS 0.015619f
C1051 VTAIL.n54 VSUBS 0.014751f
C1052 VTAIL.n55 VSUBS 0.027452f
C1053 VTAIL.n56 VSUBS 0.027452f
C1054 VTAIL.n57 VSUBS 0.014751f
C1055 VTAIL.n58 VSUBS 0.015619f
C1056 VTAIL.n59 VSUBS 0.034867f
C1057 VTAIL.n60 VSUBS 0.034867f
C1058 VTAIL.n61 VSUBS 0.015619f
C1059 VTAIL.n62 VSUBS 0.014751f
C1060 VTAIL.n63 VSUBS 0.027452f
C1061 VTAIL.n64 VSUBS 0.027452f
C1062 VTAIL.n65 VSUBS 0.014751f
C1063 VTAIL.n66 VSUBS 0.015619f
C1064 VTAIL.n67 VSUBS 0.034867f
C1065 VTAIL.n68 VSUBS 0.034867f
C1066 VTAIL.n69 VSUBS 0.015619f
C1067 VTAIL.n70 VSUBS 0.014751f
C1068 VTAIL.n71 VSUBS 0.027452f
C1069 VTAIL.n72 VSUBS 0.027452f
C1070 VTAIL.n73 VSUBS 0.014751f
C1071 VTAIL.n74 VSUBS 0.014751f
C1072 VTAIL.n75 VSUBS 0.015619f
C1073 VTAIL.n76 VSUBS 0.034867f
C1074 VTAIL.n77 VSUBS 0.034867f
C1075 VTAIL.n78 VSUBS 0.034867f
C1076 VTAIL.n79 VSUBS 0.015185f
C1077 VTAIL.n80 VSUBS 0.014751f
C1078 VTAIL.n81 VSUBS 0.027452f
C1079 VTAIL.n82 VSUBS 0.027452f
C1080 VTAIL.n83 VSUBS 0.014751f
C1081 VTAIL.n84 VSUBS 0.015619f
C1082 VTAIL.n85 VSUBS 0.034867f
C1083 VTAIL.n86 VSUBS 0.087189f
C1084 VTAIL.n87 VSUBS 0.015619f
C1085 VTAIL.n88 VSUBS 0.014751f
C1086 VTAIL.n89 VSUBS 0.070954f
C1087 VTAIL.n90 VSUBS 0.044189f
C1088 VTAIL.n91 VSUBS 0.290007f
C1089 VTAIL.t10 VSUBS 0.353165f
C1090 VTAIL.t11 VSUBS 0.353165f
C1091 VTAIL.n92 VSUBS 2.764f
C1092 VTAIL.n93 VSUBS 2.6848f
C1093 VTAIL.t3 VSUBS 0.353165f
C1094 VTAIL.t4 VSUBS 0.353165f
C1095 VTAIL.n94 VSUBS 2.76402f
C1096 VTAIL.n95 VSUBS 2.68478f
C1097 VTAIL.n96 VSUBS 0.03098f
C1098 VTAIL.n97 VSUBS 0.027452f
C1099 VTAIL.n98 VSUBS 0.014751f
C1100 VTAIL.n99 VSUBS 0.034867f
C1101 VTAIL.n100 VSUBS 0.015619f
C1102 VTAIL.n101 VSUBS 0.027452f
C1103 VTAIL.n102 VSUBS 0.015185f
C1104 VTAIL.n103 VSUBS 0.034867f
C1105 VTAIL.n104 VSUBS 0.014751f
C1106 VTAIL.n105 VSUBS 0.015619f
C1107 VTAIL.n106 VSUBS 0.027452f
C1108 VTAIL.n107 VSUBS 0.014751f
C1109 VTAIL.n108 VSUBS 0.034867f
C1110 VTAIL.n109 VSUBS 0.015619f
C1111 VTAIL.n110 VSUBS 0.027452f
C1112 VTAIL.n111 VSUBS 0.014751f
C1113 VTAIL.n112 VSUBS 0.034867f
C1114 VTAIL.n113 VSUBS 0.015619f
C1115 VTAIL.n114 VSUBS 0.027452f
C1116 VTAIL.n115 VSUBS 0.014751f
C1117 VTAIL.n116 VSUBS 0.034867f
C1118 VTAIL.n117 VSUBS 0.015619f
C1119 VTAIL.n118 VSUBS 0.027452f
C1120 VTAIL.n119 VSUBS 0.014751f
C1121 VTAIL.n120 VSUBS 0.034867f
C1122 VTAIL.n121 VSUBS 0.015619f
C1123 VTAIL.n122 VSUBS 0.027452f
C1124 VTAIL.n123 VSUBS 0.014751f
C1125 VTAIL.n124 VSUBS 0.02615f
C1126 VTAIL.n125 VSUBS 0.022181f
C1127 VTAIL.t5 VSUBS 0.07473f
C1128 VTAIL.n126 VSUBS 0.203875f
C1129 VTAIL.n127 VSUBS 1.91237f
C1130 VTAIL.n128 VSUBS 0.014751f
C1131 VTAIL.n129 VSUBS 0.015619f
C1132 VTAIL.n130 VSUBS 0.034867f
C1133 VTAIL.n131 VSUBS 0.034867f
C1134 VTAIL.n132 VSUBS 0.015619f
C1135 VTAIL.n133 VSUBS 0.014751f
C1136 VTAIL.n134 VSUBS 0.027452f
C1137 VTAIL.n135 VSUBS 0.027452f
C1138 VTAIL.n136 VSUBS 0.014751f
C1139 VTAIL.n137 VSUBS 0.015619f
C1140 VTAIL.n138 VSUBS 0.034867f
C1141 VTAIL.n139 VSUBS 0.034867f
C1142 VTAIL.n140 VSUBS 0.015619f
C1143 VTAIL.n141 VSUBS 0.014751f
C1144 VTAIL.n142 VSUBS 0.027452f
C1145 VTAIL.n143 VSUBS 0.027452f
C1146 VTAIL.n144 VSUBS 0.014751f
C1147 VTAIL.n145 VSUBS 0.015619f
C1148 VTAIL.n146 VSUBS 0.034867f
C1149 VTAIL.n147 VSUBS 0.034867f
C1150 VTAIL.n148 VSUBS 0.015619f
C1151 VTAIL.n149 VSUBS 0.014751f
C1152 VTAIL.n150 VSUBS 0.027452f
C1153 VTAIL.n151 VSUBS 0.027452f
C1154 VTAIL.n152 VSUBS 0.014751f
C1155 VTAIL.n153 VSUBS 0.015619f
C1156 VTAIL.n154 VSUBS 0.034867f
C1157 VTAIL.n155 VSUBS 0.034867f
C1158 VTAIL.n156 VSUBS 0.015619f
C1159 VTAIL.n157 VSUBS 0.014751f
C1160 VTAIL.n158 VSUBS 0.027452f
C1161 VTAIL.n159 VSUBS 0.027452f
C1162 VTAIL.n160 VSUBS 0.014751f
C1163 VTAIL.n161 VSUBS 0.015619f
C1164 VTAIL.n162 VSUBS 0.034867f
C1165 VTAIL.n163 VSUBS 0.034867f
C1166 VTAIL.n164 VSUBS 0.015619f
C1167 VTAIL.n165 VSUBS 0.014751f
C1168 VTAIL.n166 VSUBS 0.027452f
C1169 VTAIL.n167 VSUBS 0.027452f
C1170 VTAIL.n168 VSUBS 0.014751f
C1171 VTAIL.n169 VSUBS 0.015619f
C1172 VTAIL.n170 VSUBS 0.034867f
C1173 VTAIL.n171 VSUBS 0.034867f
C1174 VTAIL.n172 VSUBS 0.034867f
C1175 VTAIL.n173 VSUBS 0.015185f
C1176 VTAIL.n174 VSUBS 0.014751f
C1177 VTAIL.n175 VSUBS 0.027452f
C1178 VTAIL.n176 VSUBS 0.027452f
C1179 VTAIL.n177 VSUBS 0.014751f
C1180 VTAIL.n178 VSUBS 0.015619f
C1181 VTAIL.n179 VSUBS 0.034867f
C1182 VTAIL.n180 VSUBS 0.087189f
C1183 VTAIL.n181 VSUBS 0.015619f
C1184 VTAIL.n182 VSUBS 0.014751f
C1185 VTAIL.n183 VSUBS 0.070954f
C1186 VTAIL.n184 VSUBS 0.044189f
C1187 VTAIL.n185 VSUBS 0.290007f
C1188 VTAIL.t6 VSUBS 0.353165f
C1189 VTAIL.t9 VSUBS 0.353165f
C1190 VTAIL.n186 VSUBS 2.76402f
C1191 VTAIL.n187 VSUBS 0.891258f
C1192 VTAIL.n188 VSUBS 0.03098f
C1193 VTAIL.n189 VSUBS 0.027452f
C1194 VTAIL.n190 VSUBS 0.014751f
C1195 VTAIL.n191 VSUBS 0.034867f
C1196 VTAIL.n192 VSUBS 0.015619f
C1197 VTAIL.n193 VSUBS 0.027452f
C1198 VTAIL.n194 VSUBS 0.015185f
C1199 VTAIL.n195 VSUBS 0.034867f
C1200 VTAIL.n196 VSUBS 0.014751f
C1201 VTAIL.n197 VSUBS 0.015619f
C1202 VTAIL.n198 VSUBS 0.027452f
C1203 VTAIL.n199 VSUBS 0.014751f
C1204 VTAIL.n200 VSUBS 0.034867f
C1205 VTAIL.n201 VSUBS 0.015619f
C1206 VTAIL.n202 VSUBS 0.027452f
C1207 VTAIL.n203 VSUBS 0.014751f
C1208 VTAIL.n204 VSUBS 0.034867f
C1209 VTAIL.n205 VSUBS 0.015619f
C1210 VTAIL.n206 VSUBS 0.027452f
C1211 VTAIL.n207 VSUBS 0.014751f
C1212 VTAIL.n208 VSUBS 0.034867f
C1213 VTAIL.n209 VSUBS 0.015619f
C1214 VTAIL.n210 VSUBS 0.027452f
C1215 VTAIL.n211 VSUBS 0.014751f
C1216 VTAIL.n212 VSUBS 0.034867f
C1217 VTAIL.n213 VSUBS 0.015619f
C1218 VTAIL.n214 VSUBS 0.027452f
C1219 VTAIL.n215 VSUBS 0.014751f
C1220 VTAIL.n216 VSUBS 0.02615f
C1221 VTAIL.n217 VSUBS 0.022181f
C1222 VTAIL.t8 VSUBS 0.07473f
C1223 VTAIL.n218 VSUBS 0.203875f
C1224 VTAIL.n219 VSUBS 1.91237f
C1225 VTAIL.n220 VSUBS 0.014751f
C1226 VTAIL.n221 VSUBS 0.015619f
C1227 VTAIL.n222 VSUBS 0.034867f
C1228 VTAIL.n223 VSUBS 0.034867f
C1229 VTAIL.n224 VSUBS 0.015619f
C1230 VTAIL.n225 VSUBS 0.014751f
C1231 VTAIL.n226 VSUBS 0.027452f
C1232 VTAIL.n227 VSUBS 0.027452f
C1233 VTAIL.n228 VSUBS 0.014751f
C1234 VTAIL.n229 VSUBS 0.015619f
C1235 VTAIL.n230 VSUBS 0.034867f
C1236 VTAIL.n231 VSUBS 0.034867f
C1237 VTAIL.n232 VSUBS 0.015619f
C1238 VTAIL.n233 VSUBS 0.014751f
C1239 VTAIL.n234 VSUBS 0.027452f
C1240 VTAIL.n235 VSUBS 0.027452f
C1241 VTAIL.n236 VSUBS 0.014751f
C1242 VTAIL.n237 VSUBS 0.015619f
C1243 VTAIL.n238 VSUBS 0.034867f
C1244 VTAIL.n239 VSUBS 0.034867f
C1245 VTAIL.n240 VSUBS 0.015619f
C1246 VTAIL.n241 VSUBS 0.014751f
C1247 VTAIL.n242 VSUBS 0.027452f
C1248 VTAIL.n243 VSUBS 0.027452f
C1249 VTAIL.n244 VSUBS 0.014751f
C1250 VTAIL.n245 VSUBS 0.015619f
C1251 VTAIL.n246 VSUBS 0.034867f
C1252 VTAIL.n247 VSUBS 0.034867f
C1253 VTAIL.n248 VSUBS 0.015619f
C1254 VTAIL.n249 VSUBS 0.014751f
C1255 VTAIL.n250 VSUBS 0.027452f
C1256 VTAIL.n251 VSUBS 0.027452f
C1257 VTAIL.n252 VSUBS 0.014751f
C1258 VTAIL.n253 VSUBS 0.015619f
C1259 VTAIL.n254 VSUBS 0.034867f
C1260 VTAIL.n255 VSUBS 0.034867f
C1261 VTAIL.n256 VSUBS 0.015619f
C1262 VTAIL.n257 VSUBS 0.014751f
C1263 VTAIL.n258 VSUBS 0.027452f
C1264 VTAIL.n259 VSUBS 0.027452f
C1265 VTAIL.n260 VSUBS 0.014751f
C1266 VTAIL.n261 VSUBS 0.015619f
C1267 VTAIL.n262 VSUBS 0.034867f
C1268 VTAIL.n263 VSUBS 0.034867f
C1269 VTAIL.n264 VSUBS 0.034867f
C1270 VTAIL.n265 VSUBS 0.015185f
C1271 VTAIL.n266 VSUBS 0.014751f
C1272 VTAIL.n267 VSUBS 0.027452f
C1273 VTAIL.n268 VSUBS 0.027452f
C1274 VTAIL.n269 VSUBS 0.014751f
C1275 VTAIL.n270 VSUBS 0.015619f
C1276 VTAIL.n271 VSUBS 0.034867f
C1277 VTAIL.n272 VSUBS 0.087189f
C1278 VTAIL.n273 VSUBS 0.015619f
C1279 VTAIL.n274 VSUBS 0.014751f
C1280 VTAIL.n275 VSUBS 0.070954f
C1281 VTAIL.n276 VSUBS 0.044189f
C1282 VTAIL.n277 VSUBS 1.93636f
C1283 VTAIL.n278 VSUBS 0.03098f
C1284 VTAIL.n279 VSUBS 0.027452f
C1285 VTAIL.n280 VSUBS 0.014751f
C1286 VTAIL.n281 VSUBS 0.034867f
C1287 VTAIL.n282 VSUBS 0.015619f
C1288 VTAIL.n283 VSUBS 0.027452f
C1289 VTAIL.n284 VSUBS 0.015185f
C1290 VTAIL.n285 VSUBS 0.034867f
C1291 VTAIL.n286 VSUBS 0.015619f
C1292 VTAIL.n287 VSUBS 0.027452f
C1293 VTAIL.n288 VSUBS 0.014751f
C1294 VTAIL.n289 VSUBS 0.034867f
C1295 VTAIL.n290 VSUBS 0.015619f
C1296 VTAIL.n291 VSUBS 0.027452f
C1297 VTAIL.n292 VSUBS 0.014751f
C1298 VTAIL.n293 VSUBS 0.034867f
C1299 VTAIL.n294 VSUBS 0.015619f
C1300 VTAIL.n295 VSUBS 0.027452f
C1301 VTAIL.n296 VSUBS 0.014751f
C1302 VTAIL.n297 VSUBS 0.034867f
C1303 VTAIL.n298 VSUBS 0.015619f
C1304 VTAIL.n299 VSUBS 0.027452f
C1305 VTAIL.n300 VSUBS 0.014751f
C1306 VTAIL.n301 VSUBS 0.034867f
C1307 VTAIL.n302 VSUBS 0.015619f
C1308 VTAIL.n303 VSUBS 0.027452f
C1309 VTAIL.n304 VSUBS 0.014751f
C1310 VTAIL.n305 VSUBS 0.02615f
C1311 VTAIL.n306 VSUBS 0.022181f
C1312 VTAIL.t2 VSUBS 0.07473f
C1313 VTAIL.n307 VSUBS 0.203875f
C1314 VTAIL.n308 VSUBS 1.91237f
C1315 VTAIL.n309 VSUBS 0.014751f
C1316 VTAIL.n310 VSUBS 0.015619f
C1317 VTAIL.n311 VSUBS 0.034867f
C1318 VTAIL.n312 VSUBS 0.034867f
C1319 VTAIL.n313 VSUBS 0.015619f
C1320 VTAIL.n314 VSUBS 0.014751f
C1321 VTAIL.n315 VSUBS 0.027452f
C1322 VTAIL.n316 VSUBS 0.027452f
C1323 VTAIL.n317 VSUBS 0.014751f
C1324 VTAIL.n318 VSUBS 0.015619f
C1325 VTAIL.n319 VSUBS 0.034867f
C1326 VTAIL.n320 VSUBS 0.034867f
C1327 VTAIL.n321 VSUBS 0.015619f
C1328 VTAIL.n322 VSUBS 0.014751f
C1329 VTAIL.n323 VSUBS 0.027452f
C1330 VTAIL.n324 VSUBS 0.027452f
C1331 VTAIL.n325 VSUBS 0.014751f
C1332 VTAIL.n326 VSUBS 0.015619f
C1333 VTAIL.n327 VSUBS 0.034867f
C1334 VTAIL.n328 VSUBS 0.034867f
C1335 VTAIL.n329 VSUBS 0.015619f
C1336 VTAIL.n330 VSUBS 0.014751f
C1337 VTAIL.n331 VSUBS 0.027452f
C1338 VTAIL.n332 VSUBS 0.027452f
C1339 VTAIL.n333 VSUBS 0.014751f
C1340 VTAIL.n334 VSUBS 0.015619f
C1341 VTAIL.n335 VSUBS 0.034867f
C1342 VTAIL.n336 VSUBS 0.034867f
C1343 VTAIL.n337 VSUBS 0.015619f
C1344 VTAIL.n338 VSUBS 0.014751f
C1345 VTAIL.n339 VSUBS 0.027452f
C1346 VTAIL.n340 VSUBS 0.027452f
C1347 VTAIL.n341 VSUBS 0.014751f
C1348 VTAIL.n342 VSUBS 0.015619f
C1349 VTAIL.n343 VSUBS 0.034867f
C1350 VTAIL.n344 VSUBS 0.034867f
C1351 VTAIL.n345 VSUBS 0.015619f
C1352 VTAIL.n346 VSUBS 0.014751f
C1353 VTAIL.n347 VSUBS 0.027452f
C1354 VTAIL.n348 VSUBS 0.027452f
C1355 VTAIL.n349 VSUBS 0.014751f
C1356 VTAIL.n350 VSUBS 0.014751f
C1357 VTAIL.n351 VSUBS 0.015619f
C1358 VTAIL.n352 VSUBS 0.034867f
C1359 VTAIL.n353 VSUBS 0.034867f
C1360 VTAIL.n354 VSUBS 0.034867f
C1361 VTAIL.n355 VSUBS 0.015185f
C1362 VTAIL.n356 VSUBS 0.014751f
C1363 VTAIL.n357 VSUBS 0.027452f
C1364 VTAIL.n358 VSUBS 0.027452f
C1365 VTAIL.n359 VSUBS 0.014751f
C1366 VTAIL.n360 VSUBS 0.015619f
C1367 VTAIL.n361 VSUBS 0.034867f
C1368 VTAIL.n362 VSUBS 0.087189f
C1369 VTAIL.n363 VSUBS 0.015619f
C1370 VTAIL.n364 VSUBS 0.014751f
C1371 VTAIL.n365 VSUBS 0.070954f
C1372 VTAIL.n366 VSUBS 0.044189f
C1373 VTAIL.n367 VSUBS 1.89442f
C1374 VDD1.n0 VSUBS 0.030673f
C1375 VDD1.n1 VSUBS 0.02718f
C1376 VDD1.n2 VSUBS 0.014605f
C1377 VDD1.n3 VSUBS 0.034522f
C1378 VDD1.n4 VSUBS 0.015465f
C1379 VDD1.n5 VSUBS 0.02718f
C1380 VDD1.n6 VSUBS 0.015035f
C1381 VDD1.n7 VSUBS 0.034522f
C1382 VDD1.n8 VSUBS 0.014605f
C1383 VDD1.n9 VSUBS 0.015465f
C1384 VDD1.n10 VSUBS 0.02718f
C1385 VDD1.n11 VSUBS 0.014605f
C1386 VDD1.n12 VSUBS 0.034522f
C1387 VDD1.n13 VSUBS 0.015465f
C1388 VDD1.n14 VSUBS 0.02718f
C1389 VDD1.n15 VSUBS 0.014605f
C1390 VDD1.n16 VSUBS 0.034522f
C1391 VDD1.n17 VSUBS 0.015465f
C1392 VDD1.n18 VSUBS 0.02718f
C1393 VDD1.n19 VSUBS 0.014605f
C1394 VDD1.n20 VSUBS 0.034522f
C1395 VDD1.n21 VSUBS 0.015465f
C1396 VDD1.n22 VSUBS 0.02718f
C1397 VDD1.n23 VSUBS 0.014605f
C1398 VDD1.n24 VSUBS 0.034522f
C1399 VDD1.n25 VSUBS 0.015465f
C1400 VDD1.n26 VSUBS 0.02718f
C1401 VDD1.n27 VSUBS 0.014605f
C1402 VDD1.n28 VSUBS 0.025891f
C1403 VDD1.n29 VSUBS 0.021961f
C1404 VDD1.t3 VSUBS 0.073991f
C1405 VDD1.n30 VSUBS 0.201858f
C1406 VDD1.n31 VSUBS 1.89345f
C1407 VDD1.n32 VSUBS 0.014605f
C1408 VDD1.n33 VSUBS 0.015465f
C1409 VDD1.n34 VSUBS 0.034522f
C1410 VDD1.n35 VSUBS 0.034522f
C1411 VDD1.n36 VSUBS 0.015465f
C1412 VDD1.n37 VSUBS 0.014605f
C1413 VDD1.n38 VSUBS 0.02718f
C1414 VDD1.n39 VSUBS 0.02718f
C1415 VDD1.n40 VSUBS 0.014605f
C1416 VDD1.n41 VSUBS 0.015465f
C1417 VDD1.n42 VSUBS 0.034522f
C1418 VDD1.n43 VSUBS 0.034522f
C1419 VDD1.n44 VSUBS 0.015465f
C1420 VDD1.n45 VSUBS 0.014605f
C1421 VDD1.n46 VSUBS 0.02718f
C1422 VDD1.n47 VSUBS 0.02718f
C1423 VDD1.n48 VSUBS 0.014605f
C1424 VDD1.n49 VSUBS 0.015465f
C1425 VDD1.n50 VSUBS 0.034522f
C1426 VDD1.n51 VSUBS 0.034522f
C1427 VDD1.n52 VSUBS 0.015465f
C1428 VDD1.n53 VSUBS 0.014605f
C1429 VDD1.n54 VSUBS 0.02718f
C1430 VDD1.n55 VSUBS 0.02718f
C1431 VDD1.n56 VSUBS 0.014605f
C1432 VDD1.n57 VSUBS 0.015465f
C1433 VDD1.n58 VSUBS 0.034522f
C1434 VDD1.n59 VSUBS 0.034522f
C1435 VDD1.n60 VSUBS 0.015465f
C1436 VDD1.n61 VSUBS 0.014605f
C1437 VDD1.n62 VSUBS 0.02718f
C1438 VDD1.n63 VSUBS 0.02718f
C1439 VDD1.n64 VSUBS 0.014605f
C1440 VDD1.n65 VSUBS 0.015465f
C1441 VDD1.n66 VSUBS 0.034522f
C1442 VDD1.n67 VSUBS 0.034522f
C1443 VDD1.n68 VSUBS 0.015465f
C1444 VDD1.n69 VSUBS 0.014605f
C1445 VDD1.n70 VSUBS 0.02718f
C1446 VDD1.n71 VSUBS 0.02718f
C1447 VDD1.n72 VSUBS 0.014605f
C1448 VDD1.n73 VSUBS 0.015465f
C1449 VDD1.n74 VSUBS 0.034522f
C1450 VDD1.n75 VSUBS 0.034522f
C1451 VDD1.n76 VSUBS 0.034522f
C1452 VDD1.n77 VSUBS 0.015035f
C1453 VDD1.n78 VSUBS 0.014605f
C1454 VDD1.n79 VSUBS 0.02718f
C1455 VDD1.n80 VSUBS 0.02718f
C1456 VDD1.n81 VSUBS 0.014605f
C1457 VDD1.n82 VSUBS 0.015465f
C1458 VDD1.n83 VSUBS 0.034522f
C1459 VDD1.n84 VSUBS 0.086326f
C1460 VDD1.n85 VSUBS 0.015465f
C1461 VDD1.n86 VSUBS 0.014605f
C1462 VDD1.n87 VSUBS 0.070252f
C1463 VDD1.n88 VSUBS 0.066599f
C1464 VDD1.n89 VSUBS 0.030673f
C1465 VDD1.n90 VSUBS 0.02718f
C1466 VDD1.n91 VSUBS 0.014605f
C1467 VDD1.n92 VSUBS 0.034522f
C1468 VDD1.n93 VSUBS 0.015465f
C1469 VDD1.n94 VSUBS 0.02718f
C1470 VDD1.n95 VSUBS 0.015035f
C1471 VDD1.n96 VSUBS 0.034522f
C1472 VDD1.n97 VSUBS 0.015465f
C1473 VDD1.n98 VSUBS 0.02718f
C1474 VDD1.n99 VSUBS 0.014605f
C1475 VDD1.n100 VSUBS 0.034522f
C1476 VDD1.n101 VSUBS 0.015465f
C1477 VDD1.n102 VSUBS 0.02718f
C1478 VDD1.n103 VSUBS 0.014605f
C1479 VDD1.n104 VSUBS 0.034522f
C1480 VDD1.n105 VSUBS 0.015465f
C1481 VDD1.n106 VSUBS 0.02718f
C1482 VDD1.n107 VSUBS 0.014605f
C1483 VDD1.n108 VSUBS 0.034522f
C1484 VDD1.n109 VSUBS 0.015465f
C1485 VDD1.n110 VSUBS 0.02718f
C1486 VDD1.n111 VSUBS 0.014605f
C1487 VDD1.n112 VSUBS 0.034522f
C1488 VDD1.n113 VSUBS 0.015465f
C1489 VDD1.n114 VSUBS 0.02718f
C1490 VDD1.n115 VSUBS 0.014605f
C1491 VDD1.n116 VSUBS 0.025891f
C1492 VDD1.n117 VSUBS 0.021961f
C1493 VDD1.t0 VSUBS 0.073991f
C1494 VDD1.n118 VSUBS 0.201858f
C1495 VDD1.n119 VSUBS 1.89345f
C1496 VDD1.n120 VSUBS 0.014605f
C1497 VDD1.n121 VSUBS 0.015465f
C1498 VDD1.n122 VSUBS 0.034522f
C1499 VDD1.n123 VSUBS 0.034522f
C1500 VDD1.n124 VSUBS 0.015465f
C1501 VDD1.n125 VSUBS 0.014605f
C1502 VDD1.n126 VSUBS 0.02718f
C1503 VDD1.n127 VSUBS 0.02718f
C1504 VDD1.n128 VSUBS 0.014605f
C1505 VDD1.n129 VSUBS 0.015465f
C1506 VDD1.n130 VSUBS 0.034522f
C1507 VDD1.n131 VSUBS 0.034522f
C1508 VDD1.n132 VSUBS 0.015465f
C1509 VDD1.n133 VSUBS 0.014605f
C1510 VDD1.n134 VSUBS 0.02718f
C1511 VDD1.n135 VSUBS 0.02718f
C1512 VDD1.n136 VSUBS 0.014605f
C1513 VDD1.n137 VSUBS 0.015465f
C1514 VDD1.n138 VSUBS 0.034522f
C1515 VDD1.n139 VSUBS 0.034522f
C1516 VDD1.n140 VSUBS 0.015465f
C1517 VDD1.n141 VSUBS 0.014605f
C1518 VDD1.n142 VSUBS 0.02718f
C1519 VDD1.n143 VSUBS 0.02718f
C1520 VDD1.n144 VSUBS 0.014605f
C1521 VDD1.n145 VSUBS 0.015465f
C1522 VDD1.n146 VSUBS 0.034522f
C1523 VDD1.n147 VSUBS 0.034522f
C1524 VDD1.n148 VSUBS 0.015465f
C1525 VDD1.n149 VSUBS 0.014605f
C1526 VDD1.n150 VSUBS 0.02718f
C1527 VDD1.n151 VSUBS 0.02718f
C1528 VDD1.n152 VSUBS 0.014605f
C1529 VDD1.n153 VSUBS 0.015465f
C1530 VDD1.n154 VSUBS 0.034522f
C1531 VDD1.n155 VSUBS 0.034522f
C1532 VDD1.n156 VSUBS 0.015465f
C1533 VDD1.n157 VSUBS 0.014605f
C1534 VDD1.n158 VSUBS 0.02718f
C1535 VDD1.n159 VSUBS 0.02718f
C1536 VDD1.n160 VSUBS 0.014605f
C1537 VDD1.n161 VSUBS 0.014605f
C1538 VDD1.n162 VSUBS 0.015465f
C1539 VDD1.n163 VSUBS 0.034522f
C1540 VDD1.n164 VSUBS 0.034522f
C1541 VDD1.n165 VSUBS 0.034522f
C1542 VDD1.n166 VSUBS 0.015035f
C1543 VDD1.n167 VSUBS 0.014605f
C1544 VDD1.n168 VSUBS 0.02718f
C1545 VDD1.n169 VSUBS 0.02718f
C1546 VDD1.n170 VSUBS 0.014605f
C1547 VDD1.n171 VSUBS 0.015465f
C1548 VDD1.n172 VSUBS 0.034522f
C1549 VDD1.n173 VSUBS 0.086326f
C1550 VDD1.n174 VSUBS 0.015465f
C1551 VDD1.n175 VSUBS 0.014605f
C1552 VDD1.n176 VSUBS 0.070252f
C1553 VDD1.n177 VSUBS 0.06604f
C1554 VDD1.t1 VSUBS 0.349671f
C1555 VDD1.t5 VSUBS 0.349671f
C1556 VDD1.n178 VSUBS 2.88823f
C1557 VDD1.n179 VSUBS 3.12926f
C1558 VDD1.t4 VSUBS 0.349671f
C1559 VDD1.t2 VSUBS 0.349671f
C1560 VDD1.n180 VSUBS 2.88482f
C1561 VDD1.n181 VSUBS 3.37006f
C1562 VP.n0 VSUBS 0.037743f
C1563 VP.t4 VSUBS 2.69879f
C1564 VP.n1 VSUBS 0.051631f
C1565 VP.n2 VSUBS 0.037743f
C1566 VP.t0 VSUBS 2.69879f
C1567 VP.n3 VSUBS 0.059045f
C1568 VP.n4 VSUBS 0.037743f
C1569 VP.t3 VSUBS 2.69879f
C1570 VP.n5 VSUBS 0.051631f
C1571 VP.t5 VSUBS 2.83033f
C1572 VP.n6 VSUBS 1.04658f
C1573 VP.t2 VSUBS 2.69879f
C1574 VP.n7 VSUBS 1.02716f
C1575 VP.n8 VSUBS 0.053244f
C1576 VP.n9 VSUBS 0.241019f
C1577 VP.n10 VSUBS 0.037743f
C1578 VP.n11 VSUBS 0.037743f
C1579 VP.n12 VSUBS 0.059045f
C1580 VP.n13 VSUBS 0.048357f
C1581 VP.n14 VSUBS 1.0356f
C1582 VP.n15 VSUBS 1.93212f
C1583 VP.n16 VSUBS 1.96035f
C1584 VP.t1 VSUBS 2.69879f
C1585 VP.n17 VSUBS 1.0356f
C1586 VP.n18 VSUBS 0.048357f
C1587 VP.n19 VSUBS 0.037743f
C1588 VP.n20 VSUBS 0.037743f
C1589 VP.n21 VSUBS 0.037743f
C1590 VP.n22 VSUBS 0.051631f
C1591 VP.n23 VSUBS 0.053244f
C1592 VP.n24 VSUBS 0.953306f
C1593 VP.n25 VSUBS 0.053244f
C1594 VP.n26 VSUBS 0.037743f
C1595 VP.n27 VSUBS 0.037743f
C1596 VP.n28 VSUBS 0.037743f
C1597 VP.n29 VSUBS 0.059045f
C1598 VP.n30 VSUBS 0.048357f
C1599 VP.n31 VSUBS 1.0356f
C1600 VP.n32 VSUBS 0.037198f
.ends

