* NGSPICE file created from diff_pair_sample_0924.ext - technology: sky130A

.subckt diff_pair_sample_0924 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t1 VP.t0 VTAIL.t3 w_n2142_n2734# sky130_fd_pr__pfet_01v8 ad=3.4437 pd=18.44 as=3.4437 ps=18.44 w=8.83 l=2.6
X1 B.t11 B.t9 B.t10 w_n2142_n2734# sky130_fd_pr__pfet_01v8 ad=3.4437 pd=18.44 as=0 ps=0 w=8.83 l=2.6
X2 VDD1.t0 VP.t1 VTAIL.t2 w_n2142_n2734# sky130_fd_pr__pfet_01v8 ad=3.4437 pd=18.44 as=3.4437 ps=18.44 w=8.83 l=2.6
X3 VDD2.t1 VN.t0 VTAIL.t0 w_n2142_n2734# sky130_fd_pr__pfet_01v8 ad=3.4437 pd=18.44 as=3.4437 ps=18.44 w=8.83 l=2.6
X4 VDD2.t0 VN.t1 VTAIL.t1 w_n2142_n2734# sky130_fd_pr__pfet_01v8 ad=3.4437 pd=18.44 as=3.4437 ps=18.44 w=8.83 l=2.6
X5 B.t8 B.t6 B.t7 w_n2142_n2734# sky130_fd_pr__pfet_01v8 ad=3.4437 pd=18.44 as=0 ps=0 w=8.83 l=2.6
X6 B.t5 B.t3 B.t4 w_n2142_n2734# sky130_fd_pr__pfet_01v8 ad=3.4437 pd=18.44 as=0 ps=0 w=8.83 l=2.6
X7 B.t2 B.t0 B.t1 w_n2142_n2734# sky130_fd_pr__pfet_01v8 ad=3.4437 pd=18.44 as=0 ps=0 w=8.83 l=2.6
R0 VP.n0 VP.t1 173.274
R1 VP.n0 VP.t0 131.018
R2 VP VP.n0 0.336784
R3 VTAIL.n186 VTAIL.n144 756.745
R4 VTAIL.n42 VTAIL.n0 756.745
R5 VTAIL.n138 VTAIL.n96 756.745
R6 VTAIL.n90 VTAIL.n48 756.745
R7 VTAIL.n161 VTAIL.n160 585
R8 VTAIL.n163 VTAIL.n162 585
R9 VTAIL.n156 VTAIL.n155 585
R10 VTAIL.n169 VTAIL.n168 585
R11 VTAIL.n171 VTAIL.n170 585
R12 VTAIL.n152 VTAIL.n151 585
R13 VTAIL.n177 VTAIL.n176 585
R14 VTAIL.n179 VTAIL.n178 585
R15 VTAIL.n148 VTAIL.n147 585
R16 VTAIL.n185 VTAIL.n184 585
R17 VTAIL.n187 VTAIL.n186 585
R18 VTAIL.n17 VTAIL.n16 585
R19 VTAIL.n19 VTAIL.n18 585
R20 VTAIL.n12 VTAIL.n11 585
R21 VTAIL.n25 VTAIL.n24 585
R22 VTAIL.n27 VTAIL.n26 585
R23 VTAIL.n8 VTAIL.n7 585
R24 VTAIL.n33 VTAIL.n32 585
R25 VTAIL.n35 VTAIL.n34 585
R26 VTAIL.n4 VTAIL.n3 585
R27 VTAIL.n41 VTAIL.n40 585
R28 VTAIL.n43 VTAIL.n42 585
R29 VTAIL.n139 VTAIL.n138 585
R30 VTAIL.n137 VTAIL.n136 585
R31 VTAIL.n100 VTAIL.n99 585
R32 VTAIL.n131 VTAIL.n130 585
R33 VTAIL.n129 VTAIL.n128 585
R34 VTAIL.n104 VTAIL.n103 585
R35 VTAIL.n123 VTAIL.n122 585
R36 VTAIL.n121 VTAIL.n120 585
R37 VTAIL.n108 VTAIL.n107 585
R38 VTAIL.n115 VTAIL.n114 585
R39 VTAIL.n113 VTAIL.n112 585
R40 VTAIL.n91 VTAIL.n90 585
R41 VTAIL.n89 VTAIL.n88 585
R42 VTAIL.n52 VTAIL.n51 585
R43 VTAIL.n83 VTAIL.n82 585
R44 VTAIL.n81 VTAIL.n80 585
R45 VTAIL.n56 VTAIL.n55 585
R46 VTAIL.n75 VTAIL.n74 585
R47 VTAIL.n73 VTAIL.n72 585
R48 VTAIL.n60 VTAIL.n59 585
R49 VTAIL.n67 VTAIL.n66 585
R50 VTAIL.n65 VTAIL.n64 585
R51 VTAIL.n159 VTAIL.t1 327.469
R52 VTAIL.n15 VTAIL.t3 327.469
R53 VTAIL.n111 VTAIL.t2 327.469
R54 VTAIL.n63 VTAIL.t0 327.469
R55 VTAIL.n162 VTAIL.n161 171.744
R56 VTAIL.n162 VTAIL.n155 171.744
R57 VTAIL.n169 VTAIL.n155 171.744
R58 VTAIL.n170 VTAIL.n169 171.744
R59 VTAIL.n170 VTAIL.n151 171.744
R60 VTAIL.n177 VTAIL.n151 171.744
R61 VTAIL.n178 VTAIL.n177 171.744
R62 VTAIL.n178 VTAIL.n147 171.744
R63 VTAIL.n185 VTAIL.n147 171.744
R64 VTAIL.n186 VTAIL.n185 171.744
R65 VTAIL.n18 VTAIL.n17 171.744
R66 VTAIL.n18 VTAIL.n11 171.744
R67 VTAIL.n25 VTAIL.n11 171.744
R68 VTAIL.n26 VTAIL.n25 171.744
R69 VTAIL.n26 VTAIL.n7 171.744
R70 VTAIL.n33 VTAIL.n7 171.744
R71 VTAIL.n34 VTAIL.n33 171.744
R72 VTAIL.n34 VTAIL.n3 171.744
R73 VTAIL.n41 VTAIL.n3 171.744
R74 VTAIL.n42 VTAIL.n41 171.744
R75 VTAIL.n138 VTAIL.n137 171.744
R76 VTAIL.n137 VTAIL.n99 171.744
R77 VTAIL.n130 VTAIL.n99 171.744
R78 VTAIL.n130 VTAIL.n129 171.744
R79 VTAIL.n129 VTAIL.n103 171.744
R80 VTAIL.n122 VTAIL.n103 171.744
R81 VTAIL.n122 VTAIL.n121 171.744
R82 VTAIL.n121 VTAIL.n107 171.744
R83 VTAIL.n114 VTAIL.n107 171.744
R84 VTAIL.n114 VTAIL.n113 171.744
R85 VTAIL.n90 VTAIL.n89 171.744
R86 VTAIL.n89 VTAIL.n51 171.744
R87 VTAIL.n82 VTAIL.n51 171.744
R88 VTAIL.n82 VTAIL.n81 171.744
R89 VTAIL.n81 VTAIL.n55 171.744
R90 VTAIL.n74 VTAIL.n55 171.744
R91 VTAIL.n74 VTAIL.n73 171.744
R92 VTAIL.n73 VTAIL.n59 171.744
R93 VTAIL.n66 VTAIL.n59 171.744
R94 VTAIL.n66 VTAIL.n65 171.744
R95 VTAIL.n161 VTAIL.t1 85.8723
R96 VTAIL.n17 VTAIL.t3 85.8723
R97 VTAIL.n113 VTAIL.t2 85.8723
R98 VTAIL.n65 VTAIL.t0 85.8723
R99 VTAIL.n191 VTAIL.n190 31.2157
R100 VTAIL.n47 VTAIL.n46 31.2157
R101 VTAIL.n143 VTAIL.n142 31.2157
R102 VTAIL.n95 VTAIL.n94 31.2157
R103 VTAIL.n95 VTAIL.n47 25.0307
R104 VTAIL.n191 VTAIL.n143 22.5048
R105 VTAIL.n160 VTAIL.n159 16.3894
R106 VTAIL.n16 VTAIL.n15 16.3894
R107 VTAIL.n112 VTAIL.n111 16.3894
R108 VTAIL.n64 VTAIL.n63 16.3894
R109 VTAIL.n163 VTAIL.n158 12.8005
R110 VTAIL.n19 VTAIL.n14 12.8005
R111 VTAIL.n115 VTAIL.n110 12.8005
R112 VTAIL.n67 VTAIL.n62 12.8005
R113 VTAIL.n164 VTAIL.n156 12.0247
R114 VTAIL.n20 VTAIL.n12 12.0247
R115 VTAIL.n116 VTAIL.n108 12.0247
R116 VTAIL.n68 VTAIL.n60 12.0247
R117 VTAIL.n168 VTAIL.n167 11.249
R118 VTAIL.n24 VTAIL.n23 11.249
R119 VTAIL.n120 VTAIL.n119 11.249
R120 VTAIL.n72 VTAIL.n71 11.249
R121 VTAIL.n171 VTAIL.n154 10.4732
R122 VTAIL.n27 VTAIL.n10 10.4732
R123 VTAIL.n123 VTAIL.n106 10.4732
R124 VTAIL.n75 VTAIL.n58 10.4732
R125 VTAIL.n172 VTAIL.n152 9.69747
R126 VTAIL.n28 VTAIL.n8 9.69747
R127 VTAIL.n124 VTAIL.n104 9.69747
R128 VTAIL.n76 VTAIL.n56 9.69747
R129 VTAIL.n190 VTAIL.n189 9.45567
R130 VTAIL.n46 VTAIL.n45 9.45567
R131 VTAIL.n142 VTAIL.n141 9.45567
R132 VTAIL.n94 VTAIL.n93 9.45567
R133 VTAIL.n183 VTAIL.n182 9.3005
R134 VTAIL.n146 VTAIL.n145 9.3005
R135 VTAIL.n189 VTAIL.n188 9.3005
R136 VTAIL.n150 VTAIL.n149 9.3005
R137 VTAIL.n175 VTAIL.n174 9.3005
R138 VTAIL.n173 VTAIL.n172 9.3005
R139 VTAIL.n154 VTAIL.n153 9.3005
R140 VTAIL.n167 VTAIL.n166 9.3005
R141 VTAIL.n165 VTAIL.n164 9.3005
R142 VTAIL.n158 VTAIL.n157 9.3005
R143 VTAIL.n181 VTAIL.n180 9.3005
R144 VTAIL.n39 VTAIL.n38 9.3005
R145 VTAIL.n2 VTAIL.n1 9.3005
R146 VTAIL.n45 VTAIL.n44 9.3005
R147 VTAIL.n6 VTAIL.n5 9.3005
R148 VTAIL.n31 VTAIL.n30 9.3005
R149 VTAIL.n29 VTAIL.n28 9.3005
R150 VTAIL.n10 VTAIL.n9 9.3005
R151 VTAIL.n23 VTAIL.n22 9.3005
R152 VTAIL.n21 VTAIL.n20 9.3005
R153 VTAIL.n14 VTAIL.n13 9.3005
R154 VTAIL.n37 VTAIL.n36 9.3005
R155 VTAIL.n98 VTAIL.n97 9.3005
R156 VTAIL.n135 VTAIL.n134 9.3005
R157 VTAIL.n133 VTAIL.n132 9.3005
R158 VTAIL.n102 VTAIL.n101 9.3005
R159 VTAIL.n127 VTAIL.n126 9.3005
R160 VTAIL.n125 VTAIL.n124 9.3005
R161 VTAIL.n106 VTAIL.n105 9.3005
R162 VTAIL.n119 VTAIL.n118 9.3005
R163 VTAIL.n117 VTAIL.n116 9.3005
R164 VTAIL.n110 VTAIL.n109 9.3005
R165 VTAIL.n141 VTAIL.n140 9.3005
R166 VTAIL.n50 VTAIL.n49 9.3005
R167 VTAIL.n93 VTAIL.n92 9.3005
R168 VTAIL.n87 VTAIL.n86 9.3005
R169 VTAIL.n85 VTAIL.n84 9.3005
R170 VTAIL.n54 VTAIL.n53 9.3005
R171 VTAIL.n79 VTAIL.n78 9.3005
R172 VTAIL.n77 VTAIL.n76 9.3005
R173 VTAIL.n58 VTAIL.n57 9.3005
R174 VTAIL.n71 VTAIL.n70 9.3005
R175 VTAIL.n69 VTAIL.n68 9.3005
R176 VTAIL.n62 VTAIL.n61 9.3005
R177 VTAIL.n176 VTAIL.n175 8.92171
R178 VTAIL.n190 VTAIL.n144 8.92171
R179 VTAIL.n32 VTAIL.n31 8.92171
R180 VTAIL.n46 VTAIL.n0 8.92171
R181 VTAIL.n142 VTAIL.n96 8.92171
R182 VTAIL.n128 VTAIL.n127 8.92171
R183 VTAIL.n94 VTAIL.n48 8.92171
R184 VTAIL.n80 VTAIL.n79 8.92171
R185 VTAIL.n179 VTAIL.n150 8.14595
R186 VTAIL.n188 VTAIL.n187 8.14595
R187 VTAIL.n35 VTAIL.n6 8.14595
R188 VTAIL.n44 VTAIL.n43 8.14595
R189 VTAIL.n140 VTAIL.n139 8.14595
R190 VTAIL.n131 VTAIL.n102 8.14595
R191 VTAIL.n92 VTAIL.n91 8.14595
R192 VTAIL.n83 VTAIL.n54 8.14595
R193 VTAIL.n180 VTAIL.n148 7.3702
R194 VTAIL.n184 VTAIL.n146 7.3702
R195 VTAIL.n36 VTAIL.n4 7.3702
R196 VTAIL.n40 VTAIL.n2 7.3702
R197 VTAIL.n136 VTAIL.n98 7.3702
R198 VTAIL.n132 VTAIL.n100 7.3702
R199 VTAIL.n88 VTAIL.n50 7.3702
R200 VTAIL.n84 VTAIL.n52 7.3702
R201 VTAIL.n183 VTAIL.n148 6.59444
R202 VTAIL.n184 VTAIL.n183 6.59444
R203 VTAIL.n39 VTAIL.n4 6.59444
R204 VTAIL.n40 VTAIL.n39 6.59444
R205 VTAIL.n136 VTAIL.n135 6.59444
R206 VTAIL.n135 VTAIL.n100 6.59444
R207 VTAIL.n88 VTAIL.n87 6.59444
R208 VTAIL.n87 VTAIL.n52 6.59444
R209 VTAIL.n180 VTAIL.n179 5.81868
R210 VTAIL.n187 VTAIL.n146 5.81868
R211 VTAIL.n36 VTAIL.n35 5.81868
R212 VTAIL.n43 VTAIL.n2 5.81868
R213 VTAIL.n139 VTAIL.n98 5.81868
R214 VTAIL.n132 VTAIL.n131 5.81868
R215 VTAIL.n91 VTAIL.n50 5.81868
R216 VTAIL.n84 VTAIL.n83 5.81868
R217 VTAIL.n176 VTAIL.n150 5.04292
R218 VTAIL.n188 VTAIL.n144 5.04292
R219 VTAIL.n32 VTAIL.n6 5.04292
R220 VTAIL.n44 VTAIL.n0 5.04292
R221 VTAIL.n140 VTAIL.n96 5.04292
R222 VTAIL.n128 VTAIL.n102 5.04292
R223 VTAIL.n92 VTAIL.n48 5.04292
R224 VTAIL.n80 VTAIL.n54 5.04292
R225 VTAIL.n175 VTAIL.n152 4.26717
R226 VTAIL.n31 VTAIL.n8 4.26717
R227 VTAIL.n127 VTAIL.n104 4.26717
R228 VTAIL.n79 VTAIL.n56 4.26717
R229 VTAIL.n111 VTAIL.n109 3.70987
R230 VTAIL.n63 VTAIL.n61 3.70987
R231 VTAIL.n159 VTAIL.n157 3.70987
R232 VTAIL.n15 VTAIL.n13 3.70987
R233 VTAIL.n172 VTAIL.n171 3.49141
R234 VTAIL.n28 VTAIL.n27 3.49141
R235 VTAIL.n124 VTAIL.n123 3.49141
R236 VTAIL.n76 VTAIL.n75 3.49141
R237 VTAIL.n168 VTAIL.n154 2.71565
R238 VTAIL.n24 VTAIL.n10 2.71565
R239 VTAIL.n120 VTAIL.n106 2.71565
R240 VTAIL.n72 VTAIL.n58 2.71565
R241 VTAIL.n167 VTAIL.n156 1.93989
R242 VTAIL.n23 VTAIL.n12 1.93989
R243 VTAIL.n119 VTAIL.n108 1.93989
R244 VTAIL.n71 VTAIL.n60 1.93989
R245 VTAIL.n143 VTAIL.n95 1.73326
R246 VTAIL.n164 VTAIL.n163 1.16414
R247 VTAIL.n20 VTAIL.n19 1.16414
R248 VTAIL.n116 VTAIL.n115 1.16414
R249 VTAIL.n68 VTAIL.n67 1.16414
R250 VTAIL VTAIL.n47 1.15998
R251 VTAIL VTAIL.n191 0.573776
R252 VTAIL.n160 VTAIL.n158 0.388379
R253 VTAIL.n16 VTAIL.n14 0.388379
R254 VTAIL.n112 VTAIL.n110 0.388379
R255 VTAIL.n64 VTAIL.n62 0.388379
R256 VTAIL.n165 VTAIL.n157 0.155672
R257 VTAIL.n166 VTAIL.n165 0.155672
R258 VTAIL.n166 VTAIL.n153 0.155672
R259 VTAIL.n173 VTAIL.n153 0.155672
R260 VTAIL.n174 VTAIL.n173 0.155672
R261 VTAIL.n174 VTAIL.n149 0.155672
R262 VTAIL.n181 VTAIL.n149 0.155672
R263 VTAIL.n182 VTAIL.n181 0.155672
R264 VTAIL.n182 VTAIL.n145 0.155672
R265 VTAIL.n189 VTAIL.n145 0.155672
R266 VTAIL.n21 VTAIL.n13 0.155672
R267 VTAIL.n22 VTAIL.n21 0.155672
R268 VTAIL.n22 VTAIL.n9 0.155672
R269 VTAIL.n29 VTAIL.n9 0.155672
R270 VTAIL.n30 VTAIL.n29 0.155672
R271 VTAIL.n30 VTAIL.n5 0.155672
R272 VTAIL.n37 VTAIL.n5 0.155672
R273 VTAIL.n38 VTAIL.n37 0.155672
R274 VTAIL.n38 VTAIL.n1 0.155672
R275 VTAIL.n45 VTAIL.n1 0.155672
R276 VTAIL.n141 VTAIL.n97 0.155672
R277 VTAIL.n134 VTAIL.n97 0.155672
R278 VTAIL.n134 VTAIL.n133 0.155672
R279 VTAIL.n133 VTAIL.n101 0.155672
R280 VTAIL.n126 VTAIL.n101 0.155672
R281 VTAIL.n126 VTAIL.n125 0.155672
R282 VTAIL.n125 VTAIL.n105 0.155672
R283 VTAIL.n118 VTAIL.n105 0.155672
R284 VTAIL.n118 VTAIL.n117 0.155672
R285 VTAIL.n117 VTAIL.n109 0.155672
R286 VTAIL.n93 VTAIL.n49 0.155672
R287 VTAIL.n86 VTAIL.n49 0.155672
R288 VTAIL.n86 VTAIL.n85 0.155672
R289 VTAIL.n85 VTAIL.n53 0.155672
R290 VTAIL.n78 VTAIL.n53 0.155672
R291 VTAIL.n78 VTAIL.n77 0.155672
R292 VTAIL.n77 VTAIL.n57 0.155672
R293 VTAIL.n70 VTAIL.n57 0.155672
R294 VTAIL.n70 VTAIL.n69 0.155672
R295 VTAIL.n69 VTAIL.n61 0.155672
R296 VDD1.n42 VDD1.n0 756.745
R297 VDD1.n89 VDD1.n47 756.745
R298 VDD1.n43 VDD1.n42 585
R299 VDD1.n41 VDD1.n40 585
R300 VDD1.n4 VDD1.n3 585
R301 VDD1.n35 VDD1.n34 585
R302 VDD1.n33 VDD1.n32 585
R303 VDD1.n8 VDD1.n7 585
R304 VDD1.n27 VDD1.n26 585
R305 VDD1.n25 VDD1.n24 585
R306 VDD1.n12 VDD1.n11 585
R307 VDD1.n19 VDD1.n18 585
R308 VDD1.n17 VDD1.n16 585
R309 VDD1.n64 VDD1.n63 585
R310 VDD1.n66 VDD1.n65 585
R311 VDD1.n59 VDD1.n58 585
R312 VDD1.n72 VDD1.n71 585
R313 VDD1.n74 VDD1.n73 585
R314 VDD1.n55 VDD1.n54 585
R315 VDD1.n80 VDD1.n79 585
R316 VDD1.n82 VDD1.n81 585
R317 VDD1.n51 VDD1.n50 585
R318 VDD1.n88 VDD1.n87 585
R319 VDD1.n90 VDD1.n89 585
R320 VDD1.n15 VDD1.t0 327.469
R321 VDD1.n62 VDD1.t1 327.469
R322 VDD1.n42 VDD1.n41 171.744
R323 VDD1.n41 VDD1.n3 171.744
R324 VDD1.n34 VDD1.n3 171.744
R325 VDD1.n34 VDD1.n33 171.744
R326 VDD1.n33 VDD1.n7 171.744
R327 VDD1.n26 VDD1.n7 171.744
R328 VDD1.n26 VDD1.n25 171.744
R329 VDD1.n25 VDD1.n11 171.744
R330 VDD1.n18 VDD1.n11 171.744
R331 VDD1.n18 VDD1.n17 171.744
R332 VDD1.n65 VDD1.n64 171.744
R333 VDD1.n65 VDD1.n58 171.744
R334 VDD1.n72 VDD1.n58 171.744
R335 VDD1.n73 VDD1.n72 171.744
R336 VDD1.n73 VDD1.n54 171.744
R337 VDD1.n80 VDD1.n54 171.744
R338 VDD1.n81 VDD1.n80 171.744
R339 VDD1.n81 VDD1.n50 171.744
R340 VDD1.n88 VDD1.n50 171.744
R341 VDD1.n89 VDD1.n88 171.744
R342 VDD1.n17 VDD1.t0 85.8723
R343 VDD1.n64 VDD1.t1 85.8723
R344 VDD1 VDD1.n93 85.374
R345 VDD1 VDD1.n46 48.5841
R346 VDD1.n16 VDD1.n15 16.3894
R347 VDD1.n63 VDD1.n62 16.3894
R348 VDD1.n19 VDD1.n14 12.8005
R349 VDD1.n66 VDD1.n61 12.8005
R350 VDD1.n20 VDD1.n12 12.0247
R351 VDD1.n67 VDD1.n59 12.0247
R352 VDD1.n24 VDD1.n23 11.249
R353 VDD1.n71 VDD1.n70 11.249
R354 VDD1.n27 VDD1.n10 10.4732
R355 VDD1.n74 VDD1.n57 10.4732
R356 VDD1.n28 VDD1.n8 9.69747
R357 VDD1.n75 VDD1.n55 9.69747
R358 VDD1.n46 VDD1.n45 9.45567
R359 VDD1.n93 VDD1.n92 9.45567
R360 VDD1.n2 VDD1.n1 9.3005
R361 VDD1.n39 VDD1.n38 9.3005
R362 VDD1.n37 VDD1.n36 9.3005
R363 VDD1.n6 VDD1.n5 9.3005
R364 VDD1.n31 VDD1.n30 9.3005
R365 VDD1.n29 VDD1.n28 9.3005
R366 VDD1.n10 VDD1.n9 9.3005
R367 VDD1.n23 VDD1.n22 9.3005
R368 VDD1.n21 VDD1.n20 9.3005
R369 VDD1.n14 VDD1.n13 9.3005
R370 VDD1.n45 VDD1.n44 9.3005
R371 VDD1.n86 VDD1.n85 9.3005
R372 VDD1.n49 VDD1.n48 9.3005
R373 VDD1.n92 VDD1.n91 9.3005
R374 VDD1.n53 VDD1.n52 9.3005
R375 VDD1.n78 VDD1.n77 9.3005
R376 VDD1.n76 VDD1.n75 9.3005
R377 VDD1.n57 VDD1.n56 9.3005
R378 VDD1.n70 VDD1.n69 9.3005
R379 VDD1.n68 VDD1.n67 9.3005
R380 VDD1.n61 VDD1.n60 9.3005
R381 VDD1.n84 VDD1.n83 9.3005
R382 VDD1.n46 VDD1.n0 8.92171
R383 VDD1.n32 VDD1.n31 8.92171
R384 VDD1.n79 VDD1.n78 8.92171
R385 VDD1.n93 VDD1.n47 8.92171
R386 VDD1.n44 VDD1.n43 8.14595
R387 VDD1.n35 VDD1.n6 8.14595
R388 VDD1.n82 VDD1.n53 8.14595
R389 VDD1.n91 VDD1.n90 8.14595
R390 VDD1.n40 VDD1.n2 7.3702
R391 VDD1.n36 VDD1.n4 7.3702
R392 VDD1.n83 VDD1.n51 7.3702
R393 VDD1.n87 VDD1.n49 7.3702
R394 VDD1.n40 VDD1.n39 6.59444
R395 VDD1.n39 VDD1.n4 6.59444
R396 VDD1.n86 VDD1.n51 6.59444
R397 VDD1.n87 VDD1.n86 6.59444
R398 VDD1.n43 VDD1.n2 5.81868
R399 VDD1.n36 VDD1.n35 5.81868
R400 VDD1.n83 VDD1.n82 5.81868
R401 VDD1.n90 VDD1.n49 5.81868
R402 VDD1.n44 VDD1.n0 5.04292
R403 VDD1.n32 VDD1.n6 5.04292
R404 VDD1.n79 VDD1.n53 5.04292
R405 VDD1.n91 VDD1.n47 5.04292
R406 VDD1.n31 VDD1.n8 4.26717
R407 VDD1.n78 VDD1.n55 4.26717
R408 VDD1.n15 VDD1.n13 3.70987
R409 VDD1.n62 VDD1.n60 3.70987
R410 VDD1.n28 VDD1.n27 3.49141
R411 VDD1.n75 VDD1.n74 3.49141
R412 VDD1.n24 VDD1.n10 2.71565
R413 VDD1.n71 VDD1.n57 2.71565
R414 VDD1.n23 VDD1.n12 1.93989
R415 VDD1.n70 VDD1.n59 1.93989
R416 VDD1.n20 VDD1.n19 1.16414
R417 VDD1.n67 VDD1.n66 1.16414
R418 VDD1.n16 VDD1.n14 0.388379
R419 VDD1.n63 VDD1.n61 0.388379
R420 VDD1.n45 VDD1.n1 0.155672
R421 VDD1.n38 VDD1.n1 0.155672
R422 VDD1.n38 VDD1.n37 0.155672
R423 VDD1.n37 VDD1.n5 0.155672
R424 VDD1.n30 VDD1.n5 0.155672
R425 VDD1.n30 VDD1.n29 0.155672
R426 VDD1.n29 VDD1.n9 0.155672
R427 VDD1.n22 VDD1.n9 0.155672
R428 VDD1.n22 VDD1.n21 0.155672
R429 VDD1.n21 VDD1.n13 0.155672
R430 VDD1.n68 VDD1.n60 0.155672
R431 VDD1.n69 VDD1.n68 0.155672
R432 VDD1.n69 VDD1.n56 0.155672
R433 VDD1.n76 VDD1.n56 0.155672
R434 VDD1.n77 VDD1.n76 0.155672
R435 VDD1.n77 VDD1.n52 0.155672
R436 VDD1.n84 VDD1.n52 0.155672
R437 VDD1.n85 VDD1.n84 0.155672
R438 VDD1.n85 VDD1.n48 0.155672
R439 VDD1.n92 VDD1.n48 0.155672
R440 B.n284 B.n283 585
R441 B.n282 B.n83 585
R442 B.n281 B.n280 585
R443 B.n279 B.n84 585
R444 B.n278 B.n277 585
R445 B.n276 B.n85 585
R446 B.n275 B.n274 585
R447 B.n273 B.n86 585
R448 B.n272 B.n271 585
R449 B.n270 B.n87 585
R450 B.n269 B.n268 585
R451 B.n267 B.n88 585
R452 B.n266 B.n265 585
R453 B.n264 B.n89 585
R454 B.n263 B.n262 585
R455 B.n261 B.n90 585
R456 B.n260 B.n259 585
R457 B.n258 B.n91 585
R458 B.n257 B.n256 585
R459 B.n255 B.n92 585
R460 B.n254 B.n253 585
R461 B.n252 B.n93 585
R462 B.n251 B.n250 585
R463 B.n249 B.n94 585
R464 B.n248 B.n247 585
R465 B.n246 B.n95 585
R466 B.n245 B.n244 585
R467 B.n243 B.n96 585
R468 B.n242 B.n241 585
R469 B.n240 B.n97 585
R470 B.n239 B.n238 585
R471 B.n237 B.n98 585
R472 B.n235 B.n234 585
R473 B.n233 B.n101 585
R474 B.n232 B.n231 585
R475 B.n230 B.n102 585
R476 B.n229 B.n228 585
R477 B.n227 B.n103 585
R478 B.n226 B.n225 585
R479 B.n224 B.n104 585
R480 B.n223 B.n222 585
R481 B.n221 B.n105 585
R482 B.n220 B.n219 585
R483 B.n215 B.n106 585
R484 B.n214 B.n213 585
R485 B.n212 B.n107 585
R486 B.n211 B.n210 585
R487 B.n209 B.n108 585
R488 B.n208 B.n207 585
R489 B.n206 B.n109 585
R490 B.n205 B.n204 585
R491 B.n203 B.n110 585
R492 B.n202 B.n201 585
R493 B.n200 B.n111 585
R494 B.n199 B.n198 585
R495 B.n197 B.n112 585
R496 B.n196 B.n195 585
R497 B.n194 B.n113 585
R498 B.n193 B.n192 585
R499 B.n191 B.n114 585
R500 B.n190 B.n189 585
R501 B.n188 B.n115 585
R502 B.n187 B.n186 585
R503 B.n185 B.n116 585
R504 B.n184 B.n183 585
R505 B.n182 B.n117 585
R506 B.n181 B.n180 585
R507 B.n179 B.n118 585
R508 B.n178 B.n177 585
R509 B.n176 B.n119 585
R510 B.n175 B.n174 585
R511 B.n173 B.n120 585
R512 B.n172 B.n171 585
R513 B.n170 B.n121 585
R514 B.n285 B.n82 585
R515 B.n287 B.n286 585
R516 B.n288 B.n81 585
R517 B.n290 B.n289 585
R518 B.n291 B.n80 585
R519 B.n293 B.n292 585
R520 B.n294 B.n79 585
R521 B.n296 B.n295 585
R522 B.n297 B.n78 585
R523 B.n299 B.n298 585
R524 B.n300 B.n77 585
R525 B.n302 B.n301 585
R526 B.n303 B.n76 585
R527 B.n305 B.n304 585
R528 B.n306 B.n75 585
R529 B.n308 B.n307 585
R530 B.n309 B.n74 585
R531 B.n311 B.n310 585
R532 B.n312 B.n73 585
R533 B.n314 B.n313 585
R534 B.n315 B.n72 585
R535 B.n317 B.n316 585
R536 B.n318 B.n71 585
R537 B.n320 B.n319 585
R538 B.n321 B.n70 585
R539 B.n323 B.n322 585
R540 B.n324 B.n69 585
R541 B.n326 B.n325 585
R542 B.n327 B.n68 585
R543 B.n329 B.n328 585
R544 B.n330 B.n67 585
R545 B.n332 B.n331 585
R546 B.n333 B.n66 585
R547 B.n335 B.n334 585
R548 B.n336 B.n65 585
R549 B.n338 B.n337 585
R550 B.n339 B.n64 585
R551 B.n341 B.n340 585
R552 B.n342 B.n63 585
R553 B.n344 B.n343 585
R554 B.n345 B.n62 585
R555 B.n347 B.n346 585
R556 B.n348 B.n61 585
R557 B.n350 B.n349 585
R558 B.n351 B.n60 585
R559 B.n353 B.n352 585
R560 B.n354 B.n59 585
R561 B.n356 B.n355 585
R562 B.n357 B.n58 585
R563 B.n359 B.n358 585
R564 B.n360 B.n57 585
R565 B.n362 B.n361 585
R566 B.n474 B.n473 585
R567 B.n472 B.n15 585
R568 B.n471 B.n470 585
R569 B.n469 B.n16 585
R570 B.n468 B.n467 585
R571 B.n466 B.n17 585
R572 B.n465 B.n464 585
R573 B.n463 B.n18 585
R574 B.n462 B.n461 585
R575 B.n460 B.n19 585
R576 B.n459 B.n458 585
R577 B.n457 B.n20 585
R578 B.n456 B.n455 585
R579 B.n454 B.n21 585
R580 B.n453 B.n452 585
R581 B.n451 B.n22 585
R582 B.n450 B.n449 585
R583 B.n448 B.n23 585
R584 B.n447 B.n446 585
R585 B.n445 B.n24 585
R586 B.n444 B.n443 585
R587 B.n442 B.n25 585
R588 B.n441 B.n440 585
R589 B.n439 B.n26 585
R590 B.n438 B.n437 585
R591 B.n436 B.n27 585
R592 B.n435 B.n434 585
R593 B.n433 B.n28 585
R594 B.n432 B.n431 585
R595 B.n430 B.n29 585
R596 B.n429 B.n428 585
R597 B.n427 B.n30 585
R598 B.n426 B.n425 585
R599 B.n424 B.n31 585
R600 B.n423 B.n422 585
R601 B.n421 B.n35 585
R602 B.n420 B.n419 585
R603 B.n418 B.n36 585
R604 B.n417 B.n416 585
R605 B.n415 B.n37 585
R606 B.n414 B.n413 585
R607 B.n412 B.n38 585
R608 B.n410 B.n409 585
R609 B.n408 B.n41 585
R610 B.n407 B.n406 585
R611 B.n405 B.n42 585
R612 B.n404 B.n403 585
R613 B.n402 B.n43 585
R614 B.n401 B.n400 585
R615 B.n399 B.n44 585
R616 B.n398 B.n397 585
R617 B.n396 B.n45 585
R618 B.n395 B.n394 585
R619 B.n393 B.n46 585
R620 B.n392 B.n391 585
R621 B.n390 B.n47 585
R622 B.n389 B.n388 585
R623 B.n387 B.n48 585
R624 B.n386 B.n385 585
R625 B.n384 B.n49 585
R626 B.n383 B.n382 585
R627 B.n381 B.n50 585
R628 B.n380 B.n379 585
R629 B.n378 B.n51 585
R630 B.n377 B.n376 585
R631 B.n375 B.n52 585
R632 B.n374 B.n373 585
R633 B.n372 B.n53 585
R634 B.n371 B.n370 585
R635 B.n369 B.n54 585
R636 B.n368 B.n367 585
R637 B.n366 B.n55 585
R638 B.n365 B.n364 585
R639 B.n363 B.n56 585
R640 B.n475 B.n14 585
R641 B.n477 B.n476 585
R642 B.n478 B.n13 585
R643 B.n480 B.n479 585
R644 B.n481 B.n12 585
R645 B.n483 B.n482 585
R646 B.n484 B.n11 585
R647 B.n486 B.n485 585
R648 B.n487 B.n10 585
R649 B.n489 B.n488 585
R650 B.n490 B.n9 585
R651 B.n492 B.n491 585
R652 B.n493 B.n8 585
R653 B.n495 B.n494 585
R654 B.n496 B.n7 585
R655 B.n498 B.n497 585
R656 B.n499 B.n6 585
R657 B.n501 B.n500 585
R658 B.n502 B.n5 585
R659 B.n504 B.n503 585
R660 B.n505 B.n4 585
R661 B.n507 B.n506 585
R662 B.n508 B.n3 585
R663 B.n510 B.n509 585
R664 B.n511 B.n0 585
R665 B.n2 B.n1 585
R666 B.n134 B.n133 585
R667 B.n136 B.n135 585
R668 B.n137 B.n132 585
R669 B.n139 B.n138 585
R670 B.n140 B.n131 585
R671 B.n142 B.n141 585
R672 B.n143 B.n130 585
R673 B.n145 B.n144 585
R674 B.n146 B.n129 585
R675 B.n148 B.n147 585
R676 B.n149 B.n128 585
R677 B.n151 B.n150 585
R678 B.n152 B.n127 585
R679 B.n154 B.n153 585
R680 B.n155 B.n126 585
R681 B.n157 B.n156 585
R682 B.n158 B.n125 585
R683 B.n160 B.n159 585
R684 B.n161 B.n124 585
R685 B.n163 B.n162 585
R686 B.n164 B.n123 585
R687 B.n166 B.n165 585
R688 B.n167 B.n122 585
R689 B.n169 B.n168 585
R690 B.n170 B.n169 487.695
R691 B.n283 B.n82 487.695
R692 B.n361 B.n56 487.695
R693 B.n475 B.n474 487.695
R694 B.n99 B.t7 375.627
R695 B.n39 B.t11 375.627
R696 B.n216 B.t4 375.627
R697 B.n32 B.t2 375.627
R698 B.n100 B.t8 318.803
R699 B.n40 B.t10 318.803
R700 B.n217 B.t5 318.803
R701 B.n33 B.t1 318.803
R702 B.n216 B.t3 289.894
R703 B.n99 B.t6 289.894
R704 B.n39 B.t9 289.894
R705 B.n32 B.t0 289.894
R706 B.n513 B.n512 256.663
R707 B.n512 B.n511 235.042
R708 B.n512 B.n2 235.042
R709 B.n171 B.n170 163.367
R710 B.n171 B.n120 163.367
R711 B.n175 B.n120 163.367
R712 B.n176 B.n175 163.367
R713 B.n177 B.n176 163.367
R714 B.n177 B.n118 163.367
R715 B.n181 B.n118 163.367
R716 B.n182 B.n181 163.367
R717 B.n183 B.n182 163.367
R718 B.n183 B.n116 163.367
R719 B.n187 B.n116 163.367
R720 B.n188 B.n187 163.367
R721 B.n189 B.n188 163.367
R722 B.n189 B.n114 163.367
R723 B.n193 B.n114 163.367
R724 B.n194 B.n193 163.367
R725 B.n195 B.n194 163.367
R726 B.n195 B.n112 163.367
R727 B.n199 B.n112 163.367
R728 B.n200 B.n199 163.367
R729 B.n201 B.n200 163.367
R730 B.n201 B.n110 163.367
R731 B.n205 B.n110 163.367
R732 B.n206 B.n205 163.367
R733 B.n207 B.n206 163.367
R734 B.n207 B.n108 163.367
R735 B.n211 B.n108 163.367
R736 B.n212 B.n211 163.367
R737 B.n213 B.n212 163.367
R738 B.n213 B.n106 163.367
R739 B.n220 B.n106 163.367
R740 B.n221 B.n220 163.367
R741 B.n222 B.n221 163.367
R742 B.n222 B.n104 163.367
R743 B.n226 B.n104 163.367
R744 B.n227 B.n226 163.367
R745 B.n228 B.n227 163.367
R746 B.n228 B.n102 163.367
R747 B.n232 B.n102 163.367
R748 B.n233 B.n232 163.367
R749 B.n234 B.n233 163.367
R750 B.n234 B.n98 163.367
R751 B.n239 B.n98 163.367
R752 B.n240 B.n239 163.367
R753 B.n241 B.n240 163.367
R754 B.n241 B.n96 163.367
R755 B.n245 B.n96 163.367
R756 B.n246 B.n245 163.367
R757 B.n247 B.n246 163.367
R758 B.n247 B.n94 163.367
R759 B.n251 B.n94 163.367
R760 B.n252 B.n251 163.367
R761 B.n253 B.n252 163.367
R762 B.n253 B.n92 163.367
R763 B.n257 B.n92 163.367
R764 B.n258 B.n257 163.367
R765 B.n259 B.n258 163.367
R766 B.n259 B.n90 163.367
R767 B.n263 B.n90 163.367
R768 B.n264 B.n263 163.367
R769 B.n265 B.n264 163.367
R770 B.n265 B.n88 163.367
R771 B.n269 B.n88 163.367
R772 B.n270 B.n269 163.367
R773 B.n271 B.n270 163.367
R774 B.n271 B.n86 163.367
R775 B.n275 B.n86 163.367
R776 B.n276 B.n275 163.367
R777 B.n277 B.n276 163.367
R778 B.n277 B.n84 163.367
R779 B.n281 B.n84 163.367
R780 B.n282 B.n281 163.367
R781 B.n283 B.n282 163.367
R782 B.n361 B.n360 163.367
R783 B.n360 B.n359 163.367
R784 B.n359 B.n58 163.367
R785 B.n355 B.n58 163.367
R786 B.n355 B.n354 163.367
R787 B.n354 B.n353 163.367
R788 B.n353 B.n60 163.367
R789 B.n349 B.n60 163.367
R790 B.n349 B.n348 163.367
R791 B.n348 B.n347 163.367
R792 B.n347 B.n62 163.367
R793 B.n343 B.n62 163.367
R794 B.n343 B.n342 163.367
R795 B.n342 B.n341 163.367
R796 B.n341 B.n64 163.367
R797 B.n337 B.n64 163.367
R798 B.n337 B.n336 163.367
R799 B.n336 B.n335 163.367
R800 B.n335 B.n66 163.367
R801 B.n331 B.n66 163.367
R802 B.n331 B.n330 163.367
R803 B.n330 B.n329 163.367
R804 B.n329 B.n68 163.367
R805 B.n325 B.n68 163.367
R806 B.n325 B.n324 163.367
R807 B.n324 B.n323 163.367
R808 B.n323 B.n70 163.367
R809 B.n319 B.n70 163.367
R810 B.n319 B.n318 163.367
R811 B.n318 B.n317 163.367
R812 B.n317 B.n72 163.367
R813 B.n313 B.n72 163.367
R814 B.n313 B.n312 163.367
R815 B.n312 B.n311 163.367
R816 B.n311 B.n74 163.367
R817 B.n307 B.n74 163.367
R818 B.n307 B.n306 163.367
R819 B.n306 B.n305 163.367
R820 B.n305 B.n76 163.367
R821 B.n301 B.n76 163.367
R822 B.n301 B.n300 163.367
R823 B.n300 B.n299 163.367
R824 B.n299 B.n78 163.367
R825 B.n295 B.n78 163.367
R826 B.n295 B.n294 163.367
R827 B.n294 B.n293 163.367
R828 B.n293 B.n80 163.367
R829 B.n289 B.n80 163.367
R830 B.n289 B.n288 163.367
R831 B.n288 B.n287 163.367
R832 B.n287 B.n82 163.367
R833 B.n474 B.n15 163.367
R834 B.n470 B.n15 163.367
R835 B.n470 B.n469 163.367
R836 B.n469 B.n468 163.367
R837 B.n468 B.n17 163.367
R838 B.n464 B.n17 163.367
R839 B.n464 B.n463 163.367
R840 B.n463 B.n462 163.367
R841 B.n462 B.n19 163.367
R842 B.n458 B.n19 163.367
R843 B.n458 B.n457 163.367
R844 B.n457 B.n456 163.367
R845 B.n456 B.n21 163.367
R846 B.n452 B.n21 163.367
R847 B.n452 B.n451 163.367
R848 B.n451 B.n450 163.367
R849 B.n450 B.n23 163.367
R850 B.n446 B.n23 163.367
R851 B.n446 B.n445 163.367
R852 B.n445 B.n444 163.367
R853 B.n444 B.n25 163.367
R854 B.n440 B.n25 163.367
R855 B.n440 B.n439 163.367
R856 B.n439 B.n438 163.367
R857 B.n438 B.n27 163.367
R858 B.n434 B.n27 163.367
R859 B.n434 B.n433 163.367
R860 B.n433 B.n432 163.367
R861 B.n432 B.n29 163.367
R862 B.n428 B.n29 163.367
R863 B.n428 B.n427 163.367
R864 B.n427 B.n426 163.367
R865 B.n426 B.n31 163.367
R866 B.n422 B.n31 163.367
R867 B.n422 B.n421 163.367
R868 B.n421 B.n420 163.367
R869 B.n420 B.n36 163.367
R870 B.n416 B.n36 163.367
R871 B.n416 B.n415 163.367
R872 B.n415 B.n414 163.367
R873 B.n414 B.n38 163.367
R874 B.n409 B.n38 163.367
R875 B.n409 B.n408 163.367
R876 B.n408 B.n407 163.367
R877 B.n407 B.n42 163.367
R878 B.n403 B.n42 163.367
R879 B.n403 B.n402 163.367
R880 B.n402 B.n401 163.367
R881 B.n401 B.n44 163.367
R882 B.n397 B.n44 163.367
R883 B.n397 B.n396 163.367
R884 B.n396 B.n395 163.367
R885 B.n395 B.n46 163.367
R886 B.n391 B.n46 163.367
R887 B.n391 B.n390 163.367
R888 B.n390 B.n389 163.367
R889 B.n389 B.n48 163.367
R890 B.n385 B.n48 163.367
R891 B.n385 B.n384 163.367
R892 B.n384 B.n383 163.367
R893 B.n383 B.n50 163.367
R894 B.n379 B.n50 163.367
R895 B.n379 B.n378 163.367
R896 B.n378 B.n377 163.367
R897 B.n377 B.n52 163.367
R898 B.n373 B.n52 163.367
R899 B.n373 B.n372 163.367
R900 B.n372 B.n371 163.367
R901 B.n371 B.n54 163.367
R902 B.n367 B.n54 163.367
R903 B.n367 B.n366 163.367
R904 B.n366 B.n365 163.367
R905 B.n365 B.n56 163.367
R906 B.n476 B.n475 163.367
R907 B.n476 B.n13 163.367
R908 B.n480 B.n13 163.367
R909 B.n481 B.n480 163.367
R910 B.n482 B.n481 163.367
R911 B.n482 B.n11 163.367
R912 B.n486 B.n11 163.367
R913 B.n487 B.n486 163.367
R914 B.n488 B.n487 163.367
R915 B.n488 B.n9 163.367
R916 B.n492 B.n9 163.367
R917 B.n493 B.n492 163.367
R918 B.n494 B.n493 163.367
R919 B.n494 B.n7 163.367
R920 B.n498 B.n7 163.367
R921 B.n499 B.n498 163.367
R922 B.n500 B.n499 163.367
R923 B.n500 B.n5 163.367
R924 B.n504 B.n5 163.367
R925 B.n505 B.n504 163.367
R926 B.n506 B.n505 163.367
R927 B.n506 B.n3 163.367
R928 B.n510 B.n3 163.367
R929 B.n511 B.n510 163.367
R930 B.n134 B.n2 163.367
R931 B.n135 B.n134 163.367
R932 B.n135 B.n132 163.367
R933 B.n139 B.n132 163.367
R934 B.n140 B.n139 163.367
R935 B.n141 B.n140 163.367
R936 B.n141 B.n130 163.367
R937 B.n145 B.n130 163.367
R938 B.n146 B.n145 163.367
R939 B.n147 B.n146 163.367
R940 B.n147 B.n128 163.367
R941 B.n151 B.n128 163.367
R942 B.n152 B.n151 163.367
R943 B.n153 B.n152 163.367
R944 B.n153 B.n126 163.367
R945 B.n157 B.n126 163.367
R946 B.n158 B.n157 163.367
R947 B.n159 B.n158 163.367
R948 B.n159 B.n124 163.367
R949 B.n163 B.n124 163.367
R950 B.n164 B.n163 163.367
R951 B.n165 B.n164 163.367
R952 B.n165 B.n122 163.367
R953 B.n169 B.n122 163.367
R954 B.n218 B.n217 59.5399
R955 B.n236 B.n100 59.5399
R956 B.n411 B.n40 59.5399
R957 B.n34 B.n33 59.5399
R958 B.n217 B.n216 56.8247
R959 B.n100 B.n99 56.8247
R960 B.n40 B.n39 56.8247
R961 B.n33 B.n32 56.8247
R962 B.n473 B.n14 31.6883
R963 B.n363 B.n362 31.6883
R964 B.n285 B.n284 31.6883
R965 B.n168 B.n121 31.6883
R966 B B.n513 18.0485
R967 B.n477 B.n14 10.6151
R968 B.n478 B.n477 10.6151
R969 B.n479 B.n478 10.6151
R970 B.n479 B.n12 10.6151
R971 B.n483 B.n12 10.6151
R972 B.n484 B.n483 10.6151
R973 B.n485 B.n484 10.6151
R974 B.n485 B.n10 10.6151
R975 B.n489 B.n10 10.6151
R976 B.n490 B.n489 10.6151
R977 B.n491 B.n490 10.6151
R978 B.n491 B.n8 10.6151
R979 B.n495 B.n8 10.6151
R980 B.n496 B.n495 10.6151
R981 B.n497 B.n496 10.6151
R982 B.n497 B.n6 10.6151
R983 B.n501 B.n6 10.6151
R984 B.n502 B.n501 10.6151
R985 B.n503 B.n502 10.6151
R986 B.n503 B.n4 10.6151
R987 B.n507 B.n4 10.6151
R988 B.n508 B.n507 10.6151
R989 B.n509 B.n508 10.6151
R990 B.n509 B.n0 10.6151
R991 B.n473 B.n472 10.6151
R992 B.n472 B.n471 10.6151
R993 B.n471 B.n16 10.6151
R994 B.n467 B.n16 10.6151
R995 B.n467 B.n466 10.6151
R996 B.n466 B.n465 10.6151
R997 B.n465 B.n18 10.6151
R998 B.n461 B.n18 10.6151
R999 B.n461 B.n460 10.6151
R1000 B.n460 B.n459 10.6151
R1001 B.n459 B.n20 10.6151
R1002 B.n455 B.n20 10.6151
R1003 B.n455 B.n454 10.6151
R1004 B.n454 B.n453 10.6151
R1005 B.n453 B.n22 10.6151
R1006 B.n449 B.n22 10.6151
R1007 B.n449 B.n448 10.6151
R1008 B.n448 B.n447 10.6151
R1009 B.n447 B.n24 10.6151
R1010 B.n443 B.n24 10.6151
R1011 B.n443 B.n442 10.6151
R1012 B.n442 B.n441 10.6151
R1013 B.n441 B.n26 10.6151
R1014 B.n437 B.n26 10.6151
R1015 B.n437 B.n436 10.6151
R1016 B.n436 B.n435 10.6151
R1017 B.n435 B.n28 10.6151
R1018 B.n431 B.n28 10.6151
R1019 B.n431 B.n430 10.6151
R1020 B.n430 B.n429 10.6151
R1021 B.n429 B.n30 10.6151
R1022 B.n425 B.n424 10.6151
R1023 B.n424 B.n423 10.6151
R1024 B.n423 B.n35 10.6151
R1025 B.n419 B.n35 10.6151
R1026 B.n419 B.n418 10.6151
R1027 B.n418 B.n417 10.6151
R1028 B.n417 B.n37 10.6151
R1029 B.n413 B.n37 10.6151
R1030 B.n413 B.n412 10.6151
R1031 B.n410 B.n41 10.6151
R1032 B.n406 B.n41 10.6151
R1033 B.n406 B.n405 10.6151
R1034 B.n405 B.n404 10.6151
R1035 B.n404 B.n43 10.6151
R1036 B.n400 B.n43 10.6151
R1037 B.n400 B.n399 10.6151
R1038 B.n399 B.n398 10.6151
R1039 B.n398 B.n45 10.6151
R1040 B.n394 B.n45 10.6151
R1041 B.n394 B.n393 10.6151
R1042 B.n393 B.n392 10.6151
R1043 B.n392 B.n47 10.6151
R1044 B.n388 B.n47 10.6151
R1045 B.n388 B.n387 10.6151
R1046 B.n387 B.n386 10.6151
R1047 B.n386 B.n49 10.6151
R1048 B.n382 B.n49 10.6151
R1049 B.n382 B.n381 10.6151
R1050 B.n381 B.n380 10.6151
R1051 B.n380 B.n51 10.6151
R1052 B.n376 B.n51 10.6151
R1053 B.n376 B.n375 10.6151
R1054 B.n375 B.n374 10.6151
R1055 B.n374 B.n53 10.6151
R1056 B.n370 B.n53 10.6151
R1057 B.n370 B.n369 10.6151
R1058 B.n369 B.n368 10.6151
R1059 B.n368 B.n55 10.6151
R1060 B.n364 B.n55 10.6151
R1061 B.n364 B.n363 10.6151
R1062 B.n362 B.n57 10.6151
R1063 B.n358 B.n57 10.6151
R1064 B.n358 B.n357 10.6151
R1065 B.n357 B.n356 10.6151
R1066 B.n356 B.n59 10.6151
R1067 B.n352 B.n59 10.6151
R1068 B.n352 B.n351 10.6151
R1069 B.n351 B.n350 10.6151
R1070 B.n350 B.n61 10.6151
R1071 B.n346 B.n61 10.6151
R1072 B.n346 B.n345 10.6151
R1073 B.n345 B.n344 10.6151
R1074 B.n344 B.n63 10.6151
R1075 B.n340 B.n63 10.6151
R1076 B.n340 B.n339 10.6151
R1077 B.n339 B.n338 10.6151
R1078 B.n338 B.n65 10.6151
R1079 B.n334 B.n65 10.6151
R1080 B.n334 B.n333 10.6151
R1081 B.n333 B.n332 10.6151
R1082 B.n332 B.n67 10.6151
R1083 B.n328 B.n67 10.6151
R1084 B.n328 B.n327 10.6151
R1085 B.n327 B.n326 10.6151
R1086 B.n326 B.n69 10.6151
R1087 B.n322 B.n69 10.6151
R1088 B.n322 B.n321 10.6151
R1089 B.n321 B.n320 10.6151
R1090 B.n320 B.n71 10.6151
R1091 B.n316 B.n71 10.6151
R1092 B.n316 B.n315 10.6151
R1093 B.n315 B.n314 10.6151
R1094 B.n314 B.n73 10.6151
R1095 B.n310 B.n73 10.6151
R1096 B.n310 B.n309 10.6151
R1097 B.n309 B.n308 10.6151
R1098 B.n308 B.n75 10.6151
R1099 B.n304 B.n75 10.6151
R1100 B.n304 B.n303 10.6151
R1101 B.n303 B.n302 10.6151
R1102 B.n302 B.n77 10.6151
R1103 B.n298 B.n77 10.6151
R1104 B.n298 B.n297 10.6151
R1105 B.n297 B.n296 10.6151
R1106 B.n296 B.n79 10.6151
R1107 B.n292 B.n79 10.6151
R1108 B.n292 B.n291 10.6151
R1109 B.n291 B.n290 10.6151
R1110 B.n290 B.n81 10.6151
R1111 B.n286 B.n81 10.6151
R1112 B.n286 B.n285 10.6151
R1113 B.n133 B.n1 10.6151
R1114 B.n136 B.n133 10.6151
R1115 B.n137 B.n136 10.6151
R1116 B.n138 B.n137 10.6151
R1117 B.n138 B.n131 10.6151
R1118 B.n142 B.n131 10.6151
R1119 B.n143 B.n142 10.6151
R1120 B.n144 B.n143 10.6151
R1121 B.n144 B.n129 10.6151
R1122 B.n148 B.n129 10.6151
R1123 B.n149 B.n148 10.6151
R1124 B.n150 B.n149 10.6151
R1125 B.n150 B.n127 10.6151
R1126 B.n154 B.n127 10.6151
R1127 B.n155 B.n154 10.6151
R1128 B.n156 B.n155 10.6151
R1129 B.n156 B.n125 10.6151
R1130 B.n160 B.n125 10.6151
R1131 B.n161 B.n160 10.6151
R1132 B.n162 B.n161 10.6151
R1133 B.n162 B.n123 10.6151
R1134 B.n166 B.n123 10.6151
R1135 B.n167 B.n166 10.6151
R1136 B.n168 B.n167 10.6151
R1137 B.n172 B.n121 10.6151
R1138 B.n173 B.n172 10.6151
R1139 B.n174 B.n173 10.6151
R1140 B.n174 B.n119 10.6151
R1141 B.n178 B.n119 10.6151
R1142 B.n179 B.n178 10.6151
R1143 B.n180 B.n179 10.6151
R1144 B.n180 B.n117 10.6151
R1145 B.n184 B.n117 10.6151
R1146 B.n185 B.n184 10.6151
R1147 B.n186 B.n185 10.6151
R1148 B.n186 B.n115 10.6151
R1149 B.n190 B.n115 10.6151
R1150 B.n191 B.n190 10.6151
R1151 B.n192 B.n191 10.6151
R1152 B.n192 B.n113 10.6151
R1153 B.n196 B.n113 10.6151
R1154 B.n197 B.n196 10.6151
R1155 B.n198 B.n197 10.6151
R1156 B.n198 B.n111 10.6151
R1157 B.n202 B.n111 10.6151
R1158 B.n203 B.n202 10.6151
R1159 B.n204 B.n203 10.6151
R1160 B.n204 B.n109 10.6151
R1161 B.n208 B.n109 10.6151
R1162 B.n209 B.n208 10.6151
R1163 B.n210 B.n209 10.6151
R1164 B.n210 B.n107 10.6151
R1165 B.n214 B.n107 10.6151
R1166 B.n215 B.n214 10.6151
R1167 B.n219 B.n215 10.6151
R1168 B.n223 B.n105 10.6151
R1169 B.n224 B.n223 10.6151
R1170 B.n225 B.n224 10.6151
R1171 B.n225 B.n103 10.6151
R1172 B.n229 B.n103 10.6151
R1173 B.n230 B.n229 10.6151
R1174 B.n231 B.n230 10.6151
R1175 B.n231 B.n101 10.6151
R1176 B.n235 B.n101 10.6151
R1177 B.n238 B.n237 10.6151
R1178 B.n238 B.n97 10.6151
R1179 B.n242 B.n97 10.6151
R1180 B.n243 B.n242 10.6151
R1181 B.n244 B.n243 10.6151
R1182 B.n244 B.n95 10.6151
R1183 B.n248 B.n95 10.6151
R1184 B.n249 B.n248 10.6151
R1185 B.n250 B.n249 10.6151
R1186 B.n250 B.n93 10.6151
R1187 B.n254 B.n93 10.6151
R1188 B.n255 B.n254 10.6151
R1189 B.n256 B.n255 10.6151
R1190 B.n256 B.n91 10.6151
R1191 B.n260 B.n91 10.6151
R1192 B.n261 B.n260 10.6151
R1193 B.n262 B.n261 10.6151
R1194 B.n262 B.n89 10.6151
R1195 B.n266 B.n89 10.6151
R1196 B.n267 B.n266 10.6151
R1197 B.n268 B.n267 10.6151
R1198 B.n268 B.n87 10.6151
R1199 B.n272 B.n87 10.6151
R1200 B.n273 B.n272 10.6151
R1201 B.n274 B.n273 10.6151
R1202 B.n274 B.n85 10.6151
R1203 B.n278 B.n85 10.6151
R1204 B.n279 B.n278 10.6151
R1205 B.n280 B.n279 10.6151
R1206 B.n280 B.n83 10.6151
R1207 B.n284 B.n83 10.6151
R1208 B.n34 B.n30 9.36635
R1209 B.n411 B.n410 9.36635
R1210 B.n219 B.n218 9.36635
R1211 B.n237 B.n236 9.36635
R1212 B.n513 B.n0 8.11757
R1213 B.n513 B.n1 8.11757
R1214 B.n425 B.n34 1.24928
R1215 B.n412 B.n411 1.24928
R1216 B.n218 B.n105 1.24928
R1217 B.n236 B.n235 1.24928
R1218 VN VN.t0 173.369
R1219 VN VN.t1 131.355
R1220 VDD2.n89 VDD2.n47 756.745
R1221 VDD2.n42 VDD2.n0 756.745
R1222 VDD2.n90 VDD2.n89 585
R1223 VDD2.n88 VDD2.n87 585
R1224 VDD2.n51 VDD2.n50 585
R1225 VDD2.n82 VDD2.n81 585
R1226 VDD2.n80 VDD2.n79 585
R1227 VDD2.n55 VDD2.n54 585
R1228 VDD2.n74 VDD2.n73 585
R1229 VDD2.n72 VDD2.n71 585
R1230 VDD2.n59 VDD2.n58 585
R1231 VDD2.n66 VDD2.n65 585
R1232 VDD2.n64 VDD2.n63 585
R1233 VDD2.n17 VDD2.n16 585
R1234 VDD2.n19 VDD2.n18 585
R1235 VDD2.n12 VDD2.n11 585
R1236 VDD2.n25 VDD2.n24 585
R1237 VDD2.n27 VDD2.n26 585
R1238 VDD2.n8 VDD2.n7 585
R1239 VDD2.n33 VDD2.n32 585
R1240 VDD2.n35 VDD2.n34 585
R1241 VDD2.n4 VDD2.n3 585
R1242 VDD2.n41 VDD2.n40 585
R1243 VDD2.n43 VDD2.n42 585
R1244 VDD2.n62 VDD2.t1 327.469
R1245 VDD2.n15 VDD2.t0 327.469
R1246 VDD2.n89 VDD2.n88 171.744
R1247 VDD2.n88 VDD2.n50 171.744
R1248 VDD2.n81 VDD2.n50 171.744
R1249 VDD2.n81 VDD2.n80 171.744
R1250 VDD2.n80 VDD2.n54 171.744
R1251 VDD2.n73 VDD2.n54 171.744
R1252 VDD2.n73 VDD2.n72 171.744
R1253 VDD2.n72 VDD2.n58 171.744
R1254 VDD2.n65 VDD2.n58 171.744
R1255 VDD2.n65 VDD2.n64 171.744
R1256 VDD2.n18 VDD2.n17 171.744
R1257 VDD2.n18 VDD2.n11 171.744
R1258 VDD2.n25 VDD2.n11 171.744
R1259 VDD2.n26 VDD2.n25 171.744
R1260 VDD2.n26 VDD2.n7 171.744
R1261 VDD2.n33 VDD2.n7 171.744
R1262 VDD2.n34 VDD2.n33 171.744
R1263 VDD2.n34 VDD2.n3 171.744
R1264 VDD2.n41 VDD2.n3 171.744
R1265 VDD2.n42 VDD2.n41 171.744
R1266 VDD2.n64 VDD2.t1 85.8723
R1267 VDD2.n17 VDD2.t0 85.8723
R1268 VDD2.n94 VDD2.n46 84.2177
R1269 VDD2.n94 VDD2.n93 47.8944
R1270 VDD2.n63 VDD2.n62 16.3894
R1271 VDD2.n16 VDD2.n15 16.3894
R1272 VDD2.n66 VDD2.n61 12.8005
R1273 VDD2.n19 VDD2.n14 12.8005
R1274 VDD2.n67 VDD2.n59 12.0247
R1275 VDD2.n20 VDD2.n12 12.0247
R1276 VDD2.n71 VDD2.n70 11.249
R1277 VDD2.n24 VDD2.n23 11.249
R1278 VDD2.n74 VDD2.n57 10.4732
R1279 VDD2.n27 VDD2.n10 10.4732
R1280 VDD2.n75 VDD2.n55 9.69747
R1281 VDD2.n28 VDD2.n8 9.69747
R1282 VDD2.n93 VDD2.n92 9.45567
R1283 VDD2.n46 VDD2.n45 9.45567
R1284 VDD2.n49 VDD2.n48 9.3005
R1285 VDD2.n86 VDD2.n85 9.3005
R1286 VDD2.n84 VDD2.n83 9.3005
R1287 VDD2.n53 VDD2.n52 9.3005
R1288 VDD2.n78 VDD2.n77 9.3005
R1289 VDD2.n76 VDD2.n75 9.3005
R1290 VDD2.n57 VDD2.n56 9.3005
R1291 VDD2.n70 VDD2.n69 9.3005
R1292 VDD2.n68 VDD2.n67 9.3005
R1293 VDD2.n61 VDD2.n60 9.3005
R1294 VDD2.n92 VDD2.n91 9.3005
R1295 VDD2.n39 VDD2.n38 9.3005
R1296 VDD2.n2 VDD2.n1 9.3005
R1297 VDD2.n45 VDD2.n44 9.3005
R1298 VDD2.n6 VDD2.n5 9.3005
R1299 VDD2.n31 VDD2.n30 9.3005
R1300 VDD2.n29 VDD2.n28 9.3005
R1301 VDD2.n10 VDD2.n9 9.3005
R1302 VDD2.n23 VDD2.n22 9.3005
R1303 VDD2.n21 VDD2.n20 9.3005
R1304 VDD2.n14 VDD2.n13 9.3005
R1305 VDD2.n37 VDD2.n36 9.3005
R1306 VDD2.n93 VDD2.n47 8.92171
R1307 VDD2.n79 VDD2.n78 8.92171
R1308 VDD2.n32 VDD2.n31 8.92171
R1309 VDD2.n46 VDD2.n0 8.92171
R1310 VDD2.n91 VDD2.n90 8.14595
R1311 VDD2.n82 VDD2.n53 8.14595
R1312 VDD2.n35 VDD2.n6 8.14595
R1313 VDD2.n44 VDD2.n43 8.14595
R1314 VDD2.n87 VDD2.n49 7.3702
R1315 VDD2.n83 VDD2.n51 7.3702
R1316 VDD2.n36 VDD2.n4 7.3702
R1317 VDD2.n40 VDD2.n2 7.3702
R1318 VDD2.n87 VDD2.n86 6.59444
R1319 VDD2.n86 VDD2.n51 6.59444
R1320 VDD2.n39 VDD2.n4 6.59444
R1321 VDD2.n40 VDD2.n39 6.59444
R1322 VDD2.n90 VDD2.n49 5.81868
R1323 VDD2.n83 VDD2.n82 5.81868
R1324 VDD2.n36 VDD2.n35 5.81868
R1325 VDD2.n43 VDD2.n2 5.81868
R1326 VDD2.n91 VDD2.n47 5.04292
R1327 VDD2.n79 VDD2.n53 5.04292
R1328 VDD2.n32 VDD2.n6 5.04292
R1329 VDD2.n44 VDD2.n0 5.04292
R1330 VDD2.n78 VDD2.n55 4.26717
R1331 VDD2.n31 VDD2.n8 4.26717
R1332 VDD2.n62 VDD2.n60 3.70987
R1333 VDD2.n15 VDD2.n13 3.70987
R1334 VDD2.n75 VDD2.n74 3.49141
R1335 VDD2.n28 VDD2.n27 3.49141
R1336 VDD2.n71 VDD2.n57 2.71565
R1337 VDD2.n24 VDD2.n10 2.71565
R1338 VDD2.n70 VDD2.n59 1.93989
R1339 VDD2.n23 VDD2.n12 1.93989
R1340 VDD2.n67 VDD2.n66 1.16414
R1341 VDD2.n20 VDD2.n19 1.16414
R1342 VDD2 VDD2.n94 0.690155
R1343 VDD2.n63 VDD2.n61 0.388379
R1344 VDD2.n16 VDD2.n14 0.388379
R1345 VDD2.n92 VDD2.n48 0.155672
R1346 VDD2.n85 VDD2.n48 0.155672
R1347 VDD2.n85 VDD2.n84 0.155672
R1348 VDD2.n84 VDD2.n52 0.155672
R1349 VDD2.n77 VDD2.n52 0.155672
R1350 VDD2.n77 VDD2.n76 0.155672
R1351 VDD2.n76 VDD2.n56 0.155672
R1352 VDD2.n69 VDD2.n56 0.155672
R1353 VDD2.n69 VDD2.n68 0.155672
R1354 VDD2.n68 VDD2.n60 0.155672
R1355 VDD2.n21 VDD2.n13 0.155672
R1356 VDD2.n22 VDD2.n21 0.155672
R1357 VDD2.n22 VDD2.n9 0.155672
R1358 VDD2.n29 VDD2.n9 0.155672
R1359 VDD2.n30 VDD2.n29 0.155672
R1360 VDD2.n30 VDD2.n5 0.155672
R1361 VDD2.n37 VDD2.n5 0.155672
R1362 VDD2.n38 VDD2.n37 0.155672
R1363 VDD2.n38 VDD2.n1 0.155672
R1364 VDD2.n45 VDD2.n1 0.155672
C0 w_n2142_n2734# VN 2.8945f
C1 VP VN 4.865149f
C2 w_n2142_n2734# VTAIL 2.30634f
C3 VP VTAIL 1.93403f
C4 B VN 1.01269f
C5 VP w_n2142_n2734# 3.16735f
C6 VDD1 VN 0.148122f
C7 VDD2 VN 2.11105f
C8 B VTAIL 2.94729f
C9 B w_n2142_n2734# 7.92025f
C10 B VP 1.46126f
C11 VDD1 VTAIL 4.22944f
C12 VDD2 VTAIL 4.28079f
C13 VDD1 w_n2142_n2734# 1.56097f
C14 VDD1 VP 2.29377f
C15 VDD2 w_n2142_n2734# 1.58685f
C16 VDD2 VP 0.332813f
C17 VDD1 B 1.455f
C18 VDD2 B 1.48508f
C19 VDD2 VDD1 0.67424f
C20 VN VTAIL 1.91979f
C21 VDD2 VSUBS 0.791391f
C22 VDD1 VSUBS 3.330133f
C23 VTAIL VSUBS 0.844205f
C24 VN VSUBS 6.42282f
C25 VP VSUBS 1.558709f
C26 B VSUBS 3.641315f
C27 w_n2142_n2734# VSUBS 72.511f
C28 VDD2.n0 VSUBS 0.023494f
C29 VDD2.n1 VSUBS 0.020586f
C30 VDD2.n2 VSUBS 0.011062f
C31 VDD2.n3 VSUBS 0.026147f
C32 VDD2.n4 VSUBS 0.011713f
C33 VDD2.n5 VSUBS 0.020586f
C34 VDD2.n6 VSUBS 0.011062f
C35 VDD2.n7 VSUBS 0.026147f
C36 VDD2.n8 VSUBS 0.011713f
C37 VDD2.n9 VSUBS 0.020586f
C38 VDD2.n10 VSUBS 0.011062f
C39 VDD2.n11 VSUBS 0.026147f
C40 VDD2.n12 VSUBS 0.011713f
C41 VDD2.n13 VSUBS 0.737678f
C42 VDD2.n14 VSUBS 0.011062f
C43 VDD2.t0 VSUBS 0.055747f
C44 VDD2.n15 VSUBS 0.107737f
C45 VDD2.n16 VSUBS 0.016633f
C46 VDD2.n17 VSUBS 0.01961f
C47 VDD2.n18 VSUBS 0.026147f
C48 VDD2.n19 VSUBS 0.011713f
C49 VDD2.n20 VSUBS 0.011062f
C50 VDD2.n21 VSUBS 0.020586f
C51 VDD2.n22 VSUBS 0.020586f
C52 VDD2.n23 VSUBS 0.011062f
C53 VDD2.n24 VSUBS 0.011713f
C54 VDD2.n25 VSUBS 0.026147f
C55 VDD2.n26 VSUBS 0.026147f
C56 VDD2.n27 VSUBS 0.011713f
C57 VDD2.n28 VSUBS 0.011062f
C58 VDD2.n29 VSUBS 0.020586f
C59 VDD2.n30 VSUBS 0.020586f
C60 VDD2.n31 VSUBS 0.011062f
C61 VDD2.n32 VSUBS 0.011713f
C62 VDD2.n33 VSUBS 0.026147f
C63 VDD2.n34 VSUBS 0.026147f
C64 VDD2.n35 VSUBS 0.011713f
C65 VDD2.n36 VSUBS 0.011062f
C66 VDD2.n37 VSUBS 0.020586f
C67 VDD2.n38 VSUBS 0.020586f
C68 VDD2.n39 VSUBS 0.011062f
C69 VDD2.n40 VSUBS 0.011713f
C70 VDD2.n41 VSUBS 0.026147f
C71 VDD2.n42 VSUBS 0.066275f
C72 VDD2.n43 VSUBS 0.011713f
C73 VDD2.n44 VSUBS 0.011062f
C74 VDD2.n45 VSUBS 0.046178f
C75 VDD2.n46 VSUBS 0.522394f
C76 VDD2.n47 VSUBS 0.023494f
C77 VDD2.n48 VSUBS 0.020586f
C78 VDD2.n49 VSUBS 0.011062f
C79 VDD2.n50 VSUBS 0.026147f
C80 VDD2.n51 VSUBS 0.011713f
C81 VDD2.n52 VSUBS 0.020586f
C82 VDD2.n53 VSUBS 0.011062f
C83 VDD2.n54 VSUBS 0.026147f
C84 VDD2.n55 VSUBS 0.011713f
C85 VDD2.n56 VSUBS 0.020586f
C86 VDD2.n57 VSUBS 0.011062f
C87 VDD2.n58 VSUBS 0.026147f
C88 VDD2.n59 VSUBS 0.011713f
C89 VDD2.n60 VSUBS 0.737678f
C90 VDD2.n61 VSUBS 0.011062f
C91 VDD2.t1 VSUBS 0.055747f
C92 VDD2.n62 VSUBS 0.107737f
C93 VDD2.n63 VSUBS 0.016633f
C94 VDD2.n64 VSUBS 0.01961f
C95 VDD2.n65 VSUBS 0.026147f
C96 VDD2.n66 VSUBS 0.011713f
C97 VDD2.n67 VSUBS 0.011062f
C98 VDD2.n68 VSUBS 0.020586f
C99 VDD2.n69 VSUBS 0.020586f
C100 VDD2.n70 VSUBS 0.011062f
C101 VDD2.n71 VSUBS 0.011713f
C102 VDD2.n72 VSUBS 0.026147f
C103 VDD2.n73 VSUBS 0.026147f
C104 VDD2.n74 VSUBS 0.011713f
C105 VDD2.n75 VSUBS 0.011062f
C106 VDD2.n76 VSUBS 0.020586f
C107 VDD2.n77 VSUBS 0.020586f
C108 VDD2.n78 VSUBS 0.011062f
C109 VDD2.n79 VSUBS 0.011713f
C110 VDD2.n80 VSUBS 0.026147f
C111 VDD2.n81 VSUBS 0.026147f
C112 VDD2.n82 VSUBS 0.011713f
C113 VDD2.n83 VSUBS 0.011062f
C114 VDD2.n84 VSUBS 0.020586f
C115 VDD2.n85 VSUBS 0.020586f
C116 VDD2.n86 VSUBS 0.011062f
C117 VDD2.n87 VSUBS 0.011713f
C118 VDD2.n88 VSUBS 0.026147f
C119 VDD2.n89 VSUBS 0.066275f
C120 VDD2.n90 VSUBS 0.011713f
C121 VDD2.n91 VSUBS 0.011062f
C122 VDD2.n92 VSUBS 0.046178f
C123 VDD2.n93 VSUBS 0.047644f
C124 VDD2.n94 VSUBS 2.23434f
C125 VN.t1 VSUBS 2.61229f
C126 VN.t0 VSUBS 3.17511f
C127 B.n0 VSUBS 0.005949f
C128 B.n1 VSUBS 0.005949f
C129 B.n2 VSUBS 0.008798f
C130 B.n3 VSUBS 0.006742f
C131 B.n4 VSUBS 0.006742f
C132 B.n5 VSUBS 0.006742f
C133 B.n6 VSUBS 0.006742f
C134 B.n7 VSUBS 0.006742f
C135 B.n8 VSUBS 0.006742f
C136 B.n9 VSUBS 0.006742f
C137 B.n10 VSUBS 0.006742f
C138 B.n11 VSUBS 0.006742f
C139 B.n12 VSUBS 0.006742f
C140 B.n13 VSUBS 0.006742f
C141 B.n14 VSUBS 0.015237f
C142 B.n15 VSUBS 0.006742f
C143 B.n16 VSUBS 0.006742f
C144 B.n17 VSUBS 0.006742f
C145 B.n18 VSUBS 0.006742f
C146 B.n19 VSUBS 0.006742f
C147 B.n20 VSUBS 0.006742f
C148 B.n21 VSUBS 0.006742f
C149 B.n22 VSUBS 0.006742f
C150 B.n23 VSUBS 0.006742f
C151 B.n24 VSUBS 0.006742f
C152 B.n25 VSUBS 0.006742f
C153 B.n26 VSUBS 0.006742f
C154 B.n27 VSUBS 0.006742f
C155 B.n28 VSUBS 0.006742f
C156 B.n29 VSUBS 0.006742f
C157 B.n30 VSUBS 0.006346f
C158 B.n31 VSUBS 0.006742f
C159 B.t1 VSUBS 0.138232f
C160 B.t2 VSUBS 0.166609f
C161 B.t0 VSUBS 1.02549f
C162 B.n32 VSUBS 0.272763f
C163 B.n33 VSUBS 0.197196f
C164 B.n34 VSUBS 0.015621f
C165 B.n35 VSUBS 0.006742f
C166 B.n36 VSUBS 0.006742f
C167 B.n37 VSUBS 0.006742f
C168 B.n38 VSUBS 0.006742f
C169 B.t10 VSUBS 0.138234f
C170 B.t11 VSUBS 0.166611f
C171 B.t9 VSUBS 1.02549f
C172 B.n39 VSUBS 0.272761f
C173 B.n40 VSUBS 0.197194f
C174 B.n41 VSUBS 0.006742f
C175 B.n42 VSUBS 0.006742f
C176 B.n43 VSUBS 0.006742f
C177 B.n44 VSUBS 0.006742f
C178 B.n45 VSUBS 0.006742f
C179 B.n46 VSUBS 0.006742f
C180 B.n47 VSUBS 0.006742f
C181 B.n48 VSUBS 0.006742f
C182 B.n49 VSUBS 0.006742f
C183 B.n50 VSUBS 0.006742f
C184 B.n51 VSUBS 0.006742f
C185 B.n52 VSUBS 0.006742f
C186 B.n53 VSUBS 0.006742f
C187 B.n54 VSUBS 0.006742f
C188 B.n55 VSUBS 0.006742f
C189 B.n56 VSUBS 0.015698f
C190 B.n57 VSUBS 0.006742f
C191 B.n58 VSUBS 0.006742f
C192 B.n59 VSUBS 0.006742f
C193 B.n60 VSUBS 0.006742f
C194 B.n61 VSUBS 0.006742f
C195 B.n62 VSUBS 0.006742f
C196 B.n63 VSUBS 0.006742f
C197 B.n64 VSUBS 0.006742f
C198 B.n65 VSUBS 0.006742f
C199 B.n66 VSUBS 0.006742f
C200 B.n67 VSUBS 0.006742f
C201 B.n68 VSUBS 0.006742f
C202 B.n69 VSUBS 0.006742f
C203 B.n70 VSUBS 0.006742f
C204 B.n71 VSUBS 0.006742f
C205 B.n72 VSUBS 0.006742f
C206 B.n73 VSUBS 0.006742f
C207 B.n74 VSUBS 0.006742f
C208 B.n75 VSUBS 0.006742f
C209 B.n76 VSUBS 0.006742f
C210 B.n77 VSUBS 0.006742f
C211 B.n78 VSUBS 0.006742f
C212 B.n79 VSUBS 0.006742f
C213 B.n80 VSUBS 0.006742f
C214 B.n81 VSUBS 0.006742f
C215 B.n82 VSUBS 0.015237f
C216 B.n83 VSUBS 0.006742f
C217 B.n84 VSUBS 0.006742f
C218 B.n85 VSUBS 0.006742f
C219 B.n86 VSUBS 0.006742f
C220 B.n87 VSUBS 0.006742f
C221 B.n88 VSUBS 0.006742f
C222 B.n89 VSUBS 0.006742f
C223 B.n90 VSUBS 0.006742f
C224 B.n91 VSUBS 0.006742f
C225 B.n92 VSUBS 0.006742f
C226 B.n93 VSUBS 0.006742f
C227 B.n94 VSUBS 0.006742f
C228 B.n95 VSUBS 0.006742f
C229 B.n96 VSUBS 0.006742f
C230 B.n97 VSUBS 0.006742f
C231 B.n98 VSUBS 0.006742f
C232 B.t8 VSUBS 0.138234f
C233 B.t7 VSUBS 0.166611f
C234 B.t6 VSUBS 1.02549f
C235 B.n99 VSUBS 0.272761f
C236 B.n100 VSUBS 0.197194f
C237 B.n101 VSUBS 0.006742f
C238 B.n102 VSUBS 0.006742f
C239 B.n103 VSUBS 0.006742f
C240 B.n104 VSUBS 0.006742f
C241 B.n105 VSUBS 0.003768f
C242 B.n106 VSUBS 0.006742f
C243 B.n107 VSUBS 0.006742f
C244 B.n108 VSUBS 0.006742f
C245 B.n109 VSUBS 0.006742f
C246 B.n110 VSUBS 0.006742f
C247 B.n111 VSUBS 0.006742f
C248 B.n112 VSUBS 0.006742f
C249 B.n113 VSUBS 0.006742f
C250 B.n114 VSUBS 0.006742f
C251 B.n115 VSUBS 0.006742f
C252 B.n116 VSUBS 0.006742f
C253 B.n117 VSUBS 0.006742f
C254 B.n118 VSUBS 0.006742f
C255 B.n119 VSUBS 0.006742f
C256 B.n120 VSUBS 0.006742f
C257 B.n121 VSUBS 0.015698f
C258 B.n122 VSUBS 0.006742f
C259 B.n123 VSUBS 0.006742f
C260 B.n124 VSUBS 0.006742f
C261 B.n125 VSUBS 0.006742f
C262 B.n126 VSUBS 0.006742f
C263 B.n127 VSUBS 0.006742f
C264 B.n128 VSUBS 0.006742f
C265 B.n129 VSUBS 0.006742f
C266 B.n130 VSUBS 0.006742f
C267 B.n131 VSUBS 0.006742f
C268 B.n132 VSUBS 0.006742f
C269 B.n133 VSUBS 0.006742f
C270 B.n134 VSUBS 0.006742f
C271 B.n135 VSUBS 0.006742f
C272 B.n136 VSUBS 0.006742f
C273 B.n137 VSUBS 0.006742f
C274 B.n138 VSUBS 0.006742f
C275 B.n139 VSUBS 0.006742f
C276 B.n140 VSUBS 0.006742f
C277 B.n141 VSUBS 0.006742f
C278 B.n142 VSUBS 0.006742f
C279 B.n143 VSUBS 0.006742f
C280 B.n144 VSUBS 0.006742f
C281 B.n145 VSUBS 0.006742f
C282 B.n146 VSUBS 0.006742f
C283 B.n147 VSUBS 0.006742f
C284 B.n148 VSUBS 0.006742f
C285 B.n149 VSUBS 0.006742f
C286 B.n150 VSUBS 0.006742f
C287 B.n151 VSUBS 0.006742f
C288 B.n152 VSUBS 0.006742f
C289 B.n153 VSUBS 0.006742f
C290 B.n154 VSUBS 0.006742f
C291 B.n155 VSUBS 0.006742f
C292 B.n156 VSUBS 0.006742f
C293 B.n157 VSUBS 0.006742f
C294 B.n158 VSUBS 0.006742f
C295 B.n159 VSUBS 0.006742f
C296 B.n160 VSUBS 0.006742f
C297 B.n161 VSUBS 0.006742f
C298 B.n162 VSUBS 0.006742f
C299 B.n163 VSUBS 0.006742f
C300 B.n164 VSUBS 0.006742f
C301 B.n165 VSUBS 0.006742f
C302 B.n166 VSUBS 0.006742f
C303 B.n167 VSUBS 0.006742f
C304 B.n168 VSUBS 0.015237f
C305 B.n169 VSUBS 0.015237f
C306 B.n170 VSUBS 0.015698f
C307 B.n171 VSUBS 0.006742f
C308 B.n172 VSUBS 0.006742f
C309 B.n173 VSUBS 0.006742f
C310 B.n174 VSUBS 0.006742f
C311 B.n175 VSUBS 0.006742f
C312 B.n176 VSUBS 0.006742f
C313 B.n177 VSUBS 0.006742f
C314 B.n178 VSUBS 0.006742f
C315 B.n179 VSUBS 0.006742f
C316 B.n180 VSUBS 0.006742f
C317 B.n181 VSUBS 0.006742f
C318 B.n182 VSUBS 0.006742f
C319 B.n183 VSUBS 0.006742f
C320 B.n184 VSUBS 0.006742f
C321 B.n185 VSUBS 0.006742f
C322 B.n186 VSUBS 0.006742f
C323 B.n187 VSUBS 0.006742f
C324 B.n188 VSUBS 0.006742f
C325 B.n189 VSUBS 0.006742f
C326 B.n190 VSUBS 0.006742f
C327 B.n191 VSUBS 0.006742f
C328 B.n192 VSUBS 0.006742f
C329 B.n193 VSUBS 0.006742f
C330 B.n194 VSUBS 0.006742f
C331 B.n195 VSUBS 0.006742f
C332 B.n196 VSUBS 0.006742f
C333 B.n197 VSUBS 0.006742f
C334 B.n198 VSUBS 0.006742f
C335 B.n199 VSUBS 0.006742f
C336 B.n200 VSUBS 0.006742f
C337 B.n201 VSUBS 0.006742f
C338 B.n202 VSUBS 0.006742f
C339 B.n203 VSUBS 0.006742f
C340 B.n204 VSUBS 0.006742f
C341 B.n205 VSUBS 0.006742f
C342 B.n206 VSUBS 0.006742f
C343 B.n207 VSUBS 0.006742f
C344 B.n208 VSUBS 0.006742f
C345 B.n209 VSUBS 0.006742f
C346 B.n210 VSUBS 0.006742f
C347 B.n211 VSUBS 0.006742f
C348 B.n212 VSUBS 0.006742f
C349 B.n213 VSUBS 0.006742f
C350 B.n214 VSUBS 0.006742f
C351 B.n215 VSUBS 0.006742f
C352 B.t5 VSUBS 0.138232f
C353 B.t4 VSUBS 0.166609f
C354 B.t3 VSUBS 1.02549f
C355 B.n216 VSUBS 0.272763f
C356 B.n217 VSUBS 0.197196f
C357 B.n218 VSUBS 0.015621f
C358 B.n219 VSUBS 0.006346f
C359 B.n220 VSUBS 0.006742f
C360 B.n221 VSUBS 0.006742f
C361 B.n222 VSUBS 0.006742f
C362 B.n223 VSUBS 0.006742f
C363 B.n224 VSUBS 0.006742f
C364 B.n225 VSUBS 0.006742f
C365 B.n226 VSUBS 0.006742f
C366 B.n227 VSUBS 0.006742f
C367 B.n228 VSUBS 0.006742f
C368 B.n229 VSUBS 0.006742f
C369 B.n230 VSUBS 0.006742f
C370 B.n231 VSUBS 0.006742f
C371 B.n232 VSUBS 0.006742f
C372 B.n233 VSUBS 0.006742f
C373 B.n234 VSUBS 0.006742f
C374 B.n235 VSUBS 0.003768f
C375 B.n236 VSUBS 0.015621f
C376 B.n237 VSUBS 0.006346f
C377 B.n238 VSUBS 0.006742f
C378 B.n239 VSUBS 0.006742f
C379 B.n240 VSUBS 0.006742f
C380 B.n241 VSUBS 0.006742f
C381 B.n242 VSUBS 0.006742f
C382 B.n243 VSUBS 0.006742f
C383 B.n244 VSUBS 0.006742f
C384 B.n245 VSUBS 0.006742f
C385 B.n246 VSUBS 0.006742f
C386 B.n247 VSUBS 0.006742f
C387 B.n248 VSUBS 0.006742f
C388 B.n249 VSUBS 0.006742f
C389 B.n250 VSUBS 0.006742f
C390 B.n251 VSUBS 0.006742f
C391 B.n252 VSUBS 0.006742f
C392 B.n253 VSUBS 0.006742f
C393 B.n254 VSUBS 0.006742f
C394 B.n255 VSUBS 0.006742f
C395 B.n256 VSUBS 0.006742f
C396 B.n257 VSUBS 0.006742f
C397 B.n258 VSUBS 0.006742f
C398 B.n259 VSUBS 0.006742f
C399 B.n260 VSUBS 0.006742f
C400 B.n261 VSUBS 0.006742f
C401 B.n262 VSUBS 0.006742f
C402 B.n263 VSUBS 0.006742f
C403 B.n264 VSUBS 0.006742f
C404 B.n265 VSUBS 0.006742f
C405 B.n266 VSUBS 0.006742f
C406 B.n267 VSUBS 0.006742f
C407 B.n268 VSUBS 0.006742f
C408 B.n269 VSUBS 0.006742f
C409 B.n270 VSUBS 0.006742f
C410 B.n271 VSUBS 0.006742f
C411 B.n272 VSUBS 0.006742f
C412 B.n273 VSUBS 0.006742f
C413 B.n274 VSUBS 0.006742f
C414 B.n275 VSUBS 0.006742f
C415 B.n276 VSUBS 0.006742f
C416 B.n277 VSUBS 0.006742f
C417 B.n278 VSUBS 0.006742f
C418 B.n279 VSUBS 0.006742f
C419 B.n280 VSUBS 0.006742f
C420 B.n281 VSUBS 0.006742f
C421 B.n282 VSUBS 0.006742f
C422 B.n283 VSUBS 0.015698f
C423 B.n284 VSUBS 0.014877f
C424 B.n285 VSUBS 0.016058f
C425 B.n286 VSUBS 0.006742f
C426 B.n287 VSUBS 0.006742f
C427 B.n288 VSUBS 0.006742f
C428 B.n289 VSUBS 0.006742f
C429 B.n290 VSUBS 0.006742f
C430 B.n291 VSUBS 0.006742f
C431 B.n292 VSUBS 0.006742f
C432 B.n293 VSUBS 0.006742f
C433 B.n294 VSUBS 0.006742f
C434 B.n295 VSUBS 0.006742f
C435 B.n296 VSUBS 0.006742f
C436 B.n297 VSUBS 0.006742f
C437 B.n298 VSUBS 0.006742f
C438 B.n299 VSUBS 0.006742f
C439 B.n300 VSUBS 0.006742f
C440 B.n301 VSUBS 0.006742f
C441 B.n302 VSUBS 0.006742f
C442 B.n303 VSUBS 0.006742f
C443 B.n304 VSUBS 0.006742f
C444 B.n305 VSUBS 0.006742f
C445 B.n306 VSUBS 0.006742f
C446 B.n307 VSUBS 0.006742f
C447 B.n308 VSUBS 0.006742f
C448 B.n309 VSUBS 0.006742f
C449 B.n310 VSUBS 0.006742f
C450 B.n311 VSUBS 0.006742f
C451 B.n312 VSUBS 0.006742f
C452 B.n313 VSUBS 0.006742f
C453 B.n314 VSUBS 0.006742f
C454 B.n315 VSUBS 0.006742f
C455 B.n316 VSUBS 0.006742f
C456 B.n317 VSUBS 0.006742f
C457 B.n318 VSUBS 0.006742f
C458 B.n319 VSUBS 0.006742f
C459 B.n320 VSUBS 0.006742f
C460 B.n321 VSUBS 0.006742f
C461 B.n322 VSUBS 0.006742f
C462 B.n323 VSUBS 0.006742f
C463 B.n324 VSUBS 0.006742f
C464 B.n325 VSUBS 0.006742f
C465 B.n326 VSUBS 0.006742f
C466 B.n327 VSUBS 0.006742f
C467 B.n328 VSUBS 0.006742f
C468 B.n329 VSUBS 0.006742f
C469 B.n330 VSUBS 0.006742f
C470 B.n331 VSUBS 0.006742f
C471 B.n332 VSUBS 0.006742f
C472 B.n333 VSUBS 0.006742f
C473 B.n334 VSUBS 0.006742f
C474 B.n335 VSUBS 0.006742f
C475 B.n336 VSUBS 0.006742f
C476 B.n337 VSUBS 0.006742f
C477 B.n338 VSUBS 0.006742f
C478 B.n339 VSUBS 0.006742f
C479 B.n340 VSUBS 0.006742f
C480 B.n341 VSUBS 0.006742f
C481 B.n342 VSUBS 0.006742f
C482 B.n343 VSUBS 0.006742f
C483 B.n344 VSUBS 0.006742f
C484 B.n345 VSUBS 0.006742f
C485 B.n346 VSUBS 0.006742f
C486 B.n347 VSUBS 0.006742f
C487 B.n348 VSUBS 0.006742f
C488 B.n349 VSUBS 0.006742f
C489 B.n350 VSUBS 0.006742f
C490 B.n351 VSUBS 0.006742f
C491 B.n352 VSUBS 0.006742f
C492 B.n353 VSUBS 0.006742f
C493 B.n354 VSUBS 0.006742f
C494 B.n355 VSUBS 0.006742f
C495 B.n356 VSUBS 0.006742f
C496 B.n357 VSUBS 0.006742f
C497 B.n358 VSUBS 0.006742f
C498 B.n359 VSUBS 0.006742f
C499 B.n360 VSUBS 0.006742f
C500 B.n361 VSUBS 0.015237f
C501 B.n362 VSUBS 0.015237f
C502 B.n363 VSUBS 0.015698f
C503 B.n364 VSUBS 0.006742f
C504 B.n365 VSUBS 0.006742f
C505 B.n366 VSUBS 0.006742f
C506 B.n367 VSUBS 0.006742f
C507 B.n368 VSUBS 0.006742f
C508 B.n369 VSUBS 0.006742f
C509 B.n370 VSUBS 0.006742f
C510 B.n371 VSUBS 0.006742f
C511 B.n372 VSUBS 0.006742f
C512 B.n373 VSUBS 0.006742f
C513 B.n374 VSUBS 0.006742f
C514 B.n375 VSUBS 0.006742f
C515 B.n376 VSUBS 0.006742f
C516 B.n377 VSUBS 0.006742f
C517 B.n378 VSUBS 0.006742f
C518 B.n379 VSUBS 0.006742f
C519 B.n380 VSUBS 0.006742f
C520 B.n381 VSUBS 0.006742f
C521 B.n382 VSUBS 0.006742f
C522 B.n383 VSUBS 0.006742f
C523 B.n384 VSUBS 0.006742f
C524 B.n385 VSUBS 0.006742f
C525 B.n386 VSUBS 0.006742f
C526 B.n387 VSUBS 0.006742f
C527 B.n388 VSUBS 0.006742f
C528 B.n389 VSUBS 0.006742f
C529 B.n390 VSUBS 0.006742f
C530 B.n391 VSUBS 0.006742f
C531 B.n392 VSUBS 0.006742f
C532 B.n393 VSUBS 0.006742f
C533 B.n394 VSUBS 0.006742f
C534 B.n395 VSUBS 0.006742f
C535 B.n396 VSUBS 0.006742f
C536 B.n397 VSUBS 0.006742f
C537 B.n398 VSUBS 0.006742f
C538 B.n399 VSUBS 0.006742f
C539 B.n400 VSUBS 0.006742f
C540 B.n401 VSUBS 0.006742f
C541 B.n402 VSUBS 0.006742f
C542 B.n403 VSUBS 0.006742f
C543 B.n404 VSUBS 0.006742f
C544 B.n405 VSUBS 0.006742f
C545 B.n406 VSUBS 0.006742f
C546 B.n407 VSUBS 0.006742f
C547 B.n408 VSUBS 0.006742f
C548 B.n409 VSUBS 0.006742f
C549 B.n410 VSUBS 0.006346f
C550 B.n411 VSUBS 0.015621f
C551 B.n412 VSUBS 0.003768f
C552 B.n413 VSUBS 0.006742f
C553 B.n414 VSUBS 0.006742f
C554 B.n415 VSUBS 0.006742f
C555 B.n416 VSUBS 0.006742f
C556 B.n417 VSUBS 0.006742f
C557 B.n418 VSUBS 0.006742f
C558 B.n419 VSUBS 0.006742f
C559 B.n420 VSUBS 0.006742f
C560 B.n421 VSUBS 0.006742f
C561 B.n422 VSUBS 0.006742f
C562 B.n423 VSUBS 0.006742f
C563 B.n424 VSUBS 0.006742f
C564 B.n425 VSUBS 0.003768f
C565 B.n426 VSUBS 0.006742f
C566 B.n427 VSUBS 0.006742f
C567 B.n428 VSUBS 0.006742f
C568 B.n429 VSUBS 0.006742f
C569 B.n430 VSUBS 0.006742f
C570 B.n431 VSUBS 0.006742f
C571 B.n432 VSUBS 0.006742f
C572 B.n433 VSUBS 0.006742f
C573 B.n434 VSUBS 0.006742f
C574 B.n435 VSUBS 0.006742f
C575 B.n436 VSUBS 0.006742f
C576 B.n437 VSUBS 0.006742f
C577 B.n438 VSUBS 0.006742f
C578 B.n439 VSUBS 0.006742f
C579 B.n440 VSUBS 0.006742f
C580 B.n441 VSUBS 0.006742f
C581 B.n442 VSUBS 0.006742f
C582 B.n443 VSUBS 0.006742f
C583 B.n444 VSUBS 0.006742f
C584 B.n445 VSUBS 0.006742f
C585 B.n446 VSUBS 0.006742f
C586 B.n447 VSUBS 0.006742f
C587 B.n448 VSUBS 0.006742f
C588 B.n449 VSUBS 0.006742f
C589 B.n450 VSUBS 0.006742f
C590 B.n451 VSUBS 0.006742f
C591 B.n452 VSUBS 0.006742f
C592 B.n453 VSUBS 0.006742f
C593 B.n454 VSUBS 0.006742f
C594 B.n455 VSUBS 0.006742f
C595 B.n456 VSUBS 0.006742f
C596 B.n457 VSUBS 0.006742f
C597 B.n458 VSUBS 0.006742f
C598 B.n459 VSUBS 0.006742f
C599 B.n460 VSUBS 0.006742f
C600 B.n461 VSUBS 0.006742f
C601 B.n462 VSUBS 0.006742f
C602 B.n463 VSUBS 0.006742f
C603 B.n464 VSUBS 0.006742f
C604 B.n465 VSUBS 0.006742f
C605 B.n466 VSUBS 0.006742f
C606 B.n467 VSUBS 0.006742f
C607 B.n468 VSUBS 0.006742f
C608 B.n469 VSUBS 0.006742f
C609 B.n470 VSUBS 0.006742f
C610 B.n471 VSUBS 0.006742f
C611 B.n472 VSUBS 0.006742f
C612 B.n473 VSUBS 0.015698f
C613 B.n474 VSUBS 0.015698f
C614 B.n475 VSUBS 0.015237f
C615 B.n476 VSUBS 0.006742f
C616 B.n477 VSUBS 0.006742f
C617 B.n478 VSUBS 0.006742f
C618 B.n479 VSUBS 0.006742f
C619 B.n480 VSUBS 0.006742f
C620 B.n481 VSUBS 0.006742f
C621 B.n482 VSUBS 0.006742f
C622 B.n483 VSUBS 0.006742f
C623 B.n484 VSUBS 0.006742f
C624 B.n485 VSUBS 0.006742f
C625 B.n486 VSUBS 0.006742f
C626 B.n487 VSUBS 0.006742f
C627 B.n488 VSUBS 0.006742f
C628 B.n489 VSUBS 0.006742f
C629 B.n490 VSUBS 0.006742f
C630 B.n491 VSUBS 0.006742f
C631 B.n492 VSUBS 0.006742f
C632 B.n493 VSUBS 0.006742f
C633 B.n494 VSUBS 0.006742f
C634 B.n495 VSUBS 0.006742f
C635 B.n496 VSUBS 0.006742f
C636 B.n497 VSUBS 0.006742f
C637 B.n498 VSUBS 0.006742f
C638 B.n499 VSUBS 0.006742f
C639 B.n500 VSUBS 0.006742f
C640 B.n501 VSUBS 0.006742f
C641 B.n502 VSUBS 0.006742f
C642 B.n503 VSUBS 0.006742f
C643 B.n504 VSUBS 0.006742f
C644 B.n505 VSUBS 0.006742f
C645 B.n506 VSUBS 0.006742f
C646 B.n507 VSUBS 0.006742f
C647 B.n508 VSUBS 0.006742f
C648 B.n509 VSUBS 0.006742f
C649 B.n510 VSUBS 0.006742f
C650 B.n511 VSUBS 0.008798f
C651 B.n512 VSUBS 0.009373f
C652 B.n513 VSUBS 0.018638f
C653 VDD1.n0 VSUBS 0.023581f
C654 VDD1.n1 VSUBS 0.020662f
C655 VDD1.n2 VSUBS 0.011103f
C656 VDD1.n3 VSUBS 0.026244f
C657 VDD1.n4 VSUBS 0.011756f
C658 VDD1.n5 VSUBS 0.020662f
C659 VDD1.n6 VSUBS 0.011103f
C660 VDD1.n7 VSUBS 0.026244f
C661 VDD1.n8 VSUBS 0.011756f
C662 VDD1.n9 VSUBS 0.020662f
C663 VDD1.n10 VSUBS 0.011103f
C664 VDD1.n11 VSUBS 0.026244f
C665 VDD1.n12 VSUBS 0.011756f
C666 VDD1.n13 VSUBS 0.740408f
C667 VDD1.n14 VSUBS 0.011103f
C668 VDD1.t0 VSUBS 0.055953f
C669 VDD1.n15 VSUBS 0.108136f
C670 VDD1.n16 VSUBS 0.016695f
C671 VDD1.n17 VSUBS 0.019683f
C672 VDD1.n18 VSUBS 0.026244f
C673 VDD1.n19 VSUBS 0.011756f
C674 VDD1.n20 VSUBS 0.011103f
C675 VDD1.n21 VSUBS 0.020662f
C676 VDD1.n22 VSUBS 0.020662f
C677 VDD1.n23 VSUBS 0.011103f
C678 VDD1.n24 VSUBS 0.011756f
C679 VDD1.n25 VSUBS 0.026244f
C680 VDD1.n26 VSUBS 0.026244f
C681 VDD1.n27 VSUBS 0.011756f
C682 VDD1.n28 VSUBS 0.011103f
C683 VDD1.n29 VSUBS 0.020662f
C684 VDD1.n30 VSUBS 0.020662f
C685 VDD1.n31 VSUBS 0.011103f
C686 VDD1.n32 VSUBS 0.011756f
C687 VDD1.n33 VSUBS 0.026244f
C688 VDD1.n34 VSUBS 0.026244f
C689 VDD1.n35 VSUBS 0.011756f
C690 VDD1.n36 VSUBS 0.011103f
C691 VDD1.n37 VSUBS 0.020662f
C692 VDD1.n38 VSUBS 0.020662f
C693 VDD1.n39 VSUBS 0.011103f
C694 VDD1.n40 VSUBS 0.011756f
C695 VDD1.n41 VSUBS 0.026244f
C696 VDD1.n42 VSUBS 0.066521f
C697 VDD1.n43 VSUBS 0.011756f
C698 VDD1.n44 VSUBS 0.011103f
C699 VDD1.n45 VSUBS 0.046349f
C700 VDD1.n46 VSUBS 0.049025f
C701 VDD1.n47 VSUBS 0.023581f
C702 VDD1.n48 VSUBS 0.020662f
C703 VDD1.n49 VSUBS 0.011103f
C704 VDD1.n50 VSUBS 0.026244f
C705 VDD1.n51 VSUBS 0.011756f
C706 VDD1.n52 VSUBS 0.020662f
C707 VDD1.n53 VSUBS 0.011103f
C708 VDD1.n54 VSUBS 0.026244f
C709 VDD1.n55 VSUBS 0.011756f
C710 VDD1.n56 VSUBS 0.020662f
C711 VDD1.n57 VSUBS 0.011103f
C712 VDD1.n58 VSUBS 0.026244f
C713 VDD1.n59 VSUBS 0.011756f
C714 VDD1.n60 VSUBS 0.740408f
C715 VDD1.n61 VSUBS 0.011103f
C716 VDD1.t1 VSUBS 0.055953f
C717 VDD1.n62 VSUBS 0.108136f
C718 VDD1.n63 VSUBS 0.016695f
C719 VDD1.n64 VSUBS 0.019683f
C720 VDD1.n65 VSUBS 0.026244f
C721 VDD1.n66 VSUBS 0.011756f
C722 VDD1.n67 VSUBS 0.011103f
C723 VDD1.n68 VSUBS 0.020662f
C724 VDD1.n69 VSUBS 0.020662f
C725 VDD1.n70 VSUBS 0.011103f
C726 VDD1.n71 VSUBS 0.011756f
C727 VDD1.n72 VSUBS 0.026244f
C728 VDD1.n73 VSUBS 0.026244f
C729 VDD1.n74 VSUBS 0.011756f
C730 VDD1.n75 VSUBS 0.011103f
C731 VDD1.n76 VSUBS 0.020662f
C732 VDD1.n77 VSUBS 0.020662f
C733 VDD1.n78 VSUBS 0.011103f
C734 VDD1.n79 VSUBS 0.011756f
C735 VDD1.n80 VSUBS 0.026244f
C736 VDD1.n81 VSUBS 0.026244f
C737 VDD1.n82 VSUBS 0.011756f
C738 VDD1.n83 VSUBS 0.011103f
C739 VDD1.n84 VSUBS 0.020662f
C740 VDD1.n85 VSUBS 0.020662f
C741 VDD1.n86 VSUBS 0.011103f
C742 VDD1.n87 VSUBS 0.011756f
C743 VDD1.n88 VSUBS 0.026244f
C744 VDD1.n89 VSUBS 0.066521f
C745 VDD1.n90 VSUBS 0.011756f
C746 VDD1.n91 VSUBS 0.011103f
C747 VDD1.n92 VSUBS 0.046349f
C748 VDD1.n93 VSUBS 0.562887f
C749 VTAIL.n0 VSUBS 0.027427f
C750 VTAIL.n1 VSUBS 0.024033f
C751 VTAIL.n2 VSUBS 0.012914f
C752 VTAIL.n3 VSUBS 0.030525f
C753 VTAIL.n4 VSUBS 0.013674f
C754 VTAIL.n5 VSUBS 0.024033f
C755 VTAIL.n6 VSUBS 0.012914f
C756 VTAIL.n7 VSUBS 0.030525f
C757 VTAIL.n8 VSUBS 0.013674f
C758 VTAIL.n9 VSUBS 0.024033f
C759 VTAIL.n10 VSUBS 0.012914f
C760 VTAIL.n11 VSUBS 0.030525f
C761 VTAIL.n12 VSUBS 0.013674f
C762 VTAIL.n13 VSUBS 0.861182f
C763 VTAIL.n14 VSUBS 0.012914f
C764 VTAIL.t3 VSUBS 0.06508f
C765 VTAIL.n15 VSUBS 0.125775f
C766 VTAIL.n16 VSUBS 0.019418f
C767 VTAIL.n17 VSUBS 0.022893f
C768 VTAIL.n18 VSUBS 0.030525f
C769 VTAIL.n19 VSUBS 0.013674f
C770 VTAIL.n20 VSUBS 0.012914f
C771 VTAIL.n21 VSUBS 0.024033f
C772 VTAIL.n22 VSUBS 0.024033f
C773 VTAIL.n23 VSUBS 0.012914f
C774 VTAIL.n24 VSUBS 0.013674f
C775 VTAIL.n25 VSUBS 0.030525f
C776 VTAIL.n26 VSUBS 0.030525f
C777 VTAIL.n27 VSUBS 0.013674f
C778 VTAIL.n28 VSUBS 0.012914f
C779 VTAIL.n29 VSUBS 0.024033f
C780 VTAIL.n30 VSUBS 0.024033f
C781 VTAIL.n31 VSUBS 0.012914f
C782 VTAIL.n32 VSUBS 0.013674f
C783 VTAIL.n33 VSUBS 0.030525f
C784 VTAIL.n34 VSUBS 0.030525f
C785 VTAIL.n35 VSUBS 0.013674f
C786 VTAIL.n36 VSUBS 0.012914f
C787 VTAIL.n37 VSUBS 0.024033f
C788 VTAIL.n38 VSUBS 0.024033f
C789 VTAIL.n39 VSUBS 0.012914f
C790 VTAIL.n40 VSUBS 0.013674f
C791 VTAIL.n41 VSUBS 0.030525f
C792 VTAIL.n42 VSUBS 0.077371f
C793 VTAIL.n43 VSUBS 0.013674f
C794 VTAIL.n44 VSUBS 0.012914f
C795 VTAIL.n45 VSUBS 0.053909f
C796 VTAIL.n46 VSUBS 0.039013f
C797 VTAIL.n47 VSUBS 1.41652f
C798 VTAIL.n48 VSUBS 0.027427f
C799 VTAIL.n49 VSUBS 0.024033f
C800 VTAIL.n50 VSUBS 0.012914f
C801 VTAIL.n51 VSUBS 0.030525f
C802 VTAIL.n52 VSUBS 0.013674f
C803 VTAIL.n53 VSUBS 0.024033f
C804 VTAIL.n54 VSUBS 0.012914f
C805 VTAIL.n55 VSUBS 0.030525f
C806 VTAIL.n56 VSUBS 0.013674f
C807 VTAIL.n57 VSUBS 0.024033f
C808 VTAIL.n58 VSUBS 0.012914f
C809 VTAIL.n59 VSUBS 0.030525f
C810 VTAIL.n60 VSUBS 0.013674f
C811 VTAIL.n61 VSUBS 0.861182f
C812 VTAIL.n62 VSUBS 0.012914f
C813 VTAIL.t0 VSUBS 0.06508f
C814 VTAIL.n63 VSUBS 0.125775f
C815 VTAIL.n64 VSUBS 0.019418f
C816 VTAIL.n65 VSUBS 0.022893f
C817 VTAIL.n66 VSUBS 0.030525f
C818 VTAIL.n67 VSUBS 0.013674f
C819 VTAIL.n68 VSUBS 0.012914f
C820 VTAIL.n69 VSUBS 0.024033f
C821 VTAIL.n70 VSUBS 0.024033f
C822 VTAIL.n71 VSUBS 0.012914f
C823 VTAIL.n72 VSUBS 0.013674f
C824 VTAIL.n73 VSUBS 0.030525f
C825 VTAIL.n74 VSUBS 0.030525f
C826 VTAIL.n75 VSUBS 0.013674f
C827 VTAIL.n76 VSUBS 0.012914f
C828 VTAIL.n77 VSUBS 0.024033f
C829 VTAIL.n78 VSUBS 0.024033f
C830 VTAIL.n79 VSUBS 0.012914f
C831 VTAIL.n80 VSUBS 0.013674f
C832 VTAIL.n81 VSUBS 0.030525f
C833 VTAIL.n82 VSUBS 0.030525f
C834 VTAIL.n83 VSUBS 0.013674f
C835 VTAIL.n84 VSUBS 0.012914f
C836 VTAIL.n85 VSUBS 0.024033f
C837 VTAIL.n86 VSUBS 0.024033f
C838 VTAIL.n87 VSUBS 0.012914f
C839 VTAIL.n88 VSUBS 0.013674f
C840 VTAIL.n89 VSUBS 0.030525f
C841 VTAIL.n90 VSUBS 0.077371f
C842 VTAIL.n91 VSUBS 0.013674f
C843 VTAIL.n92 VSUBS 0.012914f
C844 VTAIL.n93 VSUBS 0.053909f
C845 VTAIL.n94 VSUBS 0.039013f
C846 VTAIL.n95 VSUBS 1.46092f
C847 VTAIL.n96 VSUBS 0.027427f
C848 VTAIL.n97 VSUBS 0.024033f
C849 VTAIL.n98 VSUBS 0.012914f
C850 VTAIL.n99 VSUBS 0.030525f
C851 VTAIL.n100 VSUBS 0.013674f
C852 VTAIL.n101 VSUBS 0.024033f
C853 VTAIL.n102 VSUBS 0.012914f
C854 VTAIL.n103 VSUBS 0.030525f
C855 VTAIL.n104 VSUBS 0.013674f
C856 VTAIL.n105 VSUBS 0.024033f
C857 VTAIL.n106 VSUBS 0.012914f
C858 VTAIL.n107 VSUBS 0.030525f
C859 VTAIL.n108 VSUBS 0.013674f
C860 VTAIL.n109 VSUBS 0.861182f
C861 VTAIL.n110 VSUBS 0.012914f
C862 VTAIL.t2 VSUBS 0.06508f
C863 VTAIL.n111 VSUBS 0.125775f
C864 VTAIL.n112 VSUBS 0.019418f
C865 VTAIL.n113 VSUBS 0.022893f
C866 VTAIL.n114 VSUBS 0.030525f
C867 VTAIL.n115 VSUBS 0.013674f
C868 VTAIL.n116 VSUBS 0.012914f
C869 VTAIL.n117 VSUBS 0.024033f
C870 VTAIL.n118 VSUBS 0.024033f
C871 VTAIL.n119 VSUBS 0.012914f
C872 VTAIL.n120 VSUBS 0.013674f
C873 VTAIL.n121 VSUBS 0.030525f
C874 VTAIL.n122 VSUBS 0.030525f
C875 VTAIL.n123 VSUBS 0.013674f
C876 VTAIL.n124 VSUBS 0.012914f
C877 VTAIL.n125 VSUBS 0.024033f
C878 VTAIL.n126 VSUBS 0.024033f
C879 VTAIL.n127 VSUBS 0.012914f
C880 VTAIL.n128 VSUBS 0.013674f
C881 VTAIL.n129 VSUBS 0.030525f
C882 VTAIL.n130 VSUBS 0.030525f
C883 VTAIL.n131 VSUBS 0.013674f
C884 VTAIL.n132 VSUBS 0.012914f
C885 VTAIL.n133 VSUBS 0.024033f
C886 VTAIL.n134 VSUBS 0.024033f
C887 VTAIL.n135 VSUBS 0.012914f
C888 VTAIL.n136 VSUBS 0.013674f
C889 VTAIL.n137 VSUBS 0.030525f
C890 VTAIL.n138 VSUBS 0.077371f
C891 VTAIL.n139 VSUBS 0.013674f
C892 VTAIL.n140 VSUBS 0.012914f
C893 VTAIL.n141 VSUBS 0.053909f
C894 VTAIL.n142 VSUBS 0.039013f
C895 VTAIL.n143 VSUBS 1.26532f
C896 VTAIL.n144 VSUBS 0.027427f
C897 VTAIL.n145 VSUBS 0.024033f
C898 VTAIL.n146 VSUBS 0.012914f
C899 VTAIL.n147 VSUBS 0.030525f
C900 VTAIL.n148 VSUBS 0.013674f
C901 VTAIL.n149 VSUBS 0.024033f
C902 VTAIL.n150 VSUBS 0.012914f
C903 VTAIL.n151 VSUBS 0.030525f
C904 VTAIL.n152 VSUBS 0.013674f
C905 VTAIL.n153 VSUBS 0.024033f
C906 VTAIL.n154 VSUBS 0.012914f
C907 VTAIL.n155 VSUBS 0.030525f
C908 VTAIL.n156 VSUBS 0.013674f
C909 VTAIL.n157 VSUBS 0.861182f
C910 VTAIL.n158 VSUBS 0.012914f
C911 VTAIL.t1 VSUBS 0.06508f
C912 VTAIL.n159 VSUBS 0.125775f
C913 VTAIL.n160 VSUBS 0.019418f
C914 VTAIL.n161 VSUBS 0.022893f
C915 VTAIL.n162 VSUBS 0.030525f
C916 VTAIL.n163 VSUBS 0.013674f
C917 VTAIL.n164 VSUBS 0.012914f
C918 VTAIL.n165 VSUBS 0.024033f
C919 VTAIL.n166 VSUBS 0.024033f
C920 VTAIL.n167 VSUBS 0.012914f
C921 VTAIL.n168 VSUBS 0.013674f
C922 VTAIL.n169 VSUBS 0.030525f
C923 VTAIL.n170 VSUBS 0.030525f
C924 VTAIL.n171 VSUBS 0.013674f
C925 VTAIL.n172 VSUBS 0.012914f
C926 VTAIL.n173 VSUBS 0.024033f
C927 VTAIL.n174 VSUBS 0.024033f
C928 VTAIL.n175 VSUBS 0.012914f
C929 VTAIL.n176 VSUBS 0.013674f
C930 VTAIL.n177 VSUBS 0.030525f
C931 VTAIL.n178 VSUBS 0.030525f
C932 VTAIL.n179 VSUBS 0.013674f
C933 VTAIL.n180 VSUBS 0.012914f
C934 VTAIL.n181 VSUBS 0.024033f
C935 VTAIL.n182 VSUBS 0.024033f
C936 VTAIL.n183 VSUBS 0.012914f
C937 VTAIL.n184 VSUBS 0.013674f
C938 VTAIL.n185 VSUBS 0.030525f
C939 VTAIL.n186 VSUBS 0.077371f
C940 VTAIL.n187 VSUBS 0.013674f
C941 VTAIL.n188 VSUBS 0.012914f
C942 VTAIL.n189 VSUBS 0.053909f
C943 VTAIL.n190 VSUBS 0.039013f
C944 VTAIL.n191 VSUBS 1.17553f
C945 VP.t1 VSUBS 3.34814f
C946 VP.t0 VSUBS 2.75607f
C947 VP.n0 VSUBS 4.20515f
.ends

