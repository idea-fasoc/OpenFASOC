* NGSPICE file created from diff_pair_sample_1003.ext - technology: sky130A

.subckt diff_pair_sample_1003 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t7 VN.t0 VDD2.t2 w_n3442_n3268# sky130_fd_pr__pfet_01v8 ad=4.485 pd=23.78 as=1.8975 ps=11.83 w=11.5 l=3.79
X1 B.t11 B.t9 B.t10 w_n3442_n3268# sky130_fd_pr__pfet_01v8 ad=4.485 pd=23.78 as=0 ps=0 w=11.5 l=3.79
X2 B.t8 B.t6 B.t7 w_n3442_n3268# sky130_fd_pr__pfet_01v8 ad=4.485 pd=23.78 as=0 ps=0 w=11.5 l=3.79
X3 VTAIL.t6 VN.t1 VDD2.t1 w_n3442_n3268# sky130_fd_pr__pfet_01v8 ad=4.485 pd=23.78 as=1.8975 ps=11.83 w=11.5 l=3.79
X4 VDD1.t3 VP.t0 VTAIL.t2 w_n3442_n3268# sky130_fd_pr__pfet_01v8 ad=1.8975 pd=11.83 as=4.485 ps=23.78 w=11.5 l=3.79
X5 VTAIL.t3 VP.t1 VDD1.t2 w_n3442_n3268# sky130_fd_pr__pfet_01v8 ad=4.485 pd=23.78 as=1.8975 ps=11.83 w=11.5 l=3.79
X6 B.t5 B.t3 B.t4 w_n3442_n3268# sky130_fd_pr__pfet_01v8 ad=4.485 pd=23.78 as=0 ps=0 w=11.5 l=3.79
X7 VDD2.t0 VN.t2 VTAIL.t5 w_n3442_n3268# sky130_fd_pr__pfet_01v8 ad=1.8975 pd=11.83 as=4.485 ps=23.78 w=11.5 l=3.79
X8 VTAIL.t0 VP.t2 VDD1.t1 w_n3442_n3268# sky130_fd_pr__pfet_01v8 ad=4.485 pd=23.78 as=1.8975 ps=11.83 w=11.5 l=3.79
X9 B.t2 B.t0 B.t1 w_n3442_n3268# sky130_fd_pr__pfet_01v8 ad=4.485 pd=23.78 as=0 ps=0 w=11.5 l=3.79
X10 VDD2.t3 VN.t3 VTAIL.t4 w_n3442_n3268# sky130_fd_pr__pfet_01v8 ad=1.8975 pd=11.83 as=4.485 ps=23.78 w=11.5 l=3.79
X11 VDD1.t0 VP.t3 VTAIL.t1 w_n3442_n3268# sky130_fd_pr__pfet_01v8 ad=1.8975 pd=11.83 as=4.485 ps=23.78 w=11.5 l=3.79
R0 VN.n1 VN.t2 107.081
R1 VN.n0 VN.t0 107.081
R2 VN.n0 VN.t3 105.731
R3 VN.n1 VN.t1 105.731
R4 VN VN.n1 51.6504
R5 VN VN.n0 1.85871
R6 VDD2.n2 VDD2.n0 121.005
R7 VDD2.n2 VDD2.n1 76.7222
R8 VDD2.n1 VDD2.t1 2.82702
R9 VDD2.n1 VDD2.t0 2.82702
R10 VDD2.n0 VDD2.t2 2.82702
R11 VDD2.n0 VDD2.t3 2.82702
R12 VDD2 VDD2.n2 0.0586897
R13 VTAIL.n490 VTAIL.n434 756.745
R14 VTAIL.n56 VTAIL.n0 756.745
R15 VTAIL.n118 VTAIL.n62 756.745
R16 VTAIL.n180 VTAIL.n124 756.745
R17 VTAIL.n428 VTAIL.n372 756.745
R18 VTAIL.n366 VTAIL.n310 756.745
R19 VTAIL.n304 VTAIL.n248 756.745
R20 VTAIL.n242 VTAIL.n186 756.745
R21 VTAIL.n455 VTAIL.n454 585
R22 VTAIL.n457 VTAIL.n456 585
R23 VTAIL.n450 VTAIL.n449 585
R24 VTAIL.n463 VTAIL.n462 585
R25 VTAIL.n465 VTAIL.n464 585
R26 VTAIL.n446 VTAIL.n445 585
R27 VTAIL.n472 VTAIL.n471 585
R28 VTAIL.n473 VTAIL.n444 585
R29 VTAIL.n475 VTAIL.n474 585
R30 VTAIL.n442 VTAIL.n441 585
R31 VTAIL.n481 VTAIL.n480 585
R32 VTAIL.n483 VTAIL.n482 585
R33 VTAIL.n438 VTAIL.n437 585
R34 VTAIL.n489 VTAIL.n488 585
R35 VTAIL.n491 VTAIL.n490 585
R36 VTAIL.n21 VTAIL.n20 585
R37 VTAIL.n23 VTAIL.n22 585
R38 VTAIL.n16 VTAIL.n15 585
R39 VTAIL.n29 VTAIL.n28 585
R40 VTAIL.n31 VTAIL.n30 585
R41 VTAIL.n12 VTAIL.n11 585
R42 VTAIL.n38 VTAIL.n37 585
R43 VTAIL.n39 VTAIL.n10 585
R44 VTAIL.n41 VTAIL.n40 585
R45 VTAIL.n8 VTAIL.n7 585
R46 VTAIL.n47 VTAIL.n46 585
R47 VTAIL.n49 VTAIL.n48 585
R48 VTAIL.n4 VTAIL.n3 585
R49 VTAIL.n55 VTAIL.n54 585
R50 VTAIL.n57 VTAIL.n56 585
R51 VTAIL.n83 VTAIL.n82 585
R52 VTAIL.n85 VTAIL.n84 585
R53 VTAIL.n78 VTAIL.n77 585
R54 VTAIL.n91 VTAIL.n90 585
R55 VTAIL.n93 VTAIL.n92 585
R56 VTAIL.n74 VTAIL.n73 585
R57 VTAIL.n100 VTAIL.n99 585
R58 VTAIL.n101 VTAIL.n72 585
R59 VTAIL.n103 VTAIL.n102 585
R60 VTAIL.n70 VTAIL.n69 585
R61 VTAIL.n109 VTAIL.n108 585
R62 VTAIL.n111 VTAIL.n110 585
R63 VTAIL.n66 VTAIL.n65 585
R64 VTAIL.n117 VTAIL.n116 585
R65 VTAIL.n119 VTAIL.n118 585
R66 VTAIL.n145 VTAIL.n144 585
R67 VTAIL.n147 VTAIL.n146 585
R68 VTAIL.n140 VTAIL.n139 585
R69 VTAIL.n153 VTAIL.n152 585
R70 VTAIL.n155 VTAIL.n154 585
R71 VTAIL.n136 VTAIL.n135 585
R72 VTAIL.n162 VTAIL.n161 585
R73 VTAIL.n163 VTAIL.n134 585
R74 VTAIL.n165 VTAIL.n164 585
R75 VTAIL.n132 VTAIL.n131 585
R76 VTAIL.n171 VTAIL.n170 585
R77 VTAIL.n173 VTAIL.n172 585
R78 VTAIL.n128 VTAIL.n127 585
R79 VTAIL.n179 VTAIL.n178 585
R80 VTAIL.n181 VTAIL.n180 585
R81 VTAIL.n429 VTAIL.n428 585
R82 VTAIL.n427 VTAIL.n426 585
R83 VTAIL.n376 VTAIL.n375 585
R84 VTAIL.n421 VTAIL.n420 585
R85 VTAIL.n419 VTAIL.n418 585
R86 VTAIL.n380 VTAIL.n379 585
R87 VTAIL.n384 VTAIL.n382 585
R88 VTAIL.n413 VTAIL.n412 585
R89 VTAIL.n411 VTAIL.n410 585
R90 VTAIL.n386 VTAIL.n385 585
R91 VTAIL.n405 VTAIL.n404 585
R92 VTAIL.n403 VTAIL.n402 585
R93 VTAIL.n390 VTAIL.n389 585
R94 VTAIL.n397 VTAIL.n396 585
R95 VTAIL.n395 VTAIL.n394 585
R96 VTAIL.n367 VTAIL.n366 585
R97 VTAIL.n365 VTAIL.n364 585
R98 VTAIL.n314 VTAIL.n313 585
R99 VTAIL.n359 VTAIL.n358 585
R100 VTAIL.n357 VTAIL.n356 585
R101 VTAIL.n318 VTAIL.n317 585
R102 VTAIL.n322 VTAIL.n320 585
R103 VTAIL.n351 VTAIL.n350 585
R104 VTAIL.n349 VTAIL.n348 585
R105 VTAIL.n324 VTAIL.n323 585
R106 VTAIL.n343 VTAIL.n342 585
R107 VTAIL.n341 VTAIL.n340 585
R108 VTAIL.n328 VTAIL.n327 585
R109 VTAIL.n335 VTAIL.n334 585
R110 VTAIL.n333 VTAIL.n332 585
R111 VTAIL.n305 VTAIL.n304 585
R112 VTAIL.n303 VTAIL.n302 585
R113 VTAIL.n252 VTAIL.n251 585
R114 VTAIL.n297 VTAIL.n296 585
R115 VTAIL.n295 VTAIL.n294 585
R116 VTAIL.n256 VTAIL.n255 585
R117 VTAIL.n260 VTAIL.n258 585
R118 VTAIL.n289 VTAIL.n288 585
R119 VTAIL.n287 VTAIL.n286 585
R120 VTAIL.n262 VTAIL.n261 585
R121 VTAIL.n281 VTAIL.n280 585
R122 VTAIL.n279 VTAIL.n278 585
R123 VTAIL.n266 VTAIL.n265 585
R124 VTAIL.n273 VTAIL.n272 585
R125 VTAIL.n271 VTAIL.n270 585
R126 VTAIL.n243 VTAIL.n242 585
R127 VTAIL.n241 VTAIL.n240 585
R128 VTAIL.n190 VTAIL.n189 585
R129 VTAIL.n235 VTAIL.n234 585
R130 VTAIL.n233 VTAIL.n232 585
R131 VTAIL.n194 VTAIL.n193 585
R132 VTAIL.n198 VTAIL.n196 585
R133 VTAIL.n227 VTAIL.n226 585
R134 VTAIL.n225 VTAIL.n224 585
R135 VTAIL.n200 VTAIL.n199 585
R136 VTAIL.n219 VTAIL.n218 585
R137 VTAIL.n217 VTAIL.n216 585
R138 VTAIL.n204 VTAIL.n203 585
R139 VTAIL.n211 VTAIL.n210 585
R140 VTAIL.n209 VTAIL.n208 585
R141 VTAIL.n453 VTAIL.t4 329.036
R142 VTAIL.n19 VTAIL.t7 329.036
R143 VTAIL.n81 VTAIL.t1 329.036
R144 VTAIL.n143 VTAIL.t0 329.036
R145 VTAIL.n393 VTAIL.t2 329.036
R146 VTAIL.n331 VTAIL.t3 329.036
R147 VTAIL.n269 VTAIL.t5 329.036
R148 VTAIL.n207 VTAIL.t6 329.036
R149 VTAIL.n456 VTAIL.n455 171.744
R150 VTAIL.n456 VTAIL.n449 171.744
R151 VTAIL.n463 VTAIL.n449 171.744
R152 VTAIL.n464 VTAIL.n463 171.744
R153 VTAIL.n464 VTAIL.n445 171.744
R154 VTAIL.n472 VTAIL.n445 171.744
R155 VTAIL.n473 VTAIL.n472 171.744
R156 VTAIL.n474 VTAIL.n473 171.744
R157 VTAIL.n474 VTAIL.n441 171.744
R158 VTAIL.n481 VTAIL.n441 171.744
R159 VTAIL.n482 VTAIL.n481 171.744
R160 VTAIL.n482 VTAIL.n437 171.744
R161 VTAIL.n489 VTAIL.n437 171.744
R162 VTAIL.n490 VTAIL.n489 171.744
R163 VTAIL.n22 VTAIL.n21 171.744
R164 VTAIL.n22 VTAIL.n15 171.744
R165 VTAIL.n29 VTAIL.n15 171.744
R166 VTAIL.n30 VTAIL.n29 171.744
R167 VTAIL.n30 VTAIL.n11 171.744
R168 VTAIL.n38 VTAIL.n11 171.744
R169 VTAIL.n39 VTAIL.n38 171.744
R170 VTAIL.n40 VTAIL.n39 171.744
R171 VTAIL.n40 VTAIL.n7 171.744
R172 VTAIL.n47 VTAIL.n7 171.744
R173 VTAIL.n48 VTAIL.n47 171.744
R174 VTAIL.n48 VTAIL.n3 171.744
R175 VTAIL.n55 VTAIL.n3 171.744
R176 VTAIL.n56 VTAIL.n55 171.744
R177 VTAIL.n84 VTAIL.n83 171.744
R178 VTAIL.n84 VTAIL.n77 171.744
R179 VTAIL.n91 VTAIL.n77 171.744
R180 VTAIL.n92 VTAIL.n91 171.744
R181 VTAIL.n92 VTAIL.n73 171.744
R182 VTAIL.n100 VTAIL.n73 171.744
R183 VTAIL.n101 VTAIL.n100 171.744
R184 VTAIL.n102 VTAIL.n101 171.744
R185 VTAIL.n102 VTAIL.n69 171.744
R186 VTAIL.n109 VTAIL.n69 171.744
R187 VTAIL.n110 VTAIL.n109 171.744
R188 VTAIL.n110 VTAIL.n65 171.744
R189 VTAIL.n117 VTAIL.n65 171.744
R190 VTAIL.n118 VTAIL.n117 171.744
R191 VTAIL.n146 VTAIL.n145 171.744
R192 VTAIL.n146 VTAIL.n139 171.744
R193 VTAIL.n153 VTAIL.n139 171.744
R194 VTAIL.n154 VTAIL.n153 171.744
R195 VTAIL.n154 VTAIL.n135 171.744
R196 VTAIL.n162 VTAIL.n135 171.744
R197 VTAIL.n163 VTAIL.n162 171.744
R198 VTAIL.n164 VTAIL.n163 171.744
R199 VTAIL.n164 VTAIL.n131 171.744
R200 VTAIL.n171 VTAIL.n131 171.744
R201 VTAIL.n172 VTAIL.n171 171.744
R202 VTAIL.n172 VTAIL.n127 171.744
R203 VTAIL.n179 VTAIL.n127 171.744
R204 VTAIL.n180 VTAIL.n179 171.744
R205 VTAIL.n428 VTAIL.n427 171.744
R206 VTAIL.n427 VTAIL.n375 171.744
R207 VTAIL.n420 VTAIL.n375 171.744
R208 VTAIL.n420 VTAIL.n419 171.744
R209 VTAIL.n419 VTAIL.n379 171.744
R210 VTAIL.n384 VTAIL.n379 171.744
R211 VTAIL.n412 VTAIL.n384 171.744
R212 VTAIL.n412 VTAIL.n411 171.744
R213 VTAIL.n411 VTAIL.n385 171.744
R214 VTAIL.n404 VTAIL.n385 171.744
R215 VTAIL.n404 VTAIL.n403 171.744
R216 VTAIL.n403 VTAIL.n389 171.744
R217 VTAIL.n396 VTAIL.n389 171.744
R218 VTAIL.n396 VTAIL.n395 171.744
R219 VTAIL.n366 VTAIL.n365 171.744
R220 VTAIL.n365 VTAIL.n313 171.744
R221 VTAIL.n358 VTAIL.n313 171.744
R222 VTAIL.n358 VTAIL.n357 171.744
R223 VTAIL.n357 VTAIL.n317 171.744
R224 VTAIL.n322 VTAIL.n317 171.744
R225 VTAIL.n350 VTAIL.n322 171.744
R226 VTAIL.n350 VTAIL.n349 171.744
R227 VTAIL.n349 VTAIL.n323 171.744
R228 VTAIL.n342 VTAIL.n323 171.744
R229 VTAIL.n342 VTAIL.n341 171.744
R230 VTAIL.n341 VTAIL.n327 171.744
R231 VTAIL.n334 VTAIL.n327 171.744
R232 VTAIL.n334 VTAIL.n333 171.744
R233 VTAIL.n304 VTAIL.n303 171.744
R234 VTAIL.n303 VTAIL.n251 171.744
R235 VTAIL.n296 VTAIL.n251 171.744
R236 VTAIL.n296 VTAIL.n295 171.744
R237 VTAIL.n295 VTAIL.n255 171.744
R238 VTAIL.n260 VTAIL.n255 171.744
R239 VTAIL.n288 VTAIL.n260 171.744
R240 VTAIL.n288 VTAIL.n287 171.744
R241 VTAIL.n287 VTAIL.n261 171.744
R242 VTAIL.n280 VTAIL.n261 171.744
R243 VTAIL.n280 VTAIL.n279 171.744
R244 VTAIL.n279 VTAIL.n265 171.744
R245 VTAIL.n272 VTAIL.n265 171.744
R246 VTAIL.n272 VTAIL.n271 171.744
R247 VTAIL.n242 VTAIL.n241 171.744
R248 VTAIL.n241 VTAIL.n189 171.744
R249 VTAIL.n234 VTAIL.n189 171.744
R250 VTAIL.n234 VTAIL.n233 171.744
R251 VTAIL.n233 VTAIL.n193 171.744
R252 VTAIL.n198 VTAIL.n193 171.744
R253 VTAIL.n226 VTAIL.n198 171.744
R254 VTAIL.n226 VTAIL.n225 171.744
R255 VTAIL.n225 VTAIL.n199 171.744
R256 VTAIL.n218 VTAIL.n199 171.744
R257 VTAIL.n218 VTAIL.n217 171.744
R258 VTAIL.n217 VTAIL.n203 171.744
R259 VTAIL.n210 VTAIL.n203 171.744
R260 VTAIL.n210 VTAIL.n209 171.744
R261 VTAIL.n455 VTAIL.t4 85.8723
R262 VTAIL.n21 VTAIL.t7 85.8723
R263 VTAIL.n83 VTAIL.t1 85.8723
R264 VTAIL.n145 VTAIL.t0 85.8723
R265 VTAIL.n395 VTAIL.t2 85.8723
R266 VTAIL.n333 VTAIL.t3 85.8723
R267 VTAIL.n271 VTAIL.t5 85.8723
R268 VTAIL.n209 VTAIL.t6 85.8723
R269 VTAIL.n495 VTAIL.n494 34.1247
R270 VTAIL.n61 VTAIL.n60 34.1247
R271 VTAIL.n123 VTAIL.n122 34.1247
R272 VTAIL.n185 VTAIL.n184 34.1247
R273 VTAIL.n433 VTAIL.n432 34.1247
R274 VTAIL.n371 VTAIL.n370 34.1247
R275 VTAIL.n309 VTAIL.n308 34.1247
R276 VTAIL.n247 VTAIL.n246 34.1247
R277 VTAIL.n495 VTAIL.n433 25.8324
R278 VTAIL.n247 VTAIL.n185 25.8324
R279 VTAIL.n475 VTAIL.n442 13.1884
R280 VTAIL.n41 VTAIL.n8 13.1884
R281 VTAIL.n103 VTAIL.n70 13.1884
R282 VTAIL.n165 VTAIL.n132 13.1884
R283 VTAIL.n382 VTAIL.n380 13.1884
R284 VTAIL.n320 VTAIL.n318 13.1884
R285 VTAIL.n258 VTAIL.n256 13.1884
R286 VTAIL.n196 VTAIL.n194 13.1884
R287 VTAIL.n476 VTAIL.n444 12.8005
R288 VTAIL.n480 VTAIL.n479 12.8005
R289 VTAIL.n42 VTAIL.n10 12.8005
R290 VTAIL.n46 VTAIL.n45 12.8005
R291 VTAIL.n104 VTAIL.n72 12.8005
R292 VTAIL.n108 VTAIL.n107 12.8005
R293 VTAIL.n166 VTAIL.n134 12.8005
R294 VTAIL.n170 VTAIL.n169 12.8005
R295 VTAIL.n418 VTAIL.n417 12.8005
R296 VTAIL.n414 VTAIL.n413 12.8005
R297 VTAIL.n356 VTAIL.n355 12.8005
R298 VTAIL.n352 VTAIL.n351 12.8005
R299 VTAIL.n294 VTAIL.n293 12.8005
R300 VTAIL.n290 VTAIL.n289 12.8005
R301 VTAIL.n232 VTAIL.n231 12.8005
R302 VTAIL.n228 VTAIL.n227 12.8005
R303 VTAIL.n471 VTAIL.n470 12.0247
R304 VTAIL.n483 VTAIL.n440 12.0247
R305 VTAIL.n37 VTAIL.n36 12.0247
R306 VTAIL.n49 VTAIL.n6 12.0247
R307 VTAIL.n99 VTAIL.n98 12.0247
R308 VTAIL.n111 VTAIL.n68 12.0247
R309 VTAIL.n161 VTAIL.n160 12.0247
R310 VTAIL.n173 VTAIL.n130 12.0247
R311 VTAIL.n421 VTAIL.n378 12.0247
R312 VTAIL.n410 VTAIL.n383 12.0247
R313 VTAIL.n359 VTAIL.n316 12.0247
R314 VTAIL.n348 VTAIL.n321 12.0247
R315 VTAIL.n297 VTAIL.n254 12.0247
R316 VTAIL.n286 VTAIL.n259 12.0247
R317 VTAIL.n235 VTAIL.n192 12.0247
R318 VTAIL.n224 VTAIL.n197 12.0247
R319 VTAIL.n469 VTAIL.n446 11.249
R320 VTAIL.n484 VTAIL.n438 11.249
R321 VTAIL.n35 VTAIL.n12 11.249
R322 VTAIL.n50 VTAIL.n4 11.249
R323 VTAIL.n97 VTAIL.n74 11.249
R324 VTAIL.n112 VTAIL.n66 11.249
R325 VTAIL.n159 VTAIL.n136 11.249
R326 VTAIL.n174 VTAIL.n128 11.249
R327 VTAIL.n422 VTAIL.n376 11.249
R328 VTAIL.n409 VTAIL.n386 11.249
R329 VTAIL.n360 VTAIL.n314 11.249
R330 VTAIL.n347 VTAIL.n324 11.249
R331 VTAIL.n298 VTAIL.n252 11.249
R332 VTAIL.n285 VTAIL.n262 11.249
R333 VTAIL.n236 VTAIL.n190 11.249
R334 VTAIL.n223 VTAIL.n200 11.249
R335 VTAIL.n454 VTAIL.n453 10.7239
R336 VTAIL.n20 VTAIL.n19 10.7239
R337 VTAIL.n82 VTAIL.n81 10.7239
R338 VTAIL.n144 VTAIL.n143 10.7239
R339 VTAIL.n394 VTAIL.n393 10.7239
R340 VTAIL.n332 VTAIL.n331 10.7239
R341 VTAIL.n270 VTAIL.n269 10.7239
R342 VTAIL.n208 VTAIL.n207 10.7239
R343 VTAIL.n466 VTAIL.n465 10.4732
R344 VTAIL.n488 VTAIL.n487 10.4732
R345 VTAIL.n32 VTAIL.n31 10.4732
R346 VTAIL.n54 VTAIL.n53 10.4732
R347 VTAIL.n94 VTAIL.n93 10.4732
R348 VTAIL.n116 VTAIL.n115 10.4732
R349 VTAIL.n156 VTAIL.n155 10.4732
R350 VTAIL.n178 VTAIL.n177 10.4732
R351 VTAIL.n426 VTAIL.n425 10.4732
R352 VTAIL.n406 VTAIL.n405 10.4732
R353 VTAIL.n364 VTAIL.n363 10.4732
R354 VTAIL.n344 VTAIL.n343 10.4732
R355 VTAIL.n302 VTAIL.n301 10.4732
R356 VTAIL.n282 VTAIL.n281 10.4732
R357 VTAIL.n240 VTAIL.n239 10.4732
R358 VTAIL.n220 VTAIL.n219 10.4732
R359 VTAIL.n462 VTAIL.n448 9.69747
R360 VTAIL.n491 VTAIL.n436 9.69747
R361 VTAIL.n28 VTAIL.n14 9.69747
R362 VTAIL.n57 VTAIL.n2 9.69747
R363 VTAIL.n90 VTAIL.n76 9.69747
R364 VTAIL.n119 VTAIL.n64 9.69747
R365 VTAIL.n152 VTAIL.n138 9.69747
R366 VTAIL.n181 VTAIL.n126 9.69747
R367 VTAIL.n429 VTAIL.n374 9.69747
R368 VTAIL.n402 VTAIL.n388 9.69747
R369 VTAIL.n367 VTAIL.n312 9.69747
R370 VTAIL.n340 VTAIL.n326 9.69747
R371 VTAIL.n305 VTAIL.n250 9.69747
R372 VTAIL.n278 VTAIL.n264 9.69747
R373 VTAIL.n243 VTAIL.n188 9.69747
R374 VTAIL.n216 VTAIL.n202 9.69747
R375 VTAIL.n494 VTAIL.n493 9.45567
R376 VTAIL.n60 VTAIL.n59 9.45567
R377 VTAIL.n122 VTAIL.n121 9.45567
R378 VTAIL.n184 VTAIL.n183 9.45567
R379 VTAIL.n432 VTAIL.n431 9.45567
R380 VTAIL.n370 VTAIL.n369 9.45567
R381 VTAIL.n308 VTAIL.n307 9.45567
R382 VTAIL.n246 VTAIL.n245 9.45567
R383 VTAIL.n493 VTAIL.n492 9.3005
R384 VTAIL.n436 VTAIL.n435 9.3005
R385 VTAIL.n487 VTAIL.n486 9.3005
R386 VTAIL.n485 VTAIL.n484 9.3005
R387 VTAIL.n440 VTAIL.n439 9.3005
R388 VTAIL.n479 VTAIL.n478 9.3005
R389 VTAIL.n452 VTAIL.n451 9.3005
R390 VTAIL.n459 VTAIL.n458 9.3005
R391 VTAIL.n461 VTAIL.n460 9.3005
R392 VTAIL.n448 VTAIL.n447 9.3005
R393 VTAIL.n467 VTAIL.n466 9.3005
R394 VTAIL.n469 VTAIL.n468 9.3005
R395 VTAIL.n470 VTAIL.n443 9.3005
R396 VTAIL.n477 VTAIL.n476 9.3005
R397 VTAIL.n59 VTAIL.n58 9.3005
R398 VTAIL.n2 VTAIL.n1 9.3005
R399 VTAIL.n53 VTAIL.n52 9.3005
R400 VTAIL.n51 VTAIL.n50 9.3005
R401 VTAIL.n6 VTAIL.n5 9.3005
R402 VTAIL.n45 VTAIL.n44 9.3005
R403 VTAIL.n18 VTAIL.n17 9.3005
R404 VTAIL.n25 VTAIL.n24 9.3005
R405 VTAIL.n27 VTAIL.n26 9.3005
R406 VTAIL.n14 VTAIL.n13 9.3005
R407 VTAIL.n33 VTAIL.n32 9.3005
R408 VTAIL.n35 VTAIL.n34 9.3005
R409 VTAIL.n36 VTAIL.n9 9.3005
R410 VTAIL.n43 VTAIL.n42 9.3005
R411 VTAIL.n121 VTAIL.n120 9.3005
R412 VTAIL.n64 VTAIL.n63 9.3005
R413 VTAIL.n115 VTAIL.n114 9.3005
R414 VTAIL.n113 VTAIL.n112 9.3005
R415 VTAIL.n68 VTAIL.n67 9.3005
R416 VTAIL.n107 VTAIL.n106 9.3005
R417 VTAIL.n80 VTAIL.n79 9.3005
R418 VTAIL.n87 VTAIL.n86 9.3005
R419 VTAIL.n89 VTAIL.n88 9.3005
R420 VTAIL.n76 VTAIL.n75 9.3005
R421 VTAIL.n95 VTAIL.n94 9.3005
R422 VTAIL.n97 VTAIL.n96 9.3005
R423 VTAIL.n98 VTAIL.n71 9.3005
R424 VTAIL.n105 VTAIL.n104 9.3005
R425 VTAIL.n183 VTAIL.n182 9.3005
R426 VTAIL.n126 VTAIL.n125 9.3005
R427 VTAIL.n177 VTAIL.n176 9.3005
R428 VTAIL.n175 VTAIL.n174 9.3005
R429 VTAIL.n130 VTAIL.n129 9.3005
R430 VTAIL.n169 VTAIL.n168 9.3005
R431 VTAIL.n142 VTAIL.n141 9.3005
R432 VTAIL.n149 VTAIL.n148 9.3005
R433 VTAIL.n151 VTAIL.n150 9.3005
R434 VTAIL.n138 VTAIL.n137 9.3005
R435 VTAIL.n157 VTAIL.n156 9.3005
R436 VTAIL.n159 VTAIL.n158 9.3005
R437 VTAIL.n160 VTAIL.n133 9.3005
R438 VTAIL.n167 VTAIL.n166 9.3005
R439 VTAIL.n392 VTAIL.n391 9.3005
R440 VTAIL.n399 VTAIL.n398 9.3005
R441 VTAIL.n401 VTAIL.n400 9.3005
R442 VTAIL.n388 VTAIL.n387 9.3005
R443 VTAIL.n407 VTAIL.n406 9.3005
R444 VTAIL.n409 VTAIL.n408 9.3005
R445 VTAIL.n383 VTAIL.n381 9.3005
R446 VTAIL.n415 VTAIL.n414 9.3005
R447 VTAIL.n431 VTAIL.n430 9.3005
R448 VTAIL.n374 VTAIL.n373 9.3005
R449 VTAIL.n425 VTAIL.n424 9.3005
R450 VTAIL.n423 VTAIL.n422 9.3005
R451 VTAIL.n378 VTAIL.n377 9.3005
R452 VTAIL.n417 VTAIL.n416 9.3005
R453 VTAIL.n330 VTAIL.n329 9.3005
R454 VTAIL.n337 VTAIL.n336 9.3005
R455 VTAIL.n339 VTAIL.n338 9.3005
R456 VTAIL.n326 VTAIL.n325 9.3005
R457 VTAIL.n345 VTAIL.n344 9.3005
R458 VTAIL.n347 VTAIL.n346 9.3005
R459 VTAIL.n321 VTAIL.n319 9.3005
R460 VTAIL.n353 VTAIL.n352 9.3005
R461 VTAIL.n369 VTAIL.n368 9.3005
R462 VTAIL.n312 VTAIL.n311 9.3005
R463 VTAIL.n363 VTAIL.n362 9.3005
R464 VTAIL.n361 VTAIL.n360 9.3005
R465 VTAIL.n316 VTAIL.n315 9.3005
R466 VTAIL.n355 VTAIL.n354 9.3005
R467 VTAIL.n268 VTAIL.n267 9.3005
R468 VTAIL.n275 VTAIL.n274 9.3005
R469 VTAIL.n277 VTAIL.n276 9.3005
R470 VTAIL.n264 VTAIL.n263 9.3005
R471 VTAIL.n283 VTAIL.n282 9.3005
R472 VTAIL.n285 VTAIL.n284 9.3005
R473 VTAIL.n259 VTAIL.n257 9.3005
R474 VTAIL.n291 VTAIL.n290 9.3005
R475 VTAIL.n307 VTAIL.n306 9.3005
R476 VTAIL.n250 VTAIL.n249 9.3005
R477 VTAIL.n301 VTAIL.n300 9.3005
R478 VTAIL.n299 VTAIL.n298 9.3005
R479 VTAIL.n254 VTAIL.n253 9.3005
R480 VTAIL.n293 VTAIL.n292 9.3005
R481 VTAIL.n206 VTAIL.n205 9.3005
R482 VTAIL.n213 VTAIL.n212 9.3005
R483 VTAIL.n215 VTAIL.n214 9.3005
R484 VTAIL.n202 VTAIL.n201 9.3005
R485 VTAIL.n221 VTAIL.n220 9.3005
R486 VTAIL.n223 VTAIL.n222 9.3005
R487 VTAIL.n197 VTAIL.n195 9.3005
R488 VTAIL.n229 VTAIL.n228 9.3005
R489 VTAIL.n245 VTAIL.n244 9.3005
R490 VTAIL.n188 VTAIL.n187 9.3005
R491 VTAIL.n239 VTAIL.n238 9.3005
R492 VTAIL.n237 VTAIL.n236 9.3005
R493 VTAIL.n192 VTAIL.n191 9.3005
R494 VTAIL.n231 VTAIL.n230 9.3005
R495 VTAIL.n461 VTAIL.n450 8.92171
R496 VTAIL.n492 VTAIL.n434 8.92171
R497 VTAIL.n27 VTAIL.n16 8.92171
R498 VTAIL.n58 VTAIL.n0 8.92171
R499 VTAIL.n89 VTAIL.n78 8.92171
R500 VTAIL.n120 VTAIL.n62 8.92171
R501 VTAIL.n151 VTAIL.n140 8.92171
R502 VTAIL.n182 VTAIL.n124 8.92171
R503 VTAIL.n430 VTAIL.n372 8.92171
R504 VTAIL.n401 VTAIL.n390 8.92171
R505 VTAIL.n368 VTAIL.n310 8.92171
R506 VTAIL.n339 VTAIL.n328 8.92171
R507 VTAIL.n306 VTAIL.n248 8.92171
R508 VTAIL.n277 VTAIL.n266 8.92171
R509 VTAIL.n244 VTAIL.n186 8.92171
R510 VTAIL.n215 VTAIL.n204 8.92171
R511 VTAIL.n458 VTAIL.n457 8.14595
R512 VTAIL.n24 VTAIL.n23 8.14595
R513 VTAIL.n86 VTAIL.n85 8.14595
R514 VTAIL.n148 VTAIL.n147 8.14595
R515 VTAIL.n398 VTAIL.n397 8.14595
R516 VTAIL.n336 VTAIL.n335 8.14595
R517 VTAIL.n274 VTAIL.n273 8.14595
R518 VTAIL.n212 VTAIL.n211 8.14595
R519 VTAIL.n454 VTAIL.n452 7.3702
R520 VTAIL.n20 VTAIL.n18 7.3702
R521 VTAIL.n82 VTAIL.n80 7.3702
R522 VTAIL.n144 VTAIL.n142 7.3702
R523 VTAIL.n394 VTAIL.n392 7.3702
R524 VTAIL.n332 VTAIL.n330 7.3702
R525 VTAIL.n270 VTAIL.n268 7.3702
R526 VTAIL.n208 VTAIL.n206 7.3702
R527 VTAIL.n457 VTAIL.n452 5.81868
R528 VTAIL.n23 VTAIL.n18 5.81868
R529 VTAIL.n85 VTAIL.n80 5.81868
R530 VTAIL.n147 VTAIL.n142 5.81868
R531 VTAIL.n397 VTAIL.n392 5.81868
R532 VTAIL.n335 VTAIL.n330 5.81868
R533 VTAIL.n273 VTAIL.n268 5.81868
R534 VTAIL.n211 VTAIL.n206 5.81868
R535 VTAIL.n458 VTAIL.n450 5.04292
R536 VTAIL.n494 VTAIL.n434 5.04292
R537 VTAIL.n24 VTAIL.n16 5.04292
R538 VTAIL.n60 VTAIL.n0 5.04292
R539 VTAIL.n86 VTAIL.n78 5.04292
R540 VTAIL.n122 VTAIL.n62 5.04292
R541 VTAIL.n148 VTAIL.n140 5.04292
R542 VTAIL.n184 VTAIL.n124 5.04292
R543 VTAIL.n432 VTAIL.n372 5.04292
R544 VTAIL.n398 VTAIL.n390 5.04292
R545 VTAIL.n370 VTAIL.n310 5.04292
R546 VTAIL.n336 VTAIL.n328 5.04292
R547 VTAIL.n308 VTAIL.n248 5.04292
R548 VTAIL.n274 VTAIL.n266 5.04292
R549 VTAIL.n246 VTAIL.n186 5.04292
R550 VTAIL.n212 VTAIL.n204 5.04292
R551 VTAIL.n462 VTAIL.n461 4.26717
R552 VTAIL.n492 VTAIL.n491 4.26717
R553 VTAIL.n28 VTAIL.n27 4.26717
R554 VTAIL.n58 VTAIL.n57 4.26717
R555 VTAIL.n90 VTAIL.n89 4.26717
R556 VTAIL.n120 VTAIL.n119 4.26717
R557 VTAIL.n152 VTAIL.n151 4.26717
R558 VTAIL.n182 VTAIL.n181 4.26717
R559 VTAIL.n430 VTAIL.n429 4.26717
R560 VTAIL.n402 VTAIL.n401 4.26717
R561 VTAIL.n368 VTAIL.n367 4.26717
R562 VTAIL.n340 VTAIL.n339 4.26717
R563 VTAIL.n306 VTAIL.n305 4.26717
R564 VTAIL.n278 VTAIL.n277 4.26717
R565 VTAIL.n244 VTAIL.n243 4.26717
R566 VTAIL.n216 VTAIL.n215 4.26717
R567 VTAIL.n309 VTAIL.n247 3.55222
R568 VTAIL.n433 VTAIL.n371 3.55222
R569 VTAIL.n185 VTAIL.n123 3.55222
R570 VTAIL.n465 VTAIL.n448 3.49141
R571 VTAIL.n488 VTAIL.n436 3.49141
R572 VTAIL.n31 VTAIL.n14 3.49141
R573 VTAIL.n54 VTAIL.n2 3.49141
R574 VTAIL.n93 VTAIL.n76 3.49141
R575 VTAIL.n116 VTAIL.n64 3.49141
R576 VTAIL.n155 VTAIL.n138 3.49141
R577 VTAIL.n178 VTAIL.n126 3.49141
R578 VTAIL.n426 VTAIL.n374 3.49141
R579 VTAIL.n405 VTAIL.n388 3.49141
R580 VTAIL.n364 VTAIL.n312 3.49141
R581 VTAIL.n343 VTAIL.n326 3.49141
R582 VTAIL.n302 VTAIL.n250 3.49141
R583 VTAIL.n281 VTAIL.n264 3.49141
R584 VTAIL.n240 VTAIL.n188 3.49141
R585 VTAIL.n219 VTAIL.n202 3.49141
R586 VTAIL.n466 VTAIL.n446 2.71565
R587 VTAIL.n487 VTAIL.n438 2.71565
R588 VTAIL.n32 VTAIL.n12 2.71565
R589 VTAIL.n53 VTAIL.n4 2.71565
R590 VTAIL.n94 VTAIL.n74 2.71565
R591 VTAIL.n115 VTAIL.n66 2.71565
R592 VTAIL.n156 VTAIL.n136 2.71565
R593 VTAIL.n177 VTAIL.n128 2.71565
R594 VTAIL.n425 VTAIL.n376 2.71565
R595 VTAIL.n406 VTAIL.n386 2.71565
R596 VTAIL.n363 VTAIL.n314 2.71565
R597 VTAIL.n344 VTAIL.n324 2.71565
R598 VTAIL.n301 VTAIL.n252 2.71565
R599 VTAIL.n282 VTAIL.n262 2.71565
R600 VTAIL.n239 VTAIL.n190 2.71565
R601 VTAIL.n220 VTAIL.n200 2.71565
R602 VTAIL.n453 VTAIL.n451 2.41282
R603 VTAIL.n19 VTAIL.n17 2.41282
R604 VTAIL.n81 VTAIL.n79 2.41282
R605 VTAIL.n143 VTAIL.n141 2.41282
R606 VTAIL.n393 VTAIL.n391 2.41282
R607 VTAIL.n331 VTAIL.n329 2.41282
R608 VTAIL.n269 VTAIL.n267 2.41282
R609 VTAIL.n207 VTAIL.n205 2.41282
R610 VTAIL.n471 VTAIL.n469 1.93989
R611 VTAIL.n484 VTAIL.n483 1.93989
R612 VTAIL.n37 VTAIL.n35 1.93989
R613 VTAIL.n50 VTAIL.n49 1.93989
R614 VTAIL.n99 VTAIL.n97 1.93989
R615 VTAIL.n112 VTAIL.n111 1.93989
R616 VTAIL.n161 VTAIL.n159 1.93989
R617 VTAIL.n174 VTAIL.n173 1.93989
R618 VTAIL.n422 VTAIL.n421 1.93989
R619 VTAIL.n410 VTAIL.n409 1.93989
R620 VTAIL.n360 VTAIL.n359 1.93989
R621 VTAIL.n348 VTAIL.n347 1.93989
R622 VTAIL.n298 VTAIL.n297 1.93989
R623 VTAIL.n286 VTAIL.n285 1.93989
R624 VTAIL.n236 VTAIL.n235 1.93989
R625 VTAIL.n224 VTAIL.n223 1.93989
R626 VTAIL VTAIL.n61 1.83455
R627 VTAIL VTAIL.n495 1.71817
R628 VTAIL.n470 VTAIL.n444 1.16414
R629 VTAIL.n480 VTAIL.n440 1.16414
R630 VTAIL.n36 VTAIL.n10 1.16414
R631 VTAIL.n46 VTAIL.n6 1.16414
R632 VTAIL.n98 VTAIL.n72 1.16414
R633 VTAIL.n108 VTAIL.n68 1.16414
R634 VTAIL.n160 VTAIL.n134 1.16414
R635 VTAIL.n170 VTAIL.n130 1.16414
R636 VTAIL.n418 VTAIL.n378 1.16414
R637 VTAIL.n413 VTAIL.n383 1.16414
R638 VTAIL.n356 VTAIL.n316 1.16414
R639 VTAIL.n351 VTAIL.n321 1.16414
R640 VTAIL.n294 VTAIL.n254 1.16414
R641 VTAIL.n289 VTAIL.n259 1.16414
R642 VTAIL.n232 VTAIL.n192 1.16414
R643 VTAIL.n227 VTAIL.n197 1.16414
R644 VTAIL.n371 VTAIL.n309 0.470328
R645 VTAIL.n123 VTAIL.n61 0.470328
R646 VTAIL.n476 VTAIL.n475 0.388379
R647 VTAIL.n479 VTAIL.n442 0.388379
R648 VTAIL.n42 VTAIL.n41 0.388379
R649 VTAIL.n45 VTAIL.n8 0.388379
R650 VTAIL.n104 VTAIL.n103 0.388379
R651 VTAIL.n107 VTAIL.n70 0.388379
R652 VTAIL.n166 VTAIL.n165 0.388379
R653 VTAIL.n169 VTAIL.n132 0.388379
R654 VTAIL.n417 VTAIL.n380 0.388379
R655 VTAIL.n414 VTAIL.n382 0.388379
R656 VTAIL.n355 VTAIL.n318 0.388379
R657 VTAIL.n352 VTAIL.n320 0.388379
R658 VTAIL.n293 VTAIL.n256 0.388379
R659 VTAIL.n290 VTAIL.n258 0.388379
R660 VTAIL.n231 VTAIL.n194 0.388379
R661 VTAIL.n228 VTAIL.n196 0.388379
R662 VTAIL.n459 VTAIL.n451 0.155672
R663 VTAIL.n460 VTAIL.n459 0.155672
R664 VTAIL.n460 VTAIL.n447 0.155672
R665 VTAIL.n467 VTAIL.n447 0.155672
R666 VTAIL.n468 VTAIL.n467 0.155672
R667 VTAIL.n468 VTAIL.n443 0.155672
R668 VTAIL.n477 VTAIL.n443 0.155672
R669 VTAIL.n478 VTAIL.n477 0.155672
R670 VTAIL.n478 VTAIL.n439 0.155672
R671 VTAIL.n485 VTAIL.n439 0.155672
R672 VTAIL.n486 VTAIL.n485 0.155672
R673 VTAIL.n486 VTAIL.n435 0.155672
R674 VTAIL.n493 VTAIL.n435 0.155672
R675 VTAIL.n25 VTAIL.n17 0.155672
R676 VTAIL.n26 VTAIL.n25 0.155672
R677 VTAIL.n26 VTAIL.n13 0.155672
R678 VTAIL.n33 VTAIL.n13 0.155672
R679 VTAIL.n34 VTAIL.n33 0.155672
R680 VTAIL.n34 VTAIL.n9 0.155672
R681 VTAIL.n43 VTAIL.n9 0.155672
R682 VTAIL.n44 VTAIL.n43 0.155672
R683 VTAIL.n44 VTAIL.n5 0.155672
R684 VTAIL.n51 VTAIL.n5 0.155672
R685 VTAIL.n52 VTAIL.n51 0.155672
R686 VTAIL.n52 VTAIL.n1 0.155672
R687 VTAIL.n59 VTAIL.n1 0.155672
R688 VTAIL.n87 VTAIL.n79 0.155672
R689 VTAIL.n88 VTAIL.n87 0.155672
R690 VTAIL.n88 VTAIL.n75 0.155672
R691 VTAIL.n95 VTAIL.n75 0.155672
R692 VTAIL.n96 VTAIL.n95 0.155672
R693 VTAIL.n96 VTAIL.n71 0.155672
R694 VTAIL.n105 VTAIL.n71 0.155672
R695 VTAIL.n106 VTAIL.n105 0.155672
R696 VTAIL.n106 VTAIL.n67 0.155672
R697 VTAIL.n113 VTAIL.n67 0.155672
R698 VTAIL.n114 VTAIL.n113 0.155672
R699 VTAIL.n114 VTAIL.n63 0.155672
R700 VTAIL.n121 VTAIL.n63 0.155672
R701 VTAIL.n149 VTAIL.n141 0.155672
R702 VTAIL.n150 VTAIL.n149 0.155672
R703 VTAIL.n150 VTAIL.n137 0.155672
R704 VTAIL.n157 VTAIL.n137 0.155672
R705 VTAIL.n158 VTAIL.n157 0.155672
R706 VTAIL.n158 VTAIL.n133 0.155672
R707 VTAIL.n167 VTAIL.n133 0.155672
R708 VTAIL.n168 VTAIL.n167 0.155672
R709 VTAIL.n168 VTAIL.n129 0.155672
R710 VTAIL.n175 VTAIL.n129 0.155672
R711 VTAIL.n176 VTAIL.n175 0.155672
R712 VTAIL.n176 VTAIL.n125 0.155672
R713 VTAIL.n183 VTAIL.n125 0.155672
R714 VTAIL.n431 VTAIL.n373 0.155672
R715 VTAIL.n424 VTAIL.n373 0.155672
R716 VTAIL.n424 VTAIL.n423 0.155672
R717 VTAIL.n423 VTAIL.n377 0.155672
R718 VTAIL.n416 VTAIL.n377 0.155672
R719 VTAIL.n416 VTAIL.n415 0.155672
R720 VTAIL.n415 VTAIL.n381 0.155672
R721 VTAIL.n408 VTAIL.n381 0.155672
R722 VTAIL.n408 VTAIL.n407 0.155672
R723 VTAIL.n407 VTAIL.n387 0.155672
R724 VTAIL.n400 VTAIL.n387 0.155672
R725 VTAIL.n400 VTAIL.n399 0.155672
R726 VTAIL.n399 VTAIL.n391 0.155672
R727 VTAIL.n369 VTAIL.n311 0.155672
R728 VTAIL.n362 VTAIL.n311 0.155672
R729 VTAIL.n362 VTAIL.n361 0.155672
R730 VTAIL.n361 VTAIL.n315 0.155672
R731 VTAIL.n354 VTAIL.n315 0.155672
R732 VTAIL.n354 VTAIL.n353 0.155672
R733 VTAIL.n353 VTAIL.n319 0.155672
R734 VTAIL.n346 VTAIL.n319 0.155672
R735 VTAIL.n346 VTAIL.n345 0.155672
R736 VTAIL.n345 VTAIL.n325 0.155672
R737 VTAIL.n338 VTAIL.n325 0.155672
R738 VTAIL.n338 VTAIL.n337 0.155672
R739 VTAIL.n337 VTAIL.n329 0.155672
R740 VTAIL.n307 VTAIL.n249 0.155672
R741 VTAIL.n300 VTAIL.n249 0.155672
R742 VTAIL.n300 VTAIL.n299 0.155672
R743 VTAIL.n299 VTAIL.n253 0.155672
R744 VTAIL.n292 VTAIL.n253 0.155672
R745 VTAIL.n292 VTAIL.n291 0.155672
R746 VTAIL.n291 VTAIL.n257 0.155672
R747 VTAIL.n284 VTAIL.n257 0.155672
R748 VTAIL.n284 VTAIL.n283 0.155672
R749 VTAIL.n283 VTAIL.n263 0.155672
R750 VTAIL.n276 VTAIL.n263 0.155672
R751 VTAIL.n276 VTAIL.n275 0.155672
R752 VTAIL.n275 VTAIL.n267 0.155672
R753 VTAIL.n245 VTAIL.n187 0.155672
R754 VTAIL.n238 VTAIL.n187 0.155672
R755 VTAIL.n238 VTAIL.n237 0.155672
R756 VTAIL.n237 VTAIL.n191 0.155672
R757 VTAIL.n230 VTAIL.n191 0.155672
R758 VTAIL.n230 VTAIL.n229 0.155672
R759 VTAIL.n229 VTAIL.n195 0.155672
R760 VTAIL.n222 VTAIL.n195 0.155672
R761 VTAIL.n222 VTAIL.n221 0.155672
R762 VTAIL.n221 VTAIL.n201 0.155672
R763 VTAIL.n214 VTAIL.n201 0.155672
R764 VTAIL.n214 VTAIL.n213 0.155672
R765 VTAIL.n213 VTAIL.n205 0.155672
R766 B.n390 B.n389 585
R767 B.n388 B.n119 585
R768 B.n387 B.n386 585
R769 B.n385 B.n120 585
R770 B.n384 B.n383 585
R771 B.n382 B.n121 585
R772 B.n381 B.n380 585
R773 B.n379 B.n122 585
R774 B.n378 B.n377 585
R775 B.n376 B.n123 585
R776 B.n375 B.n374 585
R777 B.n373 B.n124 585
R778 B.n372 B.n371 585
R779 B.n370 B.n125 585
R780 B.n369 B.n368 585
R781 B.n367 B.n126 585
R782 B.n366 B.n365 585
R783 B.n364 B.n127 585
R784 B.n363 B.n362 585
R785 B.n361 B.n128 585
R786 B.n360 B.n359 585
R787 B.n358 B.n129 585
R788 B.n357 B.n356 585
R789 B.n355 B.n130 585
R790 B.n354 B.n353 585
R791 B.n352 B.n131 585
R792 B.n351 B.n350 585
R793 B.n349 B.n132 585
R794 B.n348 B.n347 585
R795 B.n346 B.n133 585
R796 B.n345 B.n344 585
R797 B.n343 B.n134 585
R798 B.n342 B.n341 585
R799 B.n340 B.n135 585
R800 B.n339 B.n338 585
R801 B.n337 B.n136 585
R802 B.n336 B.n335 585
R803 B.n334 B.n137 585
R804 B.n333 B.n332 585
R805 B.n331 B.n138 585
R806 B.n330 B.n329 585
R807 B.n325 B.n139 585
R808 B.n324 B.n323 585
R809 B.n322 B.n140 585
R810 B.n321 B.n320 585
R811 B.n319 B.n141 585
R812 B.n318 B.n317 585
R813 B.n316 B.n142 585
R814 B.n315 B.n314 585
R815 B.n313 B.n143 585
R816 B.n311 B.n310 585
R817 B.n309 B.n146 585
R818 B.n308 B.n307 585
R819 B.n306 B.n147 585
R820 B.n305 B.n304 585
R821 B.n303 B.n148 585
R822 B.n302 B.n301 585
R823 B.n300 B.n149 585
R824 B.n299 B.n298 585
R825 B.n297 B.n150 585
R826 B.n296 B.n295 585
R827 B.n294 B.n151 585
R828 B.n293 B.n292 585
R829 B.n291 B.n152 585
R830 B.n290 B.n289 585
R831 B.n288 B.n153 585
R832 B.n287 B.n286 585
R833 B.n285 B.n154 585
R834 B.n284 B.n283 585
R835 B.n282 B.n155 585
R836 B.n281 B.n280 585
R837 B.n279 B.n156 585
R838 B.n278 B.n277 585
R839 B.n276 B.n157 585
R840 B.n275 B.n274 585
R841 B.n273 B.n158 585
R842 B.n272 B.n271 585
R843 B.n270 B.n159 585
R844 B.n269 B.n268 585
R845 B.n267 B.n160 585
R846 B.n266 B.n265 585
R847 B.n264 B.n161 585
R848 B.n263 B.n262 585
R849 B.n261 B.n162 585
R850 B.n260 B.n259 585
R851 B.n258 B.n163 585
R852 B.n257 B.n256 585
R853 B.n255 B.n164 585
R854 B.n254 B.n253 585
R855 B.n252 B.n165 585
R856 B.n391 B.n118 585
R857 B.n393 B.n392 585
R858 B.n394 B.n117 585
R859 B.n396 B.n395 585
R860 B.n397 B.n116 585
R861 B.n399 B.n398 585
R862 B.n400 B.n115 585
R863 B.n402 B.n401 585
R864 B.n403 B.n114 585
R865 B.n405 B.n404 585
R866 B.n406 B.n113 585
R867 B.n408 B.n407 585
R868 B.n409 B.n112 585
R869 B.n411 B.n410 585
R870 B.n412 B.n111 585
R871 B.n414 B.n413 585
R872 B.n415 B.n110 585
R873 B.n417 B.n416 585
R874 B.n418 B.n109 585
R875 B.n420 B.n419 585
R876 B.n421 B.n108 585
R877 B.n423 B.n422 585
R878 B.n424 B.n107 585
R879 B.n426 B.n425 585
R880 B.n427 B.n106 585
R881 B.n429 B.n428 585
R882 B.n430 B.n105 585
R883 B.n432 B.n431 585
R884 B.n433 B.n104 585
R885 B.n435 B.n434 585
R886 B.n436 B.n103 585
R887 B.n438 B.n437 585
R888 B.n439 B.n102 585
R889 B.n441 B.n440 585
R890 B.n442 B.n101 585
R891 B.n444 B.n443 585
R892 B.n445 B.n100 585
R893 B.n447 B.n446 585
R894 B.n448 B.n99 585
R895 B.n450 B.n449 585
R896 B.n451 B.n98 585
R897 B.n453 B.n452 585
R898 B.n454 B.n97 585
R899 B.n456 B.n455 585
R900 B.n457 B.n96 585
R901 B.n459 B.n458 585
R902 B.n460 B.n95 585
R903 B.n462 B.n461 585
R904 B.n463 B.n94 585
R905 B.n465 B.n464 585
R906 B.n466 B.n93 585
R907 B.n468 B.n467 585
R908 B.n469 B.n92 585
R909 B.n471 B.n470 585
R910 B.n472 B.n91 585
R911 B.n474 B.n473 585
R912 B.n475 B.n90 585
R913 B.n477 B.n476 585
R914 B.n478 B.n89 585
R915 B.n480 B.n479 585
R916 B.n481 B.n88 585
R917 B.n483 B.n482 585
R918 B.n484 B.n87 585
R919 B.n486 B.n485 585
R920 B.n487 B.n86 585
R921 B.n489 B.n488 585
R922 B.n490 B.n85 585
R923 B.n492 B.n491 585
R924 B.n493 B.n84 585
R925 B.n495 B.n494 585
R926 B.n496 B.n83 585
R927 B.n498 B.n497 585
R928 B.n499 B.n82 585
R929 B.n501 B.n500 585
R930 B.n502 B.n81 585
R931 B.n504 B.n503 585
R932 B.n505 B.n80 585
R933 B.n507 B.n506 585
R934 B.n508 B.n79 585
R935 B.n510 B.n509 585
R936 B.n511 B.n78 585
R937 B.n513 B.n512 585
R938 B.n514 B.n77 585
R939 B.n516 B.n515 585
R940 B.n517 B.n76 585
R941 B.n519 B.n518 585
R942 B.n520 B.n75 585
R943 B.n522 B.n521 585
R944 B.n523 B.n74 585
R945 B.n525 B.n524 585
R946 B.n661 B.n24 585
R947 B.n660 B.n659 585
R948 B.n658 B.n25 585
R949 B.n657 B.n656 585
R950 B.n655 B.n26 585
R951 B.n654 B.n653 585
R952 B.n652 B.n27 585
R953 B.n651 B.n650 585
R954 B.n649 B.n28 585
R955 B.n648 B.n647 585
R956 B.n646 B.n29 585
R957 B.n645 B.n644 585
R958 B.n643 B.n30 585
R959 B.n642 B.n641 585
R960 B.n640 B.n31 585
R961 B.n639 B.n638 585
R962 B.n637 B.n32 585
R963 B.n636 B.n635 585
R964 B.n634 B.n33 585
R965 B.n633 B.n632 585
R966 B.n631 B.n34 585
R967 B.n630 B.n629 585
R968 B.n628 B.n35 585
R969 B.n627 B.n626 585
R970 B.n625 B.n36 585
R971 B.n624 B.n623 585
R972 B.n622 B.n37 585
R973 B.n621 B.n620 585
R974 B.n619 B.n38 585
R975 B.n618 B.n617 585
R976 B.n616 B.n39 585
R977 B.n615 B.n614 585
R978 B.n613 B.n40 585
R979 B.n612 B.n611 585
R980 B.n610 B.n41 585
R981 B.n609 B.n608 585
R982 B.n607 B.n42 585
R983 B.n606 B.n605 585
R984 B.n604 B.n43 585
R985 B.n603 B.n602 585
R986 B.n601 B.n600 585
R987 B.n599 B.n47 585
R988 B.n598 B.n597 585
R989 B.n596 B.n48 585
R990 B.n595 B.n594 585
R991 B.n593 B.n49 585
R992 B.n592 B.n591 585
R993 B.n590 B.n50 585
R994 B.n589 B.n588 585
R995 B.n587 B.n51 585
R996 B.n585 B.n584 585
R997 B.n583 B.n54 585
R998 B.n582 B.n581 585
R999 B.n580 B.n55 585
R1000 B.n579 B.n578 585
R1001 B.n577 B.n56 585
R1002 B.n576 B.n575 585
R1003 B.n574 B.n57 585
R1004 B.n573 B.n572 585
R1005 B.n571 B.n58 585
R1006 B.n570 B.n569 585
R1007 B.n568 B.n59 585
R1008 B.n567 B.n566 585
R1009 B.n565 B.n60 585
R1010 B.n564 B.n563 585
R1011 B.n562 B.n61 585
R1012 B.n561 B.n560 585
R1013 B.n559 B.n62 585
R1014 B.n558 B.n557 585
R1015 B.n556 B.n63 585
R1016 B.n555 B.n554 585
R1017 B.n553 B.n64 585
R1018 B.n552 B.n551 585
R1019 B.n550 B.n65 585
R1020 B.n549 B.n548 585
R1021 B.n547 B.n66 585
R1022 B.n546 B.n545 585
R1023 B.n544 B.n67 585
R1024 B.n543 B.n542 585
R1025 B.n541 B.n68 585
R1026 B.n540 B.n539 585
R1027 B.n538 B.n69 585
R1028 B.n537 B.n536 585
R1029 B.n535 B.n70 585
R1030 B.n534 B.n533 585
R1031 B.n532 B.n71 585
R1032 B.n531 B.n530 585
R1033 B.n529 B.n72 585
R1034 B.n528 B.n527 585
R1035 B.n526 B.n73 585
R1036 B.n663 B.n662 585
R1037 B.n664 B.n23 585
R1038 B.n666 B.n665 585
R1039 B.n667 B.n22 585
R1040 B.n669 B.n668 585
R1041 B.n670 B.n21 585
R1042 B.n672 B.n671 585
R1043 B.n673 B.n20 585
R1044 B.n675 B.n674 585
R1045 B.n676 B.n19 585
R1046 B.n678 B.n677 585
R1047 B.n679 B.n18 585
R1048 B.n681 B.n680 585
R1049 B.n682 B.n17 585
R1050 B.n684 B.n683 585
R1051 B.n685 B.n16 585
R1052 B.n687 B.n686 585
R1053 B.n688 B.n15 585
R1054 B.n690 B.n689 585
R1055 B.n691 B.n14 585
R1056 B.n693 B.n692 585
R1057 B.n694 B.n13 585
R1058 B.n696 B.n695 585
R1059 B.n697 B.n12 585
R1060 B.n699 B.n698 585
R1061 B.n700 B.n11 585
R1062 B.n702 B.n701 585
R1063 B.n703 B.n10 585
R1064 B.n705 B.n704 585
R1065 B.n706 B.n9 585
R1066 B.n708 B.n707 585
R1067 B.n709 B.n8 585
R1068 B.n711 B.n710 585
R1069 B.n712 B.n7 585
R1070 B.n714 B.n713 585
R1071 B.n715 B.n6 585
R1072 B.n717 B.n716 585
R1073 B.n718 B.n5 585
R1074 B.n720 B.n719 585
R1075 B.n721 B.n4 585
R1076 B.n723 B.n722 585
R1077 B.n724 B.n3 585
R1078 B.n726 B.n725 585
R1079 B.n727 B.n0 585
R1080 B.n2 B.n1 585
R1081 B.n188 B.n187 585
R1082 B.n189 B.n186 585
R1083 B.n191 B.n190 585
R1084 B.n192 B.n185 585
R1085 B.n194 B.n193 585
R1086 B.n195 B.n184 585
R1087 B.n197 B.n196 585
R1088 B.n198 B.n183 585
R1089 B.n200 B.n199 585
R1090 B.n201 B.n182 585
R1091 B.n203 B.n202 585
R1092 B.n204 B.n181 585
R1093 B.n206 B.n205 585
R1094 B.n207 B.n180 585
R1095 B.n209 B.n208 585
R1096 B.n210 B.n179 585
R1097 B.n212 B.n211 585
R1098 B.n213 B.n178 585
R1099 B.n215 B.n214 585
R1100 B.n216 B.n177 585
R1101 B.n218 B.n217 585
R1102 B.n219 B.n176 585
R1103 B.n221 B.n220 585
R1104 B.n222 B.n175 585
R1105 B.n224 B.n223 585
R1106 B.n225 B.n174 585
R1107 B.n227 B.n226 585
R1108 B.n228 B.n173 585
R1109 B.n230 B.n229 585
R1110 B.n231 B.n172 585
R1111 B.n233 B.n232 585
R1112 B.n234 B.n171 585
R1113 B.n236 B.n235 585
R1114 B.n237 B.n170 585
R1115 B.n239 B.n238 585
R1116 B.n240 B.n169 585
R1117 B.n242 B.n241 585
R1118 B.n243 B.n168 585
R1119 B.n245 B.n244 585
R1120 B.n246 B.n167 585
R1121 B.n248 B.n247 585
R1122 B.n249 B.n166 585
R1123 B.n251 B.n250 585
R1124 B.n250 B.n165 482.89
R1125 B.n391 B.n390 482.89
R1126 B.n524 B.n73 482.89
R1127 B.n662 B.n661 482.89
R1128 B.n326 B.t10 446.678
R1129 B.n52 B.t8 446.678
R1130 B.n144 B.t4 446.678
R1131 B.n44 B.t2 446.678
R1132 B.n327 B.t11 366.776
R1133 B.n53 B.t7 366.776
R1134 B.n145 B.t5 366.776
R1135 B.n45 B.t1 366.776
R1136 B.n144 B.t3 282.462
R1137 B.n326 B.t9 282.462
R1138 B.n52 B.t6 282.462
R1139 B.n44 B.t0 282.462
R1140 B.n729 B.n728 256.663
R1141 B.n728 B.n727 235.042
R1142 B.n728 B.n2 235.042
R1143 B.n254 B.n165 163.367
R1144 B.n255 B.n254 163.367
R1145 B.n256 B.n255 163.367
R1146 B.n256 B.n163 163.367
R1147 B.n260 B.n163 163.367
R1148 B.n261 B.n260 163.367
R1149 B.n262 B.n261 163.367
R1150 B.n262 B.n161 163.367
R1151 B.n266 B.n161 163.367
R1152 B.n267 B.n266 163.367
R1153 B.n268 B.n267 163.367
R1154 B.n268 B.n159 163.367
R1155 B.n272 B.n159 163.367
R1156 B.n273 B.n272 163.367
R1157 B.n274 B.n273 163.367
R1158 B.n274 B.n157 163.367
R1159 B.n278 B.n157 163.367
R1160 B.n279 B.n278 163.367
R1161 B.n280 B.n279 163.367
R1162 B.n280 B.n155 163.367
R1163 B.n284 B.n155 163.367
R1164 B.n285 B.n284 163.367
R1165 B.n286 B.n285 163.367
R1166 B.n286 B.n153 163.367
R1167 B.n290 B.n153 163.367
R1168 B.n291 B.n290 163.367
R1169 B.n292 B.n291 163.367
R1170 B.n292 B.n151 163.367
R1171 B.n296 B.n151 163.367
R1172 B.n297 B.n296 163.367
R1173 B.n298 B.n297 163.367
R1174 B.n298 B.n149 163.367
R1175 B.n302 B.n149 163.367
R1176 B.n303 B.n302 163.367
R1177 B.n304 B.n303 163.367
R1178 B.n304 B.n147 163.367
R1179 B.n308 B.n147 163.367
R1180 B.n309 B.n308 163.367
R1181 B.n310 B.n309 163.367
R1182 B.n310 B.n143 163.367
R1183 B.n315 B.n143 163.367
R1184 B.n316 B.n315 163.367
R1185 B.n317 B.n316 163.367
R1186 B.n317 B.n141 163.367
R1187 B.n321 B.n141 163.367
R1188 B.n322 B.n321 163.367
R1189 B.n323 B.n322 163.367
R1190 B.n323 B.n139 163.367
R1191 B.n330 B.n139 163.367
R1192 B.n331 B.n330 163.367
R1193 B.n332 B.n331 163.367
R1194 B.n332 B.n137 163.367
R1195 B.n336 B.n137 163.367
R1196 B.n337 B.n336 163.367
R1197 B.n338 B.n337 163.367
R1198 B.n338 B.n135 163.367
R1199 B.n342 B.n135 163.367
R1200 B.n343 B.n342 163.367
R1201 B.n344 B.n343 163.367
R1202 B.n344 B.n133 163.367
R1203 B.n348 B.n133 163.367
R1204 B.n349 B.n348 163.367
R1205 B.n350 B.n349 163.367
R1206 B.n350 B.n131 163.367
R1207 B.n354 B.n131 163.367
R1208 B.n355 B.n354 163.367
R1209 B.n356 B.n355 163.367
R1210 B.n356 B.n129 163.367
R1211 B.n360 B.n129 163.367
R1212 B.n361 B.n360 163.367
R1213 B.n362 B.n361 163.367
R1214 B.n362 B.n127 163.367
R1215 B.n366 B.n127 163.367
R1216 B.n367 B.n366 163.367
R1217 B.n368 B.n367 163.367
R1218 B.n368 B.n125 163.367
R1219 B.n372 B.n125 163.367
R1220 B.n373 B.n372 163.367
R1221 B.n374 B.n373 163.367
R1222 B.n374 B.n123 163.367
R1223 B.n378 B.n123 163.367
R1224 B.n379 B.n378 163.367
R1225 B.n380 B.n379 163.367
R1226 B.n380 B.n121 163.367
R1227 B.n384 B.n121 163.367
R1228 B.n385 B.n384 163.367
R1229 B.n386 B.n385 163.367
R1230 B.n386 B.n119 163.367
R1231 B.n390 B.n119 163.367
R1232 B.n524 B.n523 163.367
R1233 B.n523 B.n522 163.367
R1234 B.n522 B.n75 163.367
R1235 B.n518 B.n75 163.367
R1236 B.n518 B.n517 163.367
R1237 B.n517 B.n516 163.367
R1238 B.n516 B.n77 163.367
R1239 B.n512 B.n77 163.367
R1240 B.n512 B.n511 163.367
R1241 B.n511 B.n510 163.367
R1242 B.n510 B.n79 163.367
R1243 B.n506 B.n79 163.367
R1244 B.n506 B.n505 163.367
R1245 B.n505 B.n504 163.367
R1246 B.n504 B.n81 163.367
R1247 B.n500 B.n81 163.367
R1248 B.n500 B.n499 163.367
R1249 B.n499 B.n498 163.367
R1250 B.n498 B.n83 163.367
R1251 B.n494 B.n83 163.367
R1252 B.n494 B.n493 163.367
R1253 B.n493 B.n492 163.367
R1254 B.n492 B.n85 163.367
R1255 B.n488 B.n85 163.367
R1256 B.n488 B.n487 163.367
R1257 B.n487 B.n486 163.367
R1258 B.n486 B.n87 163.367
R1259 B.n482 B.n87 163.367
R1260 B.n482 B.n481 163.367
R1261 B.n481 B.n480 163.367
R1262 B.n480 B.n89 163.367
R1263 B.n476 B.n89 163.367
R1264 B.n476 B.n475 163.367
R1265 B.n475 B.n474 163.367
R1266 B.n474 B.n91 163.367
R1267 B.n470 B.n91 163.367
R1268 B.n470 B.n469 163.367
R1269 B.n469 B.n468 163.367
R1270 B.n468 B.n93 163.367
R1271 B.n464 B.n93 163.367
R1272 B.n464 B.n463 163.367
R1273 B.n463 B.n462 163.367
R1274 B.n462 B.n95 163.367
R1275 B.n458 B.n95 163.367
R1276 B.n458 B.n457 163.367
R1277 B.n457 B.n456 163.367
R1278 B.n456 B.n97 163.367
R1279 B.n452 B.n97 163.367
R1280 B.n452 B.n451 163.367
R1281 B.n451 B.n450 163.367
R1282 B.n450 B.n99 163.367
R1283 B.n446 B.n99 163.367
R1284 B.n446 B.n445 163.367
R1285 B.n445 B.n444 163.367
R1286 B.n444 B.n101 163.367
R1287 B.n440 B.n101 163.367
R1288 B.n440 B.n439 163.367
R1289 B.n439 B.n438 163.367
R1290 B.n438 B.n103 163.367
R1291 B.n434 B.n103 163.367
R1292 B.n434 B.n433 163.367
R1293 B.n433 B.n432 163.367
R1294 B.n432 B.n105 163.367
R1295 B.n428 B.n105 163.367
R1296 B.n428 B.n427 163.367
R1297 B.n427 B.n426 163.367
R1298 B.n426 B.n107 163.367
R1299 B.n422 B.n107 163.367
R1300 B.n422 B.n421 163.367
R1301 B.n421 B.n420 163.367
R1302 B.n420 B.n109 163.367
R1303 B.n416 B.n109 163.367
R1304 B.n416 B.n415 163.367
R1305 B.n415 B.n414 163.367
R1306 B.n414 B.n111 163.367
R1307 B.n410 B.n111 163.367
R1308 B.n410 B.n409 163.367
R1309 B.n409 B.n408 163.367
R1310 B.n408 B.n113 163.367
R1311 B.n404 B.n113 163.367
R1312 B.n404 B.n403 163.367
R1313 B.n403 B.n402 163.367
R1314 B.n402 B.n115 163.367
R1315 B.n398 B.n115 163.367
R1316 B.n398 B.n397 163.367
R1317 B.n397 B.n396 163.367
R1318 B.n396 B.n117 163.367
R1319 B.n392 B.n117 163.367
R1320 B.n392 B.n391 163.367
R1321 B.n661 B.n660 163.367
R1322 B.n660 B.n25 163.367
R1323 B.n656 B.n25 163.367
R1324 B.n656 B.n655 163.367
R1325 B.n655 B.n654 163.367
R1326 B.n654 B.n27 163.367
R1327 B.n650 B.n27 163.367
R1328 B.n650 B.n649 163.367
R1329 B.n649 B.n648 163.367
R1330 B.n648 B.n29 163.367
R1331 B.n644 B.n29 163.367
R1332 B.n644 B.n643 163.367
R1333 B.n643 B.n642 163.367
R1334 B.n642 B.n31 163.367
R1335 B.n638 B.n31 163.367
R1336 B.n638 B.n637 163.367
R1337 B.n637 B.n636 163.367
R1338 B.n636 B.n33 163.367
R1339 B.n632 B.n33 163.367
R1340 B.n632 B.n631 163.367
R1341 B.n631 B.n630 163.367
R1342 B.n630 B.n35 163.367
R1343 B.n626 B.n35 163.367
R1344 B.n626 B.n625 163.367
R1345 B.n625 B.n624 163.367
R1346 B.n624 B.n37 163.367
R1347 B.n620 B.n37 163.367
R1348 B.n620 B.n619 163.367
R1349 B.n619 B.n618 163.367
R1350 B.n618 B.n39 163.367
R1351 B.n614 B.n39 163.367
R1352 B.n614 B.n613 163.367
R1353 B.n613 B.n612 163.367
R1354 B.n612 B.n41 163.367
R1355 B.n608 B.n41 163.367
R1356 B.n608 B.n607 163.367
R1357 B.n607 B.n606 163.367
R1358 B.n606 B.n43 163.367
R1359 B.n602 B.n43 163.367
R1360 B.n602 B.n601 163.367
R1361 B.n601 B.n47 163.367
R1362 B.n597 B.n47 163.367
R1363 B.n597 B.n596 163.367
R1364 B.n596 B.n595 163.367
R1365 B.n595 B.n49 163.367
R1366 B.n591 B.n49 163.367
R1367 B.n591 B.n590 163.367
R1368 B.n590 B.n589 163.367
R1369 B.n589 B.n51 163.367
R1370 B.n584 B.n51 163.367
R1371 B.n584 B.n583 163.367
R1372 B.n583 B.n582 163.367
R1373 B.n582 B.n55 163.367
R1374 B.n578 B.n55 163.367
R1375 B.n578 B.n577 163.367
R1376 B.n577 B.n576 163.367
R1377 B.n576 B.n57 163.367
R1378 B.n572 B.n57 163.367
R1379 B.n572 B.n571 163.367
R1380 B.n571 B.n570 163.367
R1381 B.n570 B.n59 163.367
R1382 B.n566 B.n59 163.367
R1383 B.n566 B.n565 163.367
R1384 B.n565 B.n564 163.367
R1385 B.n564 B.n61 163.367
R1386 B.n560 B.n61 163.367
R1387 B.n560 B.n559 163.367
R1388 B.n559 B.n558 163.367
R1389 B.n558 B.n63 163.367
R1390 B.n554 B.n63 163.367
R1391 B.n554 B.n553 163.367
R1392 B.n553 B.n552 163.367
R1393 B.n552 B.n65 163.367
R1394 B.n548 B.n65 163.367
R1395 B.n548 B.n547 163.367
R1396 B.n547 B.n546 163.367
R1397 B.n546 B.n67 163.367
R1398 B.n542 B.n67 163.367
R1399 B.n542 B.n541 163.367
R1400 B.n541 B.n540 163.367
R1401 B.n540 B.n69 163.367
R1402 B.n536 B.n69 163.367
R1403 B.n536 B.n535 163.367
R1404 B.n535 B.n534 163.367
R1405 B.n534 B.n71 163.367
R1406 B.n530 B.n71 163.367
R1407 B.n530 B.n529 163.367
R1408 B.n529 B.n528 163.367
R1409 B.n528 B.n73 163.367
R1410 B.n662 B.n23 163.367
R1411 B.n666 B.n23 163.367
R1412 B.n667 B.n666 163.367
R1413 B.n668 B.n667 163.367
R1414 B.n668 B.n21 163.367
R1415 B.n672 B.n21 163.367
R1416 B.n673 B.n672 163.367
R1417 B.n674 B.n673 163.367
R1418 B.n674 B.n19 163.367
R1419 B.n678 B.n19 163.367
R1420 B.n679 B.n678 163.367
R1421 B.n680 B.n679 163.367
R1422 B.n680 B.n17 163.367
R1423 B.n684 B.n17 163.367
R1424 B.n685 B.n684 163.367
R1425 B.n686 B.n685 163.367
R1426 B.n686 B.n15 163.367
R1427 B.n690 B.n15 163.367
R1428 B.n691 B.n690 163.367
R1429 B.n692 B.n691 163.367
R1430 B.n692 B.n13 163.367
R1431 B.n696 B.n13 163.367
R1432 B.n697 B.n696 163.367
R1433 B.n698 B.n697 163.367
R1434 B.n698 B.n11 163.367
R1435 B.n702 B.n11 163.367
R1436 B.n703 B.n702 163.367
R1437 B.n704 B.n703 163.367
R1438 B.n704 B.n9 163.367
R1439 B.n708 B.n9 163.367
R1440 B.n709 B.n708 163.367
R1441 B.n710 B.n709 163.367
R1442 B.n710 B.n7 163.367
R1443 B.n714 B.n7 163.367
R1444 B.n715 B.n714 163.367
R1445 B.n716 B.n715 163.367
R1446 B.n716 B.n5 163.367
R1447 B.n720 B.n5 163.367
R1448 B.n721 B.n720 163.367
R1449 B.n722 B.n721 163.367
R1450 B.n722 B.n3 163.367
R1451 B.n726 B.n3 163.367
R1452 B.n727 B.n726 163.367
R1453 B.n188 B.n2 163.367
R1454 B.n189 B.n188 163.367
R1455 B.n190 B.n189 163.367
R1456 B.n190 B.n185 163.367
R1457 B.n194 B.n185 163.367
R1458 B.n195 B.n194 163.367
R1459 B.n196 B.n195 163.367
R1460 B.n196 B.n183 163.367
R1461 B.n200 B.n183 163.367
R1462 B.n201 B.n200 163.367
R1463 B.n202 B.n201 163.367
R1464 B.n202 B.n181 163.367
R1465 B.n206 B.n181 163.367
R1466 B.n207 B.n206 163.367
R1467 B.n208 B.n207 163.367
R1468 B.n208 B.n179 163.367
R1469 B.n212 B.n179 163.367
R1470 B.n213 B.n212 163.367
R1471 B.n214 B.n213 163.367
R1472 B.n214 B.n177 163.367
R1473 B.n218 B.n177 163.367
R1474 B.n219 B.n218 163.367
R1475 B.n220 B.n219 163.367
R1476 B.n220 B.n175 163.367
R1477 B.n224 B.n175 163.367
R1478 B.n225 B.n224 163.367
R1479 B.n226 B.n225 163.367
R1480 B.n226 B.n173 163.367
R1481 B.n230 B.n173 163.367
R1482 B.n231 B.n230 163.367
R1483 B.n232 B.n231 163.367
R1484 B.n232 B.n171 163.367
R1485 B.n236 B.n171 163.367
R1486 B.n237 B.n236 163.367
R1487 B.n238 B.n237 163.367
R1488 B.n238 B.n169 163.367
R1489 B.n242 B.n169 163.367
R1490 B.n243 B.n242 163.367
R1491 B.n244 B.n243 163.367
R1492 B.n244 B.n167 163.367
R1493 B.n248 B.n167 163.367
R1494 B.n249 B.n248 163.367
R1495 B.n250 B.n249 163.367
R1496 B.n145 B.n144 79.9035
R1497 B.n327 B.n326 79.9035
R1498 B.n53 B.n52 79.9035
R1499 B.n45 B.n44 79.9035
R1500 B.n312 B.n145 59.5399
R1501 B.n328 B.n327 59.5399
R1502 B.n586 B.n53 59.5399
R1503 B.n46 B.n45 59.5399
R1504 B.n663 B.n24 31.3761
R1505 B.n526 B.n525 31.3761
R1506 B.n389 B.n118 31.3761
R1507 B.n252 B.n251 31.3761
R1508 B B.n729 18.0485
R1509 B.n664 B.n663 10.6151
R1510 B.n665 B.n664 10.6151
R1511 B.n665 B.n22 10.6151
R1512 B.n669 B.n22 10.6151
R1513 B.n670 B.n669 10.6151
R1514 B.n671 B.n670 10.6151
R1515 B.n671 B.n20 10.6151
R1516 B.n675 B.n20 10.6151
R1517 B.n676 B.n675 10.6151
R1518 B.n677 B.n676 10.6151
R1519 B.n677 B.n18 10.6151
R1520 B.n681 B.n18 10.6151
R1521 B.n682 B.n681 10.6151
R1522 B.n683 B.n682 10.6151
R1523 B.n683 B.n16 10.6151
R1524 B.n687 B.n16 10.6151
R1525 B.n688 B.n687 10.6151
R1526 B.n689 B.n688 10.6151
R1527 B.n689 B.n14 10.6151
R1528 B.n693 B.n14 10.6151
R1529 B.n694 B.n693 10.6151
R1530 B.n695 B.n694 10.6151
R1531 B.n695 B.n12 10.6151
R1532 B.n699 B.n12 10.6151
R1533 B.n700 B.n699 10.6151
R1534 B.n701 B.n700 10.6151
R1535 B.n701 B.n10 10.6151
R1536 B.n705 B.n10 10.6151
R1537 B.n706 B.n705 10.6151
R1538 B.n707 B.n706 10.6151
R1539 B.n707 B.n8 10.6151
R1540 B.n711 B.n8 10.6151
R1541 B.n712 B.n711 10.6151
R1542 B.n713 B.n712 10.6151
R1543 B.n713 B.n6 10.6151
R1544 B.n717 B.n6 10.6151
R1545 B.n718 B.n717 10.6151
R1546 B.n719 B.n718 10.6151
R1547 B.n719 B.n4 10.6151
R1548 B.n723 B.n4 10.6151
R1549 B.n724 B.n723 10.6151
R1550 B.n725 B.n724 10.6151
R1551 B.n725 B.n0 10.6151
R1552 B.n659 B.n24 10.6151
R1553 B.n659 B.n658 10.6151
R1554 B.n658 B.n657 10.6151
R1555 B.n657 B.n26 10.6151
R1556 B.n653 B.n26 10.6151
R1557 B.n653 B.n652 10.6151
R1558 B.n652 B.n651 10.6151
R1559 B.n651 B.n28 10.6151
R1560 B.n647 B.n28 10.6151
R1561 B.n647 B.n646 10.6151
R1562 B.n646 B.n645 10.6151
R1563 B.n645 B.n30 10.6151
R1564 B.n641 B.n30 10.6151
R1565 B.n641 B.n640 10.6151
R1566 B.n640 B.n639 10.6151
R1567 B.n639 B.n32 10.6151
R1568 B.n635 B.n32 10.6151
R1569 B.n635 B.n634 10.6151
R1570 B.n634 B.n633 10.6151
R1571 B.n633 B.n34 10.6151
R1572 B.n629 B.n34 10.6151
R1573 B.n629 B.n628 10.6151
R1574 B.n628 B.n627 10.6151
R1575 B.n627 B.n36 10.6151
R1576 B.n623 B.n36 10.6151
R1577 B.n623 B.n622 10.6151
R1578 B.n622 B.n621 10.6151
R1579 B.n621 B.n38 10.6151
R1580 B.n617 B.n38 10.6151
R1581 B.n617 B.n616 10.6151
R1582 B.n616 B.n615 10.6151
R1583 B.n615 B.n40 10.6151
R1584 B.n611 B.n40 10.6151
R1585 B.n611 B.n610 10.6151
R1586 B.n610 B.n609 10.6151
R1587 B.n609 B.n42 10.6151
R1588 B.n605 B.n42 10.6151
R1589 B.n605 B.n604 10.6151
R1590 B.n604 B.n603 10.6151
R1591 B.n600 B.n599 10.6151
R1592 B.n599 B.n598 10.6151
R1593 B.n598 B.n48 10.6151
R1594 B.n594 B.n48 10.6151
R1595 B.n594 B.n593 10.6151
R1596 B.n593 B.n592 10.6151
R1597 B.n592 B.n50 10.6151
R1598 B.n588 B.n50 10.6151
R1599 B.n588 B.n587 10.6151
R1600 B.n585 B.n54 10.6151
R1601 B.n581 B.n54 10.6151
R1602 B.n581 B.n580 10.6151
R1603 B.n580 B.n579 10.6151
R1604 B.n579 B.n56 10.6151
R1605 B.n575 B.n56 10.6151
R1606 B.n575 B.n574 10.6151
R1607 B.n574 B.n573 10.6151
R1608 B.n573 B.n58 10.6151
R1609 B.n569 B.n58 10.6151
R1610 B.n569 B.n568 10.6151
R1611 B.n568 B.n567 10.6151
R1612 B.n567 B.n60 10.6151
R1613 B.n563 B.n60 10.6151
R1614 B.n563 B.n562 10.6151
R1615 B.n562 B.n561 10.6151
R1616 B.n561 B.n62 10.6151
R1617 B.n557 B.n62 10.6151
R1618 B.n557 B.n556 10.6151
R1619 B.n556 B.n555 10.6151
R1620 B.n555 B.n64 10.6151
R1621 B.n551 B.n64 10.6151
R1622 B.n551 B.n550 10.6151
R1623 B.n550 B.n549 10.6151
R1624 B.n549 B.n66 10.6151
R1625 B.n545 B.n66 10.6151
R1626 B.n545 B.n544 10.6151
R1627 B.n544 B.n543 10.6151
R1628 B.n543 B.n68 10.6151
R1629 B.n539 B.n68 10.6151
R1630 B.n539 B.n538 10.6151
R1631 B.n538 B.n537 10.6151
R1632 B.n537 B.n70 10.6151
R1633 B.n533 B.n70 10.6151
R1634 B.n533 B.n532 10.6151
R1635 B.n532 B.n531 10.6151
R1636 B.n531 B.n72 10.6151
R1637 B.n527 B.n72 10.6151
R1638 B.n527 B.n526 10.6151
R1639 B.n525 B.n74 10.6151
R1640 B.n521 B.n74 10.6151
R1641 B.n521 B.n520 10.6151
R1642 B.n520 B.n519 10.6151
R1643 B.n519 B.n76 10.6151
R1644 B.n515 B.n76 10.6151
R1645 B.n515 B.n514 10.6151
R1646 B.n514 B.n513 10.6151
R1647 B.n513 B.n78 10.6151
R1648 B.n509 B.n78 10.6151
R1649 B.n509 B.n508 10.6151
R1650 B.n508 B.n507 10.6151
R1651 B.n507 B.n80 10.6151
R1652 B.n503 B.n80 10.6151
R1653 B.n503 B.n502 10.6151
R1654 B.n502 B.n501 10.6151
R1655 B.n501 B.n82 10.6151
R1656 B.n497 B.n82 10.6151
R1657 B.n497 B.n496 10.6151
R1658 B.n496 B.n495 10.6151
R1659 B.n495 B.n84 10.6151
R1660 B.n491 B.n84 10.6151
R1661 B.n491 B.n490 10.6151
R1662 B.n490 B.n489 10.6151
R1663 B.n489 B.n86 10.6151
R1664 B.n485 B.n86 10.6151
R1665 B.n485 B.n484 10.6151
R1666 B.n484 B.n483 10.6151
R1667 B.n483 B.n88 10.6151
R1668 B.n479 B.n88 10.6151
R1669 B.n479 B.n478 10.6151
R1670 B.n478 B.n477 10.6151
R1671 B.n477 B.n90 10.6151
R1672 B.n473 B.n90 10.6151
R1673 B.n473 B.n472 10.6151
R1674 B.n472 B.n471 10.6151
R1675 B.n471 B.n92 10.6151
R1676 B.n467 B.n92 10.6151
R1677 B.n467 B.n466 10.6151
R1678 B.n466 B.n465 10.6151
R1679 B.n465 B.n94 10.6151
R1680 B.n461 B.n94 10.6151
R1681 B.n461 B.n460 10.6151
R1682 B.n460 B.n459 10.6151
R1683 B.n459 B.n96 10.6151
R1684 B.n455 B.n96 10.6151
R1685 B.n455 B.n454 10.6151
R1686 B.n454 B.n453 10.6151
R1687 B.n453 B.n98 10.6151
R1688 B.n449 B.n98 10.6151
R1689 B.n449 B.n448 10.6151
R1690 B.n448 B.n447 10.6151
R1691 B.n447 B.n100 10.6151
R1692 B.n443 B.n100 10.6151
R1693 B.n443 B.n442 10.6151
R1694 B.n442 B.n441 10.6151
R1695 B.n441 B.n102 10.6151
R1696 B.n437 B.n102 10.6151
R1697 B.n437 B.n436 10.6151
R1698 B.n436 B.n435 10.6151
R1699 B.n435 B.n104 10.6151
R1700 B.n431 B.n104 10.6151
R1701 B.n431 B.n430 10.6151
R1702 B.n430 B.n429 10.6151
R1703 B.n429 B.n106 10.6151
R1704 B.n425 B.n106 10.6151
R1705 B.n425 B.n424 10.6151
R1706 B.n424 B.n423 10.6151
R1707 B.n423 B.n108 10.6151
R1708 B.n419 B.n108 10.6151
R1709 B.n419 B.n418 10.6151
R1710 B.n418 B.n417 10.6151
R1711 B.n417 B.n110 10.6151
R1712 B.n413 B.n110 10.6151
R1713 B.n413 B.n412 10.6151
R1714 B.n412 B.n411 10.6151
R1715 B.n411 B.n112 10.6151
R1716 B.n407 B.n112 10.6151
R1717 B.n407 B.n406 10.6151
R1718 B.n406 B.n405 10.6151
R1719 B.n405 B.n114 10.6151
R1720 B.n401 B.n114 10.6151
R1721 B.n401 B.n400 10.6151
R1722 B.n400 B.n399 10.6151
R1723 B.n399 B.n116 10.6151
R1724 B.n395 B.n116 10.6151
R1725 B.n395 B.n394 10.6151
R1726 B.n394 B.n393 10.6151
R1727 B.n393 B.n118 10.6151
R1728 B.n187 B.n1 10.6151
R1729 B.n187 B.n186 10.6151
R1730 B.n191 B.n186 10.6151
R1731 B.n192 B.n191 10.6151
R1732 B.n193 B.n192 10.6151
R1733 B.n193 B.n184 10.6151
R1734 B.n197 B.n184 10.6151
R1735 B.n198 B.n197 10.6151
R1736 B.n199 B.n198 10.6151
R1737 B.n199 B.n182 10.6151
R1738 B.n203 B.n182 10.6151
R1739 B.n204 B.n203 10.6151
R1740 B.n205 B.n204 10.6151
R1741 B.n205 B.n180 10.6151
R1742 B.n209 B.n180 10.6151
R1743 B.n210 B.n209 10.6151
R1744 B.n211 B.n210 10.6151
R1745 B.n211 B.n178 10.6151
R1746 B.n215 B.n178 10.6151
R1747 B.n216 B.n215 10.6151
R1748 B.n217 B.n216 10.6151
R1749 B.n217 B.n176 10.6151
R1750 B.n221 B.n176 10.6151
R1751 B.n222 B.n221 10.6151
R1752 B.n223 B.n222 10.6151
R1753 B.n223 B.n174 10.6151
R1754 B.n227 B.n174 10.6151
R1755 B.n228 B.n227 10.6151
R1756 B.n229 B.n228 10.6151
R1757 B.n229 B.n172 10.6151
R1758 B.n233 B.n172 10.6151
R1759 B.n234 B.n233 10.6151
R1760 B.n235 B.n234 10.6151
R1761 B.n235 B.n170 10.6151
R1762 B.n239 B.n170 10.6151
R1763 B.n240 B.n239 10.6151
R1764 B.n241 B.n240 10.6151
R1765 B.n241 B.n168 10.6151
R1766 B.n245 B.n168 10.6151
R1767 B.n246 B.n245 10.6151
R1768 B.n247 B.n246 10.6151
R1769 B.n247 B.n166 10.6151
R1770 B.n251 B.n166 10.6151
R1771 B.n253 B.n252 10.6151
R1772 B.n253 B.n164 10.6151
R1773 B.n257 B.n164 10.6151
R1774 B.n258 B.n257 10.6151
R1775 B.n259 B.n258 10.6151
R1776 B.n259 B.n162 10.6151
R1777 B.n263 B.n162 10.6151
R1778 B.n264 B.n263 10.6151
R1779 B.n265 B.n264 10.6151
R1780 B.n265 B.n160 10.6151
R1781 B.n269 B.n160 10.6151
R1782 B.n270 B.n269 10.6151
R1783 B.n271 B.n270 10.6151
R1784 B.n271 B.n158 10.6151
R1785 B.n275 B.n158 10.6151
R1786 B.n276 B.n275 10.6151
R1787 B.n277 B.n276 10.6151
R1788 B.n277 B.n156 10.6151
R1789 B.n281 B.n156 10.6151
R1790 B.n282 B.n281 10.6151
R1791 B.n283 B.n282 10.6151
R1792 B.n283 B.n154 10.6151
R1793 B.n287 B.n154 10.6151
R1794 B.n288 B.n287 10.6151
R1795 B.n289 B.n288 10.6151
R1796 B.n289 B.n152 10.6151
R1797 B.n293 B.n152 10.6151
R1798 B.n294 B.n293 10.6151
R1799 B.n295 B.n294 10.6151
R1800 B.n295 B.n150 10.6151
R1801 B.n299 B.n150 10.6151
R1802 B.n300 B.n299 10.6151
R1803 B.n301 B.n300 10.6151
R1804 B.n301 B.n148 10.6151
R1805 B.n305 B.n148 10.6151
R1806 B.n306 B.n305 10.6151
R1807 B.n307 B.n306 10.6151
R1808 B.n307 B.n146 10.6151
R1809 B.n311 B.n146 10.6151
R1810 B.n314 B.n313 10.6151
R1811 B.n314 B.n142 10.6151
R1812 B.n318 B.n142 10.6151
R1813 B.n319 B.n318 10.6151
R1814 B.n320 B.n319 10.6151
R1815 B.n320 B.n140 10.6151
R1816 B.n324 B.n140 10.6151
R1817 B.n325 B.n324 10.6151
R1818 B.n329 B.n325 10.6151
R1819 B.n333 B.n138 10.6151
R1820 B.n334 B.n333 10.6151
R1821 B.n335 B.n334 10.6151
R1822 B.n335 B.n136 10.6151
R1823 B.n339 B.n136 10.6151
R1824 B.n340 B.n339 10.6151
R1825 B.n341 B.n340 10.6151
R1826 B.n341 B.n134 10.6151
R1827 B.n345 B.n134 10.6151
R1828 B.n346 B.n345 10.6151
R1829 B.n347 B.n346 10.6151
R1830 B.n347 B.n132 10.6151
R1831 B.n351 B.n132 10.6151
R1832 B.n352 B.n351 10.6151
R1833 B.n353 B.n352 10.6151
R1834 B.n353 B.n130 10.6151
R1835 B.n357 B.n130 10.6151
R1836 B.n358 B.n357 10.6151
R1837 B.n359 B.n358 10.6151
R1838 B.n359 B.n128 10.6151
R1839 B.n363 B.n128 10.6151
R1840 B.n364 B.n363 10.6151
R1841 B.n365 B.n364 10.6151
R1842 B.n365 B.n126 10.6151
R1843 B.n369 B.n126 10.6151
R1844 B.n370 B.n369 10.6151
R1845 B.n371 B.n370 10.6151
R1846 B.n371 B.n124 10.6151
R1847 B.n375 B.n124 10.6151
R1848 B.n376 B.n375 10.6151
R1849 B.n377 B.n376 10.6151
R1850 B.n377 B.n122 10.6151
R1851 B.n381 B.n122 10.6151
R1852 B.n382 B.n381 10.6151
R1853 B.n383 B.n382 10.6151
R1854 B.n383 B.n120 10.6151
R1855 B.n387 B.n120 10.6151
R1856 B.n388 B.n387 10.6151
R1857 B.n389 B.n388 10.6151
R1858 B.n603 B.n46 9.36635
R1859 B.n586 B.n585 9.36635
R1860 B.n312 B.n311 9.36635
R1861 B.n328 B.n138 9.36635
R1862 B.n729 B.n0 8.11757
R1863 B.n729 B.n1 8.11757
R1864 B.n600 B.n46 1.24928
R1865 B.n587 B.n586 1.24928
R1866 B.n313 B.n312 1.24928
R1867 B.n329 B.n328 1.24928
R1868 VP.n21 VP.n20 161.3
R1869 VP.n19 VP.n1 161.3
R1870 VP.n18 VP.n17 161.3
R1871 VP.n16 VP.n2 161.3
R1872 VP.n15 VP.n14 161.3
R1873 VP.n13 VP.n3 161.3
R1874 VP.n12 VP.n11 161.3
R1875 VP.n10 VP.n4 161.3
R1876 VP.n9 VP.n8 161.3
R1877 VP.n5 VP.t1 107.081
R1878 VP.n5 VP.t0 105.731
R1879 VP.n7 VP.n6 87.2945
R1880 VP.n22 VP.n0 87.2945
R1881 VP.n7 VP.t2 73.1271
R1882 VP.n0 VP.t3 73.1271
R1883 VP.n6 VP.n5 51.4851
R1884 VP.n14 VP.n13 40.577
R1885 VP.n14 VP.n2 40.577
R1886 VP.n8 VP.n4 24.5923
R1887 VP.n12 VP.n4 24.5923
R1888 VP.n13 VP.n12 24.5923
R1889 VP.n18 VP.n2 24.5923
R1890 VP.n19 VP.n18 24.5923
R1891 VP.n20 VP.n19 24.5923
R1892 VP.n8 VP.n7 2.95152
R1893 VP.n20 VP.n0 2.95152
R1894 VP.n9 VP.n6 0.354861
R1895 VP.n22 VP.n21 0.354861
R1896 VP VP.n22 0.267071
R1897 VP.n10 VP.n9 0.189894
R1898 VP.n11 VP.n10 0.189894
R1899 VP.n11 VP.n3 0.189894
R1900 VP.n15 VP.n3 0.189894
R1901 VP.n16 VP.n15 0.189894
R1902 VP.n17 VP.n16 0.189894
R1903 VP.n17 VP.n1 0.189894
R1904 VP.n21 VP.n1 0.189894
R1905 VDD1 VDD1.n1 121.531
R1906 VDD1 VDD1.n0 76.7804
R1907 VDD1.n0 VDD1.t2 2.82702
R1908 VDD1.n0 VDD1.t3 2.82702
R1909 VDD1.n1 VDD1.t1 2.82702
R1910 VDD1.n1 VDD1.t0 2.82702
C0 VDD2 VDD1 1.31506f
C1 VDD2 VN 4.83908f
C2 VDD1 VTAIL 5.64032f
C3 VTAIL VN 4.94569f
C4 VDD1 w_n3442_n3268# 1.65919f
C5 VN w_n3442_n3268# 6.03587f
C6 VDD2 VP 0.470216f
C7 VTAIL VP 4.9598f
C8 B VDD1 1.45922f
C9 B VN 1.33333f
C10 VP w_n3442_n3268# 6.48136f
C11 VDD2 VTAIL 5.702509f
C12 VDD2 w_n3442_n3268# 1.74154f
C13 B VP 2.07815f
C14 VTAIL w_n3442_n3268# 3.90352f
C15 VDD1 VN 0.150264f
C16 B VDD2 1.53106f
C17 B VTAIL 5.25055f
C18 B w_n3442_n3268# 10.569f
C19 VDD1 VP 5.15799f
C20 VP VN 6.95183f
C21 VDD2 VSUBS 1.125853f
C22 VDD1 VSUBS 6.386f
C23 VTAIL VSUBS 1.352534f
C24 VN VSUBS 6.11212f
C25 VP VSUBS 2.894112f
C26 B VSUBS 5.258322f
C27 w_n3442_n3268# VSUBS 0.138575p
C28 VDD1.t2 VSUBS 0.252407f
C29 VDD1.t3 VSUBS 0.252407f
C30 VDD1.n0 VSUBS 1.96255f
C31 VDD1.t1 VSUBS 0.252407f
C32 VDD1.t0 VSUBS 0.252407f
C33 VDD1.n1 VSUBS 2.742f
C34 VP.t3 VSUBS 3.68444f
C35 VP.n0 VSUBS 1.40883f
C36 VP.n1 VSUBS 0.031065f
C37 VP.n2 VSUBS 0.061416f
C38 VP.n3 VSUBS 0.031065f
C39 VP.n4 VSUBS 0.057607f
C40 VP.t1 VSUBS 4.17528f
C41 VP.t0 VSUBS 4.15671f
C42 VP.n5 VSUBS 4.49055f
C43 VP.n6 VSUBS 1.87056f
C44 VP.t2 VSUBS 3.68444f
C45 VP.n7 VSUBS 1.40883f
C46 VP.n8 VSUBS 0.03258f
C47 VP.n9 VSUBS 0.05013f
C48 VP.n10 VSUBS 0.031065f
C49 VP.n11 VSUBS 0.031065f
C50 VP.n12 VSUBS 0.057607f
C51 VP.n13 VSUBS 0.061416f
C52 VP.n14 VSUBS 0.02509f
C53 VP.n15 VSUBS 0.031065f
C54 VP.n16 VSUBS 0.031065f
C55 VP.n17 VSUBS 0.031065f
C56 VP.n18 VSUBS 0.057607f
C57 VP.n19 VSUBS 0.057607f
C58 VP.n20 VSUBS 0.03258f
C59 VP.n21 VSUBS 0.05013f
C60 VP.n22 VSUBS 0.095077f
C61 B.n0 VSUBS 0.006275f
C62 B.n1 VSUBS 0.006275f
C63 B.n2 VSUBS 0.00928f
C64 B.n3 VSUBS 0.007112f
C65 B.n4 VSUBS 0.007112f
C66 B.n5 VSUBS 0.007112f
C67 B.n6 VSUBS 0.007112f
C68 B.n7 VSUBS 0.007112f
C69 B.n8 VSUBS 0.007112f
C70 B.n9 VSUBS 0.007112f
C71 B.n10 VSUBS 0.007112f
C72 B.n11 VSUBS 0.007112f
C73 B.n12 VSUBS 0.007112f
C74 B.n13 VSUBS 0.007112f
C75 B.n14 VSUBS 0.007112f
C76 B.n15 VSUBS 0.007112f
C77 B.n16 VSUBS 0.007112f
C78 B.n17 VSUBS 0.007112f
C79 B.n18 VSUBS 0.007112f
C80 B.n19 VSUBS 0.007112f
C81 B.n20 VSUBS 0.007112f
C82 B.n21 VSUBS 0.007112f
C83 B.n22 VSUBS 0.007112f
C84 B.n23 VSUBS 0.007112f
C85 B.n24 VSUBS 0.016648f
C86 B.n25 VSUBS 0.007112f
C87 B.n26 VSUBS 0.007112f
C88 B.n27 VSUBS 0.007112f
C89 B.n28 VSUBS 0.007112f
C90 B.n29 VSUBS 0.007112f
C91 B.n30 VSUBS 0.007112f
C92 B.n31 VSUBS 0.007112f
C93 B.n32 VSUBS 0.007112f
C94 B.n33 VSUBS 0.007112f
C95 B.n34 VSUBS 0.007112f
C96 B.n35 VSUBS 0.007112f
C97 B.n36 VSUBS 0.007112f
C98 B.n37 VSUBS 0.007112f
C99 B.n38 VSUBS 0.007112f
C100 B.n39 VSUBS 0.007112f
C101 B.n40 VSUBS 0.007112f
C102 B.n41 VSUBS 0.007112f
C103 B.n42 VSUBS 0.007112f
C104 B.n43 VSUBS 0.007112f
C105 B.t1 VSUBS 0.203319f
C106 B.t2 VSUBS 0.246863f
C107 B.t0 VSUBS 2.0694f
C108 B.n44 VSUBS 0.394253f
C109 B.n45 VSUBS 0.253565f
C110 B.n46 VSUBS 0.016477f
C111 B.n47 VSUBS 0.007112f
C112 B.n48 VSUBS 0.007112f
C113 B.n49 VSUBS 0.007112f
C114 B.n50 VSUBS 0.007112f
C115 B.n51 VSUBS 0.007112f
C116 B.t7 VSUBS 0.203322f
C117 B.t8 VSUBS 0.246865f
C118 B.t6 VSUBS 2.0694f
C119 B.n52 VSUBS 0.394251f
C120 B.n53 VSUBS 0.253562f
C121 B.n54 VSUBS 0.007112f
C122 B.n55 VSUBS 0.007112f
C123 B.n56 VSUBS 0.007112f
C124 B.n57 VSUBS 0.007112f
C125 B.n58 VSUBS 0.007112f
C126 B.n59 VSUBS 0.007112f
C127 B.n60 VSUBS 0.007112f
C128 B.n61 VSUBS 0.007112f
C129 B.n62 VSUBS 0.007112f
C130 B.n63 VSUBS 0.007112f
C131 B.n64 VSUBS 0.007112f
C132 B.n65 VSUBS 0.007112f
C133 B.n66 VSUBS 0.007112f
C134 B.n67 VSUBS 0.007112f
C135 B.n68 VSUBS 0.007112f
C136 B.n69 VSUBS 0.007112f
C137 B.n70 VSUBS 0.007112f
C138 B.n71 VSUBS 0.007112f
C139 B.n72 VSUBS 0.007112f
C140 B.n73 VSUBS 0.016648f
C141 B.n74 VSUBS 0.007112f
C142 B.n75 VSUBS 0.007112f
C143 B.n76 VSUBS 0.007112f
C144 B.n77 VSUBS 0.007112f
C145 B.n78 VSUBS 0.007112f
C146 B.n79 VSUBS 0.007112f
C147 B.n80 VSUBS 0.007112f
C148 B.n81 VSUBS 0.007112f
C149 B.n82 VSUBS 0.007112f
C150 B.n83 VSUBS 0.007112f
C151 B.n84 VSUBS 0.007112f
C152 B.n85 VSUBS 0.007112f
C153 B.n86 VSUBS 0.007112f
C154 B.n87 VSUBS 0.007112f
C155 B.n88 VSUBS 0.007112f
C156 B.n89 VSUBS 0.007112f
C157 B.n90 VSUBS 0.007112f
C158 B.n91 VSUBS 0.007112f
C159 B.n92 VSUBS 0.007112f
C160 B.n93 VSUBS 0.007112f
C161 B.n94 VSUBS 0.007112f
C162 B.n95 VSUBS 0.007112f
C163 B.n96 VSUBS 0.007112f
C164 B.n97 VSUBS 0.007112f
C165 B.n98 VSUBS 0.007112f
C166 B.n99 VSUBS 0.007112f
C167 B.n100 VSUBS 0.007112f
C168 B.n101 VSUBS 0.007112f
C169 B.n102 VSUBS 0.007112f
C170 B.n103 VSUBS 0.007112f
C171 B.n104 VSUBS 0.007112f
C172 B.n105 VSUBS 0.007112f
C173 B.n106 VSUBS 0.007112f
C174 B.n107 VSUBS 0.007112f
C175 B.n108 VSUBS 0.007112f
C176 B.n109 VSUBS 0.007112f
C177 B.n110 VSUBS 0.007112f
C178 B.n111 VSUBS 0.007112f
C179 B.n112 VSUBS 0.007112f
C180 B.n113 VSUBS 0.007112f
C181 B.n114 VSUBS 0.007112f
C182 B.n115 VSUBS 0.007112f
C183 B.n116 VSUBS 0.007112f
C184 B.n117 VSUBS 0.007112f
C185 B.n118 VSUBS 0.016648f
C186 B.n119 VSUBS 0.007112f
C187 B.n120 VSUBS 0.007112f
C188 B.n121 VSUBS 0.007112f
C189 B.n122 VSUBS 0.007112f
C190 B.n123 VSUBS 0.007112f
C191 B.n124 VSUBS 0.007112f
C192 B.n125 VSUBS 0.007112f
C193 B.n126 VSUBS 0.007112f
C194 B.n127 VSUBS 0.007112f
C195 B.n128 VSUBS 0.007112f
C196 B.n129 VSUBS 0.007112f
C197 B.n130 VSUBS 0.007112f
C198 B.n131 VSUBS 0.007112f
C199 B.n132 VSUBS 0.007112f
C200 B.n133 VSUBS 0.007112f
C201 B.n134 VSUBS 0.007112f
C202 B.n135 VSUBS 0.007112f
C203 B.n136 VSUBS 0.007112f
C204 B.n137 VSUBS 0.007112f
C205 B.n138 VSUBS 0.006693f
C206 B.n139 VSUBS 0.007112f
C207 B.n140 VSUBS 0.007112f
C208 B.n141 VSUBS 0.007112f
C209 B.n142 VSUBS 0.007112f
C210 B.n143 VSUBS 0.007112f
C211 B.t5 VSUBS 0.203319f
C212 B.t4 VSUBS 0.246863f
C213 B.t3 VSUBS 2.0694f
C214 B.n144 VSUBS 0.394253f
C215 B.n145 VSUBS 0.253565f
C216 B.n146 VSUBS 0.007112f
C217 B.n147 VSUBS 0.007112f
C218 B.n148 VSUBS 0.007112f
C219 B.n149 VSUBS 0.007112f
C220 B.n150 VSUBS 0.007112f
C221 B.n151 VSUBS 0.007112f
C222 B.n152 VSUBS 0.007112f
C223 B.n153 VSUBS 0.007112f
C224 B.n154 VSUBS 0.007112f
C225 B.n155 VSUBS 0.007112f
C226 B.n156 VSUBS 0.007112f
C227 B.n157 VSUBS 0.007112f
C228 B.n158 VSUBS 0.007112f
C229 B.n159 VSUBS 0.007112f
C230 B.n160 VSUBS 0.007112f
C231 B.n161 VSUBS 0.007112f
C232 B.n162 VSUBS 0.007112f
C233 B.n163 VSUBS 0.007112f
C234 B.n164 VSUBS 0.007112f
C235 B.n165 VSUBS 0.016648f
C236 B.n166 VSUBS 0.007112f
C237 B.n167 VSUBS 0.007112f
C238 B.n168 VSUBS 0.007112f
C239 B.n169 VSUBS 0.007112f
C240 B.n170 VSUBS 0.007112f
C241 B.n171 VSUBS 0.007112f
C242 B.n172 VSUBS 0.007112f
C243 B.n173 VSUBS 0.007112f
C244 B.n174 VSUBS 0.007112f
C245 B.n175 VSUBS 0.007112f
C246 B.n176 VSUBS 0.007112f
C247 B.n177 VSUBS 0.007112f
C248 B.n178 VSUBS 0.007112f
C249 B.n179 VSUBS 0.007112f
C250 B.n180 VSUBS 0.007112f
C251 B.n181 VSUBS 0.007112f
C252 B.n182 VSUBS 0.007112f
C253 B.n183 VSUBS 0.007112f
C254 B.n184 VSUBS 0.007112f
C255 B.n185 VSUBS 0.007112f
C256 B.n186 VSUBS 0.007112f
C257 B.n187 VSUBS 0.007112f
C258 B.n188 VSUBS 0.007112f
C259 B.n189 VSUBS 0.007112f
C260 B.n190 VSUBS 0.007112f
C261 B.n191 VSUBS 0.007112f
C262 B.n192 VSUBS 0.007112f
C263 B.n193 VSUBS 0.007112f
C264 B.n194 VSUBS 0.007112f
C265 B.n195 VSUBS 0.007112f
C266 B.n196 VSUBS 0.007112f
C267 B.n197 VSUBS 0.007112f
C268 B.n198 VSUBS 0.007112f
C269 B.n199 VSUBS 0.007112f
C270 B.n200 VSUBS 0.007112f
C271 B.n201 VSUBS 0.007112f
C272 B.n202 VSUBS 0.007112f
C273 B.n203 VSUBS 0.007112f
C274 B.n204 VSUBS 0.007112f
C275 B.n205 VSUBS 0.007112f
C276 B.n206 VSUBS 0.007112f
C277 B.n207 VSUBS 0.007112f
C278 B.n208 VSUBS 0.007112f
C279 B.n209 VSUBS 0.007112f
C280 B.n210 VSUBS 0.007112f
C281 B.n211 VSUBS 0.007112f
C282 B.n212 VSUBS 0.007112f
C283 B.n213 VSUBS 0.007112f
C284 B.n214 VSUBS 0.007112f
C285 B.n215 VSUBS 0.007112f
C286 B.n216 VSUBS 0.007112f
C287 B.n217 VSUBS 0.007112f
C288 B.n218 VSUBS 0.007112f
C289 B.n219 VSUBS 0.007112f
C290 B.n220 VSUBS 0.007112f
C291 B.n221 VSUBS 0.007112f
C292 B.n222 VSUBS 0.007112f
C293 B.n223 VSUBS 0.007112f
C294 B.n224 VSUBS 0.007112f
C295 B.n225 VSUBS 0.007112f
C296 B.n226 VSUBS 0.007112f
C297 B.n227 VSUBS 0.007112f
C298 B.n228 VSUBS 0.007112f
C299 B.n229 VSUBS 0.007112f
C300 B.n230 VSUBS 0.007112f
C301 B.n231 VSUBS 0.007112f
C302 B.n232 VSUBS 0.007112f
C303 B.n233 VSUBS 0.007112f
C304 B.n234 VSUBS 0.007112f
C305 B.n235 VSUBS 0.007112f
C306 B.n236 VSUBS 0.007112f
C307 B.n237 VSUBS 0.007112f
C308 B.n238 VSUBS 0.007112f
C309 B.n239 VSUBS 0.007112f
C310 B.n240 VSUBS 0.007112f
C311 B.n241 VSUBS 0.007112f
C312 B.n242 VSUBS 0.007112f
C313 B.n243 VSUBS 0.007112f
C314 B.n244 VSUBS 0.007112f
C315 B.n245 VSUBS 0.007112f
C316 B.n246 VSUBS 0.007112f
C317 B.n247 VSUBS 0.007112f
C318 B.n248 VSUBS 0.007112f
C319 B.n249 VSUBS 0.007112f
C320 B.n250 VSUBS 0.015773f
C321 B.n251 VSUBS 0.015773f
C322 B.n252 VSUBS 0.016648f
C323 B.n253 VSUBS 0.007112f
C324 B.n254 VSUBS 0.007112f
C325 B.n255 VSUBS 0.007112f
C326 B.n256 VSUBS 0.007112f
C327 B.n257 VSUBS 0.007112f
C328 B.n258 VSUBS 0.007112f
C329 B.n259 VSUBS 0.007112f
C330 B.n260 VSUBS 0.007112f
C331 B.n261 VSUBS 0.007112f
C332 B.n262 VSUBS 0.007112f
C333 B.n263 VSUBS 0.007112f
C334 B.n264 VSUBS 0.007112f
C335 B.n265 VSUBS 0.007112f
C336 B.n266 VSUBS 0.007112f
C337 B.n267 VSUBS 0.007112f
C338 B.n268 VSUBS 0.007112f
C339 B.n269 VSUBS 0.007112f
C340 B.n270 VSUBS 0.007112f
C341 B.n271 VSUBS 0.007112f
C342 B.n272 VSUBS 0.007112f
C343 B.n273 VSUBS 0.007112f
C344 B.n274 VSUBS 0.007112f
C345 B.n275 VSUBS 0.007112f
C346 B.n276 VSUBS 0.007112f
C347 B.n277 VSUBS 0.007112f
C348 B.n278 VSUBS 0.007112f
C349 B.n279 VSUBS 0.007112f
C350 B.n280 VSUBS 0.007112f
C351 B.n281 VSUBS 0.007112f
C352 B.n282 VSUBS 0.007112f
C353 B.n283 VSUBS 0.007112f
C354 B.n284 VSUBS 0.007112f
C355 B.n285 VSUBS 0.007112f
C356 B.n286 VSUBS 0.007112f
C357 B.n287 VSUBS 0.007112f
C358 B.n288 VSUBS 0.007112f
C359 B.n289 VSUBS 0.007112f
C360 B.n290 VSUBS 0.007112f
C361 B.n291 VSUBS 0.007112f
C362 B.n292 VSUBS 0.007112f
C363 B.n293 VSUBS 0.007112f
C364 B.n294 VSUBS 0.007112f
C365 B.n295 VSUBS 0.007112f
C366 B.n296 VSUBS 0.007112f
C367 B.n297 VSUBS 0.007112f
C368 B.n298 VSUBS 0.007112f
C369 B.n299 VSUBS 0.007112f
C370 B.n300 VSUBS 0.007112f
C371 B.n301 VSUBS 0.007112f
C372 B.n302 VSUBS 0.007112f
C373 B.n303 VSUBS 0.007112f
C374 B.n304 VSUBS 0.007112f
C375 B.n305 VSUBS 0.007112f
C376 B.n306 VSUBS 0.007112f
C377 B.n307 VSUBS 0.007112f
C378 B.n308 VSUBS 0.007112f
C379 B.n309 VSUBS 0.007112f
C380 B.n310 VSUBS 0.007112f
C381 B.n311 VSUBS 0.006693f
C382 B.n312 VSUBS 0.016477f
C383 B.n313 VSUBS 0.003974f
C384 B.n314 VSUBS 0.007112f
C385 B.n315 VSUBS 0.007112f
C386 B.n316 VSUBS 0.007112f
C387 B.n317 VSUBS 0.007112f
C388 B.n318 VSUBS 0.007112f
C389 B.n319 VSUBS 0.007112f
C390 B.n320 VSUBS 0.007112f
C391 B.n321 VSUBS 0.007112f
C392 B.n322 VSUBS 0.007112f
C393 B.n323 VSUBS 0.007112f
C394 B.n324 VSUBS 0.007112f
C395 B.n325 VSUBS 0.007112f
C396 B.t11 VSUBS 0.203322f
C397 B.t10 VSUBS 0.246865f
C398 B.t9 VSUBS 2.0694f
C399 B.n326 VSUBS 0.394251f
C400 B.n327 VSUBS 0.253562f
C401 B.n328 VSUBS 0.016477f
C402 B.n329 VSUBS 0.003974f
C403 B.n330 VSUBS 0.007112f
C404 B.n331 VSUBS 0.007112f
C405 B.n332 VSUBS 0.007112f
C406 B.n333 VSUBS 0.007112f
C407 B.n334 VSUBS 0.007112f
C408 B.n335 VSUBS 0.007112f
C409 B.n336 VSUBS 0.007112f
C410 B.n337 VSUBS 0.007112f
C411 B.n338 VSUBS 0.007112f
C412 B.n339 VSUBS 0.007112f
C413 B.n340 VSUBS 0.007112f
C414 B.n341 VSUBS 0.007112f
C415 B.n342 VSUBS 0.007112f
C416 B.n343 VSUBS 0.007112f
C417 B.n344 VSUBS 0.007112f
C418 B.n345 VSUBS 0.007112f
C419 B.n346 VSUBS 0.007112f
C420 B.n347 VSUBS 0.007112f
C421 B.n348 VSUBS 0.007112f
C422 B.n349 VSUBS 0.007112f
C423 B.n350 VSUBS 0.007112f
C424 B.n351 VSUBS 0.007112f
C425 B.n352 VSUBS 0.007112f
C426 B.n353 VSUBS 0.007112f
C427 B.n354 VSUBS 0.007112f
C428 B.n355 VSUBS 0.007112f
C429 B.n356 VSUBS 0.007112f
C430 B.n357 VSUBS 0.007112f
C431 B.n358 VSUBS 0.007112f
C432 B.n359 VSUBS 0.007112f
C433 B.n360 VSUBS 0.007112f
C434 B.n361 VSUBS 0.007112f
C435 B.n362 VSUBS 0.007112f
C436 B.n363 VSUBS 0.007112f
C437 B.n364 VSUBS 0.007112f
C438 B.n365 VSUBS 0.007112f
C439 B.n366 VSUBS 0.007112f
C440 B.n367 VSUBS 0.007112f
C441 B.n368 VSUBS 0.007112f
C442 B.n369 VSUBS 0.007112f
C443 B.n370 VSUBS 0.007112f
C444 B.n371 VSUBS 0.007112f
C445 B.n372 VSUBS 0.007112f
C446 B.n373 VSUBS 0.007112f
C447 B.n374 VSUBS 0.007112f
C448 B.n375 VSUBS 0.007112f
C449 B.n376 VSUBS 0.007112f
C450 B.n377 VSUBS 0.007112f
C451 B.n378 VSUBS 0.007112f
C452 B.n379 VSUBS 0.007112f
C453 B.n380 VSUBS 0.007112f
C454 B.n381 VSUBS 0.007112f
C455 B.n382 VSUBS 0.007112f
C456 B.n383 VSUBS 0.007112f
C457 B.n384 VSUBS 0.007112f
C458 B.n385 VSUBS 0.007112f
C459 B.n386 VSUBS 0.007112f
C460 B.n387 VSUBS 0.007112f
C461 B.n388 VSUBS 0.007112f
C462 B.n389 VSUBS 0.015773f
C463 B.n390 VSUBS 0.016648f
C464 B.n391 VSUBS 0.015773f
C465 B.n392 VSUBS 0.007112f
C466 B.n393 VSUBS 0.007112f
C467 B.n394 VSUBS 0.007112f
C468 B.n395 VSUBS 0.007112f
C469 B.n396 VSUBS 0.007112f
C470 B.n397 VSUBS 0.007112f
C471 B.n398 VSUBS 0.007112f
C472 B.n399 VSUBS 0.007112f
C473 B.n400 VSUBS 0.007112f
C474 B.n401 VSUBS 0.007112f
C475 B.n402 VSUBS 0.007112f
C476 B.n403 VSUBS 0.007112f
C477 B.n404 VSUBS 0.007112f
C478 B.n405 VSUBS 0.007112f
C479 B.n406 VSUBS 0.007112f
C480 B.n407 VSUBS 0.007112f
C481 B.n408 VSUBS 0.007112f
C482 B.n409 VSUBS 0.007112f
C483 B.n410 VSUBS 0.007112f
C484 B.n411 VSUBS 0.007112f
C485 B.n412 VSUBS 0.007112f
C486 B.n413 VSUBS 0.007112f
C487 B.n414 VSUBS 0.007112f
C488 B.n415 VSUBS 0.007112f
C489 B.n416 VSUBS 0.007112f
C490 B.n417 VSUBS 0.007112f
C491 B.n418 VSUBS 0.007112f
C492 B.n419 VSUBS 0.007112f
C493 B.n420 VSUBS 0.007112f
C494 B.n421 VSUBS 0.007112f
C495 B.n422 VSUBS 0.007112f
C496 B.n423 VSUBS 0.007112f
C497 B.n424 VSUBS 0.007112f
C498 B.n425 VSUBS 0.007112f
C499 B.n426 VSUBS 0.007112f
C500 B.n427 VSUBS 0.007112f
C501 B.n428 VSUBS 0.007112f
C502 B.n429 VSUBS 0.007112f
C503 B.n430 VSUBS 0.007112f
C504 B.n431 VSUBS 0.007112f
C505 B.n432 VSUBS 0.007112f
C506 B.n433 VSUBS 0.007112f
C507 B.n434 VSUBS 0.007112f
C508 B.n435 VSUBS 0.007112f
C509 B.n436 VSUBS 0.007112f
C510 B.n437 VSUBS 0.007112f
C511 B.n438 VSUBS 0.007112f
C512 B.n439 VSUBS 0.007112f
C513 B.n440 VSUBS 0.007112f
C514 B.n441 VSUBS 0.007112f
C515 B.n442 VSUBS 0.007112f
C516 B.n443 VSUBS 0.007112f
C517 B.n444 VSUBS 0.007112f
C518 B.n445 VSUBS 0.007112f
C519 B.n446 VSUBS 0.007112f
C520 B.n447 VSUBS 0.007112f
C521 B.n448 VSUBS 0.007112f
C522 B.n449 VSUBS 0.007112f
C523 B.n450 VSUBS 0.007112f
C524 B.n451 VSUBS 0.007112f
C525 B.n452 VSUBS 0.007112f
C526 B.n453 VSUBS 0.007112f
C527 B.n454 VSUBS 0.007112f
C528 B.n455 VSUBS 0.007112f
C529 B.n456 VSUBS 0.007112f
C530 B.n457 VSUBS 0.007112f
C531 B.n458 VSUBS 0.007112f
C532 B.n459 VSUBS 0.007112f
C533 B.n460 VSUBS 0.007112f
C534 B.n461 VSUBS 0.007112f
C535 B.n462 VSUBS 0.007112f
C536 B.n463 VSUBS 0.007112f
C537 B.n464 VSUBS 0.007112f
C538 B.n465 VSUBS 0.007112f
C539 B.n466 VSUBS 0.007112f
C540 B.n467 VSUBS 0.007112f
C541 B.n468 VSUBS 0.007112f
C542 B.n469 VSUBS 0.007112f
C543 B.n470 VSUBS 0.007112f
C544 B.n471 VSUBS 0.007112f
C545 B.n472 VSUBS 0.007112f
C546 B.n473 VSUBS 0.007112f
C547 B.n474 VSUBS 0.007112f
C548 B.n475 VSUBS 0.007112f
C549 B.n476 VSUBS 0.007112f
C550 B.n477 VSUBS 0.007112f
C551 B.n478 VSUBS 0.007112f
C552 B.n479 VSUBS 0.007112f
C553 B.n480 VSUBS 0.007112f
C554 B.n481 VSUBS 0.007112f
C555 B.n482 VSUBS 0.007112f
C556 B.n483 VSUBS 0.007112f
C557 B.n484 VSUBS 0.007112f
C558 B.n485 VSUBS 0.007112f
C559 B.n486 VSUBS 0.007112f
C560 B.n487 VSUBS 0.007112f
C561 B.n488 VSUBS 0.007112f
C562 B.n489 VSUBS 0.007112f
C563 B.n490 VSUBS 0.007112f
C564 B.n491 VSUBS 0.007112f
C565 B.n492 VSUBS 0.007112f
C566 B.n493 VSUBS 0.007112f
C567 B.n494 VSUBS 0.007112f
C568 B.n495 VSUBS 0.007112f
C569 B.n496 VSUBS 0.007112f
C570 B.n497 VSUBS 0.007112f
C571 B.n498 VSUBS 0.007112f
C572 B.n499 VSUBS 0.007112f
C573 B.n500 VSUBS 0.007112f
C574 B.n501 VSUBS 0.007112f
C575 B.n502 VSUBS 0.007112f
C576 B.n503 VSUBS 0.007112f
C577 B.n504 VSUBS 0.007112f
C578 B.n505 VSUBS 0.007112f
C579 B.n506 VSUBS 0.007112f
C580 B.n507 VSUBS 0.007112f
C581 B.n508 VSUBS 0.007112f
C582 B.n509 VSUBS 0.007112f
C583 B.n510 VSUBS 0.007112f
C584 B.n511 VSUBS 0.007112f
C585 B.n512 VSUBS 0.007112f
C586 B.n513 VSUBS 0.007112f
C587 B.n514 VSUBS 0.007112f
C588 B.n515 VSUBS 0.007112f
C589 B.n516 VSUBS 0.007112f
C590 B.n517 VSUBS 0.007112f
C591 B.n518 VSUBS 0.007112f
C592 B.n519 VSUBS 0.007112f
C593 B.n520 VSUBS 0.007112f
C594 B.n521 VSUBS 0.007112f
C595 B.n522 VSUBS 0.007112f
C596 B.n523 VSUBS 0.007112f
C597 B.n524 VSUBS 0.015773f
C598 B.n525 VSUBS 0.015773f
C599 B.n526 VSUBS 0.016648f
C600 B.n527 VSUBS 0.007112f
C601 B.n528 VSUBS 0.007112f
C602 B.n529 VSUBS 0.007112f
C603 B.n530 VSUBS 0.007112f
C604 B.n531 VSUBS 0.007112f
C605 B.n532 VSUBS 0.007112f
C606 B.n533 VSUBS 0.007112f
C607 B.n534 VSUBS 0.007112f
C608 B.n535 VSUBS 0.007112f
C609 B.n536 VSUBS 0.007112f
C610 B.n537 VSUBS 0.007112f
C611 B.n538 VSUBS 0.007112f
C612 B.n539 VSUBS 0.007112f
C613 B.n540 VSUBS 0.007112f
C614 B.n541 VSUBS 0.007112f
C615 B.n542 VSUBS 0.007112f
C616 B.n543 VSUBS 0.007112f
C617 B.n544 VSUBS 0.007112f
C618 B.n545 VSUBS 0.007112f
C619 B.n546 VSUBS 0.007112f
C620 B.n547 VSUBS 0.007112f
C621 B.n548 VSUBS 0.007112f
C622 B.n549 VSUBS 0.007112f
C623 B.n550 VSUBS 0.007112f
C624 B.n551 VSUBS 0.007112f
C625 B.n552 VSUBS 0.007112f
C626 B.n553 VSUBS 0.007112f
C627 B.n554 VSUBS 0.007112f
C628 B.n555 VSUBS 0.007112f
C629 B.n556 VSUBS 0.007112f
C630 B.n557 VSUBS 0.007112f
C631 B.n558 VSUBS 0.007112f
C632 B.n559 VSUBS 0.007112f
C633 B.n560 VSUBS 0.007112f
C634 B.n561 VSUBS 0.007112f
C635 B.n562 VSUBS 0.007112f
C636 B.n563 VSUBS 0.007112f
C637 B.n564 VSUBS 0.007112f
C638 B.n565 VSUBS 0.007112f
C639 B.n566 VSUBS 0.007112f
C640 B.n567 VSUBS 0.007112f
C641 B.n568 VSUBS 0.007112f
C642 B.n569 VSUBS 0.007112f
C643 B.n570 VSUBS 0.007112f
C644 B.n571 VSUBS 0.007112f
C645 B.n572 VSUBS 0.007112f
C646 B.n573 VSUBS 0.007112f
C647 B.n574 VSUBS 0.007112f
C648 B.n575 VSUBS 0.007112f
C649 B.n576 VSUBS 0.007112f
C650 B.n577 VSUBS 0.007112f
C651 B.n578 VSUBS 0.007112f
C652 B.n579 VSUBS 0.007112f
C653 B.n580 VSUBS 0.007112f
C654 B.n581 VSUBS 0.007112f
C655 B.n582 VSUBS 0.007112f
C656 B.n583 VSUBS 0.007112f
C657 B.n584 VSUBS 0.007112f
C658 B.n585 VSUBS 0.006693f
C659 B.n586 VSUBS 0.016477f
C660 B.n587 VSUBS 0.003974f
C661 B.n588 VSUBS 0.007112f
C662 B.n589 VSUBS 0.007112f
C663 B.n590 VSUBS 0.007112f
C664 B.n591 VSUBS 0.007112f
C665 B.n592 VSUBS 0.007112f
C666 B.n593 VSUBS 0.007112f
C667 B.n594 VSUBS 0.007112f
C668 B.n595 VSUBS 0.007112f
C669 B.n596 VSUBS 0.007112f
C670 B.n597 VSUBS 0.007112f
C671 B.n598 VSUBS 0.007112f
C672 B.n599 VSUBS 0.007112f
C673 B.n600 VSUBS 0.003974f
C674 B.n601 VSUBS 0.007112f
C675 B.n602 VSUBS 0.007112f
C676 B.n603 VSUBS 0.006693f
C677 B.n604 VSUBS 0.007112f
C678 B.n605 VSUBS 0.007112f
C679 B.n606 VSUBS 0.007112f
C680 B.n607 VSUBS 0.007112f
C681 B.n608 VSUBS 0.007112f
C682 B.n609 VSUBS 0.007112f
C683 B.n610 VSUBS 0.007112f
C684 B.n611 VSUBS 0.007112f
C685 B.n612 VSUBS 0.007112f
C686 B.n613 VSUBS 0.007112f
C687 B.n614 VSUBS 0.007112f
C688 B.n615 VSUBS 0.007112f
C689 B.n616 VSUBS 0.007112f
C690 B.n617 VSUBS 0.007112f
C691 B.n618 VSUBS 0.007112f
C692 B.n619 VSUBS 0.007112f
C693 B.n620 VSUBS 0.007112f
C694 B.n621 VSUBS 0.007112f
C695 B.n622 VSUBS 0.007112f
C696 B.n623 VSUBS 0.007112f
C697 B.n624 VSUBS 0.007112f
C698 B.n625 VSUBS 0.007112f
C699 B.n626 VSUBS 0.007112f
C700 B.n627 VSUBS 0.007112f
C701 B.n628 VSUBS 0.007112f
C702 B.n629 VSUBS 0.007112f
C703 B.n630 VSUBS 0.007112f
C704 B.n631 VSUBS 0.007112f
C705 B.n632 VSUBS 0.007112f
C706 B.n633 VSUBS 0.007112f
C707 B.n634 VSUBS 0.007112f
C708 B.n635 VSUBS 0.007112f
C709 B.n636 VSUBS 0.007112f
C710 B.n637 VSUBS 0.007112f
C711 B.n638 VSUBS 0.007112f
C712 B.n639 VSUBS 0.007112f
C713 B.n640 VSUBS 0.007112f
C714 B.n641 VSUBS 0.007112f
C715 B.n642 VSUBS 0.007112f
C716 B.n643 VSUBS 0.007112f
C717 B.n644 VSUBS 0.007112f
C718 B.n645 VSUBS 0.007112f
C719 B.n646 VSUBS 0.007112f
C720 B.n647 VSUBS 0.007112f
C721 B.n648 VSUBS 0.007112f
C722 B.n649 VSUBS 0.007112f
C723 B.n650 VSUBS 0.007112f
C724 B.n651 VSUBS 0.007112f
C725 B.n652 VSUBS 0.007112f
C726 B.n653 VSUBS 0.007112f
C727 B.n654 VSUBS 0.007112f
C728 B.n655 VSUBS 0.007112f
C729 B.n656 VSUBS 0.007112f
C730 B.n657 VSUBS 0.007112f
C731 B.n658 VSUBS 0.007112f
C732 B.n659 VSUBS 0.007112f
C733 B.n660 VSUBS 0.007112f
C734 B.n661 VSUBS 0.016648f
C735 B.n662 VSUBS 0.015773f
C736 B.n663 VSUBS 0.015773f
C737 B.n664 VSUBS 0.007112f
C738 B.n665 VSUBS 0.007112f
C739 B.n666 VSUBS 0.007112f
C740 B.n667 VSUBS 0.007112f
C741 B.n668 VSUBS 0.007112f
C742 B.n669 VSUBS 0.007112f
C743 B.n670 VSUBS 0.007112f
C744 B.n671 VSUBS 0.007112f
C745 B.n672 VSUBS 0.007112f
C746 B.n673 VSUBS 0.007112f
C747 B.n674 VSUBS 0.007112f
C748 B.n675 VSUBS 0.007112f
C749 B.n676 VSUBS 0.007112f
C750 B.n677 VSUBS 0.007112f
C751 B.n678 VSUBS 0.007112f
C752 B.n679 VSUBS 0.007112f
C753 B.n680 VSUBS 0.007112f
C754 B.n681 VSUBS 0.007112f
C755 B.n682 VSUBS 0.007112f
C756 B.n683 VSUBS 0.007112f
C757 B.n684 VSUBS 0.007112f
C758 B.n685 VSUBS 0.007112f
C759 B.n686 VSUBS 0.007112f
C760 B.n687 VSUBS 0.007112f
C761 B.n688 VSUBS 0.007112f
C762 B.n689 VSUBS 0.007112f
C763 B.n690 VSUBS 0.007112f
C764 B.n691 VSUBS 0.007112f
C765 B.n692 VSUBS 0.007112f
C766 B.n693 VSUBS 0.007112f
C767 B.n694 VSUBS 0.007112f
C768 B.n695 VSUBS 0.007112f
C769 B.n696 VSUBS 0.007112f
C770 B.n697 VSUBS 0.007112f
C771 B.n698 VSUBS 0.007112f
C772 B.n699 VSUBS 0.007112f
C773 B.n700 VSUBS 0.007112f
C774 B.n701 VSUBS 0.007112f
C775 B.n702 VSUBS 0.007112f
C776 B.n703 VSUBS 0.007112f
C777 B.n704 VSUBS 0.007112f
C778 B.n705 VSUBS 0.007112f
C779 B.n706 VSUBS 0.007112f
C780 B.n707 VSUBS 0.007112f
C781 B.n708 VSUBS 0.007112f
C782 B.n709 VSUBS 0.007112f
C783 B.n710 VSUBS 0.007112f
C784 B.n711 VSUBS 0.007112f
C785 B.n712 VSUBS 0.007112f
C786 B.n713 VSUBS 0.007112f
C787 B.n714 VSUBS 0.007112f
C788 B.n715 VSUBS 0.007112f
C789 B.n716 VSUBS 0.007112f
C790 B.n717 VSUBS 0.007112f
C791 B.n718 VSUBS 0.007112f
C792 B.n719 VSUBS 0.007112f
C793 B.n720 VSUBS 0.007112f
C794 B.n721 VSUBS 0.007112f
C795 B.n722 VSUBS 0.007112f
C796 B.n723 VSUBS 0.007112f
C797 B.n724 VSUBS 0.007112f
C798 B.n725 VSUBS 0.007112f
C799 B.n726 VSUBS 0.007112f
C800 B.n727 VSUBS 0.00928f
C801 B.n728 VSUBS 0.009886f
C802 B.n729 VSUBS 0.019659f
C803 VTAIL.n0 VSUBS 0.027795f
C804 VTAIL.n1 VSUBS 0.024816f
C805 VTAIL.n2 VSUBS 0.013335f
C806 VTAIL.n3 VSUBS 0.031519f
C807 VTAIL.n4 VSUBS 0.014119f
C808 VTAIL.n5 VSUBS 0.024816f
C809 VTAIL.n6 VSUBS 0.013335f
C810 VTAIL.n7 VSUBS 0.031519f
C811 VTAIL.n8 VSUBS 0.013727f
C812 VTAIL.n9 VSUBS 0.024816f
C813 VTAIL.n10 VSUBS 0.014119f
C814 VTAIL.n11 VSUBS 0.031519f
C815 VTAIL.n12 VSUBS 0.014119f
C816 VTAIL.n13 VSUBS 0.024816f
C817 VTAIL.n14 VSUBS 0.013335f
C818 VTAIL.n15 VSUBS 0.031519f
C819 VTAIL.n16 VSUBS 0.014119f
C820 VTAIL.n17 VSUBS 1.16491f
C821 VTAIL.n18 VSUBS 0.013335f
C822 VTAIL.t7 VSUBS 0.067883f
C823 VTAIL.n19 VSUBS 0.189834f
C824 VTAIL.n20 VSUBS 0.02371f
C825 VTAIL.n21 VSUBS 0.023639f
C826 VTAIL.n22 VSUBS 0.031519f
C827 VTAIL.n23 VSUBS 0.014119f
C828 VTAIL.n24 VSUBS 0.013335f
C829 VTAIL.n25 VSUBS 0.024816f
C830 VTAIL.n26 VSUBS 0.024816f
C831 VTAIL.n27 VSUBS 0.013335f
C832 VTAIL.n28 VSUBS 0.014119f
C833 VTAIL.n29 VSUBS 0.031519f
C834 VTAIL.n30 VSUBS 0.031519f
C835 VTAIL.n31 VSUBS 0.014119f
C836 VTAIL.n32 VSUBS 0.013335f
C837 VTAIL.n33 VSUBS 0.024816f
C838 VTAIL.n34 VSUBS 0.024816f
C839 VTAIL.n35 VSUBS 0.013335f
C840 VTAIL.n36 VSUBS 0.013335f
C841 VTAIL.n37 VSUBS 0.014119f
C842 VTAIL.n38 VSUBS 0.031519f
C843 VTAIL.n39 VSUBS 0.031519f
C844 VTAIL.n40 VSUBS 0.031519f
C845 VTAIL.n41 VSUBS 0.013727f
C846 VTAIL.n42 VSUBS 0.013335f
C847 VTAIL.n43 VSUBS 0.024816f
C848 VTAIL.n44 VSUBS 0.024816f
C849 VTAIL.n45 VSUBS 0.013335f
C850 VTAIL.n46 VSUBS 0.014119f
C851 VTAIL.n47 VSUBS 0.031519f
C852 VTAIL.n48 VSUBS 0.031519f
C853 VTAIL.n49 VSUBS 0.014119f
C854 VTAIL.n50 VSUBS 0.013335f
C855 VTAIL.n51 VSUBS 0.024816f
C856 VTAIL.n52 VSUBS 0.024816f
C857 VTAIL.n53 VSUBS 0.013335f
C858 VTAIL.n54 VSUBS 0.014119f
C859 VTAIL.n55 VSUBS 0.031519f
C860 VTAIL.n56 VSUBS 0.078101f
C861 VTAIL.n57 VSUBS 0.014119f
C862 VTAIL.n58 VSUBS 0.013335f
C863 VTAIL.n59 VSUBS 0.060751f
C864 VTAIL.n60 VSUBS 0.039457f
C865 VTAIL.n61 VSUBS 0.207334f
C866 VTAIL.n62 VSUBS 0.027795f
C867 VTAIL.n63 VSUBS 0.024816f
C868 VTAIL.n64 VSUBS 0.013335f
C869 VTAIL.n65 VSUBS 0.031519f
C870 VTAIL.n66 VSUBS 0.014119f
C871 VTAIL.n67 VSUBS 0.024816f
C872 VTAIL.n68 VSUBS 0.013335f
C873 VTAIL.n69 VSUBS 0.031519f
C874 VTAIL.n70 VSUBS 0.013727f
C875 VTAIL.n71 VSUBS 0.024816f
C876 VTAIL.n72 VSUBS 0.014119f
C877 VTAIL.n73 VSUBS 0.031519f
C878 VTAIL.n74 VSUBS 0.014119f
C879 VTAIL.n75 VSUBS 0.024816f
C880 VTAIL.n76 VSUBS 0.013335f
C881 VTAIL.n77 VSUBS 0.031519f
C882 VTAIL.n78 VSUBS 0.014119f
C883 VTAIL.n79 VSUBS 1.16491f
C884 VTAIL.n80 VSUBS 0.013335f
C885 VTAIL.t1 VSUBS 0.067883f
C886 VTAIL.n81 VSUBS 0.189834f
C887 VTAIL.n82 VSUBS 0.02371f
C888 VTAIL.n83 VSUBS 0.023639f
C889 VTAIL.n84 VSUBS 0.031519f
C890 VTAIL.n85 VSUBS 0.014119f
C891 VTAIL.n86 VSUBS 0.013335f
C892 VTAIL.n87 VSUBS 0.024816f
C893 VTAIL.n88 VSUBS 0.024816f
C894 VTAIL.n89 VSUBS 0.013335f
C895 VTAIL.n90 VSUBS 0.014119f
C896 VTAIL.n91 VSUBS 0.031519f
C897 VTAIL.n92 VSUBS 0.031519f
C898 VTAIL.n93 VSUBS 0.014119f
C899 VTAIL.n94 VSUBS 0.013335f
C900 VTAIL.n95 VSUBS 0.024816f
C901 VTAIL.n96 VSUBS 0.024816f
C902 VTAIL.n97 VSUBS 0.013335f
C903 VTAIL.n98 VSUBS 0.013335f
C904 VTAIL.n99 VSUBS 0.014119f
C905 VTAIL.n100 VSUBS 0.031519f
C906 VTAIL.n101 VSUBS 0.031519f
C907 VTAIL.n102 VSUBS 0.031519f
C908 VTAIL.n103 VSUBS 0.013727f
C909 VTAIL.n104 VSUBS 0.013335f
C910 VTAIL.n105 VSUBS 0.024816f
C911 VTAIL.n106 VSUBS 0.024816f
C912 VTAIL.n107 VSUBS 0.013335f
C913 VTAIL.n108 VSUBS 0.014119f
C914 VTAIL.n109 VSUBS 0.031519f
C915 VTAIL.n110 VSUBS 0.031519f
C916 VTAIL.n111 VSUBS 0.014119f
C917 VTAIL.n112 VSUBS 0.013335f
C918 VTAIL.n113 VSUBS 0.024816f
C919 VTAIL.n114 VSUBS 0.024816f
C920 VTAIL.n115 VSUBS 0.013335f
C921 VTAIL.n116 VSUBS 0.014119f
C922 VTAIL.n117 VSUBS 0.031519f
C923 VTAIL.n118 VSUBS 0.078101f
C924 VTAIL.n119 VSUBS 0.014119f
C925 VTAIL.n120 VSUBS 0.013335f
C926 VTAIL.n121 VSUBS 0.060751f
C927 VTAIL.n122 VSUBS 0.039457f
C928 VTAIL.n123 VSUBS 0.344683f
C929 VTAIL.n124 VSUBS 0.027795f
C930 VTAIL.n125 VSUBS 0.024816f
C931 VTAIL.n126 VSUBS 0.013335f
C932 VTAIL.n127 VSUBS 0.031519f
C933 VTAIL.n128 VSUBS 0.014119f
C934 VTAIL.n129 VSUBS 0.024816f
C935 VTAIL.n130 VSUBS 0.013335f
C936 VTAIL.n131 VSUBS 0.031519f
C937 VTAIL.n132 VSUBS 0.013727f
C938 VTAIL.n133 VSUBS 0.024816f
C939 VTAIL.n134 VSUBS 0.014119f
C940 VTAIL.n135 VSUBS 0.031519f
C941 VTAIL.n136 VSUBS 0.014119f
C942 VTAIL.n137 VSUBS 0.024816f
C943 VTAIL.n138 VSUBS 0.013335f
C944 VTAIL.n139 VSUBS 0.031519f
C945 VTAIL.n140 VSUBS 0.014119f
C946 VTAIL.n141 VSUBS 1.16491f
C947 VTAIL.n142 VSUBS 0.013335f
C948 VTAIL.t0 VSUBS 0.067883f
C949 VTAIL.n143 VSUBS 0.189834f
C950 VTAIL.n144 VSUBS 0.02371f
C951 VTAIL.n145 VSUBS 0.023639f
C952 VTAIL.n146 VSUBS 0.031519f
C953 VTAIL.n147 VSUBS 0.014119f
C954 VTAIL.n148 VSUBS 0.013335f
C955 VTAIL.n149 VSUBS 0.024816f
C956 VTAIL.n150 VSUBS 0.024816f
C957 VTAIL.n151 VSUBS 0.013335f
C958 VTAIL.n152 VSUBS 0.014119f
C959 VTAIL.n153 VSUBS 0.031519f
C960 VTAIL.n154 VSUBS 0.031519f
C961 VTAIL.n155 VSUBS 0.014119f
C962 VTAIL.n156 VSUBS 0.013335f
C963 VTAIL.n157 VSUBS 0.024816f
C964 VTAIL.n158 VSUBS 0.024816f
C965 VTAIL.n159 VSUBS 0.013335f
C966 VTAIL.n160 VSUBS 0.013335f
C967 VTAIL.n161 VSUBS 0.014119f
C968 VTAIL.n162 VSUBS 0.031519f
C969 VTAIL.n163 VSUBS 0.031519f
C970 VTAIL.n164 VSUBS 0.031519f
C971 VTAIL.n165 VSUBS 0.013727f
C972 VTAIL.n166 VSUBS 0.013335f
C973 VTAIL.n167 VSUBS 0.024816f
C974 VTAIL.n168 VSUBS 0.024816f
C975 VTAIL.n169 VSUBS 0.013335f
C976 VTAIL.n170 VSUBS 0.014119f
C977 VTAIL.n171 VSUBS 0.031519f
C978 VTAIL.n172 VSUBS 0.031519f
C979 VTAIL.n173 VSUBS 0.014119f
C980 VTAIL.n174 VSUBS 0.013335f
C981 VTAIL.n175 VSUBS 0.024816f
C982 VTAIL.n176 VSUBS 0.024816f
C983 VTAIL.n177 VSUBS 0.013335f
C984 VTAIL.n178 VSUBS 0.014119f
C985 VTAIL.n179 VSUBS 0.031519f
C986 VTAIL.n180 VSUBS 0.078101f
C987 VTAIL.n181 VSUBS 0.014119f
C988 VTAIL.n182 VSUBS 0.013335f
C989 VTAIL.n183 VSUBS 0.060751f
C990 VTAIL.n184 VSUBS 0.039457f
C991 VTAIL.n185 VSUBS 1.72094f
C992 VTAIL.n186 VSUBS 0.027795f
C993 VTAIL.n187 VSUBS 0.024816f
C994 VTAIL.n188 VSUBS 0.013335f
C995 VTAIL.n189 VSUBS 0.031519f
C996 VTAIL.n190 VSUBS 0.014119f
C997 VTAIL.n191 VSUBS 0.024816f
C998 VTAIL.n192 VSUBS 0.013335f
C999 VTAIL.n193 VSUBS 0.031519f
C1000 VTAIL.n194 VSUBS 0.013727f
C1001 VTAIL.n195 VSUBS 0.024816f
C1002 VTAIL.n196 VSUBS 0.013727f
C1003 VTAIL.n197 VSUBS 0.013335f
C1004 VTAIL.n198 VSUBS 0.031519f
C1005 VTAIL.n199 VSUBS 0.031519f
C1006 VTAIL.n200 VSUBS 0.014119f
C1007 VTAIL.n201 VSUBS 0.024816f
C1008 VTAIL.n202 VSUBS 0.013335f
C1009 VTAIL.n203 VSUBS 0.031519f
C1010 VTAIL.n204 VSUBS 0.014119f
C1011 VTAIL.n205 VSUBS 1.16491f
C1012 VTAIL.n206 VSUBS 0.013335f
C1013 VTAIL.t6 VSUBS 0.067883f
C1014 VTAIL.n207 VSUBS 0.189834f
C1015 VTAIL.n208 VSUBS 0.02371f
C1016 VTAIL.n209 VSUBS 0.023639f
C1017 VTAIL.n210 VSUBS 0.031519f
C1018 VTAIL.n211 VSUBS 0.014119f
C1019 VTAIL.n212 VSUBS 0.013335f
C1020 VTAIL.n213 VSUBS 0.024816f
C1021 VTAIL.n214 VSUBS 0.024816f
C1022 VTAIL.n215 VSUBS 0.013335f
C1023 VTAIL.n216 VSUBS 0.014119f
C1024 VTAIL.n217 VSUBS 0.031519f
C1025 VTAIL.n218 VSUBS 0.031519f
C1026 VTAIL.n219 VSUBS 0.014119f
C1027 VTAIL.n220 VSUBS 0.013335f
C1028 VTAIL.n221 VSUBS 0.024816f
C1029 VTAIL.n222 VSUBS 0.024816f
C1030 VTAIL.n223 VSUBS 0.013335f
C1031 VTAIL.n224 VSUBS 0.014119f
C1032 VTAIL.n225 VSUBS 0.031519f
C1033 VTAIL.n226 VSUBS 0.031519f
C1034 VTAIL.n227 VSUBS 0.014119f
C1035 VTAIL.n228 VSUBS 0.013335f
C1036 VTAIL.n229 VSUBS 0.024816f
C1037 VTAIL.n230 VSUBS 0.024816f
C1038 VTAIL.n231 VSUBS 0.013335f
C1039 VTAIL.n232 VSUBS 0.014119f
C1040 VTAIL.n233 VSUBS 0.031519f
C1041 VTAIL.n234 VSUBS 0.031519f
C1042 VTAIL.n235 VSUBS 0.014119f
C1043 VTAIL.n236 VSUBS 0.013335f
C1044 VTAIL.n237 VSUBS 0.024816f
C1045 VTAIL.n238 VSUBS 0.024816f
C1046 VTAIL.n239 VSUBS 0.013335f
C1047 VTAIL.n240 VSUBS 0.014119f
C1048 VTAIL.n241 VSUBS 0.031519f
C1049 VTAIL.n242 VSUBS 0.078101f
C1050 VTAIL.n243 VSUBS 0.014119f
C1051 VTAIL.n244 VSUBS 0.013335f
C1052 VTAIL.n245 VSUBS 0.060751f
C1053 VTAIL.n246 VSUBS 0.039457f
C1054 VTAIL.n247 VSUBS 1.72094f
C1055 VTAIL.n248 VSUBS 0.027795f
C1056 VTAIL.n249 VSUBS 0.024816f
C1057 VTAIL.n250 VSUBS 0.013335f
C1058 VTAIL.n251 VSUBS 0.031519f
C1059 VTAIL.n252 VSUBS 0.014119f
C1060 VTAIL.n253 VSUBS 0.024816f
C1061 VTAIL.n254 VSUBS 0.013335f
C1062 VTAIL.n255 VSUBS 0.031519f
C1063 VTAIL.n256 VSUBS 0.013727f
C1064 VTAIL.n257 VSUBS 0.024816f
C1065 VTAIL.n258 VSUBS 0.013727f
C1066 VTAIL.n259 VSUBS 0.013335f
C1067 VTAIL.n260 VSUBS 0.031519f
C1068 VTAIL.n261 VSUBS 0.031519f
C1069 VTAIL.n262 VSUBS 0.014119f
C1070 VTAIL.n263 VSUBS 0.024816f
C1071 VTAIL.n264 VSUBS 0.013335f
C1072 VTAIL.n265 VSUBS 0.031519f
C1073 VTAIL.n266 VSUBS 0.014119f
C1074 VTAIL.n267 VSUBS 1.16491f
C1075 VTAIL.n268 VSUBS 0.013335f
C1076 VTAIL.t5 VSUBS 0.067883f
C1077 VTAIL.n269 VSUBS 0.189834f
C1078 VTAIL.n270 VSUBS 0.02371f
C1079 VTAIL.n271 VSUBS 0.023639f
C1080 VTAIL.n272 VSUBS 0.031519f
C1081 VTAIL.n273 VSUBS 0.014119f
C1082 VTAIL.n274 VSUBS 0.013335f
C1083 VTAIL.n275 VSUBS 0.024816f
C1084 VTAIL.n276 VSUBS 0.024816f
C1085 VTAIL.n277 VSUBS 0.013335f
C1086 VTAIL.n278 VSUBS 0.014119f
C1087 VTAIL.n279 VSUBS 0.031519f
C1088 VTAIL.n280 VSUBS 0.031519f
C1089 VTAIL.n281 VSUBS 0.014119f
C1090 VTAIL.n282 VSUBS 0.013335f
C1091 VTAIL.n283 VSUBS 0.024816f
C1092 VTAIL.n284 VSUBS 0.024816f
C1093 VTAIL.n285 VSUBS 0.013335f
C1094 VTAIL.n286 VSUBS 0.014119f
C1095 VTAIL.n287 VSUBS 0.031519f
C1096 VTAIL.n288 VSUBS 0.031519f
C1097 VTAIL.n289 VSUBS 0.014119f
C1098 VTAIL.n290 VSUBS 0.013335f
C1099 VTAIL.n291 VSUBS 0.024816f
C1100 VTAIL.n292 VSUBS 0.024816f
C1101 VTAIL.n293 VSUBS 0.013335f
C1102 VTAIL.n294 VSUBS 0.014119f
C1103 VTAIL.n295 VSUBS 0.031519f
C1104 VTAIL.n296 VSUBS 0.031519f
C1105 VTAIL.n297 VSUBS 0.014119f
C1106 VTAIL.n298 VSUBS 0.013335f
C1107 VTAIL.n299 VSUBS 0.024816f
C1108 VTAIL.n300 VSUBS 0.024816f
C1109 VTAIL.n301 VSUBS 0.013335f
C1110 VTAIL.n302 VSUBS 0.014119f
C1111 VTAIL.n303 VSUBS 0.031519f
C1112 VTAIL.n304 VSUBS 0.078101f
C1113 VTAIL.n305 VSUBS 0.014119f
C1114 VTAIL.n306 VSUBS 0.013335f
C1115 VTAIL.n307 VSUBS 0.060751f
C1116 VTAIL.n308 VSUBS 0.039457f
C1117 VTAIL.n309 VSUBS 0.344683f
C1118 VTAIL.n310 VSUBS 0.027795f
C1119 VTAIL.n311 VSUBS 0.024816f
C1120 VTAIL.n312 VSUBS 0.013335f
C1121 VTAIL.n313 VSUBS 0.031519f
C1122 VTAIL.n314 VSUBS 0.014119f
C1123 VTAIL.n315 VSUBS 0.024816f
C1124 VTAIL.n316 VSUBS 0.013335f
C1125 VTAIL.n317 VSUBS 0.031519f
C1126 VTAIL.n318 VSUBS 0.013727f
C1127 VTAIL.n319 VSUBS 0.024816f
C1128 VTAIL.n320 VSUBS 0.013727f
C1129 VTAIL.n321 VSUBS 0.013335f
C1130 VTAIL.n322 VSUBS 0.031519f
C1131 VTAIL.n323 VSUBS 0.031519f
C1132 VTAIL.n324 VSUBS 0.014119f
C1133 VTAIL.n325 VSUBS 0.024816f
C1134 VTAIL.n326 VSUBS 0.013335f
C1135 VTAIL.n327 VSUBS 0.031519f
C1136 VTAIL.n328 VSUBS 0.014119f
C1137 VTAIL.n329 VSUBS 1.16491f
C1138 VTAIL.n330 VSUBS 0.013335f
C1139 VTAIL.t3 VSUBS 0.067883f
C1140 VTAIL.n331 VSUBS 0.189834f
C1141 VTAIL.n332 VSUBS 0.02371f
C1142 VTAIL.n333 VSUBS 0.023639f
C1143 VTAIL.n334 VSUBS 0.031519f
C1144 VTAIL.n335 VSUBS 0.014119f
C1145 VTAIL.n336 VSUBS 0.013335f
C1146 VTAIL.n337 VSUBS 0.024816f
C1147 VTAIL.n338 VSUBS 0.024816f
C1148 VTAIL.n339 VSUBS 0.013335f
C1149 VTAIL.n340 VSUBS 0.014119f
C1150 VTAIL.n341 VSUBS 0.031519f
C1151 VTAIL.n342 VSUBS 0.031519f
C1152 VTAIL.n343 VSUBS 0.014119f
C1153 VTAIL.n344 VSUBS 0.013335f
C1154 VTAIL.n345 VSUBS 0.024816f
C1155 VTAIL.n346 VSUBS 0.024816f
C1156 VTAIL.n347 VSUBS 0.013335f
C1157 VTAIL.n348 VSUBS 0.014119f
C1158 VTAIL.n349 VSUBS 0.031519f
C1159 VTAIL.n350 VSUBS 0.031519f
C1160 VTAIL.n351 VSUBS 0.014119f
C1161 VTAIL.n352 VSUBS 0.013335f
C1162 VTAIL.n353 VSUBS 0.024816f
C1163 VTAIL.n354 VSUBS 0.024816f
C1164 VTAIL.n355 VSUBS 0.013335f
C1165 VTAIL.n356 VSUBS 0.014119f
C1166 VTAIL.n357 VSUBS 0.031519f
C1167 VTAIL.n358 VSUBS 0.031519f
C1168 VTAIL.n359 VSUBS 0.014119f
C1169 VTAIL.n360 VSUBS 0.013335f
C1170 VTAIL.n361 VSUBS 0.024816f
C1171 VTAIL.n362 VSUBS 0.024816f
C1172 VTAIL.n363 VSUBS 0.013335f
C1173 VTAIL.n364 VSUBS 0.014119f
C1174 VTAIL.n365 VSUBS 0.031519f
C1175 VTAIL.n366 VSUBS 0.078101f
C1176 VTAIL.n367 VSUBS 0.014119f
C1177 VTAIL.n368 VSUBS 0.013335f
C1178 VTAIL.n369 VSUBS 0.060751f
C1179 VTAIL.n370 VSUBS 0.039457f
C1180 VTAIL.n371 VSUBS 0.344683f
C1181 VTAIL.n372 VSUBS 0.027795f
C1182 VTAIL.n373 VSUBS 0.024816f
C1183 VTAIL.n374 VSUBS 0.013335f
C1184 VTAIL.n375 VSUBS 0.031519f
C1185 VTAIL.n376 VSUBS 0.014119f
C1186 VTAIL.n377 VSUBS 0.024816f
C1187 VTAIL.n378 VSUBS 0.013335f
C1188 VTAIL.n379 VSUBS 0.031519f
C1189 VTAIL.n380 VSUBS 0.013727f
C1190 VTAIL.n381 VSUBS 0.024816f
C1191 VTAIL.n382 VSUBS 0.013727f
C1192 VTAIL.n383 VSUBS 0.013335f
C1193 VTAIL.n384 VSUBS 0.031519f
C1194 VTAIL.n385 VSUBS 0.031519f
C1195 VTAIL.n386 VSUBS 0.014119f
C1196 VTAIL.n387 VSUBS 0.024816f
C1197 VTAIL.n388 VSUBS 0.013335f
C1198 VTAIL.n389 VSUBS 0.031519f
C1199 VTAIL.n390 VSUBS 0.014119f
C1200 VTAIL.n391 VSUBS 1.16491f
C1201 VTAIL.n392 VSUBS 0.013335f
C1202 VTAIL.t2 VSUBS 0.067883f
C1203 VTAIL.n393 VSUBS 0.189834f
C1204 VTAIL.n394 VSUBS 0.02371f
C1205 VTAIL.n395 VSUBS 0.023639f
C1206 VTAIL.n396 VSUBS 0.031519f
C1207 VTAIL.n397 VSUBS 0.014119f
C1208 VTAIL.n398 VSUBS 0.013335f
C1209 VTAIL.n399 VSUBS 0.024816f
C1210 VTAIL.n400 VSUBS 0.024816f
C1211 VTAIL.n401 VSUBS 0.013335f
C1212 VTAIL.n402 VSUBS 0.014119f
C1213 VTAIL.n403 VSUBS 0.031519f
C1214 VTAIL.n404 VSUBS 0.031519f
C1215 VTAIL.n405 VSUBS 0.014119f
C1216 VTAIL.n406 VSUBS 0.013335f
C1217 VTAIL.n407 VSUBS 0.024816f
C1218 VTAIL.n408 VSUBS 0.024816f
C1219 VTAIL.n409 VSUBS 0.013335f
C1220 VTAIL.n410 VSUBS 0.014119f
C1221 VTAIL.n411 VSUBS 0.031519f
C1222 VTAIL.n412 VSUBS 0.031519f
C1223 VTAIL.n413 VSUBS 0.014119f
C1224 VTAIL.n414 VSUBS 0.013335f
C1225 VTAIL.n415 VSUBS 0.024816f
C1226 VTAIL.n416 VSUBS 0.024816f
C1227 VTAIL.n417 VSUBS 0.013335f
C1228 VTAIL.n418 VSUBS 0.014119f
C1229 VTAIL.n419 VSUBS 0.031519f
C1230 VTAIL.n420 VSUBS 0.031519f
C1231 VTAIL.n421 VSUBS 0.014119f
C1232 VTAIL.n422 VSUBS 0.013335f
C1233 VTAIL.n423 VSUBS 0.024816f
C1234 VTAIL.n424 VSUBS 0.024816f
C1235 VTAIL.n425 VSUBS 0.013335f
C1236 VTAIL.n426 VSUBS 0.014119f
C1237 VTAIL.n427 VSUBS 0.031519f
C1238 VTAIL.n428 VSUBS 0.078101f
C1239 VTAIL.n429 VSUBS 0.014119f
C1240 VTAIL.n430 VSUBS 0.013335f
C1241 VTAIL.n431 VSUBS 0.060751f
C1242 VTAIL.n432 VSUBS 0.039457f
C1243 VTAIL.n433 VSUBS 1.72094f
C1244 VTAIL.n434 VSUBS 0.027795f
C1245 VTAIL.n435 VSUBS 0.024816f
C1246 VTAIL.n436 VSUBS 0.013335f
C1247 VTAIL.n437 VSUBS 0.031519f
C1248 VTAIL.n438 VSUBS 0.014119f
C1249 VTAIL.n439 VSUBS 0.024816f
C1250 VTAIL.n440 VSUBS 0.013335f
C1251 VTAIL.n441 VSUBS 0.031519f
C1252 VTAIL.n442 VSUBS 0.013727f
C1253 VTAIL.n443 VSUBS 0.024816f
C1254 VTAIL.n444 VSUBS 0.014119f
C1255 VTAIL.n445 VSUBS 0.031519f
C1256 VTAIL.n446 VSUBS 0.014119f
C1257 VTAIL.n447 VSUBS 0.024816f
C1258 VTAIL.n448 VSUBS 0.013335f
C1259 VTAIL.n449 VSUBS 0.031519f
C1260 VTAIL.n450 VSUBS 0.014119f
C1261 VTAIL.n451 VSUBS 1.16491f
C1262 VTAIL.n452 VSUBS 0.013335f
C1263 VTAIL.t4 VSUBS 0.067883f
C1264 VTAIL.n453 VSUBS 0.189834f
C1265 VTAIL.n454 VSUBS 0.02371f
C1266 VTAIL.n455 VSUBS 0.023639f
C1267 VTAIL.n456 VSUBS 0.031519f
C1268 VTAIL.n457 VSUBS 0.014119f
C1269 VTAIL.n458 VSUBS 0.013335f
C1270 VTAIL.n459 VSUBS 0.024816f
C1271 VTAIL.n460 VSUBS 0.024816f
C1272 VTAIL.n461 VSUBS 0.013335f
C1273 VTAIL.n462 VSUBS 0.014119f
C1274 VTAIL.n463 VSUBS 0.031519f
C1275 VTAIL.n464 VSUBS 0.031519f
C1276 VTAIL.n465 VSUBS 0.014119f
C1277 VTAIL.n466 VSUBS 0.013335f
C1278 VTAIL.n467 VSUBS 0.024816f
C1279 VTAIL.n468 VSUBS 0.024816f
C1280 VTAIL.n469 VSUBS 0.013335f
C1281 VTAIL.n470 VSUBS 0.013335f
C1282 VTAIL.n471 VSUBS 0.014119f
C1283 VTAIL.n472 VSUBS 0.031519f
C1284 VTAIL.n473 VSUBS 0.031519f
C1285 VTAIL.n474 VSUBS 0.031519f
C1286 VTAIL.n475 VSUBS 0.013727f
C1287 VTAIL.n476 VSUBS 0.013335f
C1288 VTAIL.n477 VSUBS 0.024816f
C1289 VTAIL.n478 VSUBS 0.024816f
C1290 VTAIL.n479 VSUBS 0.013335f
C1291 VTAIL.n480 VSUBS 0.014119f
C1292 VTAIL.n481 VSUBS 0.031519f
C1293 VTAIL.n482 VSUBS 0.031519f
C1294 VTAIL.n483 VSUBS 0.014119f
C1295 VTAIL.n484 VSUBS 0.013335f
C1296 VTAIL.n485 VSUBS 0.024816f
C1297 VTAIL.n486 VSUBS 0.024816f
C1298 VTAIL.n487 VSUBS 0.013335f
C1299 VTAIL.n488 VSUBS 0.014119f
C1300 VTAIL.n489 VSUBS 0.031519f
C1301 VTAIL.n490 VSUBS 0.078101f
C1302 VTAIL.n491 VSUBS 0.014119f
C1303 VTAIL.n492 VSUBS 0.013335f
C1304 VTAIL.n493 VSUBS 0.060751f
C1305 VTAIL.n494 VSUBS 0.039457f
C1306 VTAIL.n495 VSUBS 1.57429f
C1307 VDD2.t2 VSUBS 0.247749f
C1308 VDD2.t3 VSUBS 0.247749f
C1309 VDD2.n0 VSUBS 2.66605f
C1310 VDD2.t1 VSUBS 0.247749f
C1311 VDD2.t0 VSUBS 0.247749f
C1312 VDD2.n1 VSUBS 1.92571f
C1313 VDD2.n2 VSUBS 4.59938f
C1314 VN.t3 VSUBS 3.65108f
C1315 VN.t0 VSUBS 3.66739f
C1316 VN.n0 VSUBS 2.17794f
C1317 VN.t1 VSUBS 3.65108f
C1318 VN.t2 VSUBS 3.66739f
C1319 VN.n1 VSUBS 3.95532f
.ends

