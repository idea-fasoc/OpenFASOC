* NGSPICE file created from diff_pair_sample_1024.ext - technology: sky130A

.subckt diff_pair_sample_1024 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t6 VN.t0 VDD2.t0 w_n2560_n4264# sky130_fd_pr__pfet_01v8 ad=6.4272 pd=33.74 as=2.7192 ps=16.81 w=16.48 l=2.32
X1 VTAIL.t5 VN.t1 VDD2.t1 w_n2560_n4264# sky130_fd_pr__pfet_01v8 ad=6.4272 pd=33.74 as=2.7192 ps=16.81 w=16.48 l=2.32
X2 VDD1.t3 VP.t0 VTAIL.t2 w_n2560_n4264# sky130_fd_pr__pfet_01v8 ad=2.7192 pd=16.81 as=6.4272 ps=33.74 w=16.48 l=2.32
X3 B.t11 B.t9 B.t10 w_n2560_n4264# sky130_fd_pr__pfet_01v8 ad=6.4272 pd=33.74 as=0 ps=0 w=16.48 l=2.32
X4 VTAIL.t7 VP.t1 VDD1.t2 w_n2560_n4264# sky130_fd_pr__pfet_01v8 ad=6.4272 pd=33.74 as=2.7192 ps=16.81 w=16.48 l=2.32
X5 VDD2.t2 VN.t2 VTAIL.t4 w_n2560_n4264# sky130_fd_pr__pfet_01v8 ad=2.7192 pd=16.81 as=6.4272 ps=33.74 w=16.48 l=2.32
X6 B.t8 B.t6 B.t7 w_n2560_n4264# sky130_fd_pr__pfet_01v8 ad=6.4272 pd=33.74 as=0 ps=0 w=16.48 l=2.32
X7 VTAIL.t1 VP.t2 VDD1.t1 w_n2560_n4264# sky130_fd_pr__pfet_01v8 ad=6.4272 pd=33.74 as=2.7192 ps=16.81 w=16.48 l=2.32
X8 VDD1.t0 VP.t3 VTAIL.t0 w_n2560_n4264# sky130_fd_pr__pfet_01v8 ad=2.7192 pd=16.81 as=6.4272 ps=33.74 w=16.48 l=2.32
X9 B.t5 B.t3 B.t4 w_n2560_n4264# sky130_fd_pr__pfet_01v8 ad=6.4272 pd=33.74 as=0 ps=0 w=16.48 l=2.32
X10 B.t2 B.t0 B.t1 w_n2560_n4264# sky130_fd_pr__pfet_01v8 ad=6.4272 pd=33.74 as=0 ps=0 w=16.48 l=2.32
X11 VDD2.t3 VN.t3 VTAIL.t3 w_n2560_n4264# sky130_fd_pr__pfet_01v8 ad=2.7192 pd=16.81 as=6.4272 ps=33.74 w=16.48 l=2.32
R0 VN.n0 VN.t1 207.739
R1 VN.n1 VN.t2 207.739
R2 VN.n0 VN.t3 207.083
R3 VN.n1 VN.t0 207.083
R4 VN VN.n1 54.6313
R5 VN VN.n0 5.49868
R6 VDD2.n2 VDD2.n0 115.142
R7 VDD2.n2 VDD2.n1 70.367
R8 VDD2.n1 VDD2.t0 1.97289
R9 VDD2.n1 VDD2.t2 1.97289
R10 VDD2.n0 VDD2.t1 1.97289
R11 VDD2.n0 VDD2.t3 1.97289
R12 VDD2 VDD2.n2 0.0586897
R13 VTAIL.n5 VTAIL.t1 55.6608
R14 VTAIL.n4 VTAIL.t4 55.6608
R15 VTAIL.n3 VTAIL.t6 55.6608
R16 VTAIL.n7 VTAIL.t3 55.6606
R17 VTAIL.n0 VTAIL.t5 55.6606
R18 VTAIL.n1 VTAIL.t0 55.6606
R19 VTAIL.n2 VTAIL.t7 55.6606
R20 VTAIL.n6 VTAIL.t2 55.6606
R21 VTAIL.n7 VTAIL.n6 28.8583
R22 VTAIL.n3 VTAIL.n2 28.8583
R23 VTAIL.n4 VTAIL.n3 2.28498
R24 VTAIL.n6 VTAIL.n5 2.28498
R25 VTAIL.n2 VTAIL.n1 2.28498
R26 VTAIL VTAIL.n0 1.20093
R27 VTAIL VTAIL.n7 1.08455
R28 VTAIL.n5 VTAIL.n4 0.470328
R29 VTAIL.n1 VTAIL.n0 0.470328
R30 VP.n3 VP.t2 207.739
R31 VP.n3 VP.t0 207.083
R32 VP.n5 VP.t1 171.194
R33 VP.n13 VP.t3 171.194
R34 VP.n12 VP.n0 161.3
R35 VP.n11 VP.n10 161.3
R36 VP.n9 VP.n1 161.3
R37 VP.n8 VP.n7 161.3
R38 VP.n6 VP.n2 161.3
R39 VP.n5 VP.n4 94.9235
R40 VP.n14 VP.n13 94.9235
R41 VP.n4 VP.n3 54.3524
R42 VP.n7 VP.n1 40.577
R43 VP.n11 VP.n1 40.577
R44 VP.n7 VP.n6 24.5923
R45 VP.n12 VP.n11 24.5923
R46 VP.n6 VP.n5 15.9852
R47 VP.n13 VP.n12 15.9852
R48 VP.n4 VP.n2 0.278335
R49 VP.n14 VP.n0 0.278335
R50 VP.n8 VP.n2 0.189894
R51 VP.n9 VP.n8 0.189894
R52 VP.n10 VP.n9 0.189894
R53 VP.n10 VP.n0 0.189894
R54 VP VP.n14 0.153485
R55 VDD1 VDD1.n1 115.666
R56 VDD1 VDD1.n0 70.4252
R57 VDD1.n0 VDD1.t1 1.97289
R58 VDD1.n0 VDD1.t3 1.97289
R59 VDD1.n1 VDD1.t2 1.97289
R60 VDD1.n1 VDD1.t0 1.97289
R61 B.n416 B.n113 585
R62 B.n415 B.n414 585
R63 B.n413 B.n114 585
R64 B.n412 B.n411 585
R65 B.n410 B.n115 585
R66 B.n409 B.n408 585
R67 B.n407 B.n116 585
R68 B.n406 B.n405 585
R69 B.n404 B.n117 585
R70 B.n403 B.n402 585
R71 B.n401 B.n118 585
R72 B.n400 B.n399 585
R73 B.n398 B.n119 585
R74 B.n397 B.n396 585
R75 B.n395 B.n120 585
R76 B.n394 B.n393 585
R77 B.n392 B.n121 585
R78 B.n391 B.n390 585
R79 B.n389 B.n122 585
R80 B.n388 B.n387 585
R81 B.n386 B.n123 585
R82 B.n385 B.n384 585
R83 B.n383 B.n124 585
R84 B.n382 B.n381 585
R85 B.n380 B.n125 585
R86 B.n379 B.n378 585
R87 B.n377 B.n126 585
R88 B.n376 B.n375 585
R89 B.n374 B.n127 585
R90 B.n373 B.n372 585
R91 B.n371 B.n128 585
R92 B.n370 B.n369 585
R93 B.n368 B.n129 585
R94 B.n367 B.n366 585
R95 B.n365 B.n130 585
R96 B.n364 B.n363 585
R97 B.n362 B.n131 585
R98 B.n361 B.n360 585
R99 B.n359 B.n132 585
R100 B.n358 B.n357 585
R101 B.n356 B.n133 585
R102 B.n355 B.n354 585
R103 B.n353 B.n134 585
R104 B.n352 B.n351 585
R105 B.n350 B.n135 585
R106 B.n349 B.n348 585
R107 B.n347 B.n136 585
R108 B.n346 B.n345 585
R109 B.n344 B.n137 585
R110 B.n343 B.n342 585
R111 B.n341 B.n138 585
R112 B.n340 B.n339 585
R113 B.n338 B.n139 585
R114 B.n337 B.n336 585
R115 B.n335 B.n140 585
R116 B.n334 B.n333 585
R117 B.n329 B.n141 585
R118 B.n328 B.n327 585
R119 B.n326 B.n142 585
R120 B.n325 B.n324 585
R121 B.n323 B.n143 585
R122 B.n322 B.n321 585
R123 B.n320 B.n144 585
R124 B.n319 B.n318 585
R125 B.n316 B.n145 585
R126 B.n315 B.n314 585
R127 B.n313 B.n148 585
R128 B.n312 B.n311 585
R129 B.n310 B.n149 585
R130 B.n309 B.n308 585
R131 B.n307 B.n150 585
R132 B.n306 B.n305 585
R133 B.n304 B.n151 585
R134 B.n303 B.n302 585
R135 B.n301 B.n152 585
R136 B.n300 B.n299 585
R137 B.n298 B.n153 585
R138 B.n297 B.n296 585
R139 B.n295 B.n154 585
R140 B.n294 B.n293 585
R141 B.n292 B.n155 585
R142 B.n291 B.n290 585
R143 B.n289 B.n156 585
R144 B.n288 B.n287 585
R145 B.n286 B.n157 585
R146 B.n285 B.n284 585
R147 B.n283 B.n158 585
R148 B.n282 B.n281 585
R149 B.n280 B.n159 585
R150 B.n279 B.n278 585
R151 B.n277 B.n160 585
R152 B.n276 B.n275 585
R153 B.n274 B.n161 585
R154 B.n273 B.n272 585
R155 B.n271 B.n162 585
R156 B.n270 B.n269 585
R157 B.n268 B.n163 585
R158 B.n267 B.n266 585
R159 B.n265 B.n164 585
R160 B.n264 B.n263 585
R161 B.n262 B.n165 585
R162 B.n261 B.n260 585
R163 B.n259 B.n166 585
R164 B.n258 B.n257 585
R165 B.n256 B.n167 585
R166 B.n255 B.n254 585
R167 B.n253 B.n168 585
R168 B.n252 B.n251 585
R169 B.n250 B.n169 585
R170 B.n249 B.n248 585
R171 B.n247 B.n170 585
R172 B.n246 B.n245 585
R173 B.n244 B.n171 585
R174 B.n243 B.n242 585
R175 B.n241 B.n172 585
R176 B.n240 B.n239 585
R177 B.n238 B.n173 585
R178 B.n237 B.n236 585
R179 B.n235 B.n174 585
R180 B.n418 B.n417 585
R181 B.n419 B.n112 585
R182 B.n421 B.n420 585
R183 B.n422 B.n111 585
R184 B.n424 B.n423 585
R185 B.n425 B.n110 585
R186 B.n427 B.n426 585
R187 B.n428 B.n109 585
R188 B.n430 B.n429 585
R189 B.n431 B.n108 585
R190 B.n433 B.n432 585
R191 B.n434 B.n107 585
R192 B.n436 B.n435 585
R193 B.n437 B.n106 585
R194 B.n439 B.n438 585
R195 B.n440 B.n105 585
R196 B.n442 B.n441 585
R197 B.n443 B.n104 585
R198 B.n445 B.n444 585
R199 B.n446 B.n103 585
R200 B.n448 B.n447 585
R201 B.n449 B.n102 585
R202 B.n451 B.n450 585
R203 B.n452 B.n101 585
R204 B.n454 B.n453 585
R205 B.n455 B.n100 585
R206 B.n457 B.n456 585
R207 B.n458 B.n99 585
R208 B.n460 B.n459 585
R209 B.n461 B.n98 585
R210 B.n463 B.n462 585
R211 B.n464 B.n97 585
R212 B.n466 B.n465 585
R213 B.n467 B.n96 585
R214 B.n469 B.n468 585
R215 B.n470 B.n95 585
R216 B.n472 B.n471 585
R217 B.n473 B.n94 585
R218 B.n475 B.n474 585
R219 B.n476 B.n93 585
R220 B.n478 B.n477 585
R221 B.n479 B.n92 585
R222 B.n481 B.n480 585
R223 B.n482 B.n91 585
R224 B.n484 B.n483 585
R225 B.n485 B.n90 585
R226 B.n487 B.n486 585
R227 B.n488 B.n89 585
R228 B.n490 B.n489 585
R229 B.n491 B.n88 585
R230 B.n493 B.n492 585
R231 B.n494 B.n87 585
R232 B.n496 B.n495 585
R233 B.n497 B.n86 585
R234 B.n499 B.n498 585
R235 B.n500 B.n85 585
R236 B.n502 B.n501 585
R237 B.n503 B.n84 585
R238 B.n505 B.n504 585
R239 B.n506 B.n83 585
R240 B.n508 B.n507 585
R241 B.n509 B.n82 585
R242 B.n511 B.n510 585
R243 B.n512 B.n81 585
R244 B.n693 B.n692 585
R245 B.n691 B.n18 585
R246 B.n690 B.n689 585
R247 B.n688 B.n19 585
R248 B.n687 B.n686 585
R249 B.n685 B.n20 585
R250 B.n684 B.n683 585
R251 B.n682 B.n21 585
R252 B.n681 B.n680 585
R253 B.n679 B.n22 585
R254 B.n678 B.n677 585
R255 B.n676 B.n23 585
R256 B.n675 B.n674 585
R257 B.n673 B.n24 585
R258 B.n672 B.n671 585
R259 B.n670 B.n25 585
R260 B.n669 B.n668 585
R261 B.n667 B.n26 585
R262 B.n666 B.n665 585
R263 B.n664 B.n27 585
R264 B.n663 B.n662 585
R265 B.n661 B.n28 585
R266 B.n660 B.n659 585
R267 B.n658 B.n29 585
R268 B.n657 B.n656 585
R269 B.n655 B.n30 585
R270 B.n654 B.n653 585
R271 B.n652 B.n31 585
R272 B.n651 B.n650 585
R273 B.n649 B.n32 585
R274 B.n648 B.n647 585
R275 B.n646 B.n33 585
R276 B.n645 B.n644 585
R277 B.n643 B.n34 585
R278 B.n642 B.n641 585
R279 B.n640 B.n35 585
R280 B.n639 B.n638 585
R281 B.n637 B.n36 585
R282 B.n636 B.n635 585
R283 B.n634 B.n37 585
R284 B.n633 B.n632 585
R285 B.n631 B.n38 585
R286 B.n630 B.n629 585
R287 B.n628 B.n39 585
R288 B.n627 B.n626 585
R289 B.n625 B.n40 585
R290 B.n624 B.n623 585
R291 B.n622 B.n41 585
R292 B.n621 B.n620 585
R293 B.n619 B.n42 585
R294 B.n618 B.n617 585
R295 B.n616 B.n43 585
R296 B.n615 B.n614 585
R297 B.n613 B.n44 585
R298 B.n612 B.n611 585
R299 B.n609 B.n45 585
R300 B.n608 B.n607 585
R301 B.n606 B.n48 585
R302 B.n605 B.n604 585
R303 B.n603 B.n49 585
R304 B.n602 B.n601 585
R305 B.n600 B.n50 585
R306 B.n599 B.n598 585
R307 B.n597 B.n51 585
R308 B.n595 B.n594 585
R309 B.n593 B.n54 585
R310 B.n592 B.n591 585
R311 B.n590 B.n55 585
R312 B.n589 B.n588 585
R313 B.n587 B.n56 585
R314 B.n586 B.n585 585
R315 B.n584 B.n57 585
R316 B.n583 B.n582 585
R317 B.n581 B.n58 585
R318 B.n580 B.n579 585
R319 B.n578 B.n59 585
R320 B.n577 B.n576 585
R321 B.n575 B.n60 585
R322 B.n574 B.n573 585
R323 B.n572 B.n61 585
R324 B.n571 B.n570 585
R325 B.n569 B.n62 585
R326 B.n568 B.n567 585
R327 B.n566 B.n63 585
R328 B.n565 B.n564 585
R329 B.n563 B.n64 585
R330 B.n562 B.n561 585
R331 B.n560 B.n65 585
R332 B.n559 B.n558 585
R333 B.n557 B.n66 585
R334 B.n556 B.n555 585
R335 B.n554 B.n67 585
R336 B.n553 B.n552 585
R337 B.n551 B.n68 585
R338 B.n550 B.n549 585
R339 B.n548 B.n69 585
R340 B.n547 B.n546 585
R341 B.n545 B.n70 585
R342 B.n544 B.n543 585
R343 B.n542 B.n71 585
R344 B.n541 B.n540 585
R345 B.n539 B.n72 585
R346 B.n538 B.n537 585
R347 B.n536 B.n73 585
R348 B.n535 B.n534 585
R349 B.n533 B.n74 585
R350 B.n532 B.n531 585
R351 B.n530 B.n75 585
R352 B.n529 B.n528 585
R353 B.n527 B.n76 585
R354 B.n526 B.n525 585
R355 B.n524 B.n77 585
R356 B.n523 B.n522 585
R357 B.n521 B.n78 585
R358 B.n520 B.n519 585
R359 B.n518 B.n79 585
R360 B.n517 B.n516 585
R361 B.n515 B.n80 585
R362 B.n514 B.n513 585
R363 B.n694 B.n17 585
R364 B.n696 B.n695 585
R365 B.n697 B.n16 585
R366 B.n699 B.n698 585
R367 B.n700 B.n15 585
R368 B.n702 B.n701 585
R369 B.n703 B.n14 585
R370 B.n705 B.n704 585
R371 B.n706 B.n13 585
R372 B.n708 B.n707 585
R373 B.n709 B.n12 585
R374 B.n711 B.n710 585
R375 B.n712 B.n11 585
R376 B.n714 B.n713 585
R377 B.n715 B.n10 585
R378 B.n717 B.n716 585
R379 B.n718 B.n9 585
R380 B.n720 B.n719 585
R381 B.n721 B.n8 585
R382 B.n723 B.n722 585
R383 B.n724 B.n7 585
R384 B.n726 B.n725 585
R385 B.n727 B.n6 585
R386 B.n729 B.n728 585
R387 B.n730 B.n5 585
R388 B.n732 B.n731 585
R389 B.n733 B.n4 585
R390 B.n735 B.n734 585
R391 B.n736 B.n3 585
R392 B.n738 B.n737 585
R393 B.n739 B.n0 585
R394 B.n2 B.n1 585
R395 B.n190 B.n189 585
R396 B.n192 B.n191 585
R397 B.n193 B.n188 585
R398 B.n195 B.n194 585
R399 B.n196 B.n187 585
R400 B.n198 B.n197 585
R401 B.n199 B.n186 585
R402 B.n201 B.n200 585
R403 B.n202 B.n185 585
R404 B.n204 B.n203 585
R405 B.n205 B.n184 585
R406 B.n207 B.n206 585
R407 B.n208 B.n183 585
R408 B.n210 B.n209 585
R409 B.n211 B.n182 585
R410 B.n213 B.n212 585
R411 B.n214 B.n181 585
R412 B.n216 B.n215 585
R413 B.n217 B.n180 585
R414 B.n219 B.n218 585
R415 B.n220 B.n179 585
R416 B.n222 B.n221 585
R417 B.n223 B.n178 585
R418 B.n225 B.n224 585
R419 B.n226 B.n177 585
R420 B.n228 B.n227 585
R421 B.n229 B.n176 585
R422 B.n231 B.n230 585
R423 B.n232 B.n175 585
R424 B.n234 B.n233 585
R425 B.n235 B.n234 511.721
R426 B.n418 B.n113 511.721
R427 B.n514 B.n81 511.721
R428 B.n692 B.n17 511.721
R429 B.n146 B.t6 378.774
R430 B.n330 B.t3 378.774
R431 B.n52 B.t9 378.774
R432 B.n46 B.t0 378.774
R433 B.n741 B.n740 256.663
R434 B.n740 B.n739 235.042
R435 B.n740 B.n2 235.042
R436 B.n236 B.n235 163.367
R437 B.n236 B.n173 163.367
R438 B.n240 B.n173 163.367
R439 B.n241 B.n240 163.367
R440 B.n242 B.n241 163.367
R441 B.n242 B.n171 163.367
R442 B.n246 B.n171 163.367
R443 B.n247 B.n246 163.367
R444 B.n248 B.n247 163.367
R445 B.n248 B.n169 163.367
R446 B.n252 B.n169 163.367
R447 B.n253 B.n252 163.367
R448 B.n254 B.n253 163.367
R449 B.n254 B.n167 163.367
R450 B.n258 B.n167 163.367
R451 B.n259 B.n258 163.367
R452 B.n260 B.n259 163.367
R453 B.n260 B.n165 163.367
R454 B.n264 B.n165 163.367
R455 B.n265 B.n264 163.367
R456 B.n266 B.n265 163.367
R457 B.n266 B.n163 163.367
R458 B.n270 B.n163 163.367
R459 B.n271 B.n270 163.367
R460 B.n272 B.n271 163.367
R461 B.n272 B.n161 163.367
R462 B.n276 B.n161 163.367
R463 B.n277 B.n276 163.367
R464 B.n278 B.n277 163.367
R465 B.n278 B.n159 163.367
R466 B.n282 B.n159 163.367
R467 B.n283 B.n282 163.367
R468 B.n284 B.n283 163.367
R469 B.n284 B.n157 163.367
R470 B.n288 B.n157 163.367
R471 B.n289 B.n288 163.367
R472 B.n290 B.n289 163.367
R473 B.n290 B.n155 163.367
R474 B.n294 B.n155 163.367
R475 B.n295 B.n294 163.367
R476 B.n296 B.n295 163.367
R477 B.n296 B.n153 163.367
R478 B.n300 B.n153 163.367
R479 B.n301 B.n300 163.367
R480 B.n302 B.n301 163.367
R481 B.n302 B.n151 163.367
R482 B.n306 B.n151 163.367
R483 B.n307 B.n306 163.367
R484 B.n308 B.n307 163.367
R485 B.n308 B.n149 163.367
R486 B.n312 B.n149 163.367
R487 B.n313 B.n312 163.367
R488 B.n314 B.n313 163.367
R489 B.n314 B.n145 163.367
R490 B.n319 B.n145 163.367
R491 B.n320 B.n319 163.367
R492 B.n321 B.n320 163.367
R493 B.n321 B.n143 163.367
R494 B.n325 B.n143 163.367
R495 B.n326 B.n325 163.367
R496 B.n327 B.n326 163.367
R497 B.n327 B.n141 163.367
R498 B.n334 B.n141 163.367
R499 B.n335 B.n334 163.367
R500 B.n336 B.n335 163.367
R501 B.n336 B.n139 163.367
R502 B.n340 B.n139 163.367
R503 B.n341 B.n340 163.367
R504 B.n342 B.n341 163.367
R505 B.n342 B.n137 163.367
R506 B.n346 B.n137 163.367
R507 B.n347 B.n346 163.367
R508 B.n348 B.n347 163.367
R509 B.n348 B.n135 163.367
R510 B.n352 B.n135 163.367
R511 B.n353 B.n352 163.367
R512 B.n354 B.n353 163.367
R513 B.n354 B.n133 163.367
R514 B.n358 B.n133 163.367
R515 B.n359 B.n358 163.367
R516 B.n360 B.n359 163.367
R517 B.n360 B.n131 163.367
R518 B.n364 B.n131 163.367
R519 B.n365 B.n364 163.367
R520 B.n366 B.n365 163.367
R521 B.n366 B.n129 163.367
R522 B.n370 B.n129 163.367
R523 B.n371 B.n370 163.367
R524 B.n372 B.n371 163.367
R525 B.n372 B.n127 163.367
R526 B.n376 B.n127 163.367
R527 B.n377 B.n376 163.367
R528 B.n378 B.n377 163.367
R529 B.n378 B.n125 163.367
R530 B.n382 B.n125 163.367
R531 B.n383 B.n382 163.367
R532 B.n384 B.n383 163.367
R533 B.n384 B.n123 163.367
R534 B.n388 B.n123 163.367
R535 B.n389 B.n388 163.367
R536 B.n390 B.n389 163.367
R537 B.n390 B.n121 163.367
R538 B.n394 B.n121 163.367
R539 B.n395 B.n394 163.367
R540 B.n396 B.n395 163.367
R541 B.n396 B.n119 163.367
R542 B.n400 B.n119 163.367
R543 B.n401 B.n400 163.367
R544 B.n402 B.n401 163.367
R545 B.n402 B.n117 163.367
R546 B.n406 B.n117 163.367
R547 B.n407 B.n406 163.367
R548 B.n408 B.n407 163.367
R549 B.n408 B.n115 163.367
R550 B.n412 B.n115 163.367
R551 B.n413 B.n412 163.367
R552 B.n414 B.n413 163.367
R553 B.n414 B.n113 163.367
R554 B.n510 B.n81 163.367
R555 B.n510 B.n509 163.367
R556 B.n509 B.n508 163.367
R557 B.n508 B.n83 163.367
R558 B.n504 B.n83 163.367
R559 B.n504 B.n503 163.367
R560 B.n503 B.n502 163.367
R561 B.n502 B.n85 163.367
R562 B.n498 B.n85 163.367
R563 B.n498 B.n497 163.367
R564 B.n497 B.n496 163.367
R565 B.n496 B.n87 163.367
R566 B.n492 B.n87 163.367
R567 B.n492 B.n491 163.367
R568 B.n491 B.n490 163.367
R569 B.n490 B.n89 163.367
R570 B.n486 B.n89 163.367
R571 B.n486 B.n485 163.367
R572 B.n485 B.n484 163.367
R573 B.n484 B.n91 163.367
R574 B.n480 B.n91 163.367
R575 B.n480 B.n479 163.367
R576 B.n479 B.n478 163.367
R577 B.n478 B.n93 163.367
R578 B.n474 B.n93 163.367
R579 B.n474 B.n473 163.367
R580 B.n473 B.n472 163.367
R581 B.n472 B.n95 163.367
R582 B.n468 B.n95 163.367
R583 B.n468 B.n467 163.367
R584 B.n467 B.n466 163.367
R585 B.n466 B.n97 163.367
R586 B.n462 B.n97 163.367
R587 B.n462 B.n461 163.367
R588 B.n461 B.n460 163.367
R589 B.n460 B.n99 163.367
R590 B.n456 B.n99 163.367
R591 B.n456 B.n455 163.367
R592 B.n455 B.n454 163.367
R593 B.n454 B.n101 163.367
R594 B.n450 B.n101 163.367
R595 B.n450 B.n449 163.367
R596 B.n449 B.n448 163.367
R597 B.n448 B.n103 163.367
R598 B.n444 B.n103 163.367
R599 B.n444 B.n443 163.367
R600 B.n443 B.n442 163.367
R601 B.n442 B.n105 163.367
R602 B.n438 B.n105 163.367
R603 B.n438 B.n437 163.367
R604 B.n437 B.n436 163.367
R605 B.n436 B.n107 163.367
R606 B.n432 B.n107 163.367
R607 B.n432 B.n431 163.367
R608 B.n431 B.n430 163.367
R609 B.n430 B.n109 163.367
R610 B.n426 B.n109 163.367
R611 B.n426 B.n425 163.367
R612 B.n425 B.n424 163.367
R613 B.n424 B.n111 163.367
R614 B.n420 B.n111 163.367
R615 B.n420 B.n419 163.367
R616 B.n419 B.n418 163.367
R617 B.n692 B.n691 163.367
R618 B.n691 B.n690 163.367
R619 B.n690 B.n19 163.367
R620 B.n686 B.n19 163.367
R621 B.n686 B.n685 163.367
R622 B.n685 B.n684 163.367
R623 B.n684 B.n21 163.367
R624 B.n680 B.n21 163.367
R625 B.n680 B.n679 163.367
R626 B.n679 B.n678 163.367
R627 B.n678 B.n23 163.367
R628 B.n674 B.n23 163.367
R629 B.n674 B.n673 163.367
R630 B.n673 B.n672 163.367
R631 B.n672 B.n25 163.367
R632 B.n668 B.n25 163.367
R633 B.n668 B.n667 163.367
R634 B.n667 B.n666 163.367
R635 B.n666 B.n27 163.367
R636 B.n662 B.n27 163.367
R637 B.n662 B.n661 163.367
R638 B.n661 B.n660 163.367
R639 B.n660 B.n29 163.367
R640 B.n656 B.n29 163.367
R641 B.n656 B.n655 163.367
R642 B.n655 B.n654 163.367
R643 B.n654 B.n31 163.367
R644 B.n650 B.n31 163.367
R645 B.n650 B.n649 163.367
R646 B.n649 B.n648 163.367
R647 B.n648 B.n33 163.367
R648 B.n644 B.n33 163.367
R649 B.n644 B.n643 163.367
R650 B.n643 B.n642 163.367
R651 B.n642 B.n35 163.367
R652 B.n638 B.n35 163.367
R653 B.n638 B.n637 163.367
R654 B.n637 B.n636 163.367
R655 B.n636 B.n37 163.367
R656 B.n632 B.n37 163.367
R657 B.n632 B.n631 163.367
R658 B.n631 B.n630 163.367
R659 B.n630 B.n39 163.367
R660 B.n626 B.n39 163.367
R661 B.n626 B.n625 163.367
R662 B.n625 B.n624 163.367
R663 B.n624 B.n41 163.367
R664 B.n620 B.n41 163.367
R665 B.n620 B.n619 163.367
R666 B.n619 B.n618 163.367
R667 B.n618 B.n43 163.367
R668 B.n614 B.n43 163.367
R669 B.n614 B.n613 163.367
R670 B.n613 B.n612 163.367
R671 B.n612 B.n45 163.367
R672 B.n607 B.n45 163.367
R673 B.n607 B.n606 163.367
R674 B.n606 B.n605 163.367
R675 B.n605 B.n49 163.367
R676 B.n601 B.n49 163.367
R677 B.n601 B.n600 163.367
R678 B.n600 B.n599 163.367
R679 B.n599 B.n51 163.367
R680 B.n594 B.n51 163.367
R681 B.n594 B.n593 163.367
R682 B.n593 B.n592 163.367
R683 B.n592 B.n55 163.367
R684 B.n588 B.n55 163.367
R685 B.n588 B.n587 163.367
R686 B.n587 B.n586 163.367
R687 B.n586 B.n57 163.367
R688 B.n582 B.n57 163.367
R689 B.n582 B.n581 163.367
R690 B.n581 B.n580 163.367
R691 B.n580 B.n59 163.367
R692 B.n576 B.n59 163.367
R693 B.n576 B.n575 163.367
R694 B.n575 B.n574 163.367
R695 B.n574 B.n61 163.367
R696 B.n570 B.n61 163.367
R697 B.n570 B.n569 163.367
R698 B.n569 B.n568 163.367
R699 B.n568 B.n63 163.367
R700 B.n564 B.n63 163.367
R701 B.n564 B.n563 163.367
R702 B.n563 B.n562 163.367
R703 B.n562 B.n65 163.367
R704 B.n558 B.n65 163.367
R705 B.n558 B.n557 163.367
R706 B.n557 B.n556 163.367
R707 B.n556 B.n67 163.367
R708 B.n552 B.n67 163.367
R709 B.n552 B.n551 163.367
R710 B.n551 B.n550 163.367
R711 B.n550 B.n69 163.367
R712 B.n546 B.n69 163.367
R713 B.n546 B.n545 163.367
R714 B.n545 B.n544 163.367
R715 B.n544 B.n71 163.367
R716 B.n540 B.n71 163.367
R717 B.n540 B.n539 163.367
R718 B.n539 B.n538 163.367
R719 B.n538 B.n73 163.367
R720 B.n534 B.n73 163.367
R721 B.n534 B.n533 163.367
R722 B.n533 B.n532 163.367
R723 B.n532 B.n75 163.367
R724 B.n528 B.n75 163.367
R725 B.n528 B.n527 163.367
R726 B.n527 B.n526 163.367
R727 B.n526 B.n77 163.367
R728 B.n522 B.n77 163.367
R729 B.n522 B.n521 163.367
R730 B.n521 B.n520 163.367
R731 B.n520 B.n79 163.367
R732 B.n516 B.n79 163.367
R733 B.n516 B.n515 163.367
R734 B.n515 B.n514 163.367
R735 B.n696 B.n17 163.367
R736 B.n697 B.n696 163.367
R737 B.n698 B.n697 163.367
R738 B.n698 B.n15 163.367
R739 B.n702 B.n15 163.367
R740 B.n703 B.n702 163.367
R741 B.n704 B.n703 163.367
R742 B.n704 B.n13 163.367
R743 B.n708 B.n13 163.367
R744 B.n709 B.n708 163.367
R745 B.n710 B.n709 163.367
R746 B.n710 B.n11 163.367
R747 B.n714 B.n11 163.367
R748 B.n715 B.n714 163.367
R749 B.n716 B.n715 163.367
R750 B.n716 B.n9 163.367
R751 B.n720 B.n9 163.367
R752 B.n721 B.n720 163.367
R753 B.n722 B.n721 163.367
R754 B.n722 B.n7 163.367
R755 B.n726 B.n7 163.367
R756 B.n727 B.n726 163.367
R757 B.n728 B.n727 163.367
R758 B.n728 B.n5 163.367
R759 B.n732 B.n5 163.367
R760 B.n733 B.n732 163.367
R761 B.n734 B.n733 163.367
R762 B.n734 B.n3 163.367
R763 B.n738 B.n3 163.367
R764 B.n739 B.n738 163.367
R765 B.n189 B.n2 163.367
R766 B.n192 B.n189 163.367
R767 B.n193 B.n192 163.367
R768 B.n194 B.n193 163.367
R769 B.n194 B.n187 163.367
R770 B.n198 B.n187 163.367
R771 B.n199 B.n198 163.367
R772 B.n200 B.n199 163.367
R773 B.n200 B.n185 163.367
R774 B.n204 B.n185 163.367
R775 B.n205 B.n204 163.367
R776 B.n206 B.n205 163.367
R777 B.n206 B.n183 163.367
R778 B.n210 B.n183 163.367
R779 B.n211 B.n210 163.367
R780 B.n212 B.n211 163.367
R781 B.n212 B.n181 163.367
R782 B.n216 B.n181 163.367
R783 B.n217 B.n216 163.367
R784 B.n218 B.n217 163.367
R785 B.n218 B.n179 163.367
R786 B.n222 B.n179 163.367
R787 B.n223 B.n222 163.367
R788 B.n224 B.n223 163.367
R789 B.n224 B.n177 163.367
R790 B.n228 B.n177 163.367
R791 B.n229 B.n228 163.367
R792 B.n230 B.n229 163.367
R793 B.n230 B.n175 163.367
R794 B.n234 B.n175 163.367
R795 B.n330 B.t4 160.865
R796 B.n52 B.t11 160.865
R797 B.n146 B.t7 160.845
R798 B.n46 B.t2 160.845
R799 B.n331 B.t5 109.472
R800 B.n53 B.t10 109.472
R801 B.n147 B.t8 109.451
R802 B.n47 B.t1 109.451
R803 B.n317 B.n147 59.5399
R804 B.n332 B.n331 59.5399
R805 B.n596 B.n53 59.5399
R806 B.n610 B.n47 59.5399
R807 B.n147 B.n146 51.3944
R808 B.n331 B.n330 51.3944
R809 B.n53 B.n52 51.3944
R810 B.n47 B.n46 51.3944
R811 B.n694 B.n693 33.2493
R812 B.n513 B.n512 33.2493
R813 B.n417 B.n416 33.2493
R814 B.n233 B.n174 33.2493
R815 B B.n741 18.0485
R816 B.n695 B.n694 10.6151
R817 B.n695 B.n16 10.6151
R818 B.n699 B.n16 10.6151
R819 B.n700 B.n699 10.6151
R820 B.n701 B.n700 10.6151
R821 B.n701 B.n14 10.6151
R822 B.n705 B.n14 10.6151
R823 B.n706 B.n705 10.6151
R824 B.n707 B.n706 10.6151
R825 B.n707 B.n12 10.6151
R826 B.n711 B.n12 10.6151
R827 B.n712 B.n711 10.6151
R828 B.n713 B.n712 10.6151
R829 B.n713 B.n10 10.6151
R830 B.n717 B.n10 10.6151
R831 B.n718 B.n717 10.6151
R832 B.n719 B.n718 10.6151
R833 B.n719 B.n8 10.6151
R834 B.n723 B.n8 10.6151
R835 B.n724 B.n723 10.6151
R836 B.n725 B.n724 10.6151
R837 B.n725 B.n6 10.6151
R838 B.n729 B.n6 10.6151
R839 B.n730 B.n729 10.6151
R840 B.n731 B.n730 10.6151
R841 B.n731 B.n4 10.6151
R842 B.n735 B.n4 10.6151
R843 B.n736 B.n735 10.6151
R844 B.n737 B.n736 10.6151
R845 B.n737 B.n0 10.6151
R846 B.n693 B.n18 10.6151
R847 B.n689 B.n18 10.6151
R848 B.n689 B.n688 10.6151
R849 B.n688 B.n687 10.6151
R850 B.n687 B.n20 10.6151
R851 B.n683 B.n20 10.6151
R852 B.n683 B.n682 10.6151
R853 B.n682 B.n681 10.6151
R854 B.n681 B.n22 10.6151
R855 B.n677 B.n22 10.6151
R856 B.n677 B.n676 10.6151
R857 B.n676 B.n675 10.6151
R858 B.n675 B.n24 10.6151
R859 B.n671 B.n24 10.6151
R860 B.n671 B.n670 10.6151
R861 B.n670 B.n669 10.6151
R862 B.n669 B.n26 10.6151
R863 B.n665 B.n26 10.6151
R864 B.n665 B.n664 10.6151
R865 B.n664 B.n663 10.6151
R866 B.n663 B.n28 10.6151
R867 B.n659 B.n28 10.6151
R868 B.n659 B.n658 10.6151
R869 B.n658 B.n657 10.6151
R870 B.n657 B.n30 10.6151
R871 B.n653 B.n30 10.6151
R872 B.n653 B.n652 10.6151
R873 B.n652 B.n651 10.6151
R874 B.n651 B.n32 10.6151
R875 B.n647 B.n32 10.6151
R876 B.n647 B.n646 10.6151
R877 B.n646 B.n645 10.6151
R878 B.n645 B.n34 10.6151
R879 B.n641 B.n34 10.6151
R880 B.n641 B.n640 10.6151
R881 B.n640 B.n639 10.6151
R882 B.n639 B.n36 10.6151
R883 B.n635 B.n36 10.6151
R884 B.n635 B.n634 10.6151
R885 B.n634 B.n633 10.6151
R886 B.n633 B.n38 10.6151
R887 B.n629 B.n38 10.6151
R888 B.n629 B.n628 10.6151
R889 B.n628 B.n627 10.6151
R890 B.n627 B.n40 10.6151
R891 B.n623 B.n40 10.6151
R892 B.n623 B.n622 10.6151
R893 B.n622 B.n621 10.6151
R894 B.n621 B.n42 10.6151
R895 B.n617 B.n42 10.6151
R896 B.n617 B.n616 10.6151
R897 B.n616 B.n615 10.6151
R898 B.n615 B.n44 10.6151
R899 B.n611 B.n44 10.6151
R900 B.n609 B.n608 10.6151
R901 B.n608 B.n48 10.6151
R902 B.n604 B.n48 10.6151
R903 B.n604 B.n603 10.6151
R904 B.n603 B.n602 10.6151
R905 B.n602 B.n50 10.6151
R906 B.n598 B.n50 10.6151
R907 B.n598 B.n597 10.6151
R908 B.n595 B.n54 10.6151
R909 B.n591 B.n54 10.6151
R910 B.n591 B.n590 10.6151
R911 B.n590 B.n589 10.6151
R912 B.n589 B.n56 10.6151
R913 B.n585 B.n56 10.6151
R914 B.n585 B.n584 10.6151
R915 B.n584 B.n583 10.6151
R916 B.n583 B.n58 10.6151
R917 B.n579 B.n58 10.6151
R918 B.n579 B.n578 10.6151
R919 B.n578 B.n577 10.6151
R920 B.n577 B.n60 10.6151
R921 B.n573 B.n60 10.6151
R922 B.n573 B.n572 10.6151
R923 B.n572 B.n571 10.6151
R924 B.n571 B.n62 10.6151
R925 B.n567 B.n62 10.6151
R926 B.n567 B.n566 10.6151
R927 B.n566 B.n565 10.6151
R928 B.n565 B.n64 10.6151
R929 B.n561 B.n64 10.6151
R930 B.n561 B.n560 10.6151
R931 B.n560 B.n559 10.6151
R932 B.n559 B.n66 10.6151
R933 B.n555 B.n66 10.6151
R934 B.n555 B.n554 10.6151
R935 B.n554 B.n553 10.6151
R936 B.n553 B.n68 10.6151
R937 B.n549 B.n68 10.6151
R938 B.n549 B.n548 10.6151
R939 B.n548 B.n547 10.6151
R940 B.n547 B.n70 10.6151
R941 B.n543 B.n70 10.6151
R942 B.n543 B.n542 10.6151
R943 B.n542 B.n541 10.6151
R944 B.n541 B.n72 10.6151
R945 B.n537 B.n72 10.6151
R946 B.n537 B.n536 10.6151
R947 B.n536 B.n535 10.6151
R948 B.n535 B.n74 10.6151
R949 B.n531 B.n74 10.6151
R950 B.n531 B.n530 10.6151
R951 B.n530 B.n529 10.6151
R952 B.n529 B.n76 10.6151
R953 B.n525 B.n76 10.6151
R954 B.n525 B.n524 10.6151
R955 B.n524 B.n523 10.6151
R956 B.n523 B.n78 10.6151
R957 B.n519 B.n78 10.6151
R958 B.n519 B.n518 10.6151
R959 B.n518 B.n517 10.6151
R960 B.n517 B.n80 10.6151
R961 B.n513 B.n80 10.6151
R962 B.n512 B.n511 10.6151
R963 B.n511 B.n82 10.6151
R964 B.n507 B.n82 10.6151
R965 B.n507 B.n506 10.6151
R966 B.n506 B.n505 10.6151
R967 B.n505 B.n84 10.6151
R968 B.n501 B.n84 10.6151
R969 B.n501 B.n500 10.6151
R970 B.n500 B.n499 10.6151
R971 B.n499 B.n86 10.6151
R972 B.n495 B.n86 10.6151
R973 B.n495 B.n494 10.6151
R974 B.n494 B.n493 10.6151
R975 B.n493 B.n88 10.6151
R976 B.n489 B.n88 10.6151
R977 B.n489 B.n488 10.6151
R978 B.n488 B.n487 10.6151
R979 B.n487 B.n90 10.6151
R980 B.n483 B.n90 10.6151
R981 B.n483 B.n482 10.6151
R982 B.n482 B.n481 10.6151
R983 B.n481 B.n92 10.6151
R984 B.n477 B.n92 10.6151
R985 B.n477 B.n476 10.6151
R986 B.n476 B.n475 10.6151
R987 B.n475 B.n94 10.6151
R988 B.n471 B.n94 10.6151
R989 B.n471 B.n470 10.6151
R990 B.n470 B.n469 10.6151
R991 B.n469 B.n96 10.6151
R992 B.n465 B.n96 10.6151
R993 B.n465 B.n464 10.6151
R994 B.n464 B.n463 10.6151
R995 B.n463 B.n98 10.6151
R996 B.n459 B.n98 10.6151
R997 B.n459 B.n458 10.6151
R998 B.n458 B.n457 10.6151
R999 B.n457 B.n100 10.6151
R1000 B.n453 B.n100 10.6151
R1001 B.n453 B.n452 10.6151
R1002 B.n452 B.n451 10.6151
R1003 B.n451 B.n102 10.6151
R1004 B.n447 B.n102 10.6151
R1005 B.n447 B.n446 10.6151
R1006 B.n446 B.n445 10.6151
R1007 B.n445 B.n104 10.6151
R1008 B.n441 B.n104 10.6151
R1009 B.n441 B.n440 10.6151
R1010 B.n440 B.n439 10.6151
R1011 B.n439 B.n106 10.6151
R1012 B.n435 B.n106 10.6151
R1013 B.n435 B.n434 10.6151
R1014 B.n434 B.n433 10.6151
R1015 B.n433 B.n108 10.6151
R1016 B.n429 B.n108 10.6151
R1017 B.n429 B.n428 10.6151
R1018 B.n428 B.n427 10.6151
R1019 B.n427 B.n110 10.6151
R1020 B.n423 B.n110 10.6151
R1021 B.n423 B.n422 10.6151
R1022 B.n422 B.n421 10.6151
R1023 B.n421 B.n112 10.6151
R1024 B.n417 B.n112 10.6151
R1025 B.n190 B.n1 10.6151
R1026 B.n191 B.n190 10.6151
R1027 B.n191 B.n188 10.6151
R1028 B.n195 B.n188 10.6151
R1029 B.n196 B.n195 10.6151
R1030 B.n197 B.n196 10.6151
R1031 B.n197 B.n186 10.6151
R1032 B.n201 B.n186 10.6151
R1033 B.n202 B.n201 10.6151
R1034 B.n203 B.n202 10.6151
R1035 B.n203 B.n184 10.6151
R1036 B.n207 B.n184 10.6151
R1037 B.n208 B.n207 10.6151
R1038 B.n209 B.n208 10.6151
R1039 B.n209 B.n182 10.6151
R1040 B.n213 B.n182 10.6151
R1041 B.n214 B.n213 10.6151
R1042 B.n215 B.n214 10.6151
R1043 B.n215 B.n180 10.6151
R1044 B.n219 B.n180 10.6151
R1045 B.n220 B.n219 10.6151
R1046 B.n221 B.n220 10.6151
R1047 B.n221 B.n178 10.6151
R1048 B.n225 B.n178 10.6151
R1049 B.n226 B.n225 10.6151
R1050 B.n227 B.n226 10.6151
R1051 B.n227 B.n176 10.6151
R1052 B.n231 B.n176 10.6151
R1053 B.n232 B.n231 10.6151
R1054 B.n233 B.n232 10.6151
R1055 B.n237 B.n174 10.6151
R1056 B.n238 B.n237 10.6151
R1057 B.n239 B.n238 10.6151
R1058 B.n239 B.n172 10.6151
R1059 B.n243 B.n172 10.6151
R1060 B.n244 B.n243 10.6151
R1061 B.n245 B.n244 10.6151
R1062 B.n245 B.n170 10.6151
R1063 B.n249 B.n170 10.6151
R1064 B.n250 B.n249 10.6151
R1065 B.n251 B.n250 10.6151
R1066 B.n251 B.n168 10.6151
R1067 B.n255 B.n168 10.6151
R1068 B.n256 B.n255 10.6151
R1069 B.n257 B.n256 10.6151
R1070 B.n257 B.n166 10.6151
R1071 B.n261 B.n166 10.6151
R1072 B.n262 B.n261 10.6151
R1073 B.n263 B.n262 10.6151
R1074 B.n263 B.n164 10.6151
R1075 B.n267 B.n164 10.6151
R1076 B.n268 B.n267 10.6151
R1077 B.n269 B.n268 10.6151
R1078 B.n269 B.n162 10.6151
R1079 B.n273 B.n162 10.6151
R1080 B.n274 B.n273 10.6151
R1081 B.n275 B.n274 10.6151
R1082 B.n275 B.n160 10.6151
R1083 B.n279 B.n160 10.6151
R1084 B.n280 B.n279 10.6151
R1085 B.n281 B.n280 10.6151
R1086 B.n281 B.n158 10.6151
R1087 B.n285 B.n158 10.6151
R1088 B.n286 B.n285 10.6151
R1089 B.n287 B.n286 10.6151
R1090 B.n287 B.n156 10.6151
R1091 B.n291 B.n156 10.6151
R1092 B.n292 B.n291 10.6151
R1093 B.n293 B.n292 10.6151
R1094 B.n293 B.n154 10.6151
R1095 B.n297 B.n154 10.6151
R1096 B.n298 B.n297 10.6151
R1097 B.n299 B.n298 10.6151
R1098 B.n299 B.n152 10.6151
R1099 B.n303 B.n152 10.6151
R1100 B.n304 B.n303 10.6151
R1101 B.n305 B.n304 10.6151
R1102 B.n305 B.n150 10.6151
R1103 B.n309 B.n150 10.6151
R1104 B.n310 B.n309 10.6151
R1105 B.n311 B.n310 10.6151
R1106 B.n311 B.n148 10.6151
R1107 B.n315 B.n148 10.6151
R1108 B.n316 B.n315 10.6151
R1109 B.n318 B.n144 10.6151
R1110 B.n322 B.n144 10.6151
R1111 B.n323 B.n322 10.6151
R1112 B.n324 B.n323 10.6151
R1113 B.n324 B.n142 10.6151
R1114 B.n328 B.n142 10.6151
R1115 B.n329 B.n328 10.6151
R1116 B.n333 B.n329 10.6151
R1117 B.n337 B.n140 10.6151
R1118 B.n338 B.n337 10.6151
R1119 B.n339 B.n338 10.6151
R1120 B.n339 B.n138 10.6151
R1121 B.n343 B.n138 10.6151
R1122 B.n344 B.n343 10.6151
R1123 B.n345 B.n344 10.6151
R1124 B.n345 B.n136 10.6151
R1125 B.n349 B.n136 10.6151
R1126 B.n350 B.n349 10.6151
R1127 B.n351 B.n350 10.6151
R1128 B.n351 B.n134 10.6151
R1129 B.n355 B.n134 10.6151
R1130 B.n356 B.n355 10.6151
R1131 B.n357 B.n356 10.6151
R1132 B.n357 B.n132 10.6151
R1133 B.n361 B.n132 10.6151
R1134 B.n362 B.n361 10.6151
R1135 B.n363 B.n362 10.6151
R1136 B.n363 B.n130 10.6151
R1137 B.n367 B.n130 10.6151
R1138 B.n368 B.n367 10.6151
R1139 B.n369 B.n368 10.6151
R1140 B.n369 B.n128 10.6151
R1141 B.n373 B.n128 10.6151
R1142 B.n374 B.n373 10.6151
R1143 B.n375 B.n374 10.6151
R1144 B.n375 B.n126 10.6151
R1145 B.n379 B.n126 10.6151
R1146 B.n380 B.n379 10.6151
R1147 B.n381 B.n380 10.6151
R1148 B.n381 B.n124 10.6151
R1149 B.n385 B.n124 10.6151
R1150 B.n386 B.n385 10.6151
R1151 B.n387 B.n386 10.6151
R1152 B.n387 B.n122 10.6151
R1153 B.n391 B.n122 10.6151
R1154 B.n392 B.n391 10.6151
R1155 B.n393 B.n392 10.6151
R1156 B.n393 B.n120 10.6151
R1157 B.n397 B.n120 10.6151
R1158 B.n398 B.n397 10.6151
R1159 B.n399 B.n398 10.6151
R1160 B.n399 B.n118 10.6151
R1161 B.n403 B.n118 10.6151
R1162 B.n404 B.n403 10.6151
R1163 B.n405 B.n404 10.6151
R1164 B.n405 B.n116 10.6151
R1165 B.n409 B.n116 10.6151
R1166 B.n410 B.n409 10.6151
R1167 B.n411 B.n410 10.6151
R1168 B.n411 B.n114 10.6151
R1169 B.n415 B.n114 10.6151
R1170 B.n416 B.n415 10.6151
R1171 B.n741 B.n0 8.11757
R1172 B.n741 B.n1 8.11757
R1173 B.n610 B.n609 6.5566
R1174 B.n597 B.n596 6.5566
R1175 B.n318 B.n317 6.5566
R1176 B.n333 B.n332 6.5566
R1177 B.n611 B.n610 4.05904
R1178 B.n596 B.n595 4.05904
R1179 B.n317 B.n316 4.05904
R1180 B.n332 B.n140 4.05904
C0 w_n2560_n4264# VTAIL 4.98864f
C1 VDD2 VN 6.27307f
C2 w_n2560_n4264# VP 4.69123f
C3 VDD1 VN 0.148911f
C4 VDD2 VTAIL 6.54292f
C5 VN B 1.11171f
C6 VDD1 VTAIL 6.49059f
C7 VDD2 VP 0.376653f
C8 VDD1 VP 6.50014f
C9 B VTAIL 6.261f
C10 w_n2560_n4264# VDD2 1.5664f
C11 B VP 1.65535f
C12 VDD1 w_n2560_n4264# 1.51654f
C13 w_n2560_n4264# B 10.158f
C14 VDD1 VDD2 0.962074f
C15 VN VTAIL 5.94535f
C16 VN VP 6.81418f
C17 VDD2 B 1.38198f
C18 VDD1 B 1.33444f
C19 w_n2560_n4264# VN 4.36284f
C20 VTAIL VP 5.95945f
C21 VDD2 VSUBS 0.999097f
C22 VDD1 VSUBS 6.14233f
C23 VTAIL VSUBS 1.395836f
C24 VN VSUBS 5.508759f
C25 VP VSUBS 2.30473f
C26 B VSUBS 4.407817f
C27 w_n2560_n4264# VSUBS 0.133663p
C28 B.n0 VSUBS 0.005637f
C29 B.n1 VSUBS 0.005637f
C30 B.n2 VSUBS 0.008337f
C31 B.n3 VSUBS 0.006388f
C32 B.n4 VSUBS 0.006388f
C33 B.n5 VSUBS 0.006388f
C34 B.n6 VSUBS 0.006388f
C35 B.n7 VSUBS 0.006388f
C36 B.n8 VSUBS 0.006388f
C37 B.n9 VSUBS 0.006388f
C38 B.n10 VSUBS 0.006388f
C39 B.n11 VSUBS 0.006388f
C40 B.n12 VSUBS 0.006388f
C41 B.n13 VSUBS 0.006388f
C42 B.n14 VSUBS 0.006388f
C43 B.n15 VSUBS 0.006388f
C44 B.n16 VSUBS 0.006388f
C45 B.n17 VSUBS 0.014827f
C46 B.n18 VSUBS 0.006388f
C47 B.n19 VSUBS 0.006388f
C48 B.n20 VSUBS 0.006388f
C49 B.n21 VSUBS 0.006388f
C50 B.n22 VSUBS 0.006388f
C51 B.n23 VSUBS 0.006388f
C52 B.n24 VSUBS 0.006388f
C53 B.n25 VSUBS 0.006388f
C54 B.n26 VSUBS 0.006388f
C55 B.n27 VSUBS 0.006388f
C56 B.n28 VSUBS 0.006388f
C57 B.n29 VSUBS 0.006388f
C58 B.n30 VSUBS 0.006388f
C59 B.n31 VSUBS 0.006388f
C60 B.n32 VSUBS 0.006388f
C61 B.n33 VSUBS 0.006388f
C62 B.n34 VSUBS 0.006388f
C63 B.n35 VSUBS 0.006388f
C64 B.n36 VSUBS 0.006388f
C65 B.n37 VSUBS 0.006388f
C66 B.n38 VSUBS 0.006388f
C67 B.n39 VSUBS 0.006388f
C68 B.n40 VSUBS 0.006388f
C69 B.n41 VSUBS 0.006388f
C70 B.n42 VSUBS 0.006388f
C71 B.n43 VSUBS 0.006388f
C72 B.n44 VSUBS 0.006388f
C73 B.n45 VSUBS 0.006388f
C74 B.t1 VSUBS 0.504497f
C75 B.t2 VSUBS 0.522257f
C76 B.t0 VSUBS 1.54393f
C77 B.n46 VSUBS 0.271108f
C78 B.n47 VSUBS 0.064693f
C79 B.n48 VSUBS 0.006388f
C80 B.n49 VSUBS 0.006388f
C81 B.n50 VSUBS 0.006388f
C82 B.n51 VSUBS 0.006388f
C83 B.t10 VSUBS 0.504481f
C84 B.t11 VSUBS 0.522243f
C85 B.t9 VSUBS 1.54393f
C86 B.n52 VSUBS 0.271121f
C87 B.n53 VSUBS 0.064709f
C88 B.n54 VSUBS 0.006388f
C89 B.n55 VSUBS 0.006388f
C90 B.n56 VSUBS 0.006388f
C91 B.n57 VSUBS 0.006388f
C92 B.n58 VSUBS 0.006388f
C93 B.n59 VSUBS 0.006388f
C94 B.n60 VSUBS 0.006388f
C95 B.n61 VSUBS 0.006388f
C96 B.n62 VSUBS 0.006388f
C97 B.n63 VSUBS 0.006388f
C98 B.n64 VSUBS 0.006388f
C99 B.n65 VSUBS 0.006388f
C100 B.n66 VSUBS 0.006388f
C101 B.n67 VSUBS 0.006388f
C102 B.n68 VSUBS 0.006388f
C103 B.n69 VSUBS 0.006388f
C104 B.n70 VSUBS 0.006388f
C105 B.n71 VSUBS 0.006388f
C106 B.n72 VSUBS 0.006388f
C107 B.n73 VSUBS 0.006388f
C108 B.n74 VSUBS 0.006388f
C109 B.n75 VSUBS 0.006388f
C110 B.n76 VSUBS 0.006388f
C111 B.n77 VSUBS 0.006388f
C112 B.n78 VSUBS 0.006388f
C113 B.n79 VSUBS 0.006388f
C114 B.n80 VSUBS 0.006388f
C115 B.n81 VSUBS 0.014827f
C116 B.n82 VSUBS 0.006388f
C117 B.n83 VSUBS 0.006388f
C118 B.n84 VSUBS 0.006388f
C119 B.n85 VSUBS 0.006388f
C120 B.n86 VSUBS 0.006388f
C121 B.n87 VSUBS 0.006388f
C122 B.n88 VSUBS 0.006388f
C123 B.n89 VSUBS 0.006388f
C124 B.n90 VSUBS 0.006388f
C125 B.n91 VSUBS 0.006388f
C126 B.n92 VSUBS 0.006388f
C127 B.n93 VSUBS 0.006388f
C128 B.n94 VSUBS 0.006388f
C129 B.n95 VSUBS 0.006388f
C130 B.n96 VSUBS 0.006388f
C131 B.n97 VSUBS 0.006388f
C132 B.n98 VSUBS 0.006388f
C133 B.n99 VSUBS 0.006388f
C134 B.n100 VSUBS 0.006388f
C135 B.n101 VSUBS 0.006388f
C136 B.n102 VSUBS 0.006388f
C137 B.n103 VSUBS 0.006388f
C138 B.n104 VSUBS 0.006388f
C139 B.n105 VSUBS 0.006388f
C140 B.n106 VSUBS 0.006388f
C141 B.n107 VSUBS 0.006388f
C142 B.n108 VSUBS 0.006388f
C143 B.n109 VSUBS 0.006388f
C144 B.n110 VSUBS 0.006388f
C145 B.n111 VSUBS 0.006388f
C146 B.n112 VSUBS 0.006388f
C147 B.n113 VSUBS 0.015424f
C148 B.n114 VSUBS 0.006388f
C149 B.n115 VSUBS 0.006388f
C150 B.n116 VSUBS 0.006388f
C151 B.n117 VSUBS 0.006388f
C152 B.n118 VSUBS 0.006388f
C153 B.n119 VSUBS 0.006388f
C154 B.n120 VSUBS 0.006388f
C155 B.n121 VSUBS 0.006388f
C156 B.n122 VSUBS 0.006388f
C157 B.n123 VSUBS 0.006388f
C158 B.n124 VSUBS 0.006388f
C159 B.n125 VSUBS 0.006388f
C160 B.n126 VSUBS 0.006388f
C161 B.n127 VSUBS 0.006388f
C162 B.n128 VSUBS 0.006388f
C163 B.n129 VSUBS 0.006388f
C164 B.n130 VSUBS 0.006388f
C165 B.n131 VSUBS 0.006388f
C166 B.n132 VSUBS 0.006388f
C167 B.n133 VSUBS 0.006388f
C168 B.n134 VSUBS 0.006388f
C169 B.n135 VSUBS 0.006388f
C170 B.n136 VSUBS 0.006388f
C171 B.n137 VSUBS 0.006388f
C172 B.n138 VSUBS 0.006388f
C173 B.n139 VSUBS 0.006388f
C174 B.n140 VSUBS 0.004416f
C175 B.n141 VSUBS 0.006388f
C176 B.n142 VSUBS 0.006388f
C177 B.n143 VSUBS 0.006388f
C178 B.n144 VSUBS 0.006388f
C179 B.n145 VSUBS 0.006388f
C180 B.t8 VSUBS 0.504497f
C181 B.t7 VSUBS 0.522257f
C182 B.t6 VSUBS 1.54393f
C183 B.n146 VSUBS 0.271108f
C184 B.n147 VSUBS 0.064693f
C185 B.n148 VSUBS 0.006388f
C186 B.n149 VSUBS 0.006388f
C187 B.n150 VSUBS 0.006388f
C188 B.n151 VSUBS 0.006388f
C189 B.n152 VSUBS 0.006388f
C190 B.n153 VSUBS 0.006388f
C191 B.n154 VSUBS 0.006388f
C192 B.n155 VSUBS 0.006388f
C193 B.n156 VSUBS 0.006388f
C194 B.n157 VSUBS 0.006388f
C195 B.n158 VSUBS 0.006388f
C196 B.n159 VSUBS 0.006388f
C197 B.n160 VSUBS 0.006388f
C198 B.n161 VSUBS 0.006388f
C199 B.n162 VSUBS 0.006388f
C200 B.n163 VSUBS 0.006388f
C201 B.n164 VSUBS 0.006388f
C202 B.n165 VSUBS 0.006388f
C203 B.n166 VSUBS 0.006388f
C204 B.n167 VSUBS 0.006388f
C205 B.n168 VSUBS 0.006388f
C206 B.n169 VSUBS 0.006388f
C207 B.n170 VSUBS 0.006388f
C208 B.n171 VSUBS 0.006388f
C209 B.n172 VSUBS 0.006388f
C210 B.n173 VSUBS 0.006388f
C211 B.n174 VSUBS 0.015424f
C212 B.n175 VSUBS 0.006388f
C213 B.n176 VSUBS 0.006388f
C214 B.n177 VSUBS 0.006388f
C215 B.n178 VSUBS 0.006388f
C216 B.n179 VSUBS 0.006388f
C217 B.n180 VSUBS 0.006388f
C218 B.n181 VSUBS 0.006388f
C219 B.n182 VSUBS 0.006388f
C220 B.n183 VSUBS 0.006388f
C221 B.n184 VSUBS 0.006388f
C222 B.n185 VSUBS 0.006388f
C223 B.n186 VSUBS 0.006388f
C224 B.n187 VSUBS 0.006388f
C225 B.n188 VSUBS 0.006388f
C226 B.n189 VSUBS 0.006388f
C227 B.n190 VSUBS 0.006388f
C228 B.n191 VSUBS 0.006388f
C229 B.n192 VSUBS 0.006388f
C230 B.n193 VSUBS 0.006388f
C231 B.n194 VSUBS 0.006388f
C232 B.n195 VSUBS 0.006388f
C233 B.n196 VSUBS 0.006388f
C234 B.n197 VSUBS 0.006388f
C235 B.n198 VSUBS 0.006388f
C236 B.n199 VSUBS 0.006388f
C237 B.n200 VSUBS 0.006388f
C238 B.n201 VSUBS 0.006388f
C239 B.n202 VSUBS 0.006388f
C240 B.n203 VSUBS 0.006388f
C241 B.n204 VSUBS 0.006388f
C242 B.n205 VSUBS 0.006388f
C243 B.n206 VSUBS 0.006388f
C244 B.n207 VSUBS 0.006388f
C245 B.n208 VSUBS 0.006388f
C246 B.n209 VSUBS 0.006388f
C247 B.n210 VSUBS 0.006388f
C248 B.n211 VSUBS 0.006388f
C249 B.n212 VSUBS 0.006388f
C250 B.n213 VSUBS 0.006388f
C251 B.n214 VSUBS 0.006388f
C252 B.n215 VSUBS 0.006388f
C253 B.n216 VSUBS 0.006388f
C254 B.n217 VSUBS 0.006388f
C255 B.n218 VSUBS 0.006388f
C256 B.n219 VSUBS 0.006388f
C257 B.n220 VSUBS 0.006388f
C258 B.n221 VSUBS 0.006388f
C259 B.n222 VSUBS 0.006388f
C260 B.n223 VSUBS 0.006388f
C261 B.n224 VSUBS 0.006388f
C262 B.n225 VSUBS 0.006388f
C263 B.n226 VSUBS 0.006388f
C264 B.n227 VSUBS 0.006388f
C265 B.n228 VSUBS 0.006388f
C266 B.n229 VSUBS 0.006388f
C267 B.n230 VSUBS 0.006388f
C268 B.n231 VSUBS 0.006388f
C269 B.n232 VSUBS 0.006388f
C270 B.n233 VSUBS 0.014827f
C271 B.n234 VSUBS 0.014827f
C272 B.n235 VSUBS 0.015424f
C273 B.n236 VSUBS 0.006388f
C274 B.n237 VSUBS 0.006388f
C275 B.n238 VSUBS 0.006388f
C276 B.n239 VSUBS 0.006388f
C277 B.n240 VSUBS 0.006388f
C278 B.n241 VSUBS 0.006388f
C279 B.n242 VSUBS 0.006388f
C280 B.n243 VSUBS 0.006388f
C281 B.n244 VSUBS 0.006388f
C282 B.n245 VSUBS 0.006388f
C283 B.n246 VSUBS 0.006388f
C284 B.n247 VSUBS 0.006388f
C285 B.n248 VSUBS 0.006388f
C286 B.n249 VSUBS 0.006388f
C287 B.n250 VSUBS 0.006388f
C288 B.n251 VSUBS 0.006388f
C289 B.n252 VSUBS 0.006388f
C290 B.n253 VSUBS 0.006388f
C291 B.n254 VSUBS 0.006388f
C292 B.n255 VSUBS 0.006388f
C293 B.n256 VSUBS 0.006388f
C294 B.n257 VSUBS 0.006388f
C295 B.n258 VSUBS 0.006388f
C296 B.n259 VSUBS 0.006388f
C297 B.n260 VSUBS 0.006388f
C298 B.n261 VSUBS 0.006388f
C299 B.n262 VSUBS 0.006388f
C300 B.n263 VSUBS 0.006388f
C301 B.n264 VSUBS 0.006388f
C302 B.n265 VSUBS 0.006388f
C303 B.n266 VSUBS 0.006388f
C304 B.n267 VSUBS 0.006388f
C305 B.n268 VSUBS 0.006388f
C306 B.n269 VSUBS 0.006388f
C307 B.n270 VSUBS 0.006388f
C308 B.n271 VSUBS 0.006388f
C309 B.n272 VSUBS 0.006388f
C310 B.n273 VSUBS 0.006388f
C311 B.n274 VSUBS 0.006388f
C312 B.n275 VSUBS 0.006388f
C313 B.n276 VSUBS 0.006388f
C314 B.n277 VSUBS 0.006388f
C315 B.n278 VSUBS 0.006388f
C316 B.n279 VSUBS 0.006388f
C317 B.n280 VSUBS 0.006388f
C318 B.n281 VSUBS 0.006388f
C319 B.n282 VSUBS 0.006388f
C320 B.n283 VSUBS 0.006388f
C321 B.n284 VSUBS 0.006388f
C322 B.n285 VSUBS 0.006388f
C323 B.n286 VSUBS 0.006388f
C324 B.n287 VSUBS 0.006388f
C325 B.n288 VSUBS 0.006388f
C326 B.n289 VSUBS 0.006388f
C327 B.n290 VSUBS 0.006388f
C328 B.n291 VSUBS 0.006388f
C329 B.n292 VSUBS 0.006388f
C330 B.n293 VSUBS 0.006388f
C331 B.n294 VSUBS 0.006388f
C332 B.n295 VSUBS 0.006388f
C333 B.n296 VSUBS 0.006388f
C334 B.n297 VSUBS 0.006388f
C335 B.n298 VSUBS 0.006388f
C336 B.n299 VSUBS 0.006388f
C337 B.n300 VSUBS 0.006388f
C338 B.n301 VSUBS 0.006388f
C339 B.n302 VSUBS 0.006388f
C340 B.n303 VSUBS 0.006388f
C341 B.n304 VSUBS 0.006388f
C342 B.n305 VSUBS 0.006388f
C343 B.n306 VSUBS 0.006388f
C344 B.n307 VSUBS 0.006388f
C345 B.n308 VSUBS 0.006388f
C346 B.n309 VSUBS 0.006388f
C347 B.n310 VSUBS 0.006388f
C348 B.n311 VSUBS 0.006388f
C349 B.n312 VSUBS 0.006388f
C350 B.n313 VSUBS 0.006388f
C351 B.n314 VSUBS 0.006388f
C352 B.n315 VSUBS 0.006388f
C353 B.n316 VSUBS 0.004416f
C354 B.n317 VSUBS 0.014802f
C355 B.n318 VSUBS 0.005167f
C356 B.n319 VSUBS 0.006388f
C357 B.n320 VSUBS 0.006388f
C358 B.n321 VSUBS 0.006388f
C359 B.n322 VSUBS 0.006388f
C360 B.n323 VSUBS 0.006388f
C361 B.n324 VSUBS 0.006388f
C362 B.n325 VSUBS 0.006388f
C363 B.n326 VSUBS 0.006388f
C364 B.n327 VSUBS 0.006388f
C365 B.n328 VSUBS 0.006388f
C366 B.n329 VSUBS 0.006388f
C367 B.t5 VSUBS 0.504481f
C368 B.t4 VSUBS 0.522243f
C369 B.t3 VSUBS 1.54393f
C370 B.n330 VSUBS 0.271121f
C371 B.n331 VSUBS 0.064709f
C372 B.n332 VSUBS 0.014802f
C373 B.n333 VSUBS 0.005167f
C374 B.n334 VSUBS 0.006388f
C375 B.n335 VSUBS 0.006388f
C376 B.n336 VSUBS 0.006388f
C377 B.n337 VSUBS 0.006388f
C378 B.n338 VSUBS 0.006388f
C379 B.n339 VSUBS 0.006388f
C380 B.n340 VSUBS 0.006388f
C381 B.n341 VSUBS 0.006388f
C382 B.n342 VSUBS 0.006388f
C383 B.n343 VSUBS 0.006388f
C384 B.n344 VSUBS 0.006388f
C385 B.n345 VSUBS 0.006388f
C386 B.n346 VSUBS 0.006388f
C387 B.n347 VSUBS 0.006388f
C388 B.n348 VSUBS 0.006388f
C389 B.n349 VSUBS 0.006388f
C390 B.n350 VSUBS 0.006388f
C391 B.n351 VSUBS 0.006388f
C392 B.n352 VSUBS 0.006388f
C393 B.n353 VSUBS 0.006388f
C394 B.n354 VSUBS 0.006388f
C395 B.n355 VSUBS 0.006388f
C396 B.n356 VSUBS 0.006388f
C397 B.n357 VSUBS 0.006388f
C398 B.n358 VSUBS 0.006388f
C399 B.n359 VSUBS 0.006388f
C400 B.n360 VSUBS 0.006388f
C401 B.n361 VSUBS 0.006388f
C402 B.n362 VSUBS 0.006388f
C403 B.n363 VSUBS 0.006388f
C404 B.n364 VSUBS 0.006388f
C405 B.n365 VSUBS 0.006388f
C406 B.n366 VSUBS 0.006388f
C407 B.n367 VSUBS 0.006388f
C408 B.n368 VSUBS 0.006388f
C409 B.n369 VSUBS 0.006388f
C410 B.n370 VSUBS 0.006388f
C411 B.n371 VSUBS 0.006388f
C412 B.n372 VSUBS 0.006388f
C413 B.n373 VSUBS 0.006388f
C414 B.n374 VSUBS 0.006388f
C415 B.n375 VSUBS 0.006388f
C416 B.n376 VSUBS 0.006388f
C417 B.n377 VSUBS 0.006388f
C418 B.n378 VSUBS 0.006388f
C419 B.n379 VSUBS 0.006388f
C420 B.n380 VSUBS 0.006388f
C421 B.n381 VSUBS 0.006388f
C422 B.n382 VSUBS 0.006388f
C423 B.n383 VSUBS 0.006388f
C424 B.n384 VSUBS 0.006388f
C425 B.n385 VSUBS 0.006388f
C426 B.n386 VSUBS 0.006388f
C427 B.n387 VSUBS 0.006388f
C428 B.n388 VSUBS 0.006388f
C429 B.n389 VSUBS 0.006388f
C430 B.n390 VSUBS 0.006388f
C431 B.n391 VSUBS 0.006388f
C432 B.n392 VSUBS 0.006388f
C433 B.n393 VSUBS 0.006388f
C434 B.n394 VSUBS 0.006388f
C435 B.n395 VSUBS 0.006388f
C436 B.n396 VSUBS 0.006388f
C437 B.n397 VSUBS 0.006388f
C438 B.n398 VSUBS 0.006388f
C439 B.n399 VSUBS 0.006388f
C440 B.n400 VSUBS 0.006388f
C441 B.n401 VSUBS 0.006388f
C442 B.n402 VSUBS 0.006388f
C443 B.n403 VSUBS 0.006388f
C444 B.n404 VSUBS 0.006388f
C445 B.n405 VSUBS 0.006388f
C446 B.n406 VSUBS 0.006388f
C447 B.n407 VSUBS 0.006388f
C448 B.n408 VSUBS 0.006388f
C449 B.n409 VSUBS 0.006388f
C450 B.n410 VSUBS 0.006388f
C451 B.n411 VSUBS 0.006388f
C452 B.n412 VSUBS 0.006388f
C453 B.n413 VSUBS 0.006388f
C454 B.n414 VSUBS 0.006388f
C455 B.n415 VSUBS 0.006388f
C456 B.n416 VSUBS 0.014683f
C457 B.n417 VSUBS 0.015569f
C458 B.n418 VSUBS 0.014827f
C459 B.n419 VSUBS 0.006388f
C460 B.n420 VSUBS 0.006388f
C461 B.n421 VSUBS 0.006388f
C462 B.n422 VSUBS 0.006388f
C463 B.n423 VSUBS 0.006388f
C464 B.n424 VSUBS 0.006388f
C465 B.n425 VSUBS 0.006388f
C466 B.n426 VSUBS 0.006388f
C467 B.n427 VSUBS 0.006388f
C468 B.n428 VSUBS 0.006388f
C469 B.n429 VSUBS 0.006388f
C470 B.n430 VSUBS 0.006388f
C471 B.n431 VSUBS 0.006388f
C472 B.n432 VSUBS 0.006388f
C473 B.n433 VSUBS 0.006388f
C474 B.n434 VSUBS 0.006388f
C475 B.n435 VSUBS 0.006388f
C476 B.n436 VSUBS 0.006388f
C477 B.n437 VSUBS 0.006388f
C478 B.n438 VSUBS 0.006388f
C479 B.n439 VSUBS 0.006388f
C480 B.n440 VSUBS 0.006388f
C481 B.n441 VSUBS 0.006388f
C482 B.n442 VSUBS 0.006388f
C483 B.n443 VSUBS 0.006388f
C484 B.n444 VSUBS 0.006388f
C485 B.n445 VSUBS 0.006388f
C486 B.n446 VSUBS 0.006388f
C487 B.n447 VSUBS 0.006388f
C488 B.n448 VSUBS 0.006388f
C489 B.n449 VSUBS 0.006388f
C490 B.n450 VSUBS 0.006388f
C491 B.n451 VSUBS 0.006388f
C492 B.n452 VSUBS 0.006388f
C493 B.n453 VSUBS 0.006388f
C494 B.n454 VSUBS 0.006388f
C495 B.n455 VSUBS 0.006388f
C496 B.n456 VSUBS 0.006388f
C497 B.n457 VSUBS 0.006388f
C498 B.n458 VSUBS 0.006388f
C499 B.n459 VSUBS 0.006388f
C500 B.n460 VSUBS 0.006388f
C501 B.n461 VSUBS 0.006388f
C502 B.n462 VSUBS 0.006388f
C503 B.n463 VSUBS 0.006388f
C504 B.n464 VSUBS 0.006388f
C505 B.n465 VSUBS 0.006388f
C506 B.n466 VSUBS 0.006388f
C507 B.n467 VSUBS 0.006388f
C508 B.n468 VSUBS 0.006388f
C509 B.n469 VSUBS 0.006388f
C510 B.n470 VSUBS 0.006388f
C511 B.n471 VSUBS 0.006388f
C512 B.n472 VSUBS 0.006388f
C513 B.n473 VSUBS 0.006388f
C514 B.n474 VSUBS 0.006388f
C515 B.n475 VSUBS 0.006388f
C516 B.n476 VSUBS 0.006388f
C517 B.n477 VSUBS 0.006388f
C518 B.n478 VSUBS 0.006388f
C519 B.n479 VSUBS 0.006388f
C520 B.n480 VSUBS 0.006388f
C521 B.n481 VSUBS 0.006388f
C522 B.n482 VSUBS 0.006388f
C523 B.n483 VSUBS 0.006388f
C524 B.n484 VSUBS 0.006388f
C525 B.n485 VSUBS 0.006388f
C526 B.n486 VSUBS 0.006388f
C527 B.n487 VSUBS 0.006388f
C528 B.n488 VSUBS 0.006388f
C529 B.n489 VSUBS 0.006388f
C530 B.n490 VSUBS 0.006388f
C531 B.n491 VSUBS 0.006388f
C532 B.n492 VSUBS 0.006388f
C533 B.n493 VSUBS 0.006388f
C534 B.n494 VSUBS 0.006388f
C535 B.n495 VSUBS 0.006388f
C536 B.n496 VSUBS 0.006388f
C537 B.n497 VSUBS 0.006388f
C538 B.n498 VSUBS 0.006388f
C539 B.n499 VSUBS 0.006388f
C540 B.n500 VSUBS 0.006388f
C541 B.n501 VSUBS 0.006388f
C542 B.n502 VSUBS 0.006388f
C543 B.n503 VSUBS 0.006388f
C544 B.n504 VSUBS 0.006388f
C545 B.n505 VSUBS 0.006388f
C546 B.n506 VSUBS 0.006388f
C547 B.n507 VSUBS 0.006388f
C548 B.n508 VSUBS 0.006388f
C549 B.n509 VSUBS 0.006388f
C550 B.n510 VSUBS 0.006388f
C551 B.n511 VSUBS 0.006388f
C552 B.n512 VSUBS 0.014827f
C553 B.n513 VSUBS 0.015424f
C554 B.n514 VSUBS 0.015424f
C555 B.n515 VSUBS 0.006388f
C556 B.n516 VSUBS 0.006388f
C557 B.n517 VSUBS 0.006388f
C558 B.n518 VSUBS 0.006388f
C559 B.n519 VSUBS 0.006388f
C560 B.n520 VSUBS 0.006388f
C561 B.n521 VSUBS 0.006388f
C562 B.n522 VSUBS 0.006388f
C563 B.n523 VSUBS 0.006388f
C564 B.n524 VSUBS 0.006388f
C565 B.n525 VSUBS 0.006388f
C566 B.n526 VSUBS 0.006388f
C567 B.n527 VSUBS 0.006388f
C568 B.n528 VSUBS 0.006388f
C569 B.n529 VSUBS 0.006388f
C570 B.n530 VSUBS 0.006388f
C571 B.n531 VSUBS 0.006388f
C572 B.n532 VSUBS 0.006388f
C573 B.n533 VSUBS 0.006388f
C574 B.n534 VSUBS 0.006388f
C575 B.n535 VSUBS 0.006388f
C576 B.n536 VSUBS 0.006388f
C577 B.n537 VSUBS 0.006388f
C578 B.n538 VSUBS 0.006388f
C579 B.n539 VSUBS 0.006388f
C580 B.n540 VSUBS 0.006388f
C581 B.n541 VSUBS 0.006388f
C582 B.n542 VSUBS 0.006388f
C583 B.n543 VSUBS 0.006388f
C584 B.n544 VSUBS 0.006388f
C585 B.n545 VSUBS 0.006388f
C586 B.n546 VSUBS 0.006388f
C587 B.n547 VSUBS 0.006388f
C588 B.n548 VSUBS 0.006388f
C589 B.n549 VSUBS 0.006388f
C590 B.n550 VSUBS 0.006388f
C591 B.n551 VSUBS 0.006388f
C592 B.n552 VSUBS 0.006388f
C593 B.n553 VSUBS 0.006388f
C594 B.n554 VSUBS 0.006388f
C595 B.n555 VSUBS 0.006388f
C596 B.n556 VSUBS 0.006388f
C597 B.n557 VSUBS 0.006388f
C598 B.n558 VSUBS 0.006388f
C599 B.n559 VSUBS 0.006388f
C600 B.n560 VSUBS 0.006388f
C601 B.n561 VSUBS 0.006388f
C602 B.n562 VSUBS 0.006388f
C603 B.n563 VSUBS 0.006388f
C604 B.n564 VSUBS 0.006388f
C605 B.n565 VSUBS 0.006388f
C606 B.n566 VSUBS 0.006388f
C607 B.n567 VSUBS 0.006388f
C608 B.n568 VSUBS 0.006388f
C609 B.n569 VSUBS 0.006388f
C610 B.n570 VSUBS 0.006388f
C611 B.n571 VSUBS 0.006388f
C612 B.n572 VSUBS 0.006388f
C613 B.n573 VSUBS 0.006388f
C614 B.n574 VSUBS 0.006388f
C615 B.n575 VSUBS 0.006388f
C616 B.n576 VSUBS 0.006388f
C617 B.n577 VSUBS 0.006388f
C618 B.n578 VSUBS 0.006388f
C619 B.n579 VSUBS 0.006388f
C620 B.n580 VSUBS 0.006388f
C621 B.n581 VSUBS 0.006388f
C622 B.n582 VSUBS 0.006388f
C623 B.n583 VSUBS 0.006388f
C624 B.n584 VSUBS 0.006388f
C625 B.n585 VSUBS 0.006388f
C626 B.n586 VSUBS 0.006388f
C627 B.n587 VSUBS 0.006388f
C628 B.n588 VSUBS 0.006388f
C629 B.n589 VSUBS 0.006388f
C630 B.n590 VSUBS 0.006388f
C631 B.n591 VSUBS 0.006388f
C632 B.n592 VSUBS 0.006388f
C633 B.n593 VSUBS 0.006388f
C634 B.n594 VSUBS 0.006388f
C635 B.n595 VSUBS 0.004416f
C636 B.n596 VSUBS 0.014802f
C637 B.n597 VSUBS 0.005167f
C638 B.n598 VSUBS 0.006388f
C639 B.n599 VSUBS 0.006388f
C640 B.n600 VSUBS 0.006388f
C641 B.n601 VSUBS 0.006388f
C642 B.n602 VSUBS 0.006388f
C643 B.n603 VSUBS 0.006388f
C644 B.n604 VSUBS 0.006388f
C645 B.n605 VSUBS 0.006388f
C646 B.n606 VSUBS 0.006388f
C647 B.n607 VSUBS 0.006388f
C648 B.n608 VSUBS 0.006388f
C649 B.n609 VSUBS 0.005167f
C650 B.n610 VSUBS 0.014802f
C651 B.n611 VSUBS 0.004416f
C652 B.n612 VSUBS 0.006388f
C653 B.n613 VSUBS 0.006388f
C654 B.n614 VSUBS 0.006388f
C655 B.n615 VSUBS 0.006388f
C656 B.n616 VSUBS 0.006388f
C657 B.n617 VSUBS 0.006388f
C658 B.n618 VSUBS 0.006388f
C659 B.n619 VSUBS 0.006388f
C660 B.n620 VSUBS 0.006388f
C661 B.n621 VSUBS 0.006388f
C662 B.n622 VSUBS 0.006388f
C663 B.n623 VSUBS 0.006388f
C664 B.n624 VSUBS 0.006388f
C665 B.n625 VSUBS 0.006388f
C666 B.n626 VSUBS 0.006388f
C667 B.n627 VSUBS 0.006388f
C668 B.n628 VSUBS 0.006388f
C669 B.n629 VSUBS 0.006388f
C670 B.n630 VSUBS 0.006388f
C671 B.n631 VSUBS 0.006388f
C672 B.n632 VSUBS 0.006388f
C673 B.n633 VSUBS 0.006388f
C674 B.n634 VSUBS 0.006388f
C675 B.n635 VSUBS 0.006388f
C676 B.n636 VSUBS 0.006388f
C677 B.n637 VSUBS 0.006388f
C678 B.n638 VSUBS 0.006388f
C679 B.n639 VSUBS 0.006388f
C680 B.n640 VSUBS 0.006388f
C681 B.n641 VSUBS 0.006388f
C682 B.n642 VSUBS 0.006388f
C683 B.n643 VSUBS 0.006388f
C684 B.n644 VSUBS 0.006388f
C685 B.n645 VSUBS 0.006388f
C686 B.n646 VSUBS 0.006388f
C687 B.n647 VSUBS 0.006388f
C688 B.n648 VSUBS 0.006388f
C689 B.n649 VSUBS 0.006388f
C690 B.n650 VSUBS 0.006388f
C691 B.n651 VSUBS 0.006388f
C692 B.n652 VSUBS 0.006388f
C693 B.n653 VSUBS 0.006388f
C694 B.n654 VSUBS 0.006388f
C695 B.n655 VSUBS 0.006388f
C696 B.n656 VSUBS 0.006388f
C697 B.n657 VSUBS 0.006388f
C698 B.n658 VSUBS 0.006388f
C699 B.n659 VSUBS 0.006388f
C700 B.n660 VSUBS 0.006388f
C701 B.n661 VSUBS 0.006388f
C702 B.n662 VSUBS 0.006388f
C703 B.n663 VSUBS 0.006388f
C704 B.n664 VSUBS 0.006388f
C705 B.n665 VSUBS 0.006388f
C706 B.n666 VSUBS 0.006388f
C707 B.n667 VSUBS 0.006388f
C708 B.n668 VSUBS 0.006388f
C709 B.n669 VSUBS 0.006388f
C710 B.n670 VSUBS 0.006388f
C711 B.n671 VSUBS 0.006388f
C712 B.n672 VSUBS 0.006388f
C713 B.n673 VSUBS 0.006388f
C714 B.n674 VSUBS 0.006388f
C715 B.n675 VSUBS 0.006388f
C716 B.n676 VSUBS 0.006388f
C717 B.n677 VSUBS 0.006388f
C718 B.n678 VSUBS 0.006388f
C719 B.n679 VSUBS 0.006388f
C720 B.n680 VSUBS 0.006388f
C721 B.n681 VSUBS 0.006388f
C722 B.n682 VSUBS 0.006388f
C723 B.n683 VSUBS 0.006388f
C724 B.n684 VSUBS 0.006388f
C725 B.n685 VSUBS 0.006388f
C726 B.n686 VSUBS 0.006388f
C727 B.n687 VSUBS 0.006388f
C728 B.n688 VSUBS 0.006388f
C729 B.n689 VSUBS 0.006388f
C730 B.n690 VSUBS 0.006388f
C731 B.n691 VSUBS 0.006388f
C732 B.n692 VSUBS 0.015424f
C733 B.n693 VSUBS 0.015424f
C734 B.n694 VSUBS 0.014827f
C735 B.n695 VSUBS 0.006388f
C736 B.n696 VSUBS 0.006388f
C737 B.n697 VSUBS 0.006388f
C738 B.n698 VSUBS 0.006388f
C739 B.n699 VSUBS 0.006388f
C740 B.n700 VSUBS 0.006388f
C741 B.n701 VSUBS 0.006388f
C742 B.n702 VSUBS 0.006388f
C743 B.n703 VSUBS 0.006388f
C744 B.n704 VSUBS 0.006388f
C745 B.n705 VSUBS 0.006388f
C746 B.n706 VSUBS 0.006388f
C747 B.n707 VSUBS 0.006388f
C748 B.n708 VSUBS 0.006388f
C749 B.n709 VSUBS 0.006388f
C750 B.n710 VSUBS 0.006388f
C751 B.n711 VSUBS 0.006388f
C752 B.n712 VSUBS 0.006388f
C753 B.n713 VSUBS 0.006388f
C754 B.n714 VSUBS 0.006388f
C755 B.n715 VSUBS 0.006388f
C756 B.n716 VSUBS 0.006388f
C757 B.n717 VSUBS 0.006388f
C758 B.n718 VSUBS 0.006388f
C759 B.n719 VSUBS 0.006388f
C760 B.n720 VSUBS 0.006388f
C761 B.n721 VSUBS 0.006388f
C762 B.n722 VSUBS 0.006388f
C763 B.n723 VSUBS 0.006388f
C764 B.n724 VSUBS 0.006388f
C765 B.n725 VSUBS 0.006388f
C766 B.n726 VSUBS 0.006388f
C767 B.n727 VSUBS 0.006388f
C768 B.n728 VSUBS 0.006388f
C769 B.n729 VSUBS 0.006388f
C770 B.n730 VSUBS 0.006388f
C771 B.n731 VSUBS 0.006388f
C772 B.n732 VSUBS 0.006388f
C773 B.n733 VSUBS 0.006388f
C774 B.n734 VSUBS 0.006388f
C775 B.n735 VSUBS 0.006388f
C776 B.n736 VSUBS 0.006388f
C777 B.n737 VSUBS 0.006388f
C778 B.n738 VSUBS 0.006388f
C779 B.n739 VSUBS 0.008337f
C780 B.n740 VSUBS 0.008881f
C781 B.n741 VSUBS 0.01766f
C782 VDD1.t1 VSUBS 0.347833f
C783 VDD1.t3 VSUBS 0.347833f
C784 VDD1.n0 VSUBS 2.86135f
C785 VDD1.t2 VSUBS 0.347833f
C786 VDD1.t0 VSUBS 0.347833f
C787 VDD1.n1 VSUBS 3.76053f
C788 VP.n0 VSUBS 0.043935f
C789 VP.t3 VSUBS 3.49867f
C790 VP.n1 VSUBS 0.026917f
C791 VP.n2 VSUBS 0.043935f
C792 VP.t1 VSUBS 3.49867f
C793 VP.t0 VSUBS 3.74383f
C794 VP.t2 VSUBS 3.74825f
C795 VP.n3 VSUBS 4.2936f
C796 VP.n4 VSUBS 2.01886f
C797 VP.n5 VSUBS 1.33036f
C798 VP.n6 VSUBS 0.051123f
C799 VP.n7 VSUBS 0.065888f
C800 VP.n8 VSUBS 0.033327f
C801 VP.n9 VSUBS 0.033327f
C802 VP.n10 VSUBS 0.033327f
C803 VP.n11 VSUBS 0.065888f
C804 VP.n12 VSUBS 0.051123f
C805 VP.n13 VSUBS 1.33036f
C806 VP.n14 VSUBS 0.046276f
C807 VTAIL.t5 VSUBS 2.962f
C808 VTAIL.n0 VSUBS 0.754769f
C809 VTAIL.t0 VSUBS 2.962f
C810 VTAIL.n1 VSUBS 0.832979f
C811 VTAIL.t7 VSUBS 2.962f
C812 VTAIL.n2 VSUBS 2.29301f
C813 VTAIL.t6 VSUBS 2.96201f
C814 VTAIL.n3 VSUBS 2.29301f
C815 VTAIL.t4 VSUBS 2.96201f
C816 VTAIL.n4 VSUBS 0.832974f
C817 VTAIL.t1 VSUBS 2.96201f
C818 VTAIL.n5 VSUBS 0.832974f
C819 VTAIL.t2 VSUBS 2.962f
C820 VTAIL.n6 VSUBS 2.29301f
C821 VTAIL.t3 VSUBS 2.962f
C822 VTAIL.n7 VSUBS 2.20641f
C823 VDD2.t1 VSUBS 0.345101f
C824 VDD2.t3 VSUBS 0.345101f
C825 VDD2.n0 VSUBS 3.7043f
C826 VDD2.t0 VSUBS 0.345101f
C827 VDD2.t2 VSUBS 0.345101f
C828 VDD2.n1 VSUBS 2.83828f
C829 VDD2.n2 VSUBS 4.67625f
C830 VN.t1 VSUBS 3.64743f
C831 VN.t3 VSUBS 3.64313f
C832 VN.n0 VSUBS 2.38382f
C833 VN.t2 VSUBS 3.64743f
C834 VN.t0 VSUBS 3.64313f
C835 VN.n1 VSUBS 4.19488f
.ends

