* NGSPICE file created from diff_pair_sample_1578.ext - technology: sky130A

.subckt diff_pair_sample_1578 VTAIL VN VP B VDD2 VDD1
X0 B.t19 B.t17 B.t18 B.t14 sky130_fd_pr__nfet_01v8 ad=1.3572 pd=7.74 as=0 ps=0 w=3.48 l=2.77
X1 VDD1.t5 VP.t0 VTAIL.t11 B.t0 sky130_fd_pr__nfet_01v8 ad=0.5742 pd=3.81 as=1.3572 ps=7.74 w=3.48 l=2.77
X2 VDD2.t5 VN.t0 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=1.3572 pd=7.74 as=0.5742 ps=3.81 w=3.48 l=2.77
X3 VDD2.t4 VN.t1 VTAIL.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=1.3572 pd=7.74 as=0.5742 ps=3.81 w=3.48 l=2.77
X4 B.t16 B.t13 B.t15 B.t14 sky130_fd_pr__nfet_01v8 ad=1.3572 pd=7.74 as=0 ps=0 w=3.48 l=2.77
X5 VTAIL.t8 VP.t1 VDD1.t4 B.t1 sky130_fd_pr__nfet_01v8 ad=0.5742 pd=3.81 as=0.5742 ps=3.81 w=3.48 l=2.77
X6 VTAIL.t5 VN.t2 VDD2.t3 B.t5 sky130_fd_pr__nfet_01v8 ad=0.5742 pd=3.81 as=0.5742 ps=3.81 w=3.48 l=2.77
X7 B.t12 B.t10 B.t11 B.t7 sky130_fd_pr__nfet_01v8 ad=1.3572 pd=7.74 as=0 ps=0 w=3.48 l=2.77
X8 VDD2.t2 VN.t3 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=0.5742 pd=3.81 as=1.3572 ps=7.74 w=3.48 l=2.77
X9 VTAIL.t1 VN.t4 VDD2.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=0.5742 pd=3.81 as=0.5742 ps=3.81 w=3.48 l=2.77
X10 VDD1.t3 VP.t2 VTAIL.t6 B.t4 sky130_fd_pr__nfet_01v8 ad=1.3572 pd=7.74 as=0.5742 ps=3.81 w=3.48 l=2.77
X11 VDD1.t2 VP.t3 VTAIL.t7 B.t3 sky130_fd_pr__nfet_01v8 ad=1.3572 pd=7.74 as=0.5742 ps=3.81 w=3.48 l=2.77
X12 B.t9 B.t6 B.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=1.3572 pd=7.74 as=0 ps=0 w=3.48 l=2.77
X13 VDD2.t0 VN.t5 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=0.5742 pd=3.81 as=1.3572 ps=7.74 w=3.48 l=2.77
X14 VTAIL.t9 VP.t4 VDD1.t1 B.t5 sky130_fd_pr__nfet_01v8 ad=0.5742 pd=3.81 as=0.5742 ps=3.81 w=3.48 l=2.77
X15 VDD1.t0 VP.t5 VTAIL.t10 B.t2 sky130_fd_pr__nfet_01v8 ad=0.5742 pd=3.81 as=1.3572 ps=7.74 w=3.48 l=2.77
R0 B.n583 B.n582 585
R1 B.n584 B.n583 585
R2 B.n192 B.n105 585
R3 B.n191 B.n190 585
R4 B.n189 B.n188 585
R5 B.n187 B.n186 585
R6 B.n185 B.n184 585
R7 B.n183 B.n182 585
R8 B.n181 B.n180 585
R9 B.n179 B.n178 585
R10 B.n177 B.n176 585
R11 B.n175 B.n174 585
R12 B.n173 B.n172 585
R13 B.n171 B.n170 585
R14 B.n169 B.n168 585
R15 B.n167 B.n166 585
R16 B.n165 B.n164 585
R17 B.n163 B.n162 585
R18 B.n161 B.n160 585
R19 B.n159 B.n158 585
R20 B.n157 B.n156 585
R21 B.n155 B.n154 585
R22 B.n153 B.n152 585
R23 B.n151 B.n150 585
R24 B.n149 B.n148 585
R25 B.n147 B.n146 585
R26 B.n145 B.n144 585
R27 B.n142 B.n141 585
R28 B.n140 B.n139 585
R29 B.n138 B.n137 585
R30 B.n136 B.n135 585
R31 B.n134 B.n133 585
R32 B.n132 B.n131 585
R33 B.n130 B.n129 585
R34 B.n128 B.n127 585
R35 B.n126 B.n125 585
R36 B.n124 B.n123 585
R37 B.n122 B.n121 585
R38 B.n120 B.n119 585
R39 B.n118 B.n117 585
R40 B.n116 B.n115 585
R41 B.n114 B.n113 585
R42 B.n112 B.n111 585
R43 B.n82 B.n81 585
R44 B.n581 B.n83 585
R45 B.n585 B.n83 585
R46 B.n580 B.n579 585
R47 B.n579 B.n79 585
R48 B.n578 B.n78 585
R49 B.n591 B.n78 585
R50 B.n577 B.n77 585
R51 B.n592 B.n77 585
R52 B.n576 B.n76 585
R53 B.n593 B.n76 585
R54 B.n575 B.n574 585
R55 B.n574 B.n72 585
R56 B.n573 B.n71 585
R57 B.n599 B.n71 585
R58 B.n572 B.n70 585
R59 B.n600 B.n70 585
R60 B.n571 B.n69 585
R61 B.n601 B.n69 585
R62 B.n570 B.n569 585
R63 B.n569 B.n65 585
R64 B.n568 B.n64 585
R65 B.n607 B.n64 585
R66 B.n567 B.n63 585
R67 B.n608 B.n63 585
R68 B.n566 B.n62 585
R69 B.n609 B.n62 585
R70 B.n565 B.n564 585
R71 B.n564 B.n58 585
R72 B.n563 B.n57 585
R73 B.n615 B.n57 585
R74 B.n562 B.n56 585
R75 B.n616 B.n56 585
R76 B.n561 B.n55 585
R77 B.n617 B.n55 585
R78 B.n560 B.n559 585
R79 B.n559 B.n51 585
R80 B.n558 B.n50 585
R81 B.n623 B.n50 585
R82 B.n557 B.n49 585
R83 B.n624 B.n49 585
R84 B.n556 B.n48 585
R85 B.n625 B.n48 585
R86 B.n555 B.n554 585
R87 B.n554 B.n44 585
R88 B.n553 B.n43 585
R89 B.n631 B.n43 585
R90 B.n552 B.n42 585
R91 B.n632 B.n42 585
R92 B.n551 B.n41 585
R93 B.n633 B.n41 585
R94 B.n550 B.n549 585
R95 B.n549 B.n37 585
R96 B.n548 B.n36 585
R97 B.n639 B.n36 585
R98 B.n547 B.n35 585
R99 B.n640 B.n35 585
R100 B.n546 B.n34 585
R101 B.n641 B.n34 585
R102 B.n545 B.n544 585
R103 B.n544 B.n33 585
R104 B.n543 B.n29 585
R105 B.n647 B.n29 585
R106 B.n542 B.n28 585
R107 B.n648 B.n28 585
R108 B.n541 B.n27 585
R109 B.n649 B.n27 585
R110 B.n540 B.n539 585
R111 B.n539 B.n23 585
R112 B.n538 B.n22 585
R113 B.n655 B.n22 585
R114 B.n537 B.n21 585
R115 B.n656 B.n21 585
R116 B.n536 B.n20 585
R117 B.n657 B.n20 585
R118 B.n535 B.n534 585
R119 B.n534 B.n16 585
R120 B.n533 B.n15 585
R121 B.n663 B.n15 585
R122 B.n532 B.n14 585
R123 B.n664 B.n14 585
R124 B.n531 B.n13 585
R125 B.n665 B.n13 585
R126 B.n530 B.n529 585
R127 B.n529 B.n12 585
R128 B.n528 B.n527 585
R129 B.n528 B.n8 585
R130 B.n526 B.n7 585
R131 B.n672 B.n7 585
R132 B.n525 B.n6 585
R133 B.n673 B.n6 585
R134 B.n524 B.n5 585
R135 B.n674 B.n5 585
R136 B.n523 B.n522 585
R137 B.n522 B.n4 585
R138 B.n521 B.n193 585
R139 B.n521 B.n520 585
R140 B.n511 B.n194 585
R141 B.n195 B.n194 585
R142 B.n513 B.n512 585
R143 B.n514 B.n513 585
R144 B.n510 B.n200 585
R145 B.n200 B.n199 585
R146 B.n509 B.n508 585
R147 B.n508 B.n507 585
R148 B.n202 B.n201 585
R149 B.n203 B.n202 585
R150 B.n500 B.n499 585
R151 B.n501 B.n500 585
R152 B.n498 B.n208 585
R153 B.n208 B.n207 585
R154 B.n497 B.n496 585
R155 B.n496 B.n495 585
R156 B.n210 B.n209 585
R157 B.n211 B.n210 585
R158 B.n488 B.n487 585
R159 B.n489 B.n488 585
R160 B.n486 B.n216 585
R161 B.n216 B.n215 585
R162 B.n485 B.n484 585
R163 B.n484 B.n483 585
R164 B.n218 B.n217 585
R165 B.n476 B.n218 585
R166 B.n475 B.n474 585
R167 B.n477 B.n475 585
R168 B.n473 B.n223 585
R169 B.n223 B.n222 585
R170 B.n472 B.n471 585
R171 B.n471 B.n470 585
R172 B.n225 B.n224 585
R173 B.n226 B.n225 585
R174 B.n463 B.n462 585
R175 B.n464 B.n463 585
R176 B.n461 B.n231 585
R177 B.n231 B.n230 585
R178 B.n460 B.n459 585
R179 B.n459 B.n458 585
R180 B.n233 B.n232 585
R181 B.n234 B.n233 585
R182 B.n451 B.n450 585
R183 B.n452 B.n451 585
R184 B.n449 B.n239 585
R185 B.n239 B.n238 585
R186 B.n448 B.n447 585
R187 B.n447 B.n446 585
R188 B.n241 B.n240 585
R189 B.n242 B.n241 585
R190 B.n439 B.n438 585
R191 B.n440 B.n439 585
R192 B.n437 B.n247 585
R193 B.n247 B.n246 585
R194 B.n436 B.n435 585
R195 B.n435 B.n434 585
R196 B.n249 B.n248 585
R197 B.n250 B.n249 585
R198 B.n427 B.n426 585
R199 B.n428 B.n427 585
R200 B.n425 B.n255 585
R201 B.n255 B.n254 585
R202 B.n424 B.n423 585
R203 B.n423 B.n422 585
R204 B.n257 B.n256 585
R205 B.n258 B.n257 585
R206 B.n415 B.n414 585
R207 B.n416 B.n415 585
R208 B.n413 B.n262 585
R209 B.n266 B.n262 585
R210 B.n412 B.n411 585
R211 B.n411 B.n410 585
R212 B.n264 B.n263 585
R213 B.n265 B.n264 585
R214 B.n403 B.n402 585
R215 B.n404 B.n403 585
R216 B.n401 B.n271 585
R217 B.n271 B.n270 585
R218 B.n400 B.n399 585
R219 B.n399 B.n398 585
R220 B.n273 B.n272 585
R221 B.n274 B.n273 585
R222 B.n391 B.n390 585
R223 B.n392 B.n391 585
R224 B.n277 B.n276 585
R225 B.n307 B.n306 585
R226 B.n308 B.n304 585
R227 B.n304 B.n278 585
R228 B.n310 B.n309 585
R229 B.n312 B.n303 585
R230 B.n315 B.n314 585
R231 B.n316 B.n302 585
R232 B.n318 B.n317 585
R233 B.n320 B.n301 585
R234 B.n323 B.n322 585
R235 B.n324 B.n300 585
R236 B.n326 B.n325 585
R237 B.n328 B.n299 585
R238 B.n331 B.n330 585
R239 B.n332 B.n298 585
R240 B.n334 B.n333 585
R241 B.n336 B.n297 585
R242 B.n339 B.n338 585
R243 B.n340 B.n293 585
R244 B.n342 B.n341 585
R245 B.n344 B.n292 585
R246 B.n347 B.n346 585
R247 B.n348 B.n291 585
R248 B.n350 B.n349 585
R249 B.n352 B.n290 585
R250 B.n355 B.n354 585
R251 B.n357 B.n287 585
R252 B.n359 B.n358 585
R253 B.n361 B.n286 585
R254 B.n364 B.n363 585
R255 B.n365 B.n285 585
R256 B.n367 B.n366 585
R257 B.n369 B.n284 585
R258 B.n372 B.n371 585
R259 B.n373 B.n283 585
R260 B.n375 B.n374 585
R261 B.n377 B.n282 585
R262 B.n380 B.n379 585
R263 B.n381 B.n281 585
R264 B.n383 B.n382 585
R265 B.n385 B.n280 585
R266 B.n388 B.n387 585
R267 B.n389 B.n279 585
R268 B.n394 B.n393 585
R269 B.n393 B.n392 585
R270 B.n395 B.n275 585
R271 B.n275 B.n274 585
R272 B.n397 B.n396 585
R273 B.n398 B.n397 585
R274 B.n269 B.n268 585
R275 B.n270 B.n269 585
R276 B.n406 B.n405 585
R277 B.n405 B.n404 585
R278 B.n407 B.n267 585
R279 B.n267 B.n265 585
R280 B.n409 B.n408 585
R281 B.n410 B.n409 585
R282 B.n261 B.n260 585
R283 B.n266 B.n261 585
R284 B.n418 B.n417 585
R285 B.n417 B.n416 585
R286 B.n419 B.n259 585
R287 B.n259 B.n258 585
R288 B.n421 B.n420 585
R289 B.n422 B.n421 585
R290 B.n253 B.n252 585
R291 B.n254 B.n253 585
R292 B.n430 B.n429 585
R293 B.n429 B.n428 585
R294 B.n431 B.n251 585
R295 B.n251 B.n250 585
R296 B.n433 B.n432 585
R297 B.n434 B.n433 585
R298 B.n245 B.n244 585
R299 B.n246 B.n245 585
R300 B.n442 B.n441 585
R301 B.n441 B.n440 585
R302 B.n443 B.n243 585
R303 B.n243 B.n242 585
R304 B.n445 B.n444 585
R305 B.n446 B.n445 585
R306 B.n237 B.n236 585
R307 B.n238 B.n237 585
R308 B.n454 B.n453 585
R309 B.n453 B.n452 585
R310 B.n455 B.n235 585
R311 B.n235 B.n234 585
R312 B.n457 B.n456 585
R313 B.n458 B.n457 585
R314 B.n229 B.n228 585
R315 B.n230 B.n229 585
R316 B.n466 B.n465 585
R317 B.n465 B.n464 585
R318 B.n467 B.n227 585
R319 B.n227 B.n226 585
R320 B.n469 B.n468 585
R321 B.n470 B.n469 585
R322 B.n221 B.n220 585
R323 B.n222 B.n221 585
R324 B.n479 B.n478 585
R325 B.n478 B.n477 585
R326 B.n480 B.n219 585
R327 B.n476 B.n219 585
R328 B.n482 B.n481 585
R329 B.n483 B.n482 585
R330 B.n214 B.n213 585
R331 B.n215 B.n214 585
R332 B.n491 B.n490 585
R333 B.n490 B.n489 585
R334 B.n492 B.n212 585
R335 B.n212 B.n211 585
R336 B.n494 B.n493 585
R337 B.n495 B.n494 585
R338 B.n206 B.n205 585
R339 B.n207 B.n206 585
R340 B.n503 B.n502 585
R341 B.n502 B.n501 585
R342 B.n504 B.n204 585
R343 B.n204 B.n203 585
R344 B.n506 B.n505 585
R345 B.n507 B.n506 585
R346 B.n198 B.n197 585
R347 B.n199 B.n198 585
R348 B.n516 B.n515 585
R349 B.n515 B.n514 585
R350 B.n517 B.n196 585
R351 B.n196 B.n195 585
R352 B.n519 B.n518 585
R353 B.n520 B.n519 585
R354 B.n3 B.n0 585
R355 B.n4 B.n3 585
R356 B.n671 B.n1 585
R357 B.n672 B.n671 585
R358 B.n670 B.n669 585
R359 B.n670 B.n8 585
R360 B.n668 B.n9 585
R361 B.n12 B.n9 585
R362 B.n667 B.n666 585
R363 B.n666 B.n665 585
R364 B.n11 B.n10 585
R365 B.n664 B.n11 585
R366 B.n662 B.n661 585
R367 B.n663 B.n662 585
R368 B.n660 B.n17 585
R369 B.n17 B.n16 585
R370 B.n659 B.n658 585
R371 B.n658 B.n657 585
R372 B.n19 B.n18 585
R373 B.n656 B.n19 585
R374 B.n654 B.n653 585
R375 B.n655 B.n654 585
R376 B.n652 B.n24 585
R377 B.n24 B.n23 585
R378 B.n651 B.n650 585
R379 B.n650 B.n649 585
R380 B.n26 B.n25 585
R381 B.n648 B.n26 585
R382 B.n646 B.n645 585
R383 B.n647 B.n646 585
R384 B.n644 B.n30 585
R385 B.n33 B.n30 585
R386 B.n643 B.n642 585
R387 B.n642 B.n641 585
R388 B.n32 B.n31 585
R389 B.n640 B.n32 585
R390 B.n638 B.n637 585
R391 B.n639 B.n638 585
R392 B.n636 B.n38 585
R393 B.n38 B.n37 585
R394 B.n635 B.n634 585
R395 B.n634 B.n633 585
R396 B.n40 B.n39 585
R397 B.n632 B.n40 585
R398 B.n630 B.n629 585
R399 B.n631 B.n630 585
R400 B.n628 B.n45 585
R401 B.n45 B.n44 585
R402 B.n627 B.n626 585
R403 B.n626 B.n625 585
R404 B.n47 B.n46 585
R405 B.n624 B.n47 585
R406 B.n622 B.n621 585
R407 B.n623 B.n622 585
R408 B.n620 B.n52 585
R409 B.n52 B.n51 585
R410 B.n619 B.n618 585
R411 B.n618 B.n617 585
R412 B.n54 B.n53 585
R413 B.n616 B.n54 585
R414 B.n614 B.n613 585
R415 B.n615 B.n614 585
R416 B.n612 B.n59 585
R417 B.n59 B.n58 585
R418 B.n611 B.n610 585
R419 B.n610 B.n609 585
R420 B.n61 B.n60 585
R421 B.n608 B.n61 585
R422 B.n606 B.n605 585
R423 B.n607 B.n606 585
R424 B.n604 B.n66 585
R425 B.n66 B.n65 585
R426 B.n603 B.n602 585
R427 B.n602 B.n601 585
R428 B.n68 B.n67 585
R429 B.n600 B.n68 585
R430 B.n598 B.n597 585
R431 B.n599 B.n598 585
R432 B.n596 B.n73 585
R433 B.n73 B.n72 585
R434 B.n595 B.n594 585
R435 B.n594 B.n593 585
R436 B.n75 B.n74 585
R437 B.n592 B.n75 585
R438 B.n590 B.n589 585
R439 B.n591 B.n590 585
R440 B.n588 B.n80 585
R441 B.n80 B.n79 585
R442 B.n587 B.n586 585
R443 B.n586 B.n585 585
R444 B.n675 B.n674 585
R445 B.n673 B.n2 585
R446 B.n586 B.n82 487.695
R447 B.n583 B.n83 487.695
R448 B.n391 B.n279 487.695
R449 B.n393 B.n277 487.695
R450 B.n584 B.n104 256.663
R451 B.n584 B.n103 256.663
R452 B.n584 B.n102 256.663
R453 B.n584 B.n101 256.663
R454 B.n584 B.n100 256.663
R455 B.n584 B.n99 256.663
R456 B.n584 B.n98 256.663
R457 B.n584 B.n97 256.663
R458 B.n584 B.n96 256.663
R459 B.n584 B.n95 256.663
R460 B.n584 B.n94 256.663
R461 B.n584 B.n93 256.663
R462 B.n584 B.n92 256.663
R463 B.n584 B.n91 256.663
R464 B.n584 B.n90 256.663
R465 B.n584 B.n89 256.663
R466 B.n584 B.n88 256.663
R467 B.n584 B.n87 256.663
R468 B.n584 B.n86 256.663
R469 B.n584 B.n85 256.663
R470 B.n584 B.n84 256.663
R471 B.n305 B.n278 256.663
R472 B.n311 B.n278 256.663
R473 B.n313 B.n278 256.663
R474 B.n319 B.n278 256.663
R475 B.n321 B.n278 256.663
R476 B.n327 B.n278 256.663
R477 B.n329 B.n278 256.663
R478 B.n335 B.n278 256.663
R479 B.n337 B.n278 256.663
R480 B.n343 B.n278 256.663
R481 B.n345 B.n278 256.663
R482 B.n351 B.n278 256.663
R483 B.n353 B.n278 256.663
R484 B.n360 B.n278 256.663
R485 B.n362 B.n278 256.663
R486 B.n368 B.n278 256.663
R487 B.n370 B.n278 256.663
R488 B.n376 B.n278 256.663
R489 B.n378 B.n278 256.663
R490 B.n384 B.n278 256.663
R491 B.n386 B.n278 256.663
R492 B.n677 B.n676 256.663
R493 B.n109 B.t17 238.567
R494 B.n106 B.t13 238.567
R495 B.n288 B.t6 238.567
R496 B.n294 B.t10 238.567
R497 B.n113 B.n112 163.367
R498 B.n117 B.n116 163.367
R499 B.n121 B.n120 163.367
R500 B.n125 B.n124 163.367
R501 B.n129 B.n128 163.367
R502 B.n133 B.n132 163.367
R503 B.n137 B.n136 163.367
R504 B.n141 B.n140 163.367
R505 B.n146 B.n145 163.367
R506 B.n150 B.n149 163.367
R507 B.n154 B.n153 163.367
R508 B.n158 B.n157 163.367
R509 B.n162 B.n161 163.367
R510 B.n166 B.n165 163.367
R511 B.n170 B.n169 163.367
R512 B.n174 B.n173 163.367
R513 B.n178 B.n177 163.367
R514 B.n182 B.n181 163.367
R515 B.n186 B.n185 163.367
R516 B.n190 B.n189 163.367
R517 B.n583 B.n105 163.367
R518 B.n391 B.n273 163.367
R519 B.n399 B.n273 163.367
R520 B.n399 B.n271 163.367
R521 B.n403 B.n271 163.367
R522 B.n403 B.n264 163.367
R523 B.n411 B.n264 163.367
R524 B.n411 B.n262 163.367
R525 B.n415 B.n262 163.367
R526 B.n415 B.n257 163.367
R527 B.n423 B.n257 163.367
R528 B.n423 B.n255 163.367
R529 B.n427 B.n255 163.367
R530 B.n427 B.n249 163.367
R531 B.n435 B.n249 163.367
R532 B.n435 B.n247 163.367
R533 B.n439 B.n247 163.367
R534 B.n439 B.n241 163.367
R535 B.n447 B.n241 163.367
R536 B.n447 B.n239 163.367
R537 B.n451 B.n239 163.367
R538 B.n451 B.n233 163.367
R539 B.n459 B.n233 163.367
R540 B.n459 B.n231 163.367
R541 B.n463 B.n231 163.367
R542 B.n463 B.n225 163.367
R543 B.n471 B.n225 163.367
R544 B.n471 B.n223 163.367
R545 B.n475 B.n223 163.367
R546 B.n475 B.n218 163.367
R547 B.n484 B.n218 163.367
R548 B.n484 B.n216 163.367
R549 B.n488 B.n216 163.367
R550 B.n488 B.n210 163.367
R551 B.n496 B.n210 163.367
R552 B.n496 B.n208 163.367
R553 B.n500 B.n208 163.367
R554 B.n500 B.n202 163.367
R555 B.n508 B.n202 163.367
R556 B.n508 B.n200 163.367
R557 B.n513 B.n200 163.367
R558 B.n513 B.n194 163.367
R559 B.n521 B.n194 163.367
R560 B.n522 B.n521 163.367
R561 B.n522 B.n5 163.367
R562 B.n6 B.n5 163.367
R563 B.n7 B.n6 163.367
R564 B.n528 B.n7 163.367
R565 B.n529 B.n528 163.367
R566 B.n529 B.n13 163.367
R567 B.n14 B.n13 163.367
R568 B.n15 B.n14 163.367
R569 B.n534 B.n15 163.367
R570 B.n534 B.n20 163.367
R571 B.n21 B.n20 163.367
R572 B.n22 B.n21 163.367
R573 B.n539 B.n22 163.367
R574 B.n539 B.n27 163.367
R575 B.n28 B.n27 163.367
R576 B.n29 B.n28 163.367
R577 B.n544 B.n29 163.367
R578 B.n544 B.n34 163.367
R579 B.n35 B.n34 163.367
R580 B.n36 B.n35 163.367
R581 B.n549 B.n36 163.367
R582 B.n549 B.n41 163.367
R583 B.n42 B.n41 163.367
R584 B.n43 B.n42 163.367
R585 B.n554 B.n43 163.367
R586 B.n554 B.n48 163.367
R587 B.n49 B.n48 163.367
R588 B.n50 B.n49 163.367
R589 B.n559 B.n50 163.367
R590 B.n559 B.n55 163.367
R591 B.n56 B.n55 163.367
R592 B.n57 B.n56 163.367
R593 B.n564 B.n57 163.367
R594 B.n564 B.n62 163.367
R595 B.n63 B.n62 163.367
R596 B.n64 B.n63 163.367
R597 B.n569 B.n64 163.367
R598 B.n569 B.n69 163.367
R599 B.n70 B.n69 163.367
R600 B.n71 B.n70 163.367
R601 B.n574 B.n71 163.367
R602 B.n574 B.n76 163.367
R603 B.n77 B.n76 163.367
R604 B.n78 B.n77 163.367
R605 B.n579 B.n78 163.367
R606 B.n579 B.n83 163.367
R607 B.n306 B.n304 163.367
R608 B.n310 B.n304 163.367
R609 B.n314 B.n312 163.367
R610 B.n318 B.n302 163.367
R611 B.n322 B.n320 163.367
R612 B.n326 B.n300 163.367
R613 B.n330 B.n328 163.367
R614 B.n334 B.n298 163.367
R615 B.n338 B.n336 163.367
R616 B.n342 B.n293 163.367
R617 B.n346 B.n344 163.367
R618 B.n350 B.n291 163.367
R619 B.n354 B.n352 163.367
R620 B.n359 B.n287 163.367
R621 B.n363 B.n361 163.367
R622 B.n367 B.n285 163.367
R623 B.n371 B.n369 163.367
R624 B.n375 B.n283 163.367
R625 B.n379 B.n377 163.367
R626 B.n383 B.n281 163.367
R627 B.n387 B.n385 163.367
R628 B.n393 B.n275 163.367
R629 B.n397 B.n275 163.367
R630 B.n397 B.n269 163.367
R631 B.n405 B.n269 163.367
R632 B.n405 B.n267 163.367
R633 B.n409 B.n267 163.367
R634 B.n409 B.n261 163.367
R635 B.n417 B.n261 163.367
R636 B.n417 B.n259 163.367
R637 B.n421 B.n259 163.367
R638 B.n421 B.n253 163.367
R639 B.n429 B.n253 163.367
R640 B.n429 B.n251 163.367
R641 B.n433 B.n251 163.367
R642 B.n433 B.n245 163.367
R643 B.n441 B.n245 163.367
R644 B.n441 B.n243 163.367
R645 B.n445 B.n243 163.367
R646 B.n445 B.n237 163.367
R647 B.n453 B.n237 163.367
R648 B.n453 B.n235 163.367
R649 B.n457 B.n235 163.367
R650 B.n457 B.n229 163.367
R651 B.n465 B.n229 163.367
R652 B.n465 B.n227 163.367
R653 B.n469 B.n227 163.367
R654 B.n469 B.n221 163.367
R655 B.n478 B.n221 163.367
R656 B.n478 B.n219 163.367
R657 B.n482 B.n219 163.367
R658 B.n482 B.n214 163.367
R659 B.n490 B.n214 163.367
R660 B.n490 B.n212 163.367
R661 B.n494 B.n212 163.367
R662 B.n494 B.n206 163.367
R663 B.n502 B.n206 163.367
R664 B.n502 B.n204 163.367
R665 B.n506 B.n204 163.367
R666 B.n506 B.n198 163.367
R667 B.n515 B.n198 163.367
R668 B.n515 B.n196 163.367
R669 B.n519 B.n196 163.367
R670 B.n519 B.n3 163.367
R671 B.n675 B.n3 163.367
R672 B.n671 B.n2 163.367
R673 B.n671 B.n670 163.367
R674 B.n670 B.n9 163.367
R675 B.n666 B.n9 163.367
R676 B.n666 B.n11 163.367
R677 B.n662 B.n11 163.367
R678 B.n662 B.n17 163.367
R679 B.n658 B.n17 163.367
R680 B.n658 B.n19 163.367
R681 B.n654 B.n19 163.367
R682 B.n654 B.n24 163.367
R683 B.n650 B.n24 163.367
R684 B.n650 B.n26 163.367
R685 B.n646 B.n26 163.367
R686 B.n646 B.n30 163.367
R687 B.n642 B.n30 163.367
R688 B.n642 B.n32 163.367
R689 B.n638 B.n32 163.367
R690 B.n638 B.n38 163.367
R691 B.n634 B.n38 163.367
R692 B.n634 B.n40 163.367
R693 B.n630 B.n40 163.367
R694 B.n630 B.n45 163.367
R695 B.n626 B.n45 163.367
R696 B.n626 B.n47 163.367
R697 B.n622 B.n47 163.367
R698 B.n622 B.n52 163.367
R699 B.n618 B.n52 163.367
R700 B.n618 B.n54 163.367
R701 B.n614 B.n54 163.367
R702 B.n614 B.n59 163.367
R703 B.n610 B.n59 163.367
R704 B.n610 B.n61 163.367
R705 B.n606 B.n61 163.367
R706 B.n606 B.n66 163.367
R707 B.n602 B.n66 163.367
R708 B.n602 B.n68 163.367
R709 B.n598 B.n68 163.367
R710 B.n598 B.n73 163.367
R711 B.n594 B.n73 163.367
R712 B.n594 B.n75 163.367
R713 B.n590 B.n75 163.367
R714 B.n590 B.n80 163.367
R715 B.n586 B.n80 163.367
R716 B.n392 B.n278 162.079
R717 B.n585 B.n584 162.079
R718 B.n106 B.t15 134.323
R719 B.n288 B.t9 134.323
R720 B.n109 B.t18 134.321
R721 B.n294 B.t12 134.321
R722 B.n392 B.n274 85.4374
R723 B.n398 B.n274 85.4374
R724 B.n398 B.n270 85.4374
R725 B.n404 B.n270 85.4374
R726 B.n404 B.n265 85.4374
R727 B.n410 B.n265 85.4374
R728 B.n410 B.n266 85.4374
R729 B.n416 B.n258 85.4374
R730 B.n422 B.n258 85.4374
R731 B.n422 B.n254 85.4374
R732 B.n428 B.n254 85.4374
R733 B.n428 B.n250 85.4374
R734 B.n434 B.n250 85.4374
R735 B.n434 B.n246 85.4374
R736 B.n440 B.n246 85.4374
R737 B.n440 B.n242 85.4374
R738 B.n446 B.n242 85.4374
R739 B.n446 B.n238 85.4374
R740 B.n452 B.n238 85.4374
R741 B.n458 B.n234 85.4374
R742 B.n458 B.n230 85.4374
R743 B.n464 B.n230 85.4374
R744 B.n464 B.n226 85.4374
R745 B.n470 B.n226 85.4374
R746 B.n470 B.n222 85.4374
R747 B.n477 B.n222 85.4374
R748 B.n477 B.n476 85.4374
R749 B.n483 B.n215 85.4374
R750 B.n489 B.n215 85.4374
R751 B.n489 B.n211 85.4374
R752 B.n495 B.n211 85.4374
R753 B.n495 B.n207 85.4374
R754 B.n501 B.n207 85.4374
R755 B.n501 B.n203 85.4374
R756 B.n507 B.n203 85.4374
R757 B.n514 B.n199 85.4374
R758 B.n514 B.n195 85.4374
R759 B.n520 B.n195 85.4374
R760 B.n520 B.n4 85.4374
R761 B.n674 B.n4 85.4374
R762 B.n674 B.n673 85.4374
R763 B.n673 B.n672 85.4374
R764 B.n672 B.n8 85.4374
R765 B.n12 B.n8 85.4374
R766 B.n665 B.n12 85.4374
R767 B.n665 B.n664 85.4374
R768 B.n663 B.n16 85.4374
R769 B.n657 B.n16 85.4374
R770 B.n657 B.n656 85.4374
R771 B.n656 B.n655 85.4374
R772 B.n655 B.n23 85.4374
R773 B.n649 B.n23 85.4374
R774 B.n649 B.n648 85.4374
R775 B.n648 B.n647 85.4374
R776 B.n641 B.n33 85.4374
R777 B.n641 B.n640 85.4374
R778 B.n640 B.n639 85.4374
R779 B.n639 B.n37 85.4374
R780 B.n633 B.n37 85.4374
R781 B.n633 B.n632 85.4374
R782 B.n632 B.n631 85.4374
R783 B.n631 B.n44 85.4374
R784 B.n625 B.n624 85.4374
R785 B.n624 B.n623 85.4374
R786 B.n623 B.n51 85.4374
R787 B.n617 B.n51 85.4374
R788 B.n617 B.n616 85.4374
R789 B.n616 B.n615 85.4374
R790 B.n615 B.n58 85.4374
R791 B.n609 B.n58 85.4374
R792 B.n609 B.n608 85.4374
R793 B.n608 B.n607 85.4374
R794 B.n607 B.n65 85.4374
R795 B.n601 B.n65 85.4374
R796 B.n600 B.n599 85.4374
R797 B.n599 B.n72 85.4374
R798 B.n593 B.n72 85.4374
R799 B.n593 B.n592 85.4374
R800 B.n592 B.n591 85.4374
R801 B.n591 B.n79 85.4374
R802 B.n585 B.n79 85.4374
R803 B.t3 B.n234 76.6424
R804 B.t0 B.n44 76.6424
R805 B.n107 B.t16 74.2027
R806 B.n289 B.t8 74.2027
R807 B.n110 B.t19 74.1998
R808 B.n295 B.t11 74.1998
R809 B.n84 B.n82 71.676
R810 B.n113 B.n85 71.676
R811 B.n117 B.n86 71.676
R812 B.n121 B.n87 71.676
R813 B.n125 B.n88 71.676
R814 B.n129 B.n89 71.676
R815 B.n133 B.n90 71.676
R816 B.n137 B.n91 71.676
R817 B.n141 B.n92 71.676
R818 B.n146 B.n93 71.676
R819 B.n150 B.n94 71.676
R820 B.n154 B.n95 71.676
R821 B.n158 B.n96 71.676
R822 B.n162 B.n97 71.676
R823 B.n166 B.n98 71.676
R824 B.n170 B.n99 71.676
R825 B.n174 B.n100 71.676
R826 B.n178 B.n101 71.676
R827 B.n182 B.n102 71.676
R828 B.n186 B.n103 71.676
R829 B.n190 B.n104 71.676
R830 B.n105 B.n104 71.676
R831 B.n189 B.n103 71.676
R832 B.n185 B.n102 71.676
R833 B.n181 B.n101 71.676
R834 B.n177 B.n100 71.676
R835 B.n173 B.n99 71.676
R836 B.n169 B.n98 71.676
R837 B.n165 B.n97 71.676
R838 B.n161 B.n96 71.676
R839 B.n157 B.n95 71.676
R840 B.n153 B.n94 71.676
R841 B.n149 B.n93 71.676
R842 B.n145 B.n92 71.676
R843 B.n140 B.n91 71.676
R844 B.n136 B.n90 71.676
R845 B.n132 B.n89 71.676
R846 B.n128 B.n88 71.676
R847 B.n124 B.n87 71.676
R848 B.n120 B.n86 71.676
R849 B.n116 B.n85 71.676
R850 B.n112 B.n84 71.676
R851 B.n305 B.n277 71.676
R852 B.n311 B.n310 71.676
R853 B.n314 B.n313 71.676
R854 B.n319 B.n318 71.676
R855 B.n322 B.n321 71.676
R856 B.n327 B.n326 71.676
R857 B.n330 B.n329 71.676
R858 B.n335 B.n334 71.676
R859 B.n338 B.n337 71.676
R860 B.n343 B.n342 71.676
R861 B.n346 B.n345 71.676
R862 B.n351 B.n350 71.676
R863 B.n354 B.n353 71.676
R864 B.n360 B.n359 71.676
R865 B.n363 B.n362 71.676
R866 B.n368 B.n367 71.676
R867 B.n371 B.n370 71.676
R868 B.n376 B.n375 71.676
R869 B.n379 B.n378 71.676
R870 B.n384 B.n383 71.676
R871 B.n387 B.n386 71.676
R872 B.n306 B.n305 71.676
R873 B.n312 B.n311 71.676
R874 B.n313 B.n302 71.676
R875 B.n320 B.n319 71.676
R876 B.n321 B.n300 71.676
R877 B.n328 B.n327 71.676
R878 B.n329 B.n298 71.676
R879 B.n336 B.n335 71.676
R880 B.n337 B.n293 71.676
R881 B.n344 B.n343 71.676
R882 B.n345 B.n291 71.676
R883 B.n352 B.n351 71.676
R884 B.n353 B.n287 71.676
R885 B.n361 B.n360 71.676
R886 B.n362 B.n285 71.676
R887 B.n369 B.n368 71.676
R888 B.n370 B.n283 71.676
R889 B.n377 B.n376 71.676
R890 B.n378 B.n281 71.676
R891 B.n385 B.n384 71.676
R892 B.n386 B.n279 71.676
R893 B.n676 B.n675 71.676
R894 B.n676 B.n2 71.676
R895 B.n266 B.t7 66.591
R896 B.n483 B.t5 66.591
R897 B.n647 B.t1 66.591
R898 B.t14 B.n600 66.591
R899 B.n110 B.n109 60.1217
R900 B.n107 B.n106 60.1217
R901 B.n289 B.n288 60.1217
R902 B.n295 B.n294 60.1217
R903 B.n143 B.n110 59.5399
R904 B.n108 B.n107 59.5399
R905 B.n356 B.n289 59.5399
R906 B.n296 B.n295 59.5399
R907 B.t2 B.n199 56.5396
R908 B.n664 B.t4 56.5396
R909 B.n394 B.n276 31.6883
R910 B.n390 B.n389 31.6883
R911 B.n582 B.n581 31.6883
R912 B.n587 B.n81 31.6883
R913 B.n507 B.t2 28.8983
R914 B.t4 B.n663 28.8983
R915 B.n416 B.t7 18.8469
R916 B.n476 B.t5 18.8469
R917 B.n33 B.t1 18.8469
R918 B.n601 B.t14 18.8469
R919 B B.n677 18.0485
R920 B.n395 B.n394 10.6151
R921 B.n396 B.n395 10.6151
R922 B.n396 B.n268 10.6151
R923 B.n406 B.n268 10.6151
R924 B.n407 B.n406 10.6151
R925 B.n408 B.n407 10.6151
R926 B.n408 B.n260 10.6151
R927 B.n418 B.n260 10.6151
R928 B.n419 B.n418 10.6151
R929 B.n420 B.n419 10.6151
R930 B.n420 B.n252 10.6151
R931 B.n430 B.n252 10.6151
R932 B.n431 B.n430 10.6151
R933 B.n432 B.n431 10.6151
R934 B.n432 B.n244 10.6151
R935 B.n442 B.n244 10.6151
R936 B.n443 B.n442 10.6151
R937 B.n444 B.n443 10.6151
R938 B.n444 B.n236 10.6151
R939 B.n454 B.n236 10.6151
R940 B.n455 B.n454 10.6151
R941 B.n456 B.n455 10.6151
R942 B.n456 B.n228 10.6151
R943 B.n466 B.n228 10.6151
R944 B.n467 B.n466 10.6151
R945 B.n468 B.n467 10.6151
R946 B.n468 B.n220 10.6151
R947 B.n479 B.n220 10.6151
R948 B.n480 B.n479 10.6151
R949 B.n481 B.n480 10.6151
R950 B.n481 B.n213 10.6151
R951 B.n491 B.n213 10.6151
R952 B.n492 B.n491 10.6151
R953 B.n493 B.n492 10.6151
R954 B.n493 B.n205 10.6151
R955 B.n503 B.n205 10.6151
R956 B.n504 B.n503 10.6151
R957 B.n505 B.n504 10.6151
R958 B.n505 B.n197 10.6151
R959 B.n516 B.n197 10.6151
R960 B.n517 B.n516 10.6151
R961 B.n518 B.n517 10.6151
R962 B.n518 B.n0 10.6151
R963 B.n307 B.n276 10.6151
R964 B.n308 B.n307 10.6151
R965 B.n309 B.n308 10.6151
R966 B.n309 B.n303 10.6151
R967 B.n315 B.n303 10.6151
R968 B.n316 B.n315 10.6151
R969 B.n317 B.n316 10.6151
R970 B.n317 B.n301 10.6151
R971 B.n323 B.n301 10.6151
R972 B.n324 B.n323 10.6151
R973 B.n325 B.n324 10.6151
R974 B.n325 B.n299 10.6151
R975 B.n331 B.n299 10.6151
R976 B.n332 B.n331 10.6151
R977 B.n333 B.n332 10.6151
R978 B.n333 B.n297 10.6151
R979 B.n340 B.n339 10.6151
R980 B.n341 B.n340 10.6151
R981 B.n341 B.n292 10.6151
R982 B.n347 B.n292 10.6151
R983 B.n348 B.n347 10.6151
R984 B.n349 B.n348 10.6151
R985 B.n349 B.n290 10.6151
R986 B.n355 B.n290 10.6151
R987 B.n358 B.n357 10.6151
R988 B.n358 B.n286 10.6151
R989 B.n364 B.n286 10.6151
R990 B.n365 B.n364 10.6151
R991 B.n366 B.n365 10.6151
R992 B.n366 B.n284 10.6151
R993 B.n372 B.n284 10.6151
R994 B.n373 B.n372 10.6151
R995 B.n374 B.n373 10.6151
R996 B.n374 B.n282 10.6151
R997 B.n380 B.n282 10.6151
R998 B.n381 B.n380 10.6151
R999 B.n382 B.n381 10.6151
R1000 B.n382 B.n280 10.6151
R1001 B.n388 B.n280 10.6151
R1002 B.n389 B.n388 10.6151
R1003 B.n390 B.n272 10.6151
R1004 B.n400 B.n272 10.6151
R1005 B.n401 B.n400 10.6151
R1006 B.n402 B.n401 10.6151
R1007 B.n402 B.n263 10.6151
R1008 B.n412 B.n263 10.6151
R1009 B.n413 B.n412 10.6151
R1010 B.n414 B.n413 10.6151
R1011 B.n414 B.n256 10.6151
R1012 B.n424 B.n256 10.6151
R1013 B.n425 B.n424 10.6151
R1014 B.n426 B.n425 10.6151
R1015 B.n426 B.n248 10.6151
R1016 B.n436 B.n248 10.6151
R1017 B.n437 B.n436 10.6151
R1018 B.n438 B.n437 10.6151
R1019 B.n438 B.n240 10.6151
R1020 B.n448 B.n240 10.6151
R1021 B.n449 B.n448 10.6151
R1022 B.n450 B.n449 10.6151
R1023 B.n450 B.n232 10.6151
R1024 B.n460 B.n232 10.6151
R1025 B.n461 B.n460 10.6151
R1026 B.n462 B.n461 10.6151
R1027 B.n462 B.n224 10.6151
R1028 B.n472 B.n224 10.6151
R1029 B.n473 B.n472 10.6151
R1030 B.n474 B.n473 10.6151
R1031 B.n474 B.n217 10.6151
R1032 B.n485 B.n217 10.6151
R1033 B.n486 B.n485 10.6151
R1034 B.n487 B.n486 10.6151
R1035 B.n487 B.n209 10.6151
R1036 B.n497 B.n209 10.6151
R1037 B.n498 B.n497 10.6151
R1038 B.n499 B.n498 10.6151
R1039 B.n499 B.n201 10.6151
R1040 B.n509 B.n201 10.6151
R1041 B.n510 B.n509 10.6151
R1042 B.n512 B.n510 10.6151
R1043 B.n512 B.n511 10.6151
R1044 B.n511 B.n193 10.6151
R1045 B.n523 B.n193 10.6151
R1046 B.n524 B.n523 10.6151
R1047 B.n525 B.n524 10.6151
R1048 B.n526 B.n525 10.6151
R1049 B.n527 B.n526 10.6151
R1050 B.n530 B.n527 10.6151
R1051 B.n531 B.n530 10.6151
R1052 B.n532 B.n531 10.6151
R1053 B.n533 B.n532 10.6151
R1054 B.n535 B.n533 10.6151
R1055 B.n536 B.n535 10.6151
R1056 B.n537 B.n536 10.6151
R1057 B.n538 B.n537 10.6151
R1058 B.n540 B.n538 10.6151
R1059 B.n541 B.n540 10.6151
R1060 B.n542 B.n541 10.6151
R1061 B.n543 B.n542 10.6151
R1062 B.n545 B.n543 10.6151
R1063 B.n546 B.n545 10.6151
R1064 B.n547 B.n546 10.6151
R1065 B.n548 B.n547 10.6151
R1066 B.n550 B.n548 10.6151
R1067 B.n551 B.n550 10.6151
R1068 B.n552 B.n551 10.6151
R1069 B.n553 B.n552 10.6151
R1070 B.n555 B.n553 10.6151
R1071 B.n556 B.n555 10.6151
R1072 B.n557 B.n556 10.6151
R1073 B.n558 B.n557 10.6151
R1074 B.n560 B.n558 10.6151
R1075 B.n561 B.n560 10.6151
R1076 B.n562 B.n561 10.6151
R1077 B.n563 B.n562 10.6151
R1078 B.n565 B.n563 10.6151
R1079 B.n566 B.n565 10.6151
R1080 B.n567 B.n566 10.6151
R1081 B.n568 B.n567 10.6151
R1082 B.n570 B.n568 10.6151
R1083 B.n571 B.n570 10.6151
R1084 B.n572 B.n571 10.6151
R1085 B.n573 B.n572 10.6151
R1086 B.n575 B.n573 10.6151
R1087 B.n576 B.n575 10.6151
R1088 B.n577 B.n576 10.6151
R1089 B.n578 B.n577 10.6151
R1090 B.n580 B.n578 10.6151
R1091 B.n581 B.n580 10.6151
R1092 B.n669 B.n1 10.6151
R1093 B.n669 B.n668 10.6151
R1094 B.n668 B.n667 10.6151
R1095 B.n667 B.n10 10.6151
R1096 B.n661 B.n10 10.6151
R1097 B.n661 B.n660 10.6151
R1098 B.n660 B.n659 10.6151
R1099 B.n659 B.n18 10.6151
R1100 B.n653 B.n18 10.6151
R1101 B.n653 B.n652 10.6151
R1102 B.n652 B.n651 10.6151
R1103 B.n651 B.n25 10.6151
R1104 B.n645 B.n25 10.6151
R1105 B.n645 B.n644 10.6151
R1106 B.n644 B.n643 10.6151
R1107 B.n643 B.n31 10.6151
R1108 B.n637 B.n31 10.6151
R1109 B.n637 B.n636 10.6151
R1110 B.n636 B.n635 10.6151
R1111 B.n635 B.n39 10.6151
R1112 B.n629 B.n39 10.6151
R1113 B.n629 B.n628 10.6151
R1114 B.n628 B.n627 10.6151
R1115 B.n627 B.n46 10.6151
R1116 B.n621 B.n46 10.6151
R1117 B.n621 B.n620 10.6151
R1118 B.n620 B.n619 10.6151
R1119 B.n619 B.n53 10.6151
R1120 B.n613 B.n53 10.6151
R1121 B.n613 B.n612 10.6151
R1122 B.n612 B.n611 10.6151
R1123 B.n611 B.n60 10.6151
R1124 B.n605 B.n60 10.6151
R1125 B.n605 B.n604 10.6151
R1126 B.n604 B.n603 10.6151
R1127 B.n603 B.n67 10.6151
R1128 B.n597 B.n67 10.6151
R1129 B.n597 B.n596 10.6151
R1130 B.n596 B.n595 10.6151
R1131 B.n595 B.n74 10.6151
R1132 B.n589 B.n74 10.6151
R1133 B.n589 B.n588 10.6151
R1134 B.n588 B.n587 10.6151
R1135 B.n111 B.n81 10.6151
R1136 B.n114 B.n111 10.6151
R1137 B.n115 B.n114 10.6151
R1138 B.n118 B.n115 10.6151
R1139 B.n119 B.n118 10.6151
R1140 B.n122 B.n119 10.6151
R1141 B.n123 B.n122 10.6151
R1142 B.n126 B.n123 10.6151
R1143 B.n127 B.n126 10.6151
R1144 B.n130 B.n127 10.6151
R1145 B.n131 B.n130 10.6151
R1146 B.n134 B.n131 10.6151
R1147 B.n135 B.n134 10.6151
R1148 B.n138 B.n135 10.6151
R1149 B.n139 B.n138 10.6151
R1150 B.n142 B.n139 10.6151
R1151 B.n147 B.n144 10.6151
R1152 B.n148 B.n147 10.6151
R1153 B.n151 B.n148 10.6151
R1154 B.n152 B.n151 10.6151
R1155 B.n155 B.n152 10.6151
R1156 B.n156 B.n155 10.6151
R1157 B.n159 B.n156 10.6151
R1158 B.n160 B.n159 10.6151
R1159 B.n164 B.n163 10.6151
R1160 B.n167 B.n164 10.6151
R1161 B.n168 B.n167 10.6151
R1162 B.n171 B.n168 10.6151
R1163 B.n172 B.n171 10.6151
R1164 B.n175 B.n172 10.6151
R1165 B.n176 B.n175 10.6151
R1166 B.n179 B.n176 10.6151
R1167 B.n180 B.n179 10.6151
R1168 B.n183 B.n180 10.6151
R1169 B.n184 B.n183 10.6151
R1170 B.n187 B.n184 10.6151
R1171 B.n188 B.n187 10.6151
R1172 B.n191 B.n188 10.6151
R1173 B.n192 B.n191 10.6151
R1174 B.n582 B.n192 10.6151
R1175 B.n452 B.t3 8.79547
R1176 B.n625 B.t0 8.79547
R1177 B.n677 B.n0 8.11757
R1178 B.n677 B.n1 8.11757
R1179 B.n339 B.n296 6.5566
R1180 B.n356 B.n355 6.5566
R1181 B.n144 B.n143 6.5566
R1182 B.n160 B.n108 6.5566
R1183 B.n297 B.n296 4.05904
R1184 B.n357 B.n356 4.05904
R1185 B.n143 B.n142 4.05904
R1186 B.n163 B.n108 4.05904
R1187 VP.n13 VP.n12 161.3
R1188 VP.n14 VP.n9 161.3
R1189 VP.n16 VP.n15 161.3
R1190 VP.n17 VP.n8 161.3
R1191 VP.n19 VP.n18 161.3
R1192 VP.n20 VP.n7 161.3
R1193 VP.n43 VP.n0 161.3
R1194 VP.n42 VP.n41 161.3
R1195 VP.n40 VP.n1 161.3
R1196 VP.n39 VP.n38 161.3
R1197 VP.n37 VP.n2 161.3
R1198 VP.n36 VP.n35 161.3
R1199 VP.n34 VP.n3 161.3
R1200 VP.n33 VP.n32 161.3
R1201 VP.n31 VP.n4 161.3
R1202 VP.n30 VP.n29 161.3
R1203 VP.n28 VP.n5 161.3
R1204 VP.n27 VP.n26 161.3
R1205 VP.n25 VP.n6 161.3
R1206 VP.n24 VP.n23 105.99
R1207 VP.n45 VP.n44 105.99
R1208 VP.n22 VP.n21 105.99
R1209 VP.n11 VP.t2 64.3576
R1210 VP.n11 VP.n10 49.0286
R1211 VP.n30 VP.n5 45.4209
R1212 VP.n38 VP.n1 45.4209
R1213 VP.n15 VP.n8 45.4209
R1214 VP.n23 VP.n22 42.8709
R1215 VP.n31 VP.n30 35.7332
R1216 VP.n38 VP.n37 35.7332
R1217 VP.n15 VP.n14 35.7332
R1218 VP.n3 VP.t4 30.2778
R1219 VP.n24 VP.t3 30.2778
R1220 VP.n44 VP.t5 30.2778
R1221 VP.n10 VP.t1 30.2778
R1222 VP.n21 VP.t0 30.2778
R1223 VP.n26 VP.n25 24.5923
R1224 VP.n26 VP.n5 24.5923
R1225 VP.n32 VP.n31 24.5923
R1226 VP.n32 VP.n3 24.5923
R1227 VP.n36 VP.n3 24.5923
R1228 VP.n37 VP.n36 24.5923
R1229 VP.n42 VP.n1 24.5923
R1230 VP.n43 VP.n42 24.5923
R1231 VP.n19 VP.n8 24.5923
R1232 VP.n20 VP.n19 24.5923
R1233 VP.n13 VP.n10 24.5923
R1234 VP.n14 VP.n13 24.5923
R1235 VP.n12 VP.n11 4.96469
R1236 VP.n25 VP.n24 4.91887
R1237 VP.n44 VP.n43 4.91887
R1238 VP.n21 VP.n20 4.91887
R1239 VP.n22 VP.n7 0.278335
R1240 VP.n23 VP.n6 0.278335
R1241 VP.n45 VP.n0 0.278335
R1242 VP.n12 VP.n9 0.189894
R1243 VP.n16 VP.n9 0.189894
R1244 VP.n17 VP.n16 0.189894
R1245 VP.n18 VP.n17 0.189894
R1246 VP.n18 VP.n7 0.189894
R1247 VP.n27 VP.n6 0.189894
R1248 VP.n28 VP.n27 0.189894
R1249 VP.n29 VP.n28 0.189894
R1250 VP.n29 VP.n4 0.189894
R1251 VP.n33 VP.n4 0.189894
R1252 VP.n34 VP.n33 0.189894
R1253 VP.n35 VP.n34 0.189894
R1254 VP.n35 VP.n2 0.189894
R1255 VP.n39 VP.n2 0.189894
R1256 VP.n40 VP.n39 0.189894
R1257 VP.n41 VP.n40 0.189894
R1258 VP.n41 VP.n0 0.189894
R1259 VP VP.n45 0.153485
R1260 VTAIL.n7 VTAIL.t2 64.3714
R1261 VTAIL.n11 VTAIL.t0 64.3714
R1262 VTAIL.n2 VTAIL.t10 64.3714
R1263 VTAIL.n10 VTAIL.t11 64.3714
R1264 VTAIL.n9 VTAIL.n8 58.6819
R1265 VTAIL.n6 VTAIL.n5 58.6819
R1266 VTAIL.n1 VTAIL.n0 58.6816
R1267 VTAIL.n4 VTAIL.n3 58.6816
R1268 VTAIL.n6 VTAIL.n4 20.7117
R1269 VTAIL.n11 VTAIL.n10 18.0393
R1270 VTAIL.n0 VTAIL.t4 5.69016
R1271 VTAIL.n0 VTAIL.t1 5.69016
R1272 VTAIL.n3 VTAIL.t7 5.69016
R1273 VTAIL.n3 VTAIL.t9 5.69016
R1274 VTAIL.n8 VTAIL.t6 5.69016
R1275 VTAIL.n8 VTAIL.t8 5.69016
R1276 VTAIL.n5 VTAIL.t3 5.69016
R1277 VTAIL.n5 VTAIL.t5 5.69016
R1278 VTAIL.n7 VTAIL.n6 2.67291
R1279 VTAIL.n10 VTAIL.n9 2.67291
R1280 VTAIL.n4 VTAIL.n2 2.67291
R1281 VTAIL VTAIL.n11 1.94662
R1282 VTAIL.n9 VTAIL.n7 1.80653
R1283 VTAIL.n2 VTAIL.n1 1.80653
R1284 VTAIL VTAIL.n1 0.726793
R1285 VDD1 VDD1.t3 83.1127
R1286 VDD1.n1 VDD1.t2 82.9991
R1287 VDD1.n1 VDD1.n0 75.9732
R1288 VDD1.n3 VDD1.n2 75.3605
R1289 VDD1.n3 VDD1.n1 37.3199
R1290 VDD1.n2 VDD1.t4 5.69016
R1291 VDD1.n2 VDD1.t5 5.69016
R1292 VDD1.n0 VDD1.t1 5.69016
R1293 VDD1.n0 VDD1.t0 5.69016
R1294 VDD1 VDD1.n3 0.610414
R1295 VN.n29 VN.n16 161.3
R1296 VN.n28 VN.n27 161.3
R1297 VN.n26 VN.n17 161.3
R1298 VN.n25 VN.n24 161.3
R1299 VN.n23 VN.n18 161.3
R1300 VN.n22 VN.n21 161.3
R1301 VN.n13 VN.n0 161.3
R1302 VN.n12 VN.n11 161.3
R1303 VN.n10 VN.n1 161.3
R1304 VN.n9 VN.n8 161.3
R1305 VN.n7 VN.n2 161.3
R1306 VN.n6 VN.n5 161.3
R1307 VN.n15 VN.n14 105.99
R1308 VN.n31 VN.n30 105.99
R1309 VN.n4 VN.t1 64.3576
R1310 VN.n20 VN.t5 64.3576
R1311 VN.n20 VN.n19 49.0286
R1312 VN.n4 VN.n3 49.0286
R1313 VN.n8 VN.n1 45.4209
R1314 VN.n24 VN.n17 45.4209
R1315 VN VN.n31 43.1497
R1316 VN.n8 VN.n7 35.7332
R1317 VN.n24 VN.n23 35.7332
R1318 VN.n3 VN.t4 30.2778
R1319 VN.n14 VN.t3 30.2778
R1320 VN.n19 VN.t2 30.2778
R1321 VN.n30 VN.t0 30.2778
R1322 VN.n6 VN.n3 24.5923
R1323 VN.n7 VN.n6 24.5923
R1324 VN.n12 VN.n1 24.5923
R1325 VN.n13 VN.n12 24.5923
R1326 VN.n23 VN.n22 24.5923
R1327 VN.n22 VN.n19 24.5923
R1328 VN.n29 VN.n28 24.5923
R1329 VN.n28 VN.n17 24.5923
R1330 VN.n21 VN.n20 4.96469
R1331 VN.n5 VN.n4 4.96469
R1332 VN.n14 VN.n13 4.91887
R1333 VN.n30 VN.n29 4.91887
R1334 VN.n31 VN.n16 0.278335
R1335 VN.n15 VN.n0 0.278335
R1336 VN.n27 VN.n16 0.189894
R1337 VN.n27 VN.n26 0.189894
R1338 VN.n26 VN.n25 0.189894
R1339 VN.n25 VN.n18 0.189894
R1340 VN.n21 VN.n18 0.189894
R1341 VN.n5 VN.n2 0.189894
R1342 VN.n9 VN.n2 0.189894
R1343 VN.n10 VN.n9 0.189894
R1344 VN.n11 VN.n10 0.189894
R1345 VN.n11 VN.n0 0.189894
R1346 VN VN.n15 0.153485
R1347 VDD2.n1 VDD2.t4 82.9991
R1348 VDD2.n2 VDD2.t5 81.0502
R1349 VDD2.n1 VDD2.n0 75.9732
R1350 VDD2 VDD2.n3 75.9704
R1351 VDD2.n2 VDD2.n1 35.4006
R1352 VDD2.n3 VDD2.t3 5.69016
R1353 VDD2.n3 VDD2.t0 5.69016
R1354 VDD2.n0 VDD2.t1 5.69016
R1355 VDD2.n0 VDD2.t2 5.69016
R1356 VDD2 VDD2.n2 2.063
C0 VP VDD2 0.477589f
C1 VP VN 5.51456f
C2 VN VDD2 2.25371f
C3 VP VTAIL 3.04762f
C4 VP VDD1 2.57297f
C5 VTAIL VDD2 4.80014f
C6 VTAIL VN 3.03346f
C7 VDD1 VDD2 1.47142f
C8 VDD1 VN 0.155857f
C9 VTAIL VDD1 4.74613f
C10 VDD2 B 4.596719f
C11 VDD1 B 4.913896f
C12 VTAIL B 4.135751f
C13 VN B 12.604481f
C14 VP B 11.224395f
C15 VDD2.t4 B 0.608843f
C16 VDD2.t1 B 0.061652f
C17 VDD2.t2 B 0.061652f
C18 VDD2.n0 B 0.476254f
C19 VDD2.n1 B 2.17104f
C20 VDD2.t5 B 0.600356f
C21 VDD2.n2 B 1.91403f
C22 VDD2.t3 B 0.061652f
C23 VDD2.t0 B 0.061652f
C24 VDD2.n3 B 0.47623f
C25 VN.n0 B 0.037131f
C26 VN.t3 B 0.688006f
C27 VN.n1 B 0.053886f
C28 VN.n2 B 0.028166f
C29 VN.t4 B 0.688006f
C30 VN.n3 B 0.379177f
C31 VN.t1 B 0.934671f
C32 VN.n4 B 0.348297f
C33 VN.n5 B 0.294678f
C34 VN.n6 B 0.052231f
C35 VN.n7 B 0.056572f
C36 VN.n8 B 0.023659f
C37 VN.n9 B 0.028166f
C38 VN.n10 B 0.028166f
C39 VN.n11 B 0.028166f
C40 VN.n12 B 0.052231f
C41 VN.n13 B 0.031603f
C42 VN.n14 B 0.371787f
C43 VN.n15 B 0.050931f
C44 VN.n16 B 0.037131f
C45 VN.t0 B 0.688006f
C46 VN.n17 B 0.053886f
C47 VN.n18 B 0.028166f
C48 VN.t2 B 0.688006f
C49 VN.n19 B 0.379177f
C50 VN.t5 B 0.934671f
C51 VN.n20 B 0.348297f
C52 VN.n21 B 0.294678f
C53 VN.n22 B 0.052231f
C54 VN.n23 B 0.056572f
C55 VN.n24 B 0.023659f
C56 VN.n25 B 0.028166f
C57 VN.n26 B 0.028166f
C58 VN.n27 B 0.028166f
C59 VN.n28 B 0.052231f
C60 VN.n29 B 0.031603f
C61 VN.n30 B 0.371787f
C62 VN.n31 B 1.25929f
C63 VDD1.t3 B 0.61947f
C64 VDD1.t2 B 0.618776f
C65 VDD1.t1 B 0.062658f
C66 VDD1.t0 B 0.062658f
C67 VDD1.n0 B 0.484025f
C68 VDD1.n1 B 2.31553f
C69 VDD1.t4 B 0.062658f
C70 VDD1.t5 B 0.062658f
C71 VDD1.n2 B 0.480598f
C72 VDD1.n3 B 1.96857f
C73 VTAIL.t4 B 0.083965f
C74 VTAIL.t1 B 0.083965f
C75 VTAIL.n0 B 0.579568f
C76 VTAIL.n1 B 0.504704f
C77 VTAIL.t10 B 0.744516f
C78 VTAIL.n2 B 0.760217f
C79 VTAIL.t7 B 0.083965f
C80 VTAIL.t9 B 0.083965f
C81 VTAIL.n3 B 0.579568f
C82 VTAIL.n4 B 1.75423f
C83 VTAIL.t3 B 0.083965f
C84 VTAIL.t5 B 0.083965f
C85 VTAIL.n5 B 0.57957f
C86 VTAIL.n6 B 1.75423f
C87 VTAIL.t2 B 0.744521f
C88 VTAIL.n7 B 0.760212f
C89 VTAIL.t6 B 0.083965f
C90 VTAIL.t8 B 0.083965f
C91 VTAIL.n8 B 0.57957f
C92 VTAIL.n9 B 0.696167f
C93 VTAIL.t11 B 0.744516f
C94 VTAIL.n10 B 1.55536f
C95 VTAIL.t0 B 0.744516f
C96 VTAIL.n11 B 1.4839f
C97 VP.n0 B 0.038303f
C98 VP.t5 B 0.709719f
C99 VP.n1 B 0.055587f
C100 VP.n2 B 0.029055f
C101 VP.t4 B 0.709719f
C102 VP.n3 B 0.315513f
C103 VP.n4 B 0.029055f
C104 VP.n5 B 0.055587f
C105 VP.n6 B 0.038303f
C106 VP.t3 B 0.709719f
C107 VP.n7 B 0.038303f
C108 VP.t0 B 0.709719f
C109 VP.n8 B 0.055587f
C110 VP.n9 B 0.029055f
C111 VP.t1 B 0.709719f
C112 VP.n10 B 0.391144f
C113 VP.t2 B 0.964169f
C114 VP.n11 B 0.359289f
C115 VP.n12 B 0.303978f
C116 VP.n13 B 0.053879f
C117 VP.n14 B 0.058357f
C118 VP.n15 B 0.024406f
C119 VP.n16 B 0.029055f
C120 VP.n17 B 0.029055f
C121 VP.n18 B 0.029055f
C122 VP.n19 B 0.053879f
C123 VP.n20 B 0.0326f
C124 VP.n21 B 0.38352f
C125 VP.n22 B 1.28301f
C126 VP.n23 B 1.30745f
C127 VP.n24 B 0.38352f
C128 VP.n25 B 0.0326f
C129 VP.n26 B 0.053879f
C130 VP.n27 B 0.029055f
C131 VP.n28 B 0.029055f
C132 VP.n29 B 0.029055f
C133 VP.n30 B 0.024406f
C134 VP.n31 B 0.058357f
C135 VP.n32 B 0.053879f
C136 VP.n33 B 0.029055f
C137 VP.n34 B 0.029055f
C138 VP.n35 B 0.029055f
C139 VP.n36 B 0.053879f
C140 VP.n37 B 0.058357f
C141 VP.n38 B 0.024406f
C142 VP.n39 B 0.029055f
C143 VP.n40 B 0.029055f
C144 VP.n41 B 0.029055f
C145 VP.n42 B 0.053879f
C146 VP.n43 B 0.0326f
C147 VP.n44 B 0.38352f
C148 VP.n45 B 0.052539f
.ends

