* NGSPICE file created from diff_pair_sample_0763.ext - technology: sky130A

.subckt diff_pair_sample_0763 VTAIL VN VP B VDD2 VDD1
X0 B.t11 B.t9 B.t10 w_n2420_n3730# sky130_fd_pr__pfet_01v8 ad=5.3859 pd=28.4 as=0 ps=0 w=13.81 l=1.12
X1 VTAIL.t15 VP.t0 VDD1.t7 w_n2420_n3730# sky130_fd_pr__pfet_01v8 ad=5.3859 pd=28.4 as=2.27865 ps=14.14 w=13.81 l=1.12
X2 VDD2.t7 VN.t0 VTAIL.t3 w_n2420_n3730# sky130_fd_pr__pfet_01v8 ad=2.27865 pd=14.14 as=2.27865 ps=14.14 w=13.81 l=1.12
X3 VDD1.t2 VP.t1 VTAIL.t14 w_n2420_n3730# sky130_fd_pr__pfet_01v8 ad=2.27865 pd=14.14 as=2.27865 ps=14.14 w=13.81 l=1.12
X4 VDD1.t4 VP.t2 VTAIL.t13 w_n2420_n3730# sky130_fd_pr__pfet_01v8 ad=2.27865 pd=14.14 as=2.27865 ps=14.14 w=13.81 l=1.12
X5 VTAIL.t12 VP.t3 VDD1.t3 w_n2420_n3730# sky130_fd_pr__pfet_01v8 ad=2.27865 pd=14.14 as=2.27865 ps=14.14 w=13.81 l=1.12
X6 VDD1.t1 VP.t4 VTAIL.t11 w_n2420_n3730# sky130_fd_pr__pfet_01v8 ad=2.27865 pd=14.14 as=5.3859 ps=28.4 w=13.81 l=1.12
X7 VDD2.t6 VN.t1 VTAIL.t6 w_n2420_n3730# sky130_fd_pr__pfet_01v8 ad=2.27865 pd=14.14 as=5.3859 ps=28.4 w=13.81 l=1.12
X8 B.t8 B.t6 B.t7 w_n2420_n3730# sky130_fd_pr__pfet_01v8 ad=5.3859 pd=28.4 as=0 ps=0 w=13.81 l=1.12
X9 VTAIL.t0 VN.t2 VDD2.t5 w_n2420_n3730# sky130_fd_pr__pfet_01v8 ad=5.3859 pd=28.4 as=2.27865 ps=14.14 w=13.81 l=1.12
X10 B.t5 B.t3 B.t4 w_n2420_n3730# sky130_fd_pr__pfet_01v8 ad=5.3859 pd=28.4 as=0 ps=0 w=13.81 l=1.12
X11 VTAIL.t10 VP.t5 VDD1.t5 w_n2420_n3730# sky130_fd_pr__pfet_01v8 ad=2.27865 pd=14.14 as=2.27865 ps=14.14 w=13.81 l=1.12
X12 VDD2.t4 VN.t3 VTAIL.t4 w_n2420_n3730# sky130_fd_pr__pfet_01v8 ad=2.27865 pd=14.14 as=5.3859 ps=28.4 w=13.81 l=1.12
X13 VTAIL.t2 VN.t4 VDD2.t3 w_n2420_n3730# sky130_fd_pr__pfet_01v8 ad=2.27865 pd=14.14 as=2.27865 ps=14.14 w=13.81 l=1.12
X14 VTAIL.t7 VN.t5 VDD2.t2 w_n2420_n3730# sky130_fd_pr__pfet_01v8 ad=2.27865 pd=14.14 as=2.27865 ps=14.14 w=13.81 l=1.12
X15 VDD2.t1 VN.t6 VTAIL.t5 w_n2420_n3730# sky130_fd_pr__pfet_01v8 ad=2.27865 pd=14.14 as=2.27865 ps=14.14 w=13.81 l=1.12
X16 B.t2 B.t0 B.t1 w_n2420_n3730# sky130_fd_pr__pfet_01v8 ad=5.3859 pd=28.4 as=0 ps=0 w=13.81 l=1.12
X17 VTAIL.t1 VN.t7 VDD2.t0 w_n2420_n3730# sky130_fd_pr__pfet_01v8 ad=5.3859 pd=28.4 as=2.27865 ps=14.14 w=13.81 l=1.12
X18 VDD1.t0 VP.t6 VTAIL.t9 w_n2420_n3730# sky130_fd_pr__pfet_01v8 ad=2.27865 pd=14.14 as=5.3859 ps=28.4 w=13.81 l=1.12
X19 VTAIL.t8 VP.t7 VDD1.t6 w_n2420_n3730# sky130_fd_pr__pfet_01v8 ad=5.3859 pd=28.4 as=2.27865 ps=14.14 w=13.81 l=1.12
R0 B.n370 B.n369 585
R1 B.n368 B.n103 585
R2 B.n367 B.n366 585
R3 B.n365 B.n104 585
R4 B.n364 B.n363 585
R5 B.n362 B.n105 585
R6 B.n361 B.n360 585
R7 B.n359 B.n106 585
R8 B.n358 B.n357 585
R9 B.n356 B.n107 585
R10 B.n355 B.n354 585
R11 B.n353 B.n108 585
R12 B.n352 B.n351 585
R13 B.n350 B.n109 585
R14 B.n349 B.n348 585
R15 B.n347 B.n110 585
R16 B.n346 B.n345 585
R17 B.n344 B.n111 585
R18 B.n343 B.n342 585
R19 B.n341 B.n112 585
R20 B.n340 B.n339 585
R21 B.n338 B.n113 585
R22 B.n337 B.n336 585
R23 B.n335 B.n114 585
R24 B.n334 B.n333 585
R25 B.n332 B.n115 585
R26 B.n331 B.n330 585
R27 B.n329 B.n116 585
R28 B.n328 B.n327 585
R29 B.n326 B.n117 585
R30 B.n325 B.n324 585
R31 B.n323 B.n118 585
R32 B.n322 B.n321 585
R33 B.n320 B.n119 585
R34 B.n319 B.n318 585
R35 B.n317 B.n120 585
R36 B.n316 B.n315 585
R37 B.n314 B.n121 585
R38 B.n313 B.n312 585
R39 B.n311 B.n122 585
R40 B.n310 B.n309 585
R41 B.n308 B.n123 585
R42 B.n307 B.n306 585
R43 B.n305 B.n124 585
R44 B.n304 B.n303 585
R45 B.n302 B.n125 585
R46 B.n301 B.n300 585
R47 B.n299 B.n298 585
R48 B.n297 B.n129 585
R49 B.n296 B.n295 585
R50 B.n294 B.n130 585
R51 B.n293 B.n292 585
R52 B.n291 B.n131 585
R53 B.n290 B.n289 585
R54 B.n288 B.n132 585
R55 B.n287 B.n286 585
R56 B.n284 B.n133 585
R57 B.n283 B.n282 585
R58 B.n281 B.n136 585
R59 B.n280 B.n279 585
R60 B.n278 B.n137 585
R61 B.n277 B.n276 585
R62 B.n275 B.n138 585
R63 B.n274 B.n273 585
R64 B.n272 B.n139 585
R65 B.n271 B.n270 585
R66 B.n269 B.n140 585
R67 B.n268 B.n267 585
R68 B.n266 B.n141 585
R69 B.n265 B.n264 585
R70 B.n263 B.n142 585
R71 B.n262 B.n261 585
R72 B.n260 B.n143 585
R73 B.n259 B.n258 585
R74 B.n257 B.n144 585
R75 B.n256 B.n255 585
R76 B.n254 B.n145 585
R77 B.n253 B.n252 585
R78 B.n251 B.n146 585
R79 B.n250 B.n249 585
R80 B.n248 B.n147 585
R81 B.n247 B.n246 585
R82 B.n245 B.n148 585
R83 B.n244 B.n243 585
R84 B.n242 B.n149 585
R85 B.n241 B.n240 585
R86 B.n239 B.n150 585
R87 B.n238 B.n237 585
R88 B.n236 B.n151 585
R89 B.n235 B.n234 585
R90 B.n233 B.n152 585
R91 B.n232 B.n231 585
R92 B.n230 B.n153 585
R93 B.n229 B.n228 585
R94 B.n227 B.n154 585
R95 B.n226 B.n225 585
R96 B.n224 B.n155 585
R97 B.n223 B.n222 585
R98 B.n221 B.n156 585
R99 B.n220 B.n219 585
R100 B.n218 B.n157 585
R101 B.n217 B.n216 585
R102 B.n215 B.n158 585
R103 B.n371 B.n102 585
R104 B.n373 B.n372 585
R105 B.n374 B.n101 585
R106 B.n376 B.n375 585
R107 B.n377 B.n100 585
R108 B.n379 B.n378 585
R109 B.n380 B.n99 585
R110 B.n382 B.n381 585
R111 B.n383 B.n98 585
R112 B.n385 B.n384 585
R113 B.n386 B.n97 585
R114 B.n388 B.n387 585
R115 B.n389 B.n96 585
R116 B.n391 B.n390 585
R117 B.n392 B.n95 585
R118 B.n394 B.n393 585
R119 B.n395 B.n94 585
R120 B.n397 B.n396 585
R121 B.n398 B.n93 585
R122 B.n400 B.n399 585
R123 B.n401 B.n92 585
R124 B.n403 B.n402 585
R125 B.n404 B.n91 585
R126 B.n406 B.n405 585
R127 B.n407 B.n90 585
R128 B.n409 B.n408 585
R129 B.n410 B.n89 585
R130 B.n412 B.n411 585
R131 B.n413 B.n88 585
R132 B.n415 B.n414 585
R133 B.n416 B.n87 585
R134 B.n418 B.n417 585
R135 B.n419 B.n86 585
R136 B.n421 B.n420 585
R137 B.n422 B.n85 585
R138 B.n424 B.n423 585
R139 B.n425 B.n84 585
R140 B.n427 B.n426 585
R141 B.n428 B.n83 585
R142 B.n430 B.n429 585
R143 B.n431 B.n82 585
R144 B.n433 B.n432 585
R145 B.n434 B.n81 585
R146 B.n436 B.n435 585
R147 B.n437 B.n80 585
R148 B.n439 B.n438 585
R149 B.n440 B.n79 585
R150 B.n442 B.n441 585
R151 B.n443 B.n78 585
R152 B.n445 B.n444 585
R153 B.n446 B.n77 585
R154 B.n448 B.n447 585
R155 B.n449 B.n76 585
R156 B.n451 B.n450 585
R157 B.n452 B.n75 585
R158 B.n454 B.n453 585
R159 B.n455 B.n74 585
R160 B.n457 B.n456 585
R161 B.n458 B.n73 585
R162 B.n460 B.n459 585
R163 B.n616 B.n615 585
R164 B.n614 B.n17 585
R165 B.n613 B.n612 585
R166 B.n611 B.n18 585
R167 B.n610 B.n609 585
R168 B.n608 B.n19 585
R169 B.n607 B.n606 585
R170 B.n605 B.n20 585
R171 B.n604 B.n603 585
R172 B.n602 B.n21 585
R173 B.n601 B.n600 585
R174 B.n599 B.n22 585
R175 B.n598 B.n597 585
R176 B.n596 B.n23 585
R177 B.n595 B.n594 585
R178 B.n593 B.n24 585
R179 B.n592 B.n591 585
R180 B.n590 B.n25 585
R181 B.n589 B.n588 585
R182 B.n587 B.n26 585
R183 B.n586 B.n585 585
R184 B.n584 B.n27 585
R185 B.n583 B.n582 585
R186 B.n581 B.n28 585
R187 B.n580 B.n579 585
R188 B.n578 B.n29 585
R189 B.n577 B.n576 585
R190 B.n575 B.n30 585
R191 B.n574 B.n573 585
R192 B.n572 B.n31 585
R193 B.n571 B.n570 585
R194 B.n569 B.n32 585
R195 B.n568 B.n567 585
R196 B.n566 B.n33 585
R197 B.n565 B.n564 585
R198 B.n563 B.n34 585
R199 B.n562 B.n561 585
R200 B.n560 B.n35 585
R201 B.n559 B.n558 585
R202 B.n557 B.n36 585
R203 B.n556 B.n555 585
R204 B.n554 B.n37 585
R205 B.n553 B.n552 585
R206 B.n551 B.n38 585
R207 B.n550 B.n549 585
R208 B.n548 B.n39 585
R209 B.n547 B.n546 585
R210 B.n545 B.n544 585
R211 B.n543 B.n43 585
R212 B.n542 B.n541 585
R213 B.n540 B.n44 585
R214 B.n539 B.n538 585
R215 B.n537 B.n45 585
R216 B.n536 B.n535 585
R217 B.n534 B.n46 585
R218 B.n533 B.n532 585
R219 B.n530 B.n47 585
R220 B.n529 B.n528 585
R221 B.n527 B.n50 585
R222 B.n526 B.n525 585
R223 B.n524 B.n51 585
R224 B.n523 B.n522 585
R225 B.n521 B.n52 585
R226 B.n520 B.n519 585
R227 B.n518 B.n53 585
R228 B.n517 B.n516 585
R229 B.n515 B.n54 585
R230 B.n514 B.n513 585
R231 B.n512 B.n55 585
R232 B.n511 B.n510 585
R233 B.n509 B.n56 585
R234 B.n508 B.n507 585
R235 B.n506 B.n57 585
R236 B.n505 B.n504 585
R237 B.n503 B.n58 585
R238 B.n502 B.n501 585
R239 B.n500 B.n59 585
R240 B.n499 B.n498 585
R241 B.n497 B.n60 585
R242 B.n496 B.n495 585
R243 B.n494 B.n61 585
R244 B.n493 B.n492 585
R245 B.n491 B.n62 585
R246 B.n490 B.n489 585
R247 B.n488 B.n63 585
R248 B.n487 B.n486 585
R249 B.n485 B.n64 585
R250 B.n484 B.n483 585
R251 B.n482 B.n65 585
R252 B.n481 B.n480 585
R253 B.n479 B.n66 585
R254 B.n478 B.n477 585
R255 B.n476 B.n67 585
R256 B.n475 B.n474 585
R257 B.n473 B.n68 585
R258 B.n472 B.n471 585
R259 B.n470 B.n69 585
R260 B.n469 B.n468 585
R261 B.n467 B.n70 585
R262 B.n466 B.n465 585
R263 B.n464 B.n71 585
R264 B.n463 B.n462 585
R265 B.n461 B.n72 585
R266 B.n617 B.n16 585
R267 B.n619 B.n618 585
R268 B.n620 B.n15 585
R269 B.n622 B.n621 585
R270 B.n623 B.n14 585
R271 B.n625 B.n624 585
R272 B.n626 B.n13 585
R273 B.n628 B.n627 585
R274 B.n629 B.n12 585
R275 B.n631 B.n630 585
R276 B.n632 B.n11 585
R277 B.n634 B.n633 585
R278 B.n635 B.n10 585
R279 B.n637 B.n636 585
R280 B.n638 B.n9 585
R281 B.n640 B.n639 585
R282 B.n641 B.n8 585
R283 B.n643 B.n642 585
R284 B.n644 B.n7 585
R285 B.n646 B.n645 585
R286 B.n647 B.n6 585
R287 B.n649 B.n648 585
R288 B.n650 B.n5 585
R289 B.n652 B.n651 585
R290 B.n653 B.n4 585
R291 B.n655 B.n654 585
R292 B.n656 B.n3 585
R293 B.n658 B.n657 585
R294 B.n659 B.n0 585
R295 B.n2 B.n1 585
R296 B.n173 B.n172 585
R297 B.n175 B.n174 585
R298 B.n176 B.n171 585
R299 B.n178 B.n177 585
R300 B.n179 B.n170 585
R301 B.n181 B.n180 585
R302 B.n182 B.n169 585
R303 B.n184 B.n183 585
R304 B.n185 B.n168 585
R305 B.n187 B.n186 585
R306 B.n188 B.n167 585
R307 B.n190 B.n189 585
R308 B.n191 B.n166 585
R309 B.n193 B.n192 585
R310 B.n194 B.n165 585
R311 B.n196 B.n195 585
R312 B.n197 B.n164 585
R313 B.n199 B.n198 585
R314 B.n200 B.n163 585
R315 B.n202 B.n201 585
R316 B.n203 B.n162 585
R317 B.n205 B.n204 585
R318 B.n206 B.n161 585
R319 B.n208 B.n207 585
R320 B.n209 B.n160 585
R321 B.n211 B.n210 585
R322 B.n212 B.n159 585
R323 B.n214 B.n213 585
R324 B.n215 B.n214 526.135
R325 B.n371 B.n370 526.135
R326 B.n461 B.n460 526.135
R327 B.n617 B.n616 526.135
R328 B.n134 B.t0 500.839
R329 B.n126 B.t3 500.839
R330 B.n48 B.t9 500.839
R331 B.n40 B.t6 500.839
R332 B.n661 B.n660 256.663
R333 B.n660 B.n659 235.042
R334 B.n660 B.n2 235.042
R335 B.n216 B.n215 163.367
R336 B.n216 B.n157 163.367
R337 B.n220 B.n157 163.367
R338 B.n221 B.n220 163.367
R339 B.n222 B.n221 163.367
R340 B.n222 B.n155 163.367
R341 B.n226 B.n155 163.367
R342 B.n227 B.n226 163.367
R343 B.n228 B.n227 163.367
R344 B.n228 B.n153 163.367
R345 B.n232 B.n153 163.367
R346 B.n233 B.n232 163.367
R347 B.n234 B.n233 163.367
R348 B.n234 B.n151 163.367
R349 B.n238 B.n151 163.367
R350 B.n239 B.n238 163.367
R351 B.n240 B.n239 163.367
R352 B.n240 B.n149 163.367
R353 B.n244 B.n149 163.367
R354 B.n245 B.n244 163.367
R355 B.n246 B.n245 163.367
R356 B.n246 B.n147 163.367
R357 B.n250 B.n147 163.367
R358 B.n251 B.n250 163.367
R359 B.n252 B.n251 163.367
R360 B.n252 B.n145 163.367
R361 B.n256 B.n145 163.367
R362 B.n257 B.n256 163.367
R363 B.n258 B.n257 163.367
R364 B.n258 B.n143 163.367
R365 B.n262 B.n143 163.367
R366 B.n263 B.n262 163.367
R367 B.n264 B.n263 163.367
R368 B.n264 B.n141 163.367
R369 B.n268 B.n141 163.367
R370 B.n269 B.n268 163.367
R371 B.n270 B.n269 163.367
R372 B.n270 B.n139 163.367
R373 B.n274 B.n139 163.367
R374 B.n275 B.n274 163.367
R375 B.n276 B.n275 163.367
R376 B.n276 B.n137 163.367
R377 B.n280 B.n137 163.367
R378 B.n281 B.n280 163.367
R379 B.n282 B.n281 163.367
R380 B.n282 B.n133 163.367
R381 B.n287 B.n133 163.367
R382 B.n288 B.n287 163.367
R383 B.n289 B.n288 163.367
R384 B.n289 B.n131 163.367
R385 B.n293 B.n131 163.367
R386 B.n294 B.n293 163.367
R387 B.n295 B.n294 163.367
R388 B.n295 B.n129 163.367
R389 B.n299 B.n129 163.367
R390 B.n300 B.n299 163.367
R391 B.n300 B.n125 163.367
R392 B.n304 B.n125 163.367
R393 B.n305 B.n304 163.367
R394 B.n306 B.n305 163.367
R395 B.n306 B.n123 163.367
R396 B.n310 B.n123 163.367
R397 B.n311 B.n310 163.367
R398 B.n312 B.n311 163.367
R399 B.n312 B.n121 163.367
R400 B.n316 B.n121 163.367
R401 B.n317 B.n316 163.367
R402 B.n318 B.n317 163.367
R403 B.n318 B.n119 163.367
R404 B.n322 B.n119 163.367
R405 B.n323 B.n322 163.367
R406 B.n324 B.n323 163.367
R407 B.n324 B.n117 163.367
R408 B.n328 B.n117 163.367
R409 B.n329 B.n328 163.367
R410 B.n330 B.n329 163.367
R411 B.n330 B.n115 163.367
R412 B.n334 B.n115 163.367
R413 B.n335 B.n334 163.367
R414 B.n336 B.n335 163.367
R415 B.n336 B.n113 163.367
R416 B.n340 B.n113 163.367
R417 B.n341 B.n340 163.367
R418 B.n342 B.n341 163.367
R419 B.n342 B.n111 163.367
R420 B.n346 B.n111 163.367
R421 B.n347 B.n346 163.367
R422 B.n348 B.n347 163.367
R423 B.n348 B.n109 163.367
R424 B.n352 B.n109 163.367
R425 B.n353 B.n352 163.367
R426 B.n354 B.n353 163.367
R427 B.n354 B.n107 163.367
R428 B.n358 B.n107 163.367
R429 B.n359 B.n358 163.367
R430 B.n360 B.n359 163.367
R431 B.n360 B.n105 163.367
R432 B.n364 B.n105 163.367
R433 B.n365 B.n364 163.367
R434 B.n366 B.n365 163.367
R435 B.n366 B.n103 163.367
R436 B.n370 B.n103 163.367
R437 B.n460 B.n73 163.367
R438 B.n456 B.n73 163.367
R439 B.n456 B.n455 163.367
R440 B.n455 B.n454 163.367
R441 B.n454 B.n75 163.367
R442 B.n450 B.n75 163.367
R443 B.n450 B.n449 163.367
R444 B.n449 B.n448 163.367
R445 B.n448 B.n77 163.367
R446 B.n444 B.n77 163.367
R447 B.n444 B.n443 163.367
R448 B.n443 B.n442 163.367
R449 B.n442 B.n79 163.367
R450 B.n438 B.n79 163.367
R451 B.n438 B.n437 163.367
R452 B.n437 B.n436 163.367
R453 B.n436 B.n81 163.367
R454 B.n432 B.n81 163.367
R455 B.n432 B.n431 163.367
R456 B.n431 B.n430 163.367
R457 B.n430 B.n83 163.367
R458 B.n426 B.n83 163.367
R459 B.n426 B.n425 163.367
R460 B.n425 B.n424 163.367
R461 B.n424 B.n85 163.367
R462 B.n420 B.n85 163.367
R463 B.n420 B.n419 163.367
R464 B.n419 B.n418 163.367
R465 B.n418 B.n87 163.367
R466 B.n414 B.n87 163.367
R467 B.n414 B.n413 163.367
R468 B.n413 B.n412 163.367
R469 B.n412 B.n89 163.367
R470 B.n408 B.n89 163.367
R471 B.n408 B.n407 163.367
R472 B.n407 B.n406 163.367
R473 B.n406 B.n91 163.367
R474 B.n402 B.n91 163.367
R475 B.n402 B.n401 163.367
R476 B.n401 B.n400 163.367
R477 B.n400 B.n93 163.367
R478 B.n396 B.n93 163.367
R479 B.n396 B.n395 163.367
R480 B.n395 B.n394 163.367
R481 B.n394 B.n95 163.367
R482 B.n390 B.n95 163.367
R483 B.n390 B.n389 163.367
R484 B.n389 B.n388 163.367
R485 B.n388 B.n97 163.367
R486 B.n384 B.n97 163.367
R487 B.n384 B.n383 163.367
R488 B.n383 B.n382 163.367
R489 B.n382 B.n99 163.367
R490 B.n378 B.n99 163.367
R491 B.n378 B.n377 163.367
R492 B.n377 B.n376 163.367
R493 B.n376 B.n101 163.367
R494 B.n372 B.n101 163.367
R495 B.n372 B.n371 163.367
R496 B.n616 B.n17 163.367
R497 B.n612 B.n17 163.367
R498 B.n612 B.n611 163.367
R499 B.n611 B.n610 163.367
R500 B.n610 B.n19 163.367
R501 B.n606 B.n19 163.367
R502 B.n606 B.n605 163.367
R503 B.n605 B.n604 163.367
R504 B.n604 B.n21 163.367
R505 B.n600 B.n21 163.367
R506 B.n600 B.n599 163.367
R507 B.n599 B.n598 163.367
R508 B.n598 B.n23 163.367
R509 B.n594 B.n23 163.367
R510 B.n594 B.n593 163.367
R511 B.n593 B.n592 163.367
R512 B.n592 B.n25 163.367
R513 B.n588 B.n25 163.367
R514 B.n588 B.n587 163.367
R515 B.n587 B.n586 163.367
R516 B.n586 B.n27 163.367
R517 B.n582 B.n27 163.367
R518 B.n582 B.n581 163.367
R519 B.n581 B.n580 163.367
R520 B.n580 B.n29 163.367
R521 B.n576 B.n29 163.367
R522 B.n576 B.n575 163.367
R523 B.n575 B.n574 163.367
R524 B.n574 B.n31 163.367
R525 B.n570 B.n31 163.367
R526 B.n570 B.n569 163.367
R527 B.n569 B.n568 163.367
R528 B.n568 B.n33 163.367
R529 B.n564 B.n33 163.367
R530 B.n564 B.n563 163.367
R531 B.n563 B.n562 163.367
R532 B.n562 B.n35 163.367
R533 B.n558 B.n35 163.367
R534 B.n558 B.n557 163.367
R535 B.n557 B.n556 163.367
R536 B.n556 B.n37 163.367
R537 B.n552 B.n37 163.367
R538 B.n552 B.n551 163.367
R539 B.n551 B.n550 163.367
R540 B.n550 B.n39 163.367
R541 B.n546 B.n39 163.367
R542 B.n546 B.n545 163.367
R543 B.n545 B.n43 163.367
R544 B.n541 B.n43 163.367
R545 B.n541 B.n540 163.367
R546 B.n540 B.n539 163.367
R547 B.n539 B.n45 163.367
R548 B.n535 B.n45 163.367
R549 B.n535 B.n534 163.367
R550 B.n534 B.n533 163.367
R551 B.n533 B.n47 163.367
R552 B.n528 B.n47 163.367
R553 B.n528 B.n527 163.367
R554 B.n527 B.n526 163.367
R555 B.n526 B.n51 163.367
R556 B.n522 B.n51 163.367
R557 B.n522 B.n521 163.367
R558 B.n521 B.n520 163.367
R559 B.n520 B.n53 163.367
R560 B.n516 B.n53 163.367
R561 B.n516 B.n515 163.367
R562 B.n515 B.n514 163.367
R563 B.n514 B.n55 163.367
R564 B.n510 B.n55 163.367
R565 B.n510 B.n509 163.367
R566 B.n509 B.n508 163.367
R567 B.n508 B.n57 163.367
R568 B.n504 B.n57 163.367
R569 B.n504 B.n503 163.367
R570 B.n503 B.n502 163.367
R571 B.n502 B.n59 163.367
R572 B.n498 B.n59 163.367
R573 B.n498 B.n497 163.367
R574 B.n497 B.n496 163.367
R575 B.n496 B.n61 163.367
R576 B.n492 B.n61 163.367
R577 B.n492 B.n491 163.367
R578 B.n491 B.n490 163.367
R579 B.n490 B.n63 163.367
R580 B.n486 B.n63 163.367
R581 B.n486 B.n485 163.367
R582 B.n485 B.n484 163.367
R583 B.n484 B.n65 163.367
R584 B.n480 B.n65 163.367
R585 B.n480 B.n479 163.367
R586 B.n479 B.n478 163.367
R587 B.n478 B.n67 163.367
R588 B.n474 B.n67 163.367
R589 B.n474 B.n473 163.367
R590 B.n473 B.n472 163.367
R591 B.n472 B.n69 163.367
R592 B.n468 B.n69 163.367
R593 B.n468 B.n467 163.367
R594 B.n467 B.n466 163.367
R595 B.n466 B.n71 163.367
R596 B.n462 B.n71 163.367
R597 B.n462 B.n461 163.367
R598 B.n618 B.n617 163.367
R599 B.n618 B.n15 163.367
R600 B.n622 B.n15 163.367
R601 B.n623 B.n622 163.367
R602 B.n624 B.n623 163.367
R603 B.n624 B.n13 163.367
R604 B.n628 B.n13 163.367
R605 B.n629 B.n628 163.367
R606 B.n630 B.n629 163.367
R607 B.n630 B.n11 163.367
R608 B.n634 B.n11 163.367
R609 B.n635 B.n634 163.367
R610 B.n636 B.n635 163.367
R611 B.n636 B.n9 163.367
R612 B.n640 B.n9 163.367
R613 B.n641 B.n640 163.367
R614 B.n642 B.n641 163.367
R615 B.n642 B.n7 163.367
R616 B.n646 B.n7 163.367
R617 B.n647 B.n646 163.367
R618 B.n648 B.n647 163.367
R619 B.n648 B.n5 163.367
R620 B.n652 B.n5 163.367
R621 B.n653 B.n652 163.367
R622 B.n654 B.n653 163.367
R623 B.n654 B.n3 163.367
R624 B.n658 B.n3 163.367
R625 B.n659 B.n658 163.367
R626 B.n173 B.n2 163.367
R627 B.n174 B.n173 163.367
R628 B.n174 B.n171 163.367
R629 B.n178 B.n171 163.367
R630 B.n179 B.n178 163.367
R631 B.n180 B.n179 163.367
R632 B.n180 B.n169 163.367
R633 B.n184 B.n169 163.367
R634 B.n185 B.n184 163.367
R635 B.n186 B.n185 163.367
R636 B.n186 B.n167 163.367
R637 B.n190 B.n167 163.367
R638 B.n191 B.n190 163.367
R639 B.n192 B.n191 163.367
R640 B.n192 B.n165 163.367
R641 B.n196 B.n165 163.367
R642 B.n197 B.n196 163.367
R643 B.n198 B.n197 163.367
R644 B.n198 B.n163 163.367
R645 B.n202 B.n163 163.367
R646 B.n203 B.n202 163.367
R647 B.n204 B.n203 163.367
R648 B.n204 B.n161 163.367
R649 B.n208 B.n161 163.367
R650 B.n209 B.n208 163.367
R651 B.n210 B.n209 163.367
R652 B.n210 B.n159 163.367
R653 B.n214 B.n159 163.367
R654 B.n126 B.t4 138.941
R655 B.n48 B.t11 138.941
R656 B.n134 B.t1 138.924
R657 B.n40 B.t8 138.924
R658 B.n127 B.t5 110.82
R659 B.n49 B.t10 110.82
R660 B.n135 B.t2 110.802
R661 B.n41 B.t7 110.802
R662 B.n285 B.n135 59.5399
R663 B.n128 B.n127 59.5399
R664 B.n531 B.n49 59.5399
R665 B.n42 B.n41 59.5399
R666 B.n615 B.n16 34.1859
R667 B.n459 B.n72 34.1859
R668 B.n369 B.n102 34.1859
R669 B.n213 B.n158 34.1859
R670 B.n135 B.n134 28.1217
R671 B.n127 B.n126 28.1217
R672 B.n49 B.n48 28.1217
R673 B.n41 B.n40 28.1217
R674 B B.n661 18.0485
R675 B.n619 B.n16 10.6151
R676 B.n620 B.n619 10.6151
R677 B.n621 B.n620 10.6151
R678 B.n621 B.n14 10.6151
R679 B.n625 B.n14 10.6151
R680 B.n626 B.n625 10.6151
R681 B.n627 B.n626 10.6151
R682 B.n627 B.n12 10.6151
R683 B.n631 B.n12 10.6151
R684 B.n632 B.n631 10.6151
R685 B.n633 B.n632 10.6151
R686 B.n633 B.n10 10.6151
R687 B.n637 B.n10 10.6151
R688 B.n638 B.n637 10.6151
R689 B.n639 B.n638 10.6151
R690 B.n639 B.n8 10.6151
R691 B.n643 B.n8 10.6151
R692 B.n644 B.n643 10.6151
R693 B.n645 B.n644 10.6151
R694 B.n645 B.n6 10.6151
R695 B.n649 B.n6 10.6151
R696 B.n650 B.n649 10.6151
R697 B.n651 B.n650 10.6151
R698 B.n651 B.n4 10.6151
R699 B.n655 B.n4 10.6151
R700 B.n656 B.n655 10.6151
R701 B.n657 B.n656 10.6151
R702 B.n657 B.n0 10.6151
R703 B.n615 B.n614 10.6151
R704 B.n614 B.n613 10.6151
R705 B.n613 B.n18 10.6151
R706 B.n609 B.n18 10.6151
R707 B.n609 B.n608 10.6151
R708 B.n608 B.n607 10.6151
R709 B.n607 B.n20 10.6151
R710 B.n603 B.n20 10.6151
R711 B.n603 B.n602 10.6151
R712 B.n602 B.n601 10.6151
R713 B.n601 B.n22 10.6151
R714 B.n597 B.n22 10.6151
R715 B.n597 B.n596 10.6151
R716 B.n596 B.n595 10.6151
R717 B.n595 B.n24 10.6151
R718 B.n591 B.n24 10.6151
R719 B.n591 B.n590 10.6151
R720 B.n590 B.n589 10.6151
R721 B.n589 B.n26 10.6151
R722 B.n585 B.n26 10.6151
R723 B.n585 B.n584 10.6151
R724 B.n584 B.n583 10.6151
R725 B.n583 B.n28 10.6151
R726 B.n579 B.n28 10.6151
R727 B.n579 B.n578 10.6151
R728 B.n578 B.n577 10.6151
R729 B.n577 B.n30 10.6151
R730 B.n573 B.n30 10.6151
R731 B.n573 B.n572 10.6151
R732 B.n572 B.n571 10.6151
R733 B.n571 B.n32 10.6151
R734 B.n567 B.n32 10.6151
R735 B.n567 B.n566 10.6151
R736 B.n566 B.n565 10.6151
R737 B.n565 B.n34 10.6151
R738 B.n561 B.n34 10.6151
R739 B.n561 B.n560 10.6151
R740 B.n560 B.n559 10.6151
R741 B.n559 B.n36 10.6151
R742 B.n555 B.n36 10.6151
R743 B.n555 B.n554 10.6151
R744 B.n554 B.n553 10.6151
R745 B.n553 B.n38 10.6151
R746 B.n549 B.n38 10.6151
R747 B.n549 B.n548 10.6151
R748 B.n548 B.n547 10.6151
R749 B.n544 B.n543 10.6151
R750 B.n543 B.n542 10.6151
R751 B.n542 B.n44 10.6151
R752 B.n538 B.n44 10.6151
R753 B.n538 B.n537 10.6151
R754 B.n537 B.n536 10.6151
R755 B.n536 B.n46 10.6151
R756 B.n532 B.n46 10.6151
R757 B.n530 B.n529 10.6151
R758 B.n529 B.n50 10.6151
R759 B.n525 B.n50 10.6151
R760 B.n525 B.n524 10.6151
R761 B.n524 B.n523 10.6151
R762 B.n523 B.n52 10.6151
R763 B.n519 B.n52 10.6151
R764 B.n519 B.n518 10.6151
R765 B.n518 B.n517 10.6151
R766 B.n517 B.n54 10.6151
R767 B.n513 B.n54 10.6151
R768 B.n513 B.n512 10.6151
R769 B.n512 B.n511 10.6151
R770 B.n511 B.n56 10.6151
R771 B.n507 B.n56 10.6151
R772 B.n507 B.n506 10.6151
R773 B.n506 B.n505 10.6151
R774 B.n505 B.n58 10.6151
R775 B.n501 B.n58 10.6151
R776 B.n501 B.n500 10.6151
R777 B.n500 B.n499 10.6151
R778 B.n499 B.n60 10.6151
R779 B.n495 B.n60 10.6151
R780 B.n495 B.n494 10.6151
R781 B.n494 B.n493 10.6151
R782 B.n493 B.n62 10.6151
R783 B.n489 B.n62 10.6151
R784 B.n489 B.n488 10.6151
R785 B.n488 B.n487 10.6151
R786 B.n487 B.n64 10.6151
R787 B.n483 B.n64 10.6151
R788 B.n483 B.n482 10.6151
R789 B.n482 B.n481 10.6151
R790 B.n481 B.n66 10.6151
R791 B.n477 B.n66 10.6151
R792 B.n477 B.n476 10.6151
R793 B.n476 B.n475 10.6151
R794 B.n475 B.n68 10.6151
R795 B.n471 B.n68 10.6151
R796 B.n471 B.n470 10.6151
R797 B.n470 B.n469 10.6151
R798 B.n469 B.n70 10.6151
R799 B.n465 B.n70 10.6151
R800 B.n465 B.n464 10.6151
R801 B.n464 B.n463 10.6151
R802 B.n463 B.n72 10.6151
R803 B.n459 B.n458 10.6151
R804 B.n458 B.n457 10.6151
R805 B.n457 B.n74 10.6151
R806 B.n453 B.n74 10.6151
R807 B.n453 B.n452 10.6151
R808 B.n452 B.n451 10.6151
R809 B.n451 B.n76 10.6151
R810 B.n447 B.n76 10.6151
R811 B.n447 B.n446 10.6151
R812 B.n446 B.n445 10.6151
R813 B.n445 B.n78 10.6151
R814 B.n441 B.n78 10.6151
R815 B.n441 B.n440 10.6151
R816 B.n440 B.n439 10.6151
R817 B.n439 B.n80 10.6151
R818 B.n435 B.n80 10.6151
R819 B.n435 B.n434 10.6151
R820 B.n434 B.n433 10.6151
R821 B.n433 B.n82 10.6151
R822 B.n429 B.n82 10.6151
R823 B.n429 B.n428 10.6151
R824 B.n428 B.n427 10.6151
R825 B.n427 B.n84 10.6151
R826 B.n423 B.n84 10.6151
R827 B.n423 B.n422 10.6151
R828 B.n422 B.n421 10.6151
R829 B.n421 B.n86 10.6151
R830 B.n417 B.n86 10.6151
R831 B.n417 B.n416 10.6151
R832 B.n416 B.n415 10.6151
R833 B.n415 B.n88 10.6151
R834 B.n411 B.n88 10.6151
R835 B.n411 B.n410 10.6151
R836 B.n410 B.n409 10.6151
R837 B.n409 B.n90 10.6151
R838 B.n405 B.n90 10.6151
R839 B.n405 B.n404 10.6151
R840 B.n404 B.n403 10.6151
R841 B.n403 B.n92 10.6151
R842 B.n399 B.n92 10.6151
R843 B.n399 B.n398 10.6151
R844 B.n398 B.n397 10.6151
R845 B.n397 B.n94 10.6151
R846 B.n393 B.n94 10.6151
R847 B.n393 B.n392 10.6151
R848 B.n392 B.n391 10.6151
R849 B.n391 B.n96 10.6151
R850 B.n387 B.n96 10.6151
R851 B.n387 B.n386 10.6151
R852 B.n386 B.n385 10.6151
R853 B.n385 B.n98 10.6151
R854 B.n381 B.n98 10.6151
R855 B.n381 B.n380 10.6151
R856 B.n380 B.n379 10.6151
R857 B.n379 B.n100 10.6151
R858 B.n375 B.n100 10.6151
R859 B.n375 B.n374 10.6151
R860 B.n374 B.n373 10.6151
R861 B.n373 B.n102 10.6151
R862 B.n172 B.n1 10.6151
R863 B.n175 B.n172 10.6151
R864 B.n176 B.n175 10.6151
R865 B.n177 B.n176 10.6151
R866 B.n177 B.n170 10.6151
R867 B.n181 B.n170 10.6151
R868 B.n182 B.n181 10.6151
R869 B.n183 B.n182 10.6151
R870 B.n183 B.n168 10.6151
R871 B.n187 B.n168 10.6151
R872 B.n188 B.n187 10.6151
R873 B.n189 B.n188 10.6151
R874 B.n189 B.n166 10.6151
R875 B.n193 B.n166 10.6151
R876 B.n194 B.n193 10.6151
R877 B.n195 B.n194 10.6151
R878 B.n195 B.n164 10.6151
R879 B.n199 B.n164 10.6151
R880 B.n200 B.n199 10.6151
R881 B.n201 B.n200 10.6151
R882 B.n201 B.n162 10.6151
R883 B.n205 B.n162 10.6151
R884 B.n206 B.n205 10.6151
R885 B.n207 B.n206 10.6151
R886 B.n207 B.n160 10.6151
R887 B.n211 B.n160 10.6151
R888 B.n212 B.n211 10.6151
R889 B.n213 B.n212 10.6151
R890 B.n217 B.n158 10.6151
R891 B.n218 B.n217 10.6151
R892 B.n219 B.n218 10.6151
R893 B.n219 B.n156 10.6151
R894 B.n223 B.n156 10.6151
R895 B.n224 B.n223 10.6151
R896 B.n225 B.n224 10.6151
R897 B.n225 B.n154 10.6151
R898 B.n229 B.n154 10.6151
R899 B.n230 B.n229 10.6151
R900 B.n231 B.n230 10.6151
R901 B.n231 B.n152 10.6151
R902 B.n235 B.n152 10.6151
R903 B.n236 B.n235 10.6151
R904 B.n237 B.n236 10.6151
R905 B.n237 B.n150 10.6151
R906 B.n241 B.n150 10.6151
R907 B.n242 B.n241 10.6151
R908 B.n243 B.n242 10.6151
R909 B.n243 B.n148 10.6151
R910 B.n247 B.n148 10.6151
R911 B.n248 B.n247 10.6151
R912 B.n249 B.n248 10.6151
R913 B.n249 B.n146 10.6151
R914 B.n253 B.n146 10.6151
R915 B.n254 B.n253 10.6151
R916 B.n255 B.n254 10.6151
R917 B.n255 B.n144 10.6151
R918 B.n259 B.n144 10.6151
R919 B.n260 B.n259 10.6151
R920 B.n261 B.n260 10.6151
R921 B.n261 B.n142 10.6151
R922 B.n265 B.n142 10.6151
R923 B.n266 B.n265 10.6151
R924 B.n267 B.n266 10.6151
R925 B.n267 B.n140 10.6151
R926 B.n271 B.n140 10.6151
R927 B.n272 B.n271 10.6151
R928 B.n273 B.n272 10.6151
R929 B.n273 B.n138 10.6151
R930 B.n277 B.n138 10.6151
R931 B.n278 B.n277 10.6151
R932 B.n279 B.n278 10.6151
R933 B.n279 B.n136 10.6151
R934 B.n283 B.n136 10.6151
R935 B.n284 B.n283 10.6151
R936 B.n286 B.n132 10.6151
R937 B.n290 B.n132 10.6151
R938 B.n291 B.n290 10.6151
R939 B.n292 B.n291 10.6151
R940 B.n292 B.n130 10.6151
R941 B.n296 B.n130 10.6151
R942 B.n297 B.n296 10.6151
R943 B.n298 B.n297 10.6151
R944 B.n302 B.n301 10.6151
R945 B.n303 B.n302 10.6151
R946 B.n303 B.n124 10.6151
R947 B.n307 B.n124 10.6151
R948 B.n308 B.n307 10.6151
R949 B.n309 B.n308 10.6151
R950 B.n309 B.n122 10.6151
R951 B.n313 B.n122 10.6151
R952 B.n314 B.n313 10.6151
R953 B.n315 B.n314 10.6151
R954 B.n315 B.n120 10.6151
R955 B.n319 B.n120 10.6151
R956 B.n320 B.n319 10.6151
R957 B.n321 B.n320 10.6151
R958 B.n321 B.n118 10.6151
R959 B.n325 B.n118 10.6151
R960 B.n326 B.n325 10.6151
R961 B.n327 B.n326 10.6151
R962 B.n327 B.n116 10.6151
R963 B.n331 B.n116 10.6151
R964 B.n332 B.n331 10.6151
R965 B.n333 B.n332 10.6151
R966 B.n333 B.n114 10.6151
R967 B.n337 B.n114 10.6151
R968 B.n338 B.n337 10.6151
R969 B.n339 B.n338 10.6151
R970 B.n339 B.n112 10.6151
R971 B.n343 B.n112 10.6151
R972 B.n344 B.n343 10.6151
R973 B.n345 B.n344 10.6151
R974 B.n345 B.n110 10.6151
R975 B.n349 B.n110 10.6151
R976 B.n350 B.n349 10.6151
R977 B.n351 B.n350 10.6151
R978 B.n351 B.n108 10.6151
R979 B.n355 B.n108 10.6151
R980 B.n356 B.n355 10.6151
R981 B.n357 B.n356 10.6151
R982 B.n357 B.n106 10.6151
R983 B.n361 B.n106 10.6151
R984 B.n362 B.n361 10.6151
R985 B.n363 B.n362 10.6151
R986 B.n363 B.n104 10.6151
R987 B.n367 B.n104 10.6151
R988 B.n368 B.n367 10.6151
R989 B.n369 B.n368 10.6151
R990 B.n661 B.n0 8.11757
R991 B.n661 B.n1 8.11757
R992 B.n544 B.n42 6.5566
R993 B.n532 B.n531 6.5566
R994 B.n286 B.n285 6.5566
R995 B.n298 B.n128 6.5566
R996 B.n547 B.n42 4.05904
R997 B.n531 B.n530 4.05904
R998 B.n285 B.n284 4.05904
R999 B.n301 B.n128 4.05904
R1000 VP.n7 VP.t7 355.313
R1001 VP.n17 VP.t0 332.452
R1002 VP.n29 VP.t4 332.452
R1003 VP.n15 VP.t6 332.452
R1004 VP.n22 VP.t2 297.163
R1005 VP.n1 VP.t3 297.163
R1006 VP.n5 VP.t5 297.163
R1007 VP.n8 VP.t1 297.163
R1008 VP.n9 VP.n6 161.3
R1009 VP.n11 VP.n10 161.3
R1010 VP.n13 VP.n12 161.3
R1011 VP.n14 VP.n4 161.3
R1012 VP.n28 VP.n0 161.3
R1013 VP.n27 VP.n26 161.3
R1014 VP.n25 VP.n24 161.3
R1015 VP.n23 VP.n2 161.3
R1016 VP.n21 VP.n20 161.3
R1017 VP.n19 VP.n3 161.3
R1018 VP.n16 VP.n15 80.6037
R1019 VP.n30 VP.n29 80.6037
R1020 VP.n18 VP.n17 80.6037
R1021 VP.n24 VP.n23 56.5193
R1022 VP.n10 VP.n9 56.5193
R1023 VP.n17 VP.n3 49.9132
R1024 VP.n29 VP.n28 49.9132
R1025 VP.n15 VP.n14 49.9132
R1026 VP.n18 VP.n16 45.5317
R1027 VP.n8 VP.n7 33.7295
R1028 VP.n7 VP.n6 28.2143
R1029 VP.n21 VP.n3 24.4675
R1030 VP.n28 VP.n27 24.4675
R1031 VP.n14 VP.n13 24.4675
R1032 VP.n23 VP.n22 23.2442
R1033 VP.n24 VP.n1 23.2442
R1034 VP.n10 VP.n5 23.2442
R1035 VP.n9 VP.n8 23.2442
R1036 VP.n22 VP.n21 1.22385
R1037 VP.n27 VP.n1 1.22385
R1038 VP.n13 VP.n5 1.22385
R1039 VP.n16 VP.n4 0.285035
R1040 VP.n19 VP.n18 0.285035
R1041 VP.n30 VP.n0 0.285035
R1042 VP.n11 VP.n6 0.189894
R1043 VP.n12 VP.n11 0.189894
R1044 VP.n12 VP.n4 0.189894
R1045 VP.n20 VP.n19 0.189894
R1046 VP.n20 VP.n2 0.189894
R1047 VP.n25 VP.n2 0.189894
R1048 VP.n26 VP.n25 0.189894
R1049 VP.n26 VP.n0 0.189894
R1050 VP VP.n30 0.146778
R1051 VDD1 VDD1.n0 70.497
R1052 VDD1.n3 VDD1.n2 70.3834
R1053 VDD1.n3 VDD1.n1 70.3834
R1054 VDD1.n5 VDD1.n4 69.8138
R1055 VDD1.n5 VDD1.n3 41.8285
R1056 VDD1.n4 VDD1.t5 2.35423
R1057 VDD1.n4 VDD1.t0 2.35423
R1058 VDD1.n0 VDD1.t6 2.35423
R1059 VDD1.n0 VDD1.t2 2.35423
R1060 VDD1.n2 VDD1.t3 2.35423
R1061 VDD1.n2 VDD1.t1 2.35423
R1062 VDD1.n1 VDD1.t7 2.35423
R1063 VDD1.n1 VDD1.t4 2.35423
R1064 VDD1 VDD1.n5 0.56731
R1065 VTAIL.n14 VTAIL.t9 55.4888
R1066 VTAIL.n11 VTAIL.t8 55.4887
R1067 VTAIL.n10 VTAIL.t6 55.4887
R1068 VTAIL.n7 VTAIL.t0 55.4887
R1069 VTAIL.n15 VTAIL.t4 55.4886
R1070 VTAIL.n2 VTAIL.t1 55.4886
R1071 VTAIL.n3 VTAIL.t11 55.4886
R1072 VTAIL.n6 VTAIL.t15 55.4886
R1073 VTAIL.n13 VTAIL.n12 53.135
R1074 VTAIL.n9 VTAIL.n8 53.135
R1075 VTAIL.n1 VTAIL.n0 53.135
R1076 VTAIL.n5 VTAIL.n4 53.135
R1077 VTAIL.n15 VTAIL.n14 25.5221
R1078 VTAIL.n7 VTAIL.n6 25.5221
R1079 VTAIL.n0 VTAIL.t5 2.35423
R1080 VTAIL.n0 VTAIL.t2 2.35423
R1081 VTAIL.n4 VTAIL.t13 2.35423
R1082 VTAIL.n4 VTAIL.t12 2.35423
R1083 VTAIL.n12 VTAIL.t14 2.35423
R1084 VTAIL.n12 VTAIL.t10 2.35423
R1085 VTAIL.n8 VTAIL.t3 2.35423
R1086 VTAIL.n8 VTAIL.t7 2.35423
R1087 VTAIL.n9 VTAIL.n7 1.2505
R1088 VTAIL.n10 VTAIL.n9 1.2505
R1089 VTAIL.n13 VTAIL.n11 1.2505
R1090 VTAIL.n14 VTAIL.n13 1.2505
R1091 VTAIL.n6 VTAIL.n5 1.2505
R1092 VTAIL.n5 VTAIL.n3 1.2505
R1093 VTAIL.n2 VTAIL.n1 1.2505
R1094 VTAIL VTAIL.n15 1.19231
R1095 VTAIL.n11 VTAIL.n10 0.470328
R1096 VTAIL.n3 VTAIL.n2 0.470328
R1097 VTAIL VTAIL.n1 0.0586897
R1098 VN.n3 VN.t7 355.313
R1099 VN.n16 VN.t1 355.313
R1100 VN.n11 VN.t3 332.452
R1101 VN.n24 VN.t2 332.452
R1102 VN.n4 VN.t6 297.163
R1103 VN.n1 VN.t4 297.163
R1104 VN.n17 VN.t5 297.163
R1105 VN.n14 VN.t0 297.163
R1106 VN.n23 VN.n13 161.3
R1107 VN.n22 VN.n21 161.3
R1108 VN.n20 VN.n19 161.3
R1109 VN.n18 VN.n15 161.3
R1110 VN.n10 VN.n0 161.3
R1111 VN.n9 VN.n8 161.3
R1112 VN.n7 VN.n6 161.3
R1113 VN.n5 VN.n2 161.3
R1114 VN.n25 VN.n24 80.6037
R1115 VN.n12 VN.n11 80.6037
R1116 VN.n6 VN.n5 56.5193
R1117 VN.n19 VN.n18 56.5193
R1118 VN.n11 VN.n10 49.9132
R1119 VN.n24 VN.n23 49.9132
R1120 VN VN.n25 45.8172
R1121 VN.n4 VN.n3 33.7295
R1122 VN.n17 VN.n16 33.7295
R1123 VN.n16 VN.n15 28.2143
R1124 VN.n3 VN.n2 28.2143
R1125 VN.n10 VN.n9 24.4675
R1126 VN.n23 VN.n22 24.4675
R1127 VN.n5 VN.n4 23.2442
R1128 VN.n6 VN.n1 23.2442
R1129 VN.n18 VN.n17 23.2442
R1130 VN.n19 VN.n14 23.2442
R1131 VN.n9 VN.n1 1.22385
R1132 VN.n22 VN.n14 1.22385
R1133 VN.n25 VN.n13 0.285035
R1134 VN.n12 VN.n0 0.285035
R1135 VN.n21 VN.n13 0.189894
R1136 VN.n21 VN.n20 0.189894
R1137 VN.n20 VN.n15 0.189894
R1138 VN.n7 VN.n2 0.189894
R1139 VN.n8 VN.n7 0.189894
R1140 VN.n8 VN.n0 0.189894
R1141 VN VN.n12 0.146778
R1142 VDD2.n2 VDD2.n1 70.3834
R1143 VDD2.n2 VDD2.n0 70.3834
R1144 VDD2 VDD2.n5 70.3806
R1145 VDD2.n4 VDD2.n3 69.8138
R1146 VDD2.n4 VDD2.n2 41.2455
R1147 VDD2.n5 VDD2.t2 2.35423
R1148 VDD2.n5 VDD2.t6 2.35423
R1149 VDD2.n3 VDD2.t5 2.35423
R1150 VDD2.n3 VDD2.t7 2.35423
R1151 VDD2.n1 VDD2.t3 2.35423
R1152 VDD2.n1 VDD2.t4 2.35423
R1153 VDD2.n0 VDD2.t0 2.35423
R1154 VDD2.n0 VDD2.t1 2.35423
R1155 VDD2 VDD2.n4 0.68369
C0 VDD1 VDD2 1.03659f
C1 B VTAIL 4.6757f
C2 VDD1 VTAIL 10.201401f
C3 VP B 1.41277f
C4 w_n2420_n3730# B 8.35751f
C5 VP VDD1 7.99734f
C6 VDD2 VTAIL 10.2459f
C7 w_n2420_n3730# VDD1 1.50755f
C8 VP VDD2 0.362239f
C9 w_n2420_n3730# VDD2 1.55999f
C10 VP VTAIL 7.64763f
C11 w_n2420_n3730# VTAIL 4.59766f
C12 B VN 0.901323f
C13 w_n2420_n3730# VP 4.84735f
C14 VDD1 VN 0.149109f
C15 VN VDD2 7.78486f
C16 VN VTAIL 7.63352f
C17 VDD1 B 1.24714f
C18 VP VN 6.18619f
C19 B VDD2 1.2968f
C20 w_n2420_n3730# VN 4.53755f
C21 VDD2 VSUBS 1.47046f
C22 VDD1 VSUBS 1.853095f
C23 VTAIL VSUBS 1.12194f
C24 VN VSUBS 5.14442f
C25 VP VSUBS 2.159324f
C26 B VSUBS 3.506472f
C27 w_n2420_n3730# VSUBS 0.110846p
C28 VDD2.t0 VSUBS 0.279469f
C29 VDD2.t1 VSUBS 0.279469f
C30 VDD2.n0 VSUBS 2.22654f
C31 VDD2.t3 VSUBS 0.279469f
C32 VDD2.t4 VSUBS 0.279469f
C33 VDD2.n1 VSUBS 2.22654f
C34 VDD2.n2 VSUBS 3.17154f
C35 VDD2.t5 VSUBS 0.279469f
C36 VDD2.t7 VSUBS 0.279469f
C37 VDD2.n3 VSUBS 2.22116f
C38 VDD2.n4 VSUBS 2.93073f
C39 VDD2.t2 VSUBS 0.279469f
C40 VDD2.t6 VSUBS 0.279469f
C41 VDD2.n5 VSUBS 2.22651f
C42 VN.n0 VSUBS 0.057647f
C43 VN.t4 VSUBS 1.82741f
C44 VN.n1 VSUBS 0.663951f
C45 VN.n2 VSUBS 0.22639f
C46 VN.t6 VSUBS 1.82741f
C47 VN.t7 VSUBS 1.9498f
C48 VN.n3 VSUBS 0.721581f
C49 VN.n4 VSUBS 0.733087f
C50 VN.n5 VSUBS 0.061076f
C51 VN.n6 VSUBS 0.061076f
C52 VN.n7 VSUBS 0.043201f
C53 VN.n8 VSUBS 0.043201f
C54 VN.n9 VSUBS 0.04275f
C55 VN.n10 VSUBS 0.054719f
C56 VN.t3 VSUBS 1.90154f
C57 VN.n11 VSUBS 0.739377f
C58 VN.n12 VSUBS 0.04046f
C59 VN.n13 VSUBS 0.057647f
C60 VN.t0 VSUBS 1.82741f
C61 VN.n14 VSUBS 0.663951f
C62 VN.n15 VSUBS 0.22639f
C63 VN.t5 VSUBS 1.82741f
C64 VN.t1 VSUBS 1.9498f
C65 VN.n16 VSUBS 0.721581f
C66 VN.n17 VSUBS 0.733087f
C67 VN.n18 VSUBS 0.061076f
C68 VN.n19 VSUBS 0.061076f
C69 VN.n20 VSUBS 0.043201f
C70 VN.n21 VSUBS 0.043201f
C71 VN.n22 VSUBS 0.04275f
C72 VN.n23 VSUBS 0.054719f
C73 VN.t2 VSUBS 1.90154f
C74 VN.n24 VSUBS 0.739377f
C75 VN.n25 VSUBS 2.07227f
C76 VTAIL.t5 VSUBS 0.260623f
C77 VTAIL.t2 VSUBS 0.260623f
C78 VTAIL.n0 VSUBS 1.9255f
C79 VTAIL.n1 VSUBS 0.683344f
C80 VTAIL.t1 VSUBS 2.53551f
C81 VTAIL.n2 VSUBS 0.815802f
C82 VTAIL.t11 VSUBS 2.53551f
C83 VTAIL.n3 VSUBS 0.815802f
C84 VTAIL.t13 VSUBS 0.260623f
C85 VTAIL.t12 VSUBS 0.260623f
C86 VTAIL.n4 VSUBS 1.9255f
C87 VTAIL.n5 VSUBS 0.775057f
C88 VTAIL.t15 VSUBS 2.53551f
C89 VTAIL.n6 VSUBS 2.11637f
C90 VTAIL.t0 VSUBS 2.53553f
C91 VTAIL.n7 VSUBS 2.11636f
C92 VTAIL.t3 VSUBS 0.260623f
C93 VTAIL.t7 VSUBS 0.260623f
C94 VTAIL.n8 VSUBS 1.9255f
C95 VTAIL.n9 VSUBS 0.775052f
C96 VTAIL.t6 VSUBS 2.53553f
C97 VTAIL.n10 VSUBS 0.815784f
C98 VTAIL.t8 VSUBS 2.53553f
C99 VTAIL.n11 VSUBS 0.815784f
C100 VTAIL.t14 VSUBS 0.260623f
C101 VTAIL.t10 VSUBS 0.260623f
C102 VTAIL.n12 VSUBS 1.9255f
C103 VTAIL.n13 VSUBS 0.775052f
C104 VTAIL.t9 VSUBS 2.53552f
C105 VTAIL.n14 VSUBS 2.11636f
C106 VTAIL.t4 VSUBS 2.53551f
C107 VTAIL.n15 VSUBS 2.1119f
C108 VDD1.t6 VSUBS 0.281097f
C109 VDD1.t2 VSUBS 0.281097f
C110 VDD1.n0 VSUBS 2.24066f
C111 VDD1.t7 VSUBS 0.281097f
C112 VDD1.t4 VSUBS 0.281097f
C113 VDD1.n1 VSUBS 2.23951f
C114 VDD1.t3 VSUBS 0.281097f
C115 VDD1.t1 VSUBS 0.281097f
C116 VDD1.n2 VSUBS 2.23951f
C117 VDD1.n3 VSUBS 3.24456f
C118 VDD1.t5 VSUBS 0.281097f
C119 VDD1.t0 VSUBS 0.281097f
C120 VDD1.n4 VSUBS 2.2341f
C121 VDD1.n5 VSUBS 2.97874f
C122 VP.n0 VSUBS 0.058888f
C123 VP.t3 VSUBS 1.86676f
C124 VP.n1 VSUBS 0.678249f
C125 VP.n2 VSUBS 0.044131f
C126 VP.t2 VSUBS 1.86676f
C127 VP.n3 VSUBS 0.055897f
C128 VP.n4 VSUBS 0.058888f
C129 VP.t6 VSUBS 1.94249f
C130 VP.t5 VSUBS 1.86676f
C131 VP.n5 VSUBS 0.678249f
C132 VP.n6 VSUBS 0.231266f
C133 VP.t1 VSUBS 1.86676f
C134 VP.t7 VSUBS 1.99179f
C135 VP.n7 VSUBS 0.737119f
C136 VP.n8 VSUBS 0.748873f
C137 VP.n9 VSUBS 0.062392f
C138 VP.n10 VSUBS 0.062392f
C139 VP.n11 VSUBS 0.044131f
C140 VP.n12 VSUBS 0.044131f
C141 VP.n13 VSUBS 0.043671f
C142 VP.n14 VSUBS 0.055897f
C143 VP.n15 VSUBS 0.755298f
C144 VP.n16 VSUBS 2.09247f
C145 VP.t0 VSUBS 1.94249f
C146 VP.n17 VSUBS 0.755298f
C147 VP.n18 VSUBS 2.12731f
C148 VP.n19 VSUBS 0.058888f
C149 VP.n20 VSUBS 0.044131f
C150 VP.n21 VSUBS 0.043671f
C151 VP.n22 VSUBS 0.678249f
C152 VP.n23 VSUBS 0.062392f
C153 VP.n24 VSUBS 0.062392f
C154 VP.n25 VSUBS 0.044131f
C155 VP.n26 VSUBS 0.044131f
C156 VP.n27 VSUBS 0.043671f
C157 VP.n28 VSUBS 0.055897f
C158 VP.t4 VSUBS 1.94249f
C159 VP.n29 VSUBS 0.755298f
C160 VP.n30 VSUBS 0.041331f
C161 B.n0 VSUBS 0.006687f
C162 B.n1 VSUBS 0.006687f
C163 B.n2 VSUBS 0.00989f
C164 B.n3 VSUBS 0.007579f
C165 B.n4 VSUBS 0.007579f
C166 B.n5 VSUBS 0.007579f
C167 B.n6 VSUBS 0.007579f
C168 B.n7 VSUBS 0.007579f
C169 B.n8 VSUBS 0.007579f
C170 B.n9 VSUBS 0.007579f
C171 B.n10 VSUBS 0.007579f
C172 B.n11 VSUBS 0.007579f
C173 B.n12 VSUBS 0.007579f
C174 B.n13 VSUBS 0.007579f
C175 B.n14 VSUBS 0.007579f
C176 B.n15 VSUBS 0.007579f
C177 B.n16 VSUBS 0.01808f
C178 B.n17 VSUBS 0.007579f
C179 B.n18 VSUBS 0.007579f
C180 B.n19 VSUBS 0.007579f
C181 B.n20 VSUBS 0.007579f
C182 B.n21 VSUBS 0.007579f
C183 B.n22 VSUBS 0.007579f
C184 B.n23 VSUBS 0.007579f
C185 B.n24 VSUBS 0.007579f
C186 B.n25 VSUBS 0.007579f
C187 B.n26 VSUBS 0.007579f
C188 B.n27 VSUBS 0.007579f
C189 B.n28 VSUBS 0.007579f
C190 B.n29 VSUBS 0.007579f
C191 B.n30 VSUBS 0.007579f
C192 B.n31 VSUBS 0.007579f
C193 B.n32 VSUBS 0.007579f
C194 B.n33 VSUBS 0.007579f
C195 B.n34 VSUBS 0.007579f
C196 B.n35 VSUBS 0.007579f
C197 B.n36 VSUBS 0.007579f
C198 B.n37 VSUBS 0.007579f
C199 B.n38 VSUBS 0.007579f
C200 B.n39 VSUBS 0.007579f
C201 B.t7 VSUBS 0.49413f
C202 B.t8 VSUBS 0.506357f
C203 B.t6 VSUBS 0.708853f
C204 B.n40 VSUBS 0.199151f
C205 B.n41 VSUBS 0.071209f
C206 B.n42 VSUBS 0.017559f
C207 B.n43 VSUBS 0.007579f
C208 B.n44 VSUBS 0.007579f
C209 B.n45 VSUBS 0.007579f
C210 B.n46 VSUBS 0.007579f
C211 B.n47 VSUBS 0.007579f
C212 B.t10 VSUBS 0.494118f
C213 B.t11 VSUBS 0.506346f
C214 B.t9 VSUBS 0.708853f
C215 B.n48 VSUBS 0.199162f
C216 B.n49 VSUBS 0.071221f
C217 B.n50 VSUBS 0.007579f
C218 B.n51 VSUBS 0.007579f
C219 B.n52 VSUBS 0.007579f
C220 B.n53 VSUBS 0.007579f
C221 B.n54 VSUBS 0.007579f
C222 B.n55 VSUBS 0.007579f
C223 B.n56 VSUBS 0.007579f
C224 B.n57 VSUBS 0.007579f
C225 B.n58 VSUBS 0.007579f
C226 B.n59 VSUBS 0.007579f
C227 B.n60 VSUBS 0.007579f
C228 B.n61 VSUBS 0.007579f
C229 B.n62 VSUBS 0.007579f
C230 B.n63 VSUBS 0.007579f
C231 B.n64 VSUBS 0.007579f
C232 B.n65 VSUBS 0.007579f
C233 B.n66 VSUBS 0.007579f
C234 B.n67 VSUBS 0.007579f
C235 B.n68 VSUBS 0.007579f
C236 B.n69 VSUBS 0.007579f
C237 B.n70 VSUBS 0.007579f
C238 B.n71 VSUBS 0.007579f
C239 B.n72 VSUBS 0.018476f
C240 B.n73 VSUBS 0.007579f
C241 B.n74 VSUBS 0.007579f
C242 B.n75 VSUBS 0.007579f
C243 B.n76 VSUBS 0.007579f
C244 B.n77 VSUBS 0.007579f
C245 B.n78 VSUBS 0.007579f
C246 B.n79 VSUBS 0.007579f
C247 B.n80 VSUBS 0.007579f
C248 B.n81 VSUBS 0.007579f
C249 B.n82 VSUBS 0.007579f
C250 B.n83 VSUBS 0.007579f
C251 B.n84 VSUBS 0.007579f
C252 B.n85 VSUBS 0.007579f
C253 B.n86 VSUBS 0.007579f
C254 B.n87 VSUBS 0.007579f
C255 B.n88 VSUBS 0.007579f
C256 B.n89 VSUBS 0.007579f
C257 B.n90 VSUBS 0.007579f
C258 B.n91 VSUBS 0.007579f
C259 B.n92 VSUBS 0.007579f
C260 B.n93 VSUBS 0.007579f
C261 B.n94 VSUBS 0.007579f
C262 B.n95 VSUBS 0.007579f
C263 B.n96 VSUBS 0.007579f
C264 B.n97 VSUBS 0.007579f
C265 B.n98 VSUBS 0.007579f
C266 B.n99 VSUBS 0.007579f
C267 B.n100 VSUBS 0.007579f
C268 B.n101 VSUBS 0.007579f
C269 B.n102 VSUBS 0.018935f
C270 B.n103 VSUBS 0.007579f
C271 B.n104 VSUBS 0.007579f
C272 B.n105 VSUBS 0.007579f
C273 B.n106 VSUBS 0.007579f
C274 B.n107 VSUBS 0.007579f
C275 B.n108 VSUBS 0.007579f
C276 B.n109 VSUBS 0.007579f
C277 B.n110 VSUBS 0.007579f
C278 B.n111 VSUBS 0.007579f
C279 B.n112 VSUBS 0.007579f
C280 B.n113 VSUBS 0.007579f
C281 B.n114 VSUBS 0.007579f
C282 B.n115 VSUBS 0.007579f
C283 B.n116 VSUBS 0.007579f
C284 B.n117 VSUBS 0.007579f
C285 B.n118 VSUBS 0.007579f
C286 B.n119 VSUBS 0.007579f
C287 B.n120 VSUBS 0.007579f
C288 B.n121 VSUBS 0.007579f
C289 B.n122 VSUBS 0.007579f
C290 B.n123 VSUBS 0.007579f
C291 B.n124 VSUBS 0.007579f
C292 B.n125 VSUBS 0.007579f
C293 B.t5 VSUBS 0.494118f
C294 B.t4 VSUBS 0.506346f
C295 B.t3 VSUBS 0.708853f
C296 B.n126 VSUBS 0.199162f
C297 B.n127 VSUBS 0.071221f
C298 B.n128 VSUBS 0.017559f
C299 B.n129 VSUBS 0.007579f
C300 B.n130 VSUBS 0.007579f
C301 B.n131 VSUBS 0.007579f
C302 B.n132 VSUBS 0.007579f
C303 B.n133 VSUBS 0.007579f
C304 B.t2 VSUBS 0.49413f
C305 B.t1 VSUBS 0.506357f
C306 B.t0 VSUBS 0.708853f
C307 B.n134 VSUBS 0.199151f
C308 B.n135 VSUBS 0.071209f
C309 B.n136 VSUBS 0.007579f
C310 B.n137 VSUBS 0.007579f
C311 B.n138 VSUBS 0.007579f
C312 B.n139 VSUBS 0.007579f
C313 B.n140 VSUBS 0.007579f
C314 B.n141 VSUBS 0.007579f
C315 B.n142 VSUBS 0.007579f
C316 B.n143 VSUBS 0.007579f
C317 B.n144 VSUBS 0.007579f
C318 B.n145 VSUBS 0.007579f
C319 B.n146 VSUBS 0.007579f
C320 B.n147 VSUBS 0.007579f
C321 B.n148 VSUBS 0.007579f
C322 B.n149 VSUBS 0.007579f
C323 B.n150 VSUBS 0.007579f
C324 B.n151 VSUBS 0.007579f
C325 B.n152 VSUBS 0.007579f
C326 B.n153 VSUBS 0.007579f
C327 B.n154 VSUBS 0.007579f
C328 B.n155 VSUBS 0.007579f
C329 B.n156 VSUBS 0.007579f
C330 B.n157 VSUBS 0.007579f
C331 B.n158 VSUBS 0.018476f
C332 B.n159 VSUBS 0.007579f
C333 B.n160 VSUBS 0.007579f
C334 B.n161 VSUBS 0.007579f
C335 B.n162 VSUBS 0.007579f
C336 B.n163 VSUBS 0.007579f
C337 B.n164 VSUBS 0.007579f
C338 B.n165 VSUBS 0.007579f
C339 B.n166 VSUBS 0.007579f
C340 B.n167 VSUBS 0.007579f
C341 B.n168 VSUBS 0.007579f
C342 B.n169 VSUBS 0.007579f
C343 B.n170 VSUBS 0.007579f
C344 B.n171 VSUBS 0.007579f
C345 B.n172 VSUBS 0.007579f
C346 B.n173 VSUBS 0.007579f
C347 B.n174 VSUBS 0.007579f
C348 B.n175 VSUBS 0.007579f
C349 B.n176 VSUBS 0.007579f
C350 B.n177 VSUBS 0.007579f
C351 B.n178 VSUBS 0.007579f
C352 B.n179 VSUBS 0.007579f
C353 B.n180 VSUBS 0.007579f
C354 B.n181 VSUBS 0.007579f
C355 B.n182 VSUBS 0.007579f
C356 B.n183 VSUBS 0.007579f
C357 B.n184 VSUBS 0.007579f
C358 B.n185 VSUBS 0.007579f
C359 B.n186 VSUBS 0.007579f
C360 B.n187 VSUBS 0.007579f
C361 B.n188 VSUBS 0.007579f
C362 B.n189 VSUBS 0.007579f
C363 B.n190 VSUBS 0.007579f
C364 B.n191 VSUBS 0.007579f
C365 B.n192 VSUBS 0.007579f
C366 B.n193 VSUBS 0.007579f
C367 B.n194 VSUBS 0.007579f
C368 B.n195 VSUBS 0.007579f
C369 B.n196 VSUBS 0.007579f
C370 B.n197 VSUBS 0.007579f
C371 B.n198 VSUBS 0.007579f
C372 B.n199 VSUBS 0.007579f
C373 B.n200 VSUBS 0.007579f
C374 B.n201 VSUBS 0.007579f
C375 B.n202 VSUBS 0.007579f
C376 B.n203 VSUBS 0.007579f
C377 B.n204 VSUBS 0.007579f
C378 B.n205 VSUBS 0.007579f
C379 B.n206 VSUBS 0.007579f
C380 B.n207 VSUBS 0.007579f
C381 B.n208 VSUBS 0.007579f
C382 B.n209 VSUBS 0.007579f
C383 B.n210 VSUBS 0.007579f
C384 B.n211 VSUBS 0.007579f
C385 B.n212 VSUBS 0.007579f
C386 B.n213 VSUBS 0.01808f
C387 B.n214 VSUBS 0.01808f
C388 B.n215 VSUBS 0.018476f
C389 B.n216 VSUBS 0.007579f
C390 B.n217 VSUBS 0.007579f
C391 B.n218 VSUBS 0.007579f
C392 B.n219 VSUBS 0.007579f
C393 B.n220 VSUBS 0.007579f
C394 B.n221 VSUBS 0.007579f
C395 B.n222 VSUBS 0.007579f
C396 B.n223 VSUBS 0.007579f
C397 B.n224 VSUBS 0.007579f
C398 B.n225 VSUBS 0.007579f
C399 B.n226 VSUBS 0.007579f
C400 B.n227 VSUBS 0.007579f
C401 B.n228 VSUBS 0.007579f
C402 B.n229 VSUBS 0.007579f
C403 B.n230 VSUBS 0.007579f
C404 B.n231 VSUBS 0.007579f
C405 B.n232 VSUBS 0.007579f
C406 B.n233 VSUBS 0.007579f
C407 B.n234 VSUBS 0.007579f
C408 B.n235 VSUBS 0.007579f
C409 B.n236 VSUBS 0.007579f
C410 B.n237 VSUBS 0.007579f
C411 B.n238 VSUBS 0.007579f
C412 B.n239 VSUBS 0.007579f
C413 B.n240 VSUBS 0.007579f
C414 B.n241 VSUBS 0.007579f
C415 B.n242 VSUBS 0.007579f
C416 B.n243 VSUBS 0.007579f
C417 B.n244 VSUBS 0.007579f
C418 B.n245 VSUBS 0.007579f
C419 B.n246 VSUBS 0.007579f
C420 B.n247 VSUBS 0.007579f
C421 B.n248 VSUBS 0.007579f
C422 B.n249 VSUBS 0.007579f
C423 B.n250 VSUBS 0.007579f
C424 B.n251 VSUBS 0.007579f
C425 B.n252 VSUBS 0.007579f
C426 B.n253 VSUBS 0.007579f
C427 B.n254 VSUBS 0.007579f
C428 B.n255 VSUBS 0.007579f
C429 B.n256 VSUBS 0.007579f
C430 B.n257 VSUBS 0.007579f
C431 B.n258 VSUBS 0.007579f
C432 B.n259 VSUBS 0.007579f
C433 B.n260 VSUBS 0.007579f
C434 B.n261 VSUBS 0.007579f
C435 B.n262 VSUBS 0.007579f
C436 B.n263 VSUBS 0.007579f
C437 B.n264 VSUBS 0.007579f
C438 B.n265 VSUBS 0.007579f
C439 B.n266 VSUBS 0.007579f
C440 B.n267 VSUBS 0.007579f
C441 B.n268 VSUBS 0.007579f
C442 B.n269 VSUBS 0.007579f
C443 B.n270 VSUBS 0.007579f
C444 B.n271 VSUBS 0.007579f
C445 B.n272 VSUBS 0.007579f
C446 B.n273 VSUBS 0.007579f
C447 B.n274 VSUBS 0.007579f
C448 B.n275 VSUBS 0.007579f
C449 B.n276 VSUBS 0.007579f
C450 B.n277 VSUBS 0.007579f
C451 B.n278 VSUBS 0.007579f
C452 B.n279 VSUBS 0.007579f
C453 B.n280 VSUBS 0.007579f
C454 B.n281 VSUBS 0.007579f
C455 B.n282 VSUBS 0.007579f
C456 B.n283 VSUBS 0.007579f
C457 B.n284 VSUBS 0.005238f
C458 B.n285 VSUBS 0.017559f
C459 B.n286 VSUBS 0.00613f
C460 B.n287 VSUBS 0.007579f
C461 B.n288 VSUBS 0.007579f
C462 B.n289 VSUBS 0.007579f
C463 B.n290 VSUBS 0.007579f
C464 B.n291 VSUBS 0.007579f
C465 B.n292 VSUBS 0.007579f
C466 B.n293 VSUBS 0.007579f
C467 B.n294 VSUBS 0.007579f
C468 B.n295 VSUBS 0.007579f
C469 B.n296 VSUBS 0.007579f
C470 B.n297 VSUBS 0.007579f
C471 B.n298 VSUBS 0.00613f
C472 B.n299 VSUBS 0.007579f
C473 B.n300 VSUBS 0.007579f
C474 B.n301 VSUBS 0.005238f
C475 B.n302 VSUBS 0.007579f
C476 B.n303 VSUBS 0.007579f
C477 B.n304 VSUBS 0.007579f
C478 B.n305 VSUBS 0.007579f
C479 B.n306 VSUBS 0.007579f
C480 B.n307 VSUBS 0.007579f
C481 B.n308 VSUBS 0.007579f
C482 B.n309 VSUBS 0.007579f
C483 B.n310 VSUBS 0.007579f
C484 B.n311 VSUBS 0.007579f
C485 B.n312 VSUBS 0.007579f
C486 B.n313 VSUBS 0.007579f
C487 B.n314 VSUBS 0.007579f
C488 B.n315 VSUBS 0.007579f
C489 B.n316 VSUBS 0.007579f
C490 B.n317 VSUBS 0.007579f
C491 B.n318 VSUBS 0.007579f
C492 B.n319 VSUBS 0.007579f
C493 B.n320 VSUBS 0.007579f
C494 B.n321 VSUBS 0.007579f
C495 B.n322 VSUBS 0.007579f
C496 B.n323 VSUBS 0.007579f
C497 B.n324 VSUBS 0.007579f
C498 B.n325 VSUBS 0.007579f
C499 B.n326 VSUBS 0.007579f
C500 B.n327 VSUBS 0.007579f
C501 B.n328 VSUBS 0.007579f
C502 B.n329 VSUBS 0.007579f
C503 B.n330 VSUBS 0.007579f
C504 B.n331 VSUBS 0.007579f
C505 B.n332 VSUBS 0.007579f
C506 B.n333 VSUBS 0.007579f
C507 B.n334 VSUBS 0.007579f
C508 B.n335 VSUBS 0.007579f
C509 B.n336 VSUBS 0.007579f
C510 B.n337 VSUBS 0.007579f
C511 B.n338 VSUBS 0.007579f
C512 B.n339 VSUBS 0.007579f
C513 B.n340 VSUBS 0.007579f
C514 B.n341 VSUBS 0.007579f
C515 B.n342 VSUBS 0.007579f
C516 B.n343 VSUBS 0.007579f
C517 B.n344 VSUBS 0.007579f
C518 B.n345 VSUBS 0.007579f
C519 B.n346 VSUBS 0.007579f
C520 B.n347 VSUBS 0.007579f
C521 B.n348 VSUBS 0.007579f
C522 B.n349 VSUBS 0.007579f
C523 B.n350 VSUBS 0.007579f
C524 B.n351 VSUBS 0.007579f
C525 B.n352 VSUBS 0.007579f
C526 B.n353 VSUBS 0.007579f
C527 B.n354 VSUBS 0.007579f
C528 B.n355 VSUBS 0.007579f
C529 B.n356 VSUBS 0.007579f
C530 B.n357 VSUBS 0.007579f
C531 B.n358 VSUBS 0.007579f
C532 B.n359 VSUBS 0.007579f
C533 B.n360 VSUBS 0.007579f
C534 B.n361 VSUBS 0.007579f
C535 B.n362 VSUBS 0.007579f
C536 B.n363 VSUBS 0.007579f
C537 B.n364 VSUBS 0.007579f
C538 B.n365 VSUBS 0.007579f
C539 B.n366 VSUBS 0.007579f
C540 B.n367 VSUBS 0.007579f
C541 B.n368 VSUBS 0.007579f
C542 B.n369 VSUBS 0.017621f
C543 B.n370 VSUBS 0.018476f
C544 B.n371 VSUBS 0.01808f
C545 B.n372 VSUBS 0.007579f
C546 B.n373 VSUBS 0.007579f
C547 B.n374 VSUBS 0.007579f
C548 B.n375 VSUBS 0.007579f
C549 B.n376 VSUBS 0.007579f
C550 B.n377 VSUBS 0.007579f
C551 B.n378 VSUBS 0.007579f
C552 B.n379 VSUBS 0.007579f
C553 B.n380 VSUBS 0.007579f
C554 B.n381 VSUBS 0.007579f
C555 B.n382 VSUBS 0.007579f
C556 B.n383 VSUBS 0.007579f
C557 B.n384 VSUBS 0.007579f
C558 B.n385 VSUBS 0.007579f
C559 B.n386 VSUBS 0.007579f
C560 B.n387 VSUBS 0.007579f
C561 B.n388 VSUBS 0.007579f
C562 B.n389 VSUBS 0.007579f
C563 B.n390 VSUBS 0.007579f
C564 B.n391 VSUBS 0.007579f
C565 B.n392 VSUBS 0.007579f
C566 B.n393 VSUBS 0.007579f
C567 B.n394 VSUBS 0.007579f
C568 B.n395 VSUBS 0.007579f
C569 B.n396 VSUBS 0.007579f
C570 B.n397 VSUBS 0.007579f
C571 B.n398 VSUBS 0.007579f
C572 B.n399 VSUBS 0.007579f
C573 B.n400 VSUBS 0.007579f
C574 B.n401 VSUBS 0.007579f
C575 B.n402 VSUBS 0.007579f
C576 B.n403 VSUBS 0.007579f
C577 B.n404 VSUBS 0.007579f
C578 B.n405 VSUBS 0.007579f
C579 B.n406 VSUBS 0.007579f
C580 B.n407 VSUBS 0.007579f
C581 B.n408 VSUBS 0.007579f
C582 B.n409 VSUBS 0.007579f
C583 B.n410 VSUBS 0.007579f
C584 B.n411 VSUBS 0.007579f
C585 B.n412 VSUBS 0.007579f
C586 B.n413 VSUBS 0.007579f
C587 B.n414 VSUBS 0.007579f
C588 B.n415 VSUBS 0.007579f
C589 B.n416 VSUBS 0.007579f
C590 B.n417 VSUBS 0.007579f
C591 B.n418 VSUBS 0.007579f
C592 B.n419 VSUBS 0.007579f
C593 B.n420 VSUBS 0.007579f
C594 B.n421 VSUBS 0.007579f
C595 B.n422 VSUBS 0.007579f
C596 B.n423 VSUBS 0.007579f
C597 B.n424 VSUBS 0.007579f
C598 B.n425 VSUBS 0.007579f
C599 B.n426 VSUBS 0.007579f
C600 B.n427 VSUBS 0.007579f
C601 B.n428 VSUBS 0.007579f
C602 B.n429 VSUBS 0.007579f
C603 B.n430 VSUBS 0.007579f
C604 B.n431 VSUBS 0.007579f
C605 B.n432 VSUBS 0.007579f
C606 B.n433 VSUBS 0.007579f
C607 B.n434 VSUBS 0.007579f
C608 B.n435 VSUBS 0.007579f
C609 B.n436 VSUBS 0.007579f
C610 B.n437 VSUBS 0.007579f
C611 B.n438 VSUBS 0.007579f
C612 B.n439 VSUBS 0.007579f
C613 B.n440 VSUBS 0.007579f
C614 B.n441 VSUBS 0.007579f
C615 B.n442 VSUBS 0.007579f
C616 B.n443 VSUBS 0.007579f
C617 B.n444 VSUBS 0.007579f
C618 B.n445 VSUBS 0.007579f
C619 B.n446 VSUBS 0.007579f
C620 B.n447 VSUBS 0.007579f
C621 B.n448 VSUBS 0.007579f
C622 B.n449 VSUBS 0.007579f
C623 B.n450 VSUBS 0.007579f
C624 B.n451 VSUBS 0.007579f
C625 B.n452 VSUBS 0.007579f
C626 B.n453 VSUBS 0.007579f
C627 B.n454 VSUBS 0.007579f
C628 B.n455 VSUBS 0.007579f
C629 B.n456 VSUBS 0.007579f
C630 B.n457 VSUBS 0.007579f
C631 B.n458 VSUBS 0.007579f
C632 B.n459 VSUBS 0.01808f
C633 B.n460 VSUBS 0.01808f
C634 B.n461 VSUBS 0.018476f
C635 B.n462 VSUBS 0.007579f
C636 B.n463 VSUBS 0.007579f
C637 B.n464 VSUBS 0.007579f
C638 B.n465 VSUBS 0.007579f
C639 B.n466 VSUBS 0.007579f
C640 B.n467 VSUBS 0.007579f
C641 B.n468 VSUBS 0.007579f
C642 B.n469 VSUBS 0.007579f
C643 B.n470 VSUBS 0.007579f
C644 B.n471 VSUBS 0.007579f
C645 B.n472 VSUBS 0.007579f
C646 B.n473 VSUBS 0.007579f
C647 B.n474 VSUBS 0.007579f
C648 B.n475 VSUBS 0.007579f
C649 B.n476 VSUBS 0.007579f
C650 B.n477 VSUBS 0.007579f
C651 B.n478 VSUBS 0.007579f
C652 B.n479 VSUBS 0.007579f
C653 B.n480 VSUBS 0.007579f
C654 B.n481 VSUBS 0.007579f
C655 B.n482 VSUBS 0.007579f
C656 B.n483 VSUBS 0.007579f
C657 B.n484 VSUBS 0.007579f
C658 B.n485 VSUBS 0.007579f
C659 B.n486 VSUBS 0.007579f
C660 B.n487 VSUBS 0.007579f
C661 B.n488 VSUBS 0.007579f
C662 B.n489 VSUBS 0.007579f
C663 B.n490 VSUBS 0.007579f
C664 B.n491 VSUBS 0.007579f
C665 B.n492 VSUBS 0.007579f
C666 B.n493 VSUBS 0.007579f
C667 B.n494 VSUBS 0.007579f
C668 B.n495 VSUBS 0.007579f
C669 B.n496 VSUBS 0.007579f
C670 B.n497 VSUBS 0.007579f
C671 B.n498 VSUBS 0.007579f
C672 B.n499 VSUBS 0.007579f
C673 B.n500 VSUBS 0.007579f
C674 B.n501 VSUBS 0.007579f
C675 B.n502 VSUBS 0.007579f
C676 B.n503 VSUBS 0.007579f
C677 B.n504 VSUBS 0.007579f
C678 B.n505 VSUBS 0.007579f
C679 B.n506 VSUBS 0.007579f
C680 B.n507 VSUBS 0.007579f
C681 B.n508 VSUBS 0.007579f
C682 B.n509 VSUBS 0.007579f
C683 B.n510 VSUBS 0.007579f
C684 B.n511 VSUBS 0.007579f
C685 B.n512 VSUBS 0.007579f
C686 B.n513 VSUBS 0.007579f
C687 B.n514 VSUBS 0.007579f
C688 B.n515 VSUBS 0.007579f
C689 B.n516 VSUBS 0.007579f
C690 B.n517 VSUBS 0.007579f
C691 B.n518 VSUBS 0.007579f
C692 B.n519 VSUBS 0.007579f
C693 B.n520 VSUBS 0.007579f
C694 B.n521 VSUBS 0.007579f
C695 B.n522 VSUBS 0.007579f
C696 B.n523 VSUBS 0.007579f
C697 B.n524 VSUBS 0.007579f
C698 B.n525 VSUBS 0.007579f
C699 B.n526 VSUBS 0.007579f
C700 B.n527 VSUBS 0.007579f
C701 B.n528 VSUBS 0.007579f
C702 B.n529 VSUBS 0.007579f
C703 B.n530 VSUBS 0.005238f
C704 B.n531 VSUBS 0.017559f
C705 B.n532 VSUBS 0.00613f
C706 B.n533 VSUBS 0.007579f
C707 B.n534 VSUBS 0.007579f
C708 B.n535 VSUBS 0.007579f
C709 B.n536 VSUBS 0.007579f
C710 B.n537 VSUBS 0.007579f
C711 B.n538 VSUBS 0.007579f
C712 B.n539 VSUBS 0.007579f
C713 B.n540 VSUBS 0.007579f
C714 B.n541 VSUBS 0.007579f
C715 B.n542 VSUBS 0.007579f
C716 B.n543 VSUBS 0.007579f
C717 B.n544 VSUBS 0.00613f
C718 B.n545 VSUBS 0.007579f
C719 B.n546 VSUBS 0.007579f
C720 B.n547 VSUBS 0.005238f
C721 B.n548 VSUBS 0.007579f
C722 B.n549 VSUBS 0.007579f
C723 B.n550 VSUBS 0.007579f
C724 B.n551 VSUBS 0.007579f
C725 B.n552 VSUBS 0.007579f
C726 B.n553 VSUBS 0.007579f
C727 B.n554 VSUBS 0.007579f
C728 B.n555 VSUBS 0.007579f
C729 B.n556 VSUBS 0.007579f
C730 B.n557 VSUBS 0.007579f
C731 B.n558 VSUBS 0.007579f
C732 B.n559 VSUBS 0.007579f
C733 B.n560 VSUBS 0.007579f
C734 B.n561 VSUBS 0.007579f
C735 B.n562 VSUBS 0.007579f
C736 B.n563 VSUBS 0.007579f
C737 B.n564 VSUBS 0.007579f
C738 B.n565 VSUBS 0.007579f
C739 B.n566 VSUBS 0.007579f
C740 B.n567 VSUBS 0.007579f
C741 B.n568 VSUBS 0.007579f
C742 B.n569 VSUBS 0.007579f
C743 B.n570 VSUBS 0.007579f
C744 B.n571 VSUBS 0.007579f
C745 B.n572 VSUBS 0.007579f
C746 B.n573 VSUBS 0.007579f
C747 B.n574 VSUBS 0.007579f
C748 B.n575 VSUBS 0.007579f
C749 B.n576 VSUBS 0.007579f
C750 B.n577 VSUBS 0.007579f
C751 B.n578 VSUBS 0.007579f
C752 B.n579 VSUBS 0.007579f
C753 B.n580 VSUBS 0.007579f
C754 B.n581 VSUBS 0.007579f
C755 B.n582 VSUBS 0.007579f
C756 B.n583 VSUBS 0.007579f
C757 B.n584 VSUBS 0.007579f
C758 B.n585 VSUBS 0.007579f
C759 B.n586 VSUBS 0.007579f
C760 B.n587 VSUBS 0.007579f
C761 B.n588 VSUBS 0.007579f
C762 B.n589 VSUBS 0.007579f
C763 B.n590 VSUBS 0.007579f
C764 B.n591 VSUBS 0.007579f
C765 B.n592 VSUBS 0.007579f
C766 B.n593 VSUBS 0.007579f
C767 B.n594 VSUBS 0.007579f
C768 B.n595 VSUBS 0.007579f
C769 B.n596 VSUBS 0.007579f
C770 B.n597 VSUBS 0.007579f
C771 B.n598 VSUBS 0.007579f
C772 B.n599 VSUBS 0.007579f
C773 B.n600 VSUBS 0.007579f
C774 B.n601 VSUBS 0.007579f
C775 B.n602 VSUBS 0.007579f
C776 B.n603 VSUBS 0.007579f
C777 B.n604 VSUBS 0.007579f
C778 B.n605 VSUBS 0.007579f
C779 B.n606 VSUBS 0.007579f
C780 B.n607 VSUBS 0.007579f
C781 B.n608 VSUBS 0.007579f
C782 B.n609 VSUBS 0.007579f
C783 B.n610 VSUBS 0.007579f
C784 B.n611 VSUBS 0.007579f
C785 B.n612 VSUBS 0.007579f
C786 B.n613 VSUBS 0.007579f
C787 B.n614 VSUBS 0.007579f
C788 B.n615 VSUBS 0.018476f
C789 B.n616 VSUBS 0.018476f
C790 B.n617 VSUBS 0.01808f
C791 B.n618 VSUBS 0.007579f
C792 B.n619 VSUBS 0.007579f
C793 B.n620 VSUBS 0.007579f
C794 B.n621 VSUBS 0.007579f
C795 B.n622 VSUBS 0.007579f
C796 B.n623 VSUBS 0.007579f
C797 B.n624 VSUBS 0.007579f
C798 B.n625 VSUBS 0.007579f
C799 B.n626 VSUBS 0.007579f
C800 B.n627 VSUBS 0.007579f
C801 B.n628 VSUBS 0.007579f
C802 B.n629 VSUBS 0.007579f
C803 B.n630 VSUBS 0.007579f
C804 B.n631 VSUBS 0.007579f
C805 B.n632 VSUBS 0.007579f
C806 B.n633 VSUBS 0.007579f
C807 B.n634 VSUBS 0.007579f
C808 B.n635 VSUBS 0.007579f
C809 B.n636 VSUBS 0.007579f
C810 B.n637 VSUBS 0.007579f
C811 B.n638 VSUBS 0.007579f
C812 B.n639 VSUBS 0.007579f
C813 B.n640 VSUBS 0.007579f
C814 B.n641 VSUBS 0.007579f
C815 B.n642 VSUBS 0.007579f
C816 B.n643 VSUBS 0.007579f
C817 B.n644 VSUBS 0.007579f
C818 B.n645 VSUBS 0.007579f
C819 B.n646 VSUBS 0.007579f
C820 B.n647 VSUBS 0.007579f
C821 B.n648 VSUBS 0.007579f
C822 B.n649 VSUBS 0.007579f
C823 B.n650 VSUBS 0.007579f
C824 B.n651 VSUBS 0.007579f
C825 B.n652 VSUBS 0.007579f
C826 B.n653 VSUBS 0.007579f
C827 B.n654 VSUBS 0.007579f
C828 B.n655 VSUBS 0.007579f
C829 B.n656 VSUBS 0.007579f
C830 B.n657 VSUBS 0.007579f
C831 B.n658 VSUBS 0.007579f
C832 B.n659 VSUBS 0.00989f
C833 B.n660 VSUBS 0.010535f
C834 B.n661 VSUBS 0.02095f
.ends

