* NGSPICE file created from diff_pair_sample_0305.ext - technology: sky130A

.subckt diff_pair_sample_0305 VTAIL VN VP B VDD2 VDD1
X0 B.t11 B.t9 B.t10 w_n4340_n4328# sky130_fd_pr__pfet_01v8 ad=6.552 pd=34.38 as=0 ps=0 w=16.8 l=3.04
X1 VTAIL.t15 VP.t0 VDD1.t6 w_n4340_n4328# sky130_fd_pr__pfet_01v8 ad=2.772 pd=17.13 as=2.772 ps=17.13 w=16.8 l=3.04
X2 VTAIL.t7 VN.t0 VDD2.t7 w_n4340_n4328# sky130_fd_pr__pfet_01v8 ad=6.552 pd=34.38 as=2.772 ps=17.13 w=16.8 l=3.04
X3 VTAIL.t5 VN.t1 VDD2.t6 w_n4340_n4328# sky130_fd_pr__pfet_01v8 ad=6.552 pd=34.38 as=2.772 ps=17.13 w=16.8 l=3.04
X4 VDD1.t4 VP.t1 VTAIL.t14 w_n4340_n4328# sky130_fd_pr__pfet_01v8 ad=2.772 pd=17.13 as=2.772 ps=17.13 w=16.8 l=3.04
X5 VTAIL.t3 VN.t2 VDD2.t5 w_n4340_n4328# sky130_fd_pr__pfet_01v8 ad=2.772 pd=17.13 as=2.772 ps=17.13 w=16.8 l=3.04
X6 B.t8 B.t6 B.t7 w_n4340_n4328# sky130_fd_pr__pfet_01v8 ad=6.552 pd=34.38 as=0 ps=0 w=16.8 l=3.04
X7 VDD2.t4 VN.t3 VTAIL.t1 w_n4340_n4328# sky130_fd_pr__pfet_01v8 ad=2.772 pd=17.13 as=6.552 ps=34.38 w=16.8 l=3.04
X8 VDD1.t1 VP.t2 VTAIL.t13 w_n4340_n4328# sky130_fd_pr__pfet_01v8 ad=2.772 pd=17.13 as=6.552 ps=34.38 w=16.8 l=3.04
X9 B.t5 B.t3 B.t4 w_n4340_n4328# sky130_fd_pr__pfet_01v8 ad=6.552 pd=34.38 as=0 ps=0 w=16.8 l=3.04
X10 VTAIL.t12 VP.t3 VDD1.t0 w_n4340_n4328# sky130_fd_pr__pfet_01v8 ad=6.552 pd=34.38 as=2.772 ps=17.13 w=16.8 l=3.04
X11 VTAIL.t11 VP.t4 VDD1.t2 w_n4340_n4328# sky130_fd_pr__pfet_01v8 ad=2.772 pd=17.13 as=2.772 ps=17.13 w=16.8 l=3.04
X12 B.t2 B.t0 B.t1 w_n4340_n4328# sky130_fd_pr__pfet_01v8 ad=6.552 pd=34.38 as=0 ps=0 w=16.8 l=3.04
X13 VTAIL.t6 VN.t4 VDD2.t3 w_n4340_n4328# sky130_fd_pr__pfet_01v8 ad=2.772 pd=17.13 as=2.772 ps=17.13 w=16.8 l=3.04
X14 VDD2.t2 VN.t5 VTAIL.t2 w_n4340_n4328# sky130_fd_pr__pfet_01v8 ad=2.772 pd=17.13 as=2.772 ps=17.13 w=16.8 l=3.04
X15 VDD1.t3 VP.t5 VTAIL.t10 w_n4340_n4328# sky130_fd_pr__pfet_01v8 ad=2.772 pd=17.13 as=6.552 ps=34.38 w=16.8 l=3.04
X16 VDD1.t5 VP.t6 VTAIL.t9 w_n4340_n4328# sky130_fd_pr__pfet_01v8 ad=2.772 pd=17.13 as=2.772 ps=17.13 w=16.8 l=3.04
X17 VDD2.t1 VN.t6 VTAIL.t4 w_n4340_n4328# sky130_fd_pr__pfet_01v8 ad=2.772 pd=17.13 as=6.552 ps=34.38 w=16.8 l=3.04
X18 VTAIL.t8 VP.t7 VDD1.t7 w_n4340_n4328# sky130_fd_pr__pfet_01v8 ad=6.552 pd=34.38 as=2.772 ps=17.13 w=16.8 l=3.04
X19 VDD2.t0 VN.t7 VTAIL.t0 w_n4340_n4328# sky130_fd_pr__pfet_01v8 ad=2.772 pd=17.13 as=2.772 ps=17.13 w=16.8 l=3.04
R0 B.n513 B.n154 585
R1 B.n512 B.n511 585
R2 B.n510 B.n155 585
R3 B.n509 B.n508 585
R4 B.n507 B.n156 585
R5 B.n506 B.n505 585
R6 B.n504 B.n157 585
R7 B.n503 B.n502 585
R8 B.n501 B.n158 585
R9 B.n500 B.n499 585
R10 B.n498 B.n159 585
R11 B.n497 B.n496 585
R12 B.n495 B.n160 585
R13 B.n494 B.n493 585
R14 B.n492 B.n161 585
R15 B.n491 B.n490 585
R16 B.n489 B.n162 585
R17 B.n488 B.n487 585
R18 B.n486 B.n163 585
R19 B.n485 B.n484 585
R20 B.n483 B.n164 585
R21 B.n482 B.n481 585
R22 B.n480 B.n165 585
R23 B.n479 B.n478 585
R24 B.n477 B.n166 585
R25 B.n476 B.n475 585
R26 B.n474 B.n167 585
R27 B.n473 B.n472 585
R28 B.n471 B.n168 585
R29 B.n470 B.n469 585
R30 B.n468 B.n169 585
R31 B.n467 B.n466 585
R32 B.n465 B.n170 585
R33 B.n464 B.n463 585
R34 B.n462 B.n171 585
R35 B.n461 B.n460 585
R36 B.n459 B.n172 585
R37 B.n458 B.n457 585
R38 B.n456 B.n173 585
R39 B.n455 B.n454 585
R40 B.n453 B.n174 585
R41 B.n452 B.n451 585
R42 B.n450 B.n175 585
R43 B.n449 B.n448 585
R44 B.n447 B.n176 585
R45 B.n446 B.n445 585
R46 B.n444 B.n177 585
R47 B.n443 B.n442 585
R48 B.n441 B.n178 585
R49 B.n440 B.n439 585
R50 B.n438 B.n179 585
R51 B.n437 B.n436 585
R52 B.n435 B.n180 585
R53 B.n434 B.n433 585
R54 B.n432 B.n181 585
R55 B.n431 B.n430 585
R56 B.n428 B.n182 585
R57 B.n427 B.n426 585
R58 B.n425 B.n185 585
R59 B.n424 B.n423 585
R60 B.n422 B.n186 585
R61 B.n421 B.n420 585
R62 B.n419 B.n187 585
R63 B.n418 B.n417 585
R64 B.n416 B.n188 585
R65 B.n414 B.n413 585
R66 B.n412 B.n191 585
R67 B.n411 B.n410 585
R68 B.n409 B.n192 585
R69 B.n408 B.n407 585
R70 B.n406 B.n193 585
R71 B.n405 B.n404 585
R72 B.n403 B.n194 585
R73 B.n402 B.n401 585
R74 B.n400 B.n195 585
R75 B.n399 B.n398 585
R76 B.n397 B.n196 585
R77 B.n396 B.n395 585
R78 B.n394 B.n197 585
R79 B.n393 B.n392 585
R80 B.n391 B.n198 585
R81 B.n390 B.n389 585
R82 B.n388 B.n199 585
R83 B.n387 B.n386 585
R84 B.n385 B.n200 585
R85 B.n384 B.n383 585
R86 B.n382 B.n201 585
R87 B.n381 B.n380 585
R88 B.n379 B.n202 585
R89 B.n378 B.n377 585
R90 B.n376 B.n203 585
R91 B.n375 B.n374 585
R92 B.n373 B.n204 585
R93 B.n372 B.n371 585
R94 B.n370 B.n205 585
R95 B.n369 B.n368 585
R96 B.n367 B.n206 585
R97 B.n366 B.n365 585
R98 B.n364 B.n207 585
R99 B.n363 B.n362 585
R100 B.n361 B.n208 585
R101 B.n360 B.n359 585
R102 B.n358 B.n209 585
R103 B.n357 B.n356 585
R104 B.n355 B.n210 585
R105 B.n354 B.n353 585
R106 B.n352 B.n211 585
R107 B.n351 B.n350 585
R108 B.n349 B.n212 585
R109 B.n348 B.n347 585
R110 B.n346 B.n213 585
R111 B.n345 B.n344 585
R112 B.n343 B.n214 585
R113 B.n342 B.n341 585
R114 B.n340 B.n215 585
R115 B.n339 B.n338 585
R116 B.n337 B.n216 585
R117 B.n336 B.n335 585
R118 B.n334 B.n217 585
R119 B.n333 B.n332 585
R120 B.n331 B.n218 585
R121 B.n515 B.n514 585
R122 B.n516 B.n153 585
R123 B.n518 B.n517 585
R124 B.n519 B.n152 585
R125 B.n521 B.n520 585
R126 B.n522 B.n151 585
R127 B.n524 B.n523 585
R128 B.n525 B.n150 585
R129 B.n527 B.n526 585
R130 B.n528 B.n149 585
R131 B.n530 B.n529 585
R132 B.n531 B.n148 585
R133 B.n533 B.n532 585
R134 B.n534 B.n147 585
R135 B.n536 B.n535 585
R136 B.n537 B.n146 585
R137 B.n539 B.n538 585
R138 B.n540 B.n145 585
R139 B.n542 B.n541 585
R140 B.n543 B.n144 585
R141 B.n545 B.n544 585
R142 B.n546 B.n143 585
R143 B.n548 B.n547 585
R144 B.n549 B.n142 585
R145 B.n551 B.n550 585
R146 B.n552 B.n141 585
R147 B.n554 B.n553 585
R148 B.n555 B.n140 585
R149 B.n557 B.n556 585
R150 B.n558 B.n139 585
R151 B.n560 B.n559 585
R152 B.n561 B.n138 585
R153 B.n563 B.n562 585
R154 B.n564 B.n137 585
R155 B.n566 B.n565 585
R156 B.n567 B.n136 585
R157 B.n569 B.n568 585
R158 B.n570 B.n135 585
R159 B.n572 B.n571 585
R160 B.n573 B.n134 585
R161 B.n575 B.n574 585
R162 B.n576 B.n133 585
R163 B.n578 B.n577 585
R164 B.n579 B.n132 585
R165 B.n581 B.n580 585
R166 B.n582 B.n131 585
R167 B.n584 B.n583 585
R168 B.n585 B.n130 585
R169 B.n587 B.n586 585
R170 B.n588 B.n129 585
R171 B.n590 B.n589 585
R172 B.n591 B.n128 585
R173 B.n593 B.n592 585
R174 B.n594 B.n127 585
R175 B.n596 B.n595 585
R176 B.n597 B.n126 585
R177 B.n599 B.n598 585
R178 B.n600 B.n125 585
R179 B.n602 B.n601 585
R180 B.n603 B.n124 585
R181 B.n605 B.n604 585
R182 B.n606 B.n123 585
R183 B.n608 B.n607 585
R184 B.n609 B.n122 585
R185 B.n611 B.n610 585
R186 B.n612 B.n121 585
R187 B.n614 B.n613 585
R188 B.n615 B.n120 585
R189 B.n617 B.n616 585
R190 B.n618 B.n119 585
R191 B.n620 B.n619 585
R192 B.n621 B.n118 585
R193 B.n623 B.n622 585
R194 B.n624 B.n117 585
R195 B.n626 B.n625 585
R196 B.n627 B.n116 585
R197 B.n629 B.n628 585
R198 B.n630 B.n115 585
R199 B.n632 B.n631 585
R200 B.n633 B.n114 585
R201 B.n635 B.n634 585
R202 B.n636 B.n113 585
R203 B.n638 B.n637 585
R204 B.n639 B.n112 585
R205 B.n641 B.n640 585
R206 B.n642 B.n111 585
R207 B.n644 B.n643 585
R208 B.n645 B.n110 585
R209 B.n647 B.n646 585
R210 B.n648 B.n109 585
R211 B.n650 B.n649 585
R212 B.n651 B.n108 585
R213 B.n653 B.n652 585
R214 B.n654 B.n107 585
R215 B.n656 B.n655 585
R216 B.n657 B.n106 585
R217 B.n659 B.n658 585
R218 B.n660 B.n105 585
R219 B.n662 B.n661 585
R220 B.n663 B.n104 585
R221 B.n665 B.n664 585
R222 B.n666 B.n103 585
R223 B.n668 B.n667 585
R224 B.n669 B.n102 585
R225 B.n671 B.n670 585
R226 B.n672 B.n101 585
R227 B.n674 B.n673 585
R228 B.n675 B.n100 585
R229 B.n677 B.n676 585
R230 B.n678 B.n99 585
R231 B.n680 B.n679 585
R232 B.n681 B.n98 585
R233 B.n683 B.n682 585
R234 B.n684 B.n97 585
R235 B.n686 B.n685 585
R236 B.n687 B.n96 585
R237 B.n870 B.n869 585
R238 B.n868 B.n31 585
R239 B.n867 B.n866 585
R240 B.n865 B.n32 585
R241 B.n864 B.n863 585
R242 B.n862 B.n33 585
R243 B.n861 B.n860 585
R244 B.n859 B.n34 585
R245 B.n858 B.n857 585
R246 B.n856 B.n35 585
R247 B.n855 B.n854 585
R248 B.n853 B.n36 585
R249 B.n852 B.n851 585
R250 B.n850 B.n37 585
R251 B.n849 B.n848 585
R252 B.n847 B.n38 585
R253 B.n846 B.n845 585
R254 B.n844 B.n39 585
R255 B.n843 B.n842 585
R256 B.n841 B.n40 585
R257 B.n840 B.n839 585
R258 B.n838 B.n41 585
R259 B.n837 B.n836 585
R260 B.n835 B.n42 585
R261 B.n834 B.n833 585
R262 B.n832 B.n43 585
R263 B.n831 B.n830 585
R264 B.n829 B.n44 585
R265 B.n828 B.n827 585
R266 B.n826 B.n45 585
R267 B.n825 B.n824 585
R268 B.n823 B.n46 585
R269 B.n822 B.n821 585
R270 B.n820 B.n47 585
R271 B.n819 B.n818 585
R272 B.n817 B.n48 585
R273 B.n816 B.n815 585
R274 B.n814 B.n49 585
R275 B.n813 B.n812 585
R276 B.n811 B.n50 585
R277 B.n810 B.n809 585
R278 B.n808 B.n51 585
R279 B.n807 B.n806 585
R280 B.n805 B.n52 585
R281 B.n804 B.n803 585
R282 B.n802 B.n53 585
R283 B.n801 B.n800 585
R284 B.n799 B.n54 585
R285 B.n798 B.n797 585
R286 B.n796 B.n55 585
R287 B.n795 B.n794 585
R288 B.n793 B.n56 585
R289 B.n792 B.n791 585
R290 B.n790 B.n57 585
R291 B.n789 B.n788 585
R292 B.n787 B.n58 585
R293 B.n786 B.n785 585
R294 B.n784 B.n59 585
R295 B.n783 B.n782 585
R296 B.n781 B.n63 585
R297 B.n780 B.n779 585
R298 B.n778 B.n64 585
R299 B.n777 B.n776 585
R300 B.n775 B.n65 585
R301 B.n774 B.n773 585
R302 B.n771 B.n66 585
R303 B.n770 B.n769 585
R304 B.n768 B.n69 585
R305 B.n767 B.n766 585
R306 B.n765 B.n70 585
R307 B.n764 B.n763 585
R308 B.n762 B.n71 585
R309 B.n761 B.n760 585
R310 B.n759 B.n72 585
R311 B.n758 B.n757 585
R312 B.n756 B.n73 585
R313 B.n755 B.n754 585
R314 B.n753 B.n74 585
R315 B.n752 B.n751 585
R316 B.n750 B.n75 585
R317 B.n749 B.n748 585
R318 B.n747 B.n76 585
R319 B.n746 B.n745 585
R320 B.n744 B.n77 585
R321 B.n743 B.n742 585
R322 B.n741 B.n78 585
R323 B.n740 B.n739 585
R324 B.n738 B.n79 585
R325 B.n737 B.n736 585
R326 B.n735 B.n80 585
R327 B.n734 B.n733 585
R328 B.n732 B.n81 585
R329 B.n731 B.n730 585
R330 B.n729 B.n82 585
R331 B.n728 B.n727 585
R332 B.n726 B.n83 585
R333 B.n725 B.n724 585
R334 B.n723 B.n84 585
R335 B.n722 B.n721 585
R336 B.n720 B.n85 585
R337 B.n719 B.n718 585
R338 B.n717 B.n86 585
R339 B.n716 B.n715 585
R340 B.n714 B.n87 585
R341 B.n713 B.n712 585
R342 B.n711 B.n88 585
R343 B.n710 B.n709 585
R344 B.n708 B.n89 585
R345 B.n707 B.n706 585
R346 B.n705 B.n90 585
R347 B.n704 B.n703 585
R348 B.n702 B.n91 585
R349 B.n701 B.n700 585
R350 B.n699 B.n92 585
R351 B.n698 B.n697 585
R352 B.n696 B.n93 585
R353 B.n695 B.n694 585
R354 B.n693 B.n94 585
R355 B.n692 B.n691 585
R356 B.n690 B.n95 585
R357 B.n689 B.n688 585
R358 B.n871 B.n30 585
R359 B.n873 B.n872 585
R360 B.n874 B.n29 585
R361 B.n876 B.n875 585
R362 B.n877 B.n28 585
R363 B.n879 B.n878 585
R364 B.n880 B.n27 585
R365 B.n882 B.n881 585
R366 B.n883 B.n26 585
R367 B.n885 B.n884 585
R368 B.n886 B.n25 585
R369 B.n888 B.n887 585
R370 B.n889 B.n24 585
R371 B.n891 B.n890 585
R372 B.n892 B.n23 585
R373 B.n894 B.n893 585
R374 B.n895 B.n22 585
R375 B.n897 B.n896 585
R376 B.n898 B.n21 585
R377 B.n900 B.n899 585
R378 B.n901 B.n20 585
R379 B.n903 B.n902 585
R380 B.n904 B.n19 585
R381 B.n906 B.n905 585
R382 B.n907 B.n18 585
R383 B.n909 B.n908 585
R384 B.n910 B.n17 585
R385 B.n912 B.n911 585
R386 B.n913 B.n16 585
R387 B.n915 B.n914 585
R388 B.n916 B.n15 585
R389 B.n918 B.n917 585
R390 B.n919 B.n14 585
R391 B.n921 B.n920 585
R392 B.n922 B.n13 585
R393 B.n924 B.n923 585
R394 B.n925 B.n12 585
R395 B.n927 B.n926 585
R396 B.n928 B.n11 585
R397 B.n930 B.n929 585
R398 B.n931 B.n10 585
R399 B.n933 B.n932 585
R400 B.n934 B.n9 585
R401 B.n936 B.n935 585
R402 B.n937 B.n8 585
R403 B.n939 B.n938 585
R404 B.n940 B.n7 585
R405 B.n942 B.n941 585
R406 B.n943 B.n6 585
R407 B.n945 B.n944 585
R408 B.n946 B.n5 585
R409 B.n948 B.n947 585
R410 B.n949 B.n4 585
R411 B.n951 B.n950 585
R412 B.n952 B.n3 585
R413 B.n954 B.n953 585
R414 B.n955 B.n0 585
R415 B.n2 B.n1 585
R416 B.n247 B.n246 585
R417 B.n249 B.n248 585
R418 B.n250 B.n245 585
R419 B.n252 B.n251 585
R420 B.n253 B.n244 585
R421 B.n255 B.n254 585
R422 B.n256 B.n243 585
R423 B.n258 B.n257 585
R424 B.n259 B.n242 585
R425 B.n261 B.n260 585
R426 B.n262 B.n241 585
R427 B.n264 B.n263 585
R428 B.n265 B.n240 585
R429 B.n267 B.n266 585
R430 B.n268 B.n239 585
R431 B.n270 B.n269 585
R432 B.n271 B.n238 585
R433 B.n273 B.n272 585
R434 B.n274 B.n237 585
R435 B.n276 B.n275 585
R436 B.n277 B.n236 585
R437 B.n279 B.n278 585
R438 B.n280 B.n235 585
R439 B.n282 B.n281 585
R440 B.n283 B.n234 585
R441 B.n285 B.n284 585
R442 B.n286 B.n233 585
R443 B.n288 B.n287 585
R444 B.n289 B.n232 585
R445 B.n291 B.n290 585
R446 B.n292 B.n231 585
R447 B.n294 B.n293 585
R448 B.n295 B.n230 585
R449 B.n297 B.n296 585
R450 B.n298 B.n229 585
R451 B.n300 B.n299 585
R452 B.n301 B.n228 585
R453 B.n303 B.n302 585
R454 B.n304 B.n227 585
R455 B.n306 B.n305 585
R456 B.n307 B.n226 585
R457 B.n309 B.n308 585
R458 B.n310 B.n225 585
R459 B.n312 B.n311 585
R460 B.n313 B.n224 585
R461 B.n315 B.n314 585
R462 B.n316 B.n223 585
R463 B.n318 B.n317 585
R464 B.n319 B.n222 585
R465 B.n321 B.n320 585
R466 B.n322 B.n221 585
R467 B.n324 B.n323 585
R468 B.n325 B.n220 585
R469 B.n327 B.n326 585
R470 B.n328 B.n219 585
R471 B.n330 B.n329 585
R472 B.n329 B.n218 530.939
R473 B.n515 B.n154 530.939
R474 B.n689 B.n96 530.939
R475 B.n871 B.n870 530.939
R476 B.n183 B.t4 527.399
R477 B.n67 B.t8 527.399
R478 B.n189 B.t10 527.399
R479 B.n60 B.t2 527.399
R480 B.n184 B.t5 462.041
R481 B.n68 B.t7 462.041
R482 B.n190 B.t11 462.041
R483 B.n61 B.t1 462.041
R484 B.n189 B.t9 341.81
R485 B.n183 B.t3 341.81
R486 B.n67 B.t6 341.81
R487 B.n60 B.t0 341.81
R488 B.n957 B.n956 256.663
R489 B.n956 B.n955 235.042
R490 B.n956 B.n2 235.042
R491 B.n333 B.n218 163.367
R492 B.n334 B.n333 163.367
R493 B.n335 B.n334 163.367
R494 B.n335 B.n216 163.367
R495 B.n339 B.n216 163.367
R496 B.n340 B.n339 163.367
R497 B.n341 B.n340 163.367
R498 B.n341 B.n214 163.367
R499 B.n345 B.n214 163.367
R500 B.n346 B.n345 163.367
R501 B.n347 B.n346 163.367
R502 B.n347 B.n212 163.367
R503 B.n351 B.n212 163.367
R504 B.n352 B.n351 163.367
R505 B.n353 B.n352 163.367
R506 B.n353 B.n210 163.367
R507 B.n357 B.n210 163.367
R508 B.n358 B.n357 163.367
R509 B.n359 B.n358 163.367
R510 B.n359 B.n208 163.367
R511 B.n363 B.n208 163.367
R512 B.n364 B.n363 163.367
R513 B.n365 B.n364 163.367
R514 B.n365 B.n206 163.367
R515 B.n369 B.n206 163.367
R516 B.n370 B.n369 163.367
R517 B.n371 B.n370 163.367
R518 B.n371 B.n204 163.367
R519 B.n375 B.n204 163.367
R520 B.n376 B.n375 163.367
R521 B.n377 B.n376 163.367
R522 B.n377 B.n202 163.367
R523 B.n381 B.n202 163.367
R524 B.n382 B.n381 163.367
R525 B.n383 B.n382 163.367
R526 B.n383 B.n200 163.367
R527 B.n387 B.n200 163.367
R528 B.n388 B.n387 163.367
R529 B.n389 B.n388 163.367
R530 B.n389 B.n198 163.367
R531 B.n393 B.n198 163.367
R532 B.n394 B.n393 163.367
R533 B.n395 B.n394 163.367
R534 B.n395 B.n196 163.367
R535 B.n399 B.n196 163.367
R536 B.n400 B.n399 163.367
R537 B.n401 B.n400 163.367
R538 B.n401 B.n194 163.367
R539 B.n405 B.n194 163.367
R540 B.n406 B.n405 163.367
R541 B.n407 B.n406 163.367
R542 B.n407 B.n192 163.367
R543 B.n411 B.n192 163.367
R544 B.n412 B.n411 163.367
R545 B.n413 B.n412 163.367
R546 B.n413 B.n188 163.367
R547 B.n418 B.n188 163.367
R548 B.n419 B.n418 163.367
R549 B.n420 B.n419 163.367
R550 B.n420 B.n186 163.367
R551 B.n424 B.n186 163.367
R552 B.n425 B.n424 163.367
R553 B.n426 B.n425 163.367
R554 B.n426 B.n182 163.367
R555 B.n431 B.n182 163.367
R556 B.n432 B.n431 163.367
R557 B.n433 B.n432 163.367
R558 B.n433 B.n180 163.367
R559 B.n437 B.n180 163.367
R560 B.n438 B.n437 163.367
R561 B.n439 B.n438 163.367
R562 B.n439 B.n178 163.367
R563 B.n443 B.n178 163.367
R564 B.n444 B.n443 163.367
R565 B.n445 B.n444 163.367
R566 B.n445 B.n176 163.367
R567 B.n449 B.n176 163.367
R568 B.n450 B.n449 163.367
R569 B.n451 B.n450 163.367
R570 B.n451 B.n174 163.367
R571 B.n455 B.n174 163.367
R572 B.n456 B.n455 163.367
R573 B.n457 B.n456 163.367
R574 B.n457 B.n172 163.367
R575 B.n461 B.n172 163.367
R576 B.n462 B.n461 163.367
R577 B.n463 B.n462 163.367
R578 B.n463 B.n170 163.367
R579 B.n467 B.n170 163.367
R580 B.n468 B.n467 163.367
R581 B.n469 B.n468 163.367
R582 B.n469 B.n168 163.367
R583 B.n473 B.n168 163.367
R584 B.n474 B.n473 163.367
R585 B.n475 B.n474 163.367
R586 B.n475 B.n166 163.367
R587 B.n479 B.n166 163.367
R588 B.n480 B.n479 163.367
R589 B.n481 B.n480 163.367
R590 B.n481 B.n164 163.367
R591 B.n485 B.n164 163.367
R592 B.n486 B.n485 163.367
R593 B.n487 B.n486 163.367
R594 B.n487 B.n162 163.367
R595 B.n491 B.n162 163.367
R596 B.n492 B.n491 163.367
R597 B.n493 B.n492 163.367
R598 B.n493 B.n160 163.367
R599 B.n497 B.n160 163.367
R600 B.n498 B.n497 163.367
R601 B.n499 B.n498 163.367
R602 B.n499 B.n158 163.367
R603 B.n503 B.n158 163.367
R604 B.n504 B.n503 163.367
R605 B.n505 B.n504 163.367
R606 B.n505 B.n156 163.367
R607 B.n509 B.n156 163.367
R608 B.n510 B.n509 163.367
R609 B.n511 B.n510 163.367
R610 B.n511 B.n154 163.367
R611 B.n685 B.n96 163.367
R612 B.n685 B.n684 163.367
R613 B.n684 B.n683 163.367
R614 B.n683 B.n98 163.367
R615 B.n679 B.n98 163.367
R616 B.n679 B.n678 163.367
R617 B.n678 B.n677 163.367
R618 B.n677 B.n100 163.367
R619 B.n673 B.n100 163.367
R620 B.n673 B.n672 163.367
R621 B.n672 B.n671 163.367
R622 B.n671 B.n102 163.367
R623 B.n667 B.n102 163.367
R624 B.n667 B.n666 163.367
R625 B.n666 B.n665 163.367
R626 B.n665 B.n104 163.367
R627 B.n661 B.n104 163.367
R628 B.n661 B.n660 163.367
R629 B.n660 B.n659 163.367
R630 B.n659 B.n106 163.367
R631 B.n655 B.n106 163.367
R632 B.n655 B.n654 163.367
R633 B.n654 B.n653 163.367
R634 B.n653 B.n108 163.367
R635 B.n649 B.n108 163.367
R636 B.n649 B.n648 163.367
R637 B.n648 B.n647 163.367
R638 B.n647 B.n110 163.367
R639 B.n643 B.n110 163.367
R640 B.n643 B.n642 163.367
R641 B.n642 B.n641 163.367
R642 B.n641 B.n112 163.367
R643 B.n637 B.n112 163.367
R644 B.n637 B.n636 163.367
R645 B.n636 B.n635 163.367
R646 B.n635 B.n114 163.367
R647 B.n631 B.n114 163.367
R648 B.n631 B.n630 163.367
R649 B.n630 B.n629 163.367
R650 B.n629 B.n116 163.367
R651 B.n625 B.n116 163.367
R652 B.n625 B.n624 163.367
R653 B.n624 B.n623 163.367
R654 B.n623 B.n118 163.367
R655 B.n619 B.n118 163.367
R656 B.n619 B.n618 163.367
R657 B.n618 B.n617 163.367
R658 B.n617 B.n120 163.367
R659 B.n613 B.n120 163.367
R660 B.n613 B.n612 163.367
R661 B.n612 B.n611 163.367
R662 B.n611 B.n122 163.367
R663 B.n607 B.n122 163.367
R664 B.n607 B.n606 163.367
R665 B.n606 B.n605 163.367
R666 B.n605 B.n124 163.367
R667 B.n601 B.n124 163.367
R668 B.n601 B.n600 163.367
R669 B.n600 B.n599 163.367
R670 B.n599 B.n126 163.367
R671 B.n595 B.n126 163.367
R672 B.n595 B.n594 163.367
R673 B.n594 B.n593 163.367
R674 B.n593 B.n128 163.367
R675 B.n589 B.n128 163.367
R676 B.n589 B.n588 163.367
R677 B.n588 B.n587 163.367
R678 B.n587 B.n130 163.367
R679 B.n583 B.n130 163.367
R680 B.n583 B.n582 163.367
R681 B.n582 B.n581 163.367
R682 B.n581 B.n132 163.367
R683 B.n577 B.n132 163.367
R684 B.n577 B.n576 163.367
R685 B.n576 B.n575 163.367
R686 B.n575 B.n134 163.367
R687 B.n571 B.n134 163.367
R688 B.n571 B.n570 163.367
R689 B.n570 B.n569 163.367
R690 B.n569 B.n136 163.367
R691 B.n565 B.n136 163.367
R692 B.n565 B.n564 163.367
R693 B.n564 B.n563 163.367
R694 B.n563 B.n138 163.367
R695 B.n559 B.n138 163.367
R696 B.n559 B.n558 163.367
R697 B.n558 B.n557 163.367
R698 B.n557 B.n140 163.367
R699 B.n553 B.n140 163.367
R700 B.n553 B.n552 163.367
R701 B.n552 B.n551 163.367
R702 B.n551 B.n142 163.367
R703 B.n547 B.n142 163.367
R704 B.n547 B.n546 163.367
R705 B.n546 B.n545 163.367
R706 B.n545 B.n144 163.367
R707 B.n541 B.n144 163.367
R708 B.n541 B.n540 163.367
R709 B.n540 B.n539 163.367
R710 B.n539 B.n146 163.367
R711 B.n535 B.n146 163.367
R712 B.n535 B.n534 163.367
R713 B.n534 B.n533 163.367
R714 B.n533 B.n148 163.367
R715 B.n529 B.n148 163.367
R716 B.n529 B.n528 163.367
R717 B.n528 B.n527 163.367
R718 B.n527 B.n150 163.367
R719 B.n523 B.n150 163.367
R720 B.n523 B.n522 163.367
R721 B.n522 B.n521 163.367
R722 B.n521 B.n152 163.367
R723 B.n517 B.n152 163.367
R724 B.n517 B.n516 163.367
R725 B.n516 B.n515 163.367
R726 B.n870 B.n31 163.367
R727 B.n866 B.n31 163.367
R728 B.n866 B.n865 163.367
R729 B.n865 B.n864 163.367
R730 B.n864 B.n33 163.367
R731 B.n860 B.n33 163.367
R732 B.n860 B.n859 163.367
R733 B.n859 B.n858 163.367
R734 B.n858 B.n35 163.367
R735 B.n854 B.n35 163.367
R736 B.n854 B.n853 163.367
R737 B.n853 B.n852 163.367
R738 B.n852 B.n37 163.367
R739 B.n848 B.n37 163.367
R740 B.n848 B.n847 163.367
R741 B.n847 B.n846 163.367
R742 B.n846 B.n39 163.367
R743 B.n842 B.n39 163.367
R744 B.n842 B.n841 163.367
R745 B.n841 B.n840 163.367
R746 B.n840 B.n41 163.367
R747 B.n836 B.n41 163.367
R748 B.n836 B.n835 163.367
R749 B.n835 B.n834 163.367
R750 B.n834 B.n43 163.367
R751 B.n830 B.n43 163.367
R752 B.n830 B.n829 163.367
R753 B.n829 B.n828 163.367
R754 B.n828 B.n45 163.367
R755 B.n824 B.n45 163.367
R756 B.n824 B.n823 163.367
R757 B.n823 B.n822 163.367
R758 B.n822 B.n47 163.367
R759 B.n818 B.n47 163.367
R760 B.n818 B.n817 163.367
R761 B.n817 B.n816 163.367
R762 B.n816 B.n49 163.367
R763 B.n812 B.n49 163.367
R764 B.n812 B.n811 163.367
R765 B.n811 B.n810 163.367
R766 B.n810 B.n51 163.367
R767 B.n806 B.n51 163.367
R768 B.n806 B.n805 163.367
R769 B.n805 B.n804 163.367
R770 B.n804 B.n53 163.367
R771 B.n800 B.n53 163.367
R772 B.n800 B.n799 163.367
R773 B.n799 B.n798 163.367
R774 B.n798 B.n55 163.367
R775 B.n794 B.n55 163.367
R776 B.n794 B.n793 163.367
R777 B.n793 B.n792 163.367
R778 B.n792 B.n57 163.367
R779 B.n788 B.n57 163.367
R780 B.n788 B.n787 163.367
R781 B.n787 B.n786 163.367
R782 B.n786 B.n59 163.367
R783 B.n782 B.n59 163.367
R784 B.n782 B.n781 163.367
R785 B.n781 B.n780 163.367
R786 B.n780 B.n64 163.367
R787 B.n776 B.n64 163.367
R788 B.n776 B.n775 163.367
R789 B.n775 B.n774 163.367
R790 B.n774 B.n66 163.367
R791 B.n769 B.n66 163.367
R792 B.n769 B.n768 163.367
R793 B.n768 B.n767 163.367
R794 B.n767 B.n70 163.367
R795 B.n763 B.n70 163.367
R796 B.n763 B.n762 163.367
R797 B.n762 B.n761 163.367
R798 B.n761 B.n72 163.367
R799 B.n757 B.n72 163.367
R800 B.n757 B.n756 163.367
R801 B.n756 B.n755 163.367
R802 B.n755 B.n74 163.367
R803 B.n751 B.n74 163.367
R804 B.n751 B.n750 163.367
R805 B.n750 B.n749 163.367
R806 B.n749 B.n76 163.367
R807 B.n745 B.n76 163.367
R808 B.n745 B.n744 163.367
R809 B.n744 B.n743 163.367
R810 B.n743 B.n78 163.367
R811 B.n739 B.n78 163.367
R812 B.n739 B.n738 163.367
R813 B.n738 B.n737 163.367
R814 B.n737 B.n80 163.367
R815 B.n733 B.n80 163.367
R816 B.n733 B.n732 163.367
R817 B.n732 B.n731 163.367
R818 B.n731 B.n82 163.367
R819 B.n727 B.n82 163.367
R820 B.n727 B.n726 163.367
R821 B.n726 B.n725 163.367
R822 B.n725 B.n84 163.367
R823 B.n721 B.n84 163.367
R824 B.n721 B.n720 163.367
R825 B.n720 B.n719 163.367
R826 B.n719 B.n86 163.367
R827 B.n715 B.n86 163.367
R828 B.n715 B.n714 163.367
R829 B.n714 B.n713 163.367
R830 B.n713 B.n88 163.367
R831 B.n709 B.n88 163.367
R832 B.n709 B.n708 163.367
R833 B.n708 B.n707 163.367
R834 B.n707 B.n90 163.367
R835 B.n703 B.n90 163.367
R836 B.n703 B.n702 163.367
R837 B.n702 B.n701 163.367
R838 B.n701 B.n92 163.367
R839 B.n697 B.n92 163.367
R840 B.n697 B.n696 163.367
R841 B.n696 B.n695 163.367
R842 B.n695 B.n94 163.367
R843 B.n691 B.n94 163.367
R844 B.n691 B.n690 163.367
R845 B.n690 B.n689 163.367
R846 B.n872 B.n871 163.367
R847 B.n872 B.n29 163.367
R848 B.n876 B.n29 163.367
R849 B.n877 B.n876 163.367
R850 B.n878 B.n877 163.367
R851 B.n878 B.n27 163.367
R852 B.n882 B.n27 163.367
R853 B.n883 B.n882 163.367
R854 B.n884 B.n883 163.367
R855 B.n884 B.n25 163.367
R856 B.n888 B.n25 163.367
R857 B.n889 B.n888 163.367
R858 B.n890 B.n889 163.367
R859 B.n890 B.n23 163.367
R860 B.n894 B.n23 163.367
R861 B.n895 B.n894 163.367
R862 B.n896 B.n895 163.367
R863 B.n896 B.n21 163.367
R864 B.n900 B.n21 163.367
R865 B.n901 B.n900 163.367
R866 B.n902 B.n901 163.367
R867 B.n902 B.n19 163.367
R868 B.n906 B.n19 163.367
R869 B.n907 B.n906 163.367
R870 B.n908 B.n907 163.367
R871 B.n908 B.n17 163.367
R872 B.n912 B.n17 163.367
R873 B.n913 B.n912 163.367
R874 B.n914 B.n913 163.367
R875 B.n914 B.n15 163.367
R876 B.n918 B.n15 163.367
R877 B.n919 B.n918 163.367
R878 B.n920 B.n919 163.367
R879 B.n920 B.n13 163.367
R880 B.n924 B.n13 163.367
R881 B.n925 B.n924 163.367
R882 B.n926 B.n925 163.367
R883 B.n926 B.n11 163.367
R884 B.n930 B.n11 163.367
R885 B.n931 B.n930 163.367
R886 B.n932 B.n931 163.367
R887 B.n932 B.n9 163.367
R888 B.n936 B.n9 163.367
R889 B.n937 B.n936 163.367
R890 B.n938 B.n937 163.367
R891 B.n938 B.n7 163.367
R892 B.n942 B.n7 163.367
R893 B.n943 B.n942 163.367
R894 B.n944 B.n943 163.367
R895 B.n944 B.n5 163.367
R896 B.n948 B.n5 163.367
R897 B.n949 B.n948 163.367
R898 B.n950 B.n949 163.367
R899 B.n950 B.n3 163.367
R900 B.n954 B.n3 163.367
R901 B.n955 B.n954 163.367
R902 B.n246 B.n2 163.367
R903 B.n249 B.n246 163.367
R904 B.n250 B.n249 163.367
R905 B.n251 B.n250 163.367
R906 B.n251 B.n244 163.367
R907 B.n255 B.n244 163.367
R908 B.n256 B.n255 163.367
R909 B.n257 B.n256 163.367
R910 B.n257 B.n242 163.367
R911 B.n261 B.n242 163.367
R912 B.n262 B.n261 163.367
R913 B.n263 B.n262 163.367
R914 B.n263 B.n240 163.367
R915 B.n267 B.n240 163.367
R916 B.n268 B.n267 163.367
R917 B.n269 B.n268 163.367
R918 B.n269 B.n238 163.367
R919 B.n273 B.n238 163.367
R920 B.n274 B.n273 163.367
R921 B.n275 B.n274 163.367
R922 B.n275 B.n236 163.367
R923 B.n279 B.n236 163.367
R924 B.n280 B.n279 163.367
R925 B.n281 B.n280 163.367
R926 B.n281 B.n234 163.367
R927 B.n285 B.n234 163.367
R928 B.n286 B.n285 163.367
R929 B.n287 B.n286 163.367
R930 B.n287 B.n232 163.367
R931 B.n291 B.n232 163.367
R932 B.n292 B.n291 163.367
R933 B.n293 B.n292 163.367
R934 B.n293 B.n230 163.367
R935 B.n297 B.n230 163.367
R936 B.n298 B.n297 163.367
R937 B.n299 B.n298 163.367
R938 B.n299 B.n228 163.367
R939 B.n303 B.n228 163.367
R940 B.n304 B.n303 163.367
R941 B.n305 B.n304 163.367
R942 B.n305 B.n226 163.367
R943 B.n309 B.n226 163.367
R944 B.n310 B.n309 163.367
R945 B.n311 B.n310 163.367
R946 B.n311 B.n224 163.367
R947 B.n315 B.n224 163.367
R948 B.n316 B.n315 163.367
R949 B.n317 B.n316 163.367
R950 B.n317 B.n222 163.367
R951 B.n321 B.n222 163.367
R952 B.n322 B.n321 163.367
R953 B.n323 B.n322 163.367
R954 B.n323 B.n220 163.367
R955 B.n327 B.n220 163.367
R956 B.n328 B.n327 163.367
R957 B.n329 B.n328 163.367
R958 B.n190 B.n189 65.3581
R959 B.n184 B.n183 65.3581
R960 B.n68 B.n67 65.3581
R961 B.n61 B.n60 65.3581
R962 B.n415 B.n190 59.5399
R963 B.n429 B.n184 59.5399
R964 B.n772 B.n68 59.5399
R965 B.n62 B.n61 59.5399
R966 B.n869 B.n30 34.4981
R967 B.n688 B.n687 34.4981
R968 B.n514 B.n513 34.4981
R969 B.n331 B.n330 34.4981
R970 B B.n957 18.0485
R971 B.n873 B.n30 10.6151
R972 B.n874 B.n873 10.6151
R973 B.n875 B.n874 10.6151
R974 B.n875 B.n28 10.6151
R975 B.n879 B.n28 10.6151
R976 B.n880 B.n879 10.6151
R977 B.n881 B.n880 10.6151
R978 B.n881 B.n26 10.6151
R979 B.n885 B.n26 10.6151
R980 B.n886 B.n885 10.6151
R981 B.n887 B.n886 10.6151
R982 B.n887 B.n24 10.6151
R983 B.n891 B.n24 10.6151
R984 B.n892 B.n891 10.6151
R985 B.n893 B.n892 10.6151
R986 B.n893 B.n22 10.6151
R987 B.n897 B.n22 10.6151
R988 B.n898 B.n897 10.6151
R989 B.n899 B.n898 10.6151
R990 B.n899 B.n20 10.6151
R991 B.n903 B.n20 10.6151
R992 B.n904 B.n903 10.6151
R993 B.n905 B.n904 10.6151
R994 B.n905 B.n18 10.6151
R995 B.n909 B.n18 10.6151
R996 B.n910 B.n909 10.6151
R997 B.n911 B.n910 10.6151
R998 B.n911 B.n16 10.6151
R999 B.n915 B.n16 10.6151
R1000 B.n916 B.n915 10.6151
R1001 B.n917 B.n916 10.6151
R1002 B.n917 B.n14 10.6151
R1003 B.n921 B.n14 10.6151
R1004 B.n922 B.n921 10.6151
R1005 B.n923 B.n922 10.6151
R1006 B.n923 B.n12 10.6151
R1007 B.n927 B.n12 10.6151
R1008 B.n928 B.n927 10.6151
R1009 B.n929 B.n928 10.6151
R1010 B.n929 B.n10 10.6151
R1011 B.n933 B.n10 10.6151
R1012 B.n934 B.n933 10.6151
R1013 B.n935 B.n934 10.6151
R1014 B.n935 B.n8 10.6151
R1015 B.n939 B.n8 10.6151
R1016 B.n940 B.n939 10.6151
R1017 B.n941 B.n940 10.6151
R1018 B.n941 B.n6 10.6151
R1019 B.n945 B.n6 10.6151
R1020 B.n946 B.n945 10.6151
R1021 B.n947 B.n946 10.6151
R1022 B.n947 B.n4 10.6151
R1023 B.n951 B.n4 10.6151
R1024 B.n952 B.n951 10.6151
R1025 B.n953 B.n952 10.6151
R1026 B.n953 B.n0 10.6151
R1027 B.n869 B.n868 10.6151
R1028 B.n868 B.n867 10.6151
R1029 B.n867 B.n32 10.6151
R1030 B.n863 B.n32 10.6151
R1031 B.n863 B.n862 10.6151
R1032 B.n862 B.n861 10.6151
R1033 B.n861 B.n34 10.6151
R1034 B.n857 B.n34 10.6151
R1035 B.n857 B.n856 10.6151
R1036 B.n856 B.n855 10.6151
R1037 B.n855 B.n36 10.6151
R1038 B.n851 B.n36 10.6151
R1039 B.n851 B.n850 10.6151
R1040 B.n850 B.n849 10.6151
R1041 B.n849 B.n38 10.6151
R1042 B.n845 B.n38 10.6151
R1043 B.n845 B.n844 10.6151
R1044 B.n844 B.n843 10.6151
R1045 B.n843 B.n40 10.6151
R1046 B.n839 B.n40 10.6151
R1047 B.n839 B.n838 10.6151
R1048 B.n838 B.n837 10.6151
R1049 B.n837 B.n42 10.6151
R1050 B.n833 B.n42 10.6151
R1051 B.n833 B.n832 10.6151
R1052 B.n832 B.n831 10.6151
R1053 B.n831 B.n44 10.6151
R1054 B.n827 B.n44 10.6151
R1055 B.n827 B.n826 10.6151
R1056 B.n826 B.n825 10.6151
R1057 B.n825 B.n46 10.6151
R1058 B.n821 B.n46 10.6151
R1059 B.n821 B.n820 10.6151
R1060 B.n820 B.n819 10.6151
R1061 B.n819 B.n48 10.6151
R1062 B.n815 B.n48 10.6151
R1063 B.n815 B.n814 10.6151
R1064 B.n814 B.n813 10.6151
R1065 B.n813 B.n50 10.6151
R1066 B.n809 B.n50 10.6151
R1067 B.n809 B.n808 10.6151
R1068 B.n808 B.n807 10.6151
R1069 B.n807 B.n52 10.6151
R1070 B.n803 B.n52 10.6151
R1071 B.n803 B.n802 10.6151
R1072 B.n802 B.n801 10.6151
R1073 B.n801 B.n54 10.6151
R1074 B.n797 B.n54 10.6151
R1075 B.n797 B.n796 10.6151
R1076 B.n796 B.n795 10.6151
R1077 B.n795 B.n56 10.6151
R1078 B.n791 B.n56 10.6151
R1079 B.n791 B.n790 10.6151
R1080 B.n790 B.n789 10.6151
R1081 B.n789 B.n58 10.6151
R1082 B.n785 B.n784 10.6151
R1083 B.n784 B.n783 10.6151
R1084 B.n783 B.n63 10.6151
R1085 B.n779 B.n63 10.6151
R1086 B.n779 B.n778 10.6151
R1087 B.n778 B.n777 10.6151
R1088 B.n777 B.n65 10.6151
R1089 B.n773 B.n65 10.6151
R1090 B.n771 B.n770 10.6151
R1091 B.n770 B.n69 10.6151
R1092 B.n766 B.n69 10.6151
R1093 B.n766 B.n765 10.6151
R1094 B.n765 B.n764 10.6151
R1095 B.n764 B.n71 10.6151
R1096 B.n760 B.n71 10.6151
R1097 B.n760 B.n759 10.6151
R1098 B.n759 B.n758 10.6151
R1099 B.n758 B.n73 10.6151
R1100 B.n754 B.n73 10.6151
R1101 B.n754 B.n753 10.6151
R1102 B.n753 B.n752 10.6151
R1103 B.n752 B.n75 10.6151
R1104 B.n748 B.n75 10.6151
R1105 B.n748 B.n747 10.6151
R1106 B.n747 B.n746 10.6151
R1107 B.n746 B.n77 10.6151
R1108 B.n742 B.n77 10.6151
R1109 B.n742 B.n741 10.6151
R1110 B.n741 B.n740 10.6151
R1111 B.n740 B.n79 10.6151
R1112 B.n736 B.n79 10.6151
R1113 B.n736 B.n735 10.6151
R1114 B.n735 B.n734 10.6151
R1115 B.n734 B.n81 10.6151
R1116 B.n730 B.n81 10.6151
R1117 B.n730 B.n729 10.6151
R1118 B.n729 B.n728 10.6151
R1119 B.n728 B.n83 10.6151
R1120 B.n724 B.n83 10.6151
R1121 B.n724 B.n723 10.6151
R1122 B.n723 B.n722 10.6151
R1123 B.n722 B.n85 10.6151
R1124 B.n718 B.n85 10.6151
R1125 B.n718 B.n717 10.6151
R1126 B.n717 B.n716 10.6151
R1127 B.n716 B.n87 10.6151
R1128 B.n712 B.n87 10.6151
R1129 B.n712 B.n711 10.6151
R1130 B.n711 B.n710 10.6151
R1131 B.n710 B.n89 10.6151
R1132 B.n706 B.n89 10.6151
R1133 B.n706 B.n705 10.6151
R1134 B.n705 B.n704 10.6151
R1135 B.n704 B.n91 10.6151
R1136 B.n700 B.n91 10.6151
R1137 B.n700 B.n699 10.6151
R1138 B.n699 B.n698 10.6151
R1139 B.n698 B.n93 10.6151
R1140 B.n694 B.n93 10.6151
R1141 B.n694 B.n693 10.6151
R1142 B.n693 B.n692 10.6151
R1143 B.n692 B.n95 10.6151
R1144 B.n688 B.n95 10.6151
R1145 B.n687 B.n686 10.6151
R1146 B.n686 B.n97 10.6151
R1147 B.n682 B.n97 10.6151
R1148 B.n682 B.n681 10.6151
R1149 B.n681 B.n680 10.6151
R1150 B.n680 B.n99 10.6151
R1151 B.n676 B.n99 10.6151
R1152 B.n676 B.n675 10.6151
R1153 B.n675 B.n674 10.6151
R1154 B.n674 B.n101 10.6151
R1155 B.n670 B.n101 10.6151
R1156 B.n670 B.n669 10.6151
R1157 B.n669 B.n668 10.6151
R1158 B.n668 B.n103 10.6151
R1159 B.n664 B.n103 10.6151
R1160 B.n664 B.n663 10.6151
R1161 B.n663 B.n662 10.6151
R1162 B.n662 B.n105 10.6151
R1163 B.n658 B.n105 10.6151
R1164 B.n658 B.n657 10.6151
R1165 B.n657 B.n656 10.6151
R1166 B.n656 B.n107 10.6151
R1167 B.n652 B.n107 10.6151
R1168 B.n652 B.n651 10.6151
R1169 B.n651 B.n650 10.6151
R1170 B.n650 B.n109 10.6151
R1171 B.n646 B.n109 10.6151
R1172 B.n646 B.n645 10.6151
R1173 B.n645 B.n644 10.6151
R1174 B.n644 B.n111 10.6151
R1175 B.n640 B.n111 10.6151
R1176 B.n640 B.n639 10.6151
R1177 B.n639 B.n638 10.6151
R1178 B.n638 B.n113 10.6151
R1179 B.n634 B.n113 10.6151
R1180 B.n634 B.n633 10.6151
R1181 B.n633 B.n632 10.6151
R1182 B.n632 B.n115 10.6151
R1183 B.n628 B.n115 10.6151
R1184 B.n628 B.n627 10.6151
R1185 B.n627 B.n626 10.6151
R1186 B.n626 B.n117 10.6151
R1187 B.n622 B.n117 10.6151
R1188 B.n622 B.n621 10.6151
R1189 B.n621 B.n620 10.6151
R1190 B.n620 B.n119 10.6151
R1191 B.n616 B.n119 10.6151
R1192 B.n616 B.n615 10.6151
R1193 B.n615 B.n614 10.6151
R1194 B.n614 B.n121 10.6151
R1195 B.n610 B.n121 10.6151
R1196 B.n610 B.n609 10.6151
R1197 B.n609 B.n608 10.6151
R1198 B.n608 B.n123 10.6151
R1199 B.n604 B.n123 10.6151
R1200 B.n604 B.n603 10.6151
R1201 B.n603 B.n602 10.6151
R1202 B.n602 B.n125 10.6151
R1203 B.n598 B.n125 10.6151
R1204 B.n598 B.n597 10.6151
R1205 B.n597 B.n596 10.6151
R1206 B.n596 B.n127 10.6151
R1207 B.n592 B.n127 10.6151
R1208 B.n592 B.n591 10.6151
R1209 B.n591 B.n590 10.6151
R1210 B.n590 B.n129 10.6151
R1211 B.n586 B.n129 10.6151
R1212 B.n586 B.n585 10.6151
R1213 B.n585 B.n584 10.6151
R1214 B.n584 B.n131 10.6151
R1215 B.n580 B.n131 10.6151
R1216 B.n580 B.n579 10.6151
R1217 B.n579 B.n578 10.6151
R1218 B.n578 B.n133 10.6151
R1219 B.n574 B.n133 10.6151
R1220 B.n574 B.n573 10.6151
R1221 B.n573 B.n572 10.6151
R1222 B.n572 B.n135 10.6151
R1223 B.n568 B.n135 10.6151
R1224 B.n568 B.n567 10.6151
R1225 B.n567 B.n566 10.6151
R1226 B.n566 B.n137 10.6151
R1227 B.n562 B.n137 10.6151
R1228 B.n562 B.n561 10.6151
R1229 B.n561 B.n560 10.6151
R1230 B.n560 B.n139 10.6151
R1231 B.n556 B.n139 10.6151
R1232 B.n556 B.n555 10.6151
R1233 B.n555 B.n554 10.6151
R1234 B.n554 B.n141 10.6151
R1235 B.n550 B.n141 10.6151
R1236 B.n550 B.n549 10.6151
R1237 B.n549 B.n548 10.6151
R1238 B.n548 B.n143 10.6151
R1239 B.n544 B.n143 10.6151
R1240 B.n544 B.n543 10.6151
R1241 B.n543 B.n542 10.6151
R1242 B.n542 B.n145 10.6151
R1243 B.n538 B.n145 10.6151
R1244 B.n538 B.n537 10.6151
R1245 B.n537 B.n536 10.6151
R1246 B.n536 B.n147 10.6151
R1247 B.n532 B.n147 10.6151
R1248 B.n532 B.n531 10.6151
R1249 B.n531 B.n530 10.6151
R1250 B.n530 B.n149 10.6151
R1251 B.n526 B.n149 10.6151
R1252 B.n526 B.n525 10.6151
R1253 B.n525 B.n524 10.6151
R1254 B.n524 B.n151 10.6151
R1255 B.n520 B.n151 10.6151
R1256 B.n520 B.n519 10.6151
R1257 B.n519 B.n518 10.6151
R1258 B.n518 B.n153 10.6151
R1259 B.n514 B.n153 10.6151
R1260 B.n247 B.n1 10.6151
R1261 B.n248 B.n247 10.6151
R1262 B.n248 B.n245 10.6151
R1263 B.n252 B.n245 10.6151
R1264 B.n253 B.n252 10.6151
R1265 B.n254 B.n253 10.6151
R1266 B.n254 B.n243 10.6151
R1267 B.n258 B.n243 10.6151
R1268 B.n259 B.n258 10.6151
R1269 B.n260 B.n259 10.6151
R1270 B.n260 B.n241 10.6151
R1271 B.n264 B.n241 10.6151
R1272 B.n265 B.n264 10.6151
R1273 B.n266 B.n265 10.6151
R1274 B.n266 B.n239 10.6151
R1275 B.n270 B.n239 10.6151
R1276 B.n271 B.n270 10.6151
R1277 B.n272 B.n271 10.6151
R1278 B.n272 B.n237 10.6151
R1279 B.n276 B.n237 10.6151
R1280 B.n277 B.n276 10.6151
R1281 B.n278 B.n277 10.6151
R1282 B.n278 B.n235 10.6151
R1283 B.n282 B.n235 10.6151
R1284 B.n283 B.n282 10.6151
R1285 B.n284 B.n283 10.6151
R1286 B.n284 B.n233 10.6151
R1287 B.n288 B.n233 10.6151
R1288 B.n289 B.n288 10.6151
R1289 B.n290 B.n289 10.6151
R1290 B.n290 B.n231 10.6151
R1291 B.n294 B.n231 10.6151
R1292 B.n295 B.n294 10.6151
R1293 B.n296 B.n295 10.6151
R1294 B.n296 B.n229 10.6151
R1295 B.n300 B.n229 10.6151
R1296 B.n301 B.n300 10.6151
R1297 B.n302 B.n301 10.6151
R1298 B.n302 B.n227 10.6151
R1299 B.n306 B.n227 10.6151
R1300 B.n307 B.n306 10.6151
R1301 B.n308 B.n307 10.6151
R1302 B.n308 B.n225 10.6151
R1303 B.n312 B.n225 10.6151
R1304 B.n313 B.n312 10.6151
R1305 B.n314 B.n313 10.6151
R1306 B.n314 B.n223 10.6151
R1307 B.n318 B.n223 10.6151
R1308 B.n319 B.n318 10.6151
R1309 B.n320 B.n319 10.6151
R1310 B.n320 B.n221 10.6151
R1311 B.n324 B.n221 10.6151
R1312 B.n325 B.n324 10.6151
R1313 B.n326 B.n325 10.6151
R1314 B.n326 B.n219 10.6151
R1315 B.n330 B.n219 10.6151
R1316 B.n332 B.n331 10.6151
R1317 B.n332 B.n217 10.6151
R1318 B.n336 B.n217 10.6151
R1319 B.n337 B.n336 10.6151
R1320 B.n338 B.n337 10.6151
R1321 B.n338 B.n215 10.6151
R1322 B.n342 B.n215 10.6151
R1323 B.n343 B.n342 10.6151
R1324 B.n344 B.n343 10.6151
R1325 B.n344 B.n213 10.6151
R1326 B.n348 B.n213 10.6151
R1327 B.n349 B.n348 10.6151
R1328 B.n350 B.n349 10.6151
R1329 B.n350 B.n211 10.6151
R1330 B.n354 B.n211 10.6151
R1331 B.n355 B.n354 10.6151
R1332 B.n356 B.n355 10.6151
R1333 B.n356 B.n209 10.6151
R1334 B.n360 B.n209 10.6151
R1335 B.n361 B.n360 10.6151
R1336 B.n362 B.n361 10.6151
R1337 B.n362 B.n207 10.6151
R1338 B.n366 B.n207 10.6151
R1339 B.n367 B.n366 10.6151
R1340 B.n368 B.n367 10.6151
R1341 B.n368 B.n205 10.6151
R1342 B.n372 B.n205 10.6151
R1343 B.n373 B.n372 10.6151
R1344 B.n374 B.n373 10.6151
R1345 B.n374 B.n203 10.6151
R1346 B.n378 B.n203 10.6151
R1347 B.n379 B.n378 10.6151
R1348 B.n380 B.n379 10.6151
R1349 B.n380 B.n201 10.6151
R1350 B.n384 B.n201 10.6151
R1351 B.n385 B.n384 10.6151
R1352 B.n386 B.n385 10.6151
R1353 B.n386 B.n199 10.6151
R1354 B.n390 B.n199 10.6151
R1355 B.n391 B.n390 10.6151
R1356 B.n392 B.n391 10.6151
R1357 B.n392 B.n197 10.6151
R1358 B.n396 B.n197 10.6151
R1359 B.n397 B.n396 10.6151
R1360 B.n398 B.n397 10.6151
R1361 B.n398 B.n195 10.6151
R1362 B.n402 B.n195 10.6151
R1363 B.n403 B.n402 10.6151
R1364 B.n404 B.n403 10.6151
R1365 B.n404 B.n193 10.6151
R1366 B.n408 B.n193 10.6151
R1367 B.n409 B.n408 10.6151
R1368 B.n410 B.n409 10.6151
R1369 B.n410 B.n191 10.6151
R1370 B.n414 B.n191 10.6151
R1371 B.n417 B.n416 10.6151
R1372 B.n417 B.n187 10.6151
R1373 B.n421 B.n187 10.6151
R1374 B.n422 B.n421 10.6151
R1375 B.n423 B.n422 10.6151
R1376 B.n423 B.n185 10.6151
R1377 B.n427 B.n185 10.6151
R1378 B.n428 B.n427 10.6151
R1379 B.n430 B.n181 10.6151
R1380 B.n434 B.n181 10.6151
R1381 B.n435 B.n434 10.6151
R1382 B.n436 B.n435 10.6151
R1383 B.n436 B.n179 10.6151
R1384 B.n440 B.n179 10.6151
R1385 B.n441 B.n440 10.6151
R1386 B.n442 B.n441 10.6151
R1387 B.n442 B.n177 10.6151
R1388 B.n446 B.n177 10.6151
R1389 B.n447 B.n446 10.6151
R1390 B.n448 B.n447 10.6151
R1391 B.n448 B.n175 10.6151
R1392 B.n452 B.n175 10.6151
R1393 B.n453 B.n452 10.6151
R1394 B.n454 B.n453 10.6151
R1395 B.n454 B.n173 10.6151
R1396 B.n458 B.n173 10.6151
R1397 B.n459 B.n458 10.6151
R1398 B.n460 B.n459 10.6151
R1399 B.n460 B.n171 10.6151
R1400 B.n464 B.n171 10.6151
R1401 B.n465 B.n464 10.6151
R1402 B.n466 B.n465 10.6151
R1403 B.n466 B.n169 10.6151
R1404 B.n470 B.n169 10.6151
R1405 B.n471 B.n470 10.6151
R1406 B.n472 B.n471 10.6151
R1407 B.n472 B.n167 10.6151
R1408 B.n476 B.n167 10.6151
R1409 B.n477 B.n476 10.6151
R1410 B.n478 B.n477 10.6151
R1411 B.n478 B.n165 10.6151
R1412 B.n482 B.n165 10.6151
R1413 B.n483 B.n482 10.6151
R1414 B.n484 B.n483 10.6151
R1415 B.n484 B.n163 10.6151
R1416 B.n488 B.n163 10.6151
R1417 B.n489 B.n488 10.6151
R1418 B.n490 B.n489 10.6151
R1419 B.n490 B.n161 10.6151
R1420 B.n494 B.n161 10.6151
R1421 B.n495 B.n494 10.6151
R1422 B.n496 B.n495 10.6151
R1423 B.n496 B.n159 10.6151
R1424 B.n500 B.n159 10.6151
R1425 B.n501 B.n500 10.6151
R1426 B.n502 B.n501 10.6151
R1427 B.n502 B.n157 10.6151
R1428 B.n506 B.n157 10.6151
R1429 B.n507 B.n506 10.6151
R1430 B.n508 B.n507 10.6151
R1431 B.n508 B.n155 10.6151
R1432 B.n512 B.n155 10.6151
R1433 B.n513 B.n512 10.6151
R1434 B.n957 B.n0 8.11757
R1435 B.n957 B.n1 8.11757
R1436 B.n785 B.n62 6.5566
R1437 B.n773 B.n772 6.5566
R1438 B.n416 B.n415 6.5566
R1439 B.n429 B.n428 6.5566
R1440 B.n62 B.n58 4.05904
R1441 B.n772 B.n771 4.05904
R1442 B.n415 B.n414 4.05904
R1443 B.n430 B.n429 4.05904
R1444 VP.n19 VP.t7 166.341
R1445 VP.n21 VP.n18 161.3
R1446 VP.n23 VP.n22 161.3
R1447 VP.n24 VP.n17 161.3
R1448 VP.n26 VP.n25 161.3
R1449 VP.n27 VP.n16 161.3
R1450 VP.n29 VP.n28 161.3
R1451 VP.n31 VP.n30 161.3
R1452 VP.n32 VP.n14 161.3
R1453 VP.n34 VP.n33 161.3
R1454 VP.n35 VP.n13 161.3
R1455 VP.n37 VP.n36 161.3
R1456 VP.n38 VP.n12 161.3
R1457 VP.n40 VP.n39 161.3
R1458 VP.n75 VP.n74 161.3
R1459 VP.n73 VP.n1 161.3
R1460 VP.n72 VP.n71 161.3
R1461 VP.n70 VP.n2 161.3
R1462 VP.n69 VP.n68 161.3
R1463 VP.n67 VP.n3 161.3
R1464 VP.n66 VP.n65 161.3
R1465 VP.n64 VP.n63 161.3
R1466 VP.n62 VP.n5 161.3
R1467 VP.n61 VP.n60 161.3
R1468 VP.n59 VP.n6 161.3
R1469 VP.n58 VP.n57 161.3
R1470 VP.n56 VP.n7 161.3
R1471 VP.n54 VP.n53 161.3
R1472 VP.n52 VP.n8 161.3
R1473 VP.n51 VP.n50 161.3
R1474 VP.n49 VP.n9 161.3
R1475 VP.n48 VP.n47 161.3
R1476 VP.n46 VP.n10 161.3
R1477 VP.n45 VP.n44 161.3
R1478 VP.n43 VP.t3 133.185
R1479 VP.n55 VP.t6 133.185
R1480 VP.n4 VP.t4 133.185
R1481 VP.n0 VP.t5 133.185
R1482 VP.n11 VP.t2 133.185
R1483 VP.n15 VP.t0 133.185
R1484 VP.n20 VP.t1 133.185
R1485 VP.n43 VP.n42 75.2445
R1486 VP.n76 VP.n0 75.2445
R1487 VP.n41 VP.n11 75.2445
R1488 VP.n42 VP.n41 56.6435
R1489 VP.n61 VP.n6 56.5617
R1490 VP.n26 VP.n17 56.5617
R1491 VP.n20 VP.n19 52.6903
R1492 VP.n49 VP.n48 52.2023
R1493 VP.n72 VP.n2 52.2023
R1494 VP.n37 VP.n13 52.2023
R1495 VP.n50 VP.n49 28.9518
R1496 VP.n68 VP.n2 28.9518
R1497 VP.n33 VP.n13 28.9518
R1498 VP.n44 VP.n10 24.5923
R1499 VP.n48 VP.n10 24.5923
R1500 VP.n50 VP.n8 24.5923
R1501 VP.n54 VP.n8 24.5923
R1502 VP.n57 VP.n56 24.5923
R1503 VP.n57 VP.n6 24.5923
R1504 VP.n62 VP.n61 24.5923
R1505 VP.n63 VP.n62 24.5923
R1506 VP.n67 VP.n66 24.5923
R1507 VP.n68 VP.n67 24.5923
R1508 VP.n73 VP.n72 24.5923
R1509 VP.n74 VP.n73 24.5923
R1510 VP.n38 VP.n37 24.5923
R1511 VP.n39 VP.n38 24.5923
R1512 VP.n27 VP.n26 24.5923
R1513 VP.n28 VP.n27 24.5923
R1514 VP.n32 VP.n31 24.5923
R1515 VP.n33 VP.n32 24.5923
R1516 VP.n22 VP.n21 24.5923
R1517 VP.n22 VP.n17 24.5923
R1518 VP.n56 VP.n55 21.3954
R1519 VP.n63 VP.n4 21.3954
R1520 VP.n28 VP.n15 21.3954
R1521 VP.n21 VP.n20 21.3954
R1522 VP.n44 VP.n43 15.0015
R1523 VP.n74 VP.n0 15.0015
R1524 VP.n39 VP.n11 15.0015
R1525 VP.n19 VP.n18 4.13669
R1526 VP.n55 VP.n54 3.19744
R1527 VP.n66 VP.n4 3.19744
R1528 VP.n31 VP.n15 3.19744
R1529 VP.n41 VP.n40 0.354861
R1530 VP.n45 VP.n42 0.354861
R1531 VP.n76 VP.n75 0.354861
R1532 VP VP.n76 0.267071
R1533 VP.n23 VP.n18 0.189894
R1534 VP.n24 VP.n23 0.189894
R1535 VP.n25 VP.n24 0.189894
R1536 VP.n25 VP.n16 0.189894
R1537 VP.n29 VP.n16 0.189894
R1538 VP.n30 VP.n29 0.189894
R1539 VP.n30 VP.n14 0.189894
R1540 VP.n34 VP.n14 0.189894
R1541 VP.n35 VP.n34 0.189894
R1542 VP.n36 VP.n35 0.189894
R1543 VP.n36 VP.n12 0.189894
R1544 VP.n40 VP.n12 0.189894
R1545 VP.n46 VP.n45 0.189894
R1546 VP.n47 VP.n46 0.189894
R1547 VP.n47 VP.n9 0.189894
R1548 VP.n51 VP.n9 0.189894
R1549 VP.n52 VP.n51 0.189894
R1550 VP.n53 VP.n52 0.189894
R1551 VP.n53 VP.n7 0.189894
R1552 VP.n58 VP.n7 0.189894
R1553 VP.n59 VP.n58 0.189894
R1554 VP.n60 VP.n59 0.189894
R1555 VP.n60 VP.n5 0.189894
R1556 VP.n64 VP.n5 0.189894
R1557 VP.n65 VP.n64 0.189894
R1558 VP.n65 VP.n3 0.189894
R1559 VP.n69 VP.n3 0.189894
R1560 VP.n70 VP.n69 0.189894
R1561 VP.n71 VP.n70 0.189894
R1562 VP.n71 VP.n1 0.189894
R1563 VP.n75 VP.n1 0.189894
R1564 VDD1 VDD1.n0 70.9028
R1565 VDD1.n3 VDD1.n2 70.7891
R1566 VDD1.n3 VDD1.n1 70.7891
R1567 VDD1.n5 VDD1.n4 69.3918
R1568 VDD1.n5 VDD1.n3 51.8543
R1569 VDD1.n4 VDD1.t6 1.93532
R1570 VDD1.n4 VDD1.t1 1.93532
R1571 VDD1.n0 VDD1.t7 1.93532
R1572 VDD1.n0 VDD1.t4 1.93532
R1573 VDD1.n2 VDD1.t2 1.93532
R1574 VDD1.n2 VDD1.t3 1.93532
R1575 VDD1.n1 VDD1.t0 1.93532
R1576 VDD1.n1 VDD1.t5 1.93532
R1577 VDD1 VDD1.n5 1.3949
R1578 VTAIL.n754 VTAIL.n666 756.745
R1579 VTAIL.n90 VTAIL.n2 756.745
R1580 VTAIL.n184 VTAIL.n96 756.745
R1581 VTAIL.n280 VTAIL.n192 756.745
R1582 VTAIL.n660 VTAIL.n572 756.745
R1583 VTAIL.n564 VTAIL.n476 756.745
R1584 VTAIL.n470 VTAIL.n382 756.745
R1585 VTAIL.n374 VTAIL.n286 756.745
R1586 VTAIL.n697 VTAIL.n696 585
R1587 VTAIL.n694 VTAIL.n693 585
R1588 VTAIL.n703 VTAIL.n702 585
R1589 VTAIL.n705 VTAIL.n704 585
R1590 VTAIL.n690 VTAIL.n689 585
R1591 VTAIL.n711 VTAIL.n710 585
R1592 VTAIL.n713 VTAIL.n712 585
R1593 VTAIL.n686 VTAIL.n685 585
R1594 VTAIL.n719 VTAIL.n718 585
R1595 VTAIL.n721 VTAIL.n720 585
R1596 VTAIL.n682 VTAIL.n681 585
R1597 VTAIL.n727 VTAIL.n726 585
R1598 VTAIL.n729 VTAIL.n728 585
R1599 VTAIL.n678 VTAIL.n677 585
R1600 VTAIL.n735 VTAIL.n734 585
R1601 VTAIL.n738 VTAIL.n737 585
R1602 VTAIL.n736 VTAIL.n674 585
R1603 VTAIL.n743 VTAIL.n673 585
R1604 VTAIL.n745 VTAIL.n744 585
R1605 VTAIL.n747 VTAIL.n746 585
R1606 VTAIL.n670 VTAIL.n669 585
R1607 VTAIL.n753 VTAIL.n752 585
R1608 VTAIL.n755 VTAIL.n754 585
R1609 VTAIL.n33 VTAIL.n32 585
R1610 VTAIL.n30 VTAIL.n29 585
R1611 VTAIL.n39 VTAIL.n38 585
R1612 VTAIL.n41 VTAIL.n40 585
R1613 VTAIL.n26 VTAIL.n25 585
R1614 VTAIL.n47 VTAIL.n46 585
R1615 VTAIL.n49 VTAIL.n48 585
R1616 VTAIL.n22 VTAIL.n21 585
R1617 VTAIL.n55 VTAIL.n54 585
R1618 VTAIL.n57 VTAIL.n56 585
R1619 VTAIL.n18 VTAIL.n17 585
R1620 VTAIL.n63 VTAIL.n62 585
R1621 VTAIL.n65 VTAIL.n64 585
R1622 VTAIL.n14 VTAIL.n13 585
R1623 VTAIL.n71 VTAIL.n70 585
R1624 VTAIL.n74 VTAIL.n73 585
R1625 VTAIL.n72 VTAIL.n10 585
R1626 VTAIL.n79 VTAIL.n9 585
R1627 VTAIL.n81 VTAIL.n80 585
R1628 VTAIL.n83 VTAIL.n82 585
R1629 VTAIL.n6 VTAIL.n5 585
R1630 VTAIL.n89 VTAIL.n88 585
R1631 VTAIL.n91 VTAIL.n90 585
R1632 VTAIL.n127 VTAIL.n126 585
R1633 VTAIL.n124 VTAIL.n123 585
R1634 VTAIL.n133 VTAIL.n132 585
R1635 VTAIL.n135 VTAIL.n134 585
R1636 VTAIL.n120 VTAIL.n119 585
R1637 VTAIL.n141 VTAIL.n140 585
R1638 VTAIL.n143 VTAIL.n142 585
R1639 VTAIL.n116 VTAIL.n115 585
R1640 VTAIL.n149 VTAIL.n148 585
R1641 VTAIL.n151 VTAIL.n150 585
R1642 VTAIL.n112 VTAIL.n111 585
R1643 VTAIL.n157 VTAIL.n156 585
R1644 VTAIL.n159 VTAIL.n158 585
R1645 VTAIL.n108 VTAIL.n107 585
R1646 VTAIL.n165 VTAIL.n164 585
R1647 VTAIL.n168 VTAIL.n167 585
R1648 VTAIL.n166 VTAIL.n104 585
R1649 VTAIL.n173 VTAIL.n103 585
R1650 VTAIL.n175 VTAIL.n174 585
R1651 VTAIL.n177 VTAIL.n176 585
R1652 VTAIL.n100 VTAIL.n99 585
R1653 VTAIL.n183 VTAIL.n182 585
R1654 VTAIL.n185 VTAIL.n184 585
R1655 VTAIL.n223 VTAIL.n222 585
R1656 VTAIL.n220 VTAIL.n219 585
R1657 VTAIL.n229 VTAIL.n228 585
R1658 VTAIL.n231 VTAIL.n230 585
R1659 VTAIL.n216 VTAIL.n215 585
R1660 VTAIL.n237 VTAIL.n236 585
R1661 VTAIL.n239 VTAIL.n238 585
R1662 VTAIL.n212 VTAIL.n211 585
R1663 VTAIL.n245 VTAIL.n244 585
R1664 VTAIL.n247 VTAIL.n246 585
R1665 VTAIL.n208 VTAIL.n207 585
R1666 VTAIL.n253 VTAIL.n252 585
R1667 VTAIL.n255 VTAIL.n254 585
R1668 VTAIL.n204 VTAIL.n203 585
R1669 VTAIL.n261 VTAIL.n260 585
R1670 VTAIL.n264 VTAIL.n263 585
R1671 VTAIL.n262 VTAIL.n200 585
R1672 VTAIL.n269 VTAIL.n199 585
R1673 VTAIL.n271 VTAIL.n270 585
R1674 VTAIL.n273 VTAIL.n272 585
R1675 VTAIL.n196 VTAIL.n195 585
R1676 VTAIL.n279 VTAIL.n278 585
R1677 VTAIL.n281 VTAIL.n280 585
R1678 VTAIL.n661 VTAIL.n660 585
R1679 VTAIL.n659 VTAIL.n658 585
R1680 VTAIL.n576 VTAIL.n575 585
R1681 VTAIL.n653 VTAIL.n652 585
R1682 VTAIL.n651 VTAIL.n650 585
R1683 VTAIL.n649 VTAIL.n579 585
R1684 VTAIL.n583 VTAIL.n580 585
R1685 VTAIL.n644 VTAIL.n643 585
R1686 VTAIL.n642 VTAIL.n641 585
R1687 VTAIL.n585 VTAIL.n584 585
R1688 VTAIL.n636 VTAIL.n635 585
R1689 VTAIL.n634 VTAIL.n633 585
R1690 VTAIL.n589 VTAIL.n588 585
R1691 VTAIL.n628 VTAIL.n627 585
R1692 VTAIL.n626 VTAIL.n625 585
R1693 VTAIL.n593 VTAIL.n592 585
R1694 VTAIL.n620 VTAIL.n619 585
R1695 VTAIL.n618 VTAIL.n617 585
R1696 VTAIL.n597 VTAIL.n596 585
R1697 VTAIL.n612 VTAIL.n611 585
R1698 VTAIL.n610 VTAIL.n609 585
R1699 VTAIL.n601 VTAIL.n600 585
R1700 VTAIL.n604 VTAIL.n603 585
R1701 VTAIL.n565 VTAIL.n564 585
R1702 VTAIL.n563 VTAIL.n562 585
R1703 VTAIL.n480 VTAIL.n479 585
R1704 VTAIL.n557 VTAIL.n556 585
R1705 VTAIL.n555 VTAIL.n554 585
R1706 VTAIL.n553 VTAIL.n483 585
R1707 VTAIL.n487 VTAIL.n484 585
R1708 VTAIL.n548 VTAIL.n547 585
R1709 VTAIL.n546 VTAIL.n545 585
R1710 VTAIL.n489 VTAIL.n488 585
R1711 VTAIL.n540 VTAIL.n539 585
R1712 VTAIL.n538 VTAIL.n537 585
R1713 VTAIL.n493 VTAIL.n492 585
R1714 VTAIL.n532 VTAIL.n531 585
R1715 VTAIL.n530 VTAIL.n529 585
R1716 VTAIL.n497 VTAIL.n496 585
R1717 VTAIL.n524 VTAIL.n523 585
R1718 VTAIL.n522 VTAIL.n521 585
R1719 VTAIL.n501 VTAIL.n500 585
R1720 VTAIL.n516 VTAIL.n515 585
R1721 VTAIL.n514 VTAIL.n513 585
R1722 VTAIL.n505 VTAIL.n504 585
R1723 VTAIL.n508 VTAIL.n507 585
R1724 VTAIL.n471 VTAIL.n470 585
R1725 VTAIL.n469 VTAIL.n468 585
R1726 VTAIL.n386 VTAIL.n385 585
R1727 VTAIL.n463 VTAIL.n462 585
R1728 VTAIL.n461 VTAIL.n460 585
R1729 VTAIL.n459 VTAIL.n389 585
R1730 VTAIL.n393 VTAIL.n390 585
R1731 VTAIL.n454 VTAIL.n453 585
R1732 VTAIL.n452 VTAIL.n451 585
R1733 VTAIL.n395 VTAIL.n394 585
R1734 VTAIL.n446 VTAIL.n445 585
R1735 VTAIL.n444 VTAIL.n443 585
R1736 VTAIL.n399 VTAIL.n398 585
R1737 VTAIL.n438 VTAIL.n437 585
R1738 VTAIL.n436 VTAIL.n435 585
R1739 VTAIL.n403 VTAIL.n402 585
R1740 VTAIL.n430 VTAIL.n429 585
R1741 VTAIL.n428 VTAIL.n427 585
R1742 VTAIL.n407 VTAIL.n406 585
R1743 VTAIL.n422 VTAIL.n421 585
R1744 VTAIL.n420 VTAIL.n419 585
R1745 VTAIL.n411 VTAIL.n410 585
R1746 VTAIL.n414 VTAIL.n413 585
R1747 VTAIL.n375 VTAIL.n374 585
R1748 VTAIL.n373 VTAIL.n372 585
R1749 VTAIL.n290 VTAIL.n289 585
R1750 VTAIL.n367 VTAIL.n366 585
R1751 VTAIL.n365 VTAIL.n364 585
R1752 VTAIL.n363 VTAIL.n293 585
R1753 VTAIL.n297 VTAIL.n294 585
R1754 VTAIL.n358 VTAIL.n357 585
R1755 VTAIL.n356 VTAIL.n355 585
R1756 VTAIL.n299 VTAIL.n298 585
R1757 VTAIL.n350 VTAIL.n349 585
R1758 VTAIL.n348 VTAIL.n347 585
R1759 VTAIL.n303 VTAIL.n302 585
R1760 VTAIL.n342 VTAIL.n341 585
R1761 VTAIL.n340 VTAIL.n339 585
R1762 VTAIL.n307 VTAIL.n306 585
R1763 VTAIL.n334 VTAIL.n333 585
R1764 VTAIL.n332 VTAIL.n331 585
R1765 VTAIL.n311 VTAIL.n310 585
R1766 VTAIL.n326 VTAIL.n325 585
R1767 VTAIL.n324 VTAIL.n323 585
R1768 VTAIL.n315 VTAIL.n314 585
R1769 VTAIL.n318 VTAIL.n317 585
R1770 VTAIL.t13 VTAIL.n602 327.466
R1771 VTAIL.t8 VTAIL.n506 327.466
R1772 VTAIL.t1 VTAIL.n412 327.466
R1773 VTAIL.t7 VTAIL.n316 327.466
R1774 VTAIL.t4 VTAIL.n695 327.466
R1775 VTAIL.t5 VTAIL.n31 327.466
R1776 VTAIL.t10 VTAIL.n125 327.466
R1777 VTAIL.t12 VTAIL.n221 327.466
R1778 VTAIL.n696 VTAIL.n693 171.744
R1779 VTAIL.n703 VTAIL.n693 171.744
R1780 VTAIL.n704 VTAIL.n703 171.744
R1781 VTAIL.n704 VTAIL.n689 171.744
R1782 VTAIL.n711 VTAIL.n689 171.744
R1783 VTAIL.n712 VTAIL.n711 171.744
R1784 VTAIL.n712 VTAIL.n685 171.744
R1785 VTAIL.n719 VTAIL.n685 171.744
R1786 VTAIL.n720 VTAIL.n719 171.744
R1787 VTAIL.n720 VTAIL.n681 171.744
R1788 VTAIL.n727 VTAIL.n681 171.744
R1789 VTAIL.n728 VTAIL.n727 171.744
R1790 VTAIL.n728 VTAIL.n677 171.744
R1791 VTAIL.n735 VTAIL.n677 171.744
R1792 VTAIL.n737 VTAIL.n735 171.744
R1793 VTAIL.n737 VTAIL.n736 171.744
R1794 VTAIL.n736 VTAIL.n673 171.744
R1795 VTAIL.n745 VTAIL.n673 171.744
R1796 VTAIL.n746 VTAIL.n745 171.744
R1797 VTAIL.n746 VTAIL.n669 171.744
R1798 VTAIL.n753 VTAIL.n669 171.744
R1799 VTAIL.n754 VTAIL.n753 171.744
R1800 VTAIL.n32 VTAIL.n29 171.744
R1801 VTAIL.n39 VTAIL.n29 171.744
R1802 VTAIL.n40 VTAIL.n39 171.744
R1803 VTAIL.n40 VTAIL.n25 171.744
R1804 VTAIL.n47 VTAIL.n25 171.744
R1805 VTAIL.n48 VTAIL.n47 171.744
R1806 VTAIL.n48 VTAIL.n21 171.744
R1807 VTAIL.n55 VTAIL.n21 171.744
R1808 VTAIL.n56 VTAIL.n55 171.744
R1809 VTAIL.n56 VTAIL.n17 171.744
R1810 VTAIL.n63 VTAIL.n17 171.744
R1811 VTAIL.n64 VTAIL.n63 171.744
R1812 VTAIL.n64 VTAIL.n13 171.744
R1813 VTAIL.n71 VTAIL.n13 171.744
R1814 VTAIL.n73 VTAIL.n71 171.744
R1815 VTAIL.n73 VTAIL.n72 171.744
R1816 VTAIL.n72 VTAIL.n9 171.744
R1817 VTAIL.n81 VTAIL.n9 171.744
R1818 VTAIL.n82 VTAIL.n81 171.744
R1819 VTAIL.n82 VTAIL.n5 171.744
R1820 VTAIL.n89 VTAIL.n5 171.744
R1821 VTAIL.n90 VTAIL.n89 171.744
R1822 VTAIL.n126 VTAIL.n123 171.744
R1823 VTAIL.n133 VTAIL.n123 171.744
R1824 VTAIL.n134 VTAIL.n133 171.744
R1825 VTAIL.n134 VTAIL.n119 171.744
R1826 VTAIL.n141 VTAIL.n119 171.744
R1827 VTAIL.n142 VTAIL.n141 171.744
R1828 VTAIL.n142 VTAIL.n115 171.744
R1829 VTAIL.n149 VTAIL.n115 171.744
R1830 VTAIL.n150 VTAIL.n149 171.744
R1831 VTAIL.n150 VTAIL.n111 171.744
R1832 VTAIL.n157 VTAIL.n111 171.744
R1833 VTAIL.n158 VTAIL.n157 171.744
R1834 VTAIL.n158 VTAIL.n107 171.744
R1835 VTAIL.n165 VTAIL.n107 171.744
R1836 VTAIL.n167 VTAIL.n165 171.744
R1837 VTAIL.n167 VTAIL.n166 171.744
R1838 VTAIL.n166 VTAIL.n103 171.744
R1839 VTAIL.n175 VTAIL.n103 171.744
R1840 VTAIL.n176 VTAIL.n175 171.744
R1841 VTAIL.n176 VTAIL.n99 171.744
R1842 VTAIL.n183 VTAIL.n99 171.744
R1843 VTAIL.n184 VTAIL.n183 171.744
R1844 VTAIL.n222 VTAIL.n219 171.744
R1845 VTAIL.n229 VTAIL.n219 171.744
R1846 VTAIL.n230 VTAIL.n229 171.744
R1847 VTAIL.n230 VTAIL.n215 171.744
R1848 VTAIL.n237 VTAIL.n215 171.744
R1849 VTAIL.n238 VTAIL.n237 171.744
R1850 VTAIL.n238 VTAIL.n211 171.744
R1851 VTAIL.n245 VTAIL.n211 171.744
R1852 VTAIL.n246 VTAIL.n245 171.744
R1853 VTAIL.n246 VTAIL.n207 171.744
R1854 VTAIL.n253 VTAIL.n207 171.744
R1855 VTAIL.n254 VTAIL.n253 171.744
R1856 VTAIL.n254 VTAIL.n203 171.744
R1857 VTAIL.n261 VTAIL.n203 171.744
R1858 VTAIL.n263 VTAIL.n261 171.744
R1859 VTAIL.n263 VTAIL.n262 171.744
R1860 VTAIL.n262 VTAIL.n199 171.744
R1861 VTAIL.n271 VTAIL.n199 171.744
R1862 VTAIL.n272 VTAIL.n271 171.744
R1863 VTAIL.n272 VTAIL.n195 171.744
R1864 VTAIL.n279 VTAIL.n195 171.744
R1865 VTAIL.n280 VTAIL.n279 171.744
R1866 VTAIL.n660 VTAIL.n659 171.744
R1867 VTAIL.n659 VTAIL.n575 171.744
R1868 VTAIL.n652 VTAIL.n575 171.744
R1869 VTAIL.n652 VTAIL.n651 171.744
R1870 VTAIL.n651 VTAIL.n579 171.744
R1871 VTAIL.n583 VTAIL.n579 171.744
R1872 VTAIL.n643 VTAIL.n583 171.744
R1873 VTAIL.n643 VTAIL.n642 171.744
R1874 VTAIL.n642 VTAIL.n584 171.744
R1875 VTAIL.n635 VTAIL.n584 171.744
R1876 VTAIL.n635 VTAIL.n634 171.744
R1877 VTAIL.n634 VTAIL.n588 171.744
R1878 VTAIL.n627 VTAIL.n588 171.744
R1879 VTAIL.n627 VTAIL.n626 171.744
R1880 VTAIL.n626 VTAIL.n592 171.744
R1881 VTAIL.n619 VTAIL.n592 171.744
R1882 VTAIL.n619 VTAIL.n618 171.744
R1883 VTAIL.n618 VTAIL.n596 171.744
R1884 VTAIL.n611 VTAIL.n596 171.744
R1885 VTAIL.n611 VTAIL.n610 171.744
R1886 VTAIL.n610 VTAIL.n600 171.744
R1887 VTAIL.n603 VTAIL.n600 171.744
R1888 VTAIL.n564 VTAIL.n563 171.744
R1889 VTAIL.n563 VTAIL.n479 171.744
R1890 VTAIL.n556 VTAIL.n479 171.744
R1891 VTAIL.n556 VTAIL.n555 171.744
R1892 VTAIL.n555 VTAIL.n483 171.744
R1893 VTAIL.n487 VTAIL.n483 171.744
R1894 VTAIL.n547 VTAIL.n487 171.744
R1895 VTAIL.n547 VTAIL.n546 171.744
R1896 VTAIL.n546 VTAIL.n488 171.744
R1897 VTAIL.n539 VTAIL.n488 171.744
R1898 VTAIL.n539 VTAIL.n538 171.744
R1899 VTAIL.n538 VTAIL.n492 171.744
R1900 VTAIL.n531 VTAIL.n492 171.744
R1901 VTAIL.n531 VTAIL.n530 171.744
R1902 VTAIL.n530 VTAIL.n496 171.744
R1903 VTAIL.n523 VTAIL.n496 171.744
R1904 VTAIL.n523 VTAIL.n522 171.744
R1905 VTAIL.n522 VTAIL.n500 171.744
R1906 VTAIL.n515 VTAIL.n500 171.744
R1907 VTAIL.n515 VTAIL.n514 171.744
R1908 VTAIL.n514 VTAIL.n504 171.744
R1909 VTAIL.n507 VTAIL.n504 171.744
R1910 VTAIL.n470 VTAIL.n469 171.744
R1911 VTAIL.n469 VTAIL.n385 171.744
R1912 VTAIL.n462 VTAIL.n385 171.744
R1913 VTAIL.n462 VTAIL.n461 171.744
R1914 VTAIL.n461 VTAIL.n389 171.744
R1915 VTAIL.n393 VTAIL.n389 171.744
R1916 VTAIL.n453 VTAIL.n393 171.744
R1917 VTAIL.n453 VTAIL.n452 171.744
R1918 VTAIL.n452 VTAIL.n394 171.744
R1919 VTAIL.n445 VTAIL.n394 171.744
R1920 VTAIL.n445 VTAIL.n444 171.744
R1921 VTAIL.n444 VTAIL.n398 171.744
R1922 VTAIL.n437 VTAIL.n398 171.744
R1923 VTAIL.n437 VTAIL.n436 171.744
R1924 VTAIL.n436 VTAIL.n402 171.744
R1925 VTAIL.n429 VTAIL.n402 171.744
R1926 VTAIL.n429 VTAIL.n428 171.744
R1927 VTAIL.n428 VTAIL.n406 171.744
R1928 VTAIL.n421 VTAIL.n406 171.744
R1929 VTAIL.n421 VTAIL.n420 171.744
R1930 VTAIL.n420 VTAIL.n410 171.744
R1931 VTAIL.n413 VTAIL.n410 171.744
R1932 VTAIL.n374 VTAIL.n373 171.744
R1933 VTAIL.n373 VTAIL.n289 171.744
R1934 VTAIL.n366 VTAIL.n289 171.744
R1935 VTAIL.n366 VTAIL.n365 171.744
R1936 VTAIL.n365 VTAIL.n293 171.744
R1937 VTAIL.n297 VTAIL.n293 171.744
R1938 VTAIL.n357 VTAIL.n297 171.744
R1939 VTAIL.n357 VTAIL.n356 171.744
R1940 VTAIL.n356 VTAIL.n298 171.744
R1941 VTAIL.n349 VTAIL.n298 171.744
R1942 VTAIL.n349 VTAIL.n348 171.744
R1943 VTAIL.n348 VTAIL.n302 171.744
R1944 VTAIL.n341 VTAIL.n302 171.744
R1945 VTAIL.n341 VTAIL.n340 171.744
R1946 VTAIL.n340 VTAIL.n306 171.744
R1947 VTAIL.n333 VTAIL.n306 171.744
R1948 VTAIL.n333 VTAIL.n332 171.744
R1949 VTAIL.n332 VTAIL.n310 171.744
R1950 VTAIL.n325 VTAIL.n310 171.744
R1951 VTAIL.n325 VTAIL.n324 171.744
R1952 VTAIL.n324 VTAIL.n314 171.744
R1953 VTAIL.n317 VTAIL.n314 171.744
R1954 VTAIL.n696 VTAIL.t4 85.8723
R1955 VTAIL.n32 VTAIL.t5 85.8723
R1956 VTAIL.n126 VTAIL.t10 85.8723
R1957 VTAIL.n222 VTAIL.t12 85.8723
R1958 VTAIL.n603 VTAIL.t13 85.8723
R1959 VTAIL.n507 VTAIL.t8 85.8723
R1960 VTAIL.n413 VTAIL.t1 85.8723
R1961 VTAIL.n317 VTAIL.t7 85.8723
R1962 VTAIL.n571 VTAIL.n570 52.7133
R1963 VTAIL.n381 VTAIL.n380 52.7133
R1964 VTAIL.n1 VTAIL.n0 52.7131
R1965 VTAIL.n191 VTAIL.n190 52.7131
R1966 VTAIL.n759 VTAIL.n758 32.1853
R1967 VTAIL.n95 VTAIL.n94 32.1853
R1968 VTAIL.n189 VTAIL.n188 32.1853
R1969 VTAIL.n285 VTAIL.n284 32.1853
R1970 VTAIL.n665 VTAIL.n664 32.1853
R1971 VTAIL.n569 VTAIL.n568 32.1853
R1972 VTAIL.n475 VTAIL.n474 32.1853
R1973 VTAIL.n379 VTAIL.n378 32.1853
R1974 VTAIL.n759 VTAIL.n665 29.7548
R1975 VTAIL.n379 VTAIL.n285 29.7548
R1976 VTAIL.n697 VTAIL.n695 16.3895
R1977 VTAIL.n33 VTAIL.n31 16.3895
R1978 VTAIL.n127 VTAIL.n125 16.3895
R1979 VTAIL.n223 VTAIL.n221 16.3895
R1980 VTAIL.n604 VTAIL.n602 16.3895
R1981 VTAIL.n508 VTAIL.n506 16.3895
R1982 VTAIL.n414 VTAIL.n412 16.3895
R1983 VTAIL.n318 VTAIL.n316 16.3895
R1984 VTAIL.n744 VTAIL.n743 13.1884
R1985 VTAIL.n80 VTAIL.n79 13.1884
R1986 VTAIL.n174 VTAIL.n173 13.1884
R1987 VTAIL.n270 VTAIL.n269 13.1884
R1988 VTAIL.n650 VTAIL.n649 13.1884
R1989 VTAIL.n554 VTAIL.n553 13.1884
R1990 VTAIL.n460 VTAIL.n459 13.1884
R1991 VTAIL.n364 VTAIL.n363 13.1884
R1992 VTAIL.n698 VTAIL.n694 12.8005
R1993 VTAIL.n742 VTAIL.n674 12.8005
R1994 VTAIL.n747 VTAIL.n672 12.8005
R1995 VTAIL.n34 VTAIL.n30 12.8005
R1996 VTAIL.n78 VTAIL.n10 12.8005
R1997 VTAIL.n83 VTAIL.n8 12.8005
R1998 VTAIL.n128 VTAIL.n124 12.8005
R1999 VTAIL.n172 VTAIL.n104 12.8005
R2000 VTAIL.n177 VTAIL.n102 12.8005
R2001 VTAIL.n224 VTAIL.n220 12.8005
R2002 VTAIL.n268 VTAIL.n200 12.8005
R2003 VTAIL.n273 VTAIL.n198 12.8005
R2004 VTAIL.n653 VTAIL.n578 12.8005
R2005 VTAIL.n648 VTAIL.n580 12.8005
R2006 VTAIL.n605 VTAIL.n601 12.8005
R2007 VTAIL.n557 VTAIL.n482 12.8005
R2008 VTAIL.n552 VTAIL.n484 12.8005
R2009 VTAIL.n509 VTAIL.n505 12.8005
R2010 VTAIL.n463 VTAIL.n388 12.8005
R2011 VTAIL.n458 VTAIL.n390 12.8005
R2012 VTAIL.n415 VTAIL.n411 12.8005
R2013 VTAIL.n367 VTAIL.n292 12.8005
R2014 VTAIL.n362 VTAIL.n294 12.8005
R2015 VTAIL.n319 VTAIL.n315 12.8005
R2016 VTAIL.n702 VTAIL.n701 12.0247
R2017 VTAIL.n739 VTAIL.n738 12.0247
R2018 VTAIL.n748 VTAIL.n670 12.0247
R2019 VTAIL.n38 VTAIL.n37 12.0247
R2020 VTAIL.n75 VTAIL.n74 12.0247
R2021 VTAIL.n84 VTAIL.n6 12.0247
R2022 VTAIL.n132 VTAIL.n131 12.0247
R2023 VTAIL.n169 VTAIL.n168 12.0247
R2024 VTAIL.n178 VTAIL.n100 12.0247
R2025 VTAIL.n228 VTAIL.n227 12.0247
R2026 VTAIL.n265 VTAIL.n264 12.0247
R2027 VTAIL.n274 VTAIL.n196 12.0247
R2028 VTAIL.n654 VTAIL.n576 12.0247
R2029 VTAIL.n645 VTAIL.n644 12.0247
R2030 VTAIL.n609 VTAIL.n608 12.0247
R2031 VTAIL.n558 VTAIL.n480 12.0247
R2032 VTAIL.n549 VTAIL.n548 12.0247
R2033 VTAIL.n513 VTAIL.n512 12.0247
R2034 VTAIL.n464 VTAIL.n386 12.0247
R2035 VTAIL.n455 VTAIL.n454 12.0247
R2036 VTAIL.n419 VTAIL.n418 12.0247
R2037 VTAIL.n368 VTAIL.n290 12.0247
R2038 VTAIL.n359 VTAIL.n358 12.0247
R2039 VTAIL.n323 VTAIL.n322 12.0247
R2040 VTAIL.n705 VTAIL.n692 11.249
R2041 VTAIL.n734 VTAIL.n676 11.249
R2042 VTAIL.n752 VTAIL.n751 11.249
R2043 VTAIL.n41 VTAIL.n28 11.249
R2044 VTAIL.n70 VTAIL.n12 11.249
R2045 VTAIL.n88 VTAIL.n87 11.249
R2046 VTAIL.n135 VTAIL.n122 11.249
R2047 VTAIL.n164 VTAIL.n106 11.249
R2048 VTAIL.n182 VTAIL.n181 11.249
R2049 VTAIL.n231 VTAIL.n218 11.249
R2050 VTAIL.n260 VTAIL.n202 11.249
R2051 VTAIL.n278 VTAIL.n277 11.249
R2052 VTAIL.n658 VTAIL.n657 11.249
R2053 VTAIL.n641 VTAIL.n582 11.249
R2054 VTAIL.n612 VTAIL.n599 11.249
R2055 VTAIL.n562 VTAIL.n561 11.249
R2056 VTAIL.n545 VTAIL.n486 11.249
R2057 VTAIL.n516 VTAIL.n503 11.249
R2058 VTAIL.n468 VTAIL.n467 11.249
R2059 VTAIL.n451 VTAIL.n392 11.249
R2060 VTAIL.n422 VTAIL.n409 11.249
R2061 VTAIL.n372 VTAIL.n371 11.249
R2062 VTAIL.n355 VTAIL.n296 11.249
R2063 VTAIL.n326 VTAIL.n313 11.249
R2064 VTAIL.n706 VTAIL.n690 10.4732
R2065 VTAIL.n733 VTAIL.n678 10.4732
R2066 VTAIL.n755 VTAIL.n668 10.4732
R2067 VTAIL.n42 VTAIL.n26 10.4732
R2068 VTAIL.n69 VTAIL.n14 10.4732
R2069 VTAIL.n91 VTAIL.n4 10.4732
R2070 VTAIL.n136 VTAIL.n120 10.4732
R2071 VTAIL.n163 VTAIL.n108 10.4732
R2072 VTAIL.n185 VTAIL.n98 10.4732
R2073 VTAIL.n232 VTAIL.n216 10.4732
R2074 VTAIL.n259 VTAIL.n204 10.4732
R2075 VTAIL.n281 VTAIL.n194 10.4732
R2076 VTAIL.n661 VTAIL.n574 10.4732
R2077 VTAIL.n640 VTAIL.n585 10.4732
R2078 VTAIL.n613 VTAIL.n597 10.4732
R2079 VTAIL.n565 VTAIL.n478 10.4732
R2080 VTAIL.n544 VTAIL.n489 10.4732
R2081 VTAIL.n517 VTAIL.n501 10.4732
R2082 VTAIL.n471 VTAIL.n384 10.4732
R2083 VTAIL.n450 VTAIL.n395 10.4732
R2084 VTAIL.n423 VTAIL.n407 10.4732
R2085 VTAIL.n375 VTAIL.n288 10.4732
R2086 VTAIL.n354 VTAIL.n299 10.4732
R2087 VTAIL.n327 VTAIL.n311 10.4732
R2088 VTAIL.n710 VTAIL.n709 9.69747
R2089 VTAIL.n730 VTAIL.n729 9.69747
R2090 VTAIL.n756 VTAIL.n666 9.69747
R2091 VTAIL.n46 VTAIL.n45 9.69747
R2092 VTAIL.n66 VTAIL.n65 9.69747
R2093 VTAIL.n92 VTAIL.n2 9.69747
R2094 VTAIL.n140 VTAIL.n139 9.69747
R2095 VTAIL.n160 VTAIL.n159 9.69747
R2096 VTAIL.n186 VTAIL.n96 9.69747
R2097 VTAIL.n236 VTAIL.n235 9.69747
R2098 VTAIL.n256 VTAIL.n255 9.69747
R2099 VTAIL.n282 VTAIL.n192 9.69747
R2100 VTAIL.n662 VTAIL.n572 9.69747
R2101 VTAIL.n637 VTAIL.n636 9.69747
R2102 VTAIL.n617 VTAIL.n616 9.69747
R2103 VTAIL.n566 VTAIL.n476 9.69747
R2104 VTAIL.n541 VTAIL.n540 9.69747
R2105 VTAIL.n521 VTAIL.n520 9.69747
R2106 VTAIL.n472 VTAIL.n382 9.69747
R2107 VTAIL.n447 VTAIL.n446 9.69747
R2108 VTAIL.n427 VTAIL.n426 9.69747
R2109 VTAIL.n376 VTAIL.n286 9.69747
R2110 VTAIL.n351 VTAIL.n350 9.69747
R2111 VTAIL.n331 VTAIL.n330 9.69747
R2112 VTAIL.n758 VTAIL.n757 9.45567
R2113 VTAIL.n94 VTAIL.n93 9.45567
R2114 VTAIL.n188 VTAIL.n187 9.45567
R2115 VTAIL.n284 VTAIL.n283 9.45567
R2116 VTAIL.n664 VTAIL.n663 9.45567
R2117 VTAIL.n568 VTAIL.n567 9.45567
R2118 VTAIL.n474 VTAIL.n473 9.45567
R2119 VTAIL.n378 VTAIL.n377 9.45567
R2120 VTAIL.n757 VTAIL.n756 9.3005
R2121 VTAIL.n668 VTAIL.n667 9.3005
R2122 VTAIL.n751 VTAIL.n750 9.3005
R2123 VTAIL.n749 VTAIL.n748 9.3005
R2124 VTAIL.n672 VTAIL.n671 9.3005
R2125 VTAIL.n717 VTAIL.n716 9.3005
R2126 VTAIL.n715 VTAIL.n714 9.3005
R2127 VTAIL.n688 VTAIL.n687 9.3005
R2128 VTAIL.n709 VTAIL.n708 9.3005
R2129 VTAIL.n707 VTAIL.n706 9.3005
R2130 VTAIL.n692 VTAIL.n691 9.3005
R2131 VTAIL.n701 VTAIL.n700 9.3005
R2132 VTAIL.n699 VTAIL.n698 9.3005
R2133 VTAIL.n684 VTAIL.n683 9.3005
R2134 VTAIL.n723 VTAIL.n722 9.3005
R2135 VTAIL.n725 VTAIL.n724 9.3005
R2136 VTAIL.n680 VTAIL.n679 9.3005
R2137 VTAIL.n731 VTAIL.n730 9.3005
R2138 VTAIL.n733 VTAIL.n732 9.3005
R2139 VTAIL.n676 VTAIL.n675 9.3005
R2140 VTAIL.n740 VTAIL.n739 9.3005
R2141 VTAIL.n742 VTAIL.n741 9.3005
R2142 VTAIL.n93 VTAIL.n92 9.3005
R2143 VTAIL.n4 VTAIL.n3 9.3005
R2144 VTAIL.n87 VTAIL.n86 9.3005
R2145 VTAIL.n85 VTAIL.n84 9.3005
R2146 VTAIL.n8 VTAIL.n7 9.3005
R2147 VTAIL.n53 VTAIL.n52 9.3005
R2148 VTAIL.n51 VTAIL.n50 9.3005
R2149 VTAIL.n24 VTAIL.n23 9.3005
R2150 VTAIL.n45 VTAIL.n44 9.3005
R2151 VTAIL.n43 VTAIL.n42 9.3005
R2152 VTAIL.n28 VTAIL.n27 9.3005
R2153 VTAIL.n37 VTAIL.n36 9.3005
R2154 VTAIL.n35 VTAIL.n34 9.3005
R2155 VTAIL.n20 VTAIL.n19 9.3005
R2156 VTAIL.n59 VTAIL.n58 9.3005
R2157 VTAIL.n61 VTAIL.n60 9.3005
R2158 VTAIL.n16 VTAIL.n15 9.3005
R2159 VTAIL.n67 VTAIL.n66 9.3005
R2160 VTAIL.n69 VTAIL.n68 9.3005
R2161 VTAIL.n12 VTAIL.n11 9.3005
R2162 VTAIL.n76 VTAIL.n75 9.3005
R2163 VTAIL.n78 VTAIL.n77 9.3005
R2164 VTAIL.n187 VTAIL.n186 9.3005
R2165 VTAIL.n98 VTAIL.n97 9.3005
R2166 VTAIL.n181 VTAIL.n180 9.3005
R2167 VTAIL.n179 VTAIL.n178 9.3005
R2168 VTAIL.n102 VTAIL.n101 9.3005
R2169 VTAIL.n147 VTAIL.n146 9.3005
R2170 VTAIL.n145 VTAIL.n144 9.3005
R2171 VTAIL.n118 VTAIL.n117 9.3005
R2172 VTAIL.n139 VTAIL.n138 9.3005
R2173 VTAIL.n137 VTAIL.n136 9.3005
R2174 VTAIL.n122 VTAIL.n121 9.3005
R2175 VTAIL.n131 VTAIL.n130 9.3005
R2176 VTAIL.n129 VTAIL.n128 9.3005
R2177 VTAIL.n114 VTAIL.n113 9.3005
R2178 VTAIL.n153 VTAIL.n152 9.3005
R2179 VTAIL.n155 VTAIL.n154 9.3005
R2180 VTAIL.n110 VTAIL.n109 9.3005
R2181 VTAIL.n161 VTAIL.n160 9.3005
R2182 VTAIL.n163 VTAIL.n162 9.3005
R2183 VTAIL.n106 VTAIL.n105 9.3005
R2184 VTAIL.n170 VTAIL.n169 9.3005
R2185 VTAIL.n172 VTAIL.n171 9.3005
R2186 VTAIL.n283 VTAIL.n282 9.3005
R2187 VTAIL.n194 VTAIL.n193 9.3005
R2188 VTAIL.n277 VTAIL.n276 9.3005
R2189 VTAIL.n275 VTAIL.n274 9.3005
R2190 VTAIL.n198 VTAIL.n197 9.3005
R2191 VTAIL.n243 VTAIL.n242 9.3005
R2192 VTAIL.n241 VTAIL.n240 9.3005
R2193 VTAIL.n214 VTAIL.n213 9.3005
R2194 VTAIL.n235 VTAIL.n234 9.3005
R2195 VTAIL.n233 VTAIL.n232 9.3005
R2196 VTAIL.n218 VTAIL.n217 9.3005
R2197 VTAIL.n227 VTAIL.n226 9.3005
R2198 VTAIL.n225 VTAIL.n224 9.3005
R2199 VTAIL.n210 VTAIL.n209 9.3005
R2200 VTAIL.n249 VTAIL.n248 9.3005
R2201 VTAIL.n251 VTAIL.n250 9.3005
R2202 VTAIL.n206 VTAIL.n205 9.3005
R2203 VTAIL.n257 VTAIL.n256 9.3005
R2204 VTAIL.n259 VTAIL.n258 9.3005
R2205 VTAIL.n202 VTAIL.n201 9.3005
R2206 VTAIL.n266 VTAIL.n265 9.3005
R2207 VTAIL.n268 VTAIL.n267 9.3005
R2208 VTAIL.n630 VTAIL.n629 9.3005
R2209 VTAIL.n632 VTAIL.n631 9.3005
R2210 VTAIL.n587 VTAIL.n586 9.3005
R2211 VTAIL.n638 VTAIL.n637 9.3005
R2212 VTAIL.n640 VTAIL.n639 9.3005
R2213 VTAIL.n582 VTAIL.n581 9.3005
R2214 VTAIL.n646 VTAIL.n645 9.3005
R2215 VTAIL.n648 VTAIL.n647 9.3005
R2216 VTAIL.n663 VTAIL.n662 9.3005
R2217 VTAIL.n574 VTAIL.n573 9.3005
R2218 VTAIL.n657 VTAIL.n656 9.3005
R2219 VTAIL.n655 VTAIL.n654 9.3005
R2220 VTAIL.n578 VTAIL.n577 9.3005
R2221 VTAIL.n591 VTAIL.n590 9.3005
R2222 VTAIL.n624 VTAIL.n623 9.3005
R2223 VTAIL.n622 VTAIL.n621 9.3005
R2224 VTAIL.n595 VTAIL.n594 9.3005
R2225 VTAIL.n616 VTAIL.n615 9.3005
R2226 VTAIL.n614 VTAIL.n613 9.3005
R2227 VTAIL.n599 VTAIL.n598 9.3005
R2228 VTAIL.n608 VTAIL.n607 9.3005
R2229 VTAIL.n606 VTAIL.n605 9.3005
R2230 VTAIL.n534 VTAIL.n533 9.3005
R2231 VTAIL.n536 VTAIL.n535 9.3005
R2232 VTAIL.n491 VTAIL.n490 9.3005
R2233 VTAIL.n542 VTAIL.n541 9.3005
R2234 VTAIL.n544 VTAIL.n543 9.3005
R2235 VTAIL.n486 VTAIL.n485 9.3005
R2236 VTAIL.n550 VTAIL.n549 9.3005
R2237 VTAIL.n552 VTAIL.n551 9.3005
R2238 VTAIL.n567 VTAIL.n566 9.3005
R2239 VTAIL.n478 VTAIL.n477 9.3005
R2240 VTAIL.n561 VTAIL.n560 9.3005
R2241 VTAIL.n559 VTAIL.n558 9.3005
R2242 VTAIL.n482 VTAIL.n481 9.3005
R2243 VTAIL.n495 VTAIL.n494 9.3005
R2244 VTAIL.n528 VTAIL.n527 9.3005
R2245 VTAIL.n526 VTAIL.n525 9.3005
R2246 VTAIL.n499 VTAIL.n498 9.3005
R2247 VTAIL.n520 VTAIL.n519 9.3005
R2248 VTAIL.n518 VTAIL.n517 9.3005
R2249 VTAIL.n503 VTAIL.n502 9.3005
R2250 VTAIL.n512 VTAIL.n511 9.3005
R2251 VTAIL.n510 VTAIL.n509 9.3005
R2252 VTAIL.n440 VTAIL.n439 9.3005
R2253 VTAIL.n442 VTAIL.n441 9.3005
R2254 VTAIL.n397 VTAIL.n396 9.3005
R2255 VTAIL.n448 VTAIL.n447 9.3005
R2256 VTAIL.n450 VTAIL.n449 9.3005
R2257 VTAIL.n392 VTAIL.n391 9.3005
R2258 VTAIL.n456 VTAIL.n455 9.3005
R2259 VTAIL.n458 VTAIL.n457 9.3005
R2260 VTAIL.n473 VTAIL.n472 9.3005
R2261 VTAIL.n384 VTAIL.n383 9.3005
R2262 VTAIL.n467 VTAIL.n466 9.3005
R2263 VTAIL.n465 VTAIL.n464 9.3005
R2264 VTAIL.n388 VTAIL.n387 9.3005
R2265 VTAIL.n401 VTAIL.n400 9.3005
R2266 VTAIL.n434 VTAIL.n433 9.3005
R2267 VTAIL.n432 VTAIL.n431 9.3005
R2268 VTAIL.n405 VTAIL.n404 9.3005
R2269 VTAIL.n426 VTAIL.n425 9.3005
R2270 VTAIL.n424 VTAIL.n423 9.3005
R2271 VTAIL.n409 VTAIL.n408 9.3005
R2272 VTAIL.n418 VTAIL.n417 9.3005
R2273 VTAIL.n416 VTAIL.n415 9.3005
R2274 VTAIL.n344 VTAIL.n343 9.3005
R2275 VTAIL.n346 VTAIL.n345 9.3005
R2276 VTAIL.n301 VTAIL.n300 9.3005
R2277 VTAIL.n352 VTAIL.n351 9.3005
R2278 VTAIL.n354 VTAIL.n353 9.3005
R2279 VTAIL.n296 VTAIL.n295 9.3005
R2280 VTAIL.n360 VTAIL.n359 9.3005
R2281 VTAIL.n362 VTAIL.n361 9.3005
R2282 VTAIL.n377 VTAIL.n376 9.3005
R2283 VTAIL.n288 VTAIL.n287 9.3005
R2284 VTAIL.n371 VTAIL.n370 9.3005
R2285 VTAIL.n369 VTAIL.n368 9.3005
R2286 VTAIL.n292 VTAIL.n291 9.3005
R2287 VTAIL.n305 VTAIL.n304 9.3005
R2288 VTAIL.n338 VTAIL.n337 9.3005
R2289 VTAIL.n336 VTAIL.n335 9.3005
R2290 VTAIL.n309 VTAIL.n308 9.3005
R2291 VTAIL.n330 VTAIL.n329 9.3005
R2292 VTAIL.n328 VTAIL.n327 9.3005
R2293 VTAIL.n313 VTAIL.n312 9.3005
R2294 VTAIL.n322 VTAIL.n321 9.3005
R2295 VTAIL.n320 VTAIL.n319 9.3005
R2296 VTAIL.n713 VTAIL.n688 8.92171
R2297 VTAIL.n726 VTAIL.n680 8.92171
R2298 VTAIL.n49 VTAIL.n24 8.92171
R2299 VTAIL.n62 VTAIL.n16 8.92171
R2300 VTAIL.n143 VTAIL.n118 8.92171
R2301 VTAIL.n156 VTAIL.n110 8.92171
R2302 VTAIL.n239 VTAIL.n214 8.92171
R2303 VTAIL.n252 VTAIL.n206 8.92171
R2304 VTAIL.n633 VTAIL.n587 8.92171
R2305 VTAIL.n620 VTAIL.n595 8.92171
R2306 VTAIL.n537 VTAIL.n491 8.92171
R2307 VTAIL.n524 VTAIL.n499 8.92171
R2308 VTAIL.n443 VTAIL.n397 8.92171
R2309 VTAIL.n430 VTAIL.n405 8.92171
R2310 VTAIL.n347 VTAIL.n301 8.92171
R2311 VTAIL.n334 VTAIL.n309 8.92171
R2312 VTAIL.n714 VTAIL.n686 8.14595
R2313 VTAIL.n725 VTAIL.n682 8.14595
R2314 VTAIL.n50 VTAIL.n22 8.14595
R2315 VTAIL.n61 VTAIL.n18 8.14595
R2316 VTAIL.n144 VTAIL.n116 8.14595
R2317 VTAIL.n155 VTAIL.n112 8.14595
R2318 VTAIL.n240 VTAIL.n212 8.14595
R2319 VTAIL.n251 VTAIL.n208 8.14595
R2320 VTAIL.n632 VTAIL.n589 8.14595
R2321 VTAIL.n621 VTAIL.n593 8.14595
R2322 VTAIL.n536 VTAIL.n493 8.14595
R2323 VTAIL.n525 VTAIL.n497 8.14595
R2324 VTAIL.n442 VTAIL.n399 8.14595
R2325 VTAIL.n431 VTAIL.n403 8.14595
R2326 VTAIL.n346 VTAIL.n303 8.14595
R2327 VTAIL.n335 VTAIL.n307 8.14595
R2328 VTAIL.n718 VTAIL.n717 7.3702
R2329 VTAIL.n722 VTAIL.n721 7.3702
R2330 VTAIL.n54 VTAIL.n53 7.3702
R2331 VTAIL.n58 VTAIL.n57 7.3702
R2332 VTAIL.n148 VTAIL.n147 7.3702
R2333 VTAIL.n152 VTAIL.n151 7.3702
R2334 VTAIL.n244 VTAIL.n243 7.3702
R2335 VTAIL.n248 VTAIL.n247 7.3702
R2336 VTAIL.n629 VTAIL.n628 7.3702
R2337 VTAIL.n625 VTAIL.n624 7.3702
R2338 VTAIL.n533 VTAIL.n532 7.3702
R2339 VTAIL.n529 VTAIL.n528 7.3702
R2340 VTAIL.n439 VTAIL.n438 7.3702
R2341 VTAIL.n435 VTAIL.n434 7.3702
R2342 VTAIL.n343 VTAIL.n342 7.3702
R2343 VTAIL.n339 VTAIL.n338 7.3702
R2344 VTAIL.n718 VTAIL.n684 6.59444
R2345 VTAIL.n721 VTAIL.n684 6.59444
R2346 VTAIL.n54 VTAIL.n20 6.59444
R2347 VTAIL.n57 VTAIL.n20 6.59444
R2348 VTAIL.n148 VTAIL.n114 6.59444
R2349 VTAIL.n151 VTAIL.n114 6.59444
R2350 VTAIL.n244 VTAIL.n210 6.59444
R2351 VTAIL.n247 VTAIL.n210 6.59444
R2352 VTAIL.n628 VTAIL.n591 6.59444
R2353 VTAIL.n625 VTAIL.n591 6.59444
R2354 VTAIL.n532 VTAIL.n495 6.59444
R2355 VTAIL.n529 VTAIL.n495 6.59444
R2356 VTAIL.n438 VTAIL.n401 6.59444
R2357 VTAIL.n435 VTAIL.n401 6.59444
R2358 VTAIL.n342 VTAIL.n305 6.59444
R2359 VTAIL.n339 VTAIL.n305 6.59444
R2360 VTAIL.n717 VTAIL.n686 5.81868
R2361 VTAIL.n722 VTAIL.n682 5.81868
R2362 VTAIL.n53 VTAIL.n22 5.81868
R2363 VTAIL.n58 VTAIL.n18 5.81868
R2364 VTAIL.n147 VTAIL.n116 5.81868
R2365 VTAIL.n152 VTAIL.n112 5.81868
R2366 VTAIL.n243 VTAIL.n212 5.81868
R2367 VTAIL.n248 VTAIL.n208 5.81868
R2368 VTAIL.n629 VTAIL.n589 5.81868
R2369 VTAIL.n624 VTAIL.n593 5.81868
R2370 VTAIL.n533 VTAIL.n493 5.81868
R2371 VTAIL.n528 VTAIL.n497 5.81868
R2372 VTAIL.n439 VTAIL.n399 5.81868
R2373 VTAIL.n434 VTAIL.n403 5.81868
R2374 VTAIL.n343 VTAIL.n303 5.81868
R2375 VTAIL.n338 VTAIL.n307 5.81868
R2376 VTAIL.n714 VTAIL.n713 5.04292
R2377 VTAIL.n726 VTAIL.n725 5.04292
R2378 VTAIL.n50 VTAIL.n49 5.04292
R2379 VTAIL.n62 VTAIL.n61 5.04292
R2380 VTAIL.n144 VTAIL.n143 5.04292
R2381 VTAIL.n156 VTAIL.n155 5.04292
R2382 VTAIL.n240 VTAIL.n239 5.04292
R2383 VTAIL.n252 VTAIL.n251 5.04292
R2384 VTAIL.n633 VTAIL.n632 5.04292
R2385 VTAIL.n621 VTAIL.n620 5.04292
R2386 VTAIL.n537 VTAIL.n536 5.04292
R2387 VTAIL.n525 VTAIL.n524 5.04292
R2388 VTAIL.n443 VTAIL.n442 5.04292
R2389 VTAIL.n431 VTAIL.n430 5.04292
R2390 VTAIL.n347 VTAIL.n346 5.04292
R2391 VTAIL.n335 VTAIL.n334 5.04292
R2392 VTAIL.n710 VTAIL.n688 4.26717
R2393 VTAIL.n729 VTAIL.n680 4.26717
R2394 VTAIL.n758 VTAIL.n666 4.26717
R2395 VTAIL.n46 VTAIL.n24 4.26717
R2396 VTAIL.n65 VTAIL.n16 4.26717
R2397 VTAIL.n94 VTAIL.n2 4.26717
R2398 VTAIL.n140 VTAIL.n118 4.26717
R2399 VTAIL.n159 VTAIL.n110 4.26717
R2400 VTAIL.n188 VTAIL.n96 4.26717
R2401 VTAIL.n236 VTAIL.n214 4.26717
R2402 VTAIL.n255 VTAIL.n206 4.26717
R2403 VTAIL.n284 VTAIL.n192 4.26717
R2404 VTAIL.n664 VTAIL.n572 4.26717
R2405 VTAIL.n636 VTAIL.n587 4.26717
R2406 VTAIL.n617 VTAIL.n595 4.26717
R2407 VTAIL.n568 VTAIL.n476 4.26717
R2408 VTAIL.n540 VTAIL.n491 4.26717
R2409 VTAIL.n521 VTAIL.n499 4.26717
R2410 VTAIL.n474 VTAIL.n382 4.26717
R2411 VTAIL.n446 VTAIL.n397 4.26717
R2412 VTAIL.n427 VTAIL.n405 4.26717
R2413 VTAIL.n378 VTAIL.n286 4.26717
R2414 VTAIL.n350 VTAIL.n301 4.26717
R2415 VTAIL.n331 VTAIL.n309 4.26717
R2416 VTAIL.n699 VTAIL.n695 3.70982
R2417 VTAIL.n35 VTAIL.n31 3.70982
R2418 VTAIL.n129 VTAIL.n125 3.70982
R2419 VTAIL.n225 VTAIL.n221 3.70982
R2420 VTAIL.n606 VTAIL.n602 3.70982
R2421 VTAIL.n510 VTAIL.n506 3.70982
R2422 VTAIL.n416 VTAIL.n412 3.70982
R2423 VTAIL.n320 VTAIL.n316 3.70982
R2424 VTAIL.n709 VTAIL.n690 3.49141
R2425 VTAIL.n730 VTAIL.n678 3.49141
R2426 VTAIL.n756 VTAIL.n755 3.49141
R2427 VTAIL.n45 VTAIL.n26 3.49141
R2428 VTAIL.n66 VTAIL.n14 3.49141
R2429 VTAIL.n92 VTAIL.n91 3.49141
R2430 VTAIL.n139 VTAIL.n120 3.49141
R2431 VTAIL.n160 VTAIL.n108 3.49141
R2432 VTAIL.n186 VTAIL.n185 3.49141
R2433 VTAIL.n235 VTAIL.n216 3.49141
R2434 VTAIL.n256 VTAIL.n204 3.49141
R2435 VTAIL.n282 VTAIL.n281 3.49141
R2436 VTAIL.n662 VTAIL.n661 3.49141
R2437 VTAIL.n637 VTAIL.n585 3.49141
R2438 VTAIL.n616 VTAIL.n597 3.49141
R2439 VTAIL.n566 VTAIL.n565 3.49141
R2440 VTAIL.n541 VTAIL.n489 3.49141
R2441 VTAIL.n520 VTAIL.n501 3.49141
R2442 VTAIL.n472 VTAIL.n471 3.49141
R2443 VTAIL.n447 VTAIL.n395 3.49141
R2444 VTAIL.n426 VTAIL.n407 3.49141
R2445 VTAIL.n376 VTAIL.n375 3.49141
R2446 VTAIL.n351 VTAIL.n299 3.49141
R2447 VTAIL.n330 VTAIL.n311 3.49141
R2448 VTAIL.n381 VTAIL.n379 2.90567
R2449 VTAIL.n475 VTAIL.n381 2.90567
R2450 VTAIL.n571 VTAIL.n569 2.90567
R2451 VTAIL.n665 VTAIL.n571 2.90567
R2452 VTAIL.n285 VTAIL.n191 2.90567
R2453 VTAIL.n191 VTAIL.n189 2.90567
R2454 VTAIL.n95 VTAIL.n1 2.90567
R2455 VTAIL VTAIL.n759 2.84748
R2456 VTAIL.n706 VTAIL.n705 2.71565
R2457 VTAIL.n734 VTAIL.n733 2.71565
R2458 VTAIL.n752 VTAIL.n668 2.71565
R2459 VTAIL.n42 VTAIL.n41 2.71565
R2460 VTAIL.n70 VTAIL.n69 2.71565
R2461 VTAIL.n88 VTAIL.n4 2.71565
R2462 VTAIL.n136 VTAIL.n135 2.71565
R2463 VTAIL.n164 VTAIL.n163 2.71565
R2464 VTAIL.n182 VTAIL.n98 2.71565
R2465 VTAIL.n232 VTAIL.n231 2.71565
R2466 VTAIL.n260 VTAIL.n259 2.71565
R2467 VTAIL.n278 VTAIL.n194 2.71565
R2468 VTAIL.n658 VTAIL.n574 2.71565
R2469 VTAIL.n641 VTAIL.n640 2.71565
R2470 VTAIL.n613 VTAIL.n612 2.71565
R2471 VTAIL.n562 VTAIL.n478 2.71565
R2472 VTAIL.n545 VTAIL.n544 2.71565
R2473 VTAIL.n517 VTAIL.n516 2.71565
R2474 VTAIL.n468 VTAIL.n384 2.71565
R2475 VTAIL.n451 VTAIL.n450 2.71565
R2476 VTAIL.n423 VTAIL.n422 2.71565
R2477 VTAIL.n372 VTAIL.n288 2.71565
R2478 VTAIL.n355 VTAIL.n354 2.71565
R2479 VTAIL.n327 VTAIL.n326 2.71565
R2480 VTAIL.n702 VTAIL.n692 1.93989
R2481 VTAIL.n738 VTAIL.n676 1.93989
R2482 VTAIL.n751 VTAIL.n670 1.93989
R2483 VTAIL.n38 VTAIL.n28 1.93989
R2484 VTAIL.n74 VTAIL.n12 1.93989
R2485 VTAIL.n87 VTAIL.n6 1.93989
R2486 VTAIL.n132 VTAIL.n122 1.93989
R2487 VTAIL.n168 VTAIL.n106 1.93989
R2488 VTAIL.n181 VTAIL.n100 1.93989
R2489 VTAIL.n228 VTAIL.n218 1.93989
R2490 VTAIL.n264 VTAIL.n202 1.93989
R2491 VTAIL.n277 VTAIL.n196 1.93989
R2492 VTAIL.n657 VTAIL.n576 1.93989
R2493 VTAIL.n644 VTAIL.n582 1.93989
R2494 VTAIL.n609 VTAIL.n599 1.93989
R2495 VTAIL.n561 VTAIL.n480 1.93989
R2496 VTAIL.n548 VTAIL.n486 1.93989
R2497 VTAIL.n513 VTAIL.n503 1.93989
R2498 VTAIL.n467 VTAIL.n386 1.93989
R2499 VTAIL.n454 VTAIL.n392 1.93989
R2500 VTAIL.n419 VTAIL.n409 1.93989
R2501 VTAIL.n371 VTAIL.n290 1.93989
R2502 VTAIL.n358 VTAIL.n296 1.93989
R2503 VTAIL.n323 VTAIL.n313 1.93989
R2504 VTAIL.n0 VTAIL.t2 1.93532
R2505 VTAIL.n0 VTAIL.t3 1.93532
R2506 VTAIL.n190 VTAIL.t9 1.93532
R2507 VTAIL.n190 VTAIL.t11 1.93532
R2508 VTAIL.n570 VTAIL.t14 1.93532
R2509 VTAIL.n570 VTAIL.t15 1.93532
R2510 VTAIL.n380 VTAIL.t0 1.93532
R2511 VTAIL.n380 VTAIL.t6 1.93532
R2512 VTAIL.n701 VTAIL.n694 1.16414
R2513 VTAIL.n739 VTAIL.n674 1.16414
R2514 VTAIL.n748 VTAIL.n747 1.16414
R2515 VTAIL.n37 VTAIL.n30 1.16414
R2516 VTAIL.n75 VTAIL.n10 1.16414
R2517 VTAIL.n84 VTAIL.n83 1.16414
R2518 VTAIL.n131 VTAIL.n124 1.16414
R2519 VTAIL.n169 VTAIL.n104 1.16414
R2520 VTAIL.n178 VTAIL.n177 1.16414
R2521 VTAIL.n227 VTAIL.n220 1.16414
R2522 VTAIL.n265 VTAIL.n200 1.16414
R2523 VTAIL.n274 VTAIL.n273 1.16414
R2524 VTAIL.n654 VTAIL.n653 1.16414
R2525 VTAIL.n645 VTAIL.n580 1.16414
R2526 VTAIL.n608 VTAIL.n601 1.16414
R2527 VTAIL.n558 VTAIL.n557 1.16414
R2528 VTAIL.n549 VTAIL.n484 1.16414
R2529 VTAIL.n512 VTAIL.n505 1.16414
R2530 VTAIL.n464 VTAIL.n463 1.16414
R2531 VTAIL.n455 VTAIL.n390 1.16414
R2532 VTAIL.n418 VTAIL.n411 1.16414
R2533 VTAIL.n368 VTAIL.n367 1.16414
R2534 VTAIL.n359 VTAIL.n294 1.16414
R2535 VTAIL.n322 VTAIL.n315 1.16414
R2536 VTAIL.n569 VTAIL.n475 0.470328
R2537 VTAIL.n189 VTAIL.n95 0.470328
R2538 VTAIL.n698 VTAIL.n697 0.388379
R2539 VTAIL.n743 VTAIL.n742 0.388379
R2540 VTAIL.n744 VTAIL.n672 0.388379
R2541 VTAIL.n34 VTAIL.n33 0.388379
R2542 VTAIL.n79 VTAIL.n78 0.388379
R2543 VTAIL.n80 VTAIL.n8 0.388379
R2544 VTAIL.n128 VTAIL.n127 0.388379
R2545 VTAIL.n173 VTAIL.n172 0.388379
R2546 VTAIL.n174 VTAIL.n102 0.388379
R2547 VTAIL.n224 VTAIL.n223 0.388379
R2548 VTAIL.n269 VTAIL.n268 0.388379
R2549 VTAIL.n270 VTAIL.n198 0.388379
R2550 VTAIL.n650 VTAIL.n578 0.388379
R2551 VTAIL.n649 VTAIL.n648 0.388379
R2552 VTAIL.n605 VTAIL.n604 0.388379
R2553 VTAIL.n554 VTAIL.n482 0.388379
R2554 VTAIL.n553 VTAIL.n552 0.388379
R2555 VTAIL.n509 VTAIL.n508 0.388379
R2556 VTAIL.n460 VTAIL.n388 0.388379
R2557 VTAIL.n459 VTAIL.n458 0.388379
R2558 VTAIL.n415 VTAIL.n414 0.388379
R2559 VTAIL.n364 VTAIL.n292 0.388379
R2560 VTAIL.n363 VTAIL.n362 0.388379
R2561 VTAIL.n319 VTAIL.n318 0.388379
R2562 VTAIL.n700 VTAIL.n699 0.155672
R2563 VTAIL.n700 VTAIL.n691 0.155672
R2564 VTAIL.n707 VTAIL.n691 0.155672
R2565 VTAIL.n708 VTAIL.n707 0.155672
R2566 VTAIL.n708 VTAIL.n687 0.155672
R2567 VTAIL.n715 VTAIL.n687 0.155672
R2568 VTAIL.n716 VTAIL.n715 0.155672
R2569 VTAIL.n716 VTAIL.n683 0.155672
R2570 VTAIL.n723 VTAIL.n683 0.155672
R2571 VTAIL.n724 VTAIL.n723 0.155672
R2572 VTAIL.n724 VTAIL.n679 0.155672
R2573 VTAIL.n731 VTAIL.n679 0.155672
R2574 VTAIL.n732 VTAIL.n731 0.155672
R2575 VTAIL.n732 VTAIL.n675 0.155672
R2576 VTAIL.n740 VTAIL.n675 0.155672
R2577 VTAIL.n741 VTAIL.n740 0.155672
R2578 VTAIL.n741 VTAIL.n671 0.155672
R2579 VTAIL.n749 VTAIL.n671 0.155672
R2580 VTAIL.n750 VTAIL.n749 0.155672
R2581 VTAIL.n750 VTAIL.n667 0.155672
R2582 VTAIL.n757 VTAIL.n667 0.155672
R2583 VTAIL.n36 VTAIL.n35 0.155672
R2584 VTAIL.n36 VTAIL.n27 0.155672
R2585 VTAIL.n43 VTAIL.n27 0.155672
R2586 VTAIL.n44 VTAIL.n43 0.155672
R2587 VTAIL.n44 VTAIL.n23 0.155672
R2588 VTAIL.n51 VTAIL.n23 0.155672
R2589 VTAIL.n52 VTAIL.n51 0.155672
R2590 VTAIL.n52 VTAIL.n19 0.155672
R2591 VTAIL.n59 VTAIL.n19 0.155672
R2592 VTAIL.n60 VTAIL.n59 0.155672
R2593 VTAIL.n60 VTAIL.n15 0.155672
R2594 VTAIL.n67 VTAIL.n15 0.155672
R2595 VTAIL.n68 VTAIL.n67 0.155672
R2596 VTAIL.n68 VTAIL.n11 0.155672
R2597 VTAIL.n76 VTAIL.n11 0.155672
R2598 VTAIL.n77 VTAIL.n76 0.155672
R2599 VTAIL.n77 VTAIL.n7 0.155672
R2600 VTAIL.n85 VTAIL.n7 0.155672
R2601 VTAIL.n86 VTAIL.n85 0.155672
R2602 VTAIL.n86 VTAIL.n3 0.155672
R2603 VTAIL.n93 VTAIL.n3 0.155672
R2604 VTAIL.n130 VTAIL.n129 0.155672
R2605 VTAIL.n130 VTAIL.n121 0.155672
R2606 VTAIL.n137 VTAIL.n121 0.155672
R2607 VTAIL.n138 VTAIL.n137 0.155672
R2608 VTAIL.n138 VTAIL.n117 0.155672
R2609 VTAIL.n145 VTAIL.n117 0.155672
R2610 VTAIL.n146 VTAIL.n145 0.155672
R2611 VTAIL.n146 VTAIL.n113 0.155672
R2612 VTAIL.n153 VTAIL.n113 0.155672
R2613 VTAIL.n154 VTAIL.n153 0.155672
R2614 VTAIL.n154 VTAIL.n109 0.155672
R2615 VTAIL.n161 VTAIL.n109 0.155672
R2616 VTAIL.n162 VTAIL.n161 0.155672
R2617 VTAIL.n162 VTAIL.n105 0.155672
R2618 VTAIL.n170 VTAIL.n105 0.155672
R2619 VTAIL.n171 VTAIL.n170 0.155672
R2620 VTAIL.n171 VTAIL.n101 0.155672
R2621 VTAIL.n179 VTAIL.n101 0.155672
R2622 VTAIL.n180 VTAIL.n179 0.155672
R2623 VTAIL.n180 VTAIL.n97 0.155672
R2624 VTAIL.n187 VTAIL.n97 0.155672
R2625 VTAIL.n226 VTAIL.n225 0.155672
R2626 VTAIL.n226 VTAIL.n217 0.155672
R2627 VTAIL.n233 VTAIL.n217 0.155672
R2628 VTAIL.n234 VTAIL.n233 0.155672
R2629 VTAIL.n234 VTAIL.n213 0.155672
R2630 VTAIL.n241 VTAIL.n213 0.155672
R2631 VTAIL.n242 VTAIL.n241 0.155672
R2632 VTAIL.n242 VTAIL.n209 0.155672
R2633 VTAIL.n249 VTAIL.n209 0.155672
R2634 VTAIL.n250 VTAIL.n249 0.155672
R2635 VTAIL.n250 VTAIL.n205 0.155672
R2636 VTAIL.n257 VTAIL.n205 0.155672
R2637 VTAIL.n258 VTAIL.n257 0.155672
R2638 VTAIL.n258 VTAIL.n201 0.155672
R2639 VTAIL.n266 VTAIL.n201 0.155672
R2640 VTAIL.n267 VTAIL.n266 0.155672
R2641 VTAIL.n267 VTAIL.n197 0.155672
R2642 VTAIL.n275 VTAIL.n197 0.155672
R2643 VTAIL.n276 VTAIL.n275 0.155672
R2644 VTAIL.n276 VTAIL.n193 0.155672
R2645 VTAIL.n283 VTAIL.n193 0.155672
R2646 VTAIL.n663 VTAIL.n573 0.155672
R2647 VTAIL.n656 VTAIL.n573 0.155672
R2648 VTAIL.n656 VTAIL.n655 0.155672
R2649 VTAIL.n655 VTAIL.n577 0.155672
R2650 VTAIL.n647 VTAIL.n577 0.155672
R2651 VTAIL.n647 VTAIL.n646 0.155672
R2652 VTAIL.n646 VTAIL.n581 0.155672
R2653 VTAIL.n639 VTAIL.n581 0.155672
R2654 VTAIL.n639 VTAIL.n638 0.155672
R2655 VTAIL.n638 VTAIL.n586 0.155672
R2656 VTAIL.n631 VTAIL.n586 0.155672
R2657 VTAIL.n631 VTAIL.n630 0.155672
R2658 VTAIL.n630 VTAIL.n590 0.155672
R2659 VTAIL.n623 VTAIL.n590 0.155672
R2660 VTAIL.n623 VTAIL.n622 0.155672
R2661 VTAIL.n622 VTAIL.n594 0.155672
R2662 VTAIL.n615 VTAIL.n594 0.155672
R2663 VTAIL.n615 VTAIL.n614 0.155672
R2664 VTAIL.n614 VTAIL.n598 0.155672
R2665 VTAIL.n607 VTAIL.n598 0.155672
R2666 VTAIL.n607 VTAIL.n606 0.155672
R2667 VTAIL.n567 VTAIL.n477 0.155672
R2668 VTAIL.n560 VTAIL.n477 0.155672
R2669 VTAIL.n560 VTAIL.n559 0.155672
R2670 VTAIL.n559 VTAIL.n481 0.155672
R2671 VTAIL.n551 VTAIL.n481 0.155672
R2672 VTAIL.n551 VTAIL.n550 0.155672
R2673 VTAIL.n550 VTAIL.n485 0.155672
R2674 VTAIL.n543 VTAIL.n485 0.155672
R2675 VTAIL.n543 VTAIL.n542 0.155672
R2676 VTAIL.n542 VTAIL.n490 0.155672
R2677 VTAIL.n535 VTAIL.n490 0.155672
R2678 VTAIL.n535 VTAIL.n534 0.155672
R2679 VTAIL.n534 VTAIL.n494 0.155672
R2680 VTAIL.n527 VTAIL.n494 0.155672
R2681 VTAIL.n527 VTAIL.n526 0.155672
R2682 VTAIL.n526 VTAIL.n498 0.155672
R2683 VTAIL.n519 VTAIL.n498 0.155672
R2684 VTAIL.n519 VTAIL.n518 0.155672
R2685 VTAIL.n518 VTAIL.n502 0.155672
R2686 VTAIL.n511 VTAIL.n502 0.155672
R2687 VTAIL.n511 VTAIL.n510 0.155672
R2688 VTAIL.n473 VTAIL.n383 0.155672
R2689 VTAIL.n466 VTAIL.n383 0.155672
R2690 VTAIL.n466 VTAIL.n465 0.155672
R2691 VTAIL.n465 VTAIL.n387 0.155672
R2692 VTAIL.n457 VTAIL.n387 0.155672
R2693 VTAIL.n457 VTAIL.n456 0.155672
R2694 VTAIL.n456 VTAIL.n391 0.155672
R2695 VTAIL.n449 VTAIL.n391 0.155672
R2696 VTAIL.n449 VTAIL.n448 0.155672
R2697 VTAIL.n448 VTAIL.n396 0.155672
R2698 VTAIL.n441 VTAIL.n396 0.155672
R2699 VTAIL.n441 VTAIL.n440 0.155672
R2700 VTAIL.n440 VTAIL.n400 0.155672
R2701 VTAIL.n433 VTAIL.n400 0.155672
R2702 VTAIL.n433 VTAIL.n432 0.155672
R2703 VTAIL.n432 VTAIL.n404 0.155672
R2704 VTAIL.n425 VTAIL.n404 0.155672
R2705 VTAIL.n425 VTAIL.n424 0.155672
R2706 VTAIL.n424 VTAIL.n408 0.155672
R2707 VTAIL.n417 VTAIL.n408 0.155672
R2708 VTAIL.n417 VTAIL.n416 0.155672
R2709 VTAIL.n377 VTAIL.n287 0.155672
R2710 VTAIL.n370 VTAIL.n287 0.155672
R2711 VTAIL.n370 VTAIL.n369 0.155672
R2712 VTAIL.n369 VTAIL.n291 0.155672
R2713 VTAIL.n361 VTAIL.n291 0.155672
R2714 VTAIL.n361 VTAIL.n360 0.155672
R2715 VTAIL.n360 VTAIL.n295 0.155672
R2716 VTAIL.n353 VTAIL.n295 0.155672
R2717 VTAIL.n353 VTAIL.n352 0.155672
R2718 VTAIL.n352 VTAIL.n300 0.155672
R2719 VTAIL.n345 VTAIL.n300 0.155672
R2720 VTAIL.n345 VTAIL.n344 0.155672
R2721 VTAIL.n344 VTAIL.n304 0.155672
R2722 VTAIL.n337 VTAIL.n304 0.155672
R2723 VTAIL.n337 VTAIL.n336 0.155672
R2724 VTAIL.n336 VTAIL.n308 0.155672
R2725 VTAIL.n329 VTAIL.n308 0.155672
R2726 VTAIL.n329 VTAIL.n328 0.155672
R2727 VTAIL.n328 VTAIL.n312 0.155672
R2728 VTAIL.n321 VTAIL.n312 0.155672
R2729 VTAIL.n321 VTAIL.n320 0.155672
R2730 VTAIL VTAIL.n1 0.0586897
R2731 VN.n39 VN.t3 166.341
R2732 VN.n8 VN.t1 166.341
R2733 VN.n60 VN.n59 161.3
R2734 VN.n58 VN.n32 161.3
R2735 VN.n57 VN.n56 161.3
R2736 VN.n55 VN.n33 161.3
R2737 VN.n54 VN.n53 161.3
R2738 VN.n52 VN.n34 161.3
R2739 VN.n51 VN.n50 161.3
R2740 VN.n49 VN.n48 161.3
R2741 VN.n47 VN.n36 161.3
R2742 VN.n46 VN.n45 161.3
R2743 VN.n44 VN.n37 161.3
R2744 VN.n43 VN.n42 161.3
R2745 VN.n41 VN.n38 161.3
R2746 VN.n29 VN.n28 161.3
R2747 VN.n27 VN.n1 161.3
R2748 VN.n26 VN.n25 161.3
R2749 VN.n24 VN.n2 161.3
R2750 VN.n23 VN.n22 161.3
R2751 VN.n21 VN.n3 161.3
R2752 VN.n20 VN.n19 161.3
R2753 VN.n18 VN.n17 161.3
R2754 VN.n16 VN.n5 161.3
R2755 VN.n15 VN.n14 161.3
R2756 VN.n13 VN.n6 161.3
R2757 VN.n12 VN.n11 161.3
R2758 VN.n10 VN.n7 161.3
R2759 VN.n9 VN.t5 133.185
R2760 VN.n4 VN.t2 133.185
R2761 VN.n0 VN.t6 133.185
R2762 VN.n40 VN.t4 133.185
R2763 VN.n35 VN.t7 133.185
R2764 VN.n31 VN.t0 133.185
R2765 VN.n30 VN.n0 75.2445
R2766 VN.n61 VN.n31 75.2445
R2767 VN VN.n61 56.8087
R2768 VN.n15 VN.n6 56.5617
R2769 VN.n46 VN.n37 56.5617
R2770 VN.n9 VN.n8 52.6903
R2771 VN.n40 VN.n39 52.6903
R2772 VN.n26 VN.n2 52.2023
R2773 VN.n57 VN.n33 52.2023
R2774 VN.n22 VN.n2 28.9518
R2775 VN.n53 VN.n33 28.9518
R2776 VN.n11 VN.n10 24.5923
R2777 VN.n11 VN.n6 24.5923
R2778 VN.n16 VN.n15 24.5923
R2779 VN.n17 VN.n16 24.5923
R2780 VN.n21 VN.n20 24.5923
R2781 VN.n22 VN.n21 24.5923
R2782 VN.n27 VN.n26 24.5923
R2783 VN.n28 VN.n27 24.5923
R2784 VN.n42 VN.n37 24.5923
R2785 VN.n42 VN.n41 24.5923
R2786 VN.n53 VN.n52 24.5923
R2787 VN.n52 VN.n51 24.5923
R2788 VN.n48 VN.n47 24.5923
R2789 VN.n47 VN.n46 24.5923
R2790 VN.n59 VN.n58 24.5923
R2791 VN.n58 VN.n57 24.5923
R2792 VN.n10 VN.n9 21.3954
R2793 VN.n17 VN.n4 21.3954
R2794 VN.n41 VN.n40 21.3954
R2795 VN.n48 VN.n35 21.3954
R2796 VN.n28 VN.n0 15.0015
R2797 VN.n59 VN.n31 15.0015
R2798 VN.n8 VN.n7 4.13672
R2799 VN.n39 VN.n38 4.13672
R2800 VN.n20 VN.n4 3.19744
R2801 VN.n51 VN.n35 3.19744
R2802 VN.n61 VN.n60 0.354861
R2803 VN.n30 VN.n29 0.354861
R2804 VN VN.n30 0.267071
R2805 VN.n60 VN.n32 0.189894
R2806 VN.n56 VN.n32 0.189894
R2807 VN.n56 VN.n55 0.189894
R2808 VN.n55 VN.n54 0.189894
R2809 VN.n54 VN.n34 0.189894
R2810 VN.n50 VN.n34 0.189894
R2811 VN.n50 VN.n49 0.189894
R2812 VN.n49 VN.n36 0.189894
R2813 VN.n45 VN.n36 0.189894
R2814 VN.n45 VN.n44 0.189894
R2815 VN.n44 VN.n43 0.189894
R2816 VN.n43 VN.n38 0.189894
R2817 VN.n12 VN.n7 0.189894
R2818 VN.n13 VN.n12 0.189894
R2819 VN.n14 VN.n13 0.189894
R2820 VN.n14 VN.n5 0.189894
R2821 VN.n18 VN.n5 0.189894
R2822 VN.n19 VN.n18 0.189894
R2823 VN.n19 VN.n3 0.189894
R2824 VN.n23 VN.n3 0.189894
R2825 VN.n24 VN.n23 0.189894
R2826 VN.n25 VN.n24 0.189894
R2827 VN.n25 VN.n1 0.189894
R2828 VN.n29 VN.n1 0.189894
R2829 VDD2.n2 VDD2.n1 70.7891
R2830 VDD2.n2 VDD2.n0 70.7891
R2831 VDD2 VDD2.n5 70.7862
R2832 VDD2.n4 VDD2.n3 69.392
R2833 VDD2.n4 VDD2.n2 51.2713
R2834 VDD2.n5 VDD2.t3 1.93532
R2835 VDD2.n5 VDD2.t4 1.93532
R2836 VDD2.n3 VDD2.t7 1.93532
R2837 VDD2.n3 VDD2.t0 1.93532
R2838 VDD2.n1 VDD2.t5 1.93532
R2839 VDD2.n1 VDD2.t1 1.93532
R2840 VDD2.n0 VDD2.t6 1.93532
R2841 VDD2.n0 VDD2.t2 1.93532
R2842 VDD2 VDD2.n4 1.51128
C0 VDD1 VDD2 2.00621f
C1 B w_n4340_n4328# 12.135099f
C2 VP w_n4340_n4328# 9.608179f
C3 B VP 2.33712f
C4 VN w_n4340_n4328# 9.04346f
C5 VTAIL w_n4340_n4328# 5.31438f
C6 VN B 1.38811f
C7 VTAIL B 6.78812f
C8 VN VP 9.088019f
C9 VDD1 w_n4340_n4328# 2.22506f
C10 VDD2 w_n4340_n4328# 2.35823f
C11 VTAIL VP 12.6797f
C12 VDD1 B 1.9124f
C13 VDD2 B 2.02227f
C14 VN VTAIL 12.6656f
C15 VDD1 VP 12.7537f
C16 VDD2 VP 0.566769f
C17 VDD1 VN 0.152801f
C18 VDD2 VN 12.3413f
C19 VDD1 VTAIL 9.69417f
C20 VDD2 VTAIL 9.751539f
C21 VDD2 VSUBS 2.320287f
C22 VDD1 VSUBS 2.94915f
C23 VTAIL VSUBS 1.626563f
C24 VN VSUBS 7.4973f
C25 VP VSUBS 4.218628f
C26 B VSUBS 5.90122f
C27 w_n4340_n4328# VSUBS 0.229933p
C28 VDD2.t6 VSUBS 0.414116f
C29 VDD2.t2 VSUBS 0.414116f
C30 VDD2.n0 VSUBS 3.43084f
C31 VDD2.t5 VSUBS 0.414116f
C32 VDD2.t1 VSUBS 0.414116f
C33 VDD2.n1 VSUBS 3.43084f
C34 VDD2.n2 VSUBS 5.48183f
C35 VDD2.t7 VSUBS 0.414116f
C36 VDD2.t0 VSUBS 0.414116f
C37 VDD2.n3 VSUBS 3.41002f
C38 VDD2.n4 VSUBS 4.67707f
C39 VDD2.t3 VSUBS 0.414116f
C40 VDD2.t4 VSUBS 0.414116f
C41 VDD2.n5 VSUBS 3.43078f
C42 VN.t6 VSUBS 3.40075f
C43 VN.n0 VSUBS 1.26707f
C44 VN.n1 VSUBS 0.024241f
C45 VN.n2 VSUBS 0.024427f
C46 VN.n3 VSUBS 0.024241f
C47 VN.t2 VSUBS 3.40075f
C48 VN.n4 VSUBS 1.17872f
C49 VN.n5 VSUBS 0.024241f
C50 VN.n6 VSUBS 0.035238f
C51 VN.n7 VSUBS 0.276912f
C52 VN.t5 VSUBS 3.40075f
C53 VN.t1 VSUBS 3.66849f
C54 VN.n8 VSUBS 1.21221f
C55 VN.n9 VSUBS 1.26474f
C56 VN.n10 VSUBS 0.042068f
C57 VN.n11 VSUBS 0.044953f
C58 VN.n12 VSUBS 0.024241f
C59 VN.n13 VSUBS 0.024241f
C60 VN.n14 VSUBS 0.024241f
C61 VN.n15 VSUBS 0.035238f
C62 VN.n16 VSUBS 0.044953f
C63 VN.n17 VSUBS 0.042068f
C64 VN.n18 VSUBS 0.024241f
C65 VN.n19 VSUBS 0.024241f
C66 VN.n20 VSUBS 0.025646f
C67 VN.n21 VSUBS 0.044953f
C68 VN.n22 VSUBS 0.047693f
C69 VN.n23 VSUBS 0.024241f
C70 VN.n24 VSUBS 0.024241f
C71 VN.n25 VSUBS 0.024241f
C72 VN.n26 VSUBS 0.04331f
C73 VN.n27 VSUBS 0.044953f
C74 VN.n28 VSUBS 0.036298f
C75 VN.n29 VSUBS 0.039119f
C76 VN.n30 VSUBS 0.055803f
C77 VN.t0 VSUBS 3.40075f
C78 VN.n31 VSUBS 1.26707f
C79 VN.n32 VSUBS 0.024241f
C80 VN.n33 VSUBS 0.024427f
C81 VN.n34 VSUBS 0.024241f
C82 VN.t7 VSUBS 3.40075f
C83 VN.n35 VSUBS 1.17872f
C84 VN.n36 VSUBS 0.024241f
C85 VN.n37 VSUBS 0.035238f
C86 VN.n38 VSUBS 0.276912f
C87 VN.t4 VSUBS 3.40075f
C88 VN.t3 VSUBS 3.66849f
C89 VN.n39 VSUBS 1.21221f
C90 VN.n40 VSUBS 1.26474f
C91 VN.n41 VSUBS 0.042068f
C92 VN.n42 VSUBS 0.044953f
C93 VN.n43 VSUBS 0.024241f
C94 VN.n44 VSUBS 0.024241f
C95 VN.n45 VSUBS 0.024241f
C96 VN.n46 VSUBS 0.035238f
C97 VN.n47 VSUBS 0.044953f
C98 VN.n48 VSUBS 0.042068f
C99 VN.n49 VSUBS 0.024241f
C100 VN.n50 VSUBS 0.024241f
C101 VN.n51 VSUBS 0.025646f
C102 VN.n52 VSUBS 0.044953f
C103 VN.n53 VSUBS 0.047693f
C104 VN.n54 VSUBS 0.024241f
C105 VN.n55 VSUBS 0.024241f
C106 VN.n56 VSUBS 0.024241f
C107 VN.n57 VSUBS 0.04331f
C108 VN.n58 VSUBS 0.044953f
C109 VN.n59 VSUBS 0.036298f
C110 VN.n60 VSUBS 0.039119f
C111 VN.n61 VSUBS 1.64681f
C112 VTAIL.t2 VSUBS 0.320615f
C113 VTAIL.t3 VSUBS 0.320615f
C114 VTAIL.n0 VSUBS 2.49217f
C115 VTAIL.n1 VSUBS 0.817754f
C116 VTAIL.n2 VSUBS 0.025616f
C117 VTAIL.n3 VSUBS 0.02415f
C118 VTAIL.n4 VSUBS 0.012977f
C119 VTAIL.n5 VSUBS 0.030674f
C120 VTAIL.n6 VSUBS 0.013741f
C121 VTAIL.n7 VSUBS 0.02415f
C122 VTAIL.n8 VSUBS 0.012977f
C123 VTAIL.n9 VSUBS 0.030674f
C124 VTAIL.n10 VSUBS 0.013741f
C125 VTAIL.n11 VSUBS 0.02415f
C126 VTAIL.n12 VSUBS 0.012977f
C127 VTAIL.n13 VSUBS 0.030674f
C128 VTAIL.n14 VSUBS 0.013741f
C129 VTAIL.n15 VSUBS 0.02415f
C130 VTAIL.n16 VSUBS 0.012977f
C131 VTAIL.n17 VSUBS 0.030674f
C132 VTAIL.n18 VSUBS 0.013741f
C133 VTAIL.n19 VSUBS 0.02415f
C134 VTAIL.n20 VSUBS 0.012977f
C135 VTAIL.n21 VSUBS 0.030674f
C136 VTAIL.n22 VSUBS 0.013741f
C137 VTAIL.n23 VSUBS 0.02415f
C138 VTAIL.n24 VSUBS 0.012977f
C139 VTAIL.n25 VSUBS 0.030674f
C140 VTAIL.n26 VSUBS 0.013741f
C141 VTAIL.n27 VSUBS 0.02415f
C142 VTAIL.n28 VSUBS 0.012977f
C143 VTAIL.n29 VSUBS 0.030674f
C144 VTAIL.n30 VSUBS 0.013741f
C145 VTAIL.n31 VSUBS 0.18306f
C146 VTAIL.t5 VSUBS 0.065774f
C147 VTAIL.n32 VSUBS 0.023005f
C148 VTAIL.n33 VSUBS 0.019513f
C149 VTAIL.n34 VSUBS 0.012977f
C150 VTAIL.n35 VSUBS 1.73938f
C151 VTAIL.n36 VSUBS 0.02415f
C152 VTAIL.n37 VSUBS 0.012977f
C153 VTAIL.n38 VSUBS 0.013741f
C154 VTAIL.n39 VSUBS 0.030674f
C155 VTAIL.n40 VSUBS 0.030674f
C156 VTAIL.n41 VSUBS 0.013741f
C157 VTAIL.n42 VSUBS 0.012977f
C158 VTAIL.n43 VSUBS 0.02415f
C159 VTAIL.n44 VSUBS 0.02415f
C160 VTAIL.n45 VSUBS 0.012977f
C161 VTAIL.n46 VSUBS 0.013741f
C162 VTAIL.n47 VSUBS 0.030674f
C163 VTAIL.n48 VSUBS 0.030674f
C164 VTAIL.n49 VSUBS 0.013741f
C165 VTAIL.n50 VSUBS 0.012977f
C166 VTAIL.n51 VSUBS 0.02415f
C167 VTAIL.n52 VSUBS 0.02415f
C168 VTAIL.n53 VSUBS 0.012977f
C169 VTAIL.n54 VSUBS 0.013741f
C170 VTAIL.n55 VSUBS 0.030674f
C171 VTAIL.n56 VSUBS 0.030674f
C172 VTAIL.n57 VSUBS 0.013741f
C173 VTAIL.n58 VSUBS 0.012977f
C174 VTAIL.n59 VSUBS 0.02415f
C175 VTAIL.n60 VSUBS 0.02415f
C176 VTAIL.n61 VSUBS 0.012977f
C177 VTAIL.n62 VSUBS 0.013741f
C178 VTAIL.n63 VSUBS 0.030674f
C179 VTAIL.n64 VSUBS 0.030674f
C180 VTAIL.n65 VSUBS 0.013741f
C181 VTAIL.n66 VSUBS 0.012977f
C182 VTAIL.n67 VSUBS 0.02415f
C183 VTAIL.n68 VSUBS 0.02415f
C184 VTAIL.n69 VSUBS 0.012977f
C185 VTAIL.n70 VSUBS 0.013741f
C186 VTAIL.n71 VSUBS 0.030674f
C187 VTAIL.n72 VSUBS 0.030674f
C188 VTAIL.n73 VSUBS 0.030674f
C189 VTAIL.n74 VSUBS 0.013741f
C190 VTAIL.n75 VSUBS 0.012977f
C191 VTAIL.n76 VSUBS 0.02415f
C192 VTAIL.n77 VSUBS 0.02415f
C193 VTAIL.n78 VSUBS 0.012977f
C194 VTAIL.n79 VSUBS 0.013359f
C195 VTAIL.n80 VSUBS 0.013359f
C196 VTAIL.n81 VSUBS 0.030674f
C197 VTAIL.n82 VSUBS 0.030674f
C198 VTAIL.n83 VSUBS 0.013741f
C199 VTAIL.n84 VSUBS 0.012977f
C200 VTAIL.n85 VSUBS 0.02415f
C201 VTAIL.n86 VSUBS 0.02415f
C202 VTAIL.n87 VSUBS 0.012977f
C203 VTAIL.n88 VSUBS 0.013741f
C204 VTAIL.n89 VSUBS 0.030674f
C205 VTAIL.n90 VSUBS 0.071124f
C206 VTAIL.n91 VSUBS 0.013741f
C207 VTAIL.n92 VSUBS 0.012977f
C208 VTAIL.n93 VSUBS 0.055822f
C209 VTAIL.n94 VSUBS 0.035628f
C210 VTAIL.n95 VSUBS 0.283259f
C211 VTAIL.n96 VSUBS 0.025616f
C212 VTAIL.n97 VSUBS 0.02415f
C213 VTAIL.n98 VSUBS 0.012977f
C214 VTAIL.n99 VSUBS 0.030674f
C215 VTAIL.n100 VSUBS 0.013741f
C216 VTAIL.n101 VSUBS 0.02415f
C217 VTAIL.n102 VSUBS 0.012977f
C218 VTAIL.n103 VSUBS 0.030674f
C219 VTAIL.n104 VSUBS 0.013741f
C220 VTAIL.n105 VSUBS 0.02415f
C221 VTAIL.n106 VSUBS 0.012977f
C222 VTAIL.n107 VSUBS 0.030674f
C223 VTAIL.n108 VSUBS 0.013741f
C224 VTAIL.n109 VSUBS 0.02415f
C225 VTAIL.n110 VSUBS 0.012977f
C226 VTAIL.n111 VSUBS 0.030674f
C227 VTAIL.n112 VSUBS 0.013741f
C228 VTAIL.n113 VSUBS 0.02415f
C229 VTAIL.n114 VSUBS 0.012977f
C230 VTAIL.n115 VSUBS 0.030674f
C231 VTAIL.n116 VSUBS 0.013741f
C232 VTAIL.n117 VSUBS 0.02415f
C233 VTAIL.n118 VSUBS 0.012977f
C234 VTAIL.n119 VSUBS 0.030674f
C235 VTAIL.n120 VSUBS 0.013741f
C236 VTAIL.n121 VSUBS 0.02415f
C237 VTAIL.n122 VSUBS 0.012977f
C238 VTAIL.n123 VSUBS 0.030674f
C239 VTAIL.n124 VSUBS 0.013741f
C240 VTAIL.n125 VSUBS 0.18306f
C241 VTAIL.t10 VSUBS 0.065774f
C242 VTAIL.n126 VSUBS 0.023005f
C243 VTAIL.n127 VSUBS 0.019513f
C244 VTAIL.n128 VSUBS 0.012977f
C245 VTAIL.n129 VSUBS 1.73938f
C246 VTAIL.n130 VSUBS 0.02415f
C247 VTAIL.n131 VSUBS 0.012977f
C248 VTAIL.n132 VSUBS 0.013741f
C249 VTAIL.n133 VSUBS 0.030674f
C250 VTAIL.n134 VSUBS 0.030674f
C251 VTAIL.n135 VSUBS 0.013741f
C252 VTAIL.n136 VSUBS 0.012977f
C253 VTAIL.n137 VSUBS 0.02415f
C254 VTAIL.n138 VSUBS 0.02415f
C255 VTAIL.n139 VSUBS 0.012977f
C256 VTAIL.n140 VSUBS 0.013741f
C257 VTAIL.n141 VSUBS 0.030674f
C258 VTAIL.n142 VSUBS 0.030674f
C259 VTAIL.n143 VSUBS 0.013741f
C260 VTAIL.n144 VSUBS 0.012977f
C261 VTAIL.n145 VSUBS 0.02415f
C262 VTAIL.n146 VSUBS 0.02415f
C263 VTAIL.n147 VSUBS 0.012977f
C264 VTAIL.n148 VSUBS 0.013741f
C265 VTAIL.n149 VSUBS 0.030674f
C266 VTAIL.n150 VSUBS 0.030674f
C267 VTAIL.n151 VSUBS 0.013741f
C268 VTAIL.n152 VSUBS 0.012977f
C269 VTAIL.n153 VSUBS 0.02415f
C270 VTAIL.n154 VSUBS 0.02415f
C271 VTAIL.n155 VSUBS 0.012977f
C272 VTAIL.n156 VSUBS 0.013741f
C273 VTAIL.n157 VSUBS 0.030674f
C274 VTAIL.n158 VSUBS 0.030674f
C275 VTAIL.n159 VSUBS 0.013741f
C276 VTAIL.n160 VSUBS 0.012977f
C277 VTAIL.n161 VSUBS 0.02415f
C278 VTAIL.n162 VSUBS 0.02415f
C279 VTAIL.n163 VSUBS 0.012977f
C280 VTAIL.n164 VSUBS 0.013741f
C281 VTAIL.n165 VSUBS 0.030674f
C282 VTAIL.n166 VSUBS 0.030674f
C283 VTAIL.n167 VSUBS 0.030674f
C284 VTAIL.n168 VSUBS 0.013741f
C285 VTAIL.n169 VSUBS 0.012977f
C286 VTAIL.n170 VSUBS 0.02415f
C287 VTAIL.n171 VSUBS 0.02415f
C288 VTAIL.n172 VSUBS 0.012977f
C289 VTAIL.n173 VSUBS 0.013359f
C290 VTAIL.n174 VSUBS 0.013359f
C291 VTAIL.n175 VSUBS 0.030674f
C292 VTAIL.n176 VSUBS 0.030674f
C293 VTAIL.n177 VSUBS 0.013741f
C294 VTAIL.n178 VSUBS 0.012977f
C295 VTAIL.n179 VSUBS 0.02415f
C296 VTAIL.n180 VSUBS 0.02415f
C297 VTAIL.n181 VSUBS 0.012977f
C298 VTAIL.n182 VSUBS 0.013741f
C299 VTAIL.n183 VSUBS 0.030674f
C300 VTAIL.n184 VSUBS 0.071124f
C301 VTAIL.n185 VSUBS 0.013741f
C302 VTAIL.n186 VSUBS 0.012977f
C303 VTAIL.n187 VSUBS 0.055822f
C304 VTAIL.n188 VSUBS 0.035628f
C305 VTAIL.n189 VSUBS 0.283259f
C306 VTAIL.t9 VSUBS 0.320615f
C307 VTAIL.t11 VSUBS 0.320615f
C308 VTAIL.n190 VSUBS 2.49217f
C309 VTAIL.n191 VSUBS 1.0393f
C310 VTAIL.n192 VSUBS 0.025616f
C311 VTAIL.n193 VSUBS 0.02415f
C312 VTAIL.n194 VSUBS 0.012977f
C313 VTAIL.n195 VSUBS 0.030674f
C314 VTAIL.n196 VSUBS 0.013741f
C315 VTAIL.n197 VSUBS 0.02415f
C316 VTAIL.n198 VSUBS 0.012977f
C317 VTAIL.n199 VSUBS 0.030674f
C318 VTAIL.n200 VSUBS 0.013741f
C319 VTAIL.n201 VSUBS 0.02415f
C320 VTAIL.n202 VSUBS 0.012977f
C321 VTAIL.n203 VSUBS 0.030674f
C322 VTAIL.n204 VSUBS 0.013741f
C323 VTAIL.n205 VSUBS 0.02415f
C324 VTAIL.n206 VSUBS 0.012977f
C325 VTAIL.n207 VSUBS 0.030674f
C326 VTAIL.n208 VSUBS 0.013741f
C327 VTAIL.n209 VSUBS 0.02415f
C328 VTAIL.n210 VSUBS 0.012977f
C329 VTAIL.n211 VSUBS 0.030674f
C330 VTAIL.n212 VSUBS 0.013741f
C331 VTAIL.n213 VSUBS 0.02415f
C332 VTAIL.n214 VSUBS 0.012977f
C333 VTAIL.n215 VSUBS 0.030674f
C334 VTAIL.n216 VSUBS 0.013741f
C335 VTAIL.n217 VSUBS 0.02415f
C336 VTAIL.n218 VSUBS 0.012977f
C337 VTAIL.n219 VSUBS 0.030674f
C338 VTAIL.n220 VSUBS 0.013741f
C339 VTAIL.n221 VSUBS 0.18306f
C340 VTAIL.t12 VSUBS 0.065774f
C341 VTAIL.n222 VSUBS 0.023005f
C342 VTAIL.n223 VSUBS 0.019513f
C343 VTAIL.n224 VSUBS 0.012977f
C344 VTAIL.n225 VSUBS 1.73938f
C345 VTAIL.n226 VSUBS 0.02415f
C346 VTAIL.n227 VSUBS 0.012977f
C347 VTAIL.n228 VSUBS 0.013741f
C348 VTAIL.n229 VSUBS 0.030674f
C349 VTAIL.n230 VSUBS 0.030674f
C350 VTAIL.n231 VSUBS 0.013741f
C351 VTAIL.n232 VSUBS 0.012977f
C352 VTAIL.n233 VSUBS 0.02415f
C353 VTAIL.n234 VSUBS 0.02415f
C354 VTAIL.n235 VSUBS 0.012977f
C355 VTAIL.n236 VSUBS 0.013741f
C356 VTAIL.n237 VSUBS 0.030674f
C357 VTAIL.n238 VSUBS 0.030674f
C358 VTAIL.n239 VSUBS 0.013741f
C359 VTAIL.n240 VSUBS 0.012977f
C360 VTAIL.n241 VSUBS 0.02415f
C361 VTAIL.n242 VSUBS 0.02415f
C362 VTAIL.n243 VSUBS 0.012977f
C363 VTAIL.n244 VSUBS 0.013741f
C364 VTAIL.n245 VSUBS 0.030674f
C365 VTAIL.n246 VSUBS 0.030674f
C366 VTAIL.n247 VSUBS 0.013741f
C367 VTAIL.n248 VSUBS 0.012977f
C368 VTAIL.n249 VSUBS 0.02415f
C369 VTAIL.n250 VSUBS 0.02415f
C370 VTAIL.n251 VSUBS 0.012977f
C371 VTAIL.n252 VSUBS 0.013741f
C372 VTAIL.n253 VSUBS 0.030674f
C373 VTAIL.n254 VSUBS 0.030674f
C374 VTAIL.n255 VSUBS 0.013741f
C375 VTAIL.n256 VSUBS 0.012977f
C376 VTAIL.n257 VSUBS 0.02415f
C377 VTAIL.n258 VSUBS 0.02415f
C378 VTAIL.n259 VSUBS 0.012977f
C379 VTAIL.n260 VSUBS 0.013741f
C380 VTAIL.n261 VSUBS 0.030674f
C381 VTAIL.n262 VSUBS 0.030674f
C382 VTAIL.n263 VSUBS 0.030674f
C383 VTAIL.n264 VSUBS 0.013741f
C384 VTAIL.n265 VSUBS 0.012977f
C385 VTAIL.n266 VSUBS 0.02415f
C386 VTAIL.n267 VSUBS 0.02415f
C387 VTAIL.n268 VSUBS 0.012977f
C388 VTAIL.n269 VSUBS 0.013359f
C389 VTAIL.n270 VSUBS 0.013359f
C390 VTAIL.n271 VSUBS 0.030674f
C391 VTAIL.n272 VSUBS 0.030674f
C392 VTAIL.n273 VSUBS 0.013741f
C393 VTAIL.n274 VSUBS 0.012977f
C394 VTAIL.n275 VSUBS 0.02415f
C395 VTAIL.n276 VSUBS 0.02415f
C396 VTAIL.n277 VSUBS 0.012977f
C397 VTAIL.n278 VSUBS 0.013741f
C398 VTAIL.n279 VSUBS 0.030674f
C399 VTAIL.n280 VSUBS 0.071124f
C400 VTAIL.n281 VSUBS 0.013741f
C401 VTAIL.n282 VSUBS 0.012977f
C402 VTAIL.n283 VSUBS 0.055822f
C403 VTAIL.n284 VSUBS 0.035628f
C404 VTAIL.n285 VSUBS 1.92783f
C405 VTAIL.n286 VSUBS 0.025616f
C406 VTAIL.n287 VSUBS 0.02415f
C407 VTAIL.n288 VSUBS 0.012977f
C408 VTAIL.n289 VSUBS 0.030674f
C409 VTAIL.n290 VSUBS 0.013741f
C410 VTAIL.n291 VSUBS 0.02415f
C411 VTAIL.n292 VSUBS 0.012977f
C412 VTAIL.n293 VSUBS 0.030674f
C413 VTAIL.n294 VSUBS 0.013741f
C414 VTAIL.n295 VSUBS 0.02415f
C415 VTAIL.n296 VSUBS 0.012977f
C416 VTAIL.n297 VSUBS 0.030674f
C417 VTAIL.n298 VSUBS 0.030674f
C418 VTAIL.n299 VSUBS 0.013741f
C419 VTAIL.n300 VSUBS 0.02415f
C420 VTAIL.n301 VSUBS 0.012977f
C421 VTAIL.n302 VSUBS 0.030674f
C422 VTAIL.n303 VSUBS 0.013741f
C423 VTAIL.n304 VSUBS 0.02415f
C424 VTAIL.n305 VSUBS 0.012977f
C425 VTAIL.n306 VSUBS 0.030674f
C426 VTAIL.n307 VSUBS 0.013741f
C427 VTAIL.n308 VSUBS 0.02415f
C428 VTAIL.n309 VSUBS 0.012977f
C429 VTAIL.n310 VSUBS 0.030674f
C430 VTAIL.n311 VSUBS 0.013741f
C431 VTAIL.n312 VSUBS 0.02415f
C432 VTAIL.n313 VSUBS 0.012977f
C433 VTAIL.n314 VSUBS 0.030674f
C434 VTAIL.n315 VSUBS 0.013741f
C435 VTAIL.n316 VSUBS 0.18306f
C436 VTAIL.t7 VSUBS 0.065774f
C437 VTAIL.n317 VSUBS 0.023005f
C438 VTAIL.n318 VSUBS 0.019513f
C439 VTAIL.n319 VSUBS 0.012977f
C440 VTAIL.n320 VSUBS 1.73938f
C441 VTAIL.n321 VSUBS 0.02415f
C442 VTAIL.n322 VSUBS 0.012977f
C443 VTAIL.n323 VSUBS 0.013741f
C444 VTAIL.n324 VSUBS 0.030674f
C445 VTAIL.n325 VSUBS 0.030674f
C446 VTAIL.n326 VSUBS 0.013741f
C447 VTAIL.n327 VSUBS 0.012977f
C448 VTAIL.n328 VSUBS 0.02415f
C449 VTAIL.n329 VSUBS 0.02415f
C450 VTAIL.n330 VSUBS 0.012977f
C451 VTAIL.n331 VSUBS 0.013741f
C452 VTAIL.n332 VSUBS 0.030674f
C453 VTAIL.n333 VSUBS 0.030674f
C454 VTAIL.n334 VSUBS 0.013741f
C455 VTAIL.n335 VSUBS 0.012977f
C456 VTAIL.n336 VSUBS 0.02415f
C457 VTAIL.n337 VSUBS 0.02415f
C458 VTAIL.n338 VSUBS 0.012977f
C459 VTAIL.n339 VSUBS 0.013741f
C460 VTAIL.n340 VSUBS 0.030674f
C461 VTAIL.n341 VSUBS 0.030674f
C462 VTAIL.n342 VSUBS 0.013741f
C463 VTAIL.n343 VSUBS 0.012977f
C464 VTAIL.n344 VSUBS 0.02415f
C465 VTAIL.n345 VSUBS 0.02415f
C466 VTAIL.n346 VSUBS 0.012977f
C467 VTAIL.n347 VSUBS 0.013741f
C468 VTAIL.n348 VSUBS 0.030674f
C469 VTAIL.n349 VSUBS 0.030674f
C470 VTAIL.n350 VSUBS 0.013741f
C471 VTAIL.n351 VSUBS 0.012977f
C472 VTAIL.n352 VSUBS 0.02415f
C473 VTAIL.n353 VSUBS 0.02415f
C474 VTAIL.n354 VSUBS 0.012977f
C475 VTAIL.n355 VSUBS 0.013741f
C476 VTAIL.n356 VSUBS 0.030674f
C477 VTAIL.n357 VSUBS 0.030674f
C478 VTAIL.n358 VSUBS 0.013741f
C479 VTAIL.n359 VSUBS 0.012977f
C480 VTAIL.n360 VSUBS 0.02415f
C481 VTAIL.n361 VSUBS 0.02415f
C482 VTAIL.n362 VSUBS 0.012977f
C483 VTAIL.n363 VSUBS 0.013359f
C484 VTAIL.n364 VSUBS 0.013359f
C485 VTAIL.n365 VSUBS 0.030674f
C486 VTAIL.n366 VSUBS 0.030674f
C487 VTAIL.n367 VSUBS 0.013741f
C488 VTAIL.n368 VSUBS 0.012977f
C489 VTAIL.n369 VSUBS 0.02415f
C490 VTAIL.n370 VSUBS 0.02415f
C491 VTAIL.n371 VSUBS 0.012977f
C492 VTAIL.n372 VSUBS 0.013741f
C493 VTAIL.n373 VSUBS 0.030674f
C494 VTAIL.n374 VSUBS 0.071124f
C495 VTAIL.n375 VSUBS 0.013741f
C496 VTAIL.n376 VSUBS 0.012977f
C497 VTAIL.n377 VSUBS 0.055822f
C498 VTAIL.n378 VSUBS 0.035628f
C499 VTAIL.n379 VSUBS 1.92783f
C500 VTAIL.t0 VSUBS 0.320615f
C501 VTAIL.t6 VSUBS 0.320615f
C502 VTAIL.n380 VSUBS 2.49219f
C503 VTAIL.n381 VSUBS 1.03928f
C504 VTAIL.n382 VSUBS 0.025616f
C505 VTAIL.n383 VSUBS 0.02415f
C506 VTAIL.n384 VSUBS 0.012977f
C507 VTAIL.n385 VSUBS 0.030674f
C508 VTAIL.n386 VSUBS 0.013741f
C509 VTAIL.n387 VSUBS 0.02415f
C510 VTAIL.n388 VSUBS 0.012977f
C511 VTAIL.n389 VSUBS 0.030674f
C512 VTAIL.n390 VSUBS 0.013741f
C513 VTAIL.n391 VSUBS 0.02415f
C514 VTAIL.n392 VSUBS 0.012977f
C515 VTAIL.n393 VSUBS 0.030674f
C516 VTAIL.n394 VSUBS 0.030674f
C517 VTAIL.n395 VSUBS 0.013741f
C518 VTAIL.n396 VSUBS 0.02415f
C519 VTAIL.n397 VSUBS 0.012977f
C520 VTAIL.n398 VSUBS 0.030674f
C521 VTAIL.n399 VSUBS 0.013741f
C522 VTAIL.n400 VSUBS 0.02415f
C523 VTAIL.n401 VSUBS 0.012977f
C524 VTAIL.n402 VSUBS 0.030674f
C525 VTAIL.n403 VSUBS 0.013741f
C526 VTAIL.n404 VSUBS 0.02415f
C527 VTAIL.n405 VSUBS 0.012977f
C528 VTAIL.n406 VSUBS 0.030674f
C529 VTAIL.n407 VSUBS 0.013741f
C530 VTAIL.n408 VSUBS 0.02415f
C531 VTAIL.n409 VSUBS 0.012977f
C532 VTAIL.n410 VSUBS 0.030674f
C533 VTAIL.n411 VSUBS 0.013741f
C534 VTAIL.n412 VSUBS 0.18306f
C535 VTAIL.t1 VSUBS 0.065774f
C536 VTAIL.n413 VSUBS 0.023005f
C537 VTAIL.n414 VSUBS 0.019513f
C538 VTAIL.n415 VSUBS 0.012977f
C539 VTAIL.n416 VSUBS 1.73938f
C540 VTAIL.n417 VSUBS 0.02415f
C541 VTAIL.n418 VSUBS 0.012977f
C542 VTAIL.n419 VSUBS 0.013741f
C543 VTAIL.n420 VSUBS 0.030674f
C544 VTAIL.n421 VSUBS 0.030674f
C545 VTAIL.n422 VSUBS 0.013741f
C546 VTAIL.n423 VSUBS 0.012977f
C547 VTAIL.n424 VSUBS 0.02415f
C548 VTAIL.n425 VSUBS 0.02415f
C549 VTAIL.n426 VSUBS 0.012977f
C550 VTAIL.n427 VSUBS 0.013741f
C551 VTAIL.n428 VSUBS 0.030674f
C552 VTAIL.n429 VSUBS 0.030674f
C553 VTAIL.n430 VSUBS 0.013741f
C554 VTAIL.n431 VSUBS 0.012977f
C555 VTAIL.n432 VSUBS 0.02415f
C556 VTAIL.n433 VSUBS 0.02415f
C557 VTAIL.n434 VSUBS 0.012977f
C558 VTAIL.n435 VSUBS 0.013741f
C559 VTAIL.n436 VSUBS 0.030674f
C560 VTAIL.n437 VSUBS 0.030674f
C561 VTAIL.n438 VSUBS 0.013741f
C562 VTAIL.n439 VSUBS 0.012977f
C563 VTAIL.n440 VSUBS 0.02415f
C564 VTAIL.n441 VSUBS 0.02415f
C565 VTAIL.n442 VSUBS 0.012977f
C566 VTAIL.n443 VSUBS 0.013741f
C567 VTAIL.n444 VSUBS 0.030674f
C568 VTAIL.n445 VSUBS 0.030674f
C569 VTAIL.n446 VSUBS 0.013741f
C570 VTAIL.n447 VSUBS 0.012977f
C571 VTAIL.n448 VSUBS 0.02415f
C572 VTAIL.n449 VSUBS 0.02415f
C573 VTAIL.n450 VSUBS 0.012977f
C574 VTAIL.n451 VSUBS 0.013741f
C575 VTAIL.n452 VSUBS 0.030674f
C576 VTAIL.n453 VSUBS 0.030674f
C577 VTAIL.n454 VSUBS 0.013741f
C578 VTAIL.n455 VSUBS 0.012977f
C579 VTAIL.n456 VSUBS 0.02415f
C580 VTAIL.n457 VSUBS 0.02415f
C581 VTAIL.n458 VSUBS 0.012977f
C582 VTAIL.n459 VSUBS 0.013359f
C583 VTAIL.n460 VSUBS 0.013359f
C584 VTAIL.n461 VSUBS 0.030674f
C585 VTAIL.n462 VSUBS 0.030674f
C586 VTAIL.n463 VSUBS 0.013741f
C587 VTAIL.n464 VSUBS 0.012977f
C588 VTAIL.n465 VSUBS 0.02415f
C589 VTAIL.n466 VSUBS 0.02415f
C590 VTAIL.n467 VSUBS 0.012977f
C591 VTAIL.n468 VSUBS 0.013741f
C592 VTAIL.n469 VSUBS 0.030674f
C593 VTAIL.n470 VSUBS 0.071124f
C594 VTAIL.n471 VSUBS 0.013741f
C595 VTAIL.n472 VSUBS 0.012977f
C596 VTAIL.n473 VSUBS 0.055822f
C597 VTAIL.n474 VSUBS 0.035628f
C598 VTAIL.n475 VSUBS 0.283259f
C599 VTAIL.n476 VSUBS 0.025616f
C600 VTAIL.n477 VSUBS 0.02415f
C601 VTAIL.n478 VSUBS 0.012977f
C602 VTAIL.n479 VSUBS 0.030674f
C603 VTAIL.n480 VSUBS 0.013741f
C604 VTAIL.n481 VSUBS 0.02415f
C605 VTAIL.n482 VSUBS 0.012977f
C606 VTAIL.n483 VSUBS 0.030674f
C607 VTAIL.n484 VSUBS 0.013741f
C608 VTAIL.n485 VSUBS 0.02415f
C609 VTAIL.n486 VSUBS 0.012977f
C610 VTAIL.n487 VSUBS 0.030674f
C611 VTAIL.n488 VSUBS 0.030674f
C612 VTAIL.n489 VSUBS 0.013741f
C613 VTAIL.n490 VSUBS 0.02415f
C614 VTAIL.n491 VSUBS 0.012977f
C615 VTAIL.n492 VSUBS 0.030674f
C616 VTAIL.n493 VSUBS 0.013741f
C617 VTAIL.n494 VSUBS 0.02415f
C618 VTAIL.n495 VSUBS 0.012977f
C619 VTAIL.n496 VSUBS 0.030674f
C620 VTAIL.n497 VSUBS 0.013741f
C621 VTAIL.n498 VSUBS 0.02415f
C622 VTAIL.n499 VSUBS 0.012977f
C623 VTAIL.n500 VSUBS 0.030674f
C624 VTAIL.n501 VSUBS 0.013741f
C625 VTAIL.n502 VSUBS 0.02415f
C626 VTAIL.n503 VSUBS 0.012977f
C627 VTAIL.n504 VSUBS 0.030674f
C628 VTAIL.n505 VSUBS 0.013741f
C629 VTAIL.n506 VSUBS 0.18306f
C630 VTAIL.t8 VSUBS 0.065774f
C631 VTAIL.n507 VSUBS 0.023005f
C632 VTAIL.n508 VSUBS 0.019513f
C633 VTAIL.n509 VSUBS 0.012977f
C634 VTAIL.n510 VSUBS 1.73938f
C635 VTAIL.n511 VSUBS 0.02415f
C636 VTAIL.n512 VSUBS 0.012977f
C637 VTAIL.n513 VSUBS 0.013741f
C638 VTAIL.n514 VSUBS 0.030674f
C639 VTAIL.n515 VSUBS 0.030674f
C640 VTAIL.n516 VSUBS 0.013741f
C641 VTAIL.n517 VSUBS 0.012977f
C642 VTAIL.n518 VSUBS 0.02415f
C643 VTAIL.n519 VSUBS 0.02415f
C644 VTAIL.n520 VSUBS 0.012977f
C645 VTAIL.n521 VSUBS 0.013741f
C646 VTAIL.n522 VSUBS 0.030674f
C647 VTAIL.n523 VSUBS 0.030674f
C648 VTAIL.n524 VSUBS 0.013741f
C649 VTAIL.n525 VSUBS 0.012977f
C650 VTAIL.n526 VSUBS 0.02415f
C651 VTAIL.n527 VSUBS 0.02415f
C652 VTAIL.n528 VSUBS 0.012977f
C653 VTAIL.n529 VSUBS 0.013741f
C654 VTAIL.n530 VSUBS 0.030674f
C655 VTAIL.n531 VSUBS 0.030674f
C656 VTAIL.n532 VSUBS 0.013741f
C657 VTAIL.n533 VSUBS 0.012977f
C658 VTAIL.n534 VSUBS 0.02415f
C659 VTAIL.n535 VSUBS 0.02415f
C660 VTAIL.n536 VSUBS 0.012977f
C661 VTAIL.n537 VSUBS 0.013741f
C662 VTAIL.n538 VSUBS 0.030674f
C663 VTAIL.n539 VSUBS 0.030674f
C664 VTAIL.n540 VSUBS 0.013741f
C665 VTAIL.n541 VSUBS 0.012977f
C666 VTAIL.n542 VSUBS 0.02415f
C667 VTAIL.n543 VSUBS 0.02415f
C668 VTAIL.n544 VSUBS 0.012977f
C669 VTAIL.n545 VSUBS 0.013741f
C670 VTAIL.n546 VSUBS 0.030674f
C671 VTAIL.n547 VSUBS 0.030674f
C672 VTAIL.n548 VSUBS 0.013741f
C673 VTAIL.n549 VSUBS 0.012977f
C674 VTAIL.n550 VSUBS 0.02415f
C675 VTAIL.n551 VSUBS 0.02415f
C676 VTAIL.n552 VSUBS 0.012977f
C677 VTAIL.n553 VSUBS 0.013359f
C678 VTAIL.n554 VSUBS 0.013359f
C679 VTAIL.n555 VSUBS 0.030674f
C680 VTAIL.n556 VSUBS 0.030674f
C681 VTAIL.n557 VSUBS 0.013741f
C682 VTAIL.n558 VSUBS 0.012977f
C683 VTAIL.n559 VSUBS 0.02415f
C684 VTAIL.n560 VSUBS 0.02415f
C685 VTAIL.n561 VSUBS 0.012977f
C686 VTAIL.n562 VSUBS 0.013741f
C687 VTAIL.n563 VSUBS 0.030674f
C688 VTAIL.n564 VSUBS 0.071124f
C689 VTAIL.n565 VSUBS 0.013741f
C690 VTAIL.n566 VSUBS 0.012977f
C691 VTAIL.n567 VSUBS 0.055822f
C692 VTAIL.n568 VSUBS 0.035628f
C693 VTAIL.n569 VSUBS 0.283259f
C694 VTAIL.t14 VSUBS 0.320615f
C695 VTAIL.t15 VSUBS 0.320615f
C696 VTAIL.n570 VSUBS 2.49219f
C697 VTAIL.n571 VSUBS 1.03928f
C698 VTAIL.n572 VSUBS 0.025616f
C699 VTAIL.n573 VSUBS 0.02415f
C700 VTAIL.n574 VSUBS 0.012977f
C701 VTAIL.n575 VSUBS 0.030674f
C702 VTAIL.n576 VSUBS 0.013741f
C703 VTAIL.n577 VSUBS 0.02415f
C704 VTAIL.n578 VSUBS 0.012977f
C705 VTAIL.n579 VSUBS 0.030674f
C706 VTAIL.n580 VSUBS 0.013741f
C707 VTAIL.n581 VSUBS 0.02415f
C708 VTAIL.n582 VSUBS 0.012977f
C709 VTAIL.n583 VSUBS 0.030674f
C710 VTAIL.n584 VSUBS 0.030674f
C711 VTAIL.n585 VSUBS 0.013741f
C712 VTAIL.n586 VSUBS 0.02415f
C713 VTAIL.n587 VSUBS 0.012977f
C714 VTAIL.n588 VSUBS 0.030674f
C715 VTAIL.n589 VSUBS 0.013741f
C716 VTAIL.n590 VSUBS 0.02415f
C717 VTAIL.n591 VSUBS 0.012977f
C718 VTAIL.n592 VSUBS 0.030674f
C719 VTAIL.n593 VSUBS 0.013741f
C720 VTAIL.n594 VSUBS 0.02415f
C721 VTAIL.n595 VSUBS 0.012977f
C722 VTAIL.n596 VSUBS 0.030674f
C723 VTAIL.n597 VSUBS 0.013741f
C724 VTAIL.n598 VSUBS 0.02415f
C725 VTAIL.n599 VSUBS 0.012977f
C726 VTAIL.n600 VSUBS 0.030674f
C727 VTAIL.n601 VSUBS 0.013741f
C728 VTAIL.n602 VSUBS 0.18306f
C729 VTAIL.t13 VSUBS 0.065774f
C730 VTAIL.n603 VSUBS 0.023005f
C731 VTAIL.n604 VSUBS 0.019513f
C732 VTAIL.n605 VSUBS 0.012977f
C733 VTAIL.n606 VSUBS 1.73938f
C734 VTAIL.n607 VSUBS 0.02415f
C735 VTAIL.n608 VSUBS 0.012977f
C736 VTAIL.n609 VSUBS 0.013741f
C737 VTAIL.n610 VSUBS 0.030674f
C738 VTAIL.n611 VSUBS 0.030674f
C739 VTAIL.n612 VSUBS 0.013741f
C740 VTAIL.n613 VSUBS 0.012977f
C741 VTAIL.n614 VSUBS 0.02415f
C742 VTAIL.n615 VSUBS 0.02415f
C743 VTAIL.n616 VSUBS 0.012977f
C744 VTAIL.n617 VSUBS 0.013741f
C745 VTAIL.n618 VSUBS 0.030674f
C746 VTAIL.n619 VSUBS 0.030674f
C747 VTAIL.n620 VSUBS 0.013741f
C748 VTAIL.n621 VSUBS 0.012977f
C749 VTAIL.n622 VSUBS 0.02415f
C750 VTAIL.n623 VSUBS 0.02415f
C751 VTAIL.n624 VSUBS 0.012977f
C752 VTAIL.n625 VSUBS 0.013741f
C753 VTAIL.n626 VSUBS 0.030674f
C754 VTAIL.n627 VSUBS 0.030674f
C755 VTAIL.n628 VSUBS 0.013741f
C756 VTAIL.n629 VSUBS 0.012977f
C757 VTAIL.n630 VSUBS 0.02415f
C758 VTAIL.n631 VSUBS 0.02415f
C759 VTAIL.n632 VSUBS 0.012977f
C760 VTAIL.n633 VSUBS 0.013741f
C761 VTAIL.n634 VSUBS 0.030674f
C762 VTAIL.n635 VSUBS 0.030674f
C763 VTAIL.n636 VSUBS 0.013741f
C764 VTAIL.n637 VSUBS 0.012977f
C765 VTAIL.n638 VSUBS 0.02415f
C766 VTAIL.n639 VSUBS 0.02415f
C767 VTAIL.n640 VSUBS 0.012977f
C768 VTAIL.n641 VSUBS 0.013741f
C769 VTAIL.n642 VSUBS 0.030674f
C770 VTAIL.n643 VSUBS 0.030674f
C771 VTAIL.n644 VSUBS 0.013741f
C772 VTAIL.n645 VSUBS 0.012977f
C773 VTAIL.n646 VSUBS 0.02415f
C774 VTAIL.n647 VSUBS 0.02415f
C775 VTAIL.n648 VSUBS 0.012977f
C776 VTAIL.n649 VSUBS 0.013359f
C777 VTAIL.n650 VSUBS 0.013359f
C778 VTAIL.n651 VSUBS 0.030674f
C779 VTAIL.n652 VSUBS 0.030674f
C780 VTAIL.n653 VSUBS 0.013741f
C781 VTAIL.n654 VSUBS 0.012977f
C782 VTAIL.n655 VSUBS 0.02415f
C783 VTAIL.n656 VSUBS 0.02415f
C784 VTAIL.n657 VSUBS 0.012977f
C785 VTAIL.n658 VSUBS 0.013741f
C786 VTAIL.n659 VSUBS 0.030674f
C787 VTAIL.n660 VSUBS 0.071124f
C788 VTAIL.n661 VSUBS 0.013741f
C789 VTAIL.n662 VSUBS 0.012977f
C790 VTAIL.n663 VSUBS 0.055822f
C791 VTAIL.n664 VSUBS 0.035628f
C792 VTAIL.n665 VSUBS 1.92783f
C793 VTAIL.n666 VSUBS 0.025616f
C794 VTAIL.n667 VSUBS 0.02415f
C795 VTAIL.n668 VSUBS 0.012977f
C796 VTAIL.n669 VSUBS 0.030674f
C797 VTAIL.n670 VSUBS 0.013741f
C798 VTAIL.n671 VSUBS 0.02415f
C799 VTAIL.n672 VSUBS 0.012977f
C800 VTAIL.n673 VSUBS 0.030674f
C801 VTAIL.n674 VSUBS 0.013741f
C802 VTAIL.n675 VSUBS 0.02415f
C803 VTAIL.n676 VSUBS 0.012977f
C804 VTAIL.n677 VSUBS 0.030674f
C805 VTAIL.n678 VSUBS 0.013741f
C806 VTAIL.n679 VSUBS 0.02415f
C807 VTAIL.n680 VSUBS 0.012977f
C808 VTAIL.n681 VSUBS 0.030674f
C809 VTAIL.n682 VSUBS 0.013741f
C810 VTAIL.n683 VSUBS 0.02415f
C811 VTAIL.n684 VSUBS 0.012977f
C812 VTAIL.n685 VSUBS 0.030674f
C813 VTAIL.n686 VSUBS 0.013741f
C814 VTAIL.n687 VSUBS 0.02415f
C815 VTAIL.n688 VSUBS 0.012977f
C816 VTAIL.n689 VSUBS 0.030674f
C817 VTAIL.n690 VSUBS 0.013741f
C818 VTAIL.n691 VSUBS 0.02415f
C819 VTAIL.n692 VSUBS 0.012977f
C820 VTAIL.n693 VSUBS 0.030674f
C821 VTAIL.n694 VSUBS 0.013741f
C822 VTAIL.n695 VSUBS 0.18306f
C823 VTAIL.t4 VSUBS 0.065774f
C824 VTAIL.n696 VSUBS 0.023005f
C825 VTAIL.n697 VSUBS 0.019513f
C826 VTAIL.n698 VSUBS 0.012977f
C827 VTAIL.n699 VSUBS 1.73938f
C828 VTAIL.n700 VSUBS 0.02415f
C829 VTAIL.n701 VSUBS 0.012977f
C830 VTAIL.n702 VSUBS 0.013741f
C831 VTAIL.n703 VSUBS 0.030674f
C832 VTAIL.n704 VSUBS 0.030674f
C833 VTAIL.n705 VSUBS 0.013741f
C834 VTAIL.n706 VSUBS 0.012977f
C835 VTAIL.n707 VSUBS 0.02415f
C836 VTAIL.n708 VSUBS 0.02415f
C837 VTAIL.n709 VSUBS 0.012977f
C838 VTAIL.n710 VSUBS 0.013741f
C839 VTAIL.n711 VSUBS 0.030674f
C840 VTAIL.n712 VSUBS 0.030674f
C841 VTAIL.n713 VSUBS 0.013741f
C842 VTAIL.n714 VSUBS 0.012977f
C843 VTAIL.n715 VSUBS 0.02415f
C844 VTAIL.n716 VSUBS 0.02415f
C845 VTAIL.n717 VSUBS 0.012977f
C846 VTAIL.n718 VSUBS 0.013741f
C847 VTAIL.n719 VSUBS 0.030674f
C848 VTAIL.n720 VSUBS 0.030674f
C849 VTAIL.n721 VSUBS 0.013741f
C850 VTAIL.n722 VSUBS 0.012977f
C851 VTAIL.n723 VSUBS 0.02415f
C852 VTAIL.n724 VSUBS 0.02415f
C853 VTAIL.n725 VSUBS 0.012977f
C854 VTAIL.n726 VSUBS 0.013741f
C855 VTAIL.n727 VSUBS 0.030674f
C856 VTAIL.n728 VSUBS 0.030674f
C857 VTAIL.n729 VSUBS 0.013741f
C858 VTAIL.n730 VSUBS 0.012977f
C859 VTAIL.n731 VSUBS 0.02415f
C860 VTAIL.n732 VSUBS 0.02415f
C861 VTAIL.n733 VSUBS 0.012977f
C862 VTAIL.n734 VSUBS 0.013741f
C863 VTAIL.n735 VSUBS 0.030674f
C864 VTAIL.n736 VSUBS 0.030674f
C865 VTAIL.n737 VSUBS 0.030674f
C866 VTAIL.n738 VSUBS 0.013741f
C867 VTAIL.n739 VSUBS 0.012977f
C868 VTAIL.n740 VSUBS 0.02415f
C869 VTAIL.n741 VSUBS 0.02415f
C870 VTAIL.n742 VSUBS 0.012977f
C871 VTAIL.n743 VSUBS 0.013359f
C872 VTAIL.n744 VSUBS 0.013359f
C873 VTAIL.n745 VSUBS 0.030674f
C874 VTAIL.n746 VSUBS 0.030674f
C875 VTAIL.n747 VSUBS 0.013741f
C876 VTAIL.n748 VSUBS 0.012977f
C877 VTAIL.n749 VSUBS 0.02415f
C878 VTAIL.n750 VSUBS 0.02415f
C879 VTAIL.n751 VSUBS 0.012977f
C880 VTAIL.n752 VSUBS 0.013741f
C881 VTAIL.n753 VSUBS 0.030674f
C882 VTAIL.n754 VSUBS 0.071124f
C883 VTAIL.n755 VSUBS 0.013741f
C884 VTAIL.n756 VSUBS 0.012977f
C885 VTAIL.n757 VSUBS 0.055822f
C886 VTAIL.n758 VSUBS 0.035628f
C887 VTAIL.n759 VSUBS 1.92331f
C888 VDD1.t7 VSUBS 0.386399f
C889 VDD1.t4 VSUBS 0.386399f
C890 VDD1.n0 VSUBS 3.20299f
C891 VDD1.t0 VSUBS 0.386399f
C892 VDD1.t5 VSUBS 0.386399f
C893 VDD1.n1 VSUBS 3.20121f
C894 VDD1.t2 VSUBS 0.386399f
C895 VDD1.t3 VSUBS 0.386399f
C896 VDD1.n2 VSUBS 3.20121f
C897 VDD1.n3 VSUBS 5.17507f
C898 VDD1.t6 VSUBS 0.386399f
C899 VDD1.t1 VSUBS 0.386399f
C900 VDD1.n4 VSUBS 3.18178f
C901 VDD1.n5 VSUBS 4.40051f
C902 VP.t5 VSUBS 3.67193f
C903 VP.n0 VSUBS 1.36811f
C904 VP.n1 VSUBS 0.026174f
C905 VP.n2 VSUBS 0.026375f
C906 VP.n3 VSUBS 0.026174f
C907 VP.t4 VSUBS 3.67193f
C908 VP.n4 VSUBS 1.27271f
C909 VP.n5 VSUBS 0.026174f
C910 VP.n6 VSUBS 0.038048f
C911 VP.n7 VSUBS 0.026174f
C912 VP.t6 VSUBS 3.67193f
C913 VP.n8 VSUBS 0.048538f
C914 VP.n9 VSUBS 0.026174f
C915 VP.n10 VSUBS 0.048538f
C916 VP.t2 VSUBS 3.67193f
C917 VP.n11 VSUBS 1.36811f
C918 VP.n12 VSUBS 0.026174f
C919 VP.n13 VSUBS 0.026375f
C920 VP.n14 VSUBS 0.026174f
C921 VP.t0 VSUBS 3.67193f
C922 VP.n15 VSUBS 1.27271f
C923 VP.n16 VSUBS 0.026174f
C924 VP.n17 VSUBS 0.038048f
C925 VP.n18 VSUBS 0.298994f
C926 VP.t1 VSUBS 3.67193f
C927 VP.t7 VSUBS 3.96102f
C928 VP.n19 VSUBS 1.30887f
C929 VP.n20 VSUBS 1.36559f
C930 VP.n21 VSUBS 0.045423f
C931 VP.n22 VSUBS 0.048538f
C932 VP.n23 VSUBS 0.026174f
C933 VP.n24 VSUBS 0.026174f
C934 VP.n25 VSUBS 0.026174f
C935 VP.n26 VSUBS 0.038048f
C936 VP.n27 VSUBS 0.048538f
C937 VP.n28 VSUBS 0.045423f
C938 VP.n29 VSUBS 0.026174f
C939 VP.n30 VSUBS 0.026174f
C940 VP.n31 VSUBS 0.027691f
C941 VP.n32 VSUBS 0.048538f
C942 VP.n33 VSUBS 0.051496f
C943 VP.n34 VSUBS 0.026174f
C944 VP.n35 VSUBS 0.026174f
C945 VP.n36 VSUBS 0.026174f
C946 VP.n37 VSUBS 0.046763f
C947 VP.n38 VSUBS 0.048538f
C948 VP.n39 VSUBS 0.039193f
C949 VP.n40 VSUBS 0.042238f
C950 VP.n41 VSUBS 1.76784f
C951 VP.n42 VSUBS 1.7845f
C952 VP.t3 VSUBS 3.67193f
C953 VP.n43 VSUBS 1.36811f
C954 VP.n44 VSUBS 0.039193f
C955 VP.n45 VSUBS 0.042238f
C956 VP.n46 VSUBS 0.026174f
C957 VP.n47 VSUBS 0.026174f
C958 VP.n48 VSUBS 0.046763f
C959 VP.n49 VSUBS 0.026375f
C960 VP.n50 VSUBS 0.051496f
C961 VP.n51 VSUBS 0.026174f
C962 VP.n52 VSUBS 0.026174f
C963 VP.n53 VSUBS 0.026174f
C964 VP.n54 VSUBS 0.027691f
C965 VP.n55 VSUBS 1.27271f
C966 VP.n56 VSUBS 0.045423f
C967 VP.n57 VSUBS 0.048538f
C968 VP.n58 VSUBS 0.026174f
C969 VP.n59 VSUBS 0.026174f
C970 VP.n60 VSUBS 0.026174f
C971 VP.n61 VSUBS 0.038048f
C972 VP.n62 VSUBS 0.048538f
C973 VP.n63 VSUBS 0.045423f
C974 VP.n64 VSUBS 0.026174f
C975 VP.n65 VSUBS 0.026174f
C976 VP.n66 VSUBS 0.027691f
C977 VP.n67 VSUBS 0.048538f
C978 VP.n68 VSUBS 0.051496f
C979 VP.n69 VSUBS 0.026174f
C980 VP.n70 VSUBS 0.026174f
C981 VP.n71 VSUBS 0.026174f
C982 VP.n72 VSUBS 0.046763f
C983 VP.n73 VSUBS 0.048538f
C984 VP.n74 VSUBS 0.039193f
C985 VP.n75 VSUBS 0.042238f
C986 VP.n76 VSUBS 0.060252f
C987 B.n0 VSUBS 0.006421f
C988 B.n1 VSUBS 0.006421f
C989 B.n2 VSUBS 0.009496f
C990 B.n3 VSUBS 0.007277f
C991 B.n4 VSUBS 0.007277f
C992 B.n5 VSUBS 0.007277f
C993 B.n6 VSUBS 0.007277f
C994 B.n7 VSUBS 0.007277f
C995 B.n8 VSUBS 0.007277f
C996 B.n9 VSUBS 0.007277f
C997 B.n10 VSUBS 0.007277f
C998 B.n11 VSUBS 0.007277f
C999 B.n12 VSUBS 0.007277f
C1000 B.n13 VSUBS 0.007277f
C1001 B.n14 VSUBS 0.007277f
C1002 B.n15 VSUBS 0.007277f
C1003 B.n16 VSUBS 0.007277f
C1004 B.n17 VSUBS 0.007277f
C1005 B.n18 VSUBS 0.007277f
C1006 B.n19 VSUBS 0.007277f
C1007 B.n20 VSUBS 0.007277f
C1008 B.n21 VSUBS 0.007277f
C1009 B.n22 VSUBS 0.007277f
C1010 B.n23 VSUBS 0.007277f
C1011 B.n24 VSUBS 0.007277f
C1012 B.n25 VSUBS 0.007277f
C1013 B.n26 VSUBS 0.007277f
C1014 B.n27 VSUBS 0.007277f
C1015 B.n28 VSUBS 0.007277f
C1016 B.n29 VSUBS 0.007277f
C1017 B.n30 VSUBS 0.017171f
C1018 B.n31 VSUBS 0.007277f
C1019 B.n32 VSUBS 0.007277f
C1020 B.n33 VSUBS 0.007277f
C1021 B.n34 VSUBS 0.007277f
C1022 B.n35 VSUBS 0.007277f
C1023 B.n36 VSUBS 0.007277f
C1024 B.n37 VSUBS 0.007277f
C1025 B.n38 VSUBS 0.007277f
C1026 B.n39 VSUBS 0.007277f
C1027 B.n40 VSUBS 0.007277f
C1028 B.n41 VSUBS 0.007277f
C1029 B.n42 VSUBS 0.007277f
C1030 B.n43 VSUBS 0.007277f
C1031 B.n44 VSUBS 0.007277f
C1032 B.n45 VSUBS 0.007277f
C1033 B.n46 VSUBS 0.007277f
C1034 B.n47 VSUBS 0.007277f
C1035 B.n48 VSUBS 0.007277f
C1036 B.n49 VSUBS 0.007277f
C1037 B.n50 VSUBS 0.007277f
C1038 B.n51 VSUBS 0.007277f
C1039 B.n52 VSUBS 0.007277f
C1040 B.n53 VSUBS 0.007277f
C1041 B.n54 VSUBS 0.007277f
C1042 B.n55 VSUBS 0.007277f
C1043 B.n56 VSUBS 0.007277f
C1044 B.n57 VSUBS 0.007277f
C1045 B.n58 VSUBS 0.00503f
C1046 B.n59 VSUBS 0.007277f
C1047 B.t1 VSUBS 0.334914f
C1048 B.t2 VSUBS 0.374345f
C1049 B.t0 VSUBS 2.39297f
C1050 B.n60 VSUBS 0.586561f
C1051 B.n61 VSUBS 0.328563f
C1052 B.n62 VSUBS 0.01686f
C1053 B.n63 VSUBS 0.007277f
C1054 B.n64 VSUBS 0.007277f
C1055 B.n65 VSUBS 0.007277f
C1056 B.n66 VSUBS 0.007277f
C1057 B.t7 VSUBS 0.334918f
C1058 B.t8 VSUBS 0.374348f
C1059 B.t6 VSUBS 2.39297f
C1060 B.n67 VSUBS 0.586557f
C1061 B.n68 VSUBS 0.32856f
C1062 B.n69 VSUBS 0.007277f
C1063 B.n70 VSUBS 0.007277f
C1064 B.n71 VSUBS 0.007277f
C1065 B.n72 VSUBS 0.007277f
C1066 B.n73 VSUBS 0.007277f
C1067 B.n74 VSUBS 0.007277f
C1068 B.n75 VSUBS 0.007277f
C1069 B.n76 VSUBS 0.007277f
C1070 B.n77 VSUBS 0.007277f
C1071 B.n78 VSUBS 0.007277f
C1072 B.n79 VSUBS 0.007277f
C1073 B.n80 VSUBS 0.007277f
C1074 B.n81 VSUBS 0.007277f
C1075 B.n82 VSUBS 0.007277f
C1076 B.n83 VSUBS 0.007277f
C1077 B.n84 VSUBS 0.007277f
C1078 B.n85 VSUBS 0.007277f
C1079 B.n86 VSUBS 0.007277f
C1080 B.n87 VSUBS 0.007277f
C1081 B.n88 VSUBS 0.007277f
C1082 B.n89 VSUBS 0.007277f
C1083 B.n90 VSUBS 0.007277f
C1084 B.n91 VSUBS 0.007277f
C1085 B.n92 VSUBS 0.007277f
C1086 B.n93 VSUBS 0.007277f
C1087 B.n94 VSUBS 0.007277f
C1088 B.n95 VSUBS 0.007277f
C1089 B.n96 VSUBS 0.017171f
C1090 B.n97 VSUBS 0.007277f
C1091 B.n98 VSUBS 0.007277f
C1092 B.n99 VSUBS 0.007277f
C1093 B.n100 VSUBS 0.007277f
C1094 B.n101 VSUBS 0.007277f
C1095 B.n102 VSUBS 0.007277f
C1096 B.n103 VSUBS 0.007277f
C1097 B.n104 VSUBS 0.007277f
C1098 B.n105 VSUBS 0.007277f
C1099 B.n106 VSUBS 0.007277f
C1100 B.n107 VSUBS 0.007277f
C1101 B.n108 VSUBS 0.007277f
C1102 B.n109 VSUBS 0.007277f
C1103 B.n110 VSUBS 0.007277f
C1104 B.n111 VSUBS 0.007277f
C1105 B.n112 VSUBS 0.007277f
C1106 B.n113 VSUBS 0.007277f
C1107 B.n114 VSUBS 0.007277f
C1108 B.n115 VSUBS 0.007277f
C1109 B.n116 VSUBS 0.007277f
C1110 B.n117 VSUBS 0.007277f
C1111 B.n118 VSUBS 0.007277f
C1112 B.n119 VSUBS 0.007277f
C1113 B.n120 VSUBS 0.007277f
C1114 B.n121 VSUBS 0.007277f
C1115 B.n122 VSUBS 0.007277f
C1116 B.n123 VSUBS 0.007277f
C1117 B.n124 VSUBS 0.007277f
C1118 B.n125 VSUBS 0.007277f
C1119 B.n126 VSUBS 0.007277f
C1120 B.n127 VSUBS 0.007277f
C1121 B.n128 VSUBS 0.007277f
C1122 B.n129 VSUBS 0.007277f
C1123 B.n130 VSUBS 0.007277f
C1124 B.n131 VSUBS 0.007277f
C1125 B.n132 VSUBS 0.007277f
C1126 B.n133 VSUBS 0.007277f
C1127 B.n134 VSUBS 0.007277f
C1128 B.n135 VSUBS 0.007277f
C1129 B.n136 VSUBS 0.007277f
C1130 B.n137 VSUBS 0.007277f
C1131 B.n138 VSUBS 0.007277f
C1132 B.n139 VSUBS 0.007277f
C1133 B.n140 VSUBS 0.007277f
C1134 B.n141 VSUBS 0.007277f
C1135 B.n142 VSUBS 0.007277f
C1136 B.n143 VSUBS 0.007277f
C1137 B.n144 VSUBS 0.007277f
C1138 B.n145 VSUBS 0.007277f
C1139 B.n146 VSUBS 0.007277f
C1140 B.n147 VSUBS 0.007277f
C1141 B.n148 VSUBS 0.007277f
C1142 B.n149 VSUBS 0.007277f
C1143 B.n150 VSUBS 0.007277f
C1144 B.n151 VSUBS 0.007277f
C1145 B.n152 VSUBS 0.007277f
C1146 B.n153 VSUBS 0.007277f
C1147 B.n154 VSUBS 0.018144f
C1148 B.n155 VSUBS 0.007277f
C1149 B.n156 VSUBS 0.007277f
C1150 B.n157 VSUBS 0.007277f
C1151 B.n158 VSUBS 0.007277f
C1152 B.n159 VSUBS 0.007277f
C1153 B.n160 VSUBS 0.007277f
C1154 B.n161 VSUBS 0.007277f
C1155 B.n162 VSUBS 0.007277f
C1156 B.n163 VSUBS 0.007277f
C1157 B.n164 VSUBS 0.007277f
C1158 B.n165 VSUBS 0.007277f
C1159 B.n166 VSUBS 0.007277f
C1160 B.n167 VSUBS 0.007277f
C1161 B.n168 VSUBS 0.007277f
C1162 B.n169 VSUBS 0.007277f
C1163 B.n170 VSUBS 0.007277f
C1164 B.n171 VSUBS 0.007277f
C1165 B.n172 VSUBS 0.007277f
C1166 B.n173 VSUBS 0.007277f
C1167 B.n174 VSUBS 0.007277f
C1168 B.n175 VSUBS 0.007277f
C1169 B.n176 VSUBS 0.007277f
C1170 B.n177 VSUBS 0.007277f
C1171 B.n178 VSUBS 0.007277f
C1172 B.n179 VSUBS 0.007277f
C1173 B.n180 VSUBS 0.007277f
C1174 B.n181 VSUBS 0.007277f
C1175 B.n182 VSUBS 0.007277f
C1176 B.t5 VSUBS 0.334918f
C1177 B.t4 VSUBS 0.374348f
C1178 B.t3 VSUBS 2.39297f
C1179 B.n183 VSUBS 0.586557f
C1180 B.n184 VSUBS 0.32856f
C1181 B.n185 VSUBS 0.007277f
C1182 B.n186 VSUBS 0.007277f
C1183 B.n187 VSUBS 0.007277f
C1184 B.n188 VSUBS 0.007277f
C1185 B.t11 VSUBS 0.334914f
C1186 B.t10 VSUBS 0.374345f
C1187 B.t9 VSUBS 2.39297f
C1188 B.n189 VSUBS 0.586561f
C1189 B.n190 VSUBS 0.328563f
C1190 B.n191 VSUBS 0.007277f
C1191 B.n192 VSUBS 0.007277f
C1192 B.n193 VSUBS 0.007277f
C1193 B.n194 VSUBS 0.007277f
C1194 B.n195 VSUBS 0.007277f
C1195 B.n196 VSUBS 0.007277f
C1196 B.n197 VSUBS 0.007277f
C1197 B.n198 VSUBS 0.007277f
C1198 B.n199 VSUBS 0.007277f
C1199 B.n200 VSUBS 0.007277f
C1200 B.n201 VSUBS 0.007277f
C1201 B.n202 VSUBS 0.007277f
C1202 B.n203 VSUBS 0.007277f
C1203 B.n204 VSUBS 0.007277f
C1204 B.n205 VSUBS 0.007277f
C1205 B.n206 VSUBS 0.007277f
C1206 B.n207 VSUBS 0.007277f
C1207 B.n208 VSUBS 0.007277f
C1208 B.n209 VSUBS 0.007277f
C1209 B.n210 VSUBS 0.007277f
C1210 B.n211 VSUBS 0.007277f
C1211 B.n212 VSUBS 0.007277f
C1212 B.n213 VSUBS 0.007277f
C1213 B.n214 VSUBS 0.007277f
C1214 B.n215 VSUBS 0.007277f
C1215 B.n216 VSUBS 0.007277f
C1216 B.n217 VSUBS 0.007277f
C1217 B.n218 VSUBS 0.018144f
C1218 B.n219 VSUBS 0.007277f
C1219 B.n220 VSUBS 0.007277f
C1220 B.n221 VSUBS 0.007277f
C1221 B.n222 VSUBS 0.007277f
C1222 B.n223 VSUBS 0.007277f
C1223 B.n224 VSUBS 0.007277f
C1224 B.n225 VSUBS 0.007277f
C1225 B.n226 VSUBS 0.007277f
C1226 B.n227 VSUBS 0.007277f
C1227 B.n228 VSUBS 0.007277f
C1228 B.n229 VSUBS 0.007277f
C1229 B.n230 VSUBS 0.007277f
C1230 B.n231 VSUBS 0.007277f
C1231 B.n232 VSUBS 0.007277f
C1232 B.n233 VSUBS 0.007277f
C1233 B.n234 VSUBS 0.007277f
C1234 B.n235 VSUBS 0.007277f
C1235 B.n236 VSUBS 0.007277f
C1236 B.n237 VSUBS 0.007277f
C1237 B.n238 VSUBS 0.007277f
C1238 B.n239 VSUBS 0.007277f
C1239 B.n240 VSUBS 0.007277f
C1240 B.n241 VSUBS 0.007277f
C1241 B.n242 VSUBS 0.007277f
C1242 B.n243 VSUBS 0.007277f
C1243 B.n244 VSUBS 0.007277f
C1244 B.n245 VSUBS 0.007277f
C1245 B.n246 VSUBS 0.007277f
C1246 B.n247 VSUBS 0.007277f
C1247 B.n248 VSUBS 0.007277f
C1248 B.n249 VSUBS 0.007277f
C1249 B.n250 VSUBS 0.007277f
C1250 B.n251 VSUBS 0.007277f
C1251 B.n252 VSUBS 0.007277f
C1252 B.n253 VSUBS 0.007277f
C1253 B.n254 VSUBS 0.007277f
C1254 B.n255 VSUBS 0.007277f
C1255 B.n256 VSUBS 0.007277f
C1256 B.n257 VSUBS 0.007277f
C1257 B.n258 VSUBS 0.007277f
C1258 B.n259 VSUBS 0.007277f
C1259 B.n260 VSUBS 0.007277f
C1260 B.n261 VSUBS 0.007277f
C1261 B.n262 VSUBS 0.007277f
C1262 B.n263 VSUBS 0.007277f
C1263 B.n264 VSUBS 0.007277f
C1264 B.n265 VSUBS 0.007277f
C1265 B.n266 VSUBS 0.007277f
C1266 B.n267 VSUBS 0.007277f
C1267 B.n268 VSUBS 0.007277f
C1268 B.n269 VSUBS 0.007277f
C1269 B.n270 VSUBS 0.007277f
C1270 B.n271 VSUBS 0.007277f
C1271 B.n272 VSUBS 0.007277f
C1272 B.n273 VSUBS 0.007277f
C1273 B.n274 VSUBS 0.007277f
C1274 B.n275 VSUBS 0.007277f
C1275 B.n276 VSUBS 0.007277f
C1276 B.n277 VSUBS 0.007277f
C1277 B.n278 VSUBS 0.007277f
C1278 B.n279 VSUBS 0.007277f
C1279 B.n280 VSUBS 0.007277f
C1280 B.n281 VSUBS 0.007277f
C1281 B.n282 VSUBS 0.007277f
C1282 B.n283 VSUBS 0.007277f
C1283 B.n284 VSUBS 0.007277f
C1284 B.n285 VSUBS 0.007277f
C1285 B.n286 VSUBS 0.007277f
C1286 B.n287 VSUBS 0.007277f
C1287 B.n288 VSUBS 0.007277f
C1288 B.n289 VSUBS 0.007277f
C1289 B.n290 VSUBS 0.007277f
C1290 B.n291 VSUBS 0.007277f
C1291 B.n292 VSUBS 0.007277f
C1292 B.n293 VSUBS 0.007277f
C1293 B.n294 VSUBS 0.007277f
C1294 B.n295 VSUBS 0.007277f
C1295 B.n296 VSUBS 0.007277f
C1296 B.n297 VSUBS 0.007277f
C1297 B.n298 VSUBS 0.007277f
C1298 B.n299 VSUBS 0.007277f
C1299 B.n300 VSUBS 0.007277f
C1300 B.n301 VSUBS 0.007277f
C1301 B.n302 VSUBS 0.007277f
C1302 B.n303 VSUBS 0.007277f
C1303 B.n304 VSUBS 0.007277f
C1304 B.n305 VSUBS 0.007277f
C1305 B.n306 VSUBS 0.007277f
C1306 B.n307 VSUBS 0.007277f
C1307 B.n308 VSUBS 0.007277f
C1308 B.n309 VSUBS 0.007277f
C1309 B.n310 VSUBS 0.007277f
C1310 B.n311 VSUBS 0.007277f
C1311 B.n312 VSUBS 0.007277f
C1312 B.n313 VSUBS 0.007277f
C1313 B.n314 VSUBS 0.007277f
C1314 B.n315 VSUBS 0.007277f
C1315 B.n316 VSUBS 0.007277f
C1316 B.n317 VSUBS 0.007277f
C1317 B.n318 VSUBS 0.007277f
C1318 B.n319 VSUBS 0.007277f
C1319 B.n320 VSUBS 0.007277f
C1320 B.n321 VSUBS 0.007277f
C1321 B.n322 VSUBS 0.007277f
C1322 B.n323 VSUBS 0.007277f
C1323 B.n324 VSUBS 0.007277f
C1324 B.n325 VSUBS 0.007277f
C1325 B.n326 VSUBS 0.007277f
C1326 B.n327 VSUBS 0.007277f
C1327 B.n328 VSUBS 0.007277f
C1328 B.n329 VSUBS 0.017171f
C1329 B.n330 VSUBS 0.017171f
C1330 B.n331 VSUBS 0.018144f
C1331 B.n332 VSUBS 0.007277f
C1332 B.n333 VSUBS 0.007277f
C1333 B.n334 VSUBS 0.007277f
C1334 B.n335 VSUBS 0.007277f
C1335 B.n336 VSUBS 0.007277f
C1336 B.n337 VSUBS 0.007277f
C1337 B.n338 VSUBS 0.007277f
C1338 B.n339 VSUBS 0.007277f
C1339 B.n340 VSUBS 0.007277f
C1340 B.n341 VSUBS 0.007277f
C1341 B.n342 VSUBS 0.007277f
C1342 B.n343 VSUBS 0.007277f
C1343 B.n344 VSUBS 0.007277f
C1344 B.n345 VSUBS 0.007277f
C1345 B.n346 VSUBS 0.007277f
C1346 B.n347 VSUBS 0.007277f
C1347 B.n348 VSUBS 0.007277f
C1348 B.n349 VSUBS 0.007277f
C1349 B.n350 VSUBS 0.007277f
C1350 B.n351 VSUBS 0.007277f
C1351 B.n352 VSUBS 0.007277f
C1352 B.n353 VSUBS 0.007277f
C1353 B.n354 VSUBS 0.007277f
C1354 B.n355 VSUBS 0.007277f
C1355 B.n356 VSUBS 0.007277f
C1356 B.n357 VSUBS 0.007277f
C1357 B.n358 VSUBS 0.007277f
C1358 B.n359 VSUBS 0.007277f
C1359 B.n360 VSUBS 0.007277f
C1360 B.n361 VSUBS 0.007277f
C1361 B.n362 VSUBS 0.007277f
C1362 B.n363 VSUBS 0.007277f
C1363 B.n364 VSUBS 0.007277f
C1364 B.n365 VSUBS 0.007277f
C1365 B.n366 VSUBS 0.007277f
C1366 B.n367 VSUBS 0.007277f
C1367 B.n368 VSUBS 0.007277f
C1368 B.n369 VSUBS 0.007277f
C1369 B.n370 VSUBS 0.007277f
C1370 B.n371 VSUBS 0.007277f
C1371 B.n372 VSUBS 0.007277f
C1372 B.n373 VSUBS 0.007277f
C1373 B.n374 VSUBS 0.007277f
C1374 B.n375 VSUBS 0.007277f
C1375 B.n376 VSUBS 0.007277f
C1376 B.n377 VSUBS 0.007277f
C1377 B.n378 VSUBS 0.007277f
C1378 B.n379 VSUBS 0.007277f
C1379 B.n380 VSUBS 0.007277f
C1380 B.n381 VSUBS 0.007277f
C1381 B.n382 VSUBS 0.007277f
C1382 B.n383 VSUBS 0.007277f
C1383 B.n384 VSUBS 0.007277f
C1384 B.n385 VSUBS 0.007277f
C1385 B.n386 VSUBS 0.007277f
C1386 B.n387 VSUBS 0.007277f
C1387 B.n388 VSUBS 0.007277f
C1388 B.n389 VSUBS 0.007277f
C1389 B.n390 VSUBS 0.007277f
C1390 B.n391 VSUBS 0.007277f
C1391 B.n392 VSUBS 0.007277f
C1392 B.n393 VSUBS 0.007277f
C1393 B.n394 VSUBS 0.007277f
C1394 B.n395 VSUBS 0.007277f
C1395 B.n396 VSUBS 0.007277f
C1396 B.n397 VSUBS 0.007277f
C1397 B.n398 VSUBS 0.007277f
C1398 B.n399 VSUBS 0.007277f
C1399 B.n400 VSUBS 0.007277f
C1400 B.n401 VSUBS 0.007277f
C1401 B.n402 VSUBS 0.007277f
C1402 B.n403 VSUBS 0.007277f
C1403 B.n404 VSUBS 0.007277f
C1404 B.n405 VSUBS 0.007277f
C1405 B.n406 VSUBS 0.007277f
C1406 B.n407 VSUBS 0.007277f
C1407 B.n408 VSUBS 0.007277f
C1408 B.n409 VSUBS 0.007277f
C1409 B.n410 VSUBS 0.007277f
C1410 B.n411 VSUBS 0.007277f
C1411 B.n412 VSUBS 0.007277f
C1412 B.n413 VSUBS 0.007277f
C1413 B.n414 VSUBS 0.00503f
C1414 B.n415 VSUBS 0.01686f
C1415 B.n416 VSUBS 0.005886f
C1416 B.n417 VSUBS 0.007277f
C1417 B.n418 VSUBS 0.007277f
C1418 B.n419 VSUBS 0.007277f
C1419 B.n420 VSUBS 0.007277f
C1420 B.n421 VSUBS 0.007277f
C1421 B.n422 VSUBS 0.007277f
C1422 B.n423 VSUBS 0.007277f
C1423 B.n424 VSUBS 0.007277f
C1424 B.n425 VSUBS 0.007277f
C1425 B.n426 VSUBS 0.007277f
C1426 B.n427 VSUBS 0.007277f
C1427 B.n428 VSUBS 0.005886f
C1428 B.n429 VSUBS 0.01686f
C1429 B.n430 VSUBS 0.00503f
C1430 B.n431 VSUBS 0.007277f
C1431 B.n432 VSUBS 0.007277f
C1432 B.n433 VSUBS 0.007277f
C1433 B.n434 VSUBS 0.007277f
C1434 B.n435 VSUBS 0.007277f
C1435 B.n436 VSUBS 0.007277f
C1436 B.n437 VSUBS 0.007277f
C1437 B.n438 VSUBS 0.007277f
C1438 B.n439 VSUBS 0.007277f
C1439 B.n440 VSUBS 0.007277f
C1440 B.n441 VSUBS 0.007277f
C1441 B.n442 VSUBS 0.007277f
C1442 B.n443 VSUBS 0.007277f
C1443 B.n444 VSUBS 0.007277f
C1444 B.n445 VSUBS 0.007277f
C1445 B.n446 VSUBS 0.007277f
C1446 B.n447 VSUBS 0.007277f
C1447 B.n448 VSUBS 0.007277f
C1448 B.n449 VSUBS 0.007277f
C1449 B.n450 VSUBS 0.007277f
C1450 B.n451 VSUBS 0.007277f
C1451 B.n452 VSUBS 0.007277f
C1452 B.n453 VSUBS 0.007277f
C1453 B.n454 VSUBS 0.007277f
C1454 B.n455 VSUBS 0.007277f
C1455 B.n456 VSUBS 0.007277f
C1456 B.n457 VSUBS 0.007277f
C1457 B.n458 VSUBS 0.007277f
C1458 B.n459 VSUBS 0.007277f
C1459 B.n460 VSUBS 0.007277f
C1460 B.n461 VSUBS 0.007277f
C1461 B.n462 VSUBS 0.007277f
C1462 B.n463 VSUBS 0.007277f
C1463 B.n464 VSUBS 0.007277f
C1464 B.n465 VSUBS 0.007277f
C1465 B.n466 VSUBS 0.007277f
C1466 B.n467 VSUBS 0.007277f
C1467 B.n468 VSUBS 0.007277f
C1468 B.n469 VSUBS 0.007277f
C1469 B.n470 VSUBS 0.007277f
C1470 B.n471 VSUBS 0.007277f
C1471 B.n472 VSUBS 0.007277f
C1472 B.n473 VSUBS 0.007277f
C1473 B.n474 VSUBS 0.007277f
C1474 B.n475 VSUBS 0.007277f
C1475 B.n476 VSUBS 0.007277f
C1476 B.n477 VSUBS 0.007277f
C1477 B.n478 VSUBS 0.007277f
C1478 B.n479 VSUBS 0.007277f
C1479 B.n480 VSUBS 0.007277f
C1480 B.n481 VSUBS 0.007277f
C1481 B.n482 VSUBS 0.007277f
C1482 B.n483 VSUBS 0.007277f
C1483 B.n484 VSUBS 0.007277f
C1484 B.n485 VSUBS 0.007277f
C1485 B.n486 VSUBS 0.007277f
C1486 B.n487 VSUBS 0.007277f
C1487 B.n488 VSUBS 0.007277f
C1488 B.n489 VSUBS 0.007277f
C1489 B.n490 VSUBS 0.007277f
C1490 B.n491 VSUBS 0.007277f
C1491 B.n492 VSUBS 0.007277f
C1492 B.n493 VSUBS 0.007277f
C1493 B.n494 VSUBS 0.007277f
C1494 B.n495 VSUBS 0.007277f
C1495 B.n496 VSUBS 0.007277f
C1496 B.n497 VSUBS 0.007277f
C1497 B.n498 VSUBS 0.007277f
C1498 B.n499 VSUBS 0.007277f
C1499 B.n500 VSUBS 0.007277f
C1500 B.n501 VSUBS 0.007277f
C1501 B.n502 VSUBS 0.007277f
C1502 B.n503 VSUBS 0.007277f
C1503 B.n504 VSUBS 0.007277f
C1504 B.n505 VSUBS 0.007277f
C1505 B.n506 VSUBS 0.007277f
C1506 B.n507 VSUBS 0.007277f
C1507 B.n508 VSUBS 0.007277f
C1508 B.n509 VSUBS 0.007277f
C1509 B.n510 VSUBS 0.007277f
C1510 B.n511 VSUBS 0.007277f
C1511 B.n512 VSUBS 0.007277f
C1512 B.n513 VSUBS 0.01733f
C1513 B.n514 VSUBS 0.017985f
C1514 B.n515 VSUBS 0.017171f
C1515 B.n516 VSUBS 0.007277f
C1516 B.n517 VSUBS 0.007277f
C1517 B.n518 VSUBS 0.007277f
C1518 B.n519 VSUBS 0.007277f
C1519 B.n520 VSUBS 0.007277f
C1520 B.n521 VSUBS 0.007277f
C1521 B.n522 VSUBS 0.007277f
C1522 B.n523 VSUBS 0.007277f
C1523 B.n524 VSUBS 0.007277f
C1524 B.n525 VSUBS 0.007277f
C1525 B.n526 VSUBS 0.007277f
C1526 B.n527 VSUBS 0.007277f
C1527 B.n528 VSUBS 0.007277f
C1528 B.n529 VSUBS 0.007277f
C1529 B.n530 VSUBS 0.007277f
C1530 B.n531 VSUBS 0.007277f
C1531 B.n532 VSUBS 0.007277f
C1532 B.n533 VSUBS 0.007277f
C1533 B.n534 VSUBS 0.007277f
C1534 B.n535 VSUBS 0.007277f
C1535 B.n536 VSUBS 0.007277f
C1536 B.n537 VSUBS 0.007277f
C1537 B.n538 VSUBS 0.007277f
C1538 B.n539 VSUBS 0.007277f
C1539 B.n540 VSUBS 0.007277f
C1540 B.n541 VSUBS 0.007277f
C1541 B.n542 VSUBS 0.007277f
C1542 B.n543 VSUBS 0.007277f
C1543 B.n544 VSUBS 0.007277f
C1544 B.n545 VSUBS 0.007277f
C1545 B.n546 VSUBS 0.007277f
C1546 B.n547 VSUBS 0.007277f
C1547 B.n548 VSUBS 0.007277f
C1548 B.n549 VSUBS 0.007277f
C1549 B.n550 VSUBS 0.007277f
C1550 B.n551 VSUBS 0.007277f
C1551 B.n552 VSUBS 0.007277f
C1552 B.n553 VSUBS 0.007277f
C1553 B.n554 VSUBS 0.007277f
C1554 B.n555 VSUBS 0.007277f
C1555 B.n556 VSUBS 0.007277f
C1556 B.n557 VSUBS 0.007277f
C1557 B.n558 VSUBS 0.007277f
C1558 B.n559 VSUBS 0.007277f
C1559 B.n560 VSUBS 0.007277f
C1560 B.n561 VSUBS 0.007277f
C1561 B.n562 VSUBS 0.007277f
C1562 B.n563 VSUBS 0.007277f
C1563 B.n564 VSUBS 0.007277f
C1564 B.n565 VSUBS 0.007277f
C1565 B.n566 VSUBS 0.007277f
C1566 B.n567 VSUBS 0.007277f
C1567 B.n568 VSUBS 0.007277f
C1568 B.n569 VSUBS 0.007277f
C1569 B.n570 VSUBS 0.007277f
C1570 B.n571 VSUBS 0.007277f
C1571 B.n572 VSUBS 0.007277f
C1572 B.n573 VSUBS 0.007277f
C1573 B.n574 VSUBS 0.007277f
C1574 B.n575 VSUBS 0.007277f
C1575 B.n576 VSUBS 0.007277f
C1576 B.n577 VSUBS 0.007277f
C1577 B.n578 VSUBS 0.007277f
C1578 B.n579 VSUBS 0.007277f
C1579 B.n580 VSUBS 0.007277f
C1580 B.n581 VSUBS 0.007277f
C1581 B.n582 VSUBS 0.007277f
C1582 B.n583 VSUBS 0.007277f
C1583 B.n584 VSUBS 0.007277f
C1584 B.n585 VSUBS 0.007277f
C1585 B.n586 VSUBS 0.007277f
C1586 B.n587 VSUBS 0.007277f
C1587 B.n588 VSUBS 0.007277f
C1588 B.n589 VSUBS 0.007277f
C1589 B.n590 VSUBS 0.007277f
C1590 B.n591 VSUBS 0.007277f
C1591 B.n592 VSUBS 0.007277f
C1592 B.n593 VSUBS 0.007277f
C1593 B.n594 VSUBS 0.007277f
C1594 B.n595 VSUBS 0.007277f
C1595 B.n596 VSUBS 0.007277f
C1596 B.n597 VSUBS 0.007277f
C1597 B.n598 VSUBS 0.007277f
C1598 B.n599 VSUBS 0.007277f
C1599 B.n600 VSUBS 0.007277f
C1600 B.n601 VSUBS 0.007277f
C1601 B.n602 VSUBS 0.007277f
C1602 B.n603 VSUBS 0.007277f
C1603 B.n604 VSUBS 0.007277f
C1604 B.n605 VSUBS 0.007277f
C1605 B.n606 VSUBS 0.007277f
C1606 B.n607 VSUBS 0.007277f
C1607 B.n608 VSUBS 0.007277f
C1608 B.n609 VSUBS 0.007277f
C1609 B.n610 VSUBS 0.007277f
C1610 B.n611 VSUBS 0.007277f
C1611 B.n612 VSUBS 0.007277f
C1612 B.n613 VSUBS 0.007277f
C1613 B.n614 VSUBS 0.007277f
C1614 B.n615 VSUBS 0.007277f
C1615 B.n616 VSUBS 0.007277f
C1616 B.n617 VSUBS 0.007277f
C1617 B.n618 VSUBS 0.007277f
C1618 B.n619 VSUBS 0.007277f
C1619 B.n620 VSUBS 0.007277f
C1620 B.n621 VSUBS 0.007277f
C1621 B.n622 VSUBS 0.007277f
C1622 B.n623 VSUBS 0.007277f
C1623 B.n624 VSUBS 0.007277f
C1624 B.n625 VSUBS 0.007277f
C1625 B.n626 VSUBS 0.007277f
C1626 B.n627 VSUBS 0.007277f
C1627 B.n628 VSUBS 0.007277f
C1628 B.n629 VSUBS 0.007277f
C1629 B.n630 VSUBS 0.007277f
C1630 B.n631 VSUBS 0.007277f
C1631 B.n632 VSUBS 0.007277f
C1632 B.n633 VSUBS 0.007277f
C1633 B.n634 VSUBS 0.007277f
C1634 B.n635 VSUBS 0.007277f
C1635 B.n636 VSUBS 0.007277f
C1636 B.n637 VSUBS 0.007277f
C1637 B.n638 VSUBS 0.007277f
C1638 B.n639 VSUBS 0.007277f
C1639 B.n640 VSUBS 0.007277f
C1640 B.n641 VSUBS 0.007277f
C1641 B.n642 VSUBS 0.007277f
C1642 B.n643 VSUBS 0.007277f
C1643 B.n644 VSUBS 0.007277f
C1644 B.n645 VSUBS 0.007277f
C1645 B.n646 VSUBS 0.007277f
C1646 B.n647 VSUBS 0.007277f
C1647 B.n648 VSUBS 0.007277f
C1648 B.n649 VSUBS 0.007277f
C1649 B.n650 VSUBS 0.007277f
C1650 B.n651 VSUBS 0.007277f
C1651 B.n652 VSUBS 0.007277f
C1652 B.n653 VSUBS 0.007277f
C1653 B.n654 VSUBS 0.007277f
C1654 B.n655 VSUBS 0.007277f
C1655 B.n656 VSUBS 0.007277f
C1656 B.n657 VSUBS 0.007277f
C1657 B.n658 VSUBS 0.007277f
C1658 B.n659 VSUBS 0.007277f
C1659 B.n660 VSUBS 0.007277f
C1660 B.n661 VSUBS 0.007277f
C1661 B.n662 VSUBS 0.007277f
C1662 B.n663 VSUBS 0.007277f
C1663 B.n664 VSUBS 0.007277f
C1664 B.n665 VSUBS 0.007277f
C1665 B.n666 VSUBS 0.007277f
C1666 B.n667 VSUBS 0.007277f
C1667 B.n668 VSUBS 0.007277f
C1668 B.n669 VSUBS 0.007277f
C1669 B.n670 VSUBS 0.007277f
C1670 B.n671 VSUBS 0.007277f
C1671 B.n672 VSUBS 0.007277f
C1672 B.n673 VSUBS 0.007277f
C1673 B.n674 VSUBS 0.007277f
C1674 B.n675 VSUBS 0.007277f
C1675 B.n676 VSUBS 0.007277f
C1676 B.n677 VSUBS 0.007277f
C1677 B.n678 VSUBS 0.007277f
C1678 B.n679 VSUBS 0.007277f
C1679 B.n680 VSUBS 0.007277f
C1680 B.n681 VSUBS 0.007277f
C1681 B.n682 VSUBS 0.007277f
C1682 B.n683 VSUBS 0.007277f
C1683 B.n684 VSUBS 0.007277f
C1684 B.n685 VSUBS 0.007277f
C1685 B.n686 VSUBS 0.007277f
C1686 B.n687 VSUBS 0.017171f
C1687 B.n688 VSUBS 0.018144f
C1688 B.n689 VSUBS 0.018144f
C1689 B.n690 VSUBS 0.007277f
C1690 B.n691 VSUBS 0.007277f
C1691 B.n692 VSUBS 0.007277f
C1692 B.n693 VSUBS 0.007277f
C1693 B.n694 VSUBS 0.007277f
C1694 B.n695 VSUBS 0.007277f
C1695 B.n696 VSUBS 0.007277f
C1696 B.n697 VSUBS 0.007277f
C1697 B.n698 VSUBS 0.007277f
C1698 B.n699 VSUBS 0.007277f
C1699 B.n700 VSUBS 0.007277f
C1700 B.n701 VSUBS 0.007277f
C1701 B.n702 VSUBS 0.007277f
C1702 B.n703 VSUBS 0.007277f
C1703 B.n704 VSUBS 0.007277f
C1704 B.n705 VSUBS 0.007277f
C1705 B.n706 VSUBS 0.007277f
C1706 B.n707 VSUBS 0.007277f
C1707 B.n708 VSUBS 0.007277f
C1708 B.n709 VSUBS 0.007277f
C1709 B.n710 VSUBS 0.007277f
C1710 B.n711 VSUBS 0.007277f
C1711 B.n712 VSUBS 0.007277f
C1712 B.n713 VSUBS 0.007277f
C1713 B.n714 VSUBS 0.007277f
C1714 B.n715 VSUBS 0.007277f
C1715 B.n716 VSUBS 0.007277f
C1716 B.n717 VSUBS 0.007277f
C1717 B.n718 VSUBS 0.007277f
C1718 B.n719 VSUBS 0.007277f
C1719 B.n720 VSUBS 0.007277f
C1720 B.n721 VSUBS 0.007277f
C1721 B.n722 VSUBS 0.007277f
C1722 B.n723 VSUBS 0.007277f
C1723 B.n724 VSUBS 0.007277f
C1724 B.n725 VSUBS 0.007277f
C1725 B.n726 VSUBS 0.007277f
C1726 B.n727 VSUBS 0.007277f
C1727 B.n728 VSUBS 0.007277f
C1728 B.n729 VSUBS 0.007277f
C1729 B.n730 VSUBS 0.007277f
C1730 B.n731 VSUBS 0.007277f
C1731 B.n732 VSUBS 0.007277f
C1732 B.n733 VSUBS 0.007277f
C1733 B.n734 VSUBS 0.007277f
C1734 B.n735 VSUBS 0.007277f
C1735 B.n736 VSUBS 0.007277f
C1736 B.n737 VSUBS 0.007277f
C1737 B.n738 VSUBS 0.007277f
C1738 B.n739 VSUBS 0.007277f
C1739 B.n740 VSUBS 0.007277f
C1740 B.n741 VSUBS 0.007277f
C1741 B.n742 VSUBS 0.007277f
C1742 B.n743 VSUBS 0.007277f
C1743 B.n744 VSUBS 0.007277f
C1744 B.n745 VSUBS 0.007277f
C1745 B.n746 VSUBS 0.007277f
C1746 B.n747 VSUBS 0.007277f
C1747 B.n748 VSUBS 0.007277f
C1748 B.n749 VSUBS 0.007277f
C1749 B.n750 VSUBS 0.007277f
C1750 B.n751 VSUBS 0.007277f
C1751 B.n752 VSUBS 0.007277f
C1752 B.n753 VSUBS 0.007277f
C1753 B.n754 VSUBS 0.007277f
C1754 B.n755 VSUBS 0.007277f
C1755 B.n756 VSUBS 0.007277f
C1756 B.n757 VSUBS 0.007277f
C1757 B.n758 VSUBS 0.007277f
C1758 B.n759 VSUBS 0.007277f
C1759 B.n760 VSUBS 0.007277f
C1760 B.n761 VSUBS 0.007277f
C1761 B.n762 VSUBS 0.007277f
C1762 B.n763 VSUBS 0.007277f
C1763 B.n764 VSUBS 0.007277f
C1764 B.n765 VSUBS 0.007277f
C1765 B.n766 VSUBS 0.007277f
C1766 B.n767 VSUBS 0.007277f
C1767 B.n768 VSUBS 0.007277f
C1768 B.n769 VSUBS 0.007277f
C1769 B.n770 VSUBS 0.007277f
C1770 B.n771 VSUBS 0.00503f
C1771 B.n772 VSUBS 0.01686f
C1772 B.n773 VSUBS 0.005886f
C1773 B.n774 VSUBS 0.007277f
C1774 B.n775 VSUBS 0.007277f
C1775 B.n776 VSUBS 0.007277f
C1776 B.n777 VSUBS 0.007277f
C1777 B.n778 VSUBS 0.007277f
C1778 B.n779 VSUBS 0.007277f
C1779 B.n780 VSUBS 0.007277f
C1780 B.n781 VSUBS 0.007277f
C1781 B.n782 VSUBS 0.007277f
C1782 B.n783 VSUBS 0.007277f
C1783 B.n784 VSUBS 0.007277f
C1784 B.n785 VSUBS 0.005886f
C1785 B.n786 VSUBS 0.007277f
C1786 B.n787 VSUBS 0.007277f
C1787 B.n788 VSUBS 0.007277f
C1788 B.n789 VSUBS 0.007277f
C1789 B.n790 VSUBS 0.007277f
C1790 B.n791 VSUBS 0.007277f
C1791 B.n792 VSUBS 0.007277f
C1792 B.n793 VSUBS 0.007277f
C1793 B.n794 VSUBS 0.007277f
C1794 B.n795 VSUBS 0.007277f
C1795 B.n796 VSUBS 0.007277f
C1796 B.n797 VSUBS 0.007277f
C1797 B.n798 VSUBS 0.007277f
C1798 B.n799 VSUBS 0.007277f
C1799 B.n800 VSUBS 0.007277f
C1800 B.n801 VSUBS 0.007277f
C1801 B.n802 VSUBS 0.007277f
C1802 B.n803 VSUBS 0.007277f
C1803 B.n804 VSUBS 0.007277f
C1804 B.n805 VSUBS 0.007277f
C1805 B.n806 VSUBS 0.007277f
C1806 B.n807 VSUBS 0.007277f
C1807 B.n808 VSUBS 0.007277f
C1808 B.n809 VSUBS 0.007277f
C1809 B.n810 VSUBS 0.007277f
C1810 B.n811 VSUBS 0.007277f
C1811 B.n812 VSUBS 0.007277f
C1812 B.n813 VSUBS 0.007277f
C1813 B.n814 VSUBS 0.007277f
C1814 B.n815 VSUBS 0.007277f
C1815 B.n816 VSUBS 0.007277f
C1816 B.n817 VSUBS 0.007277f
C1817 B.n818 VSUBS 0.007277f
C1818 B.n819 VSUBS 0.007277f
C1819 B.n820 VSUBS 0.007277f
C1820 B.n821 VSUBS 0.007277f
C1821 B.n822 VSUBS 0.007277f
C1822 B.n823 VSUBS 0.007277f
C1823 B.n824 VSUBS 0.007277f
C1824 B.n825 VSUBS 0.007277f
C1825 B.n826 VSUBS 0.007277f
C1826 B.n827 VSUBS 0.007277f
C1827 B.n828 VSUBS 0.007277f
C1828 B.n829 VSUBS 0.007277f
C1829 B.n830 VSUBS 0.007277f
C1830 B.n831 VSUBS 0.007277f
C1831 B.n832 VSUBS 0.007277f
C1832 B.n833 VSUBS 0.007277f
C1833 B.n834 VSUBS 0.007277f
C1834 B.n835 VSUBS 0.007277f
C1835 B.n836 VSUBS 0.007277f
C1836 B.n837 VSUBS 0.007277f
C1837 B.n838 VSUBS 0.007277f
C1838 B.n839 VSUBS 0.007277f
C1839 B.n840 VSUBS 0.007277f
C1840 B.n841 VSUBS 0.007277f
C1841 B.n842 VSUBS 0.007277f
C1842 B.n843 VSUBS 0.007277f
C1843 B.n844 VSUBS 0.007277f
C1844 B.n845 VSUBS 0.007277f
C1845 B.n846 VSUBS 0.007277f
C1846 B.n847 VSUBS 0.007277f
C1847 B.n848 VSUBS 0.007277f
C1848 B.n849 VSUBS 0.007277f
C1849 B.n850 VSUBS 0.007277f
C1850 B.n851 VSUBS 0.007277f
C1851 B.n852 VSUBS 0.007277f
C1852 B.n853 VSUBS 0.007277f
C1853 B.n854 VSUBS 0.007277f
C1854 B.n855 VSUBS 0.007277f
C1855 B.n856 VSUBS 0.007277f
C1856 B.n857 VSUBS 0.007277f
C1857 B.n858 VSUBS 0.007277f
C1858 B.n859 VSUBS 0.007277f
C1859 B.n860 VSUBS 0.007277f
C1860 B.n861 VSUBS 0.007277f
C1861 B.n862 VSUBS 0.007277f
C1862 B.n863 VSUBS 0.007277f
C1863 B.n864 VSUBS 0.007277f
C1864 B.n865 VSUBS 0.007277f
C1865 B.n866 VSUBS 0.007277f
C1866 B.n867 VSUBS 0.007277f
C1867 B.n868 VSUBS 0.007277f
C1868 B.n869 VSUBS 0.018144f
C1869 B.n870 VSUBS 0.018144f
C1870 B.n871 VSUBS 0.017171f
C1871 B.n872 VSUBS 0.007277f
C1872 B.n873 VSUBS 0.007277f
C1873 B.n874 VSUBS 0.007277f
C1874 B.n875 VSUBS 0.007277f
C1875 B.n876 VSUBS 0.007277f
C1876 B.n877 VSUBS 0.007277f
C1877 B.n878 VSUBS 0.007277f
C1878 B.n879 VSUBS 0.007277f
C1879 B.n880 VSUBS 0.007277f
C1880 B.n881 VSUBS 0.007277f
C1881 B.n882 VSUBS 0.007277f
C1882 B.n883 VSUBS 0.007277f
C1883 B.n884 VSUBS 0.007277f
C1884 B.n885 VSUBS 0.007277f
C1885 B.n886 VSUBS 0.007277f
C1886 B.n887 VSUBS 0.007277f
C1887 B.n888 VSUBS 0.007277f
C1888 B.n889 VSUBS 0.007277f
C1889 B.n890 VSUBS 0.007277f
C1890 B.n891 VSUBS 0.007277f
C1891 B.n892 VSUBS 0.007277f
C1892 B.n893 VSUBS 0.007277f
C1893 B.n894 VSUBS 0.007277f
C1894 B.n895 VSUBS 0.007277f
C1895 B.n896 VSUBS 0.007277f
C1896 B.n897 VSUBS 0.007277f
C1897 B.n898 VSUBS 0.007277f
C1898 B.n899 VSUBS 0.007277f
C1899 B.n900 VSUBS 0.007277f
C1900 B.n901 VSUBS 0.007277f
C1901 B.n902 VSUBS 0.007277f
C1902 B.n903 VSUBS 0.007277f
C1903 B.n904 VSUBS 0.007277f
C1904 B.n905 VSUBS 0.007277f
C1905 B.n906 VSUBS 0.007277f
C1906 B.n907 VSUBS 0.007277f
C1907 B.n908 VSUBS 0.007277f
C1908 B.n909 VSUBS 0.007277f
C1909 B.n910 VSUBS 0.007277f
C1910 B.n911 VSUBS 0.007277f
C1911 B.n912 VSUBS 0.007277f
C1912 B.n913 VSUBS 0.007277f
C1913 B.n914 VSUBS 0.007277f
C1914 B.n915 VSUBS 0.007277f
C1915 B.n916 VSUBS 0.007277f
C1916 B.n917 VSUBS 0.007277f
C1917 B.n918 VSUBS 0.007277f
C1918 B.n919 VSUBS 0.007277f
C1919 B.n920 VSUBS 0.007277f
C1920 B.n921 VSUBS 0.007277f
C1921 B.n922 VSUBS 0.007277f
C1922 B.n923 VSUBS 0.007277f
C1923 B.n924 VSUBS 0.007277f
C1924 B.n925 VSUBS 0.007277f
C1925 B.n926 VSUBS 0.007277f
C1926 B.n927 VSUBS 0.007277f
C1927 B.n928 VSUBS 0.007277f
C1928 B.n929 VSUBS 0.007277f
C1929 B.n930 VSUBS 0.007277f
C1930 B.n931 VSUBS 0.007277f
C1931 B.n932 VSUBS 0.007277f
C1932 B.n933 VSUBS 0.007277f
C1933 B.n934 VSUBS 0.007277f
C1934 B.n935 VSUBS 0.007277f
C1935 B.n936 VSUBS 0.007277f
C1936 B.n937 VSUBS 0.007277f
C1937 B.n938 VSUBS 0.007277f
C1938 B.n939 VSUBS 0.007277f
C1939 B.n940 VSUBS 0.007277f
C1940 B.n941 VSUBS 0.007277f
C1941 B.n942 VSUBS 0.007277f
C1942 B.n943 VSUBS 0.007277f
C1943 B.n944 VSUBS 0.007277f
C1944 B.n945 VSUBS 0.007277f
C1945 B.n946 VSUBS 0.007277f
C1946 B.n947 VSUBS 0.007277f
C1947 B.n948 VSUBS 0.007277f
C1948 B.n949 VSUBS 0.007277f
C1949 B.n950 VSUBS 0.007277f
C1950 B.n951 VSUBS 0.007277f
C1951 B.n952 VSUBS 0.007277f
C1952 B.n953 VSUBS 0.007277f
C1953 B.n954 VSUBS 0.007277f
C1954 B.n955 VSUBS 0.009496f
C1955 B.n956 VSUBS 0.010116f
C1956 B.n957 VSUBS 0.020116f
.ends

