* NGSPICE file created from diff_pair_sample_0901.ext - technology: sky130A

.subckt diff_pair_sample_0901 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t9 VP.t0 VTAIL.t12 w_n4570_n2674# sky130_fd_pr__pfet_01v8 ad=1.40745 pd=8.86 as=3.3267 ps=17.84 w=8.53 l=2.67
X1 VTAIL.t11 VP.t1 VDD1.t8 w_n4570_n2674# sky130_fd_pr__pfet_01v8 ad=1.40745 pd=8.86 as=1.40745 ps=8.86 w=8.53 l=2.67
X2 VDD2.t9 VN.t0 VTAIL.t5 w_n4570_n2674# sky130_fd_pr__pfet_01v8 ad=3.3267 pd=17.84 as=1.40745 ps=8.86 w=8.53 l=2.67
X3 VTAIL.t1 VN.t1 VDD2.t8 w_n4570_n2674# sky130_fd_pr__pfet_01v8 ad=1.40745 pd=8.86 as=1.40745 ps=8.86 w=8.53 l=2.67
X4 VDD1.t7 VP.t2 VTAIL.t10 w_n4570_n2674# sky130_fd_pr__pfet_01v8 ad=1.40745 pd=8.86 as=1.40745 ps=8.86 w=8.53 l=2.67
X5 VTAIL.t15 VP.t3 VDD1.t6 w_n4570_n2674# sky130_fd_pr__pfet_01v8 ad=1.40745 pd=8.86 as=1.40745 ps=8.86 w=8.53 l=2.67
X6 VTAIL.t2 VN.t2 VDD2.t7 w_n4570_n2674# sky130_fd_pr__pfet_01v8 ad=1.40745 pd=8.86 as=1.40745 ps=8.86 w=8.53 l=2.67
X7 VTAIL.t4 VN.t3 VDD2.t6 w_n4570_n2674# sky130_fd_pr__pfet_01v8 ad=1.40745 pd=8.86 as=1.40745 ps=8.86 w=8.53 l=2.67
X8 VDD2.t5 VN.t4 VTAIL.t6 w_n4570_n2674# sky130_fd_pr__pfet_01v8 ad=1.40745 pd=8.86 as=3.3267 ps=17.84 w=8.53 l=2.67
X9 VTAIL.t14 VP.t4 VDD1.t5 w_n4570_n2674# sky130_fd_pr__pfet_01v8 ad=1.40745 pd=8.86 as=1.40745 ps=8.86 w=8.53 l=2.67
X10 VDD2.t4 VN.t5 VTAIL.t9 w_n4570_n2674# sky130_fd_pr__pfet_01v8 ad=1.40745 pd=8.86 as=3.3267 ps=17.84 w=8.53 l=2.67
X11 VDD1.t4 VP.t5 VTAIL.t18 w_n4570_n2674# sky130_fd_pr__pfet_01v8 ad=3.3267 pd=17.84 as=1.40745 ps=8.86 w=8.53 l=2.67
X12 B.t11 B.t9 B.t10 w_n4570_n2674# sky130_fd_pr__pfet_01v8 ad=3.3267 pd=17.84 as=0 ps=0 w=8.53 l=2.67
X13 VTAIL.t3 VN.t6 VDD2.t3 w_n4570_n2674# sky130_fd_pr__pfet_01v8 ad=1.40745 pd=8.86 as=1.40745 ps=8.86 w=8.53 l=2.67
X14 VDD1.t3 VP.t6 VTAIL.t17 w_n4570_n2674# sky130_fd_pr__pfet_01v8 ad=1.40745 pd=8.86 as=1.40745 ps=8.86 w=8.53 l=2.67
X15 B.t8 B.t6 B.t7 w_n4570_n2674# sky130_fd_pr__pfet_01v8 ad=3.3267 pd=17.84 as=0 ps=0 w=8.53 l=2.67
X16 VDD2.t2 VN.t7 VTAIL.t0 w_n4570_n2674# sky130_fd_pr__pfet_01v8 ad=1.40745 pd=8.86 as=1.40745 ps=8.86 w=8.53 l=2.67
X17 B.t5 B.t3 B.t4 w_n4570_n2674# sky130_fd_pr__pfet_01v8 ad=3.3267 pd=17.84 as=0 ps=0 w=8.53 l=2.67
X18 VDD1.t2 VP.t7 VTAIL.t16 w_n4570_n2674# sky130_fd_pr__pfet_01v8 ad=3.3267 pd=17.84 as=1.40745 ps=8.86 w=8.53 l=2.67
X19 B.t2 B.t0 B.t1 w_n4570_n2674# sky130_fd_pr__pfet_01v8 ad=3.3267 pd=17.84 as=0 ps=0 w=8.53 l=2.67
X20 VDD2.t1 VN.t8 VTAIL.t8 w_n4570_n2674# sky130_fd_pr__pfet_01v8 ad=3.3267 pd=17.84 as=1.40745 ps=8.86 w=8.53 l=2.67
X21 VTAIL.t13 VP.t8 VDD1.t1 w_n4570_n2674# sky130_fd_pr__pfet_01v8 ad=1.40745 pd=8.86 as=1.40745 ps=8.86 w=8.53 l=2.67
X22 VDD2.t0 VN.t9 VTAIL.t7 w_n4570_n2674# sky130_fd_pr__pfet_01v8 ad=1.40745 pd=8.86 as=1.40745 ps=8.86 w=8.53 l=2.67
X23 VDD1.t0 VP.t9 VTAIL.t19 w_n4570_n2674# sky130_fd_pr__pfet_01v8 ad=1.40745 pd=8.86 as=3.3267 ps=17.84 w=8.53 l=2.67
R0 VP.n25 VP.n24 161.3
R1 VP.n26 VP.n21 161.3
R2 VP.n28 VP.n27 161.3
R3 VP.n29 VP.n20 161.3
R4 VP.n31 VP.n30 161.3
R5 VP.n32 VP.n19 161.3
R6 VP.n34 VP.n33 161.3
R7 VP.n35 VP.n18 161.3
R8 VP.n37 VP.n36 161.3
R9 VP.n38 VP.n17 161.3
R10 VP.n40 VP.n39 161.3
R11 VP.n41 VP.n16 161.3
R12 VP.n43 VP.n42 161.3
R13 VP.n44 VP.n15 161.3
R14 VP.n46 VP.n45 161.3
R15 VP.n47 VP.n14 161.3
R16 VP.n49 VP.n48 161.3
R17 VP.n86 VP.n85 161.3
R18 VP.n84 VP.n1 161.3
R19 VP.n83 VP.n82 161.3
R20 VP.n81 VP.n2 161.3
R21 VP.n80 VP.n79 161.3
R22 VP.n78 VP.n3 161.3
R23 VP.n77 VP.n76 161.3
R24 VP.n75 VP.n4 161.3
R25 VP.n74 VP.n73 161.3
R26 VP.n72 VP.n5 161.3
R27 VP.n71 VP.n70 161.3
R28 VP.n69 VP.n6 161.3
R29 VP.n68 VP.n67 161.3
R30 VP.n66 VP.n7 161.3
R31 VP.n65 VP.n64 161.3
R32 VP.n63 VP.n8 161.3
R33 VP.n62 VP.n61 161.3
R34 VP.n60 VP.n9 161.3
R35 VP.n59 VP.n58 161.3
R36 VP.n57 VP.n10 161.3
R37 VP.n56 VP.n55 161.3
R38 VP.n54 VP.n11 161.3
R39 VP.n53 VP.n52 161.3
R40 VP.n22 VP.t7 109.144
R41 VP.n0 VP.t9 76.9941
R42 VP.n78 VP.t4 76.9941
R43 VP.n6 VP.t6 76.9941
R44 VP.n60 VP.t3 76.9941
R45 VP.n12 VP.t5 76.9941
R46 VP.n23 VP.t8 76.9941
R47 VP.n19 VP.t2 76.9941
R48 VP.n41 VP.t1 76.9941
R49 VP.n13 VP.t0 76.9941
R50 VP.n50 VP.n13 65.6004
R51 VP.n87 VP.n0 65.6004
R52 VP.n51 VP.n12 65.6004
R53 VP.n51 VP.n50 50.9766
R54 VP.n23 VP.n22 48.9289
R55 VP.n55 VP.n54 40.4934
R56 VP.n55 VP.n10 40.4934
R57 VP.n65 VP.n8 40.4934
R58 VP.n66 VP.n65 40.4934
R59 VP.n73 VP.n72 40.4934
R60 VP.n73 VP.n4 40.4934
R61 VP.n83 VP.n2 40.4934
R62 VP.n84 VP.n83 40.4934
R63 VP.n47 VP.n46 40.4934
R64 VP.n46 VP.n15 40.4934
R65 VP.n36 VP.n17 40.4934
R66 VP.n36 VP.n35 40.4934
R67 VP.n29 VP.n28 40.4934
R68 VP.n28 VP.n21 40.4934
R69 VP.n53 VP.n12 24.4675
R70 VP.n54 VP.n53 24.4675
R71 VP.n59 VP.n10 24.4675
R72 VP.n60 VP.n59 24.4675
R73 VP.n61 VP.n60 24.4675
R74 VP.n61 VP.n8 24.4675
R75 VP.n67 VP.n66 24.4675
R76 VP.n67 VP.n6 24.4675
R77 VP.n71 VP.n6 24.4675
R78 VP.n72 VP.n71 24.4675
R79 VP.n77 VP.n4 24.4675
R80 VP.n78 VP.n77 24.4675
R81 VP.n79 VP.n78 24.4675
R82 VP.n79 VP.n2 24.4675
R83 VP.n85 VP.n84 24.4675
R84 VP.n85 VP.n0 24.4675
R85 VP.n48 VP.n47 24.4675
R86 VP.n48 VP.n13 24.4675
R87 VP.n40 VP.n17 24.4675
R88 VP.n41 VP.n40 24.4675
R89 VP.n42 VP.n41 24.4675
R90 VP.n42 VP.n15 24.4675
R91 VP.n30 VP.n29 24.4675
R92 VP.n30 VP.n19 24.4675
R93 VP.n34 VP.n19 24.4675
R94 VP.n35 VP.n34 24.4675
R95 VP.n24 VP.n23 24.4675
R96 VP.n24 VP.n21 24.4675
R97 VP.n25 VP.n22 5.18913
R98 VP.n50 VP.n49 0.354971
R99 VP.n52 VP.n51 0.354971
R100 VP.n87 VP.n86 0.354971
R101 VP VP.n87 0.26696
R102 VP.n26 VP.n25 0.189894
R103 VP.n27 VP.n26 0.189894
R104 VP.n27 VP.n20 0.189894
R105 VP.n31 VP.n20 0.189894
R106 VP.n32 VP.n31 0.189894
R107 VP.n33 VP.n32 0.189894
R108 VP.n33 VP.n18 0.189894
R109 VP.n37 VP.n18 0.189894
R110 VP.n38 VP.n37 0.189894
R111 VP.n39 VP.n38 0.189894
R112 VP.n39 VP.n16 0.189894
R113 VP.n43 VP.n16 0.189894
R114 VP.n44 VP.n43 0.189894
R115 VP.n45 VP.n44 0.189894
R116 VP.n45 VP.n14 0.189894
R117 VP.n49 VP.n14 0.189894
R118 VP.n52 VP.n11 0.189894
R119 VP.n56 VP.n11 0.189894
R120 VP.n57 VP.n56 0.189894
R121 VP.n58 VP.n57 0.189894
R122 VP.n58 VP.n9 0.189894
R123 VP.n62 VP.n9 0.189894
R124 VP.n63 VP.n62 0.189894
R125 VP.n64 VP.n63 0.189894
R126 VP.n64 VP.n7 0.189894
R127 VP.n68 VP.n7 0.189894
R128 VP.n69 VP.n68 0.189894
R129 VP.n70 VP.n69 0.189894
R130 VP.n70 VP.n5 0.189894
R131 VP.n74 VP.n5 0.189894
R132 VP.n75 VP.n74 0.189894
R133 VP.n76 VP.n75 0.189894
R134 VP.n76 VP.n3 0.189894
R135 VP.n80 VP.n3 0.189894
R136 VP.n81 VP.n80 0.189894
R137 VP.n82 VP.n81 0.189894
R138 VP.n82 VP.n1 0.189894
R139 VP.n86 VP.n1 0.189894
R140 VTAIL.n192 VTAIL.n152 756.745
R141 VTAIL.n42 VTAIL.n2 756.745
R142 VTAIL.n146 VTAIL.n106 756.745
R143 VTAIL.n96 VTAIL.n56 756.745
R144 VTAIL.n167 VTAIL.n166 585
R145 VTAIL.n164 VTAIL.n163 585
R146 VTAIL.n173 VTAIL.n172 585
R147 VTAIL.n175 VTAIL.n174 585
R148 VTAIL.n160 VTAIL.n159 585
R149 VTAIL.n181 VTAIL.n180 585
R150 VTAIL.n184 VTAIL.n183 585
R151 VTAIL.n182 VTAIL.n156 585
R152 VTAIL.n189 VTAIL.n155 585
R153 VTAIL.n191 VTAIL.n190 585
R154 VTAIL.n193 VTAIL.n192 585
R155 VTAIL.n17 VTAIL.n16 585
R156 VTAIL.n14 VTAIL.n13 585
R157 VTAIL.n23 VTAIL.n22 585
R158 VTAIL.n25 VTAIL.n24 585
R159 VTAIL.n10 VTAIL.n9 585
R160 VTAIL.n31 VTAIL.n30 585
R161 VTAIL.n34 VTAIL.n33 585
R162 VTAIL.n32 VTAIL.n6 585
R163 VTAIL.n39 VTAIL.n5 585
R164 VTAIL.n41 VTAIL.n40 585
R165 VTAIL.n43 VTAIL.n42 585
R166 VTAIL.n147 VTAIL.n146 585
R167 VTAIL.n145 VTAIL.n144 585
R168 VTAIL.n143 VTAIL.n109 585
R169 VTAIL.n113 VTAIL.n110 585
R170 VTAIL.n138 VTAIL.n137 585
R171 VTAIL.n136 VTAIL.n135 585
R172 VTAIL.n115 VTAIL.n114 585
R173 VTAIL.n130 VTAIL.n129 585
R174 VTAIL.n128 VTAIL.n127 585
R175 VTAIL.n119 VTAIL.n118 585
R176 VTAIL.n122 VTAIL.n121 585
R177 VTAIL.n97 VTAIL.n96 585
R178 VTAIL.n95 VTAIL.n94 585
R179 VTAIL.n93 VTAIL.n59 585
R180 VTAIL.n63 VTAIL.n60 585
R181 VTAIL.n88 VTAIL.n87 585
R182 VTAIL.n86 VTAIL.n85 585
R183 VTAIL.n65 VTAIL.n64 585
R184 VTAIL.n80 VTAIL.n79 585
R185 VTAIL.n78 VTAIL.n77 585
R186 VTAIL.n69 VTAIL.n68 585
R187 VTAIL.n72 VTAIL.n71 585
R188 VTAIL.t12 VTAIL.n120 329.039
R189 VTAIL.t9 VTAIL.n70 329.039
R190 VTAIL.t6 VTAIL.n165 329.038
R191 VTAIL.t19 VTAIL.n15 329.038
R192 VTAIL.n166 VTAIL.n163 171.744
R193 VTAIL.n173 VTAIL.n163 171.744
R194 VTAIL.n174 VTAIL.n173 171.744
R195 VTAIL.n174 VTAIL.n159 171.744
R196 VTAIL.n181 VTAIL.n159 171.744
R197 VTAIL.n183 VTAIL.n181 171.744
R198 VTAIL.n183 VTAIL.n182 171.744
R199 VTAIL.n182 VTAIL.n155 171.744
R200 VTAIL.n191 VTAIL.n155 171.744
R201 VTAIL.n192 VTAIL.n191 171.744
R202 VTAIL.n16 VTAIL.n13 171.744
R203 VTAIL.n23 VTAIL.n13 171.744
R204 VTAIL.n24 VTAIL.n23 171.744
R205 VTAIL.n24 VTAIL.n9 171.744
R206 VTAIL.n31 VTAIL.n9 171.744
R207 VTAIL.n33 VTAIL.n31 171.744
R208 VTAIL.n33 VTAIL.n32 171.744
R209 VTAIL.n32 VTAIL.n5 171.744
R210 VTAIL.n41 VTAIL.n5 171.744
R211 VTAIL.n42 VTAIL.n41 171.744
R212 VTAIL.n146 VTAIL.n145 171.744
R213 VTAIL.n145 VTAIL.n109 171.744
R214 VTAIL.n113 VTAIL.n109 171.744
R215 VTAIL.n137 VTAIL.n113 171.744
R216 VTAIL.n137 VTAIL.n136 171.744
R217 VTAIL.n136 VTAIL.n114 171.744
R218 VTAIL.n129 VTAIL.n114 171.744
R219 VTAIL.n129 VTAIL.n128 171.744
R220 VTAIL.n128 VTAIL.n118 171.744
R221 VTAIL.n121 VTAIL.n118 171.744
R222 VTAIL.n96 VTAIL.n95 171.744
R223 VTAIL.n95 VTAIL.n59 171.744
R224 VTAIL.n63 VTAIL.n59 171.744
R225 VTAIL.n87 VTAIL.n63 171.744
R226 VTAIL.n87 VTAIL.n86 171.744
R227 VTAIL.n86 VTAIL.n64 171.744
R228 VTAIL.n79 VTAIL.n64 171.744
R229 VTAIL.n79 VTAIL.n78 171.744
R230 VTAIL.n78 VTAIL.n68 171.744
R231 VTAIL.n71 VTAIL.n68 171.744
R232 VTAIL.n166 VTAIL.t6 85.8723
R233 VTAIL.n16 VTAIL.t19 85.8723
R234 VTAIL.n121 VTAIL.t12 85.8723
R235 VTAIL.n71 VTAIL.t9 85.8723
R236 VTAIL.n105 VTAIL.n104 63.8194
R237 VTAIL.n103 VTAIL.n102 63.8194
R238 VTAIL.n55 VTAIL.n54 63.8194
R239 VTAIL.n53 VTAIL.n52 63.8194
R240 VTAIL.n199 VTAIL.n198 63.8192
R241 VTAIL.n1 VTAIL.n0 63.8192
R242 VTAIL.n49 VTAIL.n48 63.8192
R243 VTAIL.n51 VTAIL.n50 63.8192
R244 VTAIL.n197 VTAIL.n196 32.3793
R245 VTAIL.n47 VTAIL.n46 32.3793
R246 VTAIL.n151 VTAIL.n150 32.3793
R247 VTAIL.n101 VTAIL.n100 32.3793
R248 VTAIL.n53 VTAIL.n51 24.8927
R249 VTAIL.n197 VTAIL.n151 22.3065
R250 VTAIL.n190 VTAIL.n189 13.1884
R251 VTAIL.n40 VTAIL.n39 13.1884
R252 VTAIL.n144 VTAIL.n143 13.1884
R253 VTAIL.n94 VTAIL.n93 13.1884
R254 VTAIL.n188 VTAIL.n156 12.8005
R255 VTAIL.n193 VTAIL.n154 12.8005
R256 VTAIL.n38 VTAIL.n6 12.8005
R257 VTAIL.n43 VTAIL.n4 12.8005
R258 VTAIL.n147 VTAIL.n108 12.8005
R259 VTAIL.n142 VTAIL.n110 12.8005
R260 VTAIL.n97 VTAIL.n58 12.8005
R261 VTAIL.n92 VTAIL.n60 12.8005
R262 VTAIL.n185 VTAIL.n184 12.0247
R263 VTAIL.n194 VTAIL.n152 12.0247
R264 VTAIL.n35 VTAIL.n34 12.0247
R265 VTAIL.n44 VTAIL.n2 12.0247
R266 VTAIL.n148 VTAIL.n106 12.0247
R267 VTAIL.n139 VTAIL.n138 12.0247
R268 VTAIL.n98 VTAIL.n56 12.0247
R269 VTAIL.n89 VTAIL.n88 12.0247
R270 VTAIL.n180 VTAIL.n158 11.249
R271 VTAIL.n30 VTAIL.n8 11.249
R272 VTAIL.n135 VTAIL.n112 11.249
R273 VTAIL.n85 VTAIL.n62 11.249
R274 VTAIL.n167 VTAIL.n165 10.7239
R275 VTAIL.n17 VTAIL.n15 10.7239
R276 VTAIL.n122 VTAIL.n120 10.7239
R277 VTAIL.n72 VTAIL.n70 10.7239
R278 VTAIL.n179 VTAIL.n160 10.4732
R279 VTAIL.n29 VTAIL.n10 10.4732
R280 VTAIL.n134 VTAIL.n115 10.4732
R281 VTAIL.n84 VTAIL.n65 10.4732
R282 VTAIL.n176 VTAIL.n175 9.69747
R283 VTAIL.n26 VTAIL.n25 9.69747
R284 VTAIL.n131 VTAIL.n130 9.69747
R285 VTAIL.n81 VTAIL.n80 9.69747
R286 VTAIL.n196 VTAIL.n195 9.45567
R287 VTAIL.n46 VTAIL.n45 9.45567
R288 VTAIL.n150 VTAIL.n149 9.45567
R289 VTAIL.n100 VTAIL.n99 9.45567
R290 VTAIL.n195 VTAIL.n194 9.3005
R291 VTAIL.n154 VTAIL.n153 9.3005
R292 VTAIL.n169 VTAIL.n168 9.3005
R293 VTAIL.n171 VTAIL.n170 9.3005
R294 VTAIL.n162 VTAIL.n161 9.3005
R295 VTAIL.n177 VTAIL.n176 9.3005
R296 VTAIL.n179 VTAIL.n178 9.3005
R297 VTAIL.n158 VTAIL.n157 9.3005
R298 VTAIL.n186 VTAIL.n185 9.3005
R299 VTAIL.n188 VTAIL.n187 9.3005
R300 VTAIL.n45 VTAIL.n44 9.3005
R301 VTAIL.n4 VTAIL.n3 9.3005
R302 VTAIL.n19 VTAIL.n18 9.3005
R303 VTAIL.n21 VTAIL.n20 9.3005
R304 VTAIL.n12 VTAIL.n11 9.3005
R305 VTAIL.n27 VTAIL.n26 9.3005
R306 VTAIL.n29 VTAIL.n28 9.3005
R307 VTAIL.n8 VTAIL.n7 9.3005
R308 VTAIL.n36 VTAIL.n35 9.3005
R309 VTAIL.n38 VTAIL.n37 9.3005
R310 VTAIL.n124 VTAIL.n123 9.3005
R311 VTAIL.n126 VTAIL.n125 9.3005
R312 VTAIL.n117 VTAIL.n116 9.3005
R313 VTAIL.n132 VTAIL.n131 9.3005
R314 VTAIL.n134 VTAIL.n133 9.3005
R315 VTAIL.n112 VTAIL.n111 9.3005
R316 VTAIL.n140 VTAIL.n139 9.3005
R317 VTAIL.n142 VTAIL.n141 9.3005
R318 VTAIL.n149 VTAIL.n148 9.3005
R319 VTAIL.n108 VTAIL.n107 9.3005
R320 VTAIL.n74 VTAIL.n73 9.3005
R321 VTAIL.n76 VTAIL.n75 9.3005
R322 VTAIL.n67 VTAIL.n66 9.3005
R323 VTAIL.n82 VTAIL.n81 9.3005
R324 VTAIL.n84 VTAIL.n83 9.3005
R325 VTAIL.n62 VTAIL.n61 9.3005
R326 VTAIL.n90 VTAIL.n89 9.3005
R327 VTAIL.n92 VTAIL.n91 9.3005
R328 VTAIL.n99 VTAIL.n98 9.3005
R329 VTAIL.n58 VTAIL.n57 9.3005
R330 VTAIL.n172 VTAIL.n162 8.92171
R331 VTAIL.n22 VTAIL.n12 8.92171
R332 VTAIL.n127 VTAIL.n117 8.92171
R333 VTAIL.n77 VTAIL.n67 8.92171
R334 VTAIL.n171 VTAIL.n164 8.14595
R335 VTAIL.n21 VTAIL.n14 8.14595
R336 VTAIL.n126 VTAIL.n119 8.14595
R337 VTAIL.n76 VTAIL.n69 8.14595
R338 VTAIL.n168 VTAIL.n167 7.3702
R339 VTAIL.n18 VTAIL.n17 7.3702
R340 VTAIL.n123 VTAIL.n122 7.3702
R341 VTAIL.n73 VTAIL.n72 7.3702
R342 VTAIL.n168 VTAIL.n164 5.81868
R343 VTAIL.n18 VTAIL.n14 5.81868
R344 VTAIL.n123 VTAIL.n119 5.81868
R345 VTAIL.n73 VTAIL.n69 5.81868
R346 VTAIL.n172 VTAIL.n171 5.04292
R347 VTAIL.n22 VTAIL.n21 5.04292
R348 VTAIL.n127 VTAIL.n126 5.04292
R349 VTAIL.n77 VTAIL.n76 5.04292
R350 VTAIL.n175 VTAIL.n162 4.26717
R351 VTAIL.n25 VTAIL.n12 4.26717
R352 VTAIL.n130 VTAIL.n117 4.26717
R353 VTAIL.n80 VTAIL.n67 4.26717
R354 VTAIL.n198 VTAIL.t0 3.81117
R355 VTAIL.n198 VTAIL.t1 3.81117
R356 VTAIL.n0 VTAIL.t8 3.81117
R357 VTAIL.n0 VTAIL.t4 3.81117
R358 VTAIL.n48 VTAIL.t17 3.81117
R359 VTAIL.n48 VTAIL.t14 3.81117
R360 VTAIL.n50 VTAIL.t18 3.81117
R361 VTAIL.n50 VTAIL.t15 3.81117
R362 VTAIL.n104 VTAIL.t10 3.81117
R363 VTAIL.n104 VTAIL.t11 3.81117
R364 VTAIL.n102 VTAIL.t16 3.81117
R365 VTAIL.n102 VTAIL.t13 3.81117
R366 VTAIL.n54 VTAIL.t7 3.81117
R367 VTAIL.n54 VTAIL.t3 3.81117
R368 VTAIL.n52 VTAIL.t5 3.81117
R369 VTAIL.n52 VTAIL.t2 3.81117
R370 VTAIL.n176 VTAIL.n160 3.49141
R371 VTAIL.n26 VTAIL.n10 3.49141
R372 VTAIL.n131 VTAIL.n115 3.49141
R373 VTAIL.n81 VTAIL.n65 3.49141
R374 VTAIL.n180 VTAIL.n179 2.71565
R375 VTAIL.n30 VTAIL.n29 2.71565
R376 VTAIL.n135 VTAIL.n134 2.71565
R377 VTAIL.n85 VTAIL.n84 2.71565
R378 VTAIL.n55 VTAIL.n53 2.58671
R379 VTAIL.n101 VTAIL.n55 2.58671
R380 VTAIL.n105 VTAIL.n103 2.58671
R381 VTAIL.n151 VTAIL.n105 2.58671
R382 VTAIL.n51 VTAIL.n49 2.58671
R383 VTAIL.n49 VTAIL.n47 2.58671
R384 VTAIL.n199 VTAIL.n197 2.58671
R385 VTAIL.n169 VTAIL.n165 2.41285
R386 VTAIL.n19 VTAIL.n15 2.41285
R387 VTAIL.n124 VTAIL.n120 2.41285
R388 VTAIL.n74 VTAIL.n70 2.41285
R389 VTAIL VTAIL.n1 1.99834
R390 VTAIL.n184 VTAIL.n158 1.93989
R391 VTAIL.n196 VTAIL.n152 1.93989
R392 VTAIL.n34 VTAIL.n8 1.93989
R393 VTAIL.n46 VTAIL.n2 1.93989
R394 VTAIL.n150 VTAIL.n106 1.93989
R395 VTAIL.n138 VTAIL.n112 1.93989
R396 VTAIL.n100 VTAIL.n56 1.93989
R397 VTAIL.n88 VTAIL.n62 1.93989
R398 VTAIL.n103 VTAIL.n101 1.76343
R399 VTAIL.n47 VTAIL.n1 1.76343
R400 VTAIL.n185 VTAIL.n156 1.16414
R401 VTAIL.n194 VTAIL.n193 1.16414
R402 VTAIL.n35 VTAIL.n6 1.16414
R403 VTAIL.n44 VTAIL.n43 1.16414
R404 VTAIL.n148 VTAIL.n147 1.16414
R405 VTAIL.n139 VTAIL.n110 1.16414
R406 VTAIL.n98 VTAIL.n97 1.16414
R407 VTAIL.n89 VTAIL.n60 1.16414
R408 VTAIL VTAIL.n199 0.588862
R409 VTAIL.n189 VTAIL.n188 0.388379
R410 VTAIL.n190 VTAIL.n154 0.388379
R411 VTAIL.n39 VTAIL.n38 0.388379
R412 VTAIL.n40 VTAIL.n4 0.388379
R413 VTAIL.n144 VTAIL.n108 0.388379
R414 VTAIL.n143 VTAIL.n142 0.388379
R415 VTAIL.n94 VTAIL.n58 0.388379
R416 VTAIL.n93 VTAIL.n92 0.388379
R417 VTAIL.n170 VTAIL.n169 0.155672
R418 VTAIL.n170 VTAIL.n161 0.155672
R419 VTAIL.n177 VTAIL.n161 0.155672
R420 VTAIL.n178 VTAIL.n177 0.155672
R421 VTAIL.n178 VTAIL.n157 0.155672
R422 VTAIL.n186 VTAIL.n157 0.155672
R423 VTAIL.n187 VTAIL.n186 0.155672
R424 VTAIL.n187 VTAIL.n153 0.155672
R425 VTAIL.n195 VTAIL.n153 0.155672
R426 VTAIL.n20 VTAIL.n19 0.155672
R427 VTAIL.n20 VTAIL.n11 0.155672
R428 VTAIL.n27 VTAIL.n11 0.155672
R429 VTAIL.n28 VTAIL.n27 0.155672
R430 VTAIL.n28 VTAIL.n7 0.155672
R431 VTAIL.n36 VTAIL.n7 0.155672
R432 VTAIL.n37 VTAIL.n36 0.155672
R433 VTAIL.n37 VTAIL.n3 0.155672
R434 VTAIL.n45 VTAIL.n3 0.155672
R435 VTAIL.n149 VTAIL.n107 0.155672
R436 VTAIL.n141 VTAIL.n107 0.155672
R437 VTAIL.n141 VTAIL.n140 0.155672
R438 VTAIL.n140 VTAIL.n111 0.155672
R439 VTAIL.n133 VTAIL.n111 0.155672
R440 VTAIL.n133 VTAIL.n132 0.155672
R441 VTAIL.n132 VTAIL.n116 0.155672
R442 VTAIL.n125 VTAIL.n116 0.155672
R443 VTAIL.n125 VTAIL.n124 0.155672
R444 VTAIL.n99 VTAIL.n57 0.155672
R445 VTAIL.n91 VTAIL.n57 0.155672
R446 VTAIL.n91 VTAIL.n90 0.155672
R447 VTAIL.n90 VTAIL.n61 0.155672
R448 VTAIL.n83 VTAIL.n61 0.155672
R449 VTAIL.n83 VTAIL.n82 0.155672
R450 VTAIL.n82 VTAIL.n66 0.155672
R451 VTAIL.n75 VTAIL.n66 0.155672
R452 VTAIL.n75 VTAIL.n74 0.155672
R453 VDD1.n40 VDD1.n0 756.745
R454 VDD1.n87 VDD1.n47 756.745
R455 VDD1.n41 VDD1.n40 585
R456 VDD1.n39 VDD1.n38 585
R457 VDD1.n37 VDD1.n3 585
R458 VDD1.n7 VDD1.n4 585
R459 VDD1.n32 VDD1.n31 585
R460 VDD1.n30 VDD1.n29 585
R461 VDD1.n9 VDD1.n8 585
R462 VDD1.n24 VDD1.n23 585
R463 VDD1.n22 VDD1.n21 585
R464 VDD1.n13 VDD1.n12 585
R465 VDD1.n16 VDD1.n15 585
R466 VDD1.n62 VDD1.n61 585
R467 VDD1.n59 VDD1.n58 585
R468 VDD1.n68 VDD1.n67 585
R469 VDD1.n70 VDD1.n69 585
R470 VDD1.n55 VDD1.n54 585
R471 VDD1.n76 VDD1.n75 585
R472 VDD1.n79 VDD1.n78 585
R473 VDD1.n77 VDD1.n51 585
R474 VDD1.n84 VDD1.n50 585
R475 VDD1.n86 VDD1.n85 585
R476 VDD1.n88 VDD1.n87 585
R477 VDD1.t2 VDD1.n14 329.039
R478 VDD1.t4 VDD1.n60 329.038
R479 VDD1.n40 VDD1.n39 171.744
R480 VDD1.n39 VDD1.n3 171.744
R481 VDD1.n7 VDD1.n3 171.744
R482 VDD1.n31 VDD1.n7 171.744
R483 VDD1.n31 VDD1.n30 171.744
R484 VDD1.n30 VDD1.n8 171.744
R485 VDD1.n23 VDD1.n8 171.744
R486 VDD1.n23 VDD1.n22 171.744
R487 VDD1.n22 VDD1.n12 171.744
R488 VDD1.n15 VDD1.n12 171.744
R489 VDD1.n61 VDD1.n58 171.744
R490 VDD1.n68 VDD1.n58 171.744
R491 VDD1.n69 VDD1.n68 171.744
R492 VDD1.n69 VDD1.n54 171.744
R493 VDD1.n76 VDD1.n54 171.744
R494 VDD1.n78 VDD1.n76 171.744
R495 VDD1.n78 VDD1.n77 171.744
R496 VDD1.n77 VDD1.n50 171.744
R497 VDD1.n86 VDD1.n50 171.744
R498 VDD1.n87 VDD1.n86 171.744
R499 VDD1.n15 VDD1.t2 85.8723
R500 VDD1.n61 VDD1.t4 85.8723
R501 VDD1.n95 VDD1.n94 82.3823
R502 VDD1.n46 VDD1.n45 80.4982
R503 VDD1.n97 VDD1.n96 80.498
R504 VDD1.n93 VDD1.n92 80.498
R505 VDD1.n46 VDD1.n44 51.6443
R506 VDD1.n93 VDD1.n91 51.6443
R507 VDD1.n97 VDD1.n95 45.2293
R508 VDD1.n38 VDD1.n37 13.1884
R509 VDD1.n85 VDD1.n84 13.1884
R510 VDD1.n41 VDD1.n2 12.8005
R511 VDD1.n36 VDD1.n4 12.8005
R512 VDD1.n83 VDD1.n51 12.8005
R513 VDD1.n88 VDD1.n49 12.8005
R514 VDD1.n42 VDD1.n0 12.0247
R515 VDD1.n33 VDD1.n32 12.0247
R516 VDD1.n80 VDD1.n79 12.0247
R517 VDD1.n89 VDD1.n47 12.0247
R518 VDD1.n29 VDD1.n6 11.249
R519 VDD1.n75 VDD1.n53 11.249
R520 VDD1.n16 VDD1.n14 10.7239
R521 VDD1.n62 VDD1.n60 10.7239
R522 VDD1.n28 VDD1.n9 10.4732
R523 VDD1.n74 VDD1.n55 10.4732
R524 VDD1.n25 VDD1.n24 9.69747
R525 VDD1.n71 VDD1.n70 9.69747
R526 VDD1.n44 VDD1.n43 9.45567
R527 VDD1.n91 VDD1.n90 9.45567
R528 VDD1.n18 VDD1.n17 9.3005
R529 VDD1.n20 VDD1.n19 9.3005
R530 VDD1.n11 VDD1.n10 9.3005
R531 VDD1.n26 VDD1.n25 9.3005
R532 VDD1.n28 VDD1.n27 9.3005
R533 VDD1.n6 VDD1.n5 9.3005
R534 VDD1.n34 VDD1.n33 9.3005
R535 VDD1.n36 VDD1.n35 9.3005
R536 VDD1.n43 VDD1.n42 9.3005
R537 VDD1.n2 VDD1.n1 9.3005
R538 VDD1.n90 VDD1.n89 9.3005
R539 VDD1.n49 VDD1.n48 9.3005
R540 VDD1.n64 VDD1.n63 9.3005
R541 VDD1.n66 VDD1.n65 9.3005
R542 VDD1.n57 VDD1.n56 9.3005
R543 VDD1.n72 VDD1.n71 9.3005
R544 VDD1.n74 VDD1.n73 9.3005
R545 VDD1.n53 VDD1.n52 9.3005
R546 VDD1.n81 VDD1.n80 9.3005
R547 VDD1.n83 VDD1.n82 9.3005
R548 VDD1.n21 VDD1.n11 8.92171
R549 VDD1.n67 VDD1.n57 8.92171
R550 VDD1.n20 VDD1.n13 8.14595
R551 VDD1.n66 VDD1.n59 8.14595
R552 VDD1.n17 VDD1.n16 7.3702
R553 VDD1.n63 VDD1.n62 7.3702
R554 VDD1.n17 VDD1.n13 5.81868
R555 VDD1.n63 VDD1.n59 5.81868
R556 VDD1.n21 VDD1.n20 5.04292
R557 VDD1.n67 VDD1.n66 5.04292
R558 VDD1.n24 VDD1.n11 4.26717
R559 VDD1.n70 VDD1.n57 4.26717
R560 VDD1.n96 VDD1.t8 3.81117
R561 VDD1.n96 VDD1.t9 3.81117
R562 VDD1.n45 VDD1.t1 3.81117
R563 VDD1.n45 VDD1.t7 3.81117
R564 VDD1.n94 VDD1.t5 3.81117
R565 VDD1.n94 VDD1.t0 3.81117
R566 VDD1.n92 VDD1.t6 3.81117
R567 VDD1.n92 VDD1.t3 3.81117
R568 VDD1.n25 VDD1.n9 3.49141
R569 VDD1.n71 VDD1.n55 3.49141
R570 VDD1.n29 VDD1.n28 2.71565
R571 VDD1.n75 VDD1.n74 2.71565
R572 VDD1.n18 VDD1.n14 2.41285
R573 VDD1.n64 VDD1.n60 2.41285
R574 VDD1.n44 VDD1.n0 1.93989
R575 VDD1.n32 VDD1.n6 1.93989
R576 VDD1.n79 VDD1.n53 1.93989
R577 VDD1.n91 VDD1.n47 1.93989
R578 VDD1 VDD1.n97 1.88197
R579 VDD1.n42 VDD1.n41 1.16414
R580 VDD1.n33 VDD1.n4 1.16414
R581 VDD1.n80 VDD1.n51 1.16414
R582 VDD1.n89 VDD1.n88 1.16414
R583 VDD1 VDD1.n46 0.705241
R584 VDD1.n95 VDD1.n93 0.591706
R585 VDD1.n38 VDD1.n2 0.388379
R586 VDD1.n37 VDD1.n36 0.388379
R587 VDD1.n84 VDD1.n83 0.388379
R588 VDD1.n85 VDD1.n49 0.388379
R589 VDD1.n43 VDD1.n1 0.155672
R590 VDD1.n35 VDD1.n1 0.155672
R591 VDD1.n35 VDD1.n34 0.155672
R592 VDD1.n34 VDD1.n5 0.155672
R593 VDD1.n27 VDD1.n5 0.155672
R594 VDD1.n27 VDD1.n26 0.155672
R595 VDD1.n26 VDD1.n10 0.155672
R596 VDD1.n19 VDD1.n10 0.155672
R597 VDD1.n19 VDD1.n18 0.155672
R598 VDD1.n65 VDD1.n64 0.155672
R599 VDD1.n65 VDD1.n56 0.155672
R600 VDD1.n72 VDD1.n56 0.155672
R601 VDD1.n73 VDD1.n72 0.155672
R602 VDD1.n73 VDD1.n52 0.155672
R603 VDD1.n81 VDD1.n52 0.155672
R604 VDD1.n82 VDD1.n81 0.155672
R605 VDD1.n82 VDD1.n48 0.155672
R606 VDD1.n90 VDD1.n48 0.155672
R607 VN.n74 VN.n73 161.3
R608 VN.n72 VN.n39 161.3
R609 VN.n71 VN.n70 161.3
R610 VN.n69 VN.n40 161.3
R611 VN.n68 VN.n67 161.3
R612 VN.n66 VN.n41 161.3
R613 VN.n65 VN.n64 161.3
R614 VN.n63 VN.n42 161.3
R615 VN.n62 VN.n61 161.3
R616 VN.n60 VN.n43 161.3
R617 VN.n59 VN.n58 161.3
R618 VN.n57 VN.n44 161.3
R619 VN.n56 VN.n55 161.3
R620 VN.n54 VN.n45 161.3
R621 VN.n53 VN.n52 161.3
R622 VN.n51 VN.n46 161.3
R623 VN.n50 VN.n49 161.3
R624 VN.n36 VN.n35 161.3
R625 VN.n34 VN.n1 161.3
R626 VN.n33 VN.n32 161.3
R627 VN.n31 VN.n2 161.3
R628 VN.n30 VN.n29 161.3
R629 VN.n28 VN.n3 161.3
R630 VN.n27 VN.n26 161.3
R631 VN.n25 VN.n4 161.3
R632 VN.n24 VN.n23 161.3
R633 VN.n22 VN.n5 161.3
R634 VN.n21 VN.n20 161.3
R635 VN.n19 VN.n6 161.3
R636 VN.n18 VN.n17 161.3
R637 VN.n16 VN.n7 161.3
R638 VN.n15 VN.n14 161.3
R639 VN.n13 VN.n8 161.3
R640 VN.n12 VN.n11 161.3
R641 VN.n9 VN.t8 109.144
R642 VN.n47 VN.t5 109.144
R643 VN.n0 VN.t4 76.9941
R644 VN.n28 VN.t1 76.9941
R645 VN.n6 VN.t7 76.9941
R646 VN.n10 VN.t3 76.9941
R647 VN.n38 VN.t0 76.9941
R648 VN.n66 VN.t2 76.9941
R649 VN.n44 VN.t9 76.9941
R650 VN.n48 VN.t6 76.9941
R651 VN.n75 VN.n38 65.6004
R652 VN.n37 VN.n0 65.6004
R653 VN VN.n75 51.142
R654 VN.n48 VN.n47 48.9288
R655 VN.n10 VN.n9 48.9288
R656 VN.n15 VN.n8 40.4934
R657 VN.n16 VN.n15 40.4934
R658 VN.n23 VN.n22 40.4934
R659 VN.n23 VN.n4 40.4934
R660 VN.n33 VN.n2 40.4934
R661 VN.n34 VN.n33 40.4934
R662 VN.n53 VN.n46 40.4934
R663 VN.n54 VN.n53 40.4934
R664 VN.n61 VN.n60 40.4934
R665 VN.n61 VN.n42 40.4934
R666 VN.n71 VN.n40 40.4934
R667 VN.n72 VN.n71 40.4934
R668 VN.n11 VN.n10 24.4675
R669 VN.n11 VN.n8 24.4675
R670 VN.n17 VN.n16 24.4675
R671 VN.n17 VN.n6 24.4675
R672 VN.n21 VN.n6 24.4675
R673 VN.n22 VN.n21 24.4675
R674 VN.n27 VN.n4 24.4675
R675 VN.n28 VN.n27 24.4675
R676 VN.n29 VN.n28 24.4675
R677 VN.n29 VN.n2 24.4675
R678 VN.n35 VN.n34 24.4675
R679 VN.n35 VN.n0 24.4675
R680 VN.n49 VN.n46 24.4675
R681 VN.n49 VN.n48 24.4675
R682 VN.n60 VN.n59 24.4675
R683 VN.n59 VN.n44 24.4675
R684 VN.n55 VN.n44 24.4675
R685 VN.n55 VN.n54 24.4675
R686 VN.n67 VN.n40 24.4675
R687 VN.n67 VN.n66 24.4675
R688 VN.n66 VN.n65 24.4675
R689 VN.n65 VN.n42 24.4675
R690 VN.n73 VN.n38 24.4675
R691 VN.n73 VN.n72 24.4675
R692 VN.n50 VN.n47 5.18917
R693 VN.n12 VN.n9 5.18917
R694 VN.n75 VN.n74 0.354971
R695 VN.n37 VN.n36 0.354971
R696 VN VN.n37 0.26696
R697 VN.n74 VN.n39 0.189894
R698 VN.n70 VN.n39 0.189894
R699 VN.n70 VN.n69 0.189894
R700 VN.n69 VN.n68 0.189894
R701 VN.n68 VN.n41 0.189894
R702 VN.n64 VN.n41 0.189894
R703 VN.n64 VN.n63 0.189894
R704 VN.n63 VN.n62 0.189894
R705 VN.n62 VN.n43 0.189894
R706 VN.n58 VN.n43 0.189894
R707 VN.n58 VN.n57 0.189894
R708 VN.n57 VN.n56 0.189894
R709 VN.n56 VN.n45 0.189894
R710 VN.n52 VN.n45 0.189894
R711 VN.n52 VN.n51 0.189894
R712 VN.n51 VN.n50 0.189894
R713 VN.n13 VN.n12 0.189894
R714 VN.n14 VN.n13 0.189894
R715 VN.n14 VN.n7 0.189894
R716 VN.n18 VN.n7 0.189894
R717 VN.n19 VN.n18 0.189894
R718 VN.n20 VN.n19 0.189894
R719 VN.n20 VN.n5 0.189894
R720 VN.n24 VN.n5 0.189894
R721 VN.n25 VN.n24 0.189894
R722 VN.n26 VN.n25 0.189894
R723 VN.n26 VN.n3 0.189894
R724 VN.n30 VN.n3 0.189894
R725 VN.n31 VN.n30 0.189894
R726 VN.n32 VN.n31 0.189894
R727 VN.n32 VN.n1 0.189894
R728 VN.n36 VN.n1 0.189894
R729 VDD2.n89 VDD2.n49 756.745
R730 VDD2.n40 VDD2.n0 756.745
R731 VDD2.n90 VDD2.n89 585
R732 VDD2.n88 VDD2.n87 585
R733 VDD2.n86 VDD2.n52 585
R734 VDD2.n56 VDD2.n53 585
R735 VDD2.n81 VDD2.n80 585
R736 VDD2.n79 VDD2.n78 585
R737 VDD2.n58 VDD2.n57 585
R738 VDD2.n73 VDD2.n72 585
R739 VDD2.n71 VDD2.n70 585
R740 VDD2.n62 VDD2.n61 585
R741 VDD2.n65 VDD2.n64 585
R742 VDD2.n15 VDD2.n14 585
R743 VDD2.n12 VDD2.n11 585
R744 VDD2.n21 VDD2.n20 585
R745 VDD2.n23 VDD2.n22 585
R746 VDD2.n8 VDD2.n7 585
R747 VDD2.n29 VDD2.n28 585
R748 VDD2.n32 VDD2.n31 585
R749 VDD2.n30 VDD2.n4 585
R750 VDD2.n37 VDD2.n3 585
R751 VDD2.n39 VDD2.n38 585
R752 VDD2.n41 VDD2.n40 585
R753 VDD2.t9 VDD2.n63 329.039
R754 VDD2.t1 VDD2.n13 329.038
R755 VDD2.n89 VDD2.n88 171.744
R756 VDD2.n88 VDD2.n52 171.744
R757 VDD2.n56 VDD2.n52 171.744
R758 VDD2.n80 VDD2.n56 171.744
R759 VDD2.n80 VDD2.n79 171.744
R760 VDD2.n79 VDD2.n57 171.744
R761 VDD2.n72 VDD2.n57 171.744
R762 VDD2.n72 VDD2.n71 171.744
R763 VDD2.n71 VDD2.n61 171.744
R764 VDD2.n64 VDD2.n61 171.744
R765 VDD2.n14 VDD2.n11 171.744
R766 VDD2.n21 VDD2.n11 171.744
R767 VDD2.n22 VDD2.n21 171.744
R768 VDD2.n22 VDD2.n7 171.744
R769 VDD2.n29 VDD2.n7 171.744
R770 VDD2.n31 VDD2.n29 171.744
R771 VDD2.n31 VDD2.n30 171.744
R772 VDD2.n30 VDD2.n3 171.744
R773 VDD2.n39 VDD2.n3 171.744
R774 VDD2.n40 VDD2.n39 171.744
R775 VDD2.n64 VDD2.t9 85.8723
R776 VDD2.n14 VDD2.t1 85.8723
R777 VDD2.n48 VDD2.n47 82.3823
R778 VDD2 VDD2.n97 82.3795
R779 VDD2.n96 VDD2.n95 80.4982
R780 VDD2.n46 VDD2.n45 80.498
R781 VDD2.n46 VDD2.n44 51.6443
R782 VDD2.n94 VDD2.n93 49.0581
R783 VDD2.n94 VDD2.n48 43.3532
R784 VDD2.n87 VDD2.n86 13.1884
R785 VDD2.n38 VDD2.n37 13.1884
R786 VDD2.n90 VDD2.n51 12.8005
R787 VDD2.n85 VDD2.n53 12.8005
R788 VDD2.n36 VDD2.n4 12.8005
R789 VDD2.n41 VDD2.n2 12.8005
R790 VDD2.n91 VDD2.n49 12.0247
R791 VDD2.n82 VDD2.n81 12.0247
R792 VDD2.n33 VDD2.n32 12.0247
R793 VDD2.n42 VDD2.n0 12.0247
R794 VDD2.n78 VDD2.n55 11.249
R795 VDD2.n28 VDD2.n6 11.249
R796 VDD2.n65 VDD2.n63 10.7239
R797 VDD2.n15 VDD2.n13 10.7239
R798 VDD2.n77 VDD2.n58 10.4732
R799 VDD2.n27 VDD2.n8 10.4732
R800 VDD2.n74 VDD2.n73 9.69747
R801 VDD2.n24 VDD2.n23 9.69747
R802 VDD2.n93 VDD2.n92 9.45567
R803 VDD2.n44 VDD2.n43 9.45567
R804 VDD2.n67 VDD2.n66 9.3005
R805 VDD2.n69 VDD2.n68 9.3005
R806 VDD2.n60 VDD2.n59 9.3005
R807 VDD2.n75 VDD2.n74 9.3005
R808 VDD2.n77 VDD2.n76 9.3005
R809 VDD2.n55 VDD2.n54 9.3005
R810 VDD2.n83 VDD2.n82 9.3005
R811 VDD2.n85 VDD2.n84 9.3005
R812 VDD2.n92 VDD2.n91 9.3005
R813 VDD2.n51 VDD2.n50 9.3005
R814 VDD2.n43 VDD2.n42 9.3005
R815 VDD2.n2 VDD2.n1 9.3005
R816 VDD2.n17 VDD2.n16 9.3005
R817 VDD2.n19 VDD2.n18 9.3005
R818 VDD2.n10 VDD2.n9 9.3005
R819 VDD2.n25 VDD2.n24 9.3005
R820 VDD2.n27 VDD2.n26 9.3005
R821 VDD2.n6 VDD2.n5 9.3005
R822 VDD2.n34 VDD2.n33 9.3005
R823 VDD2.n36 VDD2.n35 9.3005
R824 VDD2.n70 VDD2.n60 8.92171
R825 VDD2.n20 VDD2.n10 8.92171
R826 VDD2.n69 VDD2.n62 8.14595
R827 VDD2.n19 VDD2.n12 8.14595
R828 VDD2.n66 VDD2.n65 7.3702
R829 VDD2.n16 VDD2.n15 7.3702
R830 VDD2.n66 VDD2.n62 5.81868
R831 VDD2.n16 VDD2.n12 5.81868
R832 VDD2.n70 VDD2.n69 5.04292
R833 VDD2.n20 VDD2.n19 5.04292
R834 VDD2.n73 VDD2.n60 4.26717
R835 VDD2.n23 VDD2.n10 4.26717
R836 VDD2.n97 VDD2.t3 3.81117
R837 VDD2.n97 VDD2.t4 3.81117
R838 VDD2.n95 VDD2.t7 3.81117
R839 VDD2.n95 VDD2.t0 3.81117
R840 VDD2.n47 VDD2.t8 3.81117
R841 VDD2.n47 VDD2.t5 3.81117
R842 VDD2.n45 VDD2.t6 3.81117
R843 VDD2.n45 VDD2.t2 3.81117
R844 VDD2.n74 VDD2.n58 3.49141
R845 VDD2.n24 VDD2.n8 3.49141
R846 VDD2.n78 VDD2.n77 2.71565
R847 VDD2.n28 VDD2.n27 2.71565
R848 VDD2.n96 VDD2.n94 2.58671
R849 VDD2.n67 VDD2.n63 2.41285
R850 VDD2.n17 VDD2.n13 2.41285
R851 VDD2.n93 VDD2.n49 1.93989
R852 VDD2.n81 VDD2.n55 1.93989
R853 VDD2.n32 VDD2.n6 1.93989
R854 VDD2.n44 VDD2.n0 1.93989
R855 VDD2.n91 VDD2.n90 1.16414
R856 VDD2.n82 VDD2.n53 1.16414
R857 VDD2.n33 VDD2.n4 1.16414
R858 VDD2.n42 VDD2.n41 1.16414
R859 VDD2 VDD2.n96 0.705241
R860 VDD2.n48 VDD2.n46 0.591706
R861 VDD2.n87 VDD2.n51 0.388379
R862 VDD2.n86 VDD2.n85 0.388379
R863 VDD2.n37 VDD2.n36 0.388379
R864 VDD2.n38 VDD2.n2 0.388379
R865 VDD2.n92 VDD2.n50 0.155672
R866 VDD2.n84 VDD2.n50 0.155672
R867 VDD2.n84 VDD2.n83 0.155672
R868 VDD2.n83 VDD2.n54 0.155672
R869 VDD2.n76 VDD2.n54 0.155672
R870 VDD2.n76 VDD2.n75 0.155672
R871 VDD2.n75 VDD2.n59 0.155672
R872 VDD2.n68 VDD2.n59 0.155672
R873 VDD2.n68 VDD2.n67 0.155672
R874 VDD2.n18 VDD2.n17 0.155672
R875 VDD2.n18 VDD2.n9 0.155672
R876 VDD2.n25 VDD2.n9 0.155672
R877 VDD2.n26 VDD2.n25 0.155672
R878 VDD2.n26 VDD2.n5 0.155672
R879 VDD2.n34 VDD2.n5 0.155672
R880 VDD2.n35 VDD2.n34 0.155672
R881 VDD2.n35 VDD2.n1 0.155672
R882 VDD2.n43 VDD2.n1 0.155672
R883 B.n590 B.n589 585
R884 B.n591 B.n72 585
R885 B.n593 B.n592 585
R886 B.n594 B.n71 585
R887 B.n596 B.n595 585
R888 B.n597 B.n70 585
R889 B.n599 B.n598 585
R890 B.n600 B.n69 585
R891 B.n602 B.n601 585
R892 B.n603 B.n68 585
R893 B.n605 B.n604 585
R894 B.n606 B.n67 585
R895 B.n608 B.n607 585
R896 B.n609 B.n66 585
R897 B.n611 B.n610 585
R898 B.n612 B.n65 585
R899 B.n614 B.n613 585
R900 B.n615 B.n64 585
R901 B.n617 B.n616 585
R902 B.n618 B.n63 585
R903 B.n620 B.n619 585
R904 B.n621 B.n62 585
R905 B.n623 B.n622 585
R906 B.n624 B.n61 585
R907 B.n626 B.n625 585
R908 B.n627 B.n60 585
R909 B.n629 B.n628 585
R910 B.n630 B.n59 585
R911 B.n632 B.n631 585
R912 B.n633 B.n58 585
R913 B.n635 B.n634 585
R914 B.n637 B.n55 585
R915 B.n639 B.n638 585
R916 B.n640 B.n54 585
R917 B.n642 B.n641 585
R918 B.n643 B.n53 585
R919 B.n645 B.n644 585
R920 B.n646 B.n52 585
R921 B.n648 B.n647 585
R922 B.n649 B.n51 585
R923 B.n651 B.n650 585
R924 B.n653 B.n652 585
R925 B.n654 B.n47 585
R926 B.n656 B.n655 585
R927 B.n657 B.n46 585
R928 B.n659 B.n658 585
R929 B.n660 B.n45 585
R930 B.n662 B.n661 585
R931 B.n663 B.n44 585
R932 B.n665 B.n664 585
R933 B.n666 B.n43 585
R934 B.n668 B.n667 585
R935 B.n669 B.n42 585
R936 B.n671 B.n670 585
R937 B.n672 B.n41 585
R938 B.n674 B.n673 585
R939 B.n675 B.n40 585
R940 B.n677 B.n676 585
R941 B.n678 B.n39 585
R942 B.n680 B.n679 585
R943 B.n681 B.n38 585
R944 B.n683 B.n682 585
R945 B.n684 B.n37 585
R946 B.n686 B.n685 585
R947 B.n687 B.n36 585
R948 B.n689 B.n688 585
R949 B.n690 B.n35 585
R950 B.n692 B.n691 585
R951 B.n693 B.n34 585
R952 B.n695 B.n694 585
R953 B.n696 B.n33 585
R954 B.n698 B.n697 585
R955 B.n588 B.n73 585
R956 B.n587 B.n586 585
R957 B.n585 B.n74 585
R958 B.n584 B.n583 585
R959 B.n582 B.n75 585
R960 B.n581 B.n580 585
R961 B.n579 B.n76 585
R962 B.n578 B.n577 585
R963 B.n576 B.n77 585
R964 B.n575 B.n574 585
R965 B.n573 B.n78 585
R966 B.n572 B.n571 585
R967 B.n570 B.n79 585
R968 B.n569 B.n568 585
R969 B.n567 B.n80 585
R970 B.n566 B.n565 585
R971 B.n564 B.n81 585
R972 B.n563 B.n562 585
R973 B.n561 B.n82 585
R974 B.n560 B.n559 585
R975 B.n558 B.n83 585
R976 B.n557 B.n556 585
R977 B.n555 B.n84 585
R978 B.n554 B.n553 585
R979 B.n552 B.n85 585
R980 B.n551 B.n550 585
R981 B.n549 B.n86 585
R982 B.n548 B.n547 585
R983 B.n546 B.n87 585
R984 B.n545 B.n544 585
R985 B.n543 B.n88 585
R986 B.n542 B.n541 585
R987 B.n540 B.n89 585
R988 B.n539 B.n538 585
R989 B.n537 B.n90 585
R990 B.n536 B.n535 585
R991 B.n534 B.n91 585
R992 B.n533 B.n532 585
R993 B.n531 B.n92 585
R994 B.n530 B.n529 585
R995 B.n528 B.n93 585
R996 B.n527 B.n526 585
R997 B.n525 B.n94 585
R998 B.n524 B.n523 585
R999 B.n522 B.n95 585
R1000 B.n521 B.n520 585
R1001 B.n519 B.n96 585
R1002 B.n518 B.n517 585
R1003 B.n516 B.n97 585
R1004 B.n515 B.n514 585
R1005 B.n513 B.n98 585
R1006 B.n512 B.n511 585
R1007 B.n510 B.n99 585
R1008 B.n509 B.n508 585
R1009 B.n507 B.n100 585
R1010 B.n506 B.n505 585
R1011 B.n504 B.n101 585
R1012 B.n503 B.n502 585
R1013 B.n501 B.n102 585
R1014 B.n500 B.n499 585
R1015 B.n498 B.n103 585
R1016 B.n497 B.n496 585
R1017 B.n495 B.n104 585
R1018 B.n494 B.n493 585
R1019 B.n492 B.n105 585
R1020 B.n491 B.n490 585
R1021 B.n489 B.n106 585
R1022 B.n488 B.n487 585
R1023 B.n486 B.n107 585
R1024 B.n485 B.n484 585
R1025 B.n483 B.n108 585
R1026 B.n482 B.n481 585
R1027 B.n480 B.n109 585
R1028 B.n479 B.n478 585
R1029 B.n477 B.n110 585
R1030 B.n476 B.n475 585
R1031 B.n474 B.n111 585
R1032 B.n473 B.n472 585
R1033 B.n471 B.n112 585
R1034 B.n470 B.n469 585
R1035 B.n468 B.n113 585
R1036 B.n467 B.n466 585
R1037 B.n465 B.n114 585
R1038 B.n464 B.n463 585
R1039 B.n462 B.n115 585
R1040 B.n461 B.n460 585
R1041 B.n459 B.n116 585
R1042 B.n458 B.n457 585
R1043 B.n456 B.n117 585
R1044 B.n455 B.n454 585
R1045 B.n453 B.n118 585
R1046 B.n452 B.n451 585
R1047 B.n450 B.n119 585
R1048 B.n449 B.n448 585
R1049 B.n447 B.n120 585
R1050 B.n446 B.n445 585
R1051 B.n444 B.n121 585
R1052 B.n443 B.n442 585
R1053 B.n441 B.n122 585
R1054 B.n440 B.n439 585
R1055 B.n438 B.n123 585
R1056 B.n437 B.n436 585
R1057 B.n435 B.n124 585
R1058 B.n434 B.n433 585
R1059 B.n432 B.n125 585
R1060 B.n431 B.n430 585
R1061 B.n429 B.n126 585
R1062 B.n428 B.n427 585
R1063 B.n426 B.n127 585
R1064 B.n425 B.n424 585
R1065 B.n423 B.n128 585
R1066 B.n422 B.n421 585
R1067 B.n420 B.n129 585
R1068 B.n419 B.n418 585
R1069 B.n417 B.n130 585
R1070 B.n416 B.n415 585
R1071 B.n414 B.n131 585
R1072 B.n413 B.n412 585
R1073 B.n411 B.n132 585
R1074 B.n410 B.n409 585
R1075 B.n408 B.n133 585
R1076 B.n407 B.n406 585
R1077 B.n405 B.n134 585
R1078 B.n296 B.n295 585
R1079 B.n297 B.n174 585
R1080 B.n299 B.n298 585
R1081 B.n300 B.n173 585
R1082 B.n302 B.n301 585
R1083 B.n303 B.n172 585
R1084 B.n305 B.n304 585
R1085 B.n306 B.n171 585
R1086 B.n308 B.n307 585
R1087 B.n309 B.n170 585
R1088 B.n311 B.n310 585
R1089 B.n312 B.n169 585
R1090 B.n314 B.n313 585
R1091 B.n315 B.n168 585
R1092 B.n317 B.n316 585
R1093 B.n318 B.n167 585
R1094 B.n320 B.n319 585
R1095 B.n321 B.n166 585
R1096 B.n323 B.n322 585
R1097 B.n324 B.n165 585
R1098 B.n326 B.n325 585
R1099 B.n327 B.n164 585
R1100 B.n329 B.n328 585
R1101 B.n330 B.n163 585
R1102 B.n332 B.n331 585
R1103 B.n333 B.n162 585
R1104 B.n335 B.n334 585
R1105 B.n336 B.n161 585
R1106 B.n338 B.n337 585
R1107 B.n339 B.n160 585
R1108 B.n341 B.n340 585
R1109 B.n343 B.n157 585
R1110 B.n345 B.n344 585
R1111 B.n346 B.n156 585
R1112 B.n348 B.n347 585
R1113 B.n349 B.n155 585
R1114 B.n351 B.n350 585
R1115 B.n352 B.n154 585
R1116 B.n354 B.n353 585
R1117 B.n355 B.n153 585
R1118 B.n357 B.n356 585
R1119 B.n359 B.n358 585
R1120 B.n360 B.n149 585
R1121 B.n362 B.n361 585
R1122 B.n363 B.n148 585
R1123 B.n365 B.n364 585
R1124 B.n366 B.n147 585
R1125 B.n368 B.n367 585
R1126 B.n369 B.n146 585
R1127 B.n371 B.n370 585
R1128 B.n372 B.n145 585
R1129 B.n374 B.n373 585
R1130 B.n375 B.n144 585
R1131 B.n377 B.n376 585
R1132 B.n378 B.n143 585
R1133 B.n380 B.n379 585
R1134 B.n381 B.n142 585
R1135 B.n383 B.n382 585
R1136 B.n384 B.n141 585
R1137 B.n386 B.n385 585
R1138 B.n387 B.n140 585
R1139 B.n389 B.n388 585
R1140 B.n390 B.n139 585
R1141 B.n392 B.n391 585
R1142 B.n393 B.n138 585
R1143 B.n395 B.n394 585
R1144 B.n396 B.n137 585
R1145 B.n398 B.n397 585
R1146 B.n399 B.n136 585
R1147 B.n401 B.n400 585
R1148 B.n402 B.n135 585
R1149 B.n404 B.n403 585
R1150 B.n294 B.n175 585
R1151 B.n293 B.n292 585
R1152 B.n291 B.n176 585
R1153 B.n290 B.n289 585
R1154 B.n288 B.n177 585
R1155 B.n287 B.n286 585
R1156 B.n285 B.n178 585
R1157 B.n284 B.n283 585
R1158 B.n282 B.n179 585
R1159 B.n281 B.n280 585
R1160 B.n279 B.n180 585
R1161 B.n278 B.n277 585
R1162 B.n276 B.n181 585
R1163 B.n275 B.n274 585
R1164 B.n273 B.n182 585
R1165 B.n272 B.n271 585
R1166 B.n270 B.n183 585
R1167 B.n269 B.n268 585
R1168 B.n267 B.n184 585
R1169 B.n266 B.n265 585
R1170 B.n264 B.n185 585
R1171 B.n263 B.n262 585
R1172 B.n261 B.n186 585
R1173 B.n260 B.n259 585
R1174 B.n258 B.n187 585
R1175 B.n257 B.n256 585
R1176 B.n255 B.n188 585
R1177 B.n254 B.n253 585
R1178 B.n252 B.n189 585
R1179 B.n251 B.n250 585
R1180 B.n249 B.n190 585
R1181 B.n248 B.n247 585
R1182 B.n246 B.n191 585
R1183 B.n245 B.n244 585
R1184 B.n243 B.n192 585
R1185 B.n242 B.n241 585
R1186 B.n240 B.n193 585
R1187 B.n239 B.n238 585
R1188 B.n237 B.n194 585
R1189 B.n236 B.n235 585
R1190 B.n234 B.n195 585
R1191 B.n233 B.n232 585
R1192 B.n231 B.n196 585
R1193 B.n230 B.n229 585
R1194 B.n228 B.n197 585
R1195 B.n227 B.n226 585
R1196 B.n225 B.n198 585
R1197 B.n224 B.n223 585
R1198 B.n222 B.n199 585
R1199 B.n221 B.n220 585
R1200 B.n219 B.n200 585
R1201 B.n218 B.n217 585
R1202 B.n216 B.n201 585
R1203 B.n215 B.n214 585
R1204 B.n213 B.n202 585
R1205 B.n212 B.n211 585
R1206 B.n210 B.n203 585
R1207 B.n209 B.n208 585
R1208 B.n207 B.n204 585
R1209 B.n206 B.n205 585
R1210 B.n2 B.n0 585
R1211 B.n789 B.n1 585
R1212 B.n788 B.n787 585
R1213 B.n786 B.n3 585
R1214 B.n785 B.n784 585
R1215 B.n783 B.n4 585
R1216 B.n782 B.n781 585
R1217 B.n780 B.n5 585
R1218 B.n779 B.n778 585
R1219 B.n777 B.n6 585
R1220 B.n776 B.n775 585
R1221 B.n774 B.n7 585
R1222 B.n773 B.n772 585
R1223 B.n771 B.n8 585
R1224 B.n770 B.n769 585
R1225 B.n768 B.n9 585
R1226 B.n767 B.n766 585
R1227 B.n765 B.n10 585
R1228 B.n764 B.n763 585
R1229 B.n762 B.n11 585
R1230 B.n761 B.n760 585
R1231 B.n759 B.n12 585
R1232 B.n758 B.n757 585
R1233 B.n756 B.n13 585
R1234 B.n755 B.n754 585
R1235 B.n753 B.n14 585
R1236 B.n752 B.n751 585
R1237 B.n750 B.n15 585
R1238 B.n749 B.n748 585
R1239 B.n747 B.n16 585
R1240 B.n746 B.n745 585
R1241 B.n744 B.n17 585
R1242 B.n743 B.n742 585
R1243 B.n741 B.n18 585
R1244 B.n740 B.n739 585
R1245 B.n738 B.n19 585
R1246 B.n737 B.n736 585
R1247 B.n735 B.n20 585
R1248 B.n734 B.n733 585
R1249 B.n732 B.n21 585
R1250 B.n731 B.n730 585
R1251 B.n729 B.n22 585
R1252 B.n728 B.n727 585
R1253 B.n726 B.n23 585
R1254 B.n725 B.n724 585
R1255 B.n723 B.n24 585
R1256 B.n722 B.n721 585
R1257 B.n720 B.n25 585
R1258 B.n719 B.n718 585
R1259 B.n717 B.n26 585
R1260 B.n716 B.n715 585
R1261 B.n714 B.n27 585
R1262 B.n713 B.n712 585
R1263 B.n711 B.n28 585
R1264 B.n710 B.n709 585
R1265 B.n708 B.n29 585
R1266 B.n707 B.n706 585
R1267 B.n705 B.n30 585
R1268 B.n704 B.n703 585
R1269 B.n702 B.n31 585
R1270 B.n701 B.n700 585
R1271 B.n699 B.n32 585
R1272 B.n791 B.n790 585
R1273 B.n296 B.n175 540.549
R1274 B.n699 B.n698 540.549
R1275 B.n405 B.n404 540.549
R1276 B.n590 B.n73 540.549
R1277 B.n150 B.t8 371.168
R1278 B.n56 B.t1 371.168
R1279 B.n158 B.t11 371.168
R1280 B.n48 B.t4 371.168
R1281 B.n151 B.t7 312.986
R1282 B.n57 B.t2 312.986
R1283 B.n159 B.t10 312.986
R1284 B.n49 B.t5 312.986
R1285 B.n150 B.t6 285.144
R1286 B.n158 B.t9 285.144
R1287 B.n48 B.t3 285.144
R1288 B.n56 B.t0 285.144
R1289 B.n292 B.n175 163.367
R1290 B.n292 B.n291 163.367
R1291 B.n291 B.n290 163.367
R1292 B.n290 B.n177 163.367
R1293 B.n286 B.n177 163.367
R1294 B.n286 B.n285 163.367
R1295 B.n285 B.n284 163.367
R1296 B.n284 B.n179 163.367
R1297 B.n280 B.n179 163.367
R1298 B.n280 B.n279 163.367
R1299 B.n279 B.n278 163.367
R1300 B.n278 B.n181 163.367
R1301 B.n274 B.n181 163.367
R1302 B.n274 B.n273 163.367
R1303 B.n273 B.n272 163.367
R1304 B.n272 B.n183 163.367
R1305 B.n268 B.n183 163.367
R1306 B.n268 B.n267 163.367
R1307 B.n267 B.n266 163.367
R1308 B.n266 B.n185 163.367
R1309 B.n262 B.n185 163.367
R1310 B.n262 B.n261 163.367
R1311 B.n261 B.n260 163.367
R1312 B.n260 B.n187 163.367
R1313 B.n256 B.n187 163.367
R1314 B.n256 B.n255 163.367
R1315 B.n255 B.n254 163.367
R1316 B.n254 B.n189 163.367
R1317 B.n250 B.n189 163.367
R1318 B.n250 B.n249 163.367
R1319 B.n249 B.n248 163.367
R1320 B.n248 B.n191 163.367
R1321 B.n244 B.n191 163.367
R1322 B.n244 B.n243 163.367
R1323 B.n243 B.n242 163.367
R1324 B.n242 B.n193 163.367
R1325 B.n238 B.n193 163.367
R1326 B.n238 B.n237 163.367
R1327 B.n237 B.n236 163.367
R1328 B.n236 B.n195 163.367
R1329 B.n232 B.n195 163.367
R1330 B.n232 B.n231 163.367
R1331 B.n231 B.n230 163.367
R1332 B.n230 B.n197 163.367
R1333 B.n226 B.n197 163.367
R1334 B.n226 B.n225 163.367
R1335 B.n225 B.n224 163.367
R1336 B.n224 B.n199 163.367
R1337 B.n220 B.n199 163.367
R1338 B.n220 B.n219 163.367
R1339 B.n219 B.n218 163.367
R1340 B.n218 B.n201 163.367
R1341 B.n214 B.n201 163.367
R1342 B.n214 B.n213 163.367
R1343 B.n213 B.n212 163.367
R1344 B.n212 B.n203 163.367
R1345 B.n208 B.n203 163.367
R1346 B.n208 B.n207 163.367
R1347 B.n207 B.n206 163.367
R1348 B.n206 B.n2 163.367
R1349 B.n790 B.n2 163.367
R1350 B.n790 B.n789 163.367
R1351 B.n789 B.n788 163.367
R1352 B.n788 B.n3 163.367
R1353 B.n784 B.n3 163.367
R1354 B.n784 B.n783 163.367
R1355 B.n783 B.n782 163.367
R1356 B.n782 B.n5 163.367
R1357 B.n778 B.n5 163.367
R1358 B.n778 B.n777 163.367
R1359 B.n777 B.n776 163.367
R1360 B.n776 B.n7 163.367
R1361 B.n772 B.n7 163.367
R1362 B.n772 B.n771 163.367
R1363 B.n771 B.n770 163.367
R1364 B.n770 B.n9 163.367
R1365 B.n766 B.n9 163.367
R1366 B.n766 B.n765 163.367
R1367 B.n765 B.n764 163.367
R1368 B.n764 B.n11 163.367
R1369 B.n760 B.n11 163.367
R1370 B.n760 B.n759 163.367
R1371 B.n759 B.n758 163.367
R1372 B.n758 B.n13 163.367
R1373 B.n754 B.n13 163.367
R1374 B.n754 B.n753 163.367
R1375 B.n753 B.n752 163.367
R1376 B.n752 B.n15 163.367
R1377 B.n748 B.n15 163.367
R1378 B.n748 B.n747 163.367
R1379 B.n747 B.n746 163.367
R1380 B.n746 B.n17 163.367
R1381 B.n742 B.n17 163.367
R1382 B.n742 B.n741 163.367
R1383 B.n741 B.n740 163.367
R1384 B.n740 B.n19 163.367
R1385 B.n736 B.n19 163.367
R1386 B.n736 B.n735 163.367
R1387 B.n735 B.n734 163.367
R1388 B.n734 B.n21 163.367
R1389 B.n730 B.n21 163.367
R1390 B.n730 B.n729 163.367
R1391 B.n729 B.n728 163.367
R1392 B.n728 B.n23 163.367
R1393 B.n724 B.n23 163.367
R1394 B.n724 B.n723 163.367
R1395 B.n723 B.n722 163.367
R1396 B.n722 B.n25 163.367
R1397 B.n718 B.n25 163.367
R1398 B.n718 B.n717 163.367
R1399 B.n717 B.n716 163.367
R1400 B.n716 B.n27 163.367
R1401 B.n712 B.n27 163.367
R1402 B.n712 B.n711 163.367
R1403 B.n711 B.n710 163.367
R1404 B.n710 B.n29 163.367
R1405 B.n706 B.n29 163.367
R1406 B.n706 B.n705 163.367
R1407 B.n705 B.n704 163.367
R1408 B.n704 B.n31 163.367
R1409 B.n700 B.n31 163.367
R1410 B.n700 B.n699 163.367
R1411 B.n297 B.n296 163.367
R1412 B.n298 B.n297 163.367
R1413 B.n298 B.n173 163.367
R1414 B.n302 B.n173 163.367
R1415 B.n303 B.n302 163.367
R1416 B.n304 B.n303 163.367
R1417 B.n304 B.n171 163.367
R1418 B.n308 B.n171 163.367
R1419 B.n309 B.n308 163.367
R1420 B.n310 B.n309 163.367
R1421 B.n310 B.n169 163.367
R1422 B.n314 B.n169 163.367
R1423 B.n315 B.n314 163.367
R1424 B.n316 B.n315 163.367
R1425 B.n316 B.n167 163.367
R1426 B.n320 B.n167 163.367
R1427 B.n321 B.n320 163.367
R1428 B.n322 B.n321 163.367
R1429 B.n322 B.n165 163.367
R1430 B.n326 B.n165 163.367
R1431 B.n327 B.n326 163.367
R1432 B.n328 B.n327 163.367
R1433 B.n328 B.n163 163.367
R1434 B.n332 B.n163 163.367
R1435 B.n333 B.n332 163.367
R1436 B.n334 B.n333 163.367
R1437 B.n334 B.n161 163.367
R1438 B.n338 B.n161 163.367
R1439 B.n339 B.n338 163.367
R1440 B.n340 B.n339 163.367
R1441 B.n340 B.n157 163.367
R1442 B.n345 B.n157 163.367
R1443 B.n346 B.n345 163.367
R1444 B.n347 B.n346 163.367
R1445 B.n347 B.n155 163.367
R1446 B.n351 B.n155 163.367
R1447 B.n352 B.n351 163.367
R1448 B.n353 B.n352 163.367
R1449 B.n353 B.n153 163.367
R1450 B.n357 B.n153 163.367
R1451 B.n358 B.n357 163.367
R1452 B.n358 B.n149 163.367
R1453 B.n362 B.n149 163.367
R1454 B.n363 B.n362 163.367
R1455 B.n364 B.n363 163.367
R1456 B.n364 B.n147 163.367
R1457 B.n368 B.n147 163.367
R1458 B.n369 B.n368 163.367
R1459 B.n370 B.n369 163.367
R1460 B.n370 B.n145 163.367
R1461 B.n374 B.n145 163.367
R1462 B.n375 B.n374 163.367
R1463 B.n376 B.n375 163.367
R1464 B.n376 B.n143 163.367
R1465 B.n380 B.n143 163.367
R1466 B.n381 B.n380 163.367
R1467 B.n382 B.n381 163.367
R1468 B.n382 B.n141 163.367
R1469 B.n386 B.n141 163.367
R1470 B.n387 B.n386 163.367
R1471 B.n388 B.n387 163.367
R1472 B.n388 B.n139 163.367
R1473 B.n392 B.n139 163.367
R1474 B.n393 B.n392 163.367
R1475 B.n394 B.n393 163.367
R1476 B.n394 B.n137 163.367
R1477 B.n398 B.n137 163.367
R1478 B.n399 B.n398 163.367
R1479 B.n400 B.n399 163.367
R1480 B.n400 B.n135 163.367
R1481 B.n404 B.n135 163.367
R1482 B.n406 B.n405 163.367
R1483 B.n406 B.n133 163.367
R1484 B.n410 B.n133 163.367
R1485 B.n411 B.n410 163.367
R1486 B.n412 B.n411 163.367
R1487 B.n412 B.n131 163.367
R1488 B.n416 B.n131 163.367
R1489 B.n417 B.n416 163.367
R1490 B.n418 B.n417 163.367
R1491 B.n418 B.n129 163.367
R1492 B.n422 B.n129 163.367
R1493 B.n423 B.n422 163.367
R1494 B.n424 B.n423 163.367
R1495 B.n424 B.n127 163.367
R1496 B.n428 B.n127 163.367
R1497 B.n429 B.n428 163.367
R1498 B.n430 B.n429 163.367
R1499 B.n430 B.n125 163.367
R1500 B.n434 B.n125 163.367
R1501 B.n435 B.n434 163.367
R1502 B.n436 B.n435 163.367
R1503 B.n436 B.n123 163.367
R1504 B.n440 B.n123 163.367
R1505 B.n441 B.n440 163.367
R1506 B.n442 B.n441 163.367
R1507 B.n442 B.n121 163.367
R1508 B.n446 B.n121 163.367
R1509 B.n447 B.n446 163.367
R1510 B.n448 B.n447 163.367
R1511 B.n448 B.n119 163.367
R1512 B.n452 B.n119 163.367
R1513 B.n453 B.n452 163.367
R1514 B.n454 B.n453 163.367
R1515 B.n454 B.n117 163.367
R1516 B.n458 B.n117 163.367
R1517 B.n459 B.n458 163.367
R1518 B.n460 B.n459 163.367
R1519 B.n460 B.n115 163.367
R1520 B.n464 B.n115 163.367
R1521 B.n465 B.n464 163.367
R1522 B.n466 B.n465 163.367
R1523 B.n466 B.n113 163.367
R1524 B.n470 B.n113 163.367
R1525 B.n471 B.n470 163.367
R1526 B.n472 B.n471 163.367
R1527 B.n472 B.n111 163.367
R1528 B.n476 B.n111 163.367
R1529 B.n477 B.n476 163.367
R1530 B.n478 B.n477 163.367
R1531 B.n478 B.n109 163.367
R1532 B.n482 B.n109 163.367
R1533 B.n483 B.n482 163.367
R1534 B.n484 B.n483 163.367
R1535 B.n484 B.n107 163.367
R1536 B.n488 B.n107 163.367
R1537 B.n489 B.n488 163.367
R1538 B.n490 B.n489 163.367
R1539 B.n490 B.n105 163.367
R1540 B.n494 B.n105 163.367
R1541 B.n495 B.n494 163.367
R1542 B.n496 B.n495 163.367
R1543 B.n496 B.n103 163.367
R1544 B.n500 B.n103 163.367
R1545 B.n501 B.n500 163.367
R1546 B.n502 B.n501 163.367
R1547 B.n502 B.n101 163.367
R1548 B.n506 B.n101 163.367
R1549 B.n507 B.n506 163.367
R1550 B.n508 B.n507 163.367
R1551 B.n508 B.n99 163.367
R1552 B.n512 B.n99 163.367
R1553 B.n513 B.n512 163.367
R1554 B.n514 B.n513 163.367
R1555 B.n514 B.n97 163.367
R1556 B.n518 B.n97 163.367
R1557 B.n519 B.n518 163.367
R1558 B.n520 B.n519 163.367
R1559 B.n520 B.n95 163.367
R1560 B.n524 B.n95 163.367
R1561 B.n525 B.n524 163.367
R1562 B.n526 B.n525 163.367
R1563 B.n526 B.n93 163.367
R1564 B.n530 B.n93 163.367
R1565 B.n531 B.n530 163.367
R1566 B.n532 B.n531 163.367
R1567 B.n532 B.n91 163.367
R1568 B.n536 B.n91 163.367
R1569 B.n537 B.n536 163.367
R1570 B.n538 B.n537 163.367
R1571 B.n538 B.n89 163.367
R1572 B.n542 B.n89 163.367
R1573 B.n543 B.n542 163.367
R1574 B.n544 B.n543 163.367
R1575 B.n544 B.n87 163.367
R1576 B.n548 B.n87 163.367
R1577 B.n549 B.n548 163.367
R1578 B.n550 B.n549 163.367
R1579 B.n550 B.n85 163.367
R1580 B.n554 B.n85 163.367
R1581 B.n555 B.n554 163.367
R1582 B.n556 B.n555 163.367
R1583 B.n556 B.n83 163.367
R1584 B.n560 B.n83 163.367
R1585 B.n561 B.n560 163.367
R1586 B.n562 B.n561 163.367
R1587 B.n562 B.n81 163.367
R1588 B.n566 B.n81 163.367
R1589 B.n567 B.n566 163.367
R1590 B.n568 B.n567 163.367
R1591 B.n568 B.n79 163.367
R1592 B.n572 B.n79 163.367
R1593 B.n573 B.n572 163.367
R1594 B.n574 B.n573 163.367
R1595 B.n574 B.n77 163.367
R1596 B.n578 B.n77 163.367
R1597 B.n579 B.n578 163.367
R1598 B.n580 B.n579 163.367
R1599 B.n580 B.n75 163.367
R1600 B.n584 B.n75 163.367
R1601 B.n585 B.n584 163.367
R1602 B.n586 B.n585 163.367
R1603 B.n586 B.n73 163.367
R1604 B.n698 B.n33 163.367
R1605 B.n694 B.n33 163.367
R1606 B.n694 B.n693 163.367
R1607 B.n693 B.n692 163.367
R1608 B.n692 B.n35 163.367
R1609 B.n688 B.n35 163.367
R1610 B.n688 B.n687 163.367
R1611 B.n687 B.n686 163.367
R1612 B.n686 B.n37 163.367
R1613 B.n682 B.n37 163.367
R1614 B.n682 B.n681 163.367
R1615 B.n681 B.n680 163.367
R1616 B.n680 B.n39 163.367
R1617 B.n676 B.n39 163.367
R1618 B.n676 B.n675 163.367
R1619 B.n675 B.n674 163.367
R1620 B.n674 B.n41 163.367
R1621 B.n670 B.n41 163.367
R1622 B.n670 B.n669 163.367
R1623 B.n669 B.n668 163.367
R1624 B.n668 B.n43 163.367
R1625 B.n664 B.n43 163.367
R1626 B.n664 B.n663 163.367
R1627 B.n663 B.n662 163.367
R1628 B.n662 B.n45 163.367
R1629 B.n658 B.n45 163.367
R1630 B.n658 B.n657 163.367
R1631 B.n657 B.n656 163.367
R1632 B.n656 B.n47 163.367
R1633 B.n652 B.n47 163.367
R1634 B.n652 B.n651 163.367
R1635 B.n651 B.n51 163.367
R1636 B.n647 B.n51 163.367
R1637 B.n647 B.n646 163.367
R1638 B.n646 B.n645 163.367
R1639 B.n645 B.n53 163.367
R1640 B.n641 B.n53 163.367
R1641 B.n641 B.n640 163.367
R1642 B.n640 B.n639 163.367
R1643 B.n639 B.n55 163.367
R1644 B.n634 B.n55 163.367
R1645 B.n634 B.n633 163.367
R1646 B.n633 B.n632 163.367
R1647 B.n632 B.n59 163.367
R1648 B.n628 B.n59 163.367
R1649 B.n628 B.n627 163.367
R1650 B.n627 B.n626 163.367
R1651 B.n626 B.n61 163.367
R1652 B.n622 B.n61 163.367
R1653 B.n622 B.n621 163.367
R1654 B.n621 B.n620 163.367
R1655 B.n620 B.n63 163.367
R1656 B.n616 B.n63 163.367
R1657 B.n616 B.n615 163.367
R1658 B.n615 B.n614 163.367
R1659 B.n614 B.n65 163.367
R1660 B.n610 B.n65 163.367
R1661 B.n610 B.n609 163.367
R1662 B.n609 B.n608 163.367
R1663 B.n608 B.n67 163.367
R1664 B.n604 B.n67 163.367
R1665 B.n604 B.n603 163.367
R1666 B.n603 B.n602 163.367
R1667 B.n602 B.n69 163.367
R1668 B.n598 B.n69 163.367
R1669 B.n598 B.n597 163.367
R1670 B.n597 B.n596 163.367
R1671 B.n596 B.n71 163.367
R1672 B.n592 B.n71 163.367
R1673 B.n592 B.n591 163.367
R1674 B.n591 B.n590 163.367
R1675 B.n152 B.n151 59.5399
R1676 B.n342 B.n159 59.5399
R1677 B.n50 B.n49 59.5399
R1678 B.n636 B.n57 59.5399
R1679 B.n151 B.n150 58.1823
R1680 B.n159 B.n158 58.1823
R1681 B.n49 B.n48 58.1823
R1682 B.n57 B.n56 58.1823
R1683 B.n697 B.n32 35.1225
R1684 B.n589 B.n588 35.1225
R1685 B.n403 B.n134 35.1225
R1686 B.n295 B.n294 35.1225
R1687 B B.n791 18.0485
R1688 B.n697 B.n696 10.6151
R1689 B.n696 B.n695 10.6151
R1690 B.n695 B.n34 10.6151
R1691 B.n691 B.n34 10.6151
R1692 B.n691 B.n690 10.6151
R1693 B.n690 B.n689 10.6151
R1694 B.n689 B.n36 10.6151
R1695 B.n685 B.n36 10.6151
R1696 B.n685 B.n684 10.6151
R1697 B.n684 B.n683 10.6151
R1698 B.n683 B.n38 10.6151
R1699 B.n679 B.n38 10.6151
R1700 B.n679 B.n678 10.6151
R1701 B.n678 B.n677 10.6151
R1702 B.n677 B.n40 10.6151
R1703 B.n673 B.n40 10.6151
R1704 B.n673 B.n672 10.6151
R1705 B.n672 B.n671 10.6151
R1706 B.n671 B.n42 10.6151
R1707 B.n667 B.n42 10.6151
R1708 B.n667 B.n666 10.6151
R1709 B.n666 B.n665 10.6151
R1710 B.n665 B.n44 10.6151
R1711 B.n661 B.n44 10.6151
R1712 B.n661 B.n660 10.6151
R1713 B.n660 B.n659 10.6151
R1714 B.n659 B.n46 10.6151
R1715 B.n655 B.n46 10.6151
R1716 B.n655 B.n654 10.6151
R1717 B.n654 B.n653 10.6151
R1718 B.n650 B.n649 10.6151
R1719 B.n649 B.n648 10.6151
R1720 B.n648 B.n52 10.6151
R1721 B.n644 B.n52 10.6151
R1722 B.n644 B.n643 10.6151
R1723 B.n643 B.n642 10.6151
R1724 B.n642 B.n54 10.6151
R1725 B.n638 B.n54 10.6151
R1726 B.n638 B.n637 10.6151
R1727 B.n635 B.n58 10.6151
R1728 B.n631 B.n58 10.6151
R1729 B.n631 B.n630 10.6151
R1730 B.n630 B.n629 10.6151
R1731 B.n629 B.n60 10.6151
R1732 B.n625 B.n60 10.6151
R1733 B.n625 B.n624 10.6151
R1734 B.n624 B.n623 10.6151
R1735 B.n623 B.n62 10.6151
R1736 B.n619 B.n62 10.6151
R1737 B.n619 B.n618 10.6151
R1738 B.n618 B.n617 10.6151
R1739 B.n617 B.n64 10.6151
R1740 B.n613 B.n64 10.6151
R1741 B.n613 B.n612 10.6151
R1742 B.n612 B.n611 10.6151
R1743 B.n611 B.n66 10.6151
R1744 B.n607 B.n66 10.6151
R1745 B.n607 B.n606 10.6151
R1746 B.n606 B.n605 10.6151
R1747 B.n605 B.n68 10.6151
R1748 B.n601 B.n68 10.6151
R1749 B.n601 B.n600 10.6151
R1750 B.n600 B.n599 10.6151
R1751 B.n599 B.n70 10.6151
R1752 B.n595 B.n70 10.6151
R1753 B.n595 B.n594 10.6151
R1754 B.n594 B.n593 10.6151
R1755 B.n593 B.n72 10.6151
R1756 B.n589 B.n72 10.6151
R1757 B.n407 B.n134 10.6151
R1758 B.n408 B.n407 10.6151
R1759 B.n409 B.n408 10.6151
R1760 B.n409 B.n132 10.6151
R1761 B.n413 B.n132 10.6151
R1762 B.n414 B.n413 10.6151
R1763 B.n415 B.n414 10.6151
R1764 B.n415 B.n130 10.6151
R1765 B.n419 B.n130 10.6151
R1766 B.n420 B.n419 10.6151
R1767 B.n421 B.n420 10.6151
R1768 B.n421 B.n128 10.6151
R1769 B.n425 B.n128 10.6151
R1770 B.n426 B.n425 10.6151
R1771 B.n427 B.n426 10.6151
R1772 B.n427 B.n126 10.6151
R1773 B.n431 B.n126 10.6151
R1774 B.n432 B.n431 10.6151
R1775 B.n433 B.n432 10.6151
R1776 B.n433 B.n124 10.6151
R1777 B.n437 B.n124 10.6151
R1778 B.n438 B.n437 10.6151
R1779 B.n439 B.n438 10.6151
R1780 B.n439 B.n122 10.6151
R1781 B.n443 B.n122 10.6151
R1782 B.n444 B.n443 10.6151
R1783 B.n445 B.n444 10.6151
R1784 B.n445 B.n120 10.6151
R1785 B.n449 B.n120 10.6151
R1786 B.n450 B.n449 10.6151
R1787 B.n451 B.n450 10.6151
R1788 B.n451 B.n118 10.6151
R1789 B.n455 B.n118 10.6151
R1790 B.n456 B.n455 10.6151
R1791 B.n457 B.n456 10.6151
R1792 B.n457 B.n116 10.6151
R1793 B.n461 B.n116 10.6151
R1794 B.n462 B.n461 10.6151
R1795 B.n463 B.n462 10.6151
R1796 B.n463 B.n114 10.6151
R1797 B.n467 B.n114 10.6151
R1798 B.n468 B.n467 10.6151
R1799 B.n469 B.n468 10.6151
R1800 B.n469 B.n112 10.6151
R1801 B.n473 B.n112 10.6151
R1802 B.n474 B.n473 10.6151
R1803 B.n475 B.n474 10.6151
R1804 B.n475 B.n110 10.6151
R1805 B.n479 B.n110 10.6151
R1806 B.n480 B.n479 10.6151
R1807 B.n481 B.n480 10.6151
R1808 B.n481 B.n108 10.6151
R1809 B.n485 B.n108 10.6151
R1810 B.n486 B.n485 10.6151
R1811 B.n487 B.n486 10.6151
R1812 B.n487 B.n106 10.6151
R1813 B.n491 B.n106 10.6151
R1814 B.n492 B.n491 10.6151
R1815 B.n493 B.n492 10.6151
R1816 B.n493 B.n104 10.6151
R1817 B.n497 B.n104 10.6151
R1818 B.n498 B.n497 10.6151
R1819 B.n499 B.n498 10.6151
R1820 B.n499 B.n102 10.6151
R1821 B.n503 B.n102 10.6151
R1822 B.n504 B.n503 10.6151
R1823 B.n505 B.n504 10.6151
R1824 B.n505 B.n100 10.6151
R1825 B.n509 B.n100 10.6151
R1826 B.n510 B.n509 10.6151
R1827 B.n511 B.n510 10.6151
R1828 B.n511 B.n98 10.6151
R1829 B.n515 B.n98 10.6151
R1830 B.n516 B.n515 10.6151
R1831 B.n517 B.n516 10.6151
R1832 B.n517 B.n96 10.6151
R1833 B.n521 B.n96 10.6151
R1834 B.n522 B.n521 10.6151
R1835 B.n523 B.n522 10.6151
R1836 B.n523 B.n94 10.6151
R1837 B.n527 B.n94 10.6151
R1838 B.n528 B.n527 10.6151
R1839 B.n529 B.n528 10.6151
R1840 B.n529 B.n92 10.6151
R1841 B.n533 B.n92 10.6151
R1842 B.n534 B.n533 10.6151
R1843 B.n535 B.n534 10.6151
R1844 B.n535 B.n90 10.6151
R1845 B.n539 B.n90 10.6151
R1846 B.n540 B.n539 10.6151
R1847 B.n541 B.n540 10.6151
R1848 B.n541 B.n88 10.6151
R1849 B.n545 B.n88 10.6151
R1850 B.n546 B.n545 10.6151
R1851 B.n547 B.n546 10.6151
R1852 B.n547 B.n86 10.6151
R1853 B.n551 B.n86 10.6151
R1854 B.n552 B.n551 10.6151
R1855 B.n553 B.n552 10.6151
R1856 B.n553 B.n84 10.6151
R1857 B.n557 B.n84 10.6151
R1858 B.n558 B.n557 10.6151
R1859 B.n559 B.n558 10.6151
R1860 B.n559 B.n82 10.6151
R1861 B.n563 B.n82 10.6151
R1862 B.n564 B.n563 10.6151
R1863 B.n565 B.n564 10.6151
R1864 B.n565 B.n80 10.6151
R1865 B.n569 B.n80 10.6151
R1866 B.n570 B.n569 10.6151
R1867 B.n571 B.n570 10.6151
R1868 B.n571 B.n78 10.6151
R1869 B.n575 B.n78 10.6151
R1870 B.n576 B.n575 10.6151
R1871 B.n577 B.n576 10.6151
R1872 B.n577 B.n76 10.6151
R1873 B.n581 B.n76 10.6151
R1874 B.n582 B.n581 10.6151
R1875 B.n583 B.n582 10.6151
R1876 B.n583 B.n74 10.6151
R1877 B.n587 B.n74 10.6151
R1878 B.n588 B.n587 10.6151
R1879 B.n295 B.n174 10.6151
R1880 B.n299 B.n174 10.6151
R1881 B.n300 B.n299 10.6151
R1882 B.n301 B.n300 10.6151
R1883 B.n301 B.n172 10.6151
R1884 B.n305 B.n172 10.6151
R1885 B.n306 B.n305 10.6151
R1886 B.n307 B.n306 10.6151
R1887 B.n307 B.n170 10.6151
R1888 B.n311 B.n170 10.6151
R1889 B.n312 B.n311 10.6151
R1890 B.n313 B.n312 10.6151
R1891 B.n313 B.n168 10.6151
R1892 B.n317 B.n168 10.6151
R1893 B.n318 B.n317 10.6151
R1894 B.n319 B.n318 10.6151
R1895 B.n319 B.n166 10.6151
R1896 B.n323 B.n166 10.6151
R1897 B.n324 B.n323 10.6151
R1898 B.n325 B.n324 10.6151
R1899 B.n325 B.n164 10.6151
R1900 B.n329 B.n164 10.6151
R1901 B.n330 B.n329 10.6151
R1902 B.n331 B.n330 10.6151
R1903 B.n331 B.n162 10.6151
R1904 B.n335 B.n162 10.6151
R1905 B.n336 B.n335 10.6151
R1906 B.n337 B.n336 10.6151
R1907 B.n337 B.n160 10.6151
R1908 B.n341 B.n160 10.6151
R1909 B.n344 B.n343 10.6151
R1910 B.n344 B.n156 10.6151
R1911 B.n348 B.n156 10.6151
R1912 B.n349 B.n348 10.6151
R1913 B.n350 B.n349 10.6151
R1914 B.n350 B.n154 10.6151
R1915 B.n354 B.n154 10.6151
R1916 B.n355 B.n354 10.6151
R1917 B.n356 B.n355 10.6151
R1918 B.n360 B.n359 10.6151
R1919 B.n361 B.n360 10.6151
R1920 B.n361 B.n148 10.6151
R1921 B.n365 B.n148 10.6151
R1922 B.n366 B.n365 10.6151
R1923 B.n367 B.n366 10.6151
R1924 B.n367 B.n146 10.6151
R1925 B.n371 B.n146 10.6151
R1926 B.n372 B.n371 10.6151
R1927 B.n373 B.n372 10.6151
R1928 B.n373 B.n144 10.6151
R1929 B.n377 B.n144 10.6151
R1930 B.n378 B.n377 10.6151
R1931 B.n379 B.n378 10.6151
R1932 B.n379 B.n142 10.6151
R1933 B.n383 B.n142 10.6151
R1934 B.n384 B.n383 10.6151
R1935 B.n385 B.n384 10.6151
R1936 B.n385 B.n140 10.6151
R1937 B.n389 B.n140 10.6151
R1938 B.n390 B.n389 10.6151
R1939 B.n391 B.n390 10.6151
R1940 B.n391 B.n138 10.6151
R1941 B.n395 B.n138 10.6151
R1942 B.n396 B.n395 10.6151
R1943 B.n397 B.n396 10.6151
R1944 B.n397 B.n136 10.6151
R1945 B.n401 B.n136 10.6151
R1946 B.n402 B.n401 10.6151
R1947 B.n403 B.n402 10.6151
R1948 B.n294 B.n293 10.6151
R1949 B.n293 B.n176 10.6151
R1950 B.n289 B.n176 10.6151
R1951 B.n289 B.n288 10.6151
R1952 B.n288 B.n287 10.6151
R1953 B.n287 B.n178 10.6151
R1954 B.n283 B.n178 10.6151
R1955 B.n283 B.n282 10.6151
R1956 B.n282 B.n281 10.6151
R1957 B.n281 B.n180 10.6151
R1958 B.n277 B.n180 10.6151
R1959 B.n277 B.n276 10.6151
R1960 B.n276 B.n275 10.6151
R1961 B.n275 B.n182 10.6151
R1962 B.n271 B.n182 10.6151
R1963 B.n271 B.n270 10.6151
R1964 B.n270 B.n269 10.6151
R1965 B.n269 B.n184 10.6151
R1966 B.n265 B.n184 10.6151
R1967 B.n265 B.n264 10.6151
R1968 B.n264 B.n263 10.6151
R1969 B.n263 B.n186 10.6151
R1970 B.n259 B.n186 10.6151
R1971 B.n259 B.n258 10.6151
R1972 B.n258 B.n257 10.6151
R1973 B.n257 B.n188 10.6151
R1974 B.n253 B.n188 10.6151
R1975 B.n253 B.n252 10.6151
R1976 B.n252 B.n251 10.6151
R1977 B.n251 B.n190 10.6151
R1978 B.n247 B.n190 10.6151
R1979 B.n247 B.n246 10.6151
R1980 B.n246 B.n245 10.6151
R1981 B.n245 B.n192 10.6151
R1982 B.n241 B.n192 10.6151
R1983 B.n241 B.n240 10.6151
R1984 B.n240 B.n239 10.6151
R1985 B.n239 B.n194 10.6151
R1986 B.n235 B.n194 10.6151
R1987 B.n235 B.n234 10.6151
R1988 B.n234 B.n233 10.6151
R1989 B.n233 B.n196 10.6151
R1990 B.n229 B.n196 10.6151
R1991 B.n229 B.n228 10.6151
R1992 B.n228 B.n227 10.6151
R1993 B.n227 B.n198 10.6151
R1994 B.n223 B.n198 10.6151
R1995 B.n223 B.n222 10.6151
R1996 B.n222 B.n221 10.6151
R1997 B.n221 B.n200 10.6151
R1998 B.n217 B.n200 10.6151
R1999 B.n217 B.n216 10.6151
R2000 B.n216 B.n215 10.6151
R2001 B.n215 B.n202 10.6151
R2002 B.n211 B.n202 10.6151
R2003 B.n211 B.n210 10.6151
R2004 B.n210 B.n209 10.6151
R2005 B.n209 B.n204 10.6151
R2006 B.n205 B.n204 10.6151
R2007 B.n205 B.n0 10.6151
R2008 B.n787 B.n1 10.6151
R2009 B.n787 B.n786 10.6151
R2010 B.n786 B.n785 10.6151
R2011 B.n785 B.n4 10.6151
R2012 B.n781 B.n4 10.6151
R2013 B.n781 B.n780 10.6151
R2014 B.n780 B.n779 10.6151
R2015 B.n779 B.n6 10.6151
R2016 B.n775 B.n6 10.6151
R2017 B.n775 B.n774 10.6151
R2018 B.n774 B.n773 10.6151
R2019 B.n773 B.n8 10.6151
R2020 B.n769 B.n8 10.6151
R2021 B.n769 B.n768 10.6151
R2022 B.n768 B.n767 10.6151
R2023 B.n767 B.n10 10.6151
R2024 B.n763 B.n10 10.6151
R2025 B.n763 B.n762 10.6151
R2026 B.n762 B.n761 10.6151
R2027 B.n761 B.n12 10.6151
R2028 B.n757 B.n12 10.6151
R2029 B.n757 B.n756 10.6151
R2030 B.n756 B.n755 10.6151
R2031 B.n755 B.n14 10.6151
R2032 B.n751 B.n14 10.6151
R2033 B.n751 B.n750 10.6151
R2034 B.n750 B.n749 10.6151
R2035 B.n749 B.n16 10.6151
R2036 B.n745 B.n16 10.6151
R2037 B.n745 B.n744 10.6151
R2038 B.n744 B.n743 10.6151
R2039 B.n743 B.n18 10.6151
R2040 B.n739 B.n18 10.6151
R2041 B.n739 B.n738 10.6151
R2042 B.n738 B.n737 10.6151
R2043 B.n737 B.n20 10.6151
R2044 B.n733 B.n20 10.6151
R2045 B.n733 B.n732 10.6151
R2046 B.n732 B.n731 10.6151
R2047 B.n731 B.n22 10.6151
R2048 B.n727 B.n22 10.6151
R2049 B.n727 B.n726 10.6151
R2050 B.n726 B.n725 10.6151
R2051 B.n725 B.n24 10.6151
R2052 B.n721 B.n24 10.6151
R2053 B.n721 B.n720 10.6151
R2054 B.n720 B.n719 10.6151
R2055 B.n719 B.n26 10.6151
R2056 B.n715 B.n26 10.6151
R2057 B.n715 B.n714 10.6151
R2058 B.n714 B.n713 10.6151
R2059 B.n713 B.n28 10.6151
R2060 B.n709 B.n28 10.6151
R2061 B.n709 B.n708 10.6151
R2062 B.n708 B.n707 10.6151
R2063 B.n707 B.n30 10.6151
R2064 B.n703 B.n30 10.6151
R2065 B.n703 B.n702 10.6151
R2066 B.n702 B.n701 10.6151
R2067 B.n701 B.n32 10.6151
R2068 B.n653 B.n50 9.36635
R2069 B.n636 B.n635 9.36635
R2070 B.n342 B.n341 9.36635
R2071 B.n359 B.n152 9.36635
R2072 B.n791 B.n0 2.81026
R2073 B.n791 B.n1 2.81026
R2074 B.n650 B.n50 1.24928
R2075 B.n637 B.n636 1.24928
R2076 B.n343 B.n342 1.24928
R2077 B.n356 B.n152 1.24928
C0 VTAIL VP 8.62165f
C1 w_n4570_n2674# VDD1 2.56777f
C2 VP w_n4570_n2674# 10.3478f
C3 VTAIL VDD2 8.881701f
C4 B VN 1.26039f
C5 VDD2 w_n4570_n2674# 2.71495f
C6 B VDD1 2.23309f
C7 VDD1 VN 0.153079f
C8 VTAIL w_n4570_n2674# 2.72374f
C9 VP B 2.26165f
C10 VP VN 7.86351f
C11 VDD2 B 2.35373f
C12 VP VDD1 8.21732f
C13 VDD2 VN 7.78185f
C14 VTAIL B 2.97883f
C15 VTAIL VN 8.60742f
C16 VDD2 VDD1 2.21649f
C17 B w_n4570_n2674# 9.69193f
C18 VDD2 VP 0.591796f
C19 w_n4570_n2674# VN 9.75263f
C20 VTAIL VDD1 8.82942f
C21 VDD2 VSUBS 2.140133f
C22 VDD1 VSUBS 1.902505f
C23 VTAIL VSUBS 1.202159f
C24 VN VSUBS 7.73959f
C25 VP VSUBS 4.214962f
C26 B VSUBS 5.163039f
C27 w_n4570_n2674# VSUBS 0.151413p
C28 B.n0 VSUBS 0.006651f
C29 B.n1 VSUBS 0.006651f
C30 B.n2 VSUBS 0.010518f
C31 B.n3 VSUBS 0.010518f
C32 B.n4 VSUBS 0.010518f
C33 B.n5 VSUBS 0.010518f
C34 B.n6 VSUBS 0.010518f
C35 B.n7 VSUBS 0.010518f
C36 B.n8 VSUBS 0.010518f
C37 B.n9 VSUBS 0.010518f
C38 B.n10 VSUBS 0.010518f
C39 B.n11 VSUBS 0.010518f
C40 B.n12 VSUBS 0.010518f
C41 B.n13 VSUBS 0.010518f
C42 B.n14 VSUBS 0.010518f
C43 B.n15 VSUBS 0.010518f
C44 B.n16 VSUBS 0.010518f
C45 B.n17 VSUBS 0.010518f
C46 B.n18 VSUBS 0.010518f
C47 B.n19 VSUBS 0.010518f
C48 B.n20 VSUBS 0.010518f
C49 B.n21 VSUBS 0.010518f
C50 B.n22 VSUBS 0.010518f
C51 B.n23 VSUBS 0.010518f
C52 B.n24 VSUBS 0.010518f
C53 B.n25 VSUBS 0.010518f
C54 B.n26 VSUBS 0.010518f
C55 B.n27 VSUBS 0.010518f
C56 B.n28 VSUBS 0.010518f
C57 B.n29 VSUBS 0.010518f
C58 B.n30 VSUBS 0.010518f
C59 B.n31 VSUBS 0.010518f
C60 B.n32 VSUBS 0.025423f
C61 B.n33 VSUBS 0.010518f
C62 B.n34 VSUBS 0.010518f
C63 B.n35 VSUBS 0.010518f
C64 B.n36 VSUBS 0.010518f
C65 B.n37 VSUBS 0.010518f
C66 B.n38 VSUBS 0.010518f
C67 B.n39 VSUBS 0.010518f
C68 B.n40 VSUBS 0.010518f
C69 B.n41 VSUBS 0.010518f
C70 B.n42 VSUBS 0.010518f
C71 B.n43 VSUBS 0.010518f
C72 B.n44 VSUBS 0.010518f
C73 B.n45 VSUBS 0.010518f
C74 B.n46 VSUBS 0.010518f
C75 B.n47 VSUBS 0.010518f
C76 B.t5 VSUBS 0.205752f
C77 B.t4 VSUBS 0.250688f
C78 B.t3 VSUBS 1.59256f
C79 B.n48 VSUBS 0.413202f
C80 B.n49 VSUBS 0.301664f
C81 B.n50 VSUBS 0.02437f
C82 B.n51 VSUBS 0.010518f
C83 B.n52 VSUBS 0.010518f
C84 B.n53 VSUBS 0.010518f
C85 B.n54 VSUBS 0.010518f
C86 B.n55 VSUBS 0.010518f
C87 B.t2 VSUBS 0.205756f
C88 B.t1 VSUBS 0.250691f
C89 B.t0 VSUBS 1.59256f
C90 B.n56 VSUBS 0.413199f
C91 B.n57 VSUBS 0.301661f
C92 B.n58 VSUBS 0.010518f
C93 B.n59 VSUBS 0.010518f
C94 B.n60 VSUBS 0.010518f
C95 B.n61 VSUBS 0.010518f
C96 B.n62 VSUBS 0.010518f
C97 B.n63 VSUBS 0.010518f
C98 B.n64 VSUBS 0.010518f
C99 B.n65 VSUBS 0.010518f
C100 B.n66 VSUBS 0.010518f
C101 B.n67 VSUBS 0.010518f
C102 B.n68 VSUBS 0.010518f
C103 B.n69 VSUBS 0.010518f
C104 B.n70 VSUBS 0.010518f
C105 B.n71 VSUBS 0.010518f
C106 B.n72 VSUBS 0.010518f
C107 B.n73 VSUBS 0.025423f
C108 B.n74 VSUBS 0.010518f
C109 B.n75 VSUBS 0.010518f
C110 B.n76 VSUBS 0.010518f
C111 B.n77 VSUBS 0.010518f
C112 B.n78 VSUBS 0.010518f
C113 B.n79 VSUBS 0.010518f
C114 B.n80 VSUBS 0.010518f
C115 B.n81 VSUBS 0.010518f
C116 B.n82 VSUBS 0.010518f
C117 B.n83 VSUBS 0.010518f
C118 B.n84 VSUBS 0.010518f
C119 B.n85 VSUBS 0.010518f
C120 B.n86 VSUBS 0.010518f
C121 B.n87 VSUBS 0.010518f
C122 B.n88 VSUBS 0.010518f
C123 B.n89 VSUBS 0.010518f
C124 B.n90 VSUBS 0.010518f
C125 B.n91 VSUBS 0.010518f
C126 B.n92 VSUBS 0.010518f
C127 B.n93 VSUBS 0.010518f
C128 B.n94 VSUBS 0.010518f
C129 B.n95 VSUBS 0.010518f
C130 B.n96 VSUBS 0.010518f
C131 B.n97 VSUBS 0.010518f
C132 B.n98 VSUBS 0.010518f
C133 B.n99 VSUBS 0.010518f
C134 B.n100 VSUBS 0.010518f
C135 B.n101 VSUBS 0.010518f
C136 B.n102 VSUBS 0.010518f
C137 B.n103 VSUBS 0.010518f
C138 B.n104 VSUBS 0.010518f
C139 B.n105 VSUBS 0.010518f
C140 B.n106 VSUBS 0.010518f
C141 B.n107 VSUBS 0.010518f
C142 B.n108 VSUBS 0.010518f
C143 B.n109 VSUBS 0.010518f
C144 B.n110 VSUBS 0.010518f
C145 B.n111 VSUBS 0.010518f
C146 B.n112 VSUBS 0.010518f
C147 B.n113 VSUBS 0.010518f
C148 B.n114 VSUBS 0.010518f
C149 B.n115 VSUBS 0.010518f
C150 B.n116 VSUBS 0.010518f
C151 B.n117 VSUBS 0.010518f
C152 B.n118 VSUBS 0.010518f
C153 B.n119 VSUBS 0.010518f
C154 B.n120 VSUBS 0.010518f
C155 B.n121 VSUBS 0.010518f
C156 B.n122 VSUBS 0.010518f
C157 B.n123 VSUBS 0.010518f
C158 B.n124 VSUBS 0.010518f
C159 B.n125 VSUBS 0.010518f
C160 B.n126 VSUBS 0.010518f
C161 B.n127 VSUBS 0.010518f
C162 B.n128 VSUBS 0.010518f
C163 B.n129 VSUBS 0.010518f
C164 B.n130 VSUBS 0.010518f
C165 B.n131 VSUBS 0.010518f
C166 B.n132 VSUBS 0.010518f
C167 B.n133 VSUBS 0.010518f
C168 B.n134 VSUBS 0.025423f
C169 B.n135 VSUBS 0.010518f
C170 B.n136 VSUBS 0.010518f
C171 B.n137 VSUBS 0.010518f
C172 B.n138 VSUBS 0.010518f
C173 B.n139 VSUBS 0.010518f
C174 B.n140 VSUBS 0.010518f
C175 B.n141 VSUBS 0.010518f
C176 B.n142 VSUBS 0.010518f
C177 B.n143 VSUBS 0.010518f
C178 B.n144 VSUBS 0.010518f
C179 B.n145 VSUBS 0.010518f
C180 B.n146 VSUBS 0.010518f
C181 B.n147 VSUBS 0.010518f
C182 B.n148 VSUBS 0.010518f
C183 B.n149 VSUBS 0.010518f
C184 B.t7 VSUBS 0.205756f
C185 B.t8 VSUBS 0.250691f
C186 B.t6 VSUBS 1.59256f
C187 B.n150 VSUBS 0.413199f
C188 B.n151 VSUBS 0.301661f
C189 B.n152 VSUBS 0.02437f
C190 B.n153 VSUBS 0.010518f
C191 B.n154 VSUBS 0.010518f
C192 B.n155 VSUBS 0.010518f
C193 B.n156 VSUBS 0.010518f
C194 B.n157 VSUBS 0.010518f
C195 B.t10 VSUBS 0.205752f
C196 B.t11 VSUBS 0.250688f
C197 B.t9 VSUBS 1.59256f
C198 B.n158 VSUBS 0.413202f
C199 B.n159 VSUBS 0.301664f
C200 B.n160 VSUBS 0.010518f
C201 B.n161 VSUBS 0.010518f
C202 B.n162 VSUBS 0.010518f
C203 B.n163 VSUBS 0.010518f
C204 B.n164 VSUBS 0.010518f
C205 B.n165 VSUBS 0.010518f
C206 B.n166 VSUBS 0.010518f
C207 B.n167 VSUBS 0.010518f
C208 B.n168 VSUBS 0.010518f
C209 B.n169 VSUBS 0.010518f
C210 B.n170 VSUBS 0.010518f
C211 B.n171 VSUBS 0.010518f
C212 B.n172 VSUBS 0.010518f
C213 B.n173 VSUBS 0.010518f
C214 B.n174 VSUBS 0.010518f
C215 B.n175 VSUBS 0.025423f
C216 B.n176 VSUBS 0.010518f
C217 B.n177 VSUBS 0.010518f
C218 B.n178 VSUBS 0.010518f
C219 B.n179 VSUBS 0.010518f
C220 B.n180 VSUBS 0.010518f
C221 B.n181 VSUBS 0.010518f
C222 B.n182 VSUBS 0.010518f
C223 B.n183 VSUBS 0.010518f
C224 B.n184 VSUBS 0.010518f
C225 B.n185 VSUBS 0.010518f
C226 B.n186 VSUBS 0.010518f
C227 B.n187 VSUBS 0.010518f
C228 B.n188 VSUBS 0.010518f
C229 B.n189 VSUBS 0.010518f
C230 B.n190 VSUBS 0.010518f
C231 B.n191 VSUBS 0.010518f
C232 B.n192 VSUBS 0.010518f
C233 B.n193 VSUBS 0.010518f
C234 B.n194 VSUBS 0.010518f
C235 B.n195 VSUBS 0.010518f
C236 B.n196 VSUBS 0.010518f
C237 B.n197 VSUBS 0.010518f
C238 B.n198 VSUBS 0.010518f
C239 B.n199 VSUBS 0.010518f
C240 B.n200 VSUBS 0.010518f
C241 B.n201 VSUBS 0.010518f
C242 B.n202 VSUBS 0.010518f
C243 B.n203 VSUBS 0.010518f
C244 B.n204 VSUBS 0.010518f
C245 B.n205 VSUBS 0.010518f
C246 B.n206 VSUBS 0.010518f
C247 B.n207 VSUBS 0.010518f
C248 B.n208 VSUBS 0.010518f
C249 B.n209 VSUBS 0.010518f
C250 B.n210 VSUBS 0.010518f
C251 B.n211 VSUBS 0.010518f
C252 B.n212 VSUBS 0.010518f
C253 B.n213 VSUBS 0.010518f
C254 B.n214 VSUBS 0.010518f
C255 B.n215 VSUBS 0.010518f
C256 B.n216 VSUBS 0.010518f
C257 B.n217 VSUBS 0.010518f
C258 B.n218 VSUBS 0.010518f
C259 B.n219 VSUBS 0.010518f
C260 B.n220 VSUBS 0.010518f
C261 B.n221 VSUBS 0.010518f
C262 B.n222 VSUBS 0.010518f
C263 B.n223 VSUBS 0.010518f
C264 B.n224 VSUBS 0.010518f
C265 B.n225 VSUBS 0.010518f
C266 B.n226 VSUBS 0.010518f
C267 B.n227 VSUBS 0.010518f
C268 B.n228 VSUBS 0.010518f
C269 B.n229 VSUBS 0.010518f
C270 B.n230 VSUBS 0.010518f
C271 B.n231 VSUBS 0.010518f
C272 B.n232 VSUBS 0.010518f
C273 B.n233 VSUBS 0.010518f
C274 B.n234 VSUBS 0.010518f
C275 B.n235 VSUBS 0.010518f
C276 B.n236 VSUBS 0.010518f
C277 B.n237 VSUBS 0.010518f
C278 B.n238 VSUBS 0.010518f
C279 B.n239 VSUBS 0.010518f
C280 B.n240 VSUBS 0.010518f
C281 B.n241 VSUBS 0.010518f
C282 B.n242 VSUBS 0.010518f
C283 B.n243 VSUBS 0.010518f
C284 B.n244 VSUBS 0.010518f
C285 B.n245 VSUBS 0.010518f
C286 B.n246 VSUBS 0.010518f
C287 B.n247 VSUBS 0.010518f
C288 B.n248 VSUBS 0.010518f
C289 B.n249 VSUBS 0.010518f
C290 B.n250 VSUBS 0.010518f
C291 B.n251 VSUBS 0.010518f
C292 B.n252 VSUBS 0.010518f
C293 B.n253 VSUBS 0.010518f
C294 B.n254 VSUBS 0.010518f
C295 B.n255 VSUBS 0.010518f
C296 B.n256 VSUBS 0.010518f
C297 B.n257 VSUBS 0.010518f
C298 B.n258 VSUBS 0.010518f
C299 B.n259 VSUBS 0.010518f
C300 B.n260 VSUBS 0.010518f
C301 B.n261 VSUBS 0.010518f
C302 B.n262 VSUBS 0.010518f
C303 B.n263 VSUBS 0.010518f
C304 B.n264 VSUBS 0.010518f
C305 B.n265 VSUBS 0.010518f
C306 B.n266 VSUBS 0.010518f
C307 B.n267 VSUBS 0.010518f
C308 B.n268 VSUBS 0.010518f
C309 B.n269 VSUBS 0.010518f
C310 B.n270 VSUBS 0.010518f
C311 B.n271 VSUBS 0.010518f
C312 B.n272 VSUBS 0.010518f
C313 B.n273 VSUBS 0.010518f
C314 B.n274 VSUBS 0.010518f
C315 B.n275 VSUBS 0.010518f
C316 B.n276 VSUBS 0.010518f
C317 B.n277 VSUBS 0.010518f
C318 B.n278 VSUBS 0.010518f
C319 B.n279 VSUBS 0.010518f
C320 B.n280 VSUBS 0.010518f
C321 B.n281 VSUBS 0.010518f
C322 B.n282 VSUBS 0.010518f
C323 B.n283 VSUBS 0.010518f
C324 B.n284 VSUBS 0.010518f
C325 B.n285 VSUBS 0.010518f
C326 B.n286 VSUBS 0.010518f
C327 B.n287 VSUBS 0.010518f
C328 B.n288 VSUBS 0.010518f
C329 B.n289 VSUBS 0.010518f
C330 B.n290 VSUBS 0.010518f
C331 B.n291 VSUBS 0.010518f
C332 B.n292 VSUBS 0.010518f
C333 B.n293 VSUBS 0.010518f
C334 B.n294 VSUBS 0.025423f
C335 B.n295 VSUBS 0.02624f
C336 B.n296 VSUBS 0.02624f
C337 B.n297 VSUBS 0.010518f
C338 B.n298 VSUBS 0.010518f
C339 B.n299 VSUBS 0.010518f
C340 B.n300 VSUBS 0.010518f
C341 B.n301 VSUBS 0.010518f
C342 B.n302 VSUBS 0.010518f
C343 B.n303 VSUBS 0.010518f
C344 B.n304 VSUBS 0.010518f
C345 B.n305 VSUBS 0.010518f
C346 B.n306 VSUBS 0.010518f
C347 B.n307 VSUBS 0.010518f
C348 B.n308 VSUBS 0.010518f
C349 B.n309 VSUBS 0.010518f
C350 B.n310 VSUBS 0.010518f
C351 B.n311 VSUBS 0.010518f
C352 B.n312 VSUBS 0.010518f
C353 B.n313 VSUBS 0.010518f
C354 B.n314 VSUBS 0.010518f
C355 B.n315 VSUBS 0.010518f
C356 B.n316 VSUBS 0.010518f
C357 B.n317 VSUBS 0.010518f
C358 B.n318 VSUBS 0.010518f
C359 B.n319 VSUBS 0.010518f
C360 B.n320 VSUBS 0.010518f
C361 B.n321 VSUBS 0.010518f
C362 B.n322 VSUBS 0.010518f
C363 B.n323 VSUBS 0.010518f
C364 B.n324 VSUBS 0.010518f
C365 B.n325 VSUBS 0.010518f
C366 B.n326 VSUBS 0.010518f
C367 B.n327 VSUBS 0.010518f
C368 B.n328 VSUBS 0.010518f
C369 B.n329 VSUBS 0.010518f
C370 B.n330 VSUBS 0.010518f
C371 B.n331 VSUBS 0.010518f
C372 B.n332 VSUBS 0.010518f
C373 B.n333 VSUBS 0.010518f
C374 B.n334 VSUBS 0.010518f
C375 B.n335 VSUBS 0.010518f
C376 B.n336 VSUBS 0.010518f
C377 B.n337 VSUBS 0.010518f
C378 B.n338 VSUBS 0.010518f
C379 B.n339 VSUBS 0.010518f
C380 B.n340 VSUBS 0.010518f
C381 B.n341 VSUBS 0.0099f
C382 B.n342 VSUBS 0.02437f
C383 B.n343 VSUBS 0.005878f
C384 B.n344 VSUBS 0.010518f
C385 B.n345 VSUBS 0.010518f
C386 B.n346 VSUBS 0.010518f
C387 B.n347 VSUBS 0.010518f
C388 B.n348 VSUBS 0.010518f
C389 B.n349 VSUBS 0.010518f
C390 B.n350 VSUBS 0.010518f
C391 B.n351 VSUBS 0.010518f
C392 B.n352 VSUBS 0.010518f
C393 B.n353 VSUBS 0.010518f
C394 B.n354 VSUBS 0.010518f
C395 B.n355 VSUBS 0.010518f
C396 B.n356 VSUBS 0.005878f
C397 B.n357 VSUBS 0.010518f
C398 B.n358 VSUBS 0.010518f
C399 B.n359 VSUBS 0.0099f
C400 B.n360 VSUBS 0.010518f
C401 B.n361 VSUBS 0.010518f
C402 B.n362 VSUBS 0.010518f
C403 B.n363 VSUBS 0.010518f
C404 B.n364 VSUBS 0.010518f
C405 B.n365 VSUBS 0.010518f
C406 B.n366 VSUBS 0.010518f
C407 B.n367 VSUBS 0.010518f
C408 B.n368 VSUBS 0.010518f
C409 B.n369 VSUBS 0.010518f
C410 B.n370 VSUBS 0.010518f
C411 B.n371 VSUBS 0.010518f
C412 B.n372 VSUBS 0.010518f
C413 B.n373 VSUBS 0.010518f
C414 B.n374 VSUBS 0.010518f
C415 B.n375 VSUBS 0.010518f
C416 B.n376 VSUBS 0.010518f
C417 B.n377 VSUBS 0.010518f
C418 B.n378 VSUBS 0.010518f
C419 B.n379 VSUBS 0.010518f
C420 B.n380 VSUBS 0.010518f
C421 B.n381 VSUBS 0.010518f
C422 B.n382 VSUBS 0.010518f
C423 B.n383 VSUBS 0.010518f
C424 B.n384 VSUBS 0.010518f
C425 B.n385 VSUBS 0.010518f
C426 B.n386 VSUBS 0.010518f
C427 B.n387 VSUBS 0.010518f
C428 B.n388 VSUBS 0.010518f
C429 B.n389 VSUBS 0.010518f
C430 B.n390 VSUBS 0.010518f
C431 B.n391 VSUBS 0.010518f
C432 B.n392 VSUBS 0.010518f
C433 B.n393 VSUBS 0.010518f
C434 B.n394 VSUBS 0.010518f
C435 B.n395 VSUBS 0.010518f
C436 B.n396 VSUBS 0.010518f
C437 B.n397 VSUBS 0.010518f
C438 B.n398 VSUBS 0.010518f
C439 B.n399 VSUBS 0.010518f
C440 B.n400 VSUBS 0.010518f
C441 B.n401 VSUBS 0.010518f
C442 B.n402 VSUBS 0.010518f
C443 B.n403 VSUBS 0.02624f
C444 B.n404 VSUBS 0.02624f
C445 B.n405 VSUBS 0.025423f
C446 B.n406 VSUBS 0.010518f
C447 B.n407 VSUBS 0.010518f
C448 B.n408 VSUBS 0.010518f
C449 B.n409 VSUBS 0.010518f
C450 B.n410 VSUBS 0.010518f
C451 B.n411 VSUBS 0.010518f
C452 B.n412 VSUBS 0.010518f
C453 B.n413 VSUBS 0.010518f
C454 B.n414 VSUBS 0.010518f
C455 B.n415 VSUBS 0.010518f
C456 B.n416 VSUBS 0.010518f
C457 B.n417 VSUBS 0.010518f
C458 B.n418 VSUBS 0.010518f
C459 B.n419 VSUBS 0.010518f
C460 B.n420 VSUBS 0.010518f
C461 B.n421 VSUBS 0.010518f
C462 B.n422 VSUBS 0.010518f
C463 B.n423 VSUBS 0.010518f
C464 B.n424 VSUBS 0.010518f
C465 B.n425 VSUBS 0.010518f
C466 B.n426 VSUBS 0.010518f
C467 B.n427 VSUBS 0.010518f
C468 B.n428 VSUBS 0.010518f
C469 B.n429 VSUBS 0.010518f
C470 B.n430 VSUBS 0.010518f
C471 B.n431 VSUBS 0.010518f
C472 B.n432 VSUBS 0.010518f
C473 B.n433 VSUBS 0.010518f
C474 B.n434 VSUBS 0.010518f
C475 B.n435 VSUBS 0.010518f
C476 B.n436 VSUBS 0.010518f
C477 B.n437 VSUBS 0.010518f
C478 B.n438 VSUBS 0.010518f
C479 B.n439 VSUBS 0.010518f
C480 B.n440 VSUBS 0.010518f
C481 B.n441 VSUBS 0.010518f
C482 B.n442 VSUBS 0.010518f
C483 B.n443 VSUBS 0.010518f
C484 B.n444 VSUBS 0.010518f
C485 B.n445 VSUBS 0.010518f
C486 B.n446 VSUBS 0.010518f
C487 B.n447 VSUBS 0.010518f
C488 B.n448 VSUBS 0.010518f
C489 B.n449 VSUBS 0.010518f
C490 B.n450 VSUBS 0.010518f
C491 B.n451 VSUBS 0.010518f
C492 B.n452 VSUBS 0.010518f
C493 B.n453 VSUBS 0.010518f
C494 B.n454 VSUBS 0.010518f
C495 B.n455 VSUBS 0.010518f
C496 B.n456 VSUBS 0.010518f
C497 B.n457 VSUBS 0.010518f
C498 B.n458 VSUBS 0.010518f
C499 B.n459 VSUBS 0.010518f
C500 B.n460 VSUBS 0.010518f
C501 B.n461 VSUBS 0.010518f
C502 B.n462 VSUBS 0.010518f
C503 B.n463 VSUBS 0.010518f
C504 B.n464 VSUBS 0.010518f
C505 B.n465 VSUBS 0.010518f
C506 B.n466 VSUBS 0.010518f
C507 B.n467 VSUBS 0.010518f
C508 B.n468 VSUBS 0.010518f
C509 B.n469 VSUBS 0.010518f
C510 B.n470 VSUBS 0.010518f
C511 B.n471 VSUBS 0.010518f
C512 B.n472 VSUBS 0.010518f
C513 B.n473 VSUBS 0.010518f
C514 B.n474 VSUBS 0.010518f
C515 B.n475 VSUBS 0.010518f
C516 B.n476 VSUBS 0.010518f
C517 B.n477 VSUBS 0.010518f
C518 B.n478 VSUBS 0.010518f
C519 B.n479 VSUBS 0.010518f
C520 B.n480 VSUBS 0.010518f
C521 B.n481 VSUBS 0.010518f
C522 B.n482 VSUBS 0.010518f
C523 B.n483 VSUBS 0.010518f
C524 B.n484 VSUBS 0.010518f
C525 B.n485 VSUBS 0.010518f
C526 B.n486 VSUBS 0.010518f
C527 B.n487 VSUBS 0.010518f
C528 B.n488 VSUBS 0.010518f
C529 B.n489 VSUBS 0.010518f
C530 B.n490 VSUBS 0.010518f
C531 B.n491 VSUBS 0.010518f
C532 B.n492 VSUBS 0.010518f
C533 B.n493 VSUBS 0.010518f
C534 B.n494 VSUBS 0.010518f
C535 B.n495 VSUBS 0.010518f
C536 B.n496 VSUBS 0.010518f
C537 B.n497 VSUBS 0.010518f
C538 B.n498 VSUBS 0.010518f
C539 B.n499 VSUBS 0.010518f
C540 B.n500 VSUBS 0.010518f
C541 B.n501 VSUBS 0.010518f
C542 B.n502 VSUBS 0.010518f
C543 B.n503 VSUBS 0.010518f
C544 B.n504 VSUBS 0.010518f
C545 B.n505 VSUBS 0.010518f
C546 B.n506 VSUBS 0.010518f
C547 B.n507 VSUBS 0.010518f
C548 B.n508 VSUBS 0.010518f
C549 B.n509 VSUBS 0.010518f
C550 B.n510 VSUBS 0.010518f
C551 B.n511 VSUBS 0.010518f
C552 B.n512 VSUBS 0.010518f
C553 B.n513 VSUBS 0.010518f
C554 B.n514 VSUBS 0.010518f
C555 B.n515 VSUBS 0.010518f
C556 B.n516 VSUBS 0.010518f
C557 B.n517 VSUBS 0.010518f
C558 B.n518 VSUBS 0.010518f
C559 B.n519 VSUBS 0.010518f
C560 B.n520 VSUBS 0.010518f
C561 B.n521 VSUBS 0.010518f
C562 B.n522 VSUBS 0.010518f
C563 B.n523 VSUBS 0.010518f
C564 B.n524 VSUBS 0.010518f
C565 B.n525 VSUBS 0.010518f
C566 B.n526 VSUBS 0.010518f
C567 B.n527 VSUBS 0.010518f
C568 B.n528 VSUBS 0.010518f
C569 B.n529 VSUBS 0.010518f
C570 B.n530 VSUBS 0.010518f
C571 B.n531 VSUBS 0.010518f
C572 B.n532 VSUBS 0.010518f
C573 B.n533 VSUBS 0.010518f
C574 B.n534 VSUBS 0.010518f
C575 B.n535 VSUBS 0.010518f
C576 B.n536 VSUBS 0.010518f
C577 B.n537 VSUBS 0.010518f
C578 B.n538 VSUBS 0.010518f
C579 B.n539 VSUBS 0.010518f
C580 B.n540 VSUBS 0.010518f
C581 B.n541 VSUBS 0.010518f
C582 B.n542 VSUBS 0.010518f
C583 B.n543 VSUBS 0.010518f
C584 B.n544 VSUBS 0.010518f
C585 B.n545 VSUBS 0.010518f
C586 B.n546 VSUBS 0.010518f
C587 B.n547 VSUBS 0.010518f
C588 B.n548 VSUBS 0.010518f
C589 B.n549 VSUBS 0.010518f
C590 B.n550 VSUBS 0.010518f
C591 B.n551 VSUBS 0.010518f
C592 B.n552 VSUBS 0.010518f
C593 B.n553 VSUBS 0.010518f
C594 B.n554 VSUBS 0.010518f
C595 B.n555 VSUBS 0.010518f
C596 B.n556 VSUBS 0.010518f
C597 B.n557 VSUBS 0.010518f
C598 B.n558 VSUBS 0.010518f
C599 B.n559 VSUBS 0.010518f
C600 B.n560 VSUBS 0.010518f
C601 B.n561 VSUBS 0.010518f
C602 B.n562 VSUBS 0.010518f
C603 B.n563 VSUBS 0.010518f
C604 B.n564 VSUBS 0.010518f
C605 B.n565 VSUBS 0.010518f
C606 B.n566 VSUBS 0.010518f
C607 B.n567 VSUBS 0.010518f
C608 B.n568 VSUBS 0.010518f
C609 B.n569 VSUBS 0.010518f
C610 B.n570 VSUBS 0.010518f
C611 B.n571 VSUBS 0.010518f
C612 B.n572 VSUBS 0.010518f
C613 B.n573 VSUBS 0.010518f
C614 B.n574 VSUBS 0.010518f
C615 B.n575 VSUBS 0.010518f
C616 B.n576 VSUBS 0.010518f
C617 B.n577 VSUBS 0.010518f
C618 B.n578 VSUBS 0.010518f
C619 B.n579 VSUBS 0.010518f
C620 B.n580 VSUBS 0.010518f
C621 B.n581 VSUBS 0.010518f
C622 B.n582 VSUBS 0.010518f
C623 B.n583 VSUBS 0.010518f
C624 B.n584 VSUBS 0.010518f
C625 B.n585 VSUBS 0.010518f
C626 B.n586 VSUBS 0.010518f
C627 B.n587 VSUBS 0.010518f
C628 B.n588 VSUBS 0.026579f
C629 B.n589 VSUBS 0.025085f
C630 B.n590 VSUBS 0.02624f
C631 B.n591 VSUBS 0.010518f
C632 B.n592 VSUBS 0.010518f
C633 B.n593 VSUBS 0.010518f
C634 B.n594 VSUBS 0.010518f
C635 B.n595 VSUBS 0.010518f
C636 B.n596 VSUBS 0.010518f
C637 B.n597 VSUBS 0.010518f
C638 B.n598 VSUBS 0.010518f
C639 B.n599 VSUBS 0.010518f
C640 B.n600 VSUBS 0.010518f
C641 B.n601 VSUBS 0.010518f
C642 B.n602 VSUBS 0.010518f
C643 B.n603 VSUBS 0.010518f
C644 B.n604 VSUBS 0.010518f
C645 B.n605 VSUBS 0.010518f
C646 B.n606 VSUBS 0.010518f
C647 B.n607 VSUBS 0.010518f
C648 B.n608 VSUBS 0.010518f
C649 B.n609 VSUBS 0.010518f
C650 B.n610 VSUBS 0.010518f
C651 B.n611 VSUBS 0.010518f
C652 B.n612 VSUBS 0.010518f
C653 B.n613 VSUBS 0.010518f
C654 B.n614 VSUBS 0.010518f
C655 B.n615 VSUBS 0.010518f
C656 B.n616 VSUBS 0.010518f
C657 B.n617 VSUBS 0.010518f
C658 B.n618 VSUBS 0.010518f
C659 B.n619 VSUBS 0.010518f
C660 B.n620 VSUBS 0.010518f
C661 B.n621 VSUBS 0.010518f
C662 B.n622 VSUBS 0.010518f
C663 B.n623 VSUBS 0.010518f
C664 B.n624 VSUBS 0.010518f
C665 B.n625 VSUBS 0.010518f
C666 B.n626 VSUBS 0.010518f
C667 B.n627 VSUBS 0.010518f
C668 B.n628 VSUBS 0.010518f
C669 B.n629 VSUBS 0.010518f
C670 B.n630 VSUBS 0.010518f
C671 B.n631 VSUBS 0.010518f
C672 B.n632 VSUBS 0.010518f
C673 B.n633 VSUBS 0.010518f
C674 B.n634 VSUBS 0.010518f
C675 B.n635 VSUBS 0.0099f
C676 B.n636 VSUBS 0.02437f
C677 B.n637 VSUBS 0.005878f
C678 B.n638 VSUBS 0.010518f
C679 B.n639 VSUBS 0.010518f
C680 B.n640 VSUBS 0.010518f
C681 B.n641 VSUBS 0.010518f
C682 B.n642 VSUBS 0.010518f
C683 B.n643 VSUBS 0.010518f
C684 B.n644 VSUBS 0.010518f
C685 B.n645 VSUBS 0.010518f
C686 B.n646 VSUBS 0.010518f
C687 B.n647 VSUBS 0.010518f
C688 B.n648 VSUBS 0.010518f
C689 B.n649 VSUBS 0.010518f
C690 B.n650 VSUBS 0.005878f
C691 B.n651 VSUBS 0.010518f
C692 B.n652 VSUBS 0.010518f
C693 B.n653 VSUBS 0.0099f
C694 B.n654 VSUBS 0.010518f
C695 B.n655 VSUBS 0.010518f
C696 B.n656 VSUBS 0.010518f
C697 B.n657 VSUBS 0.010518f
C698 B.n658 VSUBS 0.010518f
C699 B.n659 VSUBS 0.010518f
C700 B.n660 VSUBS 0.010518f
C701 B.n661 VSUBS 0.010518f
C702 B.n662 VSUBS 0.010518f
C703 B.n663 VSUBS 0.010518f
C704 B.n664 VSUBS 0.010518f
C705 B.n665 VSUBS 0.010518f
C706 B.n666 VSUBS 0.010518f
C707 B.n667 VSUBS 0.010518f
C708 B.n668 VSUBS 0.010518f
C709 B.n669 VSUBS 0.010518f
C710 B.n670 VSUBS 0.010518f
C711 B.n671 VSUBS 0.010518f
C712 B.n672 VSUBS 0.010518f
C713 B.n673 VSUBS 0.010518f
C714 B.n674 VSUBS 0.010518f
C715 B.n675 VSUBS 0.010518f
C716 B.n676 VSUBS 0.010518f
C717 B.n677 VSUBS 0.010518f
C718 B.n678 VSUBS 0.010518f
C719 B.n679 VSUBS 0.010518f
C720 B.n680 VSUBS 0.010518f
C721 B.n681 VSUBS 0.010518f
C722 B.n682 VSUBS 0.010518f
C723 B.n683 VSUBS 0.010518f
C724 B.n684 VSUBS 0.010518f
C725 B.n685 VSUBS 0.010518f
C726 B.n686 VSUBS 0.010518f
C727 B.n687 VSUBS 0.010518f
C728 B.n688 VSUBS 0.010518f
C729 B.n689 VSUBS 0.010518f
C730 B.n690 VSUBS 0.010518f
C731 B.n691 VSUBS 0.010518f
C732 B.n692 VSUBS 0.010518f
C733 B.n693 VSUBS 0.010518f
C734 B.n694 VSUBS 0.010518f
C735 B.n695 VSUBS 0.010518f
C736 B.n696 VSUBS 0.010518f
C737 B.n697 VSUBS 0.02624f
C738 B.n698 VSUBS 0.02624f
C739 B.n699 VSUBS 0.025423f
C740 B.n700 VSUBS 0.010518f
C741 B.n701 VSUBS 0.010518f
C742 B.n702 VSUBS 0.010518f
C743 B.n703 VSUBS 0.010518f
C744 B.n704 VSUBS 0.010518f
C745 B.n705 VSUBS 0.010518f
C746 B.n706 VSUBS 0.010518f
C747 B.n707 VSUBS 0.010518f
C748 B.n708 VSUBS 0.010518f
C749 B.n709 VSUBS 0.010518f
C750 B.n710 VSUBS 0.010518f
C751 B.n711 VSUBS 0.010518f
C752 B.n712 VSUBS 0.010518f
C753 B.n713 VSUBS 0.010518f
C754 B.n714 VSUBS 0.010518f
C755 B.n715 VSUBS 0.010518f
C756 B.n716 VSUBS 0.010518f
C757 B.n717 VSUBS 0.010518f
C758 B.n718 VSUBS 0.010518f
C759 B.n719 VSUBS 0.010518f
C760 B.n720 VSUBS 0.010518f
C761 B.n721 VSUBS 0.010518f
C762 B.n722 VSUBS 0.010518f
C763 B.n723 VSUBS 0.010518f
C764 B.n724 VSUBS 0.010518f
C765 B.n725 VSUBS 0.010518f
C766 B.n726 VSUBS 0.010518f
C767 B.n727 VSUBS 0.010518f
C768 B.n728 VSUBS 0.010518f
C769 B.n729 VSUBS 0.010518f
C770 B.n730 VSUBS 0.010518f
C771 B.n731 VSUBS 0.010518f
C772 B.n732 VSUBS 0.010518f
C773 B.n733 VSUBS 0.010518f
C774 B.n734 VSUBS 0.010518f
C775 B.n735 VSUBS 0.010518f
C776 B.n736 VSUBS 0.010518f
C777 B.n737 VSUBS 0.010518f
C778 B.n738 VSUBS 0.010518f
C779 B.n739 VSUBS 0.010518f
C780 B.n740 VSUBS 0.010518f
C781 B.n741 VSUBS 0.010518f
C782 B.n742 VSUBS 0.010518f
C783 B.n743 VSUBS 0.010518f
C784 B.n744 VSUBS 0.010518f
C785 B.n745 VSUBS 0.010518f
C786 B.n746 VSUBS 0.010518f
C787 B.n747 VSUBS 0.010518f
C788 B.n748 VSUBS 0.010518f
C789 B.n749 VSUBS 0.010518f
C790 B.n750 VSUBS 0.010518f
C791 B.n751 VSUBS 0.010518f
C792 B.n752 VSUBS 0.010518f
C793 B.n753 VSUBS 0.010518f
C794 B.n754 VSUBS 0.010518f
C795 B.n755 VSUBS 0.010518f
C796 B.n756 VSUBS 0.010518f
C797 B.n757 VSUBS 0.010518f
C798 B.n758 VSUBS 0.010518f
C799 B.n759 VSUBS 0.010518f
C800 B.n760 VSUBS 0.010518f
C801 B.n761 VSUBS 0.010518f
C802 B.n762 VSUBS 0.010518f
C803 B.n763 VSUBS 0.010518f
C804 B.n764 VSUBS 0.010518f
C805 B.n765 VSUBS 0.010518f
C806 B.n766 VSUBS 0.010518f
C807 B.n767 VSUBS 0.010518f
C808 B.n768 VSUBS 0.010518f
C809 B.n769 VSUBS 0.010518f
C810 B.n770 VSUBS 0.010518f
C811 B.n771 VSUBS 0.010518f
C812 B.n772 VSUBS 0.010518f
C813 B.n773 VSUBS 0.010518f
C814 B.n774 VSUBS 0.010518f
C815 B.n775 VSUBS 0.010518f
C816 B.n776 VSUBS 0.010518f
C817 B.n777 VSUBS 0.010518f
C818 B.n778 VSUBS 0.010518f
C819 B.n779 VSUBS 0.010518f
C820 B.n780 VSUBS 0.010518f
C821 B.n781 VSUBS 0.010518f
C822 B.n782 VSUBS 0.010518f
C823 B.n783 VSUBS 0.010518f
C824 B.n784 VSUBS 0.010518f
C825 B.n785 VSUBS 0.010518f
C826 B.n786 VSUBS 0.010518f
C827 B.n787 VSUBS 0.010518f
C828 B.n788 VSUBS 0.010518f
C829 B.n789 VSUBS 0.010518f
C830 B.n790 VSUBS 0.010518f
C831 B.n791 VSUBS 0.023817f
C832 VDD2.n0 VSUBS 0.032469f
C833 VDD2.n1 VSUBS 0.032019f
C834 VDD2.n2 VSUBS 0.017205f
C835 VDD2.n3 VSUBS 0.040668f
C836 VDD2.n4 VSUBS 0.018218f
C837 VDD2.n5 VSUBS 0.032019f
C838 VDD2.n6 VSUBS 0.017205f
C839 VDD2.n7 VSUBS 0.040668f
C840 VDD2.n8 VSUBS 0.018218f
C841 VDD2.n9 VSUBS 0.032019f
C842 VDD2.n10 VSUBS 0.017205f
C843 VDD2.n11 VSUBS 0.040668f
C844 VDD2.n12 VSUBS 0.018218f
C845 VDD2.n13 VSUBS 0.201984f
C846 VDD2.t1 VSUBS 0.087323f
C847 VDD2.n14 VSUBS 0.030501f
C848 VDD2.n15 VSUBS 0.030592f
C849 VDD2.n16 VSUBS 0.017205f
C850 VDD2.n17 VSUBS 1.08625f
C851 VDD2.n18 VSUBS 0.032019f
C852 VDD2.n19 VSUBS 0.017205f
C853 VDD2.n20 VSUBS 0.018218f
C854 VDD2.n21 VSUBS 0.040668f
C855 VDD2.n22 VSUBS 0.040668f
C856 VDD2.n23 VSUBS 0.018218f
C857 VDD2.n24 VSUBS 0.017205f
C858 VDD2.n25 VSUBS 0.032019f
C859 VDD2.n26 VSUBS 0.032019f
C860 VDD2.n27 VSUBS 0.017205f
C861 VDD2.n28 VSUBS 0.018218f
C862 VDD2.n29 VSUBS 0.040668f
C863 VDD2.n30 VSUBS 0.040668f
C864 VDD2.n31 VSUBS 0.040668f
C865 VDD2.n32 VSUBS 0.018218f
C866 VDD2.n33 VSUBS 0.017205f
C867 VDD2.n34 VSUBS 0.032019f
C868 VDD2.n35 VSUBS 0.032019f
C869 VDD2.n36 VSUBS 0.017205f
C870 VDD2.n37 VSUBS 0.017712f
C871 VDD2.n38 VSUBS 0.017712f
C872 VDD2.n39 VSUBS 0.040668f
C873 VDD2.n40 VSUBS 0.089212f
C874 VDD2.n41 VSUBS 0.018218f
C875 VDD2.n42 VSUBS 0.017205f
C876 VDD2.n43 VSUBS 0.074447f
C877 VDD2.n44 VSUBS 0.083034f
C878 VDD2.t6 VSUBS 0.215828f
C879 VDD2.t2 VSUBS 0.215828f
C880 VDD2.n45 VSUBS 1.57882f
C881 VDD2.n46 VSUBS 1.19764f
C882 VDD2.t8 VSUBS 0.215828f
C883 VDD2.t5 VSUBS 0.215828f
C884 VDD2.n47 VSUBS 1.60239f
C885 VDD2.n48 VSUBS 3.78585f
C886 VDD2.n49 VSUBS 0.032469f
C887 VDD2.n50 VSUBS 0.032019f
C888 VDD2.n51 VSUBS 0.017205f
C889 VDD2.n52 VSUBS 0.040668f
C890 VDD2.n53 VSUBS 0.018218f
C891 VDD2.n54 VSUBS 0.032019f
C892 VDD2.n55 VSUBS 0.017205f
C893 VDD2.n56 VSUBS 0.040668f
C894 VDD2.n57 VSUBS 0.040668f
C895 VDD2.n58 VSUBS 0.018218f
C896 VDD2.n59 VSUBS 0.032019f
C897 VDD2.n60 VSUBS 0.017205f
C898 VDD2.n61 VSUBS 0.040668f
C899 VDD2.n62 VSUBS 0.018218f
C900 VDD2.n63 VSUBS 0.201984f
C901 VDD2.t9 VSUBS 0.087323f
C902 VDD2.n64 VSUBS 0.030501f
C903 VDD2.n65 VSUBS 0.030592f
C904 VDD2.n66 VSUBS 0.017205f
C905 VDD2.n67 VSUBS 1.08625f
C906 VDD2.n68 VSUBS 0.032019f
C907 VDD2.n69 VSUBS 0.017205f
C908 VDD2.n70 VSUBS 0.018218f
C909 VDD2.n71 VSUBS 0.040668f
C910 VDD2.n72 VSUBS 0.040668f
C911 VDD2.n73 VSUBS 0.018218f
C912 VDD2.n74 VSUBS 0.017205f
C913 VDD2.n75 VSUBS 0.032019f
C914 VDD2.n76 VSUBS 0.032019f
C915 VDD2.n77 VSUBS 0.017205f
C916 VDD2.n78 VSUBS 0.018218f
C917 VDD2.n79 VSUBS 0.040668f
C918 VDD2.n80 VSUBS 0.040668f
C919 VDD2.n81 VSUBS 0.018218f
C920 VDD2.n82 VSUBS 0.017205f
C921 VDD2.n83 VSUBS 0.032019f
C922 VDD2.n84 VSUBS 0.032019f
C923 VDD2.n85 VSUBS 0.017205f
C924 VDD2.n86 VSUBS 0.017712f
C925 VDD2.n87 VSUBS 0.017712f
C926 VDD2.n88 VSUBS 0.040668f
C927 VDD2.n89 VSUBS 0.089212f
C928 VDD2.n90 VSUBS 0.018218f
C929 VDD2.n91 VSUBS 0.017205f
C930 VDD2.n92 VSUBS 0.074447f
C931 VDD2.n93 VSUBS 0.066572f
C932 VDD2.n94 VSUBS 3.39235f
C933 VDD2.t7 VSUBS 0.215828f
C934 VDD2.t0 VSUBS 0.215828f
C935 VDD2.n95 VSUBS 1.57882f
C936 VDD2.n96 VSUBS 0.895821f
C937 VDD2.t3 VSUBS 0.215828f
C938 VDD2.t4 VSUBS 0.215828f
C939 VDD2.n97 VSUBS 1.60234f
C940 VN.t4 VSUBS 1.9051f
C941 VN.n0 VSUBS 0.809587f
C942 VN.n1 VSUBS 0.031062f
C943 VN.n2 VSUBS 0.061735f
C944 VN.n3 VSUBS 0.031062f
C945 VN.t1 VSUBS 1.9051f
C946 VN.n4 VSUBS 0.061735f
C947 VN.n5 VSUBS 0.031062f
C948 VN.t7 VSUBS 1.9051f
C949 VN.n6 VSUBS 0.718748f
C950 VN.n7 VSUBS 0.031062f
C951 VN.n8 VSUBS 0.061735f
C952 VN.t8 VSUBS 2.16719f
C953 VN.n9 VSUBS 0.75913f
C954 VN.t3 VSUBS 1.9051f
C955 VN.n10 VSUBS 0.798627f
C956 VN.n11 VSUBS 0.057891f
C957 VN.n12 VSUBS 0.321382f
C958 VN.n13 VSUBS 0.031062f
C959 VN.n14 VSUBS 0.031062f
C960 VN.n15 VSUBS 0.025111f
C961 VN.n16 VSUBS 0.061735f
C962 VN.n17 VSUBS 0.057891f
C963 VN.n18 VSUBS 0.031062f
C964 VN.n19 VSUBS 0.031062f
C965 VN.n20 VSUBS 0.031062f
C966 VN.n21 VSUBS 0.057891f
C967 VN.n22 VSUBS 0.061735f
C968 VN.n23 VSUBS 0.025111f
C969 VN.n24 VSUBS 0.031062f
C970 VN.n25 VSUBS 0.031062f
C971 VN.n26 VSUBS 0.031062f
C972 VN.n27 VSUBS 0.057891f
C973 VN.n28 VSUBS 0.718748f
C974 VN.n29 VSUBS 0.057891f
C975 VN.n30 VSUBS 0.031062f
C976 VN.n31 VSUBS 0.031062f
C977 VN.n32 VSUBS 0.031062f
C978 VN.n33 VSUBS 0.025111f
C979 VN.n34 VSUBS 0.061735f
C980 VN.n35 VSUBS 0.057891f
C981 VN.n36 VSUBS 0.050133f
C982 VN.n37 VSUBS 0.055147f
C983 VN.t0 VSUBS 1.9051f
C984 VN.n38 VSUBS 0.809587f
C985 VN.n39 VSUBS 0.031062f
C986 VN.n40 VSUBS 0.061735f
C987 VN.n41 VSUBS 0.031062f
C988 VN.t2 VSUBS 1.9051f
C989 VN.n42 VSUBS 0.061735f
C990 VN.n43 VSUBS 0.031062f
C991 VN.t9 VSUBS 1.9051f
C992 VN.n44 VSUBS 0.718748f
C993 VN.n45 VSUBS 0.031062f
C994 VN.n46 VSUBS 0.061735f
C995 VN.t5 VSUBS 2.16719f
C996 VN.n47 VSUBS 0.75913f
C997 VN.t6 VSUBS 1.9051f
C998 VN.n48 VSUBS 0.798627f
C999 VN.n49 VSUBS 0.057891f
C1000 VN.n50 VSUBS 0.321382f
C1001 VN.n51 VSUBS 0.031062f
C1002 VN.n52 VSUBS 0.031062f
C1003 VN.n53 VSUBS 0.025111f
C1004 VN.n54 VSUBS 0.061735f
C1005 VN.n55 VSUBS 0.057891f
C1006 VN.n56 VSUBS 0.031062f
C1007 VN.n57 VSUBS 0.031062f
C1008 VN.n58 VSUBS 0.031062f
C1009 VN.n59 VSUBS 0.057891f
C1010 VN.n60 VSUBS 0.061735f
C1011 VN.n61 VSUBS 0.025111f
C1012 VN.n62 VSUBS 0.031062f
C1013 VN.n63 VSUBS 0.031062f
C1014 VN.n64 VSUBS 0.031062f
C1015 VN.n65 VSUBS 0.057891f
C1016 VN.n66 VSUBS 0.718748f
C1017 VN.n67 VSUBS 0.057891f
C1018 VN.n68 VSUBS 0.031062f
C1019 VN.n69 VSUBS 0.031062f
C1020 VN.n70 VSUBS 0.031062f
C1021 VN.n71 VSUBS 0.025111f
C1022 VN.n72 VSUBS 0.061735f
C1023 VN.n73 VSUBS 0.057891f
C1024 VN.n74 VSUBS 0.050133f
C1025 VN.n75 VSUBS 1.8069f
C1026 VDD1.n0 VSUBS 0.03231f
C1027 VDD1.n1 VSUBS 0.031862f
C1028 VDD1.n2 VSUBS 0.017121f
C1029 VDD1.n3 VSUBS 0.040468f
C1030 VDD1.n4 VSUBS 0.018128f
C1031 VDD1.n5 VSUBS 0.031862f
C1032 VDD1.n6 VSUBS 0.017121f
C1033 VDD1.n7 VSUBS 0.040468f
C1034 VDD1.n8 VSUBS 0.040468f
C1035 VDD1.n9 VSUBS 0.018128f
C1036 VDD1.n10 VSUBS 0.031862f
C1037 VDD1.n11 VSUBS 0.017121f
C1038 VDD1.n12 VSUBS 0.040468f
C1039 VDD1.n13 VSUBS 0.018128f
C1040 VDD1.n14 VSUBS 0.200993f
C1041 VDD1.t2 VSUBS 0.086894f
C1042 VDD1.n15 VSUBS 0.030351f
C1043 VDD1.n16 VSUBS 0.030442f
C1044 VDD1.n17 VSUBS 0.017121f
C1045 VDD1.n18 VSUBS 1.08092f
C1046 VDD1.n19 VSUBS 0.031862f
C1047 VDD1.n20 VSUBS 0.017121f
C1048 VDD1.n21 VSUBS 0.018128f
C1049 VDD1.n22 VSUBS 0.040468f
C1050 VDD1.n23 VSUBS 0.040468f
C1051 VDD1.n24 VSUBS 0.018128f
C1052 VDD1.n25 VSUBS 0.017121f
C1053 VDD1.n26 VSUBS 0.031862f
C1054 VDD1.n27 VSUBS 0.031862f
C1055 VDD1.n28 VSUBS 0.017121f
C1056 VDD1.n29 VSUBS 0.018128f
C1057 VDD1.n30 VSUBS 0.040468f
C1058 VDD1.n31 VSUBS 0.040468f
C1059 VDD1.n32 VSUBS 0.018128f
C1060 VDD1.n33 VSUBS 0.017121f
C1061 VDD1.n34 VSUBS 0.031862f
C1062 VDD1.n35 VSUBS 0.031862f
C1063 VDD1.n36 VSUBS 0.017121f
C1064 VDD1.n37 VSUBS 0.017625f
C1065 VDD1.n38 VSUBS 0.017625f
C1066 VDD1.n39 VSUBS 0.040468f
C1067 VDD1.n40 VSUBS 0.088774f
C1068 VDD1.n41 VSUBS 0.018128f
C1069 VDD1.n42 VSUBS 0.017121f
C1070 VDD1.n43 VSUBS 0.074082f
C1071 VDD1.n44 VSUBS 0.082627f
C1072 VDD1.t1 VSUBS 0.21477f
C1073 VDD1.t7 VSUBS 0.21477f
C1074 VDD1.n45 VSUBS 1.57108f
C1075 VDD1.n46 VSUBS 1.20216f
C1076 VDD1.n47 VSUBS 0.03231f
C1077 VDD1.n48 VSUBS 0.031862f
C1078 VDD1.n49 VSUBS 0.017121f
C1079 VDD1.n50 VSUBS 0.040468f
C1080 VDD1.n51 VSUBS 0.018128f
C1081 VDD1.n52 VSUBS 0.031862f
C1082 VDD1.n53 VSUBS 0.017121f
C1083 VDD1.n54 VSUBS 0.040468f
C1084 VDD1.n55 VSUBS 0.018128f
C1085 VDD1.n56 VSUBS 0.031862f
C1086 VDD1.n57 VSUBS 0.017121f
C1087 VDD1.n58 VSUBS 0.040468f
C1088 VDD1.n59 VSUBS 0.018128f
C1089 VDD1.n60 VSUBS 0.200993f
C1090 VDD1.t4 VSUBS 0.086894f
C1091 VDD1.n61 VSUBS 0.030351f
C1092 VDD1.n62 VSUBS 0.030442f
C1093 VDD1.n63 VSUBS 0.017121f
C1094 VDD1.n64 VSUBS 1.08092f
C1095 VDD1.n65 VSUBS 0.031862f
C1096 VDD1.n66 VSUBS 0.017121f
C1097 VDD1.n67 VSUBS 0.018128f
C1098 VDD1.n68 VSUBS 0.040468f
C1099 VDD1.n69 VSUBS 0.040468f
C1100 VDD1.n70 VSUBS 0.018128f
C1101 VDD1.n71 VSUBS 0.017121f
C1102 VDD1.n72 VSUBS 0.031862f
C1103 VDD1.n73 VSUBS 0.031862f
C1104 VDD1.n74 VSUBS 0.017121f
C1105 VDD1.n75 VSUBS 0.018128f
C1106 VDD1.n76 VSUBS 0.040468f
C1107 VDD1.n77 VSUBS 0.040468f
C1108 VDD1.n78 VSUBS 0.040468f
C1109 VDD1.n79 VSUBS 0.018128f
C1110 VDD1.n80 VSUBS 0.017121f
C1111 VDD1.n81 VSUBS 0.031862f
C1112 VDD1.n82 VSUBS 0.031862f
C1113 VDD1.n83 VSUBS 0.017121f
C1114 VDD1.n84 VSUBS 0.017625f
C1115 VDD1.n85 VSUBS 0.017625f
C1116 VDD1.n86 VSUBS 0.040468f
C1117 VDD1.n87 VSUBS 0.088774f
C1118 VDD1.n88 VSUBS 0.018128f
C1119 VDD1.n89 VSUBS 0.017121f
C1120 VDD1.n90 VSUBS 0.074082f
C1121 VDD1.n91 VSUBS 0.082627f
C1122 VDD1.t6 VSUBS 0.21477f
C1123 VDD1.t3 VSUBS 0.21477f
C1124 VDD1.n92 VSUBS 1.57107f
C1125 VDD1.n93 VSUBS 1.19177f
C1126 VDD1.t5 VSUBS 0.21477f
C1127 VDD1.t0 VSUBS 0.21477f
C1128 VDD1.n94 VSUBS 1.59454f
C1129 VDD1.n95 VSUBS 3.92571f
C1130 VDD1.t8 VSUBS 0.21477f
C1131 VDD1.t9 VSUBS 0.21477f
C1132 VDD1.n96 VSUBS 1.57107f
C1133 VDD1.n97 VSUBS 4.03294f
C1134 VTAIL.t8 VSUBS 0.207258f
C1135 VTAIL.t4 VSUBS 0.207258f
C1136 VTAIL.n0 VSUBS 1.37804f
C1137 VTAIL.n1 VSUBS 1.00309f
C1138 VTAIL.n2 VSUBS 0.03118f
C1139 VTAIL.n3 VSUBS 0.030747f
C1140 VTAIL.n4 VSUBS 0.016522f
C1141 VTAIL.n5 VSUBS 0.039053f
C1142 VTAIL.n6 VSUBS 0.017494f
C1143 VTAIL.n7 VSUBS 0.030747f
C1144 VTAIL.n8 VSUBS 0.016522f
C1145 VTAIL.n9 VSUBS 0.039053f
C1146 VTAIL.n10 VSUBS 0.017494f
C1147 VTAIL.n11 VSUBS 0.030747f
C1148 VTAIL.n12 VSUBS 0.016522f
C1149 VTAIL.n13 VSUBS 0.039053f
C1150 VTAIL.n14 VSUBS 0.017494f
C1151 VTAIL.n15 VSUBS 0.193963f
C1152 VTAIL.t19 VSUBS 0.083855f
C1153 VTAIL.n16 VSUBS 0.029289f
C1154 VTAIL.n17 VSUBS 0.029377f
C1155 VTAIL.n18 VSUBS 0.016522f
C1156 VTAIL.n19 VSUBS 1.04311f
C1157 VTAIL.n20 VSUBS 0.030747f
C1158 VTAIL.n21 VSUBS 0.016522f
C1159 VTAIL.n22 VSUBS 0.017494f
C1160 VTAIL.n23 VSUBS 0.039053f
C1161 VTAIL.n24 VSUBS 0.039053f
C1162 VTAIL.n25 VSUBS 0.017494f
C1163 VTAIL.n26 VSUBS 0.016522f
C1164 VTAIL.n27 VSUBS 0.030747f
C1165 VTAIL.n28 VSUBS 0.030747f
C1166 VTAIL.n29 VSUBS 0.016522f
C1167 VTAIL.n30 VSUBS 0.017494f
C1168 VTAIL.n31 VSUBS 0.039053f
C1169 VTAIL.n32 VSUBS 0.039053f
C1170 VTAIL.n33 VSUBS 0.039053f
C1171 VTAIL.n34 VSUBS 0.017494f
C1172 VTAIL.n35 VSUBS 0.016522f
C1173 VTAIL.n36 VSUBS 0.030747f
C1174 VTAIL.n37 VSUBS 0.030747f
C1175 VTAIL.n38 VSUBS 0.016522f
C1176 VTAIL.n39 VSUBS 0.017008f
C1177 VTAIL.n40 VSUBS 0.017008f
C1178 VTAIL.n41 VSUBS 0.039053f
C1179 VTAIL.n42 VSUBS 0.085669f
C1180 VTAIL.n43 VSUBS 0.017494f
C1181 VTAIL.n44 VSUBS 0.016522f
C1182 VTAIL.n45 VSUBS 0.071491f
C1183 VTAIL.n46 VSUBS 0.042701f
C1184 VTAIL.n47 VSUBS 0.457388f
C1185 VTAIL.t17 VSUBS 0.207258f
C1186 VTAIL.t14 VSUBS 0.207258f
C1187 VTAIL.n48 VSUBS 1.37804f
C1188 VTAIL.n49 VSUBS 1.14295f
C1189 VTAIL.t18 VSUBS 0.207258f
C1190 VTAIL.t15 VSUBS 0.207258f
C1191 VTAIL.n50 VSUBS 1.37804f
C1192 VTAIL.n51 VSUBS 2.54539f
C1193 VTAIL.t5 VSUBS 0.207258f
C1194 VTAIL.t2 VSUBS 0.207258f
C1195 VTAIL.n52 VSUBS 1.37805f
C1196 VTAIL.n53 VSUBS 2.54538f
C1197 VTAIL.t7 VSUBS 0.207258f
C1198 VTAIL.t3 VSUBS 0.207258f
C1199 VTAIL.n54 VSUBS 1.37805f
C1200 VTAIL.n55 VSUBS 1.14294f
C1201 VTAIL.n56 VSUBS 0.03118f
C1202 VTAIL.n57 VSUBS 0.030747f
C1203 VTAIL.n58 VSUBS 0.016522f
C1204 VTAIL.n59 VSUBS 0.039053f
C1205 VTAIL.n60 VSUBS 0.017494f
C1206 VTAIL.n61 VSUBS 0.030747f
C1207 VTAIL.n62 VSUBS 0.016522f
C1208 VTAIL.n63 VSUBS 0.039053f
C1209 VTAIL.n64 VSUBS 0.039053f
C1210 VTAIL.n65 VSUBS 0.017494f
C1211 VTAIL.n66 VSUBS 0.030747f
C1212 VTAIL.n67 VSUBS 0.016522f
C1213 VTAIL.n68 VSUBS 0.039053f
C1214 VTAIL.n69 VSUBS 0.017494f
C1215 VTAIL.n70 VSUBS 0.193963f
C1216 VTAIL.t9 VSUBS 0.083855f
C1217 VTAIL.n71 VSUBS 0.029289f
C1218 VTAIL.n72 VSUBS 0.029377f
C1219 VTAIL.n73 VSUBS 0.016522f
C1220 VTAIL.n74 VSUBS 1.04311f
C1221 VTAIL.n75 VSUBS 0.030747f
C1222 VTAIL.n76 VSUBS 0.016522f
C1223 VTAIL.n77 VSUBS 0.017494f
C1224 VTAIL.n78 VSUBS 0.039053f
C1225 VTAIL.n79 VSUBS 0.039053f
C1226 VTAIL.n80 VSUBS 0.017494f
C1227 VTAIL.n81 VSUBS 0.016522f
C1228 VTAIL.n82 VSUBS 0.030747f
C1229 VTAIL.n83 VSUBS 0.030747f
C1230 VTAIL.n84 VSUBS 0.016522f
C1231 VTAIL.n85 VSUBS 0.017494f
C1232 VTAIL.n86 VSUBS 0.039053f
C1233 VTAIL.n87 VSUBS 0.039053f
C1234 VTAIL.n88 VSUBS 0.017494f
C1235 VTAIL.n89 VSUBS 0.016522f
C1236 VTAIL.n90 VSUBS 0.030747f
C1237 VTAIL.n91 VSUBS 0.030747f
C1238 VTAIL.n92 VSUBS 0.016522f
C1239 VTAIL.n93 VSUBS 0.017008f
C1240 VTAIL.n94 VSUBS 0.017008f
C1241 VTAIL.n95 VSUBS 0.039053f
C1242 VTAIL.n96 VSUBS 0.085669f
C1243 VTAIL.n97 VSUBS 0.017494f
C1244 VTAIL.n98 VSUBS 0.016522f
C1245 VTAIL.n99 VSUBS 0.071491f
C1246 VTAIL.n100 VSUBS 0.042701f
C1247 VTAIL.n101 VSUBS 0.457388f
C1248 VTAIL.t16 VSUBS 0.207258f
C1249 VTAIL.t13 VSUBS 0.207258f
C1250 VTAIL.n102 VSUBS 1.37805f
C1251 VTAIL.n103 VSUBS 1.06138f
C1252 VTAIL.t10 VSUBS 0.207258f
C1253 VTAIL.t11 VSUBS 0.207258f
C1254 VTAIL.n104 VSUBS 1.37805f
C1255 VTAIL.n105 VSUBS 1.14294f
C1256 VTAIL.n106 VSUBS 0.03118f
C1257 VTAIL.n107 VSUBS 0.030747f
C1258 VTAIL.n108 VSUBS 0.016522f
C1259 VTAIL.n109 VSUBS 0.039053f
C1260 VTAIL.n110 VSUBS 0.017494f
C1261 VTAIL.n111 VSUBS 0.030747f
C1262 VTAIL.n112 VSUBS 0.016522f
C1263 VTAIL.n113 VSUBS 0.039053f
C1264 VTAIL.n114 VSUBS 0.039053f
C1265 VTAIL.n115 VSUBS 0.017494f
C1266 VTAIL.n116 VSUBS 0.030747f
C1267 VTAIL.n117 VSUBS 0.016522f
C1268 VTAIL.n118 VSUBS 0.039053f
C1269 VTAIL.n119 VSUBS 0.017494f
C1270 VTAIL.n120 VSUBS 0.193963f
C1271 VTAIL.t12 VSUBS 0.083855f
C1272 VTAIL.n121 VSUBS 0.029289f
C1273 VTAIL.n122 VSUBS 0.029377f
C1274 VTAIL.n123 VSUBS 0.016522f
C1275 VTAIL.n124 VSUBS 1.04311f
C1276 VTAIL.n125 VSUBS 0.030747f
C1277 VTAIL.n126 VSUBS 0.016522f
C1278 VTAIL.n127 VSUBS 0.017494f
C1279 VTAIL.n128 VSUBS 0.039053f
C1280 VTAIL.n129 VSUBS 0.039053f
C1281 VTAIL.n130 VSUBS 0.017494f
C1282 VTAIL.n131 VSUBS 0.016522f
C1283 VTAIL.n132 VSUBS 0.030747f
C1284 VTAIL.n133 VSUBS 0.030747f
C1285 VTAIL.n134 VSUBS 0.016522f
C1286 VTAIL.n135 VSUBS 0.017494f
C1287 VTAIL.n136 VSUBS 0.039053f
C1288 VTAIL.n137 VSUBS 0.039053f
C1289 VTAIL.n138 VSUBS 0.017494f
C1290 VTAIL.n139 VSUBS 0.016522f
C1291 VTAIL.n140 VSUBS 0.030747f
C1292 VTAIL.n141 VSUBS 0.030747f
C1293 VTAIL.n142 VSUBS 0.016522f
C1294 VTAIL.n143 VSUBS 0.017008f
C1295 VTAIL.n144 VSUBS 0.017008f
C1296 VTAIL.n145 VSUBS 0.039053f
C1297 VTAIL.n146 VSUBS 0.085669f
C1298 VTAIL.n147 VSUBS 0.017494f
C1299 VTAIL.n148 VSUBS 0.016522f
C1300 VTAIL.n149 VSUBS 0.071491f
C1301 VTAIL.n150 VSUBS 0.042701f
C1302 VTAIL.n151 VSUBS 1.68516f
C1303 VTAIL.n152 VSUBS 0.03118f
C1304 VTAIL.n153 VSUBS 0.030747f
C1305 VTAIL.n154 VSUBS 0.016522f
C1306 VTAIL.n155 VSUBS 0.039053f
C1307 VTAIL.n156 VSUBS 0.017494f
C1308 VTAIL.n157 VSUBS 0.030747f
C1309 VTAIL.n158 VSUBS 0.016522f
C1310 VTAIL.n159 VSUBS 0.039053f
C1311 VTAIL.n160 VSUBS 0.017494f
C1312 VTAIL.n161 VSUBS 0.030747f
C1313 VTAIL.n162 VSUBS 0.016522f
C1314 VTAIL.n163 VSUBS 0.039053f
C1315 VTAIL.n164 VSUBS 0.017494f
C1316 VTAIL.n165 VSUBS 0.193963f
C1317 VTAIL.t6 VSUBS 0.083855f
C1318 VTAIL.n166 VSUBS 0.029289f
C1319 VTAIL.n167 VSUBS 0.029377f
C1320 VTAIL.n168 VSUBS 0.016522f
C1321 VTAIL.n169 VSUBS 1.04311f
C1322 VTAIL.n170 VSUBS 0.030747f
C1323 VTAIL.n171 VSUBS 0.016522f
C1324 VTAIL.n172 VSUBS 0.017494f
C1325 VTAIL.n173 VSUBS 0.039053f
C1326 VTAIL.n174 VSUBS 0.039053f
C1327 VTAIL.n175 VSUBS 0.017494f
C1328 VTAIL.n176 VSUBS 0.016522f
C1329 VTAIL.n177 VSUBS 0.030747f
C1330 VTAIL.n178 VSUBS 0.030747f
C1331 VTAIL.n179 VSUBS 0.016522f
C1332 VTAIL.n180 VSUBS 0.017494f
C1333 VTAIL.n181 VSUBS 0.039053f
C1334 VTAIL.n182 VSUBS 0.039053f
C1335 VTAIL.n183 VSUBS 0.039053f
C1336 VTAIL.n184 VSUBS 0.017494f
C1337 VTAIL.n185 VSUBS 0.016522f
C1338 VTAIL.n186 VSUBS 0.030747f
C1339 VTAIL.n187 VSUBS 0.030747f
C1340 VTAIL.n188 VSUBS 0.016522f
C1341 VTAIL.n189 VSUBS 0.017008f
C1342 VTAIL.n190 VSUBS 0.017008f
C1343 VTAIL.n191 VSUBS 0.039053f
C1344 VTAIL.n192 VSUBS 0.085669f
C1345 VTAIL.n193 VSUBS 0.017494f
C1346 VTAIL.n194 VSUBS 0.016522f
C1347 VTAIL.n195 VSUBS 0.071491f
C1348 VTAIL.n196 VSUBS 0.042701f
C1349 VTAIL.n197 VSUBS 1.68516f
C1350 VTAIL.t0 VSUBS 0.207258f
C1351 VTAIL.t1 VSUBS 0.207258f
C1352 VTAIL.n198 VSUBS 1.37804f
C1353 VTAIL.n199 VSUBS 0.945016f
C1354 VP.t9 VSUBS 2.08654f
C1355 VP.n0 VSUBS 0.886695f
C1356 VP.n1 VSUBS 0.03402f
C1357 VP.n2 VSUBS 0.067615f
C1358 VP.n3 VSUBS 0.03402f
C1359 VP.t4 VSUBS 2.08654f
C1360 VP.n4 VSUBS 0.067615f
C1361 VP.n5 VSUBS 0.03402f
C1362 VP.t6 VSUBS 2.08654f
C1363 VP.n6 VSUBS 0.787205f
C1364 VP.n7 VSUBS 0.03402f
C1365 VP.n8 VSUBS 0.067615f
C1366 VP.n9 VSUBS 0.03402f
C1367 VP.t3 VSUBS 2.08654f
C1368 VP.n10 VSUBS 0.067615f
C1369 VP.n11 VSUBS 0.03402f
C1370 VP.t5 VSUBS 2.08654f
C1371 VP.n12 VSUBS 0.886695f
C1372 VP.t0 VSUBS 2.08654f
C1373 VP.n13 VSUBS 0.886695f
C1374 VP.n14 VSUBS 0.03402f
C1375 VP.n15 VSUBS 0.067615f
C1376 VP.n16 VSUBS 0.03402f
C1377 VP.t1 VSUBS 2.08654f
C1378 VP.n17 VSUBS 0.067615f
C1379 VP.n18 VSUBS 0.03402f
C1380 VP.t2 VSUBS 2.08654f
C1381 VP.n19 VSUBS 0.787205f
C1382 VP.n20 VSUBS 0.03402f
C1383 VP.n21 VSUBS 0.067615f
C1384 VP.t7 VSUBS 2.3736f
C1385 VP.n22 VSUBS 0.831433f
C1386 VP.t8 VSUBS 2.08654f
C1387 VP.n23 VSUBS 0.874691f
C1388 VP.n24 VSUBS 0.063405f
C1389 VP.n25 VSUBS 0.351993f
C1390 VP.n26 VSUBS 0.03402f
C1391 VP.n27 VSUBS 0.03402f
C1392 VP.n28 VSUBS 0.027502f
C1393 VP.n29 VSUBS 0.067615f
C1394 VP.n30 VSUBS 0.063405f
C1395 VP.n31 VSUBS 0.03402f
C1396 VP.n32 VSUBS 0.03402f
C1397 VP.n33 VSUBS 0.03402f
C1398 VP.n34 VSUBS 0.063405f
C1399 VP.n35 VSUBS 0.067615f
C1400 VP.n36 VSUBS 0.027502f
C1401 VP.n37 VSUBS 0.03402f
C1402 VP.n38 VSUBS 0.03402f
C1403 VP.n39 VSUBS 0.03402f
C1404 VP.n40 VSUBS 0.063405f
C1405 VP.n41 VSUBS 0.787205f
C1406 VP.n42 VSUBS 0.063405f
C1407 VP.n43 VSUBS 0.03402f
C1408 VP.n44 VSUBS 0.03402f
C1409 VP.n45 VSUBS 0.03402f
C1410 VP.n46 VSUBS 0.027502f
C1411 VP.n47 VSUBS 0.067615f
C1412 VP.n48 VSUBS 0.063405f
C1413 VP.n49 VSUBS 0.054908f
C1414 VP.n50 VSUBS 1.96516f
C1415 VP.n51 VSUBS 1.98915f
C1416 VP.n52 VSUBS 0.054908f
C1417 VP.n53 VSUBS 0.063405f
C1418 VP.n54 VSUBS 0.067615f
C1419 VP.n55 VSUBS 0.027502f
C1420 VP.n56 VSUBS 0.03402f
C1421 VP.n57 VSUBS 0.03402f
C1422 VP.n58 VSUBS 0.03402f
C1423 VP.n59 VSUBS 0.063405f
C1424 VP.n60 VSUBS 0.787205f
C1425 VP.n61 VSUBS 0.063405f
C1426 VP.n62 VSUBS 0.03402f
C1427 VP.n63 VSUBS 0.03402f
C1428 VP.n64 VSUBS 0.03402f
C1429 VP.n65 VSUBS 0.027502f
C1430 VP.n66 VSUBS 0.067615f
C1431 VP.n67 VSUBS 0.063405f
C1432 VP.n68 VSUBS 0.03402f
C1433 VP.n69 VSUBS 0.03402f
C1434 VP.n70 VSUBS 0.03402f
C1435 VP.n71 VSUBS 0.063405f
C1436 VP.n72 VSUBS 0.067615f
C1437 VP.n73 VSUBS 0.027502f
C1438 VP.n74 VSUBS 0.03402f
C1439 VP.n75 VSUBS 0.03402f
C1440 VP.n76 VSUBS 0.03402f
C1441 VP.n77 VSUBS 0.063405f
C1442 VP.n78 VSUBS 0.787205f
C1443 VP.n79 VSUBS 0.063405f
C1444 VP.n80 VSUBS 0.03402f
C1445 VP.n81 VSUBS 0.03402f
C1446 VP.n82 VSUBS 0.03402f
C1447 VP.n83 VSUBS 0.027502f
C1448 VP.n84 VSUBS 0.067615f
C1449 VP.n85 VSUBS 0.063405f
C1450 VP.n86 VSUBS 0.054908f
C1451 VP.n87 VSUBS 0.0604f
.ends

