* NGSPICE file created from diff_pair_sample_0595.ext - technology: sky130A

.subckt diff_pair_sample_0595 VTAIL VN VP B VDD2 VDD1
X0 B.t17 B.t15 B.t16 B.t12 sky130_fd_pr__nfet_01v8 ad=2.9367 pd=15.84 as=0 ps=0 w=7.53 l=0.75
X1 B.t14 B.t11 B.t13 B.t12 sky130_fd_pr__nfet_01v8 ad=2.9367 pd=15.84 as=0 ps=0 w=7.53 l=0.75
X2 VDD1.t3 VP.t0 VTAIL.t7 B.t3 sky130_fd_pr__nfet_01v8 ad=1.24245 pd=7.86 as=2.9367 ps=15.84 w=7.53 l=0.75
X3 VTAIL.t6 VP.t1 VDD1.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=2.9367 pd=15.84 as=1.24245 ps=7.86 w=7.53 l=0.75
X4 B.t10 B.t8 B.t9 B.t5 sky130_fd_pr__nfet_01v8 ad=2.9367 pd=15.84 as=0 ps=0 w=7.53 l=0.75
X5 VDD2.t3 VN.t0 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=1.24245 pd=7.86 as=2.9367 ps=15.84 w=7.53 l=0.75
X6 VTAIL.t3 VN.t1 VDD2.t2 B.t1 sky130_fd_pr__nfet_01v8 ad=2.9367 pd=15.84 as=1.24245 ps=7.86 w=7.53 l=0.75
X7 VDD1.t1 VP.t2 VTAIL.t5 B.t0 sky130_fd_pr__nfet_01v8 ad=1.24245 pd=7.86 as=2.9367 ps=15.84 w=7.53 l=0.75
X8 VDD2.t1 VN.t2 VTAIL.t2 B.t3 sky130_fd_pr__nfet_01v8 ad=1.24245 pd=7.86 as=2.9367 ps=15.84 w=7.53 l=0.75
X9 VTAIL.t1 VN.t3 VDD2.t0 B.t2 sky130_fd_pr__nfet_01v8 ad=2.9367 pd=15.84 as=1.24245 ps=7.86 w=7.53 l=0.75
X10 B.t7 B.t4 B.t6 B.t5 sky130_fd_pr__nfet_01v8 ad=2.9367 pd=15.84 as=0 ps=0 w=7.53 l=0.75
X11 VTAIL.t4 VP.t3 VDD1.t0 B.t1 sky130_fd_pr__nfet_01v8 ad=2.9367 pd=15.84 as=1.24245 ps=7.86 w=7.53 l=0.75
R0 B.n488 B.n487 585
R1 B.n489 B.n488 585
R2 B.n206 B.n69 585
R3 B.n205 B.n204 585
R4 B.n203 B.n202 585
R5 B.n201 B.n200 585
R6 B.n199 B.n198 585
R7 B.n197 B.n196 585
R8 B.n195 B.n194 585
R9 B.n193 B.n192 585
R10 B.n191 B.n190 585
R11 B.n189 B.n188 585
R12 B.n187 B.n186 585
R13 B.n185 B.n184 585
R14 B.n183 B.n182 585
R15 B.n181 B.n180 585
R16 B.n179 B.n178 585
R17 B.n177 B.n176 585
R18 B.n175 B.n174 585
R19 B.n173 B.n172 585
R20 B.n171 B.n170 585
R21 B.n169 B.n168 585
R22 B.n167 B.n166 585
R23 B.n165 B.n164 585
R24 B.n163 B.n162 585
R25 B.n161 B.n160 585
R26 B.n159 B.n158 585
R27 B.n157 B.n156 585
R28 B.n155 B.n154 585
R29 B.n153 B.n152 585
R30 B.n151 B.n150 585
R31 B.n149 B.n148 585
R32 B.n147 B.n146 585
R33 B.n145 B.n144 585
R34 B.n143 B.n142 585
R35 B.n141 B.n140 585
R36 B.n139 B.n138 585
R37 B.n137 B.n136 585
R38 B.n135 B.n134 585
R39 B.n132 B.n131 585
R40 B.n130 B.n129 585
R41 B.n128 B.n127 585
R42 B.n126 B.n125 585
R43 B.n124 B.n123 585
R44 B.n122 B.n121 585
R45 B.n120 B.n119 585
R46 B.n118 B.n117 585
R47 B.n116 B.n115 585
R48 B.n114 B.n113 585
R49 B.n112 B.n111 585
R50 B.n110 B.n109 585
R51 B.n108 B.n107 585
R52 B.n106 B.n105 585
R53 B.n104 B.n103 585
R54 B.n102 B.n101 585
R55 B.n100 B.n99 585
R56 B.n98 B.n97 585
R57 B.n96 B.n95 585
R58 B.n94 B.n93 585
R59 B.n92 B.n91 585
R60 B.n90 B.n89 585
R61 B.n88 B.n87 585
R62 B.n86 B.n85 585
R63 B.n84 B.n83 585
R64 B.n82 B.n81 585
R65 B.n80 B.n79 585
R66 B.n78 B.n77 585
R67 B.n76 B.n75 585
R68 B.n486 B.n35 585
R69 B.n490 B.n35 585
R70 B.n485 B.n34 585
R71 B.n491 B.n34 585
R72 B.n484 B.n483 585
R73 B.n483 B.n30 585
R74 B.n482 B.n29 585
R75 B.n497 B.n29 585
R76 B.n481 B.n28 585
R77 B.n498 B.n28 585
R78 B.n480 B.n27 585
R79 B.n499 B.n27 585
R80 B.n479 B.n478 585
R81 B.n478 B.n23 585
R82 B.n477 B.n22 585
R83 B.n505 B.n22 585
R84 B.n476 B.n21 585
R85 B.n506 B.n21 585
R86 B.n475 B.n20 585
R87 B.n507 B.n20 585
R88 B.n474 B.n473 585
R89 B.n473 B.n16 585
R90 B.n472 B.n15 585
R91 B.n513 B.n15 585
R92 B.n471 B.n14 585
R93 B.n514 B.n14 585
R94 B.n470 B.n13 585
R95 B.n515 B.n13 585
R96 B.n469 B.n468 585
R97 B.n468 B.n12 585
R98 B.n467 B.n466 585
R99 B.n467 B.n8 585
R100 B.n465 B.n7 585
R101 B.n522 B.n7 585
R102 B.n464 B.n6 585
R103 B.n523 B.n6 585
R104 B.n463 B.n5 585
R105 B.n524 B.n5 585
R106 B.n462 B.n461 585
R107 B.n461 B.n4 585
R108 B.n460 B.n207 585
R109 B.n460 B.n459 585
R110 B.n449 B.n208 585
R111 B.n452 B.n208 585
R112 B.n451 B.n450 585
R113 B.n453 B.n451 585
R114 B.n448 B.n213 585
R115 B.n213 B.n212 585
R116 B.n447 B.n446 585
R117 B.n446 B.n445 585
R118 B.n215 B.n214 585
R119 B.n216 B.n215 585
R120 B.n438 B.n437 585
R121 B.n439 B.n438 585
R122 B.n436 B.n221 585
R123 B.n221 B.n220 585
R124 B.n435 B.n434 585
R125 B.n434 B.n433 585
R126 B.n223 B.n222 585
R127 B.n224 B.n223 585
R128 B.n426 B.n425 585
R129 B.n427 B.n426 585
R130 B.n424 B.n228 585
R131 B.n232 B.n228 585
R132 B.n423 B.n422 585
R133 B.n422 B.n421 585
R134 B.n230 B.n229 585
R135 B.n231 B.n230 585
R136 B.n414 B.n413 585
R137 B.n415 B.n414 585
R138 B.n412 B.n237 585
R139 B.n237 B.n236 585
R140 B.n406 B.n405 585
R141 B.n404 B.n272 585
R142 B.n403 B.n271 585
R143 B.n408 B.n271 585
R144 B.n402 B.n401 585
R145 B.n400 B.n399 585
R146 B.n398 B.n397 585
R147 B.n396 B.n395 585
R148 B.n394 B.n393 585
R149 B.n392 B.n391 585
R150 B.n390 B.n389 585
R151 B.n388 B.n387 585
R152 B.n386 B.n385 585
R153 B.n384 B.n383 585
R154 B.n382 B.n381 585
R155 B.n380 B.n379 585
R156 B.n378 B.n377 585
R157 B.n376 B.n375 585
R158 B.n374 B.n373 585
R159 B.n372 B.n371 585
R160 B.n370 B.n369 585
R161 B.n368 B.n367 585
R162 B.n366 B.n365 585
R163 B.n364 B.n363 585
R164 B.n362 B.n361 585
R165 B.n360 B.n359 585
R166 B.n358 B.n357 585
R167 B.n356 B.n355 585
R168 B.n354 B.n353 585
R169 B.n352 B.n351 585
R170 B.n350 B.n349 585
R171 B.n348 B.n347 585
R172 B.n346 B.n345 585
R173 B.n344 B.n343 585
R174 B.n342 B.n341 585
R175 B.n340 B.n339 585
R176 B.n338 B.n337 585
R177 B.n336 B.n335 585
R178 B.n334 B.n333 585
R179 B.n331 B.n330 585
R180 B.n329 B.n328 585
R181 B.n327 B.n326 585
R182 B.n325 B.n324 585
R183 B.n323 B.n322 585
R184 B.n321 B.n320 585
R185 B.n319 B.n318 585
R186 B.n317 B.n316 585
R187 B.n315 B.n314 585
R188 B.n313 B.n312 585
R189 B.n311 B.n310 585
R190 B.n309 B.n308 585
R191 B.n307 B.n306 585
R192 B.n305 B.n304 585
R193 B.n303 B.n302 585
R194 B.n301 B.n300 585
R195 B.n299 B.n298 585
R196 B.n297 B.n296 585
R197 B.n295 B.n294 585
R198 B.n293 B.n292 585
R199 B.n291 B.n290 585
R200 B.n289 B.n288 585
R201 B.n287 B.n286 585
R202 B.n285 B.n284 585
R203 B.n283 B.n282 585
R204 B.n281 B.n280 585
R205 B.n279 B.n278 585
R206 B.n239 B.n238 585
R207 B.n411 B.n410 585
R208 B.n235 B.n234 585
R209 B.n236 B.n235 585
R210 B.n417 B.n416 585
R211 B.n416 B.n415 585
R212 B.n418 B.n233 585
R213 B.n233 B.n231 585
R214 B.n420 B.n419 585
R215 B.n421 B.n420 585
R216 B.n227 B.n226 585
R217 B.n232 B.n227 585
R218 B.n429 B.n428 585
R219 B.n428 B.n427 585
R220 B.n430 B.n225 585
R221 B.n225 B.n224 585
R222 B.n432 B.n431 585
R223 B.n433 B.n432 585
R224 B.n219 B.n218 585
R225 B.n220 B.n219 585
R226 B.n441 B.n440 585
R227 B.n440 B.n439 585
R228 B.n442 B.n217 585
R229 B.n217 B.n216 585
R230 B.n444 B.n443 585
R231 B.n445 B.n444 585
R232 B.n211 B.n210 585
R233 B.n212 B.n211 585
R234 B.n455 B.n454 585
R235 B.n454 B.n453 585
R236 B.n456 B.n209 585
R237 B.n452 B.n209 585
R238 B.n458 B.n457 585
R239 B.n459 B.n458 585
R240 B.n3 B.n0 585
R241 B.n4 B.n3 585
R242 B.n521 B.n1 585
R243 B.n522 B.n521 585
R244 B.n520 B.n519 585
R245 B.n520 B.n8 585
R246 B.n518 B.n9 585
R247 B.n12 B.n9 585
R248 B.n517 B.n516 585
R249 B.n516 B.n515 585
R250 B.n11 B.n10 585
R251 B.n514 B.n11 585
R252 B.n512 B.n511 585
R253 B.n513 B.n512 585
R254 B.n510 B.n17 585
R255 B.n17 B.n16 585
R256 B.n509 B.n508 585
R257 B.n508 B.n507 585
R258 B.n19 B.n18 585
R259 B.n506 B.n19 585
R260 B.n504 B.n503 585
R261 B.n505 B.n504 585
R262 B.n502 B.n24 585
R263 B.n24 B.n23 585
R264 B.n501 B.n500 585
R265 B.n500 B.n499 585
R266 B.n26 B.n25 585
R267 B.n498 B.n26 585
R268 B.n496 B.n495 585
R269 B.n497 B.n496 585
R270 B.n494 B.n31 585
R271 B.n31 B.n30 585
R272 B.n493 B.n492 585
R273 B.n492 B.n491 585
R274 B.n33 B.n32 585
R275 B.n490 B.n33 585
R276 B.n525 B.n524 585
R277 B.n523 B.n2 585
R278 B.n75 B.n33 482.89
R279 B.n488 B.n35 482.89
R280 B.n410 B.n237 482.89
R281 B.n406 B.n235 482.89
R282 B.n70 B.t11 445.086
R283 B.n276 B.t4 445.086
R284 B.n73 B.t15 444.676
R285 B.n273 B.t8 444.676
R286 B.n489 B.n68 256.663
R287 B.n489 B.n67 256.663
R288 B.n489 B.n66 256.663
R289 B.n489 B.n65 256.663
R290 B.n489 B.n64 256.663
R291 B.n489 B.n63 256.663
R292 B.n489 B.n62 256.663
R293 B.n489 B.n61 256.663
R294 B.n489 B.n60 256.663
R295 B.n489 B.n59 256.663
R296 B.n489 B.n58 256.663
R297 B.n489 B.n57 256.663
R298 B.n489 B.n56 256.663
R299 B.n489 B.n55 256.663
R300 B.n489 B.n54 256.663
R301 B.n489 B.n53 256.663
R302 B.n489 B.n52 256.663
R303 B.n489 B.n51 256.663
R304 B.n489 B.n50 256.663
R305 B.n489 B.n49 256.663
R306 B.n489 B.n48 256.663
R307 B.n489 B.n47 256.663
R308 B.n489 B.n46 256.663
R309 B.n489 B.n45 256.663
R310 B.n489 B.n44 256.663
R311 B.n489 B.n43 256.663
R312 B.n489 B.n42 256.663
R313 B.n489 B.n41 256.663
R314 B.n489 B.n40 256.663
R315 B.n489 B.n39 256.663
R316 B.n489 B.n38 256.663
R317 B.n489 B.n37 256.663
R318 B.n489 B.n36 256.663
R319 B.n408 B.n407 256.663
R320 B.n408 B.n240 256.663
R321 B.n408 B.n241 256.663
R322 B.n408 B.n242 256.663
R323 B.n408 B.n243 256.663
R324 B.n408 B.n244 256.663
R325 B.n408 B.n245 256.663
R326 B.n408 B.n246 256.663
R327 B.n408 B.n247 256.663
R328 B.n408 B.n248 256.663
R329 B.n408 B.n249 256.663
R330 B.n408 B.n250 256.663
R331 B.n408 B.n251 256.663
R332 B.n408 B.n252 256.663
R333 B.n408 B.n253 256.663
R334 B.n408 B.n254 256.663
R335 B.n408 B.n255 256.663
R336 B.n408 B.n256 256.663
R337 B.n408 B.n257 256.663
R338 B.n408 B.n258 256.663
R339 B.n408 B.n259 256.663
R340 B.n408 B.n260 256.663
R341 B.n408 B.n261 256.663
R342 B.n408 B.n262 256.663
R343 B.n408 B.n263 256.663
R344 B.n408 B.n264 256.663
R345 B.n408 B.n265 256.663
R346 B.n408 B.n266 256.663
R347 B.n408 B.n267 256.663
R348 B.n408 B.n268 256.663
R349 B.n408 B.n269 256.663
R350 B.n408 B.n270 256.663
R351 B.n409 B.n408 256.663
R352 B.n527 B.n526 256.663
R353 B.n79 B.n78 163.367
R354 B.n83 B.n82 163.367
R355 B.n87 B.n86 163.367
R356 B.n91 B.n90 163.367
R357 B.n95 B.n94 163.367
R358 B.n99 B.n98 163.367
R359 B.n103 B.n102 163.367
R360 B.n107 B.n106 163.367
R361 B.n111 B.n110 163.367
R362 B.n115 B.n114 163.367
R363 B.n119 B.n118 163.367
R364 B.n123 B.n122 163.367
R365 B.n127 B.n126 163.367
R366 B.n131 B.n130 163.367
R367 B.n136 B.n135 163.367
R368 B.n140 B.n139 163.367
R369 B.n144 B.n143 163.367
R370 B.n148 B.n147 163.367
R371 B.n152 B.n151 163.367
R372 B.n156 B.n155 163.367
R373 B.n160 B.n159 163.367
R374 B.n164 B.n163 163.367
R375 B.n168 B.n167 163.367
R376 B.n172 B.n171 163.367
R377 B.n176 B.n175 163.367
R378 B.n180 B.n179 163.367
R379 B.n184 B.n183 163.367
R380 B.n188 B.n187 163.367
R381 B.n192 B.n191 163.367
R382 B.n196 B.n195 163.367
R383 B.n200 B.n199 163.367
R384 B.n204 B.n203 163.367
R385 B.n488 B.n69 163.367
R386 B.n414 B.n237 163.367
R387 B.n414 B.n230 163.367
R388 B.n422 B.n230 163.367
R389 B.n422 B.n228 163.367
R390 B.n426 B.n228 163.367
R391 B.n426 B.n223 163.367
R392 B.n434 B.n223 163.367
R393 B.n434 B.n221 163.367
R394 B.n438 B.n221 163.367
R395 B.n438 B.n215 163.367
R396 B.n446 B.n215 163.367
R397 B.n446 B.n213 163.367
R398 B.n451 B.n213 163.367
R399 B.n451 B.n208 163.367
R400 B.n460 B.n208 163.367
R401 B.n461 B.n460 163.367
R402 B.n461 B.n5 163.367
R403 B.n6 B.n5 163.367
R404 B.n7 B.n6 163.367
R405 B.n467 B.n7 163.367
R406 B.n468 B.n467 163.367
R407 B.n468 B.n13 163.367
R408 B.n14 B.n13 163.367
R409 B.n15 B.n14 163.367
R410 B.n473 B.n15 163.367
R411 B.n473 B.n20 163.367
R412 B.n21 B.n20 163.367
R413 B.n22 B.n21 163.367
R414 B.n478 B.n22 163.367
R415 B.n478 B.n27 163.367
R416 B.n28 B.n27 163.367
R417 B.n29 B.n28 163.367
R418 B.n483 B.n29 163.367
R419 B.n483 B.n34 163.367
R420 B.n35 B.n34 163.367
R421 B.n272 B.n271 163.367
R422 B.n401 B.n271 163.367
R423 B.n399 B.n398 163.367
R424 B.n395 B.n394 163.367
R425 B.n391 B.n390 163.367
R426 B.n387 B.n386 163.367
R427 B.n383 B.n382 163.367
R428 B.n379 B.n378 163.367
R429 B.n375 B.n374 163.367
R430 B.n371 B.n370 163.367
R431 B.n367 B.n366 163.367
R432 B.n363 B.n362 163.367
R433 B.n359 B.n358 163.367
R434 B.n355 B.n354 163.367
R435 B.n351 B.n350 163.367
R436 B.n347 B.n346 163.367
R437 B.n343 B.n342 163.367
R438 B.n339 B.n338 163.367
R439 B.n335 B.n334 163.367
R440 B.n330 B.n329 163.367
R441 B.n326 B.n325 163.367
R442 B.n322 B.n321 163.367
R443 B.n318 B.n317 163.367
R444 B.n314 B.n313 163.367
R445 B.n310 B.n309 163.367
R446 B.n306 B.n305 163.367
R447 B.n302 B.n301 163.367
R448 B.n298 B.n297 163.367
R449 B.n294 B.n293 163.367
R450 B.n290 B.n289 163.367
R451 B.n286 B.n285 163.367
R452 B.n282 B.n281 163.367
R453 B.n278 B.n239 163.367
R454 B.n416 B.n235 163.367
R455 B.n416 B.n233 163.367
R456 B.n420 B.n233 163.367
R457 B.n420 B.n227 163.367
R458 B.n428 B.n227 163.367
R459 B.n428 B.n225 163.367
R460 B.n432 B.n225 163.367
R461 B.n432 B.n219 163.367
R462 B.n440 B.n219 163.367
R463 B.n440 B.n217 163.367
R464 B.n444 B.n217 163.367
R465 B.n444 B.n211 163.367
R466 B.n454 B.n211 163.367
R467 B.n454 B.n209 163.367
R468 B.n458 B.n209 163.367
R469 B.n458 B.n3 163.367
R470 B.n525 B.n3 163.367
R471 B.n521 B.n2 163.367
R472 B.n521 B.n520 163.367
R473 B.n520 B.n9 163.367
R474 B.n516 B.n9 163.367
R475 B.n516 B.n11 163.367
R476 B.n512 B.n11 163.367
R477 B.n512 B.n17 163.367
R478 B.n508 B.n17 163.367
R479 B.n508 B.n19 163.367
R480 B.n504 B.n19 163.367
R481 B.n504 B.n24 163.367
R482 B.n500 B.n24 163.367
R483 B.n500 B.n26 163.367
R484 B.n496 B.n26 163.367
R485 B.n496 B.n31 163.367
R486 B.n492 B.n31 163.367
R487 B.n492 B.n33 163.367
R488 B.n408 B.n236 114.252
R489 B.n490 B.n489 114.252
R490 B.n70 B.t13 90.8734
R491 B.n276 B.t7 90.8734
R492 B.n73 B.t16 90.8646
R493 B.n273 B.t10 90.8646
R494 B.n75 B.n36 71.676
R495 B.n79 B.n37 71.676
R496 B.n83 B.n38 71.676
R497 B.n87 B.n39 71.676
R498 B.n91 B.n40 71.676
R499 B.n95 B.n41 71.676
R500 B.n99 B.n42 71.676
R501 B.n103 B.n43 71.676
R502 B.n107 B.n44 71.676
R503 B.n111 B.n45 71.676
R504 B.n115 B.n46 71.676
R505 B.n119 B.n47 71.676
R506 B.n123 B.n48 71.676
R507 B.n127 B.n49 71.676
R508 B.n131 B.n50 71.676
R509 B.n136 B.n51 71.676
R510 B.n140 B.n52 71.676
R511 B.n144 B.n53 71.676
R512 B.n148 B.n54 71.676
R513 B.n152 B.n55 71.676
R514 B.n156 B.n56 71.676
R515 B.n160 B.n57 71.676
R516 B.n164 B.n58 71.676
R517 B.n168 B.n59 71.676
R518 B.n172 B.n60 71.676
R519 B.n176 B.n61 71.676
R520 B.n180 B.n62 71.676
R521 B.n184 B.n63 71.676
R522 B.n188 B.n64 71.676
R523 B.n192 B.n65 71.676
R524 B.n196 B.n66 71.676
R525 B.n200 B.n67 71.676
R526 B.n204 B.n68 71.676
R527 B.n69 B.n68 71.676
R528 B.n203 B.n67 71.676
R529 B.n199 B.n66 71.676
R530 B.n195 B.n65 71.676
R531 B.n191 B.n64 71.676
R532 B.n187 B.n63 71.676
R533 B.n183 B.n62 71.676
R534 B.n179 B.n61 71.676
R535 B.n175 B.n60 71.676
R536 B.n171 B.n59 71.676
R537 B.n167 B.n58 71.676
R538 B.n163 B.n57 71.676
R539 B.n159 B.n56 71.676
R540 B.n155 B.n55 71.676
R541 B.n151 B.n54 71.676
R542 B.n147 B.n53 71.676
R543 B.n143 B.n52 71.676
R544 B.n139 B.n51 71.676
R545 B.n135 B.n50 71.676
R546 B.n130 B.n49 71.676
R547 B.n126 B.n48 71.676
R548 B.n122 B.n47 71.676
R549 B.n118 B.n46 71.676
R550 B.n114 B.n45 71.676
R551 B.n110 B.n44 71.676
R552 B.n106 B.n43 71.676
R553 B.n102 B.n42 71.676
R554 B.n98 B.n41 71.676
R555 B.n94 B.n40 71.676
R556 B.n90 B.n39 71.676
R557 B.n86 B.n38 71.676
R558 B.n82 B.n37 71.676
R559 B.n78 B.n36 71.676
R560 B.n407 B.n406 71.676
R561 B.n401 B.n240 71.676
R562 B.n398 B.n241 71.676
R563 B.n394 B.n242 71.676
R564 B.n390 B.n243 71.676
R565 B.n386 B.n244 71.676
R566 B.n382 B.n245 71.676
R567 B.n378 B.n246 71.676
R568 B.n374 B.n247 71.676
R569 B.n370 B.n248 71.676
R570 B.n366 B.n249 71.676
R571 B.n362 B.n250 71.676
R572 B.n358 B.n251 71.676
R573 B.n354 B.n252 71.676
R574 B.n350 B.n253 71.676
R575 B.n346 B.n254 71.676
R576 B.n342 B.n255 71.676
R577 B.n338 B.n256 71.676
R578 B.n334 B.n257 71.676
R579 B.n329 B.n258 71.676
R580 B.n325 B.n259 71.676
R581 B.n321 B.n260 71.676
R582 B.n317 B.n261 71.676
R583 B.n313 B.n262 71.676
R584 B.n309 B.n263 71.676
R585 B.n305 B.n264 71.676
R586 B.n301 B.n265 71.676
R587 B.n297 B.n266 71.676
R588 B.n293 B.n267 71.676
R589 B.n289 B.n268 71.676
R590 B.n285 B.n269 71.676
R591 B.n281 B.n270 71.676
R592 B.n409 B.n239 71.676
R593 B.n407 B.n272 71.676
R594 B.n399 B.n240 71.676
R595 B.n395 B.n241 71.676
R596 B.n391 B.n242 71.676
R597 B.n387 B.n243 71.676
R598 B.n383 B.n244 71.676
R599 B.n379 B.n245 71.676
R600 B.n375 B.n246 71.676
R601 B.n371 B.n247 71.676
R602 B.n367 B.n248 71.676
R603 B.n363 B.n249 71.676
R604 B.n359 B.n250 71.676
R605 B.n355 B.n251 71.676
R606 B.n351 B.n252 71.676
R607 B.n347 B.n253 71.676
R608 B.n343 B.n254 71.676
R609 B.n339 B.n255 71.676
R610 B.n335 B.n256 71.676
R611 B.n330 B.n257 71.676
R612 B.n326 B.n258 71.676
R613 B.n322 B.n259 71.676
R614 B.n318 B.n260 71.676
R615 B.n314 B.n261 71.676
R616 B.n310 B.n262 71.676
R617 B.n306 B.n263 71.676
R618 B.n302 B.n264 71.676
R619 B.n298 B.n265 71.676
R620 B.n294 B.n266 71.676
R621 B.n290 B.n267 71.676
R622 B.n286 B.n268 71.676
R623 B.n282 B.n269 71.676
R624 B.n278 B.n270 71.676
R625 B.n410 B.n409 71.676
R626 B.n526 B.n525 71.676
R627 B.n526 B.n2 71.676
R628 B.n71 B.t14 69.9279
R629 B.n277 B.t6 69.9279
R630 B.n74 B.t17 69.9192
R631 B.n274 B.t9 69.9192
R632 B.n133 B.n74 59.5399
R633 B.n72 B.n71 59.5399
R634 B.n332 B.n277 59.5399
R635 B.n275 B.n274 59.5399
R636 B.n415 B.n236 58.4152
R637 B.n415 B.n231 58.4152
R638 B.n421 B.n231 58.4152
R639 B.n421 B.n232 58.4152
R640 B.n427 B.n224 58.4152
R641 B.n433 B.n224 58.4152
R642 B.n433 B.n220 58.4152
R643 B.n439 B.n220 58.4152
R644 B.n439 B.n216 58.4152
R645 B.n445 B.n216 58.4152
R646 B.n453 B.n212 58.4152
R647 B.n453 B.n452 58.4152
R648 B.n459 B.n4 58.4152
R649 B.n524 B.n4 58.4152
R650 B.n524 B.n523 58.4152
R651 B.n523 B.n522 58.4152
R652 B.n522 B.n8 58.4152
R653 B.n515 B.n12 58.4152
R654 B.n515 B.n514 58.4152
R655 B.n513 B.n16 58.4152
R656 B.n507 B.n16 58.4152
R657 B.n507 B.n506 58.4152
R658 B.n506 B.n505 58.4152
R659 B.n505 B.n23 58.4152
R660 B.n499 B.n23 58.4152
R661 B.n498 B.n497 58.4152
R662 B.n497 B.n30 58.4152
R663 B.n491 B.n30 58.4152
R664 B.n491 B.n490 58.4152
R665 B.t2 B.n212 50.6838
R666 B.n514 B.t3 50.6838
R667 B.n232 B.t5 43.8115
R668 B.t12 B.n498 43.8115
R669 B.n459 B.t0 40.3754
R670 B.t1 B.n8 40.3754
R671 B.n405 B.n234 31.3761
R672 B.n412 B.n411 31.3761
R673 B.n487 B.n486 31.3761
R674 B.n76 B.n32 31.3761
R675 B.n74 B.n73 20.946
R676 B.n71 B.n70 20.946
R677 B.n277 B.n276 20.946
R678 B.n274 B.n273 20.946
R679 B B.n527 18.0485
R680 B.n452 B.t0 18.0403
R681 B.n12 B.t1 18.0403
R682 B.n427 B.t5 14.6042
R683 B.n499 B.t12 14.6042
R684 B.n417 B.n234 10.6151
R685 B.n418 B.n417 10.6151
R686 B.n419 B.n418 10.6151
R687 B.n419 B.n226 10.6151
R688 B.n429 B.n226 10.6151
R689 B.n430 B.n429 10.6151
R690 B.n431 B.n430 10.6151
R691 B.n431 B.n218 10.6151
R692 B.n441 B.n218 10.6151
R693 B.n442 B.n441 10.6151
R694 B.n443 B.n442 10.6151
R695 B.n443 B.n210 10.6151
R696 B.n455 B.n210 10.6151
R697 B.n456 B.n455 10.6151
R698 B.n457 B.n456 10.6151
R699 B.n457 B.n0 10.6151
R700 B.n405 B.n404 10.6151
R701 B.n404 B.n403 10.6151
R702 B.n403 B.n402 10.6151
R703 B.n402 B.n400 10.6151
R704 B.n400 B.n397 10.6151
R705 B.n397 B.n396 10.6151
R706 B.n396 B.n393 10.6151
R707 B.n393 B.n392 10.6151
R708 B.n392 B.n389 10.6151
R709 B.n389 B.n388 10.6151
R710 B.n388 B.n385 10.6151
R711 B.n385 B.n384 10.6151
R712 B.n384 B.n381 10.6151
R713 B.n381 B.n380 10.6151
R714 B.n380 B.n377 10.6151
R715 B.n377 B.n376 10.6151
R716 B.n376 B.n373 10.6151
R717 B.n373 B.n372 10.6151
R718 B.n372 B.n369 10.6151
R719 B.n369 B.n368 10.6151
R720 B.n368 B.n365 10.6151
R721 B.n365 B.n364 10.6151
R722 B.n364 B.n361 10.6151
R723 B.n361 B.n360 10.6151
R724 B.n360 B.n357 10.6151
R725 B.n357 B.n356 10.6151
R726 B.n356 B.n353 10.6151
R727 B.n353 B.n352 10.6151
R728 B.n349 B.n348 10.6151
R729 B.n348 B.n345 10.6151
R730 B.n345 B.n344 10.6151
R731 B.n344 B.n341 10.6151
R732 B.n341 B.n340 10.6151
R733 B.n340 B.n337 10.6151
R734 B.n337 B.n336 10.6151
R735 B.n336 B.n333 10.6151
R736 B.n331 B.n328 10.6151
R737 B.n328 B.n327 10.6151
R738 B.n327 B.n324 10.6151
R739 B.n324 B.n323 10.6151
R740 B.n323 B.n320 10.6151
R741 B.n320 B.n319 10.6151
R742 B.n319 B.n316 10.6151
R743 B.n316 B.n315 10.6151
R744 B.n315 B.n312 10.6151
R745 B.n312 B.n311 10.6151
R746 B.n311 B.n308 10.6151
R747 B.n308 B.n307 10.6151
R748 B.n307 B.n304 10.6151
R749 B.n304 B.n303 10.6151
R750 B.n303 B.n300 10.6151
R751 B.n300 B.n299 10.6151
R752 B.n299 B.n296 10.6151
R753 B.n296 B.n295 10.6151
R754 B.n295 B.n292 10.6151
R755 B.n292 B.n291 10.6151
R756 B.n291 B.n288 10.6151
R757 B.n288 B.n287 10.6151
R758 B.n287 B.n284 10.6151
R759 B.n284 B.n283 10.6151
R760 B.n283 B.n280 10.6151
R761 B.n280 B.n279 10.6151
R762 B.n279 B.n238 10.6151
R763 B.n411 B.n238 10.6151
R764 B.n413 B.n412 10.6151
R765 B.n413 B.n229 10.6151
R766 B.n423 B.n229 10.6151
R767 B.n424 B.n423 10.6151
R768 B.n425 B.n424 10.6151
R769 B.n425 B.n222 10.6151
R770 B.n435 B.n222 10.6151
R771 B.n436 B.n435 10.6151
R772 B.n437 B.n436 10.6151
R773 B.n437 B.n214 10.6151
R774 B.n447 B.n214 10.6151
R775 B.n448 B.n447 10.6151
R776 B.n450 B.n448 10.6151
R777 B.n450 B.n449 10.6151
R778 B.n449 B.n207 10.6151
R779 B.n462 B.n207 10.6151
R780 B.n463 B.n462 10.6151
R781 B.n464 B.n463 10.6151
R782 B.n465 B.n464 10.6151
R783 B.n466 B.n465 10.6151
R784 B.n469 B.n466 10.6151
R785 B.n470 B.n469 10.6151
R786 B.n471 B.n470 10.6151
R787 B.n472 B.n471 10.6151
R788 B.n474 B.n472 10.6151
R789 B.n475 B.n474 10.6151
R790 B.n476 B.n475 10.6151
R791 B.n477 B.n476 10.6151
R792 B.n479 B.n477 10.6151
R793 B.n480 B.n479 10.6151
R794 B.n481 B.n480 10.6151
R795 B.n482 B.n481 10.6151
R796 B.n484 B.n482 10.6151
R797 B.n485 B.n484 10.6151
R798 B.n486 B.n485 10.6151
R799 B.n519 B.n1 10.6151
R800 B.n519 B.n518 10.6151
R801 B.n518 B.n517 10.6151
R802 B.n517 B.n10 10.6151
R803 B.n511 B.n10 10.6151
R804 B.n511 B.n510 10.6151
R805 B.n510 B.n509 10.6151
R806 B.n509 B.n18 10.6151
R807 B.n503 B.n18 10.6151
R808 B.n503 B.n502 10.6151
R809 B.n502 B.n501 10.6151
R810 B.n501 B.n25 10.6151
R811 B.n495 B.n25 10.6151
R812 B.n495 B.n494 10.6151
R813 B.n494 B.n493 10.6151
R814 B.n493 B.n32 10.6151
R815 B.n77 B.n76 10.6151
R816 B.n80 B.n77 10.6151
R817 B.n81 B.n80 10.6151
R818 B.n84 B.n81 10.6151
R819 B.n85 B.n84 10.6151
R820 B.n88 B.n85 10.6151
R821 B.n89 B.n88 10.6151
R822 B.n92 B.n89 10.6151
R823 B.n93 B.n92 10.6151
R824 B.n96 B.n93 10.6151
R825 B.n97 B.n96 10.6151
R826 B.n100 B.n97 10.6151
R827 B.n101 B.n100 10.6151
R828 B.n104 B.n101 10.6151
R829 B.n105 B.n104 10.6151
R830 B.n108 B.n105 10.6151
R831 B.n109 B.n108 10.6151
R832 B.n112 B.n109 10.6151
R833 B.n113 B.n112 10.6151
R834 B.n116 B.n113 10.6151
R835 B.n117 B.n116 10.6151
R836 B.n120 B.n117 10.6151
R837 B.n121 B.n120 10.6151
R838 B.n124 B.n121 10.6151
R839 B.n125 B.n124 10.6151
R840 B.n128 B.n125 10.6151
R841 B.n129 B.n128 10.6151
R842 B.n132 B.n129 10.6151
R843 B.n137 B.n134 10.6151
R844 B.n138 B.n137 10.6151
R845 B.n141 B.n138 10.6151
R846 B.n142 B.n141 10.6151
R847 B.n145 B.n142 10.6151
R848 B.n146 B.n145 10.6151
R849 B.n149 B.n146 10.6151
R850 B.n150 B.n149 10.6151
R851 B.n154 B.n153 10.6151
R852 B.n157 B.n154 10.6151
R853 B.n158 B.n157 10.6151
R854 B.n161 B.n158 10.6151
R855 B.n162 B.n161 10.6151
R856 B.n165 B.n162 10.6151
R857 B.n166 B.n165 10.6151
R858 B.n169 B.n166 10.6151
R859 B.n170 B.n169 10.6151
R860 B.n173 B.n170 10.6151
R861 B.n174 B.n173 10.6151
R862 B.n177 B.n174 10.6151
R863 B.n178 B.n177 10.6151
R864 B.n181 B.n178 10.6151
R865 B.n182 B.n181 10.6151
R866 B.n185 B.n182 10.6151
R867 B.n186 B.n185 10.6151
R868 B.n189 B.n186 10.6151
R869 B.n190 B.n189 10.6151
R870 B.n193 B.n190 10.6151
R871 B.n194 B.n193 10.6151
R872 B.n197 B.n194 10.6151
R873 B.n198 B.n197 10.6151
R874 B.n201 B.n198 10.6151
R875 B.n202 B.n201 10.6151
R876 B.n205 B.n202 10.6151
R877 B.n206 B.n205 10.6151
R878 B.n487 B.n206 10.6151
R879 B.n527 B.n0 8.11757
R880 B.n527 B.n1 8.11757
R881 B.n445 B.t2 7.73186
R882 B.t3 B.n513 7.73186
R883 B.n349 B.n275 6.4005
R884 B.n333 B.n332 6.4005
R885 B.n134 B.n133 6.4005
R886 B.n150 B.n72 6.4005
R887 B.n352 B.n275 4.21513
R888 B.n332 B.n331 4.21513
R889 B.n133 B.n132 4.21513
R890 B.n153 B.n72 4.21513
R891 VP.n1 VP.t3 315.659
R892 VP.n1 VP.t0 315.61
R893 VP.n3 VP.t1 294.663
R894 VP.n5 VP.t2 294.663
R895 VP.n6 VP.n5 161.3
R896 VP.n4 VP.n0 161.3
R897 VP.n3 VP.n2 161.3
R898 VP.n2 VP.n1 81.8742
R899 VP.n4 VP.n3 24.1005
R900 VP.n5 VP.n4 24.1005
R901 VP.n2 VP.n0 0.189894
R902 VP.n6 VP.n0 0.189894
R903 VP VP.n6 0.0516364
R904 VTAIL.n5 VTAIL.t4 51.9874
R905 VTAIL.n4 VTAIL.t0 51.9874
R906 VTAIL.n3 VTAIL.t1 51.9874
R907 VTAIL.n7 VTAIL.t2 51.9872
R908 VTAIL.n0 VTAIL.t3 51.9872
R909 VTAIL.n1 VTAIL.t5 51.9872
R910 VTAIL.n2 VTAIL.t6 51.9872
R911 VTAIL.n6 VTAIL.t7 51.9872
R912 VTAIL.n7 VTAIL.n6 19.7893
R913 VTAIL.n3 VTAIL.n2 19.7893
R914 VTAIL.n4 VTAIL.n3 0.931535
R915 VTAIL.n6 VTAIL.n5 0.931535
R916 VTAIL.n2 VTAIL.n1 0.931535
R917 VTAIL VTAIL.n0 0.524207
R918 VTAIL.n5 VTAIL.n4 0.470328
R919 VTAIL.n1 VTAIL.n0 0.470328
R920 VTAIL VTAIL.n7 0.407828
R921 VDD1 VDD1.n1 99.5606
R922 VDD1 VDD1.n0 66.0947
R923 VDD1.n0 VDD1.t0 2.62998
R924 VDD1.n0 VDD1.t3 2.62998
R925 VDD1.n1 VDD1.t2 2.62998
R926 VDD1.n1 VDD1.t1 2.62998
R927 VN.n0 VN.t1 315.659
R928 VN.n1 VN.t0 315.659
R929 VN.n0 VN.t2 315.61
R930 VN.n1 VN.t3 315.61
R931 VN VN.n1 82.2549
R932 VN VN.n0 44.7132
R933 VDD2.n2 VDD2.n0 99.0358
R934 VDD2.n2 VDD2.n1 66.0365
R935 VDD2.n1 VDD2.t0 2.62998
R936 VDD2.n1 VDD2.t3 2.62998
R937 VDD2.n0 VDD2.t2 2.62998
R938 VDD2.n0 VDD2.t1 2.62998
R939 VDD2 VDD2.n2 0.0586897
C0 VDD1 VN 0.147136f
C1 VDD1 VP 2.28199f
C2 VDD2 VTAIL 4.75705f
C3 VN VTAIL 1.94918f
C4 VDD2 VN 2.153f
C5 VP VTAIL 1.96329f
C6 VDD2 VP 0.276396f
C7 VDD1 VTAIL 4.71524f
C8 VDD2 VDD1 0.577924f
C9 VP VN 4.03075f
C10 VDD2 B 2.378547f
C11 VDD1 B 5.4876f
C12 VTAIL B 6.282812f
C13 VN B 6.90346f
C14 VP B 4.700194f
C15 VDD2.t2 B 0.167537f
C16 VDD2.t1 B 0.167537f
C17 VDD2.n0 B 1.88176f
C18 VDD2.t0 B 0.167537f
C19 VDD2.t3 B 0.167537f
C20 VDD2.n1 B 1.44339f
C21 VDD2.n2 B 2.91417f
C22 VN.t1 B 0.620527f
C23 VN.t2 B 0.620479f
C24 VN.n0 B 0.49397f
C25 VN.t0 B 0.620527f
C26 VN.t3 B 0.620479f
C27 VN.n1 B 1.10888f
C28 VDD1.t0 B 0.165085f
C29 VDD1.t3 B 0.165085f
C30 VDD1.n0 B 1.42254f
C31 VDD1.t2 B 0.165085f
C32 VDD1.t1 B 0.165085f
C33 VDD1.n1 B 1.8779f
C34 VTAIL.t3 B 0.761497f
C35 VTAIL.n0 B 0.188531f
C36 VTAIL.t5 B 0.761497f
C37 VTAIL.n1 B 0.204675f
C38 VTAIL.t6 B 0.761497f
C39 VTAIL.n2 B 0.647331f
C40 VTAIL.t1 B 0.761499f
C41 VTAIL.n3 B 0.647329f
C42 VTAIL.t0 B 0.761499f
C43 VTAIL.n4 B 0.204673f
C44 VTAIL.t4 B 0.761499f
C45 VTAIL.n5 B 0.204673f
C46 VTAIL.t7 B 0.761497f
C47 VTAIL.n6 B 0.647331f
C48 VTAIL.t2 B 0.761497f
C49 VTAIL.n7 B 0.626574f
C50 VP.n0 B 0.038002f
C51 VP.t0 B 0.635833f
C52 VP.t3 B 0.635882f
C53 VP.n1 B 1.1214f
C54 VP.n2 B 2.04563f
C55 VP.t1 B 0.617965f
C56 VP.n3 B 0.266481f
C57 VP.n4 B 0.008623f
C58 VP.t2 B 0.617965f
C59 VP.n5 B 0.266481f
C60 VP.n6 B 0.02945f
.ends

