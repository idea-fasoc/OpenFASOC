* NGSPICE file created from diff_pair_sample_1772.ext - technology: sky130A

.subckt diff_pair_sample_1772 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t10 VN.t0 VDD2.t3 w_n4154_n1626# sky130_fd_pr__pfet_01v8 ad=0.54285 pd=3.62 as=0.54285 ps=3.62 w=3.29 l=3.65
X1 VTAIL.t0 VP.t0 VDD1.t5 w_n4154_n1626# sky130_fd_pr__pfet_01v8 ad=0.54285 pd=3.62 as=0.54285 ps=3.62 w=3.29 l=3.65
X2 B.t11 B.t9 B.t10 w_n4154_n1626# sky130_fd_pr__pfet_01v8 ad=1.2831 pd=7.36 as=0 ps=0 w=3.29 l=3.65
X3 VTAIL.t11 VP.t1 VDD1.t4 w_n4154_n1626# sky130_fd_pr__pfet_01v8 ad=0.54285 pd=3.62 as=0.54285 ps=3.62 w=3.29 l=3.65
X4 VDD2.t4 VN.t1 VTAIL.t9 w_n4154_n1626# sky130_fd_pr__pfet_01v8 ad=1.2831 pd=7.36 as=0.54285 ps=3.62 w=3.29 l=3.65
X5 VTAIL.t8 VN.t2 VDD2.t0 w_n4154_n1626# sky130_fd_pr__pfet_01v8 ad=0.54285 pd=3.62 as=0.54285 ps=3.62 w=3.29 l=3.65
X6 VDD2.t5 VN.t3 VTAIL.t7 w_n4154_n1626# sky130_fd_pr__pfet_01v8 ad=1.2831 pd=7.36 as=0.54285 ps=3.62 w=3.29 l=3.65
X7 VDD2.t2 VN.t4 VTAIL.t6 w_n4154_n1626# sky130_fd_pr__pfet_01v8 ad=0.54285 pd=3.62 as=1.2831 ps=7.36 w=3.29 l=3.65
X8 VDD2.t1 VN.t5 VTAIL.t5 w_n4154_n1626# sky130_fd_pr__pfet_01v8 ad=0.54285 pd=3.62 as=1.2831 ps=7.36 w=3.29 l=3.65
X9 VDD1.t3 VP.t2 VTAIL.t1 w_n4154_n1626# sky130_fd_pr__pfet_01v8 ad=0.54285 pd=3.62 as=1.2831 ps=7.36 w=3.29 l=3.65
X10 VDD1.t2 VP.t3 VTAIL.t2 w_n4154_n1626# sky130_fd_pr__pfet_01v8 ad=1.2831 pd=7.36 as=0.54285 ps=3.62 w=3.29 l=3.65
X11 VDD1.t1 VP.t4 VTAIL.t4 w_n4154_n1626# sky130_fd_pr__pfet_01v8 ad=1.2831 pd=7.36 as=0.54285 ps=3.62 w=3.29 l=3.65
X12 B.t8 B.t6 B.t7 w_n4154_n1626# sky130_fd_pr__pfet_01v8 ad=1.2831 pd=7.36 as=0 ps=0 w=3.29 l=3.65
X13 B.t5 B.t3 B.t4 w_n4154_n1626# sky130_fd_pr__pfet_01v8 ad=1.2831 pd=7.36 as=0 ps=0 w=3.29 l=3.65
X14 VDD1.t0 VP.t5 VTAIL.t3 w_n4154_n1626# sky130_fd_pr__pfet_01v8 ad=0.54285 pd=3.62 as=1.2831 ps=7.36 w=3.29 l=3.65
X15 B.t2 B.t0 B.t1 w_n4154_n1626# sky130_fd_pr__pfet_01v8 ad=1.2831 pd=7.36 as=0 ps=0 w=3.29 l=3.65
R0 VN.n38 VN.n37 161.3
R1 VN.n36 VN.n21 161.3
R2 VN.n35 VN.n34 161.3
R3 VN.n33 VN.n22 161.3
R4 VN.n32 VN.n31 161.3
R5 VN.n30 VN.n23 161.3
R6 VN.n29 VN.n28 161.3
R7 VN.n27 VN.n24 161.3
R8 VN.n18 VN.n17 161.3
R9 VN.n16 VN.n1 161.3
R10 VN.n15 VN.n14 161.3
R11 VN.n13 VN.n2 161.3
R12 VN.n12 VN.n11 161.3
R13 VN.n10 VN.n3 161.3
R14 VN.n9 VN.n8 161.3
R15 VN.n7 VN.n4 161.3
R16 VN.n19 VN.n0 78.8126
R17 VN.n39 VN.n20 78.8126
R18 VN.n26 VN.n25 62.412
R19 VN.n6 VN.n5 62.412
R20 VN.n11 VN.n2 56.5193
R21 VN.n31 VN.n22 56.5193
R22 VN.n26 VN.t5 55.3043
R23 VN.n6 VN.t1 55.3043
R24 VN VN.n39 46.5056
R25 VN.n9 VN.n4 24.4675
R26 VN.n10 VN.n9 24.4675
R27 VN.n11 VN.n10 24.4675
R28 VN.n15 VN.n2 24.4675
R29 VN.n16 VN.n15 24.4675
R30 VN.n17 VN.n16 24.4675
R31 VN.n31 VN.n30 24.4675
R32 VN.n30 VN.n29 24.4675
R33 VN.n29 VN.n24 24.4675
R34 VN.n37 VN.n36 24.4675
R35 VN.n36 VN.n35 24.4675
R36 VN.n35 VN.n22 24.4675
R37 VN.n5 VN.t0 21.7235
R38 VN.n0 VN.t4 21.7235
R39 VN.n25 VN.t2 21.7235
R40 VN.n20 VN.t3 21.7235
R41 VN.n5 VN.n4 12.234
R42 VN.n25 VN.n24 12.234
R43 VN.n17 VN.n0 11.2553
R44 VN.n37 VN.n20 11.2553
R45 VN.n27 VN.n26 3.1161
R46 VN.n7 VN.n6 3.1161
R47 VN.n39 VN.n38 0.354971
R48 VN.n19 VN.n18 0.354971
R49 VN VN.n19 0.26696
R50 VN.n38 VN.n21 0.189894
R51 VN.n34 VN.n21 0.189894
R52 VN.n34 VN.n33 0.189894
R53 VN.n33 VN.n32 0.189894
R54 VN.n32 VN.n23 0.189894
R55 VN.n28 VN.n23 0.189894
R56 VN.n28 VN.n27 0.189894
R57 VN.n8 VN.n7 0.189894
R58 VN.n8 VN.n3 0.189894
R59 VN.n12 VN.n3 0.189894
R60 VN.n13 VN.n12 0.189894
R61 VN.n14 VN.n13 0.189894
R62 VN.n14 VN.n1 0.189894
R63 VN.n18 VN.n1 0.189894
R64 VDD2.n27 VDD2.n17 756.745
R65 VDD2.n10 VDD2.n0 756.745
R66 VDD2.n28 VDD2.n27 585
R67 VDD2.n26 VDD2.n25 585
R68 VDD2.n21 VDD2.n20 585
R69 VDD2.n4 VDD2.n3 585
R70 VDD2.n9 VDD2.n8 585
R71 VDD2.n11 VDD2.n10 585
R72 VDD2.n22 VDD2.t5 336.901
R73 VDD2.n5 VDD2.t4 336.901
R74 VDD2.n27 VDD2.n26 171.744
R75 VDD2.n26 VDD2.n20 171.744
R76 VDD2.n9 VDD2.n3 171.744
R77 VDD2.n10 VDD2.n9 171.744
R78 VDD2.n16 VDD2.n15 131.951
R79 VDD2 VDD2.n33 131.947
R80 VDD2.t5 VDD2.n20 85.8723
R81 VDD2.t4 VDD2.n3 85.8723
R82 VDD2.n16 VDD2.n14 54.679
R83 VDD2.n32 VDD2.n31 52.1611
R84 VDD2.n32 VDD2.n16 37.7024
R85 VDD2.n22 VDD2.n21 16.193
R86 VDD2.n5 VDD2.n4 16.193
R87 VDD2.n25 VDD2.n24 12.8005
R88 VDD2.n8 VDD2.n7 12.8005
R89 VDD2.n28 VDD2.n19 12.0247
R90 VDD2.n11 VDD2.n2 12.0247
R91 VDD2.n29 VDD2.n17 11.249
R92 VDD2.n12 VDD2.n0 11.249
R93 VDD2.n33 VDD2.t0 9.88044
R94 VDD2.n33 VDD2.t1 9.88044
R95 VDD2.n15 VDD2.t3 9.88044
R96 VDD2.n15 VDD2.t2 9.88044
R97 VDD2.n31 VDD2.n30 9.45567
R98 VDD2.n14 VDD2.n13 9.45567
R99 VDD2.n30 VDD2.n29 9.3005
R100 VDD2.n19 VDD2.n18 9.3005
R101 VDD2.n24 VDD2.n23 9.3005
R102 VDD2.n13 VDD2.n12 9.3005
R103 VDD2.n2 VDD2.n1 9.3005
R104 VDD2.n7 VDD2.n6 9.3005
R105 VDD2.n23 VDD2.n22 3.91276
R106 VDD2.n6 VDD2.n5 3.91276
R107 VDD2.n31 VDD2.n17 2.71565
R108 VDD2.n14 VDD2.n0 2.71565
R109 VDD2 VDD2.n32 2.63197
R110 VDD2.n29 VDD2.n28 1.93989
R111 VDD2.n12 VDD2.n11 1.93989
R112 VDD2.n25 VDD2.n19 1.16414
R113 VDD2.n8 VDD2.n2 1.16414
R114 VDD2.n24 VDD2.n21 0.388379
R115 VDD2.n7 VDD2.n4 0.388379
R116 VDD2.n30 VDD2.n18 0.155672
R117 VDD2.n23 VDD2.n18 0.155672
R118 VDD2.n6 VDD2.n1 0.155672
R119 VDD2.n13 VDD2.n1 0.155672
R120 VTAIL.n66 VTAIL.n56 756.745
R121 VTAIL.n12 VTAIL.n2 756.745
R122 VTAIL.n50 VTAIL.n40 756.745
R123 VTAIL.n32 VTAIL.n22 756.745
R124 VTAIL.n60 VTAIL.n59 585
R125 VTAIL.n65 VTAIL.n64 585
R126 VTAIL.n67 VTAIL.n66 585
R127 VTAIL.n6 VTAIL.n5 585
R128 VTAIL.n11 VTAIL.n10 585
R129 VTAIL.n13 VTAIL.n12 585
R130 VTAIL.n51 VTAIL.n50 585
R131 VTAIL.n49 VTAIL.n48 585
R132 VTAIL.n44 VTAIL.n43 585
R133 VTAIL.n33 VTAIL.n32 585
R134 VTAIL.n31 VTAIL.n30 585
R135 VTAIL.n26 VTAIL.n25 585
R136 VTAIL.n61 VTAIL.t6 336.901
R137 VTAIL.n7 VTAIL.t1 336.901
R138 VTAIL.n45 VTAIL.t3 336.901
R139 VTAIL.n27 VTAIL.t5 336.901
R140 VTAIL.n65 VTAIL.n59 171.744
R141 VTAIL.n66 VTAIL.n65 171.744
R142 VTAIL.n11 VTAIL.n5 171.744
R143 VTAIL.n12 VTAIL.n11 171.744
R144 VTAIL.n50 VTAIL.n49 171.744
R145 VTAIL.n49 VTAIL.n43 171.744
R146 VTAIL.n32 VTAIL.n31 171.744
R147 VTAIL.n31 VTAIL.n25 171.744
R148 VTAIL.n39 VTAIL.n38 114.469
R149 VTAIL.n21 VTAIL.n20 114.469
R150 VTAIL.n1 VTAIL.n0 114.469
R151 VTAIL.n19 VTAIL.n18 114.469
R152 VTAIL.t6 VTAIL.n59 85.8723
R153 VTAIL.t1 VTAIL.n5 85.8723
R154 VTAIL.t3 VTAIL.n43 85.8723
R155 VTAIL.t5 VTAIL.n25 85.8723
R156 VTAIL.n71 VTAIL.n70 35.4823
R157 VTAIL.n17 VTAIL.n16 35.4823
R158 VTAIL.n55 VTAIL.n54 35.4823
R159 VTAIL.n37 VTAIL.n36 35.4823
R160 VTAIL.n21 VTAIL.n19 22.0652
R161 VTAIL.n71 VTAIL.n55 18.6341
R162 VTAIL.n61 VTAIL.n60 16.193
R163 VTAIL.n7 VTAIL.n6 16.193
R164 VTAIL.n45 VTAIL.n44 16.193
R165 VTAIL.n27 VTAIL.n26 16.193
R166 VTAIL.n64 VTAIL.n63 12.8005
R167 VTAIL.n10 VTAIL.n9 12.8005
R168 VTAIL.n48 VTAIL.n47 12.8005
R169 VTAIL.n30 VTAIL.n29 12.8005
R170 VTAIL.n67 VTAIL.n58 12.0247
R171 VTAIL.n13 VTAIL.n4 12.0247
R172 VTAIL.n51 VTAIL.n42 12.0247
R173 VTAIL.n33 VTAIL.n24 12.0247
R174 VTAIL.n68 VTAIL.n56 11.249
R175 VTAIL.n14 VTAIL.n2 11.249
R176 VTAIL.n52 VTAIL.n40 11.249
R177 VTAIL.n34 VTAIL.n22 11.249
R178 VTAIL.n0 VTAIL.t9 9.88044
R179 VTAIL.n0 VTAIL.t10 9.88044
R180 VTAIL.n18 VTAIL.t2 9.88044
R181 VTAIL.n18 VTAIL.t0 9.88044
R182 VTAIL.n38 VTAIL.t4 9.88044
R183 VTAIL.n38 VTAIL.t11 9.88044
R184 VTAIL.n20 VTAIL.t7 9.88044
R185 VTAIL.n20 VTAIL.t8 9.88044
R186 VTAIL.n70 VTAIL.n69 9.45567
R187 VTAIL.n16 VTAIL.n15 9.45567
R188 VTAIL.n54 VTAIL.n53 9.45567
R189 VTAIL.n36 VTAIL.n35 9.45567
R190 VTAIL.n69 VTAIL.n68 9.3005
R191 VTAIL.n58 VTAIL.n57 9.3005
R192 VTAIL.n63 VTAIL.n62 9.3005
R193 VTAIL.n15 VTAIL.n14 9.3005
R194 VTAIL.n4 VTAIL.n3 9.3005
R195 VTAIL.n9 VTAIL.n8 9.3005
R196 VTAIL.n53 VTAIL.n52 9.3005
R197 VTAIL.n42 VTAIL.n41 9.3005
R198 VTAIL.n47 VTAIL.n46 9.3005
R199 VTAIL.n35 VTAIL.n34 9.3005
R200 VTAIL.n24 VTAIL.n23 9.3005
R201 VTAIL.n29 VTAIL.n28 9.3005
R202 VTAIL.n46 VTAIL.n45 3.91276
R203 VTAIL.n28 VTAIL.n27 3.91276
R204 VTAIL.n62 VTAIL.n61 3.91276
R205 VTAIL.n8 VTAIL.n7 3.91276
R206 VTAIL.n37 VTAIL.n21 3.43153
R207 VTAIL.n55 VTAIL.n39 3.43153
R208 VTAIL.n19 VTAIL.n17 3.43153
R209 VTAIL.n70 VTAIL.n56 2.71565
R210 VTAIL.n16 VTAIL.n2 2.71565
R211 VTAIL.n54 VTAIL.n40 2.71565
R212 VTAIL.n36 VTAIL.n22 2.71565
R213 VTAIL VTAIL.n71 2.51559
R214 VTAIL.n39 VTAIL.n37 2.18584
R215 VTAIL.n17 VTAIL.n1 2.18584
R216 VTAIL.n68 VTAIL.n67 1.93989
R217 VTAIL.n14 VTAIL.n13 1.93989
R218 VTAIL.n52 VTAIL.n51 1.93989
R219 VTAIL.n34 VTAIL.n33 1.93989
R220 VTAIL.n64 VTAIL.n58 1.16414
R221 VTAIL.n10 VTAIL.n4 1.16414
R222 VTAIL.n48 VTAIL.n42 1.16414
R223 VTAIL.n30 VTAIL.n24 1.16414
R224 VTAIL VTAIL.n1 0.916448
R225 VTAIL.n63 VTAIL.n60 0.388379
R226 VTAIL.n9 VTAIL.n6 0.388379
R227 VTAIL.n47 VTAIL.n44 0.388379
R228 VTAIL.n29 VTAIL.n26 0.388379
R229 VTAIL.n62 VTAIL.n57 0.155672
R230 VTAIL.n69 VTAIL.n57 0.155672
R231 VTAIL.n8 VTAIL.n3 0.155672
R232 VTAIL.n15 VTAIL.n3 0.155672
R233 VTAIL.n53 VTAIL.n41 0.155672
R234 VTAIL.n46 VTAIL.n41 0.155672
R235 VTAIL.n35 VTAIL.n23 0.155672
R236 VTAIL.n28 VTAIL.n23 0.155672
R237 VP.n16 VP.n13 161.3
R238 VP.n18 VP.n17 161.3
R239 VP.n19 VP.n12 161.3
R240 VP.n21 VP.n20 161.3
R241 VP.n22 VP.n11 161.3
R242 VP.n24 VP.n23 161.3
R243 VP.n25 VP.n10 161.3
R244 VP.n27 VP.n26 161.3
R245 VP.n55 VP.n54 161.3
R246 VP.n53 VP.n1 161.3
R247 VP.n52 VP.n51 161.3
R248 VP.n50 VP.n2 161.3
R249 VP.n49 VP.n48 161.3
R250 VP.n47 VP.n3 161.3
R251 VP.n46 VP.n45 161.3
R252 VP.n44 VP.n4 161.3
R253 VP.n43 VP.n42 161.3
R254 VP.n40 VP.n5 161.3
R255 VP.n39 VP.n38 161.3
R256 VP.n37 VP.n6 161.3
R257 VP.n36 VP.n35 161.3
R258 VP.n34 VP.n7 161.3
R259 VP.n33 VP.n32 161.3
R260 VP.n31 VP.n8 161.3
R261 VP.n30 VP.n29 78.8126
R262 VP.n56 VP.n0 78.8126
R263 VP.n28 VP.n9 78.8126
R264 VP.n15 VP.n14 62.412
R265 VP.n35 VP.n6 56.5193
R266 VP.n48 VP.n2 56.5193
R267 VP.n20 VP.n11 56.5193
R268 VP.n15 VP.t4 55.3041
R269 VP.n30 VP.n28 46.3402
R270 VP.n33 VP.n8 24.4675
R271 VP.n34 VP.n33 24.4675
R272 VP.n35 VP.n34 24.4675
R273 VP.n39 VP.n6 24.4675
R274 VP.n40 VP.n39 24.4675
R275 VP.n42 VP.n40 24.4675
R276 VP.n46 VP.n4 24.4675
R277 VP.n47 VP.n46 24.4675
R278 VP.n48 VP.n47 24.4675
R279 VP.n52 VP.n2 24.4675
R280 VP.n53 VP.n52 24.4675
R281 VP.n54 VP.n53 24.4675
R282 VP.n24 VP.n11 24.4675
R283 VP.n25 VP.n24 24.4675
R284 VP.n26 VP.n25 24.4675
R285 VP.n18 VP.n13 24.4675
R286 VP.n19 VP.n18 24.4675
R287 VP.n20 VP.n19 24.4675
R288 VP.n29 VP.t3 21.7235
R289 VP.n41 VP.t0 21.7235
R290 VP.n0 VP.t2 21.7235
R291 VP.n9 VP.t5 21.7235
R292 VP.n14 VP.t1 21.7235
R293 VP.n42 VP.n41 12.234
R294 VP.n41 VP.n4 12.234
R295 VP.n14 VP.n13 12.234
R296 VP.n29 VP.n8 11.2553
R297 VP.n54 VP.n0 11.2553
R298 VP.n26 VP.n9 11.2553
R299 VP.n16 VP.n15 3.11608
R300 VP.n28 VP.n27 0.354971
R301 VP.n31 VP.n30 0.354971
R302 VP.n56 VP.n55 0.354971
R303 VP VP.n56 0.26696
R304 VP.n17 VP.n16 0.189894
R305 VP.n17 VP.n12 0.189894
R306 VP.n21 VP.n12 0.189894
R307 VP.n22 VP.n21 0.189894
R308 VP.n23 VP.n22 0.189894
R309 VP.n23 VP.n10 0.189894
R310 VP.n27 VP.n10 0.189894
R311 VP.n32 VP.n31 0.189894
R312 VP.n32 VP.n7 0.189894
R313 VP.n36 VP.n7 0.189894
R314 VP.n37 VP.n36 0.189894
R315 VP.n38 VP.n37 0.189894
R316 VP.n38 VP.n5 0.189894
R317 VP.n43 VP.n5 0.189894
R318 VP.n44 VP.n43 0.189894
R319 VP.n45 VP.n44 0.189894
R320 VP.n45 VP.n3 0.189894
R321 VP.n49 VP.n3 0.189894
R322 VP.n50 VP.n49 0.189894
R323 VP.n51 VP.n50 0.189894
R324 VP.n51 VP.n1 0.189894
R325 VP.n55 VP.n1 0.189894
R326 VDD1.n10 VDD1.n0 756.745
R327 VDD1.n25 VDD1.n15 756.745
R328 VDD1.n11 VDD1.n10 585
R329 VDD1.n9 VDD1.n8 585
R330 VDD1.n4 VDD1.n3 585
R331 VDD1.n19 VDD1.n18 585
R332 VDD1.n24 VDD1.n23 585
R333 VDD1.n26 VDD1.n25 585
R334 VDD1.n5 VDD1.t1 336.901
R335 VDD1.n20 VDD1.t2 336.901
R336 VDD1.n10 VDD1.n9 171.744
R337 VDD1.n9 VDD1.n3 171.744
R338 VDD1.n24 VDD1.n18 171.744
R339 VDD1.n25 VDD1.n24 171.744
R340 VDD1.n31 VDD1.n30 131.951
R341 VDD1.n33 VDD1.n32 131.148
R342 VDD1.t1 VDD1.n3 85.8723
R343 VDD1.t2 VDD1.n18 85.8723
R344 VDD1 VDD1.n14 54.7926
R345 VDD1.n31 VDD1.n29 54.679
R346 VDD1.n33 VDD1.n31 40.0009
R347 VDD1.n5 VDD1.n4 16.193
R348 VDD1.n20 VDD1.n19 16.193
R349 VDD1.n8 VDD1.n7 12.8005
R350 VDD1.n23 VDD1.n22 12.8005
R351 VDD1.n11 VDD1.n2 12.0247
R352 VDD1.n26 VDD1.n17 12.0247
R353 VDD1.n12 VDD1.n0 11.249
R354 VDD1.n27 VDD1.n15 11.249
R355 VDD1.n32 VDD1.t4 9.88044
R356 VDD1.n32 VDD1.t0 9.88044
R357 VDD1.n30 VDD1.t5 9.88044
R358 VDD1.n30 VDD1.t3 9.88044
R359 VDD1.n14 VDD1.n13 9.45567
R360 VDD1.n29 VDD1.n28 9.45567
R361 VDD1.n13 VDD1.n12 9.3005
R362 VDD1.n2 VDD1.n1 9.3005
R363 VDD1.n7 VDD1.n6 9.3005
R364 VDD1.n28 VDD1.n27 9.3005
R365 VDD1.n17 VDD1.n16 9.3005
R366 VDD1.n22 VDD1.n21 9.3005
R367 VDD1.n6 VDD1.n5 3.91276
R368 VDD1.n21 VDD1.n20 3.91276
R369 VDD1.n14 VDD1.n0 2.71565
R370 VDD1.n29 VDD1.n15 2.71565
R371 VDD1.n12 VDD1.n11 1.93989
R372 VDD1.n27 VDD1.n26 1.93989
R373 VDD1.n8 VDD1.n2 1.16414
R374 VDD1.n23 VDD1.n17 1.16414
R375 VDD1 VDD1.n33 0.800069
R376 VDD1.n7 VDD1.n4 0.388379
R377 VDD1.n22 VDD1.n19 0.388379
R378 VDD1.n13 VDD1.n1 0.155672
R379 VDD1.n6 VDD1.n1 0.155672
R380 VDD1.n21 VDD1.n16 0.155672
R381 VDD1.n28 VDD1.n16 0.155672
R382 B.n476 B.n55 585
R383 B.n478 B.n477 585
R384 B.n479 B.n54 585
R385 B.n481 B.n480 585
R386 B.n482 B.n53 585
R387 B.n484 B.n483 585
R388 B.n485 B.n52 585
R389 B.n487 B.n486 585
R390 B.n488 B.n51 585
R391 B.n490 B.n489 585
R392 B.n491 B.n50 585
R393 B.n493 B.n492 585
R394 B.n494 B.n49 585
R395 B.n496 B.n495 585
R396 B.n497 B.n45 585
R397 B.n499 B.n498 585
R398 B.n500 B.n44 585
R399 B.n502 B.n501 585
R400 B.n503 B.n43 585
R401 B.n505 B.n504 585
R402 B.n506 B.n42 585
R403 B.n508 B.n507 585
R404 B.n509 B.n41 585
R405 B.n511 B.n510 585
R406 B.n512 B.n40 585
R407 B.n514 B.n513 585
R408 B.n516 B.n37 585
R409 B.n518 B.n517 585
R410 B.n519 B.n36 585
R411 B.n521 B.n520 585
R412 B.n522 B.n35 585
R413 B.n524 B.n523 585
R414 B.n525 B.n34 585
R415 B.n527 B.n526 585
R416 B.n528 B.n33 585
R417 B.n530 B.n529 585
R418 B.n531 B.n32 585
R419 B.n533 B.n532 585
R420 B.n534 B.n31 585
R421 B.n536 B.n535 585
R422 B.n537 B.n30 585
R423 B.n539 B.n538 585
R424 B.n475 B.n474 585
R425 B.n473 B.n56 585
R426 B.n472 B.n471 585
R427 B.n470 B.n57 585
R428 B.n469 B.n468 585
R429 B.n467 B.n58 585
R430 B.n466 B.n465 585
R431 B.n464 B.n59 585
R432 B.n463 B.n462 585
R433 B.n461 B.n60 585
R434 B.n460 B.n459 585
R435 B.n458 B.n61 585
R436 B.n457 B.n456 585
R437 B.n455 B.n62 585
R438 B.n454 B.n453 585
R439 B.n452 B.n63 585
R440 B.n451 B.n450 585
R441 B.n449 B.n64 585
R442 B.n448 B.n447 585
R443 B.n446 B.n65 585
R444 B.n445 B.n444 585
R445 B.n443 B.n66 585
R446 B.n442 B.n441 585
R447 B.n440 B.n67 585
R448 B.n439 B.n438 585
R449 B.n437 B.n68 585
R450 B.n436 B.n435 585
R451 B.n434 B.n69 585
R452 B.n433 B.n432 585
R453 B.n431 B.n70 585
R454 B.n430 B.n429 585
R455 B.n428 B.n71 585
R456 B.n427 B.n426 585
R457 B.n425 B.n72 585
R458 B.n424 B.n423 585
R459 B.n422 B.n73 585
R460 B.n421 B.n420 585
R461 B.n419 B.n74 585
R462 B.n418 B.n417 585
R463 B.n416 B.n75 585
R464 B.n415 B.n414 585
R465 B.n413 B.n76 585
R466 B.n412 B.n411 585
R467 B.n410 B.n77 585
R468 B.n409 B.n408 585
R469 B.n407 B.n78 585
R470 B.n406 B.n405 585
R471 B.n404 B.n79 585
R472 B.n403 B.n402 585
R473 B.n401 B.n80 585
R474 B.n400 B.n399 585
R475 B.n398 B.n81 585
R476 B.n397 B.n396 585
R477 B.n395 B.n82 585
R478 B.n394 B.n393 585
R479 B.n392 B.n83 585
R480 B.n391 B.n390 585
R481 B.n389 B.n84 585
R482 B.n388 B.n387 585
R483 B.n386 B.n85 585
R484 B.n385 B.n384 585
R485 B.n383 B.n86 585
R486 B.n382 B.n381 585
R487 B.n380 B.n87 585
R488 B.n379 B.n378 585
R489 B.n377 B.n88 585
R490 B.n376 B.n375 585
R491 B.n374 B.n89 585
R492 B.n373 B.n372 585
R493 B.n371 B.n90 585
R494 B.n370 B.n369 585
R495 B.n368 B.n91 585
R496 B.n367 B.n366 585
R497 B.n365 B.n92 585
R498 B.n364 B.n363 585
R499 B.n362 B.n93 585
R500 B.n361 B.n360 585
R501 B.n359 B.n94 585
R502 B.n358 B.n357 585
R503 B.n356 B.n95 585
R504 B.n355 B.n354 585
R505 B.n353 B.n96 585
R506 B.n352 B.n351 585
R507 B.n350 B.n97 585
R508 B.n349 B.n348 585
R509 B.n347 B.n98 585
R510 B.n346 B.n345 585
R511 B.n344 B.n99 585
R512 B.n343 B.n342 585
R513 B.n341 B.n100 585
R514 B.n340 B.n339 585
R515 B.n338 B.n101 585
R516 B.n337 B.n336 585
R517 B.n335 B.n102 585
R518 B.n334 B.n333 585
R519 B.n332 B.n103 585
R520 B.n331 B.n330 585
R521 B.n329 B.n104 585
R522 B.n328 B.n327 585
R523 B.n326 B.n105 585
R524 B.n325 B.n324 585
R525 B.n323 B.n106 585
R526 B.n322 B.n321 585
R527 B.n320 B.n107 585
R528 B.n319 B.n318 585
R529 B.n317 B.n108 585
R530 B.n316 B.n315 585
R531 B.n314 B.n109 585
R532 B.n313 B.n312 585
R533 B.n311 B.n110 585
R534 B.n310 B.n309 585
R535 B.n245 B.n136 585
R536 B.n247 B.n246 585
R537 B.n248 B.n135 585
R538 B.n250 B.n249 585
R539 B.n251 B.n134 585
R540 B.n253 B.n252 585
R541 B.n254 B.n133 585
R542 B.n256 B.n255 585
R543 B.n257 B.n132 585
R544 B.n259 B.n258 585
R545 B.n260 B.n131 585
R546 B.n262 B.n261 585
R547 B.n263 B.n130 585
R548 B.n265 B.n264 585
R549 B.n266 B.n129 585
R550 B.n268 B.n267 585
R551 B.n270 B.n126 585
R552 B.n272 B.n271 585
R553 B.n273 B.n125 585
R554 B.n275 B.n274 585
R555 B.n276 B.n124 585
R556 B.n278 B.n277 585
R557 B.n279 B.n123 585
R558 B.n281 B.n280 585
R559 B.n282 B.n122 585
R560 B.n284 B.n283 585
R561 B.n286 B.n285 585
R562 B.n287 B.n118 585
R563 B.n289 B.n288 585
R564 B.n290 B.n117 585
R565 B.n292 B.n291 585
R566 B.n293 B.n116 585
R567 B.n295 B.n294 585
R568 B.n296 B.n115 585
R569 B.n298 B.n297 585
R570 B.n299 B.n114 585
R571 B.n301 B.n300 585
R572 B.n302 B.n113 585
R573 B.n304 B.n303 585
R574 B.n305 B.n112 585
R575 B.n307 B.n306 585
R576 B.n308 B.n111 585
R577 B.n244 B.n243 585
R578 B.n242 B.n137 585
R579 B.n241 B.n240 585
R580 B.n239 B.n138 585
R581 B.n238 B.n237 585
R582 B.n236 B.n139 585
R583 B.n235 B.n234 585
R584 B.n233 B.n140 585
R585 B.n232 B.n231 585
R586 B.n230 B.n141 585
R587 B.n229 B.n228 585
R588 B.n227 B.n142 585
R589 B.n226 B.n225 585
R590 B.n224 B.n143 585
R591 B.n223 B.n222 585
R592 B.n221 B.n144 585
R593 B.n220 B.n219 585
R594 B.n218 B.n145 585
R595 B.n217 B.n216 585
R596 B.n215 B.n146 585
R597 B.n214 B.n213 585
R598 B.n212 B.n147 585
R599 B.n211 B.n210 585
R600 B.n209 B.n148 585
R601 B.n208 B.n207 585
R602 B.n206 B.n149 585
R603 B.n205 B.n204 585
R604 B.n203 B.n150 585
R605 B.n202 B.n201 585
R606 B.n200 B.n151 585
R607 B.n199 B.n198 585
R608 B.n197 B.n152 585
R609 B.n196 B.n195 585
R610 B.n194 B.n153 585
R611 B.n193 B.n192 585
R612 B.n191 B.n154 585
R613 B.n190 B.n189 585
R614 B.n188 B.n155 585
R615 B.n187 B.n186 585
R616 B.n185 B.n156 585
R617 B.n184 B.n183 585
R618 B.n182 B.n157 585
R619 B.n181 B.n180 585
R620 B.n179 B.n158 585
R621 B.n178 B.n177 585
R622 B.n176 B.n159 585
R623 B.n175 B.n174 585
R624 B.n173 B.n160 585
R625 B.n172 B.n171 585
R626 B.n170 B.n161 585
R627 B.n169 B.n168 585
R628 B.n167 B.n162 585
R629 B.n166 B.n165 585
R630 B.n164 B.n163 585
R631 B.n2 B.n0 585
R632 B.n621 B.n1 585
R633 B.n620 B.n619 585
R634 B.n618 B.n3 585
R635 B.n617 B.n616 585
R636 B.n615 B.n4 585
R637 B.n614 B.n613 585
R638 B.n612 B.n5 585
R639 B.n611 B.n610 585
R640 B.n609 B.n6 585
R641 B.n608 B.n607 585
R642 B.n606 B.n7 585
R643 B.n605 B.n604 585
R644 B.n603 B.n8 585
R645 B.n602 B.n601 585
R646 B.n600 B.n9 585
R647 B.n599 B.n598 585
R648 B.n597 B.n10 585
R649 B.n596 B.n595 585
R650 B.n594 B.n11 585
R651 B.n593 B.n592 585
R652 B.n591 B.n12 585
R653 B.n590 B.n589 585
R654 B.n588 B.n13 585
R655 B.n587 B.n586 585
R656 B.n585 B.n14 585
R657 B.n584 B.n583 585
R658 B.n582 B.n15 585
R659 B.n581 B.n580 585
R660 B.n579 B.n16 585
R661 B.n578 B.n577 585
R662 B.n576 B.n17 585
R663 B.n575 B.n574 585
R664 B.n573 B.n18 585
R665 B.n572 B.n571 585
R666 B.n570 B.n19 585
R667 B.n569 B.n568 585
R668 B.n567 B.n20 585
R669 B.n566 B.n565 585
R670 B.n564 B.n21 585
R671 B.n563 B.n562 585
R672 B.n561 B.n22 585
R673 B.n560 B.n559 585
R674 B.n558 B.n23 585
R675 B.n557 B.n556 585
R676 B.n555 B.n24 585
R677 B.n554 B.n553 585
R678 B.n552 B.n25 585
R679 B.n551 B.n550 585
R680 B.n549 B.n26 585
R681 B.n548 B.n547 585
R682 B.n546 B.n27 585
R683 B.n545 B.n544 585
R684 B.n543 B.n28 585
R685 B.n542 B.n541 585
R686 B.n540 B.n29 585
R687 B.n623 B.n622 585
R688 B.n243 B.n136 454.062
R689 B.n538 B.n29 454.062
R690 B.n309 B.n308 454.062
R691 B.n476 B.n475 454.062
R692 B.n119 B.t2 304.495
R693 B.n46 B.t4 304.495
R694 B.n127 B.t8 304.495
R695 B.n38 B.t10 304.495
R696 B.n119 B.t0 230.946
R697 B.n127 B.t6 230.946
R698 B.n38 B.t9 230.946
R699 B.n46 B.t3 230.946
R700 B.n120 B.t1 227.306
R701 B.n47 B.t5 227.306
R702 B.n128 B.t7 227.306
R703 B.n39 B.t11 227.306
R704 B.n243 B.n242 163.367
R705 B.n242 B.n241 163.367
R706 B.n241 B.n138 163.367
R707 B.n237 B.n138 163.367
R708 B.n237 B.n236 163.367
R709 B.n236 B.n235 163.367
R710 B.n235 B.n140 163.367
R711 B.n231 B.n140 163.367
R712 B.n231 B.n230 163.367
R713 B.n230 B.n229 163.367
R714 B.n229 B.n142 163.367
R715 B.n225 B.n142 163.367
R716 B.n225 B.n224 163.367
R717 B.n224 B.n223 163.367
R718 B.n223 B.n144 163.367
R719 B.n219 B.n144 163.367
R720 B.n219 B.n218 163.367
R721 B.n218 B.n217 163.367
R722 B.n217 B.n146 163.367
R723 B.n213 B.n146 163.367
R724 B.n213 B.n212 163.367
R725 B.n212 B.n211 163.367
R726 B.n211 B.n148 163.367
R727 B.n207 B.n148 163.367
R728 B.n207 B.n206 163.367
R729 B.n206 B.n205 163.367
R730 B.n205 B.n150 163.367
R731 B.n201 B.n150 163.367
R732 B.n201 B.n200 163.367
R733 B.n200 B.n199 163.367
R734 B.n199 B.n152 163.367
R735 B.n195 B.n152 163.367
R736 B.n195 B.n194 163.367
R737 B.n194 B.n193 163.367
R738 B.n193 B.n154 163.367
R739 B.n189 B.n154 163.367
R740 B.n189 B.n188 163.367
R741 B.n188 B.n187 163.367
R742 B.n187 B.n156 163.367
R743 B.n183 B.n156 163.367
R744 B.n183 B.n182 163.367
R745 B.n182 B.n181 163.367
R746 B.n181 B.n158 163.367
R747 B.n177 B.n158 163.367
R748 B.n177 B.n176 163.367
R749 B.n176 B.n175 163.367
R750 B.n175 B.n160 163.367
R751 B.n171 B.n160 163.367
R752 B.n171 B.n170 163.367
R753 B.n170 B.n169 163.367
R754 B.n169 B.n162 163.367
R755 B.n165 B.n162 163.367
R756 B.n165 B.n164 163.367
R757 B.n164 B.n2 163.367
R758 B.n622 B.n2 163.367
R759 B.n622 B.n621 163.367
R760 B.n621 B.n620 163.367
R761 B.n620 B.n3 163.367
R762 B.n616 B.n3 163.367
R763 B.n616 B.n615 163.367
R764 B.n615 B.n614 163.367
R765 B.n614 B.n5 163.367
R766 B.n610 B.n5 163.367
R767 B.n610 B.n609 163.367
R768 B.n609 B.n608 163.367
R769 B.n608 B.n7 163.367
R770 B.n604 B.n7 163.367
R771 B.n604 B.n603 163.367
R772 B.n603 B.n602 163.367
R773 B.n602 B.n9 163.367
R774 B.n598 B.n9 163.367
R775 B.n598 B.n597 163.367
R776 B.n597 B.n596 163.367
R777 B.n596 B.n11 163.367
R778 B.n592 B.n11 163.367
R779 B.n592 B.n591 163.367
R780 B.n591 B.n590 163.367
R781 B.n590 B.n13 163.367
R782 B.n586 B.n13 163.367
R783 B.n586 B.n585 163.367
R784 B.n585 B.n584 163.367
R785 B.n584 B.n15 163.367
R786 B.n580 B.n15 163.367
R787 B.n580 B.n579 163.367
R788 B.n579 B.n578 163.367
R789 B.n578 B.n17 163.367
R790 B.n574 B.n17 163.367
R791 B.n574 B.n573 163.367
R792 B.n573 B.n572 163.367
R793 B.n572 B.n19 163.367
R794 B.n568 B.n19 163.367
R795 B.n568 B.n567 163.367
R796 B.n567 B.n566 163.367
R797 B.n566 B.n21 163.367
R798 B.n562 B.n21 163.367
R799 B.n562 B.n561 163.367
R800 B.n561 B.n560 163.367
R801 B.n560 B.n23 163.367
R802 B.n556 B.n23 163.367
R803 B.n556 B.n555 163.367
R804 B.n555 B.n554 163.367
R805 B.n554 B.n25 163.367
R806 B.n550 B.n25 163.367
R807 B.n550 B.n549 163.367
R808 B.n549 B.n548 163.367
R809 B.n548 B.n27 163.367
R810 B.n544 B.n27 163.367
R811 B.n544 B.n543 163.367
R812 B.n543 B.n542 163.367
R813 B.n542 B.n29 163.367
R814 B.n247 B.n136 163.367
R815 B.n248 B.n247 163.367
R816 B.n249 B.n248 163.367
R817 B.n249 B.n134 163.367
R818 B.n253 B.n134 163.367
R819 B.n254 B.n253 163.367
R820 B.n255 B.n254 163.367
R821 B.n255 B.n132 163.367
R822 B.n259 B.n132 163.367
R823 B.n260 B.n259 163.367
R824 B.n261 B.n260 163.367
R825 B.n261 B.n130 163.367
R826 B.n265 B.n130 163.367
R827 B.n266 B.n265 163.367
R828 B.n267 B.n266 163.367
R829 B.n267 B.n126 163.367
R830 B.n272 B.n126 163.367
R831 B.n273 B.n272 163.367
R832 B.n274 B.n273 163.367
R833 B.n274 B.n124 163.367
R834 B.n278 B.n124 163.367
R835 B.n279 B.n278 163.367
R836 B.n280 B.n279 163.367
R837 B.n280 B.n122 163.367
R838 B.n284 B.n122 163.367
R839 B.n285 B.n284 163.367
R840 B.n285 B.n118 163.367
R841 B.n289 B.n118 163.367
R842 B.n290 B.n289 163.367
R843 B.n291 B.n290 163.367
R844 B.n291 B.n116 163.367
R845 B.n295 B.n116 163.367
R846 B.n296 B.n295 163.367
R847 B.n297 B.n296 163.367
R848 B.n297 B.n114 163.367
R849 B.n301 B.n114 163.367
R850 B.n302 B.n301 163.367
R851 B.n303 B.n302 163.367
R852 B.n303 B.n112 163.367
R853 B.n307 B.n112 163.367
R854 B.n308 B.n307 163.367
R855 B.n309 B.n110 163.367
R856 B.n313 B.n110 163.367
R857 B.n314 B.n313 163.367
R858 B.n315 B.n314 163.367
R859 B.n315 B.n108 163.367
R860 B.n319 B.n108 163.367
R861 B.n320 B.n319 163.367
R862 B.n321 B.n320 163.367
R863 B.n321 B.n106 163.367
R864 B.n325 B.n106 163.367
R865 B.n326 B.n325 163.367
R866 B.n327 B.n326 163.367
R867 B.n327 B.n104 163.367
R868 B.n331 B.n104 163.367
R869 B.n332 B.n331 163.367
R870 B.n333 B.n332 163.367
R871 B.n333 B.n102 163.367
R872 B.n337 B.n102 163.367
R873 B.n338 B.n337 163.367
R874 B.n339 B.n338 163.367
R875 B.n339 B.n100 163.367
R876 B.n343 B.n100 163.367
R877 B.n344 B.n343 163.367
R878 B.n345 B.n344 163.367
R879 B.n345 B.n98 163.367
R880 B.n349 B.n98 163.367
R881 B.n350 B.n349 163.367
R882 B.n351 B.n350 163.367
R883 B.n351 B.n96 163.367
R884 B.n355 B.n96 163.367
R885 B.n356 B.n355 163.367
R886 B.n357 B.n356 163.367
R887 B.n357 B.n94 163.367
R888 B.n361 B.n94 163.367
R889 B.n362 B.n361 163.367
R890 B.n363 B.n362 163.367
R891 B.n363 B.n92 163.367
R892 B.n367 B.n92 163.367
R893 B.n368 B.n367 163.367
R894 B.n369 B.n368 163.367
R895 B.n369 B.n90 163.367
R896 B.n373 B.n90 163.367
R897 B.n374 B.n373 163.367
R898 B.n375 B.n374 163.367
R899 B.n375 B.n88 163.367
R900 B.n379 B.n88 163.367
R901 B.n380 B.n379 163.367
R902 B.n381 B.n380 163.367
R903 B.n381 B.n86 163.367
R904 B.n385 B.n86 163.367
R905 B.n386 B.n385 163.367
R906 B.n387 B.n386 163.367
R907 B.n387 B.n84 163.367
R908 B.n391 B.n84 163.367
R909 B.n392 B.n391 163.367
R910 B.n393 B.n392 163.367
R911 B.n393 B.n82 163.367
R912 B.n397 B.n82 163.367
R913 B.n398 B.n397 163.367
R914 B.n399 B.n398 163.367
R915 B.n399 B.n80 163.367
R916 B.n403 B.n80 163.367
R917 B.n404 B.n403 163.367
R918 B.n405 B.n404 163.367
R919 B.n405 B.n78 163.367
R920 B.n409 B.n78 163.367
R921 B.n410 B.n409 163.367
R922 B.n411 B.n410 163.367
R923 B.n411 B.n76 163.367
R924 B.n415 B.n76 163.367
R925 B.n416 B.n415 163.367
R926 B.n417 B.n416 163.367
R927 B.n417 B.n74 163.367
R928 B.n421 B.n74 163.367
R929 B.n422 B.n421 163.367
R930 B.n423 B.n422 163.367
R931 B.n423 B.n72 163.367
R932 B.n427 B.n72 163.367
R933 B.n428 B.n427 163.367
R934 B.n429 B.n428 163.367
R935 B.n429 B.n70 163.367
R936 B.n433 B.n70 163.367
R937 B.n434 B.n433 163.367
R938 B.n435 B.n434 163.367
R939 B.n435 B.n68 163.367
R940 B.n439 B.n68 163.367
R941 B.n440 B.n439 163.367
R942 B.n441 B.n440 163.367
R943 B.n441 B.n66 163.367
R944 B.n445 B.n66 163.367
R945 B.n446 B.n445 163.367
R946 B.n447 B.n446 163.367
R947 B.n447 B.n64 163.367
R948 B.n451 B.n64 163.367
R949 B.n452 B.n451 163.367
R950 B.n453 B.n452 163.367
R951 B.n453 B.n62 163.367
R952 B.n457 B.n62 163.367
R953 B.n458 B.n457 163.367
R954 B.n459 B.n458 163.367
R955 B.n459 B.n60 163.367
R956 B.n463 B.n60 163.367
R957 B.n464 B.n463 163.367
R958 B.n465 B.n464 163.367
R959 B.n465 B.n58 163.367
R960 B.n469 B.n58 163.367
R961 B.n470 B.n469 163.367
R962 B.n471 B.n470 163.367
R963 B.n471 B.n56 163.367
R964 B.n475 B.n56 163.367
R965 B.n538 B.n537 163.367
R966 B.n537 B.n536 163.367
R967 B.n536 B.n31 163.367
R968 B.n532 B.n31 163.367
R969 B.n532 B.n531 163.367
R970 B.n531 B.n530 163.367
R971 B.n530 B.n33 163.367
R972 B.n526 B.n33 163.367
R973 B.n526 B.n525 163.367
R974 B.n525 B.n524 163.367
R975 B.n524 B.n35 163.367
R976 B.n520 B.n35 163.367
R977 B.n520 B.n519 163.367
R978 B.n519 B.n518 163.367
R979 B.n518 B.n37 163.367
R980 B.n513 B.n37 163.367
R981 B.n513 B.n512 163.367
R982 B.n512 B.n511 163.367
R983 B.n511 B.n41 163.367
R984 B.n507 B.n41 163.367
R985 B.n507 B.n506 163.367
R986 B.n506 B.n505 163.367
R987 B.n505 B.n43 163.367
R988 B.n501 B.n43 163.367
R989 B.n501 B.n500 163.367
R990 B.n500 B.n499 163.367
R991 B.n499 B.n45 163.367
R992 B.n495 B.n45 163.367
R993 B.n495 B.n494 163.367
R994 B.n494 B.n493 163.367
R995 B.n493 B.n50 163.367
R996 B.n489 B.n50 163.367
R997 B.n489 B.n488 163.367
R998 B.n488 B.n487 163.367
R999 B.n487 B.n52 163.367
R1000 B.n483 B.n52 163.367
R1001 B.n483 B.n482 163.367
R1002 B.n482 B.n481 163.367
R1003 B.n481 B.n54 163.367
R1004 B.n477 B.n54 163.367
R1005 B.n477 B.n476 163.367
R1006 B.n120 B.n119 77.1884
R1007 B.n128 B.n127 77.1884
R1008 B.n39 B.n38 77.1884
R1009 B.n47 B.n46 77.1884
R1010 B.n121 B.n120 59.5399
R1011 B.n269 B.n128 59.5399
R1012 B.n515 B.n39 59.5399
R1013 B.n48 B.n47 59.5399
R1014 B.n474 B.n55 29.5029
R1015 B.n540 B.n539 29.5029
R1016 B.n310 B.n111 29.5029
R1017 B.n245 B.n244 29.5029
R1018 B B.n623 18.0485
R1019 B.n539 B.n30 10.6151
R1020 B.n535 B.n30 10.6151
R1021 B.n535 B.n534 10.6151
R1022 B.n534 B.n533 10.6151
R1023 B.n533 B.n32 10.6151
R1024 B.n529 B.n32 10.6151
R1025 B.n529 B.n528 10.6151
R1026 B.n528 B.n527 10.6151
R1027 B.n527 B.n34 10.6151
R1028 B.n523 B.n34 10.6151
R1029 B.n523 B.n522 10.6151
R1030 B.n522 B.n521 10.6151
R1031 B.n521 B.n36 10.6151
R1032 B.n517 B.n36 10.6151
R1033 B.n517 B.n516 10.6151
R1034 B.n514 B.n40 10.6151
R1035 B.n510 B.n40 10.6151
R1036 B.n510 B.n509 10.6151
R1037 B.n509 B.n508 10.6151
R1038 B.n508 B.n42 10.6151
R1039 B.n504 B.n42 10.6151
R1040 B.n504 B.n503 10.6151
R1041 B.n503 B.n502 10.6151
R1042 B.n502 B.n44 10.6151
R1043 B.n498 B.n497 10.6151
R1044 B.n497 B.n496 10.6151
R1045 B.n496 B.n49 10.6151
R1046 B.n492 B.n49 10.6151
R1047 B.n492 B.n491 10.6151
R1048 B.n491 B.n490 10.6151
R1049 B.n490 B.n51 10.6151
R1050 B.n486 B.n51 10.6151
R1051 B.n486 B.n485 10.6151
R1052 B.n485 B.n484 10.6151
R1053 B.n484 B.n53 10.6151
R1054 B.n480 B.n53 10.6151
R1055 B.n480 B.n479 10.6151
R1056 B.n479 B.n478 10.6151
R1057 B.n478 B.n55 10.6151
R1058 B.n311 B.n310 10.6151
R1059 B.n312 B.n311 10.6151
R1060 B.n312 B.n109 10.6151
R1061 B.n316 B.n109 10.6151
R1062 B.n317 B.n316 10.6151
R1063 B.n318 B.n317 10.6151
R1064 B.n318 B.n107 10.6151
R1065 B.n322 B.n107 10.6151
R1066 B.n323 B.n322 10.6151
R1067 B.n324 B.n323 10.6151
R1068 B.n324 B.n105 10.6151
R1069 B.n328 B.n105 10.6151
R1070 B.n329 B.n328 10.6151
R1071 B.n330 B.n329 10.6151
R1072 B.n330 B.n103 10.6151
R1073 B.n334 B.n103 10.6151
R1074 B.n335 B.n334 10.6151
R1075 B.n336 B.n335 10.6151
R1076 B.n336 B.n101 10.6151
R1077 B.n340 B.n101 10.6151
R1078 B.n341 B.n340 10.6151
R1079 B.n342 B.n341 10.6151
R1080 B.n342 B.n99 10.6151
R1081 B.n346 B.n99 10.6151
R1082 B.n347 B.n346 10.6151
R1083 B.n348 B.n347 10.6151
R1084 B.n348 B.n97 10.6151
R1085 B.n352 B.n97 10.6151
R1086 B.n353 B.n352 10.6151
R1087 B.n354 B.n353 10.6151
R1088 B.n354 B.n95 10.6151
R1089 B.n358 B.n95 10.6151
R1090 B.n359 B.n358 10.6151
R1091 B.n360 B.n359 10.6151
R1092 B.n360 B.n93 10.6151
R1093 B.n364 B.n93 10.6151
R1094 B.n365 B.n364 10.6151
R1095 B.n366 B.n365 10.6151
R1096 B.n366 B.n91 10.6151
R1097 B.n370 B.n91 10.6151
R1098 B.n371 B.n370 10.6151
R1099 B.n372 B.n371 10.6151
R1100 B.n372 B.n89 10.6151
R1101 B.n376 B.n89 10.6151
R1102 B.n377 B.n376 10.6151
R1103 B.n378 B.n377 10.6151
R1104 B.n378 B.n87 10.6151
R1105 B.n382 B.n87 10.6151
R1106 B.n383 B.n382 10.6151
R1107 B.n384 B.n383 10.6151
R1108 B.n384 B.n85 10.6151
R1109 B.n388 B.n85 10.6151
R1110 B.n389 B.n388 10.6151
R1111 B.n390 B.n389 10.6151
R1112 B.n390 B.n83 10.6151
R1113 B.n394 B.n83 10.6151
R1114 B.n395 B.n394 10.6151
R1115 B.n396 B.n395 10.6151
R1116 B.n396 B.n81 10.6151
R1117 B.n400 B.n81 10.6151
R1118 B.n401 B.n400 10.6151
R1119 B.n402 B.n401 10.6151
R1120 B.n402 B.n79 10.6151
R1121 B.n406 B.n79 10.6151
R1122 B.n407 B.n406 10.6151
R1123 B.n408 B.n407 10.6151
R1124 B.n408 B.n77 10.6151
R1125 B.n412 B.n77 10.6151
R1126 B.n413 B.n412 10.6151
R1127 B.n414 B.n413 10.6151
R1128 B.n414 B.n75 10.6151
R1129 B.n418 B.n75 10.6151
R1130 B.n419 B.n418 10.6151
R1131 B.n420 B.n419 10.6151
R1132 B.n420 B.n73 10.6151
R1133 B.n424 B.n73 10.6151
R1134 B.n425 B.n424 10.6151
R1135 B.n426 B.n425 10.6151
R1136 B.n426 B.n71 10.6151
R1137 B.n430 B.n71 10.6151
R1138 B.n431 B.n430 10.6151
R1139 B.n432 B.n431 10.6151
R1140 B.n432 B.n69 10.6151
R1141 B.n436 B.n69 10.6151
R1142 B.n437 B.n436 10.6151
R1143 B.n438 B.n437 10.6151
R1144 B.n438 B.n67 10.6151
R1145 B.n442 B.n67 10.6151
R1146 B.n443 B.n442 10.6151
R1147 B.n444 B.n443 10.6151
R1148 B.n444 B.n65 10.6151
R1149 B.n448 B.n65 10.6151
R1150 B.n449 B.n448 10.6151
R1151 B.n450 B.n449 10.6151
R1152 B.n450 B.n63 10.6151
R1153 B.n454 B.n63 10.6151
R1154 B.n455 B.n454 10.6151
R1155 B.n456 B.n455 10.6151
R1156 B.n456 B.n61 10.6151
R1157 B.n460 B.n61 10.6151
R1158 B.n461 B.n460 10.6151
R1159 B.n462 B.n461 10.6151
R1160 B.n462 B.n59 10.6151
R1161 B.n466 B.n59 10.6151
R1162 B.n467 B.n466 10.6151
R1163 B.n468 B.n467 10.6151
R1164 B.n468 B.n57 10.6151
R1165 B.n472 B.n57 10.6151
R1166 B.n473 B.n472 10.6151
R1167 B.n474 B.n473 10.6151
R1168 B.n246 B.n245 10.6151
R1169 B.n246 B.n135 10.6151
R1170 B.n250 B.n135 10.6151
R1171 B.n251 B.n250 10.6151
R1172 B.n252 B.n251 10.6151
R1173 B.n252 B.n133 10.6151
R1174 B.n256 B.n133 10.6151
R1175 B.n257 B.n256 10.6151
R1176 B.n258 B.n257 10.6151
R1177 B.n258 B.n131 10.6151
R1178 B.n262 B.n131 10.6151
R1179 B.n263 B.n262 10.6151
R1180 B.n264 B.n263 10.6151
R1181 B.n264 B.n129 10.6151
R1182 B.n268 B.n129 10.6151
R1183 B.n271 B.n270 10.6151
R1184 B.n271 B.n125 10.6151
R1185 B.n275 B.n125 10.6151
R1186 B.n276 B.n275 10.6151
R1187 B.n277 B.n276 10.6151
R1188 B.n277 B.n123 10.6151
R1189 B.n281 B.n123 10.6151
R1190 B.n282 B.n281 10.6151
R1191 B.n283 B.n282 10.6151
R1192 B.n287 B.n286 10.6151
R1193 B.n288 B.n287 10.6151
R1194 B.n288 B.n117 10.6151
R1195 B.n292 B.n117 10.6151
R1196 B.n293 B.n292 10.6151
R1197 B.n294 B.n293 10.6151
R1198 B.n294 B.n115 10.6151
R1199 B.n298 B.n115 10.6151
R1200 B.n299 B.n298 10.6151
R1201 B.n300 B.n299 10.6151
R1202 B.n300 B.n113 10.6151
R1203 B.n304 B.n113 10.6151
R1204 B.n305 B.n304 10.6151
R1205 B.n306 B.n305 10.6151
R1206 B.n306 B.n111 10.6151
R1207 B.n244 B.n137 10.6151
R1208 B.n240 B.n137 10.6151
R1209 B.n240 B.n239 10.6151
R1210 B.n239 B.n238 10.6151
R1211 B.n238 B.n139 10.6151
R1212 B.n234 B.n139 10.6151
R1213 B.n234 B.n233 10.6151
R1214 B.n233 B.n232 10.6151
R1215 B.n232 B.n141 10.6151
R1216 B.n228 B.n141 10.6151
R1217 B.n228 B.n227 10.6151
R1218 B.n227 B.n226 10.6151
R1219 B.n226 B.n143 10.6151
R1220 B.n222 B.n143 10.6151
R1221 B.n222 B.n221 10.6151
R1222 B.n221 B.n220 10.6151
R1223 B.n220 B.n145 10.6151
R1224 B.n216 B.n145 10.6151
R1225 B.n216 B.n215 10.6151
R1226 B.n215 B.n214 10.6151
R1227 B.n214 B.n147 10.6151
R1228 B.n210 B.n147 10.6151
R1229 B.n210 B.n209 10.6151
R1230 B.n209 B.n208 10.6151
R1231 B.n208 B.n149 10.6151
R1232 B.n204 B.n149 10.6151
R1233 B.n204 B.n203 10.6151
R1234 B.n203 B.n202 10.6151
R1235 B.n202 B.n151 10.6151
R1236 B.n198 B.n151 10.6151
R1237 B.n198 B.n197 10.6151
R1238 B.n197 B.n196 10.6151
R1239 B.n196 B.n153 10.6151
R1240 B.n192 B.n153 10.6151
R1241 B.n192 B.n191 10.6151
R1242 B.n191 B.n190 10.6151
R1243 B.n190 B.n155 10.6151
R1244 B.n186 B.n155 10.6151
R1245 B.n186 B.n185 10.6151
R1246 B.n185 B.n184 10.6151
R1247 B.n184 B.n157 10.6151
R1248 B.n180 B.n157 10.6151
R1249 B.n180 B.n179 10.6151
R1250 B.n179 B.n178 10.6151
R1251 B.n178 B.n159 10.6151
R1252 B.n174 B.n159 10.6151
R1253 B.n174 B.n173 10.6151
R1254 B.n173 B.n172 10.6151
R1255 B.n172 B.n161 10.6151
R1256 B.n168 B.n161 10.6151
R1257 B.n168 B.n167 10.6151
R1258 B.n167 B.n166 10.6151
R1259 B.n166 B.n163 10.6151
R1260 B.n163 B.n0 10.6151
R1261 B.n619 B.n1 10.6151
R1262 B.n619 B.n618 10.6151
R1263 B.n618 B.n617 10.6151
R1264 B.n617 B.n4 10.6151
R1265 B.n613 B.n4 10.6151
R1266 B.n613 B.n612 10.6151
R1267 B.n612 B.n611 10.6151
R1268 B.n611 B.n6 10.6151
R1269 B.n607 B.n6 10.6151
R1270 B.n607 B.n606 10.6151
R1271 B.n606 B.n605 10.6151
R1272 B.n605 B.n8 10.6151
R1273 B.n601 B.n8 10.6151
R1274 B.n601 B.n600 10.6151
R1275 B.n600 B.n599 10.6151
R1276 B.n599 B.n10 10.6151
R1277 B.n595 B.n10 10.6151
R1278 B.n595 B.n594 10.6151
R1279 B.n594 B.n593 10.6151
R1280 B.n593 B.n12 10.6151
R1281 B.n589 B.n12 10.6151
R1282 B.n589 B.n588 10.6151
R1283 B.n588 B.n587 10.6151
R1284 B.n587 B.n14 10.6151
R1285 B.n583 B.n14 10.6151
R1286 B.n583 B.n582 10.6151
R1287 B.n582 B.n581 10.6151
R1288 B.n581 B.n16 10.6151
R1289 B.n577 B.n16 10.6151
R1290 B.n577 B.n576 10.6151
R1291 B.n576 B.n575 10.6151
R1292 B.n575 B.n18 10.6151
R1293 B.n571 B.n18 10.6151
R1294 B.n571 B.n570 10.6151
R1295 B.n570 B.n569 10.6151
R1296 B.n569 B.n20 10.6151
R1297 B.n565 B.n20 10.6151
R1298 B.n565 B.n564 10.6151
R1299 B.n564 B.n563 10.6151
R1300 B.n563 B.n22 10.6151
R1301 B.n559 B.n22 10.6151
R1302 B.n559 B.n558 10.6151
R1303 B.n558 B.n557 10.6151
R1304 B.n557 B.n24 10.6151
R1305 B.n553 B.n24 10.6151
R1306 B.n553 B.n552 10.6151
R1307 B.n552 B.n551 10.6151
R1308 B.n551 B.n26 10.6151
R1309 B.n547 B.n26 10.6151
R1310 B.n547 B.n546 10.6151
R1311 B.n546 B.n545 10.6151
R1312 B.n545 B.n28 10.6151
R1313 B.n541 B.n28 10.6151
R1314 B.n541 B.n540 10.6151
R1315 B.n516 B.n515 9.36635
R1316 B.n498 B.n48 9.36635
R1317 B.n269 B.n268 9.36635
R1318 B.n286 B.n121 9.36635
R1319 B.n623 B.n0 2.81026
R1320 B.n623 B.n1 2.81026
R1321 B.n515 B.n514 1.24928
R1322 B.n48 B.n44 1.24928
R1323 B.n270 B.n269 1.24928
R1324 B.n283 B.n121 1.24928
C0 VDD1 B 1.66336f
C1 VP B 2.20467f
C2 VDD2 w_n4154_n1626# 2.06744f
C3 VTAIL VN 3.32284f
C4 VDD2 VDD1 1.81666f
C5 VP VDD2 0.552502f
C6 w_n4154_n1626# VN 7.96186f
C7 VDD2 B 1.7629f
C8 VTAIL w_n4154_n1626# 1.86773f
C9 VDD1 VN 0.157127f
C10 VTAIL VDD1 5.28253f
C11 VP VN 6.33803f
C12 VP VTAIL 3.33703f
C13 B VN 1.29818f
C14 VTAIL B 1.94818f
C15 w_n4154_n1626# VDD1 1.94926f
C16 VP w_n4154_n1626# 8.499969f
C17 VDD2 VN 2.24179f
C18 VTAIL VDD2 5.34269f
C19 VP VDD1 2.63436f
C20 w_n4154_n1626# B 8.725441f
C21 VDD2 VSUBS 1.762395f
C22 VDD1 VSUBS 1.818268f
C23 VTAIL VSUBS 0.66579f
C24 VN VSUBS 6.82621f
C25 VP VSUBS 3.182844f
C26 B VSUBS 4.643898f
C27 w_n4154_n1626# VSUBS 85.3896f
C28 B.n0 VSUBS 0.005866f
C29 B.n1 VSUBS 0.005866f
C30 B.n2 VSUBS 0.009276f
C31 B.n3 VSUBS 0.009276f
C32 B.n4 VSUBS 0.009276f
C33 B.n5 VSUBS 0.009276f
C34 B.n6 VSUBS 0.009276f
C35 B.n7 VSUBS 0.009276f
C36 B.n8 VSUBS 0.009276f
C37 B.n9 VSUBS 0.009276f
C38 B.n10 VSUBS 0.009276f
C39 B.n11 VSUBS 0.009276f
C40 B.n12 VSUBS 0.009276f
C41 B.n13 VSUBS 0.009276f
C42 B.n14 VSUBS 0.009276f
C43 B.n15 VSUBS 0.009276f
C44 B.n16 VSUBS 0.009276f
C45 B.n17 VSUBS 0.009276f
C46 B.n18 VSUBS 0.009276f
C47 B.n19 VSUBS 0.009276f
C48 B.n20 VSUBS 0.009276f
C49 B.n21 VSUBS 0.009276f
C50 B.n22 VSUBS 0.009276f
C51 B.n23 VSUBS 0.009276f
C52 B.n24 VSUBS 0.009276f
C53 B.n25 VSUBS 0.009276f
C54 B.n26 VSUBS 0.009276f
C55 B.n27 VSUBS 0.009276f
C56 B.n28 VSUBS 0.009276f
C57 B.n29 VSUBS 0.019601f
C58 B.n30 VSUBS 0.009276f
C59 B.n31 VSUBS 0.009276f
C60 B.n32 VSUBS 0.009276f
C61 B.n33 VSUBS 0.009276f
C62 B.n34 VSUBS 0.009276f
C63 B.n35 VSUBS 0.009276f
C64 B.n36 VSUBS 0.009276f
C65 B.n37 VSUBS 0.009276f
C66 B.t11 VSUBS 0.064468f
C67 B.t10 VSUBS 0.095935f
C68 B.t9 VSUBS 0.778307f
C69 B.n38 VSUBS 0.164417f
C70 B.n39 VSUBS 0.13736f
C71 B.n40 VSUBS 0.009276f
C72 B.n41 VSUBS 0.009276f
C73 B.n42 VSUBS 0.009276f
C74 B.n43 VSUBS 0.009276f
C75 B.n44 VSUBS 0.005184f
C76 B.n45 VSUBS 0.009276f
C77 B.t5 VSUBS 0.064469f
C78 B.t4 VSUBS 0.095935f
C79 B.t3 VSUBS 0.778307f
C80 B.n46 VSUBS 0.164416f
C81 B.n47 VSUBS 0.137359f
C82 B.n48 VSUBS 0.021493f
C83 B.n49 VSUBS 0.009276f
C84 B.n50 VSUBS 0.009276f
C85 B.n51 VSUBS 0.009276f
C86 B.n52 VSUBS 0.009276f
C87 B.n53 VSUBS 0.009276f
C88 B.n54 VSUBS 0.009276f
C89 B.n55 VSUBS 0.019838f
C90 B.n56 VSUBS 0.009276f
C91 B.n57 VSUBS 0.009276f
C92 B.n58 VSUBS 0.009276f
C93 B.n59 VSUBS 0.009276f
C94 B.n60 VSUBS 0.009276f
C95 B.n61 VSUBS 0.009276f
C96 B.n62 VSUBS 0.009276f
C97 B.n63 VSUBS 0.009276f
C98 B.n64 VSUBS 0.009276f
C99 B.n65 VSUBS 0.009276f
C100 B.n66 VSUBS 0.009276f
C101 B.n67 VSUBS 0.009276f
C102 B.n68 VSUBS 0.009276f
C103 B.n69 VSUBS 0.009276f
C104 B.n70 VSUBS 0.009276f
C105 B.n71 VSUBS 0.009276f
C106 B.n72 VSUBS 0.009276f
C107 B.n73 VSUBS 0.009276f
C108 B.n74 VSUBS 0.009276f
C109 B.n75 VSUBS 0.009276f
C110 B.n76 VSUBS 0.009276f
C111 B.n77 VSUBS 0.009276f
C112 B.n78 VSUBS 0.009276f
C113 B.n79 VSUBS 0.009276f
C114 B.n80 VSUBS 0.009276f
C115 B.n81 VSUBS 0.009276f
C116 B.n82 VSUBS 0.009276f
C117 B.n83 VSUBS 0.009276f
C118 B.n84 VSUBS 0.009276f
C119 B.n85 VSUBS 0.009276f
C120 B.n86 VSUBS 0.009276f
C121 B.n87 VSUBS 0.009276f
C122 B.n88 VSUBS 0.009276f
C123 B.n89 VSUBS 0.009276f
C124 B.n90 VSUBS 0.009276f
C125 B.n91 VSUBS 0.009276f
C126 B.n92 VSUBS 0.009276f
C127 B.n93 VSUBS 0.009276f
C128 B.n94 VSUBS 0.009276f
C129 B.n95 VSUBS 0.009276f
C130 B.n96 VSUBS 0.009276f
C131 B.n97 VSUBS 0.009276f
C132 B.n98 VSUBS 0.009276f
C133 B.n99 VSUBS 0.009276f
C134 B.n100 VSUBS 0.009276f
C135 B.n101 VSUBS 0.009276f
C136 B.n102 VSUBS 0.009276f
C137 B.n103 VSUBS 0.009276f
C138 B.n104 VSUBS 0.009276f
C139 B.n105 VSUBS 0.009276f
C140 B.n106 VSUBS 0.009276f
C141 B.n107 VSUBS 0.009276f
C142 B.n108 VSUBS 0.009276f
C143 B.n109 VSUBS 0.009276f
C144 B.n110 VSUBS 0.009276f
C145 B.n111 VSUBS 0.021051f
C146 B.n112 VSUBS 0.009276f
C147 B.n113 VSUBS 0.009276f
C148 B.n114 VSUBS 0.009276f
C149 B.n115 VSUBS 0.009276f
C150 B.n116 VSUBS 0.009276f
C151 B.n117 VSUBS 0.009276f
C152 B.n118 VSUBS 0.009276f
C153 B.t1 VSUBS 0.064469f
C154 B.t2 VSUBS 0.095935f
C155 B.t0 VSUBS 0.778307f
C156 B.n119 VSUBS 0.164416f
C157 B.n120 VSUBS 0.137359f
C158 B.n121 VSUBS 0.021493f
C159 B.n122 VSUBS 0.009276f
C160 B.n123 VSUBS 0.009276f
C161 B.n124 VSUBS 0.009276f
C162 B.n125 VSUBS 0.009276f
C163 B.n126 VSUBS 0.009276f
C164 B.t7 VSUBS 0.064468f
C165 B.t8 VSUBS 0.095935f
C166 B.t6 VSUBS 0.778307f
C167 B.n127 VSUBS 0.164417f
C168 B.n128 VSUBS 0.13736f
C169 B.n129 VSUBS 0.009276f
C170 B.n130 VSUBS 0.009276f
C171 B.n131 VSUBS 0.009276f
C172 B.n132 VSUBS 0.009276f
C173 B.n133 VSUBS 0.009276f
C174 B.n134 VSUBS 0.009276f
C175 B.n135 VSUBS 0.009276f
C176 B.n136 VSUBS 0.021051f
C177 B.n137 VSUBS 0.009276f
C178 B.n138 VSUBS 0.009276f
C179 B.n139 VSUBS 0.009276f
C180 B.n140 VSUBS 0.009276f
C181 B.n141 VSUBS 0.009276f
C182 B.n142 VSUBS 0.009276f
C183 B.n143 VSUBS 0.009276f
C184 B.n144 VSUBS 0.009276f
C185 B.n145 VSUBS 0.009276f
C186 B.n146 VSUBS 0.009276f
C187 B.n147 VSUBS 0.009276f
C188 B.n148 VSUBS 0.009276f
C189 B.n149 VSUBS 0.009276f
C190 B.n150 VSUBS 0.009276f
C191 B.n151 VSUBS 0.009276f
C192 B.n152 VSUBS 0.009276f
C193 B.n153 VSUBS 0.009276f
C194 B.n154 VSUBS 0.009276f
C195 B.n155 VSUBS 0.009276f
C196 B.n156 VSUBS 0.009276f
C197 B.n157 VSUBS 0.009276f
C198 B.n158 VSUBS 0.009276f
C199 B.n159 VSUBS 0.009276f
C200 B.n160 VSUBS 0.009276f
C201 B.n161 VSUBS 0.009276f
C202 B.n162 VSUBS 0.009276f
C203 B.n163 VSUBS 0.009276f
C204 B.n164 VSUBS 0.009276f
C205 B.n165 VSUBS 0.009276f
C206 B.n166 VSUBS 0.009276f
C207 B.n167 VSUBS 0.009276f
C208 B.n168 VSUBS 0.009276f
C209 B.n169 VSUBS 0.009276f
C210 B.n170 VSUBS 0.009276f
C211 B.n171 VSUBS 0.009276f
C212 B.n172 VSUBS 0.009276f
C213 B.n173 VSUBS 0.009276f
C214 B.n174 VSUBS 0.009276f
C215 B.n175 VSUBS 0.009276f
C216 B.n176 VSUBS 0.009276f
C217 B.n177 VSUBS 0.009276f
C218 B.n178 VSUBS 0.009276f
C219 B.n179 VSUBS 0.009276f
C220 B.n180 VSUBS 0.009276f
C221 B.n181 VSUBS 0.009276f
C222 B.n182 VSUBS 0.009276f
C223 B.n183 VSUBS 0.009276f
C224 B.n184 VSUBS 0.009276f
C225 B.n185 VSUBS 0.009276f
C226 B.n186 VSUBS 0.009276f
C227 B.n187 VSUBS 0.009276f
C228 B.n188 VSUBS 0.009276f
C229 B.n189 VSUBS 0.009276f
C230 B.n190 VSUBS 0.009276f
C231 B.n191 VSUBS 0.009276f
C232 B.n192 VSUBS 0.009276f
C233 B.n193 VSUBS 0.009276f
C234 B.n194 VSUBS 0.009276f
C235 B.n195 VSUBS 0.009276f
C236 B.n196 VSUBS 0.009276f
C237 B.n197 VSUBS 0.009276f
C238 B.n198 VSUBS 0.009276f
C239 B.n199 VSUBS 0.009276f
C240 B.n200 VSUBS 0.009276f
C241 B.n201 VSUBS 0.009276f
C242 B.n202 VSUBS 0.009276f
C243 B.n203 VSUBS 0.009276f
C244 B.n204 VSUBS 0.009276f
C245 B.n205 VSUBS 0.009276f
C246 B.n206 VSUBS 0.009276f
C247 B.n207 VSUBS 0.009276f
C248 B.n208 VSUBS 0.009276f
C249 B.n209 VSUBS 0.009276f
C250 B.n210 VSUBS 0.009276f
C251 B.n211 VSUBS 0.009276f
C252 B.n212 VSUBS 0.009276f
C253 B.n213 VSUBS 0.009276f
C254 B.n214 VSUBS 0.009276f
C255 B.n215 VSUBS 0.009276f
C256 B.n216 VSUBS 0.009276f
C257 B.n217 VSUBS 0.009276f
C258 B.n218 VSUBS 0.009276f
C259 B.n219 VSUBS 0.009276f
C260 B.n220 VSUBS 0.009276f
C261 B.n221 VSUBS 0.009276f
C262 B.n222 VSUBS 0.009276f
C263 B.n223 VSUBS 0.009276f
C264 B.n224 VSUBS 0.009276f
C265 B.n225 VSUBS 0.009276f
C266 B.n226 VSUBS 0.009276f
C267 B.n227 VSUBS 0.009276f
C268 B.n228 VSUBS 0.009276f
C269 B.n229 VSUBS 0.009276f
C270 B.n230 VSUBS 0.009276f
C271 B.n231 VSUBS 0.009276f
C272 B.n232 VSUBS 0.009276f
C273 B.n233 VSUBS 0.009276f
C274 B.n234 VSUBS 0.009276f
C275 B.n235 VSUBS 0.009276f
C276 B.n236 VSUBS 0.009276f
C277 B.n237 VSUBS 0.009276f
C278 B.n238 VSUBS 0.009276f
C279 B.n239 VSUBS 0.009276f
C280 B.n240 VSUBS 0.009276f
C281 B.n241 VSUBS 0.009276f
C282 B.n242 VSUBS 0.009276f
C283 B.n243 VSUBS 0.019601f
C284 B.n244 VSUBS 0.019601f
C285 B.n245 VSUBS 0.021051f
C286 B.n246 VSUBS 0.009276f
C287 B.n247 VSUBS 0.009276f
C288 B.n248 VSUBS 0.009276f
C289 B.n249 VSUBS 0.009276f
C290 B.n250 VSUBS 0.009276f
C291 B.n251 VSUBS 0.009276f
C292 B.n252 VSUBS 0.009276f
C293 B.n253 VSUBS 0.009276f
C294 B.n254 VSUBS 0.009276f
C295 B.n255 VSUBS 0.009276f
C296 B.n256 VSUBS 0.009276f
C297 B.n257 VSUBS 0.009276f
C298 B.n258 VSUBS 0.009276f
C299 B.n259 VSUBS 0.009276f
C300 B.n260 VSUBS 0.009276f
C301 B.n261 VSUBS 0.009276f
C302 B.n262 VSUBS 0.009276f
C303 B.n263 VSUBS 0.009276f
C304 B.n264 VSUBS 0.009276f
C305 B.n265 VSUBS 0.009276f
C306 B.n266 VSUBS 0.009276f
C307 B.n267 VSUBS 0.009276f
C308 B.n268 VSUBS 0.008731f
C309 B.n269 VSUBS 0.021493f
C310 B.n270 VSUBS 0.005184f
C311 B.n271 VSUBS 0.009276f
C312 B.n272 VSUBS 0.009276f
C313 B.n273 VSUBS 0.009276f
C314 B.n274 VSUBS 0.009276f
C315 B.n275 VSUBS 0.009276f
C316 B.n276 VSUBS 0.009276f
C317 B.n277 VSUBS 0.009276f
C318 B.n278 VSUBS 0.009276f
C319 B.n279 VSUBS 0.009276f
C320 B.n280 VSUBS 0.009276f
C321 B.n281 VSUBS 0.009276f
C322 B.n282 VSUBS 0.009276f
C323 B.n283 VSUBS 0.005184f
C324 B.n284 VSUBS 0.009276f
C325 B.n285 VSUBS 0.009276f
C326 B.n286 VSUBS 0.008731f
C327 B.n287 VSUBS 0.009276f
C328 B.n288 VSUBS 0.009276f
C329 B.n289 VSUBS 0.009276f
C330 B.n290 VSUBS 0.009276f
C331 B.n291 VSUBS 0.009276f
C332 B.n292 VSUBS 0.009276f
C333 B.n293 VSUBS 0.009276f
C334 B.n294 VSUBS 0.009276f
C335 B.n295 VSUBS 0.009276f
C336 B.n296 VSUBS 0.009276f
C337 B.n297 VSUBS 0.009276f
C338 B.n298 VSUBS 0.009276f
C339 B.n299 VSUBS 0.009276f
C340 B.n300 VSUBS 0.009276f
C341 B.n301 VSUBS 0.009276f
C342 B.n302 VSUBS 0.009276f
C343 B.n303 VSUBS 0.009276f
C344 B.n304 VSUBS 0.009276f
C345 B.n305 VSUBS 0.009276f
C346 B.n306 VSUBS 0.009276f
C347 B.n307 VSUBS 0.009276f
C348 B.n308 VSUBS 0.021051f
C349 B.n309 VSUBS 0.019601f
C350 B.n310 VSUBS 0.019601f
C351 B.n311 VSUBS 0.009276f
C352 B.n312 VSUBS 0.009276f
C353 B.n313 VSUBS 0.009276f
C354 B.n314 VSUBS 0.009276f
C355 B.n315 VSUBS 0.009276f
C356 B.n316 VSUBS 0.009276f
C357 B.n317 VSUBS 0.009276f
C358 B.n318 VSUBS 0.009276f
C359 B.n319 VSUBS 0.009276f
C360 B.n320 VSUBS 0.009276f
C361 B.n321 VSUBS 0.009276f
C362 B.n322 VSUBS 0.009276f
C363 B.n323 VSUBS 0.009276f
C364 B.n324 VSUBS 0.009276f
C365 B.n325 VSUBS 0.009276f
C366 B.n326 VSUBS 0.009276f
C367 B.n327 VSUBS 0.009276f
C368 B.n328 VSUBS 0.009276f
C369 B.n329 VSUBS 0.009276f
C370 B.n330 VSUBS 0.009276f
C371 B.n331 VSUBS 0.009276f
C372 B.n332 VSUBS 0.009276f
C373 B.n333 VSUBS 0.009276f
C374 B.n334 VSUBS 0.009276f
C375 B.n335 VSUBS 0.009276f
C376 B.n336 VSUBS 0.009276f
C377 B.n337 VSUBS 0.009276f
C378 B.n338 VSUBS 0.009276f
C379 B.n339 VSUBS 0.009276f
C380 B.n340 VSUBS 0.009276f
C381 B.n341 VSUBS 0.009276f
C382 B.n342 VSUBS 0.009276f
C383 B.n343 VSUBS 0.009276f
C384 B.n344 VSUBS 0.009276f
C385 B.n345 VSUBS 0.009276f
C386 B.n346 VSUBS 0.009276f
C387 B.n347 VSUBS 0.009276f
C388 B.n348 VSUBS 0.009276f
C389 B.n349 VSUBS 0.009276f
C390 B.n350 VSUBS 0.009276f
C391 B.n351 VSUBS 0.009276f
C392 B.n352 VSUBS 0.009276f
C393 B.n353 VSUBS 0.009276f
C394 B.n354 VSUBS 0.009276f
C395 B.n355 VSUBS 0.009276f
C396 B.n356 VSUBS 0.009276f
C397 B.n357 VSUBS 0.009276f
C398 B.n358 VSUBS 0.009276f
C399 B.n359 VSUBS 0.009276f
C400 B.n360 VSUBS 0.009276f
C401 B.n361 VSUBS 0.009276f
C402 B.n362 VSUBS 0.009276f
C403 B.n363 VSUBS 0.009276f
C404 B.n364 VSUBS 0.009276f
C405 B.n365 VSUBS 0.009276f
C406 B.n366 VSUBS 0.009276f
C407 B.n367 VSUBS 0.009276f
C408 B.n368 VSUBS 0.009276f
C409 B.n369 VSUBS 0.009276f
C410 B.n370 VSUBS 0.009276f
C411 B.n371 VSUBS 0.009276f
C412 B.n372 VSUBS 0.009276f
C413 B.n373 VSUBS 0.009276f
C414 B.n374 VSUBS 0.009276f
C415 B.n375 VSUBS 0.009276f
C416 B.n376 VSUBS 0.009276f
C417 B.n377 VSUBS 0.009276f
C418 B.n378 VSUBS 0.009276f
C419 B.n379 VSUBS 0.009276f
C420 B.n380 VSUBS 0.009276f
C421 B.n381 VSUBS 0.009276f
C422 B.n382 VSUBS 0.009276f
C423 B.n383 VSUBS 0.009276f
C424 B.n384 VSUBS 0.009276f
C425 B.n385 VSUBS 0.009276f
C426 B.n386 VSUBS 0.009276f
C427 B.n387 VSUBS 0.009276f
C428 B.n388 VSUBS 0.009276f
C429 B.n389 VSUBS 0.009276f
C430 B.n390 VSUBS 0.009276f
C431 B.n391 VSUBS 0.009276f
C432 B.n392 VSUBS 0.009276f
C433 B.n393 VSUBS 0.009276f
C434 B.n394 VSUBS 0.009276f
C435 B.n395 VSUBS 0.009276f
C436 B.n396 VSUBS 0.009276f
C437 B.n397 VSUBS 0.009276f
C438 B.n398 VSUBS 0.009276f
C439 B.n399 VSUBS 0.009276f
C440 B.n400 VSUBS 0.009276f
C441 B.n401 VSUBS 0.009276f
C442 B.n402 VSUBS 0.009276f
C443 B.n403 VSUBS 0.009276f
C444 B.n404 VSUBS 0.009276f
C445 B.n405 VSUBS 0.009276f
C446 B.n406 VSUBS 0.009276f
C447 B.n407 VSUBS 0.009276f
C448 B.n408 VSUBS 0.009276f
C449 B.n409 VSUBS 0.009276f
C450 B.n410 VSUBS 0.009276f
C451 B.n411 VSUBS 0.009276f
C452 B.n412 VSUBS 0.009276f
C453 B.n413 VSUBS 0.009276f
C454 B.n414 VSUBS 0.009276f
C455 B.n415 VSUBS 0.009276f
C456 B.n416 VSUBS 0.009276f
C457 B.n417 VSUBS 0.009276f
C458 B.n418 VSUBS 0.009276f
C459 B.n419 VSUBS 0.009276f
C460 B.n420 VSUBS 0.009276f
C461 B.n421 VSUBS 0.009276f
C462 B.n422 VSUBS 0.009276f
C463 B.n423 VSUBS 0.009276f
C464 B.n424 VSUBS 0.009276f
C465 B.n425 VSUBS 0.009276f
C466 B.n426 VSUBS 0.009276f
C467 B.n427 VSUBS 0.009276f
C468 B.n428 VSUBS 0.009276f
C469 B.n429 VSUBS 0.009276f
C470 B.n430 VSUBS 0.009276f
C471 B.n431 VSUBS 0.009276f
C472 B.n432 VSUBS 0.009276f
C473 B.n433 VSUBS 0.009276f
C474 B.n434 VSUBS 0.009276f
C475 B.n435 VSUBS 0.009276f
C476 B.n436 VSUBS 0.009276f
C477 B.n437 VSUBS 0.009276f
C478 B.n438 VSUBS 0.009276f
C479 B.n439 VSUBS 0.009276f
C480 B.n440 VSUBS 0.009276f
C481 B.n441 VSUBS 0.009276f
C482 B.n442 VSUBS 0.009276f
C483 B.n443 VSUBS 0.009276f
C484 B.n444 VSUBS 0.009276f
C485 B.n445 VSUBS 0.009276f
C486 B.n446 VSUBS 0.009276f
C487 B.n447 VSUBS 0.009276f
C488 B.n448 VSUBS 0.009276f
C489 B.n449 VSUBS 0.009276f
C490 B.n450 VSUBS 0.009276f
C491 B.n451 VSUBS 0.009276f
C492 B.n452 VSUBS 0.009276f
C493 B.n453 VSUBS 0.009276f
C494 B.n454 VSUBS 0.009276f
C495 B.n455 VSUBS 0.009276f
C496 B.n456 VSUBS 0.009276f
C497 B.n457 VSUBS 0.009276f
C498 B.n458 VSUBS 0.009276f
C499 B.n459 VSUBS 0.009276f
C500 B.n460 VSUBS 0.009276f
C501 B.n461 VSUBS 0.009276f
C502 B.n462 VSUBS 0.009276f
C503 B.n463 VSUBS 0.009276f
C504 B.n464 VSUBS 0.009276f
C505 B.n465 VSUBS 0.009276f
C506 B.n466 VSUBS 0.009276f
C507 B.n467 VSUBS 0.009276f
C508 B.n468 VSUBS 0.009276f
C509 B.n469 VSUBS 0.009276f
C510 B.n470 VSUBS 0.009276f
C511 B.n471 VSUBS 0.009276f
C512 B.n472 VSUBS 0.009276f
C513 B.n473 VSUBS 0.009276f
C514 B.n474 VSUBS 0.020815f
C515 B.n475 VSUBS 0.019601f
C516 B.n476 VSUBS 0.021051f
C517 B.n477 VSUBS 0.009276f
C518 B.n478 VSUBS 0.009276f
C519 B.n479 VSUBS 0.009276f
C520 B.n480 VSUBS 0.009276f
C521 B.n481 VSUBS 0.009276f
C522 B.n482 VSUBS 0.009276f
C523 B.n483 VSUBS 0.009276f
C524 B.n484 VSUBS 0.009276f
C525 B.n485 VSUBS 0.009276f
C526 B.n486 VSUBS 0.009276f
C527 B.n487 VSUBS 0.009276f
C528 B.n488 VSUBS 0.009276f
C529 B.n489 VSUBS 0.009276f
C530 B.n490 VSUBS 0.009276f
C531 B.n491 VSUBS 0.009276f
C532 B.n492 VSUBS 0.009276f
C533 B.n493 VSUBS 0.009276f
C534 B.n494 VSUBS 0.009276f
C535 B.n495 VSUBS 0.009276f
C536 B.n496 VSUBS 0.009276f
C537 B.n497 VSUBS 0.009276f
C538 B.n498 VSUBS 0.008731f
C539 B.n499 VSUBS 0.009276f
C540 B.n500 VSUBS 0.009276f
C541 B.n501 VSUBS 0.009276f
C542 B.n502 VSUBS 0.009276f
C543 B.n503 VSUBS 0.009276f
C544 B.n504 VSUBS 0.009276f
C545 B.n505 VSUBS 0.009276f
C546 B.n506 VSUBS 0.009276f
C547 B.n507 VSUBS 0.009276f
C548 B.n508 VSUBS 0.009276f
C549 B.n509 VSUBS 0.009276f
C550 B.n510 VSUBS 0.009276f
C551 B.n511 VSUBS 0.009276f
C552 B.n512 VSUBS 0.009276f
C553 B.n513 VSUBS 0.009276f
C554 B.n514 VSUBS 0.005184f
C555 B.n515 VSUBS 0.021493f
C556 B.n516 VSUBS 0.008731f
C557 B.n517 VSUBS 0.009276f
C558 B.n518 VSUBS 0.009276f
C559 B.n519 VSUBS 0.009276f
C560 B.n520 VSUBS 0.009276f
C561 B.n521 VSUBS 0.009276f
C562 B.n522 VSUBS 0.009276f
C563 B.n523 VSUBS 0.009276f
C564 B.n524 VSUBS 0.009276f
C565 B.n525 VSUBS 0.009276f
C566 B.n526 VSUBS 0.009276f
C567 B.n527 VSUBS 0.009276f
C568 B.n528 VSUBS 0.009276f
C569 B.n529 VSUBS 0.009276f
C570 B.n530 VSUBS 0.009276f
C571 B.n531 VSUBS 0.009276f
C572 B.n532 VSUBS 0.009276f
C573 B.n533 VSUBS 0.009276f
C574 B.n534 VSUBS 0.009276f
C575 B.n535 VSUBS 0.009276f
C576 B.n536 VSUBS 0.009276f
C577 B.n537 VSUBS 0.009276f
C578 B.n538 VSUBS 0.021051f
C579 B.n539 VSUBS 0.021051f
C580 B.n540 VSUBS 0.019601f
C581 B.n541 VSUBS 0.009276f
C582 B.n542 VSUBS 0.009276f
C583 B.n543 VSUBS 0.009276f
C584 B.n544 VSUBS 0.009276f
C585 B.n545 VSUBS 0.009276f
C586 B.n546 VSUBS 0.009276f
C587 B.n547 VSUBS 0.009276f
C588 B.n548 VSUBS 0.009276f
C589 B.n549 VSUBS 0.009276f
C590 B.n550 VSUBS 0.009276f
C591 B.n551 VSUBS 0.009276f
C592 B.n552 VSUBS 0.009276f
C593 B.n553 VSUBS 0.009276f
C594 B.n554 VSUBS 0.009276f
C595 B.n555 VSUBS 0.009276f
C596 B.n556 VSUBS 0.009276f
C597 B.n557 VSUBS 0.009276f
C598 B.n558 VSUBS 0.009276f
C599 B.n559 VSUBS 0.009276f
C600 B.n560 VSUBS 0.009276f
C601 B.n561 VSUBS 0.009276f
C602 B.n562 VSUBS 0.009276f
C603 B.n563 VSUBS 0.009276f
C604 B.n564 VSUBS 0.009276f
C605 B.n565 VSUBS 0.009276f
C606 B.n566 VSUBS 0.009276f
C607 B.n567 VSUBS 0.009276f
C608 B.n568 VSUBS 0.009276f
C609 B.n569 VSUBS 0.009276f
C610 B.n570 VSUBS 0.009276f
C611 B.n571 VSUBS 0.009276f
C612 B.n572 VSUBS 0.009276f
C613 B.n573 VSUBS 0.009276f
C614 B.n574 VSUBS 0.009276f
C615 B.n575 VSUBS 0.009276f
C616 B.n576 VSUBS 0.009276f
C617 B.n577 VSUBS 0.009276f
C618 B.n578 VSUBS 0.009276f
C619 B.n579 VSUBS 0.009276f
C620 B.n580 VSUBS 0.009276f
C621 B.n581 VSUBS 0.009276f
C622 B.n582 VSUBS 0.009276f
C623 B.n583 VSUBS 0.009276f
C624 B.n584 VSUBS 0.009276f
C625 B.n585 VSUBS 0.009276f
C626 B.n586 VSUBS 0.009276f
C627 B.n587 VSUBS 0.009276f
C628 B.n588 VSUBS 0.009276f
C629 B.n589 VSUBS 0.009276f
C630 B.n590 VSUBS 0.009276f
C631 B.n591 VSUBS 0.009276f
C632 B.n592 VSUBS 0.009276f
C633 B.n593 VSUBS 0.009276f
C634 B.n594 VSUBS 0.009276f
C635 B.n595 VSUBS 0.009276f
C636 B.n596 VSUBS 0.009276f
C637 B.n597 VSUBS 0.009276f
C638 B.n598 VSUBS 0.009276f
C639 B.n599 VSUBS 0.009276f
C640 B.n600 VSUBS 0.009276f
C641 B.n601 VSUBS 0.009276f
C642 B.n602 VSUBS 0.009276f
C643 B.n603 VSUBS 0.009276f
C644 B.n604 VSUBS 0.009276f
C645 B.n605 VSUBS 0.009276f
C646 B.n606 VSUBS 0.009276f
C647 B.n607 VSUBS 0.009276f
C648 B.n608 VSUBS 0.009276f
C649 B.n609 VSUBS 0.009276f
C650 B.n610 VSUBS 0.009276f
C651 B.n611 VSUBS 0.009276f
C652 B.n612 VSUBS 0.009276f
C653 B.n613 VSUBS 0.009276f
C654 B.n614 VSUBS 0.009276f
C655 B.n615 VSUBS 0.009276f
C656 B.n616 VSUBS 0.009276f
C657 B.n617 VSUBS 0.009276f
C658 B.n618 VSUBS 0.009276f
C659 B.n619 VSUBS 0.009276f
C660 B.n620 VSUBS 0.009276f
C661 B.n621 VSUBS 0.009276f
C662 B.n622 VSUBS 0.009276f
C663 B.n623 VSUBS 0.021005f
C664 VDD1.n0 VSUBS 0.025327f
C665 VDD1.n1 VSUBS 0.023048f
C666 VDD1.n2 VSUBS 0.012385f
C667 VDD1.n3 VSUBS 0.021956f
C668 VDD1.n4 VSUBS 0.018073f
C669 VDD1.t1 VSUBS 0.06618f
C670 VDD1.n5 VSUBS 0.085296f
C671 VDD1.n6 VSUBS 0.240367f
C672 VDD1.n7 VSUBS 0.012385f
C673 VDD1.n8 VSUBS 0.013114f
C674 VDD1.n9 VSUBS 0.029274f
C675 VDD1.n10 VSUBS 0.070874f
C676 VDD1.n11 VSUBS 0.013114f
C677 VDD1.n12 VSUBS 0.012385f
C678 VDD1.n13 VSUBS 0.058628f
C679 VDD1.n14 VSUBS 0.063341f
C680 VDD1.n15 VSUBS 0.025327f
C681 VDD1.n16 VSUBS 0.023048f
C682 VDD1.n17 VSUBS 0.012385f
C683 VDD1.n18 VSUBS 0.021956f
C684 VDD1.n19 VSUBS 0.018073f
C685 VDD1.t2 VSUBS 0.06618f
C686 VDD1.n20 VSUBS 0.085296f
C687 VDD1.n21 VSUBS 0.240367f
C688 VDD1.n22 VSUBS 0.012385f
C689 VDD1.n23 VSUBS 0.013114f
C690 VDD1.n24 VSUBS 0.029274f
C691 VDD1.n25 VSUBS 0.070874f
C692 VDD1.n26 VSUBS 0.013114f
C693 VDD1.n27 VSUBS 0.012385f
C694 VDD1.n28 VSUBS 0.058628f
C695 VDD1.n29 VSUBS 0.062482f
C696 VDD1.t5 VSUBS 0.059923f
C697 VDD1.t3 VSUBS 0.059923f
C698 VDD1.n30 VSUBS 0.329586f
C699 VDD1.n31 VSUBS 2.64983f
C700 VDD1.t4 VSUBS 0.059923f
C701 VDD1.t0 VSUBS 0.059923f
C702 VDD1.n32 VSUBS 0.325771f
C703 VDD1.n33 VSUBS 2.33846f
C704 VP.t2 VSUBS 1.47069f
C705 VP.n0 VSUBS 0.78909f
C706 VP.n1 VSUBS 0.048628f
C707 VP.n2 VSUBS 0.072343f
C708 VP.n3 VSUBS 0.048628f
C709 VP.n4 VSUBS 0.068258f
C710 VP.n5 VSUBS 0.048628f
C711 VP.n6 VSUBS 0.069633f
C712 VP.n7 VSUBS 0.048628f
C713 VP.n8 VSUBS 0.066468f
C714 VP.t5 VSUBS 1.47069f
C715 VP.n9 VSUBS 0.78909f
C716 VP.n10 VSUBS 0.048628f
C717 VP.n11 VSUBS 0.072343f
C718 VP.n12 VSUBS 0.048628f
C719 VP.n13 VSUBS 0.068258f
C720 VP.t4 VSUBS 2.05708f
C721 VP.t1 VSUBS 1.47069f
C722 VP.n14 VSUBS 0.760284f
C723 VP.n15 VSUBS 0.772437f
C724 VP.n16 VSUBS 0.60833f
C725 VP.n17 VSUBS 0.048628f
C726 VP.n18 VSUBS 0.09063f
C727 VP.n19 VSUBS 0.09063f
C728 VP.n20 VSUBS 0.069633f
C729 VP.n21 VSUBS 0.048628f
C730 VP.n22 VSUBS 0.048628f
C731 VP.n23 VSUBS 0.048628f
C732 VP.n24 VSUBS 0.09063f
C733 VP.n25 VSUBS 0.09063f
C734 VP.n26 VSUBS 0.066468f
C735 VP.n27 VSUBS 0.078485f
C736 VP.n28 VSUBS 2.49306f
C737 VP.t3 VSUBS 1.47069f
C738 VP.n29 VSUBS 0.78909f
C739 VP.n30 VSUBS 2.53078f
C740 VP.n31 VSUBS 0.078485f
C741 VP.n32 VSUBS 0.048628f
C742 VP.n33 VSUBS 0.09063f
C743 VP.n34 VSUBS 0.09063f
C744 VP.n35 VSUBS 0.072343f
C745 VP.n36 VSUBS 0.048628f
C746 VP.n37 VSUBS 0.048628f
C747 VP.n38 VSUBS 0.048628f
C748 VP.n39 VSUBS 0.09063f
C749 VP.n40 VSUBS 0.09063f
C750 VP.t0 VSUBS 1.47069f
C751 VP.n41 VSUBS 0.590244f
C752 VP.n42 VSUBS 0.068258f
C753 VP.n43 VSUBS 0.048628f
C754 VP.n44 VSUBS 0.048628f
C755 VP.n45 VSUBS 0.048628f
C756 VP.n46 VSUBS 0.09063f
C757 VP.n47 VSUBS 0.09063f
C758 VP.n48 VSUBS 0.069633f
C759 VP.n49 VSUBS 0.048628f
C760 VP.n50 VSUBS 0.048628f
C761 VP.n51 VSUBS 0.048628f
C762 VP.n52 VSUBS 0.09063f
C763 VP.n53 VSUBS 0.09063f
C764 VP.n54 VSUBS 0.066468f
C765 VP.n55 VSUBS 0.078485f
C766 VP.n56 VSUBS 0.131714f
C767 VTAIL.t9 VSUBS 0.084312f
C768 VTAIL.t10 VSUBS 0.084312f
C769 VTAIL.n0 VSUBS 0.397133f
C770 VTAIL.n1 VSUBS 0.767615f
C771 VTAIL.n2 VSUBS 0.035635f
C772 VTAIL.n3 VSUBS 0.032429f
C773 VTAIL.n4 VSUBS 0.017426f
C774 VTAIL.n5 VSUBS 0.030892f
C775 VTAIL.n6 VSUBS 0.025429f
C776 VTAIL.t1 VSUBS 0.093116f
C777 VTAIL.n7 VSUBS 0.120012f
C778 VTAIL.n8 VSUBS 0.338199f
C779 VTAIL.n9 VSUBS 0.017426f
C780 VTAIL.n10 VSUBS 0.018451f
C781 VTAIL.n11 VSUBS 0.041189f
C782 VTAIL.n12 VSUBS 0.099721f
C783 VTAIL.n13 VSUBS 0.018451f
C784 VTAIL.n14 VSUBS 0.017426f
C785 VTAIL.n15 VSUBS 0.08249f
C786 VTAIL.n16 VSUBS 0.050371f
C787 VTAIL.n17 VSUBS 0.618839f
C788 VTAIL.t2 VSUBS 0.084312f
C789 VTAIL.t0 VSUBS 0.084312f
C790 VTAIL.n18 VSUBS 0.397133f
C791 VTAIL.n19 VSUBS 2.256f
C792 VTAIL.t7 VSUBS 0.084312f
C793 VTAIL.t8 VSUBS 0.084312f
C794 VTAIL.n20 VSUBS 0.397135f
C795 VTAIL.n21 VSUBS 2.256f
C796 VTAIL.n22 VSUBS 0.035635f
C797 VTAIL.n23 VSUBS 0.032429f
C798 VTAIL.n24 VSUBS 0.017426f
C799 VTAIL.n25 VSUBS 0.030892f
C800 VTAIL.n26 VSUBS 0.025429f
C801 VTAIL.t5 VSUBS 0.093116f
C802 VTAIL.n27 VSUBS 0.120012f
C803 VTAIL.n28 VSUBS 0.338199f
C804 VTAIL.n29 VSUBS 0.017426f
C805 VTAIL.n30 VSUBS 0.018451f
C806 VTAIL.n31 VSUBS 0.041189f
C807 VTAIL.n32 VSUBS 0.099721f
C808 VTAIL.n33 VSUBS 0.018451f
C809 VTAIL.n34 VSUBS 0.017426f
C810 VTAIL.n35 VSUBS 0.08249f
C811 VTAIL.n36 VSUBS 0.050371f
C812 VTAIL.n37 VSUBS 0.618839f
C813 VTAIL.t4 VSUBS 0.084312f
C814 VTAIL.t11 VSUBS 0.084312f
C815 VTAIL.n38 VSUBS 0.397135f
C816 VTAIL.n39 VSUBS 1.03043f
C817 VTAIL.n40 VSUBS 0.035635f
C818 VTAIL.n41 VSUBS 0.032429f
C819 VTAIL.n42 VSUBS 0.017426f
C820 VTAIL.n43 VSUBS 0.030892f
C821 VTAIL.n44 VSUBS 0.025429f
C822 VTAIL.t3 VSUBS 0.093116f
C823 VTAIL.n45 VSUBS 0.120012f
C824 VTAIL.n46 VSUBS 0.338199f
C825 VTAIL.n47 VSUBS 0.017426f
C826 VTAIL.n48 VSUBS 0.018451f
C827 VTAIL.n49 VSUBS 0.041189f
C828 VTAIL.n50 VSUBS 0.099721f
C829 VTAIL.n51 VSUBS 0.018451f
C830 VTAIL.n52 VSUBS 0.017426f
C831 VTAIL.n53 VSUBS 0.08249f
C832 VTAIL.n54 VSUBS 0.050371f
C833 VTAIL.n55 VSUBS 1.48589f
C834 VTAIL.n56 VSUBS 0.035635f
C835 VTAIL.n57 VSUBS 0.032429f
C836 VTAIL.n58 VSUBS 0.017426f
C837 VTAIL.n59 VSUBS 0.030892f
C838 VTAIL.n60 VSUBS 0.025429f
C839 VTAIL.t6 VSUBS 0.093116f
C840 VTAIL.n61 VSUBS 0.120012f
C841 VTAIL.n62 VSUBS 0.338199f
C842 VTAIL.n63 VSUBS 0.017426f
C843 VTAIL.n64 VSUBS 0.018451f
C844 VTAIL.n65 VSUBS 0.041189f
C845 VTAIL.n66 VSUBS 0.099721f
C846 VTAIL.n67 VSUBS 0.018451f
C847 VTAIL.n68 VSUBS 0.017426f
C848 VTAIL.n69 VSUBS 0.08249f
C849 VTAIL.n70 VSUBS 0.050371f
C850 VTAIL.n71 VSUBS 1.39018f
C851 VDD2.n0 VSUBS 0.031112f
C852 VDD2.n1 VSUBS 0.028313f
C853 VDD2.n2 VSUBS 0.015214f
C854 VDD2.n3 VSUBS 0.026971f
C855 VDD2.n4 VSUBS 0.022201f
C856 VDD2.t4 VSUBS 0.081298f
C857 VDD2.n5 VSUBS 0.10478f
C858 VDD2.n6 VSUBS 0.295274f
C859 VDD2.n7 VSUBS 0.015214f
C860 VDD2.n8 VSUBS 0.016109f
C861 VDD2.n9 VSUBS 0.035961f
C862 VDD2.n10 VSUBS 0.087064f
C863 VDD2.n11 VSUBS 0.016109f
C864 VDD2.n12 VSUBS 0.015214f
C865 VDD2.n13 VSUBS 0.07202f
C866 VDD2.n14 VSUBS 0.076755f
C867 VDD2.t3 VSUBS 0.073611f
C868 VDD2.t2 VSUBS 0.073611f
C869 VDD2.n15 VSUBS 0.404872f
C870 VDD2.n16 VSUBS 3.09457f
C871 VDD2.n17 VSUBS 0.031112f
C872 VDD2.n18 VSUBS 0.028313f
C873 VDD2.n19 VSUBS 0.015214f
C874 VDD2.n20 VSUBS 0.026971f
C875 VDD2.n21 VSUBS 0.022201f
C876 VDD2.t5 VSUBS 0.081298f
C877 VDD2.n22 VSUBS 0.10478f
C878 VDD2.n23 VSUBS 0.295274f
C879 VDD2.n24 VSUBS 0.015214f
C880 VDD2.n25 VSUBS 0.016109f
C881 VDD2.n26 VSUBS 0.035961f
C882 VDD2.n27 VSUBS 0.087064f
C883 VDD2.n28 VSUBS 0.016109f
C884 VDD2.n29 VSUBS 0.015214f
C885 VDD2.n30 VSUBS 0.07202f
C886 VDD2.n31 VSUBS 0.063481f
C887 VDD2.n32 VSUBS 2.45731f
C888 VDD2.t0 VSUBS 0.073611f
C889 VDD2.t1 VSUBS 0.073611f
C890 VDD2.n33 VSUBS 0.404849f
C891 VN.t4 VSUBS 1.26782f
C892 VN.n0 VSUBS 0.68024f
C893 VN.n1 VSUBS 0.04192f
C894 VN.n2 VSUBS 0.062364f
C895 VN.n3 VSUBS 0.04192f
C896 VN.n4 VSUBS 0.058842f
C897 VN.t0 VSUBS 1.26782f
C898 VN.n5 VSUBS 0.655407f
C899 VN.t1 VSUBS 1.77332f
C900 VN.n6 VSUBS 0.665883f
C901 VN.n7 VSUBS 0.524413f
C902 VN.n8 VSUBS 0.04192f
C903 VN.n9 VSUBS 0.078128f
C904 VN.n10 VSUBS 0.078128f
C905 VN.n11 VSUBS 0.060027f
C906 VN.n12 VSUBS 0.04192f
C907 VN.n13 VSUBS 0.04192f
C908 VN.n14 VSUBS 0.04192f
C909 VN.n15 VSUBS 0.078128f
C910 VN.n16 VSUBS 0.078128f
C911 VN.n17 VSUBS 0.057299f
C912 VN.n18 VSUBS 0.067658f
C913 VN.n19 VSUBS 0.113544f
C914 VN.t3 VSUBS 1.26782f
C915 VN.n20 VSUBS 0.68024f
C916 VN.n21 VSUBS 0.04192f
C917 VN.n22 VSUBS 0.062364f
C918 VN.n23 VSUBS 0.04192f
C919 VN.n24 VSUBS 0.058842f
C920 VN.t5 VSUBS 1.77332f
C921 VN.t2 VSUBS 1.26782f
C922 VN.n25 VSUBS 0.655407f
C923 VN.n26 VSUBS 0.665883f
C924 VN.n27 VSUBS 0.524413f
C925 VN.n28 VSUBS 0.04192f
C926 VN.n29 VSUBS 0.078128f
C927 VN.n30 VSUBS 0.078128f
C928 VN.n31 VSUBS 0.060027f
C929 VN.n32 VSUBS 0.04192f
C930 VN.n33 VSUBS 0.04192f
C931 VN.n34 VSUBS 0.04192f
C932 VN.n35 VSUBS 0.078128f
C933 VN.n36 VSUBS 0.078128f
C934 VN.n37 VSUBS 0.057299f
C935 VN.n38 VSUBS 0.067658f
C936 VN.n39 VSUBS 2.16675f
.ends

