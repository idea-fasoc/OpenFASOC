* NGSPICE file created from diff_pair_sample_0815.ext - technology: sky130A

.subckt diff_pair_sample_0815 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t5 VN.t0 VTAIL.t11 w_n4194_n4126# sky130_fd_pr__pfet_01v8 ad=2.60535 pd=16.12 as=6.1581 ps=32.36 w=15.79 l=3.7
X1 VTAIL.t6 VN.t1 VDD2.t4 w_n4194_n4126# sky130_fd_pr__pfet_01v8 ad=2.60535 pd=16.12 as=2.60535 ps=16.12 w=15.79 l=3.7
X2 VDD1.t5 VP.t0 VTAIL.t1 w_n4194_n4126# sky130_fd_pr__pfet_01v8 ad=2.60535 pd=16.12 as=6.1581 ps=32.36 w=15.79 l=3.7
X3 VDD1.t4 VP.t1 VTAIL.t5 w_n4194_n4126# sky130_fd_pr__pfet_01v8 ad=6.1581 pd=32.36 as=2.60535 ps=16.12 w=15.79 l=3.7
X4 VTAIL.t4 VP.t2 VDD1.t3 w_n4194_n4126# sky130_fd_pr__pfet_01v8 ad=2.60535 pd=16.12 as=2.60535 ps=16.12 w=15.79 l=3.7
X5 VDD1.t2 VP.t3 VTAIL.t3 w_n4194_n4126# sky130_fd_pr__pfet_01v8 ad=6.1581 pd=32.36 as=2.60535 ps=16.12 w=15.79 l=3.7
X6 B.t11 B.t9 B.t10 w_n4194_n4126# sky130_fd_pr__pfet_01v8 ad=6.1581 pd=32.36 as=0 ps=0 w=15.79 l=3.7
X7 VDD2.t3 VN.t2 VTAIL.t7 w_n4194_n4126# sky130_fd_pr__pfet_01v8 ad=2.60535 pd=16.12 as=6.1581 ps=32.36 w=15.79 l=3.7
X8 VDD2.t2 VN.t3 VTAIL.t8 w_n4194_n4126# sky130_fd_pr__pfet_01v8 ad=6.1581 pd=32.36 as=2.60535 ps=16.12 w=15.79 l=3.7
X9 B.t8 B.t6 B.t7 w_n4194_n4126# sky130_fd_pr__pfet_01v8 ad=6.1581 pd=32.36 as=0 ps=0 w=15.79 l=3.7
X10 B.t5 B.t3 B.t4 w_n4194_n4126# sky130_fd_pr__pfet_01v8 ad=6.1581 pd=32.36 as=0 ps=0 w=15.79 l=3.7
X11 VTAIL.t0 VP.t4 VDD1.t1 w_n4194_n4126# sky130_fd_pr__pfet_01v8 ad=2.60535 pd=16.12 as=2.60535 ps=16.12 w=15.79 l=3.7
X12 B.t2 B.t0 B.t1 w_n4194_n4126# sky130_fd_pr__pfet_01v8 ad=6.1581 pd=32.36 as=0 ps=0 w=15.79 l=3.7
X13 VDD1.t0 VP.t5 VTAIL.t2 w_n4194_n4126# sky130_fd_pr__pfet_01v8 ad=2.60535 pd=16.12 as=6.1581 ps=32.36 w=15.79 l=3.7
X14 VDD2.t1 VN.t4 VTAIL.t9 w_n4194_n4126# sky130_fd_pr__pfet_01v8 ad=6.1581 pd=32.36 as=2.60535 ps=16.12 w=15.79 l=3.7
X15 VTAIL.t10 VN.t5 VDD2.t0 w_n4194_n4126# sky130_fd_pr__pfet_01v8 ad=2.60535 pd=16.12 as=2.60535 ps=16.12 w=15.79 l=3.7
R0 VN.n38 VN.n37 161.3
R1 VN.n36 VN.n21 161.3
R2 VN.n35 VN.n34 161.3
R3 VN.n33 VN.n22 161.3
R4 VN.n32 VN.n31 161.3
R5 VN.n30 VN.n23 161.3
R6 VN.n29 VN.n28 161.3
R7 VN.n27 VN.n24 161.3
R8 VN.n18 VN.n17 161.3
R9 VN.n16 VN.n1 161.3
R10 VN.n15 VN.n14 161.3
R11 VN.n13 VN.n2 161.3
R12 VN.n12 VN.n11 161.3
R13 VN.n10 VN.n3 161.3
R14 VN.n9 VN.n8 161.3
R15 VN.n7 VN.n4 161.3
R16 VN.n6 VN.t3 135.38
R17 VN.n26 VN.t2 135.38
R18 VN.n5 VN.t5 102.849
R19 VN.n0 VN.t0 102.849
R20 VN.n25 VN.t1 102.849
R21 VN.n20 VN.t4 102.849
R22 VN.n19 VN.n0 88.5994
R23 VN.n39 VN.n20 88.5994
R24 VN VN.n39 56.0321
R25 VN.n26 VN.n25 50.4814
R26 VN.n6 VN.n5 50.4814
R27 VN.n11 VN.n2 41.9503
R28 VN.n31 VN.n22 41.9503
R29 VN.n11 VN.n10 39.0365
R30 VN.n31 VN.n30 39.0365
R31 VN.n5 VN.n4 24.4675
R32 VN.n9 VN.n4 24.4675
R33 VN.n10 VN.n9 24.4675
R34 VN.n15 VN.n2 24.4675
R35 VN.n16 VN.n15 24.4675
R36 VN.n17 VN.n16 24.4675
R37 VN.n30 VN.n29 24.4675
R38 VN.n29 VN.n24 24.4675
R39 VN.n25 VN.n24 24.4675
R40 VN.n37 VN.n36 24.4675
R41 VN.n36 VN.n35 24.4675
R42 VN.n35 VN.n22 24.4675
R43 VN.n7 VN.n6 2.49445
R44 VN.n27 VN.n26 2.49445
R45 VN.n17 VN.n0 1.46852
R46 VN.n37 VN.n20 1.46852
R47 VN.n39 VN.n38 0.354971
R48 VN.n19 VN.n18 0.354971
R49 VN VN.n19 0.26696
R50 VN.n38 VN.n21 0.189894
R51 VN.n34 VN.n21 0.189894
R52 VN.n34 VN.n33 0.189894
R53 VN.n33 VN.n32 0.189894
R54 VN.n32 VN.n23 0.189894
R55 VN.n28 VN.n23 0.189894
R56 VN.n28 VN.n27 0.189894
R57 VN.n8 VN.n7 0.189894
R58 VN.n8 VN.n3 0.189894
R59 VN.n12 VN.n3 0.189894
R60 VN.n13 VN.n12 0.189894
R61 VN.n14 VN.n13 0.189894
R62 VN.n14 VN.n1 0.189894
R63 VN.n18 VN.n1 0.189894
R64 VTAIL.n7 VTAIL.t7 56.7611
R65 VTAIL.n10 VTAIL.t1 56.761
R66 VTAIL.n11 VTAIL.t11 56.7609
R67 VTAIL.n2 VTAIL.t2 56.7609
R68 VTAIL.n9 VTAIL.n8 54.7026
R69 VTAIL.n6 VTAIL.n5 54.7026
R70 VTAIL.n1 VTAIL.n0 54.7023
R71 VTAIL.n4 VTAIL.n3 54.7023
R72 VTAIL.n6 VTAIL.n4 32.9272
R73 VTAIL.n11 VTAIL.n10 29.4531
R74 VTAIL.n7 VTAIL.n6 3.47464
R75 VTAIL.n10 VTAIL.n9 3.47464
R76 VTAIL.n4 VTAIL.n2 3.47464
R77 VTAIL VTAIL.n11 2.54791
R78 VTAIL.n9 VTAIL.n7 2.2074
R79 VTAIL.n2 VTAIL.n1 2.2074
R80 VTAIL.n0 VTAIL.t8 2.05908
R81 VTAIL.n0 VTAIL.t10 2.05908
R82 VTAIL.n3 VTAIL.t3 2.05908
R83 VTAIL.n3 VTAIL.t4 2.05908
R84 VTAIL.n8 VTAIL.t5 2.05908
R85 VTAIL.n8 VTAIL.t0 2.05908
R86 VTAIL.n5 VTAIL.t9 2.05908
R87 VTAIL.n5 VTAIL.t6 2.05908
R88 VTAIL VTAIL.n1 0.927224
R89 VDD2.n1 VDD2.t2 75.99
R90 VDD2.n2 VDD2.t1 73.4399
R91 VDD2.n1 VDD2.n0 72.1943
R92 VDD2 VDD2.n3 72.1915
R93 VDD2.n2 VDD2.n1 48.6183
R94 VDD2 VDD2.n2 2.66429
R95 VDD2.n3 VDD2.t4 2.05908
R96 VDD2.n3 VDD2.t3 2.05908
R97 VDD2.n0 VDD2.t0 2.05908
R98 VDD2.n0 VDD2.t5 2.05908
R99 VP.n16 VP.n13 161.3
R100 VP.n18 VP.n17 161.3
R101 VP.n19 VP.n12 161.3
R102 VP.n21 VP.n20 161.3
R103 VP.n22 VP.n11 161.3
R104 VP.n24 VP.n23 161.3
R105 VP.n25 VP.n10 161.3
R106 VP.n27 VP.n26 161.3
R107 VP.n56 VP.n55 161.3
R108 VP.n54 VP.n1 161.3
R109 VP.n53 VP.n52 161.3
R110 VP.n51 VP.n2 161.3
R111 VP.n50 VP.n49 161.3
R112 VP.n48 VP.n3 161.3
R113 VP.n47 VP.n46 161.3
R114 VP.n45 VP.n4 161.3
R115 VP.n44 VP.n43 161.3
R116 VP.n42 VP.n5 161.3
R117 VP.n41 VP.n40 161.3
R118 VP.n39 VP.n6 161.3
R119 VP.n38 VP.n37 161.3
R120 VP.n36 VP.n7 161.3
R121 VP.n35 VP.n34 161.3
R122 VP.n33 VP.n8 161.3
R123 VP.n32 VP.n31 161.3
R124 VP.n15 VP.t1 135.38
R125 VP.n43 VP.t2 102.849
R126 VP.n30 VP.t3 102.849
R127 VP.n0 VP.t5 102.849
R128 VP.n14 VP.t4 102.849
R129 VP.n9 VP.t0 102.849
R130 VP.n30 VP.n29 88.5994
R131 VP.n57 VP.n0 88.5994
R132 VP.n28 VP.n9 88.5994
R133 VP.n29 VP.n28 55.8668
R134 VP.n15 VP.n14 50.4814
R135 VP.n37 VP.n36 41.9503
R136 VP.n49 VP.n2 41.9503
R137 VP.n20 VP.n11 41.9503
R138 VP.n37 VP.n6 39.0365
R139 VP.n49 VP.n48 39.0365
R140 VP.n20 VP.n19 39.0365
R141 VP.n31 VP.n8 24.4675
R142 VP.n35 VP.n8 24.4675
R143 VP.n36 VP.n35 24.4675
R144 VP.n41 VP.n6 24.4675
R145 VP.n42 VP.n41 24.4675
R146 VP.n43 VP.n42 24.4675
R147 VP.n43 VP.n4 24.4675
R148 VP.n47 VP.n4 24.4675
R149 VP.n48 VP.n47 24.4675
R150 VP.n53 VP.n2 24.4675
R151 VP.n54 VP.n53 24.4675
R152 VP.n55 VP.n54 24.4675
R153 VP.n24 VP.n11 24.4675
R154 VP.n25 VP.n24 24.4675
R155 VP.n26 VP.n25 24.4675
R156 VP.n14 VP.n13 24.4675
R157 VP.n18 VP.n13 24.4675
R158 VP.n19 VP.n18 24.4675
R159 VP.n16 VP.n15 2.49444
R160 VP.n31 VP.n30 1.46852
R161 VP.n55 VP.n0 1.46852
R162 VP.n26 VP.n9 1.46852
R163 VP.n28 VP.n27 0.354971
R164 VP.n32 VP.n29 0.354971
R165 VP.n57 VP.n56 0.354971
R166 VP VP.n57 0.26696
R167 VP.n17 VP.n16 0.189894
R168 VP.n17 VP.n12 0.189894
R169 VP.n21 VP.n12 0.189894
R170 VP.n22 VP.n21 0.189894
R171 VP.n23 VP.n22 0.189894
R172 VP.n23 VP.n10 0.189894
R173 VP.n27 VP.n10 0.189894
R174 VP.n33 VP.n32 0.189894
R175 VP.n34 VP.n33 0.189894
R176 VP.n34 VP.n7 0.189894
R177 VP.n38 VP.n7 0.189894
R178 VP.n39 VP.n38 0.189894
R179 VP.n40 VP.n39 0.189894
R180 VP.n40 VP.n5 0.189894
R181 VP.n44 VP.n5 0.189894
R182 VP.n45 VP.n44 0.189894
R183 VP.n46 VP.n45 0.189894
R184 VP.n46 VP.n3 0.189894
R185 VP.n50 VP.n3 0.189894
R186 VP.n51 VP.n50 0.189894
R187 VP.n52 VP.n51 0.189894
R188 VP.n52 VP.n1 0.189894
R189 VP.n56 VP.n1 0.189894
R190 VDD1 VDD1.t4 76.1036
R191 VDD1.n1 VDD1.t2 75.99
R192 VDD1.n1 VDD1.n0 72.1943
R193 VDD1.n3 VDD1.n2 71.3812
R194 VDD1.n3 VDD1.n1 50.9384
R195 VDD1.n2 VDD1.t1 2.05908
R196 VDD1.n2 VDD1.t5 2.05908
R197 VDD1.n0 VDD1.t3 2.05908
R198 VDD1.n0 VDD1.t0 2.05908
R199 VDD1 VDD1.n3 0.810845
R200 B.n491 B.n490 585
R201 B.n489 B.n148 585
R202 B.n488 B.n487 585
R203 B.n486 B.n149 585
R204 B.n485 B.n484 585
R205 B.n483 B.n150 585
R206 B.n482 B.n481 585
R207 B.n480 B.n151 585
R208 B.n479 B.n478 585
R209 B.n477 B.n152 585
R210 B.n476 B.n475 585
R211 B.n474 B.n153 585
R212 B.n473 B.n472 585
R213 B.n471 B.n154 585
R214 B.n470 B.n469 585
R215 B.n468 B.n155 585
R216 B.n467 B.n466 585
R217 B.n465 B.n156 585
R218 B.n464 B.n463 585
R219 B.n462 B.n157 585
R220 B.n461 B.n460 585
R221 B.n459 B.n158 585
R222 B.n458 B.n457 585
R223 B.n456 B.n159 585
R224 B.n455 B.n454 585
R225 B.n453 B.n160 585
R226 B.n452 B.n451 585
R227 B.n450 B.n161 585
R228 B.n449 B.n448 585
R229 B.n447 B.n162 585
R230 B.n446 B.n445 585
R231 B.n444 B.n163 585
R232 B.n443 B.n442 585
R233 B.n441 B.n164 585
R234 B.n440 B.n439 585
R235 B.n438 B.n165 585
R236 B.n437 B.n436 585
R237 B.n435 B.n166 585
R238 B.n434 B.n433 585
R239 B.n432 B.n167 585
R240 B.n431 B.n430 585
R241 B.n429 B.n168 585
R242 B.n428 B.n427 585
R243 B.n426 B.n169 585
R244 B.n425 B.n424 585
R245 B.n423 B.n170 585
R246 B.n422 B.n421 585
R247 B.n420 B.n171 585
R248 B.n419 B.n418 585
R249 B.n417 B.n172 585
R250 B.n416 B.n415 585
R251 B.n414 B.n173 585
R252 B.n413 B.n412 585
R253 B.n411 B.n410 585
R254 B.n409 B.n177 585
R255 B.n408 B.n407 585
R256 B.n406 B.n178 585
R257 B.n405 B.n404 585
R258 B.n403 B.n179 585
R259 B.n402 B.n401 585
R260 B.n400 B.n180 585
R261 B.n399 B.n398 585
R262 B.n396 B.n181 585
R263 B.n395 B.n394 585
R264 B.n393 B.n184 585
R265 B.n392 B.n391 585
R266 B.n390 B.n185 585
R267 B.n389 B.n388 585
R268 B.n387 B.n186 585
R269 B.n386 B.n385 585
R270 B.n384 B.n187 585
R271 B.n383 B.n382 585
R272 B.n381 B.n188 585
R273 B.n380 B.n379 585
R274 B.n378 B.n189 585
R275 B.n377 B.n376 585
R276 B.n375 B.n190 585
R277 B.n374 B.n373 585
R278 B.n372 B.n191 585
R279 B.n371 B.n370 585
R280 B.n369 B.n192 585
R281 B.n368 B.n367 585
R282 B.n366 B.n193 585
R283 B.n365 B.n364 585
R284 B.n363 B.n194 585
R285 B.n362 B.n361 585
R286 B.n360 B.n195 585
R287 B.n359 B.n358 585
R288 B.n357 B.n196 585
R289 B.n356 B.n355 585
R290 B.n354 B.n197 585
R291 B.n353 B.n352 585
R292 B.n351 B.n198 585
R293 B.n350 B.n349 585
R294 B.n348 B.n199 585
R295 B.n347 B.n346 585
R296 B.n345 B.n200 585
R297 B.n344 B.n343 585
R298 B.n342 B.n201 585
R299 B.n341 B.n340 585
R300 B.n339 B.n202 585
R301 B.n338 B.n337 585
R302 B.n336 B.n203 585
R303 B.n335 B.n334 585
R304 B.n333 B.n204 585
R305 B.n332 B.n331 585
R306 B.n330 B.n205 585
R307 B.n329 B.n328 585
R308 B.n327 B.n206 585
R309 B.n326 B.n325 585
R310 B.n324 B.n207 585
R311 B.n323 B.n322 585
R312 B.n321 B.n208 585
R313 B.n320 B.n319 585
R314 B.n318 B.n209 585
R315 B.n492 B.n147 585
R316 B.n494 B.n493 585
R317 B.n495 B.n146 585
R318 B.n497 B.n496 585
R319 B.n498 B.n145 585
R320 B.n500 B.n499 585
R321 B.n501 B.n144 585
R322 B.n503 B.n502 585
R323 B.n504 B.n143 585
R324 B.n506 B.n505 585
R325 B.n507 B.n142 585
R326 B.n509 B.n508 585
R327 B.n510 B.n141 585
R328 B.n512 B.n511 585
R329 B.n513 B.n140 585
R330 B.n515 B.n514 585
R331 B.n516 B.n139 585
R332 B.n518 B.n517 585
R333 B.n519 B.n138 585
R334 B.n521 B.n520 585
R335 B.n522 B.n137 585
R336 B.n524 B.n523 585
R337 B.n525 B.n136 585
R338 B.n527 B.n526 585
R339 B.n528 B.n135 585
R340 B.n530 B.n529 585
R341 B.n531 B.n134 585
R342 B.n533 B.n532 585
R343 B.n534 B.n133 585
R344 B.n536 B.n535 585
R345 B.n537 B.n132 585
R346 B.n539 B.n538 585
R347 B.n540 B.n131 585
R348 B.n542 B.n541 585
R349 B.n543 B.n130 585
R350 B.n545 B.n544 585
R351 B.n546 B.n129 585
R352 B.n548 B.n547 585
R353 B.n549 B.n128 585
R354 B.n551 B.n550 585
R355 B.n552 B.n127 585
R356 B.n554 B.n553 585
R357 B.n555 B.n126 585
R358 B.n557 B.n556 585
R359 B.n558 B.n125 585
R360 B.n560 B.n559 585
R361 B.n561 B.n124 585
R362 B.n563 B.n562 585
R363 B.n564 B.n123 585
R364 B.n566 B.n565 585
R365 B.n567 B.n122 585
R366 B.n569 B.n568 585
R367 B.n570 B.n121 585
R368 B.n572 B.n571 585
R369 B.n573 B.n120 585
R370 B.n575 B.n574 585
R371 B.n576 B.n119 585
R372 B.n578 B.n577 585
R373 B.n579 B.n118 585
R374 B.n581 B.n580 585
R375 B.n582 B.n117 585
R376 B.n584 B.n583 585
R377 B.n585 B.n116 585
R378 B.n587 B.n586 585
R379 B.n588 B.n115 585
R380 B.n590 B.n589 585
R381 B.n591 B.n114 585
R382 B.n593 B.n592 585
R383 B.n594 B.n113 585
R384 B.n596 B.n595 585
R385 B.n597 B.n112 585
R386 B.n599 B.n598 585
R387 B.n600 B.n111 585
R388 B.n602 B.n601 585
R389 B.n603 B.n110 585
R390 B.n605 B.n604 585
R391 B.n606 B.n109 585
R392 B.n608 B.n607 585
R393 B.n609 B.n108 585
R394 B.n611 B.n610 585
R395 B.n612 B.n107 585
R396 B.n614 B.n613 585
R397 B.n615 B.n106 585
R398 B.n617 B.n616 585
R399 B.n618 B.n105 585
R400 B.n620 B.n619 585
R401 B.n621 B.n104 585
R402 B.n623 B.n622 585
R403 B.n624 B.n103 585
R404 B.n626 B.n625 585
R405 B.n627 B.n102 585
R406 B.n629 B.n628 585
R407 B.n630 B.n101 585
R408 B.n632 B.n631 585
R409 B.n633 B.n100 585
R410 B.n635 B.n634 585
R411 B.n636 B.n99 585
R412 B.n638 B.n637 585
R413 B.n639 B.n98 585
R414 B.n641 B.n640 585
R415 B.n642 B.n97 585
R416 B.n644 B.n643 585
R417 B.n645 B.n96 585
R418 B.n647 B.n646 585
R419 B.n648 B.n95 585
R420 B.n650 B.n649 585
R421 B.n651 B.n94 585
R422 B.n653 B.n652 585
R423 B.n654 B.n93 585
R424 B.n656 B.n655 585
R425 B.n657 B.n92 585
R426 B.n659 B.n658 585
R427 B.n833 B.n832 585
R428 B.n831 B.n30 585
R429 B.n830 B.n829 585
R430 B.n828 B.n31 585
R431 B.n827 B.n826 585
R432 B.n825 B.n32 585
R433 B.n824 B.n823 585
R434 B.n822 B.n33 585
R435 B.n821 B.n820 585
R436 B.n819 B.n34 585
R437 B.n818 B.n817 585
R438 B.n816 B.n35 585
R439 B.n815 B.n814 585
R440 B.n813 B.n36 585
R441 B.n812 B.n811 585
R442 B.n810 B.n37 585
R443 B.n809 B.n808 585
R444 B.n807 B.n38 585
R445 B.n806 B.n805 585
R446 B.n804 B.n39 585
R447 B.n803 B.n802 585
R448 B.n801 B.n40 585
R449 B.n800 B.n799 585
R450 B.n798 B.n41 585
R451 B.n797 B.n796 585
R452 B.n795 B.n42 585
R453 B.n794 B.n793 585
R454 B.n792 B.n43 585
R455 B.n791 B.n790 585
R456 B.n789 B.n44 585
R457 B.n788 B.n787 585
R458 B.n786 B.n45 585
R459 B.n785 B.n784 585
R460 B.n783 B.n46 585
R461 B.n782 B.n781 585
R462 B.n780 B.n47 585
R463 B.n779 B.n778 585
R464 B.n777 B.n48 585
R465 B.n776 B.n775 585
R466 B.n774 B.n49 585
R467 B.n773 B.n772 585
R468 B.n771 B.n50 585
R469 B.n770 B.n769 585
R470 B.n768 B.n51 585
R471 B.n767 B.n766 585
R472 B.n765 B.n52 585
R473 B.n764 B.n763 585
R474 B.n762 B.n53 585
R475 B.n761 B.n760 585
R476 B.n759 B.n54 585
R477 B.n758 B.n757 585
R478 B.n756 B.n55 585
R479 B.n755 B.n754 585
R480 B.n753 B.n752 585
R481 B.n751 B.n59 585
R482 B.n750 B.n749 585
R483 B.n748 B.n60 585
R484 B.n747 B.n746 585
R485 B.n745 B.n61 585
R486 B.n744 B.n743 585
R487 B.n742 B.n62 585
R488 B.n741 B.n740 585
R489 B.n738 B.n63 585
R490 B.n737 B.n736 585
R491 B.n735 B.n66 585
R492 B.n734 B.n733 585
R493 B.n732 B.n67 585
R494 B.n731 B.n730 585
R495 B.n729 B.n68 585
R496 B.n728 B.n727 585
R497 B.n726 B.n69 585
R498 B.n725 B.n724 585
R499 B.n723 B.n70 585
R500 B.n722 B.n721 585
R501 B.n720 B.n71 585
R502 B.n719 B.n718 585
R503 B.n717 B.n72 585
R504 B.n716 B.n715 585
R505 B.n714 B.n73 585
R506 B.n713 B.n712 585
R507 B.n711 B.n74 585
R508 B.n710 B.n709 585
R509 B.n708 B.n75 585
R510 B.n707 B.n706 585
R511 B.n705 B.n76 585
R512 B.n704 B.n703 585
R513 B.n702 B.n77 585
R514 B.n701 B.n700 585
R515 B.n699 B.n78 585
R516 B.n698 B.n697 585
R517 B.n696 B.n79 585
R518 B.n695 B.n694 585
R519 B.n693 B.n80 585
R520 B.n692 B.n691 585
R521 B.n690 B.n81 585
R522 B.n689 B.n688 585
R523 B.n687 B.n82 585
R524 B.n686 B.n685 585
R525 B.n684 B.n83 585
R526 B.n683 B.n682 585
R527 B.n681 B.n84 585
R528 B.n680 B.n679 585
R529 B.n678 B.n85 585
R530 B.n677 B.n676 585
R531 B.n675 B.n86 585
R532 B.n674 B.n673 585
R533 B.n672 B.n87 585
R534 B.n671 B.n670 585
R535 B.n669 B.n88 585
R536 B.n668 B.n667 585
R537 B.n666 B.n89 585
R538 B.n665 B.n664 585
R539 B.n663 B.n90 585
R540 B.n662 B.n661 585
R541 B.n660 B.n91 585
R542 B.n834 B.n29 585
R543 B.n836 B.n835 585
R544 B.n837 B.n28 585
R545 B.n839 B.n838 585
R546 B.n840 B.n27 585
R547 B.n842 B.n841 585
R548 B.n843 B.n26 585
R549 B.n845 B.n844 585
R550 B.n846 B.n25 585
R551 B.n848 B.n847 585
R552 B.n849 B.n24 585
R553 B.n851 B.n850 585
R554 B.n852 B.n23 585
R555 B.n854 B.n853 585
R556 B.n855 B.n22 585
R557 B.n857 B.n856 585
R558 B.n858 B.n21 585
R559 B.n860 B.n859 585
R560 B.n861 B.n20 585
R561 B.n863 B.n862 585
R562 B.n864 B.n19 585
R563 B.n866 B.n865 585
R564 B.n867 B.n18 585
R565 B.n869 B.n868 585
R566 B.n870 B.n17 585
R567 B.n872 B.n871 585
R568 B.n873 B.n16 585
R569 B.n875 B.n874 585
R570 B.n876 B.n15 585
R571 B.n878 B.n877 585
R572 B.n879 B.n14 585
R573 B.n881 B.n880 585
R574 B.n882 B.n13 585
R575 B.n884 B.n883 585
R576 B.n885 B.n12 585
R577 B.n887 B.n886 585
R578 B.n888 B.n11 585
R579 B.n890 B.n889 585
R580 B.n891 B.n10 585
R581 B.n893 B.n892 585
R582 B.n894 B.n9 585
R583 B.n896 B.n895 585
R584 B.n897 B.n8 585
R585 B.n899 B.n898 585
R586 B.n900 B.n7 585
R587 B.n902 B.n901 585
R588 B.n903 B.n6 585
R589 B.n905 B.n904 585
R590 B.n906 B.n5 585
R591 B.n908 B.n907 585
R592 B.n909 B.n4 585
R593 B.n911 B.n910 585
R594 B.n912 B.n3 585
R595 B.n914 B.n913 585
R596 B.n915 B.n0 585
R597 B.n2 B.n1 585
R598 B.n237 B.n236 585
R599 B.n239 B.n238 585
R600 B.n240 B.n235 585
R601 B.n242 B.n241 585
R602 B.n243 B.n234 585
R603 B.n245 B.n244 585
R604 B.n246 B.n233 585
R605 B.n248 B.n247 585
R606 B.n249 B.n232 585
R607 B.n251 B.n250 585
R608 B.n252 B.n231 585
R609 B.n254 B.n253 585
R610 B.n255 B.n230 585
R611 B.n257 B.n256 585
R612 B.n258 B.n229 585
R613 B.n260 B.n259 585
R614 B.n261 B.n228 585
R615 B.n263 B.n262 585
R616 B.n264 B.n227 585
R617 B.n266 B.n265 585
R618 B.n267 B.n226 585
R619 B.n269 B.n268 585
R620 B.n270 B.n225 585
R621 B.n272 B.n271 585
R622 B.n273 B.n224 585
R623 B.n275 B.n274 585
R624 B.n276 B.n223 585
R625 B.n278 B.n277 585
R626 B.n279 B.n222 585
R627 B.n281 B.n280 585
R628 B.n282 B.n221 585
R629 B.n284 B.n283 585
R630 B.n285 B.n220 585
R631 B.n287 B.n286 585
R632 B.n288 B.n219 585
R633 B.n290 B.n289 585
R634 B.n291 B.n218 585
R635 B.n293 B.n292 585
R636 B.n294 B.n217 585
R637 B.n296 B.n295 585
R638 B.n297 B.n216 585
R639 B.n299 B.n298 585
R640 B.n300 B.n215 585
R641 B.n302 B.n301 585
R642 B.n303 B.n214 585
R643 B.n305 B.n304 585
R644 B.n306 B.n213 585
R645 B.n308 B.n307 585
R646 B.n309 B.n212 585
R647 B.n311 B.n310 585
R648 B.n312 B.n211 585
R649 B.n314 B.n313 585
R650 B.n315 B.n210 585
R651 B.n317 B.n316 585
R652 B.n316 B.n209 511.721
R653 B.n490 B.n147 511.721
R654 B.n658 B.n91 511.721
R655 B.n832 B.n29 511.721
R656 B.n182 B.t9 312.113
R657 B.n174 B.t3 312.113
R658 B.n64 B.t6 312.113
R659 B.n56 B.t0 312.113
R660 B.n917 B.n916 256.663
R661 B.n916 B.n915 235.042
R662 B.n916 B.n2 235.042
R663 B.n174 B.t4 187.52
R664 B.n64 B.t8 187.52
R665 B.n182 B.t10 187.5
R666 B.n56 B.t2 187.5
R667 B.n320 B.n209 163.367
R668 B.n321 B.n320 163.367
R669 B.n322 B.n321 163.367
R670 B.n322 B.n207 163.367
R671 B.n326 B.n207 163.367
R672 B.n327 B.n326 163.367
R673 B.n328 B.n327 163.367
R674 B.n328 B.n205 163.367
R675 B.n332 B.n205 163.367
R676 B.n333 B.n332 163.367
R677 B.n334 B.n333 163.367
R678 B.n334 B.n203 163.367
R679 B.n338 B.n203 163.367
R680 B.n339 B.n338 163.367
R681 B.n340 B.n339 163.367
R682 B.n340 B.n201 163.367
R683 B.n344 B.n201 163.367
R684 B.n345 B.n344 163.367
R685 B.n346 B.n345 163.367
R686 B.n346 B.n199 163.367
R687 B.n350 B.n199 163.367
R688 B.n351 B.n350 163.367
R689 B.n352 B.n351 163.367
R690 B.n352 B.n197 163.367
R691 B.n356 B.n197 163.367
R692 B.n357 B.n356 163.367
R693 B.n358 B.n357 163.367
R694 B.n358 B.n195 163.367
R695 B.n362 B.n195 163.367
R696 B.n363 B.n362 163.367
R697 B.n364 B.n363 163.367
R698 B.n364 B.n193 163.367
R699 B.n368 B.n193 163.367
R700 B.n369 B.n368 163.367
R701 B.n370 B.n369 163.367
R702 B.n370 B.n191 163.367
R703 B.n374 B.n191 163.367
R704 B.n375 B.n374 163.367
R705 B.n376 B.n375 163.367
R706 B.n376 B.n189 163.367
R707 B.n380 B.n189 163.367
R708 B.n381 B.n380 163.367
R709 B.n382 B.n381 163.367
R710 B.n382 B.n187 163.367
R711 B.n386 B.n187 163.367
R712 B.n387 B.n386 163.367
R713 B.n388 B.n387 163.367
R714 B.n388 B.n185 163.367
R715 B.n392 B.n185 163.367
R716 B.n393 B.n392 163.367
R717 B.n394 B.n393 163.367
R718 B.n394 B.n181 163.367
R719 B.n399 B.n181 163.367
R720 B.n400 B.n399 163.367
R721 B.n401 B.n400 163.367
R722 B.n401 B.n179 163.367
R723 B.n405 B.n179 163.367
R724 B.n406 B.n405 163.367
R725 B.n407 B.n406 163.367
R726 B.n407 B.n177 163.367
R727 B.n411 B.n177 163.367
R728 B.n412 B.n411 163.367
R729 B.n412 B.n173 163.367
R730 B.n416 B.n173 163.367
R731 B.n417 B.n416 163.367
R732 B.n418 B.n417 163.367
R733 B.n418 B.n171 163.367
R734 B.n422 B.n171 163.367
R735 B.n423 B.n422 163.367
R736 B.n424 B.n423 163.367
R737 B.n424 B.n169 163.367
R738 B.n428 B.n169 163.367
R739 B.n429 B.n428 163.367
R740 B.n430 B.n429 163.367
R741 B.n430 B.n167 163.367
R742 B.n434 B.n167 163.367
R743 B.n435 B.n434 163.367
R744 B.n436 B.n435 163.367
R745 B.n436 B.n165 163.367
R746 B.n440 B.n165 163.367
R747 B.n441 B.n440 163.367
R748 B.n442 B.n441 163.367
R749 B.n442 B.n163 163.367
R750 B.n446 B.n163 163.367
R751 B.n447 B.n446 163.367
R752 B.n448 B.n447 163.367
R753 B.n448 B.n161 163.367
R754 B.n452 B.n161 163.367
R755 B.n453 B.n452 163.367
R756 B.n454 B.n453 163.367
R757 B.n454 B.n159 163.367
R758 B.n458 B.n159 163.367
R759 B.n459 B.n458 163.367
R760 B.n460 B.n459 163.367
R761 B.n460 B.n157 163.367
R762 B.n464 B.n157 163.367
R763 B.n465 B.n464 163.367
R764 B.n466 B.n465 163.367
R765 B.n466 B.n155 163.367
R766 B.n470 B.n155 163.367
R767 B.n471 B.n470 163.367
R768 B.n472 B.n471 163.367
R769 B.n472 B.n153 163.367
R770 B.n476 B.n153 163.367
R771 B.n477 B.n476 163.367
R772 B.n478 B.n477 163.367
R773 B.n478 B.n151 163.367
R774 B.n482 B.n151 163.367
R775 B.n483 B.n482 163.367
R776 B.n484 B.n483 163.367
R777 B.n484 B.n149 163.367
R778 B.n488 B.n149 163.367
R779 B.n489 B.n488 163.367
R780 B.n490 B.n489 163.367
R781 B.n658 B.n657 163.367
R782 B.n657 B.n656 163.367
R783 B.n656 B.n93 163.367
R784 B.n652 B.n93 163.367
R785 B.n652 B.n651 163.367
R786 B.n651 B.n650 163.367
R787 B.n650 B.n95 163.367
R788 B.n646 B.n95 163.367
R789 B.n646 B.n645 163.367
R790 B.n645 B.n644 163.367
R791 B.n644 B.n97 163.367
R792 B.n640 B.n97 163.367
R793 B.n640 B.n639 163.367
R794 B.n639 B.n638 163.367
R795 B.n638 B.n99 163.367
R796 B.n634 B.n99 163.367
R797 B.n634 B.n633 163.367
R798 B.n633 B.n632 163.367
R799 B.n632 B.n101 163.367
R800 B.n628 B.n101 163.367
R801 B.n628 B.n627 163.367
R802 B.n627 B.n626 163.367
R803 B.n626 B.n103 163.367
R804 B.n622 B.n103 163.367
R805 B.n622 B.n621 163.367
R806 B.n621 B.n620 163.367
R807 B.n620 B.n105 163.367
R808 B.n616 B.n105 163.367
R809 B.n616 B.n615 163.367
R810 B.n615 B.n614 163.367
R811 B.n614 B.n107 163.367
R812 B.n610 B.n107 163.367
R813 B.n610 B.n609 163.367
R814 B.n609 B.n608 163.367
R815 B.n608 B.n109 163.367
R816 B.n604 B.n109 163.367
R817 B.n604 B.n603 163.367
R818 B.n603 B.n602 163.367
R819 B.n602 B.n111 163.367
R820 B.n598 B.n111 163.367
R821 B.n598 B.n597 163.367
R822 B.n597 B.n596 163.367
R823 B.n596 B.n113 163.367
R824 B.n592 B.n113 163.367
R825 B.n592 B.n591 163.367
R826 B.n591 B.n590 163.367
R827 B.n590 B.n115 163.367
R828 B.n586 B.n115 163.367
R829 B.n586 B.n585 163.367
R830 B.n585 B.n584 163.367
R831 B.n584 B.n117 163.367
R832 B.n580 B.n117 163.367
R833 B.n580 B.n579 163.367
R834 B.n579 B.n578 163.367
R835 B.n578 B.n119 163.367
R836 B.n574 B.n119 163.367
R837 B.n574 B.n573 163.367
R838 B.n573 B.n572 163.367
R839 B.n572 B.n121 163.367
R840 B.n568 B.n121 163.367
R841 B.n568 B.n567 163.367
R842 B.n567 B.n566 163.367
R843 B.n566 B.n123 163.367
R844 B.n562 B.n123 163.367
R845 B.n562 B.n561 163.367
R846 B.n561 B.n560 163.367
R847 B.n560 B.n125 163.367
R848 B.n556 B.n125 163.367
R849 B.n556 B.n555 163.367
R850 B.n555 B.n554 163.367
R851 B.n554 B.n127 163.367
R852 B.n550 B.n127 163.367
R853 B.n550 B.n549 163.367
R854 B.n549 B.n548 163.367
R855 B.n548 B.n129 163.367
R856 B.n544 B.n129 163.367
R857 B.n544 B.n543 163.367
R858 B.n543 B.n542 163.367
R859 B.n542 B.n131 163.367
R860 B.n538 B.n131 163.367
R861 B.n538 B.n537 163.367
R862 B.n537 B.n536 163.367
R863 B.n536 B.n133 163.367
R864 B.n532 B.n133 163.367
R865 B.n532 B.n531 163.367
R866 B.n531 B.n530 163.367
R867 B.n530 B.n135 163.367
R868 B.n526 B.n135 163.367
R869 B.n526 B.n525 163.367
R870 B.n525 B.n524 163.367
R871 B.n524 B.n137 163.367
R872 B.n520 B.n137 163.367
R873 B.n520 B.n519 163.367
R874 B.n519 B.n518 163.367
R875 B.n518 B.n139 163.367
R876 B.n514 B.n139 163.367
R877 B.n514 B.n513 163.367
R878 B.n513 B.n512 163.367
R879 B.n512 B.n141 163.367
R880 B.n508 B.n141 163.367
R881 B.n508 B.n507 163.367
R882 B.n507 B.n506 163.367
R883 B.n506 B.n143 163.367
R884 B.n502 B.n143 163.367
R885 B.n502 B.n501 163.367
R886 B.n501 B.n500 163.367
R887 B.n500 B.n145 163.367
R888 B.n496 B.n145 163.367
R889 B.n496 B.n495 163.367
R890 B.n495 B.n494 163.367
R891 B.n494 B.n147 163.367
R892 B.n832 B.n831 163.367
R893 B.n831 B.n830 163.367
R894 B.n830 B.n31 163.367
R895 B.n826 B.n31 163.367
R896 B.n826 B.n825 163.367
R897 B.n825 B.n824 163.367
R898 B.n824 B.n33 163.367
R899 B.n820 B.n33 163.367
R900 B.n820 B.n819 163.367
R901 B.n819 B.n818 163.367
R902 B.n818 B.n35 163.367
R903 B.n814 B.n35 163.367
R904 B.n814 B.n813 163.367
R905 B.n813 B.n812 163.367
R906 B.n812 B.n37 163.367
R907 B.n808 B.n37 163.367
R908 B.n808 B.n807 163.367
R909 B.n807 B.n806 163.367
R910 B.n806 B.n39 163.367
R911 B.n802 B.n39 163.367
R912 B.n802 B.n801 163.367
R913 B.n801 B.n800 163.367
R914 B.n800 B.n41 163.367
R915 B.n796 B.n41 163.367
R916 B.n796 B.n795 163.367
R917 B.n795 B.n794 163.367
R918 B.n794 B.n43 163.367
R919 B.n790 B.n43 163.367
R920 B.n790 B.n789 163.367
R921 B.n789 B.n788 163.367
R922 B.n788 B.n45 163.367
R923 B.n784 B.n45 163.367
R924 B.n784 B.n783 163.367
R925 B.n783 B.n782 163.367
R926 B.n782 B.n47 163.367
R927 B.n778 B.n47 163.367
R928 B.n778 B.n777 163.367
R929 B.n777 B.n776 163.367
R930 B.n776 B.n49 163.367
R931 B.n772 B.n49 163.367
R932 B.n772 B.n771 163.367
R933 B.n771 B.n770 163.367
R934 B.n770 B.n51 163.367
R935 B.n766 B.n51 163.367
R936 B.n766 B.n765 163.367
R937 B.n765 B.n764 163.367
R938 B.n764 B.n53 163.367
R939 B.n760 B.n53 163.367
R940 B.n760 B.n759 163.367
R941 B.n759 B.n758 163.367
R942 B.n758 B.n55 163.367
R943 B.n754 B.n55 163.367
R944 B.n754 B.n753 163.367
R945 B.n753 B.n59 163.367
R946 B.n749 B.n59 163.367
R947 B.n749 B.n748 163.367
R948 B.n748 B.n747 163.367
R949 B.n747 B.n61 163.367
R950 B.n743 B.n61 163.367
R951 B.n743 B.n742 163.367
R952 B.n742 B.n741 163.367
R953 B.n741 B.n63 163.367
R954 B.n736 B.n63 163.367
R955 B.n736 B.n735 163.367
R956 B.n735 B.n734 163.367
R957 B.n734 B.n67 163.367
R958 B.n730 B.n67 163.367
R959 B.n730 B.n729 163.367
R960 B.n729 B.n728 163.367
R961 B.n728 B.n69 163.367
R962 B.n724 B.n69 163.367
R963 B.n724 B.n723 163.367
R964 B.n723 B.n722 163.367
R965 B.n722 B.n71 163.367
R966 B.n718 B.n71 163.367
R967 B.n718 B.n717 163.367
R968 B.n717 B.n716 163.367
R969 B.n716 B.n73 163.367
R970 B.n712 B.n73 163.367
R971 B.n712 B.n711 163.367
R972 B.n711 B.n710 163.367
R973 B.n710 B.n75 163.367
R974 B.n706 B.n75 163.367
R975 B.n706 B.n705 163.367
R976 B.n705 B.n704 163.367
R977 B.n704 B.n77 163.367
R978 B.n700 B.n77 163.367
R979 B.n700 B.n699 163.367
R980 B.n699 B.n698 163.367
R981 B.n698 B.n79 163.367
R982 B.n694 B.n79 163.367
R983 B.n694 B.n693 163.367
R984 B.n693 B.n692 163.367
R985 B.n692 B.n81 163.367
R986 B.n688 B.n81 163.367
R987 B.n688 B.n687 163.367
R988 B.n687 B.n686 163.367
R989 B.n686 B.n83 163.367
R990 B.n682 B.n83 163.367
R991 B.n682 B.n681 163.367
R992 B.n681 B.n680 163.367
R993 B.n680 B.n85 163.367
R994 B.n676 B.n85 163.367
R995 B.n676 B.n675 163.367
R996 B.n675 B.n674 163.367
R997 B.n674 B.n87 163.367
R998 B.n670 B.n87 163.367
R999 B.n670 B.n669 163.367
R1000 B.n669 B.n668 163.367
R1001 B.n668 B.n89 163.367
R1002 B.n664 B.n89 163.367
R1003 B.n664 B.n663 163.367
R1004 B.n663 B.n662 163.367
R1005 B.n662 B.n91 163.367
R1006 B.n836 B.n29 163.367
R1007 B.n837 B.n836 163.367
R1008 B.n838 B.n837 163.367
R1009 B.n838 B.n27 163.367
R1010 B.n842 B.n27 163.367
R1011 B.n843 B.n842 163.367
R1012 B.n844 B.n843 163.367
R1013 B.n844 B.n25 163.367
R1014 B.n848 B.n25 163.367
R1015 B.n849 B.n848 163.367
R1016 B.n850 B.n849 163.367
R1017 B.n850 B.n23 163.367
R1018 B.n854 B.n23 163.367
R1019 B.n855 B.n854 163.367
R1020 B.n856 B.n855 163.367
R1021 B.n856 B.n21 163.367
R1022 B.n860 B.n21 163.367
R1023 B.n861 B.n860 163.367
R1024 B.n862 B.n861 163.367
R1025 B.n862 B.n19 163.367
R1026 B.n866 B.n19 163.367
R1027 B.n867 B.n866 163.367
R1028 B.n868 B.n867 163.367
R1029 B.n868 B.n17 163.367
R1030 B.n872 B.n17 163.367
R1031 B.n873 B.n872 163.367
R1032 B.n874 B.n873 163.367
R1033 B.n874 B.n15 163.367
R1034 B.n878 B.n15 163.367
R1035 B.n879 B.n878 163.367
R1036 B.n880 B.n879 163.367
R1037 B.n880 B.n13 163.367
R1038 B.n884 B.n13 163.367
R1039 B.n885 B.n884 163.367
R1040 B.n886 B.n885 163.367
R1041 B.n886 B.n11 163.367
R1042 B.n890 B.n11 163.367
R1043 B.n891 B.n890 163.367
R1044 B.n892 B.n891 163.367
R1045 B.n892 B.n9 163.367
R1046 B.n896 B.n9 163.367
R1047 B.n897 B.n896 163.367
R1048 B.n898 B.n897 163.367
R1049 B.n898 B.n7 163.367
R1050 B.n902 B.n7 163.367
R1051 B.n903 B.n902 163.367
R1052 B.n904 B.n903 163.367
R1053 B.n904 B.n5 163.367
R1054 B.n908 B.n5 163.367
R1055 B.n909 B.n908 163.367
R1056 B.n910 B.n909 163.367
R1057 B.n910 B.n3 163.367
R1058 B.n914 B.n3 163.367
R1059 B.n915 B.n914 163.367
R1060 B.n237 B.n2 163.367
R1061 B.n238 B.n237 163.367
R1062 B.n238 B.n235 163.367
R1063 B.n242 B.n235 163.367
R1064 B.n243 B.n242 163.367
R1065 B.n244 B.n243 163.367
R1066 B.n244 B.n233 163.367
R1067 B.n248 B.n233 163.367
R1068 B.n249 B.n248 163.367
R1069 B.n250 B.n249 163.367
R1070 B.n250 B.n231 163.367
R1071 B.n254 B.n231 163.367
R1072 B.n255 B.n254 163.367
R1073 B.n256 B.n255 163.367
R1074 B.n256 B.n229 163.367
R1075 B.n260 B.n229 163.367
R1076 B.n261 B.n260 163.367
R1077 B.n262 B.n261 163.367
R1078 B.n262 B.n227 163.367
R1079 B.n266 B.n227 163.367
R1080 B.n267 B.n266 163.367
R1081 B.n268 B.n267 163.367
R1082 B.n268 B.n225 163.367
R1083 B.n272 B.n225 163.367
R1084 B.n273 B.n272 163.367
R1085 B.n274 B.n273 163.367
R1086 B.n274 B.n223 163.367
R1087 B.n278 B.n223 163.367
R1088 B.n279 B.n278 163.367
R1089 B.n280 B.n279 163.367
R1090 B.n280 B.n221 163.367
R1091 B.n284 B.n221 163.367
R1092 B.n285 B.n284 163.367
R1093 B.n286 B.n285 163.367
R1094 B.n286 B.n219 163.367
R1095 B.n290 B.n219 163.367
R1096 B.n291 B.n290 163.367
R1097 B.n292 B.n291 163.367
R1098 B.n292 B.n217 163.367
R1099 B.n296 B.n217 163.367
R1100 B.n297 B.n296 163.367
R1101 B.n298 B.n297 163.367
R1102 B.n298 B.n215 163.367
R1103 B.n302 B.n215 163.367
R1104 B.n303 B.n302 163.367
R1105 B.n304 B.n303 163.367
R1106 B.n304 B.n213 163.367
R1107 B.n308 B.n213 163.367
R1108 B.n309 B.n308 163.367
R1109 B.n310 B.n309 163.367
R1110 B.n310 B.n211 163.367
R1111 B.n314 B.n211 163.367
R1112 B.n315 B.n314 163.367
R1113 B.n316 B.n315 163.367
R1114 B.n175 B.t5 109.362
R1115 B.n65 B.t7 109.362
R1116 B.n183 B.t11 109.343
R1117 B.n57 B.t1 109.343
R1118 B.n183 B.n182 78.1581
R1119 B.n175 B.n174 78.1581
R1120 B.n65 B.n64 78.1581
R1121 B.n57 B.n56 78.1581
R1122 B.n397 B.n183 59.5399
R1123 B.n176 B.n175 59.5399
R1124 B.n739 B.n65 59.5399
R1125 B.n58 B.n57 59.5399
R1126 B.n834 B.n833 33.2493
R1127 B.n660 B.n659 33.2493
R1128 B.n492 B.n491 33.2493
R1129 B.n318 B.n317 33.2493
R1130 B B.n917 18.0485
R1131 B.n835 B.n834 10.6151
R1132 B.n835 B.n28 10.6151
R1133 B.n839 B.n28 10.6151
R1134 B.n840 B.n839 10.6151
R1135 B.n841 B.n840 10.6151
R1136 B.n841 B.n26 10.6151
R1137 B.n845 B.n26 10.6151
R1138 B.n846 B.n845 10.6151
R1139 B.n847 B.n846 10.6151
R1140 B.n847 B.n24 10.6151
R1141 B.n851 B.n24 10.6151
R1142 B.n852 B.n851 10.6151
R1143 B.n853 B.n852 10.6151
R1144 B.n853 B.n22 10.6151
R1145 B.n857 B.n22 10.6151
R1146 B.n858 B.n857 10.6151
R1147 B.n859 B.n858 10.6151
R1148 B.n859 B.n20 10.6151
R1149 B.n863 B.n20 10.6151
R1150 B.n864 B.n863 10.6151
R1151 B.n865 B.n864 10.6151
R1152 B.n865 B.n18 10.6151
R1153 B.n869 B.n18 10.6151
R1154 B.n870 B.n869 10.6151
R1155 B.n871 B.n870 10.6151
R1156 B.n871 B.n16 10.6151
R1157 B.n875 B.n16 10.6151
R1158 B.n876 B.n875 10.6151
R1159 B.n877 B.n876 10.6151
R1160 B.n877 B.n14 10.6151
R1161 B.n881 B.n14 10.6151
R1162 B.n882 B.n881 10.6151
R1163 B.n883 B.n882 10.6151
R1164 B.n883 B.n12 10.6151
R1165 B.n887 B.n12 10.6151
R1166 B.n888 B.n887 10.6151
R1167 B.n889 B.n888 10.6151
R1168 B.n889 B.n10 10.6151
R1169 B.n893 B.n10 10.6151
R1170 B.n894 B.n893 10.6151
R1171 B.n895 B.n894 10.6151
R1172 B.n895 B.n8 10.6151
R1173 B.n899 B.n8 10.6151
R1174 B.n900 B.n899 10.6151
R1175 B.n901 B.n900 10.6151
R1176 B.n901 B.n6 10.6151
R1177 B.n905 B.n6 10.6151
R1178 B.n906 B.n905 10.6151
R1179 B.n907 B.n906 10.6151
R1180 B.n907 B.n4 10.6151
R1181 B.n911 B.n4 10.6151
R1182 B.n912 B.n911 10.6151
R1183 B.n913 B.n912 10.6151
R1184 B.n913 B.n0 10.6151
R1185 B.n833 B.n30 10.6151
R1186 B.n829 B.n30 10.6151
R1187 B.n829 B.n828 10.6151
R1188 B.n828 B.n827 10.6151
R1189 B.n827 B.n32 10.6151
R1190 B.n823 B.n32 10.6151
R1191 B.n823 B.n822 10.6151
R1192 B.n822 B.n821 10.6151
R1193 B.n821 B.n34 10.6151
R1194 B.n817 B.n34 10.6151
R1195 B.n817 B.n816 10.6151
R1196 B.n816 B.n815 10.6151
R1197 B.n815 B.n36 10.6151
R1198 B.n811 B.n36 10.6151
R1199 B.n811 B.n810 10.6151
R1200 B.n810 B.n809 10.6151
R1201 B.n809 B.n38 10.6151
R1202 B.n805 B.n38 10.6151
R1203 B.n805 B.n804 10.6151
R1204 B.n804 B.n803 10.6151
R1205 B.n803 B.n40 10.6151
R1206 B.n799 B.n40 10.6151
R1207 B.n799 B.n798 10.6151
R1208 B.n798 B.n797 10.6151
R1209 B.n797 B.n42 10.6151
R1210 B.n793 B.n42 10.6151
R1211 B.n793 B.n792 10.6151
R1212 B.n792 B.n791 10.6151
R1213 B.n791 B.n44 10.6151
R1214 B.n787 B.n44 10.6151
R1215 B.n787 B.n786 10.6151
R1216 B.n786 B.n785 10.6151
R1217 B.n785 B.n46 10.6151
R1218 B.n781 B.n46 10.6151
R1219 B.n781 B.n780 10.6151
R1220 B.n780 B.n779 10.6151
R1221 B.n779 B.n48 10.6151
R1222 B.n775 B.n48 10.6151
R1223 B.n775 B.n774 10.6151
R1224 B.n774 B.n773 10.6151
R1225 B.n773 B.n50 10.6151
R1226 B.n769 B.n50 10.6151
R1227 B.n769 B.n768 10.6151
R1228 B.n768 B.n767 10.6151
R1229 B.n767 B.n52 10.6151
R1230 B.n763 B.n52 10.6151
R1231 B.n763 B.n762 10.6151
R1232 B.n762 B.n761 10.6151
R1233 B.n761 B.n54 10.6151
R1234 B.n757 B.n54 10.6151
R1235 B.n757 B.n756 10.6151
R1236 B.n756 B.n755 10.6151
R1237 B.n752 B.n751 10.6151
R1238 B.n751 B.n750 10.6151
R1239 B.n750 B.n60 10.6151
R1240 B.n746 B.n60 10.6151
R1241 B.n746 B.n745 10.6151
R1242 B.n745 B.n744 10.6151
R1243 B.n744 B.n62 10.6151
R1244 B.n740 B.n62 10.6151
R1245 B.n738 B.n737 10.6151
R1246 B.n737 B.n66 10.6151
R1247 B.n733 B.n66 10.6151
R1248 B.n733 B.n732 10.6151
R1249 B.n732 B.n731 10.6151
R1250 B.n731 B.n68 10.6151
R1251 B.n727 B.n68 10.6151
R1252 B.n727 B.n726 10.6151
R1253 B.n726 B.n725 10.6151
R1254 B.n725 B.n70 10.6151
R1255 B.n721 B.n70 10.6151
R1256 B.n721 B.n720 10.6151
R1257 B.n720 B.n719 10.6151
R1258 B.n719 B.n72 10.6151
R1259 B.n715 B.n72 10.6151
R1260 B.n715 B.n714 10.6151
R1261 B.n714 B.n713 10.6151
R1262 B.n713 B.n74 10.6151
R1263 B.n709 B.n74 10.6151
R1264 B.n709 B.n708 10.6151
R1265 B.n708 B.n707 10.6151
R1266 B.n707 B.n76 10.6151
R1267 B.n703 B.n76 10.6151
R1268 B.n703 B.n702 10.6151
R1269 B.n702 B.n701 10.6151
R1270 B.n701 B.n78 10.6151
R1271 B.n697 B.n78 10.6151
R1272 B.n697 B.n696 10.6151
R1273 B.n696 B.n695 10.6151
R1274 B.n695 B.n80 10.6151
R1275 B.n691 B.n80 10.6151
R1276 B.n691 B.n690 10.6151
R1277 B.n690 B.n689 10.6151
R1278 B.n689 B.n82 10.6151
R1279 B.n685 B.n82 10.6151
R1280 B.n685 B.n684 10.6151
R1281 B.n684 B.n683 10.6151
R1282 B.n683 B.n84 10.6151
R1283 B.n679 B.n84 10.6151
R1284 B.n679 B.n678 10.6151
R1285 B.n678 B.n677 10.6151
R1286 B.n677 B.n86 10.6151
R1287 B.n673 B.n86 10.6151
R1288 B.n673 B.n672 10.6151
R1289 B.n672 B.n671 10.6151
R1290 B.n671 B.n88 10.6151
R1291 B.n667 B.n88 10.6151
R1292 B.n667 B.n666 10.6151
R1293 B.n666 B.n665 10.6151
R1294 B.n665 B.n90 10.6151
R1295 B.n661 B.n90 10.6151
R1296 B.n661 B.n660 10.6151
R1297 B.n659 B.n92 10.6151
R1298 B.n655 B.n92 10.6151
R1299 B.n655 B.n654 10.6151
R1300 B.n654 B.n653 10.6151
R1301 B.n653 B.n94 10.6151
R1302 B.n649 B.n94 10.6151
R1303 B.n649 B.n648 10.6151
R1304 B.n648 B.n647 10.6151
R1305 B.n647 B.n96 10.6151
R1306 B.n643 B.n96 10.6151
R1307 B.n643 B.n642 10.6151
R1308 B.n642 B.n641 10.6151
R1309 B.n641 B.n98 10.6151
R1310 B.n637 B.n98 10.6151
R1311 B.n637 B.n636 10.6151
R1312 B.n636 B.n635 10.6151
R1313 B.n635 B.n100 10.6151
R1314 B.n631 B.n100 10.6151
R1315 B.n631 B.n630 10.6151
R1316 B.n630 B.n629 10.6151
R1317 B.n629 B.n102 10.6151
R1318 B.n625 B.n102 10.6151
R1319 B.n625 B.n624 10.6151
R1320 B.n624 B.n623 10.6151
R1321 B.n623 B.n104 10.6151
R1322 B.n619 B.n104 10.6151
R1323 B.n619 B.n618 10.6151
R1324 B.n618 B.n617 10.6151
R1325 B.n617 B.n106 10.6151
R1326 B.n613 B.n106 10.6151
R1327 B.n613 B.n612 10.6151
R1328 B.n612 B.n611 10.6151
R1329 B.n611 B.n108 10.6151
R1330 B.n607 B.n108 10.6151
R1331 B.n607 B.n606 10.6151
R1332 B.n606 B.n605 10.6151
R1333 B.n605 B.n110 10.6151
R1334 B.n601 B.n110 10.6151
R1335 B.n601 B.n600 10.6151
R1336 B.n600 B.n599 10.6151
R1337 B.n599 B.n112 10.6151
R1338 B.n595 B.n112 10.6151
R1339 B.n595 B.n594 10.6151
R1340 B.n594 B.n593 10.6151
R1341 B.n593 B.n114 10.6151
R1342 B.n589 B.n114 10.6151
R1343 B.n589 B.n588 10.6151
R1344 B.n588 B.n587 10.6151
R1345 B.n587 B.n116 10.6151
R1346 B.n583 B.n116 10.6151
R1347 B.n583 B.n582 10.6151
R1348 B.n582 B.n581 10.6151
R1349 B.n581 B.n118 10.6151
R1350 B.n577 B.n118 10.6151
R1351 B.n577 B.n576 10.6151
R1352 B.n576 B.n575 10.6151
R1353 B.n575 B.n120 10.6151
R1354 B.n571 B.n120 10.6151
R1355 B.n571 B.n570 10.6151
R1356 B.n570 B.n569 10.6151
R1357 B.n569 B.n122 10.6151
R1358 B.n565 B.n122 10.6151
R1359 B.n565 B.n564 10.6151
R1360 B.n564 B.n563 10.6151
R1361 B.n563 B.n124 10.6151
R1362 B.n559 B.n124 10.6151
R1363 B.n559 B.n558 10.6151
R1364 B.n558 B.n557 10.6151
R1365 B.n557 B.n126 10.6151
R1366 B.n553 B.n126 10.6151
R1367 B.n553 B.n552 10.6151
R1368 B.n552 B.n551 10.6151
R1369 B.n551 B.n128 10.6151
R1370 B.n547 B.n128 10.6151
R1371 B.n547 B.n546 10.6151
R1372 B.n546 B.n545 10.6151
R1373 B.n545 B.n130 10.6151
R1374 B.n541 B.n130 10.6151
R1375 B.n541 B.n540 10.6151
R1376 B.n540 B.n539 10.6151
R1377 B.n539 B.n132 10.6151
R1378 B.n535 B.n132 10.6151
R1379 B.n535 B.n534 10.6151
R1380 B.n534 B.n533 10.6151
R1381 B.n533 B.n134 10.6151
R1382 B.n529 B.n134 10.6151
R1383 B.n529 B.n528 10.6151
R1384 B.n528 B.n527 10.6151
R1385 B.n527 B.n136 10.6151
R1386 B.n523 B.n136 10.6151
R1387 B.n523 B.n522 10.6151
R1388 B.n522 B.n521 10.6151
R1389 B.n521 B.n138 10.6151
R1390 B.n517 B.n138 10.6151
R1391 B.n517 B.n516 10.6151
R1392 B.n516 B.n515 10.6151
R1393 B.n515 B.n140 10.6151
R1394 B.n511 B.n140 10.6151
R1395 B.n511 B.n510 10.6151
R1396 B.n510 B.n509 10.6151
R1397 B.n509 B.n142 10.6151
R1398 B.n505 B.n142 10.6151
R1399 B.n505 B.n504 10.6151
R1400 B.n504 B.n503 10.6151
R1401 B.n503 B.n144 10.6151
R1402 B.n499 B.n144 10.6151
R1403 B.n499 B.n498 10.6151
R1404 B.n498 B.n497 10.6151
R1405 B.n497 B.n146 10.6151
R1406 B.n493 B.n146 10.6151
R1407 B.n493 B.n492 10.6151
R1408 B.n236 B.n1 10.6151
R1409 B.n239 B.n236 10.6151
R1410 B.n240 B.n239 10.6151
R1411 B.n241 B.n240 10.6151
R1412 B.n241 B.n234 10.6151
R1413 B.n245 B.n234 10.6151
R1414 B.n246 B.n245 10.6151
R1415 B.n247 B.n246 10.6151
R1416 B.n247 B.n232 10.6151
R1417 B.n251 B.n232 10.6151
R1418 B.n252 B.n251 10.6151
R1419 B.n253 B.n252 10.6151
R1420 B.n253 B.n230 10.6151
R1421 B.n257 B.n230 10.6151
R1422 B.n258 B.n257 10.6151
R1423 B.n259 B.n258 10.6151
R1424 B.n259 B.n228 10.6151
R1425 B.n263 B.n228 10.6151
R1426 B.n264 B.n263 10.6151
R1427 B.n265 B.n264 10.6151
R1428 B.n265 B.n226 10.6151
R1429 B.n269 B.n226 10.6151
R1430 B.n270 B.n269 10.6151
R1431 B.n271 B.n270 10.6151
R1432 B.n271 B.n224 10.6151
R1433 B.n275 B.n224 10.6151
R1434 B.n276 B.n275 10.6151
R1435 B.n277 B.n276 10.6151
R1436 B.n277 B.n222 10.6151
R1437 B.n281 B.n222 10.6151
R1438 B.n282 B.n281 10.6151
R1439 B.n283 B.n282 10.6151
R1440 B.n283 B.n220 10.6151
R1441 B.n287 B.n220 10.6151
R1442 B.n288 B.n287 10.6151
R1443 B.n289 B.n288 10.6151
R1444 B.n289 B.n218 10.6151
R1445 B.n293 B.n218 10.6151
R1446 B.n294 B.n293 10.6151
R1447 B.n295 B.n294 10.6151
R1448 B.n295 B.n216 10.6151
R1449 B.n299 B.n216 10.6151
R1450 B.n300 B.n299 10.6151
R1451 B.n301 B.n300 10.6151
R1452 B.n301 B.n214 10.6151
R1453 B.n305 B.n214 10.6151
R1454 B.n306 B.n305 10.6151
R1455 B.n307 B.n306 10.6151
R1456 B.n307 B.n212 10.6151
R1457 B.n311 B.n212 10.6151
R1458 B.n312 B.n311 10.6151
R1459 B.n313 B.n312 10.6151
R1460 B.n313 B.n210 10.6151
R1461 B.n317 B.n210 10.6151
R1462 B.n319 B.n318 10.6151
R1463 B.n319 B.n208 10.6151
R1464 B.n323 B.n208 10.6151
R1465 B.n324 B.n323 10.6151
R1466 B.n325 B.n324 10.6151
R1467 B.n325 B.n206 10.6151
R1468 B.n329 B.n206 10.6151
R1469 B.n330 B.n329 10.6151
R1470 B.n331 B.n330 10.6151
R1471 B.n331 B.n204 10.6151
R1472 B.n335 B.n204 10.6151
R1473 B.n336 B.n335 10.6151
R1474 B.n337 B.n336 10.6151
R1475 B.n337 B.n202 10.6151
R1476 B.n341 B.n202 10.6151
R1477 B.n342 B.n341 10.6151
R1478 B.n343 B.n342 10.6151
R1479 B.n343 B.n200 10.6151
R1480 B.n347 B.n200 10.6151
R1481 B.n348 B.n347 10.6151
R1482 B.n349 B.n348 10.6151
R1483 B.n349 B.n198 10.6151
R1484 B.n353 B.n198 10.6151
R1485 B.n354 B.n353 10.6151
R1486 B.n355 B.n354 10.6151
R1487 B.n355 B.n196 10.6151
R1488 B.n359 B.n196 10.6151
R1489 B.n360 B.n359 10.6151
R1490 B.n361 B.n360 10.6151
R1491 B.n361 B.n194 10.6151
R1492 B.n365 B.n194 10.6151
R1493 B.n366 B.n365 10.6151
R1494 B.n367 B.n366 10.6151
R1495 B.n367 B.n192 10.6151
R1496 B.n371 B.n192 10.6151
R1497 B.n372 B.n371 10.6151
R1498 B.n373 B.n372 10.6151
R1499 B.n373 B.n190 10.6151
R1500 B.n377 B.n190 10.6151
R1501 B.n378 B.n377 10.6151
R1502 B.n379 B.n378 10.6151
R1503 B.n379 B.n188 10.6151
R1504 B.n383 B.n188 10.6151
R1505 B.n384 B.n383 10.6151
R1506 B.n385 B.n384 10.6151
R1507 B.n385 B.n186 10.6151
R1508 B.n389 B.n186 10.6151
R1509 B.n390 B.n389 10.6151
R1510 B.n391 B.n390 10.6151
R1511 B.n391 B.n184 10.6151
R1512 B.n395 B.n184 10.6151
R1513 B.n396 B.n395 10.6151
R1514 B.n398 B.n180 10.6151
R1515 B.n402 B.n180 10.6151
R1516 B.n403 B.n402 10.6151
R1517 B.n404 B.n403 10.6151
R1518 B.n404 B.n178 10.6151
R1519 B.n408 B.n178 10.6151
R1520 B.n409 B.n408 10.6151
R1521 B.n410 B.n409 10.6151
R1522 B.n414 B.n413 10.6151
R1523 B.n415 B.n414 10.6151
R1524 B.n415 B.n172 10.6151
R1525 B.n419 B.n172 10.6151
R1526 B.n420 B.n419 10.6151
R1527 B.n421 B.n420 10.6151
R1528 B.n421 B.n170 10.6151
R1529 B.n425 B.n170 10.6151
R1530 B.n426 B.n425 10.6151
R1531 B.n427 B.n426 10.6151
R1532 B.n427 B.n168 10.6151
R1533 B.n431 B.n168 10.6151
R1534 B.n432 B.n431 10.6151
R1535 B.n433 B.n432 10.6151
R1536 B.n433 B.n166 10.6151
R1537 B.n437 B.n166 10.6151
R1538 B.n438 B.n437 10.6151
R1539 B.n439 B.n438 10.6151
R1540 B.n439 B.n164 10.6151
R1541 B.n443 B.n164 10.6151
R1542 B.n444 B.n443 10.6151
R1543 B.n445 B.n444 10.6151
R1544 B.n445 B.n162 10.6151
R1545 B.n449 B.n162 10.6151
R1546 B.n450 B.n449 10.6151
R1547 B.n451 B.n450 10.6151
R1548 B.n451 B.n160 10.6151
R1549 B.n455 B.n160 10.6151
R1550 B.n456 B.n455 10.6151
R1551 B.n457 B.n456 10.6151
R1552 B.n457 B.n158 10.6151
R1553 B.n461 B.n158 10.6151
R1554 B.n462 B.n461 10.6151
R1555 B.n463 B.n462 10.6151
R1556 B.n463 B.n156 10.6151
R1557 B.n467 B.n156 10.6151
R1558 B.n468 B.n467 10.6151
R1559 B.n469 B.n468 10.6151
R1560 B.n469 B.n154 10.6151
R1561 B.n473 B.n154 10.6151
R1562 B.n474 B.n473 10.6151
R1563 B.n475 B.n474 10.6151
R1564 B.n475 B.n152 10.6151
R1565 B.n479 B.n152 10.6151
R1566 B.n480 B.n479 10.6151
R1567 B.n481 B.n480 10.6151
R1568 B.n481 B.n150 10.6151
R1569 B.n485 B.n150 10.6151
R1570 B.n486 B.n485 10.6151
R1571 B.n487 B.n486 10.6151
R1572 B.n487 B.n148 10.6151
R1573 B.n491 B.n148 10.6151
R1574 B.n917 B.n0 8.11757
R1575 B.n917 B.n1 8.11757
R1576 B.n752 B.n58 6.5566
R1577 B.n740 B.n739 6.5566
R1578 B.n398 B.n397 6.5566
R1579 B.n410 B.n176 6.5566
R1580 B.n755 B.n58 4.05904
R1581 B.n739 B.n738 4.05904
R1582 B.n397 B.n396 4.05904
R1583 B.n413 B.n176 4.05904
C0 VN VDD2 9.24823f
C1 VDD1 B 2.68465f
C2 B VTAIL 5.0045f
C3 VDD2 w_n4194_n4126# 2.93258f
C4 VN w_n4194_n4126# 8.29415f
C5 B VDD2 2.78512f
C6 VN B 1.44382f
C7 VDD1 VP 9.644279f
C8 VTAIL VP 9.50584f
C9 B w_n4194_n4126# 12.2579f
C10 VDD1 VTAIL 9.32955f
C11 VDD2 VP 0.551271f
C12 VN VP 8.701099f
C13 VDD1 VDD2 1.83528f
C14 VDD2 VTAIL 9.38805f
C15 VP w_n4194_n4126# 8.83944f
C16 VDD1 VN 0.152066f
C17 VN VTAIL 9.491199f
C18 VDD1 w_n4194_n4126# 2.81234f
C19 B VP 2.35977f
C20 VTAIL w_n4194_n4126# 3.57569f
C21 VDD2 VSUBS 2.28482f
C22 VDD1 VSUBS 2.87058f
C23 VTAIL VSUBS 1.534909f
C24 VN VSUBS 7.03474f
C25 VP VSUBS 3.919866f
C26 B VSUBS 6.04359f
C27 w_n4194_n4126# VSUBS 0.212032p
C28 B.n0 VSUBS 0.006692f
C29 B.n1 VSUBS 0.006692f
C30 B.n2 VSUBS 0.009897f
C31 B.n3 VSUBS 0.007584f
C32 B.n4 VSUBS 0.007584f
C33 B.n5 VSUBS 0.007584f
C34 B.n6 VSUBS 0.007584f
C35 B.n7 VSUBS 0.007584f
C36 B.n8 VSUBS 0.007584f
C37 B.n9 VSUBS 0.007584f
C38 B.n10 VSUBS 0.007584f
C39 B.n11 VSUBS 0.007584f
C40 B.n12 VSUBS 0.007584f
C41 B.n13 VSUBS 0.007584f
C42 B.n14 VSUBS 0.007584f
C43 B.n15 VSUBS 0.007584f
C44 B.n16 VSUBS 0.007584f
C45 B.n17 VSUBS 0.007584f
C46 B.n18 VSUBS 0.007584f
C47 B.n19 VSUBS 0.007584f
C48 B.n20 VSUBS 0.007584f
C49 B.n21 VSUBS 0.007584f
C50 B.n22 VSUBS 0.007584f
C51 B.n23 VSUBS 0.007584f
C52 B.n24 VSUBS 0.007584f
C53 B.n25 VSUBS 0.007584f
C54 B.n26 VSUBS 0.007584f
C55 B.n27 VSUBS 0.007584f
C56 B.n28 VSUBS 0.007584f
C57 B.n29 VSUBS 0.01756f
C58 B.n30 VSUBS 0.007584f
C59 B.n31 VSUBS 0.007584f
C60 B.n32 VSUBS 0.007584f
C61 B.n33 VSUBS 0.007584f
C62 B.n34 VSUBS 0.007584f
C63 B.n35 VSUBS 0.007584f
C64 B.n36 VSUBS 0.007584f
C65 B.n37 VSUBS 0.007584f
C66 B.n38 VSUBS 0.007584f
C67 B.n39 VSUBS 0.007584f
C68 B.n40 VSUBS 0.007584f
C69 B.n41 VSUBS 0.007584f
C70 B.n42 VSUBS 0.007584f
C71 B.n43 VSUBS 0.007584f
C72 B.n44 VSUBS 0.007584f
C73 B.n45 VSUBS 0.007584f
C74 B.n46 VSUBS 0.007584f
C75 B.n47 VSUBS 0.007584f
C76 B.n48 VSUBS 0.007584f
C77 B.n49 VSUBS 0.007584f
C78 B.n50 VSUBS 0.007584f
C79 B.n51 VSUBS 0.007584f
C80 B.n52 VSUBS 0.007584f
C81 B.n53 VSUBS 0.007584f
C82 B.n54 VSUBS 0.007584f
C83 B.n55 VSUBS 0.007584f
C84 B.t1 VSUBS 0.571933f
C85 B.t2 VSUBS 0.602007f
C86 B.t0 VSUBS 2.9024f
C87 B.n56 VSUBS 0.36039f
C88 B.n57 VSUBS 0.082964f
C89 B.n58 VSUBS 0.017572f
C90 B.n59 VSUBS 0.007584f
C91 B.n60 VSUBS 0.007584f
C92 B.n61 VSUBS 0.007584f
C93 B.n62 VSUBS 0.007584f
C94 B.n63 VSUBS 0.007584f
C95 B.t7 VSUBS 0.571916f
C96 B.t8 VSUBS 0.601994f
C97 B.t6 VSUBS 2.9024f
C98 B.n64 VSUBS 0.360403f
C99 B.n65 VSUBS 0.082982f
C100 B.n66 VSUBS 0.007584f
C101 B.n67 VSUBS 0.007584f
C102 B.n68 VSUBS 0.007584f
C103 B.n69 VSUBS 0.007584f
C104 B.n70 VSUBS 0.007584f
C105 B.n71 VSUBS 0.007584f
C106 B.n72 VSUBS 0.007584f
C107 B.n73 VSUBS 0.007584f
C108 B.n74 VSUBS 0.007584f
C109 B.n75 VSUBS 0.007584f
C110 B.n76 VSUBS 0.007584f
C111 B.n77 VSUBS 0.007584f
C112 B.n78 VSUBS 0.007584f
C113 B.n79 VSUBS 0.007584f
C114 B.n80 VSUBS 0.007584f
C115 B.n81 VSUBS 0.007584f
C116 B.n82 VSUBS 0.007584f
C117 B.n83 VSUBS 0.007584f
C118 B.n84 VSUBS 0.007584f
C119 B.n85 VSUBS 0.007584f
C120 B.n86 VSUBS 0.007584f
C121 B.n87 VSUBS 0.007584f
C122 B.n88 VSUBS 0.007584f
C123 B.n89 VSUBS 0.007584f
C124 B.n90 VSUBS 0.007584f
C125 B.n91 VSUBS 0.018354f
C126 B.n92 VSUBS 0.007584f
C127 B.n93 VSUBS 0.007584f
C128 B.n94 VSUBS 0.007584f
C129 B.n95 VSUBS 0.007584f
C130 B.n96 VSUBS 0.007584f
C131 B.n97 VSUBS 0.007584f
C132 B.n98 VSUBS 0.007584f
C133 B.n99 VSUBS 0.007584f
C134 B.n100 VSUBS 0.007584f
C135 B.n101 VSUBS 0.007584f
C136 B.n102 VSUBS 0.007584f
C137 B.n103 VSUBS 0.007584f
C138 B.n104 VSUBS 0.007584f
C139 B.n105 VSUBS 0.007584f
C140 B.n106 VSUBS 0.007584f
C141 B.n107 VSUBS 0.007584f
C142 B.n108 VSUBS 0.007584f
C143 B.n109 VSUBS 0.007584f
C144 B.n110 VSUBS 0.007584f
C145 B.n111 VSUBS 0.007584f
C146 B.n112 VSUBS 0.007584f
C147 B.n113 VSUBS 0.007584f
C148 B.n114 VSUBS 0.007584f
C149 B.n115 VSUBS 0.007584f
C150 B.n116 VSUBS 0.007584f
C151 B.n117 VSUBS 0.007584f
C152 B.n118 VSUBS 0.007584f
C153 B.n119 VSUBS 0.007584f
C154 B.n120 VSUBS 0.007584f
C155 B.n121 VSUBS 0.007584f
C156 B.n122 VSUBS 0.007584f
C157 B.n123 VSUBS 0.007584f
C158 B.n124 VSUBS 0.007584f
C159 B.n125 VSUBS 0.007584f
C160 B.n126 VSUBS 0.007584f
C161 B.n127 VSUBS 0.007584f
C162 B.n128 VSUBS 0.007584f
C163 B.n129 VSUBS 0.007584f
C164 B.n130 VSUBS 0.007584f
C165 B.n131 VSUBS 0.007584f
C166 B.n132 VSUBS 0.007584f
C167 B.n133 VSUBS 0.007584f
C168 B.n134 VSUBS 0.007584f
C169 B.n135 VSUBS 0.007584f
C170 B.n136 VSUBS 0.007584f
C171 B.n137 VSUBS 0.007584f
C172 B.n138 VSUBS 0.007584f
C173 B.n139 VSUBS 0.007584f
C174 B.n140 VSUBS 0.007584f
C175 B.n141 VSUBS 0.007584f
C176 B.n142 VSUBS 0.007584f
C177 B.n143 VSUBS 0.007584f
C178 B.n144 VSUBS 0.007584f
C179 B.n145 VSUBS 0.007584f
C180 B.n146 VSUBS 0.007584f
C181 B.n147 VSUBS 0.01756f
C182 B.n148 VSUBS 0.007584f
C183 B.n149 VSUBS 0.007584f
C184 B.n150 VSUBS 0.007584f
C185 B.n151 VSUBS 0.007584f
C186 B.n152 VSUBS 0.007584f
C187 B.n153 VSUBS 0.007584f
C188 B.n154 VSUBS 0.007584f
C189 B.n155 VSUBS 0.007584f
C190 B.n156 VSUBS 0.007584f
C191 B.n157 VSUBS 0.007584f
C192 B.n158 VSUBS 0.007584f
C193 B.n159 VSUBS 0.007584f
C194 B.n160 VSUBS 0.007584f
C195 B.n161 VSUBS 0.007584f
C196 B.n162 VSUBS 0.007584f
C197 B.n163 VSUBS 0.007584f
C198 B.n164 VSUBS 0.007584f
C199 B.n165 VSUBS 0.007584f
C200 B.n166 VSUBS 0.007584f
C201 B.n167 VSUBS 0.007584f
C202 B.n168 VSUBS 0.007584f
C203 B.n169 VSUBS 0.007584f
C204 B.n170 VSUBS 0.007584f
C205 B.n171 VSUBS 0.007584f
C206 B.n172 VSUBS 0.007584f
C207 B.n173 VSUBS 0.007584f
C208 B.t5 VSUBS 0.571916f
C209 B.t4 VSUBS 0.601994f
C210 B.t3 VSUBS 2.9024f
C211 B.n174 VSUBS 0.360403f
C212 B.n175 VSUBS 0.082982f
C213 B.n176 VSUBS 0.017572f
C214 B.n177 VSUBS 0.007584f
C215 B.n178 VSUBS 0.007584f
C216 B.n179 VSUBS 0.007584f
C217 B.n180 VSUBS 0.007584f
C218 B.n181 VSUBS 0.007584f
C219 B.t11 VSUBS 0.571933f
C220 B.t10 VSUBS 0.602007f
C221 B.t9 VSUBS 2.9024f
C222 B.n182 VSUBS 0.36039f
C223 B.n183 VSUBS 0.082964f
C224 B.n184 VSUBS 0.007584f
C225 B.n185 VSUBS 0.007584f
C226 B.n186 VSUBS 0.007584f
C227 B.n187 VSUBS 0.007584f
C228 B.n188 VSUBS 0.007584f
C229 B.n189 VSUBS 0.007584f
C230 B.n190 VSUBS 0.007584f
C231 B.n191 VSUBS 0.007584f
C232 B.n192 VSUBS 0.007584f
C233 B.n193 VSUBS 0.007584f
C234 B.n194 VSUBS 0.007584f
C235 B.n195 VSUBS 0.007584f
C236 B.n196 VSUBS 0.007584f
C237 B.n197 VSUBS 0.007584f
C238 B.n198 VSUBS 0.007584f
C239 B.n199 VSUBS 0.007584f
C240 B.n200 VSUBS 0.007584f
C241 B.n201 VSUBS 0.007584f
C242 B.n202 VSUBS 0.007584f
C243 B.n203 VSUBS 0.007584f
C244 B.n204 VSUBS 0.007584f
C245 B.n205 VSUBS 0.007584f
C246 B.n206 VSUBS 0.007584f
C247 B.n207 VSUBS 0.007584f
C248 B.n208 VSUBS 0.007584f
C249 B.n209 VSUBS 0.018354f
C250 B.n210 VSUBS 0.007584f
C251 B.n211 VSUBS 0.007584f
C252 B.n212 VSUBS 0.007584f
C253 B.n213 VSUBS 0.007584f
C254 B.n214 VSUBS 0.007584f
C255 B.n215 VSUBS 0.007584f
C256 B.n216 VSUBS 0.007584f
C257 B.n217 VSUBS 0.007584f
C258 B.n218 VSUBS 0.007584f
C259 B.n219 VSUBS 0.007584f
C260 B.n220 VSUBS 0.007584f
C261 B.n221 VSUBS 0.007584f
C262 B.n222 VSUBS 0.007584f
C263 B.n223 VSUBS 0.007584f
C264 B.n224 VSUBS 0.007584f
C265 B.n225 VSUBS 0.007584f
C266 B.n226 VSUBS 0.007584f
C267 B.n227 VSUBS 0.007584f
C268 B.n228 VSUBS 0.007584f
C269 B.n229 VSUBS 0.007584f
C270 B.n230 VSUBS 0.007584f
C271 B.n231 VSUBS 0.007584f
C272 B.n232 VSUBS 0.007584f
C273 B.n233 VSUBS 0.007584f
C274 B.n234 VSUBS 0.007584f
C275 B.n235 VSUBS 0.007584f
C276 B.n236 VSUBS 0.007584f
C277 B.n237 VSUBS 0.007584f
C278 B.n238 VSUBS 0.007584f
C279 B.n239 VSUBS 0.007584f
C280 B.n240 VSUBS 0.007584f
C281 B.n241 VSUBS 0.007584f
C282 B.n242 VSUBS 0.007584f
C283 B.n243 VSUBS 0.007584f
C284 B.n244 VSUBS 0.007584f
C285 B.n245 VSUBS 0.007584f
C286 B.n246 VSUBS 0.007584f
C287 B.n247 VSUBS 0.007584f
C288 B.n248 VSUBS 0.007584f
C289 B.n249 VSUBS 0.007584f
C290 B.n250 VSUBS 0.007584f
C291 B.n251 VSUBS 0.007584f
C292 B.n252 VSUBS 0.007584f
C293 B.n253 VSUBS 0.007584f
C294 B.n254 VSUBS 0.007584f
C295 B.n255 VSUBS 0.007584f
C296 B.n256 VSUBS 0.007584f
C297 B.n257 VSUBS 0.007584f
C298 B.n258 VSUBS 0.007584f
C299 B.n259 VSUBS 0.007584f
C300 B.n260 VSUBS 0.007584f
C301 B.n261 VSUBS 0.007584f
C302 B.n262 VSUBS 0.007584f
C303 B.n263 VSUBS 0.007584f
C304 B.n264 VSUBS 0.007584f
C305 B.n265 VSUBS 0.007584f
C306 B.n266 VSUBS 0.007584f
C307 B.n267 VSUBS 0.007584f
C308 B.n268 VSUBS 0.007584f
C309 B.n269 VSUBS 0.007584f
C310 B.n270 VSUBS 0.007584f
C311 B.n271 VSUBS 0.007584f
C312 B.n272 VSUBS 0.007584f
C313 B.n273 VSUBS 0.007584f
C314 B.n274 VSUBS 0.007584f
C315 B.n275 VSUBS 0.007584f
C316 B.n276 VSUBS 0.007584f
C317 B.n277 VSUBS 0.007584f
C318 B.n278 VSUBS 0.007584f
C319 B.n279 VSUBS 0.007584f
C320 B.n280 VSUBS 0.007584f
C321 B.n281 VSUBS 0.007584f
C322 B.n282 VSUBS 0.007584f
C323 B.n283 VSUBS 0.007584f
C324 B.n284 VSUBS 0.007584f
C325 B.n285 VSUBS 0.007584f
C326 B.n286 VSUBS 0.007584f
C327 B.n287 VSUBS 0.007584f
C328 B.n288 VSUBS 0.007584f
C329 B.n289 VSUBS 0.007584f
C330 B.n290 VSUBS 0.007584f
C331 B.n291 VSUBS 0.007584f
C332 B.n292 VSUBS 0.007584f
C333 B.n293 VSUBS 0.007584f
C334 B.n294 VSUBS 0.007584f
C335 B.n295 VSUBS 0.007584f
C336 B.n296 VSUBS 0.007584f
C337 B.n297 VSUBS 0.007584f
C338 B.n298 VSUBS 0.007584f
C339 B.n299 VSUBS 0.007584f
C340 B.n300 VSUBS 0.007584f
C341 B.n301 VSUBS 0.007584f
C342 B.n302 VSUBS 0.007584f
C343 B.n303 VSUBS 0.007584f
C344 B.n304 VSUBS 0.007584f
C345 B.n305 VSUBS 0.007584f
C346 B.n306 VSUBS 0.007584f
C347 B.n307 VSUBS 0.007584f
C348 B.n308 VSUBS 0.007584f
C349 B.n309 VSUBS 0.007584f
C350 B.n310 VSUBS 0.007584f
C351 B.n311 VSUBS 0.007584f
C352 B.n312 VSUBS 0.007584f
C353 B.n313 VSUBS 0.007584f
C354 B.n314 VSUBS 0.007584f
C355 B.n315 VSUBS 0.007584f
C356 B.n316 VSUBS 0.01756f
C357 B.n317 VSUBS 0.01756f
C358 B.n318 VSUBS 0.018354f
C359 B.n319 VSUBS 0.007584f
C360 B.n320 VSUBS 0.007584f
C361 B.n321 VSUBS 0.007584f
C362 B.n322 VSUBS 0.007584f
C363 B.n323 VSUBS 0.007584f
C364 B.n324 VSUBS 0.007584f
C365 B.n325 VSUBS 0.007584f
C366 B.n326 VSUBS 0.007584f
C367 B.n327 VSUBS 0.007584f
C368 B.n328 VSUBS 0.007584f
C369 B.n329 VSUBS 0.007584f
C370 B.n330 VSUBS 0.007584f
C371 B.n331 VSUBS 0.007584f
C372 B.n332 VSUBS 0.007584f
C373 B.n333 VSUBS 0.007584f
C374 B.n334 VSUBS 0.007584f
C375 B.n335 VSUBS 0.007584f
C376 B.n336 VSUBS 0.007584f
C377 B.n337 VSUBS 0.007584f
C378 B.n338 VSUBS 0.007584f
C379 B.n339 VSUBS 0.007584f
C380 B.n340 VSUBS 0.007584f
C381 B.n341 VSUBS 0.007584f
C382 B.n342 VSUBS 0.007584f
C383 B.n343 VSUBS 0.007584f
C384 B.n344 VSUBS 0.007584f
C385 B.n345 VSUBS 0.007584f
C386 B.n346 VSUBS 0.007584f
C387 B.n347 VSUBS 0.007584f
C388 B.n348 VSUBS 0.007584f
C389 B.n349 VSUBS 0.007584f
C390 B.n350 VSUBS 0.007584f
C391 B.n351 VSUBS 0.007584f
C392 B.n352 VSUBS 0.007584f
C393 B.n353 VSUBS 0.007584f
C394 B.n354 VSUBS 0.007584f
C395 B.n355 VSUBS 0.007584f
C396 B.n356 VSUBS 0.007584f
C397 B.n357 VSUBS 0.007584f
C398 B.n358 VSUBS 0.007584f
C399 B.n359 VSUBS 0.007584f
C400 B.n360 VSUBS 0.007584f
C401 B.n361 VSUBS 0.007584f
C402 B.n362 VSUBS 0.007584f
C403 B.n363 VSUBS 0.007584f
C404 B.n364 VSUBS 0.007584f
C405 B.n365 VSUBS 0.007584f
C406 B.n366 VSUBS 0.007584f
C407 B.n367 VSUBS 0.007584f
C408 B.n368 VSUBS 0.007584f
C409 B.n369 VSUBS 0.007584f
C410 B.n370 VSUBS 0.007584f
C411 B.n371 VSUBS 0.007584f
C412 B.n372 VSUBS 0.007584f
C413 B.n373 VSUBS 0.007584f
C414 B.n374 VSUBS 0.007584f
C415 B.n375 VSUBS 0.007584f
C416 B.n376 VSUBS 0.007584f
C417 B.n377 VSUBS 0.007584f
C418 B.n378 VSUBS 0.007584f
C419 B.n379 VSUBS 0.007584f
C420 B.n380 VSUBS 0.007584f
C421 B.n381 VSUBS 0.007584f
C422 B.n382 VSUBS 0.007584f
C423 B.n383 VSUBS 0.007584f
C424 B.n384 VSUBS 0.007584f
C425 B.n385 VSUBS 0.007584f
C426 B.n386 VSUBS 0.007584f
C427 B.n387 VSUBS 0.007584f
C428 B.n388 VSUBS 0.007584f
C429 B.n389 VSUBS 0.007584f
C430 B.n390 VSUBS 0.007584f
C431 B.n391 VSUBS 0.007584f
C432 B.n392 VSUBS 0.007584f
C433 B.n393 VSUBS 0.007584f
C434 B.n394 VSUBS 0.007584f
C435 B.n395 VSUBS 0.007584f
C436 B.n396 VSUBS 0.005242f
C437 B.n397 VSUBS 0.017572f
C438 B.n398 VSUBS 0.006134f
C439 B.n399 VSUBS 0.007584f
C440 B.n400 VSUBS 0.007584f
C441 B.n401 VSUBS 0.007584f
C442 B.n402 VSUBS 0.007584f
C443 B.n403 VSUBS 0.007584f
C444 B.n404 VSUBS 0.007584f
C445 B.n405 VSUBS 0.007584f
C446 B.n406 VSUBS 0.007584f
C447 B.n407 VSUBS 0.007584f
C448 B.n408 VSUBS 0.007584f
C449 B.n409 VSUBS 0.007584f
C450 B.n410 VSUBS 0.006134f
C451 B.n411 VSUBS 0.007584f
C452 B.n412 VSUBS 0.007584f
C453 B.n413 VSUBS 0.005242f
C454 B.n414 VSUBS 0.007584f
C455 B.n415 VSUBS 0.007584f
C456 B.n416 VSUBS 0.007584f
C457 B.n417 VSUBS 0.007584f
C458 B.n418 VSUBS 0.007584f
C459 B.n419 VSUBS 0.007584f
C460 B.n420 VSUBS 0.007584f
C461 B.n421 VSUBS 0.007584f
C462 B.n422 VSUBS 0.007584f
C463 B.n423 VSUBS 0.007584f
C464 B.n424 VSUBS 0.007584f
C465 B.n425 VSUBS 0.007584f
C466 B.n426 VSUBS 0.007584f
C467 B.n427 VSUBS 0.007584f
C468 B.n428 VSUBS 0.007584f
C469 B.n429 VSUBS 0.007584f
C470 B.n430 VSUBS 0.007584f
C471 B.n431 VSUBS 0.007584f
C472 B.n432 VSUBS 0.007584f
C473 B.n433 VSUBS 0.007584f
C474 B.n434 VSUBS 0.007584f
C475 B.n435 VSUBS 0.007584f
C476 B.n436 VSUBS 0.007584f
C477 B.n437 VSUBS 0.007584f
C478 B.n438 VSUBS 0.007584f
C479 B.n439 VSUBS 0.007584f
C480 B.n440 VSUBS 0.007584f
C481 B.n441 VSUBS 0.007584f
C482 B.n442 VSUBS 0.007584f
C483 B.n443 VSUBS 0.007584f
C484 B.n444 VSUBS 0.007584f
C485 B.n445 VSUBS 0.007584f
C486 B.n446 VSUBS 0.007584f
C487 B.n447 VSUBS 0.007584f
C488 B.n448 VSUBS 0.007584f
C489 B.n449 VSUBS 0.007584f
C490 B.n450 VSUBS 0.007584f
C491 B.n451 VSUBS 0.007584f
C492 B.n452 VSUBS 0.007584f
C493 B.n453 VSUBS 0.007584f
C494 B.n454 VSUBS 0.007584f
C495 B.n455 VSUBS 0.007584f
C496 B.n456 VSUBS 0.007584f
C497 B.n457 VSUBS 0.007584f
C498 B.n458 VSUBS 0.007584f
C499 B.n459 VSUBS 0.007584f
C500 B.n460 VSUBS 0.007584f
C501 B.n461 VSUBS 0.007584f
C502 B.n462 VSUBS 0.007584f
C503 B.n463 VSUBS 0.007584f
C504 B.n464 VSUBS 0.007584f
C505 B.n465 VSUBS 0.007584f
C506 B.n466 VSUBS 0.007584f
C507 B.n467 VSUBS 0.007584f
C508 B.n468 VSUBS 0.007584f
C509 B.n469 VSUBS 0.007584f
C510 B.n470 VSUBS 0.007584f
C511 B.n471 VSUBS 0.007584f
C512 B.n472 VSUBS 0.007584f
C513 B.n473 VSUBS 0.007584f
C514 B.n474 VSUBS 0.007584f
C515 B.n475 VSUBS 0.007584f
C516 B.n476 VSUBS 0.007584f
C517 B.n477 VSUBS 0.007584f
C518 B.n478 VSUBS 0.007584f
C519 B.n479 VSUBS 0.007584f
C520 B.n480 VSUBS 0.007584f
C521 B.n481 VSUBS 0.007584f
C522 B.n482 VSUBS 0.007584f
C523 B.n483 VSUBS 0.007584f
C524 B.n484 VSUBS 0.007584f
C525 B.n485 VSUBS 0.007584f
C526 B.n486 VSUBS 0.007584f
C527 B.n487 VSUBS 0.007584f
C528 B.n488 VSUBS 0.007584f
C529 B.n489 VSUBS 0.007584f
C530 B.n490 VSUBS 0.018354f
C531 B.n491 VSUBS 0.017474f
C532 B.n492 VSUBS 0.01844f
C533 B.n493 VSUBS 0.007584f
C534 B.n494 VSUBS 0.007584f
C535 B.n495 VSUBS 0.007584f
C536 B.n496 VSUBS 0.007584f
C537 B.n497 VSUBS 0.007584f
C538 B.n498 VSUBS 0.007584f
C539 B.n499 VSUBS 0.007584f
C540 B.n500 VSUBS 0.007584f
C541 B.n501 VSUBS 0.007584f
C542 B.n502 VSUBS 0.007584f
C543 B.n503 VSUBS 0.007584f
C544 B.n504 VSUBS 0.007584f
C545 B.n505 VSUBS 0.007584f
C546 B.n506 VSUBS 0.007584f
C547 B.n507 VSUBS 0.007584f
C548 B.n508 VSUBS 0.007584f
C549 B.n509 VSUBS 0.007584f
C550 B.n510 VSUBS 0.007584f
C551 B.n511 VSUBS 0.007584f
C552 B.n512 VSUBS 0.007584f
C553 B.n513 VSUBS 0.007584f
C554 B.n514 VSUBS 0.007584f
C555 B.n515 VSUBS 0.007584f
C556 B.n516 VSUBS 0.007584f
C557 B.n517 VSUBS 0.007584f
C558 B.n518 VSUBS 0.007584f
C559 B.n519 VSUBS 0.007584f
C560 B.n520 VSUBS 0.007584f
C561 B.n521 VSUBS 0.007584f
C562 B.n522 VSUBS 0.007584f
C563 B.n523 VSUBS 0.007584f
C564 B.n524 VSUBS 0.007584f
C565 B.n525 VSUBS 0.007584f
C566 B.n526 VSUBS 0.007584f
C567 B.n527 VSUBS 0.007584f
C568 B.n528 VSUBS 0.007584f
C569 B.n529 VSUBS 0.007584f
C570 B.n530 VSUBS 0.007584f
C571 B.n531 VSUBS 0.007584f
C572 B.n532 VSUBS 0.007584f
C573 B.n533 VSUBS 0.007584f
C574 B.n534 VSUBS 0.007584f
C575 B.n535 VSUBS 0.007584f
C576 B.n536 VSUBS 0.007584f
C577 B.n537 VSUBS 0.007584f
C578 B.n538 VSUBS 0.007584f
C579 B.n539 VSUBS 0.007584f
C580 B.n540 VSUBS 0.007584f
C581 B.n541 VSUBS 0.007584f
C582 B.n542 VSUBS 0.007584f
C583 B.n543 VSUBS 0.007584f
C584 B.n544 VSUBS 0.007584f
C585 B.n545 VSUBS 0.007584f
C586 B.n546 VSUBS 0.007584f
C587 B.n547 VSUBS 0.007584f
C588 B.n548 VSUBS 0.007584f
C589 B.n549 VSUBS 0.007584f
C590 B.n550 VSUBS 0.007584f
C591 B.n551 VSUBS 0.007584f
C592 B.n552 VSUBS 0.007584f
C593 B.n553 VSUBS 0.007584f
C594 B.n554 VSUBS 0.007584f
C595 B.n555 VSUBS 0.007584f
C596 B.n556 VSUBS 0.007584f
C597 B.n557 VSUBS 0.007584f
C598 B.n558 VSUBS 0.007584f
C599 B.n559 VSUBS 0.007584f
C600 B.n560 VSUBS 0.007584f
C601 B.n561 VSUBS 0.007584f
C602 B.n562 VSUBS 0.007584f
C603 B.n563 VSUBS 0.007584f
C604 B.n564 VSUBS 0.007584f
C605 B.n565 VSUBS 0.007584f
C606 B.n566 VSUBS 0.007584f
C607 B.n567 VSUBS 0.007584f
C608 B.n568 VSUBS 0.007584f
C609 B.n569 VSUBS 0.007584f
C610 B.n570 VSUBS 0.007584f
C611 B.n571 VSUBS 0.007584f
C612 B.n572 VSUBS 0.007584f
C613 B.n573 VSUBS 0.007584f
C614 B.n574 VSUBS 0.007584f
C615 B.n575 VSUBS 0.007584f
C616 B.n576 VSUBS 0.007584f
C617 B.n577 VSUBS 0.007584f
C618 B.n578 VSUBS 0.007584f
C619 B.n579 VSUBS 0.007584f
C620 B.n580 VSUBS 0.007584f
C621 B.n581 VSUBS 0.007584f
C622 B.n582 VSUBS 0.007584f
C623 B.n583 VSUBS 0.007584f
C624 B.n584 VSUBS 0.007584f
C625 B.n585 VSUBS 0.007584f
C626 B.n586 VSUBS 0.007584f
C627 B.n587 VSUBS 0.007584f
C628 B.n588 VSUBS 0.007584f
C629 B.n589 VSUBS 0.007584f
C630 B.n590 VSUBS 0.007584f
C631 B.n591 VSUBS 0.007584f
C632 B.n592 VSUBS 0.007584f
C633 B.n593 VSUBS 0.007584f
C634 B.n594 VSUBS 0.007584f
C635 B.n595 VSUBS 0.007584f
C636 B.n596 VSUBS 0.007584f
C637 B.n597 VSUBS 0.007584f
C638 B.n598 VSUBS 0.007584f
C639 B.n599 VSUBS 0.007584f
C640 B.n600 VSUBS 0.007584f
C641 B.n601 VSUBS 0.007584f
C642 B.n602 VSUBS 0.007584f
C643 B.n603 VSUBS 0.007584f
C644 B.n604 VSUBS 0.007584f
C645 B.n605 VSUBS 0.007584f
C646 B.n606 VSUBS 0.007584f
C647 B.n607 VSUBS 0.007584f
C648 B.n608 VSUBS 0.007584f
C649 B.n609 VSUBS 0.007584f
C650 B.n610 VSUBS 0.007584f
C651 B.n611 VSUBS 0.007584f
C652 B.n612 VSUBS 0.007584f
C653 B.n613 VSUBS 0.007584f
C654 B.n614 VSUBS 0.007584f
C655 B.n615 VSUBS 0.007584f
C656 B.n616 VSUBS 0.007584f
C657 B.n617 VSUBS 0.007584f
C658 B.n618 VSUBS 0.007584f
C659 B.n619 VSUBS 0.007584f
C660 B.n620 VSUBS 0.007584f
C661 B.n621 VSUBS 0.007584f
C662 B.n622 VSUBS 0.007584f
C663 B.n623 VSUBS 0.007584f
C664 B.n624 VSUBS 0.007584f
C665 B.n625 VSUBS 0.007584f
C666 B.n626 VSUBS 0.007584f
C667 B.n627 VSUBS 0.007584f
C668 B.n628 VSUBS 0.007584f
C669 B.n629 VSUBS 0.007584f
C670 B.n630 VSUBS 0.007584f
C671 B.n631 VSUBS 0.007584f
C672 B.n632 VSUBS 0.007584f
C673 B.n633 VSUBS 0.007584f
C674 B.n634 VSUBS 0.007584f
C675 B.n635 VSUBS 0.007584f
C676 B.n636 VSUBS 0.007584f
C677 B.n637 VSUBS 0.007584f
C678 B.n638 VSUBS 0.007584f
C679 B.n639 VSUBS 0.007584f
C680 B.n640 VSUBS 0.007584f
C681 B.n641 VSUBS 0.007584f
C682 B.n642 VSUBS 0.007584f
C683 B.n643 VSUBS 0.007584f
C684 B.n644 VSUBS 0.007584f
C685 B.n645 VSUBS 0.007584f
C686 B.n646 VSUBS 0.007584f
C687 B.n647 VSUBS 0.007584f
C688 B.n648 VSUBS 0.007584f
C689 B.n649 VSUBS 0.007584f
C690 B.n650 VSUBS 0.007584f
C691 B.n651 VSUBS 0.007584f
C692 B.n652 VSUBS 0.007584f
C693 B.n653 VSUBS 0.007584f
C694 B.n654 VSUBS 0.007584f
C695 B.n655 VSUBS 0.007584f
C696 B.n656 VSUBS 0.007584f
C697 B.n657 VSUBS 0.007584f
C698 B.n658 VSUBS 0.01756f
C699 B.n659 VSUBS 0.01756f
C700 B.n660 VSUBS 0.018354f
C701 B.n661 VSUBS 0.007584f
C702 B.n662 VSUBS 0.007584f
C703 B.n663 VSUBS 0.007584f
C704 B.n664 VSUBS 0.007584f
C705 B.n665 VSUBS 0.007584f
C706 B.n666 VSUBS 0.007584f
C707 B.n667 VSUBS 0.007584f
C708 B.n668 VSUBS 0.007584f
C709 B.n669 VSUBS 0.007584f
C710 B.n670 VSUBS 0.007584f
C711 B.n671 VSUBS 0.007584f
C712 B.n672 VSUBS 0.007584f
C713 B.n673 VSUBS 0.007584f
C714 B.n674 VSUBS 0.007584f
C715 B.n675 VSUBS 0.007584f
C716 B.n676 VSUBS 0.007584f
C717 B.n677 VSUBS 0.007584f
C718 B.n678 VSUBS 0.007584f
C719 B.n679 VSUBS 0.007584f
C720 B.n680 VSUBS 0.007584f
C721 B.n681 VSUBS 0.007584f
C722 B.n682 VSUBS 0.007584f
C723 B.n683 VSUBS 0.007584f
C724 B.n684 VSUBS 0.007584f
C725 B.n685 VSUBS 0.007584f
C726 B.n686 VSUBS 0.007584f
C727 B.n687 VSUBS 0.007584f
C728 B.n688 VSUBS 0.007584f
C729 B.n689 VSUBS 0.007584f
C730 B.n690 VSUBS 0.007584f
C731 B.n691 VSUBS 0.007584f
C732 B.n692 VSUBS 0.007584f
C733 B.n693 VSUBS 0.007584f
C734 B.n694 VSUBS 0.007584f
C735 B.n695 VSUBS 0.007584f
C736 B.n696 VSUBS 0.007584f
C737 B.n697 VSUBS 0.007584f
C738 B.n698 VSUBS 0.007584f
C739 B.n699 VSUBS 0.007584f
C740 B.n700 VSUBS 0.007584f
C741 B.n701 VSUBS 0.007584f
C742 B.n702 VSUBS 0.007584f
C743 B.n703 VSUBS 0.007584f
C744 B.n704 VSUBS 0.007584f
C745 B.n705 VSUBS 0.007584f
C746 B.n706 VSUBS 0.007584f
C747 B.n707 VSUBS 0.007584f
C748 B.n708 VSUBS 0.007584f
C749 B.n709 VSUBS 0.007584f
C750 B.n710 VSUBS 0.007584f
C751 B.n711 VSUBS 0.007584f
C752 B.n712 VSUBS 0.007584f
C753 B.n713 VSUBS 0.007584f
C754 B.n714 VSUBS 0.007584f
C755 B.n715 VSUBS 0.007584f
C756 B.n716 VSUBS 0.007584f
C757 B.n717 VSUBS 0.007584f
C758 B.n718 VSUBS 0.007584f
C759 B.n719 VSUBS 0.007584f
C760 B.n720 VSUBS 0.007584f
C761 B.n721 VSUBS 0.007584f
C762 B.n722 VSUBS 0.007584f
C763 B.n723 VSUBS 0.007584f
C764 B.n724 VSUBS 0.007584f
C765 B.n725 VSUBS 0.007584f
C766 B.n726 VSUBS 0.007584f
C767 B.n727 VSUBS 0.007584f
C768 B.n728 VSUBS 0.007584f
C769 B.n729 VSUBS 0.007584f
C770 B.n730 VSUBS 0.007584f
C771 B.n731 VSUBS 0.007584f
C772 B.n732 VSUBS 0.007584f
C773 B.n733 VSUBS 0.007584f
C774 B.n734 VSUBS 0.007584f
C775 B.n735 VSUBS 0.007584f
C776 B.n736 VSUBS 0.007584f
C777 B.n737 VSUBS 0.007584f
C778 B.n738 VSUBS 0.005242f
C779 B.n739 VSUBS 0.017572f
C780 B.n740 VSUBS 0.006134f
C781 B.n741 VSUBS 0.007584f
C782 B.n742 VSUBS 0.007584f
C783 B.n743 VSUBS 0.007584f
C784 B.n744 VSUBS 0.007584f
C785 B.n745 VSUBS 0.007584f
C786 B.n746 VSUBS 0.007584f
C787 B.n747 VSUBS 0.007584f
C788 B.n748 VSUBS 0.007584f
C789 B.n749 VSUBS 0.007584f
C790 B.n750 VSUBS 0.007584f
C791 B.n751 VSUBS 0.007584f
C792 B.n752 VSUBS 0.006134f
C793 B.n753 VSUBS 0.007584f
C794 B.n754 VSUBS 0.007584f
C795 B.n755 VSUBS 0.005242f
C796 B.n756 VSUBS 0.007584f
C797 B.n757 VSUBS 0.007584f
C798 B.n758 VSUBS 0.007584f
C799 B.n759 VSUBS 0.007584f
C800 B.n760 VSUBS 0.007584f
C801 B.n761 VSUBS 0.007584f
C802 B.n762 VSUBS 0.007584f
C803 B.n763 VSUBS 0.007584f
C804 B.n764 VSUBS 0.007584f
C805 B.n765 VSUBS 0.007584f
C806 B.n766 VSUBS 0.007584f
C807 B.n767 VSUBS 0.007584f
C808 B.n768 VSUBS 0.007584f
C809 B.n769 VSUBS 0.007584f
C810 B.n770 VSUBS 0.007584f
C811 B.n771 VSUBS 0.007584f
C812 B.n772 VSUBS 0.007584f
C813 B.n773 VSUBS 0.007584f
C814 B.n774 VSUBS 0.007584f
C815 B.n775 VSUBS 0.007584f
C816 B.n776 VSUBS 0.007584f
C817 B.n777 VSUBS 0.007584f
C818 B.n778 VSUBS 0.007584f
C819 B.n779 VSUBS 0.007584f
C820 B.n780 VSUBS 0.007584f
C821 B.n781 VSUBS 0.007584f
C822 B.n782 VSUBS 0.007584f
C823 B.n783 VSUBS 0.007584f
C824 B.n784 VSUBS 0.007584f
C825 B.n785 VSUBS 0.007584f
C826 B.n786 VSUBS 0.007584f
C827 B.n787 VSUBS 0.007584f
C828 B.n788 VSUBS 0.007584f
C829 B.n789 VSUBS 0.007584f
C830 B.n790 VSUBS 0.007584f
C831 B.n791 VSUBS 0.007584f
C832 B.n792 VSUBS 0.007584f
C833 B.n793 VSUBS 0.007584f
C834 B.n794 VSUBS 0.007584f
C835 B.n795 VSUBS 0.007584f
C836 B.n796 VSUBS 0.007584f
C837 B.n797 VSUBS 0.007584f
C838 B.n798 VSUBS 0.007584f
C839 B.n799 VSUBS 0.007584f
C840 B.n800 VSUBS 0.007584f
C841 B.n801 VSUBS 0.007584f
C842 B.n802 VSUBS 0.007584f
C843 B.n803 VSUBS 0.007584f
C844 B.n804 VSUBS 0.007584f
C845 B.n805 VSUBS 0.007584f
C846 B.n806 VSUBS 0.007584f
C847 B.n807 VSUBS 0.007584f
C848 B.n808 VSUBS 0.007584f
C849 B.n809 VSUBS 0.007584f
C850 B.n810 VSUBS 0.007584f
C851 B.n811 VSUBS 0.007584f
C852 B.n812 VSUBS 0.007584f
C853 B.n813 VSUBS 0.007584f
C854 B.n814 VSUBS 0.007584f
C855 B.n815 VSUBS 0.007584f
C856 B.n816 VSUBS 0.007584f
C857 B.n817 VSUBS 0.007584f
C858 B.n818 VSUBS 0.007584f
C859 B.n819 VSUBS 0.007584f
C860 B.n820 VSUBS 0.007584f
C861 B.n821 VSUBS 0.007584f
C862 B.n822 VSUBS 0.007584f
C863 B.n823 VSUBS 0.007584f
C864 B.n824 VSUBS 0.007584f
C865 B.n825 VSUBS 0.007584f
C866 B.n826 VSUBS 0.007584f
C867 B.n827 VSUBS 0.007584f
C868 B.n828 VSUBS 0.007584f
C869 B.n829 VSUBS 0.007584f
C870 B.n830 VSUBS 0.007584f
C871 B.n831 VSUBS 0.007584f
C872 B.n832 VSUBS 0.018354f
C873 B.n833 VSUBS 0.018354f
C874 B.n834 VSUBS 0.01756f
C875 B.n835 VSUBS 0.007584f
C876 B.n836 VSUBS 0.007584f
C877 B.n837 VSUBS 0.007584f
C878 B.n838 VSUBS 0.007584f
C879 B.n839 VSUBS 0.007584f
C880 B.n840 VSUBS 0.007584f
C881 B.n841 VSUBS 0.007584f
C882 B.n842 VSUBS 0.007584f
C883 B.n843 VSUBS 0.007584f
C884 B.n844 VSUBS 0.007584f
C885 B.n845 VSUBS 0.007584f
C886 B.n846 VSUBS 0.007584f
C887 B.n847 VSUBS 0.007584f
C888 B.n848 VSUBS 0.007584f
C889 B.n849 VSUBS 0.007584f
C890 B.n850 VSUBS 0.007584f
C891 B.n851 VSUBS 0.007584f
C892 B.n852 VSUBS 0.007584f
C893 B.n853 VSUBS 0.007584f
C894 B.n854 VSUBS 0.007584f
C895 B.n855 VSUBS 0.007584f
C896 B.n856 VSUBS 0.007584f
C897 B.n857 VSUBS 0.007584f
C898 B.n858 VSUBS 0.007584f
C899 B.n859 VSUBS 0.007584f
C900 B.n860 VSUBS 0.007584f
C901 B.n861 VSUBS 0.007584f
C902 B.n862 VSUBS 0.007584f
C903 B.n863 VSUBS 0.007584f
C904 B.n864 VSUBS 0.007584f
C905 B.n865 VSUBS 0.007584f
C906 B.n866 VSUBS 0.007584f
C907 B.n867 VSUBS 0.007584f
C908 B.n868 VSUBS 0.007584f
C909 B.n869 VSUBS 0.007584f
C910 B.n870 VSUBS 0.007584f
C911 B.n871 VSUBS 0.007584f
C912 B.n872 VSUBS 0.007584f
C913 B.n873 VSUBS 0.007584f
C914 B.n874 VSUBS 0.007584f
C915 B.n875 VSUBS 0.007584f
C916 B.n876 VSUBS 0.007584f
C917 B.n877 VSUBS 0.007584f
C918 B.n878 VSUBS 0.007584f
C919 B.n879 VSUBS 0.007584f
C920 B.n880 VSUBS 0.007584f
C921 B.n881 VSUBS 0.007584f
C922 B.n882 VSUBS 0.007584f
C923 B.n883 VSUBS 0.007584f
C924 B.n884 VSUBS 0.007584f
C925 B.n885 VSUBS 0.007584f
C926 B.n886 VSUBS 0.007584f
C927 B.n887 VSUBS 0.007584f
C928 B.n888 VSUBS 0.007584f
C929 B.n889 VSUBS 0.007584f
C930 B.n890 VSUBS 0.007584f
C931 B.n891 VSUBS 0.007584f
C932 B.n892 VSUBS 0.007584f
C933 B.n893 VSUBS 0.007584f
C934 B.n894 VSUBS 0.007584f
C935 B.n895 VSUBS 0.007584f
C936 B.n896 VSUBS 0.007584f
C937 B.n897 VSUBS 0.007584f
C938 B.n898 VSUBS 0.007584f
C939 B.n899 VSUBS 0.007584f
C940 B.n900 VSUBS 0.007584f
C941 B.n901 VSUBS 0.007584f
C942 B.n902 VSUBS 0.007584f
C943 B.n903 VSUBS 0.007584f
C944 B.n904 VSUBS 0.007584f
C945 B.n905 VSUBS 0.007584f
C946 B.n906 VSUBS 0.007584f
C947 B.n907 VSUBS 0.007584f
C948 B.n908 VSUBS 0.007584f
C949 B.n909 VSUBS 0.007584f
C950 B.n910 VSUBS 0.007584f
C951 B.n911 VSUBS 0.007584f
C952 B.n912 VSUBS 0.007584f
C953 B.n913 VSUBS 0.007584f
C954 B.n914 VSUBS 0.007584f
C955 B.n915 VSUBS 0.009897f
C956 B.n916 VSUBS 0.010543f
C957 B.n917 VSUBS 0.020966f
C958 VDD1.t4 VSUBS 3.69658f
C959 VDD1.t2 VSUBS 3.69497f
C960 VDD1.t3 VSUBS 0.344687f
C961 VDD1.t0 VSUBS 0.344687f
C962 VDD1.n0 VSUBS 2.83215f
C963 VDD1.n1 VSUBS 4.78341f
C964 VDD1.t1 VSUBS 0.344687f
C965 VDD1.t5 VSUBS 0.344687f
C966 VDD1.n2 VSUBS 2.82176f
C967 VDD1.n3 VSUBS 4.04141f
C968 VP.t5 VSUBS 4.04577f
C969 VP.n0 VSUBS 1.49146f
C970 VP.n1 VSUBS 0.025243f
C971 VP.n2 VSUBS 0.049757f
C972 VP.n3 VSUBS 0.025243f
C973 VP.n4 VSUBS 0.047047f
C974 VP.n5 VSUBS 0.025243f
C975 VP.t2 VSUBS 4.04577f
C976 VP.n6 VSUBS 0.050514f
C977 VP.n7 VSUBS 0.025243f
C978 VP.n8 VSUBS 0.047047f
C979 VP.t0 VSUBS 4.04577f
C980 VP.n9 VSUBS 1.49146f
C981 VP.n10 VSUBS 0.025243f
C982 VP.n11 VSUBS 0.049757f
C983 VP.n12 VSUBS 0.025243f
C984 VP.n13 VSUBS 0.047047f
C985 VP.t1 VSUBS 4.430049f
C986 VP.t4 VSUBS 4.04577f
C987 VP.n14 VSUBS 1.50417f
C988 VP.n15 VSUBS 1.43333f
C989 VP.n16 VSUBS 0.322033f
C990 VP.n17 VSUBS 0.025243f
C991 VP.n18 VSUBS 0.047047f
C992 VP.n19 VSUBS 0.050514f
C993 VP.n20 VSUBS 0.020481f
C994 VP.n21 VSUBS 0.025243f
C995 VP.n22 VSUBS 0.025243f
C996 VP.n23 VSUBS 0.025243f
C997 VP.n24 VSUBS 0.047047f
C998 VP.n25 VSUBS 0.047047f
C999 VP.n26 VSUBS 0.025213f
C1000 VP.n27 VSUBS 0.040742f
C1001 VP.n28 VSUBS 1.69295f
C1002 VP.n29 VSUBS 1.7092f
C1003 VP.t3 VSUBS 4.04577f
C1004 VP.n30 VSUBS 1.49146f
C1005 VP.n31 VSUBS 0.025213f
C1006 VP.n32 VSUBS 0.040742f
C1007 VP.n33 VSUBS 0.025243f
C1008 VP.n34 VSUBS 0.025243f
C1009 VP.n35 VSUBS 0.047047f
C1010 VP.n36 VSUBS 0.049757f
C1011 VP.n37 VSUBS 0.020481f
C1012 VP.n38 VSUBS 0.025243f
C1013 VP.n39 VSUBS 0.025243f
C1014 VP.n40 VSUBS 0.025243f
C1015 VP.n41 VSUBS 0.047047f
C1016 VP.n42 VSUBS 0.047047f
C1017 VP.n43 VSUBS 1.42472f
C1018 VP.n44 VSUBS 0.025243f
C1019 VP.n45 VSUBS 0.025243f
C1020 VP.n46 VSUBS 0.025243f
C1021 VP.n47 VSUBS 0.047047f
C1022 VP.n48 VSUBS 0.050514f
C1023 VP.n49 VSUBS 0.020481f
C1024 VP.n50 VSUBS 0.025243f
C1025 VP.n51 VSUBS 0.025243f
C1026 VP.n52 VSUBS 0.025243f
C1027 VP.n53 VSUBS 0.047047f
C1028 VP.n54 VSUBS 0.047047f
C1029 VP.n55 VSUBS 0.025213f
C1030 VP.n56 VSUBS 0.040742f
C1031 VP.n57 VSUBS 0.077131f
C1032 VDD2.t2 VSUBS 3.69528f
C1033 VDD2.t0 VSUBS 0.344716f
C1034 VDD2.t5 VSUBS 0.344716f
C1035 VDD2.n0 VSUBS 2.83238f
C1036 VDD2.n1 VSUBS 4.61066f
C1037 VDD2.t1 VSUBS 3.66635f
C1038 VDD2.n2 VSUBS 4.06436f
C1039 VDD2.t4 VSUBS 0.344716f
C1040 VDD2.t3 VSUBS 0.344716f
C1041 VDD2.n3 VSUBS 2.83233f
C1042 VTAIL.t8 VSUBS 0.358789f
C1043 VTAIL.t10 VSUBS 0.358789f
C1044 VTAIL.n0 VSUBS 2.77122f
C1045 VTAIL.n1 VSUBS 0.967135f
C1046 VTAIL.t2 VSUBS 3.62674f
C1047 VTAIL.n2 VSUBS 1.32615f
C1048 VTAIL.t3 VSUBS 0.358789f
C1049 VTAIL.t4 VSUBS 0.358789f
C1050 VTAIL.n3 VSUBS 2.77122f
C1051 VTAIL.n4 VSUBS 3.29425f
C1052 VTAIL.t9 VSUBS 0.358789f
C1053 VTAIL.t6 VSUBS 0.358789f
C1054 VTAIL.n5 VSUBS 2.77122f
C1055 VTAIL.n6 VSUBS 3.29425f
C1056 VTAIL.t7 VSUBS 3.62677f
C1057 VTAIL.n7 VSUBS 1.32613f
C1058 VTAIL.t5 VSUBS 0.358789f
C1059 VTAIL.t0 VSUBS 0.358789f
C1060 VTAIL.n8 VSUBS 2.77122f
C1061 VTAIL.n9 VSUBS 1.20315f
C1062 VTAIL.t1 VSUBS 3.62674f
C1063 VTAIL.n10 VSUBS 3.09536f
C1064 VTAIL.t11 VSUBS 3.62674f
C1065 VTAIL.n11 VSUBS 3.0095f
C1066 VN.t0 VSUBS 3.70007f
C1067 VN.n0 VSUBS 1.36401f
C1068 VN.n1 VSUBS 0.023086f
C1069 VN.n2 VSUBS 0.045506f
C1070 VN.n3 VSUBS 0.023086f
C1071 VN.n4 VSUBS 0.043027f
C1072 VN.t5 VSUBS 3.70007f
C1073 VN.n5 VSUBS 1.37564f
C1074 VN.t3 VSUBS 4.05151f
C1075 VN.n6 VSUBS 1.31085f
C1076 VN.n7 VSUBS 0.294515f
C1077 VN.n8 VSUBS 0.023086f
C1078 VN.n9 VSUBS 0.043027f
C1079 VN.n10 VSUBS 0.046198f
C1080 VN.n11 VSUBS 0.018731f
C1081 VN.n12 VSUBS 0.023086f
C1082 VN.n13 VSUBS 0.023086f
C1083 VN.n14 VSUBS 0.023086f
C1084 VN.n15 VSUBS 0.043027f
C1085 VN.n16 VSUBS 0.043027f
C1086 VN.n17 VSUBS 0.023059f
C1087 VN.n18 VSUBS 0.037261f
C1088 VN.n19 VSUBS 0.07054f
C1089 VN.t4 VSUBS 3.70007f
C1090 VN.n20 VSUBS 1.36401f
C1091 VN.n21 VSUBS 0.023086f
C1092 VN.n22 VSUBS 0.045506f
C1093 VN.n23 VSUBS 0.023086f
C1094 VN.n24 VSUBS 0.043027f
C1095 VN.t2 VSUBS 4.05151f
C1096 VN.t1 VSUBS 3.70007f
C1097 VN.n25 VSUBS 1.37564f
C1098 VN.n26 VSUBS 1.31085f
C1099 VN.n27 VSUBS 0.294515f
C1100 VN.n28 VSUBS 0.023086f
C1101 VN.n29 VSUBS 0.043027f
C1102 VN.n30 VSUBS 0.046198f
C1103 VN.n31 VSUBS 0.018731f
C1104 VN.n32 VSUBS 0.023086f
C1105 VN.n33 VSUBS 0.023086f
C1106 VN.n34 VSUBS 0.023086f
C1107 VN.n35 VSUBS 0.043027f
C1108 VN.n36 VSUBS 0.043027f
C1109 VN.n37 VSUBS 0.023059f
C1110 VN.n38 VSUBS 0.037261f
C1111 VN.n39 VSUBS 1.5574f
.ends

