* NGSPICE file created from diff_pair_sample_1363.ext - technology: sky130A

.subckt diff_pair_sample_1363 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t7 VN.t0 VTAIL.t8 B.t0 sky130_fd_pr__nfet_01v8 ad=0.41745 pd=2.86 as=0.9867 ps=5.84 w=2.53 l=2.84
X1 VTAIL.t10 VN.t1 VDD2.t6 B.t3 sky130_fd_pr__nfet_01v8 ad=0.41745 pd=2.86 as=0.41745 ps=2.86 w=2.53 l=2.84
X2 VTAIL.t9 VN.t2 VDD2.t5 B.t1 sky130_fd_pr__nfet_01v8 ad=0.9867 pd=5.84 as=0.41745 ps=2.86 w=2.53 l=2.84
X3 VTAIL.t7 VP.t0 VDD1.t7 B.t7 sky130_fd_pr__nfet_01v8 ad=0.9867 pd=5.84 as=0.41745 ps=2.86 w=2.53 l=2.84
X4 VDD1.t6 VP.t1 VTAIL.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=0.41745 pd=2.86 as=0.41745 ps=2.86 w=2.53 l=2.84
X5 VDD2.t4 VN.t3 VTAIL.t14 B.t6 sky130_fd_pr__nfet_01v8 ad=0.41745 pd=2.86 as=0.41745 ps=2.86 w=2.53 l=2.84
X6 VTAIL.t4 VP.t2 VDD1.t5 B.t4 sky130_fd_pr__nfet_01v8 ad=0.41745 pd=2.86 as=0.41745 ps=2.86 w=2.53 l=2.84
X7 VTAIL.t3 VP.t3 VDD1.t4 B.t3 sky130_fd_pr__nfet_01v8 ad=0.41745 pd=2.86 as=0.41745 ps=2.86 w=2.53 l=2.84
X8 VDD1.t3 VP.t4 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=0.41745 pd=2.86 as=0.9867 ps=5.84 w=2.53 l=2.84
X9 B.t21 B.t19 B.t20 B.t13 sky130_fd_pr__nfet_01v8 ad=0.9867 pd=5.84 as=0 ps=0 w=2.53 l=2.84
X10 VDD2.t3 VN.t4 VTAIL.t15 B.t5 sky130_fd_pr__nfet_01v8 ad=0.41745 pd=2.86 as=0.41745 ps=2.86 w=2.53 l=2.84
X11 VTAIL.t12 VN.t5 VDD2.t2 B.t7 sky130_fd_pr__nfet_01v8 ad=0.9867 pd=5.84 as=0.41745 ps=2.86 w=2.53 l=2.84
X12 VDD2.t1 VN.t6 VTAIL.t11 B.t2 sky130_fd_pr__nfet_01v8 ad=0.41745 pd=2.86 as=0.9867 ps=5.84 w=2.53 l=2.84
X13 VDD1.t2 VP.t5 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=0.41745 pd=2.86 as=0.9867 ps=5.84 w=2.53 l=2.84
X14 VTAIL.t13 VN.t7 VDD2.t0 B.t4 sky130_fd_pr__nfet_01v8 ad=0.41745 pd=2.86 as=0.41745 ps=2.86 w=2.53 l=2.84
X15 B.t18 B.t16 B.t17 B.t9 sky130_fd_pr__nfet_01v8 ad=0.9867 pd=5.84 as=0 ps=0 w=2.53 l=2.84
X16 VTAIL.t1 VP.t6 VDD1.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=0.9867 pd=5.84 as=0.41745 ps=2.86 w=2.53 l=2.84
X17 B.t15 B.t12 B.t14 B.t13 sky130_fd_pr__nfet_01v8 ad=0.9867 pd=5.84 as=0 ps=0 w=2.53 l=2.84
X18 VDD1.t0 VP.t7 VTAIL.t6 B.t6 sky130_fd_pr__nfet_01v8 ad=0.41745 pd=2.86 as=0.41745 ps=2.86 w=2.53 l=2.84
X19 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=0.9867 pd=5.84 as=0 ps=0 w=2.53 l=2.84
R0 VN.n59 VN.n31 161.3
R1 VN.n58 VN.n57 161.3
R2 VN.n56 VN.n32 161.3
R3 VN.n55 VN.n54 161.3
R4 VN.n53 VN.n33 161.3
R5 VN.n52 VN.n51 161.3
R6 VN.n50 VN.n34 161.3
R7 VN.n49 VN.n48 161.3
R8 VN.n47 VN.n35 161.3
R9 VN.n46 VN.n45 161.3
R10 VN.n44 VN.n37 161.3
R11 VN.n43 VN.n42 161.3
R12 VN.n41 VN.n38 161.3
R13 VN.n28 VN.n0 161.3
R14 VN.n27 VN.n26 161.3
R15 VN.n25 VN.n1 161.3
R16 VN.n24 VN.n23 161.3
R17 VN.n22 VN.n2 161.3
R18 VN.n21 VN.n20 161.3
R19 VN.n19 VN.n3 161.3
R20 VN.n18 VN.n17 161.3
R21 VN.n15 VN.n4 161.3
R22 VN.n14 VN.n13 161.3
R23 VN.n12 VN.n5 161.3
R24 VN.n11 VN.n10 161.3
R25 VN.n9 VN.n6 161.3
R26 VN.n30 VN.n29 110.511
R27 VN.n61 VN.n60 110.511
R28 VN.n8 VN.n7 57.3183
R29 VN.n40 VN.n39 57.3183
R30 VN.n14 VN.n5 56.5193
R31 VN.n46 VN.n37 56.5193
R32 VN.n7 VN.t5 53.5387
R33 VN.n39 VN.t6 53.5387
R34 VN.n23 VN.n22 48.2635
R35 VN.n54 VN.n53 48.2635
R36 VN VN.n61 45.0512
R37 VN.n23 VN.n1 32.7233
R38 VN.n54 VN.n32 32.7233
R39 VN.n10 VN.n9 24.4675
R40 VN.n10 VN.n5 24.4675
R41 VN.n15 VN.n14 24.4675
R42 VN.n17 VN.n15 24.4675
R43 VN.n21 VN.n3 24.4675
R44 VN.n22 VN.n21 24.4675
R45 VN.n27 VN.n1 24.4675
R46 VN.n28 VN.n27 24.4675
R47 VN.n42 VN.n37 24.4675
R48 VN.n42 VN.n41 24.4675
R49 VN.n53 VN.n52 24.4675
R50 VN.n52 VN.n34 24.4675
R51 VN.n48 VN.n47 24.4675
R52 VN.n47 VN.n46 24.4675
R53 VN.n59 VN.n58 24.4675
R54 VN.n58 VN.n32 24.4675
R55 VN.n8 VN.t4 21.4699
R56 VN.n16 VN.t1 21.4699
R57 VN.n29 VN.t0 21.4699
R58 VN.n40 VN.t7 21.4699
R59 VN.n36 VN.t3 21.4699
R60 VN.n60 VN.t2 21.4699
R61 VN.n9 VN.n8 16.3934
R62 VN.n17 VN.n16 16.3934
R63 VN.n41 VN.n40 16.3934
R64 VN.n48 VN.n36 16.3934
R65 VN.n16 VN.n3 8.07461
R66 VN.n36 VN.n34 8.07461
R67 VN.n39 VN.n38 5.19262
R68 VN.n7 VN.n6 5.19262
R69 VN.n61 VN.n31 0.278367
R70 VN.n30 VN.n0 0.278367
R71 VN.n29 VN.n28 0.24517
R72 VN.n60 VN.n59 0.24517
R73 VN.n57 VN.n31 0.189894
R74 VN.n57 VN.n56 0.189894
R75 VN.n56 VN.n55 0.189894
R76 VN.n55 VN.n33 0.189894
R77 VN.n51 VN.n33 0.189894
R78 VN.n51 VN.n50 0.189894
R79 VN.n50 VN.n49 0.189894
R80 VN.n49 VN.n35 0.189894
R81 VN.n45 VN.n35 0.189894
R82 VN.n45 VN.n44 0.189894
R83 VN.n44 VN.n43 0.189894
R84 VN.n43 VN.n38 0.189894
R85 VN.n11 VN.n6 0.189894
R86 VN.n12 VN.n11 0.189894
R87 VN.n13 VN.n12 0.189894
R88 VN.n13 VN.n4 0.189894
R89 VN.n18 VN.n4 0.189894
R90 VN.n19 VN.n18 0.189894
R91 VN.n20 VN.n19 0.189894
R92 VN.n20 VN.n2 0.189894
R93 VN.n24 VN.n2 0.189894
R94 VN.n25 VN.n24 0.189894
R95 VN.n26 VN.n25 0.189894
R96 VN.n26 VN.n0 0.189894
R97 VN VN.n30 0.153454
R98 VTAIL.n98 VTAIL.n92 289.615
R99 VTAIL.n8 VTAIL.n2 289.615
R100 VTAIL.n20 VTAIL.n14 289.615
R101 VTAIL.n34 VTAIL.n28 289.615
R102 VTAIL.n86 VTAIL.n80 289.615
R103 VTAIL.n72 VTAIL.n66 289.615
R104 VTAIL.n60 VTAIL.n54 289.615
R105 VTAIL.n46 VTAIL.n40 289.615
R106 VTAIL.n97 VTAIL.n96 185
R107 VTAIL.n99 VTAIL.n98 185
R108 VTAIL.n7 VTAIL.n6 185
R109 VTAIL.n9 VTAIL.n8 185
R110 VTAIL.n19 VTAIL.n18 185
R111 VTAIL.n21 VTAIL.n20 185
R112 VTAIL.n33 VTAIL.n32 185
R113 VTAIL.n35 VTAIL.n34 185
R114 VTAIL.n87 VTAIL.n86 185
R115 VTAIL.n85 VTAIL.n84 185
R116 VTAIL.n73 VTAIL.n72 185
R117 VTAIL.n71 VTAIL.n70 185
R118 VTAIL.n61 VTAIL.n60 185
R119 VTAIL.n59 VTAIL.n58 185
R120 VTAIL.n47 VTAIL.n46 185
R121 VTAIL.n45 VTAIL.n44 185
R122 VTAIL.n95 VTAIL.t8 151.613
R123 VTAIL.n5 VTAIL.t12 151.613
R124 VTAIL.n17 VTAIL.t2 151.613
R125 VTAIL.n31 VTAIL.t1 151.613
R126 VTAIL.n83 VTAIL.t0 151.613
R127 VTAIL.n69 VTAIL.t7 151.613
R128 VTAIL.n57 VTAIL.t11 151.613
R129 VTAIL.n43 VTAIL.t9 151.613
R130 VTAIL.n98 VTAIL.n97 104.615
R131 VTAIL.n8 VTAIL.n7 104.615
R132 VTAIL.n20 VTAIL.n19 104.615
R133 VTAIL.n34 VTAIL.n33 104.615
R134 VTAIL.n86 VTAIL.n85 104.615
R135 VTAIL.n72 VTAIL.n71 104.615
R136 VTAIL.n60 VTAIL.n59 104.615
R137 VTAIL.n46 VTAIL.n45 104.615
R138 VTAIL.n79 VTAIL.n78 70.8017
R139 VTAIL.n53 VTAIL.n52 70.8017
R140 VTAIL.n1 VTAIL.n0 70.8016
R141 VTAIL.n27 VTAIL.n26 70.8016
R142 VTAIL.n97 VTAIL.t8 52.3082
R143 VTAIL.n7 VTAIL.t12 52.3082
R144 VTAIL.n19 VTAIL.t2 52.3082
R145 VTAIL.n33 VTAIL.t1 52.3082
R146 VTAIL.n85 VTAIL.t0 52.3082
R147 VTAIL.n71 VTAIL.t7 52.3082
R148 VTAIL.n59 VTAIL.t11 52.3082
R149 VTAIL.n45 VTAIL.t9 52.3082
R150 VTAIL.n103 VTAIL.n102 34.7066
R151 VTAIL.n13 VTAIL.n12 34.7066
R152 VTAIL.n25 VTAIL.n24 34.7066
R153 VTAIL.n39 VTAIL.n38 34.7066
R154 VTAIL.n91 VTAIL.n90 34.7066
R155 VTAIL.n77 VTAIL.n76 34.7066
R156 VTAIL.n65 VTAIL.n64 34.7066
R157 VTAIL.n51 VTAIL.n50 34.7066
R158 VTAIL.n103 VTAIL.n91 17.2807
R159 VTAIL.n51 VTAIL.n39 17.2807
R160 VTAIL.n96 VTAIL.n95 15.3979
R161 VTAIL.n6 VTAIL.n5 15.3979
R162 VTAIL.n18 VTAIL.n17 15.3979
R163 VTAIL.n32 VTAIL.n31 15.3979
R164 VTAIL.n84 VTAIL.n83 15.3979
R165 VTAIL.n70 VTAIL.n69 15.3979
R166 VTAIL.n58 VTAIL.n57 15.3979
R167 VTAIL.n44 VTAIL.n43 15.3979
R168 VTAIL.n99 VTAIL.n94 12.8005
R169 VTAIL.n9 VTAIL.n4 12.8005
R170 VTAIL.n21 VTAIL.n16 12.8005
R171 VTAIL.n35 VTAIL.n30 12.8005
R172 VTAIL.n87 VTAIL.n82 12.8005
R173 VTAIL.n73 VTAIL.n68 12.8005
R174 VTAIL.n61 VTAIL.n56 12.8005
R175 VTAIL.n47 VTAIL.n42 12.8005
R176 VTAIL.n100 VTAIL.n92 12.0247
R177 VTAIL.n10 VTAIL.n2 12.0247
R178 VTAIL.n22 VTAIL.n14 12.0247
R179 VTAIL.n36 VTAIL.n28 12.0247
R180 VTAIL.n88 VTAIL.n80 12.0247
R181 VTAIL.n74 VTAIL.n66 12.0247
R182 VTAIL.n62 VTAIL.n54 12.0247
R183 VTAIL.n48 VTAIL.n40 12.0247
R184 VTAIL.n102 VTAIL.n101 9.45567
R185 VTAIL.n12 VTAIL.n11 9.45567
R186 VTAIL.n24 VTAIL.n23 9.45567
R187 VTAIL.n38 VTAIL.n37 9.45567
R188 VTAIL.n90 VTAIL.n89 9.45567
R189 VTAIL.n76 VTAIL.n75 9.45567
R190 VTAIL.n64 VTAIL.n63 9.45567
R191 VTAIL.n50 VTAIL.n49 9.45567
R192 VTAIL.n101 VTAIL.n100 9.3005
R193 VTAIL.n94 VTAIL.n93 9.3005
R194 VTAIL.n11 VTAIL.n10 9.3005
R195 VTAIL.n4 VTAIL.n3 9.3005
R196 VTAIL.n23 VTAIL.n22 9.3005
R197 VTAIL.n16 VTAIL.n15 9.3005
R198 VTAIL.n37 VTAIL.n36 9.3005
R199 VTAIL.n30 VTAIL.n29 9.3005
R200 VTAIL.n89 VTAIL.n88 9.3005
R201 VTAIL.n82 VTAIL.n81 9.3005
R202 VTAIL.n75 VTAIL.n74 9.3005
R203 VTAIL.n68 VTAIL.n67 9.3005
R204 VTAIL.n63 VTAIL.n62 9.3005
R205 VTAIL.n56 VTAIL.n55 9.3005
R206 VTAIL.n49 VTAIL.n48 9.3005
R207 VTAIL.n42 VTAIL.n41 9.3005
R208 VTAIL.n0 VTAIL.t15 7.82659
R209 VTAIL.n0 VTAIL.t10 7.82659
R210 VTAIL.n26 VTAIL.t6 7.82659
R211 VTAIL.n26 VTAIL.t4 7.82659
R212 VTAIL.n78 VTAIL.t5 7.82659
R213 VTAIL.n78 VTAIL.t3 7.82659
R214 VTAIL.n52 VTAIL.t14 7.82659
R215 VTAIL.n52 VTAIL.t13 7.82659
R216 VTAIL.n95 VTAIL.n93 4.69785
R217 VTAIL.n5 VTAIL.n3 4.69785
R218 VTAIL.n17 VTAIL.n15 4.69785
R219 VTAIL.n31 VTAIL.n29 4.69785
R220 VTAIL.n83 VTAIL.n81 4.69785
R221 VTAIL.n69 VTAIL.n67 4.69785
R222 VTAIL.n57 VTAIL.n55 4.69785
R223 VTAIL.n43 VTAIL.n41 4.69785
R224 VTAIL.n53 VTAIL.n51 2.73326
R225 VTAIL.n65 VTAIL.n53 2.73326
R226 VTAIL.n79 VTAIL.n77 2.73326
R227 VTAIL.n91 VTAIL.n79 2.73326
R228 VTAIL.n39 VTAIL.n27 2.73326
R229 VTAIL.n27 VTAIL.n25 2.73326
R230 VTAIL.n13 VTAIL.n1 2.73326
R231 VTAIL VTAIL.n103 2.67507
R232 VTAIL.n102 VTAIL.n92 1.93989
R233 VTAIL.n12 VTAIL.n2 1.93989
R234 VTAIL.n24 VTAIL.n14 1.93989
R235 VTAIL.n38 VTAIL.n28 1.93989
R236 VTAIL.n90 VTAIL.n80 1.93989
R237 VTAIL.n76 VTAIL.n66 1.93989
R238 VTAIL.n64 VTAIL.n54 1.93989
R239 VTAIL.n50 VTAIL.n40 1.93989
R240 VTAIL.n100 VTAIL.n99 1.16414
R241 VTAIL.n10 VTAIL.n9 1.16414
R242 VTAIL.n22 VTAIL.n21 1.16414
R243 VTAIL.n36 VTAIL.n35 1.16414
R244 VTAIL.n88 VTAIL.n87 1.16414
R245 VTAIL.n74 VTAIL.n73 1.16414
R246 VTAIL.n62 VTAIL.n61 1.16414
R247 VTAIL.n48 VTAIL.n47 1.16414
R248 VTAIL.n77 VTAIL.n65 0.470328
R249 VTAIL.n25 VTAIL.n13 0.470328
R250 VTAIL.n96 VTAIL.n94 0.388379
R251 VTAIL.n6 VTAIL.n4 0.388379
R252 VTAIL.n18 VTAIL.n16 0.388379
R253 VTAIL.n32 VTAIL.n30 0.388379
R254 VTAIL.n84 VTAIL.n82 0.388379
R255 VTAIL.n70 VTAIL.n68 0.388379
R256 VTAIL.n58 VTAIL.n56 0.388379
R257 VTAIL.n44 VTAIL.n42 0.388379
R258 VTAIL.n101 VTAIL.n93 0.155672
R259 VTAIL.n11 VTAIL.n3 0.155672
R260 VTAIL.n23 VTAIL.n15 0.155672
R261 VTAIL.n37 VTAIL.n29 0.155672
R262 VTAIL.n89 VTAIL.n81 0.155672
R263 VTAIL.n75 VTAIL.n67 0.155672
R264 VTAIL.n63 VTAIL.n55 0.155672
R265 VTAIL.n49 VTAIL.n41 0.155672
R266 VTAIL VTAIL.n1 0.0586897
R267 VDD2.n2 VDD2.n1 88.7914
R268 VDD2.n2 VDD2.n0 88.7914
R269 VDD2 VDD2.n5 88.7886
R270 VDD2.n4 VDD2.n3 87.4805
R271 VDD2.n4 VDD2.n2 38.1937
R272 VDD2.n5 VDD2.t0 7.82659
R273 VDD2.n5 VDD2.t1 7.82659
R274 VDD2.n3 VDD2.t5 7.82659
R275 VDD2.n3 VDD2.t4 7.82659
R276 VDD2.n1 VDD2.t6 7.82659
R277 VDD2.n1 VDD2.t7 7.82659
R278 VDD2.n0 VDD2.t2 7.82659
R279 VDD2.n0 VDD2.t3 7.82659
R280 VDD2 VDD2.n4 1.42507
R281 B.n561 B.n560 585
R282 B.n561 B.n100 585
R283 B.n564 B.n563 585
R284 B.n565 B.n123 585
R285 B.n567 B.n566 585
R286 B.n569 B.n122 585
R287 B.n572 B.n571 585
R288 B.n573 B.n121 585
R289 B.n575 B.n574 585
R290 B.n577 B.n120 585
R291 B.n580 B.n579 585
R292 B.n581 B.n119 585
R293 B.n583 B.n582 585
R294 B.n585 B.n118 585
R295 B.n588 B.n587 585
R296 B.n590 B.n115 585
R297 B.n592 B.n591 585
R298 B.n594 B.n114 585
R299 B.n597 B.n596 585
R300 B.n598 B.n113 585
R301 B.n600 B.n599 585
R302 B.n602 B.n112 585
R303 B.n604 B.n603 585
R304 B.n606 B.n605 585
R305 B.n609 B.n608 585
R306 B.n610 B.n107 585
R307 B.n612 B.n611 585
R308 B.n614 B.n106 585
R309 B.n617 B.n616 585
R310 B.n618 B.n105 585
R311 B.n620 B.n619 585
R312 B.n622 B.n104 585
R313 B.n625 B.n624 585
R314 B.n626 B.n103 585
R315 B.n628 B.n627 585
R316 B.n630 B.n102 585
R317 B.n633 B.n632 585
R318 B.n634 B.n101 585
R319 B.n559 B.n99 585
R320 B.n637 B.n99 585
R321 B.n558 B.n98 585
R322 B.n638 B.n98 585
R323 B.n557 B.n97 585
R324 B.n639 B.n97 585
R325 B.n556 B.n555 585
R326 B.n555 B.n93 585
R327 B.n554 B.n92 585
R328 B.n645 B.n92 585
R329 B.n553 B.n91 585
R330 B.n646 B.n91 585
R331 B.n552 B.n90 585
R332 B.n647 B.n90 585
R333 B.n551 B.n550 585
R334 B.n550 B.n89 585
R335 B.n549 B.n85 585
R336 B.n653 B.n85 585
R337 B.n548 B.n84 585
R338 B.n654 B.n84 585
R339 B.n547 B.n83 585
R340 B.n655 B.n83 585
R341 B.n546 B.n545 585
R342 B.n545 B.n79 585
R343 B.n544 B.n78 585
R344 B.n661 B.n78 585
R345 B.n543 B.n77 585
R346 B.n662 B.n77 585
R347 B.n542 B.n76 585
R348 B.n663 B.n76 585
R349 B.n541 B.n540 585
R350 B.n540 B.n72 585
R351 B.n539 B.n71 585
R352 B.n669 B.n71 585
R353 B.n538 B.n70 585
R354 B.n670 B.n70 585
R355 B.n537 B.n69 585
R356 B.n671 B.n69 585
R357 B.n536 B.n535 585
R358 B.n535 B.n65 585
R359 B.n534 B.n64 585
R360 B.n677 B.n64 585
R361 B.n533 B.n63 585
R362 B.n678 B.n63 585
R363 B.n532 B.n62 585
R364 B.n679 B.n62 585
R365 B.n531 B.n530 585
R366 B.n530 B.n58 585
R367 B.n529 B.n57 585
R368 B.n685 B.n57 585
R369 B.n528 B.n56 585
R370 B.n686 B.n56 585
R371 B.n527 B.n55 585
R372 B.n687 B.n55 585
R373 B.n526 B.n525 585
R374 B.n525 B.n51 585
R375 B.n524 B.n50 585
R376 B.n693 B.n50 585
R377 B.n523 B.n49 585
R378 B.n694 B.n49 585
R379 B.n522 B.n48 585
R380 B.n695 B.n48 585
R381 B.n521 B.n520 585
R382 B.n520 B.n44 585
R383 B.n519 B.n43 585
R384 B.n701 B.n43 585
R385 B.n518 B.n42 585
R386 B.n702 B.n42 585
R387 B.n517 B.n41 585
R388 B.n703 B.n41 585
R389 B.n516 B.n515 585
R390 B.n515 B.n37 585
R391 B.n514 B.n36 585
R392 B.n709 B.n36 585
R393 B.n513 B.n35 585
R394 B.n710 B.n35 585
R395 B.n512 B.n34 585
R396 B.n711 B.n34 585
R397 B.n511 B.n510 585
R398 B.n510 B.n30 585
R399 B.n509 B.n29 585
R400 B.n717 B.n29 585
R401 B.n508 B.n28 585
R402 B.n718 B.n28 585
R403 B.n507 B.n27 585
R404 B.n719 B.n27 585
R405 B.n506 B.n505 585
R406 B.n505 B.n23 585
R407 B.n504 B.n22 585
R408 B.n725 B.n22 585
R409 B.n503 B.n21 585
R410 B.n726 B.n21 585
R411 B.n502 B.n20 585
R412 B.n727 B.n20 585
R413 B.n501 B.n500 585
R414 B.n500 B.n16 585
R415 B.n499 B.n15 585
R416 B.n733 B.n15 585
R417 B.n498 B.n14 585
R418 B.n734 B.n14 585
R419 B.n497 B.n13 585
R420 B.n735 B.n13 585
R421 B.n496 B.n495 585
R422 B.n495 B.n12 585
R423 B.n494 B.n493 585
R424 B.n494 B.n8 585
R425 B.n492 B.n7 585
R426 B.n742 B.n7 585
R427 B.n491 B.n6 585
R428 B.n743 B.n6 585
R429 B.n490 B.n5 585
R430 B.n744 B.n5 585
R431 B.n489 B.n488 585
R432 B.n488 B.n4 585
R433 B.n487 B.n124 585
R434 B.n487 B.n486 585
R435 B.n477 B.n125 585
R436 B.n126 B.n125 585
R437 B.n479 B.n478 585
R438 B.n480 B.n479 585
R439 B.n476 B.n131 585
R440 B.n131 B.n130 585
R441 B.n475 B.n474 585
R442 B.n474 B.n473 585
R443 B.n133 B.n132 585
R444 B.n134 B.n133 585
R445 B.n466 B.n465 585
R446 B.n467 B.n466 585
R447 B.n464 B.n139 585
R448 B.n139 B.n138 585
R449 B.n463 B.n462 585
R450 B.n462 B.n461 585
R451 B.n141 B.n140 585
R452 B.n142 B.n141 585
R453 B.n454 B.n453 585
R454 B.n455 B.n454 585
R455 B.n452 B.n147 585
R456 B.n147 B.n146 585
R457 B.n451 B.n450 585
R458 B.n450 B.n449 585
R459 B.n149 B.n148 585
R460 B.n150 B.n149 585
R461 B.n442 B.n441 585
R462 B.n443 B.n442 585
R463 B.n440 B.n155 585
R464 B.n155 B.n154 585
R465 B.n439 B.n438 585
R466 B.n438 B.n437 585
R467 B.n157 B.n156 585
R468 B.n158 B.n157 585
R469 B.n430 B.n429 585
R470 B.n431 B.n430 585
R471 B.n428 B.n163 585
R472 B.n163 B.n162 585
R473 B.n427 B.n426 585
R474 B.n426 B.n425 585
R475 B.n165 B.n164 585
R476 B.n166 B.n165 585
R477 B.n418 B.n417 585
R478 B.n419 B.n418 585
R479 B.n416 B.n170 585
R480 B.n174 B.n170 585
R481 B.n415 B.n414 585
R482 B.n414 B.n413 585
R483 B.n172 B.n171 585
R484 B.n173 B.n172 585
R485 B.n406 B.n405 585
R486 B.n407 B.n406 585
R487 B.n404 B.n179 585
R488 B.n179 B.n178 585
R489 B.n403 B.n402 585
R490 B.n402 B.n401 585
R491 B.n181 B.n180 585
R492 B.n182 B.n181 585
R493 B.n394 B.n393 585
R494 B.n395 B.n394 585
R495 B.n392 B.n187 585
R496 B.n187 B.n186 585
R497 B.n391 B.n390 585
R498 B.n390 B.n389 585
R499 B.n189 B.n188 585
R500 B.n190 B.n189 585
R501 B.n382 B.n381 585
R502 B.n383 B.n382 585
R503 B.n380 B.n195 585
R504 B.n195 B.n194 585
R505 B.n379 B.n378 585
R506 B.n378 B.n377 585
R507 B.n197 B.n196 585
R508 B.n198 B.n197 585
R509 B.n370 B.n369 585
R510 B.n371 B.n370 585
R511 B.n368 B.n203 585
R512 B.n203 B.n202 585
R513 B.n367 B.n366 585
R514 B.n366 B.n365 585
R515 B.n205 B.n204 585
R516 B.n206 B.n205 585
R517 B.n358 B.n357 585
R518 B.n359 B.n358 585
R519 B.n356 B.n211 585
R520 B.n211 B.n210 585
R521 B.n355 B.n354 585
R522 B.n354 B.n353 585
R523 B.n213 B.n212 585
R524 B.n346 B.n213 585
R525 B.n345 B.n344 585
R526 B.n347 B.n345 585
R527 B.n343 B.n218 585
R528 B.n218 B.n217 585
R529 B.n342 B.n341 585
R530 B.n341 B.n340 585
R531 B.n220 B.n219 585
R532 B.n221 B.n220 585
R533 B.n333 B.n332 585
R534 B.n334 B.n333 585
R535 B.n331 B.n226 585
R536 B.n226 B.n225 585
R537 B.n330 B.n329 585
R538 B.n329 B.n328 585
R539 B.n325 B.n230 585
R540 B.n324 B.n323 585
R541 B.n321 B.n231 585
R542 B.n321 B.n229 585
R543 B.n320 B.n319 585
R544 B.n318 B.n317 585
R545 B.n316 B.n233 585
R546 B.n314 B.n313 585
R547 B.n312 B.n234 585
R548 B.n311 B.n310 585
R549 B.n308 B.n235 585
R550 B.n306 B.n305 585
R551 B.n304 B.n236 585
R552 B.n303 B.n302 585
R553 B.n300 B.n237 585
R554 B.n298 B.n297 585
R555 B.n296 B.n238 585
R556 B.n295 B.n294 585
R557 B.n292 B.n242 585
R558 B.n290 B.n289 585
R559 B.n288 B.n243 585
R560 B.n287 B.n286 585
R561 B.n284 B.n244 585
R562 B.n282 B.n281 585
R563 B.n279 B.n245 585
R564 B.n278 B.n277 585
R565 B.n275 B.n248 585
R566 B.n273 B.n272 585
R567 B.n271 B.n249 585
R568 B.n270 B.n269 585
R569 B.n267 B.n250 585
R570 B.n265 B.n264 585
R571 B.n263 B.n251 585
R572 B.n262 B.n261 585
R573 B.n259 B.n252 585
R574 B.n257 B.n256 585
R575 B.n255 B.n254 585
R576 B.n228 B.n227 585
R577 B.n327 B.n326 585
R578 B.n328 B.n327 585
R579 B.n224 B.n223 585
R580 B.n225 B.n224 585
R581 B.n336 B.n335 585
R582 B.n335 B.n334 585
R583 B.n337 B.n222 585
R584 B.n222 B.n221 585
R585 B.n339 B.n338 585
R586 B.n340 B.n339 585
R587 B.n216 B.n215 585
R588 B.n217 B.n216 585
R589 B.n349 B.n348 585
R590 B.n348 B.n347 585
R591 B.n350 B.n214 585
R592 B.n346 B.n214 585
R593 B.n352 B.n351 585
R594 B.n353 B.n352 585
R595 B.n209 B.n208 585
R596 B.n210 B.n209 585
R597 B.n361 B.n360 585
R598 B.n360 B.n359 585
R599 B.n362 B.n207 585
R600 B.n207 B.n206 585
R601 B.n364 B.n363 585
R602 B.n365 B.n364 585
R603 B.n201 B.n200 585
R604 B.n202 B.n201 585
R605 B.n373 B.n372 585
R606 B.n372 B.n371 585
R607 B.n374 B.n199 585
R608 B.n199 B.n198 585
R609 B.n376 B.n375 585
R610 B.n377 B.n376 585
R611 B.n193 B.n192 585
R612 B.n194 B.n193 585
R613 B.n385 B.n384 585
R614 B.n384 B.n383 585
R615 B.n386 B.n191 585
R616 B.n191 B.n190 585
R617 B.n388 B.n387 585
R618 B.n389 B.n388 585
R619 B.n185 B.n184 585
R620 B.n186 B.n185 585
R621 B.n397 B.n396 585
R622 B.n396 B.n395 585
R623 B.n398 B.n183 585
R624 B.n183 B.n182 585
R625 B.n400 B.n399 585
R626 B.n401 B.n400 585
R627 B.n177 B.n176 585
R628 B.n178 B.n177 585
R629 B.n409 B.n408 585
R630 B.n408 B.n407 585
R631 B.n410 B.n175 585
R632 B.n175 B.n173 585
R633 B.n412 B.n411 585
R634 B.n413 B.n412 585
R635 B.n169 B.n168 585
R636 B.n174 B.n169 585
R637 B.n421 B.n420 585
R638 B.n420 B.n419 585
R639 B.n422 B.n167 585
R640 B.n167 B.n166 585
R641 B.n424 B.n423 585
R642 B.n425 B.n424 585
R643 B.n161 B.n160 585
R644 B.n162 B.n161 585
R645 B.n433 B.n432 585
R646 B.n432 B.n431 585
R647 B.n434 B.n159 585
R648 B.n159 B.n158 585
R649 B.n436 B.n435 585
R650 B.n437 B.n436 585
R651 B.n153 B.n152 585
R652 B.n154 B.n153 585
R653 B.n445 B.n444 585
R654 B.n444 B.n443 585
R655 B.n446 B.n151 585
R656 B.n151 B.n150 585
R657 B.n448 B.n447 585
R658 B.n449 B.n448 585
R659 B.n145 B.n144 585
R660 B.n146 B.n145 585
R661 B.n457 B.n456 585
R662 B.n456 B.n455 585
R663 B.n458 B.n143 585
R664 B.n143 B.n142 585
R665 B.n460 B.n459 585
R666 B.n461 B.n460 585
R667 B.n137 B.n136 585
R668 B.n138 B.n137 585
R669 B.n469 B.n468 585
R670 B.n468 B.n467 585
R671 B.n470 B.n135 585
R672 B.n135 B.n134 585
R673 B.n472 B.n471 585
R674 B.n473 B.n472 585
R675 B.n129 B.n128 585
R676 B.n130 B.n129 585
R677 B.n482 B.n481 585
R678 B.n481 B.n480 585
R679 B.n483 B.n127 585
R680 B.n127 B.n126 585
R681 B.n485 B.n484 585
R682 B.n486 B.n485 585
R683 B.n3 B.n0 585
R684 B.n4 B.n3 585
R685 B.n741 B.n1 585
R686 B.n742 B.n741 585
R687 B.n740 B.n739 585
R688 B.n740 B.n8 585
R689 B.n738 B.n9 585
R690 B.n12 B.n9 585
R691 B.n737 B.n736 585
R692 B.n736 B.n735 585
R693 B.n11 B.n10 585
R694 B.n734 B.n11 585
R695 B.n732 B.n731 585
R696 B.n733 B.n732 585
R697 B.n730 B.n17 585
R698 B.n17 B.n16 585
R699 B.n729 B.n728 585
R700 B.n728 B.n727 585
R701 B.n19 B.n18 585
R702 B.n726 B.n19 585
R703 B.n724 B.n723 585
R704 B.n725 B.n724 585
R705 B.n722 B.n24 585
R706 B.n24 B.n23 585
R707 B.n721 B.n720 585
R708 B.n720 B.n719 585
R709 B.n26 B.n25 585
R710 B.n718 B.n26 585
R711 B.n716 B.n715 585
R712 B.n717 B.n716 585
R713 B.n714 B.n31 585
R714 B.n31 B.n30 585
R715 B.n713 B.n712 585
R716 B.n712 B.n711 585
R717 B.n33 B.n32 585
R718 B.n710 B.n33 585
R719 B.n708 B.n707 585
R720 B.n709 B.n708 585
R721 B.n706 B.n38 585
R722 B.n38 B.n37 585
R723 B.n705 B.n704 585
R724 B.n704 B.n703 585
R725 B.n40 B.n39 585
R726 B.n702 B.n40 585
R727 B.n700 B.n699 585
R728 B.n701 B.n700 585
R729 B.n698 B.n45 585
R730 B.n45 B.n44 585
R731 B.n697 B.n696 585
R732 B.n696 B.n695 585
R733 B.n47 B.n46 585
R734 B.n694 B.n47 585
R735 B.n692 B.n691 585
R736 B.n693 B.n692 585
R737 B.n690 B.n52 585
R738 B.n52 B.n51 585
R739 B.n689 B.n688 585
R740 B.n688 B.n687 585
R741 B.n54 B.n53 585
R742 B.n686 B.n54 585
R743 B.n684 B.n683 585
R744 B.n685 B.n684 585
R745 B.n682 B.n59 585
R746 B.n59 B.n58 585
R747 B.n681 B.n680 585
R748 B.n680 B.n679 585
R749 B.n61 B.n60 585
R750 B.n678 B.n61 585
R751 B.n676 B.n675 585
R752 B.n677 B.n676 585
R753 B.n674 B.n66 585
R754 B.n66 B.n65 585
R755 B.n673 B.n672 585
R756 B.n672 B.n671 585
R757 B.n68 B.n67 585
R758 B.n670 B.n68 585
R759 B.n668 B.n667 585
R760 B.n669 B.n668 585
R761 B.n666 B.n73 585
R762 B.n73 B.n72 585
R763 B.n665 B.n664 585
R764 B.n664 B.n663 585
R765 B.n75 B.n74 585
R766 B.n662 B.n75 585
R767 B.n660 B.n659 585
R768 B.n661 B.n660 585
R769 B.n658 B.n80 585
R770 B.n80 B.n79 585
R771 B.n657 B.n656 585
R772 B.n656 B.n655 585
R773 B.n82 B.n81 585
R774 B.n654 B.n82 585
R775 B.n652 B.n651 585
R776 B.n653 B.n652 585
R777 B.n650 B.n86 585
R778 B.n89 B.n86 585
R779 B.n649 B.n648 585
R780 B.n648 B.n647 585
R781 B.n88 B.n87 585
R782 B.n646 B.n88 585
R783 B.n644 B.n643 585
R784 B.n645 B.n644 585
R785 B.n642 B.n94 585
R786 B.n94 B.n93 585
R787 B.n641 B.n640 585
R788 B.n640 B.n639 585
R789 B.n96 B.n95 585
R790 B.n638 B.n96 585
R791 B.n636 B.n635 585
R792 B.n637 B.n636 585
R793 B.n745 B.n744 585
R794 B.n743 B.n2 585
R795 B.n636 B.n101 545.355
R796 B.n561 B.n99 545.355
R797 B.n329 B.n228 545.355
R798 B.n327 B.n230 545.355
R799 B.n562 B.n100 256.663
R800 B.n568 B.n100 256.663
R801 B.n570 B.n100 256.663
R802 B.n576 B.n100 256.663
R803 B.n578 B.n100 256.663
R804 B.n584 B.n100 256.663
R805 B.n586 B.n100 256.663
R806 B.n593 B.n100 256.663
R807 B.n595 B.n100 256.663
R808 B.n601 B.n100 256.663
R809 B.n111 B.n100 256.663
R810 B.n607 B.n100 256.663
R811 B.n613 B.n100 256.663
R812 B.n615 B.n100 256.663
R813 B.n621 B.n100 256.663
R814 B.n623 B.n100 256.663
R815 B.n629 B.n100 256.663
R816 B.n631 B.n100 256.663
R817 B.n322 B.n229 256.663
R818 B.n232 B.n229 256.663
R819 B.n315 B.n229 256.663
R820 B.n309 B.n229 256.663
R821 B.n307 B.n229 256.663
R822 B.n301 B.n229 256.663
R823 B.n299 B.n229 256.663
R824 B.n293 B.n229 256.663
R825 B.n291 B.n229 256.663
R826 B.n285 B.n229 256.663
R827 B.n283 B.n229 256.663
R828 B.n276 B.n229 256.663
R829 B.n274 B.n229 256.663
R830 B.n268 B.n229 256.663
R831 B.n266 B.n229 256.663
R832 B.n260 B.n229 256.663
R833 B.n258 B.n229 256.663
R834 B.n253 B.n229 256.663
R835 B.n747 B.n746 256.663
R836 B.n108 B.t12 229.852
R837 B.n116 B.t19 229.852
R838 B.n246 B.t8 229.852
R839 B.n239 B.t16 229.852
R840 B.n328 B.n229 195.9
R841 B.n637 B.n100 195.9
R842 B.n116 B.t20 184.76
R843 B.n246 B.t11 184.76
R844 B.n108 B.t14 184.76
R845 B.n239 B.t18 184.76
R846 B.n632 B.n630 163.367
R847 B.n628 B.n103 163.367
R848 B.n624 B.n622 163.367
R849 B.n620 B.n105 163.367
R850 B.n616 B.n614 163.367
R851 B.n612 B.n107 163.367
R852 B.n608 B.n606 163.367
R853 B.n603 B.n602 163.367
R854 B.n600 B.n113 163.367
R855 B.n596 B.n594 163.367
R856 B.n592 B.n115 163.367
R857 B.n587 B.n585 163.367
R858 B.n583 B.n119 163.367
R859 B.n579 B.n577 163.367
R860 B.n575 B.n121 163.367
R861 B.n571 B.n569 163.367
R862 B.n567 B.n123 163.367
R863 B.n563 B.n561 163.367
R864 B.n329 B.n226 163.367
R865 B.n333 B.n226 163.367
R866 B.n333 B.n220 163.367
R867 B.n341 B.n220 163.367
R868 B.n341 B.n218 163.367
R869 B.n345 B.n218 163.367
R870 B.n345 B.n213 163.367
R871 B.n354 B.n213 163.367
R872 B.n354 B.n211 163.367
R873 B.n358 B.n211 163.367
R874 B.n358 B.n205 163.367
R875 B.n366 B.n205 163.367
R876 B.n366 B.n203 163.367
R877 B.n370 B.n203 163.367
R878 B.n370 B.n197 163.367
R879 B.n378 B.n197 163.367
R880 B.n378 B.n195 163.367
R881 B.n382 B.n195 163.367
R882 B.n382 B.n189 163.367
R883 B.n390 B.n189 163.367
R884 B.n390 B.n187 163.367
R885 B.n394 B.n187 163.367
R886 B.n394 B.n181 163.367
R887 B.n402 B.n181 163.367
R888 B.n402 B.n179 163.367
R889 B.n406 B.n179 163.367
R890 B.n406 B.n172 163.367
R891 B.n414 B.n172 163.367
R892 B.n414 B.n170 163.367
R893 B.n418 B.n170 163.367
R894 B.n418 B.n165 163.367
R895 B.n426 B.n165 163.367
R896 B.n426 B.n163 163.367
R897 B.n430 B.n163 163.367
R898 B.n430 B.n157 163.367
R899 B.n438 B.n157 163.367
R900 B.n438 B.n155 163.367
R901 B.n442 B.n155 163.367
R902 B.n442 B.n149 163.367
R903 B.n450 B.n149 163.367
R904 B.n450 B.n147 163.367
R905 B.n454 B.n147 163.367
R906 B.n454 B.n141 163.367
R907 B.n462 B.n141 163.367
R908 B.n462 B.n139 163.367
R909 B.n466 B.n139 163.367
R910 B.n466 B.n133 163.367
R911 B.n474 B.n133 163.367
R912 B.n474 B.n131 163.367
R913 B.n479 B.n131 163.367
R914 B.n479 B.n125 163.367
R915 B.n487 B.n125 163.367
R916 B.n488 B.n487 163.367
R917 B.n488 B.n5 163.367
R918 B.n6 B.n5 163.367
R919 B.n7 B.n6 163.367
R920 B.n494 B.n7 163.367
R921 B.n495 B.n494 163.367
R922 B.n495 B.n13 163.367
R923 B.n14 B.n13 163.367
R924 B.n15 B.n14 163.367
R925 B.n500 B.n15 163.367
R926 B.n500 B.n20 163.367
R927 B.n21 B.n20 163.367
R928 B.n22 B.n21 163.367
R929 B.n505 B.n22 163.367
R930 B.n505 B.n27 163.367
R931 B.n28 B.n27 163.367
R932 B.n29 B.n28 163.367
R933 B.n510 B.n29 163.367
R934 B.n510 B.n34 163.367
R935 B.n35 B.n34 163.367
R936 B.n36 B.n35 163.367
R937 B.n515 B.n36 163.367
R938 B.n515 B.n41 163.367
R939 B.n42 B.n41 163.367
R940 B.n43 B.n42 163.367
R941 B.n520 B.n43 163.367
R942 B.n520 B.n48 163.367
R943 B.n49 B.n48 163.367
R944 B.n50 B.n49 163.367
R945 B.n525 B.n50 163.367
R946 B.n525 B.n55 163.367
R947 B.n56 B.n55 163.367
R948 B.n57 B.n56 163.367
R949 B.n530 B.n57 163.367
R950 B.n530 B.n62 163.367
R951 B.n63 B.n62 163.367
R952 B.n64 B.n63 163.367
R953 B.n535 B.n64 163.367
R954 B.n535 B.n69 163.367
R955 B.n70 B.n69 163.367
R956 B.n71 B.n70 163.367
R957 B.n540 B.n71 163.367
R958 B.n540 B.n76 163.367
R959 B.n77 B.n76 163.367
R960 B.n78 B.n77 163.367
R961 B.n545 B.n78 163.367
R962 B.n545 B.n83 163.367
R963 B.n84 B.n83 163.367
R964 B.n85 B.n84 163.367
R965 B.n550 B.n85 163.367
R966 B.n550 B.n90 163.367
R967 B.n91 B.n90 163.367
R968 B.n92 B.n91 163.367
R969 B.n555 B.n92 163.367
R970 B.n555 B.n97 163.367
R971 B.n98 B.n97 163.367
R972 B.n99 B.n98 163.367
R973 B.n323 B.n321 163.367
R974 B.n321 B.n320 163.367
R975 B.n317 B.n316 163.367
R976 B.n314 B.n234 163.367
R977 B.n310 B.n308 163.367
R978 B.n306 B.n236 163.367
R979 B.n302 B.n300 163.367
R980 B.n298 B.n238 163.367
R981 B.n294 B.n292 163.367
R982 B.n290 B.n243 163.367
R983 B.n286 B.n284 163.367
R984 B.n282 B.n245 163.367
R985 B.n277 B.n275 163.367
R986 B.n273 B.n249 163.367
R987 B.n269 B.n267 163.367
R988 B.n265 B.n251 163.367
R989 B.n261 B.n259 163.367
R990 B.n257 B.n254 163.367
R991 B.n327 B.n224 163.367
R992 B.n335 B.n224 163.367
R993 B.n335 B.n222 163.367
R994 B.n339 B.n222 163.367
R995 B.n339 B.n216 163.367
R996 B.n348 B.n216 163.367
R997 B.n348 B.n214 163.367
R998 B.n352 B.n214 163.367
R999 B.n352 B.n209 163.367
R1000 B.n360 B.n209 163.367
R1001 B.n360 B.n207 163.367
R1002 B.n364 B.n207 163.367
R1003 B.n364 B.n201 163.367
R1004 B.n372 B.n201 163.367
R1005 B.n372 B.n199 163.367
R1006 B.n376 B.n199 163.367
R1007 B.n376 B.n193 163.367
R1008 B.n384 B.n193 163.367
R1009 B.n384 B.n191 163.367
R1010 B.n388 B.n191 163.367
R1011 B.n388 B.n185 163.367
R1012 B.n396 B.n185 163.367
R1013 B.n396 B.n183 163.367
R1014 B.n400 B.n183 163.367
R1015 B.n400 B.n177 163.367
R1016 B.n408 B.n177 163.367
R1017 B.n408 B.n175 163.367
R1018 B.n412 B.n175 163.367
R1019 B.n412 B.n169 163.367
R1020 B.n420 B.n169 163.367
R1021 B.n420 B.n167 163.367
R1022 B.n424 B.n167 163.367
R1023 B.n424 B.n161 163.367
R1024 B.n432 B.n161 163.367
R1025 B.n432 B.n159 163.367
R1026 B.n436 B.n159 163.367
R1027 B.n436 B.n153 163.367
R1028 B.n444 B.n153 163.367
R1029 B.n444 B.n151 163.367
R1030 B.n448 B.n151 163.367
R1031 B.n448 B.n145 163.367
R1032 B.n456 B.n145 163.367
R1033 B.n456 B.n143 163.367
R1034 B.n460 B.n143 163.367
R1035 B.n460 B.n137 163.367
R1036 B.n468 B.n137 163.367
R1037 B.n468 B.n135 163.367
R1038 B.n472 B.n135 163.367
R1039 B.n472 B.n129 163.367
R1040 B.n481 B.n129 163.367
R1041 B.n481 B.n127 163.367
R1042 B.n485 B.n127 163.367
R1043 B.n485 B.n3 163.367
R1044 B.n745 B.n3 163.367
R1045 B.n741 B.n2 163.367
R1046 B.n741 B.n740 163.367
R1047 B.n740 B.n9 163.367
R1048 B.n736 B.n9 163.367
R1049 B.n736 B.n11 163.367
R1050 B.n732 B.n11 163.367
R1051 B.n732 B.n17 163.367
R1052 B.n728 B.n17 163.367
R1053 B.n728 B.n19 163.367
R1054 B.n724 B.n19 163.367
R1055 B.n724 B.n24 163.367
R1056 B.n720 B.n24 163.367
R1057 B.n720 B.n26 163.367
R1058 B.n716 B.n26 163.367
R1059 B.n716 B.n31 163.367
R1060 B.n712 B.n31 163.367
R1061 B.n712 B.n33 163.367
R1062 B.n708 B.n33 163.367
R1063 B.n708 B.n38 163.367
R1064 B.n704 B.n38 163.367
R1065 B.n704 B.n40 163.367
R1066 B.n700 B.n40 163.367
R1067 B.n700 B.n45 163.367
R1068 B.n696 B.n45 163.367
R1069 B.n696 B.n47 163.367
R1070 B.n692 B.n47 163.367
R1071 B.n692 B.n52 163.367
R1072 B.n688 B.n52 163.367
R1073 B.n688 B.n54 163.367
R1074 B.n684 B.n54 163.367
R1075 B.n684 B.n59 163.367
R1076 B.n680 B.n59 163.367
R1077 B.n680 B.n61 163.367
R1078 B.n676 B.n61 163.367
R1079 B.n676 B.n66 163.367
R1080 B.n672 B.n66 163.367
R1081 B.n672 B.n68 163.367
R1082 B.n668 B.n68 163.367
R1083 B.n668 B.n73 163.367
R1084 B.n664 B.n73 163.367
R1085 B.n664 B.n75 163.367
R1086 B.n660 B.n75 163.367
R1087 B.n660 B.n80 163.367
R1088 B.n656 B.n80 163.367
R1089 B.n656 B.n82 163.367
R1090 B.n652 B.n82 163.367
R1091 B.n652 B.n86 163.367
R1092 B.n648 B.n86 163.367
R1093 B.n648 B.n88 163.367
R1094 B.n644 B.n88 163.367
R1095 B.n644 B.n94 163.367
R1096 B.n640 B.n94 163.367
R1097 B.n640 B.n96 163.367
R1098 B.n636 B.n96 163.367
R1099 B.n117 B.t21 123.281
R1100 B.n247 B.t10 123.281
R1101 B.n109 B.t15 123.281
R1102 B.n240 B.t17 123.281
R1103 B.n328 B.n225 95.8365
R1104 B.n334 B.n225 95.8365
R1105 B.n334 B.n221 95.8365
R1106 B.n340 B.n221 95.8365
R1107 B.n340 B.n217 95.8365
R1108 B.n347 B.n217 95.8365
R1109 B.n347 B.n346 95.8365
R1110 B.n353 B.n210 95.8365
R1111 B.n359 B.n210 95.8365
R1112 B.n359 B.n206 95.8365
R1113 B.n365 B.n206 95.8365
R1114 B.n365 B.n202 95.8365
R1115 B.n371 B.n202 95.8365
R1116 B.n371 B.n198 95.8365
R1117 B.n377 B.n198 95.8365
R1118 B.n377 B.n194 95.8365
R1119 B.n383 B.n194 95.8365
R1120 B.n383 B.n190 95.8365
R1121 B.n389 B.n190 95.8365
R1122 B.n395 B.n186 95.8365
R1123 B.n395 B.n182 95.8365
R1124 B.n401 B.n182 95.8365
R1125 B.n401 B.n178 95.8365
R1126 B.n407 B.n178 95.8365
R1127 B.n407 B.n173 95.8365
R1128 B.n413 B.n173 95.8365
R1129 B.n413 B.n174 95.8365
R1130 B.n419 B.n166 95.8365
R1131 B.n425 B.n166 95.8365
R1132 B.n425 B.n162 95.8365
R1133 B.n431 B.n162 95.8365
R1134 B.n431 B.n158 95.8365
R1135 B.n437 B.n158 95.8365
R1136 B.n437 B.n154 95.8365
R1137 B.n443 B.n154 95.8365
R1138 B.n449 B.n150 95.8365
R1139 B.n449 B.n146 95.8365
R1140 B.n455 B.n146 95.8365
R1141 B.n455 B.n142 95.8365
R1142 B.n461 B.n142 95.8365
R1143 B.n461 B.n138 95.8365
R1144 B.n467 B.n138 95.8365
R1145 B.n467 B.n134 95.8365
R1146 B.n473 B.n134 95.8365
R1147 B.n480 B.n130 95.8365
R1148 B.n480 B.n126 95.8365
R1149 B.n486 B.n126 95.8365
R1150 B.n486 B.n4 95.8365
R1151 B.n744 B.n4 95.8365
R1152 B.n744 B.n743 95.8365
R1153 B.n743 B.n742 95.8365
R1154 B.n742 B.n8 95.8365
R1155 B.n12 B.n8 95.8365
R1156 B.n735 B.n12 95.8365
R1157 B.n735 B.n734 95.8365
R1158 B.n733 B.n16 95.8365
R1159 B.n727 B.n16 95.8365
R1160 B.n727 B.n726 95.8365
R1161 B.n726 B.n725 95.8365
R1162 B.n725 B.n23 95.8365
R1163 B.n719 B.n23 95.8365
R1164 B.n719 B.n718 95.8365
R1165 B.n718 B.n717 95.8365
R1166 B.n717 B.n30 95.8365
R1167 B.n711 B.n710 95.8365
R1168 B.n710 B.n709 95.8365
R1169 B.n709 B.n37 95.8365
R1170 B.n703 B.n37 95.8365
R1171 B.n703 B.n702 95.8365
R1172 B.n702 B.n701 95.8365
R1173 B.n701 B.n44 95.8365
R1174 B.n695 B.n44 95.8365
R1175 B.n694 B.n693 95.8365
R1176 B.n693 B.n51 95.8365
R1177 B.n687 B.n51 95.8365
R1178 B.n687 B.n686 95.8365
R1179 B.n686 B.n685 95.8365
R1180 B.n685 B.n58 95.8365
R1181 B.n679 B.n58 95.8365
R1182 B.n679 B.n678 95.8365
R1183 B.n677 B.n65 95.8365
R1184 B.n671 B.n65 95.8365
R1185 B.n671 B.n670 95.8365
R1186 B.n670 B.n669 95.8365
R1187 B.n669 B.n72 95.8365
R1188 B.n663 B.n72 95.8365
R1189 B.n663 B.n662 95.8365
R1190 B.n662 B.n661 95.8365
R1191 B.n661 B.n79 95.8365
R1192 B.n655 B.n79 95.8365
R1193 B.n655 B.n654 95.8365
R1194 B.n654 B.n653 95.8365
R1195 B.n647 B.n89 95.8365
R1196 B.n647 B.n646 95.8365
R1197 B.n646 B.n645 95.8365
R1198 B.n645 B.n93 95.8365
R1199 B.n639 B.n93 95.8365
R1200 B.n639 B.n638 95.8365
R1201 B.n638 B.n637 95.8365
R1202 B.n443 B.t4 87.3804
R1203 B.n711 B.t5 87.3804
R1204 B.t2 B.n130 73.2869
R1205 B.n734 B.t7 73.2869
R1206 B.n631 B.n101 71.676
R1207 B.n630 B.n629 71.676
R1208 B.n623 B.n103 71.676
R1209 B.n622 B.n621 71.676
R1210 B.n615 B.n105 71.676
R1211 B.n614 B.n613 71.676
R1212 B.n607 B.n107 71.676
R1213 B.n606 B.n111 71.676
R1214 B.n602 B.n601 71.676
R1215 B.n595 B.n113 71.676
R1216 B.n594 B.n593 71.676
R1217 B.n586 B.n115 71.676
R1218 B.n585 B.n584 71.676
R1219 B.n578 B.n119 71.676
R1220 B.n577 B.n576 71.676
R1221 B.n570 B.n121 71.676
R1222 B.n569 B.n568 71.676
R1223 B.n562 B.n123 71.676
R1224 B.n563 B.n562 71.676
R1225 B.n568 B.n567 71.676
R1226 B.n571 B.n570 71.676
R1227 B.n576 B.n575 71.676
R1228 B.n579 B.n578 71.676
R1229 B.n584 B.n583 71.676
R1230 B.n587 B.n586 71.676
R1231 B.n593 B.n592 71.676
R1232 B.n596 B.n595 71.676
R1233 B.n601 B.n600 71.676
R1234 B.n603 B.n111 71.676
R1235 B.n608 B.n607 71.676
R1236 B.n613 B.n612 71.676
R1237 B.n616 B.n615 71.676
R1238 B.n621 B.n620 71.676
R1239 B.n624 B.n623 71.676
R1240 B.n629 B.n628 71.676
R1241 B.n632 B.n631 71.676
R1242 B.n322 B.n230 71.676
R1243 B.n320 B.n232 71.676
R1244 B.n316 B.n315 71.676
R1245 B.n309 B.n234 71.676
R1246 B.n308 B.n307 71.676
R1247 B.n301 B.n236 71.676
R1248 B.n300 B.n299 71.676
R1249 B.n293 B.n238 71.676
R1250 B.n292 B.n291 71.676
R1251 B.n285 B.n243 71.676
R1252 B.n284 B.n283 71.676
R1253 B.n276 B.n245 71.676
R1254 B.n275 B.n274 71.676
R1255 B.n268 B.n249 71.676
R1256 B.n267 B.n266 71.676
R1257 B.n260 B.n251 71.676
R1258 B.n259 B.n258 71.676
R1259 B.n254 B.n253 71.676
R1260 B.n323 B.n322 71.676
R1261 B.n317 B.n232 71.676
R1262 B.n315 B.n314 71.676
R1263 B.n310 B.n309 71.676
R1264 B.n307 B.n306 71.676
R1265 B.n302 B.n301 71.676
R1266 B.n299 B.n298 71.676
R1267 B.n294 B.n293 71.676
R1268 B.n291 B.n290 71.676
R1269 B.n286 B.n285 71.676
R1270 B.n283 B.n282 71.676
R1271 B.n277 B.n276 71.676
R1272 B.n274 B.n273 71.676
R1273 B.n269 B.n268 71.676
R1274 B.n266 B.n265 71.676
R1275 B.n261 B.n260 71.676
R1276 B.n258 B.n257 71.676
R1277 B.n253 B.n228 71.676
R1278 B.n746 B.n745 71.676
R1279 B.n746 B.n2 71.676
R1280 B.n346 B.t9 70.4682
R1281 B.t1 B.n186 70.4682
R1282 B.n678 B.t0 70.4682
R1283 B.n89 B.t13 70.4682
R1284 B.n109 B.n108 61.4793
R1285 B.n117 B.n116 61.4793
R1286 B.n247 B.n246 61.4793
R1287 B.n240 B.n239 61.4793
R1288 B.n110 B.n109 59.5399
R1289 B.n589 B.n117 59.5399
R1290 B.n280 B.n247 59.5399
R1291 B.n241 B.n240 59.5399
R1292 B.n174 B.t6 56.3746
R1293 B.t3 B.n694 56.3746
R1294 B.n419 B.t6 39.4624
R1295 B.n695 B.t3 39.4624
R1296 B.n560 B.n559 35.4346
R1297 B.n326 B.n325 35.4346
R1298 B.n330 B.n227 35.4346
R1299 B.n635 B.n634 35.4346
R1300 B.n353 B.t9 25.3689
R1301 B.n389 B.t1 25.3689
R1302 B.t0 B.n677 25.3689
R1303 B.n653 B.t13 25.3689
R1304 B.n473 B.t2 22.5501
R1305 B.t7 B.n733 22.5501
R1306 B B.n747 18.0485
R1307 B.n326 B.n223 10.6151
R1308 B.n336 B.n223 10.6151
R1309 B.n337 B.n336 10.6151
R1310 B.n338 B.n337 10.6151
R1311 B.n338 B.n215 10.6151
R1312 B.n349 B.n215 10.6151
R1313 B.n350 B.n349 10.6151
R1314 B.n351 B.n350 10.6151
R1315 B.n351 B.n208 10.6151
R1316 B.n361 B.n208 10.6151
R1317 B.n362 B.n361 10.6151
R1318 B.n363 B.n362 10.6151
R1319 B.n363 B.n200 10.6151
R1320 B.n373 B.n200 10.6151
R1321 B.n374 B.n373 10.6151
R1322 B.n375 B.n374 10.6151
R1323 B.n375 B.n192 10.6151
R1324 B.n385 B.n192 10.6151
R1325 B.n386 B.n385 10.6151
R1326 B.n387 B.n386 10.6151
R1327 B.n387 B.n184 10.6151
R1328 B.n397 B.n184 10.6151
R1329 B.n398 B.n397 10.6151
R1330 B.n399 B.n398 10.6151
R1331 B.n399 B.n176 10.6151
R1332 B.n409 B.n176 10.6151
R1333 B.n410 B.n409 10.6151
R1334 B.n411 B.n410 10.6151
R1335 B.n411 B.n168 10.6151
R1336 B.n421 B.n168 10.6151
R1337 B.n422 B.n421 10.6151
R1338 B.n423 B.n422 10.6151
R1339 B.n423 B.n160 10.6151
R1340 B.n433 B.n160 10.6151
R1341 B.n434 B.n433 10.6151
R1342 B.n435 B.n434 10.6151
R1343 B.n435 B.n152 10.6151
R1344 B.n445 B.n152 10.6151
R1345 B.n446 B.n445 10.6151
R1346 B.n447 B.n446 10.6151
R1347 B.n447 B.n144 10.6151
R1348 B.n457 B.n144 10.6151
R1349 B.n458 B.n457 10.6151
R1350 B.n459 B.n458 10.6151
R1351 B.n459 B.n136 10.6151
R1352 B.n469 B.n136 10.6151
R1353 B.n470 B.n469 10.6151
R1354 B.n471 B.n470 10.6151
R1355 B.n471 B.n128 10.6151
R1356 B.n482 B.n128 10.6151
R1357 B.n483 B.n482 10.6151
R1358 B.n484 B.n483 10.6151
R1359 B.n484 B.n0 10.6151
R1360 B.n325 B.n324 10.6151
R1361 B.n324 B.n231 10.6151
R1362 B.n319 B.n231 10.6151
R1363 B.n319 B.n318 10.6151
R1364 B.n318 B.n233 10.6151
R1365 B.n313 B.n233 10.6151
R1366 B.n313 B.n312 10.6151
R1367 B.n312 B.n311 10.6151
R1368 B.n311 B.n235 10.6151
R1369 B.n305 B.n235 10.6151
R1370 B.n305 B.n304 10.6151
R1371 B.n304 B.n303 10.6151
R1372 B.n303 B.n237 10.6151
R1373 B.n297 B.n296 10.6151
R1374 B.n296 B.n295 10.6151
R1375 B.n295 B.n242 10.6151
R1376 B.n289 B.n242 10.6151
R1377 B.n289 B.n288 10.6151
R1378 B.n288 B.n287 10.6151
R1379 B.n287 B.n244 10.6151
R1380 B.n281 B.n244 10.6151
R1381 B.n279 B.n278 10.6151
R1382 B.n278 B.n248 10.6151
R1383 B.n272 B.n248 10.6151
R1384 B.n272 B.n271 10.6151
R1385 B.n271 B.n270 10.6151
R1386 B.n270 B.n250 10.6151
R1387 B.n264 B.n250 10.6151
R1388 B.n264 B.n263 10.6151
R1389 B.n263 B.n262 10.6151
R1390 B.n262 B.n252 10.6151
R1391 B.n256 B.n252 10.6151
R1392 B.n256 B.n255 10.6151
R1393 B.n255 B.n227 10.6151
R1394 B.n331 B.n330 10.6151
R1395 B.n332 B.n331 10.6151
R1396 B.n332 B.n219 10.6151
R1397 B.n342 B.n219 10.6151
R1398 B.n343 B.n342 10.6151
R1399 B.n344 B.n343 10.6151
R1400 B.n344 B.n212 10.6151
R1401 B.n355 B.n212 10.6151
R1402 B.n356 B.n355 10.6151
R1403 B.n357 B.n356 10.6151
R1404 B.n357 B.n204 10.6151
R1405 B.n367 B.n204 10.6151
R1406 B.n368 B.n367 10.6151
R1407 B.n369 B.n368 10.6151
R1408 B.n369 B.n196 10.6151
R1409 B.n379 B.n196 10.6151
R1410 B.n380 B.n379 10.6151
R1411 B.n381 B.n380 10.6151
R1412 B.n381 B.n188 10.6151
R1413 B.n391 B.n188 10.6151
R1414 B.n392 B.n391 10.6151
R1415 B.n393 B.n392 10.6151
R1416 B.n393 B.n180 10.6151
R1417 B.n403 B.n180 10.6151
R1418 B.n404 B.n403 10.6151
R1419 B.n405 B.n404 10.6151
R1420 B.n405 B.n171 10.6151
R1421 B.n415 B.n171 10.6151
R1422 B.n416 B.n415 10.6151
R1423 B.n417 B.n416 10.6151
R1424 B.n417 B.n164 10.6151
R1425 B.n427 B.n164 10.6151
R1426 B.n428 B.n427 10.6151
R1427 B.n429 B.n428 10.6151
R1428 B.n429 B.n156 10.6151
R1429 B.n439 B.n156 10.6151
R1430 B.n440 B.n439 10.6151
R1431 B.n441 B.n440 10.6151
R1432 B.n441 B.n148 10.6151
R1433 B.n451 B.n148 10.6151
R1434 B.n452 B.n451 10.6151
R1435 B.n453 B.n452 10.6151
R1436 B.n453 B.n140 10.6151
R1437 B.n463 B.n140 10.6151
R1438 B.n464 B.n463 10.6151
R1439 B.n465 B.n464 10.6151
R1440 B.n465 B.n132 10.6151
R1441 B.n475 B.n132 10.6151
R1442 B.n476 B.n475 10.6151
R1443 B.n478 B.n476 10.6151
R1444 B.n478 B.n477 10.6151
R1445 B.n477 B.n124 10.6151
R1446 B.n489 B.n124 10.6151
R1447 B.n490 B.n489 10.6151
R1448 B.n491 B.n490 10.6151
R1449 B.n492 B.n491 10.6151
R1450 B.n493 B.n492 10.6151
R1451 B.n496 B.n493 10.6151
R1452 B.n497 B.n496 10.6151
R1453 B.n498 B.n497 10.6151
R1454 B.n499 B.n498 10.6151
R1455 B.n501 B.n499 10.6151
R1456 B.n502 B.n501 10.6151
R1457 B.n503 B.n502 10.6151
R1458 B.n504 B.n503 10.6151
R1459 B.n506 B.n504 10.6151
R1460 B.n507 B.n506 10.6151
R1461 B.n508 B.n507 10.6151
R1462 B.n509 B.n508 10.6151
R1463 B.n511 B.n509 10.6151
R1464 B.n512 B.n511 10.6151
R1465 B.n513 B.n512 10.6151
R1466 B.n514 B.n513 10.6151
R1467 B.n516 B.n514 10.6151
R1468 B.n517 B.n516 10.6151
R1469 B.n518 B.n517 10.6151
R1470 B.n519 B.n518 10.6151
R1471 B.n521 B.n519 10.6151
R1472 B.n522 B.n521 10.6151
R1473 B.n523 B.n522 10.6151
R1474 B.n524 B.n523 10.6151
R1475 B.n526 B.n524 10.6151
R1476 B.n527 B.n526 10.6151
R1477 B.n528 B.n527 10.6151
R1478 B.n529 B.n528 10.6151
R1479 B.n531 B.n529 10.6151
R1480 B.n532 B.n531 10.6151
R1481 B.n533 B.n532 10.6151
R1482 B.n534 B.n533 10.6151
R1483 B.n536 B.n534 10.6151
R1484 B.n537 B.n536 10.6151
R1485 B.n538 B.n537 10.6151
R1486 B.n539 B.n538 10.6151
R1487 B.n541 B.n539 10.6151
R1488 B.n542 B.n541 10.6151
R1489 B.n543 B.n542 10.6151
R1490 B.n544 B.n543 10.6151
R1491 B.n546 B.n544 10.6151
R1492 B.n547 B.n546 10.6151
R1493 B.n548 B.n547 10.6151
R1494 B.n549 B.n548 10.6151
R1495 B.n551 B.n549 10.6151
R1496 B.n552 B.n551 10.6151
R1497 B.n553 B.n552 10.6151
R1498 B.n554 B.n553 10.6151
R1499 B.n556 B.n554 10.6151
R1500 B.n557 B.n556 10.6151
R1501 B.n558 B.n557 10.6151
R1502 B.n559 B.n558 10.6151
R1503 B.n739 B.n1 10.6151
R1504 B.n739 B.n738 10.6151
R1505 B.n738 B.n737 10.6151
R1506 B.n737 B.n10 10.6151
R1507 B.n731 B.n10 10.6151
R1508 B.n731 B.n730 10.6151
R1509 B.n730 B.n729 10.6151
R1510 B.n729 B.n18 10.6151
R1511 B.n723 B.n18 10.6151
R1512 B.n723 B.n722 10.6151
R1513 B.n722 B.n721 10.6151
R1514 B.n721 B.n25 10.6151
R1515 B.n715 B.n25 10.6151
R1516 B.n715 B.n714 10.6151
R1517 B.n714 B.n713 10.6151
R1518 B.n713 B.n32 10.6151
R1519 B.n707 B.n32 10.6151
R1520 B.n707 B.n706 10.6151
R1521 B.n706 B.n705 10.6151
R1522 B.n705 B.n39 10.6151
R1523 B.n699 B.n39 10.6151
R1524 B.n699 B.n698 10.6151
R1525 B.n698 B.n697 10.6151
R1526 B.n697 B.n46 10.6151
R1527 B.n691 B.n46 10.6151
R1528 B.n691 B.n690 10.6151
R1529 B.n690 B.n689 10.6151
R1530 B.n689 B.n53 10.6151
R1531 B.n683 B.n53 10.6151
R1532 B.n683 B.n682 10.6151
R1533 B.n682 B.n681 10.6151
R1534 B.n681 B.n60 10.6151
R1535 B.n675 B.n60 10.6151
R1536 B.n675 B.n674 10.6151
R1537 B.n674 B.n673 10.6151
R1538 B.n673 B.n67 10.6151
R1539 B.n667 B.n67 10.6151
R1540 B.n667 B.n666 10.6151
R1541 B.n666 B.n665 10.6151
R1542 B.n665 B.n74 10.6151
R1543 B.n659 B.n74 10.6151
R1544 B.n659 B.n658 10.6151
R1545 B.n658 B.n657 10.6151
R1546 B.n657 B.n81 10.6151
R1547 B.n651 B.n81 10.6151
R1548 B.n651 B.n650 10.6151
R1549 B.n650 B.n649 10.6151
R1550 B.n649 B.n87 10.6151
R1551 B.n643 B.n87 10.6151
R1552 B.n643 B.n642 10.6151
R1553 B.n642 B.n641 10.6151
R1554 B.n641 B.n95 10.6151
R1555 B.n635 B.n95 10.6151
R1556 B.n634 B.n633 10.6151
R1557 B.n633 B.n102 10.6151
R1558 B.n627 B.n102 10.6151
R1559 B.n627 B.n626 10.6151
R1560 B.n626 B.n625 10.6151
R1561 B.n625 B.n104 10.6151
R1562 B.n619 B.n104 10.6151
R1563 B.n619 B.n618 10.6151
R1564 B.n618 B.n617 10.6151
R1565 B.n617 B.n106 10.6151
R1566 B.n611 B.n106 10.6151
R1567 B.n611 B.n610 10.6151
R1568 B.n610 B.n609 10.6151
R1569 B.n605 B.n604 10.6151
R1570 B.n604 B.n112 10.6151
R1571 B.n599 B.n112 10.6151
R1572 B.n599 B.n598 10.6151
R1573 B.n598 B.n597 10.6151
R1574 B.n597 B.n114 10.6151
R1575 B.n591 B.n114 10.6151
R1576 B.n591 B.n590 10.6151
R1577 B.n588 B.n118 10.6151
R1578 B.n582 B.n118 10.6151
R1579 B.n582 B.n581 10.6151
R1580 B.n581 B.n580 10.6151
R1581 B.n580 B.n120 10.6151
R1582 B.n574 B.n120 10.6151
R1583 B.n574 B.n573 10.6151
R1584 B.n573 B.n572 10.6151
R1585 B.n572 B.n122 10.6151
R1586 B.n566 B.n122 10.6151
R1587 B.n566 B.n565 10.6151
R1588 B.n565 B.n564 10.6151
R1589 B.n564 B.n560 10.6151
R1590 B.t4 B.n150 8.45662
R1591 B.t5 B.n30 8.45662
R1592 B.n747 B.n0 8.11757
R1593 B.n747 B.n1 8.11757
R1594 B.n297 B.n241 6.5566
R1595 B.n281 B.n280 6.5566
R1596 B.n605 B.n110 6.5566
R1597 B.n590 B.n589 6.5566
R1598 B.n241 B.n237 4.05904
R1599 B.n280 B.n279 4.05904
R1600 B.n609 B.n110 4.05904
R1601 B.n589 B.n588 4.05904
R1602 VP.n19 VP.n16 161.3
R1603 VP.n21 VP.n20 161.3
R1604 VP.n22 VP.n15 161.3
R1605 VP.n24 VP.n23 161.3
R1606 VP.n25 VP.n14 161.3
R1607 VP.n28 VP.n27 161.3
R1608 VP.n29 VP.n13 161.3
R1609 VP.n31 VP.n30 161.3
R1610 VP.n32 VP.n12 161.3
R1611 VP.n34 VP.n33 161.3
R1612 VP.n35 VP.n11 161.3
R1613 VP.n37 VP.n36 161.3
R1614 VP.n38 VP.n10 161.3
R1615 VP.n74 VP.n0 161.3
R1616 VP.n73 VP.n72 161.3
R1617 VP.n71 VP.n1 161.3
R1618 VP.n70 VP.n69 161.3
R1619 VP.n68 VP.n2 161.3
R1620 VP.n67 VP.n66 161.3
R1621 VP.n65 VP.n3 161.3
R1622 VP.n64 VP.n63 161.3
R1623 VP.n61 VP.n4 161.3
R1624 VP.n60 VP.n59 161.3
R1625 VP.n58 VP.n5 161.3
R1626 VP.n57 VP.n56 161.3
R1627 VP.n55 VP.n6 161.3
R1628 VP.n53 VP.n52 161.3
R1629 VP.n51 VP.n7 161.3
R1630 VP.n50 VP.n49 161.3
R1631 VP.n48 VP.n8 161.3
R1632 VP.n47 VP.n46 161.3
R1633 VP.n45 VP.n9 161.3
R1634 VP.n44 VP.n43 161.3
R1635 VP.n42 VP.n41 110.511
R1636 VP.n76 VP.n75 110.511
R1637 VP.n40 VP.n39 110.511
R1638 VP.n18 VP.n17 57.3183
R1639 VP.n60 VP.n5 56.5193
R1640 VP.n24 VP.n15 56.5193
R1641 VP.n17 VP.t0 53.5387
R1642 VP.n49 VP.n48 48.2635
R1643 VP.n69 VP.n68 48.2635
R1644 VP.n33 VP.n32 48.2635
R1645 VP.n41 VP.n40 44.7723
R1646 VP.n48 VP.n47 32.7233
R1647 VP.n69 VP.n1 32.7233
R1648 VP.n33 VP.n11 32.7233
R1649 VP.n43 VP.n9 24.4675
R1650 VP.n47 VP.n9 24.4675
R1651 VP.n49 VP.n7 24.4675
R1652 VP.n53 VP.n7 24.4675
R1653 VP.n56 VP.n55 24.4675
R1654 VP.n56 VP.n5 24.4675
R1655 VP.n61 VP.n60 24.4675
R1656 VP.n63 VP.n61 24.4675
R1657 VP.n67 VP.n3 24.4675
R1658 VP.n68 VP.n67 24.4675
R1659 VP.n73 VP.n1 24.4675
R1660 VP.n74 VP.n73 24.4675
R1661 VP.n37 VP.n11 24.4675
R1662 VP.n38 VP.n37 24.4675
R1663 VP.n25 VP.n24 24.4675
R1664 VP.n27 VP.n25 24.4675
R1665 VP.n31 VP.n13 24.4675
R1666 VP.n32 VP.n31 24.4675
R1667 VP.n20 VP.n19 24.4675
R1668 VP.n20 VP.n15 24.4675
R1669 VP.n42 VP.t6 21.4699
R1670 VP.n54 VP.t7 21.4699
R1671 VP.n62 VP.t2 21.4699
R1672 VP.n75 VP.t5 21.4699
R1673 VP.n39 VP.t4 21.4699
R1674 VP.n26 VP.t3 21.4699
R1675 VP.n18 VP.t1 21.4699
R1676 VP.n55 VP.n54 16.3934
R1677 VP.n63 VP.n62 16.3934
R1678 VP.n27 VP.n26 16.3934
R1679 VP.n19 VP.n18 16.3934
R1680 VP.n54 VP.n53 8.07461
R1681 VP.n62 VP.n3 8.07461
R1682 VP.n26 VP.n13 8.07461
R1683 VP.n17 VP.n16 5.19262
R1684 VP.n40 VP.n10 0.278367
R1685 VP.n44 VP.n41 0.278367
R1686 VP.n76 VP.n0 0.278367
R1687 VP.n43 VP.n42 0.24517
R1688 VP.n75 VP.n74 0.24517
R1689 VP.n39 VP.n38 0.24517
R1690 VP.n21 VP.n16 0.189894
R1691 VP.n22 VP.n21 0.189894
R1692 VP.n23 VP.n22 0.189894
R1693 VP.n23 VP.n14 0.189894
R1694 VP.n28 VP.n14 0.189894
R1695 VP.n29 VP.n28 0.189894
R1696 VP.n30 VP.n29 0.189894
R1697 VP.n30 VP.n12 0.189894
R1698 VP.n34 VP.n12 0.189894
R1699 VP.n35 VP.n34 0.189894
R1700 VP.n36 VP.n35 0.189894
R1701 VP.n36 VP.n10 0.189894
R1702 VP.n45 VP.n44 0.189894
R1703 VP.n46 VP.n45 0.189894
R1704 VP.n46 VP.n8 0.189894
R1705 VP.n50 VP.n8 0.189894
R1706 VP.n51 VP.n50 0.189894
R1707 VP.n52 VP.n51 0.189894
R1708 VP.n52 VP.n6 0.189894
R1709 VP.n57 VP.n6 0.189894
R1710 VP.n58 VP.n57 0.189894
R1711 VP.n59 VP.n58 0.189894
R1712 VP.n59 VP.n4 0.189894
R1713 VP.n64 VP.n4 0.189894
R1714 VP.n65 VP.n64 0.189894
R1715 VP.n66 VP.n65 0.189894
R1716 VP.n66 VP.n2 0.189894
R1717 VP.n70 VP.n2 0.189894
R1718 VP.n71 VP.n70 0.189894
R1719 VP.n72 VP.n71 0.189894
R1720 VP.n72 VP.n0 0.189894
R1721 VP VP.n76 0.153454
R1722 VDD1 VDD1.n0 88.9051
R1723 VDD1.n3 VDD1.n2 88.7914
R1724 VDD1.n3 VDD1.n1 88.7914
R1725 VDD1.n5 VDD1.n4 87.4804
R1726 VDD1.n5 VDD1.n3 38.7768
R1727 VDD1.n4 VDD1.t4 7.82659
R1728 VDD1.n4 VDD1.t3 7.82659
R1729 VDD1.n0 VDD1.t7 7.82659
R1730 VDD1.n0 VDD1.t6 7.82659
R1731 VDD1.n2 VDD1.t5 7.82659
R1732 VDD1.n2 VDD1.t2 7.82659
R1733 VDD1.n1 VDD1.t1 7.82659
R1734 VDD1.n1 VDD1.t0 7.82659
R1735 VDD1 VDD1.n5 1.30869
C0 VN VP 6.21097f
C1 VTAIL VP 3.4171f
C2 VTAIL VN 3.40299f
C3 VDD1 VP 2.6227f
C4 VDD2 VP 0.551336f
C5 VDD1 VN 0.157281f
C6 VDD2 VN 2.23143f
C7 VDD1 VTAIL 5.098721f
C8 VDD2 VTAIL 5.15475f
C9 VDD2 VDD1 1.90095f
C10 VDD2 B 4.808663f
C11 VDD1 B 5.28228f
C12 VTAIL B 4.516549f
C13 VN B 15.616529f
C14 VP B 14.128262f
C15 VDD1.t7 B 0.049694f
C16 VDD1.t6 B 0.049694f
C17 VDD1.n0 B 0.361366f
C18 VDD1.t1 B 0.049694f
C19 VDD1.t0 B 0.049694f
C20 VDD1.n1 B 0.360575f
C21 VDD1.t5 B 0.049694f
C22 VDD1.t2 B 0.049694f
C23 VDD1.n2 B 0.360575f
C24 VDD1.n3 B 2.83672f
C25 VDD1.t4 B 0.049694f
C26 VDD1.t3 B 0.049694f
C27 VDD1.n4 B 0.352934f
C28 VDD1.n5 B 2.2937f
C29 VP.n0 B 0.038392f
C30 VP.t5 B 0.509116f
C31 VP.n1 B 0.058732f
C32 VP.n2 B 0.02912f
C33 VP.n3 B 0.036319f
C34 VP.n4 B 0.02912f
C35 VP.n5 B 0.04251f
C36 VP.n6 B 0.02912f
C37 VP.t7 B 0.509116f
C38 VP.n7 B 0.054273f
C39 VP.n8 B 0.02912f
C40 VP.n9 B 0.054273f
C41 VP.n10 B 0.038392f
C42 VP.t4 B 0.509116f
C43 VP.n11 B 0.058732f
C44 VP.n12 B 0.02912f
C45 VP.n13 B 0.036319f
C46 VP.n14 B 0.02912f
C47 VP.n15 B 0.04251f
C48 VP.n16 B 0.30689f
C49 VP.t1 B 0.509116f
C50 VP.t0 B 0.759037f
C51 VP.n17 B 0.307196f
C52 VP.n18 B 0.31691f
C53 VP.n19 B 0.045429f
C54 VP.n20 B 0.054273f
C55 VP.n21 B 0.02912f
C56 VP.n22 B 0.02912f
C57 VP.n23 B 0.02912f
C58 VP.n24 B 0.04251f
C59 VP.n25 B 0.054273f
C60 VP.t3 B 0.509116f
C61 VP.n26 B 0.222249f
C62 VP.n27 B 0.045429f
C63 VP.n28 B 0.02912f
C64 VP.n29 B 0.02912f
C65 VP.n30 B 0.02912f
C66 VP.n31 B 0.054273f
C67 VP.n32 B 0.054534f
C68 VP.n33 B 0.026026f
C69 VP.n34 B 0.02912f
C70 VP.n35 B 0.02912f
C71 VP.n36 B 0.02912f
C72 VP.n37 B 0.054273f
C73 VP.n38 B 0.027744f
C74 VP.n39 B 0.313928f
C75 VP.n40 B 1.37971f
C76 VP.n41 B 1.40309f
C77 VP.t6 B 0.509116f
C78 VP.n42 B 0.313928f
C79 VP.n43 B 0.027744f
C80 VP.n44 B 0.038392f
C81 VP.n45 B 0.02912f
C82 VP.n46 B 0.02912f
C83 VP.n47 B 0.058732f
C84 VP.n48 B 0.026026f
C85 VP.n49 B 0.054534f
C86 VP.n50 B 0.02912f
C87 VP.n51 B 0.02912f
C88 VP.n52 B 0.02912f
C89 VP.n53 B 0.036319f
C90 VP.n54 B 0.222249f
C91 VP.n55 B 0.045429f
C92 VP.n56 B 0.054273f
C93 VP.n57 B 0.02912f
C94 VP.n58 B 0.02912f
C95 VP.n59 B 0.02912f
C96 VP.n60 B 0.04251f
C97 VP.n61 B 0.054273f
C98 VP.t2 B 0.509116f
C99 VP.n62 B 0.222249f
C100 VP.n63 B 0.045429f
C101 VP.n64 B 0.02912f
C102 VP.n65 B 0.02912f
C103 VP.n66 B 0.02912f
C104 VP.n67 B 0.054273f
C105 VP.n68 B 0.054534f
C106 VP.n69 B 0.026026f
C107 VP.n70 B 0.02912f
C108 VP.n71 B 0.02912f
C109 VP.n72 B 0.02912f
C110 VP.n73 B 0.054273f
C111 VP.n74 B 0.027744f
C112 VP.n75 B 0.313928f
C113 VP.n76 B 0.056344f
C114 VDD2.t2 B 0.048334f
C115 VDD2.t3 B 0.048334f
C116 VDD2.n0 B 0.350708f
C117 VDD2.t6 B 0.048334f
C118 VDD2.t7 B 0.048334f
C119 VDD2.n1 B 0.350708f
C120 VDD2.n2 B 2.70866f
C121 VDD2.t5 B 0.048334f
C122 VDD2.t4 B 0.048334f
C123 VDD2.n3 B 0.343277f
C124 VDD2.n4 B 2.20113f
C125 VDD2.t0 B 0.048334f
C126 VDD2.t1 B 0.048334f
C127 VDD2.n5 B 0.350682f
C128 VTAIL.t15 B 0.060324f
C129 VTAIL.t10 B 0.060324f
C130 VTAIL.n0 B 0.377404f
C131 VTAIL.n1 B 0.503701f
C132 VTAIL.n2 B 0.040986f
C133 VTAIL.n3 B 0.229948f
C134 VTAIL.n4 B 0.016214f
C135 VTAIL.t12 B 0.066601f
C136 VTAIL.n5 B 0.107458f
C137 VTAIL.n6 B 0.021694f
C138 VTAIL.n7 B 0.028742f
C139 VTAIL.n8 B 0.080443f
C140 VTAIL.n9 B 0.017167f
C141 VTAIL.n10 B 0.016214f
C142 VTAIL.n11 B 0.075102f
C143 VTAIL.n12 B 0.044911f
C144 VTAIL.n13 B 0.340167f
C145 VTAIL.n14 B 0.040986f
C146 VTAIL.n15 B 0.229948f
C147 VTAIL.n16 B 0.016214f
C148 VTAIL.t2 B 0.066601f
C149 VTAIL.n17 B 0.107458f
C150 VTAIL.n18 B 0.021694f
C151 VTAIL.n19 B 0.028742f
C152 VTAIL.n20 B 0.080443f
C153 VTAIL.n21 B 0.017167f
C154 VTAIL.n22 B 0.016214f
C155 VTAIL.n23 B 0.075102f
C156 VTAIL.n24 B 0.044911f
C157 VTAIL.n25 B 0.340167f
C158 VTAIL.t6 B 0.060324f
C159 VTAIL.t4 B 0.060324f
C160 VTAIL.n26 B 0.377404f
C161 VTAIL.n27 B 0.763733f
C162 VTAIL.n28 B 0.040986f
C163 VTAIL.n29 B 0.229948f
C164 VTAIL.n30 B 0.016214f
C165 VTAIL.t1 B 0.066601f
C166 VTAIL.n31 B 0.107458f
C167 VTAIL.n32 B 0.021694f
C168 VTAIL.n33 B 0.028742f
C169 VTAIL.n34 B 0.080443f
C170 VTAIL.n35 B 0.017167f
C171 VTAIL.n36 B 0.016214f
C172 VTAIL.n37 B 0.075102f
C173 VTAIL.n38 B 0.044911f
C174 VTAIL.n39 B 1.18209f
C175 VTAIL.n40 B 0.040986f
C176 VTAIL.n41 B 0.229948f
C177 VTAIL.n42 B 0.016214f
C178 VTAIL.t9 B 0.066601f
C179 VTAIL.n43 B 0.107458f
C180 VTAIL.n44 B 0.021694f
C181 VTAIL.n45 B 0.028742f
C182 VTAIL.n46 B 0.080443f
C183 VTAIL.n47 B 0.017167f
C184 VTAIL.n48 B 0.016214f
C185 VTAIL.n49 B 0.075102f
C186 VTAIL.n50 B 0.044911f
C187 VTAIL.n51 B 1.18209f
C188 VTAIL.t14 B 0.060324f
C189 VTAIL.t13 B 0.060324f
C190 VTAIL.n52 B 0.377406f
C191 VTAIL.n53 B 0.76373f
C192 VTAIL.n54 B 0.040986f
C193 VTAIL.n55 B 0.229948f
C194 VTAIL.n56 B 0.016214f
C195 VTAIL.t11 B 0.066601f
C196 VTAIL.n57 B 0.107458f
C197 VTAIL.n58 B 0.021694f
C198 VTAIL.n59 B 0.028742f
C199 VTAIL.n60 B 0.080443f
C200 VTAIL.n61 B 0.017167f
C201 VTAIL.n62 B 0.016214f
C202 VTAIL.n63 B 0.075102f
C203 VTAIL.n64 B 0.044911f
C204 VTAIL.n65 B 0.340167f
C205 VTAIL.n66 B 0.040986f
C206 VTAIL.n67 B 0.229948f
C207 VTAIL.n68 B 0.016214f
C208 VTAIL.t7 B 0.066601f
C209 VTAIL.n69 B 0.107458f
C210 VTAIL.n70 B 0.021694f
C211 VTAIL.n71 B 0.028742f
C212 VTAIL.n72 B 0.080443f
C213 VTAIL.n73 B 0.017167f
C214 VTAIL.n74 B 0.016214f
C215 VTAIL.n75 B 0.075102f
C216 VTAIL.n76 B 0.044911f
C217 VTAIL.n77 B 0.340167f
C218 VTAIL.t5 B 0.060324f
C219 VTAIL.t3 B 0.060324f
C220 VTAIL.n78 B 0.377406f
C221 VTAIL.n79 B 0.76373f
C222 VTAIL.n80 B 0.040986f
C223 VTAIL.n81 B 0.229948f
C224 VTAIL.n82 B 0.016214f
C225 VTAIL.t0 B 0.066601f
C226 VTAIL.n83 B 0.107458f
C227 VTAIL.n84 B 0.021694f
C228 VTAIL.n85 B 0.028742f
C229 VTAIL.n86 B 0.080443f
C230 VTAIL.n87 B 0.017167f
C231 VTAIL.n88 B 0.016214f
C232 VTAIL.n89 B 0.075102f
C233 VTAIL.n90 B 0.044911f
C234 VTAIL.n91 B 1.18209f
C235 VTAIL.n92 B 0.040986f
C236 VTAIL.n93 B 0.229948f
C237 VTAIL.n94 B 0.016214f
C238 VTAIL.t8 B 0.066601f
C239 VTAIL.n95 B 0.107458f
C240 VTAIL.n96 B 0.021694f
C241 VTAIL.n97 B 0.028742f
C242 VTAIL.n98 B 0.080443f
C243 VTAIL.n99 B 0.017167f
C244 VTAIL.n100 B 0.016214f
C245 VTAIL.n101 B 0.075102f
C246 VTAIL.n102 B 0.044911f
C247 VTAIL.n103 B 1.17643f
C248 VN.n0 B 0.037009f
C249 VN.t0 B 0.490777f
C250 VN.n1 B 0.056617f
C251 VN.n2 B 0.028071f
C252 VN.n3 B 0.035011f
C253 VN.n4 B 0.028071f
C254 VN.n5 B 0.040979f
C255 VN.n6 B 0.295835f
C256 VN.t4 B 0.490777f
C257 VN.t5 B 0.731696f
C258 VN.n7 B 0.29613f
C259 VN.n8 B 0.305495f
C260 VN.n9 B 0.043793f
C261 VN.n10 B 0.052318f
C262 VN.n11 B 0.028071f
C263 VN.n12 B 0.028071f
C264 VN.n13 B 0.028071f
C265 VN.n14 B 0.040979f
C266 VN.n15 B 0.052318f
C267 VN.t1 B 0.490777f
C268 VN.n16 B 0.214244f
C269 VN.n17 B 0.043793f
C270 VN.n18 B 0.028071f
C271 VN.n19 B 0.028071f
C272 VN.n20 B 0.028071f
C273 VN.n21 B 0.052318f
C274 VN.n22 B 0.05257f
C275 VN.n23 B 0.025088f
C276 VN.n24 B 0.028071f
C277 VN.n25 B 0.028071f
C278 VN.n26 B 0.028071f
C279 VN.n27 B 0.052318f
C280 VN.n28 B 0.026745f
C281 VN.n29 B 0.30262f
C282 VN.n30 B 0.054314f
C283 VN.n31 B 0.037009f
C284 VN.t2 B 0.490777f
C285 VN.n32 B 0.056617f
C286 VN.n33 B 0.028071f
C287 VN.n34 B 0.035011f
C288 VN.n35 B 0.028071f
C289 VN.t3 B 0.490777f
C290 VN.n36 B 0.214244f
C291 VN.n37 B 0.040979f
C292 VN.n38 B 0.295835f
C293 VN.t7 B 0.490777f
C294 VN.t6 B 0.731696f
C295 VN.n39 B 0.29613f
C296 VN.n40 B 0.305495f
C297 VN.n41 B 0.043793f
C298 VN.n42 B 0.052318f
C299 VN.n43 B 0.028071f
C300 VN.n44 B 0.028071f
C301 VN.n45 B 0.028071f
C302 VN.n46 B 0.040979f
C303 VN.n47 B 0.052318f
C304 VN.n48 B 0.043793f
C305 VN.n49 B 0.028071f
C306 VN.n50 B 0.028071f
C307 VN.n51 B 0.028071f
C308 VN.n52 B 0.052318f
C309 VN.n53 B 0.05257f
C310 VN.n54 B 0.025088f
C311 VN.n55 B 0.028071f
C312 VN.n56 B 0.028071f
C313 VN.n57 B 0.028071f
C314 VN.n58 B 0.052318f
C315 VN.n59 B 0.026745f
C316 VN.n60 B 0.30262f
C317 VN.n61 B 1.34538f
.ends

