* NGSPICE file created from diff_pair_sample_0685.ext - technology: sky130A

.subckt diff_pair_sample_0685 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t9 VP.t0 VTAIL.t15 w_n2146_n1476# sky130_fd_pr__pfet_01v8 ad=0.4191 pd=2.87 as=0.9906 ps=5.86 w=2.54 l=0.65
X1 VDD2.t9 VN.t0 VTAIL.t0 w_n2146_n1476# sky130_fd_pr__pfet_01v8 ad=0.4191 pd=2.87 as=0.4191 ps=2.87 w=2.54 l=0.65
X2 VDD1.t8 VP.t1 VTAIL.t13 w_n2146_n1476# sky130_fd_pr__pfet_01v8 ad=0.4191 pd=2.87 as=0.4191 ps=2.87 w=2.54 l=0.65
X3 VTAIL.t19 VN.t1 VDD2.t8 w_n2146_n1476# sky130_fd_pr__pfet_01v8 ad=0.4191 pd=2.87 as=0.4191 ps=2.87 w=2.54 l=0.65
X4 VDD2.t7 VN.t2 VTAIL.t1 w_n2146_n1476# sky130_fd_pr__pfet_01v8 ad=0.9906 pd=5.86 as=0.4191 ps=2.87 w=2.54 l=0.65
X5 VDD1.t7 VP.t2 VTAIL.t9 w_n2146_n1476# sky130_fd_pr__pfet_01v8 ad=0.4191 pd=2.87 as=0.9906 ps=5.86 w=2.54 l=0.65
X6 B.t11 B.t9 B.t10 w_n2146_n1476# sky130_fd_pr__pfet_01v8 ad=0.9906 pd=5.86 as=0 ps=0 w=2.54 l=0.65
X7 VDD1.t6 VP.t3 VTAIL.t17 w_n2146_n1476# sky130_fd_pr__pfet_01v8 ad=0.9906 pd=5.86 as=0.4191 ps=2.87 w=2.54 l=0.65
X8 VDD2.t6 VN.t3 VTAIL.t8 w_n2146_n1476# sky130_fd_pr__pfet_01v8 ad=0.9906 pd=5.86 as=0.4191 ps=2.87 w=2.54 l=0.65
X9 VTAIL.t7 VN.t4 VDD2.t5 w_n2146_n1476# sky130_fd_pr__pfet_01v8 ad=0.4191 pd=2.87 as=0.4191 ps=2.87 w=2.54 l=0.65
X10 VTAIL.t16 VP.t4 VDD1.t5 w_n2146_n1476# sky130_fd_pr__pfet_01v8 ad=0.4191 pd=2.87 as=0.4191 ps=2.87 w=2.54 l=0.65
X11 VDD2.t4 VN.t5 VTAIL.t4 w_n2146_n1476# sky130_fd_pr__pfet_01v8 ad=0.4191 pd=2.87 as=0.9906 ps=5.86 w=2.54 l=0.65
X12 VTAIL.t6 VN.t6 VDD2.t3 w_n2146_n1476# sky130_fd_pr__pfet_01v8 ad=0.4191 pd=2.87 as=0.4191 ps=2.87 w=2.54 l=0.65
X13 VTAIL.t18 VP.t5 VDD1.t4 w_n2146_n1476# sky130_fd_pr__pfet_01v8 ad=0.4191 pd=2.87 as=0.4191 ps=2.87 w=2.54 l=0.65
X14 VTAIL.t2 VN.t7 VDD2.t2 w_n2146_n1476# sky130_fd_pr__pfet_01v8 ad=0.4191 pd=2.87 as=0.4191 ps=2.87 w=2.54 l=0.65
X15 VTAIL.t11 VP.t6 VDD1.t3 w_n2146_n1476# sky130_fd_pr__pfet_01v8 ad=0.4191 pd=2.87 as=0.4191 ps=2.87 w=2.54 l=0.65
X16 B.t8 B.t6 B.t7 w_n2146_n1476# sky130_fd_pr__pfet_01v8 ad=0.9906 pd=5.86 as=0 ps=0 w=2.54 l=0.65
X17 B.t5 B.t3 B.t4 w_n2146_n1476# sky130_fd_pr__pfet_01v8 ad=0.9906 pd=5.86 as=0 ps=0 w=2.54 l=0.65
X18 VDD1.t2 VP.t7 VTAIL.t10 w_n2146_n1476# sky130_fd_pr__pfet_01v8 ad=0.4191 pd=2.87 as=0.4191 ps=2.87 w=2.54 l=0.65
X19 B.t2 B.t0 B.t1 w_n2146_n1476# sky130_fd_pr__pfet_01v8 ad=0.9906 pd=5.86 as=0 ps=0 w=2.54 l=0.65
X20 VDD1.t1 VP.t8 VTAIL.t14 w_n2146_n1476# sky130_fd_pr__pfet_01v8 ad=0.9906 pd=5.86 as=0.4191 ps=2.87 w=2.54 l=0.65
X21 VDD2.t1 VN.t8 VTAIL.t3 w_n2146_n1476# sky130_fd_pr__pfet_01v8 ad=0.4191 pd=2.87 as=0.4191 ps=2.87 w=2.54 l=0.65
X22 VDD2.t0 VN.t9 VTAIL.t5 w_n2146_n1476# sky130_fd_pr__pfet_01v8 ad=0.4191 pd=2.87 as=0.9906 ps=5.86 w=2.54 l=0.65
X23 VTAIL.t12 VP.t9 VDD1.t0 w_n2146_n1476# sky130_fd_pr__pfet_01v8 ad=0.4191 pd=2.87 as=0.4191 ps=2.87 w=2.54 l=0.65
R0 VP.n4 VP.t3 181.433
R1 VP.n17 VP.n16 161.3
R2 VP.n9 VP.n8 161.3
R3 VP.n11 VP.n10 161.3
R4 VP.n10 VP.t8 154.612
R5 VP.n1 VP.t6 154.612
R6 VP.n14 VP.t1 154.612
R7 VP.n15 VP.t5 154.612
R8 VP.n16 VP.t2 154.612
R9 VP.n8 VP.t0 154.612
R10 VP.n7 VP.t4 154.612
R11 VP.n6 VP.t7 154.612
R12 VP.n5 VP.t9 154.612
R13 VP.n6 VP.n3 80.6037
R14 VP.n7 VP.n2 80.6037
R15 VP.n15 VP.n0 80.6037
R16 VP.n14 VP.n13 80.6037
R17 VP.n12 VP.n1 80.6037
R18 VP.n10 VP.n1 48.2005
R19 VP.n14 VP.n1 48.2005
R20 VP.n15 VP.n14 48.2005
R21 VP.n16 VP.n15 48.2005
R22 VP.n8 VP.n7 48.2005
R23 VP.n7 VP.n6 48.2005
R24 VP.n6 VP.n5 48.2005
R25 VP.n4 VP.n3 45.2318
R26 VP.n11 VP.n9 35.4475
R27 VP.n5 VP.n4 13.3799
R28 VP.n3 VP.n2 0.380177
R29 VP.n13 VP.n12 0.380177
R30 VP.n13 VP.n0 0.380177
R31 VP.n9 VP.n2 0.285035
R32 VP.n12 VP.n11 0.285035
R33 VP.n17 VP.n0 0.285035
R34 VP VP.n17 0.0516364
R35 VTAIL.n56 VTAIL.n50 756.745
R36 VTAIL.n8 VTAIL.n2 756.745
R37 VTAIL.n44 VTAIL.n38 756.745
R38 VTAIL.n28 VTAIL.n22 756.745
R39 VTAIL.n55 VTAIL.n54 585
R40 VTAIL.n57 VTAIL.n56 585
R41 VTAIL.n7 VTAIL.n6 585
R42 VTAIL.n9 VTAIL.n8 585
R43 VTAIL.n45 VTAIL.n44 585
R44 VTAIL.n43 VTAIL.n42 585
R45 VTAIL.n29 VTAIL.n28 585
R46 VTAIL.n27 VTAIL.n26 585
R47 VTAIL.n53 VTAIL.t5 355.474
R48 VTAIL.n5 VTAIL.t9 355.474
R49 VTAIL.n41 VTAIL.t15 355.474
R50 VTAIL.n25 VTAIL.t4 355.474
R51 VTAIL.n56 VTAIL.n55 171.744
R52 VTAIL.n8 VTAIL.n7 171.744
R53 VTAIL.n44 VTAIL.n43 171.744
R54 VTAIL.n28 VTAIL.n27 171.744
R55 VTAIL.n37 VTAIL.n36 137.756
R56 VTAIL.n35 VTAIL.n34 137.756
R57 VTAIL.n21 VTAIL.n20 137.756
R58 VTAIL.n19 VTAIL.n18 137.756
R59 VTAIL.n63 VTAIL.n62 137.756
R60 VTAIL.n1 VTAIL.n0 137.756
R61 VTAIL.n15 VTAIL.n14 137.756
R62 VTAIL.n17 VTAIL.n16 137.756
R63 VTAIL.n55 VTAIL.t5 85.8723
R64 VTAIL.n7 VTAIL.t9 85.8723
R65 VTAIL.n43 VTAIL.t15 85.8723
R66 VTAIL.n27 VTAIL.t4 85.8723
R67 VTAIL.n61 VTAIL.n60 34.9005
R68 VTAIL.n13 VTAIL.n12 34.9005
R69 VTAIL.n49 VTAIL.n48 34.9005
R70 VTAIL.n33 VTAIL.n32 34.9005
R71 VTAIL.n19 VTAIL.n17 16.2462
R72 VTAIL.n54 VTAIL.n53 15.8418
R73 VTAIL.n6 VTAIL.n5 15.8418
R74 VTAIL.n42 VTAIL.n41 15.8418
R75 VTAIL.n26 VTAIL.n25 15.8418
R76 VTAIL.n61 VTAIL.n49 15.4014
R77 VTAIL.n57 VTAIL.n52 12.8005
R78 VTAIL.n9 VTAIL.n4 12.8005
R79 VTAIL.n45 VTAIL.n40 12.8005
R80 VTAIL.n29 VTAIL.n24 12.8005
R81 VTAIL.n62 VTAIL.t0 12.7977
R82 VTAIL.n62 VTAIL.t7 12.7977
R83 VTAIL.n0 VTAIL.t1 12.7977
R84 VTAIL.n0 VTAIL.t6 12.7977
R85 VTAIL.n14 VTAIL.t13 12.7977
R86 VTAIL.n14 VTAIL.t18 12.7977
R87 VTAIL.n16 VTAIL.t14 12.7977
R88 VTAIL.n16 VTAIL.t11 12.7977
R89 VTAIL.n36 VTAIL.t10 12.7977
R90 VTAIL.n36 VTAIL.t16 12.7977
R91 VTAIL.n34 VTAIL.t17 12.7977
R92 VTAIL.n34 VTAIL.t12 12.7977
R93 VTAIL.n20 VTAIL.t3 12.7977
R94 VTAIL.n20 VTAIL.t19 12.7977
R95 VTAIL.n18 VTAIL.t8 12.7977
R96 VTAIL.n18 VTAIL.t2 12.7977
R97 VTAIL.n58 VTAIL.n50 12.0247
R98 VTAIL.n10 VTAIL.n2 12.0247
R99 VTAIL.n46 VTAIL.n38 12.0247
R100 VTAIL.n30 VTAIL.n22 12.0247
R101 VTAIL.n60 VTAIL.n59 9.45567
R102 VTAIL.n12 VTAIL.n11 9.45567
R103 VTAIL.n48 VTAIL.n47 9.45567
R104 VTAIL.n32 VTAIL.n31 9.45567
R105 VTAIL.n59 VTAIL.n58 9.3005
R106 VTAIL.n52 VTAIL.n51 9.3005
R107 VTAIL.n11 VTAIL.n10 9.3005
R108 VTAIL.n4 VTAIL.n3 9.3005
R109 VTAIL.n47 VTAIL.n46 9.3005
R110 VTAIL.n40 VTAIL.n39 9.3005
R111 VTAIL.n31 VTAIL.n30 9.3005
R112 VTAIL.n24 VTAIL.n23 9.3005
R113 VTAIL.n41 VTAIL.n39 4.29255
R114 VTAIL.n25 VTAIL.n23 4.29255
R115 VTAIL.n53 VTAIL.n51 4.29255
R116 VTAIL.n5 VTAIL.n3 4.29255
R117 VTAIL.n60 VTAIL.n50 1.93989
R118 VTAIL.n12 VTAIL.n2 1.93989
R119 VTAIL.n48 VTAIL.n38 1.93989
R120 VTAIL.n32 VTAIL.n22 1.93989
R121 VTAIL.n58 VTAIL.n57 1.16414
R122 VTAIL.n10 VTAIL.n9 1.16414
R123 VTAIL.n46 VTAIL.n45 1.16414
R124 VTAIL.n30 VTAIL.n29 1.16414
R125 VTAIL.n35 VTAIL.n33 0.892741
R126 VTAIL.n13 VTAIL.n1 0.892741
R127 VTAIL.n21 VTAIL.n19 0.845328
R128 VTAIL.n33 VTAIL.n21 0.845328
R129 VTAIL.n37 VTAIL.n35 0.845328
R130 VTAIL.n49 VTAIL.n37 0.845328
R131 VTAIL.n17 VTAIL.n15 0.845328
R132 VTAIL.n15 VTAIL.n13 0.845328
R133 VTAIL.n63 VTAIL.n61 0.845328
R134 VTAIL VTAIL.n1 0.69231
R135 VTAIL.n54 VTAIL.n52 0.388379
R136 VTAIL.n6 VTAIL.n4 0.388379
R137 VTAIL.n42 VTAIL.n40 0.388379
R138 VTAIL.n26 VTAIL.n24 0.388379
R139 VTAIL.n59 VTAIL.n51 0.155672
R140 VTAIL.n11 VTAIL.n3 0.155672
R141 VTAIL.n47 VTAIL.n39 0.155672
R142 VTAIL.n31 VTAIL.n23 0.155672
R143 VTAIL VTAIL.n63 0.153517
R144 VDD1.n6 VDD1.n0 756.745
R145 VDD1.n19 VDD1.n13 756.745
R146 VDD1.n7 VDD1.n6 585
R147 VDD1.n5 VDD1.n4 585
R148 VDD1.n18 VDD1.n17 585
R149 VDD1.n20 VDD1.n19 585
R150 VDD1.n3 VDD1.t6 355.474
R151 VDD1.n16 VDD1.t1 355.474
R152 VDD1.n6 VDD1.n5 171.744
R153 VDD1.n19 VDD1.n18 171.744
R154 VDD1.n27 VDD1.n26 155.013
R155 VDD1.n12 VDD1.n11 154.435
R156 VDD1.n29 VDD1.n28 154.435
R157 VDD1.n25 VDD1.n24 154.435
R158 VDD1.n5 VDD1.t6 85.8723
R159 VDD1.n18 VDD1.t1 85.8723
R160 VDD1.n12 VDD1.n10 52.4241
R161 VDD1.n25 VDD1.n23 52.4241
R162 VDD1.n29 VDD1.n27 30.9233
R163 VDD1.n4 VDD1.n3 15.8418
R164 VDD1.n17 VDD1.n16 15.8418
R165 VDD1.n7 VDD1.n2 12.8005
R166 VDD1.n20 VDD1.n15 12.8005
R167 VDD1.n28 VDD1.t5 12.7977
R168 VDD1.n28 VDD1.t9 12.7977
R169 VDD1.n11 VDD1.t0 12.7977
R170 VDD1.n11 VDD1.t2 12.7977
R171 VDD1.n26 VDD1.t4 12.7977
R172 VDD1.n26 VDD1.t7 12.7977
R173 VDD1.n24 VDD1.t3 12.7977
R174 VDD1.n24 VDD1.t8 12.7977
R175 VDD1.n8 VDD1.n0 12.0247
R176 VDD1.n21 VDD1.n13 12.0247
R177 VDD1.n10 VDD1.n9 9.45567
R178 VDD1.n23 VDD1.n22 9.45567
R179 VDD1.n9 VDD1.n8 9.3005
R180 VDD1.n2 VDD1.n1 9.3005
R181 VDD1.n22 VDD1.n21 9.3005
R182 VDD1.n15 VDD1.n14 9.3005
R183 VDD1.n3 VDD1.n1 4.29255
R184 VDD1.n16 VDD1.n14 4.29255
R185 VDD1.n10 VDD1.n0 1.93989
R186 VDD1.n23 VDD1.n13 1.93989
R187 VDD1.n8 VDD1.n7 1.16414
R188 VDD1.n21 VDD1.n20 1.16414
R189 VDD1 VDD1.n29 0.575931
R190 VDD1.n4 VDD1.n2 0.388379
R191 VDD1.n17 VDD1.n15 0.388379
R192 VDD1 VDD1.n12 0.269897
R193 VDD1.n27 VDD1.n25 0.156361
R194 VDD1.n9 VDD1.n1 0.155672
R195 VDD1.n22 VDD1.n14 0.155672
R196 VN.n2 VN.t2 181.433
R197 VN.n10 VN.t5 181.433
R198 VN.n7 VN.n6 161.3
R199 VN.n15 VN.n14 161.3
R200 VN.n1 VN.t6 154.612
R201 VN.n4 VN.t0 154.612
R202 VN.n5 VN.t4 154.612
R203 VN.n6 VN.t9 154.612
R204 VN.n9 VN.t1 154.612
R205 VN.n12 VN.t8 154.612
R206 VN.n13 VN.t7 154.612
R207 VN.n14 VN.t3 154.612
R208 VN.n13 VN.n8 80.6037
R209 VN.n12 VN.n11 80.6037
R210 VN.n5 VN.n0 80.6037
R211 VN.n4 VN.n3 80.6037
R212 VN.n4 VN.n1 48.2005
R213 VN.n5 VN.n4 48.2005
R214 VN.n6 VN.n5 48.2005
R215 VN.n12 VN.n9 48.2005
R216 VN.n13 VN.n12 48.2005
R217 VN.n14 VN.n13 48.2005
R218 VN.n11 VN.n10 45.2318
R219 VN.n3 VN.n2 45.2318
R220 VN VN.n15 35.8282
R221 VN.n10 VN.n9 13.3799
R222 VN.n2 VN.n1 13.3799
R223 VN.n11 VN.n8 0.380177
R224 VN.n3 VN.n0 0.380177
R225 VN.n15 VN.n8 0.285035
R226 VN.n7 VN.n0 0.285035
R227 VN VN.n7 0.0516364
R228 VDD2.n21 VDD2.n15 756.745
R229 VDD2.n6 VDD2.n0 756.745
R230 VDD2.n22 VDD2.n21 585
R231 VDD2.n20 VDD2.n19 585
R232 VDD2.n5 VDD2.n4 585
R233 VDD2.n7 VDD2.n6 585
R234 VDD2.n18 VDD2.t6 355.474
R235 VDD2.n3 VDD2.t7 355.474
R236 VDD2.n21 VDD2.n20 171.744
R237 VDD2.n6 VDD2.n5 171.744
R238 VDD2.n14 VDD2.n13 155.013
R239 VDD2 VDD2.n29 155.011
R240 VDD2.n28 VDD2.n27 154.435
R241 VDD2.n12 VDD2.n11 154.435
R242 VDD2.n20 VDD2.t6 85.8723
R243 VDD2.n5 VDD2.t7 85.8723
R244 VDD2.n12 VDD2.n10 52.4241
R245 VDD2.n26 VDD2.n25 51.5793
R246 VDD2.n26 VDD2.n14 29.9179
R247 VDD2.n19 VDD2.n18 15.8418
R248 VDD2.n4 VDD2.n3 15.8418
R249 VDD2.n22 VDD2.n17 12.8005
R250 VDD2.n7 VDD2.n2 12.8005
R251 VDD2.n29 VDD2.t8 12.7977
R252 VDD2.n29 VDD2.t4 12.7977
R253 VDD2.n27 VDD2.t2 12.7977
R254 VDD2.n27 VDD2.t1 12.7977
R255 VDD2.n13 VDD2.t5 12.7977
R256 VDD2.n13 VDD2.t0 12.7977
R257 VDD2.n11 VDD2.t3 12.7977
R258 VDD2.n11 VDD2.t9 12.7977
R259 VDD2.n23 VDD2.n15 12.0247
R260 VDD2.n8 VDD2.n0 12.0247
R261 VDD2.n25 VDD2.n24 9.45567
R262 VDD2.n10 VDD2.n9 9.45567
R263 VDD2.n24 VDD2.n23 9.3005
R264 VDD2.n17 VDD2.n16 9.3005
R265 VDD2.n9 VDD2.n8 9.3005
R266 VDD2.n2 VDD2.n1 9.3005
R267 VDD2.n18 VDD2.n16 4.29255
R268 VDD2.n3 VDD2.n1 4.29255
R269 VDD2.n25 VDD2.n15 1.93989
R270 VDD2.n10 VDD2.n0 1.93989
R271 VDD2.n23 VDD2.n22 1.16414
R272 VDD2.n8 VDD2.n7 1.16414
R273 VDD2.n28 VDD2.n26 0.845328
R274 VDD2.n19 VDD2.n17 0.388379
R275 VDD2.n4 VDD2.n2 0.388379
R276 VDD2 VDD2.n28 0.269897
R277 VDD2.n14 VDD2.n12 0.156361
R278 VDD2.n24 VDD2.n16 0.155672
R279 VDD2.n9 VDD2.n1 0.155672
R280 B.n191 B.n190 585
R281 B.n189 B.n64 585
R282 B.n188 B.n187 585
R283 B.n186 B.n65 585
R284 B.n185 B.n184 585
R285 B.n183 B.n66 585
R286 B.n182 B.n181 585
R287 B.n180 B.n67 585
R288 B.n179 B.n178 585
R289 B.n177 B.n68 585
R290 B.n176 B.n175 585
R291 B.n174 B.n69 585
R292 B.n173 B.n172 585
R293 B.n171 B.n70 585
R294 B.n170 B.n169 585
R295 B.n165 B.n71 585
R296 B.n164 B.n163 585
R297 B.n162 B.n72 585
R298 B.n161 B.n160 585
R299 B.n159 B.n73 585
R300 B.n158 B.n157 585
R301 B.n156 B.n74 585
R302 B.n155 B.n154 585
R303 B.n152 B.n75 585
R304 B.n151 B.n150 585
R305 B.n149 B.n78 585
R306 B.n148 B.n147 585
R307 B.n146 B.n79 585
R308 B.n145 B.n144 585
R309 B.n143 B.n80 585
R310 B.n142 B.n141 585
R311 B.n140 B.n81 585
R312 B.n139 B.n138 585
R313 B.n137 B.n82 585
R314 B.n136 B.n135 585
R315 B.n134 B.n83 585
R316 B.n133 B.n132 585
R317 B.n192 B.n63 585
R318 B.n194 B.n193 585
R319 B.n195 B.n62 585
R320 B.n197 B.n196 585
R321 B.n198 B.n61 585
R322 B.n200 B.n199 585
R323 B.n201 B.n60 585
R324 B.n203 B.n202 585
R325 B.n204 B.n59 585
R326 B.n206 B.n205 585
R327 B.n207 B.n58 585
R328 B.n209 B.n208 585
R329 B.n210 B.n57 585
R330 B.n212 B.n211 585
R331 B.n213 B.n56 585
R332 B.n215 B.n214 585
R333 B.n216 B.n55 585
R334 B.n218 B.n217 585
R335 B.n219 B.n54 585
R336 B.n221 B.n220 585
R337 B.n222 B.n53 585
R338 B.n224 B.n223 585
R339 B.n225 B.n52 585
R340 B.n227 B.n226 585
R341 B.n228 B.n51 585
R342 B.n230 B.n229 585
R343 B.n231 B.n50 585
R344 B.n233 B.n232 585
R345 B.n234 B.n49 585
R346 B.n236 B.n235 585
R347 B.n237 B.n48 585
R348 B.n239 B.n238 585
R349 B.n240 B.n47 585
R350 B.n242 B.n241 585
R351 B.n243 B.n46 585
R352 B.n245 B.n244 585
R353 B.n246 B.n45 585
R354 B.n248 B.n247 585
R355 B.n249 B.n44 585
R356 B.n251 B.n250 585
R357 B.n252 B.n43 585
R358 B.n254 B.n253 585
R359 B.n255 B.n42 585
R360 B.n257 B.n256 585
R361 B.n258 B.n41 585
R362 B.n260 B.n259 585
R363 B.n261 B.n40 585
R364 B.n263 B.n262 585
R365 B.n264 B.n39 585
R366 B.n266 B.n265 585
R367 B.n267 B.n38 585
R368 B.n269 B.n268 585
R369 B.n326 B.n325 585
R370 B.n324 B.n15 585
R371 B.n323 B.n322 585
R372 B.n321 B.n16 585
R373 B.n320 B.n319 585
R374 B.n318 B.n17 585
R375 B.n317 B.n316 585
R376 B.n315 B.n18 585
R377 B.n314 B.n313 585
R378 B.n312 B.n19 585
R379 B.n311 B.n310 585
R380 B.n309 B.n20 585
R381 B.n308 B.n307 585
R382 B.n306 B.n21 585
R383 B.n304 B.n303 585
R384 B.n302 B.n24 585
R385 B.n301 B.n300 585
R386 B.n299 B.n25 585
R387 B.n298 B.n297 585
R388 B.n296 B.n26 585
R389 B.n295 B.n294 585
R390 B.n293 B.n27 585
R391 B.n292 B.n291 585
R392 B.n290 B.n289 585
R393 B.n288 B.n31 585
R394 B.n287 B.n286 585
R395 B.n285 B.n32 585
R396 B.n284 B.n283 585
R397 B.n282 B.n33 585
R398 B.n281 B.n280 585
R399 B.n279 B.n34 585
R400 B.n278 B.n277 585
R401 B.n276 B.n35 585
R402 B.n275 B.n274 585
R403 B.n273 B.n36 585
R404 B.n272 B.n271 585
R405 B.n270 B.n37 585
R406 B.n327 B.n14 585
R407 B.n329 B.n328 585
R408 B.n330 B.n13 585
R409 B.n332 B.n331 585
R410 B.n333 B.n12 585
R411 B.n335 B.n334 585
R412 B.n336 B.n11 585
R413 B.n338 B.n337 585
R414 B.n339 B.n10 585
R415 B.n341 B.n340 585
R416 B.n342 B.n9 585
R417 B.n344 B.n343 585
R418 B.n345 B.n8 585
R419 B.n347 B.n346 585
R420 B.n348 B.n7 585
R421 B.n350 B.n349 585
R422 B.n351 B.n6 585
R423 B.n353 B.n352 585
R424 B.n354 B.n5 585
R425 B.n356 B.n355 585
R426 B.n357 B.n4 585
R427 B.n359 B.n358 585
R428 B.n360 B.n3 585
R429 B.n362 B.n361 585
R430 B.n363 B.n0 585
R431 B.n2 B.n1 585
R432 B.n97 B.n96 585
R433 B.n98 B.n95 585
R434 B.n100 B.n99 585
R435 B.n101 B.n94 585
R436 B.n103 B.n102 585
R437 B.n104 B.n93 585
R438 B.n106 B.n105 585
R439 B.n107 B.n92 585
R440 B.n109 B.n108 585
R441 B.n110 B.n91 585
R442 B.n112 B.n111 585
R443 B.n113 B.n90 585
R444 B.n115 B.n114 585
R445 B.n116 B.n89 585
R446 B.n118 B.n117 585
R447 B.n119 B.n88 585
R448 B.n121 B.n120 585
R449 B.n122 B.n87 585
R450 B.n124 B.n123 585
R451 B.n125 B.n86 585
R452 B.n127 B.n126 585
R453 B.n128 B.n85 585
R454 B.n130 B.n129 585
R455 B.n131 B.n84 585
R456 B.n132 B.n131 497.305
R457 B.n190 B.n63 497.305
R458 B.n268 B.n37 497.305
R459 B.n327 B.n326 497.305
R460 B.n76 B.t9 297.803
R461 B.n166 B.t3 297.803
R462 B.n28 B.t0 297.803
R463 B.n22 B.t6 297.803
R464 B.n365 B.n364 256.663
R465 B.n166 B.t4 244.034
R466 B.n28 B.t2 244.034
R467 B.n76 B.t10 244.034
R468 B.n22 B.t8 244.034
R469 B.n364 B.n363 235.042
R470 B.n364 B.n2 235.042
R471 B.n167 B.t5 225.028
R472 B.n29 B.t1 225.028
R473 B.n77 B.t11 225.026
R474 B.n23 B.t7 225.026
R475 B.n132 B.n83 163.367
R476 B.n136 B.n83 163.367
R477 B.n137 B.n136 163.367
R478 B.n138 B.n137 163.367
R479 B.n138 B.n81 163.367
R480 B.n142 B.n81 163.367
R481 B.n143 B.n142 163.367
R482 B.n144 B.n143 163.367
R483 B.n144 B.n79 163.367
R484 B.n148 B.n79 163.367
R485 B.n149 B.n148 163.367
R486 B.n150 B.n149 163.367
R487 B.n150 B.n75 163.367
R488 B.n155 B.n75 163.367
R489 B.n156 B.n155 163.367
R490 B.n157 B.n156 163.367
R491 B.n157 B.n73 163.367
R492 B.n161 B.n73 163.367
R493 B.n162 B.n161 163.367
R494 B.n163 B.n162 163.367
R495 B.n163 B.n71 163.367
R496 B.n170 B.n71 163.367
R497 B.n171 B.n170 163.367
R498 B.n172 B.n171 163.367
R499 B.n172 B.n69 163.367
R500 B.n176 B.n69 163.367
R501 B.n177 B.n176 163.367
R502 B.n178 B.n177 163.367
R503 B.n178 B.n67 163.367
R504 B.n182 B.n67 163.367
R505 B.n183 B.n182 163.367
R506 B.n184 B.n183 163.367
R507 B.n184 B.n65 163.367
R508 B.n188 B.n65 163.367
R509 B.n189 B.n188 163.367
R510 B.n190 B.n189 163.367
R511 B.n268 B.n267 163.367
R512 B.n267 B.n266 163.367
R513 B.n266 B.n39 163.367
R514 B.n262 B.n39 163.367
R515 B.n262 B.n261 163.367
R516 B.n261 B.n260 163.367
R517 B.n260 B.n41 163.367
R518 B.n256 B.n41 163.367
R519 B.n256 B.n255 163.367
R520 B.n255 B.n254 163.367
R521 B.n254 B.n43 163.367
R522 B.n250 B.n43 163.367
R523 B.n250 B.n249 163.367
R524 B.n249 B.n248 163.367
R525 B.n248 B.n45 163.367
R526 B.n244 B.n45 163.367
R527 B.n244 B.n243 163.367
R528 B.n243 B.n242 163.367
R529 B.n242 B.n47 163.367
R530 B.n238 B.n47 163.367
R531 B.n238 B.n237 163.367
R532 B.n237 B.n236 163.367
R533 B.n236 B.n49 163.367
R534 B.n232 B.n49 163.367
R535 B.n232 B.n231 163.367
R536 B.n231 B.n230 163.367
R537 B.n230 B.n51 163.367
R538 B.n226 B.n51 163.367
R539 B.n226 B.n225 163.367
R540 B.n225 B.n224 163.367
R541 B.n224 B.n53 163.367
R542 B.n220 B.n53 163.367
R543 B.n220 B.n219 163.367
R544 B.n219 B.n218 163.367
R545 B.n218 B.n55 163.367
R546 B.n214 B.n55 163.367
R547 B.n214 B.n213 163.367
R548 B.n213 B.n212 163.367
R549 B.n212 B.n57 163.367
R550 B.n208 B.n57 163.367
R551 B.n208 B.n207 163.367
R552 B.n207 B.n206 163.367
R553 B.n206 B.n59 163.367
R554 B.n202 B.n59 163.367
R555 B.n202 B.n201 163.367
R556 B.n201 B.n200 163.367
R557 B.n200 B.n61 163.367
R558 B.n196 B.n61 163.367
R559 B.n196 B.n195 163.367
R560 B.n195 B.n194 163.367
R561 B.n194 B.n63 163.367
R562 B.n326 B.n15 163.367
R563 B.n322 B.n15 163.367
R564 B.n322 B.n321 163.367
R565 B.n321 B.n320 163.367
R566 B.n320 B.n17 163.367
R567 B.n316 B.n17 163.367
R568 B.n316 B.n315 163.367
R569 B.n315 B.n314 163.367
R570 B.n314 B.n19 163.367
R571 B.n310 B.n19 163.367
R572 B.n310 B.n309 163.367
R573 B.n309 B.n308 163.367
R574 B.n308 B.n21 163.367
R575 B.n303 B.n21 163.367
R576 B.n303 B.n302 163.367
R577 B.n302 B.n301 163.367
R578 B.n301 B.n25 163.367
R579 B.n297 B.n25 163.367
R580 B.n297 B.n296 163.367
R581 B.n296 B.n295 163.367
R582 B.n295 B.n27 163.367
R583 B.n291 B.n27 163.367
R584 B.n291 B.n290 163.367
R585 B.n290 B.n31 163.367
R586 B.n286 B.n31 163.367
R587 B.n286 B.n285 163.367
R588 B.n285 B.n284 163.367
R589 B.n284 B.n33 163.367
R590 B.n280 B.n33 163.367
R591 B.n280 B.n279 163.367
R592 B.n279 B.n278 163.367
R593 B.n278 B.n35 163.367
R594 B.n274 B.n35 163.367
R595 B.n274 B.n273 163.367
R596 B.n273 B.n272 163.367
R597 B.n272 B.n37 163.367
R598 B.n328 B.n327 163.367
R599 B.n328 B.n13 163.367
R600 B.n332 B.n13 163.367
R601 B.n333 B.n332 163.367
R602 B.n334 B.n333 163.367
R603 B.n334 B.n11 163.367
R604 B.n338 B.n11 163.367
R605 B.n339 B.n338 163.367
R606 B.n340 B.n339 163.367
R607 B.n340 B.n9 163.367
R608 B.n344 B.n9 163.367
R609 B.n345 B.n344 163.367
R610 B.n346 B.n345 163.367
R611 B.n346 B.n7 163.367
R612 B.n350 B.n7 163.367
R613 B.n351 B.n350 163.367
R614 B.n352 B.n351 163.367
R615 B.n352 B.n5 163.367
R616 B.n356 B.n5 163.367
R617 B.n357 B.n356 163.367
R618 B.n358 B.n357 163.367
R619 B.n358 B.n3 163.367
R620 B.n362 B.n3 163.367
R621 B.n363 B.n362 163.367
R622 B.n96 B.n2 163.367
R623 B.n96 B.n95 163.367
R624 B.n100 B.n95 163.367
R625 B.n101 B.n100 163.367
R626 B.n102 B.n101 163.367
R627 B.n102 B.n93 163.367
R628 B.n106 B.n93 163.367
R629 B.n107 B.n106 163.367
R630 B.n108 B.n107 163.367
R631 B.n108 B.n91 163.367
R632 B.n112 B.n91 163.367
R633 B.n113 B.n112 163.367
R634 B.n114 B.n113 163.367
R635 B.n114 B.n89 163.367
R636 B.n118 B.n89 163.367
R637 B.n119 B.n118 163.367
R638 B.n120 B.n119 163.367
R639 B.n120 B.n87 163.367
R640 B.n124 B.n87 163.367
R641 B.n125 B.n124 163.367
R642 B.n126 B.n125 163.367
R643 B.n126 B.n85 163.367
R644 B.n130 B.n85 163.367
R645 B.n131 B.n130 163.367
R646 B.n153 B.n77 59.5399
R647 B.n168 B.n167 59.5399
R648 B.n30 B.n29 59.5399
R649 B.n305 B.n23 59.5399
R650 B.n325 B.n14 32.3127
R651 B.n270 B.n269 32.3127
R652 B.n192 B.n191 32.3127
R653 B.n133 B.n84 32.3127
R654 B.n77 B.n76 19.0066
R655 B.n167 B.n166 19.0066
R656 B.n29 B.n28 19.0066
R657 B.n23 B.n22 19.0066
R658 B B.n365 18.0485
R659 B.n329 B.n14 10.6151
R660 B.n330 B.n329 10.6151
R661 B.n331 B.n330 10.6151
R662 B.n331 B.n12 10.6151
R663 B.n335 B.n12 10.6151
R664 B.n336 B.n335 10.6151
R665 B.n337 B.n336 10.6151
R666 B.n337 B.n10 10.6151
R667 B.n341 B.n10 10.6151
R668 B.n342 B.n341 10.6151
R669 B.n343 B.n342 10.6151
R670 B.n343 B.n8 10.6151
R671 B.n347 B.n8 10.6151
R672 B.n348 B.n347 10.6151
R673 B.n349 B.n348 10.6151
R674 B.n349 B.n6 10.6151
R675 B.n353 B.n6 10.6151
R676 B.n354 B.n353 10.6151
R677 B.n355 B.n354 10.6151
R678 B.n355 B.n4 10.6151
R679 B.n359 B.n4 10.6151
R680 B.n360 B.n359 10.6151
R681 B.n361 B.n360 10.6151
R682 B.n361 B.n0 10.6151
R683 B.n325 B.n324 10.6151
R684 B.n324 B.n323 10.6151
R685 B.n323 B.n16 10.6151
R686 B.n319 B.n16 10.6151
R687 B.n319 B.n318 10.6151
R688 B.n318 B.n317 10.6151
R689 B.n317 B.n18 10.6151
R690 B.n313 B.n18 10.6151
R691 B.n313 B.n312 10.6151
R692 B.n312 B.n311 10.6151
R693 B.n311 B.n20 10.6151
R694 B.n307 B.n20 10.6151
R695 B.n307 B.n306 10.6151
R696 B.n304 B.n24 10.6151
R697 B.n300 B.n24 10.6151
R698 B.n300 B.n299 10.6151
R699 B.n299 B.n298 10.6151
R700 B.n298 B.n26 10.6151
R701 B.n294 B.n26 10.6151
R702 B.n294 B.n293 10.6151
R703 B.n293 B.n292 10.6151
R704 B.n289 B.n288 10.6151
R705 B.n288 B.n287 10.6151
R706 B.n287 B.n32 10.6151
R707 B.n283 B.n32 10.6151
R708 B.n283 B.n282 10.6151
R709 B.n282 B.n281 10.6151
R710 B.n281 B.n34 10.6151
R711 B.n277 B.n34 10.6151
R712 B.n277 B.n276 10.6151
R713 B.n276 B.n275 10.6151
R714 B.n275 B.n36 10.6151
R715 B.n271 B.n36 10.6151
R716 B.n271 B.n270 10.6151
R717 B.n269 B.n38 10.6151
R718 B.n265 B.n38 10.6151
R719 B.n265 B.n264 10.6151
R720 B.n264 B.n263 10.6151
R721 B.n263 B.n40 10.6151
R722 B.n259 B.n40 10.6151
R723 B.n259 B.n258 10.6151
R724 B.n258 B.n257 10.6151
R725 B.n257 B.n42 10.6151
R726 B.n253 B.n42 10.6151
R727 B.n253 B.n252 10.6151
R728 B.n252 B.n251 10.6151
R729 B.n251 B.n44 10.6151
R730 B.n247 B.n44 10.6151
R731 B.n247 B.n246 10.6151
R732 B.n246 B.n245 10.6151
R733 B.n245 B.n46 10.6151
R734 B.n241 B.n46 10.6151
R735 B.n241 B.n240 10.6151
R736 B.n240 B.n239 10.6151
R737 B.n239 B.n48 10.6151
R738 B.n235 B.n48 10.6151
R739 B.n235 B.n234 10.6151
R740 B.n234 B.n233 10.6151
R741 B.n233 B.n50 10.6151
R742 B.n229 B.n50 10.6151
R743 B.n229 B.n228 10.6151
R744 B.n228 B.n227 10.6151
R745 B.n227 B.n52 10.6151
R746 B.n223 B.n52 10.6151
R747 B.n223 B.n222 10.6151
R748 B.n222 B.n221 10.6151
R749 B.n221 B.n54 10.6151
R750 B.n217 B.n54 10.6151
R751 B.n217 B.n216 10.6151
R752 B.n216 B.n215 10.6151
R753 B.n215 B.n56 10.6151
R754 B.n211 B.n56 10.6151
R755 B.n211 B.n210 10.6151
R756 B.n210 B.n209 10.6151
R757 B.n209 B.n58 10.6151
R758 B.n205 B.n58 10.6151
R759 B.n205 B.n204 10.6151
R760 B.n204 B.n203 10.6151
R761 B.n203 B.n60 10.6151
R762 B.n199 B.n60 10.6151
R763 B.n199 B.n198 10.6151
R764 B.n198 B.n197 10.6151
R765 B.n197 B.n62 10.6151
R766 B.n193 B.n62 10.6151
R767 B.n193 B.n192 10.6151
R768 B.n97 B.n1 10.6151
R769 B.n98 B.n97 10.6151
R770 B.n99 B.n98 10.6151
R771 B.n99 B.n94 10.6151
R772 B.n103 B.n94 10.6151
R773 B.n104 B.n103 10.6151
R774 B.n105 B.n104 10.6151
R775 B.n105 B.n92 10.6151
R776 B.n109 B.n92 10.6151
R777 B.n110 B.n109 10.6151
R778 B.n111 B.n110 10.6151
R779 B.n111 B.n90 10.6151
R780 B.n115 B.n90 10.6151
R781 B.n116 B.n115 10.6151
R782 B.n117 B.n116 10.6151
R783 B.n117 B.n88 10.6151
R784 B.n121 B.n88 10.6151
R785 B.n122 B.n121 10.6151
R786 B.n123 B.n122 10.6151
R787 B.n123 B.n86 10.6151
R788 B.n127 B.n86 10.6151
R789 B.n128 B.n127 10.6151
R790 B.n129 B.n128 10.6151
R791 B.n129 B.n84 10.6151
R792 B.n134 B.n133 10.6151
R793 B.n135 B.n134 10.6151
R794 B.n135 B.n82 10.6151
R795 B.n139 B.n82 10.6151
R796 B.n140 B.n139 10.6151
R797 B.n141 B.n140 10.6151
R798 B.n141 B.n80 10.6151
R799 B.n145 B.n80 10.6151
R800 B.n146 B.n145 10.6151
R801 B.n147 B.n146 10.6151
R802 B.n147 B.n78 10.6151
R803 B.n151 B.n78 10.6151
R804 B.n152 B.n151 10.6151
R805 B.n154 B.n74 10.6151
R806 B.n158 B.n74 10.6151
R807 B.n159 B.n158 10.6151
R808 B.n160 B.n159 10.6151
R809 B.n160 B.n72 10.6151
R810 B.n164 B.n72 10.6151
R811 B.n165 B.n164 10.6151
R812 B.n169 B.n165 10.6151
R813 B.n173 B.n70 10.6151
R814 B.n174 B.n173 10.6151
R815 B.n175 B.n174 10.6151
R816 B.n175 B.n68 10.6151
R817 B.n179 B.n68 10.6151
R818 B.n180 B.n179 10.6151
R819 B.n181 B.n180 10.6151
R820 B.n181 B.n66 10.6151
R821 B.n185 B.n66 10.6151
R822 B.n186 B.n185 10.6151
R823 B.n187 B.n186 10.6151
R824 B.n187 B.n64 10.6151
R825 B.n191 B.n64 10.6151
R826 B.n365 B.n0 8.11757
R827 B.n365 B.n1 8.11757
R828 B.n305 B.n304 6.5566
R829 B.n292 B.n30 6.5566
R830 B.n154 B.n153 6.5566
R831 B.n169 B.n168 6.5566
R832 B.n306 B.n305 4.05904
R833 B.n289 B.n30 4.05904
R834 B.n153 B.n152 4.05904
R835 B.n168 B.n70 4.05904
C0 VDD2 B 1.03691f
C1 B VTAIL 0.998932f
C2 B VN 0.67615f
C3 VDD2 VTAIL 5.08743f
C4 B VDD1 0.994443f
C5 VP B 1.12454f
C6 B w_n2146_n1476# 4.61117f
C7 VDD2 VN 1.69484f
C8 VTAIL VN 1.9835f
C9 VDD2 VDD1 0.939453f
C10 VTAIL VDD1 5.04836f
C11 VP VDD2 0.340574f
C12 VP VTAIL 1.99771f
C13 VDD2 w_n2146_n1476# 1.35846f
C14 w_n2146_n1476# VTAIL 1.50872f
C15 VDD1 VN 0.155081f
C16 VP VN 3.77198f
C17 VP VDD1 1.87819f
C18 w_n2146_n1476# VN 3.78162f
C19 w_n2146_n1476# VDD1 1.31705f
C20 VP w_n2146_n1476# 4.05184f
C21 VDD2 VSUBS 0.798392f
C22 VDD1 VSUBS 0.812947f
C23 VTAIL VSUBS 0.318573f
C24 VN VSUBS 3.60538f
C25 VP VSUBS 1.292803f
C26 B VSUBS 2.044042f
C27 w_n2146_n1476# VSUBS 40.2504f
C28 B.n0 VSUBS 0.00719f
C29 B.n1 VSUBS 0.00719f
C30 B.n2 VSUBS 0.010633f
C31 B.n3 VSUBS 0.008148f
C32 B.n4 VSUBS 0.008148f
C33 B.n5 VSUBS 0.008148f
C34 B.n6 VSUBS 0.008148f
C35 B.n7 VSUBS 0.008148f
C36 B.n8 VSUBS 0.008148f
C37 B.n9 VSUBS 0.008148f
C38 B.n10 VSUBS 0.008148f
C39 B.n11 VSUBS 0.008148f
C40 B.n12 VSUBS 0.008148f
C41 B.n13 VSUBS 0.008148f
C42 B.n14 VSUBS 0.018612f
C43 B.n15 VSUBS 0.008148f
C44 B.n16 VSUBS 0.008148f
C45 B.n17 VSUBS 0.008148f
C46 B.n18 VSUBS 0.008148f
C47 B.n19 VSUBS 0.008148f
C48 B.n20 VSUBS 0.008148f
C49 B.n21 VSUBS 0.008148f
C50 B.t7 VSUBS 0.045883f
C51 B.t8 VSUBS 0.051626f
C52 B.t6 VSUBS 0.088954f
C53 B.n22 VSUBS 0.091372f
C54 B.n23 VSUBS 0.085368f
C55 B.n24 VSUBS 0.008148f
C56 B.n25 VSUBS 0.008148f
C57 B.n26 VSUBS 0.008148f
C58 B.n27 VSUBS 0.008148f
C59 B.t1 VSUBS 0.045883f
C60 B.t2 VSUBS 0.051627f
C61 B.t0 VSUBS 0.088954f
C62 B.n28 VSUBS 0.091371f
C63 B.n29 VSUBS 0.085368f
C64 B.n30 VSUBS 0.018879f
C65 B.n31 VSUBS 0.008148f
C66 B.n32 VSUBS 0.008148f
C67 B.n33 VSUBS 0.008148f
C68 B.n34 VSUBS 0.008148f
C69 B.n35 VSUBS 0.008148f
C70 B.n36 VSUBS 0.008148f
C71 B.n37 VSUBS 0.019253f
C72 B.n38 VSUBS 0.008148f
C73 B.n39 VSUBS 0.008148f
C74 B.n40 VSUBS 0.008148f
C75 B.n41 VSUBS 0.008148f
C76 B.n42 VSUBS 0.008148f
C77 B.n43 VSUBS 0.008148f
C78 B.n44 VSUBS 0.008148f
C79 B.n45 VSUBS 0.008148f
C80 B.n46 VSUBS 0.008148f
C81 B.n47 VSUBS 0.008148f
C82 B.n48 VSUBS 0.008148f
C83 B.n49 VSUBS 0.008148f
C84 B.n50 VSUBS 0.008148f
C85 B.n51 VSUBS 0.008148f
C86 B.n52 VSUBS 0.008148f
C87 B.n53 VSUBS 0.008148f
C88 B.n54 VSUBS 0.008148f
C89 B.n55 VSUBS 0.008148f
C90 B.n56 VSUBS 0.008148f
C91 B.n57 VSUBS 0.008148f
C92 B.n58 VSUBS 0.008148f
C93 B.n59 VSUBS 0.008148f
C94 B.n60 VSUBS 0.008148f
C95 B.n61 VSUBS 0.008148f
C96 B.n62 VSUBS 0.008148f
C97 B.n63 VSUBS 0.018612f
C98 B.n64 VSUBS 0.008148f
C99 B.n65 VSUBS 0.008148f
C100 B.n66 VSUBS 0.008148f
C101 B.n67 VSUBS 0.008148f
C102 B.n68 VSUBS 0.008148f
C103 B.n69 VSUBS 0.008148f
C104 B.n70 VSUBS 0.005632f
C105 B.n71 VSUBS 0.008148f
C106 B.n72 VSUBS 0.008148f
C107 B.n73 VSUBS 0.008148f
C108 B.n74 VSUBS 0.008148f
C109 B.n75 VSUBS 0.008148f
C110 B.t11 VSUBS 0.045883f
C111 B.t10 VSUBS 0.051626f
C112 B.t9 VSUBS 0.088954f
C113 B.n76 VSUBS 0.091372f
C114 B.n77 VSUBS 0.085368f
C115 B.n78 VSUBS 0.008148f
C116 B.n79 VSUBS 0.008148f
C117 B.n80 VSUBS 0.008148f
C118 B.n81 VSUBS 0.008148f
C119 B.n82 VSUBS 0.008148f
C120 B.n83 VSUBS 0.008148f
C121 B.n84 VSUBS 0.018612f
C122 B.n85 VSUBS 0.008148f
C123 B.n86 VSUBS 0.008148f
C124 B.n87 VSUBS 0.008148f
C125 B.n88 VSUBS 0.008148f
C126 B.n89 VSUBS 0.008148f
C127 B.n90 VSUBS 0.008148f
C128 B.n91 VSUBS 0.008148f
C129 B.n92 VSUBS 0.008148f
C130 B.n93 VSUBS 0.008148f
C131 B.n94 VSUBS 0.008148f
C132 B.n95 VSUBS 0.008148f
C133 B.n96 VSUBS 0.008148f
C134 B.n97 VSUBS 0.008148f
C135 B.n98 VSUBS 0.008148f
C136 B.n99 VSUBS 0.008148f
C137 B.n100 VSUBS 0.008148f
C138 B.n101 VSUBS 0.008148f
C139 B.n102 VSUBS 0.008148f
C140 B.n103 VSUBS 0.008148f
C141 B.n104 VSUBS 0.008148f
C142 B.n105 VSUBS 0.008148f
C143 B.n106 VSUBS 0.008148f
C144 B.n107 VSUBS 0.008148f
C145 B.n108 VSUBS 0.008148f
C146 B.n109 VSUBS 0.008148f
C147 B.n110 VSUBS 0.008148f
C148 B.n111 VSUBS 0.008148f
C149 B.n112 VSUBS 0.008148f
C150 B.n113 VSUBS 0.008148f
C151 B.n114 VSUBS 0.008148f
C152 B.n115 VSUBS 0.008148f
C153 B.n116 VSUBS 0.008148f
C154 B.n117 VSUBS 0.008148f
C155 B.n118 VSUBS 0.008148f
C156 B.n119 VSUBS 0.008148f
C157 B.n120 VSUBS 0.008148f
C158 B.n121 VSUBS 0.008148f
C159 B.n122 VSUBS 0.008148f
C160 B.n123 VSUBS 0.008148f
C161 B.n124 VSUBS 0.008148f
C162 B.n125 VSUBS 0.008148f
C163 B.n126 VSUBS 0.008148f
C164 B.n127 VSUBS 0.008148f
C165 B.n128 VSUBS 0.008148f
C166 B.n129 VSUBS 0.008148f
C167 B.n130 VSUBS 0.008148f
C168 B.n131 VSUBS 0.018612f
C169 B.n132 VSUBS 0.019253f
C170 B.n133 VSUBS 0.019253f
C171 B.n134 VSUBS 0.008148f
C172 B.n135 VSUBS 0.008148f
C173 B.n136 VSUBS 0.008148f
C174 B.n137 VSUBS 0.008148f
C175 B.n138 VSUBS 0.008148f
C176 B.n139 VSUBS 0.008148f
C177 B.n140 VSUBS 0.008148f
C178 B.n141 VSUBS 0.008148f
C179 B.n142 VSUBS 0.008148f
C180 B.n143 VSUBS 0.008148f
C181 B.n144 VSUBS 0.008148f
C182 B.n145 VSUBS 0.008148f
C183 B.n146 VSUBS 0.008148f
C184 B.n147 VSUBS 0.008148f
C185 B.n148 VSUBS 0.008148f
C186 B.n149 VSUBS 0.008148f
C187 B.n150 VSUBS 0.008148f
C188 B.n151 VSUBS 0.008148f
C189 B.n152 VSUBS 0.005632f
C190 B.n153 VSUBS 0.018879f
C191 B.n154 VSUBS 0.006591f
C192 B.n155 VSUBS 0.008148f
C193 B.n156 VSUBS 0.008148f
C194 B.n157 VSUBS 0.008148f
C195 B.n158 VSUBS 0.008148f
C196 B.n159 VSUBS 0.008148f
C197 B.n160 VSUBS 0.008148f
C198 B.n161 VSUBS 0.008148f
C199 B.n162 VSUBS 0.008148f
C200 B.n163 VSUBS 0.008148f
C201 B.n164 VSUBS 0.008148f
C202 B.n165 VSUBS 0.008148f
C203 B.t5 VSUBS 0.045883f
C204 B.t4 VSUBS 0.051627f
C205 B.t3 VSUBS 0.088954f
C206 B.n166 VSUBS 0.091371f
C207 B.n167 VSUBS 0.085368f
C208 B.n168 VSUBS 0.018879f
C209 B.n169 VSUBS 0.006591f
C210 B.n170 VSUBS 0.008148f
C211 B.n171 VSUBS 0.008148f
C212 B.n172 VSUBS 0.008148f
C213 B.n173 VSUBS 0.008148f
C214 B.n174 VSUBS 0.008148f
C215 B.n175 VSUBS 0.008148f
C216 B.n176 VSUBS 0.008148f
C217 B.n177 VSUBS 0.008148f
C218 B.n178 VSUBS 0.008148f
C219 B.n179 VSUBS 0.008148f
C220 B.n180 VSUBS 0.008148f
C221 B.n181 VSUBS 0.008148f
C222 B.n182 VSUBS 0.008148f
C223 B.n183 VSUBS 0.008148f
C224 B.n184 VSUBS 0.008148f
C225 B.n185 VSUBS 0.008148f
C226 B.n186 VSUBS 0.008148f
C227 B.n187 VSUBS 0.008148f
C228 B.n188 VSUBS 0.008148f
C229 B.n189 VSUBS 0.008148f
C230 B.n190 VSUBS 0.019253f
C231 B.n191 VSUBS 0.01828f
C232 B.n192 VSUBS 0.019586f
C233 B.n193 VSUBS 0.008148f
C234 B.n194 VSUBS 0.008148f
C235 B.n195 VSUBS 0.008148f
C236 B.n196 VSUBS 0.008148f
C237 B.n197 VSUBS 0.008148f
C238 B.n198 VSUBS 0.008148f
C239 B.n199 VSUBS 0.008148f
C240 B.n200 VSUBS 0.008148f
C241 B.n201 VSUBS 0.008148f
C242 B.n202 VSUBS 0.008148f
C243 B.n203 VSUBS 0.008148f
C244 B.n204 VSUBS 0.008148f
C245 B.n205 VSUBS 0.008148f
C246 B.n206 VSUBS 0.008148f
C247 B.n207 VSUBS 0.008148f
C248 B.n208 VSUBS 0.008148f
C249 B.n209 VSUBS 0.008148f
C250 B.n210 VSUBS 0.008148f
C251 B.n211 VSUBS 0.008148f
C252 B.n212 VSUBS 0.008148f
C253 B.n213 VSUBS 0.008148f
C254 B.n214 VSUBS 0.008148f
C255 B.n215 VSUBS 0.008148f
C256 B.n216 VSUBS 0.008148f
C257 B.n217 VSUBS 0.008148f
C258 B.n218 VSUBS 0.008148f
C259 B.n219 VSUBS 0.008148f
C260 B.n220 VSUBS 0.008148f
C261 B.n221 VSUBS 0.008148f
C262 B.n222 VSUBS 0.008148f
C263 B.n223 VSUBS 0.008148f
C264 B.n224 VSUBS 0.008148f
C265 B.n225 VSUBS 0.008148f
C266 B.n226 VSUBS 0.008148f
C267 B.n227 VSUBS 0.008148f
C268 B.n228 VSUBS 0.008148f
C269 B.n229 VSUBS 0.008148f
C270 B.n230 VSUBS 0.008148f
C271 B.n231 VSUBS 0.008148f
C272 B.n232 VSUBS 0.008148f
C273 B.n233 VSUBS 0.008148f
C274 B.n234 VSUBS 0.008148f
C275 B.n235 VSUBS 0.008148f
C276 B.n236 VSUBS 0.008148f
C277 B.n237 VSUBS 0.008148f
C278 B.n238 VSUBS 0.008148f
C279 B.n239 VSUBS 0.008148f
C280 B.n240 VSUBS 0.008148f
C281 B.n241 VSUBS 0.008148f
C282 B.n242 VSUBS 0.008148f
C283 B.n243 VSUBS 0.008148f
C284 B.n244 VSUBS 0.008148f
C285 B.n245 VSUBS 0.008148f
C286 B.n246 VSUBS 0.008148f
C287 B.n247 VSUBS 0.008148f
C288 B.n248 VSUBS 0.008148f
C289 B.n249 VSUBS 0.008148f
C290 B.n250 VSUBS 0.008148f
C291 B.n251 VSUBS 0.008148f
C292 B.n252 VSUBS 0.008148f
C293 B.n253 VSUBS 0.008148f
C294 B.n254 VSUBS 0.008148f
C295 B.n255 VSUBS 0.008148f
C296 B.n256 VSUBS 0.008148f
C297 B.n257 VSUBS 0.008148f
C298 B.n258 VSUBS 0.008148f
C299 B.n259 VSUBS 0.008148f
C300 B.n260 VSUBS 0.008148f
C301 B.n261 VSUBS 0.008148f
C302 B.n262 VSUBS 0.008148f
C303 B.n263 VSUBS 0.008148f
C304 B.n264 VSUBS 0.008148f
C305 B.n265 VSUBS 0.008148f
C306 B.n266 VSUBS 0.008148f
C307 B.n267 VSUBS 0.008148f
C308 B.n268 VSUBS 0.018612f
C309 B.n269 VSUBS 0.018612f
C310 B.n270 VSUBS 0.019253f
C311 B.n271 VSUBS 0.008148f
C312 B.n272 VSUBS 0.008148f
C313 B.n273 VSUBS 0.008148f
C314 B.n274 VSUBS 0.008148f
C315 B.n275 VSUBS 0.008148f
C316 B.n276 VSUBS 0.008148f
C317 B.n277 VSUBS 0.008148f
C318 B.n278 VSUBS 0.008148f
C319 B.n279 VSUBS 0.008148f
C320 B.n280 VSUBS 0.008148f
C321 B.n281 VSUBS 0.008148f
C322 B.n282 VSUBS 0.008148f
C323 B.n283 VSUBS 0.008148f
C324 B.n284 VSUBS 0.008148f
C325 B.n285 VSUBS 0.008148f
C326 B.n286 VSUBS 0.008148f
C327 B.n287 VSUBS 0.008148f
C328 B.n288 VSUBS 0.008148f
C329 B.n289 VSUBS 0.005632f
C330 B.n290 VSUBS 0.008148f
C331 B.n291 VSUBS 0.008148f
C332 B.n292 VSUBS 0.006591f
C333 B.n293 VSUBS 0.008148f
C334 B.n294 VSUBS 0.008148f
C335 B.n295 VSUBS 0.008148f
C336 B.n296 VSUBS 0.008148f
C337 B.n297 VSUBS 0.008148f
C338 B.n298 VSUBS 0.008148f
C339 B.n299 VSUBS 0.008148f
C340 B.n300 VSUBS 0.008148f
C341 B.n301 VSUBS 0.008148f
C342 B.n302 VSUBS 0.008148f
C343 B.n303 VSUBS 0.008148f
C344 B.n304 VSUBS 0.006591f
C345 B.n305 VSUBS 0.018879f
C346 B.n306 VSUBS 0.005632f
C347 B.n307 VSUBS 0.008148f
C348 B.n308 VSUBS 0.008148f
C349 B.n309 VSUBS 0.008148f
C350 B.n310 VSUBS 0.008148f
C351 B.n311 VSUBS 0.008148f
C352 B.n312 VSUBS 0.008148f
C353 B.n313 VSUBS 0.008148f
C354 B.n314 VSUBS 0.008148f
C355 B.n315 VSUBS 0.008148f
C356 B.n316 VSUBS 0.008148f
C357 B.n317 VSUBS 0.008148f
C358 B.n318 VSUBS 0.008148f
C359 B.n319 VSUBS 0.008148f
C360 B.n320 VSUBS 0.008148f
C361 B.n321 VSUBS 0.008148f
C362 B.n322 VSUBS 0.008148f
C363 B.n323 VSUBS 0.008148f
C364 B.n324 VSUBS 0.008148f
C365 B.n325 VSUBS 0.019253f
C366 B.n326 VSUBS 0.019253f
C367 B.n327 VSUBS 0.018612f
C368 B.n328 VSUBS 0.008148f
C369 B.n329 VSUBS 0.008148f
C370 B.n330 VSUBS 0.008148f
C371 B.n331 VSUBS 0.008148f
C372 B.n332 VSUBS 0.008148f
C373 B.n333 VSUBS 0.008148f
C374 B.n334 VSUBS 0.008148f
C375 B.n335 VSUBS 0.008148f
C376 B.n336 VSUBS 0.008148f
C377 B.n337 VSUBS 0.008148f
C378 B.n338 VSUBS 0.008148f
C379 B.n339 VSUBS 0.008148f
C380 B.n340 VSUBS 0.008148f
C381 B.n341 VSUBS 0.008148f
C382 B.n342 VSUBS 0.008148f
C383 B.n343 VSUBS 0.008148f
C384 B.n344 VSUBS 0.008148f
C385 B.n345 VSUBS 0.008148f
C386 B.n346 VSUBS 0.008148f
C387 B.n347 VSUBS 0.008148f
C388 B.n348 VSUBS 0.008148f
C389 B.n349 VSUBS 0.008148f
C390 B.n350 VSUBS 0.008148f
C391 B.n351 VSUBS 0.008148f
C392 B.n352 VSUBS 0.008148f
C393 B.n353 VSUBS 0.008148f
C394 B.n354 VSUBS 0.008148f
C395 B.n355 VSUBS 0.008148f
C396 B.n356 VSUBS 0.008148f
C397 B.n357 VSUBS 0.008148f
C398 B.n358 VSUBS 0.008148f
C399 B.n359 VSUBS 0.008148f
C400 B.n360 VSUBS 0.008148f
C401 B.n361 VSUBS 0.008148f
C402 B.n362 VSUBS 0.008148f
C403 B.n363 VSUBS 0.010633f
C404 B.n364 VSUBS 0.011327f
C405 B.n365 VSUBS 0.022525f
C406 VDD2.n0 VSUBS 0.019978f
C407 VDD2.n1 VSUBS 0.134228f
C408 VDD2.n2 VSUBS 0.010041f
C409 VDD2.t7 VSUBS 0.053449f
C410 VDD2.n3 VSUBS 0.062862f
C411 VDD2.n4 VSUBS 0.013994f
C412 VDD2.n5 VSUBS 0.0178f
C413 VDD2.n6 VSUBS 0.055569f
C414 VDD2.n7 VSUBS 0.010631f
C415 VDD2.n8 VSUBS 0.010041f
C416 VDD2.n9 VSUBS 0.046764f
C417 VDD2.n10 VSUBS 0.042276f
C418 VDD2.t3 VSUBS 0.037505f
C419 VDD2.t9 VSUBS 0.037505f
C420 VDD2.n11 VSUBS 0.18387f
C421 VDD2.n12 VSUBS 0.371034f
C422 VDD2.t5 VSUBS 0.037505f
C423 VDD2.t0 VSUBS 0.037505f
C424 VDD2.n13 VSUBS 0.185043f
C425 VDD2.n14 VSUBS 1.05695f
C426 VDD2.n15 VSUBS 0.019978f
C427 VDD2.n16 VSUBS 0.134228f
C428 VDD2.n17 VSUBS 0.010041f
C429 VDD2.t6 VSUBS 0.053449f
C430 VDD2.n18 VSUBS 0.062862f
C431 VDD2.n19 VSUBS 0.013994f
C432 VDD2.n20 VSUBS 0.0178f
C433 VDD2.n21 VSUBS 0.055569f
C434 VDD2.n22 VSUBS 0.010631f
C435 VDD2.n23 VSUBS 0.010041f
C436 VDD2.n24 VSUBS 0.046764f
C437 VDD2.n25 VSUBS 0.040844f
C438 VDD2.n26 VSUBS 1.0294f
C439 VDD2.t2 VSUBS 0.037505f
C440 VDD2.t1 VSUBS 0.037505f
C441 VDD2.n27 VSUBS 0.183871f
C442 VDD2.n28 VSUBS 0.28763f
C443 VDD2.t8 VSUBS 0.037505f
C444 VDD2.t4 VSUBS 0.037505f
C445 VDD2.n29 VSUBS 0.185034f
C446 VN.n0 VSUBS 0.078509f
C447 VN.t6 VSUBS 0.236117f
C448 VN.n1 VSUBS 0.159627f
C449 VN.t2 VSUBS 0.258154f
C450 VN.n2 VSUBS 0.128359f
C451 VN.n3 VSUBS 0.250773f
C452 VN.t0 VSUBS 0.236117f
C453 VN.n4 VSUBS 0.159627f
C454 VN.t4 VSUBS 0.236117f
C455 VN.n5 VSUBS 0.159627f
C456 VN.t9 VSUBS 0.236117f
C457 VN.n6 VSUBS 0.148932f
C458 VN.n7 VSUBS 0.052288f
C459 VN.n8 VSUBS 0.078509f
C460 VN.t1 VSUBS 0.236117f
C461 VN.n9 VSUBS 0.159627f
C462 VN.t8 VSUBS 0.236117f
C463 VN.t5 VSUBS 0.258154f
C464 VN.n10 VSUBS 0.128359f
C465 VN.n11 VSUBS 0.250773f
C466 VN.n12 VSUBS 0.159627f
C467 VN.t7 VSUBS 0.236117f
C468 VN.n13 VSUBS 0.159627f
C469 VN.t3 VSUBS 0.236117f
C470 VN.n14 VSUBS 0.148932f
C471 VN.n15 VSUBS 1.48613f
C472 VDD1.n0 VSUBS 0.019325f
C473 VDD1.n1 VSUBS 0.129839f
C474 VDD1.n2 VSUBS 0.009712f
C475 VDD1.t6 VSUBS 0.051701f
C476 VDD1.n3 VSUBS 0.060806f
C477 VDD1.n4 VSUBS 0.013536f
C478 VDD1.n5 VSUBS 0.017218f
C479 VDD1.n6 VSUBS 0.053753f
C480 VDD1.n7 VSUBS 0.010284f
C481 VDD1.n8 VSUBS 0.009712f
C482 VDD1.n9 VSUBS 0.045235f
C483 VDD1.n10 VSUBS 0.040894f
C484 VDD1.t0 VSUBS 0.036279f
C485 VDD1.t2 VSUBS 0.036279f
C486 VDD1.n11 VSUBS 0.177859f
C487 VDD1.n12 VSUBS 0.362825f
C488 VDD1.n13 VSUBS 0.019325f
C489 VDD1.n14 VSUBS 0.129839f
C490 VDD1.n15 VSUBS 0.009712f
C491 VDD1.t1 VSUBS 0.051701f
C492 VDD1.n16 VSUBS 0.060806f
C493 VDD1.n17 VSUBS 0.013536f
C494 VDD1.n18 VSUBS 0.017218f
C495 VDD1.n19 VSUBS 0.053753f
C496 VDD1.n20 VSUBS 0.010284f
C497 VDD1.n21 VSUBS 0.009712f
C498 VDD1.n22 VSUBS 0.045235f
C499 VDD1.n23 VSUBS 0.040894f
C500 VDD1.t3 VSUBS 0.036279f
C501 VDD1.t8 VSUBS 0.036279f
C502 VDD1.n24 VSUBS 0.177858f
C503 VDD1.n25 VSUBS 0.358902f
C504 VDD1.t4 VSUBS 0.036279f
C505 VDD1.t7 VSUBS 0.036279f
C506 VDD1.n26 VSUBS 0.178993f
C507 VDD1.n27 VSUBS 1.07409f
C508 VDD1.t5 VSUBS 0.036279f
C509 VDD1.t9 VSUBS 0.036279f
C510 VDD1.n28 VSUBS 0.177858f
C511 VDD1.n29 VSUBS 1.22815f
C512 VTAIL.t1 VSUBS 0.044914f
C513 VTAIL.t6 VSUBS 0.044914f
C514 VTAIL.n0 VSUBS 0.18873f
C515 VTAIL.n1 VSUBS 0.37937f
C516 VTAIL.n2 VSUBS 0.023924f
C517 VTAIL.n3 VSUBS 0.160743f
C518 VTAIL.n4 VSUBS 0.012024f
C519 VTAIL.t9 VSUBS 0.064007f
C520 VTAIL.n5 VSUBS 0.075279f
C521 VTAIL.n6 VSUBS 0.016758f
C522 VTAIL.n7 VSUBS 0.021316f
C523 VTAIL.n8 VSUBS 0.066546f
C524 VTAIL.n9 VSUBS 0.012731f
C525 VTAIL.n10 VSUBS 0.012024f
C526 VTAIL.n11 VSUBS 0.056002f
C527 VTAIL.n12 VSUBS 0.033492f
C528 VTAIL.n13 VSUBS 0.146778f
C529 VTAIL.t13 VSUBS 0.044914f
C530 VTAIL.t18 VSUBS 0.044914f
C531 VTAIL.n14 VSUBS 0.18873f
C532 VTAIL.n15 VSUBS 0.386984f
C533 VTAIL.t14 VSUBS 0.044914f
C534 VTAIL.t11 VSUBS 0.044914f
C535 VTAIL.n16 VSUBS 0.18873f
C536 VTAIL.n17 VSUBS 0.909735f
C537 VTAIL.t8 VSUBS 0.044914f
C538 VTAIL.t2 VSUBS 0.044914f
C539 VTAIL.n18 VSUBS 0.188731f
C540 VTAIL.n19 VSUBS 0.909734f
C541 VTAIL.t3 VSUBS 0.044914f
C542 VTAIL.t19 VSUBS 0.044914f
C543 VTAIL.n20 VSUBS 0.188731f
C544 VTAIL.n21 VSUBS 0.386983f
C545 VTAIL.n22 VSUBS 0.023924f
C546 VTAIL.n23 VSUBS 0.160743f
C547 VTAIL.n24 VSUBS 0.012024f
C548 VTAIL.t4 VSUBS 0.064007f
C549 VTAIL.n25 VSUBS 0.075279f
C550 VTAIL.n26 VSUBS 0.016758f
C551 VTAIL.n27 VSUBS 0.021316f
C552 VTAIL.n28 VSUBS 0.066546f
C553 VTAIL.n29 VSUBS 0.012731f
C554 VTAIL.n30 VSUBS 0.012024f
C555 VTAIL.n31 VSUBS 0.056002f
C556 VTAIL.n32 VSUBS 0.033492f
C557 VTAIL.n33 VSUBS 0.146778f
C558 VTAIL.t17 VSUBS 0.044914f
C559 VTAIL.t12 VSUBS 0.044914f
C560 VTAIL.n34 VSUBS 0.188731f
C561 VTAIL.n35 VSUBS 0.390401f
C562 VTAIL.t10 VSUBS 0.044914f
C563 VTAIL.t16 VSUBS 0.044914f
C564 VTAIL.n36 VSUBS 0.188731f
C565 VTAIL.n37 VSUBS 0.386983f
C566 VTAIL.n38 VSUBS 0.023924f
C567 VTAIL.n39 VSUBS 0.160743f
C568 VTAIL.n40 VSUBS 0.012024f
C569 VTAIL.t15 VSUBS 0.064007f
C570 VTAIL.n41 VSUBS 0.075279f
C571 VTAIL.n42 VSUBS 0.016758f
C572 VTAIL.n43 VSUBS 0.021316f
C573 VTAIL.n44 VSUBS 0.066546f
C574 VTAIL.n45 VSUBS 0.012731f
C575 VTAIL.n46 VSUBS 0.012024f
C576 VTAIL.n47 VSUBS 0.056002f
C577 VTAIL.n48 VSUBS 0.033492f
C578 VTAIL.n49 VSUBS 0.605196f
C579 VTAIL.n50 VSUBS 0.023924f
C580 VTAIL.n51 VSUBS 0.160743f
C581 VTAIL.n52 VSUBS 0.012024f
C582 VTAIL.t5 VSUBS 0.064007f
C583 VTAIL.n53 VSUBS 0.075279f
C584 VTAIL.n54 VSUBS 0.016758f
C585 VTAIL.n55 VSUBS 0.021316f
C586 VTAIL.n56 VSUBS 0.066546f
C587 VTAIL.n57 VSUBS 0.012731f
C588 VTAIL.n58 VSUBS 0.012024f
C589 VTAIL.n59 VSUBS 0.056002f
C590 VTAIL.n60 VSUBS 0.033492f
C591 VTAIL.n61 VSUBS 0.605196f
C592 VTAIL.t0 VSUBS 0.044914f
C593 VTAIL.t7 VSUBS 0.044914f
C594 VTAIL.n62 VSUBS 0.18873f
C595 VTAIL.n63 VSUBS 0.337103f
C596 VP.n0 VSUBS 0.082325f
C597 VP.t6 VSUBS 0.247596f
C598 VP.n1 VSUBS 0.167388f
C599 VP.n2 VSUBS 0.082325f
C600 VP.t0 VSUBS 0.247596f
C601 VP.t4 VSUBS 0.247596f
C602 VP.t7 VSUBS 0.247596f
C603 VP.n3 VSUBS 0.262965f
C604 VP.t9 VSUBS 0.247596f
C605 VP.t3 VSUBS 0.270705f
C606 VP.n4 VSUBS 0.134599f
C607 VP.n5 VSUBS 0.167388f
C608 VP.n6 VSUBS 0.167388f
C609 VP.n7 VSUBS 0.167388f
C610 VP.n8 VSUBS 0.156172f
C611 VP.n9 VSUBS 1.52555f
C612 VP.t8 VSUBS 0.247596f
C613 VP.n10 VSUBS 0.156172f
C614 VP.n11 VSUBS 1.57582f
C615 VP.n12 VSUBS 0.082325f
C616 VP.n13 VSUBS 0.098852f
C617 VP.t1 VSUBS 0.247596f
C618 VP.n14 VSUBS 0.167388f
C619 VP.t5 VSUBS 0.247596f
C620 VP.n15 VSUBS 0.167388f
C621 VP.t2 VSUBS 0.247596f
C622 VP.n16 VSUBS 0.156172f
C623 VP.n17 VSUBS 0.05483f
.ends

