* NGSPICE file created from diff_pair_sample_1048.ext - technology: sky130A

.subckt diff_pair_sample_1048 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t15 VN.t0 VDD2.t0 B.t3 sky130_fd_pr__nfet_01v8 ad=0.3705 pd=2.68 as=0.15675 ps=1.28 w=0.95 l=2.71
X1 VDD1.t7 VP.t0 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=0.15675 pd=1.28 as=0.15675 ps=1.28 w=0.95 l=2.71
X2 VDD1.t6 VP.t1 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=0.15675 pd=1.28 as=0.3705 ps=2.68 w=0.95 l=2.71
X3 VTAIL.t14 VN.t1 VDD2.t6 B.t6 sky130_fd_pr__nfet_01v8 ad=0.15675 pd=1.28 as=0.15675 ps=1.28 w=0.95 l=2.71
X4 VDD2.t4 VN.t2 VTAIL.t13 B.t2 sky130_fd_pr__nfet_01v8 ad=0.15675 pd=1.28 as=0.3705 ps=2.68 w=0.95 l=2.71
X5 B.t21 B.t19 B.t20 B.t16 sky130_fd_pr__nfet_01v8 ad=0.3705 pd=2.68 as=0 ps=0 w=0.95 l=2.71
X6 VTAIL.t3 VP.t2 VDD1.t5 B.t3 sky130_fd_pr__nfet_01v8 ad=0.3705 pd=2.68 as=0.15675 ps=1.28 w=0.95 l=2.71
X7 B.t18 B.t15 B.t17 B.t16 sky130_fd_pr__nfet_01v8 ad=0.3705 pd=2.68 as=0 ps=0 w=0.95 l=2.71
X8 VTAIL.t12 VN.t3 VDD2.t2 B.t4 sky130_fd_pr__nfet_01v8 ad=0.15675 pd=1.28 as=0.15675 ps=1.28 w=0.95 l=2.71
X9 VTAIL.t4 VP.t3 VDD1.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=0.15675 pd=1.28 as=0.15675 ps=1.28 w=0.95 l=2.71
X10 VTAIL.t11 VN.t4 VDD2.t5 B.t0 sky130_fd_pr__nfet_01v8 ad=0.3705 pd=2.68 as=0.15675 ps=1.28 w=0.95 l=2.71
X11 VTAIL.t6 VP.t4 VDD1.t3 B.t6 sky130_fd_pr__nfet_01v8 ad=0.15675 pd=1.28 as=0.15675 ps=1.28 w=0.95 l=2.71
X12 VDD2.t7 VN.t5 VTAIL.t10 B.t7 sky130_fd_pr__nfet_01v8 ad=0.15675 pd=1.28 as=0.3705 ps=2.68 w=0.95 l=2.71
X13 B.t14 B.t12 B.t13 B.t9 sky130_fd_pr__nfet_01v8 ad=0.3705 pd=2.68 as=0 ps=0 w=0.95 l=2.71
X14 VTAIL.t0 VP.t5 VDD1.t2 B.t0 sky130_fd_pr__nfet_01v8 ad=0.3705 pd=2.68 as=0.15675 ps=1.28 w=0.95 l=2.71
X15 VDD1.t1 VP.t6 VTAIL.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=0.15675 pd=1.28 as=0.15675 ps=1.28 w=0.95 l=2.71
X16 VDD1.t0 VP.t7 VTAIL.t7 B.t7 sky130_fd_pr__nfet_01v8 ad=0.15675 pd=1.28 as=0.3705 ps=2.68 w=0.95 l=2.71
X17 VDD2.t1 VN.t6 VTAIL.t9 B.t5 sky130_fd_pr__nfet_01v8 ad=0.15675 pd=1.28 as=0.15675 ps=1.28 w=0.95 l=2.71
X18 VDD2.t3 VN.t7 VTAIL.t8 B.t1 sky130_fd_pr__nfet_01v8 ad=0.15675 pd=1.28 as=0.15675 ps=1.28 w=0.95 l=2.71
X19 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=0.3705 pd=2.68 as=0 ps=0 w=0.95 l=2.71
R0 VN.n59 VN.n31 161.3
R1 VN.n58 VN.n57 161.3
R2 VN.n56 VN.n32 161.3
R3 VN.n55 VN.n54 161.3
R4 VN.n53 VN.n33 161.3
R5 VN.n52 VN.n51 161.3
R6 VN.n50 VN.n49 161.3
R7 VN.n48 VN.n35 161.3
R8 VN.n47 VN.n46 161.3
R9 VN.n45 VN.n36 161.3
R10 VN.n44 VN.n43 161.3
R11 VN.n42 VN.n37 161.3
R12 VN.n41 VN.n40 161.3
R13 VN.n28 VN.n0 161.3
R14 VN.n27 VN.n26 161.3
R15 VN.n25 VN.n1 161.3
R16 VN.n24 VN.n23 161.3
R17 VN.n22 VN.n2 161.3
R18 VN.n21 VN.n20 161.3
R19 VN.n19 VN.n18 161.3
R20 VN.n17 VN.n4 161.3
R21 VN.n16 VN.n15 161.3
R22 VN.n14 VN.n5 161.3
R23 VN.n13 VN.n12 161.3
R24 VN.n11 VN.n6 161.3
R25 VN.n10 VN.n9 161.3
R26 VN.n30 VN.n29 107.82
R27 VN.n61 VN.n60 107.82
R28 VN.n8 VN.n7 72.3368
R29 VN.n39 VN.n38 72.3368
R30 VN.n23 VN.n1 44.3785
R31 VN.n54 VN.n32 44.3785
R32 VN VN.n61 43.2557
R33 VN.n12 VN.n5 40.4934
R34 VN.n16 VN.n5 40.4934
R35 VN.n43 VN.n36 40.4934
R36 VN.n47 VN.n36 40.4934
R37 VN.n8 VN.t0 39.5494
R38 VN.n39 VN.t5 39.5494
R39 VN.n23 VN.n22 36.6083
R40 VN.n54 VN.n53 36.6083
R41 VN.n11 VN.n10 24.4675
R42 VN.n12 VN.n11 24.4675
R43 VN.n17 VN.n16 24.4675
R44 VN.n18 VN.n17 24.4675
R45 VN.n22 VN.n21 24.4675
R46 VN.n27 VN.n1 24.4675
R47 VN.n28 VN.n27 24.4675
R48 VN.n43 VN.n42 24.4675
R49 VN.n42 VN.n41 24.4675
R50 VN.n53 VN.n52 24.4675
R51 VN.n49 VN.n48 24.4675
R52 VN.n48 VN.n47 24.4675
R53 VN.n59 VN.n58 24.4675
R54 VN.n58 VN.n32 24.4675
R55 VN.n21 VN.n3 23.4888
R56 VN.n52 VN.n34 23.4888
R57 VN.n7 VN.t6 8.44884
R58 VN.n3 VN.t3 8.44884
R59 VN.n29 VN.t2 8.44884
R60 VN.n38 VN.t1 8.44884
R61 VN.n34 VN.t7 8.44884
R62 VN.n60 VN.t4 8.44884
R63 VN.n40 VN.n39 7.30997
R64 VN.n9 VN.n8 7.30997
R65 VN.n29 VN.n28 2.93654
R66 VN.n60 VN.n59 2.93654
R67 VN.n10 VN.n7 0.97918
R68 VN.n18 VN.n3 0.97918
R69 VN.n41 VN.n38 0.97918
R70 VN.n49 VN.n34 0.97918
R71 VN.n61 VN.n31 0.278367
R72 VN.n30 VN.n0 0.278367
R73 VN.n57 VN.n31 0.189894
R74 VN.n57 VN.n56 0.189894
R75 VN.n56 VN.n55 0.189894
R76 VN.n55 VN.n33 0.189894
R77 VN.n51 VN.n33 0.189894
R78 VN.n51 VN.n50 0.189894
R79 VN.n50 VN.n35 0.189894
R80 VN.n46 VN.n35 0.189894
R81 VN.n46 VN.n45 0.189894
R82 VN.n45 VN.n44 0.189894
R83 VN.n44 VN.n37 0.189894
R84 VN.n40 VN.n37 0.189894
R85 VN.n9 VN.n6 0.189894
R86 VN.n13 VN.n6 0.189894
R87 VN.n14 VN.n13 0.189894
R88 VN.n15 VN.n14 0.189894
R89 VN.n15 VN.n4 0.189894
R90 VN.n19 VN.n4 0.189894
R91 VN.n20 VN.n19 0.189894
R92 VN.n20 VN.n2 0.189894
R93 VN.n24 VN.n2 0.189894
R94 VN.n25 VN.n24 0.189894
R95 VN.n26 VN.n25 0.189894
R96 VN.n26 VN.n0 0.189894
R97 VN VN.n30 0.153454
R98 VDD2.n2 VDD2.n1 240.417
R99 VDD2.n2 VDD2.n0 240.417
R100 VDD2 VDD2.n5 240.416
R101 VDD2.n4 VDD2.n3 239.163
R102 VDD2.n4 VDD2.n2 36.3274
R103 VDD2.n5 VDD2.t6 20.8426
R104 VDD2.n5 VDD2.t7 20.8426
R105 VDD2.n3 VDD2.t5 20.8426
R106 VDD2.n3 VDD2.t3 20.8426
R107 VDD2.n1 VDD2.t2 20.8426
R108 VDD2.n1 VDD2.t4 20.8426
R109 VDD2.n0 VDD2.t0 20.8426
R110 VDD2.n0 VDD2.t1 20.8426
R111 VDD2 VDD2.n4 1.36903
R112 VTAIL.n14 VTAIL.t2 243.327
R113 VTAIL.n11 VTAIL.t3 243.327
R114 VTAIL.n10 VTAIL.t10 243.327
R115 VTAIL.n7 VTAIL.t11 243.327
R116 VTAIL.n15 VTAIL.t13 243.326
R117 VTAIL.n2 VTAIL.t15 243.326
R118 VTAIL.n3 VTAIL.t7 243.326
R119 VTAIL.n6 VTAIL.t0 243.326
R120 VTAIL.n13 VTAIL.n12 222.484
R121 VTAIL.n9 VTAIL.n8 222.484
R122 VTAIL.n1 VTAIL.n0 222.483
R123 VTAIL.n5 VTAIL.n4 222.483
R124 VTAIL.n0 VTAIL.t9 20.8426
R125 VTAIL.n0 VTAIL.t12 20.8426
R126 VTAIL.n4 VTAIL.t1 20.8426
R127 VTAIL.n4 VTAIL.t6 20.8426
R128 VTAIL.n12 VTAIL.t5 20.8426
R129 VTAIL.n12 VTAIL.t4 20.8426
R130 VTAIL.n8 VTAIL.t8 20.8426
R131 VTAIL.n8 VTAIL.t14 20.8426
R132 VTAIL.n15 VTAIL.n14 15.8065
R133 VTAIL.n7 VTAIL.n6 15.8065
R134 VTAIL.n9 VTAIL.n7 2.62119
R135 VTAIL.n10 VTAIL.n9 2.62119
R136 VTAIL.n13 VTAIL.n11 2.62119
R137 VTAIL.n14 VTAIL.n13 2.62119
R138 VTAIL.n6 VTAIL.n5 2.62119
R139 VTAIL.n5 VTAIL.n3 2.62119
R140 VTAIL.n2 VTAIL.n1 2.62119
R141 VTAIL VTAIL.n15 2.563
R142 VTAIL.n11 VTAIL.n10 0.470328
R143 VTAIL.n3 VTAIL.n2 0.470328
R144 VTAIL VTAIL.n1 0.0586897
R145 B.n577 B.n576 585
R146 B.n170 B.n111 585
R147 B.n169 B.n168 585
R148 B.n167 B.n166 585
R149 B.n165 B.n164 585
R150 B.n163 B.n162 585
R151 B.n161 B.n160 585
R152 B.n159 B.n158 585
R153 B.n157 B.n156 585
R154 B.n154 B.n153 585
R155 B.n152 B.n151 585
R156 B.n150 B.n149 585
R157 B.n148 B.n147 585
R158 B.n146 B.n145 585
R159 B.n144 B.n143 585
R160 B.n142 B.n141 585
R161 B.n140 B.n139 585
R162 B.n138 B.n137 585
R163 B.n136 B.n135 585
R164 B.n133 B.n132 585
R165 B.n131 B.n130 585
R166 B.n129 B.n128 585
R167 B.n127 B.n126 585
R168 B.n125 B.n124 585
R169 B.n123 B.n122 585
R170 B.n121 B.n120 585
R171 B.n119 B.n118 585
R172 B.n117 B.n116 585
R173 B.n575 B.n97 585
R174 B.n580 B.n97 585
R175 B.n574 B.n96 585
R176 B.n581 B.n96 585
R177 B.n573 B.n572 585
R178 B.n572 B.n92 585
R179 B.n571 B.n91 585
R180 B.n587 B.n91 585
R181 B.n570 B.n90 585
R182 B.n588 B.n90 585
R183 B.n569 B.n89 585
R184 B.n589 B.n89 585
R185 B.n568 B.n567 585
R186 B.n567 B.n85 585
R187 B.n566 B.n84 585
R188 B.n595 B.n84 585
R189 B.n565 B.n83 585
R190 B.n596 B.n83 585
R191 B.n564 B.n82 585
R192 B.n597 B.n82 585
R193 B.n563 B.n562 585
R194 B.n562 B.n78 585
R195 B.n561 B.n77 585
R196 B.n603 B.n77 585
R197 B.n560 B.n76 585
R198 B.n604 B.n76 585
R199 B.n559 B.n75 585
R200 B.n605 B.n75 585
R201 B.n558 B.n557 585
R202 B.n557 B.n71 585
R203 B.n556 B.n70 585
R204 B.n611 B.n70 585
R205 B.n555 B.n69 585
R206 B.n612 B.n69 585
R207 B.n554 B.n68 585
R208 B.n613 B.n68 585
R209 B.n553 B.n552 585
R210 B.n552 B.n64 585
R211 B.n551 B.n63 585
R212 B.n619 B.n63 585
R213 B.n550 B.n62 585
R214 B.n620 B.n62 585
R215 B.n549 B.n61 585
R216 B.n621 B.n61 585
R217 B.n548 B.n547 585
R218 B.n547 B.n57 585
R219 B.n546 B.n56 585
R220 B.n627 B.n56 585
R221 B.n545 B.n55 585
R222 B.n628 B.n55 585
R223 B.n544 B.n54 585
R224 B.n629 B.n54 585
R225 B.n543 B.n542 585
R226 B.n542 B.n50 585
R227 B.n541 B.n49 585
R228 B.n635 B.n49 585
R229 B.n540 B.n48 585
R230 B.n636 B.n48 585
R231 B.n539 B.n47 585
R232 B.n637 B.n47 585
R233 B.n538 B.n537 585
R234 B.n537 B.n43 585
R235 B.n536 B.n42 585
R236 B.n643 B.n42 585
R237 B.n535 B.n41 585
R238 B.n644 B.n41 585
R239 B.n534 B.n40 585
R240 B.n645 B.n40 585
R241 B.n533 B.n532 585
R242 B.n532 B.n36 585
R243 B.n531 B.n35 585
R244 B.n651 B.n35 585
R245 B.n530 B.n34 585
R246 B.n652 B.n34 585
R247 B.n529 B.n33 585
R248 B.n653 B.n33 585
R249 B.n528 B.n527 585
R250 B.n527 B.n29 585
R251 B.n526 B.n28 585
R252 B.n659 B.n28 585
R253 B.n525 B.n27 585
R254 B.n660 B.n27 585
R255 B.n524 B.n26 585
R256 B.n661 B.n26 585
R257 B.n523 B.n522 585
R258 B.n522 B.n22 585
R259 B.n521 B.n21 585
R260 B.n667 B.n21 585
R261 B.n520 B.n20 585
R262 B.n668 B.n20 585
R263 B.n519 B.n19 585
R264 B.n669 B.n19 585
R265 B.n518 B.n517 585
R266 B.n517 B.n18 585
R267 B.n516 B.n14 585
R268 B.n675 B.n14 585
R269 B.n515 B.n13 585
R270 B.n676 B.n13 585
R271 B.n514 B.n12 585
R272 B.n677 B.n12 585
R273 B.n513 B.n512 585
R274 B.n512 B.n8 585
R275 B.n511 B.n7 585
R276 B.n683 B.n7 585
R277 B.n510 B.n6 585
R278 B.n684 B.n6 585
R279 B.n509 B.n5 585
R280 B.n685 B.n5 585
R281 B.n508 B.n507 585
R282 B.n507 B.n4 585
R283 B.n506 B.n171 585
R284 B.n506 B.n505 585
R285 B.n496 B.n172 585
R286 B.n173 B.n172 585
R287 B.n498 B.n497 585
R288 B.n499 B.n498 585
R289 B.n495 B.n178 585
R290 B.n178 B.n177 585
R291 B.n494 B.n493 585
R292 B.n493 B.n492 585
R293 B.n180 B.n179 585
R294 B.n485 B.n180 585
R295 B.n484 B.n483 585
R296 B.n486 B.n484 585
R297 B.n482 B.n185 585
R298 B.n185 B.n184 585
R299 B.n481 B.n480 585
R300 B.n480 B.n479 585
R301 B.n187 B.n186 585
R302 B.n188 B.n187 585
R303 B.n472 B.n471 585
R304 B.n473 B.n472 585
R305 B.n470 B.n193 585
R306 B.n193 B.n192 585
R307 B.n469 B.n468 585
R308 B.n468 B.n467 585
R309 B.n195 B.n194 585
R310 B.n196 B.n195 585
R311 B.n460 B.n459 585
R312 B.n461 B.n460 585
R313 B.n458 B.n201 585
R314 B.n201 B.n200 585
R315 B.n457 B.n456 585
R316 B.n456 B.n455 585
R317 B.n203 B.n202 585
R318 B.n204 B.n203 585
R319 B.n448 B.n447 585
R320 B.n449 B.n448 585
R321 B.n446 B.n209 585
R322 B.n209 B.n208 585
R323 B.n445 B.n444 585
R324 B.n444 B.n443 585
R325 B.n211 B.n210 585
R326 B.n212 B.n211 585
R327 B.n436 B.n435 585
R328 B.n437 B.n436 585
R329 B.n434 B.n217 585
R330 B.n217 B.n216 585
R331 B.n433 B.n432 585
R332 B.n432 B.n431 585
R333 B.n219 B.n218 585
R334 B.n220 B.n219 585
R335 B.n424 B.n423 585
R336 B.n425 B.n424 585
R337 B.n422 B.n225 585
R338 B.n225 B.n224 585
R339 B.n421 B.n420 585
R340 B.n420 B.n419 585
R341 B.n227 B.n226 585
R342 B.n228 B.n227 585
R343 B.n412 B.n411 585
R344 B.n413 B.n412 585
R345 B.n410 B.n232 585
R346 B.n236 B.n232 585
R347 B.n409 B.n408 585
R348 B.n408 B.n407 585
R349 B.n234 B.n233 585
R350 B.n235 B.n234 585
R351 B.n400 B.n399 585
R352 B.n401 B.n400 585
R353 B.n398 B.n241 585
R354 B.n241 B.n240 585
R355 B.n397 B.n396 585
R356 B.n396 B.n395 585
R357 B.n243 B.n242 585
R358 B.n244 B.n243 585
R359 B.n388 B.n387 585
R360 B.n389 B.n388 585
R361 B.n386 B.n249 585
R362 B.n249 B.n248 585
R363 B.n385 B.n384 585
R364 B.n384 B.n383 585
R365 B.n251 B.n250 585
R366 B.n252 B.n251 585
R367 B.n376 B.n375 585
R368 B.n377 B.n376 585
R369 B.n374 B.n257 585
R370 B.n257 B.n256 585
R371 B.n373 B.n372 585
R372 B.n372 B.n371 585
R373 B.n259 B.n258 585
R374 B.n260 B.n259 585
R375 B.n364 B.n363 585
R376 B.n365 B.n364 585
R377 B.n362 B.n265 585
R378 B.n265 B.n264 585
R379 B.n361 B.n360 585
R380 B.n360 B.n359 585
R381 B.n267 B.n266 585
R382 B.n268 B.n267 585
R383 B.n352 B.n351 585
R384 B.n353 B.n352 585
R385 B.n350 B.n273 585
R386 B.n273 B.n272 585
R387 B.n345 B.n344 585
R388 B.n343 B.n289 585
R389 B.n342 B.n288 585
R390 B.n347 B.n288 585
R391 B.n341 B.n340 585
R392 B.n339 B.n338 585
R393 B.n337 B.n336 585
R394 B.n335 B.n334 585
R395 B.n333 B.n332 585
R396 B.n331 B.n330 585
R397 B.n329 B.n328 585
R398 B.n327 B.n326 585
R399 B.n325 B.n324 585
R400 B.n323 B.n322 585
R401 B.n321 B.n320 585
R402 B.n319 B.n318 585
R403 B.n317 B.n316 585
R404 B.n315 B.n314 585
R405 B.n313 B.n312 585
R406 B.n311 B.n310 585
R407 B.n309 B.n308 585
R408 B.n307 B.n306 585
R409 B.n305 B.n304 585
R410 B.n303 B.n302 585
R411 B.n301 B.n300 585
R412 B.n299 B.n298 585
R413 B.n297 B.n296 585
R414 B.n275 B.n274 585
R415 B.n349 B.n348 585
R416 B.n348 B.n347 585
R417 B.n271 B.n270 585
R418 B.n272 B.n271 585
R419 B.n355 B.n354 585
R420 B.n354 B.n353 585
R421 B.n356 B.n269 585
R422 B.n269 B.n268 585
R423 B.n358 B.n357 585
R424 B.n359 B.n358 585
R425 B.n263 B.n262 585
R426 B.n264 B.n263 585
R427 B.n367 B.n366 585
R428 B.n366 B.n365 585
R429 B.n368 B.n261 585
R430 B.n261 B.n260 585
R431 B.n370 B.n369 585
R432 B.n371 B.n370 585
R433 B.n255 B.n254 585
R434 B.n256 B.n255 585
R435 B.n379 B.n378 585
R436 B.n378 B.n377 585
R437 B.n380 B.n253 585
R438 B.n253 B.n252 585
R439 B.n382 B.n381 585
R440 B.n383 B.n382 585
R441 B.n247 B.n246 585
R442 B.n248 B.n247 585
R443 B.n391 B.n390 585
R444 B.n390 B.n389 585
R445 B.n392 B.n245 585
R446 B.n245 B.n244 585
R447 B.n394 B.n393 585
R448 B.n395 B.n394 585
R449 B.n239 B.n238 585
R450 B.n240 B.n239 585
R451 B.n403 B.n402 585
R452 B.n402 B.n401 585
R453 B.n404 B.n237 585
R454 B.n237 B.n235 585
R455 B.n406 B.n405 585
R456 B.n407 B.n406 585
R457 B.n231 B.n230 585
R458 B.n236 B.n231 585
R459 B.n415 B.n414 585
R460 B.n414 B.n413 585
R461 B.n416 B.n229 585
R462 B.n229 B.n228 585
R463 B.n418 B.n417 585
R464 B.n419 B.n418 585
R465 B.n223 B.n222 585
R466 B.n224 B.n223 585
R467 B.n427 B.n426 585
R468 B.n426 B.n425 585
R469 B.n428 B.n221 585
R470 B.n221 B.n220 585
R471 B.n430 B.n429 585
R472 B.n431 B.n430 585
R473 B.n215 B.n214 585
R474 B.n216 B.n215 585
R475 B.n439 B.n438 585
R476 B.n438 B.n437 585
R477 B.n440 B.n213 585
R478 B.n213 B.n212 585
R479 B.n442 B.n441 585
R480 B.n443 B.n442 585
R481 B.n207 B.n206 585
R482 B.n208 B.n207 585
R483 B.n451 B.n450 585
R484 B.n450 B.n449 585
R485 B.n452 B.n205 585
R486 B.n205 B.n204 585
R487 B.n454 B.n453 585
R488 B.n455 B.n454 585
R489 B.n199 B.n198 585
R490 B.n200 B.n199 585
R491 B.n463 B.n462 585
R492 B.n462 B.n461 585
R493 B.n464 B.n197 585
R494 B.n197 B.n196 585
R495 B.n466 B.n465 585
R496 B.n467 B.n466 585
R497 B.n191 B.n190 585
R498 B.n192 B.n191 585
R499 B.n475 B.n474 585
R500 B.n474 B.n473 585
R501 B.n476 B.n189 585
R502 B.n189 B.n188 585
R503 B.n478 B.n477 585
R504 B.n479 B.n478 585
R505 B.n183 B.n182 585
R506 B.n184 B.n183 585
R507 B.n488 B.n487 585
R508 B.n487 B.n486 585
R509 B.n489 B.n181 585
R510 B.n485 B.n181 585
R511 B.n491 B.n490 585
R512 B.n492 B.n491 585
R513 B.n176 B.n175 585
R514 B.n177 B.n176 585
R515 B.n501 B.n500 585
R516 B.n500 B.n499 585
R517 B.n502 B.n174 585
R518 B.n174 B.n173 585
R519 B.n504 B.n503 585
R520 B.n505 B.n504 585
R521 B.n2 B.n0 585
R522 B.n4 B.n2 585
R523 B.n3 B.n1 585
R524 B.n684 B.n3 585
R525 B.n682 B.n681 585
R526 B.n683 B.n682 585
R527 B.n680 B.n9 585
R528 B.n9 B.n8 585
R529 B.n679 B.n678 585
R530 B.n678 B.n677 585
R531 B.n11 B.n10 585
R532 B.n676 B.n11 585
R533 B.n674 B.n673 585
R534 B.n675 B.n674 585
R535 B.n672 B.n15 585
R536 B.n18 B.n15 585
R537 B.n671 B.n670 585
R538 B.n670 B.n669 585
R539 B.n17 B.n16 585
R540 B.n668 B.n17 585
R541 B.n666 B.n665 585
R542 B.n667 B.n666 585
R543 B.n664 B.n23 585
R544 B.n23 B.n22 585
R545 B.n663 B.n662 585
R546 B.n662 B.n661 585
R547 B.n25 B.n24 585
R548 B.n660 B.n25 585
R549 B.n658 B.n657 585
R550 B.n659 B.n658 585
R551 B.n656 B.n30 585
R552 B.n30 B.n29 585
R553 B.n655 B.n654 585
R554 B.n654 B.n653 585
R555 B.n32 B.n31 585
R556 B.n652 B.n32 585
R557 B.n650 B.n649 585
R558 B.n651 B.n650 585
R559 B.n648 B.n37 585
R560 B.n37 B.n36 585
R561 B.n647 B.n646 585
R562 B.n646 B.n645 585
R563 B.n39 B.n38 585
R564 B.n644 B.n39 585
R565 B.n642 B.n641 585
R566 B.n643 B.n642 585
R567 B.n640 B.n44 585
R568 B.n44 B.n43 585
R569 B.n639 B.n638 585
R570 B.n638 B.n637 585
R571 B.n46 B.n45 585
R572 B.n636 B.n46 585
R573 B.n634 B.n633 585
R574 B.n635 B.n634 585
R575 B.n632 B.n51 585
R576 B.n51 B.n50 585
R577 B.n631 B.n630 585
R578 B.n630 B.n629 585
R579 B.n53 B.n52 585
R580 B.n628 B.n53 585
R581 B.n626 B.n625 585
R582 B.n627 B.n626 585
R583 B.n624 B.n58 585
R584 B.n58 B.n57 585
R585 B.n623 B.n622 585
R586 B.n622 B.n621 585
R587 B.n60 B.n59 585
R588 B.n620 B.n60 585
R589 B.n618 B.n617 585
R590 B.n619 B.n618 585
R591 B.n616 B.n65 585
R592 B.n65 B.n64 585
R593 B.n615 B.n614 585
R594 B.n614 B.n613 585
R595 B.n67 B.n66 585
R596 B.n612 B.n67 585
R597 B.n610 B.n609 585
R598 B.n611 B.n610 585
R599 B.n608 B.n72 585
R600 B.n72 B.n71 585
R601 B.n607 B.n606 585
R602 B.n606 B.n605 585
R603 B.n74 B.n73 585
R604 B.n604 B.n74 585
R605 B.n602 B.n601 585
R606 B.n603 B.n602 585
R607 B.n600 B.n79 585
R608 B.n79 B.n78 585
R609 B.n599 B.n598 585
R610 B.n598 B.n597 585
R611 B.n81 B.n80 585
R612 B.n596 B.n81 585
R613 B.n594 B.n593 585
R614 B.n595 B.n594 585
R615 B.n592 B.n86 585
R616 B.n86 B.n85 585
R617 B.n591 B.n590 585
R618 B.n590 B.n589 585
R619 B.n88 B.n87 585
R620 B.n588 B.n88 585
R621 B.n586 B.n585 585
R622 B.n587 B.n586 585
R623 B.n584 B.n93 585
R624 B.n93 B.n92 585
R625 B.n583 B.n582 585
R626 B.n582 B.n581 585
R627 B.n95 B.n94 585
R628 B.n580 B.n95 585
R629 B.n687 B.n686 585
R630 B.n686 B.n685 585
R631 B.n345 B.n271 454.062
R632 B.n116 B.n95 454.062
R633 B.n348 B.n273 454.062
R634 B.n577 B.n97 454.062
R635 B.n293 B.t21 292.921
R636 B.n290 B.t18 292.921
R637 B.n114 B.t10 292.921
R638 B.n112 B.t13 292.921
R639 B.n579 B.n578 256.663
R640 B.n579 B.n110 256.663
R641 B.n579 B.n109 256.663
R642 B.n579 B.n108 256.663
R643 B.n579 B.n107 256.663
R644 B.n579 B.n106 256.663
R645 B.n579 B.n105 256.663
R646 B.n579 B.n104 256.663
R647 B.n579 B.n103 256.663
R648 B.n579 B.n102 256.663
R649 B.n579 B.n101 256.663
R650 B.n579 B.n100 256.663
R651 B.n579 B.n99 256.663
R652 B.n579 B.n98 256.663
R653 B.n347 B.n346 256.663
R654 B.n347 B.n276 256.663
R655 B.n347 B.n277 256.663
R656 B.n347 B.n278 256.663
R657 B.n347 B.n279 256.663
R658 B.n347 B.n280 256.663
R659 B.n347 B.n281 256.663
R660 B.n347 B.n282 256.663
R661 B.n347 B.n283 256.663
R662 B.n347 B.n284 256.663
R663 B.n347 B.n285 256.663
R664 B.n347 B.n286 256.663
R665 B.n347 B.n287 256.663
R666 B.n294 B.t20 233.964
R667 B.n291 B.t17 233.964
R668 B.n115 B.t11 233.964
R669 B.n113 B.t14 233.964
R670 B.n293 B.t19 209.102
R671 B.n290 B.t15 209.102
R672 B.n114 B.t8 209.102
R673 B.n112 B.t12 209.102
R674 B.n347 B.n272 196.145
R675 B.n580 B.n579 196.145
R676 B.n354 B.n271 163.367
R677 B.n354 B.n269 163.367
R678 B.n358 B.n269 163.367
R679 B.n358 B.n263 163.367
R680 B.n366 B.n263 163.367
R681 B.n366 B.n261 163.367
R682 B.n370 B.n261 163.367
R683 B.n370 B.n255 163.367
R684 B.n378 B.n255 163.367
R685 B.n378 B.n253 163.367
R686 B.n382 B.n253 163.367
R687 B.n382 B.n247 163.367
R688 B.n390 B.n247 163.367
R689 B.n390 B.n245 163.367
R690 B.n394 B.n245 163.367
R691 B.n394 B.n239 163.367
R692 B.n402 B.n239 163.367
R693 B.n402 B.n237 163.367
R694 B.n406 B.n237 163.367
R695 B.n406 B.n231 163.367
R696 B.n414 B.n231 163.367
R697 B.n414 B.n229 163.367
R698 B.n418 B.n229 163.367
R699 B.n418 B.n223 163.367
R700 B.n426 B.n223 163.367
R701 B.n426 B.n221 163.367
R702 B.n430 B.n221 163.367
R703 B.n430 B.n215 163.367
R704 B.n438 B.n215 163.367
R705 B.n438 B.n213 163.367
R706 B.n442 B.n213 163.367
R707 B.n442 B.n207 163.367
R708 B.n450 B.n207 163.367
R709 B.n450 B.n205 163.367
R710 B.n454 B.n205 163.367
R711 B.n454 B.n199 163.367
R712 B.n462 B.n199 163.367
R713 B.n462 B.n197 163.367
R714 B.n466 B.n197 163.367
R715 B.n466 B.n191 163.367
R716 B.n474 B.n191 163.367
R717 B.n474 B.n189 163.367
R718 B.n478 B.n189 163.367
R719 B.n478 B.n183 163.367
R720 B.n487 B.n183 163.367
R721 B.n487 B.n181 163.367
R722 B.n491 B.n181 163.367
R723 B.n491 B.n176 163.367
R724 B.n500 B.n176 163.367
R725 B.n500 B.n174 163.367
R726 B.n504 B.n174 163.367
R727 B.n504 B.n2 163.367
R728 B.n686 B.n2 163.367
R729 B.n686 B.n3 163.367
R730 B.n682 B.n3 163.367
R731 B.n682 B.n9 163.367
R732 B.n678 B.n9 163.367
R733 B.n678 B.n11 163.367
R734 B.n674 B.n11 163.367
R735 B.n674 B.n15 163.367
R736 B.n670 B.n15 163.367
R737 B.n670 B.n17 163.367
R738 B.n666 B.n17 163.367
R739 B.n666 B.n23 163.367
R740 B.n662 B.n23 163.367
R741 B.n662 B.n25 163.367
R742 B.n658 B.n25 163.367
R743 B.n658 B.n30 163.367
R744 B.n654 B.n30 163.367
R745 B.n654 B.n32 163.367
R746 B.n650 B.n32 163.367
R747 B.n650 B.n37 163.367
R748 B.n646 B.n37 163.367
R749 B.n646 B.n39 163.367
R750 B.n642 B.n39 163.367
R751 B.n642 B.n44 163.367
R752 B.n638 B.n44 163.367
R753 B.n638 B.n46 163.367
R754 B.n634 B.n46 163.367
R755 B.n634 B.n51 163.367
R756 B.n630 B.n51 163.367
R757 B.n630 B.n53 163.367
R758 B.n626 B.n53 163.367
R759 B.n626 B.n58 163.367
R760 B.n622 B.n58 163.367
R761 B.n622 B.n60 163.367
R762 B.n618 B.n60 163.367
R763 B.n618 B.n65 163.367
R764 B.n614 B.n65 163.367
R765 B.n614 B.n67 163.367
R766 B.n610 B.n67 163.367
R767 B.n610 B.n72 163.367
R768 B.n606 B.n72 163.367
R769 B.n606 B.n74 163.367
R770 B.n602 B.n74 163.367
R771 B.n602 B.n79 163.367
R772 B.n598 B.n79 163.367
R773 B.n598 B.n81 163.367
R774 B.n594 B.n81 163.367
R775 B.n594 B.n86 163.367
R776 B.n590 B.n86 163.367
R777 B.n590 B.n88 163.367
R778 B.n586 B.n88 163.367
R779 B.n586 B.n93 163.367
R780 B.n582 B.n93 163.367
R781 B.n582 B.n95 163.367
R782 B.n289 B.n288 163.367
R783 B.n340 B.n288 163.367
R784 B.n338 B.n337 163.367
R785 B.n334 B.n333 163.367
R786 B.n330 B.n329 163.367
R787 B.n326 B.n325 163.367
R788 B.n322 B.n321 163.367
R789 B.n318 B.n317 163.367
R790 B.n314 B.n313 163.367
R791 B.n310 B.n309 163.367
R792 B.n306 B.n305 163.367
R793 B.n302 B.n301 163.367
R794 B.n298 B.n297 163.367
R795 B.n348 B.n275 163.367
R796 B.n352 B.n273 163.367
R797 B.n352 B.n267 163.367
R798 B.n360 B.n267 163.367
R799 B.n360 B.n265 163.367
R800 B.n364 B.n265 163.367
R801 B.n364 B.n259 163.367
R802 B.n372 B.n259 163.367
R803 B.n372 B.n257 163.367
R804 B.n376 B.n257 163.367
R805 B.n376 B.n251 163.367
R806 B.n384 B.n251 163.367
R807 B.n384 B.n249 163.367
R808 B.n388 B.n249 163.367
R809 B.n388 B.n243 163.367
R810 B.n396 B.n243 163.367
R811 B.n396 B.n241 163.367
R812 B.n400 B.n241 163.367
R813 B.n400 B.n234 163.367
R814 B.n408 B.n234 163.367
R815 B.n408 B.n232 163.367
R816 B.n412 B.n232 163.367
R817 B.n412 B.n227 163.367
R818 B.n420 B.n227 163.367
R819 B.n420 B.n225 163.367
R820 B.n424 B.n225 163.367
R821 B.n424 B.n219 163.367
R822 B.n432 B.n219 163.367
R823 B.n432 B.n217 163.367
R824 B.n436 B.n217 163.367
R825 B.n436 B.n211 163.367
R826 B.n444 B.n211 163.367
R827 B.n444 B.n209 163.367
R828 B.n448 B.n209 163.367
R829 B.n448 B.n203 163.367
R830 B.n456 B.n203 163.367
R831 B.n456 B.n201 163.367
R832 B.n460 B.n201 163.367
R833 B.n460 B.n195 163.367
R834 B.n468 B.n195 163.367
R835 B.n468 B.n193 163.367
R836 B.n472 B.n193 163.367
R837 B.n472 B.n187 163.367
R838 B.n480 B.n187 163.367
R839 B.n480 B.n185 163.367
R840 B.n484 B.n185 163.367
R841 B.n484 B.n180 163.367
R842 B.n493 B.n180 163.367
R843 B.n493 B.n178 163.367
R844 B.n498 B.n178 163.367
R845 B.n498 B.n172 163.367
R846 B.n506 B.n172 163.367
R847 B.n507 B.n506 163.367
R848 B.n507 B.n5 163.367
R849 B.n6 B.n5 163.367
R850 B.n7 B.n6 163.367
R851 B.n512 B.n7 163.367
R852 B.n512 B.n12 163.367
R853 B.n13 B.n12 163.367
R854 B.n14 B.n13 163.367
R855 B.n517 B.n14 163.367
R856 B.n517 B.n19 163.367
R857 B.n20 B.n19 163.367
R858 B.n21 B.n20 163.367
R859 B.n522 B.n21 163.367
R860 B.n522 B.n26 163.367
R861 B.n27 B.n26 163.367
R862 B.n28 B.n27 163.367
R863 B.n527 B.n28 163.367
R864 B.n527 B.n33 163.367
R865 B.n34 B.n33 163.367
R866 B.n35 B.n34 163.367
R867 B.n532 B.n35 163.367
R868 B.n532 B.n40 163.367
R869 B.n41 B.n40 163.367
R870 B.n42 B.n41 163.367
R871 B.n537 B.n42 163.367
R872 B.n537 B.n47 163.367
R873 B.n48 B.n47 163.367
R874 B.n49 B.n48 163.367
R875 B.n542 B.n49 163.367
R876 B.n542 B.n54 163.367
R877 B.n55 B.n54 163.367
R878 B.n56 B.n55 163.367
R879 B.n547 B.n56 163.367
R880 B.n547 B.n61 163.367
R881 B.n62 B.n61 163.367
R882 B.n63 B.n62 163.367
R883 B.n552 B.n63 163.367
R884 B.n552 B.n68 163.367
R885 B.n69 B.n68 163.367
R886 B.n70 B.n69 163.367
R887 B.n557 B.n70 163.367
R888 B.n557 B.n75 163.367
R889 B.n76 B.n75 163.367
R890 B.n77 B.n76 163.367
R891 B.n562 B.n77 163.367
R892 B.n562 B.n82 163.367
R893 B.n83 B.n82 163.367
R894 B.n84 B.n83 163.367
R895 B.n567 B.n84 163.367
R896 B.n567 B.n89 163.367
R897 B.n90 B.n89 163.367
R898 B.n91 B.n90 163.367
R899 B.n572 B.n91 163.367
R900 B.n572 B.n96 163.367
R901 B.n97 B.n96 163.367
R902 B.n120 B.n119 163.367
R903 B.n124 B.n123 163.367
R904 B.n128 B.n127 163.367
R905 B.n132 B.n131 163.367
R906 B.n137 B.n136 163.367
R907 B.n141 B.n140 163.367
R908 B.n145 B.n144 163.367
R909 B.n149 B.n148 163.367
R910 B.n153 B.n152 163.367
R911 B.n158 B.n157 163.367
R912 B.n162 B.n161 163.367
R913 B.n166 B.n165 163.367
R914 B.n168 B.n111 163.367
R915 B.n353 B.n272 120.162
R916 B.n353 B.n268 120.162
R917 B.n359 B.n268 120.162
R918 B.n359 B.n264 120.162
R919 B.n365 B.n264 120.162
R920 B.n365 B.n260 120.162
R921 B.n371 B.n260 120.162
R922 B.n377 B.n256 120.162
R923 B.n377 B.n252 120.162
R924 B.n383 B.n252 120.162
R925 B.n383 B.n248 120.162
R926 B.n389 B.n248 120.162
R927 B.n389 B.n244 120.162
R928 B.n395 B.n244 120.162
R929 B.n395 B.n240 120.162
R930 B.n401 B.n240 120.162
R931 B.n401 B.n235 120.162
R932 B.n407 B.n235 120.162
R933 B.n407 B.n236 120.162
R934 B.n413 B.n228 120.162
R935 B.n419 B.n228 120.162
R936 B.n419 B.n224 120.162
R937 B.n425 B.n224 120.162
R938 B.n425 B.n220 120.162
R939 B.n431 B.n220 120.162
R940 B.n431 B.n216 120.162
R941 B.n437 B.n216 120.162
R942 B.n443 B.n212 120.162
R943 B.n443 B.n208 120.162
R944 B.n449 B.n208 120.162
R945 B.n449 B.n204 120.162
R946 B.n455 B.n204 120.162
R947 B.n455 B.n200 120.162
R948 B.n461 B.n200 120.162
R949 B.n467 B.n196 120.162
R950 B.n467 B.n192 120.162
R951 B.n473 B.n192 120.162
R952 B.n473 B.n188 120.162
R953 B.n479 B.n188 120.162
R954 B.n479 B.n184 120.162
R955 B.n486 B.n184 120.162
R956 B.n486 B.n485 120.162
R957 B.n492 B.n177 120.162
R958 B.n499 B.n177 120.162
R959 B.n499 B.n173 120.162
R960 B.n505 B.n173 120.162
R961 B.n505 B.n4 120.162
R962 B.n685 B.n4 120.162
R963 B.n685 B.n684 120.162
R964 B.n684 B.n683 120.162
R965 B.n683 B.n8 120.162
R966 B.n677 B.n8 120.162
R967 B.n677 B.n676 120.162
R968 B.n676 B.n675 120.162
R969 B.n669 B.n18 120.162
R970 B.n669 B.n668 120.162
R971 B.n668 B.n667 120.162
R972 B.n667 B.n22 120.162
R973 B.n661 B.n22 120.162
R974 B.n661 B.n660 120.162
R975 B.n660 B.n659 120.162
R976 B.n659 B.n29 120.162
R977 B.n653 B.n652 120.162
R978 B.n652 B.n651 120.162
R979 B.n651 B.n36 120.162
R980 B.n645 B.n36 120.162
R981 B.n645 B.n644 120.162
R982 B.n644 B.n643 120.162
R983 B.n643 B.n43 120.162
R984 B.n637 B.n636 120.162
R985 B.n636 B.n635 120.162
R986 B.n635 B.n50 120.162
R987 B.n629 B.n50 120.162
R988 B.n629 B.n628 120.162
R989 B.n628 B.n627 120.162
R990 B.n627 B.n57 120.162
R991 B.n621 B.n57 120.162
R992 B.n620 B.n619 120.162
R993 B.n619 B.n64 120.162
R994 B.n613 B.n64 120.162
R995 B.n613 B.n612 120.162
R996 B.n612 B.n611 120.162
R997 B.n611 B.n71 120.162
R998 B.n605 B.n71 120.162
R999 B.n605 B.n604 120.162
R1000 B.n604 B.n603 120.162
R1001 B.n603 B.n78 120.162
R1002 B.n597 B.n78 120.162
R1003 B.n597 B.n596 120.162
R1004 B.n595 B.n85 120.162
R1005 B.n589 B.n85 120.162
R1006 B.n589 B.n588 120.162
R1007 B.n588 B.n587 120.162
R1008 B.n587 B.n92 120.162
R1009 B.n581 B.n92 120.162
R1010 B.n581 B.n580 120.162
R1011 B.n461 B.t6 118.394
R1012 B.n653 B.t5 118.394
R1013 B.n371 B.t16 114.859
R1014 B.t1 B.n212 114.859
R1015 B.t4 B.n43 114.859
R1016 B.t9 B.n595 114.859
R1017 B.n485 B.t7 111.326
R1018 B.n18 B.t3 111.326
R1019 B.n413 B.t0 107.791
R1020 B.n621 B.t2 107.791
R1021 B.n346 B.n345 71.676
R1022 B.n340 B.n276 71.676
R1023 B.n337 B.n277 71.676
R1024 B.n333 B.n278 71.676
R1025 B.n329 B.n279 71.676
R1026 B.n325 B.n280 71.676
R1027 B.n321 B.n281 71.676
R1028 B.n317 B.n282 71.676
R1029 B.n313 B.n283 71.676
R1030 B.n309 B.n284 71.676
R1031 B.n305 B.n285 71.676
R1032 B.n301 B.n286 71.676
R1033 B.n297 B.n287 71.676
R1034 B.n116 B.n98 71.676
R1035 B.n120 B.n99 71.676
R1036 B.n124 B.n100 71.676
R1037 B.n128 B.n101 71.676
R1038 B.n132 B.n102 71.676
R1039 B.n137 B.n103 71.676
R1040 B.n141 B.n104 71.676
R1041 B.n145 B.n105 71.676
R1042 B.n149 B.n106 71.676
R1043 B.n153 B.n107 71.676
R1044 B.n158 B.n108 71.676
R1045 B.n162 B.n109 71.676
R1046 B.n166 B.n110 71.676
R1047 B.n578 B.n111 71.676
R1048 B.n578 B.n577 71.676
R1049 B.n168 B.n110 71.676
R1050 B.n165 B.n109 71.676
R1051 B.n161 B.n108 71.676
R1052 B.n157 B.n107 71.676
R1053 B.n152 B.n106 71.676
R1054 B.n148 B.n105 71.676
R1055 B.n144 B.n104 71.676
R1056 B.n140 B.n103 71.676
R1057 B.n136 B.n102 71.676
R1058 B.n131 B.n101 71.676
R1059 B.n127 B.n100 71.676
R1060 B.n123 B.n99 71.676
R1061 B.n119 B.n98 71.676
R1062 B.n346 B.n289 71.676
R1063 B.n338 B.n276 71.676
R1064 B.n334 B.n277 71.676
R1065 B.n330 B.n278 71.676
R1066 B.n326 B.n279 71.676
R1067 B.n322 B.n280 71.676
R1068 B.n318 B.n281 71.676
R1069 B.n314 B.n282 71.676
R1070 B.n310 B.n283 71.676
R1071 B.n306 B.n284 71.676
R1072 B.n302 B.n285 71.676
R1073 B.n298 B.n286 71.676
R1074 B.n287 B.n275 71.676
R1075 B.n295 B.n294 59.5399
R1076 B.n292 B.n291 59.5399
R1077 B.n134 B.n115 59.5399
R1078 B.n155 B.n113 59.5399
R1079 B.n294 B.n293 58.9581
R1080 B.n291 B.n290 58.9581
R1081 B.n115 B.n114 58.9581
R1082 B.n113 B.n112 58.9581
R1083 B.n117 B.n94 29.5029
R1084 B.n350 B.n349 29.5029
R1085 B.n344 B.n270 29.5029
R1086 B.n576 B.n575 29.5029
R1087 B B.n687 18.0485
R1088 B.n236 B.t0 12.37
R1089 B.t2 B.n620 12.37
R1090 B.n118 B.n117 10.6151
R1091 B.n121 B.n118 10.6151
R1092 B.n122 B.n121 10.6151
R1093 B.n125 B.n122 10.6151
R1094 B.n126 B.n125 10.6151
R1095 B.n129 B.n126 10.6151
R1096 B.n130 B.n129 10.6151
R1097 B.n133 B.n130 10.6151
R1098 B.n138 B.n135 10.6151
R1099 B.n139 B.n138 10.6151
R1100 B.n142 B.n139 10.6151
R1101 B.n143 B.n142 10.6151
R1102 B.n146 B.n143 10.6151
R1103 B.n147 B.n146 10.6151
R1104 B.n150 B.n147 10.6151
R1105 B.n151 B.n150 10.6151
R1106 B.n154 B.n151 10.6151
R1107 B.n159 B.n156 10.6151
R1108 B.n160 B.n159 10.6151
R1109 B.n163 B.n160 10.6151
R1110 B.n164 B.n163 10.6151
R1111 B.n167 B.n164 10.6151
R1112 B.n169 B.n167 10.6151
R1113 B.n170 B.n169 10.6151
R1114 B.n576 B.n170 10.6151
R1115 B.n351 B.n350 10.6151
R1116 B.n351 B.n266 10.6151
R1117 B.n361 B.n266 10.6151
R1118 B.n362 B.n361 10.6151
R1119 B.n363 B.n362 10.6151
R1120 B.n363 B.n258 10.6151
R1121 B.n373 B.n258 10.6151
R1122 B.n374 B.n373 10.6151
R1123 B.n375 B.n374 10.6151
R1124 B.n375 B.n250 10.6151
R1125 B.n385 B.n250 10.6151
R1126 B.n386 B.n385 10.6151
R1127 B.n387 B.n386 10.6151
R1128 B.n387 B.n242 10.6151
R1129 B.n397 B.n242 10.6151
R1130 B.n398 B.n397 10.6151
R1131 B.n399 B.n398 10.6151
R1132 B.n399 B.n233 10.6151
R1133 B.n409 B.n233 10.6151
R1134 B.n410 B.n409 10.6151
R1135 B.n411 B.n410 10.6151
R1136 B.n411 B.n226 10.6151
R1137 B.n421 B.n226 10.6151
R1138 B.n422 B.n421 10.6151
R1139 B.n423 B.n422 10.6151
R1140 B.n423 B.n218 10.6151
R1141 B.n433 B.n218 10.6151
R1142 B.n434 B.n433 10.6151
R1143 B.n435 B.n434 10.6151
R1144 B.n435 B.n210 10.6151
R1145 B.n445 B.n210 10.6151
R1146 B.n446 B.n445 10.6151
R1147 B.n447 B.n446 10.6151
R1148 B.n447 B.n202 10.6151
R1149 B.n457 B.n202 10.6151
R1150 B.n458 B.n457 10.6151
R1151 B.n459 B.n458 10.6151
R1152 B.n459 B.n194 10.6151
R1153 B.n469 B.n194 10.6151
R1154 B.n470 B.n469 10.6151
R1155 B.n471 B.n470 10.6151
R1156 B.n471 B.n186 10.6151
R1157 B.n481 B.n186 10.6151
R1158 B.n482 B.n481 10.6151
R1159 B.n483 B.n482 10.6151
R1160 B.n483 B.n179 10.6151
R1161 B.n494 B.n179 10.6151
R1162 B.n495 B.n494 10.6151
R1163 B.n497 B.n495 10.6151
R1164 B.n497 B.n496 10.6151
R1165 B.n496 B.n171 10.6151
R1166 B.n508 B.n171 10.6151
R1167 B.n509 B.n508 10.6151
R1168 B.n510 B.n509 10.6151
R1169 B.n511 B.n510 10.6151
R1170 B.n513 B.n511 10.6151
R1171 B.n514 B.n513 10.6151
R1172 B.n515 B.n514 10.6151
R1173 B.n516 B.n515 10.6151
R1174 B.n518 B.n516 10.6151
R1175 B.n519 B.n518 10.6151
R1176 B.n520 B.n519 10.6151
R1177 B.n521 B.n520 10.6151
R1178 B.n523 B.n521 10.6151
R1179 B.n524 B.n523 10.6151
R1180 B.n525 B.n524 10.6151
R1181 B.n526 B.n525 10.6151
R1182 B.n528 B.n526 10.6151
R1183 B.n529 B.n528 10.6151
R1184 B.n530 B.n529 10.6151
R1185 B.n531 B.n530 10.6151
R1186 B.n533 B.n531 10.6151
R1187 B.n534 B.n533 10.6151
R1188 B.n535 B.n534 10.6151
R1189 B.n536 B.n535 10.6151
R1190 B.n538 B.n536 10.6151
R1191 B.n539 B.n538 10.6151
R1192 B.n540 B.n539 10.6151
R1193 B.n541 B.n540 10.6151
R1194 B.n543 B.n541 10.6151
R1195 B.n544 B.n543 10.6151
R1196 B.n545 B.n544 10.6151
R1197 B.n546 B.n545 10.6151
R1198 B.n548 B.n546 10.6151
R1199 B.n549 B.n548 10.6151
R1200 B.n550 B.n549 10.6151
R1201 B.n551 B.n550 10.6151
R1202 B.n553 B.n551 10.6151
R1203 B.n554 B.n553 10.6151
R1204 B.n555 B.n554 10.6151
R1205 B.n556 B.n555 10.6151
R1206 B.n558 B.n556 10.6151
R1207 B.n559 B.n558 10.6151
R1208 B.n560 B.n559 10.6151
R1209 B.n561 B.n560 10.6151
R1210 B.n563 B.n561 10.6151
R1211 B.n564 B.n563 10.6151
R1212 B.n565 B.n564 10.6151
R1213 B.n566 B.n565 10.6151
R1214 B.n568 B.n566 10.6151
R1215 B.n569 B.n568 10.6151
R1216 B.n570 B.n569 10.6151
R1217 B.n571 B.n570 10.6151
R1218 B.n573 B.n571 10.6151
R1219 B.n574 B.n573 10.6151
R1220 B.n575 B.n574 10.6151
R1221 B.n344 B.n343 10.6151
R1222 B.n343 B.n342 10.6151
R1223 B.n342 B.n341 10.6151
R1224 B.n341 B.n339 10.6151
R1225 B.n339 B.n336 10.6151
R1226 B.n336 B.n335 10.6151
R1227 B.n335 B.n332 10.6151
R1228 B.n332 B.n331 10.6151
R1229 B.n328 B.n327 10.6151
R1230 B.n327 B.n324 10.6151
R1231 B.n324 B.n323 10.6151
R1232 B.n323 B.n320 10.6151
R1233 B.n320 B.n319 10.6151
R1234 B.n319 B.n316 10.6151
R1235 B.n316 B.n315 10.6151
R1236 B.n315 B.n312 10.6151
R1237 B.n312 B.n311 10.6151
R1238 B.n308 B.n307 10.6151
R1239 B.n307 B.n304 10.6151
R1240 B.n304 B.n303 10.6151
R1241 B.n303 B.n300 10.6151
R1242 B.n300 B.n299 10.6151
R1243 B.n299 B.n296 10.6151
R1244 B.n296 B.n274 10.6151
R1245 B.n349 B.n274 10.6151
R1246 B.n355 B.n270 10.6151
R1247 B.n356 B.n355 10.6151
R1248 B.n357 B.n356 10.6151
R1249 B.n357 B.n262 10.6151
R1250 B.n367 B.n262 10.6151
R1251 B.n368 B.n367 10.6151
R1252 B.n369 B.n368 10.6151
R1253 B.n369 B.n254 10.6151
R1254 B.n379 B.n254 10.6151
R1255 B.n380 B.n379 10.6151
R1256 B.n381 B.n380 10.6151
R1257 B.n381 B.n246 10.6151
R1258 B.n391 B.n246 10.6151
R1259 B.n392 B.n391 10.6151
R1260 B.n393 B.n392 10.6151
R1261 B.n393 B.n238 10.6151
R1262 B.n403 B.n238 10.6151
R1263 B.n404 B.n403 10.6151
R1264 B.n405 B.n404 10.6151
R1265 B.n405 B.n230 10.6151
R1266 B.n415 B.n230 10.6151
R1267 B.n416 B.n415 10.6151
R1268 B.n417 B.n416 10.6151
R1269 B.n417 B.n222 10.6151
R1270 B.n427 B.n222 10.6151
R1271 B.n428 B.n427 10.6151
R1272 B.n429 B.n428 10.6151
R1273 B.n429 B.n214 10.6151
R1274 B.n439 B.n214 10.6151
R1275 B.n440 B.n439 10.6151
R1276 B.n441 B.n440 10.6151
R1277 B.n441 B.n206 10.6151
R1278 B.n451 B.n206 10.6151
R1279 B.n452 B.n451 10.6151
R1280 B.n453 B.n452 10.6151
R1281 B.n453 B.n198 10.6151
R1282 B.n463 B.n198 10.6151
R1283 B.n464 B.n463 10.6151
R1284 B.n465 B.n464 10.6151
R1285 B.n465 B.n190 10.6151
R1286 B.n475 B.n190 10.6151
R1287 B.n476 B.n475 10.6151
R1288 B.n477 B.n476 10.6151
R1289 B.n477 B.n182 10.6151
R1290 B.n488 B.n182 10.6151
R1291 B.n489 B.n488 10.6151
R1292 B.n490 B.n489 10.6151
R1293 B.n490 B.n175 10.6151
R1294 B.n501 B.n175 10.6151
R1295 B.n502 B.n501 10.6151
R1296 B.n503 B.n502 10.6151
R1297 B.n503 B.n0 10.6151
R1298 B.n681 B.n1 10.6151
R1299 B.n681 B.n680 10.6151
R1300 B.n680 B.n679 10.6151
R1301 B.n679 B.n10 10.6151
R1302 B.n673 B.n10 10.6151
R1303 B.n673 B.n672 10.6151
R1304 B.n672 B.n671 10.6151
R1305 B.n671 B.n16 10.6151
R1306 B.n665 B.n16 10.6151
R1307 B.n665 B.n664 10.6151
R1308 B.n664 B.n663 10.6151
R1309 B.n663 B.n24 10.6151
R1310 B.n657 B.n24 10.6151
R1311 B.n657 B.n656 10.6151
R1312 B.n656 B.n655 10.6151
R1313 B.n655 B.n31 10.6151
R1314 B.n649 B.n31 10.6151
R1315 B.n649 B.n648 10.6151
R1316 B.n648 B.n647 10.6151
R1317 B.n647 B.n38 10.6151
R1318 B.n641 B.n38 10.6151
R1319 B.n641 B.n640 10.6151
R1320 B.n640 B.n639 10.6151
R1321 B.n639 B.n45 10.6151
R1322 B.n633 B.n45 10.6151
R1323 B.n633 B.n632 10.6151
R1324 B.n632 B.n631 10.6151
R1325 B.n631 B.n52 10.6151
R1326 B.n625 B.n52 10.6151
R1327 B.n625 B.n624 10.6151
R1328 B.n624 B.n623 10.6151
R1329 B.n623 B.n59 10.6151
R1330 B.n617 B.n59 10.6151
R1331 B.n617 B.n616 10.6151
R1332 B.n616 B.n615 10.6151
R1333 B.n615 B.n66 10.6151
R1334 B.n609 B.n66 10.6151
R1335 B.n609 B.n608 10.6151
R1336 B.n608 B.n607 10.6151
R1337 B.n607 B.n73 10.6151
R1338 B.n601 B.n73 10.6151
R1339 B.n601 B.n600 10.6151
R1340 B.n600 B.n599 10.6151
R1341 B.n599 B.n80 10.6151
R1342 B.n593 B.n80 10.6151
R1343 B.n593 B.n592 10.6151
R1344 B.n592 B.n591 10.6151
R1345 B.n591 B.n87 10.6151
R1346 B.n585 B.n87 10.6151
R1347 B.n585 B.n584 10.6151
R1348 B.n584 B.n583 10.6151
R1349 B.n583 B.n94 10.6151
R1350 B.n134 B.n133 9.36635
R1351 B.n156 B.n155 9.36635
R1352 B.n331 B.n292 9.36635
R1353 B.n308 B.n295 9.36635
R1354 B.n492 B.t7 8.83584
R1355 B.n675 B.t3 8.83584
R1356 B.t16 B.n256 5.3017
R1357 B.n437 B.t1 5.3017
R1358 B.n637 B.t4 5.3017
R1359 B.n596 B.t9 5.3017
R1360 B.n687 B.n0 2.81026
R1361 B.n687 B.n1 2.81026
R1362 B.t6 B.n196 1.76757
R1363 B.t5 B.n29 1.76757
R1364 B.n135 B.n134 1.24928
R1365 B.n155 B.n154 1.24928
R1366 B.n328 B.n292 1.24928
R1367 B.n311 B.n295 1.24928
R1368 VP.n21 VP.n20 161.3
R1369 VP.n22 VP.n17 161.3
R1370 VP.n24 VP.n23 161.3
R1371 VP.n25 VP.n16 161.3
R1372 VP.n27 VP.n26 161.3
R1373 VP.n28 VP.n15 161.3
R1374 VP.n30 VP.n29 161.3
R1375 VP.n32 VP.n31 161.3
R1376 VP.n33 VP.n13 161.3
R1377 VP.n35 VP.n34 161.3
R1378 VP.n36 VP.n12 161.3
R1379 VP.n38 VP.n37 161.3
R1380 VP.n39 VP.n11 161.3
R1381 VP.n72 VP.n0 161.3
R1382 VP.n71 VP.n70 161.3
R1383 VP.n69 VP.n1 161.3
R1384 VP.n68 VP.n67 161.3
R1385 VP.n66 VP.n2 161.3
R1386 VP.n65 VP.n64 161.3
R1387 VP.n63 VP.n62 161.3
R1388 VP.n61 VP.n4 161.3
R1389 VP.n60 VP.n59 161.3
R1390 VP.n58 VP.n5 161.3
R1391 VP.n57 VP.n56 161.3
R1392 VP.n55 VP.n6 161.3
R1393 VP.n54 VP.n53 161.3
R1394 VP.n52 VP.n51 161.3
R1395 VP.n50 VP.n8 161.3
R1396 VP.n49 VP.n48 161.3
R1397 VP.n47 VP.n9 161.3
R1398 VP.n46 VP.n45 161.3
R1399 VP.n44 VP.n10 161.3
R1400 VP.n43 VP.n42 107.82
R1401 VP.n74 VP.n73 107.82
R1402 VP.n41 VP.n40 107.82
R1403 VP.n19 VP.n18 72.3368
R1404 VP.n49 VP.n9 44.3785
R1405 VP.n67 VP.n1 44.3785
R1406 VP.n34 VP.n12 44.3785
R1407 VP.n42 VP.n41 42.9769
R1408 VP.n56 VP.n5 40.4934
R1409 VP.n60 VP.n5 40.4934
R1410 VP.n27 VP.n16 40.4934
R1411 VP.n23 VP.n16 40.4934
R1412 VP.n19 VP.t2 39.5494
R1413 VP.n50 VP.n49 36.6083
R1414 VP.n67 VP.n66 36.6083
R1415 VP.n34 VP.n33 36.6083
R1416 VP.n45 VP.n44 24.4675
R1417 VP.n45 VP.n9 24.4675
R1418 VP.n51 VP.n50 24.4675
R1419 VP.n55 VP.n54 24.4675
R1420 VP.n56 VP.n55 24.4675
R1421 VP.n61 VP.n60 24.4675
R1422 VP.n62 VP.n61 24.4675
R1423 VP.n66 VP.n65 24.4675
R1424 VP.n71 VP.n1 24.4675
R1425 VP.n72 VP.n71 24.4675
R1426 VP.n38 VP.n12 24.4675
R1427 VP.n39 VP.n38 24.4675
R1428 VP.n28 VP.n27 24.4675
R1429 VP.n29 VP.n28 24.4675
R1430 VP.n33 VP.n32 24.4675
R1431 VP.n22 VP.n21 24.4675
R1432 VP.n23 VP.n22 24.4675
R1433 VP.n51 VP.n7 23.4888
R1434 VP.n65 VP.n3 23.4888
R1435 VP.n32 VP.n14 23.4888
R1436 VP.n43 VP.t5 8.44884
R1437 VP.n7 VP.t0 8.44884
R1438 VP.n3 VP.t4 8.44884
R1439 VP.n73 VP.t7 8.44884
R1440 VP.n40 VP.t1 8.44884
R1441 VP.n14 VP.t3 8.44884
R1442 VP.n18 VP.t6 8.44884
R1443 VP.n20 VP.n19 7.30997
R1444 VP.n44 VP.n43 2.93654
R1445 VP.n73 VP.n72 2.93654
R1446 VP.n40 VP.n39 2.93654
R1447 VP.n54 VP.n7 0.97918
R1448 VP.n62 VP.n3 0.97918
R1449 VP.n29 VP.n14 0.97918
R1450 VP.n21 VP.n18 0.97918
R1451 VP.n41 VP.n11 0.278367
R1452 VP.n42 VP.n10 0.278367
R1453 VP.n74 VP.n0 0.278367
R1454 VP.n20 VP.n17 0.189894
R1455 VP.n24 VP.n17 0.189894
R1456 VP.n25 VP.n24 0.189894
R1457 VP.n26 VP.n25 0.189894
R1458 VP.n26 VP.n15 0.189894
R1459 VP.n30 VP.n15 0.189894
R1460 VP.n31 VP.n30 0.189894
R1461 VP.n31 VP.n13 0.189894
R1462 VP.n35 VP.n13 0.189894
R1463 VP.n36 VP.n35 0.189894
R1464 VP.n37 VP.n36 0.189894
R1465 VP.n37 VP.n11 0.189894
R1466 VP.n46 VP.n10 0.189894
R1467 VP.n47 VP.n46 0.189894
R1468 VP.n48 VP.n47 0.189894
R1469 VP.n48 VP.n8 0.189894
R1470 VP.n52 VP.n8 0.189894
R1471 VP.n53 VP.n52 0.189894
R1472 VP.n53 VP.n6 0.189894
R1473 VP.n57 VP.n6 0.189894
R1474 VP.n58 VP.n57 0.189894
R1475 VP.n59 VP.n58 0.189894
R1476 VP.n59 VP.n4 0.189894
R1477 VP.n63 VP.n4 0.189894
R1478 VP.n64 VP.n63 0.189894
R1479 VP.n64 VP.n2 0.189894
R1480 VP.n68 VP.n2 0.189894
R1481 VP.n69 VP.n68 0.189894
R1482 VP.n70 VP.n69 0.189894
R1483 VP.n70 VP.n0 0.189894
R1484 VP VP.n74 0.153454
R1485 VDD1 VDD1.n0 240.531
R1486 VDD1.n3 VDD1.n2 240.417
R1487 VDD1.n3 VDD1.n1 240.417
R1488 VDD1.n5 VDD1.n4 239.163
R1489 VDD1.n5 VDD1.n3 36.9104
R1490 VDD1.n4 VDD1.t4 20.8426
R1491 VDD1.n4 VDD1.t6 20.8426
R1492 VDD1.n0 VDD1.t5 20.8426
R1493 VDD1.n0 VDD1.t1 20.8426
R1494 VDD1.n2 VDD1.t3 20.8426
R1495 VDD1.n2 VDD1.t0 20.8426
R1496 VDD1.n1 VDD1.t2 20.8426
R1497 VDD1.n1 VDD1.t7 20.8426
R1498 VDD1 VDD1.n5 1.25266
C0 VTAIL VN 2.46448f
C1 VDD1 VTAIL 4.46352f
C2 VTAIL VP 2.47859f
C3 VDD1 VN 0.158775f
C4 VN VP 5.76194f
C5 VTAIL VDD2 4.51867f
C6 VDD1 VP 1.50609f
C7 VN VDD2 1.12855f
C8 VDD1 VDD2 1.83226f
C9 VP VDD2 0.540181f
C10 VDD2 B 4.40628f
C11 VDD1 B 4.836695f
C12 VTAIL B 3.419684f
C13 VN B 15.00364f
C14 VP B 13.488044f
C15 VDD1.t5 B 0.014211f
C16 VDD1.t1 B 0.014211f
C17 VDD1.n0 B 0.05733f
C18 VDD1.t2 B 0.014211f
C19 VDD1.t7 B 0.014211f
C20 VDD1.n1 B 0.057118f
C21 VDD1.t3 B 0.014211f
C22 VDD1.t0 B 0.014211f
C23 VDD1.n2 B 0.057118f
C24 VDD1.n3 B 2.01785f
C25 VDD1.t4 B 0.014211f
C26 VDD1.t6 B 0.014211f
C27 VDD1.n4 B 0.055173f
C28 VDD1.n5 B 1.60486f
C29 VP.n0 B 0.040475f
C30 VP.t7 B 0.143782f
C31 VP.n1 B 0.059497f
C32 VP.n2 B 0.0307f
C33 VP.t4 B 0.143782f
C34 VP.n3 B 0.102083f
C35 VP.n4 B 0.0307f
C36 VP.n5 B 0.024818f
C37 VP.n6 B 0.0307f
C38 VP.t0 B 0.143782f
C39 VP.n7 B 0.102083f
C40 VP.n8 B 0.0307f
C41 VP.n9 B 0.059497f
C42 VP.n10 B 0.040475f
C43 VP.t5 B 0.143782f
C44 VP.n11 B 0.040475f
C45 VP.t1 B 0.143782f
C46 VP.n12 B 0.059497f
C47 VP.n13 B 0.0307f
C48 VP.t3 B 0.143782f
C49 VP.n14 B 0.102083f
C50 VP.n15 B 0.0307f
C51 VP.n16 B 0.024818f
C52 VP.n17 B 0.0307f
C53 VP.t6 B 0.143782f
C54 VP.n18 B 0.182356f
C55 VP.t2 B 0.374835f
C56 VP.n19 B 0.195694f
C57 VP.n20 B 0.299817f
C58 VP.n21 B 0.030099f
C59 VP.n22 B 0.057218f
C60 VP.n23 B 0.061017f
C61 VP.n24 B 0.0307f
C62 VP.n25 B 0.0307f
C63 VP.n26 B 0.0307f
C64 VP.n27 B 0.061017f
C65 VP.n28 B 0.057218f
C66 VP.n29 B 0.030099f
C67 VP.n30 B 0.0307f
C68 VP.n31 B 0.0307f
C69 VP.n32 B 0.056088f
C70 VP.n33 B 0.0619f
C71 VP.n34 B 0.025455f
C72 VP.n35 B 0.0307f
C73 VP.n36 B 0.0307f
C74 VP.n37 B 0.0307f
C75 VP.n38 B 0.057218f
C76 VP.n39 B 0.032359f
C77 VP.n40 B 0.197878f
C78 VP.n41 B 1.36097f
C79 VP.n42 B 1.38665f
C80 VP.n43 B 0.197878f
C81 VP.n44 B 0.032359f
C82 VP.n45 B 0.057218f
C83 VP.n46 B 0.0307f
C84 VP.n47 B 0.0307f
C85 VP.n48 B 0.0307f
C86 VP.n49 B 0.025455f
C87 VP.n50 B 0.0619f
C88 VP.n51 B 0.056088f
C89 VP.n52 B 0.0307f
C90 VP.n53 B 0.0307f
C91 VP.n54 B 0.030099f
C92 VP.n55 B 0.057218f
C93 VP.n56 B 0.061017f
C94 VP.n57 B 0.0307f
C95 VP.n58 B 0.0307f
C96 VP.n59 B 0.0307f
C97 VP.n60 B 0.061017f
C98 VP.n61 B 0.057218f
C99 VP.n62 B 0.030099f
C100 VP.n63 B 0.0307f
C101 VP.n64 B 0.0307f
C102 VP.n65 B 0.056088f
C103 VP.n66 B 0.0619f
C104 VP.n67 B 0.025455f
C105 VP.n68 B 0.0307f
C106 VP.n69 B 0.0307f
C107 VP.n70 B 0.0307f
C108 VP.n71 B 0.057218f
C109 VP.n72 B 0.032359f
C110 VP.n73 B 0.197878f
C111 VP.n74 B 0.056123f
C112 VTAIL.t9 B 0.02902f
C113 VTAIL.t12 B 0.02902f
C114 VTAIL.n0 B 0.093591f
C115 VTAIL.n1 B 0.562045f
C116 VTAIL.t15 B 0.160427f
C117 VTAIL.n2 B 0.625629f
C118 VTAIL.t7 B 0.160427f
C119 VTAIL.n3 B 0.625629f
C120 VTAIL.t1 B 0.02902f
C121 VTAIL.t6 B 0.02902f
C122 VTAIL.n4 B 0.093591f
C123 VTAIL.n5 B 0.88123f
C124 VTAIL.t0 B 0.160427f
C125 VTAIL.n6 B 1.52066f
C126 VTAIL.t11 B 0.160427f
C127 VTAIL.n7 B 1.52066f
C128 VTAIL.t8 B 0.02902f
C129 VTAIL.t14 B 0.02902f
C130 VTAIL.n8 B 0.093591f
C131 VTAIL.n9 B 0.88123f
C132 VTAIL.t10 B 0.160427f
C133 VTAIL.n10 B 0.625628f
C134 VTAIL.t3 B 0.160427f
C135 VTAIL.n11 B 0.625628f
C136 VTAIL.t5 B 0.02902f
C137 VTAIL.t4 B 0.02902f
C138 VTAIL.n12 B 0.093591f
C139 VTAIL.n13 B 0.88123f
C140 VTAIL.t2 B 0.160427f
C141 VTAIL.n14 B 1.52066f
C142 VTAIL.t13 B 0.160427f
C143 VTAIL.n15 B 1.51341f
C144 VDD2.t0 B 0.014435f
C145 VDD2.t1 B 0.014435f
C146 VDD2.n0 B 0.058019f
C147 VDD2.t2 B 0.014435f
C148 VDD2.t4 B 0.014435f
C149 VDD2.n1 B 0.058019f
C150 VDD2.n2 B 2.00954f
C151 VDD2.t5 B 0.014435f
C152 VDD2.t3 B 0.014435f
C153 VDD2.n3 B 0.056043f
C154 VDD2.n4 B 1.60654f
C155 VDD2.t6 B 0.014435f
C156 VDD2.t7 B 0.014435f
C157 VDD2.n5 B 0.058012f
C158 VN.n0 B 0.040266f
C159 VN.t2 B 0.143038f
C160 VN.n1 B 0.059189f
C161 VN.n2 B 0.030542f
C162 VN.t3 B 0.143038f
C163 VN.n3 B 0.101555f
C164 VN.n4 B 0.030542f
C165 VN.n5 B 0.02469f
C166 VN.n6 B 0.030542f
C167 VN.t6 B 0.143038f
C168 VN.n7 B 0.181413f
C169 VN.t0 B 0.372896f
C170 VN.n8 B 0.194682f
C171 VN.n9 B 0.298266f
C172 VN.n10 B 0.029943f
C173 VN.n11 B 0.056922f
C174 VN.n12 B 0.060701f
C175 VN.n13 B 0.030542f
C176 VN.n14 B 0.030542f
C177 VN.n15 B 0.030542f
C178 VN.n16 B 0.060701f
C179 VN.n17 B 0.056922f
C180 VN.n18 B 0.029943f
C181 VN.n19 B 0.030542f
C182 VN.n20 B 0.030542f
C183 VN.n21 B 0.055798f
C184 VN.n22 B 0.06158f
C185 VN.n23 B 0.025323f
C186 VN.n24 B 0.030542f
C187 VN.n25 B 0.030542f
C188 VN.n26 B 0.030542f
C189 VN.n27 B 0.056922f
C190 VN.n28 B 0.032192f
C191 VN.n29 B 0.196854f
C192 VN.n30 B 0.055833f
C193 VN.n31 B 0.040266f
C194 VN.t4 B 0.143038f
C195 VN.n32 B 0.059189f
C196 VN.n33 B 0.030542f
C197 VN.t7 B 0.143038f
C198 VN.n34 B 0.101555f
C199 VN.n35 B 0.030542f
C200 VN.n36 B 0.02469f
C201 VN.n37 B 0.030542f
C202 VN.t1 B 0.143038f
C203 VN.n38 B 0.181413f
C204 VN.t5 B 0.372896f
C205 VN.n39 B 0.194682f
C206 VN.n40 B 0.298266f
C207 VN.n41 B 0.029943f
C208 VN.n42 B 0.056922f
C209 VN.n43 B 0.060701f
C210 VN.n44 B 0.030542f
C211 VN.n45 B 0.030542f
C212 VN.n46 B 0.030542f
C213 VN.n47 B 0.060701f
C214 VN.n48 B 0.056922f
C215 VN.n49 B 0.029943f
C216 VN.n50 B 0.030542f
C217 VN.n51 B 0.030542f
C218 VN.n52 B 0.055798f
C219 VN.n53 B 0.06158f
C220 VN.n54 B 0.025323f
C221 VN.n55 B 0.030542f
C222 VN.n56 B 0.030542f
C223 VN.n57 B 0.030542f
C224 VN.n58 B 0.056922f
C225 VN.n59 B 0.032192f
C226 VN.n60 B 0.196854f
C227 VN.n61 B 1.37077f
.ends

