* NGSPICE file created from diff_pair_sample_1099.ext - technology: sky130A

.subckt diff_pair_sample_1099 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t14 VN.t0 VDD2.t4 B.t0 sky130_fd_pr__nfet_01v8 ad=0.91905 pd=5.9 as=0.91905 ps=5.9 w=5.57 l=1.61
X1 VDD2.t0 VN.t1 VTAIL.t13 B.t19 sky130_fd_pr__nfet_01v8 ad=0.91905 pd=5.9 as=0.91905 ps=5.9 w=5.57 l=1.61
X2 B.t18 B.t16 B.t17 B.t6 sky130_fd_pr__nfet_01v8 ad=2.1723 pd=11.92 as=0 ps=0 w=5.57 l=1.61
X3 VDD1.t7 VP.t0 VTAIL.t5 B.t19 sky130_fd_pr__nfet_01v8 ad=0.91905 pd=5.9 as=0.91905 ps=5.9 w=5.57 l=1.61
X4 VDD1.t6 VP.t1 VTAIL.t15 B.t21 sky130_fd_pr__nfet_01v8 ad=0.91905 pd=5.9 as=0.91905 ps=5.9 w=5.57 l=1.61
X5 VTAIL.t12 VN.t2 VDD2.t6 B.t20 sky130_fd_pr__nfet_01v8 ad=0.91905 pd=5.9 as=0.91905 ps=5.9 w=5.57 l=1.61
X6 VDD2.t2 VN.t3 VTAIL.t11 B.t21 sky130_fd_pr__nfet_01v8 ad=0.91905 pd=5.9 as=0.91905 ps=5.9 w=5.57 l=1.61
X7 VTAIL.t6 VP.t2 VDD1.t5 B.t20 sky130_fd_pr__nfet_01v8 ad=0.91905 pd=5.9 as=0.91905 ps=5.9 w=5.57 l=1.61
X8 VTAIL.t4 VP.t3 VDD1.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=2.1723 pd=11.92 as=0.91905 ps=5.9 w=5.57 l=1.61
X9 VTAIL.t2 VP.t4 VDD1.t3 B.t2 sky130_fd_pr__nfet_01v8 ad=2.1723 pd=11.92 as=0.91905 ps=5.9 w=5.57 l=1.61
X10 B.t15 B.t13 B.t14 B.t10 sky130_fd_pr__nfet_01v8 ad=2.1723 pd=11.92 as=0 ps=0 w=5.57 l=1.61
X11 VDD2.t5 VN.t4 VTAIL.t10 B.t3 sky130_fd_pr__nfet_01v8 ad=0.91905 pd=5.9 as=2.1723 ps=11.92 w=5.57 l=1.61
X12 VDD1.t2 VP.t5 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=0.91905 pd=5.9 as=2.1723 ps=11.92 w=5.57 l=1.61
X13 VDD2.t1 VN.t5 VTAIL.t9 B.t1 sky130_fd_pr__nfet_01v8 ad=0.91905 pd=5.9 as=2.1723 ps=11.92 w=5.57 l=1.61
X14 VTAIL.t0 VP.t6 VDD1.t1 B.t0 sky130_fd_pr__nfet_01v8 ad=0.91905 pd=5.9 as=0.91905 ps=5.9 w=5.57 l=1.61
X15 B.t12 B.t9 B.t11 B.t10 sky130_fd_pr__nfet_01v8 ad=2.1723 pd=11.92 as=0 ps=0 w=5.57 l=1.61
X16 B.t8 B.t5 B.t7 B.t6 sky130_fd_pr__nfet_01v8 ad=2.1723 pd=11.92 as=0 ps=0 w=5.57 l=1.61
X17 VTAIL.t8 VN.t6 VDD2.t7 B.t4 sky130_fd_pr__nfet_01v8 ad=2.1723 pd=11.92 as=0.91905 ps=5.9 w=5.57 l=1.61
X18 VTAIL.t7 VN.t7 VDD2.t3 B.t2 sky130_fd_pr__nfet_01v8 ad=2.1723 pd=11.92 as=0.91905 ps=5.9 w=5.57 l=1.61
X19 VDD1.t0 VP.t7 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=0.91905 pd=5.9 as=2.1723 ps=11.92 w=5.57 l=1.61
R0 VN.n20 VN.n19 177.939
R1 VN.n41 VN.n40 177.939
R2 VN.n39 VN.n21 161.3
R3 VN.n38 VN.n37 161.3
R4 VN.n36 VN.n22 161.3
R5 VN.n35 VN.n34 161.3
R6 VN.n32 VN.n23 161.3
R7 VN.n31 VN.n30 161.3
R8 VN.n29 VN.n24 161.3
R9 VN.n28 VN.n27 161.3
R10 VN.n18 VN.n0 161.3
R11 VN.n17 VN.n16 161.3
R12 VN.n15 VN.n1 161.3
R13 VN.n14 VN.n13 161.3
R14 VN.n11 VN.n2 161.3
R15 VN.n10 VN.n9 161.3
R16 VN.n8 VN.n3 161.3
R17 VN.n7 VN.n6 161.3
R18 VN.n4 VN.t7 115.96
R19 VN.n25 VN.t5 115.96
R20 VN.n5 VN.t3 83.3775
R21 VN.n12 VN.t0 83.3775
R22 VN.n19 VN.t4 83.3775
R23 VN.n26 VN.t2 83.3775
R24 VN.n33 VN.t1 83.3775
R25 VN.n40 VN.t6 83.3775
R26 VN.n10 VN.n3 56.5193
R27 VN.n17 VN.n1 56.5193
R28 VN.n31 VN.n24 56.5193
R29 VN.n38 VN.n22 56.5193
R30 VN.n5 VN.n4 55.3922
R31 VN.n26 VN.n25 55.3922
R32 VN VN.n41 41.6918
R33 VN.n6 VN.n3 24.4675
R34 VN.n11 VN.n10 24.4675
R35 VN.n13 VN.n1 24.4675
R36 VN.n18 VN.n17 24.4675
R37 VN.n27 VN.n24 24.4675
R38 VN.n34 VN.n22 24.4675
R39 VN.n32 VN.n31 24.4675
R40 VN.n39 VN.n38 24.4675
R41 VN.n28 VN.n25 17.9992
R42 VN.n7 VN.n4 17.9992
R43 VN.n13 VN.n12 13.702
R44 VN.n34 VN.n33 13.702
R45 VN.n6 VN.n5 10.766
R46 VN.n12 VN.n11 10.766
R47 VN.n27 VN.n26 10.766
R48 VN.n33 VN.n32 10.766
R49 VN.n19 VN.n18 7.82994
R50 VN.n40 VN.n39 7.82994
R51 VN.n41 VN.n21 0.189894
R52 VN.n37 VN.n21 0.189894
R53 VN.n37 VN.n36 0.189894
R54 VN.n36 VN.n35 0.189894
R55 VN.n35 VN.n23 0.189894
R56 VN.n30 VN.n23 0.189894
R57 VN.n30 VN.n29 0.189894
R58 VN.n29 VN.n28 0.189894
R59 VN.n8 VN.n7 0.189894
R60 VN.n9 VN.n8 0.189894
R61 VN.n9 VN.n2 0.189894
R62 VN.n14 VN.n2 0.189894
R63 VN.n15 VN.n14 0.189894
R64 VN.n16 VN.n15 0.189894
R65 VN.n16 VN.n0 0.189894
R66 VN.n20 VN.n0 0.189894
R67 VN VN.n20 0.0516364
R68 VDD2.n2 VDD2.n1 67.2931
R69 VDD2.n2 VDD2.n0 67.2931
R70 VDD2 VDD2.n5 67.2903
R71 VDD2.n4 VDD2.n3 66.5124
R72 VDD2.n4 VDD2.n2 36.0429
R73 VDD2.n5 VDD2.t6 3.55526
R74 VDD2.n5 VDD2.t1 3.55526
R75 VDD2.n3 VDD2.t7 3.55526
R76 VDD2.n3 VDD2.t0 3.55526
R77 VDD2.n1 VDD2.t4 3.55526
R78 VDD2.n1 VDD2.t5 3.55526
R79 VDD2.n0 VDD2.t3 3.55526
R80 VDD2.n0 VDD2.t2 3.55526
R81 VDD2 VDD2.n4 0.894897
R82 VTAIL.n11 VTAIL.t2 53.3884
R83 VTAIL.n10 VTAIL.t9 53.3884
R84 VTAIL.n7 VTAIL.t8 53.3884
R85 VTAIL.n15 VTAIL.t10 53.3882
R86 VTAIL.n2 VTAIL.t7 53.3882
R87 VTAIL.n3 VTAIL.t1 53.3882
R88 VTAIL.n6 VTAIL.t4 53.3882
R89 VTAIL.n14 VTAIL.t3 53.3882
R90 VTAIL.n13 VTAIL.n12 49.8337
R91 VTAIL.n9 VTAIL.n8 49.8337
R92 VTAIL.n1 VTAIL.n0 49.8334
R93 VTAIL.n5 VTAIL.n4 49.8334
R94 VTAIL.n15 VTAIL.n14 18.841
R95 VTAIL.n7 VTAIL.n6 18.841
R96 VTAIL.n0 VTAIL.t11 3.55526
R97 VTAIL.n0 VTAIL.t14 3.55526
R98 VTAIL.n4 VTAIL.t5 3.55526
R99 VTAIL.n4 VTAIL.t6 3.55526
R100 VTAIL.n12 VTAIL.t15 3.55526
R101 VTAIL.n12 VTAIL.t0 3.55526
R102 VTAIL.n8 VTAIL.t13 3.55526
R103 VTAIL.n8 VTAIL.t12 3.55526
R104 VTAIL.n9 VTAIL.n7 1.67291
R105 VTAIL.n10 VTAIL.n9 1.67291
R106 VTAIL.n13 VTAIL.n11 1.67291
R107 VTAIL.n14 VTAIL.n13 1.67291
R108 VTAIL.n6 VTAIL.n5 1.67291
R109 VTAIL.n5 VTAIL.n3 1.67291
R110 VTAIL.n2 VTAIL.n1 1.67291
R111 VTAIL VTAIL.n15 1.61472
R112 VTAIL.n11 VTAIL.n10 0.470328
R113 VTAIL.n3 VTAIL.n2 0.470328
R114 VTAIL VTAIL.n1 0.0586897
R115 B.n579 B.n578 585
R116 B.n580 B.n579 585
R117 B.n207 B.n96 585
R118 B.n206 B.n205 585
R119 B.n204 B.n203 585
R120 B.n202 B.n201 585
R121 B.n200 B.n199 585
R122 B.n198 B.n197 585
R123 B.n196 B.n195 585
R124 B.n194 B.n193 585
R125 B.n192 B.n191 585
R126 B.n190 B.n189 585
R127 B.n188 B.n187 585
R128 B.n186 B.n185 585
R129 B.n184 B.n183 585
R130 B.n182 B.n181 585
R131 B.n180 B.n179 585
R132 B.n178 B.n177 585
R133 B.n176 B.n175 585
R134 B.n174 B.n173 585
R135 B.n172 B.n171 585
R136 B.n170 B.n169 585
R137 B.n168 B.n167 585
R138 B.n166 B.n165 585
R139 B.n164 B.n163 585
R140 B.n162 B.n161 585
R141 B.n160 B.n159 585
R142 B.n158 B.n157 585
R143 B.n156 B.n155 585
R144 B.n154 B.n153 585
R145 B.n152 B.n151 585
R146 B.n150 B.n149 585
R147 B.n148 B.n147 585
R148 B.n145 B.n144 585
R149 B.n143 B.n142 585
R150 B.n141 B.n140 585
R151 B.n139 B.n138 585
R152 B.n137 B.n136 585
R153 B.n135 B.n134 585
R154 B.n133 B.n132 585
R155 B.n131 B.n130 585
R156 B.n129 B.n128 585
R157 B.n127 B.n126 585
R158 B.n125 B.n124 585
R159 B.n123 B.n122 585
R160 B.n121 B.n120 585
R161 B.n119 B.n118 585
R162 B.n117 B.n116 585
R163 B.n115 B.n114 585
R164 B.n113 B.n112 585
R165 B.n111 B.n110 585
R166 B.n109 B.n108 585
R167 B.n107 B.n106 585
R168 B.n105 B.n104 585
R169 B.n103 B.n102 585
R170 B.n67 B.n66 585
R171 B.n577 B.n68 585
R172 B.n581 B.n68 585
R173 B.n576 B.n575 585
R174 B.n575 B.n64 585
R175 B.n574 B.n63 585
R176 B.n587 B.n63 585
R177 B.n573 B.n62 585
R178 B.n588 B.n62 585
R179 B.n572 B.n61 585
R180 B.n589 B.n61 585
R181 B.n571 B.n570 585
R182 B.n570 B.n57 585
R183 B.n569 B.n56 585
R184 B.n595 B.n56 585
R185 B.n568 B.n55 585
R186 B.n596 B.n55 585
R187 B.n567 B.n54 585
R188 B.n597 B.n54 585
R189 B.n566 B.n565 585
R190 B.n565 B.n50 585
R191 B.n564 B.n49 585
R192 B.n603 B.n49 585
R193 B.n563 B.n48 585
R194 B.n604 B.n48 585
R195 B.n562 B.n47 585
R196 B.n605 B.n47 585
R197 B.n561 B.n560 585
R198 B.n560 B.n43 585
R199 B.n559 B.n42 585
R200 B.n611 B.n42 585
R201 B.n558 B.n41 585
R202 B.n612 B.n41 585
R203 B.n557 B.n40 585
R204 B.n613 B.n40 585
R205 B.n556 B.n555 585
R206 B.n555 B.n36 585
R207 B.n554 B.n35 585
R208 B.n619 B.n35 585
R209 B.n553 B.n34 585
R210 B.n620 B.n34 585
R211 B.n552 B.n33 585
R212 B.n621 B.n33 585
R213 B.n551 B.n550 585
R214 B.n550 B.n29 585
R215 B.n549 B.n28 585
R216 B.n627 B.n28 585
R217 B.n548 B.n27 585
R218 B.n628 B.n27 585
R219 B.n547 B.n26 585
R220 B.n629 B.n26 585
R221 B.n546 B.n545 585
R222 B.n545 B.n22 585
R223 B.n544 B.n21 585
R224 B.n635 B.n21 585
R225 B.n543 B.n20 585
R226 B.n636 B.n20 585
R227 B.n542 B.n19 585
R228 B.n637 B.n19 585
R229 B.n541 B.n540 585
R230 B.n540 B.n15 585
R231 B.n539 B.n14 585
R232 B.n643 B.n14 585
R233 B.n538 B.n13 585
R234 B.n644 B.n13 585
R235 B.n537 B.n12 585
R236 B.n645 B.n12 585
R237 B.n536 B.n535 585
R238 B.n535 B.n534 585
R239 B.n533 B.n532 585
R240 B.n533 B.n8 585
R241 B.n531 B.n7 585
R242 B.n652 B.n7 585
R243 B.n530 B.n6 585
R244 B.n653 B.n6 585
R245 B.n529 B.n5 585
R246 B.n654 B.n5 585
R247 B.n528 B.n527 585
R248 B.n527 B.n4 585
R249 B.n526 B.n208 585
R250 B.n526 B.n525 585
R251 B.n516 B.n209 585
R252 B.n210 B.n209 585
R253 B.n518 B.n517 585
R254 B.n519 B.n518 585
R255 B.n515 B.n215 585
R256 B.n215 B.n214 585
R257 B.n514 B.n513 585
R258 B.n513 B.n512 585
R259 B.n217 B.n216 585
R260 B.n218 B.n217 585
R261 B.n505 B.n504 585
R262 B.n506 B.n505 585
R263 B.n503 B.n223 585
R264 B.n223 B.n222 585
R265 B.n502 B.n501 585
R266 B.n501 B.n500 585
R267 B.n225 B.n224 585
R268 B.n226 B.n225 585
R269 B.n493 B.n492 585
R270 B.n494 B.n493 585
R271 B.n491 B.n231 585
R272 B.n231 B.n230 585
R273 B.n490 B.n489 585
R274 B.n489 B.n488 585
R275 B.n233 B.n232 585
R276 B.n234 B.n233 585
R277 B.n481 B.n480 585
R278 B.n482 B.n481 585
R279 B.n479 B.n239 585
R280 B.n239 B.n238 585
R281 B.n478 B.n477 585
R282 B.n477 B.n476 585
R283 B.n241 B.n240 585
R284 B.n242 B.n241 585
R285 B.n469 B.n468 585
R286 B.n470 B.n469 585
R287 B.n467 B.n247 585
R288 B.n247 B.n246 585
R289 B.n466 B.n465 585
R290 B.n465 B.n464 585
R291 B.n249 B.n248 585
R292 B.n250 B.n249 585
R293 B.n457 B.n456 585
R294 B.n458 B.n457 585
R295 B.n455 B.n255 585
R296 B.n255 B.n254 585
R297 B.n454 B.n453 585
R298 B.n453 B.n452 585
R299 B.n257 B.n256 585
R300 B.n258 B.n257 585
R301 B.n445 B.n444 585
R302 B.n446 B.n445 585
R303 B.n443 B.n263 585
R304 B.n263 B.n262 585
R305 B.n442 B.n441 585
R306 B.n441 B.n440 585
R307 B.n265 B.n264 585
R308 B.n266 B.n265 585
R309 B.n433 B.n432 585
R310 B.n434 B.n433 585
R311 B.n431 B.n271 585
R312 B.n271 B.n270 585
R313 B.n430 B.n429 585
R314 B.n429 B.n428 585
R315 B.n273 B.n272 585
R316 B.n274 B.n273 585
R317 B.n421 B.n420 585
R318 B.n422 B.n421 585
R319 B.n277 B.n276 585
R320 B.n310 B.n309 585
R321 B.n311 B.n307 585
R322 B.n307 B.n278 585
R323 B.n313 B.n312 585
R324 B.n315 B.n306 585
R325 B.n318 B.n317 585
R326 B.n319 B.n305 585
R327 B.n321 B.n320 585
R328 B.n323 B.n304 585
R329 B.n326 B.n325 585
R330 B.n327 B.n303 585
R331 B.n329 B.n328 585
R332 B.n331 B.n302 585
R333 B.n334 B.n333 585
R334 B.n335 B.n301 585
R335 B.n337 B.n336 585
R336 B.n339 B.n300 585
R337 B.n342 B.n341 585
R338 B.n343 B.n299 585
R339 B.n345 B.n344 585
R340 B.n347 B.n298 585
R341 B.n350 B.n349 585
R342 B.n351 B.n295 585
R343 B.n354 B.n353 585
R344 B.n356 B.n294 585
R345 B.n359 B.n358 585
R346 B.n360 B.n293 585
R347 B.n362 B.n361 585
R348 B.n364 B.n292 585
R349 B.n367 B.n366 585
R350 B.n368 B.n291 585
R351 B.n373 B.n372 585
R352 B.n375 B.n290 585
R353 B.n378 B.n377 585
R354 B.n379 B.n289 585
R355 B.n381 B.n380 585
R356 B.n383 B.n288 585
R357 B.n386 B.n385 585
R358 B.n387 B.n287 585
R359 B.n389 B.n388 585
R360 B.n391 B.n286 585
R361 B.n394 B.n393 585
R362 B.n395 B.n285 585
R363 B.n397 B.n396 585
R364 B.n399 B.n284 585
R365 B.n402 B.n401 585
R366 B.n403 B.n283 585
R367 B.n405 B.n404 585
R368 B.n407 B.n282 585
R369 B.n410 B.n409 585
R370 B.n411 B.n281 585
R371 B.n413 B.n412 585
R372 B.n415 B.n280 585
R373 B.n418 B.n417 585
R374 B.n419 B.n279 585
R375 B.n424 B.n423 585
R376 B.n423 B.n422 585
R377 B.n425 B.n275 585
R378 B.n275 B.n274 585
R379 B.n427 B.n426 585
R380 B.n428 B.n427 585
R381 B.n269 B.n268 585
R382 B.n270 B.n269 585
R383 B.n436 B.n435 585
R384 B.n435 B.n434 585
R385 B.n437 B.n267 585
R386 B.n267 B.n266 585
R387 B.n439 B.n438 585
R388 B.n440 B.n439 585
R389 B.n261 B.n260 585
R390 B.n262 B.n261 585
R391 B.n448 B.n447 585
R392 B.n447 B.n446 585
R393 B.n449 B.n259 585
R394 B.n259 B.n258 585
R395 B.n451 B.n450 585
R396 B.n452 B.n451 585
R397 B.n253 B.n252 585
R398 B.n254 B.n253 585
R399 B.n460 B.n459 585
R400 B.n459 B.n458 585
R401 B.n461 B.n251 585
R402 B.n251 B.n250 585
R403 B.n463 B.n462 585
R404 B.n464 B.n463 585
R405 B.n245 B.n244 585
R406 B.n246 B.n245 585
R407 B.n472 B.n471 585
R408 B.n471 B.n470 585
R409 B.n473 B.n243 585
R410 B.n243 B.n242 585
R411 B.n475 B.n474 585
R412 B.n476 B.n475 585
R413 B.n237 B.n236 585
R414 B.n238 B.n237 585
R415 B.n484 B.n483 585
R416 B.n483 B.n482 585
R417 B.n485 B.n235 585
R418 B.n235 B.n234 585
R419 B.n487 B.n486 585
R420 B.n488 B.n487 585
R421 B.n229 B.n228 585
R422 B.n230 B.n229 585
R423 B.n496 B.n495 585
R424 B.n495 B.n494 585
R425 B.n497 B.n227 585
R426 B.n227 B.n226 585
R427 B.n499 B.n498 585
R428 B.n500 B.n499 585
R429 B.n221 B.n220 585
R430 B.n222 B.n221 585
R431 B.n508 B.n507 585
R432 B.n507 B.n506 585
R433 B.n509 B.n219 585
R434 B.n219 B.n218 585
R435 B.n511 B.n510 585
R436 B.n512 B.n511 585
R437 B.n213 B.n212 585
R438 B.n214 B.n213 585
R439 B.n521 B.n520 585
R440 B.n520 B.n519 585
R441 B.n522 B.n211 585
R442 B.n211 B.n210 585
R443 B.n524 B.n523 585
R444 B.n525 B.n524 585
R445 B.n3 B.n0 585
R446 B.n4 B.n3 585
R447 B.n651 B.n1 585
R448 B.n652 B.n651 585
R449 B.n650 B.n649 585
R450 B.n650 B.n8 585
R451 B.n648 B.n9 585
R452 B.n534 B.n9 585
R453 B.n647 B.n646 585
R454 B.n646 B.n645 585
R455 B.n11 B.n10 585
R456 B.n644 B.n11 585
R457 B.n642 B.n641 585
R458 B.n643 B.n642 585
R459 B.n640 B.n16 585
R460 B.n16 B.n15 585
R461 B.n639 B.n638 585
R462 B.n638 B.n637 585
R463 B.n18 B.n17 585
R464 B.n636 B.n18 585
R465 B.n634 B.n633 585
R466 B.n635 B.n634 585
R467 B.n632 B.n23 585
R468 B.n23 B.n22 585
R469 B.n631 B.n630 585
R470 B.n630 B.n629 585
R471 B.n25 B.n24 585
R472 B.n628 B.n25 585
R473 B.n626 B.n625 585
R474 B.n627 B.n626 585
R475 B.n624 B.n30 585
R476 B.n30 B.n29 585
R477 B.n623 B.n622 585
R478 B.n622 B.n621 585
R479 B.n32 B.n31 585
R480 B.n620 B.n32 585
R481 B.n618 B.n617 585
R482 B.n619 B.n618 585
R483 B.n616 B.n37 585
R484 B.n37 B.n36 585
R485 B.n615 B.n614 585
R486 B.n614 B.n613 585
R487 B.n39 B.n38 585
R488 B.n612 B.n39 585
R489 B.n610 B.n609 585
R490 B.n611 B.n610 585
R491 B.n608 B.n44 585
R492 B.n44 B.n43 585
R493 B.n607 B.n606 585
R494 B.n606 B.n605 585
R495 B.n46 B.n45 585
R496 B.n604 B.n46 585
R497 B.n602 B.n601 585
R498 B.n603 B.n602 585
R499 B.n600 B.n51 585
R500 B.n51 B.n50 585
R501 B.n599 B.n598 585
R502 B.n598 B.n597 585
R503 B.n53 B.n52 585
R504 B.n596 B.n53 585
R505 B.n594 B.n593 585
R506 B.n595 B.n594 585
R507 B.n592 B.n58 585
R508 B.n58 B.n57 585
R509 B.n591 B.n590 585
R510 B.n590 B.n589 585
R511 B.n60 B.n59 585
R512 B.n588 B.n60 585
R513 B.n586 B.n585 585
R514 B.n587 B.n586 585
R515 B.n584 B.n65 585
R516 B.n65 B.n64 585
R517 B.n583 B.n582 585
R518 B.n582 B.n581 585
R519 B.n655 B.n654 585
R520 B.n653 B.n2 585
R521 B.n582 B.n67 521.33
R522 B.n579 B.n68 521.33
R523 B.n421 B.n279 521.33
R524 B.n423 B.n277 521.33
R525 B.n100 B.t13 289.204
R526 B.n97 B.t9 289.204
R527 B.n369 B.t5 289.204
R528 B.n296 B.t16 289.204
R529 B.n580 B.n95 256.663
R530 B.n580 B.n94 256.663
R531 B.n580 B.n93 256.663
R532 B.n580 B.n92 256.663
R533 B.n580 B.n91 256.663
R534 B.n580 B.n90 256.663
R535 B.n580 B.n89 256.663
R536 B.n580 B.n88 256.663
R537 B.n580 B.n87 256.663
R538 B.n580 B.n86 256.663
R539 B.n580 B.n85 256.663
R540 B.n580 B.n84 256.663
R541 B.n580 B.n83 256.663
R542 B.n580 B.n82 256.663
R543 B.n580 B.n81 256.663
R544 B.n580 B.n80 256.663
R545 B.n580 B.n79 256.663
R546 B.n580 B.n78 256.663
R547 B.n580 B.n77 256.663
R548 B.n580 B.n76 256.663
R549 B.n580 B.n75 256.663
R550 B.n580 B.n74 256.663
R551 B.n580 B.n73 256.663
R552 B.n580 B.n72 256.663
R553 B.n580 B.n71 256.663
R554 B.n580 B.n70 256.663
R555 B.n580 B.n69 256.663
R556 B.n308 B.n278 256.663
R557 B.n314 B.n278 256.663
R558 B.n316 B.n278 256.663
R559 B.n322 B.n278 256.663
R560 B.n324 B.n278 256.663
R561 B.n330 B.n278 256.663
R562 B.n332 B.n278 256.663
R563 B.n338 B.n278 256.663
R564 B.n340 B.n278 256.663
R565 B.n346 B.n278 256.663
R566 B.n348 B.n278 256.663
R567 B.n355 B.n278 256.663
R568 B.n357 B.n278 256.663
R569 B.n363 B.n278 256.663
R570 B.n365 B.n278 256.663
R571 B.n374 B.n278 256.663
R572 B.n376 B.n278 256.663
R573 B.n382 B.n278 256.663
R574 B.n384 B.n278 256.663
R575 B.n390 B.n278 256.663
R576 B.n392 B.n278 256.663
R577 B.n398 B.n278 256.663
R578 B.n400 B.n278 256.663
R579 B.n406 B.n278 256.663
R580 B.n408 B.n278 256.663
R581 B.n414 B.n278 256.663
R582 B.n416 B.n278 256.663
R583 B.n657 B.n656 256.663
R584 B.n104 B.n103 163.367
R585 B.n108 B.n107 163.367
R586 B.n112 B.n111 163.367
R587 B.n116 B.n115 163.367
R588 B.n120 B.n119 163.367
R589 B.n124 B.n123 163.367
R590 B.n128 B.n127 163.367
R591 B.n132 B.n131 163.367
R592 B.n136 B.n135 163.367
R593 B.n140 B.n139 163.367
R594 B.n144 B.n143 163.367
R595 B.n149 B.n148 163.367
R596 B.n153 B.n152 163.367
R597 B.n157 B.n156 163.367
R598 B.n161 B.n160 163.367
R599 B.n165 B.n164 163.367
R600 B.n169 B.n168 163.367
R601 B.n173 B.n172 163.367
R602 B.n177 B.n176 163.367
R603 B.n181 B.n180 163.367
R604 B.n185 B.n184 163.367
R605 B.n189 B.n188 163.367
R606 B.n193 B.n192 163.367
R607 B.n197 B.n196 163.367
R608 B.n201 B.n200 163.367
R609 B.n205 B.n204 163.367
R610 B.n579 B.n96 163.367
R611 B.n421 B.n273 163.367
R612 B.n429 B.n273 163.367
R613 B.n429 B.n271 163.367
R614 B.n433 B.n271 163.367
R615 B.n433 B.n265 163.367
R616 B.n441 B.n265 163.367
R617 B.n441 B.n263 163.367
R618 B.n445 B.n263 163.367
R619 B.n445 B.n257 163.367
R620 B.n453 B.n257 163.367
R621 B.n453 B.n255 163.367
R622 B.n457 B.n255 163.367
R623 B.n457 B.n249 163.367
R624 B.n465 B.n249 163.367
R625 B.n465 B.n247 163.367
R626 B.n469 B.n247 163.367
R627 B.n469 B.n241 163.367
R628 B.n477 B.n241 163.367
R629 B.n477 B.n239 163.367
R630 B.n481 B.n239 163.367
R631 B.n481 B.n233 163.367
R632 B.n489 B.n233 163.367
R633 B.n489 B.n231 163.367
R634 B.n493 B.n231 163.367
R635 B.n493 B.n225 163.367
R636 B.n501 B.n225 163.367
R637 B.n501 B.n223 163.367
R638 B.n505 B.n223 163.367
R639 B.n505 B.n217 163.367
R640 B.n513 B.n217 163.367
R641 B.n513 B.n215 163.367
R642 B.n518 B.n215 163.367
R643 B.n518 B.n209 163.367
R644 B.n526 B.n209 163.367
R645 B.n527 B.n526 163.367
R646 B.n527 B.n5 163.367
R647 B.n6 B.n5 163.367
R648 B.n7 B.n6 163.367
R649 B.n533 B.n7 163.367
R650 B.n535 B.n533 163.367
R651 B.n535 B.n12 163.367
R652 B.n13 B.n12 163.367
R653 B.n14 B.n13 163.367
R654 B.n540 B.n14 163.367
R655 B.n540 B.n19 163.367
R656 B.n20 B.n19 163.367
R657 B.n21 B.n20 163.367
R658 B.n545 B.n21 163.367
R659 B.n545 B.n26 163.367
R660 B.n27 B.n26 163.367
R661 B.n28 B.n27 163.367
R662 B.n550 B.n28 163.367
R663 B.n550 B.n33 163.367
R664 B.n34 B.n33 163.367
R665 B.n35 B.n34 163.367
R666 B.n555 B.n35 163.367
R667 B.n555 B.n40 163.367
R668 B.n41 B.n40 163.367
R669 B.n42 B.n41 163.367
R670 B.n560 B.n42 163.367
R671 B.n560 B.n47 163.367
R672 B.n48 B.n47 163.367
R673 B.n49 B.n48 163.367
R674 B.n565 B.n49 163.367
R675 B.n565 B.n54 163.367
R676 B.n55 B.n54 163.367
R677 B.n56 B.n55 163.367
R678 B.n570 B.n56 163.367
R679 B.n570 B.n61 163.367
R680 B.n62 B.n61 163.367
R681 B.n63 B.n62 163.367
R682 B.n575 B.n63 163.367
R683 B.n575 B.n68 163.367
R684 B.n309 B.n307 163.367
R685 B.n313 B.n307 163.367
R686 B.n317 B.n315 163.367
R687 B.n321 B.n305 163.367
R688 B.n325 B.n323 163.367
R689 B.n329 B.n303 163.367
R690 B.n333 B.n331 163.367
R691 B.n337 B.n301 163.367
R692 B.n341 B.n339 163.367
R693 B.n345 B.n299 163.367
R694 B.n349 B.n347 163.367
R695 B.n354 B.n295 163.367
R696 B.n358 B.n356 163.367
R697 B.n362 B.n293 163.367
R698 B.n366 B.n364 163.367
R699 B.n373 B.n291 163.367
R700 B.n377 B.n375 163.367
R701 B.n381 B.n289 163.367
R702 B.n385 B.n383 163.367
R703 B.n389 B.n287 163.367
R704 B.n393 B.n391 163.367
R705 B.n397 B.n285 163.367
R706 B.n401 B.n399 163.367
R707 B.n405 B.n283 163.367
R708 B.n409 B.n407 163.367
R709 B.n413 B.n281 163.367
R710 B.n417 B.n415 163.367
R711 B.n423 B.n275 163.367
R712 B.n427 B.n275 163.367
R713 B.n427 B.n269 163.367
R714 B.n435 B.n269 163.367
R715 B.n435 B.n267 163.367
R716 B.n439 B.n267 163.367
R717 B.n439 B.n261 163.367
R718 B.n447 B.n261 163.367
R719 B.n447 B.n259 163.367
R720 B.n451 B.n259 163.367
R721 B.n451 B.n253 163.367
R722 B.n459 B.n253 163.367
R723 B.n459 B.n251 163.367
R724 B.n463 B.n251 163.367
R725 B.n463 B.n245 163.367
R726 B.n471 B.n245 163.367
R727 B.n471 B.n243 163.367
R728 B.n475 B.n243 163.367
R729 B.n475 B.n237 163.367
R730 B.n483 B.n237 163.367
R731 B.n483 B.n235 163.367
R732 B.n487 B.n235 163.367
R733 B.n487 B.n229 163.367
R734 B.n495 B.n229 163.367
R735 B.n495 B.n227 163.367
R736 B.n499 B.n227 163.367
R737 B.n499 B.n221 163.367
R738 B.n507 B.n221 163.367
R739 B.n507 B.n219 163.367
R740 B.n511 B.n219 163.367
R741 B.n511 B.n213 163.367
R742 B.n520 B.n213 163.367
R743 B.n520 B.n211 163.367
R744 B.n524 B.n211 163.367
R745 B.n524 B.n3 163.367
R746 B.n655 B.n3 163.367
R747 B.n651 B.n2 163.367
R748 B.n651 B.n650 163.367
R749 B.n650 B.n9 163.367
R750 B.n646 B.n9 163.367
R751 B.n646 B.n11 163.367
R752 B.n642 B.n11 163.367
R753 B.n642 B.n16 163.367
R754 B.n638 B.n16 163.367
R755 B.n638 B.n18 163.367
R756 B.n634 B.n18 163.367
R757 B.n634 B.n23 163.367
R758 B.n630 B.n23 163.367
R759 B.n630 B.n25 163.367
R760 B.n626 B.n25 163.367
R761 B.n626 B.n30 163.367
R762 B.n622 B.n30 163.367
R763 B.n622 B.n32 163.367
R764 B.n618 B.n32 163.367
R765 B.n618 B.n37 163.367
R766 B.n614 B.n37 163.367
R767 B.n614 B.n39 163.367
R768 B.n610 B.n39 163.367
R769 B.n610 B.n44 163.367
R770 B.n606 B.n44 163.367
R771 B.n606 B.n46 163.367
R772 B.n602 B.n46 163.367
R773 B.n602 B.n51 163.367
R774 B.n598 B.n51 163.367
R775 B.n598 B.n53 163.367
R776 B.n594 B.n53 163.367
R777 B.n594 B.n58 163.367
R778 B.n590 B.n58 163.367
R779 B.n590 B.n60 163.367
R780 B.n586 B.n60 163.367
R781 B.n586 B.n65 163.367
R782 B.n582 B.n65 163.367
R783 B.n422 B.n278 134.901
R784 B.n581 B.n580 134.901
R785 B.n97 B.t11 109.865
R786 B.n369 B.t8 109.865
R787 B.n100 B.t14 109.859
R788 B.n296 B.t18 109.859
R789 B.n98 B.t12 72.2403
R790 B.n370 B.t7 72.2403
R791 B.n101 B.t15 72.2345
R792 B.n297 B.t17 72.2345
R793 B.n69 B.n67 71.676
R794 B.n104 B.n70 71.676
R795 B.n108 B.n71 71.676
R796 B.n112 B.n72 71.676
R797 B.n116 B.n73 71.676
R798 B.n120 B.n74 71.676
R799 B.n124 B.n75 71.676
R800 B.n128 B.n76 71.676
R801 B.n132 B.n77 71.676
R802 B.n136 B.n78 71.676
R803 B.n140 B.n79 71.676
R804 B.n144 B.n80 71.676
R805 B.n149 B.n81 71.676
R806 B.n153 B.n82 71.676
R807 B.n157 B.n83 71.676
R808 B.n161 B.n84 71.676
R809 B.n165 B.n85 71.676
R810 B.n169 B.n86 71.676
R811 B.n173 B.n87 71.676
R812 B.n177 B.n88 71.676
R813 B.n181 B.n89 71.676
R814 B.n185 B.n90 71.676
R815 B.n189 B.n91 71.676
R816 B.n193 B.n92 71.676
R817 B.n197 B.n93 71.676
R818 B.n201 B.n94 71.676
R819 B.n205 B.n95 71.676
R820 B.n96 B.n95 71.676
R821 B.n204 B.n94 71.676
R822 B.n200 B.n93 71.676
R823 B.n196 B.n92 71.676
R824 B.n192 B.n91 71.676
R825 B.n188 B.n90 71.676
R826 B.n184 B.n89 71.676
R827 B.n180 B.n88 71.676
R828 B.n176 B.n87 71.676
R829 B.n172 B.n86 71.676
R830 B.n168 B.n85 71.676
R831 B.n164 B.n84 71.676
R832 B.n160 B.n83 71.676
R833 B.n156 B.n82 71.676
R834 B.n152 B.n81 71.676
R835 B.n148 B.n80 71.676
R836 B.n143 B.n79 71.676
R837 B.n139 B.n78 71.676
R838 B.n135 B.n77 71.676
R839 B.n131 B.n76 71.676
R840 B.n127 B.n75 71.676
R841 B.n123 B.n74 71.676
R842 B.n119 B.n73 71.676
R843 B.n115 B.n72 71.676
R844 B.n111 B.n71 71.676
R845 B.n107 B.n70 71.676
R846 B.n103 B.n69 71.676
R847 B.n308 B.n277 71.676
R848 B.n314 B.n313 71.676
R849 B.n317 B.n316 71.676
R850 B.n322 B.n321 71.676
R851 B.n325 B.n324 71.676
R852 B.n330 B.n329 71.676
R853 B.n333 B.n332 71.676
R854 B.n338 B.n337 71.676
R855 B.n341 B.n340 71.676
R856 B.n346 B.n345 71.676
R857 B.n349 B.n348 71.676
R858 B.n355 B.n354 71.676
R859 B.n358 B.n357 71.676
R860 B.n363 B.n362 71.676
R861 B.n366 B.n365 71.676
R862 B.n374 B.n373 71.676
R863 B.n377 B.n376 71.676
R864 B.n382 B.n381 71.676
R865 B.n385 B.n384 71.676
R866 B.n390 B.n389 71.676
R867 B.n393 B.n392 71.676
R868 B.n398 B.n397 71.676
R869 B.n401 B.n400 71.676
R870 B.n406 B.n405 71.676
R871 B.n409 B.n408 71.676
R872 B.n414 B.n413 71.676
R873 B.n417 B.n416 71.676
R874 B.n309 B.n308 71.676
R875 B.n315 B.n314 71.676
R876 B.n316 B.n305 71.676
R877 B.n323 B.n322 71.676
R878 B.n324 B.n303 71.676
R879 B.n331 B.n330 71.676
R880 B.n332 B.n301 71.676
R881 B.n339 B.n338 71.676
R882 B.n340 B.n299 71.676
R883 B.n347 B.n346 71.676
R884 B.n348 B.n295 71.676
R885 B.n356 B.n355 71.676
R886 B.n357 B.n293 71.676
R887 B.n364 B.n363 71.676
R888 B.n365 B.n291 71.676
R889 B.n375 B.n374 71.676
R890 B.n376 B.n289 71.676
R891 B.n383 B.n382 71.676
R892 B.n384 B.n287 71.676
R893 B.n391 B.n390 71.676
R894 B.n392 B.n285 71.676
R895 B.n399 B.n398 71.676
R896 B.n400 B.n283 71.676
R897 B.n407 B.n406 71.676
R898 B.n408 B.n281 71.676
R899 B.n415 B.n414 71.676
R900 B.n416 B.n279 71.676
R901 B.n656 B.n655 71.676
R902 B.n656 B.n2 71.676
R903 B.n422 B.n274 68.9724
R904 B.n428 B.n274 68.9724
R905 B.n428 B.n270 68.9724
R906 B.n434 B.n270 68.9724
R907 B.n434 B.n266 68.9724
R908 B.n440 B.n266 68.9724
R909 B.n446 B.n262 68.9724
R910 B.n446 B.n258 68.9724
R911 B.n452 B.n258 68.9724
R912 B.n452 B.n254 68.9724
R913 B.n458 B.n254 68.9724
R914 B.n458 B.n250 68.9724
R915 B.n464 B.n250 68.9724
R916 B.n470 B.n246 68.9724
R917 B.n470 B.n242 68.9724
R918 B.n476 B.n242 68.9724
R919 B.n476 B.n238 68.9724
R920 B.n482 B.n238 68.9724
R921 B.n488 B.n234 68.9724
R922 B.n488 B.n230 68.9724
R923 B.n494 B.n230 68.9724
R924 B.n494 B.n226 68.9724
R925 B.n500 B.n226 68.9724
R926 B.n506 B.n222 68.9724
R927 B.n506 B.n218 68.9724
R928 B.n512 B.n218 68.9724
R929 B.n512 B.n214 68.9724
R930 B.n519 B.n214 68.9724
R931 B.n525 B.n210 68.9724
R932 B.n525 B.n4 68.9724
R933 B.n654 B.n4 68.9724
R934 B.n654 B.n653 68.9724
R935 B.n653 B.n652 68.9724
R936 B.n652 B.n8 68.9724
R937 B.n534 B.n8 68.9724
R938 B.n645 B.n644 68.9724
R939 B.n644 B.n643 68.9724
R940 B.n643 B.n15 68.9724
R941 B.n637 B.n15 68.9724
R942 B.n637 B.n636 68.9724
R943 B.n635 B.n22 68.9724
R944 B.n629 B.n22 68.9724
R945 B.n629 B.n628 68.9724
R946 B.n628 B.n627 68.9724
R947 B.n627 B.n29 68.9724
R948 B.n621 B.n620 68.9724
R949 B.n620 B.n619 68.9724
R950 B.n619 B.n36 68.9724
R951 B.n613 B.n36 68.9724
R952 B.n613 B.n612 68.9724
R953 B.n611 B.n43 68.9724
R954 B.n605 B.n43 68.9724
R955 B.n605 B.n604 68.9724
R956 B.n604 B.n603 68.9724
R957 B.n603 B.n50 68.9724
R958 B.n597 B.n50 68.9724
R959 B.n597 B.n596 68.9724
R960 B.n595 B.n57 68.9724
R961 B.n589 B.n57 68.9724
R962 B.n589 B.n588 68.9724
R963 B.n588 B.n587 68.9724
R964 B.n587 B.n64 68.9724
R965 B.n581 B.n64 68.9724
R966 B.t6 B.n262 67.9581
R967 B.n596 B.t10 67.9581
R968 B.t1 B.n210 65.9295
R969 B.n534 B.t2 65.9295
R970 B.n464 B.t4 63.9009
R971 B.t3 B.n611 63.9009
R972 B.n146 B.n101 59.5399
R973 B.n99 B.n98 59.5399
R974 B.n371 B.n370 59.5399
R975 B.n352 B.n297 59.5399
R976 B.t20 B.n222 45.6437
R977 B.n636 B.t21 45.6437
R978 B.n482 B.t19 43.6151
R979 B.n621 B.t0 43.6151
R980 B.n101 B.n100 37.6247
R981 B.n98 B.n97 37.6247
R982 B.n370 B.n369 37.6247
R983 B.n297 B.n296 37.6247
R984 B.n424 B.n276 33.8737
R985 B.n420 B.n419 33.8737
R986 B.n578 B.n577 33.8737
R987 B.n583 B.n66 33.8737
R988 B.t19 B.n234 25.3578
R989 B.t0 B.n29 25.3578
R990 B.n500 B.t20 23.3292
R991 B.t21 B.n635 23.3292
R992 B B.n657 18.0485
R993 B.n425 B.n424 10.6151
R994 B.n426 B.n425 10.6151
R995 B.n426 B.n268 10.6151
R996 B.n436 B.n268 10.6151
R997 B.n437 B.n436 10.6151
R998 B.n438 B.n437 10.6151
R999 B.n438 B.n260 10.6151
R1000 B.n448 B.n260 10.6151
R1001 B.n449 B.n448 10.6151
R1002 B.n450 B.n449 10.6151
R1003 B.n450 B.n252 10.6151
R1004 B.n460 B.n252 10.6151
R1005 B.n461 B.n460 10.6151
R1006 B.n462 B.n461 10.6151
R1007 B.n462 B.n244 10.6151
R1008 B.n472 B.n244 10.6151
R1009 B.n473 B.n472 10.6151
R1010 B.n474 B.n473 10.6151
R1011 B.n474 B.n236 10.6151
R1012 B.n484 B.n236 10.6151
R1013 B.n485 B.n484 10.6151
R1014 B.n486 B.n485 10.6151
R1015 B.n486 B.n228 10.6151
R1016 B.n496 B.n228 10.6151
R1017 B.n497 B.n496 10.6151
R1018 B.n498 B.n497 10.6151
R1019 B.n498 B.n220 10.6151
R1020 B.n508 B.n220 10.6151
R1021 B.n509 B.n508 10.6151
R1022 B.n510 B.n509 10.6151
R1023 B.n510 B.n212 10.6151
R1024 B.n521 B.n212 10.6151
R1025 B.n522 B.n521 10.6151
R1026 B.n523 B.n522 10.6151
R1027 B.n523 B.n0 10.6151
R1028 B.n310 B.n276 10.6151
R1029 B.n311 B.n310 10.6151
R1030 B.n312 B.n311 10.6151
R1031 B.n312 B.n306 10.6151
R1032 B.n318 B.n306 10.6151
R1033 B.n319 B.n318 10.6151
R1034 B.n320 B.n319 10.6151
R1035 B.n320 B.n304 10.6151
R1036 B.n326 B.n304 10.6151
R1037 B.n327 B.n326 10.6151
R1038 B.n328 B.n327 10.6151
R1039 B.n328 B.n302 10.6151
R1040 B.n334 B.n302 10.6151
R1041 B.n335 B.n334 10.6151
R1042 B.n336 B.n335 10.6151
R1043 B.n336 B.n300 10.6151
R1044 B.n342 B.n300 10.6151
R1045 B.n343 B.n342 10.6151
R1046 B.n344 B.n343 10.6151
R1047 B.n344 B.n298 10.6151
R1048 B.n350 B.n298 10.6151
R1049 B.n351 B.n350 10.6151
R1050 B.n353 B.n294 10.6151
R1051 B.n359 B.n294 10.6151
R1052 B.n360 B.n359 10.6151
R1053 B.n361 B.n360 10.6151
R1054 B.n361 B.n292 10.6151
R1055 B.n367 B.n292 10.6151
R1056 B.n368 B.n367 10.6151
R1057 B.n372 B.n368 10.6151
R1058 B.n378 B.n290 10.6151
R1059 B.n379 B.n378 10.6151
R1060 B.n380 B.n379 10.6151
R1061 B.n380 B.n288 10.6151
R1062 B.n386 B.n288 10.6151
R1063 B.n387 B.n386 10.6151
R1064 B.n388 B.n387 10.6151
R1065 B.n388 B.n286 10.6151
R1066 B.n394 B.n286 10.6151
R1067 B.n395 B.n394 10.6151
R1068 B.n396 B.n395 10.6151
R1069 B.n396 B.n284 10.6151
R1070 B.n402 B.n284 10.6151
R1071 B.n403 B.n402 10.6151
R1072 B.n404 B.n403 10.6151
R1073 B.n404 B.n282 10.6151
R1074 B.n410 B.n282 10.6151
R1075 B.n411 B.n410 10.6151
R1076 B.n412 B.n411 10.6151
R1077 B.n412 B.n280 10.6151
R1078 B.n418 B.n280 10.6151
R1079 B.n419 B.n418 10.6151
R1080 B.n420 B.n272 10.6151
R1081 B.n430 B.n272 10.6151
R1082 B.n431 B.n430 10.6151
R1083 B.n432 B.n431 10.6151
R1084 B.n432 B.n264 10.6151
R1085 B.n442 B.n264 10.6151
R1086 B.n443 B.n442 10.6151
R1087 B.n444 B.n443 10.6151
R1088 B.n444 B.n256 10.6151
R1089 B.n454 B.n256 10.6151
R1090 B.n455 B.n454 10.6151
R1091 B.n456 B.n455 10.6151
R1092 B.n456 B.n248 10.6151
R1093 B.n466 B.n248 10.6151
R1094 B.n467 B.n466 10.6151
R1095 B.n468 B.n467 10.6151
R1096 B.n468 B.n240 10.6151
R1097 B.n478 B.n240 10.6151
R1098 B.n479 B.n478 10.6151
R1099 B.n480 B.n479 10.6151
R1100 B.n480 B.n232 10.6151
R1101 B.n490 B.n232 10.6151
R1102 B.n491 B.n490 10.6151
R1103 B.n492 B.n491 10.6151
R1104 B.n492 B.n224 10.6151
R1105 B.n502 B.n224 10.6151
R1106 B.n503 B.n502 10.6151
R1107 B.n504 B.n503 10.6151
R1108 B.n504 B.n216 10.6151
R1109 B.n514 B.n216 10.6151
R1110 B.n515 B.n514 10.6151
R1111 B.n517 B.n515 10.6151
R1112 B.n517 B.n516 10.6151
R1113 B.n516 B.n208 10.6151
R1114 B.n528 B.n208 10.6151
R1115 B.n529 B.n528 10.6151
R1116 B.n530 B.n529 10.6151
R1117 B.n531 B.n530 10.6151
R1118 B.n532 B.n531 10.6151
R1119 B.n536 B.n532 10.6151
R1120 B.n537 B.n536 10.6151
R1121 B.n538 B.n537 10.6151
R1122 B.n539 B.n538 10.6151
R1123 B.n541 B.n539 10.6151
R1124 B.n542 B.n541 10.6151
R1125 B.n543 B.n542 10.6151
R1126 B.n544 B.n543 10.6151
R1127 B.n546 B.n544 10.6151
R1128 B.n547 B.n546 10.6151
R1129 B.n548 B.n547 10.6151
R1130 B.n549 B.n548 10.6151
R1131 B.n551 B.n549 10.6151
R1132 B.n552 B.n551 10.6151
R1133 B.n553 B.n552 10.6151
R1134 B.n554 B.n553 10.6151
R1135 B.n556 B.n554 10.6151
R1136 B.n557 B.n556 10.6151
R1137 B.n558 B.n557 10.6151
R1138 B.n559 B.n558 10.6151
R1139 B.n561 B.n559 10.6151
R1140 B.n562 B.n561 10.6151
R1141 B.n563 B.n562 10.6151
R1142 B.n564 B.n563 10.6151
R1143 B.n566 B.n564 10.6151
R1144 B.n567 B.n566 10.6151
R1145 B.n568 B.n567 10.6151
R1146 B.n569 B.n568 10.6151
R1147 B.n571 B.n569 10.6151
R1148 B.n572 B.n571 10.6151
R1149 B.n573 B.n572 10.6151
R1150 B.n574 B.n573 10.6151
R1151 B.n576 B.n574 10.6151
R1152 B.n577 B.n576 10.6151
R1153 B.n649 B.n1 10.6151
R1154 B.n649 B.n648 10.6151
R1155 B.n648 B.n647 10.6151
R1156 B.n647 B.n10 10.6151
R1157 B.n641 B.n10 10.6151
R1158 B.n641 B.n640 10.6151
R1159 B.n640 B.n639 10.6151
R1160 B.n639 B.n17 10.6151
R1161 B.n633 B.n17 10.6151
R1162 B.n633 B.n632 10.6151
R1163 B.n632 B.n631 10.6151
R1164 B.n631 B.n24 10.6151
R1165 B.n625 B.n24 10.6151
R1166 B.n625 B.n624 10.6151
R1167 B.n624 B.n623 10.6151
R1168 B.n623 B.n31 10.6151
R1169 B.n617 B.n31 10.6151
R1170 B.n617 B.n616 10.6151
R1171 B.n616 B.n615 10.6151
R1172 B.n615 B.n38 10.6151
R1173 B.n609 B.n38 10.6151
R1174 B.n609 B.n608 10.6151
R1175 B.n608 B.n607 10.6151
R1176 B.n607 B.n45 10.6151
R1177 B.n601 B.n45 10.6151
R1178 B.n601 B.n600 10.6151
R1179 B.n600 B.n599 10.6151
R1180 B.n599 B.n52 10.6151
R1181 B.n593 B.n52 10.6151
R1182 B.n593 B.n592 10.6151
R1183 B.n592 B.n591 10.6151
R1184 B.n591 B.n59 10.6151
R1185 B.n585 B.n59 10.6151
R1186 B.n585 B.n584 10.6151
R1187 B.n584 B.n583 10.6151
R1188 B.n102 B.n66 10.6151
R1189 B.n105 B.n102 10.6151
R1190 B.n106 B.n105 10.6151
R1191 B.n109 B.n106 10.6151
R1192 B.n110 B.n109 10.6151
R1193 B.n113 B.n110 10.6151
R1194 B.n114 B.n113 10.6151
R1195 B.n117 B.n114 10.6151
R1196 B.n118 B.n117 10.6151
R1197 B.n121 B.n118 10.6151
R1198 B.n122 B.n121 10.6151
R1199 B.n125 B.n122 10.6151
R1200 B.n126 B.n125 10.6151
R1201 B.n129 B.n126 10.6151
R1202 B.n130 B.n129 10.6151
R1203 B.n133 B.n130 10.6151
R1204 B.n134 B.n133 10.6151
R1205 B.n137 B.n134 10.6151
R1206 B.n138 B.n137 10.6151
R1207 B.n141 B.n138 10.6151
R1208 B.n142 B.n141 10.6151
R1209 B.n145 B.n142 10.6151
R1210 B.n150 B.n147 10.6151
R1211 B.n151 B.n150 10.6151
R1212 B.n154 B.n151 10.6151
R1213 B.n155 B.n154 10.6151
R1214 B.n158 B.n155 10.6151
R1215 B.n159 B.n158 10.6151
R1216 B.n162 B.n159 10.6151
R1217 B.n163 B.n162 10.6151
R1218 B.n167 B.n166 10.6151
R1219 B.n170 B.n167 10.6151
R1220 B.n171 B.n170 10.6151
R1221 B.n174 B.n171 10.6151
R1222 B.n175 B.n174 10.6151
R1223 B.n178 B.n175 10.6151
R1224 B.n179 B.n178 10.6151
R1225 B.n182 B.n179 10.6151
R1226 B.n183 B.n182 10.6151
R1227 B.n186 B.n183 10.6151
R1228 B.n187 B.n186 10.6151
R1229 B.n190 B.n187 10.6151
R1230 B.n191 B.n190 10.6151
R1231 B.n194 B.n191 10.6151
R1232 B.n195 B.n194 10.6151
R1233 B.n198 B.n195 10.6151
R1234 B.n199 B.n198 10.6151
R1235 B.n202 B.n199 10.6151
R1236 B.n203 B.n202 10.6151
R1237 B.n206 B.n203 10.6151
R1238 B.n207 B.n206 10.6151
R1239 B.n578 B.n207 10.6151
R1240 B.n657 B.n0 8.11757
R1241 B.n657 B.n1 8.11757
R1242 B.n353 B.n352 6.5566
R1243 B.n372 B.n371 6.5566
R1244 B.n147 B.n146 6.5566
R1245 B.n163 B.n99 6.5566
R1246 B.t4 B.n246 5.07196
R1247 B.n612 B.t3 5.07196
R1248 B.n352 B.n351 4.05904
R1249 B.n371 B.n290 4.05904
R1250 B.n146 B.n145 4.05904
R1251 B.n166 B.n99 4.05904
R1252 B.n519 B.t1 3.04338
R1253 B.n645 B.t2 3.04338
R1254 B.n440 B.t6 1.01479
R1255 B.t10 B.n595 1.01479
R1256 VP.n28 VP.n27 177.939
R1257 VP.n50 VP.n49 177.939
R1258 VP.n26 VP.n25 177.939
R1259 VP.n13 VP.n12 161.3
R1260 VP.n14 VP.n9 161.3
R1261 VP.n16 VP.n15 161.3
R1262 VP.n17 VP.n8 161.3
R1263 VP.n20 VP.n19 161.3
R1264 VP.n21 VP.n7 161.3
R1265 VP.n23 VP.n22 161.3
R1266 VP.n24 VP.n6 161.3
R1267 VP.n48 VP.n0 161.3
R1268 VP.n47 VP.n46 161.3
R1269 VP.n45 VP.n1 161.3
R1270 VP.n44 VP.n43 161.3
R1271 VP.n41 VP.n2 161.3
R1272 VP.n40 VP.n39 161.3
R1273 VP.n38 VP.n3 161.3
R1274 VP.n37 VP.n36 161.3
R1275 VP.n34 VP.n4 161.3
R1276 VP.n33 VP.n32 161.3
R1277 VP.n31 VP.n5 161.3
R1278 VP.n30 VP.n29 161.3
R1279 VP.n10 VP.t4 115.96
R1280 VP.n28 VP.t3 83.3775
R1281 VP.n35 VP.t0 83.3775
R1282 VP.n42 VP.t2 83.3775
R1283 VP.n49 VP.t7 83.3775
R1284 VP.n25 VP.t5 83.3775
R1285 VP.n18 VP.t6 83.3775
R1286 VP.n11 VP.t1 83.3775
R1287 VP.n33 VP.n5 56.5193
R1288 VP.n40 VP.n3 56.5193
R1289 VP.n47 VP.n1 56.5193
R1290 VP.n23 VP.n7 56.5193
R1291 VP.n16 VP.n9 56.5193
R1292 VP.n11 VP.n10 55.3922
R1293 VP.n27 VP.n26 41.3111
R1294 VP.n29 VP.n5 24.4675
R1295 VP.n34 VP.n33 24.4675
R1296 VP.n36 VP.n3 24.4675
R1297 VP.n41 VP.n40 24.4675
R1298 VP.n43 VP.n1 24.4675
R1299 VP.n48 VP.n47 24.4675
R1300 VP.n24 VP.n23 24.4675
R1301 VP.n17 VP.n16 24.4675
R1302 VP.n19 VP.n7 24.4675
R1303 VP.n12 VP.n9 24.4675
R1304 VP.n13 VP.n10 17.9991
R1305 VP.n35 VP.n34 13.702
R1306 VP.n43 VP.n42 13.702
R1307 VP.n19 VP.n18 13.702
R1308 VP.n36 VP.n35 10.766
R1309 VP.n42 VP.n41 10.766
R1310 VP.n18 VP.n17 10.766
R1311 VP.n12 VP.n11 10.766
R1312 VP.n29 VP.n28 7.82994
R1313 VP.n49 VP.n48 7.82994
R1314 VP.n25 VP.n24 7.82994
R1315 VP.n14 VP.n13 0.189894
R1316 VP.n15 VP.n14 0.189894
R1317 VP.n15 VP.n8 0.189894
R1318 VP.n20 VP.n8 0.189894
R1319 VP.n21 VP.n20 0.189894
R1320 VP.n22 VP.n21 0.189894
R1321 VP.n22 VP.n6 0.189894
R1322 VP.n26 VP.n6 0.189894
R1323 VP.n30 VP.n27 0.189894
R1324 VP.n31 VP.n30 0.189894
R1325 VP.n32 VP.n31 0.189894
R1326 VP.n32 VP.n4 0.189894
R1327 VP.n37 VP.n4 0.189894
R1328 VP.n38 VP.n37 0.189894
R1329 VP.n39 VP.n38 0.189894
R1330 VP.n39 VP.n2 0.189894
R1331 VP.n44 VP.n2 0.189894
R1332 VP.n45 VP.n44 0.189894
R1333 VP.n46 VP.n45 0.189894
R1334 VP.n46 VP.n0 0.189894
R1335 VP.n50 VP.n0 0.189894
R1336 VP VP.n50 0.0516364
R1337 VDD1 VDD1.n0 67.4068
R1338 VDD1.n3 VDD1.n2 67.2931
R1339 VDD1.n3 VDD1.n1 67.2931
R1340 VDD1.n5 VDD1.n4 66.5123
R1341 VDD1.n5 VDD1.n3 36.6259
R1342 VDD1.n4 VDD1.t1 3.55526
R1343 VDD1.n4 VDD1.t2 3.55526
R1344 VDD1.n0 VDD1.t3 3.55526
R1345 VDD1.n0 VDD1.t6 3.55526
R1346 VDD1.n2 VDD1.t5 3.55526
R1347 VDD1.n2 VDD1.t0 3.55526
R1348 VDD1.n1 VDD1.t4 3.55526
R1349 VDD1.n1 VDD1.t7 3.55526
R1350 VDD1 VDD1.n5 0.778517
C0 VN VDD2 3.81181f
C1 VP VTAIL 4.28478f
C2 VDD1 VDD2 1.26555f
C3 VN VDD1 0.150011f
C4 VP VDD2 0.414397f
C5 VP VN 5.26052f
C6 VDD2 VTAIL 5.54571f
C7 VN VTAIL 4.27067f
C8 VP VDD1 4.0753f
C9 VDD1 VTAIL 5.497931f
C10 VDD2 B 3.887634f
C11 VDD1 B 4.226163f
C12 VTAIL B 5.718674f
C13 VN B 11.07413f
C14 VP B 9.62326f
C15 VDD1.t3 B 0.110426f
C16 VDD1.t6 B 0.110426f
C17 VDD1.n0 B 0.917607f
C18 VDD1.t4 B 0.110426f
C19 VDD1.t7 B 0.110426f
C20 VDD1.n1 B 0.916806f
C21 VDD1.t5 B 0.110426f
C22 VDD1.t0 B 0.110426f
C23 VDD1.n2 B 0.916806f
C24 VDD1.n3 B 2.36641f
C25 VDD1.t1 B 0.110426f
C26 VDD1.t2 B 0.110426f
C27 VDD1.n4 B 0.912028f
C28 VDD1.n5 B 2.13719f
C29 VP.n0 B 0.033073f
C30 VP.t7 B 0.78143f
C31 VP.n1 B 0.04275f
C32 VP.n2 B 0.033073f
C33 VP.t2 B 0.78143f
C34 VP.n3 B 0.04828f
C35 VP.n4 B 0.033073f
C36 VP.t0 B 0.78143f
C37 VP.n5 B 0.05381f
C38 VP.n6 B 0.033073f
C39 VP.t5 B 0.78143f
C40 VP.n7 B 0.04275f
C41 VP.n8 B 0.033073f
C42 VP.t6 B 0.78143f
C43 VP.n9 B 0.04828f
C44 VP.t4 B 0.905882f
C45 VP.n10 B 0.380183f
C46 VP.t1 B 0.78143f
C47 VP.n11 B 0.370433f
C48 VP.n12 B 0.044597f
C49 VP.n13 B 0.210939f
C50 VP.n14 B 0.033073f
C51 VP.n15 B 0.033073f
C52 VP.n16 B 0.04828f
C53 VP.n17 B 0.044597f
C54 VP.n18 B 0.307489f
C55 VP.n19 B 0.048249f
C56 VP.n20 B 0.033073f
C57 VP.n21 B 0.033073f
C58 VP.n22 B 0.033073f
C59 VP.n23 B 0.05381f
C60 VP.n24 B 0.040946f
C61 VP.n25 B 0.378261f
C62 VP.n26 B 1.33512f
C63 VP.n27 B 1.36389f
C64 VP.t3 B 0.78143f
C65 VP.n28 B 0.378261f
C66 VP.n29 B 0.040946f
C67 VP.n30 B 0.033073f
C68 VP.n31 B 0.033073f
C69 VP.n32 B 0.033073f
C70 VP.n33 B 0.04275f
C71 VP.n34 B 0.048249f
C72 VP.n35 B 0.307489f
C73 VP.n36 B 0.044597f
C74 VP.n37 B 0.033073f
C75 VP.n38 B 0.033073f
C76 VP.n39 B 0.033073f
C77 VP.n40 B 0.04828f
C78 VP.n41 B 0.044597f
C79 VP.n42 B 0.307489f
C80 VP.n43 B 0.048249f
C81 VP.n44 B 0.033073f
C82 VP.n45 B 0.033073f
C83 VP.n46 B 0.033073f
C84 VP.n47 B 0.05381f
C85 VP.n48 B 0.040946f
C86 VP.n49 B 0.378261f
C87 VP.n50 B 0.03293f
C88 VTAIL.t11 B 0.098246f
C89 VTAIL.t14 B 0.098246f
C90 VTAIL.n0 B 0.752551f
C91 VTAIL.n1 B 0.333204f
C92 VTAIL.t7 B 0.959089f
C93 VTAIL.n2 B 0.424216f
C94 VTAIL.t1 B 0.959089f
C95 VTAIL.n3 B 0.424216f
C96 VTAIL.t5 B 0.098246f
C97 VTAIL.t6 B 0.098246f
C98 VTAIL.n4 B 0.752551f
C99 VTAIL.n5 B 0.449302f
C100 VTAIL.t4 B 0.959089f
C101 VTAIL.n6 B 1.15926f
C102 VTAIL.t8 B 0.959093f
C103 VTAIL.n7 B 1.15926f
C104 VTAIL.t13 B 0.098246f
C105 VTAIL.t12 B 0.098246f
C106 VTAIL.n8 B 0.752555f
C107 VTAIL.n9 B 0.449298f
C108 VTAIL.t9 B 0.959093f
C109 VTAIL.n10 B 0.424212f
C110 VTAIL.t2 B 0.959093f
C111 VTAIL.n11 B 0.424212f
C112 VTAIL.t15 B 0.098246f
C113 VTAIL.t0 B 0.098246f
C114 VTAIL.n12 B 0.752555f
C115 VTAIL.n13 B 0.449298f
C116 VTAIL.t3 B 0.959089f
C117 VTAIL.n14 B 1.15926f
C118 VTAIL.t10 B 0.959089f
C119 VTAIL.n15 B 1.15507f
C120 VDD2.t3 B 0.108018f
C121 VDD2.t2 B 0.108018f
C122 VDD2.n0 B 0.896812f
C123 VDD2.t4 B 0.108018f
C124 VDD2.t5 B 0.108018f
C125 VDD2.n1 B 0.896812f
C126 VDD2.n2 B 2.26288f
C127 VDD2.t7 B 0.108018f
C128 VDD2.t0 B 0.108018f
C129 VDD2.n3 B 0.892142f
C130 VDD2.n4 B 2.06107f
C131 VDD2.t6 B 0.108018f
C132 VDD2.t1 B 0.108018f
C133 VDD2.n5 B 0.896783f
C134 VN.n0 B 0.032239f
C135 VN.t4 B 0.761734f
C136 VN.n1 B 0.041673f
C137 VN.n2 B 0.032239f
C138 VN.t0 B 0.761734f
C139 VN.n3 B 0.047063f
C140 VN.t7 B 0.883049f
C141 VN.n4 B 0.3706f
C142 VN.t3 B 0.761734f
C143 VN.n5 B 0.361096f
C144 VN.n6 B 0.043473f
C145 VN.n7 B 0.205622f
C146 VN.n8 B 0.032239f
C147 VN.n9 B 0.032239f
C148 VN.n10 B 0.047063f
C149 VN.n11 B 0.043473f
C150 VN.n12 B 0.299738f
C151 VN.n13 B 0.047033f
C152 VN.n14 B 0.032239f
C153 VN.n15 B 0.032239f
C154 VN.n16 B 0.032239f
C155 VN.n17 B 0.052453f
C156 VN.n18 B 0.039914f
C157 VN.n19 B 0.368726f
C158 VN.n20 B 0.0321f
C159 VN.n21 B 0.032239f
C160 VN.t6 B 0.761734f
C161 VN.n22 B 0.041673f
C162 VN.n23 B 0.032239f
C163 VN.t1 B 0.761734f
C164 VN.n24 B 0.047063f
C165 VN.t5 B 0.883049f
C166 VN.n25 B 0.3706f
C167 VN.t2 B 0.761734f
C168 VN.n26 B 0.361096f
C169 VN.n27 B 0.043473f
C170 VN.n28 B 0.205622f
C171 VN.n29 B 0.032239f
C172 VN.n30 B 0.032239f
C173 VN.n31 B 0.047063f
C174 VN.n32 B 0.043473f
C175 VN.n33 B 0.299738f
C176 VN.n34 B 0.047033f
C177 VN.n35 B 0.032239f
C178 VN.n36 B 0.032239f
C179 VN.n37 B 0.032239f
C180 VN.n38 B 0.052453f
C181 VN.n39 B 0.039914f
C182 VN.n40 B 0.368726f
C183 VN.n41 B 1.32265f
.ends

