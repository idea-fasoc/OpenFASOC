* NGSPICE file created from diff_pair_sample_0911.ext - technology: sky130A

.subckt diff_pair_sample_0911 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t12 VP.t0 VDD1.t3 w_n3540_n1870# sky130_fd_pr__pfet_01v8 ad=0.74415 pd=4.84 as=0.74415 ps=4.84 w=4.51 l=2.24
X1 B.t11 B.t9 B.t10 w_n3540_n1870# sky130_fd_pr__pfet_01v8 ad=1.7589 pd=9.8 as=0 ps=0 w=4.51 l=2.24
X2 VDD1.t0 VP.t1 VTAIL.t11 w_n3540_n1870# sky130_fd_pr__pfet_01v8 ad=0.74415 pd=4.84 as=1.7589 ps=9.8 w=4.51 l=2.24
X3 VTAIL.t15 VN.t0 VDD2.t7 w_n3540_n1870# sky130_fd_pr__pfet_01v8 ad=1.7589 pd=9.8 as=0.74415 ps=4.84 w=4.51 l=2.24
X4 VTAIL.t13 VN.t1 VDD2.t6 w_n3540_n1870# sky130_fd_pr__pfet_01v8 ad=0.74415 pd=4.84 as=0.74415 ps=4.84 w=4.51 l=2.24
X5 VDD2.t5 VN.t2 VTAIL.t3 w_n3540_n1870# sky130_fd_pr__pfet_01v8 ad=0.74415 pd=4.84 as=0.74415 ps=4.84 w=4.51 l=2.24
X6 VDD2.t4 VN.t3 VTAIL.t1 w_n3540_n1870# sky130_fd_pr__pfet_01v8 ad=0.74415 pd=4.84 as=1.7589 ps=9.8 w=4.51 l=2.24
X7 VTAIL.t0 VN.t4 VDD2.t3 w_n3540_n1870# sky130_fd_pr__pfet_01v8 ad=1.7589 pd=9.8 as=0.74415 ps=4.84 w=4.51 l=2.24
X8 VTAIL.t10 VP.t2 VDD1.t7 w_n3540_n1870# sky130_fd_pr__pfet_01v8 ad=1.7589 pd=9.8 as=0.74415 ps=4.84 w=4.51 l=2.24
X9 VDD2.t2 VN.t5 VTAIL.t2 w_n3540_n1870# sky130_fd_pr__pfet_01v8 ad=0.74415 pd=4.84 as=1.7589 ps=9.8 w=4.51 l=2.24
X10 B.t8 B.t6 B.t7 w_n3540_n1870# sky130_fd_pr__pfet_01v8 ad=1.7589 pd=9.8 as=0 ps=0 w=4.51 l=2.24
X11 VTAIL.t9 VP.t3 VDD1.t5 w_n3540_n1870# sky130_fd_pr__pfet_01v8 ad=0.74415 pd=4.84 as=0.74415 ps=4.84 w=4.51 l=2.24
X12 VDD1.t1 VP.t4 VTAIL.t8 w_n3540_n1870# sky130_fd_pr__pfet_01v8 ad=0.74415 pd=4.84 as=0.74415 ps=4.84 w=4.51 l=2.24
X13 VDD2.t1 VN.t6 VTAIL.t14 w_n3540_n1870# sky130_fd_pr__pfet_01v8 ad=0.74415 pd=4.84 as=0.74415 ps=4.84 w=4.51 l=2.24
X14 VDD1.t2 VP.t5 VTAIL.t7 w_n3540_n1870# sky130_fd_pr__pfet_01v8 ad=0.74415 pd=4.84 as=0.74415 ps=4.84 w=4.51 l=2.24
X15 B.t5 B.t3 B.t4 w_n3540_n1870# sky130_fd_pr__pfet_01v8 ad=1.7589 pd=9.8 as=0 ps=0 w=4.51 l=2.24
X16 VTAIL.t4 VN.t7 VDD2.t0 w_n3540_n1870# sky130_fd_pr__pfet_01v8 ad=0.74415 pd=4.84 as=0.74415 ps=4.84 w=4.51 l=2.24
X17 VTAIL.t6 VP.t6 VDD1.t6 w_n3540_n1870# sky130_fd_pr__pfet_01v8 ad=1.7589 pd=9.8 as=0.74415 ps=4.84 w=4.51 l=2.24
X18 B.t2 B.t0 B.t1 w_n3540_n1870# sky130_fd_pr__pfet_01v8 ad=1.7589 pd=9.8 as=0 ps=0 w=4.51 l=2.24
X19 VDD1.t4 VP.t7 VTAIL.t5 w_n3540_n1870# sky130_fd_pr__pfet_01v8 ad=0.74415 pd=4.84 as=1.7589 ps=9.8 w=4.51 l=2.24
R0 VP.n16 VP.n15 161.3
R1 VP.n17 VP.n12 161.3
R2 VP.n19 VP.n18 161.3
R3 VP.n20 VP.n11 161.3
R4 VP.n22 VP.n21 161.3
R5 VP.n24 VP.n10 161.3
R6 VP.n26 VP.n25 161.3
R7 VP.n27 VP.n9 161.3
R8 VP.n29 VP.n28 161.3
R9 VP.n30 VP.n8 161.3
R10 VP.n58 VP.n0 161.3
R11 VP.n57 VP.n56 161.3
R12 VP.n55 VP.n1 161.3
R13 VP.n54 VP.n53 161.3
R14 VP.n52 VP.n2 161.3
R15 VP.n50 VP.n49 161.3
R16 VP.n48 VP.n3 161.3
R17 VP.n47 VP.n46 161.3
R18 VP.n45 VP.n4 161.3
R19 VP.n44 VP.n43 161.3
R20 VP.n42 VP.n41 161.3
R21 VP.n40 VP.n6 161.3
R22 VP.n39 VP.n38 161.3
R23 VP.n37 VP.n7 161.3
R24 VP.n36 VP.n35 161.3
R25 VP.n34 VP.n33 93.3849
R26 VP.n60 VP.n59 93.3849
R27 VP.n32 VP.n31 93.3849
R28 VP.n14 VP.t2 81.9516
R29 VP.n14 VP.n13 57.3618
R30 VP.n34 VP.t6 48.5233
R31 VP.n5 VP.t5 48.5233
R32 VP.n51 VP.t0 48.5233
R33 VP.n59 VP.t7 48.5233
R34 VP.n31 VP.t1 48.5233
R35 VP.n23 VP.t3 48.5233
R36 VP.n13 VP.t4 48.5233
R37 VP.n39 VP.n7 47.2923
R38 VP.n57 VP.n1 47.2923
R39 VP.n29 VP.n9 47.2923
R40 VP.n33 VP.n32 43.5829
R41 VP.n46 VP.n45 40.4934
R42 VP.n46 VP.n3 40.4934
R43 VP.n18 VP.n11 40.4934
R44 VP.n18 VP.n17 40.4934
R45 VP.n40 VP.n39 33.6945
R46 VP.n53 VP.n1 33.6945
R47 VP.n25 VP.n9 33.6945
R48 VP.n35 VP.n7 24.4675
R49 VP.n41 VP.n40 24.4675
R50 VP.n45 VP.n44 24.4675
R51 VP.n50 VP.n3 24.4675
R52 VP.n53 VP.n52 24.4675
R53 VP.n58 VP.n57 24.4675
R54 VP.n30 VP.n29 24.4675
R55 VP.n22 VP.n11 24.4675
R56 VP.n25 VP.n24 24.4675
R57 VP.n17 VP.n16 24.4675
R58 VP.n35 VP.n34 17.3721
R59 VP.n59 VP.n58 17.3721
R60 VP.n31 VP.n30 17.3721
R61 VP.n44 VP.n5 13.9467
R62 VP.n51 VP.n50 13.9467
R63 VP.n23 VP.n22 13.9467
R64 VP.n16 VP.n13 13.9467
R65 VP.n41 VP.n5 10.5213
R66 VP.n52 VP.n51 10.5213
R67 VP.n24 VP.n23 10.5213
R68 VP.n15 VP.n14 9.22138
R69 VP.n32 VP.n8 0.278367
R70 VP.n36 VP.n33 0.278367
R71 VP.n60 VP.n0 0.278367
R72 VP.n15 VP.n12 0.189894
R73 VP.n19 VP.n12 0.189894
R74 VP.n20 VP.n19 0.189894
R75 VP.n21 VP.n20 0.189894
R76 VP.n21 VP.n10 0.189894
R77 VP.n26 VP.n10 0.189894
R78 VP.n27 VP.n26 0.189894
R79 VP.n28 VP.n27 0.189894
R80 VP.n28 VP.n8 0.189894
R81 VP.n37 VP.n36 0.189894
R82 VP.n38 VP.n37 0.189894
R83 VP.n38 VP.n6 0.189894
R84 VP.n42 VP.n6 0.189894
R85 VP.n43 VP.n42 0.189894
R86 VP.n43 VP.n4 0.189894
R87 VP.n47 VP.n4 0.189894
R88 VP.n48 VP.n47 0.189894
R89 VP.n49 VP.n48 0.189894
R90 VP.n49 VP.n2 0.189894
R91 VP.n54 VP.n2 0.189894
R92 VP.n55 VP.n54 0.189894
R93 VP.n56 VP.n55 0.189894
R94 VP.n56 VP.n0 0.189894
R95 VP VP.n60 0.153454
R96 VDD1 VDD1.n0 104.276
R97 VDD1.n3 VDD1.n2 104.162
R98 VDD1.n3 VDD1.n1 104.162
R99 VDD1.n5 VDD1.n4 103.109
R100 VDD1.n5 VDD1.n3 38.1561
R101 VDD1.n4 VDD1.t5 7.20782
R102 VDD1.n4 VDD1.t0 7.20782
R103 VDD1.n0 VDD1.t7 7.20782
R104 VDD1.n0 VDD1.t1 7.20782
R105 VDD1.n2 VDD1.t3 7.20782
R106 VDD1.n2 VDD1.t4 7.20782
R107 VDD1.n1 VDD1.t6 7.20782
R108 VDD1.n1 VDD1.t2 7.20782
R109 VDD1 VDD1.n5 1.05007
R110 VTAIL.n194 VTAIL.n176 756.745
R111 VTAIL.n20 VTAIL.n2 756.745
R112 VTAIL.n44 VTAIL.n26 756.745
R113 VTAIL.n70 VTAIL.n52 756.745
R114 VTAIL.n170 VTAIL.n152 756.745
R115 VTAIL.n144 VTAIL.n126 756.745
R116 VTAIL.n120 VTAIL.n102 756.745
R117 VTAIL.n94 VTAIL.n76 756.745
R118 VTAIL.n185 VTAIL.n184 585
R119 VTAIL.n187 VTAIL.n186 585
R120 VTAIL.n180 VTAIL.n179 585
R121 VTAIL.n193 VTAIL.n192 585
R122 VTAIL.n195 VTAIL.n194 585
R123 VTAIL.n11 VTAIL.n10 585
R124 VTAIL.n13 VTAIL.n12 585
R125 VTAIL.n6 VTAIL.n5 585
R126 VTAIL.n19 VTAIL.n18 585
R127 VTAIL.n21 VTAIL.n20 585
R128 VTAIL.n35 VTAIL.n34 585
R129 VTAIL.n37 VTAIL.n36 585
R130 VTAIL.n30 VTAIL.n29 585
R131 VTAIL.n43 VTAIL.n42 585
R132 VTAIL.n45 VTAIL.n44 585
R133 VTAIL.n61 VTAIL.n60 585
R134 VTAIL.n63 VTAIL.n62 585
R135 VTAIL.n56 VTAIL.n55 585
R136 VTAIL.n69 VTAIL.n68 585
R137 VTAIL.n71 VTAIL.n70 585
R138 VTAIL.n171 VTAIL.n170 585
R139 VTAIL.n169 VTAIL.n168 585
R140 VTAIL.n156 VTAIL.n155 585
R141 VTAIL.n163 VTAIL.n162 585
R142 VTAIL.n161 VTAIL.n160 585
R143 VTAIL.n145 VTAIL.n144 585
R144 VTAIL.n143 VTAIL.n142 585
R145 VTAIL.n130 VTAIL.n129 585
R146 VTAIL.n137 VTAIL.n136 585
R147 VTAIL.n135 VTAIL.n134 585
R148 VTAIL.n121 VTAIL.n120 585
R149 VTAIL.n119 VTAIL.n118 585
R150 VTAIL.n106 VTAIL.n105 585
R151 VTAIL.n113 VTAIL.n112 585
R152 VTAIL.n111 VTAIL.n110 585
R153 VTAIL.n95 VTAIL.n94 585
R154 VTAIL.n93 VTAIL.n92 585
R155 VTAIL.n80 VTAIL.n79 585
R156 VTAIL.n87 VTAIL.n86 585
R157 VTAIL.n85 VTAIL.n84 585
R158 VTAIL.n183 VTAIL.t2 328.587
R159 VTAIL.n9 VTAIL.t0 328.587
R160 VTAIL.n33 VTAIL.t5 328.587
R161 VTAIL.n59 VTAIL.t6 328.587
R162 VTAIL.n159 VTAIL.t11 328.587
R163 VTAIL.n133 VTAIL.t10 328.587
R164 VTAIL.n109 VTAIL.t1 328.587
R165 VTAIL.n83 VTAIL.t15 328.587
R166 VTAIL.n186 VTAIL.n185 171.744
R167 VTAIL.n186 VTAIL.n179 171.744
R168 VTAIL.n193 VTAIL.n179 171.744
R169 VTAIL.n194 VTAIL.n193 171.744
R170 VTAIL.n12 VTAIL.n11 171.744
R171 VTAIL.n12 VTAIL.n5 171.744
R172 VTAIL.n19 VTAIL.n5 171.744
R173 VTAIL.n20 VTAIL.n19 171.744
R174 VTAIL.n36 VTAIL.n35 171.744
R175 VTAIL.n36 VTAIL.n29 171.744
R176 VTAIL.n43 VTAIL.n29 171.744
R177 VTAIL.n44 VTAIL.n43 171.744
R178 VTAIL.n62 VTAIL.n61 171.744
R179 VTAIL.n62 VTAIL.n55 171.744
R180 VTAIL.n69 VTAIL.n55 171.744
R181 VTAIL.n70 VTAIL.n69 171.744
R182 VTAIL.n170 VTAIL.n169 171.744
R183 VTAIL.n169 VTAIL.n155 171.744
R184 VTAIL.n162 VTAIL.n155 171.744
R185 VTAIL.n162 VTAIL.n161 171.744
R186 VTAIL.n144 VTAIL.n143 171.744
R187 VTAIL.n143 VTAIL.n129 171.744
R188 VTAIL.n136 VTAIL.n129 171.744
R189 VTAIL.n136 VTAIL.n135 171.744
R190 VTAIL.n120 VTAIL.n119 171.744
R191 VTAIL.n119 VTAIL.n105 171.744
R192 VTAIL.n112 VTAIL.n105 171.744
R193 VTAIL.n112 VTAIL.n111 171.744
R194 VTAIL.n94 VTAIL.n93 171.744
R195 VTAIL.n93 VTAIL.n79 171.744
R196 VTAIL.n86 VTAIL.n79 171.744
R197 VTAIL.n86 VTAIL.n85 171.744
R198 VTAIL.n151 VTAIL.n150 86.4313
R199 VTAIL.n101 VTAIL.n100 86.4313
R200 VTAIL.n1 VTAIL.n0 86.4312
R201 VTAIL.n51 VTAIL.n50 86.4312
R202 VTAIL.n185 VTAIL.t2 85.8723
R203 VTAIL.n11 VTAIL.t0 85.8723
R204 VTAIL.n35 VTAIL.t5 85.8723
R205 VTAIL.n61 VTAIL.t6 85.8723
R206 VTAIL.n161 VTAIL.t11 85.8723
R207 VTAIL.n135 VTAIL.t10 85.8723
R208 VTAIL.n111 VTAIL.t1 85.8723
R209 VTAIL.n85 VTAIL.t15 85.8723
R210 VTAIL.n199 VTAIL.n198 31.2157
R211 VTAIL.n25 VTAIL.n24 31.2157
R212 VTAIL.n49 VTAIL.n48 31.2157
R213 VTAIL.n75 VTAIL.n74 31.2157
R214 VTAIL.n175 VTAIL.n174 31.2157
R215 VTAIL.n149 VTAIL.n148 31.2157
R216 VTAIL.n125 VTAIL.n124 31.2157
R217 VTAIL.n99 VTAIL.n98 31.2157
R218 VTAIL.n199 VTAIL.n175 18.4703
R219 VTAIL.n99 VTAIL.n75 18.4703
R220 VTAIL.n184 VTAIL.n183 16.3651
R221 VTAIL.n10 VTAIL.n9 16.3651
R222 VTAIL.n34 VTAIL.n33 16.3651
R223 VTAIL.n60 VTAIL.n59 16.3651
R224 VTAIL.n160 VTAIL.n159 16.3651
R225 VTAIL.n134 VTAIL.n133 16.3651
R226 VTAIL.n110 VTAIL.n109 16.3651
R227 VTAIL.n84 VTAIL.n83 16.3651
R228 VTAIL.n187 VTAIL.n182 12.8005
R229 VTAIL.n13 VTAIL.n8 12.8005
R230 VTAIL.n37 VTAIL.n32 12.8005
R231 VTAIL.n63 VTAIL.n58 12.8005
R232 VTAIL.n163 VTAIL.n158 12.8005
R233 VTAIL.n137 VTAIL.n132 12.8005
R234 VTAIL.n113 VTAIL.n108 12.8005
R235 VTAIL.n87 VTAIL.n82 12.8005
R236 VTAIL.n188 VTAIL.n180 12.0247
R237 VTAIL.n14 VTAIL.n6 12.0247
R238 VTAIL.n38 VTAIL.n30 12.0247
R239 VTAIL.n64 VTAIL.n56 12.0247
R240 VTAIL.n164 VTAIL.n156 12.0247
R241 VTAIL.n138 VTAIL.n130 12.0247
R242 VTAIL.n114 VTAIL.n106 12.0247
R243 VTAIL.n88 VTAIL.n80 12.0247
R244 VTAIL.n192 VTAIL.n191 11.249
R245 VTAIL.n18 VTAIL.n17 11.249
R246 VTAIL.n42 VTAIL.n41 11.249
R247 VTAIL.n68 VTAIL.n67 11.249
R248 VTAIL.n168 VTAIL.n167 11.249
R249 VTAIL.n142 VTAIL.n141 11.249
R250 VTAIL.n118 VTAIL.n117 11.249
R251 VTAIL.n92 VTAIL.n91 11.249
R252 VTAIL.n195 VTAIL.n178 10.4732
R253 VTAIL.n21 VTAIL.n4 10.4732
R254 VTAIL.n45 VTAIL.n28 10.4732
R255 VTAIL.n71 VTAIL.n54 10.4732
R256 VTAIL.n171 VTAIL.n154 10.4732
R257 VTAIL.n145 VTAIL.n128 10.4732
R258 VTAIL.n121 VTAIL.n104 10.4732
R259 VTAIL.n95 VTAIL.n78 10.4732
R260 VTAIL.n196 VTAIL.n176 9.69747
R261 VTAIL.n22 VTAIL.n2 9.69747
R262 VTAIL.n46 VTAIL.n26 9.69747
R263 VTAIL.n72 VTAIL.n52 9.69747
R264 VTAIL.n172 VTAIL.n152 9.69747
R265 VTAIL.n146 VTAIL.n126 9.69747
R266 VTAIL.n122 VTAIL.n102 9.69747
R267 VTAIL.n96 VTAIL.n76 9.69747
R268 VTAIL.n198 VTAIL.n197 9.45567
R269 VTAIL.n24 VTAIL.n23 9.45567
R270 VTAIL.n48 VTAIL.n47 9.45567
R271 VTAIL.n74 VTAIL.n73 9.45567
R272 VTAIL.n174 VTAIL.n173 9.45567
R273 VTAIL.n148 VTAIL.n147 9.45567
R274 VTAIL.n124 VTAIL.n123 9.45567
R275 VTAIL.n98 VTAIL.n97 9.45567
R276 VTAIL.n197 VTAIL.n196 9.3005
R277 VTAIL.n178 VTAIL.n177 9.3005
R278 VTAIL.n191 VTAIL.n190 9.3005
R279 VTAIL.n189 VTAIL.n188 9.3005
R280 VTAIL.n182 VTAIL.n181 9.3005
R281 VTAIL.n23 VTAIL.n22 9.3005
R282 VTAIL.n4 VTAIL.n3 9.3005
R283 VTAIL.n17 VTAIL.n16 9.3005
R284 VTAIL.n15 VTAIL.n14 9.3005
R285 VTAIL.n8 VTAIL.n7 9.3005
R286 VTAIL.n47 VTAIL.n46 9.3005
R287 VTAIL.n28 VTAIL.n27 9.3005
R288 VTAIL.n41 VTAIL.n40 9.3005
R289 VTAIL.n39 VTAIL.n38 9.3005
R290 VTAIL.n32 VTAIL.n31 9.3005
R291 VTAIL.n73 VTAIL.n72 9.3005
R292 VTAIL.n54 VTAIL.n53 9.3005
R293 VTAIL.n67 VTAIL.n66 9.3005
R294 VTAIL.n65 VTAIL.n64 9.3005
R295 VTAIL.n58 VTAIL.n57 9.3005
R296 VTAIL.n173 VTAIL.n172 9.3005
R297 VTAIL.n154 VTAIL.n153 9.3005
R298 VTAIL.n167 VTAIL.n166 9.3005
R299 VTAIL.n165 VTAIL.n164 9.3005
R300 VTAIL.n158 VTAIL.n157 9.3005
R301 VTAIL.n147 VTAIL.n146 9.3005
R302 VTAIL.n128 VTAIL.n127 9.3005
R303 VTAIL.n141 VTAIL.n140 9.3005
R304 VTAIL.n139 VTAIL.n138 9.3005
R305 VTAIL.n132 VTAIL.n131 9.3005
R306 VTAIL.n123 VTAIL.n122 9.3005
R307 VTAIL.n104 VTAIL.n103 9.3005
R308 VTAIL.n117 VTAIL.n116 9.3005
R309 VTAIL.n115 VTAIL.n114 9.3005
R310 VTAIL.n108 VTAIL.n107 9.3005
R311 VTAIL.n97 VTAIL.n96 9.3005
R312 VTAIL.n78 VTAIL.n77 9.3005
R313 VTAIL.n91 VTAIL.n90 9.3005
R314 VTAIL.n89 VTAIL.n88 9.3005
R315 VTAIL.n82 VTAIL.n81 9.3005
R316 VTAIL.n0 VTAIL.t14 7.20782
R317 VTAIL.n0 VTAIL.t4 7.20782
R318 VTAIL.n50 VTAIL.t7 7.20782
R319 VTAIL.n50 VTAIL.t12 7.20782
R320 VTAIL.n150 VTAIL.t8 7.20782
R321 VTAIL.n150 VTAIL.t9 7.20782
R322 VTAIL.n100 VTAIL.t3 7.20782
R323 VTAIL.n100 VTAIL.t13 7.20782
R324 VTAIL.n198 VTAIL.n176 4.26717
R325 VTAIL.n24 VTAIL.n2 4.26717
R326 VTAIL.n48 VTAIL.n26 4.26717
R327 VTAIL.n74 VTAIL.n52 4.26717
R328 VTAIL.n174 VTAIL.n152 4.26717
R329 VTAIL.n148 VTAIL.n126 4.26717
R330 VTAIL.n124 VTAIL.n102 4.26717
R331 VTAIL.n98 VTAIL.n76 4.26717
R332 VTAIL.n183 VTAIL.n181 3.73474
R333 VTAIL.n9 VTAIL.n7 3.73474
R334 VTAIL.n33 VTAIL.n31 3.73474
R335 VTAIL.n59 VTAIL.n57 3.73474
R336 VTAIL.n159 VTAIL.n157 3.73474
R337 VTAIL.n133 VTAIL.n131 3.73474
R338 VTAIL.n109 VTAIL.n107 3.73474
R339 VTAIL.n83 VTAIL.n81 3.73474
R340 VTAIL.n196 VTAIL.n195 3.49141
R341 VTAIL.n22 VTAIL.n21 3.49141
R342 VTAIL.n46 VTAIL.n45 3.49141
R343 VTAIL.n72 VTAIL.n71 3.49141
R344 VTAIL.n172 VTAIL.n171 3.49141
R345 VTAIL.n146 VTAIL.n145 3.49141
R346 VTAIL.n122 VTAIL.n121 3.49141
R347 VTAIL.n96 VTAIL.n95 3.49141
R348 VTAIL.n192 VTAIL.n178 2.71565
R349 VTAIL.n18 VTAIL.n4 2.71565
R350 VTAIL.n42 VTAIL.n28 2.71565
R351 VTAIL.n68 VTAIL.n54 2.71565
R352 VTAIL.n168 VTAIL.n154 2.71565
R353 VTAIL.n142 VTAIL.n128 2.71565
R354 VTAIL.n118 VTAIL.n104 2.71565
R355 VTAIL.n92 VTAIL.n78 2.71565
R356 VTAIL.n101 VTAIL.n99 2.21602
R357 VTAIL.n125 VTAIL.n101 2.21602
R358 VTAIL.n151 VTAIL.n149 2.21602
R359 VTAIL.n175 VTAIL.n151 2.21602
R360 VTAIL.n75 VTAIL.n51 2.21602
R361 VTAIL.n51 VTAIL.n49 2.21602
R362 VTAIL.n25 VTAIL.n1 2.21602
R363 VTAIL VTAIL.n199 2.15783
R364 VTAIL.n191 VTAIL.n180 1.93989
R365 VTAIL.n17 VTAIL.n6 1.93989
R366 VTAIL.n41 VTAIL.n30 1.93989
R367 VTAIL.n67 VTAIL.n56 1.93989
R368 VTAIL.n167 VTAIL.n156 1.93989
R369 VTAIL.n141 VTAIL.n130 1.93989
R370 VTAIL.n117 VTAIL.n106 1.93989
R371 VTAIL.n91 VTAIL.n80 1.93989
R372 VTAIL.n188 VTAIL.n187 1.16414
R373 VTAIL.n14 VTAIL.n13 1.16414
R374 VTAIL.n38 VTAIL.n37 1.16414
R375 VTAIL.n64 VTAIL.n63 1.16414
R376 VTAIL.n164 VTAIL.n163 1.16414
R377 VTAIL.n138 VTAIL.n137 1.16414
R378 VTAIL.n114 VTAIL.n113 1.16414
R379 VTAIL.n88 VTAIL.n87 1.16414
R380 VTAIL.n149 VTAIL.n125 0.470328
R381 VTAIL.n49 VTAIL.n25 0.470328
R382 VTAIL.n184 VTAIL.n182 0.388379
R383 VTAIL.n10 VTAIL.n8 0.388379
R384 VTAIL.n34 VTAIL.n32 0.388379
R385 VTAIL.n60 VTAIL.n58 0.388379
R386 VTAIL.n160 VTAIL.n158 0.388379
R387 VTAIL.n134 VTAIL.n132 0.388379
R388 VTAIL.n110 VTAIL.n108 0.388379
R389 VTAIL.n84 VTAIL.n82 0.388379
R390 VTAIL.n189 VTAIL.n181 0.155672
R391 VTAIL.n190 VTAIL.n189 0.155672
R392 VTAIL.n190 VTAIL.n177 0.155672
R393 VTAIL.n197 VTAIL.n177 0.155672
R394 VTAIL.n15 VTAIL.n7 0.155672
R395 VTAIL.n16 VTAIL.n15 0.155672
R396 VTAIL.n16 VTAIL.n3 0.155672
R397 VTAIL.n23 VTAIL.n3 0.155672
R398 VTAIL.n39 VTAIL.n31 0.155672
R399 VTAIL.n40 VTAIL.n39 0.155672
R400 VTAIL.n40 VTAIL.n27 0.155672
R401 VTAIL.n47 VTAIL.n27 0.155672
R402 VTAIL.n65 VTAIL.n57 0.155672
R403 VTAIL.n66 VTAIL.n65 0.155672
R404 VTAIL.n66 VTAIL.n53 0.155672
R405 VTAIL.n73 VTAIL.n53 0.155672
R406 VTAIL.n173 VTAIL.n153 0.155672
R407 VTAIL.n166 VTAIL.n153 0.155672
R408 VTAIL.n166 VTAIL.n165 0.155672
R409 VTAIL.n165 VTAIL.n157 0.155672
R410 VTAIL.n147 VTAIL.n127 0.155672
R411 VTAIL.n140 VTAIL.n127 0.155672
R412 VTAIL.n140 VTAIL.n139 0.155672
R413 VTAIL.n139 VTAIL.n131 0.155672
R414 VTAIL.n123 VTAIL.n103 0.155672
R415 VTAIL.n116 VTAIL.n103 0.155672
R416 VTAIL.n116 VTAIL.n115 0.155672
R417 VTAIL.n115 VTAIL.n107 0.155672
R418 VTAIL.n97 VTAIL.n77 0.155672
R419 VTAIL.n90 VTAIL.n77 0.155672
R420 VTAIL.n90 VTAIL.n89 0.155672
R421 VTAIL.n89 VTAIL.n81 0.155672
R422 VTAIL VTAIL.n1 0.0586897
R423 B.n434 B.n53 585
R424 B.n436 B.n435 585
R425 B.n437 B.n52 585
R426 B.n439 B.n438 585
R427 B.n440 B.n51 585
R428 B.n442 B.n441 585
R429 B.n443 B.n50 585
R430 B.n445 B.n444 585
R431 B.n446 B.n49 585
R432 B.n448 B.n447 585
R433 B.n449 B.n48 585
R434 B.n451 B.n450 585
R435 B.n452 B.n47 585
R436 B.n454 B.n453 585
R437 B.n455 B.n46 585
R438 B.n457 B.n456 585
R439 B.n458 B.n45 585
R440 B.n460 B.n459 585
R441 B.n461 B.n44 585
R442 B.n463 B.n462 585
R443 B.n465 B.n41 585
R444 B.n467 B.n466 585
R445 B.n468 B.n40 585
R446 B.n470 B.n469 585
R447 B.n471 B.n39 585
R448 B.n473 B.n472 585
R449 B.n474 B.n38 585
R450 B.n476 B.n475 585
R451 B.n477 B.n35 585
R452 B.n480 B.n479 585
R453 B.n481 B.n34 585
R454 B.n483 B.n482 585
R455 B.n484 B.n33 585
R456 B.n486 B.n485 585
R457 B.n487 B.n32 585
R458 B.n489 B.n488 585
R459 B.n490 B.n31 585
R460 B.n492 B.n491 585
R461 B.n493 B.n30 585
R462 B.n495 B.n494 585
R463 B.n496 B.n29 585
R464 B.n498 B.n497 585
R465 B.n499 B.n28 585
R466 B.n501 B.n500 585
R467 B.n502 B.n27 585
R468 B.n504 B.n503 585
R469 B.n505 B.n26 585
R470 B.n507 B.n506 585
R471 B.n508 B.n25 585
R472 B.n433 B.n432 585
R473 B.n431 B.n54 585
R474 B.n430 B.n429 585
R475 B.n428 B.n55 585
R476 B.n427 B.n426 585
R477 B.n425 B.n56 585
R478 B.n424 B.n423 585
R479 B.n422 B.n57 585
R480 B.n421 B.n420 585
R481 B.n419 B.n58 585
R482 B.n418 B.n417 585
R483 B.n416 B.n59 585
R484 B.n415 B.n414 585
R485 B.n413 B.n60 585
R486 B.n412 B.n411 585
R487 B.n410 B.n61 585
R488 B.n409 B.n408 585
R489 B.n407 B.n62 585
R490 B.n406 B.n405 585
R491 B.n404 B.n63 585
R492 B.n403 B.n402 585
R493 B.n401 B.n64 585
R494 B.n400 B.n399 585
R495 B.n398 B.n65 585
R496 B.n397 B.n396 585
R497 B.n395 B.n66 585
R498 B.n394 B.n393 585
R499 B.n392 B.n67 585
R500 B.n391 B.n390 585
R501 B.n389 B.n68 585
R502 B.n388 B.n387 585
R503 B.n386 B.n69 585
R504 B.n385 B.n384 585
R505 B.n383 B.n70 585
R506 B.n382 B.n381 585
R507 B.n380 B.n71 585
R508 B.n379 B.n378 585
R509 B.n377 B.n72 585
R510 B.n376 B.n375 585
R511 B.n374 B.n73 585
R512 B.n373 B.n372 585
R513 B.n371 B.n74 585
R514 B.n370 B.n369 585
R515 B.n368 B.n75 585
R516 B.n367 B.n366 585
R517 B.n365 B.n76 585
R518 B.n364 B.n363 585
R519 B.n362 B.n77 585
R520 B.n361 B.n360 585
R521 B.n359 B.n78 585
R522 B.n358 B.n357 585
R523 B.n356 B.n79 585
R524 B.n355 B.n354 585
R525 B.n353 B.n80 585
R526 B.n352 B.n351 585
R527 B.n350 B.n81 585
R528 B.n349 B.n348 585
R529 B.n347 B.n82 585
R530 B.n346 B.n345 585
R531 B.n344 B.n83 585
R532 B.n343 B.n342 585
R533 B.n341 B.n84 585
R534 B.n340 B.n339 585
R535 B.n338 B.n85 585
R536 B.n337 B.n336 585
R537 B.n335 B.n86 585
R538 B.n334 B.n333 585
R539 B.n332 B.n87 585
R540 B.n331 B.n330 585
R541 B.n329 B.n88 585
R542 B.n328 B.n327 585
R543 B.n326 B.n89 585
R544 B.n325 B.n324 585
R545 B.n323 B.n90 585
R546 B.n322 B.n321 585
R547 B.n320 B.n91 585
R548 B.n319 B.n318 585
R549 B.n317 B.n92 585
R550 B.n316 B.n315 585
R551 B.n314 B.n93 585
R552 B.n313 B.n312 585
R553 B.n311 B.n94 585
R554 B.n310 B.n309 585
R555 B.n308 B.n95 585
R556 B.n307 B.n306 585
R557 B.n305 B.n96 585
R558 B.n304 B.n303 585
R559 B.n302 B.n97 585
R560 B.n301 B.n300 585
R561 B.n299 B.n98 585
R562 B.n298 B.n297 585
R563 B.n296 B.n99 585
R564 B.n295 B.n294 585
R565 B.n220 B.n219 585
R566 B.n221 B.n128 585
R567 B.n223 B.n222 585
R568 B.n224 B.n127 585
R569 B.n226 B.n225 585
R570 B.n227 B.n126 585
R571 B.n229 B.n228 585
R572 B.n230 B.n125 585
R573 B.n232 B.n231 585
R574 B.n233 B.n124 585
R575 B.n235 B.n234 585
R576 B.n236 B.n123 585
R577 B.n238 B.n237 585
R578 B.n239 B.n122 585
R579 B.n241 B.n240 585
R580 B.n242 B.n121 585
R581 B.n244 B.n243 585
R582 B.n245 B.n120 585
R583 B.n247 B.n246 585
R584 B.n248 B.n117 585
R585 B.n251 B.n250 585
R586 B.n252 B.n116 585
R587 B.n254 B.n253 585
R588 B.n255 B.n115 585
R589 B.n257 B.n256 585
R590 B.n258 B.n114 585
R591 B.n260 B.n259 585
R592 B.n261 B.n113 585
R593 B.n263 B.n262 585
R594 B.n265 B.n264 585
R595 B.n266 B.n109 585
R596 B.n268 B.n267 585
R597 B.n269 B.n108 585
R598 B.n271 B.n270 585
R599 B.n272 B.n107 585
R600 B.n274 B.n273 585
R601 B.n275 B.n106 585
R602 B.n277 B.n276 585
R603 B.n278 B.n105 585
R604 B.n280 B.n279 585
R605 B.n281 B.n104 585
R606 B.n283 B.n282 585
R607 B.n284 B.n103 585
R608 B.n286 B.n285 585
R609 B.n287 B.n102 585
R610 B.n289 B.n288 585
R611 B.n290 B.n101 585
R612 B.n292 B.n291 585
R613 B.n293 B.n100 585
R614 B.n218 B.n129 585
R615 B.n217 B.n216 585
R616 B.n215 B.n130 585
R617 B.n214 B.n213 585
R618 B.n212 B.n131 585
R619 B.n211 B.n210 585
R620 B.n209 B.n132 585
R621 B.n208 B.n207 585
R622 B.n206 B.n133 585
R623 B.n205 B.n204 585
R624 B.n203 B.n134 585
R625 B.n202 B.n201 585
R626 B.n200 B.n135 585
R627 B.n199 B.n198 585
R628 B.n197 B.n136 585
R629 B.n196 B.n195 585
R630 B.n194 B.n137 585
R631 B.n193 B.n192 585
R632 B.n191 B.n138 585
R633 B.n190 B.n189 585
R634 B.n188 B.n139 585
R635 B.n187 B.n186 585
R636 B.n185 B.n140 585
R637 B.n184 B.n183 585
R638 B.n182 B.n141 585
R639 B.n181 B.n180 585
R640 B.n179 B.n142 585
R641 B.n178 B.n177 585
R642 B.n176 B.n143 585
R643 B.n175 B.n174 585
R644 B.n173 B.n144 585
R645 B.n172 B.n171 585
R646 B.n170 B.n145 585
R647 B.n169 B.n168 585
R648 B.n167 B.n146 585
R649 B.n166 B.n165 585
R650 B.n164 B.n147 585
R651 B.n163 B.n162 585
R652 B.n161 B.n148 585
R653 B.n160 B.n159 585
R654 B.n158 B.n149 585
R655 B.n157 B.n156 585
R656 B.n155 B.n150 585
R657 B.n154 B.n153 585
R658 B.n152 B.n151 585
R659 B.n2 B.n0 585
R660 B.n577 B.n1 585
R661 B.n576 B.n575 585
R662 B.n574 B.n3 585
R663 B.n573 B.n572 585
R664 B.n571 B.n4 585
R665 B.n570 B.n569 585
R666 B.n568 B.n5 585
R667 B.n567 B.n566 585
R668 B.n565 B.n6 585
R669 B.n564 B.n563 585
R670 B.n562 B.n7 585
R671 B.n561 B.n560 585
R672 B.n559 B.n8 585
R673 B.n558 B.n557 585
R674 B.n556 B.n9 585
R675 B.n555 B.n554 585
R676 B.n553 B.n10 585
R677 B.n552 B.n551 585
R678 B.n550 B.n11 585
R679 B.n549 B.n548 585
R680 B.n547 B.n12 585
R681 B.n546 B.n545 585
R682 B.n544 B.n13 585
R683 B.n543 B.n542 585
R684 B.n541 B.n14 585
R685 B.n540 B.n539 585
R686 B.n538 B.n15 585
R687 B.n537 B.n536 585
R688 B.n535 B.n16 585
R689 B.n534 B.n533 585
R690 B.n532 B.n17 585
R691 B.n531 B.n530 585
R692 B.n529 B.n18 585
R693 B.n528 B.n527 585
R694 B.n526 B.n19 585
R695 B.n525 B.n524 585
R696 B.n523 B.n20 585
R697 B.n522 B.n521 585
R698 B.n520 B.n21 585
R699 B.n519 B.n518 585
R700 B.n517 B.n22 585
R701 B.n516 B.n515 585
R702 B.n514 B.n23 585
R703 B.n513 B.n512 585
R704 B.n511 B.n24 585
R705 B.n510 B.n509 585
R706 B.n579 B.n578 585
R707 B.n220 B.n129 463.671
R708 B.n510 B.n25 463.671
R709 B.n294 B.n293 463.671
R710 B.n432 B.n53 463.671
R711 B.n110 B.t11 292.442
R712 B.n42 B.t7 292.442
R713 B.n118 B.t2 292.442
R714 B.n36 B.t4 292.442
R715 B.n110 B.t9 255.953
R716 B.n118 B.t0 255.953
R717 B.n36 B.t3 255.953
R718 B.n42 B.t6 255.953
R719 B.n111 B.t10 242.6
R720 B.n43 B.t8 242.6
R721 B.n119 B.t1 242.6
R722 B.n37 B.t5 242.6
R723 B.n216 B.n129 163.367
R724 B.n216 B.n215 163.367
R725 B.n215 B.n214 163.367
R726 B.n214 B.n131 163.367
R727 B.n210 B.n131 163.367
R728 B.n210 B.n209 163.367
R729 B.n209 B.n208 163.367
R730 B.n208 B.n133 163.367
R731 B.n204 B.n133 163.367
R732 B.n204 B.n203 163.367
R733 B.n203 B.n202 163.367
R734 B.n202 B.n135 163.367
R735 B.n198 B.n135 163.367
R736 B.n198 B.n197 163.367
R737 B.n197 B.n196 163.367
R738 B.n196 B.n137 163.367
R739 B.n192 B.n137 163.367
R740 B.n192 B.n191 163.367
R741 B.n191 B.n190 163.367
R742 B.n190 B.n139 163.367
R743 B.n186 B.n139 163.367
R744 B.n186 B.n185 163.367
R745 B.n185 B.n184 163.367
R746 B.n184 B.n141 163.367
R747 B.n180 B.n141 163.367
R748 B.n180 B.n179 163.367
R749 B.n179 B.n178 163.367
R750 B.n178 B.n143 163.367
R751 B.n174 B.n143 163.367
R752 B.n174 B.n173 163.367
R753 B.n173 B.n172 163.367
R754 B.n172 B.n145 163.367
R755 B.n168 B.n145 163.367
R756 B.n168 B.n167 163.367
R757 B.n167 B.n166 163.367
R758 B.n166 B.n147 163.367
R759 B.n162 B.n147 163.367
R760 B.n162 B.n161 163.367
R761 B.n161 B.n160 163.367
R762 B.n160 B.n149 163.367
R763 B.n156 B.n149 163.367
R764 B.n156 B.n155 163.367
R765 B.n155 B.n154 163.367
R766 B.n154 B.n151 163.367
R767 B.n151 B.n2 163.367
R768 B.n578 B.n2 163.367
R769 B.n578 B.n577 163.367
R770 B.n577 B.n576 163.367
R771 B.n576 B.n3 163.367
R772 B.n572 B.n3 163.367
R773 B.n572 B.n571 163.367
R774 B.n571 B.n570 163.367
R775 B.n570 B.n5 163.367
R776 B.n566 B.n5 163.367
R777 B.n566 B.n565 163.367
R778 B.n565 B.n564 163.367
R779 B.n564 B.n7 163.367
R780 B.n560 B.n7 163.367
R781 B.n560 B.n559 163.367
R782 B.n559 B.n558 163.367
R783 B.n558 B.n9 163.367
R784 B.n554 B.n9 163.367
R785 B.n554 B.n553 163.367
R786 B.n553 B.n552 163.367
R787 B.n552 B.n11 163.367
R788 B.n548 B.n11 163.367
R789 B.n548 B.n547 163.367
R790 B.n547 B.n546 163.367
R791 B.n546 B.n13 163.367
R792 B.n542 B.n13 163.367
R793 B.n542 B.n541 163.367
R794 B.n541 B.n540 163.367
R795 B.n540 B.n15 163.367
R796 B.n536 B.n15 163.367
R797 B.n536 B.n535 163.367
R798 B.n535 B.n534 163.367
R799 B.n534 B.n17 163.367
R800 B.n530 B.n17 163.367
R801 B.n530 B.n529 163.367
R802 B.n529 B.n528 163.367
R803 B.n528 B.n19 163.367
R804 B.n524 B.n19 163.367
R805 B.n524 B.n523 163.367
R806 B.n523 B.n522 163.367
R807 B.n522 B.n21 163.367
R808 B.n518 B.n21 163.367
R809 B.n518 B.n517 163.367
R810 B.n517 B.n516 163.367
R811 B.n516 B.n23 163.367
R812 B.n512 B.n23 163.367
R813 B.n512 B.n511 163.367
R814 B.n511 B.n510 163.367
R815 B.n221 B.n220 163.367
R816 B.n222 B.n221 163.367
R817 B.n222 B.n127 163.367
R818 B.n226 B.n127 163.367
R819 B.n227 B.n226 163.367
R820 B.n228 B.n227 163.367
R821 B.n228 B.n125 163.367
R822 B.n232 B.n125 163.367
R823 B.n233 B.n232 163.367
R824 B.n234 B.n233 163.367
R825 B.n234 B.n123 163.367
R826 B.n238 B.n123 163.367
R827 B.n239 B.n238 163.367
R828 B.n240 B.n239 163.367
R829 B.n240 B.n121 163.367
R830 B.n244 B.n121 163.367
R831 B.n245 B.n244 163.367
R832 B.n246 B.n245 163.367
R833 B.n246 B.n117 163.367
R834 B.n251 B.n117 163.367
R835 B.n252 B.n251 163.367
R836 B.n253 B.n252 163.367
R837 B.n253 B.n115 163.367
R838 B.n257 B.n115 163.367
R839 B.n258 B.n257 163.367
R840 B.n259 B.n258 163.367
R841 B.n259 B.n113 163.367
R842 B.n263 B.n113 163.367
R843 B.n264 B.n263 163.367
R844 B.n264 B.n109 163.367
R845 B.n268 B.n109 163.367
R846 B.n269 B.n268 163.367
R847 B.n270 B.n269 163.367
R848 B.n270 B.n107 163.367
R849 B.n274 B.n107 163.367
R850 B.n275 B.n274 163.367
R851 B.n276 B.n275 163.367
R852 B.n276 B.n105 163.367
R853 B.n280 B.n105 163.367
R854 B.n281 B.n280 163.367
R855 B.n282 B.n281 163.367
R856 B.n282 B.n103 163.367
R857 B.n286 B.n103 163.367
R858 B.n287 B.n286 163.367
R859 B.n288 B.n287 163.367
R860 B.n288 B.n101 163.367
R861 B.n292 B.n101 163.367
R862 B.n293 B.n292 163.367
R863 B.n294 B.n99 163.367
R864 B.n298 B.n99 163.367
R865 B.n299 B.n298 163.367
R866 B.n300 B.n299 163.367
R867 B.n300 B.n97 163.367
R868 B.n304 B.n97 163.367
R869 B.n305 B.n304 163.367
R870 B.n306 B.n305 163.367
R871 B.n306 B.n95 163.367
R872 B.n310 B.n95 163.367
R873 B.n311 B.n310 163.367
R874 B.n312 B.n311 163.367
R875 B.n312 B.n93 163.367
R876 B.n316 B.n93 163.367
R877 B.n317 B.n316 163.367
R878 B.n318 B.n317 163.367
R879 B.n318 B.n91 163.367
R880 B.n322 B.n91 163.367
R881 B.n323 B.n322 163.367
R882 B.n324 B.n323 163.367
R883 B.n324 B.n89 163.367
R884 B.n328 B.n89 163.367
R885 B.n329 B.n328 163.367
R886 B.n330 B.n329 163.367
R887 B.n330 B.n87 163.367
R888 B.n334 B.n87 163.367
R889 B.n335 B.n334 163.367
R890 B.n336 B.n335 163.367
R891 B.n336 B.n85 163.367
R892 B.n340 B.n85 163.367
R893 B.n341 B.n340 163.367
R894 B.n342 B.n341 163.367
R895 B.n342 B.n83 163.367
R896 B.n346 B.n83 163.367
R897 B.n347 B.n346 163.367
R898 B.n348 B.n347 163.367
R899 B.n348 B.n81 163.367
R900 B.n352 B.n81 163.367
R901 B.n353 B.n352 163.367
R902 B.n354 B.n353 163.367
R903 B.n354 B.n79 163.367
R904 B.n358 B.n79 163.367
R905 B.n359 B.n358 163.367
R906 B.n360 B.n359 163.367
R907 B.n360 B.n77 163.367
R908 B.n364 B.n77 163.367
R909 B.n365 B.n364 163.367
R910 B.n366 B.n365 163.367
R911 B.n366 B.n75 163.367
R912 B.n370 B.n75 163.367
R913 B.n371 B.n370 163.367
R914 B.n372 B.n371 163.367
R915 B.n372 B.n73 163.367
R916 B.n376 B.n73 163.367
R917 B.n377 B.n376 163.367
R918 B.n378 B.n377 163.367
R919 B.n378 B.n71 163.367
R920 B.n382 B.n71 163.367
R921 B.n383 B.n382 163.367
R922 B.n384 B.n383 163.367
R923 B.n384 B.n69 163.367
R924 B.n388 B.n69 163.367
R925 B.n389 B.n388 163.367
R926 B.n390 B.n389 163.367
R927 B.n390 B.n67 163.367
R928 B.n394 B.n67 163.367
R929 B.n395 B.n394 163.367
R930 B.n396 B.n395 163.367
R931 B.n396 B.n65 163.367
R932 B.n400 B.n65 163.367
R933 B.n401 B.n400 163.367
R934 B.n402 B.n401 163.367
R935 B.n402 B.n63 163.367
R936 B.n406 B.n63 163.367
R937 B.n407 B.n406 163.367
R938 B.n408 B.n407 163.367
R939 B.n408 B.n61 163.367
R940 B.n412 B.n61 163.367
R941 B.n413 B.n412 163.367
R942 B.n414 B.n413 163.367
R943 B.n414 B.n59 163.367
R944 B.n418 B.n59 163.367
R945 B.n419 B.n418 163.367
R946 B.n420 B.n419 163.367
R947 B.n420 B.n57 163.367
R948 B.n424 B.n57 163.367
R949 B.n425 B.n424 163.367
R950 B.n426 B.n425 163.367
R951 B.n426 B.n55 163.367
R952 B.n430 B.n55 163.367
R953 B.n431 B.n430 163.367
R954 B.n432 B.n431 163.367
R955 B.n506 B.n25 163.367
R956 B.n506 B.n505 163.367
R957 B.n505 B.n504 163.367
R958 B.n504 B.n27 163.367
R959 B.n500 B.n27 163.367
R960 B.n500 B.n499 163.367
R961 B.n499 B.n498 163.367
R962 B.n498 B.n29 163.367
R963 B.n494 B.n29 163.367
R964 B.n494 B.n493 163.367
R965 B.n493 B.n492 163.367
R966 B.n492 B.n31 163.367
R967 B.n488 B.n31 163.367
R968 B.n488 B.n487 163.367
R969 B.n487 B.n486 163.367
R970 B.n486 B.n33 163.367
R971 B.n482 B.n33 163.367
R972 B.n482 B.n481 163.367
R973 B.n481 B.n480 163.367
R974 B.n480 B.n35 163.367
R975 B.n475 B.n35 163.367
R976 B.n475 B.n474 163.367
R977 B.n474 B.n473 163.367
R978 B.n473 B.n39 163.367
R979 B.n469 B.n39 163.367
R980 B.n469 B.n468 163.367
R981 B.n468 B.n467 163.367
R982 B.n467 B.n41 163.367
R983 B.n462 B.n41 163.367
R984 B.n462 B.n461 163.367
R985 B.n461 B.n460 163.367
R986 B.n460 B.n45 163.367
R987 B.n456 B.n45 163.367
R988 B.n456 B.n455 163.367
R989 B.n455 B.n454 163.367
R990 B.n454 B.n47 163.367
R991 B.n450 B.n47 163.367
R992 B.n450 B.n449 163.367
R993 B.n449 B.n448 163.367
R994 B.n448 B.n49 163.367
R995 B.n444 B.n49 163.367
R996 B.n444 B.n443 163.367
R997 B.n443 B.n442 163.367
R998 B.n442 B.n51 163.367
R999 B.n438 B.n51 163.367
R1000 B.n438 B.n437 163.367
R1001 B.n437 B.n436 163.367
R1002 B.n436 B.n53 163.367
R1003 B.n112 B.n111 59.5399
R1004 B.n249 B.n119 59.5399
R1005 B.n478 B.n37 59.5399
R1006 B.n464 B.n43 59.5399
R1007 B.n111 B.n110 49.8429
R1008 B.n119 B.n118 49.8429
R1009 B.n37 B.n36 49.8429
R1010 B.n43 B.n42 49.8429
R1011 B.n509 B.n508 30.1273
R1012 B.n434 B.n433 30.1273
R1013 B.n295 B.n100 30.1273
R1014 B.n219 B.n218 30.1273
R1015 B B.n579 18.0485
R1016 B.n508 B.n507 10.6151
R1017 B.n507 B.n26 10.6151
R1018 B.n503 B.n26 10.6151
R1019 B.n503 B.n502 10.6151
R1020 B.n502 B.n501 10.6151
R1021 B.n501 B.n28 10.6151
R1022 B.n497 B.n28 10.6151
R1023 B.n497 B.n496 10.6151
R1024 B.n496 B.n495 10.6151
R1025 B.n495 B.n30 10.6151
R1026 B.n491 B.n30 10.6151
R1027 B.n491 B.n490 10.6151
R1028 B.n490 B.n489 10.6151
R1029 B.n489 B.n32 10.6151
R1030 B.n485 B.n32 10.6151
R1031 B.n485 B.n484 10.6151
R1032 B.n484 B.n483 10.6151
R1033 B.n483 B.n34 10.6151
R1034 B.n479 B.n34 10.6151
R1035 B.n477 B.n476 10.6151
R1036 B.n476 B.n38 10.6151
R1037 B.n472 B.n38 10.6151
R1038 B.n472 B.n471 10.6151
R1039 B.n471 B.n470 10.6151
R1040 B.n470 B.n40 10.6151
R1041 B.n466 B.n40 10.6151
R1042 B.n466 B.n465 10.6151
R1043 B.n463 B.n44 10.6151
R1044 B.n459 B.n44 10.6151
R1045 B.n459 B.n458 10.6151
R1046 B.n458 B.n457 10.6151
R1047 B.n457 B.n46 10.6151
R1048 B.n453 B.n46 10.6151
R1049 B.n453 B.n452 10.6151
R1050 B.n452 B.n451 10.6151
R1051 B.n451 B.n48 10.6151
R1052 B.n447 B.n48 10.6151
R1053 B.n447 B.n446 10.6151
R1054 B.n446 B.n445 10.6151
R1055 B.n445 B.n50 10.6151
R1056 B.n441 B.n50 10.6151
R1057 B.n441 B.n440 10.6151
R1058 B.n440 B.n439 10.6151
R1059 B.n439 B.n52 10.6151
R1060 B.n435 B.n52 10.6151
R1061 B.n435 B.n434 10.6151
R1062 B.n296 B.n295 10.6151
R1063 B.n297 B.n296 10.6151
R1064 B.n297 B.n98 10.6151
R1065 B.n301 B.n98 10.6151
R1066 B.n302 B.n301 10.6151
R1067 B.n303 B.n302 10.6151
R1068 B.n303 B.n96 10.6151
R1069 B.n307 B.n96 10.6151
R1070 B.n308 B.n307 10.6151
R1071 B.n309 B.n308 10.6151
R1072 B.n309 B.n94 10.6151
R1073 B.n313 B.n94 10.6151
R1074 B.n314 B.n313 10.6151
R1075 B.n315 B.n314 10.6151
R1076 B.n315 B.n92 10.6151
R1077 B.n319 B.n92 10.6151
R1078 B.n320 B.n319 10.6151
R1079 B.n321 B.n320 10.6151
R1080 B.n321 B.n90 10.6151
R1081 B.n325 B.n90 10.6151
R1082 B.n326 B.n325 10.6151
R1083 B.n327 B.n326 10.6151
R1084 B.n327 B.n88 10.6151
R1085 B.n331 B.n88 10.6151
R1086 B.n332 B.n331 10.6151
R1087 B.n333 B.n332 10.6151
R1088 B.n333 B.n86 10.6151
R1089 B.n337 B.n86 10.6151
R1090 B.n338 B.n337 10.6151
R1091 B.n339 B.n338 10.6151
R1092 B.n339 B.n84 10.6151
R1093 B.n343 B.n84 10.6151
R1094 B.n344 B.n343 10.6151
R1095 B.n345 B.n344 10.6151
R1096 B.n345 B.n82 10.6151
R1097 B.n349 B.n82 10.6151
R1098 B.n350 B.n349 10.6151
R1099 B.n351 B.n350 10.6151
R1100 B.n351 B.n80 10.6151
R1101 B.n355 B.n80 10.6151
R1102 B.n356 B.n355 10.6151
R1103 B.n357 B.n356 10.6151
R1104 B.n357 B.n78 10.6151
R1105 B.n361 B.n78 10.6151
R1106 B.n362 B.n361 10.6151
R1107 B.n363 B.n362 10.6151
R1108 B.n363 B.n76 10.6151
R1109 B.n367 B.n76 10.6151
R1110 B.n368 B.n367 10.6151
R1111 B.n369 B.n368 10.6151
R1112 B.n369 B.n74 10.6151
R1113 B.n373 B.n74 10.6151
R1114 B.n374 B.n373 10.6151
R1115 B.n375 B.n374 10.6151
R1116 B.n375 B.n72 10.6151
R1117 B.n379 B.n72 10.6151
R1118 B.n380 B.n379 10.6151
R1119 B.n381 B.n380 10.6151
R1120 B.n381 B.n70 10.6151
R1121 B.n385 B.n70 10.6151
R1122 B.n386 B.n385 10.6151
R1123 B.n387 B.n386 10.6151
R1124 B.n387 B.n68 10.6151
R1125 B.n391 B.n68 10.6151
R1126 B.n392 B.n391 10.6151
R1127 B.n393 B.n392 10.6151
R1128 B.n393 B.n66 10.6151
R1129 B.n397 B.n66 10.6151
R1130 B.n398 B.n397 10.6151
R1131 B.n399 B.n398 10.6151
R1132 B.n399 B.n64 10.6151
R1133 B.n403 B.n64 10.6151
R1134 B.n404 B.n403 10.6151
R1135 B.n405 B.n404 10.6151
R1136 B.n405 B.n62 10.6151
R1137 B.n409 B.n62 10.6151
R1138 B.n410 B.n409 10.6151
R1139 B.n411 B.n410 10.6151
R1140 B.n411 B.n60 10.6151
R1141 B.n415 B.n60 10.6151
R1142 B.n416 B.n415 10.6151
R1143 B.n417 B.n416 10.6151
R1144 B.n417 B.n58 10.6151
R1145 B.n421 B.n58 10.6151
R1146 B.n422 B.n421 10.6151
R1147 B.n423 B.n422 10.6151
R1148 B.n423 B.n56 10.6151
R1149 B.n427 B.n56 10.6151
R1150 B.n428 B.n427 10.6151
R1151 B.n429 B.n428 10.6151
R1152 B.n429 B.n54 10.6151
R1153 B.n433 B.n54 10.6151
R1154 B.n219 B.n128 10.6151
R1155 B.n223 B.n128 10.6151
R1156 B.n224 B.n223 10.6151
R1157 B.n225 B.n224 10.6151
R1158 B.n225 B.n126 10.6151
R1159 B.n229 B.n126 10.6151
R1160 B.n230 B.n229 10.6151
R1161 B.n231 B.n230 10.6151
R1162 B.n231 B.n124 10.6151
R1163 B.n235 B.n124 10.6151
R1164 B.n236 B.n235 10.6151
R1165 B.n237 B.n236 10.6151
R1166 B.n237 B.n122 10.6151
R1167 B.n241 B.n122 10.6151
R1168 B.n242 B.n241 10.6151
R1169 B.n243 B.n242 10.6151
R1170 B.n243 B.n120 10.6151
R1171 B.n247 B.n120 10.6151
R1172 B.n248 B.n247 10.6151
R1173 B.n250 B.n116 10.6151
R1174 B.n254 B.n116 10.6151
R1175 B.n255 B.n254 10.6151
R1176 B.n256 B.n255 10.6151
R1177 B.n256 B.n114 10.6151
R1178 B.n260 B.n114 10.6151
R1179 B.n261 B.n260 10.6151
R1180 B.n262 B.n261 10.6151
R1181 B.n266 B.n265 10.6151
R1182 B.n267 B.n266 10.6151
R1183 B.n267 B.n108 10.6151
R1184 B.n271 B.n108 10.6151
R1185 B.n272 B.n271 10.6151
R1186 B.n273 B.n272 10.6151
R1187 B.n273 B.n106 10.6151
R1188 B.n277 B.n106 10.6151
R1189 B.n278 B.n277 10.6151
R1190 B.n279 B.n278 10.6151
R1191 B.n279 B.n104 10.6151
R1192 B.n283 B.n104 10.6151
R1193 B.n284 B.n283 10.6151
R1194 B.n285 B.n284 10.6151
R1195 B.n285 B.n102 10.6151
R1196 B.n289 B.n102 10.6151
R1197 B.n290 B.n289 10.6151
R1198 B.n291 B.n290 10.6151
R1199 B.n291 B.n100 10.6151
R1200 B.n218 B.n217 10.6151
R1201 B.n217 B.n130 10.6151
R1202 B.n213 B.n130 10.6151
R1203 B.n213 B.n212 10.6151
R1204 B.n212 B.n211 10.6151
R1205 B.n211 B.n132 10.6151
R1206 B.n207 B.n132 10.6151
R1207 B.n207 B.n206 10.6151
R1208 B.n206 B.n205 10.6151
R1209 B.n205 B.n134 10.6151
R1210 B.n201 B.n134 10.6151
R1211 B.n201 B.n200 10.6151
R1212 B.n200 B.n199 10.6151
R1213 B.n199 B.n136 10.6151
R1214 B.n195 B.n136 10.6151
R1215 B.n195 B.n194 10.6151
R1216 B.n194 B.n193 10.6151
R1217 B.n193 B.n138 10.6151
R1218 B.n189 B.n138 10.6151
R1219 B.n189 B.n188 10.6151
R1220 B.n188 B.n187 10.6151
R1221 B.n187 B.n140 10.6151
R1222 B.n183 B.n140 10.6151
R1223 B.n183 B.n182 10.6151
R1224 B.n182 B.n181 10.6151
R1225 B.n181 B.n142 10.6151
R1226 B.n177 B.n142 10.6151
R1227 B.n177 B.n176 10.6151
R1228 B.n176 B.n175 10.6151
R1229 B.n175 B.n144 10.6151
R1230 B.n171 B.n144 10.6151
R1231 B.n171 B.n170 10.6151
R1232 B.n170 B.n169 10.6151
R1233 B.n169 B.n146 10.6151
R1234 B.n165 B.n146 10.6151
R1235 B.n165 B.n164 10.6151
R1236 B.n164 B.n163 10.6151
R1237 B.n163 B.n148 10.6151
R1238 B.n159 B.n148 10.6151
R1239 B.n159 B.n158 10.6151
R1240 B.n158 B.n157 10.6151
R1241 B.n157 B.n150 10.6151
R1242 B.n153 B.n150 10.6151
R1243 B.n153 B.n152 10.6151
R1244 B.n152 B.n0 10.6151
R1245 B.n575 B.n1 10.6151
R1246 B.n575 B.n574 10.6151
R1247 B.n574 B.n573 10.6151
R1248 B.n573 B.n4 10.6151
R1249 B.n569 B.n4 10.6151
R1250 B.n569 B.n568 10.6151
R1251 B.n568 B.n567 10.6151
R1252 B.n567 B.n6 10.6151
R1253 B.n563 B.n6 10.6151
R1254 B.n563 B.n562 10.6151
R1255 B.n562 B.n561 10.6151
R1256 B.n561 B.n8 10.6151
R1257 B.n557 B.n8 10.6151
R1258 B.n557 B.n556 10.6151
R1259 B.n556 B.n555 10.6151
R1260 B.n555 B.n10 10.6151
R1261 B.n551 B.n10 10.6151
R1262 B.n551 B.n550 10.6151
R1263 B.n550 B.n549 10.6151
R1264 B.n549 B.n12 10.6151
R1265 B.n545 B.n12 10.6151
R1266 B.n545 B.n544 10.6151
R1267 B.n544 B.n543 10.6151
R1268 B.n543 B.n14 10.6151
R1269 B.n539 B.n14 10.6151
R1270 B.n539 B.n538 10.6151
R1271 B.n538 B.n537 10.6151
R1272 B.n537 B.n16 10.6151
R1273 B.n533 B.n16 10.6151
R1274 B.n533 B.n532 10.6151
R1275 B.n532 B.n531 10.6151
R1276 B.n531 B.n18 10.6151
R1277 B.n527 B.n18 10.6151
R1278 B.n527 B.n526 10.6151
R1279 B.n526 B.n525 10.6151
R1280 B.n525 B.n20 10.6151
R1281 B.n521 B.n20 10.6151
R1282 B.n521 B.n520 10.6151
R1283 B.n520 B.n519 10.6151
R1284 B.n519 B.n22 10.6151
R1285 B.n515 B.n22 10.6151
R1286 B.n515 B.n514 10.6151
R1287 B.n514 B.n513 10.6151
R1288 B.n513 B.n24 10.6151
R1289 B.n509 B.n24 10.6151
R1290 B.n478 B.n477 6.5566
R1291 B.n465 B.n464 6.5566
R1292 B.n250 B.n249 6.5566
R1293 B.n262 B.n112 6.5566
R1294 B.n479 B.n478 4.05904
R1295 B.n464 B.n463 4.05904
R1296 B.n249 B.n248 4.05904
R1297 B.n265 B.n112 4.05904
R1298 B.n579 B.n0 2.81026
R1299 B.n579 B.n1 2.81026
R1300 VN.n47 VN.n25 161.3
R1301 VN.n46 VN.n45 161.3
R1302 VN.n44 VN.n26 161.3
R1303 VN.n43 VN.n42 161.3
R1304 VN.n41 VN.n27 161.3
R1305 VN.n39 VN.n38 161.3
R1306 VN.n37 VN.n28 161.3
R1307 VN.n36 VN.n35 161.3
R1308 VN.n34 VN.n29 161.3
R1309 VN.n33 VN.n32 161.3
R1310 VN.n22 VN.n0 161.3
R1311 VN.n21 VN.n20 161.3
R1312 VN.n19 VN.n1 161.3
R1313 VN.n18 VN.n17 161.3
R1314 VN.n16 VN.n2 161.3
R1315 VN.n14 VN.n13 161.3
R1316 VN.n12 VN.n3 161.3
R1317 VN.n11 VN.n10 161.3
R1318 VN.n9 VN.n4 161.3
R1319 VN.n8 VN.n7 161.3
R1320 VN.n24 VN.n23 93.3849
R1321 VN.n49 VN.n48 93.3849
R1322 VN.n6 VN.t4 81.9516
R1323 VN.n31 VN.t3 81.9516
R1324 VN.n6 VN.n5 57.3618
R1325 VN.n31 VN.n30 57.3618
R1326 VN.n5 VN.t6 48.5233
R1327 VN.n15 VN.t7 48.5233
R1328 VN.n23 VN.t5 48.5233
R1329 VN.n30 VN.t1 48.5233
R1330 VN.n40 VN.t2 48.5233
R1331 VN.n48 VN.t0 48.5233
R1332 VN.n21 VN.n1 47.2923
R1333 VN.n46 VN.n26 47.2923
R1334 VN VN.n49 43.8618
R1335 VN.n10 VN.n9 40.4934
R1336 VN.n10 VN.n3 40.4934
R1337 VN.n35 VN.n34 40.4934
R1338 VN.n35 VN.n28 40.4934
R1339 VN.n17 VN.n1 33.6945
R1340 VN.n42 VN.n26 33.6945
R1341 VN.n9 VN.n8 24.4675
R1342 VN.n14 VN.n3 24.4675
R1343 VN.n17 VN.n16 24.4675
R1344 VN.n22 VN.n21 24.4675
R1345 VN.n34 VN.n33 24.4675
R1346 VN.n42 VN.n41 24.4675
R1347 VN.n39 VN.n28 24.4675
R1348 VN.n47 VN.n46 24.4675
R1349 VN.n23 VN.n22 17.3721
R1350 VN.n48 VN.n47 17.3721
R1351 VN.n8 VN.n5 13.9467
R1352 VN.n15 VN.n14 13.9467
R1353 VN.n33 VN.n30 13.9467
R1354 VN.n40 VN.n39 13.9467
R1355 VN.n16 VN.n15 10.5213
R1356 VN.n41 VN.n40 10.5213
R1357 VN.n32 VN.n31 9.22138
R1358 VN.n7 VN.n6 9.22138
R1359 VN.n49 VN.n25 0.278367
R1360 VN.n24 VN.n0 0.278367
R1361 VN.n45 VN.n25 0.189894
R1362 VN.n45 VN.n44 0.189894
R1363 VN.n44 VN.n43 0.189894
R1364 VN.n43 VN.n27 0.189894
R1365 VN.n38 VN.n27 0.189894
R1366 VN.n38 VN.n37 0.189894
R1367 VN.n37 VN.n36 0.189894
R1368 VN.n36 VN.n29 0.189894
R1369 VN.n32 VN.n29 0.189894
R1370 VN.n7 VN.n4 0.189894
R1371 VN.n11 VN.n4 0.189894
R1372 VN.n12 VN.n11 0.189894
R1373 VN.n13 VN.n12 0.189894
R1374 VN.n13 VN.n2 0.189894
R1375 VN.n18 VN.n2 0.189894
R1376 VN.n19 VN.n18 0.189894
R1377 VN.n20 VN.n19 0.189894
R1378 VN.n20 VN.n0 0.189894
R1379 VN VN.n24 0.153454
R1380 VDD2.n2 VDD2.n1 104.162
R1381 VDD2.n2 VDD2.n0 104.162
R1382 VDD2 VDD2.n5 104.159
R1383 VDD2.n4 VDD2.n3 103.111
R1384 VDD2.n4 VDD2.n2 37.5731
R1385 VDD2.n5 VDD2.t6 7.20782
R1386 VDD2.n5 VDD2.t4 7.20782
R1387 VDD2.n3 VDD2.t7 7.20782
R1388 VDD2.n3 VDD2.t5 7.20782
R1389 VDD2.n1 VDD2.t0 7.20782
R1390 VDD2.n1 VDD2.t2 7.20782
R1391 VDD2.n0 VDD2.t3 7.20782
R1392 VDD2.n0 VDD2.t1 7.20782
R1393 VDD2 VDD2.n4 1.16645
C0 VTAIL VDD2 5.37134f
C1 VTAIL VDD1 5.31934f
C2 VP w_n3540_n1870# 7.43224f
C3 VN VP 5.84007f
C4 VP VDD2 0.485595f
C5 VP VDD1 3.77698f
C6 VTAIL VP 4.23652f
C7 w_n3540_n1870# B 7.47734f
C8 VN B 1.07686f
C9 B VDD2 1.42363f
C10 B VDD1 1.33881f
C11 VN w_n3540_n1870# 6.97396f
C12 VTAIL B 2.38445f
C13 w_n3540_n1870# VDD2 1.73147f
C14 VN VDD2 3.44799f
C15 w_n3540_n1870# VDD1 1.63218f
C16 VN VDD1 0.154841f
C17 VDD1 VDD2 1.58822f
C18 VP B 1.84344f
C19 VTAIL w_n3540_n1870# 2.46007f
C20 VTAIL VN 4.22241f
C21 VDD2 VSUBS 1.412093f
C22 VDD1 VSUBS 2.006672f
C23 VTAIL VSUBS 0.622669f
C24 VN VSUBS 5.9794f
C25 VP VSUBS 2.711438f
C26 B VSUBS 3.746848f
C27 w_n3540_n1870# VSUBS 83.1334f
C28 VDD2.t3 VSUBS 0.08652f
C29 VDD2.t1 VSUBS 0.08652f
C30 VDD2.n0 VSUBS 0.531948f
C31 VDD2.t0 VSUBS 0.08652f
C32 VDD2.t2 VSUBS 0.08652f
C33 VDD2.n1 VSUBS 0.531948f
C34 VDD2.n2 VSUBS 2.85797f
C35 VDD2.t7 VSUBS 0.08652f
C36 VDD2.t5 VSUBS 0.08652f
C37 VDD2.n3 VSUBS 0.525632f
C38 VDD2.n4 VSUBS 2.33683f
C39 VDD2.t6 VSUBS 0.08652f
C40 VDD2.t4 VSUBS 0.08652f
C41 VDD2.n5 VSUBS 0.531923f
C42 VN.n0 VSUBS 0.055986f
C43 VN.t5 VSUBS 1.11339f
C44 VN.n1 VSUBS 0.037079f
C45 VN.n2 VSUBS 0.042465f
C46 VN.t7 VSUBS 1.11339f
C47 VN.n3 VSUBS 0.084399f
C48 VN.n4 VSUBS 0.042465f
C49 VN.t6 VSUBS 1.11339f
C50 VN.n5 VSUBS 0.553054f
C51 VN.t4 VSUBS 1.38907f
C52 VN.n6 VSUBS 0.532746f
C53 VN.n7 VSUBS 0.363181f
C54 VN.n8 VSUBS 0.06234f
C55 VN.n9 VSUBS 0.084399f
C56 VN.n10 VSUBS 0.034329f
C57 VN.n11 VSUBS 0.042465f
C58 VN.n12 VSUBS 0.042465f
C59 VN.n13 VSUBS 0.042465f
C60 VN.n14 VSUBS 0.06234f
C61 VN.n15 VSUBS 0.43982f
C62 VN.n16 VSUBS 0.05687f
C63 VN.n17 VSUBS 0.085775f
C64 VN.n18 VSUBS 0.042465f
C65 VN.n19 VSUBS 0.042465f
C66 VN.n20 VSUBS 0.042465f
C67 VN.n21 VSUBS 0.080272f
C68 VN.n22 VSUBS 0.06781f
C69 VN.n23 VSUBS 0.579027f
C70 VN.n24 VSUBS 0.056426f
C71 VN.n25 VSUBS 0.055986f
C72 VN.t0 VSUBS 1.11339f
C73 VN.n26 VSUBS 0.037079f
C74 VN.n27 VSUBS 0.042465f
C75 VN.t2 VSUBS 1.11339f
C76 VN.n28 VSUBS 0.084399f
C77 VN.n29 VSUBS 0.042465f
C78 VN.t1 VSUBS 1.11339f
C79 VN.n30 VSUBS 0.553054f
C80 VN.t3 VSUBS 1.38907f
C81 VN.n31 VSUBS 0.532746f
C82 VN.n32 VSUBS 0.363181f
C83 VN.n33 VSUBS 0.06234f
C84 VN.n34 VSUBS 0.084399f
C85 VN.n35 VSUBS 0.034329f
C86 VN.n36 VSUBS 0.042465f
C87 VN.n37 VSUBS 0.042465f
C88 VN.n38 VSUBS 0.042465f
C89 VN.n39 VSUBS 0.06234f
C90 VN.n40 VSUBS 0.43982f
C91 VN.n41 VSUBS 0.05687f
C92 VN.n42 VSUBS 0.085775f
C93 VN.n43 VSUBS 0.042465f
C94 VN.n44 VSUBS 0.042465f
C95 VN.n45 VSUBS 0.042465f
C96 VN.n46 VSUBS 0.080272f
C97 VN.n47 VSUBS 0.06781f
C98 VN.n48 VSUBS 0.579027f
C99 VN.n49 VSUBS 1.92761f
C100 B.n0 VSUBS 0.00562f
C101 B.n1 VSUBS 0.00562f
C102 B.n2 VSUBS 0.008888f
C103 B.n3 VSUBS 0.008888f
C104 B.n4 VSUBS 0.008888f
C105 B.n5 VSUBS 0.008888f
C106 B.n6 VSUBS 0.008888f
C107 B.n7 VSUBS 0.008888f
C108 B.n8 VSUBS 0.008888f
C109 B.n9 VSUBS 0.008888f
C110 B.n10 VSUBS 0.008888f
C111 B.n11 VSUBS 0.008888f
C112 B.n12 VSUBS 0.008888f
C113 B.n13 VSUBS 0.008888f
C114 B.n14 VSUBS 0.008888f
C115 B.n15 VSUBS 0.008888f
C116 B.n16 VSUBS 0.008888f
C117 B.n17 VSUBS 0.008888f
C118 B.n18 VSUBS 0.008888f
C119 B.n19 VSUBS 0.008888f
C120 B.n20 VSUBS 0.008888f
C121 B.n21 VSUBS 0.008888f
C122 B.n22 VSUBS 0.008888f
C123 B.n23 VSUBS 0.008888f
C124 B.n24 VSUBS 0.008888f
C125 B.n25 VSUBS 0.020306f
C126 B.n26 VSUBS 0.008888f
C127 B.n27 VSUBS 0.008888f
C128 B.n28 VSUBS 0.008888f
C129 B.n29 VSUBS 0.008888f
C130 B.n30 VSUBS 0.008888f
C131 B.n31 VSUBS 0.008888f
C132 B.n32 VSUBS 0.008888f
C133 B.n33 VSUBS 0.008888f
C134 B.n34 VSUBS 0.008888f
C135 B.n35 VSUBS 0.008888f
C136 B.t5 VSUBS 0.082442f
C137 B.t4 VSUBS 0.10747f
C138 B.t3 VSUBS 0.610431f
C139 B.n36 VSUBS 0.189495f
C140 B.n37 VSUBS 0.159526f
C141 B.n38 VSUBS 0.008888f
C142 B.n39 VSUBS 0.008888f
C143 B.n40 VSUBS 0.008888f
C144 B.n41 VSUBS 0.008888f
C145 B.t8 VSUBS 0.082443f
C146 B.t7 VSUBS 0.107471f
C147 B.t6 VSUBS 0.610431f
C148 B.n42 VSUBS 0.189494f
C149 B.n43 VSUBS 0.159524f
C150 B.n44 VSUBS 0.008888f
C151 B.n45 VSUBS 0.008888f
C152 B.n46 VSUBS 0.008888f
C153 B.n47 VSUBS 0.008888f
C154 B.n48 VSUBS 0.008888f
C155 B.n49 VSUBS 0.008888f
C156 B.n50 VSUBS 0.008888f
C157 B.n51 VSUBS 0.008888f
C158 B.n52 VSUBS 0.008888f
C159 B.n53 VSUBS 0.020306f
C160 B.n54 VSUBS 0.008888f
C161 B.n55 VSUBS 0.008888f
C162 B.n56 VSUBS 0.008888f
C163 B.n57 VSUBS 0.008888f
C164 B.n58 VSUBS 0.008888f
C165 B.n59 VSUBS 0.008888f
C166 B.n60 VSUBS 0.008888f
C167 B.n61 VSUBS 0.008888f
C168 B.n62 VSUBS 0.008888f
C169 B.n63 VSUBS 0.008888f
C170 B.n64 VSUBS 0.008888f
C171 B.n65 VSUBS 0.008888f
C172 B.n66 VSUBS 0.008888f
C173 B.n67 VSUBS 0.008888f
C174 B.n68 VSUBS 0.008888f
C175 B.n69 VSUBS 0.008888f
C176 B.n70 VSUBS 0.008888f
C177 B.n71 VSUBS 0.008888f
C178 B.n72 VSUBS 0.008888f
C179 B.n73 VSUBS 0.008888f
C180 B.n74 VSUBS 0.008888f
C181 B.n75 VSUBS 0.008888f
C182 B.n76 VSUBS 0.008888f
C183 B.n77 VSUBS 0.008888f
C184 B.n78 VSUBS 0.008888f
C185 B.n79 VSUBS 0.008888f
C186 B.n80 VSUBS 0.008888f
C187 B.n81 VSUBS 0.008888f
C188 B.n82 VSUBS 0.008888f
C189 B.n83 VSUBS 0.008888f
C190 B.n84 VSUBS 0.008888f
C191 B.n85 VSUBS 0.008888f
C192 B.n86 VSUBS 0.008888f
C193 B.n87 VSUBS 0.008888f
C194 B.n88 VSUBS 0.008888f
C195 B.n89 VSUBS 0.008888f
C196 B.n90 VSUBS 0.008888f
C197 B.n91 VSUBS 0.008888f
C198 B.n92 VSUBS 0.008888f
C199 B.n93 VSUBS 0.008888f
C200 B.n94 VSUBS 0.008888f
C201 B.n95 VSUBS 0.008888f
C202 B.n96 VSUBS 0.008888f
C203 B.n97 VSUBS 0.008888f
C204 B.n98 VSUBS 0.008888f
C205 B.n99 VSUBS 0.008888f
C206 B.n100 VSUBS 0.020306f
C207 B.n101 VSUBS 0.008888f
C208 B.n102 VSUBS 0.008888f
C209 B.n103 VSUBS 0.008888f
C210 B.n104 VSUBS 0.008888f
C211 B.n105 VSUBS 0.008888f
C212 B.n106 VSUBS 0.008888f
C213 B.n107 VSUBS 0.008888f
C214 B.n108 VSUBS 0.008888f
C215 B.n109 VSUBS 0.008888f
C216 B.t10 VSUBS 0.082443f
C217 B.t11 VSUBS 0.107471f
C218 B.t9 VSUBS 0.610431f
C219 B.n110 VSUBS 0.189494f
C220 B.n111 VSUBS 0.159524f
C221 B.n112 VSUBS 0.020593f
C222 B.n113 VSUBS 0.008888f
C223 B.n114 VSUBS 0.008888f
C224 B.n115 VSUBS 0.008888f
C225 B.n116 VSUBS 0.008888f
C226 B.n117 VSUBS 0.008888f
C227 B.t1 VSUBS 0.082442f
C228 B.t2 VSUBS 0.10747f
C229 B.t0 VSUBS 0.610431f
C230 B.n118 VSUBS 0.189495f
C231 B.n119 VSUBS 0.159526f
C232 B.n120 VSUBS 0.008888f
C233 B.n121 VSUBS 0.008888f
C234 B.n122 VSUBS 0.008888f
C235 B.n123 VSUBS 0.008888f
C236 B.n124 VSUBS 0.008888f
C237 B.n125 VSUBS 0.008888f
C238 B.n126 VSUBS 0.008888f
C239 B.n127 VSUBS 0.008888f
C240 B.n128 VSUBS 0.008888f
C241 B.n129 VSUBS 0.019168f
C242 B.n130 VSUBS 0.008888f
C243 B.n131 VSUBS 0.008888f
C244 B.n132 VSUBS 0.008888f
C245 B.n133 VSUBS 0.008888f
C246 B.n134 VSUBS 0.008888f
C247 B.n135 VSUBS 0.008888f
C248 B.n136 VSUBS 0.008888f
C249 B.n137 VSUBS 0.008888f
C250 B.n138 VSUBS 0.008888f
C251 B.n139 VSUBS 0.008888f
C252 B.n140 VSUBS 0.008888f
C253 B.n141 VSUBS 0.008888f
C254 B.n142 VSUBS 0.008888f
C255 B.n143 VSUBS 0.008888f
C256 B.n144 VSUBS 0.008888f
C257 B.n145 VSUBS 0.008888f
C258 B.n146 VSUBS 0.008888f
C259 B.n147 VSUBS 0.008888f
C260 B.n148 VSUBS 0.008888f
C261 B.n149 VSUBS 0.008888f
C262 B.n150 VSUBS 0.008888f
C263 B.n151 VSUBS 0.008888f
C264 B.n152 VSUBS 0.008888f
C265 B.n153 VSUBS 0.008888f
C266 B.n154 VSUBS 0.008888f
C267 B.n155 VSUBS 0.008888f
C268 B.n156 VSUBS 0.008888f
C269 B.n157 VSUBS 0.008888f
C270 B.n158 VSUBS 0.008888f
C271 B.n159 VSUBS 0.008888f
C272 B.n160 VSUBS 0.008888f
C273 B.n161 VSUBS 0.008888f
C274 B.n162 VSUBS 0.008888f
C275 B.n163 VSUBS 0.008888f
C276 B.n164 VSUBS 0.008888f
C277 B.n165 VSUBS 0.008888f
C278 B.n166 VSUBS 0.008888f
C279 B.n167 VSUBS 0.008888f
C280 B.n168 VSUBS 0.008888f
C281 B.n169 VSUBS 0.008888f
C282 B.n170 VSUBS 0.008888f
C283 B.n171 VSUBS 0.008888f
C284 B.n172 VSUBS 0.008888f
C285 B.n173 VSUBS 0.008888f
C286 B.n174 VSUBS 0.008888f
C287 B.n175 VSUBS 0.008888f
C288 B.n176 VSUBS 0.008888f
C289 B.n177 VSUBS 0.008888f
C290 B.n178 VSUBS 0.008888f
C291 B.n179 VSUBS 0.008888f
C292 B.n180 VSUBS 0.008888f
C293 B.n181 VSUBS 0.008888f
C294 B.n182 VSUBS 0.008888f
C295 B.n183 VSUBS 0.008888f
C296 B.n184 VSUBS 0.008888f
C297 B.n185 VSUBS 0.008888f
C298 B.n186 VSUBS 0.008888f
C299 B.n187 VSUBS 0.008888f
C300 B.n188 VSUBS 0.008888f
C301 B.n189 VSUBS 0.008888f
C302 B.n190 VSUBS 0.008888f
C303 B.n191 VSUBS 0.008888f
C304 B.n192 VSUBS 0.008888f
C305 B.n193 VSUBS 0.008888f
C306 B.n194 VSUBS 0.008888f
C307 B.n195 VSUBS 0.008888f
C308 B.n196 VSUBS 0.008888f
C309 B.n197 VSUBS 0.008888f
C310 B.n198 VSUBS 0.008888f
C311 B.n199 VSUBS 0.008888f
C312 B.n200 VSUBS 0.008888f
C313 B.n201 VSUBS 0.008888f
C314 B.n202 VSUBS 0.008888f
C315 B.n203 VSUBS 0.008888f
C316 B.n204 VSUBS 0.008888f
C317 B.n205 VSUBS 0.008888f
C318 B.n206 VSUBS 0.008888f
C319 B.n207 VSUBS 0.008888f
C320 B.n208 VSUBS 0.008888f
C321 B.n209 VSUBS 0.008888f
C322 B.n210 VSUBS 0.008888f
C323 B.n211 VSUBS 0.008888f
C324 B.n212 VSUBS 0.008888f
C325 B.n213 VSUBS 0.008888f
C326 B.n214 VSUBS 0.008888f
C327 B.n215 VSUBS 0.008888f
C328 B.n216 VSUBS 0.008888f
C329 B.n217 VSUBS 0.008888f
C330 B.n218 VSUBS 0.019168f
C331 B.n219 VSUBS 0.020306f
C332 B.n220 VSUBS 0.020306f
C333 B.n221 VSUBS 0.008888f
C334 B.n222 VSUBS 0.008888f
C335 B.n223 VSUBS 0.008888f
C336 B.n224 VSUBS 0.008888f
C337 B.n225 VSUBS 0.008888f
C338 B.n226 VSUBS 0.008888f
C339 B.n227 VSUBS 0.008888f
C340 B.n228 VSUBS 0.008888f
C341 B.n229 VSUBS 0.008888f
C342 B.n230 VSUBS 0.008888f
C343 B.n231 VSUBS 0.008888f
C344 B.n232 VSUBS 0.008888f
C345 B.n233 VSUBS 0.008888f
C346 B.n234 VSUBS 0.008888f
C347 B.n235 VSUBS 0.008888f
C348 B.n236 VSUBS 0.008888f
C349 B.n237 VSUBS 0.008888f
C350 B.n238 VSUBS 0.008888f
C351 B.n239 VSUBS 0.008888f
C352 B.n240 VSUBS 0.008888f
C353 B.n241 VSUBS 0.008888f
C354 B.n242 VSUBS 0.008888f
C355 B.n243 VSUBS 0.008888f
C356 B.n244 VSUBS 0.008888f
C357 B.n245 VSUBS 0.008888f
C358 B.n246 VSUBS 0.008888f
C359 B.n247 VSUBS 0.008888f
C360 B.n248 VSUBS 0.006143f
C361 B.n249 VSUBS 0.020593f
C362 B.n250 VSUBS 0.007189f
C363 B.n251 VSUBS 0.008888f
C364 B.n252 VSUBS 0.008888f
C365 B.n253 VSUBS 0.008888f
C366 B.n254 VSUBS 0.008888f
C367 B.n255 VSUBS 0.008888f
C368 B.n256 VSUBS 0.008888f
C369 B.n257 VSUBS 0.008888f
C370 B.n258 VSUBS 0.008888f
C371 B.n259 VSUBS 0.008888f
C372 B.n260 VSUBS 0.008888f
C373 B.n261 VSUBS 0.008888f
C374 B.n262 VSUBS 0.007189f
C375 B.n263 VSUBS 0.008888f
C376 B.n264 VSUBS 0.008888f
C377 B.n265 VSUBS 0.006143f
C378 B.n266 VSUBS 0.008888f
C379 B.n267 VSUBS 0.008888f
C380 B.n268 VSUBS 0.008888f
C381 B.n269 VSUBS 0.008888f
C382 B.n270 VSUBS 0.008888f
C383 B.n271 VSUBS 0.008888f
C384 B.n272 VSUBS 0.008888f
C385 B.n273 VSUBS 0.008888f
C386 B.n274 VSUBS 0.008888f
C387 B.n275 VSUBS 0.008888f
C388 B.n276 VSUBS 0.008888f
C389 B.n277 VSUBS 0.008888f
C390 B.n278 VSUBS 0.008888f
C391 B.n279 VSUBS 0.008888f
C392 B.n280 VSUBS 0.008888f
C393 B.n281 VSUBS 0.008888f
C394 B.n282 VSUBS 0.008888f
C395 B.n283 VSUBS 0.008888f
C396 B.n284 VSUBS 0.008888f
C397 B.n285 VSUBS 0.008888f
C398 B.n286 VSUBS 0.008888f
C399 B.n287 VSUBS 0.008888f
C400 B.n288 VSUBS 0.008888f
C401 B.n289 VSUBS 0.008888f
C402 B.n290 VSUBS 0.008888f
C403 B.n291 VSUBS 0.008888f
C404 B.n292 VSUBS 0.008888f
C405 B.n293 VSUBS 0.020306f
C406 B.n294 VSUBS 0.019168f
C407 B.n295 VSUBS 0.019168f
C408 B.n296 VSUBS 0.008888f
C409 B.n297 VSUBS 0.008888f
C410 B.n298 VSUBS 0.008888f
C411 B.n299 VSUBS 0.008888f
C412 B.n300 VSUBS 0.008888f
C413 B.n301 VSUBS 0.008888f
C414 B.n302 VSUBS 0.008888f
C415 B.n303 VSUBS 0.008888f
C416 B.n304 VSUBS 0.008888f
C417 B.n305 VSUBS 0.008888f
C418 B.n306 VSUBS 0.008888f
C419 B.n307 VSUBS 0.008888f
C420 B.n308 VSUBS 0.008888f
C421 B.n309 VSUBS 0.008888f
C422 B.n310 VSUBS 0.008888f
C423 B.n311 VSUBS 0.008888f
C424 B.n312 VSUBS 0.008888f
C425 B.n313 VSUBS 0.008888f
C426 B.n314 VSUBS 0.008888f
C427 B.n315 VSUBS 0.008888f
C428 B.n316 VSUBS 0.008888f
C429 B.n317 VSUBS 0.008888f
C430 B.n318 VSUBS 0.008888f
C431 B.n319 VSUBS 0.008888f
C432 B.n320 VSUBS 0.008888f
C433 B.n321 VSUBS 0.008888f
C434 B.n322 VSUBS 0.008888f
C435 B.n323 VSUBS 0.008888f
C436 B.n324 VSUBS 0.008888f
C437 B.n325 VSUBS 0.008888f
C438 B.n326 VSUBS 0.008888f
C439 B.n327 VSUBS 0.008888f
C440 B.n328 VSUBS 0.008888f
C441 B.n329 VSUBS 0.008888f
C442 B.n330 VSUBS 0.008888f
C443 B.n331 VSUBS 0.008888f
C444 B.n332 VSUBS 0.008888f
C445 B.n333 VSUBS 0.008888f
C446 B.n334 VSUBS 0.008888f
C447 B.n335 VSUBS 0.008888f
C448 B.n336 VSUBS 0.008888f
C449 B.n337 VSUBS 0.008888f
C450 B.n338 VSUBS 0.008888f
C451 B.n339 VSUBS 0.008888f
C452 B.n340 VSUBS 0.008888f
C453 B.n341 VSUBS 0.008888f
C454 B.n342 VSUBS 0.008888f
C455 B.n343 VSUBS 0.008888f
C456 B.n344 VSUBS 0.008888f
C457 B.n345 VSUBS 0.008888f
C458 B.n346 VSUBS 0.008888f
C459 B.n347 VSUBS 0.008888f
C460 B.n348 VSUBS 0.008888f
C461 B.n349 VSUBS 0.008888f
C462 B.n350 VSUBS 0.008888f
C463 B.n351 VSUBS 0.008888f
C464 B.n352 VSUBS 0.008888f
C465 B.n353 VSUBS 0.008888f
C466 B.n354 VSUBS 0.008888f
C467 B.n355 VSUBS 0.008888f
C468 B.n356 VSUBS 0.008888f
C469 B.n357 VSUBS 0.008888f
C470 B.n358 VSUBS 0.008888f
C471 B.n359 VSUBS 0.008888f
C472 B.n360 VSUBS 0.008888f
C473 B.n361 VSUBS 0.008888f
C474 B.n362 VSUBS 0.008888f
C475 B.n363 VSUBS 0.008888f
C476 B.n364 VSUBS 0.008888f
C477 B.n365 VSUBS 0.008888f
C478 B.n366 VSUBS 0.008888f
C479 B.n367 VSUBS 0.008888f
C480 B.n368 VSUBS 0.008888f
C481 B.n369 VSUBS 0.008888f
C482 B.n370 VSUBS 0.008888f
C483 B.n371 VSUBS 0.008888f
C484 B.n372 VSUBS 0.008888f
C485 B.n373 VSUBS 0.008888f
C486 B.n374 VSUBS 0.008888f
C487 B.n375 VSUBS 0.008888f
C488 B.n376 VSUBS 0.008888f
C489 B.n377 VSUBS 0.008888f
C490 B.n378 VSUBS 0.008888f
C491 B.n379 VSUBS 0.008888f
C492 B.n380 VSUBS 0.008888f
C493 B.n381 VSUBS 0.008888f
C494 B.n382 VSUBS 0.008888f
C495 B.n383 VSUBS 0.008888f
C496 B.n384 VSUBS 0.008888f
C497 B.n385 VSUBS 0.008888f
C498 B.n386 VSUBS 0.008888f
C499 B.n387 VSUBS 0.008888f
C500 B.n388 VSUBS 0.008888f
C501 B.n389 VSUBS 0.008888f
C502 B.n390 VSUBS 0.008888f
C503 B.n391 VSUBS 0.008888f
C504 B.n392 VSUBS 0.008888f
C505 B.n393 VSUBS 0.008888f
C506 B.n394 VSUBS 0.008888f
C507 B.n395 VSUBS 0.008888f
C508 B.n396 VSUBS 0.008888f
C509 B.n397 VSUBS 0.008888f
C510 B.n398 VSUBS 0.008888f
C511 B.n399 VSUBS 0.008888f
C512 B.n400 VSUBS 0.008888f
C513 B.n401 VSUBS 0.008888f
C514 B.n402 VSUBS 0.008888f
C515 B.n403 VSUBS 0.008888f
C516 B.n404 VSUBS 0.008888f
C517 B.n405 VSUBS 0.008888f
C518 B.n406 VSUBS 0.008888f
C519 B.n407 VSUBS 0.008888f
C520 B.n408 VSUBS 0.008888f
C521 B.n409 VSUBS 0.008888f
C522 B.n410 VSUBS 0.008888f
C523 B.n411 VSUBS 0.008888f
C524 B.n412 VSUBS 0.008888f
C525 B.n413 VSUBS 0.008888f
C526 B.n414 VSUBS 0.008888f
C527 B.n415 VSUBS 0.008888f
C528 B.n416 VSUBS 0.008888f
C529 B.n417 VSUBS 0.008888f
C530 B.n418 VSUBS 0.008888f
C531 B.n419 VSUBS 0.008888f
C532 B.n420 VSUBS 0.008888f
C533 B.n421 VSUBS 0.008888f
C534 B.n422 VSUBS 0.008888f
C535 B.n423 VSUBS 0.008888f
C536 B.n424 VSUBS 0.008888f
C537 B.n425 VSUBS 0.008888f
C538 B.n426 VSUBS 0.008888f
C539 B.n427 VSUBS 0.008888f
C540 B.n428 VSUBS 0.008888f
C541 B.n429 VSUBS 0.008888f
C542 B.n430 VSUBS 0.008888f
C543 B.n431 VSUBS 0.008888f
C544 B.n432 VSUBS 0.019168f
C545 B.n433 VSUBS 0.020306f
C546 B.n434 VSUBS 0.019168f
C547 B.n435 VSUBS 0.008888f
C548 B.n436 VSUBS 0.008888f
C549 B.n437 VSUBS 0.008888f
C550 B.n438 VSUBS 0.008888f
C551 B.n439 VSUBS 0.008888f
C552 B.n440 VSUBS 0.008888f
C553 B.n441 VSUBS 0.008888f
C554 B.n442 VSUBS 0.008888f
C555 B.n443 VSUBS 0.008888f
C556 B.n444 VSUBS 0.008888f
C557 B.n445 VSUBS 0.008888f
C558 B.n446 VSUBS 0.008888f
C559 B.n447 VSUBS 0.008888f
C560 B.n448 VSUBS 0.008888f
C561 B.n449 VSUBS 0.008888f
C562 B.n450 VSUBS 0.008888f
C563 B.n451 VSUBS 0.008888f
C564 B.n452 VSUBS 0.008888f
C565 B.n453 VSUBS 0.008888f
C566 B.n454 VSUBS 0.008888f
C567 B.n455 VSUBS 0.008888f
C568 B.n456 VSUBS 0.008888f
C569 B.n457 VSUBS 0.008888f
C570 B.n458 VSUBS 0.008888f
C571 B.n459 VSUBS 0.008888f
C572 B.n460 VSUBS 0.008888f
C573 B.n461 VSUBS 0.008888f
C574 B.n462 VSUBS 0.008888f
C575 B.n463 VSUBS 0.006143f
C576 B.n464 VSUBS 0.020593f
C577 B.n465 VSUBS 0.007189f
C578 B.n466 VSUBS 0.008888f
C579 B.n467 VSUBS 0.008888f
C580 B.n468 VSUBS 0.008888f
C581 B.n469 VSUBS 0.008888f
C582 B.n470 VSUBS 0.008888f
C583 B.n471 VSUBS 0.008888f
C584 B.n472 VSUBS 0.008888f
C585 B.n473 VSUBS 0.008888f
C586 B.n474 VSUBS 0.008888f
C587 B.n475 VSUBS 0.008888f
C588 B.n476 VSUBS 0.008888f
C589 B.n477 VSUBS 0.007189f
C590 B.n478 VSUBS 0.020593f
C591 B.n479 VSUBS 0.006143f
C592 B.n480 VSUBS 0.008888f
C593 B.n481 VSUBS 0.008888f
C594 B.n482 VSUBS 0.008888f
C595 B.n483 VSUBS 0.008888f
C596 B.n484 VSUBS 0.008888f
C597 B.n485 VSUBS 0.008888f
C598 B.n486 VSUBS 0.008888f
C599 B.n487 VSUBS 0.008888f
C600 B.n488 VSUBS 0.008888f
C601 B.n489 VSUBS 0.008888f
C602 B.n490 VSUBS 0.008888f
C603 B.n491 VSUBS 0.008888f
C604 B.n492 VSUBS 0.008888f
C605 B.n493 VSUBS 0.008888f
C606 B.n494 VSUBS 0.008888f
C607 B.n495 VSUBS 0.008888f
C608 B.n496 VSUBS 0.008888f
C609 B.n497 VSUBS 0.008888f
C610 B.n498 VSUBS 0.008888f
C611 B.n499 VSUBS 0.008888f
C612 B.n500 VSUBS 0.008888f
C613 B.n501 VSUBS 0.008888f
C614 B.n502 VSUBS 0.008888f
C615 B.n503 VSUBS 0.008888f
C616 B.n504 VSUBS 0.008888f
C617 B.n505 VSUBS 0.008888f
C618 B.n506 VSUBS 0.008888f
C619 B.n507 VSUBS 0.008888f
C620 B.n508 VSUBS 0.020306f
C621 B.n509 VSUBS 0.019168f
C622 B.n510 VSUBS 0.019168f
C623 B.n511 VSUBS 0.008888f
C624 B.n512 VSUBS 0.008888f
C625 B.n513 VSUBS 0.008888f
C626 B.n514 VSUBS 0.008888f
C627 B.n515 VSUBS 0.008888f
C628 B.n516 VSUBS 0.008888f
C629 B.n517 VSUBS 0.008888f
C630 B.n518 VSUBS 0.008888f
C631 B.n519 VSUBS 0.008888f
C632 B.n520 VSUBS 0.008888f
C633 B.n521 VSUBS 0.008888f
C634 B.n522 VSUBS 0.008888f
C635 B.n523 VSUBS 0.008888f
C636 B.n524 VSUBS 0.008888f
C637 B.n525 VSUBS 0.008888f
C638 B.n526 VSUBS 0.008888f
C639 B.n527 VSUBS 0.008888f
C640 B.n528 VSUBS 0.008888f
C641 B.n529 VSUBS 0.008888f
C642 B.n530 VSUBS 0.008888f
C643 B.n531 VSUBS 0.008888f
C644 B.n532 VSUBS 0.008888f
C645 B.n533 VSUBS 0.008888f
C646 B.n534 VSUBS 0.008888f
C647 B.n535 VSUBS 0.008888f
C648 B.n536 VSUBS 0.008888f
C649 B.n537 VSUBS 0.008888f
C650 B.n538 VSUBS 0.008888f
C651 B.n539 VSUBS 0.008888f
C652 B.n540 VSUBS 0.008888f
C653 B.n541 VSUBS 0.008888f
C654 B.n542 VSUBS 0.008888f
C655 B.n543 VSUBS 0.008888f
C656 B.n544 VSUBS 0.008888f
C657 B.n545 VSUBS 0.008888f
C658 B.n546 VSUBS 0.008888f
C659 B.n547 VSUBS 0.008888f
C660 B.n548 VSUBS 0.008888f
C661 B.n549 VSUBS 0.008888f
C662 B.n550 VSUBS 0.008888f
C663 B.n551 VSUBS 0.008888f
C664 B.n552 VSUBS 0.008888f
C665 B.n553 VSUBS 0.008888f
C666 B.n554 VSUBS 0.008888f
C667 B.n555 VSUBS 0.008888f
C668 B.n556 VSUBS 0.008888f
C669 B.n557 VSUBS 0.008888f
C670 B.n558 VSUBS 0.008888f
C671 B.n559 VSUBS 0.008888f
C672 B.n560 VSUBS 0.008888f
C673 B.n561 VSUBS 0.008888f
C674 B.n562 VSUBS 0.008888f
C675 B.n563 VSUBS 0.008888f
C676 B.n564 VSUBS 0.008888f
C677 B.n565 VSUBS 0.008888f
C678 B.n566 VSUBS 0.008888f
C679 B.n567 VSUBS 0.008888f
C680 B.n568 VSUBS 0.008888f
C681 B.n569 VSUBS 0.008888f
C682 B.n570 VSUBS 0.008888f
C683 B.n571 VSUBS 0.008888f
C684 B.n572 VSUBS 0.008888f
C685 B.n573 VSUBS 0.008888f
C686 B.n574 VSUBS 0.008888f
C687 B.n575 VSUBS 0.008888f
C688 B.n576 VSUBS 0.008888f
C689 B.n577 VSUBS 0.008888f
C690 B.n578 VSUBS 0.008888f
C691 B.n579 VSUBS 0.020126f
C692 VTAIL.t14 VSUBS 0.10956f
C693 VTAIL.t4 VSUBS 0.10956f
C694 VTAIL.n0 VSUBS 0.578914f
C695 VTAIL.n1 VSUBS 0.725224f
C696 VTAIL.n2 VSUBS 0.031955f
C697 VTAIL.n3 VSUBS 0.030741f
C698 VTAIL.n4 VSUBS 0.016519f
C699 VTAIL.n5 VSUBS 0.039045f
C700 VTAIL.n6 VSUBS 0.017491f
C701 VTAIL.n7 VSUBS 0.49589f
C702 VTAIL.n8 VSUBS 0.016519f
C703 VTAIL.t0 VSUBS 0.084543f
C704 VTAIL.n9 VSUBS 0.122977f
C705 VTAIL.n10 VSUBS 0.024736f
C706 VTAIL.n11 VSUBS 0.029284f
C707 VTAIL.n12 VSUBS 0.039045f
C708 VTAIL.n13 VSUBS 0.017491f
C709 VTAIL.n14 VSUBS 0.016519f
C710 VTAIL.n15 VSUBS 0.030741f
C711 VTAIL.n16 VSUBS 0.030741f
C712 VTAIL.n17 VSUBS 0.016519f
C713 VTAIL.n18 VSUBS 0.017491f
C714 VTAIL.n19 VSUBS 0.039045f
C715 VTAIL.n20 VSUBS 0.088315f
C716 VTAIL.n21 VSUBS 0.017491f
C717 VTAIL.n22 VSUBS 0.016519f
C718 VTAIL.n23 VSUBS 0.068957f
C719 VTAIL.n24 VSUBS 0.044072f
C720 VTAIL.n25 VSUBS 0.291068f
C721 VTAIL.n26 VSUBS 0.031955f
C722 VTAIL.n27 VSUBS 0.030741f
C723 VTAIL.n28 VSUBS 0.016519f
C724 VTAIL.n29 VSUBS 0.039045f
C725 VTAIL.n30 VSUBS 0.017491f
C726 VTAIL.n31 VSUBS 0.49589f
C727 VTAIL.n32 VSUBS 0.016519f
C728 VTAIL.t5 VSUBS 0.084543f
C729 VTAIL.n33 VSUBS 0.122977f
C730 VTAIL.n34 VSUBS 0.024736f
C731 VTAIL.n35 VSUBS 0.029284f
C732 VTAIL.n36 VSUBS 0.039045f
C733 VTAIL.n37 VSUBS 0.017491f
C734 VTAIL.n38 VSUBS 0.016519f
C735 VTAIL.n39 VSUBS 0.030741f
C736 VTAIL.n40 VSUBS 0.030741f
C737 VTAIL.n41 VSUBS 0.016519f
C738 VTAIL.n42 VSUBS 0.017491f
C739 VTAIL.n43 VSUBS 0.039045f
C740 VTAIL.n44 VSUBS 0.088315f
C741 VTAIL.n45 VSUBS 0.017491f
C742 VTAIL.n46 VSUBS 0.016519f
C743 VTAIL.n47 VSUBS 0.068957f
C744 VTAIL.n48 VSUBS 0.044072f
C745 VTAIL.n49 VSUBS 0.291068f
C746 VTAIL.t7 VSUBS 0.10956f
C747 VTAIL.t12 VSUBS 0.10956f
C748 VTAIL.n50 VSUBS 0.578914f
C749 VTAIL.n51 VSUBS 0.938918f
C750 VTAIL.n52 VSUBS 0.031955f
C751 VTAIL.n53 VSUBS 0.030741f
C752 VTAIL.n54 VSUBS 0.016519f
C753 VTAIL.n55 VSUBS 0.039045f
C754 VTAIL.n56 VSUBS 0.017491f
C755 VTAIL.n57 VSUBS 0.49589f
C756 VTAIL.n58 VSUBS 0.016519f
C757 VTAIL.t6 VSUBS 0.084543f
C758 VTAIL.n59 VSUBS 0.122977f
C759 VTAIL.n60 VSUBS 0.024736f
C760 VTAIL.n61 VSUBS 0.029284f
C761 VTAIL.n62 VSUBS 0.039045f
C762 VTAIL.n63 VSUBS 0.017491f
C763 VTAIL.n64 VSUBS 0.016519f
C764 VTAIL.n65 VSUBS 0.030741f
C765 VTAIL.n66 VSUBS 0.030741f
C766 VTAIL.n67 VSUBS 0.016519f
C767 VTAIL.n68 VSUBS 0.017491f
C768 VTAIL.n69 VSUBS 0.039045f
C769 VTAIL.n70 VSUBS 0.088315f
C770 VTAIL.n71 VSUBS 0.017491f
C771 VTAIL.n72 VSUBS 0.016519f
C772 VTAIL.n73 VSUBS 0.068957f
C773 VTAIL.n74 VSUBS 0.044072f
C774 VTAIL.n75 VSUBS 1.26669f
C775 VTAIL.n76 VSUBS 0.031955f
C776 VTAIL.n77 VSUBS 0.030741f
C777 VTAIL.n78 VSUBS 0.016519f
C778 VTAIL.n79 VSUBS 0.039045f
C779 VTAIL.n80 VSUBS 0.017491f
C780 VTAIL.n81 VSUBS 0.49589f
C781 VTAIL.n82 VSUBS 0.016519f
C782 VTAIL.t15 VSUBS 0.084543f
C783 VTAIL.n83 VSUBS 0.122977f
C784 VTAIL.n84 VSUBS 0.024736f
C785 VTAIL.n85 VSUBS 0.029284f
C786 VTAIL.n86 VSUBS 0.039045f
C787 VTAIL.n87 VSUBS 0.017491f
C788 VTAIL.n88 VSUBS 0.016519f
C789 VTAIL.n89 VSUBS 0.030741f
C790 VTAIL.n90 VSUBS 0.030741f
C791 VTAIL.n91 VSUBS 0.016519f
C792 VTAIL.n92 VSUBS 0.017491f
C793 VTAIL.n93 VSUBS 0.039045f
C794 VTAIL.n94 VSUBS 0.088315f
C795 VTAIL.n95 VSUBS 0.017491f
C796 VTAIL.n96 VSUBS 0.016519f
C797 VTAIL.n97 VSUBS 0.068957f
C798 VTAIL.n98 VSUBS 0.044072f
C799 VTAIL.n99 VSUBS 1.26669f
C800 VTAIL.t3 VSUBS 0.10956f
C801 VTAIL.t13 VSUBS 0.10956f
C802 VTAIL.n100 VSUBS 0.578918f
C803 VTAIL.n101 VSUBS 0.938914f
C804 VTAIL.n102 VSUBS 0.031955f
C805 VTAIL.n103 VSUBS 0.030741f
C806 VTAIL.n104 VSUBS 0.016519f
C807 VTAIL.n105 VSUBS 0.039045f
C808 VTAIL.n106 VSUBS 0.017491f
C809 VTAIL.n107 VSUBS 0.49589f
C810 VTAIL.n108 VSUBS 0.016519f
C811 VTAIL.t1 VSUBS 0.084543f
C812 VTAIL.n109 VSUBS 0.122977f
C813 VTAIL.n110 VSUBS 0.024736f
C814 VTAIL.n111 VSUBS 0.029284f
C815 VTAIL.n112 VSUBS 0.039045f
C816 VTAIL.n113 VSUBS 0.017491f
C817 VTAIL.n114 VSUBS 0.016519f
C818 VTAIL.n115 VSUBS 0.030741f
C819 VTAIL.n116 VSUBS 0.030741f
C820 VTAIL.n117 VSUBS 0.016519f
C821 VTAIL.n118 VSUBS 0.017491f
C822 VTAIL.n119 VSUBS 0.039045f
C823 VTAIL.n120 VSUBS 0.088315f
C824 VTAIL.n121 VSUBS 0.017491f
C825 VTAIL.n122 VSUBS 0.016519f
C826 VTAIL.n123 VSUBS 0.068957f
C827 VTAIL.n124 VSUBS 0.044072f
C828 VTAIL.n125 VSUBS 0.291068f
C829 VTAIL.n126 VSUBS 0.031955f
C830 VTAIL.n127 VSUBS 0.030741f
C831 VTAIL.n128 VSUBS 0.016519f
C832 VTAIL.n129 VSUBS 0.039045f
C833 VTAIL.n130 VSUBS 0.017491f
C834 VTAIL.n131 VSUBS 0.49589f
C835 VTAIL.n132 VSUBS 0.016519f
C836 VTAIL.t10 VSUBS 0.084543f
C837 VTAIL.n133 VSUBS 0.122977f
C838 VTAIL.n134 VSUBS 0.024736f
C839 VTAIL.n135 VSUBS 0.029284f
C840 VTAIL.n136 VSUBS 0.039045f
C841 VTAIL.n137 VSUBS 0.017491f
C842 VTAIL.n138 VSUBS 0.016519f
C843 VTAIL.n139 VSUBS 0.030741f
C844 VTAIL.n140 VSUBS 0.030741f
C845 VTAIL.n141 VSUBS 0.016519f
C846 VTAIL.n142 VSUBS 0.017491f
C847 VTAIL.n143 VSUBS 0.039045f
C848 VTAIL.n144 VSUBS 0.088315f
C849 VTAIL.n145 VSUBS 0.017491f
C850 VTAIL.n146 VSUBS 0.016519f
C851 VTAIL.n147 VSUBS 0.068957f
C852 VTAIL.n148 VSUBS 0.044072f
C853 VTAIL.n149 VSUBS 0.291068f
C854 VTAIL.t8 VSUBS 0.10956f
C855 VTAIL.t9 VSUBS 0.10956f
C856 VTAIL.n150 VSUBS 0.578918f
C857 VTAIL.n151 VSUBS 0.938914f
C858 VTAIL.n152 VSUBS 0.031955f
C859 VTAIL.n153 VSUBS 0.030741f
C860 VTAIL.n154 VSUBS 0.016519f
C861 VTAIL.n155 VSUBS 0.039045f
C862 VTAIL.n156 VSUBS 0.017491f
C863 VTAIL.n157 VSUBS 0.49589f
C864 VTAIL.n158 VSUBS 0.016519f
C865 VTAIL.t11 VSUBS 0.084543f
C866 VTAIL.n159 VSUBS 0.122977f
C867 VTAIL.n160 VSUBS 0.024736f
C868 VTAIL.n161 VSUBS 0.029284f
C869 VTAIL.n162 VSUBS 0.039045f
C870 VTAIL.n163 VSUBS 0.017491f
C871 VTAIL.n164 VSUBS 0.016519f
C872 VTAIL.n165 VSUBS 0.030741f
C873 VTAIL.n166 VSUBS 0.030741f
C874 VTAIL.n167 VSUBS 0.016519f
C875 VTAIL.n168 VSUBS 0.017491f
C876 VTAIL.n169 VSUBS 0.039045f
C877 VTAIL.n170 VSUBS 0.088315f
C878 VTAIL.n171 VSUBS 0.017491f
C879 VTAIL.n172 VSUBS 0.016519f
C880 VTAIL.n173 VSUBS 0.068957f
C881 VTAIL.n174 VSUBS 0.044072f
C882 VTAIL.n175 VSUBS 1.26669f
C883 VTAIL.n176 VSUBS 0.031955f
C884 VTAIL.n177 VSUBS 0.030741f
C885 VTAIL.n178 VSUBS 0.016519f
C886 VTAIL.n179 VSUBS 0.039045f
C887 VTAIL.n180 VSUBS 0.017491f
C888 VTAIL.n181 VSUBS 0.49589f
C889 VTAIL.n182 VSUBS 0.016519f
C890 VTAIL.t2 VSUBS 0.084543f
C891 VTAIL.n183 VSUBS 0.122977f
C892 VTAIL.n184 VSUBS 0.024736f
C893 VTAIL.n185 VSUBS 0.029284f
C894 VTAIL.n186 VSUBS 0.039045f
C895 VTAIL.n187 VSUBS 0.017491f
C896 VTAIL.n188 VSUBS 0.016519f
C897 VTAIL.n189 VSUBS 0.030741f
C898 VTAIL.n190 VSUBS 0.030741f
C899 VTAIL.n191 VSUBS 0.016519f
C900 VTAIL.n192 VSUBS 0.017491f
C901 VTAIL.n193 VSUBS 0.039045f
C902 VTAIL.n194 VSUBS 0.088315f
C903 VTAIL.n195 VSUBS 0.017491f
C904 VTAIL.n196 VSUBS 0.016519f
C905 VTAIL.n197 VSUBS 0.068957f
C906 VTAIL.n198 VSUBS 0.044072f
C907 VTAIL.n199 VSUBS 1.26093f
C908 VDD1.t7 VSUBS 0.088567f
C909 VDD1.t1 VSUBS 0.088567f
C910 VDD1.n0 VSUBS 0.545322f
C911 VDD1.t6 VSUBS 0.088567f
C912 VDD1.t2 VSUBS 0.088567f
C913 VDD1.n1 VSUBS 0.544534f
C914 VDD1.t3 VSUBS 0.088567f
C915 VDD1.t4 VSUBS 0.088567f
C916 VDD1.n2 VSUBS 0.544534f
C917 VDD1.n3 VSUBS 2.97777f
C918 VDD1.t5 VSUBS 0.088567f
C919 VDD1.t0 VSUBS 0.088567f
C920 VDD1.n4 VSUBS 0.538066f
C921 VDD1.n5 VSUBS 2.42242f
C922 VP.n0 VSUBS 0.058352f
C923 VP.t7 VSUBS 1.16045f
C924 VP.n1 VSUBS 0.038646f
C925 VP.n2 VSUBS 0.04426f
C926 VP.t0 VSUBS 1.16045f
C927 VP.n3 VSUBS 0.087966f
C928 VP.n4 VSUBS 0.04426f
C929 VP.t5 VSUBS 1.16045f
C930 VP.n5 VSUBS 0.458409f
C931 VP.n6 VSUBS 0.04426f
C932 VP.n7 VSUBS 0.083665f
C933 VP.n8 VSUBS 0.058352f
C934 VP.t1 VSUBS 1.16045f
C935 VP.n9 VSUBS 0.038646f
C936 VP.n10 VSUBS 0.04426f
C937 VP.t3 VSUBS 1.16045f
C938 VP.n11 VSUBS 0.087966f
C939 VP.n12 VSUBS 0.04426f
C940 VP.t4 VSUBS 1.16045f
C941 VP.n13 VSUBS 0.576429f
C942 VP.t2 VSUBS 1.44778f
C943 VP.n14 VSUBS 0.555262f
C944 VP.n15 VSUBS 0.378532f
C945 VP.n16 VSUBS 0.064975f
C946 VP.n17 VSUBS 0.087966f
C947 VP.n18 VSUBS 0.03578f
C948 VP.n19 VSUBS 0.04426f
C949 VP.n20 VSUBS 0.04426f
C950 VP.n21 VSUBS 0.04426f
C951 VP.n22 VSUBS 0.064975f
C952 VP.n23 VSUBS 0.458409f
C953 VP.n24 VSUBS 0.059273f
C954 VP.n25 VSUBS 0.0894f
C955 VP.n26 VSUBS 0.04426f
C956 VP.n27 VSUBS 0.04426f
C957 VP.n28 VSUBS 0.04426f
C958 VP.n29 VSUBS 0.083665f
C959 VP.n30 VSUBS 0.070676f
C960 VP.n31 VSUBS 0.6035f
C961 VP.n32 VSUBS 1.98474f
C962 VP.n33 VSUBS 2.02125f
C963 VP.t6 VSUBS 1.16045f
C964 VP.n34 VSUBS 0.6035f
C965 VP.n35 VSUBS 0.070676f
C966 VP.n36 VSUBS 0.058352f
C967 VP.n37 VSUBS 0.04426f
C968 VP.n38 VSUBS 0.04426f
C969 VP.n39 VSUBS 0.038646f
C970 VP.n40 VSUBS 0.0894f
C971 VP.n41 VSUBS 0.059273f
C972 VP.n42 VSUBS 0.04426f
C973 VP.n43 VSUBS 0.04426f
C974 VP.n44 VSUBS 0.064975f
C975 VP.n45 VSUBS 0.087966f
C976 VP.n46 VSUBS 0.03578f
C977 VP.n47 VSUBS 0.04426f
C978 VP.n48 VSUBS 0.04426f
C979 VP.n49 VSUBS 0.04426f
C980 VP.n50 VSUBS 0.064975f
C981 VP.n51 VSUBS 0.458409f
C982 VP.n52 VSUBS 0.059273f
C983 VP.n53 VSUBS 0.0894f
C984 VP.n54 VSUBS 0.04426f
C985 VP.n55 VSUBS 0.04426f
C986 VP.n56 VSUBS 0.04426f
C987 VP.n57 VSUBS 0.083665f
C988 VP.n58 VSUBS 0.070676f
C989 VP.n59 VSUBS 0.6035f
C990 VP.n60 VSUBS 0.058811f
.ends

