* NGSPICE file created from diff_pair_sample_0096.ext - technology: sky130A

.subckt diff_pair_sample_0096 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t15 VN.t0 VDD2.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=1.9305 pd=12.03 as=1.9305 ps=12.03 w=11.7 l=0.19
X1 VTAIL.t14 VN.t1 VDD2.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=1.9305 pd=12.03 as=1.9305 ps=12.03 w=11.7 l=0.19
X2 VTAIL.t2 VP.t0 VDD1.t7 B.t2 sky130_fd_pr__nfet_01v8 ad=4.563 pd=24.18 as=1.9305 ps=12.03 w=11.7 l=0.19
X3 B.t21 B.t19 B.t20 B.t9 sky130_fd_pr__nfet_01v8 ad=4.563 pd=24.18 as=0 ps=0 w=11.7 l=0.19
X4 VDD1.t6 VP.t1 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=1.9305 pd=12.03 as=4.563 ps=24.18 w=11.7 l=0.19
X5 VDD2.t2 VN.t2 VTAIL.t13 B.t5 sky130_fd_pr__nfet_01v8 ad=1.9305 pd=12.03 as=1.9305 ps=12.03 w=11.7 l=0.19
X6 VDD2.t7 VN.t3 VTAIL.t12 B.t0 sky130_fd_pr__nfet_01v8 ad=1.9305 pd=12.03 as=1.9305 ps=12.03 w=11.7 l=0.19
X7 VTAIL.t4 VP.t2 VDD1.t5 B.t4 sky130_fd_pr__nfet_01v8 ad=1.9305 pd=12.03 as=1.9305 ps=12.03 w=11.7 l=0.19
X8 B.t18 B.t16 B.t17 B.t13 sky130_fd_pr__nfet_01v8 ad=4.563 pd=24.18 as=0 ps=0 w=11.7 l=0.19
X9 VDD2.t0 VN.t4 VTAIL.t11 B.t1 sky130_fd_pr__nfet_01v8 ad=1.9305 pd=12.03 as=4.563 ps=24.18 w=11.7 l=0.19
X10 B.t15 B.t12 B.t14 B.t13 sky130_fd_pr__nfet_01v8 ad=4.563 pd=24.18 as=0 ps=0 w=11.7 l=0.19
X11 VDD1.t4 VP.t3 VTAIL.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=1.9305 pd=12.03 as=1.9305 ps=12.03 w=11.7 l=0.19
X12 VTAIL.t6 VP.t4 VDD1.t3 B.t6 sky130_fd_pr__nfet_01v8 ad=4.563 pd=24.18 as=1.9305 ps=12.03 w=11.7 l=0.19
X13 VDD2.t1 VN.t5 VTAIL.t10 B.t7 sky130_fd_pr__nfet_01v8 ad=1.9305 pd=12.03 as=4.563 ps=24.18 w=11.7 l=0.19
X14 VDD1.t2 VP.t5 VTAIL.t7 B.t7 sky130_fd_pr__nfet_01v8 ad=1.9305 pd=12.03 as=4.563 ps=24.18 w=11.7 l=0.19
X15 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=4.563 pd=24.18 as=0 ps=0 w=11.7 l=0.19
X16 VTAIL.t9 VN.t6 VDD2.t5 B.t6 sky130_fd_pr__nfet_01v8 ad=4.563 pd=24.18 as=1.9305 ps=12.03 w=11.7 l=0.19
X17 VTAIL.t8 VN.t7 VDD2.t6 B.t2 sky130_fd_pr__nfet_01v8 ad=4.563 pd=24.18 as=1.9305 ps=12.03 w=11.7 l=0.19
X18 VDD1.t1 VP.t6 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=1.9305 pd=12.03 as=1.9305 ps=12.03 w=11.7 l=0.19
X19 VTAIL.t3 VP.t7 VDD1.t0 B.t3 sky130_fd_pr__nfet_01v8 ad=1.9305 pd=12.03 as=1.9305 ps=12.03 w=11.7 l=0.19
R0 VN.n5 VN.t4 1689.84
R1 VN.n1 VN.t7 1689.84
R2 VN.n12 VN.t6 1689.84
R3 VN.n8 VN.t5 1689.84
R4 VN.n4 VN.t1 1648.95
R5 VN.n2 VN.t2 1648.95
R6 VN.n11 VN.t3 1648.95
R7 VN.n9 VN.t0 1648.95
R8 VN.n8 VN.n7 161.489
R9 VN.n1 VN.n0 161.489
R10 VN.n6 VN.n5 161.3
R11 VN.n13 VN.n12 161.3
R12 VN.n10 VN.n7 161.3
R13 VN.n3 VN.n0 161.3
R14 VN VN.n13 39.813
R15 VN.n3 VN.n2 37.9763
R16 VN.n4 VN.n3 37.9763
R17 VN.n11 VN.n10 37.9763
R18 VN.n10 VN.n9 37.9763
R19 VN.n2 VN.n1 35.055
R20 VN.n5 VN.n4 35.055
R21 VN.n12 VN.n11 35.055
R22 VN.n9 VN.n8 35.055
R23 VN.n13 VN.n7 0.189894
R24 VN.n6 VN.n0 0.189894
R25 VN VN.n6 0.0516364
R26 VDD2.n2 VDD2.n1 60.985
R27 VDD2.n2 VDD2.n0 60.985
R28 VDD2 VDD2.n5 60.9822
R29 VDD2.n4 VDD2.n3 60.8164
R30 VDD2.n4 VDD2.n2 35.8187
R31 VDD2.n5 VDD2.t4 1.69281
R32 VDD2.n5 VDD2.t1 1.69281
R33 VDD2.n3 VDD2.t5 1.69281
R34 VDD2.n3 VDD2.t7 1.69281
R35 VDD2.n1 VDD2.t3 1.69281
R36 VDD2.n1 VDD2.t0 1.69281
R37 VDD2.n0 VDD2.t6 1.69281
R38 VDD2.n0 VDD2.t2 1.69281
R39 VDD2 VDD2.n4 0.282828
R40 VTAIL.n11 VTAIL.t2 45.8299
R41 VTAIL.n10 VTAIL.t10 45.8299
R42 VTAIL.n7 VTAIL.t9 45.8299
R43 VTAIL.n15 VTAIL.t11 45.8297
R44 VTAIL.n2 VTAIL.t8 45.8297
R45 VTAIL.n3 VTAIL.t7 45.8297
R46 VTAIL.n6 VTAIL.t6 45.8297
R47 VTAIL.n14 VTAIL.t1 45.8297
R48 VTAIL.n13 VTAIL.n12 44.1376
R49 VTAIL.n9 VTAIL.n8 44.1376
R50 VTAIL.n1 VTAIL.n0 44.1374
R51 VTAIL.n5 VTAIL.n4 44.1374
R52 VTAIL.n15 VTAIL.n14 22.9014
R53 VTAIL.n7 VTAIL.n6 22.9014
R54 VTAIL.n0 VTAIL.t13 1.69281
R55 VTAIL.n0 VTAIL.t14 1.69281
R56 VTAIL.n4 VTAIL.t0 1.69281
R57 VTAIL.n4 VTAIL.t4 1.69281
R58 VTAIL.n12 VTAIL.t5 1.69281
R59 VTAIL.n12 VTAIL.t3 1.69281
R60 VTAIL.n8 VTAIL.t12 1.69281
R61 VTAIL.n8 VTAIL.t15 1.69281
R62 VTAIL.n11 VTAIL.n10 0.470328
R63 VTAIL.n3 VTAIL.n2 0.470328
R64 VTAIL.n9 VTAIL.n7 0.448776
R65 VTAIL.n10 VTAIL.n9 0.448776
R66 VTAIL.n13 VTAIL.n11 0.448776
R67 VTAIL.n14 VTAIL.n13 0.448776
R68 VTAIL.n6 VTAIL.n5 0.448776
R69 VTAIL.n5 VTAIL.n3 0.448776
R70 VTAIL.n2 VTAIL.n1 0.448776
R71 VTAIL VTAIL.n15 0.390586
R72 VTAIL VTAIL.n1 0.0586897
R73 B.n83 B.t12 1723.57
R74 B.n80 B.t16 1723.57
R75 B.n342 B.t19 1723.57
R76 B.n339 B.t8 1723.57
R77 B.n592 B.n591 585
R78 B.n593 B.n592 585
R79 B.n264 B.n79 585
R80 B.n263 B.n262 585
R81 B.n261 B.n260 585
R82 B.n259 B.n258 585
R83 B.n257 B.n256 585
R84 B.n255 B.n254 585
R85 B.n253 B.n252 585
R86 B.n251 B.n250 585
R87 B.n249 B.n248 585
R88 B.n247 B.n246 585
R89 B.n245 B.n244 585
R90 B.n243 B.n242 585
R91 B.n241 B.n240 585
R92 B.n239 B.n238 585
R93 B.n237 B.n236 585
R94 B.n235 B.n234 585
R95 B.n233 B.n232 585
R96 B.n231 B.n230 585
R97 B.n229 B.n228 585
R98 B.n227 B.n226 585
R99 B.n225 B.n224 585
R100 B.n223 B.n222 585
R101 B.n221 B.n220 585
R102 B.n219 B.n218 585
R103 B.n217 B.n216 585
R104 B.n215 B.n214 585
R105 B.n213 B.n212 585
R106 B.n211 B.n210 585
R107 B.n209 B.n208 585
R108 B.n207 B.n206 585
R109 B.n205 B.n204 585
R110 B.n203 B.n202 585
R111 B.n201 B.n200 585
R112 B.n199 B.n198 585
R113 B.n197 B.n196 585
R114 B.n195 B.n194 585
R115 B.n193 B.n192 585
R116 B.n191 B.n190 585
R117 B.n189 B.n188 585
R118 B.n187 B.n186 585
R119 B.n185 B.n184 585
R120 B.n183 B.n182 585
R121 B.n181 B.n180 585
R122 B.n179 B.n178 585
R123 B.n177 B.n176 585
R124 B.n175 B.n174 585
R125 B.n173 B.n172 585
R126 B.n171 B.n170 585
R127 B.n169 B.n168 585
R128 B.n166 B.n165 585
R129 B.n164 B.n163 585
R130 B.n162 B.n161 585
R131 B.n160 B.n159 585
R132 B.n158 B.n157 585
R133 B.n156 B.n155 585
R134 B.n154 B.n153 585
R135 B.n152 B.n151 585
R136 B.n150 B.n149 585
R137 B.n148 B.n147 585
R138 B.n146 B.n145 585
R139 B.n144 B.n143 585
R140 B.n142 B.n141 585
R141 B.n140 B.n139 585
R142 B.n138 B.n137 585
R143 B.n136 B.n135 585
R144 B.n134 B.n133 585
R145 B.n132 B.n131 585
R146 B.n130 B.n129 585
R147 B.n128 B.n127 585
R148 B.n126 B.n125 585
R149 B.n124 B.n123 585
R150 B.n122 B.n121 585
R151 B.n120 B.n119 585
R152 B.n118 B.n117 585
R153 B.n116 B.n115 585
R154 B.n114 B.n113 585
R155 B.n112 B.n111 585
R156 B.n110 B.n109 585
R157 B.n108 B.n107 585
R158 B.n106 B.n105 585
R159 B.n104 B.n103 585
R160 B.n102 B.n101 585
R161 B.n100 B.n99 585
R162 B.n98 B.n97 585
R163 B.n96 B.n95 585
R164 B.n94 B.n93 585
R165 B.n92 B.n91 585
R166 B.n90 B.n89 585
R167 B.n88 B.n87 585
R168 B.n86 B.n85 585
R169 B.n590 B.n33 585
R170 B.n594 B.n33 585
R171 B.n589 B.n32 585
R172 B.n595 B.n32 585
R173 B.n588 B.n587 585
R174 B.n587 B.n28 585
R175 B.n586 B.n27 585
R176 B.n601 B.n27 585
R177 B.n585 B.n26 585
R178 B.n602 B.n26 585
R179 B.n584 B.n25 585
R180 B.n603 B.n25 585
R181 B.n583 B.n582 585
R182 B.n582 B.n21 585
R183 B.n581 B.n20 585
R184 B.n609 B.n20 585
R185 B.n580 B.n19 585
R186 B.n610 B.n19 585
R187 B.n579 B.n18 585
R188 B.n611 B.n18 585
R189 B.n578 B.n577 585
R190 B.n577 B.n17 585
R191 B.n576 B.n12 585
R192 B.n617 B.n12 585
R193 B.n575 B.n11 585
R194 B.n618 B.n11 585
R195 B.n574 B.n10 585
R196 B.n619 B.n10 585
R197 B.n573 B.n7 585
R198 B.n622 B.n7 585
R199 B.n572 B.n6 585
R200 B.n623 B.n6 585
R201 B.n571 B.n5 585
R202 B.n624 B.n5 585
R203 B.n570 B.n569 585
R204 B.n569 B.n4 585
R205 B.n568 B.n265 585
R206 B.n568 B.n567 585
R207 B.n558 B.n266 585
R208 B.n267 B.n266 585
R209 B.n560 B.n559 585
R210 B.n561 B.n560 585
R211 B.n557 B.n271 585
R212 B.n274 B.n271 585
R213 B.n556 B.n555 585
R214 B.n555 B.n554 585
R215 B.n273 B.n272 585
R216 B.n547 B.n273 585
R217 B.n546 B.n545 585
R218 B.n548 B.n546 585
R219 B.n544 B.n279 585
R220 B.n279 B.n278 585
R221 B.n543 B.n542 585
R222 B.n542 B.n541 585
R223 B.n281 B.n280 585
R224 B.n282 B.n281 585
R225 B.n534 B.n533 585
R226 B.n535 B.n534 585
R227 B.n532 B.n287 585
R228 B.n287 B.n286 585
R229 B.n531 B.n530 585
R230 B.n530 B.n529 585
R231 B.n289 B.n288 585
R232 B.n290 B.n289 585
R233 B.n525 B.n524 585
R234 B.n293 B.n292 585
R235 B.n521 B.n520 585
R236 B.n522 B.n521 585
R237 B.n519 B.n338 585
R238 B.n518 B.n517 585
R239 B.n516 B.n515 585
R240 B.n514 B.n513 585
R241 B.n512 B.n511 585
R242 B.n510 B.n509 585
R243 B.n508 B.n507 585
R244 B.n506 B.n505 585
R245 B.n504 B.n503 585
R246 B.n502 B.n501 585
R247 B.n500 B.n499 585
R248 B.n498 B.n497 585
R249 B.n496 B.n495 585
R250 B.n494 B.n493 585
R251 B.n492 B.n491 585
R252 B.n490 B.n489 585
R253 B.n488 B.n487 585
R254 B.n486 B.n485 585
R255 B.n484 B.n483 585
R256 B.n482 B.n481 585
R257 B.n480 B.n479 585
R258 B.n478 B.n477 585
R259 B.n476 B.n475 585
R260 B.n474 B.n473 585
R261 B.n472 B.n471 585
R262 B.n470 B.n469 585
R263 B.n468 B.n467 585
R264 B.n466 B.n465 585
R265 B.n464 B.n463 585
R266 B.n462 B.n461 585
R267 B.n460 B.n459 585
R268 B.n458 B.n457 585
R269 B.n456 B.n455 585
R270 B.n454 B.n453 585
R271 B.n452 B.n451 585
R272 B.n450 B.n449 585
R273 B.n448 B.n447 585
R274 B.n446 B.n445 585
R275 B.n444 B.n443 585
R276 B.n442 B.n441 585
R277 B.n440 B.n439 585
R278 B.n438 B.n437 585
R279 B.n436 B.n435 585
R280 B.n434 B.n433 585
R281 B.n432 B.n431 585
R282 B.n430 B.n429 585
R283 B.n428 B.n427 585
R284 B.n425 B.n424 585
R285 B.n423 B.n422 585
R286 B.n421 B.n420 585
R287 B.n419 B.n418 585
R288 B.n417 B.n416 585
R289 B.n415 B.n414 585
R290 B.n413 B.n412 585
R291 B.n411 B.n410 585
R292 B.n409 B.n408 585
R293 B.n407 B.n406 585
R294 B.n405 B.n404 585
R295 B.n403 B.n402 585
R296 B.n401 B.n400 585
R297 B.n399 B.n398 585
R298 B.n397 B.n396 585
R299 B.n395 B.n394 585
R300 B.n393 B.n392 585
R301 B.n391 B.n390 585
R302 B.n389 B.n388 585
R303 B.n387 B.n386 585
R304 B.n385 B.n384 585
R305 B.n383 B.n382 585
R306 B.n381 B.n380 585
R307 B.n379 B.n378 585
R308 B.n377 B.n376 585
R309 B.n375 B.n374 585
R310 B.n373 B.n372 585
R311 B.n371 B.n370 585
R312 B.n369 B.n368 585
R313 B.n367 B.n366 585
R314 B.n365 B.n364 585
R315 B.n363 B.n362 585
R316 B.n361 B.n360 585
R317 B.n359 B.n358 585
R318 B.n357 B.n356 585
R319 B.n355 B.n354 585
R320 B.n353 B.n352 585
R321 B.n351 B.n350 585
R322 B.n349 B.n348 585
R323 B.n347 B.n346 585
R324 B.n345 B.n344 585
R325 B.n526 B.n291 585
R326 B.n291 B.n290 585
R327 B.n528 B.n527 585
R328 B.n529 B.n528 585
R329 B.n285 B.n284 585
R330 B.n286 B.n285 585
R331 B.n537 B.n536 585
R332 B.n536 B.n535 585
R333 B.n538 B.n283 585
R334 B.n283 B.n282 585
R335 B.n540 B.n539 585
R336 B.n541 B.n540 585
R337 B.n277 B.n276 585
R338 B.n278 B.n277 585
R339 B.n550 B.n549 585
R340 B.n549 B.n548 585
R341 B.n551 B.n275 585
R342 B.n547 B.n275 585
R343 B.n553 B.n552 585
R344 B.n554 B.n553 585
R345 B.n270 B.n269 585
R346 B.n274 B.n270 585
R347 B.n563 B.n562 585
R348 B.n562 B.n561 585
R349 B.n564 B.n268 585
R350 B.n268 B.n267 585
R351 B.n566 B.n565 585
R352 B.n567 B.n566 585
R353 B.n3 B.n0 585
R354 B.n4 B.n3 585
R355 B.n621 B.n1 585
R356 B.n622 B.n621 585
R357 B.n620 B.n9 585
R358 B.n620 B.n619 585
R359 B.n14 B.n8 585
R360 B.n618 B.n8 585
R361 B.n616 B.n615 585
R362 B.n617 B.n616 585
R363 B.n614 B.n13 585
R364 B.n17 B.n13 585
R365 B.n613 B.n612 585
R366 B.n612 B.n611 585
R367 B.n16 B.n15 585
R368 B.n610 B.n16 585
R369 B.n608 B.n607 585
R370 B.n609 B.n608 585
R371 B.n606 B.n22 585
R372 B.n22 B.n21 585
R373 B.n605 B.n604 585
R374 B.n604 B.n603 585
R375 B.n24 B.n23 585
R376 B.n602 B.n24 585
R377 B.n600 B.n599 585
R378 B.n601 B.n600 585
R379 B.n598 B.n29 585
R380 B.n29 B.n28 585
R381 B.n597 B.n596 585
R382 B.n596 B.n595 585
R383 B.n31 B.n30 585
R384 B.n594 B.n31 585
R385 B.n625 B.n624 585
R386 B.n623 B.n2 585
R387 B.n85 B.n31 545.355
R388 B.n592 B.n33 545.355
R389 B.n344 B.n289 545.355
R390 B.n524 B.n291 545.355
R391 B.n593 B.n78 256.663
R392 B.n593 B.n77 256.663
R393 B.n593 B.n76 256.663
R394 B.n593 B.n75 256.663
R395 B.n593 B.n74 256.663
R396 B.n593 B.n73 256.663
R397 B.n593 B.n72 256.663
R398 B.n593 B.n71 256.663
R399 B.n593 B.n70 256.663
R400 B.n593 B.n69 256.663
R401 B.n593 B.n68 256.663
R402 B.n593 B.n67 256.663
R403 B.n593 B.n66 256.663
R404 B.n593 B.n65 256.663
R405 B.n593 B.n64 256.663
R406 B.n593 B.n63 256.663
R407 B.n593 B.n62 256.663
R408 B.n593 B.n61 256.663
R409 B.n593 B.n60 256.663
R410 B.n593 B.n59 256.663
R411 B.n593 B.n58 256.663
R412 B.n593 B.n57 256.663
R413 B.n593 B.n56 256.663
R414 B.n593 B.n55 256.663
R415 B.n593 B.n54 256.663
R416 B.n593 B.n53 256.663
R417 B.n593 B.n52 256.663
R418 B.n593 B.n51 256.663
R419 B.n593 B.n50 256.663
R420 B.n593 B.n49 256.663
R421 B.n593 B.n48 256.663
R422 B.n593 B.n47 256.663
R423 B.n593 B.n46 256.663
R424 B.n593 B.n45 256.663
R425 B.n593 B.n44 256.663
R426 B.n593 B.n43 256.663
R427 B.n593 B.n42 256.663
R428 B.n593 B.n41 256.663
R429 B.n593 B.n40 256.663
R430 B.n593 B.n39 256.663
R431 B.n593 B.n38 256.663
R432 B.n593 B.n37 256.663
R433 B.n593 B.n36 256.663
R434 B.n593 B.n35 256.663
R435 B.n593 B.n34 256.663
R436 B.n523 B.n522 256.663
R437 B.n522 B.n294 256.663
R438 B.n522 B.n295 256.663
R439 B.n522 B.n296 256.663
R440 B.n522 B.n297 256.663
R441 B.n522 B.n298 256.663
R442 B.n522 B.n299 256.663
R443 B.n522 B.n300 256.663
R444 B.n522 B.n301 256.663
R445 B.n522 B.n302 256.663
R446 B.n522 B.n303 256.663
R447 B.n522 B.n304 256.663
R448 B.n522 B.n305 256.663
R449 B.n522 B.n306 256.663
R450 B.n522 B.n307 256.663
R451 B.n522 B.n308 256.663
R452 B.n522 B.n309 256.663
R453 B.n522 B.n310 256.663
R454 B.n522 B.n311 256.663
R455 B.n522 B.n312 256.663
R456 B.n522 B.n313 256.663
R457 B.n522 B.n314 256.663
R458 B.n522 B.n315 256.663
R459 B.n522 B.n316 256.663
R460 B.n522 B.n317 256.663
R461 B.n522 B.n318 256.663
R462 B.n522 B.n319 256.663
R463 B.n522 B.n320 256.663
R464 B.n522 B.n321 256.663
R465 B.n522 B.n322 256.663
R466 B.n522 B.n323 256.663
R467 B.n522 B.n324 256.663
R468 B.n522 B.n325 256.663
R469 B.n522 B.n326 256.663
R470 B.n522 B.n327 256.663
R471 B.n522 B.n328 256.663
R472 B.n522 B.n329 256.663
R473 B.n522 B.n330 256.663
R474 B.n522 B.n331 256.663
R475 B.n522 B.n332 256.663
R476 B.n522 B.n333 256.663
R477 B.n522 B.n334 256.663
R478 B.n522 B.n335 256.663
R479 B.n522 B.n336 256.663
R480 B.n522 B.n337 256.663
R481 B.n627 B.n626 256.663
R482 B.n89 B.n88 163.367
R483 B.n93 B.n92 163.367
R484 B.n97 B.n96 163.367
R485 B.n101 B.n100 163.367
R486 B.n105 B.n104 163.367
R487 B.n109 B.n108 163.367
R488 B.n113 B.n112 163.367
R489 B.n117 B.n116 163.367
R490 B.n121 B.n120 163.367
R491 B.n125 B.n124 163.367
R492 B.n129 B.n128 163.367
R493 B.n133 B.n132 163.367
R494 B.n137 B.n136 163.367
R495 B.n141 B.n140 163.367
R496 B.n145 B.n144 163.367
R497 B.n149 B.n148 163.367
R498 B.n153 B.n152 163.367
R499 B.n157 B.n156 163.367
R500 B.n161 B.n160 163.367
R501 B.n165 B.n164 163.367
R502 B.n170 B.n169 163.367
R503 B.n174 B.n173 163.367
R504 B.n178 B.n177 163.367
R505 B.n182 B.n181 163.367
R506 B.n186 B.n185 163.367
R507 B.n190 B.n189 163.367
R508 B.n194 B.n193 163.367
R509 B.n198 B.n197 163.367
R510 B.n202 B.n201 163.367
R511 B.n206 B.n205 163.367
R512 B.n210 B.n209 163.367
R513 B.n214 B.n213 163.367
R514 B.n218 B.n217 163.367
R515 B.n222 B.n221 163.367
R516 B.n226 B.n225 163.367
R517 B.n230 B.n229 163.367
R518 B.n234 B.n233 163.367
R519 B.n238 B.n237 163.367
R520 B.n242 B.n241 163.367
R521 B.n246 B.n245 163.367
R522 B.n250 B.n249 163.367
R523 B.n254 B.n253 163.367
R524 B.n258 B.n257 163.367
R525 B.n262 B.n261 163.367
R526 B.n592 B.n79 163.367
R527 B.n530 B.n289 163.367
R528 B.n530 B.n287 163.367
R529 B.n534 B.n287 163.367
R530 B.n534 B.n281 163.367
R531 B.n542 B.n281 163.367
R532 B.n542 B.n279 163.367
R533 B.n546 B.n279 163.367
R534 B.n546 B.n273 163.367
R535 B.n555 B.n273 163.367
R536 B.n555 B.n271 163.367
R537 B.n560 B.n271 163.367
R538 B.n560 B.n266 163.367
R539 B.n568 B.n266 163.367
R540 B.n569 B.n568 163.367
R541 B.n569 B.n5 163.367
R542 B.n6 B.n5 163.367
R543 B.n7 B.n6 163.367
R544 B.n10 B.n7 163.367
R545 B.n11 B.n10 163.367
R546 B.n12 B.n11 163.367
R547 B.n577 B.n12 163.367
R548 B.n577 B.n18 163.367
R549 B.n19 B.n18 163.367
R550 B.n20 B.n19 163.367
R551 B.n582 B.n20 163.367
R552 B.n582 B.n25 163.367
R553 B.n26 B.n25 163.367
R554 B.n27 B.n26 163.367
R555 B.n587 B.n27 163.367
R556 B.n587 B.n32 163.367
R557 B.n33 B.n32 163.367
R558 B.n521 B.n293 163.367
R559 B.n521 B.n338 163.367
R560 B.n517 B.n516 163.367
R561 B.n513 B.n512 163.367
R562 B.n509 B.n508 163.367
R563 B.n505 B.n504 163.367
R564 B.n501 B.n500 163.367
R565 B.n497 B.n496 163.367
R566 B.n493 B.n492 163.367
R567 B.n489 B.n488 163.367
R568 B.n485 B.n484 163.367
R569 B.n481 B.n480 163.367
R570 B.n477 B.n476 163.367
R571 B.n473 B.n472 163.367
R572 B.n469 B.n468 163.367
R573 B.n465 B.n464 163.367
R574 B.n461 B.n460 163.367
R575 B.n457 B.n456 163.367
R576 B.n453 B.n452 163.367
R577 B.n449 B.n448 163.367
R578 B.n445 B.n444 163.367
R579 B.n441 B.n440 163.367
R580 B.n437 B.n436 163.367
R581 B.n433 B.n432 163.367
R582 B.n429 B.n428 163.367
R583 B.n424 B.n423 163.367
R584 B.n420 B.n419 163.367
R585 B.n416 B.n415 163.367
R586 B.n412 B.n411 163.367
R587 B.n408 B.n407 163.367
R588 B.n404 B.n403 163.367
R589 B.n400 B.n399 163.367
R590 B.n396 B.n395 163.367
R591 B.n392 B.n391 163.367
R592 B.n388 B.n387 163.367
R593 B.n384 B.n383 163.367
R594 B.n380 B.n379 163.367
R595 B.n376 B.n375 163.367
R596 B.n372 B.n371 163.367
R597 B.n368 B.n367 163.367
R598 B.n364 B.n363 163.367
R599 B.n360 B.n359 163.367
R600 B.n356 B.n355 163.367
R601 B.n352 B.n351 163.367
R602 B.n348 B.n347 163.367
R603 B.n528 B.n291 163.367
R604 B.n528 B.n285 163.367
R605 B.n536 B.n285 163.367
R606 B.n536 B.n283 163.367
R607 B.n540 B.n283 163.367
R608 B.n540 B.n277 163.367
R609 B.n549 B.n277 163.367
R610 B.n549 B.n275 163.367
R611 B.n553 B.n275 163.367
R612 B.n553 B.n270 163.367
R613 B.n562 B.n270 163.367
R614 B.n562 B.n268 163.367
R615 B.n566 B.n268 163.367
R616 B.n566 B.n3 163.367
R617 B.n625 B.n3 163.367
R618 B.n621 B.n2 163.367
R619 B.n621 B.n620 163.367
R620 B.n620 B.n8 163.367
R621 B.n616 B.n8 163.367
R622 B.n616 B.n13 163.367
R623 B.n612 B.n13 163.367
R624 B.n612 B.n16 163.367
R625 B.n608 B.n16 163.367
R626 B.n608 B.n22 163.367
R627 B.n604 B.n22 163.367
R628 B.n604 B.n24 163.367
R629 B.n600 B.n24 163.367
R630 B.n600 B.n29 163.367
R631 B.n596 B.n29 163.367
R632 B.n596 B.n31 163.367
R633 B.n522 B.n290 91.3702
R634 B.n594 B.n593 91.3702
R635 B.n80 B.t17 80.6317
R636 B.n342 B.t21 80.6317
R637 B.n83 B.t14 80.617
R638 B.n339 B.t11 80.617
R639 B.n85 B.n34 71.676
R640 B.n89 B.n35 71.676
R641 B.n93 B.n36 71.676
R642 B.n97 B.n37 71.676
R643 B.n101 B.n38 71.676
R644 B.n105 B.n39 71.676
R645 B.n109 B.n40 71.676
R646 B.n113 B.n41 71.676
R647 B.n117 B.n42 71.676
R648 B.n121 B.n43 71.676
R649 B.n125 B.n44 71.676
R650 B.n129 B.n45 71.676
R651 B.n133 B.n46 71.676
R652 B.n137 B.n47 71.676
R653 B.n141 B.n48 71.676
R654 B.n145 B.n49 71.676
R655 B.n149 B.n50 71.676
R656 B.n153 B.n51 71.676
R657 B.n157 B.n52 71.676
R658 B.n161 B.n53 71.676
R659 B.n165 B.n54 71.676
R660 B.n170 B.n55 71.676
R661 B.n174 B.n56 71.676
R662 B.n178 B.n57 71.676
R663 B.n182 B.n58 71.676
R664 B.n186 B.n59 71.676
R665 B.n190 B.n60 71.676
R666 B.n194 B.n61 71.676
R667 B.n198 B.n62 71.676
R668 B.n202 B.n63 71.676
R669 B.n206 B.n64 71.676
R670 B.n210 B.n65 71.676
R671 B.n214 B.n66 71.676
R672 B.n218 B.n67 71.676
R673 B.n222 B.n68 71.676
R674 B.n226 B.n69 71.676
R675 B.n230 B.n70 71.676
R676 B.n234 B.n71 71.676
R677 B.n238 B.n72 71.676
R678 B.n242 B.n73 71.676
R679 B.n246 B.n74 71.676
R680 B.n250 B.n75 71.676
R681 B.n254 B.n76 71.676
R682 B.n258 B.n77 71.676
R683 B.n262 B.n78 71.676
R684 B.n79 B.n78 71.676
R685 B.n261 B.n77 71.676
R686 B.n257 B.n76 71.676
R687 B.n253 B.n75 71.676
R688 B.n249 B.n74 71.676
R689 B.n245 B.n73 71.676
R690 B.n241 B.n72 71.676
R691 B.n237 B.n71 71.676
R692 B.n233 B.n70 71.676
R693 B.n229 B.n69 71.676
R694 B.n225 B.n68 71.676
R695 B.n221 B.n67 71.676
R696 B.n217 B.n66 71.676
R697 B.n213 B.n65 71.676
R698 B.n209 B.n64 71.676
R699 B.n205 B.n63 71.676
R700 B.n201 B.n62 71.676
R701 B.n197 B.n61 71.676
R702 B.n193 B.n60 71.676
R703 B.n189 B.n59 71.676
R704 B.n185 B.n58 71.676
R705 B.n181 B.n57 71.676
R706 B.n177 B.n56 71.676
R707 B.n173 B.n55 71.676
R708 B.n169 B.n54 71.676
R709 B.n164 B.n53 71.676
R710 B.n160 B.n52 71.676
R711 B.n156 B.n51 71.676
R712 B.n152 B.n50 71.676
R713 B.n148 B.n49 71.676
R714 B.n144 B.n48 71.676
R715 B.n140 B.n47 71.676
R716 B.n136 B.n46 71.676
R717 B.n132 B.n45 71.676
R718 B.n128 B.n44 71.676
R719 B.n124 B.n43 71.676
R720 B.n120 B.n42 71.676
R721 B.n116 B.n41 71.676
R722 B.n112 B.n40 71.676
R723 B.n108 B.n39 71.676
R724 B.n104 B.n38 71.676
R725 B.n100 B.n37 71.676
R726 B.n96 B.n36 71.676
R727 B.n92 B.n35 71.676
R728 B.n88 B.n34 71.676
R729 B.n524 B.n523 71.676
R730 B.n338 B.n294 71.676
R731 B.n516 B.n295 71.676
R732 B.n512 B.n296 71.676
R733 B.n508 B.n297 71.676
R734 B.n504 B.n298 71.676
R735 B.n500 B.n299 71.676
R736 B.n496 B.n300 71.676
R737 B.n492 B.n301 71.676
R738 B.n488 B.n302 71.676
R739 B.n484 B.n303 71.676
R740 B.n480 B.n304 71.676
R741 B.n476 B.n305 71.676
R742 B.n472 B.n306 71.676
R743 B.n468 B.n307 71.676
R744 B.n464 B.n308 71.676
R745 B.n460 B.n309 71.676
R746 B.n456 B.n310 71.676
R747 B.n452 B.n311 71.676
R748 B.n448 B.n312 71.676
R749 B.n444 B.n313 71.676
R750 B.n440 B.n314 71.676
R751 B.n436 B.n315 71.676
R752 B.n432 B.n316 71.676
R753 B.n428 B.n317 71.676
R754 B.n423 B.n318 71.676
R755 B.n419 B.n319 71.676
R756 B.n415 B.n320 71.676
R757 B.n411 B.n321 71.676
R758 B.n407 B.n322 71.676
R759 B.n403 B.n323 71.676
R760 B.n399 B.n324 71.676
R761 B.n395 B.n325 71.676
R762 B.n391 B.n326 71.676
R763 B.n387 B.n327 71.676
R764 B.n383 B.n328 71.676
R765 B.n379 B.n329 71.676
R766 B.n375 B.n330 71.676
R767 B.n371 B.n331 71.676
R768 B.n367 B.n332 71.676
R769 B.n363 B.n333 71.676
R770 B.n359 B.n334 71.676
R771 B.n355 B.n335 71.676
R772 B.n351 B.n336 71.676
R773 B.n347 B.n337 71.676
R774 B.n523 B.n293 71.676
R775 B.n517 B.n294 71.676
R776 B.n513 B.n295 71.676
R777 B.n509 B.n296 71.676
R778 B.n505 B.n297 71.676
R779 B.n501 B.n298 71.676
R780 B.n497 B.n299 71.676
R781 B.n493 B.n300 71.676
R782 B.n489 B.n301 71.676
R783 B.n485 B.n302 71.676
R784 B.n481 B.n303 71.676
R785 B.n477 B.n304 71.676
R786 B.n473 B.n305 71.676
R787 B.n469 B.n306 71.676
R788 B.n465 B.n307 71.676
R789 B.n461 B.n308 71.676
R790 B.n457 B.n309 71.676
R791 B.n453 B.n310 71.676
R792 B.n449 B.n311 71.676
R793 B.n445 B.n312 71.676
R794 B.n441 B.n313 71.676
R795 B.n437 B.n314 71.676
R796 B.n433 B.n315 71.676
R797 B.n429 B.n316 71.676
R798 B.n424 B.n317 71.676
R799 B.n420 B.n318 71.676
R800 B.n416 B.n319 71.676
R801 B.n412 B.n320 71.676
R802 B.n408 B.n321 71.676
R803 B.n404 B.n322 71.676
R804 B.n400 B.n323 71.676
R805 B.n396 B.n324 71.676
R806 B.n392 B.n325 71.676
R807 B.n388 B.n326 71.676
R808 B.n384 B.n327 71.676
R809 B.n380 B.n328 71.676
R810 B.n376 B.n329 71.676
R811 B.n372 B.n330 71.676
R812 B.n368 B.n331 71.676
R813 B.n364 B.n332 71.676
R814 B.n360 B.n333 71.676
R815 B.n356 B.n334 71.676
R816 B.n352 B.n335 71.676
R817 B.n348 B.n336 71.676
R818 B.n344 B.n337 71.676
R819 B.n626 B.n625 71.676
R820 B.n626 B.n2 71.676
R821 B.n81 B.t18 70.5468
R822 B.n343 B.t20 70.5468
R823 B.n84 B.t15 70.5321
R824 B.n340 B.t10 70.5321
R825 B.n167 B.n84 59.5399
R826 B.n82 B.n81 59.5399
R827 B.n426 B.n343 59.5399
R828 B.n341 B.n340 59.5399
R829 B.n529 B.n290 44.0653
R830 B.n529 B.n286 44.0653
R831 B.n535 B.n286 44.0653
R832 B.n541 B.n282 44.0653
R833 B.n541 B.n278 44.0653
R834 B.n548 B.n278 44.0653
R835 B.n548 B.n547 44.0653
R836 B.n554 B.n274 44.0653
R837 B.n567 B.n267 44.0653
R838 B.n624 B.n4 44.0653
R839 B.n624 B.n623 44.0653
R840 B.n623 B.n622 44.0653
R841 B.n619 B.n618 44.0653
R842 B.n611 B.n17 44.0653
R843 B.n610 B.n609 44.0653
R844 B.n609 B.n21 44.0653
R845 B.n603 B.n21 44.0653
R846 B.n603 B.n602 44.0653
R847 B.n601 B.n28 44.0653
R848 B.n595 B.n28 44.0653
R849 B.n595 B.n594 44.0653
R850 B.n561 B.t0 40.8252
R851 B.n617 B.t3 40.8252
R852 B.t7 B.n4 38.2332
R853 B.n622 B.t2 38.2332
R854 B.n535 B.t9 35.6411
R855 B.t13 B.n601 35.6411
R856 B.n526 B.n525 35.4346
R857 B.n345 B.n288 35.4346
R858 B.n591 B.n590 35.4346
R859 B.n86 B.n30 35.4346
R860 B.n561 B.t4 26.569
R861 B.t5 B.n617 26.569
R862 B.n547 B.t6 23.9769
R863 B.t1 B.n610 23.9769
R864 B.n554 B.t6 20.0889
R865 B.n611 B.t1 20.0889
R866 B B.n627 18.0485
R867 B.t4 B.n267 17.4968
R868 B.n618 B.t5 17.4968
R869 B.n527 B.n526 10.6151
R870 B.n527 B.n284 10.6151
R871 B.n537 B.n284 10.6151
R872 B.n538 B.n537 10.6151
R873 B.n539 B.n538 10.6151
R874 B.n539 B.n276 10.6151
R875 B.n550 B.n276 10.6151
R876 B.n551 B.n550 10.6151
R877 B.n552 B.n551 10.6151
R878 B.n552 B.n269 10.6151
R879 B.n563 B.n269 10.6151
R880 B.n564 B.n563 10.6151
R881 B.n565 B.n564 10.6151
R882 B.n565 B.n0 10.6151
R883 B.n525 B.n292 10.6151
R884 B.n520 B.n292 10.6151
R885 B.n520 B.n519 10.6151
R886 B.n519 B.n518 10.6151
R887 B.n518 B.n515 10.6151
R888 B.n515 B.n514 10.6151
R889 B.n514 B.n511 10.6151
R890 B.n511 B.n510 10.6151
R891 B.n510 B.n507 10.6151
R892 B.n507 B.n506 10.6151
R893 B.n506 B.n503 10.6151
R894 B.n503 B.n502 10.6151
R895 B.n502 B.n499 10.6151
R896 B.n499 B.n498 10.6151
R897 B.n498 B.n495 10.6151
R898 B.n495 B.n494 10.6151
R899 B.n494 B.n491 10.6151
R900 B.n491 B.n490 10.6151
R901 B.n490 B.n487 10.6151
R902 B.n487 B.n486 10.6151
R903 B.n486 B.n483 10.6151
R904 B.n483 B.n482 10.6151
R905 B.n482 B.n479 10.6151
R906 B.n479 B.n478 10.6151
R907 B.n478 B.n475 10.6151
R908 B.n475 B.n474 10.6151
R909 B.n474 B.n471 10.6151
R910 B.n471 B.n470 10.6151
R911 B.n470 B.n467 10.6151
R912 B.n467 B.n466 10.6151
R913 B.n466 B.n463 10.6151
R914 B.n463 B.n462 10.6151
R915 B.n462 B.n459 10.6151
R916 B.n459 B.n458 10.6151
R917 B.n458 B.n455 10.6151
R918 B.n455 B.n454 10.6151
R919 B.n454 B.n451 10.6151
R920 B.n451 B.n450 10.6151
R921 B.n450 B.n447 10.6151
R922 B.n447 B.n446 10.6151
R923 B.n443 B.n442 10.6151
R924 B.n442 B.n439 10.6151
R925 B.n439 B.n438 10.6151
R926 B.n438 B.n435 10.6151
R927 B.n435 B.n434 10.6151
R928 B.n434 B.n431 10.6151
R929 B.n431 B.n430 10.6151
R930 B.n430 B.n427 10.6151
R931 B.n425 B.n422 10.6151
R932 B.n422 B.n421 10.6151
R933 B.n421 B.n418 10.6151
R934 B.n418 B.n417 10.6151
R935 B.n417 B.n414 10.6151
R936 B.n414 B.n413 10.6151
R937 B.n413 B.n410 10.6151
R938 B.n410 B.n409 10.6151
R939 B.n409 B.n406 10.6151
R940 B.n406 B.n405 10.6151
R941 B.n405 B.n402 10.6151
R942 B.n402 B.n401 10.6151
R943 B.n401 B.n398 10.6151
R944 B.n398 B.n397 10.6151
R945 B.n397 B.n394 10.6151
R946 B.n394 B.n393 10.6151
R947 B.n393 B.n390 10.6151
R948 B.n390 B.n389 10.6151
R949 B.n389 B.n386 10.6151
R950 B.n386 B.n385 10.6151
R951 B.n385 B.n382 10.6151
R952 B.n382 B.n381 10.6151
R953 B.n381 B.n378 10.6151
R954 B.n378 B.n377 10.6151
R955 B.n377 B.n374 10.6151
R956 B.n374 B.n373 10.6151
R957 B.n373 B.n370 10.6151
R958 B.n370 B.n369 10.6151
R959 B.n369 B.n366 10.6151
R960 B.n366 B.n365 10.6151
R961 B.n365 B.n362 10.6151
R962 B.n362 B.n361 10.6151
R963 B.n361 B.n358 10.6151
R964 B.n358 B.n357 10.6151
R965 B.n357 B.n354 10.6151
R966 B.n354 B.n353 10.6151
R967 B.n353 B.n350 10.6151
R968 B.n350 B.n349 10.6151
R969 B.n349 B.n346 10.6151
R970 B.n346 B.n345 10.6151
R971 B.n531 B.n288 10.6151
R972 B.n532 B.n531 10.6151
R973 B.n533 B.n532 10.6151
R974 B.n533 B.n280 10.6151
R975 B.n543 B.n280 10.6151
R976 B.n544 B.n543 10.6151
R977 B.n545 B.n544 10.6151
R978 B.n545 B.n272 10.6151
R979 B.n556 B.n272 10.6151
R980 B.n557 B.n556 10.6151
R981 B.n559 B.n557 10.6151
R982 B.n559 B.n558 10.6151
R983 B.n558 B.n265 10.6151
R984 B.n570 B.n265 10.6151
R985 B.n571 B.n570 10.6151
R986 B.n572 B.n571 10.6151
R987 B.n573 B.n572 10.6151
R988 B.n574 B.n573 10.6151
R989 B.n575 B.n574 10.6151
R990 B.n576 B.n575 10.6151
R991 B.n578 B.n576 10.6151
R992 B.n579 B.n578 10.6151
R993 B.n580 B.n579 10.6151
R994 B.n581 B.n580 10.6151
R995 B.n583 B.n581 10.6151
R996 B.n584 B.n583 10.6151
R997 B.n585 B.n584 10.6151
R998 B.n586 B.n585 10.6151
R999 B.n588 B.n586 10.6151
R1000 B.n589 B.n588 10.6151
R1001 B.n590 B.n589 10.6151
R1002 B.n9 B.n1 10.6151
R1003 B.n14 B.n9 10.6151
R1004 B.n615 B.n14 10.6151
R1005 B.n615 B.n614 10.6151
R1006 B.n614 B.n613 10.6151
R1007 B.n613 B.n15 10.6151
R1008 B.n607 B.n15 10.6151
R1009 B.n607 B.n606 10.6151
R1010 B.n606 B.n605 10.6151
R1011 B.n605 B.n23 10.6151
R1012 B.n599 B.n23 10.6151
R1013 B.n599 B.n598 10.6151
R1014 B.n598 B.n597 10.6151
R1015 B.n597 B.n30 10.6151
R1016 B.n87 B.n86 10.6151
R1017 B.n90 B.n87 10.6151
R1018 B.n91 B.n90 10.6151
R1019 B.n94 B.n91 10.6151
R1020 B.n95 B.n94 10.6151
R1021 B.n98 B.n95 10.6151
R1022 B.n99 B.n98 10.6151
R1023 B.n102 B.n99 10.6151
R1024 B.n103 B.n102 10.6151
R1025 B.n106 B.n103 10.6151
R1026 B.n107 B.n106 10.6151
R1027 B.n110 B.n107 10.6151
R1028 B.n111 B.n110 10.6151
R1029 B.n114 B.n111 10.6151
R1030 B.n115 B.n114 10.6151
R1031 B.n118 B.n115 10.6151
R1032 B.n119 B.n118 10.6151
R1033 B.n122 B.n119 10.6151
R1034 B.n123 B.n122 10.6151
R1035 B.n126 B.n123 10.6151
R1036 B.n127 B.n126 10.6151
R1037 B.n130 B.n127 10.6151
R1038 B.n131 B.n130 10.6151
R1039 B.n134 B.n131 10.6151
R1040 B.n135 B.n134 10.6151
R1041 B.n138 B.n135 10.6151
R1042 B.n139 B.n138 10.6151
R1043 B.n142 B.n139 10.6151
R1044 B.n143 B.n142 10.6151
R1045 B.n146 B.n143 10.6151
R1046 B.n147 B.n146 10.6151
R1047 B.n150 B.n147 10.6151
R1048 B.n151 B.n150 10.6151
R1049 B.n154 B.n151 10.6151
R1050 B.n155 B.n154 10.6151
R1051 B.n158 B.n155 10.6151
R1052 B.n159 B.n158 10.6151
R1053 B.n162 B.n159 10.6151
R1054 B.n163 B.n162 10.6151
R1055 B.n166 B.n163 10.6151
R1056 B.n171 B.n168 10.6151
R1057 B.n172 B.n171 10.6151
R1058 B.n175 B.n172 10.6151
R1059 B.n176 B.n175 10.6151
R1060 B.n179 B.n176 10.6151
R1061 B.n180 B.n179 10.6151
R1062 B.n183 B.n180 10.6151
R1063 B.n184 B.n183 10.6151
R1064 B.n188 B.n187 10.6151
R1065 B.n191 B.n188 10.6151
R1066 B.n192 B.n191 10.6151
R1067 B.n195 B.n192 10.6151
R1068 B.n196 B.n195 10.6151
R1069 B.n199 B.n196 10.6151
R1070 B.n200 B.n199 10.6151
R1071 B.n203 B.n200 10.6151
R1072 B.n204 B.n203 10.6151
R1073 B.n207 B.n204 10.6151
R1074 B.n208 B.n207 10.6151
R1075 B.n211 B.n208 10.6151
R1076 B.n212 B.n211 10.6151
R1077 B.n215 B.n212 10.6151
R1078 B.n216 B.n215 10.6151
R1079 B.n219 B.n216 10.6151
R1080 B.n220 B.n219 10.6151
R1081 B.n223 B.n220 10.6151
R1082 B.n224 B.n223 10.6151
R1083 B.n227 B.n224 10.6151
R1084 B.n228 B.n227 10.6151
R1085 B.n231 B.n228 10.6151
R1086 B.n232 B.n231 10.6151
R1087 B.n235 B.n232 10.6151
R1088 B.n236 B.n235 10.6151
R1089 B.n239 B.n236 10.6151
R1090 B.n240 B.n239 10.6151
R1091 B.n243 B.n240 10.6151
R1092 B.n244 B.n243 10.6151
R1093 B.n247 B.n244 10.6151
R1094 B.n248 B.n247 10.6151
R1095 B.n251 B.n248 10.6151
R1096 B.n252 B.n251 10.6151
R1097 B.n255 B.n252 10.6151
R1098 B.n256 B.n255 10.6151
R1099 B.n259 B.n256 10.6151
R1100 B.n260 B.n259 10.6151
R1101 B.n263 B.n260 10.6151
R1102 B.n264 B.n263 10.6151
R1103 B.n591 B.n264 10.6151
R1104 B.n84 B.n83 10.0853
R1105 B.n81 B.n80 10.0853
R1106 B.n343 B.n342 10.0853
R1107 B.n340 B.n339 10.0853
R1108 B.t9 B.n282 8.42465
R1109 B.n602 B.t13 8.42465
R1110 B.n627 B.n0 8.11757
R1111 B.n627 B.n1 8.11757
R1112 B.n443 B.n341 6.5566
R1113 B.n427 B.n426 6.5566
R1114 B.n168 B.n167 6.5566
R1115 B.n184 B.n82 6.5566
R1116 B.n567 B.t7 5.83261
R1117 B.n619 B.t2 5.83261
R1118 B.n446 B.n341 4.05904
R1119 B.n426 B.n425 4.05904
R1120 B.n167 B.n166 4.05904
R1121 B.n187 B.n82 4.05904
R1122 B.n274 B.t0 3.24056
R1123 B.n17 B.t3 3.24056
R1124 VP.n13 VP.t5 1689.84
R1125 VP.n9 VP.t4 1689.84
R1126 VP.n2 VP.t0 1689.84
R1127 VP.n6 VP.t1 1689.84
R1128 VP.n12 VP.t2 1648.95
R1129 VP.n10 VP.t6 1648.95
R1130 VP.n3 VP.t3 1648.95
R1131 VP.n5 VP.t7 1648.95
R1132 VP.n2 VP.n1 161.489
R1133 VP.n14 VP.n13 161.3
R1134 VP.n4 VP.n1 161.3
R1135 VP.n7 VP.n6 161.3
R1136 VP.n11 VP.n0 161.3
R1137 VP.n9 VP.n8 161.3
R1138 VP.n8 VP.n7 39.4323
R1139 VP.n11 VP.n10 37.9763
R1140 VP.n12 VP.n11 37.9763
R1141 VP.n4 VP.n3 37.9763
R1142 VP.n5 VP.n4 37.9763
R1143 VP.n10 VP.n9 35.055
R1144 VP.n13 VP.n12 35.055
R1145 VP.n3 VP.n2 35.055
R1146 VP.n6 VP.n5 35.055
R1147 VP.n7 VP.n1 0.189894
R1148 VP.n8 VP.n0 0.189894
R1149 VP.n14 VP.n0 0.189894
R1150 VP VP.n14 0.0516364
R1151 VDD1 VDD1.n0 61.0987
R1152 VDD1.n3 VDD1.n2 60.985
R1153 VDD1.n3 VDD1.n1 60.985
R1154 VDD1.n5 VDD1.n4 60.8162
R1155 VDD1.n5 VDD1.n3 36.4018
R1156 VDD1.n4 VDD1.t0 1.69281
R1157 VDD1.n4 VDD1.t6 1.69281
R1158 VDD1.n0 VDD1.t7 1.69281
R1159 VDD1.n0 VDD1.t4 1.69281
R1160 VDD1.n2 VDD1.t5 1.69281
R1161 VDD1.n2 VDD1.t2 1.69281
R1162 VDD1.n1 VDD1.t3 1.69281
R1163 VDD1.n1 VDD1.t1 1.69281
R1164 VDD1 VDD1.n5 0.166448
C0 VDD2 VN 2.47725f
C1 VP VTAIL 2.00177f
C2 VDD1 VTAIL 19.4498f
C3 VDD2 VTAIL 19.488f
C4 VN VTAIL 1.98767f
C5 VP VDD1 2.59292f
C6 VDD2 VP 0.263052f
C7 VN VP 4.65873f
C8 VDD2 VDD1 0.577749f
C9 VN VDD1 0.147201f
C10 VDD2 B 3.052441f
C11 VDD1 B 3.218363f
C12 VTAIL B 8.159462f
C13 VN B 6.47092f
C14 VP B 4.618447f
C15 VDD1.t7 B 0.352691f
C16 VDD1.t4 B 0.352691f
C17 VDD1.n0 B 3.13763f
C18 VDD1.t3 B 0.352691f
C19 VDD1.t1 B 0.352691f
C20 VDD1.n1 B 3.13682f
C21 VDD1.t5 B 0.352691f
C22 VDD1.t2 B 0.352691f
C23 VDD1.n2 B 3.13682f
C24 VDD1.n3 B 2.9195f
C25 VDD1.t0 B 0.352691f
C26 VDD1.t6 B 0.352691f
C27 VDD1.n4 B 3.13567f
C28 VDD1.n5 B 3.23642f
C29 VP.n0 B 0.060968f
C30 VP.t2 B 0.383068f
C31 VP.t6 B 0.383068f
C32 VP.t4 B 0.3869f
C33 VP.n1 B 0.13125f
C34 VP.t7 B 0.383068f
C35 VP.t3 B 0.383068f
C36 VP.t0 B 0.3869f
C37 VP.n2 B 0.175569f
C38 VP.n3 B 0.159469f
C39 VP.n4 B 0.020977f
C40 VP.n5 B 0.159469f
C41 VP.t1 B 0.3869f
C42 VP.n6 B 0.175486f
C43 VP.n7 B 2.25997f
C44 VP.n8 B 2.31571f
C45 VP.n9 B 0.175486f
C46 VP.n10 B 0.159469f
C47 VP.n11 B 0.020977f
C48 VP.n12 B 0.159469f
C49 VP.t5 B 0.3869f
C50 VP.n13 B 0.175486f
C51 VP.n14 B 0.047248f
C52 VTAIL.t13 B 0.241647f
C53 VTAIL.t14 B 0.241647f
C54 VTAIL.n0 B 2.06814f
C55 VTAIL.n1 B 0.304793f
C56 VTAIL.t8 B 2.6354f
C57 VTAIL.n2 B 0.431242f
C58 VTAIL.t7 B 2.6354f
C59 VTAIL.n3 B 0.431242f
C60 VTAIL.t0 B 0.241647f
C61 VTAIL.t4 B 0.241647f
C62 VTAIL.n4 B 2.06814f
C63 VTAIL.n5 B 0.337645f
C64 VTAIL.t6 B 2.6354f
C65 VTAIL.n6 B 1.63388f
C66 VTAIL.t9 B 2.63541f
C67 VTAIL.n7 B 1.63387f
C68 VTAIL.t12 B 0.241647f
C69 VTAIL.t15 B 0.241647f
C70 VTAIL.n8 B 2.06815f
C71 VTAIL.n9 B 0.337638f
C72 VTAIL.t10 B 2.63541f
C73 VTAIL.n10 B 0.431235f
C74 VTAIL.t2 B 2.63541f
C75 VTAIL.n11 B 0.431235f
C76 VTAIL.t5 B 0.241647f
C77 VTAIL.t3 B 0.241647f
C78 VTAIL.n12 B 2.06815f
C79 VTAIL.n13 B 0.337638f
C80 VTAIL.t1 B 2.6354f
C81 VTAIL.n14 B 1.63388f
C82 VTAIL.t11 B 2.6354f
C83 VTAIL.n15 B 1.62898f
C84 VDD2.t6 B 0.354964f
C85 VDD2.t2 B 0.354964f
C86 VDD2.n0 B 3.15704f
C87 VDD2.t3 B 0.354964f
C88 VDD2.t0 B 0.354964f
C89 VDD2.n1 B 3.15704f
C90 VDD2.n2 B 2.8557f
C91 VDD2.t5 B 0.354964f
C92 VDD2.t7 B 0.354964f
C93 VDD2.n3 B 3.15589f
C94 VDD2.n4 B 3.21248f
C95 VDD2.t4 B 0.354964f
C96 VDD2.t1 B 0.354964f
C97 VDD2.n5 B 3.157f
C98 VN.n0 B 0.100685f
C99 VN.t1 B 0.293861f
C100 VN.t2 B 0.293861f
C101 VN.t7 B 0.296801f
C102 VN.n1 B 0.134683f
C103 VN.n2 B 0.122333f
C104 VN.n3 B 0.016092f
C105 VN.n4 B 0.122333f
C106 VN.t4 B 0.296801f
C107 VN.n5 B 0.13462f
C108 VN.n6 B 0.036245f
C109 VN.n7 B 0.100685f
C110 VN.t6 B 0.296801f
C111 VN.t3 B 0.293861f
C112 VN.t0 B 0.293861f
C113 VN.t5 B 0.296801f
C114 VN.n8 B 0.134683f
C115 VN.n9 B 0.122333f
C116 VN.n10 B 0.016092f
C117 VN.n11 B 0.122333f
C118 VN.n12 B 0.13462f
C119 VN.n13 B 1.76451f
.ends

