* NGSPICE file created from diff_pair_sample_0004.ext - technology: sky130A

.subckt diff_pair_sample_0004 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t7 VP.t0 VDD1.t0 w_n3334_n4204# sky130_fd_pr__pfet_01v8 ad=6.3102 pd=33.14 as=2.6697 ps=16.51 w=16.18 l=3.61
X1 VDD2.t3 VN.t0 VTAIL.t3 w_n3334_n4204# sky130_fd_pr__pfet_01v8 ad=2.6697 pd=16.51 as=6.3102 ps=33.14 w=16.18 l=3.61
X2 B.t11 B.t9 B.t10 w_n3334_n4204# sky130_fd_pr__pfet_01v8 ad=6.3102 pd=33.14 as=0 ps=0 w=16.18 l=3.61
X3 B.t8 B.t6 B.t7 w_n3334_n4204# sky130_fd_pr__pfet_01v8 ad=6.3102 pd=33.14 as=0 ps=0 w=16.18 l=3.61
X4 B.t5 B.t3 B.t4 w_n3334_n4204# sky130_fd_pr__pfet_01v8 ad=6.3102 pd=33.14 as=0 ps=0 w=16.18 l=3.61
X5 VDD2.t2 VN.t1 VTAIL.t1 w_n3334_n4204# sky130_fd_pr__pfet_01v8 ad=2.6697 pd=16.51 as=6.3102 ps=33.14 w=16.18 l=3.61
X6 VDD1.t2 VP.t1 VTAIL.t6 w_n3334_n4204# sky130_fd_pr__pfet_01v8 ad=2.6697 pd=16.51 as=6.3102 ps=33.14 w=16.18 l=3.61
X7 VDD1.t1 VP.t2 VTAIL.t5 w_n3334_n4204# sky130_fd_pr__pfet_01v8 ad=2.6697 pd=16.51 as=6.3102 ps=33.14 w=16.18 l=3.61
X8 VTAIL.t4 VP.t3 VDD1.t3 w_n3334_n4204# sky130_fd_pr__pfet_01v8 ad=6.3102 pd=33.14 as=2.6697 ps=16.51 w=16.18 l=3.61
X9 B.t2 B.t0 B.t1 w_n3334_n4204# sky130_fd_pr__pfet_01v8 ad=6.3102 pd=33.14 as=0 ps=0 w=16.18 l=3.61
X10 VTAIL.t2 VN.t2 VDD2.t1 w_n3334_n4204# sky130_fd_pr__pfet_01v8 ad=6.3102 pd=33.14 as=2.6697 ps=16.51 w=16.18 l=3.61
X11 VTAIL.t0 VN.t3 VDD2.t0 w_n3334_n4204# sky130_fd_pr__pfet_01v8 ad=6.3102 pd=33.14 as=2.6697 ps=16.51 w=16.18 l=3.61
R0 VP.n19 VP.n18 161.3
R1 VP.n17 VP.n1 161.3
R2 VP.n16 VP.n15 161.3
R3 VP.n14 VP.n2 161.3
R4 VP.n13 VP.n12 161.3
R5 VP.n11 VP.n3 161.3
R6 VP.n10 VP.n9 161.3
R7 VP.n8 VP.n4 161.3
R8 VP.n5 VP.t0 143.006
R9 VP.n5 VP.t2 141.76
R10 VP.n6 VP.t3 108.016
R11 VP.n0 VP.t1 108.016
R12 VP.n7 VP.n6 79.4252
R13 VP.n20 VP.n0 79.4252
R14 VP.n12 VP.n2 56.5617
R15 VP.n7 VP.n5 54.7607
R16 VP.n10 VP.n4 24.5923
R17 VP.n11 VP.n10 24.5923
R18 VP.n12 VP.n11 24.5923
R19 VP.n16 VP.n2 24.5923
R20 VP.n17 VP.n16 24.5923
R21 VP.n18 VP.n17 24.5923
R22 VP.n6 VP.n4 10.8209
R23 VP.n18 VP.n0 10.8209
R24 VP.n8 VP.n7 0.354861
R25 VP.n20 VP.n19 0.354861
R26 VP VP.n20 0.267071
R27 VP.n9 VP.n8 0.189894
R28 VP.n9 VP.n3 0.189894
R29 VP.n13 VP.n3 0.189894
R30 VP.n14 VP.n13 0.189894
R31 VP.n15 VP.n14 0.189894
R32 VP.n15 VP.n1 0.189894
R33 VP.n19 VP.n1 0.189894
R34 VDD1 VDD1.n1 120.118
R35 VDD1 VDD1.n0 71.7995
R36 VDD1.n0 VDD1.t0 2.00946
R37 VDD1.n0 VDD1.t1 2.00946
R38 VDD1.n1 VDD1.t3 2.00946
R39 VDD1.n1 VDD1.t2 2.00946
R40 VTAIL.n714 VTAIL.n630 756.745
R41 VTAIL.n84 VTAIL.n0 756.745
R42 VTAIL.n174 VTAIL.n90 756.745
R43 VTAIL.n264 VTAIL.n180 756.745
R44 VTAIL.n624 VTAIL.n540 756.745
R45 VTAIL.n534 VTAIL.n450 756.745
R46 VTAIL.n444 VTAIL.n360 756.745
R47 VTAIL.n354 VTAIL.n270 756.745
R48 VTAIL.n658 VTAIL.n657 585
R49 VTAIL.n663 VTAIL.n662 585
R50 VTAIL.n665 VTAIL.n664 585
R51 VTAIL.n654 VTAIL.n653 585
R52 VTAIL.n671 VTAIL.n670 585
R53 VTAIL.n673 VTAIL.n672 585
R54 VTAIL.n650 VTAIL.n649 585
R55 VTAIL.n679 VTAIL.n678 585
R56 VTAIL.n681 VTAIL.n680 585
R57 VTAIL.n646 VTAIL.n645 585
R58 VTAIL.n687 VTAIL.n686 585
R59 VTAIL.n689 VTAIL.n688 585
R60 VTAIL.n642 VTAIL.n641 585
R61 VTAIL.n695 VTAIL.n694 585
R62 VTAIL.n697 VTAIL.n696 585
R63 VTAIL.n638 VTAIL.n637 585
R64 VTAIL.n704 VTAIL.n703 585
R65 VTAIL.n705 VTAIL.n636 585
R66 VTAIL.n707 VTAIL.n706 585
R67 VTAIL.n634 VTAIL.n633 585
R68 VTAIL.n713 VTAIL.n712 585
R69 VTAIL.n715 VTAIL.n714 585
R70 VTAIL.n28 VTAIL.n27 585
R71 VTAIL.n33 VTAIL.n32 585
R72 VTAIL.n35 VTAIL.n34 585
R73 VTAIL.n24 VTAIL.n23 585
R74 VTAIL.n41 VTAIL.n40 585
R75 VTAIL.n43 VTAIL.n42 585
R76 VTAIL.n20 VTAIL.n19 585
R77 VTAIL.n49 VTAIL.n48 585
R78 VTAIL.n51 VTAIL.n50 585
R79 VTAIL.n16 VTAIL.n15 585
R80 VTAIL.n57 VTAIL.n56 585
R81 VTAIL.n59 VTAIL.n58 585
R82 VTAIL.n12 VTAIL.n11 585
R83 VTAIL.n65 VTAIL.n64 585
R84 VTAIL.n67 VTAIL.n66 585
R85 VTAIL.n8 VTAIL.n7 585
R86 VTAIL.n74 VTAIL.n73 585
R87 VTAIL.n75 VTAIL.n6 585
R88 VTAIL.n77 VTAIL.n76 585
R89 VTAIL.n4 VTAIL.n3 585
R90 VTAIL.n83 VTAIL.n82 585
R91 VTAIL.n85 VTAIL.n84 585
R92 VTAIL.n118 VTAIL.n117 585
R93 VTAIL.n123 VTAIL.n122 585
R94 VTAIL.n125 VTAIL.n124 585
R95 VTAIL.n114 VTAIL.n113 585
R96 VTAIL.n131 VTAIL.n130 585
R97 VTAIL.n133 VTAIL.n132 585
R98 VTAIL.n110 VTAIL.n109 585
R99 VTAIL.n139 VTAIL.n138 585
R100 VTAIL.n141 VTAIL.n140 585
R101 VTAIL.n106 VTAIL.n105 585
R102 VTAIL.n147 VTAIL.n146 585
R103 VTAIL.n149 VTAIL.n148 585
R104 VTAIL.n102 VTAIL.n101 585
R105 VTAIL.n155 VTAIL.n154 585
R106 VTAIL.n157 VTAIL.n156 585
R107 VTAIL.n98 VTAIL.n97 585
R108 VTAIL.n164 VTAIL.n163 585
R109 VTAIL.n165 VTAIL.n96 585
R110 VTAIL.n167 VTAIL.n166 585
R111 VTAIL.n94 VTAIL.n93 585
R112 VTAIL.n173 VTAIL.n172 585
R113 VTAIL.n175 VTAIL.n174 585
R114 VTAIL.n208 VTAIL.n207 585
R115 VTAIL.n213 VTAIL.n212 585
R116 VTAIL.n215 VTAIL.n214 585
R117 VTAIL.n204 VTAIL.n203 585
R118 VTAIL.n221 VTAIL.n220 585
R119 VTAIL.n223 VTAIL.n222 585
R120 VTAIL.n200 VTAIL.n199 585
R121 VTAIL.n229 VTAIL.n228 585
R122 VTAIL.n231 VTAIL.n230 585
R123 VTAIL.n196 VTAIL.n195 585
R124 VTAIL.n237 VTAIL.n236 585
R125 VTAIL.n239 VTAIL.n238 585
R126 VTAIL.n192 VTAIL.n191 585
R127 VTAIL.n245 VTAIL.n244 585
R128 VTAIL.n247 VTAIL.n246 585
R129 VTAIL.n188 VTAIL.n187 585
R130 VTAIL.n254 VTAIL.n253 585
R131 VTAIL.n255 VTAIL.n186 585
R132 VTAIL.n257 VTAIL.n256 585
R133 VTAIL.n184 VTAIL.n183 585
R134 VTAIL.n263 VTAIL.n262 585
R135 VTAIL.n265 VTAIL.n264 585
R136 VTAIL.n625 VTAIL.n624 585
R137 VTAIL.n623 VTAIL.n622 585
R138 VTAIL.n544 VTAIL.n543 585
R139 VTAIL.n617 VTAIL.n616 585
R140 VTAIL.n615 VTAIL.n546 585
R141 VTAIL.n614 VTAIL.n613 585
R142 VTAIL.n549 VTAIL.n547 585
R143 VTAIL.n608 VTAIL.n607 585
R144 VTAIL.n606 VTAIL.n605 585
R145 VTAIL.n553 VTAIL.n552 585
R146 VTAIL.n600 VTAIL.n599 585
R147 VTAIL.n598 VTAIL.n597 585
R148 VTAIL.n557 VTAIL.n556 585
R149 VTAIL.n592 VTAIL.n591 585
R150 VTAIL.n590 VTAIL.n589 585
R151 VTAIL.n561 VTAIL.n560 585
R152 VTAIL.n584 VTAIL.n583 585
R153 VTAIL.n582 VTAIL.n581 585
R154 VTAIL.n565 VTAIL.n564 585
R155 VTAIL.n576 VTAIL.n575 585
R156 VTAIL.n574 VTAIL.n573 585
R157 VTAIL.n569 VTAIL.n568 585
R158 VTAIL.n535 VTAIL.n534 585
R159 VTAIL.n533 VTAIL.n532 585
R160 VTAIL.n454 VTAIL.n453 585
R161 VTAIL.n527 VTAIL.n526 585
R162 VTAIL.n525 VTAIL.n456 585
R163 VTAIL.n524 VTAIL.n523 585
R164 VTAIL.n459 VTAIL.n457 585
R165 VTAIL.n518 VTAIL.n517 585
R166 VTAIL.n516 VTAIL.n515 585
R167 VTAIL.n463 VTAIL.n462 585
R168 VTAIL.n510 VTAIL.n509 585
R169 VTAIL.n508 VTAIL.n507 585
R170 VTAIL.n467 VTAIL.n466 585
R171 VTAIL.n502 VTAIL.n501 585
R172 VTAIL.n500 VTAIL.n499 585
R173 VTAIL.n471 VTAIL.n470 585
R174 VTAIL.n494 VTAIL.n493 585
R175 VTAIL.n492 VTAIL.n491 585
R176 VTAIL.n475 VTAIL.n474 585
R177 VTAIL.n486 VTAIL.n485 585
R178 VTAIL.n484 VTAIL.n483 585
R179 VTAIL.n479 VTAIL.n478 585
R180 VTAIL.n445 VTAIL.n444 585
R181 VTAIL.n443 VTAIL.n442 585
R182 VTAIL.n364 VTAIL.n363 585
R183 VTAIL.n437 VTAIL.n436 585
R184 VTAIL.n435 VTAIL.n366 585
R185 VTAIL.n434 VTAIL.n433 585
R186 VTAIL.n369 VTAIL.n367 585
R187 VTAIL.n428 VTAIL.n427 585
R188 VTAIL.n426 VTAIL.n425 585
R189 VTAIL.n373 VTAIL.n372 585
R190 VTAIL.n420 VTAIL.n419 585
R191 VTAIL.n418 VTAIL.n417 585
R192 VTAIL.n377 VTAIL.n376 585
R193 VTAIL.n412 VTAIL.n411 585
R194 VTAIL.n410 VTAIL.n409 585
R195 VTAIL.n381 VTAIL.n380 585
R196 VTAIL.n404 VTAIL.n403 585
R197 VTAIL.n402 VTAIL.n401 585
R198 VTAIL.n385 VTAIL.n384 585
R199 VTAIL.n396 VTAIL.n395 585
R200 VTAIL.n394 VTAIL.n393 585
R201 VTAIL.n389 VTAIL.n388 585
R202 VTAIL.n355 VTAIL.n354 585
R203 VTAIL.n353 VTAIL.n352 585
R204 VTAIL.n274 VTAIL.n273 585
R205 VTAIL.n347 VTAIL.n346 585
R206 VTAIL.n345 VTAIL.n276 585
R207 VTAIL.n344 VTAIL.n343 585
R208 VTAIL.n279 VTAIL.n277 585
R209 VTAIL.n338 VTAIL.n337 585
R210 VTAIL.n336 VTAIL.n335 585
R211 VTAIL.n283 VTAIL.n282 585
R212 VTAIL.n330 VTAIL.n329 585
R213 VTAIL.n328 VTAIL.n327 585
R214 VTAIL.n287 VTAIL.n286 585
R215 VTAIL.n322 VTAIL.n321 585
R216 VTAIL.n320 VTAIL.n319 585
R217 VTAIL.n291 VTAIL.n290 585
R218 VTAIL.n314 VTAIL.n313 585
R219 VTAIL.n312 VTAIL.n311 585
R220 VTAIL.n295 VTAIL.n294 585
R221 VTAIL.n306 VTAIL.n305 585
R222 VTAIL.n304 VTAIL.n303 585
R223 VTAIL.n299 VTAIL.n298 585
R224 VTAIL.n659 VTAIL.t3 327.466
R225 VTAIL.n29 VTAIL.t0 327.466
R226 VTAIL.n119 VTAIL.t6 327.466
R227 VTAIL.n209 VTAIL.t4 327.466
R228 VTAIL.n570 VTAIL.t5 327.466
R229 VTAIL.n480 VTAIL.t7 327.466
R230 VTAIL.n390 VTAIL.t1 327.466
R231 VTAIL.n300 VTAIL.t2 327.466
R232 VTAIL.n663 VTAIL.n657 171.744
R233 VTAIL.n664 VTAIL.n663 171.744
R234 VTAIL.n664 VTAIL.n653 171.744
R235 VTAIL.n671 VTAIL.n653 171.744
R236 VTAIL.n672 VTAIL.n671 171.744
R237 VTAIL.n672 VTAIL.n649 171.744
R238 VTAIL.n679 VTAIL.n649 171.744
R239 VTAIL.n680 VTAIL.n679 171.744
R240 VTAIL.n680 VTAIL.n645 171.744
R241 VTAIL.n687 VTAIL.n645 171.744
R242 VTAIL.n688 VTAIL.n687 171.744
R243 VTAIL.n688 VTAIL.n641 171.744
R244 VTAIL.n695 VTAIL.n641 171.744
R245 VTAIL.n696 VTAIL.n695 171.744
R246 VTAIL.n696 VTAIL.n637 171.744
R247 VTAIL.n704 VTAIL.n637 171.744
R248 VTAIL.n705 VTAIL.n704 171.744
R249 VTAIL.n706 VTAIL.n705 171.744
R250 VTAIL.n706 VTAIL.n633 171.744
R251 VTAIL.n713 VTAIL.n633 171.744
R252 VTAIL.n714 VTAIL.n713 171.744
R253 VTAIL.n33 VTAIL.n27 171.744
R254 VTAIL.n34 VTAIL.n33 171.744
R255 VTAIL.n34 VTAIL.n23 171.744
R256 VTAIL.n41 VTAIL.n23 171.744
R257 VTAIL.n42 VTAIL.n41 171.744
R258 VTAIL.n42 VTAIL.n19 171.744
R259 VTAIL.n49 VTAIL.n19 171.744
R260 VTAIL.n50 VTAIL.n49 171.744
R261 VTAIL.n50 VTAIL.n15 171.744
R262 VTAIL.n57 VTAIL.n15 171.744
R263 VTAIL.n58 VTAIL.n57 171.744
R264 VTAIL.n58 VTAIL.n11 171.744
R265 VTAIL.n65 VTAIL.n11 171.744
R266 VTAIL.n66 VTAIL.n65 171.744
R267 VTAIL.n66 VTAIL.n7 171.744
R268 VTAIL.n74 VTAIL.n7 171.744
R269 VTAIL.n75 VTAIL.n74 171.744
R270 VTAIL.n76 VTAIL.n75 171.744
R271 VTAIL.n76 VTAIL.n3 171.744
R272 VTAIL.n83 VTAIL.n3 171.744
R273 VTAIL.n84 VTAIL.n83 171.744
R274 VTAIL.n123 VTAIL.n117 171.744
R275 VTAIL.n124 VTAIL.n123 171.744
R276 VTAIL.n124 VTAIL.n113 171.744
R277 VTAIL.n131 VTAIL.n113 171.744
R278 VTAIL.n132 VTAIL.n131 171.744
R279 VTAIL.n132 VTAIL.n109 171.744
R280 VTAIL.n139 VTAIL.n109 171.744
R281 VTAIL.n140 VTAIL.n139 171.744
R282 VTAIL.n140 VTAIL.n105 171.744
R283 VTAIL.n147 VTAIL.n105 171.744
R284 VTAIL.n148 VTAIL.n147 171.744
R285 VTAIL.n148 VTAIL.n101 171.744
R286 VTAIL.n155 VTAIL.n101 171.744
R287 VTAIL.n156 VTAIL.n155 171.744
R288 VTAIL.n156 VTAIL.n97 171.744
R289 VTAIL.n164 VTAIL.n97 171.744
R290 VTAIL.n165 VTAIL.n164 171.744
R291 VTAIL.n166 VTAIL.n165 171.744
R292 VTAIL.n166 VTAIL.n93 171.744
R293 VTAIL.n173 VTAIL.n93 171.744
R294 VTAIL.n174 VTAIL.n173 171.744
R295 VTAIL.n213 VTAIL.n207 171.744
R296 VTAIL.n214 VTAIL.n213 171.744
R297 VTAIL.n214 VTAIL.n203 171.744
R298 VTAIL.n221 VTAIL.n203 171.744
R299 VTAIL.n222 VTAIL.n221 171.744
R300 VTAIL.n222 VTAIL.n199 171.744
R301 VTAIL.n229 VTAIL.n199 171.744
R302 VTAIL.n230 VTAIL.n229 171.744
R303 VTAIL.n230 VTAIL.n195 171.744
R304 VTAIL.n237 VTAIL.n195 171.744
R305 VTAIL.n238 VTAIL.n237 171.744
R306 VTAIL.n238 VTAIL.n191 171.744
R307 VTAIL.n245 VTAIL.n191 171.744
R308 VTAIL.n246 VTAIL.n245 171.744
R309 VTAIL.n246 VTAIL.n187 171.744
R310 VTAIL.n254 VTAIL.n187 171.744
R311 VTAIL.n255 VTAIL.n254 171.744
R312 VTAIL.n256 VTAIL.n255 171.744
R313 VTAIL.n256 VTAIL.n183 171.744
R314 VTAIL.n263 VTAIL.n183 171.744
R315 VTAIL.n264 VTAIL.n263 171.744
R316 VTAIL.n624 VTAIL.n623 171.744
R317 VTAIL.n623 VTAIL.n543 171.744
R318 VTAIL.n616 VTAIL.n543 171.744
R319 VTAIL.n616 VTAIL.n615 171.744
R320 VTAIL.n615 VTAIL.n614 171.744
R321 VTAIL.n614 VTAIL.n547 171.744
R322 VTAIL.n607 VTAIL.n547 171.744
R323 VTAIL.n607 VTAIL.n606 171.744
R324 VTAIL.n606 VTAIL.n552 171.744
R325 VTAIL.n599 VTAIL.n552 171.744
R326 VTAIL.n599 VTAIL.n598 171.744
R327 VTAIL.n598 VTAIL.n556 171.744
R328 VTAIL.n591 VTAIL.n556 171.744
R329 VTAIL.n591 VTAIL.n590 171.744
R330 VTAIL.n590 VTAIL.n560 171.744
R331 VTAIL.n583 VTAIL.n560 171.744
R332 VTAIL.n583 VTAIL.n582 171.744
R333 VTAIL.n582 VTAIL.n564 171.744
R334 VTAIL.n575 VTAIL.n564 171.744
R335 VTAIL.n575 VTAIL.n574 171.744
R336 VTAIL.n574 VTAIL.n568 171.744
R337 VTAIL.n534 VTAIL.n533 171.744
R338 VTAIL.n533 VTAIL.n453 171.744
R339 VTAIL.n526 VTAIL.n453 171.744
R340 VTAIL.n526 VTAIL.n525 171.744
R341 VTAIL.n525 VTAIL.n524 171.744
R342 VTAIL.n524 VTAIL.n457 171.744
R343 VTAIL.n517 VTAIL.n457 171.744
R344 VTAIL.n517 VTAIL.n516 171.744
R345 VTAIL.n516 VTAIL.n462 171.744
R346 VTAIL.n509 VTAIL.n462 171.744
R347 VTAIL.n509 VTAIL.n508 171.744
R348 VTAIL.n508 VTAIL.n466 171.744
R349 VTAIL.n501 VTAIL.n466 171.744
R350 VTAIL.n501 VTAIL.n500 171.744
R351 VTAIL.n500 VTAIL.n470 171.744
R352 VTAIL.n493 VTAIL.n470 171.744
R353 VTAIL.n493 VTAIL.n492 171.744
R354 VTAIL.n492 VTAIL.n474 171.744
R355 VTAIL.n485 VTAIL.n474 171.744
R356 VTAIL.n485 VTAIL.n484 171.744
R357 VTAIL.n484 VTAIL.n478 171.744
R358 VTAIL.n444 VTAIL.n443 171.744
R359 VTAIL.n443 VTAIL.n363 171.744
R360 VTAIL.n436 VTAIL.n363 171.744
R361 VTAIL.n436 VTAIL.n435 171.744
R362 VTAIL.n435 VTAIL.n434 171.744
R363 VTAIL.n434 VTAIL.n367 171.744
R364 VTAIL.n427 VTAIL.n367 171.744
R365 VTAIL.n427 VTAIL.n426 171.744
R366 VTAIL.n426 VTAIL.n372 171.744
R367 VTAIL.n419 VTAIL.n372 171.744
R368 VTAIL.n419 VTAIL.n418 171.744
R369 VTAIL.n418 VTAIL.n376 171.744
R370 VTAIL.n411 VTAIL.n376 171.744
R371 VTAIL.n411 VTAIL.n410 171.744
R372 VTAIL.n410 VTAIL.n380 171.744
R373 VTAIL.n403 VTAIL.n380 171.744
R374 VTAIL.n403 VTAIL.n402 171.744
R375 VTAIL.n402 VTAIL.n384 171.744
R376 VTAIL.n395 VTAIL.n384 171.744
R377 VTAIL.n395 VTAIL.n394 171.744
R378 VTAIL.n394 VTAIL.n388 171.744
R379 VTAIL.n354 VTAIL.n353 171.744
R380 VTAIL.n353 VTAIL.n273 171.744
R381 VTAIL.n346 VTAIL.n273 171.744
R382 VTAIL.n346 VTAIL.n345 171.744
R383 VTAIL.n345 VTAIL.n344 171.744
R384 VTAIL.n344 VTAIL.n277 171.744
R385 VTAIL.n337 VTAIL.n277 171.744
R386 VTAIL.n337 VTAIL.n336 171.744
R387 VTAIL.n336 VTAIL.n282 171.744
R388 VTAIL.n329 VTAIL.n282 171.744
R389 VTAIL.n329 VTAIL.n328 171.744
R390 VTAIL.n328 VTAIL.n286 171.744
R391 VTAIL.n321 VTAIL.n286 171.744
R392 VTAIL.n321 VTAIL.n320 171.744
R393 VTAIL.n320 VTAIL.n290 171.744
R394 VTAIL.n313 VTAIL.n290 171.744
R395 VTAIL.n313 VTAIL.n312 171.744
R396 VTAIL.n312 VTAIL.n294 171.744
R397 VTAIL.n305 VTAIL.n294 171.744
R398 VTAIL.n305 VTAIL.n304 171.744
R399 VTAIL.n304 VTAIL.n298 171.744
R400 VTAIL.t3 VTAIL.n657 85.8723
R401 VTAIL.t0 VTAIL.n27 85.8723
R402 VTAIL.t6 VTAIL.n117 85.8723
R403 VTAIL.t4 VTAIL.n207 85.8723
R404 VTAIL.t5 VTAIL.n568 85.8723
R405 VTAIL.t7 VTAIL.n478 85.8723
R406 VTAIL.t1 VTAIL.n388 85.8723
R407 VTAIL.t2 VTAIL.n298 85.8723
R408 VTAIL.n719 VTAIL.n718 34.1247
R409 VTAIL.n89 VTAIL.n88 34.1247
R410 VTAIL.n179 VTAIL.n178 34.1247
R411 VTAIL.n269 VTAIL.n268 34.1247
R412 VTAIL.n629 VTAIL.n628 34.1247
R413 VTAIL.n539 VTAIL.n538 34.1247
R414 VTAIL.n449 VTAIL.n448 34.1247
R415 VTAIL.n359 VTAIL.n358 34.1247
R416 VTAIL.n719 VTAIL.n629 29.7117
R417 VTAIL.n359 VTAIL.n269 29.7117
R418 VTAIL.n659 VTAIL.n658 16.3895
R419 VTAIL.n29 VTAIL.n28 16.3895
R420 VTAIL.n119 VTAIL.n118 16.3895
R421 VTAIL.n209 VTAIL.n208 16.3895
R422 VTAIL.n570 VTAIL.n569 16.3895
R423 VTAIL.n480 VTAIL.n479 16.3895
R424 VTAIL.n390 VTAIL.n389 16.3895
R425 VTAIL.n300 VTAIL.n299 16.3895
R426 VTAIL.n707 VTAIL.n636 13.1884
R427 VTAIL.n77 VTAIL.n6 13.1884
R428 VTAIL.n167 VTAIL.n96 13.1884
R429 VTAIL.n257 VTAIL.n186 13.1884
R430 VTAIL.n617 VTAIL.n546 13.1884
R431 VTAIL.n527 VTAIL.n456 13.1884
R432 VTAIL.n437 VTAIL.n366 13.1884
R433 VTAIL.n347 VTAIL.n276 13.1884
R434 VTAIL.n662 VTAIL.n661 12.8005
R435 VTAIL.n703 VTAIL.n702 12.8005
R436 VTAIL.n708 VTAIL.n634 12.8005
R437 VTAIL.n32 VTAIL.n31 12.8005
R438 VTAIL.n73 VTAIL.n72 12.8005
R439 VTAIL.n78 VTAIL.n4 12.8005
R440 VTAIL.n122 VTAIL.n121 12.8005
R441 VTAIL.n163 VTAIL.n162 12.8005
R442 VTAIL.n168 VTAIL.n94 12.8005
R443 VTAIL.n212 VTAIL.n211 12.8005
R444 VTAIL.n253 VTAIL.n252 12.8005
R445 VTAIL.n258 VTAIL.n184 12.8005
R446 VTAIL.n618 VTAIL.n544 12.8005
R447 VTAIL.n613 VTAIL.n548 12.8005
R448 VTAIL.n573 VTAIL.n572 12.8005
R449 VTAIL.n528 VTAIL.n454 12.8005
R450 VTAIL.n523 VTAIL.n458 12.8005
R451 VTAIL.n483 VTAIL.n482 12.8005
R452 VTAIL.n438 VTAIL.n364 12.8005
R453 VTAIL.n433 VTAIL.n368 12.8005
R454 VTAIL.n393 VTAIL.n392 12.8005
R455 VTAIL.n348 VTAIL.n274 12.8005
R456 VTAIL.n343 VTAIL.n278 12.8005
R457 VTAIL.n303 VTAIL.n302 12.8005
R458 VTAIL.n665 VTAIL.n656 12.0247
R459 VTAIL.n701 VTAIL.n638 12.0247
R460 VTAIL.n712 VTAIL.n711 12.0247
R461 VTAIL.n35 VTAIL.n26 12.0247
R462 VTAIL.n71 VTAIL.n8 12.0247
R463 VTAIL.n82 VTAIL.n81 12.0247
R464 VTAIL.n125 VTAIL.n116 12.0247
R465 VTAIL.n161 VTAIL.n98 12.0247
R466 VTAIL.n172 VTAIL.n171 12.0247
R467 VTAIL.n215 VTAIL.n206 12.0247
R468 VTAIL.n251 VTAIL.n188 12.0247
R469 VTAIL.n262 VTAIL.n261 12.0247
R470 VTAIL.n622 VTAIL.n621 12.0247
R471 VTAIL.n612 VTAIL.n549 12.0247
R472 VTAIL.n576 VTAIL.n567 12.0247
R473 VTAIL.n532 VTAIL.n531 12.0247
R474 VTAIL.n522 VTAIL.n459 12.0247
R475 VTAIL.n486 VTAIL.n477 12.0247
R476 VTAIL.n442 VTAIL.n441 12.0247
R477 VTAIL.n432 VTAIL.n369 12.0247
R478 VTAIL.n396 VTAIL.n387 12.0247
R479 VTAIL.n352 VTAIL.n351 12.0247
R480 VTAIL.n342 VTAIL.n279 12.0247
R481 VTAIL.n306 VTAIL.n297 12.0247
R482 VTAIL.n666 VTAIL.n654 11.249
R483 VTAIL.n698 VTAIL.n697 11.249
R484 VTAIL.n715 VTAIL.n632 11.249
R485 VTAIL.n36 VTAIL.n24 11.249
R486 VTAIL.n68 VTAIL.n67 11.249
R487 VTAIL.n85 VTAIL.n2 11.249
R488 VTAIL.n126 VTAIL.n114 11.249
R489 VTAIL.n158 VTAIL.n157 11.249
R490 VTAIL.n175 VTAIL.n92 11.249
R491 VTAIL.n216 VTAIL.n204 11.249
R492 VTAIL.n248 VTAIL.n247 11.249
R493 VTAIL.n265 VTAIL.n182 11.249
R494 VTAIL.n625 VTAIL.n542 11.249
R495 VTAIL.n609 VTAIL.n608 11.249
R496 VTAIL.n577 VTAIL.n565 11.249
R497 VTAIL.n535 VTAIL.n452 11.249
R498 VTAIL.n519 VTAIL.n518 11.249
R499 VTAIL.n487 VTAIL.n475 11.249
R500 VTAIL.n445 VTAIL.n362 11.249
R501 VTAIL.n429 VTAIL.n428 11.249
R502 VTAIL.n397 VTAIL.n385 11.249
R503 VTAIL.n355 VTAIL.n272 11.249
R504 VTAIL.n339 VTAIL.n338 11.249
R505 VTAIL.n307 VTAIL.n295 11.249
R506 VTAIL.n670 VTAIL.n669 10.4732
R507 VTAIL.n694 VTAIL.n640 10.4732
R508 VTAIL.n716 VTAIL.n630 10.4732
R509 VTAIL.n40 VTAIL.n39 10.4732
R510 VTAIL.n64 VTAIL.n10 10.4732
R511 VTAIL.n86 VTAIL.n0 10.4732
R512 VTAIL.n130 VTAIL.n129 10.4732
R513 VTAIL.n154 VTAIL.n100 10.4732
R514 VTAIL.n176 VTAIL.n90 10.4732
R515 VTAIL.n220 VTAIL.n219 10.4732
R516 VTAIL.n244 VTAIL.n190 10.4732
R517 VTAIL.n266 VTAIL.n180 10.4732
R518 VTAIL.n626 VTAIL.n540 10.4732
R519 VTAIL.n605 VTAIL.n551 10.4732
R520 VTAIL.n581 VTAIL.n580 10.4732
R521 VTAIL.n536 VTAIL.n450 10.4732
R522 VTAIL.n515 VTAIL.n461 10.4732
R523 VTAIL.n491 VTAIL.n490 10.4732
R524 VTAIL.n446 VTAIL.n360 10.4732
R525 VTAIL.n425 VTAIL.n371 10.4732
R526 VTAIL.n401 VTAIL.n400 10.4732
R527 VTAIL.n356 VTAIL.n270 10.4732
R528 VTAIL.n335 VTAIL.n281 10.4732
R529 VTAIL.n311 VTAIL.n310 10.4732
R530 VTAIL.n673 VTAIL.n652 9.69747
R531 VTAIL.n693 VTAIL.n642 9.69747
R532 VTAIL.n43 VTAIL.n22 9.69747
R533 VTAIL.n63 VTAIL.n12 9.69747
R534 VTAIL.n133 VTAIL.n112 9.69747
R535 VTAIL.n153 VTAIL.n102 9.69747
R536 VTAIL.n223 VTAIL.n202 9.69747
R537 VTAIL.n243 VTAIL.n192 9.69747
R538 VTAIL.n604 VTAIL.n553 9.69747
R539 VTAIL.n584 VTAIL.n563 9.69747
R540 VTAIL.n514 VTAIL.n463 9.69747
R541 VTAIL.n494 VTAIL.n473 9.69747
R542 VTAIL.n424 VTAIL.n373 9.69747
R543 VTAIL.n404 VTAIL.n383 9.69747
R544 VTAIL.n334 VTAIL.n283 9.69747
R545 VTAIL.n314 VTAIL.n293 9.69747
R546 VTAIL.n718 VTAIL.n717 9.45567
R547 VTAIL.n88 VTAIL.n87 9.45567
R548 VTAIL.n178 VTAIL.n177 9.45567
R549 VTAIL.n268 VTAIL.n267 9.45567
R550 VTAIL.n628 VTAIL.n627 9.45567
R551 VTAIL.n538 VTAIL.n537 9.45567
R552 VTAIL.n448 VTAIL.n447 9.45567
R553 VTAIL.n358 VTAIL.n357 9.45567
R554 VTAIL.n717 VTAIL.n716 9.3005
R555 VTAIL.n632 VTAIL.n631 9.3005
R556 VTAIL.n711 VTAIL.n710 9.3005
R557 VTAIL.n709 VTAIL.n708 9.3005
R558 VTAIL.n648 VTAIL.n647 9.3005
R559 VTAIL.n677 VTAIL.n676 9.3005
R560 VTAIL.n675 VTAIL.n674 9.3005
R561 VTAIL.n652 VTAIL.n651 9.3005
R562 VTAIL.n669 VTAIL.n668 9.3005
R563 VTAIL.n667 VTAIL.n666 9.3005
R564 VTAIL.n656 VTAIL.n655 9.3005
R565 VTAIL.n661 VTAIL.n660 9.3005
R566 VTAIL.n683 VTAIL.n682 9.3005
R567 VTAIL.n685 VTAIL.n684 9.3005
R568 VTAIL.n644 VTAIL.n643 9.3005
R569 VTAIL.n691 VTAIL.n690 9.3005
R570 VTAIL.n693 VTAIL.n692 9.3005
R571 VTAIL.n640 VTAIL.n639 9.3005
R572 VTAIL.n699 VTAIL.n698 9.3005
R573 VTAIL.n701 VTAIL.n700 9.3005
R574 VTAIL.n702 VTAIL.n635 9.3005
R575 VTAIL.n87 VTAIL.n86 9.3005
R576 VTAIL.n2 VTAIL.n1 9.3005
R577 VTAIL.n81 VTAIL.n80 9.3005
R578 VTAIL.n79 VTAIL.n78 9.3005
R579 VTAIL.n18 VTAIL.n17 9.3005
R580 VTAIL.n47 VTAIL.n46 9.3005
R581 VTAIL.n45 VTAIL.n44 9.3005
R582 VTAIL.n22 VTAIL.n21 9.3005
R583 VTAIL.n39 VTAIL.n38 9.3005
R584 VTAIL.n37 VTAIL.n36 9.3005
R585 VTAIL.n26 VTAIL.n25 9.3005
R586 VTAIL.n31 VTAIL.n30 9.3005
R587 VTAIL.n53 VTAIL.n52 9.3005
R588 VTAIL.n55 VTAIL.n54 9.3005
R589 VTAIL.n14 VTAIL.n13 9.3005
R590 VTAIL.n61 VTAIL.n60 9.3005
R591 VTAIL.n63 VTAIL.n62 9.3005
R592 VTAIL.n10 VTAIL.n9 9.3005
R593 VTAIL.n69 VTAIL.n68 9.3005
R594 VTAIL.n71 VTAIL.n70 9.3005
R595 VTAIL.n72 VTAIL.n5 9.3005
R596 VTAIL.n177 VTAIL.n176 9.3005
R597 VTAIL.n92 VTAIL.n91 9.3005
R598 VTAIL.n171 VTAIL.n170 9.3005
R599 VTAIL.n169 VTAIL.n168 9.3005
R600 VTAIL.n108 VTAIL.n107 9.3005
R601 VTAIL.n137 VTAIL.n136 9.3005
R602 VTAIL.n135 VTAIL.n134 9.3005
R603 VTAIL.n112 VTAIL.n111 9.3005
R604 VTAIL.n129 VTAIL.n128 9.3005
R605 VTAIL.n127 VTAIL.n126 9.3005
R606 VTAIL.n116 VTAIL.n115 9.3005
R607 VTAIL.n121 VTAIL.n120 9.3005
R608 VTAIL.n143 VTAIL.n142 9.3005
R609 VTAIL.n145 VTAIL.n144 9.3005
R610 VTAIL.n104 VTAIL.n103 9.3005
R611 VTAIL.n151 VTAIL.n150 9.3005
R612 VTAIL.n153 VTAIL.n152 9.3005
R613 VTAIL.n100 VTAIL.n99 9.3005
R614 VTAIL.n159 VTAIL.n158 9.3005
R615 VTAIL.n161 VTAIL.n160 9.3005
R616 VTAIL.n162 VTAIL.n95 9.3005
R617 VTAIL.n267 VTAIL.n266 9.3005
R618 VTAIL.n182 VTAIL.n181 9.3005
R619 VTAIL.n261 VTAIL.n260 9.3005
R620 VTAIL.n259 VTAIL.n258 9.3005
R621 VTAIL.n198 VTAIL.n197 9.3005
R622 VTAIL.n227 VTAIL.n226 9.3005
R623 VTAIL.n225 VTAIL.n224 9.3005
R624 VTAIL.n202 VTAIL.n201 9.3005
R625 VTAIL.n219 VTAIL.n218 9.3005
R626 VTAIL.n217 VTAIL.n216 9.3005
R627 VTAIL.n206 VTAIL.n205 9.3005
R628 VTAIL.n211 VTAIL.n210 9.3005
R629 VTAIL.n233 VTAIL.n232 9.3005
R630 VTAIL.n235 VTAIL.n234 9.3005
R631 VTAIL.n194 VTAIL.n193 9.3005
R632 VTAIL.n241 VTAIL.n240 9.3005
R633 VTAIL.n243 VTAIL.n242 9.3005
R634 VTAIL.n190 VTAIL.n189 9.3005
R635 VTAIL.n249 VTAIL.n248 9.3005
R636 VTAIL.n251 VTAIL.n250 9.3005
R637 VTAIL.n252 VTAIL.n185 9.3005
R638 VTAIL.n596 VTAIL.n595 9.3005
R639 VTAIL.n555 VTAIL.n554 9.3005
R640 VTAIL.n602 VTAIL.n601 9.3005
R641 VTAIL.n604 VTAIL.n603 9.3005
R642 VTAIL.n551 VTAIL.n550 9.3005
R643 VTAIL.n610 VTAIL.n609 9.3005
R644 VTAIL.n612 VTAIL.n611 9.3005
R645 VTAIL.n548 VTAIL.n545 9.3005
R646 VTAIL.n627 VTAIL.n626 9.3005
R647 VTAIL.n542 VTAIL.n541 9.3005
R648 VTAIL.n621 VTAIL.n620 9.3005
R649 VTAIL.n619 VTAIL.n618 9.3005
R650 VTAIL.n594 VTAIL.n593 9.3005
R651 VTAIL.n559 VTAIL.n558 9.3005
R652 VTAIL.n588 VTAIL.n587 9.3005
R653 VTAIL.n586 VTAIL.n585 9.3005
R654 VTAIL.n563 VTAIL.n562 9.3005
R655 VTAIL.n580 VTAIL.n579 9.3005
R656 VTAIL.n578 VTAIL.n577 9.3005
R657 VTAIL.n567 VTAIL.n566 9.3005
R658 VTAIL.n572 VTAIL.n571 9.3005
R659 VTAIL.n506 VTAIL.n505 9.3005
R660 VTAIL.n465 VTAIL.n464 9.3005
R661 VTAIL.n512 VTAIL.n511 9.3005
R662 VTAIL.n514 VTAIL.n513 9.3005
R663 VTAIL.n461 VTAIL.n460 9.3005
R664 VTAIL.n520 VTAIL.n519 9.3005
R665 VTAIL.n522 VTAIL.n521 9.3005
R666 VTAIL.n458 VTAIL.n455 9.3005
R667 VTAIL.n537 VTAIL.n536 9.3005
R668 VTAIL.n452 VTAIL.n451 9.3005
R669 VTAIL.n531 VTAIL.n530 9.3005
R670 VTAIL.n529 VTAIL.n528 9.3005
R671 VTAIL.n504 VTAIL.n503 9.3005
R672 VTAIL.n469 VTAIL.n468 9.3005
R673 VTAIL.n498 VTAIL.n497 9.3005
R674 VTAIL.n496 VTAIL.n495 9.3005
R675 VTAIL.n473 VTAIL.n472 9.3005
R676 VTAIL.n490 VTAIL.n489 9.3005
R677 VTAIL.n488 VTAIL.n487 9.3005
R678 VTAIL.n477 VTAIL.n476 9.3005
R679 VTAIL.n482 VTAIL.n481 9.3005
R680 VTAIL.n416 VTAIL.n415 9.3005
R681 VTAIL.n375 VTAIL.n374 9.3005
R682 VTAIL.n422 VTAIL.n421 9.3005
R683 VTAIL.n424 VTAIL.n423 9.3005
R684 VTAIL.n371 VTAIL.n370 9.3005
R685 VTAIL.n430 VTAIL.n429 9.3005
R686 VTAIL.n432 VTAIL.n431 9.3005
R687 VTAIL.n368 VTAIL.n365 9.3005
R688 VTAIL.n447 VTAIL.n446 9.3005
R689 VTAIL.n362 VTAIL.n361 9.3005
R690 VTAIL.n441 VTAIL.n440 9.3005
R691 VTAIL.n439 VTAIL.n438 9.3005
R692 VTAIL.n414 VTAIL.n413 9.3005
R693 VTAIL.n379 VTAIL.n378 9.3005
R694 VTAIL.n408 VTAIL.n407 9.3005
R695 VTAIL.n406 VTAIL.n405 9.3005
R696 VTAIL.n383 VTAIL.n382 9.3005
R697 VTAIL.n400 VTAIL.n399 9.3005
R698 VTAIL.n398 VTAIL.n397 9.3005
R699 VTAIL.n387 VTAIL.n386 9.3005
R700 VTAIL.n392 VTAIL.n391 9.3005
R701 VTAIL.n326 VTAIL.n325 9.3005
R702 VTAIL.n285 VTAIL.n284 9.3005
R703 VTAIL.n332 VTAIL.n331 9.3005
R704 VTAIL.n334 VTAIL.n333 9.3005
R705 VTAIL.n281 VTAIL.n280 9.3005
R706 VTAIL.n340 VTAIL.n339 9.3005
R707 VTAIL.n342 VTAIL.n341 9.3005
R708 VTAIL.n278 VTAIL.n275 9.3005
R709 VTAIL.n357 VTAIL.n356 9.3005
R710 VTAIL.n272 VTAIL.n271 9.3005
R711 VTAIL.n351 VTAIL.n350 9.3005
R712 VTAIL.n349 VTAIL.n348 9.3005
R713 VTAIL.n324 VTAIL.n323 9.3005
R714 VTAIL.n289 VTAIL.n288 9.3005
R715 VTAIL.n318 VTAIL.n317 9.3005
R716 VTAIL.n316 VTAIL.n315 9.3005
R717 VTAIL.n293 VTAIL.n292 9.3005
R718 VTAIL.n310 VTAIL.n309 9.3005
R719 VTAIL.n308 VTAIL.n307 9.3005
R720 VTAIL.n297 VTAIL.n296 9.3005
R721 VTAIL.n302 VTAIL.n301 9.3005
R722 VTAIL.n674 VTAIL.n650 8.92171
R723 VTAIL.n690 VTAIL.n689 8.92171
R724 VTAIL.n44 VTAIL.n20 8.92171
R725 VTAIL.n60 VTAIL.n59 8.92171
R726 VTAIL.n134 VTAIL.n110 8.92171
R727 VTAIL.n150 VTAIL.n149 8.92171
R728 VTAIL.n224 VTAIL.n200 8.92171
R729 VTAIL.n240 VTAIL.n239 8.92171
R730 VTAIL.n601 VTAIL.n600 8.92171
R731 VTAIL.n585 VTAIL.n561 8.92171
R732 VTAIL.n511 VTAIL.n510 8.92171
R733 VTAIL.n495 VTAIL.n471 8.92171
R734 VTAIL.n421 VTAIL.n420 8.92171
R735 VTAIL.n405 VTAIL.n381 8.92171
R736 VTAIL.n331 VTAIL.n330 8.92171
R737 VTAIL.n315 VTAIL.n291 8.92171
R738 VTAIL.n678 VTAIL.n677 8.14595
R739 VTAIL.n686 VTAIL.n644 8.14595
R740 VTAIL.n48 VTAIL.n47 8.14595
R741 VTAIL.n56 VTAIL.n14 8.14595
R742 VTAIL.n138 VTAIL.n137 8.14595
R743 VTAIL.n146 VTAIL.n104 8.14595
R744 VTAIL.n228 VTAIL.n227 8.14595
R745 VTAIL.n236 VTAIL.n194 8.14595
R746 VTAIL.n597 VTAIL.n555 8.14595
R747 VTAIL.n589 VTAIL.n588 8.14595
R748 VTAIL.n507 VTAIL.n465 8.14595
R749 VTAIL.n499 VTAIL.n498 8.14595
R750 VTAIL.n417 VTAIL.n375 8.14595
R751 VTAIL.n409 VTAIL.n408 8.14595
R752 VTAIL.n327 VTAIL.n285 8.14595
R753 VTAIL.n319 VTAIL.n318 8.14595
R754 VTAIL.n681 VTAIL.n648 7.3702
R755 VTAIL.n685 VTAIL.n646 7.3702
R756 VTAIL.n51 VTAIL.n18 7.3702
R757 VTAIL.n55 VTAIL.n16 7.3702
R758 VTAIL.n141 VTAIL.n108 7.3702
R759 VTAIL.n145 VTAIL.n106 7.3702
R760 VTAIL.n231 VTAIL.n198 7.3702
R761 VTAIL.n235 VTAIL.n196 7.3702
R762 VTAIL.n596 VTAIL.n557 7.3702
R763 VTAIL.n592 VTAIL.n559 7.3702
R764 VTAIL.n506 VTAIL.n467 7.3702
R765 VTAIL.n502 VTAIL.n469 7.3702
R766 VTAIL.n416 VTAIL.n377 7.3702
R767 VTAIL.n412 VTAIL.n379 7.3702
R768 VTAIL.n326 VTAIL.n287 7.3702
R769 VTAIL.n322 VTAIL.n289 7.3702
R770 VTAIL.n682 VTAIL.n681 6.59444
R771 VTAIL.n682 VTAIL.n646 6.59444
R772 VTAIL.n52 VTAIL.n51 6.59444
R773 VTAIL.n52 VTAIL.n16 6.59444
R774 VTAIL.n142 VTAIL.n141 6.59444
R775 VTAIL.n142 VTAIL.n106 6.59444
R776 VTAIL.n232 VTAIL.n231 6.59444
R777 VTAIL.n232 VTAIL.n196 6.59444
R778 VTAIL.n593 VTAIL.n557 6.59444
R779 VTAIL.n593 VTAIL.n592 6.59444
R780 VTAIL.n503 VTAIL.n467 6.59444
R781 VTAIL.n503 VTAIL.n502 6.59444
R782 VTAIL.n413 VTAIL.n377 6.59444
R783 VTAIL.n413 VTAIL.n412 6.59444
R784 VTAIL.n323 VTAIL.n287 6.59444
R785 VTAIL.n323 VTAIL.n322 6.59444
R786 VTAIL.n678 VTAIL.n648 5.81868
R787 VTAIL.n686 VTAIL.n685 5.81868
R788 VTAIL.n48 VTAIL.n18 5.81868
R789 VTAIL.n56 VTAIL.n55 5.81868
R790 VTAIL.n138 VTAIL.n108 5.81868
R791 VTAIL.n146 VTAIL.n145 5.81868
R792 VTAIL.n228 VTAIL.n198 5.81868
R793 VTAIL.n236 VTAIL.n235 5.81868
R794 VTAIL.n597 VTAIL.n596 5.81868
R795 VTAIL.n589 VTAIL.n559 5.81868
R796 VTAIL.n507 VTAIL.n506 5.81868
R797 VTAIL.n499 VTAIL.n469 5.81868
R798 VTAIL.n417 VTAIL.n416 5.81868
R799 VTAIL.n409 VTAIL.n379 5.81868
R800 VTAIL.n327 VTAIL.n326 5.81868
R801 VTAIL.n319 VTAIL.n289 5.81868
R802 VTAIL.n677 VTAIL.n650 5.04292
R803 VTAIL.n689 VTAIL.n644 5.04292
R804 VTAIL.n47 VTAIL.n20 5.04292
R805 VTAIL.n59 VTAIL.n14 5.04292
R806 VTAIL.n137 VTAIL.n110 5.04292
R807 VTAIL.n149 VTAIL.n104 5.04292
R808 VTAIL.n227 VTAIL.n200 5.04292
R809 VTAIL.n239 VTAIL.n194 5.04292
R810 VTAIL.n600 VTAIL.n555 5.04292
R811 VTAIL.n588 VTAIL.n561 5.04292
R812 VTAIL.n510 VTAIL.n465 5.04292
R813 VTAIL.n498 VTAIL.n471 5.04292
R814 VTAIL.n420 VTAIL.n375 5.04292
R815 VTAIL.n408 VTAIL.n381 5.04292
R816 VTAIL.n330 VTAIL.n285 5.04292
R817 VTAIL.n318 VTAIL.n291 5.04292
R818 VTAIL.n674 VTAIL.n673 4.26717
R819 VTAIL.n690 VTAIL.n642 4.26717
R820 VTAIL.n44 VTAIL.n43 4.26717
R821 VTAIL.n60 VTAIL.n12 4.26717
R822 VTAIL.n134 VTAIL.n133 4.26717
R823 VTAIL.n150 VTAIL.n102 4.26717
R824 VTAIL.n224 VTAIL.n223 4.26717
R825 VTAIL.n240 VTAIL.n192 4.26717
R826 VTAIL.n601 VTAIL.n553 4.26717
R827 VTAIL.n585 VTAIL.n584 4.26717
R828 VTAIL.n511 VTAIL.n463 4.26717
R829 VTAIL.n495 VTAIL.n494 4.26717
R830 VTAIL.n421 VTAIL.n373 4.26717
R831 VTAIL.n405 VTAIL.n404 4.26717
R832 VTAIL.n331 VTAIL.n283 4.26717
R833 VTAIL.n315 VTAIL.n314 4.26717
R834 VTAIL.n660 VTAIL.n659 3.70982
R835 VTAIL.n30 VTAIL.n29 3.70982
R836 VTAIL.n120 VTAIL.n119 3.70982
R837 VTAIL.n210 VTAIL.n209 3.70982
R838 VTAIL.n571 VTAIL.n570 3.70982
R839 VTAIL.n481 VTAIL.n480 3.70982
R840 VTAIL.n391 VTAIL.n390 3.70982
R841 VTAIL.n301 VTAIL.n300 3.70982
R842 VTAIL.n670 VTAIL.n652 3.49141
R843 VTAIL.n694 VTAIL.n693 3.49141
R844 VTAIL.n718 VTAIL.n630 3.49141
R845 VTAIL.n40 VTAIL.n22 3.49141
R846 VTAIL.n64 VTAIL.n63 3.49141
R847 VTAIL.n88 VTAIL.n0 3.49141
R848 VTAIL.n130 VTAIL.n112 3.49141
R849 VTAIL.n154 VTAIL.n153 3.49141
R850 VTAIL.n178 VTAIL.n90 3.49141
R851 VTAIL.n220 VTAIL.n202 3.49141
R852 VTAIL.n244 VTAIL.n243 3.49141
R853 VTAIL.n268 VTAIL.n180 3.49141
R854 VTAIL.n628 VTAIL.n540 3.49141
R855 VTAIL.n605 VTAIL.n604 3.49141
R856 VTAIL.n581 VTAIL.n563 3.49141
R857 VTAIL.n538 VTAIL.n450 3.49141
R858 VTAIL.n515 VTAIL.n514 3.49141
R859 VTAIL.n491 VTAIL.n473 3.49141
R860 VTAIL.n448 VTAIL.n360 3.49141
R861 VTAIL.n425 VTAIL.n424 3.49141
R862 VTAIL.n401 VTAIL.n383 3.49141
R863 VTAIL.n358 VTAIL.n270 3.49141
R864 VTAIL.n335 VTAIL.n334 3.49141
R865 VTAIL.n311 VTAIL.n293 3.49141
R866 VTAIL.n449 VTAIL.n359 3.39705
R867 VTAIL.n629 VTAIL.n539 3.39705
R868 VTAIL.n269 VTAIL.n179 3.39705
R869 VTAIL.n669 VTAIL.n654 2.71565
R870 VTAIL.n697 VTAIL.n640 2.71565
R871 VTAIL.n716 VTAIL.n715 2.71565
R872 VTAIL.n39 VTAIL.n24 2.71565
R873 VTAIL.n67 VTAIL.n10 2.71565
R874 VTAIL.n86 VTAIL.n85 2.71565
R875 VTAIL.n129 VTAIL.n114 2.71565
R876 VTAIL.n157 VTAIL.n100 2.71565
R877 VTAIL.n176 VTAIL.n175 2.71565
R878 VTAIL.n219 VTAIL.n204 2.71565
R879 VTAIL.n247 VTAIL.n190 2.71565
R880 VTAIL.n266 VTAIL.n265 2.71565
R881 VTAIL.n626 VTAIL.n625 2.71565
R882 VTAIL.n608 VTAIL.n551 2.71565
R883 VTAIL.n580 VTAIL.n565 2.71565
R884 VTAIL.n536 VTAIL.n535 2.71565
R885 VTAIL.n518 VTAIL.n461 2.71565
R886 VTAIL.n490 VTAIL.n475 2.71565
R887 VTAIL.n446 VTAIL.n445 2.71565
R888 VTAIL.n428 VTAIL.n371 2.71565
R889 VTAIL.n400 VTAIL.n385 2.71565
R890 VTAIL.n356 VTAIL.n355 2.71565
R891 VTAIL.n338 VTAIL.n281 2.71565
R892 VTAIL.n310 VTAIL.n295 2.71565
R893 VTAIL.n666 VTAIL.n665 1.93989
R894 VTAIL.n698 VTAIL.n638 1.93989
R895 VTAIL.n712 VTAIL.n632 1.93989
R896 VTAIL.n36 VTAIL.n35 1.93989
R897 VTAIL.n68 VTAIL.n8 1.93989
R898 VTAIL.n82 VTAIL.n2 1.93989
R899 VTAIL.n126 VTAIL.n125 1.93989
R900 VTAIL.n158 VTAIL.n98 1.93989
R901 VTAIL.n172 VTAIL.n92 1.93989
R902 VTAIL.n216 VTAIL.n215 1.93989
R903 VTAIL.n248 VTAIL.n188 1.93989
R904 VTAIL.n262 VTAIL.n182 1.93989
R905 VTAIL.n622 VTAIL.n542 1.93989
R906 VTAIL.n609 VTAIL.n549 1.93989
R907 VTAIL.n577 VTAIL.n576 1.93989
R908 VTAIL.n532 VTAIL.n452 1.93989
R909 VTAIL.n519 VTAIL.n459 1.93989
R910 VTAIL.n487 VTAIL.n486 1.93989
R911 VTAIL.n442 VTAIL.n362 1.93989
R912 VTAIL.n429 VTAIL.n369 1.93989
R913 VTAIL.n397 VTAIL.n396 1.93989
R914 VTAIL.n352 VTAIL.n272 1.93989
R915 VTAIL.n339 VTAIL.n279 1.93989
R916 VTAIL.n307 VTAIL.n306 1.93989
R917 VTAIL VTAIL.n89 1.75697
R918 VTAIL VTAIL.n719 1.64059
R919 VTAIL.n662 VTAIL.n656 1.16414
R920 VTAIL.n703 VTAIL.n701 1.16414
R921 VTAIL.n711 VTAIL.n634 1.16414
R922 VTAIL.n32 VTAIL.n26 1.16414
R923 VTAIL.n73 VTAIL.n71 1.16414
R924 VTAIL.n81 VTAIL.n4 1.16414
R925 VTAIL.n122 VTAIL.n116 1.16414
R926 VTAIL.n163 VTAIL.n161 1.16414
R927 VTAIL.n171 VTAIL.n94 1.16414
R928 VTAIL.n212 VTAIL.n206 1.16414
R929 VTAIL.n253 VTAIL.n251 1.16414
R930 VTAIL.n261 VTAIL.n184 1.16414
R931 VTAIL.n621 VTAIL.n544 1.16414
R932 VTAIL.n613 VTAIL.n612 1.16414
R933 VTAIL.n573 VTAIL.n567 1.16414
R934 VTAIL.n531 VTAIL.n454 1.16414
R935 VTAIL.n523 VTAIL.n522 1.16414
R936 VTAIL.n483 VTAIL.n477 1.16414
R937 VTAIL.n441 VTAIL.n364 1.16414
R938 VTAIL.n433 VTAIL.n432 1.16414
R939 VTAIL.n393 VTAIL.n387 1.16414
R940 VTAIL.n351 VTAIL.n274 1.16414
R941 VTAIL.n343 VTAIL.n342 1.16414
R942 VTAIL.n303 VTAIL.n297 1.16414
R943 VTAIL.n539 VTAIL.n449 0.470328
R944 VTAIL.n179 VTAIL.n89 0.470328
R945 VTAIL.n661 VTAIL.n658 0.388379
R946 VTAIL.n702 VTAIL.n636 0.388379
R947 VTAIL.n708 VTAIL.n707 0.388379
R948 VTAIL.n31 VTAIL.n28 0.388379
R949 VTAIL.n72 VTAIL.n6 0.388379
R950 VTAIL.n78 VTAIL.n77 0.388379
R951 VTAIL.n121 VTAIL.n118 0.388379
R952 VTAIL.n162 VTAIL.n96 0.388379
R953 VTAIL.n168 VTAIL.n167 0.388379
R954 VTAIL.n211 VTAIL.n208 0.388379
R955 VTAIL.n252 VTAIL.n186 0.388379
R956 VTAIL.n258 VTAIL.n257 0.388379
R957 VTAIL.n618 VTAIL.n617 0.388379
R958 VTAIL.n548 VTAIL.n546 0.388379
R959 VTAIL.n572 VTAIL.n569 0.388379
R960 VTAIL.n528 VTAIL.n527 0.388379
R961 VTAIL.n458 VTAIL.n456 0.388379
R962 VTAIL.n482 VTAIL.n479 0.388379
R963 VTAIL.n438 VTAIL.n437 0.388379
R964 VTAIL.n368 VTAIL.n366 0.388379
R965 VTAIL.n392 VTAIL.n389 0.388379
R966 VTAIL.n348 VTAIL.n347 0.388379
R967 VTAIL.n278 VTAIL.n276 0.388379
R968 VTAIL.n302 VTAIL.n299 0.388379
R969 VTAIL.n660 VTAIL.n655 0.155672
R970 VTAIL.n667 VTAIL.n655 0.155672
R971 VTAIL.n668 VTAIL.n667 0.155672
R972 VTAIL.n668 VTAIL.n651 0.155672
R973 VTAIL.n675 VTAIL.n651 0.155672
R974 VTAIL.n676 VTAIL.n675 0.155672
R975 VTAIL.n676 VTAIL.n647 0.155672
R976 VTAIL.n683 VTAIL.n647 0.155672
R977 VTAIL.n684 VTAIL.n683 0.155672
R978 VTAIL.n684 VTAIL.n643 0.155672
R979 VTAIL.n691 VTAIL.n643 0.155672
R980 VTAIL.n692 VTAIL.n691 0.155672
R981 VTAIL.n692 VTAIL.n639 0.155672
R982 VTAIL.n699 VTAIL.n639 0.155672
R983 VTAIL.n700 VTAIL.n699 0.155672
R984 VTAIL.n700 VTAIL.n635 0.155672
R985 VTAIL.n709 VTAIL.n635 0.155672
R986 VTAIL.n710 VTAIL.n709 0.155672
R987 VTAIL.n710 VTAIL.n631 0.155672
R988 VTAIL.n717 VTAIL.n631 0.155672
R989 VTAIL.n30 VTAIL.n25 0.155672
R990 VTAIL.n37 VTAIL.n25 0.155672
R991 VTAIL.n38 VTAIL.n37 0.155672
R992 VTAIL.n38 VTAIL.n21 0.155672
R993 VTAIL.n45 VTAIL.n21 0.155672
R994 VTAIL.n46 VTAIL.n45 0.155672
R995 VTAIL.n46 VTAIL.n17 0.155672
R996 VTAIL.n53 VTAIL.n17 0.155672
R997 VTAIL.n54 VTAIL.n53 0.155672
R998 VTAIL.n54 VTAIL.n13 0.155672
R999 VTAIL.n61 VTAIL.n13 0.155672
R1000 VTAIL.n62 VTAIL.n61 0.155672
R1001 VTAIL.n62 VTAIL.n9 0.155672
R1002 VTAIL.n69 VTAIL.n9 0.155672
R1003 VTAIL.n70 VTAIL.n69 0.155672
R1004 VTAIL.n70 VTAIL.n5 0.155672
R1005 VTAIL.n79 VTAIL.n5 0.155672
R1006 VTAIL.n80 VTAIL.n79 0.155672
R1007 VTAIL.n80 VTAIL.n1 0.155672
R1008 VTAIL.n87 VTAIL.n1 0.155672
R1009 VTAIL.n120 VTAIL.n115 0.155672
R1010 VTAIL.n127 VTAIL.n115 0.155672
R1011 VTAIL.n128 VTAIL.n127 0.155672
R1012 VTAIL.n128 VTAIL.n111 0.155672
R1013 VTAIL.n135 VTAIL.n111 0.155672
R1014 VTAIL.n136 VTAIL.n135 0.155672
R1015 VTAIL.n136 VTAIL.n107 0.155672
R1016 VTAIL.n143 VTAIL.n107 0.155672
R1017 VTAIL.n144 VTAIL.n143 0.155672
R1018 VTAIL.n144 VTAIL.n103 0.155672
R1019 VTAIL.n151 VTAIL.n103 0.155672
R1020 VTAIL.n152 VTAIL.n151 0.155672
R1021 VTAIL.n152 VTAIL.n99 0.155672
R1022 VTAIL.n159 VTAIL.n99 0.155672
R1023 VTAIL.n160 VTAIL.n159 0.155672
R1024 VTAIL.n160 VTAIL.n95 0.155672
R1025 VTAIL.n169 VTAIL.n95 0.155672
R1026 VTAIL.n170 VTAIL.n169 0.155672
R1027 VTAIL.n170 VTAIL.n91 0.155672
R1028 VTAIL.n177 VTAIL.n91 0.155672
R1029 VTAIL.n210 VTAIL.n205 0.155672
R1030 VTAIL.n217 VTAIL.n205 0.155672
R1031 VTAIL.n218 VTAIL.n217 0.155672
R1032 VTAIL.n218 VTAIL.n201 0.155672
R1033 VTAIL.n225 VTAIL.n201 0.155672
R1034 VTAIL.n226 VTAIL.n225 0.155672
R1035 VTAIL.n226 VTAIL.n197 0.155672
R1036 VTAIL.n233 VTAIL.n197 0.155672
R1037 VTAIL.n234 VTAIL.n233 0.155672
R1038 VTAIL.n234 VTAIL.n193 0.155672
R1039 VTAIL.n241 VTAIL.n193 0.155672
R1040 VTAIL.n242 VTAIL.n241 0.155672
R1041 VTAIL.n242 VTAIL.n189 0.155672
R1042 VTAIL.n249 VTAIL.n189 0.155672
R1043 VTAIL.n250 VTAIL.n249 0.155672
R1044 VTAIL.n250 VTAIL.n185 0.155672
R1045 VTAIL.n259 VTAIL.n185 0.155672
R1046 VTAIL.n260 VTAIL.n259 0.155672
R1047 VTAIL.n260 VTAIL.n181 0.155672
R1048 VTAIL.n267 VTAIL.n181 0.155672
R1049 VTAIL.n627 VTAIL.n541 0.155672
R1050 VTAIL.n620 VTAIL.n541 0.155672
R1051 VTAIL.n620 VTAIL.n619 0.155672
R1052 VTAIL.n619 VTAIL.n545 0.155672
R1053 VTAIL.n611 VTAIL.n545 0.155672
R1054 VTAIL.n611 VTAIL.n610 0.155672
R1055 VTAIL.n610 VTAIL.n550 0.155672
R1056 VTAIL.n603 VTAIL.n550 0.155672
R1057 VTAIL.n603 VTAIL.n602 0.155672
R1058 VTAIL.n602 VTAIL.n554 0.155672
R1059 VTAIL.n595 VTAIL.n554 0.155672
R1060 VTAIL.n595 VTAIL.n594 0.155672
R1061 VTAIL.n594 VTAIL.n558 0.155672
R1062 VTAIL.n587 VTAIL.n558 0.155672
R1063 VTAIL.n587 VTAIL.n586 0.155672
R1064 VTAIL.n586 VTAIL.n562 0.155672
R1065 VTAIL.n579 VTAIL.n562 0.155672
R1066 VTAIL.n579 VTAIL.n578 0.155672
R1067 VTAIL.n578 VTAIL.n566 0.155672
R1068 VTAIL.n571 VTAIL.n566 0.155672
R1069 VTAIL.n537 VTAIL.n451 0.155672
R1070 VTAIL.n530 VTAIL.n451 0.155672
R1071 VTAIL.n530 VTAIL.n529 0.155672
R1072 VTAIL.n529 VTAIL.n455 0.155672
R1073 VTAIL.n521 VTAIL.n455 0.155672
R1074 VTAIL.n521 VTAIL.n520 0.155672
R1075 VTAIL.n520 VTAIL.n460 0.155672
R1076 VTAIL.n513 VTAIL.n460 0.155672
R1077 VTAIL.n513 VTAIL.n512 0.155672
R1078 VTAIL.n512 VTAIL.n464 0.155672
R1079 VTAIL.n505 VTAIL.n464 0.155672
R1080 VTAIL.n505 VTAIL.n504 0.155672
R1081 VTAIL.n504 VTAIL.n468 0.155672
R1082 VTAIL.n497 VTAIL.n468 0.155672
R1083 VTAIL.n497 VTAIL.n496 0.155672
R1084 VTAIL.n496 VTAIL.n472 0.155672
R1085 VTAIL.n489 VTAIL.n472 0.155672
R1086 VTAIL.n489 VTAIL.n488 0.155672
R1087 VTAIL.n488 VTAIL.n476 0.155672
R1088 VTAIL.n481 VTAIL.n476 0.155672
R1089 VTAIL.n447 VTAIL.n361 0.155672
R1090 VTAIL.n440 VTAIL.n361 0.155672
R1091 VTAIL.n440 VTAIL.n439 0.155672
R1092 VTAIL.n439 VTAIL.n365 0.155672
R1093 VTAIL.n431 VTAIL.n365 0.155672
R1094 VTAIL.n431 VTAIL.n430 0.155672
R1095 VTAIL.n430 VTAIL.n370 0.155672
R1096 VTAIL.n423 VTAIL.n370 0.155672
R1097 VTAIL.n423 VTAIL.n422 0.155672
R1098 VTAIL.n422 VTAIL.n374 0.155672
R1099 VTAIL.n415 VTAIL.n374 0.155672
R1100 VTAIL.n415 VTAIL.n414 0.155672
R1101 VTAIL.n414 VTAIL.n378 0.155672
R1102 VTAIL.n407 VTAIL.n378 0.155672
R1103 VTAIL.n407 VTAIL.n406 0.155672
R1104 VTAIL.n406 VTAIL.n382 0.155672
R1105 VTAIL.n399 VTAIL.n382 0.155672
R1106 VTAIL.n399 VTAIL.n398 0.155672
R1107 VTAIL.n398 VTAIL.n386 0.155672
R1108 VTAIL.n391 VTAIL.n386 0.155672
R1109 VTAIL.n357 VTAIL.n271 0.155672
R1110 VTAIL.n350 VTAIL.n271 0.155672
R1111 VTAIL.n350 VTAIL.n349 0.155672
R1112 VTAIL.n349 VTAIL.n275 0.155672
R1113 VTAIL.n341 VTAIL.n275 0.155672
R1114 VTAIL.n341 VTAIL.n340 0.155672
R1115 VTAIL.n340 VTAIL.n280 0.155672
R1116 VTAIL.n333 VTAIL.n280 0.155672
R1117 VTAIL.n333 VTAIL.n332 0.155672
R1118 VTAIL.n332 VTAIL.n284 0.155672
R1119 VTAIL.n325 VTAIL.n284 0.155672
R1120 VTAIL.n325 VTAIL.n324 0.155672
R1121 VTAIL.n324 VTAIL.n288 0.155672
R1122 VTAIL.n317 VTAIL.n288 0.155672
R1123 VTAIL.n317 VTAIL.n316 0.155672
R1124 VTAIL.n316 VTAIL.n292 0.155672
R1125 VTAIL.n309 VTAIL.n292 0.155672
R1126 VTAIL.n309 VTAIL.n308 0.155672
R1127 VTAIL.n308 VTAIL.n296 0.155672
R1128 VTAIL.n301 VTAIL.n296 0.155672
R1129 VN.n1 VN.t1 143.006
R1130 VN.n0 VN.t3 143.006
R1131 VN.n0 VN.t0 141.76
R1132 VN.n1 VN.t2 141.76
R1133 VN VN.n1 54.926
R1134 VN VN.n0 2.08127
R1135 VDD2.n2 VDD2.n0 119.594
R1136 VDD2.n2 VDD2.n1 71.7413
R1137 VDD2.n1 VDD2.t1 2.00946
R1138 VDD2.n1 VDD2.t2 2.00946
R1139 VDD2.n0 VDD2.t0 2.00946
R1140 VDD2.n0 VDD2.t3 2.00946
R1141 VDD2 VDD2.n2 0.0586897
R1142 B.n586 B.n585 585
R1143 B.n587 B.n86 585
R1144 B.n589 B.n588 585
R1145 B.n590 B.n85 585
R1146 B.n592 B.n591 585
R1147 B.n593 B.n84 585
R1148 B.n595 B.n594 585
R1149 B.n596 B.n83 585
R1150 B.n598 B.n597 585
R1151 B.n599 B.n82 585
R1152 B.n601 B.n600 585
R1153 B.n602 B.n81 585
R1154 B.n604 B.n603 585
R1155 B.n605 B.n80 585
R1156 B.n607 B.n606 585
R1157 B.n608 B.n79 585
R1158 B.n610 B.n609 585
R1159 B.n611 B.n78 585
R1160 B.n613 B.n612 585
R1161 B.n614 B.n77 585
R1162 B.n616 B.n615 585
R1163 B.n617 B.n76 585
R1164 B.n619 B.n618 585
R1165 B.n620 B.n75 585
R1166 B.n622 B.n621 585
R1167 B.n623 B.n74 585
R1168 B.n625 B.n624 585
R1169 B.n626 B.n73 585
R1170 B.n628 B.n627 585
R1171 B.n629 B.n72 585
R1172 B.n631 B.n630 585
R1173 B.n632 B.n71 585
R1174 B.n634 B.n633 585
R1175 B.n635 B.n70 585
R1176 B.n637 B.n636 585
R1177 B.n638 B.n69 585
R1178 B.n640 B.n639 585
R1179 B.n641 B.n68 585
R1180 B.n643 B.n642 585
R1181 B.n644 B.n67 585
R1182 B.n646 B.n645 585
R1183 B.n647 B.n66 585
R1184 B.n649 B.n648 585
R1185 B.n650 B.n65 585
R1186 B.n652 B.n651 585
R1187 B.n653 B.n64 585
R1188 B.n655 B.n654 585
R1189 B.n656 B.n63 585
R1190 B.n658 B.n657 585
R1191 B.n659 B.n62 585
R1192 B.n661 B.n660 585
R1193 B.n662 B.n61 585
R1194 B.n664 B.n663 585
R1195 B.n665 B.n58 585
R1196 B.n668 B.n667 585
R1197 B.n669 B.n57 585
R1198 B.n671 B.n670 585
R1199 B.n672 B.n56 585
R1200 B.n674 B.n673 585
R1201 B.n675 B.n55 585
R1202 B.n677 B.n676 585
R1203 B.n678 B.n51 585
R1204 B.n680 B.n679 585
R1205 B.n681 B.n50 585
R1206 B.n683 B.n682 585
R1207 B.n684 B.n49 585
R1208 B.n686 B.n685 585
R1209 B.n687 B.n48 585
R1210 B.n689 B.n688 585
R1211 B.n690 B.n47 585
R1212 B.n692 B.n691 585
R1213 B.n693 B.n46 585
R1214 B.n695 B.n694 585
R1215 B.n696 B.n45 585
R1216 B.n698 B.n697 585
R1217 B.n699 B.n44 585
R1218 B.n701 B.n700 585
R1219 B.n702 B.n43 585
R1220 B.n704 B.n703 585
R1221 B.n705 B.n42 585
R1222 B.n707 B.n706 585
R1223 B.n708 B.n41 585
R1224 B.n710 B.n709 585
R1225 B.n711 B.n40 585
R1226 B.n713 B.n712 585
R1227 B.n714 B.n39 585
R1228 B.n716 B.n715 585
R1229 B.n717 B.n38 585
R1230 B.n719 B.n718 585
R1231 B.n720 B.n37 585
R1232 B.n722 B.n721 585
R1233 B.n723 B.n36 585
R1234 B.n725 B.n724 585
R1235 B.n726 B.n35 585
R1236 B.n728 B.n727 585
R1237 B.n729 B.n34 585
R1238 B.n731 B.n730 585
R1239 B.n732 B.n33 585
R1240 B.n734 B.n733 585
R1241 B.n735 B.n32 585
R1242 B.n737 B.n736 585
R1243 B.n738 B.n31 585
R1244 B.n740 B.n739 585
R1245 B.n741 B.n30 585
R1246 B.n743 B.n742 585
R1247 B.n744 B.n29 585
R1248 B.n746 B.n745 585
R1249 B.n747 B.n28 585
R1250 B.n749 B.n748 585
R1251 B.n750 B.n27 585
R1252 B.n752 B.n751 585
R1253 B.n753 B.n26 585
R1254 B.n755 B.n754 585
R1255 B.n756 B.n25 585
R1256 B.n758 B.n757 585
R1257 B.n759 B.n24 585
R1258 B.n761 B.n760 585
R1259 B.n584 B.n87 585
R1260 B.n583 B.n582 585
R1261 B.n581 B.n88 585
R1262 B.n580 B.n579 585
R1263 B.n578 B.n89 585
R1264 B.n577 B.n576 585
R1265 B.n575 B.n90 585
R1266 B.n574 B.n573 585
R1267 B.n572 B.n91 585
R1268 B.n571 B.n570 585
R1269 B.n569 B.n92 585
R1270 B.n568 B.n567 585
R1271 B.n566 B.n93 585
R1272 B.n565 B.n564 585
R1273 B.n563 B.n94 585
R1274 B.n562 B.n561 585
R1275 B.n560 B.n95 585
R1276 B.n559 B.n558 585
R1277 B.n557 B.n96 585
R1278 B.n556 B.n555 585
R1279 B.n554 B.n97 585
R1280 B.n553 B.n552 585
R1281 B.n551 B.n98 585
R1282 B.n550 B.n549 585
R1283 B.n548 B.n99 585
R1284 B.n547 B.n546 585
R1285 B.n545 B.n100 585
R1286 B.n544 B.n543 585
R1287 B.n542 B.n101 585
R1288 B.n541 B.n540 585
R1289 B.n539 B.n102 585
R1290 B.n538 B.n537 585
R1291 B.n536 B.n103 585
R1292 B.n535 B.n534 585
R1293 B.n533 B.n104 585
R1294 B.n532 B.n531 585
R1295 B.n530 B.n105 585
R1296 B.n529 B.n528 585
R1297 B.n527 B.n106 585
R1298 B.n526 B.n525 585
R1299 B.n524 B.n107 585
R1300 B.n523 B.n522 585
R1301 B.n521 B.n108 585
R1302 B.n520 B.n519 585
R1303 B.n518 B.n109 585
R1304 B.n517 B.n516 585
R1305 B.n515 B.n110 585
R1306 B.n514 B.n513 585
R1307 B.n512 B.n111 585
R1308 B.n511 B.n510 585
R1309 B.n509 B.n112 585
R1310 B.n508 B.n507 585
R1311 B.n506 B.n113 585
R1312 B.n505 B.n504 585
R1313 B.n503 B.n114 585
R1314 B.n502 B.n501 585
R1315 B.n500 B.n115 585
R1316 B.n499 B.n498 585
R1317 B.n497 B.n116 585
R1318 B.n496 B.n495 585
R1319 B.n494 B.n117 585
R1320 B.n493 B.n492 585
R1321 B.n491 B.n118 585
R1322 B.n490 B.n489 585
R1323 B.n488 B.n119 585
R1324 B.n487 B.n486 585
R1325 B.n485 B.n120 585
R1326 B.n484 B.n483 585
R1327 B.n482 B.n121 585
R1328 B.n481 B.n480 585
R1329 B.n479 B.n122 585
R1330 B.n478 B.n477 585
R1331 B.n476 B.n123 585
R1332 B.n475 B.n474 585
R1333 B.n473 B.n124 585
R1334 B.n472 B.n471 585
R1335 B.n470 B.n125 585
R1336 B.n469 B.n468 585
R1337 B.n467 B.n126 585
R1338 B.n466 B.n465 585
R1339 B.n464 B.n127 585
R1340 B.n463 B.n462 585
R1341 B.n461 B.n128 585
R1342 B.n460 B.n459 585
R1343 B.n458 B.n129 585
R1344 B.n457 B.n456 585
R1345 B.n455 B.n130 585
R1346 B.n276 B.n275 585
R1347 B.n277 B.n190 585
R1348 B.n279 B.n278 585
R1349 B.n280 B.n189 585
R1350 B.n282 B.n281 585
R1351 B.n283 B.n188 585
R1352 B.n285 B.n284 585
R1353 B.n286 B.n187 585
R1354 B.n288 B.n287 585
R1355 B.n289 B.n186 585
R1356 B.n291 B.n290 585
R1357 B.n292 B.n185 585
R1358 B.n294 B.n293 585
R1359 B.n295 B.n184 585
R1360 B.n297 B.n296 585
R1361 B.n298 B.n183 585
R1362 B.n300 B.n299 585
R1363 B.n301 B.n182 585
R1364 B.n303 B.n302 585
R1365 B.n304 B.n181 585
R1366 B.n306 B.n305 585
R1367 B.n307 B.n180 585
R1368 B.n309 B.n308 585
R1369 B.n310 B.n179 585
R1370 B.n312 B.n311 585
R1371 B.n313 B.n178 585
R1372 B.n315 B.n314 585
R1373 B.n316 B.n177 585
R1374 B.n318 B.n317 585
R1375 B.n319 B.n176 585
R1376 B.n321 B.n320 585
R1377 B.n322 B.n175 585
R1378 B.n324 B.n323 585
R1379 B.n325 B.n174 585
R1380 B.n327 B.n326 585
R1381 B.n328 B.n173 585
R1382 B.n330 B.n329 585
R1383 B.n331 B.n172 585
R1384 B.n333 B.n332 585
R1385 B.n334 B.n171 585
R1386 B.n336 B.n335 585
R1387 B.n337 B.n170 585
R1388 B.n339 B.n338 585
R1389 B.n340 B.n169 585
R1390 B.n342 B.n341 585
R1391 B.n343 B.n168 585
R1392 B.n345 B.n344 585
R1393 B.n346 B.n167 585
R1394 B.n348 B.n347 585
R1395 B.n349 B.n166 585
R1396 B.n351 B.n350 585
R1397 B.n352 B.n165 585
R1398 B.n354 B.n353 585
R1399 B.n355 B.n162 585
R1400 B.n358 B.n357 585
R1401 B.n359 B.n161 585
R1402 B.n361 B.n360 585
R1403 B.n362 B.n160 585
R1404 B.n364 B.n363 585
R1405 B.n365 B.n159 585
R1406 B.n367 B.n366 585
R1407 B.n368 B.n158 585
R1408 B.n373 B.n372 585
R1409 B.n374 B.n157 585
R1410 B.n376 B.n375 585
R1411 B.n377 B.n156 585
R1412 B.n379 B.n378 585
R1413 B.n380 B.n155 585
R1414 B.n382 B.n381 585
R1415 B.n383 B.n154 585
R1416 B.n385 B.n384 585
R1417 B.n386 B.n153 585
R1418 B.n388 B.n387 585
R1419 B.n389 B.n152 585
R1420 B.n391 B.n390 585
R1421 B.n392 B.n151 585
R1422 B.n394 B.n393 585
R1423 B.n395 B.n150 585
R1424 B.n397 B.n396 585
R1425 B.n398 B.n149 585
R1426 B.n400 B.n399 585
R1427 B.n401 B.n148 585
R1428 B.n403 B.n402 585
R1429 B.n404 B.n147 585
R1430 B.n406 B.n405 585
R1431 B.n407 B.n146 585
R1432 B.n409 B.n408 585
R1433 B.n410 B.n145 585
R1434 B.n412 B.n411 585
R1435 B.n413 B.n144 585
R1436 B.n415 B.n414 585
R1437 B.n416 B.n143 585
R1438 B.n418 B.n417 585
R1439 B.n419 B.n142 585
R1440 B.n421 B.n420 585
R1441 B.n422 B.n141 585
R1442 B.n424 B.n423 585
R1443 B.n425 B.n140 585
R1444 B.n427 B.n426 585
R1445 B.n428 B.n139 585
R1446 B.n430 B.n429 585
R1447 B.n431 B.n138 585
R1448 B.n433 B.n432 585
R1449 B.n434 B.n137 585
R1450 B.n436 B.n435 585
R1451 B.n437 B.n136 585
R1452 B.n439 B.n438 585
R1453 B.n440 B.n135 585
R1454 B.n442 B.n441 585
R1455 B.n443 B.n134 585
R1456 B.n445 B.n444 585
R1457 B.n446 B.n133 585
R1458 B.n448 B.n447 585
R1459 B.n449 B.n132 585
R1460 B.n451 B.n450 585
R1461 B.n452 B.n131 585
R1462 B.n454 B.n453 585
R1463 B.n274 B.n191 585
R1464 B.n273 B.n272 585
R1465 B.n271 B.n192 585
R1466 B.n270 B.n269 585
R1467 B.n268 B.n193 585
R1468 B.n267 B.n266 585
R1469 B.n265 B.n194 585
R1470 B.n264 B.n263 585
R1471 B.n262 B.n195 585
R1472 B.n261 B.n260 585
R1473 B.n259 B.n196 585
R1474 B.n258 B.n257 585
R1475 B.n256 B.n197 585
R1476 B.n255 B.n254 585
R1477 B.n253 B.n198 585
R1478 B.n252 B.n251 585
R1479 B.n250 B.n199 585
R1480 B.n249 B.n248 585
R1481 B.n247 B.n200 585
R1482 B.n246 B.n245 585
R1483 B.n244 B.n201 585
R1484 B.n243 B.n242 585
R1485 B.n241 B.n202 585
R1486 B.n240 B.n239 585
R1487 B.n238 B.n203 585
R1488 B.n237 B.n236 585
R1489 B.n235 B.n204 585
R1490 B.n234 B.n233 585
R1491 B.n232 B.n205 585
R1492 B.n231 B.n230 585
R1493 B.n229 B.n206 585
R1494 B.n228 B.n227 585
R1495 B.n226 B.n207 585
R1496 B.n225 B.n224 585
R1497 B.n223 B.n208 585
R1498 B.n222 B.n221 585
R1499 B.n220 B.n209 585
R1500 B.n219 B.n218 585
R1501 B.n217 B.n210 585
R1502 B.n216 B.n215 585
R1503 B.n214 B.n211 585
R1504 B.n213 B.n212 585
R1505 B.n2 B.n0 585
R1506 B.n825 B.n1 585
R1507 B.n824 B.n823 585
R1508 B.n822 B.n3 585
R1509 B.n821 B.n820 585
R1510 B.n819 B.n4 585
R1511 B.n818 B.n817 585
R1512 B.n816 B.n5 585
R1513 B.n815 B.n814 585
R1514 B.n813 B.n6 585
R1515 B.n812 B.n811 585
R1516 B.n810 B.n7 585
R1517 B.n809 B.n808 585
R1518 B.n807 B.n8 585
R1519 B.n806 B.n805 585
R1520 B.n804 B.n9 585
R1521 B.n803 B.n802 585
R1522 B.n801 B.n10 585
R1523 B.n800 B.n799 585
R1524 B.n798 B.n11 585
R1525 B.n797 B.n796 585
R1526 B.n795 B.n12 585
R1527 B.n794 B.n793 585
R1528 B.n792 B.n13 585
R1529 B.n791 B.n790 585
R1530 B.n789 B.n14 585
R1531 B.n788 B.n787 585
R1532 B.n786 B.n15 585
R1533 B.n785 B.n784 585
R1534 B.n783 B.n16 585
R1535 B.n782 B.n781 585
R1536 B.n780 B.n17 585
R1537 B.n779 B.n778 585
R1538 B.n777 B.n18 585
R1539 B.n776 B.n775 585
R1540 B.n774 B.n19 585
R1541 B.n773 B.n772 585
R1542 B.n771 B.n20 585
R1543 B.n770 B.n769 585
R1544 B.n768 B.n21 585
R1545 B.n767 B.n766 585
R1546 B.n765 B.n22 585
R1547 B.n764 B.n763 585
R1548 B.n762 B.n23 585
R1549 B.n827 B.n826 585
R1550 B.n369 B.t2 527.369
R1551 B.n59 B.t7 527.369
R1552 B.n163 B.t11 527.369
R1553 B.n52 B.t4 527.369
R1554 B.n275 B.n274 511.721
R1555 B.n760 B.n23 511.721
R1556 B.n453 B.n130 511.721
R1557 B.n585 B.n584 511.721
R1558 B.n370 B.t1 450.957
R1559 B.n60 B.t8 450.957
R1560 B.n164 B.t10 450.955
R1561 B.n53 B.t5 450.955
R1562 B.n369 B.t0 317.207
R1563 B.n163 B.t9 317.207
R1564 B.n52 B.t3 317.207
R1565 B.n59 B.t6 317.207
R1566 B.n274 B.n273 163.367
R1567 B.n273 B.n192 163.367
R1568 B.n269 B.n192 163.367
R1569 B.n269 B.n268 163.367
R1570 B.n268 B.n267 163.367
R1571 B.n267 B.n194 163.367
R1572 B.n263 B.n194 163.367
R1573 B.n263 B.n262 163.367
R1574 B.n262 B.n261 163.367
R1575 B.n261 B.n196 163.367
R1576 B.n257 B.n196 163.367
R1577 B.n257 B.n256 163.367
R1578 B.n256 B.n255 163.367
R1579 B.n255 B.n198 163.367
R1580 B.n251 B.n198 163.367
R1581 B.n251 B.n250 163.367
R1582 B.n250 B.n249 163.367
R1583 B.n249 B.n200 163.367
R1584 B.n245 B.n200 163.367
R1585 B.n245 B.n244 163.367
R1586 B.n244 B.n243 163.367
R1587 B.n243 B.n202 163.367
R1588 B.n239 B.n202 163.367
R1589 B.n239 B.n238 163.367
R1590 B.n238 B.n237 163.367
R1591 B.n237 B.n204 163.367
R1592 B.n233 B.n204 163.367
R1593 B.n233 B.n232 163.367
R1594 B.n232 B.n231 163.367
R1595 B.n231 B.n206 163.367
R1596 B.n227 B.n206 163.367
R1597 B.n227 B.n226 163.367
R1598 B.n226 B.n225 163.367
R1599 B.n225 B.n208 163.367
R1600 B.n221 B.n208 163.367
R1601 B.n221 B.n220 163.367
R1602 B.n220 B.n219 163.367
R1603 B.n219 B.n210 163.367
R1604 B.n215 B.n210 163.367
R1605 B.n215 B.n214 163.367
R1606 B.n214 B.n213 163.367
R1607 B.n213 B.n2 163.367
R1608 B.n826 B.n2 163.367
R1609 B.n826 B.n825 163.367
R1610 B.n825 B.n824 163.367
R1611 B.n824 B.n3 163.367
R1612 B.n820 B.n3 163.367
R1613 B.n820 B.n819 163.367
R1614 B.n819 B.n818 163.367
R1615 B.n818 B.n5 163.367
R1616 B.n814 B.n5 163.367
R1617 B.n814 B.n813 163.367
R1618 B.n813 B.n812 163.367
R1619 B.n812 B.n7 163.367
R1620 B.n808 B.n7 163.367
R1621 B.n808 B.n807 163.367
R1622 B.n807 B.n806 163.367
R1623 B.n806 B.n9 163.367
R1624 B.n802 B.n9 163.367
R1625 B.n802 B.n801 163.367
R1626 B.n801 B.n800 163.367
R1627 B.n800 B.n11 163.367
R1628 B.n796 B.n11 163.367
R1629 B.n796 B.n795 163.367
R1630 B.n795 B.n794 163.367
R1631 B.n794 B.n13 163.367
R1632 B.n790 B.n13 163.367
R1633 B.n790 B.n789 163.367
R1634 B.n789 B.n788 163.367
R1635 B.n788 B.n15 163.367
R1636 B.n784 B.n15 163.367
R1637 B.n784 B.n783 163.367
R1638 B.n783 B.n782 163.367
R1639 B.n782 B.n17 163.367
R1640 B.n778 B.n17 163.367
R1641 B.n778 B.n777 163.367
R1642 B.n777 B.n776 163.367
R1643 B.n776 B.n19 163.367
R1644 B.n772 B.n19 163.367
R1645 B.n772 B.n771 163.367
R1646 B.n771 B.n770 163.367
R1647 B.n770 B.n21 163.367
R1648 B.n766 B.n21 163.367
R1649 B.n766 B.n765 163.367
R1650 B.n765 B.n764 163.367
R1651 B.n764 B.n23 163.367
R1652 B.n275 B.n190 163.367
R1653 B.n279 B.n190 163.367
R1654 B.n280 B.n279 163.367
R1655 B.n281 B.n280 163.367
R1656 B.n281 B.n188 163.367
R1657 B.n285 B.n188 163.367
R1658 B.n286 B.n285 163.367
R1659 B.n287 B.n286 163.367
R1660 B.n287 B.n186 163.367
R1661 B.n291 B.n186 163.367
R1662 B.n292 B.n291 163.367
R1663 B.n293 B.n292 163.367
R1664 B.n293 B.n184 163.367
R1665 B.n297 B.n184 163.367
R1666 B.n298 B.n297 163.367
R1667 B.n299 B.n298 163.367
R1668 B.n299 B.n182 163.367
R1669 B.n303 B.n182 163.367
R1670 B.n304 B.n303 163.367
R1671 B.n305 B.n304 163.367
R1672 B.n305 B.n180 163.367
R1673 B.n309 B.n180 163.367
R1674 B.n310 B.n309 163.367
R1675 B.n311 B.n310 163.367
R1676 B.n311 B.n178 163.367
R1677 B.n315 B.n178 163.367
R1678 B.n316 B.n315 163.367
R1679 B.n317 B.n316 163.367
R1680 B.n317 B.n176 163.367
R1681 B.n321 B.n176 163.367
R1682 B.n322 B.n321 163.367
R1683 B.n323 B.n322 163.367
R1684 B.n323 B.n174 163.367
R1685 B.n327 B.n174 163.367
R1686 B.n328 B.n327 163.367
R1687 B.n329 B.n328 163.367
R1688 B.n329 B.n172 163.367
R1689 B.n333 B.n172 163.367
R1690 B.n334 B.n333 163.367
R1691 B.n335 B.n334 163.367
R1692 B.n335 B.n170 163.367
R1693 B.n339 B.n170 163.367
R1694 B.n340 B.n339 163.367
R1695 B.n341 B.n340 163.367
R1696 B.n341 B.n168 163.367
R1697 B.n345 B.n168 163.367
R1698 B.n346 B.n345 163.367
R1699 B.n347 B.n346 163.367
R1700 B.n347 B.n166 163.367
R1701 B.n351 B.n166 163.367
R1702 B.n352 B.n351 163.367
R1703 B.n353 B.n352 163.367
R1704 B.n353 B.n162 163.367
R1705 B.n358 B.n162 163.367
R1706 B.n359 B.n358 163.367
R1707 B.n360 B.n359 163.367
R1708 B.n360 B.n160 163.367
R1709 B.n364 B.n160 163.367
R1710 B.n365 B.n364 163.367
R1711 B.n366 B.n365 163.367
R1712 B.n366 B.n158 163.367
R1713 B.n373 B.n158 163.367
R1714 B.n374 B.n373 163.367
R1715 B.n375 B.n374 163.367
R1716 B.n375 B.n156 163.367
R1717 B.n379 B.n156 163.367
R1718 B.n380 B.n379 163.367
R1719 B.n381 B.n380 163.367
R1720 B.n381 B.n154 163.367
R1721 B.n385 B.n154 163.367
R1722 B.n386 B.n385 163.367
R1723 B.n387 B.n386 163.367
R1724 B.n387 B.n152 163.367
R1725 B.n391 B.n152 163.367
R1726 B.n392 B.n391 163.367
R1727 B.n393 B.n392 163.367
R1728 B.n393 B.n150 163.367
R1729 B.n397 B.n150 163.367
R1730 B.n398 B.n397 163.367
R1731 B.n399 B.n398 163.367
R1732 B.n399 B.n148 163.367
R1733 B.n403 B.n148 163.367
R1734 B.n404 B.n403 163.367
R1735 B.n405 B.n404 163.367
R1736 B.n405 B.n146 163.367
R1737 B.n409 B.n146 163.367
R1738 B.n410 B.n409 163.367
R1739 B.n411 B.n410 163.367
R1740 B.n411 B.n144 163.367
R1741 B.n415 B.n144 163.367
R1742 B.n416 B.n415 163.367
R1743 B.n417 B.n416 163.367
R1744 B.n417 B.n142 163.367
R1745 B.n421 B.n142 163.367
R1746 B.n422 B.n421 163.367
R1747 B.n423 B.n422 163.367
R1748 B.n423 B.n140 163.367
R1749 B.n427 B.n140 163.367
R1750 B.n428 B.n427 163.367
R1751 B.n429 B.n428 163.367
R1752 B.n429 B.n138 163.367
R1753 B.n433 B.n138 163.367
R1754 B.n434 B.n433 163.367
R1755 B.n435 B.n434 163.367
R1756 B.n435 B.n136 163.367
R1757 B.n439 B.n136 163.367
R1758 B.n440 B.n439 163.367
R1759 B.n441 B.n440 163.367
R1760 B.n441 B.n134 163.367
R1761 B.n445 B.n134 163.367
R1762 B.n446 B.n445 163.367
R1763 B.n447 B.n446 163.367
R1764 B.n447 B.n132 163.367
R1765 B.n451 B.n132 163.367
R1766 B.n452 B.n451 163.367
R1767 B.n453 B.n452 163.367
R1768 B.n457 B.n130 163.367
R1769 B.n458 B.n457 163.367
R1770 B.n459 B.n458 163.367
R1771 B.n459 B.n128 163.367
R1772 B.n463 B.n128 163.367
R1773 B.n464 B.n463 163.367
R1774 B.n465 B.n464 163.367
R1775 B.n465 B.n126 163.367
R1776 B.n469 B.n126 163.367
R1777 B.n470 B.n469 163.367
R1778 B.n471 B.n470 163.367
R1779 B.n471 B.n124 163.367
R1780 B.n475 B.n124 163.367
R1781 B.n476 B.n475 163.367
R1782 B.n477 B.n476 163.367
R1783 B.n477 B.n122 163.367
R1784 B.n481 B.n122 163.367
R1785 B.n482 B.n481 163.367
R1786 B.n483 B.n482 163.367
R1787 B.n483 B.n120 163.367
R1788 B.n487 B.n120 163.367
R1789 B.n488 B.n487 163.367
R1790 B.n489 B.n488 163.367
R1791 B.n489 B.n118 163.367
R1792 B.n493 B.n118 163.367
R1793 B.n494 B.n493 163.367
R1794 B.n495 B.n494 163.367
R1795 B.n495 B.n116 163.367
R1796 B.n499 B.n116 163.367
R1797 B.n500 B.n499 163.367
R1798 B.n501 B.n500 163.367
R1799 B.n501 B.n114 163.367
R1800 B.n505 B.n114 163.367
R1801 B.n506 B.n505 163.367
R1802 B.n507 B.n506 163.367
R1803 B.n507 B.n112 163.367
R1804 B.n511 B.n112 163.367
R1805 B.n512 B.n511 163.367
R1806 B.n513 B.n512 163.367
R1807 B.n513 B.n110 163.367
R1808 B.n517 B.n110 163.367
R1809 B.n518 B.n517 163.367
R1810 B.n519 B.n518 163.367
R1811 B.n519 B.n108 163.367
R1812 B.n523 B.n108 163.367
R1813 B.n524 B.n523 163.367
R1814 B.n525 B.n524 163.367
R1815 B.n525 B.n106 163.367
R1816 B.n529 B.n106 163.367
R1817 B.n530 B.n529 163.367
R1818 B.n531 B.n530 163.367
R1819 B.n531 B.n104 163.367
R1820 B.n535 B.n104 163.367
R1821 B.n536 B.n535 163.367
R1822 B.n537 B.n536 163.367
R1823 B.n537 B.n102 163.367
R1824 B.n541 B.n102 163.367
R1825 B.n542 B.n541 163.367
R1826 B.n543 B.n542 163.367
R1827 B.n543 B.n100 163.367
R1828 B.n547 B.n100 163.367
R1829 B.n548 B.n547 163.367
R1830 B.n549 B.n548 163.367
R1831 B.n549 B.n98 163.367
R1832 B.n553 B.n98 163.367
R1833 B.n554 B.n553 163.367
R1834 B.n555 B.n554 163.367
R1835 B.n555 B.n96 163.367
R1836 B.n559 B.n96 163.367
R1837 B.n560 B.n559 163.367
R1838 B.n561 B.n560 163.367
R1839 B.n561 B.n94 163.367
R1840 B.n565 B.n94 163.367
R1841 B.n566 B.n565 163.367
R1842 B.n567 B.n566 163.367
R1843 B.n567 B.n92 163.367
R1844 B.n571 B.n92 163.367
R1845 B.n572 B.n571 163.367
R1846 B.n573 B.n572 163.367
R1847 B.n573 B.n90 163.367
R1848 B.n577 B.n90 163.367
R1849 B.n578 B.n577 163.367
R1850 B.n579 B.n578 163.367
R1851 B.n579 B.n88 163.367
R1852 B.n583 B.n88 163.367
R1853 B.n584 B.n583 163.367
R1854 B.n760 B.n759 163.367
R1855 B.n759 B.n758 163.367
R1856 B.n758 B.n25 163.367
R1857 B.n754 B.n25 163.367
R1858 B.n754 B.n753 163.367
R1859 B.n753 B.n752 163.367
R1860 B.n752 B.n27 163.367
R1861 B.n748 B.n27 163.367
R1862 B.n748 B.n747 163.367
R1863 B.n747 B.n746 163.367
R1864 B.n746 B.n29 163.367
R1865 B.n742 B.n29 163.367
R1866 B.n742 B.n741 163.367
R1867 B.n741 B.n740 163.367
R1868 B.n740 B.n31 163.367
R1869 B.n736 B.n31 163.367
R1870 B.n736 B.n735 163.367
R1871 B.n735 B.n734 163.367
R1872 B.n734 B.n33 163.367
R1873 B.n730 B.n33 163.367
R1874 B.n730 B.n729 163.367
R1875 B.n729 B.n728 163.367
R1876 B.n728 B.n35 163.367
R1877 B.n724 B.n35 163.367
R1878 B.n724 B.n723 163.367
R1879 B.n723 B.n722 163.367
R1880 B.n722 B.n37 163.367
R1881 B.n718 B.n37 163.367
R1882 B.n718 B.n717 163.367
R1883 B.n717 B.n716 163.367
R1884 B.n716 B.n39 163.367
R1885 B.n712 B.n39 163.367
R1886 B.n712 B.n711 163.367
R1887 B.n711 B.n710 163.367
R1888 B.n710 B.n41 163.367
R1889 B.n706 B.n41 163.367
R1890 B.n706 B.n705 163.367
R1891 B.n705 B.n704 163.367
R1892 B.n704 B.n43 163.367
R1893 B.n700 B.n43 163.367
R1894 B.n700 B.n699 163.367
R1895 B.n699 B.n698 163.367
R1896 B.n698 B.n45 163.367
R1897 B.n694 B.n45 163.367
R1898 B.n694 B.n693 163.367
R1899 B.n693 B.n692 163.367
R1900 B.n692 B.n47 163.367
R1901 B.n688 B.n47 163.367
R1902 B.n688 B.n687 163.367
R1903 B.n687 B.n686 163.367
R1904 B.n686 B.n49 163.367
R1905 B.n682 B.n49 163.367
R1906 B.n682 B.n681 163.367
R1907 B.n681 B.n680 163.367
R1908 B.n680 B.n51 163.367
R1909 B.n676 B.n51 163.367
R1910 B.n676 B.n675 163.367
R1911 B.n675 B.n674 163.367
R1912 B.n674 B.n56 163.367
R1913 B.n670 B.n56 163.367
R1914 B.n670 B.n669 163.367
R1915 B.n669 B.n668 163.367
R1916 B.n668 B.n58 163.367
R1917 B.n663 B.n58 163.367
R1918 B.n663 B.n662 163.367
R1919 B.n662 B.n661 163.367
R1920 B.n661 B.n62 163.367
R1921 B.n657 B.n62 163.367
R1922 B.n657 B.n656 163.367
R1923 B.n656 B.n655 163.367
R1924 B.n655 B.n64 163.367
R1925 B.n651 B.n64 163.367
R1926 B.n651 B.n650 163.367
R1927 B.n650 B.n649 163.367
R1928 B.n649 B.n66 163.367
R1929 B.n645 B.n66 163.367
R1930 B.n645 B.n644 163.367
R1931 B.n644 B.n643 163.367
R1932 B.n643 B.n68 163.367
R1933 B.n639 B.n68 163.367
R1934 B.n639 B.n638 163.367
R1935 B.n638 B.n637 163.367
R1936 B.n637 B.n70 163.367
R1937 B.n633 B.n70 163.367
R1938 B.n633 B.n632 163.367
R1939 B.n632 B.n631 163.367
R1940 B.n631 B.n72 163.367
R1941 B.n627 B.n72 163.367
R1942 B.n627 B.n626 163.367
R1943 B.n626 B.n625 163.367
R1944 B.n625 B.n74 163.367
R1945 B.n621 B.n74 163.367
R1946 B.n621 B.n620 163.367
R1947 B.n620 B.n619 163.367
R1948 B.n619 B.n76 163.367
R1949 B.n615 B.n76 163.367
R1950 B.n615 B.n614 163.367
R1951 B.n614 B.n613 163.367
R1952 B.n613 B.n78 163.367
R1953 B.n609 B.n78 163.367
R1954 B.n609 B.n608 163.367
R1955 B.n608 B.n607 163.367
R1956 B.n607 B.n80 163.367
R1957 B.n603 B.n80 163.367
R1958 B.n603 B.n602 163.367
R1959 B.n602 B.n601 163.367
R1960 B.n601 B.n82 163.367
R1961 B.n597 B.n82 163.367
R1962 B.n597 B.n596 163.367
R1963 B.n596 B.n595 163.367
R1964 B.n595 B.n84 163.367
R1965 B.n591 B.n84 163.367
R1966 B.n591 B.n590 163.367
R1967 B.n590 B.n589 163.367
R1968 B.n589 B.n86 163.367
R1969 B.n585 B.n86 163.367
R1970 B.n370 B.n369 76.4126
R1971 B.n164 B.n163 76.4126
R1972 B.n53 B.n52 76.4126
R1973 B.n60 B.n59 76.4126
R1974 B.n371 B.n370 59.5399
R1975 B.n356 B.n164 59.5399
R1976 B.n54 B.n53 59.5399
R1977 B.n666 B.n60 59.5399
R1978 B.n762 B.n761 33.2493
R1979 B.n586 B.n87 33.2493
R1980 B.n455 B.n454 33.2493
R1981 B.n276 B.n191 33.2493
R1982 B B.n827 18.0485
R1983 B.n761 B.n24 10.6151
R1984 B.n757 B.n24 10.6151
R1985 B.n757 B.n756 10.6151
R1986 B.n756 B.n755 10.6151
R1987 B.n755 B.n26 10.6151
R1988 B.n751 B.n26 10.6151
R1989 B.n751 B.n750 10.6151
R1990 B.n750 B.n749 10.6151
R1991 B.n749 B.n28 10.6151
R1992 B.n745 B.n28 10.6151
R1993 B.n745 B.n744 10.6151
R1994 B.n744 B.n743 10.6151
R1995 B.n743 B.n30 10.6151
R1996 B.n739 B.n30 10.6151
R1997 B.n739 B.n738 10.6151
R1998 B.n738 B.n737 10.6151
R1999 B.n737 B.n32 10.6151
R2000 B.n733 B.n32 10.6151
R2001 B.n733 B.n732 10.6151
R2002 B.n732 B.n731 10.6151
R2003 B.n731 B.n34 10.6151
R2004 B.n727 B.n34 10.6151
R2005 B.n727 B.n726 10.6151
R2006 B.n726 B.n725 10.6151
R2007 B.n725 B.n36 10.6151
R2008 B.n721 B.n36 10.6151
R2009 B.n721 B.n720 10.6151
R2010 B.n720 B.n719 10.6151
R2011 B.n719 B.n38 10.6151
R2012 B.n715 B.n38 10.6151
R2013 B.n715 B.n714 10.6151
R2014 B.n714 B.n713 10.6151
R2015 B.n713 B.n40 10.6151
R2016 B.n709 B.n40 10.6151
R2017 B.n709 B.n708 10.6151
R2018 B.n708 B.n707 10.6151
R2019 B.n707 B.n42 10.6151
R2020 B.n703 B.n42 10.6151
R2021 B.n703 B.n702 10.6151
R2022 B.n702 B.n701 10.6151
R2023 B.n701 B.n44 10.6151
R2024 B.n697 B.n44 10.6151
R2025 B.n697 B.n696 10.6151
R2026 B.n696 B.n695 10.6151
R2027 B.n695 B.n46 10.6151
R2028 B.n691 B.n46 10.6151
R2029 B.n691 B.n690 10.6151
R2030 B.n690 B.n689 10.6151
R2031 B.n689 B.n48 10.6151
R2032 B.n685 B.n48 10.6151
R2033 B.n685 B.n684 10.6151
R2034 B.n684 B.n683 10.6151
R2035 B.n683 B.n50 10.6151
R2036 B.n679 B.n678 10.6151
R2037 B.n678 B.n677 10.6151
R2038 B.n677 B.n55 10.6151
R2039 B.n673 B.n55 10.6151
R2040 B.n673 B.n672 10.6151
R2041 B.n672 B.n671 10.6151
R2042 B.n671 B.n57 10.6151
R2043 B.n667 B.n57 10.6151
R2044 B.n665 B.n664 10.6151
R2045 B.n664 B.n61 10.6151
R2046 B.n660 B.n61 10.6151
R2047 B.n660 B.n659 10.6151
R2048 B.n659 B.n658 10.6151
R2049 B.n658 B.n63 10.6151
R2050 B.n654 B.n63 10.6151
R2051 B.n654 B.n653 10.6151
R2052 B.n653 B.n652 10.6151
R2053 B.n652 B.n65 10.6151
R2054 B.n648 B.n65 10.6151
R2055 B.n648 B.n647 10.6151
R2056 B.n647 B.n646 10.6151
R2057 B.n646 B.n67 10.6151
R2058 B.n642 B.n67 10.6151
R2059 B.n642 B.n641 10.6151
R2060 B.n641 B.n640 10.6151
R2061 B.n640 B.n69 10.6151
R2062 B.n636 B.n69 10.6151
R2063 B.n636 B.n635 10.6151
R2064 B.n635 B.n634 10.6151
R2065 B.n634 B.n71 10.6151
R2066 B.n630 B.n71 10.6151
R2067 B.n630 B.n629 10.6151
R2068 B.n629 B.n628 10.6151
R2069 B.n628 B.n73 10.6151
R2070 B.n624 B.n73 10.6151
R2071 B.n624 B.n623 10.6151
R2072 B.n623 B.n622 10.6151
R2073 B.n622 B.n75 10.6151
R2074 B.n618 B.n75 10.6151
R2075 B.n618 B.n617 10.6151
R2076 B.n617 B.n616 10.6151
R2077 B.n616 B.n77 10.6151
R2078 B.n612 B.n77 10.6151
R2079 B.n612 B.n611 10.6151
R2080 B.n611 B.n610 10.6151
R2081 B.n610 B.n79 10.6151
R2082 B.n606 B.n79 10.6151
R2083 B.n606 B.n605 10.6151
R2084 B.n605 B.n604 10.6151
R2085 B.n604 B.n81 10.6151
R2086 B.n600 B.n81 10.6151
R2087 B.n600 B.n599 10.6151
R2088 B.n599 B.n598 10.6151
R2089 B.n598 B.n83 10.6151
R2090 B.n594 B.n83 10.6151
R2091 B.n594 B.n593 10.6151
R2092 B.n593 B.n592 10.6151
R2093 B.n592 B.n85 10.6151
R2094 B.n588 B.n85 10.6151
R2095 B.n588 B.n587 10.6151
R2096 B.n587 B.n586 10.6151
R2097 B.n456 B.n455 10.6151
R2098 B.n456 B.n129 10.6151
R2099 B.n460 B.n129 10.6151
R2100 B.n461 B.n460 10.6151
R2101 B.n462 B.n461 10.6151
R2102 B.n462 B.n127 10.6151
R2103 B.n466 B.n127 10.6151
R2104 B.n467 B.n466 10.6151
R2105 B.n468 B.n467 10.6151
R2106 B.n468 B.n125 10.6151
R2107 B.n472 B.n125 10.6151
R2108 B.n473 B.n472 10.6151
R2109 B.n474 B.n473 10.6151
R2110 B.n474 B.n123 10.6151
R2111 B.n478 B.n123 10.6151
R2112 B.n479 B.n478 10.6151
R2113 B.n480 B.n479 10.6151
R2114 B.n480 B.n121 10.6151
R2115 B.n484 B.n121 10.6151
R2116 B.n485 B.n484 10.6151
R2117 B.n486 B.n485 10.6151
R2118 B.n486 B.n119 10.6151
R2119 B.n490 B.n119 10.6151
R2120 B.n491 B.n490 10.6151
R2121 B.n492 B.n491 10.6151
R2122 B.n492 B.n117 10.6151
R2123 B.n496 B.n117 10.6151
R2124 B.n497 B.n496 10.6151
R2125 B.n498 B.n497 10.6151
R2126 B.n498 B.n115 10.6151
R2127 B.n502 B.n115 10.6151
R2128 B.n503 B.n502 10.6151
R2129 B.n504 B.n503 10.6151
R2130 B.n504 B.n113 10.6151
R2131 B.n508 B.n113 10.6151
R2132 B.n509 B.n508 10.6151
R2133 B.n510 B.n509 10.6151
R2134 B.n510 B.n111 10.6151
R2135 B.n514 B.n111 10.6151
R2136 B.n515 B.n514 10.6151
R2137 B.n516 B.n515 10.6151
R2138 B.n516 B.n109 10.6151
R2139 B.n520 B.n109 10.6151
R2140 B.n521 B.n520 10.6151
R2141 B.n522 B.n521 10.6151
R2142 B.n522 B.n107 10.6151
R2143 B.n526 B.n107 10.6151
R2144 B.n527 B.n526 10.6151
R2145 B.n528 B.n527 10.6151
R2146 B.n528 B.n105 10.6151
R2147 B.n532 B.n105 10.6151
R2148 B.n533 B.n532 10.6151
R2149 B.n534 B.n533 10.6151
R2150 B.n534 B.n103 10.6151
R2151 B.n538 B.n103 10.6151
R2152 B.n539 B.n538 10.6151
R2153 B.n540 B.n539 10.6151
R2154 B.n540 B.n101 10.6151
R2155 B.n544 B.n101 10.6151
R2156 B.n545 B.n544 10.6151
R2157 B.n546 B.n545 10.6151
R2158 B.n546 B.n99 10.6151
R2159 B.n550 B.n99 10.6151
R2160 B.n551 B.n550 10.6151
R2161 B.n552 B.n551 10.6151
R2162 B.n552 B.n97 10.6151
R2163 B.n556 B.n97 10.6151
R2164 B.n557 B.n556 10.6151
R2165 B.n558 B.n557 10.6151
R2166 B.n558 B.n95 10.6151
R2167 B.n562 B.n95 10.6151
R2168 B.n563 B.n562 10.6151
R2169 B.n564 B.n563 10.6151
R2170 B.n564 B.n93 10.6151
R2171 B.n568 B.n93 10.6151
R2172 B.n569 B.n568 10.6151
R2173 B.n570 B.n569 10.6151
R2174 B.n570 B.n91 10.6151
R2175 B.n574 B.n91 10.6151
R2176 B.n575 B.n574 10.6151
R2177 B.n576 B.n575 10.6151
R2178 B.n576 B.n89 10.6151
R2179 B.n580 B.n89 10.6151
R2180 B.n581 B.n580 10.6151
R2181 B.n582 B.n581 10.6151
R2182 B.n582 B.n87 10.6151
R2183 B.n277 B.n276 10.6151
R2184 B.n278 B.n277 10.6151
R2185 B.n278 B.n189 10.6151
R2186 B.n282 B.n189 10.6151
R2187 B.n283 B.n282 10.6151
R2188 B.n284 B.n283 10.6151
R2189 B.n284 B.n187 10.6151
R2190 B.n288 B.n187 10.6151
R2191 B.n289 B.n288 10.6151
R2192 B.n290 B.n289 10.6151
R2193 B.n290 B.n185 10.6151
R2194 B.n294 B.n185 10.6151
R2195 B.n295 B.n294 10.6151
R2196 B.n296 B.n295 10.6151
R2197 B.n296 B.n183 10.6151
R2198 B.n300 B.n183 10.6151
R2199 B.n301 B.n300 10.6151
R2200 B.n302 B.n301 10.6151
R2201 B.n302 B.n181 10.6151
R2202 B.n306 B.n181 10.6151
R2203 B.n307 B.n306 10.6151
R2204 B.n308 B.n307 10.6151
R2205 B.n308 B.n179 10.6151
R2206 B.n312 B.n179 10.6151
R2207 B.n313 B.n312 10.6151
R2208 B.n314 B.n313 10.6151
R2209 B.n314 B.n177 10.6151
R2210 B.n318 B.n177 10.6151
R2211 B.n319 B.n318 10.6151
R2212 B.n320 B.n319 10.6151
R2213 B.n320 B.n175 10.6151
R2214 B.n324 B.n175 10.6151
R2215 B.n325 B.n324 10.6151
R2216 B.n326 B.n325 10.6151
R2217 B.n326 B.n173 10.6151
R2218 B.n330 B.n173 10.6151
R2219 B.n331 B.n330 10.6151
R2220 B.n332 B.n331 10.6151
R2221 B.n332 B.n171 10.6151
R2222 B.n336 B.n171 10.6151
R2223 B.n337 B.n336 10.6151
R2224 B.n338 B.n337 10.6151
R2225 B.n338 B.n169 10.6151
R2226 B.n342 B.n169 10.6151
R2227 B.n343 B.n342 10.6151
R2228 B.n344 B.n343 10.6151
R2229 B.n344 B.n167 10.6151
R2230 B.n348 B.n167 10.6151
R2231 B.n349 B.n348 10.6151
R2232 B.n350 B.n349 10.6151
R2233 B.n350 B.n165 10.6151
R2234 B.n354 B.n165 10.6151
R2235 B.n355 B.n354 10.6151
R2236 B.n357 B.n161 10.6151
R2237 B.n361 B.n161 10.6151
R2238 B.n362 B.n361 10.6151
R2239 B.n363 B.n362 10.6151
R2240 B.n363 B.n159 10.6151
R2241 B.n367 B.n159 10.6151
R2242 B.n368 B.n367 10.6151
R2243 B.n372 B.n368 10.6151
R2244 B.n376 B.n157 10.6151
R2245 B.n377 B.n376 10.6151
R2246 B.n378 B.n377 10.6151
R2247 B.n378 B.n155 10.6151
R2248 B.n382 B.n155 10.6151
R2249 B.n383 B.n382 10.6151
R2250 B.n384 B.n383 10.6151
R2251 B.n384 B.n153 10.6151
R2252 B.n388 B.n153 10.6151
R2253 B.n389 B.n388 10.6151
R2254 B.n390 B.n389 10.6151
R2255 B.n390 B.n151 10.6151
R2256 B.n394 B.n151 10.6151
R2257 B.n395 B.n394 10.6151
R2258 B.n396 B.n395 10.6151
R2259 B.n396 B.n149 10.6151
R2260 B.n400 B.n149 10.6151
R2261 B.n401 B.n400 10.6151
R2262 B.n402 B.n401 10.6151
R2263 B.n402 B.n147 10.6151
R2264 B.n406 B.n147 10.6151
R2265 B.n407 B.n406 10.6151
R2266 B.n408 B.n407 10.6151
R2267 B.n408 B.n145 10.6151
R2268 B.n412 B.n145 10.6151
R2269 B.n413 B.n412 10.6151
R2270 B.n414 B.n413 10.6151
R2271 B.n414 B.n143 10.6151
R2272 B.n418 B.n143 10.6151
R2273 B.n419 B.n418 10.6151
R2274 B.n420 B.n419 10.6151
R2275 B.n420 B.n141 10.6151
R2276 B.n424 B.n141 10.6151
R2277 B.n425 B.n424 10.6151
R2278 B.n426 B.n425 10.6151
R2279 B.n426 B.n139 10.6151
R2280 B.n430 B.n139 10.6151
R2281 B.n431 B.n430 10.6151
R2282 B.n432 B.n431 10.6151
R2283 B.n432 B.n137 10.6151
R2284 B.n436 B.n137 10.6151
R2285 B.n437 B.n436 10.6151
R2286 B.n438 B.n437 10.6151
R2287 B.n438 B.n135 10.6151
R2288 B.n442 B.n135 10.6151
R2289 B.n443 B.n442 10.6151
R2290 B.n444 B.n443 10.6151
R2291 B.n444 B.n133 10.6151
R2292 B.n448 B.n133 10.6151
R2293 B.n449 B.n448 10.6151
R2294 B.n450 B.n449 10.6151
R2295 B.n450 B.n131 10.6151
R2296 B.n454 B.n131 10.6151
R2297 B.n272 B.n191 10.6151
R2298 B.n272 B.n271 10.6151
R2299 B.n271 B.n270 10.6151
R2300 B.n270 B.n193 10.6151
R2301 B.n266 B.n193 10.6151
R2302 B.n266 B.n265 10.6151
R2303 B.n265 B.n264 10.6151
R2304 B.n264 B.n195 10.6151
R2305 B.n260 B.n195 10.6151
R2306 B.n260 B.n259 10.6151
R2307 B.n259 B.n258 10.6151
R2308 B.n258 B.n197 10.6151
R2309 B.n254 B.n197 10.6151
R2310 B.n254 B.n253 10.6151
R2311 B.n253 B.n252 10.6151
R2312 B.n252 B.n199 10.6151
R2313 B.n248 B.n199 10.6151
R2314 B.n248 B.n247 10.6151
R2315 B.n247 B.n246 10.6151
R2316 B.n246 B.n201 10.6151
R2317 B.n242 B.n201 10.6151
R2318 B.n242 B.n241 10.6151
R2319 B.n241 B.n240 10.6151
R2320 B.n240 B.n203 10.6151
R2321 B.n236 B.n203 10.6151
R2322 B.n236 B.n235 10.6151
R2323 B.n235 B.n234 10.6151
R2324 B.n234 B.n205 10.6151
R2325 B.n230 B.n205 10.6151
R2326 B.n230 B.n229 10.6151
R2327 B.n229 B.n228 10.6151
R2328 B.n228 B.n207 10.6151
R2329 B.n224 B.n207 10.6151
R2330 B.n224 B.n223 10.6151
R2331 B.n223 B.n222 10.6151
R2332 B.n222 B.n209 10.6151
R2333 B.n218 B.n209 10.6151
R2334 B.n218 B.n217 10.6151
R2335 B.n217 B.n216 10.6151
R2336 B.n216 B.n211 10.6151
R2337 B.n212 B.n211 10.6151
R2338 B.n212 B.n0 10.6151
R2339 B.n823 B.n1 10.6151
R2340 B.n823 B.n822 10.6151
R2341 B.n822 B.n821 10.6151
R2342 B.n821 B.n4 10.6151
R2343 B.n817 B.n4 10.6151
R2344 B.n817 B.n816 10.6151
R2345 B.n816 B.n815 10.6151
R2346 B.n815 B.n6 10.6151
R2347 B.n811 B.n6 10.6151
R2348 B.n811 B.n810 10.6151
R2349 B.n810 B.n809 10.6151
R2350 B.n809 B.n8 10.6151
R2351 B.n805 B.n8 10.6151
R2352 B.n805 B.n804 10.6151
R2353 B.n804 B.n803 10.6151
R2354 B.n803 B.n10 10.6151
R2355 B.n799 B.n10 10.6151
R2356 B.n799 B.n798 10.6151
R2357 B.n798 B.n797 10.6151
R2358 B.n797 B.n12 10.6151
R2359 B.n793 B.n12 10.6151
R2360 B.n793 B.n792 10.6151
R2361 B.n792 B.n791 10.6151
R2362 B.n791 B.n14 10.6151
R2363 B.n787 B.n14 10.6151
R2364 B.n787 B.n786 10.6151
R2365 B.n786 B.n785 10.6151
R2366 B.n785 B.n16 10.6151
R2367 B.n781 B.n16 10.6151
R2368 B.n781 B.n780 10.6151
R2369 B.n780 B.n779 10.6151
R2370 B.n779 B.n18 10.6151
R2371 B.n775 B.n18 10.6151
R2372 B.n775 B.n774 10.6151
R2373 B.n774 B.n773 10.6151
R2374 B.n773 B.n20 10.6151
R2375 B.n769 B.n20 10.6151
R2376 B.n769 B.n768 10.6151
R2377 B.n768 B.n767 10.6151
R2378 B.n767 B.n22 10.6151
R2379 B.n763 B.n22 10.6151
R2380 B.n763 B.n762 10.6151
R2381 B.n679 B.n54 6.5566
R2382 B.n667 B.n666 6.5566
R2383 B.n357 B.n356 6.5566
R2384 B.n372 B.n371 6.5566
R2385 B.n54 B.n50 4.05904
R2386 B.n666 B.n665 4.05904
R2387 B.n356 B.n355 4.05904
R2388 B.n371 B.n157 4.05904
R2389 B.n827 B.n0 2.81026
R2390 B.n827 B.n1 2.81026
C0 VP VTAIL 6.50345f
C1 VDD2 w_n3334_n4204# 1.83516f
C2 w_n3334_n4204# VN 5.89749f
C3 VP VDD1 6.93121f
C4 VTAIL VDD1 6.56333f
C5 w_n3334_n4204# VP 6.32864f
C6 VDD2 B 1.62211f
C7 w_n3334_n4204# VTAIL 4.9203f
C8 B VN 1.35406f
C9 VDD2 VN 6.62355f
C10 w_n3334_n4204# VDD1 1.75676f
C11 B VP 2.07424f
C12 VDD2 VP 0.459059f
C13 B VTAIL 6.79679f
C14 VDD2 VTAIL 6.62431f
C15 VP VN 7.68651f
C16 VN VTAIL 6.48934f
C17 B VDD1 1.55324f
C18 VDD2 VDD1 1.27025f
C19 VN VDD1 0.150399f
C20 w_n3334_n4204# B 11.6596f
C21 VDD2 VSUBS 1.208947f
C22 VDD1 VSUBS 6.82901f
C23 VTAIL VSUBS 1.531992f
C24 VN VSUBS 6.13295f
C25 VP VSUBS 2.974456f
C26 B VSUBS 5.498695f
C27 w_n3334_n4204# VSUBS 0.171674p
C28 B.n0 VSUBS 0.004014f
C29 B.n1 VSUBS 0.004014f
C30 B.n2 VSUBS 0.006347f
C31 B.n3 VSUBS 0.006347f
C32 B.n4 VSUBS 0.006347f
C33 B.n5 VSUBS 0.006347f
C34 B.n6 VSUBS 0.006347f
C35 B.n7 VSUBS 0.006347f
C36 B.n8 VSUBS 0.006347f
C37 B.n9 VSUBS 0.006347f
C38 B.n10 VSUBS 0.006347f
C39 B.n11 VSUBS 0.006347f
C40 B.n12 VSUBS 0.006347f
C41 B.n13 VSUBS 0.006347f
C42 B.n14 VSUBS 0.006347f
C43 B.n15 VSUBS 0.006347f
C44 B.n16 VSUBS 0.006347f
C45 B.n17 VSUBS 0.006347f
C46 B.n18 VSUBS 0.006347f
C47 B.n19 VSUBS 0.006347f
C48 B.n20 VSUBS 0.006347f
C49 B.n21 VSUBS 0.006347f
C50 B.n22 VSUBS 0.006347f
C51 B.n23 VSUBS 0.014875f
C52 B.n24 VSUBS 0.006347f
C53 B.n25 VSUBS 0.006347f
C54 B.n26 VSUBS 0.006347f
C55 B.n27 VSUBS 0.006347f
C56 B.n28 VSUBS 0.006347f
C57 B.n29 VSUBS 0.006347f
C58 B.n30 VSUBS 0.006347f
C59 B.n31 VSUBS 0.006347f
C60 B.n32 VSUBS 0.006347f
C61 B.n33 VSUBS 0.006347f
C62 B.n34 VSUBS 0.006347f
C63 B.n35 VSUBS 0.006347f
C64 B.n36 VSUBS 0.006347f
C65 B.n37 VSUBS 0.006347f
C66 B.n38 VSUBS 0.006347f
C67 B.n39 VSUBS 0.006347f
C68 B.n40 VSUBS 0.006347f
C69 B.n41 VSUBS 0.006347f
C70 B.n42 VSUBS 0.006347f
C71 B.n43 VSUBS 0.006347f
C72 B.n44 VSUBS 0.006347f
C73 B.n45 VSUBS 0.006347f
C74 B.n46 VSUBS 0.006347f
C75 B.n47 VSUBS 0.006347f
C76 B.n48 VSUBS 0.006347f
C77 B.n49 VSUBS 0.006347f
C78 B.n50 VSUBS 0.004387f
C79 B.n51 VSUBS 0.006347f
C80 B.t5 VSUBS 0.278809f
C81 B.t4 VSUBS 0.318316f
C82 B.t3 VSUBS 2.42097f
C83 B.n52 VSUBS 0.506264f
C84 B.n53 VSUBS 0.281712f
C85 B.n54 VSUBS 0.014706f
C86 B.n55 VSUBS 0.006347f
C87 B.n56 VSUBS 0.006347f
C88 B.n57 VSUBS 0.006347f
C89 B.n58 VSUBS 0.006347f
C90 B.t8 VSUBS 0.278812f
C91 B.t7 VSUBS 0.318318f
C92 B.t6 VSUBS 2.42097f
C93 B.n59 VSUBS 0.506262f
C94 B.n60 VSUBS 0.281708f
C95 B.n61 VSUBS 0.006347f
C96 B.n62 VSUBS 0.006347f
C97 B.n63 VSUBS 0.006347f
C98 B.n64 VSUBS 0.006347f
C99 B.n65 VSUBS 0.006347f
C100 B.n66 VSUBS 0.006347f
C101 B.n67 VSUBS 0.006347f
C102 B.n68 VSUBS 0.006347f
C103 B.n69 VSUBS 0.006347f
C104 B.n70 VSUBS 0.006347f
C105 B.n71 VSUBS 0.006347f
C106 B.n72 VSUBS 0.006347f
C107 B.n73 VSUBS 0.006347f
C108 B.n74 VSUBS 0.006347f
C109 B.n75 VSUBS 0.006347f
C110 B.n76 VSUBS 0.006347f
C111 B.n77 VSUBS 0.006347f
C112 B.n78 VSUBS 0.006347f
C113 B.n79 VSUBS 0.006347f
C114 B.n80 VSUBS 0.006347f
C115 B.n81 VSUBS 0.006347f
C116 B.n82 VSUBS 0.006347f
C117 B.n83 VSUBS 0.006347f
C118 B.n84 VSUBS 0.006347f
C119 B.n85 VSUBS 0.006347f
C120 B.n86 VSUBS 0.006347f
C121 B.n87 VSUBS 0.015612f
C122 B.n88 VSUBS 0.006347f
C123 B.n89 VSUBS 0.006347f
C124 B.n90 VSUBS 0.006347f
C125 B.n91 VSUBS 0.006347f
C126 B.n92 VSUBS 0.006347f
C127 B.n93 VSUBS 0.006347f
C128 B.n94 VSUBS 0.006347f
C129 B.n95 VSUBS 0.006347f
C130 B.n96 VSUBS 0.006347f
C131 B.n97 VSUBS 0.006347f
C132 B.n98 VSUBS 0.006347f
C133 B.n99 VSUBS 0.006347f
C134 B.n100 VSUBS 0.006347f
C135 B.n101 VSUBS 0.006347f
C136 B.n102 VSUBS 0.006347f
C137 B.n103 VSUBS 0.006347f
C138 B.n104 VSUBS 0.006347f
C139 B.n105 VSUBS 0.006347f
C140 B.n106 VSUBS 0.006347f
C141 B.n107 VSUBS 0.006347f
C142 B.n108 VSUBS 0.006347f
C143 B.n109 VSUBS 0.006347f
C144 B.n110 VSUBS 0.006347f
C145 B.n111 VSUBS 0.006347f
C146 B.n112 VSUBS 0.006347f
C147 B.n113 VSUBS 0.006347f
C148 B.n114 VSUBS 0.006347f
C149 B.n115 VSUBS 0.006347f
C150 B.n116 VSUBS 0.006347f
C151 B.n117 VSUBS 0.006347f
C152 B.n118 VSUBS 0.006347f
C153 B.n119 VSUBS 0.006347f
C154 B.n120 VSUBS 0.006347f
C155 B.n121 VSUBS 0.006347f
C156 B.n122 VSUBS 0.006347f
C157 B.n123 VSUBS 0.006347f
C158 B.n124 VSUBS 0.006347f
C159 B.n125 VSUBS 0.006347f
C160 B.n126 VSUBS 0.006347f
C161 B.n127 VSUBS 0.006347f
C162 B.n128 VSUBS 0.006347f
C163 B.n129 VSUBS 0.006347f
C164 B.n130 VSUBS 0.014875f
C165 B.n131 VSUBS 0.006347f
C166 B.n132 VSUBS 0.006347f
C167 B.n133 VSUBS 0.006347f
C168 B.n134 VSUBS 0.006347f
C169 B.n135 VSUBS 0.006347f
C170 B.n136 VSUBS 0.006347f
C171 B.n137 VSUBS 0.006347f
C172 B.n138 VSUBS 0.006347f
C173 B.n139 VSUBS 0.006347f
C174 B.n140 VSUBS 0.006347f
C175 B.n141 VSUBS 0.006347f
C176 B.n142 VSUBS 0.006347f
C177 B.n143 VSUBS 0.006347f
C178 B.n144 VSUBS 0.006347f
C179 B.n145 VSUBS 0.006347f
C180 B.n146 VSUBS 0.006347f
C181 B.n147 VSUBS 0.006347f
C182 B.n148 VSUBS 0.006347f
C183 B.n149 VSUBS 0.006347f
C184 B.n150 VSUBS 0.006347f
C185 B.n151 VSUBS 0.006347f
C186 B.n152 VSUBS 0.006347f
C187 B.n153 VSUBS 0.006347f
C188 B.n154 VSUBS 0.006347f
C189 B.n155 VSUBS 0.006347f
C190 B.n156 VSUBS 0.006347f
C191 B.n157 VSUBS 0.004387f
C192 B.n158 VSUBS 0.006347f
C193 B.n159 VSUBS 0.006347f
C194 B.n160 VSUBS 0.006347f
C195 B.n161 VSUBS 0.006347f
C196 B.n162 VSUBS 0.006347f
C197 B.t10 VSUBS 0.278809f
C198 B.t11 VSUBS 0.318316f
C199 B.t9 VSUBS 2.42097f
C200 B.n163 VSUBS 0.506264f
C201 B.n164 VSUBS 0.281712f
C202 B.n165 VSUBS 0.006347f
C203 B.n166 VSUBS 0.006347f
C204 B.n167 VSUBS 0.006347f
C205 B.n168 VSUBS 0.006347f
C206 B.n169 VSUBS 0.006347f
C207 B.n170 VSUBS 0.006347f
C208 B.n171 VSUBS 0.006347f
C209 B.n172 VSUBS 0.006347f
C210 B.n173 VSUBS 0.006347f
C211 B.n174 VSUBS 0.006347f
C212 B.n175 VSUBS 0.006347f
C213 B.n176 VSUBS 0.006347f
C214 B.n177 VSUBS 0.006347f
C215 B.n178 VSUBS 0.006347f
C216 B.n179 VSUBS 0.006347f
C217 B.n180 VSUBS 0.006347f
C218 B.n181 VSUBS 0.006347f
C219 B.n182 VSUBS 0.006347f
C220 B.n183 VSUBS 0.006347f
C221 B.n184 VSUBS 0.006347f
C222 B.n185 VSUBS 0.006347f
C223 B.n186 VSUBS 0.006347f
C224 B.n187 VSUBS 0.006347f
C225 B.n188 VSUBS 0.006347f
C226 B.n189 VSUBS 0.006347f
C227 B.n190 VSUBS 0.006347f
C228 B.n191 VSUBS 0.014875f
C229 B.n192 VSUBS 0.006347f
C230 B.n193 VSUBS 0.006347f
C231 B.n194 VSUBS 0.006347f
C232 B.n195 VSUBS 0.006347f
C233 B.n196 VSUBS 0.006347f
C234 B.n197 VSUBS 0.006347f
C235 B.n198 VSUBS 0.006347f
C236 B.n199 VSUBS 0.006347f
C237 B.n200 VSUBS 0.006347f
C238 B.n201 VSUBS 0.006347f
C239 B.n202 VSUBS 0.006347f
C240 B.n203 VSUBS 0.006347f
C241 B.n204 VSUBS 0.006347f
C242 B.n205 VSUBS 0.006347f
C243 B.n206 VSUBS 0.006347f
C244 B.n207 VSUBS 0.006347f
C245 B.n208 VSUBS 0.006347f
C246 B.n209 VSUBS 0.006347f
C247 B.n210 VSUBS 0.006347f
C248 B.n211 VSUBS 0.006347f
C249 B.n212 VSUBS 0.006347f
C250 B.n213 VSUBS 0.006347f
C251 B.n214 VSUBS 0.006347f
C252 B.n215 VSUBS 0.006347f
C253 B.n216 VSUBS 0.006347f
C254 B.n217 VSUBS 0.006347f
C255 B.n218 VSUBS 0.006347f
C256 B.n219 VSUBS 0.006347f
C257 B.n220 VSUBS 0.006347f
C258 B.n221 VSUBS 0.006347f
C259 B.n222 VSUBS 0.006347f
C260 B.n223 VSUBS 0.006347f
C261 B.n224 VSUBS 0.006347f
C262 B.n225 VSUBS 0.006347f
C263 B.n226 VSUBS 0.006347f
C264 B.n227 VSUBS 0.006347f
C265 B.n228 VSUBS 0.006347f
C266 B.n229 VSUBS 0.006347f
C267 B.n230 VSUBS 0.006347f
C268 B.n231 VSUBS 0.006347f
C269 B.n232 VSUBS 0.006347f
C270 B.n233 VSUBS 0.006347f
C271 B.n234 VSUBS 0.006347f
C272 B.n235 VSUBS 0.006347f
C273 B.n236 VSUBS 0.006347f
C274 B.n237 VSUBS 0.006347f
C275 B.n238 VSUBS 0.006347f
C276 B.n239 VSUBS 0.006347f
C277 B.n240 VSUBS 0.006347f
C278 B.n241 VSUBS 0.006347f
C279 B.n242 VSUBS 0.006347f
C280 B.n243 VSUBS 0.006347f
C281 B.n244 VSUBS 0.006347f
C282 B.n245 VSUBS 0.006347f
C283 B.n246 VSUBS 0.006347f
C284 B.n247 VSUBS 0.006347f
C285 B.n248 VSUBS 0.006347f
C286 B.n249 VSUBS 0.006347f
C287 B.n250 VSUBS 0.006347f
C288 B.n251 VSUBS 0.006347f
C289 B.n252 VSUBS 0.006347f
C290 B.n253 VSUBS 0.006347f
C291 B.n254 VSUBS 0.006347f
C292 B.n255 VSUBS 0.006347f
C293 B.n256 VSUBS 0.006347f
C294 B.n257 VSUBS 0.006347f
C295 B.n258 VSUBS 0.006347f
C296 B.n259 VSUBS 0.006347f
C297 B.n260 VSUBS 0.006347f
C298 B.n261 VSUBS 0.006347f
C299 B.n262 VSUBS 0.006347f
C300 B.n263 VSUBS 0.006347f
C301 B.n264 VSUBS 0.006347f
C302 B.n265 VSUBS 0.006347f
C303 B.n266 VSUBS 0.006347f
C304 B.n267 VSUBS 0.006347f
C305 B.n268 VSUBS 0.006347f
C306 B.n269 VSUBS 0.006347f
C307 B.n270 VSUBS 0.006347f
C308 B.n271 VSUBS 0.006347f
C309 B.n272 VSUBS 0.006347f
C310 B.n273 VSUBS 0.006347f
C311 B.n274 VSUBS 0.014875f
C312 B.n275 VSUBS 0.015181f
C313 B.n276 VSUBS 0.015181f
C314 B.n277 VSUBS 0.006347f
C315 B.n278 VSUBS 0.006347f
C316 B.n279 VSUBS 0.006347f
C317 B.n280 VSUBS 0.006347f
C318 B.n281 VSUBS 0.006347f
C319 B.n282 VSUBS 0.006347f
C320 B.n283 VSUBS 0.006347f
C321 B.n284 VSUBS 0.006347f
C322 B.n285 VSUBS 0.006347f
C323 B.n286 VSUBS 0.006347f
C324 B.n287 VSUBS 0.006347f
C325 B.n288 VSUBS 0.006347f
C326 B.n289 VSUBS 0.006347f
C327 B.n290 VSUBS 0.006347f
C328 B.n291 VSUBS 0.006347f
C329 B.n292 VSUBS 0.006347f
C330 B.n293 VSUBS 0.006347f
C331 B.n294 VSUBS 0.006347f
C332 B.n295 VSUBS 0.006347f
C333 B.n296 VSUBS 0.006347f
C334 B.n297 VSUBS 0.006347f
C335 B.n298 VSUBS 0.006347f
C336 B.n299 VSUBS 0.006347f
C337 B.n300 VSUBS 0.006347f
C338 B.n301 VSUBS 0.006347f
C339 B.n302 VSUBS 0.006347f
C340 B.n303 VSUBS 0.006347f
C341 B.n304 VSUBS 0.006347f
C342 B.n305 VSUBS 0.006347f
C343 B.n306 VSUBS 0.006347f
C344 B.n307 VSUBS 0.006347f
C345 B.n308 VSUBS 0.006347f
C346 B.n309 VSUBS 0.006347f
C347 B.n310 VSUBS 0.006347f
C348 B.n311 VSUBS 0.006347f
C349 B.n312 VSUBS 0.006347f
C350 B.n313 VSUBS 0.006347f
C351 B.n314 VSUBS 0.006347f
C352 B.n315 VSUBS 0.006347f
C353 B.n316 VSUBS 0.006347f
C354 B.n317 VSUBS 0.006347f
C355 B.n318 VSUBS 0.006347f
C356 B.n319 VSUBS 0.006347f
C357 B.n320 VSUBS 0.006347f
C358 B.n321 VSUBS 0.006347f
C359 B.n322 VSUBS 0.006347f
C360 B.n323 VSUBS 0.006347f
C361 B.n324 VSUBS 0.006347f
C362 B.n325 VSUBS 0.006347f
C363 B.n326 VSUBS 0.006347f
C364 B.n327 VSUBS 0.006347f
C365 B.n328 VSUBS 0.006347f
C366 B.n329 VSUBS 0.006347f
C367 B.n330 VSUBS 0.006347f
C368 B.n331 VSUBS 0.006347f
C369 B.n332 VSUBS 0.006347f
C370 B.n333 VSUBS 0.006347f
C371 B.n334 VSUBS 0.006347f
C372 B.n335 VSUBS 0.006347f
C373 B.n336 VSUBS 0.006347f
C374 B.n337 VSUBS 0.006347f
C375 B.n338 VSUBS 0.006347f
C376 B.n339 VSUBS 0.006347f
C377 B.n340 VSUBS 0.006347f
C378 B.n341 VSUBS 0.006347f
C379 B.n342 VSUBS 0.006347f
C380 B.n343 VSUBS 0.006347f
C381 B.n344 VSUBS 0.006347f
C382 B.n345 VSUBS 0.006347f
C383 B.n346 VSUBS 0.006347f
C384 B.n347 VSUBS 0.006347f
C385 B.n348 VSUBS 0.006347f
C386 B.n349 VSUBS 0.006347f
C387 B.n350 VSUBS 0.006347f
C388 B.n351 VSUBS 0.006347f
C389 B.n352 VSUBS 0.006347f
C390 B.n353 VSUBS 0.006347f
C391 B.n354 VSUBS 0.006347f
C392 B.n355 VSUBS 0.004387f
C393 B.n356 VSUBS 0.014706f
C394 B.n357 VSUBS 0.005134f
C395 B.n358 VSUBS 0.006347f
C396 B.n359 VSUBS 0.006347f
C397 B.n360 VSUBS 0.006347f
C398 B.n361 VSUBS 0.006347f
C399 B.n362 VSUBS 0.006347f
C400 B.n363 VSUBS 0.006347f
C401 B.n364 VSUBS 0.006347f
C402 B.n365 VSUBS 0.006347f
C403 B.n366 VSUBS 0.006347f
C404 B.n367 VSUBS 0.006347f
C405 B.n368 VSUBS 0.006347f
C406 B.t1 VSUBS 0.278812f
C407 B.t2 VSUBS 0.318318f
C408 B.t0 VSUBS 2.42097f
C409 B.n369 VSUBS 0.506262f
C410 B.n370 VSUBS 0.281708f
C411 B.n371 VSUBS 0.014706f
C412 B.n372 VSUBS 0.005134f
C413 B.n373 VSUBS 0.006347f
C414 B.n374 VSUBS 0.006347f
C415 B.n375 VSUBS 0.006347f
C416 B.n376 VSUBS 0.006347f
C417 B.n377 VSUBS 0.006347f
C418 B.n378 VSUBS 0.006347f
C419 B.n379 VSUBS 0.006347f
C420 B.n380 VSUBS 0.006347f
C421 B.n381 VSUBS 0.006347f
C422 B.n382 VSUBS 0.006347f
C423 B.n383 VSUBS 0.006347f
C424 B.n384 VSUBS 0.006347f
C425 B.n385 VSUBS 0.006347f
C426 B.n386 VSUBS 0.006347f
C427 B.n387 VSUBS 0.006347f
C428 B.n388 VSUBS 0.006347f
C429 B.n389 VSUBS 0.006347f
C430 B.n390 VSUBS 0.006347f
C431 B.n391 VSUBS 0.006347f
C432 B.n392 VSUBS 0.006347f
C433 B.n393 VSUBS 0.006347f
C434 B.n394 VSUBS 0.006347f
C435 B.n395 VSUBS 0.006347f
C436 B.n396 VSUBS 0.006347f
C437 B.n397 VSUBS 0.006347f
C438 B.n398 VSUBS 0.006347f
C439 B.n399 VSUBS 0.006347f
C440 B.n400 VSUBS 0.006347f
C441 B.n401 VSUBS 0.006347f
C442 B.n402 VSUBS 0.006347f
C443 B.n403 VSUBS 0.006347f
C444 B.n404 VSUBS 0.006347f
C445 B.n405 VSUBS 0.006347f
C446 B.n406 VSUBS 0.006347f
C447 B.n407 VSUBS 0.006347f
C448 B.n408 VSUBS 0.006347f
C449 B.n409 VSUBS 0.006347f
C450 B.n410 VSUBS 0.006347f
C451 B.n411 VSUBS 0.006347f
C452 B.n412 VSUBS 0.006347f
C453 B.n413 VSUBS 0.006347f
C454 B.n414 VSUBS 0.006347f
C455 B.n415 VSUBS 0.006347f
C456 B.n416 VSUBS 0.006347f
C457 B.n417 VSUBS 0.006347f
C458 B.n418 VSUBS 0.006347f
C459 B.n419 VSUBS 0.006347f
C460 B.n420 VSUBS 0.006347f
C461 B.n421 VSUBS 0.006347f
C462 B.n422 VSUBS 0.006347f
C463 B.n423 VSUBS 0.006347f
C464 B.n424 VSUBS 0.006347f
C465 B.n425 VSUBS 0.006347f
C466 B.n426 VSUBS 0.006347f
C467 B.n427 VSUBS 0.006347f
C468 B.n428 VSUBS 0.006347f
C469 B.n429 VSUBS 0.006347f
C470 B.n430 VSUBS 0.006347f
C471 B.n431 VSUBS 0.006347f
C472 B.n432 VSUBS 0.006347f
C473 B.n433 VSUBS 0.006347f
C474 B.n434 VSUBS 0.006347f
C475 B.n435 VSUBS 0.006347f
C476 B.n436 VSUBS 0.006347f
C477 B.n437 VSUBS 0.006347f
C478 B.n438 VSUBS 0.006347f
C479 B.n439 VSUBS 0.006347f
C480 B.n440 VSUBS 0.006347f
C481 B.n441 VSUBS 0.006347f
C482 B.n442 VSUBS 0.006347f
C483 B.n443 VSUBS 0.006347f
C484 B.n444 VSUBS 0.006347f
C485 B.n445 VSUBS 0.006347f
C486 B.n446 VSUBS 0.006347f
C487 B.n447 VSUBS 0.006347f
C488 B.n448 VSUBS 0.006347f
C489 B.n449 VSUBS 0.006347f
C490 B.n450 VSUBS 0.006347f
C491 B.n451 VSUBS 0.006347f
C492 B.n452 VSUBS 0.006347f
C493 B.n453 VSUBS 0.015181f
C494 B.n454 VSUBS 0.015181f
C495 B.n455 VSUBS 0.014875f
C496 B.n456 VSUBS 0.006347f
C497 B.n457 VSUBS 0.006347f
C498 B.n458 VSUBS 0.006347f
C499 B.n459 VSUBS 0.006347f
C500 B.n460 VSUBS 0.006347f
C501 B.n461 VSUBS 0.006347f
C502 B.n462 VSUBS 0.006347f
C503 B.n463 VSUBS 0.006347f
C504 B.n464 VSUBS 0.006347f
C505 B.n465 VSUBS 0.006347f
C506 B.n466 VSUBS 0.006347f
C507 B.n467 VSUBS 0.006347f
C508 B.n468 VSUBS 0.006347f
C509 B.n469 VSUBS 0.006347f
C510 B.n470 VSUBS 0.006347f
C511 B.n471 VSUBS 0.006347f
C512 B.n472 VSUBS 0.006347f
C513 B.n473 VSUBS 0.006347f
C514 B.n474 VSUBS 0.006347f
C515 B.n475 VSUBS 0.006347f
C516 B.n476 VSUBS 0.006347f
C517 B.n477 VSUBS 0.006347f
C518 B.n478 VSUBS 0.006347f
C519 B.n479 VSUBS 0.006347f
C520 B.n480 VSUBS 0.006347f
C521 B.n481 VSUBS 0.006347f
C522 B.n482 VSUBS 0.006347f
C523 B.n483 VSUBS 0.006347f
C524 B.n484 VSUBS 0.006347f
C525 B.n485 VSUBS 0.006347f
C526 B.n486 VSUBS 0.006347f
C527 B.n487 VSUBS 0.006347f
C528 B.n488 VSUBS 0.006347f
C529 B.n489 VSUBS 0.006347f
C530 B.n490 VSUBS 0.006347f
C531 B.n491 VSUBS 0.006347f
C532 B.n492 VSUBS 0.006347f
C533 B.n493 VSUBS 0.006347f
C534 B.n494 VSUBS 0.006347f
C535 B.n495 VSUBS 0.006347f
C536 B.n496 VSUBS 0.006347f
C537 B.n497 VSUBS 0.006347f
C538 B.n498 VSUBS 0.006347f
C539 B.n499 VSUBS 0.006347f
C540 B.n500 VSUBS 0.006347f
C541 B.n501 VSUBS 0.006347f
C542 B.n502 VSUBS 0.006347f
C543 B.n503 VSUBS 0.006347f
C544 B.n504 VSUBS 0.006347f
C545 B.n505 VSUBS 0.006347f
C546 B.n506 VSUBS 0.006347f
C547 B.n507 VSUBS 0.006347f
C548 B.n508 VSUBS 0.006347f
C549 B.n509 VSUBS 0.006347f
C550 B.n510 VSUBS 0.006347f
C551 B.n511 VSUBS 0.006347f
C552 B.n512 VSUBS 0.006347f
C553 B.n513 VSUBS 0.006347f
C554 B.n514 VSUBS 0.006347f
C555 B.n515 VSUBS 0.006347f
C556 B.n516 VSUBS 0.006347f
C557 B.n517 VSUBS 0.006347f
C558 B.n518 VSUBS 0.006347f
C559 B.n519 VSUBS 0.006347f
C560 B.n520 VSUBS 0.006347f
C561 B.n521 VSUBS 0.006347f
C562 B.n522 VSUBS 0.006347f
C563 B.n523 VSUBS 0.006347f
C564 B.n524 VSUBS 0.006347f
C565 B.n525 VSUBS 0.006347f
C566 B.n526 VSUBS 0.006347f
C567 B.n527 VSUBS 0.006347f
C568 B.n528 VSUBS 0.006347f
C569 B.n529 VSUBS 0.006347f
C570 B.n530 VSUBS 0.006347f
C571 B.n531 VSUBS 0.006347f
C572 B.n532 VSUBS 0.006347f
C573 B.n533 VSUBS 0.006347f
C574 B.n534 VSUBS 0.006347f
C575 B.n535 VSUBS 0.006347f
C576 B.n536 VSUBS 0.006347f
C577 B.n537 VSUBS 0.006347f
C578 B.n538 VSUBS 0.006347f
C579 B.n539 VSUBS 0.006347f
C580 B.n540 VSUBS 0.006347f
C581 B.n541 VSUBS 0.006347f
C582 B.n542 VSUBS 0.006347f
C583 B.n543 VSUBS 0.006347f
C584 B.n544 VSUBS 0.006347f
C585 B.n545 VSUBS 0.006347f
C586 B.n546 VSUBS 0.006347f
C587 B.n547 VSUBS 0.006347f
C588 B.n548 VSUBS 0.006347f
C589 B.n549 VSUBS 0.006347f
C590 B.n550 VSUBS 0.006347f
C591 B.n551 VSUBS 0.006347f
C592 B.n552 VSUBS 0.006347f
C593 B.n553 VSUBS 0.006347f
C594 B.n554 VSUBS 0.006347f
C595 B.n555 VSUBS 0.006347f
C596 B.n556 VSUBS 0.006347f
C597 B.n557 VSUBS 0.006347f
C598 B.n558 VSUBS 0.006347f
C599 B.n559 VSUBS 0.006347f
C600 B.n560 VSUBS 0.006347f
C601 B.n561 VSUBS 0.006347f
C602 B.n562 VSUBS 0.006347f
C603 B.n563 VSUBS 0.006347f
C604 B.n564 VSUBS 0.006347f
C605 B.n565 VSUBS 0.006347f
C606 B.n566 VSUBS 0.006347f
C607 B.n567 VSUBS 0.006347f
C608 B.n568 VSUBS 0.006347f
C609 B.n569 VSUBS 0.006347f
C610 B.n570 VSUBS 0.006347f
C611 B.n571 VSUBS 0.006347f
C612 B.n572 VSUBS 0.006347f
C613 B.n573 VSUBS 0.006347f
C614 B.n574 VSUBS 0.006347f
C615 B.n575 VSUBS 0.006347f
C616 B.n576 VSUBS 0.006347f
C617 B.n577 VSUBS 0.006347f
C618 B.n578 VSUBS 0.006347f
C619 B.n579 VSUBS 0.006347f
C620 B.n580 VSUBS 0.006347f
C621 B.n581 VSUBS 0.006347f
C622 B.n582 VSUBS 0.006347f
C623 B.n583 VSUBS 0.006347f
C624 B.n584 VSUBS 0.014875f
C625 B.n585 VSUBS 0.015181f
C626 B.n586 VSUBS 0.014444f
C627 B.n587 VSUBS 0.006347f
C628 B.n588 VSUBS 0.006347f
C629 B.n589 VSUBS 0.006347f
C630 B.n590 VSUBS 0.006347f
C631 B.n591 VSUBS 0.006347f
C632 B.n592 VSUBS 0.006347f
C633 B.n593 VSUBS 0.006347f
C634 B.n594 VSUBS 0.006347f
C635 B.n595 VSUBS 0.006347f
C636 B.n596 VSUBS 0.006347f
C637 B.n597 VSUBS 0.006347f
C638 B.n598 VSUBS 0.006347f
C639 B.n599 VSUBS 0.006347f
C640 B.n600 VSUBS 0.006347f
C641 B.n601 VSUBS 0.006347f
C642 B.n602 VSUBS 0.006347f
C643 B.n603 VSUBS 0.006347f
C644 B.n604 VSUBS 0.006347f
C645 B.n605 VSUBS 0.006347f
C646 B.n606 VSUBS 0.006347f
C647 B.n607 VSUBS 0.006347f
C648 B.n608 VSUBS 0.006347f
C649 B.n609 VSUBS 0.006347f
C650 B.n610 VSUBS 0.006347f
C651 B.n611 VSUBS 0.006347f
C652 B.n612 VSUBS 0.006347f
C653 B.n613 VSUBS 0.006347f
C654 B.n614 VSUBS 0.006347f
C655 B.n615 VSUBS 0.006347f
C656 B.n616 VSUBS 0.006347f
C657 B.n617 VSUBS 0.006347f
C658 B.n618 VSUBS 0.006347f
C659 B.n619 VSUBS 0.006347f
C660 B.n620 VSUBS 0.006347f
C661 B.n621 VSUBS 0.006347f
C662 B.n622 VSUBS 0.006347f
C663 B.n623 VSUBS 0.006347f
C664 B.n624 VSUBS 0.006347f
C665 B.n625 VSUBS 0.006347f
C666 B.n626 VSUBS 0.006347f
C667 B.n627 VSUBS 0.006347f
C668 B.n628 VSUBS 0.006347f
C669 B.n629 VSUBS 0.006347f
C670 B.n630 VSUBS 0.006347f
C671 B.n631 VSUBS 0.006347f
C672 B.n632 VSUBS 0.006347f
C673 B.n633 VSUBS 0.006347f
C674 B.n634 VSUBS 0.006347f
C675 B.n635 VSUBS 0.006347f
C676 B.n636 VSUBS 0.006347f
C677 B.n637 VSUBS 0.006347f
C678 B.n638 VSUBS 0.006347f
C679 B.n639 VSUBS 0.006347f
C680 B.n640 VSUBS 0.006347f
C681 B.n641 VSUBS 0.006347f
C682 B.n642 VSUBS 0.006347f
C683 B.n643 VSUBS 0.006347f
C684 B.n644 VSUBS 0.006347f
C685 B.n645 VSUBS 0.006347f
C686 B.n646 VSUBS 0.006347f
C687 B.n647 VSUBS 0.006347f
C688 B.n648 VSUBS 0.006347f
C689 B.n649 VSUBS 0.006347f
C690 B.n650 VSUBS 0.006347f
C691 B.n651 VSUBS 0.006347f
C692 B.n652 VSUBS 0.006347f
C693 B.n653 VSUBS 0.006347f
C694 B.n654 VSUBS 0.006347f
C695 B.n655 VSUBS 0.006347f
C696 B.n656 VSUBS 0.006347f
C697 B.n657 VSUBS 0.006347f
C698 B.n658 VSUBS 0.006347f
C699 B.n659 VSUBS 0.006347f
C700 B.n660 VSUBS 0.006347f
C701 B.n661 VSUBS 0.006347f
C702 B.n662 VSUBS 0.006347f
C703 B.n663 VSUBS 0.006347f
C704 B.n664 VSUBS 0.006347f
C705 B.n665 VSUBS 0.004387f
C706 B.n666 VSUBS 0.014706f
C707 B.n667 VSUBS 0.005134f
C708 B.n668 VSUBS 0.006347f
C709 B.n669 VSUBS 0.006347f
C710 B.n670 VSUBS 0.006347f
C711 B.n671 VSUBS 0.006347f
C712 B.n672 VSUBS 0.006347f
C713 B.n673 VSUBS 0.006347f
C714 B.n674 VSUBS 0.006347f
C715 B.n675 VSUBS 0.006347f
C716 B.n676 VSUBS 0.006347f
C717 B.n677 VSUBS 0.006347f
C718 B.n678 VSUBS 0.006347f
C719 B.n679 VSUBS 0.005134f
C720 B.n680 VSUBS 0.006347f
C721 B.n681 VSUBS 0.006347f
C722 B.n682 VSUBS 0.006347f
C723 B.n683 VSUBS 0.006347f
C724 B.n684 VSUBS 0.006347f
C725 B.n685 VSUBS 0.006347f
C726 B.n686 VSUBS 0.006347f
C727 B.n687 VSUBS 0.006347f
C728 B.n688 VSUBS 0.006347f
C729 B.n689 VSUBS 0.006347f
C730 B.n690 VSUBS 0.006347f
C731 B.n691 VSUBS 0.006347f
C732 B.n692 VSUBS 0.006347f
C733 B.n693 VSUBS 0.006347f
C734 B.n694 VSUBS 0.006347f
C735 B.n695 VSUBS 0.006347f
C736 B.n696 VSUBS 0.006347f
C737 B.n697 VSUBS 0.006347f
C738 B.n698 VSUBS 0.006347f
C739 B.n699 VSUBS 0.006347f
C740 B.n700 VSUBS 0.006347f
C741 B.n701 VSUBS 0.006347f
C742 B.n702 VSUBS 0.006347f
C743 B.n703 VSUBS 0.006347f
C744 B.n704 VSUBS 0.006347f
C745 B.n705 VSUBS 0.006347f
C746 B.n706 VSUBS 0.006347f
C747 B.n707 VSUBS 0.006347f
C748 B.n708 VSUBS 0.006347f
C749 B.n709 VSUBS 0.006347f
C750 B.n710 VSUBS 0.006347f
C751 B.n711 VSUBS 0.006347f
C752 B.n712 VSUBS 0.006347f
C753 B.n713 VSUBS 0.006347f
C754 B.n714 VSUBS 0.006347f
C755 B.n715 VSUBS 0.006347f
C756 B.n716 VSUBS 0.006347f
C757 B.n717 VSUBS 0.006347f
C758 B.n718 VSUBS 0.006347f
C759 B.n719 VSUBS 0.006347f
C760 B.n720 VSUBS 0.006347f
C761 B.n721 VSUBS 0.006347f
C762 B.n722 VSUBS 0.006347f
C763 B.n723 VSUBS 0.006347f
C764 B.n724 VSUBS 0.006347f
C765 B.n725 VSUBS 0.006347f
C766 B.n726 VSUBS 0.006347f
C767 B.n727 VSUBS 0.006347f
C768 B.n728 VSUBS 0.006347f
C769 B.n729 VSUBS 0.006347f
C770 B.n730 VSUBS 0.006347f
C771 B.n731 VSUBS 0.006347f
C772 B.n732 VSUBS 0.006347f
C773 B.n733 VSUBS 0.006347f
C774 B.n734 VSUBS 0.006347f
C775 B.n735 VSUBS 0.006347f
C776 B.n736 VSUBS 0.006347f
C777 B.n737 VSUBS 0.006347f
C778 B.n738 VSUBS 0.006347f
C779 B.n739 VSUBS 0.006347f
C780 B.n740 VSUBS 0.006347f
C781 B.n741 VSUBS 0.006347f
C782 B.n742 VSUBS 0.006347f
C783 B.n743 VSUBS 0.006347f
C784 B.n744 VSUBS 0.006347f
C785 B.n745 VSUBS 0.006347f
C786 B.n746 VSUBS 0.006347f
C787 B.n747 VSUBS 0.006347f
C788 B.n748 VSUBS 0.006347f
C789 B.n749 VSUBS 0.006347f
C790 B.n750 VSUBS 0.006347f
C791 B.n751 VSUBS 0.006347f
C792 B.n752 VSUBS 0.006347f
C793 B.n753 VSUBS 0.006347f
C794 B.n754 VSUBS 0.006347f
C795 B.n755 VSUBS 0.006347f
C796 B.n756 VSUBS 0.006347f
C797 B.n757 VSUBS 0.006347f
C798 B.n758 VSUBS 0.006347f
C799 B.n759 VSUBS 0.006347f
C800 B.n760 VSUBS 0.015181f
C801 B.n761 VSUBS 0.015181f
C802 B.n762 VSUBS 0.014875f
C803 B.n763 VSUBS 0.006347f
C804 B.n764 VSUBS 0.006347f
C805 B.n765 VSUBS 0.006347f
C806 B.n766 VSUBS 0.006347f
C807 B.n767 VSUBS 0.006347f
C808 B.n768 VSUBS 0.006347f
C809 B.n769 VSUBS 0.006347f
C810 B.n770 VSUBS 0.006347f
C811 B.n771 VSUBS 0.006347f
C812 B.n772 VSUBS 0.006347f
C813 B.n773 VSUBS 0.006347f
C814 B.n774 VSUBS 0.006347f
C815 B.n775 VSUBS 0.006347f
C816 B.n776 VSUBS 0.006347f
C817 B.n777 VSUBS 0.006347f
C818 B.n778 VSUBS 0.006347f
C819 B.n779 VSUBS 0.006347f
C820 B.n780 VSUBS 0.006347f
C821 B.n781 VSUBS 0.006347f
C822 B.n782 VSUBS 0.006347f
C823 B.n783 VSUBS 0.006347f
C824 B.n784 VSUBS 0.006347f
C825 B.n785 VSUBS 0.006347f
C826 B.n786 VSUBS 0.006347f
C827 B.n787 VSUBS 0.006347f
C828 B.n788 VSUBS 0.006347f
C829 B.n789 VSUBS 0.006347f
C830 B.n790 VSUBS 0.006347f
C831 B.n791 VSUBS 0.006347f
C832 B.n792 VSUBS 0.006347f
C833 B.n793 VSUBS 0.006347f
C834 B.n794 VSUBS 0.006347f
C835 B.n795 VSUBS 0.006347f
C836 B.n796 VSUBS 0.006347f
C837 B.n797 VSUBS 0.006347f
C838 B.n798 VSUBS 0.006347f
C839 B.n799 VSUBS 0.006347f
C840 B.n800 VSUBS 0.006347f
C841 B.n801 VSUBS 0.006347f
C842 B.n802 VSUBS 0.006347f
C843 B.n803 VSUBS 0.006347f
C844 B.n804 VSUBS 0.006347f
C845 B.n805 VSUBS 0.006347f
C846 B.n806 VSUBS 0.006347f
C847 B.n807 VSUBS 0.006347f
C848 B.n808 VSUBS 0.006347f
C849 B.n809 VSUBS 0.006347f
C850 B.n810 VSUBS 0.006347f
C851 B.n811 VSUBS 0.006347f
C852 B.n812 VSUBS 0.006347f
C853 B.n813 VSUBS 0.006347f
C854 B.n814 VSUBS 0.006347f
C855 B.n815 VSUBS 0.006347f
C856 B.n816 VSUBS 0.006347f
C857 B.n817 VSUBS 0.006347f
C858 B.n818 VSUBS 0.006347f
C859 B.n819 VSUBS 0.006347f
C860 B.n820 VSUBS 0.006347f
C861 B.n821 VSUBS 0.006347f
C862 B.n822 VSUBS 0.006347f
C863 B.n823 VSUBS 0.006347f
C864 B.n824 VSUBS 0.006347f
C865 B.n825 VSUBS 0.006347f
C866 B.n826 VSUBS 0.006347f
C867 B.n827 VSUBS 0.014372f
C868 VDD2.t0 VSUBS 0.341772f
C869 VDD2.t3 VSUBS 0.341772f
C870 VDD2.n0 VSUBS 3.73294f
C871 VDD2.t1 VSUBS 0.341772f
C872 VDD2.t2 VSUBS 0.341772f
C873 VDD2.n1 VSUBS 2.80937f
C874 VDD2.n2 VSUBS 4.9923f
C875 VN.t0 VSUBS 4.41749f
C876 VN.t3 VSUBS 4.43078f
C877 VN.n0 VSUBS 2.66955f
C878 VN.t1 VSUBS 4.43078f
C879 VN.t2 VSUBS 4.41749f
C880 VN.n1 VSUBS 4.42405f
C881 VTAIL.n0 VSUBS 0.025204f
C882 VTAIL.n1 VSUBS 0.023206f
C883 VTAIL.n2 VSUBS 0.01247f
C884 VTAIL.n3 VSUBS 0.029474f
C885 VTAIL.n4 VSUBS 0.013203f
C886 VTAIL.n5 VSUBS 0.023206f
C887 VTAIL.n6 VSUBS 0.012836f
C888 VTAIL.n7 VSUBS 0.029474f
C889 VTAIL.n8 VSUBS 0.013203f
C890 VTAIL.n9 VSUBS 0.023206f
C891 VTAIL.n10 VSUBS 0.01247f
C892 VTAIL.n11 VSUBS 0.029474f
C893 VTAIL.n12 VSUBS 0.013203f
C894 VTAIL.n13 VSUBS 0.023206f
C895 VTAIL.n14 VSUBS 0.01247f
C896 VTAIL.n15 VSUBS 0.029474f
C897 VTAIL.n16 VSUBS 0.013203f
C898 VTAIL.n17 VSUBS 0.023206f
C899 VTAIL.n18 VSUBS 0.01247f
C900 VTAIL.n19 VSUBS 0.029474f
C901 VTAIL.n20 VSUBS 0.013203f
C902 VTAIL.n21 VSUBS 0.023206f
C903 VTAIL.n22 VSUBS 0.01247f
C904 VTAIL.n23 VSUBS 0.029474f
C905 VTAIL.n24 VSUBS 0.013203f
C906 VTAIL.n25 VSUBS 0.023206f
C907 VTAIL.n26 VSUBS 0.01247f
C908 VTAIL.n27 VSUBS 0.022105f
C909 VTAIL.n28 VSUBS 0.01875f
C910 VTAIL.t0 VSUBS 0.063165f
C911 VTAIL.n29 VSUBS 0.171656f
C912 VTAIL.n30 VSUBS 1.60603f
C913 VTAIL.n31 VSUBS 0.01247f
C914 VTAIL.n32 VSUBS 0.013203f
C915 VTAIL.n33 VSUBS 0.029474f
C916 VTAIL.n34 VSUBS 0.029474f
C917 VTAIL.n35 VSUBS 0.013203f
C918 VTAIL.n36 VSUBS 0.01247f
C919 VTAIL.n37 VSUBS 0.023206f
C920 VTAIL.n38 VSUBS 0.023206f
C921 VTAIL.n39 VSUBS 0.01247f
C922 VTAIL.n40 VSUBS 0.013203f
C923 VTAIL.n41 VSUBS 0.029474f
C924 VTAIL.n42 VSUBS 0.029474f
C925 VTAIL.n43 VSUBS 0.013203f
C926 VTAIL.n44 VSUBS 0.01247f
C927 VTAIL.n45 VSUBS 0.023206f
C928 VTAIL.n46 VSUBS 0.023206f
C929 VTAIL.n47 VSUBS 0.01247f
C930 VTAIL.n48 VSUBS 0.013203f
C931 VTAIL.n49 VSUBS 0.029474f
C932 VTAIL.n50 VSUBS 0.029474f
C933 VTAIL.n51 VSUBS 0.013203f
C934 VTAIL.n52 VSUBS 0.01247f
C935 VTAIL.n53 VSUBS 0.023206f
C936 VTAIL.n54 VSUBS 0.023206f
C937 VTAIL.n55 VSUBS 0.01247f
C938 VTAIL.n56 VSUBS 0.013203f
C939 VTAIL.n57 VSUBS 0.029474f
C940 VTAIL.n58 VSUBS 0.029474f
C941 VTAIL.n59 VSUBS 0.013203f
C942 VTAIL.n60 VSUBS 0.01247f
C943 VTAIL.n61 VSUBS 0.023206f
C944 VTAIL.n62 VSUBS 0.023206f
C945 VTAIL.n63 VSUBS 0.01247f
C946 VTAIL.n64 VSUBS 0.013203f
C947 VTAIL.n65 VSUBS 0.029474f
C948 VTAIL.n66 VSUBS 0.029474f
C949 VTAIL.n67 VSUBS 0.013203f
C950 VTAIL.n68 VSUBS 0.01247f
C951 VTAIL.n69 VSUBS 0.023206f
C952 VTAIL.n70 VSUBS 0.023206f
C953 VTAIL.n71 VSUBS 0.01247f
C954 VTAIL.n72 VSUBS 0.01247f
C955 VTAIL.n73 VSUBS 0.013203f
C956 VTAIL.n74 VSUBS 0.029474f
C957 VTAIL.n75 VSUBS 0.029474f
C958 VTAIL.n76 VSUBS 0.029474f
C959 VTAIL.n77 VSUBS 0.012836f
C960 VTAIL.n78 VSUBS 0.01247f
C961 VTAIL.n79 VSUBS 0.023206f
C962 VTAIL.n80 VSUBS 0.023206f
C963 VTAIL.n81 VSUBS 0.01247f
C964 VTAIL.n82 VSUBS 0.013203f
C965 VTAIL.n83 VSUBS 0.029474f
C966 VTAIL.n84 VSUBS 0.070352f
C967 VTAIL.n85 VSUBS 0.013203f
C968 VTAIL.n86 VSUBS 0.01247f
C969 VTAIL.n87 VSUBS 0.056809f
C970 VTAIL.n88 VSUBS 0.03543f
C971 VTAIL.n89 VSUBS 0.188079f
C972 VTAIL.n90 VSUBS 0.025204f
C973 VTAIL.n91 VSUBS 0.023206f
C974 VTAIL.n92 VSUBS 0.01247f
C975 VTAIL.n93 VSUBS 0.029474f
C976 VTAIL.n94 VSUBS 0.013203f
C977 VTAIL.n95 VSUBS 0.023206f
C978 VTAIL.n96 VSUBS 0.012836f
C979 VTAIL.n97 VSUBS 0.029474f
C980 VTAIL.n98 VSUBS 0.013203f
C981 VTAIL.n99 VSUBS 0.023206f
C982 VTAIL.n100 VSUBS 0.01247f
C983 VTAIL.n101 VSUBS 0.029474f
C984 VTAIL.n102 VSUBS 0.013203f
C985 VTAIL.n103 VSUBS 0.023206f
C986 VTAIL.n104 VSUBS 0.01247f
C987 VTAIL.n105 VSUBS 0.029474f
C988 VTAIL.n106 VSUBS 0.013203f
C989 VTAIL.n107 VSUBS 0.023206f
C990 VTAIL.n108 VSUBS 0.01247f
C991 VTAIL.n109 VSUBS 0.029474f
C992 VTAIL.n110 VSUBS 0.013203f
C993 VTAIL.n111 VSUBS 0.023206f
C994 VTAIL.n112 VSUBS 0.01247f
C995 VTAIL.n113 VSUBS 0.029474f
C996 VTAIL.n114 VSUBS 0.013203f
C997 VTAIL.n115 VSUBS 0.023206f
C998 VTAIL.n116 VSUBS 0.01247f
C999 VTAIL.n117 VSUBS 0.022105f
C1000 VTAIL.n118 VSUBS 0.01875f
C1001 VTAIL.t6 VSUBS 0.063165f
C1002 VTAIL.n119 VSUBS 0.171656f
C1003 VTAIL.n120 VSUBS 1.60603f
C1004 VTAIL.n121 VSUBS 0.01247f
C1005 VTAIL.n122 VSUBS 0.013203f
C1006 VTAIL.n123 VSUBS 0.029474f
C1007 VTAIL.n124 VSUBS 0.029474f
C1008 VTAIL.n125 VSUBS 0.013203f
C1009 VTAIL.n126 VSUBS 0.01247f
C1010 VTAIL.n127 VSUBS 0.023206f
C1011 VTAIL.n128 VSUBS 0.023206f
C1012 VTAIL.n129 VSUBS 0.01247f
C1013 VTAIL.n130 VSUBS 0.013203f
C1014 VTAIL.n131 VSUBS 0.029474f
C1015 VTAIL.n132 VSUBS 0.029474f
C1016 VTAIL.n133 VSUBS 0.013203f
C1017 VTAIL.n134 VSUBS 0.01247f
C1018 VTAIL.n135 VSUBS 0.023206f
C1019 VTAIL.n136 VSUBS 0.023206f
C1020 VTAIL.n137 VSUBS 0.01247f
C1021 VTAIL.n138 VSUBS 0.013203f
C1022 VTAIL.n139 VSUBS 0.029474f
C1023 VTAIL.n140 VSUBS 0.029474f
C1024 VTAIL.n141 VSUBS 0.013203f
C1025 VTAIL.n142 VSUBS 0.01247f
C1026 VTAIL.n143 VSUBS 0.023206f
C1027 VTAIL.n144 VSUBS 0.023206f
C1028 VTAIL.n145 VSUBS 0.01247f
C1029 VTAIL.n146 VSUBS 0.013203f
C1030 VTAIL.n147 VSUBS 0.029474f
C1031 VTAIL.n148 VSUBS 0.029474f
C1032 VTAIL.n149 VSUBS 0.013203f
C1033 VTAIL.n150 VSUBS 0.01247f
C1034 VTAIL.n151 VSUBS 0.023206f
C1035 VTAIL.n152 VSUBS 0.023206f
C1036 VTAIL.n153 VSUBS 0.01247f
C1037 VTAIL.n154 VSUBS 0.013203f
C1038 VTAIL.n155 VSUBS 0.029474f
C1039 VTAIL.n156 VSUBS 0.029474f
C1040 VTAIL.n157 VSUBS 0.013203f
C1041 VTAIL.n158 VSUBS 0.01247f
C1042 VTAIL.n159 VSUBS 0.023206f
C1043 VTAIL.n160 VSUBS 0.023206f
C1044 VTAIL.n161 VSUBS 0.01247f
C1045 VTAIL.n162 VSUBS 0.01247f
C1046 VTAIL.n163 VSUBS 0.013203f
C1047 VTAIL.n164 VSUBS 0.029474f
C1048 VTAIL.n165 VSUBS 0.029474f
C1049 VTAIL.n166 VSUBS 0.029474f
C1050 VTAIL.n167 VSUBS 0.012836f
C1051 VTAIL.n168 VSUBS 0.01247f
C1052 VTAIL.n169 VSUBS 0.023206f
C1053 VTAIL.n170 VSUBS 0.023206f
C1054 VTAIL.n171 VSUBS 0.01247f
C1055 VTAIL.n172 VSUBS 0.013203f
C1056 VTAIL.n173 VSUBS 0.029474f
C1057 VTAIL.n174 VSUBS 0.070352f
C1058 VTAIL.n175 VSUBS 0.013203f
C1059 VTAIL.n176 VSUBS 0.01247f
C1060 VTAIL.n177 VSUBS 0.056809f
C1061 VTAIL.n178 VSUBS 0.03543f
C1062 VTAIL.n179 VSUBS 0.310714f
C1063 VTAIL.n180 VSUBS 0.025204f
C1064 VTAIL.n181 VSUBS 0.023206f
C1065 VTAIL.n182 VSUBS 0.01247f
C1066 VTAIL.n183 VSUBS 0.029474f
C1067 VTAIL.n184 VSUBS 0.013203f
C1068 VTAIL.n185 VSUBS 0.023206f
C1069 VTAIL.n186 VSUBS 0.012836f
C1070 VTAIL.n187 VSUBS 0.029474f
C1071 VTAIL.n188 VSUBS 0.013203f
C1072 VTAIL.n189 VSUBS 0.023206f
C1073 VTAIL.n190 VSUBS 0.01247f
C1074 VTAIL.n191 VSUBS 0.029474f
C1075 VTAIL.n192 VSUBS 0.013203f
C1076 VTAIL.n193 VSUBS 0.023206f
C1077 VTAIL.n194 VSUBS 0.01247f
C1078 VTAIL.n195 VSUBS 0.029474f
C1079 VTAIL.n196 VSUBS 0.013203f
C1080 VTAIL.n197 VSUBS 0.023206f
C1081 VTAIL.n198 VSUBS 0.01247f
C1082 VTAIL.n199 VSUBS 0.029474f
C1083 VTAIL.n200 VSUBS 0.013203f
C1084 VTAIL.n201 VSUBS 0.023206f
C1085 VTAIL.n202 VSUBS 0.01247f
C1086 VTAIL.n203 VSUBS 0.029474f
C1087 VTAIL.n204 VSUBS 0.013203f
C1088 VTAIL.n205 VSUBS 0.023206f
C1089 VTAIL.n206 VSUBS 0.01247f
C1090 VTAIL.n207 VSUBS 0.022105f
C1091 VTAIL.n208 VSUBS 0.01875f
C1092 VTAIL.t4 VSUBS 0.063165f
C1093 VTAIL.n209 VSUBS 0.171656f
C1094 VTAIL.n210 VSUBS 1.60603f
C1095 VTAIL.n211 VSUBS 0.01247f
C1096 VTAIL.n212 VSUBS 0.013203f
C1097 VTAIL.n213 VSUBS 0.029474f
C1098 VTAIL.n214 VSUBS 0.029474f
C1099 VTAIL.n215 VSUBS 0.013203f
C1100 VTAIL.n216 VSUBS 0.01247f
C1101 VTAIL.n217 VSUBS 0.023206f
C1102 VTAIL.n218 VSUBS 0.023206f
C1103 VTAIL.n219 VSUBS 0.01247f
C1104 VTAIL.n220 VSUBS 0.013203f
C1105 VTAIL.n221 VSUBS 0.029474f
C1106 VTAIL.n222 VSUBS 0.029474f
C1107 VTAIL.n223 VSUBS 0.013203f
C1108 VTAIL.n224 VSUBS 0.01247f
C1109 VTAIL.n225 VSUBS 0.023206f
C1110 VTAIL.n226 VSUBS 0.023206f
C1111 VTAIL.n227 VSUBS 0.01247f
C1112 VTAIL.n228 VSUBS 0.013203f
C1113 VTAIL.n229 VSUBS 0.029474f
C1114 VTAIL.n230 VSUBS 0.029474f
C1115 VTAIL.n231 VSUBS 0.013203f
C1116 VTAIL.n232 VSUBS 0.01247f
C1117 VTAIL.n233 VSUBS 0.023206f
C1118 VTAIL.n234 VSUBS 0.023206f
C1119 VTAIL.n235 VSUBS 0.01247f
C1120 VTAIL.n236 VSUBS 0.013203f
C1121 VTAIL.n237 VSUBS 0.029474f
C1122 VTAIL.n238 VSUBS 0.029474f
C1123 VTAIL.n239 VSUBS 0.013203f
C1124 VTAIL.n240 VSUBS 0.01247f
C1125 VTAIL.n241 VSUBS 0.023206f
C1126 VTAIL.n242 VSUBS 0.023206f
C1127 VTAIL.n243 VSUBS 0.01247f
C1128 VTAIL.n244 VSUBS 0.013203f
C1129 VTAIL.n245 VSUBS 0.029474f
C1130 VTAIL.n246 VSUBS 0.029474f
C1131 VTAIL.n247 VSUBS 0.013203f
C1132 VTAIL.n248 VSUBS 0.01247f
C1133 VTAIL.n249 VSUBS 0.023206f
C1134 VTAIL.n250 VSUBS 0.023206f
C1135 VTAIL.n251 VSUBS 0.01247f
C1136 VTAIL.n252 VSUBS 0.01247f
C1137 VTAIL.n253 VSUBS 0.013203f
C1138 VTAIL.n254 VSUBS 0.029474f
C1139 VTAIL.n255 VSUBS 0.029474f
C1140 VTAIL.n256 VSUBS 0.029474f
C1141 VTAIL.n257 VSUBS 0.012836f
C1142 VTAIL.n258 VSUBS 0.01247f
C1143 VTAIL.n259 VSUBS 0.023206f
C1144 VTAIL.n260 VSUBS 0.023206f
C1145 VTAIL.n261 VSUBS 0.01247f
C1146 VTAIL.n262 VSUBS 0.013203f
C1147 VTAIL.n263 VSUBS 0.029474f
C1148 VTAIL.n264 VSUBS 0.070352f
C1149 VTAIL.n265 VSUBS 0.013203f
C1150 VTAIL.n266 VSUBS 0.01247f
C1151 VTAIL.n267 VSUBS 0.056809f
C1152 VTAIL.n268 VSUBS 0.03543f
C1153 VTAIL.n269 VSUBS 1.88774f
C1154 VTAIL.n270 VSUBS 0.025204f
C1155 VTAIL.n271 VSUBS 0.023206f
C1156 VTAIL.n272 VSUBS 0.01247f
C1157 VTAIL.n273 VSUBS 0.029474f
C1158 VTAIL.n274 VSUBS 0.013203f
C1159 VTAIL.n275 VSUBS 0.023206f
C1160 VTAIL.n276 VSUBS 0.012836f
C1161 VTAIL.n277 VSUBS 0.029474f
C1162 VTAIL.n278 VSUBS 0.01247f
C1163 VTAIL.n279 VSUBS 0.013203f
C1164 VTAIL.n280 VSUBS 0.023206f
C1165 VTAIL.n281 VSUBS 0.01247f
C1166 VTAIL.n282 VSUBS 0.029474f
C1167 VTAIL.n283 VSUBS 0.013203f
C1168 VTAIL.n284 VSUBS 0.023206f
C1169 VTAIL.n285 VSUBS 0.01247f
C1170 VTAIL.n286 VSUBS 0.029474f
C1171 VTAIL.n287 VSUBS 0.013203f
C1172 VTAIL.n288 VSUBS 0.023206f
C1173 VTAIL.n289 VSUBS 0.01247f
C1174 VTAIL.n290 VSUBS 0.029474f
C1175 VTAIL.n291 VSUBS 0.013203f
C1176 VTAIL.n292 VSUBS 0.023206f
C1177 VTAIL.n293 VSUBS 0.01247f
C1178 VTAIL.n294 VSUBS 0.029474f
C1179 VTAIL.n295 VSUBS 0.013203f
C1180 VTAIL.n296 VSUBS 0.023206f
C1181 VTAIL.n297 VSUBS 0.01247f
C1182 VTAIL.n298 VSUBS 0.022105f
C1183 VTAIL.n299 VSUBS 0.01875f
C1184 VTAIL.t2 VSUBS 0.063165f
C1185 VTAIL.n300 VSUBS 0.171656f
C1186 VTAIL.n301 VSUBS 1.60603f
C1187 VTAIL.n302 VSUBS 0.01247f
C1188 VTAIL.n303 VSUBS 0.013203f
C1189 VTAIL.n304 VSUBS 0.029474f
C1190 VTAIL.n305 VSUBS 0.029474f
C1191 VTAIL.n306 VSUBS 0.013203f
C1192 VTAIL.n307 VSUBS 0.01247f
C1193 VTAIL.n308 VSUBS 0.023206f
C1194 VTAIL.n309 VSUBS 0.023206f
C1195 VTAIL.n310 VSUBS 0.01247f
C1196 VTAIL.n311 VSUBS 0.013203f
C1197 VTAIL.n312 VSUBS 0.029474f
C1198 VTAIL.n313 VSUBS 0.029474f
C1199 VTAIL.n314 VSUBS 0.013203f
C1200 VTAIL.n315 VSUBS 0.01247f
C1201 VTAIL.n316 VSUBS 0.023206f
C1202 VTAIL.n317 VSUBS 0.023206f
C1203 VTAIL.n318 VSUBS 0.01247f
C1204 VTAIL.n319 VSUBS 0.013203f
C1205 VTAIL.n320 VSUBS 0.029474f
C1206 VTAIL.n321 VSUBS 0.029474f
C1207 VTAIL.n322 VSUBS 0.013203f
C1208 VTAIL.n323 VSUBS 0.01247f
C1209 VTAIL.n324 VSUBS 0.023206f
C1210 VTAIL.n325 VSUBS 0.023206f
C1211 VTAIL.n326 VSUBS 0.01247f
C1212 VTAIL.n327 VSUBS 0.013203f
C1213 VTAIL.n328 VSUBS 0.029474f
C1214 VTAIL.n329 VSUBS 0.029474f
C1215 VTAIL.n330 VSUBS 0.013203f
C1216 VTAIL.n331 VSUBS 0.01247f
C1217 VTAIL.n332 VSUBS 0.023206f
C1218 VTAIL.n333 VSUBS 0.023206f
C1219 VTAIL.n334 VSUBS 0.01247f
C1220 VTAIL.n335 VSUBS 0.013203f
C1221 VTAIL.n336 VSUBS 0.029474f
C1222 VTAIL.n337 VSUBS 0.029474f
C1223 VTAIL.n338 VSUBS 0.013203f
C1224 VTAIL.n339 VSUBS 0.01247f
C1225 VTAIL.n340 VSUBS 0.023206f
C1226 VTAIL.n341 VSUBS 0.023206f
C1227 VTAIL.n342 VSUBS 0.01247f
C1228 VTAIL.n343 VSUBS 0.013203f
C1229 VTAIL.n344 VSUBS 0.029474f
C1230 VTAIL.n345 VSUBS 0.029474f
C1231 VTAIL.n346 VSUBS 0.029474f
C1232 VTAIL.n347 VSUBS 0.012836f
C1233 VTAIL.n348 VSUBS 0.01247f
C1234 VTAIL.n349 VSUBS 0.023206f
C1235 VTAIL.n350 VSUBS 0.023206f
C1236 VTAIL.n351 VSUBS 0.01247f
C1237 VTAIL.n352 VSUBS 0.013203f
C1238 VTAIL.n353 VSUBS 0.029474f
C1239 VTAIL.n354 VSUBS 0.070352f
C1240 VTAIL.n355 VSUBS 0.013203f
C1241 VTAIL.n356 VSUBS 0.01247f
C1242 VTAIL.n357 VSUBS 0.056809f
C1243 VTAIL.n358 VSUBS 0.03543f
C1244 VTAIL.n359 VSUBS 1.88774f
C1245 VTAIL.n360 VSUBS 0.025204f
C1246 VTAIL.n361 VSUBS 0.023206f
C1247 VTAIL.n362 VSUBS 0.01247f
C1248 VTAIL.n363 VSUBS 0.029474f
C1249 VTAIL.n364 VSUBS 0.013203f
C1250 VTAIL.n365 VSUBS 0.023206f
C1251 VTAIL.n366 VSUBS 0.012836f
C1252 VTAIL.n367 VSUBS 0.029474f
C1253 VTAIL.n368 VSUBS 0.01247f
C1254 VTAIL.n369 VSUBS 0.013203f
C1255 VTAIL.n370 VSUBS 0.023206f
C1256 VTAIL.n371 VSUBS 0.01247f
C1257 VTAIL.n372 VSUBS 0.029474f
C1258 VTAIL.n373 VSUBS 0.013203f
C1259 VTAIL.n374 VSUBS 0.023206f
C1260 VTAIL.n375 VSUBS 0.01247f
C1261 VTAIL.n376 VSUBS 0.029474f
C1262 VTAIL.n377 VSUBS 0.013203f
C1263 VTAIL.n378 VSUBS 0.023206f
C1264 VTAIL.n379 VSUBS 0.01247f
C1265 VTAIL.n380 VSUBS 0.029474f
C1266 VTAIL.n381 VSUBS 0.013203f
C1267 VTAIL.n382 VSUBS 0.023206f
C1268 VTAIL.n383 VSUBS 0.01247f
C1269 VTAIL.n384 VSUBS 0.029474f
C1270 VTAIL.n385 VSUBS 0.013203f
C1271 VTAIL.n386 VSUBS 0.023206f
C1272 VTAIL.n387 VSUBS 0.01247f
C1273 VTAIL.n388 VSUBS 0.022105f
C1274 VTAIL.n389 VSUBS 0.01875f
C1275 VTAIL.t1 VSUBS 0.063165f
C1276 VTAIL.n390 VSUBS 0.171656f
C1277 VTAIL.n391 VSUBS 1.60603f
C1278 VTAIL.n392 VSUBS 0.01247f
C1279 VTAIL.n393 VSUBS 0.013203f
C1280 VTAIL.n394 VSUBS 0.029474f
C1281 VTAIL.n395 VSUBS 0.029474f
C1282 VTAIL.n396 VSUBS 0.013203f
C1283 VTAIL.n397 VSUBS 0.01247f
C1284 VTAIL.n398 VSUBS 0.023206f
C1285 VTAIL.n399 VSUBS 0.023206f
C1286 VTAIL.n400 VSUBS 0.01247f
C1287 VTAIL.n401 VSUBS 0.013203f
C1288 VTAIL.n402 VSUBS 0.029474f
C1289 VTAIL.n403 VSUBS 0.029474f
C1290 VTAIL.n404 VSUBS 0.013203f
C1291 VTAIL.n405 VSUBS 0.01247f
C1292 VTAIL.n406 VSUBS 0.023206f
C1293 VTAIL.n407 VSUBS 0.023206f
C1294 VTAIL.n408 VSUBS 0.01247f
C1295 VTAIL.n409 VSUBS 0.013203f
C1296 VTAIL.n410 VSUBS 0.029474f
C1297 VTAIL.n411 VSUBS 0.029474f
C1298 VTAIL.n412 VSUBS 0.013203f
C1299 VTAIL.n413 VSUBS 0.01247f
C1300 VTAIL.n414 VSUBS 0.023206f
C1301 VTAIL.n415 VSUBS 0.023206f
C1302 VTAIL.n416 VSUBS 0.01247f
C1303 VTAIL.n417 VSUBS 0.013203f
C1304 VTAIL.n418 VSUBS 0.029474f
C1305 VTAIL.n419 VSUBS 0.029474f
C1306 VTAIL.n420 VSUBS 0.013203f
C1307 VTAIL.n421 VSUBS 0.01247f
C1308 VTAIL.n422 VSUBS 0.023206f
C1309 VTAIL.n423 VSUBS 0.023206f
C1310 VTAIL.n424 VSUBS 0.01247f
C1311 VTAIL.n425 VSUBS 0.013203f
C1312 VTAIL.n426 VSUBS 0.029474f
C1313 VTAIL.n427 VSUBS 0.029474f
C1314 VTAIL.n428 VSUBS 0.013203f
C1315 VTAIL.n429 VSUBS 0.01247f
C1316 VTAIL.n430 VSUBS 0.023206f
C1317 VTAIL.n431 VSUBS 0.023206f
C1318 VTAIL.n432 VSUBS 0.01247f
C1319 VTAIL.n433 VSUBS 0.013203f
C1320 VTAIL.n434 VSUBS 0.029474f
C1321 VTAIL.n435 VSUBS 0.029474f
C1322 VTAIL.n436 VSUBS 0.029474f
C1323 VTAIL.n437 VSUBS 0.012836f
C1324 VTAIL.n438 VSUBS 0.01247f
C1325 VTAIL.n439 VSUBS 0.023206f
C1326 VTAIL.n440 VSUBS 0.023206f
C1327 VTAIL.n441 VSUBS 0.01247f
C1328 VTAIL.n442 VSUBS 0.013203f
C1329 VTAIL.n443 VSUBS 0.029474f
C1330 VTAIL.n444 VSUBS 0.070352f
C1331 VTAIL.n445 VSUBS 0.013203f
C1332 VTAIL.n446 VSUBS 0.01247f
C1333 VTAIL.n447 VSUBS 0.056809f
C1334 VTAIL.n448 VSUBS 0.03543f
C1335 VTAIL.n449 VSUBS 0.310714f
C1336 VTAIL.n450 VSUBS 0.025204f
C1337 VTAIL.n451 VSUBS 0.023206f
C1338 VTAIL.n452 VSUBS 0.01247f
C1339 VTAIL.n453 VSUBS 0.029474f
C1340 VTAIL.n454 VSUBS 0.013203f
C1341 VTAIL.n455 VSUBS 0.023206f
C1342 VTAIL.n456 VSUBS 0.012836f
C1343 VTAIL.n457 VSUBS 0.029474f
C1344 VTAIL.n458 VSUBS 0.01247f
C1345 VTAIL.n459 VSUBS 0.013203f
C1346 VTAIL.n460 VSUBS 0.023206f
C1347 VTAIL.n461 VSUBS 0.01247f
C1348 VTAIL.n462 VSUBS 0.029474f
C1349 VTAIL.n463 VSUBS 0.013203f
C1350 VTAIL.n464 VSUBS 0.023206f
C1351 VTAIL.n465 VSUBS 0.01247f
C1352 VTAIL.n466 VSUBS 0.029474f
C1353 VTAIL.n467 VSUBS 0.013203f
C1354 VTAIL.n468 VSUBS 0.023206f
C1355 VTAIL.n469 VSUBS 0.01247f
C1356 VTAIL.n470 VSUBS 0.029474f
C1357 VTAIL.n471 VSUBS 0.013203f
C1358 VTAIL.n472 VSUBS 0.023206f
C1359 VTAIL.n473 VSUBS 0.01247f
C1360 VTAIL.n474 VSUBS 0.029474f
C1361 VTAIL.n475 VSUBS 0.013203f
C1362 VTAIL.n476 VSUBS 0.023206f
C1363 VTAIL.n477 VSUBS 0.01247f
C1364 VTAIL.n478 VSUBS 0.022105f
C1365 VTAIL.n479 VSUBS 0.01875f
C1366 VTAIL.t7 VSUBS 0.063165f
C1367 VTAIL.n480 VSUBS 0.171656f
C1368 VTAIL.n481 VSUBS 1.60603f
C1369 VTAIL.n482 VSUBS 0.01247f
C1370 VTAIL.n483 VSUBS 0.013203f
C1371 VTAIL.n484 VSUBS 0.029474f
C1372 VTAIL.n485 VSUBS 0.029474f
C1373 VTAIL.n486 VSUBS 0.013203f
C1374 VTAIL.n487 VSUBS 0.01247f
C1375 VTAIL.n488 VSUBS 0.023206f
C1376 VTAIL.n489 VSUBS 0.023206f
C1377 VTAIL.n490 VSUBS 0.01247f
C1378 VTAIL.n491 VSUBS 0.013203f
C1379 VTAIL.n492 VSUBS 0.029474f
C1380 VTAIL.n493 VSUBS 0.029474f
C1381 VTAIL.n494 VSUBS 0.013203f
C1382 VTAIL.n495 VSUBS 0.01247f
C1383 VTAIL.n496 VSUBS 0.023206f
C1384 VTAIL.n497 VSUBS 0.023206f
C1385 VTAIL.n498 VSUBS 0.01247f
C1386 VTAIL.n499 VSUBS 0.013203f
C1387 VTAIL.n500 VSUBS 0.029474f
C1388 VTAIL.n501 VSUBS 0.029474f
C1389 VTAIL.n502 VSUBS 0.013203f
C1390 VTAIL.n503 VSUBS 0.01247f
C1391 VTAIL.n504 VSUBS 0.023206f
C1392 VTAIL.n505 VSUBS 0.023206f
C1393 VTAIL.n506 VSUBS 0.01247f
C1394 VTAIL.n507 VSUBS 0.013203f
C1395 VTAIL.n508 VSUBS 0.029474f
C1396 VTAIL.n509 VSUBS 0.029474f
C1397 VTAIL.n510 VSUBS 0.013203f
C1398 VTAIL.n511 VSUBS 0.01247f
C1399 VTAIL.n512 VSUBS 0.023206f
C1400 VTAIL.n513 VSUBS 0.023206f
C1401 VTAIL.n514 VSUBS 0.01247f
C1402 VTAIL.n515 VSUBS 0.013203f
C1403 VTAIL.n516 VSUBS 0.029474f
C1404 VTAIL.n517 VSUBS 0.029474f
C1405 VTAIL.n518 VSUBS 0.013203f
C1406 VTAIL.n519 VSUBS 0.01247f
C1407 VTAIL.n520 VSUBS 0.023206f
C1408 VTAIL.n521 VSUBS 0.023206f
C1409 VTAIL.n522 VSUBS 0.01247f
C1410 VTAIL.n523 VSUBS 0.013203f
C1411 VTAIL.n524 VSUBS 0.029474f
C1412 VTAIL.n525 VSUBS 0.029474f
C1413 VTAIL.n526 VSUBS 0.029474f
C1414 VTAIL.n527 VSUBS 0.012836f
C1415 VTAIL.n528 VSUBS 0.01247f
C1416 VTAIL.n529 VSUBS 0.023206f
C1417 VTAIL.n530 VSUBS 0.023206f
C1418 VTAIL.n531 VSUBS 0.01247f
C1419 VTAIL.n532 VSUBS 0.013203f
C1420 VTAIL.n533 VSUBS 0.029474f
C1421 VTAIL.n534 VSUBS 0.070352f
C1422 VTAIL.n535 VSUBS 0.013203f
C1423 VTAIL.n536 VSUBS 0.01247f
C1424 VTAIL.n537 VSUBS 0.056809f
C1425 VTAIL.n538 VSUBS 0.03543f
C1426 VTAIL.n539 VSUBS 0.310714f
C1427 VTAIL.n540 VSUBS 0.025204f
C1428 VTAIL.n541 VSUBS 0.023206f
C1429 VTAIL.n542 VSUBS 0.01247f
C1430 VTAIL.n543 VSUBS 0.029474f
C1431 VTAIL.n544 VSUBS 0.013203f
C1432 VTAIL.n545 VSUBS 0.023206f
C1433 VTAIL.n546 VSUBS 0.012836f
C1434 VTAIL.n547 VSUBS 0.029474f
C1435 VTAIL.n548 VSUBS 0.01247f
C1436 VTAIL.n549 VSUBS 0.013203f
C1437 VTAIL.n550 VSUBS 0.023206f
C1438 VTAIL.n551 VSUBS 0.01247f
C1439 VTAIL.n552 VSUBS 0.029474f
C1440 VTAIL.n553 VSUBS 0.013203f
C1441 VTAIL.n554 VSUBS 0.023206f
C1442 VTAIL.n555 VSUBS 0.01247f
C1443 VTAIL.n556 VSUBS 0.029474f
C1444 VTAIL.n557 VSUBS 0.013203f
C1445 VTAIL.n558 VSUBS 0.023206f
C1446 VTAIL.n559 VSUBS 0.01247f
C1447 VTAIL.n560 VSUBS 0.029474f
C1448 VTAIL.n561 VSUBS 0.013203f
C1449 VTAIL.n562 VSUBS 0.023206f
C1450 VTAIL.n563 VSUBS 0.01247f
C1451 VTAIL.n564 VSUBS 0.029474f
C1452 VTAIL.n565 VSUBS 0.013203f
C1453 VTAIL.n566 VSUBS 0.023206f
C1454 VTAIL.n567 VSUBS 0.01247f
C1455 VTAIL.n568 VSUBS 0.022105f
C1456 VTAIL.n569 VSUBS 0.01875f
C1457 VTAIL.t5 VSUBS 0.063165f
C1458 VTAIL.n570 VSUBS 0.171656f
C1459 VTAIL.n571 VSUBS 1.60603f
C1460 VTAIL.n572 VSUBS 0.01247f
C1461 VTAIL.n573 VSUBS 0.013203f
C1462 VTAIL.n574 VSUBS 0.029474f
C1463 VTAIL.n575 VSUBS 0.029474f
C1464 VTAIL.n576 VSUBS 0.013203f
C1465 VTAIL.n577 VSUBS 0.01247f
C1466 VTAIL.n578 VSUBS 0.023206f
C1467 VTAIL.n579 VSUBS 0.023206f
C1468 VTAIL.n580 VSUBS 0.01247f
C1469 VTAIL.n581 VSUBS 0.013203f
C1470 VTAIL.n582 VSUBS 0.029474f
C1471 VTAIL.n583 VSUBS 0.029474f
C1472 VTAIL.n584 VSUBS 0.013203f
C1473 VTAIL.n585 VSUBS 0.01247f
C1474 VTAIL.n586 VSUBS 0.023206f
C1475 VTAIL.n587 VSUBS 0.023206f
C1476 VTAIL.n588 VSUBS 0.01247f
C1477 VTAIL.n589 VSUBS 0.013203f
C1478 VTAIL.n590 VSUBS 0.029474f
C1479 VTAIL.n591 VSUBS 0.029474f
C1480 VTAIL.n592 VSUBS 0.013203f
C1481 VTAIL.n593 VSUBS 0.01247f
C1482 VTAIL.n594 VSUBS 0.023206f
C1483 VTAIL.n595 VSUBS 0.023206f
C1484 VTAIL.n596 VSUBS 0.01247f
C1485 VTAIL.n597 VSUBS 0.013203f
C1486 VTAIL.n598 VSUBS 0.029474f
C1487 VTAIL.n599 VSUBS 0.029474f
C1488 VTAIL.n600 VSUBS 0.013203f
C1489 VTAIL.n601 VSUBS 0.01247f
C1490 VTAIL.n602 VSUBS 0.023206f
C1491 VTAIL.n603 VSUBS 0.023206f
C1492 VTAIL.n604 VSUBS 0.01247f
C1493 VTAIL.n605 VSUBS 0.013203f
C1494 VTAIL.n606 VSUBS 0.029474f
C1495 VTAIL.n607 VSUBS 0.029474f
C1496 VTAIL.n608 VSUBS 0.013203f
C1497 VTAIL.n609 VSUBS 0.01247f
C1498 VTAIL.n610 VSUBS 0.023206f
C1499 VTAIL.n611 VSUBS 0.023206f
C1500 VTAIL.n612 VSUBS 0.01247f
C1501 VTAIL.n613 VSUBS 0.013203f
C1502 VTAIL.n614 VSUBS 0.029474f
C1503 VTAIL.n615 VSUBS 0.029474f
C1504 VTAIL.n616 VSUBS 0.029474f
C1505 VTAIL.n617 VSUBS 0.012836f
C1506 VTAIL.n618 VSUBS 0.01247f
C1507 VTAIL.n619 VSUBS 0.023206f
C1508 VTAIL.n620 VSUBS 0.023206f
C1509 VTAIL.n621 VSUBS 0.01247f
C1510 VTAIL.n622 VSUBS 0.013203f
C1511 VTAIL.n623 VSUBS 0.029474f
C1512 VTAIL.n624 VSUBS 0.070352f
C1513 VTAIL.n625 VSUBS 0.013203f
C1514 VTAIL.n626 VSUBS 0.01247f
C1515 VTAIL.n627 VSUBS 0.056809f
C1516 VTAIL.n628 VSUBS 0.03543f
C1517 VTAIL.n629 VSUBS 1.88774f
C1518 VTAIL.n630 VSUBS 0.025204f
C1519 VTAIL.n631 VSUBS 0.023206f
C1520 VTAIL.n632 VSUBS 0.01247f
C1521 VTAIL.n633 VSUBS 0.029474f
C1522 VTAIL.n634 VSUBS 0.013203f
C1523 VTAIL.n635 VSUBS 0.023206f
C1524 VTAIL.n636 VSUBS 0.012836f
C1525 VTAIL.n637 VSUBS 0.029474f
C1526 VTAIL.n638 VSUBS 0.013203f
C1527 VTAIL.n639 VSUBS 0.023206f
C1528 VTAIL.n640 VSUBS 0.01247f
C1529 VTAIL.n641 VSUBS 0.029474f
C1530 VTAIL.n642 VSUBS 0.013203f
C1531 VTAIL.n643 VSUBS 0.023206f
C1532 VTAIL.n644 VSUBS 0.01247f
C1533 VTAIL.n645 VSUBS 0.029474f
C1534 VTAIL.n646 VSUBS 0.013203f
C1535 VTAIL.n647 VSUBS 0.023206f
C1536 VTAIL.n648 VSUBS 0.01247f
C1537 VTAIL.n649 VSUBS 0.029474f
C1538 VTAIL.n650 VSUBS 0.013203f
C1539 VTAIL.n651 VSUBS 0.023206f
C1540 VTAIL.n652 VSUBS 0.01247f
C1541 VTAIL.n653 VSUBS 0.029474f
C1542 VTAIL.n654 VSUBS 0.013203f
C1543 VTAIL.n655 VSUBS 0.023206f
C1544 VTAIL.n656 VSUBS 0.01247f
C1545 VTAIL.n657 VSUBS 0.022105f
C1546 VTAIL.n658 VSUBS 0.01875f
C1547 VTAIL.t3 VSUBS 0.063165f
C1548 VTAIL.n659 VSUBS 0.171656f
C1549 VTAIL.n660 VSUBS 1.60603f
C1550 VTAIL.n661 VSUBS 0.01247f
C1551 VTAIL.n662 VSUBS 0.013203f
C1552 VTAIL.n663 VSUBS 0.029474f
C1553 VTAIL.n664 VSUBS 0.029474f
C1554 VTAIL.n665 VSUBS 0.013203f
C1555 VTAIL.n666 VSUBS 0.01247f
C1556 VTAIL.n667 VSUBS 0.023206f
C1557 VTAIL.n668 VSUBS 0.023206f
C1558 VTAIL.n669 VSUBS 0.01247f
C1559 VTAIL.n670 VSUBS 0.013203f
C1560 VTAIL.n671 VSUBS 0.029474f
C1561 VTAIL.n672 VSUBS 0.029474f
C1562 VTAIL.n673 VSUBS 0.013203f
C1563 VTAIL.n674 VSUBS 0.01247f
C1564 VTAIL.n675 VSUBS 0.023206f
C1565 VTAIL.n676 VSUBS 0.023206f
C1566 VTAIL.n677 VSUBS 0.01247f
C1567 VTAIL.n678 VSUBS 0.013203f
C1568 VTAIL.n679 VSUBS 0.029474f
C1569 VTAIL.n680 VSUBS 0.029474f
C1570 VTAIL.n681 VSUBS 0.013203f
C1571 VTAIL.n682 VSUBS 0.01247f
C1572 VTAIL.n683 VSUBS 0.023206f
C1573 VTAIL.n684 VSUBS 0.023206f
C1574 VTAIL.n685 VSUBS 0.01247f
C1575 VTAIL.n686 VSUBS 0.013203f
C1576 VTAIL.n687 VSUBS 0.029474f
C1577 VTAIL.n688 VSUBS 0.029474f
C1578 VTAIL.n689 VSUBS 0.013203f
C1579 VTAIL.n690 VSUBS 0.01247f
C1580 VTAIL.n691 VSUBS 0.023206f
C1581 VTAIL.n692 VSUBS 0.023206f
C1582 VTAIL.n693 VSUBS 0.01247f
C1583 VTAIL.n694 VSUBS 0.013203f
C1584 VTAIL.n695 VSUBS 0.029474f
C1585 VTAIL.n696 VSUBS 0.029474f
C1586 VTAIL.n697 VSUBS 0.013203f
C1587 VTAIL.n698 VSUBS 0.01247f
C1588 VTAIL.n699 VSUBS 0.023206f
C1589 VTAIL.n700 VSUBS 0.023206f
C1590 VTAIL.n701 VSUBS 0.01247f
C1591 VTAIL.n702 VSUBS 0.01247f
C1592 VTAIL.n703 VSUBS 0.013203f
C1593 VTAIL.n704 VSUBS 0.029474f
C1594 VTAIL.n705 VSUBS 0.029474f
C1595 VTAIL.n706 VSUBS 0.029474f
C1596 VTAIL.n707 VSUBS 0.012836f
C1597 VTAIL.n708 VSUBS 0.01247f
C1598 VTAIL.n709 VSUBS 0.023206f
C1599 VTAIL.n710 VSUBS 0.023206f
C1600 VTAIL.n711 VSUBS 0.01247f
C1601 VTAIL.n712 VSUBS 0.013203f
C1602 VTAIL.n713 VSUBS 0.029474f
C1603 VTAIL.n714 VSUBS 0.070352f
C1604 VTAIL.n715 VSUBS 0.013203f
C1605 VTAIL.n716 VSUBS 0.01247f
C1606 VTAIL.n717 VSUBS 0.056809f
C1607 VTAIL.n718 VSUBS 0.03543f
C1608 VTAIL.n719 VSUBS 1.7564f
C1609 VDD1.t0 VSUBS 0.346945f
C1610 VDD1.t1 VSUBS 0.346945f
C1611 VDD1.n0 VSUBS 2.85256f
C1612 VDD1.t3 VSUBS 0.346945f
C1613 VDD1.t2 VSUBS 0.346945f
C1614 VDD1.n1 VSUBS 3.81696f
C1615 VP.t1 VSUBS 4.4693f
C1616 VP.n0 VSUBS 1.65786f
C1617 VP.n1 VSUBS 0.027878f
C1618 VP.n2 VSUBS 0.040524f
C1619 VP.n3 VSUBS 0.027878f
C1620 VP.n4 VSUBS 0.037404f
C1621 VP.t0 VSUBS 4.90193f
C1622 VP.t2 VSUBS 4.88724f
C1623 VP.n5 VSUBS 4.88348f
C1624 VP.t3 VSUBS 4.4693f
C1625 VP.n6 VSUBS 1.65786f
C1626 VP.n7 VSUBS 1.81648f
C1627 VP.n8 VSUBS 0.044987f
C1628 VP.n9 VSUBS 0.027878f
C1629 VP.n10 VSUBS 0.051696f
C1630 VP.n11 VSUBS 0.051696f
C1631 VP.n12 VSUBS 0.040524f
C1632 VP.n13 VSUBS 0.027878f
C1633 VP.n14 VSUBS 0.027878f
C1634 VP.n15 VSUBS 0.027878f
C1635 VP.n16 VSUBS 0.051696f
C1636 VP.n17 VSUBS 0.051696f
C1637 VP.n18 VSUBS 0.037404f
C1638 VP.n19 VSUBS 0.044987f
C1639 VP.n20 VSUBS 0.075437f
.ends

