* NGSPICE file created from diff_pair_sample_1329.ext - technology: sky130A

.subckt diff_pair_sample_1329 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t11 VP.t0 VDD1.t3 w_n3866_n4008# sky130_fd_pr__pfet_01v8 ad=2.508 pd=15.53 as=2.508 ps=15.53 w=15.2 l=3.29
X1 B.t11 B.t9 B.t10 w_n3866_n4008# sky130_fd_pr__pfet_01v8 ad=5.928 pd=31.18 as=0 ps=0 w=15.2 l=3.29
X2 B.t8 B.t6 B.t7 w_n3866_n4008# sky130_fd_pr__pfet_01v8 ad=5.928 pd=31.18 as=0 ps=0 w=15.2 l=3.29
X3 VTAIL.t2 VN.t0 VDD2.t5 w_n3866_n4008# sky130_fd_pr__pfet_01v8 ad=2.508 pd=15.53 as=2.508 ps=15.53 w=15.2 l=3.29
X4 VDD1.t5 VP.t1 VTAIL.t10 w_n3866_n4008# sky130_fd_pr__pfet_01v8 ad=5.928 pd=31.18 as=2.508 ps=15.53 w=15.2 l=3.29
X5 B.t5 B.t3 B.t4 w_n3866_n4008# sky130_fd_pr__pfet_01v8 ad=5.928 pd=31.18 as=0 ps=0 w=15.2 l=3.29
X6 B.t2 B.t0 B.t1 w_n3866_n4008# sky130_fd_pr__pfet_01v8 ad=5.928 pd=31.18 as=0 ps=0 w=15.2 l=3.29
X7 VDD1.t2 VP.t2 VTAIL.t9 w_n3866_n4008# sky130_fd_pr__pfet_01v8 ad=2.508 pd=15.53 as=5.928 ps=31.18 w=15.2 l=3.29
X8 VDD2.t4 VN.t1 VTAIL.t0 w_n3866_n4008# sky130_fd_pr__pfet_01v8 ad=2.508 pd=15.53 as=5.928 ps=31.18 w=15.2 l=3.29
X9 VTAIL.t1 VN.t2 VDD2.t3 w_n3866_n4008# sky130_fd_pr__pfet_01v8 ad=2.508 pd=15.53 as=2.508 ps=15.53 w=15.2 l=3.29
X10 VDD2.t2 VN.t3 VTAIL.t4 w_n3866_n4008# sky130_fd_pr__pfet_01v8 ad=5.928 pd=31.18 as=2.508 ps=15.53 w=15.2 l=3.29
X11 VDD1.t0 VP.t3 VTAIL.t8 w_n3866_n4008# sky130_fd_pr__pfet_01v8 ad=5.928 pd=31.18 as=2.508 ps=15.53 w=15.2 l=3.29
X12 VDD2.t1 VN.t4 VTAIL.t3 w_n3866_n4008# sky130_fd_pr__pfet_01v8 ad=5.928 pd=31.18 as=2.508 ps=15.53 w=15.2 l=3.29
X13 VDD1.t1 VP.t4 VTAIL.t7 w_n3866_n4008# sky130_fd_pr__pfet_01v8 ad=2.508 pd=15.53 as=5.928 ps=31.18 w=15.2 l=3.29
X14 VDD2.t0 VN.t5 VTAIL.t5 w_n3866_n4008# sky130_fd_pr__pfet_01v8 ad=2.508 pd=15.53 as=5.928 ps=31.18 w=15.2 l=3.29
X15 VTAIL.t6 VP.t5 VDD1.t4 w_n3866_n4008# sky130_fd_pr__pfet_01v8 ad=2.508 pd=15.53 as=2.508 ps=15.53 w=15.2 l=3.29
R0 VP.n16 VP.n15 161.3
R1 VP.n17 VP.n12 161.3
R2 VP.n19 VP.n18 161.3
R3 VP.n20 VP.n11 161.3
R4 VP.n22 VP.n21 161.3
R5 VP.n23 VP.n10 161.3
R6 VP.n25 VP.n24 161.3
R7 VP.n49 VP.n48 161.3
R8 VP.n47 VP.n1 161.3
R9 VP.n46 VP.n45 161.3
R10 VP.n44 VP.n2 161.3
R11 VP.n43 VP.n42 161.3
R12 VP.n41 VP.n3 161.3
R13 VP.n40 VP.n39 161.3
R14 VP.n38 VP.n37 161.3
R15 VP.n36 VP.n5 161.3
R16 VP.n35 VP.n34 161.3
R17 VP.n33 VP.n6 161.3
R18 VP.n32 VP.n31 161.3
R19 VP.n30 VP.n7 161.3
R20 VP.n29 VP.n28 161.3
R21 VP.n14 VP.t3 144.672
R22 VP.n8 VP.t1 111.344
R23 VP.n4 VP.t0 111.344
R24 VP.n0 VP.t2 111.344
R25 VP.n9 VP.t4 111.344
R26 VP.n13 VP.t5 111.344
R27 VP.n27 VP.n8 72.0476
R28 VP.n50 VP.n0 72.0476
R29 VP.n26 VP.n9 72.0476
R30 VP.n14 VP.n13 62.2244
R31 VP.n27 VP.n26 53.9692
R32 VP.n31 VP.n6 46.3896
R33 VP.n46 VP.n2 46.3896
R34 VP.n22 VP.n11 46.3896
R35 VP.n35 VP.n6 34.7644
R36 VP.n42 VP.n2 34.7644
R37 VP.n18 VP.n11 34.7644
R38 VP.n30 VP.n29 24.5923
R39 VP.n31 VP.n30 24.5923
R40 VP.n36 VP.n35 24.5923
R41 VP.n37 VP.n36 24.5923
R42 VP.n41 VP.n40 24.5923
R43 VP.n42 VP.n41 24.5923
R44 VP.n47 VP.n46 24.5923
R45 VP.n48 VP.n47 24.5923
R46 VP.n23 VP.n22 24.5923
R47 VP.n24 VP.n23 24.5923
R48 VP.n17 VP.n16 24.5923
R49 VP.n18 VP.n17 24.5923
R50 VP.n29 VP.n8 18.1985
R51 VP.n48 VP.n0 18.1985
R52 VP.n24 VP.n9 18.1985
R53 VP.n37 VP.n4 12.2964
R54 VP.n40 VP.n4 12.2964
R55 VP.n16 VP.n13 12.2964
R56 VP.n15 VP.n14 3.97924
R57 VP.n26 VP.n25 0.354861
R58 VP.n28 VP.n27 0.354861
R59 VP.n50 VP.n49 0.354861
R60 VP VP.n50 0.267071
R61 VP.n15 VP.n12 0.189894
R62 VP.n19 VP.n12 0.189894
R63 VP.n20 VP.n19 0.189894
R64 VP.n21 VP.n20 0.189894
R65 VP.n21 VP.n10 0.189894
R66 VP.n25 VP.n10 0.189894
R67 VP.n28 VP.n7 0.189894
R68 VP.n32 VP.n7 0.189894
R69 VP.n33 VP.n32 0.189894
R70 VP.n34 VP.n33 0.189894
R71 VP.n34 VP.n5 0.189894
R72 VP.n38 VP.n5 0.189894
R73 VP.n39 VP.n38 0.189894
R74 VP.n39 VP.n3 0.189894
R75 VP.n43 VP.n3 0.189894
R76 VP.n44 VP.n43 0.189894
R77 VP.n45 VP.n44 0.189894
R78 VP.n45 VP.n1 0.189894
R79 VP.n49 VP.n1 0.189894
R80 VDD1 VDD1.t0 78.9211
R81 VDD1.n1 VDD1.t5 78.8074
R82 VDD1.n1 VDD1.n0 75.1085
R83 VDD1.n3 VDD1.n2 74.3838
R84 VDD1.n3 VDD1.n1 49.1043
R85 VDD1.n2 VDD1.t4 2.13899
R86 VDD1.n2 VDD1.t1 2.13899
R87 VDD1.n0 VDD1.t3 2.13899
R88 VDD1.n0 VDD1.t2 2.13899
R89 VDD1 VDD1.n3 0.722483
R90 VTAIL.n7 VTAIL.t0 59.8437
R91 VTAIL.n11 VTAIL.t5 59.8434
R92 VTAIL.n2 VTAIL.t9 59.8434
R93 VTAIL.n10 VTAIL.t7 59.8434
R94 VTAIL.n9 VTAIL.n8 57.7052
R95 VTAIL.n6 VTAIL.n5 57.7052
R96 VTAIL.n1 VTAIL.n0 57.7049
R97 VTAIL.n4 VTAIL.n3 57.7049
R98 VTAIL.n6 VTAIL.n4 31.7117
R99 VTAIL.n11 VTAIL.n10 28.591
R100 VTAIL.n7 VTAIL.n6 3.12119
R101 VTAIL.n10 VTAIL.n9 3.12119
R102 VTAIL.n4 VTAIL.n2 3.12119
R103 VTAIL VTAIL.n11 2.28283
R104 VTAIL.n0 VTAIL.t4 2.13899
R105 VTAIL.n0 VTAIL.t2 2.13899
R106 VTAIL.n3 VTAIL.t10 2.13899
R107 VTAIL.n3 VTAIL.t11 2.13899
R108 VTAIL.n8 VTAIL.t8 2.13899
R109 VTAIL.n8 VTAIL.t6 2.13899
R110 VTAIL.n5 VTAIL.t3 2.13899
R111 VTAIL.n5 VTAIL.t1 2.13899
R112 VTAIL.n9 VTAIL.n7 2.03067
R113 VTAIL.n2 VTAIL.n1 2.03067
R114 VTAIL VTAIL.n1 0.838862
R115 B.n466 B.n139 585
R116 B.n465 B.n464 585
R117 B.n463 B.n140 585
R118 B.n462 B.n461 585
R119 B.n460 B.n141 585
R120 B.n459 B.n458 585
R121 B.n457 B.n142 585
R122 B.n456 B.n455 585
R123 B.n454 B.n143 585
R124 B.n453 B.n452 585
R125 B.n451 B.n144 585
R126 B.n450 B.n449 585
R127 B.n448 B.n145 585
R128 B.n447 B.n446 585
R129 B.n445 B.n146 585
R130 B.n444 B.n443 585
R131 B.n442 B.n147 585
R132 B.n441 B.n440 585
R133 B.n439 B.n148 585
R134 B.n438 B.n437 585
R135 B.n436 B.n149 585
R136 B.n435 B.n434 585
R137 B.n433 B.n150 585
R138 B.n432 B.n431 585
R139 B.n430 B.n151 585
R140 B.n429 B.n428 585
R141 B.n427 B.n152 585
R142 B.n426 B.n425 585
R143 B.n424 B.n153 585
R144 B.n423 B.n422 585
R145 B.n421 B.n154 585
R146 B.n420 B.n419 585
R147 B.n418 B.n155 585
R148 B.n417 B.n416 585
R149 B.n415 B.n156 585
R150 B.n414 B.n413 585
R151 B.n412 B.n157 585
R152 B.n411 B.n410 585
R153 B.n409 B.n158 585
R154 B.n408 B.n407 585
R155 B.n406 B.n159 585
R156 B.n405 B.n404 585
R157 B.n403 B.n160 585
R158 B.n402 B.n401 585
R159 B.n400 B.n161 585
R160 B.n399 B.n398 585
R161 B.n397 B.n162 585
R162 B.n396 B.n395 585
R163 B.n394 B.n163 585
R164 B.n393 B.n392 585
R165 B.n391 B.n164 585
R166 B.n389 B.n388 585
R167 B.n387 B.n167 585
R168 B.n386 B.n385 585
R169 B.n384 B.n168 585
R170 B.n383 B.n382 585
R171 B.n381 B.n169 585
R172 B.n380 B.n379 585
R173 B.n378 B.n170 585
R174 B.n377 B.n376 585
R175 B.n375 B.n171 585
R176 B.n374 B.n373 585
R177 B.n369 B.n172 585
R178 B.n368 B.n367 585
R179 B.n366 B.n173 585
R180 B.n365 B.n364 585
R181 B.n363 B.n174 585
R182 B.n362 B.n361 585
R183 B.n360 B.n175 585
R184 B.n359 B.n358 585
R185 B.n357 B.n176 585
R186 B.n356 B.n355 585
R187 B.n354 B.n177 585
R188 B.n353 B.n352 585
R189 B.n351 B.n178 585
R190 B.n350 B.n349 585
R191 B.n348 B.n179 585
R192 B.n347 B.n346 585
R193 B.n345 B.n180 585
R194 B.n344 B.n343 585
R195 B.n342 B.n181 585
R196 B.n341 B.n340 585
R197 B.n339 B.n182 585
R198 B.n338 B.n337 585
R199 B.n336 B.n183 585
R200 B.n335 B.n334 585
R201 B.n333 B.n184 585
R202 B.n332 B.n331 585
R203 B.n330 B.n185 585
R204 B.n329 B.n328 585
R205 B.n327 B.n186 585
R206 B.n326 B.n325 585
R207 B.n324 B.n187 585
R208 B.n323 B.n322 585
R209 B.n321 B.n188 585
R210 B.n320 B.n319 585
R211 B.n318 B.n189 585
R212 B.n317 B.n316 585
R213 B.n315 B.n190 585
R214 B.n314 B.n313 585
R215 B.n312 B.n191 585
R216 B.n311 B.n310 585
R217 B.n309 B.n192 585
R218 B.n308 B.n307 585
R219 B.n306 B.n193 585
R220 B.n305 B.n304 585
R221 B.n303 B.n194 585
R222 B.n302 B.n301 585
R223 B.n300 B.n195 585
R224 B.n299 B.n298 585
R225 B.n297 B.n196 585
R226 B.n296 B.n295 585
R227 B.n468 B.n467 585
R228 B.n469 B.n138 585
R229 B.n471 B.n470 585
R230 B.n472 B.n137 585
R231 B.n474 B.n473 585
R232 B.n475 B.n136 585
R233 B.n477 B.n476 585
R234 B.n478 B.n135 585
R235 B.n480 B.n479 585
R236 B.n481 B.n134 585
R237 B.n483 B.n482 585
R238 B.n484 B.n133 585
R239 B.n486 B.n485 585
R240 B.n487 B.n132 585
R241 B.n489 B.n488 585
R242 B.n490 B.n131 585
R243 B.n492 B.n491 585
R244 B.n493 B.n130 585
R245 B.n495 B.n494 585
R246 B.n496 B.n129 585
R247 B.n498 B.n497 585
R248 B.n499 B.n128 585
R249 B.n501 B.n500 585
R250 B.n502 B.n127 585
R251 B.n504 B.n503 585
R252 B.n505 B.n126 585
R253 B.n507 B.n506 585
R254 B.n508 B.n125 585
R255 B.n510 B.n509 585
R256 B.n511 B.n124 585
R257 B.n513 B.n512 585
R258 B.n514 B.n123 585
R259 B.n516 B.n515 585
R260 B.n517 B.n122 585
R261 B.n519 B.n518 585
R262 B.n520 B.n121 585
R263 B.n522 B.n521 585
R264 B.n523 B.n120 585
R265 B.n525 B.n524 585
R266 B.n526 B.n119 585
R267 B.n528 B.n527 585
R268 B.n529 B.n118 585
R269 B.n531 B.n530 585
R270 B.n532 B.n117 585
R271 B.n534 B.n533 585
R272 B.n535 B.n116 585
R273 B.n537 B.n536 585
R274 B.n538 B.n115 585
R275 B.n540 B.n539 585
R276 B.n541 B.n114 585
R277 B.n543 B.n542 585
R278 B.n544 B.n113 585
R279 B.n546 B.n545 585
R280 B.n547 B.n112 585
R281 B.n549 B.n548 585
R282 B.n550 B.n111 585
R283 B.n552 B.n551 585
R284 B.n553 B.n110 585
R285 B.n555 B.n554 585
R286 B.n556 B.n109 585
R287 B.n558 B.n557 585
R288 B.n559 B.n108 585
R289 B.n561 B.n560 585
R290 B.n562 B.n107 585
R291 B.n564 B.n563 585
R292 B.n565 B.n106 585
R293 B.n567 B.n566 585
R294 B.n568 B.n105 585
R295 B.n570 B.n569 585
R296 B.n571 B.n104 585
R297 B.n573 B.n572 585
R298 B.n574 B.n103 585
R299 B.n576 B.n575 585
R300 B.n577 B.n102 585
R301 B.n579 B.n578 585
R302 B.n580 B.n101 585
R303 B.n582 B.n581 585
R304 B.n583 B.n100 585
R305 B.n585 B.n584 585
R306 B.n586 B.n99 585
R307 B.n588 B.n587 585
R308 B.n589 B.n98 585
R309 B.n591 B.n590 585
R310 B.n592 B.n97 585
R311 B.n594 B.n593 585
R312 B.n595 B.n96 585
R313 B.n597 B.n596 585
R314 B.n598 B.n95 585
R315 B.n600 B.n599 585
R316 B.n601 B.n94 585
R317 B.n603 B.n602 585
R318 B.n604 B.n93 585
R319 B.n606 B.n605 585
R320 B.n607 B.n92 585
R321 B.n609 B.n608 585
R322 B.n610 B.n91 585
R323 B.n612 B.n611 585
R324 B.n613 B.n90 585
R325 B.n615 B.n614 585
R326 B.n616 B.n89 585
R327 B.n618 B.n617 585
R328 B.n619 B.n88 585
R329 B.n788 B.n27 585
R330 B.n787 B.n786 585
R331 B.n785 B.n28 585
R332 B.n784 B.n783 585
R333 B.n782 B.n29 585
R334 B.n781 B.n780 585
R335 B.n779 B.n30 585
R336 B.n778 B.n777 585
R337 B.n776 B.n31 585
R338 B.n775 B.n774 585
R339 B.n773 B.n32 585
R340 B.n772 B.n771 585
R341 B.n770 B.n33 585
R342 B.n769 B.n768 585
R343 B.n767 B.n34 585
R344 B.n766 B.n765 585
R345 B.n764 B.n35 585
R346 B.n763 B.n762 585
R347 B.n761 B.n36 585
R348 B.n760 B.n759 585
R349 B.n758 B.n37 585
R350 B.n757 B.n756 585
R351 B.n755 B.n38 585
R352 B.n754 B.n753 585
R353 B.n752 B.n39 585
R354 B.n751 B.n750 585
R355 B.n749 B.n40 585
R356 B.n748 B.n747 585
R357 B.n746 B.n41 585
R358 B.n745 B.n744 585
R359 B.n743 B.n42 585
R360 B.n742 B.n741 585
R361 B.n740 B.n43 585
R362 B.n739 B.n738 585
R363 B.n737 B.n44 585
R364 B.n736 B.n735 585
R365 B.n734 B.n45 585
R366 B.n733 B.n732 585
R367 B.n731 B.n46 585
R368 B.n730 B.n729 585
R369 B.n728 B.n47 585
R370 B.n727 B.n726 585
R371 B.n725 B.n48 585
R372 B.n724 B.n723 585
R373 B.n722 B.n49 585
R374 B.n721 B.n720 585
R375 B.n719 B.n50 585
R376 B.n718 B.n717 585
R377 B.n716 B.n51 585
R378 B.n715 B.n714 585
R379 B.n713 B.n52 585
R380 B.n712 B.n711 585
R381 B.n710 B.n53 585
R382 B.n709 B.n708 585
R383 B.n707 B.n57 585
R384 B.n706 B.n705 585
R385 B.n704 B.n58 585
R386 B.n703 B.n702 585
R387 B.n701 B.n59 585
R388 B.n700 B.n699 585
R389 B.n698 B.n60 585
R390 B.n696 B.n695 585
R391 B.n694 B.n63 585
R392 B.n693 B.n692 585
R393 B.n691 B.n64 585
R394 B.n690 B.n689 585
R395 B.n688 B.n65 585
R396 B.n687 B.n686 585
R397 B.n685 B.n66 585
R398 B.n684 B.n683 585
R399 B.n682 B.n67 585
R400 B.n681 B.n680 585
R401 B.n679 B.n68 585
R402 B.n678 B.n677 585
R403 B.n676 B.n69 585
R404 B.n675 B.n674 585
R405 B.n673 B.n70 585
R406 B.n672 B.n671 585
R407 B.n670 B.n71 585
R408 B.n669 B.n668 585
R409 B.n667 B.n72 585
R410 B.n666 B.n665 585
R411 B.n664 B.n73 585
R412 B.n663 B.n662 585
R413 B.n661 B.n74 585
R414 B.n660 B.n659 585
R415 B.n658 B.n75 585
R416 B.n657 B.n656 585
R417 B.n655 B.n76 585
R418 B.n654 B.n653 585
R419 B.n652 B.n77 585
R420 B.n651 B.n650 585
R421 B.n649 B.n78 585
R422 B.n648 B.n647 585
R423 B.n646 B.n79 585
R424 B.n645 B.n644 585
R425 B.n643 B.n80 585
R426 B.n642 B.n641 585
R427 B.n640 B.n81 585
R428 B.n639 B.n638 585
R429 B.n637 B.n82 585
R430 B.n636 B.n635 585
R431 B.n634 B.n83 585
R432 B.n633 B.n632 585
R433 B.n631 B.n84 585
R434 B.n630 B.n629 585
R435 B.n628 B.n85 585
R436 B.n627 B.n626 585
R437 B.n625 B.n86 585
R438 B.n624 B.n623 585
R439 B.n622 B.n87 585
R440 B.n621 B.n620 585
R441 B.n790 B.n789 585
R442 B.n791 B.n26 585
R443 B.n793 B.n792 585
R444 B.n794 B.n25 585
R445 B.n796 B.n795 585
R446 B.n797 B.n24 585
R447 B.n799 B.n798 585
R448 B.n800 B.n23 585
R449 B.n802 B.n801 585
R450 B.n803 B.n22 585
R451 B.n805 B.n804 585
R452 B.n806 B.n21 585
R453 B.n808 B.n807 585
R454 B.n809 B.n20 585
R455 B.n811 B.n810 585
R456 B.n812 B.n19 585
R457 B.n814 B.n813 585
R458 B.n815 B.n18 585
R459 B.n817 B.n816 585
R460 B.n818 B.n17 585
R461 B.n820 B.n819 585
R462 B.n821 B.n16 585
R463 B.n823 B.n822 585
R464 B.n824 B.n15 585
R465 B.n826 B.n825 585
R466 B.n827 B.n14 585
R467 B.n829 B.n828 585
R468 B.n830 B.n13 585
R469 B.n832 B.n831 585
R470 B.n833 B.n12 585
R471 B.n835 B.n834 585
R472 B.n836 B.n11 585
R473 B.n838 B.n837 585
R474 B.n839 B.n10 585
R475 B.n841 B.n840 585
R476 B.n842 B.n9 585
R477 B.n844 B.n843 585
R478 B.n845 B.n8 585
R479 B.n847 B.n846 585
R480 B.n848 B.n7 585
R481 B.n850 B.n849 585
R482 B.n851 B.n6 585
R483 B.n853 B.n852 585
R484 B.n854 B.n5 585
R485 B.n856 B.n855 585
R486 B.n857 B.n4 585
R487 B.n859 B.n858 585
R488 B.n860 B.n3 585
R489 B.n862 B.n861 585
R490 B.n863 B.n0 585
R491 B.n2 B.n1 585
R492 B.n222 B.n221 585
R493 B.n224 B.n223 585
R494 B.n225 B.n220 585
R495 B.n227 B.n226 585
R496 B.n228 B.n219 585
R497 B.n230 B.n229 585
R498 B.n231 B.n218 585
R499 B.n233 B.n232 585
R500 B.n234 B.n217 585
R501 B.n236 B.n235 585
R502 B.n237 B.n216 585
R503 B.n239 B.n238 585
R504 B.n240 B.n215 585
R505 B.n242 B.n241 585
R506 B.n243 B.n214 585
R507 B.n245 B.n244 585
R508 B.n246 B.n213 585
R509 B.n248 B.n247 585
R510 B.n249 B.n212 585
R511 B.n251 B.n250 585
R512 B.n252 B.n211 585
R513 B.n254 B.n253 585
R514 B.n255 B.n210 585
R515 B.n257 B.n256 585
R516 B.n258 B.n209 585
R517 B.n260 B.n259 585
R518 B.n261 B.n208 585
R519 B.n263 B.n262 585
R520 B.n264 B.n207 585
R521 B.n266 B.n265 585
R522 B.n267 B.n206 585
R523 B.n269 B.n268 585
R524 B.n270 B.n205 585
R525 B.n272 B.n271 585
R526 B.n273 B.n204 585
R527 B.n275 B.n274 585
R528 B.n276 B.n203 585
R529 B.n278 B.n277 585
R530 B.n279 B.n202 585
R531 B.n281 B.n280 585
R532 B.n282 B.n201 585
R533 B.n284 B.n283 585
R534 B.n285 B.n200 585
R535 B.n287 B.n286 585
R536 B.n288 B.n199 585
R537 B.n290 B.n289 585
R538 B.n291 B.n198 585
R539 B.n293 B.n292 585
R540 B.n294 B.n197 585
R541 B.n295 B.n294 502.111
R542 B.n467 B.n466 502.111
R543 B.n621 B.n88 502.111
R544 B.n790 B.n27 502.111
R545 B.n370 B.t9 320.238
R546 B.n165 B.t0 320.238
R547 B.n61 B.t6 320.238
R548 B.n54 B.t3 320.238
R549 B.n865 B.n864 256.663
R550 B.n864 B.n863 235.042
R551 B.n864 B.n2 235.042
R552 B.n165 B.t1 181.393
R553 B.n61 B.t8 181.393
R554 B.n370 B.t10 181.375
R555 B.n54 B.t5 181.375
R556 B.n295 B.n196 163.367
R557 B.n299 B.n196 163.367
R558 B.n300 B.n299 163.367
R559 B.n301 B.n300 163.367
R560 B.n301 B.n194 163.367
R561 B.n305 B.n194 163.367
R562 B.n306 B.n305 163.367
R563 B.n307 B.n306 163.367
R564 B.n307 B.n192 163.367
R565 B.n311 B.n192 163.367
R566 B.n312 B.n311 163.367
R567 B.n313 B.n312 163.367
R568 B.n313 B.n190 163.367
R569 B.n317 B.n190 163.367
R570 B.n318 B.n317 163.367
R571 B.n319 B.n318 163.367
R572 B.n319 B.n188 163.367
R573 B.n323 B.n188 163.367
R574 B.n324 B.n323 163.367
R575 B.n325 B.n324 163.367
R576 B.n325 B.n186 163.367
R577 B.n329 B.n186 163.367
R578 B.n330 B.n329 163.367
R579 B.n331 B.n330 163.367
R580 B.n331 B.n184 163.367
R581 B.n335 B.n184 163.367
R582 B.n336 B.n335 163.367
R583 B.n337 B.n336 163.367
R584 B.n337 B.n182 163.367
R585 B.n341 B.n182 163.367
R586 B.n342 B.n341 163.367
R587 B.n343 B.n342 163.367
R588 B.n343 B.n180 163.367
R589 B.n347 B.n180 163.367
R590 B.n348 B.n347 163.367
R591 B.n349 B.n348 163.367
R592 B.n349 B.n178 163.367
R593 B.n353 B.n178 163.367
R594 B.n354 B.n353 163.367
R595 B.n355 B.n354 163.367
R596 B.n355 B.n176 163.367
R597 B.n359 B.n176 163.367
R598 B.n360 B.n359 163.367
R599 B.n361 B.n360 163.367
R600 B.n361 B.n174 163.367
R601 B.n365 B.n174 163.367
R602 B.n366 B.n365 163.367
R603 B.n367 B.n366 163.367
R604 B.n367 B.n172 163.367
R605 B.n374 B.n172 163.367
R606 B.n375 B.n374 163.367
R607 B.n376 B.n375 163.367
R608 B.n376 B.n170 163.367
R609 B.n380 B.n170 163.367
R610 B.n381 B.n380 163.367
R611 B.n382 B.n381 163.367
R612 B.n382 B.n168 163.367
R613 B.n386 B.n168 163.367
R614 B.n387 B.n386 163.367
R615 B.n388 B.n387 163.367
R616 B.n388 B.n164 163.367
R617 B.n393 B.n164 163.367
R618 B.n394 B.n393 163.367
R619 B.n395 B.n394 163.367
R620 B.n395 B.n162 163.367
R621 B.n399 B.n162 163.367
R622 B.n400 B.n399 163.367
R623 B.n401 B.n400 163.367
R624 B.n401 B.n160 163.367
R625 B.n405 B.n160 163.367
R626 B.n406 B.n405 163.367
R627 B.n407 B.n406 163.367
R628 B.n407 B.n158 163.367
R629 B.n411 B.n158 163.367
R630 B.n412 B.n411 163.367
R631 B.n413 B.n412 163.367
R632 B.n413 B.n156 163.367
R633 B.n417 B.n156 163.367
R634 B.n418 B.n417 163.367
R635 B.n419 B.n418 163.367
R636 B.n419 B.n154 163.367
R637 B.n423 B.n154 163.367
R638 B.n424 B.n423 163.367
R639 B.n425 B.n424 163.367
R640 B.n425 B.n152 163.367
R641 B.n429 B.n152 163.367
R642 B.n430 B.n429 163.367
R643 B.n431 B.n430 163.367
R644 B.n431 B.n150 163.367
R645 B.n435 B.n150 163.367
R646 B.n436 B.n435 163.367
R647 B.n437 B.n436 163.367
R648 B.n437 B.n148 163.367
R649 B.n441 B.n148 163.367
R650 B.n442 B.n441 163.367
R651 B.n443 B.n442 163.367
R652 B.n443 B.n146 163.367
R653 B.n447 B.n146 163.367
R654 B.n448 B.n447 163.367
R655 B.n449 B.n448 163.367
R656 B.n449 B.n144 163.367
R657 B.n453 B.n144 163.367
R658 B.n454 B.n453 163.367
R659 B.n455 B.n454 163.367
R660 B.n455 B.n142 163.367
R661 B.n459 B.n142 163.367
R662 B.n460 B.n459 163.367
R663 B.n461 B.n460 163.367
R664 B.n461 B.n140 163.367
R665 B.n465 B.n140 163.367
R666 B.n466 B.n465 163.367
R667 B.n617 B.n88 163.367
R668 B.n617 B.n616 163.367
R669 B.n616 B.n615 163.367
R670 B.n615 B.n90 163.367
R671 B.n611 B.n90 163.367
R672 B.n611 B.n610 163.367
R673 B.n610 B.n609 163.367
R674 B.n609 B.n92 163.367
R675 B.n605 B.n92 163.367
R676 B.n605 B.n604 163.367
R677 B.n604 B.n603 163.367
R678 B.n603 B.n94 163.367
R679 B.n599 B.n94 163.367
R680 B.n599 B.n598 163.367
R681 B.n598 B.n597 163.367
R682 B.n597 B.n96 163.367
R683 B.n593 B.n96 163.367
R684 B.n593 B.n592 163.367
R685 B.n592 B.n591 163.367
R686 B.n591 B.n98 163.367
R687 B.n587 B.n98 163.367
R688 B.n587 B.n586 163.367
R689 B.n586 B.n585 163.367
R690 B.n585 B.n100 163.367
R691 B.n581 B.n100 163.367
R692 B.n581 B.n580 163.367
R693 B.n580 B.n579 163.367
R694 B.n579 B.n102 163.367
R695 B.n575 B.n102 163.367
R696 B.n575 B.n574 163.367
R697 B.n574 B.n573 163.367
R698 B.n573 B.n104 163.367
R699 B.n569 B.n104 163.367
R700 B.n569 B.n568 163.367
R701 B.n568 B.n567 163.367
R702 B.n567 B.n106 163.367
R703 B.n563 B.n106 163.367
R704 B.n563 B.n562 163.367
R705 B.n562 B.n561 163.367
R706 B.n561 B.n108 163.367
R707 B.n557 B.n108 163.367
R708 B.n557 B.n556 163.367
R709 B.n556 B.n555 163.367
R710 B.n555 B.n110 163.367
R711 B.n551 B.n110 163.367
R712 B.n551 B.n550 163.367
R713 B.n550 B.n549 163.367
R714 B.n549 B.n112 163.367
R715 B.n545 B.n112 163.367
R716 B.n545 B.n544 163.367
R717 B.n544 B.n543 163.367
R718 B.n543 B.n114 163.367
R719 B.n539 B.n114 163.367
R720 B.n539 B.n538 163.367
R721 B.n538 B.n537 163.367
R722 B.n537 B.n116 163.367
R723 B.n533 B.n116 163.367
R724 B.n533 B.n532 163.367
R725 B.n532 B.n531 163.367
R726 B.n531 B.n118 163.367
R727 B.n527 B.n118 163.367
R728 B.n527 B.n526 163.367
R729 B.n526 B.n525 163.367
R730 B.n525 B.n120 163.367
R731 B.n521 B.n120 163.367
R732 B.n521 B.n520 163.367
R733 B.n520 B.n519 163.367
R734 B.n519 B.n122 163.367
R735 B.n515 B.n122 163.367
R736 B.n515 B.n514 163.367
R737 B.n514 B.n513 163.367
R738 B.n513 B.n124 163.367
R739 B.n509 B.n124 163.367
R740 B.n509 B.n508 163.367
R741 B.n508 B.n507 163.367
R742 B.n507 B.n126 163.367
R743 B.n503 B.n126 163.367
R744 B.n503 B.n502 163.367
R745 B.n502 B.n501 163.367
R746 B.n501 B.n128 163.367
R747 B.n497 B.n128 163.367
R748 B.n497 B.n496 163.367
R749 B.n496 B.n495 163.367
R750 B.n495 B.n130 163.367
R751 B.n491 B.n130 163.367
R752 B.n491 B.n490 163.367
R753 B.n490 B.n489 163.367
R754 B.n489 B.n132 163.367
R755 B.n485 B.n132 163.367
R756 B.n485 B.n484 163.367
R757 B.n484 B.n483 163.367
R758 B.n483 B.n134 163.367
R759 B.n479 B.n134 163.367
R760 B.n479 B.n478 163.367
R761 B.n478 B.n477 163.367
R762 B.n477 B.n136 163.367
R763 B.n473 B.n136 163.367
R764 B.n473 B.n472 163.367
R765 B.n472 B.n471 163.367
R766 B.n471 B.n138 163.367
R767 B.n467 B.n138 163.367
R768 B.n786 B.n27 163.367
R769 B.n786 B.n785 163.367
R770 B.n785 B.n784 163.367
R771 B.n784 B.n29 163.367
R772 B.n780 B.n29 163.367
R773 B.n780 B.n779 163.367
R774 B.n779 B.n778 163.367
R775 B.n778 B.n31 163.367
R776 B.n774 B.n31 163.367
R777 B.n774 B.n773 163.367
R778 B.n773 B.n772 163.367
R779 B.n772 B.n33 163.367
R780 B.n768 B.n33 163.367
R781 B.n768 B.n767 163.367
R782 B.n767 B.n766 163.367
R783 B.n766 B.n35 163.367
R784 B.n762 B.n35 163.367
R785 B.n762 B.n761 163.367
R786 B.n761 B.n760 163.367
R787 B.n760 B.n37 163.367
R788 B.n756 B.n37 163.367
R789 B.n756 B.n755 163.367
R790 B.n755 B.n754 163.367
R791 B.n754 B.n39 163.367
R792 B.n750 B.n39 163.367
R793 B.n750 B.n749 163.367
R794 B.n749 B.n748 163.367
R795 B.n748 B.n41 163.367
R796 B.n744 B.n41 163.367
R797 B.n744 B.n743 163.367
R798 B.n743 B.n742 163.367
R799 B.n742 B.n43 163.367
R800 B.n738 B.n43 163.367
R801 B.n738 B.n737 163.367
R802 B.n737 B.n736 163.367
R803 B.n736 B.n45 163.367
R804 B.n732 B.n45 163.367
R805 B.n732 B.n731 163.367
R806 B.n731 B.n730 163.367
R807 B.n730 B.n47 163.367
R808 B.n726 B.n47 163.367
R809 B.n726 B.n725 163.367
R810 B.n725 B.n724 163.367
R811 B.n724 B.n49 163.367
R812 B.n720 B.n49 163.367
R813 B.n720 B.n719 163.367
R814 B.n719 B.n718 163.367
R815 B.n718 B.n51 163.367
R816 B.n714 B.n51 163.367
R817 B.n714 B.n713 163.367
R818 B.n713 B.n712 163.367
R819 B.n712 B.n53 163.367
R820 B.n708 B.n53 163.367
R821 B.n708 B.n707 163.367
R822 B.n707 B.n706 163.367
R823 B.n706 B.n58 163.367
R824 B.n702 B.n58 163.367
R825 B.n702 B.n701 163.367
R826 B.n701 B.n700 163.367
R827 B.n700 B.n60 163.367
R828 B.n695 B.n60 163.367
R829 B.n695 B.n694 163.367
R830 B.n694 B.n693 163.367
R831 B.n693 B.n64 163.367
R832 B.n689 B.n64 163.367
R833 B.n689 B.n688 163.367
R834 B.n688 B.n687 163.367
R835 B.n687 B.n66 163.367
R836 B.n683 B.n66 163.367
R837 B.n683 B.n682 163.367
R838 B.n682 B.n681 163.367
R839 B.n681 B.n68 163.367
R840 B.n677 B.n68 163.367
R841 B.n677 B.n676 163.367
R842 B.n676 B.n675 163.367
R843 B.n675 B.n70 163.367
R844 B.n671 B.n70 163.367
R845 B.n671 B.n670 163.367
R846 B.n670 B.n669 163.367
R847 B.n669 B.n72 163.367
R848 B.n665 B.n72 163.367
R849 B.n665 B.n664 163.367
R850 B.n664 B.n663 163.367
R851 B.n663 B.n74 163.367
R852 B.n659 B.n74 163.367
R853 B.n659 B.n658 163.367
R854 B.n658 B.n657 163.367
R855 B.n657 B.n76 163.367
R856 B.n653 B.n76 163.367
R857 B.n653 B.n652 163.367
R858 B.n652 B.n651 163.367
R859 B.n651 B.n78 163.367
R860 B.n647 B.n78 163.367
R861 B.n647 B.n646 163.367
R862 B.n646 B.n645 163.367
R863 B.n645 B.n80 163.367
R864 B.n641 B.n80 163.367
R865 B.n641 B.n640 163.367
R866 B.n640 B.n639 163.367
R867 B.n639 B.n82 163.367
R868 B.n635 B.n82 163.367
R869 B.n635 B.n634 163.367
R870 B.n634 B.n633 163.367
R871 B.n633 B.n84 163.367
R872 B.n629 B.n84 163.367
R873 B.n629 B.n628 163.367
R874 B.n628 B.n627 163.367
R875 B.n627 B.n86 163.367
R876 B.n623 B.n86 163.367
R877 B.n623 B.n622 163.367
R878 B.n622 B.n621 163.367
R879 B.n791 B.n790 163.367
R880 B.n792 B.n791 163.367
R881 B.n792 B.n25 163.367
R882 B.n796 B.n25 163.367
R883 B.n797 B.n796 163.367
R884 B.n798 B.n797 163.367
R885 B.n798 B.n23 163.367
R886 B.n802 B.n23 163.367
R887 B.n803 B.n802 163.367
R888 B.n804 B.n803 163.367
R889 B.n804 B.n21 163.367
R890 B.n808 B.n21 163.367
R891 B.n809 B.n808 163.367
R892 B.n810 B.n809 163.367
R893 B.n810 B.n19 163.367
R894 B.n814 B.n19 163.367
R895 B.n815 B.n814 163.367
R896 B.n816 B.n815 163.367
R897 B.n816 B.n17 163.367
R898 B.n820 B.n17 163.367
R899 B.n821 B.n820 163.367
R900 B.n822 B.n821 163.367
R901 B.n822 B.n15 163.367
R902 B.n826 B.n15 163.367
R903 B.n827 B.n826 163.367
R904 B.n828 B.n827 163.367
R905 B.n828 B.n13 163.367
R906 B.n832 B.n13 163.367
R907 B.n833 B.n832 163.367
R908 B.n834 B.n833 163.367
R909 B.n834 B.n11 163.367
R910 B.n838 B.n11 163.367
R911 B.n839 B.n838 163.367
R912 B.n840 B.n839 163.367
R913 B.n840 B.n9 163.367
R914 B.n844 B.n9 163.367
R915 B.n845 B.n844 163.367
R916 B.n846 B.n845 163.367
R917 B.n846 B.n7 163.367
R918 B.n850 B.n7 163.367
R919 B.n851 B.n850 163.367
R920 B.n852 B.n851 163.367
R921 B.n852 B.n5 163.367
R922 B.n856 B.n5 163.367
R923 B.n857 B.n856 163.367
R924 B.n858 B.n857 163.367
R925 B.n858 B.n3 163.367
R926 B.n862 B.n3 163.367
R927 B.n863 B.n862 163.367
R928 B.n222 B.n2 163.367
R929 B.n223 B.n222 163.367
R930 B.n223 B.n220 163.367
R931 B.n227 B.n220 163.367
R932 B.n228 B.n227 163.367
R933 B.n229 B.n228 163.367
R934 B.n229 B.n218 163.367
R935 B.n233 B.n218 163.367
R936 B.n234 B.n233 163.367
R937 B.n235 B.n234 163.367
R938 B.n235 B.n216 163.367
R939 B.n239 B.n216 163.367
R940 B.n240 B.n239 163.367
R941 B.n241 B.n240 163.367
R942 B.n241 B.n214 163.367
R943 B.n245 B.n214 163.367
R944 B.n246 B.n245 163.367
R945 B.n247 B.n246 163.367
R946 B.n247 B.n212 163.367
R947 B.n251 B.n212 163.367
R948 B.n252 B.n251 163.367
R949 B.n253 B.n252 163.367
R950 B.n253 B.n210 163.367
R951 B.n257 B.n210 163.367
R952 B.n258 B.n257 163.367
R953 B.n259 B.n258 163.367
R954 B.n259 B.n208 163.367
R955 B.n263 B.n208 163.367
R956 B.n264 B.n263 163.367
R957 B.n265 B.n264 163.367
R958 B.n265 B.n206 163.367
R959 B.n269 B.n206 163.367
R960 B.n270 B.n269 163.367
R961 B.n271 B.n270 163.367
R962 B.n271 B.n204 163.367
R963 B.n275 B.n204 163.367
R964 B.n276 B.n275 163.367
R965 B.n277 B.n276 163.367
R966 B.n277 B.n202 163.367
R967 B.n281 B.n202 163.367
R968 B.n282 B.n281 163.367
R969 B.n283 B.n282 163.367
R970 B.n283 B.n200 163.367
R971 B.n287 B.n200 163.367
R972 B.n288 B.n287 163.367
R973 B.n289 B.n288 163.367
R974 B.n289 B.n198 163.367
R975 B.n293 B.n198 163.367
R976 B.n294 B.n293 163.367
R977 B.n166 B.t2 111.188
R978 B.n62 B.t7 111.188
R979 B.n371 B.t11 111.168
R980 B.n55 B.t4 111.168
R981 B.n371 B.n370 70.2066
R982 B.n166 B.n165 70.2066
R983 B.n62 B.n61 70.2066
R984 B.n55 B.n54 70.2066
R985 B.n372 B.n371 59.5399
R986 B.n390 B.n166 59.5399
R987 B.n697 B.n62 59.5399
R988 B.n56 B.n55 59.5399
R989 B.n789 B.n788 32.6249
R990 B.n620 B.n619 32.6249
R991 B.n468 B.n139 32.6249
R992 B.n296 B.n197 32.6249
R993 B B.n865 18.0485
R994 B.n789 B.n26 10.6151
R995 B.n793 B.n26 10.6151
R996 B.n794 B.n793 10.6151
R997 B.n795 B.n794 10.6151
R998 B.n795 B.n24 10.6151
R999 B.n799 B.n24 10.6151
R1000 B.n800 B.n799 10.6151
R1001 B.n801 B.n800 10.6151
R1002 B.n801 B.n22 10.6151
R1003 B.n805 B.n22 10.6151
R1004 B.n806 B.n805 10.6151
R1005 B.n807 B.n806 10.6151
R1006 B.n807 B.n20 10.6151
R1007 B.n811 B.n20 10.6151
R1008 B.n812 B.n811 10.6151
R1009 B.n813 B.n812 10.6151
R1010 B.n813 B.n18 10.6151
R1011 B.n817 B.n18 10.6151
R1012 B.n818 B.n817 10.6151
R1013 B.n819 B.n818 10.6151
R1014 B.n819 B.n16 10.6151
R1015 B.n823 B.n16 10.6151
R1016 B.n824 B.n823 10.6151
R1017 B.n825 B.n824 10.6151
R1018 B.n825 B.n14 10.6151
R1019 B.n829 B.n14 10.6151
R1020 B.n830 B.n829 10.6151
R1021 B.n831 B.n830 10.6151
R1022 B.n831 B.n12 10.6151
R1023 B.n835 B.n12 10.6151
R1024 B.n836 B.n835 10.6151
R1025 B.n837 B.n836 10.6151
R1026 B.n837 B.n10 10.6151
R1027 B.n841 B.n10 10.6151
R1028 B.n842 B.n841 10.6151
R1029 B.n843 B.n842 10.6151
R1030 B.n843 B.n8 10.6151
R1031 B.n847 B.n8 10.6151
R1032 B.n848 B.n847 10.6151
R1033 B.n849 B.n848 10.6151
R1034 B.n849 B.n6 10.6151
R1035 B.n853 B.n6 10.6151
R1036 B.n854 B.n853 10.6151
R1037 B.n855 B.n854 10.6151
R1038 B.n855 B.n4 10.6151
R1039 B.n859 B.n4 10.6151
R1040 B.n860 B.n859 10.6151
R1041 B.n861 B.n860 10.6151
R1042 B.n861 B.n0 10.6151
R1043 B.n788 B.n787 10.6151
R1044 B.n787 B.n28 10.6151
R1045 B.n783 B.n28 10.6151
R1046 B.n783 B.n782 10.6151
R1047 B.n782 B.n781 10.6151
R1048 B.n781 B.n30 10.6151
R1049 B.n777 B.n30 10.6151
R1050 B.n777 B.n776 10.6151
R1051 B.n776 B.n775 10.6151
R1052 B.n775 B.n32 10.6151
R1053 B.n771 B.n32 10.6151
R1054 B.n771 B.n770 10.6151
R1055 B.n770 B.n769 10.6151
R1056 B.n769 B.n34 10.6151
R1057 B.n765 B.n34 10.6151
R1058 B.n765 B.n764 10.6151
R1059 B.n764 B.n763 10.6151
R1060 B.n763 B.n36 10.6151
R1061 B.n759 B.n36 10.6151
R1062 B.n759 B.n758 10.6151
R1063 B.n758 B.n757 10.6151
R1064 B.n757 B.n38 10.6151
R1065 B.n753 B.n38 10.6151
R1066 B.n753 B.n752 10.6151
R1067 B.n752 B.n751 10.6151
R1068 B.n751 B.n40 10.6151
R1069 B.n747 B.n40 10.6151
R1070 B.n747 B.n746 10.6151
R1071 B.n746 B.n745 10.6151
R1072 B.n745 B.n42 10.6151
R1073 B.n741 B.n42 10.6151
R1074 B.n741 B.n740 10.6151
R1075 B.n740 B.n739 10.6151
R1076 B.n739 B.n44 10.6151
R1077 B.n735 B.n44 10.6151
R1078 B.n735 B.n734 10.6151
R1079 B.n734 B.n733 10.6151
R1080 B.n733 B.n46 10.6151
R1081 B.n729 B.n46 10.6151
R1082 B.n729 B.n728 10.6151
R1083 B.n728 B.n727 10.6151
R1084 B.n727 B.n48 10.6151
R1085 B.n723 B.n48 10.6151
R1086 B.n723 B.n722 10.6151
R1087 B.n722 B.n721 10.6151
R1088 B.n721 B.n50 10.6151
R1089 B.n717 B.n50 10.6151
R1090 B.n717 B.n716 10.6151
R1091 B.n716 B.n715 10.6151
R1092 B.n715 B.n52 10.6151
R1093 B.n711 B.n710 10.6151
R1094 B.n710 B.n709 10.6151
R1095 B.n709 B.n57 10.6151
R1096 B.n705 B.n57 10.6151
R1097 B.n705 B.n704 10.6151
R1098 B.n704 B.n703 10.6151
R1099 B.n703 B.n59 10.6151
R1100 B.n699 B.n59 10.6151
R1101 B.n699 B.n698 10.6151
R1102 B.n696 B.n63 10.6151
R1103 B.n692 B.n63 10.6151
R1104 B.n692 B.n691 10.6151
R1105 B.n691 B.n690 10.6151
R1106 B.n690 B.n65 10.6151
R1107 B.n686 B.n65 10.6151
R1108 B.n686 B.n685 10.6151
R1109 B.n685 B.n684 10.6151
R1110 B.n684 B.n67 10.6151
R1111 B.n680 B.n67 10.6151
R1112 B.n680 B.n679 10.6151
R1113 B.n679 B.n678 10.6151
R1114 B.n678 B.n69 10.6151
R1115 B.n674 B.n69 10.6151
R1116 B.n674 B.n673 10.6151
R1117 B.n673 B.n672 10.6151
R1118 B.n672 B.n71 10.6151
R1119 B.n668 B.n71 10.6151
R1120 B.n668 B.n667 10.6151
R1121 B.n667 B.n666 10.6151
R1122 B.n666 B.n73 10.6151
R1123 B.n662 B.n73 10.6151
R1124 B.n662 B.n661 10.6151
R1125 B.n661 B.n660 10.6151
R1126 B.n660 B.n75 10.6151
R1127 B.n656 B.n75 10.6151
R1128 B.n656 B.n655 10.6151
R1129 B.n655 B.n654 10.6151
R1130 B.n654 B.n77 10.6151
R1131 B.n650 B.n77 10.6151
R1132 B.n650 B.n649 10.6151
R1133 B.n649 B.n648 10.6151
R1134 B.n648 B.n79 10.6151
R1135 B.n644 B.n79 10.6151
R1136 B.n644 B.n643 10.6151
R1137 B.n643 B.n642 10.6151
R1138 B.n642 B.n81 10.6151
R1139 B.n638 B.n81 10.6151
R1140 B.n638 B.n637 10.6151
R1141 B.n637 B.n636 10.6151
R1142 B.n636 B.n83 10.6151
R1143 B.n632 B.n83 10.6151
R1144 B.n632 B.n631 10.6151
R1145 B.n631 B.n630 10.6151
R1146 B.n630 B.n85 10.6151
R1147 B.n626 B.n85 10.6151
R1148 B.n626 B.n625 10.6151
R1149 B.n625 B.n624 10.6151
R1150 B.n624 B.n87 10.6151
R1151 B.n620 B.n87 10.6151
R1152 B.n619 B.n618 10.6151
R1153 B.n618 B.n89 10.6151
R1154 B.n614 B.n89 10.6151
R1155 B.n614 B.n613 10.6151
R1156 B.n613 B.n612 10.6151
R1157 B.n612 B.n91 10.6151
R1158 B.n608 B.n91 10.6151
R1159 B.n608 B.n607 10.6151
R1160 B.n607 B.n606 10.6151
R1161 B.n606 B.n93 10.6151
R1162 B.n602 B.n93 10.6151
R1163 B.n602 B.n601 10.6151
R1164 B.n601 B.n600 10.6151
R1165 B.n600 B.n95 10.6151
R1166 B.n596 B.n95 10.6151
R1167 B.n596 B.n595 10.6151
R1168 B.n595 B.n594 10.6151
R1169 B.n594 B.n97 10.6151
R1170 B.n590 B.n97 10.6151
R1171 B.n590 B.n589 10.6151
R1172 B.n589 B.n588 10.6151
R1173 B.n588 B.n99 10.6151
R1174 B.n584 B.n99 10.6151
R1175 B.n584 B.n583 10.6151
R1176 B.n583 B.n582 10.6151
R1177 B.n582 B.n101 10.6151
R1178 B.n578 B.n101 10.6151
R1179 B.n578 B.n577 10.6151
R1180 B.n577 B.n576 10.6151
R1181 B.n576 B.n103 10.6151
R1182 B.n572 B.n103 10.6151
R1183 B.n572 B.n571 10.6151
R1184 B.n571 B.n570 10.6151
R1185 B.n570 B.n105 10.6151
R1186 B.n566 B.n105 10.6151
R1187 B.n566 B.n565 10.6151
R1188 B.n565 B.n564 10.6151
R1189 B.n564 B.n107 10.6151
R1190 B.n560 B.n107 10.6151
R1191 B.n560 B.n559 10.6151
R1192 B.n559 B.n558 10.6151
R1193 B.n558 B.n109 10.6151
R1194 B.n554 B.n109 10.6151
R1195 B.n554 B.n553 10.6151
R1196 B.n553 B.n552 10.6151
R1197 B.n552 B.n111 10.6151
R1198 B.n548 B.n111 10.6151
R1199 B.n548 B.n547 10.6151
R1200 B.n547 B.n546 10.6151
R1201 B.n546 B.n113 10.6151
R1202 B.n542 B.n113 10.6151
R1203 B.n542 B.n541 10.6151
R1204 B.n541 B.n540 10.6151
R1205 B.n540 B.n115 10.6151
R1206 B.n536 B.n115 10.6151
R1207 B.n536 B.n535 10.6151
R1208 B.n535 B.n534 10.6151
R1209 B.n534 B.n117 10.6151
R1210 B.n530 B.n117 10.6151
R1211 B.n530 B.n529 10.6151
R1212 B.n529 B.n528 10.6151
R1213 B.n528 B.n119 10.6151
R1214 B.n524 B.n119 10.6151
R1215 B.n524 B.n523 10.6151
R1216 B.n523 B.n522 10.6151
R1217 B.n522 B.n121 10.6151
R1218 B.n518 B.n121 10.6151
R1219 B.n518 B.n517 10.6151
R1220 B.n517 B.n516 10.6151
R1221 B.n516 B.n123 10.6151
R1222 B.n512 B.n123 10.6151
R1223 B.n512 B.n511 10.6151
R1224 B.n511 B.n510 10.6151
R1225 B.n510 B.n125 10.6151
R1226 B.n506 B.n125 10.6151
R1227 B.n506 B.n505 10.6151
R1228 B.n505 B.n504 10.6151
R1229 B.n504 B.n127 10.6151
R1230 B.n500 B.n127 10.6151
R1231 B.n500 B.n499 10.6151
R1232 B.n499 B.n498 10.6151
R1233 B.n498 B.n129 10.6151
R1234 B.n494 B.n129 10.6151
R1235 B.n494 B.n493 10.6151
R1236 B.n493 B.n492 10.6151
R1237 B.n492 B.n131 10.6151
R1238 B.n488 B.n131 10.6151
R1239 B.n488 B.n487 10.6151
R1240 B.n487 B.n486 10.6151
R1241 B.n486 B.n133 10.6151
R1242 B.n482 B.n133 10.6151
R1243 B.n482 B.n481 10.6151
R1244 B.n481 B.n480 10.6151
R1245 B.n480 B.n135 10.6151
R1246 B.n476 B.n135 10.6151
R1247 B.n476 B.n475 10.6151
R1248 B.n475 B.n474 10.6151
R1249 B.n474 B.n137 10.6151
R1250 B.n470 B.n137 10.6151
R1251 B.n470 B.n469 10.6151
R1252 B.n469 B.n468 10.6151
R1253 B.n221 B.n1 10.6151
R1254 B.n224 B.n221 10.6151
R1255 B.n225 B.n224 10.6151
R1256 B.n226 B.n225 10.6151
R1257 B.n226 B.n219 10.6151
R1258 B.n230 B.n219 10.6151
R1259 B.n231 B.n230 10.6151
R1260 B.n232 B.n231 10.6151
R1261 B.n232 B.n217 10.6151
R1262 B.n236 B.n217 10.6151
R1263 B.n237 B.n236 10.6151
R1264 B.n238 B.n237 10.6151
R1265 B.n238 B.n215 10.6151
R1266 B.n242 B.n215 10.6151
R1267 B.n243 B.n242 10.6151
R1268 B.n244 B.n243 10.6151
R1269 B.n244 B.n213 10.6151
R1270 B.n248 B.n213 10.6151
R1271 B.n249 B.n248 10.6151
R1272 B.n250 B.n249 10.6151
R1273 B.n250 B.n211 10.6151
R1274 B.n254 B.n211 10.6151
R1275 B.n255 B.n254 10.6151
R1276 B.n256 B.n255 10.6151
R1277 B.n256 B.n209 10.6151
R1278 B.n260 B.n209 10.6151
R1279 B.n261 B.n260 10.6151
R1280 B.n262 B.n261 10.6151
R1281 B.n262 B.n207 10.6151
R1282 B.n266 B.n207 10.6151
R1283 B.n267 B.n266 10.6151
R1284 B.n268 B.n267 10.6151
R1285 B.n268 B.n205 10.6151
R1286 B.n272 B.n205 10.6151
R1287 B.n273 B.n272 10.6151
R1288 B.n274 B.n273 10.6151
R1289 B.n274 B.n203 10.6151
R1290 B.n278 B.n203 10.6151
R1291 B.n279 B.n278 10.6151
R1292 B.n280 B.n279 10.6151
R1293 B.n280 B.n201 10.6151
R1294 B.n284 B.n201 10.6151
R1295 B.n285 B.n284 10.6151
R1296 B.n286 B.n285 10.6151
R1297 B.n286 B.n199 10.6151
R1298 B.n290 B.n199 10.6151
R1299 B.n291 B.n290 10.6151
R1300 B.n292 B.n291 10.6151
R1301 B.n292 B.n197 10.6151
R1302 B.n297 B.n296 10.6151
R1303 B.n298 B.n297 10.6151
R1304 B.n298 B.n195 10.6151
R1305 B.n302 B.n195 10.6151
R1306 B.n303 B.n302 10.6151
R1307 B.n304 B.n303 10.6151
R1308 B.n304 B.n193 10.6151
R1309 B.n308 B.n193 10.6151
R1310 B.n309 B.n308 10.6151
R1311 B.n310 B.n309 10.6151
R1312 B.n310 B.n191 10.6151
R1313 B.n314 B.n191 10.6151
R1314 B.n315 B.n314 10.6151
R1315 B.n316 B.n315 10.6151
R1316 B.n316 B.n189 10.6151
R1317 B.n320 B.n189 10.6151
R1318 B.n321 B.n320 10.6151
R1319 B.n322 B.n321 10.6151
R1320 B.n322 B.n187 10.6151
R1321 B.n326 B.n187 10.6151
R1322 B.n327 B.n326 10.6151
R1323 B.n328 B.n327 10.6151
R1324 B.n328 B.n185 10.6151
R1325 B.n332 B.n185 10.6151
R1326 B.n333 B.n332 10.6151
R1327 B.n334 B.n333 10.6151
R1328 B.n334 B.n183 10.6151
R1329 B.n338 B.n183 10.6151
R1330 B.n339 B.n338 10.6151
R1331 B.n340 B.n339 10.6151
R1332 B.n340 B.n181 10.6151
R1333 B.n344 B.n181 10.6151
R1334 B.n345 B.n344 10.6151
R1335 B.n346 B.n345 10.6151
R1336 B.n346 B.n179 10.6151
R1337 B.n350 B.n179 10.6151
R1338 B.n351 B.n350 10.6151
R1339 B.n352 B.n351 10.6151
R1340 B.n352 B.n177 10.6151
R1341 B.n356 B.n177 10.6151
R1342 B.n357 B.n356 10.6151
R1343 B.n358 B.n357 10.6151
R1344 B.n358 B.n175 10.6151
R1345 B.n362 B.n175 10.6151
R1346 B.n363 B.n362 10.6151
R1347 B.n364 B.n363 10.6151
R1348 B.n364 B.n173 10.6151
R1349 B.n368 B.n173 10.6151
R1350 B.n369 B.n368 10.6151
R1351 B.n373 B.n369 10.6151
R1352 B.n377 B.n171 10.6151
R1353 B.n378 B.n377 10.6151
R1354 B.n379 B.n378 10.6151
R1355 B.n379 B.n169 10.6151
R1356 B.n383 B.n169 10.6151
R1357 B.n384 B.n383 10.6151
R1358 B.n385 B.n384 10.6151
R1359 B.n385 B.n167 10.6151
R1360 B.n389 B.n167 10.6151
R1361 B.n392 B.n391 10.6151
R1362 B.n392 B.n163 10.6151
R1363 B.n396 B.n163 10.6151
R1364 B.n397 B.n396 10.6151
R1365 B.n398 B.n397 10.6151
R1366 B.n398 B.n161 10.6151
R1367 B.n402 B.n161 10.6151
R1368 B.n403 B.n402 10.6151
R1369 B.n404 B.n403 10.6151
R1370 B.n404 B.n159 10.6151
R1371 B.n408 B.n159 10.6151
R1372 B.n409 B.n408 10.6151
R1373 B.n410 B.n409 10.6151
R1374 B.n410 B.n157 10.6151
R1375 B.n414 B.n157 10.6151
R1376 B.n415 B.n414 10.6151
R1377 B.n416 B.n415 10.6151
R1378 B.n416 B.n155 10.6151
R1379 B.n420 B.n155 10.6151
R1380 B.n421 B.n420 10.6151
R1381 B.n422 B.n421 10.6151
R1382 B.n422 B.n153 10.6151
R1383 B.n426 B.n153 10.6151
R1384 B.n427 B.n426 10.6151
R1385 B.n428 B.n427 10.6151
R1386 B.n428 B.n151 10.6151
R1387 B.n432 B.n151 10.6151
R1388 B.n433 B.n432 10.6151
R1389 B.n434 B.n433 10.6151
R1390 B.n434 B.n149 10.6151
R1391 B.n438 B.n149 10.6151
R1392 B.n439 B.n438 10.6151
R1393 B.n440 B.n439 10.6151
R1394 B.n440 B.n147 10.6151
R1395 B.n444 B.n147 10.6151
R1396 B.n445 B.n444 10.6151
R1397 B.n446 B.n445 10.6151
R1398 B.n446 B.n145 10.6151
R1399 B.n450 B.n145 10.6151
R1400 B.n451 B.n450 10.6151
R1401 B.n452 B.n451 10.6151
R1402 B.n452 B.n143 10.6151
R1403 B.n456 B.n143 10.6151
R1404 B.n457 B.n456 10.6151
R1405 B.n458 B.n457 10.6151
R1406 B.n458 B.n141 10.6151
R1407 B.n462 B.n141 10.6151
R1408 B.n463 B.n462 10.6151
R1409 B.n464 B.n463 10.6151
R1410 B.n464 B.n139 10.6151
R1411 B.n56 B.n52 9.36635
R1412 B.n697 B.n696 9.36635
R1413 B.n373 B.n372 9.36635
R1414 B.n391 B.n390 9.36635
R1415 B.n865 B.n0 8.11757
R1416 B.n865 B.n1 8.11757
R1417 B.n711 B.n56 1.24928
R1418 B.n698 B.n697 1.24928
R1419 B.n372 B.n171 1.24928
R1420 B.n390 B.n389 1.24928
R1421 VN.n34 VN.n33 161.3
R1422 VN.n32 VN.n19 161.3
R1423 VN.n31 VN.n30 161.3
R1424 VN.n29 VN.n20 161.3
R1425 VN.n28 VN.n27 161.3
R1426 VN.n26 VN.n21 161.3
R1427 VN.n25 VN.n24 161.3
R1428 VN.n16 VN.n15 161.3
R1429 VN.n14 VN.n1 161.3
R1430 VN.n13 VN.n12 161.3
R1431 VN.n11 VN.n2 161.3
R1432 VN.n10 VN.n9 161.3
R1433 VN.n8 VN.n3 161.3
R1434 VN.n7 VN.n6 161.3
R1435 VN.n23 VN.t1 144.672
R1436 VN.n5 VN.t3 144.672
R1437 VN.n4 VN.t0 111.344
R1438 VN.n0 VN.t5 111.344
R1439 VN.n22 VN.t2 111.344
R1440 VN.n18 VN.t4 111.344
R1441 VN.n17 VN.n0 72.0476
R1442 VN.n35 VN.n18 72.0476
R1443 VN.n5 VN.n4 62.2244
R1444 VN.n23 VN.n22 62.2244
R1445 VN VN.n35 54.1345
R1446 VN.n13 VN.n2 46.3896
R1447 VN.n31 VN.n20 46.3896
R1448 VN.n9 VN.n2 34.7644
R1449 VN.n27 VN.n20 34.7644
R1450 VN.n8 VN.n7 24.5923
R1451 VN.n9 VN.n8 24.5923
R1452 VN.n14 VN.n13 24.5923
R1453 VN.n15 VN.n14 24.5923
R1454 VN.n27 VN.n26 24.5923
R1455 VN.n26 VN.n25 24.5923
R1456 VN.n33 VN.n32 24.5923
R1457 VN.n32 VN.n31 24.5923
R1458 VN.n15 VN.n0 18.1985
R1459 VN.n33 VN.n18 18.1985
R1460 VN.n7 VN.n4 12.2964
R1461 VN.n25 VN.n22 12.2964
R1462 VN.n24 VN.n23 3.97927
R1463 VN.n6 VN.n5 3.97927
R1464 VN.n35 VN.n34 0.354861
R1465 VN.n17 VN.n16 0.354861
R1466 VN VN.n17 0.267071
R1467 VN.n34 VN.n19 0.189894
R1468 VN.n30 VN.n19 0.189894
R1469 VN.n30 VN.n29 0.189894
R1470 VN.n29 VN.n28 0.189894
R1471 VN.n28 VN.n21 0.189894
R1472 VN.n24 VN.n21 0.189894
R1473 VN.n6 VN.n3 0.189894
R1474 VN.n10 VN.n3 0.189894
R1475 VN.n11 VN.n10 0.189894
R1476 VN.n12 VN.n11 0.189894
R1477 VN.n12 VN.n1 0.189894
R1478 VN.n16 VN.n1 0.189894
R1479 VDD2.n1 VDD2.t2 78.8074
R1480 VDD2.n2 VDD2.t1 76.5224
R1481 VDD2.n1 VDD2.n0 75.1085
R1482 VDD2 VDD2.n3 75.1057
R1483 VDD2.n2 VDD2.n1 46.961
R1484 VDD2 VDD2.n2 2.39921
R1485 VDD2.n3 VDD2.t3 2.13899
R1486 VDD2.n3 VDD2.t4 2.13899
R1487 VDD2.n0 VDD2.t5 2.13899
R1488 VDD2.n0 VDD2.t0 2.13899
C0 VTAIL VN 8.941629f
C1 w_n3866_n4008# B 11.5262f
C2 VTAIL VP 8.9559f
C3 B VDD2 2.62035f
C4 w_n3866_n4008# VDD1 2.67673f
C5 VDD1 VDD2 1.6757f
C6 w_n3866_n4008# VDD2 2.78385f
C7 VP VN 8.18296f
C8 VTAIL B 4.70582f
C9 VTAIL VDD1 8.99962f
C10 w_n3866_n4008# VTAIL 3.46724f
C11 B VN 1.35475f
C12 VTAIL VDD2 9.05511f
C13 B VP 2.19594f
C14 VDD1 VN 0.151913f
C15 w_n3866_n4008# VN 7.53963f
C16 VDD1 VP 9.126821f
C17 w_n3866_n4008# VP 8.04137f
C18 VN VDD2 8.765f
C19 VP VDD2 0.517269f
C20 VDD1 B 2.52971f
C21 VDD2 VSUBS 2.15964f
C22 VDD1 VSUBS 2.7006f
C23 VTAIL VSUBS 1.43926f
C24 VN VSUBS 6.61863f
C25 VP VSUBS 3.595553f
C26 B VSUBS 5.589792f
C27 w_n3866_n4008# VSUBS 0.189975p
C28 VDD2.t2 VSUBS 3.56494f
C29 VDD2.t5 VSUBS 0.333206f
C30 VDD2.t0 VSUBS 0.333206f
C31 VDD2.n0 VSUBS 2.73293f
C32 VDD2.n1 VSUBS 4.36395f
C33 VDD2.t1 VSUBS 3.54103f
C34 VDD2.n2 VSUBS 3.88963f
C35 VDD2.t3 VSUBS 0.333206f
C36 VDD2.t4 VSUBS 0.333206f
C37 VDD2.n3 VSUBS 2.73288f
C38 VN.t5 VSUBS 3.42013f
C39 VN.n0 VSUBS 1.2914f
C40 VN.n1 VSUBS 0.024951f
C41 VN.n2 VSUBS 0.021321f
C42 VN.n3 VSUBS 0.024951f
C43 VN.t0 VSUBS 3.42013f
C44 VN.n4 VSUBS 1.27101f
C45 VN.t3 VSUBS 3.73554f
C46 VN.n5 VSUBS 1.21476f
C47 VN.n6 VSUBS 0.290986f
C48 VN.n7 VSUBS 0.034849f
C49 VN.n8 VSUBS 0.04627f
C50 VN.n9 VSUBS 0.050146f
C51 VN.n10 VSUBS 0.024951f
C52 VN.n11 VSUBS 0.024951f
C53 VN.n12 VSUBS 0.024951f
C54 VN.n13 VSUBS 0.047343f
C55 VN.n14 VSUBS 0.04627f
C56 VN.n15 VSUBS 0.040331f
C57 VN.n16 VSUBS 0.040264f
C58 VN.n17 VSUBS 0.056536f
C59 VN.t4 VSUBS 3.42013f
C60 VN.n18 VSUBS 1.2914f
C61 VN.n19 VSUBS 0.024951f
C62 VN.n20 VSUBS 0.021321f
C63 VN.n21 VSUBS 0.024951f
C64 VN.t2 VSUBS 3.42013f
C65 VN.n22 VSUBS 1.27101f
C66 VN.t1 VSUBS 3.73554f
C67 VN.n23 VSUBS 1.21476f
C68 VN.n24 VSUBS 0.290986f
C69 VN.n25 VSUBS 0.034849f
C70 VN.n26 VSUBS 0.04627f
C71 VN.n27 VSUBS 0.050146f
C72 VN.n28 VSUBS 0.024951f
C73 VN.n29 VSUBS 0.024951f
C74 VN.n30 VSUBS 0.024951f
C75 VN.n31 VSUBS 0.047343f
C76 VN.n32 VSUBS 0.04627f
C77 VN.n33 VSUBS 0.040331f
C78 VN.n34 VSUBS 0.040264f
C79 VN.n35 VSUBS 1.58856f
C80 B.n0 VSUBS 0.006911f
C81 B.n1 VSUBS 0.006911f
C82 B.n2 VSUBS 0.010221f
C83 B.n3 VSUBS 0.007832f
C84 B.n4 VSUBS 0.007832f
C85 B.n5 VSUBS 0.007832f
C86 B.n6 VSUBS 0.007832f
C87 B.n7 VSUBS 0.007832f
C88 B.n8 VSUBS 0.007832f
C89 B.n9 VSUBS 0.007832f
C90 B.n10 VSUBS 0.007832f
C91 B.n11 VSUBS 0.007832f
C92 B.n12 VSUBS 0.007832f
C93 B.n13 VSUBS 0.007832f
C94 B.n14 VSUBS 0.007832f
C95 B.n15 VSUBS 0.007832f
C96 B.n16 VSUBS 0.007832f
C97 B.n17 VSUBS 0.007832f
C98 B.n18 VSUBS 0.007832f
C99 B.n19 VSUBS 0.007832f
C100 B.n20 VSUBS 0.007832f
C101 B.n21 VSUBS 0.007832f
C102 B.n22 VSUBS 0.007832f
C103 B.n23 VSUBS 0.007832f
C104 B.n24 VSUBS 0.007832f
C105 B.n25 VSUBS 0.007832f
C106 B.n26 VSUBS 0.007832f
C107 B.n27 VSUBS 0.019048f
C108 B.n28 VSUBS 0.007832f
C109 B.n29 VSUBS 0.007832f
C110 B.n30 VSUBS 0.007832f
C111 B.n31 VSUBS 0.007832f
C112 B.n32 VSUBS 0.007832f
C113 B.n33 VSUBS 0.007832f
C114 B.n34 VSUBS 0.007832f
C115 B.n35 VSUBS 0.007832f
C116 B.n36 VSUBS 0.007832f
C117 B.n37 VSUBS 0.007832f
C118 B.n38 VSUBS 0.007832f
C119 B.n39 VSUBS 0.007832f
C120 B.n40 VSUBS 0.007832f
C121 B.n41 VSUBS 0.007832f
C122 B.n42 VSUBS 0.007832f
C123 B.n43 VSUBS 0.007832f
C124 B.n44 VSUBS 0.007832f
C125 B.n45 VSUBS 0.007832f
C126 B.n46 VSUBS 0.007832f
C127 B.n47 VSUBS 0.007832f
C128 B.n48 VSUBS 0.007832f
C129 B.n49 VSUBS 0.007832f
C130 B.n50 VSUBS 0.007832f
C131 B.n51 VSUBS 0.007832f
C132 B.n52 VSUBS 0.007371f
C133 B.n53 VSUBS 0.007832f
C134 B.t4 VSUBS 0.566802f
C135 B.t5 VSUBS 0.594888f
C136 B.t3 VSUBS 2.55172f
C137 B.n54 VSUBS 0.342118f
C138 B.n55 VSUBS 0.083728f
C139 B.n56 VSUBS 0.018146f
C140 B.n57 VSUBS 0.007832f
C141 B.n58 VSUBS 0.007832f
C142 B.n59 VSUBS 0.007832f
C143 B.n60 VSUBS 0.007832f
C144 B.t7 VSUBS 0.566786f
C145 B.t8 VSUBS 0.594875f
C146 B.t6 VSUBS 2.55172f
C147 B.n61 VSUBS 0.342131f
C148 B.n62 VSUBS 0.083744f
C149 B.n63 VSUBS 0.007832f
C150 B.n64 VSUBS 0.007832f
C151 B.n65 VSUBS 0.007832f
C152 B.n66 VSUBS 0.007832f
C153 B.n67 VSUBS 0.007832f
C154 B.n68 VSUBS 0.007832f
C155 B.n69 VSUBS 0.007832f
C156 B.n70 VSUBS 0.007832f
C157 B.n71 VSUBS 0.007832f
C158 B.n72 VSUBS 0.007832f
C159 B.n73 VSUBS 0.007832f
C160 B.n74 VSUBS 0.007832f
C161 B.n75 VSUBS 0.007832f
C162 B.n76 VSUBS 0.007832f
C163 B.n77 VSUBS 0.007832f
C164 B.n78 VSUBS 0.007832f
C165 B.n79 VSUBS 0.007832f
C166 B.n80 VSUBS 0.007832f
C167 B.n81 VSUBS 0.007832f
C168 B.n82 VSUBS 0.007832f
C169 B.n83 VSUBS 0.007832f
C170 B.n84 VSUBS 0.007832f
C171 B.n85 VSUBS 0.007832f
C172 B.n86 VSUBS 0.007832f
C173 B.n87 VSUBS 0.007832f
C174 B.n88 VSUBS 0.017579f
C175 B.n89 VSUBS 0.007832f
C176 B.n90 VSUBS 0.007832f
C177 B.n91 VSUBS 0.007832f
C178 B.n92 VSUBS 0.007832f
C179 B.n93 VSUBS 0.007832f
C180 B.n94 VSUBS 0.007832f
C181 B.n95 VSUBS 0.007832f
C182 B.n96 VSUBS 0.007832f
C183 B.n97 VSUBS 0.007832f
C184 B.n98 VSUBS 0.007832f
C185 B.n99 VSUBS 0.007832f
C186 B.n100 VSUBS 0.007832f
C187 B.n101 VSUBS 0.007832f
C188 B.n102 VSUBS 0.007832f
C189 B.n103 VSUBS 0.007832f
C190 B.n104 VSUBS 0.007832f
C191 B.n105 VSUBS 0.007832f
C192 B.n106 VSUBS 0.007832f
C193 B.n107 VSUBS 0.007832f
C194 B.n108 VSUBS 0.007832f
C195 B.n109 VSUBS 0.007832f
C196 B.n110 VSUBS 0.007832f
C197 B.n111 VSUBS 0.007832f
C198 B.n112 VSUBS 0.007832f
C199 B.n113 VSUBS 0.007832f
C200 B.n114 VSUBS 0.007832f
C201 B.n115 VSUBS 0.007832f
C202 B.n116 VSUBS 0.007832f
C203 B.n117 VSUBS 0.007832f
C204 B.n118 VSUBS 0.007832f
C205 B.n119 VSUBS 0.007832f
C206 B.n120 VSUBS 0.007832f
C207 B.n121 VSUBS 0.007832f
C208 B.n122 VSUBS 0.007832f
C209 B.n123 VSUBS 0.007832f
C210 B.n124 VSUBS 0.007832f
C211 B.n125 VSUBS 0.007832f
C212 B.n126 VSUBS 0.007832f
C213 B.n127 VSUBS 0.007832f
C214 B.n128 VSUBS 0.007832f
C215 B.n129 VSUBS 0.007832f
C216 B.n130 VSUBS 0.007832f
C217 B.n131 VSUBS 0.007832f
C218 B.n132 VSUBS 0.007832f
C219 B.n133 VSUBS 0.007832f
C220 B.n134 VSUBS 0.007832f
C221 B.n135 VSUBS 0.007832f
C222 B.n136 VSUBS 0.007832f
C223 B.n137 VSUBS 0.007832f
C224 B.n138 VSUBS 0.007832f
C225 B.n139 VSUBS 0.018121f
C226 B.n140 VSUBS 0.007832f
C227 B.n141 VSUBS 0.007832f
C228 B.n142 VSUBS 0.007832f
C229 B.n143 VSUBS 0.007832f
C230 B.n144 VSUBS 0.007832f
C231 B.n145 VSUBS 0.007832f
C232 B.n146 VSUBS 0.007832f
C233 B.n147 VSUBS 0.007832f
C234 B.n148 VSUBS 0.007832f
C235 B.n149 VSUBS 0.007832f
C236 B.n150 VSUBS 0.007832f
C237 B.n151 VSUBS 0.007832f
C238 B.n152 VSUBS 0.007832f
C239 B.n153 VSUBS 0.007832f
C240 B.n154 VSUBS 0.007832f
C241 B.n155 VSUBS 0.007832f
C242 B.n156 VSUBS 0.007832f
C243 B.n157 VSUBS 0.007832f
C244 B.n158 VSUBS 0.007832f
C245 B.n159 VSUBS 0.007832f
C246 B.n160 VSUBS 0.007832f
C247 B.n161 VSUBS 0.007832f
C248 B.n162 VSUBS 0.007832f
C249 B.n163 VSUBS 0.007832f
C250 B.n164 VSUBS 0.007832f
C251 B.t2 VSUBS 0.566786f
C252 B.t1 VSUBS 0.594875f
C253 B.t0 VSUBS 2.55172f
C254 B.n165 VSUBS 0.342131f
C255 B.n166 VSUBS 0.083744f
C256 B.n167 VSUBS 0.007832f
C257 B.n168 VSUBS 0.007832f
C258 B.n169 VSUBS 0.007832f
C259 B.n170 VSUBS 0.007832f
C260 B.n171 VSUBS 0.004377f
C261 B.n172 VSUBS 0.007832f
C262 B.n173 VSUBS 0.007832f
C263 B.n174 VSUBS 0.007832f
C264 B.n175 VSUBS 0.007832f
C265 B.n176 VSUBS 0.007832f
C266 B.n177 VSUBS 0.007832f
C267 B.n178 VSUBS 0.007832f
C268 B.n179 VSUBS 0.007832f
C269 B.n180 VSUBS 0.007832f
C270 B.n181 VSUBS 0.007832f
C271 B.n182 VSUBS 0.007832f
C272 B.n183 VSUBS 0.007832f
C273 B.n184 VSUBS 0.007832f
C274 B.n185 VSUBS 0.007832f
C275 B.n186 VSUBS 0.007832f
C276 B.n187 VSUBS 0.007832f
C277 B.n188 VSUBS 0.007832f
C278 B.n189 VSUBS 0.007832f
C279 B.n190 VSUBS 0.007832f
C280 B.n191 VSUBS 0.007832f
C281 B.n192 VSUBS 0.007832f
C282 B.n193 VSUBS 0.007832f
C283 B.n194 VSUBS 0.007832f
C284 B.n195 VSUBS 0.007832f
C285 B.n196 VSUBS 0.007832f
C286 B.n197 VSUBS 0.017579f
C287 B.n198 VSUBS 0.007832f
C288 B.n199 VSUBS 0.007832f
C289 B.n200 VSUBS 0.007832f
C290 B.n201 VSUBS 0.007832f
C291 B.n202 VSUBS 0.007832f
C292 B.n203 VSUBS 0.007832f
C293 B.n204 VSUBS 0.007832f
C294 B.n205 VSUBS 0.007832f
C295 B.n206 VSUBS 0.007832f
C296 B.n207 VSUBS 0.007832f
C297 B.n208 VSUBS 0.007832f
C298 B.n209 VSUBS 0.007832f
C299 B.n210 VSUBS 0.007832f
C300 B.n211 VSUBS 0.007832f
C301 B.n212 VSUBS 0.007832f
C302 B.n213 VSUBS 0.007832f
C303 B.n214 VSUBS 0.007832f
C304 B.n215 VSUBS 0.007832f
C305 B.n216 VSUBS 0.007832f
C306 B.n217 VSUBS 0.007832f
C307 B.n218 VSUBS 0.007832f
C308 B.n219 VSUBS 0.007832f
C309 B.n220 VSUBS 0.007832f
C310 B.n221 VSUBS 0.007832f
C311 B.n222 VSUBS 0.007832f
C312 B.n223 VSUBS 0.007832f
C313 B.n224 VSUBS 0.007832f
C314 B.n225 VSUBS 0.007832f
C315 B.n226 VSUBS 0.007832f
C316 B.n227 VSUBS 0.007832f
C317 B.n228 VSUBS 0.007832f
C318 B.n229 VSUBS 0.007832f
C319 B.n230 VSUBS 0.007832f
C320 B.n231 VSUBS 0.007832f
C321 B.n232 VSUBS 0.007832f
C322 B.n233 VSUBS 0.007832f
C323 B.n234 VSUBS 0.007832f
C324 B.n235 VSUBS 0.007832f
C325 B.n236 VSUBS 0.007832f
C326 B.n237 VSUBS 0.007832f
C327 B.n238 VSUBS 0.007832f
C328 B.n239 VSUBS 0.007832f
C329 B.n240 VSUBS 0.007832f
C330 B.n241 VSUBS 0.007832f
C331 B.n242 VSUBS 0.007832f
C332 B.n243 VSUBS 0.007832f
C333 B.n244 VSUBS 0.007832f
C334 B.n245 VSUBS 0.007832f
C335 B.n246 VSUBS 0.007832f
C336 B.n247 VSUBS 0.007832f
C337 B.n248 VSUBS 0.007832f
C338 B.n249 VSUBS 0.007832f
C339 B.n250 VSUBS 0.007832f
C340 B.n251 VSUBS 0.007832f
C341 B.n252 VSUBS 0.007832f
C342 B.n253 VSUBS 0.007832f
C343 B.n254 VSUBS 0.007832f
C344 B.n255 VSUBS 0.007832f
C345 B.n256 VSUBS 0.007832f
C346 B.n257 VSUBS 0.007832f
C347 B.n258 VSUBS 0.007832f
C348 B.n259 VSUBS 0.007832f
C349 B.n260 VSUBS 0.007832f
C350 B.n261 VSUBS 0.007832f
C351 B.n262 VSUBS 0.007832f
C352 B.n263 VSUBS 0.007832f
C353 B.n264 VSUBS 0.007832f
C354 B.n265 VSUBS 0.007832f
C355 B.n266 VSUBS 0.007832f
C356 B.n267 VSUBS 0.007832f
C357 B.n268 VSUBS 0.007832f
C358 B.n269 VSUBS 0.007832f
C359 B.n270 VSUBS 0.007832f
C360 B.n271 VSUBS 0.007832f
C361 B.n272 VSUBS 0.007832f
C362 B.n273 VSUBS 0.007832f
C363 B.n274 VSUBS 0.007832f
C364 B.n275 VSUBS 0.007832f
C365 B.n276 VSUBS 0.007832f
C366 B.n277 VSUBS 0.007832f
C367 B.n278 VSUBS 0.007832f
C368 B.n279 VSUBS 0.007832f
C369 B.n280 VSUBS 0.007832f
C370 B.n281 VSUBS 0.007832f
C371 B.n282 VSUBS 0.007832f
C372 B.n283 VSUBS 0.007832f
C373 B.n284 VSUBS 0.007832f
C374 B.n285 VSUBS 0.007832f
C375 B.n286 VSUBS 0.007832f
C376 B.n287 VSUBS 0.007832f
C377 B.n288 VSUBS 0.007832f
C378 B.n289 VSUBS 0.007832f
C379 B.n290 VSUBS 0.007832f
C380 B.n291 VSUBS 0.007832f
C381 B.n292 VSUBS 0.007832f
C382 B.n293 VSUBS 0.007832f
C383 B.n294 VSUBS 0.017579f
C384 B.n295 VSUBS 0.019048f
C385 B.n296 VSUBS 0.019048f
C386 B.n297 VSUBS 0.007832f
C387 B.n298 VSUBS 0.007832f
C388 B.n299 VSUBS 0.007832f
C389 B.n300 VSUBS 0.007832f
C390 B.n301 VSUBS 0.007832f
C391 B.n302 VSUBS 0.007832f
C392 B.n303 VSUBS 0.007832f
C393 B.n304 VSUBS 0.007832f
C394 B.n305 VSUBS 0.007832f
C395 B.n306 VSUBS 0.007832f
C396 B.n307 VSUBS 0.007832f
C397 B.n308 VSUBS 0.007832f
C398 B.n309 VSUBS 0.007832f
C399 B.n310 VSUBS 0.007832f
C400 B.n311 VSUBS 0.007832f
C401 B.n312 VSUBS 0.007832f
C402 B.n313 VSUBS 0.007832f
C403 B.n314 VSUBS 0.007832f
C404 B.n315 VSUBS 0.007832f
C405 B.n316 VSUBS 0.007832f
C406 B.n317 VSUBS 0.007832f
C407 B.n318 VSUBS 0.007832f
C408 B.n319 VSUBS 0.007832f
C409 B.n320 VSUBS 0.007832f
C410 B.n321 VSUBS 0.007832f
C411 B.n322 VSUBS 0.007832f
C412 B.n323 VSUBS 0.007832f
C413 B.n324 VSUBS 0.007832f
C414 B.n325 VSUBS 0.007832f
C415 B.n326 VSUBS 0.007832f
C416 B.n327 VSUBS 0.007832f
C417 B.n328 VSUBS 0.007832f
C418 B.n329 VSUBS 0.007832f
C419 B.n330 VSUBS 0.007832f
C420 B.n331 VSUBS 0.007832f
C421 B.n332 VSUBS 0.007832f
C422 B.n333 VSUBS 0.007832f
C423 B.n334 VSUBS 0.007832f
C424 B.n335 VSUBS 0.007832f
C425 B.n336 VSUBS 0.007832f
C426 B.n337 VSUBS 0.007832f
C427 B.n338 VSUBS 0.007832f
C428 B.n339 VSUBS 0.007832f
C429 B.n340 VSUBS 0.007832f
C430 B.n341 VSUBS 0.007832f
C431 B.n342 VSUBS 0.007832f
C432 B.n343 VSUBS 0.007832f
C433 B.n344 VSUBS 0.007832f
C434 B.n345 VSUBS 0.007832f
C435 B.n346 VSUBS 0.007832f
C436 B.n347 VSUBS 0.007832f
C437 B.n348 VSUBS 0.007832f
C438 B.n349 VSUBS 0.007832f
C439 B.n350 VSUBS 0.007832f
C440 B.n351 VSUBS 0.007832f
C441 B.n352 VSUBS 0.007832f
C442 B.n353 VSUBS 0.007832f
C443 B.n354 VSUBS 0.007832f
C444 B.n355 VSUBS 0.007832f
C445 B.n356 VSUBS 0.007832f
C446 B.n357 VSUBS 0.007832f
C447 B.n358 VSUBS 0.007832f
C448 B.n359 VSUBS 0.007832f
C449 B.n360 VSUBS 0.007832f
C450 B.n361 VSUBS 0.007832f
C451 B.n362 VSUBS 0.007832f
C452 B.n363 VSUBS 0.007832f
C453 B.n364 VSUBS 0.007832f
C454 B.n365 VSUBS 0.007832f
C455 B.n366 VSUBS 0.007832f
C456 B.n367 VSUBS 0.007832f
C457 B.n368 VSUBS 0.007832f
C458 B.n369 VSUBS 0.007832f
C459 B.t11 VSUBS 0.566802f
C460 B.t10 VSUBS 0.594888f
C461 B.t9 VSUBS 2.55172f
C462 B.n370 VSUBS 0.342118f
C463 B.n371 VSUBS 0.083728f
C464 B.n372 VSUBS 0.018146f
C465 B.n373 VSUBS 0.007371f
C466 B.n374 VSUBS 0.007832f
C467 B.n375 VSUBS 0.007832f
C468 B.n376 VSUBS 0.007832f
C469 B.n377 VSUBS 0.007832f
C470 B.n378 VSUBS 0.007832f
C471 B.n379 VSUBS 0.007832f
C472 B.n380 VSUBS 0.007832f
C473 B.n381 VSUBS 0.007832f
C474 B.n382 VSUBS 0.007832f
C475 B.n383 VSUBS 0.007832f
C476 B.n384 VSUBS 0.007832f
C477 B.n385 VSUBS 0.007832f
C478 B.n386 VSUBS 0.007832f
C479 B.n387 VSUBS 0.007832f
C480 B.n388 VSUBS 0.007832f
C481 B.n389 VSUBS 0.004377f
C482 B.n390 VSUBS 0.018146f
C483 B.n391 VSUBS 0.007371f
C484 B.n392 VSUBS 0.007832f
C485 B.n393 VSUBS 0.007832f
C486 B.n394 VSUBS 0.007832f
C487 B.n395 VSUBS 0.007832f
C488 B.n396 VSUBS 0.007832f
C489 B.n397 VSUBS 0.007832f
C490 B.n398 VSUBS 0.007832f
C491 B.n399 VSUBS 0.007832f
C492 B.n400 VSUBS 0.007832f
C493 B.n401 VSUBS 0.007832f
C494 B.n402 VSUBS 0.007832f
C495 B.n403 VSUBS 0.007832f
C496 B.n404 VSUBS 0.007832f
C497 B.n405 VSUBS 0.007832f
C498 B.n406 VSUBS 0.007832f
C499 B.n407 VSUBS 0.007832f
C500 B.n408 VSUBS 0.007832f
C501 B.n409 VSUBS 0.007832f
C502 B.n410 VSUBS 0.007832f
C503 B.n411 VSUBS 0.007832f
C504 B.n412 VSUBS 0.007832f
C505 B.n413 VSUBS 0.007832f
C506 B.n414 VSUBS 0.007832f
C507 B.n415 VSUBS 0.007832f
C508 B.n416 VSUBS 0.007832f
C509 B.n417 VSUBS 0.007832f
C510 B.n418 VSUBS 0.007832f
C511 B.n419 VSUBS 0.007832f
C512 B.n420 VSUBS 0.007832f
C513 B.n421 VSUBS 0.007832f
C514 B.n422 VSUBS 0.007832f
C515 B.n423 VSUBS 0.007832f
C516 B.n424 VSUBS 0.007832f
C517 B.n425 VSUBS 0.007832f
C518 B.n426 VSUBS 0.007832f
C519 B.n427 VSUBS 0.007832f
C520 B.n428 VSUBS 0.007832f
C521 B.n429 VSUBS 0.007832f
C522 B.n430 VSUBS 0.007832f
C523 B.n431 VSUBS 0.007832f
C524 B.n432 VSUBS 0.007832f
C525 B.n433 VSUBS 0.007832f
C526 B.n434 VSUBS 0.007832f
C527 B.n435 VSUBS 0.007832f
C528 B.n436 VSUBS 0.007832f
C529 B.n437 VSUBS 0.007832f
C530 B.n438 VSUBS 0.007832f
C531 B.n439 VSUBS 0.007832f
C532 B.n440 VSUBS 0.007832f
C533 B.n441 VSUBS 0.007832f
C534 B.n442 VSUBS 0.007832f
C535 B.n443 VSUBS 0.007832f
C536 B.n444 VSUBS 0.007832f
C537 B.n445 VSUBS 0.007832f
C538 B.n446 VSUBS 0.007832f
C539 B.n447 VSUBS 0.007832f
C540 B.n448 VSUBS 0.007832f
C541 B.n449 VSUBS 0.007832f
C542 B.n450 VSUBS 0.007832f
C543 B.n451 VSUBS 0.007832f
C544 B.n452 VSUBS 0.007832f
C545 B.n453 VSUBS 0.007832f
C546 B.n454 VSUBS 0.007832f
C547 B.n455 VSUBS 0.007832f
C548 B.n456 VSUBS 0.007832f
C549 B.n457 VSUBS 0.007832f
C550 B.n458 VSUBS 0.007832f
C551 B.n459 VSUBS 0.007832f
C552 B.n460 VSUBS 0.007832f
C553 B.n461 VSUBS 0.007832f
C554 B.n462 VSUBS 0.007832f
C555 B.n463 VSUBS 0.007832f
C556 B.n464 VSUBS 0.007832f
C557 B.n465 VSUBS 0.007832f
C558 B.n466 VSUBS 0.019048f
C559 B.n467 VSUBS 0.017579f
C560 B.n468 VSUBS 0.018506f
C561 B.n469 VSUBS 0.007832f
C562 B.n470 VSUBS 0.007832f
C563 B.n471 VSUBS 0.007832f
C564 B.n472 VSUBS 0.007832f
C565 B.n473 VSUBS 0.007832f
C566 B.n474 VSUBS 0.007832f
C567 B.n475 VSUBS 0.007832f
C568 B.n476 VSUBS 0.007832f
C569 B.n477 VSUBS 0.007832f
C570 B.n478 VSUBS 0.007832f
C571 B.n479 VSUBS 0.007832f
C572 B.n480 VSUBS 0.007832f
C573 B.n481 VSUBS 0.007832f
C574 B.n482 VSUBS 0.007832f
C575 B.n483 VSUBS 0.007832f
C576 B.n484 VSUBS 0.007832f
C577 B.n485 VSUBS 0.007832f
C578 B.n486 VSUBS 0.007832f
C579 B.n487 VSUBS 0.007832f
C580 B.n488 VSUBS 0.007832f
C581 B.n489 VSUBS 0.007832f
C582 B.n490 VSUBS 0.007832f
C583 B.n491 VSUBS 0.007832f
C584 B.n492 VSUBS 0.007832f
C585 B.n493 VSUBS 0.007832f
C586 B.n494 VSUBS 0.007832f
C587 B.n495 VSUBS 0.007832f
C588 B.n496 VSUBS 0.007832f
C589 B.n497 VSUBS 0.007832f
C590 B.n498 VSUBS 0.007832f
C591 B.n499 VSUBS 0.007832f
C592 B.n500 VSUBS 0.007832f
C593 B.n501 VSUBS 0.007832f
C594 B.n502 VSUBS 0.007832f
C595 B.n503 VSUBS 0.007832f
C596 B.n504 VSUBS 0.007832f
C597 B.n505 VSUBS 0.007832f
C598 B.n506 VSUBS 0.007832f
C599 B.n507 VSUBS 0.007832f
C600 B.n508 VSUBS 0.007832f
C601 B.n509 VSUBS 0.007832f
C602 B.n510 VSUBS 0.007832f
C603 B.n511 VSUBS 0.007832f
C604 B.n512 VSUBS 0.007832f
C605 B.n513 VSUBS 0.007832f
C606 B.n514 VSUBS 0.007832f
C607 B.n515 VSUBS 0.007832f
C608 B.n516 VSUBS 0.007832f
C609 B.n517 VSUBS 0.007832f
C610 B.n518 VSUBS 0.007832f
C611 B.n519 VSUBS 0.007832f
C612 B.n520 VSUBS 0.007832f
C613 B.n521 VSUBS 0.007832f
C614 B.n522 VSUBS 0.007832f
C615 B.n523 VSUBS 0.007832f
C616 B.n524 VSUBS 0.007832f
C617 B.n525 VSUBS 0.007832f
C618 B.n526 VSUBS 0.007832f
C619 B.n527 VSUBS 0.007832f
C620 B.n528 VSUBS 0.007832f
C621 B.n529 VSUBS 0.007832f
C622 B.n530 VSUBS 0.007832f
C623 B.n531 VSUBS 0.007832f
C624 B.n532 VSUBS 0.007832f
C625 B.n533 VSUBS 0.007832f
C626 B.n534 VSUBS 0.007832f
C627 B.n535 VSUBS 0.007832f
C628 B.n536 VSUBS 0.007832f
C629 B.n537 VSUBS 0.007832f
C630 B.n538 VSUBS 0.007832f
C631 B.n539 VSUBS 0.007832f
C632 B.n540 VSUBS 0.007832f
C633 B.n541 VSUBS 0.007832f
C634 B.n542 VSUBS 0.007832f
C635 B.n543 VSUBS 0.007832f
C636 B.n544 VSUBS 0.007832f
C637 B.n545 VSUBS 0.007832f
C638 B.n546 VSUBS 0.007832f
C639 B.n547 VSUBS 0.007832f
C640 B.n548 VSUBS 0.007832f
C641 B.n549 VSUBS 0.007832f
C642 B.n550 VSUBS 0.007832f
C643 B.n551 VSUBS 0.007832f
C644 B.n552 VSUBS 0.007832f
C645 B.n553 VSUBS 0.007832f
C646 B.n554 VSUBS 0.007832f
C647 B.n555 VSUBS 0.007832f
C648 B.n556 VSUBS 0.007832f
C649 B.n557 VSUBS 0.007832f
C650 B.n558 VSUBS 0.007832f
C651 B.n559 VSUBS 0.007832f
C652 B.n560 VSUBS 0.007832f
C653 B.n561 VSUBS 0.007832f
C654 B.n562 VSUBS 0.007832f
C655 B.n563 VSUBS 0.007832f
C656 B.n564 VSUBS 0.007832f
C657 B.n565 VSUBS 0.007832f
C658 B.n566 VSUBS 0.007832f
C659 B.n567 VSUBS 0.007832f
C660 B.n568 VSUBS 0.007832f
C661 B.n569 VSUBS 0.007832f
C662 B.n570 VSUBS 0.007832f
C663 B.n571 VSUBS 0.007832f
C664 B.n572 VSUBS 0.007832f
C665 B.n573 VSUBS 0.007832f
C666 B.n574 VSUBS 0.007832f
C667 B.n575 VSUBS 0.007832f
C668 B.n576 VSUBS 0.007832f
C669 B.n577 VSUBS 0.007832f
C670 B.n578 VSUBS 0.007832f
C671 B.n579 VSUBS 0.007832f
C672 B.n580 VSUBS 0.007832f
C673 B.n581 VSUBS 0.007832f
C674 B.n582 VSUBS 0.007832f
C675 B.n583 VSUBS 0.007832f
C676 B.n584 VSUBS 0.007832f
C677 B.n585 VSUBS 0.007832f
C678 B.n586 VSUBS 0.007832f
C679 B.n587 VSUBS 0.007832f
C680 B.n588 VSUBS 0.007832f
C681 B.n589 VSUBS 0.007832f
C682 B.n590 VSUBS 0.007832f
C683 B.n591 VSUBS 0.007832f
C684 B.n592 VSUBS 0.007832f
C685 B.n593 VSUBS 0.007832f
C686 B.n594 VSUBS 0.007832f
C687 B.n595 VSUBS 0.007832f
C688 B.n596 VSUBS 0.007832f
C689 B.n597 VSUBS 0.007832f
C690 B.n598 VSUBS 0.007832f
C691 B.n599 VSUBS 0.007832f
C692 B.n600 VSUBS 0.007832f
C693 B.n601 VSUBS 0.007832f
C694 B.n602 VSUBS 0.007832f
C695 B.n603 VSUBS 0.007832f
C696 B.n604 VSUBS 0.007832f
C697 B.n605 VSUBS 0.007832f
C698 B.n606 VSUBS 0.007832f
C699 B.n607 VSUBS 0.007832f
C700 B.n608 VSUBS 0.007832f
C701 B.n609 VSUBS 0.007832f
C702 B.n610 VSUBS 0.007832f
C703 B.n611 VSUBS 0.007832f
C704 B.n612 VSUBS 0.007832f
C705 B.n613 VSUBS 0.007832f
C706 B.n614 VSUBS 0.007832f
C707 B.n615 VSUBS 0.007832f
C708 B.n616 VSUBS 0.007832f
C709 B.n617 VSUBS 0.007832f
C710 B.n618 VSUBS 0.007832f
C711 B.n619 VSUBS 0.017579f
C712 B.n620 VSUBS 0.019048f
C713 B.n621 VSUBS 0.019048f
C714 B.n622 VSUBS 0.007832f
C715 B.n623 VSUBS 0.007832f
C716 B.n624 VSUBS 0.007832f
C717 B.n625 VSUBS 0.007832f
C718 B.n626 VSUBS 0.007832f
C719 B.n627 VSUBS 0.007832f
C720 B.n628 VSUBS 0.007832f
C721 B.n629 VSUBS 0.007832f
C722 B.n630 VSUBS 0.007832f
C723 B.n631 VSUBS 0.007832f
C724 B.n632 VSUBS 0.007832f
C725 B.n633 VSUBS 0.007832f
C726 B.n634 VSUBS 0.007832f
C727 B.n635 VSUBS 0.007832f
C728 B.n636 VSUBS 0.007832f
C729 B.n637 VSUBS 0.007832f
C730 B.n638 VSUBS 0.007832f
C731 B.n639 VSUBS 0.007832f
C732 B.n640 VSUBS 0.007832f
C733 B.n641 VSUBS 0.007832f
C734 B.n642 VSUBS 0.007832f
C735 B.n643 VSUBS 0.007832f
C736 B.n644 VSUBS 0.007832f
C737 B.n645 VSUBS 0.007832f
C738 B.n646 VSUBS 0.007832f
C739 B.n647 VSUBS 0.007832f
C740 B.n648 VSUBS 0.007832f
C741 B.n649 VSUBS 0.007832f
C742 B.n650 VSUBS 0.007832f
C743 B.n651 VSUBS 0.007832f
C744 B.n652 VSUBS 0.007832f
C745 B.n653 VSUBS 0.007832f
C746 B.n654 VSUBS 0.007832f
C747 B.n655 VSUBS 0.007832f
C748 B.n656 VSUBS 0.007832f
C749 B.n657 VSUBS 0.007832f
C750 B.n658 VSUBS 0.007832f
C751 B.n659 VSUBS 0.007832f
C752 B.n660 VSUBS 0.007832f
C753 B.n661 VSUBS 0.007832f
C754 B.n662 VSUBS 0.007832f
C755 B.n663 VSUBS 0.007832f
C756 B.n664 VSUBS 0.007832f
C757 B.n665 VSUBS 0.007832f
C758 B.n666 VSUBS 0.007832f
C759 B.n667 VSUBS 0.007832f
C760 B.n668 VSUBS 0.007832f
C761 B.n669 VSUBS 0.007832f
C762 B.n670 VSUBS 0.007832f
C763 B.n671 VSUBS 0.007832f
C764 B.n672 VSUBS 0.007832f
C765 B.n673 VSUBS 0.007832f
C766 B.n674 VSUBS 0.007832f
C767 B.n675 VSUBS 0.007832f
C768 B.n676 VSUBS 0.007832f
C769 B.n677 VSUBS 0.007832f
C770 B.n678 VSUBS 0.007832f
C771 B.n679 VSUBS 0.007832f
C772 B.n680 VSUBS 0.007832f
C773 B.n681 VSUBS 0.007832f
C774 B.n682 VSUBS 0.007832f
C775 B.n683 VSUBS 0.007832f
C776 B.n684 VSUBS 0.007832f
C777 B.n685 VSUBS 0.007832f
C778 B.n686 VSUBS 0.007832f
C779 B.n687 VSUBS 0.007832f
C780 B.n688 VSUBS 0.007832f
C781 B.n689 VSUBS 0.007832f
C782 B.n690 VSUBS 0.007832f
C783 B.n691 VSUBS 0.007832f
C784 B.n692 VSUBS 0.007832f
C785 B.n693 VSUBS 0.007832f
C786 B.n694 VSUBS 0.007832f
C787 B.n695 VSUBS 0.007832f
C788 B.n696 VSUBS 0.007371f
C789 B.n697 VSUBS 0.018146f
C790 B.n698 VSUBS 0.004377f
C791 B.n699 VSUBS 0.007832f
C792 B.n700 VSUBS 0.007832f
C793 B.n701 VSUBS 0.007832f
C794 B.n702 VSUBS 0.007832f
C795 B.n703 VSUBS 0.007832f
C796 B.n704 VSUBS 0.007832f
C797 B.n705 VSUBS 0.007832f
C798 B.n706 VSUBS 0.007832f
C799 B.n707 VSUBS 0.007832f
C800 B.n708 VSUBS 0.007832f
C801 B.n709 VSUBS 0.007832f
C802 B.n710 VSUBS 0.007832f
C803 B.n711 VSUBS 0.004377f
C804 B.n712 VSUBS 0.007832f
C805 B.n713 VSUBS 0.007832f
C806 B.n714 VSUBS 0.007832f
C807 B.n715 VSUBS 0.007832f
C808 B.n716 VSUBS 0.007832f
C809 B.n717 VSUBS 0.007832f
C810 B.n718 VSUBS 0.007832f
C811 B.n719 VSUBS 0.007832f
C812 B.n720 VSUBS 0.007832f
C813 B.n721 VSUBS 0.007832f
C814 B.n722 VSUBS 0.007832f
C815 B.n723 VSUBS 0.007832f
C816 B.n724 VSUBS 0.007832f
C817 B.n725 VSUBS 0.007832f
C818 B.n726 VSUBS 0.007832f
C819 B.n727 VSUBS 0.007832f
C820 B.n728 VSUBS 0.007832f
C821 B.n729 VSUBS 0.007832f
C822 B.n730 VSUBS 0.007832f
C823 B.n731 VSUBS 0.007832f
C824 B.n732 VSUBS 0.007832f
C825 B.n733 VSUBS 0.007832f
C826 B.n734 VSUBS 0.007832f
C827 B.n735 VSUBS 0.007832f
C828 B.n736 VSUBS 0.007832f
C829 B.n737 VSUBS 0.007832f
C830 B.n738 VSUBS 0.007832f
C831 B.n739 VSUBS 0.007832f
C832 B.n740 VSUBS 0.007832f
C833 B.n741 VSUBS 0.007832f
C834 B.n742 VSUBS 0.007832f
C835 B.n743 VSUBS 0.007832f
C836 B.n744 VSUBS 0.007832f
C837 B.n745 VSUBS 0.007832f
C838 B.n746 VSUBS 0.007832f
C839 B.n747 VSUBS 0.007832f
C840 B.n748 VSUBS 0.007832f
C841 B.n749 VSUBS 0.007832f
C842 B.n750 VSUBS 0.007832f
C843 B.n751 VSUBS 0.007832f
C844 B.n752 VSUBS 0.007832f
C845 B.n753 VSUBS 0.007832f
C846 B.n754 VSUBS 0.007832f
C847 B.n755 VSUBS 0.007832f
C848 B.n756 VSUBS 0.007832f
C849 B.n757 VSUBS 0.007832f
C850 B.n758 VSUBS 0.007832f
C851 B.n759 VSUBS 0.007832f
C852 B.n760 VSUBS 0.007832f
C853 B.n761 VSUBS 0.007832f
C854 B.n762 VSUBS 0.007832f
C855 B.n763 VSUBS 0.007832f
C856 B.n764 VSUBS 0.007832f
C857 B.n765 VSUBS 0.007832f
C858 B.n766 VSUBS 0.007832f
C859 B.n767 VSUBS 0.007832f
C860 B.n768 VSUBS 0.007832f
C861 B.n769 VSUBS 0.007832f
C862 B.n770 VSUBS 0.007832f
C863 B.n771 VSUBS 0.007832f
C864 B.n772 VSUBS 0.007832f
C865 B.n773 VSUBS 0.007832f
C866 B.n774 VSUBS 0.007832f
C867 B.n775 VSUBS 0.007832f
C868 B.n776 VSUBS 0.007832f
C869 B.n777 VSUBS 0.007832f
C870 B.n778 VSUBS 0.007832f
C871 B.n779 VSUBS 0.007832f
C872 B.n780 VSUBS 0.007832f
C873 B.n781 VSUBS 0.007832f
C874 B.n782 VSUBS 0.007832f
C875 B.n783 VSUBS 0.007832f
C876 B.n784 VSUBS 0.007832f
C877 B.n785 VSUBS 0.007832f
C878 B.n786 VSUBS 0.007832f
C879 B.n787 VSUBS 0.007832f
C880 B.n788 VSUBS 0.019048f
C881 B.n789 VSUBS 0.017579f
C882 B.n790 VSUBS 0.017579f
C883 B.n791 VSUBS 0.007832f
C884 B.n792 VSUBS 0.007832f
C885 B.n793 VSUBS 0.007832f
C886 B.n794 VSUBS 0.007832f
C887 B.n795 VSUBS 0.007832f
C888 B.n796 VSUBS 0.007832f
C889 B.n797 VSUBS 0.007832f
C890 B.n798 VSUBS 0.007832f
C891 B.n799 VSUBS 0.007832f
C892 B.n800 VSUBS 0.007832f
C893 B.n801 VSUBS 0.007832f
C894 B.n802 VSUBS 0.007832f
C895 B.n803 VSUBS 0.007832f
C896 B.n804 VSUBS 0.007832f
C897 B.n805 VSUBS 0.007832f
C898 B.n806 VSUBS 0.007832f
C899 B.n807 VSUBS 0.007832f
C900 B.n808 VSUBS 0.007832f
C901 B.n809 VSUBS 0.007832f
C902 B.n810 VSUBS 0.007832f
C903 B.n811 VSUBS 0.007832f
C904 B.n812 VSUBS 0.007832f
C905 B.n813 VSUBS 0.007832f
C906 B.n814 VSUBS 0.007832f
C907 B.n815 VSUBS 0.007832f
C908 B.n816 VSUBS 0.007832f
C909 B.n817 VSUBS 0.007832f
C910 B.n818 VSUBS 0.007832f
C911 B.n819 VSUBS 0.007832f
C912 B.n820 VSUBS 0.007832f
C913 B.n821 VSUBS 0.007832f
C914 B.n822 VSUBS 0.007832f
C915 B.n823 VSUBS 0.007832f
C916 B.n824 VSUBS 0.007832f
C917 B.n825 VSUBS 0.007832f
C918 B.n826 VSUBS 0.007832f
C919 B.n827 VSUBS 0.007832f
C920 B.n828 VSUBS 0.007832f
C921 B.n829 VSUBS 0.007832f
C922 B.n830 VSUBS 0.007832f
C923 B.n831 VSUBS 0.007832f
C924 B.n832 VSUBS 0.007832f
C925 B.n833 VSUBS 0.007832f
C926 B.n834 VSUBS 0.007832f
C927 B.n835 VSUBS 0.007832f
C928 B.n836 VSUBS 0.007832f
C929 B.n837 VSUBS 0.007832f
C930 B.n838 VSUBS 0.007832f
C931 B.n839 VSUBS 0.007832f
C932 B.n840 VSUBS 0.007832f
C933 B.n841 VSUBS 0.007832f
C934 B.n842 VSUBS 0.007832f
C935 B.n843 VSUBS 0.007832f
C936 B.n844 VSUBS 0.007832f
C937 B.n845 VSUBS 0.007832f
C938 B.n846 VSUBS 0.007832f
C939 B.n847 VSUBS 0.007832f
C940 B.n848 VSUBS 0.007832f
C941 B.n849 VSUBS 0.007832f
C942 B.n850 VSUBS 0.007832f
C943 B.n851 VSUBS 0.007832f
C944 B.n852 VSUBS 0.007832f
C945 B.n853 VSUBS 0.007832f
C946 B.n854 VSUBS 0.007832f
C947 B.n855 VSUBS 0.007832f
C948 B.n856 VSUBS 0.007832f
C949 B.n857 VSUBS 0.007832f
C950 B.n858 VSUBS 0.007832f
C951 B.n859 VSUBS 0.007832f
C952 B.n860 VSUBS 0.007832f
C953 B.n861 VSUBS 0.007832f
C954 B.n862 VSUBS 0.007832f
C955 B.n863 VSUBS 0.010221f
C956 B.n864 VSUBS 0.010887f
C957 B.n865 VSUBS 0.021651f
C958 VTAIL.t4 VSUBS 0.344498f
C959 VTAIL.t2 VSUBS 0.344498f
C960 VTAIL.n0 VSUBS 2.66404f
C961 VTAIL.n1 VSUBS 0.912999f
C962 VTAIL.t9 VSUBS 3.48712f
C963 VTAIL.n2 VSUBS 1.24038f
C964 VTAIL.t10 VSUBS 0.344498f
C965 VTAIL.t11 VSUBS 0.344498f
C966 VTAIL.n3 VSUBS 2.66404f
C967 VTAIL.n4 VSUBS 3.11366f
C968 VTAIL.t3 VSUBS 0.344498f
C969 VTAIL.t1 VSUBS 0.344498f
C970 VTAIL.n5 VSUBS 2.66405f
C971 VTAIL.n6 VSUBS 3.11365f
C972 VTAIL.t0 VSUBS 3.48712f
C973 VTAIL.n7 VSUBS 1.24038f
C974 VTAIL.t8 VSUBS 0.344498f
C975 VTAIL.t6 VSUBS 0.344498f
C976 VTAIL.n8 VSUBS 2.66405f
C977 VTAIL.n9 VSUBS 1.12392f
C978 VTAIL.t7 VSUBS 3.48712f
C979 VTAIL.n10 VSUBS 2.94172f
C980 VTAIL.t5 VSUBS 3.48712f
C981 VTAIL.n11 VSUBS 2.86424f
C982 VDD1.t0 VSUBS 3.55078f
C983 VDD1.t5 VSUBS 3.54933f
C984 VDD1.t3 VSUBS 0.331747f
C985 VDD1.t2 VSUBS 0.331747f
C986 VDD1.n0 VSUBS 2.72096f
C987 VDD1.n1 VSUBS 4.50501f
C988 VDD1.t4 VSUBS 0.331747f
C989 VDD1.t1 VSUBS 0.331747f
C990 VDD1.n2 VSUBS 2.71257f
C991 VDD1.n3 VSUBS 3.85115f
C992 VP.t2 VSUBS 3.7415f
C993 VP.n0 VSUBS 1.41274f
C994 VP.n1 VSUBS 0.027296f
C995 VP.n2 VSUBS 0.023325f
C996 VP.n3 VSUBS 0.027296f
C997 VP.t0 VSUBS 3.7415f
C998 VP.n4 VSUBS 1.30012f
C999 VP.n5 VSUBS 0.027296f
C1000 VP.n6 VSUBS 0.023325f
C1001 VP.n7 VSUBS 0.027296f
C1002 VP.t1 VSUBS 3.7415f
C1003 VP.n8 VSUBS 1.41274f
C1004 VP.t4 VSUBS 3.7415f
C1005 VP.n9 VSUBS 1.41274f
C1006 VP.n10 VSUBS 0.027296f
C1007 VP.n11 VSUBS 0.023325f
C1008 VP.n12 VSUBS 0.027296f
C1009 VP.t5 VSUBS 3.7415f
C1010 VP.n13 VSUBS 1.39044f
C1011 VP.t3 VSUBS 4.08654f
C1012 VP.n14 VSUBS 1.3289f
C1013 VP.n15 VSUBS 0.318329f
C1014 VP.n16 VSUBS 0.038123f
C1015 VP.n17 VSUBS 0.050618f
C1016 VP.n18 VSUBS 0.054858f
C1017 VP.n19 VSUBS 0.027296f
C1018 VP.n20 VSUBS 0.027296f
C1019 VP.n21 VSUBS 0.027296f
C1020 VP.n22 VSUBS 0.051792f
C1021 VP.n23 VSUBS 0.050618f
C1022 VP.n24 VSUBS 0.044121f
C1023 VP.n25 VSUBS 0.044048f
C1024 VP.n26 VSUBS 1.72695f
C1025 VP.n27 VSUBS 1.74518f
C1026 VP.n28 VSUBS 0.044048f
C1027 VP.n29 VSUBS 0.044121f
C1028 VP.n30 VSUBS 0.050618f
C1029 VP.n31 VSUBS 0.051792f
C1030 VP.n32 VSUBS 0.027296f
C1031 VP.n33 VSUBS 0.027296f
C1032 VP.n34 VSUBS 0.027296f
C1033 VP.n35 VSUBS 0.054858f
C1034 VP.n36 VSUBS 0.050618f
C1035 VP.n37 VSUBS 0.038123f
C1036 VP.n38 VSUBS 0.027296f
C1037 VP.n39 VSUBS 0.027296f
C1038 VP.n40 VSUBS 0.038123f
C1039 VP.n41 VSUBS 0.050618f
C1040 VP.n42 VSUBS 0.054858f
C1041 VP.n43 VSUBS 0.027296f
C1042 VP.n44 VSUBS 0.027296f
C1043 VP.n45 VSUBS 0.027296f
C1044 VP.n46 VSUBS 0.051792f
C1045 VP.n47 VSUBS 0.050618f
C1046 VP.n48 VSUBS 0.044121f
C1047 VP.n49 VSUBS 0.044048f
C1048 VP.n50 VSUBS 0.061849f
.ends

