* NGSPICE file created from tg_sample_0006.ext - technology: sky130A

.subckt tg_sample_0006 VIN VGN VGP VSS VCC VOUT
X0 VIN.t6 VGN.t0 VOUT.t5 VSS.t11 sky130_fd_pr__nfet_01v8 ad=1.3455 pd=7.68 as=0.56925 ps=3.78 w=3.45 l=0.62
X1 VIN.t1 VGP.t0 VOUT.t1 VCC.t11 sky130_fd_pr__pfet_01v8 ad=7.332 pd=38.38 as=3.102 ps=19.13 w=18.8 l=2.6
X2 VOUT.t7 VGP.t1 VIN.t7 VCC.t10 sky130_fd_pr__pfet_01v8 ad=3.102 pd=19.13 as=3.102 ps=19.13 w=18.8 l=2.6
X3 VSS.t7 VSS.t4 VSS.t6 VSS.t5 sky130_fd_pr__nfet_01v8 ad=1.3455 pd=7.68 as=0 ps=0 w=3.45 l=0.62
X4 VOUT.t6 VGN.t1 VIN.t5 VSS.t10 sky130_fd_pr__nfet_01v8 ad=0.56925 pd=3.78 as=1.3455 ps=7.68 w=3.45 l=0.62
X5 VCC.t7 VCC.t4 VCC.t6 VCC.t5 sky130_fd_pr__pfet_01v8 ad=7.332 pd=38.38 as=0 ps=0 w=18.8 l=2.6
X6 VIN.t4 VGN.t2 VOUT.t3 VSS.t9 sky130_fd_pr__nfet_01v8 ad=0.56925 pd=3.78 as=0.56925 ps=3.78 w=3.45 l=0.62
X7 VSS.t3 VSS.t0 VSS.t2 VSS.t1 sky130_fd_pr__nfet_01v8 ad=1.3455 pd=7.68 as=0 ps=0 w=3.45 l=0.62
X8 VOUT.t2 VGP.t2 VIN.t2 VCC.t9 sky130_fd_pr__pfet_01v8 ad=3.102 pd=19.13 as=7.332 ps=38.38 w=18.8 l=2.6
X9 VOUT.t4 VGN.t3 VIN.t3 VSS.t8 sky130_fd_pr__nfet_01v8 ad=0.56925 pd=3.78 as=0.56925 ps=3.78 w=3.45 l=0.62
X10 VCC.t3 VCC.t0 VCC.t2 VCC.t1 sky130_fd_pr__pfet_01v8 ad=7.332 pd=38.38 as=0 ps=0 w=18.8 l=2.6
X11 VIN.t0 VGP.t3 VOUT.t0 VCC.t8 sky130_fd_pr__pfet_01v8 ad=3.102 pd=19.13 as=3.102 ps=19.13 w=18.8 l=2.6
R0 VGN.n1 VGN.t1 224.674
R1 VGN.n2 VGN.t2 197.853
R2 VGN.n3 VGN.t3 197.853
R3 VGN.n4 VGN.t0 197.853
R4 VGN.n5 VGN.n4 161.3
R5 VGN.n3 VGN.n0 80.6037
R6 VGN.n3 VGN.n2 48.2005
R7 VGN.n4 VGN.n3 48.2005
R8 VGN.n1 VGN.n0 45.2318
R9 VGN.n2 VGN.n1 13.3799
R10 VGN.n5 VGN.n0 0.285035
R11 VGN VGN.n5 0.133076
R12 VOUT.n5 VOUT.n3 75.5978
R13 VOUT.n5 VOUT.n4 74.7788
R14 VOUT.n2 VOUT.n0 74.491
R15 VOUT.n2 VOUT.n1 71.965
R16 VOUT VOUT.n5 12.8798
R17 VOUT.n4 VOUT.t3 5.73963
R18 VOUT.n4 VOUT.t6 5.73963
R19 VOUT.n3 VOUT.t5 5.73963
R20 VOUT.n3 VOUT.t4 5.73963
R21 VOUT.n1 VOUT.t0 1.72949
R22 VOUT.n1 VOUT.t2 1.72949
R23 VOUT.n0 VOUT.t1 1.72949
R24 VOUT.n0 VOUT.t7 1.72949
R25 VOUT VOUT.n2 1.38412
R26 VIN.n102 VIN.n101 756.745
R27 VIN.n207 VIN.n206 756.745
R28 VIN.n35 VIN.n34 585
R29 VIN.n37 VIN.n36 585
R30 VIN.n30 VIN.n29 585
R31 VIN.n43 VIN.n42 585
R32 VIN.n45 VIN.n44 585
R33 VIN.n26 VIN.n25 585
R34 VIN.n52 VIN.n51 585
R35 VIN.n53 VIN.n24 585
R36 VIN.n55 VIN.n54 585
R37 VIN.n22 VIN.n21 585
R38 VIN.n61 VIN.n60 585
R39 VIN.n63 VIN.n62 585
R40 VIN.n18 VIN.n17 585
R41 VIN.n69 VIN.n68 585
R42 VIN.n71 VIN.n70 585
R43 VIN.n14 VIN.n13 585
R44 VIN.n77 VIN.n76 585
R45 VIN.n79 VIN.n78 585
R46 VIN.n10 VIN.n9 585
R47 VIN.n85 VIN.n84 585
R48 VIN.n87 VIN.n86 585
R49 VIN.n6 VIN.n5 585
R50 VIN.n93 VIN.n92 585
R51 VIN.n95 VIN.n94 585
R52 VIN.n2 VIN.n1 585
R53 VIN.n101 VIN.n100 585
R54 VIN.n140 VIN.n139 585
R55 VIN.n142 VIN.n141 585
R56 VIN.n135 VIN.n134 585
R57 VIN.n148 VIN.n147 585
R58 VIN.n150 VIN.n149 585
R59 VIN.n131 VIN.n130 585
R60 VIN.n157 VIN.n156 585
R61 VIN.n158 VIN.n129 585
R62 VIN.n160 VIN.n159 585
R63 VIN.n127 VIN.n126 585
R64 VIN.n166 VIN.n165 585
R65 VIN.n168 VIN.n167 585
R66 VIN.n123 VIN.n122 585
R67 VIN.n174 VIN.n173 585
R68 VIN.n176 VIN.n175 585
R69 VIN.n119 VIN.n118 585
R70 VIN.n182 VIN.n181 585
R71 VIN.n184 VIN.n183 585
R72 VIN.n115 VIN.n114 585
R73 VIN.n190 VIN.n189 585
R74 VIN.n192 VIN.n191 585
R75 VIN.n111 VIN.n110 585
R76 VIN.n198 VIN.n197 585
R77 VIN.n200 VIN.n199 585
R78 VIN.n107 VIN.n106 585
R79 VIN.n206 VIN.n205 585
R80 VIN.n138 VIN.t1 329.036
R81 VIN.n33 VIN.t2 329.036
R82 VIN.n36 VIN.n35 171.744
R83 VIN.n36 VIN.n29 171.744
R84 VIN.n43 VIN.n29 171.744
R85 VIN.n44 VIN.n43 171.744
R86 VIN.n44 VIN.n25 171.744
R87 VIN.n52 VIN.n25 171.744
R88 VIN.n53 VIN.n52 171.744
R89 VIN.n54 VIN.n53 171.744
R90 VIN.n54 VIN.n21 171.744
R91 VIN.n61 VIN.n21 171.744
R92 VIN.n62 VIN.n61 171.744
R93 VIN.n62 VIN.n17 171.744
R94 VIN.n69 VIN.n17 171.744
R95 VIN.n70 VIN.n69 171.744
R96 VIN.n70 VIN.n13 171.744
R97 VIN.n77 VIN.n13 171.744
R98 VIN.n78 VIN.n77 171.744
R99 VIN.n78 VIN.n9 171.744
R100 VIN.n85 VIN.n9 171.744
R101 VIN.n86 VIN.n85 171.744
R102 VIN.n86 VIN.n5 171.744
R103 VIN.n93 VIN.n5 171.744
R104 VIN.n94 VIN.n93 171.744
R105 VIN.n94 VIN.n1 171.744
R106 VIN.n101 VIN.n1 171.744
R107 VIN.n141 VIN.n140 171.744
R108 VIN.n141 VIN.n134 171.744
R109 VIN.n148 VIN.n134 171.744
R110 VIN.n149 VIN.n148 171.744
R111 VIN.n149 VIN.n130 171.744
R112 VIN.n157 VIN.n130 171.744
R113 VIN.n158 VIN.n157 171.744
R114 VIN.n159 VIN.n158 171.744
R115 VIN.n159 VIN.n126 171.744
R116 VIN.n166 VIN.n126 171.744
R117 VIN.n167 VIN.n166 171.744
R118 VIN.n167 VIN.n122 171.744
R119 VIN.n174 VIN.n122 171.744
R120 VIN.n175 VIN.n174 171.744
R121 VIN.n175 VIN.n118 171.744
R122 VIN.n182 VIN.n118 171.744
R123 VIN.n183 VIN.n182 171.744
R124 VIN.n183 VIN.n114 171.744
R125 VIN.n190 VIN.n114 171.744
R126 VIN.n191 VIN.n190 171.744
R127 VIN.n191 VIN.n110 171.744
R128 VIN.n198 VIN.n110 171.744
R129 VIN.n199 VIN.n198 171.744
R130 VIN.n199 VIN.n106 171.744
R131 VIN.n206 VIN.n106 171.744
R132 VIN.n35 VIN.t2 85.8723
R133 VIN.n140 VIN.t1 85.8723
R134 VIN.n210 VIN.t5 64.658
R135 VIN.n211 VIN.t6 63.8391
R136 VIN.n210 VIN.n209 58.1
R137 VIN.n104 VIN.n103 55.2864
R138 VIN.n104 VIN.n102 38.2021
R139 VIN.n208 VIN.n207 35.6763
R140 VIN.n55 VIN.n22 13.1884
R141 VIN.n160 VIN.n127 13.1884
R142 VIN VIN.n208 13.0781
R143 VIN.n56 VIN.n24 12.8005
R144 VIN.n60 VIN.n59 12.8005
R145 VIN.n100 VIN.n0 12.8005
R146 VIN.n161 VIN.n129 12.8005
R147 VIN.n165 VIN.n164 12.8005
R148 VIN.n205 VIN.n105 12.8005
R149 VIN.n51 VIN.n50 12.0247
R150 VIN.n63 VIN.n20 12.0247
R151 VIN.n99 VIN.n2 12.0247
R152 VIN.n156 VIN.n155 12.0247
R153 VIN.n168 VIN.n125 12.0247
R154 VIN.n204 VIN.n107 12.0247
R155 VIN.n49 VIN.n26 11.249
R156 VIN.n64 VIN.n18 11.249
R157 VIN.n96 VIN.n95 11.249
R158 VIN.n154 VIN.n131 11.249
R159 VIN.n169 VIN.n123 11.249
R160 VIN.n201 VIN.n200 11.249
R161 VIN.n34 VIN.n33 10.7239
R162 VIN.n139 VIN.n138 10.7239
R163 VIN.n46 VIN.n45 10.4732
R164 VIN.n68 VIN.n67 10.4732
R165 VIN.n92 VIN.n4 10.4732
R166 VIN.n151 VIN.n150 10.4732
R167 VIN.n173 VIN.n172 10.4732
R168 VIN.n197 VIN.n109 10.4732
R169 VIN.n42 VIN.n28 9.69747
R170 VIN.n71 VIN.n16 9.69747
R171 VIN.n91 VIN.n6 9.69747
R172 VIN.n147 VIN.n133 9.69747
R173 VIN.n176 VIN.n121 9.69747
R174 VIN.n196 VIN.n111 9.69747
R175 VIN.n98 VIN.n0 9.45567
R176 VIN.n203 VIN.n105 9.45567
R177 VIN.n32 VIN.n31 9.3005
R178 VIN.n39 VIN.n38 9.3005
R179 VIN.n41 VIN.n40 9.3005
R180 VIN.n28 VIN.n27 9.3005
R181 VIN.n47 VIN.n46 9.3005
R182 VIN.n49 VIN.n48 9.3005
R183 VIN.n50 VIN.n23 9.3005
R184 VIN.n57 VIN.n56 9.3005
R185 VIN.n59 VIN.n58 9.3005
R186 VIN.n20 VIN.n19 9.3005
R187 VIN.n65 VIN.n64 9.3005
R188 VIN.n67 VIN.n66 9.3005
R189 VIN.n16 VIN.n15 9.3005
R190 VIN.n73 VIN.n72 9.3005
R191 VIN.n75 VIN.n74 9.3005
R192 VIN.n12 VIN.n11 9.3005
R193 VIN.n81 VIN.n80 9.3005
R194 VIN.n83 VIN.n82 9.3005
R195 VIN.n8 VIN.n7 9.3005
R196 VIN.n89 VIN.n88 9.3005
R197 VIN.n91 VIN.n90 9.3005
R198 VIN.n4 VIN.n3 9.3005
R199 VIN.n97 VIN.n96 9.3005
R200 VIN.n99 VIN.n98 9.3005
R201 VIN.n186 VIN.n185 9.3005
R202 VIN.n188 VIN.n187 9.3005
R203 VIN.n113 VIN.n112 9.3005
R204 VIN.n194 VIN.n193 9.3005
R205 VIN.n196 VIN.n195 9.3005
R206 VIN.n109 VIN.n108 9.3005
R207 VIN.n202 VIN.n201 9.3005
R208 VIN.n204 VIN.n203 9.3005
R209 VIN.n180 VIN.n179 9.3005
R210 VIN.n178 VIN.n177 9.3005
R211 VIN.n121 VIN.n120 9.3005
R212 VIN.n172 VIN.n171 9.3005
R213 VIN.n170 VIN.n169 9.3005
R214 VIN.n125 VIN.n124 9.3005
R215 VIN.n164 VIN.n163 9.3005
R216 VIN.n137 VIN.n136 9.3005
R217 VIN.n144 VIN.n143 9.3005
R218 VIN.n146 VIN.n145 9.3005
R219 VIN.n133 VIN.n132 9.3005
R220 VIN.n152 VIN.n151 9.3005
R221 VIN.n154 VIN.n153 9.3005
R222 VIN.n155 VIN.n128 9.3005
R223 VIN.n162 VIN.n161 9.3005
R224 VIN.n117 VIN.n116 9.3005
R225 VIN.n41 VIN.n30 8.92171
R226 VIN.n72 VIN.n14 8.92171
R227 VIN.n88 VIN.n87 8.92171
R228 VIN.n146 VIN.n135 8.92171
R229 VIN.n177 VIN.n119 8.92171
R230 VIN.n193 VIN.n192 8.92171
R231 VIN.n38 VIN.n37 8.14595
R232 VIN.n76 VIN.n75 8.14595
R233 VIN.n84 VIN.n8 8.14595
R234 VIN.n143 VIN.n142 8.14595
R235 VIN.n181 VIN.n180 8.14595
R236 VIN.n189 VIN.n113 8.14595
R237 VIN.n34 VIN.n32 7.3702
R238 VIN.n79 VIN.n12 7.3702
R239 VIN.n83 VIN.n10 7.3702
R240 VIN.n139 VIN.n137 7.3702
R241 VIN.n184 VIN.n117 7.3702
R242 VIN.n188 VIN.n115 7.3702
R243 VIN.n80 VIN.n79 6.59444
R244 VIN.n80 VIN.n10 6.59444
R245 VIN.n185 VIN.n184 6.59444
R246 VIN.n185 VIN.n115 6.59444
R247 VIN.n37 VIN.n32 5.81868
R248 VIN.n76 VIN.n12 5.81868
R249 VIN.n84 VIN.n83 5.81868
R250 VIN.n142 VIN.n137 5.81868
R251 VIN.n181 VIN.n117 5.81868
R252 VIN.n189 VIN.n188 5.81868
R253 VIN.n209 VIN.t3 5.73963
R254 VIN.n209 VIN.t4 5.73963
R255 VIN.n38 VIN.n30 5.04292
R256 VIN.n75 VIN.n14 5.04292
R257 VIN.n87 VIN.n8 5.04292
R258 VIN.n143 VIN.n135 5.04292
R259 VIN.n180 VIN.n119 5.04292
R260 VIN.n192 VIN.n113 5.04292
R261 VIN.n42 VIN.n41 4.26717
R262 VIN.n72 VIN.n71 4.26717
R263 VIN.n88 VIN.n6 4.26717
R264 VIN.n147 VIN.n146 4.26717
R265 VIN.n177 VIN.n176 4.26717
R266 VIN.n193 VIN.n111 4.26717
R267 VIN.n45 VIN.n28 3.49141
R268 VIN.n68 VIN.n16 3.49141
R269 VIN.n92 VIN.n91 3.49141
R270 VIN.n150 VIN.n133 3.49141
R271 VIN.n173 VIN.n121 3.49141
R272 VIN.n197 VIN.n196 3.49141
R273 VIN.n46 VIN.n26 2.71565
R274 VIN.n67 VIN.n18 2.71565
R275 VIN.n95 VIN.n4 2.71565
R276 VIN.n151 VIN.n131 2.71565
R277 VIN.n172 VIN.n123 2.71565
R278 VIN.n200 VIN.n109 2.71565
R279 VIN.n208 VIN.n104 2.52636
R280 VIN.n33 VIN.n31 2.41282
R281 VIN.n138 VIN.n136 2.41282
R282 VIN.n51 VIN.n49 1.93989
R283 VIN.n64 VIN.n63 1.93989
R284 VIN.n96 VIN.n2 1.93989
R285 VIN.n156 VIN.n154 1.93989
R286 VIN.n169 VIN.n168 1.93989
R287 VIN.n201 VIN.n107 1.93989
R288 VIN.n103 VIN.t7 1.72949
R289 VIN.n103 VIN.t0 1.72949
R290 VIN.n50 VIN.n24 1.16414
R291 VIN.n60 VIN.n20 1.16414
R292 VIN.n100 VIN.n99 1.16414
R293 VIN.n155 VIN.n129 1.16414
R294 VIN.n165 VIN.n125 1.16414
R295 VIN.n205 VIN.n204 1.16414
R296 VIN.n211 VIN.n210 0.819465
R297 VIN.n56 VIN.n55 0.388379
R298 VIN.n59 VIN.n22 0.388379
R299 VIN.n102 VIN.n0 0.388379
R300 VIN.n161 VIN.n160 0.388379
R301 VIN.n164 VIN.n127 0.388379
R302 VIN.n207 VIN.n105 0.388379
R303 VIN.n39 VIN.n31 0.155672
R304 VIN.n40 VIN.n39 0.155672
R305 VIN.n40 VIN.n27 0.155672
R306 VIN.n47 VIN.n27 0.155672
R307 VIN.n48 VIN.n47 0.155672
R308 VIN.n48 VIN.n23 0.155672
R309 VIN.n57 VIN.n23 0.155672
R310 VIN.n58 VIN.n57 0.155672
R311 VIN.n58 VIN.n19 0.155672
R312 VIN.n65 VIN.n19 0.155672
R313 VIN.n66 VIN.n65 0.155672
R314 VIN.n66 VIN.n15 0.155672
R315 VIN.n73 VIN.n15 0.155672
R316 VIN.n74 VIN.n73 0.155672
R317 VIN.n74 VIN.n11 0.155672
R318 VIN.n81 VIN.n11 0.155672
R319 VIN.n82 VIN.n81 0.155672
R320 VIN.n82 VIN.n7 0.155672
R321 VIN.n89 VIN.n7 0.155672
R322 VIN.n90 VIN.n89 0.155672
R323 VIN.n90 VIN.n3 0.155672
R324 VIN.n97 VIN.n3 0.155672
R325 VIN.n98 VIN.n97 0.155672
R326 VIN.n144 VIN.n136 0.155672
R327 VIN.n145 VIN.n144 0.155672
R328 VIN.n145 VIN.n132 0.155672
R329 VIN.n152 VIN.n132 0.155672
R330 VIN.n153 VIN.n152 0.155672
R331 VIN.n153 VIN.n128 0.155672
R332 VIN.n162 VIN.n128 0.155672
R333 VIN.n163 VIN.n162 0.155672
R334 VIN.n163 VIN.n124 0.155672
R335 VIN.n170 VIN.n124 0.155672
R336 VIN.n171 VIN.n170 0.155672
R337 VIN.n171 VIN.n120 0.155672
R338 VIN.n178 VIN.n120 0.155672
R339 VIN.n179 VIN.n178 0.155672
R340 VIN.n179 VIN.n116 0.155672
R341 VIN.n186 VIN.n116 0.155672
R342 VIN.n187 VIN.n186 0.155672
R343 VIN.n187 VIN.n112 0.155672
R344 VIN.n194 VIN.n112 0.155672
R345 VIN.n195 VIN.n194 0.155672
R346 VIN.n195 VIN.n108 0.155672
R347 VIN.n202 VIN.n108 0.155672
R348 VIN.n203 VIN.n202 0.155672
R349 VIN VIN.n211 0.00481034
R350 VSS.n102 VSS.n56 603.013
R351 VSS.n71 VSS.n54 603.013
R352 VSS.n201 VSS.n18 603.013
R353 VSS.n203 VSS.n14 603.013
R354 VSS.n57 VSS.n56 585
R355 VSS.n56 VSS.n55 585
R356 VSS.n107 VSS.n106 585
R357 VSS.n108 VSS.n107 585
R358 VSS.n48 VSS.n47 585
R359 VSS.n49 VSS.n48 585
R360 VSS.n118 VSS.n117 585
R361 VSS.n117 VSS.n116 585
R362 VSS.n45 VSS.n44 585
R363 VSS.n44 VSS.n43 585
R364 VSS.n123 VSS.n122 585
R365 VSS.n124 VSS.n123 585
R366 VSS.n35 VSS.n34 585
R367 VSS.n36 VSS.n35 585
R368 VSS.n134 VSS.n133 585
R369 VSS.n133 VSS.n132 585
R370 VSS.n32 VSS.n31 585
R371 VSS.n31 VSS.n30 585
R372 VSS.n139 VSS.n138 585
R373 VSS.n140 VSS.n139 585
R374 VSS.n29 VSS.n28 585
R375 VSS.n141 VSS.n29 585
R376 VSS.n144 VSS.n143 585
R377 VSS.n143 VSS.n142 585
R378 VSS.n26 VSS.n25 585
R379 VSS.n25 VSS.n24 585
R380 VSS.n149 VSS.n148 585
R381 VSS.n150 VSS.n149 585
R382 VSS.n22 VSS.n21 585
R383 VSS.n151 VSS.n22 585
R384 VSS.n154 VSS.n153 585
R385 VSS.n153 VSS.n152 585
R386 VSS.n19 VSS.n17 585
R387 VSS.n17 VSS.n15 585
R388 VSS.n201 VSS.n200 585
R389 VSS.n202 VSS.n201 585
R390 VSS.n204 VSS.n203 585
R391 VSS.n203 VSS.n202 585
R392 VSS.n13 VSS.n11 585
R393 VSS.n15 VSS.n13 585
R394 VSS.n208 VSS.n10 585
R395 VSS.n152 VSS.n10 585
R396 VSS.n209 VSS.n9 585
R397 VSS.n151 VSS.n9 585
R398 VSS.n210 VSS.n8 585
R399 VSS.n150 VSS.n8 585
R400 VSS.n23 VSS.n6 585
R401 VSS.n24 VSS.n23 585
R402 VSS.n214 VSS.n5 585
R403 VSS.n142 VSS.n5 585
R404 VSS.n215 VSS.n4 585
R405 VSS.n141 VSS.n4 585
R406 VSS.n216 VSS.n3 585
R407 VSS.n140 VSS.n3 585
R408 VSS.n38 VSS.n2 585
R409 VSS.n38 VSS.n30 585
R410 VSS.n131 VSS.n130 585
R411 VSS.n132 VSS.n131 585
R412 VSS.n39 VSS.n37 585
R413 VSS.n37 VSS.n36 585
R414 VSS.n126 VSS.n125 585
R415 VSS.n125 VSS.n124 585
R416 VSS.n42 VSS.n41 585
R417 VSS.n43 VSS.n42 585
R418 VSS.n115 VSS.n114 585
R419 VSS.n116 VSS.n115 585
R420 VSS.n51 VSS.n50 585
R421 VSS.n50 VSS.n49 585
R422 VSS.n110 VSS.n109 585
R423 VSS.n109 VSS.n108 585
R424 VSS.n54 VSS.n53 585
R425 VSS.n55 VSS.n54 585
R426 VSS.n14 VSS.n12 585
R427 VSS.n172 VSS.n170 585
R428 VSS.n174 VSS.n173 585
R429 VSS.n175 VSS.n165 585
R430 VSS.n177 VSS.n176 585
R431 VSS.n179 VSS.n163 585
R432 VSS.n181 VSS.n180 585
R433 VSS.n182 VSS.n162 585
R434 VSS.n184 VSS.n183 585
R435 VSS.n186 VSS.n160 585
R436 VSS.n188 VSS.n187 585
R437 VSS.n189 VSS.n159 585
R438 VSS.n191 VSS.n190 585
R439 VSS.n193 VSS.n158 585
R440 VSS.n194 VSS.n157 585
R441 VSS.n197 VSS.n196 585
R442 VSS.n198 VSS.n18 585
R443 VSS.n18 VSS.n16 585
R444 VSS.n103 VSS.n102 585
R445 VSS.n59 VSS.n58 585
R446 VSS.n99 VSS.n98 585
R447 VSS.n100 VSS.n99 585
R448 VSS.n97 VSS.n67 585
R449 VSS.n96 VSS.n95 585
R450 VSS.n94 VSS.n93 585
R451 VSS.n92 VSS.n91 585
R452 VSS.n90 VSS.n89 585
R453 VSS.n88 VSS.n87 585
R454 VSS.n86 VSS.n85 585
R455 VSS.n84 VSS.n83 585
R456 VSS.n82 VSS.n81 585
R457 VSS.n80 VSS.n79 585
R458 VSS.n78 VSS.n77 585
R459 VSS.n76 VSS.n75 585
R460 VSS.n74 VSS.n73 585
R461 VSS.n72 VSS.n71 585
R462 VSS.n100 VSS.n55 426.336
R463 VSS.n202 VSS.n16 426.336
R464 VSS.n166 VSS.t0 338.18
R465 VSS.n68 VSS.t4 338.18
R466 VSS.n108 VSS.n55 273.293
R467 VSS.n116 VSS.n49 273.293
R468 VSS.n116 VSS.n43 273.293
R469 VSS.n124 VSS.n43 273.293
R470 VSS.n132 VSS.n36 273.293
R471 VSS.n140 VSS.n30 273.293
R472 VSS.n142 VSS.n141 273.293
R473 VSS.n150 VSS.n24 273.293
R474 VSS.n151 VSS.n150 273.293
R475 VSS.n152 VSS.n151 273.293
R476 VSS.n202 VSS.n15 273.293
R477 VSS.n171 VSS.n16 256.663
R478 VSS.n169 VSS.n16 256.663
R479 VSS.n178 VSS.n16 256.663
R480 VSS.n164 VSS.n16 256.663
R481 VSS.n185 VSS.n16 256.663
R482 VSS.n161 VSS.n16 256.663
R483 VSS.n192 VSS.n16 256.663
R484 VSS.n195 VSS.n16 256.663
R485 VSS.n101 VSS.n100 256.663
R486 VSS.n100 VSS.n60 256.663
R487 VSS.n100 VSS.n61 256.663
R488 VSS.n100 VSS.n62 256.663
R489 VSS.n100 VSS.n63 256.663
R490 VSS.n100 VSS.n64 256.663
R491 VSS.n100 VSS.n65 256.663
R492 VSS.n100 VSS.n66 256.663
R493 VSS.n107 VSS.n56 240.244
R494 VSS.n107 VSS.n48 240.244
R495 VSS.n117 VSS.n48 240.244
R496 VSS.n117 VSS.n44 240.244
R497 VSS.n123 VSS.n44 240.244
R498 VSS.n123 VSS.n35 240.244
R499 VSS.n133 VSS.n35 240.244
R500 VSS.n133 VSS.n31 240.244
R501 VSS.n139 VSS.n31 240.244
R502 VSS.n139 VSS.n29 240.244
R503 VSS.n143 VSS.n29 240.244
R504 VSS.n143 VSS.n25 240.244
R505 VSS.n149 VSS.n25 240.244
R506 VSS.n149 VSS.n22 240.244
R507 VSS.n153 VSS.n22 240.244
R508 VSS.n153 VSS.n17 240.244
R509 VSS.n201 VSS.n17 240.244
R510 VSS.n109 VSS.n54 240.244
R511 VSS.n109 VSS.n50 240.244
R512 VSS.n115 VSS.n50 240.244
R513 VSS.n115 VSS.n42 240.244
R514 VSS.n125 VSS.n42 240.244
R515 VSS.n125 VSS.n37 240.244
R516 VSS.n131 VSS.n37 240.244
R517 VSS.n131 VSS.n38 240.244
R518 VSS.n38 VSS.n3 240.244
R519 VSS.n4 VSS.n3 240.244
R520 VSS.n5 VSS.n4 240.244
R521 VSS.n23 VSS.n5 240.244
R522 VSS.n23 VSS.n8 240.244
R523 VSS.n9 VSS.n8 240.244
R524 VSS.n10 VSS.n9 240.244
R525 VSS.n13 VSS.n10 240.244
R526 VSS.n203 VSS.n13 240.244
R527 VSS.n124 VSS.t11 177.641
R528 VSS.t10 VSS.n24 177.641
R529 VSS.n99 VSS.n59 163.367
R530 VSS.n99 VSS.n67 163.367
R531 VSS.n95 VSS.n94 163.367
R532 VSS.n91 VSS.n90 163.367
R533 VSS.n87 VSS.n86 163.367
R534 VSS.n83 VSS.n82 163.367
R535 VSS.n79 VSS.n78 163.367
R536 VSS.n75 VSS.n74 163.367
R537 VSS.n196 VSS.n18 163.367
R538 VSS.n194 VSS.n193 163.367
R539 VSS.n191 VSS.n159 163.367
R540 VSS.n187 VSS.n186 163.367
R541 VSS.n184 VSS.n162 163.367
R542 VSS.n180 VSS.n179 163.367
R543 VSS.n177 VSS.n165 163.367
R544 VSS.n173 VSS.n172 163.367
R545 VSS.n108 VSS.t5 155.776
R546 VSS.t1 VSS.n15 155.776
R547 VSS.n132 VSS.t8 150.311
R548 VSS.n141 VSS.t9 150.311
R549 VSS.t8 VSS.n30 122.981
R550 VSS.t9 VSS.n140 122.981
R551 VSS.t5 VSS.n49 117.516
R552 VSS.n152 VSS.t1 117.516
R553 VSS.t11 VSS.n36 95.6527
R554 VSS.n142 VSS.t10 95.6527
R555 VSS.n166 VSS.t2 92.0917
R556 VSS.n68 VSS.t7 92.0917
R557 VSS.n167 VSS.t3 73.6675
R558 VSS.n69 VSS.t6 73.6675
R559 VSS.n102 VSS.n101 71.676
R560 VSS.n67 VSS.n60 71.676
R561 VSS.n94 VSS.n61 71.676
R562 VSS.n90 VSS.n62 71.676
R563 VSS.n86 VSS.n63 71.676
R564 VSS.n82 VSS.n64 71.676
R565 VSS.n78 VSS.n65 71.676
R566 VSS.n74 VSS.n66 71.676
R567 VSS.n195 VSS.n194 71.676
R568 VSS.n192 VSS.n191 71.676
R569 VSS.n187 VSS.n161 71.676
R570 VSS.n185 VSS.n184 71.676
R571 VSS.n180 VSS.n164 71.676
R572 VSS.n178 VSS.n177 71.676
R573 VSS.n173 VSS.n169 71.676
R574 VSS.n171 VSS.n14 71.676
R575 VSS.n172 VSS.n171 71.676
R576 VSS.n169 VSS.n165 71.676
R577 VSS.n179 VSS.n178 71.676
R578 VSS.n164 VSS.n162 71.676
R579 VSS.n186 VSS.n185 71.676
R580 VSS.n161 VSS.n159 71.676
R581 VSS.n193 VSS.n192 71.676
R582 VSS.n196 VSS.n195 71.676
R583 VSS.n101 VSS.n59 71.676
R584 VSS.n95 VSS.n60 71.676
R585 VSS.n91 VSS.n61 71.676
R586 VSS.n87 VSS.n62 71.676
R587 VSS.n83 VSS.n63 71.676
R588 VSS.n79 VSS.n64 71.676
R589 VSS.n75 VSS.n65 71.676
R590 VSS.n71 VSS.n66 71.676
R591 VSS.n168 VSS.n167 34.3278
R592 VSS.n70 VSS.n69 34.3278
R593 VSS.n199 VSS.n198 30.7676
R594 VSS.n205 VSS.n12 30.7676
R595 VSS.n104 VSS.n103 30.7676
R596 VSS.n72 VSS.n52 30.7676
R597 VSS.n106 VSS.n57 19.3944
R598 VSS.n106 VSS.n47 19.3944
R599 VSS.n118 VSS.n47 19.3944
R600 VSS.n118 VSS.n45 19.3944
R601 VSS.n122 VSS.n45 19.3944
R602 VSS.n122 VSS.n34 19.3944
R603 VSS.n134 VSS.n34 19.3944
R604 VSS.n134 VSS.n32 19.3944
R605 VSS.n138 VSS.n32 19.3944
R606 VSS.n138 VSS.n28 19.3944
R607 VSS.n144 VSS.n28 19.3944
R608 VSS.n144 VSS.n26 19.3944
R609 VSS.n148 VSS.n26 19.3944
R610 VSS.n148 VSS.n21 19.3944
R611 VSS.n154 VSS.n21 19.3944
R612 VSS.n154 VSS.n19 19.3944
R613 VSS.n200 VSS.n19 19.3944
R614 VSS.n110 VSS.n53 19.3944
R615 VSS.n110 VSS.n51 19.3944
R616 VSS.n114 VSS.n51 19.3944
R617 VSS.n114 VSS.n41 19.3944
R618 VSS.n126 VSS.n41 19.3944
R619 VSS.n126 VSS.n39 19.3944
R620 VSS.n130 VSS.n39 19.3944
R621 VSS.n130 VSS.n2 19.3944
R622 VSS.n216 VSS.n2 19.3944
R623 VSS.n216 VSS.n215 19.3944
R624 VSS.n215 VSS.n214 19.3944
R625 VSS.n214 VSS.n6 19.3944
R626 VSS.n210 VSS.n6 19.3944
R627 VSS.n210 VSS.n209 19.3944
R628 VSS.n209 VSS.n208 19.3944
R629 VSS.n208 VSS.n11 19.3944
R630 VSS.n204 VSS.n11 19.3944
R631 VSS.n167 VSS.n166 18.4247
R632 VSS.n69 VSS.n68 18.4247
R633 VSS.n198 VSS.n197 10.6151
R634 VSS.n197 VSS.n157 10.6151
R635 VSS.n158 VSS.n157 10.6151
R636 VSS.n190 VSS.n158 10.6151
R637 VSS.n190 VSS.n189 10.6151
R638 VSS.n189 VSS.n188 10.6151
R639 VSS.n188 VSS.n160 10.6151
R640 VSS.n183 VSS.n160 10.6151
R641 VSS.n183 VSS.n182 10.6151
R642 VSS.n182 VSS.n181 10.6151
R643 VSS.n181 VSS.n163 10.6151
R644 VSS.n176 VSS.n163 10.6151
R645 VSS.n176 VSS.n175 10.6151
R646 VSS.n175 VSS.n174 10.6151
R647 VSS.n170 VSS.n12 10.6151
R648 VSS.n103 VSS.n58 10.6151
R649 VSS.n98 VSS.n58 10.6151
R650 VSS.n98 VSS.n97 10.6151
R651 VSS.n97 VSS.n96 10.6151
R652 VSS.n96 VSS.n93 10.6151
R653 VSS.n93 VSS.n92 10.6151
R654 VSS.n92 VSS.n89 10.6151
R655 VSS.n89 VSS.n88 10.6151
R656 VSS.n88 VSS.n85 10.6151
R657 VSS.n85 VSS.n84 10.6151
R658 VSS.n84 VSS.n81 10.6151
R659 VSS.n81 VSS.n80 10.6151
R660 VSS.n80 VSS.n77 10.6151
R661 VSS.n77 VSS.n76 10.6151
R662 VSS.n73 VSS.n72 10.6151
R663 VSS.n170 VSS.n168 9.67855
R664 VSS.n73 VSS.n70 9.67855
R665 VSS.n215 VSS.n0 9.3005
R666 VSS.n214 VSS.n213 9.3005
R667 VSS.n212 VSS.n6 9.3005
R668 VSS.n211 VSS.n210 9.3005
R669 VSS.n209 VSS.n7 9.3005
R670 VSS.n208 VSS.n207 9.3005
R671 VSS.n206 VSS.n11 9.3005
R672 VSS.n205 VSS.n204 9.3005
R673 VSS.n104 VSS.n57 9.3005
R674 VSS.n106 VSS.n105 9.3005
R675 VSS.n47 VSS.n46 9.3005
R676 VSS.n119 VSS.n118 9.3005
R677 VSS.n120 VSS.n45 9.3005
R678 VSS.n122 VSS.n121 9.3005
R679 VSS.n34 VSS.n33 9.3005
R680 VSS.n135 VSS.n134 9.3005
R681 VSS.n136 VSS.n32 9.3005
R682 VSS.n138 VSS.n137 9.3005
R683 VSS.n28 VSS.n27 9.3005
R684 VSS.n145 VSS.n144 9.3005
R685 VSS.n146 VSS.n26 9.3005
R686 VSS.n148 VSS.n147 9.3005
R687 VSS.n21 VSS.n20 9.3005
R688 VSS.n155 VSS.n154 9.3005
R689 VSS.n156 VSS.n19 9.3005
R690 VSS.n200 VSS.n199 9.3005
R691 VSS.n111 VSS.n110 9.3005
R692 VSS.n112 VSS.n51 9.3005
R693 VSS.n114 VSS.n113 9.3005
R694 VSS.n41 VSS.n40 9.3005
R695 VSS.n127 VSS.n126 9.3005
R696 VSS.n128 VSS.n39 9.3005
R697 VSS.n130 VSS.n129 9.3005
R698 VSS.n2 VSS.n1 9.3005
R699 VSS.n53 VSS.n52 9.3005
R700 VSS VSS.n216 9.3005
R701 VSS.n174 VSS.n168 0.937085
R702 VSS.n76 VSS.n70 0.937085
R703 VSS VSS.n0 0.152939
R704 VSS.n213 VSS.n0 0.152939
R705 VSS.n213 VSS.n212 0.152939
R706 VSS.n212 VSS.n211 0.152939
R707 VSS.n211 VSS.n7 0.152939
R708 VSS.n207 VSS.n7 0.152939
R709 VSS.n207 VSS.n206 0.152939
R710 VSS.n206 VSS.n205 0.152939
R711 VSS.n105 VSS.n104 0.152939
R712 VSS.n105 VSS.n46 0.152939
R713 VSS.n119 VSS.n46 0.152939
R714 VSS.n120 VSS.n119 0.152939
R715 VSS.n121 VSS.n120 0.152939
R716 VSS.n121 VSS.n33 0.152939
R717 VSS.n135 VSS.n33 0.152939
R718 VSS.n136 VSS.n135 0.152939
R719 VSS.n137 VSS.n136 0.152939
R720 VSS.n137 VSS.n27 0.152939
R721 VSS.n145 VSS.n27 0.152939
R722 VSS.n146 VSS.n145 0.152939
R723 VSS.n147 VSS.n146 0.152939
R724 VSS.n147 VSS.n20 0.152939
R725 VSS.n155 VSS.n20 0.152939
R726 VSS.n156 VSS.n155 0.152939
R727 VSS.n199 VSS.n156 0.152939
R728 VSS.n111 VSS.n52 0.152939
R729 VSS.n112 VSS.n111 0.152939
R730 VSS.n113 VSS.n112 0.152939
R731 VSS.n113 VSS.n40 0.152939
R732 VSS.n127 VSS.n40 0.152939
R733 VSS.n128 VSS.n127 0.152939
R734 VSS.n129 VSS.n128 0.152939
R735 VSS.n129 VSS.n1 0.152939
R736 VSS VSS.n1 0.1255
R737 VGP.n7 VGP.t2 207.083
R738 VGP.n8 VGP.t3 174.262
R739 VGP.n3 VGP.t1 174.262
R740 VGP.n27 VGP.t0 174.262
R741 VGP.n26 VGP.n0 161.3
R742 VGP.n25 VGP.n24 161.3
R743 VGP.n23 VGP.n1 161.3
R744 VGP.n22 VGP.n21 161.3
R745 VGP.n20 VGP.n2 161.3
R746 VGP.n19 VGP.n18 161.3
R747 VGP.n17 VGP.n16 161.3
R748 VGP.n15 VGP.n4 161.3
R749 VGP.n14 VGP.n13 161.3
R750 VGP.n12 VGP.n5 161.3
R751 VGP.n11 VGP.n10 161.3
R752 VGP.n9 VGP.n6 161.3
R753 VGP.n28 VGP.n27 103.776
R754 VGP.n8 VGP.n7 61.9251
R755 VGP.n14 VGP.n5 56.5617
R756 VGP.n21 VGP.n1 56.5617
R757 VGP.n10 VGP.n5 24.5923
R758 VGP.n10 VGP.n9 24.5923
R759 VGP.n21 VGP.n20 24.5923
R760 VGP.n20 VGP.n19 24.5923
R761 VGP.n16 VGP.n15 24.5923
R762 VGP.n15 VGP.n14 24.5923
R763 VGP.n26 VGP.n25 24.5923
R764 VGP.n25 VGP.n1 24.5923
R765 VGP.n19 VGP.n3 14.0178
R766 VGP.n9 VGP.n8 10.575
R767 VGP.n16 VGP.n3 10.575
R768 VGP.n27 VGP.n26 7.13213
R769 VGP.n7 VGP.n6 7.0132
R770 VGP.n28 VGP.n0 0.278335
R771 VGP VGP.n28 0.219773
R772 VGP.n24 VGP.n0 0.189894
R773 VGP.n24 VGP.n23 0.189894
R774 VGP.n23 VGP.n22 0.189894
R775 VGP.n22 VGP.n2 0.189894
R776 VGP.n18 VGP.n2 0.189894
R777 VGP.n18 VGP.n17 0.189894
R778 VGP.n17 VGP.n4 0.189894
R779 VGP.n13 VGP.n4 0.189894
R780 VGP.n13 VGP.n12 0.189894
R781 VGP.n12 VGP.n11 0.189894
R782 VGP.n11 VGP.n6 0.189894
R783 VCC.n443 VCC.t2 554.835
R784 VCC.n157 VCC.t7 554.835
R785 VCC.n444 VCC.t3 498.01
R786 VCC.n158 VCC.t6 498.01
R787 VCC.n443 VCC.t0 382.308
R788 VCC.n157 VCC.t4 382.308
R789 VCC.n571 VCC.n29 354.147
R790 VCC.n569 VCC.n33 354.147
R791 VCC.n283 VCC.n126 354.147
R792 VCC.n285 VCC.n124 354.147
R793 VCC.n569 VCC.n568 185
R794 VCC.n570 VCC.n569 185
R795 VCC.n34 VCC.n32 185
R796 VCC.n32 VCC.n30 185
R797 VCC.n409 VCC.n408 185
R798 VCC.n408 VCC.n407 185
R799 VCC.n37 VCC.n36 185
R800 VCC.n406 VCC.n37 185
R801 VCC.n404 VCC.n403 185
R802 VCC.n405 VCC.n404 185
R803 VCC.n41 VCC.n40 185
R804 VCC.n40 VCC.n39 185
R805 VCC.n399 VCC.n398 185
R806 VCC.n398 VCC.n397 185
R807 VCC.n44 VCC.n43 185
R808 VCC.n396 VCC.n44 185
R809 VCC.n394 VCC.n393 185
R810 VCC.n395 VCC.n394 185
R811 VCC.n48 VCC.n47 185
R812 VCC.n47 VCC.n46 185
R813 VCC.n389 VCC.n388 185
R814 VCC.n388 VCC.n387 185
R815 VCC.n51 VCC.n50 185
R816 VCC.n386 VCC.n51 185
R817 VCC.n384 VCC.n383 185
R818 VCC.n385 VCC.n384 185
R819 VCC.n55 VCC.n54 185
R820 VCC.n54 VCC.n53 185
R821 VCC.n379 VCC.n378 185
R822 VCC.n378 VCC.n377 185
R823 VCC.n58 VCC.n57 185
R824 VCC.n376 VCC.n58 185
R825 VCC.n374 VCC.n373 185
R826 VCC.n375 VCC.n374 185
R827 VCC.n62 VCC.n61 185
R828 VCC.n61 VCC.n60 185
R829 VCC.n369 VCC.n368 185
R830 VCC.n368 VCC.n367 185
R831 VCC.n65 VCC.n64 185
R832 VCC.n366 VCC.n65 185
R833 VCC.n364 VCC.n363 185
R834 VCC.n365 VCC.n364 185
R835 VCC.n68 VCC.n67 185
R836 VCC.n67 VCC.n66 185
R837 VCC.n359 VCC.n358 185
R838 VCC.n358 VCC.n357 185
R839 VCC.n71 VCC.n70 185
R840 VCC.n348 VCC.n71 185
R841 VCC.n347 VCC.n346 185
R842 VCC.n349 VCC.n347 185
R843 VCC.n80 VCC.n79 185
R844 VCC.n79 VCC.n78 185
R845 VCC.n342 VCC.n341 185
R846 VCC.n341 VCC.n340 185
R847 VCC.n83 VCC.n82 185
R848 VCC.n84 VCC.n83 185
R849 VCC.n331 VCC.n330 185
R850 VCC.n332 VCC.n331 185
R851 VCC.n91 VCC.n90 185
R852 VCC.n96 VCC.n90 185
R853 VCC.n326 VCC.n325 185
R854 VCC.n325 VCC.n324 185
R855 VCC.n94 VCC.n93 185
R856 VCC.n95 VCC.n94 185
R857 VCC.n315 VCC.n314 185
R858 VCC.n316 VCC.n315 185
R859 VCC.n104 VCC.n103 185
R860 VCC.n103 VCC.n102 185
R861 VCC.n310 VCC.n309 185
R862 VCC.n309 VCC.n308 185
R863 VCC.n107 VCC.n106 185
R864 VCC.n108 VCC.n107 185
R865 VCC.n299 VCC.n298 185
R866 VCC.n300 VCC.n299 185
R867 VCC.n115 VCC.n114 185
R868 VCC.n120 VCC.n114 185
R869 VCC.n294 VCC.n293 185
R870 VCC.n293 VCC.n292 185
R871 VCC.n118 VCC.n117 185
R872 VCC.n119 VCC.n118 185
R873 VCC.n283 VCC.n282 185
R874 VCC.n284 VCC.n283 185
R875 VCC.n286 VCC.n285 185
R876 VCC.n285 VCC.n284 185
R877 VCC.n122 VCC.n121 185
R878 VCC.n121 VCC.n119 185
R879 VCC.n291 VCC.n290 185
R880 VCC.n292 VCC.n291 185
R881 VCC.n113 VCC.n112 185
R882 VCC.n120 VCC.n113 185
R883 VCC.n302 VCC.n301 185
R884 VCC.n301 VCC.n300 185
R885 VCC.n110 VCC.n109 185
R886 VCC.n109 VCC.n108 185
R887 VCC.n307 VCC.n306 185
R888 VCC.n308 VCC.n307 185
R889 VCC.n101 VCC.n100 185
R890 VCC.n102 VCC.n101 185
R891 VCC.n318 VCC.n317 185
R892 VCC.n317 VCC.n316 185
R893 VCC.n98 VCC.n97 185
R894 VCC.n97 VCC.n95 185
R895 VCC.n323 VCC.n322 185
R896 VCC.n324 VCC.n323 185
R897 VCC.n89 VCC.n88 185
R898 VCC.n96 VCC.n89 185
R899 VCC.n334 VCC.n333 185
R900 VCC.n333 VCC.n332 185
R901 VCC.n86 VCC.n85 185
R902 VCC.n85 VCC.n84 185
R903 VCC.n339 VCC.n338 185
R904 VCC.n340 VCC.n339 185
R905 VCC.n77 VCC.n76 185
R906 VCC.n78 VCC.n77 185
R907 VCC.n351 VCC.n350 185
R908 VCC.n350 VCC.n349 185
R909 VCC.n74 VCC.n72 185
R910 VCC.n348 VCC.n72 185
R911 VCC.n356 VCC.n355 185
R912 VCC.n357 VCC.n356 185
R913 VCC.n73 VCC.n2 185
R914 VCC.n73 VCC.n66 185
R915 VCC.n602 VCC.n3 185
R916 VCC.n365 VCC.n3 185
R917 VCC.n601 VCC.n4 185
R918 VCC.n366 VCC.n4 185
R919 VCC.n600 VCC.n5 185
R920 VCC.n367 VCC.n5 185
R921 VCC.n59 VCC.n6 185
R922 VCC.n60 VCC.n59 185
R923 VCC.n596 VCC.n8 185
R924 VCC.n375 VCC.n8 185
R925 VCC.n595 VCC.n9 185
R926 VCC.n376 VCC.n9 185
R927 VCC.n594 VCC.n10 185
R928 VCC.n377 VCC.n10 185
R929 VCC.n52 VCC.n11 185
R930 VCC.n53 VCC.n52 185
R931 VCC.n590 VCC.n13 185
R932 VCC.n385 VCC.n13 185
R933 VCC.n589 VCC.n14 185
R934 VCC.n386 VCC.n14 185
R935 VCC.n588 VCC.n15 185
R936 VCC.n387 VCC.n15 185
R937 VCC.n45 VCC.n16 185
R938 VCC.n46 VCC.n45 185
R939 VCC.n584 VCC.n18 185
R940 VCC.n395 VCC.n18 185
R941 VCC.n583 VCC.n19 185
R942 VCC.n396 VCC.n19 185
R943 VCC.n582 VCC.n20 185
R944 VCC.n397 VCC.n20 185
R945 VCC.n38 VCC.n21 185
R946 VCC.n39 VCC.n38 185
R947 VCC.n578 VCC.n23 185
R948 VCC.n405 VCC.n23 185
R949 VCC.n577 VCC.n24 185
R950 VCC.n406 VCC.n24 185
R951 VCC.n576 VCC.n25 185
R952 VCC.n407 VCC.n25 185
R953 VCC.n28 VCC.n26 185
R954 VCC.n30 VCC.n28 185
R955 VCC.n572 VCC.n571 185
R956 VCC.n571 VCC.n570 185
R957 VCC.n566 VCC.n33 185
R958 VCC.n565 VCC.n564 185
R959 VCC.n562 VCC.n412 185
R960 VCC.n560 VCC.n559 185
R961 VCC.n558 VCC.n413 185
R962 VCC.n557 VCC.n556 185
R963 VCC.n554 VCC.n414 185
R964 VCC.n552 VCC.n551 185
R965 VCC.n550 VCC.n415 185
R966 VCC.n549 VCC.n548 185
R967 VCC.n546 VCC.n416 185
R968 VCC.n544 VCC.n543 185
R969 VCC.n542 VCC.n417 185
R970 VCC.n541 VCC.n540 185
R971 VCC.n538 VCC.n418 185
R972 VCC.n536 VCC.n535 185
R973 VCC.n534 VCC.n419 185
R974 VCC.n533 VCC.n532 185
R975 VCC.n530 VCC.n420 185
R976 VCC.n528 VCC.n527 185
R977 VCC.n526 VCC.n421 185
R978 VCC.n525 VCC.n524 185
R979 VCC.n522 VCC.n422 185
R980 VCC.n520 VCC.n519 185
R981 VCC.n518 VCC.n423 185
R982 VCC.n517 VCC.n516 185
R983 VCC.n514 VCC.n424 185
R984 VCC.n512 VCC.n511 185
R985 VCC.n510 VCC.n425 185
R986 VCC.n509 VCC.n508 185
R987 VCC.n506 VCC.n426 185
R988 VCC.n504 VCC.n503 185
R989 VCC.n502 VCC.n427 185
R990 VCC.n501 VCC.n500 185
R991 VCC.n498 VCC.n428 185
R992 VCC.n496 VCC.n495 185
R993 VCC.n494 VCC.n429 185
R994 VCC.n493 VCC.n492 185
R995 VCC.n490 VCC.n430 185
R996 VCC.n488 VCC.n487 185
R997 VCC.n486 VCC.n431 185
R998 VCC.n485 VCC.n484 185
R999 VCC.n482 VCC.n432 185
R1000 VCC.n480 VCC.n479 185
R1001 VCC.n478 VCC.n433 185
R1002 VCC.n477 VCC.n476 185
R1003 VCC.n474 VCC.n434 185
R1004 VCC.n472 VCC.n471 185
R1005 VCC.n470 VCC.n435 185
R1006 VCC.n469 VCC.n468 185
R1007 VCC.n466 VCC.n436 185
R1008 VCC.n464 VCC.n463 185
R1009 VCC.n462 VCC.n437 185
R1010 VCC.n461 VCC.n460 185
R1011 VCC.n458 VCC.n438 185
R1012 VCC.n456 VCC.n455 185
R1013 VCC.n454 VCC.n439 185
R1014 VCC.n453 VCC.n452 185
R1015 VCC.n450 VCC.n440 185
R1016 VCC.n448 VCC.n447 185
R1017 VCC.n445 VCC.n442 185
R1018 VCC.n29 VCC.n27 185
R1019 VCC.n124 VCC.n123 185
R1020 VCC.n162 VCC.n160 185
R1021 VCC.n163 VCC.n156 185
R1022 VCC.n163 VCC.n125 185
R1023 VCC.n166 VCC.n165 185
R1024 VCC.n167 VCC.n155 185
R1025 VCC.n169 VCC.n168 185
R1026 VCC.n171 VCC.n154 185
R1027 VCC.n174 VCC.n173 185
R1028 VCC.n175 VCC.n153 185
R1029 VCC.n177 VCC.n176 185
R1030 VCC.n179 VCC.n152 185
R1031 VCC.n182 VCC.n181 185
R1032 VCC.n183 VCC.n151 185
R1033 VCC.n185 VCC.n184 185
R1034 VCC.n187 VCC.n150 185
R1035 VCC.n190 VCC.n189 185
R1036 VCC.n191 VCC.n149 185
R1037 VCC.n193 VCC.n192 185
R1038 VCC.n195 VCC.n148 185
R1039 VCC.n198 VCC.n197 185
R1040 VCC.n199 VCC.n147 185
R1041 VCC.n201 VCC.n200 185
R1042 VCC.n203 VCC.n146 185
R1043 VCC.n206 VCC.n205 185
R1044 VCC.n207 VCC.n145 185
R1045 VCC.n209 VCC.n208 185
R1046 VCC.n211 VCC.n144 185
R1047 VCC.n214 VCC.n213 185
R1048 VCC.n215 VCC.n143 185
R1049 VCC.n217 VCC.n216 185
R1050 VCC.n219 VCC.n142 185
R1051 VCC.n222 VCC.n221 185
R1052 VCC.n223 VCC.n141 185
R1053 VCC.n225 VCC.n224 185
R1054 VCC.n227 VCC.n140 185
R1055 VCC.n230 VCC.n229 185
R1056 VCC.n231 VCC.n139 185
R1057 VCC.n233 VCC.n232 185
R1058 VCC.n235 VCC.n138 185
R1059 VCC.n238 VCC.n237 185
R1060 VCC.n239 VCC.n137 185
R1061 VCC.n241 VCC.n240 185
R1062 VCC.n243 VCC.n136 185
R1063 VCC.n246 VCC.n245 185
R1064 VCC.n247 VCC.n135 185
R1065 VCC.n249 VCC.n248 185
R1066 VCC.n251 VCC.n134 185
R1067 VCC.n254 VCC.n253 185
R1068 VCC.n255 VCC.n133 185
R1069 VCC.n257 VCC.n256 185
R1070 VCC.n259 VCC.n132 185
R1071 VCC.n262 VCC.n261 185
R1072 VCC.n263 VCC.n131 185
R1073 VCC.n265 VCC.n264 185
R1074 VCC.n267 VCC.n130 185
R1075 VCC.n270 VCC.n269 185
R1076 VCC.n271 VCC.n129 185
R1077 VCC.n273 VCC.n272 185
R1078 VCC.n275 VCC.n128 185
R1079 VCC.n276 VCC.n127 185
R1080 VCC.n279 VCC.n278 185
R1081 VCC.n280 VCC.n126 185
R1082 VCC.n126 VCC.n125 185
R1083 VCC.n283 VCC.n118 146.341
R1084 VCC.n293 VCC.n118 146.341
R1085 VCC.n293 VCC.n114 146.341
R1086 VCC.n299 VCC.n114 146.341
R1087 VCC.n299 VCC.n107 146.341
R1088 VCC.n309 VCC.n107 146.341
R1089 VCC.n309 VCC.n103 146.341
R1090 VCC.n315 VCC.n103 146.341
R1091 VCC.n315 VCC.n94 146.341
R1092 VCC.n325 VCC.n94 146.341
R1093 VCC.n325 VCC.n90 146.341
R1094 VCC.n331 VCC.n90 146.341
R1095 VCC.n331 VCC.n83 146.341
R1096 VCC.n341 VCC.n83 146.341
R1097 VCC.n341 VCC.n79 146.341
R1098 VCC.n347 VCC.n79 146.341
R1099 VCC.n347 VCC.n71 146.341
R1100 VCC.n358 VCC.n71 146.341
R1101 VCC.n358 VCC.n67 146.341
R1102 VCC.n364 VCC.n67 146.341
R1103 VCC.n364 VCC.n65 146.341
R1104 VCC.n368 VCC.n65 146.341
R1105 VCC.n368 VCC.n61 146.341
R1106 VCC.n374 VCC.n61 146.341
R1107 VCC.n374 VCC.n58 146.341
R1108 VCC.n378 VCC.n58 146.341
R1109 VCC.n378 VCC.n54 146.341
R1110 VCC.n384 VCC.n54 146.341
R1111 VCC.n384 VCC.n51 146.341
R1112 VCC.n388 VCC.n51 146.341
R1113 VCC.n388 VCC.n47 146.341
R1114 VCC.n394 VCC.n47 146.341
R1115 VCC.n394 VCC.n44 146.341
R1116 VCC.n398 VCC.n44 146.341
R1117 VCC.n398 VCC.n40 146.341
R1118 VCC.n404 VCC.n40 146.341
R1119 VCC.n404 VCC.n37 146.341
R1120 VCC.n408 VCC.n37 146.341
R1121 VCC.n408 VCC.n32 146.341
R1122 VCC.n569 VCC.n32 146.341
R1123 VCC.n285 VCC.n121 146.341
R1124 VCC.n291 VCC.n121 146.341
R1125 VCC.n291 VCC.n113 146.341
R1126 VCC.n301 VCC.n113 146.341
R1127 VCC.n301 VCC.n109 146.341
R1128 VCC.n307 VCC.n109 146.341
R1129 VCC.n307 VCC.n101 146.341
R1130 VCC.n317 VCC.n101 146.341
R1131 VCC.n317 VCC.n97 146.341
R1132 VCC.n323 VCC.n97 146.341
R1133 VCC.n323 VCC.n89 146.341
R1134 VCC.n333 VCC.n89 146.341
R1135 VCC.n333 VCC.n85 146.341
R1136 VCC.n339 VCC.n85 146.341
R1137 VCC.n339 VCC.n77 146.341
R1138 VCC.n350 VCC.n77 146.341
R1139 VCC.n350 VCC.n72 146.341
R1140 VCC.n356 VCC.n72 146.341
R1141 VCC.n356 VCC.n73 146.341
R1142 VCC.n73 VCC.n3 146.341
R1143 VCC.n4 VCC.n3 146.341
R1144 VCC.n5 VCC.n4 146.341
R1145 VCC.n59 VCC.n5 146.341
R1146 VCC.n59 VCC.n8 146.341
R1147 VCC.n9 VCC.n8 146.341
R1148 VCC.n10 VCC.n9 146.341
R1149 VCC.n52 VCC.n10 146.341
R1150 VCC.n52 VCC.n13 146.341
R1151 VCC.n14 VCC.n13 146.341
R1152 VCC.n15 VCC.n14 146.341
R1153 VCC.n45 VCC.n15 146.341
R1154 VCC.n45 VCC.n18 146.341
R1155 VCC.n19 VCC.n18 146.341
R1156 VCC.n20 VCC.n19 146.341
R1157 VCC.n38 VCC.n20 146.341
R1158 VCC.n38 VCC.n23 146.341
R1159 VCC.n24 VCC.n23 146.341
R1160 VCC.n25 VCC.n24 146.341
R1161 VCC.n28 VCC.n25 146.341
R1162 VCC.n571 VCC.n28 146.341
R1163 VCC.n448 VCC.n442 99.5127
R1164 VCC.n452 VCC.n450 99.5127
R1165 VCC.n456 VCC.n439 99.5127
R1166 VCC.n460 VCC.n458 99.5127
R1167 VCC.n464 VCC.n437 99.5127
R1168 VCC.n468 VCC.n466 99.5127
R1169 VCC.n472 VCC.n435 99.5127
R1170 VCC.n476 VCC.n474 99.5127
R1171 VCC.n480 VCC.n433 99.5127
R1172 VCC.n484 VCC.n482 99.5127
R1173 VCC.n488 VCC.n431 99.5127
R1174 VCC.n492 VCC.n490 99.5127
R1175 VCC.n496 VCC.n429 99.5127
R1176 VCC.n500 VCC.n498 99.5127
R1177 VCC.n504 VCC.n427 99.5127
R1178 VCC.n508 VCC.n506 99.5127
R1179 VCC.n512 VCC.n425 99.5127
R1180 VCC.n516 VCC.n514 99.5127
R1181 VCC.n520 VCC.n423 99.5127
R1182 VCC.n524 VCC.n522 99.5127
R1183 VCC.n528 VCC.n421 99.5127
R1184 VCC.n532 VCC.n530 99.5127
R1185 VCC.n536 VCC.n419 99.5127
R1186 VCC.n540 VCC.n538 99.5127
R1187 VCC.n544 VCC.n417 99.5127
R1188 VCC.n548 VCC.n546 99.5127
R1189 VCC.n552 VCC.n415 99.5127
R1190 VCC.n556 VCC.n554 99.5127
R1191 VCC.n560 VCC.n413 99.5127
R1192 VCC.n564 VCC.n562 99.5127
R1193 VCC.n163 VCC.n162 99.5127
R1194 VCC.n165 VCC.n163 99.5127
R1195 VCC.n169 VCC.n155 99.5127
R1196 VCC.n173 VCC.n171 99.5127
R1197 VCC.n177 VCC.n153 99.5127
R1198 VCC.n181 VCC.n179 99.5127
R1199 VCC.n185 VCC.n151 99.5127
R1200 VCC.n189 VCC.n187 99.5127
R1201 VCC.n193 VCC.n149 99.5127
R1202 VCC.n197 VCC.n195 99.5127
R1203 VCC.n201 VCC.n147 99.5127
R1204 VCC.n205 VCC.n203 99.5127
R1205 VCC.n209 VCC.n145 99.5127
R1206 VCC.n213 VCC.n211 99.5127
R1207 VCC.n217 VCC.n143 99.5127
R1208 VCC.n221 VCC.n219 99.5127
R1209 VCC.n225 VCC.n141 99.5127
R1210 VCC.n229 VCC.n227 99.5127
R1211 VCC.n233 VCC.n139 99.5127
R1212 VCC.n237 VCC.n235 99.5127
R1213 VCC.n241 VCC.n137 99.5127
R1214 VCC.n245 VCC.n243 99.5127
R1215 VCC.n249 VCC.n135 99.5127
R1216 VCC.n253 VCC.n251 99.5127
R1217 VCC.n257 VCC.n133 99.5127
R1218 VCC.n261 VCC.n259 99.5127
R1219 VCC.n265 VCC.n131 99.5127
R1220 VCC.n269 VCC.n267 99.5127
R1221 VCC.n273 VCC.n129 99.5127
R1222 VCC.n276 VCC.n275 99.5127
R1223 VCC.n278 VCC.n126 99.5127
R1224 VCC.n563 VCC.n31 72.8958
R1225 VCC.n561 VCC.n31 72.8958
R1226 VCC.n555 VCC.n31 72.8958
R1227 VCC.n553 VCC.n31 72.8958
R1228 VCC.n547 VCC.n31 72.8958
R1229 VCC.n545 VCC.n31 72.8958
R1230 VCC.n539 VCC.n31 72.8958
R1231 VCC.n537 VCC.n31 72.8958
R1232 VCC.n531 VCC.n31 72.8958
R1233 VCC.n529 VCC.n31 72.8958
R1234 VCC.n523 VCC.n31 72.8958
R1235 VCC.n521 VCC.n31 72.8958
R1236 VCC.n515 VCC.n31 72.8958
R1237 VCC.n513 VCC.n31 72.8958
R1238 VCC.n507 VCC.n31 72.8958
R1239 VCC.n505 VCC.n31 72.8958
R1240 VCC.n499 VCC.n31 72.8958
R1241 VCC.n497 VCC.n31 72.8958
R1242 VCC.n491 VCC.n31 72.8958
R1243 VCC.n489 VCC.n31 72.8958
R1244 VCC.n483 VCC.n31 72.8958
R1245 VCC.n481 VCC.n31 72.8958
R1246 VCC.n475 VCC.n31 72.8958
R1247 VCC.n473 VCC.n31 72.8958
R1248 VCC.n467 VCC.n31 72.8958
R1249 VCC.n465 VCC.n31 72.8958
R1250 VCC.n459 VCC.n31 72.8958
R1251 VCC.n457 VCC.n31 72.8958
R1252 VCC.n451 VCC.n31 72.8958
R1253 VCC.n449 VCC.n31 72.8958
R1254 VCC.n441 VCC.n31 72.8958
R1255 VCC.n161 VCC.n125 72.8958
R1256 VCC.n164 VCC.n125 72.8958
R1257 VCC.n170 VCC.n125 72.8958
R1258 VCC.n172 VCC.n125 72.8958
R1259 VCC.n178 VCC.n125 72.8958
R1260 VCC.n180 VCC.n125 72.8958
R1261 VCC.n186 VCC.n125 72.8958
R1262 VCC.n188 VCC.n125 72.8958
R1263 VCC.n194 VCC.n125 72.8958
R1264 VCC.n196 VCC.n125 72.8958
R1265 VCC.n202 VCC.n125 72.8958
R1266 VCC.n204 VCC.n125 72.8958
R1267 VCC.n210 VCC.n125 72.8958
R1268 VCC.n212 VCC.n125 72.8958
R1269 VCC.n218 VCC.n125 72.8958
R1270 VCC.n220 VCC.n125 72.8958
R1271 VCC.n226 VCC.n125 72.8958
R1272 VCC.n228 VCC.n125 72.8958
R1273 VCC.n234 VCC.n125 72.8958
R1274 VCC.n236 VCC.n125 72.8958
R1275 VCC.n242 VCC.n125 72.8958
R1276 VCC.n244 VCC.n125 72.8958
R1277 VCC.n250 VCC.n125 72.8958
R1278 VCC.n252 VCC.n125 72.8958
R1279 VCC.n258 VCC.n125 72.8958
R1280 VCC.n260 VCC.n125 72.8958
R1281 VCC.n266 VCC.n125 72.8958
R1282 VCC.n268 VCC.n125 72.8958
R1283 VCC.n274 VCC.n125 72.8958
R1284 VCC.n277 VCC.n125 72.8958
R1285 VCC.n444 VCC.n443 56.8247
R1286 VCC.n158 VCC.n157 56.8247
R1287 VCC.n442 VCC.n441 39.2114
R1288 VCC.n450 VCC.n449 39.2114
R1289 VCC.n451 VCC.n439 39.2114
R1290 VCC.n458 VCC.n457 39.2114
R1291 VCC.n459 VCC.n437 39.2114
R1292 VCC.n466 VCC.n465 39.2114
R1293 VCC.n467 VCC.n435 39.2114
R1294 VCC.n474 VCC.n473 39.2114
R1295 VCC.n475 VCC.n433 39.2114
R1296 VCC.n482 VCC.n481 39.2114
R1297 VCC.n483 VCC.n431 39.2114
R1298 VCC.n490 VCC.n489 39.2114
R1299 VCC.n491 VCC.n429 39.2114
R1300 VCC.n498 VCC.n497 39.2114
R1301 VCC.n499 VCC.n427 39.2114
R1302 VCC.n506 VCC.n505 39.2114
R1303 VCC.n507 VCC.n425 39.2114
R1304 VCC.n514 VCC.n513 39.2114
R1305 VCC.n515 VCC.n423 39.2114
R1306 VCC.n522 VCC.n521 39.2114
R1307 VCC.n523 VCC.n421 39.2114
R1308 VCC.n530 VCC.n529 39.2114
R1309 VCC.n531 VCC.n419 39.2114
R1310 VCC.n538 VCC.n537 39.2114
R1311 VCC.n539 VCC.n417 39.2114
R1312 VCC.n546 VCC.n545 39.2114
R1313 VCC.n547 VCC.n415 39.2114
R1314 VCC.n554 VCC.n553 39.2114
R1315 VCC.n555 VCC.n413 39.2114
R1316 VCC.n562 VCC.n561 39.2114
R1317 VCC.n563 VCC.n33 39.2114
R1318 VCC.n161 VCC.n124 39.2114
R1319 VCC.n165 VCC.n164 39.2114
R1320 VCC.n170 VCC.n169 39.2114
R1321 VCC.n173 VCC.n172 39.2114
R1322 VCC.n178 VCC.n177 39.2114
R1323 VCC.n181 VCC.n180 39.2114
R1324 VCC.n186 VCC.n185 39.2114
R1325 VCC.n189 VCC.n188 39.2114
R1326 VCC.n194 VCC.n193 39.2114
R1327 VCC.n197 VCC.n196 39.2114
R1328 VCC.n202 VCC.n201 39.2114
R1329 VCC.n205 VCC.n204 39.2114
R1330 VCC.n210 VCC.n209 39.2114
R1331 VCC.n213 VCC.n212 39.2114
R1332 VCC.n218 VCC.n217 39.2114
R1333 VCC.n221 VCC.n220 39.2114
R1334 VCC.n226 VCC.n225 39.2114
R1335 VCC.n229 VCC.n228 39.2114
R1336 VCC.n234 VCC.n233 39.2114
R1337 VCC.n237 VCC.n236 39.2114
R1338 VCC.n242 VCC.n241 39.2114
R1339 VCC.n245 VCC.n244 39.2114
R1340 VCC.n250 VCC.n249 39.2114
R1341 VCC.n253 VCC.n252 39.2114
R1342 VCC.n258 VCC.n257 39.2114
R1343 VCC.n261 VCC.n260 39.2114
R1344 VCC.n266 VCC.n265 39.2114
R1345 VCC.n269 VCC.n268 39.2114
R1346 VCC.n274 VCC.n273 39.2114
R1347 VCC.n277 VCC.n276 39.2114
R1348 VCC.n564 VCC.n563 39.2114
R1349 VCC.n561 VCC.n560 39.2114
R1350 VCC.n556 VCC.n555 39.2114
R1351 VCC.n553 VCC.n552 39.2114
R1352 VCC.n548 VCC.n547 39.2114
R1353 VCC.n545 VCC.n544 39.2114
R1354 VCC.n540 VCC.n539 39.2114
R1355 VCC.n537 VCC.n536 39.2114
R1356 VCC.n532 VCC.n531 39.2114
R1357 VCC.n529 VCC.n528 39.2114
R1358 VCC.n524 VCC.n523 39.2114
R1359 VCC.n521 VCC.n520 39.2114
R1360 VCC.n516 VCC.n515 39.2114
R1361 VCC.n513 VCC.n512 39.2114
R1362 VCC.n508 VCC.n507 39.2114
R1363 VCC.n505 VCC.n504 39.2114
R1364 VCC.n500 VCC.n499 39.2114
R1365 VCC.n497 VCC.n496 39.2114
R1366 VCC.n492 VCC.n491 39.2114
R1367 VCC.n489 VCC.n488 39.2114
R1368 VCC.n484 VCC.n483 39.2114
R1369 VCC.n481 VCC.n480 39.2114
R1370 VCC.n476 VCC.n475 39.2114
R1371 VCC.n473 VCC.n472 39.2114
R1372 VCC.n468 VCC.n467 39.2114
R1373 VCC.n465 VCC.n464 39.2114
R1374 VCC.n460 VCC.n459 39.2114
R1375 VCC.n457 VCC.n456 39.2114
R1376 VCC.n452 VCC.n451 39.2114
R1377 VCC.n449 VCC.n448 39.2114
R1378 VCC.n441 VCC.n29 39.2114
R1379 VCC.n162 VCC.n161 39.2114
R1380 VCC.n164 VCC.n155 39.2114
R1381 VCC.n171 VCC.n170 39.2114
R1382 VCC.n172 VCC.n153 39.2114
R1383 VCC.n179 VCC.n178 39.2114
R1384 VCC.n180 VCC.n151 39.2114
R1385 VCC.n187 VCC.n186 39.2114
R1386 VCC.n188 VCC.n149 39.2114
R1387 VCC.n195 VCC.n194 39.2114
R1388 VCC.n196 VCC.n147 39.2114
R1389 VCC.n203 VCC.n202 39.2114
R1390 VCC.n204 VCC.n145 39.2114
R1391 VCC.n211 VCC.n210 39.2114
R1392 VCC.n212 VCC.n143 39.2114
R1393 VCC.n219 VCC.n218 39.2114
R1394 VCC.n220 VCC.n141 39.2114
R1395 VCC.n227 VCC.n226 39.2114
R1396 VCC.n228 VCC.n139 39.2114
R1397 VCC.n235 VCC.n234 39.2114
R1398 VCC.n236 VCC.n137 39.2114
R1399 VCC.n243 VCC.n242 39.2114
R1400 VCC.n244 VCC.n135 39.2114
R1401 VCC.n251 VCC.n250 39.2114
R1402 VCC.n252 VCC.n133 39.2114
R1403 VCC.n259 VCC.n258 39.2114
R1404 VCC.n260 VCC.n131 39.2114
R1405 VCC.n267 VCC.n266 39.2114
R1406 VCC.n268 VCC.n129 39.2114
R1407 VCC.n275 VCC.n274 39.2114
R1408 VCC.n278 VCC.n277 39.2114
R1409 VCC.n284 VCC.n125 34.8173
R1410 VCC.n570 VCC.n31 34.8173
R1411 VCC.n446 VCC.n444 29.2853
R1412 VCC.n159 VCC.n158 29.2853
R1413 VCC.n573 VCC.n27 27.5078
R1414 VCC.n567 VCC.n566 27.5078
R1415 VCC.n287 VCC.n123 27.5078
R1416 VCC.n281 VCC.n280 27.5078
R1417 VCC.n284 VCC.n119 20.7248
R1418 VCC.n292 VCC.n119 20.7248
R1419 VCC.n292 VCC.n120 20.7248
R1420 VCC.n300 VCC.n108 20.7248
R1421 VCC.n308 VCC.n108 20.7248
R1422 VCC.n308 VCC.n102 20.7248
R1423 VCC.n316 VCC.n102 20.7248
R1424 VCC.n316 VCC.n95 20.7248
R1425 VCC.n324 VCC.n95 20.7248
R1426 VCC.n324 VCC.n96 20.7248
R1427 VCC.n332 VCC.n84 20.7248
R1428 VCC.n340 VCC.n84 20.7248
R1429 VCC.n340 VCC.n78 20.7248
R1430 VCC.n349 VCC.n78 20.7248
R1431 VCC.n349 VCC.n348 20.7248
R1432 VCC.n357 VCC.n66 20.7248
R1433 VCC.n365 VCC.n66 20.7248
R1434 VCC.n366 VCC.n365 20.7248
R1435 VCC.n367 VCC.n366 20.7248
R1436 VCC.n375 VCC.n60 20.7248
R1437 VCC.n376 VCC.n375 20.7248
R1438 VCC.n377 VCC.n376 20.7248
R1439 VCC.n377 VCC.n53 20.7248
R1440 VCC.n385 VCC.n53 20.7248
R1441 VCC.n387 VCC.n386 20.7248
R1442 VCC.n387 VCC.n46 20.7248
R1443 VCC.n395 VCC.n46 20.7248
R1444 VCC.n396 VCC.n395 20.7248
R1445 VCC.n397 VCC.n396 20.7248
R1446 VCC.n397 VCC.n39 20.7248
R1447 VCC.n405 VCC.n39 20.7248
R1448 VCC.n407 VCC.n406 20.7248
R1449 VCC.n407 VCC.n30 20.7248
R1450 VCC.n570 VCC.n30 20.7248
R1451 VCC.n282 VCC.n117 19.3944
R1452 VCC.n294 VCC.n117 19.3944
R1453 VCC.n294 VCC.n115 19.3944
R1454 VCC.n298 VCC.n115 19.3944
R1455 VCC.n298 VCC.n106 19.3944
R1456 VCC.n310 VCC.n106 19.3944
R1457 VCC.n310 VCC.n104 19.3944
R1458 VCC.n314 VCC.n104 19.3944
R1459 VCC.n314 VCC.n93 19.3944
R1460 VCC.n326 VCC.n93 19.3944
R1461 VCC.n326 VCC.n91 19.3944
R1462 VCC.n330 VCC.n91 19.3944
R1463 VCC.n330 VCC.n82 19.3944
R1464 VCC.n342 VCC.n82 19.3944
R1465 VCC.n342 VCC.n80 19.3944
R1466 VCC.n346 VCC.n80 19.3944
R1467 VCC.n346 VCC.n70 19.3944
R1468 VCC.n359 VCC.n70 19.3944
R1469 VCC.n359 VCC.n68 19.3944
R1470 VCC.n363 VCC.n68 19.3944
R1471 VCC.n363 VCC.n64 19.3944
R1472 VCC.n369 VCC.n64 19.3944
R1473 VCC.n369 VCC.n62 19.3944
R1474 VCC.n373 VCC.n62 19.3944
R1475 VCC.n373 VCC.n57 19.3944
R1476 VCC.n379 VCC.n57 19.3944
R1477 VCC.n379 VCC.n55 19.3944
R1478 VCC.n383 VCC.n55 19.3944
R1479 VCC.n383 VCC.n50 19.3944
R1480 VCC.n389 VCC.n50 19.3944
R1481 VCC.n389 VCC.n48 19.3944
R1482 VCC.n393 VCC.n48 19.3944
R1483 VCC.n393 VCC.n43 19.3944
R1484 VCC.n399 VCC.n43 19.3944
R1485 VCC.n399 VCC.n41 19.3944
R1486 VCC.n403 VCC.n41 19.3944
R1487 VCC.n403 VCC.n36 19.3944
R1488 VCC.n409 VCC.n36 19.3944
R1489 VCC.n409 VCC.n34 19.3944
R1490 VCC.n568 VCC.n34 19.3944
R1491 VCC.n286 VCC.n122 19.3944
R1492 VCC.n290 VCC.n122 19.3944
R1493 VCC.n290 VCC.n112 19.3944
R1494 VCC.n302 VCC.n112 19.3944
R1495 VCC.n302 VCC.n110 19.3944
R1496 VCC.n306 VCC.n110 19.3944
R1497 VCC.n306 VCC.n100 19.3944
R1498 VCC.n318 VCC.n100 19.3944
R1499 VCC.n318 VCC.n98 19.3944
R1500 VCC.n322 VCC.n98 19.3944
R1501 VCC.n322 VCC.n88 19.3944
R1502 VCC.n334 VCC.n88 19.3944
R1503 VCC.n334 VCC.n86 19.3944
R1504 VCC.n338 VCC.n86 19.3944
R1505 VCC.n338 VCC.n76 19.3944
R1506 VCC.n351 VCC.n76 19.3944
R1507 VCC.n351 VCC.n74 19.3944
R1508 VCC.n355 VCC.n74 19.3944
R1509 VCC.n355 VCC.n2 19.3944
R1510 VCC.n602 VCC.n2 19.3944
R1511 VCC.n602 VCC.n601 19.3944
R1512 VCC.n601 VCC.n600 19.3944
R1513 VCC.n600 VCC.n6 19.3944
R1514 VCC.n596 VCC.n6 19.3944
R1515 VCC.n596 VCC.n595 19.3944
R1516 VCC.n595 VCC.n594 19.3944
R1517 VCC.n594 VCC.n11 19.3944
R1518 VCC.n590 VCC.n11 19.3944
R1519 VCC.n590 VCC.n589 19.3944
R1520 VCC.n589 VCC.n588 19.3944
R1521 VCC.n588 VCC.n16 19.3944
R1522 VCC.n584 VCC.n16 19.3944
R1523 VCC.n584 VCC.n583 19.3944
R1524 VCC.n583 VCC.n582 19.3944
R1525 VCC.n582 VCC.n21 19.3944
R1526 VCC.n578 VCC.n21 19.3944
R1527 VCC.n578 VCC.n577 19.3944
R1528 VCC.n577 VCC.n576 19.3944
R1529 VCC.n576 VCC.n26 19.3944
R1530 VCC.n572 VCC.n26 19.3944
R1531 VCC.n357 VCC.t10 19.2741
R1532 VCC.n367 VCC.t8 19.2741
R1533 VCC.n300 VCC.t5 17.2016
R1534 VCC.t1 VCC.n405 17.2016
R1535 VCC.n332 VCC.t11 16.3727
R1536 VCC.t9 VCC.n385 16.3727
R1537 VCC.n445 VCC.n27 10.6151
R1538 VCC.n447 VCC.n440 10.6151
R1539 VCC.n453 VCC.n440 10.6151
R1540 VCC.n454 VCC.n453 10.6151
R1541 VCC.n455 VCC.n454 10.6151
R1542 VCC.n455 VCC.n438 10.6151
R1543 VCC.n461 VCC.n438 10.6151
R1544 VCC.n462 VCC.n461 10.6151
R1545 VCC.n463 VCC.n462 10.6151
R1546 VCC.n463 VCC.n436 10.6151
R1547 VCC.n469 VCC.n436 10.6151
R1548 VCC.n470 VCC.n469 10.6151
R1549 VCC.n471 VCC.n470 10.6151
R1550 VCC.n471 VCC.n434 10.6151
R1551 VCC.n477 VCC.n434 10.6151
R1552 VCC.n478 VCC.n477 10.6151
R1553 VCC.n479 VCC.n478 10.6151
R1554 VCC.n479 VCC.n432 10.6151
R1555 VCC.n485 VCC.n432 10.6151
R1556 VCC.n486 VCC.n485 10.6151
R1557 VCC.n487 VCC.n486 10.6151
R1558 VCC.n487 VCC.n430 10.6151
R1559 VCC.n493 VCC.n430 10.6151
R1560 VCC.n494 VCC.n493 10.6151
R1561 VCC.n495 VCC.n494 10.6151
R1562 VCC.n495 VCC.n428 10.6151
R1563 VCC.n501 VCC.n428 10.6151
R1564 VCC.n502 VCC.n501 10.6151
R1565 VCC.n503 VCC.n502 10.6151
R1566 VCC.n503 VCC.n426 10.6151
R1567 VCC.n509 VCC.n426 10.6151
R1568 VCC.n510 VCC.n509 10.6151
R1569 VCC.n511 VCC.n510 10.6151
R1570 VCC.n511 VCC.n424 10.6151
R1571 VCC.n517 VCC.n424 10.6151
R1572 VCC.n518 VCC.n517 10.6151
R1573 VCC.n519 VCC.n518 10.6151
R1574 VCC.n519 VCC.n422 10.6151
R1575 VCC.n525 VCC.n422 10.6151
R1576 VCC.n526 VCC.n525 10.6151
R1577 VCC.n527 VCC.n526 10.6151
R1578 VCC.n527 VCC.n420 10.6151
R1579 VCC.n533 VCC.n420 10.6151
R1580 VCC.n534 VCC.n533 10.6151
R1581 VCC.n535 VCC.n534 10.6151
R1582 VCC.n535 VCC.n418 10.6151
R1583 VCC.n541 VCC.n418 10.6151
R1584 VCC.n542 VCC.n541 10.6151
R1585 VCC.n543 VCC.n542 10.6151
R1586 VCC.n543 VCC.n416 10.6151
R1587 VCC.n549 VCC.n416 10.6151
R1588 VCC.n550 VCC.n549 10.6151
R1589 VCC.n551 VCC.n550 10.6151
R1590 VCC.n551 VCC.n414 10.6151
R1591 VCC.n557 VCC.n414 10.6151
R1592 VCC.n558 VCC.n557 10.6151
R1593 VCC.n559 VCC.n558 10.6151
R1594 VCC.n559 VCC.n412 10.6151
R1595 VCC.n565 VCC.n412 10.6151
R1596 VCC.n566 VCC.n565 10.6151
R1597 VCC.n160 VCC.n123 10.6151
R1598 VCC.n166 VCC.n156 10.6151
R1599 VCC.n167 VCC.n166 10.6151
R1600 VCC.n168 VCC.n167 10.6151
R1601 VCC.n168 VCC.n154 10.6151
R1602 VCC.n174 VCC.n154 10.6151
R1603 VCC.n175 VCC.n174 10.6151
R1604 VCC.n176 VCC.n175 10.6151
R1605 VCC.n176 VCC.n152 10.6151
R1606 VCC.n182 VCC.n152 10.6151
R1607 VCC.n183 VCC.n182 10.6151
R1608 VCC.n184 VCC.n183 10.6151
R1609 VCC.n184 VCC.n150 10.6151
R1610 VCC.n190 VCC.n150 10.6151
R1611 VCC.n191 VCC.n190 10.6151
R1612 VCC.n192 VCC.n191 10.6151
R1613 VCC.n192 VCC.n148 10.6151
R1614 VCC.n198 VCC.n148 10.6151
R1615 VCC.n199 VCC.n198 10.6151
R1616 VCC.n200 VCC.n199 10.6151
R1617 VCC.n200 VCC.n146 10.6151
R1618 VCC.n206 VCC.n146 10.6151
R1619 VCC.n207 VCC.n206 10.6151
R1620 VCC.n208 VCC.n207 10.6151
R1621 VCC.n208 VCC.n144 10.6151
R1622 VCC.n214 VCC.n144 10.6151
R1623 VCC.n215 VCC.n214 10.6151
R1624 VCC.n216 VCC.n215 10.6151
R1625 VCC.n216 VCC.n142 10.6151
R1626 VCC.n222 VCC.n142 10.6151
R1627 VCC.n223 VCC.n222 10.6151
R1628 VCC.n224 VCC.n223 10.6151
R1629 VCC.n224 VCC.n140 10.6151
R1630 VCC.n230 VCC.n140 10.6151
R1631 VCC.n231 VCC.n230 10.6151
R1632 VCC.n232 VCC.n231 10.6151
R1633 VCC.n232 VCC.n138 10.6151
R1634 VCC.n238 VCC.n138 10.6151
R1635 VCC.n239 VCC.n238 10.6151
R1636 VCC.n240 VCC.n239 10.6151
R1637 VCC.n240 VCC.n136 10.6151
R1638 VCC.n246 VCC.n136 10.6151
R1639 VCC.n247 VCC.n246 10.6151
R1640 VCC.n248 VCC.n247 10.6151
R1641 VCC.n248 VCC.n134 10.6151
R1642 VCC.n254 VCC.n134 10.6151
R1643 VCC.n255 VCC.n254 10.6151
R1644 VCC.n256 VCC.n255 10.6151
R1645 VCC.n256 VCC.n132 10.6151
R1646 VCC.n262 VCC.n132 10.6151
R1647 VCC.n263 VCC.n262 10.6151
R1648 VCC.n264 VCC.n263 10.6151
R1649 VCC.n264 VCC.n130 10.6151
R1650 VCC.n270 VCC.n130 10.6151
R1651 VCC.n271 VCC.n270 10.6151
R1652 VCC.n272 VCC.n271 10.6151
R1653 VCC.n272 VCC.n128 10.6151
R1654 VCC.n128 VCC.n127 10.6151
R1655 VCC.n279 VCC.n127 10.6151
R1656 VCC.n280 VCC.n279 10.6151
R1657 VCC.n601 VCC.n0 9.3005
R1658 VCC.n600 VCC.n599 9.3005
R1659 VCC.n598 VCC.n6 9.3005
R1660 VCC.n597 VCC.n596 9.3005
R1661 VCC.n595 VCC.n7 9.3005
R1662 VCC.n594 VCC.n593 9.3005
R1663 VCC.n592 VCC.n11 9.3005
R1664 VCC.n591 VCC.n590 9.3005
R1665 VCC.n589 VCC.n12 9.3005
R1666 VCC.n588 VCC.n587 9.3005
R1667 VCC.n586 VCC.n16 9.3005
R1668 VCC.n585 VCC.n584 9.3005
R1669 VCC.n583 VCC.n17 9.3005
R1670 VCC.n582 VCC.n581 9.3005
R1671 VCC.n580 VCC.n21 9.3005
R1672 VCC.n579 VCC.n578 9.3005
R1673 VCC.n577 VCC.n22 9.3005
R1674 VCC.n576 VCC.n575 9.3005
R1675 VCC.n574 VCC.n26 9.3005
R1676 VCC.n573 VCC.n572 9.3005
R1677 VCC.n117 VCC.n116 9.3005
R1678 VCC.n295 VCC.n294 9.3005
R1679 VCC.n296 VCC.n115 9.3005
R1680 VCC.n298 VCC.n297 9.3005
R1681 VCC.n106 VCC.n105 9.3005
R1682 VCC.n311 VCC.n310 9.3005
R1683 VCC.n312 VCC.n104 9.3005
R1684 VCC.n314 VCC.n313 9.3005
R1685 VCC.n93 VCC.n92 9.3005
R1686 VCC.n327 VCC.n326 9.3005
R1687 VCC.n328 VCC.n91 9.3005
R1688 VCC.n330 VCC.n329 9.3005
R1689 VCC.n82 VCC.n81 9.3005
R1690 VCC.n343 VCC.n342 9.3005
R1691 VCC.n344 VCC.n80 9.3005
R1692 VCC.n346 VCC.n345 9.3005
R1693 VCC.n70 VCC.n69 9.3005
R1694 VCC.n360 VCC.n359 9.3005
R1695 VCC.n361 VCC.n68 9.3005
R1696 VCC.n363 VCC.n362 9.3005
R1697 VCC.n64 VCC.n63 9.3005
R1698 VCC.n370 VCC.n369 9.3005
R1699 VCC.n371 VCC.n62 9.3005
R1700 VCC.n373 VCC.n372 9.3005
R1701 VCC.n57 VCC.n56 9.3005
R1702 VCC.n380 VCC.n379 9.3005
R1703 VCC.n381 VCC.n55 9.3005
R1704 VCC.n383 VCC.n382 9.3005
R1705 VCC.n50 VCC.n49 9.3005
R1706 VCC.n390 VCC.n389 9.3005
R1707 VCC.n391 VCC.n48 9.3005
R1708 VCC.n393 VCC.n392 9.3005
R1709 VCC.n43 VCC.n42 9.3005
R1710 VCC.n400 VCC.n399 9.3005
R1711 VCC.n401 VCC.n41 9.3005
R1712 VCC.n403 VCC.n402 9.3005
R1713 VCC.n36 VCC.n35 9.3005
R1714 VCC.n410 VCC.n409 9.3005
R1715 VCC.n411 VCC.n34 9.3005
R1716 VCC.n568 VCC.n567 9.3005
R1717 VCC.n282 VCC.n281 9.3005
R1718 VCC.n287 VCC.n286 9.3005
R1719 VCC.n288 VCC.n122 9.3005
R1720 VCC.n290 VCC.n289 9.3005
R1721 VCC.n112 VCC.n111 9.3005
R1722 VCC.n303 VCC.n302 9.3005
R1723 VCC.n304 VCC.n110 9.3005
R1724 VCC.n306 VCC.n305 9.3005
R1725 VCC.n100 VCC.n99 9.3005
R1726 VCC.n319 VCC.n318 9.3005
R1727 VCC.n320 VCC.n98 9.3005
R1728 VCC.n322 VCC.n321 9.3005
R1729 VCC.n88 VCC.n87 9.3005
R1730 VCC.n335 VCC.n334 9.3005
R1731 VCC.n336 VCC.n86 9.3005
R1732 VCC.n338 VCC.n337 9.3005
R1733 VCC.n76 VCC.n75 9.3005
R1734 VCC.n352 VCC.n351 9.3005
R1735 VCC.n353 VCC.n74 9.3005
R1736 VCC.n355 VCC.n354 9.3005
R1737 VCC.n2 VCC.n1 9.3005
R1738 VCC.n603 VCC.n602 9.3005
R1739 VCC.n446 VCC.n445 8.89806
R1740 VCC.n160 VCC.n159 8.89806
R1741 VCC.n96 VCC.t11 4.35259
R1742 VCC.n386 VCC.t9 4.35259
R1743 VCC.n120 VCC.t5 3.52362
R1744 VCC.n406 VCC.t1 3.52362
R1745 VCC.n447 VCC.n446 1.71757
R1746 VCC.n159 VCC.n156 1.71757
R1747 VCC.n348 VCC.t10 1.4512
R1748 VCC.t8 VCC.n60 1.4512
R1749 VCC.n599 VCC.n0 0.152939
R1750 VCC.n599 VCC.n598 0.152939
R1751 VCC.n598 VCC.n597 0.152939
R1752 VCC.n597 VCC.n7 0.152939
R1753 VCC.n593 VCC.n7 0.152939
R1754 VCC.n593 VCC.n592 0.152939
R1755 VCC.n592 VCC.n591 0.152939
R1756 VCC.n591 VCC.n12 0.152939
R1757 VCC.n587 VCC.n12 0.152939
R1758 VCC.n587 VCC.n586 0.152939
R1759 VCC.n586 VCC.n585 0.152939
R1760 VCC.n585 VCC.n17 0.152939
R1761 VCC.n581 VCC.n17 0.152939
R1762 VCC.n581 VCC.n580 0.152939
R1763 VCC.n580 VCC.n579 0.152939
R1764 VCC.n579 VCC.n22 0.152939
R1765 VCC.n575 VCC.n22 0.152939
R1766 VCC.n575 VCC.n574 0.152939
R1767 VCC.n574 VCC.n573 0.152939
R1768 VCC.n281 VCC.n116 0.152939
R1769 VCC.n295 VCC.n116 0.152939
R1770 VCC.n296 VCC.n295 0.152939
R1771 VCC.n297 VCC.n296 0.152939
R1772 VCC.n297 VCC.n105 0.152939
R1773 VCC.n311 VCC.n105 0.152939
R1774 VCC.n312 VCC.n311 0.152939
R1775 VCC.n313 VCC.n312 0.152939
R1776 VCC.n313 VCC.n92 0.152939
R1777 VCC.n327 VCC.n92 0.152939
R1778 VCC.n328 VCC.n327 0.152939
R1779 VCC.n329 VCC.n328 0.152939
R1780 VCC.n329 VCC.n81 0.152939
R1781 VCC.n343 VCC.n81 0.152939
R1782 VCC.n344 VCC.n343 0.152939
R1783 VCC.n345 VCC.n344 0.152939
R1784 VCC.n345 VCC.n69 0.152939
R1785 VCC.n360 VCC.n69 0.152939
R1786 VCC.n361 VCC.n360 0.152939
R1787 VCC.n362 VCC.n361 0.152939
R1788 VCC.n362 VCC.n63 0.152939
R1789 VCC.n370 VCC.n63 0.152939
R1790 VCC.n371 VCC.n370 0.152939
R1791 VCC.n372 VCC.n371 0.152939
R1792 VCC.n372 VCC.n56 0.152939
R1793 VCC.n380 VCC.n56 0.152939
R1794 VCC.n381 VCC.n380 0.152939
R1795 VCC.n382 VCC.n381 0.152939
R1796 VCC.n382 VCC.n49 0.152939
R1797 VCC.n390 VCC.n49 0.152939
R1798 VCC.n391 VCC.n390 0.152939
R1799 VCC.n392 VCC.n391 0.152939
R1800 VCC.n392 VCC.n42 0.152939
R1801 VCC.n400 VCC.n42 0.152939
R1802 VCC.n401 VCC.n400 0.152939
R1803 VCC.n402 VCC.n401 0.152939
R1804 VCC.n402 VCC.n35 0.152939
R1805 VCC.n410 VCC.n35 0.152939
R1806 VCC.n411 VCC.n410 0.152939
R1807 VCC.n567 VCC.n411 0.152939
R1808 VCC.n288 VCC.n287 0.152939
R1809 VCC.n289 VCC.n288 0.152939
R1810 VCC.n289 VCC.n111 0.152939
R1811 VCC.n303 VCC.n111 0.152939
R1812 VCC.n304 VCC.n303 0.152939
R1813 VCC.n305 VCC.n304 0.152939
R1814 VCC.n305 VCC.n99 0.152939
R1815 VCC.n319 VCC.n99 0.152939
R1816 VCC.n320 VCC.n319 0.152939
R1817 VCC.n321 VCC.n320 0.152939
R1818 VCC.n321 VCC.n87 0.152939
R1819 VCC.n335 VCC.n87 0.152939
R1820 VCC.n336 VCC.n335 0.152939
R1821 VCC.n337 VCC.n336 0.152939
R1822 VCC.n337 VCC.n75 0.152939
R1823 VCC.n352 VCC.n75 0.152939
R1824 VCC.n353 VCC.n352 0.152939
R1825 VCC.n354 VCC.n353 0.152939
R1826 VCC.n354 VCC.n1 0.152939
R1827 VCC.n603 VCC.n1 0.13922
R1828 VCC VCC.n0 0.0767195
R1829 VCC VCC.n603 0.063
C0 VGN VGP 0.009895f
C1 VIN VCC 3.33618f
C2 VOUT VGP 6.1027f
C3 VOUT VGN 0.692745f
C4 VIN VGP 6.57638f
C5 VGN VIN 0.807714f
C6 VOUT VIN 5.17404f
C7 VGP VCC 4.24651f
C8 VGN VCC 0.009279f
C9 VOUT VCC 1.52823f
C10 VGN VSS 1.72793f
C11 VOUT VSS 1.534797f
C12 VIN VSS 2.319701f
C13 VGP VSS 1.527386f
C14 VCC VSS 64.64762f
C15 VCC.n0 VSS 0.001515f
C16 VCC.n1 VSS 0.00202f
C17 VCC.n2 VSS 0.001626f
C18 VCC.n3 VSS 0.00202f
C19 VCC.n4 VSS 0.00202f
C20 VCC.n5 VSS 0.00202f
C21 VCC.n6 VSS 0.001626f
C22 VCC.n7 VSS 0.00202f
C23 VCC.n8 VSS 0.00202f
C24 VCC.n9 VSS 0.00202f
C25 VCC.n10 VSS 0.00202f
C26 VCC.n11 VSS 0.001626f
C27 VCC.n12 VSS 0.00202f
C28 VCC.n13 VSS 0.00202f
C29 VCC.n14 VSS 0.00202f
C30 VCC.n15 VSS 0.00202f
C31 VCC.n16 VSS 0.001626f
C32 VCC.n17 VSS 0.00202f
C33 VCC.n18 VSS 0.00202f
C34 VCC.n19 VSS 0.00202f
C35 VCC.n20 VSS 0.00202f
C36 VCC.n21 VSS 0.001626f
C37 VCC.n22 VSS 0.00202f
C38 VCC.n23 VSS 0.00202f
C39 VCC.n24 VSS 0.00202f
C40 VCC.n25 VSS 0.00202f
C41 VCC.n26 VSS 0.001626f
C42 VCC.n27 VSS 0.002563f
C43 VCC.n28 VSS 0.00202f
C44 VCC.n29 VSS 0.003706f
C45 VCC.n30 VSS 0.112929f
C46 VCC.n31 VSS 0.211178f
C47 VCC.n32 VSS 0.00202f
C48 VCC.n33 VSS 0.003706f
C49 VCC.n34 VSS 0.001626f
C50 VCC.n35 VSS 0.00202f
C51 VCC.n36 VSS 0.001626f
C52 VCC.n37 VSS 0.00202f
C53 VCC.n38 VSS 0.00202f
C54 VCC.n39 VSS 0.112929f
C55 VCC.n40 VSS 0.00202f
C56 VCC.n41 VSS 0.001626f
C57 VCC.n42 VSS 0.00202f
C58 VCC.n43 VSS 0.001626f
C59 VCC.n44 VSS 0.00202f
C60 VCC.n45 VSS 0.00202f
C61 VCC.n46 VSS 0.112929f
C62 VCC.n47 VSS 0.00202f
C63 VCC.n48 VSS 0.001626f
C64 VCC.n49 VSS 0.00202f
C65 VCC.n50 VSS 0.001626f
C66 VCC.n51 VSS 0.00202f
C67 VCC.n52 VSS 0.00202f
C68 VCC.n53 VSS 0.112929f
C69 VCC.n54 VSS 0.00202f
C70 VCC.n55 VSS 0.001626f
C71 VCC.n56 VSS 0.00202f
C72 VCC.n57 VSS 0.001626f
C73 VCC.n58 VSS 0.00202f
C74 VCC.n59 VSS 0.00202f
C75 VCC.n60 VSS 0.060417f
C76 VCC.n61 VSS 0.00202f
C77 VCC.n62 VSS 0.001626f
C78 VCC.n63 VSS 0.00202f
C79 VCC.n64 VSS 0.001626f
C80 VCC.n65 VSS 0.00202f
C81 VCC.n66 VSS 0.112929f
C82 VCC.n67 VSS 0.00202f
C83 VCC.n68 VSS 0.001626f
C84 VCC.n69 VSS 0.00202f
C85 VCC.n70 VSS 0.001626f
C86 VCC.n71 VSS 0.00202f
C87 VCC.t10 VSS 0.056465f
C88 VCC.n72 VSS 0.00202f
C89 VCC.n73 VSS 0.00202f
C90 VCC.n74 VSS 0.001626f
C91 VCC.n75 VSS 0.00202f
C92 VCC.n76 VSS 0.001626f
C93 VCC.n77 VSS 0.00202f
C94 VCC.n78 VSS 0.112929f
C95 VCC.n79 VSS 0.00202f
C96 VCC.n80 VSS 0.001626f
C97 VCC.n81 VSS 0.00202f
C98 VCC.n82 VSS 0.001626f
C99 VCC.n83 VSS 0.00202f
C100 VCC.n84 VSS 0.112929f
C101 VCC.n85 VSS 0.00202f
C102 VCC.n86 VSS 0.001626f
C103 VCC.n87 VSS 0.00202f
C104 VCC.n88 VSS 0.001626f
C105 VCC.n89 VSS 0.00202f
C106 VCC.t11 VSS 0.056465f
C107 VCC.n90 VSS 0.00202f
C108 VCC.n91 VSS 0.001626f
C109 VCC.n92 VSS 0.00202f
C110 VCC.n93 VSS 0.001626f
C111 VCC.n94 VSS 0.00202f
C112 VCC.n95 VSS 0.112929f
C113 VCC.n96 VSS 0.068322f
C114 VCC.n97 VSS 0.00202f
C115 VCC.n98 VSS 0.001626f
C116 VCC.n99 VSS 0.00202f
C117 VCC.n100 VSS 0.001626f
C118 VCC.n101 VSS 0.00202f
C119 VCC.n102 VSS 0.112929f
C120 VCC.n103 VSS 0.00202f
C121 VCC.n104 VSS 0.001626f
C122 VCC.n105 VSS 0.00202f
C123 VCC.n106 VSS 0.001626f
C124 VCC.n107 VSS 0.00202f
C125 VCC.n108 VSS 0.112929f
C126 VCC.n109 VSS 0.00202f
C127 VCC.n110 VSS 0.001626f
C128 VCC.n111 VSS 0.00202f
C129 VCC.n112 VSS 0.001626f
C130 VCC.n113 VSS 0.00202f
C131 VCC.t5 VSS 0.056465f
C132 VCC.n114 VSS 0.00202f
C133 VCC.n115 VSS 0.001626f
C134 VCC.n116 VSS 0.00202f
C135 VCC.n117 VSS 0.001626f
C136 VCC.n118 VSS 0.00202f
C137 VCC.n119 VSS 0.112929f
C138 VCC.n120 VSS 0.066064f
C139 VCC.n121 VSS 0.00202f
C140 VCC.n122 VSS 0.001626f
C141 VCC.n123 VSS 0.002563f
C142 VCC.n124 VSS 0.003706f
C143 VCC.n125 VSS 0.211178f
C144 VCC.n126 VSS 0.003706f
C145 VCC.n127 VSS 0.001374f
C146 VCC.n128 VSS 0.001374f
C147 VCC.n129 VSS 0.001374f
C148 VCC.n130 VSS 0.001374f
C149 VCC.n131 VSS 0.001374f
C150 VCC.n132 VSS 0.001374f
C151 VCC.n133 VSS 0.001374f
C152 VCC.n134 VSS 0.001374f
C153 VCC.n135 VSS 0.001374f
C154 VCC.n136 VSS 0.001374f
C155 VCC.n137 VSS 0.001374f
C156 VCC.n138 VSS 0.001374f
C157 VCC.n139 VSS 0.001374f
C158 VCC.n140 VSS 0.001374f
C159 VCC.n141 VSS 0.001374f
C160 VCC.n142 VSS 0.001374f
C161 VCC.n143 VSS 0.001374f
C162 VCC.n144 VSS 0.001374f
C163 VCC.n145 VSS 0.001374f
C164 VCC.n146 VSS 0.001374f
C165 VCC.n147 VSS 0.001374f
C166 VCC.n148 VSS 0.001374f
C167 VCC.n149 VSS 0.001374f
C168 VCC.n150 VSS 0.001374f
C169 VCC.n151 VSS 0.001374f
C170 VCC.n152 VSS 0.001374f
C171 VCC.n153 VSS 0.001374f
C172 VCC.n154 VSS 0.001374f
C173 VCC.n155 VSS 0.001374f
C174 VCC.n156 VSS 7.98e-19
C175 VCC.t6 VSS 0.072685f
C176 VCC.t7 VSS 0.079284f
C177 VCC.t4 VSS 0.424228f
C178 VCC.n157 VSS 0.121117f
C179 VCC.n158 VSS 0.065124f
C180 VCC.n159 VSS 0.001914f
C181 VCC.n160 VSS 0.001263f
C182 VCC.n162 VSS 0.001374f
C183 VCC.n163 VSS 0.001374f
C184 VCC.n165 VSS 0.001374f
C185 VCC.n166 VSS 0.001374f
C186 VCC.n167 VSS 0.001374f
C187 VCC.n168 VSS 0.001374f
C188 VCC.n169 VSS 0.001374f
C189 VCC.n171 VSS 0.001374f
C190 VCC.n173 VSS 0.001374f
C191 VCC.n174 VSS 0.001374f
C192 VCC.n175 VSS 0.001374f
C193 VCC.n176 VSS 0.001374f
C194 VCC.n177 VSS 0.001374f
C195 VCC.n179 VSS 0.001374f
C196 VCC.n181 VSS 0.001374f
C197 VCC.n182 VSS 0.001374f
C198 VCC.n183 VSS 0.001374f
C199 VCC.n184 VSS 0.001374f
C200 VCC.n185 VSS 0.001374f
C201 VCC.n187 VSS 0.001374f
C202 VCC.n189 VSS 0.001374f
C203 VCC.n190 VSS 0.001374f
C204 VCC.n191 VSS 0.001374f
C205 VCC.n192 VSS 0.001374f
C206 VCC.n193 VSS 0.001374f
C207 VCC.n195 VSS 0.001374f
C208 VCC.n197 VSS 0.001374f
C209 VCC.n198 VSS 0.001374f
C210 VCC.n199 VSS 0.001374f
C211 VCC.n200 VSS 0.001374f
C212 VCC.n201 VSS 0.001374f
C213 VCC.n203 VSS 0.001374f
C214 VCC.n205 VSS 0.001374f
C215 VCC.n206 VSS 0.001374f
C216 VCC.n207 VSS 0.001374f
C217 VCC.n208 VSS 0.001374f
C218 VCC.n209 VSS 0.001374f
C219 VCC.n211 VSS 0.001374f
C220 VCC.n213 VSS 0.001374f
C221 VCC.n214 VSS 0.001374f
C222 VCC.n215 VSS 0.001374f
C223 VCC.n216 VSS 0.001374f
C224 VCC.n217 VSS 0.001374f
C225 VCC.n219 VSS 0.001374f
C226 VCC.n221 VSS 0.001374f
C227 VCC.n222 VSS 0.001374f
C228 VCC.n223 VSS 0.001374f
C229 VCC.n224 VSS 0.001374f
C230 VCC.n225 VSS 0.001374f
C231 VCC.n227 VSS 0.001374f
C232 VCC.n229 VSS 0.001374f
C233 VCC.n230 VSS 0.001374f
C234 VCC.n231 VSS 0.001374f
C235 VCC.n232 VSS 0.001374f
C236 VCC.n233 VSS 0.001374f
C237 VCC.n235 VSS 0.001374f
C238 VCC.n237 VSS 0.001374f
C239 VCC.n238 VSS 0.001374f
C240 VCC.n239 VSS 0.001374f
C241 VCC.n240 VSS 0.001374f
C242 VCC.n241 VSS 0.001374f
C243 VCC.n243 VSS 0.001374f
C244 VCC.n245 VSS 0.001374f
C245 VCC.n246 VSS 0.001374f
C246 VCC.n247 VSS 0.001374f
C247 VCC.n248 VSS 0.001374f
C248 VCC.n249 VSS 0.001374f
C249 VCC.n251 VSS 0.001374f
C250 VCC.n253 VSS 0.001374f
C251 VCC.n254 VSS 0.001374f
C252 VCC.n255 VSS 0.001374f
C253 VCC.n256 VSS 0.001374f
C254 VCC.n257 VSS 0.001374f
C255 VCC.n259 VSS 0.001374f
C256 VCC.n261 VSS 0.001374f
C257 VCC.n262 VSS 0.001374f
C258 VCC.n263 VSS 0.001374f
C259 VCC.n264 VSS 0.001374f
C260 VCC.n265 VSS 0.001374f
C261 VCC.n267 VSS 0.001374f
C262 VCC.n269 VSS 0.001374f
C263 VCC.n270 VSS 0.001374f
C264 VCC.n271 VSS 0.001374f
C265 VCC.n272 VSS 0.001374f
C266 VCC.n273 VSS 0.001374f
C267 VCC.n275 VSS 0.001374f
C268 VCC.n276 VSS 0.001374f
C269 VCC.n278 VSS 0.001374f
C270 VCC.n279 VSS 0.001374f
C271 VCC.n280 VSS 0.002563f
C272 VCC.n281 VSS 0.006507f
C273 VCC.n282 VSS 0.00135f
C274 VCC.n283 VSS 0.003708f
C275 VCC.n284 VSS 0.151325f
C276 VCC.n285 VSS 0.003708f
C277 VCC.n286 VSS 0.00135f
C278 VCC.n287 VSS 0.006507f
C279 VCC.n288 VSS 0.00202f
C280 VCC.n289 VSS 0.00202f
C281 VCC.n290 VSS 0.001626f
C282 VCC.n291 VSS 0.00202f
C283 VCC.n292 VSS 0.112929f
C284 VCC.n293 VSS 0.00202f
C285 VCC.n294 VSS 0.001626f
C286 VCC.n295 VSS 0.00202f
C287 VCC.n296 VSS 0.00202f
C288 VCC.n297 VSS 0.00202f
C289 VCC.n298 VSS 0.001626f
C290 VCC.n299 VSS 0.00202f
C291 VCC.n300 VSS 0.10333f
C292 VCC.n301 VSS 0.00202f
C293 VCC.n302 VSS 0.001626f
C294 VCC.n303 VSS 0.00202f
C295 VCC.n304 VSS 0.00202f
C296 VCC.n305 VSS 0.00202f
C297 VCC.n306 VSS 0.001626f
C298 VCC.n307 VSS 0.00202f
C299 VCC.n308 VSS 0.112929f
C300 VCC.n309 VSS 0.00202f
C301 VCC.n310 VSS 0.001626f
C302 VCC.n311 VSS 0.00202f
C303 VCC.n312 VSS 0.00202f
C304 VCC.n313 VSS 0.00202f
C305 VCC.n314 VSS 0.001626f
C306 VCC.n315 VSS 0.00202f
C307 VCC.n316 VSS 0.112929f
C308 VCC.n317 VSS 0.00202f
C309 VCC.n318 VSS 0.001626f
C310 VCC.n319 VSS 0.00202f
C311 VCC.n320 VSS 0.00202f
C312 VCC.n321 VSS 0.00202f
C313 VCC.n322 VSS 0.001626f
C314 VCC.n323 VSS 0.00202f
C315 VCC.n324 VSS 0.112929f
C316 VCC.n325 VSS 0.00202f
C317 VCC.n326 VSS 0.001626f
C318 VCC.n327 VSS 0.00202f
C319 VCC.n328 VSS 0.00202f
C320 VCC.n329 VSS 0.00202f
C321 VCC.n330 VSS 0.001626f
C322 VCC.n331 VSS 0.00202f
C323 VCC.n332 VSS 0.101072f
C324 VCC.n333 VSS 0.00202f
C325 VCC.n334 VSS 0.001626f
C326 VCC.n335 VSS 0.00202f
C327 VCC.n336 VSS 0.00202f
C328 VCC.n337 VSS 0.00202f
C329 VCC.n338 VSS 0.001626f
C330 VCC.n339 VSS 0.00202f
C331 VCC.n340 VSS 0.112929f
C332 VCC.n341 VSS 0.00202f
C333 VCC.n342 VSS 0.001626f
C334 VCC.n343 VSS 0.00202f
C335 VCC.n344 VSS 0.00202f
C336 VCC.n345 VSS 0.00202f
C337 VCC.n346 VSS 0.001626f
C338 VCC.n347 VSS 0.00202f
C339 VCC.n348 VSS 0.060417f
C340 VCC.n349 VSS 0.112929f
C341 VCC.n350 VSS 0.00202f
C342 VCC.n351 VSS 0.001626f
C343 VCC.n352 VSS 0.00202f
C344 VCC.n353 VSS 0.00202f
C345 VCC.n354 VSS 0.00202f
C346 VCC.n355 VSS 0.001626f
C347 VCC.n356 VSS 0.00202f
C348 VCC.n357 VSS 0.108977f
C349 VCC.n358 VSS 0.00202f
C350 VCC.n359 VSS 0.001626f
C351 VCC.n360 VSS 0.00202f
C352 VCC.n361 VSS 0.00202f
C353 VCC.n362 VSS 0.00202f
C354 VCC.n363 VSS 0.001626f
C355 VCC.n364 VSS 0.00202f
C356 VCC.n365 VSS 0.112929f
C357 VCC.n366 VSS 0.112929f
C358 VCC.t8 VSS 0.056465f
C359 VCC.n367 VSS 0.108977f
C360 VCC.n368 VSS 0.00202f
C361 VCC.n369 VSS 0.001626f
C362 VCC.n370 VSS 0.00202f
C363 VCC.n371 VSS 0.00202f
C364 VCC.n372 VSS 0.00202f
C365 VCC.n373 VSS 0.001626f
C366 VCC.n374 VSS 0.00202f
C367 VCC.n375 VSS 0.112929f
C368 VCC.n376 VSS 0.112929f
C369 VCC.n377 VSS 0.112929f
C370 VCC.n378 VSS 0.00202f
C371 VCC.n379 VSS 0.001626f
C372 VCC.n380 VSS 0.00202f
C373 VCC.n381 VSS 0.00202f
C374 VCC.n382 VSS 0.00202f
C375 VCC.n383 VSS 0.001626f
C376 VCC.n384 VSS 0.00202f
C377 VCC.n385 VSS 0.101072f
C378 VCC.t9 VSS 0.056465f
C379 VCC.n386 VSS 0.068322f
C380 VCC.n387 VSS 0.112929f
C381 VCC.n388 VSS 0.00202f
C382 VCC.n389 VSS 0.001626f
C383 VCC.n390 VSS 0.00202f
C384 VCC.n391 VSS 0.00202f
C385 VCC.n392 VSS 0.00202f
C386 VCC.n393 VSS 0.001626f
C387 VCC.n394 VSS 0.00202f
C388 VCC.n395 VSS 0.112929f
C389 VCC.n396 VSS 0.112929f
C390 VCC.n397 VSS 0.112929f
C391 VCC.n398 VSS 0.00202f
C392 VCC.n399 VSS 0.001626f
C393 VCC.n400 VSS 0.00202f
C394 VCC.n401 VSS 0.00202f
C395 VCC.n402 VSS 0.00202f
C396 VCC.n403 VSS 0.001626f
C397 VCC.n404 VSS 0.00202f
C398 VCC.n405 VSS 0.10333f
C399 VCC.t1 VSS 0.056465f
C400 VCC.n406 VSS 0.066064f
C401 VCC.n407 VSS 0.112929f
C402 VCC.n408 VSS 0.00202f
C403 VCC.n409 VSS 0.001626f
C404 VCC.n410 VSS 0.00202f
C405 VCC.n411 VSS 0.00202f
C406 VCC.n412 VSS 0.001374f
C407 VCC.n413 VSS 0.001374f
C408 VCC.n414 VSS 0.001374f
C409 VCC.n415 VSS 0.001374f
C410 VCC.n416 VSS 0.001374f
C411 VCC.n417 VSS 0.001374f
C412 VCC.n418 VSS 0.001374f
C413 VCC.n419 VSS 0.001374f
C414 VCC.n420 VSS 0.001374f
C415 VCC.n421 VSS 0.001374f
C416 VCC.n422 VSS 0.001374f
C417 VCC.n423 VSS 0.001374f
C418 VCC.n424 VSS 0.001374f
C419 VCC.n425 VSS 0.001374f
C420 VCC.n426 VSS 0.001374f
C421 VCC.n427 VSS 0.001374f
C422 VCC.n428 VSS 0.001374f
C423 VCC.n429 VSS 0.001374f
C424 VCC.n430 VSS 0.001374f
C425 VCC.n431 VSS 0.001374f
C426 VCC.n432 VSS 0.001374f
C427 VCC.n433 VSS 0.001374f
C428 VCC.n434 VSS 0.001374f
C429 VCC.n435 VSS 0.001374f
C430 VCC.n436 VSS 0.001374f
C431 VCC.n437 VSS 0.001374f
C432 VCC.n438 VSS 0.001374f
C433 VCC.n439 VSS 0.001374f
C434 VCC.n440 VSS 0.001374f
C435 VCC.n442 VSS 0.001374f
C436 VCC.t3 VSS 0.072685f
C437 VCC.t2 VSS 0.079284f
C438 VCC.t0 VSS 0.424228f
C439 VCC.n443 VSS 0.121117f
C440 VCC.n444 VSS 0.065124f
C441 VCC.n445 VSS 0.001263f
C442 VCC.n446 VSS 0.001914f
C443 VCC.n447 VSS 7.98e-19
C444 VCC.n448 VSS 0.001374f
C445 VCC.n450 VSS 0.001374f
C446 VCC.n452 VSS 0.001374f
C447 VCC.n453 VSS 0.001374f
C448 VCC.n454 VSS 0.001374f
C449 VCC.n455 VSS 0.001374f
C450 VCC.n456 VSS 0.001374f
C451 VCC.n458 VSS 0.001374f
C452 VCC.n460 VSS 0.001374f
C453 VCC.n461 VSS 0.001374f
C454 VCC.n462 VSS 0.001374f
C455 VCC.n463 VSS 0.001374f
C456 VCC.n464 VSS 0.001374f
C457 VCC.n466 VSS 0.001374f
C458 VCC.n468 VSS 0.001374f
C459 VCC.n469 VSS 0.001374f
C460 VCC.n470 VSS 0.001374f
C461 VCC.n471 VSS 0.001374f
C462 VCC.n472 VSS 0.001374f
C463 VCC.n474 VSS 0.001374f
C464 VCC.n476 VSS 0.001374f
C465 VCC.n477 VSS 0.001374f
C466 VCC.n478 VSS 0.001374f
C467 VCC.n479 VSS 0.001374f
C468 VCC.n480 VSS 0.001374f
C469 VCC.n482 VSS 0.001374f
C470 VCC.n484 VSS 0.001374f
C471 VCC.n485 VSS 0.001374f
C472 VCC.n486 VSS 0.001374f
C473 VCC.n487 VSS 0.001374f
C474 VCC.n488 VSS 0.001374f
C475 VCC.n490 VSS 0.001374f
C476 VCC.n492 VSS 0.001374f
C477 VCC.n493 VSS 0.001374f
C478 VCC.n494 VSS 0.001374f
C479 VCC.n495 VSS 0.001374f
C480 VCC.n496 VSS 0.001374f
C481 VCC.n498 VSS 0.001374f
C482 VCC.n500 VSS 0.001374f
C483 VCC.n501 VSS 0.001374f
C484 VCC.n502 VSS 0.001374f
C485 VCC.n503 VSS 0.001374f
C486 VCC.n504 VSS 0.001374f
C487 VCC.n506 VSS 0.001374f
C488 VCC.n508 VSS 0.001374f
C489 VCC.n509 VSS 0.001374f
C490 VCC.n510 VSS 0.001374f
C491 VCC.n511 VSS 0.001374f
C492 VCC.n512 VSS 0.001374f
C493 VCC.n514 VSS 0.001374f
C494 VCC.n516 VSS 0.001374f
C495 VCC.n517 VSS 0.001374f
C496 VCC.n518 VSS 0.001374f
C497 VCC.n519 VSS 0.001374f
C498 VCC.n520 VSS 0.001374f
C499 VCC.n522 VSS 0.001374f
C500 VCC.n524 VSS 0.001374f
C501 VCC.n525 VSS 0.001374f
C502 VCC.n526 VSS 0.001374f
C503 VCC.n527 VSS 0.001374f
C504 VCC.n528 VSS 0.001374f
C505 VCC.n530 VSS 0.001374f
C506 VCC.n532 VSS 0.001374f
C507 VCC.n533 VSS 0.001374f
C508 VCC.n534 VSS 0.001374f
C509 VCC.n535 VSS 0.001374f
C510 VCC.n536 VSS 0.001374f
C511 VCC.n538 VSS 0.001374f
C512 VCC.n540 VSS 0.001374f
C513 VCC.n541 VSS 0.001374f
C514 VCC.n542 VSS 0.001374f
C515 VCC.n543 VSS 0.001374f
C516 VCC.n544 VSS 0.001374f
C517 VCC.n546 VSS 0.001374f
C518 VCC.n548 VSS 0.001374f
C519 VCC.n549 VSS 0.001374f
C520 VCC.n550 VSS 0.001374f
C521 VCC.n551 VSS 0.001374f
C522 VCC.n552 VSS 0.001374f
C523 VCC.n554 VSS 0.001374f
C524 VCC.n556 VSS 0.001374f
C525 VCC.n557 VSS 0.001374f
C526 VCC.n558 VSS 0.001374f
C527 VCC.n559 VSS 0.001374f
C528 VCC.n560 VSS 0.001374f
C529 VCC.n562 VSS 0.001374f
C530 VCC.n564 VSS 0.001374f
C531 VCC.n565 VSS 0.001374f
C532 VCC.n566 VSS 0.002563f
C533 VCC.n567 VSS 0.006507f
C534 VCC.n568 VSS 0.00135f
C535 VCC.n569 VSS 0.003708f
C536 VCC.n570 VSS 0.151325f
C537 VCC.n571 VSS 0.003708f
C538 VCC.n572 VSS 0.00135f
C539 VCC.n573 VSS 0.006507f
C540 VCC.n574 VSS 0.00202f
C541 VCC.n575 VSS 0.00202f
C542 VCC.n576 VSS 0.001626f
C543 VCC.n577 VSS 0.001626f
C544 VCC.n578 VSS 0.001626f
C545 VCC.n579 VSS 0.00202f
C546 VCC.n580 VSS 0.00202f
C547 VCC.n581 VSS 0.00202f
C548 VCC.n582 VSS 0.001626f
C549 VCC.n583 VSS 0.001626f
C550 VCC.n584 VSS 0.001626f
C551 VCC.n585 VSS 0.00202f
C552 VCC.n586 VSS 0.00202f
C553 VCC.n587 VSS 0.00202f
C554 VCC.n588 VSS 0.001626f
C555 VCC.n589 VSS 0.001626f
C556 VCC.n590 VSS 0.001626f
C557 VCC.n591 VSS 0.00202f
C558 VCC.n592 VSS 0.00202f
C559 VCC.n593 VSS 0.00202f
C560 VCC.n594 VSS 0.001626f
C561 VCC.n595 VSS 0.001626f
C562 VCC.n596 VSS 0.001626f
C563 VCC.n597 VSS 0.00202f
C564 VCC.n598 VSS 0.00202f
C565 VCC.n599 VSS 0.00202f
C566 VCC.n600 VSS 0.001626f
C567 VCC.n601 VSS 0.001626f
C568 VCC.n602 VSS 0.001626f
C569 VCC.n603 VSS 0.001848f
C570 VGP.n0 VSS 0.028443f
C571 VGP.t0 VSS 2.90307f
C572 VGP.n1 VSS 0.035541f
C573 VGP.n2 VSS 0.021575f
C574 VGP.t1 VSS 2.90307f
C575 VGP.n3 VSS 1.00491f
C576 VGP.n4 VSS 0.021575f
C577 VGP.n5 VSS 0.031363f
C578 VGP.n6 VSS 0.208408f
C579 VGP.t3 VSS 2.90307f
C580 VGP.t2 VSS 3.08323f
C581 VGP.n7 VSS 1.04524f
C582 VGP.n8 VSS 1.06532f
C583 VGP.n9 VSS 0.028751f
C584 VGP.n10 VSS 0.040009f
C585 VGP.n11 VSS 0.021575f
C586 VGP.n12 VSS 0.021575f
C587 VGP.n13 VSS 0.021575f
C588 VGP.n14 VSS 0.031363f
C589 VGP.n15 VSS 0.040009f
C590 VGP.n16 VSS 0.028751f
C591 VGP.n17 VSS 0.021575f
C592 VGP.n18 VSS 0.021575f
C593 VGP.n19 VSS 0.031516f
C594 VGP.n20 VSS 0.040009f
C595 VGP.n21 VSS 0.027184f
C596 VGP.n22 VSS 0.021575f
C597 VGP.n23 VSS 0.021575f
C598 VGP.n24 VSS 0.021575f
C599 VGP.n25 VSS 0.040009f
C600 VGP.n26 VSS 0.025986f
C601 VGP.n27 VSS 1.07342f
C602 VGP.n28 VSS 0.042691f
C603 VIN.n0 VSS 0.011894f
C604 VIN.n1 VSS 0.026794f
C605 VIN.n2 VSS 0.012003f
C606 VIN.n3 VSS 0.021096f
C607 VIN.n4 VSS 0.011336f
C608 VIN.n5 VSS 0.026794f
C609 VIN.n6 VSS 0.012003f
C610 VIN.n7 VSS 0.021096f
C611 VIN.n8 VSS 0.011336f
C612 VIN.n9 VSS 0.026794f
C613 VIN.n10 VSS 0.012003f
C614 VIN.n11 VSS 0.021096f
C615 VIN.n12 VSS 0.011336f
C616 VIN.n13 VSS 0.026794f
C617 VIN.n14 VSS 0.012003f
C618 VIN.n15 VSS 0.021096f
C619 VIN.n16 VSS 0.011336f
C620 VIN.n17 VSS 0.026794f
C621 VIN.n18 VSS 0.012003f
C622 VIN.n19 VSS 0.021096f
C623 VIN.n20 VSS 0.011336f
C624 VIN.n21 VSS 0.026794f
C625 VIN.n22 VSS 0.011669f
C626 VIN.n23 VSS 0.021096f
C627 VIN.n24 VSS 0.012003f
C628 VIN.n25 VSS 0.026794f
C629 VIN.n26 VSS 0.012003f
C630 VIN.n27 VSS 0.021096f
C631 VIN.n28 VSS 0.011336f
C632 VIN.n29 VSS 0.026794f
C633 VIN.n30 VSS 0.012003f
C634 VIN.n31 VSS 1.66506f
C635 VIN.n32 VSS 0.011336f
C636 VIN.t2 VSS 0.058223f
C637 VIN.n33 VSS 0.231004f
C638 VIN.n34 VSS 0.020156f
C639 VIN.n35 VSS 0.020096f
C640 VIN.n36 VSS 0.026794f
C641 VIN.n37 VSS 0.012003f
C642 VIN.n38 VSS 0.011336f
C643 VIN.n39 VSS 0.021096f
C644 VIN.n40 VSS 0.021096f
C645 VIN.n41 VSS 0.011336f
C646 VIN.n42 VSS 0.012003f
C647 VIN.n43 VSS 0.026794f
C648 VIN.n44 VSS 0.026794f
C649 VIN.n45 VSS 0.012003f
C650 VIN.n46 VSS 0.011336f
C651 VIN.n47 VSS 0.021096f
C652 VIN.n48 VSS 0.021096f
C653 VIN.n49 VSS 0.011336f
C654 VIN.n50 VSS 0.011336f
C655 VIN.n51 VSS 0.012003f
C656 VIN.n52 VSS 0.026794f
C657 VIN.n53 VSS 0.026794f
C658 VIN.n54 VSS 0.026794f
C659 VIN.n55 VSS 0.011669f
C660 VIN.n56 VSS 0.011336f
C661 VIN.n57 VSS 0.021096f
C662 VIN.n58 VSS 0.021096f
C663 VIN.n59 VSS 0.011336f
C664 VIN.n60 VSS 0.012003f
C665 VIN.n61 VSS 0.026794f
C666 VIN.n62 VSS 0.026794f
C667 VIN.n63 VSS 0.012003f
C668 VIN.n64 VSS 0.011336f
C669 VIN.n65 VSS 0.021096f
C670 VIN.n66 VSS 0.021096f
C671 VIN.n67 VSS 0.011336f
C672 VIN.n68 VSS 0.012003f
C673 VIN.n69 VSS 0.026794f
C674 VIN.n70 VSS 0.026794f
C675 VIN.n71 VSS 0.012003f
C676 VIN.n72 VSS 0.011336f
C677 VIN.n73 VSS 0.021096f
C678 VIN.n74 VSS 0.021096f
C679 VIN.n75 VSS 0.011336f
C680 VIN.n76 VSS 0.012003f
C681 VIN.n77 VSS 0.026794f
C682 VIN.n78 VSS 0.026794f
C683 VIN.n79 VSS 0.012003f
C684 VIN.n80 VSS 0.011336f
C685 VIN.n81 VSS 0.021096f
C686 VIN.n82 VSS 0.021096f
C687 VIN.n83 VSS 0.011336f
C688 VIN.n84 VSS 0.012003f
C689 VIN.n85 VSS 0.026794f
C690 VIN.n86 VSS 0.026794f
C691 VIN.n87 VSS 0.012003f
C692 VIN.n88 VSS 0.011336f
C693 VIN.n89 VSS 0.021096f
C694 VIN.n90 VSS 0.021096f
C695 VIN.n91 VSS 0.011336f
C696 VIN.n92 VSS 0.012003f
C697 VIN.n93 VSS 0.026794f
C698 VIN.n94 VSS 0.026794f
C699 VIN.n95 VSS 0.012003f
C700 VIN.n96 VSS 0.011336f
C701 VIN.n97 VSS 0.021096f
C702 VIN.n98 VSS 0.054526f
C703 VIN.n99 VSS 0.011336f
C704 VIN.n100 VSS 0.012003f
C705 VIN.n101 VSS 0.06091f
C706 VIN.n102 VSS 0.053708f
C707 VIN.t7 VSS 0.313406f
C708 VIN.t0 VSS 0.313406f
C709 VIN.n103 VSS 2.51904f
C710 VIN.n104 VSS 1.01931f
C711 VIN.n105 VSS 0.011894f
C712 VIN.n106 VSS 0.026794f
C713 VIN.n107 VSS 0.012003f
C714 VIN.n108 VSS 0.021096f
C715 VIN.n109 VSS 0.011336f
C716 VIN.n110 VSS 0.026794f
C717 VIN.n111 VSS 0.012003f
C718 VIN.n112 VSS 0.021096f
C719 VIN.n113 VSS 0.011336f
C720 VIN.n114 VSS 0.026794f
C721 VIN.n115 VSS 0.012003f
C722 VIN.n116 VSS 0.021096f
C723 VIN.n117 VSS 0.011336f
C724 VIN.n118 VSS 0.026794f
C725 VIN.n119 VSS 0.012003f
C726 VIN.n120 VSS 0.021096f
C727 VIN.n121 VSS 0.011336f
C728 VIN.n122 VSS 0.026794f
C729 VIN.n123 VSS 0.012003f
C730 VIN.n124 VSS 0.021096f
C731 VIN.n125 VSS 0.011336f
C732 VIN.n126 VSS 0.026794f
C733 VIN.n127 VSS 0.011669f
C734 VIN.n128 VSS 0.021096f
C735 VIN.n129 VSS 0.012003f
C736 VIN.n130 VSS 0.026794f
C737 VIN.n131 VSS 0.012003f
C738 VIN.n132 VSS 0.021096f
C739 VIN.n133 VSS 0.011336f
C740 VIN.n134 VSS 0.026794f
C741 VIN.n135 VSS 0.012003f
C742 VIN.n136 VSS 1.66506f
C743 VIN.n137 VSS 0.011336f
C744 VIN.t1 VSS 0.058223f
C745 VIN.n138 VSS 0.231004f
C746 VIN.n139 VSS 0.020156f
C747 VIN.n140 VSS 0.020096f
C748 VIN.n141 VSS 0.026794f
C749 VIN.n142 VSS 0.012003f
C750 VIN.n143 VSS 0.011336f
C751 VIN.n144 VSS 0.021096f
C752 VIN.n145 VSS 0.021096f
C753 VIN.n146 VSS 0.011336f
C754 VIN.n147 VSS 0.012003f
C755 VIN.n148 VSS 0.026794f
C756 VIN.n149 VSS 0.026794f
C757 VIN.n150 VSS 0.012003f
C758 VIN.n151 VSS 0.011336f
C759 VIN.n152 VSS 0.021096f
C760 VIN.n153 VSS 0.021096f
C761 VIN.n154 VSS 0.011336f
C762 VIN.n155 VSS 0.011336f
C763 VIN.n156 VSS 0.012003f
C764 VIN.n157 VSS 0.026794f
C765 VIN.n158 VSS 0.026794f
C766 VIN.n159 VSS 0.026794f
C767 VIN.n160 VSS 0.011669f
C768 VIN.n161 VSS 0.011336f
C769 VIN.n162 VSS 0.021096f
C770 VIN.n163 VSS 0.021096f
C771 VIN.n164 VSS 0.011336f
C772 VIN.n165 VSS 0.012003f
C773 VIN.n166 VSS 0.026794f
C774 VIN.n167 VSS 0.026794f
C775 VIN.n168 VSS 0.012003f
C776 VIN.n169 VSS 0.011336f
C777 VIN.n170 VSS 0.021096f
C778 VIN.n171 VSS 0.021096f
C779 VIN.n172 VSS 0.011336f
C780 VIN.n173 VSS 0.012003f
C781 VIN.n174 VSS 0.026794f
C782 VIN.n175 VSS 0.026794f
C783 VIN.n176 VSS 0.012003f
C784 VIN.n177 VSS 0.011336f
C785 VIN.n178 VSS 0.021096f
C786 VIN.n179 VSS 0.021096f
C787 VIN.n180 VSS 0.011336f
C788 VIN.n181 VSS 0.012003f
C789 VIN.n182 VSS 0.026794f
C790 VIN.n183 VSS 0.026794f
C791 VIN.n184 VSS 0.012003f
C792 VIN.n185 VSS 0.011336f
C793 VIN.n186 VSS 0.021096f
C794 VIN.n187 VSS 0.021096f
C795 VIN.n188 VSS 0.011336f
C796 VIN.n189 VSS 0.012003f
C797 VIN.n190 VSS 0.026794f
C798 VIN.n191 VSS 0.026794f
C799 VIN.n192 VSS 0.012003f
C800 VIN.n193 VSS 0.011336f
C801 VIN.n194 VSS 0.021096f
C802 VIN.n195 VSS 0.021096f
C803 VIN.n196 VSS 0.011336f
C804 VIN.n197 VSS 0.012003f
C805 VIN.n198 VSS 0.026794f
C806 VIN.n199 VSS 0.026794f
C807 VIN.n200 VSS 0.012003f
C808 VIN.n201 VSS 0.011336f
C809 VIN.n202 VSS 0.021096f
C810 VIN.n203 VSS 0.054526f
C811 VIN.n204 VSS 0.011336f
C812 VIN.n205 VSS 0.012003f
C813 VIN.n206 VSS 0.06091f
C814 VIN.n207 VSS 0.040409f
C815 VIN.n208 VSS 0.455423f
C816 VIN.t5 VSS 0.511743f
C817 VIN.t3 VSS 0.057513f
C818 VIN.t4 VSS 0.057513f
C819 VIN.n209 VSS 0.395789f
C820 VIN.n210 VSS 0.569337f
C821 VIN.t6 VSS 0.508132f
C822 VIN.n211 VSS 0.27694f
C823 VOUT.t1 VSS 0.344263f
C824 VOUT.t7 VSS 0.344263f
C825 VOUT.n0 VSS 2.92552f
C826 VOUT.t0 VSS 0.344263f
C827 VOUT.t2 VSS 0.344263f
C828 VOUT.n1 VSS 2.89758f
C829 VOUT.n2 VSS 1.52471f
C830 VOUT.t5 VSS 0.063176f
C831 VOUT.t4 VSS 0.063176f
C832 VOUT.n3 VSS 0.487366f
C833 VOUT.t3 VSS 0.063176f
C834 VOUT.t6 VSS 0.063176f
C835 VOUT.n4 VSS 0.484032f
C836 VOUT.n5 VSS 1.00036f
.ends

