* NGSPICE file created from diff_pair_sample_0200.ext - technology: sky130A

.subckt diff_pair_sample_0200 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t14 VP.t0 VDD1.t4 w_n3320_n3532# sky130_fd_pr__pfet_01v8 ad=2.1153 pd=13.15 as=2.1153 ps=13.15 w=12.82 l=2.02
X1 VDD1.t2 VP.t1 VTAIL.t13 w_n3320_n3532# sky130_fd_pr__pfet_01v8 ad=2.1153 pd=13.15 as=2.1153 ps=13.15 w=12.82 l=2.02
X2 VTAIL.t6 VN.t0 VDD2.t7 w_n3320_n3532# sky130_fd_pr__pfet_01v8 ad=4.9998 pd=26.42 as=2.1153 ps=13.15 w=12.82 l=2.02
X3 VDD2.t6 VN.t1 VTAIL.t0 w_n3320_n3532# sky130_fd_pr__pfet_01v8 ad=2.1153 pd=13.15 as=4.9998 ps=26.42 w=12.82 l=2.02
X4 VTAIL.t12 VP.t2 VDD1.t1 w_n3320_n3532# sky130_fd_pr__pfet_01v8 ad=2.1153 pd=13.15 as=2.1153 ps=13.15 w=12.82 l=2.02
X5 B.t11 B.t9 B.t10 w_n3320_n3532# sky130_fd_pr__pfet_01v8 ad=4.9998 pd=26.42 as=0 ps=0 w=12.82 l=2.02
X6 VTAIL.t11 VP.t3 VDD1.t0 w_n3320_n3532# sky130_fd_pr__pfet_01v8 ad=4.9998 pd=26.42 as=2.1153 ps=13.15 w=12.82 l=2.02
X7 VDD1.t5 VP.t4 VTAIL.t10 w_n3320_n3532# sky130_fd_pr__pfet_01v8 ad=2.1153 pd=13.15 as=4.9998 ps=26.42 w=12.82 l=2.02
X8 B.t8 B.t6 B.t7 w_n3320_n3532# sky130_fd_pr__pfet_01v8 ad=4.9998 pd=26.42 as=0 ps=0 w=12.82 l=2.02
X9 VDD2.t5 VN.t2 VTAIL.t5 w_n3320_n3532# sky130_fd_pr__pfet_01v8 ad=2.1153 pd=13.15 as=4.9998 ps=26.42 w=12.82 l=2.02
X10 B.t5 B.t3 B.t4 w_n3320_n3532# sky130_fd_pr__pfet_01v8 ad=4.9998 pd=26.42 as=0 ps=0 w=12.82 l=2.02
X11 VTAIL.t1 VN.t3 VDD2.t4 w_n3320_n3532# sky130_fd_pr__pfet_01v8 ad=4.9998 pd=26.42 as=2.1153 ps=13.15 w=12.82 l=2.02
X12 VTAIL.t3 VN.t4 VDD2.t3 w_n3320_n3532# sky130_fd_pr__pfet_01v8 ad=2.1153 pd=13.15 as=2.1153 ps=13.15 w=12.82 l=2.02
X13 VDD2.t2 VN.t5 VTAIL.t4 w_n3320_n3532# sky130_fd_pr__pfet_01v8 ad=2.1153 pd=13.15 as=2.1153 ps=13.15 w=12.82 l=2.02
X14 VTAIL.t9 VP.t5 VDD1.t3 w_n3320_n3532# sky130_fd_pr__pfet_01v8 ad=4.9998 pd=26.42 as=2.1153 ps=13.15 w=12.82 l=2.02
X15 VTAIL.t2 VN.t6 VDD2.t1 w_n3320_n3532# sky130_fd_pr__pfet_01v8 ad=2.1153 pd=13.15 as=2.1153 ps=13.15 w=12.82 l=2.02
X16 B.t2 B.t0 B.t1 w_n3320_n3532# sky130_fd_pr__pfet_01v8 ad=4.9998 pd=26.42 as=0 ps=0 w=12.82 l=2.02
X17 VDD2.t0 VN.t7 VTAIL.t15 w_n3320_n3532# sky130_fd_pr__pfet_01v8 ad=2.1153 pd=13.15 as=2.1153 ps=13.15 w=12.82 l=2.02
X18 VDD1.t7 VP.t6 VTAIL.t8 w_n3320_n3532# sky130_fd_pr__pfet_01v8 ad=2.1153 pd=13.15 as=4.9998 ps=26.42 w=12.82 l=2.02
X19 VDD1.t6 VP.t7 VTAIL.t7 w_n3320_n3532# sky130_fd_pr__pfet_01v8 ad=2.1153 pd=13.15 as=2.1153 ps=13.15 w=12.82 l=2.02
R0 VP.n14 VP.t5 184.838
R1 VP.n34 VP.n33 184.427
R2 VP.n60 VP.n59 184.427
R3 VP.n32 VP.n31 184.427
R4 VP.n16 VP.n15 161.3
R5 VP.n17 VP.n12 161.3
R6 VP.n19 VP.n18 161.3
R7 VP.n20 VP.n11 161.3
R8 VP.n22 VP.n21 161.3
R9 VP.n24 VP.n10 161.3
R10 VP.n26 VP.n25 161.3
R11 VP.n27 VP.n9 161.3
R12 VP.n29 VP.n28 161.3
R13 VP.n30 VP.n8 161.3
R14 VP.n58 VP.n0 161.3
R15 VP.n57 VP.n56 161.3
R16 VP.n55 VP.n1 161.3
R17 VP.n54 VP.n53 161.3
R18 VP.n52 VP.n2 161.3
R19 VP.n50 VP.n49 161.3
R20 VP.n48 VP.n3 161.3
R21 VP.n47 VP.n46 161.3
R22 VP.n45 VP.n4 161.3
R23 VP.n44 VP.n43 161.3
R24 VP.n42 VP.n41 161.3
R25 VP.n40 VP.n6 161.3
R26 VP.n39 VP.n38 161.3
R27 VP.n37 VP.n7 161.3
R28 VP.n36 VP.n35 161.3
R29 VP.n34 VP.t3 152.952
R30 VP.n5 VP.t7 152.952
R31 VP.n51 VP.t2 152.952
R32 VP.n59 VP.t6 152.952
R33 VP.n31 VP.t4 152.952
R34 VP.n23 VP.t0 152.952
R35 VP.n13 VP.t1 152.952
R36 VP.n14 VP.n13 61.6806
R37 VP.n40 VP.n39 55.0167
R38 VP.n53 VP.n1 55.0167
R39 VP.n25 VP.n9 55.0167
R40 VP.n33 VP.n32 48.7202
R41 VP.n46 VP.n45 40.4106
R42 VP.n46 VP.n3 40.4106
R43 VP.n18 VP.n11 40.4106
R44 VP.n18 VP.n17 40.4106
R45 VP.n39 VP.n7 25.8045
R46 VP.n57 VP.n1 25.8045
R47 VP.n29 VP.n9 25.8045
R48 VP.n35 VP.n7 24.3439
R49 VP.n41 VP.n40 24.3439
R50 VP.n45 VP.n44 24.3439
R51 VP.n50 VP.n3 24.3439
R52 VP.n53 VP.n52 24.3439
R53 VP.n58 VP.n57 24.3439
R54 VP.n30 VP.n29 24.3439
R55 VP.n22 VP.n11 24.3439
R56 VP.n25 VP.n24 24.3439
R57 VP.n17 VP.n16 24.3439
R58 VP.n41 VP.n5 15.8237
R59 VP.n52 VP.n51 15.8237
R60 VP.n24 VP.n23 15.8237
R61 VP.n15 VP.n14 12.5995
R62 VP.n44 VP.n5 8.5207
R63 VP.n51 VP.n50 8.5207
R64 VP.n23 VP.n22 8.5207
R65 VP.n16 VP.n13 8.5207
R66 VP.n35 VP.n34 1.21767
R67 VP.n59 VP.n58 1.21767
R68 VP.n31 VP.n30 1.21767
R69 VP.n15 VP.n12 0.189894
R70 VP.n19 VP.n12 0.189894
R71 VP.n20 VP.n19 0.189894
R72 VP.n21 VP.n20 0.189894
R73 VP.n21 VP.n10 0.189894
R74 VP.n26 VP.n10 0.189894
R75 VP.n27 VP.n26 0.189894
R76 VP.n28 VP.n27 0.189894
R77 VP.n28 VP.n8 0.189894
R78 VP.n32 VP.n8 0.189894
R79 VP.n36 VP.n33 0.189894
R80 VP.n37 VP.n36 0.189894
R81 VP.n38 VP.n37 0.189894
R82 VP.n38 VP.n6 0.189894
R83 VP.n42 VP.n6 0.189894
R84 VP.n43 VP.n42 0.189894
R85 VP.n43 VP.n4 0.189894
R86 VP.n47 VP.n4 0.189894
R87 VP.n48 VP.n47 0.189894
R88 VP.n49 VP.n48 0.189894
R89 VP.n49 VP.n2 0.189894
R90 VP.n54 VP.n2 0.189894
R91 VP.n55 VP.n54 0.189894
R92 VP.n56 VP.n55 0.189894
R93 VP.n56 VP.n0 0.189894
R94 VP.n60 VP.n0 0.189894
R95 VP VP.n60 0.0516364
R96 VDD1 VDD1.n0 73.6946
R97 VDD1.n3 VDD1.n2 73.5811
R98 VDD1.n3 VDD1.n1 73.5811
R99 VDD1.n5 VDD1.n4 72.6233
R100 VDD1.n5 VDD1.n3 44.4664
R101 VDD1.n4 VDD1.t4 2.53599
R102 VDD1.n4 VDD1.t5 2.53599
R103 VDD1.n0 VDD1.t3 2.53599
R104 VDD1.n0 VDD1.t2 2.53599
R105 VDD1.n2 VDD1.t1 2.53599
R106 VDD1.n2 VDD1.t7 2.53599
R107 VDD1.n1 VDD1.t0 2.53599
R108 VDD1.n1 VDD1.t6 2.53599
R109 VDD1 VDD1.n5 0.955241
R110 VTAIL.n562 VTAIL.n498 756.745
R111 VTAIL.n66 VTAIL.n2 756.745
R112 VTAIL.n136 VTAIL.n72 756.745
R113 VTAIL.n208 VTAIL.n144 756.745
R114 VTAIL.n492 VTAIL.n428 756.745
R115 VTAIL.n420 VTAIL.n356 756.745
R116 VTAIL.n350 VTAIL.n286 756.745
R117 VTAIL.n278 VTAIL.n214 756.745
R118 VTAIL.n521 VTAIL.n520 585
R119 VTAIL.n518 VTAIL.n517 585
R120 VTAIL.n527 VTAIL.n526 585
R121 VTAIL.n529 VTAIL.n528 585
R122 VTAIL.n514 VTAIL.n513 585
R123 VTAIL.n535 VTAIL.n534 585
R124 VTAIL.n538 VTAIL.n537 585
R125 VTAIL.n536 VTAIL.n510 585
R126 VTAIL.n543 VTAIL.n509 585
R127 VTAIL.n545 VTAIL.n544 585
R128 VTAIL.n547 VTAIL.n546 585
R129 VTAIL.n506 VTAIL.n505 585
R130 VTAIL.n553 VTAIL.n552 585
R131 VTAIL.n555 VTAIL.n554 585
R132 VTAIL.n502 VTAIL.n501 585
R133 VTAIL.n561 VTAIL.n560 585
R134 VTAIL.n563 VTAIL.n562 585
R135 VTAIL.n25 VTAIL.n24 585
R136 VTAIL.n22 VTAIL.n21 585
R137 VTAIL.n31 VTAIL.n30 585
R138 VTAIL.n33 VTAIL.n32 585
R139 VTAIL.n18 VTAIL.n17 585
R140 VTAIL.n39 VTAIL.n38 585
R141 VTAIL.n42 VTAIL.n41 585
R142 VTAIL.n40 VTAIL.n14 585
R143 VTAIL.n47 VTAIL.n13 585
R144 VTAIL.n49 VTAIL.n48 585
R145 VTAIL.n51 VTAIL.n50 585
R146 VTAIL.n10 VTAIL.n9 585
R147 VTAIL.n57 VTAIL.n56 585
R148 VTAIL.n59 VTAIL.n58 585
R149 VTAIL.n6 VTAIL.n5 585
R150 VTAIL.n65 VTAIL.n64 585
R151 VTAIL.n67 VTAIL.n66 585
R152 VTAIL.n95 VTAIL.n94 585
R153 VTAIL.n92 VTAIL.n91 585
R154 VTAIL.n101 VTAIL.n100 585
R155 VTAIL.n103 VTAIL.n102 585
R156 VTAIL.n88 VTAIL.n87 585
R157 VTAIL.n109 VTAIL.n108 585
R158 VTAIL.n112 VTAIL.n111 585
R159 VTAIL.n110 VTAIL.n84 585
R160 VTAIL.n117 VTAIL.n83 585
R161 VTAIL.n119 VTAIL.n118 585
R162 VTAIL.n121 VTAIL.n120 585
R163 VTAIL.n80 VTAIL.n79 585
R164 VTAIL.n127 VTAIL.n126 585
R165 VTAIL.n129 VTAIL.n128 585
R166 VTAIL.n76 VTAIL.n75 585
R167 VTAIL.n135 VTAIL.n134 585
R168 VTAIL.n137 VTAIL.n136 585
R169 VTAIL.n167 VTAIL.n166 585
R170 VTAIL.n164 VTAIL.n163 585
R171 VTAIL.n173 VTAIL.n172 585
R172 VTAIL.n175 VTAIL.n174 585
R173 VTAIL.n160 VTAIL.n159 585
R174 VTAIL.n181 VTAIL.n180 585
R175 VTAIL.n184 VTAIL.n183 585
R176 VTAIL.n182 VTAIL.n156 585
R177 VTAIL.n189 VTAIL.n155 585
R178 VTAIL.n191 VTAIL.n190 585
R179 VTAIL.n193 VTAIL.n192 585
R180 VTAIL.n152 VTAIL.n151 585
R181 VTAIL.n199 VTAIL.n198 585
R182 VTAIL.n201 VTAIL.n200 585
R183 VTAIL.n148 VTAIL.n147 585
R184 VTAIL.n207 VTAIL.n206 585
R185 VTAIL.n209 VTAIL.n208 585
R186 VTAIL.n493 VTAIL.n492 585
R187 VTAIL.n491 VTAIL.n490 585
R188 VTAIL.n432 VTAIL.n431 585
R189 VTAIL.n485 VTAIL.n484 585
R190 VTAIL.n483 VTAIL.n482 585
R191 VTAIL.n436 VTAIL.n435 585
R192 VTAIL.n477 VTAIL.n476 585
R193 VTAIL.n475 VTAIL.n474 585
R194 VTAIL.n473 VTAIL.n439 585
R195 VTAIL.n443 VTAIL.n440 585
R196 VTAIL.n468 VTAIL.n467 585
R197 VTAIL.n466 VTAIL.n465 585
R198 VTAIL.n445 VTAIL.n444 585
R199 VTAIL.n460 VTAIL.n459 585
R200 VTAIL.n458 VTAIL.n457 585
R201 VTAIL.n449 VTAIL.n448 585
R202 VTAIL.n452 VTAIL.n451 585
R203 VTAIL.n421 VTAIL.n420 585
R204 VTAIL.n419 VTAIL.n418 585
R205 VTAIL.n360 VTAIL.n359 585
R206 VTAIL.n413 VTAIL.n412 585
R207 VTAIL.n411 VTAIL.n410 585
R208 VTAIL.n364 VTAIL.n363 585
R209 VTAIL.n405 VTAIL.n404 585
R210 VTAIL.n403 VTAIL.n402 585
R211 VTAIL.n401 VTAIL.n367 585
R212 VTAIL.n371 VTAIL.n368 585
R213 VTAIL.n396 VTAIL.n395 585
R214 VTAIL.n394 VTAIL.n393 585
R215 VTAIL.n373 VTAIL.n372 585
R216 VTAIL.n388 VTAIL.n387 585
R217 VTAIL.n386 VTAIL.n385 585
R218 VTAIL.n377 VTAIL.n376 585
R219 VTAIL.n380 VTAIL.n379 585
R220 VTAIL.n351 VTAIL.n350 585
R221 VTAIL.n349 VTAIL.n348 585
R222 VTAIL.n290 VTAIL.n289 585
R223 VTAIL.n343 VTAIL.n342 585
R224 VTAIL.n341 VTAIL.n340 585
R225 VTAIL.n294 VTAIL.n293 585
R226 VTAIL.n335 VTAIL.n334 585
R227 VTAIL.n333 VTAIL.n332 585
R228 VTAIL.n331 VTAIL.n297 585
R229 VTAIL.n301 VTAIL.n298 585
R230 VTAIL.n326 VTAIL.n325 585
R231 VTAIL.n324 VTAIL.n323 585
R232 VTAIL.n303 VTAIL.n302 585
R233 VTAIL.n318 VTAIL.n317 585
R234 VTAIL.n316 VTAIL.n315 585
R235 VTAIL.n307 VTAIL.n306 585
R236 VTAIL.n310 VTAIL.n309 585
R237 VTAIL.n279 VTAIL.n278 585
R238 VTAIL.n277 VTAIL.n276 585
R239 VTAIL.n218 VTAIL.n217 585
R240 VTAIL.n271 VTAIL.n270 585
R241 VTAIL.n269 VTAIL.n268 585
R242 VTAIL.n222 VTAIL.n221 585
R243 VTAIL.n263 VTAIL.n262 585
R244 VTAIL.n261 VTAIL.n260 585
R245 VTAIL.n259 VTAIL.n225 585
R246 VTAIL.n229 VTAIL.n226 585
R247 VTAIL.n254 VTAIL.n253 585
R248 VTAIL.n252 VTAIL.n251 585
R249 VTAIL.n231 VTAIL.n230 585
R250 VTAIL.n246 VTAIL.n245 585
R251 VTAIL.n244 VTAIL.n243 585
R252 VTAIL.n235 VTAIL.n234 585
R253 VTAIL.n238 VTAIL.n237 585
R254 VTAIL.t0 VTAIL.n519 329.036
R255 VTAIL.t1 VTAIL.n23 329.036
R256 VTAIL.t8 VTAIL.n93 329.036
R257 VTAIL.t11 VTAIL.n165 329.036
R258 VTAIL.t10 VTAIL.n450 329.036
R259 VTAIL.t9 VTAIL.n378 329.036
R260 VTAIL.t5 VTAIL.n308 329.036
R261 VTAIL.t6 VTAIL.n236 329.036
R262 VTAIL.n520 VTAIL.n517 171.744
R263 VTAIL.n527 VTAIL.n517 171.744
R264 VTAIL.n528 VTAIL.n527 171.744
R265 VTAIL.n528 VTAIL.n513 171.744
R266 VTAIL.n535 VTAIL.n513 171.744
R267 VTAIL.n537 VTAIL.n535 171.744
R268 VTAIL.n537 VTAIL.n536 171.744
R269 VTAIL.n536 VTAIL.n509 171.744
R270 VTAIL.n545 VTAIL.n509 171.744
R271 VTAIL.n546 VTAIL.n545 171.744
R272 VTAIL.n546 VTAIL.n505 171.744
R273 VTAIL.n553 VTAIL.n505 171.744
R274 VTAIL.n554 VTAIL.n553 171.744
R275 VTAIL.n554 VTAIL.n501 171.744
R276 VTAIL.n561 VTAIL.n501 171.744
R277 VTAIL.n562 VTAIL.n561 171.744
R278 VTAIL.n24 VTAIL.n21 171.744
R279 VTAIL.n31 VTAIL.n21 171.744
R280 VTAIL.n32 VTAIL.n31 171.744
R281 VTAIL.n32 VTAIL.n17 171.744
R282 VTAIL.n39 VTAIL.n17 171.744
R283 VTAIL.n41 VTAIL.n39 171.744
R284 VTAIL.n41 VTAIL.n40 171.744
R285 VTAIL.n40 VTAIL.n13 171.744
R286 VTAIL.n49 VTAIL.n13 171.744
R287 VTAIL.n50 VTAIL.n49 171.744
R288 VTAIL.n50 VTAIL.n9 171.744
R289 VTAIL.n57 VTAIL.n9 171.744
R290 VTAIL.n58 VTAIL.n57 171.744
R291 VTAIL.n58 VTAIL.n5 171.744
R292 VTAIL.n65 VTAIL.n5 171.744
R293 VTAIL.n66 VTAIL.n65 171.744
R294 VTAIL.n94 VTAIL.n91 171.744
R295 VTAIL.n101 VTAIL.n91 171.744
R296 VTAIL.n102 VTAIL.n101 171.744
R297 VTAIL.n102 VTAIL.n87 171.744
R298 VTAIL.n109 VTAIL.n87 171.744
R299 VTAIL.n111 VTAIL.n109 171.744
R300 VTAIL.n111 VTAIL.n110 171.744
R301 VTAIL.n110 VTAIL.n83 171.744
R302 VTAIL.n119 VTAIL.n83 171.744
R303 VTAIL.n120 VTAIL.n119 171.744
R304 VTAIL.n120 VTAIL.n79 171.744
R305 VTAIL.n127 VTAIL.n79 171.744
R306 VTAIL.n128 VTAIL.n127 171.744
R307 VTAIL.n128 VTAIL.n75 171.744
R308 VTAIL.n135 VTAIL.n75 171.744
R309 VTAIL.n136 VTAIL.n135 171.744
R310 VTAIL.n166 VTAIL.n163 171.744
R311 VTAIL.n173 VTAIL.n163 171.744
R312 VTAIL.n174 VTAIL.n173 171.744
R313 VTAIL.n174 VTAIL.n159 171.744
R314 VTAIL.n181 VTAIL.n159 171.744
R315 VTAIL.n183 VTAIL.n181 171.744
R316 VTAIL.n183 VTAIL.n182 171.744
R317 VTAIL.n182 VTAIL.n155 171.744
R318 VTAIL.n191 VTAIL.n155 171.744
R319 VTAIL.n192 VTAIL.n191 171.744
R320 VTAIL.n192 VTAIL.n151 171.744
R321 VTAIL.n199 VTAIL.n151 171.744
R322 VTAIL.n200 VTAIL.n199 171.744
R323 VTAIL.n200 VTAIL.n147 171.744
R324 VTAIL.n207 VTAIL.n147 171.744
R325 VTAIL.n208 VTAIL.n207 171.744
R326 VTAIL.n492 VTAIL.n491 171.744
R327 VTAIL.n491 VTAIL.n431 171.744
R328 VTAIL.n484 VTAIL.n431 171.744
R329 VTAIL.n484 VTAIL.n483 171.744
R330 VTAIL.n483 VTAIL.n435 171.744
R331 VTAIL.n476 VTAIL.n435 171.744
R332 VTAIL.n476 VTAIL.n475 171.744
R333 VTAIL.n475 VTAIL.n439 171.744
R334 VTAIL.n443 VTAIL.n439 171.744
R335 VTAIL.n467 VTAIL.n443 171.744
R336 VTAIL.n467 VTAIL.n466 171.744
R337 VTAIL.n466 VTAIL.n444 171.744
R338 VTAIL.n459 VTAIL.n444 171.744
R339 VTAIL.n459 VTAIL.n458 171.744
R340 VTAIL.n458 VTAIL.n448 171.744
R341 VTAIL.n451 VTAIL.n448 171.744
R342 VTAIL.n420 VTAIL.n419 171.744
R343 VTAIL.n419 VTAIL.n359 171.744
R344 VTAIL.n412 VTAIL.n359 171.744
R345 VTAIL.n412 VTAIL.n411 171.744
R346 VTAIL.n411 VTAIL.n363 171.744
R347 VTAIL.n404 VTAIL.n363 171.744
R348 VTAIL.n404 VTAIL.n403 171.744
R349 VTAIL.n403 VTAIL.n367 171.744
R350 VTAIL.n371 VTAIL.n367 171.744
R351 VTAIL.n395 VTAIL.n371 171.744
R352 VTAIL.n395 VTAIL.n394 171.744
R353 VTAIL.n394 VTAIL.n372 171.744
R354 VTAIL.n387 VTAIL.n372 171.744
R355 VTAIL.n387 VTAIL.n386 171.744
R356 VTAIL.n386 VTAIL.n376 171.744
R357 VTAIL.n379 VTAIL.n376 171.744
R358 VTAIL.n350 VTAIL.n349 171.744
R359 VTAIL.n349 VTAIL.n289 171.744
R360 VTAIL.n342 VTAIL.n289 171.744
R361 VTAIL.n342 VTAIL.n341 171.744
R362 VTAIL.n341 VTAIL.n293 171.744
R363 VTAIL.n334 VTAIL.n293 171.744
R364 VTAIL.n334 VTAIL.n333 171.744
R365 VTAIL.n333 VTAIL.n297 171.744
R366 VTAIL.n301 VTAIL.n297 171.744
R367 VTAIL.n325 VTAIL.n301 171.744
R368 VTAIL.n325 VTAIL.n324 171.744
R369 VTAIL.n324 VTAIL.n302 171.744
R370 VTAIL.n317 VTAIL.n302 171.744
R371 VTAIL.n317 VTAIL.n316 171.744
R372 VTAIL.n316 VTAIL.n306 171.744
R373 VTAIL.n309 VTAIL.n306 171.744
R374 VTAIL.n278 VTAIL.n277 171.744
R375 VTAIL.n277 VTAIL.n217 171.744
R376 VTAIL.n270 VTAIL.n217 171.744
R377 VTAIL.n270 VTAIL.n269 171.744
R378 VTAIL.n269 VTAIL.n221 171.744
R379 VTAIL.n262 VTAIL.n221 171.744
R380 VTAIL.n262 VTAIL.n261 171.744
R381 VTAIL.n261 VTAIL.n225 171.744
R382 VTAIL.n229 VTAIL.n225 171.744
R383 VTAIL.n253 VTAIL.n229 171.744
R384 VTAIL.n253 VTAIL.n252 171.744
R385 VTAIL.n252 VTAIL.n230 171.744
R386 VTAIL.n245 VTAIL.n230 171.744
R387 VTAIL.n245 VTAIL.n244 171.744
R388 VTAIL.n244 VTAIL.n234 171.744
R389 VTAIL.n237 VTAIL.n234 171.744
R390 VTAIL.n520 VTAIL.t0 85.8723
R391 VTAIL.n24 VTAIL.t1 85.8723
R392 VTAIL.n94 VTAIL.t8 85.8723
R393 VTAIL.n166 VTAIL.t11 85.8723
R394 VTAIL.n451 VTAIL.t10 85.8723
R395 VTAIL.n379 VTAIL.t9 85.8723
R396 VTAIL.n309 VTAIL.t5 85.8723
R397 VTAIL.n237 VTAIL.t6 85.8723
R398 VTAIL.n1 VTAIL.n0 55.9447
R399 VTAIL.n143 VTAIL.n142 55.9447
R400 VTAIL.n427 VTAIL.n426 55.9447
R401 VTAIL.n285 VTAIL.n284 55.9447
R402 VTAIL.n567 VTAIL.n566 31.7975
R403 VTAIL.n71 VTAIL.n70 31.7975
R404 VTAIL.n141 VTAIL.n140 31.7975
R405 VTAIL.n213 VTAIL.n212 31.7975
R406 VTAIL.n497 VTAIL.n496 31.7975
R407 VTAIL.n425 VTAIL.n424 31.7975
R408 VTAIL.n355 VTAIL.n354 31.7975
R409 VTAIL.n283 VTAIL.n282 31.7975
R410 VTAIL.n567 VTAIL.n497 25.4445
R411 VTAIL.n283 VTAIL.n213 25.4445
R412 VTAIL.n544 VTAIL.n543 13.1884
R413 VTAIL.n48 VTAIL.n47 13.1884
R414 VTAIL.n118 VTAIL.n117 13.1884
R415 VTAIL.n190 VTAIL.n189 13.1884
R416 VTAIL.n474 VTAIL.n473 13.1884
R417 VTAIL.n402 VTAIL.n401 13.1884
R418 VTAIL.n332 VTAIL.n331 13.1884
R419 VTAIL.n260 VTAIL.n259 13.1884
R420 VTAIL.n542 VTAIL.n510 12.8005
R421 VTAIL.n547 VTAIL.n508 12.8005
R422 VTAIL.n46 VTAIL.n14 12.8005
R423 VTAIL.n51 VTAIL.n12 12.8005
R424 VTAIL.n116 VTAIL.n84 12.8005
R425 VTAIL.n121 VTAIL.n82 12.8005
R426 VTAIL.n188 VTAIL.n156 12.8005
R427 VTAIL.n193 VTAIL.n154 12.8005
R428 VTAIL.n477 VTAIL.n438 12.8005
R429 VTAIL.n472 VTAIL.n440 12.8005
R430 VTAIL.n405 VTAIL.n366 12.8005
R431 VTAIL.n400 VTAIL.n368 12.8005
R432 VTAIL.n335 VTAIL.n296 12.8005
R433 VTAIL.n330 VTAIL.n298 12.8005
R434 VTAIL.n263 VTAIL.n224 12.8005
R435 VTAIL.n258 VTAIL.n226 12.8005
R436 VTAIL.n539 VTAIL.n538 12.0247
R437 VTAIL.n548 VTAIL.n506 12.0247
R438 VTAIL.n43 VTAIL.n42 12.0247
R439 VTAIL.n52 VTAIL.n10 12.0247
R440 VTAIL.n113 VTAIL.n112 12.0247
R441 VTAIL.n122 VTAIL.n80 12.0247
R442 VTAIL.n185 VTAIL.n184 12.0247
R443 VTAIL.n194 VTAIL.n152 12.0247
R444 VTAIL.n478 VTAIL.n436 12.0247
R445 VTAIL.n469 VTAIL.n468 12.0247
R446 VTAIL.n406 VTAIL.n364 12.0247
R447 VTAIL.n397 VTAIL.n396 12.0247
R448 VTAIL.n336 VTAIL.n294 12.0247
R449 VTAIL.n327 VTAIL.n326 12.0247
R450 VTAIL.n264 VTAIL.n222 12.0247
R451 VTAIL.n255 VTAIL.n254 12.0247
R452 VTAIL.n534 VTAIL.n512 11.249
R453 VTAIL.n552 VTAIL.n551 11.249
R454 VTAIL.n38 VTAIL.n16 11.249
R455 VTAIL.n56 VTAIL.n55 11.249
R456 VTAIL.n108 VTAIL.n86 11.249
R457 VTAIL.n126 VTAIL.n125 11.249
R458 VTAIL.n180 VTAIL.n158 11.249
R459 VTAIL.n198 VTAIL.n197 11.249
R460 VTAIL.n482 VTAIL.n481 11.249
R461 VTAIL.n465 VTAIL.n442 11.249
R462 VTAIL.n410 VTAIL.n409 11.249
R463 VTAIL.n393 VTAIL.n370 11.249
R464 VTAIL.n340 VTAIL.n339 11.249
R465 VTAIL.n323 VTAIL.n300 11.249
R466 VTAIL.n268 VTAIL.n267 11.249
R467 VTAIL.n251 VTAIL.n228 11.249
R468 VTAIL.n521 VTAIL.n519 10.7239
R469 VTAIL.n25 VTAIL.n23 10.7239
R470 VTAIL.n95 VTAIL.n93 10.7239
R471 VTAIL.n167 VTAIL.n165 10.7239
R472 VTAIL.n452 VTAIL.n450 10.7239
R473 VTAIL.n380 VTAIL.n378 10.7239
R474 VTAIL.n310 VTAIL.n308 10.7239
R475 VTAIL.n238 VTAIL.n236 10.7239
R476 VTAIL.n533 VTAIL.n514 10.4732
R477 VTAIL.n555 VTAIL.n504 10.4732
R478 VTAIL.n37 VTAIL.n18 10.4732
R479 VTAIL.n59 VTAIL.n8 10.4732
R480 VTAIL.n107 VTAIL.n88 10.4732
R481 VTAIL.n129 VTAIL.n78 10.4732
R482 VTAIL.n179 VTAIL.n160 10.4732
R483 VTAIL.n201 VTAIL.n150 10.4732
R484 VTAIL.n485 VTAIL.n434 10.4732
R485 VTAIL.n464 VTAIL.n445 10.4732
R486 VTAIL.n413 VTAIL.n362 10.4732
R487 VTAIL.n392 VTAIL.n373 10.4732
R488 VTAIL.n343 VTAIL.n292 10.4732
R489 VTAIL.n322 VTAIL.n303 10.4732
R490 VTAIL.n271 VTAIL.n220 10.4732
R491 VTAIL.n250 VTAIL.n231 10.4732
R492 VTAIL.n530 VTAIL.n529 9.69747
R493 VTAIL.n556 VTAIL.n502 9.69747
R494 VTAIL.n34 VTAIL.n33 9.69747
R495 VTAIL.n60 VTAIL.n6 9.69747
R496 VTAIL.n104 VTAIL.n103 9.69747
R497 VTAIL.n130 VTAIL.n76 9.69747
R498 VTAIL.n176 VTAIL.n175 9.69747
R499 VTAIL.n202 VTAIL.n148 9.69747
R500 VTAIL.n486 VTAIL.n432 9.69747
R501 VTAIL.n461 VTAIL.n460 9.69747
R502 VTAIL.n414 VTAIL.n360 9.69747
R503 VTAIL.n389 VTAIL.n388 9.69747
R504 VTAIL.n344 VTAIL.n290 9.69747
R505 VTAIL.n319 VTAIL.n318 9.69747
R506 VTAIL.n272 VTAIL.n218 9.69747
R507 VTAIL.n247 VTAIL.n246 9.69747
R508 VTAIL.n566 VTAIL.n565 9.45567
R509 VTAIL.n70 VTAIL.n69 9.45567
R510 VTAIL.n140 VTAIL.n139 9.45567
R511 VTAIL.n212 VTAIL.n211 9.45567
R512 VTAIL.n496 VTAIL.n495 9.45567
R513 VTAIL.n424 VTAIL.n423 9.45567
R514 VTAIL.n354 VTAIL.n353 9.45567
R515 VTAIL.n282 VTAIL.n281 9.45567
R516 VTAIL.n500 VTAIL.n499 9.3005
R517 VTAIL.n559 VTAIL.n558 9.3005
R518 VTAIL.n557 VTAIL.n556 9.3005
R519 VTAIL.n504 VTAIL.n503 9.3005
R520 VTAIL.n551 VTAIL.n550 9.3005
R521 VTAIL.n549 VTAIL.n548 9.3005
R522 VTAIL.n508 VTAIL.n507 9.3005
R523 VTAIL.n523 VTAIL.n522 9.3005
R524 VTAIL.n525 VTAIL.n524 9.3005
R525 VTAIL.n516 VTAIL.n515 9.3005
R526 VTAIL.n531 VTAIL.n530 9.3005
R527 VTAIL.n533 VTAIL.n532 9.3005
R528 VTAIL.n512 VTAIL.n511 9.3005
R529 VTAIL.n540 VTAIL.n539 9.3005
R530 VTAIL.n542 VTAIL.n541 9.3005
R531 VTAIL.n565 VTAIL.n564 9.3005
R532 VTAIL.n4 VTAIL.n3 9.3005
R533 VTAIL.n63 VTAIL.n62 9.3005
R534 VTAIL.n61 VTAIL.n60 9.3005
R535 VTAIL.n8 VTAIL.n7 9.3005
R536 VTAIL.n55 VTAIL.n54 9.3005
R537 VTAIL.n53 VTAIL.n52 9.3005
R538 VTAIL.n12 VTAIL.n11 9.3005
R539 VTAIL.n27 VTAIL.n26 9.3005
R540 VTAIL.n29 VTAIL.n28 9.3005
R541 VTAIL.n20 VTAIL.n19 9.3005
R542 VTAIL.n35 VTAIL.n34 9.3005
R543 VTAIL.n37 VTAIL.n36 9.3005
R544 VTAIL.n16 VTAIL.n15 9.3005
R545 VTAIL.n44 VTAIL.n43 9.3005
R546 VTAIL.n46 VTAIL.n45 9.3005
R547 VTAIL.n69 VTAIL.n68 9.3005
R548 VTAIL.n74 VTAIL.n73 9.3005
R549 VTAIL.n133 VTAIL.n132 9.3005
R550 VTAIL.n131 VTAIL.n130 9.3005
R551 VTAIL.n78 VTAIL.n77 9.3005
R552 VTAIL.n125 VTAIL.n124 9.3005
R553 VTAIL.n123 VTAIL.n122 9.3005
R554 VTAIL.n82 VTAIL.n81 9.3005
R555 VTAIL.n97 VTAIL.n96 9.3005
R556 VTAIL.n99 VTAIL.n98 9.3005
R557 VTAIL.n90 VTAIL.n89 9.3005
R558 VTAIL.n105 VTAIL.n104 9.3005
R559 VTAIL.n107 VTAIL.n106 9.3005
R560 VTAIL.n86 VTAIL.n85 9.3005
R561 VTAIL.n114 VTAIL.n113 9.3005
R562 VTAIL.n116 VTAIL.n115 9.3005
R563 VTAIL.n139 VTAIL.n138 9.3005
R564 VTAIL.n146 VTAIL.n145 9.3005
R565 VTAIL.n205 VTAIL.n204 9.3005
R566 VTAIL.n203 VTAIL.n202 9.3005
R567 VTAIL.n150 VTAIL.n149 9.3005
R568 VTAIL.n197 VTAIL.n196 9.3005
R569 VTAIL.n195 VTAIL.n194 9.3005
R570 VTAIL.n154 VTAIL.n153 9.3005
R571 VTAIL.n169 VTAIL.n168 9.3005
R572 VTAIL.n171 VTAIL.n170 9.3005
R573 VTAIL.n162 VTAIL.n161 9.3005
R574 VTAIL.n177 VTAIL.n176 9.3005
R575 VTAIL.n179 VTAIL.n178 9.3005
R576 VTAIL.n158 VTAIL.n157 9.3005
R577 VTAIL.n186 VTAIL.n185 9.3005
R578 VTAIL.n188 VTAIL.n187 9.3005
R579 VTAIL.n211 VTAIL.n210 9.3005
R580 VTAIL.n454 VTAIL.n453 9.3005
R581 VTAIL.n456 VTAIL.n455 9.3005
R582 VTAIL.n447 VTAIL.n446 9.3005
R583 VTAIL.n462 VTAIL.n461 9.3005
R584 VTAIL.n464 VTAIL.n463 9.3005
R585 VTAIL.n442 VTAIL.n441 9.3005
R586 VTAIL.n470 VTAIL.n469 9.3005
R587 VTAIL.n472 VTAIL.n471 9.3005
R588 VTAIL.n495 VTAIL.n494 9.3005
R589 VTAIL.n430 VTAIL.n429 9.3005
R590 VTAIL.n489 VTAIL.n488 9.3005
R591 VTAIL.n487 VTAIL.n486 9.3005
R592 VTAIL.n434 VTAIL.n433 9.3005
R593 VTAIL.n481 VTAIL.n480 9.3005
R594 VTAIL.n479 VTAIL.n478 9.3005
R595 VTAIL.n438 VTAIL.n437 9.3005
R596 VTAIL.n382 VTAIL.n381 9.3005
R597 VTAIL.n384 VTAIL.n383 9.3005
R598 VTAIL.n375 VTAIL.n374 9.3005
R599 VTAIL.n390 VTAIL.n389 9.3005
R600 VTAIL.n392 VTAIL.n391 9.3005
R601 VTAIL.n370 VTAIL.n369 9.3005
R602 VTAIL.n398 VTAIL.n397 9.3005
R603 VTAIL.n400 VTAIL.n399 9.3005
R604 VTAIL.n423 VTAIL.n422 9.3005
R605 VTAIL.n358 VTAIL.n357 9.3005
R606 VTAIL.n417 VTAIL.n416 9.3005
R607 VTAIL.n415 VTAIL.n414 9.3005
R608 VTAIL.n362 VTAIL.n361 9.3005
R609 VTAIL.n409 VTAIL.n408 9.3005
R610 VTAIL.n407 VTAIL.n406 9.3005
R611 VTAIL.n366 VTAIL.n365 9.3005
R612 VTAIL.n312 VTAIL.n311 9.3005
R613 VTAIL.n314 VTAIL.n313 9.3005
R614 VTAIL.n305 VTAIL.n304 9.3005
R615 VTAIL.n320 VTAIL.n319 9.3005
R616 VTAIL.n322 VTAIL.n321 9.3005
R617 VTAIL.n300 VTAIL.n299 9.3005
R618 VTAIL.n328 VTAIL.n327 9.3005
R619 VTAIL.n330 VTAIL.n329 9.3005
R620 VTAIL.n353 VTAIL.n352 9.3005
R621 VTAIL.n288 VTAIL.n287 9.3005
R622 VTAIL.n347 VTAIL.n346 9.3005
R623 VTAIL.n345 VTAIL.n344 9.3005
R624 VTAIL.n292 VTAIL.n291 9.3005
R625 VTAIL.n339 VTAIL.n338 9.3005
R626 VTAIL.n337 VTAIL.n336 9.3005
R627 VTAIL.n296 VTAIL.n295 9.3005
R628 VTAIL.n240 VTAIL.n239 9.3005
R629 VTAIL.n242 VTAIL.n241 9.3005
R630 VTAIL.n233 VTAIL.n232 9.3005
R631 VTAIL.n248 VTAIL.n247 9.3005
R632 VTAIL.n250 VTAIL.n249 9.3005
R633 VTAIL.n228 VTAIL.n227 9.3005
R634 VTAIL.n256 VTAIL.n255 9.3005
R635 VTAIL.n258 VTAIL.n257 9.3005
R636 VTAIL.n281 VTAIL.n280 9.3005
R637 VTAIL.n216 VTAIL.n215 9.3005
R638 VTAIL.n275 VTAIL.n274 9.3005
R639 VTAIL.n273 VTAIL.n272 9.3005
R640 VTAIL.n220 VTAIL.n219 9.3005
R641 VTAIL.n267 VTAIL.n266 9.3005
R642 VTAIL.n265 VTAIL.n264 9.3005
R643 VTAIL.n224 VTAIL.n223 9.3005
R644 VTAIL.n526 VTAIL.n516 8.92171
R645 VTAIL.n560 VTAIL.n559 8.92171
R646 VTAIL.n30 VTAIL.n20 8.92171
R647 VTAIL.n64 VTAIL.n63 8.92171
R648 VTAIL.n100 VTAIL.n90 8.92171
R649 VTAIL.n134 VTAIL.n133 8.92171
R650 VTAIL.n172 VTAIL.n162 8.92171
R651 VTAIL.n206 VTAIL.n205 8.92171
R652 VTAIL.n490 VTAIL.n489 8.92171
R653 VTAIL.n457 VTAIL.n447 8.92171
R654 VTAIL.n418 VTAIL.n417 8.92171
R655 VTAIL.n385 VTAIL.n375 8.92171
R656 VTAIL.n348 VTAIL.n347 8.92171
R657 VTAIL.n315 VTAIL.n305 8.92171
R658 VTAIL.n276 VTAIL.n275 8.92171
R659 VTAIL.n243 VTAIL.n233 8.92171
R660 VTAIL.n525 VTAIL.n518 8.14595
R661 VTAIL.n563 VTAIL.n500 8.14595
R662 VTAIL.n29 VTAIL.n22 8.14595
R663 VTAIL.n67 VTAIL.n4 8.14595
R664 VTAIL.n99 VTAIL.n92 8.14595
R665 VTAIL.n137 VTAIL.n74 8.14595
R666 VTAIL.n171 VTAIL.n164 8.14595
R667 VTAIL.n209 VTAIL.n146 8.14595
R668 VTAIL.n493 VTAIL.n430 8.14595
R669 VTAIL.n456 VTAIL.n449 8.14595
R670 VTAIL.n421 VTAIL.n358 8.14595
R671 VTAIL.n384 VTAIL.n377 8.14595
R672 VTAIL.n351 VTAIL.n288 8.14595
R673 VTAIL.n314 VTAIL.n307 8.14595
R674 VTAIL.n279 VTAIL.n216 8.14595
R675 VTAIL.n242 VTAIL.n235 8.14595
R676 VTAIL.n522 VTAIL.n521 7.3702
R677 VTAIL.n564 VTAIL.n498 7.3702
R678 VTAIL.n26 VTAIL.n25 7.3702
R679 VTAIL.n68 VTAIL.n2 7.3702
R680 VTAIL.n96 VTAIL.n95 7.3702
R681 VTAIL.n138 VTAIL.n72 7.3702
R682 VTAIL.n168 VTAIL.n167 7.3702
R683 VTAIL.n210 VTAIL.n144 7.3702
R684 VTAIL.n494 VTAIL.n428 7.3702
R685 VTAIL.n453 VTAIL.n452 7.3702
R686 VTAIL.n422 VTAIL.n356 7.3702
R687 VTAIL.n381 VTAIL.n380 7.3702
R688 VTAIL.n352 VTAIL.n286 7.3702
R689 VTAIL.n311 VTAIL.n310 7.3702
R690 VTAIL.n280 VTAIL.n214 7.3702
R691 VTAIL.n239 VTAIL.n238 7.3702
R692 VTAIL.n566 VTAIL.n498 6.59444
R693 VTAIL.n70 VTAIL.n2 6.59444
R694 VTAIL.n140 VTAIL.n72 6.59444
R695 VTAIL.n212 VTAIL.n144 6.59444
R696 VTAIL.n496 VTAIL.n428 6.59444
R697 VTAIL.n424 VTAIL.n356 6.59444
R698 VTAIL.n354 VTAIL.n286 6.59444
R699 VTAIL.n282 VTAIL.n214 6.59444
R700 VTAIL.n522 VTAIL.n518 5.81868
R701 VTAIL.n564 VTAIL.n563 5.81868
R702 VTAIL.n26 VTAIL.n22 5.81868
R703 VTAIL.n68 VTAIL.n67 5.81868
R704 VTAIL.n96 VTAIL.n92 5.81868
R705 VTAIL.n138 VTAIL.n137 5.81868
R706 VTAIL.n168 VTAIL.n164 5.81868
R707 VTAIL.n210 VTAIL.n209 5.81868
R708 VTAIL.n494 VTAIL.n493 5.81868
R709 VTAIL.n453 VTAIL.n449 5.81868
R710 VTAIL.n422 VTAIL.n421 5.81868
R711 VTAIL.n381 VTAIL.n377 5.81868
R712 VTAIL.n352 VTAIL.n351 5.81868
R713 VTAIL.n311 VTAIL.n307 5.81868
R714 VTAIL.n280 VTAIL.n279 5.81868
R715 VTAIL.n239 VTAIL.n235 5.81868
R716 VTAIL.n526 VTAIL.n525 5.04292
R717 VTAIL.n560 VTAIL.n500 5.04292
R718 VTAIL.n30 VTAIL.n29 5.04292
R719 VTAIL.n64 VTAIL.n4 5.04292
R720 VTAIL.n100 VTAIL.n99 5.04292
R721 VTAIL.n134 VTAIL.n74 5.04292
R722 VTAIL.n172 VTAIL.n171 5.04292
R723 VTAIL.n206 VTAIL.n146 5.04292
R724 VTAIL.n490 VTAIL.n430 5.04292
R725 VTAIL.n457 VTAIL.n456 5.04292
R726 VTAIL.n418 VTAIL.n358 5.04292
R727 VTAIL.n385 VTAIL.n384 5.04292
R728 VTAIL.n348 VTAIL.n288 5.04292
R729 VTAIL.n315 VTAIL.n314 5.04292
R730 VTAIL.n276 VTAIL.n216 5.04292
R731 VTAIL.n243 VTAIL.n242 5.04292
R732 VTAIL.n529 VTAIL.n516 4.26717
R733 VTAIL.n559 VTAIL.n502 4.26717
R734 VTAIL.n33 VTAIL.n20 4.26717
R735 VTAIL.n63 VTAIL.n6 4.26717
R736 VTAIL.n103 VTAIL.n90 4.26717
R737 VTAIL.n133 VTAIL.n76 4.26717
R738 VTAIL.n175 VTAIL.n162 4.26717
R739 VTAIL.n205 VTAIL.n148 4.26717
R740 VTAIL.n489 VTAIL.n432 4.26717
R741 VTAIL.n460 VTAIL.n447 4.26717
R742 VTAIL.n417 VTAIL.n360 4.26717
R743 VTAIL.n388 VTAIL.n375 4.26717
R744 VTAIL.n347 VTAIL.n290 4.26717
R745 VTAIL.n318 VTAIL.n305 4.26717
R746 VTAIL.n275 VTAIL.n218 4.26717
R747 VTAIL.n246 VTAIL.n233 4.26717
R748 VTAIL.n530 VTAIL.n514 3.49141
R749 VTAIL.n556 VTAIL.n555 3.49141
R750 VTAIL.n34 VTAIL.n18 3.49141
R751 VTAIL.n60 VTAIL.n59 3.49141
R752 VTAIL.n104 VTAIL.n88 3.49141
R753 VTAIL.n130 VTAIL.n129 3.49141
R754 VTAIL.n176 VTAIL.n160 3.49141
R755 VTAIL.n202 VTAIL.n201 3.49141
R756 VTAIL.n486 VTAIL.n485 3.49141
R757 VTAIL.n461 VTAIL.n445 3.49141
R758 VTAIL.n414 VTAIL.n413 3.49141
R759 VTAIL.n389 VTAIL.n373 3.49141
R760 VTAIL.n344 VTAIL.n343 3.49141
R761 VTAIL.n319 VTAIL.n303 3.49141
R762 VTAIL.n272 VTAIL.n271 3.49141
R763 VTAIL.n247 VTAIL.n231 3.49141
R764 VTAIL.n534 VTAIL.n533 2.71565
R765 VTAIL.n552 VTAIL.n504 2.71565
R766 VTAIL.n38 VTAIL.n37 2.71565
R767 VTAIL.n56 VTAIL.n8 2.71565
R768 VTAIL.n108 VTAIL.n107 2.71565
R769 VTAIL.n126 VTAIL.n78 2.71565
R770 VTAIL.n180 VTAIL.n179 2.71565
R771 VTAIL.n198 VTAIL.n150 2.71565
R772 VTAIL.n482 VTAIL.n434 2.71565
R773 VTAIL.n465 VTAIL.n464 2.71565
R774 VTAIL.n410 VTAIL.n362 2.71565
R775 VTAIL.n393 VTAIL.n392 2.71565
R776 VTAIL.n340 VTAIL.n292 2.71565
R777 VTAIL.n323 VTAIL.n322 2.71565
R778 VTAIL.n268 VTAIL.n220 2.71565
R779 VTAIL.n251 VTAIL.n250 2.71565
R780 VTAIL.n0 VTAIL.t15 2.53599
R781 VTAIL.n0 VTAIL.t2 2.53599
R782 VTAIL.n142 VTAIL.t7 2.53599
R783 VTAIL.n142 VTAIL.t12 2.53599
R784 VTAIL.n426 VTAIL.t13 2.53599
R785 VTAIL.n426 VTAIL.t14 2.53599
R786 VTAIL.n284 VTAIL.t4 2.53599
R787 VTAIL.n284 VTAIL.t3 2.53599
R788 VTAIL.n523 VTAIL.n519 2.41282
R789 VTAIL.n27 VTAIL.n23 2.41282
R790 VTAIL.n97 VTAIL.n93 2.41282
R791 VTAIL.n169 VTAIL.n165 2.41282
R792 VTAIL.n454 VTAIL.n450 2.41282
R793 VTAIL.n382 VTAIL.n378 2.41282
R794 VTAIL.n312 VTAIL.n308 2.41282
R795 VTAIL.n240 VTAIL.n236 2.41282
R796 VTAIL.n285 VTAIL.n283 2.02636
R797 VTAIL.n355 VTAIL.n285 2.02636
R798 VTAIL.n427 VTAIL.n425 2.02636
R799 VTAIL.n497 VTAIL.n427 2.02636
R800 VTAIL.n213 VTAIL.n143 2.02636
R801 VTAIL.n143 VTAIL.n141 2.02636
R802 VTAIL.n71 VTAIL.n1 2.02636
R803 VTAIL VTAIL.n567 1.96817
R804 VTAIL.n538 VTAIL.n512 1.93989
R805 VTAIL.n551 VTAIL.n506 1.93989
R806 VTAIL.n42 VTAIL.n16 1.93989
R807 VTAIL.n55 VTAIL.n10 1.93989
R808 VTAIL.n112 VTAIL.n86 1.93989
R809 VTAIL.n125 VTAIL.n80 1.93989
R810 VTAIL.n184 VTAIL.n158 1.93989
R811 VTAIL.n197 VTAIL.n152 1.93989
R812 VTAIL.n481 VTAIL.n436 1.93989
R813 VTAIL.n468 VTAIL.n442 1.93989
R814 VTAIL.n409 VTAIL.n364 1.93989
R815 VTAIL.n396 VTAIL.n370 1.93989
R816 VTAIL.n339 VTAIL.n294 1.93989
R817 VTAIL.n326 VTAIL.n300 1.93989
R818 VTAIL.n267 VTAIL.n222 1.93989
R819 VTAIL.n254 VTAIL.n228 1.93989
R820 VTAIL.n539 VTAIL.n510 1.16414
R821 VTAIL.n548 VTAIL.n547 1.16414
R822 VTAIL.n43 VTAIL.n14 1.16414
R823 VTAIL.n52 VTAIL.n51 1.16414
R824 VTAIL.n113 VTAIL.n84 1.16414
R825 VTAIL.n122 VTAIL.n121 1.16414
R826 VTAIL.n185 VTAIL.n156 1.16414
R827 VTAIL.n194 VTAIL.n193 1.16414
R828 VTAIL.n478 VTAIL.n477 1.16414
R829 VTAIL.n469 VTAIL.n440 1.16414
R830 VTAIL.n406 VTAIL.n405 1.16414
R831 VTAIL.n397 VTAIL.n368 1.16414
R832 VTAIL.n336 VTAIL.n335 1.16414
R833 VTAIL.n327 VTAIL.n298 1.16414
R834 VTAIL.n264 VTAIL.n263 1.16414
R835 VTAIL.n255 VTAIL.n226 1.16414
R836 VTAIL.n425 VTAIL.n355 0.470328
R837 VTAIL.n141 VTAIL.n71 0.470328
R838 VTAIL.n543 VTAIL.n542 0.388379
R839 VTAIL.n544 VTAIL.n508 0.388379
R840 VTAIL.n47 VTAIL.n46 0.388379
R841 VTAIL.n48 VTAIL.n12 0.388379
R842 VTAIL.n117 VTAIL.n116 0.388379
R843 VTAIL.n118 VTAIL.n82 0.388379
R844 VTAIL.n189 VTAIL.n188 0.388379
R845 VTAIL.n190 VTAIL.n154 0.388379
R846 VTAIL.n474 VTAIL.n438 0.388379
R847 VTAIL.n473 VTAIL.n472 0.388379
R848 VTAIL.n402 VTAIL.n366 0.388379
R849 VTAIL.n401 VTAIL.n400 0.388379
R850 VTAIL.n332 VTAIL.n296 0.388379
R851 VTAIL.n331 VTAIL.n330 0.388379
R852 VTAIL.n260 VTAIL.n224 0.388379
R853 VTAIL.n259 VTAIL.n258 0.388379
R854 VTAIL.n524 VTAIL.n523 0.155672
R855 VTAIL.n524 VTAIL.n515 0.155672
R856 VTAIL.n531 VTAIL.n515 0.155672
R857 VTAIL.n532 VTAIL.n531 0.155672
R858 VTAIL.n532 VTAIL.n511 0.155672
R859 VTAIL.n540 VTAIL.n511 0.155672
R860 VTAIL.n541 VTAIL.n540 0.155672
R861 VTAIL.n541 VTAIL.n507 0.155672
R862 VTAIL.n549 VTAIL.n507 0.155672
R863 VTAIL.n550 VTAIL.n549 0.155672
R864 VTAIL.n550 VTAIL.n503 0.155672
R865 VTAIL.n557 VTAIL.n503 0.155672
R866 VTAIL.n558 VTAIL.n557 0.155672
R867 VTAIL.n558 VTAIL.n499 0.155672
R868 VTAIL.n565 VTAIL.n499 0.155672
R869 VTAIL.n28 VTAIL.n27 0.155672
R870 VTAIL.n28 VTAIL.n19 0.155672
R871 VTAIL.n35 VTAIL.n19 0.155672
R872 VTAIL.n36 VTAIL.n35 0.155672
R873 VTAIL.n36 VTAIL.n15 0.155672
R874 VTAIL.n44 VTAIL.n15 0.155672
R875 VTAIL.n45 VTAIL.n44 0.155672
R876 VTAIL.n45 VTAIL.n11 0.155672
R877 VTAIL.n53 VTAIL.n11 0.155672
R878 VTAIL.n54 VTAIL.n53 0.155672
R879 VTAIL.n54 VTAIL.n7 0.155672
R880 VTAIL.n61 VTAIL.n7 0.155672
R881 VTAIL.n62 VTAIL.n61 0.155672
R882 VTAIL.n62 VTAIL.n3 0.155672
R883 VTAIL.n69 VTAIL.n3 0.155672
R884 VTAIL.n98 VTAIL.n97 0.155672
R885 VTAIL.n98 VTAIL.n89 0.155672
R886 VTAIL.n105 VTAIL.n89 0.155672
R887 VTAIL.n106 VTAIL.n105 0.155672
R888 VTAIL.n106 VTAIL.n85 0.155672
R889 VTAIL.n114 VTAIL.n85 0.155672
R890 VTAIL.n115 VTAIL.n114 0.155672
R891 VTAIL.n115 VTAIL.n81 0.155672
R892 VTAIL.n123 VTAIL.n81 0.155672
R893 VTAIL.n124 VTAIL.n123 0.155672
R894 VTAIL.n124 VTAIL.n77 0.155672
R895 VTAIL.n131 VTAIL.n77 0.155672
R896 VTAIL.n132 VTAIL.n131 0.155672
R897 VTAIL.n132 VTAIL.n73 0.155672
R898 VTAIL.n139 VTAIL.n73 0.155672
R899 VTAIL.n170 VTAIL.n169 0.155672
R900 VTAIL.n170 VTAIL.n161 0.155672
R901 VTAIL.n177 VTAIL.n161 0.155672
R902 VTAIL.n178 VTAIL.n177 0.155672
R903 VTAIL.n178 VTAIL.n157 0.155672
R904 VTAIL.n186 VTAIL.n157 0.155672
R905 VTAIL.n187 VTAIL.n186 0.155672
R906 VTAIL.n187 VTAIL.n153 0.155672
R907 VTAIL.n195 VTAIL.n153 0.155672
R908 VTAIL.n196 VTAIL.n195 0.155672
R909 VTAIL.n196 VTAIL.n149 0.155672
R910 VTAIL.n203 VTAIL.n149 0.155672
R911 VTAIL.n204 VTAIL.n203 0.155672
R912 VTAIL.n204 VTAIL.n145 0.155672
R913 VTAIL.n211 VTAIL.n145 0.155672
R914 VTAIL.n495 VTAIL.n429 0.155672
R915 VTAIL.n488 VTAIL.n429 0.155672
R916 VTAIL.n488 VTAIL.n487 0.155672
R917 VTAIL.n487 VTAIL.n433 0.155672
R918 VTAIL.n480 VTAIL.n433 0.155672
R919 VTAIL.n480 VTAIL.n479 0.155672
R920 VTAIL.n479 VTAIL.n437 0.155672
R921 VTAIL.n471 VTAIL.n437 0.155672
R922 VTAIL.n471 VTAIL.n470 0.155672
R923 VTAIL.n470 VTAIL.n441 0.155672
R924 VTAIL.n463 VTAIL.n441 0.155672
R925 VTAIL.n463 VTAIL.n462 0.155672
R926 VTAIL.n462 VTAIL.n446 0.155672
R927 VTAIL.n455 VTAIL.n446 0.155672
R928 VTAIL.n455 VTAIL.n454 0.155672
R929 VTAIL.n423 VTAIL.n357 0.155672
R930 VTAIL.n416 VTAIL.n357 0.155672
R931 VTAIL.n416 VTAIL.n415 0.155672
R932 VTAIL.n415 VTAIL.n361 0.155672
R933 VTAIL.n408 VTAIL.n361 0.155672
R934 VTAIL.n408 VTAIL.n407 0.155672
R935 VTAIL.n407 VTAIL.n365 0.155672
R936 VTAIL.n399 VTAIL.n365 0.155672
R937 VTAIL.n399 VTAIL.n398 0.155672
R938 VTAIL.n398 VTAIL.n369 0.155672
R939 VTAIL.n391 VTAIL.n369 0.155672
R940 VTAIL.n391 VTAIL.n390 0.155672
R941 VTAIL.n390 VTAIL.n374 0.155672
R942 VTAIL.n383 VTAIL.n374 0.155672
R943 VTAIL.n383 VTAIL.n382 0.155672
R944 VTAIL.n353 VTAIL.n287 0.155672
R945 VTAIL.n346 VTAIL.n287 0.155672
R946 VTAIL.n346 VTAIL.n345 0.155672
R947 VTAIL.n345 VTAIL.n291 0.155672
R948 VTAIL.n338 VTAIL.n291 0.155672
R949 VTAIL.n338 VTAIL.n337 0.155672
R950 VTAIL.n337 VTAIL.n295 0.155672
R951 VTAIL.n329 VTAIL.n295 0.155672
R952 VTAIL.n329 VTAIL.n328 0.155672
R953 VTAIL.n328 VTAIL.n299 0.155672
R954 VTAIL.n321 VTAIL.n299 0.155672
R955 VTAIL.n321 VTAIL.n320 0.155672
R956 VTAIL.n320 VTAIL.n304 0.155672
R957 VTAIL.n313 VTAIL.n304 0.155672
R958 VTAIL.n313 VTAIL.n312 0.155672
R959 VTAIL.n281 VTAIL.n215 0.155672
R960 VTAIL.n274 VTAIL.n215 0.155672
R961 VTAIL.n274 VTAIL.n273 0.155672
R962 VTAIL.n273 VTAIL.n219 0.155672
R963 VTAIL.n266 VTAIL.n219 0.155672
R964 VTAIL.n266 VTAIL.n265 0.155672
R965 VTAIL.n265 VTAIL.n223 0.155672
R966 VTAIL.n257 VTAIL.n223 0.155672
R967 VTAIL.n257 VTAIL.n256 0.155672
R968 VTAIL.n256 VTAIL.n227 0.155672
R969 VTAIL.n249 VTAIL.n227 0.155672
R970 VTAIL.n249 VTAIL.n248 0.155672
R971 VTAIL.n248 VTAIL.n232 0.155672
R972 VTAIL.n241 VTAIL.n232 0.155672
R973 VTAIL.n241 VTAIL.n240 0.155672
R974 VTAIL VTAIL.n1 0.0586897
R975 VN.n6 VN.t3 184.838
R976 VN.n31 VN.t2 184.838
R977 VN.n24 VN.n23 184.427
R978 VN.n49 VN.n48 184.427
R979 VN.n47 VN.n25 161.3
R980 VN.n46 VN.n45 161.3
R981 VN.n44 VN.n26 161.3
R982 VN.n43 VN.n42 161.3
R983 VN.n41 VN.n27 161.3
R984 VN.n39 VN.n38 161.3
R985 VN.n37 VN.n28 161.3
R986 VN.n36 VN.n35 161.3
R987 VN.n34 VN.n29 161.3
R988 VN.n33 VN.n32 161.3
R989 VN.n22 VN.n0 161.3
R990 VN.n21 VN.n20 161.3
R991 VN.n19 VN.n1 161.3
R992 VN.n18 VN.n17 161.3
R993 VN.n16 VN.n2 161.3
R994 VN.n14 VN.n13 161.3
R995 VN.n12 VN.n3 161.3
R996 VN.n11 VN.n10 161.3
R997 VN.n9 VN.n4 161.3
R998 VN.n8 VN.n7 161.3
R999 VN.n5 VN.t7 152.952
R1000 VN.n15 VN.t6 152.952
R1001 VN.n23 VN.t1 152.952
R1002 VN.n30 VN.t4 152.952
R1003 VN.n40 VN.t5 152.952
R1004 VN.n48 VN.t0 152.952
R1005 VN.n6 VN.n5 61.6806
R1006 VN.n31 VN.n30 61.6806
R1007 VN.n17 VN.n1 55.0167
R1008 VN.n42 VN.n26 55.0167
R1009 VN VN.n49 49.1009
R1010 VN.n10 VN.n9 40.4106
R1011 VN.n10 VN.n3 40.4106
R1012 VN.n35 VN.n34 40.4106
R1013 VN.n35 VN.n28 40.4106
R1014 VN.n21 VN.n1 25.8045
R1015 VN.n46 VN.n26 25.8045
R1016 VN.n9 VN.n8 24.3439
R1017 VN.n14 VN.n3 24.3439
R1018 VN.n17 VN.n16 24.3439
R1019 VN.n22 VN.n21 24.3439
R1020 VN.n34 VN.n33 24.3439
R1021 VN.n42 VN.n41 24.3439
R1022 VN.n39 VN.n28 24.3439
R1023 VN.n47 VN.n46 24.3439
R1024 VN.n16 VN.n15 15.8237
R1025 VN.n41 VN.n40 15.8237
R1026 VN.n32 VN.n31 12.5995
R1027 VN.n7 VN.n6 12.5995
R1028 VN.n8 VN.n5 8.5207
R1029 VN.n15 VN.n14 8.5207
R1030 VN.n33 VN.n30 8.5207
R1031 VN.n40 VN.n39 8.5207
R1032 VN.n23 VN.n22 1.21767
R1033 VN.n48 VN.n47 1.21767
R1034 VN.n49 VN.n25 0.189894
R1035 VN.n45 VN.n25 0.189894
R1036 VN.n45 VN.n44 0.189894
R1037 VN.n44 VN.n43 0.189894
R1038 VN.n43 VN.n27 0.189894
R1039 VN.n38 VN.n27 0.189894
R1040 VN.n38 VN.n37 0.189894
R1041 VN.n37 VN.n36 0.189894
R1042 VN.n36 VN.n29 0.189894
R1043 VN.n32 VN.n29 0.189894
R1044 VN.n7 VN.n4 0.189894
R1045 VN.n11 VN.n4 0.189894
R1046 VN.n12 VN.n11 0.189894
R1047 VN.n13 VN.n12 0.189894
R1048 VN.n13 VN.n2 0.189894
R1049 VN.n18 VN.n2 0.189894
R1050 VN.n19 VN.n18 0.189894
R1051 VN.n20 VN.n19 0.189894
R1052 VN.n20 VN.n0 0.189894
R1053 VN.n24 VN.n0 0.189894
R1054 VN VN.n24 0.0516364
R1055 VDD2.n2 VDD2.n1 73.5811
R1056 VDD2.n2 VDD2.n0 73.5811
R1057 VDD2 VDD2.n5 73.578
R1058 VDD2.n4 VDD2.n3 72.6235
R1059 VDD2.n4 VDD2.n2 43.8834
R1060 VDD2.n5 VDD2.t3 2.53599
R1061 VDD2.n5 VDD2.t5 2.53599
R1062 VDD2.n3 VDD2.t7 2.53599
R1063 VDD2.n3 VDD2.t2 2.53599
R1064 VDD2.n1 VDD2.t1 2.53599
R1065 VDD2.n1 VDD2.t6 2.53599
R1066 VDD2.n0 VDD2.t4 2.53599
R1067 VDD2.n0 VDD2.t0 2.53599
R1068 VDD2 VDD2.n4 1.07162
R1069 B.n403 B.n402 585
R1070 B.n401 B.n120 585
R1071 B.n400 B.n399 585
R1072 B.n398 B.n121 585
R1073 B.n397 B.n396 585
R1074 B.n395 B.n122 585
R1075 B.n394 B.n393 585
R1076 B.n392 B.n123 585
R1077 B.n391 B.n390 585
R1078 B.n389 B.n124 585
R1079 B.n388 B.n387 585
R1080 B.n386 B.n125 585
R1081 B.n385 B.n384 585
R1082 B.n383 B.n126 585
R1083 B.n382 B.n381 585
R1084 B.n380 B.n127 585
R1085 B.n379 B.n378 585
R1086 B.n377 B.n128 585
R1087 B.n376 B.n375 585
R1088 B.n374 B.n129 585
R1089 B.n373 B.n372 585
R1090 B.n371 B.n130 585
R1091 B.n370 B.n369 585
R1092 B.n368 B.n131 585
R1093 B.n367 B.n366 585
R1094 B.n365 B.n132 585
R1095 B.n364 B.n363 585
R1096 B.n362 B.n133 585
R1097 B.n361 B.n360 585
R1098 B.n359 B.n134 585
R1099 B.n358 B.n357 585
R1100 B.n356 B.n135 585
R1101 B.n355 B.n354 585
R1102 B.n353 B.n136 585
R1103 B.n352 B.n351 585
R1104 B.n350 B.n137 585
R1105 B.n349 B.n348 585
R1106 B.n347 B.n138 585
R1107 B.n346 B.n345 585
R1108 B.n344 B.n139 585
R1109 B.n343 B.n342 585
R1110 B.n341 B.n140 585
R1111 B.n340 B.n339 585
R1112 B.n338 B.n141 585
R1113 B.n336 B.n335 585
R1114 B.n334 B.n144 585
R1115 B.n333 B.n332 585
R1116 B.n331 B.n145 585
R1117 B.n330 B.n329 585
R1118 B.n328 B.n146 585
R1119 B.n327 B.n326 585
R1120 B.n325 B.n147 585
R1121 B.n324 B.n323 585
R1122 B.n322 B.n148 585
R1123 B.n321 B.n320 585
R1124 B.n316 B.n149 585
R1125 B.n315 B.n314 585
R1126 B.n313 B.n150 585
R1127 B.n312 B.n311 585
R1128 B.n310 B.n151 585
R1129 B.n309 B.n308 585
R1130 B.n307 B.n152 585
R1131 B.n306 B.n305 585
R1132 B.n304 B.n153 585
R1133 B.n303 B.n302 585
R1134 B.n301 B.n154 585
R1135 B.n300 B.n299 585
R1136 B.n298 B.n155 585
R1137 B.n297 B.n296 585
R1138 B.n295 B.n156 585
R1139 B.n294 B.n293 585
R1140 B.n292 B.n157 585
R1141 B.n291 B.n290 585
R1142 B.n289 B.n158 585
R1143 B.n288 B.n287 585
R1144 B.n286 B.n159 585
R1145 B.n285 B.n284 585
R1146 B.n283 B.n160 585
R1147 B.n282 B.n281 585
R1148 B.n280 B.n161 585
R1149 B.n279 B.n278 585
R1150 B.n277 B.n162 585
R1151 B.n276 B.n275 585
R1152 B.n274 B.n163 585
R1153 B.n273 B.n272 585
R1154 B.n271 B.n164 585
R1155 B.n270 B.n269 585
R1156 B.n268 B.n165 585
R1157 B.n267 B.n266 585
R1158 B.n265 B.n166 585
R1159 B.n264 B.n263 585
R1160 B.n262 B.n167 585
R1161 B.n261 B.n260 585
R1162 B.n259 B.n168 585
R1163 B.n258 B.n257 585
R1164 B.n256 B.n169 585
R1165 B.n255 B.n254 585
R1166 B.n253 B.n170 585
R1167 B.n404 B.n119 585
R1168 B.n406 B.n405 585
R1169 B.n407 B.n118 585
R1170 B.n409 B.n408 585
R1171 B.n410 B.n117 585
R1172 B.n412 B.n411 585
R1173 B.n413 B.n116 585
R1174 B.n415 B.n414 585
R1175 B.n416 B.n115 585
R1176 B.n418 B.n417 585
R1177 B.n419 B.n114 585
R1178 B.n421 B.n420 585
R1179 B.n422 B.n113 585
R1180 B.n424 B.n423 585
R1181 B.n425 B.n112 585
R1182 B.n427 B.n426 585
R1183 B.n428 B.n111 585
R1184 B.n430 B.n429 585
R1185 B.n431 B.n110 585
R1186 B.n433 B.n432 585
R1187 B.n434 B.n109 585
R1188 B.n436 B.n435 585
R1189 B.n437 B.n108 585
R1190 B.n439 B.n438 585
R1191 B.n440 B.n107 585
R1192 B.n442 B.n441 585
R1193 B.n443 B.n106 585
R1194 B.n445 B.n444 585
R1195 B.n446 B.n105 585
R1196 B.n448 B.n447 585
R1197 B.n449 B.n104 585
R1198 B.n451 B.n450 585
R1199 B.n452 B.n103 585
R1200 B.n454 B.n453 585
R1201 B.n455 B.n102 585
R1202 B.n457 B.n456 585
R1203 B.n458 B.n101 585
R1204 B.n460 B.n459 585
R1205 B.n461 B.n100 585
R1206 B.n463 B.n462 585
R1207 B.n464 B.n99 585
R1208 B.n466 B.n465 585
R1209 B.n467 B.n98 585
R1210 B.n469 B.n468 585
R1211 B.n470 B.n97 585
R1212 B.n472 B.n471 585
R1213 B.n473 B.n96 585
R1214 B.n475 B.n474 585
R1215 B.n476 B.n95 585
R1216 B.n478 B.n477 585
R1217 B.n479 B.n94 585
R1218 B.n481 B.n480 585
R1219 B.n482 B.n93 585
R1220 B.n484 B.n483 585
R1221 B.n485 B.n92 585
R1222 B.n487 B.n486 585
R1223 B.n488 B.n91 585
R1224 B.n490 B.n489 585
R1225 B.n491 B.n90 585
R1226 B.n493 B.n492 585
R1227 B.n494 B.n89 585
R1228 B.n496 B.n495 585
R1229 B.n497 B.n88 585
R1230 B.n499 B.n498 585
R1231 B.n500 B.n87 585
R1232 B.n502 B.n501 585
R1233 B.n503 B.n86 585
R1234 B.n505 B.n504 585
R1235 B.n506 B.n85 585
R1236 B.n508 B.n507 585
R1237 B.n509 B.n84 585
R1238 B.n511 B.n510 585
R1239 B.n512 B.n83 585
R1240 B.n514 B.n513 585
R1241 B.n515 B.n82 585
R1242 B.n517 B.n516 585
R1243 B.n518 B.n81 585
R1244 B.n520 B.n519 585
R1245 B.n521 B.n80 585
R1246 B.n523 B.n522 585
R1247 B.n524 B.n79 585
R1248 B.n526 B.n525 585
R1249 B.n527 B.n78 585
R1250 B.n529 B.n528 585
R1251 B.n530 B.n77 585
R1252 B.n532 B.n531 585
R1253 B.n680 B.n23 585
R1254 B.n679 B.n678 585
R1255 B.n677 B.n24 585
R1256 B.n676 B.n675 585
R1257 B.n674 B.n25 585
R1258 B.n673 B.n672 585
R1259 B.n671 B.n26 585
R1260 B.n670 B.n669 585
R1261 B.n668 B.n27 585
R1262 B.n667 B.n666 585
R1263 B.n665 B.n28 585
R1264 B.n664 B.n663 585
R1265 B.n662 B.n29 585
R1266 B.n661 B.n660 585
R1267 B.n659 B.n30 585
R1268 B.n658 B.n657 585
R1269 B.n656 B.n31 585
R1270 B.n655 B.n654 585
R1271 B.n653 B.n32 585
R1272 B.n652 B.n651 585
R1273 B.n650 B.n33 585
R1274 B.n649 B.n648 585
R1275 B.n647 B.n34 585
R1276 B.n646 B.n645 585
R1277 B.n644 B.n35 585
R1278 B.n643 B.n642 585
R1279 B.n641 B.n36 585
R1280 B.n640 B.n639 585
R1281 B.n638 B.n37 585
R1282 B.n637 B.n636 585
R1283 B.n635 B.n38 585
R1284 B.n634 B.n633 585
R1285 B.n632 B.n39 585
R1286 B.n631 B.n630 585
R1287 B.n629 B.n40 585
R1288 B.n628 B.n627 585
R1289 B.n626 B.n41 585
R1290 B.n625 B.n624 585
R1291 B.n623 B.n42 585
R1292 B.n622 B.n621 585
R1293 B.n620 B.n43 585
R1294 B.n619 B.n618 585
R1295 B.n617 B.n44 585
R1296 B.n616 B.n615 585
R1297 B.n613 B.n45 585
R1298 B.n612 B.n611 585
R1299 B.n610 B.n48 585
R1300 B.n609 B.n608 585
R1301 B.n607 B.n49 585
R1302 B.n606 B.n605 585
R1303 B.n604 B.n50 585
R1304 B.n603 B.n602 585
R1305 B.n601 B.n51 585
R1306 B.n600 B.n599 585
R1307 B.n598 B.n597 585
R1308 B.n596 B.n55 585
R1309 B.n595 B.n594 585
R1310 B.n593 B.n56 585
R1311 B.n592 B.n591 585
R1312 B.n590 B.n57 585
R1313 B.n589 B.n588 585
R1314 B.n587 B.n58 585
R1315 B.n586 B.n585 585
R1316 B.n584 B.n59 585
R1317 B.n583 B.n582 585
R1318 B.n581 B.n60 585
R1319 B.n580 B.n579 585
R1320 B.n578 B.n61 585
R1321 B.n577 B.n576 585
R1322 B.n575 B.n62 585
R1323 B.n574 B.n573 585
R1324 B.n572 B.n63 585
R1325 B.n571 B.n570 585
R1326 B.n569 B.n64 585
R1327 B.n568 B.n567 585
R1328 B.n566 B.n65 585
R1329 B.n565 B.n564 585
R1330 B.n563 B.n66 585
R1331 B.n562 B.n561 585
R1332 B.n560 B.n67 585
R1333 B.n559 B.n558 585
R1334 B.n557 B.n68 585
R1335 B.n556 B.n555 585
R1336 B.n554 B.n69 585
R1337 B.n553 B.n552 585
R1338 B.n551 B.n70 585
R1339 B.n550 B.n549 585
R1340 B.n548 B.n71 585
R1341 B.n547 B.n546 585
R1342 B.n545 B.n72 585
R1343 B.n544 B.n543 585
R1344 B.n542 B.n73 585
R1345 B.n541 B.n540 585
R1346 B.n539 B.n74 585
R1347 B.n538 B.n537 585
R1348 B.n536 B.n75 585
R1349 B.n535 B.n534 585
R1350 B.n533 B.n76 585
R1351 B.n682 B.n681 585
R1352 B.n683 B.n22 585
R1353 B.n685 B.n684 585
R1354 B.n686 B.n21 585
R1355 B.n688 B.n687 585
R1356 B.n689 B.n20 585
R1357 B.n691 B.n690 585
R1358 B.n692 B.n19 585
R1359 B.n694 B.n693 585
R1360 B.n695 B.n18 585
R1361 B.n697 B.n696 585
R1362 B.n698 B.n17 585
R1363 B.n700 B.n699 585
R1364 B.n701 B.n16 585
R1365 B.n703 B.n702 585
R1366 B.n704 B.n15 585
R1367 B.n706 B.n705 585
R1368 B.n707 B.n14 585
R1369 B.n709 B.n708 585
R1370 B.n710 B.n13 585
R1371 B.n712 B.n711 585
R1372 B.n713 B.n12 585
R1373 B.n715 B.n714 585
R1374 B.n716 B.n11 585
R1375 B.n718 B.n717 585
R1376 B.n719 B.n10 585
R1377 B.n721 B.n720 585
R1378 B.n722 B.n9 585
R1379 B.n724 B.n723 585
R1380 B.n725 B.n8 585
R1381 B.n727 B.n726 585
R1382 B.n728 B.n7 585
R1383 B.n730 B.n729 585
R1384 B.n731 B.n6 585
R1385 B.n733 B.n732 585
R1386 B.n734 B.n5 585
R1387 B.n736 B.n735 585
R1388 B.n737 B.n4 585
R1389 B.n739 B.n738 585
R1390 B.n740 B.n3 585
R1391 B.n742 B.n741 585
R1392 B.n743 B.n0 585
R1393 B.n2 B.n1 585
R1394 B.n192 B.n191 585
R1395 B.n193 B.n190 585
R1396 B.n195 B.n194 585
R1397 B.n196 B.n189 585
R1398 B.n198 B.n197 585
R1399 B.n199 B.n188 585
R1400 B.n201 B.n200 585
R1401 B.n202 B.n187 585
R1402 B.n204 B.n203 585
R1403 B.n205 B.n186 585
R1404 B.n207 B.n206 585
R1405 B.n208 B.n185 585
R1406 B.n210 B.n209 585
R1407 B.n211 B.n184 585
R1408 B.n213 B.n212 585
R1409 B.n214 B.n183 585
R1410 B.n216 B.n215 585
R1411 B.n217 B.n182 585
R1412 B.n219 B.n218 585
R1413 B.n220 B.n181 585
R1414 B.n222 B.n221 585
R1415 B.n223 B.n180 585
R1416 B.n225 B.n224 585
R1417 B.n226 B.n179 585
R1418 B.n228 B.n227 585
R1419 B.n229 B.n178 585
R1420 B.n231 B.n230 585
R1421 B.n232 B.n177 585
R1422 B.n234 B.n233 585
R1423 B.n235 B.n176 585
R1424 B.n237 B.n236 585
R1425 B.n238 B.n175 585
R1426 B.n240 B.n239 585
R1427 B.n241 B.n174 585
R1428 B.n243 B.n242 585
R1429 B.n244 B.n173 585
R1430 B.n246 B.n245 585
R1431 B.n247 B.n172 585
R1432 B.n249 B.n248 585
R1433 B.n250 B.n171 585
R1434 B.n252 B.n251 585
R1435 B.n253 B.n252 497.305
R1436 B.n402 B.n119 497.305
R1437 B.n533 B.n532 497.305
R1438 B.n682 B.n23 497.305
R1439 B.n142 B.t10 436.067
R1440 B.n52 B.t8 436.067
R1441 B.n317 B.t1 436.067
R1442 B.n46 B.t5 436.067
R1443 B.n143 B.t11 390.491
R1444 B.n53 B.t7 390.491
R1445 B.n318 B.t2 390.491
R1446 B.n47 B.t4 390.491
R1447 B.n317 B.t0 359.916
R1448 B.n142 B.t9 359.916
R1449 B.n52 B.t6 359.916
R1450 B.n46 B.t3 359.916
R1451 B.n745 B.n744 256.663
R1452 B.n744 B.n743 235.042
R1453 B.n744 B.n2 235.042
R1454 B.n254 B.n253 163.367
R1455 B.n254 B.n169 163.367
R1456 B.n258 B.n169 163.367
R1457 B.n259 B.n258 163.367
R1458 B.n260 B.n259 163.367
R1459 B.n260 B.n167 163.367
R1460 B.n264 B.n167 163.367
R1461 B.n265 B.n264 163.367
R1462 B.n266 B.n265 163.367
R1463 B.n266 B.n165 163.367
R1464 B.n270 B.n165 163.367
R1465 B.n271 B.n270 163.367
R1466 B.n272 B.n271 163.367
R1467 B.n272 B.n163 163.367
R1468 B.n276 B.n163 163.367
R1469 B.n277 B.n276 163.367
R1470 B.n278 B.n277 163.367
R1471 B.n278 B.n161 163.367
R1472 B.n282 B.n161 163.367
R1473 B.n283 B.n282 163.367
R1474 B.n284 B.n283 163.367
R1475 B.n284 B.n159 163.367
R1476 B.n288 B.n159 163.367
R1477 B.n289 B.n288 163.367
R1478 B.n290 B.n289 163.367
R1479 B.n290 B.n157 163.367
R1480 B.n294 B.n157 163.367
R1481 B.n295 B.n294 163.367
R1482 B.n296 B.n295 163.367
R1483 B.n296 B.n155 163.367
R1484 B.n300 B.n155 163.367
R1485 B.n301 B.n300 163.367
R1486 B.n302 B.n301 163.367
R1487 B.n302 B.n153 163.367
R1488 B.n306 B.n153 163.367
R1489 B.n307 B.n306 163.367
R1490 B.n308 B.n307 163.367
R1491 B.n308 B.n151 163.367
R1492 B.n312 B.n151 163.367
R1493 B.n313 B.n312 163.367
R1494 B.n314 B.n313 163.367
R1495 B.n314 B.n149 163.367
R1496 B.n321 B.n149 163.367
R1497 B.n322 B.n321 163.367
R1498 B.n323 B.n322 163.367
R1499 B.n323 B.n147 163.367
R1500 B.n327 B.n147 163.367
R1501 B.n328 B.n327 163.367
R1502 B.n329 B.n328 163.367
R1503 B.n329 B.n145 163.367
R1504 B.n333 B.n145 163.367
R1505 B.n334 B.n333 163.367
R1506 B.n335 B.n334 163.367
R1507 B.n335 B.n141 163.367
R1508 B.n340 B.n141 163.367
R1509 B.n341 B.n340 163.367
R1510 B.n342 B.n341 163.367
R1511 B.n342 B.n139 163.367
R1512 B.n346 B.n139 163.367
R1513 B.n347 B.n346 163.367
R1514 B.n348 B.n347 163.367
R1515 B.n348 B.n137 163.367
R1516 B.n352 B.n137 163.367
R1517 B.n353 B.n352 163.367
R1518 B.n354 B.n353 163.367
R1519 B.n354 B.n135 163.367
R1520 B.n358 B.n135 163.367
R1521 B.n359 B.n358 163.367
R1522 B.n360 B.n359 163.367
R1523 B.n360 B.n133 163.367
R1524 B.n364 B.n133 163.367
R1525 B.n365 B.n364 163.367
R1526 B.n366 B.n365 163.367
R1527 B.n366 B.n131 163.367
R1528 B.n370 B.n131 163.367
R1529 B.n371 B.n370 163.367
R1530 B.n372 B.n371 163.367
R1531 B.n372 B.n129 163.367
R1532 B.n376 B.n129 163.367
R1533 B.n377 B.n376 163.367
R1534 B.n378 B.n377 163.367
R1535 B.n378 B.n127 163.367
R1536 B.n382 B.n127 163.367
R1537 B.n383 B.n382 163.367
R1538 B.n384 B.n383 163.367
R1539 B.n384 B.n125 163.367
R1540 B.n388 B.n125 163.367
R1541 B.n389 B.n388 163.367
R1542 B.n390 B.n389 163.367
R1543 B.n390 B.n123 163.367
R1544 B.n394 B.n123 163.367
R1545 B.n395 B.n394 163.367
R1546 B.n396 B.n395 163.367
R1547 B.n396 B.n121 163.367
R1548 B.n400 B.n121 163.367
R1549 B.n401 B.n400 163.367
R1550 B.n402 B.n401 163.367
R1551 B.n532 B.n77 163.367
R1552 B.n528 B.n77 163.367
R1553 B.n528 B.n527 163.367
R1554 B.n527 B.n526 163.367
R1555 B.n526 B.n79 163.367
R1556 B.n522 B.n79 163.367
R1557 B.n522 B.n521 163.367
R1558 B.n521 B.n520 163.367
R1559 B.n520 B.n81 163.367
R1560 B.n516 B.n81 163.367
R1561 B.n516 B.n515 163.367
R1562 B.n515 B.n514 163.367
R1563 B.n514 B.n83 163.367
R1564 B.n510 B.n83 163.367
R1565 B.n510 B.n509 163.367
R1566 B.n509 B.n508 163.367
R1567 B.n508 B.n85 163.367
R1568 B.n504 B.n85 163.367
R1569 B.n504 B.n503 163.367
R1570 B.n503 B.n502 163.367
R1571 B.n502 B.n87 163.367
R1572 B.n498 B.n87 163.367
R1573 B.n498 B.n497 163.367
R1574 B.n497 B.n496 163.367
R1575 B.n496 B.n89 163.367
R1576 B.n492 B.n89 163.367
R1577 B.n492 B.n491 163.367
R1578 B.n491 B.n490 163.367
R1579 B.n490 B.n91 163.367
R1580 B.n486 B.n91 163.367
R1581 B.n486 B.n485 163.367
R1582 B.n485 B.n484 163.367
R1583 B.n484 B.n93 163.367
R1584 B.n480 B.n93 163.367
R1585 B.n480 B.n479 163.367
R1586 B.n479 B.n478 163.367
R1587 B.n478 B.n95 163.367
R1588 B.n474 B.n95 163.367
R1589 B.n474 B.n473 163.367
R1590 B.n473 B.n472 163.367
R1591 B.n472 B.n97 163.367
R1592 B.n468 B.n97 163.367
R1593 B.n468 B.n467 163.367
R1594 B.n467 B.n466 163.367
R1595 B.n466 B.n99 163.367
R1596 B.n462 B.n99 163.367
R1597 B.n462 B.n461 163.367
R1598 B.n461 B.n460 163.367
R1599 B.n460 B.n101 163.367
R1600 B.n456 B.n101 163.367
R1601 B.n456 B.n455 163.367
R1602 B.n455 B.n454 163.367
R1603 B.n454 B.n103 163.367
R1604 B.n450 B.n103 163.367
R1605 B.n450 B.n449 163.367
R1606 B.n449 B.n448 163.367
R1607 B.n448 B.n105 163.367
R1608 B.n444 B.n105 163.367
R1609 B.n444 B.n443 163.367
R1610 B.n443 B.n442 163.367
R1611 B.n442 B.n107 163.367
R1612 B.n438 B.n107 163.367
R1613 B.n438 B.n437 163.367
R1614 B.n437 B.n436 163.367
R1615 B.n436 B.n109 163.367
R1616 B.n432 B.n109 163.367
R1617 B.n432 B.n431 163.367
R1618 B.n431 B.n430 163.367
R1619 B.n430 B.n111 163.367
R1620 B.n426 B.n111 163.367
R1621 B.n426 B.n425 163.367
R1622 B.n425 B.n424 163.367
R1623 B.n424 B.n113 163.367
R1624 B.n420 B.n113 163.367
R1625 B.n420 B.n419 163.367
R1626 B.n419 B.n418 163.367
R1627 B.n418 B.n115 163.367
R1628 B.n414 B.n115 163.367
R1629 B.n414 B.n413 163.367
R1630 B.n413 B.n412 163.367
R1631 B.n412 B.n117 163.367
R1632 B.n408 B.n117 163.367
R1633 B.n408 B.n407 163.367
R1634 B.n407 B.n406 163.367
R1635 B.n406 B.n119 163.367
R1636 B.n678 B.n23 163.367
R1637 B.n678 B.n677 163.367
R1638 B.n677 B.n676 163.367
R1639 B.n676 B.n25 163.367
R1640 B.n672 B.n25 163.367
R1641 B.n672 B.n671 163.367
R1642 B.n671 B.n670 163.367
R1643 B.n670 B.n27 163.367
R1644 B.n666 B.n27 163.367
R1645 B.n666 B.n665 163.367
R1646 B.n665 B.n664 163.367
R1647 B.n664 B.n29 163.367
R1648 B.n660 B.n29 163.367
R1649 B.n660 B.n659 163.367
R1650 B.n659 B.n658 163.367
R1651 B.n658 B.n31 163.367
R1652 B.n654 B.n31 163.367
R1653 B.n654 B.n653 163.367
R1654 B.n653 B.n652 163.367
R1655 B.n652 B.n33 163.367
R1656 B.n648 B.n33 163.367
R1657 B.n648 B.n647 163.367
R1658 B.n647 B.n646 163.367
R1659 B.n646 B.n35 163.367
R1660 B.n642 B.n35 163.367
R1661 B.n642 B.n641 163.367
R1662 B.n641 B.n640 163.367
R1663 B.n640 B.n37 163.367
R1664 B.n636 B.n37 163.367
R1665 B.n636 B.n635 163.367
R1666 B.n635 B.n634 163.367
R1667 B.n634 B.n39 163.367
R1668 B.n630 B.n39 163.367
R1669 B.n630 B.n629 163.367
R1670 B.n629 B.n628 163.367
R1671 B.n628 B.n41 163.367
R1672 B.n624 B.n41 163.367
R1673 B.n624 B.n623 163.367
R1674 B.n623 B.n622 163.367
R1675 B.n622 B.n43 163.367
R1676 B.n618 B.n43 163.367
R1677 B.n618 B.n617 163.367
R1678 B.n617 B.n616 163.367
R1679 B.n616 B.n45 163.367
R1680 B.n611 B.n45 163.367
R1681 B.n611 B.n610 163.367
R1682 B.n610 B.n609 163.367
R1683 B.n609 B.n49 163.367
R1684 B.n605 B.n49 163.367
R1685 B.n605 B.n604 163.367
R1686 B.n604 B.n603 163.367
R1687 B.n603 B.n51 163.367
R1688 B.n599 B.n51 163.367
R1689 B.n599 B.n598 163.367
R1690 B.n598 B.n55 163.367
R1691 B.n594 B.n55 163.367
R1692 B.n594 B.n593 163.367
R1693 B.n593 B.n592 163.367
R1694 B.n592 B.n57 163.367
R1695 B.n588 B.n57 163.367
R1696 B.n588 B.n587 163.367
R1697 B.n587 B.n586 163.367
R1698 B.n586 B.n59 163.367
R1699 B.n582 B.n59 163.367
R1700 B.n582 B.n581 163.367
R1701 B.n581 B.n580 163.367
R1702 B.n580 B.n61 163.367
R1703 B.n576 B.n61 163.367
R1704 B.n576 B.n575 163.367
R1705 B.n575 B.n574 163.367
R1706 B.n574 B.n63 163.367
R1707 B.n570 B.n63 163.367
R1708 B.n570 B.n569 163.367
R1709 B.n569 B.n568 163.367
R1710 B.n568 B.n65 163.367
R1711 B.n564 B.n65 163.367
R1712 B.n564 B.n563 163.367
R1713 B.n563 B.n562 163.367
R1714 B.n562 B.n67 163.367
R1715 B.n558 B.n67 163.367
R1716 B.n558 B.n557 163.367
R1717 B.n557 B.n556 163.367
R1718 B.n556 B.n69 163.367
R1719 B.n552 B.n69 163.367
R1720 B.n552 B.n551 163.367
R1721 B.n551 B.n550 163.367
R1722 B.n550 B.n71 163.367
R1723 B.n546 B.n71 163.367
R1724 B.n546 B.n545 163.367
R1725 B.n545 B.n544 163.367
R1726 B.n544 B.n73 163.367
R1727 B.n540 B.n73 163.367
R1728 B.n540 B.n539 163.367
R1729 B.n539 B.n538 163.367
R1730 B.n538 B.n75 163.367
R1731 B.n534 B.n75 163.367
R1732 B.n534 B.n533 163.367
R1733 B.n683 B.n682 163.367
R1734 B.n684 B.n683 163.367
R1735 B.n684 B.n21 163.367
R1736 B.n688 B.n21 163.367
R1737 B.n689 B.n688 163.367
R1738 B.n690 B.n689 163.367
R1739 B.n690 B.n19 163.367
R1740 B.n694 B.n19 163.367
R1741 B.n695 B.n694 163.367
R1742 B.n696 B.n695 163.367
R1743 B.n696 B.n17 163.367
R1744 B.n700 B.n17 163.367
R1745 B.n701 B.n700 163.367
R1746 B.n702 B.n701 163.367
R1747 B.n702 B.n15 163.367
R1748 B.n706 B.n15 163.367
R1749 B.n707 B.n706 163.367
R1750 B.n708 B.n707 163.367
R1751 B.n708 B.n13 163.367
R1752 B.n712 B.n13 163.367
R1753 B.n713 B.n712 163.367
R1754 B.n714 B.n713 163.367
R1755 B.n714 B.n11 163.367
R1756 B.n718 B.n11 163.367
R1757 B.n719 B.n718 163.367
R1758 B.n720 B.n719 163.367
R1759 B.n720 B.n9 163.367
R1760 B.n724 B.n9 163.367
R1761 B.n725 B.n724 163.367
R1762 B.n726 B.n725 163.367
R1763 B.n726 B.n7 163.367
R1764 B.n730 B.n7 163.367
R1765 B.n731 B.n730 163.367
R1766 B.n732 B.n731 163.367
R1767 B.n732 B.n5 163.367
R1768 B.n736 B.n5 163.367
R1769 B.n737 B.n736 163.367
R1770 B.n738 B.n737 163.367
R1771 B.n738 B.n3 163.367
R1772 B.n742 B.n3 163.367
R1773 B.n743 B.n742 163.367
R1774 B.n192 B.n2 163.367
R1775 B.n193 B.n192 163.367
R1776 B.n194 B.n193 163.367
R1777 B.n194 B.n189 163.367
R1778 B.n198 B.n189 163.367
R1779 B.n199 B.n198 163.367
R1780 B.n200 B.n199 163.367
R1781 B.n200 B.n187 163.367
R1782 B.n204 B.n187 163.367
R1783 B.n205 B.n204 163.367
R1784 B.n206 B.n205 163.367
R1785 B.n206 B.n185 163.367
R1786 B.n210 B.n185 163.367
R1787 B.n211 B.n210 163.367
R1788 B.n212 B.n211 163.367
R1789 B.n212 B.n183 163.367
R1790 B.n216 B.n183 163.367
R1791 B.n217 B.n216 163.367
R1792 B.n218 B.n217 163.367
R1793 B.n218 B.n181 163.367
R1794 B.n222 B.n181 163.367
R1795 B.n223 B.n222 163.367
R1796 B.n224 B.n223 163.367
R1797 B.n224 B.n179 163.367
R1798 B.n228 B.n179 163.367
R1799 B.n229 B.n228 163.367
R1800 B.n230 B.n229 163.367
R1801 B.n230 B.n177 163.367
R1802 B.n234 B.n177 163.367
R1803 B.n235 B.n234 163.367
R1804 B.n236 B.n235 163.367
R1805 B.n236 B.n175 163.367
R1806 B.n240 B.n175 163.367
R1807 B.n241 B.n240 163.367
R1808 B.n242 B.n241 163.367
R1809 B.n242 B.n173 163.367
R1810 B.n246 B.n173 163.367
R1811 B.n247 B.n246 163.367
R1812 B.n248 B.n247 163.367
R1813 B.n248 B.n171 163.367
R1814 B.n252 B.n171 163.367
R1815 B.n319 B.n318 59.5399
R1816 B.n337 B.n143 59.5399
R1817 B.n54 B.n53 59.5399
R1818 B.n614 B.n47 59.5399
R1819 B.n318 B.n317 45.5763
R1820 B.n143 B.n142 45.5763
R1821 B.n53 B.n52 45.5763
R1822 B.n47 B.n46 45.5763
R1823 B.n681 B.n680 32.3127
R1824 B.n531 B.n76 32.3127
R1825 B.n404 B.n403 32.3127
R1826 B.n251 B.n170 32.3127
R1827 B B.n745 18.0485
R1828 B.n681 B.n22 10.6151
R1829 B.n685 B.n22 10.6151
R1830 B.n686 B.n685 10.6151
R1831 B.n687 B.n686 10.6151
R1832 B.n687 B.n20 10.6151
R1833 B.n691 B.n20 10.6151
R1834 B.n692 B.n691 10.6151
R1835 B.n693 B.n692 10.6151
R1836 B.n693 B.n18 10.6151
R1837 B.n697 B.n18 10.6151
R1838 B.n698 B.n697 10.6151
R1839 B.n699 B.n698 10.6151
R1840 B.n699 B.n16 10.6151
R1841 B.n703 B.n16 10.6151
R1842 B.n704 B.n703 10.6151
R1843 B.n705 B.n704 10.6151
R1844 B.n705 B.n14 10.6151
R1845 B.n709 B.n14 10.6151
R1846 B.n710 B.n709 10.6151
R1847 B.n711 B.n710 10.6151
R1848 B.n711 B.n12 10.6151
R1849 B.n715 B.n12 10.6151
R1850 B.n716 B.n715 10.6151
R1851 B.n717 B.n716 10.6151
R1852 B.n717 B.n10 10.6151
R1853 B.n721 B.n10 10.6151
R1854 B.n722 B.n721 10.6151
R1855 B.n723 B.n722 10.6151
R1856 B.n723 B.n8 10.6151
R1857 B.n727 B.n8 10.6151
R1858 B.n728 B.n727 10.6151
R1859 B.n729 B.n728 10.6151
R1860 B.n729 B.n6 10.6151
R1861 B.n733 B.n6 10.6151
R1862 B.n734 B.n733 10.6151
R1863 B.n735 B.n734 10.6151
R1864 B.n735 B.n4 10.6151
R1865 B.n739 B.n4 10.6151
R1866 B.n740 B.n739 10.6151
R1867 B.n741 B.n740 10.6151
R1868 B.n741 B.n0 10.6151
R1869 B.n680 B.n679 10.6151
R1870 B.n679 B.n24 10.6151
R1871 B.n675 B.n24 10.6151
R1872 B.n675 B.n674 10.6151
R1873 B.n674 B.n673 10.6151
R1874 B.n673 B.n26 10.6151
R1875 B.n669 B.n26 10.6151
R1876 B.n669 B.n668 10.6151
R1877 B.n668 B.n667 10.6151
R1878 B.n667 B.n28 10.6151
R1879 B.n663 B.n28 10.6151
R1880 B.n663 B.n662 10.6151
R1881 B.n662 B.n661 10.6151
R1882 B.n661 B.n30 10.6151
R1883 B.n657 B.n30 10.6151
R1884 B.n657 B.n656 10.6151
R1885 B.n656 B.n655 10.6151
R1886 B.n655 B.n32 10.6151
R1887 B.n651 B.n32 10.6151
R1888 B.n651 B.n650 10.6151
R1889 B.n650 B.n649 10.6151
R1890 B.n649 B.n34 10.6151
R1891 B.n645 B.n34 10.6151
R1892 B.n645 B.n644 10.6151
R1893 B.n644 B.n643 10.6151
R1894 B.n643 B.n36 10.6151
R1895 B.n639 B.n36 10.6151
R1896 B.n639 B.n638 10.6151
R1897 B.n638 B.n637 10.6151
R1898 B.n637 B.n38 10.6151
R1899 B.n633 B.n38 10.6151
R1900 B.n633 B.n632 10.6151
R1901 B.n632 B.n631 10.6151
R1902 B.n631 B.n40 10.6151
R1903 B.n627 B.n40 10.6151
R1904 B.n627 B.n626 10.6151
R1905 B.n626 B.n625 10.6151
R1906 B.n625 B.n42 10.6151
R1907 B.n621 B.n42 10.6151
R1908 B.n621 B.n620 10.6151
R1909 B.n620 B.n619 10.6151
R1910 B.n619 B.n44 10.6151
R1911 B.n615 B.n44 10.6151
R1912 B.n613 B.n612 10.6151
R1913 B.n612 B.n48 10.6151
R1914 B.n608 B.n48 10.6151
R1915 B.n608 B.n607 10.6151
R1916 B.n607 B.n606 10.6151
R1917 B.n606 B.n50 10.6151
R1918 B.n602 B.n50 10.6151
R1919 B.n602 B.n601 10.6151
R1920 B.n601 B.n600 10.6151
R1921 B.n597 B.n596 10.6151
R1922 B.n596 B.n595 10.6151
R1923 B.n595 B.n56 10.6151
R1924 B.n591 B.n56 10.6151
R1925 B.n591 B.n590 10.6151
R1926 B.n590 B.n589 10.6151
R1927 B.n589 B.n58 10.6151
R1928 B.n585 B.n58 10.6151
R1929 B.n585 B.n584 10.6151
R1930 B.n584 B.n583 10.6151
R1931 B.n583 B.n60 10.6151
R1932 B.n579 B.n60 10.6151
R1933 B.n579 B.n578 10.6151
R1934 B.n578 B.n577 10.6151
R1935 B.n577 B.n62 10.6151
R1936 B.n573 B.n62 10.6151
R1937 B.n573 B.n572 10.6151
R1938 B.n572 B.n571 10.6151
R1939 B.n571 B.n64 10.6151
R1940 B.n567 B.n64 10.6151
R1941 B.n567 B.n566 10.6151
R1942 B.n566 B.n565 10.6151
R1943 B.n565 B.n66 10.6151
R1944 B.n561 B.n66 10.6151
R1945 B.n561 B.n560 10.6151
R1946 B.n560 B.n559 10.6151
R1947 B.n559 B.n68 10.6151
R1948 B.n555 B.n68 10.6151
R1949 B.n555 B.n554 10.6151
R1950 B.n554 B.n553 10.6151
R1951 B.n553 B.n70 10.6151
R1952 B.n549 B.n70 10.6151
R1953 B.n549 B.n548 10.6151
R1954 B.n548 B.n547 10.6151
R1955 B.n547 B.n72 10.6151
R1956 B.n543 B.n72 10.6151
R1957 B.n543 B.n542 10.6151
R1958 B.n542 B.n541 10.6151
R1959 B.n541 B.n74 10.6151
R1960 B.n537 B.n74 10.6151
R1961 B.n537 B.n536 10.6151
R1962 B.n536 B.n535 10.6151
R1963 B.n535 B.n76 10.6151
R1964 B.n531 B.n530 10.6151
R1965 B.n530 B.n529 10.6151
R1966 B.n529 B.n78 10.6151
R1967 B.n525 B.n78 10.6151
R1968 B.n525 B.n524 10.6151
R1969 B.n524 B.n523 10.6151
R1970 B.n523 B.n80 10.6151
R1971 B.n519 B.n80 10.6151
R1972 B.n519 B.n518 10.6151
R1973 B.n518 B.n517 10.6151
R1974 B.n517 B.n82 10.6151
R1975 B.n513 B.n82 10.6151
R1976 B.n513 B.n512 10.6151
R1977 B.n512 B.n511 10.6151
R1978 B.n511 B.n84 10.6151
R1979 B.n507 B.n84 10.6151
R1980 B.n507 B.n506 10.6151
R1981 B.n506 B.n505 10.6151
R1982 B.n505 B.n86 10.6151
R1983 B.n501 B.n86 10.6151
R1984 B.n501 B.n500 10.6151
R1985 B.n500 B.n499 10.6151
R1986 B.n499 B.n88 10.6151
R1987 B.n495 B.n88 10.6151
R1988 B.n495 B.n494 10.6151
R1989 B.n494 B.n493 10.6151
R1990 B.n493 B.n90 10.6151
R1991 B.n489 B.n90 10.6151
R1992 B.n489 B.n488 10.6151
R1993 B.n488 B.n487 10.6151
R1994 B.n487 B.n92 10.6151
R1995 B.n483 B.n92 10.6151
R1996 B.n483 B.n482 10.6151
R1997 B.n482 B.n481 10.6151
R1998 B.n481 B.n94 10.6151
R1999 B.n477 B.n94 10.6151
R2000 B.n477 B.n476 10.6151
R2001 B.n476 B.n475 10.6151
R2002 B.n475 B.n96 10.6151
R2003 B.n471 B.n96 10.6151
R2004 B.n471 B.n470 10.6151
R2005 B.n470 B.n469 10.6151
R2006 B.n469 B.n98 10.6151
R2007 B.n465 B.n98 10.6151
R2008 B.n465 B.n464 10.6151
R2009 B.n464 B.n463 10.6151
R2010 B.n463 B.n100 10.6151
R2011 B.n459 B.n100 10.6151
R2012 B.n459 B.n458 10.6151
R2013 B.n458 B.n457 10.6151
R2014 B.n457 B.n102 10.6151
R2015 B.n453 B.n102 10.6151
R2016 B.n453 B.n452 10.6151
R2017 B.n452 B.n451 10.6151
R2018 B.n451 B.n104 10.6151
R2019 B.n447 B.n104 10.6151
R2020 B.n447 B.n446 10.6151
R2021 B.n446 B.n445 10.6151
R2022 B.n445 B.n106 10.6151
R2023 B.n441 B.n106 10.6151
R2024 B.n441 B.n440 10.6151
R2025 B.n440 B.n439 10.6151
R2026 B.n439 B.n108 10.6151
R2027 B.n435 B.n108 10.6151
R2028 B.n435 B.n434 10.6151
R2029 B.n434 B.n433 10.6151
R2030 B.n433 B.n110 10.6151
R2031 B.n429 B.n110 10.6151
R2032 B.n429 B.n428 10.6151
R2033 B.n428 B.n427 10.6151
R2034 B.n427 B.n112 10.6151
R2035 B.n423 B.n112 10.6151
R2036 B.n423 B.n422 10.6151
R2037 B.n422 B.n421 10.6151
R2038 B.n421 B.n114 10.6151
R2039 B.n417 B.n114 10.6151
R2040 B.n417 B.n416 10.6151
R2041 B.n416 B.n415 10.6151
R2042 B.n415 B.n116 10.6151
R2043 B.n411 B.n116 10.6151
R2044 B.n411 B.n410 10.6151
R2045 B.n410 B.n409 10.6151
R2046 B.n409 B.n118 10.6151
R2047 B.n405 B.n118 10.6151
R2048 B.n405 B.n404 10.6151
R2049 B.n191 B.n1 10.6151
R2050 B.n191 B.n190 10.6151
R2051 B.n195 B.n190 10.6151
R2052 B.n196 B.n195 10.6151
R2053 B.n197 B.n196 10.6151
R2054 B.n197 B.n188 10.6151
R2055 B.n201 B.n188 10.6151
R2056 B.n202 B.n201 10.6151
R2057 B.n203 B.n202 10.6151
R2058 B.n203 B.n186 10.6151
R2059 B.n207 B.n186 10.6151
R2060 B.n208 B.n207 10.6151
R2061 B.n209 B.n208 10.6151
R2062 B.n209 B.n184 10.6151
R2063 B.n213 B.n184 10.6151
R2064 B.n214 B.n213 10.6151
R2065 B.n215 B.n214 10.6151
R2066 B.n215 B.n182 10.6151
R2067 B.n219 B.n182 10.6151
R2068 B.n220 B.n219 10.6151
R2069 B.n221 B.n220 10.6151
R2070 B.n221 B.n180 10.6151
R2071 B.n225 B.n180 10.6151
R2072 B.n226 B.n225 10.6151
R2073 B.n227 B.n226 10.6151
R2074 B.n227 B.n178 10.6151
R2075 B.n231 B.n178 10.6151
R2076 B.n232 B.n231 10.6151
R2077 B.n233 B.n232 10.6151
R2078 B.n233 B.n176 10.6151
R2079 B.n237 B.n176 10.6151
R2080 B.n238 B.n237 10.6151
R2081 B.n239 B.n238 10.6151
R2082 B.n239 B.n174 10.6151
R2083 B.n243 B.n174 10.6151
R2084 B.n244 B.n243 10.6151
R2085 B.n245 B.n244 10.6151
R2086 B.n245 B.n172 10.6151
R2087 B.n249 B.n172 10.6151
R2088 B.n250 B.n249 10.6151
R2089 B.n251 B.n250 10.6151
R2090 B.n255 B.n170 10.6151
R2091 B.n256 B.n255 10.6151
R2092 B.n257 B.n256 10.6151
R2093 B.n257 B.n168 10.6151
R2094 B.n261 B.n168 10.6151
R2095 B.n262 B.n261 10.6151
R2096 B.n263 B.n262 10.6151
R2097 B.n263 B.n166 10.6151
R2098 B.n267 B.n166 10.6151
R2099 B.n268 B.n267 10.6151
R2100 B.n269 B.n268 10.6151
R2101 B.n269 B.n164 10.6151
R2102 B.n273 B.n164 10.6151
R2103 B.n274 B.n273 10.6151
R2104 B.n275 B.n274 10.6151
R2105 B.n275 B.n162 10.6151
R2106 B.n279 B.n162 10.6151
R2107 B.n280 B.n279 10.6151
R2108 B.n281 B.n280 10.6151
R2109 B.n281 B.n160 10.6151
R2110 B.n285 B.n160 10.6151
R2111 B.n286 B.n285 10.6151
R2112 B.n287 B.n286 10.6151
R2113 B.n287 B.n158 10.6151
R2114 B.n291 B.n158 10.6151
R2115 B.n292 B.n291 10.6151
R2116 B.n293 B.n292 10.6151
R2117 B.n293 B.n156 10.6151
R2118 B.n297 B.n156 10.6151
R2119 B.n298 B.n297 10.6151
R2120 B.n299 B.n298 10.6151
R2121 B.n299 B.n154 10.6151
R2122 B.n303 B.n154 10.6151
R2123 B.n304 B.n303 10.6151
R2124 B.n305 B.n304 10.6151
R2125 B.n305 B.n152 10.6151
R2126 B.n309 B.n152 10.6151
R2127 B.n310 B.n309 10.6151
R2128 B.n311 B.n310 10.6151
R2129 B.n311 B.n150 10.6151
R2130 B.n315 B.n150 10.6151
R2131 B.n316 B.n315 10.6151
R2132 B.n320 B.n316 10.6151
R2133 B.n324 B.n148 10.6151
R2134 B.n325 B.n324 10.6151
R2135 B.n326 B.n325 10.6151
R2136 B.n326 B.n146 10.6151
R2137 B.n330 B.n146 10.6151
R2138 B.n331 B.n330 10.6151
R2139 B.n332 B.n331 10.6151
R2140 B.n332 B.n144 10.6151
R2141 B.n336 B.n144 10.6151
R2142 B.n339 B.n338 10.6151
R2143 B.n339 B.n140 10.6151
R2144 B.n343 B.n140 10.6151
R2145 B.n344 B.n343 10.6151
R2146 B.n345 B.n344 10.6151
R2147 B.n345 B.n138 10.6151
R2148 B.n349 B.n138 10.6151
R2149 B.n350 B.n349 10.6151
R2150 B.n351 B.n350 10.6151
R2151 B.n351 B.n136 10.6151
R2152 B.n355 B.n136 10.6151
R2153 B.n356 B.n355 10.6151
R2154 B.n357 B.n356 10.6151
R2155 B.n357 B.n134 10.6151
R2156 B.n361 B.n134 10.6151
R2157 B.n362 B.n361 10.6151
R2158 B.n363 B.n362 10.6151
R2159 B.n363 B.n132 10.6151
R2160 B.n367 B.n132 10.6151
R2161 B.n368 B.n367 10.6151
R2162 B.n369 B.n368 10.6151
R2163 B.n369 B.n130 10.6151
R2164 B.n373 B.n130 10.6151
R2165 B.n374 B.n373 10.6151
R2166 B.n375 B.n374 10.6151
R2167 B.n375 B.n128 10.6151
R2168 B.n379 B.n128 10.6151
R2169 B.n380 B.n379 10.6151
R2170 B.n381 B.n380 10.6151
R2171 B.n381 B.n126 10.6151
R2172 B.n385 B.n126 10.6151
R2173 B.n386 B.n385 10.6151
R2174 B.n387 B.n386 10.6151
R2175 B.n387 B.n124 10.6151
R2176 B.n391 B.n124 10.6151
R2177 B.n392 B.n391 10.6151
R2178 B.n393 B.n392 10.6151
R2179 B.n393 B.n122 10.6151
R2180 B.n397 B.n122 10.6151
R2181 B.n398 B.n397 10.6151
R2182 B.n399 B.n398 10.6151
R2183 B.n399 B.n120 10.6151
R2184 B.n403 B.n120 10.6151
R2185 B.n615 B.n614 9.36635
R2186 B.n597 B.n54 9.36635
R2187 B.n320 B.n319 9.36635
R2188 B.n338 B.n337 9.36635
R2189 B.n745 B.n0 8.11757
R2190 B.n745 B.n1 8.11757
R2191 B.n614 B.n613 1.24928
R2192 B.n600 B.n54 1.24928
R2193 B.n319 B.n148 1.24928
R2194 B.n337 B.n336 1.24928
C0 B VTAIL 4.95779f
C1 VDD1 B 1.49554f
C2 VP VTAIL 8.947639f
C3 VDD2 B 1.57332f
C4 VDD1 VP 9.05759f
C5 B VN 1.09658f
C6 VDD2 VP 0.457635f
C7 VP VN 7.10757f
C8 VDD1 VTAIL 8.415251f
C9 VDD2 VTAIL 8.46578f
C10 VDD1 VDD2 1.47569f
C11 VN VTAIL 8.93354f
C12 VDD1 VN 0.150362f
C13 VDD2 VN 8.75142f
C14 w_n3320_n3532# B 9.45735f
C15 w_n3320_n3532# VP 7.04131f
C16 w_n3320_n3532# VTAIL 4.35628f
C17 VDD1 w_n3320_n3532# 1.78867f
C18 B VP 1.81314f
C19 VDD2 w_n3320_n3532# 1.87905f
C20 w_n3320_n3532# VN 6.61201f
C21 VDD2 VSUBS 1.671772f
C22 VDD1 VSUBS 2.213786f
C23 VTAIL VSUBS 1.27357f
C24 VN VSUBS 6.02112f
C25 VP VSUBS 3.005355f
C26 B VSUBS 4.422463f
C27 w_n3320_n3532# VSUBS 0.144181p
C28 B.n0 VSUBS 0.006157f
C29 B.n1 VSUBS 0.006157f
C30 B.n2 VSUBS 0.009106f
C31 B.n3 VSUBS 0.006978f
C32 B.n4 VSUBS 0.006978f
C33 B.n5 VSUBS 0.006978f
C34 B.n6 VSUBS 0.006978f
C35 B.n7 VSUBS 0.006978f
C36 B.n8 VSUBS 0.006978f
C37 B.n9 VSUBS 0.006978f
C38 B.n10 VSUBS 0.006978f
C39 B.n11 VSUBS 0.006978f
C40 B.n12 VSUBS 0.006978f
C41 B.n13 VSUBS 0.006978f
C42 B.n14 VSUBS 0.006978f
C43 B.n15 VSUBS 0.006978f
C44 B.n16 VSUBS 0.006978f
C45 B.n17 VSUBS 0.006978f
C46 B.n18 VSUBS 0.006978f
C47 B.n19 VSUBS 0.006978f
C48 B.n20 VSUBS 0.006978f
C49 B.n21 VSUBS 0.006978f
C50 B.n22 VSUBS 0.006978f
C51 B.n23 VSUBS 0.016854f
C52 B.n24 VSUBS 0.006978f
C53 B.n25 VSUBS 0.006978f
C54 B.n26 VSUBS 0.006978f
C55 B.n27 VSUBS 0.006978f
C56 B.n28 VSUBS 0.006978f
C57 B.n29 VSUBS 0.006978f
C58 B.n30 VSUBS 0.006978f
C59 B.n31 VSUBS 0.006978f
C60 B.n32 VSUBS 0.006978f
C61 B.n33 VSUBS 0.006978f
C62 B.n34 VSUBS 0.006978f
C63 B.n35 VSUBS 0.006978f
C64 B.n36 VSUBS 0.006978f
C65 B.n37 VSUBS 0.006978f
C66 B.n38 VSUBS 0.006978f
C67 B.n39 VSUBS 0.006978f
C68 B.n40 VSUBS 0.006978f
C69 B.n41 VSUBS 0.006978f
C70 B.n42 VSUBS 0.006978f
C71 B.n43 VSUBS 0.006978f
C72 B.n44 VSUBS 0.006978f
C73 B.n45 VSUBS 0.006978f
C74 B.t4 VSUBS 0.228804f
C75 B.t5 VSUBS 0.254912f
C76 B.t3 VSUBS 1.14988f
C77 B.n46 VSUBS 0.394968f
C78 B.n47 VSUBS 0.259753f
C79 B.n48 VSUBS 0.006978f
C80 B.n49 VSUBS 0.006978f
C81 B.n50 VSUBS 0.006978f
C82 B.n51 VSUBS 0.006978f
C83 B.t7 VSUBS 0.228807f
C84 B.t8 VSUBS 0.254915f
C85 B.t6 VSUBS 1.14988f
C86 B.n52 VSUBS 0.394966f
C87 B.n53 VSUBS 0.25975f
C88 B.n54 VSUBS 0.016167f
C89 B.n55 VSUBS 0.006978f
C90 B.n56 VSUBS 0.006978f
C91 B.n57 VSUBS 0.006978f
C92 B.n58 VSUBS 0.006978f
C93 B.n59 VSUBS 0.006978f
C94 B.n60 VSUBS 0.006978f
C95 B.n61 VSUBS 0.006978f
C96 B.n62 VSUBS 0.006978f
C97 B.n63 VSUBS 0.006978f
C98 B.n64 VSUBS 0.006978f
C99 B.n65 VSUBS 0.006978f
C100 B.n66 VSUBS 0.006978f
C101 B.n67 VSUBS 0.006978f
C102 B.n68 VSUBS 0.006978f
C103 B.n69 VSUBS 0.006978f
C104 B.n70 VSUBS 0.006978f
C105 B.n71 VSUBS 0.006978f
C106 B.n72 VSUBS 0.006978f
C107 B.n73 VSUBS 0.006978f
C108 B.n74 VSUBS 0.006978f
C109 B.n75 VSUBS 0.006978f
C110 B.n76 VSUBS 0.016854f
C111 B.n77 VSUBS 0.006978f
C112 B.n78 VSUBS 0.006978f
C113 B.n79 VSUBS 0.006978f
C114 B.n80 VSUBS 0.006978f
C115 B.n81 VSUBS 0.006978f
C116 B.n82 VSUBS 0.006978f
C117 B.n83 VSUBS 0.006978f
C118 B.n84 VSUBS 0.006978f
C119 B.n85 VSUBS 0.006978f
C120 B.n86 VSUBS 0.006978f
C121 B.n87 VSUBS 0.006978f
C122 B.n88 VSUBS 0.006978f
C123 B.n89 VSUBS 0.006978f
C124 B.n90 VSUBS 0.006978f
C125 B.n91 VSUBS 0.006978f
C126 B.n92 VSUBS 0.006978f
C127 B.n93 VSUBS 0.006978f
C128 B.n94 VSUBS 0.006978f
C129 B.n95 VSUBS 0.006978f
C130 B.n96 VSUBS 0.006978f
C131 B.n97 VSUBS 0.006978f
C132 B.n98 VSUBS 0.006978f
C133 B.n99 VSUBS 0.006978f
C134 B.n100 VSUBS 0.006978f
C135 B.n101 VSUBS 0.006978f
C136 B.n102 VSUBS 0.006978f
C137 B.n103 VSUBS 0.006978f
C138 B.n104 VSUBS 0.006978f
C139 B.n105 VSUBS 0.006978f
C140 B.n106 VSUBS 0.006978f
C141 B.n107 VSUBS 0.006978f
C142 B.n108 VSUBS 0.006978f
C143 B.n109 VSUBS 0.006978f
C144 B.n110 VSUBS 0.006978f
C145 B.n111 VSUBS 0.006978f
C146 B.n112 VSUBS 0.006978f
C147 B.n113 VSUBS 0.006978f
C148 B.n114 VSUBS 0.006978f
C149 B.n115 VSUBS 0.006978f
C150 B.n116 VSUBS 0.006978f
C151 B.n117 VSUBS 0.006978f
C152 B.n118 VSUBS 0.006978f
C153 B.n119 VSUBS 0.015573f
C154 B.n120 VSUBS 0.006978f
C155 B.n121 VSUBS 0.006978f
C156 B.n122 VSUBS 0.006978f
C157 B.n123 VSUBS 0.006978f
C158 B.n124 VSUBS 0.006978f
C159 B.n125 VSUBS 0.006978f
C160 B.n126 VSUBS 0.006978f
C161 B.n127 VSUBS 0.006978f
C162 B.n128 VSUBS 0.006978f
C163 B.n129 VSUBS 0.006978f
C164 B.n130 VSUBS 0.006978f
C165 B.n131 VSUBS 0.006978f
C166 B.n132 VSUBS 0.006978f
C167 B.n133 VSUBS 0.006978f
C168 B.n134 VSUBS 0.006978f
C169 B.n135 VSUBS 0.006978f
C170 B.n136 VSUBS 0.006978f
C171 B.n137 VSUBS 0.006978f
C172 B.n138 VSUBS 0.006978f
C173 B.n139 VSUBS 0.006978f
C174 B.n140 VSUBS 0.006978f
C175 B.n141 VSUBS 0.006978f
C176 B.t11 VSUBS 0.228807f
C177 B.t10 VSUBS 0.254915f
C178 B.t9 VSUBS 1.14988f
C179 B.n142 VSUBS 0.394966f
C180 B.n143 VSUBS 0.25975f
C181 B.n144 VSUBS 0.006978f
C182 B.n145 VSUBS 0.006978f
C183 B.n146 VSUBS 0.006978f
C184 B.n147 VSUBS 0.006978f
C185 B.n148 VSUBS 0.003899f
C186 B.n149 VSUBS 0.006978f
C187 B.n150 VSUBS 0.006978f
C188 B.n151 VSUBS 0.006978f
C189 B.n152 VSUBS 0.006978f
C190 B.n153 VSUBS 0.006978f
C191 B.n154 VSUBS 0.006978f
C192 B.n155 VSUBS 0.006978f
C193 B.n156 VSUBS 0.006978f
C194 B.n157 VSUBS 0.006978f
C195 B.n158 VSUBS 0.006978f
C196 B.n159 VSUBS 0.006978f
C197 B.n160 VSUBS 0.006978f
C198 B.n161 VSUBS 0.006978f
C199 B.n162 VSUBS 0.006978f
C200 B.n163 VSUBS 0.006978f
C201 B.n164 VSUBS 0.006978f
C202 B.n165 VSUBS 0.006978f
C203 B.n166 VSUBS 0.006978f
C204 B.n167 VSUBS 0.006978f
C205 B.n168 VSUBS 0.006978f
C206 B.n169 VSUBS 0.006978f
C207 B.n170 VSUBS 0.016854f
C208 B.n171 VSUBS 0.006978f
C209 B.n172 VSUBS 0.006978f
C210 B.n173 VSUBS 0.006978f
C211 B.n174 VSUBS 0.006978f
C212 B.n175 VSUBS 0.006978f
C213 B.n176 VSUBS 0.006978f
C214 B.n177 VSUBS 0.006978f
C215 B.n178 VSUBS 0.006978f
C216 B.n179 VSUBS 0.006978f
C217 B.n180 VSUBS 0.006978f
C218 B.n181 VSUBS 0.006978f
C219 B.n182 VSUBS 0.006978f
C220 B.n183 VSUBS 0.006978f
C221 B.n184 VSUBS 0.006978f
C222 B.n185 VSUBS 0.006978f
C223 B.n186 VSUBS 0.006978f
C224 B.n187 VSUBS 0.006978f
C225 B.n188 VSUBS 0.006978f
C226 B.n189 VSUBS 0.006978f
C227 B.n190 VSUBS 0.006978f
C228 B.n191 VSUBS 0.006978f
C229 B.n192 VSUBS 0.006978f
C230 B.n193 VSUBS 0.006978f
C231 B.n194 VSUBS 0.006978f
C232 B.n195 VSUBS 0.006978f
C233 B.n196 VSUBS 0.006978f
C234 B.n197 VSUBS 0.006978f
C235 B.n198 VSUBS 0.006978f
C236 B.n199 VSUBS 0.006978f
C237 B.n200 VSUBS 0.006978f
C238 B.n201 VSUBS 0.006978f
C239 B.n202 VSUBS 0.006978f
C240 B.n203 VSUBS 0.006978f
C241 B.n204 VSUBS 0.006978f
C242 B.n205 VSUBS 0.006978f
C243 B.n206 VSUBS 0.006978f
C244 B.n207 VSUBS 0.006978f
C245 B.n208 VSUBS 0.006978f
C246 B.n209 VSUBS 0.006978f
C247 B.n210 VSUBS 0.006978f
C248 B.n211 VSUBS 0.006978f
C249 B.n212 VSUBS 0.006978f
C250 B.n213 VSUBS 0.006978f
C251 B.n214 VSUBS 0.006978f
C252 B.n215 VSUBS 0.006978f
C253 B.n216 VSUBS 0.006978f
C254 B.n217 VSUBS 0.006978f
C255 B.n218 VSUBS 0.006978f
C256 B.n219 VSUBS 0.006978f
C257 B.n220 VSUBS 0.006978f
C258 B.n221 VSUBS 0.006978f
C259 B.n222 VSUBS 0.006978f
C260 B.n223 VSUBS 0.006978f
C261 B.n224 VSUBS 0.006978f
C262 B.n225 VSUBS 0.006978f
C263 B.n226 VSUBS 0.006978f
C264 B.n227 VSUBS 0.006978f
C265 B.n228 VSUBS 0.006978f
C266 B.n229 VSUBS 0.006978f
C267 B.n230 VSUBS 0.006978f
C268 B.n231 VSUBS 0.006978f
C269 B.n232 VSUBS 0.006978f
C270 B.n233 VSUBS 0.006978f
C271 B.n234 VSUBS 0.006978f
C272 B.n235 VSUBS 0.006978f
C273 B.n236 VSUBS 0.006978f
C274 B.n237 VSUBS 0.006978f
C275 B.n238 VSUBS 0.006978f
C276 B.n239 VSUBS 0.006978f
C277 B.n240 VSUBS 0.006978f
C278 B.n241 VSUBS 0.006978f
C279 B.n242 VSUBS 0.006978f
C280 B.n243 VSUBS 0.006978f
C281 B.n244 VSUBS 0.006978f
C282 B.n245 VSUBS 0.006978f
C283 B.n246 VSUBS 0.006978f
C284 B.n247 VSUBS 0.006978f
C285 B.n248 VSUBS 0.006978f
C286 B.n249 VSUBS 0.006978f
C287 B.n250 VSUBS 0.006978f
C288 B.n251 VSUBS 0.015573f
C289 B.n252 VSUBS 0.015573f
C290 B.n253 VSUBS 0.016854f
C291 B.n254 VSUBS 0.006978f
C292 B.n255 VSUBS 0.006978f
C293 B.n256 VSUBS 0.006978f
C294 B.n257 VSUBS 0.006978f
C295 B.n258 VSUBS 0.006978f
C296 B.n259 VSUBS 0.006978f
C297 B.n260 VSUBS 0.006978f
C298 B.n261 VSUBS 0.006978f
C299 B.n262 VSUBS 0.006978f
C300 B.n263 VSUBS 0.006978f
C301 B.n264 VSUBS 0.006978f
C302 B.n265 VSUBS 0.006978f
C303 B.n266 VSUBS 0.006978f
C304 B.n267 VSUBS 0.006978f
C305 B.n268 VSUBS 0.006978f
C306 B.n269 VSUBS 0.006978f
C307 B.n270 VSUBS 0.006978f
C308 B.n271 VSUBS 0.006978f
C309 B.n272 VSUBS 0.006978f
C310 B.n273 VSUBS 0.006978f
C311 B.n274 VSUBS 0.006978f
C312 B.n275 VSUBS 0.006978f
C313 B.n276 VSUBS 0.006978f
C314 B.n277 VSUBS 0.006978f
C315 B.n278 VSUBS 0.006978f
C316 B.n279 VSUBS 0.006978f
C317 B.n280 VSUBS 0.006978f
C318 B.n281 VSUBS 0.006978f
C319 B.n282 VSUBS 0.006978f
C320 B.n283 VSUBS 0.006978f
C321 B.n284 VSUBS 0.006978f
C322 B.n285 VSUBS 0.006978f
C323 B.n286 VSUBS 0.006978f
C324 B.n287 VSUBS 0.006978f
C325 B.n288 VSUBS 0.006978f
C326 B.n289 VSUBS 0.006978f
C327 B.n290 VSUBS 0.006978f
C328 B.n291 VSUBS 0.006978f
C329 B.n292 VSUBS 0.006978f
C330 B.n293 VSUBS 0.006978f
C331 B.n294 VSUBS 0.006978f
C332 B.n295 VSUBS 0.006978f
C333 B.n296 VSUBS 0.006978f
C334 B.n297 VSUBS 0.006978f
C335 B.n298 VSUBS 0.006978f
C336 B.n299 VSUBS 0.006978f
C337 B.n300 VSUBS 0.006978f
C338 B.n301 VSUBS 0.006978f
C339 B.n302 VSUBS 0.006978f
C340 B.n303 VSUBS 0.006978f
C341 B.n304 VSUBS 0.006978f
C342 B.n305 VSUBS 0.006978f
C343 B.n306 VSUBS 0.006978f
C344 B.n307 VSUBS 0.006978f
C345 B.n308 VSUBS 0.006978f
C346 B.n309 VSUBS 0.006978f
C347 B.n310 VSUBS 0.006978f
C348 B.n311 VSUBS 0.006978f
C349 B.n312 VSUBS 0.006978f
C350 B.n313 VSUBS 0.006978f
C351 B.n314 VSUBS 0.006978f
C352 B.n315 VSUBS 0.006978f
C353 B.n316 VSUBS 0.006978f
C354 B.t2 VSUBS 0.228804f
C355 B.t1 VSUBS 0.254912f
C356 B.t0 VSUBS 1.14988f
C357 B.n317 VSUBS 0.394968f
C358 B.n318 VSUBS 0.259753f
C359 B.n319 VSUBS 0.016167f
C360 B.n320 VSUBS 0.006567f
C361 B.n321 VSUBS 0.006978f
C362 B.n322 VSUBS 0.006978f
C363 B.n323 VSUBS 0.006978f
C364 B.n324 VSUBS 0.006978f
C365 B.n325 VSUBS 0.006978f
C366 B.n326 VSUBS 0.006978f
C367 B.n327 VSUBS 0.006978f
C368 B.n328 VSUBS 0.006978f
C369 B.n329 VSUBS 0.006978f
C370 B.n330 VSUBS 0.006978f
C371 B.n331 VSUBS 0.006978f
C372 B.n332 VSUBS 0.006978f
C373 B.n333 VSUBS 0.006978f
C374 B.n334 VSUBS 0.006978f
C375 B.n335 VSUBS 0.006978f
C376 B.n336 VSUBS 0.003899f
C377 B.n337 VSUBS 0.016167f
C378 B.n338 VSUBS 0.006567f
C379 B.n339 VSUBS 0.006978f
C380 B.n340 VSUBS 0.006978f
C381 B.n341 VSUBS 0.006978f
C382 B.n342 VSUBS 0.006978f
C383 B.n343 VSUBS 0.006978f
C384 B.n344 VSUBS 0.006978f
C385 B.n345 VSUBS 0.006978f
C386 B.n346 VSUBS 0.006978f
C387 B.n347 VSUBS 0.006978f
C388 B.n348 VSUBS 0.006978f
C389 B.n349 VSUBS 0.006978f
C390 B.n350 VSUBS 0.006978f
C391 B.n351 VSUBS 0.006978f
C392 B.n352 VSUBS 0.006978f
C393 B.n353 VSUBS 0.006978f
C394 B.n354 VSUBS 0.006978f
C395 B.n355 VSUBS 0.006978f
C396 B.n356 VSUBS 0.006978f
C397 B.n357 VSUBS 0.006978f
C398 B.n358 VSUBS 0.006978f
C399 B.n359 VSUBS 0.006978f
C400 B.n360 VSUBS 0.006978f
C401 B.n361 VSUBS 0.006978f
C402 B.n362 VSUBS 0.006978f
C403 B.n363 VSUBS 0.006978f
C404 B.n364 VSUBS 0.006978f
C405 B.n365 VSUBS 0.006978f
C406 B.n366 VSUBS 0.006978f
C407 B.n367 VSUBS 0.006978f
C408 B.n368 VSUBS 0.006978f
C409 B.n369 VSUBS 0.006978f
C410 B.n370 VSUBS 0.006978f
C411 B.n371 VSUBS 0.006978f
C412 B.n372 VSUBS 0.006978f
C413 B.n373 VSUBS 0.006978f
C414 B.n374 VSUBS 0.006978f
C415 B.n375 VSUBS 0.006978f
C416 B.n376 VSUBS 0.006978f
C417 B.n377 VSUBS 0.006978f
C418 B.n378 VSUBS 0.006978f
C419 B.n379 VSUBS 0.006978f
C420 B.n380 VSUBS 0.006978f
C421 B.n381 VSUBS 0.006978f
C422 B.n382 VSUBS 0.006978f
C423 B.n383 VSUBS 0.006978f
C424 B.n384 VSUBS 0.006978f
C425 B.n385 VSUBS 0.006978f
C426 B.n386 VSUBS 0.006978f
C427 B.n387 VSUBS 0.006978f
C428 B.n388 VSUBS 0.006978f
C429 B.n389 VSUBS 0.006978f
C430 B.n390 VSUBS 0.006978f
C431 B.n391 VSUBS 0.006978f
C432 B.n392 VSUBS 0.006978f
C433 B.n393 VSUBS 0.006978f
C434 B.n394 VSUBS 0.006978f
C435 B.n395 VSUBS 0.006978f
C436 B.n396 VSUBS 0.006978f
C437 B.n397 VSUBS 0.006978f
C438 B.n398 VSUBS 0.006978f
C439 B.n399 VSUBS 0.006978f
C440 B.n400 VSUBS 0.006978f
C441 B.n401 VSUBS 0.006978f
C442 B.n402 VSUBS 0.016854f
C443 B.n403 VSUBS 0.01602f
C444 B.n404 VSUBS 0.016407f
C445 B.n405 VSUBS 0.006978f
C446 B.n406 VSUBS 0.006978f
C447 B.n407 VSUBS 0.006978f
C448 B.n408 VSUBS 0.006978f
C449 B.n409 VSUBS 0.006978f
C450 B.n410 VSUBS 0.006978f
C451 B.n411 VSUBS 0.006978f
C452 B.n412 VSUBS 0.006978f
C453 B.n413 VSUBS 0.006978f
C454 B.n414 VSUBS 0.006978f
C455 B.n415 VSUBS 0.006978f
C456 B.n416 VSUBS 0.006978f
C457 B.n417 VSUBS 0.006978f
C458 B.n418 VSUBS 0.006978f
C459 B.n419 VSUBS 0.006978f
C460 B.n420 VSUBS 0.006978f
C461 B.n421 VSUBS 0.006978f
C462 B.n422 VSUBS 0.006978f
C463 B.n423 VSUBS 0.006978f
C464 B.n424 VSUBS 0.006978f
C465 B.n425 VSUBS 0.006978f
C466 B.n426 VSUBS 0.006978f
C467 B.n427 VSUBS 0.006978f
C468 B.n428 VSUBS 0.006978f
C469 B.n429 VSUBS 0.006978f
C470 B.n430 VSUBS 0.006978f
C471 B.n431 VSUBS 0.006978f
C472 B.n432 VSUBS 0.006978f
C473 B.n433 VSUBS 0.006978f
C474 B.n434 VSUBS 0.006978f
C475 B.n435 VSUBS 0.006978f
C476 B.n436 VSUBS 0.006978f
C477 B.n437 VSUBS 0.006978f
C478 B.n438 VSUBS 0.006978f
C479 B.n439 VSUBS 0.006978f
C480 B.n440 VSUBS 0.006978f
C481 B.n441 VSUBS 0.006978f
C482 B.n442 VSUBS 0.006978f
C483 B.n443 VSUBS 0.006978f
C484 B.n444 VSUBS 0.006978f
C485 B.n445 VSUBS 0.006978f
C486 B.n446 VSUBS 0.006978f
C487 B.n447 VSUBS 0.006978f
C488 B.n448 VSUBS 0.006978f
C489 B.n449 VSUBS 0.006978f
C490 B.n450 VSUBS 0.006978f
C491 B.n451 VSUBS 0.006978f
C492 B.n452 VSUBS 0.006978f
C493 B.n453 VSUBS 0.006978f
C494 B.n454 VSUBS 0.006978f
C495 B.n455 VSUBS 0.006978f
C496 B.n456 VSUBS 0.006978f
C497 B.n457 VSUBS 0.006978f
C498 B.n458 VSUBS 0.006978f
C499 B.n459 VSUBS 0.006978f
C500 B.n460 VSUBS 0.006978f
C501 B.n461 VSUBS 0.006978f
C502 B.n462 VSUBS 0.006978f
C503 B.n463 VSUBS 0.006978f
C504 B.n464 VSUBS 0.006978f
C505 B.n465 VSUBS 0.006978f
C506 B.n466 VSUBS 0.006978f
C507 B.n467 VSUBS 0.006978f
C508 B.n468 VSUBS 0.006978f
C509 B.n469 VSUBS 0.006978f
C510 B.n470 VSUBS 0.006978f
C511 B.n471 VSUBS 0.006978f
C512 B.n472 VSUBS 0.006978f
C513 B.n473 VSUBS 0.006978f
C514 B.n474 VSUBS 0.006978f
C515 B.n475 VSUBS 0.006978f
C516 B.n476 VSUBS 0.006978f
C517 B.n477 VSUBS 0.006978f
C518 B.n478 VSUBS 0.006978f
C519 B.n479 VSUBS 0.006978f
C520 B.n480 VSUBS 0.006978f
C521 B.n481 VSUBS 0.006978f
C522 B.n482 VSUBS 0.006978f
C523 B.n483 VSUBS 0.006978f
C524 B.n484 VSUBS 0.006978f
C525 B.n485 VSUBS 0.006978f
C526 B.n486 VSUBS 0.006978f
C527 B.n487 VSUBS 0.006978f
C528 B.n488 VSUBS 0.006978f
C529 B.n489 VSUBS 0.006978f
C530 B.n490 VSUBS 0.006978f
C531 B.n491 VSUBS 0.006978f
C532 B.n492 VSUBS 0.006978f
C533 B.n493 VSUBS 0.006978f
C534 B.n494 VSUBS 0.006978f
C535 B.n495 VSUBS 0.006978f
C536 B.n496 VSUBS 0.006978f
C537 B.n497 VSUBS 0.006978f
C538 B.n498 VSUBS 0.006978f
C539 B.n499 VSUBS 0.006978f
C540 B.n500 VSUBS 0.006978f
C541 B.n501 VSUBS 0.006978f
C542 B.n502 VSUBS 0.006978f
C543 B.n503 VSUBS 0.006978f
C544 B.n504 VSUBS 0.006978f
C545 B.n505 VSUBS 0.006978f
C546 B.n506 VSUBS 0.006978f
C547 B.n507 VSUBS 0.006978f
C548 B.n508 VSUBS 0.006978f
C549 B.n509 VSUBS 0.006978f
C550 B.n510 VSUBS 0.006978f
C551 B.n511 VSUBS 0.006978f
C552 B.n512 VSUBS 0.006978f
C553 B.n513 VSUBS 0.006978f
C554 B.n514 VSUBS 0.006978f
C555 B.n515 VSUBS 0.006978f
C556 B.n516 VSUBS 0.006978f
C557 B.n517 VSUBS 0.006978f
C558 B.n518 VSUBS 0.006978f
C559 B.n519 VSUBS 0.006978f
C560 B.n520 VSUBS 0.006978f
C561 B.n521 VSUBS 0.006978f
C562 B.n522 VSUBS 0.006978f
C563 B.n523 VSUBS 0.006978f
C564 B.n524 VSUBS 0.006978f
C565 B.n525 VSUBS 0.006978f
C566 B.n526 VSUBS 0.006978f
C567 B.n527 VSUBS 0.006978f
C568 B.n528 VSUBS 0.006978f
C569 B.n529 VSUBS 0.006978f
C570 B.n530 VSUBS 0.006978f
C571 B.n531 VSUBS 0.015573f
C572 B.n532 VSUBS 0.015573f
C573 B.n533 VSUBS 0.016854f
C574 B.n534 VSUBS 0.006978f
C575 B.n535 VSUBS 0.006978f
C576 B.n536 VSUBS 0.006978f
C577 B.n537 VSUBS 0.006978f
C578 B.n538 VSUBS 0.006978f
C579 B.n539 VSUBS 0.006978f
C580 B.n540 VSUBS 0.006978f
C581 B.n541 VSUBS 0.006978f
C582 B.n542 VSUBS 0.006978f
C583 B.n543 VSUBS 0.006978f
C584 B.n544 VSUBS 0.006978f
C585 B.n545 VSUBS 0.006978f
C586 B.n546 VSUBS 0.006978f
C587 B.n547 VSUBS 0.006978f
C588 B.n548 VSUBS 0.006978f
C589 B.n549 VSUBS 0.006978f
C590 B.n550 VSUBS 0.006978f
C591 B.n551 VSUBS 0.006978f
C592 B.n552 VSUBS 0.006978f
C593 B.n553 VSUBS 0.006978f
C594 B.n554 VSUBS 0.006978f
C595 B.n555 VSUBS 0.006978f
C596 B.n556 VSUBS 0.006978f
C597 B.n557 VSUBS 0.006978f
C598 B.n558 VSUBS 0.006978f
C599 B.n559 VSUBS 0.006978f
C600 B.n560 VSUBS 0.006978f
C601 B.n561 VSUBS 0.006978f
C602 B.n562 VSUBS 0.006978f
C603 B.n563 VSUBS 0.006978f
C604 B.n564 VSUBS 0.006978f
C605 B.n565 VSUBS 0.006978f
C606 B.n566 VSUBS 0.006978f
C607 B.n567 VSUBS 0.006978f
C608 B.n568 VSUBS 0.006978f
C609 B.n569 VSUBS 0.006978f
C610 B.n570 VSUBS 0.006978f
C611 B.n571 VSUBS 0.006978f
C612 B.n572 VSUBS 0.006978f
C613 B.n573 VSUBS 0.006978f
C614 B.n574 VSUBS 0.006978f
C615 B.n575 VSUBS 0.006978f
C616 B.n576 VSUBS 0.006978f
C617 B.n577 VSUBS 0.006978f
C618 B.n578 VSUBS 0.006978f
C619 B.n579 VSUBS 0.006978f
C620 B.n580 VSUBS 0.006978f
C621 B.n581 VSUBS 0.006978f
C622 B.n582 VSUBS 0.006978f
C623 B.n583 VSUBS 0.006978f
C624 B.n584 VSUBS 0.006978f
C625 B.n585 VSUBS 0.006978f
C626 B.n586 VSUBS 0.006978f
C627 B.n587 VSUBS 0.006978f
C628 B.n588 VSUBS 0.006978f
C629 B.n589 VSUBS 0.006978f
C630 B.n590 VSUBS 0.006978f
C631 B.n591 VSUBS 0.006978f
C632 B.n592 VSUBS 0.006978f
C633 B.n593 VSUBS 0.006978f
C634 B.n594 VSUBS 0.006978f
C635 B.n595 VSUBS 0.006978f
C636 B.n596 VSUBS 0.006978f
C637 B.n597 VSUBS 0.006567f
C638 B.n598 VSUBS 0.006978f
C639 B.n599 VSUBS 0.006978f
C640 B.n600 VSUBS 0.003899f
C641 B.n601 VSUBS 0.006978f
C642 B.n602 VSUBS 0.006978f
C643 B.n603 VSUBS 0.006978f
C644 B.n604 VSUBS 0.006978f
C645 B.n605 VSUBS 0.006978f
C646 B.n606 VSUBS 0.006978f
C647 B.n607 VSUBS 0.006978f
C648 B.n608 VSUBS 0.006978f
C649 B.n609 VSUBS 0.006978f
C650 B.n610 VSUBS 0.006978f
C651 B.n611 VSUBS 0.006978f
C652 B.n612 VSUBS 0.006978f
C653 B.n613 VSUBS 0.003899f
C654 B.n614 VSUBS 0.016167f
C655 B.n615 VSUBS 0.006567f
C656 B.n616 VSUBS 0.006978f
C657 B.n617 VSUBS 0.006978f
C658 B.n618 VSUBS 0.006978f
C659 B.n619 VSUBS 0.006978f
C660 B.n620 VSUBS 0.006978f
C661 B.n621 VSUBS 0.006978f
C662 B.n622 VSUBS 0.006978f
C663 B.n623 VSUBS 0.006978f
C664 B.n624 VSUBS 0.006978f
C665 B.n625 VSUBS 0.006978f
C666 B.n626 VSUBS 0.006978f
C667 B.n627 VSUBS 0.006978f
C668 B.n628 VSUBS 0.006978f
C669 B.n629 VSUBS 0.006978f
C670 B.n630 VSUBS 0.006978f
C671 B.n631 VSUBS 0.006978f
C672 B.n632 VSUBS 0.006978f
C673 B.n633 VSUBS 0.006978f
C674 B.n634 VSUBS 0.006978f
C675 B.n635 VSUBS 0.006978f
C676 B.n636 VSUBS 0.006978f
C677 B.n637 VSUBS 0.006978f
C678 B.n638 VSUBS 0.006978f
C679 B.n639 VSUBS 0.006978f
C680 B.n640 VSUBS 0.006978f
C681 B.n641 VSUBS 0.006978f
C682 B.n642 VSUBS 0.006978f
C683 B.n643 VSUBS 0.006978f
C684 B.n644 VSUBS 0.006978f
C685 B.n645 VSUBS 0.006978f
C686 B.n646 VSUBS 0.006978f
C687 B.n647 VSUBS 0.006978f
C688 B.n648 VSUBS 0.006978f
C689 B.n649 VSUBS 0.006978f
C690 B.n650 VSUBS 0.006978f
C691 B.n651 VSUBS 0.006978f
C692 B.n652 VSUBS 0.006978f
C693 B.n653 VSUBS 0.006978f
C694 B.n654 VSUBS 0.006978f
C695 B.n655 VSUBS 0.006978f
C696 B.n656 VSUBS 0.006978f
C697 B.n657 VSUBS 0.006978f
C698 B.n658 VSUBS 0.006978f
C699 B.n659 VSUBS 0.006978f
C700 B.n660 VSUBS 0.006978f
C701 B.n661 VSUBS 0.006978f
C702 B.n662 VSUBS 0.006978f
C703 B.n663 VSUBS 0.006978f
C704 B.n664 VSUBS 0.006978f
C705 B.n665 VSUBS 0.006978f
C706 B.n666 VSUBS 0.006978f
C707 B.n667 VSUBS 0.006978f
C708 B.n668 VSUBS 0.006978f
C709 B.n669 VSUBS 0.006978f
C710 B.n670 VSUBS 0.006978f
C711 B.n671 VSUBS 0.006978f
C712 B.n672 VSUBS 0.006978f
C713 B.n673 VSUBS 0.006978f
C714 B.n674 VSUBS 0.006978f
C715 B.n675 VSUBS 0.006978f
C716 B.n676 VSUBS 0.006978f
C717 B.n677 VSUBS 0.006978f
C718 B.n678 VSUBS 0.006978f
C719 B.n679 VSUBS 0.006978f
C720 B.n680 VSUBS 0.016854f
C721 B.n681 VSUBS 0.015573f
C722 B.n682 VSUBS 0.015573f
C723 B.n683 VSUBS 0.006978f
C724 B.n684 VSUBS 0.006978f
C725 B.n685 VSUBS 0.006978f
C726 B.n686 VSUBS 0.006978f
C727 B.n687 VSUBS 0.006978f
C728 B.n688 VSUBS 0.006978f
C729 B.n689 VSUBS 0.006978f
C730 B.n690 VSUBS 0.006978f
C731 B.n691 VSUBS 0.006978f
C732 B.n692 VSUBS 0.006978f
C733 B.n693 VSUBS 0.006978f
C734 B.n694 VSUBS 0.006978f
C735 B.n695 VSUBS 0.006978f
C736 B.n696 VSUBS 0.006978f
C737 B.n697 VSUBS 0.006978f
C738 B.n698 VSUBS 0.006978f
C739 B.n699 VSUBS 0.006978f
C740 B.n700 VSUBS 0.006978f
C741 B.n701 VSUBS 0.006978f
C742 B.n702 VSUBS 0.006978f
C743 B.n703 VSUBS 0.006978f
C744 B.n704 VSUBS 0.006978f
C745 B.n705 VSUBS 0.006978f
C746 B.n706 VSUBS 0.006978f
C747 B.n707 VSUBS 0.006978f
C748 B.n708 VSUBS 0.006978f
C749 B.n709 VSUBS 0.006978f
C750 B.n710 VSUBS 0.006978f
C751 B.n711 VSUBS 0.006978f
C752 B.n712 VSUBS 0.006978f
C753 B.n713 VSUBS 0.006978f
C754 B.n714 VSUBS 0.006978f
C755 B.n715 VSUBS 0.006978f
C756 B.n716 VSUBS 0.006978f
C757 B.n717 VSUBS 0.006978f
C758 B.n718 VSUBS 0.006978f
C759 B.n719 VSUBS 0.006978f
C760 B.n720 VSUBS 0.006978f
C761 B.n721 VSUBS 0.006978f
C762 B.n722 VSUBS 0.006978f
C763 B.n723 VSUBS 0.006978f
C764 B.n724 VSUBS 0.006978f
C765 B.n725 VSUBS 0.006978f
C766 B.n726 VSUBS 0.006978f
C767 B.n727 VSUBS 0.006978f
C768 B.n728 VSUBS 0.006978f
C769 B.n729 VSUBS 0.006978f
C770 B.n730 VSUBS 0.006978f
C771 B.n731 VSUBS 0.006978f
C772 B.n732 VSUBS 0.006978f
C773 B.n733 VSUBS 0.006978f
C774 B.n734 VSUBS 0.006978f
C775 B.n735 VSUBS 0.006978f
C776 B.n736 VSUBS 0.006978f
C777 B.n737 VSUBS 0.006978f
C778 B.n738 VSUBS 0.006978f
C779 B.n739 VSUBS 0.006978f
C780 B.n740 VSUBS 0.006978f
C781 B.n741 VSUBS 0.006978f
C782 B.n742 VSUBS 0.006978f
C783 B.n743 VSUBS 0.009106f
C784 B.n744 VSUBS 0.0097f
C785 B.n745 VSUBS 0.019289f
C786 VDD2.t4 VSUBS 0.249891f
C787 VDD2.t0 VSUBS 0.249891f
C788 VDD2.n0 VSUBS 1.97884f
C789 VDD2.t1 VSUBS 0.249891f
C790 VDD2.t6 VSUBS 0.249891f
C791 VDD2.n1 VSUBS 1.97884f
C792 VDD2.n2 VSUBS 3.48336f
C793 VDD2.t7 VSUBS 0.249891f
C794 VDD2.t2 VSUBS 0.249891f
C795 VDD2.n3 VSUBS 1.9695f
C796 VDD2.n4 VSUBS 3.04195f
C797 VDD2.t3 VSUBS 0.249891f
C798 VDD2.t5 VSUBS 0.249891f
C799 VDD2.n5 VSUBS 1.9788f
C800 VN.n0 VSUBS 0.032659f
C801 VN.t1 VSUBS 2.30859f
C802 VN.n1 VSUBS 0.037366f
C803 VN.n2 VSUBS 0.032659f
C804 VN.t6 VSUBS 2.30859f
C805 VN.n3 VSUBS 0.065257f
C806 VN.n4 VSUBS 0.032659f
C807 VN.t7 VSUBS 2.30859f
C808 VN.n5 VSUBS 0.895307f
C809 VN.t3 VSUBS 2.47914f
C810 VN.n6 VSUBS 0.903653f
C811 VN.n7 VSUBS 0.245259f
C812 VN.n8 VSUBS 0.041542f
C813 VN.n9 VSUBS 0.065257f
C814 VN.n10 VSUBS 0.026429f
C815 VN.n11 VSUBS 0.032659f
C816 VN.n12 VSUBS 0.032659f
C817 VN.n13 VSUBS 0.032659f
C818 VN.n14 VSUBS 0.041542f
C819 VN.n15 VSUBS 0.820276f
C820 VN.n16 VSUBS 0.050603f
C821 VN.n17 VSUBS 0.056796f
C822 VN.n18 VSUBS 0.032659f
C823 VN.n19 VSUBS 0.032659f
C824 VN.n20 VSUBS 0.032659f
C825 VN.n21 VSUBS 0.062781f
C826 VN.n22 VSUBS 0.03248f
C827 VN.n23 VSUBS 0.902573f
C828 VN.n24 VSUBS 0.037109f
C829 VN.n25 VSUBS 0.032659f
C830 VN.t0 VSUBS 2.30859f
C831 VN.n26 VSUBS 0.037366f
C832 VN.n27 VSUBS 0.032659f
C833 VN.t5 VSUBS 2.30859f
C834 VN.n28 VSUBS 0.065257f
C835 VN.n29 VSUBS 0.032659f
C836 VN.t4 VSUBS 2.30859f
C837 VN.n30 VSUBS 0.895307f
C838 VN.t2 VSUBS 2.47914f
C839 VN.n31 VSUBS 0.903653f
C840 VN.n32 VSUBS 0.245259f
C841 VN.n33 VSUBS 0.041542f
C842 VN.n34 VSUBS 0.065257f
C843 VN.n35 VSUBS 0.026429f
C844 VN.n36 VSUBS 0.032659f
C845 VN.n37 VSUBS 0.032659f
C846 VN.n38 VSUBS 0.032659f
C847 VN.n39 VSUBS 0.041542f
C848 VN.n40 VSUBS 0.820276f
C849 VN.n41 VSUBS 0.050603f
C850 VN.n42 VSUBS 0.056796f
C851 VN.n43 VSUBS 0.032659f
C852 VN.n44 VSUBS 0.032659f
C853 VN.n45 VSUBS 0.032659f
C854 VN.n46 VSUBS 0.062781f
C855 VN.n47 VSUBS 0.03248f
C856 VN.n48 VSUBS 0.902573f
C857 VN.n49 VSUBS 1.74034f
C858 VTAIL.t15 VSUBS 0.247318f
C859 VTAIL.t2 VSUBS 0.247318f
C860 VTAIL.n0 VSUBS 1.81161f
C861 VTAIL.n1 VSUBS 0.734534f
C862 VTAIL.n2 VSUBS 0.026929f
C863 VTAIL.n3 VSUBS 0.024413f
C864 VTAIL.n4 VSUBS 0.013118f
C865 VTAIL.n5 VSUBS 0.031007f
C866 VTAIL.n6 VSUBS 0.01389f
C867 VTAIL.n7 VSUBS 0.024413f
C868 VTAIL.n8 VSUBS 0.013118f
C869 VTAIL.n9 VSUBS 0.031007f
C870 VTAIL.n10 VSUBS 0.01389f
C871 VTAIL.n11 VSUBS 0.024413f
C872 VTAIL.n12 VSUBS 0.013118f
C873 VTAIL.n13 VSUBS 0.031007f
C874 VTAIL.n14 VSUBS 0.01389f
C875 VTAIL.n15 VSUBS 0.024413f
C876 VTAIL.n16 VSUBS 0.013118f
C877 VTAIL.n17 VSUBS 0.031007f
C878 VTAIL.n18 VSUBS 0.01389f
C879 VTAIL.n19 VSUBS 0.024413f
C880 VTAIL.n20 VSUBS 0.013118f
C881 VTAIL.n21 VSUBS 0.031007f
C882 VTAIL.n22 VSUBS 0.01389f
C883 VTAIL.n23 VSUBS 0.201314f
C884 VTAIL.t1 VSUBS 0.066882f
C885 VTAIL.n24 VSUBS 0.023255f
C886 VTAIL.n25 VSUBS 0.023325f
C887 VTAIL.n26 VSUBS 0.013118f
C888 VTAIL.n27 VSUBS 1.28719f
C889 VTAIL.n28 VSUBS 0.024413f
C890 VTAIL.n29 VSUBS 0.013118f
C891 VTAIL.n30 VSUBS 0.01389f
C892 VTAIL.n31 VSUBS 0.031007f
C893 VTAIL.n32 VSUBS 0.031007f
C894 VTAIL.n33 VSUBS 0.01389f
C895 VTAIL.n34 VSUBS 0.013118f
C896 VTAIL.n35 VSUBS 0.024413f
C897 VTAIL.n36 VSUBS 0.024413f
C898 VTAIL.n37 VSUBS 0.013118f
C899 VTAIL.n38 VSUBS 0.01389f
C900 VTAIL.n39 VSUBS 0.031007f
C901 VTAIL.n40 VSUBS 0.031007f
C902 VTAIL.n41 VSUBS 0.031007f
C903 VTAIL.n42 VSUBS 0.01389f
C904 VTAIL.n43 VSUBS 0.013118f
C905 VTAIL.n44 VSUBS 0.024413f
C906 VTAIL.n45 VSUBS 0.024413f
C907 VTAIL.n46 VSUBS 0.013118f
C908 VTAIL.n47 VSUBS 0.013504f
C909 VTAIL.n48 VSUBS 0.013504f
C910 VTAIL.n49 VSUBS 0.031007f
C911 VTAIL.n50 VSUBS 0.031007f
C912 VTAIL.n51 VSUBS 0.01389f
C913 VTAIL.n52 VSUBS 0.013118f
C914 VTAIL.n53 VSUBS 0.024413f
C915 VTAIL.n54 VSUBS 0.024413f
C916 VTAIL.n55 VSUBS 0.013118f
C917 VTAIL.n56 VSUBS 0.01389f
C918 VTAIL.n57 VSUBS 0.031007f
C919 VTAIL.n58 VSUBS 0.031007f
C920 VTAIL.n59 VSUBS 0.01389f
C921 VTAIL.n60 VSUBS 0.013118f
C922 VTAIL.n61 VSUBS 0.024413f
C923 VTAIL.n62 VSUBS 0.024413f
C924 VTAIL.n63 VSUBS 0.013118f
C925 VTAIL.n64 VSUBS 0.01389f
C926 VTAIL.n65 VSUBS 0.031007f
C927 VTAIL.n66 VSUBS 0.075422f
C928 VTAIL.n67 VSUBS 0.01389f
C929 VTAIL.n68 VSUBS 0.013118f
C930 VTAIL.n69 VSUBS 0.055762f
C931 VTAIL.n70 VSUBS 0.037924f
C932 VTAIL.n71 VSUBS 0.216792f
C933 VTAIL.n72 VSUBS 0.026929f
C934 VTAIL.n73 VSUBS 0.024413f
C935 VTAIL.n74 VSUBS 0.013118f
C936 VTAIL.n75 VSUBS 0.031007f
C937 VTAIL.n76 VSUBS 0.01389f
C938 VTAIL.n77 VSUBS 0.024413f
C939 VTAIL.n78 VSUBS 0.013118f
C940 VTAIL.n79 VSUBS 0.031007f
C941 VTAIL.n80 VSUBS 0.01389f
C942 VTAIL.n81 VSUBS 0.024413f
C943 VTAIL.n82 VSUBS 0.013118f
C944 VTAIL.n83 VSUBS 0.031007f
C945 VTAIL.n84 VSUBS 0.01389f
C946 VTAIL.n85 VSUBS 0.024413f
C947 VTAIL.n86 VSUBS 0.013118f
C948 VTAIL.n87 VSUBS 0.031007f
C949 VTAIL.n88 VSUBS 0.01389f
C950 VTAIL.n89 VSUBS 0.024413f
C951 VTAIL.n90 VSUBS 0.013118f
C952 VTAIL.n91 VSUBS 0.031007f
C953 VTAIL.n92 VSUBS 0.01389f
C954 VTAIL.n93 VSUBS 0.201314f
C955 VTAIL.t8 VSUBS 0.066882f
C956 VTAIL.n94 VSUBS 0.023255f
C957 VTAIL.n95 VSUBS 0.023325f
C958 VTAIL.n96 VSUBS 0.013118f
C959 VTAIL.n97 VSUBS 1.28719f
C960 VTAIL.n98 VSUBS 0.024413f
C961 VTAIL.n99 VSUBS 0.013118f
C962 VTAIL.n100 VSUBS 0.01389f
C963 VTAIL.n101 VSUBS 0.031007f
C964 VTAIL.n102 VSUBS 0.031007f
C965 VTAIL.n103 VSUBS 0.01389f
C966 VTAIL.n104 VSUBS 0.013118f
C967 VTAIL.n105 VSUBS 0.024413f
C968 VTAIL.n106 VSUBS 0.024413f
C969 VTAIL.n107 VSUBS 0.013118f
C970 VTAIL.n108 VSUBS 0.01389f
C971 VTAIL.n109 VSUBS 0.031007f
C972 VTAIL.n110 VSUBS 0.031007f
C973 VTAIL.n111 VSUBS 0.031007f
C974 VTAIL.n112 VSUBS 0.01389f
C975 VTAIL.n113 VSUBS 0.013118f
C976 VTAIL.n114 VSUBS 0.024413f
C977 VTAIL.n115 VSUBS 0.024413f
C978 VTAIL.n116 VSUBS 0.013118f
C979 VTAIL.n117 VSUBS 0.013504f
C980 VTAIL.n118 VSUBS 0.013504f
C981 VTAIL.n119 VSUBS 0.031007f
C982 VTAIL.n120 VSUBS 0.031007f
C983 VTAIL.n121 VSUBS 0.01389f
C984 VTAIL.n122 VSUBS 0.013118f
C985 VTAIL.n123 VSUBS 0.024413f
C986 VTAIL.n124 VSUBS 0.024413f
C987 VTAIL.n125 VSUBS 0.013118f
C988 VTAIL.n126 VSUBS 0.01389f
C989 VTAIL.n127 VSUBS 0.031007f
C990 VTAIL.n128 VSUBS 0.031007f
C991 VTAIL.n129 VSUBS 0.01389f
C992 VTAIL.n130 VSUBS 0.013118f
C993 VTAIL.n131 VSUBS 0.024413f
C994 VTAIL.n132 VSUBS 0.024413f
C995 VTAIL.n133 VSUBS 0.013118f
C996 VTAIL.n134 VSUBS 0.01389f
C997 VTAIL.n135 VSUBS 0.031007f
C998 VTAIL.n136 VSUBS 0.075422f
C999 VTAIL.n137 VSUBS 0.01389f
C1000 VTAIL.n138 VSUBS 0.013118f
C1001 VTAIL.n139 VSUBS 0.055762f
C1002 VTAIL.n140 VSUBS 0.037924f
C1003 VTAIL.n141 VSUBS 0.216792f
C1004 VTAIL.t7 VSUBS 0.247318f
C1005 VTAIL.t12 VSUBS 0.247318f
C1006 VTAIL.n142 VSUBS 1.81161f
C1007 VTAIL.n143 VSUBS 0.889316f
C1008 VTAIL.n144 VSUBS 0.026929f
C1009 VTAIL.n145 VSUBS 0.024413f
C1010 VTAIL.n146 VSUBS 0.013118f
C1011 VTAIL.n147 VSUBS 0.031007f
C1012 VTAIL.n148 VSUBS 0.01389f
C1013 VTAIL.n149 VSUBS 0.024413f
C1014 VTAIL.n150 VSUBS 0.013118f
C1015 VTAIL.n151 VSUBS 0.031007f
C1016 VTAIL.n152 VSUBS 0.01389f
C1017 VTAIL.n153 VSUBS 0.024413f
C1018 VTAIL.n154 VSUBS 0.013118f
C1019 VTAIL.n155 VSUBS 0.031007f
C1020 VTAIL.n156 VSUBS 0.01389f
C1021 VTAIL.n157 VSUBS 0.024413f
C1022 VTAIL.n158 VSUBS 0.013118f
C1023 VTAIL.n159 VSUBS 0.031007f
C1024 VTAIL.n160 VSUBS 0.01389f
C1025 VTAIL.n161 VSUBS 0.024413f
C1026 VTAIL.n162 VSUBS 0.013118f
C1027 VTAIL.n163 VSUBS 0.031007f
C1028 VTAIL.n164 VSUBS 0.01389f
C1029 VTAIL.n165 VSUBS 0.201314f
C1030 VTAIL.t11 VSUBS 0.066882f
C1031 VTAIL.n166 VSUBS 0.023255f
C1032 VTAIL.n167 VSUBS 0.023325f
C1033 VTAIL.n168 VSUBS 0.013118f
C1034 VTAIL.n169 VSUBS 1.28719f
C1035 VTAIL.n170 VSUBS 0.024413f
C1036 VTAIL.n171 VSUBS 0.013118f
C1037 VTAIL.n172 VSUBS 0.01389f
C1038 VTAIL.n173 VSUBS 0.031007f
C1039 VTAIL.n174 VSUBS 0.031007f
C1040 VTAIL.n175 VSUBS 0.01389f
C1041 VTAIL.n176 VSUBS 0.013118f
C1042 VTAIL.n177 VSUBS 0.024413f
C1043 VTAIL.n178 VSUBS 0.024413f
C1044 VTAIL.n179 VSUBS 0.013118f
C1045 VTAIL.n180 VSUBS 0.01389f
C1046 VTAIL.n181 VSUBS 0.031007f
C1047 VTAIL.n182 VSUBS 0.031007f
C1048 VTAIL.n183 VSUBS 0.031007f
C1049 VTAIL.n184 VSUBS 0.01389f
C1050 VTAIL.n185 VSUBS 0.013118f
C1051 VTAIL.n186 VSUBS 0.024413f
C1052 VTAIL.n187 VSUBS 0.024413f
C1053 VTAIL.n188 VSUBS 0.013118f
C1054 VTAIL.n189 VSUBS 0.013504f
C1055 VTAIL.n190 VSUBS 0.013504f
C1056 VTAIL.n191 VSUBS 0.031007f
C1057 VTAIL.n192 VSUBS 0.031007f
C1058 VTAIL.n193 VSUBS 0.01389f
C1059 VTAIL.n194 VSUBS 0.013118f
C1060 VTAIL.n195 VSUBS 0.024413f
C1061 VTAIL.n196 VSUBS 0.024413f
C1062 VTAIL.n197 VSUBS 0.013118f
C1063 VTAIL.n198 VSUBS 0.01389f
C1064 VTAIL.n199 VSUBS 0.031007f
C1065 VTAIL.n200 VSUBS 0.031007f
C1066 VTAIL.n201 VSUBS 0.01389f
C1067 VTAIL.n202 VSUBS 0.013118f
C1068 VTAIL.n203 VSUBS 0.024413f
C1069 VTAIL.n204 VSUBS 0.024413f
C1070 VTAIL.n205 VSUBS 0.013118f
C1071 VTAIL.n206 VSUBS 0.01389f
C1072 VTAIL.n207 VSUBS 0.031007f
C1073 VTAIL.n208 VSUBS 0.075422f
C1074 VTAIL.n209 VSUBS 0.01389f
C1075 VTAIL.n210 VSUBS 0.013118f
C1076 VTAIL.n211 VSUBS 0.055762f
C1077 VTAIL.n212 VSUBS 0.037924f
C1078 VTAIL.n213 VSUBS 1.54017f
C1079 VTAIL.n214 VSUBS 0.026929f
C1080 VTAIL.n215 VSUBS 0.024413f
C1081 VTAIL.n216 VSUBS 0.013118f
C1082 VTAIL.n217 VSUBS 0.031007f
C1083 VTAIL.n218 VSUBS 0.01389f
C1084 VTAIL.n219 VSUBS 0.024413f
C1085 VTAIL.n220 VSUBS 0.013118f
C1086 VTAIL.n221 VSUBS 0.031007f
C1087 VTAIL.n222 VSUBS 0.01389f
C1088 VTAIL.n223 VSUBS 0.024413f
C1089 VTAIL.n224 VSUBS 0.013118f
C1090 VTAIL.n225 VSUBS 0.031007f
C1091 VTAIL.n226 VSUBS 0.01389f
C1092 VTAIL.n227 VSUBS 0.024413f
C1093 VTAIL.n228 VSUBS 0.013118f
C1094 VTAIL.n229 VSUBS 0.031007f
C1095 VTAIL.n230 VSUBS 0.031007f
C1096 VTAIL.n231 VSUBS 0.01389f
C1097 VTAIL.n232 VSUBS 0.024413f
C1098 VTAIL.n233 VSUBS 0.013118f
C1099 VTAIL.n234 VSUBS 0.031007f
C1100 VTAIL.n235 VSUBS 0.01389f
C1101 VTAIL.n236 VSUBS 0.201314f
C1102 VTAIL.t6 VSUBS 0.066882f
C1103 VTAIL.n237 VSUBS 0.023255f
C1104 VTAIL.n238 VSUBS 0.023325f
C1105 VTAIL.n239 VSUBS 0.013118f
C1106 VTAIL.n240 VSUBS 1.28719f
C1107 VTAIL.n241 VSUBS 0.024413f
C1108 VTAIL.n242 VSUBS 0.013118f
C1109 VTAIL.n243 VSUBS 0.01389f
C1110 VTAIL.n244 VSUBS 0.031007f
C1111 VTAIL.n245 VSUBS 0.031007f
C1112 VTAIL.n246 VSUBS 0.01389f
C1113 VTAIL.n247 VSUBS 0.013118f
C1114 VTAIL.n248 VSUBS 0.024413f
C1115 VTAIL.n249 VSUBS 0.024413f
C1116 VTAIL.n250 VSUBS 0.013118f
C1117 VTAIL.n251 VSUBS 0.01389f
C1118 VTAIL.n252 VSUBS 0.031007f
C1119 VTAIL.n253 VSUBS 0.031007f
C1120 VTAIL.n254 VSUBS 0.01389f
C1121 VTAIL.n255 VSUBS 0.013118f
C1122 VTAIL.n256 VSUBS 0.024413f
C1123 VTAIL.n257 VSUBS 0.024413f
C1124 VTAIL.n258 VSUBS 0.013118f
C1125 VTAIL.n259 VSUBS 0.013504f
C1126 VTAIL.n260 VSUBS 0.013504f
C1127 VTAIL.n261 VSUBS 0.031007f
C1128 VTAIL.n262 VSUBS 0.031007f
C1129 VTAIL.n263 VSUBS 0.01389f
C1130 VTAIL.n264 VSUBS 0.013118f
C1131 VTAIL.n265 VSUBS 0.024413f
C1132 VTAIL.n266 VSUBS 0.024413f
C1133 VTAIL.n267 VSUBS 0.013118f
C1134 VTAIL.n268 VSUBS 0.01389f
C1135 VTAIL.n269 VSUBS 0.031007f
C1136 VTAIL.n270 VSUBS 0.031007f
C1137 VTAIL.n271 VSUBS 0.01389f
C1138 VTAIL.n272 VSUBS 0.013118f
C1139 VTAIL.n273 VSUBS 0.024413f
C1140 VTAIL.n274 VSUBS 0.024413f
C1141 VTAIL.n275 VSUBS 0.013118f
C1142 VTAIL.n276 VSUBS 0.01389f
C1143 VTAIL.n277 VSUBS 0.031007f
C1144 VTAIL.n278 VSUBS 0.075422f
C1145 VTAIL.n279 VSUBS 0.01389f
C1146 VTAIL.n280 VSUBS 0.013118f
C1147 VTAIL.n281 VSUBS 0.055762f
C1148 VTAIL.n282 VSUBS 0.037924f
C1149 VTAIL.n283 VSUBS 1.54017f
C1150 VTAIL.t4 VSUBS 0.247318f
C1151 VTAIL.t3 VSUBS 0.247318f
C1152 VTAIL.n284 VSUBS 1.81162f
C1153 VTAIL.n285 VSUBS 0.889308f
C1154 VTAIL.n286 VSUBS 0.026929f
C1155 VTAIL.n287 VSUBS 0.024413f
C1156 VTAIL.n288 VSUBS 0.013118f
C1157 VTAIL.n289 VSUBS 0.031007f
C1158 VTAIL.n290 VSUBS 0.01389f
C1159 VTAIL.n291 VSUBS 0.024413f
C1160 VTAIL.n292 VSUBS 0.013118f
C1161 VTAIL.n293 VSUBS 0.031007f
C1162 VTAIL.n294 VSUBS 0.01389f
C1163 VTAIL.n295 VSUBS 0.024413f
C1164 VTAIL.n296 VSUBS 0.013118f
C1165 VTAIL.n297 VSUBS 0.031007f
C1166 VTAIL.n298 VSUBS 0.01389f
C1167 VTAIL.n299 VSUBS 0.024413f
C1168 VTAIL.n300 VSUBS 0.013118f
C1169 VTAIL.n301 VSUBS 0.031007f
C1170 VTAIL.n302 VSUBS 0.031007f
C1171 VTAIL.n303 VSUBS 0.01389f
C1172 VTAIL.n304 VSUBS 0.024413f
C1173 VTAIL.n305 VSUBS 0.013118f
C1174 VTAIL.n306 VSUBS 0.031007f
C1175 VTAIL.n307 VSUBS 0.01389f
C1176 VTAIL.n308 VSUBS 0.201314f
C1177 VTAIL.t5 VSUBS 0.066882f
C1178 VTAIL.n309 VSUBS 0.023255f
C1179 VTAIL.n310 VSUBS 0.023325f
C1180 VTAIL.n311 VSUBS 0.013118f
C1181 VTAIL.n312 VSUBS 1.28719f
C1182 VTAIL.n313 VSUBS 0.024413f
C1183 VTAIL.n314 VSUBS 0.013118f
C1184 VTAIL.n315 VSUBS 0.01389f
C1185 VTAIL.n316 VSUBS 0.031007f
C1186 VTAIL.n317 VSUBS 0.031007f
C1187 VTAIL.n318 VSUBS 0.01389f
C1188 VTAIL.n319 VSUBS 0.013118f
C1189 VTAIL.n320 VSUBS 0.024413f
C1190 VTAIL.n321 VSUBS 0.024413f
C1191 VTAIL.n322 VSUBS 0.013118f
C1192 VTAIL.n323 VSUBS 0.01389f
C1193 VTAIL.n324 VSUBS 0.031007f
C1194 VTAIL.n325 VSUBS 0.031007f
C1195 VTAIL.n326 VSUBS 0.01389f
C1196 VTAIL.n327 VSUBS 0.013118f
C1197 VTAIL.n328 VSUBS 0.024413f
C1198 VTAIL.n329 VSUBS 0.024413f
C1199 VTAIL.n330 VSUBS 0.013118f
C1200 VTAIL.n331 VSUBS 0.013504f
C1201 VTAIL.n332 VSUBS 0.013504f
C1202 VTAIL.n333 VSUBS 0.031007f
C1203 VTAIL.n334 VSUBS 0.031007f
C1204 VTAIL.n335 VSUBS 0.01389f
C1205 VTAIL.n336 VSUBS 0.013118f
C1206 VTAIL.n337 VSUBS 0.024413f
C1207 VTAIL.n338 VSUBS 0.024413f
C1208 VTAIL.n339 VSUBS 0.013118f
C1209 VTAIL.n340 VSUBS 0.01389f
C1210 VTAIL.n341 VSUBS 0.031007f
C1211 VTAIL.n342 VSUBS 0.031007f
C1212 VTAIL.n343 VSUBS 0.01389f
C1213 VTAIL.n344 VSUBS 0.013118f
C1214 VTAIL.n345 VSUBS 0.024413f
C1215 VTAIL.n346 VSUBS 0.024413f
C1216 VTAIL.n347 VSUBS 0.013118f
C1217 VTAIL.n348 VSUBS 0.01389f
C1218 VTAIL.n349 VSUBS 0.031007f
C1219 VTAIL.n350 VSUBS 0.075422f
C1220 VTAIL.n351 VSUBS 0.01389f
C1221 VTAIL.n352 VSUBS 0.013118f
C1222 VTAIL.n353 VSUBS 0.055762f
C1223 VTAIL.n354 VSUBS 0.037924f
C1224 VTAIL.n355 VSUBS 0.216792f
C1225 VTAIL.n356 VSUBS 0.026929f
C1226 VTAIL.n357 VSUBS 0.024413f
C1227 VTAIL.n358 VSUBS 0.013118f
C1228 VTAIL.n359 VSUBS 0.031007f
C1229 VTAIL.n360 VSUBS 0.01389f
C1230 VTAIL.n361 VSUBS 0.024413f
C1231 VTAIL.n362 VSUBS 0.013118f
C1232 VTAIL.n363 VSUBS 0.031007f
C1233 VTAIL.n364 VSUBS 0.01389f
C1234 VTAIL.n365 VSUBS 0.024413f
C1235 VTAIL.n366 VSUBS 0.013118f
C1236 VTAIL.n367 VSUBS 0.031007f
C1237 VTAIL.n368 VSUBS 0.01389f
C1238 VTAIL.n369 VSUBS 0.024413f
C1239 VTAIL.n370 VSUBS 0.013118f
C1240 VTAIL.n371 VSUBS 0.031007f
C1241 VTAIL.n372 VSUBS 0.031007f
C1242 VTAIL.n373 VSUBS 0.01389f
C1243 VTAIL.n374 VSUBS 0.024413f
C1244 VTAIL.n375 VSUBS 0.013118f
C1245 VTAIL.n376 VSUBS 0.031007f
C1246 VTAIL.n377 VSUBS 0.01389f
C1247 VTAIL.n378 VSUBS 0.201314f
C1248 VTAIL.t9 VSUBS 0.066882f
C1249 VTAIL.n379 VSUBS 0.023255f
C1250 VTAIL.n380 VSUBS 0.023325f
C1251 VTAIL.n381 VSUBS 0.013118f
C1252 VTAIL.n382 VSUBS 1.28719f
C1253 VTAIL.n383 VSUBS 0.024413f
C1254 VTAIL.n384 VSUBS 0.013118f
C1255 VTAIL.n385 VSUBS 0.01389f
C1256 VTAIL.n386 VSUBS 0.031007f
C1257 VTAIL.n387 VSUBS 0.031007f
C1258 VTAIL.n388 VSUBS 0.01389f
C1259 VTAIL.n389 VSUBS 0.013118f
C1260 VTAIL.n390 VSUBS 0.024413f
C1261 VTAIL.n391 VSUBS 0.024413f
C1262 VTAIL.n392 VSUBS 0.013118f
C1263 VTAIL.n393 VSUBS 0.01389f
C1264 VTAIL.n394 VSUBS 0.031007f
C1265 VTAIL.n395 VSUBS 0.031007f
C1266 VTAIL.n396 VSUBS 0.01389f
C1267 VTAIL.n397 VSUBS 0.013118f
C1268 VTAIL.n398 VSUBS 0.024413f
C1269 VTAIL.n399 VSUBS 0.024413f
C1270 VTAIL.n400 VSUBS 0.013118f
C1271 VTAIL.n401 VSUBS 0.013504f
C1272 VTAIL.n402 VSUBS 0.013504f
C1273 VTAIL.n403 VSUBS 0.031007f
C1274 VTAIL.n404 VSUBS 0.031007f
C1275 VTAIL.n405 VSUBS 0.01389f
C1276 VTAIL.n406 VSUBS 0.013118f
C1277 VTAIL.n407 VSUBS 0.024413f
C1278 VTAIL.n408 VSUBS 0.024413f
C1279 VTAIL.n409 VSUBS 0.013118f
C1280 VTAIL.n410 VSUBS 0.01389f
C1281 VTAIL.n411 VSUBS 0.031007f
C1282 VTAIL.n412 VSUBS 0.031007f
C1283 VTAIL.n413 VSUBS 0.01389f
C1284 VTAIL.n414 VSUBS 0.013118f
C1285 VTAIL.n415 VSUBS 0.024413f
C1286 VTAIL.n416 VSUBS 0.024413f
C1287 VTAIL.n417 VSUBS 0.013118f
C1288 VTAIL.n418 VSUBS 0.01389f
C1289 VTAIL.n419 VSUBS 0.031007f
C1290 VTAIL.n420 VSUBS 0.075422f
C1291 VTAIL.n421 VSUBS 0.01389f
C1292 VTAIL.n422 VSUBS 0.013118f
C1293 VTAIL.n423 VSUBS 0.055762f
C1294 VTAIL.n424 VSUBS 0.037924f
C1295 VTAIL.n425 VSUBS 0.216792f
C1296 VTAIL.t13 VSUBS 0.247318f
C1297 VTAIL.t14 VSUBS 0.247318f
C1298 VTAIL.n426 VSUBS 1.81162f
C1299 VTAIL.n427 VSUBS 0.889308f
C1300 VTAIL.n428 VSUBS 0.026929f
C1301 VTAIL.n429 VSUBS 0.024413f
C1302 VTAIL.n430 VSUBS 0.013118f
C1303 VTAIL.n431 VSUBS 0.031007f
C1304 VTAIL.n432 VSUBS 0.01389f
C1305 VTAIL.n433 VSUBS 0.024413f
C1306 VTAIL.n434 VSUBS 0.013118f
C1307 VTAIL.n435 VSUBS 0.031007f
C1308 VTAIL.n436 VSUBS 0.01389f
C1309 VTAIL.n437 VSUBS 0.024413f
C1310 VTAIL.n438 VSUBS 0.013118f
C1311 VTAIL.n439 VSUBS 0.031007f
C1312 VTAIL.n440 VSUBS 0.01389f
C1313 VTAIL.n441 VSUBS 0.024413f
C1314 VTAIL.n442 VSUBS 0.013118f
C1315 VTAIL.n443 VSUBS 0.031007f
C1316 VTAIL.n444 VSUBS 0.031007f
C1317 VTAIL.n445 VSUBS 0.01389f
C1318 VTAIL.n446 VSUBS 0.024413f
C1319 VTAIL.n447 VSUBS 0.013118f
C1320 VTAIL.n448 VSUBS 0.031007f
C1321 VTAIL.n449 VSUBS 0.01389f
C1322 VTAIL.n450 VSUBS 0.201314f
C1323 VTAIL.t10 VSUBS 0.066882f
C1324 VTAIL.n451 VSUBS 0.023255f
C1325 VTAIL.n452 VSUBS 0.023325f
C1326 VTAIL.n453 VSUBS 0.013118f
C1327 VTAIL.n454 VSUBS 1.28719f
C1328 VTAIL.n455 VSUBS 0.024413f
C1329 VTAIL.n456 VSUBS 0.013118f
C1330 VTAIL.n457 VSUBS 0.01389f
C1331 VTAIL.n458 VSUBS 0.031007f
C1332 VTAIL.n459 VSUBS 0.031007f
C1333 VTAIL.n460 VSUBS 0.01389f
C1334 VTAIL.n461 VSUBS 0.013118f
C1335 VTAIL.n462 VSUBS 0.024413f
C1336 VTAIL.n463 VSUBS 0.024413f
C1337 VTAIL.n464 VSUBS 0.013118f
C1338 VTAIL.n465 VSUBS 0.01389f
C1339 VTAIL.n466 VSUBS 0.031007f
C1340 VTAIL.n467 VSUBS 0.031007f
C1341 VTAIL.n468 VSUBS 0.01389f
C1342 VTAIL.n469 VSUBS 0.013118f
C1343 VTAIL.n470 VSUBS 0.024413f
C1344 VTAIL.n471 VSUBS 0.024413f
C1345 VTAIL.n472 VSUBS 0.013118f
C1346 VTAIL.n473 VSUBS 0.013504f
C1347 VTAIL.n474 VSUBS 0.013504f
C1348 VTAIL.n475 VSUBS 0.031007f
C1349 VTAIL.n476 VSUBS 0.031007f
C1350 VTAIL.n477 VSUBS 0.01389f
C1351 VTAIL.n478 VSUBS 0.013118f
C1352 VTAIL.n479 VSUBS 0.024413f
C1353 VTAIL.n480 VSUBS 0.024413f
C1354 VTAIL.n481 VSUBS 0.013118f
C1355 VTAIL.n482 VSUBS 0.01389f
C1356 VTAIL.n483 VSUBS 0.031007f
C1357 VTAIL.n484 VSUBS 0.031007f
C1358 VTAIL.n485 VSUBS 0.01389f
C1359 VTAIL.n486 VSUBS 0.013118f
C1360 VTAIL.n487 VSUBS 0.024413f
C1361 VTAIL.n488 VSUBS 0.024413f
C1362 VTAIL.n489 VSUBS 0.013118f
C1363 VTAIL.n490 VSUBS 0.01389f
C1364 VTAIL.n491 VSUBS 0.031007f
C1365 VTAIL.n492 VSUBS 0.075422f
C1366 VTAIL.n493 VSUBS 0.01389f
C1367 VTAIL.n494 VSUBS 0.013118f
C1368 VTAIL.n495 VSUBS 0.055762f
C1369 VTAIL.n496 VSUBS 0.037924f
C1370 VTAIL.n497 VSUBS 1.54017f
C1371 VTAIL.n498 VSUBS 0.026929f
C1372 VTAIL.n499 VSUBS 0.024413f
C1373 VTAIL.n500 VSUBS 0.013118f
C1374 VTAIL.n501 VSUBS 0.031007f
C1375 VTAIL.n502 VSUBS 0.01389f
C1376 VTAIL.n503 VSUBS 0.024413f
C1377 VTAIL.n504 VSUBS 0.013118f
C1378 VTAIL.n505 VSUBS 0.031007f
C1379 VTAIL.n506 VSUBS 0.01389f
C1380 VTAIL.n507 VSUBS 0.024413f
C1381 VTAIL.n508 VSUBS 0.013118f
C1382 VTAIL.n509 VSUBS 0.031007f
C1383 VTAIL.n510 VSUBS 0.01389f
C1384 VTAIL.n511 VSUBS 0.024413f
C1385 VTAIL.n512 VSUBS 0.013118f
C1386 VTAIL.n513 VSUBS 0.031007f
C1387 VTAIL.n514 VSUBS 0.01389f
C1388 VTAIL.n515 VSUBS 0.024413f
C1389 VTAIL.n516 VSUBS 0.013118f
C1390 VTAIL.n517 VSUBS 0.031007f
C1391 VTAIL.n518 VSUBS 0.01389f
C1392 VTAIL.n519 VSUBS 0.201314f
C1393 VTAIL.t0 VSUBS 0.066882f
C1394 VTAIL.n520 VSUBS 0.023255f
C1395 VTAIL.n521 VSUBS 0.023325f
C1396 VTAIL.n522 VSUBS 0.013118f
C1397 VTAIL.n523 VSUBS 1.28719f
C1398 VTAIL.n524 VSUBS 0.024413f
C1399 VTAIL.n525 VSUBS 0.013118f
C1400 VTAIL.n526 VSUBS 0.01389f
C1401 VTAIL.n527 VSUBS 0.031007f
C1402 VTAIL.n528 VSUBS 0.031007f
C1403 VTAIL.n529 VSUBS 0.01389f
C1404 VTAIL.n530 VSUBS 0.013118f
C1405 VTAIL.n531 VSUBS 0.024413f
C1406 VTAIL.n532 VSUBS 0.024413f
C1407 VTAIL.n533 VSUBS 0.013118f
C1408 VTAIL.n534 VSUBS 0.01389f
C1409 VTAIL.n535 VSUBS 0.031007f
C1410 VTAIL.n536 VSUBS 0.031007f
C1411 VTAIL.n537 VSUBS 0.031007f
C1412 VTAIL.n538 VSUBS 0.01389f
C1413 VTAIL.n539 VSUBS 0.013118f
C1414 VTAIL.n540 VSUBS 0.024413f
C1415 VTAIL.n541 VSUBS 0.024413f
C1416 VTAIL.n542 VSUBS 0.013118f
C1417 VTAIL.n543 VSUBS 0.013504f
C1418 VTAIL.n544 VSUBS 0.013504f
C1419 VTAIL.n545 VSUBS 0.031007f
C1420 VTAIL.n546 VSUBS 0.031007f
C1421 VTAIL.n547 VSUBS 0.01389f
C1422 VTAIL.n548 VSUBS 0.013118f
C1423 VTAIL.n549 VSUBS 0.024413f
C1424 VTAIL.n550 VSUBS 0.024413f
C1425 VTAIL.n551 VSUBS 0.013118f
C1426 VTAIL.n552 VSUBS 0.01389f
C1427 VTAIL.n553 VSUBS 0.031007f
C1428 VTAIL.n554 VSUBS 0.031007f
C1429 VTAIL.n555 VSUBS 0.01389f
C1430 VTAIL.n556 VSUBS 0.013118f
C1431 VTAIL.n557 VSUBS 0.024413f
C1432 VTAIL.n558 VSUBS 0.024413f
C1433 VTAIL.n559 VSUBS 0.013118f
C1434 VTAIL.n560 VSUBS 0.01389f
C1435 VTAIL.n561 VSUBS 0.031007f
C1436 VTAIL.n562 VSUBS 0.075422f
C1437 VTAIL.n563 VSUBS 0.01389f
C1438 VTAIL.n564 VSUBS 0.013118f
C1439 VTAIL.n565 VSUBS 0.055762f
C1440 VTAIL.n566 VSUBS 0.037924f
C1441 VTAIL.n567 VSUBS 1.53559f
C1442 VDD1.t3 VSUBS 0.251456f
C1443 VDD1.t2 VSUBS 0.251456f
C1444 VDD1.n0 VSUBS 1.99246f
C1445 VDD1.t0 VSUBS 0.251456f
C1446 VDD1.t6 VSUBS 0.251456f
C1447 VDD1.n1 VSUBS 1.99123f
C1448 VDD1.t1 VSUBS 0.251456f
C1449 VDD1.t7 VSUBS 0.251456f
C1450 VDD1.n2 VSUBS 1.99123f
C1451 VDD1.n3 VSUBS 3.55718f
C1452 VDD1.t4 VSUBS 0.251456f
C1453 VDD1.t5 VSUBS 0.251456f
C1454 VDD1.n4 VSUBS 1.98182f
C1455 VDD1.n5 VSUBS 3.09137f
C1456 VP.n0 VSUBS 0.033436f
C1457 VP.t6 VSUBS 2.36351f
C1458 VP.n1 VSUBS 0.038255f
C1459 VP.n2 VSUBS 0.033436f
C1460 VP.t2 VSUBS 2.36351f
C1461 VP.n3 VSUBS 0.066809f
C1462 VP.n4 VSUBS 0.033436f
C1463 VP.t7 VSUBS 2.36351f
C1464 VP.n5 VSUBS 0.83979f
C1465 VP.n6 VSUBS 0.033436f
C1466 VP.n7 VSUBS 0.064275f
C1467 VP.n8 VSUBS 0.033436f
C1468 VP.t4 VSUBS 2.36351f
C1469 VP.n9 VSUBS 0.038255f
C1470 VP.n10 VSUBS 0.033436f
C1471 VP.t0 VSUBS 2.36351f
C1472 VP.n11 VSUBS 0.066809f
C1473 VP.n12 VSUBS 0.033436f
C1474 VP.t1 VSUBS 2.36351f
C1475 VP.n13 VSUBS 0.916606f
C1476 VP.t5 VSUBS 2.53811f
C1477 VP.n14 VSUBS 0.925151f
C1478 VP.n15 VSUBS 0.251093f
C1479 VP.n16 VSUBS 0.04253f
C1480 VP.n17 VSUBS 0.066809f
C1481 VP.n18 VSUBS 0.027057f
C1482 VP.n19 VSUBS 0.033436f
C1483 VP.n20 VSUBS 0.033436f
C1484 VP.n21 VSUBS 0.033436f
C1485 VP.n22 VSUBS 0.04253f
C1486 VP.n23 VSUBS 0.83979f
C1487 VP.n24 VSUBS 0.051806f
C1488 VP.n25 VSUBS 0.058147f
C1489 VP.n26 VSUBS 0.033436f
C1490 VP.n27 VSUBS 0.033436f
C1491 VP.n28 VSUBS 0.033436f
C1492 VP.n29 VSUBS 0.064275f
C1493 VP.n30 VSUBS 0.033253f
C1494 VP.n31 VSUBS 0.924045f
C1495 VP.n32 VSUBS 1.75997f
C1496 VP.n33 VSUBS 1.78457f
C1497 VP.t3 VSUBS 2.36351f
C1498 VP.n34 VSUBS 0.924045f
C1499 VP.n35 VSUBS 0.033253f
C1500 VP.n36 VSUBS 0.033436f
C1501 VP.n37 VSUBS 0.033436f
C1502 VP.n38 VSUBS 0.033436f
C1503 VP.n39 VSUBS 0.038255f
C1504 VP.n40 VSUBS 0.058147f
C1505 VP.n41 VSUBS 0.051806f
C1506 VP.n42 VSUBS 0.033436f
C1507 VP.n43 VSUBS 0.033436f
C1508 VP.n44 VSUBS 0.04253f
C1509 VP.n45 VSUBS 0.066809f
C1510 VP.n46 VSUBS 0.027057f
C1511 VP.n47 VSUBS 0.033436f
C1512 VP.n48 VSUBS 0.033436f
C1513 VP.n49 VSUBS 0.033436f
C1514 VP.n50 VSUBS 0.04253f
C1515 VP.n51 VSUBS 0.83979f
C1516 VP.n52 VSUBS 0.051806f
C1517 VP.n53 VSUBS 0.058147f
C1518 VP.n54 VSUBS 0.033436f
C1519 VP.n55 VSUBS 0.033436f
C1520 VP.n56 VSUBS 0.033436f
C1521 VP.n57 VSUBS 0.064275f
C1522 VP.n58 VSUBS 0.033253f
C1523 VP.n59 VSUBS 0.924045f
C1524 VP.n60 VSUBS 0.037992f
.ends

