* NGSPICE file created from diff_pair_sample_0830.ext - technology: sky130A

.subckt diff_pair_sample_0830 VTAIL VN VP B VDD2 VDD1
X0 B.t11 B.t9 B.t10 w_n3242_n4542# sky130_fd_pr__pfet_01v8 ad=6.9693 pd=36.52 as=0 ps=0 w=17.87 l=2.51
X1 VTAIL.t11 VN.t0 VDD2.t4 w_n3242_n4542# sky130_fd_pr__pfet_01v8 ad=2.94855 pd=18.2 as=2.94855 ps=18.2 w=17.87 l=2.51
X2 VDD1.t5 VP.t0 VTAIL.t5 w_n3242_n4542# sky130_fd_pr__pfet_01v8 ad=2.94855 pd=18.2 as=6.9693 ps=36.52 w=17.87 l=2.51
X3 VDD1.t4 VP.t1 VTAIL.t3 w_n3242_n4542# sky130_fd_pr__pfet_01v8 ad=6.9693 pd=36.52 as=2.94855 ps=18.2 w=17.87 l=2.51
X4 VDD2.t3 VN.t1 VTAIL.t10 w_n3242_n4542# sky130_fd_pr__pfet_01v8 ad=2.94855 pd=18.2 as=6.9693 ps=36.52 w=17.87 l=2.51
X5 VTAIL.t4 VP.t2 VDD1.t3 w_n3242_n4542# sky130_fd_pr__pfet_01v8 ad=2.94855 pd=18.2 as=2.94855 ps=18.2 w=17.87 l=2.51
X6 VDD2.t2 VN.t2 VTAIL.t9 w_n3242_n4542# sky130_fd_pr__pfet_01v8 ad=2.94855 pd=18.2 as=6.9693 ps=36.52 w=17.87 l=2.51
X7 B.t8 B.t6 B.t7 w_n3242_n4542# sky130_fd_pr__pfet_01v8 ad=6.9693 pd=36.52 as=0 ps=0 w=17.87 l=2.51
X8 B.t5 B.t3 B.t4 w_n3242_n4542# sky130_fd_pr__pfet_01v8 ad=6.9693 pd=36.52 as=0 ps=0 w=17.87 l=2.51
X9 VDD2.t5 VN.t3 VTAIL.t8 w_n3242_n4542# sky130_fd_pr__pfet_01v8 ad=6.9693 pd=36.52 as=2.94855 ps=18.2 w=17.87 l=2.51
X10 VTAIL.t7 VN.t4 VDD2.t0 w_n3242_n4542# sky130_fd_pr__pfet_01v8 ad=2.94855 pd=18.2 as=2.94855 ps=18.2 w=17.87 l=2.51
X11 VDD1.t2 VP.t3 VTAIL.t1 w_n3242_n4542# sky130_fd_pr__pfet_01v8 ad=2.94855 pd=18.2 as=6.9693 ps=36.52 w=17.87 l=2.51
X12 VTAIL.t0 VP.t4 VDD1.t1 w_n3242_n4542# sky130_fd_pr__pfet_01v8 ad=2.94855 pd=18.2 as=2.94855 ps=18.2 w=17.87 l=2.51
X13 VDD2.t1 VN.t5 VTAIL.t6 w_n3242_n4542# sky130_fd_pr__pfet_01v8 ad=6.9693 pd=36.52 as=2.94855 ps=18.2 w=17.87 l=2.51
X14 B.t2 B.t0 B.t1 w_n3242_n4542# sky130_fd_pr__pfet_01v8 ad=6.9693 pd=36.52 as=0 ps=0 w=17.87 l=2.51
X15 VDD1.t0 VP.t5 VTAIL.t2 w_n3242_n4542# sky130_fd_pr__pfet_01v8 ad=6.9693 pd=36.52 as=2.94855 ps=18.2 w=17.87 l=2.51
R0 B.n472 B.n471 585
R1 B.n470 B.n133 585
R2 B.n469 B.n468 585
R3 B.n467 B.n134 585
R4 B.n466 B.n465 585
R5 B.n464 B.n135 585
R6 B.n463 B.n462 585
R7 B.n461 B.n136 585
R8 B.n460 B.n459 585
R9 B.n458 B.n137 585
R10 B.n457 B.n456 585
R11 B.n455 B.n138 585
R12 B.n454 B.n453 585
R13 B.n452 B.n139 585
R14 B.n451 B.n450 585
R15 B.n449 B.n140 585
R16 B.n448 B.n447 585
R17 B.n446 B.n141 585
R18 B.n445 B.n444 585
R19 B.n443 B.n142 585
R20 B.n442 B.n441 585
R21 B.n440 B.n143 585
R22 B.n439 B.n438 585
R23 B.n437 B.n144 585
R24 B.n436 B.n435 585
R25 B.n434 B.n145 585
R26 B.n433 B.n432 585
R27 B.n431 B.n146 585
R28 B.n430 B.n429 585
R29 B.n428 B.n147 585
R30 B.n427 B.n426 585
R31 B.n425 B.n148 585
R32 B.n424 B.n423 585
R33 B.n422 B.n149 585
R34 B.n421 B.n420 585
R35 B.n419 B.n150 585
R36 B.n418 B.n417 585
R37 B.n416 B.n151 585
R38 B.n415 B.n414 585
R39 B.n413 B.n152 585
R40 B.n412 B.n411 585
R41 B.n410 B.n153 585
R42 B.n409 B.n408 585
R43 B.n407 B.n154 585
R44 B.n406 B.n405 585
R45 B.n404 B.n155 585
R46 B.n403 B.n402 585
R47 B.n401 B.n156 585
R48 B.n400 B.n399 585
R49 B.n398 B.n157 585
R50 B.n397 B.n396 585
R51 B.n395 B.n158 585
R52 B.n394 B.n393 585
R53 B.n392 B.n159 585
R54 B.n391 B.n390 585
R55 B.n389 B.n160 585
R56 B.n388 B.n387 585
R57 B.n386 B.n161 585
R58 B.n385 B.n384 585
R59 B.n383 B.n382 585
R60 B.n381 B.n165 585
R61 B.n380 B.n379 585
R62 B.n378 B.n166 585
R63 B.n377 B.n376 585
R64 B.n375 B.n167 585
R65 B.n374 B.n373 585
R66 B.n372 B.n168 585
R67 B.n371 B.n370 585
R68 B.n368 B.n169 585
R69 B.n367 B.n366 585
R70 B.n365 B.n172 585
R71 B.n364 B.n363 585
R72 B.n362 B.n173 585
R73 B.n361 B.n360 585
R74 B.n359 B.n174 585
R75 B.n358 B.n357 585
R76 B.n356 B.n175 585
R77 B.n355 B.n354 585
R78 B.n353 B.n176 585
R79 B.n352 B.n351 585
R80 B.n350 B.n177 585
R81 B.n349 B.n348 585
R82 B.n347 B.n178 585
R83 B.n346 B.n345 585
R84 B.n344 B.n179 585
R85 B.n343 B.n342 585
R86 B.n341 B.n180 585
R87 B.n340 B.n339 585
R88 B.n338 B.n181 585
R89 B.n337 B.n336 585
R90 B.n335 B.n182 585
R91 B.n334 B.n333 585
R92 B.n332 B.n183 585
R93 B.n331 B.n330 585
R94 B.n329 B.n184 585
R95 B.n328 B.n327 585
R96 B.n326 B.n185 585
R97 B.n325 B.n324 585
R98 B.n323 B.n186 585
R99 B.n322 B.n321 585
R100 B.n320 B.n187 585
R101 B.n319 B.n318 585
R102 B.n317 B.n188 585
R103 B.n316 B.n315 585
R104 B.n314 B.n189 585
R105 B.n313 B.n312 585
R106 B.n311 B.n190 585
R107 B.n310 B.n309 585
R108 B.n308 B.n191 585
R109 B.n307 B.n306 585
R110 B.n305 B.n192 585
R111 B.n304 B.n303 585
R112 B.n302 B.n193 585
R113 B.n301 B.n300 585
R114 B.n299 B.n194 585
R115 B.n298 B.n297 585
R116 B.n296 B.n195 585
R117 B.n295 B.n294 585
R118 B.n293 B.n196 585
R119 B.n292 B.n291 585
R120 B.n290 B.n197 585
R121 B.n289 B.n288 585
R122 B.n287 B.n198 585
R123 B.n286 B.n285 585
R124 B.n284 B.n199 585
R125 B.n283 B.n282 585
R126 B.n281 B.n200 585
R127 B.n473 B.n132 585
R128 B.n475 B.n474 585
R129 B.n476 B.n131 585
R130 B.n478 B.n477 585
R131 B.n479 B.n130 585
R132 B.n481 B.n480 585
R133 B.n482 B.n129 585
R134 B.n484 B.n483 585
R135 B.n485 B.n128 585
R136 B.n487 B.n486 585
R137 B.n488 B.n127 585
R138 B.n490 B.n489 585
R139 B.n491 B.n126 585
R140 B.n493 B.n492 585
R141 B.n494 B.n125 585
R142 B.n496 B.n495 585
R143 B.n497 B.n124 585
R144 B.n499 B.n498 585
R145 B.n500 B.n123 585
R146 B.n502 B.n501 585
R147 B.n503 B.n122 585
R148 B.n505 B.n504 585
R149 B.n506 B.n121 585
R150 B.n508 B.n507 585
R151 B.n509 B.n120 585
R152 B.n511 B.n510 585
R153 B.n512 B.n119 585
R154 B.n514 B.n513 585
R155 B.n515 B.n118 585
R156 B.n517 B.n516 585
R157 B.n518 B.n117 585
R158 B.n520 B.n519 585
R159 B.n521 B.n116 585
R160 B.n523 B.n522 585
R161 B.n524 B.n115 585
R162 B.n526 B.n525 585
R163 B.n527 B.n114 585
R164 B.n529 B.n528 585
R165 B.n530 B.n113 585
R166 B.n532 B.n531 585
R167 B.n533 B.n112 585
R168 B.n535 B.n534 585
R169 B.n536 B.n111 585
R170 B.n538 B.n537 585
R171 B.n539 B.n110 585
R172 B.n541 B.n540 585
R173 B.n542 B.n109 585
R174 B.n544 B.n543 585
R175 B.n545 B.n108 585
R176 B.n547 B.n546 585
R177 B.n548 B.n107 585
R178 B.n550 B.n549 585
R179 B.n551 B.n106 585
R180 B.n553 B.n552 585
R181 B.n554 B.n105 585
R182 B.n556 B.n555 585
R183 B.n557 B.n104 585
R184 B.n559 B.n558 585
R185 B.n560 B.n103 585
R186 B.n562 B.n561 585
R187 B.n563 B.n102 585
R188 B.n565 B.n564 585
R189 B.n566 B.n101 585
R190 B.n568 B.n567 585
R191 B.n569 B.n100 585
R192 B.n571 B.n570 585
R193 B.n572 B.n99 585
R194 B.n574 B.n573 585
R195 B.n575 B.n98 585
R196 B.n577 B.n576 585
R197 B.n578 B.n97 585
R198 B.n580 B.n579 585
R199 B.n581 B.n96 585
R200 B.n583 B.n582 585
R201 B.n584 B.n95 585
R202 B.n586 B.n585 585
R203 B.n587 B.n94 585
R204 B.n589 B.n588 585
R205 B.n590 B.n93 585
R206 B.n592 B.n591 585
R207 B.n593 B.n92 585
R208 B.n595 B.n594 585
R209 B.n596 B.n91 585
R210 B.n598 B.n597 585
R211 B.n790 B.n789 585
R212 B.n788 B.n23 585
R213 B.n787 B.n786 585
R214 B.n785 B.n24 585
R215 B.n784 B.n783 585
R216 B.n782 B.n25 585
R217 B.n781 B.n780 585
R218 B.n779 B.n26 585
R219 B.n778 B.n777 585
R220 B.n776 B.n27 585
R221 B.n775 B.n774 585
R222 B.n773 B.n28 585
R223 B.n772 B.n771 585
R224 B.n770 B.n29 585
R225 B.n769 B.n768 585
R226 B.n767 B.n30 585
R227 B.n766 B.n765 585
R228 B.n764 B.n31 585
R229 B.n763 B.n762 585
R230 B.n761 B.n32 585
R231 B.n760 B.n759 585
R232 B.n758 B.n33 585
R233 B.n757 B.n756 585
R234 B.n755 B.n34 585
R235 B.n754 B.n753 585
R236 B.n752 B.n35 585
R237 B.n751 B.n750 585
R238 B.n749 B.n36 585
R239 B.n748 B.n747 585
R240 B.n746 B.n37 585
R241 B.n745 B.n744 585
R242 B.n743 B.n38 585
R243 B.n742 B.n741 585
R244 B.n740 B.n39 585
R245 B.n739 B.n738 585
R246 B.n737 B.n40 585
R247 B.n736 B.n735 585
R248 B.n734 B.n41 585
R249 B.n733 B.n732 585
R250 B.n731 B.n42 585
R251 B.n730 B.n729 585
R252 B.n728 B.n43 585
R253 B.n727 B.n726 585
R254 B.n725 B.n44 585
R255 B.n724 B.n723 585
R256 B.n722 B.n45 585
R257 B.n721 B.n720 585
R258 B.n719 B.n46 585
R259 B.n718 B.n717 585
R260 B.n716 B.n47 585
R261 B.n715 B.n714 585
R262 B.n713 B.n48 585
R263 B.n712 B.n711 585
R264 B.n710 B.n49 585
R265 B.n709 B.n708 585
R266 B.n707 B.n50 585
R267 B.n706 B.n705 585
R268 B.n704 B.n51 585
R269 B.n703 B.n702 585
R270 B.n701 B.n700 585
R271 B.n699 B.n55 585
R272 B.n698 B.n697 585
R273 B.n696 B.n56 585
R274 B.n695 B.n694 585
R275 B.n693 B.n57 585
R276 B.n692 B.n691 585
R277 B.n690 B.n58 585
R278 B.n689 B.n688 585
R279 B.n686 B.n59 585
R280 B.n685 B.n684 585
R281 B.n683 B.n62 585
R282 B.n682 B.n681 585
R283 B.n680 B.n63 585
R284 B.n679 B.n678 585
R285 B.n677 B.n64 585
R286 B.n676 B.n675 585
R287 B.n674 B.n65 585
R288 B.n673 B.n672 585
R289 B.n671 B.n66 585
R290 B.n670 B.n669 585
R291 B.n668 B.n67 585
R292 B.n667 B.n666 585
R293 B.n665 B.n68 585
R294 B.n664 B.n663 585
R295 B.n662 B.n69 585
R296 B.n661 B.n660 585
R297 B.n659 B.n70 585
R298 B.n658 B.n657 585
R299 B.n656 B.n71 585
R300 B.n655 B.n654 585
R301 B.n653 B.n72 585
R302 B.n652 B.n651 585
R303 B.n650 B.n73 585
R304 B.n649 B.n648 585
R305 B.n647 B.n74 585
R306 B.n646 B.n645 585
R307 B.n644 B.n75 585
R308 B.n643 B.n642 585
R309 B.n641 B.n76 585
R310 B.n640 B.n639 585
R311 B.n638 B.n77 585
R312 B.n637 B.n636 585
R313 B.n635 B.n78 585
R314 B.n634 B.n633 585
R315 B.n632 B.n79 585
R316 B.n631 B.n630 585
R317 B.n629 B.n80 585
R318 B.n628 B.n627 585
R319 B.n626 B.n81 585
R320 B.n625 B.n624 585
R321 B.n623 B.n82 585
R322 B.n622 B.n621 585
R323 B.n620 B.n83 585
R324 B.n619 B.n618 585
R325 B.n617 B.n84 585
R326 B.n616 B.n615 585
R327 B.n614 B.n85 585
R328 B.n613 B.n612 585
R329 B.n611 B.n86 585
R330 B.n610 B.n609 585
R331 B.n608 B.n87 585
R332 B.n607 B.n606 585
R333 B.n605 B.n88 585
R334 B.n604 B.n603 585
R335 B.n602 B.n89 585
R336 B.n601 B.n600 585
R337 B.n599 B.n90 585
R338 B.n791 B.n22 585
R339 B.n793 B.n792 585
R340 B.n794 B.n21 585
R341 B.n796 B.n795 585
R342 B.n797 B.n20 585
R343 B.n799 B.n798 585
R344 B.n800 B.n19 585
R345 B.n802 B.n801 585
R346 B.n803 B.n18 585
R347 B.n805 B.n804 585
R348 B.n806 B.n17 585
R349 B.n808 B.n807 585
R350 B.n809 B.n16 585
R351 B.n811 B.n810 585
R352 B.n812 B.n15 585
R353 B.n814 B.n813 585
R354 B.n815 B.n14 585
R355 B.n817 B.n816 585
R356 B.n818 B.n13 585
R357 B.n820 B.n819 585
R358 B.n821 B.n12 585
R359 B.n823 B.n822 585
R360 B.n824 B.n11 585
R361 B.n826 B.n825 585
R362 B.n827 B.n10 585
R363 B.n829 B.n828 585
R364 B.n830 B.n9 585
R365 B.n832 B.n831 585
R366 B.n833 B.n8 585
R367 B.n835 B.n834 585
R368 B.n836 B.n7 585
R369 B.n838 B.n837 585
R370 B.n839 B.n6 585
R371 B.n841 B.n840 585
R372 B.n842 B.n5 585
R373 B.n844 B.n843 585
R374 B.n845 B.n4 585
R375 B.n847 B.n846 585
R376 B.n848 B.n3 585
R377 B.n850 B.n849 585
R378 B.n851 B.n0 585
R379 B.n2 B.n1 585
R380 B.n221 B.n220 585
R381 B.n223 B.n222 585
R382 B.n224 B.n219 585
R383 B.n226 B.n225 585
R384 B.n227 B.n218 585
R385 B.n229 B.n228 585
R386 B.n230 B.n217 585
R387 B.n232 B.n231 585
R388 B.n233 B.n216 585
R389 B.n235 B.n234 585
R390 B.n236 B.n215 585
R391 B.n238 B.n237 585
R392 B.n239 B.n214 585
R393 B.n241 B.n240 585
R394 B.n242 B.n213 585
R395 B.n244 B.n243 585
R396 B.n245 B.n212 585
R397 B.n247 B.n246 585
R398 B.n248 B.n211 585
R399 B.n250 B.n249 585
R400 B.n251 B.n210 585
R401 B.n253 B.n252 585
R402 B.n254 B.n209 585
R403 B.n256 B.n255 585
R404 B.n257 B.n208 585
R405 B.n259 B.n258 585
R406 B.n260 B.n207 585
R407 B.n262 B.n261 585
R408 B.n263 B.n206 585
R409 B.n265 B.n264 585
R410 B.n266 B.n205 585
R411 B.n268 B.n267 585
R412 B.n269 B.n204 585
R413 B.n271 B.n270 585
R414 B.n272 B.n203 585
R415 B.n274 B.n273 585
R416 B.n275 B.n202 585
R417 B.n277 B.n276 585
R418 B.n278 B.n201 585
R419 B.n280 B.n279 585
R420 B.n281 B.n280 530.939
R421 B.n473 B.n472 530.939
R422 B.n599 B.n598 530.939
R423 B.n791 B.n790 530.939
R424 B.n170 B.t9 379.488
R425 B.n162 B.t0 379.488
R426 B.n60 B.t3 379.488
R427 B.n52 B.t6 379.488
R428 B.n853 B.n852 256.663
R429 B.n852 B.n851 235.042
R430 B.n852 B.n2 235.042
R431 B.n162 B.t1 164.981
R432 B.n60 B.t5 164.981
R433 B.n170 B.t10 164.958
R434 B.n52 B.t8 164.958
R435 B.n282 B.n281 163.367
R436 B.n282 B.n199 163.367
R437 B.n286 B.n199 163.367
R438 B.n287 B.n286 163.367
R439 B.n288 B.n287 163.367
R440 B.n288 B.n197 163.367
R441 B.n292 B.n197 163.367
R442 B.n293 B.n292 163.367
R443 B.n294 B.n293 163.367
R444 B.n294 B.n195 163.367
R445 B.n298 B.n195 163.367
R446 B.n299 B.n298 163.367
R447 B.n300 B.n299 163.367
R448 B.n300 B.n193 163.367
R449 B.n304 B.n193 163.367
R450 B.n305 B.n304 163.367
R451 B.n306 B.n305 163.367
R452 B.n306 B.n191 163.367
R453 B.n310 B.n191 163.367
R454 B.n311 B.n310 163.367
R455 B.n312 B.n311 163.367
R456 B.n312 B.n189 163.367
R457 B.n316 B.n189 163.367
R458 B.n317 B.n316 163.367
R459 B.n318 B.n317 163.367
R460 B.n318 B.n187 163.367
R461 B.n322 B.n187 163.367
R462 B.n323 B.n322 163.367
R463 B.n324 B.n323 163.367
R464 B.n324 B.n185 163.367
R465 B.n328 B.n185 163.367
R466 B.n329 B.n328 163.367
R467 B.n330 B.n329 163.367
R468 B.n330 B.n183 163.367
R469 B.n334 B.n183 163.367
R470 B.n335 B.n334 163.367
R471 B.n336 B.n335 163.367
R472 B.n336 B.n181 163.367
R473 B.n340 B.n181 163.367
R474 B.n341 B.n340 163.367
R475 B.n342 B.n341 163.367
R476 B.n342 B.n179 163.367
R477 B.n346 B.n179 163.367
R478 B.n347 B.n346 163.367
R479 B.n348 B.n347 163.367
R480 B.n348 B.n177 163.367
R481 B.n352 B.n177 163.367
R482 B.n353 B.n352 163.367
R483 B.n354 B.n353 163.367
R484 B.n354 B.n175 163.367
R485 B.n358 B.n175 163.367
R486 B.n359 B.n358 163.367
R487 B.n360 B.n359 163.367
R488 B.n360 B.n173 163.367
R489 B.n364 B.n173 163.367
R490 B.n365 B.n364 163.367
R491 B.n366 B.n365 163.367
R492 B.n366 B.n169 163.367
R493 B.n371 B.n169 163.367
R494 B.n372 B.n371 163.367
R495 B.n373 B.n372 163.367
R496 B.n373 B.n167 163.367
R497 B.n377 B.n167 163.367
R498 B.n378 B.n377 163.367
R499 B.n379 B.n378 163.367
R500 B.n379 B.n165 163.367
R501 B.n383 B.n165 163.367
R502 B.n384 B.n383 163.367
R503 B.n384 B.n161 163.367
R504 B.n388 B.n161 163.367
R505 B.n389 B.n388 163.367
R506 B.n390 B.n389 163.367
R507 B.n390 B.n159 163.367
R508 B.n394 B.n159 163.367
R509 B.n395 B.n394 163.367
R510 B.n396 B.n395 163.367
R511 B.n396 B.n157 163.367
R512 B.n400 B.n157 163.367
R513 B.n401 B.n400 163.367
R514 B.n402 B.n401 163.367
R515 B.n402 B.n155 163.367
R516 B.n406 B.n155 163.367
R517 B.n407 B.n406 163.367
R518 B.n408 B.n407 163.367
R519 B.n408 B.n153 163.367
R520 B.n412 B.n153 163.367
R521 B.n413 B.n412 163.367
R522 B.n414 B.n413 163.367
R523 B.n414 B.n151 163.367
R524 B.n418 B.n151 163.367
R525 B.n419 B.n418 163.367
R526 B.n420 B.n419 163.367
R527 B.n420 B.n149 163.367
R528 B.n424 B.n149 163.367
R529 B.n425 B.n424 163.367
R530 B.n426 B.n425 163.367
R531 B.n426 B.n147 163.367
R532 B.n430 B.n147 163.367
R533 B.n431 B.n430 163.367
R534 B.n432 B.n431 163.367
R535 B.n432 B.n145 163.367
R536 B.n436 B.n145 163.367
R537 B.n437 B.n436 163.367
R538 B.n438 B.n437 163.367
R539 B.n438 B.n143 163.367
R540 B.n442 B.n143 163.367
R541 B.n443 B.n442 163.367
R542 B.n444 B.n443 163.367
R543 B.n444 B.n141 163.367
R544 B.n448 B.n141 163.367
R545 B.n449 B.n448 163.367
R546 B.n450 B.n449 163.367
R547 B.n450 B.n139 163.367
R548 B.n454 B.n139 163.367
R549 B.n455 B.n454 163.367
R550 B.n456 B.n455 163.367
R551 B.n456 B.n137 163.367
R552 B.n460 B.n137 163.367
R553 B.n461 B.n460 163.367
R554 B.n462 B.n461 163.367
R555 B.n462 B.n135 163.367
R556 B.n466 B.n135 163.367
R557 B.n467 B.n466 163.367
R558 B.n468 B.n467 163.367
R559 B.n468 B.n133 163.367
R560 B.n472 B.n133 163.367
R561 B.n598 B.n91 163.367
R562 B.n594 B.n91 163.367
R563 B.n594 B.n593 163.367
R564 B.n593 B.n592 163.367
R565 B.n592 B.n93 163.367
R566 B.n588 B.n93 163.367
R567 B.n588 B.n587 163.367
R568 B.n587 B.n586 163.367
R569 B.n586 B.n95 163.367
R570 B.n582 B.n95 163.367
R571 B.n582 B.n581 163.367
R572 B.n581 B.n580 163.367
R573 B.n580 B.n97 163.367
R574 B.n576 B.n97 163.367
R575 B.n576 B.n575 163.367
R576 B.n575 B.n574 163.367
R577 B.n574 B.n99 163.367
R578 B.n570 B.n99 163.367
R579 B.n570 B.n569 163.367
R580 B.n569 B.n568 163.367
R581 B.n568 B.n101 163.367
R582 B.n564 B.n101 163.367
R583 B.n564 B.n563 163.367
R584 B.n563 B.n562 163.367
R585 B.n562 B.n103 163.367
R586 B.n558 B.n103 163.367
R587 B.n558 B.n557 163.367
R588 B.n557 B.n556 163.367
R589 B.n556 B.n105 163.367
R590 B.n552 B.n105 163.367
R591 B.n552 B.n551 163.367
R592 B.n551 B.n550 163.367
R593 B.n550 B.n107 163.367
R594 B.n546 B.n107 163.367
R595 B.n546 B.n545 163.367
R596 B.n545 B.n544 163.367
R597 B.n544 B.n109 163.367
R598 B.n540 B.n109 163.367
R599 B.n540 B.n539 163.367
R600 B.n539 B.n538 163.367
R601 B.n538 B.n111 163.367
R602 B.n534 B.n111 163.367
R603 B.n534 B.n533 163.367
R604 B.n533 B.n532 163.367
R605 B.n532 B.n113 163.367
R606 B.n528 B.n113 163.367
R607 B.n528 B.n527 163.367
R608 B.n527 B.n526 163.367
R609 B.n526 B.n115 163.367
R610 B.n522 B.n115 163.367
R611 B.n522 B.n521 163.367
R612 B.n521 B.n520 163.367
R613 B.n520 B.n117 163.367
R614 B.n516 B.n117 163.367
R615 B.n516 B.n515 163.367
R616 B.n515 B.n514 163.367
R617 B.n514 B.n119 163.367
R618 B.n510 B.n119 163.367
R619 B.n510 B.n509 163.367
R620 B.n509 B.n508 163.367
R621 B.n508 B.n121 163.367
R622 B.n504 B.n121 163.367
R623 B.n504 B.n503 163.367
R624 B.n503 B.n502 163.367
R625 B.n502 B.n123 163.367
R626 B.n498 B.n123 163.367
R627 B.n498 B.n497 163.367
R628 B.n497 B.n496 163.367
R629 B.n496 B.n125 163.367
R630 B.n492 B.n125 163.367
R631 B.n492 B.n491 163.367
R632 B.n491 B.n490 163.367
R633 B.n490 B.n127 163.367
R634 B.n486 B.n127 163.367
R635 B.n486 B.n485 163.367
R636 B.n485 B.n484 163.367
R637 B.n484 B.n129 163.367
R638 B.n480 B.n129 163.367
R639 B.n480 B.n479 163.367
R640 B.n479 B.n478 163.367
R641 B.n478 B.n131 163.367
R642 B.n474 B.n131 163.367
R643 B.n474 B.n473 163.367
R644 B.n790 B.n23 163.367
R645 B.n786 B.n23 163.367
R646 B.n786 B.n785 163.367
R647 B.n785 B.n784 163.367
R648 B.n784 B.n25 163.367
R649 B.n780 B.n25 163.367
R650 B.n780 B.n779 163.367
R651 B.n779 B.n778 163.367
R652 B.n778 B.n27 163.367
R653 B.n774 B.n27 163.367
R654 B.n774 B.n773 163.367
R655 B.n773 B.n772 163.367
R656 B.n772 B.n29 163.367
R657 B.n768 B.n29 163.367
R658 B.n768 B.n767 163.367
R659 B.n767 B.n766 163.367
R660 B.n766 B.n31 163.367
R661 B.n762 B.n31 163.367
R662 B.n762 B.n761 163.367
R663 B.n761 B.n760 163.367
R664 B.n760 B.n33 163.367
R665 B.n756 B.n33 163.367
R666 B.n756 B.n755 163.367
R667 B.n755 B.n754 163.367
R668 B.n754 B.n35 163.367
R669 B.n750 B.n35 163.367
R670 B.n750 B.n749 163.367
R671 B.n749 B.n748 163.367
R672 B.n748 B.n37 163.367
R673 B.n744 B.n37 163.367
R674 B.n744 B.n743 163.367
R675 B.n743 B.n742 163.367
R676 B.n742 B.n39 163.367
R677 B.n738 B.n39 163.367
R678 B.n738 B.n737 163.367
R679 B.n737 B.n736 163.367
R680 B.n736 B.n41 163.367
R681 B.n732 B.n41 163.367
R682 B.n732 B.n731 163.367
R683 B.n731 B.n730 163.367
R684 B.n730 B.n43 163.367
R685 B.n726 B.n43 163.367
R686 B.n726 B.n725 163.367
R687 B.n725 B.n724 163.367
R688 B.n724 B.n45 163.367
R689 B.n720 B.n45 163.367
R690 B.n720 B.n719 163.367
R691 B.n719 B.n718 163.367
R692 B.n718 B.n47 163.367
R693 B.n714 B.n47 163.367
R694 B.n714 B.n713 163.367
R695 B.n713 B.n712 163.367
R696 B.n712 B.n49 163.367
R697 B.n708 B.n49 163.367
R698 B.n708 B.n707 163.367
R699 B.n707 B.n706 163.367
R700 B.n706 B.n51 163.367
R701 B.n702 B.n51 163.367
R702 B.n702 B.n701 163.367
R703 B.n701 B.n55 163.367
R704 B.n697 B.n55 163.367
R705 B.n697 B.n696 163.367
R706 B.n696 B.n695 163.367
R707 B.n695 B.n57 163.367
R708 B.n691 B.n57 163.367
R709 B.n691 B.n690 163.367
R710 B.n690 B.n689 163.367
R711 B.n689 B.n59 163.367
R712 B.n684 B.n59 163.367
R713 B.n684 B.n683 163.367
R714 B.n683 B.n682 163.367
R715 B.n682 B.n63 163.367
R716 B.n678 B.n63 163.367
R717 B.n678 B.n677 163.367
R718 B.n677 B.n676 163.367
R719 B.n676 B.n65 163.367
R720 B.n672 B.n65 163.367
R721 B.n672 B.n671 163.367
R722 B.n671 B.n670 163.367
R723 B.n670 B.n67 163.367
R724 B.n666 B.n67 163.367
R725 B.n666 B.n665 163.367
R726 B.n665 B.n664 163.367
R727 B.n664 B.n69 163.367
R728 B.n660 B.n69 163.367
R729 B.n660 B.n659 163.367
R730 B.n659 B.n658 163.367
R731 B.n658 B.n71 163.367
R732 B.n654 B.n71 163.367
R733 B.n654 B.n653 163.367
R734 B.n653 B.n652 163.367
R735 B.n652 B.n73 163.367
R736 B.n648 B.n73 163.367
R737 B.n648 B.n647 163.367
R738 B.n647 B.n646 163.367
R739 B.n646 B.n75 163.367
R740 B.n642 B.n75 163.367
R741 B.n642 B.n641 163.367
R742 B.n641 B.n640 163.367
R743 B.n640 B.n77 163.367
R744 B.n636 B.n77 163.367
R745 B.n636 B.n635 163.367
R746 B.n635 B.n634 163.367
R747 B.n634 B.n79 163.367
R748 B.n630 B.n79 163.367
R749 B.n630 B.n629 163.367
R750 B.n629 B.n628 163.367
R751 B.n628 B.n81 163.367
R752 B.n624 B.n81 163.367
R753 B.n624 B.n623 163.367
R754 B.n623 B.n622 163.367
R755 B.n622 B.n83 163.367
R756 B.n618 B.n83 163.367
R757 B.n618 B.n617 163.367
R758 B.n617 B.n616 163.367
R759 B.n616 B.n85 163.367
R760 B.n612 B.n85 163.367
R761 B.n612 B.n611 163.367
R762 B.n611 B.n610 163.367
R763 B.n610 B.n87 163.367
R764 B.n606 B.n87 163.367
R765 B.n606 B.n605 163.367
R766 B.n605 B.n604 163.367
R767 B.n604 B.n89 163.367
R768 B.n600 B.n89 163.367
R769 B.n600 B.n599 163.367
R770 B.n792 B.n791 163.367
R771 B.n792 B.n21 163.367
R772 B.n796 B.n21 163.367
R773 B.n797 B.n796 163.367
R774 B.n798 B.n797 163.367
R775 B.n798 B.n19 163.367
R776 B.n802 B.n19 163.367
R777 B.n803 B.n802 163.367
R778 B.n804 B.n803 163.367
R779 B.n804 B.n17 163.367
R780 B.n808 B.n17 163.367
R781 B.n809 B.n808 163.367
R782 B.n810 B.n809 163.367
R783 B.n810 B.n15 163.367
R784 B.n814 B.n15 163.367
R785 B.n815 B.n814 163.367
R786 B.n816 B.n815 163.367
R787 B.n816 B.n13 163.367
R788 B.n820 B.n13 163.367
R789 B.n821 B.n820 163.367
R790 B.n822 B.n821 163.367
R791 B.n822 B.n11 163.367
R792 B.n826 B.n11 163.367
R793 B.n827 B.n826 163.367
R794 B.n828 B.n827 163.367
R795 B.n828 B.n9 163.367
R796 B.n832 B.n9 163.367
R797 B.n833 B.n832 163.367
R798 B.n834 B.n833 163.367
R799 B.n834 B.n7 163.367
R800 B.n838 B.n7 163.367
R801 B.n839 B.n838 163.367
R802 B.n840 B.n839 163.367
R803 B.n840 B.n5 163.367
R804 B.n844 B.n5 163.367
R805 B.n845 B.n844 163.367
R806 B.n846 B.n845 163.367
R807 B.n846 B.n3 163.367
R808 B.n850 B.n3 163.367
R809 B.n851 B.n850 163.367
R810 B.n221 B.n2 163.367
R811 B.n222 B.n221 163.367
R812 B.n222 B.n219 163.367
R813 B.n226 B.n219 163.367
R814 B.n227 B.n226 163.367
R815 B.n228 B.n227 163.367
R816 B.n228 B.n217 163.367
R817 B.n232 B.n217 163.367
R818 B.n233 B.n232 163.367
R819 B.n234 B.n233 163.367
R820 B.n234 B.n215 163.367
R821 B.n238 B.n215 163.367
R822 B.n239 B.n238 163.367
R823 B.n240 B.n239 163.367
R824 B.n240 B.n213 163.367
R825 B.n244 B.n213 163.367
R826 B.n245 B.n244 163.367
R827 B.n246 B.n245 163.367
R828 B.n246 B.n211 163.367
R829 B.n250 B.n211 163.367
R830 B.n251 B.n250 163.367
R831 B.n252 B.n251 163.367
R832 B.n252 B.n209 163.367
R833 B.n256 B.n209 163.367
R834 B.n257 B.n256 163.367
R835 B.n258 B.n257 163.367
R836 B.n258 B.n207 163.367
R837 B.n262 B.n207 163.367
R838 B.n263 B.n262 163.367
R839 B.n264 B.n263 163.367
R840 B.n264 B.n205 163.367
R841 B.n268 B.n205 163.367
R842 B.n269 B.n268 163.367
R843 B.n270 B.n269 163.367
R844 B.n270 B.n203 163.367
R845 B.n274 B.n203 163.367
R846 B.n275 B.n274 163.367
R847 B.n276 B.n275 163.367
R848 B.n276 B.n201 163.367
R849 B.n280 B.n201 163.367
R850 B.n163 B.t2 109.901
R851 B.n61 B.t4 109.901
R852 B.n171 B.t11 109.879
R853 B.n53 B.t7 109.879
R854 B.n369 B.n171 59.5399
R855 B.n164 B.n163 59.5399
R856 B.n687 B.n61 59.5399
R857 B.n54 B.n53 59.5399
R858 B.n171 B.n170 55.0793
R859 B.n163 B.n162 55.0793
R860 B.n61 B.n60 55.0793
R861 B.n53 B.n52 55.0793
R862 B.n789 B.n22 34.4981
R863 B.n597 B.n90 34.4981
R864 B.n471 B.n132 34.4981
R865 B.n279 B.n200 34.4981
R866 B B.n853 18.0485
R867 B.n793 B.n22 10.6151
R868 B.n794 B.n793 10.6151
R869 B.n795 B.n794 10.6151
R870 B.n795 B.n20 10.6151
R871 B.n799 B.n20 10.6151
R872 B.n800 B.n799 10.6151
R873 B.n801 B.n800 10.6151
R874 B.n801 B.n18 10.6151
R875 B.n805 B.n18 10.6151
R876 B.n806 B.n805 10.6151
R877 B.n807 B.n806 10.6151
R878 B.n807 B.n16 10.6151
R879 B.n811 B.n16 10.6151
R880 B.n812 B.n811 10.6151
R881 B.n813 B.n812 10.6151
R882 B.n813 B.n14 10.6151
R883 B.n817 B.n14 10.6151
R884 B.n818 B.n817 10.6151
R885 B.n819 B.n818 10.6151
R886 B.n819 B.n12 10.6151
R887 B.n823 B.n12 10.6151
R888 B.n824 B.n823 10.6151
R889 B.n825 B.n824 10.6151
R890 B.n825 B.n10 10.6151
R891 B.n829 B.n10 10.6151
R892 B.n830 B.n829 10.6151
R893 B.n831 B.n830 10.6151
R894 B.n831 B.n8 10.6151
R895 B.n835 B.n8 10.6151
R896 B.n836 B.n835 10.6151
R897 B.n837 B.n836 10.6151
R898 B.n837 B.n6 10.6151
R899 B.n841 B.n6 10.6151
R900 B.n842 B.n841 10.6151
R901 B.n843 B.n842 10.6151
R902 B.n843 B.n4 10.6151
R903 B.n847 B.n4 10.6151
R904 B.n848 B.n847 10.6151
R905 B.n849 B.n848 10.6151
R906 B.n849 B.n0 10.6151
R907 B.n789 B.n788 10.6151
R908 B.n788 B.n787 10.6151
R909 B.n787 B.n24 10.6151
R910 B.n783 B.n24 10.6151
R911 B.n783 B.n782 10.6151
R912 B.n782 B.n781 10.6151
R913 B.n781 B.n26 10.6151
R914 B.n777 B.n26 10.6151
R915 B.n777 B.n776 10.6151
R916 B.n776 B.n775 10.6151
R917 B.n775 B.n28 10.6151
R918 B.n771 B.n28 10.6151
R919 B.n771 B.n770 10.6151
R920 B.n770 B.n769 10.6151
R921 B.n769 B.n30 10.6151
R922 B.n765 B.n30 10.6151
R923 B.n765 B.n764 10.6151
R924 B.n764 B.n763 10.6151
R925 B.n763 B.n32 10.6151
R926 B.n759 B.n32 10.6151
R927 B.n759 B.n758 10.6151
R928 B.n758 B.n757 10.6151
R929 B.n757 B.n34 10.6151
R930 B.n753 B.n34 10.6151
R931 B.n753 B.n752 10.6151
R932 B.n752 B.n751 10.6151
R933 B.n751 B.n36 10.6151
R934 B.n747 B.n36 10.6151
R935 B.n747 B.n746 10.6151
R936 B.n746 B.n745 10.6151
R937 B.n745 B.n38 10.6151
R938 B.n741 B.n38 10.6151
R939 B.n741 B.n740 10.6151
R940 B.n740 B.n739 10.6151
R941 B.n739 B.n40 10.6151
R942 B.n735 B.n40 10.6151
R943 B.n735 B.n734 10.6151
R944 B.n734 B.n733 10.6151
R945 B.n733 B.n42 10.6151
R946 B.n729 B.n42 10.6151
R947 B.n729 B.n728 10.6151
R948 B.n728 B.n727 10.6151
R949 B.n727 B.n44 10.6151
R950 B.n723 B.n44 10.6151
R951 B.n723 B.n722 10.6151
R952 B.n722 B.n721 10.6151
R953 B.n721 B.n46 10.6151
R954 B.n717 B.n46 10.6151
R955 B.n717 B.n716 10.6151
R956 B.n716 B.n715 10.6151
R957 B.n715 B.n48 10.6151
R958 B.n711 B.n48 10.6151
R959 B.n711 B.n710 10.6151
R960 B.n710 B.n709 10.6151
R961 B.n709 B.n50 10.6151
R962 B.n705 B.n50 10.6151
R963 B.n705 B.n704 10.6151
R964 B.n704 B.n703 10.6151
R965 B.n700 B.n699 10.6151
R966 B.n699 B.n698 10.6151
R967 B.n698 B.n56 10.6151
R968 B.n694 B.n56 10.6151
R969 B.n694 B.n693 10.6151
R970 B.n693 B.n692 10.6151
R971 B.n692 B.n58 10.6151
R972 B.n688 B.n58 10.6151
R973 B.n686 B.n685 10.6151
R974 B.n685 B.n62 10.6151
R975 B.n681 B.n62 10.6151
R976 B.n681 B.n680 10.6151
R977 B.n680 B.n679 10.6151
R978 B.n679 B.n64 10.6151
R979 B.n675 B.n64 10.6151
R980 B.n675 B.n674 10.6151
R981 B.n674 B.n673 10.6151
R982 B.n673 B.n66 10.6151
R983 B.n669 B.n66 10.6151
R984 B.n669 B.n668 10.6151
R985 B.n668 B.n667 10.6151
R986 B.n667 B.n68 10.6151
R987 B.n663 B.n68 10.6151
R988 B.n663 B.n662 10.6151
R989 B.n662 B.n661 10.6151
R990 B.n661 B.n70 10.6151
R991 B.n657 B.n70 10.6151
R992 B.n657 B.n656 10.6151
R993 B.n656 B.n655 10.6151
R994 B.n655 B.n72 10.6151
R995 B.n651 B.n72 10.6151
R996 B.n651 B.n650 10.6151
R997 B.n650 B.n649 10.6151
R998 B.n649 B.n74 10.6151
R999 B.n645 B.n74 10.6151
R1000 B.n645 B.n644 10.6151
R1001 B.n644 B.n643 10.6151
R1002 B.n643 B.n76 10.6151
R1003 B.n639 B.n76 10.6151
R1004 B.n639 B.n638 10.6151
R1005 B.n638 B.n637 10.6151
R1006 B.n637 B.n78 10.6151
R1007 B.n633 B.n78 10.6151
R1008 B.n633 B.n632 10.6151
R1009 B.n632 B.n631 10.6151
R1010 B.n631 B.n80 10.6151
R1011 B.n627 B.n80 10.6151
R1012 B.n627 B.n626 10.6151
R1013 B.n626 B.n625 10.6151
R1014 B.n625 B.n82 10.6151
R1015 B.n621 B.n82 10.6151
R1016 B.n621 B.n620 10.6151
R1017 B.n620 B.n619 10.6151
R1018 B.n619 B.n84 10.6151
R1019 B.n615 B.n84 10.6151
R1020 B.n615 B.n614 10.6151
R1021 B.n614 B.n613 10.6151
R1022 B.n613 B.n86 10.6151
R1023 B.n609 B.n86 10.6151
R1024 B.n609 B.n608 10.6151
R1025 B.n608 B.n607 10.6151
R1026 B.n607 B.n88 10.6151
R1027 B.n603 B.n88 10.6151
R1028 B.n603 B.n602 10.6151
R1029 B.n602 B.n601 10.6151
R1030 B.n601 B.n90 10.6151
R1031 B.n597 B.n596 10.6151
R1032 B.n596 B.n595 10.6151
R1033 B.n595 B.n92 10.6151
R1034 B.n591 B.n92 10.6151
R1035 B.n591 B.n590 10.6151
R1036 B.n590 B.n589 10.6151
R1037 B.n589 B.n94 10.6151
R1038 B.n585 B.n94 10.6151
R1039 B.n585 B.n584 10.6151
R1040 B.n584 B.n583 10.6151
R1041 B.n583 B.n96 10.6151
R1042 B.n579 B.n96 10.6151
R1043 B.n579 B.n578 10.6151
R1044 B.n578 B.n577 10.6151
R1045 B.n577 B.n98 10.6151
R1046 B.n573 B.n98 10.6151
R1047 B.n573 B.n572 10.6151
R1048 B.n572 B.n571 10.6151
R1049 B.n571 B.n100 10.6151
R1050 B.n567 B.n100 10.6151
R1051 B.n567 B.n566 10.6151
R1052 B.n566 B.n565 10.6151
R1053 B.n565 B.n102 10.6151
R1054 B.n561 B.n102 10.6151
R1055 B.n561 B.n560 10.6151
R1056 B.n560 B.n559 10.6151
R1057 B.n559 B.n104 10.6151
R1058 B.n555 B.n104 10.6151
R1059 B.n555 B.n554 10.6151
R1060 B.n554 B.n553 10.6151
R1061 B.n553 B.n106 10.6151
R1062 B.n549 B.n106 10.6151
R1063 B.n549 B.n548 10.6151
R1064 B.n548 B.n547 10.6151
R1065 B.n547 B.n108 10.6151
R1066 B.n543 B.n108 10.6151
R1067 B.n543 B.n542 10.6151
R1068 B.n542 B.n541 10.6151
R1069 B.n541 B.n110 10.6151
R1070 B.n537 B.n110 10.6151
R1071 B.n537 B.n536 10.6151
R1072 B.n536 B.n535 10.6151
R1073 B.n535 B.n112 10.6151
R1074 B.n531 B.n112 10.6151
R1075 B.n531 B.n530 10.6151
R1076 B.n530 B.n529 10.6151
R1077 B.n529 B.n114 10.6151
R1078 B.n525 B.n114 10.6151
R1079 B.n525 B.n524 10.6151
R1080 B.n524 B.n523 10.6151
R1081 B.n523 B.n116 10.6151
R1082 B.n519 B.n116 10.6151
R1083 B.n519 B.n518 10.6151
R1084 B.n518 B.n517 10.6151
R1085 B.n517 B.n118 10.6151
R1086 B.n513 B.n118 10.6151
R1087 B.n513 B.n512 10.6151
R1088 B.n512 B.n511 10.6151
R1089 B.n511 B.n120 10.6151
R1090 B.n507 B.n120 10.6151
R1091 B.n507 B.n506 10.6151
R1092 B.n506 B.n505 10.6151
R1093 B.n505 B.n122 10.6151
R1094 B.n501 B.n122 10.6151
R1095 B.n501 B.n500 10.6151
R1096 B.n500 B.n499 10.6151
R1097 B.n499 B.n124 10.6151
R1098 B.n495 B.n124 10.6151
R1099 B.n495 B.n494 10.6151
R1100 B.n494 B.n493 10.6151
R1101 B.n493 B.n126 10.6151
R1102 B.n489 B.n126 10.6151
R1103 B.n489 B.n488 10.6151
R1104 B.n488 B.n487 10.6151
R1105 B.n487 B.n128 10.6151
R1106 B.n483 B.n128 10.6151
R1107 B.n483 B.n482 10.6151
R1108 B.n482 B.n481 10.6151
R1109 B.n481 B.n130 10.6151
R1110 B.n477 B.n130 10.6151
R1111 B.n477 B.n476 10.6151
R1112 B.n476 B.n475 10.6151
R1113 B.n475 B.n132 10.6151
R1114 B.n220 B.n1 10.6151
R1115 B.n223 B.n220 10.6151
R1116 B.n224 B.n223 10.6151
R1117 B.n225 B.n224 10.6151
R1118 B.n225 B.n218 10.6151
R1119 B.n229 B.n218 10.6151
R1120 B.n230 B.n229 10.6151
R1121 B.n231 B.n230 10.6151
R1122 B.n231 B.n216 10.6151
R1123 B.n235 B.n216 10.6151
R1124 B.n236 B.n235 10.6151
R1125 B.n237 B.n236 10.6151
R1126 B.n237 B.n214 10.6151
R1127 B.n241 B.n214 10.6151
R1128 B.n242 B.n241 10.6151
R1129 B.n243 B.n242 10.6151
R1130 B.n243 B.n212 10.6151
R1131 B.n247 B.n212 10.6151
R1132 B.n248 B.n247 10.6151
R1133 B.n249 B.n248 10.6151
R1134 B.n249 B.n210 10.6151
R1135 B.n253 B.n210 10.6151
R1136 B.n254 B.n253 10.6151
R1137 B.n255 B.n254 10.6151
R1138 B.n255 B.n208 10.6151
R1139 B.n259 B.n208 10.6151
R1140 B.n260 B.n259 10.6151
R1141 B.n261 B.n260 10.6151
R1142 B.n261 B.n206 10.6151
R1143 B.n265 B.n206 10.6151
R1144 B.n266 B.n265 10.6151
R1145 B.n267 B.n266 10.6151
R1146 B.n267 B.n204 10.6151
R1147 B.n271 B.n204 10.6151
R1148 B.n272 B.n271 10.6151
R1149 B.n273 B.n272 10.6151
R1150 B.n273 B.n202 10.6151
R1151 B.n277 B.n202 10.6151
R1152 B.n278 B.n277 10.6151
R1153 B.n279 B.n278 10.6151
R1154 B.n283 B.n200 10.6151
R1155 B.n284 B.n283 10.6151
R1156 B.n285 B.n284 10.6151
R1157 B.n285 B.n198 10.6151
R1158 B.n289 B.n198 10.6151
R1159 B.n290 B.n289 10.6151
R1160 B.n291 B.n290 10.6151
R1161 B.n291 B.n196 10.6151
R1162 B.n295 B.n196 10.6151
R1163 B.n296 B.n295 10.6151
R1164 B.n297 B.n296 10.6151
R1165 B.n297 B.n194 10.6151
R1166 B.n301 B.n194 10.6151
R1167 B.n302 B.n301 10.6151
R1168 B.n303 B.n302 10.6151
R1169 B.n303 B.n192 10.6151
R1170 B.n307 B.n192 10.6151
R1171 B.n308 B.n307 10.6151
R1172 B.n309 B.n308 10.6151
R1173 B.n309 B.n190 10.6151
R1174 B.n313 B.n190 10.6151
R1175 B.n314 B.n313 10.6151
R1176 B.n315 B.n314 10.6151
R1177 B.n315 B.n188 10.6151
R1178 B.n319 B.n188 10.6151
R1179 B.n320 B.n319 10.6151
R1180 B.n321 B.n320 10.6151
R1181 B.n321 B.n186 10.6151
R1182 B.n325 B.n186 10.6151
R1183 B.n326 B.n325 10.6151
R1184 B.n327 B.n326 10.6151
R1185 B.n327 B.n184 10.6151
R1186 B.n331 B.n184 10.6151
R1187 B.n332 B.n331 10.6151
R1188 B.n333 B.n332 10.6151
R1189 B.n333 B.n182 10.6151
R1190 B.n337 B.n182 10.6151
R1191 B.n338 B.n337 10.6151
R1192 B.n339 B.n338 10.6151
R1193 B.n339 B.n180 10.6151
R1194 B.n343 B.n180 10.6151
R1195 B.n344 B.n343 10.6151
R1196 B.n345 B.n344 10.6151
R1197 B.n345 B.n178 10.6151
R1198 B.n349 B.n178 10.6151
R1199 B.n350 B.n349 10.6151
R1200 B.n351 B.n350 10.6151
R1201 B.n351 B.n176 10.6151
R1202 B.n355 B.n176 10.6151
R1203 B.n356 B.n355 10.6151
R1204 B.n357 B.n356 10.6151
R1205 B.n357 B.n174 10.6151
R1206 B.n361 B.n174 10.6151
R1207 B.n362 B.n361 10.6151
R1208 B.n363 B.n362 10.6151
R1209 B.n363 B.n172 10.6151
R1210 B.n367 B.n172 10.6151
R1211 B.n368 B.n367 10.6151
R1212 B.n370 B.n168 10.6151
R1213 B.n374 B.n168 10.6151
R1214 B.n375 B.n374 10.6151
R1215 B.n376 B.n375 10.6151
R1216 B.n376 B.n166 10.6151
R1217 B.n380 B.n166 10.6151
R1218 B.n381 B.n380 10.6151
R1219 B.n382 B.n381 10.6151
R1220 B.n386 B.n385 10.6151
R1221 B.n387 B.n386 10.6151
R1222 B.n387 B.n160 10.6151
R1223 B.n391 B.n160 10.6151
R1224 B.n392 B.n391 10.6151
R1225 B.n393 B.n392 10.6151
R1226 B.n393 B.n158 10.6151
R1227 B.n397 B.n158 10.6151
R1228 B.n398 B.n397 10.6151
R1229 B.n399 B.n398 10.6151
R1230 B.n399 B.n156 10.6151
R1231 B.n403 B.n156 10.6151
R1232 B.n404 B.n403 10.6151
R1233 B.n405 B.n404 10.6151
R1234 B.n405 B.n154 10.6151
R1235 B.n409 B.n154 10.6151
R1236 B.n410 B.n409 10.6151
R1237 B.n411 B.n410 10.6151
R1238 B.n411 B.n152 10.6151
R1239 B.n415 B.n152 10.6151
R1240 B.n416 B.n415 10.6151
R1241 B.n417 B.n416 10.6151
R1242 B.n417 B.n150 10.6151
R1243 B.n421 B.n150 10.6151
R1244 B.n422 B.n421 10.6151
R1245 B.n423 B.n422 10.6151
R1246 B.n423 B.n148 10.6151
R1247 B.n427 B.n148 10.6151
R1248 B.n428 B.n427 10.6151
R1249 B.n429 B.n428 10.6151
R1250 B.n429 B.n146 10.6151
R1251 B.n433 B.n146 10.6151
R1252 B.n434 B.n433 10.6151
R1253 B.n435 B.n434 10.6151
R1254 B.n435 B.n144 10.6151
R1255 B.n439 B.n144 10.6151
R1256 B.n440 B.n439 10.6151
R1257 B.n441 B.n440 10.6151
R1258 B.n441 B.n142 10.6151
R1259 B.n445 B.n142 10.6151
R1260 B.n446 B.n445 10.6151
R1261 B.n447 B.n446 10.6151
R1262 B.n447 B.n140 10.6151
R1263 B.n451 B.n140 10.6151
R1264 B.n452 B.n451 10.6151
R1265 B.n453 B.n452 10.6151
R1266 B.n453 B.n138 10.6151
R1267 B.n457 B.n138 10.6151
R1268 B.n458 B.n457 10.6151
R1269 B.n459 B.n458 10.6151
R1270 B.n459 B.n136 10.6151
R1271 B.n463 B.n136 10.6151
R1272 B.n464 B.n463 10.6151
R1273 B.n465 B.n464 10.6151
R1274 B.n465 B.n134 10.6151
R1275 B.n469 B.n134 10.6151
R1276 B.n470 B.n469 10.6151
R1277 B.n471 B.n470 10.6151
R1278 B.n853 B.n0 8.11757
R1279 B.n853 B.n1 8.11757
R1280 B.n700 B.n54 6.5566
R1281 B.n688 B.n687 6.5566
R1282 B.n370 B.n369 6.5566
R1283 B.n382 B.n164 6.5566
R1284 B.n703 B.n54 4.05904
R1285 B.n687 B.n686 4.05904
R1286 B.n369 B.n368 4.05904
R1287 B.n385 B.n164 4.05904
R1288 VN.n4 VN.t5 203.425
R1289 VN.n20 VN.t2 203.425
R1290 VN.n3 VN.t4 171.581
R1291 VN.n14 VN.t1 171.581
R1292 VN.n19 VN.t0 171.581
R1293 VN.n30 VN.t3 171.581
R1294 VN.n29 VN.n16 161.3
R1295 VN.n28 VN.n27 161.3
R1296 VN.n26 VN.n17 161.3
R1297 VN.n25 VN.n24 161.3
R1298 VN.n23 VN.n18 161.3
R1299 VN.n22 VN.n21 161.3
R1300 VN.n13 VN.n0 161.3
R1301 VN.n12 VN.n11 161.3
R1302 VN.n10 VN.n1 161.3
R1303 VN.n9 VN.n8 161.3
R1304 VN.n7 VN.n2 161.3
R1305 VN.n6 VN.n5 161.3
R1306 VN.n15 VN.n14 106.353
R1307 VN.n31 VN.n30 106.353
R1308 VN.n4 VN.n3 59.8676
R1309 VN.n20 VN.n19 59.8676
R1310 VN.n8 VN.n1 56.5193
R1311 VN.n24 VN.n17 56.5193
R1312 VN VN.n31 52.9603
R1313 VN.n7 VN.n6 24.4675
R1314 VN.n8 VN.n7 24.4675
R1315 VN.n12 VN.n1 24.4675
R1316 VN.n13 VN.n12 24.4675
R1317 VN.n24 VN.n23 24.4675
R1318 VN.n23 VN.n22 24.4675
R1319 VN.n29 VN.n28 24.4675
R1320 VN.n28 VN.n17 24.4675
R1321 VN.n6 VN.n3 12.234
R1322 VN.n22 VN.n19 12.234
R1323 VN.n21 VN.n20 7.20192
R1324 VN.n5 VN.n4 7.20192
R1325 VN.n14 VN.n13 4.40456
R1326 VN.n30 VN.n29 4.40456
R1327 VN.n31 VN.n16 0.278367
R1328 VN.n15 VN.n0 0.278367
R1329 VN.n27 VN.n16 0.189894
R1330 VN.n27 VN.n26 0.189894
R1331 VN.n26 VN.n25 0.189894
R1332 VN.n25 VN.n18 0.189894
R1333 VN.n21 VN.n18 0.189894
R1334 VN.n5 VN.n2 0.189894
R1335 VN.n9 VN.n2 0.189894
R1336 VN.n10 VN.n9 0.189894
R1337 VN.n11 VN.n10 0.189894
R1338 VN.n11 VN.n0 0.189894
R1339 VN VN.n15 0.153454
R1340 VDD2.n1 VDD2.t1 72.2563
R1341 VDD2.n2 VDD2.t5 70.4757
R1342 VDD2.n1 VDD2.n0 69.2132
R1343 VDD2 VDD2.n3 69.2104
R1344 VDD2.n2 VDD2.n1 47.0774
R1345 VDD2 VDD2.n2 1.8949
R1346 VDD2.n3 VDD2.t4 1.81947
R1347 VDD2.n3 VDD2.t2 1.81947
R1348 VDD2.n0 VDD2.t0 1.81947
R1349 VDD2.n0 VDD2.t3 1.81947
R1350 VTAIL.n7 VTAIL.t9 53.7969
R1351 VTAIL.n11 VTAIL.t10 53.7967
R1352 VTAIL.n2 VTAIL.t1 53.7967
R1353 VTAIL.n10 VTAIL.t5 53.7967
R1354 VTAIL.n9 VTAIL.n8 51.978
R1355 VTAIL.n6 VTAIL.n5 51.978
R1356 VTAIL.n1 VTAIL.n0 51.9777
R1357 VTAIL.n4 VTAIL.n3 51.9777
R1358 VTAIL.n6 VTAIL.n4 32.6686
R1359 VTAIL.n11 VTAIL.n10 30.2203
R1360 VTAIL.n7 VTAIL.n6 2.44878
R1361 VTAIL.n10 VTAIL.n9 2.44878
R1362 VTAIL.n4 VTAIL.n2 2.44878
R1363 VTAIL.n0 VTAIL.t6 1.81947
R1364 VTAIL.n0 VTAIL.t7 1.81947
R1365 VTAIL.n3 VTAIL.t2 1.81947
R1366 VTAIL.n3 VTAIL.t4 1.81947
R1367 VTAIL.n8 VTAIL.t3 1.81947
R1368 VTAIL.n8 VTAIL.t0 1.81947
R1369 VTAIL.n5 VTAIL.t8 1.81947
R1370 VTAIL.n5 VTAIL.t11 1.81947
R1371 VTAIL VTAIL.n11 1.77852
R1372 VTAIL.n9 VTAIL.n7 1.69447
R1373 VTAIL.n2 VTAIL.n1 1.69447
R1374 VTAIL VTAIL.n1 0.670759
R1375 VP.n11 VP.t1 203.425
R1376 VP.n24 VP.t5 171.581
R1377 VP.n3 VP.t2 171.581
R1378 VP.n43 VP.t3 171.581
R1379 VP.n21 VP.t0 171.581
R1380 VP.n10 VP.t4 171.581
R1381 VP.n13 VP.n12 161.3
R1382 VP.n14 VP.n9 161.3
R1383 VP.n16 VP.n15 161.3
R1384 VP.n17 VP.n8 161.3
R1385 VP.n19 VP.n18 161.3
R1386 VP.n20 VP.n7 161.3
R1387 VP.n42 VP.n0 161.3
R1388 VP.n41 VP.n40 161.3
R1389 VP.n39 VP.n1 161.3
R1390 VP.n38 VP.n37 161.3
R1391 VP.n36 VP.n2 161.3
R1392 VP.n35 VP.n34 161.3
R1393 VP.n33 VP.n32 161.3
R1394 VP.n31 VP.n4 161.3
R1395 VP.n30 VP.n29 161.3
R1396 VP.n28 VP.n5 161.3
R1397 VP.n27 VP.n26 161.3
R1398 VP.n25 VP.n6 161.3
R1399 VP.n24 VP.n23 106.353
R1400 VP.n44 VP.n43 106.353
R1401 VP.n22 VP.n21 106.353
R1402 VP.n11 VP.n10 59.8676
R1403 VP.n30 VP.n5 56.5193
R1404 VP.n37 VP.n1 56.5193
R1405 VP.n15 VP.n8 56.5193
R1406 VP.n23 VP.n22 52.6814
R1407 VP.n26 VP.n25 24.4675
R1408 VP.n26 VP.n5 24.4675
R1409 VP.n31 VP.n30 24.4675
R1410 VP.n32 VP.n31 24.4675
R1411 VP.n36 VP.n35 24.4675
R1412 VP.n37 VP.n36 24.4675
R1413 VP.n41 VP.n1 24.4675
R1414 VP.n42 VP.n41 24.4675
R1415 VP.n19 VP.n8 24.4675
R1416 VP.n20 VP.n19 24.4675
R1417 VP.n14 VP.n13 24.4675
R1418 VP.n15 VP.n14 24.4675
R1419 VP.n32 VP.n3 12.234
R1420 VP.n35 VP.n3 12.234
R1421 VP.n13 VP.n10 12.234
R1422 VP.n12 VP.n11 7.20192
R1423 VP.n25 VP.n24 4.40456
R1424 VP.n43 VP.n42 4.40456
R1425 VP.n21 VP.n20 4.40456
R1426 VP.n22 VP.n7 0.278367
R1427 VP.n23 VP.n6 0.278367
R1428 VP.n44 VP.n0 0.278367
R1429 VP.n12 VP.n9 0.189894
R1430 VP.n16 VP.n9 0.189894
R1431 VP.n17 VP.n16 0.189894
R1432 VP.n18 VP.n17 0.189894
R1433 VP.n18 VP.n7 0.189894
R1434 VP.n27 VP.n6 0.189894
R1435 VP.n28 VP.n27 0.189894
R1436 VP.n29 VP.n28 0.189894
R1437 VP.n29 VP.n4 0.189894
R1438 VP.n33 VP.n4 0.189894
R1439 VP.n34 VP.n33 0.189894
R1440 VP.n34 VP.n2 0.189894
R1441 VP.n38 VP.n2 0.189894
R1442 VP.n39 VP.n38 0.189894
R1443 VP.n40 VP.n39 0.189894
R1444 VP.n40 VP.n0 0.189894
R1445 VP VP.n44 0.153454
R1446 VDD1 VDD1.t4 72.3701
R1447 VDD1.n1 VDD1.t0 72.2563
R1448 VDD1.n1 VDD1.n0 69.2132
R1449 VDD1.n3 VDD1.n2 68.6566
R1450 VDD1.n3 VDD1.n1 48.8845
R1451 VDD1.n2 VDD1.t1 1.81947
R1452 VDD1.n2 VDD1.t5 1.81947
R1453 VDD1.n0 VDD1.t3 1.81947
R1454 VDD1.n0 VDD1.t2 1.81947
R1455 VDD1 VDD1.n3 0.554379
C0 VTAIL B 4.96403f
C1 VDD1 VDD2 1.3732f
C2 VTAIL w_n3242_n4542# 3.7918f
C3 VN VP 7.93028f
C4 VTAIL VDD2 9.922421f
C5 w_n3242_n4542# B 11.1975f
C6 VN VDD1 0.150696f
C7 VDD2 B 2.60361f
C8 VTAIL VN 9.632759f
C9 VDD2 w_n3242_n4542# 2.76164f
C10 VN B 1.21707f
C11 VN w_n3242_n4542# 6.23688f
C12 VDD1 VP 10.053599f
C13 VN VDD2 9.75731f
C14 VTAIL VP 9.64715f
C15 VP B 1.916f
C16 VTAIL VDD1 9.8737f
C17 VP w_n3242_n4542# 6.65577f
C18 VDD2 VP 0.451255f
C19 VDD1 B 2.53168f
C20 VDD1 w_n3242_n4542# 2.67946f
C21 VDD2 VSUBS 2.06198f
C22 VDD1 VSUBS 2.54445f
C23 VTAIL VSUBS 1.38368f
C24 VN VSUBS 5.99306f
C25 VP VSUBS 3.074906f
C26 B VSUBS 5.046135f
C27 w_n3242_n4542# VSUBS 0.180087p
C28 VDD1.t4 VSUBS 4.13279f
C29 VDD1.t0 VSUBS 4.13131f
C30 VDD1.t3 VSUBS 0.381979f
C31 VDD1.t2 VSUBS 0.381979f
C32 VDD1.n0 VSUBS 3.17515f
C33 VDD1.n1 VSUBS 4.27796f
C34 VDD1.t1 VSUBS 0.381979f
C35 VDD1.t5 VSUBS 0.381979f
C36 VDD1.n2 VSUBS 3.16864f
C37 VDD1.n3 VSUBS 3.78445f
C38 VP.n0 VSUBS 0.037776f
C39 VP.t3 VSUBS 3.53448f
C40 VP.n1 VSUBS 0.048215f
C41 VP.n2 VSUBS 0.028653f
C42 VP.t2 VSUBS 3.53448f
C43 VP.n3 VSUBS 1.22692f
C44 VP.n4 VSUBS 0.028653f
C45 VP.n5 VSUBS 0.048215f
C46 VP.n6 VSUBS 0.037776f
C47 VP.t5 VSUBS 3.53448f
C48 VP.n7 VSUBS 0.037776f
C49 VP.t0 VSUBS 3.53448f
C50 VP.n8 VSUBS 0.048215f
C51 VP.n9 VSUBS 0.028653f
C52 VP.t4 VSUBS 3.53448f
C53 VP.n10 VSUBS 1.30776f
C54 VP.t1 VSUBS 3.75327f
C55 VP.n11 VSUBS 1.28936f
C56 VP.n12 VSUBS 0.273696f
C57 VP.n13 VSUBS 0.040219f
C58 VP.n14 VSUBS 0.053401f
C59 VP.n15 VSUBS 0.03544f
C60 VP.n16 VSUBS 0.028653f
C61 VP.n17 VSUBS 0.028653f
C62 VP.n18 VSUBS 0.028653f
C63 VP.n19 VSUBS 0.053401f
C64 VP.n20 VSUBS 0.031782f
C65 VP.n21 VSUBS 1.31107f
C66 VP.n22 VSUBS 1.72128f
C67 VP.n23 VSUBS 1.74083f
C68 VP.n24 VSUBS 1.31107f
C69 VP.n25 VSUBS 0.031782f
C70 VP.n26 VSUBS 0.053401f
C71 VP.n27 VSUBS 0.028653f
C72 VP.n28 VSUBS 0.028653f
C73 VP.n29 VSUBS 0.028653f
C74 VP.n30 VSUBS 0.03544f
C75 VP.n31 VSUBS 0.053401f
C76 VP.n32 VSUBS 0.040219f
C77 VP.n33 VSUBS 0.028653f
C78 VP.n34 VSUBS 0.028653f
C79 VP.n35 VSUBS 0.040219f
C80 VP.n36 VSUBS 0.053401f
C81 VP.n37 VSUBS 0.03544f
C82 VP.n38 VSUBS 0.028653f
C83 VP.n39 VSUBS 0.028653f
C84 VP.n40 VSUBS 0.028653f
C85 VP.n41 VSUBS 0.053401f
C86 VP.n42 VSUBS 0.031782f
C87 VP.n43 VSUBS 1.31107f
C88 VP.n44 VSUBS 0.049313f
C89 VTAIL.t6 VSUBS 0.38869f
C90 VTAIL.t7 VSUBS 0.38869f
C91 VTAIL.n0 VSUBS 3.05138f
C92 VTAIL.n1 VSUBS 0.889375f
C93 VTAIL.t1 VSUBS 3.98557f
C94 VTAIL.n2 VSUBS 1.17294f
C95 VTAIL.t2 VSUBS 0.38869f
C96 VTAIL.t4 VSUBS 0.38869f
C97 VTAIL.n3 VSUBS 3.05138f
C98 VTAIL.n4 VSUBS 3.07131f
C99 VTAIL.t8 VSUBS 0.38869f
C100 VTAIL.t11 VSUBS 0.38869f
C101 VTAIL.n5 VSUBS 3.05138f
C102 VTAIL.n6 VSUBS 3.0713f
C103 VTAIL.t9 VSUBS 3.98557f
C104 VTAIL.n7 VSUBS 1.17294f
C105 VTAIL.t3 VSUBS 0.38869f
C106 VTAIL.t0 VSUBS 0.38869f
C107 VTAIL.n8 VSUBS 3.05138f
C108 VTAIL.n9 VSUBS 1.04706f
C109 VTAIL.t5 VSUBS 3.98557f
C110 VTAIL.n10 VSUBS 2.98004f
C111 VTAIL.t10 VSUBS 3.98557f
C112 VTAIL.n11 VSUBS 2.92059f
C113 VDD2.t1 VSUBS 4.1313f
C114 VDD2.t0 VSUBS 0.381977f
C115 VDD2.t3 VSUBS 0.381977f
C116 VDD2.n0 VSUBS 3.17514f
C117 VDD2.n1 VSUBS 4.14205f
C118 VDD2.t5 VSUBS 4.11158f
C119 VDD2.n2 VSUBS 3.82266f
C120 VDD2.t4 VSUBS 0.381977f
C121 VDD2.t2 VSUBS 0.381977f
C122 VDD2.n3 VSUBS 3.17508f
C123 VN.n0 VSUBS 0.036851f
C124 VN.t1 VSUBS 3.44799f
C125 VN.n1 VSUBS 0.047035f
C126 VN.n2 VSUBS 0.027951f
C127 VN.t4 VSUBS 3.44799f
C128 VN.n3 VSUBS 1.27576f
C129 VN.t5 VSUBS 3.66143f
C130 VN.n4 VSUBS 1.25781f
C131 VN.n5 VSUBS 0.266999f
C132 VN.n6 VSUBS 0.039235f
C133 VN.n7 VSUBS 0.052095f
C134 VN.n8 VSUBS 0.034573f
C135 VN.n9 VSUBS 0.027951f
C136 VN.n10 VSUBS 0.027951f
C137 VN.n11 VSUBS 0.027951f
C138 VN.n12 VSUBS 0.052095f
C139 VN.n13 VSUBS 0.031005f
C140 VN.n14 VSUBS 1.27899f
C141 VN.n15 VSUBS 0.048106f
C142 VN.n16 VSUBS 0.036851f
C143 VN.t3 VSUBS 3.44799f
C144 VN.n17 VSUBS 0.047035f
C145 VN.n18 VSUBS 0.027951f
C146 VN.t0 VSUBS 3.44799f
C147 VN.n19 VSUBS 1.27576f
C148 VN.t2 VSUBS 3.66143f
C149 VN.n20 VSUBS 1.25781f
C150 VN.n21 VSUBS 0.266999f
C151 VN.n22 VSUBS 0.039235f
C152 VN.n23 VSUBS 0.052095f
C153 VN.n24 VSUBS 0.034573f
C154 VN.n25 VSUBS 0.027951f
C155 VN.n26 VSUBS 0.027951f
C156 VN.n27 VSUBS 0.027951f
C157 VN.n28 VSUBS 0.052095f
C158 VN.n29 VSUBS 0.031005f
C159 VN.n30 VSUBS 1.27899f
C160 VN.n31 VSUBS 1.69406f
C161 B.n0 VSUBS 0.006382f
C162 B.n1 VSUBS 0.006382f
C163 B.n2 VSUBS 0.009438f
C164 B.n3 VSUBS 0.007233f
C165 B.n4 VSUBS 0.007233f
C166 B.n5 VSUBS 0.007233f
C167 B.n6 VSUBS 0.007233f
C168 B.n7 VSUBS 0.007233f
C169 B.n8 VSUBS 0.007233f
C170 B.n9 VSUBS 0.007233f
C171 B.n10 VSUBS 0.007233f
C172 B.n11 VSUBS 0.007233f
C173 B.n12 VSUBS 0.007233f
C174 B.n13 VSUBS 0.007233f
C175 B.n14 VSUBS 0.007233f
C176 B.n15 VSUBS 0.007233f
C177 B.n16 VSUBS 0.007233f
C178 B.n17 VSUBS 0.007233f
C179 B.n18 VSUBS 0.007233f
C180 B.n19 VSUBS 0.007233f
C181 B.n20 VSUBS 0.007233f
C182 B.n21 VSUBS 0.007233f
C183 B.n22 VSUBS 0.017264f
C184 B.n23 VSUBS 0.007233f
C185 B.n24 VSUBS 0.007233f
C186 B.n25 VSUBS 0.007233f
C187 B.n26 VSUBS 0.007233f
C188 B.n27 VSUBS 0.007233f
C189 B.n28 VSUBS 0.007233f
C190 B.n29 VSUBS 0.007233f
C191 B.n30 VSUBS 0.007233f
C192 B.n31 VSUBS 0.007233f
C193 B.n32 VSUBS 0.007233f
C194 B.n33 VSUBS 0.007233f
C195 B.n34 VSUBS 0.007233f
C196 B.n35 VSUBS 0.007233f
C197 B.n36 VSUBS 0.007233f
C198 B.n37 VSUBS 0.007233f
C199 B.n38 VSUBS 0.007233f
C200 B.n39 VSUBS 0.007233f
C201 B.n40 VSUBS 0.007233f
C202 B.n41 VSUBS 0.007233f
C203 B.n42 VSUBS 0.007233f
C204 B.n43 VSUBS 0.007233f
C205 B.n44 VSUBS 0.007233f
C206 B.n45 VSUBS 0.007233f
C207 B.n46 VSUBS 0.007233f
C208 B.n47 VSUBS 0.007233f
C209 B.n48 VSUBS 0.007233f
C210 B.n49 VSUBS 0.007233f
C211 B.n50 VSUBS 0.007233f
C212 B.n51 VSUBS 0.007233f
C213 B.t7 VSUBS 0.623048f
C214 B.t8 VSUBS 0.644349f
C215 B.t6 VSUBS 2.05141f
C216 B.n52 VSUBS 0.348303f
C217 B.n53 VSUBS 0.07411f
C218 B.n54 VSUBS 0.016758f
C219 B.n55 VSUBS 0.007233f
C220 B.n56 VSUBS 0.007233f
C221 B.n57 VSUBS 0.007233f
C222 B.n58 VSUBS 0.007233f
C223 B.n59 VSUBS 0.007233f
C224 B.t4 VSUBS 0.623026f
C225 B.t5 VSUBS 0.644331f
C226 B.t3 VSUBS 2.05141f
C227 B.n60 VSUBS 0.348321f
C228 B.n61 VSUBS 0.074132f
C229 B.n62 VSUBS 0.007233f
C230 B.n63 VSUBS 0.007233f
C231 B.n64 VSUBS 0.007233f
C232 B.n65 VSUBS 0.007233f
C233 B.n66 VSUBS 0.007233f
C234 B.n67 VSUBS 0.007233f
C235 B.n68 VSUBS 0.007233f
C236 B.n69 VSUBS 0.007233f
C237 B.n70 VSUBS 0.007233f
C238 B.n71 VSUBS 0.007233f
C239 B.n72 VSUBS 0.007233f
C240 B.n73 VSUBS 0.007233f
C241 B.n74 VSUBS 0.007233f
C242 B.n75 VSUBS 0.007233f
C243 B.n76 VSUBS 0.007233f
C244 B.n77 VSUBS 0.007233f
C245 B.n78 VSUBS 0.007233f
C246 B.n79 VSUBS 0.007233f
C247 B.n80 VSUBS 0.007233f
C248 B.n81 VSUBS 0.007233f
C249 B.n82 VSUBS 0.007233f
C250 B.n83 VSUBS 0.007233f
C251 B.n84 VSUBS 0.007233f
C252 B.n85 VSUBS 0.007233f
C253 B.n86 VSUBS 0.007233f
C254 B.n87 VSUBS 0.007233f
C255 B.n88 VSUBS 0.007233f
C256 B.n89 VSUBS 0.007233f
C257 B.n90 VSUBS 0.017836f
C258 B.n91 VSUBS 0.007233f
C259 B.n92 VSUBS 0.007233f
C260 B.n93 VSUBS 0.007233f
C261 B.n94 VSUBS 0.007233f
C262 B.n95 VSUBS 0.007233f
C263 B.n96 VSUBS 0.007233f
C264 B.n97 VSUBS 0.007233f
C265 B.n98 VSUBS 0.007233f
C266 B.n99 VSUBS 0.007233f
C267 B.n100 VSUBS 0.007233f
C268 B.n101 VSUBS 0.007233f
C269 B.n102 VSUBS 0.007233f
C270 B.n103 VSUBS 0.007233f
C271 B.n104 VSUBS 0.007233f
C272 B.n105 VSUBS 0.007233f
C273 B.n106 VSUBS 0.007233f
C274 B.n107 VSUBS 0.007233f
C275 B.n108 VSUBS 0.007233f
C276 B.n109 VSUBS 0.007233f
C277 B.n110 VSUBS 0.007233f
C278 B.n111 VSUBS 0.007233f
C279 B.n112 VSUBS 0.007233f
C280 B.n113 VSUBS 0.007233f
C281 B.n114 VSUBS 0.007233f
C282 B.n115 VSUBS 0.007233f
C283 B.n116 VSUBS 0.007233f
C284 B.n117 VSUBS 0.007233f
C285 B.n118 VSUBS 0.007233f
C286 B.n119 VSUBS 0.007233f
C287 B.n120 VSUBS 0.007233f
C288 B.n121 VSUBS 0.007233f
C289 B.n122 VSUBS 0.007233f
C290 B.n123 VSUBS 0.007233f
C291 B.n124 VSUBS 0.007233f
C292 B.n125 VSUBS 0.007233f
C293 B.n126 VSUBS 0.007233f
C294 B.n127 VSUBS 0.007233f
C295 B.n128 VSUBS 0.007233f
C296 B.n129 VSUBS 0.007233f
C297 B.n130 VSUBS 0.007233f
C298 B.n131 VSUBS 0.007233f
C299 B.n132 VSUBS 0.018073f
C300 B.n133 VSUBS 0.007233f
C301 B.n134 VSUBS 0.007233f
C302 B.n135 VSUBS 0.007233f
C303 B.n136 VSUBS 0.007233f
C304 B.n137 VSUBS 0.007233f
C305 B.n138 VSUBS 0.007233f
C306 B.n139 VSUBS 0.007233f
C307 B.n140 VSUBS 0.007233f
C308 B.n141 VSUBS 0.007233f
C309 B.n142 VSUBS 0.007233f
C310 B.n143 VSUBS 0.007233f
C311 B.n144 VSUBS 0.007233f
C312 B.n145 VSUBS 0.007233f
C313 B.n146 VSUBS 0.007233f
C314 B.n147 VSUBS 0.007233f
C315 B.n148 VSUBS 0.007233f
C316 B.n149 VSUBS 0.007233f
C317 B.n150 VSUBS 0.007233f
C318 B.n151 VSUBS 0.007233f
C319 B.n152 VSUBS 0.007233f
C320 B.n153 VSUBS 0.007233f
C321 B.n154 VSUBS 0.007233f
C322 B.n155 VSUBS 0.007233f
C323 B.n156 VSUBS 0.007233f
C324 B.n157 VSUBS 0.007233f
C325 B.n158 VSUBS 0.007233f
C326 B.n159 VSUBS 0.007233f
C327 B.n160 VSUBS 0.007233f
C328 B.n161 VSUBS 0.007233f
C329 B.t2 VSUBS 0.623026f
C330 B.t1 VSUBS 0.644331f
C331 B.t0 VSUBS 2.05141f
C332 B.n162 VSUBS 0.348321f
C333 B.n163 VSUBS 0.074132f
C334 B.n164 VSUBS 0.016758f
C335 B.n165 VSUBS 0.007233f
C336 B.n166 VSUBS 0.007233f
C337 B.n167 VSUBS 0.007233f
C338 B.n168 VSUBS 0.007233f
C339 B.n169 VSUBS 0.007233f
C340 B.t11 VSUBS 0.623048f
C341 B.t10 VSUBS 0.644349f
C342 B.t9 VSUBS 2.05141f
C343 B.n170 VSUBS 0.348303f
C344 B.n171 VSUBS 0.07411f
C345 B.n172 VSUBS 0.007233f
C346 B.n173 VSUBS 0.007233f
C347 B.n174 VSUBS 0.007233f
C348 B.n175 VSUBS 0.007233f
C349 B.n176 VSUBS 0.007233f
C350 B.n177 VSUBS 0.007233f
C351 B.n178 VSUBS 0.007233f
C352 B.n179 VSUBS 0.007233f
C353 B.n180 VSUBS 0.007233f
C354 B.n181 VSUBS 0.007233f
C355 B.n182 VSUBS 0.007233f
C356 B.n183 VSUBS 0.007233f
C357 B.n184 VSUBS 0.007233f
C358 B.n185 VSUBS 0.007233f
C359 B.n186 VSUBS 0.007233f
C360 B.n187 VSUBS 0.007233f
C361 B.n188 VSUBS 0.007233f
C362 B.n189 VSUBS 0.007233f
C363 B.n190 VSUBS 0.007233f
C364 B.n191 VSUBS 0.007233f
C365 B.n192 VSUBS 0.007233f
C366 B.n193 VSUBS 0.007233f
C367 B.n194 VSUBS 0.007233f
C368 B.n195 VSUBS 0.007233f
C369 B.n196 VSUBS 0.007233f
C370 B.n197 VSUBS 0.007233f
C371 B.n198 VSUBS 0.007233f
C372 B.n199 VSUBS 0.007233f
C373 B.n200 VSUBS 0.017836f
C374 B.n201 VSUBS 0.007233f
C375 B.n202 VSUBS 0.007233f
C376 B.n203 VSUBS 0.007233f
C377 B.n204 VSUBS 0.007233f
C378 B.n205 VSUBS 0.007233f
C379 B.n206 VSUBS 0.007233f
C380 B.n207 VSUBS 0.007233f
C381 B.n208 VSUBS 0.007233f
C382 B.n209 VSUBS 0.007233f
C383 B.n210 VSUBS 0.007233f
C384 B.n211 VSUBS 0.007233f
C385 B.n212 VSUBS 0.007233f
C386 B.n213 VSUBS 0.007233f
C387 B.n214 VSUBS 0.007233f
C388 B.n215 VSUBS 0.007233f
C389 B.n216 VSUBS 0.007233f
C390 B.n217 VSUBS 0.007233f
C391 B.n218 VSUBS 0.007233f
C392 B.n219 VSUBS 0.007233f
C393 B.n220 VSUBS 0.007233f
C394 B.n221 VSUBS 0.007233f
C395 B.n222 VSUBS 0.007233f
C396 B.n223 VSUBS 0.007233f
C397 B.n224 VSUBS 0.007233f
C398 B.n225 VSUBS 0.007233f
C399 B.n226 VSUBS 0.007233f
C400 B.n227 VSUBS 0.007233f
C401 B.n228 VSUBS 0.007233f
C402 B.n229 VSUBS 0.007233f
C403 B.n230 VSUBS 0.007233f
C404 B.n231 VSUBS 0.007233f
C405 B.n232 VSUBS 0.007233f
C406 B.n233 VSUBS 0.007233f
C407 B.n234 VSUBS 0.007233f
C408 B.n235 VSUBS 0.007233f
C409 B.n236 VSUBS 0.007233f
C410 B.n237 VSUBS 0.007233f
C411 B.n238 VSUBS 0.007233f
C412 B.n239 VSUBS 0.007233f
C413 B.n240 VSUBS 0.007233f
C414 B.n241 VSUBS 0.007233f
C415 B.n242 VSUBS 0.007233f
C416 B.n243 VSUBS 0.007233f
C417 B.n244 VSUBS 0.007233f
C418 B.n245 VSUBS 0.007233f
C419 B.n246 VSUBS 0.007233f
C420 B.n247 VSUBS 0.007233f
C421 B.n248 VSUBS 0.007233f
C422 B.n249 VSUBS 0.007233f
C423 B.n250 VSUBS 0.007233f
C424 B.n251 VSUBS 0.007233f
C425 B.n252 VSUBS 0.007233f
C426 B.n253 VSUBS 0.007233f
C427 B.n254 VSUBS 0.007233f
C428 B.n255 VSUBS 0.007233f
C429 B.n256 VSUBS 0.007233f
C430 B.n257 VSUBS 0.007233f
C431 B.n258 VSUBS 0.007233f
C432 B.n259 VSUBS 0.007233f
C433 B.n260 VSUBS 0.007233f
C434 B.n261 VSUBS 0.007233f
C435 B.n262 VSUBS 0.007233f
C436 B.n263 VSUBS 0.007233f
C437 B.n264 VSUBS 0.007233f
C438 B.n265 VSUBS 0.007233f
C439 B.n266 VSUBS 0.007233f
C440 B.n267 VSUBS 0.007233f
C441 B.n268 VSUBS 0.007233f
C442 B.n269 VSUBS 0.007233f
C443 B.n270 VSUBS 0.007233f
C444 B.n271 VSUBS 0.007233f
C445 B.n272 VSUBS 0.007233f
C446 B.n273 VSUBS 0.007233f
C447 B.n274 VSUBS 0.007233f
C448 B.n275 VSUBS 0.007233f
C449 B.n276 VSUBS 0.007233f
C450 B.n277 VSUBS 0.007233f
C451 B.n278 VSUBS 0.007233f
C452 B.n279 VSUBS 0.017264f
C453 B.n280 VSUBS 0.017264f
C454 B.n281 VSUBS 0.017836f
C455 B.n282 VSUBS 0.007233f
C456 B.n283 VSUBS 0.007233f
C457 B.n284 VSUBS 0.007233f
C458 B.n285 VSUBS 0.007233f
C459 B.n286 VSUBS 0.007233f
C460 B.n287 VSUBS 0.007233f
C461 B.n288 VSUBS 0.007233f
C462 B.n289 VSUBS 0.007233f
C463 B.n290 VSUBS 0.007233f
C464 B.n291 VSUBS 0.007233f
C465 B.n292 VSUBS 0.007233f
C466 B.n293 VSUBS 0.007233f
C467 B.n294 VSUBS 0.007233f
C468 B.n295 VSUBS 0.007233f
C469 B.n296 VSUBS 0.007233f
C470 B.n297 VSUBS 0.007233f
C471 B.n298 VSUBS 0.007233f
C472 B.n299 VSUBS 0.007233f
C473 B.n300 VSUBS 0.007233f
C474 B.n301 VSUBS 0.007233f
C475 B.n302 VSUBS 0.007233f
C476 B.n303 VSUBS 0.007233f
C477 B.n304 VSUBS 0.007233f
C478 B.n305 VSUBS 0.007233f
C479 B.n306 VSUBS 0.007233f
C480 B.n307 VSUBS 0.007233f
C481 B.n308 VSUBS 0.007233f
C482 B.n309 VSUBS 0.007233f
C483 B.n310 VSUBS 0.007233f
C484 B.n311 VSUBS 0.007233f
C485 B.n312 VSUBS 0.007233f
C486 B.n313 VSUBS 0.007233f
C487 B.n314 VSUBS 0.007233f
C488 B.n315 VSUBS 0.007233f
C489 B.n316 VSUBS 0.007233f
C490 B.n317 VSUBS 0.007233f
C491 B.n318 VSUBS 0.007233f
C492 B.n319 VSUBS 0.007233f
C493 B.n320 VSUBS 0.007233f
C494 B.n321 VSUBS 0.007233f
C495 B.n322 VSUBS 0.007233f
C496 B.n323 VSUBS 0.007233f
C497 B.n324 VSUBS 0.007233f
C498 B.n325 VSUBS 0.007233f
C499 B.n326 VSUBS 0.007233f
C500 B.n327 VSUBS 0.007233f
C501 B.n328 VSUBS 0.007233f
C502 B.n329 VSUBS 0.007233f
C503 B.n330 VSUBS 0.007233f
C504 B.n331 VSUBS 0.007233f
C505 B.n332 VSUBS 0.007233f
C506 B.n333 VSUBS 0.007233f
C507 B.n334 VSUBS 0.007233f
C508 B.n335 VSUBS 0.007233f
C509 B.n336 VSUBS 0.007233f
C510 B.n337 VSUBS 0.007233f
C511 B.n338 VSUBS 0.007233f
C512 B.n339 VSUBS 0.007233f
C513 B.n340 VSUBS 0.007233f
C514 B.n341 VSUBS 0.007233f
C515 B.n342 VSUBS 0.007233f
C516 B.n343 VSUBS 0.007233f
C517 B.n344 VSUBS 0.007233f
C518 B.n345 VSUBS 0.007233f
C519 B.n346 VSUBS 0.007233f
C520 B.n347 VSUBS 0.007233f
C521 B.n348 VSUBS 0.007233f
C522 B.n349 VSUBS 0.007233f
C523 B.n350 VSUBS 0.007233f
C524 B.n351 VSUBS 0.007233f
C525 B.n352 VSUBS 0.007233f
C526 B.n353 VSUBS 0.007233f
C527 B.n354 VSUBS 0.007233f
C528 B.n355 VSUBS 0.007233f
C529 B.n356 VSUBS 0.007233f
C530 B.n357 VSUBS 0.007233f
C531 B.n358 VSUBS 0.007233f
C532 B.n359 VSUBS 0.007233f
C533 B.n360 VSUBS 0.007233f
C534 B.n361 VSUBS 0.007233f
C535 B.n362 VSUBS 0.007233f
C536 B.n363 VSUBS 0.007233f
C537 B.n364 VSUBS 0.007233f
C538 B.n365 VSUBS 0.007233f
C539 B.n366 VSUBS 0.007233f
C540 B.n367 VSUBS 0.007233f
C541 B.n368 VSUBS 0.004999f
C542 B.n369 VSUBS 0.016758f
C543 B.n370 VSUBS 0.00585f
C544 B.n371 VSUBS 0.007233f
C545 B.n372 VSUBS 0.007233f
C546 B.n373 VSUBS 0.007233f
C547 B.n374 VSUBS 0.007233f
C548 B.n375 VSUBS 0.007233f
C549 B.n376 VSUBS 0.007233f
C550 B.n377 VSUBS 0.007233f
C551 B.n378 VSUBS 0.007233f
C552 B.n379 VSUBS 0.007233f
C553 B.n380 VSUBS 0.007233f
C554 B.n381 VSUBS 0.007233f
C555 B.n382 VSUBS 0.00585f
C556 B.n383 VSUBS 0.007233f
C557 B.n384 VSUBS 0.007233f
C558 B.n385 VSUBS 0.004999f
C559 B.n386 VSUBS 0.007233f
C560 B.n387 VSUBS 0.007233f
C561 B.n388 VSUBS 0.007233f
C562 B.n389 VSUBS 0.007233f
C563 B.n390 VSUBS 0.007233f
C564 B.n391 VSUBS 0.007233f
C565 B.n392 VSUBS 0.007233f
C566 B.n393 VSUBS 0.007233f
C567 B.n394 VSUBS 0.007233f
C568 B.n395 VSUBS 0.007233f
C569 B.n396 VSUBS 0.007233f
C570 B.n397 VSUBS 0.007233f
C571 B.n398 VSUBS 0.007233f
C572 B.n399 VSUBS 0.007233f
C573 B.n400 VSUBS 0.007233f
C574 B.n401 VSUBS 0.007233f
C575 B.n402 VSUBS 0.007233f
C576 B.n403 VSUBS 0.007233f
C577 B.n404 VSUBS 0.007233f
C578 B.n405 VSUBS 0.007233f
C579 B.n406 VSUBS 0.007233f
C580 B.n407 VSUBS 0.007233f
C581 B.n408 VSUBS 0.007233f
C582 B.n409 VSUBS 0.007233f
C583 B.n410 VSUBS 0.007233f
C584 B.n411 VSUBS 0.007233f
C585 B.n412 VSUBS 0.007233f
C586 B.n413 VSUBS 0.007233f
C587 B.n414 VSUBS 0.007233f
C588 B.n415 VSUBS 0.007233f
C589 B.n416 VSUBS 0.007233f
C590 B.n417 VSUBS 0.007233f
C591 B.n418 VSUBS 0.007233f
C592 B.n419 VSUBS 0.007233f
C593 B.n420 VSUBS 0.007233f
C594 B.n421 VSUBS 0.007233f
C595 B.n422 VSUBS 0.007233f
C596 B.n423 VSUBS 0.007233f
C597 B.n424 VSUBS 0.007233f
C598 B.n425 VSUBS 0.007233f
C599 B.n426 VSUBS 0.007233f
C600 B.n427 VSUBS 0.007233f
C601 B.n428 VSUBS 0.007233f
C602 B.n429 VSUBS 0.007233f
C603 B.n430 VSUBS 0.007233f
C604 B.n431 VSUBS 0.007233f
C605 B.n432 VSUBS 0.007233f
C606 B.n433 VSUBS 0.007233f
C607 B.n434 VSUBS 0.007233f
C608 B.n435 VSUBS 0.007233f
C609 B.n436 VSUBS 0.007233f
C610 B.n437 VSUBS 0.007233f
C611 B.n438 VSUBS 0.007233f
C612 B.n439 VSUBS 0.007233f
C613 B.n440 VSUBS 0.007233f
C614 B.n441 VSUBS 0.007233f
C615 B.n442 VSUBS 0.007233f
C616 B.n443 VSUBS 0.007233f
C617 B.n444 VSUBS 0.007233f
C618 B.n445 VSUBS 0.007233f
C619 B.n446 VSUBS 0.007233f
C620 B.n447 VSUBS 0.007233f
C621 B.n448 VSUBS 0.007233f
C622 B.n449 VSUBS 0.007233f
C623 B.n450 VSUBS 0.007233f
C624 B.n451 VSUBS 0.007233f
C625 B.n452 VSUBS 0.007233f
C626 B.n453 VSUBS 0.007233f
C627 B.n454 VSUBS 0.007233f
C628 B.n455 VSUBS 0.007233f
C629 B.n456 VSUBS 0.007233f
C630 B.n457 VSUBS 0.007233f
C631 B.n458 VSUBS 0.007233f
C632 B.n459 VSUBS 0.007233f
C633 B.n460 VSUBS 0.007233f
C634 B.n461 VSUBS 0.007233f
C635 B.n462 VSUBS 0.007233f
C636 B.n463 VSUBS 0.007233f
C637 B.n464 VSUBS 0.007233f
C638 B.n465 VSUBS 0.007233f
C639 B.n466 VSUBS 0.007233f
C640 B.n467 VSUBS 0.007233f
C641 B.n468 VSUBS 0.007233f
C642 B.n469 VSUBS 0.007233f
C643 B.n470 VSUBS 0.007233f
C644 B.n471 VSUBS 0.017027f
C645 B.n472 VSUBS 0.017836f
C646 B.n473 VSUBS 0.017264f
C647 B.n474 VSUBS 0.007233f
C648 B.n475 VSUBS 0.007233f
C649 B.n476 VSUBS 0.007233f
C650 B.n477 VSUBS 0.007233f
C651 B.n478 VSUBS 0.007233f
C652 B.n479 VSUBS 0.007233f
C653 B.n480 VSUBS 0.007233f
C654 B.n481 VSUBS 0.007233f
C655 B.n482 VSUBS 0.007233f
C656 B.n483 VSUBS 0.007233f
C657 B.n484 VSUBS 0.007233f
C658 B.n485 VSUBS 0.007233f
C659 B.n486 VSUBS 0.007233f
C660 B.n487 VSUBS 0.007233f
C661 B.n488 VSUBS 0.007233f
C662 B.n489 VSUBS 0.007233f
C663 B.n490 VSUBS 0.007233f
C664 B.n491 VSUBS 0.007233f
C665 B.n492 VSUBS 0.007233f
C666 B.n493 VSUBS 0.007233f
C667 B.n494 VSUBS 0.007233f
C668 B.n495 VSUBS 0.007233f
C669 B.n496 VSUBS 0.007233f
C670 B.n497 VSUBS 0.007233f
C671 B.n498 VSUBS 0.007233f
C672 B.n499 VSUBS 0.007233f
C673 B.n500 VSUBS 0.007233f
C674 B.n501 VSUBS 0.007233f
C675 B.n502 VSUBS 0.007233f
C676 B.n503 VSUBS 0.007233f
C677 B.n504 VSUBS 0.007233f
C678 B.n505 VSUBS 0.007233f
C679 B.n506 VSUBS 0.007233f
C680 B.n507 VSUBS 0.007233f
C681 B.n508 VSUBS 0.007233f
C682 B.n509 VSUBS 0.007233f
C683 B.n510 VSUBS 0.007233f
C684 B.n511 VSUBS 0.007233f
C685 B.n512 VSUBS 0.007233f
C686 B.n513 VSUBS 0.007233f
C687 B.n514 VSUBS 0.007233f
C688 B.n515 VSUBS 0.007233f
C689 B.n516 VSUBS 0.007233f
C690 B.n517 VSUBS 0.007233f
C691 B.n518 VSUBS 0.007233f
C692 B.n519 VSUBS 0.007233f
C693 B.n520 VSUBS 0.007233f
C694 B.n521 VSUBS 0.007233f
C695 B.n522 VSUBS 0.007233f
C696 B.n523 VSUBS 0.007233f
C697 B.n524 VSUBS 0.007233f
C698 B.n525 VSUBS 0.007233f
C699 B.n526 VSUBS 0.007233f
C700 B.n527 VSUBS 0.007233f
C701 B.n528 VSUBS 0.007233f
C702 B.n529 VSUBS 0.007233f
C703 B.n530 VSUBS 0.007233f
C704 B.n531 VSUBS 0.007233f
C705 B.n532 VSUBS 0.007233f
C706 B.n533 VSUBS 0.007233f
C707 B.n534 VSUBS 0.007233f
C708 B.n535 VSUBS 0.007233f
C709 B.n536 VSUBS 0.007233f
C710 B.n537 VSUBS 0.007233f
C711 B.n538 VSUBS 0.007233f
C712 B.n539 VSUBS 0.007233f
C713 B.n540 VSUBS 0.007233f
C714 B.n541 VSUBS 0.007233f
C715 B.n542 VSUBS 0.007233f
C716 B.n543 VSUBS 0.007233f
C717 B.n544 VSUBS 0.007233f
C718 B.n545 VSUBS 0.007233f
C719 B.n546 VSUBS 0.007233f
C720 B.n547 VSUBS 0.007233f
C721 B.n548 VSUBS 0.007233f
C722 B.n549 VSUBS 0.007233f
C723 B.n550 VSUBS 0.007233f
C724 B.n551 VSUBS 0.007233f
C725 B.n552 VSUBS 0.007233f
C726 B.n553 VSUBS 0.007233f
C727 B.n554 VSUBS 0.007233f
C728 B.n555 VSUBS 0.007233f
C729 B.n556 VSUBS 0.007233f
C730 B.n557 VSUBS 0.007233f
C731 B.n558 VSUBS 0.007233f
C732 B.n559 VSUBS 0.007233f
C733 B.n560 VSUBS 0.007233f
C734 B.n561 VSUBS 0.007233f
C735 B.n562 VSUBS 0.007233f
C736 B.n563 VSUBS 0.007233f
C737 B.n564 VSUBS 0.007233f
C738 B.n565 VSUBS 0.007233f
C739 B.n566 VSUBS 0.007233f
C740 B.n567 VSUBS 0.007233f
C741 B.n568 VSUBS 0.007233f
C742 B.n569 VSUBS 0.007233f
C743 B.n570 VSUBS 0.007233f
C744 B.n571 VSUBS 0.007233f
C745 B.n572 VSUBS 0.007233f
C746 B.n573 VSUBS 0.007233f
C747 B.n574 VSUBS 0.007233f
C748 B.n575 VSUBS 0.007233f
C749 B.n576 VSUBS 0.007233f
C750 B.n577 VSUBS 0.007233f
C751 B.n578 VSUBS 0.007233f
C752 B.n579 VSUBS 0.007233f
C753 B.n580 VSUBS 0.007233f
C754 B.n581 VSUBS 0.007233f
C755 B.n582 VSUBS 0.007233f
C756 B.n583 VSUBS 0.007233f
C757 B.n584 VSUBS 0.007233f
C758 B.n585 VSUBS 0.007233f
C759 B.n586 VSUBS 0.007233f
C760 B.n587 VSUBS 0.007233f
C761 B.n588 VSUBS 0.007233f
C762 B.n589 VSUBS 0.007233f
C763 B.n590 VSUBS 0.007233f
C764 B.n591 VSUBS 0.007233f
C765 B.n592 VSUBS 0.007233f
C766 B.n593 VSUBS 0.007233f
C767 B.n594 VSUBS 0.007233f
C768 B.n595 VSUBS 0.007233f
C769 B.n596 VSUBS 0.007233f
C770 B.n597 VSUBS 0.017264f
C771 B.n598 VSUBS 0.017264f
C772 B.n599 VSUBS 0.017836f
C773 B.n600 VSUBS 0.007233f
C774 B.n601 VSUBS 0.007233f
C775 B.n602 VSUBS 0.007233f
C776 B.n603 VSUBS 0.007233f
C777 B.n604 VSUBS 0.007233f
C778 B.n605 VSUBS 0.007233f
C779 B.n606 VSUBS 0.007233f
C780 B.n607 VSUBS 0.007233f
C781 B.n608 VSUBS 0.007233f
C782 B.n609 VSUBS 0.007233f
C783 B.n610 VSUBS 0.007233f
C784 B.n611 VSUBS 0.007233f
C785 B.n612 VSUBS 0.007233f
C786 B.n613 VSUBS 0.007233f
C787 B.n614 VSUBS 0.007233f
C788 B.n615 VSUBS 0.007233f
C789 B.n616 VSUBS 0.007233f
C790 B.n617 VSUBS 0.007233f
C791 B.n618 VSUBS 0.007233f
C792 B.n619 VSUBS 0.007233f
C793 B.n620 VSUBS 0.007233f
C794 B.n621 VSUBS 0.007233f
C795 B.n622 VSUBS 0.007233f
C796 B.n623 VSUBS 0.007233f
C797 B.n624 VSUBS 0.007233f
C798 B.n625 VSUBS 0.007233f
C799 B.n626 VSUBS 0.007233f
C800 B.n627 VSUBS 0.007233f
C801 B.n628 VSUBS 0.007233f
C802 B.n629 VSUBS 0.007233f
C803 B.n630 VSUBS 0.007233f
C804 B.n631 VSUBS 0.007233f
C805 B.n632 VSUBS 0.007233f
C806 B.n633 VSUBS 0.007233f
C807 B.n634 VSUBS 0.007233f
C808 B.n635 VSUBS 0.007233f
C809 B.n636 VSUBS 0.007233f
C810 B.n637 VSUBS 0.007233f
C811 B.n638 VSUBS 0.007233f
C812 B.n639 VSUBS 0.007233f
C813 B.n640 VSUBS 0.007233f
C814 B.n641 VSUBS 0.007233f
C815 B.n642 VSUBS 0.007233f
C816 B.n643 VSUBS 0.007233f
C817 B.n644 VSUBS 0.007233f
C818 B.n645 VSUBS 0.007233f
C819 B.n646 VSUBS 0.007233f
C820 B.n647 VSUBS 0.007233f
C821 B.n648 VSUBS 0.007233f
C822 B.n649 VSUBS 0.007233f
C823 B.n650 VSUBS 0.007233f
C824 B.n651 VSUBS 0.007233f
C825 B.n652 VSUBS 0.007233f
C826 B.n653 VSUBS 0.007233f
C827 B.n654 VSUBS 0.007233f
C828 B.n655 VSUBS 0.007233f
C829 B.n656 VSUBS 0.007233f
C830 B.n657 VSUBS 0.007233f
C831 B.n658 VSUBS 0.007233f
C832 B.n659 VSUBS 0.007233f
C833 B.n660 VSUBS 0.007233f
C834 B.n661 VSUBS 0.007233f
C835 B.n662 VSUBS 0.007233f
C836 B.n663 VSUBS 0.007233f
C837 B.n664 VSUBS 0.007233f
C838 B.n665 VSUBS 0.007233f
C839 B.n666 VSUBS 0.007233f
C840 B.n667 VSUBS 0.007233f
C841 B.n668 VSUBS 0.007233f
C842 B.n669 VSUBS 0.007233f
C843 B.n670 VSUBS 0.007233f
C844 B.n671 VSUBS 0.007233f
C845 B.n672 VSUBS 0.007233f
C846 B.n673 VSUBS 0.007233f
C847 B.n674 VSUBS 0.007233f
C848 B.n675 VSUBS 0.007233f
C849 B.n676 VSUBS 0.007233f
C850 B.n677 VSUBS 0.007233f
C851 B.n678 VSUBS 0.007233f
C852 B.n679 VSUBS 0.007233f
C853 B.n680 VSUBS 0.007233f
C854 B.n681 VSUBS 0.007233f
C855 B.n682 VSUBS 0.007233f
C856 B.n683 VSUBS 0.007233f
C857 B.n684 VSUBS 0.007233f
C858 B.n685 VSUBS 0.007233f
C859 B.n686 VSUBS 0.004999f
C860 B.n687 VSUBS 0.016758f
C861 B.n688 VSUBS 0.00585f
C862 B.n689 VSUBS 0.007233f
C863 B.n690 VSUBS 0.007233f
C864 B.n691 VSUBS 0.007233f
C865 B.n692 VSUBS 0.007233f
C866 B.n693 VSUBS 0.007233f
C867 B.n694 VSUBS 0.007233f
C868 B.n695 VSUBS 0.007233f
C869 B.n696 VSUBS 0.007233f
C870 B.n697 VSUBS 0.007233f
C871 B.n698 VSUBS 0.007233f
C872 B.n699 VSUBS 0.007233f
C873 B.n700 VSUBS 0.00585f
C874 B.n701 VSUBS 0.007233f
C875 B.n702 VSUBS 0.007233f
C876 B.n703 VSUBS 0.004999f
C877 B.n704 VSUBS 0.007233f
C878 B.n705 VSUBS 0.007233f
C879 B.n706 VSUBS 0.007233f
C880 B.n707 VSUBS 0.007233f
C881 B.n708 VSUBS 0.007233f
C882 B.n709 VSUBS 0.007233f
C883 B.n710 VSUBS 0.007233f
C884 B.n711 VSUBS 0.007233f
C885 B.n712 VSUBS 0.007233f
C886 B.n713 VSUBS 0.007233f
C887 B.n714 VSUBS 0.007233f
C888 B.n715 VSUBS 0.007233f
C889 B.n716 VSUBS 0.007233f
C890 B.n717 VSUBS 0.007233f
C891 B.n718 VSUBS 0.007233f
C892 B.n719 VSUBS 0.007233f
C893 B.n720 VSUBS 0.007233f
C894 B.n721 VSUBS 0.007233f
C895 B.n722 VSUBS 0.007233f
C896 B.n723 VSUBS 0.007233f
C897 B.n724 VSUBS 0.007233f
C898 B.n725 VSUBS 0.007233f
C899 B.n726 VSUBS 0.007233f
C900 B.n727 VSUBS 0.007233f
C901 B.n728 VSUBS 0.007233f
C902 B.n729 VSUBS 0.007233f
C903 B.n730 VSUBS 0.007233f
C904 B.n731 VSUBS 0.007233f
C905 B.n732 VSUBS 0.007233f
C906 B.n733 VSUBS 0.007233f
C907 B.n734 VSUBS 0.007233f
C908 B.n735 VSUBS 0.007233f
C909 B.n736 VSUBS 0.007233f
C910 B.n737 VSUBS 0.007233f
C911 B.n738 VSUBS 0.007233f
C912 B.n739 VSUBS 0.007233f
C913 B.n740 VSUBS 0.007233f
C914 B.n741 VSUBS 0.007233f
C915 B.n742 VSUBS 0.007233f
C916 B.n743 VSUBS 0.007233f
C917 B.n744 VSUBS 0.007233f
C918 B.n745 VSUBS 0.007233f
C919 B.n746 VSUBS 0.007233f
C920 B.n747 VSUBS 0.007233f
C921 B.n748 VSUBS 0.007233f
C922 B.n749 VSUBS 0.007233f
C923 B.n750 VSUBS 0.007233f
C924 B.n751 VSUBS 0.007233f
C925 B.n752 VSUBS 0.007233f
C926 B.n753 VSUBS 0.007233f
C927 B.n754 VSUBS 0.007233f
C928 B.n755 VSUBS 0.007233f
C929 B.n756 VSUBS 0.007233f
C930 B.n757 VSUBS 0.007233f
C931 B.n758 VSUBS 0.007233f
C932 B.n759 VSUBS 0.007233f
C933 B.n760 VSUBS 0.007233f
C934 B.n761 VSUBS 0.007233f
C935 B.n762 VSUBS 0.007233f
C936 B.n763 VSUBS 0.007233f
C937 B.n764 VSUBS 0.007233f
C938 B.n765 VSUBS 0.007233f
C939 B.n766 VSUBS 0.007233f
C940 B.n767 VSUBS 0.007233f
C941 B.n768 VSUBS 0.007233f
C942 B.n769 VSUBS 0.007233f
C943 B.n770 VSUBS 0.007233f
C944 B.n771 VSUBS 0.007233f
C945 B.n772 VSUBS 0.007233f
C946 B.n773 VSUBS 0.007233f
C947 B.n774 VSUBS 0.007233f
C948 B.n775 VSUBS 0.007233f
C949 B.n776 VSUBS 0.007233f
C950 B.n777 VSUBS 0.007233f
C951 B.n778 VSUBS 0.007233f
C952 B.n779 VSUBS 0.007233f
C953 B.n780 VSUBS 0.007233f
C954 B.n781 VSUBS 0.007233f
C955 B.n782 VSUBS 0.007233f
C956 B.n783 VSUBS 0.007233f
C957 B.n784 VSUBS 0.007233f
C958 B.n785 VSUBS 0.007233f
C959 B.n786 VSUBS 0.007233f
C960 B.n787 VSUBS 0.007233f
C961 B.n788 VSUBS 0.007233f
C962 B.n789 VSUBS 0.017836f
C963 B.n790 VSUBS 0.017836f
C964 B.n791 VSUBS 0.017264f
C965 B.n792 VSUBS 0.007233f
C966 B.n793 VSUBS 0.007233f
C967 B.n794 VSUBS 0.007233f
C968 B.n795 VSUBS 0.007233f
C969 B.n796 VSUBS 0.007233f
C970 B.n797 VSUBS 0.007233f
C971 B.n798 VSUBS 0.007233f
C972 B.n799 VSUBS 0.007233f
C973 B.n800 VSUBS 0.007233f
C974 B.n801 VSUBS 0.007233f
C975 B.n802 VSUBS 0.007233f
C976 B.n803 VSUBS 0.007233f
C977 B.n804 VSUBS 0.007233f
C978 B.n805 VSUBS 0.007233f
C979 B.n806 VSUBS 0.007233f
C980 B.n807 VSUBS 0.007233f
C981 B.n808 VSUBS 0.007233f
C982 B.n809 VSUBS 0.007233f
C983 B.n810 VSUBS 0.007233f
C984 B.n811 VSUBS 0.007233f
C985 B.n812 VSUBS 0.007233f
C986 B.n813 VSUBS 0.007233f
C987 B.n814 VSUBS 0.007233f
C988 B.n815 VSUBS 0.007233f
C989 B.n816 VSUBS 0.007233f
C990 B.n817 VSUBS 0.007233f
C991 B.n818 VSUBS 0.007233f
C992 B.n819 VSUBS 0.007233f
C993 B.n820 VSUBS 0.007233f
C994 B.n821 VSUBS 0.007233f
C995 B.n822 VSUBS 0.007233f
C996 B.n823 VSUBS 0.007233f
C997 B.n824 VSUBS 0.007233f
C998 B.n825 VSUBS 0.007233f
C999 B.n826 VSUBS 0.007233f
C1000 B.n827 VSUBS 0.007233f
C1001 B.n828 VSUBS 0.007233f
C1002 B.n829 VSUBS 0.007233f
C1003 B.n830 VSUBS 0.007233f
C1004 B.n831 VSUBS 0.007233f
C1005 B.n832 VSUBS 0.007233f
C1006 B.n833 VSUBS 0.007233f
C1007 B.n834 VSUBS 0.007233f
C1008 B.n835 VSUBS 0.007233f
C1009 B.n836 VSUBS 0.007233f
C1010 B.n837 VSUBS 0.007233f
C1011 B.n838 VSUBS 0.007233f
C1012 B.n839 VSUBS 0.007233f
C1013 B.n840 VSUBS 0.007233f
C1014 B.n841 VSUBS 0.007233f
C1015 B.n842 VSUBS 0.007233f
C1016 B.n843 VSUBS 0.007233f
C1017 B.n844 VSUBS 0.007233f
C1018 B.n845 VSUBS 0.007233f
C1019 B.n846 VSUBS 0.007233f
C1020 B.n847 VSUBS 0.007233f
C1021 B.n848 VSUBS 0.007233f
C1022 B.n849 VSUBS 0.007233f
C1023 B.n850 VSUBS 0.007233f
C1024 B.n851 VSUBS 0.009438f
C1025 B.n852 VSUBS 0.010054f
C1026 B.n853 VSUBS 0.019994f
.ends

