* NGSPICE file created from diff_pair_sample_0983.ext - technology: sky130A

.subckt diff_pair_sample_0983 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t19 VN.t0 VDD2.t3 B.t4 sky130_fd_pr__nfet_01v8 ad=2.9106 pd=17.97 as=2.9106 ps=17.97 w=17.64 l=1.48
X1 VDD1.t9 VP.t0 VTAIL.t8 B.t8 sky130_fd_pr__nfet_01v8 ad=2.9106 pd=17.97 as=6.8796 ps=36.06 w=17.64 l=1.48
X2 B.t23 B.t21 B.t22 B.t11 sky130_fd_pr__nfet_01v8 ad=6.8796 pd=36.06 as=0 ps=0 w=17.64 l=1.48
X3 VTAIL.t9 VP.t1 VDD1.t8 B.t9 sky130_fd_pr__nfet_01v8 ad=2.9106 pd=17.97 as=2.9106 ps=17.97 w=17.64 l=1.48
X4 VDD2.t2 VN.t1 VTAIL.t18 B.t7 sky130_fd_pr__nfet_01v8 ad=6.8796 pd=36.06 as=2.9106 ps=17.97 w=17.64 l=1.48
X5 VTAIL.t4 VP.t2 VDD1.t7 B.t4 sky130_fd_pr__nfet_01v8 ad=2.9106 pd=17.97 as=2.9106 ps=17.97 w=17.64 l=1.48
X6 VDD2.t7 VN.t2 VTAIL.t17 B.t8 sky130_fd_pr__nfet_01v8 ad=2.9106 pd=17.97 as=6.8796 ps=36.06 w=17.64 l=1.48
X7 B.t20 B.t18 B.t19 B.t15 sky130_fd_pr__nfet_01v8 ad=6.8796 pd=36.06 as=0 ps=0 w=17.64 l=1.48
X8 VDD1.t6 VP.t3 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=2.9106 pd=17.97 as=2.9106 ps=17.97 w=17.64 l=1.48
X9 B.t17 B.t14 B.t16 B.t15 sky130_fd_pr__nfet_01v8 ad=6.8796 pd=36.06 as=0 ps=0 w=17.64 l=1.48
X10 B.t13 B.t10 B.t12 B.t11 sky130_fd_pr__nfet_01v8 ad=6.8796 pd=36.06 as=0 ps=0 w=17.64 l=1.48
X11 VDD2.t6 VN.t3 VTAIL.t16 B.t6 sky130_fd_pr__nfet_01v8 ad=2.9106 pd=17.97 as=2.9106 ps=17.97 w=17.64 l=1.48
X12 VTAIL.t15 VN.t4 VDD2.t9 B.t9 sky130_fd_pr__nfet_01v8 ad=2.9106 pd=17.97 as=2.9106 ps=17.97 w=17.64 l=1.48
X13 VDD1.t5 VP.t4 VTAIL.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=6.8796 pd=36.06 as=2.9106 ps=17.97 w=17.64 l=1.48
X14 VDD2.t8 VN.t5 VTAIL.t14 B.t2 sky130_fd_pr__nfet_01v8 ad=2.9106 pd=17.97 as=6.8796 ps=36.06 w=17.64 l=1.48
X15 VDD1.t4 VP.t5 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=2.9106 pd=17.97 as=6.8796 ps=36.06 w=17.64 l=1.48
X16 VTAIL.t3 VP.t6 VDD1.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=2.9106 pd=17.97 as=2.9106 ps=17.97 w=17.64 l=1.48
X17 VDD2.t1 VN.t6 VTAIL.t13 B.t0 sky130_fd_pr__nfet_01v8 ad=2.9106 pd=17.97 as=2.9106 ps=17.97 w=17.64 l=1.48
X18 VTAIL.t12 VN.t7 VDD2.t0 B.t3 sky130_fd_pr__nfet_01v8 ad=2.9106 pd=17.97 as=2.9106 ps=17.97 w=17.64 l=1.48
X19 VTAIL.t11 VN.t8 VDD2.t5 B.t1 sky130_fd_pr__nfet_01v8 ad=2.9106 pd=17.97 as=2.9106 ps=17.97 w=17.64 l=1.48
X20 VTAIL.t1 VP.t7 VDD1.t2 B.t1 sky130_fd_pr__nfet_01v8 ad=2.9106 pd=17.97 as=2.9106 ps=17.97 w=17.64 l=1.48
X21 VDD2.t4 VN.t9 VTAIL.t10 B.t5 sky130_fd_pr__nfet_01v8 ad=6.8796 pd=36.06 as=2.9106 ps=17.97 w=17.64 l=1.48
X22 VDD1.t1 VP.t8 VTAIL.t6 B.t6 sky130_fd_pr__nfet_01v8 ad=2.9106 pd=17.97 as=2.9106 ps=17.97 w=17.64 l=1.48
X23 VDD1.t0 VP.t9 VTAIL.t7 B.t7 sky130_fd_pr__nfet_01v8 ad=6.8796 pd=36.06 as=2.9106 ps=17.97 w=17.64 l=1.48
R0 VN.n7 VN.t1 318.837
R1 VN.n34 VN.t5 318.837
R2 VN.n12 VN.t3 287.247
R3 VN.n6 VN.t8 287.247
R4 VN.n18 VN.t4 287.247
R5 VN.n25 VN.t2 287.247
R6 VN.n39 VN.t6 287.247
R7 VN.n33 VN.t7 287.247
R8 VN.n45 VN.t0 287.247
R9 VN.n52 VN.t9 287.247
R10 VN.n26 VN.n25 179.99
R11 VN.n53 VN.n52 179.99
R12 VN.n51 VN.n27 161.3
R13 VN.n50 VN.n49 161.3
R14 VN.n48 VN.n28 161.3
R15 VN.n47 VN.n46 161.3
R16 VN.n44 VN.n29 161.3
R17 VN.n43 VN.n42 161.3
R18 VN.n41 VN.n30 161.3
R19 VN.n40 VN.n39 161.3
R20 VN.n38 VN.n31 161.3
R21 VN.n37 VN.n36 161.3
R22 VN.n35 VN.n32 161.3
R23 VN.n24 VN.n0 161.3
R24 VN.n23 VN.n22 161.3
R25 VN.n21 VN.n1 161.3
R26 VN.n20 VN.n19 161.3
R27 VN.n17 VN.n2 161.3
R28 VN.n16 VN.n15 161.3
R29 VN.n14 VN.n3 161.3
R30 VN.n13 VN.n12 161.3
R31 VN.n11 VN.n4 161.3
R32 VN.n10 VN.n9 161.3
R33 VN.n8 VN.n5 161.3
R34 VN.n23 VN.n1 56.5617
R35 VN.n50 VN.n28 56.5617
R36 VN VN.n53 51.5365
R37 VN.n7 VN.n6 50.9283
R38 VN.n34 VN.n33 50.9283
R39 VN.n11 VN.n10 49.7803
R40 VN.n16 VN.n3 49.7803
R41 VN.n38 VN.n37 49.7803
R42 VN.n43 VN.n30 49.7803
R43 VN.n10 VN.n5 31.3737
R44 VN.n17 VN.n16 31.3737
R45 VN.n37 VN.n32 31.3737
R46 VN.n44 VN.n43 31.3737
R47 VN.n12 VN.n11 24.5923
R48 VN.n12 VN.n3 24.5923
R49 VN.n19 VN.n1 24.5923
R50 VN.n24 VN.n23 24.5923
R51 VN.n39 VN.n30 24.5923
R52 VN.n39 VN.n38 24.5923
R53 VN.n46 VN.n28 24.5923
R54 VN.n51 VN.n50 24.5923
R55 VN.n35 VN.n34 18.1684
R56 VN.n8 VN.n7 18.1684
R57 VN.n6 VN.n5 15.2474
R58 VN.n18 VN.n17 15.2474
R59 VN.n33 VN.n32 15.2474
R60 VN.n45 VN.n44 15.2474
R61 VN.n19 VN.n18 9.3454
R62 VN.n46 VN.n45 9.3454
R63 VN.n25 VN.n24 5.90254
R64 VN.n52 VN.n51 5.90254
R65 VN.n53 VN.n27 0.189894
R66 VN.n49 VN.n27 0.189894
R67 VN.n49 VN.n48 0.189894
R68 VN.n48 VN.n47 0.189894
R69 VN.n47 VN.n29 0.189894
R70 VN.n42 VN.n29 0.189894
R71 VN.n42 VN.n41 0.189894
R72 VN.n41 VN.n40 0.189894
R73 VN.n40 VN.n31 0.189894
R74 VN.n36 VN.n31 0.189894
R75 VN.n36 VN.n35 0.189894
R76 VN.n9 VN.n8 0.189894
R77 VN.n9 VN.n4 0.189894
R78 VN.n13 VN.n4 0.189894
R79 VN.n14 VN.n13 0.189894
R80 VN.n15 VN.n14 0.189894
R81 VN.n15 VN.n2 0.189894
R82 VN.n20 VN.n2 0.189894
R83 VN.n21 VN.n20 0.189894
R84 VN.n22 VN.n21 0.189894
R85 VN.n22 VN.n0 0.189894
R86 VN.n26 VN.n0 0.189894
R87 VN VN.n26 0.0516364
R88 VDD2.n193 VDD2.n101 289.615
R89 VDD2.n92 VDD2.n0 289.615
R90 VDD2.n194 VDD2.n193 185
R91 VDD2.n192 VDD2.n191 185
R92 VDD2.n105 VDD2.n104 185
R93 VDD2.n186 VDD2.n185 185
R94 VDD2.n184 VDD2.n183 185
R95 VDD2.n109 VDD2.n108 185
R96 VDD2.n113 VDD2.n111 185
R97 VDD2.n178 VDD2.n177 185
R98 VDD2.n176 VDD2.n175 185
R99 VDD2.n115 VDD2.n114 185
R100 VDD2.n170 VDD2.n169 185
R101 VDD2.n168 VDD2.n167 185
R102 VDD2.n119 VDD2.n118 185
R103 VDD2.n162 VDD2.n161 185
R104 VDD2.n160 VDD2.n159 185
R105 VDD2.n123 VDD2.n122 185
R106 VDD2.n154 VDD2.n153 185
R107 VDD2.n152 VDD2.n151 185
R108 VDD2.n127 VDD2.n126 185
R109 VDD2.n146 VDD2.n145 185
R110 VDD2.n144 VDD2.n143 185
R111 VDD2.n131 VDD2.n130 185
R112 VDD2.n138 VDD2.n137 185
R113 VDD2.n136 VDD2.n135 185
R114 VDD2.n33 VDD2.n32 185
R115 VDD2.n35 VDD2.n34 185
R116 VDD2.n28 VDD2.n27 185
R117 VDD2.n41 VDD2.n40 185
R118 VDD2.n43 VDD2.n42 185
R119 VDD2.n24 VDD2.n23 185
R120 VDD2.n49 VDD2.n48 185
R121 VDD2.n51 VDD2.n50 185
R122 VDD2.n20 VDD2.n19 185
R123 VDD2.n57 VDD2.n56 185
R124 VDD2.n59 VDD2.n58 185
R125 VDD2.n16 VDD2.n15 185
R126 VDD2.n65 VDD2.n64 185
R127 VDD2.n67 VDD2.n66 185
R128 VDD2.n12 VDD2.n11 185
R129 VDD2.n74 VDD2.n73 185
R130 VDD2.n75 VDD2.n10 185
R131 VDD2.n77 VDD2.n76 185
R132 VDD2.n8 VDD2.n7 185
R133 VDD2.n83 VDD2.n82 185
R134 VDD2.n85 VDD2.n84 185
R135 VDD2.n4 VDD2.n3 185
R136 VDD2.n91 VDD2.n90 185
R137 VDD2.n93 VDD2.n92 185
R138 VDD2.n134 VDD2.t4 147.659
R139 VDD2.n31 VDD2.t2 147.659
R140 VDD2.n193 VDD2.n192 104.615
R141 VDD2.n192 VDD2.n104 104.615
R142 VDD2.n185 VDD2.n104 104.615
R143 VDD2.n185 VDD2.n184 104.615
R144 VDD2.n184 VDD2.n108 104.615
R145 VDD2.n113 VDD2.n108 104.615
R146 VDD2.n177 VDD2.n113 104.615
R147 VDD2.n177 VDD2.n176 104.615
R148 VDD2.n176 VDD2.n114 104.615
R149 VDD2.n169 VDD2.n114 104.615
R150 VDD2.n169 VDD2.n168 104.615
R151 VDD2.n168 VDD2.n118 104.615
R152 VDD2.n161 VDD2.n118 104.615
R153 VDD2.n161 VDD2.n160 104.615
R154 VDD2.n160 VDD2.n122 104.615
R155 VDD2.n153 VDD2.n122 104.615
R156 VDD2.n153 VDD2.n152 104.615
R157 VDD2.n152 VDD2.n126 104.615
R158 VDD2.n145 VDD2.n126 104.615
R159 VDD2.n145 VDD2.n144 104.615
R160 VDD2.n144 VDD2.n130 104.615
R161 VDD2.n137 VDD2.n130 104.615
R162 VDD2.n137 VDD2.n136 104.615
R163 VDD2.n34 VDD2.n33 104.615
R164 VDD2.n34 VDD2.n27 104.615
R165 VDD2.n41 VDD2.n27 104.615
R166 VDD2.n42 VDD2.n41 104.615
R167 VDD2.n42 VDD2.n23 104.615
R168 VDD2.n49 VDD2.n23 104.615
R169 VDD2.n50 VDD2.n49 104.615
R170 VDD2.n50 VDD2.n19 104.615
R171 VDD2.n57 VDD2.n19 104.615
R172 VDD2.n58 VDD2.n57 104.615
R173 VDD2.n58 VDD2.n15 104.615
R174 VDD2.n65 VDD2.n15 104.615
R175 VDD2.n66 VDD2.n65 104.615
R176 VDD2.n66 VDD2.n11 104.615
R177 VDD2.n74 VDD2.n11 104.615
R178 VDD2.n75 VDD2.n74 104.615
R179 VDD2.n76 VDD2.n75 104.615
R180 VDD2.n76 VDD2.n7 104.615
R181 VDD2.n83 VDD2.n7 104.615
R182 VDD2.n84 VDD2.n83 104.615
R183 VDD2.n84 VDD2.n3 104.615
R184 VDD2.n91 VDD2.n3 104.615
R185 VDD2.n92 VDD2.n91 104.615
R186 VDD2.n100 VDD2.n99 64.1242
R187 VDD2 VDD2.n201 64.1213
R188 VDD2.n200 VDD2.n199 63.0094
R189 VDD2.n98 VDD2.n97 63.0093
R190 VDD2.n98 VDD2.n96 52.7518
R191 VDD2.n136 VDD2.t4 52.3082
R192 VDD2.n33 VDD2.t2 52.3082
R193 VDD2.n198 VDD2.n197 51.1914
R194 VDD2.n198 VDD2.n100 46.3338
R195 VDD2.n135 VDD2.n134 15.6677
R196 VDD2.n32 VDD2.n31 15.6677
R197 VDD2.n111 VDD2.n109 13.1884
R198 VDD2.n77 VDD2.n8 13.1884
R199 VDD2.n183 VDD2.n182 12.8005
R200 VDD2.n179 VDD2.n178 12.8005
R201 VDD2.n138 VDD2.n133 12.8005
R202 VDD2.n35 VDD2.n30 12.8005
R203 VDD2.n78 VDD2.n10 12.8005
R204 VDD2.n82 VDD2.n81 12.8005
R205 VDD2.n186 VDD2.n107 12.0247
R206 VDD2.n175 VDD2.n112 12.0247
R207 VDD2.n139 VDD2.n131 12.0247
R208 VDD2.n36 VDD2.n28 12.0247
R209 VDD2.n73 VDD2.n72 12.0247
R210 VDD2.n85 VDD2.n6 12.0247
R211 VDD2.n187 VDD2.n105 11.249
R212 VDD2.n174 VDD2.n115 11.249
R213 VDD2.n143 VDD2.n142 11.249
R214 VDD2.n40 VDD2.n39 11.249
R215 VDD2.n71 VDD2.n12 11.249
R216 VDD2.n86 VDD2.n4 11.249
R217 VDD2.n191 VDD2.n190 10.4732
R218 VDD2.n171 VDD2.n170 10.4732
R219 VDD2.n146 VDD2.n129 10.4732
R220 VDD2.n43 VDD2.n26 10.4732
R221 VDD2.n68 VDD2.n67 10.4732
R222 VDD2.n90 VDD2.n89 10.4732
R223 VDD2.n194 VDD2.n103 9.69747
R224 VDD2.n167 VDD2.n117 9.69747
R225 VDD2.n147 VDD2.n127 9.69747
R226 VDD2.n44 VDD2.n24 9.69747
R227 VDD2.n64 VDD2.n14 9.69747
R228 VDD2.n93 VDD2.n2 9.69747
R229 VDD2.n197 VDD2.n196 9.45567
R230 VDD2.n96 VDD2.n95 9.45567
R231 VDD2.n121 VDD2.n120 9.3005
R232 VDD2.n164 VDD2.n163 9.3005
R233 VDD2.n166 VDD2.n165 9.3005
R234 VDD2.n117 VDD2.n116 9.3005
R235 VDD2.n172 VDD2.n171 9.3005
R236 VDD2.n174 VDD2.n173 9.3005
R237 VDD2.n112 VDD2.n110 9.3005
R238 VDD2.n180 VDD2.n179 9.3005
R239 VDD2.n196 VDD2.n195 9.3005
R240 VDD2.n103 VDD2.n102 9.3005
R241 VDD2.n190 VDD2.n189 9.3005
R242 VDD2.n188 VDD2.n187 9.3005
R243 VDD2.n107 VDD2.n106 9.3005
R244 VDD2.n182 VDD2.n181 9.3005
R245 VDD2.n158 VDD2.n157 9.3005
R246 VDD2.n156 VDD2.n155 9.3005
R247 VDD2.n125 VDD2.n124 9.3005
R248 VDD2.n150 VDD2.n149 9.3005
R249 VDD2.n148 VDD2.n147 9.3005
R250 VDD2.n129 VDD2.n128 9.3005
R251 VDD2.n142 VDD2.n141 9.3005
R252 VDD2.n140 VDD2.n139 9.3005
R253 VDD2.n133 VDD2.n132 9.3005
R254 VDD2.n95 VDD2.n94 9.3005
R255 VDD2.n2 VDD2.n1 9.3005
R256 VDD2.n89 VDD2.n88 9.3005
R257 VDD2.n87 VDD2.n86 9.3005
R258 VDD2.n6 VDD2.n5 9.3005
R259 VDD2.n81 VDD2.n80 9.3005
R260 VDD2.n53 VDD2.n52 9.3005
R261 VDD2.n22 VDD2.n21 9.3005
R262 VDD2.n47 VDD2.n46 9.3005
R263 VDD2.n45 VDD2.n44 9.3005
R264 VDD2.n26 VDD2.n25 9.3005
R265 VDD2.n39 VDD2.n38 9.3005
R266 VDD2.n37 VDD2.n36 9.3005
R267 VDD2.n30 VDD2.n29 9.3005
R268 VDD2.n55 VDD2.n54 9.3005
R269 VDD2.n18 VDD2.n17 9.3005
R270 VDD2.n61 VDD2.n60 9.3005
R271 VDD2.n63 VDD2.n62 9.3005
R272 VDD2.n14 VDD2.n13 9.3005
R273 VDD2.n69 VDD2.n68 9.3005
R274 VDD2.n71 VDD2.n70 9.3005
R275 VDD2.n72 VDD2.n9 9.3005
R276 VDD2.n79 VDD2.n78 9.3005
R277 VDD2.n195 VDD2.n101 8.92171
R278 VDD2.n166 VDD2.n119 8.92171
R279 VDD2.n151 VDD2.n150 8.92171
R280 VDD2.n48 VDD2.n47 8.92171
R281 VDD2.n63 VDD2.n16 8.92171
R282 VDD2.n94 VDD2.n0 8.92171
R283 VDD2.n163 VDD2.n162 8.14595
R284 VDD2.n154 VDD2.n125 8.14595
R285 VDD2.n51 VDD2.n22 8.14595
R286 VDD2.n60 VDD2.n59 8.14595
R287 VDD2.n159 VDD2.n121 7.3702
R288 VDD2.n155 VDD2.n123 7.3702
R289 VDD2.n52 VDD2.n20 7.3702
R290 VDD2.n56 VDD2.n18 7.3702
R291 VDD2.n159 VDD2.n158 6.59444
R292 VDD2.n158 VDD2.n123 6.59444
R293 VDD2.n55 VDD2.n20 6.59444
R294 VDD2.n56 VDD2.n55 6.59444
R295 VDD2.n162 VDD2.n121 5.81868
R296 VDD2.n155 VDD2.n154 5.81868
R297 VDD2.n52 VDD2.n51 5.81868
R298 VDD2.n59 VDD2.n18 5.81868
R299 VDD2.n197 VDD2.n101 5.04292
R300 VDD2.n163 VDD2.n119 5.04292
R301 VDD2.n151 VDD2.n125 5.04292
R302 VDD2.n48 VDD2.n22 5.04292
R303 VDD2.n60 VDD2.n16 5.04292
R304 VDD2.n96 VDD2.n0 5.04292
R305 VDD2.n134 VDD2.n132 4.38563
R306 VDD2.n31 VDD2.n29 4.38563
R307 VDD2.n195 VDD2.n194 4.26717
R308 VDD2.n167 VDD2.n166 4.26717
R309 VDD2.n150 VDD2.n127 4.26717
R310 VDD2.n47 VDD2.n24 4.26717
R311 VDD2.n64 VDD2.n63 4.26717
R312 VDD2.n94 VDD2.n93 4.26717
R313 VDD2.n191 VDD2.n103 3.49141
R314 VDD2.n170 VDD2.n117 3.49141
R315 VDD2.n147 VDD2.n146 3.49141
R316 VDD2.n44 VDD2.n43 3.49141
R317 VDD2.n67 VDD2.n14 3.49141
R318 VDD2.n90 VDD2.n2 3.49141
R319 VDD2.n190 VDD2.n105 2.71565
R320 VDD2.n171 VDD2.n115 2.71565
R321 VDD2.n143 VDD2.n129 2.71565
R322 VDD2.n40 VDD2.n26 2.71565
R323 VDD2.n68 VDD2.n12 2.71565
R324 VDD2.n89 VDD2.n4 2.71565
R325 VDD2.n187 VDD2.n186 1.93989
R326 VDD2.n175 VDD2.n174 1.93989
R327 VDD2.n142 VDD2.n131 1.93989
R328 VDD2.n39 VDD2.n28 1.93989
R329 VDD2.n73 VDD2.n71 1.93989
R330 VDD2.n86 VDD2.n85 1.93989
R331 VDD2.n200 VDD2.n198 1.56084
R332 VDD2.n183 VDD2.n107 1.16414
R333 VDD2.n178 VDD2.n112 1.16414
R334 VDD2.n139 VDD2.n138 1.16414
R335 VDD2.n36 VDD2.n35 1.16414
R336 VDD2.n72 VDD2.n10 1.16414
R337 VDD2.n82 VDD2.n6 1.16414
R338 VDD2.n201 VDD2.t0 1.12295
R339 VDD2.n201 VDD2.t8 1.12295
R340 VDD2.n199 VDD2.t3 1.12295
R341 VDD2.n199 VDD2.t1 1.12295
R342 VDD2.n99 VDD2.t9 1.12295
R343 VDD2.n99 VDD2.t7 1.12295
R344 VDD2.n97 VDD2.t5 1.12295
R345 VDD2.n97 VDD2.t6 1.12295
R346 VDD2 VDD2.n200 0.448776
R347 VDD2.n182 VDD2.n109 0.388379
R348 VDD2.n179 VDD2.n111 0.388379
R349 VDD2.n135 VDD2.n133 0.388379
R350 VDD2.n32 VDD2.n30 0.388379
R351 VDD2.n78 VDD2.n77 0.388379
R352 VDD2.n81 VDD2.n8 0.388379
R353 VDD2.n100 VDD2.n98 0.33524
R354 VDD2.n196 VDD2.n102 0.155672
R355 VDD2.n189 VDD2.n102 0.155672
R356 VDD2.n189 VDD2.n188 0.155672
R357 VDD2.n188 VDD2.n106 0.155672
R358 VDD2.n181 VDD2.n106 0.155672
R359 VDD2.n181 VDD2.n180 0.155672
R360 VDD2.n180 VDD2.n110 0.155672
R361 VDD2.n173 VDD2.n110 0.155672
R362 VDD2.n173 VDD2.n172 0.155672
R363 VDD2.n172 VDD2.n116 0.155672
R364 VDD2.n165 VDD2.n116 0.155672
R365 VDD2.n165 VDD2.n164 0.155672
R366 VDD2.n164 VDD2.n120 0.155672
R367 VDD2.n157 VDD2.n120 0.155672
R368 VDD2.n157 VDD2.n156 0.155672
R369 VDD2.n156 VDD2.n124 0.155672
R370 VDD2.n149 VDD2.n124 0.155672
R371 VDD2.n149 VDD2.n148 0.155672
R372 VDD2.n148 VDD2.n128 0.155672
R373 VDD2.n141 VDD2.n128 0.155672
R374 VDD2.n141 VDD2.n140 0.155672
R375 VDD2.n140 VDD2.n132 0.155672
R376 VDD2.n37 VDD2.n29 0.155672
R377 VDD2.n38 VDD2.n37 0.155672
R378 VDD2.n38 VDD2.n25 0.155672
R379 VDD2.n45 VDD2.n25 0.155672
R380 VDD2.n46 VDD2.n45 0.155672
R381 VDD2.n46 VDD2.n21 0.155672
R382 VDD2.n53 VDD2.n21 0.155672
R383 VDD2.n54 VDD2.n53 0.155672
R384 VDD2.n54 VDD2.n17 0.155672
R385 VDD2.n61 VDD2.n17 0.155672
R386 VDD2.n62 VDD2.n61 0.155672
R387 VDD2.n62 VDD2.n13 0.155672
R388 VDD2.n69 VDD2.n13 0.155672
R389 VDD2.n70 VDD2.n69 0.155672
R390 VDD2.n70 VDD2.n9 0.155672
R391 VDD2.n79 VDD2.n9 0.155672
R392 VDD2.n80 VDD2.n79 0.155672
R393 VDD2.n80 VDD2.n5 0.155672
R394 VDD2.n87 VDD2.n5 0.155672
R395 VDD2.n88 VDD2.n87 0.155672
R396 VDD2.n88 VDD2.n1 0.155672
R397 VDD2.n95 VDD2.n1 0.155672
R398 VTAIL.n400 VTAIL.n308 289.615
R399 VTAIL.n94 VTAIL.n2 289.615
R400 VTAIL.n302 VTAIL.n210 289.615
R401 VTAIL.n200 VTAIL.n108 289.615
R402 VTAIL.n341 VTAIL.n340 185
R403 VTAIL.n343 VTAIL.n342 185
R404 VTAIL.n336 VTAIL.n335 185
R405 VTAIL.n349 VTAIL.n348 185
R406 VTAIL.n351 VTAIL.n350 185
R407 VTAIL.n332 VTAIL.n331 185
R408 VTAIL.n357 VTAIL.n356 185
R409 VTAIL.n359 VTAIL.n358 185
R410 VTAIL.n328 VTAIL.n327 185
R411 VTAIL.n365 VTAIL.n364 185
R412 VTAIL.n367 VTAIL.n366 185
R413 VTAIL.n324 VTAIL.n323 185
R414 VTAIL.n373 VTAIL.n372 185
R415 VTAIL.n375 VTAIL.n374 185
R416 VTAIL.n320 VTAIL.n319 185
R417 VTAIL.n382 VTAIL.n381 185
R418 VTAIL.n383 VTAIL.n318 185
R419 VTAIL.n385 VTAIL.n384 185
R420 VTAIL.n316 VTAIL.n315 185
R421 VTAIL.n391 VTAIL.n390 185
R422 VTAIL.n393 VTAIL.n392 185
R423 VTAIL.n312 VTAIL.n311 185
R424 VTAIL.n399 VTAIL.n398 185
R425 VTAIL.n401 VTAIL.n400 185
R426 VTAIL.n35 VTAIL.n34 185
R427 VTAIL.n37 VTAIL.n36 185
R428 VTAIL.n30 VTAIL.n29 185
R429 VTAIL.n43 VTAIL.n42 185
R430 VTAIL.n45 VTAIL.n44 185
R431 VTAIL.n26 VTAIL.n25 185
R432 VTAIL.n51 VTAIL.n50 185
R433 VTAIL.n53 VTAIL.n52 185
R434 VTAIL.n22 VTAIL.n21 185
R435 VTAIL.n59 VTAIL.n58 185
R436 VTAIL.n61 VTAIL.n60 185
R437 VTAIL.n18 VTAIL.n17 185
R438 VTAIL.n67 VTAIL.n66 185
R439 VTAIL.n69 VTAIL.n68 185
R440 VTAIL.n14 VTAIL.n13 185
R441 VTAIL.n76 VTAIL.n75 185
R442 VTAIL.n77 VTAIL.n12 185
R443 VTAIL.n79 VTAIL.n78 185
R444 VTAIL.n10 VTAIL.n9 185
R445 VTAIL.n85 VTAIL.n84 185
R446 VTAIL.n87 VTAIL.n86 185
R447 VTAIL.n6 VTAIL.n5 185
R448 VTAIL.n93 VTAIL.n92 185
R449 VTAIL.n95 VTAIL.n94 185
R450 VTAIL.n303 VTAIL.n302 185
R451 VTAIL.n301 VTAIL.n300 185
R452 VTAIL.n214 VTAIL.n213 185
R453 VTAIL.n295 VTAIL.n294 185
R454 VTAIL.n293 VTAIL.n292 185
R455 VTAIL.n218 VTAIL.n217 185
R456 VTAIL.n222 VTAIL.n220 185
R457 VTAIL.n287 VTAIL.n286 185
R458 VTAIL.n285 VTAIL.n284 185
R459 VTAIL.n224 VTAIL.n223 185
R460 VTAIL.n279 VTAIL.n278 185
R461 VTAIL.n277 VTAIL.n276 185
R462 VTAIL.n228 VTAIL.n227 185
R463 VTAIL.n271 VTAIL.n270 185
R464 VTAIL.n269 VTAIL.n268 185
R465 VTAIL.n232 VTAIL.n231 185
R466 VTAIL.n263 VTAIL.n262 185
R467 VTAIL.n261 VTAIL.n260 185
R468 VTAIL.n236 VTAIL.n235 185
R469 VTAIL.n255 VTAIL.n254 185
R470 VTAIL.n253 VTAIL.n252 185
R471 VTAIL.n240 VTAIL.n239 185
R472 VTAIL.n247 VTAIL.n246 185
R473 VTAIL.n245 VTAIL.n244 185
R474 VTAIL.n201 VTAIL.n200 185
R475 VTAIL.n199 VTAIL.n198 185
R476 VTAIL.n112 VTAIL.n111 185
R477 VTAIL.n193 VTAIL.n192 185
R478 VTAIL.n191 VTAIL.n190 185
R479 VTAIL.n116 VTAIL.n115 185
R480 VTAIL.n120 VTAIL.n118 185
R481 VTAIL.n185 VTAIL.n184 185
R482 VTAIL.n183 VTAIL.n182 185
R483 VTAIL.n122 VTAIL.n121 185
R484 VTAIL.n177 VTAIL.n176 185
R485 VTAIL.n175 VTAIL.n174 185
R486 VTAIL.n126 VTAIL.n125 185
R487 VTAIL.n169 VTAIL.n168 185
R488 VTAIL.n167 VTAIL.n166 185
R489 VTAIL.n130 VTAIL.n129 185
R490 VTAIL.n161 VTAIL.n160 185
R491 VTAIL.n159 VTAIL.n158 185
R492 VTAIL.n134 VTAIL.n133 185
R493 VTAIL.n153 VTAIL.n152 185
R494 VTAIL.n151 VTAIL.n150 185
R495 VTAIL.n138 VTAIL.n137 185
R496 VTAIL.n145 VTAIL.n144 185
R497 VTAIL.n143 VTAIL.n142 185
R498 VTAIL.n339 VTAIL.t17 147.659
R499 VTAIL.n33 VTAIL.t2 147.659
R500 VTAIL.n243 VTAIL.t8 147.659
R501 VTAIL.n141 VTAIL.t14 147.659
R502 VTAIL.n342 VTAIL.n341 104.615
R503 VTAIL.n342 VTAIL.n335 104.615
R504 VTAIL.n349 VTAIL.n335 104.615
R505 VTAIL.n350 VTAIL.n349 104.615
R506 VTAIL.n350 VTAIL.n331 104.615
R507 VTAIL.n357 VTAIL.n331 104.615
R508 VTAIL.n358 VTAIL.n357 104.615
R509 VTAIL.n358 VTAIL.n327 104.615
R510 VTAIL.n365 VTAIL.n327 104.615
R511 VTAIL.n366 VTAIL.n365 104.615
R512 VTAIL.n366 VTAIL.n323 104.615
R513 VTAIL.n373 VTAIL.n323 104.615
R514 VTAIL.n374 VTAIL.n373 104.615
R515 VTAIL.n374 VTAIL.n319 104.615
R516 VTAIL.n382 VTAIL.n319 104.615
R517 VTAIL.n383 VTAIL.n382 104.615
R518 VTAIL.n384 VTAIL.n383 104.615
R519 VTAIL.n384 VTAIL.n315 104.615
R520 VTAIL.n391 VTAIL.n315 104.615
R521 VTAIL.n392 VTAIL.n391 104.615
R522 VTAIL.n392 VTAIL.n311 104.615
R523 VTAIL.n399 VTAIL.n311 104.615
R524 VTAIL.n400 VTAIL.n399 104.615
R525 VTAIL.n36 VTAIL.n35 104.615
R526 VTAIL.n36 VTAIL.n29 104.615
R527 VTAIL.n43 VTAIL.n29 104.615
R528 VTAIL.n44 VTAIL.n43 104.615
R529 VTAIL.n44 VTAIL.n25 104.615
R530 VTAIL.n51 VTAIL.n25 104.615
R531 VTAIL.n52 VTAIL.n51 104.615
R532 VTAIL.n52 VTAIL.n21 104.615
R533 VTAIL.n59 VTAIL.n21 104.615
R534 VTAIL.n60 VTAIL.n59 104.615
R535 VTAIL.n60 VTAIL.n17 104.615
R536 VTAIL.n67 VTAIL.n17 104.615
R537 VTAIL.n68 VTAIL.n67 104.615
R538 VTAIL.n68 VTAIL.n13 104.615
R539 VTAIL.n76 VTAIL.n13 104.615
R540 VTAIL.n77 VTAIL.n76 104.615
R541 VTAIL.n78 VTAIL.n77 104.615
R542 VTAIL.n78 VTAIL.n9 104.615
R543 VTAIL.n85 VTAIL.n9 104.615
R544 VTAIL.n86 VTAIL.n85 104.615
R545 VTAIL.n86 VTAIL.n5 104.615
R546 VTAIL.n93 VTAIL.n5 104.615
R547 VTAIL.n94 VTAIL.n93 104.615
R548 VTAIL.n302 VTAIL.n301 104.615
R549 VTAIL.n301 VTAIL.n213 104.615
R550 VTAIL.n294 VTAIL.n213 104.615
R551 VTAIL.n294 VTAIL.n293 104.615
R552 VTAIL.n293 VTAIL.n217 104.615
R553 VTAIL.n222 VTAIL.n217 104.615
R554 VTAIL.n286 VTAIL.n222 104.615
R555 VTAIL.n286 VTAIL.n285 104.615
R556 VTAIL.n285 VTAIL.n223 104.615
R557 VTAIL.n278 VTAIL.n223 104.615
R558 VTAIL.n278 VTAIL.n277 104.615
R559 VTAIL.n277 VTAIL.n227 104.615
R560 VTAIL.n270 VTAIL.n227 104.615
R561 VTAIL.n270 VTAIL.n269 104.615
R562 VTAIL.n269 VTAIL.n231 104.615
R563 VTAIL.n262 VTAIL.n231 104.615
R564 VTAIL.n262 VTAIL.n261 104.615
R565 VTAIL.n261 VTAIL.n235 104.615
R566 VTAIL.n254 VTAIL.n235 104.615
R567 VTAIL.n254 VTAIL.n253 104.615
R568 VTAIL.n253 VTAIL.n239 104.615
R569 VTAIL.n246 VTAIL.n239 104.615
R570 VTAIL.n246 VTAIL.n245 104.615
R571 VTAIL.n200 VTAIL.n199 104.615
R572 VTAIL.n199 VTAIL.n111 104.615
R573 VTAIL.n192 VTAIL.n111 104.615
R574 VTAIL.n192 VTAIL.n191 104.615
R575 VTAIL.n191 VTAIL.n115 104.615
R576 VTAIL.n120 VTAIL.n115 104.615
R577 VTAIL.n184 VTAIL.n120 104.615
R578 VTAIL.n184 VTAIL.n183 104.615
R579 VTAIL.n183 VTAIL.n121 104.615
R580 VTAIL.n176 VTAIL.n121 104.615
R581 VTAIL.n176 VTAIL.n175 104.615
R582 VTAIL.n175 VTAIL.n125 104.615
R583 VTAIL.n168 VTAIL.n125 104.615
R584 VTAIL.n168 VTAIL.n167 104.615
R585 VTAIL.n167 VTAIL.n129 104.615
R586 VTAIL.n160 VTAIL.n129 104.615
R587 VTAIL.n160 VTAIL.n159 104.615
R588 VTAIL.n159 VTAIL.n133 104.615
R589 VTAIL.n152 VTAIL.n133 104.615
R590 VTAIL.n152 VTAIL.n151 104.615
R591 VTAIL.n151 VTAIL.n137 104.615
R592 VTAIL.n144 VTAIL.n137 104.615
R593 VTAIL.n144 VTAIL.n143 104.615
R594 VTAIL.n341 VTAIL.t17 52.3082
R595 VTAIL.n35 VTAIL.t2 52.3082
R596 VTAIL.n245 VTAIL.t8 52.3082
R597 VTAIL.n143 VTAIL.t14 52.3082
R598 VTAIL.n209 VTAIL.n208 46.3306
R599 VTAIL.n207 VTAIL.n206 46.3306
R600 VTAIL.n107 VTAIL.n106 46.3306
R601 VTAIL.n105 VTAIL.n104 46.3306
R602 VTAIL.n407 VTAIL.n406 46.3305
R603 VTAIL.n1 VTAIL.n0 46.3305
R604 VTAIL.n101 VTAIL.n100 46.3305
R605 VTAIL.n103 VTAIL.n102 46.3305
R606 VTAIL.n405 VTAIL.n404 34.5126
R607 VTAIL.n99 VTAIL.n98 34.5126
R608 VTAIL.n307 VTAIL.n306 34.5126
R609 VTAIL.n205 VTAIL.n204 34.5126
R610 VTAIL.n105 VTAIL.n103 30.6945
R611 VTAIL.n405 VTAIL.n307 29.1341
R612 VTAIL.n340 VTAIL.n339 15.6677
R613 VTAIL.n34 VTAIL.n33 15.6677
R614 VTAIL.n244 VTAIL.n243 15.6677
R615 VTAIL.n142 VTAIL.n141 15.6677
R616 VTAIL.n385 VTAIL.n316 13.1884
R617 VTAIL.n79 VTAIL.n10 13.1884
R618 VTAIL.n220 VTAIL.n218 13.1884
R619 VTAIL.n118 VTAIL.n116 13.1884
R620 VTAIL.n343 VTAIL.n338 12.8005
R621 VTAIL.n386 VTAIL.n318 12.8005
R622 VTAIL.n390 VTAIL.n389 12.8005
R623 VTAIL.n37 VTAIL.n32 12.8005
R624 VTAIL.n80 VTAIL.n12 12.8005
R625 VTAIL.n84 VTAIL.n83 12.8005
R626 VTAIL.n292 VTAIL.n291 12.8005
R627 VTAIL.n288 VTAIL.n287 12.8005
R628 VTAIL.n247 VTAIL.n242 12.8005
R629 VTAIL.n190 VTAIL.n189 12.8005
R630 VTAIL.n186 VTAIL.n185 12.8005
R631 VTAIL.n145 VTAIL.n140 12.8005
R632 VTAIL.n344 VTAIL.n336 12.0247
R633 VTAIL.n381 VTAIL.n380 12.0247
R634 VTAIL.n393 VTAIL.n314 12.0247
R635 VTAIL.n38 VTAIL.n30 12.0247
R636 VTAIL.n75 VTAIL.n74 12.0247
R637 VTAIL.n87 VTAIL.n8 12.0247
R638 VTAIL.n295 VTAIL.n216 12.0247
R639 VTAIL.n284 VTAIL.n221 12.0247
R640 VTAIL.n248 VTAIL.n240 12.0247
R641 VTAIL.n193 VTAIL.n114 12.0247
R642 VTAIL.n182 VTAIL.n119 12.0247
R643 VTAIL.n146 VTAIL.n138 12.0247
R644 VTAIL.n348 VTAIL.n347 11.249
R645 VTAIL.n379 VTAIL.n320 11.249
R646 VTAIL.n394 VTAIL.n312 11.249
R647 VTAIL.n42 VTAIL.n41 11.249
R648 VTAIL.n73 VTAIL.n14 11.249
R649 VTAIL.n88 VTAIL.n6 11.249
R650 VTAIL.n296 VTAIL.n214 11.249
R651 VTAIL.n283 VTAIL.n224 11.249
R652 VTAIL.n252 VTAIL.n251 11.249
R653 VTAIL.n194 VTAIL.n112 11.249
R654 VTAIL.n181 VTAIL.n122 11.249
R655 VTAIL.n150 VTAIL.n149 11.249
R656 VTAIL.n351 VTAIL.n334 10.4732
R657 VTAIL.n376 VTAIL.n375 10.4732
R658 VTAIL.n398 VTAIL.n397 10.4732
R659 VTAIL.n45 VTAIL.n28 10.4732
R660 VTAIL.n70 VTAIL.n69 10.4732
R661 VTAIL.n92 VTAIL.n91 10.4732
R662 VTAIL.n300 VTAIL.n299 10.4732
R663 VTAIL.n280 VTAIL.n279 10.4732
R664 VTAIL.n255 VTAIL.n238 10.4732
R665 VTAIL.n198 VTAIL.n197 10.4732
R666 VTAIL.n178 VTAIL.n177 10.4732
R667 VTAIL.n153 VTAIL.n136 10.4732
R668 VTAIL.n352 VTAIL.n332 9.69747
R669 VTAIL.n372 VTAIL.n322 9.69747
R670 VTAIL.n401 VTAIL.n310 9.69747
R671 VTAIL.n46 VTAIL.n26 9.69747
R672 VTAIL.n66 VTAIL.n16 9.69747
R673 VTAIL.n95 VTAIL.n4 9.69747
R674 VTAIL.n303 VTAIL.n212 9.69747
R675 VTAIL.n276 VTAIL.n226 9.69747
R676 VTAIL.n256 VTAIL.n236 9.69747
R677 VTAIL.n201 VTAIL.n110 9.69747
R678 VTAIL.n174 VTAIL.n124 9.69747
R679 VTAIL.n154 VTAIL.n134 9.69747
R680 VTAIL.n404 VTAIL.n403 9.45567
R681 VTAIL.n98 VTAIL.n97 9.45567
R682 VTAIL.n306 VTAIL.n305 9.45567
R683 VTAIL.n204 VTAIL.n203 9.45567
R684 VTAIL.n403 VTAIL.n402 9.3005
R685 VTAIL.n310 VTAIL.n309 9.3005
R686 VTAIL.n397 VTAIL.n396 9.3005
R687 VTAIL.n395 VTAIL.n394 9.3005
R688 VTAIL.n314 VTAIL.n313 9.3005
R689 VTAIL.n389 VTAIL.n388 9.3005
R690 VTAIL.n361 VTAIL.n360 9.3005
R691 VTAIL.n330 VTAIL.n329 9.3005
R692 VTAIL.n355 VTAIL.n354 9.3005
R693 VTAIL.n353 VTAIL.n352 9.3005
R694 VTAIL.n334 VTAIL.n333 9.3005
R695 VTAIL.n347 VTAIL.n346 9.3005
R696 VTAIL.n345 VTAIL.n344 9.3005
R697 VTAIL.n338 VTAIL.n337 9.3005
R698 VTAIL.n363 VTAIL.n362 9.3005
R699 VTAIL.n326 VTAIL.n325 9.3005
R700 VTAIL.n369 VTAIL.n368 9.3005
R701 VTAIL.n371 VTAIL.n370 9.3005
R702 VTAIL.n322 VTAIL.n321 9.3005
R703 VTAIL.n377 VTAIL.n376 9.3005
R704 VTAIL.n379 VTAIL.n378 9.3005
R705 VTAIL.n380 VTAIL.n317 9.3005
R706 VTAIL.n387 VTAIL.n386 9.3005
R707 VTAIL.n97 VTAIL.n96 9.3005
R708 VTAIL.n4 VTAIL.n3 9.3005
R709 VTAIL.n91 VTAIL.n90 9.3005
R710 VTAIL.n89 VTAIL.n88 9.3005
R711 VTAIL.n8 VTAIL.n7 9.3005
R712 VTAIL.n83 VTAIL.n82 9.3005
R713 VTAIL.n55 VTAIL.n54 9.3005
R714 VTAIL.n24 VTAIL.n23 9.3005
R715 VTAIL.n49 VTAIL.n48 9.3005
R716 VTAIL.n47 VTAIL.n46 9.3005
R717 VTAIL.n28 VTAIL.n27 9.3005
R718 VTAIL.n41 VTAIL.n40 9.3005
R719 VTAIL.n39 VTAIL.n38 9.3005
R720 VTAIL.n32 VTAIL.n31 9.3005
R721 VTAIL.n57 VTAIL.n56 9.3005
R722 VTAIL.n20 VTAIL.n19 9.3005
R723 VTAIL.n63 VTAIL.n62 9.3005
R724 VTAIL.n65 VTAIL.n64 9.3005
R725 VTAIL.n16 VTAIL.n15 9.3005
R726 VTAIL.n71 VTAIL.n70 9.3005
R727 VTAIL.n73 VTAIL.n72 9.3005
R728 VTAIL.n74 VTAIL.n11 9.3005
R729 VTAIL.n81 VTAIL.n80 9.3005
R730 VTAIL.n230 VTAIL.n229 9.3005
R731 VTAIL.n273 VTAIL.n272 9.3005
R732 VTAIL.n275 VTAIL.n274 9.3005
R733 VTAIL.n226 VTAIL.n225 9.3005
R734 VTAIL.n281 VTAIL.n280 9.3005
R735 VTAIL.n283 VTAIL.n282 9.3005
R736 VTAIL.n221 VTAIL.n219 9.3005
R737 VTAIL.n289 VTAIL.n288 9.3005
R738 VTAIL.n305 VTAIL.n304 9.3005
R739 VTAIL.n212 VTAIL.n211 9.3005
R740 VTAIL.n299 VTAIL.n298 9.3005
R741 VTAIL.n297 VTAIL.n296 9.3005
R742 VTAIL.n216 VTAIL.n215 9.3005
R743 VTAIL.n291 VTAIL.n290 9.3005
R744 VTAIL.n267 VTAIL.n266 9.3005
R745 VTAIL.n265 VTAIL.n264 9.3005
R746 VTAIL.n234 VTAIL.n233 9.3005
R747 VTAIL.n259 VTAIL.n258 9.3005
R748 VTAIL.n257 VTAIL.n256 9.3005
R749 VTAIL.n238 VTAIL.n237 9.3005
R750 VTAIL.n251 VTAIL.n250 9.3005
R751 VTAIL.n249 VTAIL.n248 9.3005
R752 VTAIL.n242 VTAIL.n241 9.3005
R753 VTAIL.n128 VTAIL.n127 9.3005
R754 VTAIL.n171 VTAIL.n170 9.3005
R755 VTAIL.n173 VTAIL.n172 9.3005
R756 VTAIL.n124 VTAIL.n123 9.3005
R757 VTAIL.n179 VTAIL.n178 9.3005
R758 VTAIL.n181 VTAIL.n180 9.3005
R759 VTAIL.n119 VTAIL.n117 9.3005
R760 VTAIL.n187 VTAIL.n186 9.3005
R761 VTAIL.n203 VTAIL.n202 9.3005
R762 VTAIL.n110 VTAIL.n109 9.3005
R763 VTAIL.n197 VTAIL.n196 9.3005
R764 VTAIL.n195 VTAIL.n194 9.3005
R765 VTAIL.n114 VTAIL.n113 9.3005
R766 VTAIL.n189 VTAIL.n188 9.3005
R767 VTAIL.n165 VTAIL.n164 9.3005
R768 VTAIL.n163 VTAIL.n162 9.3005
R769 VTAIL.n132 VTAIL.n131 9.3005
R770 VTAIL.n157 VTAIL.n156 9.3005
R771 VTAIL.n155 VTAIL.n154 9.3005
R772 VTAIL.n136 VTAIL.n135 9.3005
R773 VTAIL.n149 VTAIL.n148 9.3005
R774 VTAIL.n147 VTAIL.n146 9.3005
R775 VTAIL.n140 VTAIL.n139 9.3005
R776 VTAIL.n356 VTAIL.n355 8.92171
R777 VTAIL.n371 VTAIL.n324 8.92171
R778 VTAIL.n402 VTAIL.n308 8.92171
R779 VTAIL.n50 VTAIL.n49 8.92171
R780 VTAIL.n65 VTAIL.n18 8.92171
R781 VTAIL.n96 VTAIL.n2 8.92171
R782 VTAIL.n304 VTAIL.n210 8.92171
R783 VTAIL.n275 VTAIL.n228 8.92171
R784 VTAIL.n260 VTAIL.n259 8.92171
R785 VTAIL.n202 VTAIL.n108 8.92171
R786 VTAIL.n173 VTAIL.n126 8.92171
R787 VTAIL.n158 VTAIL.n157 8.92171
R788 VTAIL.n359 VTAIL.n330 8.14595
R789 VTAIL.n368 VTAIL.n367 8.14595
R790 VTAIL.n53 VTAIL.n24 8.14595
R791 VTAIL.n62 VTAIL.n61 8.14595
R792 VTAIL.n272 VTAIL.n271 8.14595
R793 VTAIL.n263 VTAIL.n234 8.14595
R794 VTAIL.n170 VTAIL.n169 8.14595
R795 VTAIL.n161 VTAIL.n132 8.14595
R796 VTAIL.n360 VTAIL.n328 7.3702
R797 VTAIL.n364 VTAIL.n326 7.3702
R798 VTAIL.n54 VTAIL.n22 7.3702
R799 VTAIL.n58 VTAIL.n20 7.3702
R800 VTAIL.n268 VTAIL.n230 7.3702
R801 VTAIL.n264 VTAIL.n232 7.3702
R802 VTAIL.n166 VTAIL.n128 7.3702
R803 VTAIL.n162 VTAIL.n130 7.3702
R804 VTAIL.n363 VTAIL.n328 6.59444
R805 VTAIL.n364 VTAIL.n363 6.59444
R806 VTAIL.n57 VTAIL.n22 6.59444
R807 VTAIL.n58 VTAIL.n57 6.59444
R808 VTAIL.n268 VTAIL.n267 6.59444
R809 VTAIL.n267 VTAIL.n232 6.59444
R810 VTAIL.n166 VTAIL.n165 6.59444
R811 VTAIL.n165 VTAIL.n130 6.59444
R812 VTAIL.n360 VTAIL.n359 5.81868
R813 VTAIL.n367 VTAIL.n326 5.81868
R814 VTAIL.n54 VTAIL.n53 5.81868
R815 VTAIL.n61 VTAIL.n20 5.81868
R816 VTAIL.n271 VTAIL.n230 5.81868
R817 VTAIL.n264 VTAIL.n263 5.81868
R818 VTAIL.n169 VTAIL.n128 5.81868
R819 VTAIL.n162 VTAIL.n161 5.81868
R820 VTAIL.n356 VTAIL.n330 5.04292
R821 VTAIL.n368 VTAIL.n324 5.04292
R822 VTAIL.n404 VTAIL.n308 5.04292
R823 VTAIL.n50 VTAIL.n24 5.04292
R824 VTAIL.n62 VTAIL.n18 5.04292
R825 VTAIL.n98 VTAIL.n2 5.04292
R826 VTAIL.n306 VTAIL.n210 5.04292
R827 VTAIL.n272 VTAIL.n228 5.04292
R828 VTAIL.n260 VTAIL.n234 5.04292
R829 VTAIL.n204 VTAIL.n108 5.04292
R830 VTAIL.n170 VTAIL.n126 5.04292
R831 VTAIL.n158 VTAIL.n132 5.04292
R832 VTAIL.n339 VTAIL.n337 4.38563
R833 VTAIL.n33 VTAIL.n31 4.38563
R834 VTAIL.n243 VTAIL.n241 4.38563
R835 VTAIL.n141 VTAIL.n139 4.38563
R836 VTAIL.n355 VTAIL.n332 4.26717
R837 VTAIL.n372 VTAIL.n371 4.26717
R838 VTAIL.n402 VTAIL.n401 4.26717
R839 VTAIL.n49 VTAIL.n26 4.26717
R840 VTAIL.n66 VTAIL.n65 4.26717
R841 VTAIL.n96 VTAIL.n95 4.26717
R842 VTAIL.n304 VTAIL.n303 4.26717
R843 VTAIL.n276 VTAIL.n275 4.26717
R844 VTAIL.n259 VTAIL.n236 4.26717
R845 VTAIL.n202 VTAIL.n201 4.26717
R846 VTAIL.n174 VTAIL.n173 4.26717
R847 VTAIL.n157 VTAIL.n134 4.26717
R848 VTAIL.n352 VTAIL.n351 3.49141
R849 VTAIL.n375 VTAIL.n322 3.49141
R850 VTAIL.n398 VTAIL.n310 3.49141
R851 VTAIL.n46 VTAIL.n45 3.49141
R852 VTAIL.n69 VTAIL.n16 3.49141
R853 VTAIL.n92 VTAIL.n4 3.49141
R854 VTAIL.n300 VTAIL.n212 3.49141
R855 VTAIL.n279 VTAIL.n226 3.49141
R856 VTAIL.n256 VTAIL.n255 3.49141
R857 VTAIL.n198 VTAIL.n110 3.49141
R858 VTAIL.n177 VTAIL.n124 3.49141
R859 VTAIL.n154 VTAIL.n153 3.49141
R860 VTAIL.n348 VTAIL.n334 2.71565
R861 VTAIL.n376 VTAIL.n320 2.71565
R862 VTAIL.n397 VTAIL.n312 2.71565
R863 VTAIL.n42 VTAIL.n28 2.71565
R864 VTAIL.n70 VTAIL.n14 2.71565
R865 VTAIL.n91 VTAIL.n6 2.71565
R866 VTAIL.n299 VTAIL.n214 2.71565
R867 VTAIL.n280 VTAIL.n224 2.71565
R868 VTAIL.n252 VTAIL.n238 2.71565
R869 VTAIL.n197 VTAIL.n112 2.71565
R870 VTAIL.n178 VTAIL.n122 2.71565
R871 VTAIL.n150 VTAIL.n136 2.71565
R872 VTAIL.n347 VTAIL.n336 1.93989
R873 VTAIL.n381 VTAIL.n379 1.93989
R874 VTAIL.n394 VTAIL.n393 1.93989
R875 VTAIL.n41 VTAIL.n30 1.93989
R876 VTAIL.n75 VTAIL.n73 1.93989
R877 VTAIL.n88 VTAIL.n87 1.93989
R878 VTAIL.n296 VTAIL.n295 1.93989
R879 VTAIL.n284 VTAIL.n283 1.93989
R880 VTAIL.n251 VTAIL.n240 1.93989
R881 VTAIL.n194 VTAIL.n193 1.93989
R882 VTAIL.n182 VTAIL.n181 1.93989
R883 VTAIL.n149 VTAIL.n138 1.93989
R884 VTAIL.n107 VTAIL.n105 1.56084
R885 VTAIL.n205 VTAIL.n107 1.56084
R886 VTAIL.n209 VTAIL.n207 1.56084
R887 VTAIL.n307 VTAIL.n209 1.56084
R888 VTAIL.n103 VTAIL.n101 1.56084
R889 VTAIL.n101 VTAIL.n99 1.56084
R890 VTAIL.n407 VTAIL.n405 1.56084
R891 VTAIL.n207 VTAIL.n205 1.2505
R892 VTAIL.n99 VTAIL.n1 1.2505
R893 VTAIL VTAIL.n1 1.22895
R894 VTAIL.n344 VTAIL.n343 1.16414
R895 VTAIL.n380 VTAIL.n318 1.16414
R896 VTAIL.n390 VTAIL.n314 1.16414
R897 VTAIL.n38 VTAIL.n37 1.16414
R898 VTAIL.n74 VTAIL.n12 1.16414
R899 VTAIL.n84 VTAIL.n8 1.16414
R900 VTAIL.n292 VTAIL.n216 1.16414
R901 VTAIL.n287 VTAIL.n221 1.16414
R902 VTAIL.n248 VTAIL.n247 1.16414
R903 VTAIL.n190 VTAIL.n114 1.16414
R904 VTAIL.n185 VTAIL.n119 1.16414
R905 VTAIL.n146 VTAIL.n145 1.16414
R906 VTAIL.n406 VTAIL.t16 1.12295
R907 VTAIL.n406 VTAIL.t15 1.12295
R908 VTAIL.n0 VTAIL.t18 1.12295
R909 VTAIL.n0 VTAIL.t11 1.12295
R910 VTAIL.n100 VTAIL.t0 1.12295
R911 VTAIL.n100 VTAIL.t3 1.12295
R912 VTAIL.n102 VTAIL.t5 1.12295
R913 VTAIL.n102 VTAIL.t4 1.12295
R914 VTAIL.n208 VTAIL.t6 1.12295
R915 VTAIL.n208 VTAIL.t9 1.12295
R916 VTAIL.n206 VTAIL.t7 1.12295
R917 VTAIL.n206 VTAIL.t1 1.12295
R918 VTAIL.n106 VTAIL.t13 1.12295
R919 VTAIL.n106 VTAIL.t12 1.12295
R920 VTAIL.n104 VTAIL.t10 1.12295
R921 VTAIL.n104 VTAIL.t19 1.12295
R922 VTAIL.n340 VTAIL.n338 0.388379
R923 VTAIL.n386 VTAIL.n385 0.388379
R924 VTAIL.n389 VTAIL.n316 0.388379
R925 VTAIL.n34 VTAIL.n32 0.388379
R926 VTAIL.n80 VTAIL.n79 0.388379
R927 VTAIL.n83 VTAIL.n10 0.388379
R928 VTAIL.n291 VTAIL.n218 0.388379
R929 VTAIL.n288 VTAIL.n220 0.388379
R930 VTAIL.n244 VTAIL.n242 0.388379
R931 VTAIL.n189 VTAIL.n116 0.388379
R932 VTAIL.n186 VTAIL.n118 0.388379
R933 VTAIL.n142 VTAIL.n140 0.388379
R934 VTAIL VTAIL.n407 0.332397
R935 VTAIL.n345 VTAIL.n337 0.155672
R936 VTAIL.n346 VTAIL.n345 0.155672
R937 VTAIL.n346 VTAIL.n333 0.155672
R938 VTAIL.n353 VTAIL.n333 0.155672
R939 VTAIL.n354 VTAIL.n353 0.155672
R940 VTAIL.n354 VTAIL.n329 0.155672
R941 VTAIL.n361 VTAIL.n329 0.155672
R942 VTAIL.n362 VTAIL.n361 0.155672
R943 VTAIL.n362 VTAIL.n325 0.155672
R944 VTAIL.n369 VTAIL.n325 0.155672
R945 VTAIL.n370 VTAIL.n369 0.155672
R946 VTAIL.n370 VTAIL.n321 0.155672
R947 VTAIL.n377 VTAIL.n321 0.155672
R948 VTAIL.n378 VTAIL.n377 0.155672
R949 VTAIL.n378 VTAIL.n317 0.155672
R950 VTAIL.n387 VTAIL.n317 0.155672
R951 VTAIL.n388 VTAIL.n387 0.155672
R952 VTAIL.n388 VTAIL.n313 0.155672
R953 VTAIL.n395 VTAIL.n313 0.155672
R954 VTAIL.n396 VTAIL.n395 0.155672
R955 VTAIL.n396 VTAIL.n309 0.155672
R956 VTAIL.n403 VTAIL.n309 0.155672
R957 VTAIL.n39 VTAIL.n31 0.155672
R958 VTAIL.n40 VTAIL.n39 0.155672
R959 VTAIL.n40 VTAIL.n27 0.155672
R960 VTAIL.n47 VTAIL.n27 0.155672
R961 VTAIL.n48 VTAIL.n47 0.155672
R962 VTAIL.n48 VTAIL.n23 0.155672
R963 VTAIL.n55 VTAIL.n23 0.155672
R964 VTAIL.n56 VTAIL.n55 0.155672
R965 VTAIL.n56 VTAIL.n19 0.155672
R966 VTAIL.n63 VTAIL.n19 0.155672
R967 VTAIL.n64 VTAIL.n63 0.155672
R968 VTAIL.n64 VTAIL.n15 0.155672
R969 VTAIL.n71 VTAIL.n15 0.155672
R970 VTAIL.n72 VTAIL.n71 0.155672
R971 VTAIL.n72 VTAIL.n11 0.155672
R972 VTAIL.n81 VTAIL.n11 0.155672
R973 VTAIL.n82 VTAIL.n81 0.155672
R974 VTAIL.n82 VTAIL.n7 0.155672
R975 VTAIL.n89 VTAIL.n7 0.155672
R976 VTAIL.n90 VTAIL.n89 0.155672
R977 VTAIL.n90 VTAIL.n3 0.155672
R978 VTAIL.n97 VTAIL.n3 0.155672
R979 VTAIL.n305 VTAIL.n211 0.155672
R980 VTAIL.n298 VTAIL.n211 0.155672
R981 VTAIL.n298 VTAIL.n297 0.155672
R982 VTAIL.n297 VTAIL.n215 0.155672
R983 VTAIL.n290 VTAIL.n215 0.155672
R984 VTAIL.n290 VTAIL.n289 0.155672
R985 VTAIL.n289 VTAIL.n219 0.155672
R986 VTAIL.n282 VTAIL.n219 0.155672
R987 VTAIL.n282 VTAIL.n281 0.155672
R988 VTAIL.n281 VTAIL.n225 0.155672
R989 VTAIL.n274 VTAIL.n225 0.155672
R990 VTAIL.n274 VTAIL.n273 0.155672
R991 VTAIL.n273 VTAIL.n229 0.155672
R992 VTAIL.n266 VTAIL.n229 0.155672
R993 VTAIL.n266 VTAIL.n265 0.155672
R994 VTAIL.n265 VTAIL.n233 0.155672
R995 VTAIL.n258 VTAIL.n233 0.155672
R996 VTAIL.n258 VTAIL.n257 0.155672
R997 VTAIL.n257 VTAIL.n237 0.155672
R998 VTAIL.n250 VTAIL.n237 0.155672
R999 VTAIL.n250 VTAIL.n249 0.155672
R1000 VTAIL.n249 VTAIL.n241 0.155672
R1001 VTAIL.n203 VTAIL.n109 0.155672
R1002 VTAIL.n196 VTAIL.n109 0.155672
R1003 VTAIL.n196 VTAIL.n195 0.155672
R1004 VTAIL.n195 VTAIL.n113 0.155672
R1005 VTAIL.n188 VTAIL.n113 0.155672
R1006 VTAIL.n188 VTAIL.n187 0.155672
R1007 VTAIL.n187 VTAIL.n117 0.155672
R1008 VTAIL.n180 VTAIL.n117 0.155672
R1009 VTAIL.n180 VTAIL.n179 0.155672
R1010 VTAIL.n179 VTAIL.n123 0.155672
R1011 VTAIL.n172 VTAIL.n123 0.155672
R1012 VTAIL.n172 VTAIL.n171 0.155672
R1013 VTAIL.n171 VTAIL.n127 0.155672
R1014 VTAIL.n164 VTAIL.n127 0.155672
R1015 VTAIL.n164 VTAIL.n163 0.155672
R1016 VTAIL.n163 VTAIL.n131 0.155672
R1017 VTAIL.n156 VTAIL.n131 0.155672
R1018 VTAIL.n156 VTAIL.n155 0.155672
R1019 VTAIL.n155 VTAIL.n135 0.155672
R1020 VTAIL.n148 VTAIL.n135 0.155672
R1021 VTAIL.n148 VTAIL.n147 0.155672
R1022 VTAIL.n147 VTAIL.n139 0.155672
R1023 B.n962 B.n961 585
R1024 B.n391 B.n138 585
R1025 B.n390 B.n389 585
R1026 B.n388 B.n387 585
R1027 B.n386 B.n385 585
R1028 B.n384 B.n383 585
R1029 B.n382 B.n381 585
R1030 B.n380 B.n379 585
R1031 B.n378 B.n377 585
R1032 B.n376 B.n375 585
R1033 B.n374 B.n373 585
R1034 B.n372 B.n371 585
R1035 B.n370 B.n369 585
R1036 B.n368 B.n367 585
R1037 B.n366 B.n365 585
R1038 B.n364 B.n363 585
R1039 B.n362 B.n361 585
R1040 B.n360 B.n359 585
R1041 B.n358 B.n357 585
R1042 B.n356 B.n355 585
R1043 B.n354 B.n353 585
R1044 B.n352 B.n351 585
R1045 B.n350 B.n349 585
R1046 B.n348 B.n347 585
R1047 B.n346 B.n345 585
R1048 B.n344 B.n343 585
R1049 B.n342 B.n341 585
R1050 B.n340 B.n339 585
R1051 B.n338 B.n337 585
R1052 B.n336 B.n335 585
R1053 B.n334 B.n333 585
R1054 B.n332 B.n331 585
R1055 B.n330 B.n329 585
R1056 B.n328 B.n327 585
R1057 B.n326 B.n325 585
R1058 B.n324 B.n323 585
R1059 B.n322 B.n321 585
R1060 B.n320 B.n319 585
R1061 B.n318 B.n317 585
R1062 B.n316 B.n315 585
R1063 B.n314 B.n313 585
R1064 B.n312 B.n311 585
R1065 B.n310 B.n309 585
R1066 B.n308 B.n307 585
R1067 B.n306 B.n305 585
R1068 B.n304 B.n303 585
R1069 B.n302 B.n301 585
R1070 B.n300 B.n299 585
R1071 B.n298 B.n297 585
R1072 B.n296 B.n295 585
R1073 B.n294 B.n293 585
R1074 B.n292 B.n291 585
R1075 B.n290 B.n289 585
R1076 B.n288 B.n287 585
R1077 B.n286 B.n285 585
R1078 B.n284 B.n283 585
R1079 B.n282 B.n281 585
R1080 B.n280 B.n279 585
R1081 B.n278 B.n277 585
R1082 B.n276 B.n275 585
R1083 B.n274 B.n273 585
R1084 B.n272 B.n271 585
R1085 B.n270 B.n269 585
R1086 B.n268 B.n267 585
R1087 B.n266 B.n265 585
R1088 B.n264 B.n263 585
R1089 B.n262 B.n261 585
R1090 B.n260 B.n259 585
R1091 B.n258 B.n257 585
R1092 B.n256 B.n255 585
R1093 B.n254 B.n253 585
R1094 B.n252 B.n251 585
R1095 B.n250 B.n249 585
R1096 B.n248 B.n247 585
R1097 B.n246 B.n245 585
R1098 B.n244 B.n243 585
R1099 B.n242 B.n241 585
R1100 B.n240 B.n239 585
R1101 B.n238 B.n237 585
R1102 B.n236 B.n235 585
R1103 B.n234 B.n233 585
R1104 B.n232 B.n231 585
R1105 B.n230 B.n229 585
R1106 B.n228 B.n227 585
R1107 B.n226 B.n225 585
R1108 B.n224 B.n223 585
R1109 B.n222 B.n221 585
R1110 B.n220 B.n219 585
R1111 B.n218 B.n217 585
R1112 B.n216 B.n215 585
R1113 B.n214 B.n213 585
R1114 B.n212 B.n211 585
R1115 B.n210 B.n209 585
R1116 B.n208 B.n207 585
R1117 B.n206 B.n205 585
R1118 B.n204 B.n203 585
R1119 B.n202 B.n201 585
R1120 B.n200 B.n199 585
R1121 B.n198 B.n197 585
R1122 B.n196 B.n195 585
R1123 B.n194 B.n193 585
R1124 B.n192 B.n191 585
R1125 B.n190 B.n189 585
R1126 B.n188 B.n187 585
R1127 B.n186 B.n185 585
R1128 B.n184 B.n183 585
R1129 B.n182 B.n181 585
R1130 B.n180 B.n179 585
R1131 B.n178 B.n177 585
R1132 B.n176 B.n175 585
R1133 B.n174 B.n173 585
R1134 B.n172 B.n171 585
R1135 B.n170 B.n169 585
R1136 B.n168 B.n167 585
R1137 B.n166 B.n165 585
R1138 B.n164 B.n163 585
R1139 B.n162 B.n161 585
R1140 B.n160 B.n159 585
R1141 B.n158 B.n157 585
R1142 B.n156 B.n155 585
R1143 B.n154 B.n153 585
R1144 B.n152 B.n151 585
R1145 B.n150 B.n149 585
R1146 B.n148 B.n147 585
R1147 B.n146 B.n145 585
R1148 B.n74 B.n73 585
R1149 B.n960 B.n75 585
R1150 B.n965 B.n75 585
R1151 B.n959 B.n958 585
R1152 B.n958 B.n71 585
R1153 B.n957 B.n70 585
R1154 B.n971 B.n70 585
R1155 B.n956 B.n69 585
R1156 B.n972 B.n69 585
R1157 B.n955 B.n68 585
R1158 B.n973 B.n68 585
R1159 B.n954 B.n953 585
R1160 B.n953 B.n67 585
R1161 B.n952 B.n63 585
R1162 B.n979 B.n63 585
R1163 B.n951 B.n62 585
R1164 B.n980 B.n62 585
R1165 B.n950 B.n61 585
R1166 B.n981 B.n61 585
R1167 B.n949 B.n948 585
R1168 B.n948 B.n57 585
R1169 B.n947 B.n56 585
R1170 B.n987 B.n56 585
R1171 B.n946 B.n55 585
R1172 B.n988 B.n55 585
R1173 B.n945 B.n54 585
R1174 B.n989 B.n54 585
R1175 B.n944 B.n943 585
R1176 B.n943 B.n50 585
R1177 B.n942 B.n49 585
R1178 B.n995 B.n49 585
R1179 B.n941 B.n48 585
R1180 B.n996 B.n48 585
R1181 B.n940 B.n47 585
R1182 B.n997 B.n47 585
R1183 B.n939 B.n938 585
R1184 B.n938 B.n43 585
R1185 B.n937 B.n42 585
R1186 B.n1003 B.n42 585
R1187 B.n936 B.n41 585
R1188 B.n1004 B.n41 585
R1189 B.n935 B.n40 585
R1190 B.n1005 B.n40 585
R1191 B.n934 B.n933 585
R1192 B.n933 B.n36 585
R1193 B.n932 B.n35 585
R1194 B.n1011 B.n35 585
R1195 B.n931 B.n34 585
R1196 B.n1012 B.n34 585
R1197 B.n930 B.n33 585
R1198 B.n1013 B.n33 585
R1199 B.n929 B.n928 585
R1200 B.n928 B.n32 585
R1201 B.n927 B.n28 585
R1202 B.n1019 B.n28 585
R1203 B.n926 B.n27 585
R1204 B.n1020 B.n27 585
R1205 B.n925 B.n26 585
R1206 B.n1021 B.n26 585
R1207 B.n924 B.n923 585
R1208 B.n923 B.n22 585
R1209 B.n922 B.n21 585
R1210 B.n1027 B.n21 585
R1211 B.n921 B.n20 585
R1212 B.n1028 B.n20 585
R1213 B.n920 B.n19 585
R1214 B.n1029 B.n19 585
R1215 B.n919 B.n918 585
R1216 B.n918 B.n15 585
R1217 B.n917 B.n14 585
R1218 B.n1035 B.n14 585
R1219 B.n916 B.n13 585
R1220 B.n1036 B.n13 585
R1221 B.n915 B.n12 585
R1222 B.n1037 B.n12 585
R1223 B.n914 B.n913 585
R1224 B.n913 B.n8 585
R1225 B.n912 B.n7 585
R1226 B.n1043 B.n7 585
R1227 B.n911 B.n6 585
R1228 B.n1044 B.n6 585
R1229 B.n910 B.n5 585
R1230 B.n1045 B.n5 585
R1231 B.n909 B.n908 585
R1232 B.n908 B.n4 585
R1233 B.n907 B.n392 585
R1234 B.n907 B.n906 585
R1235 B.n897 B.n393 585
R1236 B.n394 B.n393 585
R1237 B.n899 B.n898 585
R1238 B.n900 B.n899 585
R1239 B.n896 B.n398 585
R1240 B.n402 B.n398 585
R1241 B.n895 B.n894 585
R1242 B.n894 B.n893 585
R1243 B.n400 B.n399 585
R1244 B.n401 B.n400 585
R1245 B.n886 B.n885 585
R1246 B.n887 B.n886 585
R1247 B.n884 B.n407 585
R1248 B.n407 B.n406 585
R1249 B.n883 B.n882 585
R1250 B.n882 B.n881 585
R1251 B.n409 B.n408 585
R1252 B.n410 B.n409 585
R1253 B.n874 B.n873 585
R1254 B.n875 B.n874 585
R1255 B.n872 B.n415 585
R1256 B.n415 B.n414 585
R1257 B.n871 B.n870 585
R1258 B.n870 B.n869 585
R1259 B.n417 B.n416 585
R1260 B.n862 B.n417 585
R1261 B.n861 B.n860 585
R1262 B.n863 B.n861 585
R1263 B.n859 B.n422 585
R1264 B.n422 B.n421 585
R1265 B.n858 B.n857 585
R1266 B.n857 B.n856 585
R1267 B.n424 B.n423 585
R1268 B.n425 B.n424 585
R1269 B.n849 B.n848 585
R1270 B.n850 B.n849 585
R1271 B.n847 B.n429 585
R1272 B.n433 B.n429 585
R1273 B.n846 B.n845 585
R1274 B.n845 B.n844 585
R1275 B.n431 B.n430 585
R1276 B.n432 B.n431 585
R1277 B.n837 B.n836 585
R1278 B.n838 B.n837 585
R1279 B.n835 B.n438 585
R1280 B.n438 B.n437 585
R1281 B.n834 B.n833 585
R1282 B.n833 B.n832 585
R1283 B.n440 B.n439 585
R1284 B.n441 B.n440 585
R1285 B.n825 B.n824 585
R1286 B.n826 B.n825 585
R1287 B.n823 B.n446 585
R1288 B.n446 B.n445 585
R1289 B.n822 B.n821 585
R1290 B.n821 B.n820 585
R1291 B.n448 B.n447 585
R1292 B.n449 B.n448 585
R1293 B.n813 B.n812 585
R1294 B.n814 B.n813 585
R1295 B.n811 B.n454 585
R1296 B.n454 B.n453 585
R1297 B.n810 B.n809 585
R1298 B.n809 B.n808 585
R1299 B.n456 B.n455 585
R1300 B.n801 B.n456 585
R1301 B.n800 B.n799 585
R1302 B.n802 B.n800 585
R1303 B.n798 B.n461 585
R1304 B.n461 B.n460 585
R1305 B.n797 B.n796 585
R1306 B.n796 B.n795 585
R1307 B.n463 B.n462 585
R1308 B.n464 B.n463 585
R1309 B.n788 B.n787 585
R1310 B.n789 B.n788 585
R1311 B.n467 B.n466 585
R1312 B.n536 B.n534 585
R1313 B.n537 B.n533 585
R1314 B.n537 B.n468 585
R1315 B.n540 B.n539 585
R1316 B.n541 B.n532 585
R1317 B.n543 B.n542 585
R1318 B.n545 B.n531 585
R1319 B.n548 B.n547 585
R1320 B.n549 B.n530 585
R1321 B.n551 B.n550 585
R1322 B.n553 B.n529 585
R1323 B.n556 B.n555 585
R1324 B.n557 B.n528 585
R1325 B.n559 B.n558 585
R1326 B.n561 B.n527 585
R1327 B.n564 B.n563 585
R1328 B.n565 B.n526 585
R1329 B.n567 B.n566 585
R1330 B.n569 B.n525 585
R1331 B.n572 B.n571 585
R1332 B.n573 B.n524 585
R1333 B.n575 B.n574 585
R1334 B.n577 B.n523 585
R1335 B.n580 B.n579 585
R1336 B.n581 B.n522 585
R1337 B.n583 B.n582 585
R1338 B.n585 B.n521 585
R1339 B.n588 B.n587 585
R1340 B.n589 B.n520 585
R1341 B.n591 B.n590 585
R1342 B.n593 B.n519 585
R1343 B.n596 B.n595 585
R1344 B.n597 B.n518 585
R1345 B.n599 B.n598 585
R1346 B.n601 B.n517 585
R1347 B.n604 B.n603 585
R1348 B.n605 B.n516 585
R1349 B.n607 B.n606 585
R1350 B.n609 B.n515 585
R1351 B.n612 B.n611 585
R1352 B.n613 B.n514 585
R1353 B.n615 B.n614 585
R1354 B.n617 B.n513 585
R1355 B.n620 B.n619 585
R1356 B.n621 B.n512 585
R1357 B.n623 B.n622 585
R1358 B.n625 B.n511 585
R1359 B.n628 B.n627 585
R1360 B.n629 B.n510 585
R1361 B.n631 B.n630 585
R1362 B.n633 B.n509 585
R1363 B.n636 B.n635 585
R1364 B.n637 B.n508 585
R1365 B.n639 B.n638 585
R1366 B.n641 B.n507 585
R1367 B.n644 B.n643 585
R1368 B.n645 B.n506 585
R1369 B.n650 B.n649 585
R1370 B.n652 B.n505 585
R1371 B.n655 B.n654 585
R1372 B.n656 B.n504 585
R1373 B.n658 B.n657 585
R1374 B.n660 B.n503 585
R1375 B.n663 B.n662 585
R1376 B.n664 B.n502 585
R1377 B.n666 B.n665 585
R1378 B.n668 B.n501 585
R1379 B.n671 B.n670 585
R1380 B.n673 B.n498 585
R1381 B.n675 B.n674 585
R1382 B.n677 B.n497 585
R1383 B.n680 B.n679 585
R1384 B.n681 B.n496 585
R1385 B.n683 B.n682 585
R1386 B.n685 B.n495 585
R1387 B.n688 B.n687 585
R1388 B.n689 B.n494 585
R1389 B.n691 B.n690 585
R1390 B.n693 B.n493 585
R1391 B.n696 B.n695 585
R1392 B.n697 B.n492 585
R1393 B.n699 B.n698 585
R1394 B.n701 B.n491 585
R1395 B.n704 B.n703 585
R1396 B.n705 B.n490 585
R1397 B.n707 B.n706 585
R1398 B.n709 B.n489 585
R1399 B.n712 B.n711 585
R1400 B.n713 B.n488 585
R1401 B.n715 B.n714 585
R1402 B.n717 B.n487 585
R1403 B.n720 B.n719 585
R1404 B.n721 B.n486 585
R1405 B.n723 B.n722 585
R1406 B.n725 B.n485 585
R1407 B.n728 B.n727 585
R1408 B.n729 B.n484 585
R1409 B.n731 B.n730 585
R1410 B.n733 B.n483 585
R1411 B.n736 B.n735 585
R1412 B.n737 B.n482 585
R1413 B.n739 B.n738 585
R1414 B.n741 B.n481 585
R1415 B.n744 B.n743 585
R1416 B.n745 B.n480 585
R1417 B.n747 B.n746 585
R1418 B.n749 B.n479 585
R1419 B.n752 B.n751 585
R1420 B.n753 B.n478 585
R1421 B.n755 B.n754 585
R1422 B.n757 B.n477 585
R1423 B.n760 B.n759 585
R1424 B.n761 B.n476 585
R1425 B.n763 B.n762 585
R1426 B.n765 B.n475 585
R1427 B.n768 B.n767 585
R1428 B.n769 B.n474 585
R1429 B.n771 B.n770 585
R1430 B.n773 B.n473 585
R1431 B.n776 B.n775 585
R1432 B.n777 B.n472 585
R1433 B.n779 B.n778 585
R1434 B.n781 B.n471 585
R1435 B.n782 B.n470 585
R1436 B.n785 B.n784 585
R1437 B.n786 B.n469 585
R1438 B.n469 B.n468 585
R1439 B.n791 B.n790 585
R1440 B.n790 B.n789 585
R1441 B.n792 B.n465 585
R1442 B.n465 B.n464 585
R1443 B.n794 B.n793 585
R1444 B.n795 B.n794 585
R1445 B.n459 B.n458 585
R1446 B.n460 B.n459 585
R1447 B.n804 B.n803 585
R1448 B.n803 B.n802 585
R1449 B.n805 B.n457 585
R1450 B.n801 B.n457 585
R1451 B.n807 B.n806 585
R1452 B.n808 B.n807 585
R1453 B.n452 B.n451 585
R1454 B.n453 B.n452 585
R1455 B.n816 B.n815 585
R1456 B.n815 B.n814 585
R1457 B.n817 B.n450 585
R1458 B.n450 B.n449 585
R1459 B.n819 B.n818 585
R1460 B.n820 B.n819 585
R1461 B.n444 B.n443 585
R1462 B.n445 B.n444 585
R1463 B.n828 B.n827 585
R1464 B.n827 B.n826 585
R1465 B.n829 B.n442 585
R1466 B.n442 B.n441 585
R1467 B.n831 B.n830 585
R1468 B.n832 B.n831 585
R1469 B.n436 B.n435 585
R1470 B.n437 B.n436 585
R1471 B.n840 B.n839 585
R1472 B.n839 B.n838 585
R1473 B.n841 B.n434 585
R1474 B.n434 B.n432 585
R1475 B.n843 B.n842 585
R1476 B.n844 B.n843 585
R1477 B.n428 B.n427 585
R1478 B.n433 B.n428 585
R1479 B.n852 B.n851 585
R1480 B.n851 B.n850 585
R1481 B.n853 B.n426 585
R1482 B.n426 B.n425 585
R1483 B.n855 B.n854 585
R1484 B.n856 B.n855 585
R1485 B.n420 B.n419 585
R1486 B.n421 B.n420 585
R1487 B.n865 B.n864 585
R1488 B.n864 B.n863 585
R1489 B.n866 B.n418 585
R1490 B.n862 B.n418 585
R1491 B.n868 B.n867 585
R1492 B.n869 B.n868 585
R1493 B.n413 B.n412 585
R1494 B.n414 B.n413 585
R1495 B.n877 B.n876 585
R1496 B.n876 B.n875 585
R1497 B.n878 B.n411 585
R1498 B.n411 B.n410 585
R1499 B.n880 B.n879 585
R1500 B.n881 B.n880 585
R1501 B.n405 B.n404 585
R1502 B.n406 B.n405 585
R1503 B.n889 B.n888 585
R1504 B.n888 B.n887 585
R1505 B.n890 B.n403 585
R1506 B.n403 B.n401 585
R1507 B.n892 B.n891 585
R1508 B.n893 B.n892 585
R1509 B.n397 B.n396 585
R1510 B.n402 B.n397 585
R1511 B.n902 B.n901 585
R1512 B.n901 B.n900 585
R1513 B.n903 B.n395 585
R1514 B.n395 B.n394 585
R1515 B.n905 B.n904 585
R1516 B.n906 B.n905 585
R1517 B.n2 B.n0 585
R1518 B.n4 B.n2 585
R1519 B.n3 B.n1 585
R1520 B.n1044 B.n3 585
R1521 B.n1042 B.n1041 585
R1522 B.n1043 B.n1042 585
R1523 B.n1040 B.n9 585
R1524 B.n9 B.n8 585
R1525 B.n1039 B.n1038 585
R1526 B.n1038 B.n1037 585
R1527 B.n11 B.n10 585
R1528 B.n1036 B.n11 585
R1529 B.n1034 B.n1033 585
R1530 B.n1035 B.n1034 585
R1531 B.n1032 B.n16 585
R1532 B.n16 B.n15 585
R1533 B.n1031 B.n1030 585
R1534 B.n1030 B.n1029 585
R1535 B.n18 B.n17 585
R1536 B.n1028 B.n18 585
R1537 B.n1026 B.n1025 585
R1538 B.n1027 B.n1026 585
R1539 B.n1024 B.n23 585
R1540 B.n23 B.n22 585
R1541 B.n1023 B.n1022 585
R1542 B.n1022 B.n1021 585
R1543 B.n25 B.n24 585
R1544 B.n1020 B.n25 585
R1545 B.n1018 B.n1017 585
R1546 B.n1019 B.n1018 585
R1547 B.n1016 B.n29 585
R1548 B.n32 B.n29 585
R1549 B.n1015 B.n1014 585
R1550 B.n1014 B.n1013 585
R1551 B.n31 B.n30 585
R1552 B.n1012 B.n31 585
R1553 B.n1010 B.n1009 585
R1554 B.n1011 B.n1010 585
R1555 B.n1008 B.n37 585
R1556 B.n37 B.n36 585
R1557 B.n1007 B.n1006 585
R1558 B.n1006 B.n1005 585
R1559 B.n39 B.n38 585
R1560 B.n1004 B.n39 585
R1561 B.n1002 B.n1001 585
R1562 B.n1003 B.n1002 585
R1563 B.n1000 B.n44 585
R1564 B.n44 B.n43 585
R1565 B.n999 B.n998 585
R1566 B.n998 B.n997 585
R1567 B.n46 B.n45 585
R1568 B.n996 B.n46 585
R1569 B.n994 B.n993 585
R1570 B.n995 B.n994 585
R1571 B.n992 B.n51 585
R1572 B.n51 B.n50 585
R1573 B.n991 B.n990 585
R1574 B.n990 B.n989 585
R1575 B.n53 B.n52 585
R1576 B.n988 B.n53 585
R1577 B.n986 B.n985 585
R1578 B.n987 B.n986 585
R1579 B.n984 B.n58 585
R1580 B.n58 B.n57 585
R1581 B.n983 B.n982 585
R1582 B.n982 B.n981 585
R1583 B.n60 B.n59 585
R1584 B.n980 B.n60 585
R1585 B.n978 B.n977 585
R1586 B.n979 B.n978 585
R1587 B.n976 B.n64 585
R1588 B.n67 B.n64 585
R1589 B.n975 B.n974 585
R1590 B.n974 B.n973 585
R1591 B.n66 B.n65 585
R1592 B.n972 B.n66 585
R1593 B.n970 B.n969 585
R1594 B.n971 B.n970 585
R1595 B.n968 B.n72 585
R1596 B.n72 B.n71 585
R1597 B.n967 B.n966 585
R1598 B.n966 B.n965 585
R1599 B.n1047 B.n1046 585
R1600 B.n1046 B.n1045 585
R1601 B.n790 B.n467 506.916
R1602 B.n966 B.n74 506.916
R1603 B.n788 B.n469 506.916
R1604 B.n962 B.n75 506.916
R1605 B.n499 B.t14 492.611
R1606 B.n646 B.t18 492.611
R1607 B.n142 B.t10 492.611
R1608 B.n139 B.t21 492.611
R1609 B.n499 B.t17 414.69
R1610 B.n139 B.t22 414.69
R1611 B.n646 B.t20 414.69
R1612 B.n142 B.t12 414.69
R1613 B.n500 B.t16 379.587
R1614 B.n140 B.t23 379.587
R1615 B.n647 B.t19 379.587
R1616 B.n143 B.t13 379.587
R1617 B.n964 B.n963 256.663
R1618 B.n964 B.n137 256.663
R1619 B.n964 B.n136 256.663
R1620 B.n964 B.n135 256.663
R1621 B.n964 B.n134 256.663
R1622 B.n964 B.n133 256.663
R1623 B.n964 B.n132 256.663
R1624 B.n964 B.n131 256.663
R1625 B.n964 B.n130 256.663
R1626 B.n964 B.n129 256.663
R1627 B.n964 B.n128 256.663
R1628 B.n964 B.n127 256.663
R1629 B.n964 B.n126 256.663
R1630 B.n964 B.n125 256.663
R1631 B.n964 B.n124 256.663
R1632 B.n964 B.n123 256.663
R1633 B.n964 B.n122 256.663
R1634 B.n964 B.n121 256.663
R1635 B.n964 B.n120 256.663
R1636 B.n964 B.n119 256.663
R1637 B.n964 B.n118 256.663
R1638 B.n964 B.n117 256.663
R1639 B.n964 B.n116 256.663
R1640 B.n964 B.n115 256.663
R1641 B.n964 B.n114 256.663
R1642 B.n964 B.n113 256.663
R1643 B.n964 B.n112 256.663
R1644 B.n964 B.n111 256.663
R1645 B.n964 B.n110 256.663
R1646 B.n964 B.n109 256.663
R1647 B.n964 B.n108 256.663
R1648 B.n964 B.n107 256.663
R1649 B.n964 B.n106 256.663
R1650 B.n964 B.n105 256.663
R1651 B.n964 B.n104 256.663
R1652 B.n964 B.n103 256.663
R1653 B.n964 B.n102 256.663
R1654 B.n964 B.n101 256.663
R1655 B.n964 B.n100 256.663
R1656 B.n964 B.n99 256.663
R1657 B.n964 B.n98 256.663
R1658 B.n964 B.n97 256.663
R1659 B.n964 B.n96 256.663
R1660 B.n964 B.n95 256.663
R1661 B.n964 B.n94 256.663
R1662 B.n964 B.n93 256.663
R1663 B.n964 B.n92 256.663
R1664 B.n964 B.n91 256.663
R1665 B.n964 B.n90 256.663
R1666 B.n964 B.n89 256.663
R1667 B.n964 B.n88 256.663
R1668 B.n964 B.n87 256.663
R1669 B.n964 B.n86 256.663
R1670 B.n964 B.n85 256.663
R1671 B.n964 B.n84 256.663
R1672 B.n964 B.n83 256.663
R1673 B.n964 B.n82 256.663
R1674 B.n964 B.n81 256.663
R1675 B.n964 B.n80 256.663
R1676 B.n964 B.n79 256.663
R1677 B.n964 B.n78 256.663
R1678 B.n964 B.n77 256.663
R1679 B.n964 B.n76 256.663
R1680 B.n535 B.n468 256.663
R1681 B.n538 B.n468 256.663
R1682 B.n544 B.n468 256.663
R1683 B.n546 B.n468 256.663
R1684 B.n552 B.n468 256.663
R1685 B.n554 B.n468 256.663
R1686 B.n560 B.n468 256.663
R1687 B.n562 B.n468 256.663
R1688 B.n568 B.n468 256.663
R1689 B.n570 B.n468 256.663
R1690 B.n576 B.n468 256.663
R1691 B.n578 B.n468 256.663
R1692 B.n584 B.n468 256.663
R1693 B.n586 B.n468 256.663
R1694 B.n592 B.n468 256.663
R1695 B.n594 B.n468 256.663
R1696 B.n600 B.n468 256.663
R1697 B.n602 B.n468 256.663
R1698 B.n608 B.n468 256.663
R1699 B.n610 B.n468 256.663
R1700 B.n616 B.n468 256.663
R1701 B.n618 B.n468 256.663
R1702 B.n624 B.n468 256.663
R1703 B.n626 B.n468 256.663
R1704 B.n632 B.n468 256.663
R1705 B.n634 B.n468 256.663
R1706 B.n640 B.n468 256.663
R1707 B.n642 B.n468 256.663
R1708 B.n651 B.n468 256.663
R1709 B.n653 B.n468 256.663
R1710 B.n659 B.n468 256.663
R1711 B.n661 B.n468 256.663
R1712 B.n667 B.n468 256.663
R1713 B.n669 B.n468 256.663
R1714 B.n676 B.n468 256.663
R1715 B.n678 B.n468 256.663
R1716 B.n684 B.n468 256.663
R1717 B.n686 B.n468 256.663
R1718 B.n692 B.n468 256.663
R1719 B.n694 B.n468 256.663
R1720 B.n700 B.n468 256.663
R1721 B.n702 B.n468 256.663
R1722 B.n708 B.n468 256.663
R1723 B.n710 B.n468 256.663
R1724 B.n716 B.n468 256.663
R1725 B.n718 B.n468 256.663
R1726 B.n724 B.n468 256.663
R1727 B.n726 B.n468 256.663
R1728 B.n732 B.n468 256.663
R1729 B.n734 B.n468 256.663
R1730 B.n740 B.n468 256.663
R1731 B.n742 B.n468 256.663
R1732 B.n748 B.n468 256.663
R1733 B.n750 B.n468 256.663
R1734 B.n756 B.n468 256.663
R1735 B.n758 B.n468 256.663
R1736 B.n764 B.n468 256.663
R1737 B.n766 B.n468 256.663
R1738 B.n772 B.n468 256.663
R1739 B.n774 B.n468 256.663
R1740 B.n780 B.n468 256.663
R1741 B.n783 B.n468 256.663
R1742 B.n790 B.n465 163.367
R1743 B.n794 B.n465 163.367
R1744 B.n794 B.n459 163.367
R1745 B.n803 B.n459 163.367
R1746 B.n803 B.n457 163.367
R1747 B.n807 B.n457 163.367
R1748 B.n807 B.n452 163.367
R1749 B.n815 B.n452 163.367
R1750 B.n815 B.n450 163.367
R1751 B.n819 B.n450 163.367
R1752 B.n819 B.n444 163.367
R1753 B.n827 B.n444 163.367
R1754 B.n827 B.n442 163.367
R1755 B.n831 B.n442 163.367
R1756 B.n831 B.n436 163.367
R1757 B.n839 B.n436 163.367
R1758 B.n839 B.n434 163.367
R1759 B.n843 B.n434 163.367
R1760 B.n843 B.n428 163.367
R1761 B.n851 B.n428 163.367
R1762 B.n851 B.n426 163.367
R1763 B.n855 B.n426 163.367
R1764 B.n855 B.n420 163.367
R1765 B.n864 B.n420 163.367
R1766 B.n864 B.n418 163.367
R1767 B.n868 B.n418 163.367
R1768 B.n868 B.n413 163.367
R1769 B.n876 B.n413 163.367
R1770 B.n876 B.n411 163.367
R1771 B.n880 B.n411 163.367
R1772 B.n880 B.n405 163.367
R1773 B.n888 B.n405 163.367
R1774 B.n888 B.n403 163.367
R1775 B.n892 B.n403 163.367
R1776 B.n892 B.n397 163.367
R1777 B.n901 B.n397 163.367
R1778 B.n901 B.n395 163.367
R1779 B.n905 B.n395 163.367
R1780 B.n905 B.n2 163.367
R1781 B.n1046 B.n2 163.367
R1782 B.n1046 B.n3 163.367
R1783 B.n1042 B.n3 163.367
R1784 B.n1042 B.n9 163.367
R1785 B.n1038 B.n9 163.367
R1786 B.n1038 B.n11 163.367
R1787 B.n1034 B.n11 163.367
R1788 B.n1034 B.n16 163.367
R1789 B.n1030 B.n16 163.367
R1790 B.n1030 B.n18 163.367
R1791 B.n1026 B.n18 163.367
R1792 B.n1026 B.n23 163.367
R1793 B.n1022 B.n23 163.367
R1794 B.n1022 B.n25 163.367
R1795 B.n1018 B.n25 163.367
R1796 B.n1018 B.n29 163.367
R1797 B.n1014 B.n29 163.367
R1798 B.n1014 B.n31 163.367
R1799 B.n1010 B.n31 163.367
R1800 B.n1010 B.n37 163.367
R1801 B.n1006 B.n37 163.367
R1802 B.n1006 B.n39 163.367
R1803 B.n1002 B.n39 163.367
R1804 B.n1002 B.n44 163.367
R1805 B.n998 B.n44 163.367
R1806 B.n998 B.n46 163.367
R1807 B.n994 B.n46 163.367
R1808 B.n994 B.n51 163.367
R1809 B.n990 B.n51 163.367
R1810 B.n990 B.n53 163.367
R1811 B.n986 B.n53 163.367
R1812 B.n986 B.n58 163.367
R1813 B.n982 B.n58 163.367
R1814 B.n982 B.n60 163.367
R1815 B.n978 B.n60 163.367
R1816 B.n978 B.n64 163.367
R1817 B.n974 B.n64 163.367
R1818 B.n974 B.n66 163.367
R1819 B.n970 B.n66 163.367
R1820 B.n970 B.n72 163.367
R1821 B.n966 B.n72 163.367
R1822 B.n537 B.n536 163.367
R1823 B.n539 B.n537 163.367
R1824 B.n543 B.n532 163.367
R1825 B.n547 B.n545 163.367
R1826 B.n551 B.n530 163.367
R1827 B.n555 B.n553 163.367
R1828 B.n559 B.n528 163.367
R1829 B.n563 B.n561 163.367
R1830 B.n567 B.n526 163.367
R1831 B.n571 B.n569 163.367
R1832 B.n575 B.n524 163.367
R1833 B.n579 B.n577 163.367
R1834 B.n583 B.n522 163.367
R1835 B.n587 B.n585 163.367
R1836 B.n591 B.n520 163.367
R1837 B.n595 B.n593 163.367
R1838 B.n599 B.n518 163.367
R1839 B.n603 B.n601 163.367
R1840 B.n607 B.n516 163.367
R1841 B.n611 B.n609 163.367
R1842 B.n615 B.n514 163.367
R1843 B.n619 B.n617 163.367
R1844 B.n623 B.n512 163.367
R1845 B.n627 B.n625 163.367
R1846 B.n631 B.n510 163.367
R1847 B.n635 B.n633 163.367
R1848 B.n639 B.n508 163.367
R1849 B.n643 B.n641 163.367
R1850 B.n650 B.n506 163.367
R1851 B.n654 B.n652 163.367
R1852 B.n658 B.n504 163.367
R1853 B.n662 B.n660 163.367
R1854 B.n666 B.n502 163.367
R1855 B.n670 B.n668 163.367
R1856 B.n675 B.n498 163.367
R1857 B.n679 B.n677 163.367
R1858 B.n683 B.n496 163.367
R1859 B.n687 B.n685 163.367
R1860 B.n691 B.n494 163.367
R1861 B.n695 B.n693 163.367
R1862 B.n699 B.n492 163.367
R1863 B.n703 B.n701 163.367
R1864 B.n707 B.n490 163.367
R1865 B.n711 B.n709 163.367
R1866 B.n715 B.n488 163.367
R1867 B.n719 B.n717 163.367
R1868 B.n723 B.n486 163.367
R1869 B.n727 B.n725 163.367
R1870 B.n731 B.n484 163.367
R1871 B.n735 B.n733 163.367
R1872 B.n739 B.n482 163.367
R1873 B.n743 B.n741 163.367
R1874 B.n747 B.n480 163.367
R1875 B.n751 B.n749 163.367
R1876 B.n755 B.n478 163.367
R1877 B.n759 B.n757 163.367
R1878 B.n763 B.n476 163.367
R1879 B.n767 B.n765 163.367
R1880 B.n771 B.n474 163.367
R1881 B.n775 B.n773 163.367
R1882 B.n779 B.n472 163.367
R1883 B.n782 B.n781 163.367
R1884 B.n784 B.n469 163.367
R1885 B.n788 B.n463 163.367
R1886 B.n796 B.n463 163.367
R1887 B.n796 B.n461 163.367
R1888 B.n800 B.n461 163.367
R1889 B.n800 B.n456 163.367
R1890 B.n809 B.n456 163.367
R1891 B.n809 B.n454 163.367
R1892 B.n813 B.n454 163.367
R1893 B.n813 B.n448 163.367
R1894 B.n821 B.n448 163.367
R1895 B.n821 B.n446 163.367
R1896 B.n825 B.n446 163.367
R1897 B.n825 B.n440 163.367
R1898 B.n833 B.n440 163.367
R1899 B.n833 B.n438 163.367
R1900 B.n837 B.n438 163.367
R1901 B.n837 B.n431 163.367
R1902 B.n845 B.n431 163.367
R1903 B.n845 B.n429 163.367
R1904 B.n849 B.n429 163.367
R1905 B.n849 B.n424 163.367
R1906 B.n857 B.n424 163.367
R1907 B.n857 B.n422 163.367
R1908 B.n861 B.n422 163.367
R1909 B.n861 B.n417 163.367
R1910 B.n870 B.n417 163.367
R1911 B.n870 B.n415 163.367
R1912 B.n874 B.n415 163.367
R1913 B.n874 B.n409 163.367
R1914 B.n882 B.n409 163.367
R1915 B.n882 B.n407 163.367
R1916 B.n886 B.n407 163.367
R1917 B.n886 B.n400 163.367
R1918 B.n894 B.n400 163.367
R1919 B.n894 B.n398 163.367
R1920 B.n899 B.n398 163.367
R1921 B.n899 B.n393 163.367
R1922 B.n907 B.n393 163.367
R1923 B.n908 B.n907 163.367
R1924 B.n908 B.n5 163.367
R1925 B.n6 B.n5 163.367
R1926 B.n7 B.n6 163.367
R1927 B.n913 B.n7 163.367
R1928 B.n913 B.n12 163.367
R1929 B.n13 B.n12 163.367
R1930 B.n14 B.n13 163.367
R1931 B.n918 B.n14 163.367
R1932 B.n918 B.n19 163.367
R1933 B.n20 B.n19 163.367
R1934 B.n21 B.n20 163.367
R1935 B.n923 B.n21 163.367
R1936 B.n923 B.n26 163.367
R1937 B.n27 B.n26 163.367
R1938 B.n28 B.n27 163.367
R1939 B.n928 B.n28 163.367
R1940 B.n928 B.n33 163.367
R1941 B.n34 B.n33 163.367
R1942 B.n35 B.n34 163.367
R1943 B.n933 B.n35 163.367
R1944 B.n933 B.n40 163.367
R1945 B.n41 B.n40 163.367
R1946 B.n42 B.n41 163.367
R1947 B.n938 B.n42 163.367
R1948 B.n938 B.n47 163.367
R1949 B.n48 B.n47 163.367
R1950 B.n49 B.n48 163.367
R1951 B.n943 B.n49 163.367
R1952 B.n943 B.n54 163.367
R1953 B.n55 B.n54 163.367
R1954 B.n56 B.n55 163.367
R1955 B.n948 B.n56 163.367
R1956 B.n948 B.n61 163.367
R1957 B.n62 B.n61 163.367
R1958 B.n63 B.n62 163.367
R1959 B.n953 B.n63 163.367
R1960 B.n953 B.n68 163.367
R1961 B.n69 B.n68 163.367
R1962 B.n70 B.n69 163.367
R1963 B.n958 B.n70 163.367
R1964 B.n958 B.n75 163.367
R1965 B.n147 B.n146 163.367
R1966 B.n151 B.n150 163.367
R1967 B.n155 B.n154 163.367
R1968 B.n159 B.n158 163.367
R1969 B.n163 B.n162 163.367
R1970 B.n167 B.n166 163.367
R1971 B.n171 B.n170 163.367
R1972 B.n175 B.n174 163.367
R1973 B.n179 B.n178 163.367
R1974 B.n183 B.n182 163.367
R1975 B.n187 B.n186 163.367
R1976 B.n191 B.n190 163.367
R1977 B.n195 B.n194 163.367
R1978 B.n199 B.n198 163.367
R1979 B.n203 B.n202 163.367
R1980 B.n207 B.n206 163.367
R1981 B.n211 B.n210 163.367
R1982 B.n215 B.n214 163.367
R1983 B.n219 B.n218 163.367
R1984 B.n223 B.n222 163.367
R1985 B.n227 B.n226 163.367
R1986 B.n231 B.n230 163.367
R1987 B.n235 B.n234 163.367
R1988 B.n239 B.n238 163.367
R1989 B.n243 B.n242 163.367
R1990 B.n247 B.n246 163.367
R1991 B.n251 B.n250 163.367
R1992 B.n255 B.n254 163.367
R1993 B.n259 B.n258 163.367
R1994 B.n263 B.n262 163.367
R1995 B.n267 B.n266 163.367
R1996 B.n271 B.n270 163.367
R1997 B.n275 B.n274 163.367
R1998 B.n279 B.n278 163.367
R1999 B.n283 B.n282 163.367
R2000 B.n287 B.n286 163.367
R2001 B.n291 B.n290 163.367
R2002 B.n295 B.n294 163.367
R2003 B.n299 B.n298 163.367
R2004 B.n303 B.n302 163.367
R2005 B.n307 B.n306 163.367
R2006 B.n311 B.n310 163.367
R2007 B.n315 B.n314 163.367
R2008 B.n319 B.n318 163.367
R2009 B.n323 B.n322 163.367
R2010 B.n327 B.n326 163.367
R2011 B.n331 B.n330 163.367
R2012 B.n335 B.n334 163.367
R2013 B.n339 B.n338 163.367
R2014 B.n343 B.n342 163.367
R2015 B.n347 B.n346 163.367
R2016 B.n351 B.n350 163.367
R2017 B.n355 B.n354 163.367
R2018 B.n359 B.n358 163.367
R2019 B.n363 B.n362 163.367
R2020 B.n367 B.n366 163.367
R2021 B.n371 B.n370 163.367
R2022 B.n375 B.n374 163.367
R2023 B.n379 B.n378 163.367
R2024 B.n383 B.n382 163.367
R2025 B.n387 B.n386 163.367
R2026 B.n389 B.n138 163.367
R2027 B.n535 B.n467 71.676
R2028 B.n539 B.n538 71.676
R2029 B.n544 B.n543 71.676
R2030 B.n547 B.n546 71.676
R2031 B.n552 B.n551 71.676
R2032 B.n555 B.n554 71.676
R2033 B.n560 B.n559 71.676
R2034 B.n563 B.n562 71.676
R2035 B.n568 B.n567 71.676
R2036 B.n571 B.n570 71.676
R2037 B.n576 B.n575 71.676
R2038 B.n579 B.n578 71.676
R2039 B.n584 B.n583 71.676
R2040 B.n587 B.n586 71.676
R2041 B.n592 B.n591 71.676
R2042 B.n595 B.n594 71.676
R2043 B.n600 B.n599 71.676
R2044 B.n603 B.n602 71.676
R2045 B.n608 B.n607 71.676
R2046 B.n611 B.n610 71.676
R2047 B.n616 B.n615 71.676
R2048 B.n619 B.n618 71.676
R2049 B.n624 B.n623 71.676
R2050 B.n627 B.n626 71.676
R2051 B.n632 B.n631 71.676
R2052 B.n635 B.n634 71.676
R2053 B.n640 B.n639 71.676
R2054 B.n643 B.n642 71.676
R2055 B.n651 B.n650 71.676
R2056 B.n654 B.n653 71.676
R2057 B.n659 B.n658 71.676
R2058 B.n662 B.n661 71.676
R2059 B.n667 B.n666 71.676
R2060 B.n670 B.n669 71.676
R2061 B.n676 B.n675 71.676
R2062 B.n679 B.n678 71.676
R2063 B.n684 B.n683 71.676
R2064 B.n687 B.n686 71.676
R2065 B.n692 B.n691 71.676
R2066 B.n695 B.n694 71.676
R2067 B.n700 B.n699 71.676
R2068 B.n703 B.n702 71.676
R2069 B.n708 B.n707 71.676
R2070 B.n711 B.n710 71.676
R2071 B.n716 B.n715 71.676
R2072 B.n719 B.n718 71.676
R2073 B.n724 B.n723 71.676
R2074 B.n727 B.n726 71.676
R2075 B.n732 B.n731 71.676
R2076 B.n735 B.n734 71.676
R2077 B.n740 B.n739 71.676
R2078 B.n743 B.n742 71.676
R2079 B.n748 B.n747 71.676
R2080 B.n751 B.n750 71.676
R2081 B.n756 B.n755 71.676
R2082 B.n759 B.n758 71.676
R2083 B.n764 B.n763 71.676
R2084 B.n767 B.n766 71.676
R2085 B.n772 B.n771 71.676
R2086 B.n775 B.n774 71.676
R2087 B.n780 B.n779 71.676
R2088 B.n783 B.n782 71.676
R2089 B.n76 B.n74 71.676
R2090 B.n147 B.n77 71.676
R2091 B.n151 B.n78 71.676
R2092 B.n155 B.n79 71.676
R2093 B.n159 B.n80 71.676
R2094 B.n163 B.n81 71.676
R2095 B.n167 B.n82 71.676
R2096 B.n171 B.n83 71.676
R2097 B.n175 B.n84 71.676
R2098 B.n179 B.n85 71.676
R2099 B.n183 B.n86 71.676
R2100 B.n187 B.n87 71.676
R2101 B.n191 B.n88 71.676
R2102 B.n195 B.n89 71.676
R2103 B.n199 B.n90 71.676
R2104 B.n203 B.n91 71.676
R2105 B.n207 B.n92 71.676
R2106 B.n211 B.n93 71.676
R2107 B.n215 B.n94 71.676
R2108 B.n219 B.n95 71.676
R2109 B.n223 B.n96 71.676
R2110 B.n227 B.n97 71.676
R2111 B.n231 B.n98 71.676
R2112 B.n235 B.n99 71.676
R2113 B.n239 B.n100 71.676
R2114 B.n243 B.n101 71.676
R2115 B.n247 B.n102 71.676
R2116 B.n251 B.n103 71.676
R2117 B.n255 B.n104 71.676
R2118 B.n259 B.n105 71.676
R2119 B.n263 B.n106 71.676
R2120 B.n267 B.n107 71.676
R2121 B.n271 B.n108 71.676
R2122 B.n275 B.n109 71.676
R2123 B.n279 B.n110 71.676
R2124 B.n283 B.n111 71.676
R2125 B.n287 B.n112 71.676
R2126 B.n291 B.n113 71.676
R2127 B.n295 B.n114 71.676
R2128 B.n299 B.n115 71.676
R2129 B.n303 B.n116 71.676
R2130 B.n307 B.n117 71.676
R2131 B.n311 B.n118 71.676
R2132 B.n315 B.n119 71.676
R2133 B.n319 B.n120 71.676
R2134 B.n323 B.n121 71.676
R2135 B.n327 B.n122 71.676
R2136 B.n331 B.n123 71.676
R2137 B.n335 B.n124 71.676
R2138 B.n339 B.n125 71.676
R2139 B.n343 B.n126 71.676
R2140 B.n347 B.n127 71.676
R2141 B.n351 B.n128 71.676
R2142 B.n355 B.n129 71.676
R2143 B.n359 B.n130 71.676
R2144 B.n363 B.n131 71.676
R2145 B.n367 B.n132 71.676
R2146 B.n371 B.n133 71.676
R2147 B.n375 B.n134 71.676
R2148 B.n379 B.n135 71.676
R2149 B.n383 B.n136 71.676
R2150 B.n387 B.n137 71.676
R2151 B.n963 B.n138 71.676
R2152 B.n963 B.n962 71.676
R2153 B.n389 B.n137 71.676
R2154 B.n386 B.n136 71.676
R2155 B.n382 B.n135 71.676
R2156 B.n378 B.n134 71.676
R2157 B.n374 B.n133 71.676
R2158 B.n370 B.n132 71.676
R2159 B.n366 B.n131 71.676
R2160 B.n362 B.n130 71.676
R2161 B.n358 B.n129 71.676
R2162 B.n354 B.n128 71.676
R2163 B.n350 B.n127 71.676
R2164 B.n346 B.n126 71.676
R2165 B.n342 B.n125 71.676
R2166 B.n338 B.n124 71.676
R2167 B.n334 B.n123 71.676
R2168 B.n330 B.n122 71.676
R2169 B.n326 B.n121 71.676
R2170 B.n322 B.n120 71.676
R2171 B.n318 B.n119 71.676
R2172 B.n314 B.n118 71.676
R2173 B.n310 B.n117 71.676
R2174 B.n306 B.n116 71.676
R2175 B.n302 B.n115 71.676
R2176 B.n298 B.n114 71.676
R2177 B.n294 B.n113 71.676
R2178 B.n290 B.n112 71.676
R2179 B.n286 B.n111 71.676
R2180 B.n282 B.n110 71.676
R2181 B.n278 B.n109 71.676
R2182 B.n274 B.n108 71.676
R2183 B.n270 B.n107 71.676
R2184 B.n266 B.n106 71.676
R2185 B.n262 B.n105 71.676
R2186 B.n258 B.n104 71.676
R2187 B.n254 B.n103 71.676
R2188 B.n250 B.n102 71.676
R2189 B.n246 B.n101 71.676
R2190 B.n242 B.n100 71.676
R2191 B.n238 B.n99 71.676
R2192 B.n234 B.n98 71.676
R2193 B.n230 B.n97 71.676
R2194 B.n226 B.n96 71.676
R2195 B.n222 B.n95 71.676
R2196 B.n218 B.n94 71.676
R2197 B.n214 B.n93 71.676
R2198 B.n210 B.n92 71.676
R2199 B.n206 B.n91 71.676
R2200 B.n202 B.n90 71.676
R2201 B.n198 B.n89 71.676
R2202 B.n194 B.n88 71.676
R2203 B.n190 B.n87 71.676
R2204 B.n186 B.n86 71.676
R2205 B.n182 B.n85 71.676
R2206 B.n178 B.n84 71.676
R2207 B.n174 B.n83 71.676
R2208 B.n170 B.n82 71.676
R2209 B.n166 B.n81 71.676
R2210 B.n162 B.n80 71.676
R2211 B.n158 B.n79 71.676
R2212 B.n154 B.n78 71.676
R2213 B.n150 B.n77 71.676
R2214 B.n146 B.n76 71.676
R2215 B.n536 B.n535 71.676
R2216 B.n538 B.n532 71.676
R2217 B.n545 B.n544 71.676
R2218 B.n546 B.n530 71.676
R2219 B.n553 B.n552 71.676
R2220 B.n554 B.n528 71.676
R2221 B.n561 B.n560 71.676
R2222 B.n562 B.n526 71.676
R2223 B.n569 B.n568 71.676
R2224 B.n570 B.n524 71.676
R2225 B.n577 B.n576 71.676
R2226 B.n578 B.n522 71.676
R2227 B.n585 B.n584 71.676
R2228 B.n586 B.n520 71.676
R2229 B.n593 B.n592 71.676
R2230 B.n594 B.n518 71.676
R2231 B.n601 B.n600 71.676
R2232 B.n602 B.n516 71.676
R2233 B.n609 B.n608 71.676
R2234 B.n610 B.n514 71.676
R2235 B.n617 B.n616 71.676
R2236 B.n618 B.n512 71.676
R2237 B.n625 B.n624 71.676
R2238 B.n626 B.n510 71.676
R2239 B.n633 B.n632 71.676
R2240 B.n634 B.n508 71.676
R2241 B.n641 B.n640 71.676
R2242 B.n642 B.n506 71.676
R2243 B.n652 B.n651 71.676
R2244 B.n653 B.n504 71.676
R2245 B.n660 B.n659 71.676
R2246 B.n661 B.n502 71.676
R2247 B.n668 B.n667 71.676
R2248 B.n669 B.n498 71.676
R2249 B.n677 B.n676 71.676
R2250 B.n678 B.n496 71.676
R2251 B.n685 B.n684 71.676
R2252 B.n686 B.n494 71.676
R2253 B.n693 B.n692 71.676
R2254 B.n694 B.n492 71.676
R2255 B.n701 B.n700 71.676
R2256 B.n702 B.n490 71.676
R2257 B.n709 B.n708 71.676
R2258 B.n710 B.n488 71.676
R2259 B.n717 B.n716 71.676
R2260 B.n718 B.n486 71.676
R2261 B.n725 B.n724 71.676
R2262 B.n726 B.n484 71.676
R2263 B.n733 B.n732 71.676
R2264 B.n734 B.n482 71.676
R2265 B.n741 B.n740 71.676
R2266 B.n742 B.n480 71.676
R2267 B.n749 B.n748 71.676
R2268 B.n750 B.n478 71.676
R2269 B.n757 B.n756 71.676
R2270 B.n758 B.n476 71.676
R2271 B.n765 B.n764 71.676
R2272 B.n766 B.n474 71.676
R2273 B.n773 B.n772 71.676
R2274 B.n774 B.n472 71.676
R2275 B.n781 B.n780 71.676
R2276 B.n784 B.n783 71.676
R2277 B.n789 B.n468 60.9649
R2278 B.n965 B.n964 60.9649
R2279 B.n672 B.n500 59.5399
R2280 B.n648 B.n647 59.5399
R2281 B.n144 B.n143 59.5399
R2282 B.n141 B.n140 59.5399
R2283 B.n500 B.n499 35.1035
R2284 B.n647 B.n646 35.1035
R2285 B.n143 B.n142 35.1035
R2286 B.n140 B.n139 35.1035
R2287 B.n967 B.n73 32.9371
R2288 B.n961 B.n960 32.9371
R2289 B.n787 B.n786 32.9371
R2290 B.n791 B.n466 32.9371
R2291 B.n789 B.n464 32.6429
R2292 B.n795 B.n464 32.6429
R2293 B.n795 B.n460 32.6429
R2294 B.n802 B.n460 32.6429
R2295 B.n802 B.n801 32.6429
R2296 B.n808 B.n453 32.6429
R2297 B.n814 B.n453 32.6429
R2298 B.n814 B.n449 32.6429
R2299 B.n820 B.n449 32.6429
R2300 B.n820 B.n445 32.6429
R2301 B.n826 B.n445 32.6429
R2302 B.n826 B.n441 32.6429
R2303 B.n832 B.n441 32.6429
R2304 B.n838 B.n437 32.6429
R2305 B.n838 B.n432 32.6429
R2306 B.n844 B.n432 32.6429
R2307 B.n844 B.n433 32.6429
R2308 B.n850 B.n425 32.6429
R2309 B.n856 B.n425 32.6429
R2310 B.n856 B.n421 32.6429
R2311 B.n863 B.n421 32.6429
R2312 B.n863 B.n862 32.6429
R2313 B.n869 B.n414 32.6429
R2314 B.n875 B.n414 32.6429
R2315 B.n875 B.n410 32.6429
R2316 B.n881 B.n410 32.6429
R2317 B.n887 B.n406 32.6429
R2318 B.n887 B.n401 32.6429
R2319 B.n893 B.n401 32.6429
R2320 B.n893 B.n402 32.6429
R2321 B.n900 B.n394 32.6429
R2322 B.n906 B.n394 32.6429
R2323 B.n906 B.n4 32.6429
R2324 B.n1045 B.n4 32.6429
R2325 B.n1045 B.n1044 32.6429
R2326 B.n1044 B.n1043 32.6429
R2327 B.n1043 B.n8 32.6429
R2328 B.n1037 B.n8 32.6429
R2329 B.n1036 B.n1035 32.6429
R2330 B.n1035 B.n15 32.6429
R2331 B.n1029 B.n15 32.6429
R2332 B.n1029 B.n1028 32.6429
R2333 B.n1027 B.n22 32.6429
R2334 B.n1021 B.n22 32.6429
R2335 B.n1021 B.n1020 32.6429
R2336 B.n1020 B.n1019 32.6429
R2337 B.n1013 B.n32 32.6429
R2338 B.n1013 B.n1012 32.6429
R2339 B.n1012 B.n1011 32.6429
R2340 B.n1011 B.n36 32.6429
R2341 B.n1005 B.n36 32.6429
R2342 B.n1004 B.n1003 32.6429
R2343 B.n1003 B.n43 32.6429
R2344 B.n997 B.n43 32.6429
R2345 B.n997 B.n996 32.6429
R2346 B.n995 B.n50 32.6429
R2347 B.n989 B.n50 32.6429
R2348 B.n989 B.n988 32.6429
R2349 B.n988 B.n987 32.6429
R2350 B.n987 B.n57 32.6429
R2351 B.n981 B.n57 32.6429
R2352 B.n981 B.n980 32.6429
R2353 B.n980 B.n979 32.6429
R2354 B.n973 B.n67 32.6429
R2355 B.n973 B.n972 32.6429
R2356 B.n972 B.n971 32.6429
R2357 B.n971 B.n71 32.6429
R2358 B.n965 B.n71 32.6429
R2359 B.n801 B.t15 29.7627
R2360 B.n869 B.t0 29.7627
R2361 B.n1019 B.t6 29.7627
R2362 B.n67 B.t11 29.7627
R2363 B.n433 B.t4 24.9623
R2364 B.t9 B.n1004 24.9623
R2365 B.n402 B.t2 24.0022
R2366 B.t7 B.n1036 24.0022
R2367 B.t3 B.n406 19.2019
R2368 B.n1028 B.t1 19.2019
R2369 B.t5 B.n437 18.2418
R2370 B.n996 B.t8 18.2418
R2371 B B.n1047 18.0485
R2372 B.n832 B.t5 14.4015
R2373 B.t8 B.n995 14.4015
R2374 B.n881 B.t3 13.4415
R2375 B.t1 B.n1027 13.4415
R2376 B.n145 B.n73 10.6151
R2377 B.n148 B.n145 10.6151
R2378 B.n149 B.n148 10.6151
R2379 B.n152 B.n149 10.6151
R2380 B.n153 B.n152 10.6151
R2381 B.n156 B.n153 10.6151
R2382 B.n157 B.n156 10.6151
R2383 B.n160 B.n157 10.6151
R2384 B.n161 B.n160 10.6151
R2385 B.n164 B.n161 10.6151
R2386 B.n165 B.n164 10.6151
R2387 B.n168 B.n165 10.6151
R2388 B.n169 B.n168 10.6151
R2389 B.n172 B.n169 10.6151
R2390 B.n173 B.n172 10.6151
R2391 B.n176 B.n173 10.6151
R2392 B.n177 B.n176 10.6151
R2393 B.n180 B.n177 10.6151
R2394 B.n181 B.n180 10.6151
R2395 B.n184 B.n181 10.6151
R2396 B.n185 B.n184 10.6151
R2397 B.n188 B.n185 10.6151
R2398 B.n189 B.n188 10.6151
R2399 B.n192 B.n189 10.6151
R2400 B.n193 B.n192 10.6151
R2401 B.n196 B.n193 10.6151
R2402 B.n197 B.n196 10.6151
R2403 B.n200 B.n197 10.6151
R2404 B.n201 B.n200 10.6151
R2405 B.n204 B.n201 10.6151
R2406 B.n205 B.n204 10.6151
R2407 B.n208 B.n205 10.6151
R2408 B.n209 B.n208 10.6151
R2409 B.n212 B.n209 10.6151
R2410 B.n213 B.n212 10.6151
R2411 B.n216 B.n213 10.6151
R2412 B.n217 B.n216 10.6151
R2413 B.n220 B.n217 10.6151
R2414 B.n221 B.n220 10.6151
R2415 B.n224 B.n221 10.6151
R2416 B.n225 B.n224 10.6151
R2417 B.n228 B.n225 10.6151
R2418 B.n229 B.n228 10.6151
R2419 B.n232 B.n229 10.6151
R2420 B.n233 B.n232 10.6151
R2421 B.n236 B.n233 10.6151
R2422 B.n237 B.n236 10.6151
R2423 B.n240 B.n237 10.6151
R2424 B.n241 B.n240 10.6151
R2425 B.n244 B.n241 10.6151
R2426 B.n245 B.n244 10.6151
R2427 B.n248 B.n245 10.6151
R2428 B.n249 B.n248 10.6151
R2429 B.n252 B.n249 10.6151
R2430 B.n253 B.n252 10.6151
R2431 B.n256 B.n253 10.6151
R2432 B.n257 B.n256 10.6151
R2433 B.n261 B.n260 10.6151
R2434 B.n264 B.n261 10.6151
R2435 B.n265 B.n264 10.6151
R2436 B.n268 B.n265 10.6151
R2437 B.n269 B.n268 10.6151
R2438 B.n272 B.n269 10.6151
R2439 B.n273 B.n272 10.6151
R2440 B.n276 B.n273 10.6151
R2441 B.n277 B.n276 10.6151
R2442 B.n281 B.n280 10.6151
R2443 B.n284 B.n281 10.6151
R2444 B.n285 B.n284 10.6151
R2445 B.n288 B.n285 10.6151
R2446 B.n289 B.n288 10.6151
R2447 B.n292 B.n289 10.6151
R2448 B.n293 B.n292 10.6151
R2449 B.n296 B.n293 10.6151
R2450 B.n297 B.n296 10.6151
R2451 B.n300 B.n297 10.6151
R2452 B.n301 B.n300 10.6151
R2453 B.n304 B.n301 10.6151
R2454 B.n305 B.n304 10.6151
R2455 B.n308 B.n305 10.6151
R2456 B.n309 B.n308 10.6151
R2457 B.n312 B.n309 10.6151
R2458 B.n313 B.n312 10.6151
R2459 B.n316 B.n313 10.6151
R2460 B.n317 B.n316 10.6151
R2461 B.n320 B.n317 10.6151
R2462 B.n321 B.n320 10.6151
R2463 B.n324 B.n321 10.6151
R2464 B.n325 B.n324 10.6151
R2465 B.n328 B.n325 10.6151
R2466 B.n329 B.n328 10.6151
R2467 B.n332 B.n329 10.6151
R2468 B.n333 B.n332 10.6151
R2469 B.n336 B.n333 10.6151
R2470 B.n337 B.n336 10.6151
R2471 B.n340 B.n337 10.6151
R2472 B.n341 B.n340 10.6151
R2473 B.n344 B.n341 10.6151
R2474 B.n345 B.n344 10.6151
R2475 B.n348 B.n345 10.6151
R2476 B.n349 B.n348 10.6151
R2477 B.n352 B.n349 10.6151
R2478 B.n353 B.n352 10.6151
R2479 B.n356 B.n353 10.6151
R2480 B.n357 B.n356 10.6151
R2481 B.n360 B.n357 10.6151
R2482 B.n361 B.n360 10.6151
R2483 B.n364 B.n361 10.6151
R2484 B.n365 B.n364 10.6151
R2485 B.n368 B.n365 10.6151
R2486 B.n369 B.n368 10.6151
R2487 B.n372 B.n369 10.6151
R2488 B.n373 B.n372 10.6151
R2489 B.n376 B.n373 10.6151
R2490 B.n377 B.n376 10.6151
R2491 B.n380 B.n377 10.6151
R2492 B.n381 B.n380 10.6151
R2493 B.n384 B.n381 10.6151
R2494 B.n385 B.n384 10.6151
R2495 B.n388 B.n385 10.6151
R2496 B.n390 B.n388 10.6151
R2497 B.n391 B.n390 10.6151
R2498 B.n961 B.n391 10.6151
R2499 B.n787 B.n462 10.6151
R2500 B.n797 B.n462 10.6151
R2501 B.n798 B.n797 10.6151
R2502 B.n799 B.n798 10.6151
R2503 B.n799 B.n455 10.6151
R2504 B.n810 B.n455 10.6151
R2505 B.n811 B.n810 10.6151
R2506 B.n812 B.n811 10.6151
R2507 B.n812 B.n447 10.6151
R2508 B.n822 B.n447 10.6151
R2509 B.n823 B.n822 10.6151
R2510 B.n824 B.n823 10.6151
R2511 B.n824 B.n439 10.6151
R2512 B.n834 B.n439 10.6151
R2513 B.n835 B.n834 10.6151
R2514 B.n836 B.n835 10.6151
R2515 B.n836 B.n430 10.6151
R2516 B.n846 B.n430 10.6151
R2517 B.n847 B.n846 10.6151
R2518 B.n848 B.n847 10.6151
R2519 B.n848 B.n423 10.6151
R2520 B.n858 B.n423 10.6151
R2521 B.n859 B.n858 10.6151
R2522 B.n860 B.n859 10.6151
R2523 B.n860 B.n416 10.6151
R2524 B.n871 B.n416 10.6151
R2525 B.n872 B.n871 10.6151
R2526 B.n873 B.n872 10.6151
R2527 B.n873 B.n408 10.6151
R2528 B.n883 B.n408 10.6151
R2529 B.n884 B.n883 10.6151
R2530 B.n885 B.n884 10.6151
R2531 B.n885 B.n399 10.6151
R2532 B.n895 B.n399 10.6151
R2533 B.n896 B.n895 10.6151
R2534 B.n898 B.n896 10.6151
R2535 B.n898 B.n897 10.6151
R2536 B.n897 B.n392 10.6151
R2537 B.n909 B.n392 10.6151
R2538 B.n910 B.n909 10.6151
R2539 B.n911 B.n910 10.6151
R2540 B.n912 B.n911 10.6151
R2541 B.n914 B.n912 10.6151
R2542 B.n915 B.n914 10.6151
R2543 B.n916 B.n915 10.6151
R2544 B.n917 B.n916 10.6151
R2545 B.n919 B.n917 10.6151
R2546 B.n920 B.n919 10.6151
R2547 B.n921 B.n920 10.6151
R2548 B.n922 B.n921 10.6151
R2549 B.n924 B.n922 10.6151
R2550 B.n925 B.n924 10.6151
R2551 B.n926 B.n925 10.6151
R2552 B.n927 B.n926 10.6151
R2553 B.n929 B.n927 10.6151
R2554 B.n930 B.n929 10.6151
R2555 B.n931 B.n930 10.6151
R2556 B.n932 B.n931 10.6151
R2557 B.n934 B.n932 10.6151
R2558 B.n935 B.n934 10.6151
R2559 B.n936 B.n935 10.6151
R2560 B.n937 B.n936 10.6151
R2561 B.n939 B.n937 10.6151
R2562 B.n940 B.n939 10.6151
R2563 B.n941 B.n940 10.6151
R2564 B.n942 B.n941 10.6151
R2565 B.n944 B.n942 10.6151
R2566 B.n945 B.n944 10.6151
R2567 B.n946 B.n945 10.6151
R2568 B.n947 B.n946 10.6151
R2569 B.n949 B.n947 10.6151
R2570 B.n950 B.n949 10.6151
R2571 B.n951 B.n950 10.6151
R2572 B.n952 B.n951 10.6151
R2573 B.n954 B.n952 10.6151
R2574 B.n955 B.n954 10.6151
R2575 B.n956 B.n955 10.6151
R2576 B.n957 B.n956 10.6151
R2577 B.n959 B.n957 10.6151
R2578 B.n960 B.n959 10.6151
R2579 B.n534 B.n466 10.6151
R2580 B.n534 B.n533 10.6151
R2581 B.n540 B.n533 10.6151
R2582 B.n541 B.n540 10.6151
R2583 B.n542 B.n541 10.6151
R2584 B.n542 B.n531 10.6151
R2585 B.n548 B.n531 10.6151
R2586 B.n549 B.n548 10.6151
R2587 B.n550 B.n549 10.6151
R2588 B.n550 B.n529 10.6151
R2589 B.n556 B.n529 10.6151
R2590 B.n557 B.n556 10.6151
R2591 B.n558 B.n557 10.6151
R2592 B.n558 B.n527 10.6151
R2593 B.n564 B.n527 10.6151
R2594 B.n565 B.n564 10.6151
R2595 B.n566 B.n565 10.6151
R2596 B.n566 B.n525 10.6151
R2597 B.n572 B.n525 10.6151
R2598 B.n573 B.n572 10.6151
R2599 B.n574 B.n573 10.6151
R2600 B.n574 B.n523 10.6151
R2601 B.n580 B.n523 10.6151
R2602 B.n581 B.n580 10.6151
R2603 B.n582 B.n581 10.6151
R2604 B.n582 B.n521 10.6151
R2605 B.n588 B.n521 10.6151
R2606 B.n589 B.n588 10.6151
R2607 B.n590 B.n589 10.6151
R2608 B.n590 B.n519 10.6151
R2609 B.n596 B.n519 10.6151
R2610 B.n597 B.n596 10.6151
R2611 B.n598 B.n597 10.6151
R2612 B.n598 B.n517 10.6151
R2613 B.n604 B.n517 10.6151
R2614 B.n605 B.n604 10.6151
R2615 B.n606 B.n605 10.6151
R2616 B.n606 B.n515 10.6151
R2617 B.n612 B.n515 10.6151
R2618 B.n613 B.n612 10.6151
R2619 B.n614 B.n613 10.6151
R2620 B.n614 B.n513 10.6151
R2621 B.n620 B.n513 10.6151
R2622 B.n621 B.n620 10.6151
R2623 B.n622 B.n621 10.6151
R2624 B.n622 B.n511 10.6151
R2625 B.n628 B.n511 10.6151
R2626 B.n629 B.n628 10.6151
R2627 B.n630 B.n629 10.6151
R2628 B.n630 B.n509 10.6151
R2629 B.n636 B.n509 10.6151
R2630 B.n637 B.n636 10.6151
R2631 B.n638 B.n637 10.6151
R2632 B.n638 B.n507 10.6151
R2633 B.n644 B.n507 10.6151
R2634 B.n645 B.n644 10.6151
R2635 B.n649 B.n645 10.6151
R2636 B.n655 B.n505 10.6151
R2637 B.n656 B.n655 10.6151
R2638 B.n657 B.n656 10.6151
R2639 B.n657 B.n503 10.6151
R2640 B.n663 B.n503 10.6151
R2641 B.n664 B.n663 10.6151
R2642 B.n665 B.n664 10.6151
R2643 B.n665 B.n501 10.6151
R2644 B.n671 B.n501 10.6151
R2645 B.n674 B.n673 10.6151
R2646 B.n674 B.n497 10.6151
R2647 B.n680 B.n497 10.6151
R2648 B.n681 B.n680 10.6151
R2649 B.n682 B.n681 10.6151
R2650 B.n682 B.n495 10.6151
R2651 B.n688 B.n495 10.6151
R2652 B.n689 B.n688 10.6151
R2653 B.n690 B.n689 10.6151
R2654 B.n690 B.n493 10.6151
R2655 B.n696 B.n493 10.6151
R2656 B.n697 B.n696 10.6151
R2657 B.n698 B.n697 10.6151
R2658 B.n698 B.n491 10.6151
R2659 B.n704 B.n491 10.6151
R2660 B.n705 B.n704 10.6151
R2661 B.n706 B.n705 10.6151
R2662 B.n706 B.n489 10.6151
R2663 B.n712 B.n489 10.6151
R2664 B.n713 B.n712 10.6151
R2665 B.n714 B.n713 10.6151
R2666 B.n714 B.n487 10.6151
R2667 B.n720 B.n487 10.6151
R2668 B.n721 B.n720 10.6151
R2669 B.n722 B.n721 10.6151
R2670 B.n722 B.n485 10.6151
R2671 B.n728 B.n485 10.6151
R2672 B.n729 B.n728 10.6151
R2673 B.n730 B.n729 10.6151
R2674 B.n730 B.n483 10.6151
R2675 B.n736 B.n483 10.6151
R2676 B.n737 B.n736 10.6151
R2677 B.n738 B.n737 10.6151
R2678 B.n738 B.n481 10.6151
R2679 B.n744 B.n481 10.6151
R2680 B.n745 B.n744 10.6151
R2681 B.n746 B.n745 10.6151
R2682 B.n746 B.n479 10.6151
R2683 B.n752 B.n479 10.6151
R2684 B.n753 B.n752 10.6151
R2685 B.n754 B.n753 10.6151
R2686 B.n754 B.n477 10.6151
R2687 B.n760 B.n477 10.6151
R2688 B.n761 B.n760 10.6151
R2689 B.n762 B.n761 10.6151
R2690 B.n762 B.n475 10.6151
R2691 B.n768 B.n475 10.6151
R2692 B.n769 B.n768 10.6151
R2693 B.n770 B.n769 10.6151
R2694 B.n770 B.n473 10.6151
R2695 B.n776 B.n473 10.6151
R2696 B.n777 B.n776 10.6151
R2697 B.n778 B.n777 10.6151
R2698 B.n778 B.n471 10.6151
R2699 B.n471 B.n470 10.6151
R2700 B.n785 B.n470 10.6151
R2701 B.n786 B.n785 10.6151
R2702 B.n792 B.n791 10.6151
R2703 B.n793 B.n792 10.6151
R2704 B.n793 B.n458 10.6151
R2705 B.n804 B.n458 10.6151
R2706 B.n805 B.n804 10.6151
R2707 B.n806 B.n805 10.6151
R2708 B.n806 B.n451 10.6151
R2709 B.n816 B.n451 10.6151
R2710 B.n817 B.n816 10.6151
R2711 B.n818 B.n817 10.6151
R2712 B.n818 B.n443 10.6151
R2713 B.n828 B.n443 10.6151
R2714 B.n829 B.n828 10.6151
R2715 B.n830 B.n829 10.6151
R2716 B.n830 B.n435 10.6151
R2717 B.n840 B.n435 10.6151
R2718 B.n841 B.n840 10.6151
R2719 B.n842 B.n841 10.6151
R2720 B.n842 B.n427 10.6151
R2721 B.n852 B.n427 10.6151
R2722 B.n853 B.n852 10.6151
R2723 B.n854 B.n853 10.6151
R2724 B.n854 B.n419 10.6151
R2725 B.n865 B.n419 10.6151
R2726 B.n866 B.n865 10.6151
R2727 B.n867 B.n866 10.6151
R2728 B.n867 B.n412 10.6151
R2729 B.n877 B.n412 10.6151
R2730 B.n878 B.n877 10.6151
R2731 B.n879 B.n878 10.6151
R2732 B.n879 B.n404 10.6151
R2733 B.n889 B.n404 10.6151
R2734 B.n890 B.n889 10.6151
R2735 B.n891 B.n890 10.6151
R2736 B.n891 B.n396 10.6151
R2737 B.n902 B.n396 10.6151
R2738 B.n903 B.n902 10.6151
R2739 B.n904 B.n903 10.6151
R2740 B.n904 B.n0 10.6151
R2741 B.n1041 B.n1 10.6151
R2742 B.n1041 B.n1040 10.6151
R2743 B.n1040 B.n1039 10.6151
R2744 B.n1039 B.n10 10.6151
R2745 B.n1033 B.n10 10.6151
R2746 B.n1033 B.n1032 10.6151
R2747 B.n1032 B.n1031 10.6151
R2748 B.n1031 B.n17 10.6151
R2749 B.n1025 B.n17 10.6151
R2750 B.n1025 B.n1024 10.6151
R2751 B.n1024 B.n1023 10.6151
R2752 B.n1023 B.n24 10.6151
R2753 B.n1017 B.n24 10.6151
R2754 B.n1017 B.n1016 10.6151
R2755 B.n1016 B.n1015 10.6151
R2756 B.n1015 B.n30 10.6151
R2757 B.n1009 B.n30 10.6151
R2758 B.n1009 B.n1008 10.6151
R2759 B.n1008 B.n1007 10.6151
R2760 B.n1007 B.n38 10.6151
R2761 B.n1001 B.n38 10.6151
R2762 B.n1001 B.n1000 10.6151
R2763 B.n1000 B.n999 10.6151
R2764 B.n999 B.n45 10.6151
R2765 B.n993 B.n45 10.6151
R2766 B.n993 B.n992 10.6151
R2767 B.n992 B.n991 10.6151
R2768 B.n991 B.n52 10.6151
R2769 B.n985 B.n52 10.6151
R2770 B.n985 B.n984 10.6151
R2771 B.n984 B.n983 10.6151
R2772 B.n983 B.n59 10.6151
R2773 B.n977 B.n59 10.6151
R2774 B.n977 B.n976 10.6151
R2775 B.n976 B.n975 10.6151
R2776 B.n975 B.n65 10.6151
R2777 B.n969 B.n65 10.6151
R2778 B.n969 B.n968 10.6151
R2779 B.n968 B.n967 10.6151
R2780 B.n257 B.n144 9.36635
R2781 B.n280 B.n141 9.36635
R2782 B.n649 B.n648 9.36635
R2783 B.n673 B.n672 9.36635
R2784 B.n900 B.t2 8.64113
R2785 B.n1037 B.t7 8.64113
R2786 B.n850 B.t4 7.68106
R2787 B.n1005 B.t9 7.68106
R2788 B.n808 B.t15 2.88071
R2789 B.n862 B.t0 2.88071
R2790 B.n32 B.t6 2.88071
R2791 B.n979 B.t11 2.88071
R2792 B.n1047 B.n0 2.81026
R2793 B.n1047 B.n1 2.81026
R2794 B.n260 B.n144 1.24928
R2795 B.n277 B.n141 1.24928
R2796 B.n648 B.n505 1.24928
R2797 B.n672 B.n671 1.24928
R2798 VP.n15 VP.t9 318.837
R2799 VP.n48 VP.t3 287.247
R2800 VP.n35 VP.t4 287.247
R2801 VP.n41 VP.t2 287.247
R2802 VP.n54 VP.t6 287.247
R2803 VP.n61 VP.t5 287.247
R2804 VP.n20 VP.t8 287.247
R2805 VP.n33 VP.t0 287.247
R2806 VP.n26 VP.t1 287.247
R2807 VP.n14 VP.t7 287.247
R2808 VP.n36 VP.n35 179.99
R2809 VP.n62 VP.n61 179.99
R2810 VP.n34 VP.n33 179.99
R2811 VP.n16 VP.n13 161.3
R2812 VP.n18 VP.n17 161.3
R2813 VP.n19 VP.n12 161.3
R2814 VP.n21 VP.n20 161.3
R2815 VP.n22 VP.n11 161.3
R2816 VP.n24 VP.n23 161.3
R2817 VP.n25 VP.n10 161.3
R2818 VP.n28 VP.n27 161.3
R2819 VP.n29 VP.n9 161.3
R2820 VP.n31 VP.n30 161.3
R2821 VP.n32 VP.n8 161.3
R2822 VP.n60 VP.n0 161.3
R2823 VP.n59 VP.n58 161.3
R2824 VP.n57 VP.n1 161.3
R2825 VP.n56 VP.n55 161.3
R2826 VP.n53 VP.n2 161.3
R2827 VP.n52 VP.n51 161.3
R2828 VP.n50 VP.n3 161.3
R2829 VP.n49 VP.n48 161.3
R2830 VP.n47 VP.n4 161.3
R2831 VP.n46 VP.n45 161.3
R2832 VP.n44 VP.n5 161.3
R2833 VP.n43 VP.n42 161.3
R2834 VP.n40 VP.n6 161.3
R2835 VP.n39 VP.n38 161.3
R2836 VP.n37 VP.n7 161.3
R2837 VP.n40 VP.n39 56.5617
R2838 VP.n31 VP.n9 56.5617
R2839 VP.n59 VP.n1 56.5617
R2840 VP.n36 VP.n34 51.1558
R2841 VP.n15 VP.n14 50.9283
R2842 VP.n47 VP.n46 49.7803
R2843 VP.n52 VP.n3 49.7803
R2844 VP.n24 VP.n11 49.7803
R2845 VP.n19 VP.n18 49.7803
R2846 VP.n46 VP.n5 31.3737
R2847 VP.n53 VP.n52 31.3737
R2848 VP.n25 VP.n24 31.3737
R2849 VP.n18 VP.n13 31.3737
R2850 VP.n39 VP.n7 24.5923
R2851 VP.n42 VP.n40 24.5923
R2852 VP.n48 VP.n47 24.5923
R2853 VP.n48 VP.n3 24.5923
R2854 VP.n55 VP.n1 24.5923
R2855 VP.n60 VP.n59 24.5923
R2856 VP.n32 VP.n31 24.5923
R2857 VP.n27 VP.n9 24.5923
R2858 VP.n20 VP.n19 24.5923
R2859 VP.n20 VP.n11 24.5923
R2860 VP.n16 VP.n15 18.1684
R2861 VP.n41 VP.n5 15.2474
R2862 VP.n54 VP.n53 15.2474
R2863 VP.n26 VP.n25 15.2474
R2864 VP.n14 VP.n13 15.2474
R2865 VP.n42 VP.n41 9.3454
R2866 VP.n55 VP.n54 9.3454
R2867 VP.n27 VP.n26 9.3454
R2868 VP.n35 VP.n7 5.90254
R2869 VP.n61 VP.n60 5.90254
R2870 VP.n33 VP.n32 5.90254
R2871 VP.n17 VP.n16 0.189894
R2872 VP.n17 VP.n12 0.189894
R2873 VP.n21 VP.n12 0.189894
R2874 VP.n22 VP.n21 0.189894
R2875 VP.n23 VP.n22 0.189894
R2876 VP.n23 VP.n10 0.189894
R2877 VP.n28 VP.n10 0.189894
R2878 VP.n29 VP.n28 0.189894
R2879 VP.n30 VP.n29 0.189894
R2880 VP.n30 VP.n8 0.189894
R2881 VP.n34 VP.n8 0.189894
R2882 VP.n37 VP.n36 0.189894
R2883 VP.n38 VP.n37 0.189894
R2884 VP.n38 VP.n6 0.189894
R2885 VP.n43 VP.n6 0.189894
R2886 VP.n44 VP.n43 0.189894
R2887 VP.n45 VP.n44 0.189894
R2888 VP.n45 VP.n4 0.189894
R2889 VP.n49 VP.n4 0.189894
R2890 VP.n50 VP.n49 0.189894
R2891 VP.n51 VP.n50 0.189894
R2892 VP.n51 VP.n2 0.189894
R2893 VP.n56 VP.n2 0.189894
R2894 VP.n57 VP.n56 0.189894
R2895 VP.n58 VP.n57 0.189894
R2896 VP.n58 VP.n0 0.189894
R2897 VP.n62 VP.n0 0.189894
R2898 VP VP.n62 0.0516364
R2899 VDD1.n92 VDD1.n0 289.615
R2900 VDD1.n191 VDD1.n99 289.615
R2901 VDD1.n93 VDD1.n92 185
R2902 VDD1.n91 VDD1.n90 185
R2903 VDD1.n4 VDD1.n3 185
R2904 VDD1.n85 VDD1.n84 185
R2905 VDD1.n83 VDD1.n82 185
R2906 VDD1.n8 VDD1.n7 185
R2907 VDD1.n12 VDD1.n10 185
R2908 VDD1.n77 VDD1.n76 185
R2909 VDD1.n75 VDD1.n74 185
R2910 VDD1.n14 VDD1.n13 185
R2911 VDD1.n69 VDD1.n68 185
R2912 VDD1.n67 VDD1.n66 185
R2913 VDD1.n18 VDD1.n17 185
R2914 VDD1.n61 VDD1.n60 185
R2915 VDD1.n59 VDD1.n58 185
R2916 VDD1.n22 VDD1.n21 185
R2917 VDD1.n53 VDD1.n52 185
R2918 VDD1.n51 VDD1.n50 185
R2919 VDD1.n26 VDD1.n25 185
R2920 VDD1.n45 VDD1.n44 185
R2921 VDD1.n43 VDD1.n42 185
R2922 VDD1.n30 VDD1.n29 185
R2923 VDD1.n37 VDD1.n36 185
R2924 VDD1.n35 VDD1.n34 185
R2925 VDD1.n132 VDD1.n131 185
R2926 VDD1.n134 VDD1.n133 185
R2927 VDD1.n127 VDD1.n126 185
R2928 VDD1.n140 VDD1.n139 185
R2929 VDD1.n142 VDD1.n141 185
R2930 VDD1.n123 VDD1.n122 185
R2931 VDD1.n148 VDD1.n147 185
R2932 VDD1.n150 VDD1.n149 185
R2933 VDD1.n119 VDD1.n118 185
R2934 VDD1.n156 VDD1.n155 185
R2935 VDD1.n158 VDD1.n157 185
R2936 VDD1.n115 VDD1.n114 185
R2937 VDD1.n164 VDD1.n163 185
R2938 VDD1.n166 VDD1.n165 185
R2939 VDD1.n111 VDD1.n110 185
R2940 VDD1.n173 VDD1.n172 185
R2941 VDD1.n174 VDD1.n109 185
R2942 VDD1.n176 VDD1.n175 185
R2943 VDD1.n107 VDD1.n106 185
R2944 VDD1.n182 VDD1.n181 185
R2945 VDD1.n184 VDD1.n183 185
R2946 VDD1.n103 VDD1.n102 185
R2947 VDD1.n190 VDD1.n189 185
R2948 VDD1.n192 VDD1.n191 185
R2949 VDD1.n33 VDD1.t0 147.659
R2950 VDD1.n130 VDD1.t5 147.659
R2951 VDD1.n92 VDD1.n91 104.615
R2952 VDD1.n91 VDD1.n3 104.615
R2953 VDD1.n84 VDD1.n3 104.615
R2954 VDD1.n84 VDD1.n83 104.615
R2955 VDD1.n83 VDD1.n7 104.615
R2956 VDD1.n12 VDD1.n7 104.615
R2957 VDD1.n76 VDD1.n12 104.615
R2958 VDD1.n76 VDD1.n75 104.615
R2959 VDD1.n75 VDD1.n13 104.615
R2960 VDD1.n68 VDD1.n13 104.615
R2961 VDD1.n68 VDD1.n67 104.615
R2962 VDD1.n67 VDD1.n17 104.615
R2963 VDD1.n60 VDD1.n17 104.615
R2964 VDD1.n60 VDD1.n59 104.615
R2965 VDD1.n59 VDD1.n21 104.615
R2966 VDD1.n52 VDD1.n21 104.615
R2967 VDD1.n52 VDD1.n51 104.615
R2968 VDD1.n51 VDD1.n25 104.615
R2969 VDD1.n44 VDD1.n25 104.615
R2970 VDD1.n44 VDD1.n43 104.615
R2971 VDD1.n43 VDD1.n29 104.615
R2972 VDD1.n36 VDD1.n29 104.615
R2973 VDD1.n36 VDD1.n35 104.615
R2974 VDD1.n133 VDD1.n132 104.615
R2975 VDD1.n133 VDD1.n126 104.615
R2976 VDD1.n140 VDD1.n126 104.615
R2977 VDD1.n141 VDD1.n140 104.615
R2978 VDD1.n141 VDD1.n122 104.615
R2979 VDD1.n148 VDD1.n122 104.615
R2980 VDD1.n149 VDD1.n148 104.615
R2981 VDD1.n149 VDD1.n118 104.615
R2982 VDD1.n156 VDD1.n118 104.615
R2983 VDD1.n157 VDD1.n156 104.615
R2984 VDD1.n157 VDD1.n114 104.615
R2985 VDD1.n164 VDD1.n114 104.615
R2986 VDD1.n165 VDD1.n164 104.615
R2987 VDD1.n165 VDD1.n110 104.615
R2988 VDD1.n173 VDD1.n110 104.615
R2989 VDD1.n174 VDD1.n173 104.615
R2990 VDD1.n175 VDD1.n174 104.615
R2991 VDD1.n175 VDD1.n106 104.615
R2992 VDD1.n182 VDD1.n106 104.615
R2993 VDD1.n183 VDD1.n182 104.615
R2994 VDD1.n183 VDD1.n102 104.615
R2995 VDD1.n190 VDD1.n102 104.615
R2996 VDD1.n191 VDD1.n190 104.615
R2997 VDD1.n199 VDD1.n198 64.1242
R2998 VDD1.n98 VDD1.n97 63.0094
R2999 VDD1.n197 VDD1.n196 63.0093
R3000 VDD1.n201 VDD1.n200 63.0092
R3001 VDD1.n98 VDD1.n96 52.7518
R3002 VDD1.n197 VDD1.n195 52.7518
R3003 VDD1.n35 VDD1.t0 52.3082
R3004 VDD1.n132 VDD1.t5 52.3082
R3005 VDD1.n201 VDD1.n199 47.697
R3006 VDD1.n34 VDD1.n33 15.6677
R3007 VDD1.n131 VDD1.n130 15.6677
R3008 VDD1.n10 VDD1.n8 13.1884
R3009 VDD1.n176 VDD1.n107 13.1884
R3010 VDD1.n82 VDD1.n81 12.8005
R3011 VDD1.n78 VDD1.n77 12.8005
R3012 VDD1.n37 VDD1.n32 12.8005
R3013 VDD1.n134 VDD1.n129 12.8005
R3014 VDD1.n177 VDD1.n109 12.8005
R3015 VDD1.n181 VDD1.n180 12.8005
R3016 VDD1.n85 VDD1.n6 12.0247
R3017 VDD1.n74 VDD1.n11 12.0247
R3018 VDD1.n38 VDD1.n30 12.0247
R3019 VDD1.n135 VDD1.n127 12.0247
R3020 VDD1.n172 VDD1.n171 12.0247
R3021 VDD1.n184 VDD1.n105 12.0247
R3022 VDD1.n86 VDD1.n4 11.249
R3023 VDD1.n73 VDD1.n14 11.249
R3024 VDD1.n42 VDD1.n41 11.249
R3025 VDD1.n139 VDD1.n138 11.249
R3026 VDD1.n170 VDD1.n111 11.249
R3027 VDD1.n185 VDD1.n103 11.249
R3028 VDD1.n90 VDD1.n89 10.4732
R3029 VDD1.n70 VDD1.n69 10.4732
R3030 VDD1.n45 VDD1.n28 10.4732
R3031 VDD1.n142 VDD1.n125 10.4732
R3032 VDD1.n167 VDD1.n166 10.4732
R3033 VDD1.n189 VDD1.n188 10.4732
R3034 VDD1.n93 VDD1.n2 9.69747
R3035 VDD1.n66 VDD1.n16 9.69747
R3036 VDD1.n46 VDD1.n26 9.69747
R3037 VDD1.n143 VDD1.n123 9.69747
R3038 VDD1.n163 VDD1.n113 9.69747
R3039 VDD1.n192 VDD1.n101 9.69747
R3040 VDD1.n96 VDD1.n95 9.45567
R3041 VDD1.n195 VDD1.n194 9.45567
R3042 VDD1.n20 VDD1.n19 9.3005
R3043 VDD1.n63 VDD1.n62 9.3005
R3044 VDD1.n65 VDD1.n64 9.3005
R3045 VDD1.n16 VDD1.n15 9.3005
R3046 VDD1.n71 VDD1.n70 9.3005
R3047 VDD1.n73 VDD1.n72 9.3005
R3048 VDD1.n11 VDD1.n9 9.3005
R3049 VDD1.n79 VDD1.n78 9.3005
R3050 VDD1.n95 VDD1.n94 9.3005
R3051 VDD1.n2 VDD1.n1 9.3005
R3052 VDD1.n89 VDD1.n88 9.3005
R3053 VDD1.n87 VDD1.n86 9.3005
R3054 VDD1.n6 VDD1.n5 9.3005
R3055 VDD1.n81 VDD1.n80 9.3005
R3056 VDD1.n57 VDD1.n56 9.3005
R3057 VDD1.n55 VDD1.n54 9.3005
R3058 VDD1.n24 VDD1.n23 9.3005
R3059 VDD1.n49 VDD1.n48 9.3005
R3060 VDD1.n47 VDD1.n46 9.3005
R3061 VDD1.n28 VDD1.n27 9.3005
R3062 VDD1.n41 VDD1.n40 9.3005
R3063 VDD1.n39 VDD1.n38 9.3005
R3064 VDD1.n32 VDD1.n31 9.3005
R3065 VDD1.n194 VDD1.n193 9.3005
R3066 VDD1.n101 VDD1.n100 9.3005
R3067 VDD1.n188 VDD1.n187 9.3005
R3068 VDD1.n186 VDD1.n185 9.3005
R3069 VDD1.n105 VDD1.n104 9.3005
R3070 VDD1.n180 VDD1.n179 9.3005
R3071 VDD1.n152 VDD1.n151 9.3005
R3072 VDD1.n121 VDD1.n120 9.3005
R3073 VDD1.n146 VDD1.n145 9.3005
R3074 VDD1.n144 VDD1.n143 9.3005
R3075 VDD1.n125 VDD1.n124 9.3005
R3076 VDD1.n138 VDD1.n137 9.3005
R3077 VDD1.n136 VDD1.n135 9.3005
R3078 VDD1.n129 VDD1.n128 9.3005
R3079 VDD1.n154 VDD1.n153 9.3005
R3080 VDD1.n117 VDD1.n116 9.3005
R3081 VDD1.n160 VDD1.n159 9.3005
R3082 VDD1.n162 VDD1.n161 9.3005
R3083 VDD1.n113 VDD1.n112 9.3005
R3084 VDD1.n168 VDD1.n167 9.3005
R3085 VDD1.n170 VDD1.n169 9.3005
R3086 VDD1.n171 VDD1.n108 9.3005
R3087 VDD1.n178 VDD1.n177 9.3005
R3088 VDD1.n94 VDD1.n0 8.92171
R3089 VDD1.n65 VDD1.n18 8.92171
R3090 VDD1.n50 VDD1.n49 8.92171
R3091 VDD1.n147 VDD1.n146 8.92171
R3092 VDD1.n162 VDD1.n115 8.92171
R3093 VDD1.n193 VDD1.n99 8.92171
R3094 VDD1.n62 VDD1.n61 8.14595
R3095 VDD1.n53 VDD1.n24 8.14595
R3096 VDD1.n150 VDD1.n121 8.14595
R3097 VDD1.n159 VDD1.n158 8.14595
R3098 VDD1.n58 VDD1.n20 7.3702
R3099 VDD1.n54 VDD1.n22 7.3702
R3100 VDD1.n151 VDD1.n119 7.3702
R3101 VDD1.n155 VDD1.n117 7.3702
R3102 VDD1.n58 VDD1.n57 6.59444
R3103 VDD1.n57 VDD1.n22 6.59444
R3104 VDD1.n154 VDD1.n119 6.59444
R3105 VDD1.n155 VDD1.n154 6.59444
R3106 VDD1.n61 VDD1.n20 5.81868
R3107 VDD1.n54 VDD1.n53 5.81868
R3108 VDD1.n151 VDD1.n150 5.81868
R3109 VDD1.n158 VDD1.n117 5.81868
R3110 VDD1.n96 VDD1.n0 5.04292
R3111 VDD1.n62 VDD1.n18 5.04292
R3112 VDD1.n50 VDD1.n24 5.04292
R3113 VDD1.n147 VDD1.n121 5.04292
R3114 VDD1.n159 VDD1.n115 5.04292
R3115 VDD1.n195 VDD1.n99 5.04292
R3116 VDD1.n33 VDD1.n31 4.38563
R3117 VDD1.n130 VDD1.n128 4.38563
R3118 VDD1.n94 VDD1.n93 4.26717
R3119 VDD1.n66 VDD1.n65 4.26717
R3120 VDD1.n49 VDD1.n26 4.26717
R3121 VDD1.n146 VDD1.n123 4.26717
R3122 VDD1.n163 VDD1.n162 4.26717
R3123 VDD1.n193 VDD1.n192 4.26717
R3124 VDD1.n90 VDD1.n2 3.49141
R3125 VDD1.n69 VDD1.n16 3.49141
R3126 VDD1.n46 VDD1.n45 3.49141
R3127 VDD1.n143 VDD1.n142 3.49141
R3128 VDD1.n166 VDD1.n113 3.49141
R3129 VDD1.n189 VDD1.n101 3.49141
R3130 VDD1.n89 VDD1.n4 2.71565
R3131 VDD1.n70 VDD1.n14 2.71565
R3132 VDD1.n42 VDD1.n28 2.71565
R3133 VDD1.n139 VDD1.n125 2.71565
R3134 VDD1.n167 VDD1.n111 2.71565
R3135 VDD1.n188 VDD1.n103 2.71565
R3136 VDD1.n86 VDD1.n85 1.93989
R3137 VDD1.n74 VDD1.n73 1.93989
R3138 VDD1.n41 VDD1.n30 1.93989
R3139 VDD1.n138 VDD1.n127 1.93989
R3140 VDD1.n172 VDD1.n170 1.93989
R3141 VDD1.n185 VDD1.n184 1.93989
R3142 VDD1.n82 VDD1.n6 1.16414
R3143 VDD1.n77 VDD1.n11 1.16414
R3144 VDD1.n38 VDD1.n37 1.16414
R3145 VDD1.n135 VDD1.n134 1.16414
R3146 VDD1.n171 VDD1.n109 1.16414
R3147 VDD1.n181 VDD1.n105 1.16414
R3148 VDD1.n200 VDD1.t8 1.12295
R3149 VDD1.n200 VDD1.t9 1.12295
R3150 VDD1.n97 VDD1.t2 1.12295
R3151 VDD1.n97 VDD1.t1 1.12295
R3152 VDD1.n198 VDD1.t3 1.12295
R3153 VDD1.n198 VDD1.t4 1.12295
R3154 VDD1.n196 VDD1.t7 1.12295
R3155 VDD1.n196 VDD1.t6 1.12295
R3156 VDD1 VDD1.n201 1.11257
R3157 VDD1 VDD1.n98 0.448776
R3158 VDD1.n81 VDD1.n8 0.388379
R3159 VDD1.n78 VDD1.n10 0.388379
R3160 VDD1.n34 VDD1.n32 0.388379
R3161 VDD1.n131 VDD1.n129 0.388379
R3162 VDD1.n177 VDD1.n176 0.388379
R3163 VDD1.n180 VDD1.n107 0.388379
R3164 VDD1.n199 VDD1.n197 0.33524
R3165 VDD1.n95 VDD1.n1 0.155672
R3166 VDD1.n88 VDD1.n1 0.155672
R3167 VDD1.n88 VDD1.n87 0.155672
R3168 VDD1.n87 VDD1.n5 0.155672
R3169 VDD1.n80 VDD1.n5 0.155672
R3170 VDD1.n80 VDD1.n79 0.155672
R3171 VDD1.n79 VDD1.n9 0.155672
R3172 VDD1.n72 VDD1.n9 0.155672
R3173 VDD1.n72 VDD1.n71 0.155672
R3174 VDD1.n71 VDD1.n15 0.155672
R3175 VDD1.n64 VDD1.n15 0.155672
R3176 VDD1.n64 VDD1.n63 0.155672
R3177 VDD1.n63 VDD1.n19 0.155672
R3178 VDD1.n56 VDD1.n19 0.155672
R3179 VDD1.n56 VDD1.n55 0.155672
R3180 VDD1.n55 VDD1.n23 0.155672
R3181 VDD1.n48 VDD1.n23 0.155672
R3182 VDD1.n48 VDD1.n47 0.155672
R3183 VDD1.n47 VDD1.n27 0.155672
R3184 VDD1.n40 VDD1.n27 0.155672
R3185 VDD1.n40 VDD1.n39 0.155672
R3186 VDD1.n39 VDD1.n31 0.155672
R3187 VDD1.n136 VDD1.n128 0.155672
R3188 VDD1.n137 VDD1.n136 0.155672
R3189 VDD1.n137 VDD1.n124 0.155672
R3190 VDD1.n144 VDD1.n124 0.155672
R3191 VDD1.n145 VDD1.n144 0.155672
R3192 VDD1.n145 VDD1.n120 0.155672
R3193 VDD1.n152 VDD1.n120 0.155672
R3194 VDD1.n153 VDD1.n152 0.155672
R3195 VDD1.n153 VDD1.n116 0.155672
R3196 VDD1.n160 VDD1.n116 0.155672
R3197 VDD1.n161 VDD1.n160 0.155672
R3198 VDD1.n161 VDD1.n112 0.155672
R3199 VDD1.n168 VDD1.n112 0.155672
R3200 VDD1.n169 VDD1.n168 0.155672
R3201 VDD1.n169 VDD1.n108 0.155672
R3202 VDD1.n178 VDD1.n108 0.155672
R3203 VDD1.n179 VDD1.n178 0.155672
R3204 VDD1.n179 VDD1.n104 0.155672
R3205 VDD1.n186 VDD1.n104 0.155672
R3206 VDD1.n187 VDD1.n186 0.155672
R3207 VDD1.n187 VDD1.n100 0.155672
R3208 VDD1.n194 VDD1.n100 0.155672
C0 VDD1 VP 13.6101f
C1 VDD2 VP 0.441804f
C2 VN VTAIL 13.272901f
C3 VDD1 VN 0.15114f
C4 VDD1 VTAIL 14.477901f
C5 VDD2 VN 13.324901f
C6 VN VP 7.78971f
C7 VDD2 VTAIL 14.517499f
C8 VTAIL VP 13.287499f
C9 VDD1 VDD2 1.44738f
C10 VDD2 B 6.897394f
C11 VDD1 B 6.870593f
C12 VTAIL B 9.441069f
C13 VN B 13.4579f
C14 VP B 11.636939f
C15 VDD1.n0 B 0.032883f
C16 VDD1.n1 B 0.022529f
C17 VDD1.n2 B 0.012106f
C18 VDD1.n3 B 0.028615f
C19 VDD1.n4 B 0.012818f
C20 VDD1.n5 B 0.022529f
C21 VDD1.n6 B 0.012106f
C22 VDD1.n7 B 0.028615f
C23 VDD1.n8 B 0.012462f
C24 VDD1.n9 B 0.022529f
C25 VDD1.n10 B 0.012462f
C26 VDD1.n11 B 0.012106f
C27 VDD1.n12 B 0.028615f
C28 VDD1.n13 B 0.028615f
C29 VDD1.n14 B 0.012818f
C30 VDD1.n15 B 0.022529f
C31 VDD1.n16 B 0.012106f
C32 VDD1.n17 B 0.028615f
C33 VDD1.n18 B 0.012818f
C34 VDD1.n19 B 0.022529f
C35 VDD1.n20 B 0.012106f
C36 VDD1.n21 B 0.028615f
C37 VDD1.n22 B 0.012818f
C38 VDD1.n23 B 0.022529f
C39 VDD1.n24 B 0.012106f
C40 VDD1.n25 B 0.028615f
C41 VDD1.n26 B 0.012818f
C42 VDD1.n27 B 0.022529f
C43 VDD1.n28 B 0.012106f
C44 VDD1.n29 B 0.028615f
C45 VDD1.n30 B 0.012818f
C46 VDD1.n31 B 1.73838f
C47 VDD1.n32 B 0.012106f
C48 VDD1.t0 B 0.047387f
C49 VDD1.n33 B 0.161854f
C50 VDD1.n34 B 0.016904f
C51 VDD1.n35 B 0.021461f
C52 VDD1.n36 B 0.028615f
C53 VDD1.n37 B 0.012818f
C54 VDD1.n38 B 0.012106f
C55 VDD1.n39 B 0.022529f
C56 VDD1.n40 B 0.022529f
C57 VDD1.n41 B 0.012106f
C58 VDD1.n42 B 0.012818f
C59 VDD1.n43 B 0.028615f
C60 VDD1.n44 B 0.028615f
C61 VDD1.n45 B 0.012818f
C62 VDD1.n46 B 0.012106f
C63 VDD1.n47 B 0.022529f
C64 VDD1.n48 B 0.022529f
C65 VDD1.n49 B 0.012106f
C66 VDD1.n50 B 0.012818f
C67 VDD1.n51 B 0.028615f
C68 VDD1.n52 B 0.028615f
C69 VDD1.n53 B 0.012818f
C70 VDD1.n54 B 0.012106f
C71 VDD1.n55 B 0.022529f
C72 VDD1.n56 B 0.022529f
C73 VDD1.n57 B 0.012106f
C74 VDD1.n58 B 0.012818f
C75 VDD1.n59 B 0.028615f
C76 VDD1.n60 B 0.028615f
C77 VDD1.n61 B 0.012818f
C78 VDD1.n62 B 0.012106f
C79 VDD1.n63 B 0.022529f
C80 VDD1.n64 B 0.022529f
C81 VDD1.n65 B 0.012106f
C82 VDD1.n66 B 0.012818f
C83 VDD1.n67 B 0.028615f
C84 VDD1.n68 B 0.028615f
C85 VDD1.n69 B 0.012818f
C86 VDD1.n70 B 0.012106f
C87 VDD1.n71 B 0.022529f
C88 VDD1.n72 B 0.022529f
C89 VDD1.n73 B 0.012106f
C90 VDD1.n74 B 0.012818f
C91 VDD1.n75 B 0.028615f
C92 VDD1.n76 B 0.028615f
C93 VDD1.n77 B 0.012818f
C94 VDD1.n78 B 0.012106f
C95 VDD1.n79 B 0.022529f
C96 VDD1.n80 B 0.022529f
C97 VDD1.n81 B 0.012106f
C98 VDD1.n82 B 0.012818f
C99 VDD1.n83 B 0.028615f
C100 VDD1.n84 B 0.028615f
C101 VDD1.n85 B 0.012818f
C102 VDD1.n86 B 0.012106f
C103 VDD1.n87 B 0.022529f
C104 VDD1.n88 B 0.022529f
C105 VDD1.n89 B 0.012106f
C106 VDD1.n90 B 0.012818f
C107 VDD1.n91 B 0.028615f
C108 VDD1.n92 B 0.064097f
C109 VDD1.n93 B 0.012818f
C110 VDD1.n94 B 0.012106f
C111 VDD1.n95 B 0.055769f
C112 VDD1.n96 B 0.056421f
C113 VDD1.t2 B 0.314052f
C114 VDD1.t1 B 0.314052f
C115 VDD1.n97 B 2.86098f
C116 VDD1.n98 B 0.484481f
C117 VDD1.n99 B 0.032883f
C118 VDD1.n100 B 0.022529f
C119 VDD1.n101 B 0.012106f
C120 VDD1.n102 B 0.028615f
C121 VDD1.n103 B 0.012818f
C122 VDD1.n104 B 0.022529f
C123 VDD1.n105 B 0.012106f
C124 VDD1.n106 B 0.028615f
C125 VDD1.n107 B 0.012462f
C126 VDD1.n108 B 0.022529f
C127 VDD1.n109 B 0.012818f
C128 VDD1.n110 B 0.028615f
C129 VDD1.n111 B 0.012818f
C130 VDD1.n112 B 0.022529f
C131 VDD1.n113 B 0.012106f
C132 VDD1.n114 B 0.028615f
C133 VDD1.n115 B 0.012818f
C134 VDD1.n116 B 0.022529f
C135 VDD1.n117 B 0.012106f
C136 VDD1.n118 B 0.028615f
C137 VDD1.n119 B 0.012818f
C138 VDD1.n120 B 0.022529f
C139 VDD1.n121 B 0.012106f
C140 VDD1.n122 B 0.028615f
C141 VDD1.n123 B 0.012818f
C142 VDD1.n124 B 0.022529f
C143 VDD1.n125 B 0.012106f
C144 VDD1.n126 B 0.028615f
C145 VDD1.n127 B 0.012818f
C146 VDD1.n128 B 1.73838f
C147 VDD1.n129 B 0.012106f
C148 VDD1.t5 B 0.047387f
C149 VDD1.n130 B 0.161854f
C150 VDD1.n131 B 0.016904f
C151 VDD1.n132 B 0.021461f
C152 VDD1.n133 B 0.028615f
C153 VDD1.n134 B 0.012818f
C154 VDD1.n135 B 0.012106f
C155 VDD1.n136 B 0.022529f
C156 VDD1.n137 B 0.022529f
C157 VDD1.n138 B 0.012106f
C158 VDD1.n139 B 0.012818f
C159 VDD1.n140 B 0.028615f
C160 VDD1.n141 B 0.028615f
C161 VDD1.n142 B 0.012818f
C162 VDD1.n143 B 0.012106f
C163 VDD1.n144 B 0.022529f
C164 VDD1.n145 B 0.022529f
C165 VDD1.n146 B 0.012106f
C166 VDD1.n147 B 0.012818f
C167 VDD1.n148 B 0.028615f
C168 VDD1.n149 B 0.028615f
C169 VDD1.n150 B 0.012818f
C170 VDD1.n151 B 0.012106f
C171 VDD1.n152 B 0.022529f
C172 VDD1.n153 B 0.022529f
C173 VDD1.n154 B 0.012106f
C174 VDD1.n155 B 0.012818f
C175 VDD1.n156 B 0.028615f
C176 VDD1.n157 B 0.028615f
C177 VDD1.n158 B 0.012818f
C178 VDD1.n159 B 0.012106f
C179 VDD1.n160 B 0.022529f
C180 VDD1.n161 B 0.022529f
C181 VDD1.n162 B 0.012106f
C182 VDD1.n163 B 0.012818f
C183 VDD1.n164 B 0.028615f
C184 VDD1.n165 B 0.028615f
C185 VDD1.n166 B 0.012818f
C186 VDD1.n167 B 0.012106f
C187 VDD1.n168 B 0.022529f
C188 VDD1.n169 B 0.022529f
C189 VDD1.n170 B 0.012106f
C190 VDD1.n171 B 0.012106f
C191 VDD1.n172 B 0.012818f
C192 VDD1.n173 B 0.028615f
C193 VDD1.n174 B 0.028615f
C194 VDD1.n175 B 0.028615f
C195 VDD1.n176 B 0.012462f
C196 VDD1.n177 B 0.012106f
C197 VDD1.n178 B 0.022529f
C198 VDD1.n179 B 0.022529f
C199 VDD1.n180 B 0.012106f
C200 VDD1.n181 B 0.012818f
C201 VDD1.n182 B 0.028615f
C202 VDD1.n183 B 0.028615f
C203 VDD1.n184 B 0.012818f
C204 VDD1.n185 B 0.012106f
C205 VDD1.n186 B 0.022529f
C206 VDD1.n187 B 0.022529f
C207 VDD1.n188 B 0.012106f
C208 VDD1.n189 B 0.012818f
C209 VDD1.n190 B 0.028615f
C210 VDD1.n191 B 0.064097f
C211 VDD1.n192 B 0.012818f
C212 VDD1.n193 B 0.012106f
C213 VDD1.n194 B 0.055769f
C214 VDD1.n195 B 0.056421f
C215 VDD1.t7 B 0.314052f
C216 VDD1.t6 B 0.314052f
C217 VDD1.n196 B 2.86097f
C218 VDD1.n197 B 0.477808f
C219 VDD1.t3 B 0.314052f
C220 VDD1.t4 B 0.314052f
C221 VDD1.n198 B 2.86773f
C222 VDD1.n199 B 2.49213f
C223 VDD1.t8 B 0.314052f
C224 VDD1.t9 B 0.314052f
C225 VDD1.n200 B 2.86097f
C226 VDD1.n201 B 2.82854f
C227 VP.n0 B 0.029774f
C228 VP.t5 B 2.13725f
C229 VP.n1 B 0.040398f
C230 VP.n2 B 0.029774f
C231 VP.t6 B 2.13725f
C232 VP.n3 B 0.054662f
C233 VP.n4 B 0.029774f
C234 VP.t3 B 2.13725f
C235 VP.n5 B 0.049098f
C236 VP.n6 B 0.029774f
C237 VP.n7 B 0.034498f
C238 VP.n8 B 0.029774f
C239 VP.t0 B 2.13725f
C240 VP.n9 B 0.040398f
C241 VP.n10 B 0.029774f
C242 VP.t1 B 2.13725f
C243 VP.n11 B 0.054662f
C244 VP.n12 B 0.029774f
C245 VP.t8 B 2.13725f
C246 VP.n13 B 0.049098f
C247 VP.t9 B 2.223f
C248 VP.t7 B 2.13725f
C249 VP.n14 B 0.811012f
C250 VP.n15 B 0.826851f
C251 VP.n16 B 0.185904f
C252 VP.n17 B 0.029774f
C253 VP.n18 B 0.027659f
C254 VP.n19 B 0.054662f
C255 VP.n20 B 0.781353f
C256 VP.n21 B 0.029774f
C257 VP.n22 B 0.029774f
C258 VP.n23 B 0.029774f
C259 VP.n24 B 0.027659f
C260 VP.n25 B 0.049098f
C261 VP.n26 B 0.753397f
C262 VP.n27 B 0.038314f
C263 VP.n28 B 0.029774f
C264 VP.n29 B 0.029774f
C265 VP.n30 B 0.029774f
C266 VP.n31 B 0.046165f
C267 VP.n32 B 0.034498f
C268 VP.n33 B 0.807763f
C269 VP.n34 B 1.68125f
C270 VP.t4 B 2.13725f
C271 VP.n35 B 0.807763f
C272 VP.n36 B 1.70223f
C273 VP.n37 B 0.029774f
C274 VP.n38 B 0.029774f
C275 VP.n39 B 0.046165f
C276 VP.n40 B 0.040398f
C277 VP.t2 B 2.13725f
C278 VP.n41 B 0.753397f
C279 VP.n42 B 0.038314f
C280 VP.n43 B 0.029774f
C281 VP.n44 B 0.029774f
C282 VP.n45 B 0.029774f
C283 VP.n46 B 0.027659f
C284 VP.n47 B 0.054662f
C285 VP.n48 B 0.781353f
C286 VP.n49 B 0.029774f
C287 VP.n50 B 0.029774f
C288 VP.n51 B 0.029774f
C289 VP.n52 B 0.027659f
C290 VP.n53 B 0.049098f
C291 VP.n54 B 0.753397f
C292 VP.n55 B 0.038314f
C293 VP.n56 B 0.029774f
C294 VP.n57 B 0.029774f
C295 VP.n58 B 0.029774f
C296 VP.n59 B 0.046165f
C297 VP.n60 B 0.034498f
C298 VP.n61 B 0.807763f
C299 VP.n62 B 0.029373f
C300 VTAIL.t18 B 0.328682f
C301 VTAIL.t11 B 0.328682f
C302 VTAIL.n0 B 2.92632f
C303 VTAIL.n1 B 0.417393f
C304 VTAIL.n2 B 0.034415f
C305 VTAIL.n3 B 0.023579f
C306 VTAIL.n4 B 0.01267f
C307 VTAIL.n5 B 0.029948f
C308 VTAIL.n6 B 0.013416f
C309 VTAIL.n7 B 0.023579f
C310 VTAIL.n8 B 0.01267f
C311 VTAIL.n9 B 0.029948f
C312 VTAIL.n10 B 0.013043f
C313 VTAIL.n11 B 0.023579f
C314 VTAIL.n12 B 0.013416f
C315 VTAIL.n13 B 0.029948f
C316 VTAIL.n14 B 0.013416f
C317 VTAIL.n15 B 0.023579f
C318 VTAIL.n16 B 0.01267f
C319 VTAIL.n17 B 0.029948f
C320 VTAIL.n18 B 0.013416f
C321 VTAIL.n19 B 0.023579f
C322 VTAIL.n20 B 0.01267f
C323 VTAIL.n21 B 0.029948f
C324 VTAIL.n22 B 0.013416f
C325 VTAIL.n23 B 0.023579f
C326 VTAIL.n24 B 0.01267f
C327 VTAIL.n25 B 0.029948f
C328 VTAIL.n26 B 0.013416f
C329 VTAIL.n27 B 0.023579f
C330 VTAIL.n28 B 0.01267f
C331 VTAIL.n29 B 0.029948f
C332 VTAIL.n30 B 0.013416f
C333 VTAIL.n31 B 1.81936f
C334 VTAIL.n32 B 0.01267f
C335 VTAIL.t2 B 0.049594f
C336 VTAIL.n33 B 0.169394f
C337 VTAIL.n34 B 0.017691f
C338 VTAIL.n35 B 0.022461f
C339 VTAIL.n36 B 0.029948f
C340 VTAIL.n37 B 0.013416f
C341 VTAIL.n38 B 0.01267f
C342 VTAIL.n39 B 0.023579f
C343 VTAIL.n40 B 0.023579f
C344 VTAIL.n41 B 0.01267f
C345 VTAIL.n42 B 0.013416f
C346 VTAIL.n43 B 0.029948f
C347 VTAIL.n44 B 0.029948f
C348 VTAIL.n45 B 0.013416f
C349 VTAIL.n46 B 0.01267f
C350 VTAIL.n47 B 0.023579f
C351 VTAIL.n48 B 0.023579f
C352 VTAIL.n49 B 0.01267f
C353 VTAIL.n50 B 0.013416f
C354 VTAIL.n51 B 0.029948f
C355 VTAIL.n52 B 0.029948f
C356 VTAIL.n53 B 0.013416f
C357 VTAIL.n54 B 0.01267f
C358 VTAIL.n55 B 0.023579f
C359 VTAIL.n56 B 0.023579f
C360 VTAIL.n57 B 0.01267f
C361 VTAIL.n58 B 0.013416f
C362 VTAIL.n59 B 0.029948f
C363 VTAIL.n60 B 0.029948f
C364 VTAIL.n61 B 0.013416f
C365 VTAIL.n62 B 0.01267f
C366 VTAIL.n63 B 0.023579f
C367 VTAIL.n64 B 0.023579f
C368 VTAIL.n65 B 0.01267f
C369 VTAIL.n66 B 0.013416f
C370 VTAIL.n67 B 0.029948f
C371 VTAIL.n68 B 0.029948f
C372 VTAIL.n69 B 0.013416f
C373 VTAIL.n70 B 0.01267f
C374 VTAIL.n71 B 0.023579f
C375 VTAIL.n72 B 0.023579f
C376 VTAIL.n73 B 0.01267f
C377 VTAIL.n74 B 0.01267f
C378 VTAIL.n75 B 0.013416f
C379 VTAIL.n76 B 0.029948f
C380 VTAIL.n77 B 0.029948f
C381 VTAIL.n78 B 0.029948f
C382 VTAIL.n79 B 0.013043f
C383 VTAIL.n80 B 0.01267f
C384 VTAIL.n81 B 0.023579f
C385 VTAIL.n82 B 0.023579f
C386 VTAIL.n83 B 0.01267f
C387 VTAIL.n84 B 0.013416f
C388 VTAIL.n85 B 0.029948f
C389 VTAIL.n86 B 0.029948f
C390 VTAIL.n87 B 0.013416f
C391 VTAIL.n88 B 0.01267f
C392 VTAIL.n89 B 0.023579f
C393 VTAIL.n90 B 0.023579f
C394 VTAIL.n91 B 0.01267f
C395 VTAIL.n92 B 0.013416f
C396 VTAIL.n93 B 0.029948f
C397 VTAIL.n94 B 0.067083f
C398 VTAIL.n95 B 0.013416f
C399 VTAIL.n96 B 0.01267f
C400 VTAIL.n97 B 0.058367f
C401 VTAIL.n98 B 0.037882f
C402 VTAIL.n99 B 0.235843f
C403 VTAIL.t0 B 0.328682f
C404 VTAIL.t3 B 0.328682f
C405 VTAIL.n100 B 2.92632f
C406 VTAIL.n101 B 0.466189f
C407 VTAIL.t5 B 0.328682f
C408 VTAIL.t4 B 0.328682f
C409 VTAIL.n102 B 2.92632f
C410 VTAIL.n103 B 2.0604f
C411 VTAIL.t10 B 0.328682f
C412 VTAIL.t19 B 0.328682f
C413 VTAIL.n104 B 2.92633f
C414 VTAIL.n105 B 2.06038f
C415 VTAIL.t13 B 0.328682f
C416 VTAIL.t12 B 0.328682f
C417 VTAIL.n106 B 2.92633f
C418 VTAIL.n107 B 0.466176f
C419 VTAIL.n108 B 0.034415f
C420 VTAIL.n109 B 0.023579f
C421 VTAIL.n110 B 0.01267f
C422 VTAIL.n111 B 0.029948f
C423 VTAIL.n112 B 0.013416f
C424 VTAIL.n113 B 0.023579f
C425 VTAIL.n114 B 0.01267f
C426 VTAIL.n115 B 0.029948f
C427 VTAIL.n116 B 0.013043f
C428 VTAIL.n117 B 0.023579f
C429 VTAIL.n118 B 0.013043f
C430 VTAIL.n119 B 0.01267f
C431 VTAIL.n120 B 0.029948f
C432 VTAIL.n121 B 0.029948f
C433 VTAIL.n122 B 0.013416f
C434 VTAIL.n123 B 0.023579f
C435 VTAIL.n124 B 0.01267f
C436 VTAIL.n125 B 0.029948f
C437 VTAIL.n126 B 0.013416f
C438 VTAIL.n127 B 0.023579f
C439 VTAIL.n128 B 0.01267f
C440 VTAIL.n129 B 0.029948f
C441 VTAIL.n130 B 0.013416f
C442 VTAIL.n131 B 0.023579f
C443 VTAIL.n132 B 0.01267f
C444 VTAIL.n133 B 0.029948f
C445 VTAIL.n134 B 0.013416f
C446 VTAIL.n135 B 0.023579f
C447 VTAIL.n136 B 0.01267f
C448 VTAIL.n137 B 0.029948f
C449 VTAIL.n138 B 0.013416f
C450 VTAIL.n139 B 1.81936f
C451 VTAIL.n140 B 0.01267f
C452 VTAIL.t14 B 0.049594f
C453 VTAIL.n141 B 0.169394f
C454 VTAIL.n142 B 0.017691f
C455 VTAIL.n143 B 0.022461f
C456 VTAIL.n144 B 0.029948f
C457 VTAIL.n145 B 0.013416f
C458 VTAIL.n146 B 0.01267f
C459 VTAIL.n147 B 0.023579f
C460 VTAIL.n148 B 0.023579f
C461 VTAIL.n149 B 0.01267f
C462 VTAIL.n150 B 0.013416f
C463 VTAIL.n151 B 0.029948f
C464 VTAIL.n152 B 0.029948f
C465 VTAIL.n153 B 0.013416f
C466 VTAIL.n154 B 0.01267f
C467 VTAIL.n155 B 0.023579f
C468 VTAIL.n156 B 0.023579f
C469 VTAIL.n157 B 0.01267f
C470 VTAIL.n158 B 0.013416f
C471 VTAIL.n159 B 0.029948f
C472 VTAIL.n160 B 0.029948f
C473 VTAIL.n161 B 0.013416f
C474 VTAIL.n162 B 0.01267f
C475 VTAIL.n163 B 0.023579f
C476 VTAIL.n164 B 0.023579f
C477 VTAIL.n165 B 0.01267f
C478 VTAIL.n166 B 0.013416f
C479 VTAIL.n167 B 0.029948f
C480 VTAIL.n168 B 0.029948f
C481 VTAIL.n169 B 0.013416f
C482 VTAIL.n170 B 0.01267f
C483 VTAIL.n171 B 0.023579f
C484 VTAIL.n172 B 0.023579f
C485 VTAIL.n173 B 0.01267f
C486 VTAIL.n174 B 0.013416f
C487 VTAIL.n175 B 0.029948f
C488 VTAIL.n176 B 0.029948f
C489 VTAIL.n177 B 0.013416f
C490 VTAIL.n178 B 0.01267f
C491 VTAIL.n179 B 0.023579f
C492 VTAIL.n180 B 0.023579f
C493 VTAIL.n181 B 0.01267f
C494 VTAIL.n182 B 0.013416f
C495 VTAIL.n183 B 0.029948f
C496 VTAIL.n184 B 0.029948f
C497 VTAIL.n185 B 0.013416f
C498 VTAIL.n186 B 0.01267f
C499 VTAIL.n187 B 0.023579f
C500 VTAIL.n188 B 0.023579f
C501 VTAIL.n189 B 0.01267f
C502 VTAIL.n190 B 0.013416f
C503 VTAIL.n191 B 0.029948f
C504 VTAIL.n192 B 0.029948f
C505 VTAIL.n193 B 0.013416f
C506 VTAIL.n194 B 0.01267f
C507 VTAIL.n195 B 0.023579f
C508 VTAIL.n196 B 0.023579f
C509 VTAIL.n197 B 0.01267f
C510 VTAIL.n198 B 0.013416f
C511 VTAIL.n199 B 0.029948f
C512 VTAIL.n200 B 0.067083f
C513 VTAIL.n201 B 0.013416f
C514 VTAIL.n202 B 0.01267f
C515 VTAIL.n203 B 0.058367f
C516 VTAIL.n204 B 0.037882f
C517 VTAIL.n205 B 0.235843f
C518 VTAIL.t7 B 0.328682f
C519 VTAIL.t1 B 0.328682f
C520 VTAIL.n206 B 2.92633f
C521 VTAIL.n207 B 0.442597f
C522 VTAIL.t6 B 0.328682f
C523 VTAIL.t9 B 0.328682f
C524 VTAIL.n208 B 2.92633f
C525 VTAIL.n209 B 0.466176f
C526 VTAIL.n210 B 0.034415f
C527 VTAIL.n211 B 0.023579f
C528 VTAIL.n212 B 0.01267f
C529 VTAIL.n213 B 0.029948f
C530 VTAIL.n214 B 0.013416f
C531 VTAIL.n215 B 0.023579f
C532 VTAIL.n216 B 0.01267f
C533 VTAIL.n217 B 0.029948f
C534 VTAIL.n218 B 0.013043f
C535 VTAIL.n219 B 0.023579f
C536 VTAIL.n220 B 0.013043f
C537 VTAIL.n221 B 0.01267f
C538 VTAIL.n222 B 0.029948f
C539 VTAIL.n223 B 0.029948f
C540 VTAIL.n224 B 0.013416f
C541 VTAIL.n225 B 0.023579f
C542 VTAIL.n226 B 0.01267f
C543 VTAIL.n227 B 0.029948f
C544 VTAIL.n228 B 0.013416f
C545 VTAIL.n229 B 0.023579f
C546 VTAIL.n230 B 0.01267f
C547 VTAIL.n231 B 0.029948f
C548 VTAIL.n232 B 0.013416f
C549 VTAIL.n233 B 0.023579f
C550 VTAIL.n234 B 0.01267f
C551 VTAIL.n235 B 0.029948f
C552 VTAIL.n236 B 0.013416f
C553 VTAIL.n237 B 0.023579f
C554 VTAIL.n238 B 0.01267f
C555 VTAIL.n239 B 0.029948f
C556 VTAIL.n240 B 0.013416f
C557 VTAIL.n241 B 1.81936f
C558 VTAIL.n242 B 0.01267f
C559 VTAIL.t8 B 0.049594f
C560 VTAIL.n243 B 0.169394f
C561 VTAIL.n244 B 0.017691f
C562 VTAIL.n245 B 0.022461f
C563 VTAIL.n246 B 0.029948f
C564 VTAIL.n247 B 0.013416f
C565 VTAIL.n248 B 0.01267f
C566 VTAIL.n249 B 0.023579f
C567 VTAIL.n250 B 0.023579f
C568 VTAIL.n251 B 0.01267f
C569 VTAIL.n252 B 0.013416f
C570 VTAIL.n253 B 0.029948f
C571 VTAIL.n254 B 0.029948f
C572 VTAIL.n255 B 0.013416f
C573 VTAIL.n256 B 0.01267f
C574 VTAIL.n257 B 0.023579f
C575 VTAIL.n258 B 0.023579f
C576 VTAIL.n259 B 0.01267f
C577 VTAIL.n260 B 0.013416f
C578 VTAIL.n261 B 0.029948f
C579 VTAIL.n262 B 0.029948f
C580 VTAIL.n263 B 0.013416f
C581 VTAIL.n264 B 0.01267f
C582 VTAIL.n265 B 0.023579f
C583 VTAIL.n266 B 0.023579f
C584 VTAIL.n267 B 0.01267f
C585 VTAIL.n268 B 0.013416f
C586 VTAIL.n269 B 0.029948f
C587 VTAIL.n270 B 0.029948f
C588 VTAIL.n271 B 0.013416f
C589 VTAIL.n272 B 0.01267f
C590 VTAIL.n273 B 0.023579f
C591 VTAIL.n274 B 0.023579f
C592 VTAIL.n275 B 0.01267f
C593 VTAIL.n276 B 0.013416f
C594 VTAIL.n277 B 0.029948f
C595 VTAIL.n278 B 0.029948f
C596 VTAIL.n279 B 0.013416f
C597 VTAIL.n280 B 0.01267f
C598 VTAIL.n281 B 0.023579f
C599 VTAIL.n282 B 0.023579f
C600 VTAIL.n283 B 0.01267f
C601 VTAIL.n284 B 0.013416f
C602 VTAIL.n285 B 0.029948f
C603 VTAIL.n286 B 0.029948f
C604 VTAIL.n287 B 0.013416f
C605 VTAIL.n288 B 0.01267f
C606 VTAIL.n289 B 0.023579f
C607 VTAIL.n290 B 0.023579f
C608 VTAIL.n291 B 0.01267f
C609 VTAIL.n292 B 0.013416f
C610 VTAIL.n293 B 0.029948f
C611 VTAIL.n294 B 0.029948f
C612 VTAIL.n295 B 0.013416f
C613 VTAIL.n296 B 0.01267f
C614 VTAIL.n297 B 0.023579f
C615 VTAIL.n298 B 0.023579f
C616 VTAIL.n299 B 0.01267f
C617 VTAIL.n300 B 0.013416f
C618 VTAIL.n301 B 0.029948f
C619 VTAIL.n302 B 0.067083f
C620 VTAIL.n303 B 0.013416f
C621 VTAIL.n304 B 0.01267f
C622 VTAIL.n305 B 0.058367f
C623 VTAIL.n306 B 0.037882f
C624 VTAIL.n307 B 1.73508f
C625 VTAIL.n308 B 0.034415f
C626 VTAIL.n309 B 0.023579f
C627 VTAIL.n310 B 0.01267f
C628 VTAIL.n311 B 0.029948f
C629 VTAIL.n312 B 0.013416f
C630 VTAIL.n313 B 0.023579f
C631 VTAIL.n314 B 0.01267f
C632 VTAIL.n315 B 0.029948f
C633 VTAIL.n316 B 0.013043f
C634 VTAIL.n317 B 0.023579f
C635 VTAIL.n318 B 0.013416f
C636 VTAIL.n319 B 0.029948f
C637 VTAIL.n320 B 0.013416f
C638 VTAIL.n321 B 0.023579f
C639 VTAIL.n322 B 0.01267f
C640 VTAIL.n323 B 0.029948f
C641 VTAIL.n324 B 0.013416f
C642 VTAIL.n325 B 0.023579f
C643 VTAIL.n326 B 0.01267f
C644 VTAIL.n327 B 0.029948f
C645 VTAIL.n328 B 0.013416f
C646 VTAIL.n329 B 0.023579f
C647 VTAIL.n330 B 0.01267f
C648 VTAIL.n331 B 0.029948f
C649 VTAIL.n332 B 0.013416f
C650 VTAIL.n333 B 0.023579f
C651 VTAIL.n334 B 0.01267f
C652 VTAIL.n335 B 0.029948f
C653 VTAIL.n336 B 0.013416f
C654 VTAIL.n337 B 1.81936f
C655 VTAIL.n338 B 0.01267f
C656 VTAIL.t17 B 0.049594f
C657 VTAIL.n339 B 0.169394f
C658 VTAIL.n340 B 0.017691f
C659 VTAIL.n341 B 0.022461f
C660 VTAIL.n342 B 0.029948f
C661 VTAIL.n343 B 0.013416f
C662 VTAIL.n344 B 0.01267f
C663 VTAIL.n345 B 0.023579f
C664 VTAIL.n346 B 0.023579f
C665 VTAIL.n347 B 0.01267f
C666 VTAIL.n348 B 0.013416f
C667 VTAIL.n349 B 0.029948f
C668 VTAIL.n350 B 0.029948f
C669 VTAIL.n351 B 0.013416f
C670 VTAIL.n352 B 0.01267f
C671 VTAIL.n353 B 0.023579f
C672 VTAIL.n354 B 0.023579f
C673 VTAIL.n355 B 0.01267f
C674 VTAIL.n356 B 0.013416f
C675 VTAIL.n357 B 0.029948f
C676 VTAIL.n358 B 0.029948f
C677 VTAIL.n359 B 0.013416f
C678 VTAIL.n360 B 0.01267f
C679 VTAIL.n361 B 0.023579f
C680 VTAIL.n362 B 0.023579f
C681 VTAIL.n363 B 0.01267f
C682 VTAIL.n364 B 0.013416f
C683 VTAIL.n365 B 0.029948f
C684 VTAIL.n366 B 0.029948f
C685 VTAIL.n367 B 0.013416f
C686 VTAIL.n368 B 0.01267f
C687 VTAIL.n369 B 0.023579f
C688 VTAIL.n370 B 0.023579f
C689 VTAIL.n371 B 0.01267f
C690 VTAIL.n372 B 0.013416f
C691 VTAIL.n373 B 0.029948f
C692 VTAIL.n374 B 0.029948f
C693 VTAIL.n375 B 0.013416f
C694 VTAIL.n376 B 0.01267f
C695 VTAIL.n377 B 0.023579f
C696 VTAIL.n378 B 0.023579f
C697 VTAIL.n379 B 0.01267f
C698 VTAIL.n380 B 0.01267f
C699 VTAIL.n381 B 0.013416f
C700 VTAIL.n382 B 0.029948f
C701 VTAIL.n383 B 0.029948f
C702 VTAIL.n384 B 0.029948f
C703 VTAIL.n385 B 0.013043f
C704 VTAIL.n386 B 0.01267f
C705 VTAIL.n387 B 0.023579f
C706 VTAIL.n388 B 0.023579f
C707 VTAIL.n389 B 0.01267f
C708 VTAIL.n390 B 0.013416f
C709 VTAIL.n391 B 0.029948f
C710 VTAIL.n392 B 0.029948f
C711 VTAIL.n393 B 0.013416f
C712 VTAIL.n394 B 0.01267f
C713 VTAIL.n395 B 0.023579f
C714 VTAIL.n396 B 0.023579f
C715 VTAIL.n397 B 0.01267f
C716 VTAIL.n398 B 0.013416f
C717 VTAIL.n399 B 0.029948f
C718 VTAIL.n400 B 0.067083f
C719 VTAIL.n401 B 0.013416f
C720 VTAIL.n402 B 0.01267f
C721 VTAIL.n403 B 0.058367f
C722 VTAIL.n404 B 0.037882f
C723 VTAIL.n405 B 1.73508f
C724 VTAIL.t16 B 0.328682f
C725 VTAIL.t15 B 0.328682f
C726 VTAIL.n406 B 2.92632f
C727 VTAIL.n407 B 0.372855f
C728 VDD2.n0 B 0.032629f
C729 VDD2.n1 B 0.022355f
C730 VDD2.n2 B 0.012013f
C731 VDD2.n3 B 0.028394f
C732 VDD2.n4 B 0.012719f
C733 VDD2.n5 B 0.022355f
C734 VDD2.n6 B 0.012013f
C735 VDD2.n7 B 0.028394f
C736 VDD2.n8 B 0.012366f
C737 VDD2.n9 B 0.022355f
C738 VDD2.n10 B 0.012719f
C739 VDD2.n11 B 0.028394f
C740 VDD2.n12 B 0.012719f
C741 VDD2.n13 B 0.022355f
C742 VDD2.n14 B 0.012013f
C743 VDD2.n15 B 0.028394f
C744 VDD2.n16 B 0.012719f
C745 VDD2.n17 B 0.022355f
C746 VDD2.n18 B 0.012013f
C747 VDD2.n19 B 0.028394f
C748 VDD2.n20 B 0.012719f
C749 VDD2.n21 B 0.022355f
C750 VDD2.n22 B 0.012013f
C751 VDD2.n23 B 0.028394f
C752 VDD2.n24 B 0.012719f
C753 VDD2.n25 B 0.022355f
C754 VDD2.n26 B 0.012013f
C755 VDD2.n27 B 0.028394f
C756 VDD2.n28 B 0.012719f
C757 VDD2.n29 B 1.72493f
C758 VDD2.n30 B 0.012013f
C759 VDD2.t2 B 0.04702f
C760 VDD2.n31 B 0.160601f
C761 VDD2.n32 B 0.016773f
C762 VDD2.n33 B 0.021295f
C763 VDD2.n34 B 0.028394f
C764 VDD2.n35 B 0.012719f
C765 VDD2.n36 B 0.012013f
C766 VDD2.n37 B 0.022355f
C767 VDD2.n38 B 0.022355f
C768 VDD2.n39 B 0.012013f
C769 VDD2.n40 B 0.012719f
C770 VDD2.n41 B 0.028394f
C771 VDD2.n42 B 0.028394f
C772 VDD2.n43 B 0.012719f
C773 VDD2.n44 B 0.012013f
C774 VDD2.n45 B 0.022355f
C775 VDD2.n46 B 0.022355f
C776 VDD2.n47 B 0.012013f
C777 VDD2.n48 B 0.012719f
C778 VDD2.n49 B 0.028394f
C779 VDD2.n50 B 0.028394f
C780 VDD2.n51 B 0.012719f
C781 VDD2.n52 B 0.012013f
C782 VDD2.n53 B 0.022355f
C783 VDD2.n54 B 0.022355f
C784 VDD2.n55 B 0.012013f
C785 VDD2.n56 B 0.012719f
C786 VDD2.n57 B 0.028394f
C787 VDD2.n58 B 0.028394f
C788 VDD2.n59 B 0.012719f
C789 VDD2.n60 B 0.012013f
C790 VDD2.n61 B 0.022355f
C791 VDD2.n62 B 0.022355f
C792 VDD2.n63 B 0.012013f
C793 VDD2.n64 B 0.012719f
C794 VDD2.n65 B 0.028394f
C795 VDD2.n66 B 0.028394f
C796 VDD2.n67 B 0.012719f
C797 VDD2.n68 B 0.012013f
C798 VDD2.n69 B 0.022355f
C799 VDD2.n70 B 0.022355f
C800 VDD2.n71 B 0.012013f
C801 VDD2.n72 B 0.012013f
C802 VDD2.n73 B 0.012719f
C803 VDD2.n74 B 0.028394f
C804 VDD2.n75 B 0.028394f
C805 VDD2.n76 B 0.028394f
C806 VDD2.n77 B 0.012366f
C807 VDD2.n78 B 0.012013f
C808 VDD2.n79 B 0.022355f
C809 VDD2.n80 B 0.022355f
C810 VDD2.n81 B 0.012013f
C811 VDD2.n82 B 0.012719f
C812 VDD2.n83 B 0.028394f
C813 VDD2.n84 B 0.028394f
C814 VDD2.n85 B 0.012719f
C815 VDD2.n86 B 0.012013f
C816 VDD2.n87 B 0.022355f
C817 VDD2.n88 B 0.022355f
C818 VDD2.n89 B 0.012013f
C819 VDD2.n90 B 0.012719f
C820 VDD2.n91 B 0.028394f
C821 VDD2.n92 B 0.063601f
C822 VDD2.n93 B 0.012719f
C823 VDD2.n94 B 0.012013f
C824 VDD2.n95 B 0.055337f
C825 VDD2.n96 B 0.055985f
C826 VDD2.t5 B 0.311622f
C827 VDD2.t6 B 0.311622f
C828 VDD2.n97 B 2.83884f
C829 VDD2.n98 B 0.474111f
C830 VDD2.t9 B 0.311622f
C831 VDD2.t7 B 0.311622f
C832 VDD2.n99 B 2.84554f
C833 VDD2.n100 B 2.38489f
C834 VDD2.n101 B 0.032629f
C835 VDD2.n102 B 0.022355f
C836 VDD2.n103 B 0.012013f
C837 VDD2.n104 B 0.028394f
C838 VDD2.n105 B 0.012719f
C839 VDD2.n106 B 0.022355f
C840 VDD2.n107 B 0.012013f
C841 VDD2.n108 B 0.028394f
C842 VDD2.n109 B 0.012366f
C843 VDD2.n110 B 0.022355f
C844 VDD2.n111 B 0.012366f
C845 VDD2.n112 B 0.012013f
C846 VDD2.n113 B 0.028394f
C847 VDD2.n114 B 0.028394f
C848 VDD2.n115 B 0.012719f
C849 VDD2.n116 B 0.022355f
C850 VDD2.n117 B 0.012013f
C851 VDD2.n118 B 0.028394f
C852 VDD2.n119 B 0.012719f
C853 VDD2.n120 B 0.022355f
C854 VDD2.n121 B 0.012013f
C855 VDD2.n122 B 0.028394f
C856 VDD2.n123 B 0.012719f
C857 VDD2.n124 B 0.022355f
C858 VDD2.n125 B 0.012013f
C859 VDD2.n126 B 0.028394f
C860 VDD2.n127 B 0.012719f
C861 VDD2.n128 B 0.022355f
C862 VDD2.n129 B 0.012013f
C863 VDD2.n130 B 0.028394f
C864 VDD2.n131 B 0.012719f
C865 VDD2.n132 B 1.72493f
C866 VDD2.n133 B 0.012013f
C867 VDD2.t4 B 0.04702f
C868 VDD2.n134 B 0.160601f
C869 VDD2.n135 B 0.016773f
C870 VDD2.n136 B 0.021295f
C871 VDD2.n137 B 0.028394f
C872 VDD2.n138 B 0.012719f
C873 VDD2.n139 B 0.012013f
C874 VDD2.n140 B 0.022355f
C875 VDD2.n141 B 0.022355f
C876 VDD2.n142 B 0.012013f
C877 VDD2.n143 B 0.012719f
C878 VDD2.n144 B 0.028394f
C879 VDD2.n145 B 0.028394f
C880 VDD2.n146 B 0.012719f
C881 VDD2.n147 B 0.012013f
C882 VDD2.n148 B 0.022355f
C883 VDD2.n149 B 0.022355f
C884 VDD2.n150 B 0.012013f
C885 VDD2.n151 B 0.012719f
C886 VDD2.n152 B 0.028394f
C887 VDD2.n153 B 0.028394f
C888 VDD2.n154 B 0.012719f
C889 VDD2.n155 B 0.012013f
C890 VDD2.n156 B 0.022355f
C891 VDD2.n157 B 0.022355f
C892 VDD2.n158 B 0.012013f
C893 VDD2.n159 B 0.012719f
C894 VDD2.n160 B 0.028394f
C895 VDD2.n161 B 0.028394f
C896 VDD2.n162 B 0.012719f
C897 VDD2.n163 B 0.012013f
C898 VDD2.n164 B 0.022355f
C899 VDD2.n165 B 0.022355f
C900 VDD2.n166 B 0.012013f
C901 VDD2.n167 B 0.012719f
C902 VDD2.n168 B 0.028394f
C903 VDD2.n169 B 0.028394f
C904 VDD2.n170 B 0.012719f
C905 VDD2.n171 B 0.012013f
C906 VDD2.n172 B 0.022355f
C907 VDD2.n173 B 0.022355f
C908 VDD2.n174 B 0.012013f
C909 VDD2.n175 B 0.012719f
C910 VDD2.n176 B 0.028394f
C911 VDD2.n177 B 0.028394f
C912 VDD2.n178 B 0.012719f
C913 VDD2.n179 B 0.012013f
C914 VDD2.n180 B 0.022355f
C915 VDD2.n181 B 0.022355f
C916 VDD2.n182 B 0.012013f
C917 VDD2.n183 B 0.012719f
C918 VDD2.n184 B 0.028394f
C919 VDD2.n185 B 0.028394f
C920 VDD2.n186 B 0.012719f
C921 VDD2.n187 B 0.012013f
C922 VDD2.n188 B 0.022355f
C923 VDD2.n189 B 0.022355f
C924 VDD2.n190 B 0.012013f
C925 VDD2.n191 B 0.012719f
C926 VDD2.n192 B 0.028394f
C927 VDD2.n193 B 0.063601f
C928 VDD2.n194 B 0.012719f
C929 VDD2.n195 B 0.012013f
C930 VDD2.n196 B 0.055337f
C931 VDD2.n197 B 0.051325f
C932 VDD2.n198 B 2.5849f
C933 VDD2.t3 B 0.311622f
C934 VDD2.t1 B 0.311622f
C935 VDD2.n199 B 2.83884f
C936 VDD2.n200 B 0.327851f
C937 VDD2.t0 B 0.311622f
C938 VDD2.t8 B 0.311622f
C939 VDD2.n201 B 2.84551f
C940 VN.n0 B 0.029481f
C941 VN.t2 B 2.11622f
C942 VN.n1 B 0.040001f
C943 VN.n2 B 0.029481f
C944 VN.t4 B 2.11622f
C945 VN.n3 B 0.054124f
C946 VN.n4 B 0.029481f
C947 VN.t3 B 2.11622f
C948 VN.n5 B 0.048615f
C949 VN.t1 B 2.20113f
C950 VN.t8 B 2.11622f
C951 VN.n6 B 0.803032f
C952 VN.n7 B 0.818715f
C953 VN.n8 B 0.184075f
C954 VN.n9 B 0.029481f
C955 VN.n10 B 0.027387f
C956 VN.n11 B 0.054124f
C957 VN.n12 B 0.773665f
C958 VN.n13 B 0.029481f
C959 VN.n14 B 0.029481f
C960 VN.n15 B 0.029481f
C961 VN.n16 B 0.027387f
C962 VN.n17 B 0.048615f
C963 VN.n18 B 0.745984f
C964 VN.n19 B 0.037937f
C965 VN.n20 B 0.029481f
C966 VN.n21 B 0.029481f
C967 VN.n22 B 0.029481f
C968 VN.n23 B 0.04571f
C969 VN.n24 B 0.034158f
C970 VN.n25 B 0.799814f
C971 VN.n26 B 0.029084f
C972 VN.n27 B 0.029481f
C973 VN.t9 B 2.11622f
C974 VN.n28 B 0.040001f
C975 VN.n29 B 0.029481f
C976 VN.t0 B 2.11622f
C977 VN.n30 B 0.054124f
C978 VN.n31 B 0.029481f
C979 VN.t6 B 2.11622f
C980 VN.n32 B 0.048615f
C981 VN.t5 B 2.20113f
C982 VN.t7 B 2.11622f
C983 VN.n33 B 0.803032f
C984 VN.n34 B 0.818715f
C985 VN.n35 B 0.184075f
C986 VN.n36 B 0.029481f
C987 VN.n37 B 0.027387f
C988 VN.n38 B 0.054124f
C989 VN.n39 B 0.773665f
C990 VN.n40 B 0.029481f
C991 VN.n41 B 0.029481f
C992 VN.n42 B 0.029481f
C993 VN.n43 B 0.027387f
C994 VN.n44 B 0.048615f
C995 VN.n45 B 0.745984f
C996 VN.n46 B 0.037937f
C997 VN.n47 B 0.029481f
C998 VN.n48 B 0.029481f
C999 VN.n49 B 0.029481f
C1000 VN.n50 B 0.04571f
C1001 VN.n51 B 0.034158f
C1002 VN.n52 B 0.799814f
C1003 VN.n53 B 1.68385f
.ends

