* NGSPICE file created from diff_pair_sample_1445.ext - technology: sky130A

.subckt diff_pair_sample_1445 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t7 VN.t0 VDD2.t0 B.t3 sky130_fd_pr__nfet_01v8 ad=0.7332 pd=4.54 as=0.3102 ps=2.21 w=1.88 l=3.06
X1 B.t17 B.t15 B.t16 B.t9 sky130_fd_pr__nfet_01v8 ad=0.7332 pd=4.54 as=0 ps=0 w=1.88 l=3.06
X2 VDD1.t3 VP.t0 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=0.3102 pd=2.21 as=0.7332 ps=4.54 w=1.88 l=3.06
X3 B.t14 B.t12 B.t13 B.t5 sky130_fd_pr__nfet_01v8 ad=0.7332 pd=4.54 as=0 ps=0 w=1.88 l=3.06
X4 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=0.7332 pd=4.54 as=0 ps=0 w=1.88 l=3.06
X5 B.t7 B.t4 B.t6 B.t5 sky130_fd_pr__nfet_01v8 ad=0.7332 pd=4.54 as=0 ps=0 w=1.88 l=3.06
X6 VDD2.t1 VN.t1 VTAIL.t6 B.t0 sky130_fd_pr__nfet_01v8 ad=0.3102 pd=2.21 as=0.7332 ps=4.54 w=1.88 l=3.06
X7 VTAIL.t2 VP.t1 VDD1.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=0.7332 pd=4.54 as=0.3102 ps=2.21 w=1.88 l=3.06
X8 VDD2.t3 VN.t2 VTAIL.t5 B.t1 sky130_fd_pr__nfet_01v8 ad=0.3102 pd=2.21 as=0.7332 ps=4.54 w=1.88 l=3.06
X9 VTAIL.t4 VN.t3 VDD2.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=0.7332 pd=4.54 as=0.3102 ps=2.21 w=1.88 l=3.06
X10 VDD1.t1 VP.t2 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=0.3102 pd=2.21 as=0.7332 ps=4.54 w=1.88 l=3.06
X11 VTAIL.t3 VP.t3 VDD1.t0 B.t3 sky130_fd_pr__nfet_01v8 ad=0.7332 pd=4.54 as=0.3102 ps=2.21 w=1.88 l=3.06
R0 VN.n1 VN.t2 49.3753
R1 VN.n0 VN.t0 49.3753
R2 VN.n0 VN.t1 48.3688
R3 VN.n1 VN.t3 48.3688
R4 VN VN.n1 43.1976
R5 VN VN.n0 2.89075
R6 VDD2.n2 VDD2.n0 137.465
R7 VDD2.n2 VDD2.n1 103.362
R8 VDD2.n1 VDD2.t2 10.5324
R9 VDD2.n1 VDD2.t3 10.5324
R10 VDD2.n0 VDD2.t0 10.5324
R11 VDD2.n0 VDD2.t1 10.5324
R12 VDD2 VDD2.n2 0.0586897
R13 VTAIL.n58 VTAIL.n56 289.615
R14 VTAIL.n2 VTAIL.n0 289.615
R15 VTAIL.n10 VTAIL.n8 289.615
R16 VTAIL.n18 VTAIL.n16 289.615
R17 VTAIL.n50 VTAIL.n48 289.615
R18 VTAIL.n42 VTAIL.n40 289.615
R19 VTAIL.n34 VTAIL.n32 289.615
R20 VTAIL.n26 VTAIL.n24 289.615
R21 VTAIL.n59 VTAIL.n58 185
R22 VTAIL.n3 VTAIL.n2 185
R23 VTAIL.n11 VTAIL.n10 185
R24 VTAIL.n19 VTAIL.n18 185
R25 VTAIL.n51 VTAIL.n50 185
R26 VTAIL.n43 VTAIL.n42 185
R27 VTAIL.n35 VTAIL.n34 185
R28 VTAIL.n27 VTAIL.n26 185
R29 VTAIL.t6 VTAIL.n57 164.876
R30 VTAIL.t7 VTAIL.n1 164.876
R31 VTAIL.t1 VTAIL.n9 164.876
R32 VTAIL.t2 VTAIL.n17 164.876
R33 VTAIL.t0 VTAIL.n49 164.876
R34 VTAIL.t3 VTAIL.n41 164.876
R35 VTAIL.t5 VTAIL.n33 164.876
R36 VTAIL.t4 VTAIL.n25 164.876
R37 VTAIL.n58 VTAIL.t6 52.3082
R38 VTAIL.n2 VTAIL.t7 52.3082
R39 VTAIL.n10 VTAIL.t1 52.3082
R40 VTAIL.n18 VTAIL.t2 52.3082
R41 VTAIL.n50 VTAIL.t0 52.3082
R42 VTAIL.n42 VTAIL.t3 52.3082
R43 VTAIL.n34 VTAIL.t5 52.3082
R44 VTAIL.n26 VTAIL.t4 52.3082
R45 VTAIL.n63 VTAIL.n62 36.0641
R46 VTAIL.n7 VTAIL.n6 36.0641
R47 VTAIL.n15 VTAIL.n14 36.0641
R48 VTAIL.n23 VTAIL.n22 36.0641
R49 VTAIL.n55 VTAIL.n54 36.0641
R50 VTAIL.n47 VTAIL.n46 36.0641
R51 VTAIL.n39 VTAIL.n38 36.0641
R52 VTAIL.n31 VTAIL.n30 36.0641
R53 VTAIL.n63 VTAIL.n55 16.91
R54 VTAIL.n31 VTAIL.n23 16.91
R55 VTAIL.n59 VTAIL.n57 14.7318
R56 VTAIL.n3 VTAIL.n1 14.7318
R57 VTAIL.n11 VTAIL.n9 14.7318
R58 VTAIL.n19 VTAIL.n17 14.7318
R59 VTAIL.n51 VTAIL.n49 14.7318
R60 VTAIL.n43 VTAIL.n41 14.7318
R61 VTAIL.n35 VTAIL.n33 14.7318
R62 VTAIL.n27 VTAIL.n25 14.7318
R63 VTAIL.n60 VTAIL.n56 12.8005
R64 VTAIL.n4 VTAIL.n0 12.8005
R65 VTAIL.n12 VTAIL.n8 12.8005
R66 VTAIL.n20 VTAIL.n16 12.8005
R67 VTAIL.n52 VTAIL.n48 12.8005
R68 VTAIL.n44 VTAIL.n40 12.8005
R69 VTAIL.n36 VTAIL.n32 12.8005
R70 VTAIL.n28 VTAIL.n24 12.8005
R71 VTAIL.n62 VTAIL.n61 9.45567
R72 VTAIL.n6 VTAIL.n5 9.45567
R73 VTAIL.n14 VTAIL.n13 9.45567
R74 VTAIL.n22 VTAIL.n21 9.45567
R75 VTAIL.n54 VTAIL.n53 9.45567
R76 VTAIL.n46 VTAIL.n45 9.45567
R77 VTAIL.n38 VTAIL.n37 9.45567
R78 VTAIL.n30 VTAIL.n29 9.45567
R79 VTAIL.n61 VTAIL.n60 9.3005
R80 VTAIL.n5 VTAIL.n4 9.3005
R81 VTAIL.n13 VTAIL.n12 9.3005
R82 VTAIL.n21 VTAIL.n20 9.3005
R83 VTAIL.n53 VTAIL.n52 9.3005
R84 VTAIL.n45 VTAIL.n44 9.3005
R85 VTAIL.n37 VTAIL.n36 9.3005
R86 VTAIL.n29 VTAIL.n28 9.3005
R87 VTAIL.n61 VTAIL.n57 5.62509
R88 VTAIL.n5 VTAIL.n1 5.62509
R89 VTAIL.n13 VTAIL.n9 5.62509
R90 VTAIL.n21 VTAIL.n17 5.62509
R91 VTAIL.n53 VTAIL.n49 5.62509
R92 VTAIL.n45 VTAIL.n41 5.62509
R93 VTAIL.n37 VTAIL.n33 5.62509
R94 VTAIL.n29 VTAIL.n25 5.62509
R95 VTAIL.n39 VTAIL.n31 2.92291
R96 VTAIL.n55 VTAIL.n47 2.92291
R97 VTAIL.n23 VTAIL.n15 2.92291
R98 VTAIL VTAIL.n7 1.5199
R99 VTAIL VTAIL.n63 1.40352
R100 VTAIL.n62 VTAIL.n56 1.16414
R101 VTAIL.n6 VTAIL.n0 1.16414
R102 VTAIL.n14 VTAIL.n8 1.16414
R103 VTAIL.n22 VTAIL.n16 1.16414
R104 VTAIL.n54 VTAIL.n48 1.16414
R105 VTAIL.n46 VTAIL.n40 1.16414
R106 VTAIL.n38 VTAIL.n32 1.16414
R107 VTAIL.n30 VTAIL.n24 1.16414
R108 VTAIL.n47 VTAIL.n39 0.470328
R109 VTAIL.n15 VTAIL.n7 0.470328
R110 VTAIL.n60 VTAIL.n59 0.388379
R111 VTAIL.n4 VTAIL.n3 0.388379
R112 VTAIL.n12 VTAIL.n11 0.388379
R113 VTAIL.n20 VTAIL.n19 0.388379
R114 VTAIL.n52 VTAIL.n51 0.388379
R115 VTAIL.n44 VTAIL.n43 0.388379
R116 VTAIL.n36 VTAIL.n35 0.388379
R117 VTAIL.n28 VTAIL.n27 0.388379
R118 B.n417 B.n92 585
R119 B.n92 B.n71 585
R120 B.n419 B.n418 585
R121 B.n421 B.n91 585
R122 B.n424 B.n423 585
R123 B.n425 B.n90 585
R124 B.n427 B.n426 585
R125 B.n429 B.n89 585
R126 B.n432 B.n431 585
R127 B.n433 B.n88 585
R128 B.n435 B.n434 585
R129 B.n437 B.n87 585
R130 B.n440 B.n439 585
R131 B.n442 B.n84 585
R132 B.n444 B.n443 585
R133 B.n446 B.n83 585
R134 B.n449 B.n448 585
R135 B.n450 B.n82 585
R136 B.n452 B.n451 585
R137 B.n454 B.n81 585
R138 B.n457 B.n456 585
R139 B.n458 B.n78 585
R140 B.n461 B.n460 585
R141 B.n463 B.n77 585
R142 B.n466 B.n465 585
R143 B.n467 B.n76 585
R144 B.n469 B.n468 585
R145 B.n471 B.n75 585
R146 B.n474 B.n473 585
R147 B.n475 B.n74 585
R148 B.n477 B.n476 585
R149 B.n479 B.n73 585
R150 B.n482 B.n481 585
R151 B.n483 B.n72 585
R152 B.n416 B.n70 585
R153 B.n486 B.n70 585
R154 B.n415 B.n69 585
R155 B.n487 B.n69 585
R156 B.n414 B.n68 585
R157 B.n488 B.n68 585
R158 B.n413 B.n412 585
R159 B.n412 B.n64 585
R160 B.n411 B.n63 585
R161 B.n494 B.n63 585
R162 B.n410 B.n62 585
R163 B.n495 B.n62 585
R164 B.n409 B.n61 585
R165 B.n496 B.n61 585
R166 B.n408 B.n407 585
R167 B.n407 B.n57 585
R168 B.n406 B.n56 585
R169 B.n502 B.n56 585
R170 B.n405 B.n55 585
R171 B.n503 B.n55 585
R172 B.n404 B.n54 585
R173 B.n504 B.n54 585
R174 B.n403 B.n402 585
R175 B.n402 B.n50 585
R176 B.n401 B.n49 585
R177 B.n510 B.n49 585
R178 B.n400 B.n48 585
R179 B.n511 B.n48 585
R180 B.n399 B.n47 585
R181 B.n512 B.n47 585
R182 B.n398 B.n397 585
R183 B.n397 B.n43 585
R184 B.n396 B.n42 585
R185 B.n518 B.n42 585
R186 B.n395 B.n41 585
R187 B.n519 B.n41 585
R188 B.n394 B.n40 585
R189 B.n520 B.n40 585
R190 B.n393 B.n392 585
R191 B.n392 B.n36 585
R192 B.n391 B.n35 585
R193 B.n526 B.n35 585
R194 B.n390 B.n34 585
R195 B.n527 B.n34 585
R196 B.n389 B.n33 585
R197 B.n528 B.n33 585
R198 B.n388 B.n387 585
R199 B.n387 B.n29 585
R200 B.n386 B.n28 585
R201 B.n534 B.n28 585
R202 B.n385 B.n27 585
R203 B.n535 B.n27 585
R204 B.n384 B.n26 585
R205 B.n536 B.n26 585
R206 B.n383 B.n382 585
R207 B.n382 B.n22 585
R208 B.n381 B.n21 585
R209 B.n542 B.n21 585
R210 B.n380 B.n20 585
R211 B.n543 B.n20 585
R212 B.n379 B.n19 585
R213 B.n544 B.n19 585
R214 B.n378 B.n377 585
R215 B.n377 B.n18 585
R216 B.n376 B.n14 585
R217 B.n550 B.n14 585
R218 B.n375 B.n13 585
R219 B.n551 B.n13 585
R220 B.n374 B.n12 585
R221 B.n552 B.n12 585
R222 B.n373 B.n372 585
R223 B.n372 B.n8 585
R224 B.n371 B.n7 585
R225 B.n558 B.n7 585
R226 B.n370 B.n6 585
R227 B.n559 B.n6 585
R228 B.n369 B.n5 585
R229 B.n560 B.n5 585
R230 B.n368 B.n367 585
R231 B.n367 B.n4 585
R232 B.n366 B.n93 585
R233 B.n366 B.n365 585
R234 B.n356 B.n94 585
R235 B.n95 B.n94 585
R236 B.n358 B.n357 585
R237 B.n359 B.n358 585
R238 B.n355 B.n100 585
R239 B.n100 B.n99 585
R240 B.n354 B.n353 585
R241 B.n353 B.n352 585
R242 B.n102 B.n101 585
R243 B.n345 B.n102 585
R244 B.n344 B.n343 585
R245 B.n346 B.n344 585
R246 B.n342 B.n107 585
R247 B.n107 B.n106 585
R248 B.n341 B.n340 585
R249 B.n340 B.n339 585
R250 B.n109 B.n108 585
R251 B.n110 B.n109 585
R252 B.n332 B.n331 585
R253 B.n333 B.n332 585
R254 B.n330 B.n115 585
R255 B.n115 B.n114 585
R256 B.n329 B.n328 585
R257 B.n328 B.n327 585
R258 B.n117 B.n116 585
R259 B.n118 B.n117 585
R260 B.n320 B.n319 585
R261 B.n321 B.n320 585
R262 B.n318 B.n122 585
R263 B.n126 B.n122 585
R264 B.n317 B.n316 585
R265 B.n316 B.n315 585
R266 B.n124 B.n123 585
R267 B.n125 B.n124 585
R268 B.n308 B.n307 585
R269 B.n309 B.n308 585
R270 B.n306 B.n131 585
R271 B.n131 B.n130 585
R272 B.n305 B.n304 585
R273 B.n304 B.n303 585
R274 B.n133 B.n132 585
R275 B.n134 B.n133 585
R276 B.n296 B.n295 585
R277 B.n297 B.n296 585
R278 B.n294 B.n139 585
R279 B.n139 B.n138 585
R280 B.n293 B.n292 585
R281 B.n292 B.n291 585
R282 B.n141 B.n140 585
R283 B.n142 B.n141 585
R284 B.n284 B.n283 585
R285 B.n285 B.n284 585
R286 B.n282 B.n147 585
R287 B.n147 B.n146 585
R288 B.n281 B.n280 585
R289 B.n280 B.n279 585
R290 B.n149 B.n148 585
R291 B.n150 B.n149 585
R292 B.n272 B.n271 585
R293 B.n273 B.n272 585
R294 B.n270 B.n155 585
R295 B.n155 B.n154 585
R296 B.n269 B.n268 585
R297 B.n268 B.n267 585
R298 B.n157 B.n156 585
R299 B.n158 B.n157 585
R300 B.n260 B.n259 585
R301 B.n261 B.n260 585
R302 B.n258 B.n163 585
R303 B.n163 B.n162 585
R304 B.n257 B.n256 585
R305 B.n256 B.n255 585
R306 B.n252 B.n167 585
R307 B.n251 B.n250 585
R308 B.n248 B.n168 585
R309 B.n248 B.n166 585
R310 B.n247 B.n246 585
R311 B.n245 B.n244 585
R312 B.n243 B.n170 585
R313 B.n241 B.n240 585
R314 B.n239 B.n171 585
R315 B.n238 B.n237 585
R316 B.n235 B.n172 585
R317 B.n233 B.n232 585
R318 B.n231 B.n173 585
R319 B.n229 B.n228 585
R320 B.n226 B.n176 585
R321 B.n224 B.n223 585
R322 B.n222 B.n177 585
R323 B.n221 B.n220 585
R324 B.n218 B.n178 585
R325 B.n216 B.n215 585
R326 B.n214 B.n179 585
R327 B.n213 B.n212 585
R328 B.n210 B.n209 585
R329 B.n208 B.n207 585
R330 B.n206 B.n184 585
R331 B.n204 B.n203 585
R332 B.n202 B.n185 585
R333 B.n201 B.n200 585
R334 B.n198 B.n186 585
R335 B.n196 B.n195 585
R336 B.n194 B.n187 585
R337 B.n193 B.n192 585
R338 B.n190 B.n188 585
R339 B.n165 B.n164 585
R340 B.n254 B.n253 585
R341 B.n255 B.n254 585
R342 B.n161 B.n160 585
R343 B.n162 B.n161 585
R344 B.n263 B.n262 585
R345 B.n262 B.n261 585
R346 B.n264 B.n159 585
R347 B.n159 B.n158 585
R348 B.n266 B.n265 585
R349 B.n267 B.n266 585
R350 B.n153 B.n152 585
R351 B.n154 B.n153 585
R352 B.n275 B.n274 585
R353 B.n274 B.n273 585
R354 B.n276 B.n151 585
R355 B.n151 B.n150 585
R356 B.n278 B.n277 585
R357 B.n279 B.n278 585
R358 B.n145 B.n144 585
R359 B.n146 B.n145 585
R360 B.n287 B.n286 585
R361 B.n286 B.n285 585
R362 B.n288 B.n143 585
R363 B.n143 B.n142 585
R364 B.n290 B.n289 585
R365 B.n291 B.n290 585
R366 B.n137 B.n136 585
R367 B.n138 B.n137 585
R368 B.n299 B.n298 585
R369 B.n298 B.n297 585
R370 B.n300 B.n135 585
R371 B.n135 B.n134 585
R372 B.n302 B.n301 585
R373 B.n303 B.n302 585
R374 B.n129 B.n128 585
R375 B.n130 B.n129 585
R376 B.n311 B.n310 585
R377 B.n310 B.n309 585
R378 B.n312 B.n127 585
R379 B.n127 B.n125 585
R380 B.n314 B.n313 585
R381 B.n315 B.n314 585
R382 B.n121 B.n120 585
R383 B.n126 B.n121 585
R384 B.n323 B.n322 585
R385 B.n322 B.n321 585
R386 B.n324 B.n119 585
R387 B.n119 B.n118 585
R388 B.n326 B.n325 585
R389 B.n327 B.n326 585
R390 B.n113 B.n112 585
R391 B.n114 B.n113 585
R392 B.n335 B.n334 585
R393 B.n334 B.n333 585
R394 B.n336 B.n111 585
R395 B.n111 B.n110 585
R396 B.n338 B.n337 585
R397 B.n339 B.n338 585
R398 B.n105 B.n104 585
R399 B.n106 B.n105 585
R400 B.n348 B.n347 585
R401 B.n347 B.n346 585
R402 B.n349 B.n103 585
R403 B.n345 B.n103 585
R404 B.n351 B.n350 585
R405 B.n352 B.n351 585
R406 B.n98 B.n97 585
R407 B.n99 B.n98 585
R408 B.n361 B.n360 585
R409 B.n360 B.n359 585
R410 B.n362 B.n96 585
R411 B.n96 B.n95 585
R412 B.n364 B.n363 585
R413 B.n365 B.n364 585
R414 B.n2 B.n0 585
R415 B.n4 B.n2 585
R416 B.n3 B.n1 585
R417 B.n559 B.n3 585
R418 B.n557 B.n556 585
R419 B.n558 B.n557 585
R420 B.n555 B.n9 585
R421 B.n9 B.n8 585
R422 B.n554 B.n553 585
R423 B.n553 B.n552 585
R424 B.n11 B.n10 585
R425 B.n551 B.n11 585
R426 B.n549 B.n548 585
R427 B.n550 B.n549 585
R428 B.n547 B.n15 585
R429 B.n18 B.n15 585
R430 B.n546 B.n545 585
R431 B.n545 B.n544 585
R432 B.n17 B.n16 585
R433 B.n543 B.n17 585
R434 B.n541 B.n540 585
R435 B.n542 B.n541 585
R436 B.n539 B.n23 585
R437 B.n23 B.n22 585
R438 B.n538 B.n537 585
R439 B.n537 B.n536 585
R440 B.n25 B.n24 585
R441 B.n535 B.n25 585
R442 B.n533 B.n532 585
R443 B.n534 B.n533 585
R444 B.n531 B.n30 585
R445 B.n30 B.n29 585
R446 B.n530 B.n529 585
R447 B.n529 B.n528 585
R448 B.n32 B.n31 585
R449 B.n527 B.n32 585
R450 B.n525 B.n524 585
R451 B.n526 B.n525 585
R452 B.n523 B.n37 585
R453 B.n37 B.n36 585
R454 B.n522 B.n521 585
R455 B.n521 B.n520 585
R456 B.n39 B.n38 585
R457 B.n519 B.n39 585
R458 B.n517 B.n516 585
R459 B.n518 B.n517 585
R460 B.n515 B.n44 585
R461 B.n44 B.n43 585
R462 B.n514 B.n513 585
R463 B.n513 B.n512 585
R464 B.n46 B.n45 585
R465 B.n511 B.n46 585
R466 B.n509 B.n508 585
R467 B.n510 B.n509 585
R468 B.n507 B.n51 585
R469 B.n51 B.n50 585
R470 B.n506 B.n505 585
R471 B.n505 B.n504 585
R472 B.n53 B.n52 585
R473 B.n503 B.n53 585
R474 B.n501 B.n500 585
R475 B.n502 B.n501 585
R476 B.n499 B.n58 585
R477 B.n58 B.n57 585
R478 B.n498 B.n497 585
R479 B.n497 B.n496 585
R480 B.n60 B.n59 585
R481 B.n495 B.n60 585
R482 B.n493 B.n492 585
R483 B.n494 B.n493 585
R484 B.n491 B.n65 585
R485 B.n65 B.n64 585
R486 B.n490 B.n489 585
R487 B.n489 B.n488 585
R488 B.n67 B.n66 585
R489 B.n487 B.n67 585
R490 B.n485 B.n484 585
R491 B.n486 B.n485 585
R492 B.n562 B.n561 585
R493 B.n561 B.n560 585
R494 B.n254 B.n167 526.135
R495 B.n485 B.n72 526.135
R496 B.n256 B.n165 526.135
R497 B.n92 B.n70 526.135
R498 B.n420 B.n71 256.663
R499 B.n422 B.n71 256.663
R500 B.n428 B.n71 256.663
R501 B.n430 B.n71 256.663
R502 B.n436 B.n71 256.663
R503 B.n438 B.n71 256.663
R504 B.n445 B.n71 256.663
R505 B.n447 B.n71 256.663
R506 B.n453 B.n71 256.663
R507 B.n455 B.n71 256.663
R508 B.n462 B.n71 256.663
R509 B.n464 B.n71 256.663
R510 B.n470 B.n71 256.663
R511 B.n472 B.n71 256.663
R512 B.n478 B.n71 256.663
R513 B.n480 B.n71 256.663
R514 B.n249 B.n166 256.663
R515 B.n169 B.n166 256.663
R516 B.n242 B.n166 256.663
R517 B.n236 B.n166 256.663
R518 B.n234 B.n166 256.663
R519 B.n227 B.n166 256.663
R520 B.n225 B.n166 256.663
R521 B.n219 B.n166 256.663
R522 B.n217 B.n166 256.663
R523 B.n211 B.n166 256.663
R524 B.n183 B.n166 256.663
R525 B.n205 B.n166 256.663
R526 B.n199 B.n166 256.663
R527 B.n197 B.n166 256.663
R528 B.n191 B.n166 256.663
R529 B.n189 B.n166 256.663
R530 B.n180 B.t15 223.457
R531 B.n174 B.t8 223.457
R532 B.n79 B.t12 223.457
R533 B.n85 B.t4 223.457
R534 B.n255 B.n166 192.173
R535 B.n486 B.n71 192.173
R536 B.n180 B.t17 186.436
R537 B.n85 B.t6 186.436
R538 B.n174 B.t11 186.436
R539 B.n79 B.t13 186.436
R540 B.n254 B.n161 163.367
R541 B.n262 B.n161 163.367
R542 B.n262 B.n159 163.367
R543 B.n266 B.n159 163.367
R544 B.n266 B.n153 163.367
R545 B.n274 B.n153 163.367
R546 B.n274 B.n151 163.367
R547 B.n278 B.n151 163.367
R548 B.n278 B.n145 163.367
R549 B.n286 B.n145 163.367
R550 B.n286 B.n143 163.367
R551 B.n290 B.n143 163.367
R552 B.n290 B.n137 163.367
R553 B.n298 B.n137 163.367
R554 B.n298 B.n135 163.367
R555 B.n302 B.n135 163.367
R556 B.n302 B.n129 163.367
R557 B.n310 B.n129 163.367
R558 B.n310 B.n127 163.367
R559 B.n314 B.n127 163.367
R560 B.n314 B.n121 163.367
R561 B.n322 B.n121 163.367
R562 B.n322 B.n119 163.367
R563 B.n326 B.n119 163.367
R564 B.n326 B.n113 163.367
R565 B.n334 B.n113 163.367
R566 B.n334 B.n111 163.367
R567 B.n338 B.n111 163.367
R568 B.n338 B.n105 163.367
R569 B.n347 B.n105 163.367
R570 B.n347 B.n103 163.367
R571 B.n351 B.n103 163.367
R572 B.n351 B.n98 163.367
R573 B.n360 B.n98 163.367
R574 B.n360 B.n96 163.367
R575 B.n364 B.n96 163.367
R576 B.n364 B.n2 163.367
R577 B.n561 B.n2 163.367
R578 B.n561 B.n3 163.367
R579 B.n557 B.n3 163.367
R580 B.n557 B.n9 163.367
R581 B.n553 B.n9 163.367
R582 B.n553 B.n11 163.367
R583 B.n549 B.n11 163.367
R584 B.n549 B.n15 163.367
R585 B.n545 B.n15 163.367
R586 B.n545 B.n17 163.367
R587 B.n541 B.n17 163.367
R588 B.n541 B.n23 163.367
R589 B.n537 B.n23 163.367
R590 B.n537 B.n25 163.367
R591 B.n533 B.n25 163.367
R592 B.n533 B.n30 163.367
R593 B.n529 B.n30 163.367
R594 B.n529 B.n32 163.367
R595 B.n525 B.n32 163.367
R596 B.n525 B.n37 163.367
R597 B.n521 B.n37 163.367
R598 B.n521 B.n39 163.367
R599 B.n517 B.n39 163.367
R600 B.n517 B.n44 163.367
R601 B.n513 B.n44 163.367
R602 B.n513 B.n46 163.367
R603 B.n509 B.n46 163.367
R604 B.n509 B.n51 163.367
R605 B.n505 B.n51 163.367
R606 B.n505 B.n53 163.367
R607 B.n501 B.n53 163.367
R608 B.n501 B.n58 163.367
R609 B.n497 B.n58 163.367
R610 B.n497 B.n60 163.367
R611 B.n493 B.n60 163.367
R612 B.n493 B.n65 163.367
R613 B.n489 B.n65 163.367
R614 B.n489 B.n67 163.367
R615 B.n485 B.n67 163.367
R616 B.n250 B.n248 163.367
R617 B.n248 B.n247 163.367
R618 B.n244 B.n243 163.367
R619 B.n241 B.n171 163.367
R620 B.n237 B.n235 163.367
R621 B.n233 B.n173 163.367
R622 B.n228 B.n226 163.367
R623 B.n224 B.n177 163.367
R624 B.n220 B.n218 163.367
R625 B.n216 B.n179 163.367
R626 B.n212 B.n210 163.367
R627 B.n207 B.n206 163.367
R628 B.n204 B.n185 163.367
R629 B.n200 B.n198 163.367
R630 B.n196 B.n187 163.367
R631 B.n192 B.n190 163.367
R632 B.n256 B.n163 163.367
R633 B.n260 B.n163 163.367
R634 B.n260 B.n157 163.367
R635 B.n268 B.n157 163.367
R636 B.n268 B.n155 163.367
R637 B.n272 B.n155 163.367
R638 B.n272 B.n149 163.367
R639 B.n280 B.n149 163.367
R640 B.n280 B.n147 163.367
R641 B.n284 B.n147 163.367
R642 B.n284 B.n141 163.367
R643 B.n292 B.n141 163.367
R644 B.n292 B.n139 163.367
R645 B.n296 B.n139 163.367
R646 B.n296 B.n133 163.367
R647 B.n304 B.n133 163.367
R648 B.n304 B.n131 163.367
R649 B.n308 B.n131 163.367
R650 B.n308 B.n124 163.367
R651 B.n316 B.n124 163.367
R652 B.n316 B.n122 163.367
R653 B.n320 B.n122 163.367
R654 B.n320 B.n117 163.367
R655 B.n328 B.n117 163.367
R656 B.n328 B.n115 163.367
R657 B.n332 B.n115 163.367
R658 B.n332 B.n109 163.367
R659 B.n340 B.n109 163.367
R660 B.n340 B.n107 163.367
R661 B.n344 B.n107 163.367
R662 B.n344 B.n102 163.367
R663 B.n353 B.n102 163.367
R664 B.n353 B.n100 163.367
R665 B.n358 B.n100 163.367
R666 B.n358 B.n94 163.367
R667 B.n366 B.n94 163.367
R668 B.n367 B.n366 163.367
R669 B.n367 B.n5 163.367
R670 B.n6 B.n5 163.367
R671 B.n7 B.n6 163.367
R672 B.n372 B.n7 163.367
R673 B.n372 B.n12 163.367
R674 B.n13 B.n12 163.367
R675 B.n14 B.n13 163.367
R676 B.n377 B.n14 163.367
R677 B.n377 B.n19 163.367
R678 B.n20 B.n19 163.367
R679 B.n21 B.n20 163.367
R680 B.n382 B.n21 163.367
R681 B.n382 B.n26 163.367
R682 B.n27 B.n26 163.367
R683 B.n28 B.n27 163.367
R684 B.n387 B.n28 163.367
R685 B.n387 B.n33 163.367
R686 B.n34 B.n33 163.367
R687 B.n35 B.n34 163.367
R688 B.n392 B.n35 163.367
R689 B.n392 B.n40 163.367
R690 B.n41 B.n40 163.367
R691 B.n42 B.n41 163.367
R692 B.n397 B.n42 163.367
R693 B.n397 B.n47 163.367
R694 B.n48 B.n47 163.367
R695 B.n49 B.n48 163.367
R696 B.n402 B.n49 163.367
R697 B.n402 B.n54 163.367
R698 B.n55 B.n54 163.367
R699 B.n56 B.n55 163.367
R700 B.n407 B.n56 163.367
R701 B.n407 B.n61 163.367
R702 B.n62 B.n61 163.367
R703 B.n63 B.n62 163.367
R704 B.n412 B.n63 163.367
R705 B.n412 B.n68 163.367
R706 B.n69 B.n68 163.367
R707 B.n70 B.n69 163.367
R708 B.n481 B.n479 163.367
R709 B.n477 B.n74 163.367
R710 B.n473 B.n471 163.367
R711 B.n469 B.n76 163.367
R712 B.n465 B.n463 163.367
R713 B.n461 B.n78 163.367
R714 B.n456 B.n454 163.367
R715 B.n452 B.n82 163.367
R716 B.n448 B.n446 163.367
R717 B.n444 B.n84 163.367
R718 B.n439 B.n437 163.367
R719 B.n435 B.n88 163.367
R720 B.n431 B.n429 163.367
R721 B.n427 B.n90 163.367
R722 B.n423 B.n421 163.367
R723 B.n419 B.n92 163.367
R724 B.n181 B.t16 120.692
R725 B.n86 B.t7 120.692
R726 B.n175 B.t10 120.692
R727 B.n80 B.t14 120.692
R728 B.n255 B.n162 104.543
R729 B.n261 B.n162 104.543
R730 B.n261 B.n158 104.543
R731 B.n267 B.n158 104.543
R732 B.n267 B.n154 104.543
R733 B.n273 B.n154 104.543
R734 B.n273 B.n150 104.543
R735 B.n279 B.n150 104.543
R736 B.n285 B.n146 104.543
R737 B.n285 B.n142 104.543
R738 B.n291 B.n142 104.543
R739 B.n291 B.n138 104.543
R740 B.n297 B.n138 104.543
R741 B.n297 B.n134 104.543
R742 B.n303 B.n134 104.543
R743 B.n303 B.n130 104.543
R744 B.n309 B.n130 104.543
R745 B.n309 B.n125 104.543
R746 B.n315 B.n125 104.543
R747 B.n315 B.n126 104.543
R748 B.n321 B.n118 104.543
R749 B.n327 B.n118 104.543
R750 B.n327 B.n114 104.543
R751 B.n333 B.n114 104.543
R752 B.n333 B.n110 104.543
R753 B.n339 B.n110 104.543
R754 B.n339 B.n106 104.543
R755 B.n346 B.n106 104.543
R756 B.n346 B.n345 104.543
R757 B.n352 B.n99 104.543
R758 B.n359 B.n99 104.543
R759 B.n359 B.n95 104.543
R760 B.n365 B.n95 104.543
R761 B.n365 B.n4 104.543
R762 B.n560 B.n4 104.543
R763 B.n560 B.n559 104.543
R764 B.n559 B.n558 104.543
R765 B.n558 B.n8 104.543
R766 B.n552 B.n8 104.543
R767 B.n552 B.n551 104.543
R768 B.n551 B.n550 104.543
R769 B.n544 B.n18 104.543
R770 B.n544 B.n543 104.543
R771 B.n543 B.n542 104.543
R772 B.n542 B.n22 104.543
R773 B.n536 B.n22 104.543
R774 B.n536 B.n535 104.543
R775 B.n535 B.n534 104.543
R776 B.n534 B.n29 104.543
R777 B.n528 B.n29 104.543
R778 B.n527 B.n526 104.543
R779 B.n526 B.n36 104.543
R780 B.n520 B.n36 104.543
R781 B.n520 B.n519 104.543
R782 B.n519 B.n518 104.543
R783 B.n518 B.n43 104.543
R784 B.n512 B.n43 104.543
R785 B.n512 B.n511 104.543
R786 B.n511 B.n510 104.543
R787 B.n510 B.n50 104.543
R788 B.n504 B.n50 104.543
R789 B.n504 B.n503 104.543
R790 B.n502 B.n57 104.543
R791 B.n496 B.n57 104.543
R792 B.n496 B.n495 104.543
R793 B.n495 B.n494 104.543
R794 B.n494 B.n64 104.543
R795 B.n488 B.n64 104.543
R796 B.n488 B.n487 104.543
R797 B.n487 B.n486 104.543
R798 B.t9 B.n146 76.8698
R799 B.n503 B.t5 76.8698
R800 B.n249 B.n167 71.676
R801 B.n247 B.n169 71.676
R802 B.n243 B.n242 71.676
R803 B.n236 B.n171 71.676
R804 B.n235 B.n234 71.676
R805 B.n227 B.n173 71.676
R806 B.n226 B.n225 71.676
R807 B.n219 B.n177 71.676
R808 B.n218 B.n217 71.676
R809 B.n211 B.n179 71.676
R810 B.n210 B.n183 71.676
R811 B.n206 B.n205 71.676
R812 B.n199 B.n185 71.676
R813 B.n198 B.n197 71.676
R814 B.n191 B.n187 71.676
R815 B.n190 B.n189 71.676
R816 B.n480 B.n72 71.676
R817 B.n479 B.n478 71.676
R818 B.n472 B.n74 71.676
R819 B.n471 B.n470 71.676
R820 B.n464 B.n76 71.676
R821 B.n463 B.n462 71.676
R822 B.n455 B.n78 71.676
R823 B.n454 B.n453 71.676
R824 B.n447 B.n82 71.676
R825 B.n446 B.n445 71.676
R826 B.n438 B.n84 71.676
R827 B.n437 B.n436 71.676
R828 B.n430 B.n88 71.676
R829 B.n429 B.n428 71.676
R830 B.n422 B.n90 71.676
R831 B.n421 B.n420 71.676
R832 B.n420 B.n419 71.676
R833 B.n423 B.n422 71.676
R834 B.n428 B.n427 71.676
R835 B.n431 B.n430 71.676
R836 B.n436 B.n435 71.676
R837 B.n439 B.n438 71.676
R838 B.n445 B.n444 71.676
R839 B.n448 B.n447 71.676
R840 B.n453 B.n452 71.676
R841 B.n456 B.n455 71.676
R842 B.n462 B.n461 71.676
R843 B.n465 B.n464 71.676
R844 B.n470 B.n469 71.676
R845 B.n473 B.n472 71.676
R846 B.n478 B.n477 71.676
R847 B.n481 B.n480 71.676
R848 B.n250 B.n249 71.676
R849 B.n244 B.n169 71.676
R850 B.n242 B.n241 71.676
R851 B.n237 B.n236 71.676
R852 B.n234 B.n233 71.676
R853 B.n228 B.n227 71.676
R854 B.n225 B.n224 71.676
R855 B.n220 B.n219 71.676
R856 B.n217 B.n216 71.676
R857 B.n212 B.n211 71.676
R858 B.n207 B.n183 71.676
R859 B.n205 B.n204 71.676
R860 B.n200 B.n199 71.676
R861 B.n197 B.n196 71.676
R862 B.n192 B.n191 71.676
R863 B.n189 B.n165 71.676
R864 B.n181 B.n180 65.746
R865 B.n175 B.n174 65.746
R866 B.n80 B.n79 65.746
R867 B.n86 B.n85 65.746
R868 B.n352 B.t1 61.496
R869 B.n550 B.t3 61.496
R870 B.n182 B.n181 59.5399
R871 B.n230 B.n175 59.5399
R872 B.n459 B.n80 59.5399
R873 B.n441 B.n86 59.5399
R874 B.n321 B.t2 58.4212
R875 B.n528 B.t0 58.4212
R876 B.n126 B.t2 46.1221
R877 B.t0 B.n527 46.1221
R878 B.n345 B.t1 43.0473
R879 B.n18 B.t3 43.0473
R880 B.n484 B.n483 34.1859
R881 B.n417 B.n416 34.1859
R882 B.n257 B.n164 34.1859
R883 B.n253 B.n252 34.1859
R884 B.n279 B.t9 27.6735
R885 B.t5 B.n502 27.6735
R886 B B.n562 18.0485
R887 B.n483 B.n482 10.6151
R888 B.n482 B.n73 10.6151
R889 B.n476 B.n73 10.6151
R890 B.n476 B.n475 10.6151
R891 B.n475 B.n474 10.6151
R892 B.n474 B.n75 10.6151
R893 B.n468 B.n75 10.6151
R894 B.n468 B.n467 10.6151
R895 B.n467 B.n466 10.6151
R896 B.n466 B.n77 10.6151
R897 B.n460 B.n77 10.6151
R898 B.n458 B.n457 10.6151
R899 B.n457 B.n81 10.6151
R900 B.n451 B.n81 10.6151
R901 B.n451 B.n450 10.6151
R902 B.n450 B.n449 10.6151
R903 B.n449 B.n83 10.6151
R904 B.n443 B.n83 10.6151
R905 B.n443 B.n442 10.6151
R906 B.n440 B.n87 10.6151
R907 B.n434 B.n87 10.6151
R908 B.n434 B.n433 10.6151
R909 B.n433 B.n432 10.6151
R910 B.n432 B.n89 10.6151
R911 B.n426 B.n89 10.6151
R912 B.n426 B.n425 10.6151
R913 B.n425 B.n424 10.6151
R914 B.n424 B.n91 10.6151
R915 B.n418 B.n91 10.6151
R916 B.n418 B.n417 10.6151
R917 B.n258 B.n257 10.6151
R918 B.n259 B.n258 10.6151
R919 B.n259 B.n156 10.6151
R920 B.n269 B.n156 10.6151
R921 B.n270 B.n269 10.6151
R922 B.n271 B.n270 10.6151
R923 B.n271 B.n148 10.6151
R924 B.n281 B.n148 10.6151
R925 B.n282 B.n281 10.6151
R926 B.n283 B.n282 10.6151
R927 B.n283 B.n140 10.6151
R928 B.n293 B.n140 10.6151
R929 B.n294 B.n293 10.6151
R930 B.n295 B.n294 10.6151
R931 B.n295 B.n132 10.6151
R932 B.n305 B.n132 10.6151
R933 B.n306 B.n305 10.6151
R934 B.n307 B.n306 10.6151
R935 B.n307 B.n123 10.6151
R936 B.n317 B.n123 10.6151
R937 B.n318 B.n317 10.6151
R938 B.n319 B.n318 10.6151
R939 B.n319 B.n116 10.6151
R940 B.n329 B.n116 10.6151
R941 B.n330 B.n329 10.6151
R942 B.n331 B.n330 10.6151
R943 B.n331 B.n108 10.6151
R944 B.n341 B.n108 10.6151
R945 B.n342 B.n341 10.6151
R946 B.n343 B.n342 10.6151
R947 B.n343 B.n101 10.6151
R948 B.n354 B.n101 10.6151
R949 B.n355 B.n354 10.6151
R950 B.n357 B.n355 10.6151
R951 B.n357 B.n356 10.6151
R952 B.n356 B.n93 10.6151
R953 B.n368 B.n93 10.6151
R954 B.n369 B.n368 10.6151
R955 B.n370 B.n369 10.6151
R956 B.n371 B.n370 10.6151
R957 B.n373 B.n371 10.6151
R958 B.n374 B.n373 10.6151
R959 B.n375 B.n374 10.6151
R960 B.n376 B.n375 10.6151
R961 B.n378 B.n376 10.6151
R962 B.n379 B.n378 10.6151
R963 B.n380 B.n379 10.6151
R964 B.n381 B.n380 10.6151
R965 B.n383 B.n381 10.6151
R966 B.n384 B.n383 10.6151
R967 B.n385 B.n384 10.6151
R968 B.n386 B.n385 10.6151
R969 B.n388 B.n386 10.6151
R970 B.n389 B.n388 10.6151
R971 B.n390 B.n389 10.6151
R972 B.n391 B.n390 10.6151
R973 B.n393 B.n391 10.6151
R974 B.n394 B.n393 10.6151
R975 B.n395 B.n394 10.6151
R976 B.n396 B.n395 10.6151
R977 B.n398 B.n396 10.6151
R978 B.n399 B.n398 10.6151
R979 B.n400 B.n399 10.6151
R980 B.n401 B.n400 10.6151
R981 B.n403 B.n401 10.6151
R982 B.n404 B.n403 10.6151
R983 B.n405 B.n404 10.6151
R984 B.n406 B.n405 10.6151
R985 B.n408 B.n406 10.6151
R986 B.n409 B.n408 10.6151
R987 B.n410 B.n409 10.6151
R988 B.n411 B.n410 10.6151
R989 B.n413 B.n411 10.6151
R990 B.n414 B.n413 10.6151
R991 B.n415 B.n414 10.6151
R992 B.n416 B.n415 10.6151
R993 B.n252 B.n251 10.6151
R994 B.n251 B.n168 10.6151
R995 B.n246 B.n168 10.6151
R996 B.n246 B.n245 10.6151
R997 B.n245 B.n170 10.6151
R998 B.n240 B.n170 10.6151
R999 B.n240 B.n239 10.6151
R1000 B.n239 B.n238 10.6151
R1001 B.n238 B.n172 10.6151
R1002 B.n232 B.n172 10.6151
R1003 B.n232 B.n231 10.6151
R1004 B.n229 B.n176 10.6151
R1005 B.n223 B.n176 10.6151
R1006 B.n223 B.n222 10.6151
R1007 B.n222 B.n221 10.6151
R1008 B.n221 B.n178 10.6151
R1009 B.n215 B.n178 10.6151
R1010 B.n215 B.n214 10.6151
R1011 B.n214 B.n213 10.6151
R1012 B.n209 B.n208 10.6151
R1013 B.n208 B.n184 10.6151
R1014 B.n203 B.n184 10.6151
R1015 B.n203 B.n202 10.6151
R1016 B.n202 B.n201 10.6151
R1017 B.n201 B.n186 10.6151
R1018 B.n195 B.n186 10.6151
R1019 B.n195 B.n194 10.6151
R1020 B.n194 B.n193 10.6151
R1021 B.n193 B.n188 10.6151
R1022 B.n188 B.n164 10.6151
R1023 B.n253 B.n160 10.6151
R1024 B.n263 B.n160 10.6151
R1025 B.n264 B.n263 10.6151
R1026 B.n265 B.n264 10.6151
R1027 B.n265 B.n152 10.6151
R1028 B.n275 B.n152 10.6151
R1029 B.n276 B.n275 10.6151
R1030 B.n277 B.n276 10.6151
R1031 B.n277 B.n144 10.6151
R1032 B.n287 B.n144 10.6151
R1033 B.n288 B.n287 10.6151
R1034 B.n289 B.n288 10.6151
R1035 B.n289 B.n136 10.6151
R1036 B.n299 B.n136 10.6151
R1037 B.n300 B.n299 10.6151
R1038 B.n301 B.n300 10.6151
R1039 B.n301 B.n128 10.6151
R1040 B.n311 B.n128 10.6151
R1041 B.n312 B.n311 10.6151
R1042 B.n313 B.n312 10.6151
R1043 B.n313 B.n120 10.6151
R1044 B.n323 B.n120 10.6151
R1045 B.n324 B.n323 10.6151
R1046 B.n325 B.n324 10.6151
R1047 B.n325 B.n112 10.6151
R1048 B.n335 B.n112 10.6151
R1049 B.n336 B.n335 10.6151
R1050 B.n337 B.n336 10.6151
R1051 B.n337 B.n104 10.6151
R1052 B.n348 B.n104 10.6151
R1053 B.n349 B.n348 10.6151
R1054 B.n350 B.n349 10.6151
R1055 B.n350 B.n97 10.6151
R1056 B.n361 B.n97 10.6151
R1057 B.n362 B.n361 10.6151
R1058 B.n363 B.n362 10.6151
R1059 B.n363 B.n0 10.6151
R1060 B.n556 B.n1 10.6151
R1061 B.n556 B.n555 10.6151
R1062 B.n555 B.n554 10.6151
R1063 B.n554 B.n10 10.6151
R1064 B.n548 B.n10 10.6151
R1065 B.n548 B.n547 10.6151
R1066 B.n547 B.n546 10.6151
R1067 B.n546 B.n16 10.6151
R1068 B.n540 B.n16 10.6151
R1069 B.n540 B.n539 10.6151
R1070 B.n539 B.n538 10.6151
R1071 B.n538 B.n24 10.6151
R1072 B.n532 B.n24 10.6151
R1073 B.n532 B.n531 10.6151
R1074 B.n531 B.n530 10.6151
R1075 B.n530 B.n31 10.6151
R1076 B.n524 B.n31 10.6151
R1077 B.n524 B.n523 10.6151
R1078 B.n523 B.n522 10.6151
R1079 B.n522 B.n38 10.6151
R1080 B.n516 B.n38 10.6151
R1081 B.n516 B.n515 10.6151
R1082 B.n515 B.n514 10.6151
R1083 B.n514 B.n45 10.6151
R1084 B.n508 B.n45 10.6151
R1085 B.n508 B.n507 10.6151
R1086 B.n507 B.n506 10.6151
R1087 B.n506 B.n52 10.6151
R1088 B.n500 B.n52 10.6151
R1089 B.n500 B.n499 10.6151
R1090 B.n499 B.n498 10.6151
R1091 B.n498 B.n59 10.6151
R1092 B.n492 B.n59 10.6151
R1093 B.n492 B.n491 10.6151
R1094 B.n491 B.n490 10.6151
R1095 B.n490 B.n66 10.6151
R1096 B.n484 B.n66 10.6151
R1097 B.n459 B.n458 6.5566
R1098 B.n442 B.n441 6.5566
R1099 B.n230 B.n229 6.5566
R1100 B.n213 B.n182 6.5566
R1101 B.n460 B.n459 4.05904
R1102 B.n441 B.n440 4.05904
R1103 B.n231 B.n230 4.05904
R1104 B.n209 B.n182 4.05904
R1105 B.n562 B.n0 2.81026
R1106 B.n562 B.n1 2.81026
R1107 VP.n15 VP.n14 161.3
R1108 VP.n13 VP.n1 161.3
R1109 VP.n12 VP.n11 161.3
R1110 VP.n10 VP.n2 161.3
R1111 VP.n9 VP.n8 161.3
R1112 VP.n7 VP.n3 161.3
R1113 VP.n6 VP.n5 68.3588
R1114 VP.n16 VP.n0 68.3588
R1115 VP.n12 VP.n2 56.5617
R1116 VP.n4 VP.t3 49.3751
R1117 VP.n4 VP.t2 48.3688
R1118 VP.n5 VP.n4 43.0323
R1119 VP.n8 VP.n7 24.5923
R1120 VP.n8 VP.n2 24.5923
R1121 VP.n13 VP.n12 24.5923
R1122 VP.n14 VP.n13 24.5923
R1123 VP.n7 VP.n6 21.8872
R1124 VP.n14 VP.n0 21.8872
R1125 VP.n6 VP.t1 14.807
R1126 VP.n0 VP.t0 14.807
R1127 VP.n5 VP.n3 0.354861
R1128 VP.n16 VP.n15 0.354861
R1129 VP VP.n16 0.267071
R1130 VP.n9 VP.n3 0.189894
R1131 VP.n10 VP.n9 0.189894
R1132 VP.n11 VP.n10 0.189894
R1133 VP.n11 VP.n1 0.189894
R1134 VP.n15 VP.n1 0.189894
R1135 VDD1 VDD1.n1 137.989
R1136 VDD1 VDD1.n0 103.421
R1137 VDD1.n0 VDD1.t0 10.5324
R1138 VDD1.n0 VDD1.t1 10.5324
R1139 VDD1.n1 VDD1.t2 10.5324
R1140 VDD1.n1 VDD1.t3 10.5324
C0 VN VDD2 1.04068f
C1 VN VTAIL 1.72753f
C2 VN VP 4.65148f
C3 VDD1 VN 0.155777f
C4 VDD2 VTAIL 3.29774f
C5 VP VDD2 0.430939f
C6 VP VTAIL 1.74163f
C7 VDD1 VDD2 1.1391f
C8 VDD1 VTAIL 3.24045f
C9 VDD1 VP 1.31381f
C10 VDD2 B 3.188502f
C11 VDD1 B 5.72504f
C12 VTAIL B 3.757979f
C13 VN B 10.2727f
C14 VP B 8.980615f
C15 VDD1.t0 B 0.031655f
C16 VDD1.t1 B 0.031655f
C17 VDD1.n0 B 0.203516f
C18 VDD1.t2 B 0.031655f
C19 VDD1.t3 B 0.031655f
C20 VDD1.n1 B 0.415743f
C21 VP.t0 B 0.28319f
C22 VP.n0 B 0.22229f
C23 VP.n1 B 0.021351f
C24 VP.n2 B 0.031037f
C25 VP.n3 B 0.034455f
C26 VP.t1 B 0.28319f
C27 VP.t3 B 0.485934f
C28 VP.t2 B 0.479864f
C29 VP.n4 B 1.30837f
C30 VP.n5 B 0.956565f
C31 VP.n6 B 0.22229f
C32 VP.n7 B 0.037443f
C33 VP.n8 B 0.039593f
C34 VP.n9 B 0.021351f
C35 VP.n10 B 0.021351f
C36 VP.n11 B 0.021351f
C37 VP.n12 B 0.031037f
C38 VP.n13 B 0.039593f
C39 VP.n14 B 0.037443f
C40 VP.n15 B 0.034455f
C41 VP.n16 B 0.043001f
C42 VTAIL.n0 B 0.025657f
C43 VTAIL.n1 B 0.060155f
C44 VTAIL.t7 B 0.042577f
C45 VTAIL.n2 B 0.044374f
C46 VTAIL.n3 B 0.01232f
C47 VTAIL.n4 B 0.01f
C48 VTAIL.n5 B 0.118497f
C49 VTAIL.n6 B 0.028193f
C50 VTAIL.n7 B 0.138061f
C51 VTAIL.n8 B 0.025657f
C52 VTAIL.n9 B 0.060155f
C53 VTAIL.t1 B 0.042577f
C54 VTAIL.n10 B 0.044374f
C55 VTAIL.n11 B 0.01232f
C56 VTAIL.n12 B 0.01f
C57 VTAIL.n13 B 0.118497f
C58 VTAIL.n14 B 0.028193f
C59 VTAIL.n15 B 0.222196f
C60 VTAIL.n16 B 0.025657f
C61 VTAIL.n17 B 0.060155f
C62 VTAIL.t2 B 0.042577f
C63 VTAIL.n18 B 0.044374f
C64 VTAIL.n19 B 0.01232f
C65 VTAIL.n20 B 0.01f
C66 VTAIL.n21 B 0.118497f
C67 VTAIL.n22 B 0.028193f
C68 VTAIL.n23 B 0.719261f
C69 VTAIL.n24 B 0.025657f
C70 VTAIL.n25 B 0.060155f
C71 VTAIL.t4 B 0.042577f
C72 VTAIL.n26 B 0.044374f
C73 VTAIL.n27 B 0.01232f
C74 VTAIL.n28 B 0.01f
C75 VTAIL.n29 B 0.118497f
C76 VTAIL.n30 B 0.028193f
C77 VTAIL.n31 B 0.719261f
C78 VTAIL.n32 B 0.025657f
C79 VTAIL.n33 B 0.060155f
C80 VTAIL.t5 B 0.042577f
C81 VTAIL.n34 B 0.044374f
C82 VTAIL.n35 B 0.01232f
C83 VTAIL.n36 B 0.01f
C84 VTAIL.n37 B 0.118497f
C85 VTAIL.n38 B 0.028193f
C86 VTAIL.n39 B 0.222196f
C87 VTAIL.n40 B 0.025657f
C88 VTAIL.n41 B 0.060155f
C89 VTAIL.t3 B 0.042577f
C90 VTAIL.n42 B 0.044374f
C91 VTAIL.n43 B 0.01232f
C92 VTAIL.n44 B 0.01f
C93 VTAIL.n45 B 0.118497f
C94 VTAIL.n46 B 0.028193f
C95 VTAIL.n47 B 0.222196f
C96 VTAIL.n48 B 0.025657f
C97 VTAIL.n49 B 0.060155f
C98 VTAIL.t0 B 0.042577f
C99 VTAIL.n50 B 0.044374f
C100 VTAIL.n51 B 0.01232f
C101 VTAIL.n52 B 0.01f
C102 VTAIL.n53 B 0.118497f
C103 VTAIL.n54 B 0.028193f
C104 VTAIL.n55 B 0.719261f
C105 VTAIL.n56 B 0.025657f
C106 VTAIL.n57 B 0.060155f
C107 VTAIL.t6 B 0.042577f
C108 VTAIL.n58 B 0.044374f
C109 VTAIL.n59 B 0.01232f
C110 VTAIL.n60 B 0.01f
C111 VTAIL.n61 B 0.118497f
C112 VTAIL.n62 B 0.028193f
C113 VTAIL.n63 B 0.628147f
C114 VDD2.t0 B 0.033467f
C115 VDD2.t1 B 0.033467f
C116 VDD2.n0 B 0.425706f
C117 VDD2.t2 B 0.033467f
C118 VDD2.t3 B 0.033467f
C119 VDD2.n1 B 0.21495f
C120 VDD2.n2 B 2.30849f
C121 VN.t1 B 0.476819f
C122 VN.t0 B 0.482851f
C123 VN.n0 B 0.309103f
C124 VN.t2 B 0.482851f
C125 VN.t3 B 0.476819f
C126 VN.n1 B 1.30913f
.ends

