* NGSPICE file created from diff_pair_sample_0840.ext - technology: sky130A

.subckt diff_pair_sample_0840 VTAIL VN VP B VDD2 VDD1
X0 B.t17 B.t15 B.t16 B.t9 sky130_fd_pr__nfet_01v8 ad=7.7688 pd=40.62 as=0 ps=0 w=19.92 l=2.86
X1 VTAIL.t7 VN.t0 VDD2.t3 B.t2 sky130_fd_pr__nfet_01v8 ad=7.7688 pd=40.62 as=3.2868 ps=20.25 w=19.92 l=2.86
X2 B.t14 B.t12 B.t13 B.t5 sky130_fd_pr__nfet_01v8 ad=7.7688 pd=40.62 as=0 ps=0 w=19.92 l=2.86
X3 VDD2.t0 VN.t1 VTAIL.t6 B.t3 sky130_fd_pr__nfet_01v8 ad=3.2868 pd=20.25 as=7.7688 ps=40.62 w=19.92 l=2.86
X4 VDD1.t3 VP.t0 VTAIL.t3 B.t1 sky130_fd_pr__nfet_01v8 ad=3.2868 pd=20.25 as=7.7688 ps=40.62 w=19.92 l=2.86
X5 VTAIL.t0 VP.t1 VDD1.t2 B.t0 sky130_fd_pr__nfet_01v8 ad=7.7688 pd=40.62 as=3.2868 ps=20.25 w=19.92 l=2.86
X6 VTAIL.t5 VN.t2 VDD2.t1 B.t0 sky130_fd_pr__nfet_01v8 ad=7.7688 pd=40.62 as=3.2868 ps=20.25 w=19.92 l=2.86
X7 VDD1.t1 VP.t2 VTAIL.t2 B.t3 sky130_fd_pr__nfet_01v8 ad=3.2868 pd=20.25 as=7.7688 ps=40.62 w=19.92 l=2.86
X8 VDD2.t2 VN.t3 VTAIL.t4 B.t1 sky130_fd_pr__nfet_01v8 ad=3.2868 pd=20.25 as=7.7688 ps=40.62 w=19.92 l=2.86
X9 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=7.7688 pd=40.62 as=0 ps=0 w=19.92 l=2.86
X10 B.t7 B.t4 B.t6 B.t5 sky130_fd_pr__nfet_01v8 ad=7.7688 pd=40.62 as=0 ps=0 w=19.92 l=2.86
X11 VTAIL.t1 VP.t3 VDD1.t0 B.t2 sky130_fd_pr__nfet_01v8 ad=7.7688 pd=40.62 as=3.2868 ps=20.25 w=19.92 l=2.86
R0 B.n996 B.n995 585
R1 B.n997 B.n996 585
R2 B.n417 B.n138 585
R3 B.n416 B.n415 585
R4 B.n414 B.n413 585
R5 B.n412 B.n411 585
R6 B.n410 B.n409 585
R7 B.n408 B.n407 585
R8 B.n406 B.n405 585
R9 B.n404 B.n403 585
R10 B.n402 B.n401 585
R11 B.n400 B.n399 585
R12 B.n398 B.n397 585
R13 B.n396 B.n395 585
R14 B.n394 B.n393 585
R15 B.n392 B.n391 585
R16 B.n390 B.n389 585
R17 B.n388 B.n387 585
R18 B.n386 B.n385 585
R19 B.n384 B.n383 585
R20 B.n382 B.n381 585
R21 B.n380 B.n379 585
R22 B.n378 B.n377 585
R23 B.n376 B.n375 585
R24 B.n374 B.n373 585
R25 B.n372 B.n371 585
R26 B.n370 B.n369 585
R27 B.n368 B.n367 585
R28 B.n366 B.n365 585
R29 B.n364 B.n363 585
R30 B.n362 B.n361 585
R31 B.n360 B.n359 585
R32 B.n358 B.n357 585
R33 B.n356 B.n355 585
R34 B.n354 B.n353 585
R35 B.n352 B.n351 585
R36 B.n350 B.n349 585
R37 B.n348 B.n347 585
R38 B.n346 B.n345 585
R39 B.n344 B.n343 585
R40 B.n342 B.n341 585
R41 B.n340 B.n339 585
R42 B.n338 B.n337 585
R43 B.n336 B.n335 585
R44 B.n334 B.n333 585
R45 B.n332 B.n331 585
R46 B.n330 B.n329 585
R47 B.n328 B.n327 585
R48 B.n326 B.n325 585
R49 B.n324 B.n323 585
R50 B.n322 B.n321 585
R51 B.n320 B.n319 585
R52 B.n318 B.n317 585
R53 B.n316 B.n315 585
R54 B.n314 B.n313 585
R55 B.n312 B.n311 585
R56 B.n310 B.n309 585
R57 B.n308 B.n307 585
R58 B.n306 B.n305 585
R59 B.n304 B.n303 585
R60 B.n302 B.n301 585
R61 B.n300 B.n299 585
R62 B.n298 B.n297 585
R63 B.n296 B.n295 585
R64 B.n294 B.n293 585
R65 B.n292 B.n291 585
R66 B.n290 B.n289 585
R67 B.n288 B.n287 585
R68 B.n286 B.n285 585
R69 B.n284 B.n283 585
R70 B.n282 B.n281 585
R71 B.n280 B.n279 585
R72 B.n278 B.n277 585
R73 B.n276 B.n275 585
R74 B.n274 B.n273 585
R75 B.n271 B.n270 585
R76 B.n269 B.n268 585
R77 B.n267 B.n266 585
R78 B.n265 B.n264 585
R79 B.n263 B.n262 585
R80 B.n261 B.n260 585
R81 B.n259 B.n258 585
R82 B.n257 B.n256 585
R83 B.n255 B.n254 585
R84 B.n253 B.n252 585
R85 B.n251 B.n250 585
R86 B.n249 B.n248 585
R87 B.n247 B.n246 585
R88 B.n245 B.n244 585
R89 B.n243 B.n242 585
R90 B.n241 B.n240 585
R91 B.n239 B.n238 585
R92 B.n237 B.n236 585
R93 B.n235 B.n234 585
R94 B.n233 B.n232 585
R95 B.n231 B.n230 585
R96 B.n229 B.n228 585
R97 B.n227 B.n226 585
R98 B.n225 B.n224 585
R99 B.n223 B.n222 585
R100 B.n221 B.n220 585
R101 B.n219 B.n218 585
R102 B.n217 B.n216 585
R103 B.n215 B.n214 585
R104 B.n213 B.n212 585
R105 B.n211 B.n210 585
R106 B.n209 B.n208 585
R107 B.n207 B.n206 585
R108 B.n205 B.n204 585
R109 B.n203 B.n202 585
R110 B.n201 B.n200 585
R111 B.n199 B.n198 585
R112 B.n197 B.n196 585
R113 B.n195 B.n194 585
R114 B.n193 B.n192 585
R115 B.n191 B.n190 585
R116 B.n189 B.n188 585
R117 B.n187 B.n186 585
R118 B.n185 B.n184 585
R119 B.n183 B.n182 585
R120 B.n181 B.n180 585
R121 B.n179 B.n178 585
R122 B.n177 B.n176 585
R123 B.n175 B.n174 585
R124 B.n173 B.n172 585
R125 B.n171 B.n170 585
R126 B.n169 B.n168 585
R127 B.n167 B.n166 585
R128 B.n165 B.n164 585
R129 B.n163 B.n162 585
R130 B.n161 B.n160 585
R131 B.n159 B.n158 585
R132 B.n157 B.n156 585
R133 B.n155 B.n154 585
R134 B.n153 B.n152 585
R135 B.n151 B.n150 585
R136 B.n149 B.n148 585
R137 B.n147 B.n146 585
R138 B.n145 B.n144 585
R139 B.n67 B.n66 585
R140 B.n994 B.n68 585
R141 B.n998 B.n68 585
R142 B.n993 B.n992 585
R143 B.n992 B.n64 585
R144 B.n991 B.n63 585
R145 B.n1004 B.n63 585
R146 B.n990 B.n62 585
R147 B.n1005 B.n62 585
R148 B.n989 B.n61 585
R149 B.n1006 B.n61 585
R150 B.n988 B.n987 585
R151 B.n987 B.n57 585
R152 B.n986 B.n56 585
R153 B.n1012 B.n56 585
R154 B.n985 B.n55 585
R155 B.n1013 B.n55 585
R156 B.n984 B.n54 585
R157 B.n1014 B.n54 585
R158 B.n983 B.n982 585
R159 B.n982 B.n50 585
R160 B.n981 B.n49 585
R161 B.n1020 B.n49 585
R162 B.n980 B.n48 585
R163 B.n1021 B.n48 585
R164 B.n979 B.n47 585
R165 B.n1022 B.n47 585
R166 B.n978 B.n977 585
R167 B.n977 B.n43 585
R168 B.n976 B.n42 585
R169 B.n1028 B.n42 585
R170 B.n975 B.n41 585
R171 B.n1029 B.n41 585
R172 B.n974 B.n40 585
R173 B.n1030 B.n40 585
R174 B.n973 B.n972 585
R175 B.n972 B.n36 585
R176 B.n971 B.n35 585
R177 B.n1036 B.n35 585
R178 B.n970 B.n34 585
R179 B.n1037 B.n34 585
R180 B.n969 B.n33 585
R181 B.n1038 B.n33 585
R182 B.n968 B.n967 585
R183 B.n967 B.n29 585
R184 B.n966 B.n28 585
R185 B.n1044 B.n28 585
R186 B.n965 B.n27 585
R187 B.n1045 B.n27 585
R188 B.n964 B.n26 585
R189 B.n1046 B.n26 585
R190 B.n963 B.n962 585
R191 B.n962 B.n22 585
R192 B.n961 B.n21 585
R193 B.n1052 B.n21 585
R194 B.n960 B.n20 585
R195 B.n1053 B.n20 585
R196 B.n959 B.n19 585
R197 B.n1054 B.n19 585
R198 B.n958 B.n957 585
R199 B.n957 B.n18 585
R200 B.n956 B.n14 585
R201 B.n1060 B.n14 585
R202 B.n955 B.n13 585
R203 B.n1061 B.n13 585
R204 B.n954 B.n12 585
R205 B.n1062 B.n12 585
R206 B.n953 B.n952 585
R207 B.n952 B.n8 585
R208 B.n951 B.n7 585
R209 B.n1068 B.n7 585
R210 B.n950 B.n6 585
R211 B.n1069 B.n6 585
R212 B.n949 B.n5 585
R213 B.n1070 B.n5 585
R214 B.n948 B.n947 585
R215 B.n947 B.n4 585
R216 B.n946 B.n418 585
R217 B.n946 B.n945 585
R218 B.n936 B.n419 585
R219 B.n420 B.n419 585
R220 B.n938 B.n937 585
R221 B.n939 B.n938 585
R222 B.n935 B.n425 585
R223 B.n425 B.n424 585
R224 B.n934 B.n933 585
R225 B.n933 B.n932 585
R226 B.n427 B.n426 585
R227 B.n925 B.n427 585
R228 B.n924 B.n923 585
R229 B.n926 B.n924 585
R230 B.n922 B.n432 585
R231 B.n432 B.n431 585
R232 B.n921 B.n920 585
R233 B.n920 B.n919 585
R234 B.n434 B.n433 585
R235 B.n435 B.n434 585
R236 B.n912 B.n911 585
R237 B.n913 B.n912 585
R238 B.n910 B.n440 585
R239 B.n440 B.n439 585
R240 B.n909 B.n908 585
R241 B.n908 B.n907 585
R242 B.n442 B.n441 585
R243 B.n443 B.n442 585
R244 B.n900 B.n899 585
R245 B.n901 B.n900 585
R246 B.n898 B.n448 585
R247 B.n448 B.n447 585
R248 B.n897 B.n896 585
R249 B.n896 B.n895 585
R250 B.n450 B.n449 585
R251 B.n451 B.n450 585
R252 B.n888 B.n887 585
R253 B.n889 B.n888 585
R254 B.n886 B.n456 585
R255 B.n456 B.n455 585
R256 B.n885 B.n884 585
R257 B.n884 B.n883 585
R258 B.n458 B.n457 585
R259 B.n459 B.n458 585
R260 B.n876 B.n875 585
R261 B.n877 B.n876 585
R262 B.n874 B.n464 585
R263 B.n464 B.n463 585
R264 B.n873 B.n872 585
R265 B.n872 B.n871 585
R266 B.n466 B.n465 585
R267 B.n467 B.n466 585
R268 B.n864 B.n863 585
R269 B.n865 B.n864 585
R270 B.n862 B.n471 585
R271 B.n475 B.n471 585
R272 B.n861 B.n860 585
R273 B.n860 B.n859 585
R274 B.n473 B.n472 585
R275 B.n474 B.n473 585
R276 B.n852 B.n851 585
R277 B.n853 B.n852 585
R278 B.n850 B.n480 585
R279 B.n480 B.n479 585
R280 B.n849 B.n848 585
R281 B.n848 B.n847 585
R282 B.n482 B.n481 585
R283 B.n483 B.n482 585
R284 B.n840 B.n839 585
R285 B.n841 B.n840 585
R286 B.n486 B.n485 585
R287 B.n564 B.n563 585
R288 B.n565 B.n561 585
R289 B.n561 B.n487 585
R290 B.n567 B.n566 585
R291 B.n569 B.n560 585
R292 B.n572 B.n571 585
R293 B.n573 B.n559 585
R294 B.n575 B.n574 585
R295 B.n577 B.n558 585
R296 B.n580 B.n579 585
R297 B.n581 B.n557 585
R298 B.n583 B.n582 585
R299 B.n585 B.n556 585
R300 B.n588 B.n587 585
R301 B.n589 B.n555 585
R302 B.n591 B.n590 585
R303 B.n593 B.n554 585
R304 B.n596 B.n595 585
R305 B.n597 B.n553 585
R306 B.n599 B.n598 585
R307 B.n601 B.n552 585
R308 B.n604 B.n603 585
R309 B.n605 B.n551 585
R310 B.n607 B.n606 585
R311 B.n609 B.n550 585
R312 B.n612 B.n611 585
R313 B.n613 B.n549 585
R314 B.n615 B.n614 585
R315 B.n617 B.n548 585
R316 B.n620 B.n619 585
R317 B.n621 B.n547 585
R318 B.n623 B.n622 585
R319 B.n625 B.n546 585
R320 B.n628 B.n627 585
R321 B.n629 B.n545 585
R322 B.n631 B.n630 585
R323 B.n633 B.n544 585
R324 B.n636 B.n635 585
R325 B.n637 B.n543 585
R326 B.n639 B.n638 585
R327 B.n641 B.n542 585
R328 B.n644 B.n643 585
R329 B.n645 B.n541 585
R330 B.n647 B.n646 585
R331 B.n649 B.n540 585
R332 B.n652 B.n651 585
R333 B.n653 B.n539 585
R334 B.n655 B.n654 585
R335 B.n657 B.n538 585
R336 B.n660 B.n659 585
R337 B.n661 B.n537 585
R338 B.n663 B.n662 585
R339 B.n665 B.n536 585
R340 B.n668 B.n667 585
R341 B.n669 B.n535 585
R342 B.n671 B.n670 585
R343 B.n673 B.n534 585
R344 B.n676 B.n675 585
R345 B.n677 B.n533 585
R346 B.n679 B.n678 585
R347 B.n681 B.n532 585
R348 B.n684 B.n683 585
R349 B.n685 B.n531 585
R350 B.n687 B.n686 585
R351 B.n689 B.n530 585
R352 B.n692 B.n691 585
R353 B.n693 B.n526 585
R354 B.n695 B.n694 585
R355 B.n697 B.n525 585
R356 B.n700 B.n699 585
R357 B.n701 B.n524 585
R358 B.n703 B.n702 585
R359 B.n705 B.n523 585
R360 B.n708 B.n707 585
R361 B.n710 B.n520 585
R362 B.n712 B.n711 585
R363 B.n714 B.n519 585
R364 B.n717 B.n716 585
R365 B.n718 B.n518 585
R366 B.n720 B.n719 585
R367 B.n722 B.n517 585
R368 B.n725 B.n724 585
R369 B.n726 B.n516 585
R370 B.n728 B.n727 585
R371 B.n730 B.n515 585
R372 B.n733 B.n732 585
R373 B.n734 B.n514 585
R374 B.n736 B.n735 585
R375 B.n738 B.n513 585
R376 B.n741 B.n740 585
R377 B.n742 B.n512 585
R378 B.n744 B.n743 585
R379 B.n746 B.n511 585
R380 B.n749 B.n748 585
R381 B.n750 B.n510 585
R382 B.n752 B.n751 585
R383 B.n754 B.n509 585
R384 B.n757 B.n756 585
R385 B.n758 B.n508 585
R386 B.n760 B.n759 585
R387 B.n762 B.n507 585
R388 B.n765 B.n764 585
R389 B.n766 B.n506 585
R390 B.n768 B.n767 585
R391 B.n770 B.n505 585
R392 B.n773 B.n772 585
R393 B.n774 B.n504 585
R394 B.n776 B.n775 585
R395 B.n778 B.n503 585
R396 B.n781 B.n780 585
R397 B.n782 B.n502 585
R398 B.n784 B.n783 585
R399 B.n786 B.n501 585
R400 B.n789 B.n788 585
R401 B.n790 B.n500 585
R402 B.n792 B.n791 585
R403 B.n794 B.n499 585
R404 B.n797 B.n796 585
R405 B.n798 B.n498 585
R406 B.n800 B.n799 585
R407 B.n802 B.n497 585
R408 B.n805 B.n804 585
R409 B.n806 B.n496 585
R410 B.n808 B.n807 585
R411 B.n810 B.n495 585
R412 B.n813 B.n812 585
R413 B.n814 B.n494 585
R414 B.n816 B.n815 585
R415 B.n818 B.n493 585
R416 B.n821 B.n820 585
R417 B.n822 B.n492 585
R418 B.n824 B.n823 585
R419 B.n826 B.n491 585
R420 B.n829 B.n828 585
R421 B.n830 B.n490 585
R422 B.n832 B.n831 585
R423 B.n834 B.n489 585
R424 B.n837 B.n836 585
R425 B.n838 B.n488 585
R426 B.n843 B.n842 585
R427 B.n842 B.n841 585
R428 B.n844 B.n484 585
R429 B.n484 B.n483 585
R430 B.n846 B.n845 585
R431 B.n847 B.n846 585
R432 B.n478 B.n477 585
R433 B.n479 B.n478 585
R434 B.n855 B.n854 585
R435 B.n854 B.n853 585
R436 B.n856 B.n476 585
R437 B.n476 B.n474 585
R438 B.n858 B.n857 585
R439 B.n859 B.n858 585
R440 B.n470 B.n469 585
R441 B.n475 B.n470 585
R442 B.n867 B.n866 585
R443 B.n866 B.n865 585
R444 B.n868 B.n468 585
R445 B.n468 B.n467 585
R446 B.n870 B.n869 585
R447 B.n871 B.n870 585
R448 B.n462 B.n461 585
R449 B.n463 B.n462 585
R450 B.n879 B.n878 585
R451 B.n878 B.n877 585
R452 B.n880 B.n460 585
R453 B.n460 B.n459 585
R454 B.n882 B.n881 585
R455 B.n883 B.n882 585
R456 B.n454 B.n453 585
R457 B.n455 B.n454 585
R458 B.n891 B.n890 585
R459 B.n890 B.n889 585
R460 B.n892 B.n452 585
R461 B.n452 B.n451 585
R462 B.n894 B.n893 585
R463 B.n895 B.n894 585
R464 B.n446 B.n445 585
R465 B.n447 B.n446 585
R466 B.n903 B.n902 585
R467 B.n902 B.n901 585
R468 B.n904 B.n444 585
R469 B.n444 B.n443 585
R470 B.n906 B.n905 585
R471 B.n907 B.n906 585
R472 B.n438 B.n437 585
R473 B.n439 B.n438 585
R474 B.n915 B.n914 585
R475 B.n914 B.n913 585
R476 B.n916 B.n436 585
R477 B.n436 B.n435 585
R478 B.n918 B.n917 585
R479 B.n919 B.n918 585
R480 B.n430 B.n429 585
R481 B.n431 B.n430 585
R482 B.n928 B.n927 585
R483 B.n927 B.n926 585
R484 B.n929 B.n428 585
R485 B.n925 B.n428 585
R486 B.n931 B.n930 585
R487 B.n932 B.n931 585
R488 B.n423 B.n422 585
R489 B.n424 B.n423 585
R490 B.n941 B.n940 585
R491 B.n940 B.n939 585
R492 B.n942 B.n421 585
R493 B.n421 B.n420 585
R494 B.n944 B.n943 585
R495 B.n945 B.n944 585
R496 B.n2 B.n0 585
R497 B.n4 B.n2 585
R498 B.n3 B.n1 585
R499 B.n1069 B.n3 585
R500 B.n1067 B.n1066 585
R501 B.n1068 B.n1067 585
R502 B.n1065 B.n9 585
R503 B.n9 B.n8 585
R504 B.n1064 B.n1063 585
R505 B.n1063 B.n1062 585
R506 B.n11 B.n10 585
R507 B.n1061 B.n11 585
R508 B.n1059 B.n1058 585
R509 B.n1060 B.n1059 585
R510 B.n1057 B.n15 585
R511 B.n18 B.n15 585
R512 B.n1056 B.n1055 585
R513 B.n1055 B.n1054 585
R514 B.n17 B.n16 585
R515 B.n1053 B.n17 585
R516 B.n1051 B.n1050 585
R517 B.n1052 B.n1051 585
R518 B.n1049 B.n23 585
R519 B.n23 B.n22 585
R520 B.n1048 B.n1047 585
R521 B.n1047 B.n1046 585
R522 B.n25 B.n24 585
R523 B.n1045 B.n25 585
R524 B.n1043 B.n1042 585
R525 B.n1044 B.n1043 585
R526 B.n1041 B.n30 585
R527 B.n30 B.n29 585
R528 B.n1040 B.n1039 585
R529 B.n1039 B.n1038 585
R530 B.n32 B.n31 585
R531 B.n1037 B.n32 585
R532 B.n1035 B.n1034 585
R533 B.n1036 B.n1035 585
R534 B.n1033 B.n37 585
R535 B.n37 B.n36 585
R536 B.n1032 B.n1031 585
R537 B.n1031 B.n1030 585
R538 B.n39 B.n38 585
R539 B.n1029 B.n39 585
R540 B.n1027 B.n1026 585
R541 B.n1028 B.n1027 585
R542 B.n1025 B.n44 585
R543 B.n44 B.n43 585
R544 B.n1024 B.n1023 585
R545 B.n1023 B.n1022 585
R546 B.n46 B.n45 585
R547 B.n1021 B.n46 585
R548 B.n1019 B.n1018 585
R549 B.n1020 B.n1019 585
R550 B.n1017 B.n51 585
R551 B.n51 B.n50 585
R552 B.n1016 B.n1015 585
R553 B.n1015 B.n1014 585
R554 B.n53 B.n52 585
R555 B.n1013 B.n53 585
R556 B.n1011 B.n1010 585
R557 B.n1012 B.n1011 585
R558 B.n1009 B.n58 585
R559 B.n58 B.n57 585
R560 B.n1008 B.n1007 585
R561 B.n1007 B.n1006 585
R562 B.n60 B.n59 585
R563 B.n1005 B.n60 585
R564 B.n1003 B.n1002 585
R565 B.n1004 B.n1003 585
R566 B.n1001 B.n65 585
R567 B.n65 B.n64 585
R568 B.n1000 B.n999 585
R569 B.n999 B.n998 585
R570 B.n1072 B.n1071 585
R571 B.n1071 B.n1070 585
R572 B.n842 B.n486 574.183
R573 B.n999 B.n67 574.183
R574 B.n840 B.n488 574.183
R575 B.n996 B.n68 574.183
R576 B.n521 B.t4 376.265
R577 B.n527 B.t12 376.265
R578 B.n142 B.t15 376.265
R579 B.n139 B.t8 376.265
R580 B.n997 B.n137 256.663
R581 B.n997 B.n136 256.663
R582 B.n997 B.n135 256.663
R583 B.n997 B.n134 256.663
R584 B.n997 B.n133 256.663
R585 B.n997 B.n132 256.663
R586 B.n997 B.n131 256.663
R587 B.n997 B.n130 256.663
R588 B.n997 B.n129 256.663
R589 B.n997 B.n128 256.663
R590 B.n997 B.n127 256.663
R591 B.n997 B.n126 256.663
R592 B.n997 B.n125 256.663
R593 B.n997 B.n124 256.663
R594 B.n997 B.n123 256.663
R595 B.n997 B.n122 256.663
R596 B.n997 B.n121 256.663
R597 B.n997 B.n120 256.663
R598 B.n997 B.n119 256.663
R599 B.n997 B.n118 256.663
R600 B.n997 B.n117 256.663
R601 B.n997 B.n116 256.663
R602 B.n997 B.n115 256.663
R603 B.n997 B.n114 256.663
R604 B.n997 B.n113 256.663
R605 B.n997 B.n112 256.663
R606 B.n997 B.n111 256.663
R607 B.n997 B.n110 256.663
R608 B.n997 B.n109 256.663
R609 B.n997 B.n108 256.663
R610 B.n997 B.n107 256.663
R611 B.n997 B.n106 256.663
R612 B.n997 B.n105 256.663
R613 B.n997 B.n104 256.663
R614 B.n997 B.n103 256.663
R615 B.n997 B.n102 256.663
R616 B.n997 B.n101 256.663
R617 B.n997 B.n100 256.663
R618 B.n997 B.n99 256.663
R619 B.n997 B.n98 256.663
R620 B.n997 B.n97 256.663
R621 B.n997 B.n96 256.663
R622 B.n997 B.n95 256.663
R623 B.n997 B.n94 256.663
R624 B.n997 B.n93 256.663
R625 B.n997 B.n92 256.663
R626 B.n997 B.n91 256.663
R627 B.n997 B.n90 256.663
R628 B.n997 B.n89 256.663
R629 B.n997 B.n88 256.663
R630 B.n997 B.n87 256.663
R631 B.n997 B.n86 256.663
R632 B.n997 B.n85 256.663
R633 B.n997 B.n84 256.663
R634 B.n997 B.n83 256.663
R635 B.n997 B.n82 256.663
R636 B.n997 B.n81 256.663
R637 B.n997 B.n80 256.663
R638 B.n997 B.n79 256.663
R639 B.n997 B.n78 256.663
R640 B.n997 B.n77 256.663
R641 B.n997 B.n76 256.663
R642 B.n997 B.n75 256.663
R643 B.n997 B.n74 256.663
R644 B.n997 B.n73 256.663
R645 B.n997 B.n72 256.663
R646 B.n997 B.n71 256.663
R647 B.n997 B.n70 256.663
R648 B.n997 B.n69 256.663
R649 B.n562 B.n487 256.663
R650 B.n568 B.n487 256.663
R651 B.n570 B.n487 256.663
R652 B.n576 B.n487 256.663
R653 B.n578 B.n487 256.663
R654 B.n584 B.n487 256.663
R655 B.n586 B.n487 256.663
R656 B.n592 B.n487 256.663
R657 B.n594 B.n487 256.663
R658 B.n600 B.n487 256.663
R659 B.n602 B.n487 256.663
R660 B.n608 B.n487 256.663
R661 B.n610 B.n487 256.663
R662 B.n616 B.n487 256.663
R663 B.n618 B.n487 256.663
R664 B.n624 B.n487 256.663
R665 B.n626 B.n487 256.663
R666 B.n632 B.n487 256.663
R667 B.n634 B.n487 256.663
R668 B.n640 B.n487 256.663
R669 B.n642 B.n487 256.663
R670 B.n648 B.n487 256.663
R671 B.n650 B.n487 256.663
R672 B.n656 B.n487 256.663
R673 B.n658 B.n487 256.663
R674 B.n664 B.n487 256.663
R675 B.n666 B.n487 256.663
R676 B.n672 B.n487 256.663
R677 B.n674 B.n487 256.663
R678 B.n680 B.n487 256.663
R679 B.n682 B.n487 256.663
R680 B.n688 B.n487 256.663
R681 B.n690 B.n487 256.663
R682 B.n696 B.n487 256.663
R683 B.n698 B.n487 256.663
R684 B.n704 B.n487 256.663
R685 B.n706 B.n487 256.663
R686 B.n713 B.n487 256.663
R687 B.n715 B.n487 256.663
R688 B.n721 B.n487 256.663
R689 B.n723 B.n487 256.663
R690 B.n729 B.n487 256.663
R691 B.n731 B.n487 256.663
R692 B.n737 B.n487 256.663
R693 B.n739 B.n487 256.663
R694 B.n745 B.n487 256.663
R695 B.n747 B.n487 256.663
R696 B.n753 B.n487 256.663
R697 B.n755 B.n487 256.663
R698 B.n761 B.n487 256.663
R699 B.n763 B.n487 256.663
R700 B.n769 B.n487 256.663
R701 B.n771 B.n487 256.663
R702 B.n777 B.n487 256.663
R703 B.n779 B.n487 256.663
R704 B.n785 B.n487 256.663
R705 B.n787 B.n487 256.663
R706 B.n793 B.n487 256.663
R707 B.n795 B.n487 256.663
R708 B.n801 B.n487 256.663
R709 B.n803 B.n487 256.663
R710 B.n809 B.n487 256.663
R711 B.n811 B.n487 256.663
R712 B.n817 B.n487 256.663
R713 B.n819 B.n487 256.663
R714 B.n825 B.n487 256.663
R715 B.n827 B.n487 256.663
R716 B.n833 B.n487 256.663
R717 B.n835 B.n487 256.663
R718 B.n842 B.n484 163.367
R719 B.n846 B.n484 163.367
R720 B.n846 B.n478 163.367
R721 B.n854 B.n478 163.367
R722 B.n854 B.n476 163.367
R723 B.n858 B.n476 163.367
R724 B.n858 B.n470 163.367
R725 B.n866 B.n470 163.367
R726 B.n866 B.n468 163.367
R727 B.n870 B.n468 163.367
R728 B.n870 B.n462 163.367
R729 B.n878 B.n462 163.367
R730 B.n878 B.n460 163.367
R731 B.n882 B.n460 163.367
R732 B.n882 B.n454 163.367
R733 B.n890 B.n454 163.367
R734 B.n890 B.n452 163.367
R735 B.n894 B.n452 163.367
R736 B.n894 B.n446 163.367
R737 B.n902 B.n446 163.367
R738 B.n902 B.n444 163.367
R739 B.n906 B.n444 163.367
R740 B.n906 B.n438 163.367
R741 B.n914 B.n438 163.367
R742 B.n914 B.n436 163.367
R743 B.n918 B.n436 163.367
R744 B.n918 B.n430 163.367
R745 B.n927 B.n430 163.367
R746 B.n927 B.n428 163.367
R747 B.n931 B.n428 163.367
R748 B.n931 B.n423 163.367
R749 B.n940 B.n423 163.367
R750 B.n940 B.n421 163.367
R751 B.n944 B.n421 163.367
R752 B.n944 B.n2 163.367
R753 B.n1071 B.n2 163.367
R754 B.n1071 B.n3 163.367
R755 B.n1067 B.n3 163.367
R756 B.n1067 B.n9 163.367
R757 B.n1063 B.n9 163.367
R758 B.n1063 B.n11 163.367
R759 B.n1059 B.n11 163.367
R760 B.n1059 B.n15 163.367
R761 B.n1055 B.n15 163.367
R762 B.n1055 B.n17 163.367
R763 B.n1051 B.n17 163.367
R764 B.n1051 B.n23 163.367
R765 B.n1047 B.n23 163.367
R766 B.n1047 B.n25 163.367
R767 B.n1043 B.n25 163.367
R768 B.n1043 B.n30 163.367
R769 B.n1039 B.n30 163.367
R770 B.n1039 B.n32 163.367
R771 B.n1035 B.n32 163.367
R772 B.n1035 B.n37 163.367
R773 B.n1031 B.n37 163.367
R774 B.n1031 B.n39 163.367
R775 B.n1027 B.n39 163.367
R776 B.n1027 B.n44 163.367
R777 B.n1023 B.n44 163.367
R778 B.n1023 B.n46 163.367
R779 B.n1019 B.n46 163.367
R780 B.n1019 B.n51 163.367
R781 B.n1015 B.n51 163.367
R782 B.n1015 B.n53 163.367
R783 B.n1011 B.n53 163.367
R784 B.n1011 B.n58 163.367
R785 B.n1007 B.n58 163.367
R786 B.n1007 B.n60 163.367
R787 B.n1003 B.n60 163.367
R788 B.n1003 B.n65 163.367
R789 B.n999 B.n65 163.367
R790 B.n563 B.n561 163.367
R791 B.n567 B.n561 163.367
R792 B.n571 B.n569 163.367
R793 B.n575 B.n559 163.367
R794 B.n579 B.n577 163.367
R795 B.n583 B.n557 163.367
R796 B.n587 B.n585 163.367
R797 B.n591 B.n555 163.367
R798 B.n595 B.n593 163.367
R799 B.n599 B.n553 163.367
R800 B.n603 B.n601 163.367
R801 B.n607 B.n551 163.367
R802 B.n611 B.n609 163.367
R803 B.n615 B.n549 163.367
R804 B.n619 B.n617 163.367
R805 B.n623 B.n547 163.367
R806 B.n627 B.n625 163.367
R807 B.n631 B.n545 163.367
R808 B.n635 B.n633 163.367
R809 B.n639 B.n543 163.367
R810 B.n643 B.n641 163.367
R811 B.n647 B.n541 163.367
R812 B.n651 B.n649 163.367
R813 B.n655 B.n539 163.367
R814 B.n659 B.n657 163.367
R815 B.n663 B.n537 163.367
R816 B.n667 B.n665 163.367
R817 B.n671 B.n535 163.367
R818 B.n675 B.n673 163.367
R819 B.n679 B.n533 163.367
R820 B.n683 B.n681 163.367
R821 B.n687 B.n531 163.367
R822 B.n691 B.n689 163.367
R823 B.n695 B.n526 163.367
R824 B.n699 B.n697 163.367
R825 B.n703 B.n524 163.367
R826 B.n707 B.n705 163.367
R827 B.n712 B.n520 163.367
R828 B.n716 B.n714 163.367
R829 B.n720 B.n518 163.367
R830 B.n724 B.n722 163.367
R831 B.n728 B.n516 163.367
R832 B.n732 B.n730 163.367
R833 B.n736 B.n514 163.367
R834 B.n740 B.n738 163.367
R835 B.n744 B.n512 163.367
R836 B.n748 B.n746 163.367
R837 B.n752 B.n510 163.367
R838 B.n756 B.n754 163.367
R839 B.n760 B.n508 163.367
R840 B.n764 B.n762 163.367
R841 B.n768 B.n506 163.367
R842 B.n772 B.n770 163.367
R843 B.n776 B.n504 163.367
R844 B.n780 B.n778 163.367
R845 B.n784 B.n502 163.367
R846 B.n788 B.n786 163.367
R847 B.n792 B.n500 163.367
R848 B.n796 B.n794 163.367
R849 B.n800 B.n498 163.367
R850 B.n804 B.n802 163.367
R851 B.n808 B.n496 163.367
R852 B.n812 B.n810 163.367
R853 B.n816 B.n494 163.367
R854 B.n820 B.n818 163.367
R855 B.n824 B.n492 163.367
R856 B.n828 B.n826 163.367
R857 B.n832 B.n490 163.367
R858 B.n836 B.n834 163.367
R859 B.n840 B.n482 163.367
R860 B.n848 B.n482 163.367
R861 B.n848 B.n480 163.367
R862 B.n852 B.n480 163.367
R863 B.n852 B.n473 163.367
R864 B.n860 B.n473 163.367
R865 B.n860 B.n471 163.367
R866 B.n864 B.n471 163.367
R867 B.n864 B.n466 163.367
R868 B.n872 B.n466 163.367
R869 B.n872 B.n464 163.367
R870 B.n876 B.n464 163.367
R871 B.n876 B.n458 163.367
R872 B.n884 B.n458 163.367
R873 B.n884 B.n456 163.367
R874 B.n888 B.n456 163.367
R875 B.n888 B.n450 163.367
R876 B.n896 B.n450 163.367
R877 B.n896 B.n448 163.367
R878 B.n900 B.n448 163.367
R879 B.n900 B.n442 163.367
R880 B.n908 B.n442 163.367
R881 B.n908 B.n440 163.367
R882 B.n912 B.n440 163.367
R883 B.n912 B.n434 163.367
R884 B.n920 B.n434 163.367
R885 B.n920 B.n432 163.367
R886 B.n924 B.n432 163.367
R887 B.n924 B.n427 163.367
R888 B.n933 B.n427 163.367
R889 B.n933 B.n425 163.367
R890 B.n938 B.n425 163.367
R891 B.n938 B.n419 163.367
R892 B.n946 B.n419 163.367
R893 B.n947 B.n946 163.367
R894 B.n947 B.n5 163.367
R895 B.n6 B.n5 163.367
R896 B.n7 B.n6 163.367
R897 B.n952 B.n7 163.367
R898 B.n952 B.n12 163.367
R899 B.n13 B.n12 163.367
R900 B.n14 B.n13 163.367
R901 B.n957 B.n14 163.367
R902 B.n957 B.n19 163.367
R903 B.n20 B.n19 163.367
R904 B.n21 B.n20 163.367
R905 B.n962 B.n21 163.367
R906 B.n962 B.n26 163.367
R907 B.n27 B.n26 163.367
R908 B.n28 B.n27 163.367
R909 B.n967 B.n28 163.367
R910 B.n967 B.n33 163.367
R911 B.n34 B.n33 163.367
R912 B.n35 B.n34 163.367
R913 B.n972 B.n35 163.367
R914 B.n972 B.n40 163.367
R915 B.n41 B.n40 163.367
R916 B.n42 B.n41 163.367
R917 B.n977 B.n42 163.367
R918 B.n977 B.n47 163.367
R919 B.n48 B.n47 163.367
R920 B.n49 B.n48 163.367
R921 B.n982 B.n49 163.367
R922 B.n982 B.n54 163.367
R923 B.n55 B.n54 163.367
R924 B.n56 B.n55 163.367
R925 B.n987 B.n56 163.367
R926 B.n987 B.n61 163.367
R927 B.n62 B.n61 163.367
R928 B.n63 B.n62 163.367
R929 B.n992 B.n63 163.367
R930 B.n992 B.n68 163.367
R931 B.n146 B.n145 163.367
R932 B.n150 B.n149 163.367
R933 B.n154 B.n153 163.367
R934 B.n158 B.n157 163.367
R935 B.n162 B.n161 163.367
R936 B.n166 B.n165 163.367
R937 B.n170 B.n169 163.367
R938 B.n174 B.n173 163.367
R939 B.n178 B.n177 163.367
R940 B.n182 B.n181 163.367
R941 B.n186 B.n185 163.367
R942 B.n190 B.n189 163.367
R943 B.n194 B.n193 163.367
R944 B.n198 B.n197 163.367
R945 B.n202 B.n201 163.367
R946 B.n206 B.n205 163.367
R947 B.n210 B.n209 163.367
R948 B.n214 B.n213 163.367
R949 B.n218 B.n217 163.367
R950 B.n222 B.n221 163.367
R951 B.n226 B.n225 163.367
R952 B.n230 B.n229 163.367
R953 B.n234 B.n233 163.367
R954 B.n238 B.n237 163.367
R955 B.n242 B.n241 163.367
R956 B.n246 B.n245 163.367
R957 B.n250 B.n249 163.367
R958 B.n254 B.n253 163.367
R959 B.n258 B.n257 163.367
R960 B.n262 B.n261 163.367
R961 B.n266 B.n265 163.367
R962 B.n270 B.n269 163.367
R963 B.n275 B.n274 163.367
R964 B.n279 B.n278 163.367
R965 B.n283 B.n282 163.367
R966 B.n287 B.n286 163.367
R967 B.n291 B.n290 163.367
R968 B.n295 B.n294 163.367
R969 B.n299 B.n298 163.367
R970 B.n303 B.n302 163.367
R971 B.n307 B.n306 163.367
R972 B.n311 B.n310 163.367
R973 B.n315 B.n314 163.367
R974 B.n319 B.n318 163.367
R975 B.n323 B.n322 163.367
R976 B.n327 B.n326 163.367
R977 B.n331 B.n330 163.367
R978 B.n335 B.n334 163.367
R979 B.n339 B.n338 163.367
R980 B.n343 B.n342 163.367
R981 B.n347 B.n346 163.367
R982 B.n351 B.n350 163.367
R983 B.n355 B.n354 163.367
R984 B.n359 B.n358 163.367
R985 B.n363 B.n362 163.367
R986 B.n367 B.n366 163.367
R987 B.n371 B.n370 163.367
R988 B.n375 B.n374 163.367
R989 B.n379 B.n378 163.367
R990 B.n383 B.n382 163.367
R991 B.n387 B.n386 163.367
R992 B.n391 B.n390 163.367
R993 B.n395 B.n394 163.367
R994 B.n399 B.n398 163.367
R995 B.n403 B.n402 163.367
R996 B.n407 B.n406 163.367
R997 B.n411 B.n410 163.367
R998 B.n415 B.n414 163.367
R999 B.n996 B.n138 163.367
R1000 B.n521 B.t7 132.891
R1001 B.n139 B.t10 132.891
R1002 B.n527 B.t14 132.864
R1003 B.n142 B.t16 132.864
R1004 B.n562 B.n486 71.676
R1005 B.n568 B.n567 71.676
R1006 B.n571 B.n570 71.676
R1007 B.n576 B.n575 71.676
R1008 B.n579 B.n578 71.676
R1009 B.n584 B.n583 71.676
R1010 B.n587 B.n586 71.676
R1011 B.n592 B.n591 71.676
R1012 B.n595 B.n594 71.676
R1013 B.n600 B.n599 71.676
R1014 B.n603 B.n602 71.676
R1015 B.n608 B.n607 71.676
R1016 B.n611 B.n610 71.676
R1017 B.n616 B.n615 71.676
R1018 B.n619 B.n618 71.676
R1019 B.n624 B.n623 71.676
R1020 B.n627 B.n626 71.676
R1021 B.n632 B.n631 71.676
R1022 B.n635 B.n634 71.676
R1023 B.n640 B.n639 71.676
R1024 B.n643 B.n642 71.676
R1025 B.n648 B.n647 71.676
R1026 B.n651 B.n650 71.676
R1027 B.n656 B.n655 71.676
R1028 B.n659 B.n658 71.676
R1029 B.n664 B.n663 71.676
R1030 B.n667 B.n666 71.676
R1031 B.n672 B.n671 71.676
R1032 B.n675 B.n674 71.676
R1033 B.n680 B.n679 71.676
R1034 B.n683 B.n682 71.676
R1035 B.n688 B.n687 71.676
R1036 B.n691 B.n690 71.676
R1037 B.n696 B.n695 71.676
R1038 B.n699 B.n698 71.676
R1039 B.n704 B.n703 71.676
R1040 B.n707 B.n706 71.676
R1041 B.n713 B.n712 71.676
R1042 B.n716 B.n715 71.676
R1043 B.n721 B.n720 71.676
R1044 B.n724 B.n723 71.676
R1045 B.n729 B.n728 71.676
R1046 B.n732 B.n731 71.676
R1047 B.n737 B.n736 71.676
R1048 B.n740 B.n739 71.676
R1049 B.n745 B.n744 71.676
R1050 B.n748 B.n747 71.676
R1051 B.n753 B.n752 71.676
R1052 B.n756 B.n755 71.676
R1053 B.n761 B.n760 71.676
R1054 B.n764 B.n763 71.676
R1055 B.n769 B.n768 71.676
R1056 B.n772 B.n771 71.676
R1057 B.n777 B.n776 71.676
R1058 B.n780 B.n779 71.676
R1059 B.n785 B.n784 71.676
R1060 B.n788 B.n787 71.676
R1061 B.n793 B.n792 71.676
R1062 B.n796 B.n795 71.676
R1063 B.n801 B.n800 71.676
R1064 B.n804 B.n803 71.676
R1065 B.n809 B.n808 71.676
R1066 B.n812 B.n811 71.676
R1067 B.n817 B.n816 71.676
R1068 B.n820 B.n819 71.676
R1069 B.n825 B.n824 71.676
R1070 B.n828 B.n827 71.676
R1071 B.n833 B.n832 71.676
R1072 B.n836 B.n835 71.676
R1073 B.n69 B.n67 71.676
R1074 B.n146 B.n70 71.676
R1075 B.n150 B.n71 71.676
R1076 B.n154 B.n72 71.676
R1077 B.n158 B.n73 71.676
R1078 B.n162 B.n74 71.676
R1079 B.n166 B.n75 71.676
R1080 B.n170 B.n76 71.676
R1081 B.n174 B.n77 71.676
R1082 B.n178 B.n78 71.676
R1083 B.n182 B.n79 71.676
R1084 B.n186 B.n80 71.676
R1085 B.n190 B.n81 71.676
R1086 B.n194 B.n82 71.676
R1087 B.n198 B.n83 71.676
R1088 B.n202 B.n84 71.676
R1089 B.n206 B.n85 71.676
R1090 B.n210 B.n86 71.676
R1091 B.n214 B.n87 71.676
R1092 B.n218 B.n88 71.676
R1093 B.n222 B.n89 71.676
R1094 B.n226 B.n90 71.676
R1095 B.n230 B.n91 71.676
R1096 B.n234 B.n92 71.676
R1097 B.n238 B.n93 71.676
R1098 B.n242 B.n94 71.676
R1099 B.n246 B.n95 71.676
R1100 B.n250 B.n96 71.676
R1101 B.n254 B.n97 71.676
R1102 B.n258 B.n98 71.676
R1103 B.n262 B.n99 71.676
R1104 B.n266 B.n100 71.676
R1105 B.n270 B.n101 71.676
R1106 B.n275 B.n102 71.676
R1107 B.n279 B.n103 71.676
R1108 B.n283 B.n104 71.676
R1109 B.n287 B.n105 71.676
R1110 B.n291 B.n106 71.676
R1111 B.n295 B.n107 71.676
R1112 B.n299 B.n108 71.676
R1113 B.n303 B.n109 71.676
R1114 B.n307 B.n110 71.676
R1115 B.n311 B.n111 71.676
R1116 B.n315 B.n112 71.676
R1117 B.n319 B.n113 71.676
R1118 B.n323 B.n114 71.676
R1119 B.n327 B.n115 71.676
R1120 B.n331 B.n116 71.676
R1121 B.n335 B.n117 71.676
R1122 B.n339 B.n118 71.676
R1123 B.n343 B.n119 71.676
R1124 B.n347 B.n120 71.676
R1125 B.n351 B.n121 71.676
R1126 B.n355 B.n122 71.676
R1127 B.n359 B.n123 71.676
R1128 B.n363 B.n124 71.676
R1129 B.n367 B.n125 71.676
R1130 B.n371 B.n126 71.676
R1131 B.n375 B.n127 71.676
R1132 B.n379 B.n128 71.676
R1133 B.n383 B.n129 71.676
R1134 B.n387 B.n130 71.676
R1135 B.n391 B.n131 71.676
R1136 B.n395 B.n132 71.676
R1137 B.n399 B.n133 71.676
R1138 B.n403 B.n134 71.676
R1139 B.n407 B.n135 71.676
R1140 B.n411 B.n136 71.676
R1141 B.n415 B.n137 71.676
R1142 B.n138 B.n137 71.676
R1143 B.n414 B.n136 71.676
R1144 B.n410 B.n135 71.676
R1145 B.n406 B.n134 71.676
R1146 B.n402 B.n133 71.676
R1147 B.n398 B.n132 71.676
R1148 B.n394 B.n131 71.676
R1149 B.n390 B.n130 71.676
R1150 B.n386 B.n129 71.676
R1151 B.n382 B.n128 71.676
R1152 B.n378 B.n127 71.676
R1153 B.n374 B.n126 71.676
R1154 B.n370 B.n125 71.676
R1155 B.n366 B.n124 71.676
R1156 B.n362 B.n123 71.676
R1157 B.n358 B.n122 71.676
R1158 B.n354 B.n121 71.676
R1159 B.n350 B.n120 71.676
R1160 B.n346 B.n119 71.676
R1161 B.n342 B.n118 71.676
R1162 B.n338 B.n117 71.676
R1163 B.n334 B.n116 71.676
R1164 B.n330 B.n115 71.676
R1165 B.n326 B.n114 71.676
R1166 B.n322 B.n113 71.676
R1167 B.n318 B.n112 71.676
R1168 B.n314 B.n111 71.676
R1169 B.n310 B.n110 71.676
R1170 B.n306 B.n109 71.676
R1171 B.n302 B.n108 71.676
R1172 B.n298 B.n107 71.676
R1173 B.n294 B.n106 71.676
R1174 B.n290 B.n105 71.676
R1175 B.n286 B.n104 71.676
R1176 B.n282 B.n103 71.676
R1177 B.n278 B.n102 71.676
R1178 B.n274 B.n101 71.676
R1179 B.n269 B.n100 71.676
R1180 B.n265 B.n99 71.676
R1181 B.n261 B.n98 71.676
R1182 B.n257 B.n97 71.676
R1183 B.n253 B.n96 71.676
R1184 B.n249 B.n95 71.676
R1185 B.n245 B.n94 71.676
R1186 B.n241 B.n93 71.676
R1187 B.n237 B.n92 71.676
R1188 B.n233 B.n91 71.676
R1189 B.n229 B.n90 71.676
R1190 B.n225 B.n89 71.676
R1191 B.n221 B.n88 71.676
R1192 B.n217 B.n87 71.676
R1193 B.n213 B.n86 71.676
R1194 B.n209 B.n85 71.676
R1195 B.n205 B.n84 71.676
R1196 B.n201 B.n83 71.676
R1197 B.n197 B.n82 71.676
R1198 B.n193 B.n81 71.676
R1199 B.n189 B.n80 71.676
R1200 B.n185 B.n79 71.676
R1201 B.n181 B.n78 71.676
R1202 B.n177 B.n77 71.676
R1203 B.n173 B.n76 71.676
R1204 B.n169 B.n75 71.676
R1205 B.n165 B.n74 71.676
R1206 B.n161 B.n73 71.676
R1207 B.n157 B.n72 71.676
R1208 B.n153 B.n71 71.676
R1209 B.n149 B.n70 71.676
R1210 B.n145 B.n69 71.676
R1211 B.n563 B.n562 71.676
R1212 B.n569 B.n568 71.676
R1213 B.n570 B.n559 71.676
R1214 B.n577 B.n576 71.676
R1215 B.n578 B.n557 71.676
R1216 B.n585 B.n584 71.676
R1217 B.n586 B.n555 71.676
R1218 B.n593 B.n592 71.676
R1219 B.n594 B.n553 71.676
R1220 B.n601 B.n600 71.676
R1221 B.n602 B.n551 71.676
R1222 B.n609 B.n608 71.676
R1223 B.n610 B.n549 71.676
R1224 B.n617 B.n616 71.676
R1225 B.n618 B.n547 71.676
R1226 B.n625 B.n624 71.676
R1227 B.n626 B.n545 71.676
R1228 B.n633 B.n632 71.676
R1229 B.n634 B.n543 71.676
R1230 B.n641 B.n640 71.676
R1231 B.n642 B.n541 71.676
R1232 B.n649 B.n648 71.676
R1233 B.n650 B.n539 71.676
R1234 B.n657 B.n656 71.676
R1235 B.n658 B.n537 71.676
R1236 B.n665 B.n664 71.676
R1237 B.n666 B.n535 71.676
R1238 B.n673 B.n672 71.676
R1239 B.n674 B.n533 71.676
R1240 B.n681 B.n680 71.676
R1241 B.n682 B.n531 71.676
R1242 B.n689 B.n688 71.676
R1243 B.n690 B.n526 71.676
R1244 B.n697 B.n696 71.676
R1245 B.n698 B.n524 71.676
R1246 B.n705 B.n704 71.676
R1247 B.n706 B.n520 71.676
R1248 B.n714 B.n713 71.676
R1249 B.n715 B.n518 71.676
R1250 B.n722 B.n721 71.676
R1251 B.n723 B.n516 71.676
R1252 B.n730 B.n729 71.676
R1253 B.n731 B.n514 71.676
R1254 B.n738 B.n737 71.676
R1255 B.n739 B.n512 71.676
R1256 B.n746 B.n745 71.676
R1257 B.n747 B.n510 71.676
R1258 B.n754 B.n753 71.676
R1259 B.n755 B.n508 71.676
R1260 B.n762 B.n761 71.676
R1261 B.n763 B.n506 71.676
R1262 B.n770 B.n769 71.676
R1263 B.n771 B.n504 71.676
R1264 B.n778 B.n777 71.676
R1265 B.n779 B.n502 71.676
R1266 B.n786 B.n785 71.676
R1267 B.n787 B.n500 71.676
R1268 B.n794 B.n793 71.676
R1269 B.n795 B.n498 71.676
R1270 B.n802 B.n801 71.676
R1271 B.n803 B.n496 71.676
R1272 B.n810 B.n809 71.676
R1273 B.n811 B.n494 71.676
R1274 B.n818 B.n817 71.676
R1275 B.n819 B.n492 71.676
R1276 B.n826 B.n825 71.676
R1277 B.n827 B.n490 71.676
R1278 B.n834 B.n833 71.676
R1279 B.n835 B.n488 71.676
R1280 B.n522 B.t6 71.0241
R1281 B.n140 B.t11 71.0241
R1282 B.n528 B.t13 70.9974
R1283 B.n143 B.t17 70.9974
R1284 B.n522 B.n521 61.8672
R1285 B.n528 B.n527 61.8672
R1286 B.n143 B.n142 61.8672
R1287 B.n140 B.n139 61.8672
R1288 B.n841 B.n487 61.5603
R1289 B.n998 B.n997 61.5603
R1290 B.n709 B.n522 59.5399
R1291 B.n529 B.n528 59.5399
R1292 B.n272 B.n143 59.5399
R1293 B.n141 B.n140 59.5399
R1294 B.n1000 B.n66 37.3078
R1295 B.n995 B.n994 37.3078
R1296 B.n839 B.n838 37.3078
R1297 B.n843 B.n485 37.3078
R1298 B.n841 B.n483 29.6889
R1299 B.n847 B.n483 29.6889
R1300 B.n847 B.n479 29.6889
R1301 B.n853 B.n479 29.6889
R1302 B.n853 B.n474 29.6889
R1303 B.n859 B.n474 29.6889
R1304 B.n859 B.n475 29.6889
R1305 B.n865 B.n467 29.6889
R1306 B.n871 B.n467 29.6889
R1307 B.n871 B.n463 29.6889
R1308 B.n877 B.n463 29.6889
R1309 B.n877 B.n459 29.6889
R1310 B.n883 B.n459 29.6889
R1311 B.n883 B.n455 29.6889
R1312 B.n889 B.n455 29.6889
R1313 B.n889 B.n451 29.6889
R1314 B.n895 B.n451 29.6889
R1315 B.n895 B.n447 29.6889
R1316 B.n901 B.n447 29.6889
R1317 B.n907 B.n443 29.6889
R1318 B.n907 B.n439 29.6889
R1319 B.n913 B.n439 29.6889
R1320 B.n913 B.n435 29.6889
R1321 B.n919 B.n435 29.6889
R1322 B.n919 B.n431 29.6889
R1323 B.n926 B.n431 29.6889
R1324 B.n926 B.n925 29.6889
R1325 B.n932 B.n424 29.6889
R1326 B.n939 B.n424 29.6889
R1327 B.n939 B.n420 29.6889
R1328 B.n945 B.n420 29.6889
R1329 B.n945 B.n4 29.6889
R1330 B.n1070 B.n4 29.6889
R1331 B.n1070 B.n1069 29.6889
R1332 B.n1069 B.n1068 29.6889
R1333 B.n1068 B.n8 29.6889
R1334 B.n1062 B.n8 29.6889
R1335 B.n1062 B.n1061 29.6889
R1336 B.n1061 B.n1060 29.6889
R1337 B.n1054 B.n18 29.6889
R1338 B.n1054 B.n1053 29.6889
R1339 B.n1053 B.n1052 29.6889
R1340 B.n1052 B.n22 29.6889
R1341 B.n1046 B.n22 29.6889
R1342 B.n1046 B.n1045 29.6889
R1343 B.n1045 B.n1044 29.6889
R1344 B.n1044 B.n29 29.6889
R1345 B.n1038 B.n1037 29.6889
R1346 B.n1037 B.n1036 29.6889
R1347 B.n1036 B.n36 29.6889
R1348 B.n1030 B.n36 29.6889
R1349 B.n1030 B.n1029 29.6889
R1350 B.n1029 B.n1028 29.6889
R1351 B.n1028 B.n43 29.6889
R1352 B.n1022 B.n43 29.6889
R1353 B.n1022 B.n1021 29.6889
R1354 B.n1021 B.n1020 29.6889
R1355 B.n1020 B.n50 29.6889
R1356 B.n1014 B.n50 29.6889
R1357 B.n1013 B.n1012 29.6889
R1358 B.n1012 B.n57 29.6889
R1359 B.n1006 B.n57 29.6889
R1360 B.n1006 B.n1005 29.6889
R1361 B.n1005 B.n1004 29.6889
R1362 B.n1004 B.n64 29.6889
R1363 B.n998 B.n64 29.6889
R1364 B.n475 B.t5 21.8302
R1365 B.t9 B.n1013 21.8302
R1366 B.n925 B.t1 20.957
R1367 B.n18 B.t2 20.957
R1368 B.t0 B.n443 20.0838
R1369 B.t3 B.n29 20.0838
R1370 B B.n1072 18.0485
R1371 B.n144 B.n66 10.6151
R1372 B.n147 B.n144 10.6151
R1373 B.n148 B.n147 10.6151
R1374 B.n151 B.n148 10.6151
R1375 B.n152 B.n151 10.6151
R1376 B.n155 B.n152 10.6151
R1377 B.n156 B.n155 10.6151
R1378 B.n159 B.n156 10.6151
R1379 B.n160 B.n159 10.6151
R1380 B.n163 B.n160 10.6151
R1381 B.n164 B.n163 10.6151
R1382 B.n167 B.n164 10.6151
R1383 B.n168 B.n167 10.6151
R1384 B.n171 B.n168 10.6151
R1385 B.n172 B.n171 10.6151
R1386 B.n175 B.n172 10.6151
R1387 B.n176 B.n175 10.6151
R1388 B.n179 B.n176 10.6151
R1389 B.n180 B.n179 10.6151
R1390 B.n183 B.n180 10.6151
R1391 B.n184 B.n183 10.6151
R1392 B.n187 B.n184 10.6151
R1393 B.n188 B.n187 10.6151
R1394 B.n191 B.n188 10.6151
R1395 B.n192 B.n191 10.6151
R1396 B.n195 B.n192 10.6151
R1397 B.n196 B.n195 10.6151
R1398 B.n199 B.n196 10.6151
R1399 B.n200 B.n199 10.6151
R1400 B.n203 B.n200 10.6151
R1401 B.n204 B.n203 10.6151
R1402 B.n207 B.n204 10.6151
R1403 B.n208 B.n207 10.6151
R1404 B.n211 B.n208 10.6151
R1405 B.n212 B.n211 10.6151
R1406 B.n215 B.n212 10.6151
R1407 B.n216 B.n215 10.6151
R1408 B.n219 B.n216 10.6151
R1409 B.n220 B.n219 10.6151
R1410 B.n223 B.n220 10.6151
R1411 B.n224 B.n223 10.6151
R1412 B.n227 B.n224 10.6151
R1413 B.n228 B.n227 10.6151
R1414 B.n231 B.n228 10.6151
R1415 B.n232 B.n231 10.6151
R1416 B.n235 B.n232 10.6151
R1417 B.n236 B.n235 10.6151
R1418 B.n239 B.n236 10.6151
R1419 B.n240 B.n239 10.6151
R1420 B.n243 B.n240 10.6151
R1421 B.n244 B.n243 10.6151
R1422 B.n247 B.n244 10.6151
R1423 B.n248 B.n247 10.6151
R1424 B.n251 B.n248 10.6151
R1425 B.n252 B.n251 10.6151
R1426 B.n255 B.n252 10.6151
R1427 B.n256 B.n255 10.6151
R1428 B.n259 B.n256 10.6151
R1429 B.n260 B.n259 10.6151
R1430 B.n263 B.n260 10.6151
R1431 B.n264 B.n263 10.6151
R1432 B.n267 B.n264 10.6151
R1433 B.n268 B.n267 10.6151
R1434 B.n271 B.n268 10.6151
R1435 B.n276 B.n273 10.6151
R1436 B.n277 B.n276 10.6151
R1437 B.n280 B.n277 10.6151
R1438 B.n281 B.n280 10.6151
R1439 B.n284 B.n281 10.6151
R1440 B.n285 B.n284 10.6151
R1441 B.n288 B.n285 10.6151
R1442 B.n289 B.n288 10.6151
R1443 B.n293 B.n292 10.6151
R1444 B.n296 B.n293 10.6151
R1445 B.n297 B.n296 10.6151
R1446 B.n300 B.n297 10.6151
R1447 B.n301 B.n300 10.6151
R1448 B.n304 B.n301 10.6151
R1449 B.n305 B.n304 10.6151
R1450 B.n308 B.n305 10.6151
R1451 B.n309 B.n308 10.6151
R1452 B.n312 B.n309 10.6151
R1453 B.n313 B.n312 10.6151
R1454 B.n316 B.n313 10.6151
R1455 B.n317 B.n316 10.6151
R1456 B.n320 B.n317 10.6151
R1457 B.n321 B.n320 10.6151
R1458 B.n324 B.n321 10.6151
R1459 B.n325 B.n324 10.6151
R1460 B.n328 B.n325 10.6151
R1461 B.n329 B.n328 10.6151
R1462 B.n332 B.n329 10.6151
R1463 B.n333 B.n332 10.6151
R1464 B.n336 B.n333 10.6151
R1465 B.n337 B.n336 10.6151
R1466 B.n340 B.n337 10.6151
R1467 B.n341 B.n340 10.6151
R1468 B.n344 B.n341 10.6151
R1469 B.n345 B.n344 10.6151
R1470 B.n348 B.n345 10.6151
R1471 B.n349 B.n348 10.6151
R1472 B.n352 B.n349 10.6151
R1473 B.n353 B.n352 10.6151
R1474 B.n356 B.n353 10.6151
R1475 B.n357 B.n356 10.6151
R1476 B.n360 B.n357 10.6151
R1477 B.n361 B.n360 10.6151
R1478 B.n364 B.n361 10.6151
R1479 B.n365 B.n364 10.6151
R1480 B.n368 B.n365 10.6151
R1481 B.n369 B.n368 10.6151
R1482 B.n372 B.n369 10.6151
R1483 B.n373 B.n372 10.6151
R1484 B.n376 B.n373 10.6151
R1485 B.n377 B.n376 10.6151
R1486 B.n380 B.n377 10.6151
R1487 B.n381 B.n380 10.6151
R1488 B.n384 B.n381 10.6151
R1489 B.n385 B.n384 10.6151
R1490 B.n388 B.n385 10.6151
R1491 B.n389 B.n388 10.6151
R1492 B.n392 B.n389 10.6151
R1493 B.n393 B.n392 10.6151
R1494 B.n396 B.n393 10.6151
R1495 B.n397 B.n396 10.6151
R1496 B.n400 B.n397 10.6151
R1497 B.n401 B.n400 10.6151
R1498 B.n404 B.n401 10.6151
R1499 B.n405 B.n404 10.6151
R1500 B.n408 B.n405 10.6151
R1501 B.n409 B.n408 10.6151
R1502 B.n412 B.n409 10.6151
R1503 B.n413 B.n412 10.6151
R1504 B.n416 B.n413 10.6151
R1505 B.n417 B.n416 10.6151
R1506 B.n995 B.n417 10.6151
R1507 B.n839 B.n481 10.6151
R1508 B.n849 B.n481 10.6151
R1509 B.n850 B.n849 10.6151
R1510 B.n851 B.n850 10.6151
R1511 B.n851 B.n472 10.6151
R1512 B.n861 B.n472 10.6151
R1513 B.n862 B.n861 10.6151
R1514 B.n863 B.n862 10.6151
R1515 B.n863 B.n465 10.6151
R1516 B.n873 B.n465 10.6151
R1517 B.n874 B.n873 10.6151
R1518 B.n875 B.n874 10.6151
R1519 B.n875 B.n457 10.6151
R1520 B.n885 B.n457 10.6151
R1521 B.n886 B.n885 10.6151
R1522 B.n887 B.n886 10.6151
R1523 B.n887 B.n449 10.6151
R1524 B.n897 B.n449 10.6151
R1525 B.n898 B.n897 10.6151
R1526 B.n899 B.n898 10.6151
R1527 B.n899 B.n441 10.6151
R1528 B.n909 B.n441 10.6151
R1529 B.n910 B.n909 10.6151
R1530 B.n911 B.n910 10.6151
R1531 B.n911 B.n433 10.6151
R1532 B.n921 B.n433 10.6151
R1533 B.n922 B.n921 10.6151
R1534 B.n923 B.n922 10.6151
R1535 B.n923 B.n426 10.6151
R1536 B.n934 B.n426 10.6151
R1537 B.n935 B.n934 10.6151
R1538 B.n937 B.n935 10.6151
R1539 B.n937 B.n936 10.6151
R1540 B.n936 B.n418 10.6151
R1541 B.n948 B.n418 10.6151
R1542 B.n949 B.n948 10.6151
R1543 B.n950 B.n949 10.6151
R1544 B.n951 B.n950 10.6151
R1545 B.n953 B.n951 10.6151
R1546 B.n954 B.n953 10.6151
R1547 B.n955 B.n954 10.6151
R1548 B.n956 B.n955 10.6151
R1549 B.n958 B.n956 10.6151
R1550 B.n959 B.n958 10.6151
R1551 B.n960 B.n959 10.6151
R1552 B.n961 B.n960 10.6151
R1553 B.n963 B.n961 10.6151
R1554 B.n964 B.n963 10.6151
R1555 B.n965 B.n964 10.6151
R1556 B.n966 B.n965 10.6151
R1557 B.n968 B.n966 10.6151
R1558 B.n969 B.n968 10.6151
R1559 B.n970 B.n969 10.6151
R1560 B.n971 B.n970 10.6151
R1561 B.n973 B.n971 10.6151
R1562 B.n974 B.n973 10.6151
R1563 B.n975 B.n974 10.6151
R1564 B.n976 B.n975 10.6151
R1565 B.n978 B.n976 10.6151
R1566 B.n979 B.n978 10.6151
R1567 B.n980 B.n979 10.6151
R1568 B.n981 B.n980 10.6151
R1569 B.n983 B.n981 10.6151
R1570 B.n984 B.n983 10.6151
R1571 B.n985 B.n984 10.6151
R1572 B.n986 B.n985 10.6151
R1573 B.n988 B.n986 10.6151
R1574 B.n989 B.n988 10.6151
R1575 B.n990 B.n989 10.6151
R1576 B.n991 B.n990 10.6151
R1577 B.n993 B.n991 10.6151
R1578 B.n994 B.n993 10.6151
R1579 B.n564 B.n485 10.6151
R1580 B.n565 B.n564 10.6151
R1581 B.n566 B.n565 10.6151
R1582 B.n566 B.n560 10.6151
R1583 B.n572 B.n560 10.6151
R1584 B.n573 B.n572 10.6151
R1585 B.n574 B.n573 10.6151
R1586 B.n574 B.n558 10.6151
R1587 B.n580 B.n558 10.6151
R1588 B.n581 B.n580 10.6151
R1589 B.n582 B.n581 10.6151
R1590 B.n582 B.n556 10.6151
R1591 B.n588 B.n556 10.6151
R1592 B.n589 B.n588 10.6151
R1593 B.n590 B.n589 10.6151
R1594 B.n590 B.n554 10.6151
R1595 B.n596 B.n554 10.6151
R1596 B.n597 B.n596 10.6151
R1597 B.n598 B.n597 10.6151
R1598 B.n598 B.n552 10.6151
R1599 B.n604 B.n552 10.6151
R1600 B.n605 B.n604 10.6151
R1601 B.n606 B.n605 10.6151
R1602 B.n606 B.n550 10.6151
R1603 B.n612 B.n550 10.6151
R1604 B.n613 B.n612 10.6151
R1605 B.n614 B.n613 10.6151
R1606 B.n614 B.n548 10.6151
R1607 B.n620 B.n548 10.6151
R1608 B.n621 B.n620 10.6151
R1609 B.n622 B.n621 10.6151
R1610 B.n622 B.n546 10.6151
R1611 B.n628 B.n546 10.6151
R1612 B.n629 B.n628 10.6151
R1613 B.n630 B.n629 10.6151
R1614 B.n630 B.n544 10.6151
R1615 B.n636 B.n544 10.6151
R1616 B.n637 B.n636 10.6151
R1617 B.n638 B.n637 10.6151
R1618 B.n638 B.n542 10.6151
R1619 B.n644 B.n542 10.6151
R1620 B.n645 B.n644 10.6151
R1621 B.n646 B.n645 10.6151
R1622 B.n646 B.n540 10.6151
R1623 B.n652 B.n540 10.6151
R1624 B.n653 B.n652 10.6151
R1625 B.n654 B.n653 10.6151
R1626 B.n654 B.n538 10.6151
R1627 B.n660 B.n538 10.6151
R1628 B.n661 B.n660 10.6151
R1629 B.n662 B.n661 10.6151
R1630 B.n662 B.n536 10.6151
R1631 B.n668 B.n536 10.6151
R1632 B.n669 B.n668 10.6151
R1633 B.n670 B.n669 10.6151
R1634 B.n670 B.n534 10.6151
R1635 B.n676 B.n534 10.6151
R1636 B.n677 B.n676 10.6151
R1637 B.n678 B.n677 10.6151
R1638 B.n678 B.n532 10.6151
R1639 B.n684 B.n532 10.6151
R1640 B.n685 B.n684 10.6151
R1641 B.n686 B.n685 10.6151
R1642 B.n686 B.n530 10.6151
R1643 B.n693 B.n692 10.6151
R1644 B.n694 B.n693 10.6151
R1645 B.n694 B.n525 10.6151
R1646 B.n700 B.n525 10.6151
R1647 B.n701 B.n700 10.6151
R1648 B.n702 B.n701 10.6151
R1649 B.n702 B.n523 10.6151
R1650 B.n708 B.n523 10.6151
R1651 B.n711 B.n710 10.6151
R1652 B.n711 B.n519 10.6151
R1653 B.n717 B.n519 10.6151
R1654 B.n718 B.n717 10.6151
R1655 B.n719 B.n718 10.6151
R1656 B.n719 B.n517 10.6151
R1657 B.n725 B.n517 10.6151
R1658 B.n726 B.n725 10.6151
R1659 B.n727 B.n726 10.6151
R1660 B.n727 B.n515 10.6151
R1661 B.n733 B.n515 10.6151
R1662 B.n734 B.n733 10.6151
R1663 B.n735 B.n734 10.6151
R1664 B.n735 B.n513 10.6151
R1665 B.n741 B.n513 10.6151
R1666 B.n742 B.n741 10.6151
R1667 B.n743 B.n742 10.6151
R1668 B.n743 B.n511 10.6151
R1669 B.n749 B.n511 10.6151
R1670 B.n750 B.n749 10.6151
R1671 B.n751 B.n750 10.6151
R1672 B.n751 B.n509 10.6151
R1673 B.n757 B.n509 10.6151
R1674 B.n758 B.n757 10.6151
R1675 B.n759 B.n758 10.6151
R1676 B.n759 B.n507 10.6151
R1677 B.n765 B.n507 10.6151
R1678 B.n766 B.n765 10.6151
R1679 B.n767 B.n766 10.6151
R1680 B.n767 B.n505 10.6151
R1681 B.n773 B.n505 10.6151
R1682 B.n774 B.n773 10.6151
R1683 B.n775 B.n774 10.6151
R1684 B.n775 B.n503 10.6151
R1685 B.n781 B.n503 10.6151
R1686 B.n782 B.n781 10.6151
R1687 B.n783 B.n782 10.6151
R1688 B.n783 B.n501 10.6151
R1689 B.n789 B.n501 10.6151
R1690 B.n790 B.n789 10.6151
R1691 B.n791 B.n790 10.6151
R1692 B.n791 B.n499 10.6151
R1693 B.n797 B.n499 10.6151
R1694 B.n798 B.n797 10.6151
R1695 B.n799 B.n798 10.6151
R1696 B.n799 B.n497 10.6151
R1697 B.n805 B.n497 10.6151
R1698 B.n806 B.n805 10.6151
R1699 B.n807 B.n806 10.6151
R1700 B.n807 B.n495 10.6151
R1701 B.n813 B.n495 10.6151
R1702 B.n814 B.n813 10.6151
R1703 B.n815 B.n814 10.6151
R1704 B.n815 B.n493 10.6151
R1705 B.n821 B.n493 10.6151
R1706 B.n822 B.n821 10.6151
R1707 B.n823 B.n822 10.6151
R1708 B.n823 B.n491 10.6151
R1709 B.n829 B.n491 10.6151
R1710 B.n830 B.n829 10.6151
R1711 B.n831 B.n830 10.6151
R1712 B.n831 B.n489 10.6151
R1713 B.n837 B.n489 10.6151
R1714 B.n838 B.n837 10.6151
R1715 B.n844 B.n843 10.6151
R1716 B.n845 B.n844 10.6151
R1717 B.n845 B.n477 10.6151
R1718 B.n855 B.n477 10.6151
R1719 B.n856 B.n855 10.6151
R1720 B.n857 B.n856 10.6151
R1721 B.n857 B.n469 10.6151
R1722 B.n867 B.n469 10.6151
R1723 B.n868 B.n867 10.6151
R1724 B.n869 B.n868 10.6151
R1725 B.n869 B.n461 10.6151
R1726 B.n879 B.n461 10.6151
R1727 B.n880 B.n879 10.6151
R1728 B.n881 B.n880 10.6151
R1729 B.n881 B.n453 10.6151
R1730 B.n891 B.n453 10.6151
R1731 B.n892 B.n891 10.6151
R1732 B.n893 B.n892 10.6151
R1733 B.n893 B.n445 10.6151
R1734 B.n903 B.n445 10.6151
R1735 B.n904 B.n903 10.6151
R1736 B.n905 B.n904 10.6151
R1737 B.n905 B.n437 10.6151
R1738 B.n915 B.n437 10.6151
R1739 B.n916 B.n915 10.6151
R1740 B.n917 B.n916 10.6151
R1741 B.n917 B.n429 10.6151
R1742 B.n928 B.n429 10.6151
R1743 B.n929 B.n928 10.6151
R1744 B.n930 B.n929 10.6151
R1745 B.n930 B.n422 10.6151
R1746 B.n941 B.n422 10.6151
R1747 B.n942 B.n941 10.6151
R1748 B.n943 B.n942 10.6151
R1749 B.n943 B.n0 10.6151
R1750 B.n1066 B.n1 10.6151
R1751 B.n1066 B.n1065 10.6151
R1752 B.n1065 B.n1064 10.6151
R1753 B.n1064 B.n10 10.6151
R1754 B.n1058 B.n10 10.6151
R1755 B.n1058 B.n1057 10.6151
R1756 B.n1057 B.n1056 10.6151
R1757 B.n1056 B.n16 10.6151
R1758 B.n1050 B.n16 10.6151
R1759 B.n1050 B.n1049 10.6151
R1760 B.n1049 B.n1048 10.6151
R1761 B.n1048 B.n24 10.6151
R1762 B.n1042 B.n24 10.6151
R1763 B.n1042 B.n1041 10.6151
R1764 B.n1041 B.n1040 10.6151
R1765 B.n1040 B.n31 10.6151
R1766 B.n1034 B.n31 10.6151
R1767 B.n1034 B.n1033 10.6151
R1768 B.n1033 B.n1032 10.6151
R1769 B.n1032 B.n38 10.6151
R1770 B.n1026 B.n38 10.6151
R1771 B.n1026 B.n1025 10.6151
R1772 B.n1025 B.n1024 10.6151
R1773 B.n1024 B.n45 10.6151
R1774 B.n1018 B.n45 10.6151
R1775 B.n1018 B.n1017 10.6151
R1776 B.n1017 B.n1016 10.6151
R1777 B.n1016 B.n52 10.6151
R1778 B.n1010 B.n52 10.6151
R1779 B.n1010 B.n1009 10.6151
R1780 B.n1009 B.n1008 10.6151
R1781 B.n1008 B.n59 10.6151
R1782 B.n1002 B.n59 10.6151
R1783 B.n1002 B.n1001 10.6151
R1784 B.n1001 B.n1000 10.6151
R1785 B.n901 B.t0 9.60558
R1786 B.n1038 B.t3 9.60558
R1787 B.n932 B.t1 8.73239
R1788 B.n1060 B.t2 8.73239
R1789 B.n865 B.t5 7.8592
R1790 B.n1014 B.t9 7.8592
R1791 B.n273 B.n272 6.5566
R1792 B.n289 B.n141 6.5566
R1793 B.n692 B.n529 6.5566
R1794 B.n709 B.n708 6.5566
R1795 B.n272 B.n271 4.05904
R1796 B.n292 B.n141 4.05904
R1797 B.n530 B.n529 4.05904
R1798 B.n710 B.n709 4.05904
R1799 B.n1072 B.n0 2.81026
R1800 B.n1072 B.n1 2.81026
R1801 VN.n0 VN.t0 203.27
R1802 VN.n1 VN.t3 203.27
R1803 VN.n0 VN.t1 202.373
R1804 VN.n1 VN.t2 202.373
R1805 VN VN.n1 56.8395
R1806 VN VN.n0 3.43417
R1807 VDD2.n2 VDD2.n0 107.404
R1808 VDD2.n2 VDD2.n1 58.2669
R1809 VDD2.n1 VDD2.t1 0.994476
R1810 VDD2.n1 VDD2.t2 0.994476
R1811 VDD2.n0 VDD2.t3 0.994476
R1812 VDD2.n0 VDD2.t0 0.994476
R1813 VDD2 VDD2.n2 0.0586897
R1814 VTAIL.n6 VTAIL.t2 42.5821
R1815 VTAIL.n5 VTAIL.t1 42.5821
R1816 VTAIL.n4 VTAIL.t4 42.5821
R1817 VTAIL.n3 VTAIL.t5 42.5821
R1818 VTAIL.n7 VTAIL.t6 42.5819
R1819 VTAIL.n0 VTAIL.t7 42.5819
R1820 VTAIL.n1 VTAIL.t3 42.5819
R1821 VTAIL.n2 VTAIL.t0 42.5819
R1822 VTAIL.n7 VTAIL.n6 32.2893
R1823 VTAIL.n3 VTAIL.n2 32.2893
R1824 VTAIL.n4 VTAIL.n3 2.7505
R1825 VTAIL.n6 VTAIL.n5 2.7505
R1826 VTAIL.n2 VTAIL.n1 2.7505
R1827 VTAIL VTAIL.n0 1.43369
R1828 VTAIL VTAIL.n7 1.31731
R1829 VTAIL.n5 VTAIL.n4 0.470328
R1830 VTAIL.n1 VTAIL.n0 0.470328
R1831 VP.n4 VP.t3 203.27
R1832 VP.n4 VP.t2 202.373
R1833 VP.n5 VP.t1 167.857
R1834 VP.n17 VP.t0 167.857
R1835 VP.n16 VP.n0 161.3
R1836 VP.n15 VP.n14 161.3
R1837 VP.n13 VP.n1 161.3
R1838 VP.n12 VP.n11 161.3
R1839 VP.n10 VP.n2 161.3
R1840 VP.n9 VP.n8 161.3
R1841 VP.n7 VP.n3 161.3
R1842 VP.n6 VP.n5 105.981
R1843 VP.n18 VP.n17 105.981
R1844 VP.n6 VP.n4 56.5606
R1845 VP.n11 VP.n10 40.4106
R1846 VP.n11 VP.n1 40.4106
R1847 VP.n9 VP.n3 24.3439
R1848 VP.n10 VP.n9 24.3439
R1849 VP.n15 VP.n1 24.3439
R1850 VP.n16 VP.n15 24.3439
R1851 VP.n5 VP.n3 4.62575
R1852 VP.n17 VP.n16 4.62575
R1853 VP.n7 VP.n6 0.278398
R1854 VP.n18 VP.n0 0.278398
R1855 VP.n8 VP.n7 0.189894
R1856 VP.n8 VP.n2 0.189894
R1857 VP.n12 VP.n2 0.189894
R1858 VP.n13 VP.n12 0.189894
R1859 VP.n14 VP.n13 0.189894
R1860 VP.n14 VP.n0 0.189894
R1861 VP VP.n18 0.153422
R1862 VDD1 VDD1.n1 107.928
R1863 VDD1 VDD1.n0 58.3251
R1864 VDD1.n0 VDD1.t0 0.994476
R1865 VDD1.n0 VDD1.t1 0.994476
R1866 VDD1.n1 VDD1.t2 0.994476
R1867 VDD1.n1 VDD1.t3 0.994476
C0 VDD2 VDD1 1.08517f
C1 VP VTAIL 7.41413f
C2 VTAIL VN 7.40002f
C3 VP VN 7.84734f
C4 VDD1 VTAIL 7.27265f
C5 VDD1 VP 8.07172f
C6 VDD2 VTAIL 7.3286f
C7 VDD2 VP 0.410354f
C8 VDD1 VN 0.148739f
C9 VDD2 VN 7.81091f
C10 VDD2 B 4.53074f
C11 VDD1 B 9.55525f
C12 VTAIL B 15.000439f
C13 VN B 11.835761f
C14 VP B 10.015865f
C15 VDD1.t0 B 0.420907f
C16 VDD1.t1 B 0.420907f
C17 VDD1.n0 B 3.84547f
C18 VDD1.t2 B 0.420907f
C19 VDD1.t3 B 0.420907f
C20 VDD1.n1 B 4.89535f
C21 VP.n0 B 0.029982f
C22 VP.t0 B 3.56991f
C23 VP.n1 B 0.045437f
C24 VP.n2 B 0.02274f
C25 VP.n3 B 0.025559f
C26 VP.t2 B 3.80644f
C27 VP.t3 B 3.81242f
C28 VP.n4 B 3.92992f
C29 VP.t1 B 3.56991f
C30 VP.n5 B 1.30915f
C31 VP.n6 B 1.50148f
C32 VP.n7 B 0.029982f
C33 VP.n8 B 0.02274f
C34 VP.n9 B 0.042594f
C35 VP.n10 B 0.045437f
C36 VP.n11 B 0.018402f
C37 VP.n12 B 0.02274f
C38 VP.n13 B 0.02274f
C39 VP.n14 B 0.02274f
C40 VP.n15 B 0.042594f
C41 VP.n16 B 0.025559f
C42 VP.n17 B 1.30915f
C43 VP.n18 B 0.042079f
C44 VTAIL.t7 B 2.72088f
C45 VTAIL.n0 B 0.311683f
C46 VTAIL.t3 B 2.72088f
C47 VTAIL.n1 B 0.376011f
C48 VTAIL.t0 B 2.72088f
C49 VTAIL.n2 B 1.53222f
C50 VTAIL.t5 B 2.7209f
C51 VTAIL.n3 B 1.53221f
C52 VTAIL.t4 B 2.7209f
C53 VTAIL.n4 B 0.375995f
C54 VTAIL.t1 B 2.7209f
C55 VTAIL.n5 B 0.375995f
C56 VTAIL.t2 B 2.72089f
C57 VTAIL.n6 B 1.53221f
C58 VTAIL.t6 B 2.72088f
C59 VTAIL.n7 B 1.46221f
C60 VDD2.t3 B 0.415371f
C61 VDD2.t0 B 0.415371f
C62 VDD2.n0 B 4.80142f
C63 VDD2.t1 B 0.415371f
C64 VDD2.t2 B 0.415371f
C65 VDD2.n1 B 3.79442f
C66 VDD2.n2 B 4.60317f
C67 VN.t0 B 3.75818f
C68 VN.t1 B 3.75228f
C69 VN.n0 B 2.38753f
C70 VN.t3 B 3.75818f
C71 VN.t2 B 3.75228f
C72 VN.n1 B 3.8857f
.ends

