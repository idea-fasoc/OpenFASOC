* NGSPICE file created from diff_pair_sample_1482.ext - technology: sky130A

.subckt diff_pair_sample_1482 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t11 VN.t0 VDD2.t1 B.t3 sky130_fd_pr__nfet_01v8 ad=0.43725 pd=2.98 as=0.43725 ps=2.98 w=2.65 l=2.81
X1 VTAIL.t3 VP.t0 VDD1.t5 B.t3 sky130_fd_pr__nfet_01v8 ad=0.43725 pd=2.98 as=0.43725 ps=2.98 w=2.65 l=2.81
X2 VDD1.t4 VP.t1 VTAIL.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=1.0335 pd=6.08 as=0.43725 ps=2.98 w=2.65 l=2.81
X3 B.t19 B.t17 B.t18 B.t14 sky130_fd_pr__nfet_01v8 ad=1.0335 pd=6.08 as=0 ps=0 w=2.65 l=2.81
X4 VDD1.t3 VP.t2 VTAIL.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=0.43725 pd=2.98 as=1.0335 ps=6.08 w=2.65 l=2.81
X5 VDD1.t2 VP.t3 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=0.43725 pd=2.98 as=1.0335 ps=6.08 w=2.65 l=2.81
X6 VDD1.t1 VP.t4 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=1.0335 pd=6.08 as=0.43725 ps=2.98 w=2.65 l=2.81
X7 B.t16 B.t13 B.t15 B.t14 sky130_fd_pr__nfet_01v8 ad=1.0335 pd=6.08 as=0 ps=0 w=2.65 l=2.81
X8 B.t12 B.t10 B.t11 B.t7 sky130_fd_pr__nfet_01v8 ad=1.0335 pd=6.08 as=0 ps=0 w=2.65 l=2.81
X9 VTAIL.t2 VP.t5 VDD1.t0 B.t2 sky130_fd_pr__nfet_01v8 ad=0.43725 pd=2.98 as=0.43725 ps=2.98 w=2.65 l=2.81
X10 VDD2.t2 VN.t1 VTAIL.t10 B.t0 sky130_fd_pr__nfet_01v8 ad=0.43725 pd=2.98 as=1.0335 ps=6.08 w=2.65 l=2.81
X11 VTAIL.t9 VN.t2 VDD2.t5 B.t2 sky130_fd_pr__nfet_01v8 ad=0.43725 pd=2.98 as=0.43725 ps=2.98 w=2.65 l=2.81
X12 VDD2.t4 VN.t3 VTAIL.t8 B.t4 sky130_fd_pr__nfet_01v8 ad=1.0335 pd=6.08 as=0.43725 ps=2.98 w=2.65 l=2.81
X13 B.t9 B.t6 B.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=1.0335 pd=6.08 as=0 ps=0 w=2.65 l=2.81
X14 VDD2.t0 VN.t4 VTAIL.t7 B.t1 sky130_fd_pr__nfet_01v8 ad=1.0335 pd=6.08 as=0.43725 ps=2.98 w=2.65 l=2.81
X15 VDD2.t3 VN.t5 VTAIL.t6 B.t5 sky130_fd_pr__nfet_01v8 ad=0.43725 pd=2.98 as=1.0335 ps=6.08 w=2.65 l=2.81
R0 VN.n29 VN.n16 161.3
R1 VN.n28 VN.n27 161.3
R2 VN.n26 VN.n17 161.3
R3 VN.n25 VN.n24 161.3
R4 VN.n23 VN.n18 161.3
R5 VN.n22 VN.n21 161.3
R6 VN.n13 VN.n0 161.3
R7 VN.n12 VN.n11 161.3
R8 VN.n10 VN.n1 161.3
R9 VN.n9 VN.n8 161.3
R10 VN.n7 VN.n2 161.3
R11 VN.n6 VN.n5 161.3
R12 VN.n15 VN.n14 103.906
R13 VN.n31 VN.n30 103.906
R14 VN.n4 VN.t3 57.3801
R15 VN.n20 VN.t1 57.3801
R16 VN.n20 VN.n19 48.9126
R17 VN.n4 VN.n3 48.9126
R18 VN.n8 VN.n1 47.2923
R19 VN.n24 VN.n17 47.2923
R20 VN VN.n31 42.7179
R21 VN.n8 VN.n7 33.6945
R22 VN.n24 VN.n23 33.6945
R23 VN.n6 VN.n3 24.4675
R24 VN.n7 VN.n6 24.4675
R25 VN.n12 VN.n1 24.4675
R26 VN.n13 VN.n12 24.4675
R27 VN.n23 VN.n22 24.4675
R28 VN.n22 VN.n19 24.4675
R29 VN.n29 VN.n28 24.4675
R30 VN.n28 VN.n17 24.4675
R31 VN.n3 VN.t0 22.7283
R32 VN.n14 VN.t5 22.7283
R33 VN.n19 VN.t2 22.7283
R34 VN.n30 VN.t4 22.7283
R35 VN.n14 VN.n13 6.85126
R36 VN.n30 VN.n29 6.85126
R37 VN.n21 VN.n20 4.90017
R38 VN.n5 VN.n4 4.90017
R39 VN.n31 VN.n16 0.278367
R40 VN.n15 VN.n0 0.278367
R41 VN.n27 VN.n16 0.189894
R42 VN.n27 VN.n26 0.189894
R43 VN.n26 VN.n25 0.189894
R44 VN.n25 VN.n18 0.189894
R45 VN.n21 VN.n18 0.189894
R46 VN.n5 VN.n2 0.189894
R47 VN.n9 VN.n2 0.189894
R48 VN.n10 VN.n9 0.189894
R49 VN.n11 VN.n10 0.189894
R50 VN.n11 VN.n0 0.189894
R51 VN VN.n15 0.153454
R52 VDD2.n19 VDD2.n13 289.615
R53 VDD2.n6 VDD2.n0 289.615
R54 VDD2.n20 VDD2.n19 185
R55 VDD2.n18 VDD2.n17 185
R56 VDD2.n5 VDD2.n4 185
R57 VDD2.n7 VDD2.n6 185
R58 VDD2.n3 VDD2.t4 153.582
R59 VDD2.n16 VDD2.t0 153.582
R60 VDD2.n19 VDD2.n18 104.615
R61 VDD2.n6 VDD2.n5 104.615
R62 VDD2.n12 VDD2.n11 84.9062
R63 VDD2 VDD2.n25 84.9033
R64 VDD2.n18 VDD2.t0 52.3082
R65 VDD2.n5 VDD2.t4 52.3082
R66 VDD2.n12 VDD2.n10 48.7056
R67 VDD2.n24 VDD2.n23 46.7308
R68 VDD2.n24 VDD2.n12 34.7972
R69 VDD2.n17 VDD2.n16 10.1164
R70 VDD2.n4 VDD2.n3 10.1164
R71 VDD2.n23 VDD2.n22 9.45567
R72 VDD2.n10 VDD2.n9 9.45567
R73 VDD2.n22 VDD2.n21 9.3005
R74 VDD2.n15 VDD2.n14 9.3005
R75 VDD2.n2 VDD2.n1 9.3005
R76 VDD2.n9 VDD2.n8 9.3005
R77 VDD2.n23 VDD2.n13 8.92171
R78 VDD2.n10 VDD2.n0 8.92171
R79 VDD2.n21 VDD2.n20 8.14595
R80 VDD2.n8 VDD2.n7 8.14595
R81 VDD2.n25 VDD2.t5 7.4722
R82 VDD2.n25 VDD2.t2 7.4722
R83 VDD2.n11 VDD2.t1 7.4722
R84 VDD2.n11 VDD2.t3 7.4722
R85 VDD2.n17 VDD2.n15 7.3702
R86 VDD2.n4 VDD2.n2 7.3702
R87 VDD2.n20 VDD2.n15 5.81868
R88 VDD2.n7 VDD2.n2 5.81868
R89 VDD2.n21 VDD2.n13 5.04292
R90 VDD2.n8 VDD2.n0 5.04292
R91 VDD2.n16 VDD2.n14 3.00987
R92 VDD2.n3 VDD2.n1 3.00987
R93 VDD2 VDD2.n24 2.08886
R94 VDD2.n22 VDD2.n14 0.155672
R95 VDD2.n9 VDD2.n1 0.155672
R96 VTAIL.n50 VTAIL.n44 289.615
R97 VTAIL.n8 VTAIL.n2 289.615
R98 VTAIL.n38 VTAIL.n32 289.615
R99 VTAIL.n24 VTAIL.n18 289.615
R100 VTAIL.n49 VTAIL.n48 185
R101 VTAIL.n51 VTAIL.n50 185
R102 VTAIL.n7 VTAIL.n6 185
R103 VTAIL.n9 VTAIL.n8 185
R104 VTAIL.n39 VTAIL.n38 185
R105 VTAIL.n37 VTAIL.n36 185
R106 VTAIL.n25 VTAIL.n24 185
R107 VTAIL.n23 VTAIL.n22 185
R108 VTAIL.n47 VTAIL.t6 153.582
R109 VTAIL.n5 VTAIL.t0 153.582
R110 VTAIL.n35 VTAIL.t5 153.582
R111 VTAIL.n21 VTAIL.t10 153.582
R112 VTAIL.n50 VTAIL.n49 104.615
R113 VTAIL.n8 VTAIL.n7 104.615
R114 VTAIL.n38 VTAIL.n37 104.615
R115 VTAIL.n24 VTAIL.n23 104.615
R116 VTAIL.n1 VTAIL.n0 67.606
R117 VTAIL.n15 VTAIL.n14 67.606
R118 VTAIL.n31 VTAIL.n30 67.606
R119 VTAIL.n17 VTAIL.n16 67.606
R120 VTAIL.n49 VTAIL.t6 52.3082
R121 VTAIL.n7 VTAIL.t0 52.3082
R122 VTAIL.n37 VTAIL.t5 52.3082
R123 VTAIL.n23 VTAIL.t10 52.3082
R124 VTAIL.n55 VTAIL.n54 30.052
R125 VTAIL.n13 VTAIL.n12 30.052
R126 VTAIL.n43 VTAIL.n42 30.052
R127 VTAIL.n29 VTAIL.n28 30.052
R128 VTAIL.n17 VTAIL.n15 20.0652
R129 VTAIL.n55 VTAIL.n43 17.3583
R130 VTAIL.n48 VTAIL.n47 10.1164
R131 VTAIL.n6 VTAIL.n5 10.1164
R132 VTAIL.n36 VTAIL.n35 10.1164
R133 VTAIL.n22 VTAIL.n21 10.1164
R134 VTAIL.n54 VTAIL.n53 9.45567
R135 VTAIL.n12 VTAIL.n11 9.45567
R136 VTAIL.n42 VTAIL.n41 9.45567
R137 VTAIL.n28 VTAIL.n27 9.45567
R138 VTAIL.n46 VTAIL.n45 9.3005
R139 VTAIL.n53 VTAIL.n52 9.3005
R140 VTAIL.n4 VTAIL.n3 9.3005
R141 VTAIL.n11 VTAIL.n10 9.3005
R142 VTAIL.n34 VTAIL.n33 9.3005
R143 VTAIL.n41 VTAIL.n40 9.3005
R144 VTAIL.n27 VTAIL.n26 9.3005
R145 VTAIL.n20 VTAIL.n19 9.3005
R146 VTAIL.n54 VTAIL.n44 8.92171
R147 VTAIL.n12 VTAIL.n2 8.92171
R148 VTAIL.n42 VTAIL.n32 8.92171
R149 VTAIL.n28 VTAIL.n18 8.92171
R150 VTAIL.n52 VTAIL.n51 8.14595
R151 VTAIL.n10 VTAIL.n9 8.14595
R152 VTAIL.n40 VTAIL.n39 8.14595
R153 VTAIL.n26 VTAIL.n25 8.14595
R154 VTAIL.n0 VTAIL.t8 7.4722
R155 VTAIL.n0 VTAIL.t11 7.4722
R156 VTAIL.n14 VTAIL.t1 7.4722
R157 VTAIL.n14 VTAIL.t2 7.4722
R158 VTAIL.n30 VTAIL.t4 7.4722
R159 VTAIL.n30 VTAIL.t3 7.4722
R160 VTAIL.n16 VTAIL.t7 7.4722
R161 VTAIL.n16 VTAIL.t9 7.4722
R162 VTAIL.n48 VTAIL.n46 7.3702
R163 VTAIL.n6 VTAIL.n4 7.3702
R164 VTAIL.n36 VTAIL.n34 7.3702
R165 VTAIL.n22 VTAIL.n20 7.3702
R166 VTAIL.n51 VTAIL.n46 5.81868
R167 VTAIL.n9 VTAIL.n4 5.81868
R168 VTAIL.n39 VTAIL.n34 5.81868
R169 VTAIL.n25 VTAIL.n20 5.81868
R170 VTAIL.n52 VTAIL.n44 5.04292
R171 VTAIL.n10 VTAIL.n2 5.04292
R172 VTAIL.n40 VTAIL.n32 5.04292
R173 VTAIL.n26 VTAIL.n18 5.04292
R174 VTAIL.n21 VTAIL.n19 3.00987
R175 VTAIL.n47 VTAIL.n45 3.00987
R176 VTAIL.n5 VTAIL.n3 3.00987
R177 VTAIL.n35 VTAIL.n33 3.00987
R178 VTAIL.n29 VTAIL.n17 2.7074
R179 VTAIL.n43 VTAIL.n31 2.7074
R180 VTAIL.n15 VTAIL.n13 2.7074
R181 VTAIL VTAIL.n55 1.97248
R182 VTAIL.n31 VTAIL.n29 1.82378
R183 VTAIL.n13 VTAIL.n1 1.82378
R184 VTAIL VTAIL.n1 0.735414
R185 VTAIL.n53 VTAIL.n45 0.155672
R186 VTAIL.n11 VTAIL.n3 0.155672
R187 VTAIL.n41 VTAIL.n33 0.155672
R188 VTAIL.n27 VTAIL.n19 0.155672
R189 B.n563 B.n562 585
R190 B.n181 B.n102 585
R191 B.n180 B.n179 585
R192 B.n178 B.n177 585
R193 B.n176 B.n175 585
R194 B.n174 B.n173 585
R195 B.n172 B.n171 585
R196 B.n170 B.n169 585
R197 B.n168 B.n167 585
R198 B.n166 B.n165 585
R199 B.n164 B.n163 585
R200 B.n162 B.n161 585
R201 B.n160 B.n159 585
R202 B.n158 B.n157 585
R203 B.n156 B.n155 585
R204 B.n154 B.n153 585
R205 B.n152 B.n151 585
R206 B.n150 B.n149 585
R207 B.n148 B.n147 585
R208 B.n146 B.n145 585
R209 B.n144 B.n143 585
R210 B.n142 B.n141 585
R211 B.n140 B.n139 585
R212 B.n138 B.n137 585
R213 B.n136 B.n135 585
R214 B.n134 B.n133 585
R215 B.n132 B.n131 585
R216 B.n130 B.n129 585
R217 B.n128 B.n127 585
R218 B.n126 B.n125 585
R219 B.n124 B.n123 585
R220 B.n122 B.n121 585
R221 B.n120 B.n119 585
R222 B.n118 B.n117 585
R223 B.n116 B.n115 585
R224 B.n114 B.n113 585
R225 B.n112 B.n111 585
R226 B.n110 B.n109 585
R227 B.n561 B.n83 585
R228 B.n566 B.n83 585
R229 B.n560 B.n82 585
R230 B.n567 B.n82 585
R231 B.n559 B.n558 585
R232 B.n558 B.n78 585
R233 B.n557 B.n77 585
R234 B.n573 B.n77 585
R235 B.n556 B.n76 585
R236 B.n574 B.n76 585
R237 B.n555 B.n75 585
R238 B.n575 B.n75 585
R239 B.n554 B.n553 585
R240 B.n553 B.n71 585
R241 B.n552 B.n70 585
R242 B.n581 B.n70 585
R243 B.n551 B.n69 585
R244 B.n582 B.n69 585
R245 B.n550 B.n68 585
R246 B.n583 B.n68 585
R247 B.n549 B.n548 585
R248 B.n548 B.n64 585
R249 B.n547 B.n63 585
R250 B.n589 B.n63 585
R251 B.n546 B.n62 585
R252 B.n590 B.n62 585
R253 B.n545 B.n61 585
R254 B.n591 B.n61 585
R255 B.n544 B.n543 585
R256 B.n543 B.n57 585
R257 B.n542 B.n56 585
R258 B.n597 B.n56 585
R259 B.n541 B.n55 585
R260 B.n598 B.n55 585
R261 B.n540 B.n54 585
R262 B.n599 B.n54 585
R263 B.n539 B.n538 585
R264 B.n538 B.n50 585
R265 B.n537 B.n49 585
R266 B.n605 B.n49 585
R267 B.n536 B.n48 585
R268 B.n606 B.n48 585
R269 B.n535 B.n47 585
R270 B.n607 B.n47 585
R271 B.n534 B.n533 585
R272 B.n533 B.n43 585
R273 B.n532 B.n42 585
R274 B.n613 B.n42 585
R275 B.n531 B.n41 585
R276 B.n614 B.n41 585
R277 B.n530 B.n40 585
R278 B.n615 B.n40 585
R279 B.n529 B.n528 585
R280 B.n528 B.n36 585
R281 B.n527 B.n35 585
R282 B.n621 B.n35 585
R283 B.n526 B.n34 585
R284 B.n622 B.n34 585
R285 B.n525 B.n33 585
R286 B.n623 B.n33 585
R287 B.n524 B.n523 585
R288 B.n523 B.n29 585
R289 B.n522 B.n28 585
R290 B.n629 B.n28 585
R291 B.n521 B.n27 585
R292 B.n630 B.n27 585
R293 B.n520 B.n26 585
R294 B.n631 B.n26 585
R295 B.n519 B.n518 585
R296 B.n518 B.n22 585
R297 B.n517 B.n21 585
R298 B.n637 B.n21 585
R299 B.n516 B.n20 585
R300 B.n638 B.n20 585
R301 B.n515 B.n19 585
R302 B.n639 B.n19 585
R303 B.n514 B.n513 585
R304 B.n513 B.n18 585
R305 B.n512 B.n14 585
R306 B.n645 B.n14 585
R307 B.n511 B.n13 585
R308 B.n646 B.n13 585
R309 B.n510 B.n12 585
R310 B.n647 B.n12 585
R311 B.n509 B.n508 585
R312 B.n508 B.n8 585
R313 B.n507 B.n7 585
R314 B.n653 B.n7 585
R315 B.n506 B.n6 585
R316 B.n654 B.n6 585
R317 B.n505 B.n5 585
R318 B.n655 B.n5 585
R319 B.n504 B.n503 585
R320 B.n503 B.n4 585
R321 B.n502 B.n182 585
R322 B.n502 B.n501 585
R323 B.n492 B.n183 585
R324 B.n184 B.n183 585
R325 B.n494 B.n493 585
R326 B.n495 B.n494 585
R327 B.n491 B.n189 585
R328 B.n189 B.n188 585
R329 B.n490 B.n489 585
R330 B.n489 B.n488 585
R331 B.n191 B.n190 585
R332 B.n481 B.n191 585
R333 B.n480 B.n479 585
R334 B.n482 B.n480 585
R335 B.n478 B.n196 585
R336 B.n196 B.n195 585
R337 B.n477 B.n476 585
R338 B.n476 B.n475 585
R339 B.n198 B.n197 585
R340 B.n199 B.n198 585
R341 B.n468 B.n467 585
R342 B.n469 B.n468 585
R343 B.n466 B.n204 585
R344 B.n204 B.n203 585
R345 B.n465 B.n464 585
R346 B.n464 B.n463 585
R347 B.n206 B.n205 585
R348 B.n207 B.n206 585
R349 B.n456 B.n455 585
R350 B.n457 B.n456 585
R351 B.n454 B.n212 585
R352 B.n212 B.n211 585
R353 B.n453 B.n452 585
R354 B.n452 B.n451 585
R355 B.n214 B.n213 585
R356 B.n215 B.n214 585
R357 B.n444 B.n443 585
R358 B.n445 B.n444 585
R359 B.n442 B.n220 585
R360 B.n220 B.n219 585
R361 B.n441 B.n440 585
R362 B.n440 B.n439 585
R363 B.n222 B.n221 585
R364 B.n223 B.n222 585
R365 B.n432 B.n431 585
R366 B.n433 B.n432 585
R367 B.n430 B.n227 585
R368 B.n231 B.n227 585
R369 B.n429 B.n428 585
R370 B.n428 B.n427 585
R371 B.n229 B.n228 585
R372 B.n230 B.n229 585
R373 B.n420 B.n419 585
R374 B.n421 B.n420 585
R375 B.n418 B.n236 585
R376 B.n236 B.n235 585
R377 B.n417 B.n416 585
R378 B.n416 B.n415 585
R379 B.n238 B.n237 585
R380 B.n239 B.n238 585
R381 B.n408 B.n407 585
R382 B.n409 B.n408 585
R383 B.n406 B.n244 585
R384 B.n244 B.n243 585
R385 B.n405 B.n404 585
R386 B.n404 B.n403 585
R387 B.n246 B.n245 585
R388 B.n247 B.n246 585
R389 B.n396 B.n395 585
R390 B.n397 B.n396 585
R391 B.n394 B.n252 585
R392 B.n252 B.n251 585
R393 B.n393 B.n392 585
R394 B.n392 B.n391 585
R395 B.n254 B.n253 585
R396 B.n255 B.n254 585
R397 B.n384 B.n383 585
R398 B.n385 B.n384 585
R399 B.n382 B.n260 585
R400 B.n260 B.n259 585
R401 B.n381 B.n380 585
R402 B.n380 B.n379 585
R403 B.n262 B.n261 585
R404 B.n263 B.n262 585
R405 B.n372 B.n371 585
R406 B.n373 B.n372 585
R407 B.n370 B.n268 585
R408 B.n268 B.n267 585
R409 B.n365 B.n364 585
R410 B.n363 B.n289 585
R411 B.n362 B.n288 585
R412 B.n367 B.n288 585
R413 B.n361 B.n360 585
R414 B.n359 B.n358 585
R415 B.n357 B.n356 585
R416 B.n355 B.n354 585
R417 B.n353 B.n352 585
R418 B.n351 B.n350 585
R419 B.n349 B.n348 585
R420 B.n347 B.n346 585
R421 B.n345 B.n344 585
R422 B.n343 B.n342 585
R423 B.n341 B.n340 585
R424 B.n338 B.n337 585
R425 B.n336 B.n335 585
R426 B.n334 B.n333 585
R427 B.n332 B.n331 585
R428 B.n330 B.n329 585
R429 B.n328 B.n327 585
R430 B.n326 B.n325 585
R431 B.n324 B.n323 585
R432 B.n322 B.n321 585
R433 B.n320 B.n319 585
R434 B.n317 B.n316 585
R435 B.n315 B.n314 585
R436 B.n313 B.n312 585
R437 B.n311 B.n310 585
R438 B.n309 B.n308 585
R439 B.n307 B.n306 585
R440 B.n305 B.n304 585
R441 B.n303 B.n302 585
R442 B.n301 B.n300 585
R443 B.n299 B.n298 585
R444 B.n297 B.n296 585
R445 B.n295 B.n294 585
R446 B.n270 B.n269 585
R447 B.n369 B.n368 585
R448 B.n368 B.n367 585
R449 B.n266 B.n265 585
R450 B.n267 B.n266 585
R451 B.n375 B.n374 585
R452 B.n374 B.n373 585
R453 B.n376 B.n264 585
R454 B.n264 B.n263 585
R455 B.n378 B.n377 585
R456 B.n379 B.n378 585
R457 B.n258 B.n257 585
R458 B.n259 B.n258 585
R459 B.n387 B.n386 585
R460 B.n386 B.n385 585
R461 B.n388 B.n256 585
R462 B.n256 B.n255 585
R463 B.n390 B.n389 585
R464 B.n391 B.n390 585
R465 B.n250 B.n249 585
R466 B.n251 B.n250 585
R467 B.n399 B.n398 585
R468 B.n398 B.n397 585
R469 B.n400 B.n248 585
R470 B.n248 B.n247 585
R471 B.n402 B.n401 585
R472 B.n403 B.n402 585
R473 B.n242 B.n241 585
R474 B.n243 B.n242 585
R475 B.n411 B.n410 585
R476 B.n410 B.n409 585
R477 B.n412 B.n240 585
R478 B.n240 B.n239 585
R479 B.n414 B.n413 585
R480 B.n415 B.n414 585
R481 B.n234 B.n233 585
R482 B.n235 B.n234 585
R483 B.n423 B.n422 585
R484 B.n422 B.n421 585
R485 B.n424 B.n232 585
R486 B.n232 B.n230 585
R487 B.n426 B.n425 585
R488 B.n427 B.n426 585
R489 B.n226 B.n225 585
R490 B.n231 B.n226 585
R491 B.n435 B.n434 585
R492 B.n434 B.n433 585
R493 B.n436 B.n224 585
R494 B.n224 B.n223 585
R495 B.n438 B.n437 585
R496 B.n439 B.n438 585
R497 B.n218 B.n217 585
R498 B.n219 B.n218 585
R499 B.n447 B.n446 585
R500 B.n446 B.n445 585
R501 B.n448 B.n216 585
R502 B.n216 B.n215 585
R503 B.n450 B.n449 585
R504 B.n451 B.n450 585
R505 B.n210 B.n209 585
R506 B.n211 B.n210 585
R507 B.n459 B.n458 585
R508 B.n458 B.n457 585
R509 B.n460 B.n208 585
R510 B.n208 B.n207 585
R511 B.n462 B.n461 585
R512 B.n463 B.n462 585
R513 B.n202 B.n201 585
R514 B.n203 B.n202 585
R515 B.n471 B.n470 585
R516 B.n470 B.n469 585
R517 B.n472 B.n200 585
R518 B.n200 B.n199 585
R519 B.n474 B.n473 585
R520 B.n475 B.n474 585
R521 B.n194 B.n193 585
R522 B.n195 B.n194 585
R523 B.n484 B.n483 585
R524 B.n483 B.n482 585
R525 B.n485 B.n192 585
R526 B.n481 B.n192 585
R527 B.n487 B.n486 585
R528 B.n488 B.n487 585
R529 B.n187 B.n186 585
R530 B.n188 B.n187 585
R531 B.n497 B.n496 585
R532 B.n496 B.n495 585
R533 B.n498 B.n185 585
R534 B.n185 B.n184 585
R535 B.n500 B.n499 585
R536 B.n501 B.n500 585
R537 B.n2 B.n0 585
R538 B.n4 B.n2 585
R539 B.n3 B.n1 585
R540 B.n654 B.n3 585
R541 B.n652 B.n651 585
R542 B.n653 B.n652 585
R543 B.n650 B.n9 585
R544 B.n9 B.n8 585
R545 B.n649 B.n648 585
R546 B.n648 B.n647 585
R547 B.n11 B.n10 585
R548 B.n646 B.n11 585
R549 B.n644 B.n643 585
R550 B.n645 B.n644 585
R551 B.n642 B.n15 585
R552 B.n18 B.n15 585
R553 B.n641 B.n640 585
R554 B.n640 B.n639 585
R555 B.n17 B.n16 585
R556 B.n638 B.n17 585
R557 B.n636 B.n635 585
R558 B.n637 B.n636 585
R559 B.n634 B.n23 585
R560 B.n23 B.n22 585
R561 B.n633 B.n632 585
R562 B.n632 B.n631 585
R563 B.n25 B.n24 585
R564 B.n630 B.n25 585
R565 B.n628 B.n627 585
R566 B.n629 B.n628 585
R567 B.n626 B.n30 585
R568 B.n30 B.n29 585
R569 B.n625 B.n624 585
R570 B.n624 B.n623 585
R571 B.n32 B.n31 585
R572 B.n622 B.n32 585
R573 B.n620 B.n619 585
R574 B.n621 B.n620 585
R575 B.n618 B.n37 585
R576 B.n37 B.n36 585
R577 B.n617 B.n616 585
R578 B.n616 B.n615 585
R579 B.n39 B.n38 585
R580 B.n614 B.n39 585
R581 B.n612 B.n611 585
R582 B.n613 B.n612 585
R583 B.n610 B.n44 585
R584 B.n44 B.n43 585
R585 B.n609 B.n608 585
R586 B.n608 B.n607 585
R587 B.n46 B.n45 585
R588 B.n606 B.n46 585
R589 B.n604 B.n603 585
R590 B.n605 B.n604 585
R591 B.n602 B.n51 585
R592 B.n51 B.n50 585
R593 B.n601 B.n600 585
R594 B.n600 B.n599 585
R595 B.n53 B.n52 585
R596 B.n598 B.n53 585
R597 B.n596 B.n595 585
R598 B.n597 B.n596 585
R599 B.n594 B.n58 585
R600 B.n58 B.n57 585
R601 B.n593 B.n592 585
R602 B.n592 B.n591 585
R603 B.n60 B.n59 585
R604 B.n590 B.n60 585
R605 B.n588 B.n587 585
R606 B.n589 B.n588 585
R607 B.n586 B.n65 585
R608 B.n65 B.n64 585
R609 B.n585 B.n584 585
R610 B.n584 B.n583 585
R611 B.n67 B.n66 585
R612 B.n582 B.n67 585
R613 B.n580 B.n579 585
R614 B.n581 B.n580 585
R615 B.n578 B.n72 585
R616 B.n72 B.n71 585
R617 B.n577 B.n576 585
R618 B.n576 B.n575 585
R619 B.n74 B.n73 585
R620 B.n574 B.n74 585
R621 B.n572 B.n571 585
R622 B.n573 B.n572 585
R623 B.n570 B.n79 585
R624 B.n79 B.n78 585
R625 B.n569 B.n568 585
R626 B.n568 B.n567 585
R627 B.n81 B.n80 585
R628 B.n566 B.n81 585
R629 B.n657 B.n656 585
R630 B.n656 B.n655 585
R631 B.n365 B.n266 492.5
R632 B.n109 B.n81 492.5
R633 B.n368 B.n268 492.5
R634 B.n563 B.n83 492.5
R635 B.n565 B.n564 256.663
R636 B.n565 B.n101 256.663
R637 B.n565 B.n100 256.663
R638 B.n565 B.n99 256.663
R639 B.n565 B.n98 256.663
R640 B.n565 B.n97 256.663
R641 B.n565 B.n96 256.663
R642 B.n565 B.n95 256.663
R643 B.n565 B.n94 256.663
R644 B.n565 B.n93 256.663
R645 B.n565 B.n92 256.663
R646 B.n565 B.n91 256.663
R647 B.n565 B.n90 256.663
R648 B.n565 B.n89 256.663
R649 B.n565 B.n88 256.663
R650 B.n565 B.n87 256.663
R651 B.n565 B.n86 256.663
R652 B.n565 B.n85 256.663
R653 B.n565 B.n84 256.663
R654 B.n367 B.n366 256.663
R655 B.n367 B.n271 256.663
R656 B.n367 B.n272 256.663
R657 B.n367 B.n273 256.663
R658 B.n367 B.n274 256.663
R659 B.n367 B.n275 256.663
R660 B.n367 B.n276 256.663
R661 B.n367 B.n277 256.663
R662 B.n367 B.n278 256.663
R663 B.n367 B.n279 256.663
R664 B.n367 B.n280 256.663
R665 B.n367 B.n281 256.663
R666 B.n367 B.n282 256.663
R667 B.n367 B.n283 256.663
R668 B.n367 B.n284 256.663
R669 B.n367 B.n285 256.663
R670 B.n367 B.n286 256.663
R671 B.n367 B.n287 256.663
R672 B.n292 B.t17 231.071
R673 B.n290 B.t13 231.071
R674 B.n106 B.t6 231.071
R675 B.n103 B.t10 231.071
R676 B.n292 B.t19 186.506
R677 B.n103 B.t11 186.506
R678 B.n290 B.t16 186.506
R679 B.n106 B.t8 186.506
R680 B.n367 B.n267 176.279
R681 B.n566 B.n565 176.279
R682 B.n374 B.n266 163.367
R683 B.n374 B.n264 163.367
R684 B.n378 B.n264 163.367
R685 B.n378 B.n258 163.367
R686 B.n386 B.n258 163.367
R687 B.n386 B.n256 163.367
R688 B.n390 B.n256 163.367
R689 B.n390 B.n250 163.367
R690 B.n398 B.n250 163.367
R691 B.n398 B.n248 163.367
R692 B.n402 B.n248 163.367
R693 B.n402 B.n242 163.367
R694 B.n410 B.n242 163.367
R695 B.n410 B.n240 163.367
R696 B.n414 B.n240 163.367
R697 B.n414 B.n234 163.367
R698 B.n422 B.n234 163.367
R699 B.n422 B.n232 163.367
R700 B.n426 B.n232 163.367
R701 B.n426 B.n226 163.367
R702 B.n434 B.n226 163.367
R703 B.n434 B.n224 163.367
R704 B.n438 B.n224 163.367
R705 B.n438 B.n218 163.367
R706 B.n446 B.n218 163.367
R707 B.n446 B.n216 163.367
R708 B.n450 B.n216 163.367
R709 B.n450 B.n210 163.367
R710 B.n458 B.n210 163.367
R711 B.n458 B.n208 163.367
R712 B.n462 B.n208 163.367
R713 B.n462 B.n202 163.367
R714 B.n470 B.n202 163.367
R715 B.n470 B.n200 163.367
R716 B.n474 B.n200 163.367
R717 B.n474 B.n194 163.367
R718 B.n483 B.n194 163.367
R719 B.n483 B.n192 163.367
R720 B.n487 B.n192 163.367
R721 B.n487 B.n187 163.367
R722 B.n496 B.n187 163.367
R723 B.n496 B.n185 163.367
R724 B.n500 B.n185 163.367
R725 B.n500 B.n2 163.367
R726 B.n656 B.n2 163.367
R727 B.n656 B.n3 163.367
R728 B.n652 B.n3 163.367
R729 B.n652 B.n9 163.367
R730 B.n648 B.n9 163.367
R731 B.n648 B.n11 163.367
R732 B.n644 B.n11 163.367
R733 B.n644 B.n15 163.367
R734 B.n640 B.n15 163.367
R735 B.n640 B.n17 163.367
R736 B.n636 B.n17 163.367
R737 B.n636 B.n23 163.367
R738 B.n632 B.n23 163.367
R739 B.n632 B.n25 163.367
R740 B.n628 B.n25 163.367
R741 B.n628 B.n30 163.367
R742 B.n624 B.n30 163.367
R743 B.n624 B.n32 163.367
R744 B.n620 B.n32 163.367
R745 B.n620 B.n37 163.367
R746 B.n616 B.n37 163.367
R747 B.n616 B.n39 163.367
R748 B.n612 B.n39 163.367
R749 B.n612 B.n44 163.367
R750 B.n608 B.n44 163.367
R751 B.n608 B.n46 163.367
R752 B.n604 B.n46 163.367
R753 B.n604 B.n51 163.367
R754 B.n600 B.n51 163.367
R755 B.n600 B.n53 163.367
R756 B.n596 B.n53 163.367
R757 B.n596 B.n58 163.367
R758 B.n592 B.n58 163.367
R759 B.n592 B.n60 163.367
R760 B.n588 B.n60 163.367
R761 B.n588 B.n65 163.367
R762 B.n584 B.n65 163.367
R763 B.n584 B.n67 163.367
R764 B.n580 B.n67 163.367
R765 B.n580 B.n72 163.367
R766 B.n576 B.n72 163.367
R767 B.n576 B.n74 163.367
R768 B.n572 B.n74 163.367
R769 B.n572 B.n79 163.367
R770 B.n568 B.n79 163.367
R771 B.n568 B.n81 163.367
R772 B.n289 B.n288 163.367
R773 B.n360 B.n288 163.367
R774 B.n358 B.n357 163.367
R775 B.n354 B.n353 163.367
R776 B.n350 B.n349 163.367
R777 B.n346 B.n345 163.367
R778 B.n342 B.n341 163.367
R779 B.n337 B.n336 163.367
R780 B.n333 B.n332 163.367
R781 B.n329 B.n328 163.367
R782 B.n325 B.n324 163.367
R783 B.n321 B.n320 163.367
R784 B.n316 B.n315 163.367
R785 B.n312 B.n311 163.367
R786 B.n308 B.n307 163.367
R787 B.n304 B.n303 163.367
R788 B.n300 B.n299 163.367
R789 B.n296 B.n295 163.367
R790 B.n368 B.n270 163.367
R791 B.n372 B.n268 163.367
R792 B.n372 B.n262 163.367
R793 B.n380 B.n262 163.367
R794 B.n380 B.n260 163.367
R795 B.n384 B.n260 163.367
R796 B.n384 B.n254 163.367
R797 B.n392 B.n254 163.367
R798 B.n392 B.n252 163.367
R799 B.n396 B.n252 163.367
R800 B.n396 B.n246 163.367
R801 B.n404 B.n246 163.367
R802 B.n404 B.n244 163.367
R803 B.n408 B.n244 163.367
R804 B.n408 B.n238 163.367
R805 B.n416 B.n238 163.367
R806 B.n416 B.n236 163.367
R807 B.n420 B.n236 163.367
R808 B.n420 B.n229 163.367
R809 B.n428 B.n229 163.367
R810 B.n428 B.n227 163.367
R811 B.n432 B.n227 163.367
R812 B.n432 B.n222 163.367
R813 B.n440 B.n222 163.367
R814 B.n440 B.n220 163.367
R815 B.n444 B.n220 163.367
R816 B.n444 B.n214 163.367
R817 B.n452 B.n214 163.367
R818 B.n452 B.n212 163.367
R819 B.n456 B.n212 163.367
R820 B.n456 B.n206 163.367
R821 B.n464 B.n206 163.367
R822 B.n464 B.n204 163.367
R823 B.n468 B.n204 163.367
R824 B.n468 B.n198 163.367
R825 B.n476 B.n198 163.367
R826 B.n476 B.n196 163.367
R827 B.n480 B.n196 163.367
R828 B.n480 B.n191 163.367
R829 B.n489 B.n191 163.367
R830 B.n489 B.n189 163.367
R831 B.n494 B.n189 163.367
R832 B.n494 B.n183 163.367
R833 B.n502 B.n183 163.367
R834 B.n503 B.n502 163.367
R835 B.n503 B.n5 163.367
R836 B.n6 B.n5 163.367
R837 B.n7 B.n6 163.367
R838 B.n508 B.n7 163.367
R839 B.n508 B.n12 163.367
R840 B.n13 B.n12 163.367
R841 B.n14 B.n13 163.367
R842 B.n513 B.n14 163.367
R843 B.n513 B.n19 163.367
R844 B.n20 B.n19 163.367
R845 B.n21 B.n20 163.367
R846 B.n518 B.n21 163.367
R847 B.n518 B.n26 163.367
R848 B.n27 B.n26 163.367
R849 B.n28 B.n27 163.367
R850 B.n523 B.n28 163.367
R851 B.n523 B.n33 163.367
R852 B.n34 B.n33 163.367
R853 B.n35 B.n34 163.367
R854 B.n528 B.n35 163.367
R855 B.n528 B.n40 163.367
R856 B.n41 B.n40 163.367
R857 B.n42 B.n41 163.367
R858 B.n533 B.n42 163.367
R859 B.n533 B.n47 163.367
R860 B.n48 B.n47 163.367
R861 B.n49 B.n48 163.367
R862 B.n538 B.n49 163.367
R863 B.n538 B.n54 163.367
R864 B.n55 B.n54 163.367
R865 B.n56 B.n55 163.367
R866 B.n543 B.n56 163.367
R867 B.n543 B.n61 163.367
R868 B.n62 B.n61 163.367
R869 B.n63 B.n62 163.367
R870 B.n548 B.n63 163.367
R871 B.n548 B.n68 163.367
R872 B.n69 B.n68 163.367
R873 B.n70 B.n69 163.367
R874 B.n553 B.n70 163.367
R875 B.n553 B.n75 163.367
R876 B.n76 B.n75 163.367
R877 B.n77 B.n76 163.367
R878 B.n558 B.n77 163.367
R879 B.n558 B.n82 163.367
R880 B.n83 B.n82 163.367
R881 B.n113 B.n112 163.367
R882 B.n117 B.n116 163.367
R883 B.n121 B.n120 163.367
R884 B.n125 B.n124 163.367
R885 B.n129 B.n128 163.367
R886 B.n133 B.n132 163.367
R887 B.n137 B.n136 163.367
R888 B.n141 B.n140 163.367
R889 B.n145 B.n144 163.367
R890 B.n149 B.n148 163.367
R891 B.n153 B.n152 163.367
R892 B.n157 B.n156 163.367
R893 B.n161 B.n160 163.367
R894 B.n165 B.n164 163.367
R895 B.n169 B.n168 163.367
R896 B.n173 B.n172 163.367
R897 B.n177 B.n176 163.367
R898 B.n179 B.n102 163.367
R899 B.n293 B.t18 125.609
R900 B.n104 B.t12 125.609
R901 B.n291 B.t15 125.609
R902 B.n107 B.t9 125.609
R903 B.n373 B.n267 94.3854
R904 B.n373 B.n263 94.3854
R905 B.n379 B.n263 94.3854
R906 B.n379 B.n259 94.3854
R907 B.n385 B.n259 94.3854
R908 B.n385 B.n255 94.3854
R909 B.n391 B.n255 94.3854
R910 B.n397 B.n251 94.3854
R911 B.n397 B.n247 94.3854
R912 B.n403 B.n247 94.3854
R913 B.n403 B.n243 94.3854
R914 B.n409 B.n243 94.3854
R915 B.n409 B.n239 94.3854
R916 B.n415 B.n239 94.3854
R917 B.n415 B.n235 94.3854
R918 B.n421 B.n235 94.3854
R919 B.n421 B.n230 94.3854
R920 B.n427 B.n230 94.3854
R921 B.n427 B.n231 94.3854
R922 B.n433 B.n223 94.3854
R923 B.n439 B.n223 94.3854
R924 B.n439 B.n219 94.3854
R925 B.n445 B.n219 94.3854
R926 B.n445 B.n215 94.3854
R927 B.n451 B.n215 94.3854
R928 B.n451 B.n211 94.3854
R929 B.n457 B.n211 94.3854
R930 B.n463 B.n207 94.3854
R931 B.n463 B.n203 94.3854
R932 B.n469 B.n203 94.3854
R933 B.n469 B.n199 94.3854
R934 B.n475 B.n199 94.3854
R935 B.n475 B.n195 94.3854
R936 B.n482 B.n195 94.3854
R937 B.n482 B.n481 94.3854
R938 B.n488 B.n188 94.3854
R939 B.n495 B.n188 94.3854
R940 B.n495 B.n184 94.3854
R941 B.n501 B.n184 94.3854
R942 B.n501 B.n4 94.3854
R943 B.n655 B.n4 94.3854
R944 B.n655 B.n654 94.3854
R945 B.n654 B.n653 94.3854
R946 B.n653 B.n8 94.3854
R947 B.n647 B.n8 94.3854
R948 B.n647 B.n646 94.3854
R949 B.n646 B.n645 94.3854
R950 B.n639 B.n18 94.3854
R951 B.n639 B.n638 94.3854
R952 B.n638 B.n637 94.3854
R953 B.n637 B.n22 94.3854
R954 B.n631 B.n22 94.3854
R955 B.n631 B.n630 94.3854
R956 B.n630 B.n629 94.3854
R957 B.n629 B.n29 94.3854
R958 B.n623 B.n622 94.3854
R959 B.n622 B.n621 94.3854
R960 B.n621 B.n36 94.3854
R961 B.n615 B.n36 94.3854
R962 B.n615 B.n614 94.3854
R963 B.n614 B.n613 94.3854
R964 B.n613 B.n43 94.3854
R965 B.n607 B.n43 94.3854
R966 B.n606 B.n605 94.3854
R967 B.n605 B.n50 94.3854
R968 B.n599 B.n50 94.3854
R969 B.n599 B.n598 94.3854
R970 B.n598 B.n597 94.3854
R971 B.n597 B.n57 94.3854
R972 B.n591 B.n57 94.3854
R973 B.n591 B.n590 94.3854
R974 B.n590 B.n589 94.3854
R975 B.n589 B.n64 94.3854
R976 B.n583 B.n64 94.3854
R977 B.n583 B.n582 94.3854
R978 B.n581 B.n71 94.3854
R979 B.n575 B.n71 94.3854
R980 B.n575 B.n574 94.3854
R981 B.n574 B.n573 94.3854
R982 B.n573 B.n78 94.3854
R983 B.n567 B.n78 94.3854
R984 B.n567 B.n566 94.3854
R985 B.n391 B.t14 81.8932
R986 B.t7 B.n581 81.8932
R987 B.n481 B.t0 73.5652
R988 B.n18 B.t4 73.5652
R989 B.n366 B.n365 71.676
R990 B.n360 B.n271 71.676
R991 B.n357 B.n272 71.676
R992 B.n353 B.n273 71.676
R993 B.n349 B.n274 71.676
R994 B.n345 B.n275 71.676
R995 B.n341 B.n276 71.676
R996 B.n336 B.n277 71.676
R997 B.n332 B.n278 71.676
R998 B.n328 B.n279 71.676
R999 B.n324 B.n280 71.676
R1000 B.n320 B.n281 71.676
R1001 B.n315 B.n282 71.676
R1002 B.n311 B.n283 71.676
R1003 B.n307 B.n284 71.676
R1004 B.n303 B.n285 71.676
R1005 B.n299 B.n286 71.676
R1006 B.n295 B.n287 71.676
R1007 B.n109 B.n84 71.676
R1008 B.n113 B.n85 71.676
R1009 B.n117 B.n86 71.676
R1010 B.n121 B.n87 71.676
R1011 B.n125 B.n88 71.676
R1012 B.n129 B.n89 71.676
R1013 B.n133 B.n90 71.676
R1014 B.n137 B.n91 71.676
R1015 B.n141 B.n92 71.676
R1016 B.n145 B.n93 71.676
R1017 B.n149 B.n94 71.676
R1018 B.n153 B.n95 71.676
R1019 B.n157 B.n96 71.676
R1020 B.n161 B.n97 71.676
R1021 B.n165 B.n98 71.676
R1022 B.n169 B.n99 71.676
R1023 B.n173 B.n100 71.676
R1024 B.n177 B.n101 71.676
R1025 B.n564 B.n102 71.676
R1026 B.n564 B.n563 71.676
R1027 B.n179 B.n101 71.676
R1028 B.n176 B.n100 71.676
R1029 B.n172 B.n99 71.676
R1030 B.n168 B.n98 71.676
R1031 B.n164 B.n97 71.676
R1032 B.n160 B.n96 71.676
R1033 B.n156 B.n95 71.676
R1034 B.n152 B.n94 71.676
R1035 B.n148 B.n93 71.676
R1036 B.n144 B.n92 71.676
R1037 B.n140 B.n91 71.676
R1038 B.n136 B.n90 71.676
R1039 B.n132 B.n89 71.676
R1040 B.n128 B.n88 71.676
R1041 B.n124 B.n87 71.676
R1042 B.n120 B.n86 71.676
R1043 B.n116 B.n85 71.676
R1044 B.n112 B.n84 71.676
R1045 B.n366 B.n289 71.676
R1046 B.n358 B.n271 71.676
R1047 B.n354 B.n272 71.676
R1048 B.n350 B.n273 71.676
R1049 B.n346 B.n274 71.676
R1050 B.n342 B.n275 71.676
R1051 B.n337 B.n276 71.676
R1052 B.n333 B.n277 71.676
R1053 B.n329 B.n278 71.676
R1054 B.n325 B.n279 71.676
R1055 B.n321 B.n280 71.676
R1056 B.n316 B.n281 71.676
R1057 B.n312 B.n282 71.676
R1058 B.n308 B.n283 71.676
R1059 B.n304 B.n284 71.676
R1060 B.n300 B.n285 71.676
R1061 B.n296 B.n286 71.676
R1062 B.n287 B.n270 71.676
R1063 B.n433 B.t1 65.2371
R1064 B.n607 B.t5 65.2371
R1065 B.n293 B.n292 60.8975
R1066 B.n291 B.n290 60.8975
R1067 B.n107 B.n106 60.8975
R1068 B.n104 B.n103 60.8975
R1069 B.n318 B.n293 59.5399
R1070 B.n339 B.n291 59.5399
R1071 B.n108 B.n107 59.5399
R1072 B.n105 B.n104 59.5399
R1073 B.n457 B.t2 51.357
R1074 B.n623 B.t3 51.357
R1075 B.t2 B.n207 43.0289
R1076 B.t3 B.n29 43.0289
R1077 B.n110 B.n80 32.0005
R1078 B.n562 B.n561 32.0005
R1079 B.n370 B.n369 32.0005
R1080 B.n364 B.n265 32.0005
R1081 B.n231 B.t1 29.1488
R1082 B.t5 B.n606 29.1488
R1083 B.n488 B.t0 20.8207
R1084 B.n645 B.t4 20.8207
R1085 B B.n657 18.0485
R1086 B.t14 B.n251 12.4926
R1087 B.n582 B.t7 12.4926
R1088 B.n111 B.n110 10.6151
R1089 B.n114 B.n111 10.6151
R1090 B.n115 B.n114 10.6151
R1091 B.n118 B.n115 10.6151
R1092 B.n119 B.n118 10.6151
R1093 B.n122 B.n119 10.6151
R1094 B.n123 B.n122 10.6151
R1095 B.n126 B.n123 10.6151
R1096 B.n127 B.n126 10.6151
R1097 B.n130 B.n127 10.6151
R1098 B.n131 B.n130 10.6151
R1099 B.n134 B.n131 10.6151
R1100 B.n135 B.n134 10.6151
R1101 B.n139 B.n138 10.6151
R1102 B.n142 B.n139 10.6151
R1103 B.n143 B.n142 10.6151
R1104 B.n146 B.n143 10.6151
R1105 B.n147 B.n146 10.6151
R1106 B.n150 B.n147 10.6151
R1107 B.n151 B.n150 10.6151
R1108 B.n154 B.n151 10.6151
R1109 B.n155 B.n154 10.6151
R1110 B.n159 B.n158 10.6151
R1111 B.n162 B.n159 10.6151
R1112 B.n163 B.n162 10.6151
R1113 B.n166 B.n163 10.6151
R1114 B.n167 B.n166 10.6151
R1115 B.n170 B.n167 10.6151
R1116 B.n171 B.n170 10.6151
R1117 B.n174 B.n171 10.6151
R1118 B.n175 B.n174 10.6151
R1119 B.n178 B.n175 10.6151
R1120 B.n180 B.n178 10.6151
R1121 B.n181 B.n180 10.6151
R1122 B.n562 B.n181 10.6151
R1123 B.n371 B.n370 10.6151
R1124 B.n371 B.n261 10.6151
R1125 B.n381 B.n261 10.6151
R1126 B.n382 B.n381 10.6151
R1127 B.n383 B.n382 10.6151
R1128 B.n383 B.n253 10.6151
R1129 B.n393 B.n253 10.6151
R1130 B.n394 B.n393 10.6151
R1131 B.n395 B.n394 10.6151
R1132 B.n395 B.n245 10.6151
R1133 B.n405 B.n245 10.6151
R1134 B.n406 B.n405 10.6151
R1135 B.n407 B.n406 10.6151
R1136 B.n407 B.n237 10.6151
R1137 B.n417 B.n237 10.6151
R1138 B.n418 B.n417 10.6151
R1139 B.n419 B.n418 10.6151
R1140 B.n419 B.n228 10.6151
R1141 B.n429 B.n228 10.6151
R1142 B.n430 B.n429 10.6151
R1143 B.n431 B.n430 10.6151
R1144 B.n431 B.n221 10.6151
R1145 B.n441 B.n221 10.6151
R1146 B.n442 B.n441 10.6151
R1147 B.n443 B.n442 10.6151
R1148 B.n443 B.n213 10.6151
R1149 B.n453 B.n213 10.6151
R1150 B.n454 B.n453 10.6151
R1151 B.n455 B.n454 10.6151
R1152 B.n455 B.n205 10.6151
R1153 B.n465 B.n205 10.6151
R1154 B.n466 B.n465 10.6151
R1155 B.n467 B.n466 10.6151
R1156 B.n467 B.n197 10.6151
R1157 B.n477 B.n197 10.6151
R1158 B.n478 B.n477 10.6151
R1159 B.n479 B.n478 10.6151
R1160 B.n479 B.n190 10.6151
R1161 B.n490 B.n190 10.6151
R1162 B.n491 B.n490 10.6151
R1163 B.n493 B.n491 10.6151
R1164 B.n493 B.n492 10.6151
R1165 B.n492 B.n182 10.6151
R1166 B.n504 B.n182 10.6151
R1167 B.n505 B.n504 10.6151
R1168 B.n506 B.n505 10.6151
R1169 B.n507 B.n506 10.6151
R1170 B.n509 B.n507 10.6151
R1171 B.n510 B.n509 10.6151
R1172 B.n511 B.n510 10.6151
R1173 B.n512 B.n511 10.6151
R1174 B.n514 B.n512 10.6151
R1175 B.n515 B.n514 10.6151
R1176 B.n516 B.n515 10.6151
R1177 B.n517 B.n516 10.6151
R1178 B.n519 B.n517 10.6151
R1179 B.n520 B.n519 10.6151
R1180 B.n521 B.n520 10.6151
R1181 B.n522 B.n521 10.6151
R1182 B.n524 B.n522 10.6151
R1183 B.n525 B.n524 10.6151
R1184 B.n526 B.n525 10.6151
R1185 B.n527 B.n526 10.6151
R1186 B.n529 B.n527 10.6151
R1187 B.n530 B.n529 10.6151
R1188 B.n531 B.n530 10.6151
R1189 B.n532 B.n531 10.6151
R1190 B.n534 B.n532 10.6151
R1191 B.n535 B.n534 10.6151
R1192 B.n536 B.n535 10.6151
R1193 B.n537 B.n536 10.6151
R1194 B.n539 B.n537 10.6151
R1195 B.n540 B.n539 10.6151
R1196 B.n541 B.n540 10.6151
R1197 B.n542 B.n541 10.6151
R1198 B.n544 B.n542 10.6151
R1199 B.n545 B.n544 10.6151
R1200 B.n546 B.n545 10.6151
R1201 B.n547 B.n546 10.6151
R1202 B.n549 B.n547 10.6151
R1203 B.n550 B.n549 10.6151
R1204 B.n551 B.n550 10.6151
R1205 B.n552 B.n551 10.6151
R1206 B.n554 B.n552 10.6151
R1207 B.n555 B.n554 10.6151
R1208 B.n556 B.n555 10.6151
R1209 B.n557 B.n556 10.6151
R1210 B.n559 B.n557 10.6151
R1211 B.n560 B.n559 10.6151
R1212 B.n561 B.n560 10.6151
R1213 B.n364 B.n363 10.6151
R1214 B.n363 B.n362 10.6151
R1215 B.n362 B.n361 10.6151
R1216 B.n361 B.n359 10.6151
R1217 B.n359 B.n356 10.6151
R1218 B.n356 B.n355 10.6151
R1219 B.n355 B.n352 10.6151
R1220 B.n352 B.n351 10.6151
R1221 B.n351 B.n348 10.6151
R1222 B.n348 B.n347 10.6151
R1223 B.n347 B.n344 10.6151
R1224 B.n344 B.n343 10.6151
R1225 B.n343 B.n340 10.6151
R1226 B.n338 B.n335 10.6151
R1227 B.n335 B.n334 10.6151
R1228 B.n334 B.n331 10.6151
R1229 B.n331 B.n330 10.6151
R1230 B.n330 B.n327 10.6151
R1231 B.n327 B.n326 10.6151
R1232 B.n326 B.n323 10.6151
R1233 B.n323 B.n322 10.6151
R1234 B.n322 B.n319 10.6151
R1235 B.n317 B.n314 10.6151
R1236 B.n314 B.n313 10.6151
R1237 B.n313 B.n310 10.6151
R1238 B.n310 B.n309 10.6151
R1239 B.n309 B.n306 10.6151
R1240 B.n306 B.n305 10.6151
R1241 B.n305 B.n302 10.6151
R1242 B.n302 B.n301 10.6151
R1243 B.n301 B.n298 10.6151
R1244 B.n298 B.n297 10.6151
R1245 B.n297 B.n294 10.6151
R1246 B.n294 B.n269 10.6151
R1247 B.n369 B.n269 10.6151
R1248 B.n375 B.n265 10.6151
R1249 B.n376 B.n375 10.6151
R1250 B.n377 B.n376 10.6151
R1251 B.n377 B.n257 10.6151
R1252 B.n387 B.n257 10.6151
R1253 B.n388 B.n387 10.6151
R1254 B.n389 B.n388 10.6151
R1255 B.n389 B.n249 10.6151
R1256 B.n399 B.n249 10.6151
R1257 B.n400 B.n399 10.6151
R1258 B.n401 B.n400 10.6151
R1259 B.n401 B.n241 10.6151
R1260 B.n411 B.n241 10.6151
R1261 B.n412 B.n411 10.6151
R1262 B.n413 B.n412 10.6151
R1263 B.n413 B.n233 10.6151
R1264 B.n423 B.n233 10.6151
R1265 B.n424 B.n423 10.6151
R1266 B.n425 B.n424 10.6151
R1267 B.n425 B.n225 10.6151
R1268 B.n435 B.n225 10.6151
R1269 B.n436 B.n435 10.6151
R1270 B.n437 B.n436 10.6151
R1271 B.n437 B.n217 10.6151
R1272 B.n447 B.n217 10.6151
R1273 B.n448 B.n447 10.6151
R1274 B.n449 B.n448 10.6151
R1275 B.n449 B.n209 10.6151
R1276 B.n459 B.n209 10.6151
R1277 B.n460 B.n459 10.6151
R1278 B.n461 B.n460 10.6151
R1279 B.n461 B.n201 10.6151
R1280 B.n471 B.n201 10.6151
R1281 B.n472 B.n471 10.6151
R1282 B.n473 B.n472 10.6151
R1283 B.n473 B.n193 10.6151
R1284 B.n484 B.n193 10.6151
R1285 B.n485 B.n484 10.6151
R1286 B.n486 B.n485 10.6151
R1287 B.n486 B.n186 10.6151
R1288 B.n497 B.n186 10.6151
R1289 B.n498 B.n497 10.6151
R1290 B.n499 B.n498 10.6151
R1291 B.n499 B.n0 10.6151
R1292 B.n651 B.n1 10.6151
R1293 B.n651 B.n650 10.6151
R1294 B.n650 B.n649 10.6151
R1295 B.n649 B.n10 10.6151
R1296 B.n643 B.n10 10.6151
R1297 B.n643 B.n642 10.6151
R1298 B.n642 B.n641 10.6151
R1299 B.n641 B.n16 10.6151
R1300 B.n635 B.n16 10.6151
R1301 B.n635 B.n634 10.6151
R1302 B.n634 B.n633 10.6151
R1303 B.n633 B.n24 10.6151
R1304 B.n627 B.n24 10.6151
R1305 B.n627 B.n626 10.6151
R1306 B.n626 B.n625 10.6151
R1307 B.n625 B.n31 10.6151
R1308 B.n619 B.n31 10.6151
R1309 B.n619 B.n618 10.6151
R1310 B.n618 B.n617 10.6151
R1311 B.n617 B.n38 10.6151
R1312 B.n611 B.n38 10.6151
R1313 B.n611 B.n610 10.6151
R1314 B.n610 B.n609 10.6151
R1315 B.n609 B.n45 10.6151
R1316 B.n603 B.n45 10.6151
R1317 B.n603 B.n602 10.6151
R1318 B.n602 B.n601 10.6151
R1319 B.n601 B.n52 10.6151
R1320 B.n595 B.n52 10.6151
R1321 B.n595 B.n594 10.6151
R1322 B.n594 B.n593 10.6151
R1323 B.n593 B.n59 10.6151
R1324 B.n587 B.n59 10.6151
R1325 B.n587 B.n586 10.6151
R1326 B.n586 B.n585 10.6151
R1327 B.n585 B.n66 10.6151
R1328 B.n579 B.n66 10.6151
R1329 B.n579 B.n578 10.6151
R1330 B.n578 B.n577 10.6151
R1331 B.n577 B.n73 10.6151
R1332 B.n571 B.n73 10.6151
R1333 B.n571 B.n570 10.6151
R1334 B.n570 B.n569 10.6151
R1335 B.n569 B.n80 10.6151
R1336 B.n135 B.n108 9.36635
R1337 B.n158 B.n105 9.36635
R1338 B.n340 B.n339 9.36635
R1339 B.n318 B.n317 9.36635
R1340 B.n657 B.n0 2.81026
R1341 B.n657 B.n1 2.81026
R1342 B.n138 B.n108 1.24928
R1343 B.n155 B.n105 1.24928
R1344 B.n339 B.n338 1.24928
R1345 B.n319 B.n318 1.24928
R1346 VP.n13 VP.n12 161.3
R1347 VP.n14 VP.n9 161.3
R1348 VP.n16 VP.n15 161.3
R1349 VP.n17 VP.n8 161.3
R1350 VP.n19 VP.n18 161.3
R1351 VP.n20 VP.n7 161.3
R1352 VP.n43 VP.n0 161.3
R1353 VP.n42 VP.n41 161.3
R1354 VP.n40 VP.n1 161.3
R1355 VP.n39 VP.n38 161.3
R1356 VP.n37 VP.n2 161.3
R1357 VP.n36 VP.n35 161.3
R1358 VP.n34 VP.n3 161.3
R1359 VP.n33 VP.n32 161.3
R1360 VP.n31 VP.n4 161.3
R1361 VP.n30 VP.n29 161.3
R1362 VP.n28 VP.n5 161.3
R1363 VP.n27 VP.n26 161.3
R1364 VP.n25 VP.n6 161.3
R1365 VP.n24 VP.n23 103.906
R1366 VP.n45 VP.n44 103.906
R1367 VP.n22 VP.n21 103.906
R1368 VP.n11 VP.t1 57.3801
R1369 VP.n11 VP.n10 48.9126
R1370 VP.n30 VP.n5 47.2923
R1371 VP.n38 VP.n1 47.2923
R1372 VP.n15 VP.n8 47.2923
R1373 VP.n23 VP.n22 42.439
R1374 VP.n31 VP.n30 33.6945
R1375 VP.n38 VP.n37 33.6945
R1376 VP.n15 VP.n14 33.6945
R1377 VP.n26 VP.n25 24.4675
R1378 VP.n26 VP.n5 24.4675
R1379 VP.n32 VP.n31 24.4675
R1380 VP.n32 VP.n3 24.4675
R1381 VP.n36 VP.n3 24.4675
R1382 VP.n37 VP.n36 24.4675
R1383 VP.n42 VP.n1 24.4675
R1384 VP.n43 VP.n42 24.4675
R1385 VP.n19 VP.n8 24.4675
R1386 VP.n20 VP.n19 24.4675
R1387 VP.n13 VP.n10 24.4675
R1388 VP.n14 VP.n13 24.4675
R1389 VP.n3 VP.t5 22.7283
R1390 VP.n24 VP.t4 22.7283
R1391 VP.n44 VP.t3 22.7283
R1392 VP.n10 VP.t0 22.7283
R1393 VP.n21 VP.t2 22.7283
R1394 VP.n25 VP.n24 6.85126
R1395 VP.n44 VP.n43 6.85126
R1396 VP.n21 VP.n20 6.85126
R1397 VP.n12 VP.n11 4.90017
R1398 VP.n22 VP.n7 0.278367
R1399 VP.n23 VP.n6 0.278367
R1400 VP.n45 VP.n0 0.278367
R1401 VP.n12 VP.n9 0.189894
R1402 VP.n16 VP.n9 0.189894
R1403 VP.n17 VP.n16 0.189894
R1404 VP.n18 VP.n17 0.189894
R1405 VP.n18 VP.n7 0.189894
R1406 VP.n27 VP.n6 0.189894
R1407 VP.n28 VP.n27 0.189894
R1408 VP.n29 VP.n28 0.189894
R1409 VP.n29 VP.n4 0.189894
R1410 VP.n33 VP.n4 0.189894
R1411 VP.n34 VP.n33 0.189894
R1412 VP.n35 VP.n34 0.189894
R1413 VP.n35 VP.n2 0.189894
R1414 VP.n39 VP.n2 0.189894
R1415 VP.n40 VP.n39 0.189894
R1416 VP.n41 VP.n40 0.189894
R1417 VP.n41 VP.n0 0.189894
R1418 VP VP.n45 0.153454
R1419 VDD1.n6 VDD1.n0 289.615
R1420 VDD1.n17 VDD1.n11 289.615
R1421 VDD1.n7 VDD1.n6 185
R1422 VDD1.n5 VDD1.n4 185
R1423 VDD1.n16 VDD1.n15 185
R1424 VDD1.n18 VDD1.n17 185
R1425 VDD1.n14 VDD1.t1 153.582
R1426 VDD1.n3 VDD1.t4 153.582
R1427 VDD1.n6 VDD1.n5 104.615
R1428 VDD1.n17 VDD1.n16 104.615
R1429 VDD1.n23 VDD1.n22 84.9062
R1430 VDD1.n25 VDD1.n24 84.2848
R1431 VDD1.n5 VDD1.t4 52.3082
R1432 VDD1.n16 VDD1.t1 52.3082
R1433 VDD1 VDD1.n10 48.8192
R1434 VDD1.n23 VDD1.n21 48.7056
R1435 VDD1.n25 VDD1.n23 36.7337
R1436 VDD1.n4 VDD1.n3 10.1164
R1437 VDD1.n15 VDD1.n14 10.1164
R1438 VDD1.n10 VDD1.n9 9.45567
R1439 VDD1.n21 VDD1.n20 9.45567
R1440 VDD1.n9 VDD1.n8 9.3005
R1441 VDD1.n2 VDD1.n1 9.3005
R1442 VDD1.n13 VDD1.n12 9.3005
R1443 VDD1.n20 VDD1.n19 9.3005
R1444 VDD1.n10 VDD1.n0 8.92171
R1445 VDD1.n21 VDD1.n11 8.92171
R1446 VDD1.n8 VDD1.n7 8.14595
R1447 VDD1.n19 VDD1.n18 8.14595
R1448 VDD1.n24 VDD1.t5 7.4722
R1449 VDD1.n24 VDD1.t3 7.4722
R1450 VDD1.n22 VDD1.t0 7.4722
R1451 VDD1.n22 VDD1.t2 7.4722
R1452 VDD1.n4 VDD1.n2 7.3702
R1453 VDD1.n15 VDD1.n13 7.3702
R1454 VDD1.n7 VDD1.n2 5.81868
R1455 VDD1.n18 VDD1.n13 5.81868
R1456 VDD1.n8 VDD1.n0 5.04292
R1457 VDD1.n19 VDD1.n11 5.04292
R1458 VDD1.n3 VDD1.n1 3.00987
R1459 VDD1.n14 VDD1.n12 3.00987
R1460 VDD1 VDD1.n25 0.619035
R1461 VDD1.n9 VDD1.n1 0.155672
R1462 VDD1.n20 VDD1.n12 0.155672
C0 VDD1 VDD2 1.4872f
C1 VTAIL VDD1 4.4789f
C2 VTAIL VDD2 4.53337f
C3 VDD1 VN 0.156462f
C4 VDD2 VN 1.81385f
C5 VDD1 VP 2.13648f
C6 VTAIL VN 2.67356f
C7 VDD2 VP 0.481678f
C8 VTAIL VP 2.6877f
C9 VN VP 5.40364f
C10 VDD2 B 4.305495f
C11 VDD1 B 4.62102f
C12 VTAIL B 3.805978f
C13 VN B 12.465289f
C14 VP B 11.27641f
C15 VDD1.n0 B 0.033215f
C16 VDD1.n1 B 0.19801f
C17 VDD1.n2 B 0.0124f
C18 VDD1.t4 B 0.053065f
C19 VDD1.n3 B 0.085938f
C20 VDD1.n4 B 0.020068f
C21 VDD1.n5 B 0.021983f
C22 VDD1.n6 B 0.064828f
C23 VDD1.n7 B 0.01313f
C24 VDD1.n8 B 0.0124f
C25 VDD1.n9 B 0.049873f
C26 VDD1.n10 B 0.060728f
C27 VDD1.n11 B 0.033215f
C28 VDD1.n12 B 0.19801f
C29 VDD1.n13 B 0.0124f
C30 VDD1.t1 B 0.053065f
C31 VDD1.n14 B 0.085938f
C32 VDD1.n15 B 0.020068f
C33 VDD1.n16 B 0.021983f
C34 VDD1.n17 B 0.064828f
C35 VDD1.n18 B 0.01313f
C36 VDD1.n19 B 0.0124f
C37 VDD1.n20 B 0.049873f
C38 VDD1.n21 B 0.059956f
C39 VDD1.t0 B 0.048325f
C40 VDD1.t2 B 0.048325f
C41 VDD1.n22 B 0.339881f
C42 VDD1.n23 B 2.13949f
C43 VDD1.t5 B 0.048325f
C44 VDD1.t3 B 0.048325f
C45 VDD1.n24 B 0.336666f
C46 VDD1.n25 B 1.9496f
C47 VP.n0 B 0.040434f
C48 VP.t3 B 0.559517f
C49 VP.n1 B 0.057974f
C50 VP.n2 B 0.030669f
C51 VP.t5 B 0.559517f
C52 VP.n3 B 0.270501f
C53 VP.n4 B 0.030669f
C54 VP.n5 B 0.057974f
C55 VP.n6 B 0.040434f
C56 VP.t4 B 0.559517f
C57 VP.n7 B 0.040434f
C58 VP.t2 B 0.559517f
C59 VP.n8 B 0.057974f
C60 VP.n9 B 0.030669f
C61 VP.t0 B 0.559517f
C62 VP.n10 B 0.351418f
C63 VP.t1 B 0.8306f
C64 VP.n11 B 0.322855f
C65 VP.n12 B 0.322134f
C66 VP.n13 B 0.05716f
C67 VP.n14 B 0.061949f
C68 VP.n15 B 0.026779f
C69 VP.n16 B 0.030669f
C70 VP.n17 B 0.030669f
C71 VP.n18 B 0.030669f
C72 VP.n19 B 0.05716f
C73 VP.n20 B 0.036841f
C74 VP.n21 B 0.347696f
C75 VP.n22 B 1.3323f
C76 VP.n23 B 1.35828f
C77 VP.n24 B 0.347696f
C78 VP.n25 B 0.036841f
C79 VP.n26 B 0.05716f
C80 VP.n27 B 0.030669f
C81 VP.n28 B 0.030669f
C82 VP.n29 B 0.030669f
C83 VP.n30 B 0.026779f
C84 VP.n31 B 0.061949f
C85 VP.n32 B 0.05716f
C86 VP.n33 B 0.030669f
C87 VP.n34 B 0.030669f
C88 VP.n35 B 0.030669f
C89 VP.n36 B 0.05716f
C90 VP.n37 B 0.061949f
C91 VP.n38 B 0.026779f
C92 VP.n39 B 0.030669f
C93 VP.n40 B 0.030669f
C94 VP.n41 B 0.030669f
C95 VP.n42 B 0.05716f
C96 VP.n43 B 0.036841f
C97 VP.n44 B 0.347696f
C98 VP.n45 B 0.054501f
C99 VTAIL.t8 B 0.068867f
C100 VTAIL.t11 B 0.068867f
C101 VTAIL.n0 B 0.417372f
C102 VTAIL.n1 B 0.547966f
C103 VTAIL.n2 B 0.047334f
C104 VTAIL.n3 B 0.282178f
C105 VTAIL.n4 B 0.017671f
C106 VTAIL.t0 B 0.075621f
C107 VTAIL.n5 B 0.122468f
C108 VTAIL.n6 B 0.028599f
C109 VTAIL.n7 B 0.031327f
C110 VTAIL.n8 B 0.092384f
C111 VTAIL.n9 B 0.018711f
C112 VTAIL.n10 B 0.017671f
C113 VTAIL.n11 B 0.071072f
C114 VTAIL.n12 B 0.051738f
C115 VTAIL.n13 B 0.505346f
C116 VTAIL.t1 B 0.068867f
C117 VTAIL.t2 B 0.068867f
C118 VTAIL.n14 B 0.417372f
C119 VTAIL.n15 B 1.82619f
C120 VTAIL.t7 B 0.068867f
C121 VTAIL.t9 B 0.068867f
C122 VTAIL.n16 B 0.417375f
C123 VTAIL.n17 B 1.82619f
C124 VTAIL.n18 B 0.047334f
C125 VTAIL.n19 B 0.282178f
C126 VTAIL.n20 B 0.017671f
C127 VTAIL.t10 B 0.075621f
C128 VTAIL.n21 B 0.122468f
C129 VTAIL.n22 B 0.028599f
C130 VTAIL.n23 B 0.031327f
C131 VTAIL.n24 B 0.092384f
C132 VTAIL.n25 B 0.018711f
C133 VTAIL.n26 B 0.017671f
C134 VTAIL.n27 B 0.071072f
C135 VTAIL.n28 B 0.051738f
C136 VTAIL.n29 B 0.505346f
C137 VTAIL.t4 B 0.068867f
C138 VTAIL.t3 B 0.068867f
C139 VTAIL.n30 B 0.417375f
C140 VTAIL.n31 B 0.756927f
C141 VTAIL.n32 B 0.047334f
C142 VTAIL.n33 B 0.282178f
C143 VTAIL.n34 B 0.017671f
C144 VTAIL.t5 B 0.075621f
C145 VTAIL.n35 B 0.122468f
C146 VTAIL.n36 B 0.028599f
C147 VTAIL.n37 B 0.031327f
C148 VTAIL.n38 B 0.092384f
C149 VTAIL.n39 B 0.018711f
C150 VTAIL.n40 B 0.017671f
C151 VTAIL.n41 B 0.071072f
C152 VTAIL.n42 B 0.051738f
C153 VTAIL.n43 B 1.28777f
C154 VTAIL.n44 B 0.047334f
C155 VTAIL.n45 B 0.282178f
C156 VTAIL.n46 B 0.017671f
C157 VTAIL.t6 B 0.075621f
C158 VTAIL.n47 B 0.122468f
C159 VTAIL.n48 B 0.028599f
C160 VTAIL.n49 B 0.031327f
C161 VTAIL.n50 B 0.092384f
C162 VTAIL.n51 B 0.018711f
C163 VTAIL.n52 B 0.017671f
C164 VTAIL.n53 B 0.071072f
C165 VTAIL.n54 B 0.051738f
C166 VTAIL.n55 B 1.2099f
C167 VDD2.n0 B 0.022943f
C168 VDD2.n1 B 0.136773f
C169 VDD2.n2 B 0.008565f
C170 VDD2.t4 B 0.036654f
C171 VDD2.n3 B 0.059361f
C172 VDD2.n4 B 0.013862f
C173 VDD2.n5 B 0.015184f
C174 VDD2.n6 B 0.044779f
C175 VDD2.n7 B 0.009069f
C176 VDD2.n8 B 0.008565f
C177 VDD2.n9 B 0.034449f
C178 VDD2.n10 B 0.041414f
C179 VDD2.t1 B 0.03338f
C180 VDD2.t3 B 0.03338f
C181 VDD2.n11 B 0.234769f
C182 VDD2.n12 B 1.40164f
C183 VDD2.n13 B 0.022943f
C184 VDD2.n14 B 0.136773f
C185 VDD2.n15 B 0.008565f
C186 VDD2.t0 B 0.036654f
C187 VDD2.n16 B 0.059361f
C188 VDD2.n17 B 0.013862f
C189 VDD2.n18 B 0.015184f
C190 VDD2.n19 B 0.044779f
C191 VDD2.n20 B 0.009069f
C192 VDD2.n21 B 0.008565f
C193 VDD2.n22 B 0.034449f
C194 VDD2.n23 B 0.036104f
C195 VDD2.n24 B 1.19772f
C196 VDD2.t5 B 0.03338f
C197 VDD2.t2 B 0.03338f
C198 VDD2.n25 B 0.234754f
C199 VN.n0 B 0.031974f
C200 VN.t5 B 0.442452f
C201 VN.n1 B 0.045845f
C202 VN.n2 B 0.024252f
C203 VN.t0 B 0.442452f
C204 VN.n3 B 0.277893f
C205 VN.t3 B 0.656818f
C206 VN.n4 B 0.255305f
C207 VN.n5 B 0.254736f
C208 VN.n6 B 0.045201f
C209 VN.n7 B 0.048988f
C210 VN.n8 B 0.021176f
C211 VN.n9 B 0.024252f
C212 VN.n10 B 0.024252f
C213 VN.n11 B 0.024252f
C214 VN.n12 B 0.045201f
C215 VN.n13 B 0.029133f
C216 VN.n14 B 0.27495f
C217 VN.n15 B 0.043098f
C218 VN.n16 B 0.031974f
C219 VN.t4 B 0.442452f
C220 VN.n17 B 0.045845f
C221 VN.n18 B 0.024252f
C222 VN.t2 B 0.442452f
C223 VN.n19 B 0.277893f
C224 VN.t1 B 0.656818f
C225 VN.n20 B 0.255305f
C226 VN.n21 B 0.254736f
C227 VN.n22 B 0.045201f
C228 VN.n23 B 0.048988f
C229 VN.n24 B 0.021176f
C230 VN.n25 B 0.024252f
C231 VN.n26 B 0.024252f
C232 VN.n27 B 0.024252f
C233 VN.n28 B 0.045201f
C234 VN.n29 B 0.029133f
C235 VN.n30 B 0.27495f
C236 VN.n31 B 1.06695f
.ends

