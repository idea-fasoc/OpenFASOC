* NGSPICE file created from diff_pair_sample_1007.ext - technology: sky130A

.subckt diff_pair_sample_1007 VTAIL VN VP B VDD2 VDD1
X0 B.t11 B.t9 B.t10 w_n1378_n1594# sky130_fd_pr__pfet_01v8 ad=1.2207 pd=7.04 as=0 ps=0 w=3.13 l=0.18
X1 VDD1.t5 VP.t0 VTAIL.t7 w_n1378_n1594# sky130_fd_pr__pfet_01v8 ad=1.2207 pd=7.04 as=0.51645 ps=3.46 w=3.13 l=0.18
X2 B.t8 B.t6 B.t7 w_n1378_n1594# sky130_fd_pr__pfet_01v8 ad=1.2207 pd=7.04 as=0 ps=0 w=3.13 l=0.18
X3 VDD2.t5 VN.t0 VTAIL.t3 w_n1378_n1594# sky130_fd_pr__pfet_01v8 ad=0.51645 pd=3.46 as=1.2207 ps=7.04 w=3.13 l=0.18
X4 VDD2.t4 VN.t1 VTAIL.t4 w_n1378_n1594# sky130_fd_pr__pfet_01v8 ad=1.2207 pd=7.04 as=0.51645 ps=3.46 w=3.13 l=0.18
X5 VTAIL.t5 VN.t2 VDD2.t3 w_n1378_n1594# sky130_fd_pr__pfet_01v8 ad=0.51645 pd=3.46 as=0.51645 ps=3.46 w=3.13 l=0.18
X6 B.t5 B.t3 B.t4 w_n1378_n1594# sky130_fd_pr__pfet_01v8 ad=1.2207 pd=7.04 as=0 ps=0 w=3.13 l=0.18
X7 B.t2 B.t0 B.t1 w_n1378_n1594# sky130_fd_pr__pfet_01v8 ad=1.2207 pd=7.04 as=0 ps=0 w=3.13 l=0.18
X8 VDD2.t2 VN.t3 VTAIL.t2 w_n1378_n1594# sky130_fd_pr__pfet_01v8 ad=1.2207 pd=7.04 as=0.51645 ps=3.46 w=3.13 l=0.18
X9 VDD1.t4 VP.t1 VTAIL.t6 w_n1378_n1594# sky130_fd_pr__pfet_01v8 ad=1.2207 pd=7.04 as=0.51645 ps=3.46 w=3.13 l=0.18
X10 VTAIL.t8 VP.t2 VDD1.t3 w_n1378_n1594# sky130_fd_pr__pfet_01v8 ad=0.51645 pd=3.46 as=0.51645 ps=3.46 w=3.13 l=0.18
X11 VDD1.t2 VP.t3 VTAIL.t9 w_n1378_n1594# sky130_fd_pr__pfet_01v8 ad=0.51645 pd=3.46 as=1.2207 ps=7.04 w=3.13 l=0.18
X12 VDD1.t1 VP.t4 VTAIL.t10 w_n1378_n1594# sky130_fd_pr__pfet_01v8 ad=0.51645 pd=3.46 as=1.2207 ps=7.04 w=3.13 l=0.18
X13 VTAIL.t1 VN.t4 VDD2.t1 w_n1378_n1594# sky130_fd_pr__pfet_01v8 ad=0.51645 pd=3.46 as=0.51645 ps=3.46 w=3.13 l=0.18
X14 VDD2.t0 VN.t5 VTAIL.t0 w_n1378_n1594# sky130_fd_pr__pfet_01v8 ad=0.51645 pd=3.46 as=1.2207 ps=7.04 w=3.13 l=0.18
X15 VTAIL.t11 VP.t5 VDD1.t0 w_n1378_n1594# sky130_fd_pr__pfet_01v8 ad=0.51645 pd=3.46 as=0.51645 ps=3.46 w=3.13 l=0.18
R0 B.n56 B.t3 662.117
R1 B.n64 B.t9 662.117
R2 B.n18 B.t0 662.117
R3 B.n24 B.t6 662.117
R4 B.n206 B.n33 585
R5 B.n208 B.n207 585
R6 B.n209 B.n32 585
R7 B.n211 B.n210 585
R8 B.n212 B.n31 585
R9 B.n214 B.n213 585
R10 B.n215 B.n30 585
R11 B.n217 B.n216 585
R12 B.n218 B.n29 585
R13 B.n220 B.n219 585
R14 B.n221 B.n28 585
R15 B.n223 B.n222 585
R16 B.n224 B.n27 585
R17 B.n226 B.n225 585
R18 B.n227 B.n26 585
R19 B.n229 B.n228 585
R20 B.n231 B.n23 585
R21 B.n233 B.n232 585
R22 B.n234 B.n22 585
R23 B.n236 B.n235 585
R24 B.n237 B.n21 585
R25 B.n239 B.n238 585
R26 B.n240 B.n20 585
R27 B.n242 B.n241 585
R28 B.n243 B.n17 585
R29 B.n246 B.n245 585
R30 B.n247 B.n16 585
R31 B.n249 B.n248 585
R32 B.n250 B.n15 585
R33 B.n252 B.n251 585
R34 B.n253 B.n14 585
R35 B.n255 B.n254 585
R36 B.n256 B.n13 585
R37 B.n258 B.n257 585
R38 B.n259 B.n12 585
R39 B.n261 B.n260 585
R40 B.n262 B.n11 585
R41 B.n264 B.n263 585
R42 B.n265 B.n10 585
R43 B.n267 B.n266 585
R44 B.n268 B.n9 585
R45 B.n205 B.n204 585
R46 B.n203 B.n34 585
R47 B.n202 B.n201 585
R48 B.n200 B.n35 585
R49 B.n199 B.n198 585
R50 B.n197 B.n36 585
R51 B.n196 B.n195 585
R52 B.n194 B.n37 585
R53 B.n193 B.n192 585
R54 B.n191 B.n38 585
R55 B.n190 B.n189 585
R56 B.n188 B.n39 585
R57 B.n187 B.n186 585
R58 B.n185 B.n40 585
R59 B.n184 B.n183 585
R60 B.n182 B.n41 585
R61 B.n181 B.n180 585
R62 B.n179 B.n42 585
R63 B.n178 B.n177 585
R64 B.n176 B.n43 585
R65 B.n175 B.n174 585
R66 B.n173 B.n44 585
R67 B.n172 B.n171 585
R68 B.n170 B.n45 585
R69 B.n169 B.n168 585
R70 B.n167 B.n46 585
R71 B.n166 B.n165 585
R72 B.n164 B.n47 585
R73 B.n163 B.n162 585
R74 B.n100 B.n99 585
R75 B.n101 B.n72 585
R76 B.n103 B.n102 585
R77 B.n104 B.n71 585
R78 B.n106 B.n105 585
R79 B.n107 B.n70 585
R80 B.n109 B.n108 585
R81 B.n110 B.n69 585
R82 B.n112 B.n111 585
R83 B.n113 B.n68 585
R84 B.n115 B.n114 585
R85 B.n116 B.n67 585
R86 B.n118 B.n117 585
R87 B.n119 B.n66 585
R88 B.n121 B.n120 585
R89 B.n122 B.n63 585
R90 B.n125 B.n124 585
R91 B.n126 B.n62 585
R92 B.n128 B.n127 585
R93 B.n129 B.n61 585
R94 B.n131 B.n130 585
R95 B.n132 B.n60 585
R96 B.n134 B.n133 585
R97 B.n135 B.n59 585
R98 B.n137 B.n136 585
R99 B.n139 B.n138 585
R100 B.n140 B.n55 585
R101 B.n142 B.n141 585
R102 B.n143 B.n54 585
R103 B.n145 B.n144 585
R104 B.n146 B.n53 585
R105 B.n148 B.n147 585
R106 B.n149 B.n52 585
R107 B.n151 B.n150 585
R108 B.n152 B.n51 585
R109 B.n154 B.n153 585
R110 B.n155 B.n50 585
R111 B.n157 B.n156 585
R112 B.n158 B.n49 585
R113 B.n160 B.n159 585
R114 B.n161 B.n48 585
R115 B.n98 B.n73 585
R116 B.n97 B.n96 585
R117 B.n95 B.n74 585
R118 B.n94 B.n93 585
R119 B.n92 B.n75 585
R120 B.n91 B.n90 585
R121 B.n89 B.n76 585
R122 B.n88 B.n87 585
R123 B.n86 B.n77 585
R124 B.n85 B.n84 585
R125 B.n83 B.n78 585
R126 B.n82 B.n81 585
R127 B.n80 B.n79 585
R128 B.n2 B.n0 585
R129 B.n289 B.n1 585
R130 B.n288 B.n287 585
R131 B.n286 B.n3 585
R132 B.n285 B.n284 585
R133 B.n283 B.n4 585
R134 B.n282 B.n281 585
R135 B.n280 B.n5 585
R136 B.n279 B.n278 585
R137 B.n277 B.n6 585
R138 B.n276 B.n275 585
R139 B.n274 B.n7 585
R140 B.n273 B.n272 585
R141 B.n271 B.n8 585
R142 B.n270 B.n269 585
R143 B.n291 B.n290 585
R144 B.n100 B.n73 487.695
R145 B.n270 B.n9 487.695
R146 B.n162 B.n161 487.695
R147 B.n204 B.n33 487.695
R148 B.n56 B.t5 234.095
R149 B.n24 B.t7 234.095
R150 B.n64 B.t11 234.095
R151 B.n18 B.t1 234.095
R152 B.n57 B.t4 224.203
R153 B.n25 B.t8 224.203
R154 B.n65 B.t10 224.203
R155 B.n19 B.t2 224.203
R156 B.n96 B.n73 163.367
R157 B.n96 B.n95 163.367
R158 B.n95 B.n94 163.367
R159 B.n94 B.n75 163.367
R160 B.n90 B.n75 163.367
R161 B.n90 B.n89 163.367
R162 B.n89 B.n88 163.367
R163 B.n88 B.n77 163.367
R164 B.n84 B.n77 163.367
R165 B.n84 B.n83 163.367
R166 B.n83 B.n82 163.367
R167 B.n82 B.n79 163.367
R168 B.n79 B.n2 163.367
R169 B.n290 B.n2 163.367
R170 B.n290 B.n289 163.367
R171 B.n289 B.n288 163.367
R172 B.n288 B.n3 163.367
R173 B.n284 B.n3 163.367
R174 B.n284 B.n283 163.367
R175 B.n283 B.n282 163.367
R176 B.n282 B.n5 163.367
R177 B.n278 B.n5 163.367
R178 B.n278 B.n277 163.367
R179 B.n277 B.n276 163.367
R180 B.n276 B.n7 163.367
R181 B.n272 B.n7 163.367
R182 B.n272 B.n271 163.367
R183 B.n271 B.n270 163.367
R184 B.n101 B.n100 163.367
R185 B.n102 B.n101 163.367
R186 B.n102 B.n71 163.367
R187 B.n106 B.n71 163.367
R188 B.n107 B.n106 163.367
R189 B.n108 B.n107 163.367
R190 B.n108 B.n69 163.367
R191 B.n112 B.n69 163.367
R192 B.n113 B.n112 163.367
R193 B.n114 B.n113 163.367
R194 B.n114 B.n67 163.367
R195 B.n118 B.n67 163.367
R196 B.n119 B.n118 163.367
R197 B.n120 B.n119 163.367
R198 B.n120 B.n63 163.367
R199 B.n125 B.n63 163.367
R200 B.n126 B.n125 163.367
R201 B.n127 B.n126 163.367
R202 B.n127 B.n61 163.367
R203 B.n131 B.n61 163.367
R204 B.n132 B.n131 163.367
R205 B.n133 B.n132 163.367
R206 B.n133 B.n59 163.367
R207 B.n137 B.n59 163.367
R208 B.n138 B.n137 163.367
R209 B.n138 B.n55 163.367
R210 B.n142 B.n55 163.367
R211 B.n143 B.n142 163.367
R212 B.n144 B.n143 163.367
R213 B.n144 B.n53 163.367
R214 B.n148 B.n53 163.367
R215 B.n149 B.n148 163.367
R216 B.n150 B.n149 163.367
R217 B.n150 B.n51 163.367
R218 B.n154 B.n51 163.367
R219 B.n155 B.n154 163.367
R220 B.n156 B.n155 163.367
R221 B.n156 B.n49 163.367
R222 B.n160 B.n49 163.367
R223 B.n161 B.n160 163.367
R224 B.n162 B.n47 163.367
R225 B.n166 B.n47 163.367
R226 B.n167 B.n166 163.367
R227 B.n168 B.n167 163.367
R228 B.n168 B.n45 163.367
R229 B.n172 B.n45 163.367
R230 B.n173 B.n172 163.367
R231 B.n174 B.n173 163.367
R232 B.n174 B.n43 163.367
R233 B.n178 B.n43 163.367
R234 B.n179 B.n178 163.367
R235 B.n180 B.n179 163.367
R236 B.n180 B.n41 163.367
R237 B.n184 B.n41 163.367
R238 B.n185 B.n184 163.367
R239 B.n186 B.n185 163.367
R240 B.n186 B.n39 163.367
R241 B.n190 B.n39 163.367
R242 B.n191 B.n190 163.367
R243 B.n192 B.n191 163.367
R244 B.n192 B.n37 163.367
R245 B.n196 B.n37 163.367
R246 B.n197 B.n196 163.367
R247 B.n198 B.n197 163.367
R248 B.n198 B.n35 163.367
R249 B.n202 B.n35 163.367
R250 B.n203 B.n202 163.367
R251 B.n204 B.n203 163.367
R252 B.n266 B.n9 163.367
R253 B.n266 B.n265 163.367
R254 B.n265 B.n264 163.367
R255 B.n264 B.n11 163.367
R256 B.n260 B.n11 163.367
R257 B.n260 B.n259 163.367
R258 B.n259 B.n258 163.367
R259 B.n258 B.n13 163.367
R260 B.n254 B.n13 163.367
R261 B.n254 B.n253 163.367
R262 B.n253 B.n252 163.367
R263 B.n252 B.n15 163.367
R264 B.n248 B.n15 163.367
R265 B.n248 B.n247 163.367
R266 B.n247 B.n246 163.367
R267 B.n246 B.n17 163.367
R268 B.n241 B.n17 163.367
R269 B.n241 B.n240 163.367
R270 B.n240 B.n239 163.367
R271 B.n239 B.n21 163.367
R272 B.n235 B.n21 163.367
R273 B.n235 B.n234 163.367
R274 B.n234 B.n233 163.367
R275 B.n233 B.n23 163.367
R276 B.n228 B.n23 163.367
R277 B.n228 B.n227 163.367
R278 B.n227 B.n226 163.367
R279 B.n226 B.n27 163.367
R280 B.n222 B.n27 163.367
R281 B.n222 B.n221 163.367
R282 B.n221 B.n220 163.367
R283 B.n220 B.n29 163.367
R284 B.n216 B.n29 163.367
R285 B.n216 B.n215 163.367
R286 B.n215 B.n214 163.367
R287 B.n214 B.n31 163.367
R288 B.n210 B.n31 163.367
R289 B.n210 B.n209 163.367
R290 B.n209 B.n208 163.367
R291 B.n208 B.n33 163.367
R292 B.n58 B.n57 59.5399
R293 B.n123 B.n65 59.5399
R294 B.n244 B.n19 59.5399
R295 B.n230 B.n25 59.5399
R296 B.n269 B.n268 31.6883
R297 B.n206 B.n205 31.6883
R298 B.n163 B.n48 31.6883
R299 B.n99 B.n98 31.6883
R300 B B.n291 18.0485
R301 B.n268 B.n267 10.6151
R302 B.n267 B.n10 10.6151
R303 B.n263 B.n10 10.6151
R304 B.n263 B.n262 10.6151
R305 B.n262 B.n261 10.6151
R306 B.n261 B.n12 10.6151
R307 B.n257 B.n12 10.6151
R308 B.n257 B.n256 10.6151
R309 B.n256 B.n255 10.6151
R310 B.n255 B.n14 10.6151
R311 B.n251 B.n14 10.6151
R312 B.n251 B.n250 10.6151
R313 B.n250 B.n249 10.6151
R314 B.n249 B.n16 10.6151
R315 B.n245 B.n16 10.6151
R316 B.n243 B.n242 10.6151
R317 B.n242 B.n20 10.6151
R318 B.n238 B.n20 10.6151
R319 B.n238 B.n237 10.6151
R320 B.n237 B.n236 10.6151
R321 B.n236 B.n22 10.6151
R322 B.n232 B.n22 10.6151
R323 B.n232 B.n231 10.6151
R324 B.n229 B.n26 10.6151
R325 B.n225 B.n26 10.6151
R326 B.n225 B.n224 10.6151
R327 B.n224 B.n223 10.6151
R328 B.n223 B.n28 10.6151
R329 B.n219 B.n28 10.6151
R330 B.n219 B.n218 10.6151
R331 B.n218 B.n217 10.6151
R332 B.n217 B.n30 10.6151
R333 B.n213 B.n30 10.6151
R334 B.n213 B.n212 10.6151
R335 B.n212 B.n211 10.6151
R336 B.n211 B.n32 10.6151
R337 B.n207 B.n32 10.6151
R338 B.n207 B.n206 10.6151
R339 B.n164 B.n163 10.6151
R340 B.n165 B.n164 10.6151
R341 B.n165 B.n46 10.6151
R342 B.n169 B.n46 10.6151
R343 B.n170 B.n169 10.6151
R344 B.n171 B.n170 10.6151
R345 B.n171 B.n44 10.6151
R346 B.n175 B.n44 10.6151
R347 B.n176 B.n175 10.6151
R348 B.n177 B.n176 10.6151
R349 B.n177 B.n42 10.6151
R350 B.n181 B.n42 10.6151
R351 B.n182 B.n181 10.6151
R352 B.n183 B.n182 10.6151
R353 B.n183 B.n40 10.6151
R354 B.n187 B.n40 10.6151
R355 B.n188 B.n187 10.6151
R356 B.n189 B.n188 10.6151
R357 B.n189 B.n38 10.6151
R358 B.n193 B.n38 10.6151
R359 B.n194 B.n193 10.6151
R360 B.n195 B.n194 10.6151
R361 B.n195 B.n36 10.6151
R362 B.n199 B.n36 10.6151
R363 B.n200 B.n199 10.6151
R364 B.n201 B.n200 10.6151
R365 B.n201 B.n34 10.6151
R366 B.n205 B.n34 10.6151
R367 B.n99 B.n72 10.6151
R368 B.n103 B.n72 10.6151
R369 B.n104 B.n103 10.6151
R370 B.n105 B.n104 10.6151
R371 B.n105 B.n70 10.6151
R372 B.n109 B.n70 10.6151
R373 B.n110 B.n109 10.6151
R374 B.n111 B.n110 10.6151
R375 B.n111 B.n68 10.6151
R376 B.n115 B.n68 10.6151
R377 B.n116 B.n115 10.6151
R378 B.n117 B.n116 10.6151
R379 B.n117 B.n66 10.6151
R380 B.n121 B.n66 10.6151
R381 B.n122 B.n121 10.6151
R382 B.n124 B.n62 10.6151
R383 B.n128 B.n62 10.6151
R384 B.n129 B.n128 10.6151
R385 B.n130 B.n129 10.6151
R386 B.n130 B.n60 10.6151
R387 B.n134 B.n60 10.6151
R388 B.n135 B.n134 10.6151
R389 B.n136 B.n135 10.6151
R390 B.n140 B.n139 10.6151
R391 B.n141 B.n140 10.6151
R392 B.n141 B.n54 10.6151
R393 B.n145 B.n54 10.6151
R394 B.n146 B.n145 10.6151
R395 B.n147 B.n146 10.6151
R396 B.n147 B.n52 10.6151
R397 B.n151 B.n52 10.6151
R398 B.n152 B.n151 10.6151
R399 B.n153 B.n152 10.6151
R400 B.n153 B.n50 10.6151
R401 B.n157 B.n50 10.6151
R402 B.n158 B.n157 10.6151
R403 B.n159 B.n158 10.6151
R404 B.n159 B.n48 10.6151
R405 B.n98 B.n97 10.6151
R406 B.n97 B.n74 10.6151
R407 B.n93 B.n74 10.6151
R408 B.n93 B.n92 10.6151
R409 B.n92 B.n91 10.6151
R410 B.n91 B.n76 10.6151
R411 B.n87 B.n76 10.6151
R412 B.n87 B.n86 10.6151
R413 B.n86 B.n85 10.6151
R414 B.n85 B.n78 10.6151
R415 B.n81 B.n78 10.6151
R416 B.n81 B.n80 10.6151
R417 B.n80 B.n0 10.6151
R418 B.n287 B.n1 10.6151
R419 B.n287 B.n286 10.6151
R420 B.n286 B.n285 10.6151
R421 B.n285 B.n4 10.6151
R422 B.n281 B.n4 10.6151
R423 B.n281 B.n280 10.6151
R424 B.n280 B.n279 10.6151
R425 B.n279 B.n6 10.6151
R426 B.n275 B.n6 10.6151
R427 B.n275 B.n274 10.6151
R428 B.n274 B.n273 10.6151
R429 B.n273 B.n8 10.6151
R430 B.n269 B.n8 10.6151
R431 B.n57 B.n56 9.89141
R432 B.n65 B.n64 9.89141
R433 B.n19 B.n18 9.89141
R434 B.n25 B.n24 9.89141
R435 B.n244 B.n243 6.5566
R436 B.n231 B.n230 6.5566
R437 B.n124 B.n123 6.5566
R438 B.n136 B.n58 6.5566
R439 B.n245 B.n244 4.05904
R440 B.n230 B.n229 4.05904
R441 B.n123 B.n122 4.05904
R442 B.n139 B.n58 4.05904
R443 B.n291 B.n0 2.81026
R444 B.n291 B.n1 2.81026
R445 VP.n7 VP.t3 632.442
R446 VP.n5 VP.t0 632.442
R447 VP.n0 VP.t1 632.442
R448 VP.n2 VP.t4 632.442
R449 VP.n6 VP.t5 594.467
R450 VP.n1 VP.t2 594.467
R451 VP.n3 VP.n0 161.489
R452 VP.n8 VP.n7 161.3
R453 VP.n3 VP.n2 161.3
R454 VP.n5 VP.n4 161.3
R455 VP.n6 VP.n5 36.5157
R456 VP.n7 VP.n6 36.5157
R457 VP.n1 VP.n0 36.5157
R458 VP.n2 VP.n1 36.5157
R459 VP.n4 VP.n3 32.4891
R460 VP.n8 VP.n4 0.189894
R461 VP VP.n8 0.0516364
R462 VTAIL.n66 VTAIL.n56 756.745
R463 VTAIL.n12 VTAIL.n2 756.745
R464 VTAIL.n50 VTAIL.n40 756.745
R465 VTAIL.n32 VTAIL.n22 756.745
R466 VTAIL.n60 VTAIL.n59 585
R467 VTAIL.n65 VTAIL.n64 585
R468 VTAIL.n67 VTAIL.n66 585
R469 VTAIL.n6 VTAIL.n5 585
R470 VTAIL.n11 VTAIL.n10 585
R471 VTAIL.n13 VTAIL.n12 585
R472 VTAIL.n51 VTAIL.n50 585
R473 VTAIL.n49 VTAIL.n48 585
R474 VTAIL.n44 VTAIL.n43 585
R475 VTAIL.n33 VTAIL.n32 585
R476 VTAIL.n31 VTAIL.n30 585
R477 VTAIL.n26 VTAIL.n25 585
R478 VTAIL.n61 VTAIL.t0 336.901
R479 VTAIL.n7 VTAIL.t9 336.901
R480 VTAIL.n45 VTAIL.t10 336.901
R481 VTAIL.n27 VTAIL.t3 336.901
R482 VTAIL.n65 VTAIL.n59 171.744
R483 VTAIL.n66 VTAIL.n65 171.744
R484 VTAIL.n11 VTAIL.n5 171.744
R485 VTAIL.n12 VTAIL.n11 171.744
R486 VTAIL.n50 VTAIL.n49 171.744
R487 VTAIL.n49 VTAIL.n43 171.744
R488 VTAIL.n32 VTAIL.n31 171.744
R489 VTAIL.n31 VTAIL.n25 171.744
R490 VTAIL.n39 VTAIL.n38 111.367
R491 VTAIL.n21 VTAIL.n20 111.367
R492 VTAIL.n1 VTAIL.n0 111.365
R493 VTAIL.n19 VTAIL.n18 111.365
R494 VTAIL.t0 VTAIL.n59 85.8723
R495 VTAIL.t9 VTAIL.n5 85.8723
R496 VTAIL.t10 VTAIL.n43 85.8723
R497 VTAIL.t3 VTAIL.n25 85.8723
R498 VTAIL.n71 VTAIL.n70 32.3793
R499 VTAIL.n17 VTAIL.n16 32.3793
R500 VTAIL.n55 VTAIL.n54 32.3793
R501 VTAIL.n37 VTAIL.n36 32.3793
R502 VTAIL.n61 VTAIL.n60 16.193
R503 VTAIL.n7 VTAIL.n6 16.193
R504 VTAIL.n45 VTAIL.n44 16.193
R505 VTAIL.n27 VTAIL.n26 16.193
R506 VTAIL.n21 VTAIL.n19 15.9445
R507 VTAIL.n71 VTAIL.n55 15.5048
R508 VTAIL.n64 VTAIL.n63 12.8005
R509 VTAIL.n10 VTAIL.n9 12.8005
R510 VTAIL.n48 VTAIL.n47 12.8005
R511 VTAIL.n30 VTAIL.n29 12.8005
R512 VTAIL.n67 VTAIL.n58 12.0247
R513 VTAIL.n13 VTAIL.n4 12.0247
R514 VTAIL.n51 VTAIL.n42 12.0247
R515 VTAIL.n33 VTAIL.n24 12.0247
R516 VTAIL.n68 VTAIL.n56 11.249
R517 VTAIL.n14 VTAIL.n2 11.249
R518 VTAIL.n52 VTAIL.n40 11.249
R519 VTAIL.n34 VTAIL.n22 11.249
R520 VTAIL.n0 VTAIL.t4 10.3855
R521 VTAIL.n0 VTAIL.t1 10.3855
R522 VTAIL.n18 VTAIL.t7 10.3855
R523 VTAIL.n18 VTAIL.t11 10.3855
R524 VTAIL.n38 VTAIL.t6 10.3855
R525 VTAIL.n38 VTAIL.t8 10.3855
R526 VTAIL.n20 VTAIL.t2 10.3855
R527 VTAIL.n20 VTAIL.t5 10.3855
R528 VTAIL.n70 VTAIL.n69 9.45567
R529 VTAIL.n16 VTAIL.n15 9.45567
R530 VTAIL.n54 VTAIL.n53 9.45567
R531 VTAIL.n36 VTAIL.n35 9.45567
R532 VTAIL.n69 VTAIL.n68 9.3005
R533 VTAIL.n58 VTAIL.n57 9.3005
R534 VTAIL.n63 VTAIL.n62 9.3005
R535 VTAIL.n15 VTAIL.n14 9.3005
R536 VTAIL.n4 VTAIL.n3 9.3005
R537 VTAIL.n9 VTAIL.n8 9.3005
R538 VTAIL.n53 VTAIL.n52 9.3005
R539 VTAIL.n42 VTAIL.n41 9.3005
R540 VTAIL.n47 VTAIL.n46 9.3005
R541 VTAIL.n35 VTAIL.n34 9.3005
R542 VTAIL.n24 VTAIL.n23 9.3005
R543 VTAIL.n29 VTAIL.n28 9.3005
R544 VTAIL.n46 VTAIL.n45 3.91276
R545 VTAIL.n28 VTAIL.n27 3.91276
R546 VTAIL.n62 VTAIL.n61 3.91276
R547 VTAIL.n8 VTAIL.n7 3.91276
R548 VTAIL.n70 VTAIL.n56 2.71565
R549 VTAIL.n16 VTAIL.n2 2.71565
R550 VTAIL.n54 VTAIL.n40 2.71565
R551 VTAIL.n36 VTAIL.n22 2.71565
R552 VTAIL.n68 VTAIL.n67 1.93989
R553 VTAIL.n14 VTAIL.n13 1.93989
R554 VTAIL.n52 VTAIL.n51 1.93989
R555 VTAIL.n34 VTAIL.n33 1.93989
R556 VTAIL.n64 VTAIL.n58 1.16414
R557 VTAIL.n10 VTAIL.n4 1.16414
R558 VTAIL.n48 VTAIL.n42 1.16414
R559 VTAIL.n30 VTAIL.n24 1.16414
R560 VTAIL.n39 VTAIL.n37 0.690155
R561 VTAIL.n17 VTAIL.n1 0.690155
R562 VTAIL.n37 VTAIL.n21 0.440155
R563 VTAIL.n55 VTAIL.n39 0.440155
R564 VTAIL.n19 VTAIL.n17 0.440155
R565 VTAIL.n63 VTAIL.n60 0.388379
R566 VTAIL.n9 VTAIL.n6 0.388379
R567 VTAIL.n47 VTAIL.n44 0.388379
R568 VTAIL.n29 VTAIL.n26 0.388379
R569 VTAIL VTAIL.n71 0.272052
R570 VTAIL VTAIL.n1 0.168603
R571 VTAIL.n62 VTAIL.n57 0.155672
R572 VTAIL.n69 VTAIL.n57 0.155672
R573 VTAIL.n8 VTAIL.n3 0.155672
R574 VTAIL.n15 VTAIL.n3 0.155672
R575 VTAIL.n53 VTAIL.n41 0.155672
R576 VTAIL.n46 VTAIL.n41 0.155672
R577 VTAIL.n35 VTAIL.n23 0.155672
R578 VTAIL.n28 VTAIL.n23 0.155672
R579 VDD1.n10 VDD1.n0 756.745
R580 VDD1.n25 VDD1.n15 756.745
R581 VDD1.n11 VDD1.n10 585
R582 VDD1.n9 VDD1.n8 585
R583 VDD1.n4 VDD1.n3 585
R584 VDD1.n19 VDD1.n18 585
R585 VDD1.n24 VDD1.n23 585
R586 VDD1.n26 VDD1.n25 585
R587 VDD1.n5 VDD1.t4 336.901
R588 VDD1.n20 VDD1.t5 336.901
R589 VDD1.n10 VDD1.n9 171.744
R590 VDD1.n9 VDD1.n3 171.744
R591 VDD1.n24 VDD1.n18 171.744
R592 VDD1.n25 VDD1.n24 171.744
R593 VDD1.n31 VDD1.n30 128.1
R594 VDD1.n33 VDD1.n32 128.044
R595 VDD1.t4 VDD1.n3 85.8723
R596 VDD1.t5 VDD1.n18 85.8723
R597 VDD1 VDD1.n14 49.446
R598 VDD1.n31 VDD1.n29 49.3325
R599 VDD1.n33 VDD1.n31 28.6453
R600 VDD1.n5 VDD1.n4 16.193
R601 VDD1.n20 VDD1.n19 16.193
R602 VDD1.n8 VDD1.n7 12.8005
R603 VDD1.n23 VDD1.n22 12.8005
R604 VDD1.n11 VDD1.n2 12.0247
R605 VDD1.n26 VDD1.n17 12.0247
R606 VDD1.n12 VDD1.n0 11.249
R607 VDD1.n27 VDD1.n15 11.249
R608 VDD1.n32 VDD1.t3 10.3855
R609 VDD1.n32 VDD1.t1 10.3855
R610 VDD1.n30 VDD1.t0 10.3855
R611 VDD1.n30 VDD1.t2 10.3855
R612 VDD1.n14 VDD1.n13 9.45567
R613 VDD1.n29 VDD1.n28 9.45567
R614 VDD1.n13 VDD1.n12 9.3005
R615 VDD1.n2 VDD1.n1 9.3005
R616 VDD1.n7 VDD1.n6 9.3005
R617 VDD1.n28 VDD1.n27 9.3005
R618 VDD1.n17 VDD1.n16 9.3005
R619 VDD1.n22 VDD1.n21 9.3005
R620 VDD1.n6 VDD1.n5 3.91276
R621 VDD1.n21 VDD1.n20 3.91276
R622 VDD1.n14 VDD1.n0 2.71565
R623 VDD1.n29 VDD1.n15 2.71565
R624 VDD1.n12 VDD1.n11 1.93989
R625 VDD1.n27 VDD1.n26 1.93989
R626 VDD1.n8 VDD1.n2 1.16414
R627 VDD1.n23 VDD1.n17 1.16414
R628 VDD1.n7 VDD1.n4 0.388379
R629 VDD1.n22 VDD1.n19 0.388379
R630 VDD1.n13 VDD1.n1 0.155672
R631 VDD1.n6 VDD1.n1 0.155672
R632 VDD1.n21 VDD1.n16 0.155672
R633 VDD1.n28 VDD1.n16 0.155672
R634 VDD1 VDD1.n33 0.0522241
R635 VN.n2 VN.t5 632.442
R636 VN.n0 VN.t1 632.442
R637 VN.n6 VN.t3 632.442
R638 VN.n4 VN.t0 632.442
R639 VN.n1 VN.t4 594.467
R640 VN.n5 VN.t2 594.467
R641 VN.n7 VN.n4 161.489
R642 VN.n3 VN.n0 161.489
R643 VN.n3 VN.n2 161.3
R644 VN.n7 VN.n6 161.3
R645 VN.n1 VN.n0 36.5157
R646 VN.n2 VN.n1 36.5157
R647 VN.n6 VN.n5 36.5157
R648 VN.n5 VN.n4 36.5157
R649 VN VN.n7 32.8698
R650 VN VN.n3 0.0516364
R651 VDD2.n27 VDD2.n17 756.745
R652 VDD2.n10 VDD2.n0 756.745
R653 VDD2.n28 VDD2.n27 585
R654 VDD2.n26 VDD2.n25 585
R655 VDD2.n21 VDD2.n20 585
R656 VDD2.n4 VDD2.n3 585
R657 VDD2.n9 VDD2.n8 585
R658 VDD2.n11 VDD2.n10 585
R659 VDD2.n22 VDD2.t2 336.901
R660 VDD2.n5 VDD2.t4 336.901
R661 VDD2.n27 VDD2.n26 171.744
R662 VDD2.n26 VDD2.n20 171.744
R663 VDD2.n9 VDD2.n3 171.744
R664 VDD2.n10 VDD2.n9 171.744
R665 VDD2.n16 VDD2.n15 128.1
R666 VDD2 VDD2.n33 128.096
R667 VDD2.t2 VDD2.n20 85.8723
R668 VDD2.t4 VDD2.n3 85.8723
R669 VDD2.n16 VDD2.n14 49.3325
R670 VDD2.n32 VDD2.n31 49.0581
R671 VDD2.n32 VDD2.n16 27.8424
R672 VDD2.n22 VDD2.n21 16.193
R673 VDD2.n5 VDD2.n4 16.193
R674 VDD2.n25 VDD2.n24 12.8005
R675 VDD2.n8 VDD2.n7 12.8005
R676 VDD2.n28 VDD2.n19 12.0247
R677 VDD2.n11 VDD2.n2 12.0247
R678 VDD2.n29 VDD2.n17 11.249
R679 VDD2.n12 VDD2.n0 11.249
R680 VDD2.n33 VDD2.t3 10.3855
R681 VDD2.n33 VDD2.t5 10.3855
R682 VDD2.n15 VDD2.t1 10.3855
R683 VDD2.n15 VDD2.t0 10.3855
R684 VDD2.n31 VDD2.n30 9.45567
R685 VDD2.n14 VDD2.n13 9.45567
R686 VDD2.n30 VDD2.n29 9.3005
R687 VDD2.n19 VDD2.n18 9.3005
R688 VDD2.n24 VDD2.n23 9.3005
R689 VDD2.n13 VDD2.n12 9.3005
R690 VDD2.n2 VDD2.n1 9.3005
R691 VDD2.n7 VDD2.n6 9.3005
R692 VDD2.n23 VDD2.n22 3.91276
R693 VDD2.n6 VDD2.n5 3.91276
R694 VDD2.n31 VDD2.n17 2.71565
R695 VDD2.n14 VDD2.n0 2.71565
R696 VDD2.n29 VDD2.n28 1.93989
R697 VDD2.n12 VDD2.n11 1.93989
R698 VDD2.n25 VDD2.n19 1.16414
R699 VDD2.n8 VDD2.n2 1.16414
R700 VDD2 VDD2.n32 0.388431
R701 VDD2.n24 VDD2.n21 0.388379
R702 VDD2.n7 VDD2.n4 0.388379
R703 VDD2.n30 VDD2.n18 0.155672
R704 VDD2.n23 VDD2.n18 0.155672
R705 VDD2.n6 VDD2.n1 0.155672
R706 VDD2.n13 VDD2.n1 0.155672
C0 VP w_n1378_n1594# 2.01557f
C1 VDD2 VN 0.75304f
C2 VP VTAIL 0.695638f
C3 VDD1 B 0.775824f
C4 VDD1 w_n1378_n1594# 0.977408f
C5 B VN 0.539605f
C6 VDD2 B 0.793628f
C7 VDD1 VTAIL 5.54115f
C8 VN w_n1378_n1594# 1.84627f
C9 VDD2 w_n1378_n1594# 0.98575f
C10 VTAIL VN 0.681346f
C11 VDD2 VTAIL 5.57593f
C12 VDD1 VP 0.856348f
C13 B w_n1378_n1594# 3.9022f
C14 VP VN 2.94112f
C15 VTAIL B 0.92813f
C16 VP VDD2 0.257281f
C17 VTAIL w_n1378_n1594# 1.47862f
C18 VDD1 VN 0.152121f
C19 VP B 0.813225f
C20 VDD1 VDD2 0.525582f
C21 VDD2 VSUBS 0.816135f
C22 VDD1 VSUBS 0.671882f
C23 VTAIL VSUBS 0.281363f
C24 VN VSUBS 2.26273f
C25 VP VSUBS 0.675971f
C26 B VSUBS 1.428702f
C27 w_n1378_n1594# VSUBS 27.797f
C28 VDD2.n0 VSUBS 0.027276f
C29 VDD2.n1 VSUBS 0.026455f
C30 VDD2.n2 VSUBS 0.014216f
C31 VDD2.n3 VSUBS 0.025201f
C32 VDD2.n4 VSUBS 0.020744f
C33 VDD2.t4 VSUBS 0.074085f
C34 VDD2.n5 VSUBS 0.094768f
C35 VDD2.n6 VSUBS 0.260431f
C36 VDD2.n7 VSUBS 0.014216f
C37 VDD2.n8 VSUBS 0.015052f
C38 VDD2.n9 VSUBS 0.033601f
C39 VDD2.n10 VSUBS 0.075238f
C40 VDD2.n11 VSUBS 0.015052f
C41 VDD2.n12 VSUBS 0.014216f
C42 VDD2.n13 VSUBS 0.061511f
C43 VDD2.n14 VSUBS 0.056267f
C44 VDD2.t1 VSUBS 0.065435f
C45 VDD2.t0 VSUBS 0.065435f
C46 VDD2.n15 VSUBS 0.350815f
C47 VDD2.n16 VSUBS 1.29627f
C48 VDD2.n17 VSUBS 0.027276f
C49 VDD2.n18 VSUBS 0.026455f
C50 VDD2.n19 VSUBS 0.014216f
C51 VDD2.n20 VSUBS 0.025201f
C52 VDD2.n21 VSUBS 0.020744f
C53 VDD2.t2 VSUBS 0.074085f
C54 VDD2.n22 VSUBS 0.094768f
C55 VDD2.n23 VSUBS 0.260431f
C56 VDD2.n24 VSUBS 0.014216f
C57 VDD2.n25 VSUBS 0.015052f
C58 VDD2.n26 VSUBS 0.033601f
C59 VDD2.n27 VSUBS 0.075238f
C60 VDD2.n28 VSUBS 0.015052f
C61 VDD2.n29 VSUBS 0.014216f
C62 VDD2.n30 VSUBS 0.061511f
C63 VDD2.n31 VSUBS 0.05584f
C64 VDD2.n32 VSUBS 1.255f
C65 VDD2.t3 VSUBS 0.065435f
C66 VDD2.t5 VSUBS 0.065435f
C67 VDD2.n33 VSUBS 0.350802f
C68 VN.t1 VSUBS 0.066838f
C69 VN.n0 VSUBS 0.051189f
C70 VN.t4 VSUBS 0.064424f
C71 VN.n1 VSUBS 0.041665f
C72 VN.t5 VSUBS 0.066838f
C73 VN.n2 VSUBS 0.051137f
C74 VN.n3 VSUBS 0.074927f
C75 VN.t0 VSUBS 0.066838f
C76 VN.n4 VSUBS 0.051189f
C77 VN.t3 VSUBS 0.066838f
C78 VN.t2 VSUBS 0.064424f
C79 VN.n5 VSUBS 0.041665f
C80 VN.n6 VSUBS 0.051137f
C81 VN.n7 VSUBS 1.0847f
C82 VDD1.n0 VSUBS 0.026329f
C83 VDD1.n1 VSUBS 0.025537f
C84 VDD1.n2 VSUBS 0.013722f
C85 VDD1.n3 VSUBS 0.024326f
C86 VDD1.n4 VSUBS 0.020024f
C87 VDD1.t4 VSUBS 0.071514f
C88 VDD1.n5 VSUBS 0.091479f
C89 VDD1.n6 VSUBS 0.251394f
C90 VDD1.n7 VSUBS 0.013722f
C91 VDD1.n8 VSUBS 0.01453f
C92 VDD1.n9 VSUBS 0.032435f
C93 VDD1.n10 VSUBS 0.072627f
C94 VDD1.n11 VSUBS 0.01453f
C95 VDD1.n12 VSUBS 0.013722f
C96 VDD1.n13 VSUBS 0.059377f
C97 VDD1.n14 VSUBS 0.05454f
C98 VDD1.n15 VSUBS 0.026329f
C99 VDD1.n16 VSUBS 0.025537f
C100 VDD1.n17 VSUBS 0.013722f
C101 VDD1.n18 VSUBS 0.024326f
C102 VDD1.n19 VSUBS 0.020024f
C103 VDD1.t5 VSUBS 0.071514f
C104 VDD1.n20 VSUBS 0.091479f
C105 VDD1.n21 VSUBS 0.251394f
C106 VDD1.n22 VSUBS 0.013722f
C107 VDD1.n23 VSUBS 0.01453f
C108 VDD1.n24 VSUBS 0.032435f
C109 VDD1.n25 VSUBS 0.072627f
C110 VDD1.n26 VSUBS 0.01453f
C111 VDD1.n27 VSUBS 0.013722f
C112 VDD1.n28 VSUBS 0.059377f
C113 VDD1.n29 VSUBS 0.054315f
C114 VDD1.t0 VSUBS 0.063164f
C115 VDD1.t2 VSUBS 0.063164f
C116 VDD1.n30 VSUBS 0.338642f
C117 VDD1.n31 VSUBS 1.3157f
C118 VDD1.t3 VSUBS 0.063164f
C119 VDD1.t1 VSUBS 0.063164f
C120 VDD1.n32 VSUBS 0.338476f
C121 VDD1.n33 VSUBS 1.53829f
C122 VTAIL.t4 VSUBS 0.075765f
C123 VTAIL.t1 VSUBS 0.075765f
C124 VTAIL.n0 VSUBS 0.34804f
C125 VTAIL.n1 VSUBS 0.493852f
C126 VTAIL.n2 VSUBS 0.031582f
C127 VTAIL.n3 VSUBS 0.030632f
C128 VTAIL.n4 VSUBS 0.01646f
C129 VTAIL.n5 VSUBS 0.02918f
C130 VTAIL.n6 VSUBS 0.024019f
C131 VTAIL.t9 VSUBS 0.085781f
C132 VTAIL.n7 VSUBS 0.10973f
C133 VTAIL.n8 VSUBS 0.301548f
C134 VTAIL.n9 VSUBS 0.01646f
C135 VTAIL.n10 VSUBS 0.017428f
C136 VTAIL.n11 VSUBS 0.038906f
C137 VTAIL.n12 VSUBS 0.087116f
C138 VTAIL.n13 VSUBS 0.017428f
C139 VTAIL.n14 VSUBS 0.01646f
C140 VTAIL.n15 VSUBS 0.071222f
C141 VTAIL.n16 VSUBS 0.043509f
C142 VTAIL.n17 VSUBS 0.137864f
C143 VTAIL.t7 VSUBS 0.075765f
C144 VTAIL.t11 VSUBS 0.075765f
C145 VTAIL.n18 VSUBS 0.34804f
C146 VTAIL.n19 VSUBS 1.2218f
C147 VTAIL.t2 VSUBS 0.075765f
C148 VTAIL.t5 VSUBS 0.075765f
C149 VTAIL.n20 VSUBS 0.348043f
C150 VTAIL.n21 VSUBS 1.2218f
C151 VTAIL.n22 VSUBS 0.031582f
C152 VTAIL.n23 VSUBS 0.030632f
C153 VTAIL.n24 VSUBS 0.01646f
C154 VTAIL.n25 VSUBS 0.02918f
C155 VTAIL.n26 VSUBS 0.024019f
C156 VTAIL.t3 VSUBS 0.085781f
C157 VTAIL.n27 VSUBS 0.10973f
C158 VTAIL.n28 VSUBS 0.301548f
C159 VTAIL.n29 VSUBS 0.01646f
C160 VTAIL.n30 VSUBS 0.017428f
C161 VTAIL.n31 VSUBS 0.038906f
C162 VTAIL.n32 VSUBS 0.087116f
C163 VTAIL.n33 VSUBS 0.017428f
C164 VTAIL.n34 VSUBS 0.01646f
C165 VTAIL.n35 VSUBS 0.071222f
C166 VTAIL.n36 VSUBS 0.043509f
C167 VTAIL.n37 VSUBS 0.137864f
C168 VTAIL.t6 VSUBS 0.075765f
C169 VTAIL.t8 VSUBS 0.075765f
C170 VTAIL.n38 VSUBS 0.348043f
C171 VTAIL.n39 VSUBS 0.520652f
C172 VTAIL.n40 VSUBS 0.031582f
C173 VTAIL.n41 VSUBS 0.030632f
C174 VTAIL.n42 VSUBS 0.01646f
C175 VTAIL.n43 VSUBS 0.02918f
C176 VTAIL.n44 VSUBS 0.024019f
C177 VTAIL.t10 VSUBS 0.085781f
C178 VTAIL.n45 VSUBS 0.10973f
C179 VTAIL.n46 VSUBS 0.301548f
C180 VTAIL.n47 VSUBS 0.01646f
C181 VTAIL.n48 VSUBS 0.017428f
C182 VTAIL.n49 VSUBS 0.038906f
C183 VTAIL.n50 VSUBS 0.087116f
C184 VTAIL.n51 VSUBS 0.017428f
C185 VTAIL.n52 VSUBS 0.01646f
C186 VTAIL.n53 VSUBS 0.071222f
C187 VTAIL.n54 VSUBS 0.043509f
C188 VTAIL.n55 VSUBS 0.795613f
C189 VTAIL.n56 VSUBS 0.031582f
C190 VTAIL.n57 VSUBS 0.030632f
C191 VTAIL.n58 VSUBS 0.01646f
C192 VTAIL.n59 VSUBS 0.02918f
C193 VTAIL.n60 VSUBS 0.024019f
C194 VTAIL.t0 VSUBS 0.085781f
C195 VTAIL.n61 VSUBS 0.10973f
C196 VTAIL.n62 VSUBS 0.301548f
C197 VTAIL.n63 VSUBS 0.01646f
C198 VTAIL.n64 VSUBS 0.017428f
C199 VTAIL.n65 VSUBS 0.038906f
C200 VTAIL.n66 VSUBS 0.087116f
C201 VTAIL.n67 VSUBS 0.017428f
C202 VTAIL.n68 VSUBS 0.01646f
C203 VTAIL.n69 VSUBS 0.071222f
C204 VTAIL.n70 VSUBS 0.043509f
C205 VTAIL.n71 VSUBS 0.77902f
C206 VP.t1 VSUBS 0.115138f
C207 VP.n0 VSUBS 0.08818f
C208 VP.t2 VSUBS 0.110979f
C209 VP.n1 VSUBS 0.071774f
C210 VP.t4 VSUBS 0.115138f
C211 VP.n2 VSUBS 0.08809f
C212 VP.n3 VSUBS 1.82306f
C213 VP.n4 VSUBS 1.822f
C214 VP.t5 VSUBS 0.110979f
C215 VP.t0 VSUBS 0.115138f
C216 VP.n5 VSUBS 0.08809f
C217 VP.n6 VSUBS 0.071774f
C218 VP.t3 VSUBS 0.115138f
C219 VP.n7 VSUBS 0.08809f
C220 VP.n8 VSUBS 0.05273f
C221 B.n0 VSUBS 0.005173f
C222 B.n1 VSUBS 0.005173f
C223 B.n2 VSUBS 0.00818f
C224 B.n3 VSUBS 0.00818f
C225 B.n4 VSUBS 0.00818f
C226 B.n5 VSUBS 0.00818f
C227 B.n6 VSUBS 0.00818f
C228 B.n7 VSUBS 0.00818f
C229 B.n8 VSUBS 0.00818f
C230 B.n9 VSUBS 0.019482f
C231 B.n10 VSUBS 0.00818f
C232 B.n11 VSUBS 0.00818f
C233 B.n12 VSUBS 0.00818f
C234 B.n13 VSUBS 0.00818f
C235 B.n14 VSUBS 0.00818f
C236 B.n15 VSUBS 0.00818f
C237 B.n16 VSUBS 0.00818f
C238 B.n17 VSUBS 0.00818f
C239 B.t2 VSUBS 0.053707f
C240 B.t1 VSUBS 0.057468f
C241 B.t0 VSUBS 0.027549f
C242 B.n18 VSUBS 0.102114f
C243 B.n19 VSUBS 0.100704f
C244 B.n20 VSUBS 0.00818f
C245 B.n21 VSUBS 0.00818f
C246 B.n22 VSUBS 0.00818f
C247 B.n23 VSUBS 0.00818f
C248 B.t8 VSUBS 0.053707f
C249 B.t7 VSUBS 0.057469f
C250 B.t6 VSUBS 0.027549f
C251 B.n24 VSUBS 0.102113f
C252 B.n25 VSUBS 0.100703f
C253 B.n26 VSUBS 0.00818f
C254 B.n27 VSUBS 0.00818f
C255 B.n28 VSUBS 0.00818f
C256 B.n29 VSUBS 0.00818f
C257 B.n30 VSUBS 0.00818f
C258 B.n31 VSUBS 0.00818f
C259 B.n32 VSUBS 0.00818f
C260 B.n33 VSUBS 0.019482f
C261 B.n34 VSUBS 0.00818f
C262 B.n35 VSUBS 0.00818f
C263 B.n36 VSUBS 0.00818f
C264 B.n37 VSUBS 0.00818f
C265 B.n38 VSUBS 0.00818f
C266 B.n39 VSUBS 0.00818f
C267 B.n40 VSUBS 0.00818f
C268 B.n41 VSUBS 0.00818f
C269 B.n42 VSUBS 0.00818f
C270 B.n43 VSUBS 0.00818f
C271 B.n44 VSUBS 0.00818f
C272 B.n45 VSUBS 0.00818f
C273 B.n46 VSUBS 0.00818f
C274 B.n47 VSUBS 0.00818f
C275 B.n48 VSUBS 0.019482f
C276 B.n49 VSUBS 0.00818f
C277 B.n50 VSUBS 0.00818f
C278 B.n51 VSUBS 0.00818f
C279 B.n52 VSUBS 0.00818f
C280 B.n53 VSUBS 0.00818f
C281 B.n54 VSUBS 0.00818f
C282 B.n55 VSUBS 0.00818f
C283 B.t4 VSUBS 0.053707f
C284 B.t5 VSUBS 0.057469f
C285 B.t3 VSUBS 0.027549f
C286 B.n56 VSUBS 0.102113f
C287 B.n57 VSUBS 0.100703f
C288 B.n58 VSUBS 0.018952f
C289 B.n59 VSUBS 0.00818f
C290 B.n60 VSUBS 0.00818f
C291 B.n61 VSUBS 0.00818f
C292 B.n62 VSUBS 0.00818f
C293 B.n63 VSUBS 0.00818f
C294 B.t10 VSUBS 0.053707f
C295 B.t11 VSUBS 0.057468f
C296 B.t9 VSUBS 0.027549f
C297 B.n64 VSUBS 0.102114f
C298 B.n65 VSUBS 0.100704f
C299 B.n66 VSUBS 0.00818f
C300 B.n67 VSUBS 0.00818f
C301 B.n68 VSUBS 0.00818f
C302 B.n69 VSUBS 0.00818f
C303 B.n70 VSUBS 0.00818f
C304 B.n71 VSUBS 0.00818f
C305 B.n72 VSUBS 0.00818f
C306 B.n73 VSUBS 0.018049f
C307 B.n74 VSUBS 0.00818f
C308 B.n75 VSUBS 0.00818f
C309 B.n76 VSUBS 0.00818f
C310 B.n77 VSUBS 0.00818f
C311 B.n78 VSUBS 0.00818f
C312 B.n79 VSUBS 0.00818f
C313 B.n80 VSUBS 0.00818f
C314 B.n81 VSUBS 0.00818f
C315 B.n82 VSUBS 0.00818f
C316 B.n83 VSUBS 0.00818f
C317 B.n84 VSUBS 0.00818f
C318 B.n85 VSUBS 0.00818f
C319 B.n86 VSUBS 0.00818f
C320 B.n87 VSUBS 0.00818f
C321 B.n88 VSUBS 0.00818f
C322 B.n89 VSUBS 0.00818f
C323 B.n90 VSUBS 0.00818f
C324 B.n91 VSUBS 0.00818f
C325 B.n92 VSUBS 0.00818f
C326 B.n93 VSUBS 0.00818f
C327 B.n94 VSUBS 0.00818f
C328 B.n95 VSUBS 0.00818f
C329 B.n96 VSUBS 0.00818f
C330 B.n97 VSUBS 0.00818f
C331 B.n98 VSUBS 0.018049f
C332 B.n99 VSUBS 0.019482f
C333 B.n100 VSUBS 0.019482f
C334 B.n101 VSUBS 0.00818f
C335 B.n102 VSUBS 0.00818f
C336 B.n103 VSUBS 0.00818f
C337 B.n104 VSUBS 0.00818f
C338 B.n105 VSUBS 0.00818f
C339 B.n106 VSUBS 0.00818f
C340 B.n107 VSUBS 0.00818f
C341 B.n108 VSUBS 0.00818f
C342 B.n109 VSUBS 0.00818f
C343 B.n110 VSUBS 0.00818f
C344 B.n111 VSUBS 0.00818f
C345 B.n112 VSUBS 0.00818f
C346 B.n113 VSUBS 0.00818f
C347 B.n114 VSUBS 0.00818f
C348 B.n115 VSUBS 0.00818f
C349 B.n116 VSUBS 0.00818f
C350 B.n117 VSUBS 0.00818f
C351 B.n118 VSUBS 0.00818f
C352 B.n119 VSUBS 0.00818f
C353 B.n120 VSUBS 0.00818f
C354 B.n121 VSUBS 0.00818f
C355 B.n122 VSUBS 0.005654f
C356 B.n123 VSUBS 0.018952f
C357 B.n124 VSUBS 0.006616f
C358 B.n125 VSUBS 0.00818f
C359 B.n126 VSUBS 0.00818f
C360 B.n127 VSUBS 0.00818f
C361 B.n128 VSUBS 0.00818f
C362 B.n129 VSUBS 0.00818f
C363 B.n130 VSUBS 0.00818f
C364 B.n131 VSUBS 0.00818f
C365 B.n132 VSUBS 0.00818f
C366 B.n133 VSUBS 0.00818f
C367 B.n134 VSUBS 0.00818f
C368 B.n135 VSUBS 0.00818f
C369 B.n136 VSUBS 0.006616f
C370 B.n137 VSUBS 0.00818f
C371 B.n138 VSUBS 0.00818f
C372 B.n139 VSUBS 0.005654f
C373 B.n140 VSUBS 0.00818f
C374 B.n141 VSUBS 0.00818f
C375 B.n142 VSUBS 0.00818f
C376 B.n143 VSUBS 0.00818f
C377 B.n144 VSUBS 0.00818f
C378 B.n145 VSUBS 0.00818f
C379 B.n146 VSUBS 0.00818f
C380 B.n147 VSUBS 0.00818f
C381 B.n148 VSUBS 0.00818f
C382 B.n149 VSUBS 0.00818f
C383 B.n150 VSUBS 0.00818f
C384 B.n151 VSUBS 0.00818f
C385 B.n152 VSUBS 0.00818f
C386 B.n153 VSUBS 0.00818f
C387 B.n154 VSUBS 0.00818f
C388 B.n155 VSUBS 0.00818f
C389 B.n156 VSUBS 0.00818f
C390 B.n157 VSUBS 0.00818f
C391 B.n158 VSUBS 0.00818f
C392 B.n159 VSUBS 0.00818f
C393 B.n160 VSUBS 0.00818f
C394 B.n161 VSUBS 0.019482f
C395 B.n162 VSUBS 0.018049f
C396 B.n163 VSUBS 0.018049f
C397 B.n164 VSUBS 0.00818f
C398 B.n165 VSUBS 0.00818f
C399 B.n166 VSUBS 0.00818f
C400 B.n167 VSUBS 0.00818f
C401 B.n168 VSUBS 0.00818f
C402 B.n169 VSUBS 0.00818f
C403 B.n170 VSUBS 0.00818f
C404 B.n171 VSUBS 0.00818f
C405 B.n172 VSUBS 0.00818f
C406 B.n173 VSUBS 0.00818f
C407 B.n174 VSUBS 0.00818f
C408 B.n175 VSUBS 0.00818f
C409 B.n176 VSUBS 0.00818f
C410 B.n177 VSUBS 0.00818f
C411 B.n178 VSUBS 0.00818f
C412 B.n179 VSUBS 0.00818f
C413 B.n180 VSUBS 0.00818f
C414 B.n181 VSUBS 0.00818f
C415 B.n182 VSUBS 0.00818f
C416 B.n183 VSUBS 0.00818f
C417 B.n184 VSUBS 0.00818f
C418 B.n185 VSUBS 0.00818f
C419 B.n186 VSUBS 0.00818f
C420 B.n187 VSUBS 0.00818f
C421 B.n188 VSUBS 0.00818f
C422 B.n189 VSUBS 0.00818f
C423 B.n190 VSUBS 0.00818f
C424 B.n191 VSUBS 0.00818f
C425 B.n192 VSUBS 0.00818f
C426 B.n193 VSUBS 0.00818f
C427 B.n194 VSUBS 0.00818f
C428 B.n195 VSUBS 0.00818f
C429 B.n196 VSUBS 0.00818f
C430 B.n197 VSUBS 0.00818f
C431 B.n198 VSUBS 0.00818f
C432 B.n199 VSUBS 0.00818f
C433 B.n200 VSUBS 0.00818f
C434 B.n201 VSUBS 0.00818f
C435 B.n202 VSUBS 0.00818f
C436 B.n203 VSUBS 0.00818f
C437 B.n204 VSUBS 0.018049f
C438 B.n205 VSUBS 0.019045f
C439 B.n206 VSUBS 0.018486f
C440 B.n207 VSUBS 0.00818f
C441 B.n208 VSUBS 0.00818f
C442 B.n209 VSUBS 0.00818f
C443 B.n210 VSUBS 0.00818f
C444 B.n211 VSUBS 0.00818f
C445 B.n212 VSUBS 0.00818f
C446 B.n213 VSUBS 0.00818f
C447 B.n214 VSUBS 0.00818f
C448 B.n215 VSUBS 0.00818f
C449 B.n216 VSUBS 0.00818f
C450 B.n217 VSUBS 0.00818f
C451 B.n218 VSUBS 0.00818f
C452 B.n219 VSUBS 0.00818f
C453 B.n220 VSUBS 0.00818f
C454 B.n221 VSUBS 0.00818f
C455 B.n222 VSUBS 0.00818f
C456 B.n223 VSUBS 0.00818f
C457 B.n224 VSUBS 0.00818f
C458 B.n225 VSUBS 0.00818f
C459 B.n226 VSUBS 0.00818f
C460 B.n227 VSUBS 0.00818f
C461 B.n228 VSUBS 0.00818f
C462 B.n229 VSUBS 0.005654f
C463 B.n230 VSUBS 0.018952f
C464 B.n231 VSUBS 0.006616f
C465 B.n232 VSUBS 0.00818f
C466 B.n233 VSUBS 0.00818f
C467 B.n234 VSUBS 0.00818f
C468 B.n235 VSUBS 0.00818f
C469 B.n236 VSUBS 0.00818f
C470 B.n237 VSUBS 0.00818f
C471 B.n238 VSUBS 0.00818f
C472 B.n239 VSUBS 0.00818f
C473 B.n240 VSUBS 0.00818f
C474 B.n241 VSUBS 0.00818f
C475 B.n242 VSUBS 0.00818f
C476 B.n243 VSUBS 0.006616f
C477 B.n244 VSUBS 0.018952f
C478 B.n245 VSUBS 0.005654f
C479 B.n246 VSUBS 0.00818f
C480 B.n247 VSUBS 0.00818f
C481 B.n248 VSUBS 0.00818f
C482 B.n249 VSUBS 0.00818f
C483 B.n250 VSUBS 0.00818f
C484 B.n251 VSUBS 0.00818f
C485 B.n252 VSUBS 0.00818f
C486 B.n253 VSUBS 0.00818f
C487 B.n254 VSUBS 0.00818f
C488 B.n255 VSUBS 0.00818f
C489 B.n256 VSUBS 0.00818f
C490 B.n257 VSUBS 0.00818f
C491 B.n258 VSUBS 0.00818f
C492 B.n259 VSUBS 0.00818f
C493 B.n260 VSUBS 0.00818f
C494 B.n261 VSUBS 0.00818f
C495 B.n262 VSUBS 0.00818f
C496 B.n263 VSUBS 0.00818f
C497 B.n264 VSUBS 0.00818f
C498 B.n265 VSUBS 0.00818f
C499 B.n266 VSUBS 0.00818f
C500 B.n267 VSUBS 0.00818f
C501 B.n268 VSUBS 0.019482f
C502 B.n269 VSUBS 0.018049f
C503 B.n270 VSUBS 0.018049f
C504 B.n271 VSUBS 0.00818f
C505 B.n272 VSUBS 0.00818f
C506 B.n273 VSUBS 0.00818f
C507 B.n274 VSUBS 0.00818f
C508 B.n275 VSUBS 0.00818f
C509 B.n276 VSUBS 0.00818f
C510 B.n277 VSUBS 0.00818f
C511 B.n278 VSUBS 0.00818f
C512 B.n279 VSUBS 0.00818f
C513 B.n280 VSUBS 0.00818f
C514 B.n281 VSUBS 0.00818f
C515 B.n282 VSUBS 0.00818f
C516 B.n283 VSUBS 0.00818f
C517 B.n284 VSUBS 0.00818f
C518 B.n285 VSUBS 0.00818f
C519 B.n286 VSUBS 0.00818f
C520 B.n287 VSUBS 0.00818f
C521 B.n288 VSUBS 0.00818f
C522 B.n289 VSUBS 0.00818f
C523 B.n290 VSUBS 0.00818f
C524 B.n291 VSUBS 0.018522f
.ends

