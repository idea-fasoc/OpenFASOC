* NGSPICE file created from diff_pair_sample_0028.ext - technology: sky130A

.subckt diff_pair_sample_0028 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t11 VP.t0 VDD1.t1 B.t5 sky130_fd_pr__nfet_01v8 ad=1.64505 pd=10.3 as=1.64505 ps=10.3 w=9.97 l=0.83
X1 VDD1.t0 VP.t1 VTAIL.t10 B.t0 sky130_fd_pr__nfet_01v8 ad=3.8883 pd=20.72 as=1.64505 ps=10.3 w=9.97 l=0.83
X2 VDD2.t5 VN.t0 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=1.64505 pd=10.3 as=3.8883 ps=20.72 w=9.97 l=0.83
X3 VDD1.t2 VP.t2 VTAIL.t9 B.t4 sky130_fd_pr__nfet_01v8 ad=1.64505 pd=10.3 as=3.8883 ps=20.72 w=9.97 l=0.83
X4 VDD2.t4 VN.t1 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=3.8883 pd=20.72 as=1.64505 ps=10.3 w=9.97 l=0.83
X5 VDD1.t4 VP.t3 VTAIL.t8 B.t2 sky130_fd_pr__nfet_01v8 ad=3.8883 pd=20.72 as=1.64505 ps=10.3 w=9.97 l=0.83
X6 B.t19 B.t17 B.t18 B.t14 sky130_fd_pr__nfet_01v8 ad=3.8883 pd=20.72 as=0 ps=0 w=9.97 l=0.83
X7 VTAIL.t7 VP.t4 VDD1.t5 B.t3 sky130_fd_pr__nfet_01v8 ad=1.64505 pd=10.3 as=1.64505 ps=10.3 w=9.97 l=0.83
X8 VTAIL.t3 VN.t2 VDD2.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=1.64505 pd=10.3 as=1.64505 ps=10.3 w=9.97 l=0.83
X9 B.t16 B.t13 B.t15 B.t14 sky130_fd_pr__nfet_01v8 ad=3.8883 pd=20.72 as=0 ps=0 w=9.97 l=0.83
X10 VDD2.t2 VN.t3 VTAIL.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=1.64505 pd=10.3 as=3.8883 ps=20.72 w=9.97 l=0.83
X11 B.t12 B.t10 B.t11 B.t7 sky130_fd_pr__nfet_01v8 ad=3.8883 pd=20.72 as=0 ps=0 w=9.97 l=0.83
X12 B.t9 B.t6 B.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=3.8883 pd=20.72 as=0 ps=0 w=9.97 l=0.83
X13 VTAIL.t5 VN.t4 VDD2.t1 B.t5 sky130_fd_pr__nfet_01v8 ad=1.64505 pd=10.3 as=1.64505 ps=10.3 w=9.97 l=0.83
X14 VDD2.t0 VN.t5 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=3.8883 pd=20.72 as=1.64505 ps=10.3 w=9.97 l=0.83
X15 VDD1.t3 VP.t5 VTAIL.t6 B.t1 sky130_fd_pr__nfet_01v8 ad=1.64505 pd=10.3 as=3.8883 ps=20.72 w=9.97 l=0.83
R0 VP.n3 VP.t1 352.361
R1 VP.n1 VP.t3 337.111
R2 VP.n13 VP.t2 337.111
R3 VP.n6 VP.t5 337.111
R4 VP.n11 VP.t4 289.49
R5 VP.n4 VP.t0 289.49
R6 VP.n5 VP.n2 161.3
R7 VP.n12 VP.n0 161.3
R8 VP.n10 VP.n9 161.3
R9 VP.n7 VP.n6 80.6037
R10 VP.n14 VP.n13 80.6037
R11 VP.n8 VP.n1 80.6037
R12 VP.n10 VP.n1 56.2746
R13 VP.n13 VP.n12 56.2746
R14 VP.n6 VP.n5 56.2746
R15 VP.n3 VP.n2 43.9052
R16 VP.n4 VP.n3 42.6472
R17 VP.n8 VP.n7 40.3044
R18 VP.n11 VP.n10 12.234
R19 VP.n12 VP.n11 12.234
R20 VP.n5 VP.n4 12.234
R21 VP.n7 VP.n2 0.285035
R22 VP.n9 VP.n8 0.285035
R23 VP.n14 VP.n0 0.285035
R24 VP.n9 VP.n0 0.189894
R25 VP VP.n14 0.146778
R26 VDD1.n48 VDD1.n0 289.615
R27 VDD1.n101 VDD1.n53 289.615
R28 VDD1.n49 VDD1.n48 185
R29 VDD1.n47 VDD1.n46 185
R30 VDD1.n4 VDD1.n3 185
R31 VDD1.n41 VDD1.n40 185
R32 VDD1.n39 VDD1.n6 185
R33 VDD1.n38 VDD1.n37 185
R34 VDD1.n9 VDD1.n7 185
R35 VDD1.n32 VDD1.n31 185
R36 VDD1.n30 VDD1.n29 185
R37 VDD1.n13 VDD1.n12 185
R38 VDD1.n24 VDD1.n23 185
R39 VDD1.n22 VDD1.n21 185
R40 VDD1.n17 VDD1.n16 185
R41 VDD1.n69 VDD1.n68 185
R42 VDD1.n74 VDD1.n73 185
R43 VDD1.n76 VDD1.n75 185
R44 VDD1.n65 VDD1.n64 185
R45 VDD1.n82 VDD1.n81 185
R46 VDD1.n84 VDD1.n83 185
R47 VDD1.n61 VDD1.n60 185
R48 VDD1.n91 VDD1.n90 185
R49 VDD1.n92 VDD1.n59 185
R50 VDD1.n94 VDD1.n93 185
R51 VDD1.n57 VDD1.n56 185
R52 VDD1.n100 VDD1.n99 185
R53 VDD1.n102 VDD1.n101 185
R54 VDD1.n18 VDD1.t0 149.524
R55 VDD1.n70 VDD1.t4 149.524
R56 VDD1.n48 VDD1.n47 104.615
R57 VDD1.n47 VDD1.n3 104.615
R58 VDD1.n40 VDD1.n3 104.615
R59 VDD1.n40 VDD1.n39 104.615
R60 VDD1.n39 VDD1.n38 104.615
R61 VDD1.n38 VDD1.n7 104.615
R62 VDD1.n31 VDD1.n7 104.615
R63 VDD1.n31 VDD1.n30 104.615
R64 VDD1.n30 VDD1.n12 104.615
R65 VDD1.n23 VDD1.n12 104.615
R66 VDD1.n23 VDD1.n22 104.615
R67 VDD1.n22 VDD1.n16 104.615
R68 VDD1.n74 VDD1.n68 104.615
R69 VDD1.n75 VDD1.n74 104.615
R70 VDD1.n75 VDD1.n64 104.615
R71 VDD1.n82 VDD1.n64 104.615
R72 VDD1.n83 VDD1.n82 104.615
R73 VDD1.n83 VDD1.n60 104.615
R74 VDD1.n91 VDD1.n60 104.615
R75 VDD1.n92 VDD1.n91 104.615
R76 VDD1.n93 VDD1.n92 104.615
R77 VDD1.n93 VDD1.n56 104.615
R78 VDD1.n100 VDD1.n56 104.615
R79 VDD1.n101 VDD1.n100 104.615
R80 VDD1.n107 VDD1.n106 63.0287
R81 VDD1.n109 VDD1.n108 62.8341
R82 VDD1.t0 VDD1.n16 52.3082
R83 VDD1.t4 VDD1.n68 52.3082
R84 VDD1 VDD1.n52 49.8663
R85 VDD1.n107 VDD1.n105 49.7527
R86 VDD1.n109 VDD1.n107 36.6431
R87 VDD1.n41 VDD1.n6 13.1884
R88 VDD1.n94 VDD1.n59 13.1884
R89 VDD1.n42 VDD1.n4 12.8005
R90 VDD1.n37 VDD1.n8 12.8005
R91 VDD1.n90 VDD1.n89 12.8005
R92 VDD1.n95 VDD1.n57 12.8005
R93 VDD1.n46 VDD1.n45 12.0247
R94 VDD1.n36 VDD1.n9 12.0247
R95 VDD1.n88 VDD1.n61 12.0247
R96 VDD1.n99 VDD1.n98 12.0247
R97 VDD1.n49 VDD1.n2 11.249
R98 VDD1.n33 VDD1.n32 11.249
R99 VDD1.n85 VDD1.n84 11.249
R100 VDD1.n102 VDD1.n55 11.249
R101 VDD1.n50 VDD1.n0 10.4732
R102 VDD1.n29 VDD1.n11 10.4732
R103 VDD1.n81 VDD1.n63 10.4732
R104 VDD1.n103 VDD1.n53 10.4732
R105 VDD1.n18 VDD1.n17 10.2747
R106 VDD1.n70 VDD1.n69 10.2747
R107 VDD1.n28 VDD1.n13 9.69747
R108 VDD1.n80 VDD1.n65 9.69747
R109 VDD1.n52 VDD1.n51 9.45567
R110 VDD1.n105 VDD1.n104 9.45567
R111 VDD1.n20 VDD1.n19 9.3005
R112 VDD1.n15 VDD1.n14 9.3005
R113 VDD1.n26 VDD1.n25 9.3005
R114 VDD1.n28 VDD1.n27 9.3005
R115 VDD1.n11 VDD1.n10 9.3005
R116 VDD1.n34 VDD1.n33 9.3005
R117 VDD1.n36 VDD1.n35 9.3005
R118 VDD1.n8 VDD1.n5 9.3005
R119 VDD1.n51 VDD1.n50 9.3005
R120 VDD1.n2 VDD1.n1 9.3005
R121 VDD1.n45 VDD1.n44 9.3005
R122 VDD1.n43 VDD1.n42 9.3005
R123 VDD1.n104 VDD1.n103 9.3005
R124 VDD1.n55 VDD1.n54 9.3005
R125 VDD1.n98 VDD1.n97 9.3005
R126 VDD1.n96 VDD1.n95 9.3005
R127 VDD1.n72 VDD1.n71 9.3005
R128 VDD1.n67 VDD1.n66 9.3005
R129 VDD1.n78 VDD1.n77 9.3005
R130 VDD1.n80 VDD1.n79 9.3005
R131 VDD1.n63 VDD1.n62 9.3005
R132 VDD1.n86 VDD1.n85 9.3005
R133 VDD1.n88 VDD1.n87 9.3005
R134 VDD1.n89 VDD1.n58 9.3005
R135 VDD1.n25 VDD1.n24 8.92171
R136 VDD1.n77 VDD1.n76 8.92171
R137 VDD1.n21 VDD1.n15 8.14595
R138 VDD1.n73 VDD1.n67 8.14595
R139 VDD1.n20 VDD1.n17 7.3702
R140 VDD1.n72 VDD1.n69 7.3702
R141 VDD1.n21 VDD1.n20 5.81868
R142 VDD1.n73 VDD1.n72 5.81868
R143 VDD1.n24 VDD1.n15 5.04292
R144 VDD1.n76 VDD1.n67 5.04292
R145 VDD1.n25 VDD1.n13 4.26717
R146 VDD1.n77 VDD1.n65 4.26717
R147 VDD1.n52 VDD1.n0 3.49141
R148 VDD1.n29 VDD1.n28 3.49141
R149 VDD1.n81 VDD1.n80 3.49141
R150 VDD1.n105 VDD1.n53 3.49141
R151 VDD1.n19 VDD1.n18 2.84303
R152 VDD1.n71 VDD1.n70 2.84303
R153 VDD1.n50 VDD1.n49 2.71565
R154 VDD1.n32 VDD1.n11 2.71565
R155 VDD1.n84 VDD1.n63 2.71565
R156 VDD1.n103 VDD1.n102 2.71565
R157 VDD1.n108 VDD1.t1 1.98646
R158 VDD1.n108 VDD1.t3 1.98646
R159 VDD1.n106 VDD1.t5 1.98646
R160 VDD1.n106 VDD1.t2 1.98646
R161 VDD1.n46 VDD1.n2 1.93989
R162 VDD1.n33 VDD1.n9 1.93989
R163 VDD1.n85 VDD1.n61 1.93989
R164 VDD1.n99 VDD1.n55 1.93989
R165 VDD1.n45 VDD1.n4 1.16414
R166 VDD1.n37 VDD1.n36 1.16414
R167 VDD1.n90 VDD1.n88 1.16414
R168 VDD1.n98 VDD1.n57 1.16414
R169 VDD1.n42 VDD1.n41 0.388379
R170 VDD1.n8 VDD1.n6 0.388379
R171 VDD1.n89 VDD1.n59 0.388379
R172 VDD1.n95 VDD1.n94 0.388379
R173 VDD1 VDD1.n109 0.19231
R174 VDD1.n51 VDD1.n1 0.155672
R175 VDD1.n44 VDD1.n1 0.155672
R176 VDD1.n44 VDD1.n43 0.155672
R177 VDD1.n43 VDD1.n5 0.155672
R178 VDD1.n35 VDD1.n5 0.155672
R179 VDD1.n35 VDD1.n34 0.155672
R180 VDD1.n34 VDD1.n10 0.155672
R181 VDD1.n27 VDD1.n10 0.155672
R182 VDD1.n27 VDD1.n26 0.155672
R183 VDD1.n26 VDD1.n14 0.155672
R184 VDD1.n19 VDD1.n14 0.155672
R185 VDD1.n71 VDD1.n66 0.155672
R186 VDD1.n78 VDD1.n66 0.155672
R187 VDD1.n79 VDD1.n78 0.155672
R188 VDD1.n79 VDD1.n62 0.155672
R189 VDD1.n86 VDD1.n62 0.155672
R190 VDD1.n87 VDD1.n86 0.155672
R191 VDD1.n87 VDD1.n58 0.155672
R192 VDD1.n96 VDD1.n58 0.155672
R193 VDD1.n97 VDD1.n96 0.155672
R194 VDD1.n97 VDD1.n54 0.155672
R195 VDD1.n104 VDD1.n54 0.155672
R196 VTAIL.n218 VTAIL.n170 289.615
R197 VTAIL.n50 VTAIL.n2 289.615
R198 VTAIL.n164 VTAIL.n116 289.615
R199 VTAIL.n108 VTAIL.n60 289.615
R200 VTAIL.n186 VTAIL.n185 185
R201 VTAIL.n191 VTAIL.n190 185
R202 VTAIL.n193 VTAIL.n192 185
R203 VTAIL.n182 VTAIL.n181 185
R204 VTAIL.n199 VTAIL.n198 185
R205 VTAIL.n201 VTAIL.n200 185
R206 VTAIL.n178 VTAIL.n177 185
R207 VTAIL.n208 VTAIL.n207 185
R208 VTAIL.n209 VTAIL.n176 185
R209 VTAIL.n211 VTAIL.n210 185
R210 VTAIL.n174 VTAIL.n173 185
R211 VTAIL.n217 VTAIL.n216 185
R212 VTAIL.n219 VTAIL.n218 185
R213 VTAIL.n18 VTAIL.n17 185
R214 VTAIL.n23 VTAIL.n22 185
R215 VTAIL.n25 VTAIL.n24 185
R216 VTAIL.n14 VTAIL.n13 185
R217 VTAIL.n31 VTAIL.n30 185
R218 VTAIL.n33 VTAIL.n32 185
R219 VTAIL.n10 VTAIL.n9 185
R220 VTAIL.n40 VTAIL.n39 185
R221 VTAIL.n41 VTAIL.n8 185
R222 VTAIL.n43 VTAIL.n42 185
R223 VTAIL.n6 VTAIL.n5 185
R224 VTAIL.n49 VTAIL.n48 185
R225 VTAIL.n51 VTAIL.n50 185
R226 VTAIL.n165 VTAIL.n164 185
R227 VTAIL.n163 VTAIL.n162 185
R228 VTAIL.n120 VTAIL.n119 185
R229 VTAIL.n157 VTAIL.n156 185
R230 VTAIL.n155 VTAIL.n122 185
R231 VTAIL.n154 VTAIL.n153 185
R232 VTAIL.n125 VTAIL.n123 185
R233 VTAIL.n148 VTAIL.n147 185
R234 VTAIL.n146 VTAIL.n145 185
R235 VTAIL.n129 VTAIL.n128 185
R236 VTAIL.n140 VTAIL.n139 185
R237 VTAIL.n138 VTAIL.n137 185
R238 VTAIL.n133 VTAIL.n132 185
R239 VTAIL.n109 VTAIL.n108 185
R240 VTAIL.n107 VTAIL.n106 185
R241 VTAIL.n64 VTAIL.n63 185
R242 VTAIL.n101 VTAIL.n100 185
R243 VTAIL.n99 VTAIL.n66 185
R244 VTAIL.n98 VTAIL.n97 185
R245 VTAIL.n69 VTAIL.n67 185
R246 VTAIL.n92 VTAIL.n91 185
R247 VTAIL.n90 VTAIL.n89 185
R248 VTAIL.n73 VTAIL.n72 185
R249 VTAIL.n84 VTAIL.n83 185
R250 VTAIL.n82 VTAIL.n81 185
R251 VTAIL.n77 VTAIL.n76 185
R252 VTAIL.n187 VTAIL.t1 149.524
R253 VTAIL.n19 VTAIL.t9 149.524
R254 VTAIL.n134 VTAIL.t6 149.524
R255 VTAIL.n78 VTAIL.t4 149.524
R256 VTAIL.n191 VTAIL.n185 104.615
R257 VTAIL.n192 VTAIL.n191 104.615
R258 VTAIL.n192 VTAIL.n181 104.615
R259 VTAIL.n199 VTAIL.n181 104.615
R260 VTAIL.n200 VTAIL.n199 104.615
R261 VTAIL.n200 VTAIL.n177 104.615
R262 VTAIL.n208 VTAIL.n177 104.615
R263 VTAIL.n209 VTAIL.n208 104.615
R264 VTAIL.n210 VTAIL.n209 104.615
R265 VTAIL.n210 VTAIL.n173 104.615
R266 VTAIL.n217 VTAIL.n173 104.615
R267 VTAIL.n218 VTAIL.n217 104.615
R268 VTAIL.n23 VTAIL.n17 104.615
R269 VTAIL.n24 VTAIL.n23 104.615
R270 VTAIL.n24 VTAIL.n13 104.615
R271 VTAIL.n31 VTAIL.n13 104.615
R272 VTAIL.n32 VTAIL.n31 104.615
R273 VTAIL.n32 VTAIL.n9 104.615
R274 VTAIL.n40 VTAIL.n9 104.615
R275 VTAIL.n41 VTAIL.n40 104.615
R276 VTAIL.n42 VTAIL.n41 104.615
R277 VTAIL.n42 VTAIL.n5 104.615
R278 VTAIL.n49 VTAIL.n5 104.615
R279 VTAIL.n50 VTAIL.n49 104.615
R280 VTAIL.n164 VTAIL.n163 104.615
R281 VTAIL.n163 VTAIL.n119 104.615
R282 VTAIL.n156 VTAIL.n119 104.615
R283 VTAIL.n156 VTAIL.n155 104.615
R284 VTAIL.n155 VTAIL.n154 104.615
R285 VTAIL.n154 VTAIL.n123 104.615
R286 VTAIL.n147 VTAIL.n123 104.615
R287 VTAIL.n147 VTAIL.n146 104.615
R288 VTAIL.n146 VTAIL.n128 104.615
R289 VTAIL.n139 VTAIL.n128 104.615
R290 VTAIL.n139 VTAIL.n138 104.615
R291 VTAIL.n138 VTAIL.n132 104.615
R292 VTAIL.n108 VTAIL.n107 104.615
R293 VTAIL.n107 VTAIL.n63 104.615
R294 VTAIL.n100 VTAIL.n63 104.615
R295 VTAIL.n100 VTAIL.n99 104.615
R296 VTAIL.n99 VTAIL.n98 104.615
R297 VTAIL.n98 VTAIL.n67 104.615
R298 VTAIL.n91 VTAIL.n67 104.615
R299 VTAIL.n91 VTAIL.n90 104.615
R300 VTAIL.n90 VTAIL.n72 104.615
R301 VTAIL.n83 VTAIL.n72 104.615
R302 VTAIL.n83 VTAIL.n82 104.615
R303 VTAIL.n82 VTAIL.n76 104.615
R304 VTAIL.t1 VTAIL.n185 52.3082
R305 VTAIL.t9 VTAIL.n17 52.3082
R306 VTAIL.t6 VTAIL.n132 52.3082
R307 VTAIL.t4 VTAIL.n76 52.3082
R308 VTAIL.n115 VTAIL.n114 46.1555
R309 VTAIL.n59 VTAIL.n58 46.1555
R310 VTAIL.n1 VTAIL.n0 46.1553
R311 VTAIL.n57 VTAIL.n56 46.1553
R312 VTAIL.n223 VTAIL.n222 32.3793
R313 VTAIL.n55 VTAIL.n54 32.3793
R314 VTAIL.n169 VTAIL.n168 32.3793
R315 VTAIL.n113 VTAIL.n112 32.3793
R316 VTAIL.n59 VTAIL.n57 22.9617
R317 VTAIL.n223 VTAIL.n169 21.9617
R318 VTAIL.n211 VTAIL.n176 13.1884
R319 VTAIL.n43 VTAIL.n8 13.1884
R320 VTAIL.n157 VTAIL.n122 13.1884
R321 VTAIL.n101 VTAIL.n66 13.1884
R322 VTAIL.n207 VTAIL.n206 12.8005
R323 VTAIL.n212 VTAIL.n174 12.8005
R324 VTAIL.n39 VTAIL.n38 12.8005
R325 VTAIL.n44 VTAIL.n6 12.8005
R326 VTAIL.n158 VTAIL.n120 12.8005
R327 VTAIL.n153 VTAIL.n124 12.8005
R328 VTAIL.n102 VTAIL.n64 12.8005
R329 VTAIL.n97 VTAIL.n68 12.8005
R330 VTAIL.n205 VTAIL.n178 12.0247
R331 VTAIL.n216 VTAIL.n215 12.0247
R332 VTAIL.n37 VTAIL.n10 12.0247
R333 VTAIL.n48 VTAIL.n47 12.0247
R334 VTAIL.n162 VTAIL.n161 12.0247
R335 VTAIL.n152 VTAIL.n125 12.0247
R336 VTAIL.n106 VTAIL.n105 12.0247
R337 VTAIL.n96 VTAIL.n69 12.0247
R338 VTAIL.n202 VTAIL.n201 11.249
R339 VTAIL.n219 VTAIL.n172 11.249
R340 VTAIL.n34 VTAIL.n33 11.249
R341 VTAIL.n51 VTAIL.n4 11.249
R342 VTAIL.n165 VTAIL.n118 11.249
R343 VTAIL.n149 VTAIL.n148 11.249
R344 VTAIL.n109 VTAIL.n62 11.249
R345 VTAIL.n93 VTAIL.n92 11.249
R346 VTAIL.n198 VTAIL.n180 10.4732
R347 VTAIL.n220 VTAIL.n170 10.4732
R348 VTAIL.n30 VTAIL.n12 10.4732
R349 VTAIL.n52 VTAIL.n2 10.4732
R350 VTAIL.n166 VTAIL.n116 10.4732
R351 VTAIL.n145 VTAIL.n127 10.4732
R352 VTAIL.n110 VTAIL.n60 10.4732
R353 VTAIL.n89 VTAIL.n71 10.4732
R354 VTAIL.n187 VTAIL.n186 10.2747
R355 VTAIL.n19 VTAIL.n18 10.2747
R356 VTAIL.n134 VTAIL.n133 10.2747
R357 VTAIL.n78 VTAIL.n77 10.2747
R358 VTAIL.n197 VTAIL.n182 9.69747
R359 VTAIL.n29 VTAIL.n14 9.69747
R360 VTAIL.n144 VTAIL.n129 9.69747
R361 VTAIL.n88 VTAIL.n73 9.69747
R362 VTAIL.n222 VTAIL.n221 9.45567
R363 VTAIL.n54 VTAIL.n53 9.45567
R364 VTAIL.n168 VTAIL.n167 9.45567
R365 VTAIL.n112 VTAIL.n111 9.45567
R366 VTAIL.n221 VTAIL.n220 9.3005
R367 VTAIL.n172 VTAIL.n171 9.3005
R368 VTAIL.n215 VTAIL.n214 9.3005
R369 VTAIL.n213 VTAIL.n212 9.3005
R370 VTAIL.n189 VTAIL.n188 9.3005
R371 VTAIL.n184 VTAIL.n183 9.3005
R372 VTAIL.n195 VTAIL.n194 9.3005
R373 VTAIL.n197 VTAIL.n196 9.3005
R374 VTAIL.n180 VTAIL.n179 9.3005
R375 VTAIL.n203 VTAIL.n202 9.3005
R376 VTAIL.n205 VTAIL.n204 9.3005
R377 VTAIL.n206 VTAIL.n175 9.3005
R378 VTAIL.n53 VTAIL.n52 9.3005
R379 VTAIL.n4 VTAIL.n3 9.3005
R380 VTAIL.n47 VTAIL.n46 9.3005
R381 VTAIL.n45 VTAIL.n44 9.3005
R382 VTAIL.n21 VTAIL.n20 9.3005
R383 VTAIL.n16 VTAIL.n15 9.3005
R384 VTAIL.n27 VTAIL.n26 9.3005
R385 VTAIL.n29 VTAIL.n28 9.3005
R386 VTAIL.n12 VTAIL.n11 9.3005
R387 VTAIL.n35 VTAIL.n34 9.3005
R388 VTAIL.n37 VTAIL.n36 9.3005
R389 VTAIL.n38 VTAIL.n7 9.3005
R390 VTAIL.n136 VTAIL.n135 9.3005
R391 VTAIL.n131 VTAIL.n130 9.3005
R392 VTAIL.n142 VTAIL.n141 9.3005
R393 VTAIL.n144 VTAIL.n143 9.3005
R394 VTAIL.n127 VTAIL.n126 9.3005
R395 VTAIL.n150 VTAIL.n149 9.3005
R396 VTAIL.n152 VTAIL.n151 9.3005
R397 VTAIL.n124 VTAIL.n121 9.3005
R398 VTAIL.n167 VTAIL.n166 9.3005
R399 VTAIL.n118 VTAIL.n117 9.3005
R400 VTAIL.n161 VTAIL.n160 9.3005
R401 VTAIL.n159 VTAIL.n158 9.3005
R402 VTAIL.n80 VTAIL.n79 9.3005
R403 VTAIL.n75 VTAIL.n74 9.3005
R404 VTAIL.n86 VTAIL.n85 9.3005
R405 VTAIL.n88 VTAIL.n87 9.3005
R406 VTAIL.n71 VTAIL.n70 9.3005
R407 VTAIL.n94 VTAIL.n93 9.3005
R408 VTAIL.n96 VTAIL.n95 9.3005
R409 VTAIL.n68 VTAIL.n65 9.3005
R410 VTAIL.n111 VTAIL.n110 9.3005
R411 VTAIL.n62 VTAIL.n61 9.3005
R412 VTAIL.n105 VTAIL.n104 9.3005
R413 VTAIL.n103 VTAIL.n102 9.3005
R414 VTAIL.n194 VTAIL.n193 8.92171
R415 VTAIL.n26 VTAIL.n25 8.92171
R416 VTAIL.n141 VTAIL.n140 8.92171
R417 VTAIL.n85 VTAIL.n84 8.92171
R418 VTAIL.n190 VTAIL.n184 8.14595
R419 VTAIL.n22 VTAIL.n16 8.14595
R420 VTAIL.n137 VTAIL.n131 8.14595
R421 VTAIL.n81 VTAIL.n75 8.14595
R422 VTAIL.n189 VTAIL.n186 7.3702
R423 VTAIL.n21 VTAIL.n18 7.3702
R424 VTAIL.n136 VTAIL.n133 7.3702
R425 VTAIL.n80 VTAIL.n77 7.3702
R426 VTAIL.n190 VTAIL.n189 5.81868
R427 VTAIL.n22 VTAIL.n21 5.81868
R428 VTAIL.n137 VTAIL.n136 5.81868
R429 VTAIL.n81 VTAIL.n80 5.81868
R430 VTAIL.n193 VTAIL.n184 5.04292
R431 VTAIL.n25 VTAIL.n16 5.04292
R432 VTAIL.n140 VTAIL.n131 5.04292
R433 VTAIL.n84 VTAIL.n75 5.04292
R434 VTAIL.n194 VTAIL.n182 4.26717
R435 VTAIL.n26 VTAIL.n14 4.26717
R436 VTAIL.n141 VTAIL.n129 4.26717
R437 VTAIL.n85 VTAIL.n73 4.26717
R438 VTAIL.n198 VTAIL.n197 3.49141
R439 VTAIL.n222 VTAIL.n170 3.49141
R440 VTAIL.n30 VTAIL.n29 3.49141
R441 VTAIL.n54 VTAIL.n2 3.49141
R442 VTAIL.n168 VTAIL.n116 3.49141
R443 VTAIL.n145 VTAIL.n144 3.49141
R444 VTAIL.n112 VTAIL.n60 3.49141
R445 VTAIL.n89 VTAIL.n88 3.49141
R446 VTAIL.n188 VTAIL.n187 2.84303
R447 VTAIL.n20 VTAIL.n19 2.84303
R448 VTAIL.n135 VTAIL.n134 2.84303
R449 VTAIL.n79 VTAIL.n78 2.84303
R450 VTAIL.n201 VTAIL.n180 2.71565
R451 VTAIL.n220 VTAIL.n219 2.71565
R452 VTAIL.n33 VTAIL.n12 2.71565
R453 VTAIL.n52 VTAIL.n51 2.71565
R454 VTAIL.n166 VTAIL.n165 2.71565
R455 VTAIL.n148 VTAIL.n127 2.71565
R456 VTAIL.n110 VTAIL.n109 2.71565
R457 VTAIL.n92 VTAIL.n71 2.71565
R458 VTAIL.n0 VTAIL.t0 1.98646
R459 VTAIL.n0 VTAIL.t5 1.98646
R460 VTAIL.n56 VTAIL.t8 1.98646
R461 VTAIL.n56 VTAIL.t7 1.98646
R462 VTAIL.n114 VTAIL.t10 1.98646
R463 VTAIL.n114 VTAIL.t11 1.98646
R464 VTAIL.n58 VTAIL.t2 1.98646
R465 VTAIL.n58 VTAIL.t3 1.98646
R466 VTAIL.n202 VTAIL.n178 1.93989
R467 VTAIL.n216 VTAIL.n172 1.93989
R468 VTAIL.n34 VTAIL.n10 1.93989
R469 VTAIL.n48 VTAIL.n4 1.93989
R470 VTAIL.n162 VTAIL.n118 1.93989
R471 VTAIL.n149 VTAIL.n125 1.93989
R472 VTAIL.n106 VTAIL.n62 1.93989
R473 VTAIL.n93 VTAIL.n69 1.93989
R474 VTAIL.n207 VTAIL.n205 1.16414
R475 VTAIL.n215 VTAIL.n174 1.16414
R476 VTAIL.n39 VTAIL.n37 1.16414
R477 VTAIL.n47 VTAIL.n6 1.16414
R478 VTAIL.n161 VTAIL.n120 1.16414
R479 VTAIL.n153 VTAIL.n152 1.16414
R480 VTAIL.n105 VTAIL.n64 1.16414
R481 VTAIL.n97 VTAIL.n96 1.16414
R482 VTAIL.n113 VTAIL.n59 1.0005
R483 VTAIL.n169 VTAIL.n115 1.0005
R484 VTAIL.n57 VTAIL.n55 1.0005
R485 VTAIL.n115 VTAIL.n113 0.970328
R486 VTAIL.n55 VTAIL.n1 0.970328
R487 VTAIL VTAIL.n223 0.69231
R488 VTAIL.n206 VTAIL.n176 0.388379
R489 VTAIL.n212 VTAIL.n211 0.388379
R490 VTAIL.n38 VTAIL.n8 0.388379
R491 VTAIL.n44 VTAIL.n43 0.388379
R492 VTAIL.n158 VTAIL.n157 0.388379
R493 VTAIL.n124 VTAIL.n122 0.388379
R494 VTAIL.n102 VTAIL.n101 0.388379
R495 VTAIL.n68 VTAIL.n66 0.388379
R496 VTAIL VTAIL.n1 0.30869
R497 VTAIL.n188 VTAIL.n183 0.155672
R498 VTAIL.n195 VTAIL.n183 0.155672
R499 VTAIL.n196 VTAIL.n195 0.155672
R500 VTAIL.n196 VTAIL.n179 0.155672
R501 VTAIL.n203 VTAIL.n179 0.155672
R502 VTAIL.n204 VTAIL.n203 0.155672
R503 VTAIL.n204 VTAIL.n175 0.155672
R504 VTAIL.n213 VTAIL.n175 0.155672
R505 VTAIL.n214 VTAIL.n213 0.155672
R506 VTAIL.n214 VTAIL.n171 0.155672
R507 VTAIL.n221 VTAIL.n171 0.155672
R508 VTAIL.n20 VTAIL.n15 0.155672
R509 VTAIL.n27 VTAIL.n15 0.155672
R510 VTAIL.n28 VTAIL.n27 0.155672
R511 VTAIL.n28 VTAIL.n11 0.155672
R512 VTAIL.n35 VTAIL.n11 0.155672
R513 VTAIL.n36 VTAIL.n35 0.155672
R514 VTAIL.n36 VTAIL.n7 0.155672
R515 VTAIL.n45 VTAIL.n7 0.155672
R516 VTAIL.n46 VTAIL.n45 0.155672
R517 VTAIL.n46 VTAIL.n3 0.155672
R518 VTAIL.n53 VTAIL.n3 0.155672
R519 VTAIL.n167 VTAIL.n117 0.155672
R520 VTAIL.n160 VTAIL.n117 0.155672
R521 VTAIL.n160 VTAIL.n159 0.155672
R522 VTAIL.n159 VTAIL.n121 0.155672
R523 VTAIL.n151 VTAIL.n121 0.155672
R524 VTAIL.n151 VTAIL.n150 0.155672
R525 VTAIL.n150 VTAIL.n126 0.155672
R526 VTAIL.n143 VTAIL.n126 0.155672
R527 VTAIL.n143 VTAIL.n142 0.155672
R528 VTAIL.n142 VTAIL.n130 0.155672
R529 VTAIL.n135 VTAIL.n130 0.155672
R530 VTAIL.n111 VTAIL.n61 0.155672
R531 VTAIL.n104 VTAIL.n61 0.155672
R532 VTAIL.n104 VTAIL.n103 0.155672
R533 VTAIL.n103 VTAIL.n65 0.155672
R534 VTAIL.n95 VTAIL.n65 0.155672
R535 VTAIL.n95 VTAIL.n94 0.155672
R536 VTAIL.n94 VTAIL.n70 0.155672
R537 VTAIL.n87 VTAIL.n70 0.155672
R538 VTAIL.n87 VTAIL.n86 0.155672
R539 VTAIL.n86 VTAIL.n74 0.155672
R540 VTAIL.n79 VTAIL.n74 0.155672
R541 B.n590 B.n589 585
R542 B.n591 B.n590 585
R543 B.n248 B.n83 585
R544 B.n247 B.n246 585
R545 B.n245 B.n244 585
R546 B.n243 B.n242 585
R547 B.n241 B.n240 585
R548 B.n239 B.n238 585
R549 B.n237 B.n236 585
R550 B.n235 B.n234 585
R551 B.n233 B.n232 585
R552 B.n231 B.n230 585
R553 B.n229 B.n228 585
R554 B.n227 B.n226 585
R555 B.n225 B.n224 585
R556 B.n223 B.n222 585
R557 B.n221 B.n220 585
R558 B.n219 B.n218 585
R559 B.n217 B.n216 585
R560 B.n215 B.n214 585
R561 B.n213 B.n212 585
R562 B.n211 B.n210 585
R563 B.n209 B.n208 585
R564 B.n207 B.n206 585
R565 B.n205 B.n204 585
R566 B.n203 B.n202 585
R567 B.n201 B.n200 585
R568 B.n199 B.n198 585
R569 B.n197 B.n196 585
R570 B.n195 B.n194 585
R571 B.n193 B.n192 585
R572 B.n191 B.n190 585
R573 B.n189 B.n188 585
R574 B.n187 B.n186 585
R575 B.n185 B.n184 585
R576 B.n183 B.n182 585
R577 B.n181 B.n180 585
R578 B.n178 B.n177 585
R579 B.n176 B.n175 585
R580 B.n174 B.n173 585
R581 B.n172 B.n171 585
R582 B.n170 B.n169 585
R583 B.n168 B.n167 585
R584 B.n166 B.n165 585
R585 B.n164 B.n163 585
R586 B.n162 B.n161 585
R587 B.n160 B.n159 585
R588 B.n158 B.n157 585
R589 B.n156 B.n155 585
R590 B.n154 B.n153 585
R591 B.n152 B.n151 585
R592 B.n150 B.n149 585
R593 B.n148 B.n147 585
R594 B.n146 B.n145 585
R595 B.n144 B.n143 585
R596 B.n142 B.n141 585
R597 B.n140 B.n139 585
R598 B.n138 B.n137 585
R599 B.n136 B.n135 585
R600 B.n134 B.n133 585
R601 B.n132 B.n131 585
R602 B.n130 B.n129 585
R603 B.n128 B.n127 585
R604 B.n126 B.n125 585
R605 B.n124 B.n123 585
R606 B.n122 B.n121 585
R607 B.n120 B.n119 585
R608 B.n118 B.n117 585
R609 B.n116 B.n115 585
R610 B.n114 B.n113 585
R611 B.n112 B.n111 585
R612 B.n110 B.n109 585
R613 B.n108 B.n107 585
R614 B.n106 B.n105 585
R615 B.n104 B.n103 585
R616 B.n102 B.n101 585
R617 B.n100 B.n99 585
R618 B.n98 B.n97 585
R619 B.n96 B.n95 585
R620 B.n94 B.n93 585
R621 B.n92 B.n91 585
R622 B.n90 B.n89 585
R623 B.n588 B.n42 585
R624 B.n592 B.n42 585
R625 B.n587 B.n41 585
R626 B.n593 B.n41 585
R627 B.n586 B.n585 585
R628 B.n585 B.n37 585
R629 B.n584 B.n36 585
R630 B.n599 B.n36 585
R631 B.n583 B.n35 585
R632 B.n600 B.n35 585
R633 B.n582 B.n34 585
R634 B.n601 B.n34 585
R635 B.n581 B.n580 585
R636 B.n580 B.n30 585
R637 B.n579 B.n29 585
R638 B.n607 B.n29 585
R639 B.n578 B.n28 585
R640 B.n608 B.n28 585
R641 B.n577 B.n27 585
R642 B.n609 B.n27 585
R643 B.n576 B.n575 585
R644 B.n575 B.n23 585
R645 B.n574 B.n22 585
R646 B.n615 B.n22 585
R647 B.n573 B.n21 585
R648 B.n616 B.n21 585
R649 B.n572 B.n20 585
R650 B.n617 B.n20 585
R651 B.n571 B.n570 585
R652 B.n570 B.n19 585
R653 B.n569 B.n15 585
R654 B.n623 B.n15 585
R655 B.n568 B.n14 585
R656 B.n624 B.n14 585
R657 B.n567 B.n13 585
R658 B.n625 B.n13 585
R659 B.n566 B.n565 585
R660 B.n565 B.n12 585
R661 B.n564 B.n563 585
R662 B.n564 B.n8 585
R663 B.n562 B.n7 585
R664 B.n632 B.n7 585
R665 B.n561 B.n6 585
R666 B.n633 B.n6 585
R667 B.n560 B.n5 585
R668 B.n634 B.n5 585
R669 B.n559 B.n558 585
R670 B.n558 B.n4 585
R671 B.n557 B.n249 585
R672 B.n557 B.n556 585
R673 B.n546 B.n250 585
R674 B.n549 B.n250 585
R675 B.n548 B.n547 585
R676 B.n550 B.n548 585
R677 B.n545 B.n255 585
R678 B.n255 B.n254 585
R679 B.n544 B.n543 585
R680 B.n543 B.n542 585
R681 B.n257 B.n256 585
R682 B.n535 B.n257 585
R683 B.n534 B.n533 585
R684 B.n536 B.n534 585
R685 B.n532 B.n262 585
R686 B.n262 B.n261 585
R687 B.n531 B.n530 585
R688 B.n530 B.n529 585
R689 B.n264 B.n263 585
R690 B.n265 B.n264 585
R691 B.n522 B.n521 585
R692 B.n523 B.n522 585
R693 B.n520 B.n270 585
R694 B.n270 B.n269 585
R695 B.n519 B.n518 585
R696 B.n518 B.n517 585
R697 B.n272 B.n271 585
R698 B.n273 B.n272 585
R699 B.n510 B.n509 585
R700 B.n511 B.n510 585
R701 B.n508 B.n277 585
R702 B.n281 B.n277 585
R703 B.n507 B.n506 585
R704 B.n506 B.n505 585
R705 B.n279 B.n278 585
R706 B.n280 B.n279 585
R707 B.n498 B.n497 585
R708 B.n499 B.n498 585
R709 B.n496 B.n286 585
R710 B.n286 B.n285 585
R711 B.n490 B.n489 585
R712 B.n488 B.n328 585
R713 B.n487 B.n327 585
R714 B.n492 B.n327 585
R715 B.n486 B.n485 585
R716 B.n484 B.n483 585
R717 B.n482 B.n481 585
R718 B.n480 B.n479 585
R719 B.n478 B.n477 585
R720 B.n476 B.n475 585
R721 B.n474 B.n473 585
R722 B.n472 B.n471 585
R723 B.n470 B.n469 585
R724 B.n468 B.n467 585
R725 B.n466 B.n465 585
R726 B.n464 B.n463 585
R727 B.n462 B.n461 585
R728 B.n460 B.n459 585
R729 B.n458 B.n457 585
R730 B.n456 B.n455 585
R731 B.n454 B.n453 585
R732 B.n452 B.n451 585
R733 B.n450 B.n449 585
R734 B.n448 B.n447 585
R735 B.n446 B.n445 585
R736 B.n444 B.n443 585
R737 B.n442 B.n441 585
R738 B.n440 B.n439 585
R739 B.n438 B.n437 585
R740 B.n436 B.n435 585
R741 B.n434 B.n433 585
R742 B.n432 B.n431 585
R743 B.n430 B.n429 585
R744 B.n428 B.n427 585
R745 B.n426 B.n425 585
R746 B.n424 B.n423 585
R747 B.n422 B.n421 585
R748 B.n419 B.n418 585
R749 B.n417 B.n416 585
R750 B.n415 B.n414 585
R751 B.n413 B.n412 585
R752 B.n411 B.n410 585
R753 B.n409 B.n408 585
R754 B.n407 B.n406 585
R755 B.n405 B.n404 585
R756 B.n403 B.n402 585
R757 B.n401 B.n400 585
R758 B.n399 B.n398 585
R759 B.n397 B.n396 585
R760 B.n395 B.n394 585
R761 B.n393 B.n392 585
R762 B.n391 B.n390 585
R763 B.n389 B.n388 585
R764 B.n387 B.n386 585
R765 B.n385 B.n384 585
R766 B.n383 B.n382 585
R767 B.n381 B.n380 585
R768 B.n379 B.n378 585
R769 B.n377 B.n376 585
R770 B.n375 B.n374 585
R771 B.n373 B.n372 585
R772 B.n371 B.n370 585
R773 B.n369 B.n368 585
R774 B.n367 B.n366 585
R775 B.n365 B.n364 585
R776 B.n363 B.n362 585
R777 B.n361 B.n360 585
R778 B.n359 B.n358 585
R779 B.n357 B.n356 585
R780 B.n355 B.n354 585
R781 B.n353 B.n352 585
R782 B.n351 B.n350 585
R783 B.n349 B.n348 585
R784 B.n347 B.n346 585
R785 B.n345 B.n344 585
R786 B.n343 B.n342 585
R787 B.n341 B.n340 585
R788 B.n339 B.n338 585
R789 B.n337 B.n336 585
R790 B.n335 B.n334 585
R791 B.n288 B.n287 585
R792 B.n495 B.n494 585
R793 B.n284 B.n283 585
R794 B.n285 B.n284 585
R795 B.n501 B.n500 585
R796 B.n500 B.n499 585
R797 B.n502 B.n282 585
R798 B.n282 B.n280 585
R799 B.n504 B.n503 585
R800 B.n505 B.n504 585
R801 B.n276 B.n275 585
R802 B.n281 B.n276 585
R803 B.n513 B.n512 585
R804 B.n512 B.n511 585
R805 B.n514 B.n274 585
R806 B.n274 B.n273 585
R807 B.n516 B.n515 585
R808 B.n517 B.n516 585
R809 B.n268 B.n267 585
R810 B.n269 B.n268 585
R811 B.n525 B.n524 585
R812 B.n524 B.n523 585
R813 B.n526 B.n266 585
R814 B.n266 B.n265 585
R815 B.n528 B.n527 585
R816 B.n529 B.n528 585
R817 B.n260 B.n259 585
R818 B.n261 B.n260 585
R819 B.n538 B.n537 585
R820 B.n537 B.n536 585
R821 B.n539 B.n258 585
R822 B.n535 B.n258 585
R823 B.n541 B.n540 585
R824 B.n542 B.n541 585
R825 B.n253 B.n252 585
R826 B.n254 B.n253 585
R827 B.n552 B.n551 585
R828 B.n551 B.n550 585
R829 B.n553 B.n251 585
R830 B.n549 B.n251 585
R831 B.n555 B.n554 585
R832 B.n556 B.n555 585
R833 B.n3 B.n0 585
R834 B.n4 B.n3 585
R835 B.n631 B.n1 585
R836 B.n632 B.n631 585
R837 B.n630 B.n629 585
R838 B.n630 B.n8 585
R839 B.n628 B.n9 585
R840 B.n12 B.n9 585
R841 B.n627 B.n626 585
R842 B.n626 B.n625 585
R843 B.n11 B.n10 585
R844 B.n624 B.n11 585
R845 B.n622 B.n621 585
R846 B.n623 B.n622 585
R847 B.n620 B.n16 585
R848 B.n19 B.n16 585
R849 B.n619 B.n618 585
R850 B.n618 B.n617 585
R851 B.n18 B.n17 585
R852 B.n616 B.n18 585
R853 B.n614 B.n613 585
R854 B.n615 B.n614 585
R855 B.n612 B.n24 585
R856 B.n24 B.n23 585
R857 B.n611 B.n610 585
R858 B.n610 B.n609 585
R859 B.n26 B.n25 585
R860 B.n608 B.n26 585
R861 B.n606 B.n605 585
R862 B.n607 B.n606 585
R863 B.n604 B.n31 585
R864 B.n31 B.n30 585
R865 B.n603 B.n602 585
R866 B.n602 B.n601 585
R867 B.n33 B.n32 585
R868 B.n600 B.n33 585
R869 B.n598 B.n597 585
R870 B.n599 B.n598 585
R871 B.n596 B.n38 585
R872 B.n38 B.n37 585
R873 B.n595 B.n594 585
R874 B.n594 B.n593 585
R875 B.n40 B.n39 585
R876 B.n592 B.n40 585
R877 B.n635 B.n634 585
R878 B.n633 B.n2 585
R879 B.n89 B.n40 530.939
R880 B.n590 B.n42 530.939
R881 B.n494 B.n286 530.939
R882 B.n490 B.n284 530.939
R883 B.n86 B.t10 491.108
R884 B.n84 B.t6 491.108
R885 B.n331 B.t13 491.108
R886 B.n329 B.t17 491.108
R887 B.n84 B.t8 269.562
R888 B.n331 B.t16 269.562
R889 B.n86 B.t11 269.562
R890 B.n329 B.t19 269.562
R891 B.n591 B.n82 256.663
R892 B.n591 B.n81 256.663
R893 B.n591 B.n80 256.663
R894 B.n591 B.n79 256.663
R895 B.n591 B.n78 256.663
R896 B.n591 B.n77 256.663
R897 B.n591 B.n76 256.663
R898 B.n591 B.n75 256.663
R899 B.n591 B.n74 256.663
R900 B.n591 B.n73 256.663
R901 B.n591 B.n72 256.663
R902 B.n591 B.n71 256.663
R903 B.n591 B.n70 256.663
R904 B.n591 B.n69 256.663
R905 B.n591 B.n68 256.663
R906 B.n591 B.n67 256.663
R907 B.n591 B.n66 256.663
R908 B.n591 B.n65 256.663
R909 B.n591 B.n64 256.663
R910 B.n591 B.n63 256.663
R911 B.n591 B.n62 256.663
R912 B.n591 B.n61 256.663
R913 B.n591 B.n60 256.663
R914 B.n591 B.n59 256.663
R915 B.n591 B.n58 256.663
R916 B.n591 B.n57 256.663
R917 B.n591 B.n56 256.663
R918 B.n591 B.n55 256.663
R919 B.n591 B.n54 256.663
R920 B.n591 B.n53 256.663
R921 B.n591 B.n52 256.663
R922 B.n591 B.n51 256.663
R923 B.n591 B.n50 256.663
R924 B.n591 B.n49 256.663
R925 B.n591 B.n48 256.663
R926 B.n591 B.n47 256.663
R927 B.n591 B.n46 256.663
R928 B.n591 B.n45 256.663
R929 B.n591 B.n44 256.663
R930 B.n591 B.n43 256.663
R931 B.n492 B.n491 256.663
R932 B.n492 B.n289 256.663
R933 B.n492 B.n290 256.663
R934 B.n492 B.n291 256.663
R935 B.n492 B.n292 256.663
R936 B.n492 B.n293 256.663
R937 B.n492 B.n294 256.663
R938 B.n492 B.n295 256.663
R939 B.n492 B.n296 256.663
R940 B.n492 B.n297 256.663
R941 B.n492 B.n298 256.663
R942 B.n492 B.n299 256.663
R943 B.n492 B.n300 256.663
R944 B.n492 B.n301 256.663
R945 B.n492 B.n302 256.663
R946 B.n492 B.n303 256.663
R947 B.n492 B.n304 256.663
R948 B.n492 B.n305 256.663
R949 B.n492 B.n306 256.663
R950 B.n492 B.n307 256.663
R951 B.n492 B.n308 256.663
R952 B.n492 B.n309 256.663
R953 B.n492 B.n310 256.663
R954 B.n492 B.n311 256.663
R955 B.n492 B.n312 256.663
R956 B.n492 B.n313 256.663
R957 B.n492 B.n314 256.663
R958 B.n492 B.n315 256.663
R959 B.n492 B.n316 256.663
R960 B.n492 B.n317 256.663
R961 B.n492 B.n318 256.663
R962 B.n492 B.n319 256.663
R963 B.n492 B.n320 256.663
R964 B.n492 B.n321 256.663
R965 B.n492 B.n322 256.663
R966 B.n492 B.n323 256.663
R967 B.n492 B.n324 256.663
R968 B.n492 B.n325 256.663
R969 B.n492 B.n326 256.663
R970 B.n493 B.n492 256.663
R971 B.n637 B.n636 256.663
R972 B.n85 B.t9 247.065
R973 B.n332 B.t15 247.065
R974 B.n87 B.t12 247.065
R975 B.n330 B.t18 247.065
R976 B.n93 B.n92 163.367
R977 B.n97 B.n96 163.367
R978 B.n101 B.n100 163.367
R979 B.n105 B.n104 163.367
R980 B.n109 B.n108 163.367
R981 B.n113 B.n112 163.367
R982 B.n117 B.n116 163.367
R983 B.n121 B.n120 163.367
R984 B.n125 B.n124 163.367
R985 B.n129 B.n128 163.367
R986 B.n133 B.n132 163.367
R987 B.n137 B.n136 163.367
R988 B.n141 B.n140 163.367
R989 B.n145 B.n144 163.367
R990 B.n149 B.n148 163.367
R991 B.n153 B.n152 163.367
R992 B.n157 B.n156 163.367
R993 B.n161 B.n160 163.367
R994 B.n165 B.n164 163.367
R995 B.n169 B.n168 163.367
R996 B.n173 B.n172 163.367
R997 B.n177 B.n176 163.367
R998 B.n182 B.n181 163.367
R999 B.n186 B.n185 163.367
R1000 B.n190 B.n189 163.367
R1001 B.n194 B.n193 163.367
R1002 B.n198 B.n197 163.367
R1003 B.n202 B.n201 163.367
R1004 B.n206 B.n205 163.367
R1005 B.n210 B.n209 163.367
R1006 B.n214 B.n213 163.367
R1007 B.n218 B.n217 163.367
R1008 B.n222 B.n221 163.367
R1009 B.n226 B.n225 163.367
R1010 B.n230 B.n229 163.367
R1011 B.n234 B.n233 163.367
R1012 B.n238 B.n237 163.367
R1013 B.n242 B.n241 163.367
R1014 B.n246 B.n245 163.367
R1015 B.n590 B.n83 163.367
R1016 B.n498 B.n286 163.367
R1017 B.n498 B.n279 163.367
R1018 B.n506 B.n279 163.367
R1019 B.n506 B.n277 163.367
R1020 B.n510 B.n277 163.367
R1021 B.n510 B.n272 163.367
R1022 B.n518 B.n272 163.367
R1023 B.n518 B.n270 163.367
R1024 B.n522 B.n270 163.367
R1025 B.n522 B.n264 163.367
R1026 B.n530 B.n264 163.367
R1027 B.n530 B.n262 163.367
R1028 B.n534 B.n262 163.367
R1029 B.n534 B.n257 163.367
R1030 B.n543 B.n257 163.367
R1031 B.n543 B.n255 163.367
R1032 B.n548 B.n255 163.367
R1033 B.n548 B.n250 163.367
R1034 B.n557 B.n250 163.367
R1035 B.n558 B.n557 163.367
R1036 B.n558 B.n5 163.367
R1037 B.n6 B.n5 163.367
R1038 B.n7 B.n6 163.367
R1039 B.n564 B.n7 163.367
R1040 B.n565 B.n564 163.367
R1041 B.n565 B.n13 163.367
R1042 B.n14 B.n13 163.367
R1043 B.n15 B.n14 163.367
R1044 B.n570 B.n15 163.367
R1045 B.n570 B.n20 163.367
R1046 B.n21 B.n20 163.367
R1047 B.n22 B.n21 163.367
R1048 B.n575 B.n22 163.367
R1049 B.n575 B.n27 163.367
R1050 B.n28 B.n27 163.367
R1051 B.n29 B.n28 163.367
R1052 B.n580 B.n29 163.367
R1053 B.n580 B.n34 163.367
R1054 B.n35 B.n34 163.367
R1055 B.n36 B.n35 163.367
R1056 B.n585 B.n36 163.367
R1057 B.n585 B.n41 163.367
R1058 B.n42 B.n41 163.367
R1059 B.n328 B.n327 163.367
R1060 B.n485 B.n327 163.367
R1061 B.n483 B.n482 163.367
R1062 B.n479 B.n478 163.367
R1063 B.n475 B.n474 163.367
R1064 B.n471 B.n470 163.367
R1065 B.n467 B.n466 163.367
R1066 B.n463 B.n462 163.367
R1067 B.n459 B.n458 163.367
R1068 B.n455 B.n454 163.367
R1069 B.n451 B.n450 163.367
R1070 B.n447 B.n446 163.367
R1071 B.n443 B.n442 163.367
R1072 B.n439 B.n438 163.367
R1073 B.n435 B.n434 163.367
R1074 B.n431 B.n430 163.367
R1075 B.n427 B.n426 163.367
R1076 B.n423 B.n422 163.367
R1077 B.n418 B.n417 163.367
R1078 B.n414 B.n413 163.367
R1079 B.n410 B.n409 163.367
R1080 B.n406 B.n405 163.367
R1081 B.n402 B.n401 163.367
R1082 B.n398 B.n397 163.367
R1083 B.n394 B.n393 163.367
R1084 B.n390 B.n389 163.367
R1085 B.n386 B.n385 163.367
R1086 B.n382 B.n381 163.367
R1087 B.n378 B.n377 163.367
R1088 B.n374 B.n373 163.367
R1089 B.n370 B.n369 163.367
R1090 B.n366 B.n365 163.367
R1091 B.n362 B.n361 163.367
R1092 B.n358 B.n357 163.367
R1093 B.n354 B.n353 163.367
R1094 B.n350 B.n349 163.367
R1095 B.n346 B.n345 163.367
R1096 B.n342 B.n341 163.367
R1097 B.n338 B.n337 163.367
R1098 B.n334 B.n288 163.367
R1099 B.n500 B.n284 163.367
R1100 B.n500 B.n282 163.367
R1101 B.n504 B.n282 163.367
R1102 B.n504 B.n276 163.367
R1103 B.n512 B.n276 163.367
R1104 B.n512 B.n274 163.367
R1105 B.n516 B.n274 163.367
R1106 B.n516 B.n268 163.367
R1107 B.n524 B.n268 163.367
R1108 B.n524 B.n266 163.367
R1109 B.n528 B.n266 163.367
R1110 B.n528 B.n260 163.367
R1111 B.n537 B.n260 163.367
R1112 B.n537 B.n258 163.367
R1113 B.n541 B.n258 163.367
R1114 B.n541 B.n253 163.367
R1115 B.n551 B.n253 163.367
R1116 B.n551 B.n251 163.367
R1117 B.n555 B.n251 163.367
R1118 B.n555 B.n3 163.367
R1119 B.n635 B.n3 163.367
R1120 B.n631 B.n2 163.367
R1121 B.n631 B.n630 163.367
R1122 B.n630 B.n9 163.367
R1123 B.n626 B.n9 163.367
R1124 B.n626 B.n11 163.367
R1125 B.n622 B.n11 163.367
R1126 B.n622 B.n16 163.367
R1127 B.n618 B.n16 163.367
R1128 B.n618 B.n18 163.367
R1129 B.n614 B.n18 163.367
R1130 B.n614 B.n24 163.367
R1131 B.n610 B.n24 163.367
R1132 B.n610 B.n26 163.367
R1133 B.n606 B.n26 163.367
R1134 B.n606 B.n31 163.367
R1135 B.n602 B.n31 163.367
R1136 B.n602 B.n33 163.367
R1137 B.n598 B.n33 163.367
R1138 B.n598 B.n38 163.367
R1139 B.n594 B.n38 163.367
R1140 B.n594 B.n40 163.367
R1141 B.n492 B.n285 101.739
R1142 B.n592 B.n591 101.739
R1143 B.n89 B.n43 71.676
R1144 B.n93 B.n44 71.676
R1145 B.n97 B.n45 71.676
R1146 B.n101 B.n46 71.676
R1147 B.n105 B.n47 71.676
R1148 B.n109 B.n48 71.676
R1149 B.n113 B.n49 71.676
R1150 B.n117 B.n50 71.676
R1151 B.n121 B.n51 71.676
R1152 B.n125 B.n52 71.676
R1153 B.n129 B.n53 71.676
R1154 B.n133 B.n54 71.676
R1155 B.n137 B.n55 71.676
R1156 B.n141 B.n56 71.676
R1157 B.n145 B.n57 71.676
R1158 B.n149 B.n58 71.676
R1159 B.n153 B.n59 71.676
R1160 B.n157 B.n60 71.676
R1161 B.n161 B.n61 71.676
R1162 B.n165 B.n62 71.676
R1163 B.n169 B.n63 71.676
R1164 B.n173 B.n64 71.676
R1165 B.n177 B.n65 71.676
R1166 B.n182 B.n66 71.676
R1167 B.n186 B.n67 71.676
R1168 B.n190 B.n68 71.676
R1169 B.n194 B.n69 71.676
R1170 B.n198 B.n70 71.676
R1171 B.n202 B.n71 71.676
R1172 B.n206 B.n72 71.676
R1173 B.n210 B.n73 71.676
R1174 B.n214 B.n74 71.676
R1175 B.n218 B.n75 71.676
R1176 B.n222 B.n76 71.676
R1177 B.n226 B.n77 71.676
R1178 B.n230 B.n78 71.676
R1179 B.n234 B.n79 71.676
R1180 B.n238 B.n80 71.676
R1181 B.n242 B.n81 71.676
R1182 B.n246 B.n82 71.676
R1183 B.n83 B.n82 71.676
R1184 B.n245 B.n81 71.676
R1185 B.n241 B.n80 71.676
R1186 B.n237 B.n79 71.676
R1187 B.n233 B.n78 71.676
R1188 B.n229 B.n77 71.676
R1189 B.n225 B.n76 71.676
R1190 B.n221 B.n75 71.676
R1191 B.n217 B.n74 71.676
R1192 B.n213 B.n73 71.676
R1193 B.n209 B.n72 71.676
R1194 B.n205 B.n71 71.676
R1195 B.n201 B.n70 71.676
R1196 B.n197 B.n69 71.676
R1197 B.n193 B.n68 71.676
R1198 B.n189 B.n67 71.676
R1199 B.n185 B.n66 71.676
R1200 B.n181 B.n65 71.676
R1201 B.n176 B.n64 71.676
R1202 B.n172 B.n63 71.676
R1203 B.n168 B.n62 71.676
R1204 B.n164 B.n61 71.676
R1205 B.n160 B.n60 71.676
R1206 B.n156 B.n59 71.676
R1207 B.n152 B.n58 71.676
R1208 B.n148 B.n57 71.676
R1209 B.n144 B.n56 71.676
R1210 B.n140 B.n55 71.676
R1211 B.n136 B.n54 71.676
R1212 B.n132 B.n53 71.676
R1213 B.n128 B.n52 71.676
R1214 B.n124 B.n51 71.676
R1215 B.n120 B.n50 71.676
R1216 B.n116 B.n49 71.676
R1217 B.n112 B.n48 71.676
R1218 B.n108 B.n47 71.676
R1219 B.n104 B.n46 71.676
R1220 B.n100 B.n45 71.676
R1221 B.n96 B.n44 71.676
R1222 B.n92 B.n43 71.676
R1223 B.n491 B.n490 71.676
R1224 B.n485 B.n289 71.676
R1225 B.n482 B.n290 71.676
R1226 B.n478 B.n291 71.676
R1227 B.n474 B.n292 71.676
R1228 B.n470 B.n293 71.676
R1229 B.n466 B.n294 71.676
R1230 B.n462 B.n295 71.676
R1231 B.n458 B.n296 71.676
R1232 B.n454 B.n297 71.676
R1233 B.n450 B.n298 71.676
R1234 B.n446 B.n299 71.676
R1235 B.n442 B.n300 71.676
R1236 B.n438 B.n301 71.676
R1237 B.n434 B.n302 71.676
R1238 B.n430 B.n303 71.676
R1239 B.n426 B.n304 71.676
R1240 B.n422 B.n305 71.676
R1241 B.n417 B.n306 71.676
R1242 B.n413 B.n307 71.676
R1243 B.n409 B.n308 71.676
R1244 B.n405 B.n309 71.676
R1245 B.n401 B.n310 71.676
R1246 B.n397 B.n311 71.676
R1247 B.n393 B.n312 71.676
R1248 B.n389 B.n313 71.676
R1249 B.n385 B.n314 71.676
R1250 B.n381 B.n315 71.676
R1251 B.n377 B.n316 71.676
R1252 B.n373 B.n317 71.676
R1253 B.n369 B.n318 71.676
R1254 B.n365 B.n319 71.676
R1255 B.n361 B.n320 71.676
R1256 B.n357 B.n321 71.676
R1257 B.n353 B.n322 71.676
R1258 B.n349 B.n323 71.676
R1259 B.n345 B.n324 71.676
R1260 B.n341 B.n325 71.676
R1261 B.n337 B.n326 71.676
R1262 B.n493 B.n288 71.676
R1263 B.n491 B.n328 71.676
R1264 B.n483 B.n289 71.676
R1265 B.n479 B.n290 71.676
R1266 B.n475 B.n291 71.676
R1267 B.n471 B.n292 71.676
R1268 B.n467 B.n293 71.676
R1269 B.n463 B.n294 71.676
R1270 B.n459 B.n295 71.676
R1271 B.n455 B.n296 71.676
R1272 B.n451 B.n297 71.676
R1273 B.n447 B.n298 71.676
R1274 B.n443 B.n299 71.676
R1275 B.n439 B.n300 71.676
R1276 B.n435 B.n301 71.676
R1277 B.n431 B.n302 71.676
R1278 B.n427 B.n303 71.676
R1279 B.n423 B.n304 71.676
R1280 B.n418 B.n305 71.676
R1281 B.n414 B.n306 71.676
R1282 B.n410 B.n307 71.676
R1283 B.n406 B.n308 71.676
R1284 B.n402 B.n309 71.676
R1285 B.n398 B.n310 71.676
R1286 B.n394 B.n311 71.676
R1287 B.n390 B.n312 71.676
R1288 B.n386 B.n313 71.676
R1289 B.n382 B.n314 71.676
R1290 B.n378 B.n315 71.676
R1291 B.n374 B.n316 71.676
R1292 B.n370 B.n317 71.676
R1293 B.n366 B.n318 71.676
R1294 B.n362 B.n319 71.676
R1295 B.n358 B.n320 71.676
R1296 B.n354 B.n321 71.676
R1297 B.n350 B.n322 71.676
R1298 B.n346 B.n323 71.676
R1299 B.n342 B.n324 71.676
R1300 B.n338 B.n325 71.676
R1301 B.n334 B.n326 71.676
R1302 B.n494 B.n493 71.676
R1303 B.n636 B.n635 71.676
R1304 B.n636 B.n2 71.676
R1305 B.n88 B.n87 59.5399
R1306 B.n179 B.n85 59.5399
R1307 B.n333 B.n332 59.5399
R1308 B.n420 B.n330 59.5399
R1309 B.n499 B.n285 49.0658
R1310 B.n499 B.n280 49.0658
R1311 B.n505 B.n280 49.0658
R1312 B.n505 B.n281 49.0658
R1313 B.n511 B.n273 49.0658
R1314 B.n517 B.n273 49.0658
R1315 B.n517 B.n269 49.0658
R1316 B.n523 B.n269 49.0658
R1317 B.n523 B.n265 49.0658
R1318 B.n529 B.n265 49.0658
R1319 B.n536 B.n261 49.0658
R1320 B.n536 B.n535 49.0658
R1321 B.n542 B.n254 49.0658
R1322 B.n550 B.n254 49.0658
R1323 B.n550 B.n549 49.0658
R1324 B.n556 B.n4 49.0658
R1325 B.n634 B.n4 49.0658
R1326 B.n634 B.n633 49.0658
R1327 B.n633 B.n632 49.0658
R1328 B.n632 B.n8 49.0658
R1329 B.n625 B.n12 49.0658
R1330 B.n625 B.n624 49.0658
R1331 B.n624 B.n623 49.0658
R1332 B.n617 B.n19 49.0658
R1333 B.n617 B.n616 49.0658
R1334 B.n615 B.n23 49.0658
R1335 B.n609 B.n23 49.0658
R1336 B.n609 B.n608 49.0658
R1337 B.n608 B.n607 49.0658
R1338 B.n607 B.n30 49.0658
R1339 B.n601 B.n30 49.0658
R1340 B.n600 B.n599 49.0658
R1341 B.n599 B.n37 49.0658
R1342 B.n593 B.n37 49.0658
R1343 B.n593 B.n592 49.0658
R1344 B.n556 B.t4 39.6856
R1345 B.t0 B.n8 39.6856
R1346 B.n535 B.t3 38.2425
R1347 B.n19 B.t5 38.2425
R1348 B.n281 B.t14 36.7995
R1349 B.t7 B.n600 36.7995
R1350 B.n489 B.n283 34.4981
R1351 B.n496 B.n495 34.4981
R1352 B.n589 B.n588 34.4981
R1353 B.n90 B.n39 34.4981
R1354 B.t2 B.n261 31.0271
R1355 B.n616 B.t1 31.0271
R1356 B.n87 B.n86 22.4975
R1357 B.n85 B.n84 22.4975
R1358 B.n332 B.n331 22.4975
R1359 B.n330 B.n329 22.4975
R1360 B B.n637 18.0485
R1361 B.n529 B.t2 18.0392
R1362 B.t1 B.n615 18.0392
R1363 B.n511 B.t14 12.2668
R1364 B.n601 B.t7 12.2668
R1365 B.n542 B.t3 10.8237
R1366 B.n623 B.t5 10.8237
R1367 B.n501 B.n283 10.6151
R1368 B.n502 B.n501 10.6151
R1369 B.n503 B.n502 10.6151
R1370 B.n503 B.n275 10.6151
R1371 B.n513 B.n275 10.6151
R1372 B.n514 B.n513 10.6151
R1373 B.n515 B.n514 10.6151
R1374 B.n515 B.n267 10.6151
R1375 B.n525 B.n267 10.6151
R1376 B.n526 B.n525 10.6151
R1377 B.n527 B.n526 10.6151
R1378 B.n527 B.n259 10.6151
R1379 B.n538 B.n259 10.6151
R1380 B.n539 B.n538 10.6151
R1381 B.n540 B.n539 10.6151
R1382 B.n540 B.n252 10.6151
R1383 B.n552 B.n252 10.6151
R1384 B.n553 B.n552 10.6151
R1385 B.n554 B.n553 10.6151
R1386 B.n554 B.n0 10.6151
R1387 B.n489 B.n488 10.6151
R1388 B.n488 B.n487 10.6151
R1389 B.n487 B.n486 10.6151
R1390 B.n486 B.n484 10.6151
R1391 B.n484 B.n481 10.6151
R1392 B.n481 B.n480 10.6151
R1393 B.n480 B.n477 10.6151
R1394 B.n477 B.n476 10.6151
R1395 B.n476 B.n473 10.6151
R1396 B.n473 B.n472 10.6151
R1397 B.n472 B.n469 10.6151
R1398 B.n469 B.n468 10.6151
R1399 B.n468 B.n465 10.6151
R1400 B.n465 B.n464 10.6151
R1401 B.n464 B.n461 10.6151
R1402 B.n461 B.n460 10.6151
R1403 B.n460 B.n457 10.6151
R1404 B.n457 B.n456 10.6151
R1405 B.n456 B.n453 10.6151
R1406 B.n453 B.n452 10.6151
R1407 B.n452 B.n449 10.6151
R1408 B.n449 B.n448 10.6151
R1409 B.n448 B.n445 10.6151
R1410 B.n445 B.n444 10.6151
R1411 B.n444 B.n441 10.6151
R1412 B.n441 B.n440 10.6151
R1413 B.n440 B.n437 10.6151
R1414 B.n437 B.n436 10.6151
R1415 B.n436 B.n433 10.6151
R1416 B.n433 B.n432 10.6151
R1417 B.n432 B.n429 10.6151
R1418 B.n429 B.n428 10.6151
R1419 B.n428 B.n425 10.6151
R1420 B.n425 B.n424 10.6151
R1421 B.n424 B.n421 10.6151
R1422 B.n419 B.n416 10.6151
R1423 B.n416 B.n415 10.6151
R1424 B.n415 B.n412 10.6151
R1425 B.n412 B.n411 10.6151
R1426 B.n411 B.n408 10.6151
R1427 B.n408 B.n407 10.6151
R1428 B.n407 B.n404 10.6151
R1429 B.n404 B.n403 10.6151
R1430 B.n400 B.n399 10.6151
R1431 B.n399 B.n396 10.6151
R1432 B.n396 B.n395 10.6151
R1433 B.n395 B.n392 10.6151
R1434 B.n392 B.n391 10.6151
R1435 B.n391 B.n388 10.6151
R1436 B.n388 B.n387 10.6151
R1437 B.n387 B.n384 10.6151
R1438 B.n384 B.n383 10.6151
R1439 B.n383 B.n380 10.6151
R1440 B.n380 B.n379 10.6151
R1441 B.n379 B.n376 10.6151
R1442 B.n376 B.n375 10.6151
R1443 B.n375 B.n372 10.6151
R1444 B.n372 B.n371 10.6151
R1445 B.n371 B.n368 10.6151
R1446 B.n368 B.n367 10.6151
R1447 B.n367 B.n364 10.6151
R1448 B.n364 B.n363 10.6151
R1449 B.n363 B.n360 10.6151
R1450 B.n360 B.n359 10.6151
R1451 B.n359 B.n356 10.6151
R1452 B.n356 B.n355 10.6151
R1453 B.n355 B.n352 10.6151
R1454 B.n352 B.n351 10.6151
R1455 B.n351 B.n348 10.6151
R1456 B.n348 B.n347 10.6151
R1457 B.n347 B.n344 10.6151
R1458 B.n344 B.n343 10.6151
R1459 B.n343 B.n340 10.6151
R1460 B.n340 B.n339 10.6151
R1461 B.n339 B.n336 10.6151
R1462 B.n336 B.n335 10.6151
R1463 B.n335 B.n287 10.6151
R1464 B.n495 B.n287 10.6151
R1465 B.n497 B.n496 10.6151
R1466 B.n497 B.n278 10.6151
R1467 B.n507 B.n278 10.6151
R1468 B.n508 B.n507 10.6151
R1469 B.n509 B.n508 10.6151
R1470 B.n509 B.n271 10.6151
R1471 B.n519 B.n271 10.6151
R1472 B.n520 B.n519 10.6151
R1473 B.n521 B.n520 10.6151
R1474 B.n521 B.n263 10.6151
R1475 B.n531 B.n263 10.6151
R1476 B.n532 B.n531 10.6151
R1477 B.n533 B.n532 10.6151
R1478 B.n533 B.n256 10.6151
R1479 B.n544 B.n256 10.6151
R1480 B.n545 B.n544 10.6151
R1481 B.n547 B.n545 10.6151
R1482 B.n547 B.n546 10.6151
R1483 B.n546 B.n249 10.6151
R1484 B.n559 B.n249 10.6151
R1485 B.n560 B.n559 10.6151
R1486 B.n561 B.n560 10.6151
R1487 B.n562 B.n561 10.6151
R1488 B.n563 B.n562 10.6151
R1489 B.n566 B.n563 10.6151
R1490 B.n567 B.n566 10.6151
R1491 B.n568 B.n567 10.6151
R1492 B.n569 B.n568 10.6151
R1493 B.n571 B.n569 10.6151
R1494 B.n572 B.n571 10.6151
R1495 B.n573 B.n572 10.6151
R1496 B.n574 B.n573 10.6151
R1497 B.n576 B.n574 10.6151
R1498 B.n577 B.n576 10.6151
R1499 B.n578 B.n577 10.6151
R1500 B.n579 B.n578 10.6151
R1501 B.n581 B.n579 10.6151
R1502 B.n582 B.n581 10.6151
R1503 B.n583 B.n582 10.6151
R1504 B.n584 B.n583 10.6151
R1505 B.n586 B.n584 10.6151
R1506 B.n587 B.n586 10.6151
R1507 B.n588 B.n587 10.6151
R1508 B.n629 B.n1 10.6151
R1509 B.n629 B.n628 10.6151
R1510 B.n628 B.n627 10.6151
R1511 B.n627 B.n10 10.6151
R1512 B.n621 B.n10 10.6151
R1513 B.n621 B.n620 10.6151
R1514 B.n620 B.n619 10.6151
R1515 B.n619 B.n17 10.6151
R1516 B.n613 B.n17 10.6151
R1517 B.n613 B.n612 10.6151
R1518 B.n612 B.n611 10.6151
R1519 B.n611 B.n25 10.6151
R1520 B.n605 B.n25 10.6151
R1521 B.n605 B.n604 10.6151
R1522 B.n604 B.n603 10.6151
R1523 B.n603 B.n32 10.6151
R1524 B.n597 B.n32 10.6151
R1525 B.n597 B.n596 10.6151
R1526 B.n596 B.n595 10.6151
R1527 B.n595 B.n39 10.6151
R1528 B.n91 B.n90 10.6151
R1529 B.n94 B.n91 10.6151
R1530 B.n95 B.n94 10.6151
R1531 B.n98 B.n95 10.6151
R1532 B.n99 B.n98 10.6151
R1533 B.n102 B.n99 10.6151
R1534 B.n103 B.n102 10.6151
R1535 B.n106 B.n103 10.6151
R1536 B.n107 B.n106 10.6151
R1537 B.n110 B.n107 10.6151
R1538 B.n111 B.n110 10.6151
R1539 B.n114 B.n111 10.6151
R1540 B.n115 B.n114 10.6151
R1541 B.n118 B.n115 10.6151
R1542 B.n119 B.n118 10.6151
R1543 B.n122 B.n119 10.6151
R1544 B.n123 B.n122 10.6151
R1545 B.n126 B.n123 10.6151
R1546 B.n127 B.n126 10.6151
R1547 B.n130 B.n127 10.6151
R1548 B.n131 B.n130 10.6151
R1549 B.n134 B.n131 10.6151
R1550 B.n135 B.n134 10.6151
R1551 B.n138 B.n135 10.6151
R1552 B.n139 B.n138 10.6151
R1553 B.n142 B.n139 10.6151
R1554 B.n143 B.n142 10.6151
R1555 B.n146 B.n143 10.6151
R1556 B.n147 B.n146 10.6151
R1557 B.n150 B.n147 10.6151
R1558 B.n151 B.n150 10.6151
R1559 B.n154 B.n151 10.6151
R1560 B.n155 B.n154 10.6151
R1561 B.n158 B.n155 10.6151
R1562 B.n159 B.n158 10.6151
R1563 B.n163 B.n162 10.6151
R1564 B.n166 B.n163 10.6151
R1565 B.n167 B.n166 10.6151
R1566 B.n170 B.n167 10.6151
R1567 B.n171 B.n170 10.6151
R1568 B.n174 B.n171 10.6151
R1569 B.n175 B.n174 10.6151
R1570 B.n178 B.n175 10.6151
R1571 B.n183 B.n180 10.6151
R1572 B.n184 B.n183 10.6151
R1573 B.n187 B.n184 10.6151
R1574 B.n188 B.n187 10.6151
R1575 B.n191 B.n188 10.6151
R1576 B.n192 B.n191 10.6151
R1577 B.n195 B.n192 10.6151
R1578 B.n196 B.n195 10.6151
R1579 B.n199 B.n196 10.6151
R1580 B.n200 B.n199 10.6151
R1581 B.n203 B.n200 10.6151
R1582 B.n204 B.n203 10.6151
R1583 B.n207 B.n204 10.6151
R1584 B.n208 B.n207 10.6151
R1585 B.n211 B.n208 10.6151
R1586 B.n212 B.n211 10.6151
R1587 B.n215 B.n212 10.6151
R1588 B.n216 B.n215 10.6151
R1589 B.n219 B.n216 10.6151
R1590 B.n220 B.n219 10.6151
R1591 B.n223 B.n220 10.6151
R1592 B.n224 B.n223 10.6151
R1593 B.n227 B.n224 10.6151
R1594 B.n228 B.n227 10.6151
R1595 B.n231 B.n228 10.6151
R1596 B.n232 B.n231 10.6151
R1597 B.n235 B.n232 10.6151
R1598 B.n236 B.n235 10.6151
R1599 B.n239 B.n236 10.6151
R1600 B.n240 B.n239 10.6151
R1601 B.n243 B.n240 10.6151
R1602 B.n244 B.n243 10.6151
R1603 B.n247 B.n244 10.6151
R1604 B.n248 B.n247 10.6151
R1605 B.n589 B.n248 10.6151
R1606 B.n549 B.t4 9.38063
R1607 B.n12 B.t0 9.38063
R1608 B.n637 B.n0 8.11757
R1609 B.n637 B.n1 8.11757
R1610 B.n420 B.n419 6.5566
R1611 B.n403 B.n333 6.5566
R1612 B.n162 B.n88 6.5566
R1613 B.n179 B.n178 6.5566
R1614 B.n421 B.n420 4.05904
R1615 B.n400 B.n333 4.05904
R1616 B.n159 B.n88 4.05904
R1617 B.n180 B.n179 4.05904
R1618 VN.n1 VN.t1 352.361
R1619 VN.n7 VN.t3 352.361
R1620 VN.n4 VN.t0 337.111
R1621 VN.n10 VN.t5 337.111
R1622 VN.n2 VN.t4 289.49
R1623 VN.n8 VN.t2 289.49
R1624 VN.n9 VN.n6 161.3
R1625 VN.n3 VN.n0 161.3
R1626 VN.n11 VN.n10 80.6037
R1627 VN.n5 VN.n4 80.6037
R1628 VN.n4 VN.n3 56.2746
R1629 VN.n10 VN.n9 56.2746
R1630 VN.n7 VN.n6 43.9052
R1631 VN.n1 VN.n0 43.9052
R1632 VN.n2 VN.n1 42.6471
R1633 VN.n8 VN.n7 42.6471
R1634 VN VN.n11 40.59
R1635 VN.n3 VN.n2 12.234
R1636 VN.n9 VN.n8 12.234
R1637 VN.n11 VN.n6 0.285035
R1638 VN.n5 VN.n0 0.285035
R1639 VN VN.n5 0.146778
R1640 VDD2.n103 VDD2.n55 289.615
R1641 VDD2.n48 VDD2.n0 289.615
R1642 VDD2.n104 VDD2.n103 185
R1643 VDD2.n102 VDD2.n101 185
R1644 VDD2.n59 VDD2.n58 185
R1645 VDD2.n96 VDD2.n95 185
R1646 VDD2.n94 VDD2.n61 185
R1647 VDD2.n93 VDD2.n92 185
R1648 VDD2.n64 VDD2.n62 185
R1649 VDD2.n87 VDD2.n86 185
R1650 VDD2.n85 VDD2.n84 185
R1651 VDD2.n68 VDD2.n67 185
R1652 VDD2.n79 VDD2.n78 185
R1653 VDD2.n77 VDD2.n76 185
R1654 VDD2.n72 VDD2.n71 185
R1655 VDD2.n16 VDD2.n15 185
R1656 VDD2.n21 VDD2.n20 185
R1657 VDD2.n23 VDD2.n22 185
R1658 VDD2.n12 VDD2.n11 185
R1659 VDD2.n29 VDD2.n28 185
R1660 VDD2.n31 VDD2.n30 185
R1661 VDD2.n8 VDD2.n7 185
R1662 VDD2.n38 VDD2.n37 185
R1663 VDD2.n39 VDD2.n6 185
R1664 VDD2.n41 VDD2.n40 185
R1665 VDD2.n4 VDD2.n3 185
R1666 VDD2.n47 VDD2.n46 185
R1667 VDD2.n49 VDD2.n48 185
R1668 VDD2.n73 VDD2.t0 149.524
R1669 VDD2.n17 VDD2.t4 149.524
R1670 VDD2.n103 VDD2.n102 104.615
R1671 VDD2.n102 VDD2.n58 104.615
R1672 VDD2.n95 VDD2.n58 104.615
R1673 VDD2.n95 VDD2.n94 104.615
R1674 VDD2.n94 VDD2.n93 104.615
R1675 VDD2.n93 VDD2.n62 104.615
R1676 VDD2.n86 VDD2.n62 104.615
R1677 VDD2.n86 VDD2.n85 104.615
R1678 VDD2.n85 VDD2.n67 104.615
R1679 VDD2.n78 VDD2.n67 104.615
R1680 VDD2.n78 VDD2.n77 104.615
R1681 VDD2.n77 VDD2.n71 104.615
R1682 VDD2.n21 VDD2.n15 104.615
R1683 VDD2.n22 VDD2.n21 104.615
R1684 VDD2.n22 VDD2.n11 104.615
R1685 VDD2.n29 VDD2.n11 104.615
R1686 VDD2.n30 VDD2.n29 104.615
R1687 VDD2.n30 VDD2.n7 104.615
R1688 VDD2.n38 VDD2.n7 104.615
R1689 VDD2.n39 VDD2.n38 104.615
R1690 VDD2.n40 VDD2.n39 104.615
R1691 VDD2.n40 VDD2.n3 104.615
R1692 VDD2.n47 VDD2.n3 104.615
R1693 VDD2.n48 VDD2.n47 104.615
R1694 VDD2.n54 VDD2.n53 63.0287
R1695 VDD2 VDD2.n109 63.0259
R1696 VDD2.t0 VDD2.n71 52.3082
R1697 VDD2.t4 VDD2.n15 52.3082
R1698 VDD2.n54 VDD2.n52 49.7527
R1699 VDD2.n108 VDD2.n107 49.0581
R1700 VDD2.n108 VDD2.n54 35.5601
R1701 VDD2.n96 VDD2.n61 13.1884
R1702 VDD2.n41 VDD2.n6 13.1884
R1703 VDD2.n97 VDD2.n59 12.8005
R1704 VDD2.n92 VDD2.n63 12.8005
R1705 VDD2.n37 VDD2.n36 12.8005
R1706 VDD2.n42 VDD2.n4 12.8005
R1707 VDD2.n101 VDD2.n100 12.0247
R1708 VDD2.n91 VDD2.n64 12.0247
R1709 VDD2.n35 VDD2.n8 12.0247
R1710 VDD2.n46 VDD2.n45 12.0247
R1711 VDD2.n104 VDD2.n57 11.249
R1712 VDD2.n88 VDD2.n87 11.249
R1713 VDD2.n32 VDD2.n31 11.249
R1714 VDD2.n49 VDD2.n2 11.249
R1715 VDD2.n105 VDD2.n55 10.4732
R1716 VDD2.n84 VDD2.n66 10.4732
R1717 VDD2.n28 VDD2.n10 10.4732
R1718 VDD2.n50 VDD2.n0 10.4732
R1719 VDD2.n73 VDD2.n72 10.2747
R1720 VDD2.n17 VDD2.n16 10.2747
R1721 VDD2.n83 VDD2.n68 9.69747
R1722 VDD2.n27 VDD2.n12 9.69747
R1723 VDD2.n107 VDD2.n106 9.45567
R1724 VDD2.n52 VDD2.n51 9.45567
R1725 VDD2.n75 VDD2.n74 9.3005
R1726 VDD2.n70 VDD2.n69 9.3005
R1727 VDD2.n81 VDD2.n80 9.3005
R1728 VDD2.n83 VDD2.n82 9.3005
R1729 VDD2.n66 VDD2.n65 9.3005
R1730 VDD2.n89 VDD2.n88 9.3005
R1731 VDD2.n91 VDD2.n90 9.3005
R1732 VDD2.n63 VDD2.n60 9.3005
R1733 VDD2.n106 VDD2.n105 9.3005
R1734 VDD2.n57 VDD2.n56 9.3005
R1735 VDD2.n100 VDD2.n99 9.3005
R1736 VDD2.n98 VDD2.n97 9.3005
R1737 VDD2.n51 VDD2.n50 9.3005
R1738 VDD2.n2 VDD2.n1 9.3005
R1739 VDD2.n45 VDD2.n44 9.3005
R1740 VDD2.n43 VDD2.n42 9.3005
R1741 VDD2.n19 VDD2.n18 9.3005
R1742 VDD2.n14 VDD2.n13 9.3005
R1743 VDD2.n25 VDD2.n24 9.3005
R1744 VDD2.n27 VDD2.n26 9.3005
R1745 VDD2.n10 VDD2.n9 9.3005
R1746 VDD2.n33 VDD2.n32 9.3005
R1747 VDD2.n35 VDD2.n34 9.3005
R1748 VDD2.n36 VDD2.n5 9.3005
R1749 VDD2.n80 VDD2.n79 8.92171
R1750 VDD2.n24 VDD2.n23 8.92171
R1751 VDD2.n76 VDD2.n70 8.14595
R1752 VDD2.n20 VDD2.n14 8.14595
R1753 VDD2.n75 VDD2.n72 7.3702
R1754 VDD2.n19 VDD2.n16 7.3702
R1755 VDD2.n76 VDD2.n75 5.81868
R1756 VDD2.n20 VDD2.n19 5.81868
R1757 VDD2.n79 VDD2.n70 5.04292
R1758 VDD2.n23 VDD2.n14 5.04292
R1759 VDD2.n80 VDD2.n68 4.26717
R1760 VDD2.n24 VDD2.n12 4.26717
R1761 VDD2.n107 VDD2.n55 3.49141
R1762 VDD2.n84 VDD2.n83 3.49141
R1763 VDD2.n28 VDD2.n27 3.49141
R1764 VDD2.n52 VDD2.n0 3.49141
R1765 VDD2.n74 VDD2.n73 2.84303
R1766 VDD2.n18 VDD2.n17 2.84303
R1767 VDD2.n105 VDD2.n104 2.71565
R1768 VDD2.n87 VDD2.n66 2.71565
R1769 VDD2.n31 VDD2.n10 2.71565
R1770 VDD2.n50 VDD2.n49 2.71565
R1771 VDD2.n109 VDD2.t3 1.98646
R1772 VDD2.n109 VDD2.t2 1.98646
R1773 VDD2.n53 VDD2.t1 1.98646
R1774 VDD2.n53 VDD2.t5 1.98646
R1775 VDD2.n101 VDD2.n57 1.93989
R1776 VDD2.n88 VDD2.n64 1.93989
R1777 VDD2.n32 VDD2.n8 1.93989
R1778 VDD2.n46 VDD2.n2 1.93989
R1779 VDD2.n100 VDD2.n59 1.16414
R1780 VDD2.n92 VDD2.n91 1.16414
R1781 VDD2.n37 VDD2.n35 1.16414
R1782 VDD2.n45 VDD2.n4 1.16414
R1783 VDD2 VDD2.n108 0.80869
R1784 VDD2.n97 VDD2.n96 0.388379
R1785 VDD2.n63 VDD2.n61 0.388379
R1786 VDD2.n36 VDD2.n6 0.388379
R1787 VDD2.n42 VDD2.n41 0.388379
R1788 VDD2.n106 VDD2.n56 0.155672
R1789 VDD2.n99 VDD2.n56 0.155672
R1790 VDD2.n99 VDD2.n98 0.155672
R1791 VDD2.n98 VDD2.n60 0.155672
R1792 VDD2.n90 VDD2.n60 0.155672
R1793 VDD2.n90 VDD2.n89 0.155672
R1794 VDD2.n89 VDD2.n65 0.155672
R1795 VDD2.n82 VDD2.n65 0.155672
R1796 VDD2.n82 VDD2.n81 0.155672
R1797 VDD2.n81 VDD2.n69 0.155672
R1798 VDD2.n74 VDD2.n69 0.155672
R1799 VDD2.n18 VDD2.n13 0.155672
R1800 VDD2.n25 VDD2.n13 0.155672
R1801 VDD2.n26 VDD2.n25 0.155672
R1802 VDD2.n26 VDD2.n9 0.155672
R1803 VDD2.n33 VDD2.n9 0.155672
R1804 VDD2.n34 VDD2.n33 0.155672
R1805 VDD2.n34 VDD2.n5 0.155672
R1806 VDD2.n43 VDD2.n5 0.155672
R1807 VDD2.n44 VDD2.n43 0.155672
R1808 VDD2.n44 VDD2.n1 0.155672
R1809 VDD2.n51 VDD2.n1 0.155672
C0 VDD1 VP 4.11475f
C1 VDD1 VTAIL 8.1008f
C2 VN VDD2 3.95846f
C3 VN VP 4.83429f
C4 VTAIL VN 3.76225f
C5 VDD1 VN 0.148378f
C6 VDD2 VP 0.308355f
C7 VTAIL VDD2 8.13728f
C8 VTAIL VP 3.77674f
C9 VDD1 VDD2 0.757858f
C10 VDD2 B 4.230444f
C11 VDD1 B 4.259959f
C12 VTAIL B 5.759612f
C13 VN B 7.842609f
C14 VP B 6.042457f
C15 VDD2.n0 B 0.030448f
C16 VDD2.n1 B 0.02287f
C17 VDD2.n2 B 0.012289f
C18 VDD2.n3 B 0.029048f
C19 VDD2.n4 B 0.013012f
C20 VDD2.n5 B 0.02287f
C21 VDD2.n6 B 0.012651f
C22 VDD2.n7 B 0.029048f
C23 VDD2.n8 B 0.013012f
C24 VDD2.n9 B 0.02287f
C25 VDD2.n10 B 0.012289f
C26 VDD2.n11 B 0.029048f
C27 VDD2.n12 B 0.013012f
C28 VDD2.n13 B 0.02287f
C29 VDD2.n14 B 0.012289f
C30 VDD2.n15 B 0.021786f
C31 VDD2.n16 B 0.020534f
C32 VDD2.t4 B 0.048811f
C33 VDD2.n17 B 0.147069f
C34 VDD2.n18 B 0.947252f
C35 VDD2.n19 B 0.012289f
C36 VDD2.n20 B 0.013012f
C37 VDD2.n21 B 0.029048f
C38 VDD2.n22 B 0.029048f
C39 VDD2.n23 B 0.013012f
C40 VDD2.n24 B 0.012289f
C41 VDD2.n25 B 0.02287f
C42 VDD2.n26 B 0.02287f
C43 VDD2.n27 B 0.012289f
C44 VDD2.n28 B 0.013012f
C45 VDD2.n29 B 0.029048f
C46 VDD2.n30 B 0.029048f
C47 VDD2.n31 B 0.013012f
C48 VDD2.n32 B 0.012289f
C49 VDD2.n33 B 0.02287f
C50 VDD2.n34 B 0.02287f
C51 VDD2.n35 B 0.012289f
C52 VDD2.n36 B 0.012289f
C53 VDD2.n37 B 0.013012f
C54 VDD2.n38 B 0.029048f
C55 VDD2.n39 B 0.029048f
C56 VDD2.n40 B 0.029048f
C57 VDD2.n41 B 0.012651f
C58 VDD2.n42 B 0.012289f
C59 VDD2.n43 B 0.02287f
C60 VDD2.n44 B 0.02287f
C61 VDD2.n45 B 0.012289f
C62 VDD2.n46 B 0.013012f
C63 VDD2.n47 B 0.029048f
C64 VDD2.n48 B 0.059881f
C65 VDD2.n49 B 0.013012f
C66 VDD2.n50 B 0.012289f
C67 VDD2.n51 B 0.053175f
C68 VDD2.n52 B 0.050339f
C69 VDD2.t1 B 0.180184f
C70 VDD2.t5 B 0.180184f
C71 VDD2.n53 B 1.58722f
C72 VDD2.n54 B 1.63255f
C73 VDD2.n55 B 0.030448f
C74 VDD2.n56 B 0.02287f
C75 VDD2.n57 B 0.012289f
C76 VDD2.n58 B 0.029048f
C77 VDD2.n59 B 0.013012f
C78 VDD2.n60 B 0.02287f
C79 VDD2.n61 B 0.012651f
C80 VDD2.n62 B 0.029048f
C81 VDD2.n63 B 0.012289f
C82 VDD2.n64 B 0.013012f
C83 VDD2.n65 B 0.02287f
C84 VDD2.n66 B 0.012289f
C85 VDD2.n67 B 0.029048f
C86 VDD2.n68 B 0.013012f
C87 VDD2.n69 B 0.02287f
C88 VDD2.n70 B 0.012289f
C89 VDD2.n71 B 0.021786f
C90 VDD2.n72 B 0.020534f
C91 VDD2.t0 B 0.048811f
C92 VDD2.n73 B 0.147069f
C93 VDD2.n74 B 0.947252f
C94 VDD2.n75 B 0.012289f
C95 VDD2.n76 B 0.013012f
C96 VDD2.n77 B 0.029048f
C97 VDD2.n78 B 0.029048f
C98 VDD2.n79 B 0.013012f
C99 VDD2.n80 B 0.012289f
C100 VDD2.n81 B 0.02287f
C101 VDD2.n82 B 0.02287f
C102 VDD2.n83 B 0.012289f
C103 VDD2.n84 B 0.013012f
C104 VDD2.n85 B 0.029048f
C105 VDD2.n86 B 0.029048f
C106 VDD2.n87 B 0.013012f
C107 VDD2.n88 B 0.012289f
C108 VDD2.n89 B 0.02287f
C109 VDD2.n90 B 0.02287f
C110 VDD2.n91 B 0.012289f
C111 VDD2.n92 B 0.013012f
C112 VDD2.n93 B 0.029048f
C113 VDD2.n94 B 0.029048f
C114 VDD2.n95 B 0.029048f
C115 VDD2.n96 B 0.012651f
C116 VDD2.n97 B 0.012289f
C117 VDD2.n98 B 0.02287f
C118 VDD2.n99 B 0.02287f
C119 VDD2.n100 B 0.012289f
C120 VDD2.n101 B 0.013012f
C121 VDD2.n102 B 0.029048f
C122 VDD2.n103 B 0.059881f
C123 VDD2.n104 B 0.013012f
C124 VDD2.n105 B 0.012289f
C125 VDD2.n106 B 0.053175f
C126 VDD2.n107 B 0.048996f
C127 VDD2.n108 B 1.75661f
C128 VDD2.t3 B 0.180184f
C129 VDD2.t2 B 0.180184f
C130 VDD2.n109 B 1.5872f
C131 VN.n0 B 0.19151f
C132 VN.t4 B 0.974f
C133 VN.t1 B 1.04776f
C134 VN.n1 B 0.424986f
C135 VN.n2 B 0.413729f
C136 VN.n3 B 0.053075f
C137 VN.t0 B 1.02925f
C138 VN.n4 B 0.427426f
C139 VN.n5 B 0.040695f
C140 VN.n6 B 0.19151f
C141 VN.t2 B 0.974f
C142 VN.t3 B 1.04776f
C143 VN.n7 B 0.424986f
C144 VN.n8 B 0.413729f
C145 VN.n9 B 0.053075f
C146 VN.t5 B 1.02925f
C147 VN.n10 B 0.427426f
C148 VN.n11 B 1.7129f
C149 VTAIL.t0 B 0.191159f
C150 VTAIL.t5 B 0.191159f
C151 VTAIL.n0 B 1.6132f
C152 VTAIL.n1 B 0.334392f
C153 VTAIL.n2 B 0.032303f
C154 VTAIL.n3 B 0.024263f
C155 VTAIL.n4 B 0.013038f
C156 VTAIL.n5 B 0.030817f
C157 VTAIL.n6 B 0.013805f
C158 VTAIL.n7 B 0.024263f
C159 VTAIL.n8 B 0.013421f
C160 VTAIL.n9 B 0.030817f
C161 VTAIL.n10 B 0.013805f
C162 VTAIL.n11 B 0.024263f
C163 VTAIL.n12 B 0.013038f
C164 VTAIL.n13 B 0.030817f
C165 VTAIL.n14 B 0.013805f
C166 VTAIL.n15 B 0.024263f
C167 VTAIL.n16 B 0.013038f
C168 VTAIL.n17 B 0.023113f
C169 VTAIL.n18 B 0.021785f
C170 VTAIL.t9 B 0.051784f
C171 VTAIL.n19 B 0.156028f
C172 VTAIL.n20 B 1.00495f
C173 VTAIL.n21 B 0.013038f
C174 VTAIL.n22 B 0.013805f
C175 VTAIL.n23 B 0.030817f
C176 VTAIL.n24 B 0.030817f
C177 VTAIL.n25 B 0.013805f
C178 VTAIL.n26 B 0.013038f
C179 VTAIL.n27 B 0.024263f
C180 VTAIL.n28 B 0.024263f
C181 VTAIL.n29 B 0.013038f
C182 VTAIL.n30 B 0.013805f
C183 VTAIL.n31 B 0.030817f
C184 VTAIL.n32 B 0.030817f
C185 VTAIL.n33 B 0.013805f
C186 VTAIL.n34 B 0.013038f
C187 VTAIL.n35 B 0.024263f
C188 VTAIL.n36 B 0.024263f
C189 VTAIL.n37 B 0.013038f
C190 VTAIL.n38 B 0.013038f
C191 VTAIL.n39 B 0.013805f
C192 VTAIL.n40 B 0.030817f
C193 VTAIL.n41 B 0.030817f
C194 VTAIL.n42 B 0.030817f
C195 VTAIL.n43 B 0.013421f
C196 VTAIL.n44 B 0.013038f
C197 VTAIL.n45 B 0.024263f
C198 VTAIL.n46 B 0.024263f
C199 VTAIL.n47 B 0.013038f
C200 VTAIL.n48 B 0.013805f
C201 VTAIL.n49 B 0.030817f
C202 VTAIL.n50 B 0.063529f
C203 VTAIL.n51 B 0.013805f
C204 VTAIL.n52 B 0.013038f
C205 VTAIL.n53 B 0.056414f
C206 VTAIL.n54 B 0.03523f
C207 VTAIL.n55 B 0.174913f
C208 VTAIL.t8 B 0.191159f
C209 VTAIL.t7 B 0.191159f
C210 VTAIL.n56 B 1.6132f
C211 VTAIL.n57 B 1.47056f
C212 VTAIL.t2 B 0.191159f
C213 VTAIL.t3 B 0.191159f
C214 VTAIL.n58 B 1.61321f
C215 VTAIL.n59 B 1.47055f
C216 VTAIL.n60 B 0.032303f
C217 VTAIL.n61 B 0.024263f
C218 VTAIL.n62 B 0.013038f
C219 VTAIL.n63 B 0.030817f
C220 VTAIL.n64 B 0.013805f
C221 VTAIL.n65 B 0.024263f
C222 VTAIL.n66 B 0.013421f
C223 VTAIL.n67 B 0.030817f
C224 VTAIL.n68 B 0.013038f
C225 VTAIL.n69 B 0.013805f
C226 VTAIL.n70 B 0.024263f
C227 VTAIL.n71 B 0.013038f
C228 VTAIL.n72 B 0.030817f
C229 VTAIL.n73 B 0.013805f
C230 VTAIL.n74 B 0.024263f
C231 VTAIL.n75 B 0.013038f
C232 VTAIL.n76 B 0.023113f
C233 VTAIL.n77 B 0.021785f
C234 VTAIL.t4 B 0.051784f
C235 VTAIL.n78 B 0.156028f
C236 VTAIL.n79 B 1.00495f
C237 VTAIL.n80 B 0.013038f
C238 VTAIL.n81 B 0.013805f
C239 VTAIL.n82 B 0.030817f
C240 VTAIL.n83 B 0.030817f
C241 VTAIL.n84 B 0.013805f
C242 VTAIL.n85 B 0.013038f
C243 VTAIL.n86 B 0.024263f
C244 VTAIL.n87 B 0.024263f
C245 VTAIL.n88 B 0.013038f
C246 VTAIL.n89 B 0.013805f
C247 VTAIL.n90 B 0.030817f
C248 VTAIL.n91 B 0.030817f
C249 VTAIL.n92 B 0.013805f
C250 VTAIL.n93 B 0.013038f
C251 VTAIL.n94 B 0.024263f
C252 VTAIL.n95 B 0.024263f
C253 VTAIL.n96 B 0.013038f
C254 VTAIL.n97 B 0.013805f
C255 VTAIL.n98 B 0.030817f
C256 VTAIL.n99 B 0.030817f
C257 VTAIL.n100 B 0.030817f
C258 VTAIL.n101 B 0.013421f
C259 VTAIL.n102 B 0.013038f
C260 VTAIL.n103 B 0.024263f
C261 VTAIL.n104 B 0.024263f
C262 VTAIL.n105 B 0.013038f
C263 VTAIL.n106 B 0.013805f
C264 VTAIL.n107 B 0.030817f
C265 VTAIL.n108 B 0.063529f
C266 VTAIL.n109 B 0.013805f
C267 VTAIL.n110 B 0.013038f
C268 VTAIL.n111 B 0.056414f
C269 VTAIL.n112 B 0.03523f
C270 VTAIL.n113 B 0.174913f
C271 VTAIL.t10 B 0.191159f
C272 VTAIL.t11 B 0.191159f
C273 VTAIL.n114 B 1.61321f
C274 VTAIL.n115 B 0.388469f
C275 VTAIL.n116 B 0.032303f
C276 VTAIL.n117 B 0.024263f
C277 VTAIL.n118 B 0.013038f
C278 VTAIL.n119 B 0.030817f
C279 VTAIL.n120 B 0.013805f
C280 VTAIL.n121 B 0.024263f
C281 VTAIL.n122 B 0.013421f
C282 VTAIL.n123 B 0.030817f
C283 VTAIL.n124 B 0.013038f
C284 VTAIL.n125 B 0.013805f
C285 VTAIL.n126 B 0.024263f
C286 VTAIL.n127 B 0.013038f
C287 VTAIL.n128 B 0.030817f
C288 VTAIL.n129 B 0.013805f
C289 VTAIL.n130 B 0.024263f
C290 VTAIL.n131 B 0.013038f
C291 VTAIL.n132 B 0.023113f
C292 VTAIL.n133 B 0.021785f
C293 VTAIL.t6 B 0.051784f
C294 VTAIL.n134 B 0.156028f
C295 VTAIL.n135 B 1.00495f
C296 VTAIL.n136 B 0.013038f
C297 VTAIL.n137 B 0.013805f
C298 VTAIL.n138 B 0.030817f
C299 VTAIL.n139 B 0.030817f
C300 VTAIL.n140 B 0.013805f
C301 VTAIL.n141 B 0.013038f
C302 VTAIL.n142 B 0.024263f
C303 VTAIL.n143 B 0.024263f
C304 VTAIL.n144 B 0.013038f
C305 VTAIL.n145 B 0.013805f
C306 VTAIL.n146 B 0.030817f
C307 VTAIL.n147 B 0.030817f
C308 VTAIL.n148 B 0.013805f
C309 VTAIL.n149 B 0.013038f
C310 VTAIL.n150 B 0.024263f
C311 VTAIL.n151 B 0.024263f
C312 VTAIL.n152 B 0.013038f
C313 VTAIL.n153 B 0.013805f
C314 VTAIL.n154 B 0.030817f
C315 VTAIL.n155 B 0.030817f
C316 VTAIL.n156 B 0.030817f
C317 VTAIL.n157 B 0.013421f
C318 VTAIL.n158 B 0.013038f
C319 VTAIL.n159 B 0.024263f
C320 VTAIL.n160 B 0.024263f
C321 VTAIL.n161 B 0.013038f
C322 VTAIL.n162 B 0.013805f
C323 VTAIL.n163 B 0.030817f
C324 VTAIL.n164 B 0.063529f
C325 VTAIL.n165 B 0.013805f
C326 VTAIL.n166 B 0.013038f
C327 VTAIL.n167 B 0.056414f
C328 VTAIL.n168 B 0.03523f
C329 VTAIL.n169 B 1.17881f
C330 VTAIL.n170 B 0.032303f
C331 VTAIL.n171 B 0.024263f
C332 VTAIL.n172 B 0.013038f
C333 VTAIL.n173 B 0.030817f
C334 VTAIL.n174 B 0.013805f
C335 VTAIL.n175 B 0.024263f
C336 VTAIL.n176 B 0.013421f
C337 VTAIL.n177 B 0.030817f
C338 VTAIL.n178 B 0.013805f
C339 VTAIL.n179 B 0.024263f
C340 VTAIL.n180 B 0.013038f
C341 VTAIL.n181 B 0.030817f
C342 VTAIL.n182 B 0.013805f
C343 VTAIL.n183 B 0.024263f
C344 VTAIL.n184 B 0.013038f
C345 VTAIL.n185 B 0.023113f
C346 VTAIL.n186 B 0.021785f
C347 VTAIL.t1 B 0.051784f
C348 VTAIL.n187 B 0.156028f
C349 VTAIL.n188 B 1.00495f
C350 VTAIL.n189 B 0.013038f
C351 VTAIL.n190 B 0.013805f
C352 VTAIL.n191 B 0.030817f
C353 VTAIL.n192 B 0.030817f
C354 VTAIL.n193 B 0.013805f
C355 VTAIL.n194 B 0.013038f
C356 VTAIL.n195 B 0.024263f
C357 VTAIL.n196 B 0.024263f
C358 VTAIL.n197 B 0.013038f
C359 VTAIL.n198 B 0.013805f
C360 VTAIL.n199 B 0.030817f
C361 VTAIL.n200 B 0.030817f
C362 VTAIL.n201 B 0.013805f
C363 VTAIL.n202 B 0.013038f
C364 VTAIL.n203 B 0.024263f
C365 VTAIL.n204 B 0.024263f
C366 VTAIL.n205 B 0.013038f
C367 VTAIL.n206 B 0.013038f
C368 VTAIL.n207 B 0.013805f
C369 VTAIL.n208 B 0.030817f
C370 VTAIL.n209 B 0.030817f
C371 VTAIL.n210 B 0.030817f
C372 VTAIL.n211 B 0.013421f
C373 VTAIL.n212 B 0.013038f
C374 VTAIL.n213 B 0.024263f
C375 VTAIL.n214 B 0.024263f
C376 VTAIL.n215 B 0.013038f
C377 VTAIL.n216 B 0.013805f
C378 VTAIL.n217 B 0.030817f
C379 VTAIL.n218 B 0.063529f
C380 VTAIL.n219 B 0.013805f
C381 VTAIL.n220 B 0.013038f
C382 VTAIL.n221 B 0.056414f
C383 VTAIL.n222 B 0.03523f
C384 VTAIL.n223 B 1.15472f
C385 VDD1.n0 B 0.030487f
C386 VDD1.n1 B 0.022899f
C387 VDD1.n2 B 0.012305f
C388 VDD1.n3 B 0.029085f
C389 VDD1.n4 B 0.013029f
C390 VDD1.n5 B 0.022899f
C391 VDD1.n6 B 0.012667f
C392 VDD1.n7 B 0.029085f
C393 VDD1.n8 B 0.012305f
C394 VDD1.n9 B 0.013029f
C395 VDD1.n10 B 0.022899f
C396 VDD1.n11 B 0.012305f
C397 VDD1.n12 B 0.029085f
C398 VDD1.n13 B 0.013029f
C399 VDD1.n14 B 0.022899f
C400 VDD1.n15 B 0.012305f
C401 VDD1.n16 B 0.021813f
C402 VDD1.n17 B 0.020561f
C403 VDD1.t0 B 0.048873f
C404 VDD1.n18 B 0.147257f
C405 VDD1.n19 B 0.948459f
C406 VDD1.n20 B 0.012305f
C407 VDD1.n21 B 0.013029f
C408 VDD1.n22 B 0.029085f
C409 VDD1.n23 B 0.029085f
C410 VDD1.n24 B 0.013029f
C411 VDD1.n25 B 0.012305f
C412 VDD1.n26 B 0.022899f
C413 VDD1.n27 B 0.022899f
C414 VDD1.n28 B 0.012305f
C415 VDD1.n29 B 0.013029f
C416 VDD1.n30 B 0.029085f
C417 VDD1.n31 B 0.029085f
C418 VDD1.n32 B 0.013029f
C419 VDD1.n33 B 0.012305f
C420 VDD1.n34 B 0.022899f
C421 VDD1.n35 B 0.022899f
C422 VDD1.n36 B 0.012305f
C423 VDD1.n37 B 0.013029f
C424 VDD1.n38 B 0.029085f
C425 VDD1.n39 B 0.029085f
C426 VDD1.n40 B 0.029085f
C427 VDD1.n41 B 0.012667f
C428 VDD1.n42 B 0.012305f
C429 VDD1.n43 B 0.022899f
C430 VDD1.n44 B 0.022899f
C431 VDD1.n45 B 0.012305f
C432 VDD1.n46 B 0.013029f
C433 VDD1.n47 B 0.029085f
C434 VDD1.n48 B 0.059958f
C435 VDD1.n49 B 0.013029f
C436 VDD1.n50 B 0.012305f
C437 VDD1.n51 B 0.053243f
C438 VDD1.n52 B 0.050742f
C439 VDD1.n53 B 0.030487f
C440 VDD1.n54 B 0.022899f
C441 VDD1.n55 B 0.012305f
C442 VDD1.n56 B 0.029085f
C443 VDD1.n57 B 0.013029f
C444 VDD1.n58 B 0.022899f
C445 VDD1.n59 B 0.012667f
C446 VDD1.n60 B 0.029085f
C447 VDD1.n61 B 0.013029f
C448 VDD1.n62 B 0.022899f
C449 VDD1.n63 B 0.012305f
C450 VDD1.n64 B 0.029085f
C451 VDD1.n65 B 0.013029f
C452 VDD1.n66 B 0.022899f
C453 VDD1.n67 B 0.012305f
C454 VDD1.n68 B 0.021813f
C455 VDD1.n69 B 0.020561f
C456 VDD1.t4 B 0.048873f
C457 VDD1.n70 B 0.147257f
C458 VDD1.n71 B 0.948459f
C459 VDD1.n72 B 0.012305f
C460 VDD1.n73 B 0.013029f
C461 VDD1.n74 B 0.029085f
C462 VDD1.n75 B 0.029085f
C463 VDD1.n76 B 0.013029f
C464 VDD1.n77 B 0.012305f
C465 VDD1.n78 B 0.022899f
C466 VDD1.n79 B 0.022899f
C467 VDD1.n80 B 0.012305f
C468 VDD1.n81 B 0.013029f
C469 VDD1.n82 B 0.029085f
C470 VDD1.n83 B 0.029085f
C471 VDD1.n84 B 0.013029f
C472 VDD1.n85 B 0.012305f
C473 VDD1.n86 B 0.022899f
C474 VDD1.n87 B 0.022899f
C475 VDD1.n88 B 0.012305f
C476 VDD1.n89 B 0.012305f
C477 VDD1.n90 B 0.013029f
C478 VDD1.n91 B 0.029085f
C479 VDD1.n92 B 0.029085f
C480 VDD1.n93 B 0.029085f
C481 VDD1.n94 B 0.012667f
C482 VDD1.n95 B 0.012305f
C483 VDD1.n96 B 0.022899f
C484 VDD1.n97 B 0.022899f
C485 VDD1.n98 B 0.012305f
C486 VDD1.n99 B 0.013029f
C487 VDD1.n100 B 0.029085f
C488 VDD1.n101 B 0.059958f
C489 VDD1.n102 B 0.013029f
C490 VDD1.n103 B 0.012305f
C491 VDD1.n104 B 0.053243f
C492 VDD1.n105 B 0.050403f
C493 VDD1.t5 B 0.180413f
C494 VDD1.t2 B 0.180413f
C495 VDD1.n106 B 1.58924f
C496 VDD1.n107 B 1.70732f
C497 VDD1.t1 B 0.180413f
C498 VDD1.t3 B 0.180413f
C499 VDD1.n108 B 1.58835f
C500 VDD1.n109 B 1.95057f
C501 VP.n0 B 0.058727f
C502 VP.t4 B 0.986512f
C503 VP.t3 B 1.04247f
C504 VP.n1 B 0.432917f
C505 VP.n2 B 0.19397f
C506 VP.t5 B 1.04247f
C507 VP.t0 B 0.986512f
C508 VP.t1 B 1.06123f
C509 VP.n3 B 0.430445f
C510 VP.n4 B 0.419044f
C511 VP.n5 B 0.053756f
C512 VP.n6 B 0.432917f
C513 VP.n7 B 1.71003f
C514 VP.n8 B 1.74928f
C515 VP.n9 B 0.058727f
C516 VP.n10 B 0.053756f
C517 VP.n11 B 0.380708f
C518 VP.n12 B 0.053756f
C519 VP.t2 B 1.04247f
C520 VP.n13 B 0.432917f
C521 VP.n14 B 0.041218f
.ends

