* NGSPICE file created from diff_pair_sample_0640.ext - technology: sky130A

.subckt diff_pair_sample_0640 VTAIL VN VP B VDD2 VDD1
X0 B.t19 B.t17 B.t18 B.t11 sky130_fd_pr__nfet_01v8 ad=2.3634 pd=12.9 as=0 ps=0 w=6.06 l=0.24
X1 B.t16 B.t14 B.t15 B.t7 sky130_fd_pr__nfet_01v8 ad=2.3634 pd=12.9 as=0 ps=0 w=6.06 l=0.24
X2 VTAIL.t9 VP.t0 VDD1.t0 B.t4 sky130_fd_pr__nfet_01v8 ad=0.9999 pd=6.39 as=0.9999 ps=6.39 w=6.06 l=0.24
X3 B.t13 B.t10 B.t12 B.t11 sky130_fd_pr__nfet_01v8 ad=2.3634 pd=12.9 as=0 ps=0 w=6.06 l=0.24
X4 VTAIL.t10 VN.t0 VDD2.t5 B.t0 sky130_fd_pr__nfet_01v8 ad=0.9999 pd=6.39 as=0.9999 ps=6.39 w=6.06 l=0.24
X5 VTAIL.t8 VP.t1 VDD1.t2 B.t0 sky130_fd_pr__nfet_01v8 ad=0.9999 pd=6.39 as=0.9999 ps=6.39 w=6.06 l=0.24
X6 VDD1.t1 VP.t2 VTAIL.t7 B.t3 sky130_fd_pr__nfet_01v8 ad=2.3634 pd=12.9 as=0.9999 ps=6.39 w=6.06 l=0.24
X7 VDD1.t5 VP.t3 VTAIL.t6 B.t2 sky130_fd_pr__nfet_01v8 ad=0.9999 pd=6.39 as=2.3634 ps=12.9 w=6.06 l=0.24
X8 VDD2.t4 VN.t1 VTAIL.t11 B.t1 sky130_fd_pr__nfet_01v8 ad=2.3634 pd=12.9 as=0.9999 ps=6.39 w=6.06 l=0.24
X9 VDD2.t3 VN.t2 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=0.9999 pd=6.39 as=2.3634 ps=12.9 w=6.06 l=0.24
X10 VDD2.t2 VN.t3 VTAIL.t1 B.t5 sky130_fd_pr__nfet_01v8 ad=0.9999 pd=6.39 as=2.3634 ps=12.9 w=6.06 l=0.24
X11 VDD1.t4 VP.t4 VTAIL.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=0.9999 pd=6.39 as=2.3634 ps=12.9 w=6.06 l=0.24
X12 VTAIL.t3 VN.t4 VDD2.t1 B.t4 sky130_fd_pr__nfet_01v8 ad=0.9999 pd=6.39 as=0.9999 ps=6.39 w=6.06 l=0.24
X13 B.t9 B.t6 B.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=2.3634 pd=12.9 as=0 ps=0 w=6.06 l=0.24
X14 VDD1.t3 VP.t5 VTAIL.t4 B.t1 sky130_fd_pr__nfet_01v8 ad=2.3634 pd=12.9 as=0.9999 ps=6.39 w=6.06 l=0.24
X15 VDD2.t0 VN.t5 VTAIL.t0 B.t3 sky130_fd_pr__nfet_01v8 ad=2.3634 pd=12.9 as=0.9999 ps=6.39 w=6.06 l=0.24
R0 B.n236 B.t14 834.833
R1 B.n234 B.t6 834.833
R2 B.n65 B.t10 834.833
R3 B.n62 B.t17 834.833
R4 B.n420 B.n419 585
R5 B.n176 B.n60 585
R6 B.n175 B.n174 585
R7 B.n173 B.n172 585
R8 B.n171 B.n170 585
R9 B.n169 B.n168 585
R10 B.n167 B.n166 585
R11 B.n165 B.n164 585
R12 B.n163 B.n162 585
R13 B.n161 B.n160 585
R14 B.n159 B.n158 585
R15 B.n157 B.n156 585
R16 B.n155 B.n154 585
R17 B.n153 B.n152 585
R18 B.n151 B.n150 585
R19 B.n149 B.n148 585
R20 B.n147 B.n146 585
R21 B.n145 B.n144 585
R22 B.n143 B.n142 585
R23 B.n141 B.n140 585
R24 B.n139 B.n138 585
R25 B.n137 B.n136 585
R26 B.n135 B.n134 585
R27 B.n133 B.n132 585
R28 B.n131 B.n130 585
R29 B.n129 B.n128 585
R30 B.n127 B.n126 585
R31 B.n125 B.n124 585
R32 B.n123 B.n122 585
R33 B.n121 B.n120 585
R34 B.n119 B.n118 585
R35 B.n117 B.n116 585
R36 B.n115 B.n114 585
R37 B.n113 B.n112 585
R38 B.n111 B.n110 585
R39 B.n109 B.n108 585
R40 B.n107 B.n106 585
R41 B.n105 B.n104 585
R42 B.n103 B.n102 585
R43 B.n101 B.n100 585
R44 B.n99 B.n98 585
R45 B.n97 B.n96 585
R46 B.n95 B.n94 585
R47 B.n93 B.n92 585
R48 B.n91 B.n90 585
R49 B.n89 B.n88 585
R50 B.n87 B.n86 585
R51 B.n85 B.n84 585
R52 B.n83 B.n82 585
R53 B.n81 B.n80 585
R54 B.n79 B.n78 585
R55 B.n77 B.n76 585
R56 B.n75 B.n74 585
R57 B.n73 B.n72 585
R58 B.n71 B.n70 585
R59 B.n69 B.n68 585
R60 B.n32 B.n31 585
R61 B.n425 B.n424 585
R62 B.n418 B.n61 585
R63 B.n61 B.n29 585
R64 B.n417 B.n28 585
R65 B.n429 B.n28 585
R66 B.n416 B.n27 585
R67 B.n430 B.n27 585
R68 B.n415 B.n26 585
R69 B.n431 B.n26 585
R70 B.n414 B.n413 585
R71 B.n413 B.n25 585
R72 B.n412 B.n21 585
R73 B.n437 B.n21 585
R74 B.n411 B.n20 585
R75 B.n438 B.n20 585
R76 B.n410 B.n19 585
R77 B.n439 B.n19 585
R78 B.n409 B.n408 585
R79 B.n408 B.n15 585
R80 B.n407 B.n14 585
R81 B.n445 B.n14 585
R82 B.n406 B.n13 585
R83 B.n446 B.n13 585
R84 B.n405 B.n12 585
R85 B.n447 B.n12 585
R86 B.n404 B.n403 585
R87 B.n403 B.n11 585
R88 B.n402 B.n7 585
R89 B.n453 B.n7 585
R90 B.n401 B.n6 585
R91 B.n454 B.n6 585
R92 B.n400 B.n5 585
R93 B.n455 B.n5 585
R94 B.n399 B.n398 585
R95 B.n398 B.n4 585
R96 B.n397 B.n177 585
R97 B.n397 B.n396 585
R98 B.n386 B.n178 585
R99 B.n389 B.n178 585
R100 B.n388 B.n387 585
R101 B.n390 B.n388 585
R102 B.n385 B.n182 585
R103 B.n186 B.n182 585
R104 B.n384 B.n383 585
R105 B.n383 B.n382 585
R106 B.n184 B.n183 585
R107 B.n185 B.n184 585
R108 B.n375 B.n374 585
R109 B.n376 B.n375 585
R110 B.n373 B.n191 585
R111 B.n191 B.n190 585
R112 B.n372 B.n371 585
R113 B.n371 B.n370 585
R114 B.n193 B.n192 585
R115 B.n363 B.n193 585
R116 B.n362 B.n361 585
R117 B.n364 B.n362 585
R118 B.n360 B.n198 585
R119 B.n198 B.n197 585
R120 B.n359 B.n358 585
R121 B.n358 B.n357 585
R122 B.n200 B.n199 585
R123 B.n201 B.n200 585
R124 B.n353 B.n352 585
R125 B.n204 B.n203 585
R126 B.n349 B.n348 585
R127 B.n350 B.n349 585
R128 B.n347 B.n233 585
R129 B.n346 B.n345 585
R130 B.n344 B.n343 585
R131 B.n342 B.n341 585
R132 B.n340 B.n339 585
R133 B.n338 B.n337 585
R134 B.n336 B.n335 585
R135 B.n334 B.n333 585
R136 B.n332 B.n331 585
R137 B.n330 B.n329 585
R138 B.n328 B.n327 585
R139 B.n326 B.n325 585
R140 B.n324 B.n323 585
R141 B.n322 B.n321 585
R142 B.n320 B.n319 585
R143 B.n318 B.n317 585
R144 B.n316 B.n315 585
R145 B.n314 B.n313 585
R146 B.n312 B.n311 585
R147 B.n310 B.n309 585
R148 B.n308 B.n307 585
R149 B.n305 B.n304 585
R150 B.n303 B.n302 585
R151 B.n301 B.n300 585
R152 B.n299 B.n298 585
R153 B.n297 B.n296 585
R154 B.n295 B.n294 585
R155 B.n293 B.n292 585
R156 B.n291 B.n290 585
R157 B.n289 B.n288 585
R158 B.n287 B.n286 585
R159 B.n284 B.n283 585
R160 B.n282 B.n281 585
R161 B.n280 B.n279 585
R162 B.n278 B.n277 585
R163 B.n276 B.n275 585
R164 B.n274 B.n273 585
R165 B.n272 B.n271 585
R166 B.n270 B.n269 585
R167 B.n268 B.n267 585
R168 B.n266 B.n265 585
R169 B.n264 B.n263 585
R170 B.n262 B.n261 585
R171 B.n260 B.n259 585
R172 B.n258 B.n257 585
R173 B.n256 B.n255 585
R174 B.n254 B.n253 585
R175 B.n252 B.n251 585
R176 B.n250 B.n249 585
R177 B.n248 B.n247 585
R178 B.n246 B.n245 585
R179 B.n244 B.n243 585
R180 B.n242 B.n241 585
R181 B.n240 B.n239 585
R182 B.n238 B.n232 585
R183 B.n350 B.n232 585
R184 B.n354 B.n202 585
R185 B.n202 B.n201 585
R186 B.n356 B.n355 585
R187 B.n357 B.n356 585
R188 B.n196 B.n195 585
R189 B.n197 B.n196 585
R190 B.n366 B.n365 585
R191 B.n365 B.n364 585
R192 B.n367 B.n194 585
R193 B.n363 B.n194 585
R194 B.n369 B.n368 585
R195 B.n370 B.n369 585
R196 B.n189 B.n188 585
R197 B.n190 B.n189 585
R198 B.n378 B.n377 585
R199 B.n377 B.n376 585
R200 B.n379 B.n187 585
R201 B.n187 B.n185 585
R202 B.n381 B.n380 585
R203 B.n382 B.n381 585
R204 B.n181 B.n180 585
R205 B.n186 B.n181 585
R206 B.n392 B.n391 585
R207 B.n391 B.n390 585
R208 B.n393 B.n179 585
R209 B.n389 B.n179 585
R210 B.n395 B.n394 585
R211 B.n396 B.n395 585
R212 B.n2 B.n0 585
R213 B.n4 B.n2 585
R214 B.n3 B.n1 585
R215 B.n454 B.n3 585
R216 B.n452 B.n451 585
R217 B.n453 B.n452 585
R218 B.n450 B.n8 585
R219 B.n11 B.n8 585
R220 B.n449 B.n448 585
R221 B.n448 B.n447 585
R222 B.n10 B.n9 585
R223 B.n446 B.n10 585
R224 B.n444 B.n443 585
R225 B.n445 B.n444 585
R226 B.n442 B.n16 585
R227 B.n16 B.n15 585
R228 B.n441 B.n440 585
R229 B.n440 B.n439 585
R230 B.n18 B.n17 585
R231 B.n438 B.n18 585
R232 B.n436 B.n435 585
R233 B.n437 B.n436 585
R234 B.n434 B.n22 585
R235 B.n25 B.n22 585
R236 B.n433 B.n432 585
R237 B.n432 B.n431 585
R238 B.n24 B.n23 585
R239 B.n430 B.n24 585
R240 B.n428 B.n427 585
R241 B.n429 B.n428 585
R242 B.n426 B.n30 585
R243 B.n30 B.n29 585
R244 B.n457 B.n456 585
R245 B.n456 B.n455 585
R246 B.n352 B.n202 458.866
R247 B.n424 B.n30 458.866
R248 B.n232 B.n200 458.866
R249 B.n420 B.n61 458.866
R250 B.n422 B.n421 256.663
R251 B.n422 B.n59 256.663
R252 B.n422 B.n58 256.663
R253 B.n422 B.n57 256.663
R254 B.n422 B.n56 256.663
R255 B.n422 B.n55 256.663
R256 B.n422 B.n54 256.663
R257 B.n422 B.n53 256.663
R258 B.n422 B.n52 256.663
R259 B.n422 B.n51 256.663
R260 B.n422 B.n50 256.663
R261 B.n422 B.n49 256.663
R262 B.n422 B.n48 256.663
R263 B.n422 B.n47 256.663
R264 B.n422 B.n46 256.663
R265 B.n422 B.n45 256.663
R266 B.n422 B.n44 256.663
R267 B.n422 B.n43 256.663
R268 B.n422 B.n42 256.663
R269 B.n422 B.n41 256.663
R270 B.n422 B.n40 256.663
R271 B.n422 B.n39 256.663
R272 B.n422 B.n38 256.663
R273 B.n422 B.n37 256.663
R274 B.n422 B.n36 256.663
R275 B.n422 B.n35 256.663
R276 B.n422 B.n34 256.663
R277 B.n422 B.n33 256.663
R278 B.n423 B.n422 256.663
R279 B.n351 B.n350 256.663
R280 B.n350 B.n205 256.663
R281 B.n350 B.n206 256.663
R282 B.n350 B.n207 256.663
R283 B.n350 B.n208 256.663
R284 B.n350 B.n209 256.663
R285 B.n350 B.n210 256.663
R286 B.n350 B.n211 256.663
R287 B.n350 B.n212 256.663
R288 B.n350 B.n213 256.663
R289 B.n350 B.n214 256.663
R290 B.n350 B.n215 256.663
R291 B.n350 B.n216 256.663
R292 B.n350 B.n217 256.663
R293 B.n350 B.n218 256.663
R294 B.n350 B.n219 256.663
R295 B.n350 B.n220 256.663
R296 B.n350 B.n221 256.663
R297 B.n350 B.n222 256.663
R298 B.n350 B.n223 256.663
R299 B.n350 B.n224 256.663
R300 B.n350 B.n225 256.663
R301 B.n350 B.n226 256.663
R302 B.n350 B.n227 256.663
R303 B.n350 B.n228 256.663
R304 B.n350 B.n229 256.663
R305 B.n350 B.n230 256.663
R306 B.n350 B.n231 256.663
R307 B.n236 B.t16 191.204
R308 B.n62 B.t18 191.204
R309 B.n234 B.t9 191.204
R310 B.n65 B.t12 191.204
R311 B.n237 B.t15 180.15
R312 B.n63 B.t19 180.15
R313 B.n235 B.t8 180.15
R314 B.n66 B.t13 180.15
R315 B.n356 B.n202 163.367
R316 B.n356 B.n196 163.367
R317 B.n365 B.n196 163.367
R318 B.n365 B.n194 163.367
R319 B.n369 B.n194 163.367
R320 B.n369 B.n189 163.367
R321 B.n377 B.n189 163.367
R322 B.n377 B.n187 163.367
R323 B.n381 B.n187 163.367
R324 B.n381 B.n181 163.367
R325 B.n391 B.n181 163.367
R326 B.n391 B.n179 163.367
R327 B.n395 B.n179 163.367
R328 B.n395 B.n2 163.367
R329 B.n456 B.n2 163.367
R330 B.n456 B.n3 163.367
R331 B.n452 B.n3 163.367
R332 B.n452 B.n8 163.367
R333 B.n448 B.n8 163.367
R334 B.n448 B.n10 163.367
R335 B.n444 B.n10 163.367
R336 B.n444 B.n16 163.367
R337 B.n440 B.n16 163.367
R338 B.n440 B.n18 163.367
R339 B.n436 B.n18 163.367
R340 B.n436 B.n22 163.367
R341 B.n432 B.n22 163.367
R342 B.n432 B.n24 163.367
R343 B.n428 B.n24 163.367
R344 B.n428 B.n30 163.367
R345 B.n349 B.n204 163.367
R346 B.n349 B.n233 163.367
R347 B.n345 B.n344 163.367
R348 B.n341 B.n340 163.367
R349 B.n337 B.n336 163.367
R350 B.n333 B.n332 163.367
R351 B.n329 B.n328 163.367
R352 B.n325 B.n324 163.367
R353 B.n321 B.n320 163.367
R354 B.n317 B.n316 163.367
R355 B.n313 B.n312 163.367
R356 B.n309 B.n308 163.367
R357 B.n304 B.n303 163.367
R358 B.n300 B.n299 163.367
R359 B.n296 B.n295 163.367
R360 B.n292 B.n291 163.367
R361 B.n288 B.n287 163.367
R362 B.n283 B.n282 163.367
R363 B.n279 B.n278 163.367
R364 B.n275 B.n274 163.367
R365 B.n271 B.n270 163.367
R366 B.n267 B.n266 163.367
R367 B.n263 B.n262 163.367
R368 B.n259 B.n258 163.367
R369 B.n255 B.n254 163.367
R370 B.n251 B.n250 163.367
R371 B.n247 B.n246 163.367
R372 B.n243 B.n242 163.367
R373 B.n239 B.n232 163.367
R374 B.n358 B.n200 163.367
R375 B.n358 B.n198 163.367
R376 B.n362 B.n198 163.367
R377 B.n362 B.n193 163.367
R378 B.n371 B.n193 163.367
R379 B.n371 B.n191 163.367
R380 B.n375 B.n191 163.367
R381 B.n375 B.n184 163.367
R382 B.n383 B.n184 163.367
R383 B.n383 B.n182 163.367
R384 B.n388 B.n182 163.367
R385 B.n388 B.n178 163.367
R386 B.n397 B.n178 163.367
R387 B.n398 B.n397 163.367
R388 B.n398 B.n5 163.367
R389 B.n6 B.n5 163.367
R390 B.n7 B.n6 163.367
R391 B.n403 B.n7 163.367
R392 B.n403 B.n12 163.367
R393 B.n13 B.n12 163.367
R394 B.n14 B.n13 163.367
R395 B.n408 B.n14 163.367
R396 B.n408 B.n19 163.367
R397 B.n20 B.n19 163.367
R398 B.n21 B.n20 163.367
R399 B.n413 B.n21 163.367
R400 B.n413 B.n26 163.367
R401 B.n27 B.n26 163.367
R402 B.n28 B.n27 163.367
R403 B.n61 B.n28 163.367
R404 B.n68 B.n32 163.367
R405 B.n72 B.n71 163.367
R406 B.n76 B.n75 163.367
R407 B.n80 B.n79 163.367
R408 B.n84 B.n83 163.367
R409 B.n88 B.n87 163.367
R410 B.n92 B.n91 163.367
R411 B.n96 B.n95 163.367
R412 B.n100 B.n99 163.367
R413 B.n104 B.n103 163.367
R414 B.n108 B.n107 163.367
R415 B.n112 B.n111 163.367
R416 B.n116 B.n115 163.367
R417 B.n120 B.n119 163.367
R418 B.n124 B.n123 163.367
R419 B.n128 B.n127 163.367
R420 B.n132 B.n131 163.367
R421 B.n136 B.n135 163.367
R422 B.n140 B.n139 163.367
R423 B.n144 B.n143 163.367
R424 B.n148 B.n147 163.367
R425 B.n152 B.n151 163.367
R426 B.n156 B.n155 163.367
R427 B.n160 B.n159 163.367
R428 B.n164 B.n163 163.367
R429 B.n168 B.n167 163.367
R430 B.n172 B.n171 163.367
R431 B.n174 B.n60 163.367
R432 B.n350 B.n201 107.719
R433 B.n422 B.n29 107.719
R434 B.n352 B.n351 71.676
R435 B.n233 B.n205 71.676
R436 B.n344 B.n206 71.676
R437 B.n340 B.n207 71.676
R438 B.n336 B.n208 71.676
R439 B.n332 B.n209 71.676
R440 B.n328 B.n210 71.676
R441 B.n324 B.n211 71.676
R442 B.n320 B.n212 71.676
R443 B.n316 B.n213 71.676
R444 B.n312 B.n214 71.676
R445 B.n308 B.n215 71.676
R446 B.n303 B.n216 71.676
R447 B.n299 B.n217 71.676
R448 B.n295 B.n218 71.676
R449 B.n291 B.n219 71.676
R450 B.n287 B.n220 71.676
R451 B.n282 B.n221 71.676
R452 B.n278 B.n222 71.676
R453 B.n274 B.n223 71.676
R454 B.n270 B.n224 71.676
R455 B.n266 B.n225 71.676
R456 B.n262 B.n226 71.676
R457 B.n258 B.n227 71.676
R458 B.n254 B.n228 71.676
R459 B.n250 B.n229 71.676
R460 B.n246 B.n230 71.676
R461 B.n242 B.n231 71.676
R462 B.n424 B.n423 71.676
R463 B.n68 B.n33 71.676
R464 B.n72 B.n34 71.676
R465 B.n76 B.n35 71.676
R466 B.n80 B.n36 71.676
R467 B.n84 B.n37 71.676
R468 B.n88 B.n38 71.676
R469 B.n92 B.n39 71.676
R470 B.n96 B.n40 71.676
R471 B.n100 B.n41 71.676
R472 B.n104 B.n42 71.676
R473 B.n108 B.n43 71.676
R474 B.n112 B.n44 71.676
R475 B.n116 B.n45 71.676
R476 B.n120 B.n46 71.676
R477 B.n124 B.n47 71.676
R478 B.n128 B.n48 71.676
R479 B.n132 B.n49 71.676
R480 B.n136 B.n50 71.676
R481 B.n140 B.n51 71.676
R482 B.n144 B.n52 71.676
R483 B.n148 B.n53 71.676
R484 B.n152 B.n54 71.676
R485 B.n156 B.n55 71.676
R486 B.n160 B.n56 71.676
R487 B.n164 B.n57 71.676
R488 B.n168 B.n58 71.676
R489 B.n172 B.n59 71.676
R490 B.n421 B.n60 71.676
R491 B.n421 B.n420 71.676
R492 B.n174 B.n59 71.676
R493 B.n171 B.n58 71.676
R494 B.n167 B.n57 71.676
R495 B.n163 B.n56 71.676
R496 B.n159 B.n55 71.676
R497 B.n155 B.n54 71.676
R498 B.n151 B.n53 71.676
R499 B.n147 B.n52 71.676
R500 B.n143 B.n51 71.676
R501 B.n139 B.n50 71.676
R502 B.n135 B.n49 71.676
R503 B.n131 B.n48 71.676
R504 B.n127 B.n47 71.676
R505 B.n123 B.n46 71.676
R506 B.n119 B.n45 71.676
R507 B.n115 B.n44 71.676
R508 B.n111 B.n43 71.676
R509 B.n107 B.n42 71.676
R510 B.n103 B.n41 71.676
R511 B.n99 B.n40 71.676
R512 B.n95 B.n39 71.676
R513 B.n91 B.n38 71.676
R514 B.n87 B.n37 71.676
R515 B.n83 B.n36 71.676
R516 B.n79 B.n35 71.676
R517 B.n75 B.n34 71.676
R518 B.n71 B.n33 71.676
R519 B.n423 B.n32 71.676
R520 B.n351 B.n204 71.676
R521 B.n345 B.n205 71.676
R522 B.n341 B.n206 71.676
R523 B.n337 B.n207 71.676
R524 B.n333 B.n208 71.676
R525 B.n329 B.n209 71.676
R526 B.n325 B.n210 71.676
R527 B.n321 B.n211 71.676
R528 B.n317 B.n212 71.676
R529 B.n313 B.n213 71.676
R530 B.n309 B.n214 71.676
R531 B.n304 B.n215 71.676
R532 B.n300 B.n216 71.676
R533 B.n296 B.n217 71.676
R534 B.n292 B.n218 71.676
R535 B.n288 B.n219 71.676
R536 B.n283 B.n220 71.676
R537 B.n279 B.n221 71.676
R538 B.n275 B.n222 71.676
R539 B.n271 B.n223 71.676
R540 B.n267 B.n224 71.676
R541 B.n263 B.n225 71.676
R542 B.n259 B.n226 71.676
R543 B.n255 B.n227 71.676
R544 B.n251 B.n228 71.676
R545 B.n247 B.n229 71.676
R546 B.n243 B.n230 71.676
R547 B.n239 B.n231 71.676
R548 B.n357 B.n201 65.9908
R549 B.n357 B.n197 65.9908
R550 B.n364 B.n197 65.9908
R551 B.n364 B.n363 65.9908
R552 B.n370 B.n190 65.9908
R553 B.n376 B.n190 65.9908
R554 B.n376 B.n185 65.9908
R555 B.n382 B.n185 65.9908
R556 B.n390 B.n389 65.9908
R557 B.n396 B.n4 65.9908
R558 B.n455 B.n4 65.9908
R559 B.n455 B.n454 65.9908
R560 B.n454 B.n453 65.9908
R561 B.n447 B.n11 65.9908
R562 B.n445 B.n15 65.9908
R563 B.n439 B.n15 65.9908
R564 B.n439 B.n438 65.9908
R565 B.n438 B.n437 65.9908
R566 B.n431 B.n25 65.9908
R567 B.n431 B.n430 65.9908
R568 B.n430 B.n429 65.9908
R569 B.n429 B.n29 65.9908
R570 B.n285 B.n237 59.5399
R571 B.n306 B.n235 59.5399
R572 B.n67 B.n66 59.5399
R573 B.n64 B.n63 59.5399
R574 B.n186 B.t4 58.2272
R575 B.t0 B.n446 58.2272
R576 B.t3 B.n186 52.4046
R577 B.n446 B.t2 52.4046
R578 B.n370 B.t7 44.641
R579 B.n437 B.t11 44.641
R580 B.n389 B.t5 36.8774
R581 B.n11 B.t1 36.8774
R582 B.n426 B.n425 29.8151
R583 B.n238 B.n199 29.8151
R584 B.n354 B.n353 29.8151
R585 B.n419 B.n418 29.8151
R586 B.n396 B.t5 29.1139
R587 B.n453 B.t1 29.1139
R588 B.n363 B.t7 21.3503
R589 B.n25 B.t11 21.3503
R590 B B.n457 18.0485
R591 B.n382 B.t3 13.5867
R592 B.t2 B.n445 13.5867
R593 B.n237 B.n236 11.055
R594 B.n235 B.n234 11.055
R595 B.n66 B.n65 11.055
R596 B.n63 B.n62 11.055
R597 B.n425 B.n31 10.6151
R598 B.n69 B.n31 10.6151
R599 B.n70 B.n69 10.6151
R600 B.n73 B.n70 10.6151
R601 B.n74 B.n73 10.6151
R602 B.n77 B.n74 10.6151
R603 B.n78 B.n77 10.6151
R604 B.n81 B.n78 10.6151
R605 B.n82 B.n81 10.6151
R606 B.n85 B.n82 10.6151
R607 B.n86 B.n85 10.6151
R608 B.n89 B.n86 10.6151
R609 B.n90 B.n89 10.6151
R610 B.n93 B.n90 10.6151
R611 B.n94 B.n93 10.6151
R612 B.n97 B.n94 10.6151
R613 B.n98 B.n97 10.6151
R614 B.n101 B.n98 10.6151
R615 B.n102 B.n101 10.6151
R616 B.n105 B.n102 10.6151
R617 B.n106 B.n105 10.6151
R618 B.n109 B.n106 10.6151
R619 B.n110 B.n109 10.6151
R620 B.n114 B.n113 10.6151
R621 B.n117 B.n114 10.6151
R622 B.n118 B.n117 10.6151
R623 B.n121 B.n118 10.6151
R624 B.n122 B.n121 10.6151
R625 B.n125 B.n122 10.6151
R626 B.n126 B.n125 10.6151
R627 B.n129 B.n126 10.6151
R628 B.n130 B.n129 10.6151
R629 B.n134 B.n133 10.6151
R630 B.n137 B.n134 10.6151
R631 B.n138 B.n137 10.6151
R632 B.n141 B.n138 10.6151
R633 B.n142 B.n141 10.6151
R634 B.n145 B.n142 10.6151
R635 B.n146 B.n145 10.6151
R636 B.n149 B.n146 10.6151
R637 B.n150 B.n149 10.6151
R638 B.n153 B.n150 10.6151
R639 B.n154 B.n153 10.6151
R640 B.n157 B.n154 10.6151
R641 B.n158 B.n157 10.6151
R642 B.n161 B.n158 10.6151
R643 B.n162 B.n161 10.6151
R644 B.n165 B.n162 10.6151
R645 B.n166 B.n165 10.6151
R646 B.n169 B.n166 10.6151
R647 B.n170 B.n169 10.6151
R648 B.n173 B.n170 10.6151
R649 B.n175 B.n173 10.6151
R650 B.n176 B.n175 10.6151
R651 B.n419 B.n176 10.6151
R652 B.n359 B.n199 10.6151
R653 B.n360 B.n359 10.6151
R654 B.n361 B.n360 10.6151
R655 B.n361 B.n192 10.6151
R656 B.n372 B.n192 10.6151
R657 B.n373 B.n372 10.6151
R658 B.n374 B.n373 10.6151
R659 B.n374 B.n183 10.6151
R660 B.n384 B.n183 10.6151
R661 B.n385 B.n384 10.6151
R662 B.n387 B.n385 10.6151
R663 B.n387 B.n386 10.6151
R664 B.n386 B.n177 10.6151
R665 B.n399 B.n177 10.6151
R666 B.n400 B.n399 10.6151
R667 B.n401 B.n400 10.6151
R668 B.n402 B.n401 10.6151
R669 B.n404 B.n402 10.6151
R670 B.n405 B.n404 10.6151
R671 B.n406 B.n405 10.6151
R672 B.n407 B.n406 10.6151
R673 B.n409 B.n407 10.6151
R674 B.n410 B.n409 10.6151
R675 B.n411 B.n410 10.6151
R676 B.n412 B.n411 10.6151
R677 B.n414 B.n412 10.6151
R678 B.n415 B.n414 10.6151
R679 B.n416 B.n415 10.6151
R680 B.n417 B.n416 10.6151
R681 B.n418 B.n417 10.6151
R682 B.n353 B.n203 10.6151
R683 B.n348 B.n203 10.6151
R684 B.n348 B.n347 10.6151
R685 B.n347 B.n346 10.6151
R686 B.n346 B.n343 10.6151
R687 B.n343 B.n342 10.6151
R688 B.n342 B.n339 10.6151
R689 B.n339 B.n338 10.6151
R690 B.n338 B.n335 10.6151
R691 B.n335 B.n334 10.6151
R692 B.n334 B.n331 10.6151
R693 B.n331 B.n330 10.6151
R694 B.n330 B.n327 10.6151
R695 B.n327 B.n326 10.6151
R696 B.n326 B.n323 10.6151
R697 B.n323 B.n322 10.6151
R698 B.n322 B.n319 10.6151
R699 B.n319 B.n318 10.6151
R700 B.n318 B.n315 10.6151
R701 B.n315 B.n314 10.6151
R702 B.n314 B.n311 10.6151
R703 B.n311 B.n310 10.6151
R704 B.n310 B.n307 10.6151
R705 B.n305 B.n302 10.6151
R706 B.n302 B.n301 10.6151
R707 B.n301 B.n298 10.6151
R708 B.n298 B.n297 10.6151
R709 B.n297 B.n294 10.6151
R710 B.n294 B.n293 10.6151
R711 B.n293 B.n290 10.6151
R712 B.n290 B.n289 10.6151
R713 B.n289 B.n286 10.6151
R714 B.n284 B.n281 10.6151
R715 B.n281 B.n280 10.6151
R716 B.n280 B.n277 10.6151
R717 B.n277 B.n276 10.6151
R718 B.n276 B.n273 10.6151
R719 B.n273 B.n272 10.6151
R720 B.n272 B.n269 10.6151
R721 B.n269 B.n268 10.6151
R722 B.n268 B.n265 10.6151
R723 B.n265 B.n264 10.6151
R724 B.n264 B.n261 10.6151
R725 B.n261 B.n260 10.6151
R726 B.n260 B.n257 10.6151
R727 B.n257 B.n256 10.6151
R728 B.n256 B.n253 10.6151
R729 B.n253 B.n252 10.6151
R730 B.n252 B.n249 10.6151
R731 B.n249 B.n248 10.6151
R732 B.n248 B.n245 10.6151
R733 B.n245 B.n244 10.6151
R734 B.n244 B.n241 10.6151
R735 B.n241 B.n240 10.6151
R736 B.n240 B.n238 10.6151
R737 B.n355 B.n354 10.6151
R738 B.n355 B.n195 10.6151
R739 B.n366 B.n195 10.6151
R740 B.n367 B.n366 10.6151
R741 B.n368 B.n367 10.6151
R742 B.n368 B.n188 10.6151
R743 B.n378 B.n188 10.6151
R744 B.n379 B.n378 10.6151
R745 B.n380 B.n379 10.6151
R746 B.n380 B.n180 10.6151
R747 B.n392 B.n180 10.6151
R748 B.n393 B.n392 10.6151
R749 B.n394 B.n393 10.6151
R750 B.n394 B.n0 10.6151
R751 B.n451 B.n1 10.6151
R752 B.n451 B.n450 10.6151
R753 B.n450 B.n449 10.6151
R754 B.n449 B.n9 10.6151
R755 B.n443 B.n9 10.6151
R756 B.n443 B.n442 10.6151
R757 B.n442 B.n441 10.6151
R758 B.n441 B.n17 10.6151
R759 B.n435 B.n17 10.6151
R760 B.n435 B.n434 10.6151
R761 B.n434 B.n433 10.6151
R762 B.n433 B.n23 10.6151
R763 B.n427 B.n23 10.6151
R764 B.n427 B.n426 10.6151
R765 B.n110 B.n67 9.36635
R766 B.n133 B.n64 9.36635
R767 B.n307 B.n306 9.36635
R768 B.n285 B.n284 9.36635
R769 B.n390 B.t4 7.76406
R770 B.n447 B.t0 7.76406
R771 B.n457 B.n0 2.81026
R772 B.n457 B.n1 2.81026
R773 B.n113 B.n67 1.24928
R774 B.n130 B.n64 1.24928
R775 B.n306 B.n305 1.24928
R776 B.n286 B.n285 1.24928
R777 VP.n7 VP.t4 785.807
R778 VP.n5 VP.t2 785.807
R779 VP.n0 VP.t5 785.807
R780 VP.n2 VP.t3 785.807
R781 VP.n6 VP.t0 739.067
R782 VP.n1 VP.t1 739.067
R783 VP.n3 VP.n0 161.489
R784 VP.n8 VP.n7 161.3
R785 VP.n3 VP.n2 161.3
R786 VP.n5 VP.n4 161.3
R787 VP.n6 VP.n5 36.5157
R788 VP.n7 VP.n6 36.5157
R789 VP.n1 VP.n0 36.5157
R790 VP.n2 VP.n1 36.5157
R791 VP.n4 VP.n3 35.0043
R792 VP.n8 VP.n4 0.189894
R793 VP VP.n8 0.0516364
R794 VDD1.n26 VDD1.n0 289.615
R795 VDD1.n57 VDD1.n31 289.615
R796 VDD1.n27 VDD1.n26 185
R797 VDD1.n25 VDD1.n24 185
R798 VDD1.n4 VDD1.n3 185
R799 VDD1.n19 VDD1.n18 185
R800 VDD1.n17 VDD1.n16 185
R801 VDD1.n8 VDD1.n7 185
R802 VDD1.n11 VDD1.n10 185
R803 VDD1.n42 VDD1.n41 185
R804 VDD1.n39 VDD1.n38 185
R805 VDD1.n48 VDD1.n47 185
R806 VDD1.n50 VDD1.n49 185
R807 VDD1.n35 VDD1.n34 185
R808 VDD1.n56 VDD1.n55 185
R809 VDD1.n58 VDD1.n57 185
R810 VDD1.t3 VDD1.n9 147.661
R811 VDD1.t1 VDD1.n40 147.661
R812 VDD1.n26 VDD1.n25 104.615
R813 VDD1.n25 VDD1.n3 104.615
R814 VDD1.n18 VDD1.n3 104.615
R815 VDD1.n18 VDD1.n17 104.615
R816 VDD1.n17 VDD1.n7 104.615
R817 VDD1.n10 VDD1.n7 104.615
R818 VDD1.n41 VDD1.n38 104.615
R819 VDD1.n48 VDD1.n38 104.615
R820 VDD1.n49 VDD1.n48 104.615
R821 VDD1.n49 VDD1.n34 104.615
R822 VDD1.n56 VDD1.n34 104.615
R823 VDD1.n57 VDD1.n56 104.615
R824 VDD1.n63 VDD1.n62 68.4218
R825 VDD1.n65 VDD1.n64 68.3543
R826 VDD1.n10 VDD1.t3 52.3082
R827 VDD1.n41 VDD1.t1 52.3082
R828 VDD1 VDD1.n30 50.4545
R829 VDD1.n63 VDD1.n61 50.341
R830 VDD1.n65 VDD1.n63 31.3651
R831 VDD1.n11 VDD1.n9 15.6674
R832 VDD1.n42 VDD1.n40 15.6674
R833 VDD1.n12 VDD1.n8 12.8005
R834 VDD1.n43 VDD1.n39 12.8005
R835 VDD1.n16 VDD1.n15 12.0247
R836 VDD1.n47 VDD1.n46 12.0247
R837 VDD1.n19 VDD1.n6 11.249
R838 VDD1.n50 VDD1.n37 11.249
R839 VDD1.n20 VDD1.n4 10.4732
R840 VDD1.n51 VDD1.n35 10.4732
R841 VDD1.n24 VDD1.n23 9.69747
R842 VDD1.n55 VDD1.n54 9.69747
R843 VDD1.n30 VDD1.n29 9.45567
R844 VDD1.n61 VDD1.n60 9.45567
R845 VDD1.n29 VDD1.n28 9.3005
R846 VDD1.n2 VDD1.n1 9.3005
R847 VDD1.n23 VDD1.n22 9.3005
R848 VDD1.n21 VDD1.n20 9.3005
R849 VDD1.n6 VDD1.n5 9.3005
R850 VDD1.n15 VDD1.n14 9.3005
R851 VDD1.n13 VDD1.n12 9.3005
R852 VDD1.n60 VDD1.n59 9.3005
R853 VDD1.n33 VDD1.n32 9.3005
R854 VDD1.n54 VDD1.n53 9.3005
R855 VDD1.n52 VDD1.n51 9.3005
R856 VDD1.n37 VDD1.n36 9.3005
R857 VDD1.n46 VDD1.n45 9.3005
R858 VDD1.n44 VDD1.n43 9.3005
R859 VDD1.n27 VDD1.n2 8.92171
R860 VDD1.n58 VDD1.n33 8.92171
R861 VDD1.n28 VDD1.n0 8.14595
R862 VDD1.n59 VDD1.n31 8.14595
R863 VDD1.n30 VDD1.n0 5.81868
R864 VDD1.n61 VDD1.n31 5.81868
R865 VDD1.n28 VDD1.n27 5.04292
R866 VDD1.n59 VDD1.n58 5.04292
R867 VDD1.n13 VDD1.n9 4.38594
R868 VDD1.n44 VDD1.n40 4.38594
R869 VDD1.n24 VDD1.n2 4.26717
R870 VDD1.n55 VDD1.n33 4.26717
R871 VDD1.n23 VDD1.n4 3.49141
R872 VDD1.n54 VDD1.n35 3.49141
R873 VDD1.n64 VDD1.t2 3.26783
R874 VDD1.n64 VDD1.t5 3.26783
R875 VDD1.n62 VDD1.t0 3.26783
R876 VDD1.n62 VDD1.t4 3.26783
R877 VDD1.n20 VDD1.n19 2.71565
R878 VDD1.n51 VDD1.n50 2.71565
R879 VDD1.n16 VDD1.n6 1.93989
R880 VDD1.n47 VDD1.n37 1.93989
R881 VDD1.n15 VDD1.n8 1.16414
R882 VDD1.n46 VDD1.n39 1.16414
R883 VDD1.n12 VDD1.n11 0.388379
R884 VDD1.n43 VDD1.n42 0.388379
R885 VDD1.n29 VDD1.n1 0.155672
R886 VDD1.n22 VDD1.n1 0.155672
R887 VDD1.n22 VDD1.n21 0.155672
R888 VDD1.n21 VDD1.n5 0.155672
R889 VDD1.n14 VDD1.n5 0.155672
R890 VDD1.n14 VDD1.n13 0.155672
R891 VDD1.n45 VDD1.n44 0.155672
R892 VDD1.n45 VDD1.n36 0.155672
R893 VDD1.n52 VDD1.n36 0.155672
R894 VDD1.n53 VDD1.n52 0.155672
R895 VDD1.n53 VDD1.n32 0.155672
R896 VDD1.n60 VDD1.n32 0.155672
R897 VDD1 VDD1.n65 0.0651552
R898 VTAIL.n130 VTAIL.n104 289.615
R899 VTAIL.n28 VTAIL.n2 289.615
R900 VTAIL.n98 VTAIL.n72 289.615
R901 VTAIL.n64 VTAIL.n38 289.615
R902 VTAIL.n115 VTAIL.n114 185
R903 VTAIL.n112 VTAIL.n111 185
R904 VTAIL.n121 VTAIL.n120 185
R905 VTAIL.n123 VTAIL.n122 185
R906 VTAIL.n108 VTAIL.n107 185
R907 VTAIL.n129 VTAIL.n128 185
R908 VTAIL.n131 VTAIL.n130 185
R909 VTAIL.n13 VTAIL.n12 185
R910 VTAIL.n10 VTAIL.n9 185
R911 VTAIL.n19 VTAIL.n18 185
R912 VTAIL.n21 VTAIL.n20 185
R913 VTAIL.n6 VTAIL.n5 185
R914 VTAIL.n27 VTAIL.n26 185
R915 VTAIL.n29 VTAIL.n28 185
R916 VTAIL.n99 VTAIL.n98 185
R917 VTAIL.n97 VTAIL.n96 185
R918 VTAIL.n76 VTAIL.n75 185
R919 VTAIL.n91 VTAIL.n90 185
R920 VTAIL.n89 VTAIL.n88 185
R921 VTAIL.n80 VTAIL.n79 185
R922 VTAIL.n83 VTAIL.n82 185
R923 VTAIL.n65 VTAIL.n64 185
R924 VTAIL.n63 VTAIL.n62 185
R925 VTAIL.n42 VTAIL.n41 185
R926 VTAIL.n57 VTAIL.n56 185
R927 VTAIL.n55 VTAIL.n54 185
R928 VTAIL.n46 VTAIL.n45 185
R929 VTAIL.n49 VTAIL.n48 185
R930 VTAIL.t2 VTAIL.n113 147.661
R931 VTAIL.t5 VTAIL.n11 147.661
R932 VTAIL.t6 VTAIL.n81 147.661
R933 VTAIL.t1 VTAIL.n47 147.661
R934 VTAIL.n114 VTAIL.n111 104.615
R935 VTAIL.n121 VTAIL.n111 104.615
R936 VTAIL.n122 VTAIL.n121 104.615
R937 VTAIL.n122 VTAIL.n107 104.615
R938 VTAIL.n129 VTAIL.n107 104.615
R939 VTAIL.n130 VTAIL.n129 104.615
R940 VTAIL.n12 VTAIL.n9 104.615
R941 VTAIL.n19 VTAIL.n9 104.615
R942 VTAIL.n20 VTAIL.n19 104.615
R943 VTAIL.n20 VTAIL.n5 104.615
R944 VTAIL.n27 VTAIL.n5 104.615
R945 VTAIL.n28 VTAIL.n27 104.615
R946 VTAIL.n98 VTAIL.n97 104.615
R947 VTAIL.n97 VTAIL.n75 104.615
R948 VTAIL.n90 VTAIL.n75 104.615
R949 VTAIL.n90 VTAIL.n89 104.615
R950 VTAIL.n89 VTAIL.n79 104.615
R951 VTAIL.n82 VTAIL.n79 104.615
R952 VTAIL.n64 VTAIL.n63 104.615
R953 VTAIL.n63 VTAIL.n41 104.615
R954 VTAIL.n56 VTAIL.n41 104.615
R955 VTAIL.n56 VTAIL.n55 104.615
R956 VTAIL.n55 VTAIL.n45 104.615
R957 VTAIL.n48 VTAIL.n45 104.615
R958 VTAIL.n114 VTAIL.t2 52.3082
R959 VTAIL.n12 VTAIL.t5 52.3082
R960 VTAIL.n82 VTAIL.t6 52.3082
R961 VTAIL.n48 VTAIL.t1 52.3082
R962 VTAIL.n71 VTAIL.n70 51.6757
R963 VTAIL.n37 VTAIL.n36 51.6757
R964 VTAIL.n1 VTAIL.n0 51.6755
R965 VTAIL.n35 VTAIL.n34 51.6755
R966 VTAIL.n135 VTAIL.n134 33.349
R967 VTAIL.n33 VTAIL.n32 33.349
R968 VTAIL.n103 VTAIL.n102 33.349
R969 VTAIL.n69 VTAIL.n68 33.349
R970 VTAIL.n37 VTAIL.n35 18.5738
R971 VTAIL.n135 VTAIL.n103 18.0824
R972 VTAIL.n115 VTAIL.n113 15.6674
R973 VTAIL.n13 VTAIL.n11 15.6674
R974 VTAIL.n83 VTAIL.n81 15.6674
R975 VTAIL.n49 VTAIL.n47 15.6674
R976 VTAIL.n116 VTAIL.n112 12.8005
R977 VTAIL.n14 VTAIL.n10 12.8005
R978 VTAIL.n84 VTAIL.n80 12.8005
R979 VTAIL.n50 VTAIL.n46 12.8005
R980 VTAIL.n120 VTAIL.n119 12.0247
R981 VTAIL.n18 VTAIL.n17 12.0247
R982 VTAIL.n88 VTAIL.n87 12.0247
R983 VTAIL.n54 VTAIL.n53 12.0247
R984 VTAIL.n123 VTAIL.n110 11.249
R985 VTAIL.n21 VTAIL.n8 11.249
R986 VTAIL.n91 VTAIL.n78 11.249
R987 VTAIL.n57 VTAIL.n44 11.249
R988 VTAIL.n124 VTAIL.n108 10.4732
R989 VTAIL.n22 VTAIL.n6 10.4732
R990 VTAIL.n92 VTAIL.n76 10.4732
R991 VTAIL.n58 VTAIL.n42 10.4732
R992 VTAIL.n128 VTAIL.n127 9.69747
R993 VTAIL.n26 VTAIL.n25 9.69747
R994 VTAIL.n96 VTAIL.n95 9.69747
R995 VTAIL.n62 VTAIL.n61 9.69747
R996 VTAIL.n134 VTAIL.n133 9.45567
R997 VTAIL.n32 VTAIL.n31 9.45567
R998 VTAIL.n102 VTAIL.n101 9.45567
R999 VTAIL.n68 VTAIL.n67 9.45567
R1000 VTAIL.n133 VTAIL.n132 9.3005
R1001 VTAIL.n106 VTAIL.n105 9.3005
R1002 VTAIL.n127 VTAIL.n126 9.3005
R1003 VTAIL.n125 VTAIL.n124 9.3005
R1004 VTAIL.n110 VTAIL.n109 9.3005
R1005 VTAIL.n119 VTAIL.n118 9.3005
R1006 VTAIL.n117 VTAIL.n116 9.3005
R1007 VTAIL.n31 VTAIL.n30 9.3005
R1008 VTAIL.n4 VTAIL.n3 9.3005
R1009 VTAIL.n25 VTAIL.n24 9.3005
R1010 VTAIL.n23 VTAIL.n22 9.3005
R1011 VTAIL.n8 VTAIL.n7 9.3005
R1012 VTAIL.n17 VTAIL.n16 9.3005
R1013 VTAIL.n15 VTAIL.n14 9.3005
R1014 VTAIL.n101 VTAIL.n100 9.3005
R1015 VTAIL.n74 VTAIL.n73 9.3005
R1016 VTAIL.n95 VTAIL.n94 9.3005
R1017 VTAIL.n93 VTAIL.n92 9.3005
R1018 VTAIL.n78 VTAIL.n77 9.3005
R1019 VTAIL.n87 VTAIL.n86 9.3005
R1020 VTAIL.n85 VTAIL.n84 9.3005
R1021 VTAIL.n67 VTAIL.n66 9.3005
R1022 VTAIL.n40 VTAIL.n39 9.3005
R1023 VTAIL.n61 VTAIL.n60 9.3005
R1024 VTAIL.n59 VTAIL.n58 9.3005
R1025 VTAIL.n44 VTAIL.n43 9.3005
R1026 VTAIL.n53 VTAIL.n52 9.3005
R1027 VTAIL.n51 VTAIL.n50 9.3005
R1028 VTAIL.n131 VTAIL.n106 8.92171
R1029 VTAIL.n29 VTAIL.n4 8.92171
R1030 VTAIL.n99 VTAIL.n74 8.92171
R1031 VTAIL.n65 VTAIL.n40 8.92171
R1032 VTAIL.n132 VTAIL.n104 8.14595
R1033 VTAIL.n30 VTAIL.n2 8.14595
R1034 VTAIL.n100 VTAIL.n72 8.14595
R1035 VTAIL.n66 VTAIL.n38 8.14595
R1036 VTAIL.n134 VTAIL.n104 5.81868
R1037 VTAIL.n32 VTAIL.n2 5.81868
R1038 VTAIL.n102 VTAIL.n72 5.81868
R1039 VTAIL.n68 VTAIL.n38 5.81868
R1040 VTAIL.n132 VTAIL.n131 5.04292
R1041 VTAIL.n30 VTAIL.n29 5.04292
R1042 VTAIL.n100 VTAIL.n99 5.04292
R1043 VTAIL.n66 VTAIL.n65 5.04292
R1044 VTAIL.n117 VTAIL.n113 4.38594
R1045 VTAIL.n15 VTAIL.n11 4.38594
R1046 VTAIL.n85 VTAIL.n81 4.38594
R1047 VTAIL.n51 VTAIL.n47 4.38594
R1048 VTAIL.n128 VTAIL.n106 4.26717
R1049 VTAIL.n26 VTAIL.n4 4.26717
R1050 VTAIL.n96 VTAIL.n74 4.26717
R1051 VTAIL.n62 VTAIL.n40 4.26717
R1052 VTAIL.n127 VTAIL.n108 3.49141
R1053 VTAIL.n25 VTAIL.n6 3.49141
R1054 VTAIL.n95 VTAIL.n76 3.49141
R1055 VTAIL.n61 VTAIL.n42 3.49141
R1056 VTAIL.n0 VTAIL.t11 3.26783
R1057 VTAIL.n0 VTAIL.t10 3.26783
R1058 VTAIL.n34 VTAIL.t7 3.26783
R1059 VTAIL.n34 VTAIL.t9 3.26783
R1060 VTAIL.n70 VTAIL.t4 3.26783
R1061 VTAIL.n70 VTAIL.t8 3.26783
R1062 VTAIL.n36 VTAIL.t0 3.26783
R1063 VTAIL.n36 VTAIL.t3 3.26783
R1064 VTAIL.n124 VTAIL.n123 2.71565
R1065 VTAIL.n22 VTAIL.n21 2.71565
R1066 VTAIL.n92 VTAIL.n91 2.71565
R1067 VTAIL.n58 VTAIL.n57 2.71565
R1068 VTAIL.n120 VTAIL.n110 1.93989
R1069 VTAIL.n18 VTAIL.n8 1.93989
R1070 VTAIL.n88 VTAIL.n78 1.93989
R1071 VTAIL.n54 VTAIL.n44 1.93989
R1072 VTAIL.n119 VTAIL.n112 1.16414
R1073 VTAIL.n17 VTAIL.n10 1.16414
R1074 VTAIL.n87 VTAIL.n80 1.16414
R1075 VTAIL.n53 VTAIL.n46 1.16414
R1076 VTAIL.n71 VTAIL.n69 0.716017
R1077 VTAIL.n33 VTAIL.n1 0.716017
R1078 VTAIL.n69 VTAIL.n37 0.491879
R1079 VTAIL.n103 VTAIL.n71 0.491879
R1080 VTAIL.n35 VTAIL.n33 0.491879
R1081 VTAIL.n116 VTAIL.n115 0.388379
R1082 VTAIL.n14 VTAIL.n13 0.388379
R1083 VTAIL.n84 VTAIL.n83 0.388379
R1084 VTAIL.n50 VTAIL.n49 0.388379
R1085 VTAIL VTAIL.n135 0.310845
R1086 VTAIL VTAIL.n1 0.181534
R1087 VTAIL.n118 VTAIL.n117 0.155672
R1088 VTAIL.n118 VTAIL.n109 0.155672
R1089 VTAIL.n125 VTAIL.n109 0.155672
R1090 VTAIL.n126 VTAIL.n125 0.155672
R1091 VTAIL.n126 VTAIL.n105 0.155672
R1092 VTAIL.n133 VTAIL.n105 0.155672
R1093 VTAIL.n16 VTAIL.n15 0.155672
R1094 VTAIL.n16 VTAIL.n7 0.155672
R1095 VTAIL.n23 VTAIL.n7 0.155672
R1096 VTAIL.n24 VTAIL.n23 0.155672
R1097 VTAIL.n24 VTAIL.n3 0.155672
R1098 VTAIL.n31 VTAIL.n3 0.155672
R1099 VTAIL.n101 VTAIL.n73 0.155672
R1100 VTAIL.n94 VTAIL.n73 0.155672
R1101 VTAIL.n94 VTAIL.n93 0.155672
R1102 VTAIL.n93 VTAIL.n77 0.155672
R1103 VTAIL.n86 VTAIL.n77 0.155672
R1104 VTAIL.n86 VTAIL.n85 0.155672
R1105 VTAIL.n67 VTAIL.n39 0.155672
R1106 VTAIL.n60 VTAIL.n39 0.155672
R1107 VTAIL.n60 VTAIL.n59 0.155672
R1108 VTAIL.n59 VTAIL.n43 0.155672
R1109 VTAIL.n52 VTAIL.n43 0.155672
R1110 VTAIL.n52 VTAIL.n51 0.155672
R1111 VN.n2 VN.t2 785.807
R1112 VN.n0 VN.t1 785.807
R1113 VN.n6 VN.t5 785.807
R1114 VN.n4 VN.t3 785.807
R1115 VN.n1 VN.t0 739.067
R1116 VN.n5 VN.t4 739.067
R1117 VN.n7 VN.n4 161.489
R1118 VN.n3 VN.n0 161.489
R1119 VN.n3 VN.n2 161.3
R1120 VN.n7 VN.n6 161.3
R1121 VN.n1 VN.n0 36.5157
R1122 VN.n2 VN.n1 36.5157
R1123 VN.n6 VN.n5 36.5157
R1124 VN.n5 VN.n4 36.5157
R1125 VN VN.n7 35.385
R1126 VN VN.n3 0.0516364
R1127 VDD2.n59 VDD2.n33 289.615
R1128 VDD2.n26 VDD2.n0 289.615
R1129 VDD2.n60 VDD2.n59 185
R1130 VDD2.n58 VDD2.n57 185
R1131 VDD2.n37 VDD2.n36 185
R1132 VDD2.n52 VDD2.n51 185
R1133 VDD2.n50 VDD2.n49 185
R1134 VDD2.n41 VDD2.n40 185
R1135 VDD2.n44 VDD2.n43 185
R1136 VDD2.n11 VDD2.n10 185
R1137 VDD2.n8 VDD2.n7 185
R1138 VDD2.n17 VDD2.n16 185
R1139 VDD2.n19 VDD2.n18 185
R1140 VDD2.n4 VDD2.n3 185
R1141 VDD2.n25 VDD2.n24 185
R1142 VDD2.n27 VDD2.n26 185
R1143 VDD2.t0 VDD2.n42 147.661
R1144 VDD2.t4 VDD2.n9 147.661
R1145 VDD2.n59 VDD2.n58 104.615
R1146 VDD2.n58 VDD2.n36 104.615
R1147 VDD2.n51 VDD2.n36 104.615
R1148 VDD2.n51 VDD2.n50 104.615
R1149 VDD2.n50 VDD2.n40 104.615
R1150 VDD2.n43 VDD2.n40 104.615
R1151 VDD2.n10 VDD2.n7 104.615
R1152 VDD2.n17 VDD2.n7 104.615
R1153 VDD2.n18 VDD2.n17 104.615
R1154 VDD2.n18 VDD2.n3 104.615
R1155 VDD2.n25 VDD2.n3 104.615
R1156 VDD2.n26 VDD2.n25 104.615
R1157 VDD2.n32 VDD2.n31 68.4218
R1158 VDD2 VDD2.n65 68.4189
R1159 VDD2.n43 VDD2.t0 52.3082
R1160 VDD2.n10 VDD2.t4 52.3082
R1161 VDD2.n32 VDD2.n30 50.341
R1162 VDD2.n64 VDD2.n63 50.0278
R1163 VDD2.n64 VDD2.n32 30.5364
R1164 VDD2.n44 VDD2.n42 15.6674
R1165 VDD2.n11 VDD2.n9 15.6674
R1166 VDD2.n45 VDD2.n41 12.8005
R1167 VDD2.n12 VDD2.n8 12.8005
R1168 VDD2.n49 VDD2.n48 12.0247
R1169 VDD2.n16 VDD2.n15 12.0247
R1170 VDD2.n52 VDD2.n39 11.249
R1171 VDD2.n19 VDD2.n6 11.249
R1172 VDD2.n53 VDD2.n37 10.4732
R1173 VDD2.n20 VDD2.n4 10.4732
R1174 VDD2.n57 VDD2.n56 9.69747
R1175 VDD2.n24 VDD2.n23 9.69747
R1176 VDD2.n63 VDD2.n62 9.45567
R1177 VDD2.n30 VDD2.n29 9.45567
R1178 VDD2.n62 VDD2.n61 9.3005
R1179 VDD2.n35 VDD2.n34 9.3005
R1180 VDD2.n56 VDD2.n55 9.3005
R1181 VDD2.n54 VDD2.n53 9.3005
R1182 VDD2.n39 VDD2.n38 9.3005
R1183 VDD2.n48 VDD2.n47 9.3005
R1184 VDD2.n46 VDD2.n45 9.3005
R1185 VDD2.n29 VDD2.n28 9.3005
R1186 VDD2.n2 VDD2.n1 9.3005
R1187 VDD2.n23 VDD2.n22 9.3005
R1188 VDD2.n21 VDD2.n20 9.3005
R1189 VDD2.n6 VDD2.n5 9.3005
R1190 VDD2.n15 VDD2.n14 9.3005
R1191 VDD2.n13 VDD2.n12 9.3005
R1192 VDD2.n60 VDD2.n35 8.92171
R1193 VDD2.n27 VDD2.n2 8.92171
R1194 VDD2.n61 VDD2.n33 8.14595
R1195 VDD2.n28 VDD2.n0 8.14595
R1196 VDD2.n63 VDD2.n33 5.81868
R1197 VDD2.n30 VDD2.n0 5.81868
R1198 VDD2.n61 VDD2.n60 5.04292
R1199 VDD2.n28 VDD2.n27 5.04292
R1200 VDD2.n46 VDD2.n42 4.38594
R1201 VDD2.n13 VDD2.n9 4.38594
R1202 VDD2.n57 VDD2.n35 4.26717
R1203 VDD2.n24 VDD2.n2 4.26717
R1204 VDD2.n56 VDD2.n37 3.49141
R1205 VDD2.n23 VDD2.n4 3.49141
R1206 VDD2.n65 VDD2.t1 3.26783
R1207 VDD2.n65 VDD2.t2 3.26783
R1208 VDD2.n31 VDD2.t5 3.26783
R1209 VDD2.n31 VDD2.t3 3.26783
R1210 VDD2.n53 VDD2.n52 2.71565
R1211 VDD2.n20 VDD2.n19 2.71565
R1212 VDD2.n49 VDD2.n39 1.93989
R1213 VDD2.n16 VDD2.n6 1.93989
R1214 VDD2.n48 VDD2.n41 1.16414
R1215 VDD2.n15 VDD2.n8 1.16414
R1216 VDD2 VDD2.n64 0.427224
R1217 VDD2.n45 VDD2.n44 0.388379
R1218 VDD2.n12 VDD2.n11 0.388379
R1219 VDD2.n62 VDD2.n34 0.155672
R1220 VDD2.n55 VDD2.n34 0.155672
R1221 VDD2.n55 VDD2.n54 0.155672
R1222 VDD2.n54 VDD2.n38 0.155672
R1223 VDD2.n47 VDD2.n38 0.155672
R1224 VDD2.n47 VDD2.n46 0.155672
R1225 VDD2.n14 VDD2.n13 0.155672
R1226 VDD2.n14 VDD2.n5 0.155672
R1227 VDD2.n21 VDD2.n5 0.155672
R1228 VDD2.n22 VDD2.n21 0.155672
R1229 VDD2.n22 VDD2.n1 0.155672
R1230 VDD2.n29 VDD2.n1 0.155672
C0 VTAIL VDD2 8.48283f
C1 VN VTAIL 1.15955f
C2 VP VDD1 1.46535f
C3 VDD1 VDD2 0.546935f
C4 VP VDD2 0.257952f
C5 VDD1 VN 0.14766f
C6 VP VN 3.53051f
C7 VN VDD2 1.35774f
C8 VDD1 VTAIL 8.449671f
C9 VP VTAIL 1.174f
C10 VDD2 B 3.041617f
C11 VDD1 B 3.01112f
C12 VTAIL B 3.781095f
C13 VN B 5.04541f
C14 VP B 3.913881f
C15 VDD2.n0 B 0.036146f
C16 VDD2.n1 B 0.024996f
C17 VDD2.n2 B 0.013432f
C18 VDD2.n3 B 0.031748f
C19 VDD2.n4 B 0.014222f
C20 VDD2.n5 B 0.024996f
C21 VDD2.n6 B 0.013432f
C22 VDD2.n7 B 0.031748f
C23 VDD2.n8 B 0.014222f
C24 VDD2.n9 B 0.107381f
C25 VDD2.t4 B 0.051769f
C26 VDD2.n10 B 0.023811f
C27 VDD2.n11 B 0.018753f
C28 VDD2.n12 B 0.013432f
C29 VDD2.n13 B 0.601567f
C30 VDD2.n14 B 0.024996f
C31 VDD2.n15 B 0.013432f
C32 VDD2.n16 B 0.014222f
C33 VDD2.n17 B 0.031748f
C34 VDD2.n18 B 0.031748f
C35 VDD2.n19 B 0.014222f
C36 VDD2.n20 B 0.013432f
C37 VDD2.n21 B 0.024996f
C38 VDD2.n22 B 0.024996f
C39 VDD2.n23 B 0.013432f
C40 VDD2.n24 B 0.014222f
C41 VDD2.n25 B 0.031748f
C42 VDD2.n26 B 0.070518f
C43 VDD2.n27 B 0.014222f
C44 VDD2.n28 B 0.013432f
C45 VDD2.n29 B 0.059826f
C46 VDD2.n30 B 0.057422f
C47 VDD2.t5 B 0.1197f
C48 VDD2.t3 B 0.1197f
C49 VDD2.n31 B 1.00015f
C50 VDD2.n32 B 1.29822f
C51 VDD2.n33 B 0.036146f
C52 VDD2.n34 B 0.024996f
C53 VDD2.n35 B 0.013432f
C54 VDD2.n36 B 0.031748f
C55 VDD2.n37 B 0.014222f
C56 VDD2.n38 B 0.024996f
C57 VDD2.n39 B 0.013432f
C58 VDD2.n40 B 0.031748f
C59 VDD2.n41 B 0.014222f
C60 VDD2.n42 B 0.107381f
C61 VDD2.t0 B 0.051769f
C62 VDD2.n43 B 0.023811f
C63 VDD2.n44 B 0.018753f
C64 VDD2.n45 B 0.013432f
C65 VDD2.n46 B 0.601567f
C66 VDD2.n47 B 0.024996f
C67 VDD2.n48 B 0.013432f
C68 VDD2.n49 B 0.014222f
C69 VDD2.n50 B 0.031748f
C70 VDD2.n51 B 0.031748f
C71 VDD2.n52 B 0.014222f
C72 VDD2.n53 B 0.013432f
C73 VDD2.n54 B 0.024996f
C74 VDD2.n55 B 0.024996f
C75 VDD2.n56 B 0.013432f
C76 VDD2.n57 B 0.014222f
C77 VDD2.n58 B 0.031748f
C78 VDD2.n59 B 0.070518f
C79 VDD2.n60 B 0.014222f
C80 VDD2.n61 B 0.013432f
C81 VDD2.n62 B 0.059826f
C82 VDD2.n63 B 0.056947f
C83 VDD2.n64 B 1.44579f
C84 VDD2.t1 B 0.1197f
C85 VDD2.t2 B 0.1197f
C86 VDD2.n65 B 1.00013f
C87 VN.t1 B 0.145148f
C88 VN.n0 B 0.076732f
C89 VN.t0 B 0.141106f
C90 VN.n1 B 0.066697f
C91 VN.t2 B 0.145148f
C92 VN.n2 B 0.076683f
C93 VN.n3 B 0.068381f
C94 VN.t3 B 0.145148f
C95 VN.n4 B 0.076732f
C96 VN.t5 B 0.145148f
C97 VN.t4 B 0.141106f
C98 VN.n5 B 0.066697f
C99 VN.n6 B 0.076683f
C100 VN.n7 B 1.07965f
C101 VTAIL.t11 B 0.131036f
C102 VTAIL.t10 B 0.131036f
C103 VTAIL.n0 B 1.02465f
C104 VTAIL.n1 B 0.333666f
C105 VTAIL.n2 B 0.039569f
C106 VTAIL.n3 B 0.027363f
C107 VTAIL.n4 B 0.014704f
C108 VTAIL.n5 B 0.034754f
C109 VTAIL.n6 B 0.015569f
C110 VTAIL.n7 B 0.027363f
C111 VTAIL.n8 B 0.014704f
C112 VTAIL.n9 B 0.034754f
C113 VTAIL.n10 B 0.015569f
C114 VTAIL.n11 B 0.11755f
C115 VTAIL.t5 B 0.056672f
C116 VTAIL.n12 B 0.026066f
C117 VTAIL.n13 B 0.020529f
C118 VTAIL.n14 B 0.014704f
C119 VTAIL.n15 B 0.658537f
C120 VTAIL.n16 B 0.027363f
C121 VTAIL.n17 B 0.014704f
C122 VTAIL.n18 B 0.015569f
C123 VTAIL.n19 B 0.034754f
C124 VTAIL.n20 B 0.034754f
C125 VTAIL.n21 B 0.015569f
C126 VTAIL.n22 B 0.014704f
C127 VTAIL.n23 B 0.027363f
C128 VTAIL.n24 B 0.027363f
C129 VTAIL.n25 B 0.014704f
C130 VTAIL.n26 B 0.015569f
C131 VTAIL.n27 B 0.034754f
C132 VTAIL.n28 B 0.077196f
C133 VTAIL.n29 B 0.015569f
C134 VTAIL.n30 B 0.014704f
C135 VTAIL.n31 B 0.065491f
C136 VTAIL.n32 B 0.043463f
C137 VTAIL.n33 B 0.131049f
C138 VTAIL.t7 B 0.131036f
C139 VTAIL.t9 B 0.131036f
C140 VTAIL.n34 B 1.02465f
C141 VTAIL.n35 B 1.2169f
C142 VTAIL.t0 B 0.131036f
C143 VTAIL.t3 B 0.131036f
C144 VTAIL.n36 B 1.02465f
C145 VTAIL.n37 B 1.21689f
C146 VTAIL.n38 B 0.039569f
C147 VTAIL.n39 B 0.027363f
C148 VTAIL.n40 B 0.014704f
C149 VTAIL.n41 B 0.034754f
C150 VTAIL.n42 B 0.015569f
C151 VTAIL.n43 B 0.027363f
C152 VTAIL.n44 B 0.014704f
C153 VTAIL.n45 B 0.034754f
C154 VTAIL.n46 B 0.015569f
C155 VTAIL.n47 B 0.11755f
C156 VTAIL.t1 B 0.056672f
C157 VTAIL.n48 B 0.026066f
C158 VTAIL.n49 B 0.020529f
C159 VTAIL.n50 B 0.014704f
C160 VTAIL.n51 B 0.658537f
C161 VTAIL.n52 B 0.027363f
C162 VTAIL.n53 B 0.014704f
C163 VTAIL.n54 B 0.015569f
C164 VTAIL.n55 B 0.034754f
C165 VTAIL.n56 B 0.034754f
C166 VTAIL.n57 B 0.015569f
C167 VTAIL.n58 B 0.014704f
C168 VTAIL.n59 B 0.027363f
C169 VTAIL.n60 B 0.027363f
C170 VTAIL.n61 B 0.014704f
C171 VTAIL.n62 B 0.015569f
C172 VTAIL.n63 B 0.034754f
C173 VTAIL.n64 B 0.077196f
C174 VTAIL.n65 B 0.015569f
C175 VTAIL.n66 B 0.014704f
C176 VTAIL.n67 B 0.065491f
C177 VTAIL.n68 B 0.043463f
C178 VTAIL.n69 B 0.131049f
C179 VTAIL.t4 B 0.131036f
C180 VTAIL.t8 B 0.131036f
C181 VTAIL.n70 B 1.02465f
C182 VTAIL.n71 B 0.361022f
C183 VTAIL.n72 B 0.039569f
C184 VTAIL.n73 B 0.027363f
C185 VTAIL.n74 B 0.014704f
C186 VTAIL.n75 B 0.034754f
C187 VTAIL.n76 B 0.015569f
C188 VTAIL.n77 B 0.027363f
C189 VTAIL.n78 B 0.014704f
C190 VTAIL.n79 B 0.034754f
C191 VTAIL.n80 B 0.015569f
C192 VTAIL.n81 B 0.11755f
C193 VTAIL.t6 B 0.056672f
C194 VTAIL.n82 B 0.026066f
C195 VTAIL.n83 B 0.020529f
C196 VTAIL.n84 B 0.014704f
C197 VTAIL.n85 B 0.658537f
C198 VTAIL.n86 B 0.027363f
C199 VTAIL.n87 B 0.014704f
C200 VTAIL.n88 B 0.015569f
C201 VTAIL.n89 B 0.034754f
C202 VTAIL.n90 B 0.034754f
C203 VTAIL.n91 B 0.015569f
C204 VTAIL.n92 B 0.014704f
C205 VTAIL.n93 B 0.027363f
C206 VTAIL.n94 B 0.027363f
C207 VTAIL.n95 B 0.014704f
C208 VTAIL.n96 B 0.015569f
C209 VTAIL.n97 B 0.034754f
C210 VTAIL.n98 B 0.077196f
C211 VTAIL.n99 B 0.015569f
C212 VTAIL.n100 B 0.014704f
C213 VTAIL.n101 B 0.065491f
C214 VTAIL.n102 B 0.043463f
C215 VTAIL.n103 B 0.943593f
C216 VTAIL.n104 B 0.039569f
C217 VTAIL.n105 B 0.027363f
C218 VTAIL.n106 B 0.014704f
C219 VTAIL.n107 B 0.034754f
C220 VTAIL.n108 B 0.015569f
C221 VTAIL.n109 B 0.027363f
C222 VTAIL.n110 B 0.014704f
C223 VTAIL.n111 B 0.034754f
C224 VTAIL.n112 B 0.015569f
C225 VTAIL.n113 B 0.11755f
C226 VTAIL.t2 B 0.056672f
C227 VTAIL.n114 B 0.026066f
C228 VTAIL.n115 B 0.020529f
C229 VTAIL.n116 B 0.014704f
C230 VTAIL.n117 B 0.658537f
C231 VTAIL.n118 B 0.027363f
C232 VTAIL.n119 B 0.014704f
C233 VTAIL.n120 B 0.015569f
C234 VTAIL.n121 B 0.034754f
C235 VTAIL.n122 B 0.034754f
C236 VTAIL.n123 B 0.015569f
C237 VTAIL.n124 B 0.014704f
C238 VTAIL.n125 B 0.027363f
C239 VTAIL.n126 B 0.027363f
C240 VTAIL.n127 B 0.014704f
C241 VTAIL.n128 B 0.015569f
C242 VTAIL.n129 B 0.034754f
C243 VTAIL.n130 B 0.077196f
C244 VTAIL.n131 B 0.015569f
C245 VTAIL.n132 B 0.014704f
C246 VTAIL.n133 B 0.065491f
C247 VTAIL.n134 B 0.043463f
C248 VTAIL.n135 B 0.927631f
C249 VDD1.n0 B 0.035337f
C250 VDD1.n1 B 0.024436f
C251 VDD1.n2 B 0.013131f
C252 VDD1.n3 B 0.031037f
C253 VDD1.n4 B 0.013903f
C254 VDD1.n5 B 0.024436f
C255 VDD1.n6 B 0.013131f
C256 VDD1.n7 B 0.031037f
C257 VDD1.n8 B 0.013903f
C258 VDD1.n9 B 0.104977f
C259 VDD1.t3 B 0.05061f
C260 VDD1.n10 B 0.023278f
C261 VDD1.n11 B 0.018333f
C262 VDD1.n12 B 0.013131f
C263 VDD1.n13 B 0.588102f
C264 VDD1.n14 B 0.024436f
C265 VDD1.n15 B 0.013131f
C266 VDD1.n16 B 0.013903f
C267 VDD1.n17 B 0.031037f
C268 VDD1.n18 B 0.031037f
C269 VDD1.n19 B 0.013903f
C270 VDD1.n20 B 0.013131f
C271 VDD1.n21 B 0.024436f
C272 VDD1.n22 B 0.024436f
C273 VDD1.n23 B 0.013131f
C274 VDD1.n24 B 0.013903f
C275 VDD1.n25 B 0.031037f
C276 VDD1.n26 B 0.068939f
C277 VDD1.n27 B 0.013903f
C278 VDD1.n28 B 0.013131f
C279 VDD1.n29 B 0.058486f
C280 VDD1.n30 B 0.056364f
C281 VDD1.n31 B 0.035337f
C282 VDD1.n32 B 0.024436f
C283 VDD1.n33 B 0.013131f
C284 VDD1.n34 B 0.031037f
C285 VDD1.n35 B 0.013903f
C286 VDD1.n36 B 0.024436f
C287 VDD1.n37 B 0.013131f
C288 VDD1.n38 B 0.031037f
C289 VDD1.n39 B 0.013903f
C290 VDD1.n40 B 0.104977f
C291 VDD1.t1 B 0.05061f
C292 VDD1.n41 B 0.023278f
C293 VDD1.n42 B 0.018333f
C294 VDD1.n43 B 0.013131f
C295 VDD1.n44 B 0.588102f
C296 VDD1.n45 B 0.024436f
C297 VDD1.n46 B 0.013131f
C298 VDD1.n47 B 0.013903f
C299 VDD1.n48 B 0.031037f
C300 VDD1.n49 B 0.031037f
C301 VDD1.n50 B 0.013903f
C302 VDD1.n51 B 0.013131f
C303 VDD1.n52 B 0.024436f
C304 VDD1.n53 B 0.024436f
C305 VDD1.n54 B 0.013131f
C306 VDD1.n55 B 0.013903f
C307 VDD1.n56 B 0.031037f
C308 VDD1.n57 B 0.068939f
C309 VDD1.n58 B 0.013903f
C310 VDD1.n59 B 0.013131f
C311 VDD1.n60 B 0.058486f
C312 VDD1.n61 B 0.056137f
C313 VDD1.t0 B 0.117021f
C314 VDD1.t4 B 0.117021f
C315 VDD1.n62 B 0.977762f
C316 VDD1.n63 B 1.33294f
C317 VDD1.t2 B 0.117021f
C318 VDD1.t5 B 0.117021f
C319 VDD1.n64 B 0.977505f
C320 VDD1.n65 B 1.60988f
C321 VP.t5 B 0.147161f
C322 VP.n0 B 0.077796f
C323 VP.t1 B 0.143063f
C324 VP.n1 B 0.067622f
C325 VP.t3 B 0.147161f
C326 VP.n2 B 0.077746f
C327 VP.n3 B 1.07167f
C328 VP.n4 B 1.06466f
C329 VP.t0 B 0.143063f
C330 VP.t2 B 0.147161f
C331 VP.n5 B 0.077746f
C332 VP.n6 B 0.067622f
C333 VP.t4 B 0.147161f
C334 VP.n7 B 0.077746f
C335 VP.n8 B 0.026759f
.ends

