* NGSPICE file created from diff_pair_sample_0722.ext - technology: sky130A

.subckt diff_pair_sample_0722 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t5 VN.t0 VTAIL.t7 B.t4 sky130_fd_pr__nfet_01v8 ad=1.1022 pd=7.01 as=2.6052 ps=14.14 w=6.68 l=2.23
X1 B.t19 B.t17 B.t18 B.t14 sky130_fd_pr__nfet_01v8 ad=2.6052 pd=14.14 as=0 ps=0 w=6.68 l=2.23
X2 VTAIL.t11 VP.t0 VDD1.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=1.1022 pd=7.01 as=1.1022 ps=7.01 w=6.68 l=2.23
X3 VTAIL.t6 VN.t1 VDD2.t4 B.t5 sky130_fd_pr__nfet_01v8 ad=1.1022 pd=7.01 as=1.1022 ps=7.01 w=6.68 l=2.23
X4 VTAIL.t8 VN.t2 VDD2.t3 B.t1 sky130_fd_pr__nfet_01v8 ad=1.1022 pd=7.01 as=1.1022 ps=7.01 w=6.68 l=2.23
X5 B.t16 B.t13 B.t15 B.t14 sky130_fd_pr__nfet_01v8 ad=2.6052 pd=14.14 as=0 ps=0 w=6.68 l=2.23
X6 VDD1.t4 VP.t1 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=2.6052 pd=14.14 as=1.1022 ps=7.01 w=6.68 l=2.23
X7 VDD1.t3 VP.t2 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=1.1022 pd=7.01 as=2.6052 ps=14.14 w=6.68 l=2.23
X8 B.t12 B.t10 B.t11 B.t7 sky130_fd_pr__nfet_01v8 ad=2.6052 pd=14.14 as=0 ps=0 w=6.68 l=2.23
X9 VDD2.t2 VN.t3 VTAIL.t9 B.t2 sky130_fd_pr__nfet_01v8 ad=2.6052 pd=14.14 as=1.1022 ps=7.01 w=6.68 l=2.23
X10 B.t9 B.t6 B.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=2.6052 pd=14.14 as=0 ps=0 w=6.68 l=2.23
X11 VDD1.t2 VP.t3 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=2.6052 pd=14.14 as=1.1022 ps=7.01 w=6.68 l=2.23
X12 VDD2.t1 VN.t4 VTAIL.t5 B.t0 sky130_fd_pr__nfet_01v8 ad=1.1022 pd=7.01 as=2.6052 ps=14.14 w=6.68 l=2.23
X13 VDD1.t1 VP.t4 VTAIL.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=1.1022 pd=7.01 as=2.6052 ps=14.14 w=6.68 l=2.23
X14 VTAIL.t1 VP.t5 VDD1.t0 B.t1 sky130_fd_pr__nfet_01v8 ad=1.1022 pd=7.01 as=1.1022 ps=7.01 w=6.68 l=2.23
X15 VDD2.t0 VN.t5 VTAIL.t10 B.t3 sky130_fd_pr__nfet_01v8 ad=2.6052 pd=14.14 as=1.1022 ps=7.01 w=6.68 l=2.23
R0 VN.n25 VN.n14 161.3
R1 VN.n24 VN.n23 161.3
R2 VN.n22 VN.n15 161.3
R3 VN.n21 VN.n20 161.3
R4 VN.n19 VN.n16 161.3
R5 VN.n11 VN.n0 161.3
R6 VN.n10 VN.n9 161.3
R7 VN.n8 VN.n1 161.3
R8 VN.n7 VN.n6 161.3
R9 VN.n5 VN.n2 161.3
R10 VN.n3 VN.t3 105.103
R11 VN.n17 VN.t4 105.103
R12 VN.n13 VN.n12 95.6613
R13 VN.n27 VN.n26 95.6613
R14 VN.n4 VN.t2 72.1924
R15 VN.n12 VN.t0 72.1924
R16 VN.n18 VN.t1 72.1924
R17 VN.n26 VN.t5 72.1924
R18 VN.n4 VN.n3 59.417
R19 VN.n18 VN.n17 59.417
R20 VN.n10 VN.n1 43.4833
R21 VN.n24 VN.n15 43.4833
R22 VN VN.n27 43.483
R23 VN.n6 VN.n1 37.6707
R24 VN.n20 VN.n15 37.6707
R25 VN.n6 VN.n5 24.5923
R26 VN.n11 VN.n10 24.5923
R27 VN.n20 VN.n19 24.5923
R28 VN.n25 VN.n24 24.5923
R29 VN.n12 VN.n11 15.2474
R30 VN.n26 VN.n25 15.2474
R31 VN.n5 VN.n4 12.2964
R32 VN.n19 VN.n18 12.2964
R33 VN.n17 VN.n16 9.41768
R34 VN.n3 VN.n2 9.41768
R35 VN.n27 VN.n14 0.278335
R36 VN.n13 VN.n0 0.278335
R37 VN.n23 VN.n14 0.189894
R38 VN.n23 VN.n22 0.189894
R39 VN.n22 VN.n21 0.189894
R40 VN.n21 VN.n16 0.189894
R41 VN.n7 VN.n2 0.189894
R42 VN.n8 VN.n7 0.189894
R43 VN.n9 VN.n8 0.189894
R44 VN.n9 VN.n0 0.189894
R45 VN VN.n13 0.153485
R46 VTAIL.n146 VTAIL.n116 289.615
R47 VTAIL.n32 VTAIL.n2 289.615
R48 VTAIL.n110 VTAIL.n80 289.615
R49 VTAIL.n72 VTAIL.n42 289.615
R50 VTAIL.n129 VTAIL.n128 185
R51 VTAIL.n131 VTAIL.n130 185
R52 VTAIL.n124 VTAIL.n123 185
R53 VTAIL.n137 VTAIL.n136 185
R54 VTAIL.n139 VTAIL.n138 185
R55 VTAIL.n120 VTAIL.n119 185
R56 VTAIL.n145 VTAIL.n144 185
R57 VTAIL.n147 VTAIL.n146 185
R58 VTAIL.n15 VTAIL.n14 185
R59 VTAIL.n17 VTAIL.n16 185
R60 VTAIL.n10 VTAIL.n9 185
R61 VTAIL.n23 VTAIL.n22 185
R62 VTAIL.n25 VTAIL.n24 185
R63 VTAIL.n6 VTAIL.n5 185
R64 VTAIL.n31 VTAIL.n30 185
R65 VTAIL.n33 VTAIL.n32 185
R66 VTAIL.n111 VTAIL.n110 185
R67 VTAIL.n109 VTAIL.n108 185
R68 VTAIL.n84 VTAIL.n83 185
R69 VTAIL.n103 VTAIL.n102 185
R70 VTAIL.n101 VTAIL.n100 185
R71 VTAIL.n88 VTAIL.n87 185
R72 VTAIL.n95 VTAIL.n94 185
R73 VTAIL.n93 VTAIL.n92 185
R74 VTAIL.n73 VTAIL.n72 185
R75 VTAIL.n71 VTAIL.n70 185
R76 VTAIL.n46 VTAIL.n45 185
R77 VTAIL.n65 VTAIL.n64 185
R78 VTAIL.n63 VTAIL.n62 185
R79 VTAIL.n50 VTAIL.n49 185
R80 VTAIL.n57 VTAIL.n56 185
R81 VTAIL.n55 VTAIL.n54 185
R82 VTAIL.n127 VTAIL.t7 147.659
R83 VTAIL.n13 VTAIL.t0 147.659
R84 VTAIL.n91 VTAIL.t4 147.659
R85 VTAIL.n53 VTAIL.t5 147.659
R86 VTAIL.n130 VTAIL.n129 104.615
R87 VTAIL.n130 VTAIL.n123 104.615
R88 VTAIL.n137 VTAIL.n123 104.615
R89 VTAIL.n138 VTAIL.n137 104.615
R90 VTAIL.n138 VTAIL.n119 104.615
R91 VTAIL.n145 VTAIL.n119 104.615
R92 VTAIL.n146 VTAIL.n145 104.615
R93 VTAIL.n16 VTAIL.n15 104.615
R94 VTAIL.n16 VTAIL.n9 104.615
R95 VTAIL.n23 VTAIL.n9 104.615
R96 VTAIL.n24 VTAIL.n23 104.615
R97 VTAIL.n24 VTAIL.n5 104.615
R98 VTAIL.n31 VTAIL.n5 104.615
R99 VTAIL.n32 VTAIL.n31 104.615
R100 VTAIL.n110 VTAIL.n109 104.615
R101 VTAIL.n109 VTAIL.n83 104.615
R102 VTAIL.n102 VTAIL.n83 104.615
R103 VTAIL.n102 VTAIL.n101 104.615
R104 VTAIL.n101 VTAIL.n87 104.615
R105 VTAIL.n94 VTAIL.n87 104.615
R106 VTAIL.n94 VTAIL.n93 104.615
R107 VTAIL.n72 VTAIL.n71 104.615
R108 VTAIL.n71 VTAIL.n45 104.615
R109 VTAIL.n64 VTAIL.n45 104.615
R110 VTAIL.n64 VTAIL.n63 104.615
R111 VTAIL.n63 VTAIL.n49 104.615
R112 VTAIL.n56 VTAIL.n49 104.615
R113 VTAIL.n56 VTAIL.n55 104.615
R114 VTAIL.n129 VTAIL.t7 52.3082
R115 VTAIL.n15 VTAIL.t0 52.3082
R116 VTAIL.n93 VTAIL.t4 52.3082
R117 VTAIL.n55 VTAIL.t5 52.3082
R118 VTAIL.n79 VTAIL.n78 48.6196
R119 VTAIL.n41 VTAIL.n40 48.6196
R120 VTAIL.n1 VTAIL.n0 48.6194
R121 VTAIL.n39 VTAIL.n38 48.6194
R122 VTAIL.n151 VTAIL.n150 31.4096
R123 VTAIL.n37 VTAIL.n36 31.4096
R124 VTAIL.n115 VTAIL.n114 31.4096
R125 VTAIL.n77 VTAIL.n76 31.4096
R126 VTAIL.n41 VTAIL.n39 22.5393
R127 VTAIL.n151 VTAIL.n115 20.3324
R128 VTAIL.n128 VTAIL.n127 15.6676
R129 VTAIL.n14 VTAIL.n13 15.6676
R130 VTAIL.n92 VTAIL.n91 15.6676
R131 VTAIL.n54 VTAIL.n53 15.6676
R132 VTAIL.n131 VTAIL.n126 12.8005
R133 VTAIL.n17 VTAIL.n12 12.8005
R134 VTAIL.n95 VTAIL.n90 12.8005
R135 VTAIL.n57 VTAIL.n52 12.8005
R136 VTAIL.n132 VTAIL.n124 12.0247
R137 VTAIL.n18 VTAIL.n10 12.0247
R138 VTAIL.n96 VTAIL.n88 12.0247
R139 VTAIL.n58 VTAIL.n50 12.0247
R140 VTAIL.n136 VTAIL.n135 11.249
R141 VTAIL.n22 VTAIL.n21 11.249
R142 VTAIL.n100 VTAIL.n99 11.249
R143 VTAIL.n62 VTAIL.n61 11.249
R144 VTAIL.n139 VTAIL.n122 10.4732
R145 VTAIL.n25 VTAIL.n8 10.4732
R146 VTAIL.n103 VTAIL.n86 10.4732
R147 VTAIL.n65 VTAIL.n48 10.4732
R148 VTAIL.n140 VTAIL.n120 9.69747
R149 VTAIL.n26 VTAIL.n6 9.69747
R150 VTAIL.n104 VTAIL.n84 9.69747
R151 VTAIL.n66 VTAIL.n46 9.69747
R152 VTAIL.n150 VTAIL.n149 9.45567
R153 VTAIL.n36 VTAIL.n35 9.45567
R154 VTAIL.n114 VTAIL.n113 9.45567
R155 VTAIL.n76 VTAIL.n75 9.45567
R156 VTAIL.n118 VTAIL.n117 9.3005
R157 VTAIL.n143 VTAIL.n142 9.3005
R158 VTAIL.n141 VTAIL.n140 9.3005
R159 VTAIL.n122 VTAIL.n121 9.3005
R160 VTAIL.n135 VTAIL.n134 9.3005
R161 VTAIL.n133 VTAIL.n132 9.3005
R162 VTAIL.n126 VTAIL.n125 9.3005
R163 VTAIL.n149 VTAIL.n148 9.3005
R164 VTAIL.n4 VTAIL.n3 9.3005
R165 VTAIL.n29 VTAIL.n28 9.3005
R166 VTAIL.n27 VTAIL.n26 9.3005
R167 VTAIL.n8 VTAIL.n7 9.3005
R168 VTAIL.n21 VTAIL.n20 9.3005
R169 VTAIL.n19 VTAIL.n18 9.3005
R170 VTAIL.n12 VTAIL.n11 9.3005
R171 VTAIL.n35 VTAIL.n34 9.3005
R172 VTAIL.n113 VTAIL.n112 9.3005
R173 VTAIL.n82 VTAIL.n81 9.3005
R174 VTAIL.n107 VTAIL.n106 9.3005
R175 VTAIL.n105 VTAIL.n104 9.3005
R176 VTAIL.n86 VTAIL.n85 9.3005
R177 VTAIL.n99 VTAIL.n98 9.3005
R178 VTAIL.n97 VTAIL.n96 9.3005
R179 VTAIL.n90 VTAIL.n89 9.3005
R180 VTAIL.n75 VTAIL.n74 9.3005
R181 VTAIL.n44 VTAIL.n43 9.3005
R182 VTAIL.n69 VTAIL.n68 9.3005
R183 VTAIL.n67 VTAIL.n66 9.3005
R184 VTAIL.n48 VTAIL.n47 9.3005
R185 VTAIL.n61 VTAIL.n60 9.3005
R186 VTAIL.n59 VTAIL.n58 9.3005
R187 VTAIL.n52 VTAIL.n51 9.3005
R188 VTAIL.n144 VTAIL.n143 8.92171
R189 VTAIL.n30 VTAIL.n29 8.92171
R190 VTAIL.n108 VTAIL.n107 8.92171
R191 VTAIL.n70 VTAIL.n69 8.92171
R192 VTAIL.n147 VTAIL.n118 8.14595
R193 VTAIL.n33 VTAIL.n4 8.14595
R194 VTAIL.n111 VTAIL.n82 8.14595
R195 VTAIL.n73 VTAIL.n44 8.14595
R196 VTAIL.n148 VTAIL.n116 7.3702
R197 VTAIL.n34 VTAIL.n2 7.3702
R198 VTAIL.n112 VTAIL.n80 7.3702
R199 VTAIL.n74 VTAIL.n42 7.3702
R200 VTAIL.n150 VTAIL.n116 6.59444
R201 VTAIL.n36 VTAIL.n2 6.59444
R202 VTAIL.n114 VTAIL.n80 6.59444
R203 VTAIL.n76 VTAIL.n42 6.59444
R204 VTAIL.n148 VTAIL.n147 5.81868
R205 VTAIL.n34 VTAIL.n33 5.81868
R206 VTAIL.n112 VTAIL.n111 5.81868
R207 VTAIL.n74 VTAIL.n73 5.81868
R208 VTAIL.n144 VTAIL.n118 5.04292
R209 VTAIL.n30 VTAIL.n4 5.04292
R210 VTAIL.n108 VTAIL.n82 5.04292
R211 VTAIL.n70 VTAIL.n44 5.04292
R212 VTAIL.n127 VTAIL.n125 4.38571
R213 VTAIL.n13 VTAIL.n11 4.38571
R214 VTAIL.n91 VTAIL.n89 4.38571
R215 VTAIL.n53 VTAIL.n51 4.38571
R216 VTAIL.n143 VTAIL.n120 4.26717
R217 VTAIL.n29 VTAIL.n6 4.26717
R218 VTAIL.n107 VTAIL.n84 4.26717
R219 VTAIL.n69 VTAIL.n46 4.26717
R220 VTAIL.n140 VTAIL.n139 3.49141
R221 VTAIL.n26 VTAIL.n25 3.49141
R222 VTAIL.n104 VTAIL.n103 3.49141
R223 VTAIL.n66 VTAIL.n65 3.49141
R224 VTAIL.n0 VTAIL.t9 2.96457
R225 VTAIL.n0 VTAIL.t8 2.96457
R226 VTAIL.n38 VTAIL.t3 2.96457
R227 VTAIL.n38 VTAIL.t11 2.96457
R228 VTAIL.n78 VTAIL.t2 2.96457
R229 VTAIL.n78 VTAIL.t1 2.96457
R230 VTAIL.n40 VTAIL.t10 2.96457
R231 VTAIL.n40 VTAIL.t6 2.96457
R232 VTAIL.n136 VTAIL.n122 2.71565
R233 VTAIL.n22 VTAIL.n8 2.71565
R234 VTAIL.n100 VTAIL.n86 2.71565
R235 VTAIL.n62 VTAIL.n48 2.71565
R236 VTAIL.n77 VTAIL.n41 2.2074
R237 VTAIL.n115 VTAIL.n79 2.2074
R238 VTAIL.n39 VTAIL.n37 2.2074
R239 VTAIL.n135 VTAIL.n124 1.93989
R240 VTAIL.n21 VTAIL.n10 1.93989
R241 VTAIL.n99 VTAIL.n88 1.93989
R242 VTAIL.n61 VTAIL.n50 1.93989
R243 VTAIL VTAIL.n151 1.59748
R244 VTAIL.n79 VTAIL.n77 1.57378
R245 VTAIL.n37 VTAIL.n1 1.57378
R246 VTAIL.n132 VTAIL.n131 1.16414
R247 VTAIL.n18 VTAIL.n17 1.16414
R248 VTAIL.n96 VTAIL.n95 1.16414
R249 VTAIL.n58 VTAIL.n57 1.16414
R250 VTAIL VTAIL.n1 0.610414
R251 VTAIL.n128 VTAIL.n126 0.388379
R252 VTAIL.n14 VTAIL.n12 0.388379
R253 VTAIL.n92 VTAIL.n90 0.388379
R254 VTAIL.n54 VTAIL.n52 0.388379
R255 VTAIL.n133 VTAIL.n125 0.155672
R256 VTAIL.n134 VTAIL.n133 0.155672
R257 VTAIL.n134 VTAIL.n121 0.155672
R258 VTAIL.n141 VTAIL.n121 0.155672
R259 VTAIL.n142 VTAIL.n141 0.155672
R260 VTAIL.n142 VTAIL.n117 0.155672
R261 VTAIL.n149 VTAIL.n117 0.155672
R262 VTAIL.n19 VTAIL.n11 0.155672
R263 VTAIL.n20 VTAIL.n19 0.155672
R264 VTAIL.n20 VTAIL.n7 0.155672
R265 VTAIL.n27 VTAIL.n7 0.155672
R266 VTAIL.n28 VTAIL.n27 0.155672
R267 VTAIL.n28 VTAIL.n3 0.155672
R268 VTAIL.n35 VTAIL.n3 0.155672
R269 VTAIL.n113 VTAIL.n81 0.155672
R270 VTAIL.n106 VTAIL.n81 0.155672
R271 VTAIL.n106 VTAIL.n105 0.155672
R272 VTAIL.n105 VTAIL.n85 0.155672
R273 VTAIL.n98 VTAIL.n85 0.155672
R274 VTAIL.n98 VTAIL.n97 0.155672
R275 VTAIL.n97 VTAIL.n89 0.155672
R276 VTAIL.n75 VTAIL.n43 0.155672
R277 VTAIL.n68 VTAIL.n43 0.155672
R278 VTAIL.n68 VTAIL.n67 0.155672
R279 VTAIL.n67 VTAIL.n47 0.155672
R280 VTAIL.n60 VTAIL.n47 0.155672
R281 VTAIL.n60 VTAIL.n59 0.155672
R282 VTAIL.n59 VTAIL.n51 0.155672
R283 VDD2.n67 VDD2.n37 289.615
R284 VDD2.n30 VDD2.n0 289.615
R285 VDD2.n68 VDD2.n67 185
R286 VDD2.n66 VDD2.n65 185
R287 VDD2.n41 VDD2.n40 185
R288 VDD2.n60 VDD2.n59 185
R289 VDD2.n58 VDD2.n57 185
R290 VDD2.n45 VDD2.n44 185
R291 VDD2.n52 VDD2.n51 185
R292 VDD2.n50 VDD2.n49 185
R293 VDD2.n13 VDD2.n12 185
R294 VDD2.n15 VDD2.n14 185
R295 VDD2.n8 VDD2.n7 185
R296 VDD2.n21 VDD2.n20 185
R297 VDD2.n23 VDD2.n22 185
R298 VDD2.n4 VDD2.n3 185
R299 VDD2.n29 VDD2.n28 185
R300 VDD2.n31 VDD2.n30 185
R301 VDD2.n48 VDD2.t0 147.659
R302 VDD2.n11 VDD2.t2 147.659
R303 VDD2.n67 VDD2.n66 104.615
R304 VDD2.n66 VDD2.n40 104.615
R305 VDD2.n59 VDD2.n40 104.615
R306 VDD2.n59 VDD2.n58 104.615
R307 VDD2.n58 VDD2.n44 104.615
R308 VDD2.n51 VDD2.n44 104.615
R309 VDD2.n51 VDD2.n50 104.615
R310 VDD2.n14 VDD2.n13 104.615
R311 VDD2.n14 VDD2.n7 104.615
R312 VDD2.n21 VDD2.n7 104.615
R313 VDD2.n22 VDD2.n21 104.615
R314 VDD2.n22 VDD2.n3 104.615
R315 VDD2.n29 VDD2.n3 104.615
R316 VDD2.n30 VDD2.n29 104.615
R317 VDD2.n36 VDD2.n35 65.7946
R318 VDD2 VDD2.n73 65.7917
R319 VDD2.n50 VDD2.t0 52.3082
R320 VDD2.n13 VDD2.t2 52.3082
R321 VDD2.n36 VDD2.n34 49.6882
R322 VDD2.n72 VDD2.n71 48.0884
R323 VDD2.n72 VDD2.n36 36.6463
R324 VDD2.n49 VDD2.n48 15.6676
R325 VDD2.n12 VDD2.n11 15.6676
R326 VDD2.n52 VDD2.n47 12.8005
R327 VDD2.n15 VDD2.n10 12.8005
R328 VDD2.n53 VDD2.n45 12.0247
R329 VDD2.n16 VDD2.n8 12.0247
R330 VDD2.n57 VDD2.n56 11.249
R331 VDD2.n20 VDD2.n19 11.249
R332 VDD2.n60 VDD2.n43 10.4732
R333 VDD2.n23 VDD2.n6 10.4732
R334 VDD2.n61 VDD2.n41 9.69747
R335 VDD2.n24 VDD2.n4 9.69747
R336 VDD2.n71 VDD2.n70 9.45567
R337 VDD2.n34 VDD2.n33 9.45567
R338 VDD2.n70 VDD2.n69 9.3005
R339 VDD2.n39 VDD2.n38 9.3005
R340 VDD2.n64 VDD2.n63 9.3005
R341 VDD2.n62 VDD2.n61 9.3005
R342 VDD2.n43 VDD2.n42 9.3005
R343 VDD2.n56 VDD2.n55 9.3005
R344 VDD2.n54 VDD2.n53 9.3005
R345 VDD2.n47 VDD2.n46 9.3005
R346 VDD2.n2 VDD2.n1 9.3005
R347 VDD2.n27 VDD2.n26 9.3005
R348 VDD2.n25 VDD2.n24 9.3005
R349 VDD2.n6 VDD2.n5 9.3005
R350 VDD2.n19 VDD2.n18 9.3005
R351 VDD2.n17 VDD2.n16 9.3005
R352 VDD2.n10 VDD2.n9 9.3005
R353 VDD2.n33 VDD2.n32 9.3005
R354 VDD2.n65 VDD2.n64 8.92171
R355 VDD2.n28 VDD2.n27 8.92171
R356 VDD2.n68 VDD2.n39 8.14595
R357 VDD2.n31 VDD2.n2 8.14595
R358 VDD2.n69 VDD2.n37 7.3702
R359 VDD2.n32 VDD2.n0 7.3702
R360 VDD2.n71 VDD2.n37 6.59444
R361 VDD2.n34 VDD2.n0 6.59444
R362 VDD2.n69 VDD2.n68 5.81868
R363 VDD2.n32 VDD2.n31 5.81868
R364 VDD2.n65 VDD2.n39 5.04292
R365 VDD2.n28 VDD2.n2 5.04292
R366 VDD2.n48 VDD2.n46 4.38571
R367 VDD2.n11 VDD2.n9 4.38571
R368 VDD2.n64 VDD2.n41 4.26717
R369 VDD2.n27 VDD2.n4 4.26717
R370 VDD2.n61 VDD2.n60 3.49141
R371 VDD2.n24 VDD2.n23 3.49141
R372 VDD2.n73 VDD2.t4 2.96457
R373 VDD2.n73 VDD2.t1 2.96457
R374 VDD2.n35 VDD2.t3 2.96457
R375 VDD2.n35 VDD2.t5 2.96457
R376 VDD2.n57 VDD2.n43 2.71565
R377 VDD2.n20 VDD2.n6 2.71565
R378 VDD2.n56 VDD2.n45 1.93989
R379 VDD2.n19 VDD2.n8 1.93989
R380 VDD2 VDD2.n72 1.71386
R381 VDD2.n53 VDD2.n52 1.16414
R382 VDD2.n16 VDD2.n15 1.16414
R383 VDD2.n49 VDD2.n47 0.388379
R384 VDD2.n12 VDD2.n10 0.388379
R385 VDD2.n70 VDD2.n38 0.155672
R386 VDD2.n63 VDD2.n38 0.155672
R387 VDD2.n63 VDD2.n62 0.155672
R388 VDD2.n62 VDD2.n42 0.155672
R389 VDD2.n55 VDD2.n42 0.155672
R390 VDD2.n55 VDD2.n54 0.155672
R391 VDD2.n54 VDD2.n46 0.155672
R392 VDD2.n17 VDD2.n9 0.155672
R393 VDD2.n18 VDD2.n17 0.155672
R394 VDD2.n18 VDD2.n5 0.155672
R395 VDD2.n25 VDD2.n5 0.155672
R396 VDD2.n26 VDD2.n25 0.155672
R397 VDD2.n26 VDD2.n1 0.155672
R398 VDD2.n33 VDD2.n1 0.155672
R399 B.n507 B.n506 585
R400 B.n508 B.n108 585
R401 B.n510 B.n509 585
R402 B.n512 B.n107 585
R403 B.n515 B.n514 585
R404 B.n516 B.n106 585
R405 B.n518 B.n517 585
R406 B.n520 B.n105 585
R407 B.n523 B.n522 585
R408 B.n524 B.n104 585
R409 B.n526 B.n525 585
R410 B.n528 B.n103 585
R411 B.n531 B.n530 585
R412 B.n532 B.n102 585
R413 B.n534 B.n533 585
R414 B.n536 B.n101 585
R415 B.n539 B.n538 585
R416 B.n540 B.n100 585
R417 B.n542 B.n541 585
R418 B.n544 B.n99 585
R419 B.n547 B.n546 585
R420 B.n548 B.n98 585
R421 B.n550 B.n549 585
R422 B.n552 B.n97 585
R423 B.n554 B.n553 585
R424 B.n556 B.n555 585
R425 B.n559 B.n558 585
R426 B.n560 B.n92 585
R427 B.n562 B.n561 585
R428 B.n564 B.n91 585
R429 B.n567 B.n566 585
R430 B.n568 B.n90 585
R431 B.n570 B.n569 585
R432 B.n572 B.n89 585
R433 B.n574 B.n573 585
R434 B.n576 B.n575 585
R435 B.n579 B.n578 585
R436 B.n580 B.n84 585
R437 B.n582 B.n581 585
R438 B.n584 B.n83 585
R439 B.n587 B.n586 585
R440 B.n588 B.n82 585
R441 B.n590 B.n589 585
R442 B.n592 B.n81 585
R443 B.n595 B.n594 585
R444 B.n596 B.n80 585
R445 B.n598 B.n597 585
R446 B.n600 B.n79 585
R447 B.n603 B.n602 585
R448 B.n604 B.n78 585
R449 B.n606 B.n605 585
R450 B.n608 B.n77 585
R451 B.n611 B.n610 585
R452 B.n612 B.n76 585
R453 B.n614 B.n613 585
R454 B.n616 B.n75 585
R455 B.n619 B.n618 585
R456 B.n620 B.n74 585
R457 B.n622 B.n621 585
R458 B.n624 B.n73 585
R459 B.n627 B.n626 585
R460 B.n628 B.n72 585
R461 B.n504 B.n70 585
R462 B.n631 B.n70 585
R463 B.n503 B.n69 585
R464 B.n632 B.n69 585
R465 B.n502 B.n68 585
R466 B.n633 B.n68 585
R467 B.n501 B.n500 585
R468 B.n500 B.n64 585
R469 B.n499 B.n63 585
R470 B.n639 B.n63 585
R471 B.n498 B.n62 585
R472 B.n640 B.n62 585
R473 B.n497 B.n61 585
R474 B.n641 B.n61 585
R475 B.n496 B.n495 585
R476 B.n495 B.n57 585
R477 B.n494 B.n56 585
R478 B.n647 B.n56 585
R479 B.n493 B.n55 585
R480 B.n648 B.n55 585
R481 B.n492 B.n54 585
R482 B.n649 B.n54 585
R483 B.n491 B.n490 585
R484 B.n490 B.n50 585
R485 B.n489 B.n49 585
R486 B.n655 B.n49 585
R487 B.n488 B.n48 585
R488 B.n656 B.n48 585
R489 B.n487 B.n47 585
R490 B.n657 B.n47 585
R491 B.n486 B.n485 585
R492 B.n485 B.n43 585
R493 B.n484 B.n42 585
R494 B.n663 B.n42 585
R495 B.n483 B.n41 585
R496 B.n664 B.n41 585
R497 B.n482 B.n40 585
R498 B.n665 B.n40 585
R499 B.n481 B.n480 585
R500 B.n480 B.n36 585
R501 B.n479 B.n35 585
R502 B.n671 B.n35 585
R503 B.n478 B.n34 585
R504 B.n672 B.n34 585
R505 B.n477 B.n33 585
R506 B.n673 B.n33 585
R507 B.n476 B.n475 585
R508 B.n475 B.n29 585
R509 B.n474 B.n28 585
R510 B.n679 B.n28 585
R511 B.n473 B.n27 585
R512 B.n680 B.n27 585
R513 B.n472 B.n26 585
R514 B.n681 B.n26 585
R515 B.n471 B.n470 585
R516 B.n470 B.n22 585
R517 B.n469 B.n21 585
R518 B.n687 B.n21 585
R519 B.n468 B.n20 585
R520 B.n688 B.n20 585
R521 B.n467 B.n19 585
R522 B.n689 B.n19 585
R523 B.n466 B.n465 585
R524 B.n465 B.n15 585
R525 B.n464 B.n14 585
R526 B.n695 B.n14 585
R527 B.n463 B.n13 585
R528 B.n696 B.n13 585
R529 B.n462 B.n12 585
R530 B.n697 B.n12 585
R531 B.n461 B.n460 585
R532 B.n460 B.n8 585
R533 B.n459 B.n7 585
R534 B.n703 B.n7 585
R535 B.n458 B.n6 585
R536 B.n704 B.n6 585
R537 B.n457 B.n5 585
R538 B.n705 B.n5 585
R539 B.n456 B.n455 585
R540 B.n455 B.n4 585
R541 B.n454 B.n109 585
R542 B.n454 B.n453 585
R543 B.n444 B.n110 585
R544 B.n111 B.n110 585
R545 B.n446 B.n445 585
R546 B.n447 B.n446 585
R547 B.n443 B.n116 585
R548 B.n116 B.n115 585
R549 B.n442 B.n441 585
R550 B.n441 B.n440 585
R551 B.n118 B.n117 585
R552 B.n119 B.n118 585
R553 B.n433 B.n432 585
R554 B.n434 B.n433 585
R555 B.n431 B.n124 585
R556 B.n124 B.n123 585
R557 B.n430 B.n429 585
R558 B.n429 B.n428 585
R559 B.n126 B.n125 585
R560 B.n127 B.n126 585
R561 B.n421 B.n420 585
R562 B.n422 B.n421 585
R563 B.n419 B.n131 585
R564 B.n135 B.n131 585
R565 B.n418 B.n417 585
R566 B.n417 B.n416 585
R567 B.n133 B.n132 585
R568 B.n134 B.n133 585
R569 B.n409 B.n408 585
R570 B.n410 B.n409 585
R571 B.n407 B.n140 585
R572 B.n140 B.n139 585
R573 B.n406 B.n405 585
R574 B.n405 B.n404 585
R575 B.n142 B.n141 585
R576 B.n143 B.n142 585
R577 B.n397 B.n396 585
R578 B.n398 B.n397 585
R579 B.n395 B.n147 585
R580 B.n151 B.n147 585
R581 B.n394 B.n393 585
R582 B.n393 B.n392 585
R583 B.n149 B.n148 585
R584 B.n150 B.n149 585
R585 B.n385 B.n384 585
R586 B.n386 B.n385 585
R587 B.n383 B.n156 585
R588 B.n156 B.n155 585
R589 B.n382 B.n381 585
R590 B.n381 B.n380 585
R591 B.n158 B.n157 585
R592 B.n159 B.n158 585
R593 B.n373 B.n372 585
R594 B.n374 B.n373 585
R595 B.n371 B.n164 585
R596 B.n164 B.n163 585
R597 B.n370 B.n369 585
R598 B.n369 B.n368 585
R599 B.n166 B.n165 585
R600 B.n167 B.n166 585
R601 B.n361 B.n360 585
R602 B.n362 B.n361 585
R603 B.n359 B.n172 585
R604 B.n172 B.n171 585
R605 B.n358 B.n357 585
R606 B.n357 B.n356 585
R607 B.n174 B.n173 585
R608 B.n175 B.n174 585
R609 B.n349 B.n348 585
R610 B.n350 B.n349 585
R611 B.n347 B.n180 585
R612 B.n180 B.n179 585
R613 B.n346 B.n345 585
R614 B.n345 B.n344 585
R615 B.n341 B.n184 585
R616 B.n340 B.n339 585
R617 B.n337 B.n185 585
R618 B.n337 B.n183 585
R619 B.n336 B.n335 585
R620 B.n334 B.n333 585
R621 B.n332 B.n187 585
R622 B.n330 B.n329 585
R623 B.n328 B.n188 585
R624 B.n327 B.n326 585
R625 B.n324 B.n189 585
R626 B.n322 B.n321 585
R627 B.n320 B.n190 585
R628 B.n319 B.n318 585
R629 B.n316 B.n191 585
R630 B.n314 B.n313 585
R631 B.n312 B.n192 585
R632 B.n311 B.n310 585
R633 B.n308 B.n193 585
R634 B.n306 B.n305 585
R635 B.n304 B.n194 585
R636 B.n303 B.n302 585
R637 B.n300 B.n195 585
R638 B.n298 B.n297 585
R639 B.n296 B.n196 585
R640 B.n295 B.n294 585
R641 B.n292 B.n197 585
R642 B.n290 B.n289 585
R643 B.n288 B.n198 585
R644 B.n287 B.n286 585
R645 B.n284 B.n202 585
R646 B.n282 B.n281 585
R647 B.n280 B.n203 585
R648 B.n279 B.n278 585
R649 B.n276 B.n204 585
R650 B.n274 B.n273 585
R651 B.n272 B.n205 585
R652 B.n270 B.n269 585
R653 B.n267 B.n208 585
R654 B.n265 B.n264 585
R655 B.n263 B.n209 585
R656 B.n262 B.n261 585
R657 B.n259 B.n210 585
R658 B.n257 B.n256 585
R659 B.n255 B.n211 585
R660 B.n254 B.n253 585
R661 B.n251 B.n212 585
R662 B.n249 B.n248 585
R663 B.n247 B.n213 585
R664 B.n246 B.n245 585
R665 B.n243 B.n214 585
R666 B.n241 B.n240 585
R667 B.n239 B.n215 585
R668 B.n238 B.n237 585
R669 B.n235 B.n216 585
R670 B.n233 B.n232 585
R671 B.n231 B.n217 585
R672 B.n230 B.n229 585
R673 B.n227 B.n218 585
R674 B.n225 B.n224 585
R675 B.n223 B.n219 585
R676 B.n222 B.n221 585
R677 B.n182 B.n181 585
R678 B.n183 B.n182 585
R679 B.n343 B.n342 585
R680 B.n344 B.n343 585
R681 B.n178 B.n177 585
R682 B.n179 B.n178 585
R683 B.n352 B.n351 585
R684 B.n351 B.n350 585
R685 B.n353 B.n176 585
R686 B.n176 B.n175 585
R687 B.n355 B.n354 585
R688 B.n356 B.n355 585
R689 B.n170 B.n169 585
R690 B.n171 B.n170 585
R691 B.n364 B.n363 585
R692 B.n363 B.n362 585
R693 B.n365 B.n168 585
R694 B.n168 B.n167 585
R695 B.n367 B.n366 585
R696 B.n368 B.n367 585
R697 B.n162 B.n161 585
R698 B.n163 B.n162 585
R699 B.n376 B.n375 585
R700 B.n375 B.n374 585
R701 B.n377 B.n160 585
R702 B.n160 B.n159 585
R703 B.n379 B.n378 585
R704 B.n380 B.n379 585
R705 B.n154 B.n153 585
R706 B.n155 B.n154 585
R707 B.n388 B.n387 585
R708 B.n387 B.n386 585
R709 B.n389 B.n152 585
R710 B.n152 B.n150 585
R711 B.n391 B.n390 585
R712 B.n392 B.n391 585
R713 B.n146 B.n145 585
R714 B.n151 B.n146 585
R715 B.n400 B.n399 585
R716 B.n399 B.n398 585
R717 B.n401 B.n144 585
R718 B.n144 B.n143 585
R719 B.n403 B.n402 585
R720 B.n404 B.n403 585
R721 B.n138 B.n137 585
R722 B.n139 B.n138 585
R723 B.n412 B.n411 585
R724 B.n411 B.n410 585
R725 B.n413 B.n136 585
R726 B.n136 B.n134 585
R727 B.n415 B.n414 585
R728 B.n416 B.n415 585
R729 B.n130 B.n129 585
R730 B.n135 B.n130 585
R731 B.n424 B.n423 585
R732 B.n423 B.n422 585
R733 B.n425 B.n128 585
R734 B.n128 B.n127 585
R735 B.n427 B.n426 585
R736 B.n428 B.n427 585
R737 B.n122 B.n121 585
R738 B.n123 B.n122 585
R739 B.n436 B.n435 585
R740 B.n435 B.n434 585
R741 B.n437 B.n120 585
R742 B.n120 B.n119 585
R743 B.n439 B.n438 585
R744 B.n440 B.n439 585
R745 B.n114 B.n113 585
R746 B.n115 B.n114 585
R747 B.n449 B.n448 585
R748 B.n448 B.n447 585
R749 B.n450 B.n112 585
R750 B.n112 B.n111 585
R751 B.n452 B.n451 585
R752 B.n453 B.n452 585
R753 B.n2 B.n0 585
R754 B.n4 B.n2 585
R755 B.n3 B.n1 585
R756 B.n704 B.n3 585
R757 B.n702 B.n701 585
R758 B.n703 B.n702 585
R759 B.n700 B.n9 585
R760 B.n9 B.n8 585
R761 B.n699 B.n698 585
R762 B.n698 B.n697 585
R763 B.n11 B.n10 585
R764 B.n696 B.n11 585
R765 B.n694 B.n693 585
R766 B.n695 B.n694 585
R767 B.n692 B.n16 585
R768 B.n16 B.n15 585
R769 B.n691 B.n690 585
R770 B.n690 B.n689 585
R771 B.n18 B.n17 585
R772 B.n688 B.n18 585
R773 B.n686 B.n685 585
R774 B.n687 B.n686 585
R775 B.n684 B.n23 585
R776 B.n23 B.n22 585
R777 B.n683 B.n682 585
R778 B.n682 B.n681 585
R779 B.n25 B.n24 585
R780 B.n680 B.n25 585
R781 B.n678 B.n677 585
R782 B.n679 B.n678 585
R783 B.n676 B.n30 585
R784 B.n30 B.n29 585
R785 B.n675 B.n674 585
R786 B.n674 B.n673 585
R787 B.n32 B.n31 585
R788 B.n672 B.n32 585
R789 B.n670 B.n669 585
R790 B.n671 B.n670 585
R791 B.n668 B.n37 585
R792 B.n37 B.n36 585
R793 B.n667 B.n666 585
R794 B.n666 B.n665 585
R795 B.n39 B.n38 585
R796 B.n664 B.n39 585
R797 B.n662 B.n661 585
R798 B.n663 B.n662 585
R799 B.n660 B.n44 585
R800 B.n44 B.n43 585
R801 B.n659 B.n658 585
R802 B.n658 B.n657 585
R803 B.n46 B.n45 585
R804 B.n656 B.n46 585
R805 B.n654 B.n653 585
R806 B.n655 B.n654 585
R807 B.n652 B.n51 585
R808 B.n51 B.n50 585
R809 B.n651 B.n650 585
R810 B.n650 B.n649 585
R811 B.n53 B.n52 585
R812 B.n648 B.n53 585
R813 B.n646 B.n645 585
R814 B.n647 B.n646 585
R815 B.n644 B.n58 585
R816 B.n58 B.n57 585
R817 B.n643 B.n642 585
R818 B.n642 B.n641 585
R819 B.n60 B.n59 585
R820 B.n640 B.n60 585
R821 B.n638 B.n637 585
R822 B.n639 B.n638 585
R823 B.n636 B.n65 585
R824 B.n65 B.n64 585
R825 B.n635 B.n634 585
R826 B.n634 B.n633 585
R827 B.n67 B.n66 585
R828 B.n632 B.n67 585
R829 B.n630 B.n629 585
R830 B.n631 B.n630 585
R831 B.n707 B.n706 585
R832 B.n706 B.n705 585
R833 B.n343 B.n184 497.305
R834 B.n630 B.n72 497.305
R835 B.n345 B.n182 497.305
R836 B.n506 B.n70 497.305
R837 B.n206 B.t13 279.603
R838 B.n199 B.t17 279.603
R839 B.n85 B.t6 279.603
R840 B.n93 B.t10 279.603
R841 B.n505 B.n71 256.663
R842 B.n511 B.n71 256.663
R843 B.n513 B.n71 256.663
R844 B.n519 B.n71 256.663
R845 B.n521 B.n71 256.663
R846 B.n527 B.n71 256.663
R847 B.n529 B.n71 256.663
R848 B.n535 B.n71 256.663
R849 B.n537 B.n71 256.663
R850 B.n543 B.n71 256.663
R851 B.n545 B.n71 256.663
R852 B.n551 B.n71 256.663
R853 B.n96 B.n71 256.663
R854 B.n557 B.n71 256.663
R855 B.n563 B.n71 256.663
R856 B.n565 B.n71 256.663
R857 B.n571 B.n71 256.663
R858 B.n88 B.n71 256.663
R859 B.n577 B.n71 256.663
R860 B.n583 B.n71 256.663
R861 B.n585 B.n71 256.663
R862 B.n591 B.n71 256.663
R863 B.n593 B.n71 256.663
R864 B.n599 B.n71 256.663
R865 B.n601 B.n71 256.663
R866 B.n607 B.n71 256.663
R867 B.n609 B.n71 256.663
R868 B.n615 B.n71 256.663
R869 B.n617 B.n71 256.663
R870 B.n623 B.n71 256.663
R871 B.n625 B.n71 256.663
R872 B.n338 B.n183 256.663
R873 B.n186 B.n183 256.663
R874 B.n331 B.n183 256.663
R875 B.n325 B.n183 256.663
R876 B.n323 B.n183 256.663
R877 B.n317 B.n183 256.663
R878 B.n315 B.n183 256.663
R879 B.n309 B.n183 256.663
R880 B.n307 B.n183 256.663
R881 B.n301 B.n183 256.663
R882 B.n299 B.n183 256.663
R883 B.n293 B.n183 256.663
R884 B.n291 B.n183 256.663
R885 B.n285 B.n183 256.663
R886 B.n283 B.n183 256.663
R887 B.n277 B.n183 256.663
R888 B.n275 B.n183 256.663
R889 B.n268 B.n183 256.663
R890 B.n266 B.n183 256.663
R891 B.n260 B.n183 256.663
R892 B.n258 B.n183 256.663
R893 B.n252 B.n183 256.663
R894 B.n250 B.n183 256.663
R895 B.n244 B.n183 256.663
R896 B.n242 B.n183 256.663
R897 B.n236 B.n183 256.663
R898 B.n234 B.n183 256.663
R899 B.n228 B.n183 256.663
R900 B.n226 B.n183 256.663
R901 B.n220 B.n183 256.663
R902 B.n206 B.t16 240.314
R903 B.n93 B.t11 240.314
R904 B.n199 B.t19 240.314
R905 B.n85 B.t8 240.314
R906 B.n207 B.t15 190.665
R907 B.n94 B.t12 190.665
R908 B.n200 B.t18 190.665
R909 B.n86 B.t9 190.665
R910 B.n343 B.n178 163.367
R911 B.n351 B.n178 163.367
R912 B.n351 B.n176 163.367
R913 B.n355 B.n176 163.367
R914 B.n355 B.n170 163.367
R915 B.n363 B.n170 163.367
R916 B.n363 B.n168 163.367
R917 B.n367 B.n168 163.367
R918 B.n367 B.n162 163.367
R919 B.n375 B.n162 163.367
R920 B.n375 B.n160 163.367
R921 B.n379 B.n160 163.367
R922 B.n379 B.n154 163.367
R923 B.n387 B.n154 163.367
R924 B.n387 B.n152 163.367
R925 B.n391 B.n152 163.367
R926 B.n391 B.n146 163.367
R927 B.n399 B.n146 163.367
R928 B.n399 B.n144 163.367
R929 B.n403 B.n144 163.367
R930 B.n403 B.n138 163.367
R931 B.n411 B.n138 163.367
R932 B.n411 B.n136 163.367
R933 B.n415 B.n136 163.367
R934 B.n415 B.n130 163.367
R935 B.n423 B.n130 163.367
R936 B.n423 B.n128 163.367
R937 B.n427 B.n128 163.367
R938 B.n427 B.n122 163.367
R939 B.n435 B.n122 163.367
R940 B.n435 B.n120 163.367
R941 B.n439 B.n120 163.367
R942 B.n439 B.n114 163.367
R943 B.n448 B.n114 163.367
R944 B.n448 B.n112 163.367
R945 B.n452 B.n112 163.367
R946 B.n452 B.n2 163.367
R947 B.n706 B.n2 163.367
R948 B.n706 B.n3 163.367
R949 B.n702 B.n3 163.367
R950 B.n702 B.n9 163.367
R951 B.n698 B.n9 163.367
R952 B.n698 B.n11 163.367
R953 B.n694 B.n11 163.367
R954 B.n694 B.n16 163.367
R955 B.n690 B.n16 163.367
R956 B.n690 B.n18 163.367
R957 B.n686 B.n18 163.367
R958 B.n686 B.n23 163.367
R959 B.n682 B.n23 163.367
R960 B.n682 B.n25 163.367
R961 B.n678 B.n25 163.367
R962 B.n678 B.n30 163.367
R963 B.n674 B.n30 163.367
R964 B.n674 B.n32 163.367
R965 B.n670 B.n32 163.367
R966 B.n670 B.n37 163.367
R967 B.n666 B.n37 163.367
R968 B.n666 B.n39 163.367
R969 B.n662 B.n39 163.367
R970 B.n662 B.n44 163.367
R971 B.n658 B.n44 163.367
R972 B.n658 B.n46 163.367
R973 B.n654 B.n46 163.367
R974 B.n654 B.n51 163.367
R975 B.n650 B.n51 163.367
R976 B.n650 B.n53 163.367
R977 B.n646 B.n53 163.367
R978 B.n646 B.n58 163.367
R979 B.n642 B.n58 163.367
R980 B.n642 B.n60 163.367
R981 B.n638 B.n60 163.367
R982 B.n638 B.n65 163.367
R983 B.n634 B.n65 163.367
R984 B.n634 B.n67 163.367
R985 B.n630 B.n67 163.367
R986 B.n339 B.n337 163.367
R987 B.n337 B.n336 163.367
R988 B.n333 B.n332 163.367
R989 B.n330 B.n188 163.367
R990 B.n326 B.n324 163.367
R991 B.n322 B.n190 163.367
R992 B.n318 B.n316 163.367
R993 B.n314 B.n192 163.367
R994 B.n310 B.n308 163.367
R995 B.n306 B.n194 163.367
R996 B.n302 B.n300 163.367
R997 B.n298 B.n196 163.367
R998 B.n294 B.n292 163.367
R999 B.n290 B.n198 163.367
R1000 B.n286 B.n284 163.367
R1001 B.n282 B.n203 163.367
R1002 B.n278 B.n276 163.367
R1003 B.n274 B.n205 163.367
R1004 B.n269 B.n267 163.367
R1005 B.n265 B.n209 163.367
R1006 B.n261 B.n259 163.367
R1007 B.n257 B.n211 163.367
R1008 B.n253 B.n251 163.367
R1009 B.n249 B.n213 163.367
R1010 B.n245 B.n243 163.367
R1011 B.n241 B.n215 163.367
R1012 B.n237 B.n235 163.367
R1013 B.n233 B.n217 163.367
R1014 B.n229 B.n227 163.367
R1015 B.n225 B.n219 163.367
R1016 B.n221 B.n182 163.367
R1017 B.n345 B.n180 163.367
R1018 B.n349 B.n180 163.367
R1019 B.n349 B.n174 163.367
R1020 B.n357 B.n174 163.367
R1021 B.n357 B.n172 163.367
R1022 B.n361 B.n172 163.367
R1023 B.n361 B.n166 163.367
R1024 B.n369 B.n166 163.367
R1025 B.n369 B.n164 163.367
R1026 B.n373 B.n164 163.367
R1027 B.n373 B.n158 163.367
R1028 B.n381 B.n158 163.367
R1029 B.n381 B.n156 163.367
R1030 B.n385 B.n156 163.367
R1031 B.n385 B.n149 163.367
R1032 B.n393 B.n149 163.367
R1033 B.n393 B.n147 163.367
R1034 B.n397 B.n147 163.367
R1035 B.n397 B.n142 163.367
R1036 B.n405 B.n142 163.367
R1037 B.n405 B.n140 163.367
R1038 B.n409 B.n140 163.367
R1039 B.n409 B.n133 163.367
R1040 B.n417 B.n133 163.367
R1041 B.n417 B.n131 163.367
R1042 B.n421 B.n131 163.367
R1043 B.n421 B.n126 163.367
R1044 B.n429 B.n126 163.367
R1045 B.n429 B.n124 163.367
R1046 B.n433 B.n124 163.367
R1047 B.n433 B.n118 163.367
R1048 B.n441 B.n118 163.367
R1049 B.n441 B.n116 163.367
R1050 B.n446 B.n116 163.367
R1051 B.n446 B.n110 163.367
R1052 B.n454 B.n110 163.367
R1053 B.n455 B.n454 163.367
R1054 B.n455 B.n5 163.367
R1055 B.n6 B.n5 163.367
R1056 B.n7 B.n6 163.367
R1057 B.n460 B.n7 163.367
R1058 B.n460 B.n12 163.367
R1059 B.n13 B.n12 163.367
R1060 B.n14 B.n13 163.367
R1061 B.n465 B.n14 163.367
R1062 B.n465 B.n19 163.367
R1063 B.n20 B.n19 163.367
R1064 B.n21 B.n20 163.367
R1065 B.n470 B.n21 163.367
R1066 B.n470 B.n26 163.367
R1067 B.n27 B.n26 163.367
R1068 B.n28 B.n27 163.367
R1069 B.n475 B.n28 163.367
R1070 B.n475 B.n33 163.367
R1071 B.n34 B.n33 163.367
R1072 B.n35 B.n34 163.367
R1073 B.n480 B.n35 163.367
R1074 B.n480 B.n40 163.367
R1075 B.n41 B.n40 163.367
R1076 B.n42 B.n41 163.367
R1077 B.n485 B.n42 163.367
R1078 B.n485 B.n47 163.367
R1079 B.n48 B.n47 163.367
R1080 B.n49 B.n48 163.367
R1081 B.n490 B.n49 163.367
R1082 B.n490 B.n54 163.367
R1083 B.n55 B.n54 163.367
R1084 B.n56 B.n55 163.367
R1085 B.n495 B.n56 163.367
R1086 B.n495 B.n61 163.367
R1087 B.n62 B.n61 163.367
R1088 B.n63 B.n62 163.367
R1089 B.n500 B.n63 163.367
R1090 B.n500 B.n68 163.367
R1091 B.n69 B.n68 163.367
R1092 B.n70 B.n69 163.367
R1093 B.n626 B.n624 163.367
R1094 B.n622 B.n74 163.367
R1095 B.n618 B.n616 163.367
R1096 B.n614 B.n76 163.367
R1097 B.n610 B.n608 163.367
R1098 B.n606 B.n78 163.367
R1099 B.n602 B.n600 163.367
R1100 B.n598 B.n80 163.367
R1101 B.n594 B.n592 163.367
R1102 B.n590 B.n82 163.367
R1103 B.n586 B.n584 163.367
R1104 B.n582 B.n84 163.367
R1105 B.n578 B.n576 163.367
R1106 B.n573 B.n572 163.367
R1107 B.n570 B.n90 163.367
R1108 B.n566 B.n564 163.367
R1109 B.n562 B.n92 163.367
R1110 B.n558 B.n556 163.367
R1111 B.n553 B.n552 163.367
R1112 B.n550 B.n98 163.367
R1113 B.n546 B.n544 163.367
R1114 B.n542 B.n100 163.367
R1115 B.n538 B.n536 163.367
R1116 B.n534 B.n102 163.367
R1117 B.n530 B.n528 163.367
R1118 B.n526 B.n104 163.367
R1119 B.n522 B.n520 163.367
R1120 B.n518 B.n106 163.367
R1121 B.n514 B.n512 163.367
R1122 B.n510 B.n108 163.367
R1123 B.n344 B.n183 127.897
R1124 B.n631 B.n71 127.897
R1125 B.n338 B.n184 71.676
R1126 B.n336 B.n186 71.676
R1127 B.n332 B.n331 71.676
R1128 B.n325 B.n188 71.676
R1129 B.n324 B.n323 71.676
R1130 B.n317 B.n190 71.676
R1131 B.n316 B.n315 71.676
R1132 B.n309 B.n192 71.676
R1133 B.n308 B.n307 71.676
R1134 B.n301 B.n194 71.676
R1135 B.n300 B.n299 71.676
R1136 B.n293 B.n196 71.676
R1137 B.n292 B.n291 71.676
R1138 B.n285 B.n198 71.676
R1139 B.n284 B.n283 71.676
R1140 B.n277 B.n203 71.676
R1141 B.n276 B.n275 71.676
R1142 B.n268 B.n205 71.676
R1143 B.n267 B.n266 71.676
R1144 B.n260 B.n209 71.676
R1145 B.n259 B.n258 71.676
R1146 B.n252 B.n211 71.676
R1147 B.n251 B.n250 71.676
R1148 B.n244 B.n213 71.676
R1149 B.n243 B.n242 71.676
R1150 B.n236 B.n215 71.676
R1151 B.n235 B.n234 71.676
R1152 B.n228 B.n217 71.676
R1153 B.n227 B.n226 71.676
R1154 B.n220 B.n219 71.676
R1155 B.n625 B.n72 71.676
R1156 B.n624 B.n623 71.676
R1157 B.n617 B.n74 71.676
R1158 B.n616 B.n615 71.676
R1159 B.n609 B.n76 71.676
R1160 B.n608 B.n607 71.676
R1161 B.n601 B.n78 71.676
R1162 B.n600 B.n599 71.676
R1163 B.n593 B.n80 71.676
R1164 B.n592 B.n591 71.676
R1165 B.n585 B.n82 71.676
R1166 B.n584 B.n583 71.676
R1167 B.n577 B.n84 71.676
R1168 B.n576 B.n88 71.676
R1169 B.n572 B.n571 71.676
R1170 B.n565 B.n90 71.676
R1171 B.n564 B.n563 71.676
R1172 B.n557 B.n92 71.676
R1173 B.n556 B.n96 71.676
R1174 B.n552 B.n551 71.676
R1175 B.n545 B.n98 71.676
R1176 B.n544 B.n543 71.676
R1177 B.n537 B.n100 71.676
R1178 B.n536 B.n535 71.676
R1179 B.n529 B.n102 71.676
R1180 B.n528 B.n527 71.676
R1181 B.n521 B.n104 71.676
R1182 B.n520 B.n519 71.676
R1183 B.n513 B.n106 71.676
R1184 B.n512 B.n511 71.676
R1185 B.n505 B.n108 71.676
R1186 B.n506 B.n505 71.676
R1187 B.n511 B.n510 71.676
R1188 B.n514 B.n513 71.676
R1189 B.n519 B.n518 71.676
R1190 B.n522 B.n521 71.676
R1191 B.n527 B.n526 71.676
R1192 B.n530 B.n529 71.676
R1193 B.n535 B.n534 71.676
R1194 B.n538 B.n537 71.676
R1195 B.n543 B.n542 71.676
R1196 B.n546 B.n545 71.676
R1197 B.n551 B.n550 71.676
R1198 B.n553 B.n96 71.676
R1199 B.n558 B.n557 71.676
R1200 B.n563 B.n562 71.676
R1201 B.n566 B.n565 71.676
R1202 B.n571 B.n570 71.676
R1203 B.n573 B.n88 71.676
R1204 B.n578 B.n577 71.676
R1205 B.n583 B.n582 71.676
R1206 B.n586 B.n585 71.676
R1207 B.n591 B.n590 71.676
R1208 B.n594 B.n593 71.676
R1209 B.n599 B.n598 71.676
R1210 B.n602 B.n601 71.676
R1211 B.n607 B.n606 71.676
R1212 B.n610 B.n609 71.676
R1213 B.n615 B.n614 71.676
R1214 B.n618 B.n617 71.676
R1215 B.n623 B.n622 71.676
R1216 B.n626 B.n625 71.676
R1217 B.n339 B.n338 71.676
R1218 B.n333 B.n186 71.676
R1219 B.n331 B.n330 71.676
R1220 B.n326 B.n325 71.676
R1221 B.n323 B.n322 71.676
R1222 B.n318 B.n317 71.676
R1223 B.n315 B.n314 71.676
R1224 B.n310 B.n309 71.676
R1225 B.n307 B.n306 71.676
R1226 B.n302 B.n301 71.676
R1227 B.n299 B.n298 71.676
R1228 B.n294 B.n293 71.676
R1229 B.n291 B.n290 71.676
R1230 B.n286 B.n285 71.676
R1231 B.n283 B.n282 71.676
R1232 B.n278 B.n277 71.676
R1233 B.n275 B.n274 71.676
R1234 B.n269 B.n268 71.676
R1235 B.n266 B.n265 71.676
R1236 B.n261 B.n260 71.676
R1237 B.n258 B.n257 71.676
R1238 B.n253 B.n252 71.676
R1239 B.n250 B.n249 71.676
R1240 B.n245 B.n244 71.676
R1241 B.n242 B.n241 71.676
R1242 B.n237 B.n236 71.676
R1243 B.n234 B.n233 71.676
R1244 B.n229 B.n228 71.676
R1245 B.n226 B.n225 71.676
R1246 B.n221 B.n220 71.676
R1247 B.n344 B.n179 62.5685
R1248 B.n350 B.n179 62.5685
R1249 B.n350 B.n175 62.5685
R1250 B.n356 B.n175 62.5685
R1251 B.n356 B.n171 62.5685
R1252 B.n362 B.n171 62.5685
R1253 B.n368 B.n167 62.5685
R1254 B.n368 B.n163 62.5685
R1255 B.n374 B.n163 62.5685
R1256 B.n374 B.n159 62.5685
R1257 B.n380 B.n159 62.5685
R1258 B.n380 B.n155 62.5685
R1259 B.n386 B.n155 62.5685
R1260 B.n386 B.n150 62.5685
R1261 B.n392 B.n150 62.5685
R1262 B.n392 B.n151 62.5685
R1263 B.n398 B.n143 62.5685
R1264 B.n404 B.n143 62.5685
R1265 B.n404 B.n139 62.5685
R1266 B.n410 B.n139 62.5685
R1267 B.n410 B.n134 62.5685
R1268 B.n416 B.n134 62.5685
R1269 B.n416 B.n135 62.5685
R1270 B.n422 B.n127 62.5685
R1271 B.n428 B.n127 62.5685
R1272 B.n428 B.n123 62.5685
R1273 B.n434 B.n123 62.5685
R1274 B.n434 B.n119 62.5685
R1275 B.n440 B.n119 62.5685
R1276 B.n447 B.n115 62.5685
R1277 B.n447 B.n111 62.5685
R1278 B.n453 B.n111 62.5685
R1279 B.n453 B.n4 62.5685
R1280 B.n705 B.n4 62.5685
R1281 B.n705 B.n704 62.5685
R1282 B.n704 B.n703 62.5685
R1283 B.n703 B.n8 62.5685
R1284 B.n697 B.n8 62.5685
R1285 B.n697 B.n696 62.5685
R1286 B.n695 B.n15 62.5685
R1287 B.n689 B.n15 62.5685
R1288 B.n689 B.n688 62.5685
R1289 B.n688 B.n687 62.5685
R1290 B.n687 B.n22 62.5685
R1291 B.n681 B.n22 62.5685
R1292 B.n680 B.n679 62.5685
R1293 B.n679 B.n29 62.5685
R1294 B.n673 B.n29 62.5685
R1295 B.n673 B.n672 62.5685
R1296 B.n672 B.n671 62.5685
R1297 B.n671 B.n36 62.5685
R1298 B.n665 B.n36 62.5685
R1299 B.n664 B.n663 62.5685
R1300 B.n663 B.n43 62.5685
R1301 B.n657 B.n43 62.5685
R1302 B.n657 B.n656 62.5685
R1303 B.n656 B.n655 62.5685
R1304 B.n655 B.n50 62.5685
R1305 B.n649 B.n50 62.5685
R1306 B.n649 B.n648 62.5685
R1307 B.n648 B.n647 62.5685
R1308 B.n647 B.n57 62.5685
R1309 B.n641 B.n640 62.5685
R1310 B.n640 B.n639 62.5685
R1311 B.n639 B.n64 62.5685
R1312 B.n633 B.n64 62.5685
R1313 B.n633 B.n632 62.5685
R1314 B.n632 B.n631 62.5685
R1315 B.n271 B.n207 59.5399
R1316 B.n201 B.n200 59.5399
R1317 B.n87 B.n86 59.5399
R1318 B.n95 B.n94 59.5399
R1319 B.n422 B.t5 56.1276
R1320 B.n681 B.t1 56.1276
R1321 B.n362 B.t14 52.4472
R1322 B.n641 B.t7 52.4472
R1323 B.n207 B.n206 49.649
R1324 B.n200 B.n199 49.649
R1325 B.n86 B.n85 49.649
R1326 B.n94 B.n93 49.649
R1327 B.n440 B.t0 39.5655
R1328 B.t2 B.n695 39.5655
R1329 B.n151 B.t3 35.8851
R1330 B.t4 B.n664 35.8851
R1331 B.n629 B.n628 32.3127
R1332 B.n507 B.n504 32.3127
R1333 B.n346 B.n181 32.3127
R1334 B.n342 B.n341 32.3127
R1335 B.n398 B.t3 26.6839
R1336 B.n665 B.t4 26.6839
R1337 B.t0 B.n115 23.0034
R1338 B.n696 B.t2 23.0034
R1339 B B.n707 18.0485
R1340 B.n628 B.n627 10.6151
R1341 B.n627 B.n73 10.6151
R1342 B.n621 B.n73 10.6151
R1343 B.n621 B.n620 10.6151
R1344 B.n620 B.n619 10.6151
R1345 B.n619 B.n75 10.6151
R1346 B.n613 B.n75 10.6151
R1347 B.n613 B.n612 10.6151
R1348 B.n612 B.n611 10.6151
R1349 B.n611 B.n77 10.6151
R1350 B.n605 B.n77 10.6151
R1351 B.n605 B.n604 10.6151
R1352 B.n604 B.n603 10.6151
R1353 B.n603 B.n79 10.6151
R1354 B.n597 B.n79 10.6151
R1355 B.n597 B.n596 10.6151
R1356 B.n596 B.n595 10.6151
R1357 B.n595 B.n81 10.6151
R1358 B.n589 B.n81 10.6151
R1359 B.n589 B.n588 10.6151
R1360 B.n588 B.n587 10.6151
R1361 B.n587 B.n83 10.6151
R1362 B.n581 B.n83 10.6151
R1363 B.n581 B.n580 10.6151
R1364 B.n580 B.n579 10.6151
R1365 B.n575 B.n574 10.6151
R1366 B.n574 B.n89 10.6151
R1367 B.n569 B.n89 10.6151
R1368 B.n569 B.n568 10.6151
R1369 B.n568 B.n567 10.6151
R1370 B.n567 B.n91 10.6151
R1371 B.n561 B.n91 10.6151
R1372 B.n561 B.n560 10.6151
R1373 B.n560 B.n559 10.6151
R1374 B.n555 B.n554 10.6151
R1375 B.n554 B.n97 10.6151
R1376 B.n549 B.n97 10.6151
R1377 B.n549 B.n548 10.6151
R1378 B.n548 B.n547 10.6151
R1379 B.n547 B.n99 10.6151
R1380 B.n541 B.n99 10.6151
R1381 B.n541 B.n540 10.6151
R1382 B.n540 B.n539 10.6151
R1383 B.n539 B.n101 10.6151
R1384 B.n533 B.n101 10.6151
R1385 B.n533 B.n532 10.6151
R1386 B.n532 B.n531 10.6151
R1387 B.n531 B.n103 10.6151
R1388 B.n525 B.n103 10.6151
R1389 B.n525 B.n524 10.6151
R1390 B.n524 B.n523 10.6151
R1391 B.n523 B.n105 10.6151
R1392 B.n517 B.n105 10.6151
R1393 B.n517 B.n516 10.6151
R1394 B.n516 B.n515 10.6151
R1395 B.n515 B.n107 10.6151
R1396 B.n509 B.n107 10.6151
R1397 B.n509 B.n508 10.6151
R1398 B.n508 B.n507 10.6151
R1399 B.n347 B.n346 10.6151
R1400 B.n348 B.n347 10.6151
R1401 B.n348 B.n173 10.6151
R1402 B.n358 B.n173 10.6151
R1403 B.n359 B.n358 10.6151
R1404 B.n360 B.n359 10.6151
R1405 B.n360 B.n165 10.6151
R1406 B.n370 B.n165 10.6151
R1407 B.n371 B.n370 10.6151
R1408 B.n372 B.n371 10.6151
R1409 B.n372 B.n157 10.6151
R1410 B.n382 B.n157 10.6151
R1411 B.n383 B.n382 10.6151
R1412 B.n384 B.n383 10.6151
R1413 B.n384 B.n148 10.6151
R1414 B.n394 B.n148 10.6151
R1415 B.n395 B.n394 10.6151
R1416 B.n396 B.n395 10.6151
R1417 B.n396 B.n141 10.6151
R1418 B.n406 B.n141 10.6151
R1419 B.n407 B.n406 10.6151
R1420 B.n408 B.n407 10.6151
R1421 B.n408 B.n132 10.6151
R1422 B.n418 B.n132 10.6151
R1423 B.n419 B.n418 10.6151
R1424 B.n420 B.n419 10.6151
R1425 B.n420 B.n125 10.6151
R1426 B.n430 B.n125 10.6151
R1427 B.n431 B.n430 10.6151
R1428 B.n432 B.n431 10.6151
R1429 B.n432 B.n117 10.6151
R1430 B.n442 B.n117 10.6151
R1431 B.n443 B.n442 10.6151
R1432 B.n445 B.n443 10.6151
R1433 B.n445 B.n444 10.6151
R1434 B.n444 B.n109 10.6151
R1435 B.n456 B.n109 10.6151
R1436 B.n457 B.n456 10.6151
R1437 B.n458 B.n457 10.6151
R1438 B.n459 B.n458 10.6151
R1439 B.n461 B.n459 10.6151
R1440 B.n462 B.n461 10.6151
R1441 B.n463 B.n462 10.6151
R1442 B.n464 B.n463 10.6151
R1443 B.n466 B.n464 10.6151
R1444 B.n467 B.n466 10.6151
R1445 B.n468 B.n467 10.6151
R1446 B.n469 B.n468 10.6151
R1447 B.n471 B.n469 10.6151
R1448 B.n472 B.n471 10.6151
R1449 B.n473 B.n472 10.6151
R1450 B.n474 B.n473 10.6151
R1451 B.n476 B.n474 10.6151
R1452 B.n477 B.n476 10.6151
R1453 B.n478 B.n477 10.6151
R1454 B.n479 B.n478 10.6151
R1455 B.n481 B.n479 10.6151
R1456 B.n482 B.n481 10.6151
R1457 B.n483 B.n482 10.6151
R1458 B.n484 B.n483 10.6151
R1459 B.n486 B.n484 10.6151
R1460 B.n487 B.n486 10.6151
R1461 B.n488 B.n487 10.6151
R1462 B.n489 B.n488 10.6151
R1463 B.n491 B.n489 10.6151
R1464 B.n492 B.n491 10.6151
R1465 B.n493 B.n492 10.6151
R1466 B.n494 B.n493 10.6151
R1467 B.n496 B.n494 10.6151
R1468 B.n497 B.n496 10.6151
R1469 B.n498 B.n497 10.6151
R1470 B.n499 B.n498 10.6151
R1471 B.n501 B.n499 10.6151
R1472 B.n502 B.n501 10.6151
R1473 B.n503 B.n502 10.6151
R1474 B.n504 B.n503 10.6151
R1475 B.n341 B.n340 10.6151
R1476 B.n340 B.n185 10.6151
R1477 B.n335 B.n185 10.6151
R1478 B.n335 B.n334 10.6151
R1479 B.n334 B.n187 10.6151
R1480 B.n329 B.n187 10.6151
R1481 B.n329 B.n328 10.6151
R1482 B.n328 B.n327 10.6151
R1483 B.n327 B.n189 10.6151
R1484 B.n321 B.n189 10.6151
R1485 B.n321 B.n320 10.6151
R1486 B.n320 B.n319 10.6151
R1487 B.n319 B.n191 10.6151
R1488 B.n313 B.n191 10.6151
R1489 B.n313 B.n312 10.6151
R1490 B.n312 B.n311 10.6151
R1491 B.n311 B.n193 10.6151
R1492 B.n305 B.n193 10.6151
R1493 B.n305 B.n304 10.6151
R1494 B.n304 B.n303 10.6151
R1495 B.n303 B.n195 10.6151
R1496 B.n297 B.n195 10.6151
R1497 B.n297 B.n296 10.6151
R1498 B.n296 B.n295 10.6151
R1499 B.n295 B.n197 10.6151
R1500 B.n289 B.n288 10.6151
R1501 B.n288 B.n287 10.6151
R1502 B.n287 B.n202 10.6151
R1503 B.n281 B.n202 10.6151
R1504 B.n281 B.n280 10.6151
R1505 B.n280 B.n279 10.6151
R1506 B.n279 B.n204 10.6151
R1507 B.n273 B.n204 10.6151
R1508 B.n273 B.n272 10.6151
R1509 B.n270 B.n208 10.6151
R1510 B.n264 B.n208 10.6151
R1511 B.n264 B.n263 10.6151
R1512 B.n263 B.n262 10.6151
R1513 B.n262 B.n210 10.6151
R1514 B.n256 B.n210 10.6151
R1515 B.n256 B.n255 10.6151
R1516 B.n255 B.n254 10.6151
R1517 B.n254 B.n212 10.6151
R1518 B.n248 B.n212 10.6151
R1519 B.n248 B.n247 10.6151
R1520 B.n247 B.n246 10.6151
R1521 B.n246 B.n214 10.6151
R1522 B.n240 B.n214 10.6151
R1523 B.n240 B.n239 10.6151
R1524 B.n239 B.n238 10.6151
R1525 B.n238 B.n216 10.6151
R1526 B.n232 B.n216 10.6151
R1527 B.n232 B.n231 10.6151
R1528 B.n231 B.n230 10.6151
R1529 B.n230 B.n218 10.6151
R1530 B.n224 B.n218 10.6151
R1531 B.n224 B.n223 10.6151
R1532 B.n223 B.n222 10.6151
R1533 B.n222 B.n181 10.6151
R1534 B.n342 B.n177 10.6151
R1535 B.n352 B.n177 10.6151
R1536 B.n353 B.n352 10.6151
R1537 B.n354 B.n353 10.6151
R1538 B.n354 B.n169 10.6151
R1539 B.n364 B.n169 10.6151
R1540 B.n365 B.n364 10.6151
R1541 B.n366 B.n365 10.6151
R1542 B.n366 B.n161 10.6151
R1543 B.n376 B.n161 10.6151
R1544 B.n377 B.n376 10.6151
R1545 B.n378 B.n377 10.6151
R1546 B.n378 B.n153 10.6151
R1547 B.n388 B.n153 10.6151
R1548 B.n389 B.n388 10.6151
R1549 B.n390 B.n389 10.6151
R1550 B.n390 B.n145 10.6151
R1551 B.n400 B.n145 10.6151
R1552 B.n401 B.n400 10.6151
R1553 B.n402 B.n401 10.6151
R1554 B.n402 B.n137 10.6151
R1555 B.n412 B.n137 10.6151
R1556 B.n413 B.n412 10.6151
R1557 B.n414 B.n413 10.6151
R1558 B.n414 B.n129 10.6151
R1559 B.n424 B.n129 10.6151
R1560 B.n425 B.n424 10.6151
R1561 B.n426 B.n425 10.6151
R1562 B.n426 B.n121 10.6151
R1563 B.n436 B.n121 10.6151
R1564 B.n437 B.n436 10.6151
R1565 B.n438 B.n437 10.6151
R1566 B.n438 B.n113 10.6151
R1567 B.n449 B.n113 10.6151
R1568 B.n450 B.n449 10.6151
R1569 B.n451 B.n450 10.6151
R1570 B.n451 B.n0 10.6151
R1571 B.n701 B.n1 10.6151
R1572 B.n701 B.n700 10.6151
R1573 B.n700 B.n699 10.6151
R1574 B.n699 B.n10 10.6151
R1575 B.n693 B.n10 10.6151
R1576 B.n693 B.n692 10.6151
R1577 B.n692 B.n691 10.6151
R1578 B.n691 B.n17 10.6151
R1579 B.n685 B.n17 10.6151
R1580 B.n685 B.n684 10.6151
R1581 B.n684 B.n683 10.6151
R1582 B.n683 B.n24 10.6151
R1583 B.n677 B.n24 10.6151
R1584 B.n677 B.n676 10.6151
R1585 B.n676 B.n675 10.6151
R1586 B.n675 B.n31 10.6151
R1587 B.n669 B.n31 10.6151
R1588 B.n669 B.n668 10.6151
R1589 B.n668 B.n667 10.6151
R1590 B.n667 B.n38 10.6151
R1591 B.n661 B.n38 10.6151
R1592 B.n661 B.n660 10.6151
R1593 B.n660 B.n659 10.6151
R1594 B.n659 B.n45 10.6151
R1595 B.n653 B.n45 10.6151
R1596 B.n653 B.n652 10.6151
R1597 B.n652 B.n651 10.6151
R1598 B.n651 B.n52 10.6151
R1599 B.n645 B.n52 10.6151
R1600 B.n645 B.n644 10.6151
R1601 B.n644 B.n643 10.6151
R1602 B.n643 B.n59 10.6151
R1603 B.n637 B.n59 10.6151
R1604 B.n637 B.n636 10.6151
R1605 B.n636 B.n635 10.6151
R1606 B.n635 B.n66 10.6151
R1607 B.n629 B.n66 10.6151
R1608 B.t14 B.n167 10.1218
R1609 B.t7 B.n57 10.1218
R1610 B.n579 B.n87 9.36635
R1611 B.n555 B.n95 9.36635
R1612 B.n201 B.n197 9.36635
R1613 B.n271 B.n270 9.36635
R1614 B.n135 B.t5 6.44132
R1615 B.t1 B.n680 6.44132
R1616 B.n707 B.n0 2.81026
R1617 B.n707 B.n1 2.81026
R1618 B.n575 B.n87 1.24928
R1619 B.n559 B.n95 1.24928
R1620 B.n289 B.n201 1.24928
R1621 B.n272 B.n271 1.24928
R1622 VP.n11 VP.n8 161.3
R1623 VP.n13 VP.n12 161.3
R1624 VP.n14 VP.n7 161.3
R1625 VP.n16 VP.n15 161.3
R1626 VP.n17 VP.n6 161.3
R1627 VP.n36 VP.n0 161.3
R1628 VP.n35 VP.n34 161.3
R1629 VP.n33 VP.n1 161.3
R1630 VP.n32 VP.n31 161.3
R1631 VP.n30 VP.n2 161.3
R1632 VP.n28 VP.n27 161.3
R1633 VP.n26 VP.n3 161.3
R1634 VP.n25 VP.n24 161.3
R1635 VP.n23 VP.n4 161.3
R1636 VP.n22 VP.n21 161.3
R1637 VP.n9 VP.t1 105.103
R1638 VP.n20 VP.n5 95.6613
R1639 VP.n38 VP.n37 95.6613
R1640 VP.n19 VP.n18 95.6613
R1641 VP.n5 VP.t3 72.1924
R1642 VP.n29 VP.t0 72.1924
R1643 VP.n37 VP.t2 72.1924
R1644 VP.n18 VP.t4 72.1924
R1645 VP.n10 VP.t5 72.1924
R1646 VP.n10 VP.n9 59.417
R1647 VP.n24 VP.n23 43.4833
R1648 VP.n35 VP.n1 43.4833
R1649 VP.n16 VP.n7 43.4833
R1650 VP.n20 VP.n19 43.2042
R1651 VP.n24 VP.n3 37.6707
R1652 VP.n31 VP.n1 37.6707
R1653 VP.n12 VP.n7 37.6707
R1654 VP.n23 VP.n22 24.5923
R1655 VP.n28 VP.n3 24.5923
R1656 VP.n31 VP.n30 24.5923
R1657 VP.n36 VP.n35 24.5923
R1658 VP.n17 VP.n16 24.5923
R1659 VP.n12 VP.n11 24.5923
R1660 VP.n22 VP.n5 15.2474
R1661 VP.n37 VP.n36 15.2474
R1662 VP.n18 VP.n17 15.2474
R1663 VP.n29 VP.n28 12.2964
R1664 VP.n30 VP.n29 12.2964
R1665 VP.n11 VP.n10 12.2964
R1666 VP.n9 VP.n8 9.41768
R1667 VP.n19 VP.n6 0.278335
R1668 VP.n21 VP.n20 0.278335
R1669 VP.n38 VP.n0 0.278335
R1670 VP.n13 VP.n8 0.189894
R1671 VP.n14 VP.n13 0.189894
R1672 VP.n15 VP.n14 0.189894
R1673 VP.n15 VP.n6 0.189894
R1674 VP.n21 VP.n4 0.189894
R1675 VP.n25 VP.n4 0.189894
R1676 VP.n26 VP.n25 0.189894
R1677 VP.n27 VP.n26 0.189894
R1678 VP.n27 VP.n2 0.189894
R1679 VP.n32 VP.n2 0.189894
R1680 VP.n33 VP.n32 0.189894
R1681 VP.n34 VP.n33 0.189894
R1682 VP.n34 VP.n0 0.189894
R1683 VP VP.n38 0.153485
R1684 VDD1.n30 VDD1.n0 289.615
R1685 VDD1.n65 VDD1.n35 289.615
R1686 VDD1.n31 VDD1.n30 185
R1687 VDD1.n29 VDD1.n28 185
R1688 VDD1.n4 VDD1.n3 185
R1689 VDD1.n23 VDD1.n22 185
R1690 VDD1.n21 VDD1.n20 185
R1691 VDD1.n8 VDD1.n7 185
R1692 VDD1.n15 VDD1.n14 185
R1693 VDD1.n13 VDD1.n12 185
R1694 VDD1.n48 VDD1.n47 185
R1695 VDD1.n50 VDD1.n49 185
R1696 VDD1.n43 VDD1.n42 185
R1697 VDD1.n56 VDD1.n55 185
R1698 VDD1.n58 VDD1.n57 185
R1699 VDD1.n39 VDD1.n38 185
R1700 VDD1.n64 VDD1.n63 185
R1701 VDD1.n66 VDD1.n65 185
R1702 VDD1.n11 VDD1.t4 147.659
R1703 VDD1.n46 VDD1.t2 147.659
R1704 VDD1.n30 VDD1.n29 104.615
R1705 VDD1.n29 VDD1.n3 104.615
R1706 VDD1.n22 VDD1.n3 104.615
R1707 VDD1.n22 VDD1.n21 104.615
R1708 VDD1.n21 VDD1.n7 104.615
R1709 VDD1.n14 VDD1.n7 104.615
R1710 VDD1.n14 VDD1.n13 104.615
R1711 VDD1.n49 VDD1.n48 104.615
R1712 VDD1.n49 VDD1.n42 104.615
R1713 VDD1.n56 VDD1.n42 104.615
R1714 VDD1.n57 VDD1.n56 104.615
R1715 VDD1.n57 VDD1.n38 104.615
R1716 VDD1.n64 VDD1.n38 104.615
R1717 VDD1.n65 VDD1.n64 104.615
R1718 VDD1.n71 VDD1.n70 65.7946
R1719 VDD1.n73 VDD1.n72 65.2982
R1720 VDD1.n13 VDD1.t4 52.3082
R1721 VDD1.n48 VDD1.t2 52.3082
R1722 VDD1 VDD1.n34 49.8017
R1723 VDD1.n71 VDD1.n69 49.6882
R1724 VDD1.n73 VDD1.n71 38.3328
R1725 VDD1.n12 VDD1.n11 15.6676
R1726 VDD1.n47 VDD1.n46 15.6676
R1727 VDD1.n15 VDD1.n10 12.8005
R1728 VDD1.n50 VDD1.n45 12.8005
R1729 VDD1.n16 VDD1.n8 12.0247
R1730 VDD1.n51 VDD1.n43 12.0247
R1731 VDD1.n20 VDD1.n19 11.249
R1732 VDD1.n55 VDD1.n54 11.249
R1733 VDD1.n23 VDD1.n6 10.4732
R1734 VDD1.n58 VDD1.n41 10.4732
R1735 VDD1.n24 VDD1.n4 9.69747
R1736 VDD1.n59 VDD1.n39 9.69747
R1737 VDD1.n34 VDD1.n33 9.45567
R1738 VDD1.n69 VDD1.n68 9.45567
R1739 VDD1.n33 VDD1.n32 9.3005
R1740 VDD1.n2 VDD1.n1 9.3005
R1741 VDD1.n27 VDD1.n26 9.3005
R1742 VDD1.n25 VDD1.n24 9.3005
R1743 VDD1.n6 VDD1.n5 9.3005
R1744 VDD1.n19 VDD1.n18 9.3005
R1745 VDD1.n17 VDD1.n16 9.3005
R1746 VDD1.n10 VDD1.n9 9.3005
R1747 VDD1.n37 VDD1.n36 9.3005
R1748 VDD1.n62 VDD1.n61 9.3005
R1749 VDD1.n60 VDD1.n59 9.3005
R1750 VDD1.n41 VDD1.n40 9.3005
R1751 VDD1.n54 VDD1.n53 9.3005
R1752 VDD1.n52 VDD1.n51 9.3005
R1753 VDD1.n45 VDD1.n44 9.3005
R1754 VDD1.n68 VDD1.n67 9.3005
R1755 VDD1.n28 VDD1.n27 8.92171
R1756 VDD1.n63 VDD1.n62 8.92171
R1757 VDD1.n31 VDD1.n2 8.14595
R1758 VDD1.n66 VDD1.n37 8.14595
R1759 VDD1.n32 VDD1.n0 7.3702
R1760 VDD1.n67 VDD1.n35 7.3702
R1761 VDD1.n34 VDD1.n0 6.59444
R1762 VDD1.n69 VDD1.n35 6.59444
R1763 VDD1.n32 VDD1.n31 5.81868
R1764 VDD1.n67 VDD1.n66 5.81868
R1765 VDD1.n28 VDD1.n2 5.04292
R1766 VDD1.n63 VDD1.n37 5.04292
R1767 VDD1.n11 VDD1.n9 4.38571
R1768 VDD1.n46 VDD1.n44 4.38571
R1769 VDD1.n27 VDD1.n4 4.26717
R1770 VDD1.n62 VDD1.n39 4.26717
R1771 VDD1.n24 VDD1.n23 3.49141
R1772 VDD1.n59 VDD1.n58 3.49141
R1773 VDD1.n72 VDD1.t0 2.96457
R1774 VDD1.n72 VDD1.t1 2.96457
R1775 VDD1.n70 VDD1.t5 2.96457
R1776 VDD1.n70 VDD1.t3 2.96457
R1777 VDD1.n20 VDD1.n6 2.71565
R1778 VDD1.n55 VDD1.n41 2.71565
R1779 VDD1.n19 VDD1.n8 1.93989
R1780 VDD1.n54 VDD1.n43 1.93989
R1781 VDD1.n16 VDD1.n15 1.16414
R1782 VDD1.n51 VDD1.n50 1.16414
R1783 VDD1 VDD1.n73 0.494034
R1784 VDD1.n12 VDD1.n10 0.388379
R1785 VDD1.n47 VDD1.n45 0.388379
R1786 VDD1.n33 VDD1.n1 0.155672
R1787 VDD1.n26 VDD1.n1 0.155672
R1788 VDD1.n26 VDD1.n25 0.155672
R1789 VDD1.n25 VDD1.n5 0.155672
R1790 VDD1.n18 VDD1.n5 0.155672
R1791 VDD1.n18 VDD1.n17 0.155672
R1792 VDD1.n17 VDD1.n9 0.155672
R1793 VDD1.n52 VDD1.n44 0.155672
R1794 VDD1.n53 VDD1.n52 0.155672
R1795 VDD1.n53 VDD1.n40 0.155672
R1796 VDD1.n60 VDD1.n40 0.155672
R1797 VDD1.n61 VDD1.n60 0.155672
R1798 VDD1.n61 VDD1.n36 0.155672
R1799 VDD1.n68 VDD1.n36 0.155672
C0 VN VDD2 3.80073f
C1 VP VDD1 4.07473f
C2 VTAIL VDD1 5.6533f
C3 VTAIL VP 4.23729f
C4 VN VDD1 0.150396f
C5 VP VN 5.57861f
C6 VTAIL VN 4.22307f
C7 VDD1 VDD2 1.261f
C8 VP VDD2 0.426659f
C9 VTAIL VDD2 5.70264f
C10 VDD2 B 4.756391f
C11 VDD1 B 4.863807f
C12 VTAIL B 5.181212f
C13 VN B 11.255f
C14 VP B 9.895929f
C15 VDD1.n0 B 0.031337f
C16 VDD1.n1 B 0.022295f
C17 VDD1.n2 B 0.01198f
C18 VDD1.n3 B 0.028316f
C19 VDD1.n4 B 0.012685f
C20 VDD1.n5 B 0.022295f
C21 VDD1.n6 B 0.01198f
C22 VDD1.n7 B 0.028316f
C23 VDD1.n8 B 0.012685f
C24 VDD1.n9 B 0.60018f
C25 VDD1.n10 B 0.01198f
C26 VDD1.t4 B 0.046129f
C27 VDD1.n11 B 0.099055f
C28 VDD1.n12 B 0.016727f
C29 VDD1.n13 B 0.021237f
C30 VDD1.n14 B 0.028316f
C31 VDD1.n15 B 0.012685f
C32 VDD1.n16 B 0.01198f
C33 VDD1.n17 B 0.022295f
C34 VDD1.n18 B 0.022295f
C35 VDD1.n19 B 0.01198f
C36 VDD1.n20 B 0.012685f
C37 VDD1.n21 B 0.028316f
C38 VDD1.n22 B 0.028316f
C39 VDD1.n23 B 0.012685f
C40 VDD1.n24 B 0.01198f
C41 VDD1.n25 B 0.022295f
C42 VDD1.n26 B 0.022295f
C43 VDD1.n27 B 0.01198f
C44 VDD1.n28 B 0.012685f
C45 VDD1.n29 B 0.028316f
C46 VDD1.n30 B 0.0613f
C47 VDD1.n31 B 0.012685f
C48 VDD1.n32 B 0.01198f
C49 VDD1.n33 B 0.050314f
C50 VDD1.n34 B 0.055353f
C51 VDD1.n35 B 0.031337f
C52 VDD1.n36 B 0.022295f
C53 VDD1.n37 B 0.01198f
C54 VDD1.n38 B 0.028316f
C55 VDD1.n39 B 0.012685f
C56 VDD1.n40 B 0.022295f
C57 VDD1.n41 B 0.01198f
C58 VDD1.n42 B 0.028316f
C59 VDD1.n43 B 0.012685f
C60 VDD1.n44 B 0.60018f
C61 VDD1.n45 B 0.01198f
C62 VDD1.t2 B 0.046129f
C63 VDD1.n46 B 0.099055f
C64 VDD1.n47 B 0.016727f
C65 VDD1.n48 B 0.021237f
C66 VDD1.n49 B 0.028316f
C67 VDD1.n50 B 0.012685f
C68 VDD1.n51 B 0.01198f
C69 VDD1.n52 B 0.022295f
C70 VDD1.n53 B 0.022295f
C71 VDD1.n54 B 0.01198f
C72 VDD1.n55 B 0.012685f
C73 VDD1.n56 B 0.028316f
C74 VDD1.n57 B 0.028316f
C75 VDD1.n58 B 0.012685f
C76 VDD1.n59 B 0.01198f
C77 VDD1.n60 B 0.022295f
C78 VDD1.n61 B 0.022295f
C79 VDD1.n62 B 0.01198f
C80 VDD1.n63 B 0.012685f
C81 VDD1.n64 B 0.028316f
C82 VDD1.n65 B 0.0613f
C83 VDD1.n66 B 0.012685f
C84 VDD1.n67 B 0.01198f
C85 VDD1.n68 B 0.050314f
C86 VDD1.n69 B 0.054736f
C87 VDD1.t5 B 0.117687f
C88 VDD1.t3 B 0.117687f
C89 VDD1.n70 B 0.996337f
C90 VDD1.n71 B 2.05563f
C91 VDD1.t0 B 0.117687f
C92 VDD1.t1 B 0.117687f
C93 VDD1.n72 B 0.993415f
C94 VDD1.n73 B 2.02646f
C95 VP.n0 B 0.037716f
C96 VP.t2 B 1.13475f
C97 VP.n1 B 0.023437f
C98 VP.n2 B 0.028609f
C99 VP.t0 B 1.13475f
C100 VP.n3 B 0.057236f
C101 VP.n4 B 0.028609f
C102 VP.t3 B 1.13475f
C103 VP.n5 B 0.513419f
C104 VP.n6 B 0.037716f
C105 VP.t4 B 1.13475f
C106 VP.n7 B 0.023437f
C107 VP.n8 B 0.244424f
C108 VP.t5 B 1.13475f
C109 VP.t1 B 1.31622f
C110 VP.n9 B 0.486993f
C111 VP.n10 B 0.498273f
C112 VP.n11 B 0.039958f
C113 VP.n12 B 0.057236f
C114 VP.n13 B 0.028609f
C115 VP.n14 B 0.028609f
C116 VP.n15 B 0.028609f
C117 VP.n16 B 0.055557f
C118 VP.n17 B 0.043101f
C119 VP.n18 B 0.513419f
C120 VP.n19 B 1.2664f
C121 VP.n20 B 1.29027f
C122 VP.n21 B 0.037716f
C123 VP.n22 B 0.043101f
C124 VP.n23 B 0.055557f
C125 VP.n24 B 0.023437f
C126 VP.n25 B 0.028609f
C127 VP.n26 B 0.028609f
C128 VP.n27 B 0.028609f
C129 VP.n28 B 0.039958f
C130 VP.n29 B 0.424308f
C131 VP.n30 B 0.039958f
C132 VP.n31 B 0.057236f
C133 VP.n32 B 0.028609f
C134 VP.n33 B 0.028609f
C135 VP.n34 B 0.028609f
C136 VP.n35 B 0.055557f
C137 VP.n36 B 0.043101f
C138 VP.n37 B 0.513419f
C139 VP.n38 B 0.039717f
C140 VDD2.n0 B 0.030635f
C141 VDD2.n1 B 0.021795f
C142 VDD2.n2 B 0.011712f
C143 VDD2.n3 B 0.027682f
C144 VDD2.n4 B 0.012401f
C145 VDD2.n5 B 0.021795f
C146 VDD2.n6 B 0.011712f
C147 VDD2.n7 B 0.027682f
C148 VDD2.n8 B 0.012401f
C149 VDD2.n9 B 0.586737f
C150 VDD2.n10 B 0.011712f
C151 VDD2.t2 B 0.045095f
C152 VDD2.n11 B 0.096836f
C153 VDD2.n12 B 0.016353f
C154 VDD2.n13 B 0.020762f
C155 VDD2.n14 B 0.027682f
C156 VDD2.n15 B 0.012401f
C157 VDD2.n16 B 0.011712f
C158 VDD2.n17 B 0.021795f
C159 VDD2.n18 B 0.021795f
C160 VDD2.n19 B 0.011712f
C161 VDD2.n20 B 0.012401f
C162 VDD2.n21 B 0.027682f
C163 VDD2.n22 B 0.027682f
C164 VDD2.n23 B 0.012401f
C165 VDD2.n24 B 0.011712f
C166 VDD2.n25 B 0.021795f
C167 VDD2.n26 B 0.021795f
C168 VDD2.n27 B 0.011712f
C169 VDD2.n28 B 0.012401f
C170 VDD2.n29 B 0.027682f
C171 VDD2.n30 B 0.059928f
C172 VDD2.n31 B 0.012401f
C173 VDD2.n32 B 0.011712f
C174 VDD2.n33 B 0.049187f
C175 VDD2.n34 B 0.053511f
C176 VDD2.t3 B 0.115051f
C177 VDD2.t5 B 0.115051f
C178 VDD2.n35 B 0.974021f
C179 VDD2.n36 B 1.91359f
C180 VDD2.n37 B 0.030635f
C181 VDD2.n38 B 0.021795f
C182 VDD2.n39 B 0.011712f
C183 VDD2.n40 B 0.027682f
C184 VDD2.n41 B 0.012401f
C185 VDD2.n42 B 0.021795f
C186 VDD2.n43 B 0.011712f
C187 VDD2.n44 B 0.027682f
C188 VDD2.n45 B 0.012401f
C189 VDD2.n46 B 0.586737f
C190 VDD2.n47 B 0.011712f
C191 VDD2.t0 B 0.045095f
C192 VDD2.n48 B 0.096836f
C193 VDD2.n49 B 0.016353f
C194 VDD2.n50 B 0.020762f
C195 VDD2.n51 B 0.027682f
C196 VDD2.n52 B 0.012401f
C197 VDD2.n53 B 0.011712f
C198 VDD2.n54 B 0.021795f
C199 VDD2.n55 B 0.021795f
C200 VDD2.n56 B 0.011712f
C201 VDD2.n57 B 0.012401f
C202 VDD2.n58 B 0.027682f
C203 VDD2.n59 B 0.027682f
C204 VDD2.n60 B 0.012401f
C205 VDD2.n61 B 0.011712f
C206 VDD2.n62 B 0.021795f
C207 VDD2.n63 B 0.021795f
C208 VDD2.n64 B 0.011712f
C209 VDD2.n65 B 0.012401f
C210 VDD2.n66 B 0.027682f
C211 VDD2.n67 B 0.059928f
C212 VDD2.n68 B 0.012401f
C213 VDD2.n69 B 0.011712f
C214 VDD2.n70 B 0.049187f
C215 VDD2.n71 B 0.048554f
C216 VDD2.n72 B 1.78073f
C217 VDD2.t4 B 0.115051f
C218 VDD2.t1 B 0.115051f
C219 VDD2.n73 B 0.973996f
C220 VTAIL.t9 B 0.137613f
C221 VTAIL.t8 B 0.137613f
C222 VTAIL.n0 B 1.08986f
C223 VTAIL.n1 B 0.433836f
C224 VTAIL.n2 B 0.036643f
C225 VTAIL.n3 B 0.026069f
C226 VTAIL.n4 B 0.014009f
C227 VTAIL.n5 B 0.033111f
C228 VTAIL.n6 B 0.014832f
C229 VTAIL.n7 B 0.026069f
C230 VTAIL.n8 B 0.014009f
C231 VTAIL.n9 B 0.033111f
C232 VTAIL.n10 B 0.014832f
C233 VTAIL.n11 B 0.701801f
C234 VTAIL.n12 B 0.014009f
C235 VTAIL.t0 B 0.053939f
C236 VTAIL.n13 B 0.115827f
C237 VTAIL.n14 B 0.019559f
C238 VTAIL.n15 B 0.024833f
C239 VTAIL.n16 B 0.033111f
C240 VTAIL.n17 B 0.014832f
C241 VTAIL.n18 B 0.014009f
C242 VTAIL.n19 B 0.026069f
C243 VTAIL.n20 B 0.026069f
C244 VTAIL.n21 B 0.014009f
C245 VTAIL.n22 B 0.014832f
C246 VTAIL.n23 B 0.033111f
C247 VTAIL.n24 B 0.033111f
C248 VTAIL.n25 B 0.014832f
C249 VTAIL.n26 B 0.014009f
C250 VTAIL.n27 B 0.026069f
C251 VTAIL.n28 B 0.026069f
C252 VTAIL.n29 B 0.014009f
C253 VTAIL.n30 B 0.014832f
C254 VTAIL.n31 B 0.033111f
C255 VTAIL.n32 B 0.07168f
C256 VTAIL.n33 B 0.014832f
C257 VTAIL.n34 B 0.014009f
C258 VTAIL.n35 B 0.058833f
C259 VTAIL.n36 B 0.040063f
C260 VTAIL.n37 B 0.339f
C261 VTAIL.t3 B 0.137613f
C262 VTAIL.t11 B 0.137613f
C263 VTAIL.n38 B 1.08986f
C264 VTAIL.n39 B 1.64444f
C265 VTAIL.t10 B 0.137613f
C266 VTAIL.t6 B 0.137613f
C267 VTAIL.n40 B 1.08987f
C268 VTAIL.n41 B 1.64444f
C269 VTAIL.n42 B 0.036643f
C270 VTAIL.n43 B 0.026069f
C271 VTAIL.n44 B 0.014009f
C272 VTAIL.n45 B 0.033111f
C273 VTAIL.n46 B 0.014832f
C274 VTAIL.n47 B 0.026069f
C275 VTAIL.n48 B 0.014009f
C276 VTAIL.n49 B 0.033111f
C277 VTAIL.n50 B 0.014832f
C278 VTAIL.n51 B 0.701801f
C279 VTAIL.n52 B 0.014009f
C280 VTAIL.t5 B 0.053939f
C281 VTAIL.n53 B 0.115827f
C282 VTAIL.n54 B 0.019559f
C283 VTAIL.n55 B 0.024833f
C284 VTAIL.n56 B 0.033111f
C285 VTAIL.n57 B 0.014832f
C286 VTAIL.n58 B 0.014009f
C287 VTAIL.n59 B 0.026069f
C288 VTAIL.n60 B 0.026069f
C289 VTAIL.n61 B 0.014009f
C290 VTAIL.n62 B 0.014832f
C291 VTAIL.n63 B 0.033111f
C292 VTAIL.n64 B 0.033111f
C293 VTAIL.n65 B 0.014832f
C294 VTAIL.n66 B 0.014009f
C295 VTAIL.n67 B 0.026069f
C296 VTAIL.n68 B 0.026069f
C297 VTAIL.n69 B 0.014009f
C298 VTAIL.n70 B 0.014832f
C299 VTAIL.n71 B 0.033111f
C300 VTAIL.n72 B 0.07168f
C301 VTAIL.n73 B 0.014832f
C302 VTAIL.n74 B 0.014009f
C303 VTAIL.n75 B 0.058833f
C304 VTAIL.n76 B 0.040063f
C305 VTAIL.n77 B 0.339f
C306 VTAIL.t2 B 0.137613f
C307 VTAIL.t1 B 0.137613f
C308 VTAIL.n78 B 1.08987f
C309 VTAIL.n79 B 0.567977f
C310 VTAIL.n80 B 0.036643f
C311 VTAIL.n81 B 0.026069f
C312 VTAIL.n82 B 0.014009f
C313 VTAIL.n83 B 0.033111f
C314 VTAIL.n84 B 0.014832f
C315 VTAIL.n85 B 0.026069f
C316 VTAIL.n86 B 0.014009f
C317 VTAIL.n87 B 0.033111f
C318 VTAIL.n88 B 0.014832f
C319 VTAIL.n89 B 0.701801f
C320 VTAIL.n90 B 0.014009f
C321 VTAIL.t4 B 0.053939f
C322 VTAIL.n91 B 0.115827f
C323 VTAIL.n92 B 0.019559f
C324 VTAIL.n93 B 0.024833f
C325 VTAIL.n94 B 0.033111f
C326 VTAIL.n95 B 0.014832f
C327 VTAIL.n96 B 0.014009f
C328 VTAIL.n97 B 0.026069f
C329 VTAIL.n98 B 0.026069f
C330 VTAIL.n99 B 0.014009f
C331 VTAIL.n100 B 0.014832f
C332 VTAIL.n101 B 0.033111f
C333 VTAIL.n102 B 0.033111f
C334 VTAIL.n103 B 0.014832f
C335 VTAIL.n104 B 0.014009f
C336 VTAIL.n105 B 0.026069f
C337 VTAIL.n106 B 0.026069f
C338 VTAIL.n107 B 0.014009f
C339 VTAIL.n108 B 0.014832f
C340 VTAIL.n109 B 0.033111f
C341 VTAIL.n110 B 0.07168f
C342 VTAIL.n111 B 0.014832f
C343 VTAIL.n112 B 0.014009f
C344 VTAIL.n113 B 0.058833f
C345 VTAIL.n114 B 0.040063f
C346 VTAIL.n115 B 1.23008f
C347 VTAIL.n116 B 0.036643f
C348 VTAIL.n117 B 0.026069f
C349 VTAIL.n118 B 0.014009f
C350 VTAIL.n119 B 0.033111f
C351 VTAIL.n120 B 0.014832f
C352 VTAIL.n121 B 0.026069f
C353 VTAIL.n122 B 0.014009f
C354 VTAIL.n123 B 0.033111f
C355 VTAIL.n124 B 0.014832f
C356 VTAIL.n125 B 0.701801f
C357 VTAIL.n126 B 0.014009f
C358 VTAIL.t7 B 0.053939f
C359 VTAIL.n127 B 0.115827f
C360 VTAIL.n128 B 0.019559f
C361 VTAIL.n129 B 0.024833f
C362 VTAIL.n130 B 0.033111f
C363 VTAIL.n131 B 0.014832f
C364 VTAIL.n132 B 0.014009f
C365 VTAIL.n133 B 0.026069f
C366 VTAIL.n134 B 0.026069f
C367 VTAIL.n135 B 0.014009f
C368 VTAIL.n136 B 0.014832f
C369 VTAIL.n137 B 0.033111f
C370 VTAIL.n138 B 0.033111f
C371 VTAIL.n139 B 0.014832f
C372 VTAIL.n140 B 0.014009f
C373 VTAIL.n141 B 0.026069f
C374 VTAIL.n142 B 0.026069f
C375 VTAIL.n143 B 0.014009f
C376 VTAIL.n144 B 0.014832f
C377 VTAIL.n145 B 0.033111f
C378 VTAIL.n146 B 0.07168f
C379 VTAIL.n147 B 0.014832f
C380 VTAIL.n148 B 0.014009f
C381 VTAIL.n149 B 0.058833f
C382 VTAIL.n150 B 0.040063f
C383 VTAIL.n151 B 1.17884f
C384 VN.n0 B 0.036796f
C385 VN.t0 B 1.10706f
C386 VN.n1 B 0.022865f
C387 VN.n2 B 0.238458f
C388 VN.t2 B 1.10706f
C389 VN.t3 B 1.2841f
C390 VN.n3 B 0.475108f
C391 VN.n4 B 0.486112f
C392 VN.n5 B 0.038983f
C393 VN.n6 B 0.05584f
C394 VN.n7 B 0.027911f
C395 VN.n8 B 0.027911f
C396 VN.n9 B 0.027911f
C397 VN.n10 B 0.054201f
C398 VN.n11 B 0.042049f
C399 VN.n12 B 0.500889f
C400 VN.n13 B 0.038748f
C401 VN.n14 B 0.036796f
C402 VN.t5 B 1.10706f
C403 VN.n15 B 0.022865f
C404 VN.n16 B 0.238458f
C405 VN.t1 B 1.10706f
C406 VN.t4 B 1.2841f
C407 VN.n17 B 0.475108f
C408 VN.n18 B 0.486112f
C409 VN.n19 B 0.038983f
C410 VN.n20 B 0.05584f
C411 VN.n21 B 0.027911f
C412 VN.n22 B 0.027911f
C413 VN.n23 B 0.027911f
C414 VN.n24 B 0.054201f
C415 VN.n25 B 0.042049f
C416 VN.n26 B 0.500889f
C417 VN.n27 B 1.25087f
.ends

