* NGSPICE file created from diff_pair_sample_1464.ext - technology: sky130A

.subckt diff_pair_sample_1464 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t9 VP.t0 VTAIL.t13 w_n4990_n1980# sky130_fd_pr__pfet_01v8 ad=0.8349 pd=5.39 as=0.8349 ps=5.39 w=5.06 l=3.02
X1 VTAIL.t4 VN.t0 VDD2.t9 w_n4990_n1980# sky130_fd_pr__pfet_01v8 ad=0.8349 pd=5.39 as=0.8349 ps=5.39 w=5.06 l=3.02
X2 B.t11 B.t9 B.t10 w_n4990_n1980# sky130_fd_pr__pfet_01v8 ad=1.9734 pd=10.9 as=0 ps=0 w=5.06 l=3.02
X3 VDD1.t8 VP.t1 VTAIL.t10 w_n4990_n1980# sky130_fd_pr__pfet_01v8 ad=0.8349 pd=5.39 as=1.9734 ps=10.9 w=5.06 l=3.02
X4 VDD1.t7 VP.t2 VTAIL.t15 w_n4990_n1980# sky130_fd_pr__pfet_01v8 ad=0.8349 pd=5.39 as=1.9734 ps=10.9 w=5.06 l=3.02
X5 VTAIL.t3 VN.t1 VDD2.t8 w_n4990_n1980# sky130_fd_pr__pfet_01v8 ad=0.8349 pd=5.39 as=0.8349 ps=5.39 w=5.06 l=3.02
X6 VTAIL.t12 VP.t3 VDD1.t6 w_n4990_n1980# sky130_fd_pr__pfet_01v8 ad=0.8349 pd=5.39 as=0.8349 ps=5.39 w=5.06 l=3.02
X7 VDD1.t5 VP.t4 VTAIL.t6 w_n4990_n1980# sky130_fd_pr__pfet_01v8 ad=1.9734 pd=10.9 as=0.8349 ps=5.39 w=5.06 l=3.02
X8 B.t8 B.t6 B.t7 w_n4990_n1980# sky130_fd_pr__pfet_01v8 ad=1.9734 pd=10.9 as=0 ps=0 w=5.06 l=3.02
X9 VDD2.t7 VN.t2 VTAIL.t17 w_n4990_n1980# sky130_fd_pr__pfet_01v8 ad=0.8349 pd=5.39 as=0.8349 ps=5.39 w=5.06 l=3.02
X10 VDD2.t6 VN.t3 VTAIL.t18 w_n4990_n1980# sky130_fd_pr__pfet_01v8 ad=0.8349 pd=5.39 as=1.9734 ps=10.9 w=5.06 l=3.02
X11 VDD2.t5 VN.t4 VTAIL.t19 w_n4990_n1980# sky130_fd_pr__pfet_01v8 ad=0.8349 pd=5.39 as=1.9734 ps=10.9 w=5.06 l=3.02
X12 VTAIL.t5 VN.t5 VDD2.t4 w_n4990_n1980# sky130_fd_pr__pfet_01v8 ad=0.8349 pd=5.39 as=0.8349 ps=5.39 w=5.06 l=3.02
X13 VDD2.t3 VN.t6 VTAIL.t16 w_n4990_n1980# sky130_fd_pr__pfet_01v8 ad=0.8349 pd=5.39 as=0.8349 ps=5.39 w=5.06 l=3.02
X14 VDD2.t2 VN.t7 VTAIL.t2 w_n4990_n1980# sky130_fd_pr__pfet_01v8 ad=1.9734 pd=10.9 as=0.8349 ps=5.39 w=5.06 l=3.02
X15 VTAIL.t7 VP.t5 VDD1.t4 w_n4990_n1980# sky130_fd_pr__pfet_01v8 ad=0.8349 pd=5.39 as=0.8349 ps=5.39 w=5.06 l=3.02
X16 B.t5 B.t3 B.t4 w_n4990_n1980# sky130_fd_pr__pfet_01v8 ad=1.9734 pd=10.9 as=0 ps=0 w=5.06 l=3.02
X17 VDD2.t1 VN.t8 VTAIL.t0 w_n4990_n1980# sky130_fd_pr__pfet_01v8 ad=1.9734 pd=10.9 as=0.8349 ps=5.39 w=5.06 l=3.02
X18 VTAIL.t1 VN.t9 VDD2.t0 w_n4990_n1980# sky130_fd_pr__pfet_01v8 ad=0.8349 pd=5.39 as=0.8349 ps=5.39 w=5.06 l=3.02
X19 VTAIL.t11 VP.t6 VDD1.t3 w_n4990_n1980# sky130_fd_pr__pfet_01v8 ad=0.8349 pd=5.39 as=0.8349 ps=5.39 w=5.06 l=3.02
X20 B.t2 B.t0 B.t1 w_n4990_n1980# sky130_fd_pr__pfet_01v8 ad=1.9734 pd=10.9 as=0 ps=0 w=5.06 l=3.02
X21 VDD1.t2 VP.t7 VTAIL.t9 w_n4990_n1980# sky130_fd_pr__pfet_01v8 ad=0.8349 pd=5.39 as=0.8349 ps=5.39 w=5.06 l=3.02
X22 VDD1.t1 VP.t8 VTAIL.t14 w_n4990_n1980# sky130_fd_pr__pfet_01v8 ad=1.9734 pd=10.9 as=0.8349 ps=5.39 w=5.06 l=3.02
X23 VTAIL.t8 VP.t9 VDD1.t0 w_n4990_n1980# sky130_fd_pr__pfet_01v8 ad=0.8349 pd=5.39 as=0.8349 ps=5.39 w=5.06 l=3.02
R0 VP.n27 VP.n24 161.3
R1 VP.n29 VP.n28 161.3
R2 VP.n30 VP.n23 161.3
R3 VP.n32 VP.n31 161.3
R4 VP.n33 VP.n22 161.3
R5 VP.n35 VP.n34 161.3
R6 VP.n36 VP.n21 161.3
R7 VP.n39 VP.n38 161.3
R8 VP.n40 VP.n20 161.3
R9 VP.n42 VP.n41 161.3
R10 VP.n43 VP.n19 161.3
R11 VP.n45 VP.n44 161.3
R12 VP.n46 VP.n18 161.3
R13 VP.n48 VP.n47 161.3
R14 VP.n50 VP.n17 161.3
R15 VP.n52 VP.n51 161.3
R16 VP.n53 VP.n16 161.3
R17 VP.n55 VP.n54 161.3
R18 VP.n56 VP.n15 161.3
R19 VP.n58 VP.n57 161.3
R20 VP.n103 VP.n102 161.3
R21 VP.n101 VP.n1 161.3
R22 VP.n100 VP.n99 161.3
R23 VP.n98 VP.n2 161.3
R24 VP.n97 VP.n96 161.3
R25 VP.n95 VP.n3 161.3
R26 VP.n93 VP.n92 161.3
R27 VP.n91 VP.n4 161.3
R28 VP.n90 VP.n89 161.3
R29 VP.n88 VP.n5 161.3
R30 VP.n87 VP.n86 161.3
R31 VP.n85 VP.n6 161.3
R32 VP.n84 VP.n83 161.3
R33 VP.n81 VP.n7 161.3
R34 VP.n80 VP.n79 161.3
R35 VP.n78 VP.n8 161.3
R36 VP.n77 VP.n76 161.3
R37 VP.n75 VP.n9 161.3
R38 VP.n74 VP.n73 161.3
R39 VP.n72 VP.n10 161.3
R40 VP.n71 VP.n70 161.3
R41 VP.n68 VP.n11 161.3
R42 VP.n67 VP.n66 161.3
R43 VP.n65 VP.n12 161.3
R44 VP.n64 VP.n63 161.3
R45 VP.n62 VP.n13 161.3
R46 VP.n26 VP.t4 72.2149
R47 VP.n26 VP.n25 69.111
R48 VP.n61 VP.n60 68.1129
R49 VP.n104 VP.n0 68.1129
R50 VP.n59 VP.n14 68.1129
R51 VP.n67 VP.n12 56.5617
R52 VP.n100 VP.n2 56.5617
R53 VP.n55 VP.n16 56.5617
R54 VP.n60 VP.n59 50.2988
R55 VP.n76 VP.n8 47.8428
R56 VP.n88 VP.n87 47.8428
R57 VP.n43 VP.n42 47.8428
R58 VP.n31 VP.n22 47.8428
R59 VP.n61 VP.t8 40.38
R60 VP.n69 VP.t6 40.38
R61 VP.n82 VP.t7 40.38
R62 VP.n94 VP.t3 40.38
R63 VP.n0 VP.t1 40.38
R64 VP.n14 VP.t2 40.38
R65 VP.n49 VP.t5 40.38
R66 VP.n37 VP.t0 40.38
R67 VP.n25 VP.t9 40.38
R68 VP.n76 VP.n75 33.3113
R69 VP.n89 VP.n88 33.3113
R70 VP.n44 VP.n43 33.3113
R71 VP.n31 VP.n30 33.3113
R72 VP.n63 VP.n62 24.5923
R73 VP.n63 VP.n12 24.5923
R74 VP.n68 VP.n67 24.5923
R75 VP.n70 VP.n68 24.5923
R76 VP.n74 VP.n10 24.5923
R77 VP.n75 VP.n74 24.5923
R78 VP.n80 VP.n8 24.5923
R79 VP.n81 VP.n80 24.5923
R80 VP.n83 VP.n6 24.5923
R81 VP.n87 VP.n6 24.5923
R82 VP.n89 VP.n4 24.5923
R83 VP.n93 VP.n4 24.5923
R84 VP.n96 VP.n95 24.5923
R85 VP.n96 VP.n2 24.5923
R86 VP.n101 VP.n100 24.5923
R87 VP.n102 VP.n101 24.5923
R88 VP.n56 VP.n55 24.5923
R89 VP.n57 VP.n56 24.5923
R90 VP.n44 VP.n18 24.5923
R91 VP.n48 VP.n18 24.5923
R92 VP.n51 VP.n50 24.5923
R93 VP.n51 VP.n16 24.5923
R94 VP.n35 VP.n22 24.5923
R95 VP.n36 VP.n35 24.5923
R96 VP.n38 VP.n20 24.5923
R97 VP.n42 VP.n20 24.5923
R98 VP.n29 VP.n24 24.5923
R99 VP.n30 VP.n29 24.5923
R100 VP.n62 VP.n61 22.1332
R101 VP.n102 VP.n0 22.1332
R102 VP.n57 VP.n14 22.1332
R103 VP.n70 VP.n69 19.674
R104 VP.n95 VP.n94 19.674
R105 VP.n50 VP.n49 19.674
R106 VP.n82 VP.n81 12.2964
R107 VP.n83 VP.n82 12.2964
R108 VP.n37 VP.n36 12.2964
R109 VP.n38 VP.n37 12.2964
R110 VP.n27 VP.n26 5.39128
R111 VP.n69 VP.n10 4.91887
R112 VP.n94 VP.n93 4.91887
R113 VP.n49 VP.n48 4.91887
R114 VP.n25 VP.n24 4.91887
R115 VP.n59 VP.n58 0.354861
R116 VP.n60 VP.n13 0.354861
R117 VP.n104 VP.n103 0.354861
R118 VP VP.n104 0.267071
R119 VP.n28 VP.n27 0.189894
R120 VP.n28 VP.n23 0.189894
R121 VP.n32 VP.n23 0.189894
R122 VP.n33 VP.n32 0.189894
R123 VP.n34 VP.n33 0.189894
R124 VP.n34 VP.n21 0.189894
R125 VP.n39 VP.n21 0.189894
R126 VP.n40 VP.n39 0.189894
R127 VP.n41 VP.n40 0.189894
R128 VP.n41 VP.n19 0.189894
R129 VP.n45 VP.n19 0.189894
R130 VP.n46 VP.n45 0.189894
R131 VP.n47 VP.n46 0.189894
R132 VP.n47 VP.n17 0.189894
R133 VP.n52 VP.n17 0.189894
R134 VP.n53 VP.n52 0.189894
R135 VP.n54 VP.n53 0.189894
R136 VP.n54 VP.n15 0.189894
R137 VP.n58 VP.n15 0.189894
R138 VP.n64 VP.n13 0.189894
R139 VP.n65 VP.n64 0.189894
R140 VP.n66 VP.n65 0.189894
R141 VP.n66 VP.n11 0.189894
R142 VP.n71 VP.n11 0.189894
R143 VP.n72 VP.n71 0.189894
R144 VP.n73 VP.n72 0.189894
R145 VP.n73 VP.n9 0.189894
R146 VP.n77 VP.n9 0.189894
R147 VP.n78 VP.n77 0.189894
R148 VP.n79 VP.n78 0.189894
R149 VP.n79 VP.n7 0.189894
R150 VP.n84 VP.n7 0.189894
R151 VP.n85 VP.n84 0.189894
R152 VP.n86 VP.n85 0.189894
R153 VP.n86 VP.n5 0.189894
R154 VP.n90 VP.n5 0.189894
R155 VP.n91 VP.n90 0.189894
R156 VP.n92 VP.n91 0.189894
R157 VP.n92 VP.n3 0.189894
R158 VP.n97 VP.n3 0.189894
R159 VP.n98 VP.n97 0.189894
R160 VP.n99 VP.n98 0.189894
R161 VP.n99 VP.n1 0.189894
R162 VP.n103 VP.n1 0.189894
R163 VTAIL.n11 VTAIL.t19 92.901
R164 VTAIL.n16 VTAIL.t15 92.9009
R165 VTAIL.n17 VTAIL.t18 92.9009
R166 VTAIL.n2 VTAIL.t10 92.9009
R167 VTAIL.n15 VTAIL.n14 86.4772
R168 VTAIL.n13 VTAIL.n12 86.4772
R169 VTAIL.n10 VTAIL.n9 86.4772
R170 VTAIL.n8 VTAIL.n7 86.4772
R171 VTAIL.n19 VTAIL.n18 86.4769
R172 VTAIL.n1 VTAIL.n0 86.4769
R173 VTAIL.n4 VTAIL.n3 86.4769
R174 VTAIL.n6 VTAIL.n5 86.4769
R175 VTAIL.n8 VTAIL.n6 22.5048
R176 VTAIL.n17 VTAIL.n16 19.6169
R177 VTAIL.n18 VTAIL.t17 6.42441
R178 VTAIL.n18 VTAIL.t5 6.42441
R179 VTAIL.n0 VTAIL.t2 6.42441
R180 VTAIL.n0 VTAIL.t1 6.42441
R181 VTAIL.n3 VTAIL.t9 6.42441
R182 VTAIL.n3 VTAIL.t12 6.42441
R183 VTAIL.n5 VTAIL.t14 6.42441
R184 VTAIL.n5 VTAIL.t11 6.42441
R185 VTAIL.n14 VTAIL.t13 6.42441
R186 VTAIL.n14 VTAIL.t7 6.42441
R187 VTAIL.n12 VTAIL.t6 6.42441
R188 VTAIL.n12 VTAIL.t8 6.42441
R189 VTAIL.n9 VTAIL.t16 6.42441
R190 VTAIL.n9 VTAIL.t3 6.42441
R191 VTAIL.n7 VTAIL.t0 6.42441
R192 VTAIL.n7 VTAIL.t4 6.42441
R193 VTAIL.n10 VTAIL.n8 2.88843
R194 VTAIL.n11 VTAIL.n10 2.88843
R195 VTAIL.n15 VTAIL.n13 2.88843
R196 VTAIL.n16 VTAIL.n15 2.88843
R197 VTAIL.n6 VTAIL.n4 2.88843
R198 VTAIL.n4 VTAIL.n2 2.88843
R199 VTAIL.n19 VTAIL.n17 2.88843
R200 VTAIL VTAIL.n1 2.22464
R201 VTAIL.n13 VTAIL.n11 1.91429
R202 VTAIL.n2 VTAIL.n1 1.91429
R203 VTAIL VTAIL.n19 0.664293
R204 VDD1.n1 VDD1.t5 112.468
R205 VDD1.n3 VDD1.t1 112.468
R206 VDD1.n5 VDD1.n4 105.266
R207 VDD1.n1 VDD1.n0 103.156
R208 VDD1.n7 VDD1.n6 103.156
R209 VDD1.n3 VDD1.n2 103.156
R210 VDD1.n7 VDD1.n5 43.822
R211 VDD1.n6 VDD1.t4 6.42441
R212 VDD1.n6 VDD1.t7 6.42441
R213 VDD1.n0 VDD1.t0 6.42441
R214 VDD1.n0 VDD1.t9 6.42441
R215 VDD1.n4 VDD1.t6 6.42441
R216 VDD1.n4 VDD1.t8 6.42441
R217 VDD1.n2 VDD1.t3 6.42441
R218 VDD1.n2 VDD1.t2 6.42441
R219 VDD1 VDD1.n7 2.10826
R220 VDD1 VDD1.n1 0.780672
R221 VDD1.n5 VDD1.n3 0.667137
R222 VN.n90 VN.n89 161.3
R223 VN.n88 VN.n47 161.3
R224 VN.n87 VN.n86 161.3
R225 VN.n85 VN.n48 161.3
R226 VN.n84 VN.n83 161.3
R227 VN.n82 VN.n49 161.3
R228 VN.n80 VN.n79 161.3
R229 VN.n78 VN.n50 161.3
R230 VN.n77 VN.n76 161.3
R231 VN.n75 VN.n51 161.3
R232 VN.n74 VN.n73 161.3
R233 VN.n72 VN.n52 161.3
R234 VN.n71 VN.n70 161.3
R235 VN.n68 VN.n53 161.3
R236 VN.n67 VN.n66 161.3
R237 VN.n65 VN.n54 161.3
R238 VN.n64 VN.n63 161.3
R239 VN.n62 VN.n55 161.3
R240 VN.n61 VN.n60 161.3
R241 VN.n59 VN.n56 161.3
R242 VN.n44 VN.n43 161.3
R243 VN.n42 VN.n1 161.3
R244 VN.n41 VN.n40 161.3
R245 VN.n39 VN.n2 161.3
R246 VN.n38 VN.n37 161.3
R247 VN.n36 VN.n3 161.3
R248 VN.n34 VN.n33 161.3
R249 VN.n32 VN.n4 161.3
R250 VN.n31 VN.n30 161.3
R251 VN.n29 VN.n5 161.3
R252 VN.n28 VN.n27 161.3
R253 VN.n26 VN.n6 161.3
R254 VN.n25 VN.n24 161.3
R255 VN.n22 VN.n7 161.3
R256 VN.n21 VN.n20 161.3
R257 VN.n19 VN.n8 161.3
R258 VN.n18 VN.n17 161.3
R259 VN.n16 VN.n9 161.3
R260 VN.n15 VN.n14 161.3
R261 VN.n13 VN.n10 161.3
R262 VN.n58 VN.t4 72.2152
R263 VN.n12 VN.t7 72.2152
R264 VN.n58 VN.n57 69.111
R265 VN.n12 VN.n11 69.1109
R266 VN.n45 VN.n0 68.1129
R267 VN.n91 VN.n46 68.1129
R268 VN.n41 VN.n2 56.5617
R269 VN.n87 VN.n48 56.5617
R270 VN VN.n91 50.464
R271 VN.n17 VN.n8 47.8428
R272 VN.n29 VN.n28 47.8428
R273 VN.n63 VN.n54 47.8428
R274 VN.n75 VN.n74 47.8428
R275 VN.n11 VN.t9 40.38
R276 VN.n23 VN.t2 40.38
R277 VN.n35 VN.t5 40.38
R278 VN.n0 VN.t3 40.38
R279 VN.n57 VN.t1 40.38
R280 VN.n69 VN.t6 40.38
R281 VN.n81 VN.t0 40.38
R282 VN.n46 VN.t8 40.38
R283 VN.n17 VN.n16 33.3113
R284 VN.n30 VN.n29 33.3113
R285 VN.n63 VN.n62 33.3113
R286 VN.n76 VN.n75 33.3113
R287 VN.n15 VN.n10 24.5923
R288 VN.n16 VN.n15 24.5923
R289 VN.n21 VN.n8 24.5923
R290 VN.n22 VN.n21 24.5923
R291 VN.n24 VN.n6 24.5923
R292 VN.n28 VN.n6 24.5923
R293 VN.n30 VN.n4 24.5923
R294 VN.n34 VN.n4 24.5923
R295 VN.n37 VN.n36 24.5923
R296 VN.n37 VN.n2 24.5923
R297 VN.n42 VN.n41 24.5923
R298 VN.n43 VN.n42 24.5923
R299 VN.n62 VN.n61 24.5923
R300 VN.n61 VN.n56 24.5923
R301 VN.n74 VN.n52 24.5923
R302 VN.n70 VN.n52 24.5923
R303 VN.n68 VN.n67 24.5923
R304 VN.n67 VN.n54 24.5923
R305 VN.n83 VN.n48 24.5923
R306 VN.n83 VN.n82 24.5923
R307 VN.n80 VN.n50 24.5923
R308 VN.n76 VN.n50 24.5923
R309 VN.n89 VN.n88 24.5923
R310 VN.n88 VN.n87 24.5923
R311 VN.n43 VN.n0 22.1332
R312 VN.n89 VN.n46 22.1332
R313 VN.n36 VN.n35 19.674
R314 VN.n82 VN.n81 19.674
R315 VN.n23 VN.n22 12.2964
R316 VN.n24 VN.n23 12.2964
R317 VN.n70 VN.n69 12.2964
R318 VN.n69 VN.n68 12.2964
R319 VN.n59 VN.n58 5.39131
R320 VN.n13 VN.n12 5.39131
R321 VN.n11 VN.n10 4.91887
R322 VN.n35 VN.n34 4.91887
R323 VN.n57 VN.n56 4.91887
R324 VN.n81 VN.n80 4.91887
R325 VN.n91 VN.n90 0.354861
R326 VN.n45 VN.n44 0.354861
R327 VN VN.n45 0.267071
R328 VN.n90 VN.n47 0.189894
R329 VN.n86 VN.n47 0.189894
R330 VN.n86 VN.n85 0.189894
R331 VN.n85 VN.n84 0.189894
R332 VN.n84 VN.n49 0.189894
R333 VN.n79 VN.n49 0.189894
R334 VN.n79 VN.n78 0.189894
R335 VN.n78 VN.n77 0.189894
R336 VN.n77 VN.n51 0.189894
R337 VN.n73 VN.n51 0.189894
R338 VN.n73 VN.n72 0.189894
R339 VN.n72 VN.n71 0.189894
R340 VN.n71 VN.n53 0.189894
R341 VN.n66 VN.n53 0.189894
R342 VN.n66 VN.n65 0.189894
R343 VN.n65 VN.n64 0.189894
R344 VN.n64 VN.n55 0.189894
R345 VN.n60 VN.n55 0.189894
R346 VN.n60 VN.n59 0.189894
R347 VN.n14 VN.n13 0.189894
R348 VN.n14 VN.n9 0.189894
R349 VN.n18 VN.n9 0.189894
R350 VN.n19 VN.n18 0.189894
R351 VN.n20 VN.n19 0.189894
R352 VN.n20 VN.n7 0.189894
R353 VN.n25 VN.n7 0.189894
R354 VN.n26 VN.n25 0.189894
R355 VN.n27 VN.n26 0.189894
R356 VN.n27 VN.n5 0.189894
R357 VN.n31 VN.n5 0.189894
R358 VN.n32 VN.n31 0.189894
R359 VN.n33 VN.n32 0.189894
R360 VN.n33 VN.n3 0.189894
R361 VN.n38 VN.n3 0.189894
R362 VN.n39 VN.n38 0.189894
R363 VN.n40 VN.n39 0.189894
R364 VN.n40 VN.n1 0.189894
R365 VN.n44 VN.n1 0.189894
R366 VDD2.n1 VDD2.t2 112.468
R367 VDD2.n4 VDD2.t1 109.579
R368 VDD2.n3 VDD2.n2 105.266
R369 VDD2 VDD2.n7 105.263
R370 VDD2.n6 VDD2.n5 103.156
R371 VDD2.n1 VDD2.n0 103.156
R372 VDD2.n4 VDD2.n3 41.795
R373 VDD2.n7 VDD2.t8 6.42441
R374 VDD2.n7 VDD2.t5 6.42441
R375 VDD2.n5 VDD2.t9 6.42441
R376 VDD2.n5 VDD2.t3 6.42441
R377 VDD2.n2 VDD2.t4 6.42441
R378 VDD2.n2 VDD2.t6 6.42441
R379 VDD2.n0 VDD2.t0 6.42441
R380 VDD2.n0 VDD2.t7 6.42441
R381 VDD2.n6 VDD2.n4 2.88843
R382 VDD2 VDD2.n6 0.780672
R383 VDD2.n3 VDD2.n1 0.667137
R384 B.n579 B.n578 585
R385 B.n580 B.n65 585
R386 B.n582 B.n581 585
R387 B.n583 B.n64 585
R388 B.n585 B.n584 585
R389 B.n586 B.n63 585
R390 B.n588 B.n587 585
R391 B.n589 B.n62 585
R392 B.n591 B.n590 585
R393 B.n592 B.n61 585
R394 B.n594 B.n593 585
R395 B.n595 B.n60 585
R396 B.n597 B.n596 585
R397 B.n598 B.n59 585
R398 B.n600 B.n599 585
R399 B.n601 B.n58 585
R400 B.n603 B.n602 585
R401 B.n604 B.n57 585
R402 B.n606 B.n605 585
R403 B.n607 B.n56 585
R404 B.n609 B.n608 585
R405 B.n611 B.n53 585
R406 B.n613 B.n612 585
R407 B.n614 B.n52 585
R408 B.n616 B.n615 585
R409 B.n617 B.n51 585
R410 B.n619 B.n618 585
R411 B.n620 B.n50 585
R412 B.n622 B.n621 585
R413 B.n623 B.n49 585
R414 B.n625 B.n624 585
R415 B.n627 B.n626 585
R416 B.n628 B.n45 585
R417 B.n630 B.n629 585
R418 B.n631 B.n44 585
R419 B.n633 B.n632 585
R420 B.n634 B.n43 585
R421 B.n636 B.n635 585
R422 B.n637 B.n42 585
R423 B.n639 B.n638 585
R424 B.n640 B.n41 585
R425 B.n642 B.n641 585
R426 B.n643 B.n40 585
R427 B.n645 B.n644 585
R428 B.n646 B.n39 585
R429 B.n648 B.n647 585
R430 B.n649 B.n38 585
R431 B.n651 B.n650 585
R432 B.n652 B.n37 585
R433 B.n654 B.n653 585
R434 B.n655 B.n36 585
R435 B.n657 B.n656 585
R436 B.n577 B.n66 585
R437 B.n576 B.n575 585
R438 B.n574 B.n67 585
R439 B.n573 B.n572 585
R440 B.n571 B.n68 585
R441 B.n570 B.n569 585
R442 B.n568 B.n69 585
R443 B.n567 B.n566 585
R444 B.n565 B.n70 585
R445 B.n564 B.n563 585
R446 B.n562 B.n71 585
R447 B.n561 B.n560 585
R448 B.n559 B.n72 585
R449 B.n558 B.n557 585
R450 B.n556 B.n73 585
R451 B.n555 B.n554 585
R452 B.n553 B.n74 585
R453 B.n552 B.n551 585
R454 B.n550 B.n75 585
R455 B.n549 B.n548 585
R456 B.n547 B.n76 585
R457 B.n546 B.n545 585
R458 B.n544 B.n77 585
R459 B.n543 B.n542 585
R460 B.n541 B.n78 585
R461 B.n540 B.n539 585
R462 B.n538 B.n79 585
R463 B.n537 B.n536 585
R464 B.n535 B.n80 585
R465 B.n534 B.n533 585
R466 B.n532 B.n81 585
R467 B.n531 B.n530 585
R468 B.n529 B.n82 585
R469 B.n528 B.n527 585
R470 B.n526 B.n83 585
R471 B.n525 B.n524 585
R472 B.n523 B.n84 585
R473 B.n522 B.n521 585
R474 B.n520 B.n85 585
R475 B.n519 B.n518 585
R476 B.n517 B.n86 585
R477 B.n516 B.n515 585
R478 B.n514 B.n87 585
R479 B.n513 B.n512 585
R480 B.n511 B.n88 585
R481 B.n510 B.n509 585
R482 B.n508 B.n89 585
R483 B.n507 B.n506 585
R484 B.n505 B.n90 585
R485 B.n504 B.n503 585
R486 B.n502 B.n91 585
R487 B.n501 B.n500 585
R488 B.n499 B.n92 585
R489 B.n498 B.n497 585
R490 B.n496 B.n93 585
R491 B.n495 B.n494 585
R492 B.n493 B.n94 585
R493 B.n492 B.n491 585
R494 B.n490 B.n95 585
R495 B.n489 B.n488 585
R496 B.n487 B.n96 585
R497 B.n486 B.n485 585
R498 B.n484 B.n97 585
R499 B.n483 B.n482 585
R500 B.n481 B.n98 585
R501 B.n480 B.n479 585
R502 B.n478 B.n99 585
R503 B.n477 B.n476 585
R504 B.n475 B.n100 585
R505 B.n474 B.n473 585
R506 B.n472 B.n101 585
R507 B.n471 B.n470 585
R508 B.n469 B.n102 585
R509 B.n468 B.n467 585
R510 B.n466 B.n103 585
R511 B.n465 B.n464 585
R512 B.n463 B.n104 585
R513 B.n462 B.n461 585
R514 B.n460 B.n105 585
R515 B.n459 B.n458 585
R516 B.n457 B.n106 585
R517 B.n456 B.n455 585
R518 B.n454 B.n107 585
R519 B.n453 B.n452 585
R520 B.n451 B.n108 585
R521 B.n450 B.n449 585
R522 B.n448 B.n109 585
R523 B.n447 B.n446 585
R524 B.n445 B.n110 585
R525 B.n444 B.n443 585
R526 B.n442 B.n111 585
R527 B.n441 B.n440 585
R528 B.n439 B.n112 585
R529 B.n438 B.n437 585
R530 B.n436 B.n113 585
R531 B.n435 B.n434 585
R532 B.n433 B.n114 585
R533 B.n432 B.n431 585
R534 B.n430 B.n115 585
R535 B.n429 B.n428 585
R536 B.n427 B.n116 585
R537 B.n426 B.n425 585
R538 B.n424 B.n117 585
R539 B.n423 B.n422 585
R540 B.n421 B.n118 585
R541 B.n420 B.n419 585
R542 B.n418 B.n119 585
R543 B.n417 B.n416 585
R544 B.n415 B.n120 585
R545 B.n414 B.n413 585
R546 B.n412 B.n121 585
R547 B.n411 B.n410 585
R548 B.n409 B.n122 585
R549 B.n408 B.n407 585
R550 B.n406 B.n123 585
R551 B.n405 B.n404 585
R552 B.n403 B.n124 585
R553 B.n402 B.n401 585
R554 B.n400 B.n125 585
R555 B.n399 B.n398 585
R556 B.n397 B.n126 585
R557 B.n396 B.n395 585
R558 B.n394 B.n127 585
R559 B.n393 B.n392 585
R560 B.n391 B.n128 585
R561 B.n390 B.n389 585
R562 B.n388 B.n129 585
R563 B.n387 B.n386 585
R564 B.n385 B.n130 585
R565 B.n384 B.n383 585
R566 B.n382 B.n131 585
R567 B.n381 B.n380 585
R568 B.n379 B.n132 585
R569 B.n378 B.n377 585
R570 B.n376 B.n133 585
R571 B.n297 B.n296 585
R572 B.n298 B.n163 585
R573 B.n300 B.n299 585
R574 B.n301 B.n162 585
R575 B.n303 B.n302 585
R576 B.n304 B.n161 585
R577 B.n306 B.n305 585
R578 B.n307 B.n160 585
R579 B.n309 B.n308 585
R580 B.n310 B.n159 585
R581 B.n312 B.n311 585
R582 B.n313 B.n158 585
R583 B.n315 B.n314 585
R584 B.n316 B.n157 585
R585 B.n318 B.n317 585
R586 B.n319 B.n156 585
R587 B.n321 B.n320 585
R588 B.n322 B.n155 585
R589 B.n324 B.n323 585
R590 B.n325 B.n154 585
R591 B.n327 B.n326 585
R592 B.n329 B.n151 585
R593 B.n331 B.n330 585
R594 B.n332 B.n150 585
R595 B.n334 B.n333 585
R596 B.n335 B.n149 585
R597 B.n337 B.n336 585
R598 B.n338 B.n148 585
R599 B.n340 B.n339 585
R600 B.n341 B.n147 585
R601 B.n343 B.n342 585
R602 B.n345 B.n344 585
R603 B.n346 B.n143 585
R604 B.n348 B.n347 585
R605 B.n349 B.n142 585
R606 B.n351 B.n350 585
R607 B.n352 B.n141 585
R608 B.n354 B.n353 585
R609 B.n355 B.n140 585
R610 B.n357 B.n356 585
R611 B.n358 B.n139 585
R612 B.n360 B.n359 585
R613 B.n361 B.n138 585
R614 B.n363 B.n362 585
R615 B.n364 B.n137 585
R616 B.n366 B.n365 585
R617 B.n367 B.n136 585
R618 B.n369 B.n368 585
R619 B.n370 B.n135 585
R620 B.n372 B.n371 585
R621 B.n373 B.n134 585
R622 B.n375 B.n374 585
R623 B.n295 B.n164 585
R624 B.n294 B.n293 585
R625 B.n292 B.n165 585
R626 B.n291 B.n290 585
R627 B.n289 B.n166 585
R628 B.n288 B.n287 585
R629 B.n286 B.n167 585
R630 B.n285 B.n284 585
R631 B.n283 B.n168 585
R632 B.n282 B.n281 585
R633 B.n280 B.n169 585
R634 B.n279 B.n278 585
R635 B.n277 B.n170 585
R636 B.n276 B.n275 585
R637 B.n274 B.n171 585
R638 B.n273 B.n272 585
R639 B.n271 B.n172 585
R640 B.n270 B.n269 585
R641 B.n268 B.n173 585
R642 B.n267 B.n266 585
R643 B.n265 B.n174 585
R644 B.n264 B.n263 585
R645 B.n262 B.n175 585
R646 B.n261 B.n260 585
R647 B.n259 B.n176 585
R648 B.n258 B.n257 585
R649 B.n256 B.n177 585
R650 B.n255 B.n254 585
R651 B.n253 B.n178 585
R652 B.n252 B.n251 585
R653 B.n250 B.n179 585
R654 B.n249 B.n248 585
R655 B.n247 B.n180 585
R656 B.n246 B.n245 585
R657 B.n244 B.n181 585
R658 B.n243 B.n242 585
R659 B.n241 B.n182 585
R660 B.n240 B.n239 585
R661 B.n238 B.n183 585
R662 B.n237 B.n236 585
R663 B.n235 B.n184 585
R664 B.n234 B.n233 585
R665 B.n232 B.n185 585
R666 B.n231 B.n230 585
R667 B.n229 B.n186 585
R668 B.n228 B.n227 585
R669 B.n226 B.n187 585
R670 B.n225 B.n224 585
R671 B.n223 B.n188 585
R672 B.n222 B.n221 585
R673 B.n220 B.n189 585
R674 B.n219 B.n218 585
R675 B.n217 B.n190 585
R676 B.n216 B.n215 585
R677 B.n214 B.n191 585
R678 B.n213 B.n212 585
R679 B.n211 B.n192 585
R680 B.n210 B.n209 585
R681 B.n208 B.n193 585
R682 B.n207 B.n206 585
R683 B.n205 B.n194 585
R684 B.n204 B.n203 585
R685 B.n202 B.n195 585
R686 B.n201 B.n200 585
R687 B.n199 B.n196 585
R688 B.n198 B.n197 585
R689 B.n2 B.n0 585
R690 B.n757 B.n1 585
R691 B.n756 B.n755 585
R692 B.n754 B.n3 585
R693 B.n753 B.n752 585
R694 B.n751 B.n4 585
R695 B.n750 B.n749 585
R696 B.n748 B.n5 585
R697 B.n747 B.n746 585
R698 B.n745 B.n6 585
R699 B.n744 B.n743 585
R700 B.n742 B.n7 585
R701 B.n741 B.n740 585
R702 B.n739 B.n8 585
R703 B.n738 B.n737 585
R704 B.n736 B.n9 585
R705 B.n735 B.n734 585
R706 B.n733 B.n10 585
R707 B.n732 B.n731 585
R708 B.n730 B.n11 585
R709 B.n729 B.n728 585
R710 B.n727 B.n12 585
R711 B.n726 B.n725 585
R712 B.n724 B.n13 585
R713 B.n723 B.n722 585
R714 B.n721 B.n14 585
R715 B.n720 B.n719 585
R716 B.n718 B.n15 585
R717 B.n717 B.n716 585
R718 B.n715 B.n16 585
R719 B.n714 B.n713 585
R720 B.n712 B.n17 585
R721 B.n711 B.n710 585
R722 B.n709 B.n18 585
R723 B.n708 B.n707 585
R724 B.n706 B.n19 585
R725 B.n705 B.n704 585
R726 B.n703 B.n20 585
R727 B.n702 B.n701 585
R728 B.n700 B.n21 585
R729 B.n699 B.n698 585
R730 B.n697 B.n22 585
R731 B.n696 B.n695 585
R732 B.n694 B.n23 585
R733 B.n693 B.n692 585
R734 B.n691 B.n24 585
R735 B.n690 B.n689 585
R736 B.n688 B.n25 585
R737 B.n687 B.n686 585
R738 B.n685 B.n26 585
R739 B.n684 B.n683 585
R740 B.n682 B.n27 585
R741 B.n681 B.n680 585
R742 B.n679 B.n28 585
R743 B.n678 B.n677 585
R744 B.n676 B.n29 585
R745 B.n675 B.n674 585
R746 B.n673 B.n30 585
R747 B.n672 B.n671 585
R748 B.n670 B.n31 585
R749 B.n669 B.n668 585
R750 B.n667 B.n32 585
R751 B.n666 B.n665 585
R752 B.n664 B.n33 585
R753 B.n663 B.n662 585
R754 B.n661 B.n34 585
R755 B.n660 B.n659 585
R756 B.n658 B.n35 585
R757 B.n759 B.n758 585
R758 B.n296 B.n295 535.745
R759 B.n656 B.n35 535.745
R760 B.n374 B.n133 535.745
R761 B.n578 B.n577 535.745
R762 B.n144 B.t0 248.983
R763 B.n152 B.t3 248.983
R764 B.n46 B.t9 248.983
R765 B.n54 B.t6 248.983
R766 B.n144 B.t2 185.231
R767 B.n54 B.t7 185.231
R768 B.n152 B.t5 185.226
R769 B.n46 B.t10 185.226
R770 B.n295 B.n294 163.367
R771 B.n294 B.n165 163.367
R772 B.n290 B.n165 163.367
R773 B.n290 B.n289 163.367
R774 B.n289 B.n288 163.367
R775 B.n288 B.n167 163.367
R776 B.n284 B.n167 163.367
R777 B.n284 B.n283 163.367
R778 B.n283 B.n282 163.367
R779 B.n282 B.n169 163.367
R780 B.n278 B.n169 163.367
R781 B.n278 B.n277 163.367
R782 B.n277 B.n276 163.367
R783 B.n276 B.n171 163.367
R784 B.n272 B.n171 163.367
R785 B.n272 B.n271 163.367
R786 B.n271 B.n270 163.367
R787 B.n270 B.n173 163.367
R788 B.n266 B.n173 163.367
R789 B.n266 B.n265 163.367
R790 B.n265 B.n264 163.367
R791 B.n264 B.n175 163.367
R792 B.n260 B.n175 163.367
R793 B.n260 B.n259 163.367
R794 B.n259 B.n258 163.367
R795 B.n258 B.n177 163.367
R796 B.n254 B.n177 163.367
R797 B.n254 B.n253 163.367
R798 B.n253 B.n252 163.367
R799 B.n252 B.n179 163.367
R800 B.n248 B.n179 163.367
R801 B.n248 B.n247 163.367
R802 B.n247 B.n246 163.367
R803 B.n246 B.n181 163.367
R804 B.n242 B.n181 163.367
R805 B.n242 B.n241 163.367
R806 B.n241 B.n240 163.367
R807 B.n240 B.n183 163.367
R808 B.n236 B.n183 163.367
R809 B.n236 B.n235 163.367
R810 B.n235 B.n234 163.367
R811 B.n234 B.n185 163.367
R812 B.n230 B.n185 163.367
R813 B.n230 B.n229 163.367
R814 B.n229 B.n228 163.367
R815 B.n228 B.n187 163.367
R816 B.n224 B.n187 163.367
R817 B.n224 B.n223 163.367
R818 B.n223 B.n222 163.367
R819 B.n222 B.n189 163.367
R820 B.n218 B.n189 163.367
R821 B.n218 B.n217 163.367
R822 B.n217 B.n216 163.367
R823 B.n216 B.n191 163.367
R824 B.n212 B.n191 163.367
R825 B.n212 B.n211 163.367
R826 B.n211 B.n210 163.367
R827 B.n210 B.n193 163.367
R828 B.n206 B.n193 163.367
R829 B.n206 B.n205 163.367
R830 B.n205 B.n204 163.367
R831 B.n204 B.n195 163.367
R832 B.n200 B.n195 163.367
R833 B.n200 B.n199 163.367
R834 B.n199 B.n198 163.367
R835 B.n198 B.n2 163.367
R836 B.n758 B.n2 163.367
R837 B.n758 B.n757 163.367
R838 B.n757 B.n756 163.367
R839 B.n756 B.n3 163.367
R840 B.n752 B.n3 163.367
R841 B.n752 B.n751 163.367
R842 B.n751 B.n750 163.367
R843 B.n750 B.n5 163.367
R844 B.n746 B.n5 163.367
R845 B.n746 B.n745 163.367
R846 B.n745 B.n744 163.367
R847 B.n744 B.n7 163.367
R848 B.n740 B.n7 163.367
R849 B.n740 B.n739 163.367
R850 B.n739 B.n738 163.367
R851 B.n738 B.n9 163.367
R852 B.n734 B.n9 163.367
R853 B.n734 B.n733 163.367
R854 B.n733 B.n732 163.367
R855 B.n732 B.n11 163.367
R856 B.n728 B.n11 163.367
R857 B.n728 B.n727 163.367
R858 B.n727 B.n726 163.367
R859 B.n726 B.n13 163.367
R860 B.n722 B.n13 163.367
R861 B.n722 B.n721 163.367
R862 B.n721 B.n720 163.367
R863 B.n720 B.n15 163.367
R864 B.n716 B.n15 163.367
R865 B.n716 B.n715 163.367
R866 B.n715 B.n714 163.367
R867 B.n714 B.n17 163.367
R868 B.n710 B.n17 163.367
R869 B.n710 B.n709 163.367
R870 B.n709 B.n708 163.367
R871 B.n708 B.n19 163.367
R872 B.n704 B.n19 163.367
R873 B.n704 B.n703 163.367
R874 B.n703 B.n702 163.367
R875 B.n702 B.n21 163.367
R876 B.n698 B.n21 163.367
R877 B.n698 B.n697 163.367
R878 B.n697 B.n696 163.367
R879 B.n696 B.n23 163.367
R880 B.n692 B.n23 163.367
R881 B.n692 B.n691 163.367
R882 B.n691 B.n690 163.367
R883 B.n690 B.n25 163.367
R884 B.n686 B.n25 163.367
R885 B.n686 B.n685 163.367
R886 B.n685 B.n684 163.367
R887 B.n684 B.n27 163.367
R888 B.n680 B.n27 163.367
R889 B.n680 B.n679 163.367
R890 B.n679 B.n678 163.367
R891 B.n678 B.n29 163.367
R892 B.n674 B.n29 163.367
R893 B.n674 B.n673 163.367
R894 B.n673 B.n672 163.367
R895 B.n672 B.n31 163.367
R896 B.n668 B.n31 163.367
R897 B.n668 B.n667 163.367
R898 B.n667 B.n666 163.367
R899 B.n666 B.n33 163.367
R900 B.n662 B.n33 163.367
R901 B.n662 B.n661 163.367
R902 B.n661 B.n660 163.367
R903 B.n660 B.n35 163.367
R904 B.n296 B.n163 163.367
R905 B.n300 B.n163 163.367
R906 B.n301 B.n300 163.367
R907 B.n302 B.n301 163.367
R908 B.n302 B.n161 163.367
R909 B.n306 B.n161 163.367
R910 B.n307 B.n306 163.367
R911 B.n308 B.n307 163.367
R912 B.n308 B.n159 163.367
R913 B.n312 B.n159 163.367
R914 B.n313 B.n312 163.367
R915 B.n314 B.n313 163.367
R916 B.n314 B.n157 163.367
R917 B.n318 B.n157 163.367
R918 B.n319 B.n318 163.367
R919 B.n320 B.n319 163.367
R920 B.n320 B.n155 163.367
R921 B.n324 B.n155 163.367
R922 B.n325 B.n324 163.367
R923 B.n326 B.n325 163.367
R924 B.n326 B.n151 163.367
R925 B.n331 B.n151 163.367
R926 B.n332 B.n331 163.367
R927 B.n333 B.n332 163.367
R928 B.n333 B.n149 163.367
R929 B.n337 B.n149 163.367
R930 B.n338 B.n337 163.367
R931 B.n339 B.n338 163.367
R932 B.n339 B.n147 163.367
R933 B.n343 B.n147 163.367
R934 B.n344 B.n343 163.367
R935 B.n344 B.n143 163.367
R936 B.n348 B.n143 163.367
R937 B.n349 B.n348 163.367
R938 B.n350 B.n349 163.367
R939 B.n350 B.n141 163.367
R940 B.n354 B.n141 163.367
R941 B.n355 B.n354 163.367
R942 B.n356 B.n355 163.367
R943 B.n356 B.n139 163.367
R944 B.n360 B.n139 163.367
R945 B.n361 B.n360 163.367
R946 B.n362 B.n361 163.367
R947 B.n362 B.n137 163.367
R948 B.n366 B.n137 163.367
R949 B.n367 B.n366 163.367
R950 B.n368 B.n367 163.367
R951 B.n368 B.n135 163.367
R952 B.n372 B.n135 163.367
R953 B.n373 B.n372 163.367
R954 B.n374 B.n373 163.367
R955 B.n378 B.n133 163.367
R956 B.n379 B.n378 163.367
R957 B.n380 B.n379 163.367
R958 B.n380 B.n131 163.367
R959 B.n384 B.n131 163.367
R960 B.n385 B.n384 163.367
R961 B.n386 B.n385 163.367
R962 B.n386 B.n129 163.367
R963 B.n390 B.n129 163.367
R964 B.n391 B.n390 163.367
R965 B.n392 B.n391 163.367
R966 B.n392 B.n127 163.367
R967 B.n396 B.n127 163.367
R968 B.n397 B.n396 163.367
R969 B.n398 B.n397 163.367
R970 B.n398 B.n125 163.367
R971 B.n402 B.n125 163.367
R972 B.n403 B.n402 163.367
R973 B.n404 B.n403 163.367
R974 B.n404 B.n123 163.367
R975 B.n408 B.n123 163.367
R976 B.n409 B.n408 163.367
R977 B.n410 B.n409 163.367
R978 B.n410 B.n121 163.367
R979 B.n414 B.n121 163.367
R980 B.n415 B.n414 163.367
R981 B.n416 B.n415 163.367
R982 B.n416 B.n119 163.367
R983 B.n420 B.n119 163.367
R984 B.n421 B.n420 163.367
R985 B.n422 B.n421 163.367
R986 B.n422 B.n117 163.367
R987 B.n426 B.n117 163.367
R988 B.n427 B.n426 163.367
R989 B.n428 B.n427 163.367
R990 B.n428 B.n115 163.367
R991 B.n432 B.n115 163.367
R992 B.n433 B.n432 163.367
R993 B.n434 B.n433 163.367
R994 B.n434 B.n113 163.367
R995 B.n438 B.n113 163.367
R996 B.n439 B.n438 163.367
R997 B.n440 B.n439 163.367
R998 B.n440 B.n111 163.367
R999 B.n444 B.n111 163.367
R1000 B.n445 B.n444 163.367
R1001 B.n446 B.n445 163.367
R1002 B.n446 B.n109 163.367
R1003 B.n450 B.n109 163.367
R1004 B.n451 B.n450 163.367
R1005 B.n452 B.n451 163.367
R1006 B.n452 B.n107 163.367
R1007 B.n456 B.n107 163.367
R1008 B.n457 B.n456 163.367
R1009 B.n458 B.n457 163.367
R1010 B.n458 B.n105 163.367
R1011 B.n462 B.n105 163.367
R1012 B.n463 B.n462 163.367
R1013 B.n464 B.n463 163.367
R1014 B.n464 B.n103 163.367
R1015 B.n468 B.n103 163.367
R1016 B.n469 B.n468 163.367
R1017 B.n470 B.n469 163.367
R1018 B.n470 B.n101 163.367
R1019 B.n474 B.n101 163.367
R1020 B.n475 B.n474 163.367
R1021 B.n476 B.n475 163.367
R1022 B.n476 B.n99 163.367
R1023 B.n480 B.n99 163.367
R1024 B.n481 B.n480 163.367
R1025 B.n482 B.n481 163.367
R1026 B.n482 B.n97 163.367
R1027 B.n486 B.n97 163.367
R1028 B.n487 B.n486 163.367
R1029 B.n488 B.n487 163.367
R1030 B.n488 B.n95 163.367
R1031 B.n492 B.n95 163.367
R1032 B.n493 B.n492 163.367
R1033 B.n494 B.n493 163.367
R1034 B.n494 B.n93 163.367
R1035 B.n498 B.n93 163.367
R1036 B.n499 B.n498 163.367
R1037 B.n500 B.n499 163.367
R1038 B.n500 B.n91 163.367
R1039 B.n504 B.n91 163.367
R1040 B.n505 B.n504 163.367
R1041 B.n506 B.n505 163.367
R1042 B.n506 B.n89 163.367
R1043 B.n510 B.n89 163.367
R1044 B.n511 B.n510 163.367
R1045 B.n512 B.n511 163.367
R1046 B.n512 B.n87 163.367
R1047 B.n516 B.n87 163.367
R1048 B.n517 B.n516 163.367
R1049 B.n518 B.n517 163.367
R1050 B.n518 B.n85 163.367
R1051 B.n522 B.n85 163.367
R1052 B.n523 B.n522 163.367
R1053 B.n524 B.n523 163.367
R1054 B.n524 B.n83 163.367
R1055 B.n528 B.n83 163.367
R1056 B.n529 B.n528 163.367
R1057 B.n530 B.n529 163.367
R1058 B.n530 B.n81 163.367
R1059 B.n534 B.n81 163.367
R1060 B.n535 B.n534 163.367
R1061 B.n536 B.n535 163.367
R1062 B.n536 B.n79 163.367
R1063 B.n540 B.n79 163.367
R1064 B.n541 B.n540 163.367
R1065 B.n542 B.n541 163.367
R1066 B.n542 B.n77 163.367
R1067 B.n546 B.n77 163.367
R1068 B.n547 B.n546 163.367
R1069 B.n548 B.n547 163.367
R1070 B.n548 B.n75 163.367
R1071 B.n552 B.n75 163.367
R1072 B.n553 B.n552 163.367
R1073 B.n554 B.n553 163.367
R1074 B.n554 B.n73 163.367
R1075 B.n558 B.n73 163.367
R1076 B.n559 B.n558 163.367
R1077 B.n560 B.n559 163.367
R1078 B.n560 B.n71 163.367
R1079 B.n564 B.n71 163.367
R1080 B.n565 B.n564 163.367
R1081 B.n566 B.n565 163.367
R1082 B.n566 B.n69 163.367
R1083 B.n570 B.n69 163.367
R1084 B.n571 B.n570 163.367
R1085 B.n572 B.n571 163.367
R1086 B.n572 B.n67 163.367
R1087 B.n576 B.n67 163.367
R1088 B.n577 B.n576 163.367
R1089 B.n656 B.n655 163.367
R1090 B.n655 B.n654 163.367
R1091 B.n654 B.n37 163.367
R1092 B.n650 B.n37 163.367
R1093 B.n650 B.n649 163.367
R1094 B.n649 B.n648 163.367
R1095 B.n648 B.n39 163.367
R1096 B.n644 B.n39 163.367
R1097 B.n644 B.n643 163.367
R1098 B.n643 B.n642 163.367
R1099 B.n642 B.n41 163.367
R1100 B.n638 B.n41 163.367
R1101 B.n638 B.n637 163.367
R1102 B.n637 B.n636 163.367
R1103 B.n636 B.n43 163.367
R1104 B.n632 B.n43 163.367
R1105 B.n632 B.n631 163.367
R1106 B.n631 B.n630 163.367
R1107 B.n630 B.n45 163.367
R1108 B.n626 B.n45 163.367
R1109 B.n626 B.n625 163.367
R1110 B.n625 B.n49 163.367
R1111 B.n621 B.n49 163.367
R1112 B.n621 B.n620 163.367
R1113 B.n620 B.n619 163.367
R1114 B.n619 B.n51 163.367
R1115 B.n615 B.n51 163.367
R1116 B.n615 B.n614 163.367
R1117 B.n614 B.n613 163.367
R1118 B.n613 B.n53 163.367
R1119 B.n608 B.n53 163.367
R1120 B.n608 B.n607 163.367
R1121 B.n607 B.n606 163.367
R1122 B.n606 B.n57 163.367
R1123 B.n602 B.n57 163.367
R1124 B.n602 B.n601 163.367
R1125 B.n601 B.n600 163.367
R1126 B.n600 B.n59 163.367
R1127 B.n596 B.n59 163.367
R1128 B.n596 B.n595 163.367
R1129 B.n595 B.n594 163.367
R1130 B.n594 B.n61 163.367
R1131 B.n590 B.n61 163.367
R1132 B.n590 B.n589 163.367
R1133 B.n589 B.n588 163.367
R1134 B.n588 B.n63 163.367
R1135 B.n584 B.n63 163.367
R1136 B.n584 B.n583 163.367
R1137 B.n583 B.n582 163.367
R1138 B.n582 B.n65 163.367
R1139 B.n578 B.n65 163.367
R1140 B.n145 B.t1 120.26
R1141 B.n55 B.t8 120.26
R1142 B.n153 B.t4 120.257
R1143 B.n47 B.t11 120.257
R1144 B.n145 B.n144 64.9702
R1145 B.n153 B.n152 64.9702
R1146 B.n47 B.n46 64.9702
R1147 B.n55 B.n54 64.9702
R1148 B.n146 B.n145 59.5399
R1149 B.n328 B.n153 59.5399
R1150 B.n48 B.n47 59.5399
R1151 B.n610 B.n55 59.5399
R1152 B.n658 B.n657 34.8103
R1153 B.n579 B.n66 34.8103
R1154 B.n376 B.n375 34.8103
R1155 B.n297 B.n164 34.8103
R1156 B B.n759 18.0485
R1157 B.n657 B.n36 10.6151
R1158 B.n653 B.n36 10.6151
R1159 B.n653 B.n652 10.6151
R1160 B.n652 B.n651 10.6151
R1161 B.n651 B.n38 10.6151
R1162 B.n647 B.n38 10.6151
R1163 B.n647 B.n646 10.6151
R1164 B.n646 B.n645 10.6151
R1165 B.n645 B.n40 10.6151
R1166 B.n641 B.n40 10.6151
R1167 B.n641 B.n640 10.6151
R1168 B.n640 B.n639 10.6151
R1169 B.n639 B.n42 10.6151
R1170 B.n635 B.n42 10.6151
R1171 B.n635 B.n634 10.6151
R1172 B.n634 B.n633 10.6151
R1173 B.n633 B.n44 10.6151
R1174 B.n629 B.n44 10.6151
R1175 B.n629 B.n628 10.6151
R1176 B.n628 B.n627 10.6151
R1177 B.n624 B.n623 10.6151
R1178 B.n623 B.n622 10.6151
R1179 B.n622 B.n50 10.6151
R1180 B.n618 B.n50 10.6151
R1181 B.n618 B.n617 10.6151
R1182 B.n617 B.n616 10.6151
R1183 B.n616 B.n52 10.6151
R1184 B.n612 B.n52 10.6151
R1185 B.n612 B.n611 10.6151
R1186 B.n609 B.n56 10.6151
R1187 B.n605 B.n56 10.6151
R1188 B.n605 B.n604 10.6151
R1189 B.n604 B.n603 10.6151
R1190 B.n603 B.n58 10.6151
R1191 B.n599 B.n58 10.6151
R1192 B.n599 B.n598 10.6151
R1193 B.n598 B.n597 10.6151
R1194 B.n597 B.n60 10.6151
R1195 B.n593 B.n60 10.6151
R1196 B.n593 B.n592 10.6151
R1197 B.n592 B.n591 10.6151
R1198 B.n591 B.n62 10.6151
R1199 B.n587 B.n62 10.6151
R1200 B.n587 B.n586 10.6151
R1201 B.n586 B.n585 10.6151
R1202 B.n585 B.n64 10.6151
R1203 B.n581 B.n64 10.6151
R1204 B.n581 B.n580 10.6151
R1205 B.n580 B.n579 10.6151
R1206 B.n377 B.n376 10.6151
R1207 B.n377 B.n132 10.6151
R1208 B.n381 B.n132 10.6151
R1209 B.n382 B.n381 10.6151
R1210 B.n383 B.n382 10.6151
R1211 B.n383 B.n130 10.6151
R1212 B.n387 B.n130 10.6151
R1213 B.n388 B.n387 10.6151
R1214 B.n389 B.n388 10.6151
R1215 B.n389 B.n128 10.6151
R1216 B.n393 B.n128 10.6151
R1217 B.n394 B.n393 10.6151
R1218 B.n395 B.n394 10.6151
R1219 B.n395 B.n126 10.6151
R1220 B.n399 B.n126 10.6151
R1221 B.n400 B.n399 10.6151
R1222 B.n401 B.n400 10.6151
R1223 B.n401 B.n124 10.6151
R1224 B.n405 B.n124 10.6151
R1225 B.n406 B.n405 10.6151
R1226 B.n407 B.n406 10.6151
R1227 B.n407 B.n122 10.6151
R1228 B.n411 B.n122 10.6151
R1229 B.n412 B.n411 10.6151
R1230 B.n413 B.n412 10.6151
R1231 B.n413 B.n120 10.6151
R1232 B.n417 B.n120 10.6151
R1233 B.n418 B.n417 10.6151
R1234 B.n419 B.n418 10.6151
R1235 B.n419 B.n118 10.6151
R1236 B.n423 B.n118 10.6151
R1237 B.n424 B.n423 10.6151
R1238 B.n425 B.n424 10.6151
R1239 B.n425 B.n116 10.6151
R1240 B.n429 B.n116 10.6151
R1241 B.n430 B.n429 10.6151
R1242 B.n431 B.n430 10.6151
R1243 B.n431 B.n114 10.6151
R1244 B.n435 B.n114 10.6151
R1245 B.n436 B.n435 10.6151
R1246 B.n437 B.n436 10.6151
R1247 B.n437 B.n112 10.6151
R1248 B.n441 B.n112 10.6151
R1249 B.n442 B.n441 10.6151
R1250 B.n443 B.n442 10.6151
R1251 B.n443 B.n110 10.6151
R1252 B.n447 B.n110 10.6151
R1253 B.n448 B.n447 10.6151
R1254 B.n449 B.n448 10.6151
R1255 B.n449 B.n108 10.6151
R1256 B.n453 B.n108 10.6151
R1257 B.n454 B.n453 10.6151
R1258 B.n455 B.n454 10.6151
R1259 B.n455 B.n106 10.6151
R1260 B.n459 B.n106 10.6151
R1261 B.n460 B.n459 10.6151
R1262 B.n461 B.n460 10.6151
R1263 B.n461 B.n104 10.6151
R1264 B.n465 B.n104 10.6151
R1265 B.n466 B.n465 10.6151
R1266 B.n467 B.n466 10.6151
R1267 B.n467 B.n102 10.6151
R1268 B.n471 B.n102 10.6151
R1269 B.n472 B.n471 10.6151
R1270 B.n473 B.n472 10.6151
R1271 B.n473 B.n100 10.6151
R1272 B.n477 B.n100 10.6151
R1273 B.n478 B.n477 10.6151
R1274 B.n479 B.n478 10.6151
R1275 B.n479 B.n98 10.6151
R1276 B.n483 B.n98 10.6151
R1277 B.n484 B.n483 10.6151
R1278 B.n485 B.n484 10.6151
R1279 B.n485 B.n96 10.6151
R1280 B.n489 B.n96 10.6151
R1281 B.n490 B.n489 10.6151
R1282 B.n491 B.n490 10.6151
R1283 B.n491 B.n94 10.6151
R1284 B.n495 B.n94 10.6151
R1285 B.n496 B.n495 10.6151
R1286 B.n497 B.n496 10.6151
R1287 B.n497 B.n92 10.6151
R1288 B.n501 B.n92 10.6151
R1289 B.n502 B.n501 10.6151
R1290 B.n503 B.n502 10.6151
R1291 B.n503 B.n90 10.6151
R1292 B.n507 B.n90 10.6151
R1293 B.n508 B.n507 10.6151
R1294 B.n509 B.n508 10.6151
R1295 B.n509 B.n88 10.6151
R1296 B.n513 B.n88 10.6151
R1297 B.n514 B.n513 10.6151
R1298 B.n515 B.n514 10.6151
R1299 B.n515 B.n86 10.6151
R1300 B.n519 B.n86 10.6151
R1301 B.n520 B.n519 10.6151
R1302 B.n521 B.n520 10.6151
R1303 B.n521 B.n84 10.6151
R1304 B.n525 B.n84 10.6151
R1305 B.n526 B.n525 10.6151
R1306 B.n527 B.n526 10.6151
R1307 B.n527 B.n82 10.6151
R1308 B.n531 B.n82 10.6151
R1309 B.n532 B.n531 10.6151
R1310 B.n533 B.n532 10.6151
R1311 B.n533 B.n80 10.6151
R1312 B.n537 B.n80 10.6151
R1313 B.n538 B.n537 10.6151
R1314 B.n539 B.n538 10.6151
R1315 B.n539 B.n78 10.6151
R1316 B.n543 B.n78 10.6151
R1317 B.n544 B.n543 10.6151
R1318 B.n545 B.n544 10.6151
R1319 B.n545 B.n76 10.6151
R1320 B.n549 B.n76 10.6151
R1321 B.n550 B.n549 10.6151
R1322 B.n551 B.n550 10.6151
R1323 B.n551 B.n74 10.6151
R1324 B.n555 B.n74 10.6151
R1325 B.n556 B.n555 10.6151
R1326 B.n557 B.n556 10.6151
R1327 B.n557 B.n72 10.6151
R1328 B.n561 B.n72 10.6151
R1329 B.n562 B.n561 10.6151
R1330 B.n563 B.n562 10.6151
R1331 B.n563 B.n70 10.6151
R1332 B.n567 B.n70 10.6151
R1333 B.n568 B.n567 10.6151
R1334 B.n569 B.n568 10.6151
R1335 B.n569 B.n68 10.6151
R1336 B.n573 B.n68 10.6151
R1337 B.n574 B.n573 10.6151
R1338 B.n575 B.n574 10.6151
R1339 B.n575 B.n66 10.6151
R1340 B.n298 B.n297 10.6151
R1341 B.n299 B.n298 10.6151
R1342 B.n299 B.n162 10.6151
R1343 B.n303 B.n162 10.6151
R1344 B.n304 B.n303 10.6151
R1345 B.n305 B.n304 10.6151
R1346 B.n305 B.n160 10.6151
R1347 B.n309 B.n160 10.6151
R1348 B.n310 B.n309 10.6151
R1349 B.n311 B.n310 10.6151
R1350 B.n311 B.n158 10.6151
R1351 B.n315 B.n158 10.6151
R1352 B.n316 B.n315 10.6151
R1353 B.n317 B.n316 10.6151
R1354 B.n317 B.n156 10.6151
R1355 B.n321 B.n156 10.6151
R1356 B.n322 B.n321 10.6151
R1357 B.n323 B.n322 10.6151
R1358 B.n323 B.n154 10.6151
R1359 B.n327 B.n154 10.6151
R1360 B.n330 B.n329 10.6151
R1361 B.n330 B.n150 10.6151
R1362 B.n334 B.n150 10.6151
R1363 B.n335 B.n334 10.6151
R1364 B.n336 B.n335 10.6151
R1365 B.n336 B.n148 10.6151
R1366 B.n340 B.n148 10.6151
R1367 B.n341 B.n340 10.6151
R1368 B.n342 B.n341 10.6151
R1369 B.n346 B.n345 10.6151
R1370 B.n347 B.n346 10.6151
R1371 B.n347 B.n142 10.6151
R1372 B.n351 B.n142 10.6151
R1373 B.n352 B.n351 10.6151
R1374 B.n353 B.n352 10.6151
R1375 B.n353 B.n140 10.6151
R1376 B.n357 B.n140 10.6151
R1377 B.n358 B.n357 10.6151
R1378 B.n359 B.n358 10.6151
R1379 B.n359 B.n138 10.6151
R1380 B.n363 B.n138 10.6151
R1381 B.n364 B.n363 10.6151
R1382 B.n365 B.n364 10.6151
R1383 B.n365 B.n136 10.6151
R1384 B.n369 B.n136 10.6151
R1385 B.n370 B.n369 10.6151
R1386 B.n371 B.n370 10.6151
R1387 B.n371 B.n134 10.6151
R1388 B.n375 B.n134 10.6151
R1389 B.n293 B.n164 10.6151
R1390 B.n293 B.n292 10.6151
R1391 B.n292 B.n291 10.6151
R1392 B.n291 B.n166 10.6151
R1393 B.n287 B.n166 10.6151
R1394 B.n287 B.n286 10.6151
R1395 B.n286 B.n285 10.6151
R1396 B.n285 B.n168 10.6151
R1397 B.n281 B.n168 10.6151
R1398 B.n281 B.n280 10.6151
R1399 B.n280 B.n279 10.6151
R1400 B.n279 B.n170 10.6151
R1401 B.n275 B.n170 10.6151
R1402 B.n275 B.n274 10.6151
R1403 B.n274 B.n273 10.6151
R1404 B.n273 B.n172 10.6151
R1405 B.n269 B.n172 10.6151
R1406 B.n269 B.n268 10.6151
R1407 B.n268 B.n267 10.6151
R1408 B.n267 B.n174 10.6151
R1409 B.n263 B.n174 10.6151
R1410 B.n263 B.n262 10.6151
R1411 B.n262 B.n261 10.6151
R1412 B.n261 B.n176 10.6151
R1413 B.n257 B.n176 10.6151
R1414 B.n257 B.n256 10.6151
R1415 B.n256 B.n255 10.6151
R1416 B.n255 B.n178 10.6151
R1417 B.n251 B.n178 10.6151
R1418 B.n251 B.n250 10.6151
R1419 B.n250 B.n249 10.6151
R1420 B.n249 B.n180 10.6151
R1421 B.n245 B.n180 10.6151
R1422 B.n245 B.n244 10.6151
R1423 B.n244 B.n243 10.6151
R1424 B.n243 B.n182 10.6151
R1425 B.n239 B.n182 10.6151
R1426 B.n239 B.n238 10.6151
R1427 B.n238 B.n237 10.6151
R1428 B.n237 B.n184 10.6151
R1429 B.n233 B.n184 10.6151
R1430 B.n233 B.n232 10.6151
R1431 B.n232 B.n231 10.6151
R1432 B.n231 B.n186 10.6151
R1433 B.n227 B.n186 10.6151
R1434 B.n227 B.n226 10.6151
R1435 B.n226 B.n225 10.6151
R1436 B.n225 B.n188 10.6151
R1437 B.n221 B.n188 10.6151
R1438 B.n221 B.n220 10.6151
R1439 B.n220 B.n219 10.6151
R1440 B.n219 B.n190 10.6151
R1441 B.n215 B.n190 10.6151
R1442 B.n215 B.n214 10.6151
R1443 B.n214 B.n213 10.6151
R1444 B.n213 B.n192 10.6151
R1445 B.n209 B.n192 10.6151
R1446 B.n209 B.n208 10.6151
R1447 B.n208 B.n207 10.6151
R1448 B.n207 B.n194 10.6151
R1449 B.n203 B.n194 10.6151
R1450 B.n203 B.n202 10.6151
R1451 B.n202 B.n201 10.6151
R1452 B.n201 B.n196 10.6151
R1453 B.n197 B.n196 10.6151
R1454 B.n197 B.n0 10.6151
R1455 B.n755 B.n1 10.6151
R1456 B.n755 B.n754 10.6151
R1457 B.n754 B.n753 10.6151
R1458 B.n753 B.n4 10.6151
R1459 B.n749 B.n4 10.6151
R1460 B.n749 B.n748 10.6151
R1461 B.n748 B.n747 10.6151
R1462 B.n747 B.n6 10.6151
R1463 B.n743 B.n6 10.6151
R1464 B.n743 B.n742 10.6151
R1465 B.n742 B.n741 10.6151
R1466 B.n741 B.n8 10.6151
R1467 B.n737 B.n8 10.6151
R1468 B.n737 B.n736 10.6151
R1469 B.n736 B.n735 10.6151
R1470 B.n735 B.n10 10.6151
R1471 B.n731 B.n10 10.6151
R1472 B.n731 B.n730 10.6151
R1473 B.n730 B.n729 10.6151
R1474 B.n729 B.n12 10.6151
R1475 B.n725 B.n12 10.6151
R1476 B.n725 B.n724 10.6151
R1477 B.n724 B.n723 10.6151
R1478 B.n723 B.n14 10.6151
R1479 B.n719 B.n14 10.6151
R1480 B.n719 B.n718 10.6151
R1481 B.n718 B.n717 10.6151
R1482 B.n717 B.n16 10.6151
R1483 B.n713 B.n16 10.6151
R1484 B.n713 B.n712 10.6151
R1485 B.n712 B.n711 10.6151
R1486 B.n711 B.n18 10.6151
R1487 B.n707 B.n18 10.6151
R1488 B.n707 B.n706 10.6151
R1489 B.n706 B.n705 10.6151
R1490 B.n705 B.n20 10.6151
R1491 B.n701 B.n20 10.6151
R1492 B.n701 B.n700 10.6151
R1493 B.n700 B.n699 10.6151
R1494 B.n699 B.n22 10.6151
R1495 B.n695 B.n22 10.6151
R1496 B.n695 B.n694 10.6151
R1497 B.n694 B.n693 10.6151
R1498 B.n693 B.n24 10.6151
R1499 B.n689 B.n24 10.6151
R1500 B.n689 B.n688 10.6151
R1501 B.n688 B.n687 10.6151
R1502 B.n687 B.n26 10.6151
R1503 B.n683 B.n26 10.6151
R1504 B.n683 B.n682 10.6151
R1505 B.n682 B.n681 10.6151
R1506 B.n681 B.n28 10.6151
R1507 B.n677 B.n28 10.6151
R1508 B.n677 B.n676 10.6151
R1509 B.n676 B.n675 10.6151
R1510 B.n675 B.n30 10.6151
R1511 B.n671 B.n30 10.6151
R1512 B.n671 B.n670 10.6151
R1513 B.n670 B.n669 10.6151
R1514 B.n669 B.n32 10.6151
R1515 B.n665 B.n32 10.6151
R1516 B.n665 B.n664 10.6151
R1517 B.n664 B.n663 10.6151
R1518 B.n663 B.n34 10.6151
R1519 B.n659 B.n34 10.6151
R1520 B.n659 B.n658 10.6151
R1521 B.n627 B.n48 9.36635
R1522 B.n610 B.n609 9.36635
R1523 B.n328 B.n327 9.36635
R1524 B.n345 B.n146 9.36635
R1525 B.n759 B.n0 2.81026
R1526 B.n759 B.n1 2.81026
R1527 B.n624 B.n48 1.24928
R1528 B.n611 B.n610 1.24928
R1529 B.n329 B.n328 1.24928
R1530 B.n342 B.n146 1.24928
C0 VDD2 w_n4990_n1980# 2.63413f
C1 VN VP 7.72542f
C2 VTAIL VP 6.336339f
C3 B w_n4990_n1980# 9.32228f
C4 VTAIL VN 6.32217f
C5 VDD1 VP 5.41406f
C6 VDD1 VN 0.154651f
C7 VDD2 VP 0.641338f
C8 VDD2 VN 4.93469f
C9 VDD1 VTAIL 7.55561f
C10 VDD2 VTAIL 7.611169f
C11 VDD2 VDD1 2.44722f
C12 VP B 2.46122f
C13 VN B 1.36432f
C14 VTAIL B 2.27905f
C15 VDD1 B 2.09113f
C16 VDD2 B 2.22553f
C17 VP w_n4990_n1980# 11.3262f
C18 VN w_n4990_n1980# 10.6753f
C19 VTAIL w_n4990_n1980# 2.30512f
C20 VDD1 w_n4990_n1980# 2.46902f
C21 VDD2 VSUBS 2.228813f
C22 VDD1 VSUBS 1.977834f
C23 VTAIL VSUBS 0.70195f
C24 VN VSUBS 8.10526f
C25 VP VSUBS 4.205382f
C26 B VSUBS 4.983951f
C27 w_n4990_n1980# VSUBS 0.123772p
C28 B.n0 VSUBS 0.007882f
C29 B.n1 VSUBS 0.007882f
C30 B.n2 VSUBS 0.012465f
C31 B.n3 VSUBS 0.012465f
C32 B.n4 VSUBS 0.012465f
C33 B.n5 VSUBS 0.012465f
C34 B.n6 VSUBS 0.012465f
C35 B.n7 VSUBS 0.012465f
C36 B.n8 VSUBS 0.012465f
C37 B.n9 VSUBS 0.012465f
C38 B.n10 VSUBS 0.012465f
C39 B.n11 VSUBS 0.012465f
C40 B.n12 VSUBS 0.012465f
C41 B.n13 VSUBS 0.012465f
C42 B.n14 VSUBS 0.012465f
C43 B.n15 VSUBS 0.012465f
C44 B.n16 VSUBS 0.012465f
C45 B.n17 VSUBS 0.012465f
C46 B.n18 VSUBS 0.012465f
C47 B.n19 VSUBS 0.012465f
C48 B.n20 VSUBS 0.012465f
C49 B.n21 VSUBS 0.012465f
C50 B.n22 VSUBS 0.012465f
C51 B.n23 VSUBS 0.012465f
C52 B.n24 VSUBS 0.012465f
C53 B.n25 VSUBS 0.012465f
C54 B.n26 VSUBS 0.012465f
C55 B.n27 VSUBS 0.012465f
C56 B.n28 VSUBS 0.012465f
C57 B.n29 VSUBS 0.012465f
C58 B.n30 VSUBS 0.012465f
C59 B.n31 VSUBS 0.012465f
C60 B.n32 VSUBS 0.012465f
C61 B.n33 VSUBS 0.012465f
C62 B.n34 VSUBS 0.012465f
C63 B.n35 VSUBS 0.029503f
C64 B.n36 VSUBS 0.012465f
C65 B.n37 VSUBS 0.012465f
C66 B.n38 VSUBS 0.012465f
C67 B.n39 VSUBS 0.012465f
C68 B.n40 VSUBS 0.012465f
C69 B.n41 VSUBS 0.012465f
C70 B.n42 VSUBS 0.012465f
C71 B.n43 VSUBS 0.012465f
C72 B.n44 VSUBS 0.012465f
C73 B.n45 VSUBS 0.012465f
C74 B.t11 VSUBS 0.252025f
C75 B.t10 VSUBS 0.290859f
C76 B.t9 VSUBS 1.30498f
C77 B.n46 VSUBS 0.192529f
C78 B.n47 VSUBS 0.128494f
C79 B.n48 VSUBS 0.028881f
C80 B.n49 VSUBS 0.012465f
C81 B.n50 VSUBS 0.012465f
C82 B.n51 VSUBS 0.012465f
C83 B.n52 VSUBS 0.012465f
C84 B.n53 VSUBS 0.012465f
C85 B.t8 VSUBS 0.252025f
C86 B.t7 VSUBS 0.290858f
C87 B.t6 VSUBS 1.30498f
C88 B.n54 VSUBS 0.19253f
C89 B.n55 VSUBS 0.128494f
C90 B.n56 VSUBS 0.012465f
C91 B.n57 VSUBS 0.012465f
C92 B.n58 VSUBS 0.012465f
C93 B.n59 VSUBS 0.012465f
C94 B.n60 VSUBS 0.012465f
C95 B.n61 VSUBS 0.012465f
C96 B.n62 VSUBS 0.012465f
C97 B.n63 VSUBS 0.012465f
C98 B.n64 VSUBS 0.012465f
C99 B.n65 VSUBS 0.012465f
C100 B.n66 VSUBS 0.030885f
C101 B.n67 VSUBS 0.012465f
C102 B.n68 VSUBS 0.012465f
C103 B.n69 VSUBS 0.012465f
C104 B.n70 VSUBS 0.012465f
C105 B.n71 VSUBS 0.012465f
C106 B.n72 VSUBS 0.012465f
C107 B.n73 VSUBS 0.012465f
C108 B.n74 VSUBS 0.012465f
C109 B.n75 VSUBS 0.012465f
C110 B.n76 VSUBS 0.012465f
C111 B.n77 VSUBS 0.012465f
C112 B.n78 VSUBS 0.012465f
C113 B.n79 VSUBS 0.012465f
C114 B.n80 VSUBS 0.012465f
C115 B.n81 VSUBS 0.012465f
C116 B.n82 VSUBS 0.012465f
C117 B.n83 VSUBS 0.012465f
C118 B.n84 VSUBS 0.012465f
C119 B.n85 VSUBS 0.012465f
C120 B.n86 VSUBS 0.012465f
C121 B.n87 VSUBS 0.012465f
C122 B.n88 VSUBS 0.012465f
C123 B.n89 VSUBS 0.012465f
C124 B.n90 VSUBS 0.012465f
C125 B.n91 VSUBS 0.012465f
C126 B.n92 VSUBS 0.012465f
C127 B.n93 VSUBS 0.012465f
C128 B.n94 VSUBS 0.012465f
C129 B.n95 VSUBS 0.012465f
C130 B.n96 VSUBS 0.012465f
C131 B.n97 VSUBS 0.012465f
C132 B.n98 VSUBS 0.012465f
C133 B.n99 VSUBS 0.012465f
C134 B.n100 VSUBS 0.012465f
C135 B.n101 VSUBS 0.012465f
C136 B.n102 VSUBS 0.012465f
C137 B.n103 VSUBS 0.012465f
C138 B.n104 VSUBS 0.012465f
C139 B.n105 VSUBS 0.012465f
C140 B.n106 VSUBS 0.012465f
C141 B.n107 VSUBS 0.012465f
C142 B.n108 VSUBS 0.012465f
C143 B.n109 VSUBS 0.012465f
C144 B.n110 VSUBS 0.012465f
C145 B.n111 VSUBS 0.012465f
C146 B.n112 VSUBS 0.012465f
C147 B.n113 VSUBS 0.012465f
C148 B.n114 VSUBS 0.012465f
C149 B.n115 VSUBS 0.012465f
C150 B.n116 VSUBS 0.012465f
C151 B.n117 VSUBS 0.012465f
C152 B.n118 VSUBS 0.012465f
C153 B.n119 VSUBS 0.012465f
C154 B.n120 VSUBS 0.012465f
C155 B.n121 VSUBS 0.012465f
C156 B.n122 VSUBS 0.012465f
C157 B.n123 VSUBS 0.012465f
C158 B.n124 VSUBS 0.012465f
C159 B.n125 VSUBS 0.012465f
C160 B.n126 VSUBS 0.012465f
C161 B.n127 VSUBS 0.012465f
C162 B.n128 VSUBS 0.012465f
C163 B.n129 VSUBS 0.012465f
C164 B.n130 VSUBS 0.012465f
C165 B.n131 VSUBS 0.012465f
C166 B.n132 VSUBS 0.012465f
C167 B.n133 VSUBS 0.029503f
C168 B.n134 VSUBS 0.012465f
C169 B.n135 VSUBS 0.012465f
C170 B.n136 VSUBS 0.012465f
C171 B.n137 VSUBS 0.012465f
C172 B.n138 VSUBS 0.012465f
C173 B.n139 VSUBS 0.012465f
C174 B.n140 VSUBS 0.012465f
C175 B.n141 VSUBS 0.012465f
C176 B.n142 VSUBS 0.012465f
C177 B.n143 VSUBS 0.012465f
C178 B.t1 VSUBS 0.252025f
C179 B.t2 VSUBS 0.290858f
C180 B.t0 VSUBS 1.30498f
C181 B.n144 VSUBS 0.19253f
C182 B.n145 VSUBS 0.128494f
C183 B.n146 VSUBS 0.028881f
C184 B.n147 VSUBS 0.012465f
C185 B.n148 VSUBS 0.012465f
C186 B.n149 VSUBS 0.012465f
C187 B.n150 VSUBS 0.012465f
C188 B.n151 VSUBS 0.012465f
C189 B.t4 VSUBS 0.252025f
C190 B.t5 VSUBS 0.290859f
C191 B.t3 VSUBS 1.30498f
C192 B.n152 VSUBS 0.192529f
C193 B.n153 VSUBS 0.128494f
C194 B.n154 VSUBS 0.012465f
C195 B.n155 VSUBS 0.012465f
C196 B.n156 VSUBS 0.012465f
C197 B.n157 VSUBS 0.012465f
C198 B.n158 VSUBS 0.012465f
C199 B.n159 VSUBS 0.012465f
C200 B.n160 VSUBS 0.012465f
C201 B.n161 VSUBS 0.012465f
C202 B.n162 VSUBS 0.012465f
C203 B.n163 VSUBS 0.012465f
C204 B.n164 VSUBS 0.029503f
C205 B.n165 VSUBS 0.012465f
C206 B.n166 VSUBS 0.012465f
C207 B.n167 VSUBS 0.012465f
C208 B.n168 VSUBS 0.012465f
C209 B.n169 VSUBS 0.012465f
C210 B.n170 VSUBS 0.012465f
C211 B.n171 VSUBS 0.012465f
C212 B.n172 VSUBS 0.012465f
C213 B.n173 VSUBS 0.012465f
C214 B.n174 VSUBS 0.012465f
C215 B.n175 VSUBS 0.012465f
C216 B.n176 VSUBS 0.012465f
C217 B.n177 VSUBS 0.012465f
C218 B.n178 VSUBS 0.012465f
C219 B.n179 VSUBS 0.012465f
C220 B.n180 VSUBS 0.012465f
C221 B.n181 VSUBS 0.012465f
C222 B.n182 VSUBS 0.012465f
C223 B.n183 VSUBS 0.012465f
C224 B.n184 VSUBS 0.012465f
C225 B.n185 VSUBS 0.012465f
C226 B.n186 VSUBS 0.012465f
C227 B.n187 VSUBS 0.012465f
C228 B.n188 VSUBS 0.012465f
C229 B.n189 VSUBS 0.012465f
C230 B.n190 VSUBS 0.012465f
C231 B.n191 VSUBS 0.012465f
C232 B.n192 VSUBS 0.012465f
C233 B.n193 VSUBS 0.012465f
C234 B.n194 VSUBS 0.012465f
C235 B.n195 VSUBS 0.012465f
C236 B.n196 VSUBS 0.012465f
C237 B.n197 VSUBS 0.012465f
C238 B.n198 VSUBS 0.012465f
C239 B.n199 VSUBS 0.012465f
C240 B.n200 VSUBS 0.012465f
C241 B.n201 VSUBS 0.012465f
C242 B.n202 VSUBS 0.012465f
C243 B.n203 VSUBS 0.012465f
C244 B.n204 VSUBS 0.012465f
C245 B.n205 VSUBS 0.012465f
C246 B.n206 VSUBS 0.012465f
C247 B.n207 VSUBS 0.012465f
C248 B.n208 VSUBS 0.012465f
C249 B.n209 VSUBS 0.012465f
C250 B.n210 VSUBS 0.012465f
C251 B.n211 VSUBS 0.012465f
C252 B.n212 VSUBS 0.012465f
C253 B.n213 VSUBS 0.012465f
C254 B.n214 VSUBS 0.012465f
C255 B.n215 VSUBS 0.012465f
C256 B.n216 VSUBS 0.012465f
C257 B.n217 VSUBS 0.012465f
C258 B.n218 VSUBS 0.012465f
C259 B.n219 VSUBS 0.012465f
C260 B.n220 VSUBS 0.012465f
C261 B.n221 VSUBS 0.012465f
C262 B.n222 VSUBS 0.012465f
C263 B.n223 VSUBS 0.012465f
C264 B.n224 VSUBS 0.012465f
C265 B.n225 VSUBS 0.012465f
C266 B.n226 VSUBS 0.012465f
C267 B.n227 VSUBS 0.012465f
C268 B.n228 VSUBS 0.012465f
C269 B.n229 VSUBS 0.012465f
C270 B.n230 VSUBS 0.012465f
C271 B.n231 VSUBS 0.012465f
C272 B.n232 VSUBS 0.012465f
C273 B.n233 VSUBS 0.012465f
C274 B.n234 VSUBS 0.012465f
C275 B.n235 VSUBS 0.012465f
C276 B.n236 VSUBS 0.012465f
C277 B.n237 VSUBS 0.012465f
C278 B.n238 VSUBS 0.012465f
C279 B.n239 VSUBS 0.012465f
C280 B.n240 VSUBS 0.012465f
C281 B.n241 VSUBS 0.012465f
C282 B.n242 VSUBS 0.012465f
C283 B.n243 VSUBS 0.012465f
C284 B.n244 VSUBS 0.012465f
C285 B.n245 VSUBS 0.012465f
C286 B.n246 VSUBS 0.012465f
C287 B.n247 VSUBS 0.012465f
C288 B.n248 VSUBS 0.012465f
C289 B.n249 VSUBS 0.012465f
C290 B.n250 VSUBS 0.012465f
C291 B.n251 VSUBS 0.012465f
C292 B.n252 VSUBS 0.012465f
C293 B.n253 VSUBS 0.012465f
C294 B.n254 VSUBS 0.012465f
C295 B.n255 VSUBS 0.012465f
C296 B.n256 VSUBS 0.012465f
C297 B.n257 VSUBS 0.012465f
C298 B.n258 VSUBS 0.012465f
C299 B.n259 VSUBS 0.012465f
C300 B.n260 VSUBS 0.012465f
C301 B.n261 VSUBS 0.012465f
C302 B.n262 VSUBS 0.012465f
C303 B.n263 VSUBS 0.012465f
C304 B.n264 VSUBS 0.012465f
C305 B.n265 VSUBS 0.012465f
C306 B.n266 VSUBS 0.012465f
C307 B.n267 VSUBS 0.012465f
C308 B.n268 VSUBS 0.012465f
C309 B.n269 VSUBS 0.012465f
C310 B.n270 VSUBS 0.012465f
C311 B.n271 VSUBS 0.012465f
C312 B.n272 VSUBS 0.012465f
C313 B.n273 VSUBS 0.012465f
C314 B.n274 VSUBS 0.012465f
C315 B.n275 VSUBS 0.012465f
C316 B.n276 VSUBS 0.012465f
C317 B.n277 VSUBS 0.012465f
C318 B.n278 VSUBS 0.012465f
C319 B.n279 VSUBS 0.012465f
C320 B.n280 VSUBS 0.012465f
C321 B.n281 VSUBS 0.012465f
C322 B.n282 VSUBS 0.012465f
C323 B.n283 VSUBS 0.012465f
C324 B.n284 VSUBS 0.012465f
C325 B.n285 VSUBS 0.012465f
C326 B.n286 VSUBS 0.012465f
C327 B.n287 VSUBS 0.012465f
C328 B.n288 VSUBS 0.012465f
C329 B.n289 VSUBS 0.012465f
C330 B.n290 VSUBS 0.012465f
C331 B.n291 VSUBS 0.012465f
C332 B.n292 VSUBS 0.012465f
C333 B.n293 VSUBS 0.012465f
C334 B.n294 VSUBS 0.012465f
C335 B.n295 VSUBS 0.029503f
C336 B.n296 VSUBS 0.031357f
C337 B.n297 VSUBS 0.031357f
C338 B.n298 VSUBS 0.012465f
C339 B.n299 VSUBS 0.012465f
C340 B.n300 VSUBS 0.012465f
C341 B.n301 VSUBS 0.012465f
C342 B.n302 VSUBS 0.012465f
C343 B.n303 VSUBS 0.012465f
C344 B.n304 VSUBS 0.012465f
C345 B.n305 VSUBS 0.012465f
C346 B.n306 VSUBS 0.012465f
C347 B.n307 VSUBS 0.012465f
C348 B.n308 VSUBS 0.012465f
C349 B.n309 VSUBS 0.012465f
C350 B.n310 VSUBS 0.012465f
C351 B.n311 VSUBS 0.012465f
C352 B.n312 VSUBS 0.012465f
C353 B.n313 VSUBS 0.012465f
C354 B.n314 VSUBS 0.012465f
C355 B.n315 VSUBS 0.012465f
C356 B.n316 VSUBS 0.012465f
C357 B.n317 VSUBS 0.012465f
C358 B.n318 VSUBS 0.012465f
C359 B.n319 VSUBS 0.012465f
C360 B.n320 VSUBS 0.012465f
C361 B.n321 VSUBS 0.012465f
C362 B.n322 VSUBS 0.012465f
C363 B.n323 VSUBS 0.012465f
C364 B.n324 VSUBS 0.012465f
C365 B.n325 VSUBS 0.012465f
C366 B.n326 VSUBS 0.012465f
C367 B.n327 VSUBS 0.011732f
C368 B.n328 VSUBS 0.028881f
C369 B.n329 VSUBS 0.006966f
C370 B.n330 VSUBS 0.012465f
C371 B.n331 VSUBS 0.012465f
C372 B.n332 VSUBS 0.012465f
C373 B.n333 VSUBS 0.012465f
C374 B.n334 VSUBS 0.012465f
C375 B.n335 VSUBS 0.012465f
C376 B.n336 VSUBS 0.012465f
C377 B.n337 VSUBS 0.012465f
C378 B.n338 VSUBS 0.012465f
C379 B.n339 VSUBS 0.012465f
C380 B.n340 VSUBS 0.012465f
C381 B.n341 VSUBS 0.012465f
C382 B.n342 VSUBS 0.006966f
C383 B.n343 VSUBS 0.012465f
C384 B.n344 VSUBS 0.012465f
C385 B.n345 VSUBS 0.011732f
C386 B.n346 VSUBS 0.012465f
C387 B.n347 VSUBS 0.012465f
C388 B.n348 VSUBS 0.012465f
C389 B.n349 VSUBS 0.012465f
C390 B.n350 VSUBS 0.012465f
C391 B.n351 VSUBS 0.012465f
C392 B.n352 VSUBS 0.012465f
C393 B.n353 VSUBS 0.012465f
C394 B.n354 VSUBS 0.012465f
C395 B.n355 VSUBS 0.012465f
C396 B.n356 VSUBS 0.012465f
C397 B.n357 VSUBS 0.012465f
C398 B.n358 VSUBS 0.012465f
C399 B.n359 VSUBS 0.012465f
C400 B.n360 VSUBS 0.012465f
C401 B.n361 VSUBS 0.012465f
C402 B.n362 VSUBS 0.012465f
C403 B.n363 VSUBS 0.012465f
C404 B.n364 VSUBS 0.012465f
C405 B.n365 VSUBS 0.012465f
C406 B.n366 VSUBS 0.012465f
C407 B.n367 VSUBS 0.012465f
C408 B.n368 VSUBS 0.012465f
C409 B.n369 VSUBS 0.012465f
C410 B.n370 VSUBS 0.012465f
C411 B.n371 VSUBS 0.012465f
C412 B.n372 VSUBS 0.012465f
C413 B.n373 VSUBS 0.012465f
C414 B.n374 VSUBS 0.031357f
C415 B.n375 VSUBS 0.031357f
C416 B.n376 VSUBS 0.029503f
C417 B.n377 VSUBS 0.012465f
C418 B.n378 VSUBS 0.012465f
C419 B.n379 VSUBS 0.012465f
C420 B.n380 VSUBS 0.012465f
C421 B.n381 VSUBS 0.012465f
C422 B.n382 VSUBS 0.012465f
C423 B.n383 VSUBS 0.012465f
C424 B.n384 VSUBS 0.012465f
C425 B.n385 VSUBS 0.012465f
C426 B.n386 VSUBS 0.012465f
C427 B.n387 VSUBS 0.012465f
C428 B.n388 VSUBS 0.012465f
C429 B.n389 VSUBS 0.012465f
C430 B.n390 VSUBS 0.012465f
C431 B.n391 VSUBS 0.012465f
C432 B.n392 VSUBS 0.012465f
C433 B.n393 VSUBS 0.012465f
C434 B.n394 VSUBS 0.012465f
C435 B.n395 VSUBS 0.012465f
C436 B.n396 VSUBS 0.012465f
C437 B.n397 VSUBS 0.012465f
C438 B.n398 VSUBS 0.012465f
C439 B.n399 VSUBS 0.012465f
C440 B.n400 VSUBS 0.012465f
C441 B.n401 VSUBS 0.012465f
C442 B.n402 VSUBS 0.012465f
C443 B.n403 VSUBS 0.012465f
C444 B.n404 VSUBS 0.012465f
C445 B.n405 VSUBS 0.012465f
C446 B.n406 VSUBS 0.012465f
C447 B.n407 VSUBS 0.012465f
C448 B.n408 VSUBS 0.012465f
C449 B.n409 VSUBS 0.012465f
C450 B.n410 VSUBS 0.012465f
C451 B.n411 VSUBS 0.012465f
C452 B.n412 VSUBS 0.012465f
C453 B.n413 VSUBS 0.012465f
C454 B.n414 VSUBS 0.012465f
C455 B.n415 VSUBS 0.012465f
C456 B.n416 VSUBS 0.012465f
C457 B.n417 VSUBS 0.012465f
C458 B.n418 VSUBS 0.012465f
C459 B.n419 VSUBS 0.012465f
C460 B.n420 VSUBS 0.012465f
C461 B.n421 VSUBS 0.012465f
C462 B.n422 VSUBS 0.012465f
C463 B.n423 VSUBS 0.012465f
C464 B.n424 VSUBS 0.012465f
C465 B.n425 VSUBS 0.012465f
C466 B.n426 VSUBS 0.012465f
C467 B.n427 VSUBS 0.012465f
C468 B.n428 VSUBS 0.012465f
C469 B.n429 VSUBS 0.012465f
C470 B.n430 VSUBS 0.012465f
C471 B.n431 VSUBS 0.012465f
C472 B.n432 VSUBS 0.012465f
C473 B.n433 VSUBS 0.012465f
C474 B.n434 VSUBS 0.012465f
C475 B.n435 VSUBS 0.012465f
C476 B.n436 VSUBS 0.012465f
C477 B.n437 VSUBS 0.012465f
C478 B.n438 VSUBS 0.012465f
C479 B.n439 VSUBS 0.012465f
C480 B.n440 VSUBS 0.012465f
C481 B.n441 VSUBS 0.012465f
C482 B.n442 VSUBS 0.012465f
C483 B.n443 VSUBS 0.012465f
C484 B.n444 VSUBS 0.012465f
C485 B.n445 VSUBS 0.012465f
C486 B.n446 VSUBS 0.012465f
C487 B.n447 VSUBS 0.012465f
C488 B.n448 VSUBS 0.012465f
C489 B.n449 VSUBS 0.012465f
C490 B.n450 VSUBS 0.012465f
C491 B.n451 VSUBS 0.012465f
C492 B.n452 VSUBS 0.012465f
C493 B.n453 VSUBS 0.012465f
C494 B.n454 VSUBS 0.012465f
C495 B.n455 VSUBS 0.012465f
C496 B.n456 VSUBS 0.012465f
C497 B.n457 VSUBS 0.012465f
C498 B.n458 VSUBS 0.012465f
C499 B.n459 VSUBS 0.012465f
C500 B.n460 VSUBS 0.012465f
C501 B.n461 VSUBS 0.012465f
C502 B.n462 VSUBS 0.012465f
C503 B.n463 VSUBS 0.012465f
C504 B.n464 VSUBS 0.012465f
C505 B.n465 VSUBS 0.012465f
C506 B.n466 VSUBS 0.012465f
C507 B.n467 VSUBS 0.012465f
C508 B.n468 VSUBS 0.012465f
C509 B.n469 VSUBS 0.012465f
C510 B.n470 VSUBS 0.012465f
C511 B.n471 VSUBS 0.012465f
C512 B.n472 VSUBS 0.012465f
C513 B.n473 VSUBS 0.012465f
C514 B.n474 VSUBS 0.012465f
C515 B.n475 VSUBS 0.012465f
C516 B.n476 VSUBS 0.012465f
C517 B.n477 VSUBS 0.012465f
C518 B.n478 VSUBS 0.012465f
C519 B.n479 VSUBS 0.012465f
C520 B.n480 VSUBS 0.012465f
C521 B.n481 VSUBS 0.012465f
C522 B.n482 VSUBS 0.012465f
C523 B.n483 VSUBS 0.012465f
C524 B.n484 VSUBS 0.012465f
C525 B.n485 VSUBS 0.012465f
C526 B.n486 VSUBS 0.012465f
C527 B.n487 VSUBS 0.012465f
C528 B.n488 VSUBS 0.012465f
C529 B.n489 VSUBS 0.012465f
C530 B.n490 VSUBS 0.012465f
C531 B.n491 VSUBS 0.012465f
C532 B.n492 VSUBS 0.012465f
C533 B.n493 VSUBS 0.012465f
C534 B.n494 VSUBS 0.012465f
C535 B.n495 VSUBS 0.012465f
C536 B.n496 VSUBS 0.012465f
C537 B.n497 VSUBS 0.012465f
C538 B.n498 VSUBS 0.012465f
C539 B.n499 VSUBS 0.012465f
C540 B.n500 VSUBS 0.012465f
C541 B.n501 VSUBS 0.012465f
C542 B.n502 VSUBS 0.012465f
C543 B.n503 VSUBS 0.012465f
C544 B.n504 VSUBS 0.012465f
C545 B.n505 VSUBS 0.012465f
C546 B.n506 VSUBS 0.012465f
C547 B.n507 VSUBS 0.012465f
C548 B.n508 VSUBS 0.012465f
C549 B.n509 VSUBS 0.012465f
C550 B.n510 VSUBS 0.012465f
C551 B.n511 VSUBS 0.012465f
C552 B.n512 VSUBS 0.012465f
C553 B.n513 VSUBS 0.012465f
C554 B.n514 VSUBS 0.012465f
C555 B.n515 VSUBS 0.012465f
C556 B.n516 VSUBS 0.012465f
C557 B.n517 VSUBS 0.012465f
C558 B.n518 VSUBS 0.012465f
C559 B.n519 VSUBS 0.012465f
C560 B.n520 VSUBS 0.012465f
C561 B.n521 VSUBS 0.012465f
C562 B.n522 VSUBS 0.012465f
C563 B.n523 VSUBS 0.012465f
C564 B.n524 VSUBS 0.012465f
C565 B.n525 VSUBS 0.012465f
C566 B.n526 VSUBS 0.012465f
C567 B.n527 VSUBS 0.012465f
C568 B.n528 VSUBS 0.012465f
C569 B.n529 VSUBS 0.012465f
C570 B.n530 VSUBS 0.012465f
C571 B.n531 VSUBS 0.012465f
C572 B.n532 VSUBS 0.012465f
C573 B.n533 VSUBS 0.012465f
C574 B.n534 VSUBS 0.012465f
C575 B.n535 VSUBS 0.012465f
C576 B.n536 VSUBS 0.012465f
C577 B.n537 VSUBS 0.012465f
C578 B.n538 VSUBS 0.012465f
C579 B.n539 VSUBS 0.012465f
C580 B.n540 VSUBS 0.012465f
C581 B.n541 VSUBS 0.012465f
C582 B.n542 VSUBS 0.012465f
C583 B.n543 VSUBS 0.012465f
C584 B.n544 VSUBS 0.012465f
C585 B.n545 VSUBS 0.012465f
C586 B.n546 VSUBS 0.012465f
C587 B.n547 VSUBS 0.012465f
C588 B.n548 VSUBS 0.012465f
C589 B.n549 VSUBS 0.012465f
C590 B.n550 VSUBS 0.012465f
C591 B.n551 VSUBS 0.012465f
C592 B.n552 VSUBS 0.012465f
C593 B.n553 VSUBS 0.012465f
C594 B.n554 VSUBS 0.012465f
C595 B.n555 VSUBS 0.012465f
C596 B.n556 VSUBS 0.012465f
C597 B.n557 VSUBS 0.012465f
C598 B.n558 VSUBS 0.012465f
C599 B.n559 VSUBS 0.012465f
C600 B.n560 VSUBS 0.012465f
C601 B.n561 VSUBS 0.012465f
C602 B.n562 VSUBS 0.012465f
C603 B.n563 VSUBS 0.012465f
C604 B.n564 VSUBS 0.012465f
C605 B.n565 VSUBS 0.012465f
C606 B.n566 VSUBS 0.012465f
C607 B.n567 VSUBS 0.012465f
C608 B.n568 VSUBS 0.012465f
C609 B.n569 VSUBS 0.012465f
C610 B.n570 VSUBS 0.012465f
C611 B.n571 VSUBS 0.012465f
C612 B.n572 VSUBS 0.012465f
C613 B.n573 VSUBS 0.012465f
C614 B.n574 VSUBS 0.012465f
C615 B.n575 VSUBS 0.012465f
C616 B.n576 VSUBS 0.012465f
C617 B.n577 VSUBS 0.029503f
C618 B.n578 VSUBS 0.031357f
C619 B.n579 VSUBS 0.029975f
C620 B.n580 VSUBS 0.012465f
C621 B.n581 VSUBS 0.012465f
C622 B.n582 VSUBS 0.012465f
C623 B.n583 VSUBS 0.012465f
C624 B.n584 VSUBS 0.012465f
C625 B.n585 VSUBS 0.012465f
C626 B.n586 VSUBS 0.012465f
C627 B.n587 VSUBS 0.012465f
C628 B.n588 VSUBS 0.012465f
C629 B.n589 VSUBS 0.012465f
C630 B.n590 VSUBS 0.012465f
C631 B.n591 VSUBS 0.012465f
C632 B.n592 VSUBS 0.012465f
C633 B.n593 VSUBS 0.012465f
C634 B.n594 VSUBS 0.012465f
C635 B.n595 VSUBS 0.012465f
C636 B.n596 VSUBS 0.012465f
C637 B.n597 VSUBS 0.012465f
C638 B.n598 VSUBS 0.012465f
C639 B.n599 VSUBS 0.012465f
C640 B.n600 VSUBS 0.012465f
C641 B.n601 VSUBS 0.012465f
C642 B.n602 VSUBS 0.012465f
C643 B.n603 VSUBS 0.012465f
C644 B.n604 VSUBS 0.012465f
C645 B.n605 VSUBS 0.012465f
C646 B.n606 VSUBS 0.012465f
C647 B.n607 VSUBS 0.012465f
C648 B.n608 VSUBS 0.012465f
C649 B.n609 VSUBS 0.011732f
C650 B.n610 VSUBS 0.028881f
C651 B.n611 VSUBS 0.006966f
C652 B.n612 VSUBS 0.012465f
C653 B.n613 VSUBS 0.012465f
C654 B.n614 VSUBS 0.012465f
C655 B.n615 VSUBS 0.012465f
C656 B.n616 VSUBS 0.012465f
C657 B.n617 VSUBS 0.012465f
C658 B.n618 VSUBS 0.012465f
C659 B.n619 VSUBS 0.012465f
C660 B.n620 VSUBS 0.012465f
C661 B.n621 VSUBS 0.012465f
C662 B.n622 VSUBS 0.012465f
C663 B.n623 VSUBS 0.012465f
C664 B.n624 VSUBS 0.006966f
C665 B.n625 VSUBS 0.012465f
C666 B.n626 VSUBS 0.012465f
C667 B.n627 VSUBS 0.011732f
C668 B.n628 VSUBS 0.012465f
C669 B.n629 VSUBS 0.012465f
C670 B.n630 VSUBS 0.012465f
C671 B.n631 VSUBS 0.012465f
C672 B.n632 VSUBS 0.012465f
C673 B.n633 VSUBS 0.012465f
C674 B.n634 VSUBS 0.012465f
C675 B.n635 VSUBS 0.012465f
C676 B.n636 VSUBS 0.012465f
C677 B.n637 VSUBS 0.012465f
C678 B.n638 VSUBS 0.012465f
C679 B.n639 VSUBS 0.012465f
C680 B.n640 VSUBS 0.012465f
C681 B.n641 VSUBS 0.012465f
C682 B.n642 VSUBS 0.012465f
C683 B.n643 VSUBS 0.012465f
C684 B.n644 VSUBS 0.012465f
C685 B.n645 VSUBS 0.012465f
C686 B.n646 VSUBS 0.012465f
C687 B.n647 VSUBS 0.012465f
C688 B.n648 VSUBS 0.012465f
C689 B.n649 VSUBS 0.012465f
C690 B.n650 VSUBS 0.012465f
C691 B.n651 VSUBS 0.012465f
C692 B.n652 VSUBS 0.012465f
C693 B.n653 VSUBS 0.012465f
C694 B.n654 VSUBS 0.012465f
C695 B.n655 VSUBS 0.012465f
C696 B.n656 VSUBS 0.031357f
C697 B.n657 VSUBS 0.031357f
C698 B.n658 VSUBS 0.029503f
C699 B.n659 VSUBS 0.012465f
C700 B.n660 VSUBS 0.012465f
C701 B.n661 VSUBS 0.012465f
C702 B.n662 VSUBS 0.012465f
C703 B.n663 VSUBS 0.012465f
C704 B.n664 VSUBS 0.012465f
C705 B.n665 VSUBS 0.012465f
C706 B.n666 VSUBS 0.012465f
C707 B.n667 VSUBS 0.012465f
C708 B.n668 VSUBS 0.012465f
C709 B.n669 VSUBS 0.012465f
C710 B.n670 VSUBS 0.012465f
C711 B.n671 VSUBS 0.012465f
C712 B.n672 VSUBS 0.012465f
C713 B.n673 VSUBS 0.012465f
C714 B.n674 VSUBS 0.012465f
C715 B.n675 VSUBS 0.012465f
C716 B.n676 VSUBS 0.012465f
C717 B.n677 VSUBS 0.012465f
C718 B.n678 VSUBS 0.012465f
C719 B.n679 VSUBS 0.012465f
C720 B.n680 VSUBS 0.012465f
C721 B.n681 VSUBS 0.012465f
C722 B.n682 VSUBS 0.012465f
C723 B.n683 VSUBS 0.012465f
C724 B.n684 VSUBS 0.012465f
C725 B.n685 VSUBS 0.012465f
C726 B.n686 VSUBS 0.012465f
C727 B.n687 VSUBS 0.012465f
C728 B.n688 VSUBS 0.012465f
C729 B.n689 VSUBS 0.012465f
C730 B.n690 VSUBS 0.012465f
C731 B.n691 VSUBS 0.012465f
C732 B.n692 VSUBS 0.012465f
C733 B.n693 VSUBS 0.012465f
C734 B.n694 VSUBS 0.012465f
C735 B.n695 VSUBS 0.012465f
C736 B.n696 VSUBS 0.012465f
C737 B.n697 VSUBS 0.012465f
C738 B.n698 VSUBS 0.012465f
C739 B.n699 VSUBS 0.012465f
C740 B.n700 VSUBS 0.012465f
C741 B.n701 VSUBS 0.012465f
C742 B.n702 VSUBS 0.012465f
C743 B.n703 VSUBS 0.012465f
C744 B.n704 VSUBS 0.012465f
C745 B.n705 VSUBS 0.012465f
C746 B.n706 VSUBS 0.012465f
C747 B.n707 VSUBS 0.012465f
C748 B.n708 VSUBS 0.012465f
C749 B.n709 VSUBS 0.012465f
C750 B.n710 VSUBS 0.012465f
C751 B.n711 VSUBS 0.012465f
C752 B.n712 VSUBS 0.012465f
C753 B.n713 VSUBS 0.012465f
C754 B.n714 VSUBS 0.012465f
C755 B.n715 VSUBS 0.012465f
C756 B.n716 VSUBS 0.012465f
C757 B.n717 VSUBS 0.012465f
C758 B.n718 VSUBS 0.012465f
C759 B.n719 VSUBS 0.012465f
C760 B.n720 VSUBS 0.012465f
C761 B.n721 VSUBS 0.012465f
C762 B.n722 VSUBS 0.012465f
C763 B.n723 VSUBS 0.012465f
C764 B.n724 VSUBS 0.012465f
C765 B.n725 VSUBS 0.012465f
C766 B.n726 VSUBS 0.012465f
C767 B.n727 VSUBS 0.012465f
C768 B.n728 VSUBS 0.012465f
C769 B.n729 VSUBS 0.012465f
C770 B.n730 VSUBS 0.012465f
C771 B.n731 VSUBS 0.012465f
C772 B.n732 VSUBS 0.012465f
C773 B.n733 VSUBS 0.012465f
C774 B.n734 VSUBS 0.012465f
C775 B.n735 VSUBS 0.012465f
C776 B.n736 VSUBS 0.012465f
C777 B.n737 VSUBS 0.012465f
C778 B.n738 VSUBS 0.012465f
C779 B.n739 VSUBS 0.012465f
C780 B.n740 VSUBS 0.012465f
C781 B.n741 VSUBS 0.012465f
C782 B.n742 VSUBS 0.012465f
C783 B.n743 VSUBS 0.012465f
C784 B.n744 VSUBS 0.012465f
C785 B.n745 VSUBS 0.012465f
C786 B.n746 VSUBS 0.012465f
C787 B.n747 VSUBS 0.012465f
C788 B.n748 VSUBS 0.012465f
C789 B.n749 VSUBS 0.012465f
C790 B.n750 VSUBS 0.012465f
C791 B.n751 VSUBS 0.012465f
C792 B.n752 VSUBS 0.012465f
C793 B.n753 VSUBS 0.012465f
C794 B.n754 VSUBS 0.012465f
C795 B.n755 VSUBS 0.012465f
C796 B.n756 VSUBS 0.012465f
C797 B.n757 VSUBS 0.012465f
C798 B.n758 VSUBS 0.012465f
C799 B.n759 VSUBS 0.028226f
C800 VDD2.t2 VSUBS 1.24015f
C801 VDD2.t0 VSUBS 0.141728f
C802 VDD2.t7 VSUBS 0.141728f
C803 VDD2.n0 VSUBS 0.896013f
C804 VDD2.n1 VSUBS 1.87917f
C805 VDD2.t4 VSUBS 0.141728f
C806 VDD2.t6 VSUBS 0.141728f
C807 VDD2.n2 VSUBS 0.918636f
C808 VDD2.n3 VSUBS 4.08639f
C809 VDD2.t1 VSUBS 1.21567f
C810 VDD2.n4 VSUBS 4.11904f
C811 VDD2.t9 VSUBS 0.141728f
C812 VDD2.t3 VSUBS 0.141728f
C813 VDD2.n5 VSUBS 0.896017f
C814 VDD2.n6 VSUBS 0.961669f
C815 VDD2.t8 VSUBS 0.141728f
C816 VDD2.t5 VSUBS 0.141728f
C817 VDD2.n7 VSUBS 0.918591f
C818 VN.t3 VSUBS 1.42479f
C819 VN.n0 VSUBS 0.686772f
C820 VN.n1 VSUBS 0.035616f
C821 VN.n2 VSUBS 0.054237f
C822 VN.n3 VSUBS 0.035616f
C823 VN.t5 VSUBS 1.42479f
C824 VN.n4 VSUBS 0.066047f
C825 VN.n5 VSUBS 0.035616f
C826 VN.n6 VSUBS 0.066047f
C827 VN.n7 VSUBS 0.035616f
C828 VN.t2 VSUBS 1.42479f
C829 VN.n8 VSUBS 0.066681f
C830 VN.n9 VSUBS 0.035616f
C831 VN.n10 VSUBS 0.039963f
C832 VN.t9 VSUBS 1.42479f
C833 VN.n11 VSUBS 0.644788f
C834 VN.t7 VSUBS 1.76957f
C835 VN.n12 VSUBS 0.627457f
C836 VN.n13 VSUBS 0.384551f
C837 VN.n14 VSUBS 0.035616f
C838 VN.n15 VSUBS 0.066047f
C839 VN.n16 VSUBS 0.071509f
C840 VN.n17 VSUBS 0.031405f
C841 VN.n18 VSUBS 0.035616f
C842 VN.n19 VSUBS 0.035616f
C843 VN.n20 VSUBS 0.035616f
C844 VN.n21 VSUBS 0.066047f
C845 VN.n22 VSUBS 0.049744f
C846 VN.n23 VSUBS 0.541028f
C847 VN.n24 VSUBS 0.049744f
C848 VN.n25 VSUBS 0.035616f
C849 VN.n26 VSUBS 0.035616f
C850 VN.n27 VSUBS 0.035616f
C851 VN.n28 VSUBS 0.066681f
C852 VN.n29 VSUBS 0.031405f
C853 VN.n30 VSUBS 0.071509f
C854 VN.n31 VSUBS 0.035616f
C855 VN.n32 VSUBS 0.035616f
C856 VN.n33 VSUBS 0.035616f
C857 VN.n34 VSUBS 0.039963f
C858 VN.n35 VSUBS 0.541028f
C859 VN.n36 VSUBS 0.059526f
C860 VN.n37 VSUBS 0.066047f
C861 VN.n38 VSUBS 0.035616f
C862 VN.n39 VSUBS 0.035616f
C863 VN.n40 VSUBS 0.035616f
C864 VN.n41 VSUBS 0.04931f
C865 VN.n42 VSUBS 0.066047f
C866 VN.n43 VSUBS 0.062786f
C867 VN.n44 VSUBS 0.057475f
C868 VN.n45 VSUBS 0.070876f
C869 VN.t8 VSUBS 1.42479f
C870 VN.n46 VSUBS 0.686772f
C871 VN.n47 VSUBS 0.035616f
C872 VN.n48 VSUBS 0.054237f
C873 VN.n49 VSUBS 0.035616f
C874 VN.t0 VSUBS 1.42479f
C875 VN.n50 VSUBS 0.066047f
C876 VN.n51 VSUBS 0.035616f
C877 VN.n52 VSUBS 0.066047f
C878 VN.n53 VSUBS 0.035616f
C879 VN.t6 VSUBS 1.42479f
C880 VN.n54 VSUBS 0.066681f
C881 VN.n55 VSUBS 0.035616f
C882 VN.n56 VSUBS 0.039963f
C883 VN.t4 VSUBS 1.76957f
C884 VN.t1 VSUBS 1.42479f
C885 VN.n57 VSUBS 0.644788f
C886 VN.n58 VSUBS 0.627457f
C887 VN.n59 VSUBS 0.384551f
C888 VN.n60 VSUBS 0.035616f
C889 VN.n61 VSUBS 0.066047f
C890 VN.n62 VSUBS 0.071509f
C891 VN.n63 VSUBS 0.031405f
C892 VN.n64 VSUBS 0.035616f
C893 VN.n65 VSUBS 0.035616f
C894 VN.n66 VSUBS 0.035616f
C895 VN.n67 VSUBS 0.066047f
C896 VN.n68 VSUBS 0.049744f
C897 VN.n69 VSUBS 0.541028f
C898 VN.n70 VSUBS 0.049744f
C899 VN.n71 VSUBS 0.035616f
C900 VN.n72 VSUBS 0.035616f
C901 VN.n73 VSUBS 0.035616f
C902 VN.n74 VSUBS 0.066681f
C903 VN.n75 VSUBS 0.031405f
C904 VN.n76 VSUBS 0.071509f
C905 VN.n77 VSUBS 0.035616f
C906 VN.n78 VSUBS 0.035616f
C907 VN.n79 VSUBS 0.035616f
C908 VN.n80 VSUBS 0.039963f
C909 VN.n81 VSUBS 0.541028f
C910 VN.n82 VSUBS 0.059526f
C911 VN.n83 VSUBS 0.066047f
C912 VN.n84 VSUBS 0.035616f
C913 VN.n85 VSUBS 0.035616f
C914 VN.n86 VSUBS 0.035616f
C915 VN.n87 VSUBS 0.04931f
C916 VN.n88 VSUBS 0.066047f
C917 VN.n89 VSUBS 0.062786f
C918 VN.n90 VSUBS 0.057475f
C919 VN.n91 VSUBS 2.04307f
C920 VDD1.t5 VSUBS 1.25073f
C921 VDD1.t0 VSUBS 0.142936f
C922 VDD1.t9 VSUBS 0.142936f
C923 VDD1.n0 VSUBS 0.903657f
C924 VDD1.n1 VSUBS 1.90702f
C925 VDD1.t1 VSUBS 1.25073f
C926 VDD1.t3 VSUBS 0.142936f
C927 VDD1.t2 VSUBS 0.142936f
C928 VDD1.n2 VSUBS 0.903653f
C929 VDD1.n3 VSUBS 1.89519f
C930 VDD1.t6 VSUBS 0.142936f
C931 VDD1.t8 VSUBS 0.142936f
C932 VDD1.n4 VSUBS 0.926468f
C933 VDD1.n5 VSUBS 4.30757f
C934 VDD1.t4 VSUBS 0.142936f
C935 VDD1.t7 VSUBS 0.142936f
C936 VDD1.n6 VSUBS 0.903652f
C937 VDD1.n7 VSUBS 4.27519f
C938 VTAIL.t2 VSUBS 0.141075f
C939 VTAIL.t1 VSUBS 0.141075f
C940 VTAIL.n0 VSUBS 0.788986f
C941 VTAIL.n1 VSUBS 1.0656f
C942 VTAIL.t10 VSUBS 1.10233f
C943 VTAIL.n2 VSUBS 1.21247f
C944 VTAIL.t9 VSUBS 0.141075f
C945 VTAIL.t12 VSUBS 0.141075f
C946 VTAIL.n3 VSUBS 0.788986f
C947 VTAIL.n4 VSUBS 1.25181f
C948 VTAIL.t14 VSUBS 0.141075f
C949 VTAIL.t11 VSUBS 0.141075f
C950 VTAIL.n5 VSUBS 0.788986f
C951 VTAIL.n6 VSUBS 2.55528f
C952 VTAIL.t0 VSUBS 0.141075f
C953 VTAIL.t4 VSUBS 0.141075f
C954 VTAIL.n7 VSUBS 0.788991f
C955 VTAIL.n8 VSUBS 2.55527f
C956 VTAIL.t16 VSUBS 0.141075f
C957 VTAIL.t3 VSUBS 0.141075f
C958 VTAIL.n9 VSUBS 0.788991f
C959 VTAIL.n10 VSUBS 1.2518f
C960 VTAIL.t19 VSUBS 1.10233f
C961 VTAIL.n11 VSUBS 1.21247f
C962 VTAIL.t6 VSUBS 0.141075f
C963 VTAIL.t8 VSUBS 0.141075f
C964 VTAIL.n12 VSUBS 0.788991f
C965 VTAIL.n13 VSUBS 1.14106f
C966 VTAIL.t13 VSUBS 0.141075f
C967 VTAIL.t7 VSUBS 0.141075f
C968 VTAIL.n14 VSUBS 0.788991f
C969 VTAIL.n15 VSUBS 1.2518f
C970 VTAIL.t15 VSUBS 1.10233f
C971 VTAIL.n16 VSUBS 2.29837f
C972 VTAIL.t18 VSUBS 1.10233f
C973 VTAIL.n17 VSUBS 2.29837f
C974 VTAIL.t17 VSUBS 0.141075f
C975 VTAIL.t5 VSUBS 0.141075f
C976 VTAIL.n18 VSUBS 0.788986f
C977 VTAIL.n19 VSUBS 0.998959f
C978 VP.t1 VSUBS 1.60078f
C979 VP.n0 VSUBS 0.771603f
C980 VP.n1 VSUBS 0.040016f
C981 VP.n2 VSUBS 0.060937f
C982 VP.n3 VSUBS 0.040016f
C983 VP.t3 VSUBS 1.60078f
C984 VP.n4 VSUBS 0.074205f
C985 VP.n5 VSUBS 0.040016f
C986 VP.n6 VSUBS 0.074205f
C987 VP.n7 VSUBS 0.040016f
C988 VP.t7 VSUBS 1.60078f
C989 VP.n8 VSUBS 0.074917f
C990 VP.n9 VSUBS 0.040016f
C991 VP.n10 VSUBS 0.044899f
C992 VP.n11 VSUBS 0.040016f
C993 VP.n12 VSUBS 0.055401f
C994 VP.n13 VSUBS 0.064574f
C995 VP.t8 VSUBS 1.60078f
C996 VP.t2 VSUBS 1.60078f
C997 VP.n14 VSUBS 0.771603f
C998 VP.n15 VSUBS 0.040016f
C999 VP.n16 VSUBS 0.060937f
C1000 VP.n17 VSUBS 0.040016f
C1001 VP.t5 VSUBS 1.60078f
C1002 VP.n18 VSUBS 0.074205f
C1003 VP.n19 VSUBS 0.040016f
C1004 VP.n20 VSUBS 0.074205f
C1005 VP.n21 VSUBS 0.040016f
C1006 VP.t0 VSUBS 1.60078f
C1007 VP.n22 VSUBS 0.074917f
C1008 VP.n23 VSUBS 0.040016f
C1009 VP.n24 VSUBS 0.044899f
C1010 VP.t4 VSUBS 1.98815f
C1011 VP.t9 VSUBS 1.60078f
C1012 VP.n25 VSUBS 0.724433f
C1013 VP.n26 VSUBS 0.704963f
C1014 VP.n27 VSUBS 0.432053f
C1015 VP.n28 VSUBS 0.040016f
C1016 VP.n29 VSUBS 0.074205f
C1017 VP.n30 VSUBS 0.080342f
C1018 VP.n31 VSUBS 0.035284f
C1019 VP.n32 VSUBS 0.040016f
C1020 VP.n33 VSUBS 0.040016f
C1021 VP.n34 VSUBS 0.040016f
C1022 VP.n35 VSUBS 0.074205f
C1023 VP.n36 VSUBS 0.055889f
C1024 VP.n37 VSUBS 0.607857f
C1025 VP.n38 VSUBS 0.055889f
C1026 VP.n39 VSUBS 0.040016f
C1027 VP.n40 VSUBS 0.040016f
C1028 VP.n41 VSUBS 0.040016f
C1029 VP.n42 VSUBS 0.074917f
C1030 VP.n43 VSUBS 0.035284f
C1031 VP.n44 VSUBS 0.080342f
C1032 VP.n45 VSUBS 0.040016f
C1033 VP.n46 VSUBS 0.040016f
C1034 VP.n47 VSUBS 0.040016f
C1035 VP.n48 VSUBS 0.044899f
C1036 VP.n49 VSUBS 0.607857f
C1037 VP.n50 VSUBS 0.066879f
C1038 VP.n51 VSUBS 0.074205f
C1039 VP.n52 VSUBS 0.040016f
C1040 VP.n53 VSUBS 0.040016f
C1041 VP.n54 VSUBS 0.040016f
C1042 VP.n55 VSUBS 0.055401f
C1043 VP.n56 VSUBS 0.074205f
C1044 VP.n57 VSUBS 0.070542f
C1045 VP.n58 VSUBS 0.064574f
C1046 VP.n59 VSUBS 2.27911f
C1047 VP.n60 VSUBS 2.30779f
C1048 VP.n61 VSUBS 0.771603f
C1049 VP.n62 VSUBS 0.070542f
C1050 VP.n63 VSUBS 0.074205f
C1051 VP.n64 VSUBS 0.040016f
C1052 VP.n65 VSUBS 0.040016f
C1053 VP.n66 VSUBS 0.040016f
C1054 VP.n67 VSUBS 0.060937f
C1055 VP.n68 VSUBS 0.074205f
C1056 VP.t6 VSUBS 1.60078f
C1057 VP.n69 VSUBS 0.607857f
C1058 VP.n70 VSUBS 0.066879f
C1059 VP.n71 VSUBS 0.040016f
C1060 VP.n72 VSUBS 0.040016f
C1061 VP.n73 VSUBS 0.040016f
C1062 VP.n74 VSUBS 0.074205f
C1063 VP.n75 VSUBS 0.080342f
C1064 VP.n76 VSUBS 0.035284f
C1065 VP.n77 VSUBS 0.040016f
C1066 VP.n78 VSUBS 0.040016f
C1067 VP.n79 VSUBS 0.040016f
C1068 VP.n80 VSUBS 0.074205f
C1069 VP.n81 VSUBS 0.055889f
C1070 VP.n82 VSUBS 0.607857f
C1071 VP.n83 VSUBS 0.055889f
C1072 VP.n84 VSUBS 0.040016f
C1073 VP.n85 VSUBS 0.040016f
C1074 VP.n86 VSUBS 0.040016f
C1075 VP.n87 VSUBS 0.074917f
C1076 VP.n88 VSUBS 0.035284f
C1077 VP.n89 VSUBS 0.080342f
C1078 VP.n90 VSUBS 0.040016f
C1079 VP.n91 VSUBS 0.040016f
C1080 VP.n92 VSUBS 0.040016f
C1081 VP.n93 VSUBS 0.044899f
C1082 VP.n94 VSUBS 0.607857f
C1083 VP.n95 VSUBS 0.066879f
C1084 VP.n96 VSUBS 0.074205f
C1085 VP.n97 VSUBS 0.040016f
C1086 VP.n98 VSUBS 0.040016f
C1087 VP.n99 VSUBS 0.040016f
C1088 VP.n100 VSUBS 0.055401f
C1089 VP.n101 VSUBS 0.074205f
C1090 VP.n102 VSUBS 0.070542f
C1091 VP.n103 VSUBS 0.064574f
C1092 VP.n104 VSUBS 0.07963f
.ends

