* NGSPICE file created from diff_pair_sample_1341.ext - technology: sky130A

.subckt diff_pair_sample_1341 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t5 VP.t0 VTAIL.t11 B.t2 sky130_fd_pr__nfet_01v8 ad=1.551 pd=9.73 as=3.666 ps=19.58 w=9.4 l=3.86
X1 B.t19 B.t17 B.t18 B.t14 sky130_fd_pr__nfet_01v8 ad=3.666 pd=19.58 as=0 ps=0 w=9.4 l=3.86
X2 VDD1.t4 VP.t1 VTAIL.t9 B.t5 sky130_fd_pr__nfet_01v8 ad=3.666 pd=19.58 as=1.551 ps=9.73 w=9.4 l=3.86
X3 VDD1.t3 VP.t2 VTAIL.t10 B.t4 sky130_fd_pr__nfet_01v8 ad=3.666 pd=19.58 as=1.551 ps=9.73 w=9.4 l=3.86
X4 VTAIL.t6 VP.t3 VDD1.t2 B.t0 sky130_fd_pr__nfet_01v8 ad=1.551 pd=9.73 as=1.551 ps=9.73 w=9.4 l=3.86
X5 VDD1.t1 VP.t4 VTAIL.t8 B.t1 sky130_fd_pr__nfet_01v8 ad=1.551 pd=9.73 as=3.666 ps=19.58 w=9.4 l=3.86
X6 VDD2.t5 VN.t0 VTAIL.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=3.666 pd=19.58 as=1.551 ps=9.73 w=9.4 l=3.86
X7 VTAIL.t0 VN.t1 VDD2.t4 B.t0 sky130_fd_pr__nfet_01v8 ad=1.551 pd=9.73 as=1.551 ps=9.73 w=9.4 l=3.86
X8 VDD2.t3 VN.t2 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=1.551 pd=9.73 as=3.666 ps=19.58 w=9.4 l=3.86
X9 VDD2.t2 VN.t3 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=1.551 pd=9.73 as=3.666 ps=19.58 w=9.4 l=3.86
X10 B.t16 B.t13 B.t15 B.t14 sky130_fd_pr__nfet_01v8 ad=3.666 pd=19.58 as=0 ps=0 w=9.4 l=3.86
X11 VDD2.t1 VN.t4 VTAIL.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=3.666 pd=19.58 as=1.551 ps=9.73 w=9.4 l=3.86
X12 VTAIL.t3 VN.t5 VDD2.t0 B.t3 sky130_fd_pr__nfet_01v8 ad=1.551 pd=9.73 as=1.551 ps=9.73 w=9.4 l=3.86
X13 VTAIL.t7 VP.t5 VDD1.t0 B.t3 sky130_fd_pr__nfet_01v8 ad=1.551 pd=9.73 as=1.551 ps=9.73 w=9.4 l=3.86
X14 B.t12 B.t10 B.t11 B.t7 sky130_fd_pr__nfet_01v8 ad=3.666 pd=19.58 as=0 ps=0 w=9.4 l=3.86
X15 B.t9 B.t6 B.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=3.666 pd=19.58 as=0 ps=0 w=9.4 l=3.86
R0 VP.n15 VP.n14 161.3
R1 VP.n16 VP.n11 161.3
R2 VP.n18 VP.n17 161.3
R3 VP.n19 VP.n10 161.3
R4 VP.n21 VP.n20 161.3
R5 VP.n22 VP.n9 161.3
R6 VP.n24 VP.n23 161.3
R7 VP.n25 VP.n8 161.3
R8 VP.n54 VP.n0 161.3
R9 VP.n53 VP.n52 161.3
R10 VP.n51 VP.n1 161.3
R11 VP.n50 VP.n49 161.3
R12 VP.n48 VP.n2 161.3
R13 VP.n47 VP.n46 161.3
R14 VP.n45 VP.n3 161.3
R15 VP.n44 VP.n43 161.3
R16 VP.n41 VP.n4 161.3
R17 VP.n40 VP.n39 161.3
R18 VP.n38 VP.n5 161.3
R19 VP.n37 VP.n36 161.3
R20 VP.n35 VP.n6 161.3
R21 VP.n34 VP.n33 161.3
R22 VP.n32 VP.n7 161.3
R23 VP.n31 VP.n30 161.3
R24 VP.n12 VP.t1 90.8175
R25 VP.n13 VP.n12 62.6969
R26 VP.n29 VP.n28 60.5633
R27 VP.n56 VP.n55 60.5633
R28 VP.n27 VP.n26 60.5633
R29 VP.n29 VP.t2 58.6896
R30 VP.n42 VP.t5 58.6896
R31 VP.n55 VP.t0 58.6896
R32 VP.n26 VP.t4 58.6896
R33 VP.n13 VP.t3 58.6896
R34 VP.n36 VP.n35 55.5035
R35 VP.n49 VP.n48 55.5035
R36 VP.n20 VP.n19 55.5035
R37 VP.n28 VP.n27 51.8785
R38 VP.n35 VP.n34 25.3177
R39 VP.n49 VP.n1 25.3177
R40 VP.n20 VP.n9 25.3177
R41 VP.n30 VP.n7 24.3439
R42 VP.n34 VP.n7 24.3439
R43 VP.n36 VP.n5 24.3439
R44 VP.n40 VP.n5 24.3439
R45 VP.n41 VP.n40 24.3439
R46 VP.n43 VP.n3 24.3439
R47 VP.n47 VP.n3 24.3439
R48 VP.n48 VP.n47 24.3439
R49 VP.n53 VP.n1 24.3439
R50 VP.n54 VP.n53 24.3439
R51 VP.n24 VP.n9 24.3439
R52 VP.n25 VP.n24 24.3439
R53 VP.n14 VP.n11 24.3439
R54 VP.n18 VP.n11 24.3439
R55 VP.n19 VP.n18 24.3439
R56 VP.n30 VP.n29 21.4227
R57 VP.n55 VP.n54 21.4227
R58 VP.n26 VP.n25 21.4227
R59 VP.n42 VP.n41 12.1722
R60 VP.n43 VP.n42 12.1722
R61 VP.n14 VP.n13 12.1722
R62 VP.n15 VP.n12 2.65071
R63 VP.n27 VP.n8 0.417764
R64 VP.n31 VP.n28 0.417764
R65 VP.n56 VP.n0 0.417764
R66 VP VP.n56 0.394061
R67 VP.n16 VP.n15 0.189894
R68 VP.n17 VP.n16 0.189894
R69 VP.n17 VP.n10 0.189894
R70 VP.n21 VP.n10 0.189894
R71 VP.n22 VP.n21 0.189894
R72 VP.n23 VP.n22 0.189894
R73 VP.n23 VP.n8 0.189894
R74 VP.n32 VP.n31 0.189894
R75 VP.n33 VP.n32 0.189894
R76 VP.n33 VP.n6 0.189894
R77 VP.n37 VP.n6 0.189894
R78 VP.n38 VP.n37 0.189894
R79 VP.n39 VP.n38 0.189894
R80 VP.n39 VP.n4 0.189894
R81 VP.n44 VP.n4 0.189894
R82 VP.n45 VP.n44 0.189894
R83 VP.n46 VP.n45 0.189894
R84 VP.n46 VP.n2 0.189894
R85 VP.n50 VP.n2 0.189894
R86 VP.n51 VP.n50 0.189894
R87 VP.n52 VP.n51 0.189894
R88 VP.n52 VP.n0 0.189894
R89 VTAIL.n202 VTAIL.n158 289.615
R90 VTAIL.n46 VTAIL.n2 289.615
R91 VTAIL.n152 VTAIL.n108 289.615
R92 VTAIL.n100 VTAIL.n56 289.615
R93 VTAIL.n175 VTAIL.n174 185
R94 VTAIL.n177 VTAIL.n176 185
R95 VTAIL.n170 VTAIL.n169 185
R96 VTAIL.n183 VTAIL.n182 185
R97 VTAIL.n185 VTAIL.n184 185
R98 VTAIL.n166 VTAIL.n165 185
R99 VTAIL.n192 VTAIL.n191 185
R100 VTAIL.n193 VTAIL.n164 185
R101 VTAIL.n195 VTAIL.n194 185
R102 VTAIL.n162 VTAIL.n161 185
R103 VTAIL.n201 VTAIL.n200 185
R104 VTAIL.n203 VTAIL.n202 185
R105 VTAIL.n19 VTAIL.n18 185
R106 VTAIL.n21 VTAIL.n20 185
R107 VTAIL.n14 VTAIL.n13 185
R108 VTAIL.n27 VTAIL.n26 185
R109 VTAIL.n29 VTAIL.n28 185
R110 VTAIL.n10 VTAIL.n9 185
R111 VTAIL.n36 VTAIL.n35 185
R112 VTAIL.n37 VTAIL.n8 185
R113 VTAIL.n39 VTAIL.n38 185
R114 VTAIL.n6 VTAIL.n5 185
R115 VTAIL.n45 VTAIL.n44 185
R116 VTAIL.n47 VTAIL.n46 185
R117 VTAIL.n153 VTAIL.n152 185
R118 VTAIL.n151 VTAIL.n150 185
R119 VTAIL.n112 VTAIL.n111 185
R120 VTAIL.n116 VTAIL.n114 185
R121 VTAIL.n145 VTAIL.n144 185
R122 VTAIL.n143 VTAIL.n142 185
R123 VTAIL.n118 VTAIL.n117 185
R124 VTAIL.n137 VTAIL.n136 185
R125 VTAIL.n135 VTAIL.n134 185
R126 VTAIL.n122 VTAIL.n121 185
R127 VTAIL.n129 VTAIL.n128 185
R128 VTAIL.n127 VTAIL.n126 185
R129 VTAIL.n101 VTAIL.n100 185
R130 VTAIL.n99 VTAIL.n98 185
R131 VTAIL.n60 VTAIL.n59 185
R132 VTAIL.n64 VTAIL.n62 185
R133 VTAIL.n93 VTAIL.n92 185
R134 VTAIL.n91 VTAIL.n90 185
R135 VTAIL.n66 VTAIL.n65 185
R136 VTAIL.n85 VTAIL.n84 185
R137 VTAIL.n83 VTAIL.n82 185
R138 VTAIL.n70 VTAIL.n69 185
R139 VTAIL.n77 VTAIL.n76 185
R140 VTAIL.n75 VTAIL.n74 185
R141 VTAIL.n173 VTAIL.t1 149.524
R142 VTAIL.n17 VTAIL.t11 149.524
R143 VTAIL.n125 VTAIL.t8 149.524
R144 VTAIL.n73 VTAIL.t2 149.524
R145 VTAIL.n176 VTAIL.n175 104.615
R146 VTAIL.n176 VTAIL.n169 104.615
R147 VTAIL.n183 VTAIL.n169 104.615
R148 VTAIL.n184 VTAIL.n183 104.615
R149 VTAIL.n184 VTAIL.n165 104.615
R150 VTAIL.n192 VTAIL.n165 104.615
R151 VTAIL.n193 VTAIL.n192 104.615
R152 VTAIL.n194 VTAIL.n193 104.615
R153 VTAIL.n194 VTAIL.n161 104.615
R154 VTAIL.n201 VTAIL.n161 104.615
R155 VTAIL.n202 VTAIL.n201 104.615
R156 VTAIL.n20 VTAIL.n19 104.615
R157 VTAIL.n20 VTAIL.n13 104.615
R158 VTAIL.n27 VTAIL.n13 104.615
R159 VTAIL.n28 VTAIL.n27 104.615
R160 VTAIL.n28 VTAIL.n9 104.615
R161 VTAIL.n36 VTAIL.n9 104.615
R162 VTAIL.n37 VTAIL.n36 104.615
R163 VTAIL.n38 VTAIL.n37 104.615
R164 VTAIL.n38 VTAIL.n5 104.615
R165 VTAIL.n45 VTAIL.n5 104.615
R166 VTAIL.n46 VTAIL.n45 104.615
R167 VTAIL.n152 VTAIL.n151 104.615
R168 VTAIL.n151 VTAIL.n111 104.615
R169 VTAIL.n116 VTAIL.n111 104.615
R170 VTAIL.n144 VTAIL.n116 104.615
R171 VTAIL.n144 VTAIL.n143 104.615
R172 VTAIL.n143 VTAIL.n117 104.615
R173 VTAIL.n136 VTAIL.n117 104.615
R174 VTAIL.n136 VTAIL.n135 104.615
R175 VTAIL.n135 VTAIL.n121 104.615
R176 VTAIL.n128 VTAIL.n121 104.615
R177 VTAIL.n128 VTAIL.n127 104.615
R178 VTAIL.n100 VTAIL.n99 104.615
R179 VTAIL.n99 VTAIL.n59 104.615
R180 VTAIL.n64 VTAIL.n59 104.615
R181 VTAIL.n92 VTAIL.n64 104.615
R182 VTAIL.n92 VTAIL.n91 104.615
R183 VTAIL.n91 VTAIL.n65 104.615
R184 VTAIL.n84 VTAIL.n65 104.615
R185 VTAIL.n84 VTAIL.n83 104.615
R186 VTAIL.n83 VTAIL.n69 104.615
R187 VTAIL.n76 VTAIL.n69 104.615
R188 VTAIL.n76 VTAIL.n75 104.615
R189 VTAIL.n175 VTAIL.t1 52.3082
R190 VTAIL.n19 VTAIL.t11 52.3082
R191 VTAIL.n127 VTAIL.t8 52.3082
R192 VTAIL.n75 VTAIL.t2 52.3082
R193 VTAIL.n107 VTAIL.n106 49.4263
R194 VTAIL.n55 VTAIL.n54 49.4263
R195 VTAIL.n1 VTAIL.n0 49.4261
R196 VTAIL.n53 VTAIL.n52 49.4261
R197 VTAIL.n207 VTAIL.n206 35.2884
R198 VTAIL.n51 VTAIL.n50 35.2884
R199 VTAIL.n157 VTAIL.n156 35.2884
R200 VTAIL.n105 VTAIL.n104 35.2884
R201 VTAIL.n55 VTAIL.n53 27.6945
R202 VTAIL.n207 VTAIL.n157 24.0824
R203 VTAIL.n195 VTAIL.n162 13.1884
R204 VTAIL.n39 VTAIL.n6 13.1884
R205 VTAIL.n114 VTAIL.n112 13.1884
R206 VTAIL.n62 VTAIL.n60 13.1884
R207 VTAIL.n196 VTAIL.n164 12.8005
R208 VTAIL.n200 VTAIL.n199 12.8005
R209 VTAIL.n40 VTAIL.n8 12.8005
R210 VTAIL.n44 VTAIL.n43 12.8005
R211 VTAIL.n150 VTAIL.n149 12.8005
R212 VTAIL.n146 VTAIL.n145 12.8005
R213 VTAIL.n98 VTAIL.n97 12.8005
R214 VTAIL.n94 VTAIL.n93 12.8005
R215 VTAIL.n191 VTAIL.n190 12.0247
R216 VTAIL.n203 VTAIL.n160 12.0247
R217 VTAIL.n35 VTAIL.n34 12.0247
R218 VTAIL.n47 VTAIL.n4 12.0247
R219 VTAIL.n153 VTAIL.n110 12.0247
R220 VTAIL.n142 VTAIL.n115 12.0247
R221 VTAIL.n101 VTAIL.n58 12.0247
R222 VTAIL.n90 VTAIL.n63 12.0247
R223 VTAIL.n189 VTAIL.n166 11.249
R224 VTAIL.n204 VTAIL.n158 11.249
R225 VTAIL.n33 VTAIL.n10 11.249
R226 VTAIL.n48 VTAIL.n2 11.249
R227 VTAIL.n154 VTAIL.n108 11.249
R228 VTAIL.n141 VTAIL.n118 11.249
R229 VTAIL.n102 VTAIL.n56 11.249
R230 VTAIL.n89 VTAIL.n66 11.249
R231 VTAIL.n186 VTAIL.n185 10.4732
R232 VTAIL.n30 VTAIL.n29 10.4732
R233 VTAIL.n138 VTAIL.n137 10.4732
R234 VTAIL.n86 VTAIL.n85 10.4732
R235 VTAIL.n174 VTAIL.n173 10.2747
R236 VTAIL.n18 VTAIL.n17 10.2747
R237 VTAIL.n126 VTAIL.n125 10.2747
R238 VTAIL.n74 VTAIL.n73 10.2747
R239 VTAIL.n182 VTAIL.n168 9.69747
R240 VTAIL.n26 VTAIL.n12 9.69747
R241 VTAIL.n134 VTAIL.n120 9.69747
R242 VTAIL.n82 VTAIL.n68 9.69747
R243 VTAIL.n206 VTAIL.n205 9.45567
R244 VTAIL.n50 VTAIL.n49 9.45567
R245 VTAIL.n156 VTAIL.n155 9.45567
R246 VTAIL.n104 VTAIL.n103 9.45567
R247 VTAIL.n205 VTAIL.n204 9.3005
R248 VTAIL.n160 VTAIL.n159 9.3005
R249 VTAIL.n199 VTAIL.n198 9.3005
R250 VTAIL.n172 VTAIL.n171 9.3005
R251 VTAIL.n179 VTAIL.n178 9.3005
R252 VTAIL.n181 VTAIL.n180 9.3005
R253 VTAIL.n168 VTAIL.n167 9.3005
R254 VTAIL.n187 VTAIL.n186 9.3005
R255 VTAIL.n189 VTAIL.n188 9.3005
R256 VTAIL.n190 VTAIL.n163 9.3005
R257 VTAIL.n197 VTAIL.n196 9.3005
R258 VTAIL.n49 VTAIL.n48 9.3005
R259 VTAIL.n4 VTAIL.n3 9.3005
R260 VTAIL.n43 VTAIL.n42 9.3005
R261 VTAIL.n16 VTAIL.n15 9.3005
R262 VTAIL.n23 VTAIL.n22 9.3005
R263 VTAIL.n25 VTAIL.n24 9.3005
R264 VTAIL.n12 VTAIL.n11 9.3005
R265 VTAIL.n31 VTAIL.n30 9.3005
R266 VTAIL.n33 VTAIL.n32 9.3005
R267 VTAIL.n34 VTAIL.n7 9.3005
R268 VTAIL.n41 VTAIL.n40 9.3005
R269 VTAIL.n124 VTAIL.n123 9.3005
R270 VTAIL.n131 VTAIL.n130 9.3005
R271 VTAIL.n133 VTAIL.n132 9.3005
R272 VTAIL.n120 VTAIL.n119 9.3005
R273 VTAIL.n139 VTAIL.n138 9.3005
R274 VTAIL.n141 VTAIL.n140 9.3005
R275 VTAIL.n115 VTAIL.n113 9.3005
R276 VTAIL.n147 VTAIL.n146 9.3005
R277 VTAIL.n155 VTAIL.n154 9.3005
R278 VTAIL.n110 VTAIL.n109 9.3005
R279 VTAIL.n149 VTAIL.n148 9.3005
R280 VTAIL.n72 VTAIL.n71 9.3005
R281 VTAIL.n79 VTAIL.n78 9.3005
R282 VTAIL.n81 VTAIL.n80 9.3005
R283 VTAIL.n68 VTAIL.n67 9.3005
R284 VTAIL.n87 VTAIL.n86 9.3005
R285 VTAIL.n89 VTAIL.n88 9.3005
R286 VTAIL.n63 VTAIL.n61 9.3005
R287 VTAIL.n95 VTAIL.n94 9.3005
R288 VTAIL.n103 VTAIL.n102 9.3005
R289 VTAIL.n58 VTAIL.n57 9.3005
R290 VTAIL.n97 VTAIL.n96 9.3005
R291 VTAIL.n181 VTAIL.n170 8.92171
R292 VTAIL.n25 VTAIL.n14 8.92171
R293 VTAIL.n133 VTAIL.n122 8.92171
R294 VTAIL.n81 VTAIL.n70 8.92171
R295 VTAIL.n178 VTAIL.n177 8.14595
R296 VTAIL.n22 VTAIL.n21 8.14595
R297 VTAIL.n130 VTAIL.n129 8.14595
R298 VTAIL.n78 VTAIL.n77 8.14595
R299 VTAIL.n174 VTAIL.n172 7.3702
R300 VTAIL.n18 VTAIL.n16 7.3702
R301 VTAIL.n126 VTAIL.n124 7.3702
R302 VTAIL.n74 VTAIL.n72 7.3702
R303 VTAIL.n177 VTAIL.n172 5.81868
R304 VTAIL.n21 VTAIL.n16 5.81868
R305 VTAIL.n129 VTAIL.n124 5.81868
R306 VTAIL.n77 VTAIL.n72 5.81868
R307 VTAIL.n178 VTAIL.n170 5.04292
R308 VTAIL.n22 VTAIL.n14 5.04292
R309 VTAIL.n130 VTAIL.n122 5.04292
R310 VTAIL.n78 VTAIL.n70 5.04292
R311 VTAIL.n182 VTAIL.n181 4.26717
R312 VTAIL.n26 VTAIL.n25 4.26717
R313 VTAIL.n134 VTAIL.n133 4.26717
R314 VTAIL.n82 VTAIL.n81 4.26717
R315 VTAIL.n105 VTAIL.n55 3.61257
R316 VTAIL.n157 VTAIL.n107 3.61257
R317 VTAIL.n53 VTAIL.n51 3.61257
R318 VTAIL.n185 VTAIL.n168 3.49141
R319 VTAIL.n29 VTAIL.n12 3.49141
R320 VTAIL.n137 VTAIL.n120 3.49141
R321 VTAIL.n85 VTAIL.n68 3.49141
R322 VTAIL.n173 VTAIL.n171 2.84303
R323 VTAIL.n17 VTAIL.n15 2.84303
R324 VTAIL.n125 VTAIL.n123 2.84303
R325 VTAIL.n73 VTAIL.n71 2.84303
R326 VTAIL.n186 VTAIL.n166 2.71565
R327 VTAIL.n206 VTAIL.n158 2.71565
R328 VTAIL.n30 VTAIL.n10 2.71565
R329 VTAIL.n50 VTAIL.n2 2.71565
R330 VTAIL.n156 VTAIL.n108 2.71565
R331 VTAIL.n138 VTAIL.n118 2.71565
R332 VTAIL.n104 VTAIL.n56 2.71565
R333 VTAIL.n86 VTAIL.n66 2.71565
R334 VTAIL VTAIL.n207 2.65136
R335 VTAIL.n107 VTAIL.n105 2.27636
R336 VTAIL.n51 VTAIL.n1 2.27636
R337 VTAIL.n0 VTAIL.t5 2.10688
R338 VTAIL.n0 VTAIL.t0 2.10688
R339 VTAIL.n52 VTAIL.t10 2.10688
R340 VTAIL.n52 VTAIL.t7 2.10688
R341 VTAIL.n106 VTAIL.t9 2.10688
R342 VTAIL.n106 VTAIL.t6 2.10688
R343 VTAIL.n54 VTAIL.t4 2.10688
R344 VTAIL.n54 VTAIL.t3 2.10688
R345 VTAIL.n191 VTAIL.n189 1.93989
R346 VTAIL.n204 VTAIL.n203 1.93989
R347 VTAIL.n35 VTAIL.n33 1.93989
R348 VTAIL.n48 VTAIL.n47 1.93989
R349 VTAIL.n154 VTAIL.n153 1.93989
R350 VTAIL.n142 VTAIL.n141 1.93989
R351 VTAIL.n102 VTAIL.n101 1.93989
R352 VTAIL.n90 VTAIL.n89 1.93989
R353 VTAIL.n190 VTAIL.n164 1.16414
R354 VTAIL.n200 VTAIL.n160 1.16414
R355 VTAIL.n34 VTAIL.n8 1.16414
R356 VTAIL.n44 VTAIL.n4 1.16414
R357 VTAIL.n150 VTAIL.n110 1.16414
R358 VTAIL.n145 VTAIL.n115 1.16414
R359 VTAIL.n98 VTAIL.n58 1.16414
R360 VTAIL.n93 VTAIL.n63 1.16414
R361 VTAIL VTAIL.n1 0.961707
R362 VTAIL.n196 VTAIL.n195 0.388379
R363 VTAIL.n199 VTAIL.n162 0.388379
R364 VTAIL.n40 VTAIL.n39 0.388379
R365 VTAIL.n43 VTAIL.n6 0.388379
R366 VTAIL.n149 VTAIL.n112 0.388379
R367 VTAIL.n146 VTAIL.n114 0.388379
R368 VTAIL.n97 VTAIL.n60 0.388379
R369 VTAIL.n94 VTAIL.n62 0.388379
R370 VTAIL.n179 VTAIL.n171 0.155672
R371 VTAIL.n180 VTAIL.n179 0.155672
R372 VTAIL.n180 VTAIL.n167 0.155672
R373 VTAIL.n187 VTAIL.n167 0.155672
R374 VTAIL.n188 VTAIL.n187 0.155672
R375 VTAIL.n188 VTAIL.n163 0.155672
R376 VTAIL.n197 VTAIL.n163 0.155672
R377 VTAIL.n198 VTAIL.n197 0.155672
R378 VTAIL.n198 VTAIL.n159 0.155672
R379 VTAIL.n205 VTAIL.n159 0.155672
R380 VTAIL.n23 VTAIL.n15 0.155672
R381 VTAIL.n24 VTAIL.n23 0.155672
R382 VTAIL.n24 VTAIL.n11 0.155672
R383 VTAIL.n31 VTAIL.n11 0.155672
R384 VTAIL.n32 VTAIL.n31 0.155672
R385 VTAIL.n32 VTAIL.n7 0.155672
R386 VTAIL.n41 VTAIL.n7 0.155672
R387 VTAIL.n42 VTAIL.n41 0.155672
R388 VTAIL.n42 VTAIL.n3 0.155672
R389 VTAIL.n49 VTAIL.n3 0.155672
R390 VTAIL.n155 VTAIL.n109 0.155672
R391 VTAIL.n148 VTAIL.n109 0.155672
R392 VTAIL.n148 VTAIL.n147 0.155672
R393 VTAIL.n147 VTAIL.n113 0.155672
R394 VTAIL.n140 VTAIL.n113 0.155672
R395 VTAIL.n140 VTAIL.n139 0.155672
R396 VTAIL.n139 VTAIL.n119 0.155672
R397 VTAIL.n132 VTAIL.n119 0.155672
R398 VTAIL.n132 VTAIL.n131 0.155672
R399 VTAIL.n131 VTAIL.n123 0.155672
R400 VTAIL.n103 VTAIL.n57 0.155672
R401 VTAIL.n96 VTAIL.n57 0.155672
R402 VTAIL.n96 VTAIL.n95 0.155672
R403 VTAIL.n95 VTAIL.n61 0.155672
R404 VTAIL.n88 VTAIL.n61 0.155672
R405 VTAIL.n88 VTAIL.n87 0.155672
R406 VTAIL.n87 VTAIL.n67 0.155672
R407 VTAIL.n80 VTAIL.n67 0.155672
R408 VTAIL.n80 VTAIL.n79 0.155672
R409 VTAIL.n79 VTAIL.n71 0.155672
R410 VDD1.n44 VDD1.n0 289.615
R411 VDD1.n93 VDD1.n49 289.615
R412 VDD1.n45 VDD1.n44 185
R413 VDD1.n43 VDD1.n42 185
R414 VDD1.n4 VDD1.n3 185
R415 VDD1.n8 VDD1.n6 185
R416 VDD1.n37 VDD1.n36 185
R417 VDD1.n35 VDD1.n34 185
R418 VDD1.n10 VDD1.n9 185
R419 VDD1.n29 VDD1.n28 185
R420 VDD1.n27 VDD1.n26 185
R421 VDD1.n14 VDD1.n13 185
R422 VDD1.n21 VDD1.n20 185
R423 VDD1.n19 VDD1.n18 185
R424 VDD1.n66 VDD1.n65 185
R425 VDD1.n68 VDD1.n67 185
R426 VDD1.n61 VDD1.n60 185
R427 VDD1.n74 VDD1.n73 185
R428 VDD1.n76 VDD1.n75 185
R429 VDD1.n57 VDD1.n56 185
R430 VDD1.n83 VDD1.n82 185
R431 VDD1.n84 VDD1.n55 185
R432 VDD1.n86 VDD1.n85 185
R433 VDD1.n53 VDD1.n52 185
R434 VDD1.n92 VDD1.n91 185
R435 VDD1.n94 VDD1.n93 185
R436 VDD1.n17 VDD1.t4 149.524
R437 VDD1.n64 VDD1.t3 149.524
R438 VDD1.n44 VDD1.n43 104.615
R439 VDD1.n43 VDD1.n3 104.615
R440 VDD1.n8 VDD1.n3 104.615
R441 VDD1.n36 VDD1.n8 104.615
R442 VDD1.n36 VDD1.n35 104.615
R443 VDD1.n35 VDD1.n9 104.615
R444 VDD1.n28 VDD1.n9 104.615
R445 VDD1.n28 VDD1.n27 104.615
R446 VDD1.n27 VDD1.n13 104.615
R447 VDD1.n20 VDD1.n13 104.615
R448 VDD1.n20 VDD1.n19 104.615
R449 VDD1.n67 VDD1.n66 104.615
R450 VDD1.n67 VDD1.n60 104.615
R451 VDD1.n74 VDD1.n60 104.615
R452 VDD1.n75 VDD1.n74 104.615
R453 VDD1.n75 VDD1.n56 104.615
R454 VDD1.n83 VDD1.n56 104.615
R455 VDD1.n84 VDD1.n83 104.615
R456 VDD1.n85 VDD1.n84 104.615
R457 VDD1.n85 VDD1.n52 104.615
R458 VDD1.n92 VDD1.n52 104.615
R459 VDD1.n93 VDD1.n92 104.615
R460 VDD1.n99 VDD1.n98 66.9526
R461 VDD1.n101 VDD1.n100 66.1049
R462 VDD1 VDD1.n48 54.7344
R463 VDD1.n99 VDD1.n97 54.6209
R464 VDD1.n19 VDD1.t4 52.3082
R465 VDD1.n66 VDD1.t3 52.3082
R466 VDD1.n101 VDD1.n99 45.947
R467 VDD1.n6 VDD1.n4 13.1884
R468 VDD1.n86 VDD1.n53 13.1884
R469 VDD1.n42 VDD1.n41 12.8005
R470 VDD1.n38 VDD1.n37 12.8005
R471 VDD1.n87 VDD1.n55 12.8005
R472 VDD1.n91 VDD1.n90 12.8005
R473 VDD1.n45 VDD1.n2 12.0247
R474 VDD1.n34 VDD1.n7 12.0247
R475 VDD1.n82 VDD1.n81 12.0247
R476 VDD1.n94 VDD1.n51 12.0247
R477 VDD1.n46 VDD1.n0 11.249
R478 VDD1.n33 VDD1.n10 11.249
R479 VDD1.n80 VDD1.n57 11.249
R480 VDD1.n95 VDD1.n49 11.249
R481 VDD1.n30 VDD1.n29 10.4732
R482 VDD1.n77 VDD1.n76 10.4732
R483 VDD1.n18 VDD1.n17 10.2747
R484 VDD1.n65 VDD1.n64 10.2747
R485 VDD1.n26 VDD1.n12 9.69747
R486 VDD1.n73 VDD1.n59 9.69747
R487 VDD1.n48 VDD1.n47 9.45567
R488 VDD1.n97 VDD1.n96 9.45567
R489 VDD1.n16 VDD1.n15 9.3005
R490 VDD1.n23 VDD1.n22 9.3005
R491 VDD1.n25 VDD1.n24 9.3005
R492 VDD1.n12 VDD1.n11 9.3005
R493 VDD1.n31 VDD1.n30 9.3005
R494 VDD1.n33 VDD1.n32 9.3005
R495 VDD1.n7 VDD1.n5 9.3005
R496 VDD1.n39 VDD1.n38 9.3005
R497 VDD1.n47 VDD1.n46 9.3005
R498 VDD1.n2 VDD1.n1 9.3005
R499 VDD1.n41 VDD1.n40 9.3005
R500 VDD1.n96 VDD1.n95 9.3005
R501 VDD1.n51 VDD1.n50 9.3005
R502 VDD1.n90 VDD1.n89 9.3005
R503 VDD1.n63 VDD1.n62 9.3005
R504 VDD1.n70 VDD1.n69 9.3005
R505 VDD1.n72 VDD1.n71 9.3005
R506 VDD1.n59 VDD1.n58 9.3005
R507 VDD1.n78 VDD1.n77 9.3005
R508 VDD1.n80 VDD1.n79 9.3005
R509 VDD1.n81 VDD1.n54 9.3005
R510 VDD1.n88 VDD1.n87 9.3005
R511 VDD1.n25 VDD1.n14 8.92171
R512 VDD1.n72 VDD1.n61 8.92171
R513 VDD1.n22 VDD1.n21 8.14595
R514 VDD1.n69 VDD1.n68 8.14595
R515 VDD1.n18 VDD1.n16 7.3702
R516 VDD1.n65 VDD1.n63 7.3702
R517 VDD1.n21 VDD1.n16 5.81868
R518 VDD1.n68 VDD1.n63 5.81868
R519 VDD1.n22 VDD1.n14 5.04292
R520 VDD1.n69 VDD1.n61 5.04292
R521 VDD1.n26 VDD1.n25 4.26717
R522 VDD1.n73 VDD1.n72 4.26717
R523 VDD1.n29 VDD1.n12 3.49141
R524 VDD1.n76 VDD1.n59 3.49141
R525 VDD1.n17 VDD1.n15 2.84303
R526 VDD1.n64 VDD1.n62 2.84303
R527 VDD1.n48 VDD1.n0 2.71565
R528 VDD1.n30 VDD1.n10 2.71565
R529 VDD1.n77 VDD1.n57 2.71565
R530 VDD1.n97 VDD1.n49 2.71565
R531 VDD1.n100 VDD1.t2 2.10688
R532 VDD1.n100 VDD1.t1 2.10688
R533 VDD1.n98 VDD1.t0 2.10688
R534 VDD1.n98 VDD1.t5 2.10688
R535 VDD1.n46 VDD1.n45 1.93989
R536 VDD1.n34 VDD1.n33 1.93989
R537 VDD1.n82 VDD1.n80 1.93989
R538 VDD1.n95 VDD1.n94 1.93989
R539 VDD1.n42 VDD1.n2 1.16414
R540 VDD1.n37 VDD1.n7 1.16414
R541 VDD1.n81 VDD1.n55 1.16414
R542 VDD1.n91 VDD1.n51 1.16414
R543 VDD1 VDD1.n101 0.845328
R544 VDD1.n41 VDD1.n4 0.388379
R545 VDD1.n38 VDD1.n6 0.388379
R546 VDD1.n87 VDD1.n86 0.388379
R547 VDD1.n90 VDD1.n53 0.388379
R548 VDD1.n47 VDD1.n1 0.155672
R549 VDD1.n40 VDD1.n1 0.155672
R550 VDD1.n40 VDD1.n39 0.155672
R551 VDD1.n39 VDD1.n5 0.155672
R552 VDD1.n32 VDD1.n5 0.155672
R553 VDD1.n32 VDD1.n31 0.155672
R554 VDD1.n31 VDD1.n11 0.155672
R555 VDD1.n24 VDD1.n11 0.155672
R556 VDD1.n24 VDD1.n23 0.155672
R557 VDD1.n23 VDD1.n15 0.155672
R558 VDD1.n70 VDD1.n62 0.155672
R559 VDD1.n71 VDD1.n70 0.155672
R560 VDD1.n71 VDD1.n58 0.155672
R561 VDD1.n78 VDD1.n58 0.155672
R562 VDD1.n79 VDD1.n78 0.155672
R563 VDD1.n79 VDD1.n54 0.155672
R564 VDD1.n88 VDD1.n54 0.155672
R565 VDD1.n89 VDD1.n88 0.155672
R566 VDD1.n89 VDD1.n50 0.155672
R567 VDD1.n96 VDD1.n50 0.155672
R568 B.n858 B.n857 585
R569 B.n859 B.n858 585
R570 B.n301 B.n144 585
R571 B.n300 B.n299 585
R572 B.n298 B.n297 585
R573 B.n296 B.n295 585
R574 B.n294 B.n293 585
R575 B.n292 B.n291 585
R576 B.n290 B.n289 585
R577 B.n288 B.n287 585
R578 B.n286 B.n285 585
R579 B.n284 B.n283 585
R580 B.n282 B.n281 585
R581 B.n280 B.n279 585
R582 B.n278 B.n277 585
R583 B.n276 B.n275 585
R584 B.n274 B.n273 585
R585 B.n272 B.n271 585
R586 B.n270 B.n269 585
R587 B.n268 B.n267 585
R588 B.n266 B.n265 585
R589 B.n264 B.n263 585
R590 B.n262 B.n261 585
R591 B.n260 B.n259 585
R592 B.n258 B.n257 585
R593 B.n256 B.n255 585
R594 B.n254 B.n253 585
R595 B.n252 B.n251 585
R596 B.n250 B.n249 585
R597 B.n248 B.n247 585
R598 B.n246 B.n245 585
R599 B.n244 B.n243 585
R600 B.n242 B.n241 585
R601 B.n240 B.n239 585
R602 B.n238 B.n237 585
R603 B.n235 B.n234 585
R604 B.n233 B.n232 585
R605 B.n231 B.n230 585
R606 B.n229 B.n228 585
R607 B.n227 B.n226 585
R608 B.n225 B.n224 585
R609 B.n223 B.n222 585
R610 B.n221 B.n220 585
R611 B.n219 B.n218 585
R612 B.n217 B.n216 585
R613 B.n215 B.n214 585
R614 B.n213 B.n212 585
R615 B.n211 B.n210 585
R616 B.n209 B.n208 585
R617 B.n207 B.n206 585
R618 B.n205 B.n204 585
R619 B.n203 B.n202 585
R620 B.n201 B.n200 585
R621 B.n199 B.n198 585
R622 B.n197 B.n196 585
R623 B.n195 B.n194 585
R624 B.n193 B.n192 585
R625 B.n191 B.n190 585
R626 B.n189 B.n188 585
R627 B.n187 B.n186 585
R628 B.n185 B.n184 585
R629 B.n183 B.n182 585
R630 B.n181 B.n180 585
R631 B.n179 B.n178 585
R632 B.n177 B.n176 585
R633 B.n175 B.n174 585
R634 B.n173 B.n172 585
R635 B.n171 B.n170 585
R636 B.n169 B.n168 585
R637 B.n167 B.n166 585
R638 B.n165 B.n164 585
R639 B.n163 B.n162 585
R640 B.n161 B.n160 585
R641 B.n159 B.n158 585
R642 B.n157 B.n156 585
R643 B.n155 B.n154 585
R644 B.n153 B.n152 585
R645 B.n151 B.n150 585
R646 B.n856 B.n105 585
R647 B.n860 B.n105 585
R648 B.n855 B.n104 585
R649 B.n861 B.n104 585
R650 B.n854 B.n853 585
R651 B.n853 B.n100 585
R652 B.n852 B.n99 585
R653 B.n867 B.n99 585
R654 B.n851 B.n98 585
R655 B.n868 B.n98 585
R656 B.n850 B.n97 585
R657 B.n869 B.n97 585
R658 B.n849 B.n848 585
R659 B.n848 B.n93 585
R660 B.n847 B.n92 585
R661 B.n875 B.n92 585
R662 B.n846 B.n91 585
R663 B.n876 B.n91 585
R664 B.n845 B.n90 585
R665 B.n877 B.n90 585
R666 B.n844 B.n843 585
R667 B.n843 B.n86 585
R668 B.n842 B.n85 585
R669 B.n883 B.n85 585
R670 B.n841 B.n84 585
R671 B.n884 B.n84 585
R672 B.n840 B.n83 585
R673 B.n885 B.n83 585
R674 B.n839 B.n838 585
R675 B.n838 B.n79 585
R676 B.n837 B.n78 585
R677 B.n891 B.n78 585
R678 B.n836 B.n77 585
R679 B.n892 B.n77 585
R680 B.n835 B.n76 585
R681 B.n893 B.n76 585
R682 B.n834 B.n833 585
R683 B.n833 B.n72 585
R684 B.n832 B.n71 585
R685 B.n899 B.n71 585
R686 B.n831 B.n70 585
R687 B.n900 B.n70 585
R688 B.n830 B.n69 585
R689 B.n901 B.n69 585
R690 B.n829 B.n828 585
R691 B.n828 B.n65 585
R692 B.n827 B.n64 585
R693 B.n907 B.n64 585
R694 B.n826 B.n63 585
R695 B.n908 B.n63 585
R696 B.n825 B.n62 585
R697 B.n909 B.n62 585
R698 B.n824 B.n823 585
R699 B.n823 B.n58 585
R700 B.n822 B.n57 585
R701 B.n915 B.n57 585
R702 B.n821 B.n56 585
R703 B.n916 B.n56 585
R704 B.n820 B.n55 585
R705 B.n917 B.n55 585
R706 B.n819 B.n818 585
R707 B.n818 B.n51 585
R708 B.n817 B.n50 585
R709 B.n923 B.n50 585
R710 B.n816 B.n49 585
R711 B.n924 B.n49 585
R712 B.n815 B.n48 585
R713 B.n925 B.n48 585
R714 B.n814 B.n813 585
R715 B.n813 B.n44 585
R716 B.n812 B.n43 585
R717 B.n931 B.n43 585
R718 B.n811 B.n42 585
R719 B.n932 B.n42 585
R720 B.n810 B.n41 585
R721 B.n933 B.n41 585
R722 B.n809 B.n808 585
R723 B.n808 B.n37 585
R724 B.n807 B.n36 585
R725 B.n939 B.n36 585
R726 B.n806 B.n35 585
R727 B.n940 B.n35 585
R728 B.n805 B.n34 585
R729 B.n941 B.n34 585
R730 B.n804 B.n803 585
R731 B.n803 B.n30 585
R732 B.n802 B.n29 585
R733 B.n947 B.n29 585
R734 B.n801 B.n28 585
R735 B.n948 B.n28 585
R736 B.n800 B.n27 585
R737 B.n949 B.n27 585
R738 B.n799 B.n798 585
R739 B.n798 B.n23 585
R740 B.n797 B.n22 585
R741 B.n955 B.n22 585
R742 B.n796 B.n21 585
R743 B.n956 B.n21 585
R744 B.n795 B.n20 585
R745 B.n957 B.n20 585
R746 B.n794 B.n793 585
R747 B.n793 B.n16 585
R748 B.n792 B.n15 585
R749 B.n963 B.n15 585
R750 B.n791 B.n14 585
R751 B.n964 B.n14 585
R752 B.n790 B.n13 585
R753 B.n965 B.n13 585
R754 B.n789 B.n788 585
R755 B.n788 B.n12 585
R756 B.n787 B.n786 585
R757 B.n787 B.n8 585
R758 B.n785 B.n7 585
R759 B.n972 B.n7 585
R760 B.n784 B.n6 585
R761 B.n973 B.n6 585
R762 B.n783 B.n5 585
R763 B.n974 B.n5 585
R764 B.n782 B.n781 585
R765 B.n781 B.n4 585
R766 B.n780 B.n302 585
R767 B.n780 B.n779 585
R768 B.n770 B.n303 585
R769 B.n304 B.n303 585
R770 B.n772 B.n771 585
R771 B.n773 B.n772 585
R772 B.n769 B.n309 585
R773 B.n309 B.n308 585
R774 B.n768 B.n767 585
R775 B.n767 B.n766 585
R776 B.n311 B.n310 585
R777 B.n312 B.n311 585
R778 B.n759 B.n758 585
R779 B.n760 B.n759 585
R780 B.n757 B.n317 585
R781 B.n317 B.n316 585
R782 B.n756 B.n755 585
R783 B.n755 B.n754 585
R784 B.n319 B.n318 585
R785 B.n320 B.n319 585
R786 B.n747 B.n746 585
R787 B.n748 B.n747 585
R788 B.n745 B.n325 585
R789 B.n325 B.n324 585
R790 B.n744 B.n743 585
R791 B.n743 B.n742 585
R792 B.n327 B.n326 585
R793 B.n328 B.n327 585
R794 B.n735 B.n734 585
R795 B.n736 B.n735 585
R796 B.n733 B.n333 585
R797 B.n333 B.n332 585
R798 B.n732 B.n731 585
R799 B.n731 B.n730 585
R800 B.n335 B.n334 585
R801 B.n336 B.n335 585
R802 B.n723 B.n722 585
R803 B.n724 B.n723 585
R804 B.n721 B.n341 585
R805 B.n341 B.n340 585
R806 B.n720 B.n719 585
R807 B.n719 B.n718 585
R808 B.n343 B.n342 585
R809 B.n344 B.n343 585
R810 B.n711 B.n710 585
R811 B.n712 B.n711 585
R812 B.n709 B.n349 585
R813 B.n349 B.n348 585
R814 B.n708 B.n707 585
R815 B.n707 B.n706 585
R816 B.n351 B.n350 585
R817 B.n352 B.n351 585
R818 B.n699 B.n698 585
R819 B.n700 B.n699 585
R820 B.n697 B.n357 585
R821 B.n357 B.n356 585
R822 B.n696 B.n695 585
R823 B.n695 B.n694 585
R824 B.n359 B.n358 585
R825 B.n360 B.n359 585
R826 B.n687 B.n686 585
R827 B.n688 B.n687 585
R828 B.n685 B.n365 585
R829 B.n365 B.n364 585
R830 B.n684 B.n683 585
R831 B.n683 B.n682 585
R832 B.n367 B.n366 585
R833 B.n368 B.n367 585
R834 B.n675 B.n674 585
R835 B.n676 B.n675 585
R836 B.n673 B.n373 585
R837 B.n373 B.n372 585
R838 B.n672 B.n671 585
R839 B.n671 B.n670 585
R840 B.n375 B.n374 585
R841 B.n376 B.n375 585
R842 B.n663 B.n662 585
R843 B.n664 B.n663 585
R844 B.n661 B.n381 585
R845 B.n381 B.n380 585
R846 B.n660 B.n659 585
R847 B.n659 B.n658 585
R848 B.n383 B.n382 585
R849 B.n384 B.n383 585
R850 B.n651 B.n650 585
R851 B.n652 B.n651 585
R852 B.n649 B.n389 585
R853 B.n389 B.n388 585
R854 B.n648 B.n647 585
R855 B.n647 B.n646 585
R856 B.n391 B.n390 585
R857 B.n392 B.n391 585
R858 B.n639 B.n638 585
R859 B.n640 B.n639 585
R860 B.n637 B.n397 585
R861 B.n397 B.n396 585
R862 B.n636 B.n635 585
R863 B.n635 B.n634 585
R864 B.n399 B.n398 585
R865 B.n400 B.n399 585
R866 B.n627 B.n626 585
R867 B.n628 B.n627 585
R868 B.n625 B.n405 585
R869 B.n405 B.n404 585
R870 B.n624 B.n623 585
R871 B.n623 B.n622 585
R872 B.n407 B.n406 585
R873 B.n408 B.n407 585
R874 B.n615 B.n614 585
R875 B.n616 B.n615 585
R876 B.n613 B.n413 585
R877 B.n413 B.n412 585
R878 B.n607 B.n606 585
R879 B.n605 B.n453 585
R880 B.n604 B.n452 585
R881 B.n609 B.n452 585
R882 B.n603 B.n602 585
R883 B.n601 B.n600 585
R884 B.n599 B.n598 585
R885 B.n597 B.n596 585
R886 B.n595 B.n594 585
R887 B.n593 B.n592 585
R888 B.n591 B.n590 585
R889 B.n589 B.n588 585
R890 B.n587 B.n586 585
R891 B.n585 B.n584 585
R892 B.n583 B.n582 585
R893 B.n581 B.n580 585
R894 B.n579 B.n578 585
R895 B.n577 B.n576 585
R896 B.n575 B.n574 585
R897 B.n573 B.n572 585
R898 B.n571 B.n570 585
R899 B.n569 B.n568 585
R900 B.n567 B.n566 585
R901 B.n565 B.n564 585
R902 B.n563 B.n562 585
R903 B.n561 B.n560 585
R904 B.n559 B.n558 585
R905 B.n557 B.n556 585
R906 B.n555 B.n554 585
R907 B.n553 B.n552 585
R908 B.n551 B.n550 585
R909 B.n549 B.n548 585
R910 B.n547 B.n546 585
R911 B.n545 B.n544 585
R912 B.n543 B.n542 585
R913 B.n540 B.n539 585
R914 B.n538 B.n537 585
R915 B.n536 B.n535 585
R916 B.n534 B.n533 585
R917 B.n532 B.n531 585
R918 B.n530 B.n529 585
R919 B.n528 B.n527 585
R920 B.n526 B.n525 585
R921 B.n524 B.n523 585
R922 B.n522 B.n521 585
R923 B.n520 B.n519 585
R924 B.n518 B.n517 585
R925 B.n516 B.n515 585
R926 B.n514 B.n513 585
R927 B.n512 B.n511 585
R928 B.n510 B.n509 585
R929 B.n508 B.n507 585
R930 B.n506 B.n505 585
R931 B.n504 B.n503 585
R932 B.n502 B.n501 585
R933 B.n500 B.n499 585
R934 B.n498 B.n497 585
R935 B.n496 B.n495 585
R936 B.n494 B.n493 585
R937 B.n492 B.n491 585
R938 B.n490 B.n489 585
R939 B.n488 B.n487 585
R940 B.n486 B.n485 585
R941 B.n484 B.n483 585
R942 B.n482 B.n481 585
R943 B.n480 B.n479 585
R944 B.n478 B.n477 585
R945 B.n476 B.n475 585
R946 B.n474 B.n473 585
R947 B.n472 B.n471 585
R948 B.n470 B.n469 585
R949 B.n468 B.n467 585
R950 B.n466 B.n465 585
R951 B.n464 B.n463 585
R952 B.n462 B.n461 585
R953 B.n460 B.n459 585
R954 B.n415 B.n414 585
R955 B.n612 B.n611 585
R956 B.n411 B.n410 585
R957 B.n412 B.n411 585
R958 B.n618 B.n617 585
R959 B.n617 B.n616 585
R960 B.n619 B.n409 585
R961 B.n409 B.n408 585
R962 B.n621 B.n620 585
R963 B.n622 B.n621 585
R964 B.n403 B.n402 585
R965 B.n404 B.n403 585
R966 B.n630 B.n629 585
R967 B.n629 B.n628 585
R968 B.n631 B.n401 585
R969 B.n401 B.n400 585
R970 B.n633 B.n632 585
R971 B.n634 B.n633 585
R972 B.n395 B.n394 585
R973 B.n396 B.n395 585
R974 B.n642 B.n641 585
R975 B.n641 B.n640 585
R976 B.n643 B.n393 585
R977 B.n393 B.n392 585
R978 B.n645 B.n644 585
R979 B.n646 B.n645 585
R980 B.n387 B.n386 585
R981 B.n388 B.n387 585
R982 B.n654 B.n653 585
R983 B.n653 B.n652 585
R984 B.n655 B.n385 585
R985 B.n385 B.n384 585
R986 B.n657 B.n656 585
R987 B.n658 B.n657 585
R988 B.n379 B.n378 585
R989 B.n380 B.n379 585
R990 B.n666 B.n665 585
R991 B.n665 B.n664 585
R992 B.n667 B.n377 585
R993 B.n377 B.n376 585
R994 B.n669 B.n668 585
R995 B.n670 B.n669 585
R996 B.n371 B.n370 585
R997 B.n372 B.n371 585
R998 B.n678 B.n677 585
R999 B.n677 B.n676 585
R1000 B.n679 B.n369 585
R1001 B.n369 B.n368 585
R1002 B.n681 B.n680 585
R1003 B.n682 B.n681 585
R1004 B.n363 B.n362 585
R1005 B.n364 B.n363 585
R1006 B.n690 B.n689 585
R1007 B.n689 B.n688 585
R1008 B.n691 B.n361 585
R1009 B.n361 B.n360 585
R1010 B.n693 B.n692 585
R1011 B.n694 B.n693 585
R1012 B.n355 B.n354 585
R1013 B.n356 B.n355 585
R1014 B.n702 B.n701 585
R1015 B.n701 B.n700 585
R1016 B.n703 B.n353 585
R1017 B.n353 B.n352 585
R1018 B.n705 B.n704 585
R1019 B.n706 B.n705 585
R1020 B.n347 B.n346 585
R1021 B.n348 B.n347 585
R1022 B.n714 B.n713 585
R1023 B.n713 B.n712 585
R1024 B.n715 B.n345 585
R1025 B.n345 B.n344 585
R1026 B.n717 B.n716 585
R1027 B.n718 B.n717 585
R1028 B.n339 B.n338 585
R1029 B.n340 B.n339 585
R1030 B.n726 B.n725 585
R1031 B.n725 B.n724 585
R1032 B.n727 B.n337 585
R1033 B.n337 B.n336 585
R1034 B.n729 B.n728 585
R1035 B.n730 B.n729 585
R1036 B.n331 B.n330 585
R1037 B.n332 B.n331 585
R1038 B.n738 B.n737 585
R1039 B.n737 B.n736 585
R1040 B.n739 B.n329 585
R1041 B.n329 B.n328 585
R1042 B.n741 B.n740 585
R1043 B.n742 B.n741 585
R1044 B.n323 B.n322 585
R1045 B.n324 B.n323 585
R1046 B.n750 B.n749 585
R1047 B.n749 B.n748 585
R1048 B.n751 B.n321 585
R1049 B.n321 B.n320 585
R1050 B.n753 B.n752 585
R1051 B.n754 B.n753 585
R1052 B.n315 B.n314 585
R1053 B.n316 B.n315 585
R1054 B.n762 B.n761 585
R1055 B.n761 B.n760 585
R1056 B.n763 B.n313 585
R1057 B.n313 B.n312 585
R1058 B.n765 B.n764 585
R1059 B.n766 B.n765 585
R1060 B.n307 B.n306 585
R1061 B.n308 B.n307 585
R1062 B.n775 B.n774 585
R1063 B.n774 B.n773 585
R1064 B.n776 B.n305 585
R1065 B.n305 B.n304 585
R1066 B.n778 B.n777 585
R1067 B.n779 B.n778 585
R1068 B.n3 B.n0 585
R1069 B.n4 B.n3 585
R1070 B.n971 B.n1 585
R1071 B.n972 B.n971 585
R1072 B.n970 B.n969 585
R1073 B.n970 B.n8 585
R1074 B.n968 B.n9 585
R1075 B.n12 B.n9 585
R1076 B.n967 B.n966 585
R1077 B.n966 B.n965 585
R1078 B.n11 B.n10 585
R1079 B.n964 B.n11 585
R1080 B.n962 B.n961 585
R1081 B.n963 B.n962 585
R1082 B.n960 B.n17 585
R1083 B.n17 B.n16 585
R1084 B.n959 B.n958 585
R1085 B.n958 B.n957 585
R1086 B.n19 B.n18 585
R1087 B.n956 B.n19 585
R1088 B.n954 B.n953 585
R1089 B.n955 B.n954 585
R1090 B.n952 B.n24 585
R1091 B.n24 B.n23 585
R1092 B.n951 B.n950 585
R1093 B.n950 B.n949 585
R1094 B.n26 B.n25 585
R1095 B.n948 B.n26 585
R1096 B.n946 B.n945 585
R1097 B.n947 B.n946 585
R1098 B.n944 B.n31 585
R1099 B.n31 B.n30 585
R1100 B.n943 B.n942 585
R1101 B.n942 B.n941 585
R1102 B.n33 B.n32 585
R1103 B.n940 B.n33 585
R1104 B.n938 B.n937 585
R1105 B.n939 B.n938 585
R1106 B.n936 B.n38 585
R1107 B.n38 B.n37 585
R1108 B.n935 B.n934 585
R1109 B.n934 B.n933 585
R1110 B.n40 B.n39 585
R1111 B.n932 B.n40 585
R1112 B.n930 B.n929 585
R1113 B.n931 B.n930 585
R1114 B.n928 B.n45 585
R1115 B.n45 B.n44 585
R1116 B.n927 B.n926 585
R1117 B.n926 B.n925 585
R1118 B.n47 B.n46 585
R1119 B.n924 B.n47 585
R1120 B.n922 B.n921 585
R1121 B.n923 B.n922 585
R1122 B.n920 B.n52 585
R1123 B.n52 B.n51 585
R1124 B.n919 B.n918 585
R1125 B.n918 B.n917 585
R1126 B.n54 B.n53 585
R1127 B.n916 B.n54 585
R1128 B.n914 B.n913 585
R1129 B.n915 B.n914 585
R1130 B.n912 B.n59 585
R1131 B.n59 B.n58 585
R1132 B.n911 B.n910 585
R1133 B.n910 B.n909 585
R1134 B.n61 B.n60 585
R1135 B.n908 B.n61 585
R1136 B.n906 B.n905 585
R1137 B.n907 B.n906 585
R1138 B.n904 B.n66 585
R1139 B.n66 B.n65 585
R1140 B.n903 B.n902 585
R1141 B.n902 B.n901 585
R1142 B.n68 B.n67 585
R1143 B.n900 B.n68 585
R1144 B.n898 B.n897 585
R1145 B.n899 B.n898 585
R1146 B.n896 B.n73 585
R1147 B.n73 B.n72 585
R1148 B.n895 B.n894 585
R1149 B.n894 B.n893 585
R1150 B.n75 B.n74 585
R1151 B.n892 B.n75 585
R1152 B.n890 B.n889 585
R1153 B.n891 B.n890 585
R1154 B.n888 B.n80 585
R1155 B.n80 B.n79 585
R1156 B.n887 B.n886 585
R1157 B.n886 B.n885 585
R1158 B.n82 B.n81 585
R1159 B.n884 B.n82 585
R1160 B.n882 B.n881 585
R1161 B.n883 B.n882 585
R1162 B.n880 B.n87 585
R1163 B.n87 B.n86 585
R1164 B.n879 B.n878 585
R1165 B.n878 B.n877 585
R1166 B.n89 B.n88 585
R1167 B.n876 B.n89 585
R1168 B.n874 B.n873 585
R1169 B.n875 B.n874 585
R1170 B.n872 B.n94 585
R1171 B.n94 B.n93 585
R1172 B.n871 B.n870 585
R1173 B.n870 B.n869 585
R1174 B.n96 B.n95 585
R1175 B.n868 B.n96 585
R1176 B.n866 B.n865 585
R1177 B.n867 B.n866 585
R1178 B.n864 B.n101 585
R1179 B.n101 B.n100 585
R1180 B.n863 B.n862 585
R1181 B.n862 B.n861 585
R1182 B.n103 B.n102 585
R1183 B.n860 B.n103 585
R1184 B.n975 B.n974 585
R1185 B.n973 B.n2 585
R1186 B.n150 B.n103 526.135
R1187 B.n858 B.n105 526.135
R1188 B.n611 B.n413 526.135
R1189 B.n607 B.n411 526.135
R1190 B.n145 B.t15 318.748
R1191 B.n456 B.t12 318.748
R1192 B.n147 B.t18 318.748
R1193 B.n454 B.t9 318.748
R1194 B.n147 B.t17 268.079
R1195 B.n145 B.t13 268.079
R1196 B.n456 B.t10 268.079
R1197 B.n454 B.t6 268.079
R1198 B.n859 B.n143 256.663
R1199 B.n859 B.n142 256.663
R1200 B.n859 B.n141 256.663
R1201 B.n859 B.n140 256.663
R1202 B.n859 B.n139 256.663
R1203 B.n859 B.n138 256.663
R1204 B.n859 B.n137 256.663
R1205 B.n859 B.n136 256.663
R1206 B.n859 B.n135 256.663
R1207 B.n859 B.n134 256.663
R1208 B.n859 B.n133 256.663
R1209 B.n859 B.n132 256.663
R1210 B.n859 B.n131 256.663
R1211 B.n859 B.n130 256.663
R1212 B.n859 B.n129 256.663
R1213 B.n859 B.n128 256.663
R1214 B.n859 B.n127 256.663
R1215 B.n859 B.n126 256.663
R1216 B.n859 B.n125 256.663
R1217 B.n859 B.n124 256.663
R1218 B.n859 B.n123 256.663
R1219 B.n859 B.n122 256.663
R1220 B.n859 B.n121 256.663
R1221 B.n859 B.n120 256.663
R1222 B.n859 B.n119 256.663
R1223 B.n859 B.n118 256.663
R1224 B.n859 B.n117 256.663
R1225 B.n859 B.n116 256.663
R1226 B.n859 B.n115 256.663
R1227 B.n859 B.n114 256.663
R1228 B.n859 B.n113 256.663
R1229 B.n859 B.n112 256.663
R1230 B.n859 B.n111 256.663
R1231 B.n859 B.n110 256.663
R1232 B.n859 B.n109 256.663
R1233 B.n859 B.n108 256.663
R1234 B.n859 B.n107 256.663
R1235 B.n859 B.n106 256.663
R1236 B.n609 B.n608 256.663
R1237 B.n609 B.n416 256.663
R1238 B.n609 B.n417 256.663
R1239 B.n609 B.n418 256.663
R1240 B.n609 B.n419 256.663
R1241 B.n609 B.n420 256.663
R1242 B.n609 B.n421 256.663
R1243 B.n609 B.n422 256.663
R1244 B.n609 B.n423 256.663
R1245 B.n609 B.n424 256.663
R1246 B.n609 B.n425 256.663
R1247 B.n609 B.n426 256.663
R1248 B.n609 B.n427 256.663
R1249 B.n609 B.n428 256.663
R1250 B.n609 B.n429 256.663
R1251 B.n609 B.n430 256.663
R1252 B.n609 B.n431 256.663
R1253 B.n609 B.n432 256.663
R1254 B.n609 B.n433 256.663
R1255 B.n609 B.n434 256.663
R1256 B.n609 B.n435 256.663
R1257 B.n609 B.n436 256.663
R1258 B.n609 B.n437 256.663
R1259 B.n609 B.n438 256.663
R1260 B.n609 B.n439 256.663
R1261 B.n609 B.n440 256.663
R1262 B.n609 B.n441 256.663
R1263 B.n609 B.n442 256.663
R1264 B.n609 B.n443 256.663
R1265 B.n609 B.n444 256.663
R1266 B.n609 B.n445 256.663
R1267 B.n609 B.n446 256.663
R1268 B.n609 B.n447 256.663
R1269 B.n609 B.n448 256.663
R1270 B.n609 B.n449 256.663
R1271 B.n609 B.n450 256.663
R1272 B.n609 B.n451 256.663
R1273 B.n610 B.n609 256.663
R1274 B.n977 B.n976 256.663
R1275 B.n146 B.t16 237.487
R1276 B.n457 B.t11 237.487
R1277 B.n148 B.t19 237.487
R1278 B.n455 B.t8 237.487
R1279 B.n154 B.n153 163.367
R1280 B.n158 B.n157 163.367
R1281 B.n162 B.n161 163.367
R1282 B.n166 B.n165 163.367
R1283 B.n170 B.n169 163.367
R1284 B.n174 B.n173 163.367
R1285 B.n178 B.n177 163.367
R1286 B.n182 B.n181 163.367
R1287 B.n186 B.n185 163.367
R1288 B.n190 B.n189 163.367
R1289 B.n194 B.n193 163.367
R1290 B.n198 B.n197 163.367
R1291 B.n202 B.n201 163.367
R1292 B.n206 B.n205 163.367
R1293 B.n210 B.n209 163.367
R1294 B.n214 B.n213 163.367
R1295 B.n218 B.n217 163.367
R1296 B.n222 B.n221 163.367
R1297 B.n226 B.n225 163.367
R1298 B.n230 B.n229 163.367
R1299 B.n234 B.n233 163.367
R1300 B.n239 B.n238 163.367
R1301 B.n243 B.n242 163.367
R1302 B.n247 B.n246 163.367
R1303 B.n251 B.n250 163.367
R1304 B.n255 B.n254 163.367
R1305 B.n259 B.n258 163.367
R1306 B.n263 B.n262 163.367
R1307 B.n267 B.n266 163.367
R1308 B.n271 B.n270 163.367
R1309 B.n275 B.n274 163.367
R1310 B.n279 B.n278 163.367
R1311 B.n283 B.n282 163.367
R1312 B.n287 B.n286 163.367
R1313 B.n291 B.n290 163.367
R1314 B.n295 B.n294 163.367
R1315 B.n299 B.n298 163.367
R1316 B.n858 B.n144 163.367
R1317 B.n615 B.n413 163.367
R1318 B.n615 B.n407 163.367
R1319 B.n623 B.n407 163.367
R1320 B.n623 B.n405 163.367
R1321 B.n627 B.n405 163.367
R1322 B.n627 B.n399 163.367
R1323 B.n635 B.n399 163.367
R1324 B.n635 B.n397 163.367
R1325 B.n639 B.n397 163.367
R1326 B.n639 B.n391 163.367
R1327 B.n647 B.n391 163.367
R1328 B.n647 B.n389 163.367
R1329 B.n651 B.n389 163.367
R1330 B.n651 B.n383 163.367
R1331 B.n659 B.n383 163.367
R1332 B.n659 B.n381 163.367
R1333 B.n663 B.n381 163.367
R1334 B.n663 B.n375 163.367
R1335 B.n671 B.n375 163.367
R1336 B.n671 B.n373 163.367
R1337 B.n675 B.n373 163.367
R1338 B.n675 B.n367 163.367
R1339 B.n683 B.n367 163.367
R1340 B.n683 B.n365 163.367
R1341 B.n687 B.n365 163.367
R1342 B.n687 B.n359 163.367
R1343 B.n695 B.n359 163.367
R1344 B.n695 B.n357 163.367
R1345 B.n699 B.n357 163.367
R1346 B.n699 B.n351 163.367
R1347 B.n707 B.n351 163.367
R1348 B.n707 B.n349 163.367
R1349 B.n711 B.n349 163.367
R1350 B.n711 B.n343 163.367
R1351 B.n719 B.n343 163.367
R1352 B.n719 B.n341 163.367
R1353 B.n723 B.n341 163.367
R1354 B.n723 B.n335 163.367
R1355 B.n731 B.n335 163.367
R1356 B.n731 B.n333 163.367
R1357 B.n735 B.n333 163.367
R1358 B.n735 B.n327 163.367
R1359 B.n743 B.n327 163.367
R1360 B.n743 B.n325 163.367
R1361 B.n747 B.n325 163.367
R1362 B.n747 B.n319 163.367
R1363 B.n755 B.n319 163.367
R1364 B.n755 B.n317 163.367
R1365 B.n759 B.n317 163.367
R1366 B.n759 B.n311 163.367
R1367 B.n767 B.n311 163.367
R1368 B.n767 B.n309 163.367
R1369 B.n772 B.n309 163.367
R1370 B.n772 B.n303 163.367
R1371 B.n780 B.n303 163.367
R1372 B.n781 B.n780 163.367
R1373 B.n781 B.n5 163.367
R1374 B.n6 B.n5 163.367
R1375 B.n7 B.n6 163.367
R1376 B.n787 B.n7 163.367
R1377 B.n788 B.n787 163.367
R1378 B.n788 B.n13 163.367
R1379 B.n14 B.n13 163.367
R1380 B.n15 B.n14 163.367
R1381 B.n793 B.n15 163.367
R1382 B.n793 B.n20 163.367
R1383 B.n21 B.n20 163.367
R1384 B.n22 B.n21 163.367
R1385 B.n798 B.n22 163.367
R1386 B.n798 B.n27 163.367
R1387 B.n28 B.n27 163.367
R1388 B.n29 B.n28 163.367
R1389 B.n803 B.n29 163.367
R1390 B.n803 B.n34 163.367
R1391 B.n35 B.n34 163.367
R1392 B.n36 B.n35 163.367
R1393 B.n808 B.n36 163.367
R1394 B.n808 B.n41 163.367
R1395 B.n42 B.n41 163.367
R1396 B.n43 B.n42 163.367
R1397 B.n813 B.n43 163.367
R1398 B.n813 B.n48 163.367
R1399 B.n49 B.n48 163.367
R1400 B.n50 B.n49 163.367
R1401 B.n818 B.n50 163.367
R1402 B.n818 B.n55 163.367
R1403 B.n56 B.n55 163.367
R1404 B.n57 B.n56 163.367
R1405 B.n823 B.n57 163.367
R1406 B.n823 B.n62 163.367
R1407 B.n63 B.n62 163.367
R1408 B.n64 B.n63 163.367
R1409 B.n828 B.n64 163.367
R1410 B.n828 B.n69 163.367
R1411 B.n70 B.n69 163.367
R1412 B.n71 B.n70 163.367
R1413 B.n833 B.n71 163.367
R1414 B.n833 B.n76 163.367
R1415 B.n77 B.n76 163.367
R1416 B.n78 B.n77 163.367
R1417 B.n838 B.n78 163.367
R1418 B.n838 B.n83 163.367
R1419 B.n84 B.n83 163.367
R1420 B.n85 B.n84 163.367
R1421 B.n843 B.n85 163.367
R1422 B.n843 B.n90 163.367
R1423 B.n91 B.n90 163.367
R1424 B.n92 B.n91 163.367
R1425 B.n848 B.n92 163.367
R1426 B.n848 B.n97 163.367
R1427 B.n98 B.n97 163.367
R1428 B.n99 B.n98 163.367
R1429 B.n853 B.n99 163.367
R1430 B.n853 B.n104 163.367
R1431 B.n105 B.n104 163.367
R1432 B.n453 B.n452 163.367
R1433 B.n602 B.n452 163.367
R1434 B.n600 B.n599 163.367
R1435 B.n596 B.n595 163.367
R1436 B.n592 B.n591 163.367
R1437 B.n588 B.n587 163.367
R1438 B.n584 B.n583 163.367
R1439 B.n580 B.n579 163.367
R1440 B.n576 B.n575 163.367
R1441 B.n572 B.n571 163.367
R1442 B.n568 B.n567 163.367
R1443 B.n564 B.n563 163.367
R1444 B.n560 B.n559 163.367
R1445 B.n556 B.n555 163.367
R1446 B.n552 B.n551 163.367
R1447 B.n548 B.n547 163.367
R1448 B.n544 B.n543 163.367
R1449 B.n539 B.n538 163.367
R1450 B.n535 B.n534 163.367
R1451 B.n531 B.n530 163.367
R1452 B.n527 B.n526 163.367
R1453 B.n523 B.n522 163.367
R1454 B.n519 B.n518 163.367
R1455 B.n515 B.n514 163.367
R1456 B.n511 B.n510 163.367
R1457 B.n507 B.n506 163.367
R1458 B.n503 B.n502 163.367
R1459 B.n499 B.n498 163.367
R1460 B.n495 B.n494 163.367
R1461 B.n491 B.n490 163.367
R1462 B.n487 B.n486 163.367
R1463 B.n483 B.n482 163.367
R1464 B.n479 B.n478 163.367
R1465 B.n475 B.n474 163.367
R1466 B.n471 B.n470 163.367
R1467 B.n467 B.n466 163.367
R1468 B.n463 B.n462 163.367
R1469 B.n459 B.n415 163.367
R1470 B.n617 B.n411 163.367
R1471 B.n617 B.n409 163.367
R1472 B.n621 B.n409 163.367
R1473 B.n621 B.n403 163.367
R1474 B.n629 B.n403 163.367
R1475 B.n629 B.n401 163.367
R1476 B.n633 B.n401 163.367
R1477 B.n633 B.n395 163.367
R1478 B.n641 B.n395 163.367
R1479 B.n641 B.n393 163.367
R1480 B.n645 B.n393 163.367
R1481 B.n645 B.n387 163.367
R1482 B.n653 B.n387 163.367
R1483 B.n653 B.n385 163.367
R1484 B.n657 B.n385 163.367
R1485 B.n657 B.n379 163.367
R1486 B.n665 B.n379 163.367
R1487 B.n665 B.n377 163.367
R1488 B.n669 B.n377 163.367
R1489 B.n669 B.n371 163.367
R1490 B.n677 B.n371 163.367
R1491 B.n677 B.n369 163.367
R1492 B.n681 B.n369 163.367
R1493 B.n681 B.n363 163.367
R1494 B.n689 B.n363 163.367
R1495 B.n689 B.n361 163.367
R1496 B.n693 B.n361 163.367
R1497 B.n693 B.n355 163.367
R1498 B.n701 B.n355 163.367
R1499 B.n701 B.n353 163.367
R1500 B.n705 B.n353 163.367
R1501 B.n705 B.n347 163.367
R1502 B.n713 B.n347 163.367
R1503 B.n713 B.n345 163.367
R1504 B.n717 B.n345 163.367
R1505 B.n717 B.n339 163.367
R1506 B.n725 B.n339 163.367
R1507 B.n725 B.n337 163.367
R1508 B.n729 B.n337 163.367
R1509 B.n729 B.n331 163.367
R1510 B.n737 B.n331 163.367
R1511 B.n737 B.n329 163.367
R1512 B.n741 B.n329 163.367
R1513 B.n741 B.n323 163.367
R1514 B.n749 B.n323 163.367
R1515 B.n749 B.n321 163.367
R1516 B.n753 B.n321 163.367
R1517 B.n753 B.n315 163.367
R1518 B.n761 B.n315 163.367
R1519 B.n761 B.n313 163.367
R1520 B.n765 B.n313 163.367
R1521 B.n765 B.n307 163.367
R1522 B.n774 B.n307 163.367
R1523 B.n774 B.n305 163.367
R1524 B.n778 B.n305 163.367
R1525 B.n778 B.n3 163.367
R1526 B.n975 B.n3 163.367
R1527 B.n971 B.n2 163.367
R1528 B.n971 B.n970 163.367
R1529 B.n970 B.n9 163.367
R1530 B.n966 B.n9 163.367
R1531 B.n966 B.n11 163.367
R1532 B.n962 B.n11 163.367
R1533 B.n962 B.n17 163.367
R1534 B.n958 B.n17 163.367
R1535 B.n958 B.n19 163.367
R1536 B.n954 B.n19 163.367
R1537 B.n954 B.n24 163.367
R1538 B.n950 B.n24 163.367
R1539 B.n950 B.n26 163.367
R1540 B.n946 B.n26 163.367
R1541 B.n946 B.n31 163.367
R1542 B.n942 B.n31 163.367
R1543 B.n942 B.n33 163.367
R1544 B.n938 B.n33 163.367
R1545 B.n938 B.n38 163.367
R1546 B.n934 B.n38 163.367
R1547 B.n934 B.n40 163.367
R1548 B.n930 B.n40 163.367
R1549 B.n930 B.n45 163.367
R1550 B.n926 B.n45 163.367
R1551 B.n926 B.n47 163.367
R1552 B.n922 B.n47 163.367
R1553 B.n922 B.n52 163.367
R1554 B.n918 B.n52 163.367
R1555 B.n918 B.n54 163.367
R1556 B.n914 B.n54 163.367
R1557 B.n914 B.n59 163.367
R1558 B.n910 B.n59 163.367
R1559 B.n910 B.n61 163.367
R1560 B.n906 B.n61 163.367
R1561 B.n906 B.n66 163.367
R1562 B.n902 B.n66 163.367
R1563 B.n902 B.n68 163.367
R1564 B.n898 B.n68 163.367
R1565 B.n898 B.n73 163.367
R1566 B.n894 B.n73 163.367
R1567 B.n894 B.n75 163.367
R1568 B.n890 B.n75 163.367
R1569 B.n890 B.n80 163.367
R1570 B.n886 B.n80 163.367
R1571 B.n886 B.n82 163.367
R1572 B.n882 B.n82 163.367
R1573 B.n882 B.n87 163.367
R1574 B.n878 B.n87 163.367
R1575 B.n878 B.n89 163.367
R1576 B.n874 B.n89 163.367
R1577 B.n874 B.n94 163.367
R1578 B.n870 B.n94 163.367
R1579 B.n870 B.n96 163.367
R1580 B.n866 B.n96 163.367
R1581 B.n866 B.n101 163.367
R1582 B.n862 B.n101 163.367
R1583 B.n862 B.n103 163.367
R1584 B.n609 B.n412 87.7007
R1585 B.n860 B.n859 87.7007
R1586 B.n148 B.n147 81.2611
R1587 B.n146 B.n145 81.2611
R1588 B.n457 B.n456 81.2611
R1589 B.n455 B.n454 81.2611
R1590 B.n150 B.n106 71.676
R1591 B.n154 B.n107 71.676
R1592 B.n158 B.n108 71.676
R1593 B.n162 B.n109 71.676
R1594 B.n166 B.n110 71.676
R1595 B.n170 B.n111 71.676
R1596 B.n174 B.n112 71.676
R1597 B.n178 B.n113 71.676
R1598 B.n182 B.n114 71.676
R1599 B.n186 B.n115 71.676
R1600 B.n190 B.n116 71.676
R1601 B.n194 B.n117 71.676
R1602 B.n198 B.n118 71.676
R1603 B.n202 B.n119 71.676
R1604 B.n206 B.n120 71.676
R1605 B.n210 B.n121 71.676
R1606 B.n214 B.n122 71.676
R1607 B.n218 B.n123 71.676
R1608 B.n222 B.n124 71.676
R1609 B.n226 B.n125 71.676
R1610 B.n230 B.n126 71.676
R1611 B.n234 B.n127 71.676
R1612 B.n239 B.n128 71.676
R1613 B.n243 B.n129 71.676
R1614 B.n247 B.n130 71.676
R1615 B.n251 B.n131 71.676
R1616 B.n255 B.n132 71.676
R1617 B.n259 B.n133 71.676
R1618 B.n263 B.n134 71.676
R1619 B.n267 B.n135 71.676
R1620 B.n271 B.n136 71.676
R1621 B.n275 B.n137 71.676
R1622 B.n279 B.n138 71.676
R1623 B.n283 B.n139 71.676
R1624 B.n287 B.n140 71.676
R1625 B.n291 B.n141 71.676
R1626 B.n295 B.n142 71.676
R1627 B.n299 B.n143 71.676
R1628 B.n144 B.n143 71.676
R1629 B.n298 B.n142 71.676
R1630 B.n294 B.n141 71.676
R1631 B.n290 B.n140 71.676
R1632 B.n286 B.n139 71.676
R1633 B.n282 B.n138 71.676
R1634 B.n278 B.n137 71.676
R1635 B.n274 B.n136 71.676
R1636 B.n270 B.n135 71.676
R1637 B.n266 B.n134 71.676
R1638 B.n262 B.n133 71.676
R1639 B.n258 B.n132 71.676
R1640 B.n254 B.n131 71.676
R1641 B.n250 B.n130 71.676
R1642 B.n246 B.n129 71.676
R1643 B.n242 B.n128 71.676
R1644 B.n238 B.n127 71.676
R1645 B.n233 B.n126 71.676
R1646 B.n229 B.n125 71.676
R1647 B.n225 B.n124 71.676
R1648 B.n221 B.n123 71.676
R1649 B.n217 B.n122 71.676
R1650 B.n213 B.n121 71.676
R1651 B.n209 B.n120 71.676
R1652 B.n205 B.n119 71.676
R1653 B.n201 B.n118 71.676
R1654 B.n197 B.n117 71.676
R1655 B.n193 B.n116 71.676
R1656 B.n189 B.n115 71.676
R1657 B.n185 B.n114 71.676
R1658 B.n181 B.n113 71.676
R1659 B.n177 B.n112 71.676
R1660 B.n173 B.n111 71.676
R1661 B.n169 B.n110 71.676
R1662 B.n165 B.n109 71.676
R1663 B.n161 B.n108 71.676
R1664 B.n157 B.n107 71.676
R1665 B.n153 B.n106 71.676
R1666 B.n608 B.n607 71.676
R1667 B.n602 B.n416 71.676
R1668 B.n599 B.n417 71.676
R1669 B.n595 B.n418 71.676
R1670 B.n591 B.n419 71.676
R1671 B.n587 B.n420 71.676
R1672 B.n583 B.n421 71.676
R1673 B.n579 B.n422 71.676
R1674 B.n575 B.n423 71.676
R1675 B.n571 B.n424 71.676
R1676 B.n567 B.n425 71.676
R1677 B.n563 B.n426 71.676
R1678 B.n559 B.n427 71.676
R1679 B.n555 B.n428 71.676
R1680 B.n551 B.n429 71.676
R1681 B.n547 B.n430 71.676
R1682 B.n543 B.n431 71.676
R1683 B.n538 B.n432 71.676
R1684 B.n534 B.n433 71.676
R1685 B.n530 B.n434 71.676
R1686 B.n526 B.n435 71.676
R1687 B.n522 B.n436 71.676
R1688 B.n518 B.n437 71.676
R1689 B.n514 B.n438 71.676
R1690 B.n510 B.n439 71.676
R1691 B.n506 B.n440 71.676
R1692 B.n502 B.n441 71.676
R1693 B.n498 B.n442 71.676
R1694 B.n494 B.n443 71.676
R1695 B.n490 B.n444 71.676
R1696 B.n486 B.n445 71.676
R1697 B.n482 B.n446 71.676
R1698 B.n478 B.n447 71.676
R1699 B.n474 B.n448 71.676
R1700 B.n470 B.n449 71.676
R1701 B.n466 B.n450 71.676
R1702 B.n462 B.n451 71.676
R1703 B.n610 B.n415 71.676
R1704 B.n608 B.n453 71.676
R1705 B.n600 B.n416 71.676
R1706 B.n596 B.n417 71.676
R1707 B.n592 B.n418 71.676
R1708 B.n588 B.n419 71.676
R1709 B.n584 B.n420 71.676
R1710 B.n580 B.n421 71.676
R1711 B.n576 B.n422 71.676
R1712 B.n572 B.n423 71.676
R1713 B.n568 B.n424 71.676
R1714 B.n564 B.n425 71.676
R1715 B.n560 B.n426 71.676
R1716 B.n556 B.n427 71.676
R1717 B.n552 B.n428 71.676
R1718 B.n548 B.n429 71.676
R1719 B.n544 B.n430 71.676
R1720 B.n539 B.n431 71.676
R1721 B.n535 B.n432 71.676
R1722 B.n531 B.n433 71.676
R1723 B.n527 B.n434 71.676
R1724 B.n523 B.n435 71.676
R1725 B.n519 B.n436 71.676
R1726 B.n515 B.n437 71.676
R1727 B.n511 B.n438 71.676
R1728 B.n507 B.n439 71.676
R1729 B.n503 B.n440 71.676
R1730 B.n499 B.n441 71.676
R1731 B.n495 B.n442 71.676
R1732 B.n491 B.n443 71.676
R1733 B.n487 B.n444 71.676
R1734 B.n483 B.n445 71.676
R1735 B.n479 B.n446 71.676
R1736 B.n475 B.n447 71.676
R1737 B.n471 B.n448 71.676
R1738 B.n467 B.n449 71.676
R1739 B.n463 B.n450 71.676
R1740 B.n459 B.n451 71.676
R1741 B.n611 B.n610 71.676
R1742 B.n976 B.n975 71.676
R1743 B.n976 B.n2 71.676
R1744 B.n149 B.n148 59.5399
R1745 B.n236 B.n146 59.5399
R1746 B.n458 B.n457 59.5399
R1747 B.n541 B.n455 59.5399
R1748 B.n616 B.n412 50.9715
R1749 B.n616 B.n408 50.9715
R1750 B.n622 B.n408 50.9715
R1751 B.n622 B.n404 50.9715
R1752 B.n628 B.n404 50.9715
R1753 B.n628 B.n400 50.9715
R1754 B.n634 B.n400 50.9715
R1755 B.n634 B.n396 50.9715
R1756 B.n640 B.n396 50.9715
R1757 B.n646 B.n392 50.9715
R1758 B.n646 B.n388 50.9715
R1759 B.n652 B.n388 50.9715
R1760 B.n652 B.n384 50.9715
R1761 B.n658 B.n384 50.9715
R1762 B.n658 B.n380 50.9715
R1763 B.n664 B.n380 50.9715
R1764 B.n664 B.n376 50.9715
R1765 B.n670 B.n376 50.9715
R1766 B.n670 B.n372 50.9715
R1767 B.n676 B.n372 50.9715
R1768 B.n676 B.n368 50.9715
R1769 B.n682 B.n368 50.9715
R1770 B.n682 B.n364 50.9715
R1771 B.n688 B.n364 50.9715
R1772 B.n694 B.n360 50.9715
R1773 B.n694 B.n356 50.9715
R1774 B.n700 B.n356 50.9715
R1775 B.n700 B.n352 50.9715
R1776 B.n706 B.n352 50.9715
R1777 B.n706 B.n348 50.9715
R1778 B.n712 B.n348 50.9715
R1779 B.n712 B.n344 50.9715
R1780 B.n718 B.n344 50.9715
R1781 B.n718 B.n340 50.9715
R1782 B.n724 B.n340 50.9715
R1783 B.n730 B.n336 50.9715
R1784 B.n730 B.n332 50.9715
R1785 B.n736 B.n332 50.9715
R1786 B.n736 B.n328 50.9715
R1787 B.n742 B.n328 50.9715
R1788 B.n742 B.n324 50.9715
R1789 B.n748 B.n324 50.9715
R1790 B.n748 B.n320 50.9715
R1791 B.n754 B.n320 50.9715
R1792 B.n754 B.n316 50.9715
R1793 B.n760 B.n316 50.9715
R1794 B.n766 B.n312 50.9715
R1795 B.n766 B.n308 50.9715
R1796 B.n773 B.n308 50.9715
R1797 B.n773 B.n304 50.9715
R1798 B.n779 B.n304 50.9715
R1799 B.n779 B.n4 50.9715
R1800 B.n974 B.n4 50.9715
R1801 B.n974 B.n973 50.9715
R1802 B.n973 B.n972 50.9715
R1803 B.n972 B.n8 50.9715
R1804 B.n12 B.n8 50.9715
R1805 B.n965 B.n12 50.9715
R1806 B.n965 B.n964 50.9715
R1807 B.n964 B.n963 50.9715
R1808 B.n963 B.n16 50.9715
R1809 B.n957 B.n956 50.9715
R1810 B.n956 B.n955 50.9715
R1811 B.n955 B.n23 50.9715
R1812 B.n949 B.n23 50.9715
R1813 B.n949 B.n948 50.9715
R1814 B.n948 B.n947 50.9715
R1815 B.n947 B.n30 50.9715
R1816 B.n941 B.n30 50.9715
R1817 B.n941 B.n940 50.9715
R1818 B.n940 B.n939 50.9715
R1819 B.n939 B.n37 50.9715
R1820 B.n933 B.n932 50.9715
R1821 B.n932 B.n931 50.9715
R1822 B.n931 B.n44 50.9715
R1823 B.n925 B.n44 50.9715
R1824 B.n925 B.n924 50.9715
R1825 B.n924 B.n923 50.9715
R1826 B.n923 B.n51 50.9715
R1827 B.n917 B.n51 50.9715
R1828 B.n917 B.n916 50.9715
R1829 B.n916 B.n915 50.9715
R1830 B.n915 B.n58 50.9715
R1831 B.n909 B.n908 50.9715
R1832 B.n908 B.n907 50.9715
R1833 B.n907 B.n65 50.9715
R1834 B.n901 B.n65 50.9715
R1835 B.n901 B.n900 50.9715
R1836 B.n900 B.n899 50.9715
R1837 B.n899 B.n72 50.9715
R1838 B.n893 B.n72 50.9715
R1839 B.n893 B.n892 50.9715
R1840 B.n892 B.n891 50.9715
R1841 B.n891 B.n79 50.9715
R1842 B.n885 B.n79 50.9715
R1843 B.n885 B.n884 50.9715
R1844 B.n884 B.n883 50.9715
R1845 B.n883 B.n86 50.9715
R1846 B.n877 B.n876 50.9715
R1847 B.n876 B.n875 50.9715
R1848 B.n875 B.n93 50.9715
R1849 B.n869 B.n93 50.9715
R1850 B.n869 B.n868 50.9715
R1851 B.n868 B.n867 50.9715
R1852 B.n867 B.n100 50.9715
R1853 B.n861 B.n100 50.9715
R1854 B.n861 B.n860 50.9715
R1855 B.t4 B.n360 46.4741
R1856 B.t1 B.n58 46.4741
R1857 B.n760 B.t2 37.4792
R1858 B.n957 B.t5 37.4792
R1859 B.n606 B.n410 34.1859
R1860 B.n613 B.n612 34.1859
R1861 B.n857 B.n856 34.1859
R1862 B.n151 B.n102 34.1859
R1863 B.t3 B.n336 29.9835
R1864 B.t0 B.n37 29.9835
R1865 B.n640 B.t7 28.4843
R1866 B.n877 B.t14 28.4843
R1867 B.t7 B.n392 22.4877
R1868 B.t14 B.n86 22.4877
R1869 B.n724 B.t3 20.9886
R1870 B.n933 B.t0 20.9886
R1871 B B.n977 18.0485
R1872 B.t2 B.n312 13.4928
R1873 B.t5 B.n16 13.4928
R1874 B.n618 B.n410 10.6151
R1875 B.n619 B.n618 10.6151
R1876 B.n620 B.n619 10.6151
R1877 B.n620 B.n402 10.6151
R1878 B.n630 B.n402 10.6151
R1879 B.n631 B.n630 10.6151
R1880 B.n632 B.n631 10.6151
R1881 B.n632 B.n394 10.6151
R1882 B.n642 B.n394 10.6151
R1883 B.n643 B.n642 10.6151
R1884 B.n644 B.n643 10.6151
R1885 B.n644 B.n386 10.6151
R1886 B.n654 B.n386 10.6151
R1887 B.n655 B.n654 10.6151
R1888 B.n656 B.n655 10.6151
R1889 B.n656 B.n378 10.6151
R1890 B.n666 B.n378 10.6151
R1891 B.n667 B.n666 10.6151
R1892 B.n668 B.n667 10.6151
R1893 B.n668 B.n370 10.6151
R1894 B.n678 B.n370 10.6151
R1895 B.n679 B.n678 10.6151
R1896 B.n680 B.n679 10.6151
R1897 B.n680 B.n362 10.6151
R1898 B.n690 B.n362 10.6151
R1899 B.n691 B.n690 10.6151
R1900 B.n692 B.n691 10.6151
R1901 B.n692 B.n354 10.6151
R1902 B.n702 B.n354 10.6151
R1903 B.n703 B.n702 10.6151
R1904 B.n704 B.n703 10.6151
R1905 B.n704 B.n346 10.6151
R1906 B.n714 B.n346 10.6151
R1907 B.n715 B.n714 10.6151
R1908 B.n716 B.n715 10.6151
R1909 B.n716 B.n338 10.6151
R1910 B.n726 B.n338 10.6151
R1911 B.n727 B.n726 10.6151
R1912 B.n728 B.n727 10.6151
R1913 B.n728 B.n330 10.6151
R1914 B.n738 B.n330 10.6151
R1915 B.n739 B.n738 10.6151
R1916 B.n740 B.n739 10.6151
R1917 B.n740 B.n322 10.6151
R1918 B.n750 B.n322 10.6151
R1919 B.n751 B.n750 10.6151
R1920 B.n752 B.n751 10.6151
R1921 B.n752 B.n314 10.6151
R1922 B.n762 B.n314 10.6151
R1923 B.n763 B.n762 10.6151
R1924 B.n764 B.n763 10.6151
R1925 B.n764 B.n306 10.6151
R1926 B.n775 B.n306 10.6151
R1927 B.n776 B.n775 10.6151
R1928 B.n777 B.n776 10.6151
R1929 B.n777 B.n0 10.6151
R1930 B.n606 B.n605 10.6151
R1931 B.n605 B.n604 10.6151
R1932 B.n604 B.n603 10.6151
R1933 B.n603 B.n601 10.6151
R1934 B.n601 B.n598 10.6151
R1935 B.n598 B.n597 10.6151
R1936 B.n597 B.n594 10.6151
R1937 B.n594 B.n593 10.6151
R1938 B.n593 B.n590 10.6151
R1939 B.n590 B.n589 10.6151
R1940 B.n589 B.n586 10.6151
R1941 B.n586 B.n585 10.6151
R1942 B.n585 B.n582 10.6151
R1943 B.n582 B.n581 10.6151
R1944 B.n581 B.n578 10.6151
R1945 B.n578 B.n577 10.6151
R1946 B.n577 B.n574 10.6151
R1947 B.n574 B.n573 10.6151
R1948 B.n573 B.n570 10.6151
R1949 B.n570 B.n569 10.6151
R1950 B.n569 B.n566 10.6151
R1951 B.n566 B.n565 10.6151
R1952 B.n565 B.n562 10.6151
R1953 B.n562 B.n561 10.6151
R1954 B.n561 B.n558 10.6151
R1955 B.n558 B.n557 10.6151
R1956 B.n557 B.n554 10.6151
R1957 B.n554 B.n553 10.6151
R1958 B.n553 B.n550 10.6151
R1959 B.n550 B.n549 10.6151
R1960 B.n549 B.n546 10.6151
R1961 B.n546 B.n545 10.6151
R1962 B.n545 B.n542 10.6151
R1963 B.n540 B.n537 10.6151
R1964 B.n537 B.n536 10.6151
R1965 B.n536 B.n533 10.6151
R1966 B.n533 B.n532 10.6151
R1967 B.n532 B.n529 10.6151
R1968 B.n529 B.n528 10.6151
R1969 B.n528 B.n525 10.6151
R1970 B.n525 B.n524 10.6151
R1971 B.n521 B.n520 10.6151
R1972 B.n520 B.n517 10.6151
R1973 B.n517 B.n516 10.6151
R1974 B.n516 B.n513 10.6151
R1975 B.n513 B.n512 10.6151
R1976 B.n512 B.n509 10.6151
R1977 B.n509 B.n508 10.6151
R1978 B.n508 B.n505 10.6151
R1979 B.n505 B.n504 10.6151
R1980 B.n504 B.n501 10.6151
R1981 B.n501 B.n500 10.6151
R1982 B.n500 B.n497 10.6151
R1983 B.n497 B.n496 10.6151
R1984 B.n496 B.n493 10.6151
R1985 B.n493 B.n492 10.6151
R1986 B.n492 B.n489 10.6151
R1987 B.n489 B.n488 10.6151
R1988 B.n488 B.n485 10.6151
R1989 B.n485 B.n484 10.6151
R1990 B.n484 B.n481 10.6151
R1991 B.n481 B.n480 10.6151
R1992 B.n480 B.n477 10.6151
R1993 B.n477 B.n476 10.6151
R1994 B.n476 B.n473 10.6151
R1995 B.n473 B.n472 10.6151
R1996 B.n472 B.n469 10.6151
R1997 B.n469 B.n468 10.6151
R1998 B.n468 B.n465 10.6151
R1999 B.n465 B.n464 10.6151
R2000 B.n464 B.n461 10.6151
R2001 B.n461 B.n460 10.6151
R2002 B.n460 B.n414 10.6151
R2003 B.n612 B.n414 10.6151
R2004 B.n614 B.n613 10.6151
R2005 B.n614 B.n406 10.6151
R2006 B.n624 B.n406 10.6151
R2007 B.n625 B.n624 10.6151
R2008 B.n626 B.n625 10.6151
R2009 B.n626 B.n398 10.6151
R2010 B.n636 B.n398 10.6151
R2011 B.n637 B.n636 10.6151
R2012 B.n638 B.n637 10.6151
R2013 B.n638 B.n390 10.6151
R2014 B.n648 B.n390 10.6151
R2015 B.n649 B.n648 10.6151
R2016 B.n650 B.n649 10.6151
R2017 B.n650 B.n382 10.6151
R2018 B.n660 B.n382 10.6151
R2019 B.n661 B.n660 10.6151
R2020 B.n662 B.n661 10.6151
R2021 B.n662 B.n374 10.6151
R2022 B.n672 B.n374 10.6151
R2023 B.n673 B.n672 10.6151
R2024 B.n674 B.n673 10.6151
R2025 B.n674 B.n366 10.6151
R2026 B.n684 B.n366 10.6151
R2027 B.n685 B.n684 10.6151
R2028 B.n686 B.n685 10.6151
R2029 B.n686 B.n358 10.6151
R2030 B.n696 B.n358 10.6151
R2031 B.n697 B.n696 10.6151
R2032 B.n698 B.n697 10.6151
R2033 B.n698 B.n350 10.6151
R2034 B.n708 B.n350 10.6151
R2035 B.n709 B.n708 10.6151
R2036 B.n710 B.n709 10.6151
R2037 B.n710 B.n342 10.6151
R2038 B.n720 B.n342 10.6151
R2039 B.n721 B.n720 10.6151
R2040 B.n722 B.n721 10.6151
R2041 B.n722 B.n334 10.6151
R2042 B.n732 B.n334 10.6151
R2043 B.n733 B.n732 10.6151
R2044 B.n734 B.n733 10.6151
R2045 B.n734 B.n326 10.6151
R2046 B.n744 B.n326 10.6151
R2047 B.n745 B.n744 10.6151
R2048 B.n746 B.n745 10.6151
R2049 B.n746 B.n318 10.6151
R2050 B.n756 B.n318 10.6151
R2051 B.n757 B.n756 10.6151
R2052 B.n758 B.n757 10.6151
R2053 B.n758 B.n310 10.6151
R2054 B.n768 B.n310 10.6151
R2055 B.n769 B.n768 10.6151
R2056 B.n771 B.n769 10.6151
R2057 B.n771 B.n770 10.6151
R2058 B.n770 B.n302 10.6151
R2059 B.n782 B.n302 10.6151
R2060 B.n783 B.n782 10.6151
R2061 B.n784 B.n783 10.6151
R2062 B.n785 B.n784 10.6151
R2063 B.n786 B.n785 10.6151
R2064 B.n789 B.n786 10.6151
R2065 B.n790 B.n789 10.6151
R2066 B.n791 B.n790 10.6151
R2067 B.n792 B.n791 10.6151
R2068 B.n794 B.n792 10.6151
R2069 B.n795 B.n794 10.6151
R2070 B.n796 B.n795 10.6151
R2071 B.n797 B.n796 10.6151
R2072 B.n799 B.n797 10.6151
R2073 B.n800 B.n799 10.6151
R2074 B.n801 B.n800 10.6151
R2075 B.n802 B.n801 10.6151
R2076 B.n804 B.n802 10.6151
R2077 B.n805 B.n804 10.6151
R2078 B.n806 B.n805 10.6151
R2079 B.n807 B.n806 10.6151
R2080 B.n809 B.n807 10.6151
R2081 B.n810 B.n809 10.6151
R2082 B.n811 B.n810 10.6151
R2083 B.n812 B.n811 10.6151
R2084 B.n814 B.n812 10.6151
R2085 B.n815 B.n814 10.6151
R2086 B.n816 B.n815 10.6151
R2087 B.n817 B.n816 10.6151
R2088 B.n819 B.n817 10.6151
R2089 B.n820 B.n819 10.6151
R2090 B.n821 B.n820 10.6151
R2091 B.n822 B.n821 10.6151
R2092 B.n824 B.n822 10.6151
R2093 B.n825 B.n824 10.6151
R2094 B.n826 B.n825 10.6151
R2095 B.n827 B.n826 10.6151
R2096 B.n829 B.n827 10.6151
R2097 B.n830 B.n829 10.6151
R2098 B.n831 B.n830 10.6151
R2099 B.n832 B.n831 10.6151
R2100 B.n834 B.n832 10.6151
R2101 B.n835 B.n834 10.6151
R2102 B.n836 B.n835 10.6151
R2103 B.n837 B.n836 10.6151
R2104 B.n839 B.n837 10.6151
R2105 B.n840 B.n839 10.6151
R2106 B.n841 B.n840 10.6151
R2107 B.n842 B.n841 10.6151
R2108 B.n844 B.n842 10.6151
R2109 B.n845 B.n844 10.6151
R2110 B.n846 B.n845 10.6151
R2111 B.n847 B.n846 10.6151
R2112 B.n849 B.n847 10.6151
R2113 B.n850 B.n849 10.6151
R2114 B.n851 B.n850 10.6151
R2115 B.n852 B.n851 10.6151
R2116 B.n854 B.n852 10.6151
R2117 B.n855 B.n854 10.6151
R2118 B.n856 B.n855 10.6151
R2119 B.n969 B.n1 10.6151
R2120 B.n969 B.n968 10.6151
R2121 B.n968 B.n967 10.6151
R2122 B.n967 B.n10 10.6151
R2123 B.n961 B.n10 10.6151
R2124 B.n961 B.n960 10.6151
R2125 B.n960 B.n959 10.6151
R2126 B.n959 B.n18 10.6151
R2127 B.n953 B.n18 10.6151
R2128 B.n953 B.n952 10.6151
R2129 B.n952 B.n951 10.6151
R2130 B.n951 B.n25 10.6151
R2131 B.n945 B.n25 10.6151
R2132 B.n945 B.n944 10.6151
R2133 B.n944 B.n943 10.6151
R2134 B.n943 B.n32 10.6151
R2135 B.n937 B.n32 10.6151
R2136 B.n937 B.n936 10.6151
R2137 B.n936 B.n935 10.6151
R2138 B.n935 B.n39 10.6151
R2139 B.n929 B.n39 10.6151
R2140 B.n929 B.n928 10.6151
R2141 B.n928 B.n927 10.6151
R2142 B.n927 B.n46 10.6151
R2143 B.n921 B.n46 10.6151
R2144 B.n921 B.n920 10.6151
R2145 B.n920 B.n919 10.6151
R2146 B.n919 B.n53 10.6151
R2147 B.n913 B.n53 10.6151
R2148 B.n913 B.n912 10.6151
R2149 B.n912 B.n911 10.6151
R2150 B.n911 B.n60 10.6151
R2151 B.n905 B.n60 10.6151
R2152 B.n905 B.n904 10.6151
R2153 B.n904 B.n903 10.6151
R2154 B.n903 B.n67 10.6151
R2155 B.n897 B.n67 10.6151
R2156 B.n897 B.n896 10.6151
R2157 B.n896 B.n895 10.6151
R2158 B.n895 B.n74 10.6151
R2159 B.n889 B.n74 10.6151
R2160 B.n889 B.n888 10.6151
R2161 B.n888 B.n887 10.6151
R2162 B.n887 B.n81 10.6151
R2163 B.n881 B.n81 10.6151
R2164 B.n881 B.n880 10.6151
R2165 B.n880 B.n879 10.6151
R2166 B.n879 B.n88 10.6151
R2167 B.n873 B.n88 10.6151
R2168 B.n873 B.n872 10.6151
R2169 B.n872 B.n871 10.6151
R2170 B.n871 B.n95 10.6151
R2171 B.n865 B.n95 10.6151
R2172 B.n865 B.n864 10.6151
R2173 B.n864 B.n863 10.6151
R2174 B.n863 B.n102 10.6151
R2175 B.n152 B.n151 10.6151
R2176 B.n155 B.n152 10.6151
R2177 B.n156 B.n155 10.6151
R2178 B.n159 B.n156 10.6151
R2179 B.n160 B.n159 10.6151
R2180 B.n163 B.n160 10.6151
R2181 B.n164 B.n163 10.6151
R2182 B.n167 B.n164 10.6151
R2183 B.n168 B.n167 10.6151
R2184 B.n171 B.n168 10.6151
R2185 B.n172 B.n171 10.6151
R2186 B.n175 B.n172 10.6151
R2187 B.n176 B.n175 10.6151
R2188 B.n179 B.n176 10.6151
R2189 B.n180 B.n179 10.6151
R2190 B.n183 B.n180 10.6151
R2191 B.n184 B.n183 10.6151
R2192 B.n187 B.n184 10.6151
R2193 B.n188 B.n187 10.6151
R2194 B.n191 B.n188 10.6151
R2195 B.n192 B.n191 10.6151
R2196 B.n195 B.n192 10.6151
R2197 B.n196 B.n195 10.6151
R2198 B.n199 B.n196 10.6151
R2199 B.n200 B.n199 10.6151
R2200 B.n203 B.n200 10.6151
R2201 B.n204 B.n203 10.6151
R2202 B.n207 B.n204 10.6151
R2203 B.n208 B.n207 10.6151
R2204 B.n211 B.n208 10.6151
R2205 B.n212 B.n211 10.6151
R2206 B.n215 B.n212 10.6151
R2207 B.n216 B.n215 10.6151
R2208 B.n220 B.n219 10.6151
R2209 B.n223 B.n220 10.6151
R2210 B.n224 B.n223 10.6151
R2211 B.n227 B.n224 10.6151
R2212 B.n228 B.n227 10.6151
R2213 B.n231 B.n228 10.6151
R2214 B.n232 B.n231 10.6151
R2215 B.n235 B.n232 10.6151
R2216 B.n240 B.n237 10.6151
R2217 B.n241 B.n240 10.6151
R2218 B.n244 B.n241 10.6151
R2219 B.n245 B.n244 10.6151
R2220 B.n248 B.n245 10.6151
R2221 B.n249 B.n248 10.6151
R2222 B.n252 B.n249 10.6151
R2223 B.n253 B.n252 10.6151
R2224 B.n256 B.n253 10.6151
R2225 B.n257 B.n256 10.6151
R2226 B.n260 B.n257 10.6151
R2227 B.n261 B.n260 10.6151
R2228 B.n264 B.n261 10.6151
R2229 B.n265 B.n264 10.6151
R2230 B.n268 B.n265 10.6151
R2231 B.n269 B.n268 10.6151
R2232 B.n272 B.n269 10.6151
R2233 B.n273 B.n272 10.6151
R2234 B.n276 B.n273 10.6151
R2235 B.n277 B.n276 10.6151
R2236 B.n280 B.n277 10.6151
R2237 B.n281 B.n280 10.6151
R2238 B.n284 B.n281 10.6151
R2239 B.n285 B.n284 10.6151
R2240 B.n288 B.n285 10.6151
R2241 B.n289 B.n288 10.6151
R2242 B.n292 B.n289 10.6151
R2243 B.n293 B.n292 10.6151
R2244 B.n296 B.n293 10.6151
R2245 B.n297 B.n296 10.6151
R2246 B.n300 B.n297 10.6151
R2247 B.n301 B.n300 10.6151
R2248 B.n857 B.n301 10.6151
R2249 B.n977 B.n0 8.11757
R2250 B.n977 B.n1 8.11757
R2251 B.n541 B.n540 6.5566
R2252 B.n524 B.n458 6.5566
R2253 B.n219 B.n149 6.5566
R2254 B.n236 B.n235 6.5566
R2255 B.n688 B.t4 4.49794
R2256 B.n909 B.t1 4.49794
R2257 B.n542 B.n541 4.05904
R2258 B.n521 B.n458 4.05904
R2259 B.n216 B.n149 4.05904
R2260 B.n237 B.n236 4.05904
R2261 VN.n37 VN.n20 161.3
R2262 VN.n36 VN.n35 161.3
R2263 VN.n34 VN.n21 161.3
R2264 VN.n33 VN.n32 161.3
R2265 VN.n31 VN.n22 161.3
R2266 VN.n30 VN.n29 161.3
R2267 VN.n28 VN.n23 161.3
R2268 VN.n27 VN.n26 161.3
R2269 VN.n17 VN.n0 161.3
R2270 VN.n16 VN.n15 161.3
R2271 VN.n14 VN.n1 161.3
R2272 VN.n13 VN.n12 161.3
R2273 VN.n11 VN.n2 161.3
R2274 VN.n10 VN.n9 161.3
R2275 VN.n8 VN.n3 161.3
R2276 VN.n7 VN.n6 161.3
R2277 VN.n4 VN.t4 90.8179
R2278 VN.n24 VN.t2 90.8179
R2279 VN.n5 VN.n4 62.6969
R2280 VN.n25 VN.n24 62.6969
R2281 VN.n19 VN.n18 60.5633
R2282 VN.n39 VN.n38 60.5633
R2283 VN.n5 VN.t1 58.6896
R2284 VN.n18 VN.t3 58.6896
R2285 VN.n25 VN.t5 58.6896
R2286 VN.n38 VN.t0 58.6896
R2287 VN.n12 VN.n11 55.5035
R2288 VN.n32 VN.n31 55.5035
R2289 VN VN.n39 51.9168
R2290 VN.n12 VN.n1 25.3177
R2291 VN.n32 VN.n21 25.3177
R2292 VN.n6 VN.n3 24.3439
R2293 VN.n10 VN.n3 24.3439
R2294 VN.n11 VN.n10 24.3439
R2295 VN.n16 VN.n1 24.3439
R2296 VN.n17 VN.n16 24.3439
R2297 VN.n31 VN.n30 24.3439
R2298 VN.n30 VN.n23 24.3439
R2299 VN.n26 VN.n23 24.3439
R2300 VN.n37 VN.n36 24.3439
R2301 VN.n36 VN.n21 24.3439
R2302 VN.n18 VN.n17 21.4227
R2303 VN.n38 VN.n37 21.4227
R2304 VN.n6 VN.n5 12.1722
R2305 VN.n26 VN.n25 12.1722
R2306 VN.n27 VN.n24 2.65074
R2307 VN.n7 VN.n4 2.65074
R2308 VN.n39 VN.n20 0.417764
R2309 VN.n19 VN.n0 0.417764
R2310 VN VN.n19 0.394061
R2311 VN.n35 VN.n20 0.189894
R2312 VN.n35 VN.n34 0.189894
R2313 VN.n34 VN.n33 0.189894
R2314 VN.n33 VN.n22 0.189894
R2315 VN.n29 VN.n22 0.189894
R2316 VN.n29 VN.n28 0.189894
R2317 VN.n28 VN.n27 0.189894
R2318 VN.n8 VN.n7 0.189894
R2319 VN.n9 VN.n8 0.189894
R2320 VN.n9 VN.n2 0.189894
R2321 VN.n13 VN.n2 0.189894
R2322 VN.n14 VN.n13 0.189894
R2323 VN.n15 VN.n14 0.189894
R2324 VN.n15 VN.n0 0.189894
R2325 VDD2.n95 VDD2.n51 289.615
R2326 VDD2.n44 VDD2.n0 289.615
R2327 VDD2.n96 VDD2.n95 185
R2328 VDD2.n94 VDD2.n93 185
R2329 VDD2.n55 VDD2.n54 185
R2330 VDD2.n59 VDD2.n57 185
R2331 VDD2.n88 VDD2.n87 185
R2332 VDD2.n86 VDD2.n85 185
R2333 VDD2.n61 VDD2.n60 185
R2334 VDD2.n80 VDD2.n79 185
R2335 VDD2.n78 VDD2.n77 185
R2336 VDD2.n65 VDD2.n64 185
R2337 VDD2.n72 VDD2.n71 185
R2338 VDD2.n70 VDD2.n69 185
R2339 VDD2.n17 VDD2.n16 185
R2340 VDD2.n19 VDD2.n18 185
R2341 VDD2.n12 VDD2.n11 185
R2342 VDD2.n25 VDD2.n24 185
R2343 VDD2.n27 VDD2.n26 185
R2344 VDD2.n8 VDD2.n7 185
R2345 VDD2.n34 VDD2.n33 185
R2346 VDD2.n35 VDD2.n6 185
R2347 VDD2.n37 VDD2.n36 185
R2348 VDD2.n4 VDD2.n3 185
R2349 VDD2.n43 VDD2.n42 185
R2350 VDD2.n45 VDD2.n44 185
R2351 VDD2.n68 VDD2.t5 149.524
R2352 VDD2.n15 VDD2.t1 149.524
R2353 VDD2.n95 VDD2.n94 104.615
R2354 VDD2.n94 VDD2.n54 104.615
R2355 VDD2.n59 VDD2.n54 104.615
R2356 VDD2.n87 VDD2.n59 104.615
R2357 VDD2.n87 VDD2.n86 104.615
R2358 VDD2.n86 VDD2.n60 104.615
R2359 VDD2.n79 VDD2.n60 104.615
R2360 VDD2.n79 VDD2.n78 104.615
R2361 VDD2.n78 VDD2.n64 104.615
R2362 VDD2.n71 VDD2.n64 104.615
R2363 VDD2.n71 VDD2.n70 104.615
R2364 VDD2.n18 VDD2.n17 104.615
R2365 VDD2.n18 VDD2.n11 104.615
R2366 VDD2.n25 VDD2.n11 104.615
R2367 VDD2.n26 VDD2.n25 104.615
R2368 VDD2.n26 VDD2.n7 104.615
R2369 VDD2.n34 VDD2.n7 104.615
R2370 VDD2.n35 VDD2.n34 104.615
R2371 VDD2.n36 VDD2.n35 104.615
R2372 VDD2.n36 VDD2.n3 104.615
R2373 VDD2.n43 VDD2.n3 104.615
R2374 VDD2.n44 VDD2.n43 104.615
R2375 VDD2.n50 VDD2.n49 66.9526
R2376 VDD2 VDD2.n101 66.9497
R2377 VDD2.n50 VDD2.n48 54.6209
R2378 VDD2.n70 VDD2.t5 52.3082
R2379 VDD2.n17 VDD2.t1 52.3082
R2380 VDD2.n100 VDD2.n99 51.9672
R2381 VDD2.n100 VDD2.n50 43.558
R2382 VDD2.n57 VDD2.n55 13.1884
R2383 VDD2.n37 VDD2.n4 13.1884
R2384 VDD2.n93 VDD2.n92 12.8005
R2385 VDD2.n89 VDD2.n88 12.8005
R2386 VDD2.n38 VDD2.n6 12.8005
R2387 VDD2.n42 VDD2.n41 12.8005
R2388 VDD2.n96 VDD2.n53 12.0247
R2389 VDD2.n85 VDD2.n58 12.0247
R2390 VDD2.n33 VDD2.n32 12.0247
R2391 VDD2.n45 VDD2.n2 12.0247
R2392 VDD2.n97 VDD2.n51 11.249
R2393 VDD2.n84 VDD2.n61 11.249
R2394 VDD2.n31 VDD2.n8 11.249
R2395 VDD2.n46 VDD2.n0 11.249
R2396 VDD2.n81 VDD2.n80 10.4732
R2397 VDD2.n28 VDD2.n27 10.4732
R2398 VDD2.n69 VDD2.n68 10.2747
R2399 VDD2.n16 VDD2.n15 10.2747
R2400 VDD2.n77 VDD2.n63 9.69747
R2401 VDD2.n24 VDD2.n10 9.69747
R2402 VDD2.n99 VDD2.n98 9.45567
R2403 VDD2.n48 VDD2.n47 9.45567
R2404 VDD2.n67 VDD2.n66 9.3005
R2405 VDD2.n74 VDD2.n73 9.3005
R2406 VDD2.n76 VDD2.n75 9.3005
R2407 VDD2.n63 VDD2.n62 9.3005
R2408 VDD2.n82 VDD2.n81 9.3005
R2409 VDD2.n84 VDD2.n83 9.3005
R2410 VDD2.n58 VDD2.n56 9.3005
R2411 VDD2.n90 VDD2.n89 9.3005
R2412 VDD2.n98 VDD2.n97 9.3005
R2413 VDD2.n53 VDD2.n52 9.3005
R2414 VDD2.n92 VDD2.n91 9.3005
R2415 VDD2.n47 VDD2.n46 9.3005
R2416 VDD2.n2 VDD2.n1 9.3005
R2417 VDD2.n41 VDD2.n40 9.3005
R2418 VDD2.n14 VDD2.n13 9.3005
R2419 VDD2.n21 VDD2.n20 9.3005
R2420 VDD2.n23 VDD2.n22 9.3005
R2421 VDD2.n10 VDD2.n9 9.3005
R2422 VDD2.n29 VDD2.n28 9.3005
R2423 VDD2.n31 VDD2.n30 9.3005
R2424 VDD2.n32 VDD2.n5 9.3005
R2425 VDD2.n39 VDD2.n38 9.3005
R2426 VDD2.n76 VDD2.n65 8.92171
R2427 VDD2.n23 VDD2.n12 8.92171
R2428 VDD2.n73 VDD2.n72 8.14595
R2429 VDD2.n20 VDD2.n19 8.14595
R2430 VDD2.n69 VDD2.n67 7.3702
R2431 VDD2.n16 VDD2.n14 7.3702
R2432 VDD2.n72 VDD2.n67 5.81868
R2433 VDD2.n19 VDD2.n14 5.81868
R2434 VDD2.n73 VDD2.n65 5.04292
R2435 VDD2.n20 VDD2.n12 5.04292
R2436 VDD2.n77 VDD2.n76 4.26717
R2437 VDD2.n24 VDD2.n23 4.26717
R2438 VDD2.n80 VDD2.n63 3.49141
R2439 VDD2.n27 VDD2.n10 3.49141
R2440 VDD2.n68 VDD2.n66 2.84303
R2441 VDD2.n15 VDD2.n13 2.84303
R2442 VDD2 VDD2.n100 2.76774
R2443 VDD2.n99 VDD2.n51 2.71565
R2444 VDD2.n81 VDD2.n61 2.71565
R2445 VDD2.n28 VDD2.n8 2.71565
R2446 VDD2.n48 VDD2.n0 2.71565
R2447 VDD2.n101 VDD2.t0 2.10688
R2448 VDD2.n101 VDD2.t3 2.10688
R2449 VDD2.n49 VDD2.t4 2.10688
R2450 VDD2.n49 VDD2.t2 2.10688
R2451 VDD2.n97 VDD2.n96 1.93989
R2452 VDD2.n85 VDD2.n84 1.93989
R2453 VDD2.n33 VDD2.n31 1.93989
R2454 VDD2.n46 VDD2.n45 1.93989
R2455 VDD2.n93 VDD2.n53 1.16414
R2456 VDD2.n88 VDD2.n58 1.16414
R2457 VDD2.n32 VDD2.n6 1.16414
R2458 VDD2.n42 VDD2.n2 1.16414
R2459 VDD2.n92 VDD2.n55 0.388379
R2460 VDD2.n89 VDD2.n57 0.388379
R2461 VDD2.n38 VDD2.n37 0.388379
R2462 VDD2.n41 VDD2.n4 0.388379
R2463 VDD2.n98 VDD2.n52 0.155672
R2464 VDD2.n91 VDD2.n52 0.155672
R2465 VDD2.n91 VDD2.n90 0.155672
R2466 VDD2.n90 VDD2.n56 0.155672
R2467 VDD2.n83 VDD2.n56 0.155672
R2468 VDD2.n83 VDD2.n82 0.155672
R2469 VDD2.n82 VDD2.n62 0.155672
R2470 VDD2.n75 VDD2.n62 0.155672
R2471 VDD2.n75 VDD2.n74 0.155672
R2472 VDD2.n74 VDD2.n66 0.155672
R2473 VDD2.n21 VDD2.n13 0.155672
R2474 VDD2.n22 VDD2.n21 0.155672
R2475 VDD2.n22 VDD2.n9 0.155672
R2476 VDD2.n29 VDD2.n9 0.155672
R2477 VDD2.n30 VDD2.n29 0.155672
R2478 VDD2.n30 VDD2.n5 0.155672
R2479 VDD2.n39 VDD2.n5 0.155672
R2480 VDD2.n40 VDD2.n39 0.155672
R2481 VDD2.n40 VDD2.n1 0.155672
R2482 VDD2.n47 VDD2.n1 0.155672
C0 VDD1 VDD2 1.89903f
C1 VTAIL VDD2 7.429911f
C2 VDD2 VP 0.564295f
C3 VTAIL VDD1 7.36923f
C4 VDD2 VN 5.6953f
C5 VDD1 VP 6.10515f
C6 VDD1 VN 0.152202f
C7 VTAIL VP 6.29791f
C8 VTAIL VN 6.28323f
C9 VP VN 7.680161f
C10 VDD2 B 6.489043f
C11 VDD1 B 6.687339f
C12 VTAIL B 7.552317f
C13 VN B 16.447f
C14 VP B 15.179312f
C15 VDD2.n0 B 0.0302f
C16 VDD2.n1 B 0.021485f
C17 VDD2.n2 B 0.011545f
C18 VDD2.n3 B 0.027289f
C19 VDD2.n4 B 0.011885f
C20 VDD2.n5 B 0.021485f
C21 VDD2.n6 B 0.012224f
C22 VDD2.n7 B 0.027289f
C23 VDD2.n8 B 0.012224f
C24 VDD2.n9 B 0.021485f
C25 VDD2.n10 B 0.011545f
C26 VDD2.n11 B 0.027289f
C27 VDD2.n12 B 0.012224f
C28 VDD2.n13 B 0.835423f
C29 VDD2.n14 B 0.011545f
C30 VDD2.t1 B 0.045793f
C31 VDD2.n15 B 0.133468f
C32 VDD2.n16 B 0.019291f
C33 VDD2.n17 B 0.020467f
C34 VDD2.n18 B 0.027289f
C35 VDD2.n19 B 0.012224f
C36 VDD2.n20 B 0.011545f
C37 VDD2.n21 B 0.021485f
C38 VDD2.n22 B 0.021485f
C39 VDD2.n23 B 0.011545f
C40 VDD2.n24 B 0.012224f
C41 VDD2.n25 B 0.027289f
C42 VDD2.n26 B 0.027289f
C43 VDD2.n27 B 0.012224f
C44 VDD2.n28 B 0.011545f
C45 VDD2.n29 B 0.021485f
C46 VDD2.n30 B 0.021485f
C47 VDD2.n31 B 0.011545f
C48 VDD2.n32 B 0.011545f
C49 VDD2.n33 B 0.012224f
C50 VDD2.n34 B 0.027289f
C51 VDD2.n35 B 0.027289f
C52 VDD2.n36 B 0.027289f
C53 VDD2.n37 B 0.011885f
C54 VDD2.n38 B 0.011545f
C55 VDD2.n39 B 0.021485f
C56 VDD2.n40 B 0.021485f
C57 VDD2.n41 B 0.011545f
C58 VDD2.n42 B 0.012224f
C59 VDD2.n43 B 0.027289f
C60 VDD2.n44 B 0.059076f
C61 VDD2.n45 B 0.012224f
C62 VDD2.n46 B 0.011545f
C63 VDD2.n47 B 0.054359f
C64 VDD2.n48 B 0.059071f
C65 VDD2.t4 B 0.159597f
C66 VDD2.t2 B 0.159597f
C67 VDD2.n49 B 1.4072f
C68 VDD2.n50 B 2.62888f
C69 VDD2.n51 B 0.0302f
C70 VDD2.n52 B 0.021485f
C71 VDD2.n53 B 0.011545f
C72 VDD2.n54 B 0.027289f
C73 VDD2.n55 B 0.011885f
C74 VDD2.n56 B 0.021485f
C75 VDD2.n57 B 0.011885f
C76 VDD2.n58 B 0.011545f
C77 VDD2.n59 B 0.027289f
C78 VDD2.n60 B 0.027289f
C79 VDD2.n61 B 0.012224f
C80 VDD2.n62 B 0.021485f
C81 VDD2.n63 B 0.011545f
C82 VDD2.n64 B 0.027289f
C83 VDD2.n65 B 0.012224f
C84 VDD2.n66 B 0.835423f
C85 VDD2.n67 B 0.011545f
C86 VDD2.t5 B 0.045793f
C87 VDD2.n68 B 0.133468f
C88 VDD2.n69 B 0.019291f
C89 VDD2.n70 B 0.020467f
C90 VDD2.n71 B 0.027289f
C91 VDD2.n72 B 0.012224f
C92 VDD2.n73 B 0.011545f
C93 VDD2.n74 B 0.021485f
C94 VDD2.n75 B 0.021485f
C95 VDD2.n76 B 0.011545f
C96 VDD2.n77 B 0.012224f
C97 VDD2.n78 B 0.027289f
C98 VDD2.n79 B 0.027289f
C99 VDD2.n80 B 0.012224f
C100 VDD2.n81 B 0.011545f
C101 VDD2.n82 B 0.021485f
C102 VDD2.n83 B 0.021485f
C103 VDD2.n84 B 0.011545f
C104 VDD2.n85 B 0.012224f
C105 VDD2.n86 B 0.027289f
C106 VDD2.n87 B 0.027289f
C107 VDD2.n88 B 0.012224f
C108 VDD2.n89 B 0.011545f
C109 VDD2.n90 B 0.021485f
C110 VDD2.n91 B 0.021485f
C111 VDD2.n92 B 0.011545f
C112 VDD2.n93 B 0.012224f
C113 VDD2.n94 B 0.027289f
C114 VDD2.n95 B 0.059076f
C115 VDD2.n96 B 0.012224f
C116 VDD2.n97 B 0.011545f
C117 VDD2.n98 B 0.054359f
C118 VDD2.n99 B 0.047996f
C119 VDD2.n100 B 2.32768f
C120 VDD2.t0 B 0.159597f
C121 VDD2.t3 B 0.159597f
C122 VDD2.n101 B 1.40717f
C123 VN.n0 B 0.035596f
C124 VN.t3 B 1.8555f
C125 VN.n1 B 0.036082f
C126 VN.n2 B 0.018918f
C127 VN.n3 B 0.035436f
C128 VN.t4 B 2.14134f
C129 VN.n4 B 0.696023f
C130 VN.t1 B 1.8555f
C131 VN.n5 B 0.727492f
C132 VN.n6 B 0.026688f
C133 VN.n7 B 0.248841f
C134 VN.n8 B 0.018918f
C135 VN.n9 B 0.018918f
C136 VN.n10 B 0.035436f
C137 VN.n11 B 0.032686f
C138 VN.n12 B 0.022144f
C139 VN.n13 B 0.018918f
C140 VN.n14 B 0.018918f
C141 VN.n15 B 0.018918f
C142 VN.n16 B 0.035436f
C143 VN.n17 B 0.033336f
C144 VN.n18 B 0.742196f
C145 VN.n19 B 0.058061f
C146 VN.n20 B 0.035596f
C147 VN.t0 B 1.8555f
C148 VN.n21 B 0.036082f
C149 VN.n22 B 0.018918f
C150 VN.n23 B 0.035436f
C151 VN.t2 B 2.14134f
C152 VN.n24 B 0.696023f
C153 VN.t5 B 1.8555f
C154 VN.n25 B 0.727492f
C155 VN.n26 B 0.026688f
C156 VN.n27 B 0.248841f
C157 VN.n28 B 0.018918f
C158 VN.n29 B 0.018918f
C159 VN.n30 B 0.035436f
C160 VN.n31 B 0.032686f
C161 VN.n32 B 0.022144f
C162 VN.n33 B 0.018918f
C163 VN.n34 B 0.018918f
C164 VN.n35 B 0.018918f
C165 VN.n36 B 0.035436f
C166 VN.n37 B 0.033336f
C167 VN.n38 B 0.742196f
C168 VN.n39 B 1.16174f
C169 VDD1.n0 B 0.030934f
C170 VDD1.n1 B 0.022008f
C171 VDD1.n2 B 0.011826f
C172 VDD1.n3 B 0.027953f
C173 VDD1.n4 B 0.012174f
C174 VDD1.n5 B 0.022008f
C175 VDD1.n6 B 0.012174f
C176 VDD1.n7 B 0.011826f
C177 VDD1.n8 B 0.027953f
C178 VDD1.n9 B 0.027953f
C179 VDD1.n10 B 0.012522f
C180 VDD1.n11 B 0.022008f
C181 VDD1.n12 B 0.011826f
C182 VDD1.n13 B 0.027953f
C183 VDD1.n14 B 0.012522f
C184 VDD1.n15 B 0.855748f
C185 VDD1.n16 B 0.011826f
C186 VDD1.t4 B 0.046907f
C187 VDD1.n17 B 0.136715f
C188 VDD1.n18 B 0.01976f
C189 VDD1.n19 B 0.020965f
C190 VDD1.n20 B 0.027953f
C191 VDD1.n21 B 0.012522f
C192 VDD1.n22 B 0.011826f
C193 VDD1.n23 B 0.022008f
C194 VDD1.n24 B 0.022008f
C195 VDD1.n25 B 0.011826f
C196 VDD1.n26 B 0.012522f
C197 VDD1.n27 B 0.027953f
C198 VDD1.n28 B 0.027953f
C199 VDD1.n29 B 0.012522f
C200 VDD1.n30 B 0.011826f
C201 VDD1.n31 B 0.022008f
C202 VDD1.n32 B 0.022008f
C203 VDD1.n33 B 0.011826f
C204 VDD1.n34 B 0.012522f
C205 VDD1.n35 B 0.027953f
C206 VDD1.n36 B 0.027953f
C207 VDD1.n37 B 0.012522f
C208 VDD1.n38 B 0.011826f
C209 VDD1.n39 B 0.022008f
C210 VDD1.n40 B 0.022008f
C211 VDD1.n41 B 0.011826f
C212 VDD1.n42 B 0.012522f
C213 VDD1.n43 B 0.027953f
C214 VDD1.n44 B 0.060513f
C215 VDD1.n45 B 0.012522f
C216 VDD1.n46 B 0.011826f
C217 VDD1.n47 B 0.055681f
C218 VDD1.n48 B 0.061367f
C219 VDD1.n49 B 0.030934f
C220 VDD1.n50 B 0.022008f
C221 VDD1.n51 B 0.011826f
C222 VDD1.n52 B 0.027953f
C223 VDD1.n53 B 0.012174f
C224 VDD1.n54 B 0.022008f
C225 VDD1.n55 B 0.012522f
C226 VDD1.n56 B 0.027953f
C227 VDD1.n57 B 0.012522f
C228 VDD1.n58 B 0.022008f
C229 VDD1.n59 B 0.011826f
C230 VDD1.n60 B 0.027953f
C231 VDD1.n61 B 0.012522f
C232 VDD1.n62 B 0.855748f
C233 VDD1.n63 B 0.011826f
C234 VDD1.t3 B 0.046907f
C235 VDD1.n64 B 0.136715f
C236 VDD1.n65 B 0.01976f
C237 VDD1.n66 B 0.020965f
C238 VDD1.n67 B 0.027953f
C239 VDD1.n68 B 0.012522f
C240 VDD1.n69 B 0.011826f
C241 VDD1.n70 B 0.022008f
C242 VDD1.n71 B 0.022008f
C243 VDD1.n72 B 0.011826f
C244 VDD1.n73 B 0.012522f
C245 VDD1.n74 B 0.027953f
C246 VDD1.n75 B 0.027953f
C247 VDD1.n76 B 0.012522f
C248 VDD1.n77 B 0.011826f
C249 VDD1.n78 B 0.022008f
C250 VDD1.n79 B 0.022008f
C251 VDD1.n80 B 0.011826f
C252 VDD1.n81 B 0.011826f
C253 VDD1.n82 B 0.012522f
C254 VDD1.n83 B 0.027953f
C255 VDD1.n84 B 0.027953f
C256 VDD1.n85 B 0.027953f
C257 VDD1.n86 B 0.012174f
C258 VDD1.n87 B 0.011826f
C259 VDD1.n88 B 0.022008f
C260 VDD1.n89 B 0.022008f
C261 VDD1.n90 B 0.011826f
C262 VDD1.n91 B 0.012522f
C263 VDD1.n92 B 0.027953f
C264 VDD1.n93 B 0.060513f
C265 VDD1.n94 B 0.012522f
C266 VDD1.n95 B 0.011826f
C267 VDD1.n96 B 0.055681f
C268 VDD1.n97 B 0.060509f
C269 VDD1.t0 B 0.16348f
C270 VDD1.t5 B 0.16348f
C271 VDD1.n98 B 1.44144f
C272 VDD1.n99 B 2.82945f
C273 VDD1.t2 B 0.16348f
C274 VDD1.t1 B 0.16348f
C275 VDD1.n100 B 1.43508f
C276 VDD1.n101 B 2.589f
C277 VTAIL.t5 B 0.190851f
C278 VTAIL.t0 B 0.190851f
C279 VTAIL.n0 B 1.60749f
C280 VTAIL.n1 B 0.506934f
C281 VTAIL.n2 B 0.036114f
C282 VTAIL.n3 B 0.025693f
C283 VTAIL.n4 B 0.013806f
C284 VTAIL.n5 B 0.032633f
C285 VTAIL.n6 B 0.014212f
C286 VTAIL.n7 B 0.025693f
C287 VTAIL.n8 B 0.014618f
C288 VTAIL.n9 B 0.032633f
C289 VTAIL.n10 B 0.014618f
C290 VTAIL.n11 B 0.025693f
C291 VTAIL.n12 B 0.013806f
C292 VTAIL.n13 B 0.032633f
C293 VTAIL.n14 B 0.014618f
C294 VTAIL.n15 B 0.999026f
C295 VTAIL.n16 B 0.013806f
C296 VTAIL.t11 B 0.05476f
C297 VTAIL.n17 B 0.159606f
C298 VTAIL.n18 B 0.023069f
C299 VTAIL.n19 B 0.024475f
C300 VTAIL.n20 B 0.032633f
C301 VTAIL.n21 B 0.014618f
C302 VTAIL.n22 B 0.013806f
C303 VTAIL.n23 B 0.025693f
C304 VTAIL.n24 B 0.025693f
C305 VTAIL.n25 B 0.013806f
C306 VTAIL.n26 B 0.014618f
C307 VTAIL.n27 B 0.032633f
C308 VTAIL.n28 B 0.032633f
C309 VTAIL.n29 B 0.014618f
C310 VTAIL.n30 B 0.013806f
C311 VTAIL.n31 B 0.025693f
C312 VTAIL.n32 B 0.025693f
C313 VTAIL.n33 B 0.013806f
C314 VTAIL.n34 B 0.013806f
C315 VTAIL.n35 B 0.014618f
C316 VTAIL.n36 B 0.032633f
C317 VTAIL.n37 B 0.032633f
C318 VTAIL.n38 B 0.032633f
C319 VTAIL.n39 B 0.014212f
C320 VTAIL.n40 B 0.013806f
C321 VTAIL.n41 B 0.025693f
C322 VTAIL.n42 B 0.025693f
C323 VTAIL.n43 B 0.013806f
C324 VTAIL.n44 B 0.014618f
C325 VTAIL.n45 B 0.032633f
C326 VTAIL.n46 B 0.070645f
C327 VTAIL.n47 B 0.014618f
C328 VTAIL.n48 B 0.013806f
C329 VTAIL.n49 B 0.065004f
C330 VTAIL.n50 B 0.039694f
C331 VTAIL.n51 B 0.512572f
C332 VTAIL.t10 B 0.190851f
C333 VTAIL.t7 B 0.190851f
C334 VTAIL.n52 B 1.60749f
C335 VTAIL.n53 B 2.15593f
C336 VTAIL.t4 B 0.190851f
C337 VTAIL.t3 B 0.190851f
C338 VTAIL.n54 B 1.6075f
C339 VTAIL.n55 B 2.15592f
C340 VTAIL.n56 B 0.036114f
C341 VTAIL.n57 B 0.025693f
C342 VTAIL.n58 B 0.013806f
C343 VTAIL.n59 B 0.032633f
C344 VTAIL.n60 B 0.014212f
C345 VTAIL.n61 B 0.025693f
C346 VTAIL.n62 B 0.014212f
C347 VTAIL.n63 B 0.013806f
C348 VTAIL.n64 B 0.032633f
C349 VTAIL.n65 B 0.032633f
C350 VTAIL.n66 B 0.014618f
C351 VTAIL.n67 B 0.025693f
C352 VTAIL.n68 B 0.013806f
C353 VTAIL.n69 B 0.032633f
C354 VTAIL.n70 B 0.014618f
C355 VTAIL.n71 B 0.999026f
C356 VTAIL.n72 B 0.013806f
C357 VTAIL.t2 B 0.05476f
C358 VTAIL.n73 B 0.159606f
C359 VTAIL.n74 B 0.023069f
C360 VTAIL.n75 B 0.024475f
C361 VTAIL.n76 B 0.032633f
C362 VTAIL.n77 B 0.014618f
C363 VTAIL.n78 B 0.013806f
C364 VTAIL.n79 B 0.025693f
C365 VTAIL.n80 B 0.025693f
C366 VTAIL.n81 B 0.013806f
C367 VTAIL.n82 B 0.014618f
C368 VTAIL.n83 B 0.032633f
C369 VTAIL.n84 B 0.032633f
C370 VTAIL.n85 B 0.014618f
C371 VTAIL.n86 B 0.013806f
C372 VTAIL.n87 B 0.025693f
C373 VTAIL.n88 B 0.025693f
C374 VTAIL.n89 B 0.013806f
C375 VTAIL.n90 B 0.014618f
C376 VTAIL.n91 B 0.032633f
C377 VTAIL.n92 B 0.032633f
C378 VTAIL.n93 B 0.014618f
C379 VTAIL.n94 B 0.013806f
C380 VTAIL.n95 B 0.025693f
C381 VTAIL.n96 B 0.025693f
C382 VTAIL.n97 B 0.013806f
C383 VTAIL.n98 B 0.014618f
C384 VTAIL.n99 B 0.032633f
C385 VTAIL.n100 B 0.070645f
C386 VTAIL.n101 B 0.014618f
C387 VTAIL.n102 B 0.013806f
C388 VTAIL.n103 B 0.065004f
C389 VTAIL.n104 B 0.039694f
C390 VTAIL.n105 B 0.512572f
C391 VTAIL.t9 B 0.190851f
C392 VTAIL.t6 B 0.190851f
C393 VTAIL.n106 B 1.6075f
C394 VTAIL.n107 B 0.726385f
C395 VTAIL.n108 B 0.036114f
C396 VTAIL.n109 B 0.025693f
C397 VTAIL.n110 B 0.013806f
C398 VTAIL.n111 B 0.032633f
C399 VTAIL.n112 B 0.014212f
C400 VTAIL.n113 B 0.025693f
C401 VTAIL.n114 B 0.014212f
C402 VTAIL.n115 B 0.013806f
C403 VTAIL.n116 B 0.032633f
C404 VTAIL.n117 B 0.032633f
C405 VTAIL.n118 B 0.014618f
C406 VTAIL.n119 B 0.025693f
C407 VTAIL.n120 B 0.013806f
C408 VTAIL.n121 B 0.032633f
C409 VTAIL.n122 B 0.014618f
C410 VTAIL.n123 B 0.999026f
C411 VTAIL.n124 B 0.013806f
C412 VTAIL.t8 B 0.05476f
C413 VTAIL.n125 B 0.159606f
C414 VTAIL.n126 B 0.023069f
C415 VTAIL.n127 B 0.024475f
C416 VTAIL.n128 B 0.032633f
C417 VTAIL.n129 B 0.014618f
C418 VTAIL.n130 B 0.013806f
C419 VTAIL.n131 B 0.025693f
C420 VTAIL.n132 B 0.025693f
C421 VTAIL.n133 B 0.013806f
C422 VTAIL.n134 B 0.014618f
C423 VTAIL.n135 B 0.032633f
C424 VTAIL.n136 B 0.032633f
C425 VTAIL.n137 B 0.014618f
C426 VTAIL.n138 B 0.013806f
C427 VTAIL.n139 B 0.025693f
C428 VTAIL.n140 B 0.025693f
C429 VTAIL.n141 B 0.013806f
C430 VTAIL.n142 B 0.014618f
C431 VTAIL.n143 B 0.032633f
C432 VTAIL.n144 B 0.032633f
C433 VTAIL.n145 B 0.014618f
C434 VTAIL.n146 B 0.013806f
C435 VTAIL.n147 B 0.025693f
C436 VTAIL.n148 B 0.025693f
C437 VTAIL.n149 B 0.013806f
C438 VTAIL.n150 B 0.014618f
C439 VTAIL.n151 B 0.032633f
C440 VTAIL.n152 B 0.070645f
C441 VTAIL.n153 B 0.014618f
C442 VTAIL.n154 B 0.013806f
C443 VTAIL.n155 B 0.065004f
C444 VTAIL.n156 B 0.039694f
C445 VTAIL.n157 B 1.64307f
C446 VTAIL.n158 B 0.036114f
C447 VTAIL.n159 B 0.025693f
C448 VTAIL.n160 B 0.013806f
C449 VTAIL.n161 B 0.032633f
C450 VTAIL.n162 B 0.014212f
C451 VTAIL.n163 B 0.025693f
C452 VTAIL.n164 B 0.014618f
C453 VTAIL.n165 B 0.032633f
C454 VTAIL.n166 B 0.014618f
C455 VTAIL.n167 B 0.025693f
C456 VTAIL.n168 B 0.013806f
C457 VTAIL.n169 B 0.032633f
C458 VTAIL.n170 B 0.014618f
C459 VTAIL.n171 B 0.999026f
C460 VTAIL.n172 B 0.013806f
C461 VTAIL.t1 B 0.05476f
C462 VTAIL.n173 B 0.159606f
C463 VTAIL.n174 B 0.023069f
C464 VTAIL.n175 B 0.024475f
C465 VTAIL.n176 B 0.032633f
C466 VTAIL.n177 B 0.014618f
C467 VTAIL.n178 B 0.013806f
C468 VTAIL.n179 B 0.025693f
C469 VTAIL.n180 B 0.025693f
C470 VTAIL.n181 B 0.013806f
C471 VTAIL.n182 B 0.014618f
C472 VTAIL.n183 B 0.032633f
C473 VTAIL.n184 B 0.032633f
C474 VTAIL.n185 B 0.014618f
C475 VTAIL.n186 B 0.013806f
C476 VTAIL.n187 B 0.025693f
C477 VTAIL.n188 B 0.025693f
C478 VTAIL.n189 B 0.013806f
C479 VTAIL.n190 B 0.013806f
C480 VTAIL.n191 B 0.014618f
C481 VTAIL.n192 B 0.032633f
C482 VTAIL.n193 B 0.032633f
C483 VTAIL.n194 B 0.032633f
C484 VTAIL.n195 B 0.014212f
C485 VTAIL.n196 B 0.013806f
C486 VTAIL.n197 B 0.025693f
C487 VTAIL.n198 B 0.025693f
C488 VTAIL.n199 B 0.013806f
C489 VTAIL.n200 B 0.014618f
C490 VTAIL.n201 B 0.032633f
C491 VTAIL.n202 B 0.070645f
C492 VTAIL.n203 B 0.014618f
C493 VTAIL.n204 B 0.013806f
C494 VTAIL.n205 B 0.065004f
C495 VTAIL.n206 B 0.039694f
C496 VTAIL.n207 B 1.5635f
C497 VP.n0 B 0.036368f
C498 VP.t0 B 1.89573f
C499 VP.n1 B 0.036864f
C500 VP.n2 B 0.019329f
C501 VP.n3 B 0.036204f
C502 VP.n4 B 0.019329f
C503 VP.t5 B 1.89573f
C504 VP.n5 B 0.036204f
C505 VP.n6 B 0.019329f
C506 VP.n7 B 0.036204f
C507 VP.n8 B 0.036368f
C508 VP.t4 B 1.89573f
C509 VP.n9 B 0.036864f
C510 VP.n10 B 0.019329f
C511 VP.n11 B 0.036204f
C512 VP.t1 B 2.18777f
C513 VP.n12 B 0.711117f
C514 VP.t3 B 1.89573f
C515 VP.n13 B 0.743267f
C516 VP.n14 B 0.027267f
C517 VP.n15 B 0.254238f
C518 VP.n16 B 0.019329f
C519 VP.n17 B 0.019329f
C520 VP.n18 B 0.036204f
C521 VP.n19 B 0.033395f
C522 VP.n20 B 0.022624f
C523 VP.n21 B 0.019329f
C524 VP.n22 B 0.019329f
C525 VP.n23 B 0.019329f
C526 VP.n24 B 0.036204f
C527 VP.n25 B 0.034059f
C528 VP.n26 B 0.75829f
C529 VP.n27 B 1.18201f
C530 VP.n28 B 1.19536f
C531 VP.t2 B 1.89573f
C532 VP.n29 B 0.75829f
C533 VP.n30 B 0.034059f
C534 VP.n31 B 0.036368f
C535 VP.n32 B 0.019329f
C536 VP.n33 B 0.019329f
C537 VP.n34 B 0.036864f
C538 VP.n35 B 0.022624f
C539 VP.n36 B 0.033395f
C540 VP.n37 B 0.019329f
C541 VP.n38 B 0.019329f
C542 VP.n39 B 0.019329f
C543 VP.n40 B 0.036204f
C544 VP.n41 B 0.027267f
C545 VP.n42 B 0.673019f
C546 VP.n43 B 0.027267f
C547 VP.n44 B 0.019329f
C548 VP.n45 B 0.019329f
C549 VP.n46 B 0.019329f
C550 VP.n47 B 0.036204f
C551 VP.n48 B 0.033395f
C552 VP.n49 B 0.022624f
C553 VP.n50 B 0.019329f
C554 VP.n51 B 0.019329f
C555 VP.n52 B 0.019329f
C556 VP.n53 B 0.036204f
C557 VP.n54 B 0.034059f
C558 VP.n55 B 0.75829f
C559 VP.n56 B 0.05932f
.ends

