* NGSPICE file created from diff_pair_sample_0369.ext - technology: sky130A

.subckt diff_pair_sample_0369 VTAIL VN VP B VDD2 VDD1
X0 B.t17 B.t15 B.t16 B.t9 sky130_fd_pr__nfet_01v8 ad=3.6348 pd=19.42 as=0 ps=0 w=9.32 l=1.86
X1 VTAIL.t7 VN.t0 VDD2.t3 B.t0 sky130_fd_pr__nfet_01v8 ad=3.6348 pd=19.42 as=1.5378 ps=9.65 w=9.32 l=1.86
X2 B.t14 B.t12 B.t13 B.t5 sky130_fd_pr__nfet_01v8 ad=3.6348 pd=19.42 as=0 ps=0 w=9.32 l=1.86
X3 VDD1.t3 VP.t0 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=1.5378 pd=9.65 as=3.6348 ps=19.42 w=9.32 l=1.86
X4 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=3.6348 pd=19.42 as=0 ps=0 w=9.32 l=1.86
X5 VTAIL.t6 VN.t1 VDD2.t0 B.t3 sky130_fd_pr__nfet_01v8 ad=3.6348 pd=19.42 as=1.5378 ps=9.65 w=9.32 l=1.86
X6 B.t7 B.t4 B.t6 B.t5 sky130_fd_pr__nfet_01v8 ad=3.6348 pd=19.42 as=0 ps=0 w=9.32 l=1.86
X7 VTAIL.t3 VP.t1 VDD1.t2 B.t3 sky130_fd_pr__nfet_01v8 ad=3.6348 pd=19.42 as=1.5378 ps=9.65 w=9.32 l=1.86
X8 VTAIL.t0 VP.t2 VDD1.t1 B.t0 sky130_fd_pr__nfet_01v8 ad=3.6348 pd=19.42 as=1.5378 ps=9.65 w=9.32 l=1.86
X9 VDD2.t2 VN.t2 VTAIL.t5 B.t1 sky130_fd_pr__nfet_01v8 ad=1.5378 pd=9.65 as=3.6348 ps=19.42 w=9.32 l=1.86
X10 VDD2.t1 VN.t3 VTAIL.t4 B.t2 sky130_fd_pr__nfet_01v8 ad=1.5378 pd=9.65 as=3.6348 ps=19.42 w=9.32 l=1.86
X11 VDD1.t0 VP.t3 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=1.5378 pd=9.65 as=3.6348 ps=19.42 w=9.32 l=1.86
R0 B.n615 B.n614 585
R1 B.n616 B.n615 585
R2 B.n246 B.n92 585
R3 B.n245 B.n244 585
R4 B.n243 B.n242 585
R5 B.n241 B.n240 585
R6 B.n239 B.n238 585
R7 B.n237 B.n236 585
R8 B.n235 B.n234 585
R9 B.n233 B.n232 585
R10 B.n231 B.n230 585
R11 B.n229 B.n228 585
R12 B.n227 B.n226 585
R13 B.n225 B.n224 585
R14 B.n223 B.n222 585
R15 B.n221 B.n220 585
R16 B.n219 B.n218 585
R17 B.n217 B.n216 585
R18 B.n215 B.n214 585
R19 B.n213 B.n212 585
R20 B.n211 B.n210 585
R21 B.n209 B.n208 585
R22 B.n207 B.n206 585
R23 B.n205 B.n204 585
R24 B.n203 B.n202 585
R25 B.n201 B.n200 585
R26 B.n199 B.n198 585
R27 B.n197 B.n196 585
R28 B.n195 B.n194 585
R29 B.n193 B.n192 585
R30 B.n191 B.n190 585
R31 B.n189 B.n188 585
R32 B.n187 B.n186 585
R33 B.n185 B.n184 585
R34 B.n183 B.n182 585
R35 B.n180 B.n179 585
R36 B.n178 B.n177 585
R37 B.n176 B.n175 585
R38 B.n174 B.n173 585
R39 B.n172 B.n171 585
R40 B.n170 B.n169 585
R41 B.n168 B.n167 585
R42 B.n166 B.n165 585
R43 B.n164 B.n163 585
R44 B.n162 B.n161 585
R45 B.n160 B.n159 585
R46 B.n158 B.n157 585
R47 B.n156 B.n155 585
R48 B.n154 B.n153 585
R49 B.n152 B.n151 585
R50 B.n150 B.n149 585
R51 B.n148 B.n147 585
R52 B.n146 B.n145 585
R53 B.n144 B.n143 585
R54 B.n142 B.n141 585
R55 B.n140 B.n139 585
R56 B.n138 B.n137 585
R57 B.n136 B.n135 585
R58 B.n134 B.n133 585
R59 B.n132 B.n131 585
R60 B.n130 B.n129 585
R61 B.n128 B.n127 585
R62 B.n126 B.n125 585
R63 B.n124 B.n123 585
R64 B.n122 B.n121 585
R65 B.n120 B.n119 585
R66 B.n118 B.n117 585
R67 B.n116 B.n115 585
R68 B.n114 B.n113 585
R69 B.n112 B.n111 585
R70 B.n110 B.n109 585
R71 B.n108 B.n107 585
R72 B.n106 B.n105 585
R73 B.n104 B.n103 585
R74 B.n102 B.n101 585
R75 B.n100 B.n99 585
R76 B.n54 B.n53 585
R77 B.n619 B.n618 585
R78 B.n613 B.n93 585
R79 B.n93 B.n51 585
R80 B.n612 B.n50 585
R81 B.n623 B.n50 585
R82 B.n611 B.n49 585
R83 B.n624 B.n49 585
R84 B.n610 B.n48 585
R85 B.n625 B.n48 585
R86 B.n609 B.n608 585
R87 B.n608 B.n44 585
R88 B.n607 B.n43 585
R89 B.n631 B.n43 585
R90 B.n606 B.n42 585
R91 B.n632 B.n42 585
R92 B.n605 B.n41 585
R93 B.n633 B.n41 585
R94 B.n604 B.n603 585
R95 B.n603 B.n37 585
R96 B.n602 B.n36 585
R97 B.n639 B.n36 585
R98 B.n601 B.n35 585
R99 B.n640 B.n35 585
R100 B.n600 B.n34 585
R101 B.n641 B.n34 585
R102 B.n599 B.n598 585
R103 B.n598 B.n30 585
R104 B.n597 B.n29 585
R105 B.n647 B.n29 585
R106 B.n596 B.n28 585
R107 B.n648 B.n28 585
R108 B.n595 B.n27 585
R109 B.n649 B.n27 585
R110 B.n594 B.n593 585
R111 B.n593 B.n26 585
R112 B.n592 B.n22 585
R113 B.n655 B.n22 585
R114 B.n591 B.n21 585
R115 B.n656 B.n21 585
R116 B.n590 B.n20 585
R117 B.n657 B.n20 585
R118 B.n589 B.n588 585
R119 B.n588 B.n16 585
R120 B.n587 B.n15 585
R121 B.n663 B.n15 585
R122 B.n586 B.n14 585
R123 B.n664 B.n14 585
R124 B.n585 B.n13 585
R125 B.n665 B.n13 585
R126 B.n584 B.n583 585
R127 B.n583 B.n12 585
R128 B.n582 B.n581 585
R129 B.n582 B.n8 585
R130 B.n580 B.n7 585
R131 B.n672 B.n7 585
R132 B.n579 B.n6 585
R133 B.n673 B.n6 585
R134 B.n578 B.n5 585
R135 B.n674 B.n5 585
R136 B.n577 B.n576 585
R137 B.n576 B.n4 585
R138 B.n575 B.n247 585
R139 B.n575 B.n574 585
R140 B.n565 B.n248 585
R141 B.n249 B.n248 585
R142 B.n567 B.n566 585
R143 B.n568 B.n567 585
R144 B.n564 B.n253 585
R145 B.n257 B.n253 585
R146 B.n563 B.n562 585
R147 B.n562 B.n561 585
R148 B.n255 B.n254 585
R149 B.n256 B.n255 585
R150 B.n554 B.n553 585
R151 B.n555 B.n554 585
R152 B.n552 B.n262 585
R153 B.n262 B.n261 585
R154 B.n551 B.n550 585
R155 B.n550 B.n549 585
R156 B.n264 B.n263 585
R157 B.n542 B.n264 585
R158 B.n541 B.n540 585
R159 B.n543 B.n541 585
R160 B.n539 B.n269 585
R161 B.n269 B.n268 585
R162 B.n538 B.n537 585
R163 B.n537 B.n536 585
R164 B.n271 B.n270 585
R165 B.n272 B.n271 585
R166 B.n529 B.n528 585
R167 B.n530 B.n529 585
R168 B.n527 B.n277 585
R169 B.n277 B.n276 585
R170 B.n526 B.n525 585
R171 B.n525 B.n524 585
R172 B.n279 B.n278 585
R173 B.n280 B.n279 585
R174 B.n517 B.n516 585
R175 B.n518 B.n517 585
R176 B.n515 B.n284 585
R177 B.n288 B.n284 585
R178 B.n514 B.n513 585
R179 B.n513 B.n512 585
R180 B.n286 B.n285 585
R181 B.n287 B.n286 585
R182 B.n505 B.n504 585
R183 B.n506 B.n505 585
R184 B.n503 B.n293 585
R185 B.n293 B.n292 585
R186 B.n502 B.n501 585
R187 B.n501 B.n500 585
R188 B.n295 B.n294 585
R189 B.n296 B.n295 585
R190 B.n496 B.n495 585
R191 B.n299 B.n298 585
R192 B.n492 B.n491 585
R193 B.n493 B.n492 585
R194 B.n490 B.n337 585
R195 B.n489 B.n488 585
R196 B.n487 B.n486 585
R197 B.n485 B.n484 585
R198 B.n483 B.n482 585
R199 B.n481 B.n480 585
R200 B.n479 B.n478 585
R201 B.n477 B.n476 585
R202 B.n475 B.n474 585
R203 B.n473 B.n472 585
R204 B.n471 B.n470 585
R205 B.n469 B.n468 585
R206 B.n467 B.n466 585
R207 B.n465 B.n464 585
R208 B.n463 B.n462 585
R209 B.n461 B.n460 585
R210 B.n459 B.n458 585
R211 B.n457 B.n456 585
R212 B.n455 B.n454 585
R213 B.n453 B.n452 585
R214 B.n451 B.n450 585
R215 B.n449 B.n448 585
R216 B.n447 B.n446 585
R217 B.n445 B.n444 585
R218 B.n443 B.n442 585
R219 B.n441 B.n440 585
R220 B.n439 B.n438 585
R221 B.n437 B.n436 585
R222 B.n435 B.n434 585
R223 B.n433 B.n432 585
R224 B.n431 B.n430 585
R225 B.n428 B.n427 585
R226 B.n426 B.n425 585
R227 B.n424 B.n423 585
R228 B.n422 B.n421 585
R229 B.n420 B.n419 585
R230 B.n418 B.n417 585
R231 B.n416 B.n415 585
R232 B.n414 B.n413 585
R233 B.n412 B.n411 585
R234 B.n410 B.n409 585
R235 B.n408 B.n407 585
R236 B.n406 B.n405 585
R237 B.n404 B.n403 585
R238 B.n402 B.n401 585
R239 B.n400 B.n399 585
R240 B.n398 B.n397 585
R241 B.n396 B.n395 585
R242 B.n394 B.n393 585
R243 B.n392 B.n391 585
R244 B.n390 B.n389 585
R245 B.n388 B.n387 585
R246 B.n386 B.n385 585
R247 B.n384 B.n383 585
R248 B.n382 B.n381 585
R249 B.n380 B.n379 585
R250 B.n378 B.n377 585
R251 B.n376 B.n375 585
R252 B.n374 B.n373 585
R253 B.n372 B.n371 585
R254 B.n370 B.n369 585
R255 B.n368 B.n367 585
R256 B.n366 B.n365 585
R257 B.n364 B.n363 585
R258 B.n362 B.n361 585
R259 B.n360 B.n359 585
R260 B.n358 B.n357 585
R261 B.n356 B.n355 585
R262 B.n354 B.n353 585
R263 B.n352 B.n351 585
R264 B.n350 B.n349 585
R265 B.n348 B.n347 585
R266 B.n346 B.n345 585
R267 B.n344 B.n343 585
R268 B.n497 B.n297 585
R269 B.n297 B.n296 585
R270 B.n499 B.n498 585
R271 B.n500 B.n499 585
R272 B.n291 B.n290 585
R273 B.n292 B.n291 585
R274 B.n508 B.n507 585
R275 B.n507 B.n506 585
R276 B.n509 B.n289 585
R277 B.n289 B.n287 585
R278 B.n511 B.n510 585
R279 B.n512 B.n511 585
R280 B.n283 B.n282 585
R281 B.n288 B.n283 585
R282 B.n520 B.n519 585
R283 B.n519 B.n518 585
R284 B.n521 B.n281 585
R285 B.n281 B.n280 585
R286 B.n523 B.n522 585
R287 B.n524 B.n523 585
R288 B.n275 B.n274 585
R289 B.n276 B.n275 585
R290 B.n532 B.n531 585
R291 B.n531 B.n530 585
R292 B.n533 B.n273 585
R293 B.n273 B.n272 585
R294 B.n535 B.n534 585
R295 B.n536 B.n535 585
R296 B.n267 B.n266 585
R297 B.n268 B.n267 585
R298 B.n545 B.n544 585
R299 B.n544 B.n543 585
R300 B.n546 B.n265 585
R301 B.n542 B.n265 585
R302 B.n548 B.n547 585
R303 B.n549 B.n548 585
R304 B.n260 B.n259 585
R305 B.n261 B.n260 585
R306 B.n557 B.n556 585
R307 B.n556 B.n555 585
R308 B.n558 B.n258 585
R309 B.n258 B.n256 585
R310 B.n560 B.n559 585
R311 B.n561 B.n560 585
R312 B.n252 B.n251 585
R313 B.n257 B.n252 585
R314 B.n570 B.n569 585
R315 B.n569 B.n568 585
R316 B.n571 B.n250 585
R317 B.n250 B.n249 585
R318 B.n573 B.n572 585
R319 B.n574 B.n573 585
R320 B.n3 B.n0 585
R321 B.n4 B.n3 585
R322 B.n671 B.n1 585
R323 B.n672 B.n671 585
R324 B.n670 B.n669 585
R325 B.n670 B.n8 585
R326 B.n668 B.n9 585
R327 B.n12 B.n9 585
R328 B.n667 B.n666 585
R329 B.n666 B.n665 585
R330 B.n11 B.n10 585
R331 B.n664 B.n11 585
R332 B.n662 B.n661 585
R333 B.n663 B.n662 585
R334 B.n660 B.n17 585
R335 B.n17 B.n16 585
R336 B.n659 B.n658 585
R337 B.n658 B.n657 585
R338 B.n19 B.n18 585
R339 B.n656 B.n19 585
R340 B.n654 B.n653 585
R341 B.n655 B.n654 585
R342 B.n652 B.n23 585
R343 B.n26 B.n23 585
R344 B.n651 B.n650 585
R345 B.n650 B.n649 585
R346 B.n25 B.n24 585
R347 B.n648 B.n25 585
R348 B.n646 B.n645 585
R349 B.n647 B.n646 585
R350 B.n644 B.n31 585
R351 B.n31 B.n30 585
R352 B.n643 B.n642 585
R353 B.n642 B.n641 585
R354 B.n33 B.n32 585
R355 B.n640 B.n33 585
R356 B.n638 B.n637 585
R357 B.n639 B.n638 585
R358 B.n636 B.n38 585
R359 B.n38 B.n37 585
R360 B.n635 B.n634 585
R361 B.n634 B.n633 585
R362 B.n40 B.n39 585
R363 B.n632 B.n40 585
R364 B.n630 B.n629 585
R365 B.n631 B.n630 585
R366 B.n628 B.n45 585
R367 B.n45 B.n44 585
R368 B.n627 B.n626 585
R369 B.n626 B.n625 585
R370 B.n47 B.n46 585
R371 B.n624 B.n47 585
R372 B.n622 B.n621 585
R373 B.n623 B.n622 585
R374 B.n620 B.n52 585
R375 B.n52 B.n51 585
R376 B.n675 B.n674 585
R377 B.n673 B.n2 585
R378 B.n618 B.n52 492.5
R379 B.n615 B.n93 492.5
R380 B.n343 B.n295 492.5
R381 B.n495 B.n297 492.5
R382 B.n96 B.t15 327.329
R383 B.n94 B.t8 327.329
R384 B.n340 B.t12 327.329
R385 B.n338 B.t4 327.329
R386 B.n94 B.t10 278.409
R387 B.n340 B.t14 278.409
R388 B.n96 B.t16 278.409
R389 B.n338 B.t7 278.409
R390 B.n616 B.n91 256.663
R391 B.n616 B.n90 256.663
R392 B.n616 B.n89 256.663
R393 B.n616 B.n88 256.663
R394 B.n616 B.n87 256.663
R395 B.n616 B.n86 256.663
R396 B.n616 B.n85 256.663
R397 B.n616 B.n84 256.663
R398 B.n616 B.n83 256.663
R399 B.n616 B.n82 256.663
R400 B.n616 B.n81 256.663
R401 B.n616 B.n80 256.663
R402 B.n616 B.n79 256.663
R403 B.n616 B.n78 256.663
R404 B.n616 B.n77 256.663
R405 B.n616 B.n76 256.663
R406 B.n616 B.n75 256.663
R407 B.n616 B.n74 256.663
R408 B.n616 B.n73 256.663
R409 B.n616 B.n72 256.663
R410 B.n616 B.n71 256.663
R411 B.n616 B.n70 256.663
R412 B.n616 B.n69 256.663
R413 B.n616 B.n68 256.663
R414 B.n616 B.n67 256.663
R415 B.n616 B.n66 256.663
R416 B.n616 B.n65 256.663
R417 B.n616 B.n64 256.663
R418 B.n616 B.n63 256.663
R419 B.n616 B.n62 256.663
R420 B.n616 B.n61 256.663
R421 B.n616 B.n60 256.663
R422 B.n616 B.n59 256.663
R423 B.n616 B.n58 256.663
R424 B.n616 B.n57 256.663
R425 B.n616 B.n56 256.663
R426 B.n616 B.n55 256.663
R427 B.n617 B.n616 256.663
R428 B.n494 B.n493 256.663
R429 B.n493 B.n300 256.663
R430 B.n493 B.n301 256.663
R431 B.n493 B.n302 256.663
R432 B.n493 B.n303 256.663
R433 B.n493 B.n304 256.663
R434 B.n493 B.n305 256.663
R435 B.n493 B.n306 256.663
R436 B.n493 B.n307 256.663
R437 B.n493 B.n308 256.663
R438 B.n493 B.n309 256.663
R439 B.n493 B.n310 256.663
R440 B.n493 B.n311 256.663
R441 B.n493 B.n312 256.663
R442 B.n493 B.n313 256.663
R443 B.n493 B.n314 256.663
R444 B.n493 B.n315 256.663
R445 B.n493 B.n316 256.663
R446 B.n493 B.n317 256.663
R447 B.n493 B.n318 256.663
R448 B.n493 B.n319 256.663
R449 B.n493 B.n320 256.663
R450 B.n493 B.n321 256.663
R451 B.n493 B.n322 256.663
R452 B.n493 B.n323 256.663
R453 B.n493 B.n324 256.663
R454 B.n493 B.n325 256.663
R455 B.n493 B.n326 256.663
R456 B.n493 B.n327 256.663
R457 B.n493 B.n328 256.663
R458 B.n493 B.n329 256.663
R459 B.n493 B.n330 256.663
R460 B.n493 B.n331 256.663
R461 B.n493 B.n332 256.663
R462 B.n493 B.n333 256.663
R463 B.n493 B.n334 256.663
R464 B.n493 B.n335 256.663
R465 B.n493 B.n336 256.663
R466 B.n677 B.n676 256.663
R467 B.n95 B.t11 235.935
R468 B.n341 B.t13 235.935
R469 B.n97 B.t17 235.935
R470 B.n339 B.t6 235.935
R471 B.n99 B.n54 163.367
R472 B.n103 B.n102 163.367
R473 B.n107 B.n106 163.367
R474 B.n111 B.n110 163.367
R475 B.n115 B.n114 163.367
R476 B.n119 B.n118 163.367
R477 B.n123 B.n122 163.367
R478 B.n127 B.n126 163.367
R479 B.n131 B.n130 163.367
R480 B.n135 B.n134 163.367
R481 B.n139 B.n138 163.367
R482 B.n143 B.n142 163.367
R483 B.n147 B.n146 163.367
R484 B.n151 B.n150 163.367
R485 B.n155 B.n154 163.367
R486 B.n159 B.n158 163.367
R487 B.n163 B.n162 163.367
R488 B.n167 B.n166 163.367
R489 B.n171 B.n170 163.367
R490 B.n175 B.n174 163.367
R491 B.n179 B.n178 163.367
R492 B.n184 B.n183 163.367
R493 B.n188 B.n187 163.367
R494 B.n192 B.n191 163.367
R495 B.n196 B.n195 163.367
R496 B.n200 B.n199 163.367
R497 B.n204 B.n203 163.367
R498 B.n208 B.n207 163.367
R499 B.n212 B.n211 163.367
R500 B.n216 B.n215 163.367
R501 B.n220 B.n219 163.367
R502 B.n224 B.n223 163.367
R503 B.n228 B.n227 163.367
R504 B.n232 B.n231 163.367
R505 B.n236 B.n235 163.367
R506 B.n240 B.n239 163.367
R507 B.n244 B.n243 163.367
R508 B.n615 B.n92 163.367
R509 B.n501 B.n295 163.367
R510 B.n501 B.n293 163.367
R511 B.n505 B.n293 163.367
R512 B.n505 B.n286 163.367
R513 B.n513 B.n286 163.367
R514 B.n513 B.n284 163.367
R515 B.n517 B.n284 163.367
R516 B.n517 B.n279 163.367
R517 B.n525 B.n279 163.367
R518 B.n525 B.n277 163.367
R519 B.n529 B.n277 163.367
R520 B.n529 B.n271 163.367
R521 B.n537 B.n271 163.367
R522 B.n537 B.n269 163.367
R523 B.n541 B.n269 163.367
R524 B.n541 B.n264 163.367
R525 B.n550 B.n264 163.367
R526 B.n550 B.n262 163.367
R527 B.n554 B.n262 163.367
R528 B.n554 B.n255 163.367
R529 B.n562 B.n255 163.367
R530 B.n562 B.n253 163.367
R531 B.n567 B.n253 163.367
R532 B.n567 B.n248 163.367
R533 B.n575 B.n248 163.367
R534 B.n576 B.n575 163.367
R535 B.n576 B.n5 163.367
R536 B.n6 B.n5 163.367
R537 B.n7 B.n6 163.367
R538 B.n582 B.n7 163.367
R539 B.n583 B.n582 163.367
R540 B.n583 B.n13 163.367
R541 B.n14 B.n13 163.367
R542 B.n15 B.n14 163.367
R543 B.n588 B.n15 163.367
R544 B.n588 B.n20 163.367
R545 B.n21 B.n20 163.367
R546 B.n22 B.n21 163.367
R547 B.n593 B.n22 163.367
R548 B.n593 B.n27 163.367
R549 B.n28 B.n27 163.367
R550 B.n29 B.n28 163.367
R551 B.n598 B.n29 163.367
R552 B.n598 B.n34 163.367
R553 B.n35 B.n34 163.367
R554 B.n36 B.n35 163.367
R555 B.n603 B.n36 163.367
R556 B.n603 B.n41 163.367
R557 B.n42 B.n41 163.367
R558 B.n43 B.n42 163.367
R559 B.n608 B.n43 163.367
R560 B.n608 B.n48 163.367
R561 B.n49 B.n48 163.367
R562 B.n50 B.n49 163.367
R563 B.n93 B.n50 163.367
R564 B.n492 B.n299 163.367
R565 B.n492 B.n337 163.367
R566 B.n488 B.n487 163.367
R567 B.n484 B.n483 163.367
R568 B.n480 B.n479 163.367
R569 B.n476 B.n475 163.367
R570 B.n472 B.n471 163.367
R571 B.n468 B.n467 163.367
R572 B.n464 B.n463 163.367
R573 B.n460 B.n459 163.367
R574 B.n456 B.n455 163.367
R575 B.n452 B.n451 163.367
R576 B.n448 B.n447 163.367
R577 B.n444 B.n443 163.367
R578 B.n440 B.n439 163.367
R579 B.n436 B.n435 163.367
R580 B.n432 B.n431 163.367
R581 B.n427 B.n426 163.367
R582 B.n423 B.n422 163.367
R583 B.n419 B.n418 163.367
R584 B.n415 B.n414 163.367
R585 B.n411 B.n410 163.367
R586 B.n407 B.n406 163.367
R587 B.n403 B.n402 163.367
R588 B.n399 B.n398 163.367
R589 B.n395 B.n394 163.367
R590 B.n391 B.n390 163.367
R591 B.n387 B.n386 163.367
R592 B.n383 B.n382 163.367
R593 B.n379 B.n378 163.367
R594 B.n375 B.n374 163.367
R595 B.n371 B.n370 163.367
R596 B.n367 B.n366 163.367
R597 B.n363 B.n362 163.367
R598 B.n359 B.n358 163.367
R599 B.n355 B.n354 163.367
R600 B.n351 B.n350 163.367
R601 B.n347 B.n346 163.367
R602 B.n499 B.n297 163.367
R603 B.n499 B.n291 163.367
R604 B.n507 B.n291 163.367
R605 B.n507 B.n289 163.367
R606 B.n511 B.n289 163.367
R607 B.n511 B.n283 163.367
R608 B.n519 B.n283 163.367
R609 B.n519 B.n281 163.367
R610 B.n523 B.n281 163.367
R611 B.n523 B.n275 163.367
R612 B.n531 B.n275 163.367
R613 B.n531 B.n273 163.367
R614 B.n535 B.n273 163.367
R615 B.n535 B.n267 163.367
R616 B.n544 B.n267 163.367
R617 B.n544 B.n265 163.367
R618 B.n548 B.n265 163.367
R619 B.n548 B.n260 163.367
R620 B.n556 B.n260 163.367
R621 B.n556 B.n258 163.367
R622 B.n560 B.n258 163.367
R623 B.n560 B.n252 163.367
R624 B.n569 B.n252 163.367
R625 B.n569 B.n250 163.367
R626 B.n573 B.n250 163.367
R627 B.n573 B.n3 163.367
R628 B.n675 B.n3 163.367
R629 B.n671 B.n2 163.367
R630 B.n671 B.n670 163.367
R631 B.n670 B.n9 163.367
R632 B.n666 B.n9 163.367
R633 B.n666 B.n11 163.367
R634 B.n662 B.n11 163.367
R635 B.n662 B.n17 163.367
R636 B.n658 B.n17 163.367
R637 B.n658 B.n19 163.367
R638 B.n654 B.n19 163.367
R639 B.n654 B.n23 163.367
R640 B.n650 B.n23 163.367
R641 B.n650 B.n25 163.367
R642 B.n646 B.n25 163.367
R643 B.n646 B.n31 163.367
R644 B.n642 B.n31 163.367
R645 B.n642 B.n33 163.367
R646 B.n638 B.n33 163.367
R647 B.n638 B.n38 163.367
R648 B.n634 B.n38 163.367
R649 B.n634 B.n40 163.367
R650 B.n630 B.n40 163.367
R651 B.n630 B.n45 163.367
R652 B.n626 B.n45 163.367
R653 B.n626 B.n47 163.367
R654 B.n622 B.n47 163.367
R655 B.n622 B.n52 163.367
R656 B.n493 B.n296 89.6887
R657 B.n616 B.n51 89.6887
R658 B.n618 B.n617 71.676
R659 B.n99 B.n55 71.676
R660 B.n103 B.n56 71.676
R661 B.n107 B.n57 71.676
R662 B.n111 B.n58 71.676
R663 B.n115 B.n59 71.676
R664 B.n119 B.n60 71.676
R665 B.n123 B.n61 71.676
R666 B.n127 B.n62 71.676
R667 B.n131 B.n63 71.676
R668 B.n135 B.n64 71.676
R669 B.n139 B.n65 71.676
R670 B.n143 B.n66 71.676
R671 B.n147 B.n67 71.676
R672 B.n151 B.n68 71.676
R673 B.n155 B.n69 71.676
R674 B.n159 B.n70 71.676
R675 B.n163 B.n71 71.676
R676 B.n167 B.n72 71.676
R677 B.n171 B.n73 71.676
R678 B.n175 B.n74 71.676
R679 B.n179 B.n75 71.676
R680 B.n184 B.n76 71.676
R681 B.n188 B.n77 71.676
R682 B.n192 B.n78 71.676
R683 B.n196 B.n79 71.676
R684 B.n200 B.n80 71.676
R685 B.n204 B.n81 71.676
R686 B.n208 B.n82 71.676
R687 B.n212 B.n83 71.676
R688 B.n216 B.n84 71.676
R689 B.n220 B.n85 71.676
R690 B.n224 B.n86 71.676
R691 B.n228 B.n87 71.676
R692 B.n232 B.n88 71.676
R693 B.n236 B.n89 71.676
R694 B.n240 B.n90 71.676
R695 B.n244 B.n91 71.676
R696 B.n92 B.n91 71.676
R697 B.n243 B.n90 71.676
R698 B.n239 B.n89 71.676
R699 B.n235 B.n88 71.676
R700 B.n231 B.n87 71.676
R701 B.n227 B.n86 71.676
R702 B.n223 B.n85 71.676
R703 B.n219 B.n84 71.676
R704 B.n215 B.n83 71.676
R705 B.n211 B.n82 71.676
R706 B.n207 B.n81 71.676
R707 B.n203 B.n80 71.676
R708 B.n199 B.n79 71.676
R709 B.n195 B.n78 71.676
R710 B.n191 B.n77 71.676
R711 B.n187 B.n76 71.676
R712 B.n183 B.n75 71.676
R713 B.n178 B.n74 71.676
R714 B.n174 B.n73 71.676
R715 B.n170 B.n72 71.676
R716 B.n166 B.n71 71.676
R717 B.n162 B.n70 71.676
R718 B.n158 B.n69 71.676
R719 B.n154 B.n68 71.676
R720 B.n150 B.n67 71.676
R721 B.n146 B.n66 71.676
R722 B.n142 B.n65 71.676
R723 B.n138 B.n64 71.676
R724 B.n134 B.n63 71.676
R725 B.n130 B.n62 71.676
R726 B.n126 B.n61 71.676
R727 B.n122 B.n60 71.676
R728 B.n118 B.n59 71.676
R729 B.n114 B.n58 71.676
R730 B.n110 B.n57 71.676
R731 B.n106 B.n56 71.676
R732 B.n102 B.n55 71.676
R733 B.n617 B.n54 71.676
R734 B.n495 B.n494 71.676
R735 B.n337 B.n300 71.676
R736 B.n487 B.n301 71.676
R737 B.n483 B.n302 71.676
R738 B.n479 B.n303 71.676
R739 B.n475 B.n304 71.676
R740 B.n471 B.n305 71.676
R741 B.n467 B.n306 71.676
R742 B.n463 B.n307 71.676
R743 B.n459 B.n308 71.676
R744 B.n455 B.n309 71.676
R745 B.n451 B.n310 71.676
R746 B.n447 B.n311 71.676
R747 B.n443 B.n312 71.676
R748 B.n439 B.n313 71.676
R749 B.n435 B.n314 71.676
R750 B.n431 B.n315 71.676
R751 B.n426 B.n316 71.676
R752 B.n422 B.n317 71.676
R753 B.n418 B.n318 71.676
R754 B.n414 B.n319 71.676
R755 B.n410 B.n320 71.676
R756 B.n406 B.n321 71.676
R757 B.n402 B.n322 71.676
R758 B.n398 B.n323 71.676
R759 B.n394 B.n324 71.676
R760 B.n390 B.n325 71.676
R761 B.n386 B.n326 71.676
R762 B.n382 B.n327 71.676
R763 B.n378 B.n328 71.676
R764 B.n374 B.n329 71.676
R765 B.n370 B.n330 71.676
R766 B.n366 B.n331 71.676
R767 B.n362 B.n332 71.676
R768 B.n358 B.n333 71.676
R769 B.n354 B.n334 71.676
R770 B.n350 B.n335 71.676
R771 B.n346 B.n336 71.676
R772 B.n494 B.n299 71.676
R773 B.n488 B.n300 71.676
R774 B.n484 B.n301 71.676
R775 B.n480 B.n302 71.676
R776 B.n476 B.n303 71.676
R777 B.n472 B.n304 71.676
R778 B.n468 B.n305 71.676
R779 B.n464 B.n306 71.676
R780 B.n460 B.n307 71.676
R781 B.n456 B.n308 71.676
R782 B.n452 B.n309 71.676
R783 B.n448 B.n310 71.676
R784 B.n444 B.n311 71.676
R785 B.n440 B.n312 71.676
R786 B.n436 B.n313 71.676
R787 B.n432 B.n314 71.676
R788 B.n427 B.n315 71.676
R789 B.n423 B.n316 71.676
R790 B.n419 B.n317 71.676
R791 B.n415 B.n318 71.676
R792 B.n411 B.n319 71.676
R793 B.n407 B.n320 71.676
R794 B.n403 B.n321 71.676
R795 B.n399 B.n322 71.676
R796 B.n395 B.n323 71.676
R797 B.n391 B.n324 71.676
R798 B.n387 B.n325 71.676
R799 B.n383 B.n326 71.676
R800 B.n379 B.n327 71.676
R801 B.n375 B.n328 71.676
R802 B.n371 B.n329 71.676
R803 B.n367 B.n330 71.676
R804 B.n363 B.n331 71.676
R805 B.n359 B.n332 71.676
R806 B.n355 B.n333 71.676
R807 B.n351 B.n334 71.676
R808 B.n347 B.n335 71.676
R809 B.n343 B.n336 71.676
R810 B.n676 B.n675 71.676
R811 B.n676 B.n2 71.676
R812 B.n98 B.n97 59.5399
R813 B.n181 B.n95 59.5399
R814 B.n342 B.n341 59.5399
R815 B.n429 B.n339 59.5399
R816 B.n500 B.n296 51.2509
R817 B.n500 B.n292 51.2509
R818 B.n506 B.n292 51.2509
R819 B.n506 B.n287 51.2509
R820 B.n512 B.n287 51.2509
R821 B.n512 B.n288 51.2509
R822 B.n518 B.n280 51.2509
R823 B.n524 B.n280 51.2509
R824 B.n524 B.n276 51.2509
R825 B.n530 B.n276 51.2509
R826 B.n530 B.n272 51.2509
R827 B.n536 B.n272 51.2509
R828 B.n536 B.n268 51.2509
R829 B.n543 B.n268 51.2509
R830 B.n543 B.n542 51.2509
R831 B.n549 B.n261 51.2509
R832 B.n555 B.n261 51.2509
R833 B.n555 B.n256 51.2509
R834 B.n561 B.n256 51.2509
R835 B.n561 B.n257 51.2509
R836 B.n568 B.n249 51.2509
R837 B.n574 B.n249 51.2509
R838 B.n574 B.n4 51.2509
R839 B.n674 B.n4 51.2509
R840 B.n674 B.n673 51.2509
R841 B.n673 B.n672 51.2509
R842 B.n672 B.n8 51.2509
R843 B.n12 B.n8 51.2509
R844 B.n665 B.n12 51.2509
R845 B.n664 B.n663 51.2509
R846 B.n663 B.n16 51.2509
R847 B.n657 B.n16 51.2509
R848 B.n657 B.n656 51.2509
R849 B.n656 B.n655 51.2509
R850 B.n649 B.n26 51.2509
R851 B.n649 B.n648 51.2509
R852 B.n648 B.n647 51.2509
R853 B.n647 B.n30 51.2509
R854 B.n641 B.n30 51.2509
R855 B.n641 B.n640 51.2509
R856 B.n640 B.n639 51.2509
R857 B.n639 B.n37 51.2509
R858 B.n633 B.n37 51.2509
R859 B.n632 B.n631 51.2509
R860 B.n631 B.n44 51.2509
R861 B.n625 B.n44 51.2509
R862 B.n625 B.n624 51.2509
R863 B.n624 B.n623 51.2509
R864 B.n623 B.n51 51.2509
R865 B.n97 B.n96 42.4732
R866 B.n95 B.n94 42.4732
R867 B.n341 B.n340 42.4732
R868 B.n339 B.n338 42.4732
R869 B.n549 B.t0 39.192
R870 B.n655 B.t1 39.192
R871 B.n257 B.t2 34.6699
R872 B.t3 B.n664 34.6699
R873 B.n497 B.n496 32.0005
R874 B.n344 B.n294 32.0005
R875 B.n614 B.n613 32.0005
R876 B.n620 B.n619 32.0005
R877 B.n288 B.t5 30.1478
R878 B.t9 B.n632 30.1478
R879 B.n518 B.t5 21.1036
R880 B.n633 B.t9 21.1036
R881 B B.n677 18.0485
R882 B.n568 B.t2 16.5815
R883 B.n665 B.t3 16.5815
R884 B.n542 B.t0 12.0594
R885 B.n26 B.t1 12.0594
R886 B.n498 B.n497 10.6151
R887 B.n498 B.n290 10.6151
R888 B.n508 B.n290 10.6151
R889 B.n509 B.n508 10.6151
R890 B.n510 B.n509 10.6151
R891 B.n510 B.n282 10.6151
R892 B.n520 B.n282 10.6151
R893 B.n521 B.n520 10.6151
R894 B.n522 B.n521 10.6151
R895 B.n522 B.n274 10.6151
R896 B.n532 B.n274 10.6151
R897 B.n533 B.n532 10.6151
R898 B.n534 B.n533 10.6151
R899 B.n534 B.n266 10.6151
R900 B.n545 B.n266 10.6151
R901 B.n546 B.n545 10.6151
R902 B.n547 B.n546 10.6151
R903 B.n547 B.n259 10.6151
R904 B.n557 B.n259 10.6151
R905 B.n558 B.n557 10.6151
R906 B.n559 B.n558 10.6151
R907 B.n559 B.n251 10.6151
R908 B.n570 B.n251 10.6151
R909 B.n571 B.n570 10.6151
R910 B.n572 B.n571 10.6151
R911 B.n572 B.n0 10.6151
R912 B.n496 B.n298 10.6151
R913 B.n491 B.n298 10.6151
R914 B.n491 B.n490 10.6151
R915 B.n490 B.n489 10.6151
R916 B.n489 B.n486 10.6151
R917 B.n486 B.n485 10.6151
R918 B.n485 B.n482 10.6151
R919 B.n482 B.n481 10.6151
R920 B.n481 B.n478 10.6151
R921 B.n478 B.n477 10.6151
R922 B.n477 B.n474 10.6151
R923 B.n474 B.n473 10.6151
R924 B.n473 B.n470 10.6151
R925 B.n470 B.n469 10.6151
R926 B.n469 B.n466 10.6151
R927 B.n466 B.n465 10.6151
R928 B.n465 B.n462 10.6151
R929 B.n462 B.n461 10.6151
R930 B.n461 B.n458 10.6151
R931 B.n458 B.n457 10.6151
R932 B.n457 B.n454 10.6151
R933 B.n454 B.n453 10.6151
R934 B.n453 B.n450 10.6151
R935 B.n450 B.n449 10.6151
R936 B.n449 B.n446 10.6151
R937 B.n446 B.n445 10.6151
R938 B.n445 B.n442 10.6151
R939 B.n442 B.n441 10.6151
R940 B.n441 B.n438 10.6151
R941 B.n438 B.n437 10.6151
R942 B.n437 B.n434 10.6151
R943 B.n434 B.n433 10.6151
R944 B.n433 B.n430 10.6151
R945 B.n428 B.n425 10.6151
R946 B.n425 B.n424 10.6151
R947 B.n424 B.n421 10.6151
R948 B.n421 B.n420 10.6151
R949 B.n420 B.n417 10.6151
R950 B.n417 B.n416 10.6151
R951 B.n416 B.n413 10.6151
R952 B.n413 B.n412 10.6151
R953 B.n409 B.n408 10.6151
R954 B.n408 B.n405 10.6151
R955 B.n405 B.n404 10.6151
R956 B.n404 B.n401 10.6151
R957 B.n401 B.n400 10.6151
R958 B.n400 B.n397 10.6151
R959 B.n397 B.n396 10.6151
R960 B.n396 B.n393 10.6151
R961 B.n393 B.n392 10.6151
R962 B.n392 B.n389 10.6151
R963 B.n389 B.n388 10.6151
R964 B.n388 B.n385 10.6151
R965 B.n385 B.n384 10.6151
R966 B.n384 B.n381 10.6151
R967 B.n381 B.n380 10.6151
R968 B.n380 B.n377 10.6151
R969 B.n377 B.n376 10.6151
R970 B.n376 B.n373 10.6151
R971 B.n373 B.n372 10.6151
R972 B.n372 B.n369 10.6151
R973 B.n369 B.n368 10.6151
R974 B.n368 B.n365 10.6151
R975 B.n365 B.n364 10.6151
R976 B.n364 B.n361 10.6151
R977 B.n361 B.n360 10.6151
R978 B.n360 B.n357 10.6151
R979 B.n357 B.n356 10.6151
R980 B.n356 B.n353 10.6151
R981 B.n353 B.n352 10.6151
R982 B.n352 B.n349 10.6151
R983 B.n349 B.n348 10.6151
R984 B.n348 B.n345 10.6151
R985 B.n345 B.n344 10.6151
R986 B.n502 B.n294 10.6151
R987 B.n503 B.n502 10.6151
R988 B.n504 B.n503 10.6151
R989 B.n504 B.n285 10.6151
R990 B.n514 B.n285 10.6151
R991 B.n515 B.n514 10.6151
R992 B.n516 B.n515 10.6151
R993 B.n516 B.n278 10.6151
R994 B.n526 B.n278 10.6151
R995 B.n527 B.n526 10.6151
R996 B.n528 B.n527 10.6151
R997 B.n528 B.n270 10.6151
R998 B.n538 B.n270 10.6151
R999 B.n539 B.n538 10.6151
R1000 B.n540 B.n539 10.6151
R1001 B.n540 B.n263 10.6151
R1002 B.n551 B.n263 10.6151
R1003 B.n552 B.n551 10.6151
R1004 B.n553 B.n552 10.6151
R1005 B.n553 B.n254 10.6151
R1006 B.n563 B.n254 10.6151
R1007 B.n564 B.n563 10.6151
R1008 B.n566 B.n564 10.6151
R1009 B.n566 B.n565 10.6151
R1010 B.n565 B.n247 10.6151
R1011 B.n577 B.n247 10.6151
R1012 B.n578 B.n577 10.6151
R1013 B.n579 B.n578 10.6151
R1014 B.n580 B.n579 10.6151
R1015 B.n581 B.n580 10.6151
R1016 B.n584 B.n581 10.6151
R1017 B.n585 B.n584 10.6151
R1018 B.n586 B.n585 10.6151
R1019 B.n587 B.n586 10.6151
R1020 B.n589 B.n587 10.6151
R1021 B.n590 B.n589 10.6151
R1022 B.n591 B.n590 10.6151
R1023 B.n592 B.n591 10.6151
R1024 B.n594 B.n592 10.6151
R1025 B.n595 B.n594 10.6151
R1026 B.n596 B.n595 10.6151
R1027 B.n597 B.n596 10.6151
R1028 B.n599 B.n597 10.6151
R1029 B.n600 B.n599 10.6151
R1030 B.n601 B.n600 10.6151
R1031 B.n602 B.n601 10.6151
R1032 B.n604 B.n602 10.6151
R1033 B.n605 B.n604 10.6151
R1034 B.n606 B.n605 10.6151
R1035 B.n607 B.n606 10.6151
R1036 B.n609 B.n607 10.6151
R1037 B.n610 B.n609 10.6151
R1038 B.n611 B.n610 10.6151
R1039 B.n612 B.n611 10.6151
R1040 B.n613 B.n612 10.6151
R1041 B.n669 B.n1 10.6151
R1042 B.n669 B.n668 10.6151
R1043 B.n668 B.n667 10.6151
R1044 B.n667 B.n10 10.6151
R1045 B.n661 B.n10 10.6151
R1046 B.n661 B.n660 10.6151
R1047 B.n660 B.n659 10.6151
R1048 B.n659 B.n18 10.6151
R1049 B.n653 B.n18 10.6151
R1050 B.n653 B.n652 10.6151
R1051 B.n652 B.n651 10.6151
R1052 B.n651 B.n24 10.6151
R1053 B.n645 B.n24 10.6151
R1054 B.n645 B.n644 10.6151
R1055 B.n644 B.n643 10.6151
R1056 B.n643 B.n32 10.6151
R1057 B.n637 B.n32 10.6151
R1058 B.n637 B.n636 10.6151
R1059 B.n636 B.n635 10.6151
R1060 B.n635 B.n39 10.6151
R1061 B.n629 B.n39 10.6151
R1062 B.n629 B.n628 10.6151
R1063 B.n628 B.n627 10.6151
R1064 B.n627 B.n46 10.6151
R1065 B.n621 B.n46 10.6151
R1066 B.n621 B.n620 10.6151
R1067 B.n619 B.n53 10.6151
R1068 B.n100 B.n53 10.6151
R1069 B.n101 B.n100 10.6151
R1070 B.n104 B.n101 10.6151
R1071 B.n105 B.n104 10.6151
R1072 B.n108 B.n105 10.6151
R1073 B.n109 B.n108 10.6151
R1074 B.n112 B.n109 10.6151
R1075 B.n113 B.n112 10.6151
R1076 B.n116 B.n113 10.6151
R1077 B.n117 B.n116 10.6151
R1078 B.n120 B.n117 10.6151
R1079 B.n121 B.n120 10.6151
R1080 B.n124 B.n121 10.6151
R1081 B.n125 B.n124 10.6151
R1082 B.n128 B.n125 10.6151
R1083 B.n129 B.n128 10.6151
R1084 B.n132 B.n129 10.6151
R1085 B.n133 B.n132 10.6151
R1086 B.n136 B.n133 10.6151
R1087 B.n137 B.n136 10.6151
R1088 B.n140 B.n137 10.6151
R1089 B.n141 B.n140 10.6151
R1090 B.n144 B.n141 10.6151
R1091 B.n145 B.n144 10.6151
R1092 B.n148 B.n145 10.6151
R1093 B.n149 B.n148 10.6151
R1094 B.n152 B.n149 10.6151
R1095 B.n153 B.n152 10.6151
R1096 B.n156 B.n153 10.6151
R1097 B.n157 B.n156 10.6151
R1098 B.n160 B.n157 10.6151
R1099 B.n161 B.n160 10.6151
R1100 B.n165 B.n164 10.6151
R1101 B.n168 B.n165 10.6151
R1102 B.n169 B.n168 10.6151
R1103 B.n172 B.n169 10.6151
R1104 B.n173 B.n172 10.6151
R1105 B.n176 B.n173 10.6151
R1106 B.n177 B.n176 10.6151
R1107 B.n180 B.n177 10.6151
R1108 B.n185 B.n182 10.6151
R1109 B.n186 B.n185 10.6151
R1110 B.n189 B.n186 10.6151
R1111 B.n190 B.n189 10.6151
R1112 B.n193 B.n190 10.6151
R1113 B.n194 B.n193 10.6151
R1114 B.n197 B.n194 10.6151
R1115 B.n198 B.n197 10.6151
R1116 B.n201 B.n198 10.6151
R1117 B.n202 B.n201 10.6151
R1118 B.n205 B.n202 10.6151
R1119 B.n206 B.n205 10.6151
R1120 B.n209 B.n206 10.6151
R1121 B.n210 B.n209 10.6151
R1122 B.n213 B.n210 10.6151
R1123 B.n214 B.n213 10.6151
R1124 B.n217 B.n214 10.6151
R1125 B.n218 B.n217 10.6151
R1126 B.n221 B.n218 10.6151
R1127 B.n222 B.n221 10.6151
R1128 B.n225 B.n222 10.6151
R1129 B.n226 B.n225 10.6151
R1130 B.n229 B.n226 10.6151
R1131 B.n230 B.n229 10.6151
R1132 B.n233 B.n230 10.6151
R1133 B.n234 B.n233 10.6151
R1134 B.n237 B.n234 10.6151
R1135 B.n238 B.n237 10.6151
R1136 B.n241 B.n238 10.6151
R1137 B.n242 B.n241 10.6151
R1138 B.n245 B.n242 10.6151
R1139 B.n246 B.n245 10.6151
R1140 B.n614 B.n246 10.6151
R1141 B.n677 B.n0 8.11757
R1142 B.n677 B.n1 8.11757
R1143 B.n429 B.n428 6.5566
R1144 B.n412 B.n342 6.5566
R1145 B.n164 B.n98 6.5566
R1146 B.n181 B.n180 6.5566
R1147 B.n430 B.n429 4.05904
R1148 B.n409 B.n342 4.05904
R1149 B.n161 B.n98 4.05904
R1150 B.n182 B.n181 4.05904
R1151 VN.n0 VN.t1 158.103
R1152 VN.n1 VN.t3 158.103
R1153 VN.n0 VN.t2 157.668
R1154 VN.n1 VN.t0 157.668
R1155 VN VN.n1 51.5373
R1156 VN VN.n0 9.19261
R1157 VDD2.n2 VDD2.n0 101.966
R1158 VDD2.n2 VDD2.n1 64.5534
R1159 VDD2.n1 VDD2.t3 2.12496
R1160 VDD2.n1 VDD2.t1 2.12496
R1161 VDD2.n0 VDD2.t0 2.12496
R1162 VDD2.n0 VDD2.t2 2.12496
R1163 VDD2 VDD2.n2 0.0586897
R1164 VTAIL.n394 VTAIL.n350 289.615
R1165 VTAIL.n44 VTAIL.n0 289.615
R1166 VTAIL.n94 VTAIL.n50 289.615
R1167 VTAIL.n144 VTAIL.n100 289.615
R1168 VTAIL.n344 VTAIL.n300 289.615
R1169 VTAIL.n294 VTAIL.n250 289.615
R1170 VTAIL.n244 VTAIL.n200 289.615
R1171 VTAIL.n194 VTAIL.n150 289.615
R1172 VTAIL.n367 VTAIL.n366 185
R1173 VTAIL.n369 VTAIL.n368 185
R1174 VTAIL.n362 VTAIL.n361 185
R1175 VTAIL.n375 VTAIL.n374 185
R1176 VTAIL.n377 VTAIL.n376 185
R1177 VTAIL.n358 VTAIL.n357 185
R1178 VTAIL.n384 VTAIL.n383 185
R1179 VTAIL.n385 VTAIL.n356 185
R1180 VTAIL.n387 VTAIL.n386 185
R1181 VTAIL.n354 VTAIL.n353 185
R1182 VTAIL.n393 VTAIL.n392 185
R1183 VTAIL.n395 VTAIL.n394 185
R1184 VTAIL.n17 VTAIL.n16 185
R1185 VTAIL.n19 VTAIL.n18 185
R1186 VTAIL.n12 VTAIL.n11 185
R1187 VTAIL.n25 VTAIL.n24 185
R1188 VTAIL.n27 VTAIL.n26 185
R1189 VTAIL.n8 VTAIL.n7 185
R1190 VTAIL.n34 VTAIL.n33 185
R1191 VTAIL.n35 VTAIL.n6 185
R1192 VTAIL.n37 VTAIL.n36 185
R1193 VTAIL.n4 VTAIL.n3 185
R1194 VTAIL.n43 VTAIL.n42 185
R1195 VTAIL.n45 VTAIL.n44 185
R1196 VTAIL.n67 VTAIL.n66 185
R1197 VTAIL.n69 VTAIL.n68 185
R1198 VTAIL.n62 VTAIL.n61 185
R1199 VTAIL.n75 VTAIL.n74 185
R1200 VTAIL.n77 VTAIL.n76 185
R1201 VTAIL.n58 VTAIL.n57 185
R1202 VTAIL.n84 VTAIL.n83 185
R1203 VTAIL.n85 VTAIL.n56 185
R1204 VTAIL.n87 VTAIL.n86 185
R1205 VTAIL.n54 VTAIL.n53 185
R1206 VTAIL.n93 VTAIL.n92 185
R1207 VTAIL.n95 VTAIL.n94 185
R1208 VTAIL.n117 VTAIL.n116 185
R1209 VTAIL.n119 VTAIL.n118 185
R1210 VTAIL.n112 VTAIL.n111 185
R1211 VTAIL.n125 VTAIL.n124 185
R1212 VTAIL.n127 VTAIL.n126 185
R1213 VTAIL.n108 VTAIL.n107 185
R1214 VTAIL.n134 VTAIL.n133 185
R1215 VTAIL.n135 VTAIL.n106 185
R1216 VTAIL.n137 VTAIL.n136 185
R1217 VTAIL.n104 VTAIL.n103 185
R1218 VTAIL.n143 VTAIL.n142 185
R1219 VTAIL.n145 VTAIL.n144 185
R1220 VTAIL.n345 VTAIL.n344 185
R1221 VTAIL.n343 VTAIL.n342 185
R1222 VTAIL.n304 VTAIL.n303 185
R1223 VTAIL.n308 VTAIL.n306 185
R1224 VTAIL.n337 VTAIL.n336 185
R1225 VTAIL.n335 VTAIL.n334 185
R1226 VTAIL.n310 VTAIL.n309 185
R1227 VTAIL.n329 VTAIL.n328 185
R1228 VTAIL.n327 VTAIL.n326 185
R1229 VTAIL.n314 VTAIL.n313 185
R1230 VTAIL.n321 VTAIL.n320 185
R1231 VTAIL.n319 VTAIL.n318 185
R1232 VTAIL.n295 VTAIL.n294 185
R1233 VTAIL.n293 VTAIL.n292 185
R1234 VTAIL.n254 VTAIL.n253 185
R1235 VTAIL.n258 VTAIL.n256 185
R1236 VTAIL.n287 VTAIL.n286 185
R1237 VTAIL.n285 VTAIL.n284 185
R1238 VTAIL.n260 VTAIL.n259 185
R1239 VTAIL.n279 VTAIL.n278 185
R1240 VTAIL.n277 VTAIL.n276 185
R1241 VTAIL.n264 VTAIL.n263 185
R1242 VTAIL.n271 VTAIL.n270 185
R1243 VTAIL.n269 VTAIL.n268 185
R1244 VTAIL.n245 VTAIL.n244 185
R1245 VTAIL.n243 VTAIL.n242 185
R1246 VTAIL.n204 VTAIL.n203 185
R1247 VTAIL.n208 VTAIL.n206 185
R1248 VTAIL.n237 VTAIL.n236 185
R1249 VTAIL.n235 VTAIL.n234 185
R1250 VTAIL.n210 VTAIL.n209 185
R1251 VTAIL.n229 VTAIL.n228 185
R1252 VTAIL.n227 VTAIL.n226 185
R1253 VTAIL.n214 VTAIL.n213 185
R1254 VTAIL.n221 VTAIL.n220 185
R1255 VTAIL.n219 VTAIL.n218 185
R1256 VTAIL.n195 VTAIL.n194 185
R1257 VTAIL.n193 VTAIL.n192 185
R1258 VTAIL.n154 VTAIL.n153 185
R1259 VTAIL.n158 VTAIL.n156 185
R1260 VTAIL.n187 VTAIL.n186 185
R1261 VTAIL.n185 VTAIL.n184 185
R1262 VTAIL.n160 VTAIL.n159 185
R1263 VTAIL.n179 VTAIL.n178 185
R1264 VTAIL.n177 VTAIL.n176 185
R1265 VTAIL.n164 VTAIL.n163 185
R1266 VTAIL.n171 VTAIL.n170 185
R1267 VTAIL.n169 VTAIL.n168 185
R1268 VTAIL.n365 VTAIL.t5 149.524
R1269 VTAIL.n15 VTAIL.t6 149.524
R1270 VTAIL.n65 VTAIL.t2 149.524
R1271 VTAIL.n115 VTAIL.t0 149.524
R1272 VTAIL.n317 VTAIL.t1 149.524
R1273 VTAIL.n267 VTAIL.t3 149.524
R1274 VTAIL.n217 VTAIL.t4 149.524
R1275 VTAIL.n167 VTAIL.t7 149.524
R1276 VTAIL.n368 VTAIL.n367 104.615
R1277 VTAIL.n368 VTAIL.n361 104.615
R1278 VTAIL.n375 VTAIL.n361 104.615
R1279 VTAIL.n376 VTAIL.n375 104.615
R1280 VTAIL.n376 VTAIL.n357 104.615
R1281 VTAIL.n384 VTAIL.n357 104.615
R1282 VTAIL.n385 VTAIL.n384 104.615
R1283 VTAIL.n386 VTAIL.n385 104.615
R1284 VTAIL.n386 VTAIL.n353 104.615
R1285 VTAIL.n393 VTAIL.n353 104.615
R1286 VTAIL.n394 VTAIL.n393 104.615
R1287 VTAIL.n18 VTAIL.n17 104.615
R1288 VTAIL.n18 VTAIL.n11 104.615
R1289 VTAIL.n25 VTAIL.n11 104.615
R1290 VTAIL.n26 VTAIL.n25 104.615
R1291 VTAIL.n26 VTAIL.n7 104.615
R1292 VTAIL.n34 VTAIL.n7 104.615
R1293 VTAIL.n35 VTAIL.n34 104.615
R1294 VTAIL.n36 VTAIL.n35 104.615
R1295 VTAIL.n36 VTAIL.n3 104.615
R1296 VTAIL.n43 VTAIL.n3 104.615
R1297 VTAIL.n44 VTAIL.n43 104.615
R1298 VTAIL.n68 VTAIL.n67 104.615
R1299 VTAIL.n68 VTAIL.n61 104.615
R1300 VTAIL.n75 VTAIL.n61 104.615
R1301 VTAIL.n76 VTAIL.n75 104.615
R1302 VTAIL.n76 VTAIL.n57 104.615
R1303 VTAIL.n84 VTAIL.n57 104.615
R1304 VTAIL.n85 VTAIL.n84 104.615
R1305 VTAIL.n86 VTAIL.n85 104.615
R1306 VTAIL.n86 VTAIL.n53 104.615
R1307 VTAIL.n93 VTAIL.n53 104.615
R1308 VTAIL.n94 VTAIL.n93 104.615
R1309 VTAIL.n118 VTAIL.n117 104.615
R1310 VTAIL.n118 VTAIL.n111 104.615
R1311 VTAIL.n125 VTAIL.n111 104.615
R1312 VTAIL.n126 VTAIL.n125 104.615
R1313 VTAIL.n126 VTAIL.n107 104.615
R1314 VTAIL.n134 VTAIL.n107 104.615
R1315 VTAIL.n135 VTAIL.n134 104.615
R1316 VTAIL.n136 VTAIL.n135 104.615
R1317 VTAIL.n136 VTAIL.n103 104.615
R1318 VTAIL.n143 VTAIL.n103 104.615
R1319 VTAIL.n144 VTAIL.n143 104.615
R1320 VTAIL.n344 VTAIL.n343 104.615
R1321 VTAIL.n343 VTAIL.n303 104.615
R1322 VTAIL.n308 VTAIL.n303 104.615
R1323 VTAIL.n336 VTAIL.n308 104.615
R1324 VTAIL.n336 VTAIL.n335 104.615
R1325 VTAIL.n335 VTAIL.n309 104.615
R1326 VTAIL.n328 VTAIL.n309 104.615
R1327 VTAIL.n328 VTAIL.n327 104.615
R1328 VTAIL.n327 VTAIL.n313 104.615
R1329 VTAIL.n320 VTAIL.n313 104.615
R1330 VTAIL.n320 VTAIL.n319 104.615
R1331 VTAIL.n294 VTAIL.n293 104.615
R1332 VTAIL.n293 VTAIL.n253 104.615
R1333 VTAIL.n258 VTAIL.n253 104.615
R1334 VTAIL.n286 VTAIL.n258 104.615
R1335 VTAIL.n286 VTAIL.n285 104.615
R1336 VTAIL.n285 VTAIL.n259 104.615
R1337 VTAIL.n278 VTAIL.n259 104.615
R1338 VTAIL.n278 VTAIL.n277 104.615
R1339 VTAIL.n277 VTAIL.n263 104.615
R1340 VTAIL.n270 VTAIL.n263 104.615
R1341 VTAIL.n270 VTAIL.n269 104.615
R1342 VTAIL.n244 VTAIL.n243 104.615
R1343 VTAIL.n243 VTAIL.n203 104.615
R1344 VTAIL.n208 VTAIL.n203 104.615
R1345 VTAIL.n236 VTAIL.n208 104.615
R1346 VTAIL.n236 VTAIL.n235 104.615
R1347 VTAIL.n235 VTAIL.n209 104.615
R1348 VTAIL.n228 VTAIL.n209 104.615
R1349 VTAIL.n228 VTAIL.n227 104.615
R1350 VTAIL.n227 VTAIL.n213 104.615
R1351 VTAIL.n220 VTAIL.n213 104.615
R1352 VTAIL.n220 VTAIL.n219 104.615
R1353 VTAIL.n194 VTAIL.n193 104.615
R1354 VTAIL.n193 VTAIL.n153 104.615
R1355 VTAIL.n158 VTAIL.n153 104.615
R1356 VTAIL.n186 VTAIL.n158 104.615
R1357 VTAIL.n186 VTAIL.n185 104.615
R1358 VTAIL.n185 VTAIL.n159 104.615
R1359 VTAIL.n178 VTAIL.n159 104.615
R1360 VTAIL.n178 VTAIL.n177 104.615
R1361 VTAIL.n177 VTAIL.n163 104.615
R1362 VTAIL.n170 VTAIL.n163 104.615
R1363 VTAIL.n170 VTAIL.n169 104.615
R1364 VTAIL.n367 VTAIL.t5 52.3082
R1365 VTAIL.n17 VTAIL.t6 52.3082
R1366 VTAIL.n67 VTAIL.t2 52.3082
R1367 VTAIL.n117 VTAIL.t0 52.3082
R1368 VTAIL.n319 VTAIL.t1 52.3082
R1369 VTAIL.n269 VTAIL.t3 52.3082
R1370 VTAIL.n219 VTAIL.t4 52.3082
R1371 VTAIL.n169 VTAIL.t7 52.3082
R1372 VTAIL.n399 VTAIL.n398 33.7369
R1373 VTAIL.n49 VTAIL.n48 33.7369
R1374 VTAIL.n99 VTAIL.n98 33.7369
R1375 VTAIL.n149 VTAIL.n148 33.7369
R1376 VTAIL.n349 VTAIL.n348 33.7369
R1377 VTAIL.n299 VTAIL.n298 33.7369
R1378 VTAIL.n249 VTAIL.n248 33.7369
R1379 VTAIL.n199 VTAIL.n198 33.7369
R1380 VTAIL.n399 VTAIL.n349 22.2893
R1381 VTAIL.n199 VTAIL.n149 22.2893
R1382 VTAIL.n387 VTAIL.n354 13.1884
R1383 VTAIL.n37 VTAIL.n4 13.1884
R1384 VTAIL.n87 VTAIL.n54 13.1884
R1385 VTAIL.n137 VTAIL.n104 13.1884
R1386 VTAIL.n306 VTAIL.n304 13.1884
R1387 VTAIL.n256 VTAIL.n254 13.1884
R1388 VTAIL.n206 VTAIL.n204 13.1884
R1389 VTAIL.n156 VTAIL.n154 13.1884
R1390 VTAIL.n388 VTAIL.n356 12.8005
R1391 VTAIL.n392 VTAIL.n391 12.8005
R1392 VTAIL.n38 VTAIL.n6 12.8005
R1393 VTAIL.n42 VTAIL.n41 12.8005
R1394 VTAIL.n88 VTAIL.n56 12.8005
R1395 VTAIL.n92 VTAIL.n91 12.8005
R1396 VTAIL.n138 VTAIL.n106 12.8005
R1397 VTAIL.n142 VTAIL.n141 12.8005
R1398 VTAIL.n342 VTAIL.n341 12.8005
R1399 VTAIL.n338 VTAIL.n337 12.8005
R1400 VTAIL.n292 VTAIL.n291 12.8005
R1401 VTAIL.n288 VTAIL.n287 12.8005
R1402 VTAIL.n242 VTAIL.n241 12.8005
R1403 VTAIL.n238 VTAIL.n237 12.8005
R1404 VTAIL.n192 VTAIL.n191 12.8005
R1405 VTAIL.n188 VTAIL.n187 12.8005
R1406 VTAIL.n383 VTAIL.n382 12.0247
R1407 VTAIL.n395 VTAIL.n352 12.0247
R1408 VTAIL.n33 VTAIL.n32 12.0247
R1409 VTAIL.n45 VTAIL.n2 12.0247
R1410 VTAIL.n83 VTAIL.n82 12.0247
R1411 VTAIL.n95 VTAIL.n52 12.0247
R1412 VTAIL.n133 VTAIL.n132 12.0247
R1413 VTAIL.n145 VTAIL.n102 12.0247
R1414 VTAIL.n345 VTAIL.n302 12.0247
R1415 VTAIL.n334 VTAIL.n307 12.0247
R1416 VTAIL.n295 VTAIL.n252 12.0247
R1417 VTAIL.n284 VTAIL.n257 12.0247
R1418 VTAIL.n245 VTAIL.n202 12.0247
R1419 VTAIL.n234 VTAIL.n207 12.0247
R1420 VTAIL.n195 VTAIL.n152 12.0247
R1421 VTAIL.n184 VTAIL.n157 12.0247
R1422 VTAIL.n381 VTAIL.n358 11.249
R1423 VTAIL.n396 VTAIL.n350 11.249
R1424 VTAIL.n31 VTAIL.n8 11.249
R1425 VTAIL.n46 VTAIL.n0 11.249
R1426 VTAIL.n81 VTAIL.n58 11.249
R1427 VTAIL.n96 VTAIL.n50 11.249
R1428 VTAIL.n131 VTAIL.n108 11.249
R1429 VTAIL.n146 VTAIL.n100 11.249
R1430 VTAIL.n346 VTAIL.n300 11.249
R1431 VTAIL.n333 VTAIL.n310 11.249
R1432 VTAIL.n296 VTAIL.n250 11.249
R1433 VTAIL.n283 VTAIL.n260 11.249
R1434 VTAIL.n246 VTAIL.n200 11.249
R1435 VTAIL.n233 VTAIL.n210 11.249
R1436 VTAIL.n196 VTAIL.n150 11.249
R1437 VTAIL.n183 VTAIL.n160 11.249
R1438 VTAIL.n378 VTAIL.n377 10.4732
R1439 VTAIL.n28 VTAIL.n27 10.4732
R1440 VTAIL.n78 VTAIL.n77 10.4732
R1441 VTAIL.n128 VTAIL.n127 10.4732
R1442 VTAIL.n330 VTAIL.n329 10.4732
R1443 VTAIL.n280 VTAIL.n279 10.4732
R1444 VTAIL.n230 VTAIL.n229 10.4732
R1445 VTAIL.n180 VTAIL.n179 10.4732
R1446 VTAIL.n366 VTAIL.n365 10.2747
R1447 VTAIL.n16 VTAIL.n15 10.2747
R1448 VTAIL.n66 VTAIL.n65 10.2747
R1449 VTAIL.n116 VTAIL.n115 10.2747
R1450 VTAIL.n318 VTAIL.n317 10.2747
R1451 VTAIL.n268 VTAIL.n267 10.2747
R1452 VTAIL.n218 VTAIL.n217 10.2747
R1453 VTAIL.n168 VTAIL.n167 10.2747
R1454 VTAIL.n374 VTAIL.n360 9.69747
R1455 VTAIL.n24 VTAIL.n10 9.69747
R1456 VTAIL.n74 VTAIL.n60 9.69747
R1457 VTAIL.n124 VTAIL.n110 9.69747
R1458 VTAIL.n326 VTAIL.n312 9.69747
R1459 VTAIL.n276 VTAIL.n262 9.69747
R1460 VTAIL.n226 VTAIL.n212 9.69747
R1461 VTAIL.n176 VTAIL.n162 9.69747
R1462 VTAIL.n398 VTAIL.n397 9.45567
R1463 VTAIL.n48 VTAIL.n47 9.45567
R1464 VTAIL.n98 VTAIL.n97 9.45567
R1465 VTAIL.n148 VTAIL.n147 9.45567
R1466 VTAIL.n348 VTAIL.n347 9.45567
R1467 VTAIL.n298 VTAIL.n297 9.45567
R1468 VTAIL.n248 VTAIL.n247 9.45567
R1469 VTAIL.n198 VTAIL.n197 9.45567
R1470 VTAIL.n397 VTAIL.n396 9.3005
R1471 VTAIL.n352 VTAIL.n351 9.3005
R1472 VTAIL.n391 VTAIL.n390 9.3005
R1473 VTAIL.n364 VTAIL.n363 9.3005
R1474 VTAIL.n371 VTAIL.n370 9.3005
R1475 VTAIL.n373 VTAIL.n372 9.3005
R1476 VTAIL.n360 VTAIL.n359 9.3005
R1477 VTAIL.n379 VTAIL.n378 9.3005
R1478 VTAIL.n381 VTAIL.n380 9.3005
R1479 VTAIL.n382 VTAIL.n355 9.3005
R1480 VTAIL.n389 VTAIL.n388 9.3005
R1481 VTAIL.n47 VTAIL.n46 9.3005
R1482 VTAIL.n2 VTAIL.n1 9.3005
R1483 VTAIL.n41 VTAIL.n40 9.3005
R1484 VTAIL.n14 VTAIL.n13 9.3005
R1485 VTAIL.n21 VTAIL.n20 9.3005
R1486 VTAIL.n23 VTAIL.n22 9.3005
R1487 VTAIL.n10 VTAIL.n9 9.3005
R1488 VTAIL.n29 VTAIL.n28 9.3005
R1489 VTAIL.n31 VTAIL.n30 9.3005
R1490 VTAIL.n32 VTAIL.n5 9.3005
R1491 VTAIL.n39 VTAIL.n38 9.3005
R1492 VTAIL.n97 VTAIL.n96 9.3005
R1493 VTAIL.n52 VTAIL.n51 9.3005
R1494 VTAIL.n91 VTAIL.n90 9.3005
R1495 VTAIL.n64 VTAIL.n63 9.3005
R1496 VTAIL.n71 VTAIL.n70 9.3005
R1497 VTAIL.n73 VTAIL.n72 9.3005
R1498 VTAIL.n60 VTAIL.n59 9.3005
R1499 VTAIL.n79 VTAIL.n78 9.3005
R1500 VTAIL.n81 VTAIL.n80 9.3005
R1501 VTAIL.n82 VTAIL.n55 9.3005
R1502 VTAIL.n89 VTAIL.n88 9.3005
R1503 VTAIL.n147 VTAIL.n146 9.3005
R1504 VTAIL.n102 VTAIL.n101 9.3005
R1505 VTAIL.n141 VTAIL.n140 9.3005
R1506 VTAIL.n114 VTAIL.n113 9.3005
R1507 VTAIL.n121 VTAIL.n120 9.3005
R1508 VTAIL.n123 VTAIL.n122 9.3005
R1509 VTAIL.n110 VTAIL.n109 9.3005
R1510 VTAIL.n129 VTAIL.n128 9.3005
R1511 VTAIL.n131 VTAIL.n130 9.3005
R1512 VTAIL.n132 VTAIL.n105 9.3005
R1513 VTAIL.n139 VTAIL.n138 9.3005
R1514 VTAIL.n316 VTAIL.n315 9.3005
R1515 VTAIL.n323 VTAIL.n322 9.3005
R1516 VTAIL.n325 VTAIL.n324 9.3005
R1517 VTAIL.n312 VTAIL.n311 9.3005
R1518 VTAIL.n331 VTAIL.n330 9.3005
R1519 VTAIL.n333 VTAIL.n332 9.3005
R1520 VTAIL.n307 VTAIL.n305 9.3005
R1521 VTAIL.n339 VTAIL.n338 9.3005
R1522 VTAIL.n347 VTAIL.n346 9.3005
R1523 VTAIL.n302 VTAIL.n301 9.3005
R1524 VTAIL.n341 VTAIL.n340 9.3005
R1525 VTAIL.n266 VTAIL.n265 9.3005
R1526 VTAIL.n273 VTAIL.n272 9.3005
R1527 VTAIL.n275 VTAIL.n274 9.3005
R1528 VTAIL.n262 VTAIL.n261 9.3005
R1529 VTAIL.n281 VTAIL.n280 9.3005
R1530 VTAIL.n283 VTAIL.n282 9.3005
R1531 VTAIL.n257 VTAIL.n255 9.3005
R1532 VTAIL.n289 VTAIL.n288 9.3005
R1533 VTAIL.n297 VTAIL.n296 9.3005
R1534 VTAIL.n252 VTAIL.n251 9.3005
R1535 VTAIL.n291 VTAIL.n290 9.3005
R1536 VTAIL.n216 VTAIL.n215 9.3005
R1537 VTAIL.n223 VTAIL.n222 9.3005
R1538 VTAIL.n225 VTAIL.n224 9.3005
R1539 VTAIL.n212 VTAIL.n211 9.3005
R1540 VTAIL.n231 VTAIL.n230 9.3005
R1541 VTAIL.n233 VTAIL.n232 9.3005
R1542 VTAIL.n207 VTAIL.n205 9.3005
R1543 VTAIL.n239 VTAIL.n238 9.3005
R1544 VTAIL.n247 VTAIL.n246 9.3005
R1545 VTAIL.n202 VTAIL.n201 9.3005
R1546 VTAIL.n241 VTAIL.n240 9.3005
R1547 VTAIL.n166 VTAIL.n165 9.3005
R1548 VTAIL.n173 VTAIL.n172 9.3005
R1549 VTAIL.n175 VTAIL.n174 9.3005
R1550 VTAIL.n162 VTAIL.n161 9.3005
R1551 VTAIL.n181 VTAIL.n180 9.3005
R1552 VTAIL.n183 VTAIL.n182 9.3005
R1553 VTAIL.n157 VTAIL.n155 9.3005
R1554 VTAIL.n189 VTAIL.n188 9.3005
R1555 VTAIL.n197 VTAIL.n196 9.3005
R1556 VTAIL.n152 VTAIL.n151 9.3005
R1557 VTAIL.n191 VTAIL.n190 9.3005
R1558 VTAIL.n373 VTAIL.n362 8.92171
R1559 VTAIL.n23 VTAIL.n12 8.92171
R1560 VTAIL.n73 VTAIL.n62 8.92171
R1561 VTAIL.n123 VTAIL.n112 8.92171
R1562 VTAIL.n325 VTAIL.n314 8.92171
R1563 VTAIL.n275 VTAIL.n264 8.92171
R1564 VTAIL.n225 VTAIL.n214 8.92171
R1565 VTAIL.n175 VTAIL.n164 8.92171
R1566 VTAIL.n370 VTAIL.n369 8.14595
R1567 VTAIL.n20 VTAIL.n19 8.14595
R1568 VTAIL.n70 VTAIL.n69 8.14595
R1569 VTAIL.n120 VTAIL.n119 8.14595
R1570 VTAIL.n322 VTAIL.n321 8.14595
R1571 VTAIL.n272 VTAIL.n271 8.14595
R1572 VTAIL.n222 VTAIL.n221 8.14595
R1573 VTAIL.n172 VTAIL.n171 8.14595
R1574 VTAIL.n366 VTAIL.n364 7.3702
R1575 VTAIL.n16 VTAIL.n14 7.3702
R1576 VTAIL.n66 VTAIL.n64 7.3702
R1577 VTAIL.n116 VTAIL.n114 7.3702
R1578 VTAIL.n318 VTAIL.n316 7.3702
R1579 VTAIL.n268 VTAIL.n266 7.3702
R1580 VTAIL.n218 VTAIL.n216 7.3702
R1581 VTAIL.n168 VTAIL.n166 7.3702
R1582 VTAIL.n369 VTAIL.n364 5.81868
R1583 VTAIL.n19 VTAIL.n14 5.81868
R1584 VTAIL.n69 VTAIL.n64 5.81868
R1585 VTAIL.n119 VTAIL.n114 5.81868
R1586 VTAIL.n321 VTAIL.n316 5.81868
R1587 VTAIL.n271 VTAIL.n266 5.81868
R1588 VTAIL.n221 VTAIL.n216 5.81868
R1589 VTAIL.n171 VTAIL.n166 5.81868
R1590 VTAIL.n370 VTAIL.n362 5.04292
R1591 VTAIL.n20 VTAIL.n12 5.04292
R1592 VTAIL.n70 VTAIL.n62 5.04292
R1593 VTAIL.n120 VTAIL.n112 5.04292
R1594 VTAIL.n322 VTAIL.n314 5.04292
R1595 VTAIL.n272 VTAIL.n264 5.04292
R1596 VTAIL.n222 VTAIL.n214 5.04292
R1597 VTAIL.n172 VTAIL.n164 5.04292
R1598 VTAIL.n374 VTAIL.n373 4.26717
R1599 VTAIL.n24 VTAIL.n23 4.26717
R1600 VTAIL.n74 VTAIL.n73 4.26717
R1601 VTAIL.n124 VTAIL.n123 4.26717
R1602 VTAIL.n326 VTAIL.n325 4.26717
R1603 VTAIL.n276 VTAIL.n275 4.26717
R1604 VTAIL.n226 VTAIL.n225 4.26717
R1605 VTAIL.n176 VTAIL.n175 4.26717
R1606 VTAIL.n377 VTAIL.n360 3.49141
R1607 VTAIL.n27 VTAIL.n10 3.49141
R1608 VTAIL.n77 VTAIL.n60 3.49141
R1609 VTAIL.n127 VTAIL.n110 3.49141
R1610 VTAIL.n329 VTAIL.n312 3.49141
R1611 VTAIL.n279 VTAIL.n262 3.49141
R1612 VTAIL.n229 VTAIL.n212 3.49141
R1613 VTAIL.n179 VTAIL.n162 3.49141
R1614 VTAIL.n365 VTAIL.n363 2.84303
R1615 VTAIL.n15 VTAIL.n13 2.84303
R1616 VTAIL.n65 VTAIL.n63 2.84303
R1617 VTAIL.n115 VTAIL.n113 2.84303
R1618 VTAIL.n317 VTAIL.n315 2.84303
R1619 VTAIL.n267 VTAIL.n265 2.84303
R1620 VTAIL.n217 VTAIL.n215 2.84303
R1621 VTAIL.n167 VTAIL.n165 2.84303
R1622 VTAIL.n378 VTAIL.n358 2.71565
R1623 VTAIL.n398 VTAIL.n350 2.71565
R1624 VTAIL.n28 VTAIL.n8 2.71565
R1625 VTAIL.n48 VTAIL.n0 2.71565
R1626 VTAIL.n78 VTAIL.n58 2.71565
R1627 VTAIL.n98 VTAIL.n50 2.71565
R1628 VTAIL.n128 VTAIL.n108 2.71565
R1629 VTAIL.n148 VTAIL.n100 2.71565
R1630 VTAIL.n348 VTAIL.n300 2.71565
R1631 VTAIL.n330 VTAIL.n310 2.71565
R1632 VTAIL.n298 VTAIL.n250 2.71565
R1633 VTAIL.n280 VTAIL.n260 2.71565
R1634 VTAIL.n248 VTAIL.n200 2.71565
R1635 VTAIL.n230 VTAIL.n210 2.71565
R1636 VTAIL.n198 VTAIL.n150 2.71565
R1637 VTAIL.n180 VTAIL.n160 2.71565
R1638 VTAIL.n383 VTAIL.n381 1.93989
R1639 VTAIL.n396 VTAIL.n395 1.93989
R1640 VTAIL.n33 VTAIL.n31 1.93989
R1641 VTAIL.n46 VTAIL.n45 1.93989
R1642 VTAIL.n83 VTAIL.n81 1.93989
R1643 VTAIL.n96 VTAIL.n95 1.93989
R1644 VTAIL.n133 VTAIL.n131 1.93989
R1645 VTAIL.n146 VTAIL.n145 1.93989
R1646 VTAIL.n346 VTAIL.n345 1.93989
R1647 VTAIL.n334 VTAIL.n333 1.93989
R1648 VTAIL.n296 VTAIL.n295 1.93989
R1649 VTAIL.n284 VTAIL.n283 1.93989
R1650 VTAIL.n246 VTAIL.n245 1.93989
R1651 VTAIL.n234 VTAIL.n233 1.93989
R1652 VTAIL.n196 VTAIL.n195 1.93989
R1653 VTAIL.n184 VTAIL.n183 1.93989
R1654 VTAIL.n249 VTAIL.n199 1.88843
R1655 VTAIL.n349 VTAIL.n299 1.88843
R1656 VTAIL.n149 VTAIL.n99 1.88843
R1657 VTAIL.n382 VTAIL.n356 1.16414
R1658 VTAIL.n392 VTAIL.n352 1.16414
R1659 VTAIL.n32 VTAIL.n6 1.16414
R1660 VTAIL.n42 VTAIL.n2 1.16414
R1661 VTAIL.n82 VTAIL.n56 1.16414
R1662 VTAIL.n92 VTAIL.n52 1.16414
R1663 VTAIL.n132 VTAIL.n106 1.16414
R1664 VTAIL.n142 VTAIL.n102 1.16414
R1665 VTAIL.n342 VTAIL.n302 1.16414
R1666 VTAIL.n337 VTAIL.n307 1.16414
R1667 VTAIL.n292 VTAIL.n252 1.16414
R1668 VTAIL.n287 VTAIL.n257 1.16414
R1669 VTAIL.n242 VTAIL.n202 1.16414
R1670 VTAIL.n237 VTAIL.n207 1.16414
R1671 VTAIL.n192 VTAIL.n152 1.16414
R1672 VTAIL.n187 VTAIL.n157 1.16414
R1673 VTAIL VTAIL.n49 1.00266
R1674 VTAIL VTAIL.n399 0.886276
R1675 VTAIL.n299 VTAIL.n249 0.470328
R1676 VTAIL.n99 VTAIL.n49 0.470328
R1677 VTAIL.n388 VTAIL.n387 0.388379
R1678 VTAIL.n391 VTAIL.n354 0.388379
R1679 VTAIL.n38 VTAIL.n37 0.388379
R1680 VTAIL.n41 VTAIL.n4 0.388379
R1681 VTAIL.n88 VTAIL.n87 0.388379
R1682 VTAIL.n91 VTAIL.n54 0.388379
R1683 VTAIL.n138 VTAIL.n137 0.388379
R1684 VTAIL.n141 VTAIL.n104 0.388379
R1685 VTAIL.n341 VTAIL.n304 0.388379
R1686 VTAIL.n338 VTAIL.n306 0.388379
R1687 VTAIL.n291 VTAIL.n254 0.388379
R1688 VTAIL.n288 VTAIL.n256 0.388379
R1689 VTAIL.n241 VTAIL.n204 0.388379
R1690 VTAIL.n238 VTAIL.n206 0.388379
R1691 VTAIL.n191 VTAIL.n154 0.388379
R1692 VTAIL.n188 VTAIL.n156 0.388379
R1693 VTAIL.n371 VTAIL.n363 0.155672
R1694 VTAIL.n372 VTAIL.n371 0.155672
R1695 VTAIL.n372 VTAIL.n359 0.155672
R1696 VTAIL.n379 VTAIL.n359 0.155672
R1697 VTAIL.n380 VTAIL.n379 0.155672
R1698 VTAIL.n380 VTAIL.n355 0.155672
R1699 VTAIL.n389 VTAIL.n355 0.155672
R1700 VTAIL.n390 VTAIL.n389 0.155672
R1701 VTAIL.n390 VTAIL.n351 0.155672
R1702 VTAIL.n397 VTAIL.n351 0.155672
R1703 VTAIL.n21 VTAIL.n13 0.155672
R1704 VTAIL.n22 VTAIL.n21 0.155672
R1705 VTAIL.n22 VTAIL.n9 0.155672
R1706 VTAIL.n29 VTAIL.n9 0.155672
R1707 VTAIL.n30 VTAIL.n29 0.155672
R1708 VTAIL.n30 VTAIL.n5 0.155672
R1709 VTAIL.n39 VTAIL.n5 0.155672
R1710 VTAIL.n40 VTAIL.n39 0.155672
R1711 VTAIL.n40 VTAIL.n1 0.155672
R1712 VTAIL.n47 VTAIL.n1 0.155672
R1713 VTAIL.n71 VTAIL.n63 0.155672
R1714 VTAIL.n72 VTAIL.n71 0.155672
R1715 VTAIL.n72 VTAIL.n59 0.155672
R1716 VTAIL.n79 VTAIL.n59 0.155672
R1717 VTAIL.n80 VTAIL.n79 0.155672
R1718 VTAIL.n80 VTAIL.n55 0.155672
R1719 VTAIL.n89 VTAIL.n55 0.155672
R1720 VTAIL.n90 VTAIL.n89 0.155672
R1721 VTAIL.n90 VTAIL.n51 0.155672
R1722 VTAIL.n97 VTAIL.n51 0.155672
R1723 VTAIL.n121 VTAIL.n113 0.155672
R1724 VTAIL.n122 VTAIL.n121 0.155672
R1725 VTAIL.n122 VTAIL.n109 0.155672
R1726 VTAIL.n129 VTAIL.n109 0.155672
R1727 VTAIL.n130 VTAIL.n129 0.155672
R1728 VTAIL.n130 VTAIL.n105 0.155672
R1729 VTAIL.n139 VTAIL.n105 0.155672
R1730 VTAIL.n140 VTAIL.n139 0.155672
R1731 VTAIL.n140 VTAIL.n101 0.155672
R1732 VTAIL.n147 VTAIL.n101 0.155672
R1733 VTAIL.n347 VTAIL.n301 0.155672
R1734 VTAIL.n340 VTAIL.n301 0.155672
R1735 VTAIL.n340 VTAIL.n339 0.155672
R1736 VTAIL.n339 VTAIL.n305 0.155672
R1737 VTAIL.n332 VTAIL.n305 0.155672
R1738 VTAIL.n332 VTAIL.n331 0.155672
R1739 VTAIL.n331 VTAIL.n311 0.155672
R1740 VTAIL.n324 VTAIL.n311 0.155672
R1741 VTAIL.n324 VTAIL.n323 0.155672
R1742 VTAIL.n323 VTAIL.n315 0.155672
R1743 VTAIL.n297 VTAIL.n251 0.155672
R1744 VTAIL.n290 VTAIL.n251 0.155672
R1745 VTAIL.n290 VTAIL.n289 0.155672
R1746 VTAIL.n289 VTAIL.n255 0.155672
R1747 VTAIL.n282 VTAIL.n255 0.155672
R1748 VTAIL.n282 VTAIL.n281 0.155672
R1749 VTAIL.n281 VTAIL.n261 0.155672
R1750 VTAIL.n274 VTAIL.n261 0.155672
R1751 VTAIL.n274 VTAIL.n273 0.155672
R1752 VTAIL.n273 VTAIL.n265 0.155672
R1753 VTAIL.n247 VTAIL.n201 0.155672
R1754 VTAIL.n240 VTAIL.n201 0.155672
R1755 VTAIL.n240 VTAIL.n239 0.155672
R1756 VTAIL.n239 VTAIL.n205 0.155672
R1757 VTAIL.n232 VTAIL.n205 0.155672
R1758 VTAIL.n232 VTAIL.n231 0.155672
R1759 VTAIL.n231 VTAIL.n211 0.155672
R1760 VTAIL.n224 VTAIL.n211 0.155672
R1761 VTAIL.n224 VTAIL.n223 0.155672
R1762 VTAIL.n223 VTAIL.n215 0.155672
R1763 VTAIL.n197 VTAIL.n151 0.155672
R1764 VTAIL.n190 VTAIL.n151 0.155672
R1765 VTAIL.n190 VTAIL.n189 0.155672
R1766 VTAIL.n189 VTAIL.n155 0.155672
R1767 VTAIL.n182 VTAIL.n155 0.155672
R1768 VTAIL.n182 VTAIL.n181 0.155672
R1769 VTAIL.n181 VTAIL.n161 0.155672
R1770 VTAIL.n174 VTAIL.n161 0.155672
R1771 VTAIL.n174 VTAIL.n173 0.155672
R1772 VTAIL.n173 VTAIL.n165 0.155672
R1773 VP.n5 VP.n4 181.018
R1774 VP.n14 VP.n13 181.018
R1775 VP.n12 VP.n0 161.3
R1776 VP.n11 VP.n10 161.3
R1777 VP.n9 VP.n1 161.3
R1778 VP.n8 VP.n7 161.3
R1779 VP.n6 VP.n2 161.3
R1780 VP.n3 VP.t1 158.103
R1781 VP.n3 VP.t3 157.668
R1782 VP.n5 VP.t2 120.76
R1783 VP.n13 VP.t0 120.76
R1784 VP.n4 VP.n3 51.1566
R1785 VP.n7 VP.n1 40.4106
R1786 VP.n11 VP.n1 40.4106
R1787 VP.n7 VP.n6 24.3439
R1788 VP.n12 VP.n11 24.3439
R1789 VP.n6 VP.n5 4.62575
R1790 VP.n13 VP.n12 4.62575
R1791 VP.n4 VP.n2 0.189894
R1792 VP.n8 VP.n2 0.189894
R1793 VP.n9 VP.n8 0.189894
R1794 VP.n10 VP.n9 0.189894
R1795 VP.n10 VP.n0 0.189894
R1796 VP.n14 VP.n0 0.189894
R1797 VP VP.n14 0.0516364
R1798 VDD1 VDD1.n1 102.492
R1799 VDD1 VDD1.n0 64.6116
R1800 VDD1.n0 VDD1.t2 2.12496
R1801 VDD1.n0 VDD1.t0 2.12496
R1802 VDD1.n1 VDD1.t1 2.12496
R1803 VDD1.n1 VDD1.t3 2.12496
C0 VTAIL VDD1 4.67046f
C1 VDD1 VDD2 0.846722f
C2 VP VN 5.16236f
C3 VTAIL VN 3.42951f
C4 VN VDD2 3.51183f
C5 VN VDD1 0.14782f
C6 VTAIL VP 3.44362f
C7 VP VDD2 0.346706f
C8 VP VDD1 3.71017f
C9 VTAIL VDD2 4.71971f
C10 VDD2 B 3.136959f
C11 VDD1 B 6.750741f
C12 VTAIL B 8.049464f
C13 VN B 9.13375f
C14 VP B 7.164778f
C15 VDD1.t2 B 0.199405f
C16 VDD1.t0 B 0.199405f
C17 VDD1.n0 B 1.74851f
C18 VDD1.t1 B 0.199405f
C19 VDD1.t3 B 0.199405f
C20 VDD1.n1 B 2.30699f
C21 VP.n0 B 0.03263f
C22 VP.t0 B 1.52851f
C23 VP.n1 B 0.026405f
C24 VP.n2 B 0.03263f
C25 VP.t2 B 1.52851f
C26 VP.t1 B 1.69934f
C27 VP.t3 B 1.69736f
C28 VP.n3 B 2.45935f
C29 VP.n4 B 1.66525f
C30 VP.n5 B 0.63751f
C31 VP.n6 B 0.036676f
C32 VP.n7 B 0.065198f
C33 VP.n8 B 0.03263f
C34 VP.n9 B 0.03263f
C35 VP.n10 B 0.03263f
C36 VP.n11 B 0.065198f
C37 VP.n12 B 0.036676f
C38 VP.n13 B 0.63751f
C39 VP.n14 B 0.034936f
C40 VTAIL.n0 B 0.022626f
C41 VTAIL.n1 B 0.01674f
C42 VTAIL.n2 B 0.008995f
C43 VTAIL.n3 B 0.021262f
C44 VTAIL.n4 B 0.00926f
C45 VTAIL.n5 B 0.01674f
C46 VTAIL.n6 B 0.009524f
C47 VTAIL.n7 B 0.021262f
C48 VTAIL.n8 B 0.009524f
C49 VTAIL.n9 B 0.01674f
C50 VTAIL.n10 B 0.008995f
C51 VTAIL.n11 B 0.021262f
C52 VTAIL.n12 B 0.009524f
C53 VTAIL.n13 B 0.644947f
C54 VTAIL.n14 B 0.008995f
C55 VTAIL.t6 B 0.035671f
C56 VTAIL.n15 B 0.103474f
C57 VTAIL.n16 B 0.01503f
C58 VTAIL.n17 B 0.015946f
C59 VTAIL.n18 B 0.021262f
C60 VTAIL.n19 B 0.009524f
C61 VTAIL.n20 B 0.008995f
C62 VTAIL.n21 B 0.01674f
C63 VTAIL.n22 B 0.01674f
C64 VTAIL.n23 B 0.008995f
C65 VTAIL.n24 B 0.009524f
C66 VTAIL.n25 B 0.021262f
C67 VTAIL.n26 B 0.021262f
C68 VTAIL.n27 B 0.009524f
C69 VTAIL.n28 B 0.008995f
C70 VTAIL.n29 B 0.01674f
C71 VTAIL.n30 B 0.01674f
C72 VTAIL.n31 B 0.008995f
C73 VTAIL.n32 B 0.008995f
C74 VTAIL.n33 B 0.009524f
C75 VTAIL.n34 B 0.021262f
C76 VTAIL.n35 B 0.021262f
C77 VTAIL.n36 B 0.021262f
C78 VTAIL.n37 B 0.00926f
C79 VTAIL.n38 B 0.008995f
C80 VTAIL.n39 B 0.01674f
C81 VTAIL.n40 B 0.01674f
C82 VTAIL.n41 B 0.008995f
C83 VTAIL.n42 B 0.009524f
C84 VTAIL.n43 B 0.021262f
C85 VTAIL.n44 B 0.04443f
C86 VTAIL.n45 B 0.009524f
C87 VTAIL.n46 B 0.008995f
C88 VTAIL.n47 B 0.040523f
C89 VTAIL.n48 B 0.024751f
C90 VTAIL.n49 B 0.094729f
C91 VTAIL.n50 B 0.022626f
C92 VTAIL.n51 B 0.01674f
C93 VTAIL.n52 B 0.008995f
C94 VTAIL.n53 B 0.021262f
C95 VTAIL.n54 B 0.00926f
C96 VTAIL.n55 B 0.01674f
C97 VTAIL.n56 B 0.009524f
C98 VTAIL.n57 B 0.021262f
C99 VTAIL.n58 B 0.009524f
C100 VTAIL.n59 B 0.01674f
C101 VTAIL.n60 B 0.008995f
C102 VTAIL.n61 B 0.021262f
C103 VTAIL.n62 B 0.009524f
C104 VTAIL.n63 B 0.644947f
C105 VTAIL.n64 B 0.008995f
C106 VTAIL.t2 B 0.035671f
C107 VTAIL.n65 B 0.103474f
C108 VTAIL.n66 B 0.01503f
C109 VTAIL.n67 B 0.015946f
C110 VTAIL.n68 B 0.021262f
C111 VTAIL.n69 B 0.009524f
C112 VTAIL.n70 B 0.008995f
C113 VTAIL.n71 B 0.01674f
C114 VTAIL.n72 B 0.01674f
C115 VTAIL.n73 B 0.008995f
C116 VTAIL.n74 B 0.009524f
C117 VTAIL.n75 B 0.021262f
C118 VTAIL.n76 B 0.021262f
C119 VTAIL.n77 B 0.009524f
C120 VTAIL.n78 B 0.008995f
C121 VTAIL.n79 B 0.01674f
C122 VTAIL.n80 B 0.01674f
C123 VTAIL.n81 B 0.008995f
C124 VTAIL.n82 B 0.008995f
C125 VTAIL.n83 B 0.009524f
C126 VTAIL.n84 B 0.021262f
C127 VTAIL.n85 B 0.021262f
C128 VTAIL.n86 B 0.021262f
C129 VTAIL.n87 B 0.00926f
C130 VTAIL.n88 B 0.008995f
C131 VTAIL.n89 B 0.01674f
C132 VTAIL.n90 B 0.01674f
C133 VTAIL.n91 B 0.008995f
C134 VTAIL.n92 B 0.009524f
C135 VTAIL.n93 B 0.021262f
C136 VTAIL.n94 B 0.04443f
C137 VTAIL.n95 B 0.009524f
C138 VTAIL.n96 B 0.008995f
C139 VTAIL.n97 B 0.040523f
C140 VTAIL.n98 B 0.024751f
C141 VTAIL.n99 B 0.142508f
C142 VTAIL.n100 B 0.022626f
C143 VTAIL.n101 B 0.01674f
C144 VTAIL.n102 B 0.008995f
C145 VTAIL.n103 B 0.021262f
C146 VTAIL.n104 B 0.00926f
C147 VTAIL.n105 B 0.01674f
C148 VTAIL.n106 B 0.009524f
C149 VTAIL.n107 B 0.021262f
C150 VTAIL.n108 B 0.009524f
C151 VTAIL.n109 B 0.01674f
C152 VTAIL.n110 B 0.008995f
C153 VTAIL.n111 B 0.021262f
C154 VTAIL.n112 B 0.009524f
C155 VTAIL.n113 B 0.644947f
C156 VTAIL.n114 B 0.008995f
C157 VTAIL.t0 B 0.035671f
C158 VTAIL.n115 B 0.103474f
C159 VTAIL.n116 B 0.01503f
C160 VTAIL.n117 B 0.015946f
C161 VTAIL.n118 B 0.021262f
C162 VTAIL.n119 B 0.009524f
C163 VTAIL.n120 B 0.008995f
C164 VTAIL.n121 B 0.01674f
C165 VTAIL.n122 B 0.01674f
C166 VTAIL.n123 B 0.008995f
C167 VTAIL.n124 B 0.009524f
C168 VTAIL.n125 B 0.021262f
C169 VTAIL.n126 B 0.021262f
C170 VTAIL.n127 B 0.009524f
C171 VTAIL.n128 B 0.008995f
C172 VTAIL.n129 B 0.01674f
C173 VTAIL.n130 B 0.01674f
C174 VTAIL.n131 B 0.008995f
C175 VTAIL.n132 B 0.008995f
C176 VTAIL.n133 B 0.009524f
C177 VTAIL.n134 B 0.021262f
C178 VTAIL.n135 B 0.021262f
C179 VTAIL.n136 B 0.021262f
C180 VTAIL.n137 B 0.00926f
C181 VTAIL.n138 B 0.008995f
C182 VTAIL.n139 B 0.01674f
C183 VTAIL.n140 B 0.01674f
C184 VTAIL.n141 B 0.008995f
C185 VTAIL.n142 B 0.009524f
C186 VTAIL.n143 B 0.021262f
C187 VTAIL.n144 B 0.04443f
C188 VTAIL.n145 B 0.009524f
C189 VTAIL.n146 B 0.008995f
C190 VTAIL.n147 B 0.040523f
C191 VTAIL.n148 B 0.024751f
C192 VTAIL.n149 B 0.879769f
C193 VTAIL.n150 B 0.022626f
C194 VTAIL.n151 B 0.01674f
C195 VTAIL.n152 B 0.008995f
C196 VTAIL.n153 B 0.021262f
C197 VTAIL.n154 B 0.00926f
C198 VTAIL.n155 B 0.01674f
C199 VTAIL.n156 B 0.00926f
C200 VTAIL.n157 B 0.008995f
C201 VTAIL.n158 B 0.021262f
C202 VTAIL.n159 B 0.021262f
C203 VTAIL.n160 B 0.009524f
C204 VTAIL.n161 B 0.01674f
C205 VTAIL.n162 B 0.008995f
C206 VTAIL.n163 B 0.021262f
C207 VTAIL.n164 B 0.009524f
C208 VTAIL.n165 B 0.644947f
C209 VTAIL.n166 B 0.008995f
C210 VTAIL.t7 B 0.035671f
C211 VTAIL.n167 B 0.103474f
C212 VTAIL.n168 B 0.01503f
C213 VTAIL.n169 B 0.015946f
C214 VTAIL.n170 B 0.021262f
C215 VTAIL.n171 B 0.009524f
C216 VTAIL.n172 B 0.008995f
C217 VTAIL.n173 B 0.01674f
C218 VTAIL.n174 B 0.01674f
C219 VTAIL.n175 B 0.008995f
C220 VTAIL.n176 B 0.009524f
C221 VTAIL.n177 B 0.021262f
C222 VTAIL.n178 B 0.021262f
C223 VTAIL.n179 B 0.009524f
C224 VTAIL.n180 B 0.008995f
C225 VTAIL.n181 B 0.01674f
C226 VTAIL.n182 B 0.01674f
C227 VTAIL.n183 B 0.008995f
C228 VTAIL.n184 B 0.009524f
C229 VTAIL.n185 B 0.021262f
C230 VTAIL.n186 B 0.021262f
C231 VTAIL.n187 B 0.009524f
C232 VTAIL.n188 B 0.008995f
C233 VTAIL.n189 B 0.01674f
C234 VTAIL.n190 B 0.01674f
C235 VTAIL.n191 B 0.008995f
C236 VTAIL.n192 B 0.009524f
C237 VTAIL.n193 B 0.021262f
C238 VTAIL.n194 B 0.04443f
C239 VTAIL.n195 B 0.009524f
C240 VTAIL.n196 B 0.008995f
C241 VTAIL.n197 B 0.040523f
C242 VTAIL.n198 B 0.024751f
C243 VTAIL.n199 B 0.879769f
C244 VTAIL.n200 B 0.022626f
C245 VTAIL.n201 B 0.01674f
C246 VTAIL.n202 B 0.008995f
C247 VTAIL.n203 B 0.021262f
C248 VTAIL.n204 B 0.00926f
C249 VTAIL.n205 B 0.01674f
C250 VTAIL.n206 B 0.00926f
C251 VTAIL.n207 B 0.008995f
C252 VTAIL.n208 B 0.021262f
C253 VTAIL.n209 B 0.021262f
C254 VTAIL.n210 B 0.009524f
C255 VTAIL.n211 B 0.01674f
C256 VTAIL.n212 B 0.008995f
C257 VTAIL.n213 B 0.021262f
C258 VTAIL.n214 B 0.009524f
C259 VTAIL.n215 B 0.644947f
C260 VTAIL.n216 B 0.008995f
C261 VTAIL.t4 B 0.035671f
C262 VTAIL.n217 B 0.103474f
C263 VTAIL.n218 B 0.01503f
C264 VTAIL.n219 B 0.015946f
C265 VTAIL.n220 B 0.021262f
C266 VTAIL.n221 B 0.009524f
C267 VTAIL.n222 B 0.008995f
C268 VTAIL.n223 B 0.01674f
C269 VTAIL.n224 B 0.01674f
C270 VTAIL.n225 B 0.008995f
C271 VTAIL.n226 B 0.009524f
C272 VTAIL.n227 B 0.021262f
C273 VTAIL.n228 B 0.021262f
C274 VTAIL.n229 B 0.009524f
C275 VTAIL.n230 B 0.008995f
C276 VTAIL.n231 B 0.01674f
C277 VTAIL.n232 B 0.01674f
C278 VTAIL.n233 B 0.008995f
C279 VTAIL.n234 B 0.009524f
C280 VTAIL.n235 B 0.021262f
C281 VTAIL.n236 B 0.021262f
C282 VTAIL.n237 B 0.009524f
C283 VTAIL.n238 B 0.008995f
C284 VTAIL.n239 B 0.01674f
C285 VTAIL.n240 B 0.01674f
C286 VTAIL.n241 B 0.008995f
C287 VTAIL.n242 B 0.009524f
C288 VTAIL.n243 B 0.021262f
C289 VTAIL.n244 B 0.04443f
C290 VTAIL.n245 B 0.009524f
C291 VTAIL.n246 B 0.008995f
C292 VTAIL.n247 B 0.040523f
C293 VTAIL.n248 B 0.024751f
C294 VTAIL.n249 B 0.142508f
C295 VTAIL.n250 B 0.022626f
C296 VTAIL.n251 B 0.01674f
C297 VTAIL.n252 B 0.008995f
C298 VTAIL.n253 B 0.021262f
C299 VTAIL.n254 B 0.00926f
C300 VTAIL.n255 B 0.01674f
C301 VTAIL.n256 B 0.00926f
C302 VTAIL.n257 B 0.008995f
C303 VTAIL.n258 B 0.021262f
C304 VTAIL.n259 B 0.021262f
C305 VTAIL.n260 B 0.009524f
C306 VTAIL.n261 B 0.01674f
C307 VTAIL.n262 B 0.008995f
C308 VTAIL.n263 B 0.021262f
C309 VTAIL.n264 B 0.009524f
C310 VTAIL.n265 B 0.644947f
C311 VTAIL.n266 B 0.008995f
C312 VTAIL.t3 B 0.035671f
C313 VTAIL.n267 B 0.103474f
C314 VTAIL.n268 B 0.01503f
C315 VTAIL.n269 B 0.015946f
C316 VTAIL.n270 B 0.021262f
C317 VTAIL.n271 B 0.009524f
C318 VTAIL.n272 B 0.008995f
C319 VTAIL.n273 B 0.01674f
C320 VTAIL.n274 B 0.01674f
C321 VTAIL.n275 B 0.008995f
C322 VTAIL.n276 B 0.009524f
C323 VTAIL.n277 B 0.021262f
C324 VTAIL.n278 B 0.021262f
C325 VTAIL.n279 B 0.009524f
C326 VTAIL.n280 B 0.008995f
C327 VTAIL.n281 B 0.01674f
C328 VTAIL.n282 B 0.01674f
C329 VTAIL.n283 B 0.008995f
C330 VTAIL.n284 B 0.009524f
C331 VTAIL.n285 B 0.021262f
C332 VTAIL.n286 B 0.021262f
C333 VTAIL.n287 B 0.009524f
C334 VTAIL.n288 B 0.008995f
C335 VTAIL.n289 B 0.01674f
C336 VTAIL.n290 B 0.01674f
C337 VTAIL.n291 B 0.008995f
C338 VTAIL.n292 B 0.009524f
C339 VTAIL.n293 B 0.021262f
C340 VTAIL.n294 B 0.04443f
C341 VTAIL.n295 B 0.009524f
C342 VTAIL.n296 B 0.008995f
C343 VTAIL.n297 B 0.040523f
C344 VTAIL.n298 B 0.024751f
C345 VTAIL.n299 B 0.142508f
C346 VTAIL.n300 B 0.022626f
C347 VTAIL.n301 B 0.01674f
C348 VTAIL.n302 B 0.008995f
C349 VTAIL.n303 B 0.021262f
C350 VTAIL.n304 B 0.00926f
C351 VTAIL.n305 B 0.01674f
C352 VTAIL.n306 B 0.00926f
C353 VTAIL.n307 B 0.008995f
C354 VTAIL.n308 B 0.021262f
C355 VTAIL.n309 B 0.021262f
C356 VTAIL.n310 B 0.009524f
C357 VTAIL.n311 B 0.01674f
C358 VTAIL.n312 B 0.008995f
C359 VTAIL.n313 B 0.021262f
C360 VTAIL.n314 B 0.009524f
C361 VTAIL.n315 B 0.644947f
C362 VTAIL.n316 B 0.008995f
C363 VTAIL.t1 B 0.035671f
C364 VTAIL.n317 B 0.103474f
C365 VTAIL.n318 B 0.01503f
C366 VTAIL.n319 B 0.015946f
C367 VTAIL.n320 B 0.021262f
C368 VTAIL.n321 B 0.009524f
C369 VTAIL.n322 B 0.008995f
C370 VTAIL.n323 B 0.01674f
C371 VTAIL.n324 B 0.01674f
C372 VTAIL.n325 B 0.008995f
C373 VTAIL.n326 B 0.009524f
C374 VTAIL.n327 B 0.021262f
C375 VTAIL.n328 B 0.021262f
C376 VTAIL.n329 B 0.009524f
C377 VTAIL.n330 B 0.008995f
C378 VTAIL.n331 B 0.01674f
C379 VTAIL.n332 B 0.01674f
C380 VTAIL.n333 B 0.008995f
C381 VTAIL.n334 B 0.009524f
C382 VTAIL.n335 B 0.021262f
C383 VTAIL.n336 B 0.021262f
C384 VTAIL.n337 B 0.009524f
C385 VTAIL.n338 B 0.008995f
C386 VTAIL.n339 B 0.01674f
C387 VTAIL.n340 B 0.01674f
C388 VTAIL.n341 B 0.008995f
C389 VTAIL.n342 B 0.009524f
C390 VTAIL.n343 B 0.021262f
C391 VTAIL.n344 B 0.04443f
C392 VTAIL.n345 B 0.009524f
C393 VTAIL.n346 B 0.008995f
C394 VTAIL.n347 B 0.040523f
C395 VTAIL.n348 B 0.024751f
C396 VTAIL.n349 B 0.879769f
C397 VTAIL.n350 B 0.022626f
C398 VTAIL.n351 B 0.01674f
C399 VTAIL.n352 B 0.008995f
C400 VTAIL.n353 B 0.021262f
C401 VTAIL.n354 B 0.00926f
C402 VTAIL.n355 B 0.01674f
C403 VTAIL.n356 B 0.009524f
C404 VTAIL.n357 B 0.021262f
C405 VTAIL.n358 B 0.009524f
C406 VTAIL.n359 B 0.01674f
C407 VTAIL.n360 B 0.008995f
C408 VTAIL.n361 B 0.021262f
C409 VTAIL.n362 B 0.009524f
C410 VTAIL.n363 B 0.644947f
C411 VTAIL.n364 B 0.008995f
C412 VTAIL.t5 B 0.035671f
C413 VTAIL.n365 B 0.103474f
C414 VTAIL.n366 B 0.01503f
C415 VTAIL.n367 B 0.015946f
C416 VTAIL.n368 B 0.021262f
C417 VTAIL.n369 B 0.009524f
C418 VTAIL.n370 B 0.008995f
C419 VTAIL.n371 B 0.01674f
C420 VTAIL.n372 B 0.01674f
C421 VTAIL.n373 B 0.008995f
C422 VTAIL.n374 B 0.009524f
C423 VTAIL.n375 B 0.021262f
C424 VTAIL.n376 B 0.021262f
C425 VTAIL.n377 B 0.009524f
C426 VTAIL.n378 B 0.008995f
C427 VTAIL.n379 B 0.01674f
C428 VTAIL.n380 B 0.01674f
C429 VTAIL.n381 B 0.008995f
C430 VTAIL.n382 B 0.008995f
C431 VTAIL.n383 B 0.009524f
C432 VTAIL.n384 B 0.021262f
C433 VTAIL.n385 B 0.021262f
C434 VTAIL.n386 B 0.021262f
C435 VTAIL.n387 B 0.00926f
C436 VTAIL.n388 B 0.008995f
C437 VTAIL.n389 B 0.01674f
C438 VTAIL.n390 B 0.01674f
C439 VTAIL.n391 B 0.008995f
C440 VTAIL.n392 B 0.009524f
C441 VTAIL.n393 B 0.021262f
C442 VTAIL.n394 B 0.04443f
C443 VTAIL.n395 B 0.009524f
C444 VTAIL.n396 B 0.008995f
C445 VTAIL.n397 B 0.040523f
C446 VTAIL.n398 B 0.024751f
C447 VTAIL.n399 B 0.825713f
C448 VDD2.t0 B 0.197002f
C449 VDD2.t2 B 0.197002f
C450 VDD2.n0 B 2.25458f
C451 VDD2.t3 B 0.197002f
C452 VDD2.t1 B 0.197002f
C453 VDD2.n1 B 1.72709f
C454 VDD2.n2 B 3.26184f
C455 VN.t1 B 1.6655f
C456 VN.t2 B 1.66356f
C457 VN.n0 B 1.15025f
C458 VN.t3 B 1.6655f
C459 VN.t0 B 1.66356f
C460 VN.n1 B 2.42967f
.ends

