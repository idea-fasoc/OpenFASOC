* NGSPICE file created from diff_pair_sample_0855.ext - technology: sky130A

.subckt diff_pair_sample_0855 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t5 VN.t0 VTAIL.t6 w_n2938_n1294# sky130_fd_pr__pfet_01v8 ad=0.26895 pd=1.96 as=0.6357 ps=4.04 w=1.63 l=2.13
X1 VTAIL.t3 VP.t0 VDD1.t5 w_n2938_n1294# sky130_fd_pr__pfet_01v8 ad=0.26895 pd=1.96 as=0.26895 ps=1.96 w=1.63 l=2.13
X2 B.t11 B.t9 B.t10 w_n2938_n1294# sky130_fd_pr__pfet_01v8 ad=0.6357 pd=4.04 as=0 ps=0 w=1.63 l=2.13
X3 VTAIL.t9 VN.t1 VDD2.t4 w_n2938_n1294# sky130_fd_pr__pfet_01v8 ad=0.26895 pd=1.96 as=0.26895 ps=1.96 w=1.63 l=2.13
X4 B.t8 B.t6 B.t7 w_n2938_n1294# sky130_fd_pr__pfet_01v8 ad=0.6357 pd=4.04 as=0 ps=0 w=1.63 l=2.13
X5 B.t5 B.t3 B.t4 w_n2938_n1294# sky130_fd_pr__pfet_01v8 ad=0.6357 pd=4.04 as=0 ps=0 w=1.63 l=2.13
X6 VDD2.t3 VN.t2 VTAIL.t8 w_n2938_n1294# sky130_fd_pr__pfet_01v8 ad=0.26895 pd=1.96 as=0.6357 ps=4.04 w=1.63 l=2.13
X7 VDD1.t4 VP.t1 VTAIL.t4 w_n2938_n1294# sky130_fd_pr__pfet_01v8 ad=0.26895 pd=1.96 as=0.6357 ps=4.04 w=1.63 l=2.13
X8 VTAIL.t7 VN.t3 VDD2.t2 w_n2938_n1294# sky130_fd_pr__pfet_01v8 ad=0.26895 pd=1.96 as=0.26895 ps=1.96 w=1.63 l=2.13
X9 VDD2.t1 VN.t4 VTAIL.t10 w_n2938_n1294# sky130_fd_pr__pfet_01v8 ad=0.6357 pd=4.04 as=0.26895 ps=1.96 w=1.63 l=2.13
X10 VDD1.t3 VP.t2 VTAIL.t2 w_n2938_n1294# sky130_fd_pr__pfet_01v8 ad=0.6357 pd=4.04 as=0.26895 ps=1.96 w=1.63 l=2.13
X11 B.t2 B.t0 B.t1 w_n2938_n1294# sky130_fd_pr__pfet_01v8 ad=0.6357 pd=4.04 as=0 ps=0 w=1.63 l=2.13
X12 VDD1.t2 VP.t3 VTAIL.t5 w_n2938_n1294# sky130_fd_pr__pfet_01v8 ad=0.6357 pd=4.04 as=0.26895 ps=1.96 w=1.63 l=2.13
X13 VTAIL.t1 VP.t4 VDD1.t1 w_n2938_n1294# sky130_fd_pr__pfet_01v8 ad=0.26895 pd=1.96 as=0.26895 ps=1.96 w=1.63 l=2.13
X14 VDD2.t0 VN.t5 VTAIL.t11 w_n2938_n1294# sky130_fd_pr__pfet_01v8 ad=0.6357 pd=4.04 as=0.26895 ps=1.96 w=1.63 l=2.13
X15 VDD1.t0 VP.t5 VTAIL.t0 w_n2938_n1294# sky130_fd_pr__pfet_01v8 ad=0.26895 pd=1.96 as=0.6357 ps=4.04 w=1.63 l=2.13
R0 VN.n21 VN.n12 161.3
R1 VN.n20 VN.n19 161.3
R2 VN.n18 VN.n13 161.3
R3 VN.n17 VN.n16 161.3
R4 VN.n9 VN.n0 161.3
R5 VN.n8 VN.n7 161.3
R6 VN.n6 VN.n1 161.3
R7 VN.n5 VN.n4 161.3
R8 VN.n11 VN.n10 88.2468
R9 VN.n23 VN.n22 88.2468
R10 VN.n8 VN.n1 56.5193
R11 VN.n20 VN.n13 56.5193
R12 VN.n2 VN.t4 52.972
R13 VN.n14 VN.t2 52.972
R14 VN.n15 VN.n14 46.3041
R15 VN.n3 VN.n2 46.3041
R16 VN VN.n23 39.3542
R17 VN.n4 VN.n3 24.4675
R18 VN.n4 VN.n1 24.4675
R19 VN.n9 VN.n8 24.4675
R20 VN.n16 VN.n13 24.4675
R21 VN.n16 VN.n15 24.4675
R22 VN.n21 VN.n20 24.4675
R23 VN.n10 VN.n9 22.5101
R24 VN.n22 VN.n21 22.5101
R25 VN.n3 VN.t1 18.4432
R26 VN.n10 VN.t0 18.4432
R27 VN.n15 VN.t3 18.4432
R28 VN.n22 VN.t5 18.4432
R29 VN.n17 VN.n14 8.73622
R30 VN.n5 VN.n2 8.73622
R31 VN.n23 VN.n12 0.278367
R32 VN.n11 VN.n0 0.278367
R33 VN.n19 VN.n12 0.189894
R34 VN.n19 VN.n18 0.189894
R35 VN.n18 VN.n17 0.189894
R36 VN.n6 VN.n5 0.189894
R37 VN.n7 VN.n6 0.189894
R38 VN.n7 VN.n0 0.189894
R39 VN VN.n11 0.153454
R40 VTAIL.n11 VTAIL.t6 252.405
R41 VTAIL.n2 VTAIL.t4 252.405
R42 VTAIL.n10 VTAIL.t0 252.405
R43 VTAIL.n7 VTAIL.t8 252.405
R44 VTAIL.n1 VTAIL.n0 232.464
R45 VTAIL.n4 VTAIL.n3 232.464
R46 VTAIL.n9 VTAIL.n8 232.464
R47 VTAIL.n6 VTAIL.n5 232.464
R48 VTAIL.n0 VTAIL.t10 19.9422
R49 VTAIL.n0 VTAIL.t9 19.9422
R50 VTAIL.n3 VTAIL.t2 19.9422
R51 VTAIL.n3 VTAIL.t3 19.9422
R52 VTAIL.n8 VTAIL.t5 19.9422
R53 VTAIL.n8 VTAIL.t1 19.9422
R54 VTAIL.n5 VTAIL.t11 19.9422
R55 VTAIL.n5 VTAIL.t7 19.9422
R56 VTAIL.n6 VTAIL.n4 18.0134
R57 VTAIL.n11 VTAIL.n10 15.8927
R58 VTAIL.n7 VTAIL.n6 2.12119
R59 VTAIL.n10 VTAIL.n9 2.12119
R60 VTAIL.n4 VTAIL.n2 2.12119
R61 VTAIL VTAIL.n11 1.53283
R62 VTAIL.n9 VTAIL.n7 1.53067
R63 VTAIL.n2 VTAIL.n1 1.53067
R64 VTAIL VTAIL.n1 0.588862
R65 VDD2.n1 VDD2.t1 270.618
R66 VDD2.n2 VDD2.t0 269.084
R67 VDD2.n1 VDD2.n0 249.617
R68 VDD2 VDD2.n3 249.613
R69 VDD2.n2 VDD2.n1 32.0127
R70 VDD2.n3 VDD2.t2 19.9422
R71 VDD2.n3 VDD2.t3 19.9422
R72 VDD2.n0 VDD2.t4 19.9422
R73 VDD2.n0 VDD2.t5 19.9422
R74 VDD2 VDD2.n2 1.64921
R75 VP.n10 VP.n9 161.3
R76 VP.n11 VP.n6 161.3
R77 VP.n13 VP.n12 161.3
R78 VP.n14 VP.n5 161.3
R79 VP.n31 VP.n0 161.3
R80 VP.n30 VP.n29 161.3
R81 VP.n28 VP.n1 161.3
R82 VP.n27 VP.n26 161.3
R83 VP.n25 VP.n2 161.3
R84 VP.n24 VP.n23 161.3
R85 VP.n22 VP.n3 161.3
R86 VP.n21 VP.n20 161.3
R87 VP.n19 VP.n4 161.3
R88 VP.n18 VP.n17 88.2468
R89 VP.n33 VP.n32 88.2468
R90 VP.n16 VP.n15 88.2468
R91 VP.n20 VP.n3 56.5193
R92 VP.n30 VP.n1 56.5193
R93 VP.n13 VP.n6 56.5193
R94 VP.n7 VP.t3 52.972
R95 VP.n8 VP.n7 46.3041
R96 VP.n17 VP.n16 39.0753
R97 VP.n20 VP.n19 24.4675
R98 VP.n24 VP.n3 24.4675
R99 VP.n25 VP.n24 24.4675
R100 VP.n26 VP.n25 24.4675
R101 VP.n26 VP.n1 24.4675
R102 VP.n31 VP.n30 24.4675
R103 VP.n14 VP.n13 24.4675
R104 VP.n9 VP.n8 24.4675
R105 VP.n9 VP.n6 24.4675
R106 VP.n19 VP.n18 22.5101
R107 VP.n32 VP.n31 22.5101
R108 VP.n15 VP.n14 22.5101
R109 VP.n25 VP.t0 18.4432
R110 VP.n18 VP.t2 18.4432
R111 VP.n32 VP.t1 18.4432
R112 VP.n8 VP.t4 18.4432
R113 VP.n15 VP.t5 18.4432
R114 VP.n10 VP.n7 8.73622
R115 VP.n16 VP.n5 0.278367
R116 VP.n17 VP.n4 0.278367
R117 VP.n33 VP.n0 0.278367
R118 VP.n11 VP.n10 0.189894
R119 VP.n12 VP.n11 0.189894
R120 VP.n12 VP.n5 0.189894
R121 VP.n21 VP.n4 0.189894
R122 VP.n22 VP.n21 0.189894
R123 VP.n23 VP.n22 0.189894
R124 VP.n23 VP.n2 0.189894
R125 VP.n27 VP.n2 0.189894
R126 VP.n28 VP.n27 0.189894
R127 VP.n29 VP.n28 0.189894
R128 VP.n29 VP.n0 0.189894
R129 VP VP.n33 0.153454
R130 VDD1 VDD1.t2 270.733
R131 VDD1.n1 VDD1.t3 270.618
R132 VDD1.n1 VDD1.n0 249.617
R133 VDD1.n3 VDD1.n2 249.142
R134 VDD1.n3 VDD1.n1 33.6561
R135 VDD1.n2 VDD1.t1 19.9422
R136 VDD1.n2 VDD1.t0 19.9422
R137 VDD1.n0 VDD1.t5 19.9422
R138 VDD1.n0 VDD1.t4 19.9422
R139 VDD1 VDD1.n3 0.472483
R140 B.n334 B.n333 585
R141 B.n335 B.n40 585
R142 B.n337 B.n336 585
R143 B.n338 B.n39 585
R144 B.n340 B.n339 585
R145 B.n341 B.n38 585
R146 B.n343 B.n342 585
R147 B.n344 B.n37 585
R148 B.n346 B.n345 585
R149 B.n347 B.n36 585
R150 B.n349 B.n348 585
R151 B.n351 B.n33 585
R152 B.n353 B.n352 585
R153 B.n354 B.n32 585
R154 B.n356 B.n355 585
R155 B.n357 B.n31 585
R156 B.n359 B.n358 585
R157 B.n360 B.n30 585
R158 B.n362 B.n361 585
R159 B.n363 B.n29 585
R160 B.n365 B.n364 585
R161 B.n367 B.n366 585
R162 B.n368 B.n25 585
R163 B.n370 B.n369 585
R164 B.n371 B.n24 585
R165 B.n373 B.n372 585
R166 B.n374 B.n23 585
R167 B.n376 B.n375 585
R168 B.n377 B.n22 585
R169 B.n379 B.n378 585
R170 B.n380 B.n21 585
R171 B.n382 B.n381 585
R172 B.n332 B.n41 585
R173 B.n331 B.n330 585
R174 B.n329 B.n42 585
R175 B.n328 B.n327 585
R176 B.n326 B.n43 585
R177 B.n325 B.n324 585
R178 B.n323 B.n44 585
R179 B.n322 B.n321 585
R180 B.n320 B.n45 585
R181 B.n319 B.n318 585
R182 B.n317 B.n46 585
R183 B.n316 B.n315 585
R184 B.n314 B.n47 585
R185 B.n313 B.n312 585
R186 B.n311 B.n48 585
R187 B.n310 B.n309 585
R188 B.n308 B.n49 585
R189 B.n307 B.n306 585
R190 B.n305 B.n50 585
R191 B.n304 B.n303 585
R192 B.n302 B.n51 585
R193 B.n301 B.n300 585
R194 B.n299 B.n52 585
R195 B.n298 B.n297 585
R196 B.n296 B.n53 585
R197 B.n295 B.n294 585
R198 B.n293 B.n54 585
R199 B.n292 B.n291 585
R200 B.n290 B.n55 585
R201 B.n289 B.n288 585
R202 B.n287 B.n56 585
R203 B.n286 B.n285 585
R204 B.n284 B.n57 585
R205 B.n283 B.n282 585
R206 B.n281 B.n58 585
R207 B.n280 B.n279 585
R208 B.n278 B.n59 585
R209 B.n277 B.n276 585
R210 B.n275 B.n60 585
R211 B.n274 B.n273 585
R212 B.n272 B.n61 585
R213 B.n271 B.n270 585
R214 B.n269 B.n62 585
R215 B.n268 B.n267 585
R216 B.n266 B.n63 585
R217 B.n265 B.n264 585
R218 B.n263 B.n64 585
R219 B.n262 B.n261 585
R220 B.n260 B.n65 585
R221 B.n259 B.n258 585
R222 B.n257 B.n66 585
R223 B.n256 B.n255 585
R224 B.n254 B.n67 585
R225 B.n253 B.n252 585
R226 B.n251 B.n68 585
R227 B.n250 B.n249 585
R228 B.n248 B.n69 585
R229 B.n247 B.n246 585
R230 B.n245 B.n70 585
R231 B.n244 B.n243 585
R232 B.n242 B.n71 585
R233 B.n241 B.n240 585
R234 B.n239 B.n72 585
R235 B.n238 B.n237 585
R236 B.n236 B.n73 585
R237 B.n235 B.n234 585
R238 B.n233 B.n74 585
R239 B.n232 B.n231 585
R240 B.n230 B.n75 585
R241 B.n229 B.n228 585
R242 B.n227 B.n76 585
R243 B.n226 B.n225 585
R244 B.n224 B.n77 585
R245 B.n223 B.n222 585
R246 B.n221 B.n78 585
R247 B.n172 B.n171 585
R248 B.n173 B.n98 585
R249 B.n175 B.n174 585
R250 B.n176 B.n97 585
R251 B.n178 B.n177 585
R252 B.n179 B.n96 585
R253 B.n181 B.n180 585
R254 B.n182 B.n95 585
R255 B.n184 B.n183 585
R256 B.n185 B.n94 585
R257 B.n187 B.n186 585
R258 B.n189 B.n91 585
R259 B.n191 B.n190 585
R260 B.n192 B.n90 585
R261 B.n194 B.n193 585
R262 B.n195 B.n89 585
R263 B.n197 B.n196 585
R264 B.n198 B.n88 585
R265 B.n200 B.n199 585
R266 B.n201 B.n87 585
R267 B.n203 B.n202 585
R268 B.n205 B.n204 585
R269 B.n206 B.n83 585
R270 B.n208 B.n207 585
R271 B.n209 B.n82 585
R272 B.n211 B.n210 585
R273 B.n212 B.n81 585
R274 B.n214 B.n213 585
R275 B.n215 B.n80 585
R276 B.n217 B.n216 585
R277 B.n218 B.n79 585
R278 B.n220 B.n219 585
R279 B.n170 B.n99 585
R280 B.n169 B.n168 585
R281 B.n167 B.n100 585
R282 B.n166 B.n165 585
R283 B.n164 B.n101 585
R284 B.n163 B.n162 585
R285 B.n161 B.n102 585
R286 B.n160 B.n159 585
R287 B.n158 B.n103 585
R288 B.n157 B.n156 585
R289 B.n155 B.n104 585
R290 B.n154 B.n153 585
R291 B.n152 B.n105 585
R292 B.n151 B.n150 585
R293 B.n149 B.n106 585
R294 B.n148 B.n147 585
R295 B.n146 B.n107 585
R296 B.n145 B.n144 585
R297 B.n143 B.n108 585
R298 B.n142 B.n141 585
R299 B.n140 B.n109 585
R300 B.n139 B.n138 585
R301 B.n137 B.n110 585
R302 B.n136 B.n135 585
R303 B.n134 B.n111 585
R304 B.n133 B.n132 585
R305 B.n131 B.n112 585
R306 B.n130 B.n129 585
R307 B.n128 B.n113 585
R308 B.n127 B.n126 585
R309 B.n125 B.n114 585
R310 B.n124 B.n123 585
R311 B.n122 B.n115 585
R312 B.n121 B.n120 585
R313 B.n119 B.n116 585
R314 B.n118 B.n117 585
R315 B.n2 B.n0 585
R316 B.n437 B.n1 585
R317 B.n436 B.n435 585
R318 B.n434 B.n3 585
R319 B.n433 B.n432 585
R320 B.n431 B.n4 585
R321 B.n430 B.n429 585
R322 B.n428 B.n5 585
R323 B.n427 B.n426 585
R324 B.n425 B.n6 585
R325 B.n424 B.n423 585
R326 B.n422 B.n7 585
R327 B.n421 B.n420 585
R328 B.n419 B.n8 585
R329 B.n418 B.n417 585
R330 B.n416 B.n9 585
R331 B.n415 B.n414 585
R332 B.n413 B.n10 585
R333 B.n412 B.n411 585
R334 B.n410 B.n11 585
R335 B.n409 B.n408 585
R336 B.n407 B.n12 585
R337 B.n406 B.n405 585
R338 B.n404 B.n13 585
R339 B.n403 B.n402 585
R340 B.n401 B.n14 585
R341 B.n400 B.n399 585
R342 B.n398 B.n15 585
R343 B.n397 B.n396 585
R344 B.n395 B.n16 585
R345 B.n394 B.n393 585
R346 B.n392 B.n17 585
R347 B.n391 B.n390 585
R348 B.n389 B.n18 585
R349 B.n388 B.n387 585
R350 B.n386 B.n19 585
R351 B.n385 B.n384 585
R352 B.n383 B.n20 585
R353 B.n439 B.n438 585
R354 B.n172 B.n99 492.5
R355 B.n383 B.n382 492.5
R356 B.n221 B.n220 492.5
R357 B.n334 B.n41 492.5
R358 B.n84 B.t2 297.95
R359 B.n34 B.t7 297.95
R360 B.n92 B.t5 297.95
R361 B.n26 B.t10 297.95
R362 B.n85 B.t1 250.24
R363 B.n35 B.t8 250.24
R364 B.n93 B.t4 250.24
R365 B.n27 B.t11 250.24
R366 B.n84 B.t0 225.65
R367 B.n92 B.t3 225.65
R368 B.n26 B.t9 225.65
R369 B.n34 B.t6 225.65
R370 B.n168 B.n99 163.367
R371 B.n168 B.n167 163.367
R372 B.n167 B.n166 163.367
R373 B.n166 B.n101 163.367
R374 B.n162 B.n101 163.367
R375 B.n162 B.n161 163.367
R376 B.n161 B.n160 163.367
R377 B.n160 B.n103 163.367
R378 B.n156 B.n103 163.367
R379 B.n156 B.n155 163.367
R380 B.n155 B.n154 163.367
R381 B.n154 B.n105 163.367
R382 B.n150 B.n105 163.367
R383 B.n150 B.n149 163.367
R384 B.n149 B.n148 163.367
R385 B.n148 B.n107 163.367
R386 B.n144 B.n107 163.367
R387 B.n144 B.n143 163.367
R388 B.n143 B.n142 163.367
R389 B.n142 B.n109 163.367
R390 B.n138 B.n109 163.367
R391 B.n138 B.n137 163.367
R392 B.n137 B.n136 163.367
R393 B.n136 B.n111 163.367
R394 B.n132 B.n111 163.367
R395 B.n132 B.n131 163.367
R396 B.n131 B.n130 163.367
R397 B.n130 B.n113 163.367
R398 B.n126 B.n113 163.367
R399 B.n126 B.n125 163.367
R400 B.n125 B.n124 163.367
R401 B.n124 B.n115 163.367
R402 B.n120 B.n115 163.367
R403 B.n120 B.n119 163.367
R404 B.n119 B.n118 163.367
R405 B.n118 B.n2 163.367
R406 B.n438 B.n2 163.367
R407 B.n438 B.n437 163.367
R408 B.n437 B.n436 163.367
R409 B.n436 B.n3 163.367
R410 B.n432 B.n3 163.367
R411 B.n432 B.n431 163.367
R412 B.n431 B.n430 163.367
R413 B.n430 B.n5 163.367
R414 B.n426 B.n5 163.367
R415 B.n426 B.n425 163.367
R416 B.n425 B.n424 163.367
R417 B.n424 B.n7 163.367
R418 B.n420 B.n7 163.367
R419 B.n420 B.n419 163.367
R420 B.n419 B.n418 163.367
R421 B.n418 B.n9 163.367
R422 B.n414 B.n9 163.367
R423 B.n414 B.n413 163.367
R424 B.n413 B.n412 163.367
R425 B.n412 B.n11 163.367
R426 B.n408 B.n11 163.367
R427 B.n408 B.n407 163.367
R428 B.n407 B.n406 163.367
R429 B.n406 B.n13 163.367
R430 B.n402 B.n13 163.367
R431 B.n402 B.n401 163.367
R432 B.n401 B.n400 163.367
R433 B.n400 B.n15 163.367
R434 B.n396 B.n15 163.367
R435 B.n396 B.n395 163.367
R436 B.n395 B.n394 163.367
R437 B.n394 B.n17 163.367
R438 B.n390 B.n17 163.367
R439 B.n390 B.n389 163.367
R440 B.n389 B.n388 163.367
R441 B.n388 B.n19 163.367
R442 B.n384 B.n19 163.367
R443 B.n384 B.n383 163.367
R444 B.n173 B.n172 163.367
R445 B.n174 B.n173 163.367
R446 B.n174 B.n97 163.367
R447 B.n178 B.n97 163.367
R448 B.n179 B.n178 163.367
R449 B.n180 B.n179 163.367
R450 B.n180 B.n95 163.367
R451 B.n184 B.n95 163.367
R452 B.n185 B.n184 163.367
R453 B.n186 B.n185 163.367
R454 B.n186 B.n91 163.367
R455 B.n191 B.n91 163.367
R456 B.n192 B.n191 163.367
R457 B.n193 B.n192 163.367
R458 B.n193 B.n89 163.367
R459 B.n197 B.n89 163.367
R460 B.n198 B.n197 163.367
R461 B.n199 B.n198 163.367
R462 B.n199 B.n87 163.367
R463 B.n203 B.n87 163.367
R464 B.n204 B.n203 163.367
R465 B.n204 B.n83 163.367
R466 B.n208 B.n83 163.367
R467 B.n209 B.n208 163.367
R468 B.n210 B.n209 163.367
R469 B.n210 B.n81 163.367
R470 B.n214 B.n81 163.367
R471 B.n215 B.n214 163.367
R472 B.n216 B.n215 163.367
R473 B.n216 B.n79 163.367
R474 B.n220 B.n79 163.367
R475 B.n222 B.n221 163.367
R476 B.n222 B.n77 163.367
R477 B.n226 B.n77 163.367
R478 B.n227 B.n226 163.367
R479 B.n228 B.n227 163.367
R480 B.n228 B.n75 163.367
R481 B.n232 B.n75 163.367
R482 B.n233 B.n232 163.367
R483 B.n234 B.n233 163.367
R484 B.n234 B.n73 163.367
R485 B.n238 B.n73 163.367
R486 B.n239 B.n238 163.367
R487 B.n240 B.n239 163.367
R488 B.n240 B.n71 163.367
R489 B.n244 B.n71 163.367
R490 B.n245 B.n244 163.367
R491 B.n246 B.n245 163.367
R492 B.n246 B.n69 163.367
R493 B.n250 B.n69 163.367
R494 B.n251 B.n250 163.367
R495 B.n252 B.n251 163.367
R496 B.n252 B.n67 163.367
R497 B.n256 B.n67 163.367
R498 B.n257 B.n256 163.367
R499 B.n258 B.n257 163.367
R500 B.n258 B.n65 163.367
R501 B.n262 B.n65 163.367
R502 B.n263 B.n262 163.367
R503 B.n264 B.n263 163.367
R504 B.n264 B.n63 163.367
R505 B.n268 B.n63 163.367
R506 B.n269 B.n268 163.367
R507 B.n270 B.n269 163.367
R508 B.n270 B.n61 163.367
R509 B.n274 B.n61 163.367
R510 B.n275 B.n274 163.367
R511 B.n276 B.n275 163.367
R512 B.n276 B.n59 163.367
R513 B.n280 B.n59 163.367
R514 B.n281 B.n280 163.367
R515 B.n282 B.n281 163.367
R516 B.n282 B.n57 163.367
R517 B.n286 B.n57 163.367
R518 B.n287 B.n286 163.367
R519 B.n288 B.n287 163.367
R520 B.n288 B.n55 163.367
R521 B.n292 B.n55 163.367
R522 B.n293 B.n292 163.367
R523 B.n294 B.n293 163.367
R524 B.n294 B.n53 163.367
R525 B.n298 B.n53 163.367
R526 B.n299 B.n298 163.367
R527 B.n300 B.n299 163.367
R528 B.n300 B.n51 163.367
R529 B.n304 B.n51 163.367
R530 B.n305 B.n304 163.367
R531 B.n306 B.n305 163.367
R532 B.n306 B.n49 163.367
R533 B.n310 B.n49 163.367
R534 B.n311 B.n310 163.367
R535 B.n312 B.n311 163.367
R536 B.n312 B.n47 163.367
R537 B.n316 B.n47 163.367
R538 B.n317 B.n316 163.367
R539 B.n318 B.n317 163.367
R540 B.n318 B.n45 163.367
R541 B.n322 B.n45 163.367
R542 B.n323 B.n322 163.367
R543 B.n324 B.n323 163.367
R544 B.n324 B.n43 163.367
R545 B.n328 B.n43 163.367
R546 B.n329 B.n328 163.367
R547 B.n330 B.n329 163.367
R548 B.n330 B.n41 163.367
R549 B.n382 B.n21 163.367
R550 B.n378 B.n21 163.367
R551 B.n378 B.n377 163.367
R552 B.n377 B.n376 163.367
R553 B.n376 B.n23 163.367
R554 B.n372 B.n23 163.367
R555 B.n372 B.n371 163.367
R556 B.n371 B.n370 163.367
R557 B.n370 B.n25 163.367
R558 B.n366 B.n25 163.367
R559 B.n366 B.n365 163.367
R560 B.n365 B.n29 163.367
R561 B.n361 B.n29 163.367
R562 B.n361 B.n360 163.367
R563 B.n360 B.n359 163.367
R564 B.n359 B.n31 163.367
R565 B.n355 B.n31 163.367
R566 B.n355 B.n354 163.367
R567 B.n354 B.n353 163.367
R568 B.n353 B.n33 163.367
R569 B.n348 B.n33 163.367
R570 B.n348 B.n347 163.367
R571 B.n347 B.n346 163.367
R572 B.n346 B.n37 163.367
R573 B.n342 B.n37 163.367
R574 B.n342 B.n341 163.367
R575 B.n341 B.n340 163.367
R576 B.n340 B.n39 163.367
R577 B.n336 B.n39 163.367
R578 B.n336 B.n335 163.367
R579 B.n335 B.n334 163.367
R580 B.n86 B.n85 59.5399
R581 B.n188 B.n93 59.5399
R582 B.n28 B.n27 59.5399
R583 B.n350 B.n35 59.5399
R584 B.n85 B.n84 47.7096
R585 B.n93 B.n92 47.7096
R586 B.n27 B.n26 47.7096
R587 B.n35 B.n34 47.7096
R588 B.n381 B.n20 32.0005
R589 B.n333 B.n332 32.0005
R590 B.n219 B.n78 32.0005
R591 B.n171 B.n170 32.0005
R592 B B.n439 18.0485
R593 B.n381 B.n380 10.6151
R594 B.n380 B.n379 10.6151
R595 B.n379 B.n22 10.6151
R596 B.n375 B.n22 10.6151
R597 B.n375 B.n374 10.6151
R598 B.n374 B.n373 10.6151
R599 B.n373 B.n24 10.6151
R600 B.n369 B.n24 10.6151
R601 B.n369 B.n368 10.6151
R602 B.n368 B.n367 10.6151
R603 B.n364 B.n363 10.6151
R604 B.n363 B.n362 10.6151
R605 B.n362 B.n30 10.6151
R606 B.n358 B.n30 10.6151
R607 B.n358 B.n357 10.6151
R608 B.n357 B.n356 10.6151
R609 B.n356 B.n32 10.6151
R610 B.n352 B.n32 10.6151
R611 B.n352 B.n351 10.6151
R612 B.n349 B.n36 10.6151
R613 B.n345 B.n36 10.6151
R614 B.n345 B.n344 10.6151
R615 B.n344 B.n343 10.6151
R616 B.n343 B.n38 10.6151
R617 B.n339 B.n38 10.6151
R618 B.n339 B.n338 10.6151
R619 B.n338 B.n337 10.6151
R620 B.n337 B.n40 10.6151
R621 B.n333 B.n40 10.6151
R622 B.n223 B.n78 10.6151
R623 B.n224 B.n223 10.6151
R624 B.n225 B.n224 10.6151
R625 B.n225 B.n76 10.6151
R626 B.n229 B.n76 10.6151
R627 B.n230 B.n229 10.6151
R628 B.n231 B.n230 10.6151
R629 B.n231 B.n74 10.6151
R630 B.n235 B.n74 10.6151
R631 B.n236 B.n235 10.6151
R632 B.n237 B.n236 10.6151
R633 B.n237 B.n72 10.6151
R634 B.n241 B.n72 10.6151
R635 B.n242 B.n241 10.6151
R636 B.n243 B.n242 10.6151
R637 B.n243 B.n70 10.6151
R638 B.n247 B.n70 10.6151
R639 B.n248 B.n247 10.6151
R640 B.n249 B.n248 10.6151
R641 B.n249 B.n68 10.6151
R642 B.n253 B.n68 10.6151
R643 B.n254 B.n253 10.6151
R644 B.n255 B.n254 10.6151
R645 B.n255 B.n66 10.6151
R646 B.n259 B.n66 10.6151
R647 B.n260 B.n259 10.6151
R648 B.n261 B.n260 10.6151
R649 B.n261 B.n64 10.6151
R650 B.n265 B.n64 10.6151
R651 B.n266 B.n265 10.6151
R652 B.n267 B.n266 10.6151
R653 B.n267 B.n62 10.6151
R654 B.n271 B.n62 10.6151
R655 B.n272 B.n271 10.6151
R656 B.n273 B.n272 10.6151
R657 B.n273 B.n60 10.6151
R658 B.n277 B.n60 10.6151
R659 B.n278 B.n277 10.6151
R660 B.n279 B.n278 10.6151
R661 B.n279 B.n58 10.6151
R662 B.n283 B.n58 10.6151
R663 B.n284 B.n283 10.6151
R664 B.n285 B.n284 10.6151
R665 B.n285 B.n56 10.6151
R666 B.n289 B.n56 10.6151
R667 B.n290 B.n289 10.6151
R668 B.n291 B.n290 10.6151
R669 B.n291 B.n54 10.6151
R670 B.n295 B.n54 10.6151
R671 B.n296 B.n295 10.6151
R672 B.n297 B.n296 10.6151
R673 B.n297 B.n52 10.6151
R674 B.n301 B.n52 10.6151
R675 B.n302 B.n301 10.6151
R676 B.n303 B.n302 10.6151
R677 B.n303 B.n50 10.6151
R678 B.n307 B.n50 10.6151
R679 B.n308 B.n307 10.6151
R680 B.n309 B.n308 10.6151
R681 B.n309 B.n48 10.6151
R682 B.n313 B.n48 10.6151
R683 B.n314 B.n313 10.6151
R684 B.n315 B.n314 10.6151
R685 B.n315 B.n46 10.6151
R686 B.n319 B.n46 10.6151
R687 B.n320 B.n319 10.6151
R688 B.n321 B.n320 10.6151
R689 B.n321 B.n44 10.6151
R690 B.n325 B.n44 10.6151
R691 B.n326 B.n325 10.6151
R692 B.n327 B.n326 10.6151
R693 B.n327 B.n42 10.6151
R694 B.n331 B.n42 10.6151
R695 B.n332 B.n331 10.6151
R696 B.n171 B.n98 10.6151
R697 B.n175 B.n98 10.6151
R698 B.n176 B.n175 10.6151
R699 B.n177 B.n176 10.6151
R700 B.n177 B.n96 10.6151
R701 B.n181 B.n96 10.6151
R702 B.n182 B.n181 10.6151
R703 B.n183 B.n182 10.6151
R704 B.n183 B.n94 10.6151
R705 B.n187 B.n94 10.6151
R706 B.n190 B.n189 10.6151
R707 B.n190 B.n90 10.6151
R708 B.n194 B.n90 10.6151
R709 B.n195 B.n194 10.6151
R710 B.n196 B.n195 10.6151
R711 B.n196 B.n88 10.6151
R712 B.n200 B.n88 10.6151
R713 B.n201 B.n200 10.6151
R714 B.n202 B.n201 10.6151
R715 B.n206 B.n205 10.6151
R716 B.n207 B.n206 10.6151
R717 B.n207 B.n82 10.6151
R718 B.n211 B.n82 10.6151
R719 B.n212 B.n211 10.6151
R720 B.n213 B.n212 10.6151
R721 B.n213 B.n80 10.6151
R722 B.n217 B.n80 10.6151
R723 B.n218 B.n217 10.6151
R724 B.n219 B.n218 10.6151
R725 B.n170 B.n169 10.6151
R726 B.n169 B.n100 10.6151
R727 B.n165 B.n100 10.6151
R728 B.n165 B.n164 10.6151
R729 B.n164 B.n163 10.6151
R730 B.n163 B.n102 10.6151
R731 B.n159 B.n102 10.6151
R732 B.n159 B.n158 10.6151
R733 B.n158 B.n157 10.6151
R734 B.n157 B.n104 10.6151
R735 B.n153 B.n104 10.6151
R736 B.n153 B.n152 10.6151
R737 B.n152 B.n151 10.6151
R738 B.n151 B.n106 10.6151
R739 B.n147 B.n106 10.6151
R740 B.n147 B.n146 10.6151
R741 B.n146 B.n145 10.6151
R742 B.n145 B.n108 10.6151
R743 B.n141 B.n108 10.6151
R744 B.n141 B.n140 10.6151
R745 B.n140 B.n139 10.6151
R746 B.n139 B.n110 10.6151
R747 B.n135 B.n110 10.6151
R748 B.n135 B.n134 10.6151
R749 B.n134 B.n133 10.6151
R750 B.n133 B.n112 10.6151
R751 B.n129 B.n112 10.6151
R752 B.n129 B.n128 10.6151
R753 B.n128 B.n127 10.6151
R754 B.n127 B.n114 10.6151
R755 B.n123 B.n114 10.6151
R756 B.n123 B.n122 10.6151
R757 B.n122 B.n121 10.6151
R758 B.n121 B.n116 10.6151
R759 B.n117 B.n116 10.6151
R760 B.n117 B.n0 10.6151
R761 B.n435 B.n1 10.6151
R762 B.n435 B.n434 10.6151
R763 B.n434 B.n433 10.6151
R764 B.n433 B.n4 10.6151
R765 B.n429 B.n4 10.6151
R766 B.n429 B.n428 10.6151
R767 B.n428 B.n427 10.6151
R768 B.n427 B.n6 10.6151
R769 B.n423 B.n6 10.6151
R770 B.n423 B.n422 10.6151
R771 B.n422 B.n421 10.6151
R772 B.n421 B.n8 10.6151
R773 B.n417 B.n8 10.6151
R774 B.n417 B.n416 10.6151
R775 B.n416 B.n415 10.6151
R776 B.n415 B.n10 10.6151
R777 B.n411 B.n10 10.6151
R778 B.n411 B.n410 10.6151
R779 B.n410 B.n409 10.6151
R780 B.n409 B.n12 10.6151
R781 B.n405 B.n12 10.6151
R782 B.n405 B.n404 10.6151
R783 B.n404 B.n403 10.6151
R784 B.n403 B.n14 10.6151
R785 B.n399 B.n14 10.6151
R786 B.n399 B.n398 10.6151
R787 B.n398 B.n397 10.6151
R788 B.n397 B.n16 10.6151
R789 B.n393 B.n16 10.6151
R790 B.n393 B.n392 10.6151
R791 B.n392 B.n391 10.6151
R792 B.n391 B.n18 10.6151
R793 B.n387 B.n18 10.6151
R794 B.n387 B.n386 10.6151
R795 B.n386 B.n385 10.6151
R796 B.n385 B.n20 10.6151
R797 B.n367 B.n28 9.36635
R798 B.n350 B.n349 9.36635
R799 B.n188 B.n187 9.36635
R800 B.n205 B.n86 9.36635
R801 B.n439 B.n0 2.81026
R802 B.n439 B.n1 2.81026
R803 B.n364 B.n28 1.24928
R804 B.n351 B.n350 1.24928
R805 B.n189 B.n188 1.24928
R806 B.n202 B.n86 1.24928
C0 VTAIL w_n2938_n1294# 1.41187f
C1 B VN 0.925515f
C2 VTAIL VDD2 3.68761f
C3 VTAIL VDD1 3.63761f
C4 VP VTAIL 1.94673f
C5 VDD2 w_n2938_n1294# 1.51342f
C6 VDD1 w_n2938_n1294# 1.44416f
C7 VP w_n2938_n1294# 5.61261f
C8 VDD2 VDD1 1.22308f
C9 VP VDD2 0.425691f
C10 VP VDD1 1.46814f
C11 VTAIL VN 1.9326f
C12 VN w_n2938_n1294# 5.23988f
C13 VTAIL B 1.15198f
C14 B w_n2938_n1294# 6.15189f
C15 VN VDD2 1.20211f
C16 VN VDD1 0.157111f
C17 VP VN 4.55542f
C18 B VDD2 1.22104f
C19 B VDD1 1.15785f
C20 VP B 1.55424f
C21 VDD2 VSUBS 0.956195f
C22 VDD1 VSUBS 1.338434f
C23 VTAIL VSUBS 0.385182f
C24 VN VSUBS 4.8486f
C25 VP VSUBS 2.013789f
C26 B VSUBS 3.105719f
C27 w_n2938_n1294# VSUBS 48.6885f
C28 B.n0 VSUBS 0.005896f
C29 B.n1 VSUBS 0.005896f
C30 B.n2 VSUBS 0.009324f
C31 B.n3 VSUBS 0.009324f
C32 B.n4 VSUBS 0.009324f
C33 B.n5 VSUBS 0.009324f
C34 B.n6 VSUBS 0.009324f
C35 B.n7 VSUBS 0.009324f
C36 B.n8 VSUBS 0.009324f
C37 B.n9 VSUBS 0.009324f
C38 B.n10 VSUBS 0.009324f
C39 B.n11 VSUBS 0.009324f
C40 B.n12 VSUBS 0.009324f
C41 B.n13 VSUBS 0.009324f
C42 B.n14 VSUBS 0.009324f
C43 B.n15 VSUBS 0.009324f
C44 B.n16 VSUBS 0.009324f
C45 B.n17 VSUBS 0.009324f
C46 B.n18 VSUBS 0.009324f
C47 B.n19 VSUBS 0.009324f
C48 B.n20 VSUBS 0.020855f
C49 B.n21 VSUBS 0.009324f
C50 B.n22 VSUBS 0.009324f
C51 B.n23 VSUBS 0.009324f
C52 B.n24 VSUBS 0.009324f
C53 B.n25 VSUBS 0.009324f
C54 B.t11 VSUBS 0.044604f
C55 B.t10 VSUBS 0.053672f
C56 B.t9 VSUBS 0.228889f
C57 B.n26 VSUBS 0.085323f
C58 B.n27 VSUBS 0.069926f
C59 B.n28 VSUBS 0.021602f
C60 B.n29 VSUBS 0.009324f
C61 B.n30 VSUBS 0.009324f
C62 B.n31 VSUBS 0.009324f
C63 B.n32 VSUBS 0.009324f
C64 B.n33 VSUBS 0.009324f
C65 B.t8 VSUBS 0.044604f
C66 B.t7 VSUBS 0.053672f
C67 B.t6 VSUBS 0.228889f
C68 B.n34 VSUBS 0.085323f
C69 B.n35 VSUBS 0.069926f
C70 B.n36 VSUBS 0.009324f
C71 B.n37 VSUBS 0.009324f
C72 B.n38 VSUBS 0.009324f
C73 B.n39 VSUBS 0.009324f
C74 B.n40 VSUBS 0.009324f
C75 B.n41 VSUBS 0.020855f
C76 B.n42 VSUBS 0.009324f
C77 B.n43 VSUBS 0.009324f
C78 B.n44 VSUBS 0.009324f
C79 B.n45 VSUBS 0.009324f
C80 B.n46 VSUBS 0.009324f
C81 B.n47 VSUBS 0.009324f
C82 B.n48 VSUBS 0.009324f
C83 B.n49 VSUBS 0.009324f
C84 B.n50 VSUBS 0.009324f
C85 B.n51 VSUBS 0.009324f
C86 B.n52 VSUBS 0.009324f
C87 B.n53 VSUBS 0.009324f
C88 B.n54 VSUBS 0.009324f
C89 B.n55 VSUBS 0.009324f
C90 B.n56 VSUBS 0.009324f
C91 B.n57 VSUBS 0.009324f
C92 B.n58 VSUBS 0.009324f
C93 B.n59 VSUBS 0.009324f
C94 B.n60 VSUBS 0.009324f
C95 B.n61 VSUBS 0.009324f
C96 B.n62 VSUBS 0.009324f
C97 B.n63 VSUBS 0.009324f
C98 B.n64 VSUBS 0.009324f
C99 B.n65 VSUBS 0.009324f
C100 B.n66 VSUBS 0.009324f
C101 B.n67 VSUBS 0.009324f
C102 B.n68 VSUBS 0.009324f
C103 B.n69 VSUBS 0.009324f
C104 B.n70 VSUBS 0.009324f
C105 B.n71 VSUBS 0.009324f
C106 B.n72 VSUBS 0.009324f
C107 B.n73 VSUBS 0.009324f
C108 B.n74 VSUBS 0.009324f
C109 B.n75 VSUBS 0.009324f
C110 B.n76 VSUBS 0.009324f
C111 B.n77 VSUBS 0.009324f
C112 B.n78 VSUBS 0.020855f
C113 B.n79 VSUBS 0.009324f
C114 B.n80 VSUBS 0.009324f
C115 B.n81 VSUBS 0.009324f
C116 B.n82 VSUBS 0.009324f
C117 B.n83 VSUBS 0.009324f
C118 B.t1 VSUBS 0.044604f
C119 B.t2 VSUBS 0.053672f
C120 B.t0 VSUBS 0.228889f
C121 B.n84 VSUBS 0.085323f
C122 B.n85 VSUBS 0.069926f
C123 B.n86 VSUBS 0.021602f
C124 B.n87 VSUBS 0.009324f
C125 B.n88 VSUBS 0.009324f
C126 B.n89 VSUBS 0.009324f
C127 B.n90 VSUBS 0.009324f
C128 B.n91 VSUBS 0.009324f
C129 B.t4 VSUBS 0.044604f
C130 B.t5 VSUBS 0.053672f
C131 B.t3 VSUBS 0.228889f
C132 B.n92 VSUBS 0.085323f
C133 B.n93 VSUBS 0.069926f
C134 B.n94 VSUBS 0.009324f
C135 B.n95 VSUBS 0.009324f
C136 B.n96 VSUBS 0.009324f
C137 B.n97 VSUBS 0.009324f
C138 B.n98 VSUBS 0.009324f
C139 B.n99 VSUBS 0.020855f
C140 B.n100 VSUBS 0.009324f
C141 B.n101 VSUBS 0.009324f
C142 B.n102 VSUBS 0.009324f
C143 B.n103 VSUBS 0.009324f
C144 B.n104 VSUBS 0.009324f
C145 B.n105 VSUBS 0.009324f
C146 B.n106 VSUBS 0.009324f
C147 B.n107 VSUBS 0.009324f
C148 B.n108 VSUBS 0.009324f
C149 B.n109 VSUBS 0.009324f
C150 B.n110 VSUBS 0.009324f
C151 B.n111 VSUBS 0.009324f
C152 B.n112 VSUBS 0.009324f
C153 B.n113 VSUBS 0.009324f
C154 B.n114 VSUBS 0.009324f
C155 B.n115 VSUBS 0.009324f
C156 B.n116 VSUBS 0.009324f
C157 B.n117 VSUBS 0.009324f
C158 B.n118 VSUBS 0.009324f
C159 B.n119 VSUBS 0.009324f
C160 B.n120 VSUBS 0.009324f
C161 B.n121 VSUBS 0.009324f
C162 B.n122 VSUBS 0.009324f
C163 B.n123 VSUBS 0.009324f
C164 B.n124 VSUBS 0.009324f
C165 B.n125 VSUBS 0.009324f
C166 B.n126 VSUBS 0.009324f
C167 B.n127 VSUBS 0.009324f
C168 B.n128 VSUBS 0.009324f
C169 B.n129 VSUBS 0.009324f
C170 B.n130 VSUBS 0.009324f
C171 B.n131 VSUBS 0.009324f
C172 B.n132 VSUBS 0.009324f
C173 B.n133 VSUBS 0.009324f
C174 B.n134 VSUBS 0.009324f
C175 B.n135 VSUBS 0.009324f
C176 B.n136 VSUBS 0.009324f
C177 B.n137 VSUBS 0.009324f
C178 B.n138 VSUBS 0.009324f
C179 B.n139 VSUBS 0.009324f
C180 B.n140 VSUBS 0.009324f
C181 B.n141 VSUBS 0.009324f
C182 B.n142 VSUBS 0.009324f
C183 B.n143 VSUBS 0.009324f
C184 B.n144 VSUBS 0.009324f
C185 B.n145 VSUBS 0.009324f
C186 B.n146 VSUBS 0.009324f
C187 B.n147 VSUBS 0.009324f
C188 B.n148 VSUBS 0.009324f
C189 B.n149 VSUBS 0.009324f
C190 B.n150 VSUBS 0.009324f
C191 B.n151 VSUBS 0.009324f
C192 B.n152 VSUBS 0.009324f
C193 B.n153 VSUBS 0.009324f
C194 B.n154 VSUBS 0.009324f
C195 B.n155 VSUBS 0.009324f
C196 B.n156 VSUBS 0.009324f
C197 B.n157 VSUBS 0.009324f
C198 B.n158 VSUBS 0.009324f
C199 B.n159 VSUBS 0.009324f
C200 B.n160 VSUBS 0.009324f
C201 B.n161 VSUBS 0.009324f
C202 B.n162 VSUBS 0.009324f
C203 B.n163 VSUBS 0.009324f
C204 B.n164 VSUBS 0.009324f
C205 B.n165 VSUBS 0.009324f
C206 B.n166 VSUBS 0.009324f
C207 B.n167 VSUBS 0.009324f
C208 B.n168 VSUBS 0.009324f
C209 B.n169 VSUBS 0.009324f
C210 B.n170 VSUBS 0.020855f
C211 B.n171 VSUBS 0.022199f
C212 B.n172 VSUBS 0.022199f
C213 B.n173 VSUBS 0.009324f
C214 B.n174 VSUBS 0.009324f
C215 B.n175 VSUBS 0.009324f
C216 B.n176 VSUBS 0.009324f
C217 B.n177 VSUBS 0.009324f
C218 B.n178 VSUBS 0.009324f
C219 B.n179 VSUBS 0.009324f
C220 B.n180 VSUBS 0.009324f
C221 B.n181 VSUBS 0.009324f
C222 B.n182 VSUBS 0.009324f
C223 B.n183 VSUBS 0.009324f
C224 B.n184 VSUBS 0.009324f
C225 B.n185 VSUBS 0.009324f
C226 B.n186 VSUBS 0.009324f
C227 B.n187 VSUBS 0.008775f
C228 B.n188 VSUBS 0.021602f
C229 B.n189 VSUBS 0.00521f
C230 B.n190 VSUBS 0.009324f
C231 B.n191 VSUBS 0.009324f
C232 B.n192 VSUBS 0.009324f
C233 B.n193 VSUBS 0.009324f
C234 B.n194 VSUBS 0.009324f
C235 B.n195 VSUBS 0.009324f
C236 B.n196 VSUBS 0.009324f
C237 B.n197 VSUBS 0.009324f
C238 B.n198 VSUBS 0.009324f
C239 B.n199 VSUBS 0.009324f
C240 B.n200 VSUBS 0.009324f
C241 B.n201 VSUBS 0.009324f
C242 B.n202 VSUBS 0.00521f
C243 B.n203 VSUBS 0.009324f
C244 B.n204 VSUBS 0.009324f
C245 B.n205 VSUBS 0.008775f
C246 B.n206 VSUBS 0.009324f
C247 B.n207 VSUBS 0.009324f
C248 B.n208 VSUBS 0.009324f
C249 B.n209 VSUBS 0.009324f
C250 B.n210 VSUBS 0.009324f
C251 B.n211 VSUBS 0.009324f
C252 B.n212 VSUBS 0.009324f
C253 B.n213 VSUBS 0.009324f
C254 B.n214 VSUBS 0.009324f
C255 B.n215 VSUBS 0.009324f
C256 B.n216 VSUBS 0.009324f
C257 B.n217 VSUBS 0.009324f
C258 B.n218 VSUBS 0.009324f
C259 B.n219 VSUBS 0.022199f
C260 B.n220 VSUBS 0.022199f
C261 B.n221 VSUBS 0.020855f
C262 B.n222 VSUBS 0.009324f
C263 B.n223 VSUBS 0.009324f
C264 B.n224 VSUBS 0.009324f
C265 B.n225 VSUBS 0.009324f
C266 B.n226 VSUBS 0.009324f
C267 B.n227 VSUBS 0.009324f
C268 B.n228 VSUBS 0.009324f
C269 B.n229 VSUBS 0.009324f
C270 B.n230 VSUBS 0.009324f
C271 B.n231 VSUBS 0.009324f
C272 B.n232 VSUBS 0.009324f
C273 B.n233 VSUBS 0.009324f
C274 B.n234 VSUBS 0.009324f
C275 B.n235 VSUBS 0.009324f
C276 B.n236 VSUBS 0.009324f
C277 B.n237 VSUBS 0.009324f
C278 B.n238 VSUBS 0.009324f
C279 B.n239 VSUBS 0.009324f
C280 B.n240 VSUBS 0.009324f
C281 B.n241 VSUBS 0.009324f
C282 B.n242 VSUBS 0.009324f
C283 B.n243 VSUBS 0.009324f
C284 B.n244 VSUBS 0.009324f
C285 B.n245 VSUBS 0.009324f
C286 B.n246 VSUBS 0.009324f
C287 B.n247 VSUBS 0.009324f
C288 B.n248 VSUBS 0.009324f
C289 B.n249 VSUBS 0.009324f
C290 B.n250 VSUBS 0.009324f
C291 B.n251 VSUBS 0.009324f
C292 B.n252 VSUBS 0.009324f
C293 B.n253 VSUBS 0.009324f
C294 B.n254 VSUBS 0.009324f
C295 B.n255 VSUBS 0.009324f
C296 B.n256 VSUBS 0.009324f
C297 B.n257 VSUBS 0.009324f
C298 B.n258 VSUBS 0.009324f
C299 B.n259 VSUBS 0.009324f
C300 B.n260 VSUBS 0.009324f
C301 B.n261 VSUBS 0.009324f
C302 B.n262 VSUBS 0.009324f
C303 B.n263 VSUBS 0.009324f
C304 B.n264 VSUBS 0.009324f
C305 B.n265 VSUBS 0.009324f
C306 B.n266 VSUBS 0.009324f
C307 B.n267 VSUBS 0.009324f
C308 B.n268 VSUBS 0.009324f
C309 B.n269 VSUBS 0.009324f
C310 B.n270 VSUBS 0.009324f
C311 B.n271 VSUBS 0.009324f
C312 B.n272 VSUBS 0.009324f
C313 B.n273 VSUBS 0.009324f
C314 B.n274 VSUBS 0.009324f
C315 B.n275 VSUBS 0.009324f
C316 B.n276 VSUBS 0.009324f
C317 B.n277 VSUBS 0.009324f
C318 B.n278 VSUBS 0.009324f
C319 B.n279 VSUBS 0.009324f
C320 B.n280 VSUBS 0.009324f
C321 B.n281 VSUBS 0.009324f
C322 B.n282 VSUBS 0.009324f
C323 B.n283 VSUBS 0.009324f
C324 B.n284 VSUBS 0.009324f
C325 B.n285 VSUBS 0.009324f
C326 B.n286 VSUBS 0.009324f
C327 B.n287 VSUBS 0.009324f
C328 B.n288 VSUBS 0.009324f
C329 B.n289 VSUBS 0.009324f
C330 B.n290 VSUBS 0.009324f
C331 B.n291 VSUBS 0.009324f
C332 B.n292 VSUBS 0.009324f
C333 B.n293 VSUBS 0.009324f
C334 B.n294 VSUBS 0.009324f
C335 B.n295 VSUBS 0.009324f
C336 B.n296 VSUBS 0.009324f
C337 B.n297 VSUBS 0.009324f
C338 B.n298 VSUBS 0.009324f
C339 B.n299 VSUBS 0.009324f
C340 B.n300 VSUBS 0.009324f
C341 B.n301 VSUBS 0.009324f
C342 B.n302 VSUBS 0.009324f
C343 B.n303 VSUBS 0.009324f
C344 B.n304 VSUBS 0.009324f
C345 B.n305 VSUBS 0.009324f
C346 B.n306 VSUBS 0.009324f
C347 B.n307 VSUBS 0.009324f
C348 B.n308 VSUBS 0.009324f
C349 B.n309 VSUBS 0.009324f
C350 B.n310 VSUBS 0.009324f
C351 B.n311 VSUBS 0.009324f
C352 B.n312 VSUBS 0.009324f
C353 B.n313 VSUBS 0.009324f
C354 B.n314 VSUBS 0.009324f
C355 B.n315 VSUBS 0.009324f
C356 B.n316 VSUBS 0.009324f
C357 B.n317 VSUBS 0.009324f
C358 B.n318 VSUBS 0.009324f
C359 B.n319 VSUBS 0.009324f
C360 B.n320 VSUBS 0.009324f
C361 B.n321 VSUBS 0.009324f
C362 B.n322 VSUBS 0.009324f
C363 B.n323 VSUBS 0.009324f
C364 B.n324 VSUBS 0.009324f
C365 B.n325 VSUBS 0.009324f
C366 B.n326 VSUBS 0.009324f
C367 B.n327 VSUBS 0.009324f
C368 B.n328 VSUBS 0.009324f
C369 B.n329 VSUBS 0.009324f
C370 B.n330 VSUBS 0.009324f
C371 B.n331 VSUBS 0.009324f
C372 B.n332 VSUBS 0.02198f
C373 B.n333 VSUBS 0.021075f
C374 B.n334 VSUBS 0.022199f
C375 B.n335 VSUBS 0.009324f
C376 B.n336 VSUBS 0.009324f
C377 B.n337 VSUBS 0.009324f
C378 B.n338 VSUBS 0.009324f
C379 B.n339 VSUBS 0.009324f
C380 B.n340 VSUBS 0.009324f
C381 B.n341 VSUBS 0.009324f
C382 B.n342 VSUBS 0.009324f
C383 B.n343 VSUBS 0.009324f
C384 B.n344 VSUBS 0.009324f
C385 B.n345 VSUBS 0.009324f
C386 B.n346 VSUBS 0.009324f
C387 B.n347 VSUBS 0.009324f
C388 B.n348 VSUBS 0.009324f
C389 B.n349 VSUBS 0.008775f
C390 B.n350 VSUBS 0.021602f
C391 B.n351 VSUBS 0.00521f
C392 B.n352 VSUBS 0.009324f
C393 B.n353 VSUBS 0.009324f
C394 B.n354 VSUBS 0.009324f
C395 B.n355 VSUBS 0.009324f
C396 B.n356 VSUBS 0.009324f
C397 B.n357 VSUBS 0.009324f
C398 B.n358 VSUBS 0.009324f
C399 B.n359 VSUBS 0.009324f
C400 B.n360 VSUBS 0.009324f
C401 B.n361 VSUBS 0.009324f
C402 B.n362 VSUBS 0.009324f
C403 B.n363 VSUBS 0.009324f
C404 B.n364 VSUBS 0.00521f
C405 B.n365 VSUBS 0.009324f
C406 B.n366 VSUBS 0.009324f
C407 B.n367 VSUBS 0.008775f
C408 B.n368 VSUBS 0.009324f
C409 B.n369 VSUBS 0.009324f
C410 B.n370 VSUBS 0.009324f
C411 B.n371 VSUBS 0.009324f
C412 B.n372 VSUBS 0.009324f
C413 B.n373 VSUBS 0.009324f
C414 B.n374 VSUBS 0.009324f
C415 B.n375 VSUBS 0.009324f
C416 B.n376 VSUBS 0.009324f
C417 B.n377 VSUBS 0.009324f
C418 B.n378 VSUBS 0.009324f
C419 B.n379 VSUBS 0.009324f
C420 B.n380 VSUBS 0.009324f
C421 B.n381 VSUBS 0.022199f
C422 B.n382 VSUBS 0.022199f
C423 B.n383 VSUBS 0.020855f
C424 B.n384 VSUBS 0.009324f
C425 B.n385 VSUBS 0.009324f
C426 B.n386 VSUBS 0.009324f
C427 B.n387 VSUBS 0.009324f
C428 B.n388 VSUBS 0.009324f
C429 B.n389 VSUBS 0.009324f
C430 B.n390 VSUBS 0.009324f
C431 B.n391 VSUBS 0.009324f
C432 B.n392 VSUBS 0.009324f
C433 B.n393 VSUBS 0.009324f
C434 B.n394 VSUBS 0.009324f
C435 B.n395 VSUBS 0.009324f
C436 B.n396 VSUBS 0.009324f
C437 B.n397 VSUBS 0.009324f
C438 B.n398 VSUBS 0.009324f
C439 B.n399 VSUBS 0.009324f
C440 B.n400 VSUBS 0.009324f
C441 B.n401 VSUBS 0.009324f
C442 B.n402 VSUBS 0.009324f
C443 B.n403 VSUBS 0.009324f
C444 B.n404 VSUBS 0.009324f
C445 B.n405 VSUBS 0.009324f
C446 B.n406 VSUBS 0.009324f
C447 B.n407 VSUBS 0.009324f
C448 B.n408 VSUBS 0.009324f
C449 B.n409 VSUBS 0.009324f
C450 B.n410 VSUBS 0.009324f
C451 B.n411 VSUBS 0.009324f
C452 B.n412 VSUBS 0.009324f
C453 B.n413 VSUBS 0.009324f
C454 B.n414 VSUBS 0.009324f
C455 B.n415 VSUBS 0.009324f
C456 B.n416 VSUBS 0.009324f
C457 B.n417 VSUBS 0.009324f
C458 B.n418 VSUBS 0.009324f
C459 B.n419 VSUBS 0.009324f
C460 B.n420 VSUBS 0.009324f
C461 B.n421 VSUBS 0.009324f
C462 B.n422 VSUBS 0.009324f
C463 B.n423 VSUBS 0.009324f
C464 B.n424 VSUBS 0.009324f
C465 B.n425 VSUBS 0.009324f
C466 B.n426 VSUBS 0.009324f
C467 B.n427 VSUBS 0.009324f
C468 B.n428 VSUBS 0.009324f
C469 B.n429 VSUBS 0.009324f
C470 B.n430 VSUBS 0.009324f
C471 B.n431 VSUBS 0.009324f
C472 B.n432 VSUBS 0.009324f
C473 B.n433 VSUBS 0.009324f
C474 B.n434 VSUBS 0.009324f
C475 B.n435 VSUBS 0.009324f
C476 B.n436 VSUBS 0.009324f
C477 B.n437 VSUBS 0.009324f
C478 B.n438 VSUBS 0.009324f
C479 B.n439 VSUBS 0.021112f
C480 VDD1.t2 VSUBS 0.130378f
C481 VDD1.t3 VSUBS 0.130233f
C482 VDD1.t5 VSUBS 0.021229f
C483 VDD1.t4 VSUBS 0.021229f
C484 VDD1.n0 VSUBS 0.080046f
C485 VDD1.n1 VSUBS 1.47407f
C486 VDD1.t1 VSUBS 0.021229f
C487 VDD1.t0 VSUBS 0.021229f
C488 VDD1.n2 VSUBS 0.079457f
C489 VDD1.n3 VSUBS 1.24261f
C490 VP.n0 VSUBS 0.063111f
C491 VP.t1 VSUBS 0.370516f
C492 VP.n1 VSUBS 0.067213f
C493 VP.n2 VSUBS 0.047869f
C494 VP.t0 VSUBS 0.370516f
C495 VP.n3 VSUBS 0.067213f
C496 VP.n4 VSUBS 0.063111f
C497 VP.t2 VSUBS 0.370516f
C498 VP.n5 VSUBS 0.063111f
C499 VP.t5 VSUBS 0.370516f
C500 VP.n6 VSUBS 0.067213f
C501 VP.t3 VSUBS 0.673901f
C502 VP.n7 VSUBS 0.292403f
C503 VP.t4 VSUBS 0.370516f
C504 VP.n8 VSUBS 0.344629f
C505 VP.n9 VSUBS 0.089217f
C506 VP.n10 VSUBS 0.403577f
C507 VP.n11 VSUBS 0.047869f
C508 VP.n12 VSUBS 0.047869f
C509 VP.n13 VSUBS 0.072549f
C510 VP.n14 VSUBS 0.085693f
C511 VP.n15 VSUBS 0.3638f
C512 VP.n16 VSUBS 1.78512f
C513 VP.n17 VSUBS 1.82915f
C514 VP.n18 VSUBS 0.3638f
C515 VP.n19 VSUBS 0.085693f
C516 VP.n20 VSUBS 0.072549f
C517 VP.n21 VSUBS 0.047869f
C518 VP.n22 VSUBS 0.047869f
C519 VP.n23 VSUBS 0.047869f
C520 VP.n24 VSUBS 0.089217f
C521 VP.n25 VSUBS 0.244471f
C522 VP.n26 VSUBS 0.089217f
C523 VP.n27 VSUBS 0.047869f
C524 VP.n28 VSUBS 0.047869f
C525 VP.n29 VSUBS 0.047869f
C526 VP.n30 VSUBS 0.072549f
C527 VP.n31 VSUBS 0.085693f
C528 VP.n32 VSUBS 0.3638f
C529 VP.n33 VSUBS 0.054824f
C530 VDD2.t1 VSUBS 0.136153f
C531 VDD2.t4 VSUBS 0.022194f
C532 VDD2.t5 VSUBS 0.022194f
C533 VDD2.n0 VSUBS 0.083685f
C534 VDD2.n1 VSUBS 1.47089f
C535 VDD2.t0 VSUBS 0.134602f
C536 VDD2.n2 VSUBS 1.26224f
C537 VDD2.t2 VSUBS 0.022194f
C538 VDD2.t3 VSUBS 0.022194f
C539 VDD2.n3 VSUBS 0.08368f
C540 VTAIL.t10 VSUBS 0.02941f
C541 VTAIL.t9 VSUBS 0.02941f
C542 VTAIL.n0 VSUBS 0.094037f
C543 VTAIL.n1 VSUBS 0.368725f
C544 VTAIL.t4 VSUBS 0.162802f
C545 VTAIL.n2 VSUBS 0.492902f
C546 VTAIL.t2 VSUBS 0.02941f
C547 VTAIL.t3 VSUBS 0.02941f
C548 VTAIL.n3 VSUBS 0.094037f
C549 VTAIL.n4 VSUBS 1.09445f
C550 VTAIL.t11 VSUBS 0.02941f
C551 VTAIL.t7 VSUBS 0.02941f
C552 VTAIL.n5 VSUBS 0.094037f
C553 VTAIL.n6 VSUBS 1.09445f
C554 VTAIL.t8 VSUBS 0.162802f
C555 VTAIL.n7 VSUBS 0.492901f
C556 VTAIL.t5 VSUBS 0.02941f
C557 VTAIL.t1 VSUBS 0.02941f
C558 VTAIL.n8 VSUBS 0.094037f
C559 VTAIL.n9 VSUBS 0.481458f
C560 VTAIL.t0 VSUBS 0.162802f
C561 VTAIL.n10 VSUBS 0.949873f
C562 VTAIL.t6 VSUBS 0.162802f
C563 VTAIL.n11 VSUBS 0.906587f
C564 VN.n0 VSUBS 0.060239f
C565 VN.t0 VSUBS 0.353653f
C566 VN.n1 VSUBS 0.064154f
C567 VN.t4 VSUBS 0.64323f
C568 VN.n2 VSUBS 0.279095f
C569 VN.t1 VSUBS 0.353653f
C570 VN.n3 VSUBS 0.328944f
C571 VN.n4 VSUBS 0.085156f
C572 VN.n5 VSUBS 0.385209f
C573 VN.n6 VSUBS 0.045691f
C574 VN.n7 VSUBS 0.045691f
C575 VN.n8 VSUBS 0.069247f
C576 VN.n9 VSUBS 0.081793f
C577 VN.n10 VSUBS 0.347242f
C578 VN.n11 VSUBS 0.052328f
C579 VN.n12 VSUBS 0.060239f
C580 VN.t5 VSUBS 0.353653f
C581 VN.n13 VSUBS 0.064154f
C582 VN.t2 VSUBS 0.64323f
C583 VN.n14 VSUBS 0.279095f
C584 VN.t3 VSUBS 0.353653f
C585 VN.n15 VSUBS 0.328944f
C586 VN.n16 VSUBS 0.085156f
C587 VN.n17 VSUBS 0.385209f
C588 VN.n18 VSUBS 0.045691f
C589 VN.n19 VSUBS 0.045691f
C590 VN.n20 VSUBS 0.069247f
C591 VN.n21 VSUBS 0.081793f
C592 VN.n22 VSUBS 0.347242f
C593 VN.n23 VSUBS 1.72951f
.ends

