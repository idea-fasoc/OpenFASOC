* NGSPICE file created from diff_pair_sample_1006.ext - technology: sky130A

.subckt diff_pair_sample_1006 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t5 VP.t0 VTAIL.t9 w_n1682_n4180# sky130_fd_pr__pfet_01v8 ad=6.2634 pd=32.9 as=2.6499 ps=16.39 w=16.06 l=0.56
X1 VDD1.t4 VP.t1 VTAIL.t10 w_n1682_n4180# sky130_fd_pr__pfet_01v8 ad=6.2634 pd=32.9 as=2.6499 ps=16.39 w=16.06 l=0.56
X2 VDD1.t3 VP.t2 VTAIL.t6 w_n1682_n4180# sky130_fd_pr__pfet_01v8 ad=2.6499 pd=16.39 as=6.2634 ps=32.9 w=16.06 l=0.56
X3 B.t11 B.t9 B.t10 w_n1682_n4180# sky130_fd_pr__pfet_01v8 ad=6.2634 pd=32.9 as=0 ps=0 w=16.06 l=0.56
X4 VTAIL.t11 VP.t3 VDD1.t2 w_n1682_n4180# sky130_fd_pr__pfet_01v8 ad=2.6499 pd=16.39 as=2.6499 ps=16.39 w=16.06 l=0.56
X5 VDD2.t5 VN.t0 VTAIL.t3 w_n1682_n4180# sky130_fd_pr__pfet_01v8 ad=6.2634 pd=32.9 as=2.6499 ps=16.39 w=16.06 l=0.56
X6 VDD1.t1 VP.t4 VTAIL.t8 w_n1682_n4180# sky130_fd_pr__pfet_01v8 ad=2.6499 pd=16.39 as=6.2634 ps=32.9 w=16.06 l=0.56
X7 VDD2.t4 VN.t1 VTAIL.t4 w_n1682_n4180# sky130_fd_pr__pfet_01v8 ad=2.6499 pd=16.39 as=6.2634 ps=32.9 w=16.06 l=0.56
X8 B.t8 B.t6 B.t7 w_n1682_n4180# sky130_fd_pr__pfet_01v8 ad=6.2634 pd=32.9 as=0 ps=0 w=16.06 l=0.56
X9 B.t5 B.t3 B.t4 w_n1682_n4180# sky130_fd_pr__pfet_01v8 ad=6.2634 pd=32.9 as=0 ps=0 w=16.06 l=0.56
X10 VTAIL.t5 VN.t2 VDD2.t3 w_n1682_n4180# sky130_fd_pr__pfet_01v8 ad=2.6499 pd=16.39 as=2.6499 ps=16.39 w=16.06 l=0.56
X11 VTAIL.t7 VP.t5 VDD1.t0 w_n1682_n4180# sky130_fd_pr__pfet_01v8 ad=2.6499 pd=16.39 as=2.6499 ps=16.39 w=16.06 l=0.56
X12 VDD2.t2 VN.t3 VTAIL.t2 w_n1682_n4180# sky130_fd_pr__pfet_01v8 ad=6.2634 pd=32.9 as=2.6499 ps=16.39 w=16.06 l=0.56
X13 VDD2.t1 VN.t4 VTAIL.t0 w_n1682_n4180# sky130_fd_pr__pfet_01v8 ad=2.6499 pd=16.39 as=6.2634 ps=32.9 w=16.06 l=0.56
X14 B.t2 B.t0 B.t1 w_n1682_n4180# sky130_fd_pr__pfet_01v8 ad=6.2634 pd=32.9 as=0 ps=0 w=16.06 l=0.56
X15 VTAIL.t1 VN.t5 VDD2.t0 w_n1682_n4180# sky130_fd_pr__pfet_01v8 ad=2.6499 pd=16.39 as=2.6499 ps=16.39 w=16.06 l=0.56
R0 VP.n1 VP.t0 788.124
R1 VP.n6 VP.t1 761.303
R2 VP.n7 VP.t3 761.303
R3 VP.n8 VP.t4 761.303
R4 VP.n3 VP.t2 761.303
R5 VP.n2 VP.t5 761.303
R6 VP.n9 VP.n8 161.3
R7 VP.n4 VP.n3 161.3
R8 VP.n6 VP.n5 161.3
R9 VP.n7 VP.n0 80.6037
R10 VP.n7 VP.n6 48.2005
R11 VP.n8 VP.n7 48.2005
R12 VP.n3 VP.n2 48.2005
R13 VP.n4 VP.n1 45.1367
R14 VP.n5 VP.n4 43.777
R15 VP.n2 VP.n1 13.3799
R16 VP.n5 VP.n0 0.285035
R17 VP.n9 VP.n0 0.285035
R18 VP VP.n9 0.0516364
R19 VTAIL.n362 VTAIL.n278 756.745
R20 VTAIL.n86 VTAIL.n2 756.745
R21 VTAIL.n272 VTAIL.n188 756.745
R22 VTAIL.n180 VTAIL.n96 756.745
R23 VTAIL.n306 VTAIL.n305 585
R24 VTAIL.n311 VTAIL.n310 585
R25 VTAIL.n313 VTAIL.n312 585
R26 VTAIL.n302 VTAIL.n301 585
R27 VTAIL.n319 VTAIL.n318 585
R28 VTAIL.n321 VTAIL.n320 585
R29 VTAIL.n298 VTAIL.n297 585
R30 VTAIL.n327 VTAIL.n326 585
R31 VTAIL.n329 VTAIL.n328 585
R32 VTAIL.n294 VTAIL.n293 585
R33 VTAIL.n335 VTAIL.n334 585
R34 VTAIL.n337 VTAIL.n336 585
R35 VTAIL.n290 VTAIL.n289 585
R36 VTAIL.n343 VTAIL.n342 585
R37 VTAIL.n345 VTAIL.n344 585
R38 VTAIL.n286 VTAIL.n285 585
R39 VTAIL.n352 VTAIL.n351 585
R40 VTAIL.n353 VTAIL.n284 585
R41 VTAIL.n355 VTAIL.n354 585
R42 VTAIL.n282 VTAIL.n281 585
R43 VTAIL.n361 VTAIL.n360 585
R44 VTAIL.n363 VTAIL.n362 585
R45 VTAIL.n30 VTAIL.n29 585
R46 VTAIL.n35 VTAIL.n34 585
R47 VTAIL.n37 VTAIL.n36 585
R48 VTAIL.n26 VTAIL.n25 585
R49 VTAIL.n43 VTAIL.n42 585
R50 VTAIL.n45 VTAIL.n44 585
R51 VTAIL.n22 VTAIL.n21 585
R52 VTAIL.n51 VTAIL.n50 585
R53 VTAIL.n53 VTAIL.n52 585
R54 VTAIL.n18 VTAIL.n17 585
R55 VTAIL.n59 VTAIL.n58 585
R56 VTAIL.n61 VTAIL.n60 585
R57 VTAIL.n14 VTAIL.n13 585
R58 VTAIL.n67 VTAIL.n66 585
R59 VTAIL.n69 VTAIL.n68 585
R60 VTAIL.n10 VTAIL.n9 585
R61 VTAIL.n76 VTAIL.n75 585
R62 VTAIL.n77 VTAIL.n8 585
R63 VTAIL.n79 VTAIL.n78 585
R64 VTAIL.n6 VTAIL.n5 585
R65 VTAIL.n85 VTAIL.n84 585
R66 VTAIL.n87 VTAIL.n86 585
R67 VTAIL.n273 VTAIL.n272 585
R68 VTAIL.n271 VTAIL.n270 585
R69 VTAIL.n192 VTAIL.n191 585
R70 VTAIL.n265 VTAIL.n264 585
R71 VTAIL.n263 VTAIL.n194 585
R72 VTAIL.n262 VTAIL.n261 585
R73 VTAIL.n197 VTAIL.n195 585
R74 VTAIL.n256 VTAIL.n255 585
R75 VTAIL.n254 VTAIL.n253 585
R76 VTAIL.n201 VTAIL.n200 585
R77 VTAIL.n248 VTAIL.n247 585
R78 VTAIL.n246 VTAIL.n245 585
R79 VTAIL.n205 VTAIL.n204 585
R80 VTAIL.n240 VTAIL.n239 585
R81 VTAIL.n238 VTAIL.n237 585
R82 VTAIL.n209 VTAIL.n208 585
R83 VTAIL.n232 VTAIL.n231 585
R84 VTAIL.n230 VTAIL.n229 585
R85 VTAIL.n213 VTAIL.n212 585
R86 VTAIL.n224 VTAIL.n223 585
R87 VTAIL.n222 VTAIL.n221 585
R88 VTAIL.n217 VTAIL.n216 585
R89 VTAIL.n181 VTAIL.n180 585
R90 VTAIL.n179 VTAIL.n178 585
R91 VTAIL.n100 VTAIL.n99 585
R92 VTAIL.n173 VTAIL.n172 585
R93 VTAIL.n171 VTAIL.n102 585
R94 VTAIL.n170 VTAIL.n169 585
R95 VTAIL.n105 VTAIL.n103 585
R96 VTAIL.n164 VTAIL.n163 585
R97 VTAIL.n162 VTAIL.n161 585
R98 VTAIL.n109 VTAIL.n108 585
R99 VTAIL.n156 VTAIL.n155 585
R100 VTAIL.n154 VTAIL.n153 585
R101 VTAIL.n113 VTAIL.n112 585
R102 VTAIL.n148 VTAIL.n147 585
R103 VTAIL.n146 VTAIL.n145 585
R104 VTAIL.n117 VTAIL.n116 585
R105 VTAIL.n140 VTAIL.n139 585
R106 VTAIL.n138 VTAIL.n137 585
R107 VTAIL.n121 VTAIL.n120 585
R108 VTAIL.n132 VTAIL.n131 585
R109 VTAIL.n130 VTAIL.n129 585
R110 VTAIL.n125 VTAIL.n124 585
R111 VTAIL.n307 VTAIL.t0 327.466
R112 VTAIL.n31 VTAIL.t8 327.466
R113 VTAIL.n218 VTAIL.t6 327.466
R114 VTAIL.n126 VTAIL.t4 327.466
R115 VTAIL.n311 VTAIL.n305 171.744
R116 VTAIL.n312 VTAIL.n311 171.744
R117 VTAIL.n312 VTAIL.n301 171.744
R118 VTAIL.n319 VTAIL.n301 171.744
R119 VTAIL.n320 VTAIL.n319 171.744
R120 VTAIL.n320 VTAIL.n297 171.744
R121 VTAIL.n327 VTAIL.n297 171.744
R122 VTAIL.n328 VTAIL.n327 171.744
R123 VTAIL.n328 VTAIL.n293 171.744
R124 VTAIL.n335 VTAIL.n293 171.744
R125 VTAIL.n336 VTAIL.n335 171.744
R126 VTAIL.n336 VTAIL.n289 171.744
R127 VTAIL.n343 VTAIL.n289 171.744
R128 VTAIL.n344 VTAIL.n343 171.744
R129 VTAIL.n344 VTAIL.n285 171.744
R130 VTAIL.n352 VTAIL.n285 171.744
R131 VTAIL.n353 VTAIL.n352 171.744
R132 VTAIL.n354 VTAIL.n353 171.744
R133 VTAIL.n354 VTAIL.n281 171.744
R134 VTAIL.n361 VTAIL.n281 171.744
R135 VTAIL.n362 VTAIL.n361 171.744
R136 VTAIL.n35 VTAIL.n29 171.744
R137 VTAIL.n36 VTAIL.n35 171.744
R138 VTAIL.n36 VTAIL.n25 171.744
R139 VTAIL.n43 VTAIL.n25 171.744
R140 VTAIL.n44 VTAIL.n43 171.744
R141 VTAIL.n44 VTAIL.n21 171.744
R142 VTAIL.n51 VTAIL.n21 171.744
R143 VTAIL.n52 VTAIL.n51 171.744
R144 VTAIL.n52 VTAIL.n17 171.744
R145 VTAIL.n59 VTAIL.n17 171.744
R146 VTAIL.n60 VTAIL.n59 171.744
R147 VTAIL.n60 VTAIL.n13 171.744
R148 VTAIL.n67 VTAIL.n13 171.744
R149 VTAIL.n68 VTAIL.n67 171.744
R150 VTAIL.n68 VTAIL.n9 171.744
R151 VTAIL.n76 VTAIL.n9 171.744
R152 VTAIL.n77 VTAIL.n76 171.744
R153 VTAIL.n78 VTAIL.n77 171.744
R154 VTAIL.n78 VTAIL.n5 171.744
R155 VTAIL.n85 VTAIL.n5 171.744
R156 VTAIL.n86 VTAIL.n85 171.744
R157 VTAIL.n272 VTAIL.n271 171.744
R158 VTAIL.n271 VTAIL.n191 171.744
R159 VTAIL.n264 VTAIL.n191 171.744
R160 VTAIL.n264 VTAIL.n263 171.744
R161 VTAIL.n263 VTAIL.n262 171.744
R162 VTAIL.n262 VTAIL.n195 171.744
R163 VTAIL.n255 VTAIL.n195 171.744
R164 VTAIL.n255 VTAIL.n254 171.744
R165 VTAIL.n254 VTAIL.n200 171.744
R166 VTAIL.n247 VTAIL.n200 171.744
R167 VTAIL.n247 VTAIL.n246 171.744
R168 VTAIL.n246 VTAIL.n204 171.744
R169 VTAIL.n239 VTAIL.n204 171.744
R170 VTAIL.n239 VTAIL.n238 171.744
R171 VTAIL.n238 VTAIL.n208 171.744
R172 VTAIL.n231 VTAIL.n208 171.744
R173 VTAIL.n231 VTAIL.n230 171.744
R174 VTAIL.n230 VTAIL.n212 171.744
R175 VTAIL.n223 VTAIL.n212 171.744
R176 VTAIL.n223 VTAIL.n222 171.744
R177 VTAIL.n222 VTAIL.n216 171.744
R178 VTAIL.n180 VTAIL.n179 171.744
R179 VTAIL.n179 VTAIL.n99 171.744
R180 VTAIL.n172 VTAIL.n99 171.744
R181 VTAIL.n172 VTAIL.n171 171.744
R182 VTAIL.n171 VTAIL.n170 171.744
R183 VTAIL.n170 VTAIL.n103 171.744
R184 VTAIL.n163 VTAIL.n103 171.744
R185 VTAIL.n163 VTAIL.n162 171.744
R186 VTAIL.n162 VTAIL.n108 171.744
R187 VTAIL.n155 VTAIL.n108 171.744
R188 VTAIL.n155 VTAIL.n154 171.744
R189 VTAIL.n154 VTAIL.n112 171.744
R190 VTAIL.n147 VTAIL.n112 171.744
R191 VTAIL.n147 VTAIL.n146 171.744
R192 VTAIL.n146 VTAIL.n116 171.744
R193 VTAIL.n139 VTAIL.n116 171.744
R194 VTAIL.n139 VTAIL.n138 171.744
R195 VTAIL.n138 VTAIL.n120 171.744
R196 VTAIL.n131 VTAIL.n120 171.744
R197 VTAIL.n131 VTAIL.n130 171.744
R198 VTAIL.n130 VTAIL.n124 171.744
R199 VTAIL.t0 VTAIL.n305 85.8723
R200 VTAIL.t8 VTAIL.n29 85.8723
R201 VTAIL.t6 VTAIL.n216 85.8723
R202 VTAIL.t4 VTAIL.n124 85.8723
R203 VTAIL.n187 VTAIL.n186 52.7355
R204 VTAIL.n95 VTAIL.n94 52.7355
R205 VTAIL.n1 VTAIL.n0 52.7353
R206 VTAIL.n93 VTAIL.n92 52.7353
R207 VTAIL.n367 VTAIL.n366 31.7975
R208 VTAIL.n91 VTAIL.n90 31.7975
R209 VTAIL.n277 VTAIL.n276 31.7975
R210 VTAIL.n185 VTAIL.n184 31.7975
R211 VTAIL.n95 VTAIL.n93 27.7462
R212 VTAIL.n367 VTAIL.n277 26.9789
R213 VTAIL.n307 VTAIL.n306 16.3895
R214 VTAIL.n31 VTAIL.n30 16.3895
R215 VTAIL.n218 VTAIL.n217 16.3895
R216 VTAIL.n126 VTAIL.n125 16.3895
R217 VTAIL.n355 VTAIL.n284 13.1884
R218 VTAIL.n79 VTAIL.n8 13.1884
R219 VTAIL.n265 VTAIL.n194 13.1884
R220 VTAIL.n173 VTAIL.n102 13.1884
R221 VTAIL.n310 VTAIL.n309 12.8005
R222 VTAIL.n351 VTAIL.n350 12.8005
R223 VTAIL.n356 VTAIL.n282 12.8005
R224 VTAIL.n34 VTAIL.n33 12.8005
R225 VTAIL.n75 VTAIL.n74 12.8005
R226 VTAIL.n80 VTAIL.n6 12.8005
R227 VTAIL.n266 VTAIL.n192 12.8005
R228 VTAIL.n261 VTAIL.n196 12.8005
R229 VTAIL.n221 VTAIL.n220 12.8005
R230 VTAIL.n174 VTAIL.n100 12.8005
R231 VTAIL.n169 VTAIL.n104 12.8005
R232 VTAIL.n129 VTAIL.n128 12.8005
R233 VTAIL.n313 VTAIL.n304 12.0247
R234 VTAIL.n349 VTAIL.n286 12.0247
R235 VTAIL.n360 VTAIL.n359 12.0247
R236 VTAIL.n37 VTAIL.n28 12.0247
R237 VTAIL.n73 VTAIL.n10 12.0247
R238 VTAIL.n84 VTAIL.n83 12.0247
R239 VTAIL.n270 VTAIL.n269 12.0247
R240 VTAIL.n260 VTAIL.n197 12.0247
R241 VTAIL.n224 VTAIL.n215 12.0247
R242 VTAIL.n178 VTAIL.n177 12.0247
R243 VTAIL.n168 VTAIL.n105 12.0247
R244 VTAIL.n132 VTAIL.n123 12.0247
R245 VTAIL.n314 VTAIL.n302 11.249
R246 VTAIL.n346 VTAIL.n345 11.249
R247 VTAIL.n363 VTAIL.n280 11.249
R248 VTAIL.n38 VTAIL.n26 11.249
R249 VTAIL.n70 VTAIL.n69 11.249
R250 VTAIL.n87 VTAIL.n4 11.249
R251 VTAIL.n273 VTAIL.n190 11.249
R252 VTAIL.n257 VTAIL.n256 11.249
R253 VTAIL.n225 VTAIL.n213 11.249
R254 VTAIL.n181 VTAIL.n98 11.249
R255 VTAIL.n165 VTAIL.n164 11.249
R256 VTAIL.n133 VTAIL.n121 11.249
R257 VTAIL.n318 VTAIL.n317 10.4732
R258 VTAIL.n342 VTAIL.n288 10.4732
R259 VTAIL.n364 VTAIL.n278 10.4732
R260 VTAIL.n42 VTAIL.n41 10.4732
R261 VTAIL.n66 VTAIL.n12 10.4732
R262 VTAIL.n88 VTAIL.n2 10.4732
R263 VTAIL.n274 VTAIL.n188 10.4732
R264 VTAIL.n253 VTAIL.n199 10.4732
R265 VTAIL.n229 VTAIL.n228 10.4732
R266 VTAIL.n182 VTAIL.n96 10.4732
R267 VTAIL.n161 VTAIL.n107 10.4732
R268 VTAIL.n137 VTAIL.n136 10.4732
R269 VTAIL.n321 VTAIL.n300 9.69747
R270 VTAIL.n341 VTAIL.n290 9.69747
R271 VTAIL.n45 VTAIL.n24 9.69747
R272 VTAIL.n65 VTAIL.n14 9.69747
R273 VTAIL.n252 VTAIL.n201 9.69747
R274 VTAIL.n232 VTAIL.n211 9.69747
R275 VTAIL.n160 VTAIL.n109 9.69747
R276 VTAIL.n140 VTAIL.n119 9.69747
R277 VTAIL.n366 VTAIL.n365 9.45567
R278 VTAIL.n90 VTAIL.n89 9.45567
R279 VTAIL.n276 VTAIL.n275 9.45567
R280 VTAIL.n184 VTAIL.n183 9.45567
R281 VTAIL.n365 VTAIL.n364 9.3005
R282 VTAIL.n280 VTAIL.n279 9.3005
R283 VTAIL.n359 VTAIL.n358 9.3005
R284 VTAIL.n357 VTAIL.n356 9.3005
R285 VTAIL.n296 VTAIL.n295 9.3005
R286 VTAIL.n325 VTAIL.n324 9.3005
R287 VTAIL.n323 VTAIL.n322 9.3005
R288 VTAIL.n300 VTAIL.n299 9.3005
R289 VTAIL.n317 VTAIL.n316 9.3005
R290 VTAIL.n315 VTAIL.n314 9.3005
R291 VTAIL.n304 VTAIL.n303 9.3005
R292 VTAIL.n309 VTAIL.n308 9.3005
R293 VTAIL.n331 VTAIL.n330 9.3005
R294 VTAIL.n333 VTAIL.n332 9.3005
R295 VTAIL.n292 VTAIL.n291 9.3005
R296 VTAIL.n339 VTAIL.n338 9.3005
R297 VTAIL.n341 VTAIL.n340 9.3005
R298 VTAIL.n288 VTAIL.n287 9.3005
R299 VTAIL.n347 VTAIL.n346 9.3005
R300 VTAIL.n349 VTAIL.n348 9.3005
R301 VTAIL.n350 VTAIL.n283 9.3005
R302 VTAIL.n89 VTAIL.n88 9.3005
R303 VTAIL.n4 VTAIL.n3 9.3005
R304 VTAIL.n83 VTAIL.n82 9.3005
R305 VTAIL.n81 VTAIL.n80 9.3005
R306 VTAIL.n20 VTAIL.n19 9.3005
R307 VTAIL.n49 VTAIL.n48 9.3005
R308 VTAIL.n47 VTAIL.n46 9.3005
R309 VTAIL.n24 VTAIL.n23 9.3005
R310 VTAIL.n41 VTAIL.n40 9.3005
R311 VTAIL.n39 VTAIL.n38 9.3005
R312 VTAIL.n28 VTAIL.n27 9.3005
R313 VTAIL.n33 VTAIL.n32 9.3005
R314 VTAIL.n55 VTAIL.n54 9.3005
R315 VTAIL.n57 VTAIL.n56 9.3005
R316 VTAIL.n16 VTAIL.n15 9.3005
R317 VTAIL.n63 VTAIL.n62 9.3005
R318 VTAIL.n65 VTAIL.n64 9.3005
R319 VTAIL.n12 VTAIL.n11 9.3005
R320 VTAIL.n71 VTAIL.n70 9.3005
R321 VTAIL.n73 VTAIL.n72 9.3005
R322 VTAIL.n74 VTAIL.n7 9.3005
R323 VTAIL.n244 VTAIL.n243 9.3005
R324 VTAIL.n203 VTAIL.n202 9.3005
R325 VTAIL.n250 VTAIL.n249 9.3005
R326 VTAIL.n252 VTAIL.n251 9.3005
R327 VTAIL.n199 VTAIL.n198 9.3005
R328 VTAIL.n258 VTAIL.n257 9.3005
R329 VTAIL.n260 VTAIL.n259 9.3005
R330 VTAIL.n196 VTAIL.n193 9.3005
R331 VTAIL.n275 VTAIL.n274 9.3005
R332 VTAIL.n190 VTAIL.n189 9.3005
R333 VTAIL.n269 VTAIL.n268 9.3005
R334 VTAIL.n267 VTAIL.n266 9.3005
R335 VTAIL.n242 VTAIL.n241 9.3005
R336 VTAIL.n207 VTAIL.n206 9.3005
R337 VTAIL.n236 VTAIL.n235 9.3005
R338 VTAIL.n234 VTAIL.n233 9.3005
R339 VTAIL.n211 VTAIL.n210 9.3005
R340 VTAIL.n228 VTAIL.n227 9.3005
R341 VTAIL.n226 VTAIL.n225 9.3005
R342 VTAIL.n215 VTAIL.n214 9.3005
R343 VTAIL.n220 VTAIL.n219 9.3005
R344 VTAIL.n152 VTAIL.n151 9.3005
R345 VTAIL.n111 VTAIL.n110 9.3005
R346 VTAIL.n158 VTAIL.n157 9.3005
R347 VTAIL.n160 VTAIL.n159 9.3005
R348 VTAIL.n107 VTAIL.n106 9.3005
R349 VTAIL.n166 VTAIL.n165 9.3005
R350 VTAIL.n168 VTAIL.n167 9.3005
R351 VTAIL.n104 VTAIL.n101 9.3005
R352 VTAIL.n183 VTAIL.n182 9.3005
R353 VTAIL.n98 VTAIL.n97 9.3005
R354 VTAIL.n177 VTAIL.n176 9.3005
R355 VTAIL.n175 VTAIL.n174 9.3005
R356 VTAIL.n150 VTAIL.n149 9.3005
R357 VTAIL.n115 VTAIL.n114 9.3005
R358 VTAIL.n144 VTAIL.n143 9.3005
R359 VTAIL.n142 VTAIL.n141 9.3005
R360 VTAIL.n119 VTAIL.n118 9.3005
R361 VTAIL.n136 VTAIL.n135 9.3005
R362 VTAIL.n134 VTAIL.n133 9.3005
R363 VTAIL.n123 VTAIL.n122 9.3005
R364 VTAIL.n128 VTAIL.n127 9.3005
R365 VTAIL.n322 VTAIL.n298 8.92171
R366 VTAIL.n338 VTAIL.n337 8.92171
R367 VTAIL.n46 VTAIL.n22 8.92171
R368 VTAIL.n62 VTAIL.n61 8.92171
R369 VTAIL.n249 VTAIL.n248 8.92171
R370 VTAIL.n233 VTAIL.n209 8.92171
R371 VTAIL.n157 VTAIL.n156 8.92171
R372 VTAIL.n141 VTAIL.n117 8.92171
R373 VTAIL.n326 VTAIL.n325 8.14595
R374 VTAIL.n334 VTAIL.n292 8.14595
R375 VTAIL.n50 VTAIL.n49 8.14595
R376 VTAIL.n58 VTAIL.n16 8.14595
R377 VTAIL.n245 VTAIL.n203 8.14595
R378 VTAIL.n237 VTAIL.n236 8.14595
R379 VTAIL.n153 VTAIL.n111 8.14595
R380 VTAIL.n145 VTAIL.n144 8.14595
R381 VTAIL.n329 VTAIL.n296 7.3702
R382 VTAIL.n333 VTAIL.n294 7.3702
R383 VTAIL.n53 VTAIL.n20 7.3702
R384 VTAIL.n57 VTAIL.n18 7.3702
R385 VTAIL.n244 VTAIL.n205 7.3702
R386 VTAIL.n240 VTAIL.n207 7.3702
R387 VTAIL.n152 VTAIL.n113 7.3702
R388 VTAIL.n148 VTAIL.n115 7.3702
R389 VTAIL.n330 VTAIL.n329 6.59444
R390 VTAIL.n330 VTAIL.n294 6.59444
R391 VTAIL.n54 VTAIL.n53 6.59444
R392 VTAIL.n54 VTAIL.n18 6.59444
R393 VTAIL.n241 VTAIL.n205 6.59444
R394 VTAIL.n241 VTAIL.n240 6.59444
R395 VTAIL.n149 VTAIL.n113 6.59444
R396 VTAIL.n149 VTAIL.n148 6.59444
R397 VTAIL.n326 VTAIL.n296 5.81868
R398 VTAIL.n334 VTAIL.n333 5.81868
R399 VTAIL.n50 VTAIL.n20 5.81868
R400 VTAIL.n58 VTAIL.n57 5.81868
R401 VTAIL.n245 VTAIL.n244 5.81868
R402 VTAIL.n237 VTAIL.n207 5.81868
R403 VTAIL.n153 VTAIL.n152 5.81868
R404 VTAIL.n145 VTAIL.n115 5.81868
R405 VTAIL.n325 VTAIL.n298 5.04292
R406 VTAIL.n337 VTAIL.n292 5.04292
R407 VTAIL.n49 VTAIL.n22 5.04292
R408 VTAIL.n61 VTAIL.n16 5.04292
R409 VTAIL.n248 VTAIL.n203 5.04292
R410 VTAIL.n236 VTAIL.n209 5.04292
R411 VTAIL.n156 VTAIL.n111 5.04292
R412 VTAIL.n144 VTAIL.n117 5.04292
R413 VTAIL.n322 VTAIL.n321 4.26717
R414 VTAIL.n338 VTAIL.n290 4.26717
R415 VTAIL.n46 VTAIL.n45 4.26717
R416 VTAIL.n62 VTAIL.n14 4.26717
R417 VTAIL.n249 VTAIL.n201 4.26717
R418 VTAIL.n233 VTAIL.n232 4.26717
R419 VTAIL.n157 VTAIL.n109 4.26717
R420 VTAIL.n141 VTAIL.n140 4.26717
R421 VTAIL.n308 VTAIL.n307 3.70982
R422 VTAIL.n32 VTAIL.n31 3.70982
R423 VTAIL.n219 VTAIL.n218 3.70982
R424 VTAIL.n127 VTAIL.n126 3.70982
R425 VTAIL.n318 VTAIL.n300 3.49141
R426 VTAIL.n342 VTAIL.n341 3.49141
R427 VTAIL.n366 VTAIL.n278 3.49141
R428 VTAIL.n42 VTAIL.n24 3.49141
R429 VTAIL.n66 VTAIL.n65 3.49141
R430 VTAIL.n90 VTAIL.n2 3.49141
R431 VTAIL.n276 VTAIL.n188 3.49141
R432 VTAIL.n253 VTAIL.n252 3.49141
R433 VTAIL.n229 VTAIL.n211 3.49141
R434 VTAIL.n184 VTAIL.n96 3.49141
R435 VTAIL.n161 VTAIL.n160 3.49141
R436 VTAIL.n137 VTAIL.n119 3.49141
R437 VTAIL.n317 VTAIL.n302 2.71565
R438 VTAIL.n345 VTAIL.n288 2.71565
R439 VTAIL.n364 VTAIL.n363 2.71565
R440 VTAIL.n41 VTAIL.n26 2.71565
R441 VTAIL.n69 VTAIL.n12 2.71565
R442 VTAIL.n88 VTAIL.n87 2.71565
R443 VTAIL.n274 VTAIL.n273 2.71565
R444 VTAIL.n256 VTAIL.n199 2.71565
R445 VTAIL.n228 VTAIL.n213 2.71565
R446 VTAIL.n182 VTAIL.n181 2.71565
R447 VTAIL.n164 VTAIL.n107 2.71565
R448 VTAIL.n136 VTAIL.n121 2.71565
R449 VTAIL.n0 VTAIL.t2 2.02447
R450 VTAIL.n0 VTAIL.t5 2.02447
R451 VTAIL.n92 VTAIL.t10 2.02447
R452 VTAIL.n92 VTAIL.t11 2.02447
R453 VTAIL.n186 VTAIL.t9 2.02447
R454 VTAIL.n186 VTAIL.t7 2.02447
R455 VTAIL.n94 VTAIL.t3 2.02447
R456 VTAIL.n94 VTAIL.t1 2.02447
R457 VTAIL.n314 VTAIL.n313 1.93989
R458 VTAIL.n346 VTAIL.n286 1.93989
R459 VTAIL.n360 VTAIL.n280 1.93989
R460 VTAIL.n38 VTAIL.n37 1.93989
R461 VTAIL.n70 VTAIL.n10 1.93989
R462 VTAIL.n84 VTAIL.n4 1.93989
R463 VTAIL.n270 VTAIL.n190 1.93989
R464 VTAIL.n257 VTAIL.n197 1.93989
R465 VTAIL.n225 VTAIL.n224 1.93989
R466 VTAIL.n178 VTAIL.n98 1.93989
R467 VTAIL.n165 VTAIL.n105 1.93989
R468 VTAIL.n133 VTAIL.n132 1.93989
R469 VTAIL.n310 VTAIL.n304 1.16414
R470 VTAIL.n351 VTAIL.n349 1.16414
R471 VTAIL.n359 VTAIL.n282 1.16414
R472 VTAIL.n34 VTAIL.n28 1.16414
R473 VTAIL.n75 VTAIL.n73 1.16414
R474 VTAIL.n83 VTAIL.n6 1.16414
R475 VTAIL.n269 VTAIL.n192 1.16414
R476 VTAIL.n261 VTAIL.n260 1.16414
R477 VTAIL.n221 VTAIL.n215 1.16414
R478 VTAIL.n177 VTAIL.n100 1.16414
R479 VTAIL.n169 VTAIL.n168 1.16414
R480 VTAIL.n129 VTAIL.n123 1.16414
R481 VTAIL.n187 VTAIL.n185 0.853948
R482 VTAIL.n91 VTAIL.n1 0.853948
R483 VTAIL.n185 VTAIL.n95 0.767741
R484 VTAIL.n277 VTAIL.n187 0.767741
R485 VTAIL.n93 VTAIL.n91 0.767741
R486 VTAIL VTAIL.n367 0.517741
R487 VTAIL.n309 VTAIL.n306 0.388379
R488 VTAIL.n350 VTAIL.n284 0.388379
R489 VTAIL.n356 VTAIL.n355 0.388379
R490 VTAIL.n33 VTAIL.n30 0.388379
R491 VTAIL.n74 VTAIL.n8 0.388379
R492 VTAIL.n80 VTAIL.n79 0.388379
R493 VTAIL.n266 VTAIL.n265 0.388379
R494 VTAIL.n196 VTAIL.n194 0.388379
R495 VTAIL.n220 VTAIL.n217 0.388379
R496 VTAIL.n174 VTAIL.n173 0.388379
R497 VTAIL.n104 VTAIL.n102 0.388379
R498 VTAIL.n128 VTAIL.n125 0.388379
R499 VTAIL VTAIL.n1 0.2505
R500 VTAIL.n308 VTAIL.n303 0.155672
R501 VTAIL.n315 VTAIL.n303 0.155672
R502 VTAIL.n316 VTAIL.n315 0.155672
R503 VTAIL.n316 VTAIL.n299 0.155672
R504 VTAIL.n323 VTAIL.n299 0.155672
R505 VTAIL.n324 VTAIL.n323 0.155672
R506 VTAIL.n324 VTAIL.n295 0.155672
R507 VTAIL.n331 VTAIL.n295 0.155672
R508 VTAIL.n332 VTAIL.n331 0.155672
R509 VTAIL.n332 VTAIL.n291 0.155672
R510 VTAIL.n339 VTAIL.n291 0.155672
R511 VTAIL.n340 VTAIL.n339 0.155672
R512 VTAIL.n340 VTAIL.n287 0.155672
R513 VTAIL.n347 VTAIL.n287 0.155672
R514 VTAIL.n348 VTAIL.n347 0.155672
R515 VTAIL.n348 VTAIL.n283 0.155672
R516 VTAIL.n357 VTAIL.n283 0.155672
R517 VTAIL.n358 VTAIL.n357 0.155672
R518 VTAIL.n358 VTAIL.n279 0.155672
R519 VTAIL.n365 VTAIL.n279 0.155672
R520 VTAIL.n32 VTAIL.n27 0.155672
R521 VTAIL.n39 VTAIL.n27 0.155672
R522 VTAIL.n40 VTAIL.n39 0.155672
R523 VTAIL.n40 VTAIL.n23 0.155672
R524 VTAIL.n47 VTAIL.n23 0.155672
R525 VTAIL.n48 VTAIL.n47 0.155672
R526 VTAIL.n48 VTAIL.n19 0.155672
R527 VTAIL.n55 VTAIL.n19 0.155672
R528 VTAIL.n56 VTAIL.n55 0.155672
R529 VTAIL.n56 VTAIL.n15 0.155672
R530 VTAIL.n63 VTAIL.n15 0.155672
R531 VTAIL.n64 VTAIL.n63 0.155672
R532 VTAIL.n64 VTAIL.n11 0.155672
R533 VTAIL.n71 VTAIL.n11 0.155672
R534 VTAIL.n72 VTAIL.n71 0.155672
R535 VTAIL.n72 VTAIL.n7 0.155672
R536 VTAIL.n81 VTAIL.n7 0.155672
R537 VTAIL.n82 VTAIL.n81 0.155672
R538 VTAIL.n82 VTAIL.n3 0.155672
R539 VTAIL.n89 VTAIL.n3 0.155672
R540 VTAIL.n275 VTAIL.n189 0.155672
R541 VTAIL.n268 VTAIL.n189 0.155672
R542 VTAIL.n268 VTAIL.n267 0.155672
R543 VTAIL.n267 VTAIL.n193 0.155672
R544 VTAIL.n259 VTAIL.n193 0.155672
R545 VTAIL.n259 VTAIL.n258 0.155672
R546 VTAIL.n258 VTAIL.n198 0.155672
R547 VTAIL.n251 VTAIL.n198 0.155672
R548 VTAIL.n251 VTAIL.n250 0.155672
R549 VTAIL.n250 VTAIL.n202 0.155672
R550 VTAIL.n243 VTAIL.n202 0.155672
R551 VTAIL.n243 VTAIL.n242 0.155672
R552 VTAIL.n242 VTAIL.n206 0.155672
R553 VTAIL.n235 VTAIL.n206 0.155672
R554 VTAIL.n235 VTAIL.n234 0.155672
R555 VTAIL.n234 VTAIL.n210 0.155672
R556 VTAIL.n227 VTAIL.n210 0.155672
R557 VTAIL.n227 VTAIL.n226 0.155672
R558 VTAIL.n226 VTAIL.n214 0.155672
R559 VTAIL.n219 VTAIL.n214 0.155672
R560 VTAIL.n183 VTAIL.n97 0.155672
R561 VTAIL.n176 VTAIL.n97 0.155672
R562 VTAIL.n176 VTAIL.n175 0.155672
R563 VTAIL.n175 VTAIL.n101 0.155672
R564 VTAIL.n167 VTAIL.n101 0.155672
R565 VTAIL.n167 VTAIL.n166 0.155672
R566 VTAIL.n166 VTAIL.n106 0.155672
R567 VTAIL.n159 VTAIL.n106 0.155672
R568 VTAIL.n159 VTAIL.n158 0.155672
R569 VTAIL.n158 VTAIL.n110 0.155672
R570 VTAIL.n151 VTAIL.n110 0.155672
R571 VTAIL.n151 VTAIL.n150 0.155672
R572 VTAIL.n150 VTAIL.n114 0.155672
R573 VTAIL.n143 VTAIL.n114 0.155672
R574 VTAIL.n143 VTAIL.n142 0.155672
R575 VTAIL.n142 VTAIL.n118 0.155672
R576 VTAIL.n135 VTAIL.n118 0.155672
R577 VTAIL.n135 VTAIL.n134 0.155672
R578 VTAIL.n134 VTAIL.n122 0.155672
R579 VTAIL.n127 VTAIL.n122 0.155672
R580 VDD1.n84 VDD1.n0 756.745
R581 VDD1.n173 VDD1.n89 756.745
R582 VDD1.n85 VDD1.n84 585
R583 VDD1.n83 VDD1.n82 585
R584 VDD1.n4 VDD1.n3 585
R585 VDD1.n77 VDD1.n76 585
R586 VDD1.n75 VDD1.n6 585
R587 VDD1.n74 VDD1.n73 585
R588 VDD1.n9 VDD1.n7 585
R589 VDD1.n68 VDD1.n67 585
R590 VDD1.n66 VDD1.n65 585
R591 VDD1.n13 VDD1.n12 585
R592 VDD1.n60 VDD1.n59 585
R593 VDD1.n58 VDD1.n57 585
R594 VDD1.n17 VDD1.n16 585
R595 VDD1.n52 VDD1.n51 585
R596 VDD1.n50 VDD1.n49 585
R597 VDD1.n21 VDD1.n20 585
R598 VDD1.n44 VDD1.n43 585
R599 VDD1.n42 VDD1.n41 585
R600 VDD1.n25 VDD1.n24 585
R601 VDD1.n36 VDD1.n35 585
R602 VDD1.n34 VDD1.n33 585
R603 VDD1.n29 VDD1.n28 585
R604 VDD1.n117 VDD1.n116 585
R605 VDD1.n122 VDD1.n121 585
R606 VDD1.n124 VDD1.n123 585
R607 VDD1.n113 VDD1.n112 585
R608 VDD1.n130 VDD1.n129 585
R609 VDD1.n132 VDD1.n131 585
R610 VDD1.n109 VDD1.n108 585
R611 VDD1.n138 VDD1.n137 585
R612 VDD1.n140 VDD1.n139 585
R613 VDD1.n105 VDD1.n104 585
R614 VDD1.n146 VDD1.n145 585
R615 VDD1.n148 VDD1.n147 585
R616 VDD1.n101 VDD1.n100 585
R617 VDD1.n154 VDD1.n153 585
R618 VDD1.n156 VDD1.n155 585
R619 VDD1.n97 VDD1.n96 585
R620 VDD1.n163 VDD1.n162 585
R621 VDD1.n164 VDD1.n95 585
R622 VDD1.n166 VDD1.n165 585
R623 VDD1.n93 VDD1.n92 585
R624 VDD1.n172 VDD1.n171 585
R625 VDD1.n174 VDD1.n173 585
R626 VDD1.n30 VDD1.t5 327.466
R627 VDD1.n118 VDD1.t4 327.466
R628 VDD1.n84 VDD1.n83 171.744
R629 VDD1.n83 VDD1.n3 171.744
R630 VDD1.n76 VDD1.n3 171.744
R631 VDD1.n76 VDD1.n75 171.744
R632 VDD1.n75 VDD1.n74 171.744
R633 VDD1.n74 VDD1.n7 171.744
R634 VDD1.n67 VDD1.n7 171.744
R635 VDD1.n67 VDD1.n66 171.744
R636 VDD1.n66 VDD1.n12 171.744
R637 VDD1.n59 VDD1.n12 171.744
R638 VDD1.n59 VDD1.n58 171.744
R639 VDD1.n58 VDD1.n16 171.744
R640 VDD1.n51 VDD1.n16 171.744
R641 VDD1.n51 VDD1.n50 171.744
R642 VDD1.n50 VDD1.n20 171.744
R643 VDD1.n43 VDD1.n20 171.744
R644 VDD1.n43 VDD1.n42 171.744
R645 VDD1.n42 VDD1.n24 171.744
R646 VDD1.n35 VDD1.n24 171.744
R647 VDD1.n35 VDD1.n34 171.744
R648 VDD1.n34 VDD1.n28 171.744
R649 VDD1.n122 VDD1.n116 171.744
R650 VDD1.n123 VDD1.n122 171.744
R651 VDD1.n123 VDD1.n112 171.744
R652 VDD1.n130 VDD1.n112 171.744
R653 VDD1.n131 VDD1.n130 171.744
R654 VDD1.n131 VDD1.n108 171.744
R655 VDD1.n138 VDD1.n108 171.744
R656 VDD1.n139 VDD1.n138 171.744
R657 VDD1.n139 VDD1.n104 171.744
R658 VDD1.n146 VDD1.n104 171.744
R659 VDD1.n147 VDD1.n146 171.744
R660 VDD1.n147 VDD1.n100 171.744
R661 VDD1.n154 VDD1.n100 171.744
R662 VDD1.n155 VDD1.n154 171.744
R663 VDD1.n155 VDD1.n96 171.744
R664 VDD1.n163 VDD1.n96 171.744
R665 VDD1.n164 VDD1.n163 171.744
R666 VDD1.n165 VDD1.n164 171.744
R667 VDD1.n165 VDD1.n92 171.744
R668 VDD1.n172 VDD1.n92 171.744
R669 VDD1.n173 VDD1.n172 171.744
R670 VDD1.t5 VDD1.n28 85.8723
R671 VDD1.t4 VDD1.n116 85.8723
R672 VDD1.n179 VDD1.n178 69.5505
R673 VDD1.n181 VDD1.n180 69.4141
R674 VDD1 VDD1.n88 49.1099
R675 VDD1.n179 VDD1.n177 48.9963
R676 VDD1.n181 VDD1.n179 41.0203
R677 VDD1.n30 VDD1.n29 16.3895
R678 VDD1.n118 VDD1.n117 16.3895
R679 VDD1.n77 VDD1.n6 13.1884
R680 VDD1.n166 VDD1.n95 13.1884
R681 VDD1.n78 VDD1.n4 12.8005
R682 VDD1.n73 VDD1.n8 12.8005
R683 VDD1.n33 VDD1.n32 12.8005
R684 VDD1.n121 VDD1.n120 12.8005
R685 VDD1.n162 VDD1.n161 12.8005
R686 VDD1.n167 VDD1.n93 12.8005
R687 VDD1.n82 VDD1.n81 12.0247
R688 VDD1.n72 VDD1.n9 12.0247
R689 VDD1.n36 VDD1.n27 12.0247
R690 VDD1.n124 VDD1.n115 12.0247
R691 VDD1.n160 VDD1.n97 12.0247
R692 VDD1.n171 VDD1.n170 12.0247
R693 VDD1.n85 VDD1.n2 11.249
R694 VDD1.n69 VDD1.n68 11.249
R695 VDD1.n37 VDD1.n25 11.249
R696 VDD1.n125 VDD1.n113 11.249
R697 VDD1.n157 VDD1.n156 11.249
R698 VDD1.n174 VDD1.n91 11.249
R699 VDD1.n86 VDD1.n0 10.4732
R700 VDD1.n65 VDD1.n11 10.4732
R701 VDD1.n41 VDD1.n40 10.4732
R702 VDD1.n129 VDD1.n128 10.4732
R703 VDD1.n153 VDD1.n99 10.4732
R704 VDD1.n175 VDD1.n89 10.4732
R705 VDD1.n64 VDD1.n13 9.69747
R706 VDD1.n44 VDD1.n23 9.69747
R707 VDD1.n132 VDD1.n111 9.69747
R708 VDD1.n152 VDD1.n101 9.69747
R709 VDD1.n88 VDD1.n87 9.45567
R710 VDD1.n177 VDD1.n176 9.45567
R711 VDD1.n56 VDD1.n55 9.3005
R712 VDD1.n15 VDD1.n14 9.3005
R713 VDD1.n62 VDD1.n61 9.3005
R714 VDD1.n64 VDD1.n63 9.3005
R715 VDD1.n11 VDD1.n10 9.3005
R716 VDD1.n70 VDD1.n69 9.3005
R717 VDD1.n72 VDD1.n71 9.3005
R718 VDD1.n8 VDD1.n5 9.3005
R719 VDD1.n87 VDD1.n86 9.3005
R720 VDD1.n2 VDD1.n1 9.3005
R721 VDD1.n81 VDD1.n80 9.3005
R722 VDD1.n79 VDD1.n78 9.3005
R723 VDD1.n54 VDD1.n53 9.3005
R724 VDD1.n19 VDD1.n18 9.3005
R725 VDD1.n48 VDD1.n47 9.3005
R726 VDD1.n46 VDD1.n45 9.3005
R727 VDD1.n23 VDD1.n22 9.3005
R728 VDD1.n40 VDD1.n39 9.3005
R729 VDD1.n38 VDD1.n37 9.3005
R730 VDD1.n27 VDD1.n26 9.3005
R731 VDD1.n32 VDD1.n31 9.3005
R732 VDD1.n176 VDD1.n175 9.3005
R733 VDD1.n91 VDD1.n90 9.3005
R734 VDD1.n170 VDD1.n169 9.3005
R735 VDD1.n168 VDD1.n167 9.3005
R736 VDD1.n107 VDD1.n106 9.3005
R737 VDD1.n136 VDD1.n135 9.3005
R738 VDD1.n134 VDD1.n133 9.3005
R739 VDD1.n111 VDD1.n110 9.3005
R740 VDD1.n128 VDD1.n127 9.3005
R741 VDD1.n126 VDD1.n125 9.3005
R742 VDD1.n115 VDD1.n114 9.3005
R743 VDD1.n120 VDD1.n119 9.3005
R744 VDD1.n142 VDD1.n141 9.3005
R745 VDD1.n144 VDD1.n143 9.3005
R746 VDD1.n103 VDD1.n102 9.3005
R747 VDD1.n150 VDD1.n149 9.3005
R748 VDD1.n152 VDD1.n151 9.3005
R749 VDD1.n99 VDD1.n98 9.3005
R750 VDD1.n158 VDD1.n157 9.3005
R751 VDD1.n160 VDD1.n159 9.3005
R752 VDD1.n161 VDD1.n94 9.3005
R753 VDD1.n61 VDD1.n60 8.92171
R754 VDD1.n45 VDD1.n21 8.92171
R755 VDD1.n133 VDD1.n109 8.92171
R756 VDD1.n149 VDD1.n148 8.92171
R757 VDD1.n57 VDD1.n15 8.14595
R758 VDD1.n49 VDD1.n48 8.14595
R759 VDD1.n137 VDD1.n136 8.14595
R760 VDD1.n145 VDD1.n103 8.14595
R761 VDD1.n56 VDD1.n17 7.3702
R762 VDD1.n52 VDD1.n19 7.3702
R763 VDD1.n140 VDD1.n107 7.3702
R764 VDD1.n144 VDD1.n105 7.3702
R765 VDD1.n53 VDD1.n17 6.59444
R766 VDD1.n53 VDD1.n52 6.59444
R767 VDD1.n141 VDD1.n140 6.59444
R768 VDD1.n141 VDD1.n105 6.59444
R769 VDD1.n57 VDD1.n56 5.81868
R770 VDD1.n49 VDD1.n19 5.81868
R771 VDD1.n137 VDD1.n107 5.81868
R772 VDD1.n145 VDD1.n144 5.81868
R773 VDD1.n60 VDD1.n15 5.04292
R774 VDD1.n48 VDD1.n21 5.04292
R775 VDD1.n136 VDD1.n109 5.04292
R776 VDD1.n148 VDD1.n103 5.04292
R777 VDD1.n61 VDD1.n13 4.26717
R778 VDD1.n45 VDD1.n44 4.26717
R779 VDD1.n133 VDD1.n132 4.26717
R780 VDD1.n149 VDD1.n101 4.26717
R781 VDD1.n31 VDD1.n30 3.70982
R782 VDD1.n119 VDD1.n118 3.70982
R783 VDD1.n88 VDD1.n0 3.49141
R784 VDD1.n65 VDD1.n64 3.49141
R785 VDD1.n41 VDD1.n23 3.49141
R786 VDD1.n129 VDD1.n111 3.49141
R787 VDD1.n153 VDD1.n152 3.49141
R788 VDD1.n177 VDD1.n89 3.49141
R789 VDD1.n86 VDD1.n85 2.71565
R790 VDD1.n68 VDD1.n11 2.71565
R791 VDD1.n40 VDD1.n25 2.71565
R792 VDD1.n128 VDD1.n113 2.71565
R793 VDD1.n156 VDD1.n99 2.71565
R794 VDD1.n175 VDD1.n174 2.71565
R795 VDD1.n180 VDD1.t0 2.02447
R796 VDD1.n180 VDD1.t3 2.02447
R797 VDD1.n178 VDD1.t2 2.02447
R798 VDD1.n178 VDD1.t1 2.02447
R799 VDD1.n82 VDD1.n2 1.93989
R800 VDD1.n69 VDD1.n9 1.93989
R801 VDD1.n37 VDD1.n36 1.93989
R802 VDD1.n125 VDD1.n124 1.93989
R803 VDD1.n157 VDD1.n97 1.93989
R804 VDD1.n171 VDD1.n91 1.93989
R805 VDD1.n81 VDD1.n4 1.16414
R806 VDD1.n73 VDD1.n72 1.16414
R807 VDD1.n33 VDD1.n27 1.16414
R808 VDD1.n121 VDD1.n115 1.16414
R809 VDD1.n162 VDD1.n160 1.16414
R810 VDD1.n170 VDD1.n93 1.16414
R811 VDD1.n78 VDD1.n77 0.388379
R812 VDD1.n8 VDD1.n6 0.388379
R813 VDD1.n32 VDD1.n29 0.388379
R814 VDD1.n120 VDD1.n117 0.388379
R815 VDD1.n161 VDD1.n95 0.388379
R816 VDD1.n167 VDD1.n166 0.388379
R817 VDD1.n87 VDD1.n1 0.155672
R818 VDD1.n80 VDD1.n1 0.155672
R819 VDD1.n80 VDD1.n79 0.155672
R820 VDD1.n79 VDD1.n5 0.155672
R821 VDD1.n71 VDD1.n5 0.155672
R822 VDD1.n71 VDD1.n70 0.155672
R823 VDD1.n70 VDD1.n10 0.155672
R824 VDD1.n63 VDD1.n10 0.155672
R825 VDD1.n63 VDD1.n62 0.155672
R826 VDD1.n62 VDD1.n14 0.155672
R827 VDD1.n55 VDD1.n14 0.155672
R828 VDD1.n55 VDD1.n54 0.155672
R829 VDD1.n54 VDD1.n18 0.155672
R830 VDD1.n47 VDD1.n18 0.155672
R831 VDD1.n47 VDD1.n46 0.155672
R832 VDD1.n46 VDD1.n22 0.155672
R833 VDD1.n39 VDD1.n22 0.155672
R834 VDD1.n39 VDD1.n38 0.155672
R835 VDD1.n38 VDD1.n26 0.155672
R836 VDD1.n31 VDD1.n26 0.155672
R837 VDD1.n119 VDD1.n114 0.155672
R838 VDD1.n126 VDD1.n114 0.155672
R839 VDD1.n127 VDD1.n126 0.155672
R840 VDD1.n127 VDD1.n110 0.155672
R841 VDD1.n134 VDD1.n110 0.155672
R842 VDD1.n135 VDD1.n134 0.155672
R843 VDD1.n135 VDD1.n106 0.155672
R844 VDD1.n142 VDD1.n106 0.155672
R845 VDD1.n143 VDD1.n142 0.155672
R846 VDD1.n143 VDD1.n102 0.155672
R847 VDD1.n150 VDD1.n102 0.155672
R848 VDD1.n151 VDD1.n150 0.155672
R849 VDD1.n151 VDD1.n98 0.155672
R850 VDD1.n158 VDD1.n98 0.155672
R851 VDD1.n159 VDD1.n158 0.155672
R852 VDD1.n159 VDD1.n94 0.155672
R853 VDD1.n168 VDD1.n94 0.155672
R854 VDD1.n169 VDD1.n168 0.155672
R855 VDD1.n169 VDD1.n90 0.155672
R856 VDD1.n176 VDD1.n90 0.155672
R857 VDD1 VDD1.n181 0.134121
R858 B.n128 B.t9 896.27
R859 B.n120 B.t3 896.27
R860 B.n46 B.t0 896.27
R861 B.n38 B.t6 896.27
R862 B.n366 B.n93 585
R863 B.n365 B.n364 585
R864 B.n363 B.n94 585
R865 B.n362 B.n361 585
R866 B.n360 B.n95 585
R867 B.n359 B.n358 585
R868 B.n357 B.n96 585
R869 B.n356 B.n355 585
R870 B.n354 B.n97 585
R871 B.n353 B.n352 585
R872 B.n351 B.n98 585
R873 B.n350 B.n349 585
R874 B.n348 B.n99 585
R875 B.n347 B.n346 585
R876 B.n345 B.n100 585
R877 B.n344 B.n343 585
R878 B.n342 B.n101 585
R879 B.n341 B.n340 585
R880 B.n339 B.n102 585
R881 B.n338 B.n337 585
R882 B.n336 B.n103 585
R883 B.n335 B.n334 585
R884 B.n333 B.n104 585
R885 B.n332 B.n331 585
R886 B.n330 B.n105 585
R887 B.n329 B.n328 585
R888 B.n327 B.n106 585
R889 B.n326 B.n325 585
R890 B.n324 B.n107 585
R891 B.n323 B.n322 585
R892 B.n321 B.n108 585
R893 B.n320 B.n319 585
R894 B.n318 B.n109 585
R895 B.n317 B.n316 585
R896 B.n315 B.n110 585
R897 B.n314 B.n313 585
R898 B.n312 B.n111 585
R899 B.n311 B.n310 585
R900 B.n309 B.n112 585
R901 B.n308 B.n307 585
R902 B.n306 B.n113 585
R903 B.n305 B.n304 585
R904 B.n303 B.n114 585
R905 B.n302 B.n301 585
R906 B.n300 B.n115 585
R907 B.n299 B.n298 585
R908 B.n297 B.n116 585
R909 B.n296 B.n295 585
R910 B.n294 B.n117 585
R911 B.n293 B.n292 585
R912 B.n291 B.n118 585
R913 B.n290 B.n289 585
R914 B.n288 B.n119 585
R915 B.n287 B.n286 585
R916 B.n285 B.n284 585
R917 B.n283 B.n123 585
R918 B.n282 B.n281 585
R919 B.n280 B.n124 585
R920 B.n279 B.n278 585
R921 B.n277 B.n125 585
R922 B.n276 B.n275 585
R923 B.n274 B.n126 585
R924 B.n273 B.n272 585
R925 B.n270 B.n127 585
R926 B.n269 B.n268 585
R927 B.n267 B.n130 585
R928 B.n266 B.n265 585
R929 B.n264 B.n131 585
R930 B.n263 B.n262 585
R931 B.n261 B.n132 585
R932 B.n260 B.n259 585
R933 B.n258 B.n133 585
R934 B.n257 B.n256 585
R935 B.n255 B.n134 585
R936 B.n254 B.n253 585
R937 B.n252 B.n135 585
R938 B.n251 B.n250 585
R939 B.n249 B.n136 585
R940 B.n248 B.n247 585
R941 B.n246 B.n137 585
R942 B.n245 B.n244 585
R943 B.n243 B.n138 585
R944 B.n242 B.n241 585
R945 B.n240 B.n139 585
R946 B.n239 B.n238 585
R947 B.n237 B.n140 585
R948 B.n236 B.n235 585
R949 B.n234 B.n141 585
R950 B.n233 B.n232 585
R951 B.n231 B.n142 585
R952 B.n230 B.n229 585
R953 B.n228 B.n143 585
R954 B.n227 B.n226 585
R955 B.n225 B.n144 585
R956 B.n224 B.n223 585
R957 B.n222 B.n145 585
R958 B.n221 B.n220 585
R959 B.n219 B.n146 585
R960 B.n218 B.n217 585
R961 B.n216 B.n147 585
R962 B.n215 B.n214 585
R963 B.n213 B.n148 585
R964 B.n212 B.n211 585
R965 B.n210 B.n149 585
R966 B.n209 B.n208 585
R967 B.n207 B.n150 585
R968 B.n206 B.n205 585
R969 B.n204 B.n151 585
R970 B.n203 B.n202 585
R971 B.n201 B.n152 585
R972 B.n200 B.n199 585
R973 B.n198 B.n153 585
R974 B.n197 B.n196 585
R975 B.n195 B.n154 585
R976 B.n194 B.n193 585
R977 B.n192 B.n155 585
R978 B.n191 B.n190 585
R979 B.n368 B.n367 585
R980 B.n369 B.n92 585
R981 B.n371 B.n370 585
R982 B.n372 B.n91 585
R983 B.n374 B.n373 585
R984 B.n375 B.n90 585
R985 B.n377 B.n376 585
R986 B.n378 B.n89 585
R987 B.n380 B.n379 585
R988 B.n381 B.n88 585
R989 B.n383 B.n382 585
R990 B.n384 B.n87 585
R991 B.n386 B.n385 585
R992 B.n387 B.n86 585
R993 B.n389 B.n388 585
R994 B.n390 B.n85 585
R995 B.n392 B.n391 585
R996 B.n393 B.n84 585
R997 B.n395 B.n394 585
R998 B.n396 B.n83 585
R999 B.n398 B.n397 585
R1000 B.n399 B.n82 585
R1001 B.n401 B.n400 585
R1002 B.n402 B.n81 585
R1003 B.n404 B.n403 585
R1004 B.n405 B.n80 585
R1005 B.n407 B.n406 585
R1006 B.n408 B.n79 585
R1007 B.n410 B.n409 585
R1008 B.n411 B.n78 585
R1009 B.n413 B.n412 585
R1010 B.n414 B.n77 585
R1011 B.n416 B.n415 585
R1012 B.n417 B.n76 585
R1013 B.n419 B.n418 585
R1014 B.n420 B.n75 585
R1015 B.n422 B.n421 585
R1016 B.n423 B.n74 585
R1017 B.n600 B.n11 585
R1018 B.n599 B.n598 585
R1019 B.n597 B.n12 585
R1020 B.n596 B.n595 585
R1021 B.n594 B.n13 585
R1022 B.n593 B.n592 585
R1023 B.n591 B.n14 585
R1024 B.n590 B.n589 585
R1025 B.n588 B.n15 585
R1026 B.n587 B.n586 585
R1027 B.n585 B.n16 585
R1028 B.n584 B.n583 585
R1029 B.n582 B.n17 585
R1030 B.n581 B.n580 585
R1031 B.n579 B.n18 585
R1032 B.n578 B.n577 585
R1033 B.n576 B.n19 585
R1034 B.n575 B.n574 585
R1035 B.n573 B.n20 585
R1036 B.n572 B.n571 585
R1037 B.n570 B.n21 585
R1038 B.n569 B.n568 585
R1039 B.n567 B.n22 585
R1040 B.n566 B.n565 585
R1041 B.n564 B.n23 585
R1042 B.n563 B.n562 585
R1043 B.n561 B.n24 585
R1044 B.n560 B.n559 585
R1045 B.n558 B.n25 585
R1046 B.n557 B.n556 585
R1047 B.n555 B.n26 585
R1048 B.n554 B.n553 585
R1049 B.n552 B.n27 585
R1050 B.n551 B.n550 585
R1051 B.n549 B.n28 585
R1052 B.n548 B.n547 585
R1053 B.n546 B.n29 585
R1054 B.n545 B.n544 585
R1055 B.n543 B.n30 585
R1056 B.n542 B.n541 585
R1057 B.n540 B.n31 585
R1058 B.n539 B.n538 585
R1059 B.n537 B.n32 585
R1060 B.n536 B.n535 585
R1061 B.n534 B.n33 585
R1062 B.n533 B.n532 585
R1063 B.n531 B.n34 585
R1064 B.n530 B.n529 585
R1065 B.n528 B.n35 585
R1066 B.n527 B.n526 585
R1067 B.n525 B.n36 585
R1068 B.n524 B.n523 585
R1069 B.n522 B.n37 585
R1070 B.n521 B.n520 585
R1071 B.n519 B.n518 585
R1072 B.n517 B.n41 585
R1073 B.n516 B.n515 585
R1074 B.n514 B.n42 585
R1075 B.n513 B.n512 585
R1076 B.n511 B.n43 585
R1077 B.n510 B.n509 585
R1078 B.n508 B.n44 585
R1079 B.n507 B.n506 585
R1080 B.n504 B.n45 585
R1081 B.n503 B.n502 585
R1082 B.n501 B.n48 585
R1083 B.n500 B.n499 585
R1084 B.n498 B.n49 585
R1085 B.n497 B.n496 585
R1086 B.n495 B.n50 585
R1087 B.n494 B.n493 585
R1088 B.n492 B.n51 585
R1089 B.n491 B.n490 585
R1090 B.n489 B.n52 585
R1091 B.n488 B.n487 585
R1092 B.n486 B.n53 585
R1093 B.n485 B.n484 585
R1094 B.n483 B.n54 585
R1095 B.n482 B.n481 585
R1096 B.n480 B.n55 585
R1097 B.n479 B.n478 585
R1098 B.n477 B.n56 585
R1099 B.n476 B.n475 585
R1100 B.n474 B.n57 585
R1101 B.n473 B.n472 585
R1102 B.n471 B.n58 585
R1103 B.n470 B.n469 585
R1104 B.n468 B.n59 585
R1105 B.n467 B.n466 585
R1106 B.n465 B.n60 585
R1107 B.n464 B.n463 585
R1108 B.n462 B.n61 585
R1109 B.n461 B.n460 585
R1110 B.n459 B.n62 585
R1111 B.n458 B.n457 585
R1112 B.n456 B.n63 585
R1113 B.n455 B.n454 585
R1114 B.n453 B.n64 585
R1115 B.n452 B.n451 585
R1116 B.n450 B.n65 585
R1117 B.n449 B.n448 585
R1118 B.n447 B.n66 585
R1119 B.n446 B.n445 585
R1120 B.n444 B.n67 585
R1121 B.n443 B.n442 585
R1122 B.n441 B.n68 585
R1123 B.n440 B.n439 585
R1124 B.n438 B.n69 585
R1125 B.n437 B.n436 585
R1126 B.n435 B.n70 585
R1127 B.n434 B.n433 585
R1128 B.n432 B.n71 585
R1129 B.n431 B.n430 585
R1130 B.n429 B.n72 585
R1131 B.n428 B.n427 585
R1132 B.n426 B.n73 585
R1133 B.n425 B.n424 585
R1134 B.n602 B.n601 585
R1135 B.n603 B.n10 585
R1136 B.n605 B.n604 585
R1137 B.n606 B.n9 585
R1138 B.n608 B.n607 585
R1139 B.n609 B.n8 585
R1140 B.n611 B.n610 585
R1141 B.n612 B.n7 585
R1142 B.n614 B.n613 585
R1143 B.n615 B.n6 585
R1144 B.n617 B.n616 585
R1145 B.n618 B.n5 585
R1146 B.n620 B.n619 585
R1147 B.n621 B.n4 585
R1148 B.n623 B.n622 585
R1149 B.n624 B.n3 585
R1150 B.n626 B.n625 585
R1151 B.n627 B.n0 585
R1152 B.n2 B.n1 585
R1153 B.n165 B.n164 585
R1154 B.n167 B.n166 585
R1155 B.n168 B.n163 585
R1156 B.n170 B.n169 585
R1157 B.n171 B.n162 585
R1158 B.n173 B.n172 585
R1159 B.n174 B.n161 585
R1160 B.n176 B.n175 585
R1161 B.n177 B.n160 585
R1162 B.n179 B.n178 585
R1163 B.n180 B.n159 585
R1164 B.n182 B.n181 585
R1165 B.n183 B.n158 585
R1166 B.n185 B.n184 585
R1167 B.n186 B.n157 585
R1168 B.n188 B.n187 585
R1169 B.n189 B.n156 585
R1170 B.n190 B.n189 487.695
R1171 B.n368 B.n93 487.695
R1172 B.n424 B.n423 487.695
R1173 B.n602 B.n11 487.695
R1174 B.n120 B.t4 465.889
R1175 B.n46 B.t2 465.889
R1176 B.n128 B.t10 465.889
R1177 B.n38 B.t8 465.889
R1178 B.n121 B.t5 448.628
R1179 B.n47 B.t1 448.628
R1180 B.n129 B.t11 448.628
R1181 B.n39 B.t7 448.628
R1182 B.n629 B.n628 256.663
R1183 B.n628 B.n627 235.042
R1184 B.n628 B.n2 235.042
R1185 B.n190 B.n155 163.367
R1186 B.n194 B.n155 163.367
R1187 B.n195 B.n194 163.367
R1188 B.n196 B.n195 163.367
R1189 B.n196 B.n153 163.367
R1190 B.n200 B.n153 163.367
R1191 B.n201 B.n200 163.367
R1192 B.n202 B.n201 163.367
R1193 B.n202 B.n151 163.367
R1194 B.n206 B.n151 163.367
R1195 B.n207 B.n206 163.367
R1196 B.n208 B.n207 163.367
R1197 B.n208 B.n149 163.367
R1198 B.n212 B.n149 163.367
R1199 B.n213 B.n212 163.367
R1200 B.n214 B.n213 163.367
R1201 B.n214 B.n147 163.367
R1202 B.n218 B.n147 163.367
R1203 B.n219 B.n218 163.367
R1204 B.n220 B.n219 163.367
R1205 B.n220 B.n145 163.367
R1206 B.n224 B.n145 163.367
R1207 B.n225 B.n224 163.367
R1208 B.n226 B.n225 163.367
R1209 B.n226 B.n143 163.367
R1210 B.n230 B.n143 163.367
R1211 B.n231 B.n230 163.367
R1212 B.n232 B.n231 163.367
R1213 B.n232 B.n141 163.367
R1214 B.n236 B.n141 163.367
R1215 B.n237 B.n236 163.367
R1216 B.n238 B.n237 163.367
R1217 B.n238 B.n139 163.367
R1218 B.n242 B.n139 163.367
R1219 B.n243 B.n242 163.367
R1220 B.n244 B.n243 163.367
R1221 B.n244 B.n137 163.367
R1222 B.n248 B.n137 163.367
R1223 B.n249 B.n248 163.367
R1224 B.n250 B.n249 163.367
R1225 B.n250 B.n135 163.367
R1226 B.n254 B.n135 163.367
R1227 B.n255 B.n254 163.367
R1228 B.n256 B.n255 163.367
R1229 B.n256 B.n133 163.367
R1230 B.n260 B.n133 163.367
R1231 B.n261 B.n260 163.367
R1232 B.n262 B.n261 163.367
R1233 B.n262 B.n131 163.367
R1234 B.n266 B.n131 163.367
R1235 B.n267 B.n266 163.367
R1236 B.n268 B.n267 163.367
R1237 B.n268 B.n127 163.367
R1238 B.n273 B.n127 163.367
R1239 B.n274 B.n273 163.367
R1240 B.n275 B.n274 163.367
R1241 B.n275 B.n125 163.367
R1242 B.n279 B.n125 163.367
R1243 B.n280 B.n279 163.367
R1244 B.n281 B.n280 163.367
R1245 B.n281 B.n123 163.367
R1246 B.n285 B.n123 163.367
R1247 B.n286 B.n285 163.367
R1248 B.n286 B.n119 163.367
R1249 B.n290 B.n119 163.367
R1250 B.n291 B.n290 163.367
R1251 B.n292 B.n291 163.367
R1252 B.n292 B.n117 163.367
R1253 B.n296 B.n117 163.367
R1254 B.n297 B.n296 163.367
R1255 B.n298 B.n297 163.367
R1256 B.n298 B.n115 163.367
R1257 B.n302 B.n115 163.367
R1258 B.n303 B.n302 163.367
R1259 B.n304 B.n303 163.367
R1260 B.n304 B.n113 163.367
R1261 B.n308 B.n113 163.367
R1262 B.n309 B.n308 163.367
R1263 B.n310 B.n309 163.367
R1264 B.n310 B.n111 163.367
R1265 B.n314 B.n111 163.367
R1266 B.n315 B.n314 163.367
R1267 B.n316 B.n315 163.367
R1268 B.n316 B.n109 163.367
R1269 B.n320 B.n109 163.367
R1270 B.n321 B.n320 163.367
R1271 B.n322 B.n321 163.367
R1272 B.n322 B.n107 163.367
R1273 B.n326 B.n107 163.367
R1274 B.n327 B.n326 163.367
R1275 B.n328 B.n327 163.367
R1276 B.n328 B.n105 163.367
R1277 B.n332 B.n105 163.367
R1278 B.n333 B.n332 163.367
R1279 B.n334 B.n333 163.367
R1280 B.n334 B.n103 163.367
R1281 B.n338 B.n103 163.367
R1282 B.n339 B.n338 163.367
R1283 B.n340 B.n339 163.367
R1284 B.n340 B.n101 163.367
R1285 B.n344 B.n101 163.367
R1286 B.n345 B.n344 163.367
R1287 B.n346 B.n345 163.367
R1288 B.n346 B.n99 163.367
R1289 B.n350 B.n99 163.367
R1290 B.n351 B.n350 163.367
R1291 B.n352 B.n351 163.367
R1292 B.n352 B.n97 163.367
R1293 B.n356 B.n97 163.367
R1294 B.n357 B.n356 163.367
R1295 B.n358 B.n357 163.367
R1296 B.n358 B.n95 163.367
R1297 B.n362 B.n95 163.367
R1298 B.n363 B.n362 163.367
R1299 B.n364 B.n363 163.367
R1300 B.n364 B.n93 163.367
R1301 B.n423 B.n422 163.367
R1302 B.n422 B.n75 163.367
R1303 B.n418 B.n75 163.367
R1304 B.n418 B.n417 163.367
R1305 B.n417 B.n416 163.367
R1306 B.n416 B.n77 163.367
R1307 B.n412 B.n77 163.367
R1308 B.n412 B.n411 163.367
R1309 B.n411 B.n410 163.367
R1310 B.n410 B.n79 163.367
R1311 B.n406 B.n79 163.367
R1312 B.n406 B.n405 163.367
R1313 B.n405 B.n404 163.367
R1314 B.n404 B.n81 163.367
R1315 B.n400 B.n81 163.367
R1316 B.n400 B.n399 163.367
R1317 B.n399 B.n398 163.367
R1318 B.n398 B.n83 163.367
R1319 B.n394 B.n83 163.367
R1320 B.n394 B.n393 163.367
R1321 B.n393 B.n392 163.367
R1322 B.n392 B.n85 163.367
R1323 B.n388 B.n85 163.367
R1324 B.n388 B.n387 163.367
R1325 B.n387 B.n386 163.367
R1326 B.n386 B.n87 163.367
R1327 B.n382 B.n87 163.367
R1328 B.n382 B.n381 163.367
R1329 B.n381 B.n380 163.367
R1330 B.n380 B.n89 163.367
R1331 B.n376 B.n89 163.367
R1332 B.n376 B.n375 163.367
R1333 B.n375 B.n374 163.367
R1334 B.n374 B.n91 163.367
R1335 B.n370 B.n91 163.367
R1336 B.n370 B.n369 163.367
R1337 B.n369 B.n368 163.367
R1338 B.n598 B.n11 163.367
R1339 B.n598 B.n597 163.367
R1340 B.n597 B.n596 163.367
R1341 B.n596 B.n13 163.367
R1342 B.n592 B.n13 163.367
R1343 B.n592 B.n591 163.367
R1344 B.n591 B.n590 163.367
R1345 B.n590 B.n15 163.367
R1346 B.n586 B.n15 163.367
R1347 B.n586 B.n585 163.367
R1348 B.n585 B.n584 163.367
R1349 B.n584 B.n17 163.367
R1350 B.n580 B.n17 163.367
R1351 B.n580 B.n579 163.367
R1352 B.n579 B.n578 163.367
R1353 B.n578 B.n19 163.367
R1354 B.n574 B.n19 163.367
R1355 B.n574 B.n573 163.367
R1356 B.n573 B.n572 163.367
R1357 B.n572 B.n21 163.367
R1358 B.n568 B.n21 163.367
R1359 B.n568 B.n567 163.367
R1360 B.n567 B.n566 163.367
R1361 B.n566 B.n23 163.367
R1362 B.n562 B.n23 163.367
R1363 B.n562 B.n561 163.367
R1364 B.n561 B.n560 163.367
R1365 B.n560 B.n25 163.367
R1366 B.n556 B.n25 163.367
R1367 B.n556 B.n555 163.367
R1368 B.n555 B.n554 163.367
R1369 B.n554 B.n27 163.367
R1370 B.n550 B.n27 163.367
R1371 B.n550 B.n549 163.367
R1372 B.n549 B.n548 163.367
R1373 B.n548 B.n29 163.367
R1374 B.n544 B.n29 163.367
R1375 B.n544 B.n543 163.367
R1376 B.n543 B.n542 163.367
R1377 B.n542 B.n31 163.367
R1378 B.n538 B.n31 163.367
R1379 B.n538 B.n537 163.367
R1380 B.n537 B.n536 163.367
R1381 B.n536 B.n33 163.367
R1382 B.n532 B.n33 163.367
R1383 B.n532 B.n531 163.367
R1384 B.n531 B.n530 163.367
R1385 B.n530 B.n35 163.367
R1386 B.n526 B.n35 163.367
R1387 B.n526 B.n525 163.367
R1388 B.n525 B.n524 163.367
R1389 B.n524 B.n37 163.367
R1390 B.n520 B.n37 163.367
R1391 B.n520 B.n519 163.367
R1392 B.n519 B.n41 163.367
R1393 B.n515 B.n41 163.367
R1394 B.n515 B.n514 163.367
R1395 B.n514 B.n513 163.367
R1396 B.n513 B.n43 163.367
R1397 B.n509 B.n43 163.367
R1398 B.n509 B.n508 163.367
R1399 B.n508 B.n507 163.367
R1400 B.n507 B.n45 163.367
R1401 B.n502 B.n45 163.367
R1402 B.n502 B.n501 163.367
R1403 B.n501 B.n500 163.367
R1404 B.n500 B.n49 163.367
R1405 B.n496 B.n49 163.367
R1406 B.n496 B.n495 163.367
R1407 B.n495 B.n494 163.367
R1408 B.n494 B.n51 163.367
R1409 B.n490 B.n51 163.367
R1410 B.n490 B.n489 163.367
R1411 B.n489 B.n488 163.367
R1412 B.n488 B.n53 163.367
R1413 B.n484 B.n53 163.367
R1414 B.n484 B.n483 163.367
R1415 B.n483 B.n482 163.367
R1416 B.n482 B.n55 163.367
R1417 B.n478 B.n55 163.367
R1418 B.n478 B.n477 163.367
R1419 B.n477 B.n476 163.367
R1420 B.n476 B.n57 163.367
R1421 B.n472 B.n57 163.367
R1422 B.n472 B.n471 163.367
R1423 B.n471 B.n470 163.367
R1424 B.n470 B.n59 163.367
R1425 B.n466 B.n59 163.367
R1426 B.n466 B.n465 163.367
R1427 B.n465 B.n464 163.367
R1428 B.n464 B.n61 163.367
R1429 B.n460 B.n61 163.367
R1430 B.n460 B.n459 163.367
R1431 B.n459 B.n458 163.367
R1432 B.n458 B.n63 163.367
R1433 B.n454 B.n63 163.367
R1434 B.n454 B.n453 163.367
R1435 B.n453 B.n452 163.367
R1436 B.n452 B.n65 163.367
R1437 B.n448 B.n65 163.367
R1438 B.n448 B.n447 163.367
R1439 B.n447 B.n446 163.367
R1440 B.n446 B.n67 163.367
R1441 B.n442 B.n67 163.367
R1442 B.n442 B.n441 163.367
R1443 B.n441 B.n440 163.367
R1444 B.n440 B.n69 163.367
R1445 B.n436 B.n69 163.367
R1446 B.n436 B.n435 163.367
R1447 B.n435 B.n434 163.367
R1448 B.n434 B.n71 163.367
R1449 B.n430 B.n71 163.367
R1450 B.n430 B.n429 163.367
R1451 B.n429 B.n428 163.367
R1452 B.n428 B.n73 163.367
R1453 B.n424 B.n73 163.367
R1454 B.n603 B.n602 163.367
R1455 B.n604 B.n603 163.367
R1456 B.n604 B.n9 163.367
R1457 B.n608 B.n9 163.367
R1458 B.n609 B.n608 163.367
R1459 B.n610 B.n609 163.367
R1460 B.n610 B.n7 163.367
R1461 B.n614 B.n7 163.367
R1462 B.n615 B.n614 163.367
R1463 B.n616 B.n615 163.367
R1464 B.n616 B.n5 163.367
R1465 B.n620 B.n5 163.367
R1466 B.n621 B.n620 163.367
R1467 B.n622 B.n621 163.367
R1468 B.n622 B.n3 163.367
R1469 B.n626 B.n3 163.367
R1470 B.n627 B.n626 163.367
R1471 B.n165 B.n2 163.367
R1472 B.n166 B.n165 163.367
R1473 B.n166 B.n163 163.367
R1474 B.n170 B.n163 163.367
R1475 B.n171 B.n170 163.367
R1476 B.n172 B.n171 163.367
R1477 B.n172 B.n161 163.367
R1478 B.n176 B.n161 163.367
R1479 B.n177 B.n176 163.367
R1480 B.n178 B.n177 163.367
R1481 B.n178 B.n159 163.367
R1482 B.n182 B.n159 163.367
R1483 B.n183 B.n182 163.367
R1484 B.n184 B.n183 163.367
R1485 B.n184 B.n157 163.367
R1486 B.n188 B.n157 163.367
R1487 B.n189 B.n188 163.367
R1488 B.n271 B.n129 59.5399
R1489 B.n122 B.n121 59.5399
R1490 B.n505 B.n47 59.5399
R1491 B.n40 B.n39 59.5399
R1492 B.n601 B.n600 31.6883
R1493 B.n425 B.n74 31.6883
R1494 B.n367 B.n366 31.6883
R1495 B.n191 B.n156 31.6883
R1496 B B.n629 18.0485
R1497 B.n129 B.n128 17.2611
R1498 B.n121 B.n120 17.2611
R1499 B.n47 B.n46 17.2611
R1500 B.n39 B.n38 17.2611
R1501 B.n601 B.n10 10.6151
R1502 B.n605 B.n10 10.6151
R1503 B.n606 B.n605 10.6151
R1504 B.n607 B.n606 10.6151
R1505 B.n607 B.n8 10.6151
R1506 B.n611 B.n8 10.6151
R1507 B.n612 B.n611 10.6151
R1508 B.n613 B.n612 10.6151
R1509 B.n613 B.n6 10.6151
R1510 B.n617 B.n6 10.6151
R1511 B.n618 B.n617 10.6151
R1512 B.n619 B.n618 10.6151
R1513 B.n619 B.n4 10.6151
R1514 B.n623 B.n4 10.6151
R1515 B.n624 B.n623 10.6151
R1516 B.n625 B.n624 10.6151
R1517 B.n625 B.n0 10.6151
R1518 B.n600 B.n599 10.6151
R1519 B.n599 B.n12 10.6151
R1520 B.n595 B.n12 10.6151
R1521 B.n595 B.n594 10.6151
R1522 B.n594 B.n593 10.6151
R1523 B.n593 B.n14 10.6151
R1524 B.n589 B.n14 10.6151
R1525 B.n589 B.n588 10.6151
R1526 B.n588 B.n587 10.6151
R1527 B.n587 B.n16 10.6151
R1528 B.n583 B.n16 10.6151
R1529 B.n583 B.n582 10.6151
R1530 B.n582 B.n581 10.6151
R1531 B.n581 B.n18 10.6151
R1532 B.n577 B.n18 10.6151
R1533 B.n577 B.n576 10.6151
R1534 B.n576 B.n575 10.6151
R1535 B.n575 B.n20 10.6151
R1536 B.n571 B.n20 10.6151
R1537 B.n571 B.n570 10.6151
R1538 B.n570 B.n569 10.6151
R1539 B.n569 B.n22 10.6151
R1540 B.n565 B.n22 10.6151
R1541 B.n565 B.n564 10.6151
R1542 B.n564 B.n563 10.6151
R1543 B.n563 B.n24 10.6151
R1544 B.n559 B.n24 10.6151
R1545 B.n559 B.n558 10.6151
R1546 B.n558 B.n557 10.6151
R1547 B.n557 B.n26 10.6151
R1548 B.n553 B.n26 10.6151
R1549 B.n553 B.n552 10.6151
R1550 B.n552 B.n551 10.6151
R1551 B.n551 B.n28 10.6151
R1552 B.n547 B.n28 10.6151
R1553 B.n547 B.n546 10.6151
R1554 B.n546 B.n545 10.6151
R1555 B.n545 B.n30 10.6151
R1556 B.n541 B.n30 10.6151
R1557 B.n541 B.n540 10.6151
R1558 B.n540 B.n539 10.6151
R1559 B.n539 B.n32 10.6151
R1560 B.n535 B.n32 10.6151
R1561 B.n535 B.n534 10.6151
R1562 B.n534 B.n533 10.6151
R1563 B.n533 B.n34 10.6151
R1564 B.n529 B.n34 10.6151
R1565 B.n529 B.n528 10.6151
R1566 B.n528 B.n527 10.6151
R1567 B.n527 B.n36 10.6151
R1568 B.n523 B.n36 10.6151
R1569 B.n523 B.n522 10.6151
R1570 B.n522 B.n521 10.6151
R1571 B.n518 B.n517 10.6151
R1572 B.n517 B.n516 10.6151
R1573 B.n516 B.n42 10.6151
R1574 B.n512 B.n42 10.6151
R1575 B.n512 B.n511 10.6151
R1576 B.n511 B.n510 10.6151
R1577 B.n510 B.n44 10.6151
R1578 B.n506 B.n44 10.6151
R1579 B.n504 B.n503 10.6151
R1580 B.n503 B.n48 10.6151
R1581 B.n499 B.n48 10.6151
R1582 B.n499 B.n498 10.6151
R1583 B.n498 B.n497 10.6151
R1584 B.n497 B.n50 10.6151
R1585 B.n493 B.n50 10.6151
R1586 B.n493 B.n492 10.6151
R1587 B.n492 B.n491 10.6151
R1588 B.n491 B.n52 10.6151
R1589 B.n487 B.n52 10.6151
R1590 B.n487 B.n486 10.6151
R1591 B.n486 B.n485 10.6151
R1592 B.n485 B.n54 10.6151
R1593 B.n481 B.n54 10.6151
R1594 B.n481 B.n480 10.6151
R1595 B.n480 B.n479 10.6151
R1596 B.n479 B.n56 10.6151
R1597 B.n475 B.n56 10.6151
R1598 B.n475 B.n474 10.6151
R1599 B.n474 B.n473 10.6151
R1600 B.n473 B.n58 10.6151
R1601 B.n469 B.n58 10.6151
R1602 B.n469 B.n468 10.6151
R1603 B.n468 B.n467 10.6151
R1604 B.n467 B.n60 10.6151
R1605 B.n463 B.n60 10.6151
R1606 B.n463 B.n462 10.6151
R1607 B.n462 B.n461 10.6151
R1608 B.n461 B.n62 10.6151
R1609 B.n457 B.n62 10.6151
R1610 B.n457 B.n456 10.6151
R1611 B.n456 B.n455 10.6151
R1612 B.n455 B.n64 10.6151
R1613 B.n451 B.n64 10.6151
R1614 B.n451 B.n450 10.6151
R1615 B.n450 B.n449 10.6151
R1616 B.n449 B.n66 10.6151
R1617 B.n445 B.n66 10.6151
R1618 B.n445 B.n444 10.6151
R1619 B.n444 B.n443 10.6151
R1620 B.n443 B.n68 10.6151
R1621 B.n439 B.n68 10.6151
R1622 B.n439 B.n438 10.6151
R1623 B.n438 B.n437 10.6151
R1624 B.n437 B.n70 10.6151
R1625 B.n433 B.n70 10.6151
R1626 B.n433 B.n432 10.6151
R1627 B.n432 B.n431 10.6151
R1628 B.n431 B.n72 10.6151
R1629 B.n427 B.n72 10.6151
R1630 B.n427 B.n426 10.6151
R1631 B.n426 B.n425 10.6151
R1632 B.n421 B.n74 10.6151
R1633 B.n421 B.n420 10.6151
R1634 B.n420 B.n419 10.6151
R1635 B.n419 B.n76 10.6151
R1636 B.n415 B.n76 10.6151
R1637 B.n415 B.n414 10.6151
R1638 B.n414 B.n413 10.6151
R1639 B.n413 B.n78 10.6151
R1640 B.n409 B.n78 10.6151
R1641 B.n409 B.n408 10.6151
R1642 B.n408 B.n407 10.6151
R1643 B.n407 B.n80 10.6151
R1644 B.n403 B.n80 10.6151
R1645 B.n403 B.n402 10.6151
R1646 B.n402 B.n401 10.6151
R1647 B.n401 B.n82 10.6151
R1648 B.n397 B.n82 10.6151
R1649 B.n397 B.n396 10.6151
R1650 B.n396 B.n395 10.6151
R1651 B.n395 B.n84 10.6151
R1652 B.n391 B.n84 10.6151
R1653 B.n391 B.n390 10.6151
R1654 B.n390 B.n389 10.6151
R1655 B.n389 B.n86 10.6151
R1656 B.n385 B.n86 10.6151
R1657 B.n385 B.n384 10.6151
R1658 B.n384 B.n383 10.6151
R1659 B.n383 B.n88 10.6151
R1660 B.n379 B.n88 10.6151
R1661 B.n379 B.n378 10.6151
R1662 B.n378 B.n377 10.6151
R1663 B.n377 B.n90 10.6151
R1664 B.n373 B.n90 10.6151
R1665 B.n373 B.n372 10.6151
R1666 B.n372 B.n371 10.6151
R1667 B.n371 B.n92 10.6151
R1668 B.n367 B.n92 10.6151
R1669 B.n164 B.n1 10.6151
R1670 B.n167 B.n164 10.6151
R1671 B.n168 B.n167 10.6151
R1672 B.n169 B.n168 10.6151
R1673 B.n169 B.n162 10.6151
R1674 B.n173 B.n162 10.6151
R1675 B.n174 B.n173 10.6151
R1676 B.n175 B.n174 10.6151
R1677 B.n175 B.n160 10.6151
R1678 B.n179 B.n160 10.6151
R1679 B.n180 B.n179 10.6151
R1680 B.n181 B.n180 10.6151
R1681 B.n181 B.n158 10.6151
R1682 B.n185 B.n158 10.6151
R1683 B.n186 B.n185 10.6151
R1684 B.n187 B.n186 10.6151
R1685 B.n187 B.n156 10.6151
R1686 B.n192 B.n191 10.6151
R1687 B.n193 B.n192 10.6151
R1688 B.n193 B.n154 10.6151
R1689 B.n197 B.n154 10.6151
R1690 B.n198 B.n197 10.6151
R1691 B.n199 B.n198 10.6151
R1692 B.n199 B.n152 10.6151
R1693 B.n203 B.n152 10.6151
R1694 B.n204 B.n203 10.6151
R1695 B.n205 B.n204 10.6151
R1696 B.n205 B.n150 10.6151
R1697 B.n209 B.n150 10.6151
R1698 B.n210 B.n209 10.6151
R1699 B.n211 B.n210 10.6151
R1700 B.n211 B.n148 10.6151
R1701 B.n215 B.n148 10.6151
R1702 B.n216 B.n215 10.6151
R1703 B.n217 B.n216 10.6151
R1704 B.n217 B.n146 10.6151
R1705 B.n221 B.n146 10.6151
R1706 B.n222 B.n221 10.6151
R1707 B.n223 B.n222 10.6151
R1708 B.n223 B.n144 10.6151
R1709 B.n227 B.n144 10.6151
R1710 B.n228 B.n227 10.6151
R1711 B.n229 B.n228 10.6151
R1712 B.n229 B.n142 10.6151
R1713 B.n233 B.n142 10.6151
R1714 B.n234 B.n233 10.6151
R1715 B.n235 B.n234 10.6151
R1716 B.n235 B.n140 10.6151
R1717 B.n239 B.n140 10.6151
R1718 B.n240 B.n239 10.6151
R1719 B.n241 B.n240 10.6151
R1720 B.n241 B.n138 10.6151
R1721 B.n245 B.n138 10.6151
R1722 B.n246 B.n245 10.6151
R1723 B.n247 B.n246 10.6151
R1724 B.n247 B.n136 10.6151
R1725 B.n251 B.n136 10.6151
R1726 B.n252 B.n251 10.6151
R1727 B.n253 B.n252 10.6151
R1728 B.n253 B.n134 10.6151
R1729 B.n257 B.n134 10.6151
R1730 B.n258 B.n257 10.6151
R1731 B.n259 B.n258 10.6151
R1732 B.n259 B.n132 10.6151
R1733 B.n263 B.n132 10.6151
R1734 B.n264 B.n263 10.6151
R1735 B.n265 B.n264 10.6151
R1736 B.n265 B.n130 10.6151
R1737 B.n269 B.n130 10.6151
R1738 B.n270 B.n269 10.6151
R1739 B.n272 B.n126 10.6151
R1740 B.n276 B.n126 10.6151
R1741 B.n277 B.n276 10.6151
R1742 B.n278 B.n277 10.6151
R1743 B.n278 B.n124 10.6151
R1744 B.n282 B.n124 10.6151
R1745 B.n283 B.n282 10.6151
R1746 B.n284 B.n283 10.6151
R1747 B.n288 B.n287 10.6151
R1748 B.n289 B.n288 10.6151
R1749 B.n289 B.n118 10.6151
R1750 B.n293 B.n118 10.6151
R1751 B.n294 B.n293 10.6151
R1752 B.n295 B.n294 10.6151
R1753 B.n295 B.n116 10.6151
R1754 B.n299 B.n116 10.6151
R1755 B.n300 B.n299 10.6151
R1756 B.n301 B.n300 10.6151
R1757 B.n301 B.n114 10.6151
R1758 B.n305 B.n114 10.6151
R1759 B.n306 B.n305 10.6151
R1760 B.n307 B.n306 10.6151
R1761 B.n307 B.n112 10.6151
R1762 B.n311 B.n112 10.6151
R1763 B.n312 B.n311 10.6151
R1764 B.n313 B.n312 10.6151
R1765 B.n313 B.n110 10.6151
R1766 B.n317 B.n110 10.6151
R1767 B.n318 B.n317 10.6151
R1768 B.n319 B.n318 10.6151
R1769 B.n319 B.n108 10.6151
R1770 B.n323 B.n108 10.6151
R1771 B.n324 B.n323 10.6151
R1772 B.n325 B.n324 10.6151
R1773 B.n325 B.n106 10.6151
R1774 B.n329 B.n106 10.6151
R1775 B.n330 B.n329 10.6151
R1776 B.n331 B.n330 10.6151
R1777 B.n331 B.n104 10.6151
R1778 B.n335 B.n104 10.6151
R1779 B.n336 B.n335 10.6151
R1780 B.n337 B.n336 10.6151
R1781 B.n337 B.n102 10.6151
R1782 B.n341 B.n102 10.6151
R1783 B.n342 B.n341 10.6151
R1784 B.n343 B.n342 10.6151
R1785 B.n343 B.n100 10.6151
R1786 B.n347 B.n100 10.6151
R1787 B.n348 B.n347 10.6151
R1788 B.n349 B.n348 10.6151
R1789 B.n349 B.n98 10.6151
R1790 B.n353 B.n98 10.6151
R1791 B.n354 B.n353 10.6151
R1792 B.n355 B.n354 10.6151
R1793 B.n355 B.n96 10.6151
R1794 B.n359 B.n96 10.6151
R1795 B.n360 B.n359 10.6151
R1796 B.n361 B.n360 10.6151
R1797 B.n361 B.n94 10.6151
R1798 B.n365 B.n94 10.6151
R1799 B.n366 B.n365 10.6151
R1800 B.n629 B.n0 8.11757
R1801 B.n629 B.n1 8.11757
R1802 B.n518 B.n40 6.5566
R1803 B.n506 B.n505 6.5566
R1804 B.n272 B.n271 6.5566
R1805 B.n284 B.n122 6.5566
R1806 B.n521 B.n40 4.05904
R1807 B.n505 B.n504 4.05904
R1808 B.n271 B.n270 4.05904
R1809 B.n287 B.n122 4.05904
R1810 VN.n0 VN.t3 788.124
R1811 VN.n4 VN.t1 788.124
R1812 VN.n1 VN.t2 761.303
R1813 VN.n2 VN.t4 761.303
R1814 VN.n5 VN.t5 761.303
R1815 VN.n6 VN.t0 761.303
R1816 VN.n3 VN.n2 161.3
R1817 VN.n7 VN.n6 161.3
R1818 VN.n2 VN.n1 48.2005
R1819 VN.n6 VN.n5 48.2005
R1820 VN.n7 VN.n4 45.1367
R1821 VN.n3 VN.n0 45.1367
R1822 VN VN.n7 44.1577
R1823 VN.n5 VN.n4 13.3799
R1824 VN.n1 VN.n0 13.3799
R1825 VN VN.n3 0.0516364
R1826 VDD2.n175 VDD2.n91 756.745
R1827 VDD2.n84 VDD2.n0 756.745
R1828 VDD2.n176 VDD2.n175 585
R1829 VDD2.n174 VDD2.n173 585
R1830 VDD2.n95 VDD2.n94 585
R1831 VDD2.n168 VDD2.n167 585
R1832 VDD2.n166 VDD2.n97 585
R1833 VDD2.n165 VDD2.n164 585
R1834 VDD2.n100 VDD2.n98 585
R1835 VDD2.n159 VDD2.n158 585
R1836 VDD2.n157 VDD2.n156 585
R1837 VDD2.n104 VDD2.n103 585
R1838 VDD2.n151 VDD2.n150 585
R1839 VDD2.n149 VDD2.n148 585
R1840 VDD2.n108 VDD2.n107 585
R1841 VDD2.n143 VDD2.n142 585
R1842 VDD2.n141 VDD2.n140 585
R1843 VDD2.n112 VDD2.n111 585
R1844 VDD2.n135 VDD2.n134 585
R1845 VDD2.n133 VDD2.n132 585
R1846 VDD2.n116 VDD2.n115 585
R1847 VDD2.n127 VDD2.n126 585
R1848 VDD2.n125 VDD2.n124 585
R1849 VDD2.n120 VDD2.n119 585
R1850 VDD2.n28 VDD2.n27 585
R1851 VDD2.n33 VDD2.n32 585
R1852 VDD2.n35 VDD2.n34 585
R1853 VDD2.n24 VDD2.n23 585
R1854 VDD2.n41 VDD2.n40 585
R1855 VDD2.n43 VDD2.n42 585
R1856 VDD2.n20 VDD2.n19 585
R1857 VDD2.n49 VDD2.n48 585
R1858 VDD2.n51 VDD2.n50 585
R1859 VDD2.n16 VDD2.n15 585
R1860 VDD2.n57 VDD2.n56 585
R1861 VDD2.n59 VDD2.n58 585
R1862 VDD2.n12 VDD2.n11 585
R1863 VDD2.n65 VDD2.n64 585
R1864 VDD2.n67 VDD2.n66 585
R1865 VDD2.n8 VDD2.n7 585
R1866 VDD2.n74 VDD2.n73 585
R1867 VDD2.n75 VDD2.n6 585
R1868 VDD2.n77 VDD2.n76 585
R1869 VDD2.n4 VDD2.n3 585
R1870 VDD2.n83 VDD2.n82 585
R1871 VDD2.n85 VDD2.n84 585
R1872 VDD2.n121 VDD2.t5 327.466
R1873 VDD2.n29 VDD2.t2 327.466
R1874 VDD2.n175 VDD2.n174 171.744
R1875 VDD2.n174 VDD2.n94 171.744
R1876 VDD2.n167 VDD2.n94 171.744
R1877 VDD2.n167 VDD2.n166 171.744
R1878 VDD2.n166 VDD2.n165 171.744
R1879 VDD2.n165 VDD2.n98 171.744
R1880 VDD2.n158 VDD2.n98 171.744
R1881 VDD2.n158 VDD2.n157 171.744
R1882 VDD2.n157 VDD2.n103 171.744
R1883 VDD2.n150 VDD2.n103 171.744
R1884 VDD2.n150 VDD2.n149 171.744
R1885 VDD2.n149 VDD2.n107 171.744
R1886 VDD2.n142 VDD2.n107 171.744
R1887 VDD2.n142 VDD2.n141 171.744
R1888 VDD2.n141 VDD2.n111 171.744
R1889 VDD2.n134 VDD2.n111 171.744
R1890 VDD2.n134 VDD2.n133 171.744
R1891 VDD2.n133 VDD2.n115 171.744
R1892 VDD2.n126 VDD2.n115 171.744
R1893 VDD2.n126 VDD2.n125 171.744
R1894 VDD2.n125 VDD2.n119 171.744
R1895 VDD2.n33 VDD2.n27 171.744
R1896 VDD2.n34 VDD2.n33 171.744
R1897 VDD2.n34 VDD2.n23 171.744
R1898 VDD2.n41 VDD2.n23 171.744
R1899 VDD2.n42 VDD2.n41 171.744
R1900 VDD2.n42 VDD2.n19 171.744
R1901 VDD2.n49 VDD2.n19 171.744
R1902 VDD2.n50 VDD2.n49 171.744
R1903 VDD2.n50 VDD2.n15 171.744
R1904 VDD2.n57 VDD2.n15 171.744
R1905 VDD2.n58 VDD2.n57 171.744
R1906 VDD2.n58 VDD2.n11 171.744
R1907 VDD2.n65 VDD2.n11 171.744
R1908 VDD2.n66 VDD2.n65 171.744
R1909 VDD2.n66 VDD2.n7 171.744
R1910 VDD2.n74 VDD2.n7 171.744
R1911 VDD2.n75 VDD2.n74 171.744
R1912 VDD2.n76 VDD2.n75 171.744
R1913 VDD2.n76 VDD2.n3 171.744
R1914 VDD2.n83 VDD2.n3 171.744
R1915 VDD2.n84 VDD2.n83 171.744
R1916 VDD2.t5 VDD2.n119 85.8723
R1917 VDD2.t2 VDD2.n27 85.8723
R1918 VDD2.n90 VDD2.n89 69.5505
R1919 VDD2 VDD2.n181 69.5477
R1920 VDD2.n90 VDD2.n88 48.9963
R1921 VDD2.n180 VDD2.n179 48.4763
R1922 VDD2.n180 VDD2.n90 40.0537
R1923 VDD2.n121 VDD2.n120 16.3895
R1924 VDD2.n29 VDD2.n28 16.3895
R1925 VDD2.n168 VDD2.n97 13.1884
R1926 VDD2.n77 VDD2.n6 13.1884
R1927 VDD2.n169 VDD2.n95 12.8005
R1928 VDD2.n164 VDD2.n99 12.8005
R1929 VDD2.n124 VDD2.n123 12.8005
R1930 VDD2.n32 VDD2.n31 12.8005
R1931 VDD2.n73 VDD2.n72 12.8005
R1932 VDD2.n78 VDD2.n4 12.8005
R1933 VDD2.n173 VDD2.n172 12.0247
R1934 VDD2.n163 VDD2.n100 12.0247
R1935 VDD2.n127 VDD2.n118 12.0247
R1936 VDD2.n35 VDD2.n26 12.0247
R1937 VDD2.n71 VDD2.n8 12.0247
R1938 VDD2.n82 VDD2.n81 12.0247
R1939 VDD2.n176 VDD2.n93 11.249
R1940 VDD2.n160 VDD2.n159 11.249
R1941 VDD2.n128 VDD2.n116 11.249
R1942 VDD2.n36 VDD2.n24 11.249
R1943 VDD2.n68 VDD2.n67 11.249
R1944 VDD2.n85 VDD2.n2 11.249
R1945 VDD2.n177 VDD2.n91 10.4732
R1946 VDD2.n156 VDD2.n102 10.4732
R1947 VDD2.n132 VDD2.n131 10.4732
R1948 VDD2.n40 VDD2.n39 10.4732
R1949 VDD2.n64 VDD2.n10 10.4732
R1950 VDD2.n86 VDD2.n0 10.4732
R1951 VDD2.n155 VDD2.n104 9.69747
R1952 VDD2.n135 VDD2.n114 9.69747
R1953 VDD2.n43 VDD2.n22 9.69747
R1954 VDD2.n63 VDD2.n12 9.69747
R1955 VDD2.n179 VDD2.n178 9.45567
R1956 VDD2.n88 VDD2.n87 9.45567
R1957 VDD2.n147 VDD2.n146 9.3005
R1958 VDD2.n106 VDD2.n105 9.3005
R1959 VDD2.n153 VDD2.n152 9.3005
R1960 VDD2.n155 VDD2.n154 9.3005
R1961 VDD2.n102 VDD2.n101 9.3005
R1962 VDD2.n161 VDD2.n160 9.3005
R1963 VDD2.n163 VDD2.n162 9.3005
R1964 VDD2.n99 VDD2.n96 9.3005
R1965 VDD2.n178 VDD2.n177 9.3005
R1966 VDD2.n93 VDD2.n92 9.3005
R1967 VDD2.n172 VDD2.n171 9.3005
R1968 VDD2.n170 VDD2.n169 9.3005
R1969 VDD2.n145 VDD2.n144 9.3005
R1970 VDD2.n110 VDD2.n109 9.3005
R1971 VDD2.n139 VDD2.n138 9.3005
R1972 VDD2.n137 VDD2.n136 9.3005
R1973 VDD2.n114 VDD2.n113 9.3005
R1974 VDD2.n131 VDD2.n130 9.3005
R1975 VDD2.n129 VDD2.n128 9.3005
R1976 VDD2.n118 VDD2.n117 9.3005
R1977 VDD2.n123 VDD2.n122 9.3005
R1978 VDD2.n87 VDD2.n86 9.3005
R1979 VDD2.n2 VDD2.n1 9.3005
R1980 VDD2.n81 VDD2.n80 9.3005
R1981 VDD2.n79 VDD2.n78 9.3005
R1982 VDD2.n18 VDD2.n17 9.3005
R1983 VDD2.n47 VDD2.n46 9.3005
R1984 VDD2.n45 VDD2.n44 9.3005
R1985 VDD2.n22 VDD2.n21 9.3005
R1986 VDD2.n39 VDD2.n38 9.3005
R1987 VDD2.n37 VDD2.n36 9.3005
R1988 VDD2.n26 VDD2.n25 9.3005
R1989 VDD2.n31 VDD2.n30 9.3005
R1990 VDD2.n53 VDD2.n52 9.3005
R1991 VDD2.n55 VDD2.n54 9.3005
R1992 VDD2.n14 VDD2.n13 9.3005
R1993 VDD2.n61 VDD2.n60 9.3005
R1994 VDD2.n63 VDD2.n62 9.3005
R1995 VDD2.n10 VDD2.n9 9.3005
R1996 VDD2.n69 VDD2.n68 9.3005
R1997 VDD2.n71 VDD2.n70 9.3005
R1998 VDD2.n72 VDD2.n5 9.3005
R1999 VDD2.n152 VDD2.n151 8.92171
R2000 VDD2.n136 VDD2.n112 8.92171
R2001 VDD2.n44 VDD2.n20 8.92171
R2002 VDD2.n60 VDD2.n59 8.92171
R2003 VDD2.n148 VDD2.n106 8.14595
R2004 VDD2.n140 VDD2.n139 8.14595
R2005 VDD2.n48 VDD2.n47 8.14595
R2006 VDD2.n56 VDD2.n14 8.14595
R2007 VDD2.n147 VDD2.n108 7.3702
R2008 VDD2.n143 VDD2.n110 7.3702
R2009 VDD2.n51 VDD2.n18 7.3702
R2010 VDD2.n55 VDD2.n16 7.3702
R2011 VDD2.n144 VDD2.n108 6.59444
R2012 VDD2.n144 VDD2.n143 6.59444
R2013 VDD2.n52 VDD2.n51 6.59444
R2014 VDD2.n52 VDD2.n16 6.59444
R2015 VDD2.n148 VDD2.n147 5.81868
R2016 VDD2.n140 VDD2.n110 5.81868
R2017 VDD2.n48 VDD2.n18 5.81868
R2018 VDD2.n56 VDD2.n55 5.81868
R2019 VDD2.n151 VDD2.n106 5.04292
R2020 VDD2.n139 VDD2.n112 5.04292
R2021 VDD2.n47 VDD2.n20 5.04292
R2022 VDD2.n59 VDD2.n14 5.04292
R2023 VDD2.n152 VDD2.n104 4.26717
R2024 VDD2.n136 VDD2.n135 4.26717
R2025 VDD2.n44 VDD2.n43 4.26717
R2026 VDD2.n60 VDD2.n12 4.26717
R2027 VDD2.n122 VDD2.n121 3.70982
R2028 VDD2.n30 VDD2.n29 3.70982
R2029 VDD2.n179 VDD2.n91 3.49141
R2030 VDD2.n156 VDD2.n155 3.49141
R2031 VDD2.n132 VDD2.n114 3.49141
R2032 VDD2.n40 VDD2.n22 3.49141
R2033 VDD2.n64 VDD2.n63 3.49141
R2034 VDD2.n88 VDD2.n0 3.49141
R2035 VDD2.n177 VDD2.n176 2.71565
R2036 VDD2.n159 VDD2.n102 2.71565
R2037 VDD2.n131 VDD2.n116 2.71565
R2038 VDD2.n39 VDD2.n24 2.71565
R2039 VDD2.n67 VDD2.n10 2.71565
R2040 VDD2.n86 VDD2.n85 2.71565
R2041 VDD2.n181 VDD2.t0 2.02447
R2042 VDD2.n181 VDD2.t4 2.02447
R2043 VDD2.n89 VDD2.t3 2.02447
R2044 VDD2.n89 VDD2.t1 2.02447
R2045 VDD2.n173 VDD2.n93 1.93989
R2046 VDD2.n160 VDD2.n100 1.93989
R2047 VDD2.n128 VDD2.n127 1.93989
R2048 VDD2.n36 VDD2.n35 1.93989
R2049 VDD2.n68 VDD2.n8 1.93989
R2050 VDD2.n82 VDD2.n2 1.93989
R2051 VDD2.n172 VDD2.n95 1.16414
R2052 VDD2.n164 VDD2.n163 1.16414
R2053 VDD2.n124 VDD2.n118 1.16414
R2054 VDD2.n32 VDD2.n26 1.16414
R2055 VDD2.n73 VDD2.n71 1.16414
R2056 VDD2.n81 VDD2.n4 1.16414
R2057 VDD2 VDD2.n180 0.634121
R2058 VDD2.n169 VDD2.n168 0.388379
R2059 VDD2.n99 VDD2.n97 0.388379
R2060 VDD2.n123 VDD2.n120 0.388379
R2061 VDD2.n31 VDD2.n28 0.388379
R2062 VDD2.n72 VDD2.n6 0.388379
R2063 VDD2.n78 VDD2.n77 0.388379
R2064 VDD2.n178 VDD2.n92 0.155672
R2065 VDD2.n171 VDD2.n92 0.155672
R2066 VDD2.n171 VDD2.n170 0.155672
R2067 VDD2.n170 VDD2.n96 0.155672
R2068 VDD2.n162 VDD2.n96 0.155672
R2069 VDD2.n162 VDD2.n161 0.155672
R2070 VDD2.n161 VDD2.n101 0.155672
R2071 VDD2.n154 VDD2.n101 0.155672
R2072 VDD2.n154 VDD2.n153 0.155672
R2073 VDD2.n153 VDD2.n105 0.155672
R2074 VDD2.n146 VDD2.n105 0.155672
R2075 VDD2.n146 VDD2.n145 0.155672
R2076 VDD2.n145 VDD2.n109 0.155672
R2077 VDD2.n138 VDD2.n109 0.155672
R2078 VDD2.n138 VDD2.n137 0.155672
R2079 VDD2.n137 VDD2.n113 0.155672
R2080 VDD2.n130 VDD2.n113 0.155672
R2081 VDD2.n130 VDD2.n129 0.155672
R2082 VDD2.n129 VDD2.n117 0.155672
R2083 VDD2.n122 VDD2.n117 0.155672
R2084 VDD2.n30 VDD2.n25 0.155672
R2085 VDD2.n37 VDD2.n25 0.155672
R2086 VDD2.n38 VDD2.n37 0.155672
R2087 VDD2.n38 VDD2.n21 0.155672
R2088 VDD2.n45 VDD2.n21 0.155672
R2089 VDD2.n46 VDD2.n45 0.155672
R2090 VDD2.n46 VDD2.n17 0.155672
R2091 VDD2.n53 VDD2.n17 0.155672
R2092 VDD2.n54 VDD2.n53 0.155672
R2093 VDD2.n54 VDD2.n13 0.155672
R2094 VDD2.n61 VDD2.n13 0.155672
R2095 VDD2.n62 VDD2.n61 0.155672
R2096 VDD2.n62 VDD2.n9 0.155672
R2097 VDD2.n69 VDD2.n9 0.155672
R2098 VDD2.n70 VDD2.n69 0.155672
R2099 VDD2.n70 VDD2.n5 0.155672
R2100 VDD2.n79 VDD2.n5 0.155672
R2101 VDD2.n80 VDD2.n79 0.155672
R2102 VDD2.n80 VDD2.n1 0.155672
R2103 VDD2.n87 VDD2.n1 0.155672
C0 B VTAIL 3.31502f
C1 VN VTAIL 4.54535f
C2 VDD1 w_n1682_n4180# 2.07475f
C3 VP B 1.12698f
C4 VN VP 5.6938f
C5 VDD1 VDD2 0.662413f
C6 VTAIL w_n1682_n4180# 3.604f
C7 VP w_n1682_n4180# 2.97513f
C8 VTAIL VDD2 13.915501f
C9 VN B 0.783668f
C10 VP VDD2 0.286871f
C11 VDD1 VTAIL 13.8854f
C12 VDD1 VP 5.19709f
C13 B w_n1682_n4180# 7.99933f
C14 VN w_n1682_n4180# 2.76336f
C15 B VDD2 1.83376f
C16 VN VDD2 5.06478f
C17 VP VTAIL 4.56019f
C18 VDD1 B 1.80807f
C19 VDD1 VN 0.148339f
C20 w_n1682_n4180# VDD2 2.09447f
C21 VDD2 VSUBS 1.528067f
C22 VDD1 VSUBS 1.254221f
C23 VTAIL VSUBS 0.824501f
C24 VN VSUBS 4.78117f
C25 VP VSUBS 1.515979f
C26 B VSUBS 2.958539f
C27 w_n1682_n4180# VSUBS 86.12511f
C28 VDD2.n0 VSUBS 0.027926f
C29 VDD2.n1 VSUBS 0.026975f
C30 VDD2.n2 VSUBS 0.014495f
C31 VDD2.n3 VSUBS 0.034261f
C32 VDD2.n4 VSUBS 0.015348f
C33 VDD2.n5 VSUBS 0.026975f
C34 VDD2.n6 VSUBS 0.014922f
C35 VDD2.n7 VSUBS 0.034261f
C36 VDD2.n8 VSUBS 0.015348f
C37 VDD2.n9 VSUBS 0.026975f
C38 VDD2.n10 VSUBS 0.014495f
C39 VDD2.n11 VSUBS 0.034261f
C40 VDD2.n12 VSUBS 0.015348f
C41 VDD2.n13 VSUBS 0.026975f
C42 VDD2.n14 VSUBS 0.014495f
C43 VDD2.n15 VSUBS 0.034261f
C44 VDD2.n16 VSUBS 0.015348f
C45 VDD2.n17 VSUBS 0.026975f
C46 VDD2.n18 VSUBS 0.014495f
C47 VDD2.n19 VSUBS 0.034261f
C48 VDD2.n20 VSUBS 0.015348f
C49 VDD2.n21 VSUBS 0.026975f
C50 VDD2.n22 VSUBS 0.014495f
C51 VDD2.n23 VSUBS 0.034261f
C52 VDD2.n24 VSUBS 0.015348f
C53 VDD2.n25 VSUBS 0.026975f
C54 VDD2.n26 VSUBS 0.014495f
C55 VDD2.n27 VSUBS 0.025696f
C56 VDD2.n28 VSUBS 0.021796f
C57 VDD2.t2 VSUBS 0.073418f
C58 VDD2.n29 VSUBS 0.198585f
C59 VDD2.n30 VSUBS 1.85222f
C60 VDD2.n31 VSUBS 0.014495f
C61 VDD2.n32 VSUBS 0.015348f
C62 VDD2.n33 VSUBS 0.034261f
C63 VDD2.n34 VSUBS 0.034261f
C64 VDD2.n35 VSUBS 0.015348f
C65 VDD2.n36 VSUBS 0.014495f
C66 VDD2.n37 VSUBS 0.026975f
C67 VDD2.n38 VSUBS 0.026975f
C68 VDD2.n39 VSUBS 0.014495f
C69 VDD2.n40 VSUBS 0.015348f
C70 VDD2.n41 VSUBS 0.034261f
C71 VDD2.n42 VSUBS 0.034261f
C72 VDD2.n43 VSUBS 0.015348f
C73 VDD2.n44 VSUBS 0.014495f
C74 VDD2.n45 VSUBS 0.026975f
C75 VDD2.n46 VSUBS 0.026975f
C76 VDD2.n47 VSUBS 0.014495f
C77 VDD2.n48 VSUBS 0.015348f
C78 VDD2.n49 VSUBS 0.034261f
C79 VDD2.n50 VSUBS 0.034261f
C80 VDD2.n51 VSUBS 0.015348f
C81 VDD2.n52 VSUBS 0.014495f
C82 VDD2.n53 VSUBS 0.026975f
C83 VDD2.n54 VSUBS 0.026975f
C84 VDD2.n55 VSUBS 0.014495f
C85 VDD2.n56 VSUBS 0.015348f
C86 VDD2.n57 VSUBS 0.034261f
C87 VDD2.n58 VSUBS 0.034261f
C88 VDD2.n59 VSUBS 0.015348f
C89 VDD2.n60 VSUBS 0.014495f
C90 VDD2.n61 VSUBS 0.026975f
C91 VDD2.n62 VSUBS 0.026975f
C92 VDD2.n63 VSUBS 0.014495f
C93 VDD2.n64 VSUBS 0.015348f
C94 VDD2.n65 VSUBS 0.034261f
C95 VDD2.n66 VSUBS 0.034261f
C96 VDD2.n67 VSUBS 0.015348f
C97 VDD2.n68 VSUBS 0.014495f
C98 VDD2.n69 VSUBS 0.026975f
C99 VDD2.n70 VSUBS 0.026975f
C100 VDD2.n71 VSUBS 0.014495f
C101 VDD2.n72 VSUBS 0.014495f
C102 VDD2.n73 VSUBS 0.015348f
C103 VDD2.n74 VSUBS 0.034261f
C104 VDD2.n75 VSUBS 0.034261f
C105 VDD2.n76 VSUBS 0.034261f
C106 VDD2.n77 VSUBS 0.014922f
C107 VDD2.n78 VSUBS 0.014495f
C108 VDD2.n79 VSUBS 0.026975f
C109 VDD2.n80 VSUBS 0.026975f
C110 VDD2.n81 VSUBS 0.014495f
C111 VDD2.n82 VSUBS 0.015348f
C112 VDD2.n83 VSUBS 0.034261f
C113 VDD2.n84 VSUBS 0.077106f
C114 VDD2.n85 VSUBS 0.015348f
C115 VDD2.n86 VSUBS 0.014495f
C116 VDD2.n87 VSUBS 0.061615f
C117 VDD2.n88 VSUBS 0.058165f
C118 VDD2.t3 VSUBS 0.342344f
C119 VDD2.t1 VSUBS 0.342344f
C120 VDD2.n89 VSUBS 2.80204f
C121 VDD2.n90 VSUBS 2.5041f
C122 VDD2.n91 VSUBS 0.027926f
C123 VDD2.n92 VSUBS 0.026975f
C124 VDD2.n93 VSUBS 0.014495f
C125 VDD2.n94 VSUBS 0.034261f
C126 VDD2.n95 VSUBS 0.015348f
C127 VDD2.n96 VSUBS 0.026975f
C128 VDD2.n97 VSUBS 0.014922f
C129 VDD2.n98 VSUBS 0.034261f
C130 VDD2.n99 VSUBS 0.014495f
C131 VDD2.n100 VSUBS 0.015348f
C132 VDD2.n101 VSUBS 0.026975f
C133 VDD2.n102 VSUBS 0.014495f
C134 VDD2.n103 VSUBS 0.034261f
C135 VDD2.n104 VSUBS 0.015348f
C136 VDD2.n105 VSUBS 0.026975f
C137 VDD2.n106 VSUBS 0.014495f
C138 VDD2.n107 VSUBS 0.034261f
C139 VDD2.n108 VSUBS 0.015348f
C140 VDD2.n109 VSUBS 0.026975f
C141 VDD2.n110 VSUBS 0.014495f
C142 VDD2.n111 VSUBS 0.034261f
C143 VDD2.n112 VSUBS 0.015348f
C144 VDD2.n113 VSUBS 0.026975f
C145 VDD2.n114 VSUBS 0.014495f
C146 VDD2.n115 VSUBS 0.034261f
C147 VDD2.n116 VSUBS 0.015348f
C148 VDD2.n117 VSUBS 0.026975f
C149 VDD2.n118 VSUBS 0.014495f
C150 VDD2.n119 VSUBS 0.025696f
C151 VDD2.n120 VSUBS 0.021796f
C152 VDD2.t5 VSUBS 0.073418f
C153 VDD2.n121 VSUBS 0.198585f
C154 VDD2.n122 VSUBS 1.85222f
C155 VDD2.n123 VSUBS 0.014495f
C156 VDD2.n124 VSUBS 0.015348f
C157 VDD2.n125 VSUBS 0.034261f
C158 VDD2.n126 VSUBS 0.034261f
C159 VDD2.n127 VSUBS 0.015348f
C160 VDD2.n128 VSUBS 0.014495f
C161 VDD2.n129 VSUBS 0.026975f
C162 VDD2.n130 VSUBS 0.026975f
C163 VDD2.n131 VSUBS 0.014495f
C164 VDD2.n132 VSUBS 0.015348f
C165 VDD2.n133 VSUBS 0.034261f
C166 VDD2.n134 VSUBS 0.034261f
C167 VDD2.n135 VSUBS 0.015348f
C168 VDD2.n136 VSUBS 0.014495f
C169 VDD2.n137 VSUBS 0.026975f
C170 VDD2.n138 VSUBS 0.026975f
C171 VDD2.n139 VSUBS 0.014495f
C172 VDD2.n140 VSUBS 0.015348f
C173 VDD2.n141 VSUBS 0.034261f
C174 VDD2.n142 VSUBS 0.034261f
C175 VDD2.n143 VSUBS 0.015348f
C176 VDD2.n144 VSUBS 0.014495f
C177 VDD2.n145 VSUBS 0.026975f
C178 VDD2.n146 VSUBS 0.026975f
C179 VDD2.n147 VSUBS 0.014495f
C180 VDD2.n148 VSUBS 0.015348f
C181 VDD2.n149 VSUBS 0.034261f
C182 VDD2.n150 VSUBS 0.034261f
C183 VDD2.n151 VSUBS 0.015348f
C184 VDD2.n152 VSUBS 0.014495f
C185 VDD2.n153 VSUBS 0.026975f
C186 VDD2.n154 VSUBS 0.026975f
C187 VDD2.n155 VSUBS 0.014495f
C188 VDD2.n156 VSUBS 0.015348f
C189 VDD2.n157 VSUBS 0.034261f
C190 VDD2.n158 VSUBS 0.034261f
C191 VDD2.n159 VSUBS 0.015348f
C192 VDD2.n160 VSUBS 0.014495f
C193 VDD2.n161 VSUBS 0.026975f
C194 VDD2.n162 VSUBS 0.026975f
C195 VDD2.n163 VSUBS 0.014495f
C196 VDD2.n164 VSUBS 0.015348f
C197 VDD2.n165 VSUBS 0.034261f
C198 VDD2.n166 VSUBS 0.034261f
C199 VDD2.n167 VSUBS 0.034261f
C200 VDD2.n168 VSUBS 0.014922f
C201 VDD2.n169 VSUBS 0.014495f
C202 VDD2.n170 VSUBS 0.026975f
C203 VDD2.n171 VSUBS 0.026975f
C204 VDD2.n172 VSUBS 0.014495f
C205 VDD2.n173 VSUBS 0.015348f
C206 VDD2.n174 VSUBS 0.034261f
C207 VDD2.n175 VSUBS 0.077106f
C208 VDD2.n176 VSUBS 0.015348f
C209 VDD2.n177 VSUBS 0.014495f
C210 VDD2.n178 VSUBS 0.061615f
C211 VDD2.n179 VSUBS 0.057126f
C212 VDD2.n180 VSUBS 2.50329f
C213 VDD2.t0 VSUBS 0.342344f
C214 VDD2.t4 VSUBS 0.342344f
C215 VDD2.n181 VSUBS 2.802f
C216 VN.t3 VSUBS 1.51216f
C217 VN.n0 VSUBS 0.556071f
C218 VN.t2 VSUBS 1.49261f
C219 VN.n1 VSUBS 0.587672f
C220 VN.t4 VSUBS 1.49261f
C221 VN.n2 VSUBS 0.574407f
C222 VN.n3 VSUBS 0.231706f
C223 VN.t1 VSUBS 1.51216f
C224 VN.n4 VSUBS 0.556071f
C225 VN.t5 VSUBS 1.49261f
C226 VN.n5 VSUBS 0.587672f
C227 VN.t0 VSUBS 1.49261f
C228 VN.n6 VSUBS 0.574407f
C229 VN.n7 VSUBS 2.80759f
C230 B.n0 VSUBS 0.006245f
C231 B.n1 VSUBS 0.006245f
C232 B.n2 VSUBS 0.009236f
C233 B.n3 VSUBS 0.007078f
C234 B.n4 VSUBS 0.007078f
C235 B.n5 VSUBS 0.007078f
C236 B.n6 VSUBS 0.007078f
C237 B.n7 VSUBS 0.007078f
C238 B.n8 VSUBS 0.007078f
C239 B.n9 VSUBS 0.007078f
C240 B.n10 VSUBS 0.007078f
C241 B.n11 VSUBS 0.016815f
C242 B.n12 VSUBS 0.007078f
C243 B.n13 VSUBS 0.007078f
C244 B.n14 VSUBS 0.007078f
C245 B.n15 VSUBS 0.007078f
C246 B.n16 VSUBS 0.007078f
C247 B.n17 VSUBS 0.007078f
C248 B.n18 VSUBS 0.007078f
C249 B.n19 VSUBS 0.007078f
C250 B.n20 VSUBS 0.007078f
C251 B.n21 VSUBS 0.007078f
C252 B.n22 VSUBS 0.007078f
C253 B.n23 VSUBS 0.007078f
C254 B.n24 VSUBS 0.007078f
C255 B.n25 VSUBS 0.007078f
C256 B.n26 VSUBS 0.007078f
C257 B.n27 VSUBS 0.007078f
C258 B.n28 VSUBS 0.007078f
C259 B.n29 VSUBS 0.007078f
C260 B.n30 VSUBS 0.007078f
C261 B.n31 VSUBS 0.007078f
C262 B.n32 VSUBS 0.007078f
C263 B.n33 VSUBS 0.007078f
C264 B.n34 VSUBS 0.007078f
C265 B.n35 VSUBS 0.007078f
C266 B.n36 VSUBS 0.007078f
C267 B.n37 VSUBS 0.007078f
C268 B.t7 VSUBS 0.307842f
C269 B.t8 VSUBS 0.318584f
C270 B.t6 VSUBS 0.364008f
C271 B.n38 VSUBS 0.384806f
C272 B.n39 VSUBS 0.300035f
C273 B.n40 VSUBS 0.016399f
C274 B.n41 VSUBS 0.007078f
C275 B.n42 VSUBS 0.007078f
C276 B.n43 VSUBS 0.007078f
C277 B.n44 VSUBS 0.007078f
C278 B.n45 VSUBS 0.007078f
C279 B.t1 VSUBS 0.307845f
C280 B.t2 VSUBS 0.318587f
C281 B.t0 VSUBS 0.364008f
C282 B.n46 VSUBS 0.384802f
C283 B.n47 VSUBS 0.300031f
C284 B.n48 VSUBS 0.007078f
C285 B.n49 VSUBS 0.007078f
C286 B.n50 VSUBS 0.007078f
C287 B.n51 VSUBS 0.007078f
C288 B.n52 VSUBS 0.007078f
C289 B.n53 VSUBS 0.007078f
C290 B.n54 VSUBS 0.007078f
C291 B.n55 VSUBS 0.007078f
C292 B.n56 VSUBS 0.007078f
C293 B.n57 VSUBS 0.007078f
C294 B.n58 VSUBS 0.007078f
C295 B.n59 VSUBS 0.007078f
C296 B.n60 VSUBS 0.007078f
C297 B.n61 VSUBS 0.007078f
C298 B.n62 VSUBS 0.007078f
C299 B.n63 VSUBS 0.007078f
C300 B.n64 VSUBS 0.007078f
C301 B.n65 VSUBS 0.007078f
C302 B.n66 VSUBS 0.007078f
C303 B.n67 VSUBS 0.007078f
C304 B.n68 VSUBS 0.007078f
C305 B.n69 VSUBS 0.007078f
C306 B.n70 VSUBS 0.007078f
C307 B.n71 VSUBS 0.007078f
C308 B.n72 VSUBS 0.007078f
C309 B.n73 VSUBS 0.007078f
C310 B.n74 VSUBS 0.015659f
C311 B.n75 VSUBS 0.007078f
C312 B.n76 VSUBS 0.007078f
C313 B.n77 VSUBS 0.007078f
C314 B.n78 VSUBS 0.007078f
C315 B.n79 VSUBS 0.007078f
C316 B.n80 VSUBS 0.007078f
C317 B.n81 VSUBS 0.007078f
C318 B.n82 VSUBS 0.007078f
C319 B.n83 VSUBS 0.007078f
C320 B.n84 VSUBS 0.007078f
C321 B.n85 VSUBS 0.007078f
C322 B.n86 VSUBS 0.007078f
C323 B.n87 VSUBS 0.007078f
C324 B.n88 VSUBS 0.007078f
C325 B.n89 VSUBS 0.007078f
C326 B.n90 VSUBS 0.007078f
C327 B.n91 VSUBS 0.007078f
C328 B.n92 VSUBS 0.007078f
C329 B.n93 VSUBS 0.016815f
C330 B.n94 VSUBS 0.007078f
C331 B.n95 VSUBS 0.007078f
C332 B.n96 VSUBS 0.007078f
C333 B.n97 VSUBS 0.007078f
C334 B.n98 VSUBS 0.007078f
C335 B.n99 VSUBS 0.007078f
C336 B.n100 VSUBS 0.007078f
C337 B.n101 VSUBS 0.007078f
C338 B.n102 VSUBS 0.007078f
C339 B.n103 VSUBS 0.007078f
C340 B.n104 VSUBS 0.007078f
C341 B.n105 VSUBS 0.007078f
C342 B.n106 VSUBS 0.007078f
C343 B.n107 VSUBS 0.007078f
C344 B.n108 VSUBS 0.007078f
C345 B.n109 VSUBS 0.007078f
C346 B.n110 VSUBS 0.007078f
C347 B.n111 VSUBS 0.007078f
C348 B.n112 VSUBS 0.007078f
C349 B.n113 VSUBS 0.007078f
C350 B.n114 VSUBS 0.007078f
C351 B.n115 VSUBS 0.007078f
C352 B.n116 VSUBS 0.007078f
C353 B.n117 VSUBS 0.007078f
C354 B.n118 VSUBS 0.007078f
C355 B.n119 VSUBS 0.007078f
C356 B.t5 VSUBS 0.307845f
C357 B.t4 VSUBS 0.318587f
C358 B.t3 VSUBS 0.364008f
C359 B.n120 VSUBS 0.384802f
C360 B.n121 VSUBS 0.300031f
C361 B.n122 VSUBS 0.016399f
C362 B.n123 VSUBS 0.007078f
C363 B.n124 VSUBS 0.007078f
C364 B.n125 VSUBS 0.007078f
C365 B.n126 VSUBS 0.007078f
C366 B.n127 VSUBS 0.007078f
C367 B.t11 VSUBS 0.307842f
C368 B.t10 VSUBS 0.318584f
C369 B.t9 VSUBS 0.364008f
C370 B.n128 VSUBS 0.384806f
C371 B.n129 VSUBS 0.300035f
C372 B.n130 VSUBS 0.007078f
C373 B.n131 VSUBS 0.007078f
C374 B.n132 VSUBS 0.007078f
C375 B.n133 VSUBS 0.007078f
C376 B.n134 VSUBS 0.007078f
C377 B.n135 VSUBS 0.007078f
C378 B.n136 VSUBS 0.007078f
C379 B.n137 VSUBS 0.007078f
C380 B.n138 VSUBS 0.007078f
C381 B.n139 VSUBS 0.007078f
C382 B.n140 VSUBS 0.007078f
C383 B.n141 VSUBS 0.007078f
C384 B.n142 VSUBS 0.007078f
C385 B.n143 VSUBS 0.007078f
C386 B.n144 VSUBS 0.007078f
C387 B.n145 VSUBS 0.007078f
C388 B.n146 VSUBS 0.007078f
C389 B.n147 VSUBS 0.007078f
C390 B.n148 VSUBS 0.007078f
C391 B.n149 VSUBS 0.007078f
C392 B.n150 VSUBS 0.007078f
C393 B.n151 VSUBS 0.007078f
C394 B.n152 VSUBS 0.007078f
C395 B.n153 VSUBS 0.007078f
C396 B.n154 VSUBS 0.007078f
C397 B.n155 VSUBS 0.007078f
C398 B.n156 VSUBS 0.015659f
C399 B.n157 VSUBS 0.007078f
C400 B.n158 VSUBS 0.007078f
C401 B.n159 VSUBS 0.007078f
C402 B.n160 VSUBS 0.007078f
C403 B.n161 VSUBS 0.007078f
C404 B.n162 VSUBS 0.007078f
C405 B.n163 VSUBS 0.007078f
C406 B.n164 VSUBS 0.007078f
C407 B.n165 VSUBS 0.007078f
C408 B.n166 VSUBS 0.007078f
C409 B.n167 VSUBS 0.007078f
C410 B.n168 VSUBS 0.007078f
C411 B.n169 VSUBS 0.007078f
C412 B.n170 VSUBS 0.007078f
C413 B.n171 VSUBS 0.007078f
C414 B.n172 VSUBS 0.007078f
C415 B.n173 VSUBS 0.007078f
C416 B.n174 VSUBS 0.007078f
C417 B.n175 VSUBS 0.007078f
C418 B.n176 VSUBS 0.007078f
C419 B.n177 VSUBS 0.007078f
C420 B.n178 VSUBS 0.007078f
C421 B.n179 VSUBS 0.007078f
C422 B.n180 VSUBS 0.007078f
C423 B.n181 VSUBS 0.007078f
C424 B.n182 VSUBS 0.007078f
C425 B.n183 VSUBS 0.007078f
C426 B.n184 VSUBS 0.007078f
C427 B.n185 VSUBS 0.007078f
C428 B.n186 VSUBS 0.007078f
C429 B.n187 VSUBS 0.007078f
C430 B.n188 VSUBS 0.007078f
C431 B.n189 VSUBS 0.015659f
C432 B.n190 VSUBS 0.016815f
C433 B.n191 VSUBS 0.016815f
C434 B.n192 VSUBS 0.007078f
C435 B.n193 VSUBS 0.007078f
C436 B.n194 VSUBS 0.007078f
C437 B.n195 VSUBS 0.007078f
C438 B.n196 VSUBS 0.007078f
C439 B.n197 VSUBS 0.007078f
C440 B.n198 VSUBS 0.007078f
C441 B.n199 VSUBS 0.007078f
C442 B.n200 VSUBS 0.007078f
C443 B.n201 VSUBS 0.007078f
C444 B.n202 VSUBS 0.007078f
C445 B.n203 VSUBS 0.007078f
C446 B.n204 VSUBS 0.007078f
C447 B.n205 VSUBS 0.007078f
C448 B.n206 VSUBS 0.007078f
C449 B.n207 VSUBS 0.007078f
C450 B.n208 VSUBS 0.007078f
C451 B.n209 VSUBS 0.007078f
C452 B.n210 VSUBS 0.007078f
C453 B.n211 VSUBS 0.007078f
C454 B.n212 VSUBS 0.007078f
C455 B.n213 VSUBS 0.007078f
C456 B.n214 VSUBS 0.007078f
C457 B.n215 VSUBS 0.007078f
C458 B.n216 VSUBS 0.007078f
C459 B.n217 VSUBS 0.007078f
C460 B.n218 VSUBS 0.007078f
C461 B.n219 VSUBS 0.007078f
C462 B.n220 VSUBS 0.007078f
C463 B.n221 VSUBS 0.007078f
C464 B.n222 VSUBS 0.007078f
C465 B.n223 VSUBS 0.007078f
C466 B.n224 VSUBS 0.007078f
C467 B.n225 VSUBS 0.007078f
C468 B.n226 VSUBS 0.007078f
C469 B.n227 VSUBS 0.007078f
C470 B.n228 VSUBS 0.007078f
C471 B.n229 VSUBS 0.007078f
C472 B.n230 VSUBS 0.007078f
C473 B.n231 VSUBS 0.007078f
C474 B.n232 VSUBS 0.007078f
C475 B.n233 VSUBS 0.007078f
C476 B.n234 VSUBS 0.007078f
C477 B.n235 VSUBS 0.007078f
C478 B.n236 VSUBS 0.007078f
C479 B.n237 VSUBS 0.007078f
C480 B.n238 VSUBS 0.007078f
C481 B.n239 VSUBS 0.007078f
C482 B.n240 VSUBS 0.007078f
C483 B.n241 VSUBS 0.007078f
C484 B.n242 VSUBS 0.007078f
C485 B.n243 VSUBS 0.007078f
C486 B.n244 VSUBS 0.007078f
C487 B.n245 VSUBS 0.007078f
C488 B.n246 VSUBS 0.007078f
C489 B.n247 VSUBS 0.007078f
C490 B.n248 VSUBS 0.007078f
C491 B.n249 VSUBS 0.007078f
C492 B.n250 VSUBS 0.007078f
C493 B.n251 VSUBS 0.007078f
C494 B.n252 VSUBS 0.007078f
C495 B.n253 VSUBS 0.007078f
C496 B.n254 VSUBS 0.007078f
C497 B.n255 VSUBS 0.007078f
C498 B.n256 VSUBS 0.007078f
C499 B.n257 VSUBS 0.007078f
C500 B.n258 VSUBS 0.007078f
C501 B.n259 VSUBS 0.007078f
C502 B.n260 VSUBS 0.007078f
C503 B.n261 VSUBS 0.007078f
C504 B.n262 VSUBS 0.007078f
C505 B.n263 VSUBS 0.007078f
C506 B.n264 VSUBS 0.007078f
C507 B.n265 VSUBS 0.007078f
C508 B.n266 VSUBS 0.007078f
C509 B.n267 VSUBS 0.007078f
C510 B.n268 VSUBS 0.007078f
C511 B.n269 VSUBS 0.007078f
C512 B.n270 VSUBS 0.004892f
C513 B.n271 VSUBS 0.016399f
C514 B.n272 VSUBS 0.005725f
C515 B.n273 VSUBS 0.007078f
C516 B.n274 VSUBS 0.007078f
C517 B.n275 VSUBS 0.007078f
C518 B.n276 VSUBS 0.007078f
C519 B.n277 VSUBS 0.007078f
C520 B.n278 VSUBS 0.007078f
C521 B.n279 VSUBS 0.007078f
C522 B.n280 VSUBS 0.007078f
C523 B.n281 VSUBS 0.007078f
C524 B.n282 VSUBS 0.007078f
C525 B.n283 VSUBS 0.007078f
C526 B.n284 VSUBS 0.005725f
C527 B.n285 VSUBS 0.007078f
C528 B.n286 VSUBS 0.007078f
C529 B.n287 VSUBS 0.004892f
C530 B.n288 VSUBS 0.007078f
C531 B.n289 VSUBS 0.007078f
C532 B.n290 VSUBS 0.007078f
C533 B.n291 VSUBS 0.007078f
C534 B.n292 VSUBS 0.007078f
C535 B.n293 VSUBS 0.007078f
C536 B.n294 VSUBS 0.007078f
C537 B.n295 VSUBS 0.007078f
C538 B.n296 VSUBS 0.007078f
C539 B.n297 VSUBS 0.007078f
C540 B.n298 VSUBS 0.007078f
C541 B.n299 VSUBS 0.007078f
C542 B.n300 VSUBS 0.007078f
C543 B.n301 VSUBS 0.007078f
C544 B.n302 VSUBS 0.007078f
C545 B.n303 VSUBS 0.007078f
C546 B.n304 VSUBS 0.007078f
C547 B.n305 VSUBS 0.007078f
C548 B.n306 VSUBS 0.007078f
C549 B.n307 VSUBS 0.007078f
C550 B.n308 VSUBS 0.007078f
C551 B.n309 VSUBS 0.007078f
C552 B.n310 VSUBS 0.007078f
C553 B.n311 VSUBS 0.007078f
C554 B.n312 VSUBS 0.007078f
C555 B.n313 VSUBS 0.007078f
C556 B.n314 VSUBS 0.007078f
C557 B.n315 VSUBS 0.007078f
C558 B.n316 VSUBS 0.007078f
C559 B.n317 VSUBS 0.007078f
C560 B.n318 VSUBS 0.007078f
C561 B.n319 VSUBS 0.007078f
C562 B.n320 VSUBS 0.007078f
C563 B.n321 VSUBS 0.007078f
C564 B.n322 VSUBS 0.007078f
C565 B.n323 VSUBS 0.007078f
C566 B.n324 VSUBS 0.007078f
C567 B.n325 VSUBS 0.007078f
C568 B.n326 VSUBS 0.007078f
C569 B.n327 VSUBS 0.007078f
C570 B.n328 VSUBS 0.007078f
C571 B.n329 VSUBS 0.007078f
C572 B.n330 VSUBS 0.007078f
C573 B.n331 VSUBS 0.007078f
C574 B.n332 VSUBS 0.007078f
C575 B.n333 VSUBS 0.007078f
C576 B.n334 VSUBS 0.007078f
C577 B.n335 VSUBS 0.007078f
C578 B.n336 VSUBS 0.007078f
C579 B.n337 VSUBS 0.007078f
C580 B.n338 VSUBS 0.007078f
C581 B.n339 VSUBS 0.007078f
C582 B.n340 VSUBS 0.007078f
C583 B.n341 VSUBS 0.007078f
C584 B.n342 VSUBS 0.007078f
C585 B.n343 VSUBS 0.007078f
C586 B.n344 VSUBS 0.007078f
C587 B.n345 VSUBS 0.007078f
C588 B.n346 VSUBS 0.007078f
C589 B.n347 VSUBS 0.007078f
C590 B.n348 VSUBS 0.007078f
C591 B.n349 VSUBS 0.007078f
C592 B.n350 VSUBS 0.007078f
C593 B.n351 VSUBS 0.007078f
C594 B.n352 VSUBS 0.007078f
C595 B.n353 VSUBS 0.007078f
C596 B.n354 VSUBS 0.007078f
C597 B.n355 VSUBS 0.007078f
C598 B.n356 VSUBS 0.007078f
C599 B.n357 VSUBS 0.007078f
C600 B.n358 VSUBS 0.007078f
C601 B.n359 VSUBS 0.007078f
C602 B.n360 VSUBS 0.007078f
C603 B.n361 VSUBS 0.007078f
C604 B.n362 VSUBS 0.007078f
C605 B.n363 VSUBS 0.007078f
C606 B.n364 VSUBS 0.007078f
C607 B.n365 VSUBS 0.007078f
C608 B.n366 VSUBS 0.015953f
C609 B.n367 VSUBS 0.016521f
C610 B.n368 VSUBS 0.015659f
C611 B.n369 VSUBS 0.007078f
C612 B.n370 VSUBS 0.007078f
C613 B.n371 VSUBS 0.007078f
C614 B.n372 VSUBS 0.007078f
C615 B.n373 VSUBS 0.007078f
C616 B.n374 VSUBS 0.007078f
C617 B.n375 VSUBS 0.007078f
C618 B.n376 VSUBS 0.007078f
C619 B.n377 VSUBS 0.007078f
C620 B.n378 VSUBS 0.007078f
C621 B.n379 VSUBS 0.007078f
C622 B.n380 VSUBS 0.007078f
C623 B.n381 VSUBS 0.007078f
C624 B.n382 VSUBS 0.007078f
C625 B.n383 VSUBS 0.007078f
C626 B.n384 VSUBS 0.007078f
C627 B.n385 VSUBS 0.007078f
C628 B.n386 VSUBS 0.007078f
C629 B.n387 VSUBS 0.007078f
C630 B.n388 VSUBS 0.007078f
C631 B.n389 VSUBS 0.007078f
C632 B.n390 VSUBS 0.007078f
C633 B.n391 VSUBS 0.007078f
C634 B.n392 VSUBS 0.007078f
C635 B.n393 VSUBS 0.007078f
C636 B.n394 VSUBS 0.007078f
C637 B.n395 VSUBS 0.007078f
C638 B.n396 VSUBS 0.007078f
C639 B.n397 VSUBS 0.007078f
C640 B.n398 VSUBS 0.007078f
C641 B.n399 VSUBS 0.007078f
C642 B.n400 VSUBS 0.007078f
C643 B.n401 VSUBS 0.007078f
C644 B.n402 VSUBS 0.007078f
C645 B.n403 VSUBS 0.007078f
C646 B.n404 VSUBS 0.007078f
C647 B.n405 VSUBS 0.007078f
C648 B.n406 VSUBS 0.007078f
C649 B.n407 VSUBS 0.007078f
C650 B.n408 VSUBS 0.007078f
C651 B.n409 VSUBS 0.007078f
C652 B.n410 VSUBS 0.007078f
C653 B.n411 VSUBS 0.007078f
C654 B.n412 VSUBS 0.007078f
C655 B.n413 VSUBS 0.007078f
C656 B.n414 VSUBS 0.007078f
C657 B.n415 VSUBS 0.007078f
C658 B.n416 VSUBS 0.007078f
C659 B.n417 VSUBS 0.007078f
C660 B.n418 VSUBS 0.007078f
C661 B.n419 VSUBS 0.007078f
C662 B.n420 VSUBS 0.007078f
C663 B.n421 VSUBS 0.007078f
C664 B.n422 VSUBS 0.007078f
C665 B.n423 VSUBS 0.015659f
C666 B.n424 VSUBS 0.016815f
C667 B.n425 VSUBS 0.016815f
C668 B.n426 VSUBS 0.007078f
C669 B.n427 VSUBS 0.007078f
C670 B.n428 VSUBS 0.007078f
C671 B.n429 VSUBS 0.007078f
C672 B.n430 VSUBS 0.007078f
C673 B.n431 VSUBS 0.007078f
C674 B.n432 VSUBS 0.007078f
C675 B.n433 VSUBS 0.007078f
C676 B.n434 VSUBS 0.007078f
C677 B.n435 VSUBS 0.007078f
C678 B.n436 VSUBS 0.007078f
C679 B.n437 VSUBS 0.007078f
C680 B.n438 VSUBS 0.007078f
C681 B.n439 VSUBS 0.007078f
C682 B.n440 VSUBS 0.007078f
C683 B.n441 VSUBS 0.007078f
C684 B.n442 VSUBS 0.007078f
C685 B.n443 VSUBS 0.007078f
C686 B.n444 VSUBS 0.007078f
C687 B.n445 VSUBS 0.007078f
C688 B.n446 VSUBS 0.007078f
C689 B.n447 VSUBS 0.007078f
C690 B.n448 VSUBS 0.007078f
C691 B.n449 VSUBS 0.007078f
C692 B.n450 VSUBS 0.007078f
C693 B.n451 VSUBS 0.007078f
C694 B.n452 VSUBS 0.007078f
C695 B.n453 VSUBS 0.007078f
C696 B.n454 VSUBS 0.007078f
C697 B.n455 VSUBS 0.007078f
C698 B.n456 VSUBS 0.007078f
C699 B.n457 VSUBS 0.007078f
C700 B.n458 VSUBS 0.007078f
C701 B.n459 VSUBS 0.007078f
C702 B.n460 VSUBS 0.007078f
C703 B.n461 VSUBS 0.007078f
C704 B.n462 VSUBS 0.007078f
C705 B.n463 VSUBS 0.007078f
C706 B.n464 VSUBS 0.007078f
C707 B.n465 VSUBS 0.007078f
C708 B.n466 VSUBS 0.007078f
C709 B.n467 VSUBS 0.007078f
C710 B.n468 VSUBS 0.007078f
C711 B.n469 VSUBS 0.007078f
C712 B.n470 VSUBS 0.007078f
C713 B.n471 VSUBS 0.007078f
C714 B.n472 VSUBS 0.007078f
C715 B.n473 VSUBS 0.007078f
C716 B.n474 VSUBS 0.007078f
C717 B.n475 VSUBS 0.007078f
C718 B.n476 VSUBS 0.007078f
C719 B.n477 VSUBS 0.007078f
C720 B.n478 VSUBS 0.007078f
C721 B.n479 VSUBS 0.007078f
C722 B.n480 VSUBS 0.007078f
C723 B.n481 VSUBS 0.007078f
C724 B.n482 VSUBS 0.007078f
C725 B.n483 VSUBS 0.007078f
C726 B.n484 VSUBS 0.007078f
C727 B.n485 VSUBS 0.007078f
C728 B.n486 VSUBS 0.007078f
C729 B.n487 VSUBS 0.007078f
C730 B.n488 VSUBS 0.007078f
C731 B.n489 VSUBS 0.007078f
C732 B.n490 VSUBS 0.007078f
C733 B.n491 VSUBS 0.007078f
C734 B.n492 VSUBS 0.007078f
C735 B.n493 VSUBS 0.007078f
C736 B.n494 VSUBS 0.007078f
C737 B.n495 VSUBS 0.007078f
C738 B.n496 VSUBS 0.007078f
C739 B.n497 VSUBS 0.007078f
C740 B.n498 VSUBS 0.007078f
C741 B.n499 VSUBS 0.007078f
C742 B.n500 VSUBS 0.007078f
C743 B.n501 VSUBS 0.007078f
C744 B.n502 VSUBS 0.007078f
C745 B.n503 VSUBS 0.007078f
C746 B.n504 VSUBS 0.004892f
C747 B.n505 VSUBS 0.016399f
C748 B.n506 VSUBS 0.005725f
C749 B.n507 VSUBS 0.007078f
C750 B.n508 VSUBS 0.007078f
C751 B.n509 VSUBS 0.007078f
C752 B.n510 VSUBS 0.007078f
C753 B.n511 VSUBS 0.007078f
C754 B.n512 VSUBS 0.007078f
C755 B.n513 VSUBS 0.007078f
C756 B.n514 VSUBS 0.007078f
C757 B.n515 VSUBS 0.007078f
C758 B.n516 VSUBS 0.007078f
C759 B.n517 VSUBS 0.007078f
C760 B.n518 VSUBS 0.005725f
C761 B.n519 VSUBS 0.007078f
C762 B.n520 VSUBS 0.007078f
C763 B.n521 VSUBS 0.004892f
C764 B.n522 VSUBS 0.007078f
C765 B.n523 VSUBS 0.007078f
C766 B.n524 VSUBS 0.007078f
C767 B.n525 VSUBS 0.007078f
C768 B.n526 VSUBS 0.007078f
C769 B.n527 VSUBS 0.007078f
C770 B.n528 VSUBS 0.007078f
C771 B.n529 VSUBS 0.007078f
C772 B.n530 VSUBS 0.007078f
C773 B.n531 VSUBS 0.007078f
C774 B.n532 VSUBS 0.007078f
C775 B.n533 VSUBS 0.007078f
C776 B.n534 VSUBS 0.007078f
C777 B.n535 VSUBS 0.007078f
C778 B.n536 VSUBS 0.007078f
C779 B.n537 VSUBS 0.007078f
C780 B.n538 VSUBS 0.007078f
C781 B.n539 VSUBS 0.007078f
C782 B.n540 VSUBS 0.007078f
C783 B.n541 VSUBS 0.007078f
C784 B.n542 VSUBS 0.007078f
C785 B.n543 VSUBS 0.007078f
C786 B.n544 VSUBS 0.007078f
C787 B.n545 VSUBS 0.007078f
C788 B.n546 VSUBS 0.007078f
C789 B.n547 VSUBS 0.007078f
C790 B.n548 VSUBS 0.007078f
C791 B.n549 VSUBS 0.007078f
C792 B.n550 VSUBS 0.007078f
C793 B.n551 VSUBS 0.007078f
C794 B.n552 VSUBS 0.007078f
C795 B.n553 VSUBS 0.007078f
C796 B.n554 VSUBS 0.007078f
C797 B.n555 VSUBS 0.007078f
C798 B.n556 VSUBS 0.007078f
C799 B.n557 VSUBS 0.007078f
C800 B.n558 VSUBS 0.007078f
C801 B.n559 VSUBS 0.007078f
C802 B.n560 VSUBS 0.007078f
C803 B.n561 VSUBS 0.007078f
C804 B.n562 VSUBS 0.007078f
C805 B.n563 VSUBS 0.007078f
C806 B.n564 VSUBS 0.007078f
C807 B.n565 VSUBS 0.007078f
C808 B.n566 VSUBS 0.007078f
C809 B.n567 VSUBS 0.007078f
C810 B.n568 VSUBS 0.007078f
C811 B.n569 VSUBS 0.007078f
C812 B.n570 VSUBS 0.007078f
C813 B.n571 VSUBS 0.007078f
C814 B.n572 VSUBS 0.007078f
C815 B.n573 VSUBS 0.007078f
C816 B.n574 VSUBS 0.007078f
C817 B.n575 VSUBS 0.007078f
C818 B.n576 VSUBS 0.007078f
C819 B.n577 VSUBS 0.007078f
C820 B.n578 VSUBS 0.007078f
C821 B.n579 VSUBS 0.007078f
C822 B.n580 VSUBS 0.007078f
C823 B.n581 VSUBS 0.007078f
C824 B.n582 VSUBS 0.007078f
C825 B.n583 VSUBS 0.007078f
C826 B.n584 VSUBS 0.007078f
C827 B.n585 VSUBS 0.007078f
C828 B.n586 VSUBS 0.007078f
C829 B.n587 VSUBS 0.007078f
C830 B.n588 VSUBS 0.007078f
C831 B.n589 VSUBS 0.007078f
C832 B.n590 VSUBS 0.007078f
C833 B.n591 VSUBS 0.007078f
C834 B.n592 VSUBS 0.007078f
C835 B.n593 VSUBS 0.007078f
C836 B.n594 VSUBS 0.007078f
C837 B.n595 VSUBS 0.007078f
C838 B.n596 VSUBS 0.007078f
C839 B.n597 VSUBS 0.007078f
C840 B.n598 VSUBS 0.007078f
C841 B.n599 VSUBS 0.007078f
C842 B.n600 VSUBS 0.016815f
C843 B.n601 VSUBS 0.015659f
C844 B.n602 VSUBS 0.015659f
C845 B.n603 VSUBS 0.007078f
C846 B.n604 VSUBS 0.007078f
C847 B.n605 VSUBS 0.007078f
C848 B.n606 VSUBS 0.007078f
C849 B.n607 VSUBS 0.007078f
C850 B.n608 VSUBS 0.007078f
C851 B.n609 VSUBS 0.007078f
C852 B.n610 VSUBS 0.007078f
C853 B.n611 VSUBS 0.007078f
C854 B.n612 VSUBS 0.007078f
C855 B.n613 VSUBS 0.007078f
C856 B.n614 VSUBS 0.007078f
C857 B.n615 VSUBS 0.007078f
C858 B.n616 VSUBS 0.007078f
C859 B.n617 VSUBS 0.007078f
C860 B.n618 VSUBS 0.007078f
C861 B.n619 VSUBS 0.007078f
C862 B.n620 VSUBS 0.007078f
C863 B.n621 VSUBS 0.007078f
C864 B.n622 VSUBS 0.007078f
C865 B.n623 VSUBS 0.007078f
C866 B.n624 VSUBS 0.007078f
C867 B.n625 VSUBS 0.007078f
C868 B.n626 VSUBS 0.007078f
C869 B.n627 VSUBS 0.009236f
C870 B.n628 VSUBS 0.009839f
C871 B.n629 VSUBS 0.019565f
C872 VDD1.n0 VSUBS 0.027927f
C873 VDD1.n1 VSUBS 0.026976f
C874 VDD1.n2 VSUBS 0.014495f
C875 VDD1.n3 VSUBS 0.034262f
C876 VDD1.n4 VSUBS 0.015348f
C877 VDD1.n5 VSUBS 0.026976f
C878 VDD1.n6 VSUBS 0.014922f
C879 VDD1.n7 VSUBS 0.034262f
C880 VDD1.n8 VSUBS 0.014495f
C881 VDD1.n9 VSUBS 0.015348f
C882 VDD1.n10 VSUBS 0.026976f
C883 VDD1.n11 VSUBS 0.014495f
C884 VDD1.n12 VSUBS 0.034262f
C885 VDD1.n13 VSUBS 0.015348f
C886 VDD1.n14 VSUBS 0.026976f
C887 VDD1.n15 VSUBS 0.014495f
C888 VDD1.n16 VSUBS 0.034262f
C889 VDD1.n17 VSUBS 0.015348f
C890 VDD1.n18 VSUBS 0.026976f
C891 VDD1.n19 VSUBS 0.014495f
C892 VDD1.n20 VSUBS 0.034262f
C893 VDD1.n21 VSUBS 0.015348f
C894 VDD1.n22 VSUBS 0.026976f
C895 VDD1.n23 VSUBS 0.014495f
C896 VDD1.n24 VSUBS 0.034262f
C897 VDD1.n25 VSUBS 0.015348f
C898 VDD1.n26 VSUBS 0.026976f
C899 VDD1.n27 VSUBS 0.014495f
C900 VDD1.n28 VSUBS 0.025697f
C901 VDD1.n29 VSUBS 0.021796f
C902 VDD1.t5 VSUBS 0.073419f
C903 VDD1.n30 VSUBS 0.198589f
C904 VDD1.n31 VSUBS 1.85226f
C905 VDD1.n32 VSUBS 0.014495f
C906 VDD1.n33 VSUBS 0.015348f
C907 VDD1.n34 VSUBS 0.034262f
C908 VDD1.n35 VSUBS 0.034262f
C909 VDD1.n36 VSUBS 0.015348f
C910 VDD1.n37 VSUBS 0.014495f
C911 VDD1.n38 VSUBS 0.026976f
C912 VDD1.n39 VSUBS 0.026976f
C913 VDD1.n40 VSUBS 0.014495f
C914 VDD1.n41 VSUBS 0.015348f
C915 VDD1.n42 VSUBS 0.034262f
C916 VDD1.n43 VSUBS 0.034262f
C917 VDD1.n44 VSUBS 0.015348f
C918 VDD1.n45 VSUBS 0.014495f
C919 VDD1.n46 VSUBS 0.026976f
C920 VDD1.n47 VSUBS 0.026976f
C921 VDD1.n48 VSUBS 0.014495f
C922 VDD1.n49 VSUBS 0.015348f
C923 VDD1.n50 VSUBS 0.034262f
C924 VDD1.n51 VSUBS 0.034262f
C925 VDD1.n52 VSUBS 0.015348f
C926 VDD1.n53 VSUBS 0.014495f
C927 VDD1.n54 VSUBS 0.026976f
C928 VDD1.n55 VSUBS 0.026976f
C929 VDD1.n56 VSUBS 0.014495f
C930 VDD1.n57 VSUBS 0.015348f
C931 VDD1.n58 VSUBS 0.034262f
C932 VDD1.n59 VSUBS 0.034262f
C933 VDD1.n60 VSUBS 0.015348f
C934 VDD1.n61 VSUBS 0.014495f
C935 VDD1.n62 VSUBS 0.026976f
C936 VDD1.n63 VSUBS 0.026976f
C937 VDD1.n64 VSUBS 0.014495f
C938 VDD1.n65 VSUBS 0.015348f
C939 VDD1.n66 VSUBS 0.034262f
C940 VDD1.n67 VSUBS 0.034262f
C941 VDD1.n68 VSUBS 0.015348f
C942 VDD1.n69 VSUBS 0.014495f
C943 VDD1.n70 VSUBS 0.026976f
C944 VDD1.n71 VSUBS 0.026976f
C945 VDD1.n72 VSUBS 0.014495f
C946 VDD1.n73 VSUBS 0.015348f
C947 VDD1.n74 VSUBS 0.034262f
C948 VDD1.n75 VSUBS 0.034262f
C949 VDD1.n76 VSUBS 0.034262f
C950 VDD1.n77 VSUBS 0.014922f
C951 VDD1.n78 VSUBS 0.014495f
C952 VDD1.n79 VSUBS 0.026976f
C953 VDD1.n80 VSUBS 0.026976f
C954 VDD1.n81 VSUBS 0.014495f
C955 VDD1.n82 VSUBS 0.015348f
C956 VDD1.n83 VSUBS 0.034262f
C957 VDD1.n84 VSUBS 0.077108f
C958 VDD1.n85 VSUBS 0.015348f
C959 VDD1.n86 VSUBS 0.014495f
C960 VDD1.n87 VSUBS 0.061616f
C961 VDD1.n88 VSUBS 0.058502f
C962 VDD1.n89 VSUBS 0.027927f
C963 VDD1.n90 VSUBS 0.026976f
C964 VDD1.n91 VSUBS 0.014495f
C965 VDD1.n92 VSUBS 0.034262f
C966 VDD1.n93 VSUBS 0.015348f
C967 VDD1.n94 VSUBS 0.026976f
C968 VDD1.n95 VSUBS 0.014922f
C969 VDD1.n96 VSUBS 0.034262f
C970 VDD1.n97 VSUBS 0.015348f
C971 VDD1.n98 VSUBS 0.026976f
C972 VDD1.n99 VSUBS 0.014495f
C973 VDD1.n100 VSUBS 0.034262f
C974 VDD1.n101 VSUBS 0.015348f
C975 VDD1.n102 VSUBS 0.026976f
C976 VDD1.n103 VSUBS 0.014495f
C977 VDD1.n104 VSUBS 0.034262f
C978 VDD1.n105 VSUBS 0.015348f
C979 VDD1.n106 VSUBS 0.026976f
C980 VDD1.n107 VSUBS 0.014495f
C981 VDD1.n108 VSUBS 0.034262f
C982 VDD1.n109 VSUBS 0.015348f
C983 VDD1.n110 VSUBS 0.026976f
C984 VDD1.n111 VSUBS 0.014495f
C985 VDD1.n112 VSUBS 0.034262f
C986 VDD1.n113 VSUBS 0.015348f
C987 VDD1.n114 VSUBS 0.026976f
C988 VDD1.n115 VSUBS 0.014495f
C989 VDD1.n116 VSUBS 0.025697f
C990 VDD1.n117 VSUBS 0.021796f
C991 VDD1.t4 VSUBS 0.073419f
C992 VDD1.n118 VSUBS 0.198589f
C993 VDD1.n119 VSUBS 1.85226f
C994 VDD1.n120 VSUBS 0.014495f
C995 VDD1.n121 VSUBS 0.015348f
C996 VDD1.n122 VSUBS 0.034262f
C997 VDD1.n123 VSUBS 0.034262f
C998 VDD1.n124 VSUBS 0.015348f
C999 VDD1.n125 VSUBS 0.014495f
C1000 VDD1.n126 VSUBS 0.026976f
C1001 VDD1.n127 VSUBS 0.026976f
C1002 VDD1.n128 VSUBS 0.014495f
C1003 VDD1.n129 VSUBS 0.015348f
C1004 VDD1.n130 VSUBS 0.034262f
C1005 VDD1.n131 VSUBS 0.034262f
C1006 VDD1.n132 VSUBS 0.015348f
C1007 VDD1.n133 VSUBS 0.014495f
C1008 VDD1.n134 VSUBS 0.026976f
C1009 VDD1.n135 VSUBS 0.026976f
C1010 VDD1.n136 VSUBS 0.014495f
C1011 VDD1.n137 VSUBS 0.015348f
C1012 VDD1.n138 VSUBS 0.034262f
C1013 VDD1.n139 VSUBS 0.034262f
C1014 VDD1.n140 VSUBS 0.015348f
C1015 VDD1.n141 VSUBS 0.014495f
C1016 VDD1.n142 VSUBS 0.026976f
C1017 VDD1.n143 VSUBS 0.026976f
C1018 VDD1.n144 VSUBS 0.014495f
C1019 VDD1.n145 VSUBS 0.015348f
C1020 VDD1.n146 VSUBS 0.034262f
C1021 VDD1.n147 VSUBS 0.034262f
C1022 VDD1.n148 VSUBS 0.015348f
C1023 VDD1.n149 VSUBS 0.014495f
C1024 VDD1.n150 VSUBS 0.026976f
C1025 VDD1.n151 VSUBS 0.026976f
C1026 VDD1.n152 VSUBS 0.014495f
C1027 VDD1.n153 VSUBS 0.015348f
C1028 VDD1.n154 VSUBS 0.034262f
C1029 VDD1.n155 VSUBS 0.034262f
C1030 VDD1.n156 VSUBS 0.015348f
C1031 VDD1.n157 VSUBS 0.014495f
C1032 VDD1.n158 VSUBS 0.026976f
C1033 VDD1.n159 VSUBS 0.026976f
C1034 VDD1.n160 VSUBS 0.014495f
C1035 VDD1.n161 VSUBS 0.014495f
C1036 VDD1.n162 VSUBS 0.015348f
C1037 VDD1.n163 VSUBS 0.034262f
C1038 VDD1.n164 VSUBS 0.034262f
C1039 VDD1.n165 VSUBS 0.034262f
C1040 VDD1.n166 VSUBS 0.014922f
C1041 VDD1.n167 VSUBS 0.014495f
C1042 VDD1.n168 VSUBS 0.026976f
C1043 VDD1.n169 VSUBS 0.026976f
C1044 VDD1.n170 VSUBS 0.014495f
C1045 VDD1.n171 VSUBS 0.015348f
C1046 VDD1.n172 VSUBS 0.034262f
C1047 VDD1.n173 VSUBS 0.077108f
C1048 VDD1.n174 VSUBS 0.015348f
C1049 VDD1.n175 VSUBS 0.014495f
C1050 VDD1.n176 VSUBS 0.061616f
C1051 VDD1.n177 VSUBS 0.058166f
C1052 VDD1.t2 VSUBS 0.34235f
C1053 VDD1.t1 VSUBS 0.34235f
C1054 VDD1.n178 VSUBS 2.80208f
C1055 VDD1.n179 VSUBS 2.58491f
C1056 VDD1.t0 VSUBS 0.34235f
C1057 VDD1.t3 VSUBS 0.34235f
C1058 VDD1.n180 VSUBS 2.80087f
C1059 VDD1.n181 VSUBS 3.03005f
C1060 VTAIL.t2 VSUBS 0.37209f
C1061 VTAIL.t5 VSUBS 0.37209f
C1062 VTAIL.n0 VSUBS 2.86538f
C1063 VTAIL.n1 VSUBS 0.814111f
C1064 VTAIL.n2 VSUBS 0.030353f
C1065 VTAIL.n3 VSUBS 0.029319f
C1066 VTAIL.n4 VSUBS 0.015755f
C1067 VTAIL.n5 VSUBS 0.037239f
C1068 VTAIL.n6 VSUBS 0.016681f
C1069 VTAIL.n7 VSUBS 0.029319f
C1070 VTAIL.n8 VSUBS 0.016218f
C1071 VTAIL.n9 VSUBS 0.037239f
C1072 VTAIL.n10 VSUBS 0.016681f
C1073 VTAIL.n11 VSUBS 0.029319f
C1074 VTAIL.n12 VSUBS 0.015755f
C1075 VTAIL.n13 VSUBS 0.037239f
C1076 VTAIL.n14 VSUBS 0.016681f
C1077 VTAIL.n15 VSUBS 0.029319f
C1078 VTAIL.n16 VSUBS 0.015755f
C1079 VTAIL.n17 VSUBS 0.037239f
C1080 VTAIL.n18 VSUBS 0.016681f
C1081 VTAIL.n19 VSUBS 0.029319f
C1082 VTAIL.n20 VSUBS 0.015755f
C1083 VTAIL.n21 VSUBS 0.037239f
C1084 VTAIL.n22 VSUBS 0.016681f
C1085 VTAIL.n23 VSUBS 0.029319f
C1086 VTAIL.n24 VSUBS 0.015755f
C1087 VTAIL.n25 VSUBS 0.037239f
C1088 VTAIL.n26 VSUBS 0.016681f
C1089 VTAIL.n27 VSUBS 0.029319f
C1090 VTAIL.n28 VSUBS 0.015755f
C1091 VTAIL.n29 VSUBS 0.027929f
C1092 VTAIL.n30 VSUBS 0.023689f
C1093 VTAIL.t8 VSUBS 0.079797f
C1094 VTAIL.n31 VSUBS 0.21584f
C1095 VTAIL.n32 VSUBS 2.01316f
C1096 VTAIL.n33 VSUBS 0.015755f
C1097 VTAIL.n34 VSUBS 0.016681f
C1098 VTAIL.n35 VSUBS 0.037239f
C1099 VTAIL.n36 VSUBS 0.037239f
C1100 VTAIL.n37 VSUBS 0.016681f
C1101 VTAIL.n38 VSUBS 0.015755f
C1102 VTAIL.n39 VSUBS 0.029319f
C1103 VTAIL.n40 VSUBS 0.029319f
C1104 VTAIL.n41 VSUBS 0.015755f
C1105 VTAIL.n42 VSUBS 0.016681f
C1106 VTAIL.n43 VSUBS 0.037239f
C1107 VTAIL.n44 VSUBS 0.037239f
C1108 VTAIL.n45 VSUBS 0.016681f
C1109 VTAIL.n46 VSUBS 0.015755f
C1110 VTAIL.n47 VSUBS 0.029319f
C1111 VTAIL.n48 VSUBS 0.029319f
C1112 VTAIL.n49 VSUBS 0.015755f
C1113 VTAIL.n50 VSUBS 0.016681f
C1114 VTAIL.n51 VSUBS 0.037239f
C1115 VTAIL.n52 VSUBS 0.037239f
C1116 VTAIL.n53 VSUBS 0.016681f
C1117 VTAIL.n54 VSUBS 0.015755f
C1118 VTAIL.n55 VSUBS 0.029319f
C1119 VTAIL.n56 VSUBS 0.029319f
C1120 VTAIL.n57 VSUBS 0.015755f
C1121 VTAIL.n58 VSUBS 0.016681f
C1122 VTAIL.n59 VSUBS 0.037239f
C1123 VTAIL.n60 VSUBS 0.037239f
C1124 VTAIL.n61 VSUBS 0.016681f
C1125 VTAIL.n62 VSUBS 0.015755f
C1126 VTAIL.n63 VSUBS 0.029319f
C1127 VTAIL.n64 VSUBS 0.029319f
C1128 VTAIL.n65 VSUBS 0.015755f
C1129 VTAIL.n66 VSUBS 0.016681f
C1130 VTAIL.n67 VSUBS 0.037239f
C1131 VTAIL.n68 VSUBS 0.037239f
C1132 VTAIL.n69 VSUBS 0.016681f
C1133 VTAIL.n70 VSUBS 0.015755f
C1134 VTAIL.n71 VSUBS 0.029319f
C1135 VTAIL.n72 VSUBS 0.029319f
C1136 VTAIL.n73 VSUBS 0.015755f
C1137 VTAIL.n74 VSUBS 0.015755f
C1138 VTAIL.n75 VSUBS 0.016681f
C1139 VTAIL.n76 VSUBS 0.037239f
C1140 VTAIL.n77 VSUBS 0.037239f
C1141 VTAIL.n78 VSUBS 0.037239f
C1142 VTAIL.n79 VSUBS 0.016218f
C1143 VTAIL.n80 VSUBS 0.015755f
C1144 VTAIL.n81 VSUBS 0.029319f
C1145 VTAIL.n82 VSUBS 0.029319f
C1146 VTAIL.n83 VSUBS 0.015755f
C1147 VTAIL.n84 VSUBS 0.016681f
C1148 VTAIL.n85 VSUBS 0.037239f
C1149 VTAIL.n86 VSUBS 0.083806f
C1150 VTAIL.n87 VSUBS 0.016681f
C1151 VTAIL.n88 VSUBS 0.015755f
C1152 VTAIL.n89 VSUBS 0.066968f
C1153 VTAIL.n90 VSUBS 0.041839f
C1154 VTAIL.n91 VSUBS 0.177699f
C1155 VTAIL.t10 VSUBS 0.37209f
C1156 VTAIL.t11 VSUBS 0.37209f
C1157 VTAIL.n92 VSUBS 2.86538f
C1158 VTAIL.n93 VSUBS 2.63353f
C1159 VTAIL.t3 VSUBS 0.37209f
C1160 VTAIL.t1 VSUBS 0.37209f
C1161 VTAIL.n94 VSUBS 2.8654f
C1162 VTAIL.n95 VSUBS 2.63351f
C1163 VTAIL.n96 VSUBS 0.030353f
C1164 VTAIL.n97 VSUBS 0.029319f
C1165 VTAIL.n98 VSUBS 0.015755f
C1166 VTAIL.n99 VSUBS 0.037239f
C1167 VTAIL.n100 VSUBS 0.016681f
C1168 VTAIL.n101 VSUBS 0.029319f
C1169 VTAIL.n102 VSUBS 0.016218f
C1170 VTAIL.n103 VSUBS 0.037239f
C1171 VTAIL.n104 VSUBS 0.015755f
C1172 VTAIL.n105 VSUBS 0.016681f
C1173 VTAIL.n106 VSUBS 0.029319f
C1174 VTAIL.n107 VSUBS 0.015755f
C1175 VTAIL.n108 VSUBS 0.037239f
C1176 VTAIL.n109 VSUBS 0.016681f
C1177 VTAIL.n110 VSUBS 0.029319f
C1178 VTAIL.n111 VSUBS 0.015755f
C1179 VTAIL.n112 VSUBS 0.037239f
C1180 VTAIL.n113 VSUBS 0.016681f
C1181 VTAIL.n114 VSUBS 0.029319f
C1182 VTAIL.n115 VSUBS 0.015755f
C1183 VTAIL.n116 VSUBS 0.037239f
C1184 VTAIL.n117 VSUBS 0.016681f
C1185 VTAIL.n118 VSUBS 0.029319f
C1186 VTAIL.n119 VSUBS 0.015755f
C1187 VTAIL.n120 VSUBS 0.037239f
C1188 VTAIL.n121 VSUBS 0.016681f
C1189 VTAIL.n122 VSUBS 0.029319f
C1190 VTAIL.n123 VSUBS 0.015755f
C1191 VTAIL.n124 VSUBS 0.027929f
C1192 VTAIL.n125 VSUBS 0.023689f
C1193 VTAIL.t4 VSUBS 0.079797f
C1194 VTAIL.n126 VSUBS 0.21584f
C1195 VTAIL.n127 VSUBS 2.01316f
C1196 VTAIL.n128 VSUBS 0.015755f
C1197 VTAIL.n129 VSUBS 0.016681f
C1198 VTAIL.n130 VSUBS 0.037239f
C1199 VTAIL.n131 VSUBS 0.037239f
C1200 VTAIL.n132 VSUBS 0.016681f
C1201 VTAIL.n133 VSUBS 0.015755f
C1202 VTAIL.n134 VSUBS 0.029319f
C1203 VTAIL.n135 VSUBS 0.029319f
C1204 VTAIL.n136 VSUBS 0.015755f
C1205 VTAIL.n137 VSUBS 0.016681f
C1206 VTAIL.n138 VSUBS 0.037239f
C1207 VTAIL.n139 VSUBS 0.037239f
C1208 VTAIL.n140 VSUBS 0.016681f
C1209 VTAIL.n141 VSUBS 0.015755f
C1210 VTAIL.n142 VSUBS 0.029319f
C1211 VTAIL.n143 VSUBS 0.029319f
C1212 VTAIL.n144 VSUBS 0.015755f
C1213 VTAIL.n145 VSUBS 0.016681f
C1214 VTAIL.n146 VSUBS 0.037239f
C1215 VTAIL.n147 VSUBS 0.037239f
C1216 VTAIL.n148 VSUBS 0.016681f
C1217 VTAIL.n149 VSUBS 0.015755f
C1218 VTAIL.n150 VSUBS 0.029319f
C1219 VTAIL.n151 VSUBS 0.029319f
C1220 VTAIL.n152 VSUBS 0.015755f
C1221 VTAIL.n153 VSUBS 0.016681f
C1222 VTAIL.n154 VSUBS 0.037239f
C1223 VTAIL.n155 VSUBS 0.037239f
C1224 VTAIL.n156 VSUBS 0.016681f
C1225 VTAIL.n157 VSUBS 0.015755f
C1226 VTAIL.n158 VSUBS 0.029319f
C1227 VTAIL.n159 VSUBS 0.029319f
C1228 VTAIL.n160 VSUBS 0.015755f
C1229 VTAIL.n161 VSUBS 0.016681f
C1230 VTAIL.n162 VSUBS 0.037239f
C1231 VTAIL.n163 VSUBS 0.037239f
C1232 VTAIL.n164 VSUBS 0.016681f
C1233 VTAIL.n165 VSUBS 0.015755f
C1234 VTAIL.n166 VSUBS 0.029319f
C1235 VTAIL.n167 VSUBS 0.029319f
C1236 VTAIL.n168 VSUBS 0.015755f
C1237 VTAIL.n169 VSUBS 0.016681f
C1238 VTAIL.n170 VSUBS 0.037239f
C1239 VTAIL.n171 VSUBS 0.037239f
C1240 VTAIL.n172 VSUBS 0.037239f
C1241 VTAIL.n173 VSUBS 0.016218f
C1242 VTAIL.n174 VSUBS 0.015755f
C1243 VTAIL.n175 VSUBS 0.029319f
C1244 VTAIL.n176 VSUBS 0.029319f
C1245 VTAIL.n177 VSUBS 0.015755f
C1246 VTAIL.n178 VSUBS 0.016681f
C1247 VTAIL.n179 VSUBS 0.037239f
C1248 VTAIL.n180 VSUBS 0.083806f
C1249 VTAIL.n181 VSUBS 0.016681f
C1250 VTAIL.n182 VSUBS 0.015755f
C1251 VTAIL.n183 VSUBS 0.066968f
C1252 VTAIL.n184 VSUBS 0.041839f
C1253 VTAIL.n185 VSUBS 0.177699f
C1254 VTAIL.t9 VSUBS 0.37209f
C1255 VTAIL.t7 VSUBS 0.37209f
C1256 VTAIL.n186 VSUBS 2.8654f
C1257 VTAIL.n187 VSUBS 0.862957f
C1258 VTAIL.n188 VSUBS 0.030353f
C1259 VTAIL.n189 VSUBS 0.029319f
C1260 VTAIL.n190 VSUBS 0.015755f
C1261 VTAIL.n191 VSUBS 0.037239f
C1262 VTAIL.n192 VSUBS 0.016681f
C1263 VTAIL.n193 VSUBS 0.029319f
C1264 VTAIL.n194 VSUBS 0.016218f
C1265 VTAIL.n195 VSUBS 0.037239f
C1266 VTAIL.n196 VSUBS 0.015755f
C1267 VTAIL.n197 VSUBS 0.016681f
C1268 VTAIL.n198 VSUBS 0.029319f
C1269 VTAIL.n199 VSUBS 0.015755f
C1270 VTAIL.n200 VSUBS 0.037239f
C1271 VTAIL.n201 VSUBS 0.016681f
C1272 VTAIL.n202 VSUBS 0.029319f
C1273 VTAIL.n203 VSUBS 0.015755f
C1274 VTAIL.n204 VSUBS 0.037239f
C1275 VTAIL.n205 VSUBS 0.016681f
C1276 VTAIL.n206 VSUBS 0.029319f
C1277 VTAIL.n207 VSUBS 0.015755f
C1278 VTAIL.n208 VSUBS 0.037239f
C1279 VTAIL.n209 VSUBS 0.016681f
C1280 VTAIL.n210 VSUBS 0.029319f
C1281 VTAIL.n211 VSUBS 0.015755f
C1282 VTAIL.n212 VSUBS 0.037239f
C1283 VTAIL.n213 VSUBS 0.016681f
C1284 VTAIL.n214 VSUBS 0.029319f
C1285 VTAIL.n215 VSUBS 0.015755f
C1286 VTAIL.n216 VSUBS 0.027929f
C1287 VTAIL.n217 VSUBS 0.023689f
C1288 VTAIL.t6 VSUBS 0.079797f
C1289 VTAIL.n218 VSUBS 0.21584f
C1290 VTAIL.n219 VSUBS 2.01316f
C1291 VTAIL.n220 VSUBS 0.015755f
C1292 VTAIL.n221 VSUBS 0.016681f
C1293 VTAIL.n222 VSUBS 0.037239f
C1294 VTAIL.n223 VSUBS 0.037239f
C1295 VTAIL.n224 VSUBS 0.016681f
C1296 VTAIL.n225 VSUBS 0.015755f
C1297 VTAIL.n226 VSUBS 0.029319f
C1298 VTAIL.n227 VSUBS 0.029319f
C1299 VTAIL.n228 VSUBS 0.015755f
C1300 VTAIL.n229 VSUBS 0.016681f
C1301 VTAIL.n230 VSUBS 0.037239f
C1302 VTAIL.n231 VSUBS 0.037239f
C1303 VTAIL.n232 VSUBS 0.016681f
C1304 VTAIL.n233 VSUBS 0.015755f
C1305 VTAIL.n234 VSUBS 0.029319f
C1306 VTAIL.n235 VSUBS 0.029319f
C1307 VTAIL.n236 VSUBS 0.015755f
C1308 VTAIL.n237 VSUBS 0.016681f
C1309 VTAIL.n238 VSUBS 0.037239f
C1310 VTAIL.n239 VSUBS 0.037239f
C1311 VTAIL.n240 VSUBS 0.016681f
C1312 VTAIL.n241 VSUBS 0.015755f
C1313 VTAIL.n242 VSUBS 0.029319f
C1314 VTAIL.n243 VSUBS 0.029319f
C1315 VTAIL.n244 VSUBS 0.015755f
C1316 VTAIL.n245 VSUBS 0.016681f
C1317 VTAIL.n246 VSUBS 0.037239f
C1318 VTAIL.n247 VSUBS 0.037239f
C1319 VTAIL.n248 VSUBS 0.016681f
C1320 VTAIL.n249 VSUBS 0.015755f
C1321 VTAIL.n250 VSUBS 0.029319f
C1322 VTAIL.n251 VSUBS 0.029319f
C1323 VTAIL.n252 VSUBS 0.015755f
C1324 VTAIL.n253 VSUBS 0.016681f
C1325 VTAIL.n254 VSUBS 0.037239f
C1326 VTAIL.n255 VSUBS 0.037239f
C1327 VTAIL.n256 VSUBS 0.016681f
C1328 VTAIL.n257 VSUBS 0.015755f
C1329 VTAIL.n258 VSUBS 0.029319f
C1330 VTAIL.n259 VSUBS 0.029319f
C1331 VTAIL.n260 VSUBS 0.015755f
C1332 VTAIL.n261 VSUBS 0.016681f
C1333 VTAIL.n262 VSUBS 0.037239f
C1334 VTAIL.n263 VSUBS 0.037239f
C1335 VTAIL.n264 VSUBS 0.037239f
C1336 VTAIL.n265 VSUBS 0.016218f
C1337 VTAIL.n266 VSUBS 0.015755f
C1338 VTAIL.n267 VSUBS 0.029319f
C1339 VTAIL.n268 VSUBS 0.029319f
C1340 VTAIL.n269 VSUBS 0.015755f
C1341 VTAIL.n270 VSUBS 0.016681f
C1342 VTAIL.n271 VSUBS 0.037239f
C1343 VTAIL.n272 VSUBS 0.083806f
C1344 VTAIL.n273 VSUBS 0.016681f
C1345 VTAIL.n274 VSUBS 0.015755f
C1346 VTAIL.n275 VSUBS 0.066968f
C1347 VTAIL.n276 VSUBS 0.041839f
C1348 VTAIL.n277 VSUBS 1.87577f
C1349 VTAIL.n278 VSUBS 0.030353f
C1350 VTAIL.n279 VSUBS 0.029319f
C1351 VTAIL.n280 VSUBS 0.015755f
C1352 VTAIL.n281 VSUBS 0.037239f
C1353 VTAIL.n282 VSUBS 0.016681f
C1354 VTAIL.n283 VSUBS 0.029319f
C1355 VTAIL.n284 VSUBS 0.016218f
C1356 VTAIL.n285 VSUBS 0.037239f
C1357 VTAIL.n286 VSUBS 0.016681f
C1358 VTAIL.n287 VSUBS 0.029319f
C1359 VTAIL.n288 VSUBS 0.015755f
C1360 VTAIL.n289 VSUBS 0.037239f
C1361 VTAIL.n290 VSUBS 0.016681f
C1362 VTAIL.n291 VSUBS 0.029319f
C1363 VTAIL.n292 VSUBS 0.015755f
C1364 VTAIL.n293 VSUBS 0.037239f
C1365 VTAIL.n294 VSUBS 0.016681f
C1366 VTAIL.n295 VSUBS 0.029319f
C1367 VTAIL.n296 VSUBS 0.015755f
C1368 VTAIL.n297 VSUBS 0.037239f
C1369 VTAIL.n298 VSUBS 0.016681f
C1370 VTAIL.n299 VSUBS 0.029319f
C1371 VTAIL.n300 VSUBS 0.015755f
C1372 VTAIL.n301 VSUBS 0.037239f
C1373 VTAIL.n302 VSUBS 0.016681f
C1374 VTAIL.n303 VSUBS 0.029319f
C1375 VTAIL.n304 VSUBS 0.015755f
C1376 VTAIL.n305 VSUBS 0.027929f
C1377 VTAIL.n306 VSUBS 0.023689f
C1378 VTAIL.t0 VSUBS 0.079797f
C1379 VTAIL.n307 VSUBS 0.21584f
C1380 VTAIL.n308 VSUBS 2.01316f
C1381 VTAIL.n309 VSUBS 0.015755f
C1382 VTAIL.n310 VSUBS 0.016681f
C1383 VTAIL.n311 VSUBS 0.037239f
C1384 VTAIL.n312 VSUBS 0.037239f
C1385 VTAIL.n313 VSUBS 0.016681f
C1386 VTAIL.n314 VSUBS 0.015755f
C1387 VTAIL.n315 VSUBS 0.029319f
C1388 VTAIL.n316 VSUBS 0.029319f
C1389 VTAIL.n317 VSUBS 0.015755f
C1390 VTAIL.n318 VSUBS 0.016681f
C1391 VTAIL.n319 VSUBS 0.037239f
C1392 VTAIL.n320 VSUBS 0.037239f
C1393 VTAIL.n321 VSUBS 0.016681f
C1394 VTAIL.n322 VSUBS 0.015755f
C1395 VTAIL.n323 VSUBS 0.029319f
C1396 VTAIL.n324 VSUBS 0.029319f
C1397 VTAIL.n325 VSUBS 0.015755f
C1398 VTAIL.n326 VSUBS 0.016681f
C1399 VTAIL.n327 VSUBS 0.037239f
C1400 VTAIL.n328 VSUBS 0.037239f
C1401 VTAIL.n329 VSUBS 0.016681f
C1402 VTAIL.n330 VSUBS 0.015755f
C1403 VTAIL.n331 VSUBS 0.029319f
C1404 VTAIL.n332 VSUBS 0.029319f
C1405 VTAIL.n333 VSUBS 0.015755f
C1406 VTAIL.n334 VSUBS 0.016681f
C1407 VTAIL.n335 VSUBS 0.037239f
C1408 VTAIL.n336 VSUBS 0.037239f
C1409 VTAIL.n337 VSUBS 0.016681f
C1410 VTAIL.n338 VSUBS 0.015755f
C1411 VTAIL.n339 VSUBS 0.029319f
C1412 VTAIL.n340 VSUBS 0.029319f
C1413 VTAIL.n341 VSUBS 0.015755f
C1414 VTAIL.n342 VSUBS 0.016681f
C1415 VTAIL.n343 VSUBS 0.037239f
C1416 VTAIL.n344 VSUBS 0.037239f
C1417 VTAIL.n345 VSUBS 0.016681f
C1418 VTAIL.n346 VSUBS 0.015755f
C1419 VTAIL.n347 VSUBS 0.029319f
C1420 VTAIL.n348 VSUBS 0.029319f
C1421 VTAIL.n349 VSUBS 0.015755f
C1422 VTAIL.n350 VSUBS 0.015755f
C1423 VTAIL.n351 VSUBS 0.016681f
C1424 VTAIL.n352 VSUBS 0.037239f
C1425 VTAIL.n353 VSUBS 0.037239f
C1426 VTAIL.n354 VSUBS 0.037239f
C1427 VTAIL.n355 VSUBS 0.016218f
C1428 VTAIL.n356 VSUBS 0.015755f
C1429 VTAIL.n357 VSUBS 0.029319f
C1430 VTAIL.n358 VSUBS 0.029319f
C1431 VTAIL.n359 VSUBS 0.015755f
C1432 VTAIL.n360 VSUBS 0.016681f
C1433 VTAIL.n361 VSUBS 0.037239f
C1434 VTAIL.n362 VSUBS 0.083806f
C1435 VTAIL.n363 VSUBS 0.016681f
C1436 VTAIL.n364 VSUBS 0.015755f
C1437 VTAIL.n365 VSUBS 0.066968f
C1438 VTAIL.n366 VSUBS 0.041839f
C1439 VTAIL.n367 VSUBS 1.85215f
C1440 VP.n0 VSUBS 0.079902f
C1441 VP.t0 VSUBS 1.55263f
C1442 VP.n1 VSUBS 0.570952f
C1443 VP.t2 VSUBS 1.53255f
C1444 VP.t5 VSUBS 1.53255f
C1445 VP.n2 VSUBS 0.603399f
C1446 VP.n3 VSUBS 0.589779f
C1447 VP.n4 VSUBS 2.84342f
C1448 VP.n5 VSUBS 2.72153f
C1449 VP.t1 VSUBS 1.53255f
C1450 VP.n6 VSUBS 0.589779f
C1451 VP.t3 VSUBS 1.53255f
C1452 VP.n7 VSUBS 0.603399f
C1453 VP.t4 VSUBS 1.53255f
C1454 VP.n8 VSUBS 0.589779f
C1455 VP.n9 VSUBS 0.066583f
.ends

