* NGSPICE file created from diff_pair_sample_0590.ext - technology: sky130A

.subckt diff_pair_sample_0590 VTAIL VN VP B VDD2 VDD1
X0 B.t11 B.t9 B.t10 w_n3666_n3866# sky130_fd_pr__pfet_01v8 ad=5.6511 pd=29.76 as=0 ps=0 w=14.49 l=3.04
X1 VDD1.t5 VP.t0 VTAIL.t8 w_n3666_n3866# sky130_fd_pr__pfet_01v8 ad=2.39085 pd=14.82 as=5.6511 ps=29.76 w=14.49 l=3.04
X2 VTAIL.t6 VP.t1 VDD1.t4 w_n3666_n3866# sky130_fd_pr__pfet_01v8 ad=2.39085 pd=14.82 as=2.39085 ps=14.82 w=14.49 l=3.04
X3 B.t8 B.t6 B.t7 w_n3666_n3866# sky130_fd_pr__pfet_01v8 ad=5.6511 pd=29.76 as=0 ps=0 w=14.49 l=3.04
X4 VTAIL.t7 VP.t2 VDD1.t3 w_n3666_n3866# sky130_fd_pr__pfet_01v8 ad=2.39085 pd=14.82 as=2.39085 ps=14.82 w=14.49 l=3.04
X5 VDD2.t5 VN.t0 VTAIL.t4 w_n3666_n3866# sky130_fd_pr__pfet_01v8 ad=2.39085 pd=14.82 as=5.6511 ps=29.76 w=14.49 l=3.04
X6 VTAIL.t5 VN.t1 VDD2.t4 w_n3666_n3866# sky130_fd_pr__pfet_01v8 ad=2.39085 pd=14.82 as=2.39085 ps=14.82 w=14.49 l=3.04
X7 VDD1.t2 VP.t3 VTAIL.t9 w_n3666_n3866# sky130_fd_pr__pfet_01v8 ad=2.39085 pd=14.82 as=5.6511 ps=29.76 w=14.49 l=3.04
X8 VDD1.t1 VP.t4 VTAIL.t11 w_n3666_n3866# sky130_fd_pr__pfet_01v8 ad=5.6511 pd=29.76 as=2.39085 ps=14.82 w=14.49 l=3.04
X9 B.t5 B.t3 B.t4 w_n3666_n3866# sky130_fd_pr__pfet_01v8 ad=5.6511 pd=29.76 as=0 ps=0 w=14.49 l=3.04
X10 B.t2 B.t0 B.t1 w_n3666_n3866# sky130_fd_pr__pfet_01v8 ad=5.6511 pd=29.76 as=0 ps=0 w=14.49 l=3.04
X11 VTAIL.t3 VN.t2 VDD2.t3 w_n3666_n3866# sky130_fd_pr__pfet_01v8 ad=2.39085 pd=14.82 as=2.39085 ps=14.82 w=14.49 l=3.04
X12 VDD2.t2 VN.t3 VTAIL.t1 w_n3666_n3866# sky130_fd_pr__pfet_01v8 ad=5.6511 pd=29.76 as=2.39085 ps=14.82 w=14.49 l=3.04
X13 VDD2.t1 VN.t4 VTAIL.t2 w_n3666_n3866# sky130_fd_pr__pfet_01v8 ad=2.39085 pd=14.82 as=5.6511 ps=29.76 w=14.49 l=3.04
X14 VDD1.t0 VP.t5 VTAIL.t10 w_n3666_n3866# sky130_fd_pr__pfet_01v8 ad=5.6511 pd=29.76 as=2.39085 ps=14.82 w=14.49 l=3.04
X15 VDD2.t0 VN.t5 VTAIL.t0 w_n3666_n3866# sky130_fd_pr__pfet_01v8 ad=5.6511 pd=29.76 as=2.39085 ps=14.82 w=14.49 l=3.04
R0 B.n443 B.n442 585
R1 B.n441 B.n132 585
R2 B.n440 B.n439 585
R3 B.n438 B.n133 585
R4 B.n437 B.n436 585
R5 B.n435 B.n134 585
R6 B.n434 B.n433 585
R7 B.n432 B.n135 585
R8 B.n431 B.n430 585
R9 B.n429 B.n136 585
R10 B.n428 B.n427 585
R11 B.n426 B.n137 585
R12 B.n425 B.n424 585
R13 B.n423 B.n138 585
R14 B.n422 B.n421 585
R15 B.n420 B.n139 585
R16 B.n419 B.n418 585
R17 B.n417 B.n140 585
R18 B.n416 B.n415 585
R19 B.n414 B.n141 585
R20 B.n413 B.n412 585
R21 B.n411 B.n142 585
R22 B.n410 B.n409 585
R23 B.n408 B.n143 585
R24 B.n407 B.n406 585
R25 B.n405 B.n144 585
R26 B.n404 B.n403 585
R27 B.n402 B.n145 585
R28 B.n401 B.n400 585
R29 B.n399 B.n146 585
R30 B.n398 B.n397 585
R31 B.n396 B.n147 585
R32 B.n395 B.n394 585
R33 B.n393 B.n148 585
R34 B.n392 B.n391 585
R35 B.n390 B.n149 585
R36 B.n389 B.n388 585
R37 B.n387 B.n150 585
R38 B.n386 B.n385 585
R39 B.n384 B.n151 585
R40 B.n383 B.n382 585
R41 B.n381 B.n152 585
R42 B.n380 B.n379 585
R43 B.n378 B.n153 585
R44 B.n377 B.n376 585
R45 B.n375 B.n154 585
R46 B.n374 B.n373 585
R47 B.n372 B.n155 585
R48 B.n371 B.n370 585
R49 B.n369 B.n368 585
R50 B.n367 B.n159 585
R51 B.n366 B.n365 585
R52 B.n364 B.n160 585
R53 B.n363 B.n362 585
R54 B.n361 B.n161 585
R55 B.n360 B.n359 585
R56 B.n358 B.n162 585
R57 B.n357 B.n356 585
R58 B.n354 B.n163 585
R59 B.n353 B.n352 585
R60 B.n351 B.n166 585
R61 B.n350 B.n349 585
R62 B.n348 B.n167 585
R63 B.n347 B.n346 585
R64 B.n345 B.n168 585
R65 B.n344 B.n343 585
R66 B.n342 B.n169 585
R67 B.n341 B.n340 585
R68 B.n339 B.n170 585
R69 B.n338 B.n337 585
R70 B.n336 B.n171 585
R71 B.n335 B.n334 585
R72 B.n333 B.n172 585
R73 B.n332 B.n331 585
R74 B.n330 B.n173 585
R75 B.n329 B.n328 585
R76 B.n327 B.n174 585
R77 B.n326 B.n325 585
R78 B.n324 B.n175 585
R79 B.n323 B.n322 585
R80 B.n321 B.n176 585
R81 B.n320 B.n319 585
R82 B.n318 B.n177 585
R83 B.n317 B.n316 585
R84 B.n315 B.n178 585
R85 B.n314 B.n313 585
R86 B.n312 B.n179 585
R87 B.n311 B.n310 585
R88 B.n309 B.n180 585
R89 B.n308 B.n307 585
R90 B.n306 B.n181 585
R91 B.n305 B.n304 585
R92 B.n303 B.n182 585
R93 B.n302 B.n301 585
R94 B.n300 B.n183 585
R95 B.n299 B.n298 585
R96 B.n297 B.n184 585
R97 B.n296 B.n295 585
R98 B.n294 B.n185 585
R99 B.n293 B.n292 585
R100 B.n291 B.n186 585
R101 B.n290 B.n289 585
R102 B.n288 B.n187 585
R103 B.n287 B.n286 585
R104 B.n285 B.n188 585
R105 B.n284 B.n283 585
R106 B.n282 B.n189 585
R107 B.n444 B.n131 585
R108 B.n446 B.n445 585
R109 B.n447 B.n130 585
R110 B.n449 B.n448 585
R111 B.n450 B.n129 585
R112 B.n452 B.n451 585
R113 B.n453 B.n128 585
R114 B.n455 B.n454 585
R115 B.n456 B.n127 585
R116 B.n458 B.n457 585
R117 B.n459 B.n126 585
R118 B.n461 B.n460 585
R119 B.n462 B.n125 585
R120 B.n464 B.n463 585
R121 B.n465 B.n124 585
R122 B.n467 B.n466 585
R123 B.n468 B.n123 585
R124 B.n470 B.n469 585
R125 B.n471 B.n122 585
R126 B.n473 B.n472 585
R127 B.n474 B.n121 585
R128 B.n476 B.n475 585
R129 B.n477 B.n120 585
R130 B.n479 B.n478 585
R131 B.n480 B.n119 585
R132 B.n482 B.n481 585
R133 B.n483 B.n118 585
R134 B.n485 B.n484 585
R135 B.n486 B.n117 585
R136 B.n488 B.n487 585
R137 B.n489 B.n116 585
R138 B.n491 B.n490 585
R139 B.n492 B.n115 585
R140 B.n494 B.n493 585
R141 B.n495 B.n114 585
R142 B.n497 B.n496 585
R143 B.n498 B.n113 585
R144 B.n500 B.n499 585
R145 B.n501 B.n112 585
R146 B.n503 B.n502 585
R147 B.n504 B.n111 585
R148 B.n506 B.n505 585
R149 B.n507 B.n110 585
R150 B.n509 B.n508 585
R151 B.n510 B.n109 585
R152 B.n512 B.n511 585
R153 B.n513 B.n108 585
R154 B.n515 B.n514 585
R155 B.n516 B.n107 585
R156 B.n518 B.n517 585
R157 B.n519 B.n106 585
R158 B.n521 B.n520 585
R159 B.n522 B.n105 585
R160 B.n524 B.n523 585
R161 B.n525 B.n104 585
R162 B.n527 B.n526 585
R163 B.n528 B.n103 585
R164 B.n530 B.n529 585
R165 B.n531 B.n102 585
R166 B.n533 B.n532 585
R167 B.n534 B.n101 585
R168 B.n536 B.n535 585
R169 B.n537 B.n100 585
R170 B.n539 B.n538 585
R171 B.n540 B.n99 585
R172 B.n542 B.n541 585
R173 B.n543 B.n98 585
R174 B.n545 B.n544 585
R175 B.n546 B.n97 585
R176 B.n548 B.n547 585
R177 B.n549 B.n96 585
R178 B.n551 B.n550 585
R179 B.n552 B.n95 585
R180 B.n554 B.n553 585
R181 B.n555 B.n94 585
R182 B.n557 B.n556 585
R183 B.n558 B.n93 585
R184 B.n560 B.n559 585
R185 B.n561 B.n92 585
R186 B.n563 B.n562 585
R187 B.n564 B.n91 585
R188 B.n566 B.n565 585
R189 B.n567 B.n90 585
R190 B.n569 B.n568 585
R191 B.n570 B.n89 585
R192 B.n572 B.n571 585
R193 B.n573 B.n88 585
R194 B.n575 B.n574 585
R195 B.n576 B.n87 585
R196 B.n578 B.n577 585
R197 B.n579 B.n86 585
R198 B.n581 B.n580 585
R199 B.n582 B.n85 585
R200 B.n584 B.n583 585
R201 B.n585 B.n84 585
R202 B.n587 B.n586 585
R203 B.n749 B.n748 585
R204 B.n747 B.n26 585
R205 B.n746 B.n745 585
R206 B.n744 B.n27 585
R207 B.n743 B.n742 585
R208 B.n741 B.n28 585
R209 B.n740 B.n739 585
R210 B.n738 B.n29 585
R211 B.n737 B.n736 585
R212 B.n735 B.n30 585
R213 B.n734 B.n733 585
R214 B.n732 B.n31 585
R215 B.n731 B.n730 585
R216 B.n729 B.n32 585
R217 B.n728 B.n727 585
R218 B.n726 B.n33 585
R219 B.n725 B.n724 585
R220 B.n723 B.n34 585
R221 B.n722 B.n721 585
R222 B.n720 B.n35 585
R223 B.n719 B.n718 585
R224 B.n717 B.n36 585
R225 B.n716 B.n715 585
R226 B.n714 B.n37 585
R227 B.n713 B.n712 585
R228 B.n711 B.n38 585
R229 B.n710 B.n709 585
R230 B.n708 B.n39 585
R231 B.n707 B.n706 585
R232 B.n705 B.n40 585
R233 B.n704 B.n703 585
R234 B.n702 B.n41 585
R235 B.n701 B.n700 585
R236 B.n699 B.n42 585
R237 B.n698 B.n697 585
R238 B.n696 B.n43 585
R239 B.n695 B.n694 585
R240 B.n693 B.n44 585
R241 B.n692 B.n691 585
R242 B.n690 B.n45 585
R243 B.n689 B.n688 585
R244 B.n687 B.n46 585
R245 B.n686 B.n685 585
R246 B.n684 B.n47 585
R247 B.n683 B.n682 585
R248 B.n681 B.n48 585
R249 B.n680 B.n679 585
R250 B.n678 B.n49 585
R251 B.n677 B.n676 585
R252 B.n675 B.n674 585
R253 B.n673 B.n53 585
R254 B.n672 B.n671 585
R255 B.n670 B.n54 585
R256 B.n669 B.n668 585
R257 B.n667 B.n55 585
R258 B.n666 B.n665 585
R259 B.n664 B.n56 585
R260 B.n663 B.n662 585
R261 B.n660 B.n57 585
R262 B.n659 B.n658 585
R263 B.n657 B.n60 585
R264 B.n656 B.n655 585
R265 B.n654 B.n61 585
R266 B.n653 B.n652 585
R267 B.n651 B.n62 585
R268 B.n650 B.n649 585
R269 B.n648 B.n63 585
R270 B.n647 B.n646 585
R271 B.n645 B.n64 585
R272 B.n644 B.n643 585
R273 B.n642 B.n65 585
R274 B.n641 B.n640 585
R275 B.n639 B.n66 585
R276 B.n638 B.n637 585
R277 B.n636 B.n67 585
R278 B.n635 B.n634 585
R279 B.n633 B.n68 585
R280 B.n632 B.n631 585
R281 B.n630 B.n69 585
R282 B.n629 B.n628 585
R283 B.n627 B.n70 585
R284 B.n626 B.n625 585
R285 B.n624 B.n71 585
R286 B.n623 B.n622 585
R287 B.n621 B.n72 585
R288 B.n620 B.n619 585
R289 B.n618 B.n73 585
R290 B.n617 B.n616 585
R291 B.n615 B.n74 585
R292 B.n614 B.n613 585
R293 B.n612 B.n75 585
R294 B.n611 B.n610 585
R295 B.n609 B.n76 585
R296 B.n608 B.n607 585
R297 B.n606 B.n77 585
R298 B.n605 B.n604 585
R299 B.n603 B.n78 585
R300 B.n602 B.n601 585
R301 B.n600 B.n79 585
R302 B.n599 B.n598 585
R303 B.n597 B.n80 585
R304 B.n596 B.n595 585
R305 B.n594 B.n81 585
R306 B.n593 B.n592 585
R307 B.n591 B.n82 585
R308 B.n590 B.n589 585
R309 B.n588 B.n83 585
R310 B.n750 B.n25 585
R311 B.n752 B.n751 585
R312 B.n753 B.n24 585
R313 B.n755 B.n754 585
R314 B.n756 B.n23 585
R315 B.n758 B.n757 585
R316 B.n759 B.n22 585
R317 B.n761 B.n760 585
R318 B.n762 B.n21 585
R319 B.n764 B.n763 585
R320 B.n765 B.n20 585
R321 B.n767 B.n766 585
R322 B.n768 B.n19 585
R323 B.n770 B.n769 585
R324 B.n771 B.n18 585
R325 B.n773 B.n772 585
R326 B.n774 B.n17 585
R327 B.n776 B.n775 585
R328 B.n777 B.n16 585
R329 B.n779 B.n778 585
R330 B.n780 B.n15 585
R331 B.n782 B.n781 585
R332 B.n783 B.n14 585
R333 B.n785 B.n784 585
R334 B.n786 B.n13 585
R335 B.n788 B.n787 585
R336 B.n789 B.n12 585
R337 B.n791 B.n790 585
R338 B.n792 B.n11 585
R339 B.n794 B.n793 585
R340 B.n795 B.n10 585
R341 B.n797 B.n796 585
R342 B.n798 B.n9 585
R343 B.n800 B.n799 585
R344 B.n801 B.n8 585
R345 B.n803 B.n802 585
R346 B.n804 B.n7 585
R347 B.n806 B.n805 585
R348 B.n807 B.n6 585
R349 B.n809 B.n808 585
R350 B.n810 B.n5 585
R351 B.n812 B.n811 585
R352 B.n813 B.n4 585
R353 B.n815 B.n814 585
R354 B.n816 B.n3 585
R355 B.n818 B.n817 585
R356 B.n819 B.n0 585
R357 B.n2 B.n1 585
R358 B.n213 B.n212 585
R359 B.n215 B.n214 585
R360 B.n216 B.n211 585
R361 B.n218 B.n217 585
R362 B.n219 B.n210 585
R363 B.n221 B.n220 585
R364 B.n222 B.n209 585
R365 B.n224 B.n223 585
R366 B.n225 B.n208 585
R367 B.n227 B.n226 585
R368 B.n228 B.n207 585
R369 B.n230 B.n229 585
R370 B.n231 B.n206 585
R371 B.n233 B.n232 585
R372 B.n234 B.n205 585
R373 B.n236 B.n235 585
R374 B.n237 B.n204 585
R375 B.n239 B.n238 585
R376 B.n240 B.n203 585
R377 B.n242 B.n241 585
R378 B.n243 B.n202 585
R379 B.n245 B.n244 585
R380 B.n246 B.n201 585
R381 B.n248 B.n247 585
R382 B.n249 B.n200 585
R383 B.n251 B.n250 585
R384 B.n252 B.n199 585
R385 B.n254 B.n253 585
R386 B.n255 B.n198 585
R387 B.n257 B.n256 585
R388 B.n258 B.n197 585
R389 B.n260 B.n259 585
R390 B.n261 B.n196 585
R391 B.n263 B.n262 585
R392 B.n264 B.n195 585
R393 B.n266 B.n265 585
R394 B.n267 B.n194 585
R395 B.n269 B.n268 585
R396 B.n270 B.n193 585
R397 B.n272 B.n271 585
R398 B.n273 B.n192 585
R399 B.n275 B.n274 585
R400 B.n276 B.n191 585
R401 B.n278 B.n277 585
R402 B.n279 B.n190 585
R403 B.n281 B.n280 585
R404 B.n280 B.n189 578.989
R405 B.n442 B.n131 578.989
R406 B.n586 B.n83 578.989
R407 B.n748 B.n25 578.989
R408 B.n164 B.t9 323.498
R409 B.n156 B.t0 323.498
R410 B.n58 B.t6 323.498
R411 B.n50 B.t3 323.498
R412 B.n821 B.n820 256.663
R413 B.n820 B.n819 235.042
R414 B.n820 B.n2 235.042
R415 B.n156 B.t1 176.067
R416 B.n58 B.t8 176.067
R417 B.n164 B.t10 176.049
R418 B.n50 B.t5 176.049
R419 B.n284 B.n189 163.367
R420 B.n285 B.n284 163.367
R421 B.n286 B.n285 163.367
R422 B.n286 B.n187 163.367
R423 B.n290 B.n187 163.367
R424 B.n291 B.n290 163.367
R425 B.n292 B.n291 163.367
R426 B.n292 B.n185 163.367
R427 B.n296 B.n185 163.367
R428 B.n297 B.n296 163.367
R429 B.n298 B.n297 163.367
R430 B.n298 B.n183 163.367
R431 B.n302 B.n183 163.367
R432 B.n303 B.n302 163.367
R433 B.n304 B.n303 163.367
R434 B.n304 B.n181 163.367
R435 B.n308 B.n181 163.367
R436 B.n309 B.n308 163.367
R437 B.n310 B.n309 163.367
R438 B.n310 B.n179 163.367
R439 B.n314 B.n179 163.367
R440 B.n315 B.n314 163.367
R441 B.n316 B.n315 163.367
R442 B.n316 B.n177 163.367
R443 B.n320 B.n177 163.367
R444 B.n321 B.n320 163.367
R445 B.n322 B.n321 163.367
R446 B.n322 B.n175 163.367
R447 B.n326 B.n175 163.367
R448 B.n327 B.n326 163.367
R449 B.n328 B.n327 163.367
R450 B.n328 B.n173 163.367
R451 B.n332 B.n173 163.367
R452 B.n333 B.n332 163.367
R453 B.n334 B.n333 163.367
R454 B.n334 B.n171 163.367
R455 B.n338 B.n171 163.367
R456 B.n339 B.n338 163.367
R457 B.n340 B.n339 163.367
R458 B.n340 B.n169 163.367
R459 B.n344 B.n169 163.367
R460 B.n345 B.n344 163.367
R461 B.n346 B.n345 163.367
R462 B.n346 B.n167 163.367
R463 B.n350 B.n167 163.367
R464 B.n351 B.n350 163.367
R465 B.n352 B.n351 163.367
R466 B.n352 B.n163 163.367
R467 B.n357 B.n163 163.367
R468 B.n358 B.n357 163.367
R469 B.n359 B.n358 163.367
R470 B.n359 B.n161 163.367
R471 B.n363 B.n161 163.367
R472 B.n364 B.n363 163.367
R473 B.n365 B.n364 163.367
R474 B.n365 B.n159 163.367
R475 B.n369 B.n159 163.367
R476 B.n370 B.n369 163.367
R477 B.n370 B.n155 163.367
R478 B.n374 B.n155 163.367
R479 B.n375 B.n374 163.367
R480 B.n376 B.n375 163.367
R481 B.n376 B.n153 163.367
R482 B.n380 B.n153 163.367
R483 B.n381 B.n380 163.367
R484 B.n382 B.n381 163.367
R485 B.n382 B.n151 163.367
R486 B.n386 B.n151 163.367
R487 B.n387 B.n386 163.367
R488 B.n388 B.n387 163.367
R489 B.n388 B.n149 163.367
R490 B.n392 B.n149 163.367
R491 B.n393 B.n392 163.367
R492 B.n394 B.n393 163.367
R493 B.n394 B.n147 163.367
R494 B.n398 B.n147 163.367
R495 B.n399 B.n398 163.367
R496 B.n400 B.n399 163.367
R497 B.n400 B.n145 163.367
R498 B.n404 B.n145 163.367
R499 B.n405 B.n404 163.367
R500 B.n406 B.n405 163.367
R501 B.n406 B.n143 163.367
R502 B.n410 B.n143 163.367
R503 B.n411 B.n410 163.367
R504 B.n412 B.n411 163.367
R505 B.n412 B.n141 163.367
R506 B.n416 B.n141 163.367
R507 B.n417 B.n416 163.367
R508 B.n418 B.n417 163.367
R509 B.n418 B.n139 163.367
R510 B.n422 B.n139 163.367
R511 B.n423 B.n422 163.367
R512 B.n424 B.n423 163.367
R513 B.n424 B.n137 163.367
R514 B.n428 B.n137 163.367
R515 B.n429 B.n428 163.367
R516 B.n430 B.n429 163.367
R517 B.n430 B.n135 163.367
R518 B.n434 B.n135 163.367
R519 B.n435 B.n434 163.367
R520 B.n436 B.n435 163.367
R521 B.n436 B.n133 163.367
R522 B.n440 B.n133 163.367
R523 B.n441 B.n440 163.367
R524 B.n442 B.n441 163.367
R525 B.n586 B.n585 163.367
R526 B.n585 B.n584 163.367
R527 B.n584 B.n85 163.367
R528 B.n580 B.n85 163.367
R529 B.n580 B.n579 163.367
R530 B.n579 B.n578 163.367
R531 B.n578 B.n87 163.367
R532 B.n574 B.n87 163.367
R533 B.n574 B.n573 163.367
R534 B.n573 B.n572 163.367
R535 B.n572 B.n89 163.367
R536 B.n568 B.n89 163.367
R537 B.n568 B.n567 163.367
R538 B.n567 B.n566 163.367
R539 B.n566 B.n91 163.367
R540 B.n562 B.n91 163.367
R541 B.n562 B.n561 163.367
R542 B.n561 B.n560 163.367
R543 B.n560 B.n93 163.367
R544 B.n556 B.n93 163.367
R545 B.n556 B.n555 163.367
R546 B.n555 B.n554 163.367
R547 B.n554 B.n95 163.367
R548 B.n550 B.n95 163.367
R549 B.n550 B.n549 163.367
R550 B.n549 B.n548 163.367
R551 B.n548 B.n97 163.367
R552 B.n544 B.n97 163.367
R553 B.n544 B.n543 163.367
R554 B.n543 B.n542 163.367
R555 B.n542 B.n99 163.367
R556 B.n538 B.n99 163.367
R557 B.n538 B.n537 163.367
R558 B.n537 B.n536 163.367
R559 B.n536 B.n101 163.367
R560 B.n532 B.n101 163.367
R561 B.n532 B.n531 163.367
R562 B.n531 B.n530 163.367
R563 B.n530 B.n103 163.367
R564 B.n526 B.n103 163.367
R565 B.n526 B.n525 163.367
R566 B.n525 B.n524 163.367
R567 B.n524 B.n105 163.367
R568 B.n520 B.n105 163.367
R569 B.n520 B.n519 163.367
R570 B.n519 B.n518 163.367
R571 B.n518 B.n107 163.367
R572 B.n514 B.n107 163.367
R573 B.n514 B.n513 163.367
R574 B.n513 B.n512 163.367
R575 B.n512 B.n109 163.367
R576 B.n508 B.n109 163.367
R577 B.n508 B.n507 163.367
R578 B.n507 B.n506 163.367
R579 B.n506 B.n111 163.367
R580 B.n502 B.n111 163.367
R581 B.n502 B.n501 163.367
R582 B.n501 B.n500 163.367
R583 B.n500 B.n113 163.367
R584 B.n496 B.n113 163.367
R585 B.n496 B.n495 163.367
R586 B.n495 B.n494 163.367
R587 B.n494 B.n115 163.367
R588 B.n490 B.n115 163.367
R589 B.n490 B.n489 163.367
R590 B.n489 B.n488 163.367
R591 B.n488 B.n117 163.367
R592 B.n484 B.n117 163.367
R593 B.n484 B.n483 163.367
R594 B.n483 B.n482 163.367
R595 B.n482 B.n119 163.367
R596 B.n478 B.n119 163.367
R597 B.n478 B.n477 163.367
R598 B.n477 B.n476 163.367
R599 B.n476 B.n121 163.367
R600 B.n472 B.n121 163.367
R601 B.n472 B.n471 163.367
R602 B.n471 B.n470 163.367
R603 B.n470 B.n123 163.367
R604 B.n466 B.n123 163.367
R605 B.n466 B.n465 163.367
R606 B.n465 B.n464 163.367
R607 B.n464 B.n125 163.367
R608 B.n460 B.n125 163.367
R609 B.n460 B.n459 163.367
R610 B.n459 B.n458 163.367
R611 B.n458 B.n127 163.367
R612 B.n454 B.n127 163.367
R613 B.n454 B.n453 163.367
R614 B.n453 B.n452 163.367
R615 B.n452 B.n129 163.367
R616 B.n448 B.n129 163.367
R617 B.n448 B.n447 163.367
R618 B.n447 B.n446 163.367
R619 B.n446 B.n131 163.367
R620 B.n748 B.n747 163.367
R621 B.n747 B.n746 163.367
R622 B.n746 B.n27 163.367
R623 B.n742 B.n27 163.367
R624 B.n742 B.n741 163.367
R625 B.n741 B.n740 163.367
R626 B.n740 B.n29 163.367
R627 B.n736 B.n29 163.367
R628 B.n736 B.n735 163.367
R629 B.n735 B.n734 163.367
R630 B.n734 B.n31 163.367
R631 B.n730 B.n31 163.367
R632 B.n730 B.n729 163.367
R633 B.n729 B.n728 163.367
R634 B.n728 B.n33 163.367
R635 B.n724 B.n33 163.367
R636 B.n724 B.n723 163.367
R637 B.n723 B.n722 163.367
R638 B.n722 B.n35 163.367
R639 B.n718 B.n35 163.367
R640 B.n718 B.n717 163.367
R641 B.n717 B.n716 163.367
R642 B.n716 B.n37 163.367
R643 B.n712 B.n37 163.367
R644 B.n712 B.n711 163.367
R645 B.n711 B.n710 163.367
R646 B.n710 B.n39 163.367
R647 B.n706 B.n39 163.367
R648 B.n706 B.n705 163.367
R649 B.n705 B.n704 163.367
R650 B.n704 B.n41 163.367
R651 B.n700 B.n41 163.367
R652 B.n700 B.n699 163.367
R653 B.n699 B.n698 163.367
R654 B.n698 B.n43 163.367
R655 B.n694 B.n43 163.367
R656 B.n694 B.n693 163.367
R657 B.n693 B.n692 163.367
R658 B.n692 B.n45 163.367
R659 B.n688 B.n45 163.367
R660 B.n688 B.n687 163.367
R661 B.n687 B.n686 163.367
R662 B.n686 B.n47 163.367
R663 B.n682 B.n47 163.367
R664 B.n682 B.n681 163.367
R665 B.n681 B.n680 163.367
R666 B.n680 B.n49 163.367
R667 B.n676 B.n49 163.367
R668 B.n676 B.n675 163.367
R669 B.n675 B.n53 163.367
R670 B.n671 B.n53 163.367
R671 B.n671 B.n670 163.367
R672 B.n670 B.n669 163.367
R673 B.n669 B.n55 163.367
R674 B.n665 B.n55 163.367
R675 B.n665 B.n664 163.367
R676 B.n664 B.n663 163.367
R677 B.n663 B.n57 163.367
R678 B.n658 B.n57 163.367
R679 B.n658 B.n657 163.367
R680 B.n657 B.n656 163.367
R681 B.n656 B.n61 163.367
R682 B.n652 B.n61 163.367
R683 B.n652 B.n651 163.367
R684 B.n651 B.n650 163.367
R685 B.n650 B.n63 163.367
R686 B.n646 B.n63 163.367
R687 B.n646 B.n645 163.367
R688 B.n645 B.n644 163.367
R689 B.n644 B.n65 163.367
R690 B.n640 B.n65 163.367
R691 B.n640 B.n639 163.367
R692 B.n639 B.n638 163.367
R693 B.n638 B.n67 163.367
R694 B.n634 B.n67 163.367
R695 B.n634 B.n633 163.367
R696 B.n633 B.n632 163.367
R697 B.n632 B.n69 163.367
R698 B.n628 B.n69 163.367
R699 B.n628 B.n627 163.367
R700 B.n627 B.n626 163.367
R701 B.n626 B.n71 163.367
R702 B.n622 B.n71 163.367
R703 B.n622 B.n621 163.367
R704 B.n621 B.n620 163.367
R705 B.n620 B.n73 163.367
R706 B.n616 B.n73 163.367
R707 B.n616 B.n615 163.367
R708 B.n615 B.n614 163.367
R709 B.n614 B.n75 163.367
R710 B.n610 B.n75 163.367
R711 B.n610 B.n609 163.367
R712 B.n609 B.n608 163.367
R713 B.n608 B.n77 163.367
R714 B.n604 B.n77 163.367
R715 B.n604 B.n603 163.367
R716 B.n603 B.n602 163.367
R717 B.n602 B.n79 163.367
R718 B.n598 B.n79 163.367
R719 B.n598 B.n597 163.367
R720 B.n597 B.n596 163.367
R721 B.n596 B.n81 163.367
R722 B.n592 B.n81 163.367
R723 B.n592 B.n591 163.367
R724 B.n591 B.n590 163.367
R725 B.n590 B.n83 163.367
R726 B.n752 B.n25 163.367
R727 B.n753 B.n752 163.367
R728 B.n754 B.n753 163.367
R729 B.n754 B.n23 163.367
R730 B.n758 B.n23 163.367
R731 B.n759 B.n758 163.367
R732 B.n760 B.n759 163.367
R733 B.n760 B.n21 163.367
R734 B.n764 B.n21 163.367
R735 B.n765 B.n764 163.367
R736 B.n766 B.n765 163.367
R737 B.n766 B.n19 163.367
R738 B.n770 B.n19 163.367
R739 B.n771 B.n770 163.367
R740 B.n772 B.n771 163.367
R741 B.n772 B.n17 163.367
R742 B.n776 B.n17 163.367
R743 B.n777 B.n776 163.367
R744 B.n778 B.n777 163.367
R745 B.n778 B.n15 163.367
R746 B.n782 B.n15 163.367
R747 B.n783 B.n782 163.367
R748 B.n784 B.n783 163.367
R749 B.n784 B.n13 163.367
R750 B.n788 B.n13 163.367
R751 B.n789 B.n788 163.367
R752 B.n790 B.n789 163.367
R753 B.n790 B.n11 163.367
R754 B.n794 B.n11 163.367
R755 B.n795 B.n794 163.367
R756 B.n796 B.n795 163.367
R757 B.n796 B.n9 163.367
R758 B.n800 B.n9 163.367
R759 B.n801 B.n800 163.367
R760 B.n802 B.n801 163.367
R761 B.n802 B.n7 163.367
R762 B.n806 B.n7 163.367
R763 B.n807 B.n806 163.367
R764 B.n808 B.n807 163.367
R765 B.n808 B.n5 163.367
R766 B.n812 B.n5 163.367
R767 B.n813 B.n812 163.367
R768 B.n814 B.n813 163.367
R769 B.n814 B.n3 163.367
R770 B.n818 B.n3 163.367
R771 B.n819 B.n818 163.367
R772 B.n213 B.n2 163.367
R773 B.n214 B.n213 163.367
R774 B.n214 B.n211 163.367
R775 B.n218 B.n211 163.367
R776 B.n219 B.n218 163.367
R777 B.n220 B.n219 163.367
R778 B.n220 B.n209 163.367
R779 B.n224 B.n209 163.367
R780 B.n225 B.n224 163.367
R781 B.n226 B.n225 163.367
R782 B.n226 B.n207 163.367
R783 B.n230 B.n207 163.367
R784 B.n231 B.n230 163.367
R785 B.n232 B.n231 163.367
R786 B.n232 B.n205 163.367
R787 B.n236 B.n205 163.367
R788 B.n237 B.n236 163.367
R789 B.n238 B.n237 163.367
R790 B.n238 B.n203 163.367
R791 B.n242 B.n203 163.367
R792 B.n243 B.n242 163.367
R793 B.n244 B.n243 163.367
R794 B.n244 B.n201 163.367
R795 B.n248 B.n201 163.367
R796 B.n249 B.n248 163.367
R797 B.n250 B.n249 163.367
R798 B.n250 B.n199 163.367
R799 B.n254 B.n199 163.367
R800 B.n255 B.n254 163.367
R801 B.n256 B.n255 163.367
R802 B.n256 B.n197 163.367
R803 B.n260 B.n197 163.367
R804 B.n261 B.n260 163.367
R805 B.n262 B.n261 163.367
R806 B.n262 B.n195 163.367
R807 B.n266 B.n195 163.367
R808 B.n267 B.n266 163.367
R809 B.n268 B.n267 163.367
R810 B.n268 B.n193 163.367
R811 B.n272 B.n193 163.367
R812 B.n273 B.n272 163.367
R813 B.n274 B.n273 163.367
R814 B.n274 B.n191 163.367
R815 B.n278 B.n191 163.367
R816 B.n279 B.n278 163.367
R817 B.n280 B.n279 163.367
R818 B.n157 B.t2 110.71
R819 B.n59 B.t7 110.71
R820 B.n165 B.t11 110.692
R821 B.n51 B.t4 110.692
R822 B.n165 B.n164 65.3581
R823 B.n157 B.n156 65.3581
R824 B.n59 B.n58 65.3581
R825 B.n51 B.n50 65.3581
R826 B.n355 B.n165 59.5399
R827 B.n158 B.n157 59.5399
R828 B.n661 B.n59 59.5399
R829 B.n52 B.n51 59.5399
R830 B.n750 B.n749 37.62
R831 B.n588 B.n587 37.62
R832 B.n444 B.n443 37.62
R833 B.n282 B.n281 37.62
R834 B B.n821 18.0485
R835 B.n751 B.n750 10.6151
R836 B.n751 B.n24 10.6151
R837 B.n755 B.n24 10.6151
R838 B.n756 B.n755 10.6151
R839 B.n757 B.n756 10.6151
R840 B.n757 B.n22 10.6151
R841 B.n761 B.n22 10.6151
R842 B.n762 B.n761 10.6151
R843 B.n763 B.n762 10.6151
R844 B.n763 B.n20 10.6151
R845 B.n767 B.n20 10.6151
R846 B.n768 B.n767 10.6151
R847 B.n769 B.n768 10.6151
R848 B.n769 B.n18 10.6151
R849 B.n773 B.n18 10.6151
R850 B.n774 B.n773 10.6151
R851 B.n775 B.n774 10.6151
R852 B.n775 B.n16 10.6151
R853 B.n779 B.n16 10.6151
R854 B.n780 B.n779 10.6151
R855 B.n781 B.n780 10.6151
R856 B.n781 B.n14 10.6151
R857 B.n785 B.n14 10.6151
R858 B.n786 B.n785 10.6151
R859 B.n787 B.n786 10.6151
R860 B.n787 B.n12 10.6151
R861 B.n791 B.n12 10.6151
R862 B.n792 B.n791 10.6151
R863 B.n793 B.n792 10.6151
R864 B.n793 B.n10 10.6151
R865 B.n797 B.n10 10.6151
R866 B.n798 B.n797 10.6151
R867 B.n799 B.n798 10.6151
R868 B.n799 B.n8 10.6151
R869 B.n803 B.n8 10.6151
R870 B.n804 B.n803 10.6151
R871 B.n805 B.n804 10.6151
R872 B.n805 B.n6 10.6151
R873 B.n809 B.n6 10.6151
R874 B.n810 B.n809 10.6151
R875 B.n811 B.n810 10.6151
R876 B.n811 B.n4 10.6151
R877 B.n815 B.n4 10.6151
R878 B.n816 B.n815 10.6151
R879 B.n817 B.n816 10.6151
R880 B.n817 B.n0 10.6151
R881 B.n749 B.n26 10.6151
R882 B.n745 B.n26 10.6151
R883 B.n745 B.n744 10.6151
R884 B.n744 B.n743 10.6151
R885 B.n743 B.n28 10.6151
R886 B.n739 B.n28 10.6151
R887 B.n739 B.n738 10.6151
R888 B.n738 B.n737 10.6151
R889 B.n737 B.n30 10.6151
R890 B.n733 B.n30 10.6151
R891 B.n733 B.n732 10.6151
R892 B.n732 B.n731 10.6151
R893 B.n731 B.n32 10.6151
R894 B.n727 B.n32 10.6151
R895 B.n727 B.n726 10.6151
R896 B.n726 B.n725 10.6151
R897 B.n725 B.n34 10.6151
R898 B.n721 B.n34 10.6151
R899 B.n721 B.n720 10.6151
R900 B.n720 B.n719 10.6151
R901 B.n719 B.n36 10.6151
R902 B.n715 B.n36 10.6151
R903 B.n715 B.n714 10.6151
R904 B.n714 B.n713 10.6151
R905 B.n713 B.n38 10.6151
R906 B.n709 B.n38 10.6151
R907 B.n709 B.n708 10.6151
R908 B.n708 B.n707 10.6151
R909 B.n707 B.n40 10.6151
R910 B.n703 B.n40 10.6151
R911 B.n703 B.n702 10.6151
R912 B.n702 B.n701 10.6151
R913 B.n701 B.n42 10.6151
R914 B.n697 B.n42 10.6151
R915 B.n697 B.n696 10.6151
R916 B.n696 B.n695 10.6151
R917 B.n695 B.n44 10.6151
R918 B.n691 B.n44 10.6151
R919 B.n691 B.n690 10.6151
R920 B.n690 B.n689 10.6151
R921 B.n689 B.n46 10.6151
R922 B.n685 B.n46 10.6151
R923 B.n685 B.n684 10.6151
R924 B.n684 B.n683 10.6151
R925 B.n683 B.n48 10.6151
R926 B.n679 B.n48 10.6151
R927 B.n679 B.n678 10.6151
R928 B.n678 B.n677 10.6151
R929 B.n674 B.n673 10.6151
R930 B.n673 B.n672 10.6151
R931 B.n672 B.n54 10.6151
R932 B.n668 B.n54 10.6151
R933 B.n668 B.n667 10.6151
R934 B.n667 B.n666 10.6151
R935 B.n666 B.n56 10.6151
R936 B.n662 B.n56 10.6151
R937 B.n660 B.n659 10.6151
R938 B.n659 B.n60 10.6151
R939 B.n655 B.n60 10.6151
R940 B.n655 B.n654 10.6151
R941 B.n654 B.n653 10.6151
R942 B.n653 B.n62 10.6151
R943 B.n649 B.n62 10.6151
R944 B.n649 B.n648 10.6151
R945 B.n648 B.n647 10.6151
R946 B.n647 B.n64 10.6151
R947 B.n643 B.n64 10.6151
R948 B.n643 B.n642 10.6151
R949 B.n642 B.n641 10.6151
R950 B.n641 B.n66 10.6151
R951 B.n637 B.n66 10.6151
R952 B.n637 B.n636 10.6151
R953 B.n636 B.n635 10.6151
R954 B.n635 B.n68 10.6151
R955 B.n631 B.n68 10.6151
R956 B.n631 B.n630 10.6151
R957 B.n630 B.n629 10.6151
R958 B.n629 B.n70 10.6151
R959 B.n625 B.n70 10.6151
R960 B.n625 B.n624 10.6151
R961 B.n624 B.n623 10.6151
R962 B.n623 B.n72 10.6151
R963 B.n619 B.n72 10.6151
R964 B.n619 B.n618 10.6151
R965 B.n618 B.n617 10.6151
R966 B.n617 B.n74 10.6151
R967 B.n613 B.n74 10.6151
R968 B.n613 B.n612 10.6151
R969 B.n612 B.n611 10.6151
R970 B.n611 B.n76 10.6151
R971 B.n607 B.n76 10.6151
R972 B.n607 B.n606 10.6151
R973 B.n606 B.n605 10.6151
R974 B.n605 B.n78 10.6151
R975 B.n601 B.n78 10.6151
R976 B.n601 B.n600 10.6151
R977 B.n600 B.n599 10.6151
R978 B.n599 B.n80 10.6151
R979 B.n595 B.n80 10.6151
R980 B.n595 B.n594 10.6151
R981 B.n594 B.n593 10.6151
R982 B.n593 B.n82 10.6151
R983 B.n589 B.n82 10.6151
R984 B.n589 B.n588 10.6151
R985 B.n587 B.n84 10.6151
R986 B.n583 B.n84 10.6151
R987 B.n583 B.n582 10.6151
R988 B.n582 B.n581 10.6151
R989 B.n581 B.n86 10.6151
R990 B.n577 B.n86 10.6151
R991 B.n577 B.n576 10.6151
R992 B.n576 B.n575 10.6151
R993 B.n575 B.n88 10.6151
R994 B.n571 B.n88 10.6151
R995 B.n571 B.n570 10.6151
R996 B.n570 B.n569 10.6151
R997 B.n569 B.n90 10.6151
R998 B.n565 B.n90 10.6151
R999 B.n565 B.n564 10.6151
R1000 B.n564 B.n563 10.6151
R1001 B.n563 B.n92 10.6151
R1002 B.n559 B.n92 10.6151
R1003 B.n559 B.n558 10.6151
R1004 B.n558 B.n557 10.6151
R1005 B.n557 B.n94 10.6151
R1006 B.n553 B.n94 10.6151
R1007 B.n553 B.n552 10.6151
R1008 B.n552 B.n551 10.6151
R1009 B.n551 B.n96 10.6151
R1010 B.n547 B.n96 10.6151
R1011 B.n547 B.n546 10.6151
R1012 B.n546 B.n545 10.6151
R1013 B.n545 B.n98 10.6151
R1014 B.n541 B.n98 10.6151
R1015 B.n541 B.n540 10.6151
R1016 B.n540 B.n539 10.6151
R1017 B.n539 B.n100 10.6151
R1018 B.n535 B.n100 10.6151
R1019 B.n535 B.n534 10.6151
R1020 B.n534 B.n533 10.6151
R1021 B.n533 B.n102 10.6151
R1022 B.n529 B.n102 10.6151
R1023 B.n529 B.n528 10.6151
R1024 B.n528 B.n527 10.6151
R1025 B.n527 B.n104 10.6151
R1026 B.n523 B.n104 10.6151
R1027 B.n523 B.n522 10.6151
R1028 B.n522 B.n521 10.6151
R1029 B.n521 B.n106 10.6151
R1030 B.n517 B.n106 10.6151
R1031 B.n517 B.n516 10.6151
R1032 B.n516 B.n515 10.6151
R1033 B.n515 B.n108 10.6151
R1034 B.n511 B.n108 10.6151
R1035 B.n511 B.n510 10.6151
R1036 B.n510 B.n509 10.6151
R1037 B.n509 B.n110 10.6151
R1038 B.n505 B.n110 10.6151
R1039 B.n505 B.n504 10.6151
R1040 B.n504 B.n503 10.6151
R1041 B.n503 B.n112 10.6151
R1042 B.n499 B.n112 10.6151
R1043 B.n499 B.n498 10.6151
R1044 B.n498 B.n497 10.6151
R1045 B.n497 B.n114 10.6151
R1046 B.n493 B.n114 10.6151
R1047 B.n493 B.n492 10.6151
R1048 B.n492 B.n491 10.6151
R1049 B.n491 B.n116 10.6151
R1050 B.n487 B.n116 10.6151
R1051 B.n487 B.n486 10.6151
R1052 B.n486 B.n485 10.6151
R1053 B.n485 B.n118 10.6151
R1054 B.n481 B.n118 10.6151
R1055 B.n481 B.n480 10.6151
R1056 B.n480 B.n479 10.6151
R1057 B.n479 B.n120 10.6151
R1058 B.n475 B.n120 10.6151
R1059 B.n475 B.n474 10.6151
R1060 B.n474 B.n473 10.6151
R1061 B.n473 B.n122 10.6151
R1062 B.n469 B.n122 10.6151
R1063 B.n469 B.n468 10.6151
R1064 B.n468 B.n467 10.6151
R1065 B.n467 B.n124 10.6151
R1066 B.n463 B.n124 10.6151
R1067 B.n463 B.n462 10.6151
R1068 B.n462 B.n461 10.6151
R1069 B.n461 B.n126 10.6151
R1070 B.n457 B.n126 10.6151
R1071 B.n457 B.n456 10.6151
R1072 B.n456 B.n455 10.6151
R1073 B.n455 B.n128 10.6151
R1074 B.n451 B.n128 10.6151
R1075 B.n451 B.n450 10.6151
R1076 B.n450 B.n449 10.6151
R1077 B.n449 B.n130 10.6151
R1078 B.n445 B.n130 10.6151
R1079 B.n445 B.n444 10.6151
R1080 B.n212 B.n1 10.6151
R1081 B.n215 B.n212 10.6151
R1082 B.n216 B.n215 10.6151
R1083 B.n217 B.n216 10.6151
R1084 B.n217 B.n210 10.6151
R1085 B.n221 B.n210 10.6151
R1086 B.n222 B.n221 10.6151
R1087 B.n223 B.n222 10.6151
R1088 B.n223 B.n208 10.6151
R1089 B.n227 B.n208 10.6151
R1090 B.n228 B.n227 10.6151
R1091 B.n229 B.n228 10.6151
R1092 B.n229 B.n206 10.6151
R1093 B.n233 B.n206 10.6151
R1094 B.n234 B.n233 10.6151
R1095 B.n235 B.n234 10.6151
R1096 B.n235 B.n204 10.6151
R1097 B.n239 B.n204 10.6151
R1098 B.n240 B.n239 10.6151
R1099 B.n241 B.n240 10.6151
R1100 B.n241 B.n202 10.6151
R1101 B.n245 B.n202 10.6151
R1102 B.n246 B.n245 10.6151
R1103 B.n247 B.n246 10.6151
R1104 B.n247 B.n200 10.6151
R1105 B.n251 B.n200 10.6151
R1106 B.n252 B.n251 10.6151
R1107 B.n253 B.n252 10.6151
R1108 B.n253 B.n198 10.6151
R1109 B.n257 B.n198 10.6151
R1110 B.n258 B.n257 10.6151
R1111 B.n259 B.n258 10.6151
R1112 B.n259 B.n196 10.6151
R1113 B.n263 B.n196 10.6151
R1114 B.n264 B.n263 10.6151
R1115 B.n265 B.n264 10.6151
R1116 B.n265 B.n194 10.6151
R1117 B.n269 B.n194 10.6151
R1118 B.n270 B.n269 10.6151
R1119 B.n271 B.n270 10.6151
R1120 B.n271 B.n192 10.6151
R1121 B.n275 B.n192 10.6151
R1122 B.n276 B.n275 10.6151
R1123 B.n277 B.n276 10.6151
R1124 B.n277 B.n190 10.6151
R1125 B.n281 B.n190 10.6151
R1126 B.n283 B.n282 10.6151
R1127 B.n283 B.n188 10.6151
R1128 B.n287 B.n188 10.6151
R1129 B.n288 B.n287 10.6151
R1130 B.n289 B.n288 10.6151
R1131 B.n289 B.n186 10.6151
R1132 B.n293 B.n186 10.6151
R1133 B.n294 B.n293 10.6151
R1134 B.n295 B.n294 10.6151
R1135 B.n295 B.n184 10.6151
R1136 B.n299 B.n184 10.6151
R1137 B.n300 B.n299 10.6151
R1138 B.n301 B.n300 10.6151
R1139 B.n301 B.n182 10.6151
R1140 B.n305 B.n182 10.6151
R1141 B.n306 B.n305 10.6151
R1142 B.n307 B.n306 10.6151
R1143 B.n307 B.n180 10.6151
R1144 B.n311 B.n180 10.6151
R1145 B.n312 B.n311 10.6151
R1146 B.n313 B.n312 10.6151
R1147 B.n313 B.n178 10.6151
R1148 B.n317 B.n178 10.6151
R1149 B.n318 B.n317 10.6151
R1150 B.n319 B.n318 10.6151
R1151 B.n319 B.n176 10.6151
R1152 B.n323 B.n176 10.6151
R1153 B.n324 B.n323 10.6151
R1154 B.n325 B.n324 10.6151
R1155 B.n325 B.n174 10.6151
R1156 B.n329 B.n174 10.6151
R1157 B.n330 B.n329 10.6151
R1158 B.n331 B.n330 10.6151
R1159 B.n331 B.n172 10.6151
R1160 B.n335 B.n172 10.6151
R1161 B.n336 B.n335 10.6151
R1162 B.n337 B.n336 10.6151
R1163 B.n337 B.n170 10.6151
R1164 B.n341 B.n170 10.6151
R1165 B.n342 B.n341 10.6151
R1166 B.n343 B.n342 10.6151
R1167 B.n343 B.n168 10.6151
R1168 B.n347 B.n168 10.6151
R1169 B.n348 B.n347 10.6151
R1170 B.n349 B.n348 10.6151
R1171 B.n349 B.n166 10.6151
R1172 B.n353 B.n166 10.6151
R1173 B.n354 B.n353 10.6151
R1174 B.n356 B.n162 10.6151
R1175 B.n360 B.n162 10.6151
R1176 B.n361 B.n360 10.6151
R1177 B.n362 B.n361 10.6151
R1178 B.n362 B.n160 10.6151
R1179 B.n366 B.n160 10.6151
R1180 B.n367 B.n366 10.6151
R1181 B.n368 B.n367 10.6151
R1182 B.n372 B.n371 10.6151
R1183 B.n373 B.n372 10.6151
R1184 B.n373 B.n154 10.6151
R1185 B.n377 B.n154 10.6151
R1186 B.n378 B.n377 10.6151
R1187 B.n379 B.n378 10.6151
R1188 B.n379 B.n152 10.6151
R1189 B.n383 B.n152 10.6151
R1190 B.n384 B.n383 10.6151
R1191 B.n385 B.n384 10.6151
R1192 B.n385 B.n150 10.6151
R1193 B.n389 B.n150 10.6151
R1194 B.n390 B.n389 10.6151
R1195 B.n391 B.n390 10.6151
R1196 B.n391 B.n148 10.6151
R1197 B.n395 B.n148 10.6151
R1198 B.n396 B.n395 10.6151
R1199 B.n397 B.n396 10.6151
R1200 B.n397 B.n146 10.6151
R1201 B.n401 B.n146 10.6151
R1202 B.n402 B.n401 10.6151
R1203 B.n403 B.n402 10.6151
R1204 B.n403 B.n144 10.6151
R1205 B.n407 B.n144 10.6151
R1206 B.n408 B.n407 10.6151
R1207 B.n409 B.n408 10.6151
R1208 B.n409 B.n142 10.6151
R1209 B.n413 B.n142 10.6151
R1210 B.n414 B.n413 10.6151
R1211 B.n415 B.n414 10.6151
R1212 B.n415 B.n140 10.6151
R1213 B.n419 B.n140 10.6151
R1214 B.n420 B.n419 10.6151
R1215 B.n421 B.n420 10.6151
R1216 B.n421 B.n138 10.6151
R1217 B.n425 B.n138 10.6151
R1218 B.n426 B.n425 10.6151
R1219 B.n427 B.n426 10.6151
R1220 B.n427 B.n136 10.6151
R1221 B.n431 B.n136 10.6151
R1222 B.n432 B.n431 10.6151
R1223 B.n433 B.n432 10.6151
R1224 B.n433 B.n134 10.6151
R1225 B.n437 B.n134 10.6151
R1226 B.n438 B.n437 10.6151
R1227 B.n439 B.n438 10.6151
R1228 B.n439 B.n132 10.6151
R1229 B.n443 B.n132 10.6151
R1230 B.n821 B.n0 8.11757
R1231 B.n821 B.n1 8.11757
R1232 B.n674 B.n52 6.5566
R1233 B.n662 B.n661 6.5566
R1234 B.n356 B.n355 6.5566
R1235 B.n368 B.n158 6.5566
R1236 B.n677 B.n52 4.05904
R1237 B.n661 B.n660 4.05904
R1238 B.n355 B.n354 4.05904
R1239 B.n371 B.n158 4.05904
R1240 VP.n13 VP.n10 161.3
R1241 VP.n15 VP.n14 161.3
R1242 VP.n16 VP.n9 161.3
R1243 VP.n18 VP.n17 161.3
R1244 VP.n19 VP.n8 161.3
R1245 VP.n21 VP.n20 161.3
R1246 VP.n44 VP.n43 161.3
R1247 VP.n42 VP.n1 161.3
R1248 VP.n41 VP.n40 161.3
R1249 VP.n39 VP.n2 161.3
R1250 VP.n38 VP.n37 161.3
R1251 VP.n36 VP.n3 161.3
R1252 VP.n35 VP.n34 161.3
R1253 VP.n33 VP.n4 161.3
R1254 VP.n32 VP.n31 161.3
R1255 VP.n30 VP.n5 161.3
R1256 VP.n29 VP.n28 161.3
R1257 VP.n27 VP.n6 161.3
R1258 VP.n26 VP.n25 161.3
R1259 VP.n11 VP.t5 148.206
R1260 VP.n35 VP.t2 114.871
R1261 VP.n24 VP.t4 114.871
R1262 VP.n0 VP.t3 114.871
R1263 VP.n12 VP.t1 114.871
R1264 VP.n7 VP.t0 114.871
R1265 VP.n24 VP.n23 71.9618
R1266 VP.n45 VP.n0 71.9618
R1267 VP.n22 VP.n7 71.9618
R1268 VP.n30 VP.n29 56.5193
R1269 VP.n41 VP.n2 56.5193
R1270 VP.n18 VP.n9 56.5193
R1271 VP.n23 VP.n22 52.3895
R1272 VP.n12 VP.n11 49.3079
R1273 VP.n25 VP.n6 24.4675
R1274 VP.n29 VP.n6 24.4675
R1275 VP.n31 VP.n30 24.4675
R1276 VP.n31 VP.n4 24.4675
R1277 VP.n35 VP.n4 24.4675
R1278 VP.n36 VP.n35 24.4675
R1279 VP.n37 VP.n36 24.4675
R1280 VP.n37 VP.n2 24.4675
R1281 VP.n42 VP.n41 24.4675
R1282 VP.n43 VP.n42 24.4675
R1283 VP.n19 VP.n18 24.4675
R1284 VP.n20 VP.n19 24.4675
R1285 VP.n13 VP.n12 24.4675
R1286 VP.n14 VP.n13 24.4675
R1287 VP.n14 VP.n9 24.4675
R1288 VP.n25 VP.n24 18.1061
R1289 VP.n43 VP.n0 18.1061
R1290 VP.n20 VP.n7 18.1061
R1291 VP.n11 VP.n10 4.00589
R1292 VP.n22 VP.n21 0.354971
R1293 VP.n26 VP.n23 0.354971
R1294 VP.n45 VP.n44 0.354971
R1295 VP VP.n45 0.26696
R1296 VP.n15 VP.n10 0.189894
R1297 VP.n16 VP.n15 0.189894
R1298 VP.n17 VP.n16 0.189894
R1299 VP.n17 VP.n8 0.189894
R1300 VP.n21 VP.n8 0.189894
R1301 VP.n27 VP.n26 0.189894
R1302 VP.n28 VP.n27 0.189894
R1303 VP.n28 VP.n5 0.189894
R1304 VP.n32 VP.n5 0.189894
R1305 VP.n33 VP.n32 0.189894
R1306 VP.n34 VP.n33 0.189894
R1307 VP.n34 VP.n3 0.189894
R1308 VP.n38 VP.n3 0.189894
R1309 VP.n39 VP.n38 0.189894
R1310 VP.n40 VP.n39 0.189894
R1311 VP.n40 VP.n1 0.189894
R1312 VP.n44 VP.n1 0.189894
R1313 VTAIL.n7 VTAIL.t4 60.6797
R1314 VTAIL.n11 VTAIL.t2 60.6796
R1315 VTAIL.n2 VTAIL.t9 60.6796
R1316 VTAIL.n10 VTAIL.t8 60.6796
R1317 VTAIL.n9 VTAIL.n8 58.4365
R1318 VTAIL.n6 VTAIL.n5 58.4365
R1319 VTAIL.n1 VTAIL.n0 58.4363
R1320 VTAIL.n4 VTAIL.n3 58.4363
R1321 VTAIL.n6 VTAIL.n4 30.6686
R1322 VTAIL.n11 VTAIL.n10 27.7634
R1323 VTAIL.n7 VTAIL.n6 2.90567
R1324 VTAIL.n10 VTAIL.n9 2.90567
R1325 VTAIL.n4 VTAIL.n2 2.90567
R1326 VTAIL.n0 VTAIL.t1 2.24377
R1327 VTAIL.n0 VTAIL.t5 2.24377
R1328 VTAIL.n3 VTAIL.t11 2.24377
R1329 VTAIL.n3 VTAIL.t7 2.24377
R1330 VTAIL.n8 VTAIL.t10 2.24377
R1331 VTAIL.n8 VTAIL.t6 2.24377
R1332 VTAIL.n5 VTAIL.t0 2.24377
R1333 VTAIL.n5 VTAIL.t3 2.24377
R1334 VTAIL VTAIL.n11 2.12119
R1335 VTAIL.n9 VTAIL.n7 1.92291
R1336 VTAIL.n2 VTAIL.n1 1.92291
R1337 VTAIL VTAIL.n1 0.784983
R1338 VDD1 VDD1.t0 79.5956
R1339 VDD1.n1 VDD1.t1 79.4819
R1340 VDD1.n1 VDD1.n0 75.786
R1341 VDD1.n3 VDD1.n2 75.1151
R1342 VDD1.n3 VDD1.n1 47.6841
R1343 VDD1.n2 VDD1.t4 2.24377
R1344 VDD1.n2 VDD1.t5 2.24377
R1345 VDD1.n0 VDD1.t3 2.24377
R1346 VDD1.n0 VDD1.t2 2.24377
R1347 VDD1 VDD1.n3 0.668603
R1348 VN.n30 VN.n29 161.3
R1349 VN.n28 VN.n17 161.3
R1350 VN.n27 VN.n26 161.3
R1351 VN.n25 VN.n18 161.3
R1352 VN.n24 VN.n23 161.3
R1353 VN.n22 VN.n19 161.3
R1354 VN.n14 VN.n13 161.3
R1355 VN.n12 VN.n1 161.3
R1356 VN.n11 VN.n10 161.3
R1357 VN.n9 VN.n2 161.3
R1358 VN.n8 VN.n7 161.3
R1359 VN.n6 VN.n3 161.3
R1360 VN.n20 VN.t0 148.206
R1361 VN.n4 VN.t3 148.206
R1362 VN.n5 VN.t1 114.871
R1363 VN.n0 VN.t4 114.871
R1364 VN.n21 VN.t2 114.871
R1365 VN.n16 VN.t5 114.871
R1366 VN.n15 VN.n0 71.9618
R1367 VN.n31 VN.n16 71.9618
R1368 VN.n11 VN.n2 56.5193
R1369 VN.n27 VN.n18 56.5193
R1370 VN VN.n31 52.5548
R1371 VN.n5 VN.n4 49.3078
R1372 VN.n21 VN.n20 49.3078
R1373 VN.n6 VN.n5 24.4675
R1374 VN.n7 VN.n6 24.4675
R1375 VN.n7 VN.n2 24.4675
R1376 VN.n12 VN.n11 24.4675
R1377 VN.n13 VN.n12 24.4675
R1378 VN.n23 VN.n18 24.4675
R1379 VN.n23 VN.n22 24.4675
R1380 VN.n22 VN.n21 24.4675
R1381 VN.n29 VN.n28 24.4675
R1382 VN.n28 VN.n27 24.4675
R1383 VN.n13 VN.n0 18.1061
R1384 VN.n29 VN.n16 18.1061
R1385 VN.n20 VN.n19 4.00591
R1386 VN.n4 VN.n3 4.00591
R1387 VN.n31 VN.n30 0.354971
R1388 VN.n15 VN.n14 0.354971
R1389 VN VN.n15 0.26696
R1390 VN.n30 VN.n17 0.189894
R1391 VN.n26 VN.n17 0.189894
R1392 VN.n26 VN.n25 0.189894
R1393 VN.n25 VN.n24 0.189894
R1394 VN.n24 VN.n19 0.189894
R1395 VN.n8 VN.n3 0.189894
R1396 VN.n9 VN.n8 0.189894
R1397 VN.n10 VN.n9 0.189894
R1398 VN.n10 VN.n1 0.189894
R1399 VN.n14 VN.n1 0.189894
R1400 VDD2.n1 VDD2.t2 79.4819
R1401 VDD2.n2 VDD2.t0 77.3585
R1402 VDD2.n1 VDD2.n0 75.786
R1403 VDD2 VDD2.n3 75.7832
R1404 VDD2.n2 VDD2.n1 45.6485
R1405 VDD2.n3 VDD2.t3 2.24377
R1406 VDD2.n3 VDD2.t5 2.24377
R1407 VDD2.n0 VDD2.t4 2.24377
R1408 VDD2.n0 VDD2.t1 2.24377
R1409 VDD2 VDD2.n2 2.23757
C0 w_n3666_n3866# VP 7.57687f
C1 VP VDD2 0.495887f
C2 w_n3666_n3866# B 10.982201f
C3 VP VN 7.81828f
C4 w_n3666_n3866# VDD1 2.5712f
C5 B VDD2 2.49158f
C6 w_n3666_n3866# VTAIL 3.35645f
C7 VDD2 VDD1 1.57943f
C8 VTAIL VDD2 8.74802f
C9 B VN 1.2892f
C10 VN VDD1 0.151428f
C11 VTAIL VN 8.41655f
C12 B VP 2.08479f
C13 VP VDD1 8.60525f
C14 VTAIL VP 8.43083f
C15 w_n3666_n3866# VDD2 2.67032f
C16 B VDD1 2.40693f
C17 w_n3666_n3866# VN 7.10169f
C18 B VTAIL 4.44014f
C19 VTAIL VDD1 8.694309f
C20 VDD2 VN 8.264269f
C21 VDD2 VSUBS 2.074399f
C22 VDD1 VSUBS 2.5962f
C23 VTAIL VSUBS 1.369461f
C24 VN VSUBS 6.3512f
C25 VP VSUBS 3.378192f
C26 B VSUBS 5.28363f
C27 w_n3666_n3866# VSUBS 0.1739p
C28 VDD2.t2 VSUBS 3.37658f
C29 VDD2.t4 VSUBS 0.317495f
C30 VDD2.t1 VSUBS 0.317495f
C31 VDD2.n0 VSUBS 2.58741f
C32 VDD2.n1 VSUBS 4.18323f
C33 VDD2.t0 VSUBS 3.35513f
C34 VDD2.n2 VSUBS 3.74611f
C35 VDD2.t3 VSUBS 0.317495f
C36 VDD2.t5 VSUBS 0.317495f
C37 VDD2.n3 VSUBS 2.58736f
C38 VN.t4 VSUBS 3.19257f
C39 VN.n0 VSUBS 1.21602f
C40 VN.n1 VSUBS 0.026471f
C41 VN.n2 VSUBS 0.03385f
C42 VN.n3 VSUBS 0.301142f
C43 VN.t1 VSUBS 3.19257f
C44 VN.t3 VSUBS 3.4844f
C45 VN.n4 VSUBS 1.15467f
C46 VN.n5 VSUBS 1.2122f
C47 VN.n6 VSUBS 0.049335f
C48 VN.n7 VSUBS 0.049335f
C49 VN.n8 VSUBS 0.026471f
C50 VN.n9 VSUBS 0.026471f
C51 VN.n10 VSUBS 0.026471f
C52 VN.n11 VSUBS 0.043439f
C53 VN.n12 VSUBS 0.049335f
C54 VN.n13 VSUBS 0.043002f
C55 VN.n14 VSUBS 0.042723f
C56 VN.n15 VSUBS 0.057653f
C57 VN.t5 VSUBS 3.19257f
C58 VN.n16 VSUBS 1.21602f
C59 VN.n17 VSUBS 0.026471f
C60 VN.n18 VSUBS 0.03385f
C61 VN.n19 VSUBS 0.301142f
C62 VN.t2 VSUBS 3.19257f
C63 VN.t0 VSUBS 3.4844f
C64 VN.n20 VSUBS 1.15467f
C65 VN.n21 VSUBS 1.2122f
C66 VN.n22 VSUBS 0.049335f
C67 VN.n23 VSUBS 0.049335f
C68 VN.n24 VSUBS 0.026471f
C69 VN.n25 VSUBS 0.026471f
C70 VN.n26 VSUBS 0.026471f
C71 VN.n27 VSUBS 0.043439f
C72 VN.n28 VSUBS 0.049335f
C73 VN.n29 VSUBS 0.043002f
C74 VN.n30 VSUBS 0.042723f
C75 VN.n31 VSUBS 1.61251f
C76 VDD1.t0 VSUBS 3.37763f
C77 VDD1.t1 VSUBS 3.37622f
C78 VDD1.t3 VSUBS 0.317461f
C79 VDD1.t2 VSUBS 0.317461f
C80 VDD1.n0 VSUBS 2.58713f
C81 VDD1.n1 VSUBS 4.33545f
C82 VDD1.t4 VSUBS 0.317461f
C83 VDD1.t5 VSUBS 0.317461f
C84 VDD1.n2 VSUBS 2.57966f
C85 VDD1.n3 VSUBS 3.72411f
C86 VTAIL.t1 VSUBS 0.327425f
C87 VTAIL.t5 VSUBS 0.327425f
C88 VTAIL.n0 VSUBS 2.51159f
C89 VTAIL.n1 VSUBS 0.887215f
C90 VTAIL.t9 VSUBS 3.29079f
C91 VTAIL.n2 VSUBS 1.19638f
C92 VTAIL.t11 VSUBS 0.327425f
C93 VTAIL.t7 VSUBS 0.327425f
C94 VTAIL.n3 VSUBS 2.51159f
C95 VTAIL.n4 VSUBS 2.98022f
C96 VTAIL.t0 VSUBS 0.327425f
C97 VTAIL.t3 VSUBS 0.327425f
C98 VTAIL.n5 VSUBS 2.51159f
C99 VTAIL.n6 VSUBS 2.98022f
C100 VTAIL.t4 VSUBS 3.29082f
C101 VTAIL.n7 VSUBS 1.19636f
C102 VTAIL.t10 VSUBS 0.327425f
C103 VTAIL.t6 VSUBS 0.327425f
C104 VTAIL.n8 VSUBS 2.51159f
C105 VTAIL.n9 VSUBS 1.08261f
C106 VTAIL.t8 VSUBS 3.2908f
C107 VTAIL.n10 VSUBS 2.82631f
C108 VTAIL.t2 VSUBS 3.29079f
C109 VTAIL.n11 VSUBS 2.75403f
C110 VP.t3 VSUBS 3.48966f
C111 VP.n0 VSUBS 1.32918f
C112 VP.n1 VSUBS 0.028934f
C113 VP.n2 VSUBS 0.037f
C114 VP.n3 VSUBS 0.028934f
C115 VP.t2 VSUBS 3.48966f
C116 VP.n4 VSUBS 0.053926f
C117 VP.n5 VSUBS 0.028934f
C118 VP.n6 VSUBS 0.053926f
C119 VP.t0 VSUBS 3.48966f
C120 VP.n7 VSUBS 1.32918f
C121 VP.n8 VSUBS 0.028934f
C122 VP.n9 VSUBS 0.037f
C123 VP.n10 VSUBS 0.329166f
C124 VP.t1 VSUBS 3.48966f
C125 VP.t5 VSUBS 3.80865f
C126 VP.n11 VSUBS 1.26212f
C127 VP.n12 VSUBS 1.32501f
C128 VP.n13 VSUBS 0.053926f
C129 VP.n14 VSUBS 0.053926f
C130 VP.n15 VSUBS 0.028934f
C131 VP.n16 VSUBS 0.028934f
C132 VP.n17 VSUBS 0.028934f
C133 VP.n18 VSUBS 0.047482f
C134 VP.n19 VSUBS 0.053926f
C135 VP.n20 VSUBS 0.047004f
C136 VP.n21 VSUBS 0.046699f
C137 VP.n22 VSUBS 1.75091f
C138 VP.n23 VSUBS 1.77077f
C139 VP.t4 VSUBS 3.48966f
C140 VP.n24 VSUBS 1.32918f
C141 VP.n25 VSUBS 0.047004f
C142 VP.n26 VSUBS 0.046699f
C143 VP.n27 VSUBS 0.028934f
C144 VP.n28 VSUBS 0.028934f
C145 VP.n29 VSUBS 0.047482f
C146 VP.n30 VSUBS 0.037f
C147 VP.n31 VSUBS 0.053926f
C148 VP.n32 VSUBS 0.028934f
C149 VP.n33 VSUBS 0.028934f
C150 VP.n34 VSUBS 0.028934f
C151 VP.n35 VSUBS 1.24454f
C152 VP.n36 VSUBS 0.053926f
C153 VP.n37 VSUBS 0.053926f
C154 VP.n38 VSUBS 0.028934f
C155 VP.n39 VSUBS 0.028934f
C156 VP.n40 VSUBS 0.028934f
C157 VP.n41 VSUBS 0.047482f
C158 VP.n42 VSUBS 0.053926f
C159 VP.n43 VSUBS 0.047004f
C160 VP.n44 VSUBS 0.046699f
C161 VP.n45 VSUBS 0.063018f
C162 B.n0 VSUBS 0.007168f
C163 B.n1 VSUBS 0.007168f
C164 B.n2 VSUBS 0.0106f
C165 B.n3 VSUBS 0.008123f
C166 B.n4 VSUBS 0.008123f
C167 B.n5 VSUBS 0.008123f
C168 B.n6 VSUBS 0.008123f
C169 B.n7 VSUBS 0.008123f
C170 B.n8 VSUBS 0.008123f
C171 B.n9 VSUBS 0.008123f
C172 B.n10 VSUBS 0.008123f
C173 B.n11 VSUBS 0.008123f
C174 B.n12 VSUBS 0.008123f
C175 B.n13 VSUBS 0.008123f
C176 B.n14 VSUBS 0.008123f
C177 B.n15 VSUBS 0.008123f
C178 B.n16 VSUBS 0.008123f
C179 B.n17 VSUBS 0.008123f
C180 B.n18 VSUBS 0.008123f
C181 B.n19 VSUBS 0.008123f
C182 B.n20 VSUBS 0.008123f
C183 B.n21 VSUBS 0.008123f
C184 B.n22 VSUBS 0.008123f
C185 B.n23 VSUBS 0.008123f
C186 B.n24 VSUBS 0.008123f
C187 B.n25 VSUBS 0.020489f
C188 B.n26 VSUBS 0.008123f
C189 B.n27 VSUBS 0.008123f
C190 B.n28 VSUBS 0.008123f
C191 B.n29 VSUBS 0.008123f
C192 B.n30 VSUBS 0.008123f
C193 B.n31 VSUBS 0.008123f
C194 B.n32 VSUBS 0.008123f
C195 B.n33 VSUBS 0.008123f
C196 B.n34 VSUBS 0.008123f
C197 B.n35 VSUBS 0.008123f
C198 B.n36 VSUBS 0.008123f
C199 B.n37 VSUBS 0.008123f
C200 B.n38 VSUBS 0.008123f
C201 B.n39 VSUBS 0.008123f
C202 B.n40 VSUBS 0.008123f
C203 B.n41 VSUBS 0.008123f
C204 B.n42 VSUBS 0.008123f
C205 B.n43 VSUBS 0.008123f
C206 B.n44 VSUBS 0.008123f
C207 B.n45 VSUBS 0.008123f
C208 B.n46 VSUBS 0.008123f
C209 B.n47 VSUBS 0.008123f
C210 B.n48 VSUBS 0.008123f
C211 B.n49 VSUBS 0.008123f
C212 B.t4 VSUBS 0.558114f
C213 B.t5 VSUBS 0.585591f
C214 B.t3 VSUBS 2.32572f
C215 B.n50 VSUBS 0.326441f
C216 B.n51 VSUBS 0.085598f
C217 B.n52 VSUBS 0.018821f
C218 B.n53 VSUBS 0.008123f
C219 B.n54 VSUBS 0.008123f
C220 B.n55 VSUBS 0.008123f
C221 B.n56 VSUBS 0.008123f
C222 B.n57 VSUBS 0.008123f
C223 B.t7 VSUBS 0.558099f
C224 B.t8 VSUBS 0.585579f
C225 B.t6 VSUBS 2.32572f
C226 B.n58 VSUBS 0.326453f
C227 B.n59 VSUBS 0.085613f
C228 B.n60 VSUBS 0.008123f
C229 B.n61 VSUBS 0.008123f
C230 B.n62 VSUBS 0.008123f
C231 B.n63 VSUBS 0.008123f
C232 B.n64 VSUBS 0.008123f
C233 B.n65 VSUBS 0.008123f
C234 B.n66 VSUBS 0.008123f
C235 B.n67 VSUBS 0.008123f
C236 B.n68 VSUBS 0.008123f
C237 B.n69 VSUBS 0.008123f
C238 B.n70 VSUBS 0.008123f
C239 B.n71 VSUBS 0.008123f
C240 B.n72 VSUBS 0.008123f
C241 B.n73 VSUBS 0.008123f
C242 B.n74 VSUBS 0.008123f
C243 B.n75 VSUBS 0.008123f
C244 B.n76 VSUBS 0.008123f
C245 B.n77 VSUBS 0.008123f
C246 B.n78 VSUBS 0.008123f
C247 B.n79 VSUBS 0.008123f
C248 B.n80 VSUBS 0.008123f
C249 B.n81 VSUBS 0.008123f
C250 B.n82 VSUBS 0.008123f
C251 B.n83 VSUBS 0.021322f
C252 B.n84 VSUBS 0.008123f
C253 B.n85 VSUBS 0.008123f
C254 B.n86 VSUBS 0.008123f
C255 B.n87 VSUBS 0.008123f
C256 B.n88 VSUBS 0.008123f
C257 B.n89 VSUBS 0.008123f
C258 B.n90 VSUBS 0.008123f
C259 B.n91 VSUBS 0.008123f
C260 B.n92 VSUBS 0.008123f
C261 B.n93 VSUBS 0.008123f
C262 B.n94 VSUBS 0.008123f
C263 B.n95 VSUBS 0.008123f
C264 B.n96 VSUBS 0.008123f
C265 B.n97 VSUBS 0.008123f
C266 B.n98 VSUBS 0.008123f
C267 B.n99 VSUBS 0.008123f
C268 B.n100 VSUBS 0.008123f
C269 B.n101 VSUBS 0.008123f
C270 B.n102 VSUBS 0.008123f
C271 B.n103 VSUBS 0.008123f
C272 B.n104 VSUBS 0.008123f
C273 B.n105 VSUBS 0.008123f
C274 B.n106 VSUBS 0.008123f
C275 B.n107 VSUBS 0.008123f
C276 B.n108 VSUBS 0.008123f
C277 B.n109 VSUBS 0.008123f
C278 B.n110 VSUBS 0.008123f
C279 B.n111 VSUBS 0.008123f
C280 B.n112 VSUBS 0.008123f
C281 B.n113 VSUBS 0.008123f
C282 B.n114 VSUBS 0.008123f
C283 B.n115 VSUBS 0.008123f
C284 B.n116 VSUBS 0.008123f
C285 B.n117 VSUBS 0.008123f
C286 B.n118 VSUBS 0.008123f
C287 B.n119 VSUBS 0.008123f
C288 B.n120 VSUBS 0.008123f
C289 B.n121 VSUBS 0.008123f
C290 B.n122 VSUBS 0.008123f
C291 B.n123 VSUBS 0.008123f
C292 B.n124 VSUBS 0.008123f
C293 B.n125 VSUBS 0.008123f
C294 B.n126 VSUBS 0.008123f
C295 B.n127 VSUBS 0.008123f
C296 B.n128 VSUBS 0.008123f
C297 B.n129 VSUBS 0.008123f
C298 B.n130 VSUBS 0.008123f
C299 B.n131 VSUBS 0.020489f
C300 B.n132 VSUBS 0.008123f
C301 B.n133 VSUBS 0.008123f
C302 B.n134 VSUBS 0.008123f
C303 B.n135 VSUBS 0.008123f
C304 B.n136 VSUBS 0.008123f
C305 B.n137 VSUBS 0.008123f
C306 B.n138 VSUBS 0.008123f
C307 B.n139 VSUBS 0.008123f
C308 B.n140 VSUBS 0.008123f
C309 B.n141 VSUBS 0.008123f
C310 B.n142 VSUBS 0.008123f
C311 B.n143 VSUBS 0.008123f
C312 B.n144 VSUBS 0.008123f
C313 B.n145 VSUBS 0.008123f
C314 B.n146 VSUBS 0.008123f
C315 B.n147 VSUBS 0.008123f
C316 B.n148 VSUBS 0.008123f
C317 B.n149 VSUBS 0.008123f
C318 B.n150 VSUBS 0.008123f
C319 B.n151 VSUBS 0.008123f
C320 B.n152 VSUBS 0.008123f
C321 B.n153 VSUBS 0.008123f
C322 B.n154 VSUBS 0.008123f
C323 B.n155 VSUBS 0.008123f
C324 B.t2 VSUBS 0.558099f
C325 B.t1 VSUBS 0.585579f
C326 B.t0 VSUBS 2.32572f
C327 B.n156 VSUBS 0.326453f
C328 B.n157 VSUBS 0.085613f
C329 B.n158 VSUBS 0.018821f
C330 B.n159 VSUBS 0.008123f
C331 B.n160 VSUBS 0.008123f
C332 B.n161 VSUBS 0.008123f
C333 B.n162 VSUBS 0.008123f
C334 B.n163 VSUBS 0.008123f
C335 B.t11 VSUBS 0.558114f
C336 B.t10 VSUBS 0.585591f
C337 B.t9 VSUBS 2.32572f
C338 B.n164 VSUBS 0.326441f
C339 B.n165 VSUBS 0.085598f
C340 B.n166 VSUBS 0.008123f
C341 B.n167 VSUBS 0.008123f
C342 B.n168 VSUBS 0.008123f
C343 B.n169 VSUBS 0.008123f
C344 B.n170 VSUBS 0.008123f
C345 B.n171 VSUBS 0.008123f
C346 B.n172 VSUBS 0.008123f
C347 B.n173 VSUBS 0.008123f
C348 B.n174 VSUBS 0.008123f
C349 B.n175 VSUBS 0.008123f
C350 B.n176 VSUBS 0.008123f
C351 B.n177 VSUBS 0.008123f
C352 B.n178 VSUBS 0.008123f
C353 B.n179 VSUBS 0.008123f
C354 B.n180 VSUBS 0.008123f
C355 B.n181 VSUBS 0.008123f
C356 B.n182 VSUBS 0.008123f
C357 B.n183 VSUBS 0.008123f
C358 B.n184 VSUBS 0.008123f
C359 B.n185 VSUBS 0.008123f
C360 B.n186 VSUBS 0.008123f
C361 B.n187 VSUBS 0.008123f
C362 B.n188 VSUBS 0.008123f
C363 B.n189 VSUBS 0.021322f
C364 B.n190 VSUBS 0.008123f
C365 B.n191 VSUBS 0.008123f
C366 B.n192 VSUBS 0.008123f
C367 B.n193 VSUBS 0.008123f
C368 B.n194 VSUBS 0.008123f
C369 B.n195 VSUBS 0.008123f
C370 B.n196 VSUBS 0.008123f
C371 B.n197 VSUBS 0.008123f
C372 B.n198 VSUBS 0.008123f
C373 B.n199 VSUBS 0.008123f
C374 B.n200 VSUBS 0.008123f
C375 B.n201 VSUBS 0.008123f
C376 B.n202 VSUBS 0.008123f
C377 B.n203 VSUBS 0.008123f
C378 B.n204 VSUBS 0.008123f
C379 B.n205 VSUBS 0.008123f
C380 B.n206 VSUBS 0.008123f
C381 B.n207 VSUBS 0.008123f
C382 B.n208 VSUBS 0.008123f
C383 B.n209 VSUBS 0.008123f
C384 B.n210 VSUBS 0.008123f
C385 B.n211 VSUBS 0.008123f
C386 B.n212 VSUBS 0.008123f
C387 B.n213 VSUBS 0.008123f
C388 B.n214 VSUBS 0.008123f
C389 B.n215 VSUBS 0.008123f
C390 B.n216 VSUBS 0.008123f
C391 B.n217 VSUBS 0.008123f
C392 B.n218 VSUBS 0.008123f
C393 B.n219 VSUBS 0.008123f
C394 B.n220 VSUBS 0.008123f
C395 B.n221 VSUBS 0.008123f
C396 B.n222 VSUBS 0.008123f
C397 B.n223 VSUBS 0.008123f
C398 B.n224 VSUBS 0.008123f
C399 B.n225 VSUBS 0.008123f
C400 B.n226 VSUBS 0.008123f
C401 B.n227 VSUBS 0.008123f
C402 B.n228 VSUBS 0.008123f
C403 B.n229 VSUBS 0.008123f
C404 B.n230 VSUBS 0.008123f
C405 B.n231 VSUBS 0.008123f
C406 B.n232 VSUBS 0.008123f
C407 B.n233 VSUBS 0.008123f
C408 B.n234 VSUBS 0.008123f
C409 B.n235 VSUBS 0.008123f
C410 B.n236 VSUBS 0.008123f
C411 B.n237 VSUBS 0.008123f
C412 B.n238 VSUBS 0.008123f
C413 B.n239 VSUBS 0.008123f
C414 B.n240 VSUBS 0.008123f
C415 B.n241 VSUBS 0.008123f
C416 B.n242 VSUBS 0.008123f
C417 B.n243 VSUBS 0.008123f
C418 B.n244 VSUBS 0.008123f
C419 B.n245 VSUBS 0.008123f
C420 B.n246 VSUBS 0.008123f
C421 B.n247 VSUBS 0.008123f
C422 B.n248 VSUBS 0.008123f
C423 B.n249 VSUBS 0.008123f
C424 B.n250 VSUBS 0.008123f
C425 B.n251 VSUBS 0.008123f
C426 B.n252 VSUBS 0.008123f
C427 B.n253 VSUBS 0.008123f
C428 B.n254 VSUBS 0.008123f
C429 B.n255 VSUBS 0.008123f
C430 B.n256 VSUBS 0.008123f
C431 B.n257 VSUBS 0.008123f
C432 B.n258 VSUBS 0.008123f
C433 B.n259 VSUBS 0.008123f
C434 B.n260 VSUBS 0.008123f
C435 B.n261 VSUBS 0.008123f
C436 B.n262 VSUBS 0.008123f
C437 B.n263 VSUBS 0.008123f
C438 B.n264 VSUBS 0.008123f
C439 B.n265 VSUBS 0.008123f
C440 B.n266 VSUBS 0.008123f
C441 B.n267 VSUBS 0.008123f
C442 B.n268 VSUBS 0.008123f
C443 B.n269 VSUBS 0.008123f
C444 B.n270 VSUBS 0.008123f
C445 B.n271 VSUBS 0.008123f
C446 B.n272 VSUBS 0.008123f
C447 B.n273 VSUBS 0.008123f
C448 B.n274 VSUBS 0.008123f
C449 B.n275 VSUBS 0.008123f
C450 B.n276 VSUBS 0.008123f
C451 B.n277 VSUBS 0.008123f
C452 B.n278 VSUBS 0.008123f
C453 B.n279 VSUBS 0.008123f
C454 B.n280 VSUBS 0.020489f
C455 B.n281 VSUBS 0.020489f
C456 B.n282 VSUBS 0.021322f
C457 B.n283 VSUBS 0.008123f
C458 B.n284 VSUBS 0.008123f
C459 B.n285 VSUBS 0.008123f
C460 B.n286 VSUBS 0.008123f
C461 B.n287 VSUBS 0.008123f
C462 B.n288 VSUBS 0.008123f
C463 B.n289 VSUBS 0.008123f
C464 B.n290 VSUBS 0.008123f
C465 B.n291 VSUBS 0.008123f
C466 B.n292 VSUBS 0.008123f
C467 B.n293 VSUBS 0.008123f
C468 B.n294 VSUBS 0.008123f
C469 B.n295 VSUBS 0.008123f
C470 B.n296 VSUBS 0.008123f
C471 B.n297 VSUBS 0.008123f
C472 B.n298 VSUBS 0.008123f
C473 B.n299 VSUBS 0.008123f
C474 B.n300 VSUBS 0.008123f
C475 B.n301 VSUBS 0.008123f
C476 B.n302 VSUBS 0.008123f
C477 B.n303 VSUBS 0.008123f
C478 B.n304 VSUBS 0.008123f
C479 B.n305 VSUBS 0.008123f
C480 B.n306 VSUBS 0.008123f
C481 B.n307 VSUBS 0.008123f
C482 B.n308 VSUBS 0.008123f
C483 B.n309 VSUBS 0.008123f
C484 B.n310 VSUBS 0.008123f
C485 B.n311 VSUBS 0.008123f
C486 B.n312 VSUBS 0.008123f
C487 B.n313 VSUBS 0.008123f
C488 B.n314 VSUBS 0.008123f
C489 B.n315 VSUBS 0.008123f
C490 B.n316 VSUBS 0.008123f
C491 B.n317 VSUBS 0.008123f
C492 B.n318 VSUBS 0.008123f
C493 B.n319 VSUBS 0.008123f
C494 B.n320 VSUBS 0.008123f
C495 B.n321 VSUBS 0.008123f
C496 B.n322 VSUBS 0.008123f
C497 B.n323 VSUBS 0.008123f
C498 B.n324 VSUBS 0.008123f
C499 B.n325 VSUBS 0.008123f
C500 B.n326 VSUBS 0.008123f
C501 B.n327 VSUBS 0.008123f
C502 B.n328 VSUBS 0.008123f
C503 B.n329 VSUBS 0.008123f
C504 B.n330 VSUBS 0.008123f
C505 B.n331 VSUBS 0.008123f
C506 B.n332 VSUBS 0.008123f
C507 B.n333 VSUBS 0.008123f
C508 B.n334 VSUBS 0.008123f
C509 B.n335 VSUBS 0.008123f
C510 B.n336 VSUBS 0.008123f
C511 B.n337 VSUBS 0.008123f
C512 B.n338 VSUBS 0.008123f
C513 B.n339 VSUBS 0.008123f
C514 B.n340 VSUBS 0.008123f
C515 B.n341 VSUBS 0.008123f
C516 B.n342 VSUBS 0.008123f
C517 B.n343 VSUBS 0.008123f
C518 B.n344 VSUBS 0.008123f
C519 B.n345 VSUBS 0.008123f
C520 B.n346 VSUBS 0.008123f
C521 B.n347 VSUBS 0.008123f
C522 B.n348 VSUBS 0.008123f
C523 B.n349 VSUBS 0.008123f
C524 B.n350 VSUBS 0.008123f
C525 B.n351 VSUBS 0.008123f
C526 B.n352 VSUBS 0.008123f
C527 B.n353 VSUBS 0.008123f
C528 B.n354 VSUBS 0.005615f
C529 B.n355 VSUBS 0.018821f
C530 B.n356 VSUBS 0.00657f
C531 B.n357 VSUBS 0.008123f
C532 B.n358 VSUBS 0.008123f
C533 B.n359 VSUBS 0.008123f
C534 B.n360 VSUBS 0.008123f
C535 B.n361 VSUBS 0.008123f
C536 B.n362 VSUBS 0.008123f
C537 B.n363 VSUBS 0.008123f
C538 B.n364 VSUBS 0.008123f
C539 B.n365 VSUBS 0.008123f
C540 B.n366 VSUBS 0.008123f
C541 B.n367 VSUBS 0.008123f
C542 B.n368 VSUBS 0.00657f
C543 B.n369 VSUBS 0.008123f
C544 B.n370 VSUBS 0.008123f
C545 B.n371 VSUBS 0.005615f
C546 B.n372 VSUBS 0.008123f
C547 B.n373 VSUBS 0.008123f
C548 B.n374 VSUBS 0.008123f
C549 B.n375 VSUBS 0.008123f
C550 B.n376 VSUBS 0.008123f
C551 B.n377 VSUBS 0.008123f
C552 B.n378 VSUBS 0.008123f
C553 B.n379 VSUBS 0.008123f
C554 B.n380 VSUBS 0.008123f
C555 B.n381 VSUBS 0.008123f
C556 B.n382 VSUBS 0.008123f
C557 B.n383 VSUBS 0.008123f
C558 B.n384 VSUBS 0.008123f
C559 B.n385 VSUBS 0.008123f
C560 B.n386 VSUBS 0.008123f
C561 B.n387 VSUBS 0.008123f
C562 B.n388 VSUBS 0.008123f
C563 B.n389 VSUBS 0.008123f
C564 B.n390 VSUBS 0.008123f
C565 B.n391 VSUBS 0.008123f
C566 B.n392 VSUBS 0.008123f
C567 B.n393 VSUBS 0.008123f
C568 B.n394 VSUBS 0.008123f
C569 B.n395 VSUBS 0.008123f
C570 B.n396 VSUBS 0.008123f
C571 B.n397 VSUBS 0.008123f
C572 B.n398 VSUBS 0.008123f
C573 B.n399 VSUBS 0.008123f
C574 B.n400 VSUBS 0.008123f
C575 B.n401 VSUBS 0.008123f
C576 B.n402 VSUBS 0.008123f
C577 B.n403 VSUBS 0.008123f
C578 B.n404 VSUBS 0.008123f
C579 B.n405 VSUBS 0.008123f
C580 B.n406 VSUBS 0.008123f
C581 B.n407 VSUBS 0.008123f
C582 B.n408 VSUBS 0.008123f
C583 B.n409 VSUBS 0.008123f
C584 B.n410 VSUBS 0.008123f
C585 B.n411 VSUBS 0.008123f
C586 B.n412 VSUBS 0.008123f
C587 B.n413 VSUBS 0.008123f
C588 B.n414 VSUBS 0.008123f
C589 B.n415 VSUBS 0.008123f
C590 B.n416 VSUBS 0.008123f
C591 B.n417 VSUBS 0.008123f
C592 B.n418 VSUBS 0.008123f
C593 B.n419 VSUBS 0.008123f
C594 B.n420 VSUBS 0.008123f
C595 B.n421 VSUBS 0.008123f
C596 B.n422 VSUBS 0.008123f
C597 B.n423 VSUBS 0.008123f
C598 B.n424 VSUBS 0.008123f
C599 B.n425 VSUBS 0.008123f
C600 B.n426 VSUBS 0.008123f
C601 B.n427 VSUBS 0.008123f
C602 B.n428 VSUBS 0.008123f
C603 B.n429 VSUBS 0.008123f
C604 B.n430 VSUBS 0.008123f
C605 B.n431 VSUBS 0.008123f
C606 B.n432 VSUBS 0.008123f
C607 B.n433 VSUBS 0.008123f
C608 B.n434 VSUBS 0.008123f
C609 B.n435 VSUBS 0.008123f
C610 B.n436 VSUBS 0.008123f
C611 B.n437 VSUBS 0.008123f
C612 B.n438 VSUBS 0.008123f
C613 B.n439 VSUBS 0.008123f
C614 B.n440 VSUBS 0.008123f
C615 B.n441 VSUBS 0.008123f
C616 B.n442 VSUBS 0.021322f
C617 B.n443 VSUBS 0.020489f
C618 B.n444 VSUBS 0.021322f
C619 B.n445 VSUBS 0.008123f
C620 B.n446 VSUBS 0.008123f
C621 B.n447 VSUBS 0.008123f
C622 B.n448 VSUBS 0.008123f
C623 B.n449 VSUBS 0.008123f
C624 B.n450 VSUBS 0.008123f
C625 B.n451 VSUBS 0.008123f
C626 B.n452 VSUBS 0.008123f
C627 B.n453 VSUBS 0.008123f
C628 B.n454 VSUBS 0.008123f
C629 B.n455 VSUBS 0.008123f
C630 B.n456 VSUBS 0.008123f
C631 B.n457 VSUBS 0.008123f
C632 B.n458 VSUBS 0.008123f
C633 B.n459 VSUBS 0.008123f
C634 B.n460 VSUBS 0.008123f
C635 B.n461 VSUBS 0.008123f
C636 B.n462 VSUBS 0.008123f
C637 B.n463 VSUBS 0.008123f
C638 B.n464 VSUBS 0.008123f
C639 B.n465 VSUBS 0.008123f
C640 B.n466 VSUBS 0.008123f
C641 B.n467 VSUBS 0.008123f
C642 B.n468 VSUBS 0.008123f
C643 B.n469 VSUBS 0.008123f
C644 B.n470 VSUBS 0.008123f
C645 B.n471 VSUBS 0.008123f
C646 B.n472 VSUBS 0.008123f
C647 B.n473 VSUBS 0.008123f
C648 B.n474 VSUBS 0.008123f
C649 B.n475 VSUBS 0.008123f
C650 B.n476 VSUBS 0.008123f
C651 B.n477 VSUBS 0.008123f
C652 B.n478 VSUBS 0.008123f
C653 B.n479 VSUBS 0.008123f
C654 B.n480 VSUBS 0.008123f
C655 B.n481 VSUBS 0.008123f
C656 B.n482 VSUBS 0.008123f
C657 B.n483 VSUBS 0.008123f
C658 B.n484 VSUBS 0.008123f
C659 B.n485 VSUBS 0.008123f
C660 B.n486 VSUBS 0.008123f
C661 B.n487 VSUBS 0.008123f
C662 B.n488 VSUBS 0.008123f
C663 B.n489 VSUBS 0.008123f
C664 B.n490 VSUBS 0.008123f
C665 B.n491 VSUBS 0.008123f
C666 B.n492 VSUBS 0.008123f
C667 B.n493 VSUBS 0.008123f
C668 B.n494 VSUBS 0.008123f
C669 B.n495 VSUBS 0.008123f
C670 B.n496 VSUBS 0.008123f
C671 B.n497 VSUBS 0.008123f
C672 B.n498 VSUBS 0.008123f
C673 B.n499 VSUBS 0.008123f
C674 B.n500 VSUBS 0.008123f
C675 B.n501 VSUBS 0.008123f
C676 B.n502 VSUBS 0.008123f
C677 B.n503 VSUBS 0.008123f
C678 B.n504 VSUBS 0.008123f
C679 B.n505 VSUBS 0.008123f
C680 B.n506 VSUBS 0.008123f
C681 B.n507 VSUBS 0.008123f
C682 B.n508 VSUBS 0.008123f
C683 B.n509 VSUBS 0.008123f
C684 B.n510 VSUBS 0.008123f
C685 B.n511 VSUBS 0.008123f
C686 B.n512 VSUBS 0.008123f
C687 B.n513 VSUBS 0.008123f
C688 B.n514 VSUBS 0.008123f
C689 B.n515 VSUBS 0.008123f
C690 B.n516 VSUBS 0.008123f
C691 B.n517 VSUBS 0.008123f
C692 B.n518 VSUBS 0.008123f
C693 B.n519 VSUBS 0.008123f
C694 B.n520 VSUBS 0.008123f
C695 B.n521 VSUBS 0.008123f
C696 B.n522 VSUBS 0.008123f
C697 B.n523 VSUBS 0.008123f
C698 B.n524 VSUBS 0.008123f
C699 B.n525 VSUBS 0.008123f
C700 B.n526 VSUBS 0.008123f
C701 B.n527 VSUBS 0.008123f
C702 B.n528 VSUBS 0.008123f
C703 B.n529 VSUBS 0.008123f
C704 B.n530 VSUBS 0.008123f
C705 B.n531 VSUBS 0.008123f
C706 B.n532 VSUBS 0.008123f
C707 B.n533 VSUBS 0.008123f
C708 B.n534 VSUBS 0.008123f
C709 B.n535 VSUBS 0.008123f
C710 B.n536 VSUBS 0.008123f
C711 B.n537 VSUBS 0.008123f
C712 B.n538 VSUBS 0.008123f
C713 B.n539 VSUBS 0.008123f
C714 B.n540 VSUBS 0.008123f
C715 B.n541 VSUBS 0.008123f
C716 B.n542 VSUBS 0.008123f
C717 B.n543 VSUBS 0.008123f
C718 B.n544 VSUBS 0.008123f
C719 B.n545 VSUBS 0.008123f
C720 B.n546 VSUBS 0.008123f
C721 B.n547 VSUBS 0.008123f
C722 B.n548 VSUBS 0.008123f
C723 B.n549 VSUBS 0.008123f
C724 B.n550 VSUBS 0.008123f
C725 B.n551 VSUBS 0.008123f
C726 B.n552 VSUBS 0.008123f
C727 B.n553 VSUBS 0.008123f
C728 B.n554 VSUBS 0.008123f
C729 B.n555 VSUBS 0.008123f
C730 B.n556 VSUBS 0.008123f
C731 B.n557 VSUBS 0.008123f
C732 B.n558 VSUBS 0.008123f
C733 B.n559 VSUBS 0.008123f
C734 B.n560 VSUBS 0.008123f
C735 B.n561 VSUBS 0.008123f
C736 B.n562 VSUBS 0.008123f
C737 B.n563 VSUBS 0.008123f
C738 B.n564 VSUBS 0.008123f
C739 B.n565 VSUBS 0.008123f
C740 B.n566 VSUBS 0.008123f
C741 B.n567 VSUBS 0.008123f
C742 B.n568 VSUBS 0.008123f
C743 B.n569 VSUBS 0.008123f
C744 B.n570 VSUBS 0.008123f
C745 B.n571 VSUBS 0.008123f
C746 B.n572 VSUBS 0.008123f
C747 B.n573 VSUBS 0.008123f
C748 B.n574 VSUBS 0.008123f
C749 B.n575 VSUBS 0.008123f
C750 B.n576 VSUBS 0.008123f
C751 B.n577 VSUBS 0.008123f
C752 B.n578 VSUBS 0.008123f
C753 B.n579 VSUBS 0.008123f
C754 B.n580 VSUBS 0.008123f
C755 B.n581 VSUBS 0.008123f
C756 B.n582 VSUBS 0.008123f
C757 B.n583 VSUBS 0.008123f
C758 B.n584 VSUBS 0.008123f
C759 B.n585 VSUBS 0.008123f
C760 B.n586 VSUBS 0.020489f
C761 B.n587 VSUBS 0.020489f
C762 B.n588 VSUBS 0.021322f
C763 B.n589 VSUBS 0.008123f
C764 B.n590 VSUBS 0.008123f
C765 B.n591 VSUBS 0.008123f
C766 B.n592 VSUBS 0.008123f
C767 B.n593 VSUBS 0.008123f
C768 B.n594 VSUBS 0.008123f
C769 B.n595 VSUBS 0.008123f
C770 B.n596 VSUBS 0.008123f
C771 B.n597 VSUBS 0.008123f
C772 B.n598 VSUBS 0.008123f
C773 B.n599 VSUBS 0.008123f
C774 B.n600 VSUBS 0.008123f
C775 B.n601 VSUBS 0.008123f
C776 B.n602 VSUBS 0.008123f
C777 B.n603 VSUBS 0.008123f
C778 B.n604 VSUBS 0.008123f
C779 B.n605 VSUBS 0.008123f
C780 B.n606 VSUBS 0.008123f
C781 B.n607 VSUBS 0.008123f
C782 B.n608 VSUBS 0.008123f
C783 B.n609 VSUBS 0.008123f
C784 B.n610 VSUBS 0.008123f
C785 B.n611 VSUBS 0.008123f
C786 B.n612 VSUBS 0.008123f
C787 B.n613 VSUBS 0.008123f
C788 B.n614 VSUBS 0.008123f
C789 B.n615 VSUBS 0.008123f
C790 B.n616 VSUBS 0.008123f
C791 B.n617 VSUBS 0.008123f
C792 B.n618 VSUBS 0.008123f
C793 B.n619 VSUBS 0.008123f
C794 B.n620 VSUBS 0.008123f
C795 B.n621 VSUBS 0.008123f
C796 B.n622 VSUBS 0.008123f
C797 B.n623 VSUBS 0.008123f
C798 B.n624 VSUBS 0.008123f
C799 B.n625 VSUBS 0.008123f
C800 B.n626 VSUBS 0.008123f
C801 B.n627 VSUBS 0.008123f
C802 B.n628 VSUBS 0.008123f
C803 B.n629 VSUBS 0.008123f
C804 B.n630 VSUBS 0.008123f
C805 B.n631 VSUBS 0.008123f
C806 B.n632 VSUBS 0.008123f
C807 B.n633 VSUBS 0.008123f
C808 B.n634 VSUBS 0.008123f
C809 B.n635 VSUBS 0.008123f
C810 B.n636 VSUBS 0.008123f
C811 B.n637 VSUBS 0.008123f
C812 B.n638 VSUBS 0.008123f
C813 B.n639 VSUBS 0.008123f
C814 B.n640 VSUBS 0.008123f
C815 B.n641 VSUBS 0.008123f
C816 B.n642 VSUBS 0.008123f
C817 B.n643 VSUBS 0.008123f
C818 B.n644 VSUBS 0.008123f
C819 B.n645 VSUBS 0.008123f
C820 B.n646 VSUBS 0.008123f
C821 B.n647 VSUBS 0.008123f
C822 B.n648 VSUBS 0.008123f
C823 B.n649 VSUBS 0.008123f
C824 B.n650 VSUBS 0.008123f
C825 B.n651 VSUBS 0.008123f
C826 B.n652 VSUBS 0.008123f
C827 B.n653 VSUBS 0.008123f
C828 B.n654 VSUBS 0.008123f
C829 B.n655 VSUBS 0.008123f
C830 B.n656 VSUBS 0.008123f
C831 B.n657 VSUBS 0.008123f
C832 B.n658 VSUBS 0.008123f
C833 B.n659 VSUBS 0.008123f
C834 B.n660 VSUBS 0.005615f
C835 B.n661 VSUBS 0.018821f
C836 B.n662 VSUBS 0.00657f
C837 B.n663 VSUBS 0.008123f
C838 B.n664 VSUBS 0.008123f
C839 B.n665 VSUBS 0.008123f
C840 B.n666 VSUBS 0.008123f
C841 B.n667 VSUBS 0.008123f
C842 B.n668 VSUBS 0.008123f
C843 B.n669 VSUBS 0.008123f
C844 B.n670 VSUBS 0.008123f
C845 B.n671 VSUBS 0.008123f
C846 B.n672 VSUBS 0.008123f
C847 B.n673 VSUBS 0.008123f
C848 B.n674 VSUBS 0.00657f
C849 B.n675 VSUBS 0.008123f
C850 B.n676 VSUBS 0.008123f
C851 B.n677 VSUBS 0.005615f
C852 B.n678 VSUBS 0.008123f
C853 B.n679 VSUBS 0.008123f
C854 B.n680 VSUBS 0.008123f
C855 B.n681 VSUBS 0.008123f
C856 B.n682 VSUBS 0.008123f
C857 B.n683 VSUBS 0.008123f
C858 B.n684 VSUBS 0.008123f
C859 B.n685 VSUBS 0.008123f
C860 B.n686 VSUBS 0.008123f
C861 B.n687 VSUBS 0.008123f
C862 B.n688 VSUBS 0.008123f
C863 B.n689 VSUBS 0.008123f
C864 B.n690 VSUBS 0.008123f
C865 B.n691 VSUBS 0.008123f
C866 B.n692 VSUBS 0.008123f
C867 B.n693 VSUBS 0.008123f
C868 B.n694 VSUBS 0.008123f
C869 B.n695 VSUBS 0.008123f
C870 B.n696 VSUBS 0.008123f
C871 B.n697 VSUBS 0.008123f
C872 B.n698 VSUBS 0.008123f
C873 B.n699 VSUBS 0.008123f
C874 B.n700 VSUBS 0.008123f
C875 B.n701 VSUBS 0.008123f
C876 B.n702 VSUBS 0.008123f
C877 B.n703 VSUBS 0.008123f
C878 B.n704 VSUBS 0.008123f
C879 B.n705 VSUBS 0.008123f
C880 B.n706 VSUBS 0.008123f
C881 B.n707 VSUBS 0.008123f
C882 B.n708 VSUBS 0.008123f
C883 B.n709 VSUBS 0.008123f
C884 B.n710 VSUBS 0.008123f
C885 B.n711 VSUBS 0.008123f
C886 B.n712 VSUBS 0.008123f
C887 B.n713 VSUBS 0.008123f
C888 B.n714 VSUBS 0.008123f
C889 B.n715 VSUBS 0.008123f
C890 B.n716 VSUBS 0.008123f
C891 B.n717 VSUBS 0.008123f
C892 B.n718 VSUBS 0.008123f
C893 B.n719 VSUBS 0.008123f
C894 B.n720 VSUBS 0.008123f
C895 B.n721 VSUBS 0.008123f
C896 B.n722 VSUBS 0.008123f
C897 B.n723 VSUBS 0.008123f
C898 B.n724 VSUBS 0.008123f
C899 B.n725 VSUBS 0.008123f
C900 B.n726 VSUBS 0.008123f
C901 B.n727 VSUBS 0.008123f
C902 B.n728 VSUBS 0.008123f
C903 B.n729 VSUBS 0.008123f
C904 B.n730 VSUBS 0.008123f
C905 B.n731 VSUBS 0.008123f
C906 B.n732 VSUBS 0.008123f
C907 B.n733 VSUBS 0.008123f
C908 B.n734 VSUBS 0.008123f
C909 B.n735 VSUBS 0.008123f
C910 B.n736 VSUBS 0.008123f
C911 B.n737 VSUBS 0.008123f
C912 B.n738 VSUBS 0.008123f
C913 B.n739 VSUBS 0.008123f
C914 B.n740 VSUBS 0.008123f
C915 B.n741 VSUBS 0.008123f
C916 B.n742 VSUBS 0.008123f
C917 B.n743 VSUBS 0.008123f
C918 B.n744 VSUBS 0.008123f
C919 B.n745 VSUBS 0.008123f
C920 B.n746 VSUBS 0.008123f
C921 B.n747 VSUBS 0.008123f
C922 B.n748 VSUBS 0.021322f
C923 B.n749 VSUBS 0.021322f
C924 B.n750 VSUBS 0.020489f
C925 B.n751 VSUBS 0.008123f
C926 B.n752 VSUBS 0.008123f
C927 B.n753 VSUBS 0.008123f
C928 B.n754 VSUBS 0.008123f
C929 B.n755 VSUBS 0.008123f
C930 B.n756 VSUBS 0.008123f
C931 B.n757 VSUBS 0.008123f
C932 B.n758 VSUBS 0.008123f
C933 B.n759 VSUBS 0.008123f
C934 B.n760 VSUBS 0.008123f
C935 B.n761 VSUBS 0.008123f
C936 B.n762 VSUBS 0.008123f
C937 B.n763 VSUBS 0.008123f
C938 B.n764 VSUBS 0.008123f
C939 B.n765 VSUBS 0.008123f
C940 B.n766 VSUBS 0.008123f
C941 B.n767 VSUBS 0.008123f
C942 B.n768 VSUBS 0.008123f
C943 B.n769 VSUBS 0.008123f
C944 B.n770 VSUBS 0.008123f
C945 B.n771 VSUBS 0.008123f
C946 B.n772 VSUBS 0.008123f
C947 B.n773 VSUBS 0.008123f
C948 B.n774 VSUBS 0.008123f
C949 B.n775 VSUBS 0.008123f
C950 B.n776 VSUBS 0.008123f
C951 B.n777 VSUBS 0.008123f
C952 B.n778 VSUBS 0.008123f
C953 B.n779 VSUBS 0.008123f
C954 B.n780 VSUBS 0.008123f
C955 B.n781 VSUBS 0.008123f
C956 B.n782 VSUBS 0.008123f
C957 B.n783 VSUBS 0.008123f
C958 B.n784 VSUBS 0.008123f
C959 B.n785 VSUBS 0.008123f
C960 B.n786 VSUBS 0.008123f
C961 B.n787 VSUBS 0.008123f
C962 B.n788 VSUBS 0.008123f
C963 B.n789 VSUBS 0.008123f
C964 B.n790 VSUBS 0.008123f
C965 B.n791 VSUBS 0.008123f
C966 B.n792 VSUBS 0.008123f
C967 B.n793 VSUBS 0.008123f
C968 B.n794 VSUBS 0.008123f
C969 B.n795 VSUBS 0.008123f
C970 B.n796 VSUBS 0.008123f
C971 B.n797 VSUBS 0.008123f
C972 B.n798 VSUBS 0.008123f
C973 B.n799 VSUBS 0.008123f
C974 B.n800 VSUBS 0.008123f
C975 B.n801 VSUBS 0.008123f
C976 B.n802 VSUBS 0.008123f
C977 B.n803 VSUBS 0.008123f
C978 B.n804 VSUBS 0.008123f
C979 B.n805 VSUBS 0.008123f
C980 B.n806 VSUBS 0.008123f
C981 B.n807 VSUBS 0.008123f
C982 B.n808 VSUBS 0.008123f
C983 B.n809 VSUBS 0.008123f
C984 B.n810 VSUBS 0.008123f
C985 B.n811 VSUBS 0.008123f
C986 B.n812 VSUBS 0.008123f
C987 B.n813 VSUBS 0.008123f
C988 B.n814 VSUBS 0.008123f
C989 B.n815 VSUBS 0.008123f
C990 B.n816 VSUBS 0.008123f
C991 B.n817 VSUBS 0.008123f
C992 B.n818 VSUBS 0.008123f
C993 B.n819 VSUBS 0.0106f
C994 B.n820 VSUBS 0.011292f
C995 B.n821 VSUBS 0.022455f
.ends

