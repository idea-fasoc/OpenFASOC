* NGSPICE file created from diff_pair_sample_0712.ext - technology: sky130A

.subckt diff_pair_sample_0712 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t18 VN.t0 VDD2.t3 w_n3130_n2852# sky130_fd_pr__pfet_01v8 ad=1.5543 pd=9.75 as=1.5543 ps=9.75 w=9.42 l=1.47
X1 VDD1.t9 VP.t0 VTAIL.t8 w_n3130_n2852# sky130_fd_pr__pfet_01v8 ad=3.6738 pd=19.62 as=1.5543 ps=9.75 w=9.42 l=1.47
X2 VTAIL.t19 VP.t1 VDD1.t8 w_n3130_n2852# sky130_fd_pr__pfet_01v8 ad=1.5543 pd=9.75 as=1.5543 ps=9.75 w=9.42 l=1.47
X3 VDD1.t7 VP.t2 VTAIL.t4 w_n3130_n2852# sky130_fd_pr__pfet_01v8 ad=1.5543 pd=9.75 as=3.6738 ps=19.62 w=9.42 l=1.47
X4 B.t11 B.t9 B.t10 w_n3130_n2852# sky130_fd_pr__pfet_01v8 ad=3.6738 pd=19.62 as=0 ps=0 w=9.42 l=1.47
X5 VTAIL.t17 VN.t1 VDD2.t1 w_n3130_n2852# sky130_fd_pr__pfet_01v8 ad=1.5543 pd=9.75 as=1.5543 ps=9.75 w=9.42 l=1.47
X6 VDD2.t8 VN.t2 VTAIL.t16 w_n3130_n2852# sky130_fd_pr__pfet_01v8 ad=1.5543 pd=9.75 as=3.6738 ps=19.62 w=9.42 l=1.47
X7 VDD2.t6 VN.t3 VTAIL.t15 w_n3130_n2852# sky130_fd_pr__pfet_01v8 ad=3.6738 pd=19.62 as=1.5543 ps=9.75 w=9.42 l=1.47
X8 VDD1.t6 VP.t3 VTAIL.t5 w_n3130_n2852# sky130_fd_pr__pfet_01v8 ad=1.5543 pd=9.75 as=1.5543 ps=9.75 w=9.42 l=1.47
X9 VDD1.t5 VP.t4 VTAIL.t3 w_n3130_n2852# sky130_fd_pr__pfet_01v8 ad=3.6738 pd=19.62 as=1.5543 ps=9.75 w=9.42 l=1.47
X10 VDD2.t5 VN.t4 VTAIL.t14 w_n3130_n2852# sky130_fd_pr__pfet_01v8 ad=1.5543 pd=9.75 as=1.5543 ps=9.75 w=9.42 l=1.47
X11 VDD2.t4 VN.t5 VTAIL.t13 w_n3130_n2852# sky130_fd_pr__pfet_01v8 ad=1.5543 pd=9.75 as=3.6738 ps=19.62 w=9.42 l=1.47
X12 B.t8 B.t6 B.t7 w_n3130_n2852# sky130_fd_pr__pfet_01v8 ad=3.6738 pd=19.62 as=0 ps=0 w=9.42 l=1.47
X13 VDD1.t4 VP.t5 VTAIL.t6 w_n3130_n2852# sky130_fd_pr__pfet_01v8 ad=1.5543 pd=9.75 as=3.6738 ps=19.62 w=9.42 l=1.47
X14 B.t5 B.t3 B.t4 w_n3130_n2852# sky130_fd_pr__pfet_01v8 ad=3.6738 pd=19.62 as=0 ps=0 w=9.42 l=1.47
X15 VTAIL.t0 VP.t6 VDD1.t3 w_n3130_n2852# sky130_fd_pr__pfet_01v8 ad=1.5543 pd=9.75 as=1.5543 ps=9.75 w=9.42 l=1.47
X16 VDD2.t9 VN.t6 VTAIL.t12 w_n3130_n2852# sky130_fd_pr__pfet_01v8 ad=3.6738 pd=19.62 as=1.5543 ps=9.75 w=9.42 l=1.47
X17 VDD1.t2 VP.t7 VTAIL.t1 w_n3130_n2852# sky130_fd_pr__pfet_01v8 ad=1.5543 pd=9.75 as=1.5543 ps=9.75 w=9.42 l=1.47
X18 B.t2 B.t0 B.t1 w_n3130_n2852# sky130_fd_pr__pfet_01v8 ad=3.6738 pd=19.62 as=0 ps=0 w=9.42 l=1.47
X19 VTAIL.t11 VN.t7 VDD2.t0 w_n3130_n2852# sky130_fd_pr__pfet_01v8 ad=1.5543 pd=9.75 as=1.5543 ps=9.75 w=9.42 l=1.47
X20 VTAIL.t2 VP.t8 VDD1.t1 w_n3130_n2852# sky130_fd_pr__pfet_01v8 ad=1.5543 pd=9.75 as=1.5543 ps=9.75 w=9.42 l=1.47
X21 VDD2.t2 VN.t8 VTAIL.t10 w_n3130_n2852# sky130_fd_pr__pfet_01v8 ad=1.5543 pd=9.75 as=1.5543 ps=9.75 w=9.42 l=1.47
X22 VTAIL.t9 VN.t9 VDD2.t7 w_n3130_n2852# sky130_fd_pr__pfet_01v8 ad=1.5543 pd=9.75 as=1.5543 ps=9.75 w=9.42 l=1.47
X23 VTAIL.t7 VP.t9 VDD1.t0 w_n3130_n2852# sky130_fd_pr__pfet_01v8 ad=1.5543 pd=9.75 as=1.5543 ps=9.75 w=9.42 l=1.47
R0 VN.n7 VN.t6 185.481
R1 VN.n34 VN.t5 185.481
R2 VN.n26 VN.n25 180.974
R3 VN.n53 VN.n52 180.974
R4 VN.n51 VN.n27 161.3
R5 VN.n50 VN.n49 161.3
R6 VN.n48 VN.n28 161.3
R7 VN.n47 VN.n46 161.3
R8 VN.n44 VN.n29 161.3
R9 VN.n43 VN.n42 161.3
R10 VN.n41 VN.n30 161.3
R11 VN.n40 VN.n39 161.3
R12 VN.n38 VN.n31 161.3
R13 VN.n37 VN.n36 161.3
R14 VN.n35 VN.n32 161.3
R15 VN.n24 VN.n0 161.3
R16 VN.n23 VN.n22 161.3
R17 VN.n21 VN.n1 161.3
R18 VN.n20 VN.n19 161.3
R19 VN.n17 VN.n2 161.3
R20 VN.n16 VN.n15 161.3
R21 VN.n14 VN.n3 161.3
R22 VN.n13 VN.n12 161.3
R23 VN.n11 VN.n4 161.3
R24 VN.n10 VN.n9 161.3
R25 VN.n8 VN.n5 161.3
R26 VN.n12 VN.t4 154.438
R27 VN.n6 VN.t9 154.438
R28 VN.n18 VN.t0 154.438
R29 VN.n25 VN.t2 154.438
R30 VN.n39 VN.t8 154.438
R31 VN.n33 VN.t1 154.438
R32 VN.n45 VN.t7 154.438
R33 VN.n52 VN.t3 154.438
R34 VN.n23 VN.n1 56.5617
R35 VN.n50 VN.n28 56.5617
R36 VN.n7 VN.n6 51.3232
R37 VN.n34 VN.n33 51.3232
R38 VN.n11 VN.n10 50.2647
R39 VN.n16 VN.n3 50.2647
R40 VN.n38 VN.n37 50.2647
R41 VN.n43 VN.n30 50.2647
R42 VN VN.n53 45.2372
R43 VN.n10 VN.n5 30.8893
R44 VN.n17 VN.n16 30.8893
R45 VN.n37 VN.n32 30.8893
R46 VN.n44 VN.n43 30.8893
R47 VN.n12 VN.n11 24.5923
R48 VN.n12 VN.n3 24.5923
R49 VN.n19 VN.n1 24.5923
R50 VN.n24 VN.n23 24.5923
R51 VN.n39 VN.n30 24.5923
R52 VN.n39 VN.n38 24.5923
R53 VN.n46 VN.n28 24.5923
R54 VN.n51 VN.n50 24.5923
R55 VN.n35 VN.n34 18.2653
R56 VN.n8 VN.n7 18.2653
R57 VN.n6 VN.n5 14.7556
R58 VN.n18 VN.n17 14.7556
R59 VN.n33 VN.n32 14.7556
R60 VN.n45 VN.n44 14.7556
R61 VN.n19 VN.n18 9.83723
R62 VN.n46 VN.n45 9.83723
R63 VN.n25 VN.n24 4.91887
R64 VN.n52 VN.n51 4.91887
R65 VN.n53 VN.n27 0.189894
R66 VN.n49 VN.n27 0.189894
R67 VN.n49 VN.n48 0.189894
R68 VN.n48 VN.n47 0.189894
R69 VN.n47 VN.n29 0.189894
R70 VN.n42 VN.n29 0.189894
R71 VN.n42 VN.n41 0.189894
R72 VN.n41 VN.n40 0.189894
R73 VN.n40 VN.n31 0.189894
R74 VN.n36 VN.n31 0.189894
R75 VN.n36 VN.n35 0.189894
R76 VN.n9 VN.n8 0.189894
R77 VN.n9 VN.n4 0.189894
R78 VN.n13 VN.n4 0.189894
R79 VN.n14 VN.n13 0.189894
R80 VN.n15 VN.n14 0.189894
R81 VN.n15 VN.n2 0.189894
R82 VN.n20 VN.n2 0.189894
R83 VN.n21 VN.n20 0.189894
R84 VN.n22 VN.n21 0.189894
R85 VN.n22 VN.n0 0.189894
R86 VN.n26 VN.n0 0.189894
R87 VN VN.n26 0.0516364
R88 VDD2.n97 VDD2.n53 756.745
R89 VDD2.n44 VDD2.n0 756.745
R90 VDD2.n98 VDD2.n97 585
R91 VDD2.n96 VDD2.n95 585
R92 VDD2.n57 VDD2.n56 585
R93 VDD2.n61 VDD2.n59 585
R94 VDD2.n90 VDD2.n89 585
R95 VDD2.n88 VDD2.n87 585
R96 VDD2.n63 VDD2.n62 585
R97 VDD2.n82 VDD2.n81 585
R98 VDD2.n80 VDD2.n79 585
R99 VDD2.n67 VDD2.n66 585
R100 VDD2.n74 VDD2.n73 585
R101 VDD2.n72 VDD2.n71 585
R102 VDD2.n17 VDD2.n16 585
R103 VDD2.n19 VDD2.n18 585
R104 VDD2.n12 VDD2.n11 585
R105 VDD2.n25 VDD2.n24 585
R106 VDD2.n27 VDD2.n26 585
R107 VDD2.n8 VDD2.n7 585
R108 VDD2.n34 VDD2.n33 585
R109 VDD2.n35 VDD2.n6 585
R110 VDD2.n37 VDD2.n36 585
R111 VDD2.n4 VDD2.n3 585
R112 VDD2.n43 VDD2.n42 585
R113 VDD2.n45 VDD2.n44 585
R114 VDD2.n70 VDD2.t6 329.038
R115 VDD2.n15 VDD2.t9 329.038
R116 VDD2.n97 VDD2.n96 171.744
R117 VDD2.n96 VDD2.n56 171.744
R118 VDD2.n61 VDD2.n56 171.744
R119 VDD2.n89 VDD2.n61 171.744
R120 VDD2.n89 VDD2.n88 171.744
R121 VDD2.n88 VDD2.n62 171.744
R122 VDD2.n81 VDD2.n62 171.744
R123 VDD2.n81 VDD2.n80 171.744
R124 VDD2.n80 VDD2.n66 171.744
R125 VDD2.n73 VDD2.n66 171.744
R126 VDD2.n73 VDD2.n72 171.744
R127 VDD2.n18 VDD2.n17 171.744
R128 VDD2.n18 VDD2.n11 171.744
R129 VDD2.n25 VDD2.n11 171.744
R130 VDD2.n26 VDD2.n25 171.744
R131 VDD2.n26 VDD2.n7 171.744
R132 VDD2.n34 VDD2.n7 171.744
R133 VDD2.n35 VDD2.n34 171.744
R134 VDD2.n36 VDD2.n35 171.744
R135 VDD2.n36 VDD2.n3 171.744
R136 VDD2.n43 VDD2.n3 171.744
R137 VDD2.n44 VDD2.n43 171.744
R138 VDD2.n72 VDD2.t6 85.8723
R139 VDD2.n17 VDD2.t9 85.8723
R140 VDD2.n52 VDD2.n51 83.1801
R141 VDD2 VDD2.n105 83.1772
R142 VDD2.n104 VDD2.n103 82.0718
R143 VDD2.n50 VDD2.n49 82.0716
R144 VDD2.n50 VDD2.n48 53.9068
R145 VDD2.n102 VDD2.n101 52.355
R146 VDD2.n102 VDD2.n52 39.2067
R147 VDD2.n59 VDD2.n57 13.1884
R148 VDD2.n37 VDD2.n4 13.1884
R149 VDD2.n95 VDD2.n94 12.8005
R150 VDD2.n91 VDD2.n90 12.8005
R151 VDD2.n38 VDD2.n6 12.8005
R152 VDD2.n42 VDD2.n41 12.8005
R153 VDD2.n98 VDD2.n55 12.0247
R154 VDD2.n87 VDD2.n60 12.0247
R155 VDD2.n33 VDD2.n32 12.0247
R156 VDD2.n45 VDD2.n2 12.0247
R157 VDD2.n99 VDD2.n53 11.249
R158 VDD2.n86 VDD2.n63 11.249
R159 VDD2.n31 VDD2.n8 11.249
R160 VDD2.n46 VDD2.n0 11.249
R161 VDD2.n71 VDD2.n70 10.7239
R162 VDD2.n16 VDD2.n15 10.7239
R163 VDD2.n83 VDD2.n82 10.4732
R164 VDD2.n28 VDD2.n27 10.4732
R165 VDD2.n79 VDD2.n65 9.69747
R166 VDD2.n24 VDD2.n10 9.69747
R167 VDD2.n101 VDD2.n100 9.45567
R168 VDD2.n48 VDD2.n47 9.45567
R169 VDD2.n69 VDD2.n68 9.3005
R170 VDD2.n76 VDD2.n75 9.3005
R171 VDD2.n78 VDD2.n77 9.3005
R172 VDD2.n65 VDD2.n64 9.3005
R173 VDD2.n84 VDD2.n83 9.3005
R174 VDD2.n86 VDD2.n85 9.3005
R175 VDD2.n60 VDD2.n58 9.3005
R176 VDD2.n92 VDD2.n91 9.3005
R177 VDD2.n100 VDD2.n99 9.3005
R178 VDD2.n55 VDD2.n54 9.3005
R179 VDD2.n94 VDD2.n93 9.3005
R180 VDD2.n47 VDD2.n46 9.3005
R181 VDD2.n2 VDD2.n1 9.3005
R182 VDD2.n41 VDD2.n40 9.3005
R183 VDD2.n14 VDD2.n13 9.3005
R184 VDD2.n21 VDD2.n20 9.3005
R185 VDD2.n23 VDD2.n22 9.3005
R186 VDD2.n10 VDD2.n9 9.3005
R187 VDD2.n29 VDD2.n28 9.3005
R188 VDD2.n31 VDD2.n30 9.3005
R189 VDD2.n32 VDD2.n5 9.3005
R190 VDD2.n39 VDD2.n38 9.3005
R191 VDD2.n78 VDD2.n67 8.92171
R192 VDD2.n23 VDD2.n12 8.92171
R193 VDD2.n75 VDD2.n74 8.14595
R194 VDD2.n20 VDD2.n19 8.14595
R195 VDD2.n71 VDD2.n69 7.3702
R196 VDD2.n16 VDD2.n14 7.3702
R197 VDD2.n74 VDD2.n69 5.81868
R198 VDD2.n19 VDD2.n14 5.81868
R199 VDD2.n75 VDD2.n67 5.04292
R200 VDD2.n20 VDD2.n12 5.04292
R201 VDD2.n79 VDD2.n78 4.26717
R202 VDD2.n24 VDD2.n23 4.26717
R203 VDD2.n82 VDD2.n65 3.49141
R204 VDD2.n27 VDD2.n10 3.49141
R205 VDD2.n105 VDD2.t1 3.45114
R206 VDD2.n105 VDD2.t4 3.45114
R207 VDD2.n103 VDD2.t0 3.45114
R208 VDD2.n103 VDD2.t2 3.45114
R209 VDD2.n51 VDD2.t3 3.45114
R210 VDD2.n51 VDD2.t8 3.45114
R211 VDD2.n49 VDD2.t7 3.45114
R212 VDD2.n49 VDD2.t5 3.45114
R213 VDD2.n101 VDD2.n53 2.71565
R214 VDD2.n83 VDD2.n63 2.71565
R215 VDD2.n28 VDD2.n8 2.71565
R216 VDD2.n48 VDD2.n0 2.71565
R217 VDD2.n70 VDD2.n68 2.41283
R218 VDD2.n15 VDD2.n13 2.41283
R219 VDD2.n99 VDD2.n98 1.93989
R220 VDD2.n87 VDD2.n86 1.93989
R221 VDD2.n33 VDD2.n31 1.93989
R222 VDD2.n46 VDD2.n45 1.93989
R223 VDD2.n104 VDD2.n102 1.55222
R224 VDD2.n95 VDD2.n55 1.16414
R225 VDD2.n90 VDD2.n60 1.16414
R226 VDD2.n32 VDD2.n6 1.16414
R227 VDD2.n42 VDD2.n2 1.16414
R228 VDD2 VDD2.n104 0.446621
R229 VDD2.n94 VDD2.n57 0.388379
R230 VDD2.n91 VDD2.n59 0.388379
R231 VDD2.n38 VDD2.n37 0.388379
R232 VDD2.n41 VDD2.n4 0.388379
R233 VDD2.n52 VDD2.n50 0.333085
R234 VDD2.n100 VDD2.n54 0.155672
R235 VDD2.n93 VDD2.n54 0.155672
R236 VDD2.n93 VDD2.n92 0.155672
R237 VDD2.n92 VDD2.n58 0.155672
R238 VDD2.n85 VDD2.n58 0.155672
R239 VDD2.n85 VDD2.n84 0.155672
R240 VDD2.n84 VDD2.n64 0.155672
R241 VDD2.n77 VDD2.n64 0.155672
R242 VDD2.n77 VDD2.n76 0.155672
R243 VDD2.n76 VDD2.n68 0.155672
R244 VDD2.n21 VDD2.n13 0.155672
R245 VDD2.n22 VDD2.n21 0.155672
R246 VDD2.n22 VDD2.n9 0.155672
R247 VDD2.n29 VDD2.n9 0.155672
R248 VDD2.n30 VDD2.n29 0.155672
R249 VDD2.n30 VDD2.n5 0.155672
R250 VDD2.n39 VDD2.n5 0.155672
R251 VDD2.n40 VDD2.n39 0.155672
R252 VDD2.n40 VDD2.n1 0.155672
R253 VDD2.n47 VDD2.n1 0.155672
R254 VTAIL.n208 VTAIL.n164 756.745
R255 VTAIL.n46 VTAIL.n2 756.745
R256 VTAIL.n158 VTAIL.n114 756.745
R257 VTAIL.n104 VTAIL.n60 756.745
R258 VTAIL.n181 VTAIL.n180 585
R259 VTAIL.n183 VTAIL.n182 585
R260 VTAIL.n176 VTAIL.n175 585
R261 VTAIL.n189 VTAIL.n188 585
R262 VTAIL.n191 VTAIL.n190 585
R263 VTAIL.n172 VTAIL.n171 585
R264 VTAIL.n198 VTAIL.n197 585
R265 VTAIL.n199 VTAIL.n170 585
R266 VTAIL.n201 VTAIL.n200 585
R267 VTAIL.n168 VTAIL.n167 585
R268 VTAIL.n207 VTAIL.n206 585
R269 VTAIL.n209 VTAIL.n208 585
R270 VTAIL.n19 VTAIL.n18 585
R271 VTAIL.n21 VTAIL.n20 585
R272 VTAIL.n14 VTAIL.n13 585
R273 VTAIL.n27 VTAIL.n26 585
R274 VTAIL.n29 VTAIL.n28 585
R275 VTAIL.n10 VTAIL.n9 585
R276 VTAIL.n36 VTAIL.n35 585
R277 VTAIL.n37 VTAIL.n8 585
R278 VTAIL.n39 VTAIL.n38 585
R279 VTAIL.n6 VTAIL.n5 585
R280 VTAIL.n45 VTAIL.n44 585
R281 VTAIL.n47 VTAIL.n46 585
R282 VTAIL.n159 VTAIL.n158 585
R283 VTAIL.n157 VTAIL.n156 585
R284 VTAIL.n118 VTAIL.n117 585
R285 VTAIL.n122 VTAIL.n120 585
R286 VTAIL.n151 VTAIL.n150 585
R287 VTAIL.n149 VTAIL.n148 585
R288 VTAIL.n124 VTAIL.n123 585
R289 VTAIL.n143 VTAIL.n142 585
R290 VTAIL.n141 VTAIL.n140 585
R291 VTAIL.n128 VTAIL.n127 585
R292 VTAIL.n135 VTAIL.n134 585
R293 VTAIL.n133 VTAIL.n132 585
R294 VTAIL.n105 VTAIL.n104 585
R295 VTAIL.n103 VTAIL.n102 585
R296 VTAIL.n64 VTAIL.n63 585
R297 VTAIL.n68 VTAIL.n66 585
R298 VTAIL.n97 VTAIL.n96 585
R299 VTAIL.n95 VTAIL.n94 585
R300 VTAIL.n70 VTAIL.n69 585
R301 VTAIL.n89 VTAIL.n88 585
R302 VTAIL.n87 VTAIL.n86 585
R303 VTAIL.n74 VTAIL.n73 585
R304 VTAIL.n81 VTAIL.n80 585
R305 VTAIL.n79 VTAIL.n78 585
R306 VTAIL.n179 VTAIL.t16 329.038
R307 VTAIL.n17 VTAIL.t6 329.038
R308 VTAIL.n131 VTAIL.t4 329.038
R309 VTAIL.n77 VTAIL.t13 329.038
R310 VTAIL.n182 VTAIL.n181 171.744
R311 VTAIL.n182 VTAIL.n175 171.744
R312 VTAIL.n189 VTAIL.n175 171.744
R313 VTAIL.n190 VTAIL.n189 171.744
R314 VTAIL.n190 VTAIL.n171 171.744
R315 VTAIL.n198 VTAIL.n171 171.744
R316 VTAIL.n199 VTAIL.n198 171.744
R317 VTAIL.n200 VTAIL.n199 171.744
R318 VTAIL.n200 VTAIL.n167 171.744
R319 VTAIL.n207 VTAIL.n167 171.744
R320 VTAIL.n208 VTAIL.n207 171.744
R321 VTAIL.n20 VTAIL.n19 171.744
R322 VTAIL.n20 VTAIL.n13 171.744
R323 VTAIL.n27 VTAIL.n13 171.744
R324 VTAIL.n28 VTAIL.n27 171.744
R325 VTAIL.n28 VTAIL.n9 171.744
R326 VTAIL.n36 VTAIL.n9 171.744
R327 VTAIL.n37 VTAIL.n36 171.744
R328 VTAIL.n38 VTAIL.n37 171.744
R329 VTAIL.n38 VTAIL.n5 171.744
R330 VTAIL.n45 VTAIL.n5 171.744
R331 VTAIL.n46 VTAIL.n45 171.744
R332 VTAIL.n158 VTAIL.n157 171.744
R333 VTAIL.n157 VTAIL.n117 171.744
R334 VTAIL.n122 VTAIL.n117 171.744
R335 VTAIL.n150 VTAIL.n122 171.744
R336 VTAIL.n150 VTAIL.n149 171.744
R337 VTAIL.n149 VTAIL.n123 171.744
R338 VTAIL.n142 VTAIL.n123 171.744
R339 VTAIL.n142 VTAIL.n141 171.744
R340 VTAIL.n141 VTAIL.n127 171.744
R341 VTAIL.n134 VTAIL.n127 171.744
R342 VTAIL.n134 VTAIL.n133 171.744
R343 VTAIL.n104 VTAIL.n103 171.744
R344 VTAIL.n103 VTAIL.n63 171.744
R345 VTAIL.n68 VTAIL.n63 171.744
R346 VTAIL.n96 VTAIL.n68 171.744
R347 VTAIL.n96 VTAIL.n95 171.744
R348 VTAIL.n95 VTAIL.n69 171.744
R349 VTAIL.n88 VTAIL.n69 171.744
R350 VTAIL.n88 VTAIL.n87 171.744
R351 VTAIL.n87 VTAIL.n73 171.744
R352 VTAIL.n80 VTAIL.n73 171.744
R353 VTAIL.n80 VTAIL.n79 171.744
R354 VTAIL.n181 VTAIL.t16 85.8723
R355 VTAIL.n19 VTAIL.t6 85.8723
R356 VTAIL.n133 VTAIL.t4 85.8723
R357 VTAIL.n79 VTAIL.t13 85.8723
R358 VTAIL.n113 VTAIL.n112 65.393
R359 VTAIL.n111 VTAIL.n110 65.393
R360 VTAIL.n59 VTAIL.n58 65.393
R361 VTAIL.n57 VTAIL.n56 65.393
R362 VTAIL.n215 VTAIL.n214 65.3928
R363 VTAIL.n1 VTAIL.n0 65.3928
R364 VTAIL.n53 VTAIL.n52 65.3928
R365 VTAIL.n55 VTAIL.n54 65.3928
R366 VTAIL.n213 VTAIL.n212 35.6763
R367 VTAIL.n51 VTAIL.n50 35.6763
R368 VTAIL.n163 VTAIL.n162 35.6763
R369 VTAIL.n109 VTAIL.n108 35.6763
R370 VTAIL.n57 VTAIL.n55 23.591
R371 VTAIL.n213 VTAIL.n163 22.0393
R372 VTAIL.n201 VTAIL.n168 13.1884
R373 VTAIL.n39 VTAIL.n6 13.1884
R374 VTAIL.n120 VTAIL.n118 13.1884
R375 VTAIL.n66 VTAIL.n64 13.1884
R376 VTAIL.n202 VTAIL.n170 12.8005
R377 VTAIL.n206 VTAIL.n205 12.8005
R378 VTAIL.n40 VTAIL.n8 12.8005
R379 VTAIL.n44 VTAIL.n43 12.8005
R380 VTAIL.n156 VTAIL.n155 12.8005
R381 VTAIL.n152 VTAIL.n151 12.8005
R382 VTAIL.n102 VTAIL.n101 12.8005
R383 VTAIL.n98 VTAIL.n97 12.8005
R384 VTAIL.n197 VTAIL.n196 12.0247
R385 VTAIL.n209 VTAIL.n166 12.0247
R386 VTAIL.n35 VTAIL.n34 12.0247
R387 VTAIL.n47 VTAIL.n4 12.0247
R388 VTAIL.n159 VTAIL.n116 12.0247
R389 VTAIL.n148 VTAIL.n121 12.0247
R390 VTAIL.n105 VTAIL.n62 12.0247
R391 VTAIL.n94 VTAIL.n67 12.0247
R392 VTAIL.n195 VTAIL.n172 11.249
R393 VTAIL.n210 VTAIL.n164 11.249
R394 VTAIL.n33 VTAIL.n10 11.249
R395 VTAIL.n48 VTAIL.n2 11.249
R396 VTAIL.n160 VTAIL.n114 11.249
R397 VTAIL.n147 VTAIL.n124 11.249
R398 VTAIL.n106 VTAIL.n60 11.249
R399 VTAIL.n93 VTAIL.n70 11.249
R400 VTAIL.n180 VTAIL.n179 10.7239
R401 VTAIL.n18 VTAIL.n17 10.7239
R402 VTAIL.n132 VTAIL.n131 10.7239
R403 VTAIL.n78 VTAIL.n77 10.7239
R404 VTAIL.n192 VTAIL.n191 10.4732
R405 VTAIL.n30 VTAIL.n29 10.4732
R406 VTAIL.n144 VTAIL.n143 10.4732
R407 VTAIL.n90 VTAIL.n89 10.4732
R408 VTAIL.n188 VTAIL.n174 9.69747
R409 VTAIL.n26 VTAIL.n12 9.69747
R410 VTAIL.n140 VTAIL.n126 9.69747
R411 VTAIL.n86 VTAIL.n72 9.69747
R412 VTAIL.n212 VTAIL.n211 9.45567
R413 VTAIL.n50 VTAIL.n49 9.45567
R414 VTAIL.n162 VTAIL.n161 9.45567
R415 VTAIL.n108 VTAIL.n107 9.45567
R416 VTAIL.n211 VTAIL.n210 9.3005
R417 VTAIL.n166 VTAIL.n165 9.3005
R418 VTAIL.n205 VTAIL.n204 9.3005
R419 VTAIL.n178 VTAIL.n177 9.3005
R420 VTAIL.n185 VTAIL.n184 9.3005
R421 VTAIL.n187 VTAIL.n186 9.3005
R422 VTAIL.n174 VTAIL.n173 9.3005
R423 VTAIL.n193 VTAIL.n192 9.3005
R424 VTAIL.n195 VTAIL.n194 9.3005
R425 VTAIL.n196 VTAIL.n169 9.3005
R426 VTAIL.n203 VTAIL.n202 9.3005
R427 VTAIL.n49 VTAIL.n48 9.3005
R428 VTAIL.n4 VTAIL.n3 9.3005
R429 VTAIL.n43 VTAIL.n42 9.3005
R430 VTAIL.n16 VTAIL.n15 9.3005
R431 VTAIL.n23 VTAIL.n22 9.3005
R432 VTAIL.n25 VTAIL.n24 9.3005
R433 VTAIL.n12 VTAIL.n11 9.3005
R434 VTAIL.n31 VTAIL.n30 9.3005
R435 VTAIL.n33 VTAIL.n32 9.3005
R436 VTAIL.n34 VTAIL.n7 9.3005
R437 VTAIL.n41 VTAIL.n40 9.3005
R438 VTAIL.n130 VTAIL.n129 9.3005
R439 VTAIL.n137 VTAIL.n136 9.3005
R440 VTAIL.n139 VTAIL.n138 9.3005
R441 VTAIL.n126 VTAIL.n125 9.3005
R442 VTAIL.n145 VTAIL.n144 9.3005
R443 VTAIL.n147 VTAIL.n146 9.3005
R444 VTAIL.n121 VTAIL.n119 9.3005
R445 VTAIL.n153 VTAIL.n152 9.3005
R446 VTAIL.n161 VTAIL.n160 9.3005
R447 VTAIL.n116 VTAIL.n115 9.3005
R448 VTAIL.n155 VTAIL.n154 9.3005
R449 VTAIL.n76 VTAIL.n75 9.3005
R450 VTAIL.n83 VTAIL.n82 9.3005
R451 VTAIL.n85 VTAIL.n84 9.3005
R452 VTAIL.n72 VTAIL.n71 9.3005
R453 VTAIL.n91 VTAIL.n90 9.3005
R454 VTAIL.n93 VTAIL.n92 9.3005
R455 VTAIL.n67 VTAIL.n65 9.3005
R456 VTAIL.n99 VTAIL.n98 9.3005
R457 VTAIL.n107 VTAIL.n106 9.3005
R458 VTAIL.n62 VTAIL.n61 9.3005
R459 VTAIL.n101 VTAIL.n100 9.3005
R460 VTAIL.n187 VTAIL.n176 8.92171
R461 VTAIL.n25 VTAIL.n14 8.92171
R462 VTAIL.n139 VTAIL.n128 8.92171
R463 VTAIL.n85 VTAIL.n74 8.92171
R464 VTAIL.n184 VTAIL.n183 8.14595
R465 VTAIL.n22 VTAIL.n21 8.14595
R466 VTAIL.n136 VTAIL.n135 8.14595
R467 VTAIL.n82 VTAIL.n81 8.14595
R468 VTAIL.n180 VTAIL.n178 7.3702
R469 VTAIL.n18 VTAIL.n16 7.3702
R470 VTAIL.n132 VTAIL.n130 7.3702
R471 VTAIL.n78 VTAIL.n76 7.3702
R472 VTAIL.n183 VTAIL.n178 5.81868
R473 VTAIL.n21 VTAIL.n16 5.81868
R474 VTAIL.n135 VTAIL.n130 5.81868
R475 VTAIL.n81 VTAIL.n76 5.81868
R476 VTAIL.n184 VTAIL.n176 5.04292
R477 VTAIL.n22 VTAIL.n14 5.04292
R478 VTAIL.n136 VTAIL.n128 5.04292
R479 VTAIL.n82 VTAIL.n74 5.04292
R480 VTAIL.n188 VTAIL.n187 4.26717
R481 VTAIL.n26 VTAIL.n25 4.26717
R482 VTAIL.n140 VTAIL.n139 4.26717
R483 VTAIL.n86 VTAIL.n85 4.26717
R484 VTAIL.n191 VTAIL.n174 3.49141
R485 VTAIL.n29 VTAIL.n12 3.49141
R486 VTAIL.n143 VTAIL.n126 3.49141
R487 VTAIL.n89 VTAIL.n72 3.49141
R488 VTAIL.n214 VTAIL.t14 3.45114
R489 VTAIL.n214 VTAIL.t18 3.45114
R490 VTAIL.n0 VTAIL.t12 3.45114
R491 VTAIL.n0 VTAIL.t9 3.45114
R492 VTAIL.n52 VTAIL.t5 3.45114
R493 VTAIL.n52 VTAIL.t19 3.45114
R494 VTAIL.n54 VTAIL.t8 3.45114
R495 VTAIL.n54 VTAIL.t2 3.45114
R496 VTAIL.n112 VTAIL.t1 3.45114
R497 VTAIL.n112 VTAIL.t0 3.45114
R498 VTAIL.n110 VTAIL.t3 3.45114
R499 VTAIL.n110 VTAIL.t7 3.45114
R500 VTAIL.n58 VTAIL.t10 3.45114
R501 VTAIL.n58 VTAIL.t17 3.45114
R502 VTAIL.n56 VTAIL.t15 3.45114
R503 VTAIL.n56 VTAIL.t11 3.45114
R504 VTAIL.n192 VTAIL.n172 2.71565
R505 VTAIL.n212 VTAIL.n164 2.71565
R506 VTAIL.n30 VTAIL.n10 2.71565
R507 VTAIL.n50 VTAIL.n2 2.71565
R508 VTAIL.n162 VTAIL.n114 2.71565
R509 VTAIL.n144 VTAIL.n124 2.71565
R510 VTAIL.n108 VTAIL.n60 2.71565
R511 VTAIL.n90 VTAIL.n70 2.71565
R512 VTAIL.n179 VTAIL.n177 2.41283
R513 VTAIL.n17 VTAIL.n15 2.41283
R514 VTAIL.n131 VTAIL.n129 2.41283
R515 VTAIL.n77 VTAIL.n75 2.41283
R516 VTAIL.n197 VTAIL.n195 1.93989
R517 VTAIL.n210 VTAIL.n209 1.93989
R518 VTAIL.n35 VTAIL.n33 1.93989
R519 VTAIL.n48 VTAIL.n47 1.93989
R520 VTAIL.n160 VTAIL.n159 1.93989
R521 VTAIL.n148 VTAIL.n147 1.93989
R522 VTAIL.n106 VTAIL.n105 1.93989
R523 VTAIL.n94 VTAIL.n93 1.93989
R524 VTAIL.n59 VTAIL.n57 1.55222
R525 VTAIL.n109 VTAIL.n59 1.55222
R526 VTAIL.n113 VTAIL.n111 1.55222
R527 VTAIL.n163 VTAIL.n113 1.55222
R528 VTAIL.n55 VTAIL.n53 1.55222
R529 VTAIL.n53 VTAIL.n51 1.55222
R530 VTAIL.n215 VTAIL.n213 1.55222
R531 VTAIL.n111 VTAIL.n109 1.24619
R532 VTAIL.n51 VTAIL.n1 1.24619
R533 VTAIL VTAIL.n1 1.22248
R534 VTAIL.n196 VTAIL.n170 1.16414
R535 VTAIL.n206 VTAIL.n166 1.16414
R536 VTAIL.n34 VTAIL.n8 1.16414
R537 VTAIL.n44 VTAIL.n4 1.16414
R538 VTAIL.n156 VTAIL.n116 1.16414
R539 VTAIL.n151 VTAIL.n121 1.16414
R540 VTAIL.n102 VTAIL.n62 1.16414
R541 VTAIL.n97 VTAIL.n67 1.16414
R542 VTAIL.n202 VTAIL.n201 0.388379
R543 VTAIL.n205 VTAIL.n168 0.388379
R544 VTAIL.n40 VTAIL.n39 0.388379
R545 VTAIL.n43 VTAIL.n6 0.388379
R546 VTAIL.n155 VTAIL.n118 0.388379
R547 VTAIL.n152 VTAIL.n120 0.388379
R548 VTAIL.n101 VTAIL.n64 0.388379
R549 VTAIL.n98 VTAIL.n66 0.388379
R550 VTAIL VTAIL.n215 0.330241
R551 VTAIL.n185 VTAIL.n177 0.155672
R552 VTAIL.n186 VTAIL.n185 0.155672
R553 VTAIL.n186 VTAIL.n173 0.155672
R554 VTAIL.n193 VTAIL.n173 0.155672
R555 VTAIL.n194 VTAIL.n193 0.155672
R556 VTAIL.n194 VTAIL.n169 0.155672
R557 VTAIL.n203 VTAIL.n169 0.155672
R558 VTAIL.n204 VTAIL.n203 0.155672
R559 VTAIL.n204 VTAIL.n165 0.155672
R560 VTAIL.n211 VTAIL.n165 0.155672
R561 VTAIL.n23 VTAIL.n15 0.155672
R562 VTAIL.n24 VTAIL.n23 0.155672
R563 VTAIL.n24 VTAIL.n11 0.155672
R564 VTAIL.n31 VTAIL.n11 0.155672
R565 VTAIL.n32 VTAIL.n31 0.155672
R566 VTAIL.n32 VTAIL.n7 0.155672
R567 VTAIL.n41 VTAIL.n7 0.155672
R568 VTAIL.n42 VTAIL.n41 0.155672
R569 VTAIL.n42 VTAIL.n3 0.155672
R570 VTAIL.n49 VTAIL.n3 0.155672
R571 VTAIL.n161 VTAIL.n115 0.155672
R572 VTAIL.n154 VTAIL.n115 0.155672
R573 VTAIL.n154 VTAIL.n153 0.155672
R574 VTAIL.n153 VTAIL.n119 0.155672
R575 VTAIL.n146 VTAIL.n119 0.155672
R576 VTAIL.n146 VTAIL.n145 0.155672
R577 VTAIL.n145 VTAIL.n125 0.155672
R578 VTAIL.n138 VTAIL.n125 0.155672
R579 VTAIL.n138 VTAIL.n137 0.155672
R580 VTAIL.n137 VTAIL.n129 0.155672
R581 VTAIL.n107 VTAIL.n61 0.155672
R582 VTAIL.n100 VTAIL.n61 0.155672
R583 VTAIL.n100 VTAIL.n99 0.155672
R584 VTAIL.n99 VTAIL.n65 0.155672
R585 VTAIL.n92 VTAIL.n65 0.155672
R586 VTAIL.n92 VTAIL.n91 0.155672
R587 VTAIL.n91 VTAIL.n71 0.155672
R588 VTAIL.n84 VTAIL.n71 0.155672
R589 VTAIL.n84 VTAIL.n83 0.155672
R590 VTAIL.n83 VTAIL.n75 0.155672
R591 VP.n15 VP.t4 185.481
R592 VP.n36 VP.n35 180.974
R593 VP.n62 VP.n61 180.974
R594 VP.n34 VP.n33 180.974
R595 VP.n16 VP.n13 161.3
R596 VP.n18 VP.n17 161.3
R597 VP.n19 VP.n12 161.3
R598 VP.n21 VP.n20 161.3
R599 VP.n22 VP.n11 161.3
R600 VP.n24 VP.n23 161.3
R601 VP.n25 VP.n10 161.3
R602 VP.n28 VP.n27 161.3
R603 VP.n29 VP.n9 161.3
R604 VP.n31 VP.n30 161.3
R605 VP.n32 VP.n8 161.3
R606 VP.n60 VP.n0 161.3
R607 VP.n59 VP.n58 161.3
R608 VP.n57 VP.n1 161.3
R609 VP.n56 VP.n55 161.3
R610 VP.n53 VP.n2 161.3
R611 VP.n52 VP.n51 161.3
R612 VP.n50 VP.n3 161.3
R613 VP.n49 VP.n48 161.3
R614 VP.n47 VP.n4 161.3
R615 VP.n46 VP.n45 161.3
R616 VP.n44 VP.n5 161.3
R617 VP.n43 VP.n42 161.3
R618 VP.n40 VP.n6 161.3
R619 VP.n39 VP.n38 161.3
R620 VP.n37 VP.n7 161.3
R621 VP.n48 VP.t3 154.438
R622 VP.n35 VP.t0 154.438
R623 VP.n41 VP.t8 154.438
R624 VP.n54 VP.t1 154.438
R625 VP.n61 VP.t5 154.438
R626 VP.n20 VP.t7 154.438
R627 VP.n33 VP.t2 154.438
R628 VP.n26 VP.t6 154.438
R629 VP.n14 VP.t9 154.438
R630 VP.n40 VP.n39 56.5617
R631 VP.n59 VP.n1 56.5617
R632 VP.n31 VP.n9 56.5617
R633 VP.n15 VP.n14 51.3232
R634 VP.n47 VP.n46 50.2647
R635 VP.n52 VP.n3 50.2647
R636 VP.n24 VP.n11 50.2647
R637 VP.n19 VP.n18 50.2647
R638 VP.n36 VP.n34 44.8566
R639 VP.n46 VP.n5 30.8893
R640 VP.n53 VP.n52 30.8893
R641 VP.n25 VP.n24 30.8893
R642 VP.n18 VP.n13 30.8893
R643 VP.n39 VP.n7 24.5923
R644 VP.n42 VP.n40 24.5923
R645 VP.n48 VP.n47 24.5923
R646 VP.n48 VP.n3 24.5923
R647 VP.n55 VP.n1 24.5923
R648 VP.n60 VP.n59 24.5923
R649 VP.n32 VP.n31 24.5923
R650 VP.n27 VP.n9 24.5923
R651 VP.n20 VP.n19 24.5923
R652 VP.n20 VP.n11 24.5923
R653 VP.n16 VP.n15 18.2653
R654 VP.n41 VP.n5 14.7556
R655 VP.n54 VP.n53 14.7556
R656 VP.n26 VP.n25 14.7556
R657 VP.n14 VP.n13 14.7556
R658 VP.n42 VP.n41 9.83723
R659 VP.n55 VP.n54 9.83723
R660 VP.n27 VP.n26 9.83723
R661 VP.n35 VP.n7 4.91887
R662 VP.n61 VP.n60 4.91887
R663 VP.n33 VP.n32 4.91887
R664 VP.n17 VP.n16 0.189894
R665 VP.n17 VP.n12 0.189894
R666 VP.n21 VP.n12 0.189894
R667 VP.n22 VP.n21 0.189894
R668 VP.n23 VP.n22 0.189894
R669 VP.n23 VP.n10 0.189894
R670 VP.n28 VP.n10 0.189894
R671 VP.n29 VP.n28 0.189894
R672 VP.n30 VP.n29 0.189894
R673 VP.n30 VP.n8 0.189894
R674 VP.n34 VP.n8 0.189894
R675 VP.n37 VP.n36 0.189894
R676 VP.n38 VP.n37 0.189894
R677 VP.n38 VP.n6 0.189894
R678 VP.n43 VP.n6 0.189894
R679 VP.n44 VP.n43 0.189894
R680 VP.n45 VP.n44 0.189894
R681 VP.n45 VP.n4 0.189894
R682 VP.n49 VP.n4 0.189894
R683 VP.n50 VP.n49 0.189894
R684 VP.n51 VP.n50 0.189894
R685 VP.n51 VP.n2 0.189894
R686 VP.n56 VP.n2 0.189894
R687 VP.n57 VP.n56 0.189894
R688 VP.n58 VP.n57 0.189894
R689 VP.n58 VP.n0 0.189894
R690 VP.n62 VP.n0 0.189894
R691 VP VP.n62 0.0516364
R692 VDD1.n44 VDD1.n0 756.745
R693 VDD1.n95 VDD1.n51 756.745
R694 VDD1.n45 VDD1.n44 585
R695 VDD1.n43 VDD1.n42 585
R696 VDD1.n4 VDD1.n3 585
R697 VDD1.n8 VDD1.n6 585
R698 VDD1.n37 VDD1.n36 585
R699 VDD1.n35 VDD1.n34 585
R700 VDD1.n10 VDD1.n9 585
R701 VDD1.n29 VDD1.n28 585
R702 VDD1.n27 VDD1.n26 585
R703 VDD1.n14 VDD1.n13 585
R704 VDD1.n21 VDD1.n20 585
R705 VDD1.n19 VDD1.n18 585
R706 VDD1.n68 VDD1.n67 585
R707 VDD1.n70 VDD1.n69 585
R708 VDD1.n63 VDD1.n62 585
R709 VDD1.n76 VDD1.n75 585
R710 VDD1.n78 VDD1.n77 585
R711 VDD1.n59 VDD1.n58 585
R712 VDD1.n85 VDD1.n84 585
R713 VDD1.n86 VDD1.n57 585
R714 VDD1.n88 VDD1.n87 585
R715 VDD1.n55 VDD1.n54 585
R716 VDD1.n94 VDD1.n93 585
R717 VDD1.n96 VDD1.n95 585
R718 VDD1.n17 VDD1.t5 329.038
R719 VDD1.n66 VDD1.t9 329.038
R720 VDD1.n44 VDD1.n43 171.744
R721 VDD1.n43 VDD1.n3 171.744
R722 VDD1.n8 VDD1.n3 171.744
R723 VDD1.n36 VDD1.n8 171.744
R724 VDD1.n36 VDD1.n35 171.744
R725 VDD1.n35 VDD1.n9 171.744
R726 VDD1.n28 VDD1.n9 171.744
R727 VDD1.n28 VDD1.n27 171.744
R728 VDD1.n27 VDD1.n13 171.744
R729 VDD1.n20 VDD1.n13 171.744
R730 VDD1.n20 VDD1.n19 171.744
R731 VDD1.n69 VDD1.n68 171.744
R732 VDD1.n69 VDD1.n62 171.744
R733 VDD1.n76 VDD1.n62 171.744
R734 VDD1.n77 VDD1.n76 171.744
R735 VDD1.n77 VDD1.n58 171.744
R736 VDD1.n85 VDD1.n58 171.744
R737 VDD1.n86 VDD1.n85 171.744
R738 VDD1.n87 VDD1.n86 171.744
R739 VDD1.n87 VDD1.n54 171.744
R740 VDD1.n94 VDD1.n54 171.744
R741 VDD1.n95 VDD1.n94 171.744
R742 VDD1.n19 VDD1.t5 85.8723
R743 VDD1.n68 VDD1.t9 85.8723
R744 VDD1.n103 VDD1.n102 83.1801
R745 VDD1.n50 VDD1.n49 82.0718
R746 VDD1.n101 VDD1.n100 82.0716
R747 VDD1.n105 VDD1.n104 82.0716
R748 VDD1.n50 VDD1.n48 53.9068
R749 VDD1.n101 VDD1.n99 53.9068
R750 VDD1.n105 VDD1.n103 40.5656
R751 VDD1.n6 VDD1.n4 13.1884
R752 VDD1.n88 VDD1.n55 13.1884
R753 VDD1.n42 VDD1.n41 12.8005
R754 VDD1.n38 VDD1.n37 12.8005
R755 VDD1.n89 VDD1.n57 12.8005
R756 VDD1.n93 VDD1.n92 12.8005
R757 VDD1.n45 VDD1.n2 12.0247
R758 VDD1.n34 VDD1.n7 12.0247
R759 VDD1.n84 VDD1.n83 12.0247
R760 VDD1.n96 VDD1.n53 12.0247
R761 VDD1.n46 VDD1.n0 11.249
R762 VDD1.n33 VDD1.n10 11.249
R763 VDD1.n82 VDD1.n59 11.249
R764 VDD1.n97 VDD1.n51 11.249
R765 VDD1.n18 VDD1.n17 10.7239
R766 VDD1.n67 VDD1.n66 10.7239
R767 VDD1.n30 VDD1.n29 10.4732
R768 VDD1.n79 VDD1.n78 10.4732
R769 VDD1.n26 VDD1.n12 9.69747
R770 VDD1.n75 VDD1.n61 9.69747
R771 VDD1.n48 VDD1.n47 9.45567
R772 VDD1.n99 VDD1.n98 9.45567
R773 VDD1.n16 VDD1.n15 9.3005
R774 VDD1.n23 VDD1.n22 9.3005
R775 VDD1.n25 VDD1.n24 9.3005
R776 VDD1.n12 VDD1.n11 9.3005
R777 VDD1.n31 VDD1.n30 9.3005
R778 VDD1.n33 VDD1.n32 9.3005
R779 VDD1.n7 VDD1.n5 9.3005
R780 VDD1.n39 VDD1.n38 9.3005
R781 VDD1.n47 VDD1.n46 9.3005
R782 VDD1.n2 VDD1.n1 9.3005
R783 VDD1.n41 VDD1.n40 9.3005
R784 VDD1.n98 VDD1.n97 9.3005
R785 VDD1.n53 VDD1.n52 9.3005
R786 VDD1.n92 VDD1.n91 9.3005
R787 VDD1.n65 VDD1.n64 9.3005
R788 VDD1.n72 VDD1.n71 9.3005
R789 VDD1.n74 VDD1.n73 9.3005
R790 VDD1.n61 VDD1.n60 9.3005
R791 VDD1.n80 VDD1.n79 9.3005
R792 VDD1.n82 VDD1.n81 9.3005
R793 VDD1.n83 VDD1.n56 9.3005
R794 VDD1.n90 VDD1.n89 9.3005
R795 VDD1.n25 VDD1.n14 8.92171
R796 VDD1.n74 VDD1.n63 8.92171
R797 VDD1.n22 VDD1.n21 8.14595
R798 VDD1.n71 VDD1.n70 8.14595
R799 VDD1.n18 VDD1.n16 7.3702
R800 VDD1.n67 VDD1.n65 7.3702
R801 VDD1.n21 VDD1.n16 5.81868
R802 VDD1.n70 VDD1.n65 5.81868
R803 VDD1.n22 VDD1.n14 5.04292
R804 VDD1.n71 VDD1.n63 5.04292
R805 VDD1.n26 VDD1.n25 4.26717
R806 VDD1.n75 VDD1.n74 4.26717
R807 VDD1.n29 VDD1.n12 3.49141
R808 VDD1.n78 VDD1.n61 3.49141
R809 VDD1.n104 VDD1.t3 3.45114
R810 VDD1.n104 VDD1.t7 3.45114
R811 VDD1.n49 VDD1.t0 3.45114
R812 VDD1.n49 VDD1.t2 3.45114
R813 VDD1.n102 VDD1.t8 3.45114
R814 VDD1.n102 VDD1.t4 3.45114
R815 VDD1.n100 VDD1.t1 3.45114
R816 VDD1.n100 VDD1.t6 3.45114
R817 VDD1.n48 VDD1.n0 2.71565
R818 VDD1.n30 VDD1.n10 2.71565
R819 VDD1.n79 VDD1.n59 2.71565
R820 VDD1.n99 VDD1.n51 2.71565
R821 VDD1.n17 VDD1.n15 2.41283
R822 VDD1.n66 VDD1.n64 2.41283
R823 VDD1.n46 VDD1.n45 1.93989
R824 VDD1.n34 VDD1.n33 1.93989
R825 VDD1.n84 VDD1.n82 1.93989
R826 VDD1.n97 VDD1.n96 1.93989
R827 VDD1.n42 VDD1.n2 1.16414
R828 VDD1.n37 VDD1.n7 1.16414
R829 VDD1.n83 VDD1.n57 1.16414
R830 VDD1.n93 VDD1.n53 1.16414
R831 VDD1 VDD1.n105 1.1061
R832 VDD1 VDD1.n50 0.446621
R833 VDD1.n41 VDD1.n4 0.388379
R834 VDD1.n38 VDD1.n6 0.388379
R835 VDD1.n89 VDD1.n88 0.388379
R836 VDD1.n92 VDD1.n55 0.388379
R837 VDD1.n103 VDD1.n101 0.333085
R838 VDD1.n47 VDD1.n1 0.155672
R839 VDD1.n40 VDD1.n1 0.155672
R840 VDD1.n40 VDD1.n39 0.155672
R841 VDD1.n39 VDD1.n5 0.155672
R842 VDD1.n32 VDD1.n5 0.155672
R843 VDD1.n32 VDD1.n31 0.155672
R844 VDD1.n31 VDD1.n11 0.155672
R845 VDD1.n24 VDD1.n11 0.155672
R846 VDD1.n24 VDD1.n23 0.155672
R847 VDD1.n23 VDD1.n15 0.155672
R848 VDD1.n72 VDD1.n64 0.155672
R849 VDD1.n73 VDD1.n72 0.155672
R850 VDD1.n73 VDD1.n60 0.155672
R851 VDD1.n80 VDD1.n60 0.155672
R852 VDD1.n81 VDD1.n80 0.155672
R853 VDD1.n81 VDD1.n56 0.155672
R854 VDD1.n90 VDD1.n56 0.155672
R855 VDD1.n91 VDD1.n90 0.155672
R856 VDD1.n91 VDD1.n52 0.155672
R857 VDD1.n98 VDD1.n52 0.155672
R858 B.n468 B.n65 585
R859 B.n470 B.n469 585
R860 B.n471 B.n64 585
R861 B.n473 B.n472 585
R862 B.n474 B.n63 585
R863 B.n476 B.n475 585
R864 B.n477 B.n62 585
R865 B.n479 B.n478 585
R866 B.n480 B.n61 585
R867 B.n482 B.n481 585
R868 B.n483 B.n60 585
R869 B.n485 B.n484 585
R870 B.n486 B.n59 585
R871 B.n488 B.n487 585
R872 B.n489 B.n58 585
R873 B.n491 B.n490 585
R874 B.n492 B.n57 585
R875 B.n494 B.n493 585
R876 B.n495 B.n56 585
R877 B.n497 B.n496 585
R878 B.n498 B.n55 585
R879 B.n500 B.n499 585
R880 B.n501 B.n54 585
R881 B.n503 B.n502 585
R882 B.n504 B.n53 585
R883 B.n506 B.n505 585
R884 B.n507 B.n52 585
R885 B.n509 B.n508 585
R886 B.n510 B.n51 585
R887 B.n512 B.n511 585
R888 B.n513 B.n50 585
R889 B.n515 B.n514 585
R890 B.n516 B.n49 585
R891 B.n518 B.n517 585
R892 B.n520 B.n519 585
R893 B.n521 B.n45 585
R894 B.n523 B.n522 585
R895 B.n524 B.n44 585
R896 B.n526 B.n525 585
R897 B.n527 B.n43 585
R898 B.n529 B.n528 585
R899 B.n530 B.n42 585
R900 B.n532 B.n531 585
R901 B.n533 B.n39 585
R902 B.n536 B.n535 585
R903 B.n537 B.n38 585
R904 B.n539 B.n538 585
R905 B.n540 B.n37 585
R906 B.n542 B.n541 585
R907 B.n543 B.n36 585
R908 B.n545 B.n544 585
R909 B.n546 B.n35 585
R910 B.n548 B.n547 585
R911 B.n549 B.n34 585
R912 B.n551 B.n550 585
R913 B.n552 B.n33 585
R914 B.n554 B.n553 585
R915 B.n555 B.n32 585
R916 B.n557 B.n556 585
R917 B.n558 B.n31 585
R918 B.n560 B.n559 585
R919 B.n561 B.n30 585
R920 B.n563 B.n562 585
R921 B.n564 B.n29 585
R922 B.n566 B.n565 585
R923 B.n567 B.n28 585
R924 B.n569 B.n568 585
R925 B.n570 B.n27 585
R926 B.n572 B.n571 585
R927 B.n573 B.n26 585
R928 B.n575 B.n574 585
R929 B.n576 B.n25 585
R930 B.n578 B.n577 585
R931 B.n579 B.n24 585
R932 B.n581 B.n580 585
R933 B.n582 B.n23 585
R934 B.n584 B.n583 585
R935 B.n585 B.n22 585
R936 B.n467 B.n466 585
R937 B.n465 B.n66 585
R938 B.n464 B.n463 585
R939 B.n462 B.n67 585
R940 B.n461 B.n460 585
R941 B.n459 B.n68 585
R942 B.n458 B.n457 585
R943 B.n456 B.n69 585
R944 B.n455 B.n454 585
R945 B.n453 B.n70 585
R946 B.n452 B.n451 585
R947 B.n450 B.n71 585
R948 B.n449 B.n448 585
R949 B.n447 B.n72 585
R950 B.n446 B.n445 585
R951 B.n444 B.n73 585
R952 B.n443 B.n442 585
R953 B.n441 B.n74 585
R954 B.n440 B.n439 585
R955 B.n438 B.n75 585
R956 B.n437 B.n436 585
R957 B.n435 B.n76 585
R958 B.n434 B.n433 585
R959 B.n432 B.n77 585
R960 B.n431 B.n430 585
R961 B.n429 B.n78 585
R962 B.n428 B.n427 585
R963 B.n426 B.n79 585
R964 B.n425 B.n424 585
R965 B.n423 B.n80 585
R966 B.n422 B.n421 585
R967 B.n420 B.n81 585
R968 B.n419 B.n418 585
R969 B.n417 B.n82 585
R970 B.n416 B.n415 585
R971 B.n414 B.n83 585
R972 B.n413 B.n412 585
R973 B.n411 B.n84 585
R974 B.n410 B.n409 585
R975 B.n408 B.n85 585
R976 B.n407 B.n406 585
R977 B.n405 B.n86 585
R978 B.n404 B.n403 585
R979 B.n402 B.n87 585
R980 B.n401 B.n400 585
R981 B.n399 B.n88 585
R982 B.n398 B.n397 585
R983 B.n396 B.n89 585
R984 B.n395 B.n394 585
R985 B.n393 B.n90 585
R986 B.n392 B.n391 585
R987 B.n390 B.n91 585
R988 B.n389 B.n388 585
R989 B.n387 B.n92 585
R990 B.n386 B.n385 585
R991 B.n384 B.n93 585
R992 B.n383 B.n382 585
R993 B.n381 B.n94 585
R994 B.n380 B.n379 585
R995 B.n378 B.n95 585
R996 B.n377 B.n376 585
R997 B.n375 B.n96 585
R998 B.n374 B.n373 585
R999 B.n372 B.n97 585
R1000 B.n371 B.n370 585
R1001 B.n369 B.n98 585
R1002 B.n368 B.n367 585
R1003 B.n366 B.n99 585
R1004 B.n365 B.n364 585
R1005 B.n363 B.n100 585
R1006 B.n362 B.n361 585
R1007 B.n360 B.n101 585
R1008 B.n359 B.n358 585
R1009 B.n357 B.n102 585
R1010 B.n356 B.n355 585
R1011 B.n354 B.n103 585
R1012 B.n353 B.n352 585
R1013 B.n351 B.n104 585
R1014 B.n350 B.n349 585
R1015 B.n348 B.n105 585
R1016 B.n347 B.n346 585
R1017 B.n228 B.n149 585
R1018 B.n230 B.n229 585
R1019 B.n231 B.n148 585
R1020 B.n233 B.n232 585
R1021 B.n234 B.n147 585
R1022 B.n236 B.n235 585
R1023 B.n237 B.n146 585
R1024 B.n239 B.n238 585
R1025 B.n240 B.n145 585
R1026 B.n242 B.n241 585
R1027 B.n243 B.n144 585
R1028 B.n245 B.n244 585
R1029 B.n246 B.n143 585
R1030 B.n248 B.n247 585
R1031 B.n249 B.n142 585
R1032 B.n251 B.n250 585
R1033 B.n252 B.n141 585
R1034 B.n254 B.n253 585
R1035 B.n255 B.n140 585
R1036 B.n257 B.n256 585
R1037 B.n258 B.n139 585
R1038 B.n260 B.n259 585
R1039 B.n261 B.n138 585
R1040 B.n263 B.n262 585
R1041 B.n264 B.n137 585
R1042 B.n266 B.n265 585
R1043 B.n267 B.n136 585
R1044 B.n269 B.n268 585
R1045 B.n270 B.n135 585
R1046 B.n272 B.n271 585
R1047 B.n273 B.n134 585
R1048 B.n275 B.n274 585
R1049 B.n276 B.n133 585
R1050 B.n278 B.n277 585
R1051 B.n280 B.n279 585
R1052 B.n281 B.n129 585
R1053 B.n283 B.n282 585
R1054 B.n284 B.n128 585
R1055 B.n286 B.n285 585
R1056 B.n287 B.n127 585
R1057 B.n289 B.n288 585
R1058 B.n290 B.n126 585
R1059 B.n292 B.n291 585
R1060 B.n293 B.n123 585
R1061 B.n296 B.n295 585
R1062 B.n297 B.n122 585
R1063 B.n299 B.n298 585
R1064 B.n300 B.n121 585
R1065 B.n302 B.n301 585
R1066 B.n303 B.n120 585
R1067 B.n305 B.n304 585
R1068 B.n306 B.n119 585
R1069 B.n308 B.n307 585
R1070 B.n309 B.n118 585
R1071 B.n311 B.n310 585
R1072 B.n312 B.n117 585
R1073 B.n314 B.n313 585
R1074 B.n315 B.n116 585
R1075 B.n317 B.n316 585
R1076 B.n318 B.n115 585
R1077 B.n320 B.n319 585
R1078 B.n321 B.n114 585
R1079 B.n323 B.n322 585
R1080 B.n324 B.n113 585
R1081 B.n326 B.n325 585
R1082 B.n327 B.n112 585
R1083 B.n329 B.n328 585
R1084 B.n330 B.n111 585
R1085 B.n332 B.n331 585
R1086 B.n333 B.n110 585
R1087 B.n335 B.n334 585
R1088 B.n336 B.n109 585
R1089 B.n338 B.n337 585
R1090 B.n339 B.n108 585
R1091 B.n341 B.n340 585
R1092 B.n342 B.n107 585
R1093 B.n344 B.n343 585
R1094 B.n345 B.n106 585
R1095 B.n227 B.n226 585
R1096 B.n225 B.n150 585
R1097 B.n224 B.n223 585
R1098 B.n222 B.n151 585
R1099 B.n221 B.n220 585
R1100 B.n219 B.n152 585
R1101 B.n218 B.n217 585
R1102 B.n216 B.n153 585
R1103 B.n215 B.n214 585
R1104 B.n213 B.n154 585
R1105 B.n212 B.n211 585
R1106 B.n210 B.n155 585
R1107 B.n209 B.n208 585
R1108 B.n207 B.n156 585
R1109 B.n206 B.n205 585
R1110 B.n204 B.n157 585
R1111 B.n203 B.n202 585
R1112 B.n201 B.n158 585
R1113 B.n200 B.n199 585
R1114 B.n198 B.n159 585
R1115 B.n197 B.n196 585
R1116 B.n195 B.n160 585
R1117 B.n194 B.n193 585
R1118 B.n192 B.n161 585
R1119 B.n191 B.n190 585
R1120 B.n189 B.n162 585
R1121 B.n188 B.n187 585
R1122 B.n186 B.n163 585
R1123 B.n185 B.n184 585
R1124 B.n183 B.n164 585
R1125 B.n182 B.n181 585
R1126 B.n180 B.n165 585
R1127 B.n179 B.n178 585
R1128 B.n177 B.n166 585
R1129 B.n176 B.n175 585
R1130 B.n174 B.n167 585
R1131 B.n173 B.n172 585
R1132 B.n171 B.n168 585
R1133 B.n170 B.n169 585
R1134 B.n2 B.n0 585
R1135 B.n645 B.n1 585
R1136 B.n644 B.n643 585
R1137 B.n642 B.n3 585
R1138 B.n641 B.n640 585
R1139 B.n639 B.n4 585
R1140 B.n638 B.n637 585
R1141 B.n636 B.n5 585
R1142 B.n635 B.n634 585
R1143 B.n633 B.n6 585
R1144 B.n632 B.n631 585
R1145 B.n630 B.n7 585
R1146 B.n629 B.n628 585
R1147 B.n627 B.n8 585
R1148 B.n626 B.n625 585
R1149 B.n624 B.n9 585
R1150 B.n623 B.n622 585
R1151 B.n621 B.n10 585
R1152 B.n620 B.n619 585
R1153 B.n618 B.n11 585
R1154 B.n617 B.n616 585
R1155 B.n615 B.n12 585
R1156 B.n614 B.n613 585
R1157 B.n612 B.n13 585
R1158 B.n611 B.n610 585
R1159 B.n609 B.n14 585
R1160 B.n608 B.n607 585
R1161 B.n606 B.n15 585
R1162 B.n605 B.n604 585
R1163 B.n603 B.n16 585
R1164 B.n602 B.n601 585
R1165 B.n600 B.n17 585
R1166 B.n599 B.n598 585
R1167 B.n597 B.n18 585
R1168 B.n596 B.n595 585
R1169 B.n594 B.n19 585
R1170 B.n593 B.n592 585
R1171 B.n591 B.n20 585
R1172 B.n590 B.n589 585
R1173 B.n588 B.n21 585
R1174 B.n587 B.n586 585
R1175 B.n647 B.n646 585
R1176 B.n226 B.n149 449.257
R1177 B.n586 B.n585 449.257
R1178 B.n346 B.n345 449.257
R1179 B.n466 B.n65 449.257
R1180 B.n124 B.t5 364.19
R1181 B.n46 B.t1 364.19
R1182 B.n130 B.t8 364.19
R1183 B.n40 B.t10 364.19
R1184 B.n124 B.t3 359.764
R1185 B.n130 B.t6 359.764
R1186 B.n40 B.t9 359.764
R1187 B.n46 B.t0 359.764
R1188 B.n125 B.t4 329.281
R1189 B.n47 B.t2 329.281
R1190 B.n131 B.t7 329.281
R1191 B.n41 B.t11 329.281
R1192 B.n226 B.n225 163.367
R1193 B.n225 B.n224 163.367
R1194 B.n224 B.n151 163.367
R1195 B.n220 B.n151 163.367
R1196 B.n220 B.n219 163.367
R1197 B.n219 B.n218 163.367
R1198 B.n218 B.n153 163.367
R1199 B.n214 B.n153 163.367
R1200 B.n214 B.n213 163.367
R1201 B.n213 B.n212 163.367
R1202 B.n212 B.n155 163.367
R1203 B.n208 B.n155 163.367
R1204 B.n208 B.n207 163.367
R1205 B.n207 B.n206 163.367
R1206 B.n206 B.n157 163.367
R1207 B.n202 B.n157 163.367
R1208 B.n202 B.n201 163.367
R1209 B.n201 B.n200 163.367
R1210 B.n200 B.n159 163.367
R1211 B.n196 B.n159 163.367
R1212 B.n196 B.n195 163.367
R1213 B.n195 B.n194 163.367
R1214 B.n194 B.n161 163.367
R1215 B.n190 B.n161 163.367
R1216 B.n190 B.n189 163.367
R1217 B.n189 B.n188 163.367
R1218 B.n188 B.n163 163.367
R1219 B.n184 B.n163 163.367
R1220 B.n184 B.n183 163.367
R1221 B.n183 B.n182 163.367
R1222 B.n182 B.n165 163.367
R1223 B.n178 B.n165 163.367
R1224 B.n178 B.n177 163.367
R1225 B.n177 B.n176 163.367
R1226 B.n176 B.n167 163.367
R1227 B.n172 B.n167 163.367
R1228 B.n172 B.n171 163.367
R1229 B.n171 B.n170 163.367
R1230 B.n170 B.n2 163.367
R1231 B.n646 B.n2 163.367
R1232 B.n646 B.n645 163.367
R1233 B.n645 B.n644 163.367
R1234 B.n644 B.n3 163.367
R1235 B.n640 B.n3 163.367
R1236 B.n640 B.n639 163.367
R1237 B.n639 B.n638 163.367
R1238 B.n638 B.n5 163.367
R1239 B.n634 B.n5 163.367
R1240 B.n634 B.n633 163.367
R1241 B.n633 B.n632 163.367
R1242 B.n632 B.n7 163.367
R1243 B.n628 B.n7 163.367
R1244 B.n628 B.n627 163.367
R1245 B.n627 B.n626 163.367
R1246 B.n626 B.n9 163.367
R1247 B.n622 B.n9 163.367
R1248 B.n622 B.n621 163.367
R1249 B.n621 B.n620 163.367
R1250 B.n620 B.n11 163.367
R1251 B.n616 B.n11 163.367
R1252 B.n616 B.n615 163.367
R1253 B.n615 B.n614 163.367
R1254 B.n614 B.n13 163.367
R1255 B.n610 B.n13 163.367
R1256 B.n610 B.n609 163.367
R1257 B.n609 B.n608 163.367
R1258 B.n608 B.n15 163.367
R1259 B.n604 B.n15 163.367
R1260 B.n604 B.n603 163.367
R1261 B.n603 B.n602 163.367
R1262 B.n602 B.n17 163.367
R1263 B.n598 B.n17 163.367
R1264 B.n598 B.n597 163.367
R1265 B.n597 B.n596 163.367
R1266 B.n596 B.n19 163.367
R1267 B.n592 B.n19 163.367
R1268 B.n592 B.n591 163.367
R1269 B.n591 B.n590 163.367
R1270 B.n590 B.n21 163.367
R1271 B.n586 B.n21 163.367
R1272 B.n230 B.n149 163.367
R1273 B.n231 B.n230 163.367
R1274 B.n232 B.n231 163.367
R1275 B.n232 B.n147 163.367
R1276 B.n236 B.n147 163.367
R1277 B.n237 B.n236 163.367
R1278 B.n238 B.n237 163.367
R1279 B.n238 B.n145 163.367
R1280 B.n242 B.n145 163.367
R1281 B.n243 B.n242 163.367
R1282 B.n244 B.n243 163.367
R1283 B.n244 B.n143 163.367
R1284 B.n248 B.n143 163.367
R1285 B.n249 B.n248 163.367
R1286 B.n250 B.n249 163.367
R1287 B.n250 B.n141 163.367
R1288 B.n254 B.n141 163.367
R1289 B.n255 B.n254 163.367
R1290 B.n256 B.n255 163.367
R1291 B.n256 B.n139 163.367
R1292 B.n260 B.n139 163.367
R1293 B.n261 B.n260 163.367
R1294 B.n262 B.n261 163.367
R1295 B.n262 B.n137 163.367
R1296 B.n266 B.n137 163.367
R1297 B.n267 B.n266 163.367
R1298 B.n268 B.n267 163.367
R1299 B.n268 B.n135 163.367
R1300 B.n272 B.n135 163.367
R1301 B.n273 B.n272 163.367
R1302 B.n274 B.n273 163.367
R1303 B.n274 B.n133 163.367
R1304 B.n278 B.n133 163.367
R1305 B.n279 B.n278 163.367
R1306 B.n279 B.n129 163.367
R1307 B.n283 B.n129 163.367
R1308 B.n284 B.n283 163.367
R1309 B.n285 B.n284 163.367
R1310 B.n285 B.n127 163.367
R1311 B.n289 B.n127 163.367
R1312 B.n290 B.n289 163.367
R1313 B.n291 B.n290 163.367
R1314 B.n291 B.n123 163.367
R1315 B.n296 B.n123 163.367
R1316 B.n297 B.n296 163.367
R1317 B.n298 B.n297 163.367
R1318 B.n298 B.n121 163.367
R1319 B.n302 B.n121 163.367
R1320 B.n303 B.n302 163.367
R1321 B.n304 B.n303 163.367
R1322 B.n304 B.n119 163.367
R1323 B.n308 B.n119 163.367
R1324 B.n309 B.n308 163.367
R1325 B.n310 B.n309 163.367
R1326 B.n310 B.n117 163.367
R1327 B.n314 B.n117 163.367
R1328 B.n315 B.n314 163.367
R1329 B.n316 B.n315 163.367
R1330 B.n316 B.n115 163.367
R1331 B.n320 B.n115 163.367
R1332 B.n321 B.n320 163.367
R1333 B.n322 B.n321 163.367
R1334 B.n322 B.n113 163.367
R1335 B.n326 B.n113 163.367
R1336 B.n327 B.n326 163.367
R1337 B.n328 B.n327 163.367
R1338 B.n328 B.n111 163.367
R1339 B.n332 B.n111 163.367
R1340 B.n333 B.n332 163.367
R1341 B.n334 B.n333 163.367
R1342 B.n334 B.n109 163.367
R1343 B.n338 B.n109 163.367
R1344 B.n339 B.n338 163.367
R1345 B.n340 B.n339 163.367
R1346 B.n340 B.n107 163.367
R1347 B.n344 B.n107 163.367
R1348 B.n345 B.n344 163.367
R1349 B.n346 B.n105 163.367
R1350 B.n350 B.n105 163.367
R1351 B.n351 B.n350 163.367
R1352 B.n352 B.n351 163.367
R1353 B.n352 B.n103 163.367
R1354 B.n356 B.n103 163.367
R1355 B.n357 B.n356 163.367
R1356 B.n358 B.n357 163.367
R1357 B.n358 B.n101 163.367
R1358 B.n362 B.n101 163.367
R1359 B.n363 B.n362 163.367
R1360 B.n364 B.n363 163.367
R1361 B.n364 B.n99 163.367
R1362 B.n368 B.n99 163.367
R1363 B.n369 B.n368 163.367
R1364 B.n370 B.n369 163.367
R1365 B.n370 B.n97 163.367
R1366 B.n374 B.n97 163.367
R1367 B.n375 B.n374 163.367
R1368 B.n376 B.n375 163.367
R1369 B.n376 B.n95 163.367
R1370 B.n380 B.n95 163.367
R1371 B.n381 B.n380 163.367
R1372 B.n382 B.n381 163.367
R1373 B.n382 B.n93 163.367
R1374 B.n386 B.n93 163.367
R1375 B.n387 B.n386 163.367
R1376 B.n388 B.n387 163.367
R1377 B.n388 B.n91 163.367
R1378 B.n392 B.n91 163.367
R1379 B.n393 B.n392 163.367
R1380 B.n394 B.n393 163.367
R1381 B.n394 B.n89 163.367
R1382 B.n398 B.n89 163.367
R1383 B.n399 B.n398 163.367
R1384 B.n400 B.n399 163.367
R1385 B.n400 B.n87 163.367
R1386 B.n404 B.n87 163.367
R1387 B.n405 B.n404 163.367
R1388 B.n406 B.n405 163.367
R1389 B.n406 B.n85 163.367
R1390 B.n410 B.n85 163.367
R1391 B.n411 B.n410 163.367
R1392 B.n412 B.n411 163.367
R1393 B.n412 B.n83 163.367
R1394 B.n416 B.n83 163.367
R1395 B.n417 B.n416 163.367
R1396 B.n418 B.n417 163.367
R1397 B.n418 B.n81 163.367
R1398 B.n422 B.n81 163.367
R1399 B.n423 B.n422 163.367
R1400 B.n424 B.n423 163.367
R1401 B.n424 B.n79 163.367
R1402 B.n428 B.n79 163.367
R1403 B.n429 B.n428 163.367
R1404 B.n430 B.n429 163.367
R1405 B.n430 B.n77 163.367
R1406 B.n434 B.n77 163.367
R1407 B.n435 B.n434 163.367
R1408 B.n436 B.n435 163.367
R1409 B.n436 B.n75 163.367
R1410 B.n440 B.n75 163.367
R1411 B.n441 B.n440 163.367
R1412 B.n442 B.n441 163.367
R1413 B.n442 B.n73 163.367
R1414 B.n446 B.n73 163.367
R1415 B.n447 B.n446 163.367
R1416 B.n448 B.n447 163.367
R1417 B.n448 B.n71 163.367
R1418 B.n452 B.n71 163.367
R1419 B.n453 B.n452 163.367
R1420 B.n454 B.n453 163.367
R1421 B.n454 B.n69 163.367
R1422 B.n458 B.n69 163.367
R1423 B.n459 B.n458 163.367
R1424 B.n460 B.n459 163.367
R1425 B.n460 B.n67 163.367
R1426 B.n464 B.n67 163.367
R1427 B.n465 B.n464 163.367
R1428 B.n466 B.n465 163.367
R1429 B.n585 B.n584 163.367
R1430 B.n584 B.n23 163.367
R1431 B.n580 B.n23 163.367
R1432 B.n580 B.n579 163.367
R1433 B.n579 B.n578 163.367
R1434 B.n578 B.n25 163.367
R1435 B.n574 B.n25 163.367
R1436 B.n574 B.n573 163.367
R1437 B.n573 B.n572 163.367
R1438 B.n572 B.n27 163.367
R1439 B.n568 B.n27 163.367
R1440 B.n568 B.n567 163.367
R1441 B.n567 B.n566 163.367
R1442 B.n566 B.n29 163.367
R1443 B.n562 B.n29 163.367
R1444 B.n562 B.n561 163.367
R1445 B.n561 B.n560 163.367
R1446 B.n560 B.n31 163.367
R1447 B.n556 B.n31 163.367
R1448 B.n556 B.n555 163.367
R1449 B.n555 B.n554 163.367
R1450 B.n554 B.n33 163.367
R1451 B.n550 B.n33 163.367
R1452 B.n550 B.n549 163.367
R1453 B.n549 B.n548 163.367
R1454 B.n548 B.n35 163.367
R1455 B.n544 B.n35 163.367
R1456 B.n544 B.n543 163.367
R1457 B.n543 B.n542 163.367
R1458 B.n542 B.n37 163.367
R1459 B.n538 B.n37 163.367
R1460 B.n538 B.n537 163.367
R1461 B.n537 B.n536 163.367
R1462 B.n536 B.n39 163.367
R1463 B.n531 B.n39 163.367
R1464 B.n531 B.n530 163.367
R1465 B.n530 B.n529 163.367
R1466 B.n529 B.n43 163.367
R1467 B.n525 B.n43 163.367
R1468 B.n525 B.n524 163.367
R1469 B.n524 B.n523 163.367
R1470 B.n523 B.n45 163.367
R1471 B.n519 B.n45 163.367
R1472 B.n519 B.n518 163.367
R1473 B.n518 B.n49 163.367
R1474 B.n514 B.n49 163.367
R1475 B.n514 B.n513 163.367
R1476 B.n513 B.n512 163.367
R1477 B.n512 B.n51 163.367
R1478 B.n508 B.n51 163.367
R1479 B.n508 B.n507 163.367
R1480 B.n507 B.n506 163.367
R1481 B.n506 B.n53 163.367
R1482 B.n502 B.n53 163.367
R1483 B.n502 B.n501 163.367
R1484 B.n501 B.n500 163.367
R1485 B.n500 B.n55 163.367
R1486 B.n496 B.n55 163.367
R1487 B.n496 B.n495 163.367
R1488 B.n495 B.n494 163.367
R1489 B.n494 B.n57 163.367
R1490 B.n490 B.n57 163.367
R1491 B.n490 B.n489 163.367
R1492 B.n489 B.n488 163.367
R1493 B.n488 B.n59 163.367
R1494 B.n484 B.n59 163.367
R1495 B.n484 B.n483 163.367
R1496 B.n483 B.n482 163.367
R1497 B.n482 B.n61 163.367
R1498 B.n478 B.n61 163.367
R1499 B.n478 B.n477 163.367
R1500 B.n477 B.n476 163.367
R1501 B.n476 B.n63 163.367
R1502 B.n472 B.n63 163.367
R1503 B.n472 B.n471 163.367
R1504 B.n471 B.n470 163.367
R1505 B.n470 B.n65 163.367
R1506 B.n294 B.n125 59.5399
R1507 B.n132 B.n131 59.5399
R1508 B.n534 B.n41 59.5399
R1509 B.n48 B.n47 59.5399
R1510 B.n125 B.n124 34.9096
R1511 B.n131 B.n130 34.9096
R1512 B.n41 B.n40 34.9096
R1513 B.n47 B.n46 34.9096
R1514 B.n587 B.n22 29.1907
R1515 B.n468 B.n467 29.1907
R1516 B.n347 B.n106 29.1907
R1517 B.n228 B.n227 29.1907
R1518 B B.n647 18.0485
R1519 B.n583 B.n22 10.6151
R1520 B.n583 B.n582 10.6151
R1521 B.n582 B.n581 10.6151
R1522 B.n581 B.n24 10.6151
R1523 B.n577 B.n24 10.6151
R1524 B.n577 B.n576 10.6151
R1525 B.n576 B.n575 10.6151
R1526 B.n575 B.n26 10.6151
R1527 B.n571 B.n26 10.6151
R1528 B.n571 B.n570 10.6151
R1529 B.n570 B.n569 10.6151
R1530 B.n569 B.n28 10.6151
R1531 B.n565 B.n28 10.6151
R1532 B.n565 B.n564 10.6151
R1533 B.n564 B.n563 10.6151
R1534 B.n563 B.n30 10.6151
R1535 B.n559 B.n30 10.6151
R1536 B.n559 B.n558 10.6151
R1537 B.n558 B.n557 10.6151
R1538 B.n557 B.n32 10.6151
R1539 B.n553 B.n32 10.6151
R1540 B.n553 B.n552 10.6151
R1541 B.n552 B.n551 10.6151
R1542 B.n551 B.n34 10.6151
R1543 B.n547 B.n34 10.6151
R1544 B.n547 B.n546 10.6151
R1545 B.n546 B.n545 10.6151
R1546 B.n545 B.n36 10.6151
R1547 B.n541 B.n36 10.6151
R1548 B.n541 B.n540 10.6151
R1549 B.n540 B.n539 10.6151
R1550 B.n539 B.n38 10.6151
R1551 B.n535 B.n38 10.6151
R1552 B.n533 B.n532 10.6151
R1553 B.n532 B.n42 10.6151
R1554 B.n528 B.n42 10.6151
R1555 B.n528 B.n527 10.6151
R1556 B.n527 B.n526 10.6151
R1557 B.n526 B.n44 10.6151
R1558 B.n522 B.n44 10.6151
R1559 B.n522 B.n521 10.6151
R1560 B.n521 B.n520 10.6151
R1561 B.n517 B.n516 10.6151
R1562 B.n516 B.n515 10.6151
R1563 B.n515 B.n50 10.6151
R1564 B.n511 B.n50 10.6151
R1565 B.n511 B.n510 10.6151
R1566 B.n510 B.n509 10.6151
R1567 B.n509 B.n52 10.6151
R1568 B.n505 B.n52 10.6151
R1569 B.n505 B.n504 10.6151
R1570 B.n504 B.n503 10.6151
R1571 B.n503 B.n54 10.6151
R1572 B.n499 B.n54 10.6151
R1573 B.n499 B.n498 10.6151
R1574 B.n498 B.n497 10.6151
R1575 B.n497 B.n56 10.6151
R1576 B.n493 B.n56 10.6151
R1577 B.n493 B.n492 10.6151
R1578 B.n492 B.n491 10.6151
R1579 B.n491 B.n58 10.6151
R1580 B.n487 B.n58 10.6151
R1581 B.n487 B.n486 10.6151
R1582 B.n486 B.n485 10.6151
R1583 B.n485 B.n60 10.6151
R1584 B.n481 B.n60 10.6151
R1585 B.n481 B.n480 10.6151
R1586 B.n480 B.n479 10.6151
R1587 B.n479 B.n62 10.6151
R1588 B.n475 B.n62 10.6151
R1589 B.n475 B.n474 10.6151
R1590 B.n474 B.n473 10.6151
R1591 B.n473 B.n64 10.6151
R1592 B.n469 B.n64 10.6151
R1593 B.n469 B.n468 10.6151
R1594 B.n348 B.n347 10.6151
R1595 B.n349 B.n348 10.6151
R1596 B.n349 B.n104 10.6151
R1597 B.n353 B.n104 10.6151
R1598 B.n354 B.n353 10.6151
R1599 B.n355 B.n354 10.6151
R1600 B.n355 B.n102 10.6151
R1601 B.n359 B.n102 10.6151
R1602 B.n360 B.n359 10.6151
R1603 B.n361 B.n360 10.6151
R1604 B.n361 B.n100 10.6151
R1605 B.n365 B.n100 10.6151
R1606 B.n366 B.n365 10.6151
R1607 B.n367 B.n366 10.6151
R1608 B.n367 B.n98 10.6151
R1609 B.n371 B.n98 10.6151
R1610 B.n372 B.n371 10.6151
R1611 B.n373 B.n372 10.6151
R1612 B.n373 B.n96 10.6151
R1613 B.n377 B.n96 10.6151
R1614 B.n378 B.n377 10.6151
R1615 B.n379 B.n378 10.6151
R1616 B.n379 B.n94 10.6151
R1617 B.n383 B.n94 10.6151
R1618 B.n384 B.n383 10.6151
R1619 B.n385 B.n384 10.6151
R1620 B.n385 B.n92 10.6151
R1621 B.n389 B.n92 10.6151
R1622 B.n390 B.n389 10.6151
R1623 B.n391 B.n390 10.6151
R1624 B.n391 B.n90 10.6151
R1625 B.n395 B.n90 10.6151
R1626 B.n396 B.n395 10.6151
R1627 B.n397 B.n396 10.6151
R1628 B.n397 B.n88 10.6151
R1629 B.n401 B.n88 10.6151
R1630 B.n402 B.n401 10.6151
R1631 B.n403 B.n402 10.6151
R1632 B.n403 B.n86 10.6151
R1633 B.n407 B.n86 10.6151
R1634 B.n408 B.n407 10.6151
R1635 B.n409 B.n408 10.6151
R1636 B.n409 B.n84 10.6151
R1637 B.n413 B.n84 10.6151
R1638 B.n414 B.n413 10.6151
R1639 B.n415 B.n414 10.6151
R1640 B.n415 B.n82 10.6151
R1641 B.n419 B.n82 10.6151
R1642 B.n420 B.n419 10.6151
R1643 B.n421 B.n420 10.6151
R1644 B.n421 B.n80 10.6151
R1645 B.n425 B.n80 10.6151
R1646 B.n426 B.n425 10.6151
R1647 B.n427 B.n426 10.6151
R1648 B.n427 B.n78 10.6151
R1649 B.n431 B.n78 10.6151
R1650 B.n432 B.n431 10.6151
R1651 B.n433 B.n432 10.6151
R1652 B.n433 B.n76 10.6151
R1653 B.n437 B.n76 10.6151
R1654 B.n438 B.n437 10.6151
R1655 B.n439 B.n438 10.6151
R1656 B.n439 B.n74 10.6151
R1657 B.n443 B.n74 10.6151
R1658 B.n444 B.n443 10.6151
R1659 B.n445 B.n444 10.6151
R1660 B.n445 B.n72 10.6151
R1661 B.n449 B.n72 10.6151
R1662 B.n450 B.n449 10.6151
R1663 B.n451 B.n450 10.6151
R1664 B.n451 B.n70 10.6151
R1665 B.n455 B.n70 10.6151
R1666 B.n456 B.n455 10.6151
R1667 B.n457 B.n456 10.6151
R1668 B.n457 B.n68 10.6151
R1669 B.n461 B.n68 10.6151
R1670 B.n462 B.n461 10.6151
R1671 B.n463 B.n462 10.6151
R1672 B.n463 B.n66 10.6151
R1673 B.n467 B.n66 10.6151
R1674 B.n229 B.n228 10.6151
R1675 B.n229 B.n148 10.6151
R1676 B.n233 B.n148 10.6151
R1677 B.n234 B.n233 10.6151
R1678 B.n235 B.n234 10.6151
R1679 B.n235 B.n146 10.6151
R1680 B.n239 B.n146 10.6151
R1681 B.n240 B.n239 10.6151
R1682 B.n241 B.n240 10.6151
R1683 B.n241 B.n144 10.6151
R1684 B.n245 B.n144 10.6151
R1685 B.n246 B.n245 10.6151
R1686 B.n247 B.n246 10.6151
R1687 B.n247 B.n142 10.6151
R1688 B.n251 B.n142 10.6151
R1689 B.n252 B.n251 10.6151
R1690 B.n253 B.n252 10.6151
R1691 B.n253 B.n140 10.6151
R1692 B.n257 B.n140 10.6151
R1693 B.n258 B.n257 10.6151
R1694 B.n259 B.n258 10.6151
R1695 B.n259 B.n138 10.6151
R1696 B.n263 B.n138 10.6151
R1697 B.n264 B.n263 10.6151
R1698 B.n265 B.n264 10.6151
R1699 B.n265 B.n136 10.6151
R1700 B.n269 B.n136 10.6151
R1701 B.n270 B.n269 10.6151
R1702 B.n271 B.n270 10.6151
R1703 B.n271 B.n134 10.6151
R1704 B.n275 B.n134 10.6151
R1705 B.n276 B.n275 10.6151
R1706 B.n277 B.n276 10.6151
R1707 B.n281 B.n280 10.6151
R1708 B.n282 B.n281 10.6151
R1709 B.n282 B.n128 10.6151
R1710 B.n286 B.n128 10.6151
R1711 B.n287 B.n286 10.6151
R1712 B.n288 B.n287 10.6151
R1713 B.n288 B.n126 10.6151
R1714 B.n292 B.n126 10.6151
R1715 B.n293 B.n292 10.6151
R1716 B.n295 B.n122 10.6151
R1717 B.n299 B.n122 10.6151
R1718 B.n300 B.n299 10.6151
R1719 B.n301 B.n300 10.6151
R1720 B.n301 B.n120 10.6151
R1721 B.n305 B.n120 10.6151
R1722 B.n306 B.n305 10.6151
R1723 B.n307 B.n306 10.6151
R1724 B.n307 B.n118 10.6151
R1725 B.n311 B.n118 10.6151
R1726 B.n312 B.n311 10.6151
R1727 B.n313 B.n312 10.6151
R1728 B.n313 B.n116 10.6151
R1729 B.n317 B.n116 10.6151
R1730 B.n318 B.n317 10.6151
R1731 B.n319 B.n318 10.6151
R1732 B.n319 B.n114 10.6151
R1733 B.n323 B.n114 10.6151
R1734 B.n324 B.n323 10.6151
R1735 B.n325 B.n324 10.6151
R1736 B.n325 B.n112 10.6151
R1737 B.n329 B.n112 10.6151
R1738 B.n330 B.n329 10.6151
R1739 B.n331 B.n330 10.6151
R1740 B.n331 B.n110 10.6151
R1741 B.n335 B.n110 10.6151
R1742 B.n336 B.n335 10.6151
R1743 B.n337 B.n336 10.6151
R1744 B.n337 B.n108 10.6151
R1745 B.n341 B.n108 10.6151
R1746 B.n342 B.n341 10.6151
R1747 B.n343 B.n342 10.6151
R1748 B.n343 B.n106 10.6151
R1749 B.n227 B.n150 10.6151
R1750 B.n223 B.n150 10.6151
R1751 B.n223 B.n222 10.6151
R1752 B.n222 B.n221 10.6151
R1753 B.n221 B.n152 10.6151
R1754 B.n217 B.n152 10.6151
R1755 B.n217 B.n216 10.6151
R1756 B.n216 B.n215 10.6151
R1757 B.n215 B.n154 10.6151
R1758 B.n211 B.n154 10.6151
R1759 B.n211 B.n210 10.6151
R1760 B.n210 B.n209 10.6151
R1761 B.n209 B.n156 10.6151
R1762 B.n205 B.n156 10.6151
R1763 B.n205 B.n204 10.6151
R1764 B.n204 B.n203 10.6151
R1765 B.n203 B.n158 10.6151
R1766 B.n199 B.n158 10.6151
R1767 B.n199 B.n198 10.6151
R1768 B.n198 B.n197 10.6151
R1769 B.n197 B.n160 10.6151
R1770 B.n193 B.n160 10.6151
R1771 B.n193 B.n192 10.6151
R1772 B.n192 B.n191 10.6151
R1773 B.n191 B.n162 10.6151
R1774 B.n187 B.n162 10.6151
R1775 B.n187 B.n186 10.6151
R1776 B.n186 B.n185 10.6151
R1777 B.n185 B.n164 10.6151
R1778 B.n181 B.n164 10.6151
R1779 B.n181 B.n180 10.6151
R1780 B.n180 B.n179 10.6151
R1781 B.n179 B.n166 10.6151
R1782 B.n175 B.n166 10.6151
R1783 B.n175 B.n174 10.6151
R1784 B.n174 B.n173 10.6151
R1785 B.n173 B.n168 10.6151
R1786 B.n169 B.n168 10.6151
R1787 B.n169 B.n0 10.6151
R1788 B.n643 B.n1 10.6151
R1789 B.n643 B.n642 10.6151
R1790 B.n642 B.n641 10.6151
R1791 B.n641 B.n4 10.6151
R1792 B.n637 B.n4 10.6151
R1793 B.n637 B.n636 10.6151
R1794 B.n636 B.n635 10.6151
R1795 B.n635 B.n6 10.6151
R1796 B.n631 B.n6 10.6151
R1797 B.n631 B.n630 10.6151
R1798 B.n630 B.n629 10.6151
R1799 B.n629 B.n8 10.6151
R1800 B.n625 B.n8 10.6151
R1801 B.n625 B.n624 10.6151
R1802 B.n624 B.n623 10.6151
R1803 B.n623 B.n10 10.6151
R1804 B.n619 B.n10 10.6151
R1805 B.n619 B.n618 10.6151
R1806 B.n618 B.n617 10.6151
R1807 B.n617 B.n12 10.6151
R1808 B.n613 B.n12 10.6151
R1809 B.n613 B.n612 10.6151
R1810 B.n612 B.n611 10.6151
R1811 B.n611 B.n14 10.6151
R1812 B.n607 B.n14 10.6151
R1813 B.n607 B.n606 10.6151
R1814 B.n606 B.n605 10.6151
R1815 B.n605 B.n16 10.6151
R1816 B.n601 B.n16 10.6151
R1817 B.n601 B.n600 10.6151
R1818 B.n600 B.n599 10.6151
R1819 B.n599 B.n18 10.6151
R1820 B.n595 B.n18 10.6151
R1821 B.n595 B.n594 10.6151
R1822 B.n594 B.n593 10.6151
R1823 B.n593 B.n20 10.6151
R1824 B.n589 B.n20 10.6151
R1825 B.n589 B.n588 10.6151
R1826 B.n588 B.n587 10.6151
R1827 B.n535 B.n534 9.36635
R1828 B.n517 B.n48 9.36635
R1829 B.n277 B.n132 9.36635
R1830 B.n295 B.n294 9.36635
R1831 B.n647 B.n0 2.81026
R1832 B.n647 B.n1 2.81026
R1833 B.n534 B.n533 1.24928
R1834 B.n520 B.n48 1.24928
R1835 B.n280 B.n132 1.24928
R1836 B.n294 B.n293 1.24928
C0 VN VDD2 7.31922f
C1 VP VDD1 7.604259f
C2 VN VDD1 0.151126f
C3 VP B 1.64147f
C4 VN B 0.968314f
C5 w_n3130_n2852# VDD2 2.25751f
C6 VTAIL VDD2 9.399099f
C7 VDD1 w_n3130_n2852# 2.17267f
C8 VTAIL VDD1 9.35652f
C9 VP VN 6.25356f
C10 w_n3130_n2852# B 7.92289f
C11 VTAIL B 2.67812f
C12 VDD1 VDD2 1.43942f
C13 VP w_n3130_n2852# 6.70627f
C14 VP VTAIL 7.60886f
C15 VDD2 B 1.90637f
C16 VN w_n3130_n2852# 6.30225f
C17 VN VTAIL 7.5945f
C18 VDD1 B 1.83246f
C19 VP VDD2 0.439602f
C20 VTAIL w_n3130_n2852# 2.69765f
C21 VDD2 VSUBS 1.569504f
C22 VDD1 VSUBS 1.407709f
C23 VTAIL VSUBS 0.934235f
C24 VN VSUBS 5.7736f
C25 VP VSUBS 2.68907f
C26 B VSUBS 3.74483f
C27 w_n3130_n2852# VSUBS 0.110389p
C28 B.n0 VSUBS 0.004516f
C29 B.n1 VSUBS 0.004516f
C30 B.n2 VSUBS 0.007142f
C31 B.n3 VSUBS 0.007142f
C32 B.n4 VSUBS 0.007142f
C33 B.n5 VSUBS 0.007142f
C34 B.n6 VSUBS 0.007142f
C35 B.n7 VSUBS 0.007142f
C36 B.n8 VSUBS 0.007142f
C37 B.n9 VSUBS 0.007142f
C38 B.n10 VSUBS 0.007142f
C39 B.n11 VSUBS 0.007142f
C40 B.n12 VSUBS 0.007142f
C41 B.n13 VSUBS 0.007142f
C42 B.n14 VSUBS 0.007142f
C43 B.n15 VSUBS 0.007142f
C44 B.n16 VSUBS 0.007142f
C45 B.n17 VSUBS 0.007142f
C46 B.n18 VSUBS 0.007142f
C47 B.n19 VSUBS 0.007142f
C48 B.n20 VSUBS 0.007142f
C49 B.n21 VSUBS 0.007142f
C50 B.n22 VSUBS 0.016039f
C51 B.n23 VSUBS 0.007142f
C52 B.n24 VSUBS 0.007142f
C53 B.n25 VSUBS 0.007142f
C54 B.n26 VSUBS 0.007142f
C55 B.n27 VSUBS 0.007142f
C56 B.n28 VSUBS 0.007142f
C57 B.n29 VSUBS 0.007142f
C58 B.n30 VSUBS 0.007142f
C59 B.n31 VSUBS 0.007142f
C60 B.n32 VSUBS 0.007142f
C61 B.n33 VSUBS 0.007142f
C62 B.n34 VSUBS 0.007142f
C63 B.n35 VSUBS 0.007142f
C64 B.n36 VSUBS 0.007142f
C65 B.n37 VSUBS 0.007142f
C66 B.n38 VSUBS 0.007142f
C67 B.n39 VSUBS 0.007142f
C68 B.t11 VSUBS 0.158641f
C69 B.t10 VSUBS 0.178144f
C70 B.t9 VSUBS 0.627417f
C71 B.n40 VSUBS 0.28679f
C72 B.n41 VSUBS 0.213655f
C73 B.n42 VSUBS 0.007142f
C74 B.n43 VSUBS 0.007142f
C75 B.n44 VSUBS 0.007142f
C76 B.n45 VSUBS 0.007142f
C77 B.t2 VSUBS 0.158644f
C78 B.t1 VSUBS 0.178147f
C79 B.t0 VSUBS 0.627417f
C80 B.n46 VSUBS 0.286788f
C81 B.n47 VSUBS 0.213652f
C82 B.n48 VSUBS 0.016547f
C83 B.n49 VSUBS 0.007142f
C84 B.n50 VSUBS 0.007142f
C85 B.n51 VSUBS 0.007142f
C86 B.n52 VSUBS 0.007142f
C87 B.n53 VSUBS 0.007142f
C88 B.n54 VSUBS 0.007142f
C89 B.n55 VSUBS 0.007142f
C90 B.n56 VSUBS 0.007142f
C91 B.n57 VSUBS 0.007142f
C92 B.n58 VSUBS 0.007142f
C93 B.n59 VSUBS 0.007142f
C94 B.n60 VSUBS 0.007142f
C95 B.n61 VSUBS 0.007142f
C96 B.n62 VSUBS 0.007142f
C97 B.n63 VSUBS 0.007142f
C98 B.n64 VSUBS 0.007142f
C99 B.n65 VSUBS 0.016039f
C100 B.n66 VSUBS 0.007142f
C101 B.n67 VSUBS 0.007142f
C102 B.n68 VSUBS 0.007142f
C103 B.n69 VSUBS 0.007142f
C104 B.n70 VSUBS 0.007142f
C105 B.n71 VSUBS 0.007142f
C106 B.n72 VSUBS 0.007142f
C107 B.n73 VSUBS 0.007142f
C108 B.n74 VSUBS 0.007142f
C109 B.n75 VSUBS 0.007142f
C110 B.n76 VSUBS 0.007142f
C111 B.n77 VSUBS 0.007142f
C112 B.n78 VSUBS 0.007142f
C113 B.n79 VSUBS 0.007142f
C114 B.n80 VSUBS 0.007142f
C115 B.n81 VSUBS 0.007142f
C116 B.n82 VSUBS 0.007142f
C117 B.n83 VSUBS 0.007142f
C118 B.n84 VSUBS 0.007142f
C119 B.n85 VSUBS 0.007142f
C120 B.n86 VSUBS 0.007142f
C121 B.n87 VSUBS 0.007142f
C122 B.n88 VSUBS 0.007142f
C123 B.n89 VSUBS 0.007142f
C124 B.n90 VSUBS 0.007142f
C125 B.n91 VSUBS 0.007142f
C126 B.n92 VSUBS 0.007142f
C127 B.n93 VSUBS 0.007142f
C128 B.n94 VSUBS 0.007142f
C129 B.n95 VSUBS 0.007142f
C130 B.n96 VSUBS 0.007142f
C131 B.n97 VSUBS 0.007142f
C132 B.n98 VSUBS 0.007142f
C133 B.n99 VSUBS 0.007142f
C134 B.n100 VSUBS 0.007142f
C135 B.n101 VSUBS 0.007142f
C136 B.n102 VSUBS 0.007142f
C137 B.n103 VSUBS 0.007142f
C138 B.n104 VSUBS 0.007142f
C139 B.n105 VSUBS 0.007142f
C140 B.n106 VSUBS 0.016039f
C141 B.n107 VSUBS 0.007142f
C142 B.n108 VSUBS 0.007142f
C143 B.n109 VSUBS 0.007142f
C144 B.n110 VSUBS 0.007142f
C145 B.n111 VSUBS 0.007142f
C146 B.n112 VSUBS 0.007142f
C147 B.n113 VSUBS 0.007142f
C148 B.n114 VSUBS 0.007142f
C149 B.n115 VSUBS 0.007142f
C150 B.n116 VSUBS 0.007142f
C151 B.n117 VSUBS 0.007142f
C152 B.n118 VSUBS 0.007142f
C153 B.n119 VSUBS 0.007142f
C154 B.n120 VSUBS 0.007142f
C155 B.n121 VSUBS 0.007142f
C156 B.n122 VSUBS 0.007142f
C157 B.n123 VSUBS 0.007142f
C158 B.t4 VSUBS 0.158644f
C159 B.t5 VSUBS 0.178147f
C160 B.t3 VSUBS 0.627417f
C161 B.n124 VSUBS 0.286788f
C162 B.n125 VSUBS 0.213652f
C163 B.n126 VSUBS 0.007142f
C164 B.n127 VSUBS 0.007142f
C165 B.n128 VSUBS 0.007142f
C166 B.n129 VSUBS 0.007142f
C167 B.t7 VSUBS 0.158641f
C168 B.t8 VSUBS 0.178144f
C169 B.t6 VSUBS 0.627417f
C170 B.n130 VSUBS 0.28679f
C171 B.n131 VSUBS 0.213655f
C172 B.n132 VSUBS 0.016547f
C173 B.n133 VSUBS 0.007142f
C174 B.n134 VSUBS 0.007142f
C175 B.n135 VSUBS 0.007142f
C176 B.n136 VSUBS 0.007142f
C177 B.n137 VSUBS 0.007142f
C178 B.n138 VSUBS 0.007142f
C179 B.n139 VSUBS 0.007142f
C180 B.n140 VSUBS 0.007142f
C181 B.n141 VSUBS 0.007142f
C182 B.n142 VSUBS 0.007142f
C183 B.n143 VSUBS 0.007142f
C184 B.n144 VSUBS 0.007142f
C185 B.n145 VSUBS 0.007142f
C186 B.n146 VSUBS 0.007142f
C187 B.n147 VSUBS 0.007142f
C188 B.n148 VSUBS 0.007142f
C189 B.n149 VSUBS 0.016039f
C190 B.n150 VSUBS 0.007142f
C191 B.n151 VSUBS 0.007142f
C192 B.n152 VSUBS 0.007142f
C193 B.n153 VSUBS 0.007142f
C194 B.n154 VSUBS 0.007142f
C195 B.n155 VSUBS 0.007142f
C196 B.n156 VSUBS 0.007142f
C197 B.n157 VSUBS 0.007142f
C198 B.n158 VSUBS 0.007142f
C199 B.n159 VSUBS 0.007142f
C200 B.n160 VSUBS 0.007142f
C201 B.n161 VSUBS 0.007142f
C202 B.n162 VSUBS 0.007142f
C203 B.n163 VSUBS 0.007142f
C204 B.n164 VSUBS 0.007142f
C205 B.n165 VSUBS 0.007142f
C206 B.n166 VSUBS 0.007142f
C207 B.n167 VSUBS 0.007142f
C208 B.n168 VSUBS 0.007142f
C209 B.n169 VSUBS 0.007142f
C210 B.n170 VSUBS 0.007142f
C211 B.n171 VSUBS 0.007142f
C212 B.n172 VSUBS 0.007142f
C213 B.n173 VSUBS 0.007142f
C214 B.n174 VSUBS 0.007142f
C215 B.n175 VSUBS 0.007142f
C216 B.n176 VSUBS 0.007142f
C217 B.n177 VSUBS 0.007142f
C218 B.n178 VSUBS 0.007142f
C219 B.n179 VSUBS 0.007142f
C220 B.n180 VSUBS 0.007142f
C221 B.n181 VSUBS 0.007142f
C222 B.n182 VSUBS 0.007142f
C223 B.n183 VSUBS 0.007142f
C224 B.n184 VSUBS 0.007142f
C225 B.n185 VSUBS 0.007142f
C226 B.n186 VSUBS 0.007142f
C227 B.n187 VSUBS 0.007142f
C228 B.n188 VSUBS 0.007142f
C229 B.n189 VSUBS 0.007142f
C230 B.n190 VSUBS 0.007142f
C231 B.n191 VSUBS 0.007142f
C232 B.n192 VSUBS 0.007142f
C233 B.n193 VSUBS 0.007142f
C234 B.n194 VSUBS 0.007142f
C235 B.n195 VSUBS 0.007142f
C236 B.n196 VSUBS 0.007142f
C237 B.n197 VSUBS 0.007142f
C238 B.n198 VSUBS 0.007142f
C239 B.n199 VSUBS 0.007142f
C240 B.n200 VSUBS 0.007142f
C241 B.n201 VSUBS 0.007142f
C242 B.n202 VSUBS 0.007142f
C243 B.n203 VSUBS 0.007142f
C244 B.n204 VSUBS 0.007142f
C245 B.n205 VSUBS 0.007142f
C246 B.n206 VSUBS 0.007142f
C247 B.n207 VSUBS 0.007142f
C248 B.n208 VSUBS 0.007142f
C249 B.n209 VSUBS 0.007142f
C250 B.n210 VSUBS 0.007142f
C251 B.n211 VSUBS 0.007142f
C252 B.n212 VSUBS 0.007142f
C253 B.n213 VSUBS 0.007142f
C254 B.n214 VSUBS 0.007142f
C255 B.n215 VSUBS 0.007142f
C256 B.n216 VSUBS 0.007142f
C257 B.n217 VSUBS 0.007142f
C258 B.n218 VSUBS 0.007142f
C259 B.n219 VSUBS 0.007142f
C260 B.n220 VSUBS 0.007142f
C261 B.n221 VSUBS 0.007142f
C262 B.n222 VSUBS 0.007142f
C263 B.n223 VSUBS 0.007142f
C264 B.n224 VSUBS 0.007142f
C265 B.n225 VSUBS 0.007142f
C266 B.n226 VSUBS 0.015049f
C267 B.n227 VSUBS 0.015049f
C268 B.n228 VSUBS 0.016039f
C269 B.n229 VSUBS 0.007142f
C270 B.n230 VSUBS 0.007142f
C271 B.n231 VSUBS 0.007142f
C272 B.n232 VSUBS 0.007142f
C273 B.n233 VSUBS 0.007142f
C274 B.n234 VSUBS 0.007142f
C275 B.n235 VSUBS 0.007142f
C276 B.n236 VSUBS 0.007142f
C277 B.n237 VSUBS 0.007142f
C278 B.n238 VSUBS 0.007142f
C279 B.n239 VSUBS 0.007142f
C280 B.n240 VSUBS 0.007142f
C281 B.n241 VSUBS 0.007142f
C282 B.n242 VSUBS 0.007142f
C283 B.n243 VSUBS 0.007142f
C284 B.n244 VSUBS 0.007142f
C285 B.n245 VSUBS 0.007142f
C286 B.n246 VSUBS 0.007142f
C287 B.n247 VSUBS 0.007142f
C288 B.n248 VSUBS 0.007142f
C289 B.n249 VSUBS 0.007142f
C290 B.n250 VSUBS 0.007142f
C291 B.n251 VSUBS 0.007142f
C292 B.n252 VSUBS 0.007142f
C293 B.n253 VSUBS 0.007142f
C294 B.n254 VSUBS 0.007142f
C295 B.n255 VSUBS 0.007142f
C296 B.n256 VSUBS 0.007142f
C297 B.n257 VSUBS 0.007142f
C298 B.n258 VSUBS 0.007142f
C299 B.n259 VSUBS 0.007142f
C300 B.n260 VSUBS 0.007142f
C301 B.n261 VSUBS 0.007142f
C302 B.n262 VSUBS 0.007142f
C303 B.n263 VSUBS 0.007142f
C304 B.n264 VSUBS 0.007142f
C305 B.n265 VSUBS 0.007142f
C306 B.n266 VSUBS 0.007142f
C307 B.n267 VSUBS 0.007142f
C308 B.n268 VSUBS 0.007142f
C309 B.n269 VSUBS 0.007142f
C310 B.n270 VSUBS 0.007142f
C311 B.n271 VSUBS 0.007142f
C312 B.n272 VSUBS 0.007142f
C313 B.n273 VSUBS 0.007142f
C314 B.n274 VSUBS 0.007142f
C315 B.n275 VSUBS 0.007142f
C316 B.n276 VSUBS 0.007142f
C317 B.n277 VSUBS 0.006722f
C318 B.n278 VSUBS 0.007142f
C319 B.n279 VSUBS 0.007142f
C320 B.n280 VSUBS 0.003991f
C321 B.n281 VSUBS 0.007142f
C322 B.n282 VSUBS 0.007142f
C323 B.n283 VSUBS 0.007142f
C324 B.n284 VSUBS 0.007142f
C325 B.n285 VSUBS 0.007142f
C326 B.n286 VSUBS 0.007142f
C327 B.n287 VSUBS 0.007142f
C328 B.n288 VSUBS 0.007142f
C329 B.n289 VSUBS 0.007142f
C330 B.n290 VSUBS 0.007142f
C331 B.n291 VSUBS 0.007142f
C332 B.n292 VSUBS 0.007142f
C333 B.n293 VSUBS 0.003991f
C334 B.n294 VSUBS 0.016547f
C335 B.n295 VSUBS 0.006722f
C336 B.n296 VSUBS 0.007142f
C337 B.n297 VSUBS 0.007142f
C338 B.n298 VSUBS 0.007142f
C339 B.n299 VSUBS 0.007142f
C340 B.n300 VSUBS 0.007142f
C341 B.n301 VSUBS 0.007142f
C342 B.n302 VSUBS 0.007142f
C343 B.n303 VSUBS 0.007142f
C344 B.n304 VSUBS 0.007142f
C345 B.n305 VSUBS 0.007142f
C346 B.n306 VSUBS 0.007142f
C347 B.n307 VSUBS 0.007142f
C348 B.n308 VSUBS 0.007142f
C349 B.n309 VSUBS 0.007142f
C350 B.n310 VSUBS 0.007142f
C351 B.n311 VSUBS 0.007142f
C352 B.n312 VSUBS 0.007142f
C353 B.n313 VSUBS 0.007142f
C354 B.n314 VSUBS 0.007142f
C355 B.n315 VSUBS 0.007142f
C356 B.n316 VSUBS 0.007142f
C357 B.n317 VSUBS 0.007142f
C358 B.n318 VSUBS 0.007142f
C359 B.n319 VSUBS 0.007142f
C360 B.n320 VSUBS 0.007142f
C361 B.n321 VSUBS 0.007142f
C362 B.n322 VSUBS 0.007142f
C363 B.n323 VSUBS 0.007142f
C364 B.n324 VSUBS 0.007142f
C365 B.n325 VSUBS 0.007142f
C366 B.n326 VSUBS 0.007142f
C367 B.n327 VSUBS 0.007142f
C368 B.n328 VSUBS 0.007142f
C369 B.n329 VSUBS 0.007142f
C370 B.n330 VSUBS 0.007142f
C371 B.n331 VSUBS 0.007142f
C372 B.n332 VSUBS 0.007142f
C373 B.n333 VSUBS 0.007142f
C374 B.n334 VSUBS 0.007142f
C375 B.n335 VSUBS 0.007142f
C376 B.n336 VSUBS 0.007142f
C377 B.n337 VSUBS 0.007142f
C378 B.n338 VSUBS 0.007142f
C379 B.n339 VSUBS 0.007142f
C380 B.n340 VSUBS 0.007142f
C381 B.n341 VSUBS 0.007142f
C382 B.n342 VSUBS 0.007142f
C383 B.n343 VSUBS 0.007142f
C384 B.n344 VSUBS 0.007142f
C385 B.n345 VSUBS 0.016039f
C386 B.n346 VSUBS 0.015049f
C387 B.n347 VSUBS 0.015049f
C388 B.n348 VSUBS 0.007142f
C389 B.n349 VSUBS 0.007142f
C390 B.n350 VSUBS 0.007142f
C391 B.n351 VSUBS 0.007142f
C392 B.n352 VSUBS 0.007142f
C393 B.n353 VSUBS 0.007142f
C394 B.n354 VSUBS 0.007142f
C395 B.n355 VSUBS 0.007142f
C396 B.n356 VSUBS 0.007142f
C397 B.n357 VSUBS 0.007142f
C398 B.n358 VSUBS 0.007142f
C399 B.n359 VSUBS 0.007142f
C400 B.n360 VSUBS 0.007142f
C401 B.n361 VSUBS 0.007142f
C402 B.n362 VSUBS 0.007142f
C403 B.n363 VSUBS 0.007142f
C404 B.n364 VSUBS 0.007142f
C405 B.n365 VSUBS 0.007142f
C406 B.n366 VSUBS 0.007142f
C407 B.n367 VSUBS 0.007142f
C408 B.n368 VSUBS 0.007142f
C409 B.n369 VSUBS 0.007142f
C410 B.n370 VSUBS 0.007142f
C411 B.n371 VSUBS 0.007142f
C412 B.n372 VSUBS 0.007142f
C413 B.n373 VSUBS 0.007142f
C414 B.n374 VSUBS 0.007142f
C415 B.n375 VSUBS 0.007142f
C416 B.n376 VSUBS 0.007142f
C417 B.n377 VSUBS 0.007142f
C418 B.n378 VSUBS 0.007142f
C419 B.n379 VSUBS 0.007142f
C420 B.n380 VSUBS 0.007142f
C421 B.n381 VSUBS 0.007142f
C422 B.n382 VSUBS 0.007142f
C423 B.n383 VSUBS 0.007142f
C424 B.n384 VSUBS 0.007142f
C425 B.n385 VSUBS 0.007142f
C426 B.n386 VSUBS 0.007142f
C427 B.n387 VSUBS 0.007142f
C428 B.n388 VSUBS 0.007142f
C429 B.n389 VSUBS 0.007142f
C430 B.n390 VSUBS 0.007142f
C431 B.n391 VSUBS 0.007142f
C432 B.n392 VSUBS 0.007142f
C433 B.n393 VSUBS 0.007142f
C434 B.n394 VSUBS 0.007142f
C435 B.n395 VSUBS 0.007142f
C436 B.n396 VSUBS 0.007142f
C437 B.n397 VSUBS 0.007142f
C438 B.n398 VSUBS 0.007142f
C439 B.n399 VSUBS 0.007142f
C440 B.n400 VSUBS 0.007142f
C441 B.n401 VSUBS 0.007142f
C442 B.n402 VSUBS 0.007142f
C443 B.n403 VSUBS 0.007142f
C444 B.n404 VSUBS 0.007142f
C445 B.n405 VSUBS 0.007142f
C446 B.n406 VSUBS 0.007142f
C447 B.n407 VSUBS 0.007142f
C448 B.n408 VSUBS 0.007142f
C449 B.n409 VSUBS 0.007142f
C450 B.n410 VSUBS 0.007142f
C451 B.n411 VSUBS 0.007142f
C452 B.n412 VSUBS 0.007142f
C453 B.n413 VSUBS 0.007142f
C454 B.n414 VSUBS 0.007142f
C455 B.n415 VSUBS 0.007142f
C456 B.n416 VSUBS 0.007142f
C457 B.n417 VSUBS 0.007142f
C458 B.n418 VSUBS 0.007142f
C459 B.n419 VSUBS 0.007142f
C460 B.n420 VSUBS 0.007142f
C461 B.n421 VSUBS 0.007142f
C462 B.n422 VSUBS 0.007142f
C463 B.n423 VSUBS 0.007142f
C464 B.n424 VSUBS 0.007142f
C465 B.n425 VSUBS 0.007142f
C466 B.n426 VSUBS 0.007142f
C467 B.n427 VSUBS 0.007142f
C468 B.n428 VSUBS 0.007142f
C469 B.n429 VSUBS 0.007142f
C470 B.n430 VSUBS 0.007142f
C471 B.n431 VSUBS 0.007142f
C472 B.n432 VSUBS 0.007142f
C473 B.n433 VSUBS 0.007142f
C474 B.n434 VSUBS 0.007142f
C475 B.n435 VSUBS 0.007142f
C476 B.n436 VSUBS 0.007142f
C477 B.n437 VSUBS 0.007142f
C478 B.n438 VSUBS 0.007142f
C479 B.n439 VSUBS 0.007142f
C480 B.n440 VSUBS 0.007142f
C481 B.n441 VSUBS 0.007142f
C482 B.n442 VSUBS 0.007142f
C483 B.n443 VSUBS 0.007142f
C484 B.n444 VSUBS 0.007142f
C485 B.n445 VSUBS 0.007142f
C486 B.n446 VSUBS 0.007142f
C487 B.n447 VSUBS 0.007142f
C488 B.n448 VSUBS 0.007142f
C489 B.n449 VSUBS 0.007142f
C490 B.n450 VSUBS 0.007142f
C491 B.n451 VSUBS 0.007142f
C492 B.n452 VSUBS 0.007142f
C493 B.n453 VSUBS 0.007142f
C494 B.n454 VSUBS 0.007142f
C495 B.n455 VSUBS 0.007142f
C496 B.n456 VSUBS 0.007142f
C497 B.n457 VSUBS 0.007142f
C498 B.n458 VSUBS 0.007142f
C499 B.n459 VSUBS 0.007142f
C500 B.n460 VSUBS 0.007142f
C501 B.n461 VSUBS 0.007142f
C502 B.n462 VSUBS 0.007142f
C503 B.n463 VSUBS 0.007142f
C504 B.n464 VSUBS 0.007142f
C505 B.n465 VSUBS 0.007142f
C506 B.n466 VSUBS 0.015049f
C507 B.n467 VSUBS 0.015993f
C508 B.n468 VSUBS 0.015095f
C509 B.n469 VSUBS 0.007142f
C510 B.n470 VSUBS 0.007142f
C511 B.n471 VSUBS 0.007142f
C512 B.n472 VSUBS 0.007142f
C513 B.n473 VSUBS 0.007142f
C514 B.n474 VSUBS 0.007142f
C515 B.n475 VSUBS 0.007142f
C516 B.n476 VSUBS 0.007142f
C517 B.n477 VSUBS 0.007142f
C518 B.n478 VSUBS 0.007142f
C519 B.n479 VSUBS 0.007142f
C520 B.n480 VSUBS 0.007142f
C521 B.n481 VSUBS 0.007142f
C522 B.n482 VSUBS 0.007142f
C523 B.n483 VSUBS 0.007142f
C524 B.n484 VSUBS 0.007142f
C525 B.n485 VSUBS 0.007142f
C526 B.n486 VSUBS 0.007142f
C527 B.n487 VSUBS 0.007142f
C528 B.n488 VSUBS 0.007142f
C529 B.n489 VSUBS 0.007142f
C530 B.n490 VSUBS 0.007142f
C531 B.n491 VSUBS 0.007142f
C532 B.n492 VSUBS 0.007142f
C533 B.n493 VSUBS 0.007142f
C534 B.n494 VSUBS 0.007142f
C535 B.n495 VSUBS 0.007142f
C536 B.n496 VSUBS 0.007142f
C537 B.n497 VSUBS 0.007142f
C538 B.n498 VSUBS 0.007142f
C539 B.n499 VSUBS 0.007142f
C540 B.n500 VSUBS 0.007142f
C541 B.n501 VSUBS 0.007142f
C542 B.n502 VSUBS 0.007142f
C543 B.n503 VSUBS 0.007142f
C544 B.n504 VSUBS 0.007142f
C545 B.n505 VSUBS 0.007142f
C546 B.n506 VSUBS 0.007142f
C547 B.n507 VSUBS 0.007142f
C548 B.n508 VSUBS 0.007142f
C549 B.n509 VSUBS 0.007142f
C550 B.n510 VSUBS 0.007142f
C551 B.n511 VSUBS 0.007142f
C552 B.n512 VSUBS 0.007142f
C553 B.n513 VSUBS 0.007142f
C554 B.n514 VSUBS 0.007142f
C555 B.n515 VSUBS 0.007142f
C556 B.n516 VSUBS 0.007142f
C557 B.n517 VSUBS 0.006722f
C558 B.n518 VSUBS 0.007142f
C559 B.n519 VSUBS 0.007142f
C560 B.n520 VSUBS 0.003991f
C561 B.n521 VSUBS 0.007142f
C562 B.n522 VSUBS 0.007142f
C563 B.n523 VSUBS 0.007142f
C564 B.n524 VSUBS 0.007142f
C565 B.n525 VSUBS 0.007142f
C566 B.n526 VSUBS 0.007142f
C567 B.n527 VSUBS 0.007142f
C568 B.n528 VSUBS 0.007142f
C569 B.n529 VSUBS 0.007142f
C570 B.n530 VSUBS 0.007142f
C571 B.n531 VSUBS 0.007142f
C572 B.n532 VSUBS 0.007142f
C573 B.n533 VSUBS 0.003991f
C574 B.n534 VSUBS 0.016547f
C575 B.n535 VSUBS 0.006722f
C576 B.n536 VSUBS 0.007142f
C577 B.n537 VSUBS 0.007142f
C578 B.n538 VSUBS 0.007142f
C579 B.n539 VSUBS 0.007142f
C580 B.n540 VSUBS 0.007142f
C581 B.n541 VSUBS 0.007142f
C582 B.n542 VSUBS 0.007142f
C583 B.n543 VSUBS 0.007142f
C584 B.n544 VSUBS 0.007142f
C585 B.n545 VSUBS 0.007142f
C586 B.n546 VSUBS 0.007142f
C587 B.n547 VSUBS 0.007142f
C588 B.n548 VSUBS 0.007142f
C589 B.n549 VSUBS 0.007142f
C590 B.n550 VSUBS 0.007142f
C591 B.n551 VSUBS 0.007142f
C592 B.n552 VSUBS 0.007142f
C593 B.n553 VSUBS 0.007142f
C594 B.n554 VSUBS 0.007142f
C595 B.n555 VSUBS 0.007142f
C596 B.n556 VSUBS 0.007142f
C597 B.n557 VSUBS 0.007142f
C598 B.n558 VSUBS 0.007142f
C599 B.n559 VSUBS 0.007142f
C600 B.n560 VSUBS 0.007142f
C601 B.n561 VSUBS 0.007142f
C602 B.n562 VSUBS 0.007142f
C603 B.n563 VSUBS 0.007142f
C604 B.n564 VSUBS 0.007142f
C605 B.n565 VSUBS 0.007142f
C606 B.n566 VSUBS 0.007142f
C607 B.n567 VSUBS 0.007142f
C608 B.n568 VSUBS 0.007142f
C609 B.n569 VSUBS 0.007142f
C610 B.n570 VSUBS 0.007142f
C611 B.n571 VSUBS 0.007142f
C612 B.n572 VSUBS 0.007142f
C613 B.n573 VSUBS 0.007142f
C614 B.n574 VSUBS 0.007142f
C615 B.n575 VSUBS 0.007142f
C616 B.n576 VSUBS 0.007142f
C617 B.n577 VSUBS 0.007142f
C618 B.n578 VSUBS 0.007142f
C619 B.n579 VSUBS 0.007142f
C620 B.n580 VSUBS 0.007142f
C621 B.n581 VSUBS 0.007142f
C622 B.n582 VSUBS 0.007142f
C623 B.n583 VSUBS 0.007142f
C624 B.n584 VSUBS 0.007142f
C625 B.n585 VSUBS 0.016039f
C626 B.n586 VSUBS 0.015049f
C627 B.n587 VSUBS 0.015049f
C628 B.n588 VSUBS 0.007142f
C629 B.n589 VSUBS 0.007142f
C630 B.n590 VSUBS 0.007142f
C631 B.n591 VSUBS 0.007142f
C632 B.n592 VSUBS 0.007142f
C633 B.n593 VSUBS 0.007142f
C634 B.n594 VSUBS 0.007142f
C635 B.n595 VSUBS 0.007142f
C636 B.n596 VSUBS 0.007142f
C637 B.n597 VSUBS 0.007142f
C638 B.n598 VSUBS 0.007142f
C639 B.n599 VSUBS 0.007142f
C640 B.n600 VSUBS 0.007142f
C641 B.n601 VSUBS 0.007142f
C642 B.n602 VSUBS 0.007142f
C643 B.n603 VSUBS 0.007142f
C644 B.n604 VSUBS 0.007142f
C645 B.n605 VSUBS 0.007142f
C646 B.n606 VSUBS 0.007142f
C647 B.n607 VSUBS 0.007142f
C648 B.n608 VSUBS 0.007142f
C649 B.n609 VSUBS 0.007142f
C650 B.n610 VSUBS 0.007142f
C651 B.n611 VSUBS 0.007142f
C652 B.n612 VSUBS 0.007142f
C653 B.n613 VSUBS 0.007142f
C654 B.n614 VSUBS 0.007142f
C655 B.n615 VSUBS 0.007142f
C656 B.n616 VSUBS 0.007142f
C657 B.n617 VSUBS 0.007142f
C658 B.n618 VSUBS 0.007142f
C659 B.n619 VSUBS 0.007142f
C660 B.n620 VSUBS 0.007142f
C661 B.n621 VSUBS 0.007142f
C662 B.n622 VSUBS 0.007142f
C663 B.n623 VSUBS 0.007142f
C664 B.n624 VSUBS 0.007142f
C665 B.n625 VSUBS 0.007142f
C666 B.n626 VSUBS 0.007142f
C667 B.n627 VSUBS 0.007142f
C668 B.n628 VSUBS 0.007142f
C669 B.n629 VSUBS 0.007142f
C670 B.n630 VSUBS 0.007142f
C671 B.n631 VSUBS 0.007142f
C672 B.n632 VSUBS 0.007142f
C673 B.n633 VSUBS 0.007142f
C674 B.n634 VSUBS 0.007142f
C675 B.n635 VSUBS 0.007142f
C676 B.n636 VSUBS 0.007142f
C677 B.n637 VSUBS 0.007142f
C678 B.n638 VSUBS 0.007142f
C679 B.n639 VSUBS 0.007142f
C680 B.n640 VSUBS 0.007142f
C681 B.n641 VSUBS 0.007142f
C682 B.n642 VSUBS 0.007142f
C683 B.n643 VSUBS 0.007142f
C684 B.n644 VSUBS 0.007142f
C685 B.n645 VSUBS 0.007142f
C686 B.n646 VSUBS 0.007142f
C687 B.n647 VSUBS 0.016172f
C688 VDD1.n0 VSUBS 0.028512f
C689 VDD1.n1 VSUBS 0.025848f
C690 VDD1.n2 VSUBS 0.013889f
C691 VDD1.n3 VSUBS 0.03283f
C692 VDD1.n4 VSUBS 0.014298f
C693 VDD1.n5 VSUBS 0.025848f
C694 VDD1.n6 VSUBS 0.014298f
C695 VDD1.n7 VSUBS 0.013889f
C696 VDD1.n8 VSUBS 0.03283f
C697 VDD1.n9 VSUBS 0.03283f
C698 VDD1.n10 VSUBS 0.014707f
C699 VDD1.n11 VSUBS 0.025848f
C700 VDD1.n12 VSUBS 0.013889f
C701 VDD1.n13 VSUBS 0.03283f
C702 VDD1.n14 VSUBS 0.014707f
C703 VDD1.n15 VSUBS 0.977694f
C704 VDD1.n16 VSUBS 0.013889f
C705 VDD1.t5 VSUBS 0.070567f
C706 VDD1.n17 VSUBS 0.173454f
C707 VDD1.n18 VSUBS 0.024696f
C708 VDD1.n19 VSUBS 0.024622f
C709 VDD1.n20 VSUBS 0.03283f
C710 VDD1.n21 VSUBS 0.014707f
C711 VDD1.n22 VSUBS 0.013889f
C712 VDD1.n23 VSUBS 0.025848f
C713 VDD1.n24 VSUBS 0.025848f
C714 VDD1.n25 VSUBS 0.013889f
C715 VDD1.n26 VSUBS 0.014707f
C716 VDD1.n27 VSUBS 0.03283f
C717 VDD1.n28 VSUBS 0.03283f
C718 VDD1.n29 VSUBS 0.014707f
C719 VDD1.n30 VSUBS 0.013889f
C720 VDD1.n31 VSUBS 0.025848f
C721 VDD1.n32 VSUBS 0.025848f
C722 VDD1.n33 VSUBS 0.013889f
C723 VDD1.n34 VSUBS 0.014707f
C724 VDD1.n35 VSUBS 0.03283f
C725 VDD1.n36 VSUBS 0.03283f
C726 VDD1.n37 VSUBS 0.014707f
C727 VDD1.n38 VSUBS 0.013889f
C728 VDD1.n39 VSUBS 0.025848f
C729 VDD1.n40 VSUBS 0.025848f
C730 VDD1.n41 VSUBS 0.013889f
C731 VDD1.n42 VSUBS 0.014707f
C732 VDD1.n43 VSUBS 0.03283f
C733 VDD1.n44 VSUBS 0.079855f
C734 VDD1.n45 VSUBS 0.014707f
C735 VDD1.n46 VSUBS 0.013889f
C736 VDD1.n47 VSUBS 0.066102f
C737 VDD1.n48 VSUBS 0.063422f
C738 VDD1.t0 VSUBS 0.19241f
C739 VDD1.t2 VSUBS 0.19241f
C740 VDD1.n49 VSUBS 1.44524f
C741 VDD1.n50 VSUBS 0.795124f
C742 VDD1.n51 VSUBS 0.028512f
C743 VDD1.n52 VSUBS 0.025848f
C744 VDD1.n53 VSUBS 0.013889f
C745 VDD1.n54 VSUBS 0.03283f
C746 VDD1.n55 VSUBS 0.014298f
C747 VDD1.n56 VSUBS 0.025848f
C748 VDD1.n57 VSUBS 0.014707f
C749 VDD1.n58 VSUBS 0.03283f
C750 VDD1.n59 VSUBS 0.014707f
C751 VDD1.n60 VSUBS 0.025848f
C752 VDD1.n61 VSUBS 0.013889f
C753 VDD1.n62 VSUBS 0.03283f
C754 VDD1.n63 VSUBS 0.014707f
C755 VDD1.n64 VSUBS 0.977694f
C756 VDD1.n65 VSUBS 0.013889f
C757 VDD1.t9 VSUBS 0.070567f
C758 VDD1.n66 VSUBS 0.173454f
C759 VDD1.n67 VSUBS 0.024696f
C760 VDD1.n68 VSUBS 0.024622f
C761 VDD1.n69 VSUBS 0.03283f
C762 VDD1.n70 VSUBS 0.014707f
C763 VDD1.n71 VSUBS 0.013889f
C764 VDD1.n72 VSUBS 0.025848f
C765 VDD1.n73 VSUBS 0.025848f
C766 VDD1.n74 VSUBS 0.013889f
C767 VDD1.n75 VSUBS 0.014707f
C768 VDD1.n76 VSUBS 0.03283f
C769 VDD1.n77 VSUBS 0.03283f
C770 VDD1.n78 VSUBS 0.014707f
C771 VDD1.n79 VSUBS 0.013889f
C772 VDD1.n80 VSUBS 0.025848f
C773 VDD1.n81 VSUBS 0.025848f
C774 VDD1.n82 VSUBS 0.013889f
C775 VDD1.n83 VSUBS 0.013889f
C776 VDD1.n84 VSUBS 0.014707f
C777 VDD1.n85 VSUBS 0.03283f
C778 VDD1.n86 VSUBS 0.03283f
C779 VDD1.n87 VSUBS 0.03283f
C780 VDD1.n88 VSUBS 0.014298f
C781 VDD1.n89 VSUBS 0.013889f
C782 VDD1.n90 VSUBS 0.025848f
C783 VDD1.n91 VSUBS 0.025848f
C784 VDD1.n92 VSUBS 0.013889f
C785 VDD1.n93 VSUBS 0.014707f
C786 VDD1.n94 VSUBS 0.03283f
C787 VDD1.n95 VSUBS 0.079855f
C788 VDD1.n96 VSUBS 0.014707f
C789 VDD1.n97 VSUBS 0.013889f
C790 VDD1.n98 VSUBS 0.066102f
C791 VDD1.n99 VSUBS 0.063422f
C792 VDD1.t1 VSUBS 0.19241f
C793 VDD1.t6 VSUBS 0.19241f
C794 VDD1.n100 VSUBS 1.44524f
C795 VDD1.n101 VSUBS 0.787476f
C796 VDD1.t8 VSUBS 0.19241f
C797 VDD1.t4 VSUBS 0.19241f
C798 VDD1.n102 VSUBS 1.45435f
C799 VDD1.n103 VSUBS 2.56301f
C800 VDD1.t3 VSUBS 0.19241f
C801 VDD1.t7 VSUBS 0.19241f
C802 VDD1.n104 VSUBS 1.44524f
C803 VDD1.n105 VSUBS 2.82863f
C804 VP.n0 VSUBS 0.041078f
C805 VP.t5 VSUBS 1.53771f
C806 VP.n1 VSUBS 0.054031f
C807 VP.n2 VSUBS 0.041078f
C808 VP.t1 VSUBS 1.53771f
C809 VP.n3 VSUBS 0.075023f
C810 VP.n4 VSUBS 0.041078f
C811 VP.t3 VSUBS 1.53771f
C812 VP.n5 VSUBS 0.066807f
C813 VP.n6 VSUBS 0.041078f
C814 VP.n7 VSUBS 0.046091f
C815 VP.n8 VSUBS 0.041078f
C816 VP.t2 VSUBS 1.53771f
C817 VP.n9 VSUBS 0.054031f
C818 VP.n10 VSUBS 0.041078f
C819 VP.t6 VSUBS 1.53771f
C820 VP.n11 VSUBS 0.075023f
C821 VP.n12 VSUBS 0.041078f
C822 VP.t7 VSUBS 1.53771f
C823 VP.n13 VSUBS 0.066807f
C824 VP.t4 VSUBS 1.65862f
C825 VP.t9 VSUBS 1.53771f
C826 VP.n14 VSUBS 0.647362f
C827 VP.n15 VSUBS 0.665608f
C828 VP.n16 VSUBS 0.255429f
C829 VP.n17 VSUBS 0.041078f
C830 VP.n18 VSUBS 0.038731f
C831 VP.n19 VSUBS 0.075023f
C832 VP.n20 VSUBS 0.607549f
C833 VP.n21 VSUBS 0.041078f
C834 VP.n22 VSUBS 0.041078f
C835 VP.n23 VSUBS 0.041078f
C836 VP.n24 VSUBS 0.038731f
C837 VP.n25 VSUBS 0.066807f
C838 VP.n26 VSUBS 0.568979f
C839 VP.n27 VSUBS 0.053612f
C840 VP.n28 VSUBS 0.041078f
C841 VP.n29 VSUBS 0.041078f
C842 VP.n30 VSUBS 0.041078f
C843 VP.n31 VSUBS 0.065396f
C844 VP.n32 VSUBS 0.046091f
C845 VP.n33 VSUBS 0.641567f
C846 VP.n34 VSUBS 1.8965f
C847 VP.t0 VSUBS 1.53771f
C848 VP.n35 VSUBS 0.641567f
C849 VP.n36 VSUBS 1.92952f
C850 VP.n37 VSUBS 0.041078f
C851 VP.n38 VSUBS 0.041078f
C852 VP.n39 VSUBS 0.065396f
C853 VP.n40 VSUBS 0.054031f
C854 VP.t8 VSUBS 1.53771f
C855 VP.n41 VSUBS 0.568979f
C856 VP.n42 VSUBS 0.053612f
C857 VP.n43 VSUBS 0.041078f
C858 VP.n44 VSUBS 0.041078f
C859 VP.n45 VSUBS 0.041078f
C860 VP.n46 VSUBS 0.038731f
C861 VP.n47 VSUBS 0.075023f
C862 VP.n48 VSUBS 0.607549f
C863 VP.n49 VSUBS 0.041078f
C864 VP.n50 VSUBS 0.041078f
C865 VP.n51 VSUBS 0.041078f
C866 VP.n52 VSUBS 0.038731f
C867 VP.n53 VSUBS 0.066807f
C868 VP.n54 VSUBS 0.568979f
C869 VP.n55 VSUBS 0.053612f
C870 VP.n56 VSUBS 0.041078f
C871 VP.n57 VSUBS 0.041078f
C872 VP.n58 VSUBS 0.041078f
C873 VP.n59 VSUBS 0.065396f
C874 VP.n60 VSUBS 0.046091f
C875 VP.n61 VSUBS 0.641567f
C876 VP.n62 VSUBS 0.040687f
C877 VTAIL.t12 VSUBS 0.217325f
C878 VTAIL.t9 VSUBS 0.217325f
C879 VTAIL.n0 VSUBS 1.50377f
C880 VTAIL.n1 VSUBS 0.830851f
C881 VTAIL.n2 VSUBS 0.032204f
C882 VTAIL.n3 VSUBS 0.029195f
C883 VTAIL.n4 VSUBS 0.015688f
C884 VTAIL.n5 VSUBS 0.037081f
C885 VTAIL.n6 VSUBS 0.016149f
C886 VTAIL.n7 VSUBS 0.029195f
C887 VTAIL.n8 VSUBS 0.016611f
C888 VTAIL.n9 VSUBS 0.037081f
C889 VTAIL.n10 VSUBS 0.016611f
C890 VTAIL.n11 VSUBS 0.029195f
C891 VTAIL.n12 VSUBS 0.015688f
C892 VTAIL.n13 VSUBS 0.037081f
C893 VTAIL.n14 VSUBS 0.016611f
C894 VTAIL.n15 VSUBS 1.1043f
C895 VTAIL.n16 VSUBS 0.015688f
C896 VTAIL.t6 VSUBS 0.079704f
C897 VTAIL.n17 VSUBS 0.195914f
C898 VTAIL.n18 VSUBS 0.027894f
C899 VTAIL.n19 VSUBS 0.027811f
C900 VTAIL.n20 VSUBS 0.037081f
C901 VTAIL.n21 VSUBS 0.016611f
C902 VTAIL.n22 VSUBS 0.015688f
C903 VTAIL.n23 VSUBS 0.029195f
C904 VTAIL.n24 VSUBS 0.029195f
C905 VTAIL.n25 VSUBS 0.015688f
C906 VTAIL.n26 VSUBS 0.016611f
C907 VTAIL.n27 VSUBS 0.037081f
C908 VTAIL.n28 VSUBS 0.037081f
C909 VTAIL.n29 VSUBS 0.016611f
C910 VTAIL.n30 VSUBS 0.015688f
C911 VTAIL.n31 VSUBS 0.029195f
C912 VTAIL.n32 VSUBS 0.029195f
C913 VTAIL.n33 VSUBS 0.015688f
C914 VTAIL.n34 VSUBS 0.015688f
C915 VTAIL.n35 VSUBS 0.016611f
C916 VTAIL.n36 VSUBS 0.037081f
C917 VTAIL.n37 VSUBS 0.037081f
C918 VTAIL.n38 VSUBS 0.037081f
C919 VTAIL.n39 VSUBS 0.016149f
C920 VTAIL.n40 VSUBS 0.015688f
C921 VTAIL.n41 VSUBS 0.029195f
C922 VTAIL.n42 VSUBS 0.029195f
C923 VTAIL.n43 VSUBS 0.015688f
C924 VTAIL.n44 VSUBS 0.016611f
C925 VTAIL.n45 VSUBS 0.037081f
C926 VTAIL.n46 VSUBS 0.090196f
C927 VTAIL.n47 VSUBS 0.016611f
C928 VTAIL.n48 VSUBS 0.015688f
C929 VTAIL.n49 VSUBS 0.074661f
C930 VTAIL.n50 VSUBS 0.045588f
C931 VTAIL.n51 VSUBS 0.292154f
C932 VTAIL.t5 VSUBS 0.217325f
C933 VTAIL.t19 VSUBS 0.217325f
C934 VTAIL.n52 VSUBS 1.50377f
C935 VTAIL.n53 VSUBS 0.89066f
C936 VTAIL.t8 VSUBS 0.217325f
C937 VTAIL.t2 VSUBS 0.217325f
C938 VTAIL.n54 VSUBS 1.50377f
C939 VTAIL.n55 VSUBS 2.19714f
C940 VTAIL.t15 VSUBS 0.217325f
C941 VTAIL.t11 VSUBS 0.217325f
C942 VTAIL.n56 VSUBS 1.50378f
C943 VTAIL.n57 VSUBS 2.19713f
C944 VTAIL.t10 VSUBS 0.217325f
C945 VTAIL.t17 VSUBS 0.217325f
C946 VTAIL.n58 VSUBS 1.50378f
C947 VTAIL.n59 VSUBS 0.89065f
C948 VTAIL.n60 VSUBS 0.032204f
C949 VTAIL.n61 VSUBS 0.029195f
C950 VTAIL.n62 VSUBS 0.015688f
C951 VTAIL.n63 VSUBS 0.037081f
C952 VTAIL.n64 VSUBS 0.016149f
C953 VTAIL.n65 VSUBS 0.029195f
C954 VTAIL.n66 VSUBS 0.016149f
C955 VTAIL.n67 VSUBS 0.015688f
C956 VTAIL.n68 VSUBS 0.037081f
C957 VTAIL.n69 VSUBS 0.037081f
C958 VTAIL.n70 VSUBS 0.016611f
C959 VTAIL.n71 VSUBS 0.029195f
C960 VTAIL.n72 VSUBS 0.015688f
C961 VTAIL.n73 VSUBS 0.037081f
C962 VTAIL.n74 VSUBS 0.016611f
C963 VTAIL.n75 VSUBS 1.1043f
C964 VTAIL.n76 VSUBS 0.015688f
C965 VTAIL.t13 VSUBS 0.079704f
C966 VTAIL.n77 VSUBS 0.195914f
C967 VTAIL.n78 VSUBS 0.027894f
C968 VTAIL.n79 VSUBS 0.027811f
C969 VTAIL.n80 VSUBS 0.037081f
C970 VTAIL.n81 VSUBS 0.016611f
C971 VTAIL.n82 VSUBS 0.015688f
C972 VTAIL.n83 VSUBS 0.029195f
C973 VTAIL.n84 VSUBS 0.029195f
C974 VTAIL.n85 VSUBS 0.015688f
C975 VTAIL.n86 VSUBS 0.016611f
C976 VTAIL.n87 VSUBS 0.037081f
C977 VTAIL.n88 VSUBS 0.037081f
C978 VTAIL.n89 VSUBS 0.016611f
C979 VTAIL.n90 VSUBS 0.015688f
C980 VTAIL.n91 VSUBS 0.029195f
C981 VTAIL.n92 VSUBS 0.029195f
C982 VTAIL.n93 VSUBS 0.015688f
C983 VTAIL.n94 VSUBS 0.016611f
C984 VTAIL.n95 VSUBS 0.037081f
C985 VTAIL.n96 VSUBS 0.037081f
C986 VTAIL.n97 VSUBS 0.016611f
C987 VTAIL.n98 VSUBS 0.015688f
C988 VTAIL.n99 VSUBS 0.029195f
C989 VTAIL.n100 VSUBS 0.029195f
C990 VTAIL.n101 VSUBS 0.015688f
C991 VTAIL.n102 VSUBS 0.016611f
C992 VTAIL.n103 VSUBS 0.037081f
C993 VTAIL.n104 VSUBS 0.090196f
C994 VTAIL.n105 VSUBS 0.016611f
C995 VTAIL.n106 VSUBS 0.015688f
C996 VTAIL.n107 VSUBS 0.074661f
C997 VTAIL.n108 VSUBS 0.045588f
C998 VTAIL.n109 VSUBS 0.292154f
C999 VTAIL.t3 VSUBS 0.217325f
C1000 VTAIL.t7 VSUBS 0.217325f
C1001 VTAIL.n110 VSUBS 1.50378f
C1002 VTAIL.n111 VSUBS 0.861861f
C1003 VTAIL.t1 VSUBS 0.217325f
C1004 VTAIL.t0 VSUBS 0.217325f
C1005 VTAIL.n112 VSUBS 1.50378f
C1006 VTAIL.n113 VSUBS 0.89065f
C1007 VTAIL.n114 VSUBS 0.032204f
C1008 VTAIL.n115 VSUBS 0.029195f
C1009 VTAIL.n116 VSUBS 0.015688f
C1010 VTAIL.n117 VSUBS 0.037081f
C1011 VTAIL.n118 VSUBS 0.016149f
C1012 VTAIL.n119 VSUBS 0.029195f
C1013 VTAIL.n120 VSUBS 0.016149f
C1014 VTAIL.n121 VSUBS 0.015688f
C1015 VTAIL.n122 VSUBS 0.037081f
C1016 VTAIL.n123 VSUBS 0.037081f
C1017 VTAIL.n124 VSUBS 0.016611f
C1018 VTAIL.n125 VSUBS 0.029195f
C1019 VTAIL.n126 VSUBS 0.015688f
C1020 VTAIL.n127 VSUBS 0.037081f
C1021 VTAIL.n128 VSUBS 0.016611f
C1022 VTAIL.n129 VSUBS 1.1043f
C1023 VTAIL.n130 VSUBS 0.015688f
C1024 VTAIL.t4 VSUBS 0.079704f
C1025 VTAIL.n131 VSUBS 0.195914f
C1026 VTAIL.n132 VSUBS 0.027894f
C1027 VTAIL.n133 VSUBS 0.027811f
C1028 VTAIL.n134 VSUBS 0.037081f
C1029 VTAIL.n135 VSUBS 0.016611f
C1030 VTAIL.n136 VSUBS 0.015688f
C1031 VTAIL.n137 VSUBS 0.029195f
C1032 VTAIL.n138 VSUBS 0.029195f
C1033 VTAIL.n139 VSUBS 0.015688f
C1034 VTAIL.n140 VSUBS 0.016611f
C1035 VTAIL.n141 VSUBS 0.037081f
C1036 VTAIL.n142 VSUBS 0.037081f
C1037 VTAIL.n143 VSUBS 0.016611f
C1038 VTAIL.n144 VSUBS 0.015688f
C1039 VTAIL.n145 VSUBS 0.029195f
C1040 VTAIL.n146 VSUBS 0.029195f
C1041 VTAIL.n147 VSUBS 0.015688f
C1042 VTAIL.n148 VSUBS 0.016611f
C1043 VTAIL.n149 VSUBS 0.037081f
C1044 VTAIL.n150 VSUBS 0.037081f
C1045 VTAIL.n151 VSUBS 0.016611f
C1046 VTAIL.n152 VSUBS 0.015688f
C1047 VTAIL.n153 VSUBS 0.029195f
C1048 VTAIL.n154 VSUBS 0.029195f
C1049 VTAIL.n155 VSUBS 0.015688f
C1050 VTAIL.n156 VSUBS 0.016611f
C1051 VTAIL.n157 VSUBS 0.037081f
C1052 VTAIL.n158 VSUBS 0.090196f
C1053 VTAIL.n159 VSUBS 0.016611f
C1054 VTAIL.n160 VSUBS 0.015688f
C1055 VTAIL.n161 VSUBS 0.074661f
C1056 VTAIL.n162 VSUBS 0.045588f
C1057 VTAIL.n163 VSUBS 1.48145f
C1058 VTAIL.n164 VSUBS 0.032204f
C1059 VTAIL.n165 VSUBS 0.029195f
C1060 VTAIL.n166 VSUBS 0.015688f
C1061 VTAIL.n167 VSUBS 0.037081f
C1062 VTAIL.n168 VSUBS 0.016149f
C1063 VTAIL.n169 VSUBS 0.029195f
C1064 VTAIL.n170 VSUBS 0.016611f
C1065 VTAIL.n171 VSUBS 0.037081f
C1066 VTAIL.n172 VSUBS 0.016611f
C1067 VTAIL.n173 VSUBS 0.029195f
C1068 VTAIL.n174 VSUBS 0.015688f
C1069 VTAIL.n175 VSUBS 0.037081f
C1070 VTAIL.n176 VSUBS 0.016611f
C1071 VTAIL.n177 VSUBS 1.1043f
C1072 VTAIL.n178 VSUBS 0.015688f
C1073 VTAIL.t16 VSUBS 0.079704f
C1074 VTAIL.n179 VSUBS 0.195914f
C1075 VTAIL.n180 VSUBS 0.027894f
C1076 VTAIL.n181 VSUBS 0.027811f
C1077 VTAIL.n182 VSUBS 0.037081f
C1078 VTAIL.n183 VSUBS 0.016611f
C1079 VTAIL.n184 VSUBS 0.015688f
C1080 VTAIL.n185 VSUBS 0.029195f
C1081 VTAIL.n186 VSUBS 0.029195f
C1082 VTAIL.n187 VSUBS 0.015688f
C1083 VTAIL.n188 VSUBS 0.016611f
C1084 VTAIL.n189 VSUBS 0.037081f
C1085 VTAIL.n190 VSUBS 0.037081f
C1086 VTAIL.n191 VSUBS 0.016611f
C1087 VTAIL.n192 VSUBS 0.015688f
C1088 VTAIL.n193 VSUBS 0.029195f
C1089 VTAIL.n194 VSUBS 0.029195f
C1090 VTAIL.n195 VSUBS 0.015688f
C1091 VTAIL.n196 VSUBS 0.015688f
C1092 VTAIL.n197 VSUBS 0.016611f
C1093 VTAIL.n198 VSUBS 0.037081f
C1094 VTAIL.n199 VSUBS 0.037081f
C1095 VTAIL.n200 VSUBS 0.037081f
C1096 VTAIL.n201 VSUBS 0.016149f
C1097 VTAIL.n202 VSUBS 0.015688f
C1098 VTAIL.n203 VSUBS 0.029195f
C1099 VTAIL.n204 VSUBS 0.029195f
C1100 VTAIL.n205 VSUBS 0.015688f
C1101 VTAIL.n206 VSUBS 0.016611f
C1102 VTAIL.n207 VSUBS 0.037081f
C1103 VTAIL.n208 VSUBS 0.090196f
C1104 VTAIL.n209 VSUBS 0.016611f
C1105 VTAIL.n210 VSUBS 0.015688f
C1106 VTAIL.n211 VSUBS 0.074661f
C1107 VTAIL.n212 VSUBS 0.045588f
C1108 VTAIL.n213 VSUBS 1.48145f
C1109 VTAIL.t14 VSUBS 0.217325f
C1110 VTAIL.t18 VSUBS 0.217325f
C1111 VTAIL.n214 VSUBS 1.50377f
C1112 VTAIL.n215 VSUBS 0.775706f
C1113 VDD2.n0 VSUBS 0.028356f
C1114 VDD2.n1 VSUBS 0.025706f
C1115 VDD2.n2 VSUBS 0.013814f
C1116 VDD2.n3 VSUBS 0.03265f
C1117 VDD2.n4 VSUBS 0.01422f
C1118 VDD2.n5 VSUBS 0.025706f
C1119 VDD2.n6 VSUBS 0.014626f
C1120 VDD2.n7 VSUBS 0.03265f
C1121 VDD2.n8 VSUBS 0.014626f
C1122 VDD2.n9 VSUBS 0.025706f
C1123 VDD2.n10 VSUBS 0.013814f
C1124 VDD2.n11 VSUBS 0.03265f
C1125 VDD2.n12 VSUBS 0.014626f
C1126 VDD2.n13 VSUBS 0.972345f
C1127 VDD2.n14 VSUBS 0.013814f
C1128 VDD2.t9 VSUBS 0.070181f
C1129 VDD2.n15 VSUBS 0.172505f
C1130 VDD2.n16 VSUBS 0.024561f
C1131 VDD2.n17 VSUBS 0.024487f
C1132 VDD2.n18 VSUBS 0.03265f
C1133 VDD2.n19 VSUBS 0.014626f
C1134 VDD2.n20 VSUBS 0.013814f
C1135 VDD2.n21 VSUBS 0.025706f
C1136 VDD2.n22 VSUBS 0.025706f
C1137 VDD2.n23 VSUBS 0.013814f
C1138 VDD2.n24 VSUBS 0.014626f
C1139 VDD2.n25 VSUBS 0.03265f
C1140 VDD2.n26 VSUBS 0.03265f
C1141 VDD2.n27 VSUBS 0.014626f
C1142 VDD2.n28 VSUBS 0.013814f
C1143 VDD2.n29 VSUBS 0.025706f
C1144 VDD2.n30 VSUBS 0.025706f
C1145 VDD2.n31 VSUBS 0.013814f
C1146 VDD2.n32 VSUBS 0.013814f
C1147 VDD2.n33 VSUBS 0.014626f
C1148 VDD2.n34 VSUBS 0.03265f
C1149 VDD2.n35 VSUBS 0.03265f
C1150 VDD2.n36 VSUBS 0.03265f
C1151 VDD2.n37 VSUBS 0.01422f
C1152 VDD2.n38 VSUBS 0.013814f
C1153 VDD2.n39 VSUBS 0.025706f
C1154 VDD2.n40 VSUBS 0.025706f
C1155 VDD2.n41 VSUBS 0.013814f
C1156 VDD2.n42 VSUBS 0.014626f
C1157 VDD2.n43 VSUBS 0.03265f
C1158 VDD2.n44 VSUBS 0.079418f
C1159 VDD2.n45 VSUBS 0.014626f
C1160 VDD2.n46 VSUBS 0.013814f
C1161 VDD2.n47 VSUBS 0.06574f
C1162 VDD2.n48 VSUBS 0.063075f
C1163 VDD2.t7 VSUBS 0.191357f
C1164 VDD2.t5 VSUBS 0.191357f
C1165 VDD2.n49 VSUBS 1.43733f
C1166 VDD2.n50 VSUBS 0.783168f
C1167 VDD2.t3 VSUBS 0.191357f
C1168 VDD2.t8 VSUBS 0.191357f
C1169 VDD2.n51 VSUBS 1.44639f
C1170 VDD2.n52 VSUBS 2.45205f
C1171 VDD2.n53 VSUBS 0.028356f
C1172 VDD2.n54 VSUBS 0.025706f
C1173 VDD2.n55 VSUBS 0.013814f
C1174 VDD2.n56 VSUBS 0.03265f
C1175 VDD2.n57 VSUBS 0.01422f
C1176 VDD2.n58 VSUBS 0.025706f
C1177 VDD2.n59 VSUBS 0.01422f
C1178 VDD2.n60 VSUBS 0.013814f
C1179 VDD2.n61 VSUBS 0.03265f
C1180 VDD2.n62 VSUBS 0.03265f
C1181 VDD2.n63 VSUBS 0.014626f
C1182 VDD2.n64 VSUBS 0.025706f
C1183 VDD2.n65 VSUBS 0.013814f
C1184 VDD2.n66 VSUBS 0.03265f
C1185 VDD2.n67 VSUBS 0.014626f
C1186 VDD2.n68 VSUBS 0.972345f
C1187 VDD2.n69 VSUBS 0.013814f
C1188 VDD2.t6 VSUBS 0.070181f
C1189 VDD2.n70 VSUBS 0.172505f
C1190 VDD2.n71 VSUBS 0.024561f
C1191 VDD2.n72 VSUBS 0.024487f
C1192 VDD2.n73 VSUBS 0.03265f
C1193 VDD2.n74 VSUBS 0.014626f
C1194 VDD2.n75 VSUBS 0.013814f
C1195 VDD2.n76 VSUBS 0.025706f
C1196 VDD2.n77 VSUBS 0.025706f
C1197 VDD2.n78 VSUBS 0.013814f
C1198 VDD2.n79 VSUBS 0.014626f
C1199 VDD2.n80 VSUBS 0.03265f
C1200 VDD2.n81 VSUBS 0.03265f
C1201 VDD2.n82 VSUBS 0.014626f
C1202 VDD2.n83 VSUBS 0.013814f
C1203 VDD2.n84 VSUBS 0.025706f
C1204 VDD2.n85 VSUBS 0.025706f
C1205 VDD2.n86 VSUBS 0.013814f
C1206 VDD2.n87 VSUBS 0.014626f
C1207 VDD2.n88 VSUBS 0.03265f
C1208 VDD2.n89 VSUBS 0.03265f
C1209 VDD2.n90 VSUBS 0.014626f
C1210 VDD2.n91 VSUBS 0.013814f
C1211 VDD2.n92 VSUBS 0.025706f
C1212 VDD2.n93 VSUBS 0.025706f
C1213 VDD2.n94 VSUBS 0.013814f
C1214 VDD2.n95 VSUBS 0.014626f
C1215 VDD2.n96 VSUBS 0.03265f
C1216 VDD2.n97 VSUBS 0.079418f
C1217 VDD2.n98 VSUBS 0.014626f
C1218 VDD2.n99 VSUBS 0.013814f
C1219 VDD2.n100 VSUBS 0.06574f
C1220 VDD2.n101 VSUBS 0.057846f
C1221 VDD2.n102 VSUBS 2.31746f
C1222 VDD2.t0 VSUBS 0.191357f
C1223 VDD2.t2 VSUBS 0.191357f
C1224 VDD2.n103 VSUBS 1.43734f
C1225 VDD2.n104 VSUBS 0.614351f
C1226 VDD2.t1 VSUBS 0.191357f
C1227 VDD2.t4 VSUBS 0.191357f
C1228 VDD2.n105 VSUBS 1.44636f
C1229 VN.n0 VSUBS 0.039977f
C1230 VN.t2 VSUBS 1.49648f
C1231 VN.n1 VSUBS 0.052582f
C1232 VN.n2 VSUBS 0.039977f
C1233 VN.t0 VSUBS 1.49648f
C1234 VN.n3 VSUBS 0.073012f
C1235 VN.n4 VSUBS 0.039977f
C1236 VN.t4 VSUBS 1.49648f
C1237 VN.n5 VSUBS 0.065015f
C1238 VN.t6 VSUBS 1.61414f
C1239 VN.t9 VSUBS 1.49648f
C1240 VN.n6 VSUBS 0.630003f
C1241 VN.n7 VSUBS 0.64776f
C1242 VN.n8 VSUBS 0.24858f
C1243 VN.n9 VSUBS 0.039977f
C1244 VN.n10 VSUBS 0.037692f
C1245 VN.n11 VSUBS 0.073012f
C1246 VN.n12 VSUBS 0.591257f
C1247 VN.n13 VSUBS 0.039977f
C1248 VN.n14 VSUBS 0.039977f
C1249 VN.n15 VSUBS 0.039977f
C1250 VN.n16 VSUBS 0.037692f
C1251 VN.n17 VSUBS 0.065015f
C1252 VN.n18 VSUBS 0.553722f
C1253 VN.n19 VSUBS 0.052175f
C1254 VN.n20 VSUBS 0.039977f
C1255 VN.n21 VSUBS 0.039977f
C1256 VN.n22 VSUBS 0.039977f
C1257 VN.n23 VSUBS 0.063643f
C1258 VN.n24 VSUBS 0.044855f
C1259 VN.n25 VSUBS 0.624363f
C1260 VN.n26 VSUBS 0.039596f
C1261 VN.n27 VSUBS 0.039977f
C1262 VN.t3 VSUBS 1.49648f
C1263 VN.n28 VSUBS 0.052582f
C1264 VN.n29 VSUBS 0.039977f
C1265 VN.t7 VSUBS 1.49648f
C1266 VN.n30 VSUBS 0.073012f
C1267 VN.n31 VSUBS 0.039977f
C1268 VN.t8 VSUBS 1.49648f
C1269 VN.n32 VSUBS 0.065015f
C1270 VN.t5 VSUBS 1.61414f
C1271 VN.t1 VSUBS 1.49648f
C1272 VN.n33 VSUBS 0.630003f
C1273 VN.n34 VSUBS 0.64776f
C1274 VN.n35 VSUBS 0.24858f
C1275 VN.n36 VSUBS 0.039977f
C1276 VN.n37 VSUBS 0.037692f
C1277 VN.n38 VSUBS 0.073012f
C1278 VN.n39 VSUBS 0.591257f
C1279 VN.n40 VSUBS 0.039977f
C1280 VN.n41 VSUBS 0.039977f
C1281 VN.n42 VSUBS 0.039977f
C1282 VN.n43 VSUBS 0.037692f
C1283 VN.n44 VSUBS 0.065015f
C1284 VN.n45 VSUBS 0.553722f
C1285 VN.n46 VSUBS 0.052175f
C1286 VN.n47 VSUBS 0.039977f
C1287 VN.n48 VSUBS 0.039977f
C1288 VN.n49 VSUBS 0.039977f
C1289 VN.n50 VSUBS 0.063643f
C1290 VN.n51 VSUBS 0.044855f
C1291 VN.n52 VSUBS 0.624363f
C1292 VN.n53 VSUBS 1.87179f
.ends

