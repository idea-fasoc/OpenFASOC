* NGSPICE file created from tg_sample_0003.ext - technology: sky130A

.subckt tg_sample_0003 VIN VGN VGP VSS VCC VOUT
X0 VIN.t3 VGN.t0 VOUT.t2 VSS.t1 sky130_fd_pr__nfet_01v8 ad=1.1037 pd=6.44 as=0.46695 ps=3.16 w=2.83 l=1.42
X1 VCC.t9 VCC.t6 VCC.t8 VCC.t7 sky130_fd_pr__pfet_01v8 ad=1.8135 pd=10.08 as=0 ps=0 w=4.65 l=1.5
X2 VSS.t9 VSS.t6 VSS.t8 VSS.t7 sky130_fd_pr__nfet_01v8 ad=1.1037 pd=6.44 as=0 ps=0 w=2.83 l=1.42
X3 VOUT.t3 VGN.t1 VIN.t2 VSS.t0 sky130_fd_pr__nfet_01v8 ad=0.46695 pd=3.16 as=1.1037 ps=6.44 w=2.83 l=1.42
X4 VOUT.t0 VGP.t0 VIN.t0 VCC.t0 sky130_fd_pr__pfet_01v8 ad=0.76725 pd=4.98 as=1.8135 ps=10.08 w=4.65 l=1.5
X5 VSS.t5 VSS.t2 VSS.t4 VSS.t3 sky130_fd_pr__nfet_01v8 ad=1.1037 pd=6.44 as=0 ps=0 w=2.83 l=1.42
X6 VCC.t5 VCC.t2 VCC.t4 VCC.t3 sky130_fd_pr__pfet_01v8 ad=1.8135 pd=10.08 as=0 ps=0 w=4.65 l=1.5
X7 VIN.t1 VGP.t1 VOUT.t1 VCC.t1 sky130_fd_pr__pfet_01v8 ad=1.8135 pd=10.08 as=0.76725 ps=4.98 w=4.65 l=1.5
R0 VGN.n0 VGN.t1 83.207
R1 VGN.n0 VGN.t0 82.8977
R2 VGN VGN.n0 13.3738
R3 VOUT VOUT.n0 106.734
R4 VOUT VOUT.n1 93.7336
R5 VOUT.n1 VOUT.t2 6.99697
R6 VOUT.n1 VOUT.t3 6.99697
R7 VOUT.n0 VOUT.t1 6.99082
R8 VOUT.n0 VOUT.t0 6.99082
R9 VIN.n18 VIN.n0 756.745
R10 VIN.n41 VIN.n23 756.745
R11 VIN.n9 VIN.n8 585
R12 VIN.n11 VIN.n10 585
R13 VIN.n4 VIN.n3 585
R14 VIN.n17 VIN.n16 585
R15 VIN.n19 VIN.n18 585
R16 VIN.n32 VIN.n31 585
R17 VIN.n34 VIN.n33 585
R18 VIN.n27 VIN.n26 585
R19 VIN.n40 VIN.n39 585
R20 VIN.n42 VIN.n41 585
R21 VIN.n7 VIN.t0 328.587
R22 VIN.n30 VIN.t1 328.587
R23 VIN.n10 VIN.n9 171.744
R24 VIN.n10 VIN.n3 171.744
R25 VIN.n17 VIN.n3 171.744
R26 VIN.n18 VIN.n17 171.744
R27 VIN.n33 VIN.n32 171.744
R28 VIN.n33 VIN.n26 171.744
R29 VIN.n40 VIN.n26 171.744
R30 VIN.n41 VIN.n40 171.744
R31 VIN.n9 VIN.t0 85.8723
R32 VIN.n32 VIN.t1 85.8723
R33 VIN.n47 VIN.t2 74.0125
R34 VIN.n47 VIN.t3 72.5038
R35 VIN.n46 VIN.n22 35.5084
R36 VIN.n46 VIN.n45 33.9308
R37 VIN.n8 VIN.n7 16.3651
R38 VIN.n31 VIN.n30 16.3651
R39 VIN.n11 VIN.n6 12.8005
R40 VIN.n34 VIN.n29 12.8005
R41 VIN.n12 VIN.n4 12.0247
R42 VIN.n35 VIN.n27 12.0247
R43 VIN VIN.n46 11.4014
R44 VIN.n16 VIN.n15 11.249
R45 VIN.n39 VIN.n38 11.249
R46 VIN.n19 VIN.n2 10.4732
R47 VIN.n42 VIN.n25 10.4732
R48 VIN.n20 VIN.n0 9.69747
R49 VIN.n43 VIN.n23 9.69747
R50 VIN.n22 VIN.n21 9.45567
R51 VIN.n45 VIN.n44 9.45567
R52 VIN.n21 VIN.n20 9.3005
R53 VIN.n2 VIN.n1 9.3005
R54 VIN.n15 VIN.n14 9.3005
R55 VIN.n13 VIN.n12 9.3005
R56 VIN.n6 VIN.n5 9.3005
R57 VIN.n44 VIN.n43 9.3005
R58 VIN.n25 VIN.n24 9.3005
R59 VIN.n38 VIN.n37 9.3005
R60 VIN.n36 VIN.n35 9.3005
R61 VIN.n29 VIN.n28 9.3005
R62 VIN.n22 VIN.n0 4.26717
R63 VIN.n45 VIN.n23 4.26717
R64 VIN.n7 VIN.n5 3.73474
R65 VIN.n30 VIN.n28 3.73474
R66 VIN.n20 VIN.n19 3.49141
R67 VIN.n43 VIN.n42 3.49141
R68 VIN.n16 VIN.n2 2.71565
R69 VIN.n39 VIN.n25 2.71565
R70 VIN.n15 VIN.n4 1.93989
R71 VIN.n38 VIN.n27 1.93989
R72 VIN.n12 VIN.n11 1.16414
R73 VIN.n35 VIN.n34 1.16414
R74 VIN.n8 VIN.n6 0.388379
R75 VIN.n31 VIN.n29 0.388379
R76 VIN.n13 VIN.n5 0.155672
R77 VIN.n14 VIN.n13 0.155672
R78 VIN.n14 VIN.n1 0.155672
R79 VIN.n21 VIN.n1 0.155672
R80 VIN.n36 VIN.n28 0.155672
R81 VIN.n37 VIN.n36 0.155672
R82 VIN.n37 VIN.n24 0.155672
R83 VIN.n44 VIN.n24 0.155672
R84 VIN VIN.n47 0.00481034
R85 VSS.n104 VSS.n60 689.5
R86 VSS.n102 VSS.n62 689.5
R87 VSS.n204 VSS.n18 689.5
R88 VSS.n206 VSS.n14 689.5
R89 VSS.n105 VSS.n104 585
R90 VSS.n104 VSS.n103 585
R91 VSS.n58 VSS.n57 585
R92 VSS.n57 VSS.n56 585
R93 VSS.n110 VSS.n109 585
R94 VSS.n111 VSS.n110 585
R95 VSS.n49 VSS.n48 585
R96 VSS.n50 VSS.n49 585
R97 VSS.n121 VSS.n120 585
R98 VSS.n120 VSS.n119 585
R99 VSS.n45 VSS.n43 585
R100 VSS.n43 VSS.n41 585
R101 VSS.n127 VSS.n126 585
R102 VSS.n128 VSS.n127 585
R103 VSS.n46 VSS.n44 585
R104 VSS.n44 VSS.n42 585
R105 VSS.n34 VSS.n33 585
R106 VSS.n35 VSS.n34 585
R107 VSS.n139 VSS.n138 585
R108 VSS.n138 VSS.n137 585
R109 VSS.n31 VSS.n30 585
R110 VSS.n30 VSS.n29 585
R111 VSS.n144 VSS.n143 585
R112 VSS.n145 VSS.n144 585
R113 VSS.n28 VSS.n27 585
R114 VSS.n146 VSS.n28 585
R115 VSS.n150 VSS.n149 585
R116 VSS.n149 VSS.n148 585
R117 VSS.n25 VSS.n24 585
R118 VSS.n24 VSS.n23 585
R119 VSS.n155 VSS.n154 585
R120 VSS.n156 VSS.n155 585
R121 VSS.n22 VSS.n21 585
R122 VSS.n157 VSS.n22 585
R123 VSS.n161 VSS.n160 585
R124 VSS.n160 VSS.n159 585
R125 VSS.n19 VSS.n17 585
R126 VSS.n17 VSS.n15 585
R127 VSS.n204 VSS.n203 585
R128 VSS.n205 VSS.n204 585
R129 VSS.n207 VSS.n206 585
R130 VSS.n206 VSS.n205 585
R131 VSS.n208 VSS.n13 585
R132 VSS.n15 VSS.n13 585
R133 VSS.n158 VSS.n11 585
R134 VSS.n159 VSS.n158 585
R135 VSS.n212 VSS.n10 585
R136 VSS.n157 VSS.n10 585
R137 VSS.n213 VSS.n9 585
R138 VSS.n156 VSS.n9 585
R139 VSS.n214 VSS.n8 585
R140 VSS.n23 VSS.n8 585
R141 VSS.n147 VSS.n6 585
R142 VSS.n148 VSS.n147 585
R143 VSS.n218 VSS.n5 585
R144 VSS.n146 VSS.n5 585
R145 VSS.n219 VSS.n4 585
R146 VSS.n145 VSS.n4 585
R147 VSS.n220 VSS.n3 585
R148 VSS.n29 VSS.n3 585
R149 VSS.n136 VSS.n2 585
R150 VSS.n137 VSS.n136 585
R151 VSS.n135 VSS.n134 585
R152 VSS.n135 VSS.n35 585
R153 VSS.n37 VSS.n36 585
R154 VSS.n42 VSS.n36 585
R155 VSS.n130 VSS.n129 585
R156 VSS.n129 VSS.n128 585
R157 VSS.n40 VSS.n39 585
R158 VSS.n41 VSS.n40 585
R159 VSS.n118 VSS.n117 585
R160 VSS.n119 VSS.n118 585
R161 VSS.n52 VSS.n51 585
R162 VSS.n51 VSS.n50 585
R163 VSS.n113 VSS.n112 585
R164 VSS.n112 VSS.n111 585
R165 VSS.n55 VSS.n54 585
R166 VSS.n56 VSS.n55 585
R167 VSS.n102 VSS.n101 585
R168 VSS.n103 VSS.n102 585
R169 VSS.n176 VSS.n14 585
R170 VSS.n177 VSS.n173 585
R171 VSS.n180 VSS.n179 585
R172 VSS.n182 VSS.n170 585
R173 VSS.n184 VSS.n183 585
R174 VSS.n185 VSS.n169 585
R175 VSS.n187 VSS.n186 585
R176 VSS.n189 VSS.n167 585
R177 VSS.n191 VSS.n190 585
R178 VSS.n192 VSS.n166 585
R179 VSS.n194 VSS.n193 585
R180 VSS.n196 VSS.n165 585
R181 VSS.n197 VSS.n164 585
R182 VSS.n200 VSS.n199 585
R183 VSS.n201 VSS.n18 585
R184 VSS.n18 VSS.n16 585
R185 VSS.n60 VSS.n59 585
R186 VSS.n74 VSS.n73 585
R187 VSS.n75 VSS.n71 585
R188 VSS.n71 VSS.n61 585
R189 VSS.n77 VSS.n76 585
R190 VSS.n79 VSS.n70 585
R191 VSS.n82 VSS.n81 585
R192 VSS.n83 VSS.n69 585
R193 VSS.n85 VSS.n84 585
R194 VSS.n87 VSS.n68 585
R195 VSS.n90 VSS.n89 585
R196 VSS.n91 VSS.n67 585
R197 VSS.n93 VSS.n92 585
R198 VSS.n95 VSS.n66 585
R199 VSS.n98 VSS.n97 585
R200 VSS.n99 VSS.n62 585
R201 VSS.n103 VSS.n61 554.447
R202 VSS.n205 VSS.n16 554.447
R203 VSS.n103 VSS.n56 296.497
R204 VSS.n111 VSS.n56 296.497
R205 VSS.n119 VSS.n50 296.497
R206 VSS.n119 VSS.n41 296.497
R207 VSS.n128 VSS.n41 296.497
R208 VSS.n128 VSS.n42 296.497
R209 VSS.n137 VSS.n35 296.497
R210 VSS.n137 VSS.n29 296.497
R211 VSS.n145 VSS.n29 296.497
R212 VSS.n148 VSS.n146 296.497
R213 VSS.n148 VSS.n23 296.497
R214 VSS.n156 VSS.n23 296.497
R215 VSS.n157 VSS.n156 296.497
R216 VSS.n159 VSS.n15 296.497
R217 VSS.n205 VSS.n15 296.497
R218 VSS.t7 VSS.n50 275.741
R219 VSS.t3 VSS.n157 275.741
R220 VSS.n172 VSS.n16 256.663
R221 VSS.n181 VSS.n16 256.663
R222 VSS.n171 VSS.n16 256.663
R223 VSS.n188 VSS.n16 256.663
R224 VSS.n168 VSS.n16 256.663
R225 VSS.n195 VSS.n16 256.663
R226 VSS.n198 VSS.n16 256.663
R227 VSS.n72 VSS.n61 256.663
R228 VSS.n78 VSS.n61 256.663
R229 VSS.n80 VSS.n61 256.663
R230 VSS.n86 VSS.n61 256.663
R231 VSS.n88 VSS.n61 256.663
R232 VSS.n94 VSS.n61 256.663
R233 VSS.n96 VSS.n61 256.663
R234 VSS.n174 VSS.t2 253.16
R235 VSS.n63 VSS.t6 253.16
R236 VSS.n104 VSS.n57 240.244
R237 VSS.n110 VSS.n57 240.244
R238 VSS.n110 VSS.n49 240.244
R239 VSS.n120 VSS.n49 240.244
R240 VSS.n120 VSS.n43 240.244
R241 VSS.n127 VSS.n43 240.244
R242 VSS.n127 VSS.n44 240.244
R243 VSS.n44 VSS.n34 240.244
R244 VSS.n138 VSS.n34 240.244
R245 VSS.n138 VSS.n30 240.244
R246 VSS.n144 VSS.n30 240.244
R247 VSS.n144 VSS.n28 240.244
R248 VSS.n149 VSS.n28 240.244
R249 VSS.n149 VSS.n24 240.244
R250 VSS.n155 VSS.n24 240.244
R251 VSS.n155 VSS.n22 240.244
R252 VSS.n160 VSS.n22 240.244
R253 VSS.n160 VSS.n17 240.244
R254 VSS.n204 VSS.n17 240.244
R255 VSS.n102 VSS.n55 240.244
R256 VSS.n112 VSS.n55 240.244
R257 VSS.n112 VSS.n51 240.244
R258 VSS.n118 VSS.n51 240.244
R259 VSS.n118 VSS.n40 240.244
R260 VSS.n129 VSS.n40 240.244
R261 VSS.n129 VSS.n36 240.244
R262 VSS.n135 VSS.n36 240.244
R263 VSS.n136 VSS.n135 240.244
R264 VSS.n136 VSS.n3 240.244
R265 VSS.n4 VSS.n3 240.244
R266 VSS.n5 VSS.n4 240.244
R267 VSS.n147 VSS.n5 240.244
R268 VSS.n147 VSS.n8 240.244
R269 VSS.n9 VSS.n8 240.244
R270 VSS.n10 VSS.n9 240.244
R271 VSS.n158 VSS.n10 240.244
R272 VSS.n158 VSS.n13 240.244
R273 VSS.n206 VSS.n13 240.244
R274 VSS.n42 VSS.t1 222.373
R275 VSS.n146 VSS.t0 222.373
R276 VSS.n73 VSS.n71 163.367
R277 VSS.n77 VSS.n71 163.367
R278 VSS.n81 VSS.n79 163.367
R279 VSS.n85 VSS.n69 163.367
R280 VSS.n89 VSS.n87 163.367
R281 VSS.n93 VSS.n67 163.367
R282 VSS.n97 VSS.n95 163.367
R283 VSS.n199 VSS.n18 163.367
R284 VSS.n197 VSS.n196 163.367
R285 VSS.n194 VSS.n166 163.367
R286 VSS.n190 VSS.n189 163.367
R287 VSS.n187 VSS.n169 163.367
R288 VSS.n183 VSS.n182 163.367
R289 VSS.n180 VSS.n173 163.367
R290 VSS.n174 VSS.t4 111.651
R291 VSS.n63 VSS.t9 111.651
R292 VSS.n175 VSS.t5 77.7125
R293 VSS.n64 VSS.t8 77.7125
R294 VSS.t1 VSS.n35 74.1245
R295 VSS.t0 VSS.n145 74.1245
R296 VSS.n72 VSS.n60 71.676
R297 VSS.n78 VSS.n77 71.676
R298 VSS.n81 VSS.n80 71.676
R299 VSS.n86 VSS.n85 71.676
R300 VSS.n89 VSS.n88 71.676
R301 VSS.n94 VSS.n93 71.676
R302 VSS.n97 VSS.n96 71.676
R303 VSS.n198 VSS.n197 71.676
R304 VSS.n195 VSS.n194 71.676
R305 VSS.n190 VSS.n168 71.676
R306 VSS.n188 VSS.n187 71.676
R307 VSS.n183 VSS.n171 71.676
R308 VSS.n181 VSS.n180 71.676
R309 VSS.n172 VSS.n14 71.676
R310 VSS.n173 VSS.n172 71.676
R311 VSS.n182 VSS.n181 71.676
R312 VSS.n171 VSS.n169 71.676
R313 VSS.n189 VSS.n188 71.676
R314 VSS.n168 VSS.n166 71.676
R315 VSS.n196 VSS.n195 71.676
R316 VSS.n199 VSS.n198 71.676
R317 VSS.n73 VSS.n72 71.676
R318 VSS.n79 VSS.n78 71.676
R319 VSS.n80 VSS.n69 71.676
R320 VSS.n87 VSS.n86 71.676
R321 VSS.n88 VSS.n67 71.676
R322 VSS.n95 VSS.n94 71.676
R323 VSS.n96 VSS.n62 71.676
R324 VSS.n178 VSS.n175 34.5217
R325 VSS.n65 VSS.n64 34.5217
R326 VSS.n175 VSS.n174 33.9399
R327 VSS.n64 VSS.n63 33.9399
R328 VSS.n202 VSS.n201 31.5953
R329 VSS.n176 VSS.n12 31.5953
R330 VSS.n106 VSS.n59 31.5953
R331 VSS.n100 VSS.n99 31.5953
R332 VSS.n111 VSS.t7 20.7552
R333 VSS.n159 VSS.t3 20.7552
R334 VSS.n105 VSS.n58 19.3944
R335 VSS.n109 VSS.n58 19.3944
R336 VSS.n109 VSS.n48 19.3944
R337 VSS.n121 VSS.n48 19.3944
R338 VSS.n121 VSS.n45 19.3944
R339 VSS.n126 VSS.n45 19.3944
R340 VSS.n126 VSS.n46 19.3944
R341 VSS.n46 VSS.n33 19.3944
R342 VSS.n139 VSS.n33 19.3944
R343 VSS.n139 VSS.n31 19.3944
R344 VSS.n143 VSS.n31 19.3944
R345 VSS.n143 VSS.n27 19.3944
R346 VSS.n150 VSS.n27 19.3944
R347 VSS.n150 VSS.n25 19.3944
R348 VSS.n154 VSS.n25 19.3944
R349 VSS.n154 VSS.n21 19.3944
R350 VSS.n161 VSS.n21 19.3944
R351 VSS.n161 VSS.n19 19.3944
R352 VSS.n203 VSS.n19 19.3944
R353 VSS.n101 VSS.n54 19.3944
R354 VSS.n113 VSS.n54 19.3944
R355 VSS.n113 VSS.n52 19.3944
R356 VSS.n117 VSS.n52 19.3944
R357 VSS.n117 VSS.n39 19.3944
R358 VSS.n130 VSS.n39 19.3944
R359 VSS.n130 VSS.n37 19.3944
R360 VSS.n134 VSS.n37 19.3944
R361 VSS.n134 VSS.n2 19.3944
R362 VSS.n220 VSS.n2 19.3944
R363 VSS.n220 VSS.n219 19.3944
R364 VSS.n219 VSS.n218 19.3944
R365 VSS.n218 VSS.n6 19.3944
R366 VSS.n214 VSS.n6 19.3944
R367 VSS.n214 VSS.n213 19.3944
R368 VSS.n213 VSS.n212 19.3944
R369 VSS.n212 VSS.n11 19.3944
R370 VSS.n208 VSS.n11 19.3944
R371 VSS.n208 VSS.n207 19.3944
R372 VSS.n201 VSS.n200 10.6151
R373 VSS.n200 VSS.n164 10.6151
R374 VSS.n165 VSS.n164 10.6151
R375 VSS.n193 VSS.n165 10.6151
R376 VSS.n193 VSS.n192 10.6151
R377 VSS.n192 VSS.n191 10.6151
R378 VSS.n191 VSS.n167 10.6151
R379 VSS.n186 VSS.n167 10.6151
R380 VSS.n186 VSS.n185 10.6151
R381 VSS.n185 VSS.n184 10.6151
R382 VSS.n184 VSS.n170 10.6151
R383 VSS.n179 VSS.n170 10.6151
R384 VSS.n177 VSS.n176 10.6151
R385 VSS.n74 VSS.n59 10.6151
R386 VSS.n75 VSS.n74 10.6151
R387 VSS.n76 VSS.n75 10.6151
R388 VSS.n76 VSS.n70 10.6151
R389 VSS.n82 VSS.n70 10.6151
R390 VSS.n83 VSS.n82 10.6151
R391 VSS.n84 VSS.n83 10.6151
R392 VSS.n84 VSS.n68 10.6151
R393 VSS.n90 VSS.n68 10.6151
R394 VSS.n91 VSS.n90 10.6151
R395 VSS.n92 VSS.n91 10.6151
R396 VSS.n92 VSS.n66 10.6151
R397 VSS.n99 VSS.n98 10.6151
R398 VSS.n219 VSS.n0 9.3005
R399 VSS.n218 VSS.n217 9.3005
R400 VSS.n216 VSS.n6 9.3005
R401 VSS.n215 VSS.n214 9.3005
R402 VSS.n213 VSS.n7 9.3005
R403 VSS.n212 VSS.n211 9.3005
R404 VSS.n210 VSS.n11 9.3005
R405 VSS.n209 VSS.n208 9.3005
R406 VSS.n207 VSS.n12 9.3005
R407 VSS.n106 VSS.n105 9.3005
R408 VSS.n107 VSS.n58 9.3005
R409 VSS.n109 VSS.n108 9.3005
R410 VSS.n48 VSS.n47 9.3005
R411 VSS.n122 VSS.n121 9.3005
R412 VSS.n123 VSS.n45 9.3005
R413 VSS.n126 VSS.n125 9.3005
R414 VSS.n124 VSS.n46 9.3005
R415 VSS.n33 VSS.n32 9.3005
R416 VSS.n140 VSS.n139 9.3005
R417 VSS.n141 VSS.n31 9.3005
R418 VSS.n143 VSS.n142 9.3005
R419 VSS.n27 VSS.n26 9.3005
R420 VSS.n151 VSS.n150 9.3005
R421 VSS.n152 VSS.n25 9.3005
R422 VSS.n154 VSS.n153 9.3005
R423 VSS.n21 VSS.n20 9.3005
R424 VSS.n162 VSS.n161 9.3005
R425 VSS.n163 VSS.n19 9.3005
R426 VSS.n203 VSS.n202 9.3005
R427 VSS.n54 VSS.n53 9.3005
R428 VSS.n114 VSS.n113 9.3005
R429 VSS.n115 VSS.n52 9.3005
R430 VSS.n117 VSS.n116 9.3005
R431 VSS.n39 VSS.n38 9.3005
R432 VSS.n131 VSS.n130 9.3005
R433 VSS.n132 VSS.n37 9.3005
R434 VSS.n134 VSS.n133 9.3005
R435 VSS.n2 VSS.n1 9.3005
R436 VSS.n101 VSS.n100 9.3005
R437 VSS VSS.n220 9.3005
R438 VSS.n178 VSS.n177 8.74196
R439 VSS.n98 VSS.n65 8.74196
R440 VSS.n179 VSS.n178 1.87367
R441 VSS.n66 VSS.n65 1.87367
R442 VSS VSS.n0 0.152939
R443 VSS.n217 VSS.n0 0.152939
R444 VSS.n217 VSS.n216 0.152939
R445 VSS.n216 VSS.n215 0.152939
R446 VSS.n215 VSS.n7 0.152939
R447 VSS.n211 VSS.n7 0.152939
R448 VSS.n211 VSS.n210 0.152939
R449 VSS.n210 VSS.n209 0.152939
R450 VSS.n209 VSS.n12 0.152939
R451 VSS.n107 VSS.n106 0.152939
R452 VSS.n108 VSS.n107 0.152939
R453 VSS.n108 VSS.n47 0.152939
R454 VSS.n122 VSS.n47 0.152939
R455 VSS.n123 VSS.n122 0.152939
R456 VSS.n125 VSS.n123 0.152939
R457 VSS.n125 VSS.n124 0.152939
R458 VSS.n124 VSS.n32 0.152939
R459 VSS.n140 VSS.n32 0.152939
R460 VSS.n141 VSS.n140 0.152939
R461 VSS.n142 VSS.n141 0.152939
R462 VSS.n142 VSS.n26 0.152939
R463 VSS.n151 VSS.n26 0.152939
R464 VSS.n152 VSS.n151 0.152939
R465 VSS.n153 VSS.n152 0.152939
R466 VSS.n153 VSS.n20 0.152939
R467 VSS.n162 VSS.n20 0.152939
R468 VSS.n163 VSS.n162 0.152939
R469 VSS.n202 VSS.n163 0.152939
R470 VSS.n100 VSS.n53 0.152939
R471 VSS.n114 VSS.n53 0.152939
R472 VSS.n115 VSS.n114 0.152939
R473 VSS.n116 VSS.n115 0.152939
R474 VSS.n116 VSS.n38 0.152939
R475 VSS.n131 VSS.n38 0.152939
R476 VSS.n132 VSS.n131 0.152939
R477 VSS.n133 VSS.n132 0.152939
R478 VSS.n133 VSS.n1 0.152939
R479 VSS VSS.n1 0.1255
R480 VCC.n231 VCC.n14 408.293
R481 VCC.n229 VCC.n18 408.293
R482 VCC.n114 VCC.n57 408.293
R483 VCC.n112 VCC.n60 408.293
R484 VCC.n184 VCC.t4 280.805
R485 VCC.n61 VCC.t9 280.805
R486 VCC.n184 VCC.t2 280.149
R487 VCC.n61 VCC.t6 280.149
R488 VCC.n185 VCC.t5 245.315
R489 VCC.n62 VCC.t8 245.315
R490 VCC.n229 VCC.n228 185
R491 VCC.n230 VCC.n229 185
R492 VCC.n19 VCC.n17 185
R493 VCC.n17 VCC.n15 185
R494 VCC.n173 VCC.n172 185
R495 VCC.n172 VCC.n171 185
R496 VCC.n22 VCC.n21 185
R497 VCC.n169 VCC.n22 185
R498 VCC.n167 VCC.n166 185
R499 VCC.n168 VCC.n167 185
R500 VCC.n25 VCC.n24 185
R501 VCC.n24 VCC.n23 185
R502 VCC.n162 VCC.n161 185
R503 VCC.n161 VCC.n160 185
R504 VCC.n28 VCC.n27 185
R505 VCC.n158 VCC.n28 185
R506 VCC.n156 VCC.n155 185
R507 VCC.n157 VCC.n156 185
R508 VCC.n31 VCC.n30 185
R509 VCC.n30 VCC.n29 185
R510 VCC.n151 VCC.n150 185
R511 VCC.n150 VCC.n149 185
R512 VCC.n34 VCC.n33 185
R513 VCC.n35 VCC.n34 185
R514 VCC.n138 VCC.n137 185
R515 VCC.n139 VCC.n138 185
R516 VCC.n43 VCC.n42 185
R517 VCC.n140 VCC.n42 185
R518 VCC.n133 VCC.n132 185
R519 VCC.n132 VCC.n41 185
R520 VCC.n131 VCC.n45 185
R521 VCC.n131 VCC.n130 185
R522 VCC.n55 VCC.n46 185
R523 VCC.n47 VCC.n46 185
R524 VCC.n121 VCC.n120 185
R525 VCC.n122 VCC.n121 185
R526 VCC.n54 VCC.n53 185
R527 VCC.n59 VCC.n53 185
R528 VCC.n115 VCC.n114 185
R529 VCC.n114 VCC.n113 185
R530 VCC.n112 VCC.n111 185
R531 VCC.n113 VCC.n112 185
R532 VCC.n52 VCC.n51 185
R533 VCC.n59 VCC.n52 185
R534 VCC.n124 VCC.n123 185
R535 VCC.n123 VCC.n122 185
R536 VCC.n49 VCC.n48 185
R537 VCC.n48 VCC.n47 185
R538 VCC.n129 VCC.n128 185
R539 VCC.n130 VCC.n129 185
R540 VCC.n40 VCC.n39 185
R541 VCC.n41 VCC.n40 185
R542 VCC.n142 VCC.n141 185
R543 VCC.n141 VCC.n140 185
R544 VCC.n37 VCC.n36 185
R545 VCC.n139 VCC.n36 185
R546 VCC.n147 VCC.n146 185
R547 VCC.n147 VCC.n35 185
R548 VCC.n148 VCC.n2 185
R549 VCC.n149 VCC.n148 185
R550 VCC.n245 VCC.n3 185
R551 VCC.n29 VCC.n3 185
R552 VCC.n244 VCC.n4 185
R553 VCC.n157 VCC.n4 185
R554 VCC.n243 VCC.n5 185
R555 VCC.n158 VCC.n5 185
R556 VCC.n159 VCC.n6 185
R557 VCC.n160 VCC.n159 185
R558 VCC.n239 VCC.n8 185
R559 VCC.n23 VCC.n8 185
R560 VCC.n238 VCC.n9 185
R561 VCC.n168 VCC.n9 185
R562 VCC.n237 VCC.n10 185
R563 VCC.n169 VCC.n10 185
R564 VCC.n170 VCC.n11 185
R565 VCC.n171 VCC.n170 185
R566 VCC.n233 VCC.n13 185
R567 VCC.n15 VCC.n13 185
R568 VCC.n232 VCC.n231 185
R569 VCC.n231 VCC.n230 185
R570 VCC.n226 VCC.n18 185
R571 VCC.n225 VCC.n224 185
R572 VCC.n222 VCC.n176 185
R573 VCC.n220 VCC.n219 185
R574 VCC.n218 VCC.n177 185
R575 VCC.n217 VCC.n216 185
R576 VCC.n214 VCC.n178 185
R577 VCC.n212 VCC.n211 185
R578 VCC.n210 VCC.n179 185
R579 VCC.n209 VCC.n208 185
R580 VCC.n206 VCC.n180 185
R581 VCC.n204 VCC.n203 185
R582 VCC.n202 VCC.n181 185
R583 VCC.n201 VCC.n200 185
R584 VCC.n198 VCC.n182 185
R585 VCC.n196 VCC.n195 185
R586 VCC.n194 VCC.n183 185
R587 VCC.n193 VCC.n192 185
R588 VCC.n190 VCC.n189 185
R589 VCC.n188 VCC.n14 185
R590 VCC.n109 VCC.n60 185
R591 VCC.n108 VCC.n107 185
R592 VCC.n105 VCC.n104 185
R593 VCC.n105 VCC.n58 185
R594 VCC.n103 VCC.n64 185
R595 VCC.n102 VCC.n101 185
R596 VCC.n99 VCC.n65 185
R597 VCC.n97 VCC.n96 185
R598 VCC.n95 VCC.n66 185
R599 VCC.n94 VCC.n93 185
R600 VCC.n91 VCC.n67 185
R601 VCC.n89 VCC.n88 185
R602 VCC.n87 VCC.n68 185
R603 VCC.n86 VCC.n85 185
R604 VCC.n83 VCC.n69 185
R605 VCC.n81 VCC.n80 185
R606 VCC.n79 VCC.n70 185
R607 VCC.n78 VCC.n77 185
R608 VCC.n75 VCC.n71 185
R609 VCC.n73 VCC.n72 185
R610 VCC.n57 VCC.n56 185
R611 VCC.n58 VCC.n57 185
R612 VCC.n114 VCC.n53 146.341
R613 VCC.n121 VCC.n53 146.341
R614 VCC.n121 VCC.n46 146.341
R615 VCC.n131 VCC.n46 146.341
R616 VCC.n132 VCC.n131 146.341
R617 VCC.n132 VCC.n42 146.341
R618 VCC.n138 VCC.n42 146.341
R619 VCC.n138 VCC.n34 146.341
R620 VCC.n150 VCC.n34 146.341
R621 VCC.n150 VCC.n30 146.341
R622 VCC.n156 VCC.n30 146.341
R623 VCC.n156 VCC.n28 146.341
R624 VCC.n161 VCC.n28 146.341
R625 VCC.n161 VCC.n24 146.341
R626 VCC.n167 VCC.n24 146.341
R627 VCC.n167 VCC.n22 146.341
R628 VCC.n172 VCC.n22 146.341
R629 VCC.n172 VCC.n17 146.341
R630 VCC.n229 VCC.n17 146.341
R631 VCC.n112 VCC.n52 146.341
R632 VCC.n123 VCC.n52 146.341
R633 VCC.n123 VCC.n48 146.341
R634 VCC.n129 VCC.n48 146.341
R635 VCC.n129 VCC.n40 146.341
R636 VCC.n141 VCC.n40 146.341
R637 VCC.n141 VCC.n36 146.341
R638 VCC.n147 VCC.n36 146.341
R639 VCC.n148 VCC.n147 146.341
R640 VCC.n148 VCC.n3 146.341
R641 VCC.n4 VCC.n3 146.341
R642 VCC.n5 VCC.n4 146.341
R643 VCC.n159 VCC.n5 146.341
R644 VCC.n159 VCC.n8 146.341
R645 VCC.n9 VCC.n8 146.341
R646 VCC.n10 VCC.n9 146.341
R647 VCC.n170 VCC.n10 146.341
R648 VCC.n170 VCC.n13 146.341
R649 VCC.n231 VCC.n13 146.341
R650 VCC.n113 VCC.n58 104.653
R651 VCC.n230 VCC.n16 104.653
R652 VCC.n192 VCC.n190 99.5127
R653 VCC.n196 VCC.n183 99.5127
R654 VCC.n200 VCC.n198 99.5127
R655 VCC.n204 VCC.n181 99.5127
R656 VCC.n208 VCC.n206 99.5127
R657 VCC.n212 VCC.n179 99.5127
R658 VCC.n216 VCC.n214 99.5127
R659 VCC.n220 VCC.n177 99.5127
R660 VCC.n224 VCC.n222 99.5127
R661 VCC.n107 VCC.n105 99.5127
R662 VCC.n105 VCC.n64 99.5127
R663 VCC.n101 VCC.n99 99.5127
R664 VCC.n97 VCC.n66 99.5127
R665 VCC.n93 VCC.n91 99.5127
R666 VCC.n89 VCC.n68 99.5127
R667 VCC.n85 VCC.n83 99.5127
R668 VCC.n81 VCC.n70 99.5127
R669 VCC.n77 VCC.n75 99.5127
R670 VCC.n73 VCC.n57 99.5127
R671 VCC.n223 VCC.n16 72.8958
R672 VCC.n221 VCC.n16 72.8958
R673 VCC.n215 VCC.n16 72.8958
R674 VCC.n213 VCC.n16 72.8958
R675 VCC.n207 VCC.n16 72.8958
R676 VCC.n205 VCC.n16 72.8958
R677 VCC.n199 VCC.n16 72.8958
R678 VCC.n197 VCC.n16 72.8958
R679 VCC.n191 VCC.n16 72.8958
R680 VCC.n187 VCC.n16 72.8958
R681 VCC.n106 VCC.n58 72.8958
R682 VCC.n100 VCC.n58 72.8958
R683 VCC.n98 VCC.n58 72.8958
R684 VCC.n92 VCC.n58 72.8958
R685 VCC.n90 VCC.n58 72.8958
R686 VCC.n84 VCC.n58 72.8958
R687 VCC.n82 VCC.n58 72.8958
R688 VCC.n76 VCC.n58 72.8958
R689 VCC.n74 VCC.n58 72.8958
R690 VCC.n113 VCC.n59 54.2242
R691 VCC.n122 VCC.n47 54.2242
R692 VCC.n130 VCC.n47 54.2242
R693 VCC.n130 VCC.n41 54.2242
R694 VCC.n140 VCC.n41 54.2242
R695 VCC.n140 VCC.n139 54.2242
R696 VCC.n149 VCC.n35 54.2242
R697 VCC.n149 VCC.n29 54.2242
R698 VCC.n157 VCC.n29 54.2242
R699 VCC.n160 VCC.n158 54.2242
R700 VCC.n160 VCC.n23 54.2242
R701 VCC.n168 VCC.n23 54.2242
R702 VCC.n169 VCC.n168 54.2242
R703 VCC.n171 VCC.n169 54.2242
R704 VCC.n230 VCC.n15 54.2242
R705 VCC.n59 VCC.t7 45.0062
R706 VCC.t3 VCC.n15 45.0062
R707 VCC.n190 VCC.n187 39.2114
R708 VCC.n191 VCC.n183 39.2114
R709 VCC.n198 VCC.n197 39.2114
R710 VCC.n199 VCC.n181 39.2114
R711 VCC.n206 VCC.n205 39.2114
R712 VCC.n207 VCC.n179 39.2114
R713 VCC.n214 VCC.n213 39.2114
R714 VCC.n215 VCC.n177 39.2114
R715 VCC.n222 VCC.n221 39.2114
R716 VCC.n223 VCC.n18 39.2114
R717 VCC.n106 VCC.n60 39.2114
R718 VCC.n100 VCC.n64 39.2114
R719 VCC.n99 VCC.n98 39.2114
R720 VCC.n92 VCC.n66 39.2114
R721 VCC.n91 VCC.n90 39.2114
R722 VCC.n84 VCC.n68 39.2114
R723 VCC.n83 VCC.n82 39.2114
R724 VCC.n76 VCC.n70 39.2114
R725 VCC.n75 VCC.n74 39.2114
R726 VCC.n224 VCC.n223 39.2114
R727 VCC.n221 VCC.n220 39.2114
R728 VCC.n216 VCC.n215 39.2114
R729 VCC.n213 VCC.n212 39.2114
R730 VCC.n208 VCC.n207 39.2114
R731 VCC.n205 VCC.n204 39.2114
R732 VCC.n200 VCC.n199 39.2114
R733 VCC.n197 VCC.n196 39.2114
R734 VCC.n192 VCC.n191 39.2114
R735 VCC.n187 VCC.n14 39.2114
R736 VCC.n107 VCC.n106 39.2114
R737 VCC.n101 VCC.n100 39.2114
R738 VCC.n98 VCC.n97 39.2114
R739 VCC.n93 VCC.n92 39.2114
R740 VCC.n90 VCC.n89 39.2114
R741 VCC.n85 VCC.n84 39.2114
R742 VCC.n82 VCC.n81 39.2114
R743 VCC.n77 VCC.n76 39.2114
R744 VCC.n74 VCC.n73 39.2114
R745 VCC.n139 VCC.t1 36.3304
R746 VCC.n158 VCC.t0 36.3304
R747 VCC.n185 VCC.n184 35.4914
R748 VCC.n62 VCC.n61 35.4914
R749 VCC.n186 VCC.n185 29.4793
R750 VCC.n63 VCC.n62 29.4793
R751 VCC.n188 VCC.n12 29.4191
R752 VCC.n227 VCC.n226 29.4191
R753 VCC.n110 VCC.n109 29.4191
R754 VCC.n116 VCC.n56 29.4191
R755 VCC.n115 VCC.n54 19.3944
R756 VCC.n120 VCC.n54 19.3944
R757 VCC.n120 VCC.n55 19.3944
R758 VCC.n55 VCC.n45 19.3944
R759 VCC.n133 VCC.n45 19.3944
R760 VCC.n133 VCC.n43 19.3944
R761 VCC.n137 VCC.n43 19.3944
R762 VCC.n137 VCC.n33 19.3944
R763 VCC.n151 VCC.n33 19.3944
R764 VCC.n151 VCC.n31 19.3944
R765 VCC.n155 VCC.n31 19.3944
R766 VCC.n155 VCC.n27 19.3944
R767 VCC.n162 VCC.n27 19.3944
R768 VCC.n162 VCC.n25 19.3944
R769 VCC.n166 VCC.n25 19.3944
R770 VCC.n166 VCC.n21 19.3944
R771 VCC.n173 VCC.n21 19.3944
R772 VCC.n173 VCC.n19 19.3944
R773 VCC.n228 VCC.n19 19.3944
R774 VCC.n111 VCC.n51 19.3944
R775 VCC.n124 VCC.n51 19.3944
R776 VCC.n124 VCC.n49 19.3944
R777 VCC.n128 VCC.n49 19.3944
R778 VCC.n128 VCC.n39 19.3944
R779 VCC.n142 VCC.n39 19.3944
R780 VCC.n142 VCC.n37 19.3944
R781 VCC.n146 VCC.n37 19.3944
R782 VCC.n146 VCC.n2 19.3944
R783 VCC.n245 VCC.n2 19.3944
R784 VCC.n245 VCC.n244 19.3944
R785 VCC.n244 VCC.n243 19.3944
R786 VCC.n243 VCC.n6 19.3944
R787 VCC.n239 VCC.n6 19.3944
R788 VCC.n239 VCC.n238 19.3944
R789 VCC.n238 VCC.n237 19.3944
R790 VCC.n237 VCC.n11 19.3944
R791 VCC.n233 VCC.n11 19.3944
R792 VCC.n233 VCC.n232 19.3944
R793 VCC.t1 VCC.n35 17.8943
R794 VCC.t0 VCC.n157 17.8943
R795 VCC.n189 VCC.n188 10.6151
R796 VCC.n194 VCC.n193 10.6151
R797 VCC.n195 VCC.n194 10.6151
R798 VCC.n195 VCC.n182 10.6151
R799 VCC.n201 VCC.n182 10.6151
R800 VCC.n202 VCC.n201 10.6151
R801 VCC.n203 VCC.n202 10.6151
R802 VCC.n203 VCC.n180 10.6151
R803 VCC.n209 VCC.n180 10.6151
R804 VCC.n210 VCC.n209 10.6151
R805 VCC.n211 VCC.n210 10.6151
R806 VCC.n211 VCC.n178 10.6151
R807 VCC.n217 VCC.n178 10.6151
R808 VCC.n218 VCC.n217 10.6151
R809 VCC.n219 VCC.n218 10.6151
R810 VCC.n219 VCC.n176 10.6151
R811 VCC.n225 VCC.n176 10.6151
R812 VCC.n226 VCC.n225 10.6151
R813 VCC.n109 VCC.n108 10.6151
R814 VCC.n104 VCC.n103 10.6151
R815 VCC.n103 VCC.n102 10.6151
R816 VCC.n102 VCC.n65 10.6151
R817 VCC.n96 VCC.n65 10.6151
R818 VCC.n96 VCC.n95 10.6151
R819 VCC.n95 VCC.n94 10.6151
R820 VCC.n94 VCC.n67 10.6151
R821 VCC.n88 VCC.n67 10.6151
R822 VCC.n88 VCC.n87 10.6151
R823 VCC.n87 VCC.n86 10.6151
R824 VCC.n86 VCC.n69 10.6151
R825 VCC.n80 VCC.n69 10.6151
R826 VCC.n80 VCC.n79 10.6151
R827 VCC.n79 VCC.n78 10.6151
R828 VCC.n78 VCC.n71 10.6151
R829 VCC.n72 VCC.n71 10.6151
R830 VCC.n72 VCC.n56 10.6151
R831 VCC.n244 VCC.n0 9.3005
R832 VCC.n243 VCC.n242 9.3005
R833 VCC.n241 VCC.n6 9.3005
R834 VCC.n240 VCC.n239 9.3005
R835 VCC.n238 VCC.n7 9.3005
R836 VCC.n237 VCC.n236 9.3005
R837 VCC.n235 VCC.n11 9.3005
R838 VCC.n234 VCC.n233 9.3005
R839 VCC.n232 VCC.n12 9.3005
R840 VCC.n117 VCC.n54 9.3005
R841 VCC.n120 VCC.n119 9.3005
R842 VCC.n118 VCC.n55 9.3005
R843 VCC.n45 VCC.n44 9.3005
R844 VCC.n134 VCC.n133 9.3005
R845 VCC.n135 VCC.n43 9.3005
R846 VCC.n137 VCC.n136 9.3005
R847 VCC.n33 VCC.n32 9.3005
R848 VCC.n152 VCC.n151 9.3005
R849 VCC.n153 VCC.n31 9.3005
R850 VCC.n155 VCC.n154 9.3005
R851 VCC.n27 VCC.n26 9.3005
R852 VCC.n163 VCC.n162 9.3005
R853 VCC.n164 VCC.n25 9.3005
R854 VCC.n166 VCC.n165 9.3005
R855 VCC.n21 VCC.n20 9.3005
R856 VCC.n174 VCC.n173 9.3005
R857 VCC.n175 VCC.n19 9.3005
R858 VCC.n228 VCC.n227 9.3005
R859 VCC.n116 VCC.n115 9.3005
R860 VCC.n111 VCC.n110 9.3005
R861 VCC.n51 VCC.n50 9.3005
R862 VCC.n125 VCC.n124 9.3005
R863 VCC.n126 VCC.n49 9.3005
R864 VCC.n128 VCC.n127 9.3005
R865 VCC.n39 VCC.n38 9.3005
R866 VCC.n143 VCC.n142 9.3005
R867 VCC.n144 VCC.n37 9.3005
R868 VCC.n146 VCC.n145 9.3005
R869 VCC.n2 VCC.n1 9.3005
R870 VCC VCC.n245 9.3005
R871 VCC.n122 VCC.t7 9.21854
R872 VCC.n171 VCC.t3 9.21854
R873 VCC.n189 VCC.n186 6.86879
R874 VCC.n108 VCC.n63 6.86879
R875 VCC.n193 VCC.n186 3.74684
R876 VCC.n104 VCC.n63 3.74684
R877 VCC VCC.n0 0.152939
R878 VCC.n242 VCC.n0 0.152939
R879 VCC.n242 VCC.n241 0.152939
R880 VCC.n241 VCC.n240 0.152939
R881 VCC.n240 VCC.n7 0.152939
R882 VCC.n236 VCC.n7 0.152939
R883 VCC.n236 VCC.n235 0.152939
R884 VCC.n235 VCC.n234 0.152939
R885 VCC.n234 VCC.n12 0.152939
R886 VCC.n117 VCC.n116 0.152939
R887 VCC.n119 VCC.n117 0.152939
R888 VCC.n119 VCC.n118 0.152939
R889 VCC.n118 VCC.n44 0.152939
R890 VCC.n134 VCC.n44 0.152939
R891 VCC.n135 VCC.n134 0.152939
R892 VCC.n136 VCC.n135 0.152939
R893 VCC.n136 VCC.n32 0.152939
R894 VCC.n152 VCC.n32 0.152939
R895 VCC.n153 VCC.n152 0.152939
R896 VCC.n154 VCC.n153 0.152939
R897 VCC.n154 VCC.n26 0.152939
R898 VCC.n163 VCC.n26 0.152939
R899 VCC.n164 VCC.n163 0.152939
R900 VCC.n165 VCC.n164 0.152939
R901 VCC.n165 VCC.n20 0.152939
R902 VCC.n174 VCC.n20 0.152939
R903 VCC.n175 VCC.n174 0.152939
R904 VCC.n227 VCC.n175 0.152939
R905 VCC.n110 VCC.n50 0.152939
R906 VCC.n125 VCC.n50 0.152939
R907 VCC.n126 VCC.n125 0.152939
R908 VCC.n127 VCC.n126 0.152939
R909 VCC.n127 VCC.n38 0.152939
R910 VCC.n143 VCC.n38 0.152939
R911 VCC.n144 VCC.n143 0.152939
R912 VCC.n145 VCC.n144 0.152939
R913 VCC.n145 VCC.n1 0.152939
R914 VCC VCC.n1 0.1255
R915 VGP.n0 VGP.t0 111.07
R916 VGP.n0 VGP.t1 110.754
R917 VGP VGP.n0 13.1193
C0 VGP VCC 1.39871f
C1 VIN VGP 0.835111f
C2 VOUT VGP 0.689629f
C3 VGN VCC 0.010333f
C4 VGN VIN 0.572556f
C5 VGN VOUT 0.433793f
C6 VIN VCC 1.10996f
C7 VOUT VCC 0.71403f
C8 VOUT VIN 1.70878f
C9 VGN VGP 0.011363f
C10 VGN VSS 1.65915f
C11 VOUT VSS 0.766005f
C12 VIN VSS 1.15936f
C13 VGP VSS 0.405925f
C14 VCC VSS 14.7558f
.ends

