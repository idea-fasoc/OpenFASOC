* NGSPICE file created from diff_pair_sample_1369.ext - technology: sky130A

.subckt diff_pair_sample_1369 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t9 VN.t0 VTAIL.t17 B.t2 sky130_fd_pr__nfet_01v8 ad=3.2307 pd=19.91 as=7.6362 ps=39.94 w=19.58 l=3.23
X1 VDD2.t8 VN.t1 VTAIL.t11 B.t1 sky130_fd_pr__nfet_01v8 ad=3.2307 pd=19.91 as=3.2307 ps=19.91 w=19.58 l=3.23
X2 VDD2.t7 VN.t2 VTAIL.t12 B.t7 sky130_fd_pr__nfet_01v8 ad=7.6362 pd=39.94 as=3.2307 ps=19.91 w=19.58 l=3.23
X3 VDD1.t9 VP.t0 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=3.2307 pd=19.91 as=7.6362 ps=39.94 w=19.58 l=3.23
X4 B.t23 B.t21 B.t22 B.t11 sky130_fd_pr__nfet_01v8 ad=7.6362 pd=39.94 as=0 ps=0 w=19.58 l=3.23
X5 B.t20 B.t18 B.t19 B.t15 sky130_fd_pr__nfet_01v8 ad=7.6362 pd=39.94 as=0 ps=0 w=19.58 l=3.23
X6 VTAIL.t0 VP.t1 VDD1.t8 B.t0 sky130_fd_pr__nfet_01v8 ad=3.2307 pd=19.91 as=3.2307 ps=19.91 w=19.58 l=3.23
X7 VDD1.t7 VP.t2 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=3.2307 pd=19.91 as=7.6362 ps=39.94 w=19.58 l=3.23
X8 VDD2.t6 VN.t3 VTAIL.t18 B.t4 sky130_fd_pr__nfet_01v8 ad=7.6362 pd=39.94 as=3.2307 ps=19.91 w=19.58 l=3.23
X9 VTAIL.t10 VN.t4 VDD2.t5 B.t0 sky130_fd_pr__nfet_01v8 ad=3.2307 pd=19.91 as=3.2307 ps=19.91 w=19.58 l=3.23
X10 VTAIL.t14 VN.t5 VDD2.t4 B.t9 sky130_fd_pr__nfet_01v8 ad=3.2307 pd=19.91 as=3.2307 ps=19.91 w=19.58 l=3.23
X11 VTAIL.t19 VN.t6 VDD2.t3 B.t6 sky130_fd_pr__nfet_01v8 ad=3.2307 pd=19.91 as=3.2307 ps=19.91 w=19.58 l=3.23
X12 VDD2.t2 VN.t7 VTAIL.t13 B.t3 sky130_fd_pr__nfet_01v8 ad=3.2307 pd=19.91 as=7.6362 ps=39.94 w=19.58 l=3.23
X13 VTAIL.t15 VN.t8 VDD2.t1 B.t5 sky130_fd_pr__nfet_01v8 ad=3.2307 pd=19.91 as=3.2307 ps=19.91 w=19.58 l=3.23
X14 VTAIL.t5 VP.t3 VDD1.t6 B.t5 sky130_fd_pr__nfet_01v8 ad=3.2307 pd=19.91 as=3.2307 ps=19.91 w=19.58 l=3.23
X15 VTAIL.t9 VP.t4 VDD1.t5 B.t9 sky130_fd_pr__nfet_01v8 ad=3.2307 pd=19.91 as=3.2307 ps=19.91 w=19.58 l=3.23
X16 VDD1.t4 VP.t5 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=3.2307 pd=19.91 as=3.2307 ps=19.91 w=19.58 l=3.23
X17 VDD1.t3 VP.t6 VTAIL.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=7.6362 pd=39.94 as=3.2307 ps=19.91 w=19.58 l=3.23
X18 VTAIL.t6 VP.t7 VDD1.t2 B.t6 sky130_fd_pr__nfet_01v8 ad=3.2307 pd=19.91 as=3.2307 ps=19.91 w=19.58 l=3.23
X19 B.t17 B.t14 B.t16 B.t15 sky130_fd_pr__nfet_01v8 ad=7.6362 pd=39.94 as=0 ps=0 w=19.58 l=3.23
X20 VDD2.t0 VN.t9 VTAIL.t16 B.t8 sky130_fd_pr__nfet_01v8 ad=3.2307 pd=19.91 as=3.2307 ps=19.91 w=19.58 l=3.23
X21 VDD1.t1 VP.t8 VTAIL.t7 B.t7 sky130_fd_pr__nfet_01v8 ad=7.6362 pd=39.94 as=3.2307 ps=19.91 w=19.58 l=3.23
X22 B.t13 B.t10 B.t12 B.t11 sky130_fd_pr__nfet_01v8 ad=7.6362 pd=39.94 as=0 ps=0 w=19.58 l=3.23
X23 VDD1.t0 VP.t9 VTAIL.t8 B.t8 sky130_fd_pr__nfet_01v8 ad=3.2307 pd=19.91 as=3.2307 ps=19.91 w=19.58 l=3.23
R0 VN.n61 VN.t7 179.448
R1 VN.n13 VN.t2 179.448
R2 VN.n94 VN.n93 161.3
R3 VN.n92 VN.n49 161.3
R4 VN.n91 VN.n90 161.3
R5 VN.n89 VN.n50 161.3
R6 VN.n88 VN.n87 161.3
R7 VN.n86 VN.n51 161.3
R8 VN.n85 VN.n84 161.3
R9 VN.n83 VN.n82 161.3
R10 VN.n81 VN.n53 161.3
R11 VN.n80 VN.n79 161.3
R12 VN.n78 VN.n54 161.3
R13 VN.n77 VN.n76 161.3
R14 VN.n75 VN.n55 161.3
R15 VN.n74 VN.n73 161.3
R16 VN.n72 VN.n71 161.3
R17 VN.n70 VN.n57 161.3
R18 VN.n69 VN.n68 161.3
R19 VN.n67 VN.n58 161.3
R20 VN.n66 VN.n65 161.3
R21 VN.n64 VN.n59 161.3
R22 VN.n63 VN.n62 161.3
R23 VN.n46 VN.n45 161.3
R24 VN.n44 VN.n1 161.3
R25 VN.n43 VN.n42 161.3
R26 VN.n41 VN.n2 161.3
R27 VN.n40 VN.n39 161.3
R28 VN.n38 VN.n3 161.3
R29 VN.n37 VN.n36 161.3
R30 VN.n35 VN.n34 161.3
R31 VN.n33 VN.n5 161.3
R32 VN.n32 VN.n31 161.3
R33 VN.n30 VN.n6 161.3
R34 VN.n29 VN.n28 161.3
R35 VN.n27 VN.n7 161.3
R36 VN.n26 VN.n25 161.3
R37 VN.n24 VN.n23 161.3
R38 VN.n22 VN.n9 161.3
R39 VN.n21 VN.n20 161.3
R40 VN.n19 VN.n10 161.3
R41 VN.n18 VN.n17 161.3
R42 VN.n16 VN.n11 161.3
R43 VN.n15 VN.n14 161.3
R44 VN.n12 VN.t6 146.093
R45 VN.n8 VN.t1 146.093
R46 VN.n4 VN.t5 146.093
R47 VN.n0 VN.t0 146.093
R48 VN.n60 VN.t8 146.093
R49 VN.n56 VN.t9 146.093
R50 VN.n52 VN.t4 146.093
R51 VN.n48 VN.t3 146.093
R52 VN.n47 VN.n0 72.0476
R53 VN.n95 VN.n48 72.0476
R54 VN VN.n95 62.5966
R55 VN.n13 VN.n12 59.1354
R56 VN.n61 VN.n60 59.1354
R57 VN.n43 VN.n2 49.296
R58 VN.n91 VN.n50 49.296
R59 VN.n17 VN.n10 43.4833
R60 VN.n32 VN.n6 43.4833
R61 VN.n65 VN.n58 43.4833
R62 VN.n80 VN.n54 43.4833
R63 VN.n21 VN.n10 37.6707
R64 VN.n28 VN.n6 37.6707
R65 VN.n69 VN.n58 37.6707
R66 VN.n76 VN.n54 37.6707
R67 VN.n39 VN.n2 31.8581
R68 VN.n87 VN.n50 31.8581
R69 VN.n16 VN.n15 24.5923
R70 VN.n17 VN.n16 24.5923
R71 VN.n22 VN.n21 24.5923
R72 VN.n23 VN.n22 24.5923
R73 VN.n27 VN.n26 24.5923
R74 VN.n28 VN.n27 24.5923
R75 VN.n33 VN.n32 24.5923
R76 VN.n34 VN.n33 24.5923
R77 VN.n38 VN.n37 24.5923
R78 VN.n39 VN.n38 24.5923
R79 VN.n44 VN.n43 24.5923
R80 VN.n45 VN.n44 24.5923
R81 VN.n65 VN.n64 24.5923
R82 VN.n64 VN.n63 24.5923
R83 VN.n76 VN.n75 24.5923
R84 VN.n75 VN.n74 24.5923
R85 VN.n71 VN.n70 24.5923
R86 VN.n70 VN.n69 24.5923
R87 VN.n87 VN.n86 24.5923
R88 VN.n86 VN.n85 24.5923
R89 VN.n82 VN.n81 24.5923
R90 VN.n81 VN.n80 24.5923
R91 VN.n93 VN.n92 24.5923
R92 VN.n92 VN.n91 24.5923
R93 VN.n45 VN.n0 18.1985
R94 VN.n93 VN.n48 18.1985
R95 VN.n15 VN.n12 15.2474
R96 VN.n34 VN.n4 15.2474
R97 VN.n63 VN.n60 15.2474
R98 VN.n82 VN.n52 15.2474
R99 VN.n23 VN.n8 12.2964
R100 VN.n26 VN.n8 12.2964
R101 VN.n74 VN.n56 12.2964
R102 VN.n71 VN.n56 12.2964
R103 VN.n37 VN.n4 9.3454
R104 VN.n85 VN.n52 9.3454
R105 VN.n62 VN.n61 3.98083
R106 VN.n14 VN.n13 3.98083
R107 VN.n95 VN.n94 0.354861
R108 VN.n47 VN.n46 0.354861
R109 VN VN.n47 0.267071
R110 VN.n94 VN.n49 0.189894
R111 VN.n90 VN.n49 0.189894
R112 VN.n90 VN.n89 0.189894
R113 VN.n89 VN.n88 0.189894
R114 VN.n88 VN.n51 0.189894
R115 VN.n84 VN.n51 0.189894
R116 VN.n84 VN.n83 0.189894
R117 VN.n83 VN.n53 0.189894
R118 VN.n79 VN.n53 0.189894
R119 VN.n79 VN.n78 0.189894
R120 VN.n78 VN.n77 0.189894
R121 VN.n77 VN.n55 0.189894
R122 VN.n73 VN.n55 0.189894
R123 VN.n73 VN.n72 0.189894
R124 VN.n72 VN.n57 0.189894
R125 VN.n68 VN.n57 0.189894
R126 VN.n68 VN.n67 0.189894
R127 VN.n67 VN.n66 0.189894
R128 VN.n66 VN.n59 0.189894
R129 VN.n62 VN.n59 0.189894
R130 VN.n14 VN.n11 0.189894
R131 VN.n18 VN.n11 0.189894
R132 VN.n19 VN.n18 0.189894
R133 VN.n20 VN.n19 0.189894
R134 VN.n20 VN.n9 0.189894
R135 VN.n24 VN.n9 0.189894
R136 VN.n25 VN.n24 0.189894
R137 VN.n25 VN.n7 0.189894
R138 VN.n29 VN.n7 0.189894
R139 VN.n30 VN.n29 0.189894
R140 VN.n31 VN.n30 0.189894
R141 VN.n31 VN.n5 0.189894
R142 VN.n35 VN.n5 0.189894
R143 VN.n36 VN.n35 0.189894
R144 VN.n36 VN.n3 0.189894
R145 VN.n40 VN.n3 0.189894
R146 VN.n41 VN.n40 0.189894
R147 VN.n42 VN.n41 0.189894
R148 VN.n42 VN.n1 0.189894
R149 VN.n46 VN.n1 0.189894
R150 VTAIL.n448 VTAIL.n344 289.615
R151 VTAIL.n106 VTAIL.n2 289.615
R152 VTAIL.n338 VTAIL.n234 289.615
R153 VTAIL.n224 VTAIL.n120 289.615
R154 VTAIL.n381 VTAIL.n380 185
R155 VTAIL.n383 VTAIL.n382 185
R156 VTAIL.n376 VTAIL.n375 185
R157 VTAIL.n389 VTAIL.n388 185
R158 VTAIL.n391 VTAIL.n390 185
R159 VTAIL.n372 VTAIL.n371 185
R160 VTAIL.n397 VTAIL.n396 185
R161 VTAIL.n399 VTAIL.n398 185
R162 VTAIL.n368 VTAIL.n367 185
R163 VTAIL.n405 VTAIL.n404 185
R164 VTAIL.n407 VTAIL.n406 185
R165 VTAIL.n364 VTAIL.n363 185
R166 VTAIL.n413 VTAIL.n412 185
R167 VTAIL.n415 VTAIL.n414 185
R168 VTAIL.n360 VTAIL.n359 185
R169 VTAIL.n422 VTAIL.n421 185
R170 VTAIL.n423 VTAIL.n358 185
R171 VTAIL.n425 VTAIL.n424 185
R172 VTAIL.n356 VTAIL.n355 185
R173 VTAIL.n431 VTAIL.n430 185
R174 VTAIL.n433 VTAIL.n432 185
R175 VTAIL.n352 VTAIL.n351 185
R176 VTAIL.n439 VTAIL.n438 185
R177 VTAIL.n441 VTAIL.n440 185
R178 VTAIL.n348 VTAIL.n347 185
R179 VTAIL.n447 VTAIL.n446 185
R180 VTAIL.n449 VTAIL.n448 185
R181 VTAIL.n39 VTAIL.n38 185
R182 VTAIL.n41 VTAIL.n40 185
R183 VTAIL.n34 VTAIL.n33 185
R184 VTAIL.n47 VTAIL.n46 185
R185 VTAIL.n49 VTAIL.n48 185
R186 VTAIL.n30 VTAIL.n29 185
R187 VTAIL.n55 VTAIL.n54 185
R188 VTAIL.n57 VTAIL.n56 185
R189 VTAIL.n26 VTAIL.n25 185
R190 VTAIL.n63 VTAIL.n62 185
R191 VTAIL.n65 VTAIL.n64 185
R192 VTAIL.n22 VTAIL.n21 185
R193 VTAIL.n71 VTAIL.n70 185
R194 VTAIL.n73 VTAIL.n72 185
R195 VTAIL.n18 VTAIL.n17 185
R196 VTAIL.n80 VTAIL.n79 185
R197 VTAIL.n81 VTAIL.n16 185
R198 VTAIL.n83 VTAIL.n82 185
R199 VTAIL.n14 VTAIL.n13 185
R200 VTAIL.n89 VTAIL.n88 185
R201 VTAIL.n91 VTAIL.n90 185
R202 VTAIL.n10 VTAIL.n9 185
R203 VTAIL.n97 VTAIL.n96 185
R204 VTAIL.n99 VTAIL.n98 185
R205 VTAIL.n6 VTAIL.n5 185
R206 VTAIL.n105 VTAIL.n104 185
R207 VTAIL.n107 VTAIL.n106 185
R208 VTAIL.n339 VTAIL.n338 185
R209 VTAIL.n337 VTAIL.n336 185
R210 VTAIL.n238 VTAIL.n237 185
R211 VTAIL.n331 VTAIL.n330 185
R212 VTAIL.n329 VTAIL.n328 185
R213 VTAIL.n242 VTAIL.n241 185
R214 VTAIL.n323 VTAIL.n322 185
R215 VTAIL.n321 VTAIL.n320 185
R216 VTAIL.n246 VTAIL.n245 185
R217 VTAIL.n250 VTAIL.n248 185
R218 VTAIL.n315 VTAIL.n314 185
R219 VTAIL.n313 VTAIL.n312 185
R220 VTAIL.n252 VTAIL.n251 185
R221 VTAIL.n307 VTAIL.n306 185
R222 VTAIL.n305 VTAIL.n304 185
R223 VTAIL.n256 VTAIL.n255 185
R224 VTAIL.n299 VTAIL.n298 185
R225 VTAIL.n297 VTAIL.n296 185
R226 VTAIL.n260 VTAIL.n259 185
R227 VTAIL.n291 VTAIL.n290 185
R228 VTAIL.n289 VTAIL.n288 185
R229 VTAIL.n264 VTAIL.n263 185
R230 VTAIL.n283 VTAIL.n282 185
R231 VTAIL.n281 VTAIL.n280 185
R232 VTAIL.n268 VTAIL.n267 185
R233 VTAIL.n275 VTAIL.n274 185
R234 VTAIL.n273 VTAIL.n272 185
R235 VTAIL.n225 VTAIL.n224 185
R236 VTAIL.n223 VTAIL.n222 185
R237 VTAIL.n124 VTAIL.n123 185
R238 VTAIL.n217 VTAIL.n216 185
R239 VTAIL.n215 VTAIL.n214 185
R240 VTAIL.n128 VTAIL.n127 185
R241 VTAIL.n209 VTAIL.n208 185
R242 VTAIL.n207 VTAIL.n206 185
R243 VTAIL.n132 VTAIL.n131 185
R244 VTAIL.n136 VTAIL.n134 185
R245 VTAIL.n201 VTAIL.n200 185
R246 VTAIL.n199 VTAIL.n198 185
R247 VTAIL.n138 VTAIL.n137 185
R248 VTAIL.n193 VTAIL.n192 185
R249 VTAIL.n191 VTAIL.n190 185
R250 VTAIL.n142 VTAIL.n141 185
R251 VTAIL.n185 VTAIL.n184 185
R252 VTAIL.n183 VTAIL.n182 185
R253 VTAIL.n146 VTAIL.n145 185
R254 VTAIL.n177 VTAIL.n176 185
R255 VTAIL.n175 VTAIL.n174 185
R256 VTAIL.n150 VTAIL.n149 185
R257 VTAIL.n169 VTAIL.n168 185
R258 VTAIL.n167 VTAIL.n166 185
R259 VTAIL.n154 VTAIL.n153 185
R260 VTAIL.n161 VTAIL.n160 185
R261 VTAIL.n159 VTAIL.n158 185
R262 VTAIL.n379 VTAIL.t17 147.659
R263 VTAIL.n37 VTAIL.t3 147.659
R264 VTAIL.n271 VTAIL.t2 147.659
R265 VTAIL.n157 VTAIL.t13 147.659
R266 VTAIL.n382 VTAIL.n381 104.615
R267 VTAIL.n382 VTAIL.n375 104.615
R268 VTAIL.n389 VTAIL.n375 104.615
R269 VTAIL.n390 VTAIL.n389 104.615
R270 VTAIL.n390 VTAIL.n371 104.615
R271 VTAIL.n397 VTAIL.n371 104.615
R272 VTAIL.n398 VTAIL.n397 104.615
R273 VTAIL.n398 VTAIL.n367 104.615
R274 VTAIL.n405 VTAIL.n367 104.615
R275 VTAIL.n406 VTAIL.n405 104.615
R276 VTAIL.n406 VTAIL.n363 104.615
R277 VTAIL.n413 VTAIL.n363 104.615
R278 VTAIL.n414 VTAIL.n413 104.615
R279 VTAIL.n414 VTAIL.n359 104.615
R280 VTAIL.n422 VTAIL.n359 104.615
R281 VTAIL.n423 VTAIL.n422 104.615
R282 VTAIL.n424 VTAIL.n423 104.615
R283 VTAIL.n424 VTAIL.n355 104.615
R284 VTAIL.n431 VTAIL.n355 104.615
R285 VTAIL.n432 VTAIL.n431 104.615
R286 VTAIL.n432 VTAIL.n351 104.615
R287 VTAIL.n439 VTAIL.n351 104.615
R288 VTAIL.n440 VTAIL.n439 104.615
R289 VTAIL.n440 VTAIL.n347 104.615
R290 VTAIL.n447 VTAIL.n347 104.615
R291 VTAIL.n448 VTAIL.n447 104.615
R292 VTAIL.n40 VTAIL.n39 104.615
R293 VTAIL.n40 VTAIL.n33 104.615
R294 VTAIL.n47 VTAIL.n33 104.615
R295 VTAIL.n48 VTAIL.n47 104.615
R296 VTAIL.n48 VTAIL.n29 104.615
R297 VTAIL.n55 VTAIL.n29 104.615
R298 VTAIL.n56 VTAIL.n55 104.615
R299 VTAIL.n56 VTAIL.n25 104.615
R300 VTAIL.n63 VTAIL.n25 104.615
R301 VTAIL.n64 VTAIL.n63 104.615
R302 VTAIL.n64 VTAIL.n21 104.615
R303 VTAIL.n71 VTAIL.n21 104.615
R304 VTAIL.n72 VTAIL.n71 104.615
R305 VTAIL.n72 VTAIL.n17 104.615
R306 VTAIL.n80 VTAIL.n17 104.615
R307 VTAIL.n81 VTAIL.n80 104.615
R308 VTAIL.n82 VTAIL.n81 104.615
R309 VTAIL.n82 VTAIL.n13 104.615
R310 VTAIL.n89 VTAIL.n13 104.615
R311 VTAIL.n90 VTAIL.n89 104.615
R312 VTAIL.n90 VTAIL.n9 104.615
R313 VTAIL.n97 VTAIL.n9 104.615
R314 VTAIL.n98 VTAIL.n97 104.615
R315 VTAIL.n98 VTAIL.n5 104.615
R316 VTAIL.n105 VTAIL.n5 104.615
R317 VTAIL.n106 VTAIL.n105 104.615
R318 VTAIL.n338 VTAIL.n337 104.615
R319 VTAIL.n337 VTAIL.n237 104.615
R320 VTAIL.n330 VTAIL.n237 104.615
R321 VTAIL.n330 VTAIL.n329 104.615
R322 VTAIL.n329 VTAIL.n241 104.615
R323 VTAIL.n322 VTAIL.n241 104.615
R324 VTAIL.n322 VTAIL.n321 104.615
R325 VTAIL.n321 VTAIL.n245 104.615
R326 VTAIL.n250 VTAIL.n245 104.615
R327 VTAIL.n314 VTAIL.n250 104.615
R328 VTAIL.n314 VTAIL.n313 104.615
R329 VTAIL.n313 VTAIL.n251 104.615
R330 VTAIL.n306 VTAIL.n251 104.615
R331 VTAIL.n306 VTAIL.n305 104.615
R332 VTAIL.n305 VTAIL.n255 104.615
R333 VTAIL.n298 VTAIL.n255 104.615
R334 VTAIL.n298 VTAIL.n297 104.615
R335 VTAIL.n297 VTAIL.n259 104.615
R336 VTAIL.n290 VTAIL.n259 104.615
R337 VTAIL.n290 VTAIL.n289 104.615
R338 VTAIL.n289 VTAIL.n263 104.615
R339 VTAIL.n282 VTAIL.n263 104.615
R340 VTAIL.n282 VTAIL.n281 104.615
R341 VTAIL.n281 VTAIL.n267 104.615
R342 VTAIL.n274 VTAIL.n267 104.615
R343 VTAIL.n274 VTAIL.n273 104.615
R344 VTAIL.n224 VTAIL.n223 104.615
R345 VTAIL.n223 VTAIL.n123 104.615
R346 VTAIL.n216 VTAIL.n123 104.615
R347 VTAIL.n216 VTAIL.n215 104.615
R348 VTAIL.n215 VTAIL.n127 104.615
R349 VTAIL.n208 VTAIL.n127 104.615
R350 VTAIL.n208 VTAIL.n207 104.615
R351 VTAIL.n207 VTAIL.n131 104.615
R352 VTAIL.n136 VTAIL.n131 104.615
R353 VTAIL.n200 VTAIL.n136 104.615
R354 VTAIL.n200 VTAIL.n199 104.615
R355 VTAIL.n199 VTAIL.n137 104.615
R356 VTAIL.n192 VTAIL.n137 104.615
R357 VTAIL.n192 VTAIL.n191 104.615
R358 VTAIL.n191 VTAIL.n141 104.615
R359 VTAIL.n184 VTAIL.n141 104.615
R360 VTAIL.n184 VTAIL.n183 104.615
R361 VTAIL.n183 VTAIL.n145 104.615
R362 VTAIL.n176 VTAIL.n145 104.615
R363 VTAIL.n176 VTAIL.n175 104.615
R364 VTAIL.n175 VTAIL.n149 104.615
R365 VTAIL.n168 VTAIL.n149 104.615
R366 VTAIL.n168 VTAIL.n167 104.615
R367 VTAIL.n167 VTAIL.n153 104.615
R368 VTAIL.n160 VTAIL.n153 104.615
R369 VTAIL.n160 VTAIL.n159 104.615
R370 VTAIL.n381 VTAIL.t17 52.3082
R371 VTAIL.n39 VTAIL.t3 52.3082
R372 VTAIL.n273 VTAIL.t2 52.3082
R373 VTAIL.n159 VTAIL.t13 52.3082
R374 VTAIL.n233 VTAIL.n232 41.984
R375 VTAIL.n231 VTAIL.n230 41.984
R376 VTAIL.n119 VTAIL.n118 41.984
R377 VTAIL.n117 VTAIL.n116 41.984
R378 VTAIL.n455 VTAIL.n454 41.9838
R379 VTAIL.n1 VTAIL.n0 41.9838
R380 VTAIL.n113 VTAIL.n112 41.9838
R381 VTAIL.n115 VTAIL.n114 41.9838
R382 VTAIL.n117 VTAIL.n115 35.3841
R383 VTAIL.n453 VTAIL.n343 32.3152
R384 VTAIL.n453 VTAIL.n452 30.246
R385 VTAIL.n111 VTAIL.n110 30.246
R386 VTAIL.n343 VTAIL.n342 30.246
R387 VTAIL.n229 VTAIL.n228 30.246
R388 VTAIL.n380 VTAIL.n379 15.6677
R389 VTAIL.n38 VTAIL.n37 15.6677
R390 VTAIL.n272 VTAIL.n271 15.6677
R391 VTAIL.n158 VTAIL.n157 15.6677
R392 VTAIL.n425 VTAIL.n356 13.1884
R393 VTAIL.n83 VTAIL.n14 13.1884
R394 VTAIL.n248 VTAIL.n246 13.1884
R395 VTAIL.n134 VTAIL.n132 13.1884
R396 VTAIL.n383 VTAIL.n378 12.8005
R397 VTAIL.n426 VTAIL.n358 12.8005
R398 VTAIL.n430 VTAIL.n429 12.8005
R399 VTAIL.n41 VTAIL.n36 12.8005
R400 VTAIL.n84 VTAIL.n16 12.8005
R401 VTAIL.n88 VTAIL.n87 12.8005
R402 VTAIL.n320 VTAIL.n319 12.8005
R403 VTAIL.n316 VTAIL.n315 12.8005
R404 VTAIL.n275 VTAIL.n270 12.8005
R405 VTAIL.n206 VTAIL.n205 12.8005
R406 VTAIL.n202 VTAIL.n201 12.8005
R407 VTAIL.n161 VTAIL.n156 12.8005
R408 VTAIL.n384 VTAIL.n376 12.0247
R409 VTAIL.n421 VTAIL.n420 12.0247
R410 VTAIL.n433 VTAIL.n354 12.0247
R411 VTAIL.n42 VTAIL.n34 12.0247
R412 VTAIL.n79 VTAIL.n78 12.0247
R413 VTAIL.n91 VTAIL.n12 12.0247
R414 VTAIL.n323 VTAIL.n244 12.0247
R415 VTAIL.n312 VTAIL.n249 12.0247
R416 VTAIL.n276 VTAIL.n268 12.0247
R417 VTAIL.n209 VTAIL.n130 12.0247
R418 VTAIL.n198 VTAIL.n135 12.0247
R419 VTAIL.n162 VTAIL.n154 12.0247
R420 VTAIL.n388 VTAIL.n387 11.249
R421 VTAIL.n419 VTAIL.n360 11.249
R422 VTAIL.n434 VTAIL.n352 11.249
R423 VTAIL.n46 VTAIL.n45 11.249
R424 VTAIL.n77 VTAIL.n18 11.249
R425 VTAIL.n92 VTAIL.n10 11.249
R426 VTAIL.n324 VTAIL.n242 11.249
R427 VTAIL.n311 VTAIL.n252 11.249
R428 VTAIL.n280 VTAIL.n279 11.249
R429 VTAIL.n210 VTAIL.n128 11.249
R430 VTAIL.n197 VTAIL.n138 11.249
R431 VTAIL.n166 VTAIL.n165 11.249
R432 VTAIL.n391 VTAIL.n374 10.4732
R433 VTAIL.n416 VTAIL.n415 10.4732
R434 VTAIL.n438 VTAIL.n437 10.4732
R435 VTAIL.n49 VTAIL.n32 10.4732
R436 VTAIL.n74 VTAIL.n73 10.4732
R437 VTAIL.n96 VTAIL.n95 10.4732
R438 VTAIL.n328 VTAIL.n327 10.4732
R439 VTAIL.n308 VTAIL.n307 10.4732
R440 VTAIL.n283 VTAIL.n266 10.4732
R441 VTAIL.n214 VTAIL.n213 10.4732
R442 VTAIL.n194 VTAIL.n193 10.4732
R443 VTAIL.n169 VTAIL.n152 10.4732
R444 VTAIL.n392 VTAIL.n372 9.69747
R445 VTAIL.n412 VTAIL.n362 9.69747
R446 VTAIL.n441 VTAIL.n350 9.69747
R447 VTAIL.n50 VTAIL.n30 9.69747
R448 VTAIL.n70 VTAIL.n20 9.69747
R449 VTAIL.n99 VTAIL.n8 9.69747
R450 VTAIL.n331 VTAIL.n240 9.69747
R451 VTAIL.n304 VTAIL.n254 9.69747
R452 VTAIL.n284 VTAIL.n264 9.69747
R453 VTAIL.n217 VTAIL.n126 9.69747
R454 VTAIL.n190 VTAIL.n140 9.69747
R455 VTAIL.n170 VTAIL.n150 9.69747
R456 VTAIL.n452 VTAIL.n451 9.45567
R457 VTAIL.n110 VTAIL.n109 9.45567
R458 VTAIL.n342 VTAIL.n341 9.45567
R459 VTAIL.n228 VTAIL.n227 9.45567
R460 VTAIL.n451 VTAIL.n450 9.3005
R461 VTAIL.n445 VTAIL.n444 9.3005
R462 VTAIL.n443 VTAIL.n442 9.3005
R463 VTAIL.n350 VTAIL.n349 9.3005
R464 VTAIL.n437 VTAIL.n436 9.3005
R465 VTAIL.n435 VTAIL.n434 9.3005
R466 VTAIL.n354 VTAIL.n353 9.3005
R467 VTAIL.n429 VTAIL.n428 9.3005
R468 VTAIL.n401 VTAIL.n400 9.3005
R469 VTAIL.n370 VTAIL.n369 9.3005
R470 VTAIL.n395 VTAIL.n394 9.3005
R471 VTAIL.n393 VTAIL.n392 9.3005
R472 VTAIL.n374 VTAIL.n373 9.3005
R473 VTAIL.n387 VTAIL.n386 9.3005
R474 VTAIL.n385 VTAIL.n384 9.3005
R475 VTAIL.n378 VTAIL.n377 9.3005
R476 VTAIL.n403 VTAIL.n402 9.3005
R477 VTAIL.n366 VTAIL.n365 9.3005
R478 VTAIL.n409 VTAIL.n408 9.3005
R479 VTAIL.n411 VTAIL.n410 9.3005
R480 VTAIL.n362 VTAIL.n361 9.3005
R481 VTAIL.n417 VTAIL.n416 9.3005
R482 VTAIL.n419 VTAIL.n418 9.3005
R483 VTAIL.n420 VTAIL.n357 9.3005
R484 VTAIL.n427 VTAIL.n426 9.3005
R485 VTAIL.n346 VTAIL.n345 9.3005
R486 VTAIL.n109 VTAIL.n108 9.3005
R487 VTAIL.n103 VTAIL.n102 9.3005
R488 VTAIL.n101 VTAIL.n100 9.3005
R489 VTAIL.n8 VTAIL.n7 9.3005
R490 VTAIL.n95 VTAIL.n94 9.3005
R491 VTAIL.n93 VTAIL.n92 9.3005
R492 VTAIL.n12 VTAIL.n11 9.3005
R493 VTAIL.n87 VTAIL.n86 9.3005
R494 VTAIL.n59 VTAIL.n58 9.3005
R495 VTAIL.n28 VTAIL.n27 9.3005
R496 VTAIL.n53 VTAIL.n52 9.3005
R497 VTAIL.n51 VTAIL.n50 9.3005
R498 VTAIL.n32 VTAIL.n31 9.3005
R499 VTAIL.n45 VTAIL.n44 9.3005
R500 VTAIL.n43 VTAIL.n42 9.3005
R501 VTAIL.n36 VTAIL.n35 9.3005
R502 VTAIL.n61 VTAIL.n60 9.3005
R503 VTAIL.n24 VTAIL.n23 9.3005
R504 VTAIL.n67 VTAIL.n66 9.3005
R505 VTAIL.n69 VTAIL.n68 9.3005
R506 VTAIL.n20 VTAIL.n19 9.3005
R507 VTAIL.n75 VTAIL.n74 9.3005
R508 VTAIL.n77 VTAIL.n76 9.3005
R509 VTAIL.n78 VTAIL.n15 9.3005
R510 VTAIL.n85 VTAIL.n84 9.3005
R511 VTAIL.n4 VTAIL.n3 9.3005
R512 VTAIL.n258 VTAIL.n257 9.3005
R513 VTAIL.n301 VTAIL.n300 9.3005
R514 VTAIL.n303 VTAIL.n302 9.3005
R515 VTAIL.n254 VTAIL.n253 9.3005
R516 VTAIL.n309 VTAIL.n308 9.3005
R517 VTAIL.n311 VTAIL.n310 9.3005
R518 VTAIL.n249 VTAIL.n247 9.3005
R519 VTAIL.n317 VTAIL.n316 9.3005
R520 VTAIL.n341 VTAIL.n340 9.3005
R521 VTAIL.n236 VTAIL.n235 9.3005
R522 VTAIL.n335 VTAIL.n334 9.3005
R523 VTAIL.n333 VTAIL.n332 9.3005
R524 VTAIL.n240 VTAIL.n239 9.3005
R525 VTAIL.n327 VTAIL.n326 9.3005
R526 VTAIL.n325 VTAIL.n324 9.3005
R527 VTAIL.n244 VTAIL.n243 9.3005
R528 VTAIL.n319 VTAIL.n318 9.3005
R529 VTAIL.n295 VTAIL.n294 9.3005
R530 VTAIL.n293 VTAIL.n292 9.3005
R531 VTAIL.n262 VTAIL.n261 9.3005
R532 VTAIL.n287 VTAIL.n286 9.3005
R533 VTAIL.n285 VTAIL.n284 9.3005
R534 VTAIL.n266 VTAIL.n265 9.3005
R535 VTAIL.n279 VTAIL.n278 9.3005
R536 VTAIL.n277 VTAIL.n276 9.3005
R537 VTAIL.n270 VTAIL.n269 9.3005
R538 VTAIL.n144 VTAIL.n143 9.3005
R539 VTAIL.n187 VTAIL.n186 9.3005
R540 VTAIL.n189 VTAIL.n188 9.3005
R541 VTAIL.n140 VTAIL.n139 9.3005
R542 VTAIL.n195 VTAIL.n194 9.3005
R543 VTAIL.n197 VTAIL.n196 9.3005
R544 VTAIL.n135 VTAIL.n133 9.3005
R545 VTAIL.n203 VTAIL.n202 9.3005
R546 VTAIL.n227 VTAIL.n226 9.3005
R547 VTAIL.n122 VTAIL.n121 9.3005
R548 VTAIL.n221 VTAIL.n220 9.3005
R549 VTAIL.n219 VTAIL.n218 9.3005
R550 VTAIL.n126 VTAIL.n125 9.3005
R551 VTAIL.n213 VTAIL.n212 9.3005
R552 VTAIL.n211 VTAIL.n210 9.3005
R553 VTAIL.n130 VTAIL.n129 9.3005
R554 VTAIL.n205 VTAIL.n204 9.3005
R555 VTAIL.n181 VTAIL.n180 9.3005
R556 VTAIL.n179 VTAIL.n178 9.3005
R557 VTAIL.n148 VTAIL.n147 9.3005
R558 VTAIL.n173 VTAIL.n172 9.3005
R559 VTAIL.n171 VTAIL.n170 9.3005
R560 VTAIL.n152 VTAIL.n151 9.3005
R561 VTAIL.n165 VTAIL.n164 9.3005
R562 VTAIL.n163 VTAIL.n162 9.3005
R563 VTAIL.n156 VTAIL.n155 9.3005
R564 VTAIL.n396 VTAIL.n395 8.92171
R565 VTAIL.n411 VTAIL.n364 8.92171
R566 VTAIL.n442 VTAIL.n348 8.92171
R567 VTAIL.n54 VTAIL.n53 8.92171
R568 VTAIL.n69 VTAIL.n22 8.92171
R569 VTAIL.n100 VTAIL.n6 8.92171
R570 VTAIL.n332 VTAIL.n238 8.92171
R571 VTAIL.n303 VTAIL.n256 8.92171
R572 VTAIL.n288 VTAIL.n287 8.92171
R573 VTAIL.n218 VTAIL.n124 8.92171
R574 VTAIL.n189 VTAIL.n142 8.92171
R575 VTAIL.n174 VTAIL.n173 8.92171
R576 VTAIL.n399 VTAIL.n370 8.14595
R577 VTAIL.n408 VTAIL.n407 8.14595
R578 VTAIL.n446 VTAIL.n445 8.14595
R579 VTAIL.n57 VTAIL.n28 8.14595
R580 VTAIL.n66 VTAIL.n65 8.14595
R581 VTAIL.n104 VTAIL.n103 8.14595
R582 VTAIL.n336 VTAIL.n335 8.14595
R583 VTAIL.n300 VTAIL.n299 8.14595
R584 VTAIL.n291 VTAIL.n262 8.14595
R585 VTAIL.n222 VTAIL.n221 8.14595
R586 VTAIL.n186 VTAIL.n185 8.14595
R587 VTAIL.n177 VTAIL.n148 8.14595
R588 VTAIL.n400 VTAIL.n368 7.3702
R589 VTAIL.n404 VTAIL.n366 7.3702
R590 VTAIL.n449 VTAIL.n346 7.3702
R591 VTAIL.n452 VTAIL.n344 7.3702
R592 VTAIL.n58 VTAIL.n26 7.3702
R593 VTAIL.n62 VTAIL.n24 7.3702
R594 VTAIL.n107 VTAIL.n4 7.3702
R595 VTAIL.n110 VTAIL.n2 7.3702
R596 VTAIL.n342 VTAIL.n234 7.3702
R597 VTAIL.n339 VTAIL.n236 7.3702
R598 VTAIL.n296 VTAIL.n258 7.3702
R599 VTAIL.n292 VTAIL.n260 7.3702
R600 VTAIL.n228 VTAIL.n120 7.3702
R601 VTAIL.n225 VTAIL.n122 7.3702
R602 VTAIL.n182 VTAIL.n144 7.3702
R603 VTAIL.n178 VTAIL.n146 7.3702
R604 VTAIL.n403 VTAIL.n368 6.59444
R605 VTAIL.n404 VTAIL.n403 6.59444
R606 VTAIL.n450 VTAIL.n449 6.59444
R607 VTAIL.n450 VTAIL.n344 6.59444
R608 VTAIL.n61 VTAIL.n26 6.59444
R609 VTAIL.n62 VTAIL.n61 6.59444
R610 VTAIL.n108 VTAIL.n107 6.59444
R611 VTAIL.n108 VTAIL.n2 6.59444
R612 VTAIL.n340 VTAIL.n234 6.59444
R613 VTAIL.n340 VTAIL.n339 6.59444
R614 VTAIL.n296 VTAIL.n295 6.59444
R615 VTAIL.n295 VTAIL.n260 6.59444
R616 VTAIL.n226 VTAIL.n120 6.59444
R617 VTAIL.n226 VTAIL.n225 6.59444
R618 VTAIL.n182 VTAIL.n181 6.59444
R619 VTAIL.n181 VTAIL.n146 6.59444
R620 VTAIL.n400 VTAIL.n399 5.81868
R621 VTAIL.n407 VTAIL.n366 5.81868
R622 VTAIL.n446 VTAIL.n346 5.81868
R623 VTAIL.n58 VTAIL.n57 5.81868
R624 VTAIL.n65 VTAIL.n24 5.81868
R625 VTAIL.n104 VTAIL.n4 5.81868
R626 VTAIL.n336 VTAIL.n236 5.81868
R627 VTAIL.n299 VTAIL.n258 5.81868
R628 VTAIL.n292 VTAIL.n291 5.81868
R629 VTAIL.n222 VTAIL.n122 5.81868
R630 VTAIL.n185 VTAIL.n144 5.81868
R631 VTAIL.n178 VTAIL.n177 5.81868
R632 VTAIL.n396 VTAIL.n370 5.04292
R633 VTAIL.n408 VTAIL.n364 5.04292
R634 VTAIL.n445 VTAIL.n348 5.04292
R635 VTAIL.n54 VTAIL.n28 5.04292
R636 VTAIL.n66 VTAIL.n22 5.04292
R637 VTAIL.n103 VTAIL.n6 5.04292
R638 VTAIL.n335 VTAIL.n238 5.04292
R639 VTAIL.n300 VTAIL.n256 5.04292
R640 VTAIL.n288 VTAIL.n262 5.04292
R641 VTAIL.n221 VTAIL.n124 5.04292
R642 VTAIL.n186 VTAIL.n142 5.04292
R643 VTAIL.n174 VTAIL.n148 5.04292
R644 VTAIL.n379 VTAIL.n377 4.38563
R645 VTAIL.n37 VTAIL.n35 4.38563
R646 VTAIL.n271 VTAIL.n269 4.38563
R647 VTAIL.n157 VTAIL.n155 4.38563
R648 VTAIL.n395 VTAIL.n372 4.26717
R649 VTAIL.n412 VTAIL.n411 4.26717
R650 VTAIL.n442 VTAIL.n441 4.26717
R651 VTAIL.n53 VTAIL.n30 4.26717
R652 VTAIL.n70 VTAIL.n69 4.26717
R653 VTAIL.n100 VTAIL.n99 4.26717
R654 VTAIL.n332 VTAIL.n331 4.26717
R655 VTAIL.n304 VTAIL.n303 4.26717
R656 VTAIL.n287 VTAIL.n264 4.26717
R657 VTAIL.n218 VTAIL.n217 4.26717
R658 VTAIL.n190 VTAIL.n189 4.26717
R659 VTAIL.n173 VTAIL.n150 4.26717
R660 VTAIL.n392 VTAIL.n391 3.49141
R661 VTAIL.n415 VTAIL.n362 3.49141
R662 VTAIL.n438 VTAIL.n350 3.49141
R663 VTAIL.n50 VTAIL.n49 3.49141
R664 VTAIL.n73 VTAIL.n20 3.49141
R665 VTAIL.n96 VTAIL.n8 3.49141
R666 VTAIL.n328 VTAIL.n240 3.49141
R667 VTAIL.n307 VTAIL.n254 3.49141
R668 VTAIL.n284 VTAIL.n283 3.49141
R669 VTAIL.n214 VTAIL.n126 3.49141
R670 VTAIL.n193 VTAIL.n140 3.49141
R671 VTAIL.n170 VTAIL.n169 3.49141
R672 VTAIL.n119 VTAIL.n117 3.06947
R673 VTAIL.n229 VTAIL.n119 3.06947
R674 VTAIL.n233 VTAIL.n231 3.06947
R675 VTAIL.n343 VTAIL.n233 3.06947
R676 VTAIL.n115 VTAIL.n113 3.06947
R677 VTAIL.n113 VTAIL.n111 3.06947
R678 VTAIL.n455 VTAIL.n453 3.06947
R679 VTAIL.n388 VTAIL.n374 2.71565
R680 VTAIL.n416 VTAIL.n360 2.71565
R681 VTAIL.n437 VTAIL.n352 2.71565
R682 VTAIL.n46 VTAIL.n32 2.71565
R683 VTAIL.n74 VTAIL.n18 2.71565
R684 VTAIL.n95 VTAIL.n10 2.71565
R685 VTAIL.n327 VTAIL.n242 2.71565
R686 VTAIL.n308 VTAIL.n252 2.71565
R687 VTAIL.n280 VTAIL.n266 2.71565
R688 VTAIL.n213 VTAIL.n128 2.71565
R689 VTAIL.n194 VTAIL.n138 2.71565
R690 VTAIL.n166 VTAIL.n152 2.71565
R691 VTAIL VTAIL.n1 2.36041
R692 VTAIL.n231 VTAIL.n229 2.00481
R693 VTAIL.n111 VTAIL.n1 2.00481
R694 VTAIL.n387 VTAIL.n376 1.93989
R695 VTAIL.n421 VTAIL.n419 1.93989
R696 VTAIL.n434 VTAIL.n433 1.93989
R697 VTAIL.n45 VTAIL.n34 1.93989
R698 VTAIL.n79 VTAIL.n77 1.93989
R699 VTAIL.n92 VTAIL.n91 1.93989
R700 VTAIL.n324 VTAIL.n323 1.93989
R701 VTAIL.n312 VTAIL.n311 1.93989
R702 VTAIL.n279 VTAIL.n268 1.93989
R703 VTAIL.n210 VTAIL.n209 1.93989
R704 VTAIL.n198 VTAIL.n197 1.93989
R705 VTAIL.n165 VTAIL.n154 1.93989
R706 VTAIL.n384 VTAIL.n383 1.16414
R707 VTAIL.n420 VTAIL.n358 1.16414
R708 VTAIL.n430 VTAIL.n354 1.16414
R709 VTAIL.n42 VTAIL.n41 1.16414
R710 VTAIL.n78 VTAIL.n16 1.16414
R711 VTAIL.n88 VTAIL.n12 1.16414
R712 VTAIL.n320 VTAIL.n244 1.16414
R713 VTAIL.n315 VTAIL.n249 1.16414
R714 VTAIL.n276 VTAIL.n275 1.16414
R715 VTAIL.n206 VTAIL.n130 1.16414
R716 VTAIL.n201 VTAIL.n135 1.16414
R717 VTAIL.n162 VTAIL.n161 1.16414
R718 VTAIL.n454 VTAIL.t11 1.01174
R719 VTAIL.n454 VTAIL.t14 1.01174
R720 VTAIL.n0 VTAIL.t12 1.01174
R721 VTAIL.n0 VTAIL.t19 1.01174
R722 VTAIL.n112 VTAIL.t8 1.01174
R723 VTAIL.n112 VTAIL.t5 1.01174
R724 VTAIL.n114 VTAIL.t4 1.01174
R725 VTAIL.n114 VTAIL.t0 1.01174
R726 VTAIL.n232 VTAIL.t1 1.01174
R727 VTAIL.n232 VTAIL.t9 1.01174
R728 VTAIL.n230 VTAIL.t7 1.01174
R729 VTAIL.n230 VTAIL.t6 1.01174
R730 VTAIL.n118 VTAIL.t16 1.01174
R731 VTAIL.n118 VTAIL.t15 1.01174
R732 VTAIL.n116 VTAIL.t18 1.01174
R733 VTAIL.n116 VTAIL.t10 1.01174
R734 VTAIL VTAIL.n455 0.709552
R735 VTAIL.n380 VTAIL.n378 0.388379
R736 VTAIL.n426 VTAIL.n425 0.388379
R737 VTAIL.n429 VTAIL.n356 0.388379
R738 VTAIL.n38 VTAIL.n36 0.388379
R739 VTAIL.n84 VTAIL.n83 0.388379
R740 VTAIL.n87 VTAIL.n14 0.388379
R741 VTAIL.n319 VTAIL.n246 0.388379
R742 VTAIL.n316 VTAIL.n248 0.388379
R743 VTAIL.n272 VTAIL.n270 0.388379
R744 VTAIL.n205 VTAIL.n132 0.388379
R745 VTAIL.n202 VTAIL.n134 0.388379
R746 VTAIL.n158 VTAIL.n156 0.388379
R747 VTAIL.n385 VTAIL.n377 0.155672
R748 VTAIL.n386 VTAIL.n385 0.155672
R749 VTAIL.n386 VTAIL.n373 0.155672
R750 VTAIL.n393 VTAIL.n373 0.155672
R751 VTAIL.n394 VTAIL.n393 0.155672
R752 VTAIL.n394 VTAIL.n369 0.155672
R753 VTAIL.n401 VTAIL.n369 0.155672
R754 VTAIL.n402 VTAIL.n401 0.155672
R755 VTAIL.n402 VTAIL.n365 0.155672
R756 VTAIL.n409 VTAIL.n365 0.155672
R757 VTAIL.n410 VTAIL.n409 0.155672
R758 VTAIL.n410 VTAIL.n361 0.155672
R759 VTAIL.n417 VTAIL.n361 0.155672
R760 VTAIL.n418 VTAIL.n417 0.155672
R761 VTAIL.n418 VTAIL.n357 0.155672
R762 VTAIL.n427 VTAIL.n357 0.155672
R763 VTAIL.n428 VTAIL.n427 0.155672
R764 VTAIL.n428 VTAIL.n353 0.155672
R765 VTAIL.n435 VTAIL.n353 0.155672
R766 VTAIL.n436 VTAIL.n435 0.155672
R767 VTAIL.n436 VTAIL.n349 0.155672
R768 VTAIL.n443 VTAIL.n349 0.155672
R769 VTAIL.n444 VTAIL.n443 0.155672
R770 VTAIL.n444 VTAIL.n345 0.155672
R771 VTAIL.n451 VTAIL.n345 0.155672
R772 VTAIL.n43 VTAIL.n35 0.155672
R773 VTAIL.n44 VTAIL.n43 0.155672
R774 VTAIL.n44 VTAIL.n31 0.155672
R775 VTAIL.n51 VTAIL.n31 0.155672
R776 VTAIL.n52 VTAIL.n51 0.155672
R777 VTAIL.n52 VTAIL.n27 0.155672
R778 VTAIL.n59 VTAIL.n27 0.155672
R779 VTAIL.n60 VTAIL.n59 0.155672
R780 VTAIL.n60 VTAIL.n23 0.155672
R781 VTAIL.n67 VTAIL.n23 0.155672
R782 VTAIL.n68 VTAIL.n67 0.155672
R783 VTAIL.n68 VTAIL.n19 0.155672
R784 VTAIL.n75 VTAIL.n19 0.155672
R785 VTAIL.n76 VTAIL.n75 0.155672
R786 VTAIL.n76 VTAIL.n15 0.155672
R787 VTAIL.n85 VTAIL.n15 0.155672
R788 VTAIL.n86 VTAIL.n85 0.155672
R789 VTAIL.n86 VTAIL.n11 0.155672
R790 VTAIL.n93 VTAIL.n11 0.155672
R791 VTAIL.n94 VTAIL.n93 0.155672
R792 VTAIL.n94 VTAIL.n7 0.155672
R793 VTAIL.n101 VTAIL.n7 0.155672
R794 VTAIL.n102 VTAIL.n101 0.155672
R795 VTAIL.n102 VTAIL.n3 0.155672
R796 VTAIL.n109 VTAIL.n3 0.155672
R797 VTAIL.n341 VTAIL.n235 0.155672
R798 VTAIL.n334 VTAIL.n235 0.155672
R799 VTAIL.n334 VTAIL.n333 0.155672
R800 VTAIL.n333 VTAIL.n239 0.155672
R801 VTAIL.n326 VTAIL.n239 0.155672
R802 VTAIL.n326 VTAIL.n325 0.155672
R803 VTAIL.n325 VTAIL.n243 0.155672
R804 VTAIL.n318 VTAIL.n243 0.155672
R805 VTAIL.n318 VTAIL.n317 0.155672
R806 VTAIL.n317 VTAIL.n247 0.155672
R807 VTAIL.n310 VTAIL.n247 0.155672
R808 VTAIL.n310 VTAIL.n309 0.155672
R809 VTAIL.n309 VTAIL.n253 0.155672
R810 VTAIL.n302 VTAIL.n253 0.155672
R811 VTAIL.n302 VTAIL.n301 0.155672
R812 VTAIL.n301 VTAIL.n257 0.155672
R813 VTAIL.n294 VTAIL.n257 0.155672
R814 VTAIL.n294 VTAIL.n293 0.155672
R815 VTAIL.n293 VTAIL.n261 0.155672
R816 VTAIL.n286 VTAIL.n261 0.155672
R817 VTAIL.n286 VTAIL.n285 0.155672
R818 VTAIL.n285 VTAIL.n265 0.155672
R819 VTAIL.n278 VTAIL.n265 0.155672
R820 VTAIL.n278 VTAIL.n277 0.155672
R821 VTAIL.n277 VTAIL.n269 0.155672
R822 VTAIL.n227 VTAIL.n121 0.155672
R823 VTAIL.n220 VTAIL.n121 0.155672
R824 VTAIL.n220 VTAIL.n219 0.155672
R825 VTAIL.n219 VTAIL.n125 0.155672
R826 VTAIL.n212 VTAIL.n125 0.155672
R827 VTAIL.n212 VTAIL.n211 0.155672
R828 VTAIL.n211 VTAIL.n129 0.155672
R829 VTAIL.n204 VTAIL.n129 0.155672
R830 VTAIL.n204 VTAIL.n203 0.155672
R831 VTAIL.n203 VTAIL.n133 0.155672
R832 VTAIL.n196 VTAIL.n133 0.155672
R833 VTAIL.n196 VTAIL.n195 0.155672
R834 VTAIL.n195 VTAIL.n139 0.155672
R835 VTAIL.n188 VTAIL.n139 0.155672
R836 VTAIL.n188 VTAIL.n187 0.155672
R837 VTAIL.n187 VTAIL.n143 0.155672
R838 VTAIL.n180 VTAIL.n143 0.155672
R839 VTAIL.n180 VTAIL.n179 0.155672
R840 VTAIL.n179 VTAIL.n147 0.155672
R841 VTAIL.n172 VTAIL.n147 0.155672
R842 VTAIL.n172 VTAIL.n171 0.155672
R843 VTAIL.n171 VTAIL.n151 0.155672
R844 VTAIL.n164 VTAIL.n151 0.155672
R845 VTAIL.n164 VTAIL.n163 0.155672
R846 VTAIL.n163 VTAIL.n155 0.155672
R847 VDD2.n217 VDD2.n113 289.615
R848 VDD2.n104 VDD2.n0 289.615
R849 VDD2.n218 VDD2.n217 185
R850 VDD2.n216 VDD2.n215 185
R851 VDD2.n117 VDD2.n116 185
R852 VDD2.n210 VDD2.n209 185
R853 VDD2.n208 VDD2.n207 185
R854 VDD2.n121 VDD2.n120 185
R855 VDD2.n202 VDD2.n201 185
R856 VDD2.n200 VDD2.n199 185
R857 VDD2.n125 VDD2.n124 185
R858 VDD2.n129 VDD2.n127 185
R859 VDD2.n194 VDD2.n193 185
R860 VDD2.n192 VDD2.n191 185
R861 VDD2.n131 VDD2.n130 185
R862 VDD2.n186 VDD2.n185 185
R863 VDD2.n184 VDD2.n183 185
R864 VDD2.n135 VDD2.n134 185
R865 VDD2.n178 VDD2.n177 185
R866 VDD2.n176 VDD2.n175 185
R867 VDD2.n139 VDD2.n138 185
R868 VDD2.n170 VDD2.n169 185
R869 VDD2.n168 VDD2.n167 185
R870 VDD2.n143 VDD2.n142 185
R871 VDD2.n162 VDD2.n161 185
R872 VDD2.n160 VDD2.n159 185
R873 VDD2.n147 VDD2.n146 185
R874 VDD2.n154 VDD2.n153 185
R875 VDD2.n152 VDD2.n151 185
R876 VDD2.n37 VDD2.n36 185
R877 VDD2.n39 VDD2.n38 185
R878 VDD2.n32 VDD2.n31 185
R879 VDD2.n45 VDD2.n44 185
R880 VDD2.n47 VDD2.n46 185
R881 VDD2.n28 VDD2.n27 185
R882 VDD2.n53 VDD2.n52 185
R883 VDD2.n55 VDD2.n54 185
R884 VDD2.n24 VDD2.n23 185
R885 VDD2.n61 VDD2.n60 185
R886 VDD2.n63 VDD2.n62 185
R887 VDD2.n20 VDD2.n19 185
R888 VDD2.n69 VDD2.n68 185
R889 VDD2.n71 VDD2.n70 185
R890 VDD2.n16 VDD2.n15 185
R891 VDD2.n78 VDD2.n77 185
R892 VDD2.n79 VDD2.n14 185
R893 VDD2.n81 VDD2.n80 185
R894 VDD2.n12 VDD2.n11 185
R895 VDD2.n87 VDD2.n86 185
R896 VDD2.n89 VDD2.n88 185
R897 VDD2.n8 VDD2.n7 185
R898 VDD2.n95 VDD2.n94 185
R899 VDD2.n97 VDD2.n96 185
R900 VDD2.n4 VDD2.n3 185
R901 VDD2.n103 VDD2.n102 185
R902 VDD2.n105 VDD2.n104 185
R903 VDD2.n150 VDD2.t6 147.659
R904 VDD2.n35 VDD2.t7 147.659
R905 VDD2.n217 VDD2.n216 104.615
R906 VDD2.n216 VDD2.n116 104.615
R907 VDD2.n209 VDD2.n116 104.615
R908 VDD2.n209 VDD2.n208 104.615
R909 VDD2.n208 VDD2.n120 104.615
R910 VDD2.n201 VDD2.n120 104.615
R911 VDD2.n201 VDD2.n200 104.615
R912 VDD2.n200 VDD2.n124 104.615
R913 VDD2.n129 VDD2.n124 104.615
R914 VDD2.n193 VDD2.n129 104.615
R915 VDD2.n193 VDD2.n192 104.615
R916 VDD2.n192 VDD2.n130 104.615
R917 VDD2.n185 VDD2.n130 104.615
R918 VDD2.n185 VDD2.n184 104.615
R919 VDD2.n184 VDD2.n134 104.615
R920 VDD2.n177 VDD2.n134 104.615
R921 VDD2.n177 VDD2.n176 104.615
R922 VDD2.n176 VDD2.n138 104.615
R923 VDD2.n169 VDD2.n138 104.615
R924 VDD2.n169 VDD2.n168 104.615
R925 VDD2.n168 VDD2.n142 104.615
R926 VDD2.n161 VDD2.n142 104.615
R927 VDD2.n161 VDD2.n160 104.615
R928 VDD2.n160 VDD2.n146 104.615
R929 VDD2.n153 VDD2.n146 104.615
R930 VDD2.n153 VDD2.n152 104.615
R931 VDD2.n38 VDD2.n37 104.615
R932 VDD2.n38 VDD2.n31 104.615
R933 VDD2.n45 VDD2.n31 104.615
R934 VDD2.n46 VDD2.n45 104.615
R935 VDD2.n46 VDD2.n27 104.615
R936 VDD2.n53 VDD2.n27 104.615
R937 VDD2.n54 VDD2.n53 104.615
R938 VDD2.n54 VDD2.n23 104.615
R939 VDD2.n61 VDD2.n23 104.615
R940 VDD2.n62 VDD2.n61 104.615
R941 VDD2.n62 VDD2.n19 104.615
R942 VDD2.n69 VDD2.n19 104.615
R943 VDD2.n70 VDD2.n69 104.615
R944 VDD2.n70 VDD2.n15 104.615
R945 VDD2.n78 VDD2.n15 104.615
R946 VDD2.n79 VDD2.n78 104.615
R947 VDD2.n80 VDD2.n79 104.615
R948 VDD2.n80 VDD2.n11 104.615
R949 VDD2.n87 VDD2.n11 104.615
R950 VDD2.n88 VDD2.n87 104.615
R951 VDD2.n88 VDD2.n7 104.615
R952 VDD2.n95 VDD2.n7 104.615
R953 VDD2.n96 VDD2.n95 104.615
R954 VDD2.n96 VDD2.n3 104.615
R955 VDD2.n103 VDD2.n3 104.615
R956 VDD2.n104 VDD2.n103 104.615
R957 VDD2.n112 VDD2.n111 60.909
R958 VDD2 VDD2.n225 60.9061
R959 VDD2.n224 VDD2.n223 58.6628
R960 VDD2.n110 VDD2.n109 58.6626
R961 VDD2.n222 VDD2.n112 55.1722
R962 VDD2.n152 VDD2.t6 52.3082
R963 VDD2.n37 VDD2.t7 52.3082
R964 VDD2.n110 VDD2.n108 49.9937
R965 VDD2.n222 VDD2.n221 46.9247
R966 VDD2.n151 VDD2.n150 15.6677
R967 VDD2.n36 VDD2.n35 15.6677
R968 VDD2.n127 VDD2.n125 13.1884
R969 VDD2.n81 VDD2.n12 13.1884
R970 VDD2.n199 VDD2.n198 12.8005
R971 VDD2.n195 VDD2.n194 12.8005
R972 VDD2.n154 VDD2.n149 12.8005
R973 VDD2.n39 VDD2.n34 12.8005
R974 VDD2.n82 VDD2.n14 12.8005
R975 VDD2.n86 VDD2.n85 12.8005
R976 VDD2.n202 VDD2.n123 12.0247
R977 VDD2.n191 VDD2.n128 12.0247
R978 VDD2.n155 VDD2.n147 12.0247
R979 VDD2.n40 VDD2.n32 12.0247
R980 VDD2.n77 VDD2.n76 12.0247
R981 VDD2.n89 VDD2.n10 12.0247
R982 VDD2.n203 VDD2.n121 11.249
R983 VDD2.n190 VDD2.n131 11.249
R984 VDD2.n159 VDD2.n158 11.249
R985 VDD2.n44 VDD2.n43 11.249
R986 VDD2.n75 VDD2.n16 11.249
R987 VDD2.n90 VDD2.n8 11.249
R988 VDD2.n207 VDD2.n206 10.4732
R989 VDD2.n187 VDD2.n186 10.4732
R990 VDD2.n162 VDD2.n145 10.4732
R991 VDD2.n47 VDD2.n30 10.4732
R992 VDD2.n72 VDD2.n71 10.4732
R993 VDD2.n94 VDD2.n93 10.4732
R994 VDD2.n210 VDD2.n119 9.69747
R995 VDD2.n183 VDD2.n133 9.69747
R996 VDD2.n163 VDD2.n143 9.69747
R997 VDD2.n48 VDD2.n28 9.69747
R998 VDD2.n68 VDD2.n18 9.69747
R999 VDD2.n97 VDD2.n6 9.69747
R1000 VDD2.n221 VDD2.n220 9.45567
R1001 VDD2.n108 VDD2.n107 9.45567
R1002 VDD2.n137 VDD2.n136 9.3005
R1003 VDD2.n180 VDD2.n179 9.3005
R1004 VDD2.n182 VDD2.n181 9.3005
R1005 VDD2.n133 VDD2.n132 9.3005
R1006 VDD2.n188 VDD2.n187 9.3005
R1007 VDD2.n190 VDD2.n189 9.3005
R1008 VDD2.n128 VDD2.n126 9.3005
R1009 VDD2.n196 VDD2.n195 9.3005
R1010 VDD2.n220 VDD2.n219 9.3005
R1011 VDD2.n115 VDD2.n114 9.3005
R1012 VDD2.n214 VDD2.n213 9.3005
R1013 VDD2.n212 VDD2.n211 9.3005
R1014 VDD2.n119 VDD2.n118 9.3005
R1015 VDD2.n206 VDD2.n205 9.3005
R1016 VDD2.n204 VDD2.n203 9.3005
R1017 VDD2.n123 VDD2.n122 9.3005
R1018 VDD2.n198 VDD2.n197 9.3005
R1019 VDD2.n174 VDD2.n173 9.3005
R1020 VDD2.n172 VDD2.n171 9.3005
R1021 VDD2.n141 VDD2.n140 9.3005
R1022 VDD2.n166 VDD2.n165 9.3005
R1023 VDD2.n164 VDD2.n163 9.3005
R1024 VDD2.n145 VDD2.n144 9.3005
R1025 VDD2.n158 VDD2.n157 9.3005
R1026 VDD2.n156 VDD2.n155 9.3005
R1027 VDD2.n149 VDD2.n148 9.3005
R1028 VDD2.n107 VDD2.n106 9.3005
R1029 VDD2.n101 VDD2.n100 9.3005
R1030 VDD2.n99 VDD2.n98 9.3005
R1031 VDD2.n6 VDD2.n5 9.3005
R1032 VDD2.n93 VDD2.n92 9.3005
R1033 VDD2.n91 VDD2.n90 9.3005
R1034 VDD2.n10 VDD2.n9 9.3005
R1035 VDD2.n85 VDD2.n84 9.3005
R1036 VDD2.n57 VDD2.n56 9.3005
R1037 VDD2.n26 VDD2.n25 9.3005
R1038 VDD2.n51 VDD2.n50 9.3005
R1039 VDD2.n49 VDD2.n48 9.3005
R1040 VDD2.n30 VDD2.n29 9.3005
R1041 VDD2.n43 VDD2.n42 9.3005
R1042 VDD2.n41 VDD2.n40 9.3005
R1043 VDD2.n34 VDD2.n33 9.3005
R1044 VDD2.n59 VDD2.n58 9.3005
R1045 VDD2.n22 VDD2.n21 9.3005
R1046 VDD2.n65 VDD2.n64 9.3005
R1047 VDD2.n67 VDD2.n66 9.3005
R1048 VDD2.n18 VDD2.n17 9.3005
R1049 VDD2.n73 VDD2.n72 9.3005
R1050 VDD2.n75 VDD2.n74 9.3005
R1051 VDD2.n76 VDD2.n13 9.3005
R1052 VDD2.n83 VDD2.n82 9.3005
R1053 VDD2.n2 VDD2.n1 9.3005
R1054 VDD2.n211 VDD2.n117 8.92171
R1055 VDD2.n182 VDD2.n135 8.92171
R1056 VDD2.n167 VDD2.n166 8.92171
R1057 VDD2.n52 VDD2.n51 8.92171
R1058 VDD2.n67 VDD2.n20 8.92171
R1059 VDD2.n98 VDD2.n4 8.92171
R1060 VDD2.n215 VDD2.n214 8.14595
R1061 VDD2.n179 VDD2.n178 8.14595
R1062 VDD2.n170 VDD2.n141 8.14595
R1063 VDD2.n55 VDD2.n26 8.14595
R1064 VDD2.n64 VDD2.n63 8.14595
R1065 VDD2.n102 VDD2.n101 8.14595
R1066 VDD2.n221 VDD2.n113 7.3702
R1067 VDD2.n218 VDD2.n115 7.3702
R1068 VDD2.n175 VDD2.n137 7.3702
R1069 VDD2.n171 VDD2.n139 7.3702
R1070 VDD2.n56 VDD2.n24 7.3702
R1071 VDD2.n60 VDD2.n22 7.3702
R1072 VDD2.n105 VDD2.n2 7.3702
R1073 VDD2.n108 VDD2.n0 7.3702
R1074 VDD2.n219 VDD2.n113 6.59444
R1075 VDD2.n219 VDD2.n218 6.59444
R1076 VDD2.n175 VDD2.n174 6.59444
R1077 VDD2.n174 VDD2.n139 6.59444
R1078 VDD2.n59 VDD2.n24 6.59444
R1079 VDD2.n60 VDD2.n59 6.59444
R1080 VDD2.n106 VDD2.n105 6.59444
R1081 VDD2.n106 VDD2.n0 6.59444
R1082 VDD2.n215 VDD2.n115 5.81868
R1083 VDD2.n178 VDD2.n137 5.81868
R1084 VDD2.n171 VDD2.n170 5.81868
R1085 VDD2.n56 VDD2.n55 5.81868
R1086 VDD2.n63 VDD2.n22 5.81868
R1087 VDD2.n102 VDD2.n2 5.81868
R1088 VDD2.n214 VDD2.n117 5.04292
R1089 VDD2.n179 VDD2.n135 5.04292
R1090 VDD2.n167 VDD2.n141 5.04292
R1091 VDD2.n52 VDD2.n26 5.04292
R1092 VDD2.n64 VDD2.n20 5.04292
R1093 VDD2.n101 VDD2.n4 5.04292
R1094 VDD2.n150 VDD2.n148 4.38563
R1095 VDD2.n35 VDD2.n33 4.38563
R1096 VDD2.n211 VDD2.n210 4.26717
R1097 VDD2.n183 VDD2.n182 4.26717
R1098 VDD2.n166 VDD2.n143 4.26717
R1099 VDD2.n51 VDD2.n28 4.26717
R1100 VDD2.n68 VDD2.n67 4.26717
R1101 VDD2.n98 VDD2.n97 4.26717
R1102 VDD2.n207 VDD2.n119 3.49141
R1103 VDD2.n186 VDD2.n133 3.49141
R1104 VDD2.n163 VDD2.n162 3.49141
R1105 VDD2.n48 VDD2.n47 3.49141
R1106 VDD2.n71 VDD2.n18 3.49141
R1107 VDD2.n94 VDD2.n6 3.49141
R1108 VDD2.n224 VDD2.n222 3.06947
R1109 VDD2.n206 VDD2.n121 2.71565
R1110 VDD2.n187 VDD2.n131 2.71565
R1111 VDD2.n159 VDD2.n145 2.71565
R1112 VDD2.n44 VDD2.n30 2.71565
R1113 VDD2.n72 VDD2.n16 2.71565
R1114 VDD2.n93 VDD2.n8 2.71565
R1115 VDD2.n203 VDD2.n202 1.93989
R1116 VDD2.n191 VDD2.n190 1.93989
R1117 VDD2.n158 VDD2.n147 1.93989
R1118 VDD2.n43 VDD2.n32 1.93989
R1119 VDD2.n77 VDD2.n75 1.93989
R1120 VDD2.n90 VDD2.n89 1.93989
R1121 VDD2.n199 VDD2.n123 1.16414
R1122 VDD2.n194 VDD2.n128 1.16414
R1123 VDD2.n155 VDD2.n154 1.16414
R1124 VDD2.n40 VDD2.n39 1.16414
R1125 VDD2.n76 VDD2.n14 1.16414
R1126 VDD2.n86 VDD2.n10 1.16414
R1127 VDD2.n225 VDD2.t1 1.01174
R1128 VDD2.n225 VDD2.t2 1.01174
R1129 VDD2.n223 VDD2.t5 1.01174
R1130 VDD2.n223 VDD2.t0 1.01174
R1131 VDD2.n111 VDD2.t4 1.01174
R1132 VDD2.n111 VDD2.t9 1.01174
R1133 VDD2.n109 VDD2.t3 1.01174
R1134 VDD2.n109 VDD2.t8 1.01174
R1135 VDD2 VDD2.n224 0.825931
R1136 VDD2.n112 VDD2.n110 0.712395
R1137 VDD2.n198 VDD2.n125 0.388379
R1138 VDD2.n195 VDD2.n127 0.388379
R1139 VDD2.n151 VDD2.n149 0.388379
R1140 VDD2.n36 VDD2.n34 0.388379
R1141 VDD2.n82 VDD2.n81 0.388379
R1142 VDD2.n85 VDD2.n12 0.388379
R1143 VDD2.n220 VDD2.n114 0.155672
R1144 VDD2.n213 VDD2.n114 0.155672
R1145 VDD2.n213 VDD2.n212 0.155672
R1146 VDD2.n212 VDD2.n118 0.155672
R1147 VDD2.n205 VDD2.n118 0.155672
R1148 VDD2.n205 VDD2.n204 0.155672
R1149 VDD2.n204 VDD2.n122 0.155672
R1150 VDD2.n197 VDD2.n122 0.155672
R1151 VDD2.n197 VDD2.n196 0.155672
R1152 VDD2.n196 VDD2.n126 0.155672
R1153 VDD2.n189 VDD2.n126 0.155672
R1154 VDD2.n189 VDD2.n188 0.155672
R1155 VDD2.n188 VDD2.n132 0.155672
R1156 VDD2.n181 VDD2.n132 0.155672
R1157 VDD2.n181 VDD2.n180 0.155672
R1158 VDD2.n180 VDD2.n136 0.155672
R1159 VDD2.n173 VDD2.n136 0.155672
R1160 VDD2.n173 VDD2.n172 0.155672
R1161 VDD2.n172 VDD2.n140 0.155672
R1162 VDD2.n165 VDD2.n140 0.155672
R1163 VDD2.n165 VDD2.n164 0.155672
R1164 VDD2.n164 VDD2.n144 0.155672
R1165 VDD2.n157 VDD2.n144 0.155672
R1166 VDD2.n157 VDD2.n156 0.155672
R1167 VDD2.n156 VDD2.n148 0.155672
R1168 VDD2.n41 VDD2.n33 0.155672
R1169 VDD2.n42 VDD2.n41 0.155672
R1170 VDD2.n42 VDD2.n29 0.155672
R1171 VDD2.n49 VDD2.n29 0.155672
R1172 VDD2.n50 VDD2.n49 0.155672
R1173 VDD2.n50 VDD2.n25 0.155672
R1174 VDD2.n57 VDD2.n25 0.155672
R1175 VDD2.n58 VDD2.n57 0.155672
R1176 VDD2.n58 VDD2.n21 0.155672
R1177 VDD2.n65 VDD2.n21 0.155672
R1178 VDD2.n66 VDD2.n65 0.155672
R1179 VDD2.n66 VDD2.n17 0.155672
R1180 VDD2.n73 VDD2.n17 0.155672
R1181 VDD2.n74 VDD2.n73 0.155672
R1182 VDD2.n74 VDD2.n13 0.155672
R1183 VDD2.n83 VDD2.n13 0.155672
R1184 VDD2.n84 VDD2.n83 0.155672
R1185 VDD2.n84 VDD2.n9 0.155672
R1186 VDD2.n91 VDD2.n9 0.155672
R1187 VDD2.n92 VDD2.n91 0.155672
R1188 VDD2.n92 VDD2.n5 0.155672
R1189 VDD2.n99 VDD2.n5 0.155672
R1190 VDD2.n100 VDD2.n99 0.155672
R1191 VDD2.n100 VDD2.n1 0.155672
R1192 VDD2.n107 VDD2.n1 0.155672
R1193 B.n1264 B.n1263 585
R1194 B.n1265 B.n1264 585
R1195 B.n472 B.n198 585
R1196 B.n471 B.n470 585
R1197 B.n469 B.n468 585
R1198 B.n467 B.n466 585
R1199 B.n465 B.n464 585
R1200 B.n463 B.n462 585
R1201 B.n461 B.n460 585
R1202 B.n459 B.n458 585
R1203 B.n457 B.n456 585
R1204 B.n455 B.n454 585
R1205 B.n453 B.n452 585
R1206 B.n451 B.n450 585
R1207 B.n449 B.n448 585
R1208 B.n447 B.n446 585
R1209 B.n445 B.n444 585
R1210 B.n443 B.n442 585
R1211 B.n441 B.n440 585
R1212 B.n439 B.n438 585
R1213 B.n437 B.n436 585
R1214 B.n435 B.n434 585
R1215 B.n433 B.n432 585
R1216 B.n431 B.n430 585
R1217 B.n429 B.n428 585
R1218 B.n427 B.n426 585
R1219 B.n425 B.n424 585
R1220 B.n423 B.n422 585
R1221 B.n421 B.n420 585
R1222 B.n419 B.n418 585
R1223 B.n417 B.n416 585
R1224 B.n415 B.n414 585
R1225 B.n413 B.n412 585
R1226 B.n411 B.n410 585
R1227 B.n409 B.n408 585
R1228 B.n407 B.n406 585
R1229 B.n405 B.n404 585
R1230 B.n403 B.n402 585
R1231 B.n401 B.n400 585
R1232 B.n399 B.n398 585
R1233 B.n397 B.n396 585
R1234 B.n395 B.n394 585
R1235 B.n393 B.n392 585
R1236 B.n391 B.n390 585
R1237 B.n389 B.n388 585
R1238 B.n387 B.n386 585
R1239 B.n385 B.n384 585
R1240 B.n383 B.n382 585
R1241 B.n381 B.n380 585
R1242 B.n379 B.n378 585
R1243 B.n377 B.n376 585
R1244 B.n375 B.n374 585
R1245 B.n373 B.n372 585
R1246 B.n371 B.n370 585
R1247 B.n369 B.n368 585
R1248 B.n367 B.n366 585
R1249 B.n365 B.n364 585
R1250 B.n363 B.n362 585
R1251 B.n361 B.n360 585
R1252 B.n359 B.n358 585
R1253 B.n357 B.n356 585
R1254 B.n355 B.n354 585
R1255 B.n353 B.n352 585
R1256 B.n351 B.n350 585
R1257 B.n349 B.n348 585
R1258 B.n346 B.n345 585
R1259 B.n344 B.n343 585
R1260 B.n342 B.n341 585
R1261 B.n340 B.n339 585
R1262 B.n338 B.n337 585
R1263 B.n336 B.n335 585
R1264 B.n334 B.n333 585
R1265 B.n332 B.n331 585
R1266 B.n330 B.n329 585
R1267 B.n328 B.n327 585
R1268 B.n326 B.n325 585
R1269 B.n324 B.n323 585
R1270 B.n322 B.n321 585
R1271 B.n320 B.n319 585
R1272 B.n318 B.n317 585
R1273 B.n316 B.n315 585
R1274 B.n314 B.n313 585
R1275 B.n312 B.n311 585
R1276 B.n310 B.n309 585
R1277 B.n308 B.n307 585
R1278 B.n306 B.n305 585
R1279 B.n304 B.n303 585
R1280 B.n302 B.n301 585
R1281 B.n300 B.n299 585
R1282 B.n298 B.n297 585
R1283 B.n296 B.n295 585
R1284 B.n294 B.n293 585
R1285 B.n292 B.n291 585
R1286 B.n290 B.n289 585
R1287 B.n288 B.n287 585
R1288 B.n286 B.n285 585
R1289 B.n284 B.n283 585
R1290 B.n282 B.n281 585
R1291 B.n280 B.n279 585
R1292 B.n278 B.n277 585
R1293 B.n276 B.n275 585
R1294 B.n274 B.n273 585
R1295 B.n272 B.n271 585
R1296 B.n270 B.n269 585
R1297 B.n268 B.n267 585
R1298 B.n266 B.n265 585
R1299 B.n264 B.n263 585
R1300 B.n262 B.n261 585
R1301 B.n260 B.n259 585
R1302 B.n258 B.n257 585
R1303 B.n256 B.n255 585
R1304 B.n254 B.n253 585
R1305 B.n252 B.n251 585
R1306 B.n250 B.n249 585
R1307 B.n248 B.n247 585
R1308 B.n246 B.n245 585
R1309 B.n244 B.n243 585
R1310 B.n242 B.n241 585
R1311 B.n240 B.n239 585
R1312 B.n238 B.n237 585
R1313 B.n236 B.n235 585
R1314 B.n234 B.n233 585
R1315 B.n232 B.n231 585
R1316 B.n230 B.n229 585
R1317 B.n228 B.n227 585
R1318 B.n226 B.n225 585
R1319 B.n224 B.n223 585
R1320 B.n222 B.n221 585
R1321 B.n220 B.n219 585
R1322 B.n218 B.n217 585
R1323 B.n216 B.n215 585
R1324 B.n214 B.n213 585
R1325 B.n212 B.n211 585
R1326 B.n210 B.n209 585
R1327 B.n208 B.n207 585
R1328 B.n206 B.n205 585
R1329 B.n130 B.n129 585
R1330 B.n1268 B.n1267 585
R1331 B.n1262 B.n199 585
R1332 B.n199 B.n127 585
R1333 B.n1261 B.n126 585
R1334 B.n1272 B.n126 585
R1335 B.n1260 B.n125 585
R1336 B.n1273 B.n125 585
R1337 B.n1259 B.n124 585
R1338 B.n1274 B.n124 585
R1339 B.n1258 B.n1257 585
R1340 B.n1257 B.n120 585
R1341 B.n1256 B.n119 585
R1342 B.n1280 B.n119 585
R1343 B.n1255 B.n118 585
R1344 B.n1281 B.n118 585
R1345 B.n1254 B.n117 585
R1346 B.n1282 B.n117 585
R1347 B.n1253 B.n1252 585
R1348 B.n1252 B.n116 585
R1349 B.n1251 B.n112 585
R1350 B.n1288 B.n112 585
R1351 B.n1250 B.n111 585
R1352 B.n1289 B.n111 585
R1353 B.n1249 B.n110 585
R1354 B.n1290 B.n110 585
R1355 B.n1248 B.n1247 585
R1356 B.n1247 B.n106 585
R1357 B.n1246 B.n105 585
R1358 B.n1296 B.n105 585
R1359 B.n1245 B.n104 585
R1360 B.n1297 B.n104 585
R1361 B.n1244 B.n103 585
R1362 B.n1298 B.n103 585
R1363 B.n1243 B.n1242 585
R1364 B.n1242 B.n99 585
R1365 B.n1241 B.n98 585
R1366 B.n1304 B.n98 585
R1367 B.n1240 B.n97 585
R1368 B.n1305 B.n97 585
R1369 B.n1239 B.n96 585
R1370 B.n1306 B.n96 585
R1371 B.n1238 B.n1237 585
R1372 B.n1237 B.n92 585
R1373 B.n1236 B.n91 585
R1374 B.n1312 B.n91 585
R1375 B.n1235 B.n90 585
R1376 B.n1313 B.n90 585
R1377 B.n1234 B.n89 585
R1378 B.n1314 B.n89 585
R1379 B.n1233 B.n1232 585
R1380 B.n1232 B.n85 585
R1381 B.n1231 B.n84 585
R1382 B.n1320 B.n84 585
R1383 B.n1230 B.n83 585
R1384 B.n1321 B.n83 585
R1385 B.n1229 B.n82 585
R1386 B.n1322 B.n82 585
R1387 B.n1228 B.n1227 585
R1388 B.n1227 B.n78 585
R1389 B.n1226 B.n77 585
R1390 B.n1328 B.n77 585
R1391 B.n1225 B.n76 585
R1392 B.n1329 B.n76 585
R1393 B.n1224 B.n75 585
R1394 B.n1330 B.n75 585
R1395 B.n1223 B.n1222 585
R1396 B.n1222 B.n74 585
R1397 B.n1221 B.n70 585
R1398 B.n1336 B.n70 585
R1399 B.n1220 B.n69 585
R1400 B.n1337 B.n69 585
R1401 B.n1219 B.n68 585
R1402 B.n1338 B.n68 585
R1403 B.n1218 B.n1217 585
R1404 B.n1217 B.n64 585
R1405 B.n1216 B.n63 585
R1406 B.n1344 B.n63 585
R1407 B.n1215 B.n62 585
R1408 B.n1345 B.n62 585
R1409 B.n1214 B.n61 585
R1410 B.n1346 B.n61 585
R1411 B.n1213 B.n1212 585
R1412 B.n1212 B.n57 585
R1413 B.n1211 B.n56 585
R1414 B.n1352 B.n56 585
R1415 B.n1210 B.n55 585
R1416 B.n1353 B.n55 585
R1417 B.n1209 B.n54 585
R1418 B.n1354 B.n54 585
R1419 B.n1208 B.n1207 585
R1420 B.n1207 B.n50 585
R1421 B.n1206 B.n49 585
R1422 B.n1360 B.n49 585
R1423 B.n1205 B.n48 585
R1424 B.n1361 B.n48 585
R1425 B.n1204 B.n47 585
R1426 B.n1362 B.n47 585
R1427 B.n1203 B.n1202 585
R1428 B.n1202 B.n43 585
R1429 B.n1201 B.n42 585
R1430 B.n1368 B.n42 585
R1431 B.n1200 B.n41 585
R1432 B.n1369 B.n41 585
R1433 B.n1199 B.n40 585
R1434 B.n1370 B.n40 585
R1435 B.n1198 B.n1197 585
R1436 B.n1197 B.n36 585
R1437 B.n1196 B.n35 585
R1438 B.n1376 B.n35 585
R1439 B.n1195 B.n34 585
R1440 B.n1377 B.n34 585
R1441 B.n1194 B.n33 585
R1442 B.n1378 B.n33 585
R1443 B.n1193 B.n1192 585
R1444 B.n1192 B.n29 585
R1445 B.n1191 B.n28 585
R1446 B.n1384 B.n28 585
R1447 B.n1190 B.n27 585
R1448 B.n1385 B.n27 585
R1449 B.n1189 B.n26 585
R1450 B.n1386 B.n26 585
R1451 B.n1188 B.n1187 585
R1452 B.n1187 B.n22 585
R1453 B.n1186 B.n21 585
R1454 B.n1392 B.n21 585
R1455 B.n1185 B.n20 585
R1456 B.n1393 B.n20 585
R1457 B.n1184 B.n19 585
R1458 B.n1394 B.n19 585
R1459 B.n1183 B.n1182 585
R1460 B.n1182 B.n18 585
R1461 B.n1181 B.n14 585
R1462 B.n1400 B.n14 585
R1463 B.n1180 B.n13 585
R1464 B.n1401 B.n13 585
R1465 B.n1179 B.n12 585
R1466 B.n1402 B.n12 585
R1467 B.n1178 B.n1177 585
R1468 B.n1177 B.n8 585
R1469 B.n1176 B.n7 585
R1470 B.n1408 B.n7 585
R1471 B.n1175 B.n6 585
R1472 B.n1409 B.n6 585
R1473 B.n1174 B.n5 585
R1474 B.n1410 B.n5 585
R1475 B.n1173 B.n1172 585
R1476 B.n1172 B.n4 585
R1477 B.n1171 B.n473 585
R1478 B.n1171 B.n1170 585
R1479 B.n1161 B.n474 585
R1480 B.n475 B.n474 585
R1481 B.n1163 B.n1162 585
R1482 B.n1164 B.n1163 585
R1483 B.n1160 B.n480 585
R1484 B.n480 B.n479 585
R1485 B.n1159 B.n1158 585
R1486 B.n1158 B.n1157 585
R1487 B.n482 B.n481 585
R1488 B.n1150 B.n482 585
R1489 B.n1149 B.n1148 585
R1490 B.n1151 B.n1149 585
R1491 B.n1147 B.n487 585
R1492 B.n487 B.n486 585
R1493 B.n1146 B.n1145 585
R1494 B.n1145 B.n1144 585
R1495 B.n489 B.n488 585
R1496 B.n490 B.n489 585
R1497 B.n1137 B.n1136 585
R1498 B.n1138 B.n1137 585
R1499 B.n1135 B.n495 585
R1500 B.n495 B.n494 585
R1501 B.n1134 B.n1133 585
R1502 B.n1133 B.n1132 585
R1503 B.n497 B.n496 585
R1504 B.n498 B.n497 585
R1505 B.n1125 B.n1124 585
R1506 B.n1126 B.n1125 585
R1507 B.n1123 B.n503 585
R1508 B.n503 B.n502 585
R1509 B.n1122 B.n1121 585
R1510 B.n1121 B.n1120 585
R1511 B.n505 B.n504 585
R1512 B.n506 B.n505 585
R1513 B.n1113 B.n1112 585
R1514 B.n1114 B.n1113 585
R1515 B.n1111 B.n511 585
R1516 B.n511 B.n510 585
R1517 B.n1110 B.n1109 585
R1518 B.n1109 B.n1108 585
R1519 B.n513 B.n512 585
R1520 B.n514 B.n513 585
R1521 B.n1101 B.n1100 585
R1522 B.n1102 B.n1101 585
R1523 B.n1099 B.n519 585
R1524 B.n519 B.n518 585
R1525 B.n1098 B.n1097 585
R1526 B.n1097 B.n1096 585
R1527 B.n521 B.n520 585
R1528 B.n522 B.n521 585
R1529 B.n1089 B.n1088 585
R1530 B.n1090 B.n1089 585
R1531 B.n1087 B.n527 585
R1532 B.n527 B.n526 585
R1533 B.n1086 B.n1085 585
R1534 B.n1085 B.n1084 585
R1535 B.n529 B.n528 585
R1536 B.n530 B.n529 585
R1537 B.n1077 B.n1076 585
R1538 B.n1078 B.n1077 585
R1539 B.n1075 B.n535 585
R1540 B.n535 B.n534 585
R1541 B.n1074 B.n1073 585
R1542 B.n1073 B.n1072 585
R1543 B.n537 B.n536 585
R1544 B.n538 B.n537 585
R1545 B.n1065 B.n1064 585
R1546 B.n1066 B.n1065 585
R1547 B.n1063 B.n543 585
R1548 B.n543 B.n542 585
R1549 B.n1062 B.n1061 585
R1550 B.n1061 B.n1060 585
R1551 B.n545 B.n544 585
R1552 B.n1053 B.n545 585
R1553 B.n1052 B.n1051 585
R1554 B.n1054 B.n1052 585
R1555 B.n1050 B.n550 585
R1556 B.n550 B.n549 585
R1557 B.n1049 B.n1048 585
R1558 B.n1048 B.n1047 585
R1559 B.n552 B.n551 585
R1560 B.n553 B.n552 585
R1561 B.n1040 B.n1039 585
R1562 B.n1041 B.n1040 585
R1563 B.n1038 B.n558 585
R1564 B.n558 B.n557 585
R1565 B.n1037 B.n1036 585
R1566 B.n1036 B.n1035 585
R1567 B.n560 B.n559 585
R1568 B.n561 B.n560 585
R1569 B.n1028 B.n1027 585
R1570 B.n1029 B.n1028 585
R1571 B.n1026 B.n565 585
R1572 B.n569 B.n565 585
R1573 B.n1025 B.n1024 585
R1574 B.n1024 B.n1023 585
R1575 B.n567 B.n566 585
R1576 B.n568 B.n567 585
R1577 B.n1016 B.n1015 585
R1578 B.n1017 B.n1016 585
R1579 B.n1014 B.n574 585
R1580 B.n574 B.n573 585
R1581 B.n1013 B.n1012 585
R1582 B.n1012 B.n1011 585
R1583 B.n576 B.n575 585
R1584 B.n577 B.n576 585
R1585 B.n1004 B.n1003 585
R1586 B.n1005 B.n1004 585
R1587 B.n1002 B.n582 585
R1588 B.n582 B.n581 585
R1589 B.n1001 B.n1000 585
R1590 B.n1000 B.n999 585
R1591 B.n584 B.n583 585
R1592 B.n585 B.n584 585
R1593 B.n992 B.n991 585
R1594 B.n993 B.n992 585
R1595 B.n990 B.n590 585
R1596 B.n590 B.n589 585
R1597 B.n989 B.n988 585
R1598 B.n988 B.n987 585
R1599 B.n592 B.n591 585
R1600 B.n980 B.n592 585
R1601 B.n979 B.n978 585
R1602 B.n981 B.n979 585
R1603 B.n977 B.n597 585
R1604 B.n597 B.n596 585
R1605 B.n976 B.n975 585
R1606 B.n975 B.n974 585
R1607 B.n599 B.n598 585
R1608 B.n600 B.n599 585
R1609 B.n967 B.n966 585
R1610 B.n968 B.n967 585
R1611 B.n965 B.n605 585
R1612 B.n605 B.n604 585
R1613 B.n964 B.n963 585
R1614 B.n963 B.n962 585
R1615 B.n607 B.n606 585
R1616 B.n608 B.n607 585
R1617 B.n958 B.n957 585
R1618 B.n611 B.n610 585
R1619 B.n954 B.n953 585
R1620 B.n955 B.n954 585
R1621 B.n952 B.n679 585
R1622 B.n951 B.n950 585
R1623 B.n949 B.n948 585
R1624 B.n947 B.n946 585
R1625 B.n945 B.n944 585
R1626 B.n943 B.n942 585
R1627 B.n941 B.n940 585
R1628 B.n939 B.n938 585
R1629 B.n937 B.n936 585
R1630 B.n935 B.n934 585
R1631 B.n933 B.n932 585
R1632 B.n931 B.n930 585
R1633 B.n929 B.n928 585
R1634 B.n927 B.n926 585
R1635 B.n925 B.n924 585
R1636 B.n923 B.n922 585
R1637 B.n921 B.n920 585
R1638 B.n919 B.n918 585
R1639 B.n917 B.n916 585
R1640 B.n915 B.n914 585
R1641 B.n913 B.n912 585
R1642 B.n911 B.n910 585
R1643 B.n909 B.n908 585
R1644 B.n907 B.n906 585
R1645 B.n905 B.n904 585
R1646 B.n903 B.n902 585
R1647 B.n901 B.n900 585
R1648 B.n899 B.n898 585
R1649 B.n897 B.n896 585
R1650 B.n895 B.n894 585
R1651 B.n893 B.n892 585
R1652 B.n891 B.n890 585
R1653 B.n889 B.n888 585
R1654 B.n887 B.n886 585
R1655 B.n885 B.n884 585
R1656 B.n883 B.n882 585
R1657 B.n881 B.n880 585
R1658 B.n879 B.n878 585
R1659 B.n877 B.n876 585
R1660 B.n875 B.n874 585
R1661 B.n873 B.n872 585
R1662 B.n871 B.n870 585
R1663 B.n869 B.n868 585
R1664 B.n867 B.n866 585
R1665 B.n865 B.n864 585
R1666 B.n863 B.n862 585
R1667 B.n861 B.n860 585
R1668 B.n859 B.n858 585
R1669 B.n857 B.n856 585
R1670 B.n855 B.n854 585
R1671 B.n853 B.n852 585
R1672 B.n851 B.n850 585
R1673 B.n849 B.n848 585
R1674 B.n847 B.n846 585
R1675 B.n845 B.n844 585
R1676 B.n843 B.n842 585
R1677 B.n841 B.n840 585
R1678 B.n839 B.n838 585
R1679 B.n837 B.n836 585
R1680 B.n835 B.n834 585
R1681 B.n833 B.n832 585
R1682 B.n830 B.n829 585
R1683 B.n828 B.n827 585
R1684 B.n826 B.n825 585
R1685 B.n824 B.n823 585
R1686 B.n822 B.n821 585
R1687 B.n820 B.n819 585
R1688 B.n818 B.n817 585
R1689 B.n816 B.n815 585
R1690 B.n814 B.n813 585
R1691 B.n812 B.n811 585
R1692 B.n810 B.n809 585
R1693 B.n808 B.n807 585
R1694 B.n806 B.n805 585
R1695 B.n804 B.n803 585
R1696 B.n802 B.n801 585
R1697 B.n800 B.n799 585
R1698 B.n798 B.n797 585
R1699 B.n796 B.n795 585
R1700 B.n794 B.n793 585
R1701 B.n792 B.n791 585
R1702 B.n790 B.n789 585
R1703 B.n788 B.n787 585
R1704 B.n786 B.n785 585
R1705 B.n784 B.n783 585
R1706 B.n782 B.n781 585
R1707 B.n780 B.n779 585
R1708 B.n778 B.n777 585
R1709 B.n776 B.n775 585
R1710 B.n774 B.n773 585
R1711 B.n772 B.n771 585
R1712 B.n770 B.n769 585
R1713 B.n768 B.n767 585
R1714 B.n766 B.n765 585
R1715 B.n764 B.n763 585
R1716 B.n762 B.n761 585
R1717 B.n760 B.n759 585
R1718 B.n758 B.n757 585
R1719 B.n756 B.n755 585
R1720 B.n754 B.n753 585
R1721 B.n752 B.n751 585
R1722 B.n750 B.n749 585
R1723 B.n748 B.n747 585
R1724 B.n746 B.n745 585
R1725 B.n744 B.n743 585
R1726 B.n742 B.n741 585
R1727 B.n740 B.n739 585
R1728 B.n738 B.n737 585
R1729 B.n736 B.n735 585
R1730 B.n734 B.n733 585
R1731 B.n732 B.n731 585
R1732 B.n730 B.n729 585
R1733 B.n728 B.n727 585
R1734 B.n726 B.n725 585
R1735 B.n724 B.n723 585
R1736 B.n722 B.n721 585
R1737 B.n720 B.n719 585
R1738 B.n718 B.n717 585
R1739 B.n716 B.n715 585
R1740 B.n714 B.n713 585
R1741 B.n712 B.n711 585
R1742 B.n710 B.n709 585
R1743 B.n708 B.n707 585
R1744 B.n706 B.n705 585
R1745 B.n704 B.n703 585
R1746 B.n702 B.n701 585
R1747 B.n700 B.n699 585
R1748 B.n698 B.n697 585
R1749 B.n696 B.n695 585
R1750 B.n694 B.n693 585
R1751 B.n692 B.n691 585
R1752 B.n690 B.n689 585
R1753 B.n688 B.n687 585
R1754 B.n686 B.n685 585
R1755 B.n959 B.n609 585
R1756 B.n609 B.n608 585
R1757 B.n961 B.n960 585
R1758 B.n962 B.n961 585
R1759 B.n603 B.n602 585
R1760 B.n604 B.n603 585
R1761 B.n970 B.n969 585
R1762 B.n969 B.n968 585
R1763 B.n971 B.n601 585
R1764 B.n601 B.n600 585
R1765 B.n973 B.n972 585
R1766 B.n974 B.n973 585
R1767 B.n595 B.n594 585
R1768 B.n596 B.n595 585
R1769 B.n983 B.n982 585
R1770 B.n982 B.n981 585
R1771 B.n984 B.n593 585
R1772 B.n980 B.n593 585
R1773 B.n986 B.n985 585
R1774 B.n987 B.n986 585
R1775 B.n588 B.n587 585
R1776 B.n589 B.n588 585
R1777 B.n995 B.n994 585
R1778 B.n994 B.n993 585
R1779 B.n996 B.n586 585
R1780 B.n586 B.n585 585
R1781 B.n998 B.n997 585
R1782 B.n999 B.n998 585
R1783 B.n580 B.n579 585
R1784 B.n581 B.n580 585
R1785 B.n1007 B.n1006 585
R1786 B.n1006 B.n1005 585
R1787 B.n1008 B.n578 585
R1788 B.n578 B.n577 585
R1789 B.n1010 B.n1009 585
R1790 B.n1011 B.n1010 585
R1791 B.n572 B.n571 585
R1792 B.n573 B.n572 585
R1793 B.n1019 B.n1018 585
R1794 B.n1018 B.n1017 585
R1795 B.n1020 B.n570 585
R1796 B.n570 B.n568 585
R1797 B.n1022 B.n1021 585
R1798 B.n1023 B.n1022 585
R1799 B.n564 B.n563 585
R1800 B.n569 B.n564 585
R1801 B.n1031 B.n1030 585
R1802 B.n1030 B.n1029 585
R1803 B.n1032 B.n562 585
R1804 B.n562 B.n561 585
R1805 B.n1034 B.n1033 585
R1806 B.n1035 B.n1034 585
R1807 B.n556 B.n555 585
R1808 B.n557 B.n556 585
R1809 B.n1043 B.n1042 585
R1810 B.n1042 B.n1041 585
R1811 B.n1044 B.n554 585
R1812 B.n554 B.n553 585
R1813 B.n1046 B.n1045 585
R1814 B.n1047 B.n1046 585
R1815 B.n548 B.n547 585
R1816 B.n549 B.n548 585
R1817 B.n1056 B.n1055 585
R1818 B.n1055 B.n1054 585
R1819 B.n1057 B.n546 585
R1820 B.n1053 B.n546 585
R1821 B.n1059 B.n1058 585
R1822 B.n1060 B.n1059 585
R1823 B.n541 B.n540 585
R1824 B.n542 B.n541 585
R1825 B.n1068 B.n1067 585
R1826 B.n1067 B.n1066 585
R1827 B.n1069 B.n539 585
R1828 B.n539 B.n538 585
R1829 B.n1071 B.n1070 585
R1830 B.n1072 B.n1071 585
R1831 B.n533 B.n532 585
R1832 B.n534 B.n533 585
R1833 B.n1080 B.n1079 585
R1834 B.n1079 B.n1078 585
R1835 B.n1081 B.n531 585
R1836 B.n531 B.n530 585
R1837 B.n1083 B.n1082 585
R1838 B.n1084 B.n1083 585
R1839 B.n525 B.n524 585
R1840 B.n526 B.n525 585
R1841 B.n1092 B.n1091 585
R1842 B.n1091 B.n1090 585
R1843 B.n1093 B.n523 585
R1844 B.n523 B.n522 585
R1845 B.n1095 B.n1094 585
R1846 B.n1096 B.n1095 585
R1847 B.n517 B.n516 585
R1848 B.n518 B.n517 585
R1849 B.n1104 B.n1103 585
R1850 B.n1103 B.n1102 585
R1851 B.n1105 B.n515 585
R1852 B.n515 B.n514 585
R1853 B.n1107 B.n1106 585
R1854 B.n1108 B.n1107 585
R1855 B.n509 B.n508 585
R1856 B.n510 B.n509 585
R1857 B.n1116 B.n1115 585
R1858 B.n1115 B.n1114 585
R1859 B.n1117 B.n507 585
R1860 B.n507 B.n506 585
R1861 B.n1119 B.n1118 585
R1862 B.n1120 B.n1119 585
R1863 B.n501 B.n500 585
R1864 B.n502 B.n501 585
R1865 B.n1128 B.n1127 585
R1866 B.n1127 B.n1126 585
R1867 B.n1129 B.n499 585
R1868 B.n499 B.n498 585
R1869 B.n1131 B.n1130 585
R1870 B.n1132 B.n1131 585
R1871 B.n493 B.n492 585
R1872 B.n494 B.n493 585
R1873 B.n1140 B.n1139 585
R1874 B.n1139 B.n1138 585
R1875 B.n1141 B.n491 585
R1876 B.n491 B.n490 585
R1877 B.n1143 B.n1142 585
R1878 B.n1144 B.n1143 585
R1879 B.n485 B.n484 585
R1880 B.n486 B.n485 585
R1881 B.n1153 B.n1152 585
R1882 B.n1152 B.n1151 585
R1883 B.n1154 B.n483 585
R1884 B.n1150 B.n483 585
R1885 B.n1156 B.n1155 585
R1886 B.n1157 B.n1156 585
R1887 B.n478 B.n477 585
R1888 B.n479 B.n478 585
R1889 B.n1166 B.n1165 585
R1890 B.n1165 B.n1164 585
R1891 B.n1167 B.n476 585
R1892 B.n476 B.n475 585
R1893 B.n1169 B.n1168 585
R1894 B.n1170 B.n1169 585
R1895 B.n2 B.n0 585
R1896 B.n4 B.n2 585
R1897 B.n3 B.n1 585
R1898 B.n1409 B.n3 585
R1899 B.n1407 B.n1406 585
R1900 B.n1408 B.n1407 585
R1901 B.n1405 B.n9 585
R1902 B.n9 B.n8 585
R1903 B.n1404 B.n1403 585
R1904 B.n1403 B.n1402 585
R1905 B.n11 B.n10 585
R1906 B.n1401 B.n11 585
R1907 B.n1399 B.n1398 585
R1908 B.n1400 B.n1399 585
R1909 B.n1397 B.n15 585
R1910 B.n18 B.n15 585
R1911 B.n1396 B.n1395 585
R1912 B.n1395 B.n1394 585
R1913 B.n17 B.n16 585
R1914 B.n1393 B.n17 585
R1915 B.n1391 B.n1390 585
R1916 B.n1392 B.n1391 585
R1917 B.n1389 B.n23 585
R1918 B.n23 B.n22 585
R1919 B.n1388 B.n1387 585
R1920 B.n1387 B.n1386 585
R1921 B.n25 B.n24 585
R1922 B.n1385 B.n25 585
R1923 B.n1383 B.n1382 585
R1924 B.n1384 B.n1383 585
R1925 B.n1381 B.n30 585
R1926 B.n30 B.n29 585
R1927 B.n1380 B.n1379 585
R1928 B.n1379 B.n1378 585
R1929 B.n32 B.n31 585
R1930 B.n1377 B.n32 585
R1931 B.n1375 B.n1374 585
R1932 B.n1376 B.n1375 585
R1933 B.n1373 B.n37 585
R1934 B.n37 B.n36 585
R1935 B.n1372 B.n1371 585
R1936 B.n1371 B.n1370 585
R1937 B.n39 B.n38 585
R1938 B.n1369 B.n39 585
R1939 B.n1367 B.n1366 585
R1940 B.n1368 B.n1367 585
R1941 B.n1365 B.n44 585
R1942 B.n44 B.n43 585
R1943 B.n1364 B.n1363 585
R1944 B.n1363 B.n1362 585
R1945 B.n46 B.n45 585
R1946 B.n1361 B.n46 585
R1947 B.n1359 B.n1358 585
R1948 B.n1360 B.n1359 585
R1949 B.n1357 B.n51 585
R1950 B.n51 B.n50 585
R1951 B.n1356 B.n1355 585
R1952 B.n1355 B.n1354 585
R1953 B.n53 B.n52 585
R1954 B.n1353 B.n53 585
R1955 B.n1351 B.n1350 585
R1956 B.n1352 B.n1351 585
R1957 B.n1349 B.n58 585
R1958 B.n58 B.n57 585
R1959 B.n1348 B.n1347 585
R1960 B.n1347 B.n1346 585
R1961 B.n60 B.n59 585
R1962 B.n1345 B.n60 585
R1963 B.n1343 B.n1342 585
R1964 B.n1344 B.n1343 585
R1965 B.n1341 B.n65 585
R1966 B.n65 B.n64 585
R1967 B.n1340 B.n1339 585
R1968 B.n1339 B.n1338 585
R1969 B.n67 B.n66 585
R1970 B.n1337 B.n67 585
R1971 B.n1335 B.n1334 585
R1972 B.n1336 B.n1335 585
R1973 B.n1333 B.n71 585
R1974 B.n74 B.n71 585
R1975 B.n1332 B.n1331 585
R1976 B.n1331 B.n1330 585
R1977 B.n73 B.n72 585
R1978 B.n1329 B.n73 585
R1979 B.n1327 B.n1326 585
R1980 B.n1328 B.n1327 585
R1981 B.n1325 B.n79 585
R1982 B.n79 B.n78 585
R1983 B.n1324 B.n1323 585
R1984 B.n1323 B.n1322 585
R1985 B.n81 B.n80 585
R1986 B.n1321 B.n81 585
R1987 B.n1319 B.n1318 585
R1988 B.n1320 B.n1319 585
R1989 B.n1317 B.n86 585
R1990 B.n86 B.n85 585
R1991 B.n1316 B.n1315 585
R1992 B.n1315 B.n1314 585
R1993 B.n88 B.n87 585
R1994 B.n1313 B.n88 585
R1995 B.n1311 B.n1310 585
R1996 B.n1312 B.n1311 585
R1997 B.n1309 B.n93 585
R1998 B.n93 B.n92 585
R1999 B.n1308 B.n1307 585
R2000 B.n1307 B.n1306 585
R2001 B.n95 B.n94 585
R2002 B.n1305 B.n95 585
R2003 B.n1303 B.n1302 585
R2004 B.n1304 B.n1303 585
R2005 B.n1301 B.n100 585
R2006 B.n100 B.n99 585
R2007 B.n1300 B.n1299 585
R2008 B.n1299 B.n1298 585
R2009 B.n102 B.n101 585
R2010 B.n1297 B.n102 585
R2011 B.n1295 B.n1294 585
R2012 B.n1296 B.n1295 585
R2013 B.n1293 B.n107 585
R2014 B.n107 B.n106 585
R2015 B.n1292 B.n1291 585
R2016 B.n1291 B.n1290 585
R2017 B.n109 B.n108 585
R2018 B.n1289 B.n109 585
R2019 B.n1287 B.n1286 585
R2020 B.n1288 B.n1287 585
R2021 B.n1285 B.n113 585
R2022 B.n116 B.n113 585
R2023 B.n1284 B.n1283 585
R2024 B.n1283 B.n1282 585
R2025 B.n115 B.n114 585
R2026 B.n1281 B.n115 585
R2027 B.n1279 B.n1278 585
R2028 B.n1280 B.n1279 585
R2029 B.n1277 B.n121 585
R2030 B.n121 B.n120 585
R2031 B.n1276 B.n1275 585
R2032 B.n1275 B.n1274 585
R2033 B.n123 B.n122 585
R2034 B.n1273 B.n123 585
R2035 B.n1271 B.n1270 585
R2036 B.n1272 B.n1271 585
R2037 B.n1269 B.n128 585
R2038 B.n128 B.n127 585
R2039 B.n1412 B.n1411 585
R2040 B.n1411 B.n1410 585
R2041 B.n957 B.n609 521.33
R2042 B.n1267 B.n128 521.33
R2043 B.n685 B.n607 521.33
R2044 B.n1264 B.n199 521.33
R2045 B.n682 B.t23 481.827
R2046 B.n200 B.t19 481.827
R2047 B.n680 B.t13 481.827
R2048 B.n202 B.t16 481.827
R2049 B.n683 B.t22 412.784
R2050 B.n201 B.t20 412.784
R2051 B.n681 B.t12 412.784
R2052 B.n203 B.t17 412.784
R2053 B.n682 B.t21 354.926
R2054 B.n680 B.t10 354.926
R2055 B.n202 B.t14 354.926
R2056 B.n200 B.t18 354.926
R2057 B.n1265 B.n197 256.663
R2058 B.n1265 B.n196 256.663
R2059 B.n1265 B.n195 256.663
R2060 B.n1265 B.n194 256.663
R2061 B.n1265 B.n193 256.663
R2062 B.n1265 B.n192 256.663
R2063 B.n1265 B.n191 256.663
R2064 B.n1265 B.n190 256.663
R2065 B.n1265 B.n189 256.663
R2066 B.n1265 B.n188 256.663
R2067 B.n1265 B.n187 256.663
R2068 B.n1265 B.n186 256.663
R2069 B.n1265 B.n185 256.663
R2070 B.n1265 B.n184 256.663
R2071 B.n1265 B.n183 256.663
R2072 B.n1265 B.n182 256.663
R2073 B.n1265 B.n181 256.663
R2074 B.n1265 B.n180 256.663
R2075 B.n1265 B.n179 256.663
R2076 B.n1265 B.n178 256.663
R2077 B.n1265 B.n177 256.663
R2078 B.n1265 B.n176 256.663
R2079 B.n1265 B.n175 256.663
R2080 B.n1265 B.n174 256.663
R2081 B.n1265 B.n173 256.663
R2082 B.n1265 B.n172 256.663
R2083 B.n1265 B.n171 256.663
R2084 B.n1265 B.n170 256.663
R2085 B.n1265 B.n169 256.663
R2086 B.n1265 B.n168 256.663
R2087 B.n1265 B.n167 256.663
R2088 B.n1265 B.n166 256.663
R2089 B.n1265 B.n165 256.663
R2090 B.n1265 B.n164 256.663
R2091 B.n1265 B.n163 256.663
R2092 B.n1265 B.n162 256.663
R2093 B.n1265 B.n161 256.663
R2094 B.n1265 B.n160 256.663
R2095 B.n1265 B.n159 256.663
R2096 B.n1265 B.n158 256.663
R2097 B.n1265 B.n157 256.663
R2098 B.n1265 B.n156 256.663
R2099 B.n1265 B.n155 256.663
R2100 B.n1265 B.n154 256.663
R2101 B.n1265 B.n153 256.663
R2102 B.n1265 B.n152 256.663
R2103 B.n1265 B.n151 256.663
R2104 B.n1265 B.n150 256.663
R2105 B.n1265 B.n149 256.663
R2106 B.n1265 B.n148 256.663
R2107 B.n1265 B.n147 256.663
R2108 B.n1265 B.n146 256.663
R2109 B.n1265 B.n145 256.663
R2110 B.n1265 B.n144 256.663
R2111 B.n1265 B.n143 256.663
R2112 B.n1265 B.n142 256.663
R2113 B.n1265 B.n141 256.663
R2114 B.n1265 B.n140 256.663
R2115 B.n1265 B.n139 256.663
R2116 B.n1265 B.n138 256.663
R2117 B.n1265 B.n137 256.663
R2118 B.n1265 B.n136 256.663
R2119 B.n1265 B.n135 256.663
R2120 B.n1265 B.n134 256.663
R2121 B.n1265 B.n133 256.663
R2122 B.n1265 B.n132 256.663
R2123 B.n1265 B.n131 256.663
R2124 B.n1266 B.n1265 256.663
R2125 B.n956 B.n955 256.663
R2126 B.n955 B.n612 256.663
R2127 B.n955 B.n613 256.663
R2128 B.n955 B.n614 256.663
R2129 B.n955 B.n615 256.663
R2130 B.n955 B.n616 256.663
R2131 B.n955 B.n617 256.663
R2132 B.n955 B.n618 256.663
R2133 B.n955 B.n619 256.663
R2134 B.n955 B.n620 256.663
R2135 B.n955 B.n621 256.663
R2136 B.n955 B.n622 256.663
R2137 B.n955 B.n623 256.663
R2138 B.n955 B.n624 256.663
R2139 B.n955 B.n625 256.663
R2140 B.n955 B.n626 256.663
R2141 B.n955 B.n627 256.663
R2142 B.n955 B.n628 256.663
R2143 B.n955 B.n629 256.663
R2144 B.n955 B.n630 256.663
R2145 B.n955 B.n631 256.663
R2146 B.n955 B.n632 256.663
R2147 B.n955 B.n633 256.663
R2148 B.n955 B.n634 256.663
R2149 B.n955 B.n635 256.663
R2150 B.n955 B.n636 256.663
R2151 B.n955 B.n637 256.663
R2152 B.n955 B.n638 256.663
R2153 B.n955 B.n639 256.663
R2154 B.n955 B.n640 256.663
R2155 B.n955 B.n641 256.663
R2156 B.n955 B.n642 256.663
R2157 B.n955 B.n643 256.663
R2158 B.n955 B.n644 256.663
R2159 B.n955 B.n645 256.663
R2160 B.n955 B.n646 256.663
R2161 B.n955 B.n647 256.663
R2162 B.n955 B.n648 256.663
R2163 B.n955 B.n649 256.663
R2164 B.n955 B.n650 256.663
R2165 B.n955 B.n651 256.663
R2166 B.n955 B.n652 256.663
R2167 B.n955 B.n653 256.663
R2168 B.n955 B.n654 256.663
R2169 B.n955 B.n655 256.663
R2170 B.n955 B.n656 256.663
R2171 B.n955 B.n657 256.663
R2172 B.n955 B.n658 256.663
R2173 B.n955 B.n659 256.663
R2174 B.n955 B.n660 256.663
R2175 B.n955 B.n661 256.663
R2176 B.n955 B.n662 256.663
R2177 B.n955 B.n663 256.663
R2178 B.n955 B.n664 256.663
R2179 B.n955 B.n665 256.663
R2180 B.n955 B.n666 256.663
R2181 B.n955 B.n667 256.663
R2182 B.n955 B.n668 256.663
R2183 B.n955 B.n669 256.663
R2184 B.n955 B.n670 256.663
R2185 B.n955 B.n671 256.663
R2186 B.n955 B.n672 256.663
R2187 B.n955 B.n673 256.663
R2188 B.n955 B.n674 256.663
R2189 B.n955 B.n675 256.663
R2190 B.n955 B.n676 256.663
R2191 B.n955 B.n677 256.663
R2192 B.n955 B.n678 256.663
R2193 B.n961 B.n609 163.367
R2194 B.n961 B.n603 163.367
R2195 B.n969 B.n603 163.367
R2196 B.n969 B.n601 163.367
R2197 B.n973 B.n601 163.367
R2198 B.n973 B.n595 163.367
R2199 B.n982 B.n595 163.367
R2200 B.n982 B.n593 163.367
R2201 B.n986 B.n593 163.367
R2202 B.n986 B.n588 163.367
R2203 B.n994 B.n588 163.367
R2204 B.n994 B.n586 163.367
R2205 B.n998 B.n586 163.367
R2206 B.n998 B.n580 163.367
R2207 B.n1006 B.n580 163.367
R2208 B.n1006 B.n578 163.367
R2209 B.n1010 B.n578 163.367
R2210 B.n1010 B.n572 163.367
R2211 B.n1018 B.n572 163.367
R2212 B.n1018 B.n570 163.367
R2213 B.n1022 B.n570 163.367
R2214 B.n1022 B.n564 163.367
R2215 B.n1030 B.n564 163.367
R2216 B.n1030 B.n562 163.367
R2217 B.n1034 B.n562 163.367
R2218 B.n1034 B.n556 163.367
R2219 B.n1042 B.n556 163.367
R2220 B.n1042 B.n554 163.367
R2221 B.n1046 B.n554 163.367
R2222 B.n1046 B.n548 163.367
R2223 B.n1055 B.n548 163.367
R2224 B.n1055 B.n546 163.367
R2225 B.n1059 B.n546 163.367
R2226 B.n1059 B.n541 163.367
R2227 B.n1067 B.n541 163.367
R2228 B.n1067 B.n539 163.367
R2229 B.n1071 B.n539 163.367
R2230 B.n1071 B.n533 163.367
R2231 B.n1079 B.n533 163.367
R2232 B.n1079 B.n531 163.367
R2233 B.n1083 B.n531 163.367
R2234 B.n1083 B.n525 163.367
R2235 B.n1091 B.n525 163.367
R2236 B.n1091 B.n523 163.367
R2237 B.n1095 B.n523 163.367
R2238 B.n1095 B.n517 163.367
R2239 B.n1103 B.n517 163.367
R2240 B.n1103 B.n515 163.367
R2241 B.n1107 B.n515 163.367
R2242 B.n1107 B.n509 163.367
R2243 B.n1115 B.n509 163.367
R2244 B.n1115 B.n507 163.367
R2245 B.n1119 B.n507 163.367
R2246 B.n1119 B.n501 163.367
R2247 B.n1127 B.n501 163.367
R2248 B.n1127 B.n499 163.367
R2249 B.n1131 B.n499 163.367
R2250 B.n1131 B.n493 163.367
R2251 B.n1139 B.n493 163.367
R2252 B.n1139 B.n491 163.367
R2253 B.n1143 B.n491 163.367
R2254 B.n1143 B.n485 163.367
R2255 B.n1152 B.n485 163.367
R2256 B.n1152 B.n483 163.367
R2257 B.n1156 B.n483 163.367
R2258 B.n1156 B.n478 163.367
R2259 B.n1165 B.n478 163.367
R2260 B.n1165 B.n476 163.367
R2261 B.n1169 B.n476 163.367
R2262 B.n1169 B.n2 163.367
R2263 B.n1411 B.n2 163.367
R2264 B.n1411 B.n3 163.367
R2265 B.n1407 B.n3 163.367
R2266 B.n1407 B.n9 163.367
R2267 B.n1403 B.n9 163.367
R2268 B.n1403 B.n11 163.367
R2269 B.n1399 B.n11 163.367
R2270 B.n1399 B.n15 163.367
R2271 B.n1395 B.n15 163.367
R2272 B.n1395 B.n17 163.367
R2273 B.n1391 B.n17 163.367
R2274 B.n1391 B.n23 163.367
R2275 B.n1387 B.n23 163.367
R2276 B.n1387 B.n25 163.367
R2277 B.n1383 B.n25 163.367
R2278 B.n1383 B.n30 163.367
R2279 B.n1379 B.n30 163.367
R2280 B.n1379 B.n32 163.367
R2281 B.n1375 B.n32 163.367
R2282 B.n1375 B.n37 163.367
R2283 B.n1371 B.n37 163.367
R2284 B.n1371 B.n39 163.367
R2285 B.n1367 B.n39 163.367
R2286 B.n1367 B.n44 163.367
R2287 B.n1363 B.n44 163.367
R2288 B.n1363 B.n46 163.367
R2289 B.n1359 B.n46 163.367
R2290 B.n1359 B.n51 163.367
R2291 B.n1355 B.n51 163.367
R2292 B.n1355 B.n53 163.367
R2293 B.n1351 B.n53 163.367
R2294 B.n1351 B.n58 163.367
R2295 B.n1347 B.n58 163.367
R2296 B.n1347 B.n60 163.367
R2297 B.n1343 B.n60 163.367
R2298 B.n1343 B.n65 163.367
R2299 B.n1339 B.n65 163.367
R2300 B.n1339 B.n67 163.367
R2301 B.n1335 B.n67 163.367
R2302 B.n1335 B.n71 163.367
R2303 B.n1331 B.n71 163.367
R2304 B.n1331 B.n73 163.367
R2305 B.n1327 B.n73 163.367
R2306 B.n1327 B.n79 163.367
R2307 B.n1323 B.n79 163.367
R2308 B.n1323 B.n81 163.367
R2309 B.n1319 B.n81 163.367
R2310 B.n1319 B.n86 163.367
R2311 B.n1315 B.n86 163.367
R2312 B.n1315 B.n88 163.367
R2313 B.n1311 B.n88 163.367
R2314 B.n1311 B.n93 163.367
R2315 B.n1307 B.n93 163.367
R2316 B.n1307 B.n95 163.367
R2317 B.n1303 B.n95 163.367
R2318 B.n1303 B.n100 163.367
R2319 B.n1299 B.n100 163.367
R2320 B.n1299 B.n102 163.367
R2321 B.n1295 B.n102 163.367
R2322 B.n1295 B.n107 163.367
R2323 B.n1291 B.n107 163.367
R2324 B.n1291 B.n109 163.367
R2325 B.n1287 B.n109 163.367
R2326 B.n1287 B.n113 163.367
R2327 B.n1283 B.n113 163.367
R2328 B.n1283 B.n115 163.367
R2329 B.n1279 B.n115 163.367
R2330 B.n1279 B.n121 163.367
R2331 B.n1275 B.n121 163.367
R2332 B.n1275 B.n123 163.367
R2333 B.n1271 B.n123 163.367
R2334 B.n1271 B.n128 163.367
R2335 B.n954 B.n611 163.367
R2336 B.n954 B.n679 163.367
R2337 B.n950 B.n949 163.367
R2338 B.n946 B.n945 163.367
R2339 B.n942 B.n941 163.367
R2340 B.n938 B.n937 163.367
R2341 B.n934 B.n933 163.367
R2342 B.n930 B.n929 163.367
R2343 B.n926 B.n925 163.367
R2344 B.n922 B.n921 163.367
R2345 B.n918 B.n917 163.367
R2346 B.n914 B.n913 163.367
R2347 B.n910 B.n909 163.367
R2348 B.n906 B.n905 163.367
R2349 B.n902 B.n901 163.367
R2350 B.n898 B.n897 163.367
R2351 B.n894 B.n893 163.367
R2352 B.n890 B.n889 163.367
R2353 B.n886 B.n885 163.367
R2354 B.n882 B.n881 163.367
R2355 B.n878 B.n877 163.367
R2356 B.n874 B.n873 163.367
R2357 B.n870 B.n869 163.367
R2358 B.n866 B.n865 163.367
R2359 B.n862 B.n861 163.367
R2360 B.n858 B.n857 163.367
R2361 B.n854 B.n853 163.367
R2362 B.n850 B.n849 163.367
R2363 B.n846 B.n845 163.367
R2364 B.n842 B.n841 163.367
R2365 B.n838 B.n837 163.367
R2366 B.n834 B.n833 163.367
R2367 B.n829 B.n828 163.367
R2368 B.n825 B.n824 163.367
R2369 B.n821 B.n820 163.367
R2370 B.n817 B.n816 163.367
R2371 B.n813 B.n812 163.367
R2372 B.n809 B.n808 163.367
R2373 B.n805 B.n804 163.367
R2374 B.n801 B.n800 163.367
R2375 B.n797 B.n796 163.367
R2376 B.n793 B.n792 163.367
R2377 B.n789 B.n788 163.367
R2378 B.n785 B.n784 163.367
R2379 B.n781 B.n780 163.367
R2380 B.n777 B.n776 163.367
R2381 B.n773 B.n772 163.367
R2382 B.n769 B.n768 163.367
R2383 B.n765 B.n764 163.367
R2384 B.n761 B.n760 163.367
R2385 B.n757 B.n756 163.367
R2386 B.n753 B.n752 163.367
R2387 B.n749 B.n748 163.367
R2388 B.n745 B.n744 163.367
R2389 B.n741 B.n740 163.367
R2390 B.n737 B.n736 163.367
R2391 B.n733 B.n732 163.367
R2392 B.n729 B.n728 163.367
R2393 B.n725 B.n724 163.367
R2394 B.n721 B.n720 163.367
R2395 B.n717 B.n716 163.367
R2396 B.n713 B.n712 163.367
R2397 B.n709 B.n708 163.367
R2398 B.n705 B.n704 163.367
R2399 B.n701 B.n700 163.367
R2400 B.n697 B.n696 163.367
R2401 B.n693 B.n692 163.367
R2402 B.n689 B.n688 163.367
R2403 B.n963 B.n607 163.367
R2404 B.n963 B.n605 163.367
R2405 B.n967 B.n605 163.367
R2406 B.n967 B.n599 163.367
R2407 B.n975 B.n599 163.367
R2408 B.n975 B.n597 163.367
R2409 B.n979 B.n597 163.367
R2410 B.n979 B.n592 163.367
R2411 B.n988 B.n592 163.367
R2412 B.n988 B.n590 163.367
R2413 B.n992 B.n590 163.367
R2414 B.n992 B.n584 163.367
R2415 B.n1000 B.n584 163.367
R2416 B.n1000 B.n582 163.367
R2417 B.n1004 B.n582 163.367
R2418 B.n1004 B.n576 163.367
R2419 B.n1012 B.n576 163.367
R2420 B.n1012 B.n574 163.367
R2421 B.n1016 B.n574 163.367
R2422 B.n1016 B.n567 163.367
R2423 B.n1024 B.n567 163.367
R2424 B.n1024 B.n565 163.367
R2425 B.n1028 B.n565 163.367
R2426 B.n1028 B.n560 163.367
R2427 B.n1036 B.n560 163.367
R2428 B.n1036 B.n558 163.367
R2429 B.n1040 B.n558 163.367
R2430 B.n1040 B.n552 163.367
R2431 B.n1048 B.n552 163.367
R2432 B.n1048 B.n550 163.367
R2433 B.n1052 B.n550 163.367
R2434 B.n1052 B.n545 163.367
R2435 B.n1061 B.n545 163.367
R2436 B.n1061 B.n543 163.367
R2437 B.n1065 B.n543 163.367
R2438 B.n1065 B.n537 163.367
R2439 B.n1073 B.n537 163.367
R2440 B.n1073 B.n535 163.367
R2441 B.n1077 B.n535 163.367
R2442 B.n1077 B.n529 163.367
R2443 B.n1085 B.n529 163.367
R2444 B.n1085 B.n527 163.367
R2445 B.n1089 B.n527 163.367
R2446 B.n1089 B.n521 163.367
R2447 B.n1097 B.n521 163.367
R2448 B.n1097 B.n519 163.367
R2449 B.n1101 B.n519 163.367
R2450 B.n1101 B.n513 163.367
R2451 B.n1109 B.n513 163.367
R2452 B.n1109 B.n511 163.367
R2453 B.n1113 B.n511 163.367
R2454 B.n1113 B.n505 163.367
R2455 B.n1121 B.n505 163.367
R2456 B.n1121 B.n503 163.367
R2457 B.n1125 B.n503 163.367
R2458 B.n1125 B.n497 163.367
R2459 B.n1133 B.n497 163.367
R2460 B.n1133 B.n495 163.367
R2461 B.n1137 B.n495 163.367
R2462 B.n1137 B.n489 163.367
R2463 B.n1145 B.n489 163.367
R2464 B.n1145 B.n487 163.367
R2465 B.n1149 B.n487 163.367
R2466 B.n1149 B.n482 163.367
R2467 B.n1158 B.n482 163.367
R2468 B.n1158 B.n480 163.367
R2469 B.n1163 B.n480 163.367
R2470 B.n1163 B.n474 163.367
R2471 B.n1171 B.n474 163.367
R2472 B.n1172 B.n1171 163.367
R2473 B.n1172 B.n5 163.367
R2474 B.n6 B.n5 163.367
R2475 B.n7 B.n6 163.367
R2476 B.n1177 B.n7 163.367
R2477 B.n1177 B.n12 163.367
R2478 B.n13 B.n12 163.367
R2479 B.n14 B.n13 163.367
R2480 B.n1182 B.n14 163.367
R2481 B.n1182 B.n19 163.367
R2482 B.n20 B.n19 163.367
R2483 B.n21 B.n20 163.367
R2484 B.n1187 B.n21 163.367
R2485 B.n1187 B.n26 163.367
R2486 B.n27 B.n26 163.367
R2487 B.n28 B.n27 163.367
R2488 B.n1192 B.n28 163.367
R2489 B.n1192 B.n33 163.367
R2490 B.n34 B.n33 163.367
R2491 B.n35 B.n34 163.367
R2492 B.n1197 B.n35 163.367
R2493 B.n1197 B.n40 163.367
R2494 B.n41 B.n40 163.367
R2495 B.n42 B.n41 163.367
R2496 B.n1202 B.n42 163.367
R2497 B.n1202 B.n47 163.367
R2498 B.n48 B.n47 163.367
R2499 B.n49 B.n48 163.367
R2500 B.n1207 B.n49 163.367
R2501 B.n1207 B.n54 163.367
R2502 B.n55 B.n54 163.367
R2503 B.n56 B.n55 163.367
R2504 B.n1212 B.n56 163.367
R2505 B.n1212 B.n61 163.367
R2506 B.n62 B.n61 163.367
R2507 B.n63 B.n62 163.367
R2508 B.n1217 B.n63 163.367
R2509 B.n1217 B.n68 163.367
R2510 B.n69 B.n68 163.367
R2511 B.n70 B.n69 163.367
R2512 B.n1222 B.n70 163.367
R2513 B.n1222 B.n75 163.367
R2514 B.n76 B.n75 163.367
R2515 B.n77 B.n76 163.367
R2516 B.n1227 B.n77 163.367
R2517 B.n1227 B.n82 163.367
R2518 B.n83 B.n82 163.367
R2519 B.n84 B.n83 163.367
R2520 B.n1232 B.n84 163.367
R2521 B.n1232 B.n89 163.367
R2522 B.n90 B.n89 163.367
R2523 B.n91 B.n90 163.367
R2524 B.n1237 B.n91 163.367
R2525 B.n1237 B.n96 163.367
R2526 B.n97 B.n96 163.367
R2527 B.n98 B.n97 163.367
R2528 B.n1242 B.n98 163.367
R2529 B.n1242 B.n103 163.367
R2530 B.n104 B.n103 163.367
R2531 B.n105 B.n104 163.367
R2532 B.n1247 B.n105 163.367
R2533 B.n1247 B.n110 163.367
R2534 B.n111 B.n110 163.367
R2535 B.n112 B.n111 163.367
R2536 B.n1252 B.n112 163.367
R2537 B.n1252 B.n117 163.367
R2538 B.n118 B.n117 163.367
R2539 B.n119 B.n118 163.367
R2540 B.n1257 B.n119 163.367
R2541 B.n1257 B.n124 163.367
R2542 B.n125 B.n124 163.367
R2543 B.n126 B.n125 163.367
R2544 B.n199 B.n126 163.367
R2545 B.n205 B.n130 163.367
R2546 B.n209 B.n208 163.367
R2547 B.n213 B.n212 163.367
R2548 B.n217 B.n216 163.367
R2549 B.n221 B.n220 163.367
R2550 B.n225 B.n224 163.367
R2551 B.n229 B.n228 163.367
R2552 B.n233 B.n232 163.367
R2553 B.n237 B.n236 163.367
R2554 B.n241 B.n240 163.367
R2555 B.n245 B.n244 163.367
R2556 B.n249 B.n248 163.367
R2557 B.n253 B.n252 163.367
R2558 B.n257 B.n256 163.367
R2559 B.n261 B.n260 163.367
R2560 B.n265 B.n264 163.367
R2561 B.n269 B.n268 163.367
R2562 B.n273 B.n272 163.367
R2563 B.n277 B.n276 163.367
R2564 B.n281 B.n280 163.367
R2565 B.n285 B.n284 163.367
R2566 B.n289 B.n288 163.367
R2567 B.n293 B.n292 163.367
R2568 B.n297 B.n296 163.367
R2569 B.n301 B.n300 163.367
R2570 B.n305 B.n304 163.367
R2571 B.n309 B.n308 163.367
R2572 B.n313 B.n312 163.367
R2573 B.n317 B.n316 163.367
R2574 B.n321 B.n320 163.367
R2575 B.n325 B.n324 163.367
R2576 B.n329 B.n328 163.367
R2577 B.n333 B.n332 163.367
R2578 B.n337 B.n336 163.367
R2579 B.n341 B.n340 163.367
R2580 B.n345 B.n344 163.367
R2581 B.n350 B.n349 163.367
R2582 B.n354 B.n353 163.367
R2583 B.n358 B.n357 163.367
R2584 B.n362 B.n361 163.367
R2585 B.n366 B.n365 163.367
R2586 B.n370 B.n369 163.367
R2587 B.n374 B.n373 163.367
R2588 B.n378 B.n377 163.367
R2589 B.n382 B.n381 163.367
R2590 B.n386 B.n385 163.367
R2591 B.n390 B.n389 163.367
R2592 B.n394 B.n393 163.367
R2593 B.n398 B.n397 163.367
R2594 B.n402 B.n401 163.367
R2595 B.n406 B.n405 163.367
R2596 B.n410 B.n409 163.367
R2597 B.n414 B.n413 163.367
R2598 B.n418 B.n417 163.367
R2599 B.n422 B.n421 163.367
R2600 B.n426 B.n425 163.367
R2601 B.n430 B.n429 163.367
R2602 B.n434 B.n433 163.367
R2603 B.n438 B.n437 163.367
R2604 B.n442 B.n441 163.367
R2605 B.n446 B.n445 163.367
R2606 B.n450 B.n449 163.367
R2607 B.n454 B.n453 163.367
R2608 B.n458 B.n457 163.367
R2609 B.n462 B.n461 163.367
R2610 B.n466 B.n465 163.367
R2611 B.n470 B.n469 163.367
R2612 B.n1264 B.n198 163.367
R2613 B.n957 B.n956 71.676
R2614 B.n679 B.n612 71.676
R2615 B.n949 B.n613 71.676
R2616 B.n945 B.n614 71.676
R2617 B.n941 B.n615 71.676
R2618 B.n937 B.n616 71.676
R2619 B.n933 B.n617 71.676
R2620 B.n929 B.n618 71.676
R2621 B.n925 B.n619 71.676
R2622 B.n921 B.n620 71.676
R2623 B.n917 B.n621 71.676
R2624 B.n913 B.n622 71.676
R2625 B.n909 B.n623 71.676
R2626 B.n905 B.n624 71.676
R2627 B.n901 B.n625 71.676
R2628 B.n897 B.n626 71.676
R2629 B.n893 B.n627 71.676
R2630 B.n889 B.n628 71.676
R2631 B.n885 B.n629 71.676
R2632 B.n881 B.n630 71.676
R2633 B.n877 B.n631 71.676
R2634 B.n873 B.n632 71.676
R2635 B.n869 B.n633 71.676
R2636 B.n865 B.n634 71.676
R2637 B.n861 B.n635 71.676
R2638 B.n857 B.n636 71.676
R2639 B.n853 B.n637 71.676
R2640 B.n849 B.n638 71.676
R2641 B.n845 B.n639 71.676
R2642 B.n841 B.n640 71.676
R2643 B.n837 B.n641 71.676
R2644 B.n833 B.n642 71.676
R2645 B.n828 B.n643 71.676
R2646 B.n824 B.n644 71.676
R2647 B.n820 B.n645 71.676
R2648 B.n816 B.n646 71.676
R2649 B.n812 B.n647 71.676
R2650 B.n808 B.n648 71.676
R2651 B.n804 B.n649 71.676
R2652 B.n800 B.n650 71.676
R2653 B.n796 B.n651 71.676
R2654 B.n792 B.n652 71.676
R2655 B.n788 B.n653 71.676
R2656 B.n784 B.n654 71.676
R2657 B.n780 B.n655 71.676
R2658 B.n776 B.n656 71.676
R2659 B.n772 B.n657 71.676
R2660 B.n768 B.n658 71.676
R2661 B.n764 B.n659 71.676
R2662 B.n760 B.n660 71.676
R2663 B.n756 B.n661 71.676
R2664 B.n752 B.n662 71.676
R2665 B.n748 B.n663 71.676
R2666 B.n744 B.n664 71.676
R2667 B.n740 B.n665 71.676
R2668 B.n736 B.n666 71.676
R2669 B.n732 B.n667 71.676
R2670 B.n728 B.n668 71.676
R2671 B.n724 B.n669 71.676
R2672 B.n720 B.n670 71.676
R2673 B.n716 B.n671 71.676
R2674 B.n712 B.n672 71.676
R2675 B.n708 B.n673 71.676
R2676 B.n704 B.n674 71.676
R2677 B.n700 B.n675 71.676
R2678 B.n696 B.n676 71.676
R2679 B.n692 B.n677 71.676
R2680 B.n688 B.n678 71.676
R2681 B.n1267 B.n1266 71.676
R2682 B.n205 B.n131 71.676
R2683 B.n209 B.n132 71.676
R2684 B.n213 B.n133 71.676
R2685 B.n217 B.n134 71.676
R2686 B.n221 B.n135 71.676
R2687 B.n225 B.n136 71.676
R2688 B.n229 B.n137 71.676
R2689 B.n233 B.n138 71.676
R2690 B.n237 B.n139 71.676
R2691 B.n241 B.n140 71.676
R2692 B.n245 B.n141 71.676
R2693 B.n249 B.n142 71.676
R2694 B.n253 B.n143 71.676
R2695 B.n257 B.n144 71.676
R2696 B.n261 B.n145 71.676
R2697 B.n265 B.n146 71.676
R2698 B.n269 B.n147 71.676
R2699 B.n273 B.n148 71.676
R2700 B.n277 B.n149 71.676
R2701 B.n281 B.n150 71.676
R2702 B.n285 B.n151 71.676
R2703 B.n289 B.n152 71.676
R2704 B.n293 B.n153 71.676
R2705 B.n297 B.n154 71.676
R2706 B.n301 B.n155 71.676
R2707 B.n305 B.n156 71.676
R2708 B.n309 B.n157 71.676
R2709 B.n313 B.n158 71.676
R2710 B.n317 B.n159 71.676
R2711 B.n321 B.n160 71.676
R2712 B.n325 B.n161 71.676
R2713 B.n329 B.n162 71.676
R2714 B.n333 B.n163 71.676
R2715 B.n337 B.n164 71.676
R2716 B.n341 B.n165 71.676
R2717 B.n345 B.n166 71.676
R2718 B.n350 B.n167 71.676
R2719 B.n354 B.n168 71.676
R2720 B.n358 B.n169 71.676
R2721 B.n362 B.n170 71.676
R2722 B.n366 B.n171 71.676
R2723 B.n370 B.n172 71.676
R2724 B.n374 B.n173 71.676
R2725 B.n378 B.n174 71.676
R2726 B.n382 B.n175 71.676
R2727 B.n386 B.n176 71.676
R2728 B.n390 B.n177 71.676
R2729 B.n394 B.n178 71.676
R2730 B.n398 B.n179 71.676
R2731 B.n402 B.n180 71.676
R2732 B.n406 B.n181 71.676
R2733 B.n410 B.n182 71.676
R2734 B.n414 B.n183 71.676
R2735 B.n418 B.n184 71.676
R2736 B.n422 B.n185 71.676
R2737 B.n426 B.n186 71.676
R2738 B.n430 B.n187 71.676
R2739 B.n434 B.n188 71.676
R2740 B.n438 B.n189 71.676
R2741 B.n442 B.n190 71.676
R2742 B.n446 B.n191 71.676
R2743 B.n450 B.n192 71.676
R2744 B.n454 B.n193 71.676
R2745 B.n458 B.n194 71.676
R2746 B.n462 B.n195 71.676
R2747 B.n466 B.n196 71.676
R2748 B.n470 B.n197 71.676
R2749 B.n198 B.n197 71.676
R2750 B.n469 B.n196 71.676
R2751 B.n465 B.n195 71.676
R2752 B.n461 B.n194 71.676
R2753 B.n457 B.n193 71.676
R2754 B.n453 B.n192 71.676
R2755 B.n449 B.n191 71.676
R2756 B.n445 B.n190 71.676
R2757 B.n441 B.n189 71.676
R2758 B.n437 B.n188 71.676
R2759 B.n433 B.n187 71.676
R2760 B.n429 B.n186 71.676
R2761 B.n425 B.n185 71.676
R2762 B.n421 B.n184 71.676
R2763 B.n417 B.n183 71.676
R2764 B.n413 B.n182 71.676
R2765 B.n409 B.n181 71.676
R2766 B.n405 B.n180 71.676
R2767 B.n401 B.n179 71.676
R2768 B.n397 B.n178 71.676
R2769 B.n393 B.n177 71.676
R2770 B.n389 B.n176 71.676
R2771 B.n385 B.n175 71.676
R2772 B.n381 B.n174 71.676
R2773 B.n377 B.n173 71.676
R2774 B.n373 B.n172 71.676
R2775 B.n369 B.n171 71.676
R2776 B.n365 B.n170 71.676
R2777 B.n361 B.n169 71.676
R2778 B.n357 B.n168 71.676
R2779 B.n353 B.n167 71.676
R2780 B.n349 B.n166 71.676
R2781 B.n344 B.n165 71.676
R2782 B.n340 B.n164 71.676
R2783 B.n336 B.n163 71.676
R2784 B.n332 B.n162 71.676
R2785 B.n328 B.n161 71.676
R2786 B.n324 B.n160 71.676
R2787 B.n320 B.n159 71.676
R2788 B.n316 B.n158 71.676
R2789 B.n312 B.n157 71.676
R2790 B.n308 B.n156 71.676
R2791 B.n304 B.n155 71.676
R2792 B.n300 B.n154 71.676
R2793 B.n296 B.n153 71.676
R2794 B.n292 B.n152 71.676
R2795 B.n288 B.n151 71.676
R2796 B.n284 B.n150 71.676
R2797 B.n280 B.n149 71.676
R2798 B.n276 B.n148 71.676
R2799 B.n272 B.n147 71.676
R2800 B.n268 B.n146 71.676
R2801 B.n264 B.n145 71.676
R2802 B.n260 B.n144 71.676
R2803 B.n256 B.n143 71.676
R2804 B.n252 B.n142 71.676
R2805 B.n248 B.n141 71.676
R2806 B.n244 B.n140 71.676
R2807 B.n240 B.n139 71.676
R2808 B.n236 B.n138 71.676
R2809 B.n232 B.n137 71.676
R2810 B.n228 B.n136 71.676
R2811 B.n224 B.n135 71.676
R2812 B.n220 B.n134 71.676
R2813 B.n216 B.n133 71.676
R2814 B.n212 B.n132 71.676
R2815 B.n208 B.n131 71.676
R2816 B.n1266 B.n130 71.676
R2817 B.n956 B.n611 71.676
R2818 B.n950 B.n612 71.676
R2819 B.n946 B.n613 71.676
R2820 B.n942 B.n614 71.676
R2821 B.n938 B.n615 71.676
R2822 B.n934 B.n616 71.676
R2823 B.n930 B.n617 71.676
R2824 B.n926 B.n618 71.676
R2825 B.n922 B.n619 71.676
R2826 B.n918 B.n620 71.676
R2827 B.n914 B.n621 71.676
R2828 B.n910 B.n622 71.676
R2829 B.n906 B.n623 71.676
R2830 B.n902 B.n624 71.676
R2831 B.n898 B.n625 71.676
R2832 B.n894 B.n626 71.676
R2833 B.n890 B.n627 71.676
R2834 B.n886 B.n628 71.676
R2835 B.n882 B.n629 71.676
R2836 B.n878 B.n630 71.676
R2837 B.n874 B.n631 71.676
R2838 B.n870 B.n632 71.676
R2839 B.n866 B.n633 71.676
R2840 B.n862 B.n634 71.676
R2841 B.n858 B.n635 71.676
R2842 B.n854 B.n636 71.676
R2843 B.n850 B.n637 71.676
R2844 B.n846 B.n638 71.676
R2845 B.n842 B.n639 71.676
R2846 B.n838 B.n640 71.676
R2847 B.n834 B.n641 71.676
R2848 B.n829 B.n642 71.676
R2849 B.n825 B.n643 71.676
R2850 B.n821 B.n644 71.676
R2851 B.n817 B.n645 71.676
R2852 B.n813 B.n646 71.676
R2853 B.n809 B.n647 71.676
R2854 B.n805 B.n648 71.676
R2855 B.n801 B.n649 71.676
R2856 B.n797 B.n650 71.676
R2857 B.n793 B.n651 71.676
R2858 B.n789 B.n652 71.676
R2859 B.n785 B.n653 71.676
R2860 B.n781 B.n654 71.676
R2861 B.n777 B.n655 71.676
R2862 B.n773 B.n656 71.676
R2863 B.n769 B.n657 71.676
R2864 B.n765 B.n658 71.676
R2865 B.n761 B.n659 71.676
R2866 B.n757 B.n660 71.676
R2867 B.n753 B.n661 71.676
R2868 B.n749 B.n662 71.676
R2869 B.n745 B.n663 71.676
R2870 B.n741 B.n664 71.676
R2871 B.n737 B.n665 71.676
R2872 B.n733 B.n666 71.676
R2873 B.n729 B.n667 71.676
R2874 B.n725 B.n668 71.676
R2875 B.n721 B.n669 71.676
R2876 B.n717 B.n670 71.676
R2877 B.n713 B.n671 71.676
R2878 B.n709 B.n672 71.676
R2879 B.n705 B.n673 71.676
R2880 B.n701 B.n674 71.676
R2881 B.n697 B.n675 71.676
R2882 B.n693 B.n676 71.676
R2883 B.n689 B.n677 71.676
R2884 B.n685 B.n678 71.676
R2885 B.n683 B.n682 69.0429
R2886 B.n681 B.n680 69.0429
R2887 B.n203 B.n202 69.0429
R2888 B.n201 B.n200 69.0429
R2889 B.n684 B.n683 59.5399
R2890 B.n831 B.n681 59.5399
R2891 B.n204 B.n203 59.5399
R2892 B.n347 B.n201 59.5399
R2893 B.n955 B.n608 52.666
R2894 B.n1265 B.n127 52.666
R2895 B.n1269 B.n1268 33.8737
R2896 B.n1263 B.n1262 33.8737
R2897 B.n686 B.n606 33.8737
R2898 B.n959 B.n958 33.8737
R2899 B.n962 B.n608 30.095
R2900 B.n962 B.n604 30.095
R2901 B.n968 B.n604 30.095
R2902 B.n968 B.n600 30.095
R2903 B.n974 B.n600 30.095
R2904 B.n974 B.n596 30.095
R2905 B.n981 B.n596 30.095
R2906 B.n981 B.n980 30.095
R2907 B.n987 B.n589 30.095
R2908 B.n993 B.n589 30.095
R2909 B.n993 B.n585 30.095
R2910 B.n999 B.n585 30.095
R2911 B.n999 B.n581 30.095
R2912 B.n1005 B.n581 30.095
R2913 B.n1005 B.n577 30.095
R2914 B.n1011 B.n577 30.095
R2915 B.n1011 B.n573 30.095
R2916 B.n1017 B.n573 30.095
R2917 B.n1017 B.n568 30.095
R2918 B.n1023 B.n568 30.095
R2919 B.n1023 B.n569 30.095
R2920 B.n1029 B.n561 30.095
R2921 B.n1035 B.n561 30.095
R2922 B.n1035 B.n557 30.095
R2923 B.n1041 B.n557 30.095
R2924 B.n1041 B.n553 30.095
R2925 B.n1047 B.n553 30.095
R2926 B.n1047 B.n549 30.095
R2927 B.n1054 B.n549 30.095
R2928 B.n1054 B.n1053 30.095
R2929 B.n1060 B.n542 30.095
R2930 B.n1066 B.n542 30.095
R2931 B.n1066 B.n538 30.095
R2932 B.n1072 B.n538 30.095
R2933 B.n1072 B.n534 30.095
R2934 B.n1078 B.n534 30.095
R2935 B.n1078 B.n530 30.095
R2936 B.n1084 B.n530 30.095
R2937 B.n1084 B.n526 30.095
R2938 B.n1090 B.n526 30.095
R2939 B.n1096 B.n522 30.095
R2940 B.n1096 B.n518 30.095
R2941 B.n1102 B.n518 30.095
R2942 B.n1102 B.n514 30.095
R2943 B.n1108 B.n514 30.095
R2944 B.n1108 B.n510 30.095
R2945 B.n1114 B.n510 30.095
R2946 B.n1114 B.n506 30.095
R2947 B.n1120 B.n506 30.095
R2948 B.n1126 B.n502 30.095
R2949 B.n1126 B.n498 30.095
R2950 B.n1132 B.n498 30.095
R2951 B.n1132 B.n494 30.095
R2952 B.n1138 B.n494 30.095
R2953 B.n1138 B.n490 30.095
R2954 B.n1144 B.n490 30.095
R2955 B.n1144 B.n486 30.095
R2956 B.n1151 B.n486 30.095
R2957 B.n1151 B.n1150 30.095
R2958 B.n1157 B.n479 30.095
R2959 B.n1164 B.n479 30.095
R2960 B.n1164 B.n475 30.095
R2961 B.n1170 B.n475 30.095
R2962 B.n1170 B.n4 30.095
R2963 B.n1410 B.n4 30.095
R2964 B.n1410 B.n1409 30.095
R2965 B.n1409 B.n1408 30.095
R2966 B.n1408 B.n8 30.095
R2967 B.n1402 B.n8 30.095
R2968 B.n1402 B.n1401 30.095
R2969 B.n1401 B.n1400 30.095
R2970 B.n1394 B.n18 30.095
R2971 B.n1394 B.n1393 30.095
R2972 B.n1393 B.n1392 30.095
R2973 B.n1392 B.n22 30.095
R2974 B.n1386 B.n22 30.095
R2975 B.n1386 B.n1385 30.095
R2976 B.n1385 B.n1384 30.095
R2977 B.n1384 B.n29 30.095
R2978 B.n1378 B.n29 30.095
R2979 B.n1378 B.n1377 30.095
R2980 B.n1376 B.n36 30.095
R2981 B.n1370 B.n36 30.095
R2982 B.n1370 B.n1369 30.095
R2983 B.n1369 B.n1368 30.095
R2984 B.n1368 B.n43 30.095
R2985 B.n1362 B.n43 30.095
R2986 B.n1362 B.n1361 30.095
R2987 B.n1361 B.n1360 30.095
R2988 B.n1360 B.n50 30.095
R2989 B.n1354 B.n1353 30.095
R2990 B.n1353 B.n1352 30.095
R2991 B.n1352 B.n57 30.095
R2992 B.n1346 B.n57 30.095
R2993 B.n1346 B.n1345 30.095
R2994 B.n1345 B.n1344 30.095
R2995 B.n1344 B.n64 30.095
R2996 B.n1338 B.n64 30.095
R2997 B.n1338 B.n1337 30.095
R2998 B.n1337 B.n1336 30.095
R2999 B.n1330 B.n74 30.095
R3000 B.n1330 B.n1329 30.095
R3001 B.n1329 B.n1328 30.095
R3002 B.n1328 B.n78 30.095
R3003 B.n1322 B.n78 30.095
R3004 B.n1322 B.n1321 30.095
R3005 B.n1321 B.n1320 30.095
R3006 B.n1320 B.n85 30.095
R3007 B.n1314 B.n85 30.095
R3008 B.n1313 B.n1312 30.095
R3009 B.n1312 B.n92 30.095
R3010 B.n1306 B.n92 30.095
R3011 B.n1306 B.n1305 30.095
R3012 B.n1305 B.n1304 30.095
R3013 B.n1304 B.n99 30.095
R3014 B.n1298 B.n99 30.095
R3015 B.n1298 B.n1297 30.095
R3016 B.n1297 B.n1296 30.095
R3017 B.n1296 B.n106 30.095
R3018 B.n1290 B.n106 30.095
R3019 B.n1290 B.n1289 30.095
R3020 B.n1289 B.n1288 30.095
R3021 B.n1282 B.n116 30.095
R3022 B.n1282 B.n1281 30.095
R3023 B.n1281 B.n1280 30.095
R3024 B.n1280 B.n120 30.095
R3025 B.n1274 B.n120 30.095
R3026 B.n1274 B.n1273 30.095
R3027 B.n1273 B.n1272 30.095
R3028 B.n1272 B.n127 30.095
R3029 B.n1157 B.t3 25.2268
R3030 B.n1400 B.t7 25.2268
R3031 B.t8 B.n522 23.4565
R3032 B.t1 B.n50 23.4565
R3033 B.n1053 B.t0 22.5714
R3034 B.n74 B.t9 22.5714
R3035 B.n1029 B.t4 21.6863
R3036 B.n1314 B.t2 21.6863
R3037 B.n1120 B.t5 20.8011
R3038 B.t6 B.n1376 20.8011
R3039 B.n980 B.t11 18.1457
R3040 B.n116 B.t15 18.1457
R3041 B B.n1412 18.0485
R3042 B.n987 B.t11 11.9498
R3043 B.n1288 B.t15 11.9498
R3044 B.n1268 B.n129 10.6151
R3045 B.n206 B.n129 10.6151
R3046 B.n207 B.n206 10.6151
R3047 B.n210 B.n207 10.6151
R3048 B.n211 B.n210 10.6151
R3049 B.n214 B.n211 10.6151
R3050 B.n215 B.n214 10.6151
R3051 B.n218 B.n215 10.6151
R3052 B.n219 B.n218 10.6151
R3053 B.n222 B.n219 10.6151
R3054 B.n223 B.n222 10.6151
R3055 B.n226 B.n223 10.6151
R3056 B.n227 B.n226 10.6151
R3057 B.n230 B.n227 10.6151
R3058 B.n231 B.n230 10.6151
R3059 B.n234 B.n231 10.6151
R3060 B.n235 B.n234 10.6151
R3061 B.n238 B.n235 10.6151
R3062 B.n239 B.n238 10.6151
R3063 B.n242 B.n239 10.6151
R3064 B.n243 B.n242 10.6151
R3065 B.n246 B.n243 10.6151
R3066 B.n247 B.n246 10.6151
R3067 B.n250 B.n247 10.6151
R3068 B.n251 B.n250 10.6151
R3069 B.n254 B.n251 10.6151
R3070 B.n255 B.n254 10.6151
R3071 B.n258 B.n255 10.6151
R3072 B.n259 B.n258 10.6151
R3073 B.n262 B.n259 10.6151
R3074 B.n263 B.n262 10.6151
R3075 B.n266 B.n263 10.6151
R3076 B.n267 B.n266 10.6151
R3077 B.n270 B.n267 10.6151
R3078 B.n271 B.n270 10.6151
R3079 B.n274 B.n271 10.6151
R3080 B.n275 B.n274 10.6151
R3081 B.n278 B.n275 10.6151
R3082 B.n279 B.n278 10.6151
R3083 B.n282 B.n279 10.6151
R3084 B.n283 B.n282 10.6151
R3085 B.n286 B.n283 10.6151
R3086 B.n287 B.n286 10.6151
R3087 B.n290 B.n287 10.6151
R3088 B.n291 B.n290 10.6151
R3089 B.n294 B.n291 10.6151
R3090 B.n295 B.n294 10.6151
R3091 B.n298 B.n295 10.6151
R3092 B.n299 B.n298 10.6151
R3093 B.n302 B.n299 10.6151
R3094 B.n303 B.n302 10.6151
R3095 B.n306 B.n303 10.6151
R3096 B.n307 B.n306 10.6151
R3097 B.n310 B.n307 10.6151
R3098 B.n311 B.n310 10.6151
R3099 B.n314 B.n311 10.6151
R3100 B.n315 B.n314 10.6151
R3101 B.n318 B.n315 10.6151
R3102 B.n319 B.n318 10.6151
R3103 B.n322 B.n319 10.6151
R3104 B.n323 B.n322 10.6151
R3105 B.n326 B.n323 10.6151
R3106 B.n327 B.n326 10.6151
R3107 B.n331 B.n330 10.6151
R3108 B.n334 B.n331 10.6151
R3109 B.n335 B.n334 10.6151
R3110 B.n338 B.n335 10.6151
R3111 B.n339 B.n338 10.6151
R3112 B.n342 B.n339 10.6151
R3113 B.n343 B.n342 10.6151
R3114 B.n346 B.n343 10.6151
R3115 B.n351 B.n348 10.6151
R3116 B.n352 B.n351 10.6151
R3117 B.n355 B.n352 10.6151
R3118 B.n356 B.n355 10.6151
R3119 B.n359 B.n356 10.6151
R3120 B.n360 B.n359 10.6151
R3121 B.n363 B.n360 10.6151
R3122 B.n364 B.n363 10.6151
R3123 B.n367 B.n364 10.6151
R3124 B.n368 B.n367 10.6151
R3125 B.n371 B.n368 10.6151
R3126 B.n372 B.n371 10.6151
R3127 B.n375 B.n372 10.6151
R3128 B.n376 B.n375 10.6151
R3129 B.n379 B.n376 10.6151
R3130 B.n380 B.n379 10.6151
R3131 B.n383 B.n380 10.6151
R3132 B.n384 B.n383 10.6151
R3133 B.n387 B.n384 10.6151
R3134 B.n388 B.n387 10.6151
R3135 B.n391 B.n388 10.6151
R3136 B.n392 B.n391 10.6151
R3137 B.n395 B.n392 10.6151
R3138 B.n396 B.n395 10.6151
R3139 B.n399 B.n396 10.6151
R3140 B.n400 B.n399 10.6151
R3141 B.n403 B.n400 10.6151
R3142 B.n404 B.n403 10.6151
R3143 B.n407 B.n404 10.6151
R3144 B.n408 B.n407 10.6151
R3145 B.n411 B.n408 10.6151
R3146 B.n412 B.n411 10.6151
R3147 B.n415 B.n412 10.6151
R3148 B.n416 B.n415 10.6151
R3149 B.n419 B.n416 10.6151
R3150 B.n420 B.n419 10.6151
R3151 B.n423 B.n420 10.6151
R3152 B.n424 B.n423 10.6151
R3153 B.n427 B.n424 10.6151
R3154 B.n428 B.n427 10.6151
R3155 B.n431 B.n428 10.6151
R3156 B.n432 B.n431 10.6151
R3157 B.n435 B.n432 10.6151
R3158 B.n436 B.n435 10.6151
R3159 B.n439 B.n436 10.6151
R3160 B.n440 B.n439 10.6151
R3161 B.n443 B.n440 10.6151
R3162 B.n444 B.n443 10.6151
R3163 B.n447 B.n444 10.6151
R3164 B.n448 B.n447 10.6151
R3165 B.n451 B.n448 10.6151
R3166 B.n452 B.n451 10.6151
R3167 B.n455 B.n452 10.6151
R3168 B.n456 B.n455 10.6151
R3169 B.n459 B.n456 10.6151
R3170 B.n460 B.n459 10.6151
R3171 B.n463 B.n460 10.6151
R3172 B.n464 B.n463 10.6151
R3173 B.n467 B.n464 10.6151
R3174 B.n468 B.n467 10.6151
R3175 B.n471 B.n468 10.6151
R3176 B.n472 B.n471 10.6151
R3177 B.n1263 B.n472 10.6151
R3178 B.n964 B.n606 10.6151
R3179 B.n965 B.n964 10.6151
R3180 B.n966 B.n965 10.6151
R3181 B.n966 B.n598 10.6151
R3182 B.n976 B.n598 10.6151
R3183 B.n977 B.n976 10.6151
R3184 B.n978 B.n977 10.6151
R3185 B.n978 B.n591 10.6151
R3186 B.n989 B.n591 10.6151
R3187 B.n990 B.n989 10.6151
R3188 B.n991 B.n990 10.6151
R3189 B.n991 B.n583 10.6151
R3190 B.n1001 B.n583 10.6151
R3191 B.n1002 B.n1001 10.6151
R3192 B.n1003 B.n1002 10.6151
R3193 B.n1003 B.n575 10.6151
R3194 B.n1013 B.n575 10.6151
R3195 B.n1014 B.n1013 10.6151
R3196 B.n1015 B.n1014 10.6151
R3197 B.n1015 B.n566 10.6151
R3198 B.n1025 B.n566 10.6151
R3199 B.n1026 B.n1025 10.6151
R3200 B.n1027 B.n1026 10.6151
R3201 B.n1027 B.n559 10.6151
R3202 B.n1037 B.n559 10.6151
R3203 B.n1038 B.n1037 10.6151
R3204 B.n1039 B.n1038 10.6151
R3205 B.n1039 B.n551 10.6151
R3206 B.n1049 B.n551 10.6151
R3207 B.n1050 B.n1049 10.6151
R3208 B.n1051 B.n1050 10.6151
R3209 B.n1051 B.n544 10.6151
R3210 B.n1062 B.n544 10.6151
R3211 B.n1063 B.n1062 10.6151
R3212 B.n1064 B.n1063 10.6151
R3213 B.n1064 B.n536 10.6151
R3214 B.n1074 B.n536 10.6151
R3215 B.n1075 B.n1074 10.6151
R3216 B.n1076 B.n1075 10.6151
R3217 B.n1076 B.n528 10.6151
R3218 B.n1086 B.n528 10.6151
R3219 B.n1087 B.n1086 10.6151
R3220 B.n1088 B.n1087 10.6151
R3221 B.n1088 B.n520 10.6151
R3222 B.n1098 B.n520 10.6151
R3223 B.n1099 B.n1098 10.6151
R3224 B.n1100 B.n1099 10.6151
R3225 B.n1100 B.n512 10.6151
R3226 B.n1110 B.n512 10.6151
R3227 B.n1111 B.n1110 10.6151
R3228 B.n1112 B.n1111 10.6151
R3229 B.n1112 B.n504 10.6151
R3230 B.n1122 B.n504 10.6151
R3231 B.n1123 B.n1122 10.6151
R3232 B.n1124 B.n1123 10.6151
R3233 B.n1124 B.n496 10.6151
R3234 B.n1134 B.n496 10.6151
R3235 B.n1135 B.n1134 10.6151
R3236 B.n1136 B.n1135 10.6151
R3237 B.n1136 B.n488 10.6151
R3238 B.n1146 B.n488 10.6151
R3239 B.n1147 B.n1146 10.6151
R3240 B.n1148 B.n1147 10.6151
R3241 B.n1148 B.n481 10.6151
R3242 B.n1159 B.n481 10.6151
R3243 B.n1160 B.n1159 10.6151
R3244 B.n1162 B.n1160 10.6151
R3245 B.n1162 B.n1161 10.6151
R3246 B.n1161 B.n473 10.6151
R3247 B.n1173 B.n473 10.6151
R3248 B.n1174 B.n1173 10.6151
R3249 B.n1175 B.n1174 10.6151
R3250 B.n1176 B.n1175 10.6151
R3251 B.n1178 B.n1176 10.6151
R3252 B.n1179 B.n1178 10.6151
R3253 B.n1180 B.n1179 10.6151
R3254 B.n1181 B.n1180 10.6151
R3255 B.n1183 B.n1181 10.6151
R3256 B.n1184 B.n1183 10.6151
R3257 B.n1185 B.n1184 10.6151
R3258 B.n1186 B.n1185 10.6151
R3259 B.n1188 B.n1186 10.6151
R3260 B.n1189 B.n1188 10.6151
R3261 B.n1190 B.n1189 10.6151
R3262 B.n1191 B.n1190 10.6151
R3263 B.n1193 B.n1191 10.6151
R3264 B.n1194 B.n1193 10.6151
R3265 B.n1195 B.n1194 10.6151
R3266 B.n1196 B.n1195 10.6151
R3267 B.n1198 B.n1196 10.6151
R3268 B.n1199 B.n1198 10.6151
R3269 B.n1200 B.n1199 10.6151
R3270 B.n1201 B.n1200 10.6151
R3271 B.n1203 B.n1201 10.6151
R3272 B.n1204 B.n1203 10.6151
R3273 B.n1205 B.n1204 10.6151
R3274 B.n1206 B.n1205 10.6151
R3275 B.n1208 B.n1206 10.6151
R3276 B.n1209 B.n1208 10.6151
R3277 B.n1210 B.n1209 10.6151
R3278 B.n1211 B.n1210 10.6151
R3279 B.n1213 B.n1211 10.6151
R3280 B.n1214 B.n1213 10.6151
R3281 B.n1215 B.n1214 10.6151
R3282 B.n1216 B.n1215 10.6151
R3283 B.n1218 B.n1216 10.6151
R3284 B.n1219 B.n1218 10.6151
R3285 B.n1220 B.n1219 10.6151
R3286 B.n1221 B.n1220 10.6151
R3287 B.n1223 B.n1221 10.6151
R3288 B.n1224 B.n1223 10.6151
R3289 B.n1225 B.n1224 10.6151
R3290 B.n1226 B.n1225 10.6151
R3291 B.n1228 B.n1226 10.6151
R3292 B.n1229 B.n1228 10.6151
R3293 B.n1230 B.n1229 10.6151
R3294 B.n1231 B.n1230 10.6151
R3295 B.n1233 B.n1231 10.6151
R3296 B.n1234 B.n1233 10.6151
R3297 B.n1235 B.n1234 10.6151
R3298 B.n1236 B.n1235 10.6151
R3299 B.n1238 B.n1236 10.6151
R3300 B.n1239 B.n1238 10.6151
R3301 B.n1240 B.n1239 10.6151
R3302 B.n1241 B.n1240 10.6151
R3303 B.n1243 B.n1241 10.6151
R3304 B.n1244 B.n1243 10.6151
R3305 B.n1245 B.n1244 10.6151
R3306 B.n1246 B.n1245 10.6151
R3307 B.n1248 B.n1246 10.6151
R3308 B.n1249 B.n1248 10.6151
R3309 B.n1250 B.n1249 10.6151
R3310 B.n1251 B.n1250 10.6151
R3311 B.n1253 B.n1251 10.6151
R3312 B.n1254 B.n1253 10.6151
R3313 B.n1255 B.n1254 10.6151
R3314 B.n1256 B.n1255 10.6151
R3315 B.n1258 B.n1256 10.6151
R3316 B.n1259 B.n1258 10.6151
R3317 B.n1260 B.n1259 10.6151
R3318 B.n1261 B.n1260 10.6151
R3319 B.n1262 B.n1261 10.6151
R3320 B.n958 B.n610 10.6151
R3321 B.n953 B.n610 10.6151
R3322 B.n953 B.n952 10.6151
R3323 B.n952 B.n951 10.6151
R3324 B.n951 B.n948 10.6151
R3325 B.n948 B.n947 10.6151
R3326 B.n947 B.n944 10.6151
R3327 B.n944 B.n943 10.6151
R3328 B.n943 B.n940 10.6151
R3329 B.n940 B.n939 10.6151
R3330 B.n939 B.n936 10.6151
R3331 B.n936 B.n935 10.6151
R3332 B.n935 B.n932 10.6151
R3333 B.n932 B.n931 10.6151
R3334 B.n931 B.n928 10.6151
R3335 B.n928 B.n927 10.6151
R3336 B.n927 B.n924 10.6151
R3337 B.n924 B.n923 10.6151
R3338 B.n923 B.n920 10.6151
R3339 B.n920 B.n919 10.6151
R3340 B.n919 B.n916 10.6151
R3341 B.n916 B.n915 10.6151
R3342 B.n915 B.n912 10.6151
R3343 B.n912 B.n911 10.6151
R3344 B.n911 B.n908 10.6151
R3345 B.n908 B.n907 10.6151
R3346 B.n907 B.n904 10.6151
R3347 B.n904 B.n903 10.6151
R3348 B.n903 B.n900 10.6151
R3349 B.n900 B.n899 10.6151
R3350 B.n899 B.n896 10.6151
R3351 B.n896 B.n895 10.6151
R3352 B.n895 B.n892 10.6151
R3353 B.n892 B.n891 10.6151
R3354 B.n891 B.n888 10.6151
R3355 B.n888 B.n887 10.6151
R3356 B.n887 B.n884 10.6151
R3357 B.n884 B.n883 10.6151
R3358 B.n883 B.n880 10.6151
R3359 B.n880 B.n879 10.6151
R3360 B.n879 B.n876 10.6151
R3361 B.n876 B.n875 10.6151
R3362 B.n875 B.n872 10.6151
R3363 B.n872 B.n871 10.6151
R3364 B.n871 B.n868 10.6151
R3365 B.n868 B.n867 10.6151
R3366 B.n867 B.n864 10.6151
R3367 B.n864 B.n863 10.6151
R3368 B.n863 B.n860 10.6151
R3369 B.n860 B.n859 10.6151
R3370 B.n859 B.n856 10.6151
R3371 B.n856 B.n855 10.6151
R3372 B.n855 B.n852 10.6151
R3373 B.n852 B.n851 10.6151
R3374 B.n851 B.n848 10.6151
R3375 B.n848 B.n847 10.6151
R3376 B.n847 B.n844 10.6151
R3377 B.n844 B.n843 10.6151
R3378 B.n843 B.n840 10.6151
R3379 B.n840 B.n839 10.6151
R3380 B.n839 B.n836 10.6151
R3381 B.n836 B.n835 10.6151
R3382 B.n835 B.n832 10.6151
R3383 B.n830 B.n827 10.6151
R3384 B.n827 B.n826 10.6151
R3385 B.n826 B.n823 10.6151
R3386 B.n823 B.n822 10.6151
R3387 B.n822 B.n819 10.6151
R3388 B.n819 B.n818 10.6151
R3389 B.n818 B.n815 10.6151
R3390 B.n815 B.n814 10.6151
R3391 B.n811 B.n810 10.6151
R3392 B.n810 B.n807 10.6151
R3393 B.n807 B.n806 10.6151
R3394 B.n806 B.n803 10.6151
R3395 B.n803 B.n802 10.6151
R3396 B.n802 B.n799 10.6151
R3397 B.n799 B.n798 10.6151
R3398 B.n798 B.n795 10.6151
R3399 B.n795 B.n794 10.6151
R3400 B.n794 B.n791 10.6151
R3401 B.n791 B.n790 10.6151
R3402 B.n790 B.n787 10.6151
R3403 B.n787 B.n786 10.6151
R3404 B.n786 B.n783 10.6151
R3405 B.n783 B.n782 10.6151
R3406 B.n782 B.n779 10.6151
R3407 B.n779 B.n778 10.6151
R3408 B.n778 B.n775 10.6151
R3409 B.n775 B.n774 10.6151
R3410 B.n774 B.n771 10.6151
R3411 B.n771 B.n770 10.6151
R3412 B.n770 B.n767 10.6151
R3413 B.n767 B.n766 10.6151
R3414 B.n766 B.n763 10.6151
R3415 B.n763 B.n762 10.6151
R3416 B.n762 B.n759 10.6151
R3417 B.n759 B.n758 10.6151
R3418 B.n758 B.n755 10.6151
R3419 B.n755 B.n754 10.6151
R3420 B.n754 B.n751 10.6151
R3421 B.n751 B.n750 10.6151
R3422 B.n750 B.n747 10.6151
R3423 B.n747 B.n746 10.6151
R3424 B.n746 B.n743 10.6151
R3425 B.n743 B.n742 10.6151
R3426 B.n742 B.n739 10.6151
R3427 B.n739 B.n738 10.6151
R3428 B.n738 B.n735 10.6151
R3429 B.n735 B.n734 10.6151
R3430 B.n734 B.n731 10.6151
R3431 B.n731 B.n730 10.6151
R3432 B.n730 B.n727 10.6151
R3433 B.n727 B.n726 10.6151
R3434 B.n726 B.n723 10.6151
R3435 B.n723 B.n722 10.6151
R3436 B.n722 B.n719 10.6151
R3437 B.n719 B.n718 10.6151
R3438 B.n718 B.n715 10.6151
R3439 B.n715 B.n714 10.6151
R3440 B.n714 B.n711 10.6151
R3441 B.n711 B.n710 10.6151
R3442 B.n710 B.n707 10.6151
R3443 B.n707 B.n706 10.6151
R3444 B.n706 B.n703 10.6151
R3445 B.n703 B.n702 10.6151
R3446 B.n702 B.n699 10.6151
R3447 B.n699 B.n698 10.6151
R3448 B.n698 B.n695 10.6151
R3449 B.n695 B.n694 10.6151
R3450 B.n694 B.n691 10.6151
R3451 B.n691 B.n690 10.6151
R3452 B.n690 B.n687 10.6151
R3453 B.n687 B.n686 10.6151
R3454 B.n960 B.n959 10.6151
R3455 B.n960 B.n602 10.6151
R3456 B.n970 B.n602 10.6151
R3457 B.n971 B.n970 10.6151
R3458 B.n972 B.n971 10.6151
R3459 B.n972 B.n594 10.6151
R3460 B.n983 B.n594 10.6151
R3461 B.n984 B.n983 10.6151
R3462 B.n985 B.n984 10.6151
R3463 B.n985 B.n587 10.6151
R3464 B.n995 B.n587 10.6151
R3465 B.n996 B.n995 10.6151
R3466 B.n997 B.n996 10.6151
R3467 B.n997 B.n579 10.6151
R3468 B.n1007 B.n579 10.6151
R3469 B.n1008 B.n1007 10.6151
R3470 B.n1009 B.n1008 10.6151
R3471 B.n1009 B.n571 10.6151
R3472 B.n1019 B.n571 10.6151
R3473 B.n1020 B.n1019 10.6151
R3474 B.n1021 B.n1020 10.6151
R3475 B.n1021 B.n563 10.6151
R3476 B.n1031 B.n563 10.6151
R3477 B.n1032 B.n1031 10.6151
R3478 B.n1033 B.n1032 10.6151
R3479 B.n1033 B.n555 10.6151
R3480 B.n1043 B.n555 10.6151
R3481 B.n1044 B.n1043 10.6151
R3482 B.n1045 B.n1044 10.6151
R3483 B.n1045 B.n547 10.6151
R3484 B.n1056 B.n547 10.6151
R3485 B.n1057 B.n1056 10.6151
R3486 B.n1058 B.n1057 10.6151
R3487 B.n1058 B.n540 10.6151
R3488 B.n1068 B.n540 10.6151
R3489 B.n1069 B.n1068 10.6151
R3490 B.n1070 B.n1069 10.6151
R3491 B.n1070 B.n532 10.6151
R3492 B.n1080 B.n532 10.6151
R3493 B.n1081 B.n1080 10.6151
R3494 B.n1082 B.n1081 10.6151
R3495 B.n1082 B.n524 10.6151
R3496 B.n1092 B.n524 10.6151
R3497 B.n1093 B.n1092 10.6151
R3498 B.n1094 B.n1093 10.6151
R3499 B.n1094 B.n516 10.6151
R3500 B.n1104 B.n516 10.6151
R3501 B.n1105 B.n1104 10.6151
R3502 B.n1106 B.n1105 10.6151
R3503 B.n1106 B.n508 10.6151
R3504 B.n1116 B.n508 10.6151
R3505 B.n1117 B.n1116 10.6151
R3506 B.n1118 B.n1117 10.6151
R3507 B.n1118 B.n500 10.6151
R3508 B.n1128 B.n500 10.6151
R3509 B.n1129 B.n1128 10.6151
R3510 B.n1130 B.n1129 10.6151
R3511 B.n1130 B.n492 10.6151
R3512 B.n1140 B.n492 10.6151
R3513 B.n1141 B.n1140 10.6151
R3514 B.n1142 B.n1141 10.6151
R3515 B.n1142 B.n484 10.6151
R3516 B.n1153 B.n484 10.6151
R3517 B.n1154 B.n1153 10.6151
R3518 B.n1155 B.n1154 10.6151
R3519 B.n1155 B.n477 10.6151
R3520 B.n1166 B.n477 10.6151
R3521 B.n1167 B.n1166 10.6151
R3522 B.n1168 B.n1167 10.6151
R3523 B.n1168 B.n0 10.6151
R3524 B.n1406 B.n1 10.6151
R3525 B.n1406 B.n1405 10.6151
R3526 B.n1405 B.n1404 10.6151
R3527 B.n1404 B.n10 10.6151
R3528 B.n1398 B.n10 10.6151
R3529 B.n1398 B.n1397 10.6151
R3530 B.n1397 B.n1396 10.6151
R3531 B.n1396 B.n16 10.6151
R3532 B.n1390 B.n16 10.6151
R3533 B.n1390 B.n1389 10.6151
R3534 B.n1389 B.n1388 10.6151
R3535 B.n1388 B.n24 10.6151
R3536 B.n1382 B.n24 10.6151
R3537 B.n1382 B.n1381 10.6151
R3538 B.n1381 B.n1380 10.6151
R3539 B.n1380 B.n31 10.6151
R3540 B.n1374 B.n31 10.6151
R3541 B.n1374 B.n1373 10.6151
R3542 B.n1373 B.n1372 10.6151
R3543 B.n1372 B.n38 10.6151
R3544 B.n1366 B.n38 10.6151
R3545 B.n1366 B.n1365 10.6151
R3546 B.n1365 B.n1364 10.6151
R3547 B.n1364 B.n45 10.6151
R3548 B.n1358 B.n45 10.6151
R3549 B.n1358 B.n1357 10.6151
R3550 B.n1357 B.n1356 10.6151
R3551 B.n1356 B.n52 10.6151
R3552 B.n1350 B.n52 10.6151
R3553 B.n1350 B.n1349 10.6151
R3554 B.n1349 B.n1348 10.6151
R3555 B.n1348 B.n59 10.6151
R3556 B.n1342 B.n59 10.6151
R3557 B.n1342 B.n1341 10.6151
R3558 B.n1341 B.n1340 10.6151
R3559 B.n1340 B.n66 10.6151
R3560 B.n1334 B.n66 10.6151
R3561 B.n1334 B.n1333 10.6151
R3562 B.n1333 B.n1332 10.6151
R3563 B.n1332 B.n72 10.6151
R3564 B.n1326 B.n72 10.6151
R3565 B.n1326 B.n1325 10.6151
R3566 B.n1325 B.n1324 10.6151
R3567 B.n1324 B.n80 10.6151
R3568 B.n1318 B.n80 10.6151
R3569 B.n1318 B.n1317 10.6151
R3570 B.n1317 B.n1316 10.6151
R3571 B.n1316 B.n87 10.6151
R3572 B.n1310 B.n87 10.6151
R3573 B.n1310 B.n1309 10.6151
R3574 B.n1309 B.n1308 10.6151
R3575 B.n1308 B.n94 10.6151
R3576 B.n1302 B.n94 10.6151
R3577 B.n1302 B.n1301 10.6151
R3578 B.n1301 B.n1300 10.6151
R3579 B.n1300 B.n101 10.6151
R3580 B.n1294 B.n101 10.6151
R3581 B.n1294 B.n1293 10.6151
R3582 B.n1293 B.n1292 10.6151
R3583 B.n1292 B.n108 10.6151
R3584 B.n1286 B.n108 10.6151
R3585 B.n1286 B.n1285 10.6151
R3586 B.n1285 B.n1284 10.6151
R3587 B.n1284 B.n114 10.6151
R3588 B.n1278 B.n114 10.6151
R3589 B.n1278 B.n1277 10.6151
R3590 B.n1277 B.n1276 10.6151
R3591 B.n1276 B.n122 10.6151
R3592 B.n1270 B.n122 10.6151
R3593 B.n1270 B.n1269 10.6151
R3594 B.t5 B.n502 9.2944
R3595 B.n1377 B.t6 9.2944
R3596 B.n569 B.t4 8.40927
R3597 B.t2 B.n1313 8.40927
R3598 B.n1060 B.t0 7.52414
R3599 B.n1336 B.t9 7.52414
R3600 B.n1090 B.t8 6.639
R3601 B.n1354 B.t1 6.639
R3602 B.n330 B.n204 6.5566
R3603 B.n347 B.n346 6.5566
R3604 B.n831 B.n830 6.5566
R3605 B.n814 B.n684 6.5566
R3606 B.n1150 B.t3 4.86874
R3607 B.n18 B.t7 4.86874
R3608 B.n327 B.n204 4.05904
R3609 B.n348 B.n347 4.05904
R3610 B.n832 B.n831 4.05904
R3611 B.n811 B.n684 4.05904
R3612 B.n1412 B.n0 2.81026
R3613 B.n1412 B.n1 2.81026
R3614 VP.n30 VP.t8 179.447
R3615 VP.n32 VP.n31 161.3
R3616 VP.n33 VP.n28 161.3
R3617 VP.n35 VP.n34 161.3
R3618 VP.n36 VP.n27 161.3
R3619 VP.n38 VP.n37 161.3
R3620 VP.n39 VP.n26 161.3
R3621 VP.n41 VP.n40 161.3
R3622 VP.n43 VP.n42 161.3
R3623 VP.n44 VP.n24 161.3
R3624 VP.n46 VP.n45 161.3
R3625 VP.n47 VP.n23 161.3
R3626 VP.n49 VP.n48 161.3
R3627 VP.n50 VP.n22 161.3
R3628 VP.n52 VP.n51 161.3
R3629 VP.n54 VP.n53 161.3
R3630 VP.n55 VP.n20 161.3
R3631 VP.n57 VP.n56 161.3
R3632 VP.n58 VP.n19 161.3
R3633 VP.n60 VP.n59 161.3
R3634 VP.n61 VP.n18 161.3
R3635 VP.n63 VP.n62 161.3
R3636 VP.n109 VP.n108 161.3
R3637 VP.n107 VP.n1 161.3
R3638 VP.n106 VP.n105 161.3
R3639 VP.n104 VP.n2 161.3
R3640 VP.n103 VP.n102 161.3
R3641 VP.n101 VP.n3 161.3
R3642 VP.n100 VP.n99 161.3
R3643 VP.n98 VP.n97 161.3
R3644 VP.n96 VP.n5 161.3
R3645 VP.n95 VP.n94 161.3
R3646 VP.n93 VP.n6 161.3
R3647 VP.n92 VP.n91 161.3
R3648 VP.n90 VP.n7 161.3
R3649 VP.n89 VP.n88 161.3
R3650 VP.n87 VP.n86 161.3
R3651 VP.n85 VP.n9 161.3
R3652 VP.n84 VP.n83 161.3
R3653 VP.n82 VP.n10 161.3
R3654 VP.n81 VP.n80 161.3
R3655 VP.n79 VP.n11 161.3
R3656 VP.n78 VP.n77 161.3
R3657 VP.n76 VP.n75 161.3
R3658 VP.n74 VP.n13 161.3
R3659 VP.n73 VP.n72 161.3
R3660 VP.n71 VP.n14 161.3
R3661 VP.n70 VP.n69 161.3
R3662 VP.n68 VP.n15 161.3
R3663 VP.n67 VP.n66 161.3
R3664 VP.n16 VP.t6 146.093
R3665 VP.n12 VP.t1 146.093
R3666 VP.n8 VP.t9 146.093
R3667 VP.n4 VP.t3 146.093
R3668 VP.n0 VP.t0 146.093
R3669 VP.n17 VP.t2 146.093
R3670 VP.n21 VP.t4 146.093
R3671 VP.n25 VP.t5 146.093
R3672 VP.n29 VP.t7 146.093
R3673 VP.n65 VP.n16 72.0476
R3674 VP.n110 VP.n0 72.0476
R3675 VP.n64 VP.n17 72.0476
R3676 VP.n65 VP.n64 62.4314
R3677 VP.n30 VP.n29 59.1355
R3678 VP.n69 VP.n14 49.296
R3679 VP.n106 VP.n2 49.296
R3680 VP.n60 VP.n19 49.296
R3681 VP.n80 VP.n10 43.4833
R3682 VP.n95 VP.n6 43.4833
R3683 VP.n49 VP.n23 43.4833
R3684 VP.n34 VP.n27 43.4833
R3685 VP.n84 VP.n10 37.6707
R3686 VP.n91 VP.n6 37.6707
R3687 VP.n45 VP.n23 37.6707
R3688 VP.n38 VP.n27 37.6707
R3689 VP.n73 VP.n14 31.8581
R3690 VP.n102 VP.n2 31.8581
R3691 VP.n56 VP.n19 31.8581
R3692 VP.n68 VP.n67 24.5923
R3693 VP.n69 VP.n68 24.5923
R3694 VP.n74 VP.n73 24.5923
R3695 VP.n75 VP.n74 24.5923
R3696 VP.n79 VP.n78 24.5923
R3697 VP.n80 VP.n79 24.5923
R3698 VP.n85 VP.n84 24.5923
R3699 VP.n86 VP.n85 24.5923
R3700 VP.n90 VP.n89 24.5923
R3701 VP.n91 VP.n90 24.5923
R3702 VP.n96 VP.n95 24.5923
R3703 VP.n97 VP.n96 24.5923
R3704 VP.n101 VP.n100 24.5923
R3705 VP.n102 VP.n101 24.5923
R3706 VP.n107 VP.n106 24.5923
R3707 VP.n108 VP.n107 24.5923
R3708 VP.n61 VP.n60 24.5923
R3709 VP.n62 VP.n61 24.5923
R3710 VP.n50 VP.n49 24.5923
R3711 VP.n51 VP.n50 24.5923
R3712 VP.n55 VP.n54 24.5923
R3713 VP.n56 VP.n55 24.5923
R3714 VP.n39 VP.n38 24.5923
R3715 VP.n40 VP.n39 24.5923
R3716 VP.n44 VP.n43 24.5923
R3717 VP.n45 VP.n44 24.5923
R3718 VP.n33 VP.n32 24.5923
R3719 VP.n34 VP.n33 24.5923
R3720 VP.n67 VP.n16 18.1985
R3721 VP.n108 VP.n0 18.1985
R3722 VP.n62 VP.n17 18.1985
R3723 VP.n78 VP.n12 15.2474
R3724 VP.n97 VP.n4 15.2474
R3725 VP.n51 VP.n21 15.2474
R3726 VP.n32 VP.n29 15.2474
R3727 VP.n86 VP.n8 12.2964
R3728 VP.n89 VP.n8 12.2964
R3729 VP.n40 VP.n25 12.2964
R3730 VP.n43 VP.n25 12.2964
R3731 VP.n75 VP.n12 9.3454
R3732 VP.n100 VP.n4 9.3454
R3733 VP.n54 VP.n21 9.3454
R3734 VP.n31 VP.n30 3.98081
R3735 VP.n64 VP.n63 0.354861
R3736 VP.n66 VP.n65 0.354861
R3737 VP.n110 VP.n109 0.354861
R3738 VP VP.n110 0.267071
R3739 VP.n31 VP.n28 0.189894
R3740 VP.n35 VP.n28 0.189894
R3741 VP.n36 VP.n35 0.189894
R3742 VP.n37 VP.n36 0.189894
R3743 VP.n37 VP.n26 0.189894
R3744 VP.n41 VP.n26 0.189894
R3745 VP.n42 VP.n41 0.189894
R3746 VP.n42 VP.n24 0.189894
R3747 VP.n46 VP.n24 0.189894
R3748 VP.n47 VP.n46 0.189894
R3749 VP.n48 VP.n47 0.189894
R3750 VP.n48 VP.n22 0.189894
R3751 VP.n52 VP.n22 0.189894
R3752 VP.n53 VP.n52 0.189894
R3753 VP.n53 VP.n20 0.189894
R3754 VP.n57 VP.n20 0.189894
R3755 VP.n58 VP.n57 0.189894
R3756 VP.n59 VP.n58 0.189894
R3757 VP.n59 VP.n18 0.189894
R3758 VP.n63 VP.n18 0.189894
R3759 VP.n66 VP.n15 0.189894
R3760 VP.n70 VP.n15 0.189894
R3761 VP.n71 VP.n70 0.189894
R3762 VP.n72 VP.n71 0.189894
R3763 VP.n72 VP.n13 0.189894
R3764 VP.n76 VP.n13 0.189894
R3765 VP.n77 VP.n76 0.189894
R3766 VP.n77 VP.n11 0.189894
R3767 VP.n81 VP.n11 0.189894
R3768 VP.n82 VP.n81 0.189894
R3769 VP.n83 VP.n82 0.189894
R3770 VP.n83 VP.n9 0.189894
R3771 VP.n87 VP.n9 0.189894
R3772 VP.n88 VP.n87 0.189894
R3773 VP.n88 VP.n7 0.189894
R3774 VP.n92 VP.n7 0.189894
R3775 VP.n93 VP.n92 0.189894
R3776 VP.n94 VP.n93 0.189894
R3777 VP.n94 VP.n5 0.189894
R3778 VP.n98 VP.n5 0.189894
R3779 VP.n99 VP.n98 0.189894
R3780 VP.n99 VP.n3 0.189894
R3781 VP.n103 VP.n3 0.189894
R3782 VP.n104 VP.n103 0.189894
R3783 VP.n105 VP.n104 0.189894
R3784 VP.n105 VP.n1 0.189894
R3785 VP.n109 VP.n1 0.189894
R3786 VDD1.n104 VDD1.n0 289.615
R3787 VDD1.n215 VDD1.n111 289.615
R3788 VDD1.n105 VDD1.n104 185
R3789 VDD1.n103 VDD1.n102 185
R3790 VDD1.n4 VDD1.n3 185
R3791 VDD1.n97 VDD1.n96 185
R3792 VDD1.n95 VDD1.n94 185
R3793 VDD1.n8 VDD1.n7 185
R3794 VDD1.n89 VDD1.n88 185
R3795 VDD1.n87 VDD1.n86 185
R3796 VDD1.n12 VDD1.n11 185
R3797 VDD1.n16 VDD1.n14 185
R3798 VDD1.n81 VDD1.n80 185
R3799 VDD1.n79 VDD1.n78 185
R3800 VDD1.n18 VDD1.n17 185
R3801 VDD1.n73 VDD1.n72 185
R3802 VDD1.n71 VDD1.n70 185
R3803 VDD1.n22 VDD1.n21 185
R3804 VDD1.n65 VDD1.n64 185
R3805 VDD1.n63 VDD1.n62 185
R3806 VDD1.n26 VDD1.n25 185
R3807 VDD1.n57 VDD1.n56 185
R3808 VDD1.n55 VDD1.n54 185
R3809 VDD1.n30 VDD1.n29 185
R3810 VDD1.n49 VDD1.n48 185
R3811 VDD1.n47 VDD1.n46 185
R3812 VDD1.n34 VDD1.n33 185
R3813 VDD1.n41 VDD1.n40 185
R3814 VDD1.n39 VDD1.n38 185
R3815 VDD1.n148 VDD1.n147 185
R3816 VDD1.n150 VDD1.n149 185
R3817 VDD1.n143 VDD1.n142 185
R3818 VDD1.n156 VDD1.n155 185
R3819 VDD1.n158 VDD1.n157 185
R3820 VDD1.n139 VDD1.n138 185
R3821 VDD1.n164 VDD1.n163 185
R3822 VDD1.n166 VDD1.n165 185
R3823 VDD1.n135 VDD1.n134 185
R3824 VDD1.n172 VDD1.n171 185
R3825 VDD1.n174 VDD1.n173 185
R3826 VDD1.n131 VDD1.n130 185
R3827 VDD1.n180 VDD1.n179 185
R3828 VDD1.n182 VDD1.n181 185
R3829 VDD1.n127 VDD1.n126 185
R3830 VDD1.n189 VDD1.n188 185
R3831 VDD1.n190 VDD1.n125 185
R3832 VDD1.n192 VDD1.n191 185
R3833 VDD1.n123 VDD1.n122 185
R3834 VDD1.n198 VDD1.n197 185
R3835 VDD1.n200 VDD1.n199 185
R3836 VDD1.n119 VDD1.n118 185
R3837 VDD1.n206 VDD1.n205 185
R3838 VDD1.n208 VDD1.n207 185
R3839 VDD1.n115 VDD1.n114 185
R3840 VDD1.n214 VDD1.n213 185
R3841 VDD1.n216 VDD1.n215 185
R3842 VDD1.n37 VDD1.t1 147.659
R3843 VDD1.n146 VDD1.t3 147.659
R3844 VDD1.n104 VDD1.n103 104.615
R3845 VDD1.n103 VDD1.n3 104.615
R3846 VDD1.n96 VDD1.n3 104.615
R3847 VDD1.n96 VDD1.n95 104.615
R3848 VDD1.n95 VDD1.n7 104.615
R3849 VDD1.n88 VDD1.n7 104.615
R3850 VDD1.n88 VDD1.n87 104.615
R3851 VDD1.n87 VDD1.n11 104.615
R3852 VDD1.n16 VDD1.n11 104.615
R3853 VDD1.n80 VDD1.n16 104.615
R3854 VDD1.n80 VDD1.n79 104.615
R3855 VDD1.n79 VDD1.n17 104.615
R3856 VDD1.n72 VDD1.n17 104.615
R3857 VDD1.n72 VDD1.n71 104.615
R3858 VDD1.n71 VDD1.n21 104.615
R3859 VDD1.n64 VDD1.n21 104.615
R3860 VDD1.n64 VDD1.n63 104.615
R3861 VDD1.n63 VDD1.n25 104.615
R3862 VDD1.n56 VDD1.n25 104.615
R3863 VDD1.n56 VDD1.n55 104.615
R3864 VDD1.n55 VDD1.n29 104.615
R3865 VDD1.n48 VDD1.n29 104.615
R3866 VDD1.n48 VDD1.n47 104.615
R3867 VDD1.n47 VDD1.n33 104.615
R3868 VDD1.n40 VDD1.n33 104.615
R3869 VDD1.n40 VDD1.n39 104.615
R3870 VDD1.n149 VDD1.n148 104.615
R3871 VDD1.n149 VDD1.n142 104.615
R3872 VDD1.n156 VDD1.n142 104.615
R3873 VDD1.n157 VDD1.n156 104.615
R3874 VDD1.n157 VDD1.n138 104.615
R3875 VDD1.n164 VDD1.n138 104.615
R3876 VDD1.n165 VDD1.n164 104.615
R3877 VDD1.n165 VDD1.n134 104.615
R3878 VDD1.n172 VDD1.n134 104.615
R3879 VDD1.n173 VDD1.n172 104.615
R3880 VDD1.n173 VDD1.n130 104.615
R3881 VDD1.n180 VDD1.n130 104.615
R3882 VDD1.n181 VDD1.n180 104.615
R3883 VDD1.n181 VDD1.n126 104.615
R3884 VDD1.n189 VDD1.n126 104.615
R3885 VDD1.n190 VDD1.n189 104.615
R3886 VDD1.n191 VDD1.n190 104.615
R3887 VDD1.n191 VDD1.n122 104.615
R3888 VDD1.n198 VDD1.n122 104.615
R3889 VDD1.n199 VDD1.n198 104.615
R3890 VDD1.n199 VDD1.n118 104.615
R3891 VDD1.n206 VDD1.n118 104.615
R3892 VDD1.n207 VDD1.n206 104.615
R3893 VDD1.n207 VDD1.n114 104.615
R3894 VDD1.n214 VDD1.n114 104.615
R3895 VDD1.n215 VDD1.n214 104.615
R3896 VDD1.n223 VDD1.n222 60.909
R3897 VDD1.n110 VDD1.n109 58.6628
R3898 VDD1.n225 VDD1.n224 58.6626
R3899 VDD1.n221 VDD1.n220 58.6626
R3900 VDD1.n225 VDD1.n223 57.2897
R3901 VDD1.n39 VDD1.t1 52.3082
R3902 VDD1.n148 VDD1.t3 52.3082
R3903 VDD1.n110 VDD1.n108 49.9937
R3904 VDD1.n221 VDD1.n219 49.9937
R3905 VDD1.n38 VDD1.n37 15.6677
R3906 VDD1.n147 VDD1.n146 15.6677
R3907 VDD1.n14 VDD1.n12 13.1884
R3908 VDD1.n192 VDD1.n123 13.1884
R3909 VDD1.n86 VDD1.n85 12.8005
R3910 VDD1.n82 VDD1.n81 12.8005
R3911 VDD1.n41 VDD1.n36 12.8005
R3912 VDD1.n150 VDD1.n145 12.8005
R3913 VDD1.n193 VDD1.n125 12.8005
R3914 VDD1.n197 VDD1.n196 12.8005
R3915 VDD1.n89 VDD1.n10 12.0247
R3916 VDD1.n78 VDD1.n15 12.0247
R3917 VDD1.n42 VDD1.n34 12.0247
R3918 VDD1.n151 VDD1.n143 12.0247
R3919 VDD1.n188 VDD1.n187 12.0247
R3920 VDD1.n200 VDD1.n121 12.0247
R3921 VDD1.n90 VDD1.n8 11.249
R3922 VDD1.n77 VDD1.n18 11.249
R3923 VDD1.n46 VDD1.n45 11.249
R3924 VDD1.n155 VDD1.n154 11.249
R3925 VDD1.n186 VDD1.n127 11.249
R3926 VDD1.n201 VDD1.n119 11.249
R3927 VDD1.n94 VDD1.n93 10.4732
R3928 VDD1.n74 VDD1.n73 10.4732
R3929 VDD1.n49 VDD1.n32 10.4732
R3930 VDD1.n158 VDD1.n141 10.4732
R3931 VDD1.n183 VDD1.n182 10.4732
R3932 VDD1.n205 VDD1.n204 10.4732
R3933 VDD1.n97 VDD1.n6 9.69747
R3934 VDD1.n70 VDD1.n20 9.69747
R3935 VDD1.n50 VDD1.n30 9.69747
R3936 VDD1.n159 VDD1.n139 9.69747
R3937 VDD1.n179 VDD1.n129 9.69747
R3938 VDD1.n208 VDD1.n117 9.69747
R3939 VDD1.n108 VDD1.n107 9.45567
R3940 VDD1.n219 VDD1.n218 9.45567
R3941 VDD1.n24 VDD1.n23 9.3005
R3942 VDD1.n67 VDD1.n66 9.3005
R3943 VDD1.n69 VDD1.n68 9.3005
R3944 VDD1.n20 VDD1.n19 9.3005
R3945 VDD1.n75 VDD1.n74 9.3005
R3946 VDD1.n77 VDD1.n76 9.3005
R3947 VDD1.n15 VDD1.n13 9.3005
R3948 VDD1.n83 VDD1.n82 9.3005
R3949 VDD1.n107 VDD1.n106 9.3005
R3950 VDD1.n2 VDD1.n1 9.3005
R3951 VDD1.n101 VDD1.n100 9.3005
R3952 VDD1.n99 VDD1.n98 9.3005
R3953 VDD1.n6 VDD1.n5 9.3005
R3954 VDD1.n93 VDD1.n92 9.3005
R3955 VDD1.n91 VDD1.n90 9.3005
R3956 VDD1.n10 VDD1.n9 9.3005
R3957 VDD1.n85 VDD1.n84 9.3005
R3958 VDD1.n61 VDD1.n60 9.3005
R3959 VDD1.n59 VDD1.n58 9.3005
R3960 VDD1.n28 VDD1.n27 9.3005
R3961 VDD1.n53 VDD1.n52 9.3005
R3962 VDD1.n51 VDD1.n50 9.3005
R3963 VDD1.n32 VDD1.n31 9.3005
R3964 VDD1.n45 VDD1.n44 9.3005
R3965 VDD1.n43 VDD1.n42 9.3005
R3966 VDD1.n36 VDD1.n35 9.3005
R3967 VDD1.n218 VDD1.n217 9.3005
R3968 VDD1.n212 VDD1.n211 9.3005
R3969 VDD1.n210 VDD1.n209 9.3005
R3970 VDD1.n117 VDD1.n116 9.3005
R3971 VDD1.n204 VDD1.n203 9.3005
R3972 VDD1.n202 VDD1.n201 9.3005
R3973 VDD1.n121 VDD1.n120 9.3005
R3974 VDD1.n196 VDD1.n195 9.3005
R3975 VDD1.n168 VDD1.n167 9.3005
R3976 VDD1.n137 VDD1.n136 9.3005
R3977 VDD1.n162 VDD1.n161 9.3005
R3978 VDD1.n160 VDD1.n159 9.3005
R3979 VDD1.n141 VDD1.n140 9.3005
R3980 VDD1.n154 VDD1.n153 9.3005
R3981 VDD1.n152 VDD1.n151 9.3005
R3982 VDD1.n145 VDD1.n144 9.3005
R3983 VDD1.n170 VDD1.n169 9.3005
R3984 VDD1.n133 VDD1.n132 9.3005
R3985 VDD1.n176 VDD1.n175 9.3005
R3986 VDD1.n178 VDD1.n177 9.3005
R3987 VDD1.n129 VDD1.n128 9.3005
R3988 VDD1.n184 VDD1.n183 9.3005
R3989 VDD1.n186 VDD1.n185 9.3005
R3990 VDD1.n187 VDD1.n124 9.3005
R3991 VDD1.n194 VDD1.n193 9.3005
R3992 VDD1.n113 VDD1.n112 9.3005
R3993 VDD1.n98 VDD1.n4 8.92171
R3994 VDD1.n69 VDD1.n22 8.92171
R3995 VDD1.n54 VDD1.n53 8.92171
R3996 VDD1.n163 VDD1.n162 8.92171
R3997 VDD1.n178 VDD1.n131 8.92171
R3998 VDD1.n209 VDD1.n115 8.92171
R3999 VDD1.n102 VDD1.n101 8.14595
R4000 VDD1.n66 VDD1.n65 8.14595
R4001 VDD1.n57 VDD1.n28 8.14595
R4002 VDD1.n166 VDD1.n137 8.14595
R4003 VDD1.n175 VDD1.n174 8.14595
R4004 VDD1.n213 VDD1.n212 8.14595
R4005 VDD1.n108 VDD1.n0 7.3702
R4006 VDD1.n105 VDD1.n2 7.3702
R4007 VDD1.n62 VDD1.n24 7.3702
R4008 VDD1.n58 VDD1.n26 7.3702
R4009 VDD1.n167 VDD1.n135 7.3702
R4010 VDD1.n171 VDD1.n133 7.3702
R4011 VDD1.n216 VDD1.n113 7.3702
R4012 VDD1.n219 VDD1.n111 7.3702
R4013 VDD1.n106 VDD1.n0 6.59444
R4014 VDD1.n106 VDD1.n105 6.59444
R4015 VDD1.n62 VDD1.n61 6.59444
R4016 VDD1.n61 VDD1.n26 6.59444
R4017 VDD1.n170 VDD1.n135 6.59444
R4018 VDD1.n171 VDD1.n170 6.59444
R4019 VDD1.n217 VDD1.n216 6.59444
R4020 VDD1.n217 VDD1.n111 6.59444
R4021 VDD1.n102 VDD1.n2 5.81868
R4022 VDD1.n65 VDD1.n24 5.81868
R4023 VDD1.n58 VDD1.n57 5.81868
R4024 VDD1.n167 VDD1.n166 5.81868
R4025 VDD1.n174 VDD1.n133 5.81868
R4026 VDD1.n213 VDD1.n113 5.81868
R4027 VDD1.n101 VDD1.n4 5.04292
R4028 VDD1.n66 VDD1.n22 5.04292
R4029 VDD1.n54 VDD1.n28 5.04292
R4030 VDD1.n163 VDD1.n137 5.04292
R4031 VDD1.n175 VDD1.n131 5.04292
R4032 VDD1.n212 VDD1.n115 5.04292
R4033 VDD1.n37 VDD1.n35 4.38563
R4034 VDD1.n146 VDD1.n144 4.38563
R4035 VDD1.n98 VDD1.n97 4.26717
R4036 VDD1.n70 VDD1.n69 4.26717
R4037 VDD1.n53 VDD1.n30 4.26717
R4038 VDD1.n162 VDD1.n139 4.26717
R4039 VDD1.n179 VDD1.n178 4.26717
R4040 VDD1.n209 VDD1.n208 4.26717
R4041 VDD1.n94 VDD1.n6 3.49141
R4042 VDD1.n73 VDD1.n20 3.49141
R4043 VDD1.n50 VDD1.n49 3.49141
R4044 VDD1.n159 VDD1.n158 3.49141
R4045 VDD1.n182 VDD1.n129 3.49141
R4046 VDD1.n205 VDD1.n117 3.49141
R4047 VDD1.n93 VDD1.n8 2.71565
R4048 VDD1.n74 VDD1.n18 2.71565
R4049 VDD1.n46 VDD1.n32 2.71565
R4050 VDD1.n155 VDD1.n141 2.71565
R4051 VDD1.n183 VDD1.n127 2.71565
R4052 VDD1.n204 VDD1.n119 2.71565
R4053 VDD1 VDD1.n225 2.24403
R4054 VDD1.n90 VDD1.n89 1.93989
R4055 VDD1.n78 VDD1.n77 1.93989
R4056 VDD1.n45 VDD1.n34 1.93989
R4057 VDD1.n154 VDD1.n143 1.93989
R4058 VDD1.n188 VDD1.n186 1.93989
R4059 VDD1.n201 VDD1.n200 1.93989
R4060 VDD1.n86 VDD1.n10 1.16414
R4061 VDD1.n81 VDD1.n15 1.16414
R4062 VDD1.n42 VDD1.n41 1.16414
R4063 VDD1.n151 VDD1.n150 1.16414
R4064 VDD1.n187 VDD1.n125 1.16414
R4065 VDD1.n197 VDD1.n121 1.16414
R4066 VDD1.n224 VDD1.t5 1.01174
R4067 VDD1.n224 VDD1.t7 1.01174
R4068 VDD1.n109 VDD1.t2 1.01174
R4069 VDD1.n109 VDD1.t4 1.01174
R4070 VDD1.n222 VDD1.t6 1.01174
R4071 VDD1.n222 VDD1.t9 1.01174
R4072 VDD1.n220 VDD1.t8 1.01174
R4073 VDD1.n220 VDD1.t0 1.01174
R4074 VDD1 VDD1.n110 0.825931
R4075 VDD1.n223 VDD1.n221 0.712395
R4076 VDD1.n85 VDD1.n12 0.388379
R4077 VDD1.n82 VDD1.n14 0.388379
R4078 VDD1.n38 VDD1.n36 0.388379
R4079 VDD1.n147 VDD1.n145 0.388379
R4080 VDD1.n193 VDD1.n192 0.388379
R4081 VDD1.n196 VDD1.n123 0.388379
R4082 VDD1.n107 VDD1.n1 0.155672
R4083 VDD1.n100 VDD1.n1 0.155672
R4084 VDD1.n100 VDD1.n99 0.155672
R4085 VDD1.n99 VDD1.n5 0.155672
R4086 VDD1.n92 VDD1.n5 0.155672
R4087 VDD1.n92 VDD1.n91 0.155672
R4088 VDD1.n91 VDD1.n9 0.155672
R4089 VDD1.n84 VDD1.n9 0.155672
R4090 VDD1.n84 VDD1.n83 0.155672
R4091 VDD1.n83 VDD1.n13 0.155672
R4092 VDD1.n76 VDD1.n13 0.155672
R4093 VDD1.n76 VDD1.n75 0.155672
R4094 VDD1.n75 VDD1.n19 0.155672
R4095 VDD1.n68 VDD1.n19 0.155672
R4096 VDD1.n68 VDD1.n67 0.155672
R4097 VDD1.n67 VDD1.n23 0.155672
R4098 VDD1.n60 VDD1.n23 0.155672
R4099 VDD1.n60 VDD1.n59 0.155672
R4100 VDD1.n59 VDD1.n27 0.155672
R4101 VDD1.n52 VDD1.n27 0.155672
R4102 VDD1.n52 VDD1.n51 0.155672
R4103 VDD1.n51 VDD1.n31 0.155672
R4104 VDD1.n44 VDD1.n31 0.155672
R4105 VDD1.n44 VDD1.n43 0.155672
R4106 VDD1.n43 VDD1.n35 0.155672
R4107 VDD1.n152 VDD1.n144 0.155672
R4108 VDD1.n153 VDD1.n152 0.155672
R4109 VDD1.n153 VDD1.n140 0.155672
R4110 VDD1.n160 VDD1.n140 0.155672
R4111 VDD1.n161 VDD1.n160 0.155672
R4112 VDD1.n161 VDD1.n136 0.155672
R4113 VDD1.n168 VDD1.n136 0.155672
R4114 VDD1.n169 VDD1.n168 0.155672
R4115 VDD1.n169 VDD1.n132 0.155672
R4116 VDD1.n176 VDD1.n132 0.155672
R4117 VDD1.n177 VDD1.n176 0.155672
R4118 VDD1.n177 VDD1.n128 0.155672
R4119 VDD1.n184 VDD1.n128 0.155672
R4120 VDD1.n185 VDD1.n184 0.155672
R4121 VDD1.n185 VDD1.n124 0.155672
R4122 VDD1.n194 VDD1.n124 0.155672
R4123 VDD1.n195 VDD1.n194 0.155672
R4124 VDD1.n195 VDD1.n120 0.155672
R4125 VDD1.n202 VDD1.n120 0.155672
R4126 VDD1.n203 VDD1.n202 0.155672
R4127 VDD1.n203 VDD1.n116 0.155672
R4128 VDD1.n210 VDD1.n116 0.155672
R4129 VDD1.n211 VDD1.n210 0.155672
R4130 VDD1.n211 VDD1.n112 0.155672
R4131 VDD1.n218 VDD1.n112 0.155672
C0 VDD1 VDD2 2.58391f
C1 VP VN 10.7228f
C2 VP VTAIL 18.350199f
C3 VP VDD1 18.2786f
C4 VN VTAIL 18.3359f
C5 VN VDD1 0.154915f
C6 VP VDD2 0.664579f
C7 VTAIL VDD1 13.792099f
C8 VN VDD2 17.774f
C9 VTAIL VDD2 13.8464f
C10 VDD2 B 9.257039f
C11 VDD1 B 9.245883f
C12 VTAIL B 11.748511f
C13 VN B 21.739967f
C14 VP B 20.219912f
C15 VDD1.n0 B 0.033064f
C16 VDD1.n1 B 0.023751f
C17 VDD1.n2 B 0.012763f
C18 VDD1.n3 B 0.030167f
C19 VDD1.n4 B 0.013514f
C20 VDD1.n5 B 0.023751f
C21 VDD1.n6 B 0.012763f
C22 VDD1.n7 B 0.030167f
C23 VDD1.n8 B 0.013514f
C24 VDD1.n9 B 0.023751f
C25 VDD1.n10 B 0.012763f
C26 VDD1.n11 B 0.030167f
C27 VDD1.n12 B 0.013138f
C28 VDD1.n13 B 0.023751f
C29 VDD1.n14 B 0.013138f
C30 VDD1.n15 B 0.012763f
C31 VDD1.n16 B 0.030167f
C32 VDD1.n17 B 0.030167f
C33 VDD1.n18 B 0.013514f
C34 VDD1.n19 B 0.023751f
C35 VDD1.n20 B 0.012763f
C36 VDD1.n21 B 0.030167f
C37 VDD1.n22 B 0.013514f
C38 VDD1.n23 B 0.023751f
C39 VDD1.n24 B 0.012763f
C40 VDD1.n25 B 0.030167f
C41 VDD1.n26 B 0.013514f
C42 VDD1.n27 B 0.023751f
C43 VDD1.n28 B 0.012763f
C44 VDD1.n29 B 0.030167f
C45 VDD1.n30 B 0.013514f
C46 VDD1.n31 B 0.023751f
C47 VDD1.n32 B 0.012763f
C48 VDD1.n33 B 0.030167f
C49 VDD1.n34 B 0.013514f
C50 VDD1.n35 B 2.04383f
C51 VDD1.n36 B 0.012763f
C52 VDD1.t1 B 0.050114f
C53 VDD1.n37 B 0.182184f
C54 VDD1.n38 B 0.01782f
C55 VDD1.n39 B 0.022625f
C56 VDD1.n40 B 0.030167f
C57 VDD1.n41 B 0.013514f
C58 VDD1.n42 B 0.012763f
C59 VDD1.n43 B 0.023751f
C60 VDD1.n44 B 0.023751f
C61 VDD1.n45 B 0.012763f
C62 VDD1.n46 B 0.013514f
C63 VDD1.n47 B 0.030167f
C64 VDD1.n48 B 0.030167f
C65 VDD1.n49 B 0.013514f
C66 VDD1.n50 B 0.012763f
C67 VDD1.n51 B 0.023751f
C68 VDD1.n52 B 0.023751f
C69 VDD1.n53 B 0.012763f
C70 VDD1.n54 B 0.013514f
C71 VDD1.n55 B 0.030167f
C72 VDD1.n56 B 0.030167f
C73 VDD1.n57 B 0.013514f
C74 VDD1.n58 B 0.012763f
C75 VDD1.n59 B 0.023751f
C76 VDD1.n60 B 0.023751f
C77 VDD1.n61 B 0.012763f
C78 VDD1.n62 B 0.013514f
C79 VDD1.n63 B 0.030167f
C80 VDD1.n64 B 0.030167f
C81 VDD1.n65 B 0.013514f
C82 VDD1.n66 B 0.012763f
C83 VDD1.n67 B 0.023751f
C84 VDD1.n68 B 0.023751f
C85 VDD1.n69 B 0.012763f
C86 VDD1.n70 B 0.013514f
C87 VDD1.n71 B 0.030167f
C88 VDD1.n72 B 0.030167f
C89 VDD1.n73 B 0.013514f
C90 VDD1.n74 B 0.012763f
C91 VDD1.n75 B 0.023751f
C92 VDD1.n76 B 0.023751f
C93 VDD1.n77 B 0.012763f
C94 VDD1.n78 B 0.013514f
C95 VDD1.n79 B 0.030167f
C96 VDD1.n80 B 0.030167f
C97 VDD1.n81 B 0.013514f
C98 VDD1.n82 B 0.012763f
C99 VDD1.n83 B 0.023751f
C100 VDD1.n84 B 0.023751f
C101 VDD1.n85 B 0.012763f
C102 VDD1.n86 B 0.013514f
C103 VDD1.n87 B 0.030167f
C104 VDD1.n88 B 0.030167f
C105 VDD1.n89 B 0.013514f
C106 VDD1.n90 B 0.012763f
C107 VDD1.n91 B 0.023751f
C108 VDD1.n92 B 0.023751f
C109 VDD1.n93 B 0.012763f
C110 VDD1.n94 B 0.013514f
C111 VDD1.n95 B 0.030167f
C112 VDD1.n96 B 0.030167f
C113 VDD1.n97 B 0.013514f
C114 VDD1.n98 B 0.012763f
C115 VDD1.n99 B 0.023751f
C116 VDD1.n100 B 0.023751f
C117 VDD1.n101 B 0.012763f
C118 VDD1.n102 B 0.013514f
C119 VDD1.n103 B 0.030167f
C120 VDD1.n104 B 0.064739f
C121 VDD1.n105 B 0.013514f
C122 VDD1.n106 B 0.012763f
C123 VDD1.n107 B 0.051655f
C124 VDD1.n108 B 0.069603f
C125 VDD1.t2 B 0.367495f
C126 VDD1.t4 B 0.367495f
C127 VDD1.n109 B 3.35553f
C128 VDD1.n110 B 0.761363f
C129 VDD1.n111 B 0.033064f
C130 VDD1.n112 B 0.023751f
C131 VDD1.n113 B 0.012763f
C132 VDD1.n114 B 0.030167f
C133 VDD1.n115 B 0.013514f
C134 VDD1.n116 B 0.023751f
C135 VDD1.n117 B 0.012763f
C136 VDD1.n118 B 0.030167f
C137 VDD1.n119 B 0.013514f
C138 VDD1.n120 B 0.023751f
C139 VDD1.n121 B 0.012763f
C140 VDD1.n122 B 0.030167f
C141 VDD1.n123 B 0.013138f
C142 VDD1.n124 B 0.023751f
C143 VDD1.n125 B 0.013514f
C144 VDD1.n126 B 0.030167f
C145 VDD1.n127 B 0.013514f
C146 VDD1.n128 B 0.023751f
C147 VDD1.n129 B 0.012763f
C148 VDD1.n130 B 0.030167f
C149 VDD1.n131 B 0.013514f
C150 VDD1.n132 B 0.023751f
C151 VDD1.n133 B 0.012763f
C152 VDD1.n134 B 0.030167f
C153 VDD1.n135 B 0.013514f
C154 VDD1.n136 B 0.023751f
C155 VDD1.n137 B 0.012763f
C156 VDD1.n138 B 0.030167f
C157 VDD1.n139 B 0.013514f
C158 VDD1.n140 B 0.023751f
C159 VDD1.n141 B 0.012763f
C160 VDD1.n142 B 0.030167f
C161 VDD1.n143 B 0.013514f
C162 VDD1.n144 B 2.04383f
C163 VDD1.n145 B 0.012763f
C164 VDD1.t3 B 0.050114f
C165 VDD1.n146 B 0.182184f
C166 VDD1.n147 B 0.01782f
C167 VDD1.n148 B 0.022625f
C168 VDD1.n149 B 0.030167f
C169 VDD1.n150 B 0.013514f
C170 VDD1.n151 B 0.012763f
C171 VDD1.n152 B 0.023751f
C172 VDD1.n153 B 0.023751f
C173 VDD1.n154 B 0.012763f
C174 VDD1.n155 B 0.013514f
C175 VDD1.n156 B 0.030167f
C176 VDD1.n157 B 0.030167f
C177 VDD1.n158 B 0.013514f
C178 VDD1.n159 B 0.012763f
C179 VDD1.n160 B 0.023751f
C180 VDD1.n161 B 0.023751f
C181 VDD1.n162 B 0.012763f
C182 VDD1.n163 B 0.013514f
C183 VDD1.n164 B 0.030167f
C184 VDD1.n165 B 0.030167f
C185 VDD1.n166 B 0.013514f
C186 VDD1.n167 B 0.012763f
C187 VDD1.n168 B 0.023751f
C188 VDD1.n169 B 0.023751f
C189 VDD1.n170 B 0.012763f
C190 VDD1.n171 B 0.013514f
C191 VDD1.n172 B 0.030167f
C192 VDD1.n173 B 0.030167f
C193 VDD1.n174 B 0.013514f
C194 VDD1.n175 B 0.012763f
C195 VDD1.n176 B 0.023751f
C196 VDD1.n177 B 0.023751f
C197 VDD1.n178 B 0.012763f
C198 VDD1.n179 B 0.013514f
C199 VDD1.n180 B 0.030167f
C200 VDD1.n181 B 0.030167f
C201 VDD1.n182 B 0.013514f
C202 VDD1.n183 B 0.012763f
C203 VDD1.n184 B 0.023751f
C204 VDD1.n185 B 0.023751f
C205 VDD1.n186 B 0.012763f
C206 VDD1.n187 B 0.012763f
C207 VDD1.n188 B 0.013514f
C208 VDD1.n189 B 0.030167f
C209 VDD1.n190 B 0.030167f
C210 VDD1.n191 B 0.030167f
C211 VDD1.n192 B 0.013138f
C212 VDD1.n193 B 0.012763f
C213 VDD1.n194 B 0.023751f
C214 VDD1.n195 B 0.023751f
C215 VDD1.n196 B 0.012763f
C216 VDD1.n197 B 0.013514f
C217 VDD1.n198 B 0.030167f
C218 VDD1.n199 B 0.030167f
C219 VDD1.n200 B 0.013514f
C220 VDD1.n201 B 0.012763f
C221 VDD1.n202 B 0.023751f
C222 VDD1.n203 B 0.023751f
C223 VDD1.n204 B 0.012763f
C224 VDD1.n205 B 0.013514f
C225 VDD1.n206 B 0.030167f
C226 VDD1.n207 B 0.030167f
C227 VDD1.n208 B 0.013514f
C228 VDD1.n209 B 0.012763f
C229 VDD1.n210 B 0.023751f
C230 VDD1.n211 B 0.023751f
C231 VDD1.n212 B 0.012763f
C232 VDD1.n213 B 0.013514f
C233 VDD1.n214 B 0.030167f
C234 VDD1.n215 B 0.064739f
C235 VDD1.n216 B 0.013514f
C236 VDD1.n217 B 0.012763f
C237 VDD1.n218 B 0.051655f
C238 VDD1.n219 B 0.069603f
C239 VDD1.t8 B 0.367495f
C240 VDD1.t0 B 0.367495f
C241 VDD1.n220 B 3.35552f
C242 VDD1.n221 B 0.753458f
C243 VDD1.t6 B 0.367495f
C244 VDD1.t9 B 0.367495f
C245 VDD1.n222 B 3.37832f
C246 VDD1.n223 B 3.67028f
C247 VDD1.t5 B 0.367495f
C248 VDD1.t7 B 0.367495f
C249 VDD1.n224 B 3.35552f
C250 VDD1.n225 B 3.81066f
C251 VP.t0 B 3.09148f
C252 VP.n0 B 1.1366f
C253 VP.n1 B 0.017745f
C254 VP.n2 B 0.016253f
C255 VP.n3 B 0.017745f
C256 VP.t3 B 3.09148f
C257 VP.n4 B 1.06459f
C258 VP.n5 B 0.017745f
C259 VP.n6 B 0.014536f
C260 VP.n7 B 0.017745f
C261 VP.t9 B 3.09148f
C262 VP.n8 B 1.06459f
C263 VP.n9 B 0.017745f
C264 VP.n10 B 0.014536f
C265 VP.n11 B 0.017745f
C266 VP.t1 B 3.09148f
C267 VP.n12 B 1.06459f
C268 VP.n13 B 0.017745f
C269 VP.n14 B 0.016253f
C270 VP.n15 B 0.017745f
C271 VP.t6 B 3.09148f
C272 VP.n16 B 1.1366f
C273 VP.t2 B 3.09148f
C274 VP.n17 B 1.1366f
C275 VP.n18 B 0.017745f
C276 VP.n19 B 0.016253f
C277 VP.n20 B 0.017745f
C278 VP.t4 B 3.09148f
C279 VP.n21 B 1.06459f
C280 VP.n22 B 0.017745f
C281 VP.n23 B 0.014536f
C282 VP.n24 B 0.017745f
C283 VP.t5 B 3.09148f
C284 VP.n25 B 1.06459f
C285 VP.n26 B 0.017745f
C286 VP.n27 B 0.014536f
C287 VP.n28 B 0.017745f
C288 VP.t7 B 3.09148f
C289 VP.n29 B 1.1247f
C290 VP.t8 B 3.31299f
C291 VP.n30 B 1.08141f
C292 VP.n31 B 0.205688f
C293 VP.n32 B 0.026733f
C294 VP.n33 B 0.032906f
C295 VP.n34 B 0.034459f
C296 VP.n35 B 0.017745f
C297 VP.n36 B 0.017745f
C298 VP.n37 B 0.017745f
C299 VP.n38 B 0.0355f
C300 VP.n39 B 0.032906f
C301 VP.n40 B 0.024784f
C302 VP.n41 B 0.017745f
C303 VP.n42 B 0.017745f
C304 VP.n43 B 0.024784f
C305 VP.n44 B 0.032906f
C306 VP.n45 B 0.0355f
C307 VP.n46 B 0.017745f
C308 VP.n47 B 0.017745f
C309 VP.n48 B 0.017745f
C310 VP.n49 B 0.034459f
C311 VP.n50 B 0.032906f
C312 VP.n51 B 0.026733f
C313 VP.n52 B 0.017745f
C314 VP.n53 B 0.017745f
C315 VP.n54 B 0.022834f
C316 VP.n55 B 0.032906f
C317 VP.n56 B 0.035499f
C318 VP.n57 B 0.017745f
C319 VP.n58 B 0.017745f
C320 VP.n59 B 0.017745f
C321 VP.n60 B 0.032743f
C322 VP.n61 B 0.032906f
C323 VP.n62 B 0.028682f
C324 VP.n63 B 0.028635f
C325 VP.n64 B 1.36713f
C326 VP.n65 B 1.37738f
C327 VP.n66 B 0.028635f
C328 VP.n67 B 0.028682f
C329 VP.n68 B 0.032906f
C330 VP.n69 B 0.032743f
C331 VP.n70 B 0.017745f
C332 VP.n71 B 0.017745f
C333 VP.n72 B 0.017745f
C334 VP.n73 B 0.035499f
C335 VP.n74 B 0.032906f
C336 VP.n75 B 0.022834f
C337 VP.n76 B 0.017745f
C338 VP.n77 B 0.017745f
C339 VP.n78 B 0.026733f
C340 VP.n79 B 0.032906f
C341 VP.n80 B 0.034459f
C342 VP.n81 B 0.017745f
C343 VP.n82 B 0.017745f
C344 VP.n83 B 0.017745f
C345 VP.n84 B 0.0355f
C346 VP.n85 B 0.032906f
C347 VP.n86 B 0.024784f
C348 VP.n87 B 0.017745f
C349 VP.n88 B 0.017745f
C350 VP.n89 B 0.024784f
C351 VP.n90 B 0.032906f
C352 VP.n91 B 0.0355f
C353 VP.n92 B 0.017745f
C354 VP.n93 B 0.017745f
C355 VP.n94 B 0.017745f
C356 VP.n95 B 0.034459f
C357 VP.n96 B 0.032906f
C358 VP.n97 B 0.026733f
C359 VP.n98 B 0.017745f
C360 VP.n99 B 0.017745f
C361 VP.n100 B 0.022834f
C362 VP.n101 B 0.032906f
C363 VP.n102 B 0.035499f
C364 VP.n103 B 0.017745f
C365 VP.n104 B 0.017745f
C366 VP.n105 B 0.017745f
C367 VP.n106 B 0.032743f
C368 VP.n107 B 0.032906f
C369 VP.n108 B 0.028682f
C370 VP.n109 B 0.028635f
C371 VP.n110 B 0.039826f
C372 VDD2.n0 B 0.03267f
C373 VDD2.n1 B 0.023468f
C374 VDD2.n2 B 0.012611f
C375 VDD2.n3 B 0.029807f
C376 VDD2.n4 B 0.013353f
C377 VDD2.n5 B 0.023468f
C378 VDD2.n6 B 0.012611f
C379 VDD2.n7 B 0.029807f
C380 VDD2.n8 B 0.013353f
C381 VDD2.n9 B 0.023468f
C382 VDD2.n10 B 0.012611f
C383 VDD2.n11 B 0.029807f
C384 VDD2.n12 B 0.012982f
C385 VDD2.n13 B 0.023468f
C386 VDD2.n14 B 0.013353f
C387 VDD2.n15 B 0.029807f
C388 VDD2.n16 B 0.013353f
C389 VDD2.n17 B 0.023468f
C390 VDD2.n18 B 0.012611f
C391 VDD2.n19 B 0.029807f
C392 VDD2.n20 B 0.013353f
C393 VDD2.n21 B 0.023468f
C394 VDD2.n22 B 0.012611f
C395 VDD2.n23 B 0.029807f
C396 VDD2.n24 B 0.013353f
C397 VDD2.n25 B 0.023468f
C398 VDD2.n26 B 0.012611f
C399 VDD2.n27 B 0.029807f
C400 VDD2.n28 B 0.013353f
C401 VDD2.n29 B 0.023468f
C402 VDD2.n30 B 0.012611f
C403 VDD2.n31 B 0.029807f
C404 VDD2.n32 B 0.013353f
C405 VDD2.n33 B 2.01948f
C406 VDD2.n34 B 0.012611f
C407 VDD2.t7 B 0.049518f
C408 VDD2.n35 B 0.180014f
C409 VDD2.n36 B 0.017608f
C410 VDD2.n37 B 0.022356f
C411 VDD2.n38 B 0.029807f
C412 VDD2.n39 B 0.013353f
C413 VDD2.n40 B 0.012611f
C414 VDD2.n41 B 0.023468f
C415 VDD2.n42 B 0.023468f
C416 VDD2.n43 B 0.012611f
C417 VDD2.n44 B 0.013353f
C418 VDD2.n45 B 0.029807f
C419 VDD2.n46 B 0.029807f
C420 VDD2.n47 B 0.013353f
C421 VDD2.n48 B 0.012611f
C422 VDD2.n49 B 0.023468f
C423 VDD2.n50 B 0.023468f
C424 VDD2.n51 B 0.012611f
C425 VDD2.n52 B 0.013353f
C426 VDD2.n53 B 0.029807f
C427 VDD2.n54 B 0.029807f
C428 VDD2.n55 B 0.013353f
C429 VDD2.n56 B 0.012611f
C430 VDD2.n57 B 0.023468f
C431 VDD2.n58 B 0.023468f
C432 VDD2.n59 B 0.012611f
C433 VDD2.n60 B 0.013353f
C434 VDD2.n61 B 0.029807f
C435 VDD2.n62 B 0.029807f
C436 VDD2.n63 B 0.013353f
C437 VDD2.n64 B 0.012611f
C438 VDD2.n65 B 0.023468f
C439 VDD2.n66 B 0.023468f
C440 VDD2.n67 B 0.012611f
C441 VDD2.n68 B 0.013353f
C442 VDD2.n69 B 0.029807f
C443 VDD2.n70 B 0.029807f
C444 VDD2.n71 B 0.013353f
C445 VDD2.n72 B 0.012611f
C446 VDD2.n73 B 0.023468f
C447 VDD2.n74 B 0.023468f
C448 VDD2.n75 B 0.012611f
C449 VDD2.n76 B 0.012611f
C450 VDD2.n77 B 0.013353f
C451 VDD2.n78 B 0.029807f
C452 VDD2.n79 B 0.029807f
C453 VDD2.n80 B 0.029807f
C454 VDD2.n81 B 0.012982f
C455 VDD2.n82 B 0.012611f
C456 VDD2.n83 B 0.023468f
C457 VDD2.n84 B 0.023468f
C458 VDD2.n85 B 0.012611f
C459 VDD2.n86 B 0.013353f
C460 VDD2.n87 B 0.029807f
C461 VDD2.n88 B 0.029807f
C462 VDD2.n89 B 0.013353f
C463 VDD2.n90 B 0.012611f
C464 VDD2.n91 B 0.023468f
C465 VDD2.n92 B 0.023468f
C466 VDD2.n93 B 0.012611f
C467 VDD2.n94 B 0.013353f
C468 VDD2.n95 B 0.029807f
C469 VDD2.n96 B 0.029807f
C470 VDD2.n97 B 0.013353f
C471 VDD2.n98 B 0.012611f
C472 VDD2.n99 B 0.023468f
C473 VDD2.n100 B 0.023468f
C474 VDD2.n101 B 0.012611f
C475 VDD2.n102 B 0.013353f
C476 VDD2.n103 B 0.029807f
C477 VDD2.n104 B 0.063968f
C478 VDD2.n105 B 0.013353f
C479 VDD2.n106 B 0.012611f
C480 VDD2.n107 B 0.05104f
C481 VDD2.n108 B 0.068773f
C482 VDD2.t3 B 0.363118f
C483 VDD2.t8 B 0.363118f
C484 VDD2.n109 B 3.31555f
C485 VDD2.n110 B 0.744483f
C486 VDD2.t4 B 0.363118f
C487 VDD2.t9 B 0.363118f
C488 VDD2.n111 B 3.33808f
C489 VDD2.n112 B 3.48847f
C490 VDD2.n113 B 0.03267f
C491 VDD2.n114 B 0.023468f
C492 VDD2.n115 B 0.012611f
C493 VDD2.n116 B 0.029807f
C494 VDD2.n117 B 0.013353f
C495 VDD2.n118 B 0.023468f
C496 VDD2.n119 B 0.012611f
C497 VDD2.n120 B 0.029807f
C498 VDD2.n121 B 0.013353f
C499 VDD2.n122 B 0.023468f
C500 VDD2.n123 B 0.012611f
C501 VDD2.n124 B 0.029807f
C502 VDD2.n125 B 0.012982f
C503 VDD2.n126 B 0.023468f
C504 VDD2.n127 B 0.012982f
C505 VDD2.n128 B 0.012611f
C506 VDD2.n129 B 0.029807f
C507 VDD2.n130 B 0.029807f
C508 VDD2.n131 B 0.013353f
C509 VDD2.n132 B 0.023468f
C510 VDD2.n133 B 0.012611f
C511 VDD2.n134 B 0.029807f
C512 VDD2.n135 B 0.013353f
C513 VDD2.n136 B 0.023468f
C514 VDD2.n137 B 0.012611f
C515 VDD2.n138 B 0.029807f
C516 VDD2.n139 B 0.013353f
C517 VDD2.n140 B 0.023468f
C518 VDD2.n141 B 0.012611f
C519 VDD2.n142 B 0.029807f
C520 VDD2.n143 B 0.013353f
C521 VDD2.n144 B 0.023468f
C522 VDD2.n145 B 0.012611f
C523 VDD2.n146 B 0.029807f
C524 VDD2.n147 B 0.013353f
C525 VDD2.n148 B 2.01948f
C526 VDD2.n149 B 0.012611f
C527 VDD2.t6 B 0.049518f
C528 VDD2.n150 B 0.180014f
C529 VDD2.n151 B 0.017608f
C530 VDD2.n152 B 0.022356f
C531 VDD2.n153 B 0.029807f
C532 VDD2.n154 B 0.013353f
C533 VDD2.n155 B 0.012611f
C534 VDD2.n156 B 0.023468f
C535 VDD2.n157 B 0.023468f
C536 VDD2.n158 B 0.012611f
C537 VDD2.n159 B 0.013353f
C538 VDD2.n160 B 0.029807f
C539 VDD2.n161 B 0.029807f
C540 VDD2.n162 B 0.013353f
C541 VDD2.n163 B 0.012611f
C542 VDD2.n164 B 0.023468f
C543 VDD2.n165 B 0.023468f
C544 VDD2.n166 B 0.012611f
C545 VDD2.n167 B 0.013353f
C546 VDD2.n168 B 0.029807f
C547 VDD2.n169 B 0.029807f
C548 VDD2.n170 B 0.013353f
C549 VDD2.n171 B 0.012611f
C550 VDD2.n172 B 0.023468f
C551 VDD2.n173 B 0.023468f
C552 VDD2.n174 B 0.012611f
C553 VDD2.n175 B 0.013353f
C554 VDD2.n176 B 0.029807f
C555 VDD2.n177 B 0.029807f
C556 VDD2.n178 B 0.013353f
C557 VDD2.n179 B 0.012611f
C558 VDD2.n180 B 0.023468f
C559 VDD2.n181 B 0.023468f
C560 VDD2.n182 B 0.012611f
C561 VDD2.n183 B 0.013353f
C562 VDD2.n184 B 0.029807f
C563 VDD2.n185 B 0.029807f
C564 VDD2.n186 B 0.013353f
C565 VDD2.n187 B 0.012611f
C566 VDD2.n188 B 0.023468f
C567 VDD2.n189 B 0.023468f
C568 VDD2.n190 B 0.012611f
C569 VDD2.n191 B 0.013353f
C570 VDD2.n192 B 0.029807f
C571 VDD2.n193 B 0.029807f
C572 VDD2.n194 B 0.013353f
C573 VDD2.n195 B 0.012611f
C574 VDD2.n196 B 0.023468f
C575 VDD2.n197 B 0.023468f
C576 VDD2.n198 B 0.012611f
C577 VDD2.n199 B 0.013353f
C578 VDD2.n200 B 0.029807f
C579 VDD2.n201 B 0.029807f
C580 VDD2.n202 B 0.013353f
C581 VDD2.n203 B 0.012611f
C582 VDD2.n204 B 0.023468f
C583 VDD2.n205 B 0.023468f
C584 VDD2.n206 B 0.012611f
C585 VDD2.n207 B 0.013353f
C586 VDD2.n208 B 0.029807f
C587 VDD2.n209 B 0.029807f
C588 VDD2.n210 B 0.013353f
C589 VDD2.n211 B 0.012611f
C590 VDD2.n212 B 0.023468f
C591 VDD2.n213 B 0.023468f
C592 VDD2.n214 B 0.012611f
C593 VDD2.n215 B 0.013353f
C594 VDD2.n216 B 0.029807f
C595 VDD2.n217 B 0.063968f
C596 VDD2.n218 B 0.013353f
C597 VDD2.n219 B 0.012611f
C598 VDD2.n220 B 0.05104f
C599 VDD2.n221 B 0.051865f
C600 VDD2.n222 B 3.48164f
C601 VDD2.t5 B 0.363118f
C602 VDD2.t0 B 0.363118f
C603 VDD2.n223 B 3.31556f
C604 VDD2.n224 B 0.493772f
C605 VDD2.t1 B 0.363118f
C606 VDD2.t2 B 0.363118f
C607 VDD2.n225 B 3.33804f
C608 VTAIL.t12 B 0.366773f
C609 VTAIL.t19 B 0.366773f
C610 VTAIL.n0 B 3.27075f
C611 VTAIL.n1 B 0.580595f
C612 VTAIL.n2 B 0.032999f
C613 VTAIL.n3 B 0.023704f
C614 VTAIL.n4 B 0.012738f
C615 VTAIL.n5 B 0.030108f
C616 VTAIL.n6 B 0.013487f
C617 VTAIL.n7 B 0.023704f
C618 VTAIL.n8 B 0.012738f
C619 VTAIL.n9 B 0.030108f
C620 VTAIL.n10 B 0.013487f
C621 VTAIL.n11 B 0.023704f
C622 VTAIL.n12 B 0.012738f
C623 VTAIL.n13 B 0.030108f
C624 VTAIL.n14 B 0.013112f
C625 VTAIL.n15 B 0.023704f
C626 VTAIL.n16 B 0.013487f
C627 VTAIL.n17 B 0.030108f
C628 VTAIL.n18 B 0.013487f
C629 VTAIL.n19 B 0.023704f
C630 VTAIL.n20 B 0.012738f
C631 VTAIL.n21 B 0.030108f
C632 VTAIL.n22 B 0.013487f
C633 VTAIL.n23 B 0.023704f
C634 VTAIL.n24 B 0.012738f
C635 VTAIL.n25 B 0.030108f
C636 VTAIL.n26 B 0.013487f
C637 VTAIL.n27 B 0.023704f
C638 VTAIL.n28 B 0.012738f
C639 VTAIL.n29 B 0.030108f
C640 VTAIL.n30 B 0.013487f
C641 VTAIL.n31 B 0.023704f
C642 VTAIL.n32 B 0.012738f
C643 VTAIL.n33 B 0.030108f
C644 VTAIL.n34 B 0.013487f
C645 VTAIL.n35 B 2.03981f
C646 VTAIL.n36 B 0.012738f
C647 VTAIL.t3 B 0.050016f
C648 VTAIL.n37 B 0.181826f
C649 VTAIL.n38 B 0.017785f
C650 VTAIL.n39 B 0.022581f
C651 VTAIL.n40 B 0.030108f
C652 VTAIL.n41 B 0.013487f
C653 VTAIL.n42 B 0.012738f
C654 VTAIL.n43 B 0.023704f
C655 VTAIL.n44 B 0.023704f
C656 VTAIL.n45 B 0.012738f
C657 VTAIL.n46 B 0.013487f
C658 VTAIL.n47 B 0.030108f
C659 VTAIL.n48 B 0.030108f
C660 VTAIL.n49 B 0.013487f
C661 VTAIL.n50 B 0.012738f
C662 VTAIL.n51 B 0.023704f
C663 VTAIL.n52 B 0.023704f
C664 VTAIL.n53 B 0.012738f
C665 VTAIL.n54 B 0.013487f
C666 VTAIL.n55 B 0.030108f
C667 VTAIL.n56 B 0.030108f
C668 VTAIL.n57 B 0.013487f
C669 VTAIL.n58 B 0.012738f
C670 VTAIL.n59 B 0.023704f
C671 VTAIL.n60 B 0.023704f
C672 VTAIL.n61 B 0.012738f
C673 VTAIL.n62 B 0.013487f
C674 VTAIL.n63 B 0.030108f
C675 VTAIL.n64 B 0.030108f
C676 VTAIL.n65 B 0.013487f
C677 VTAIL.n66 B 0.012738f
C678 VTAIL.n67 B 0.023704f
C679 VTAIL.n68 B 0.023704f
C680 VTAIL.n69 B 0.012738f
C681 VTAIL.n70 B 0.013487f
C682 VTAIL.n71 B 0.030108f
C683 VTAIL.n72 B 0.030108f
C684 VTAIL.n73 B 0.013487f
C685 VTAIL.n74 B 0.012738f
C686 VTAIL.n75 B 0.023704f
C687 VTAIL.n76 B 0.023704f
C688 VTAIL.n77 B 0.012738f
C689 VTAIL.n78 B 0.012738f
C690 VTAIL.n79 B 0.013487f
C691 VTAIL.n80 B 0.030108f
C692 VTAIL.n81 B 0.030108f
C693 VTAIL.n82 B 0.030108f
C694 VTAIL.n83 B 0.013112f
C695 VTAIL.n84 B 0.012738f
C696 VTAIL.n85 B 0.023704f
C697 VTAIL.n86 B 0.023704f
C698 VTAIL.n87 B 0.012738f
C699 VTAIL.n88 B 0.013487f
C700 VTAIL.n89 B 0.030108f
C701 VTAIL.n90 B 0.030108f
C702 VTAIL.n91 B 0.013487f
C703 VTAIL.n92 B 0.012738f
C704 VTAIL.n93 B 0.023704f
C705 VTAIL.n94 B 0.023704f
C706 VTAIL.n95 B 0.012738f
C707 VTAIL.n96 B 0.013487f
C708 VTAIL.n97 B 0.030108f
C709 VTAIL.n98 B 0.030108f
C710 VTAIL.n99 B 0.013487f
C711 VTAIL.n100 B 0.012738f
C712 VTAIL.n101 B 0.023704f
C713 VTAIL.n102 B 0.023704f
C714 VTAIL.n103 B 0.012738f
C715 VTAIL.n104 B 0.013487f
C716 VTAIL.n105 B 0.030108f
C717 VTAIL.n106 B 0.064612f
C718 VTAIL.n107 B 0.013487f
C719 VTAIL.n108 B 0.012738f
C720 VTAIL.n109 B 0.051554f
C721 VTAIL.n110 B 0.035992f
C722 VTAIL.n111 B 0.405924f
C723 VTAIL.t8 B 0.366773f
C724 VTAIL.t5 B 0.366773f
C725 VTAIL.n112 B 3.27075f
C726 VTAIL.n113 B 0.716073f
C727 VTAIL.t4 B 0.366773f
C728 VTAIL.t0 B 0.366773f
C729 VTAIL.n114 B 3.27075f
C730 VTAIL.n115 B 2.56175f
C731 VTAIL.t18 B 0.366773f
C732 VTAIL.t10 B 0.366773f
C733 VTAIL.n116 B 3.27077f
C734 VTAIL.n117 B 2.56173f
C735 VTAIL.t16 B 0.366773f
C736 VTAIL.t15 B 0.366773f
C737 VTAIL.n118 B 3.27077f
C738 VTAIL.n119 B 0.716058f
C739 VTAIL.n120 B 0.032999f
C740 VTAIL.n121 B 0.023704f
C741 VTAIL.n122 B 0.012738f
C742 VTAIL.n123 B 0.030108f
C743 VTAIL.n124 B 0.013487f
C744 VTAIL.n125 B 0.023704f
C745 VTAIL.n126 B 0.012738f
C746 VTAIL.n127 B 0.030108f
C747 VTAIL.n128 B 0.013487f
C748 VTAIL.n129 B 0.023704f
C749 VTAIL.n130 B 0.012738f
C750 VTAIL.n131 B 0.030108f
C751 VTAIL.n132 B 0.013112f
C752 VTAIL.n133 B 0.023704f
C753 VTAIL.n134 B 0.013112f
C754 VTAIL.n135 B 0.012738f
C755 VTAIL.n136 B 0.030108f
C756 VTAIL.n137 B 0.030108f
C757 VTAIL.n138 B 0.013487f
C758 VTAIL.n139 B 0.023704f
C759 VTAIL.n140 B 0.012738f
C760 VTAIL.n141 B 0.030108f
C761 VTAIL.n142 B 0.013487f
C762 VTAIL.n143 B 0.023704f
C763 VTAIL.n144 B 0.012738f
C764 VTAIL.n145 B 0.030108f
C765 VTAIL.n146 B 0.013487f
C766 VTAIL.n147 B 0.023704f
C767 VTAIL.n148 B 0.012738f
C768 VTAIL.n149 B 0.030108f
C769 VTAIL.n150 B 0.013487f
C770 VTAIL.n151 B 0.023704f
C771 VTAIL.n152 B 0.012738f
C772 VTAIL.n153 B 0.030108f
C773 VTAIL.n154 B 0.013487f
C774 VTAIL.n155 B 2.03981f
C775 VTAIL.n156 B 0.012738f
C776 VTAIL.t13 B 0.050016f
C777 VTAIL.n157 B 0.181826f
C778 VTAIL.n158 B 0.017785f
C779 VTAIL.n159 B 0.022581f
C780 VTAIL.n160 B 0.030108f
C781 VTAIL.n161 B 0.013487f
C782 VTAIL.n162 B 0.012738f
C783 VTAIL.n163 B 0.023704f
C784 VTAIL.n164 B 0.023704f
C785 VTAIL.n165 B 0.012738f
C786 VTAIL.n166 B 0.013487f
C787 VTAIL.n167 B 0.030108f
C788 VTAIL.n168 B 0.030108f
C789 VTAIL.n169 B 0.013487f
C790 VTAIL.n170 B 0.012738f
C791 VTAIL.n171 B 0.023704f
C792 VTAIL.n172 B 0.023704f
C793 VTAIL.n173 B 0.012738f
C794 VTAIL.n174 B 0.013487f
C795 VTAIL.n175 B 0.030108f
C796 VTAIL.n176 B 0.030108f
C797 VTAIL.n177 B 0.013487f
C798 VTAIL.n178 B 0.012738f
C799 VTAIL.n179 B 0.023704f
C800 VTAIL.n180 B 0.023704f
C801 VTAIL.n181 B 0.012738f
C802 VTAIL.n182 B 0.013487f
C803 VTAIL.n183 B 0.030108f
C804 VTAIL.n184 B 0.030108f
C805 VTAIL.n185 B 0.013487f
C806 VTAIL.n186 B 0.012738f
C807 VTAIL.n187 B 0.023704f
C808 VTAIL.n188 B 0.023704f
C809 VTAIL.n189 B 0.012738f
C810 VTAIL.n190 B 0.013487f
C811 VTAIL.n191 B 0.030108f
C812 VTAIL.n192 B 0.030108f
C813 VTAIL.n193 B 0.013487f
C814 VTAIL.n194 B 0.012738f
C815 VTAIL.n195 B 0.023704f
C816 VTAIL.n196 B 0.023704f
C817 VTAIL.n197 B 0.012738f
C818 VTAIL.n198 B 0.013487f
C819 VTAIL.n199 B 0.030108f
C820 VTAIL.n200 B 0.030108f
C821 VTAIL.n201 B 0.013487f
C822 VTAIL.n202 B 0.012738f
C823 VTAIL.n203 B 0.023704f
C824 VTAIL.n204 B 0.023704f
C825 VTAIL.n205 B 0.012738f
C826 VTAIL.n206 B 0.013487f
C827 VTAIL.n207 B 0.030108f
C828 VTAIL.n208 B 0.030108f
C829 VTAIL.n209 B 0.013487f
C830 VTAIL.n210 B 0.012738f
C831 VTAIL.n211 B 0.023704f
C832 VTAIL.n212 B 0.023704f
C833 VTAIL.n213 B 0.012738f
C834 VTAIL.n214 B 0.013487f
C835 VTAIL.n215 B 0.030108f
C836 VTAIL.n216 B 0.030108f
C837 VTAIL.n217 B 0.013487f
C838 VTAIL.n218 B 0.012738f
C839 VTAIL.n219 B 0.023704f
C840 VTAIL.n220 B 0.023704f
C841 VTAIL.n221 B 0.012738f
C842 VTAIL.n222 B 0.013487f
C843 VTAIL.n223 B 0.030108f
C844 VTAIL.n224 B 0.064612f
C845 VTAIL.n225 B 0.013487f
C846 VTAIL.n226 B 0.012738f
C847 VTAIL.n227 B 0.051554f
C848 VTAIL.n228 B 0.035992f
C849 VTAIL.n229 B 0.405924f
C850 VTAIL.t7 B 0.366773f
C851 VTAIL.t6 B 0.366773f
C852 VTAIL.n230 B 3.27077f
C853 VTAIL.n231 B 0.634739f
C854 VTAIL.t1 B 0.366773f
C855 VTAIL.t9 B 0.366773f
C856 VTAIL.n232 B 3.27077f
C857 VTAIL.n233 B 0.716058f
C858 VTAIL.n234 B 0.032999f
C859 VTAIL.n235 B 0.023704f
C860 VTAIL.n236 B 0.012738f
C861 VTAIL.n237 B 0.030108f
C862 VTAIL.n238 B 0.013487f
C863 VTAIL.n239 B 0.023704f
C864 VTAIL.n240 B 0.012738f
C865 VTAIL.n241 B 0.030108f
C866 VTAIL.n242 B 0.013487f
C867 VTAIL.n243 B 0.023704f
C868 VTAIL.n244 B 0.012738f
C869 VTAIL.n245 B 0.030108f
C870 VTAIL.n246 B 0.013112f
C871 VTAIL.n247 B 0.023704f
C872 VTAIL.n248 B 0.013112f
C873 VTAIL.n249 B 0.012738f
C874 VTAIL.n250 B 0.030108f
C875 VTAIL.n251 B 0.030108f
C876 VTAIL.n252 B 0.013487f
C877 VTAIL.n253 B 0.023704f
C878 VTAIL.n254 B 0.012738f
C879 VTAIL.n255 B 0.030108f
C880 VTAIL.n256 B 0.013487f
C881 VTAIL.n257 B 0.023704f
C882 VTAIL.n258 B 0.012738f
C883 VTAIL.n259 B 0.030108f
C884 VTAIL.n260 B 0.013487f
C885 VTAIL.n261 B 0.023704f
C886 VTAIL.n262 B 0.012738f
C887 VTAIL.n263 B 0.030108f
C888 VTAIL.n264 B 0.013487f
C889 VTAIL.n265 B 0.023704f
C890 VTAIL.n266 B 0.012738f
C891 VTAIL.n267 B 0.030108f
C892 VTAIL.n268 B 0.013487f
C893 VTAIL.n269 B 2.03981f
C894 VTAIL.n270 B 0.012738f
C895 VTAIL.t2 B 0.050016f
C896 VTAIL.n271 B 0.181826f
C897 VTAIL.n272 B 0.017785f
C898 VTAIL.n273 B 0.022581f
C899 VTAIL.n274 B 0.030108f
C900 VTAIL.n275 B 0.013487f
C901 VTAIL.n276 B 0.012738f
C902 VTAIL.n277 B 0.023704f
C903 VTAIL.n278 B 0.023704f
C904 VTAIL.n279 B 0.012738f
C905 VTAIL.n280 B 0.013487f
C906 VTAIL.n281 B 0.030108f
C907 VTAIL.n282 B 0.030108f
C908 VTAIL.n283 B 0.013487f
C909 VTAIL.n284 B 0.012738f
C910 VTAIL.n285 B 0.023704f
C911 VTAIL.n286 B 0.023704f
C912 VTAIL.n287 B 0.012738f
C913 VTAIL.n288 B 0.013487f
C914 VTAIL.n289 B 0.030108f
C915 VTAIL.n290 B 0.030108f
C916 VTAIL.n291 B 0.013487f
C917 VTAIL.n292 B 0.012738f
C918 VTAIL.n293 B 0.023704f
C919 VTAIL.n294 B 0.023704f
C920 VTAIL.n295 B 0.012738f
C921 VTAIL.n296 B 0.013487f
C922 VTAIL.n297 B 0.030108f
C923 VTAIL.n298 B 0.030108f
C924 VTAIL.n299 B 0.013487f
C925 VTAIL.n300 B 0.012738f
C926 VTAIL.n301 B 0.023704f
C927 VTAIL.n302 B 0.023704f
C928 VTAIL.n303 B 0.012738f
C929 VTAIL.n304 B 0.013487f
C930 VTAIL.n305 B 0.030108f
C931 VTAIL.n306 B 0.030108f
C932 VTAIL.n307 B 0.013487f
C933 VTAIL.n308 B 0.012738f
C934 VTAIL.n309 B 0.023704f
C935 VTAIL.n310 B 0.023704f
C936 VTAIL.n311 B 0.012738f
C937 VTAIL.n312 B 0.013487f
C938 VTAIL.n313 B 0.030108f
C939 VTAIL.n314 B 0.030108f
C940 VTAIL.n315 B 0.013487f
C941 VTAIL.n316 B 0.012738f
C942 VTAIL.n317 B 0.023704f
C943 VTAIL.n318 B 0.023704f
C944 VTAIL.n319 B 0.012738f
C945 VTAIL.n320 B 0.013487f
C946 VTAIL.n321 B 0.030108f
C947 VTAIL.n322 B 0.030108f
C948 VTAIL.n323 B 0.013487f
C949 VTAIL.n324 B 0.012738f
C950 VTAIL.n325 B 0.023704f
C951 VTAIL.n326 B 0.023704f
C952 VTAIL.n327 B 0.012738f
C953 VTAIL.n328 B 0.013487f
C954 VTAIL.n329 B 0.030108f
C955 VTAIL.n330 B 0.030108f
C956 VTAIL.n331 B 0.013487f
C957 VTAIL.n332 B 0.012738f
C958 VTAIL.n333 B 0.023704f
C959 VTAIL.n334 B 0.023704f
C960 VTAIL.n335 B 0.012738f
C961 VTAIL.n336 B 0.013487f
C962 VTAIL.n337 B 0.030108f
C963 VTAIL.n338 B 0.064612f
C964 VTAIL.n339 B 0.013487f
C965 VTAIL.n340 B 0.012738f
C966 VTAIL.n341 B 0.051554f
C967 VTAIL.n342 B 0.035992f
C968 VTAIL.n343 B 2.0985f
C969 VTAIL.n344 B 0.032999f
C970 VTAIL.n345 B 0.023704f
C971 VTAIL.n346 B 0.012738f
C972 VTAIL.n347 B 0.030108f
C973 VTAIL.n348 B 0.013487f
C974 VTAIL.n349 B 0.023704f
C975 VTAIL.n350 B 0.012738f
C976 VTAIL.n351 B 0.030108f
C977 VTAIL.n352 B 0.013487f
C978 VTAIL.n353 B 0.023704f
C979 VTAIL.n354 B 0.012738f
C980 VTAIL.n355 B 0.030108f
C981 VTAIL.n356 B 0.013112f
C982 VTAIL.n357 B 0.023704f
C983 VTAIL.n358 B 0.013487f
C984 VTAIL.n359 B 0.030108f
C985 VTAIL.n360 B 0.013487f
C986 VTAIL.n361 B 0.023704f
C987 VTAIL.n362 B 0.012738f
C988 VTAIL.n363 B 0.030108f
C989 VTAIL.n364 B 0.013487f
C990 VTAIL.n365 B 0.023704f
C991 VTAIL.n366 B 0.012738f
C992 VTAIL.n367 B 0.030108f
C993 VTAIL.n368 B 0.013487f
C994 VTAIL.n369 B 0.023704f
C995 VTAIL.n370 B 0.012738f
C996 VTAIL.n371 B 0.030108f
C997 VTAIL.n372 B 0.013487f
C998 VTAIL.n373 B 0.023704f
C999 VTAIL.n374 B 0.012738f
C1000 VTAIL.n375 B 0.030108f
C1001 VTAIL.n376 B 0.013487f
C1002 VTAIL.n377 B 2.03981f
C1003 VTAIL.n378 B 0.012738f
C1004 VTAIL.t17 B 0.050016f
C1005 VTAIL.n379 B 0.181826f
C1006 VTAIL.n380 B 0.017785f
C1007 VTAIL.n381 B 0.022581f
C1008 VTAIL.n382 B 0.030108f
C1009 VTAIL.n383 B 0.013487f
C1010 VTAIL.n384 B 0.012738f
C1011 VTAIL.n385 B 0.023704f
C1012 VTAIL.n386 B 0.023704f
C1013 VTAIL.n387 B 0.012738f
C1014 VTAIL.n388 B 0.013487f
C1015 VTAIL.n389 B 0.030108f
C1016 VTAIL.n390 B 0.030108f
C1017 VTAIL.n391 B 0.013487f
C1018 VTAIL.n392 B 0.012738f
C1019 VTAIL.n393 B 0.023704f
C1020 VTAIL.n394 B 0.023704f
C1021 VTAIL.n395 B 0.012738f
C1022 VTAIL.n396 B 0.013487f
C1023 VTAIL.n397 B 0.030108f
C1024 VTAIL.n398 B 0.030108f
C1025 VTAIL.n399 B 0.013487f
C1026 VTAIL.n400 B 0.012738f
C1027 VTAIL.n401 B 0.023704f
C1028 VTAIL.n402 B 0.023704f
C1029 VTAIL.n403 B 0.012738f
C1030 VTAIL.n404 B 0.013487f
C1031 VTAIL.n405 B 0.030108f
C1032 VTAIL.n406 B 0.030108f
C1033 VTAIL.n407 B 0.013487f
C1034 VTAIL.n408 B 0.012738f
C1035 VTAIL.n409 B 0.023704f
C1036 VTAIL.n410 B 0.023704f
C1037 VTAIL.n411 B 0.012738f
C1038 VTAIL.n412 B 0.013487f
C1039 VTAIL.n413 B 0.030108f
C1040 VTAIL.n414 B 0.030108f
C1041 VTAIL.n415 B 0.013487f
C1042 VTAIL.n416 B 0.012738f
C1043 VTAIL.n417 B 0.023704f
C1044 VTAIL.n418 B 0.023704f
C1045 VTAIL.n419 B 0.012738f
C1046 VTAIL.n420 B 0.012738f
C1047 VTAIL.n421 B 0.013487f
C1048 VTAIL.n422 B 0.030108f
C1049 VTAIL.n423 B 0.030108f
C1050 VTAIL.n424 B 0.030108f
C1051 VTAIL.n425 B 0.013112f
C1052 VTAIL.n426 B 0.012738f
C1053 VTAIL.n427 B 0.023704f
C1054 VTAIL.n428 B 0.023704f
C1055 VTAIL.n429 B 0.012738f
C1056 VTAIL.n430 B 0.013487f
C1057 VTAIL.n431 B 0.030108f
C1058 VTAIL.n432 B 0.030108f
C1059 VTAIL.n433 B 0.013487f
C1060 VTAIL.n434 B 0.012738f
C1061 VTAIL.n435 B 0.023704f
C1062 VTAIL.n436 B 0.023704f
C1063 VTAIL.n437 B 0.012738f
C1064 VTAIL.n438 B 0.013487f
C1065 VTAIL.n439 B 0.030108f
C1066 VTAIL.n440 B 0.030108f
C1067 VTAIL.n441 B 0.013487f
C1068 VTAIL.n442 B 0.012738f
C1069 VTAIL.n443 B 0.023704f
C1070 VTAIL.n444 B 0.023704f
C1071 VTAIL.n445 B 0.012738f
C1072 VTAIL.n446 B 0.013487f
C1073 VTAIL.n447 B 0.030108f
C1074 VTAIL.n448 B 0.064612f
C1075 VTAIL.n449 B 0.013487f
C1076 VTAIL.n450 B 0.012738f
C1077 VTAIL.n451 B 0.051554f
C1078 VTAIL.n452 B 0.035992f
C1079 VTAIL.n453 B 2.0985f
C1080 VTAIL.t11 B 0.366773f
C1081 VTAIL.t14 B 0.366773f
C1082 VTAIL.n454 B 3.27075f
C1083 VTAIL.n455 B 0.53582f
C1084 VN.t0 B 3.05075f
C1085 VN.n0 B 1.12162f
C1086 VN.n1 B 0.017511f
C1087 VN.n2 B 0.016039f
C1088 VN.n3 B 0.017511f
C1089 VN.t5 B 3.05075f
C1090 VN.n4 B 1.05056f
C1091 VN.n5 B 0.017511f
C1092 VN.n6 B 0.014345f
C1093 VN.n7 B 0.017511f
C1094 VN.t1 B 3.05075f
C1095 VN.n8 B 1.05056f
C1096 VN.n9 B 0.017511f
C1097 VN.n10 B 0.014345f
C1098 VN.n11 B 0.017511f
C1099 VN.t6 B 3.05075f
C1100 VN.n12 B 1.10987f
C1101 VN.t2 B 3.26934f
C1102 VN.n13 B 1.06715f
C1103 VN.n14 B 0.202977f
C1104 VN.n15 B 0.026381f
C1105 VN.n16 B 0.032472f
C1106 VN.n17 B 0.034004f
C1107 VN.n18 B 0.017511f
C1108 VN.n19 B 0.017511f
C1109 VN.n20 B 0.017511f
C1110 VN.n21 B 0.035032f
C1111 VN.n22 B 0.032472f
C1112 VN.n23 B 0.024457f
C1113 VN.n24 B 0.017511f
C1114 VN.n25 B 0.017511f
C1115 VN.n26 B 0.024457f
C1116 VN.n27 B 0.032472f
C1117 VN.n28 B 0.035032f
C1118 VN.n29 B 0.017511f
C1119 VN.n30 B 0.017511f
C1120 VN.n31 B 0.017511f
C1121 VN.n32 B 0.034004f
C1122 VN.n33 B 0.032472f
C1123 VN.n34 B 0.026381f
C1124 VN.n35 B 0.017511f
C1125 VN.n36 B 0.017511f
C1126 VN.n37 B 0.022533f
C1127 VN.n38 B 0.032472f
C1128 VN.n39 B 0.035032f
C1129 VN.n40 B 0.017511f
C1130 VN.n41 B 0.017511f
C1131 VN.n42 B 0.017511f
C1132 VN.n43 B 0.032312f
C1133 VN.n44 B 0.032472f
C1134 VN.n45 B 0.028304f
C1135 VN.n46 B 0.028258f
C1136 VN.n47 B 0.039301f
C1137 VN.t3 B 3.05075f
C1138 VN.n48 B 1.12162f
C1139 VN.n49 B 0.017511f
C1140 VN.n50 B 0.016039f
C1141 VN.n51 B 0.017511f
C1142 VN.t4 B 3.05075f
C1143 VN.n52 B 1.05056f
C1144 VN.n53 B 0.017511f
C1145 VN.n54 B 0.014345f
C1146 VN.n55 B 0.017511f
C1147 VN.t9 B 3.05075f
C1148 VN.n56 B 1.05056f
C1149 VN.n57 B 0.017511f
C1150 VN.n58 B 0.014345f
C1151 VN.n59 B 0.017511f
C1152 VN.t8 B 3.05075f
C1153 VN.n60 B 1.10987f
C1154 VN.t7 B 3.26934f
C1155 VN.n61 B 1.06715f
C1156 VN.n62 B 0.202977f
C1157 VN.n63 B 0.026381f
C1158 VN.n64 B 0.032472f
C1159 VN.n65 B 0.034004f
C1160 VN.n66 B 0.017511f
C1161 VN.n67 B 0.017511f
C1162 VN.n68 B 0.017511f
C1163 VN.n69 B 0.035032f
C1164 VN.n70 B 0.032472f
C1165 VN.n71 B 0.024457f
C1166 VN.n72 B 0.017511f
C1167 VN.n73 B 0.017511f
C1168 VN.n74 B 0.024457f
C1169 VN.n75 B 0.032472f
C1170 VN.n76 B 0.035032f
C1171 VN.n77 B 0.017511f
C1172 VN.n78 B 0.017511f
C1173 VN.n79 B 0.017511f
C1174 VN.n80 B 0.034004f
C1175 VN.n81 B 0.032472f
C1176 VN.n82 B 0.026381f
C1177 VN.n83 B 0.017511f
C1178 VN.n84 B 0.017511f
C1179 VN.n85 B 0.022533f
C1180 VN.n86 B 0.032472f
C1181 VN.n87 B 0.035032f
C1182 VN.n88 B 0.017511f
C1183 VN.n89 B 0.017511f
C1184 VN.n90 B 0.017511f
C1185 VN.n91 B 0.032312f
C1186 VN.n92 B 0.032472f
C1187 VN.n93 B 0.028304f
C1188 VN.n94 B 0.028258f
C1189 VN.n95 B 1.35579f
.ends

