* NGSPICE file created from diff_pair_sample_1268.ext - technology: sky130A

.subckt diff_pair_sample_1268 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t15 VP.t0 VDD1.t4 w_n5290_n2572# sky130_fd_pr__pfet_01v8 ad=1.3233 pd=8.35 as=1.3233 ps=8.35 w=8.02 l=3.99
X1 VTAIL.t6 VN.t0 VDD2.t7 w_n5290_n2572# sky130_fd_pr__pfet_01v8 ad=3.1278 pd=16.82 as=1.3233 ps=8.35 w=8.02 l=3.99
X2 VTAIL.t0 VN.t1 VDD2.t6 w_n5290_n2572# sky130_fd_pr__pfet_01v8 ad=1.3233 pd=8.35 as=1.3233 ps=8.35 w=8.02 l=3.99
X3 B.t11 B.t9 B.t10 w_n5290_n2572# sky130_fd_pr__pfet_01v8 ad=3.1278 pd=16.82 as=0 ps=0 w=8.02 l=3.99
X4 VDD2.t5 VN.t2 VTAIL.t5 w_n5290_n2572# sky130_fd_pr__pfet_01v8 ad=1.3233 pd=8.35 as=1.3233 ps=8.35 w=8.02 l=3.99
X5 B.t8 B.t6 B.t7 w_n5290_n2572# sky130_fd_pr__pfet_01v8 ad=3.1278 pd=16.82 as=0 ps=0 w=8.02 l=3.99
X6 VTAIL.t14 VP.t1 VDD1.t5 w_n5290_n2572# sky130_fd_pr__pfet_01v8 ad=1.3233 pd=8.35 as=1.3233 ps=8.35 w=8.02 l=3.99
X7 VDD2.t4 VN.t3 VTAIL.t7 w_n5290_n2572# sky130_fd_pr__pfet_01v8 ad=1.3233 pd=8.35 as=3.1278 ps=16.82 w=8.02 l=3.99
X8 B.t5 B.t3 B.t4 w_n5290_n2572# sky130_fd_pr__pfet_01v8 ad=3.1278 pd=16.82 as=0 ps=0 w=8.02 l=3.99
X9 B.t2 B.t0 B.t1 w_n5290_n2572# sky130_fd_pr__pfet_01v8 ad=3.1278 pd=16.82 as=0 ps=0 w=8.02 l=3.99
X10 VDD1.t7 VP.t2 VTAIL.t13 w_n5290_n2572# sky130_fd_pr__pfet_01v8 ad=1.3233 pd=8.35 as=1.3233 ps=8.35 w=8.02 l=3.99
X11 VDD1.t6 VP.t3 VTAIL.t12 w_n5290_n2572# sky130_fd_pr__pfet_01v8 ad=1.3233 pd=8.35 as=3.1278 ps=16.82 w=8.02 l=3.99
X12 VTAIL.t11 VP.t4 VDD1.t2 w_n5290_n2572# sky130_fd_pr__pfet_01v8 ad=3.1278 pd=16.82 as=1.3233 ps=8.35 w=8.02 l=3.99
X13 VTAIL.t4 VN.t4 VDD2.t3 w_n5290_n2572# sky130_fd_pr__pfet_01v8 ad=1.3233 pd=8.35 as=1.3233 ps=8.35 w=8.02 l=3.99
X14 VTAIL.t10 VP.t5 VDD1.t0 w_n5290_n2572# sky130_fd_pr__pfet_01v8 ad=3.1278 pd=16.82 as=1.3233 ps=8.35 w=8.02 l=3.99
X15 VDD2.t2 VN.t5 VTAIL.t3 w_n5290_n2572# sky130_fd_pr__pfet_01v8 ad=1.3233 pd=8.35 as=1.3233 ps=8.35 w=8.02 l=3.99
X16 VDD1.t1 VP.t6 VTAIL.t9 w_n5290_n2572# sky130_fd_pr__pfet_01v8 ad=1.3233 pd=8.35 as=1.3233 ps=8.35 w=8.02 l=3.99
X17 VDD2.t1 VN.t6 VTAIL.t2 w_n5290_n2572# sky130_fd_pr__pfet_01v8 ad=1.3233 pd=8.35 as=3.1278 ps=16.82 w=8.02 l=3.99
X18 VDD1.t3 VP.t7 VTAIL.t8 w_n5290_n2572# sky130_fd_pr__pfet_01v8 ad=1.3233 pd=8.35 as=3.1278 ps=16.82 w=8.02 l=3.99
X19 VTAIL.t1 VN.t7 VDD2.t0 w_n5290_n2572# sky130_fd_pr__pfet_01v8 ad=3.1278 pd=16.82 as=1.3233 ps=8.35 w=8.02 l=3.99
R0 VP.n24 VP.n21 161.3
R1 VP.n26 VP.n25 161.3
R2 VP.n27 VP.n20 161.3
R3 VP.n29 VP.n28 161.3
R4 VP.n30 VP.n19 161.3
R5 VP.n32 VP.n31 161.3
R6 VP.n33 VP.n18 161.3
R7 VP.n35 VP.n34 161.3
R8 VP.n36 VP.n17 161.3
R9 VP.n39 VP.n38 161.3
R10 VP.n40 VP.n16 161.3
R11 VP.n42 VP.n41 161.3
R12 VP.n43 VP.n15 161.3
R13 VP.n45 VP.n44 161.3
R14 VP.n46 VP.n14 161.3
R15 VP.n48 VP.n47 161.3
R16 VP.n49 VP.n13 161.3
R17 VP.n92 VP.n0 161.3
R18 VP.n91 VP.n90 161.3
R19 VP.n89 VP.n1 161.3
R20 VP.n88 VP.n87 161.3
R21 VP.n86 VP.n2 161.3
R22 VP.n85 VP.n84 161.3
R23 VP.n83 VP.n3 161.3
R24 VP.n82 VP.n81 161.3
R25 VP.n79 VP.n4 161.3
R26 VP.n78 VP.n77 161.3
R27 VP.n76 VP.n5 161.3
R28 VP.n75 VP.n74 161.3
R29 VP.n73 VP.n6 161.3
R30 VP.n72 VP.n71 161.3
R31 VP.n70 VP.n7 161.3
R32 VP.n69 VP.n68 161.3
R33 VP.n67 VP.n8 161.3
R34 VP.n65 VP.n64 161.3
R35 VP.n63 VP.n9 161.3
R36 VP.n62 VP.n61 161.3
R37 VP.n60 VP.n10 161.3
R38 VP.n59 VP.n58 161.3
R39 VP.n57 VP.n11 161.3
R40 VP.n56 VP.n55 161.3
R41 VP.n54 VP.n12 161.3
R42 VP.n22 VP.t5 80.565
R43 VP.n23 VP.n22 67.5408
R44 VP.n53 VP.n52 58.7717
R45 VP.n94 VP.n93 58.7717
R46 VP.n51 VP.n50 58.7717
R47 VP.n60 VP.n59 56.5617
R48 VP.n87 VP.n86 56.5617
R49 VP.n44 VP.n43 56.5617
R50 VP.n52 VP.n51 54.6787
R51 VP.n53 VP.t4 48.4421
R52 VP.n66 VP.t6 48.4421
R53 VP.n80 VP.t1 48.4421
R54 VP.n93 VP.t3 48.4421
R55 VP.n50 VP.t7 48.4421
R56 VP.n37 VP.t0 48.4421
R57 VP.n23 VP.t2 48.4421
R58 VP.n73 VP.n72 40.577
R59 VP.n74 VP.n73 40.577
R60 VP.n31 VP.n30 40.577
R61 VP.n30 VP.n29 40.577
R62 VP.n55 VP.n54 24.5923
R63 VP.n55 VP.n11 24.5923
R64 VP.n59 VP.n11 24.5923
R65 VP.n61 VP.n60 24.5923
R66 VP.n61 VP.n9 24.5923
R67 VP.n65 VP.n9 24.5923
R68 VP.n68 VP.n67 24.5923
R69 VP.n68 VP.n7 24.5923
R70 VP.n72 VP.n7 24.5923
R71 VP.n74 VP.n5 24.5923
R72 VP.n78 VP.n5 24.5923
R73 VP.n79 VP.n78 24.5923
R74 VP.n81 VP.n3 24.5923
R75 VP.n85 VP.n3 24.5923
R76 VP.n86 VP.n85 24.5923
R77 VP.n87 VP.n1 24.5923
R78 VP.n91 VP.n1 24.5923
R79 VP.n92 VP.n91 24.5923
R80 VP.n44 VP.n14 24.5923
R81 VP.n48 VP.n14 24.5923
R82 VP.n49 VP.n48 24.5923
R83 VP.n31 VP.n18 24.5923
R84 VP.n35 VP.n18 24.5923
R85 VP.n36 VP.n35 24.5923
R86 VP.n38 VP.n16 24.5923
R87 VP.n42 VP.n16 24.5923
R88 VP.n43 VP.n42 24.5923
R89 VP.n25 VP.n24 24.5923
R90 VP.n25 VP.n20 24.5923
R91 VP.n29 VP.n20 24.5923
R92 VP.n54 VP.n53 23.6087
R93 VP.n93 VP.n92 23.6087
R94 VP.n50 VP.n49 23.6087
R95 VP.n66 VP.n65 16.7229
R96 VP.n81 VP.n80 16.7229
R97 VP.n38 VP.n37 16.7229
R98 VP.n67 VP.n66 7.86989
R99 VP.n80 VP.n79 7.86989
R100 VP.n37 VP.n36 7.86989
R101 VP.n24 VP.n23 7.86989
R102 VP.n22 VP.n21 2.56251
R103 VP.n51 VP.n13 0.417304
R104 VP.n52 VP.n12 0.417304
R105 VP.n94 VP.n0 0.417304
R106 VP VP.n94 0.394524
R107 VP.n26 VP.n21 0.189894
R108 VP.n27 VP.n26 0.189894
R109 VP.n28 VP.n27 0.189894
R110 VP.n28 VP.n19 0.189894
R111 VP.n32 VP.n19 0.189894
R112 VP.n33 VP.n32 0.189894
R113 VP.n34 VP.n33 0.189894
R114 VP.n34 VP.n17 0.189894
R115 VP.n39 VP.n17 0.189894
R116 VP.n40 VP.n39 0.189894
R117 VP.n41 VP.n40 0.189894
R118 VP.n41 VP.n15 0.189894
R119 VP.n45 VP.n15 0.189894
R120 VP.n46 VP.n45 0.189894
R121 VP.n47 VP.n46 0.189894
R122 VP.n47 VP.n13 0.189894
R123 VP.n56 VP.n12 0.189894
R124 VP.n57 VP.n56 0.189894
R125 VP.n58 VP.n57 0.189894
R126 VP.n58 VP.n10 0.189894
R127 VP.n62 VP.n10 0.189894
R128 VP.n63 VP.n62 0.189894
R129 VP.n64 VP.n63 0.189894
R130 VP.n64 VP.n8 0.189894
R131 VP.n69 VP.n8 0.189894
R132 VP.n70 VP.n69 0.189894
R133 VP.n71 VP.n70 0.189894
R134 VP.n71 VP.n6 0.189894
R135 VP.n75 VP.n6 0.189894
R136 VP.n76 VP.n75 0.189894
R137 VP.n77 VP.n76 0.189894
R138 VP.n77 VP.n4 0.189894
R139 VP.n82 VP.n4 0.189894
R140 VP.n83 VP.n82 0.189894
R141 VP.n84 VP.n83 0.189894
R142 VP.n84 VP.n2 0.189894
R143 VP.n88 VP.n2 0.189894
R144 VP.n89 VP.n88 0.189894
R145 VP.n90 VP.n89 0.189894
R146 VP.n90 VP.n0 0.189894
R147 VDD1 VDD1.n0 88.5462
R148 VDD1.n3 VDD1.n2 88.4325
R149 VDD1.n3 VDD1.n1 88.4325
R150 VDD1.n5 VDD1.n4 86.6257
R151 VDD1.n5 VDD1.n3 47.9707
R152 VDD1.n4 VDD1.t4 4.05349
R153 VDD1.n4 VDD1.t3 4.05349
R154 VDD1.n0 VDD1.t0 4.05349
R155 VDD1.n0 VDD1.t7 4.05349
R156 VDD1.n2 VDD1.t5 4.05349
R157 VDD1.n2 VDD1.t6 4.05349
R158 VDD1.n1 VDD1.t2 4.05349
R159 VDD1.n1 VDD1.t1 4.05349
R160 VDD1 VDD1.n5 1.80438
R161 VTAIL.n338 VTAIL.n302 756.745
R162 VTAIL.n38 VTAIL.n2 756.745
R163 VTAIL.n80 VTAIL.n44 756.745
R164 VTAIL.n124 VTAIL.n88 756.745
R165 VTAIL.n296 VTAIL.n260 756.745
R166 VTAIL.n252 VTAIL.n216 756.745
R167 VTAIL.n210 VTAIL.n174 756.745
R168 VTAIL.n166 VTAIL.n130 756.745
R169 VTAIL.n314 VTAIL.n313 585
R170 VTAIL.n319 VTAIL.n318 585
R171 VTAIL.n321 VTAIL.n320 585
R172 VTAIL.n310 VTAIL.n309 585
R173 VTAIL.n327 VTAIL.n326 585
R174 VTAIL.n329 VTAIL.n328 585
R175 VTAIL.n306 VTAIL.n305 585
R176 VTAIL.n336 VTAIL.n335 585
R177 VTAIL.n337 VTAIL.n304 585
R178 VTAIL.n339 VTAIL.n338 585
R179 VTAIL.n14 VTAIL.n13 585
R180 VTAIL.n19 VTAIL.n18 585
R181 VTAIL.n21 VTAIL.n20 585
R182 VTAIL.n10 VTAIL.n9 585
R183 VTAIL.n27 VTAIL.n26 585
R184 VTAIL.n29 VTAIL.n28 585
R185 VTAIL.n6 VTAIL.n5 585
R186 VTAIL.n36 VTAIL.n35 585
R187 VTAIL.n37 VTAIL.n4 585
R188 VTAIL.n39 VTAIL.n38 585
R189 VTAIL.n56 VTAIL.n55 585
R190 VTAIL.n61 VTAIL.n60 585
R191 VTAIL.n63 VTAIL.n62 585
R192 VTAIL.n52 VTAIL.n51 585
R193 VTAIL.n69 VTAIL.n68 585
R194 VTAIL.n71 VTAIL.n70 585
R195 VTAIL.n48 VTAIL.n47 585
R196 VTAIL.n78 VTAIL.n77 585
R197 VTAIL.n79 VTAIL.n46 585
R198 VTAIL.n81 VTAIL.n80 585
R199 VTAIL.n100 VTAIL.n99 585
R200 VTAIL.n105 VTAIL.n104 585
R201 VTAIL.n107 VTAIL.n106 585
R202 VTAIL.n96 VTAIL.n95 585
R203 VTAIL.n113 VTAIL.n112 585
R204 VTAIL.n115 VTAIL.n114 585
R205 VTAIL.n92 VTAIL.n91 585
R206 VTAIL.n122 VTAIL.n121 585
R207 VTAIL.n123 VTAIL.n90 585
R208 VTAIL.n125 VTAIL.n124 585
R209 VTAIL.n297 VTAIL.n296 585
R210 VTAIL.n295 VTAIL.n262 585
R211 VTAIL.n294 VTAIL.n293 585
R212 VTAIL.n265 VTAIL.n263 585
R213 VTAIL.n288 VTAIL.n287 585
R214 VTAIL.n286 VTAIL.n285 585
R215 VTAIL.n269 VTAIL.n268 585
R216 VTAIL.n280 VTAIL.n279 585
R217 VTAIL.n278 VTAIL.n277 585
R218 VTAIL.n273 VTAIL.n272 585
R219 VTAIL.n253 VTAIL.n252 585
R220 VTAIL.n251 VTAIL.n218 585
R221 VTAIL.n250 VTAIL.n249 585
R222 VTAIL.n221 VTAIL.n219 585
R223 VTAIL.n244 VTAIL.n243 585
R224 VTAIL.n242 VTAIL.n241 585
R225 VTAIL.n225 VTAIL.n224 585
R226 VTAIL.n236 VTAIL.n235 585
R227 VTAIL.n234 VTAIL.n233 585
R228 VTAIL.n229 VTAIL.n228 585
R229 VTAIL.n211 VTAIL.n210 585
R230 VTAIL.n209 VTAIL.n176 585
R231 VTAIL.n208 VTAIL.n207 585
R232 VTAIL.n179 VTAIL.n177 585
R233 VTAIL.n202 VTAIL.n201 585
R234 VTAIL.n200 VTAIL.n199 585
R235 VTAIL.n183 VTAIL.n182 585
R236 VTAIL.n194 VTAIL.n193 585
R237 VTAIL.n192 VTAIL.n191 585
R238 VTAIL.n187 VTAIL.n186 585
R239 VTAIL.n167 VTAIL.n166 585
R240 VTAIL.n165 VTAIL.n132 585
R241 VTAIL.n164 VTAIL.n163 585
R242 VTAIL.n135 VTAIL.n133 585
R243 VTAIL.n158 VTAIL.n157 585
R244 VTAIL.n156 VTAIL.n155 585
R245 VTAIL.n139 VTAIL.n138 585
R246 VTAIL.n150 VTAIL.n149 585
R247 VTAIL.n148 VTAIL.n147 585
R248 VTAIL.n143 VTAIL.n142 585
R249 VTAIL.n315 VTAIL.t2 329.043
R250 VTAIL.n15 VTAIL.t1 329.043
R251 VTAIL.n57 VTAIL.t12 329.043
R252 VTAIL.n101 VTAIL.t11 329.043
R253 VTAIL.n274 VTAIL.t8 329.043
R254 VTAIL.n230 VTAIL.t10 329.043
R255 VTAIL.n188 VTAIL.t7 329.043
R256 VTAIL.n144 VTAIL.t6 329.043
R257 VTAIL.n319 VTAIL.n313 171.744
R258 VTAIL.n320 VTAIL.n319 171.744
R259 VTAIL.n320 VTAIL.n309 171.744
R260 VTAIL.n327 VTAIL.n309 171.744
R261 VTAIL.n328 VTAIL.n327 171.744
R262 VTAIL.n328 VTAIL.n305 171.744
R263 VTAIL.n336 VTAIL.n305 171.744
R264 VTAIL.n337 VTAIL.n336 171.744
R265 VTAIL.n338 VTAIL.n337 171.744
R266 VTAIL.n19 VTAIL.n13 171.744
R267 VTAIL.n20 VTAIL.n19 171.744
R268 VTAIL.n20 VTAIL.n9 171.744
R269 VTAIL.n27 VTAIL.n9 171.744
R270 VTAIL.n28 VTAIL.n27 171.744
R271 VTAIL.n28 VTAIL.n5 171.744
R272 VTAIL.n36 VTAIL.n5 171.744
R273 VTAIL.n37 VTAIL.n36 171.744
R274 VTAIL.n38 VTAIL.n37 171.744
R275 VTAIL.n61 VTAIL.n55 171.744
R276 VTAIL.n62 VTAIL.n61 171.744
R277 VTAIL.n62 VTAIL.n51 171.744
R278 VTAIL.n69 VTAIL.n51 171.744
R279 VTAIL.n70 VTAIL.n69 171.744
R280 VTAIL.n70 VTAIL.n47 171.744
R281 VTAIL.n78 VTAIL.n47 171.744
R282 VTAIL.n79 VTAIL.n78 171.744
R283 VTAIL.n80 VTAIL.n79 171.744
R284 VTAIL.n105 VTAIL.n99 171.744
R285 VTAIL.n106 VTAIL.n105 171.744
R286 VTAIL.n106 VTAIL.n95 171.744
R287 VTAIL.n113 VTAIL.n95 171.744
R288 VTAIL.n114 VTAIL.n113 171.744
R289 VTAIL.n114 VTAIL.n91 171.744
R290 VTAIL.n122 VTAIL.n91 171.744
R291 VTAIL.n123 VTAIL.n122 171.744
R292 VTAIL.n124 VTAIL.n123 171.744
R293 VTAIL.n296 VTAIL.n295 171.744
R294 VTAIL.n295 VTAIL.n294 171.744
R295 VTAIL.n294 VTAIL.n263 171.744
R296 VTAIL.n287 VTAIL.n263 171.744
R297 VTAIL.n287 VTAIL.n286 171.744
R298 VTAIL.n286 VTAIL.n268 171.744
R299 VTAIL.n279 VTAIL.n268 171.744
R300 VTAIL.n279 VTAIL.n278 171.744
R301 VTAIL.n278 VTAIL.n272 171.744
R302 VTAIL.n252 VTAIL.n251 171.744
R303 VTAIL.n251 VTAIL.n250 171.744
R304 VTAIL.n250 VTAIL.n219 171.744
R305 VTAIL.n243 VTAIL.n219 171.744
R306 VTAIL.n243 VTAIL.n242 171.744
R307 VTAIL.n242 VTAIL.n224 171.744
R308 VTAIL.n235 VTAIL.n224 171.744
R309 VTAIL.n235 VTAIL.n234 171.744
R310 VTAIL.n234 VTAIL.n228 171.744
R311 VTAIL.n210 VTAIL.n209 171.744
R312 VTAIL.n209 VTAIL.n208 171.744
R313 VTAIL.n208 VTAIL.n177 171.744
R314 VTAIL.n201 VTAIL.n177 171.744
R315 VTAIL.n201 VTAIL.n200 171.744
R316 VTAIL.n200 VTAIL.n182 171.744
R317 VTAIL.n193 VTAIL.n182 171.744
R318 VTAIL.n193 VTAIL.n192 171.744
R319 VTAIL.n192 VTAIL.n186 171.744
R320 VTAIL.n166 VTAIL.n165 171.744
R321 VTAIL.n165 VTAIL.n164 171.744
R322 VTAIL.n164 VTAIL.n133 171.744
R323 VTAIL.n157 VTAIL.n133 171.744
R324 VTAIL.n157 VTAIL.n156 171.744
R325 VTAIL.n156 VTAIL.n138 171.744
R326 VTAIL.n149 VTAIL.n138 171.744
R327 VTAIL.n149 VTAIL.n148 171.744
R328 VTAIL.n148 VTAIL.n142 171.744
R329 VTAIL.t2 VTAIL.n313 85.8723
R330 VTAIL.t1 VTAIL.n13 85.8723
R331 VTAIL.t12 VTAIL.n55 85.8723
R332 VTAIL.t11 VTAIL.n99 85.8723
R333 VTAIL.t8 VTAIL.n272 85.8723
R334 VTAIL.t10 VTAIL.n228 85.8723
R335 VTAIL.t7 VTAIL.n186 85.8723
R336 VTAIL.t6 VTAIL.n142 85.8723
R337 VTAIL.n259 VTAIL.n258 69.9471
R338 VTAIL.n173 VTAIL.n172 69.9471
R339 VTAIL.n1 VTAIL.n0 69.9469
R340 VTAIL.n87 VTAIL.n86 69.9469
R341 VTAIL.n343 VTAIL.n342 36.452
R342 VTAIL.n43 VTAIL.n42 36.452
R343 VTAIL.n85 VTAIL.n84 36.452
R344 VTAIL.n129 VTAIL.n128 36.452
R345 VTAIL.n301 VTAIL.n300 36.452
R346 VTAIL.n257 VTAIL.n256 36.452
R347 VTAIL.n215 VTAIL.n214 36.452
R348 VTAIL.n171 VTAIL.n170 36.452
R349 VTAIL.n343 VTAIL.n301 23.0048
R350 VTAIL.n171 VTAIL.n129 23.0048
R351 VTAIL.n339 VTAIL.n304 13.1884
R352 VTAIL.n39 VTAIL.n4 13.1884
R353 VTAIL.n81 VTAIL.n46 13.1884
R354 VTAIL.n125 VTAIL.n90 13.1884
R355 VTAIL.n297 VTAIL.n262 13.1884
R356 VTAIL.n253 VTAIL.n218 13.1884
R357 VTAIL.n211 VTAIL.n176 13.1884
R358 VTAIL.n167 VTAIL.n132 13.1884
R359 VTAIL.n335 VTAIL.n334 12.8005
R360 VTAIL.n340 VTAIL.n302 12.8005
R361 VTAIL.n35 VTAIL.n34 12.8005
R362 VTAIL.n40 VTAIL.n2 12.8005
R363 VTAIL.n77 VTAIL.n76 12.8005
R364 VTAIL.n82 VTAIL.n44 12.8005
R365 VTAIL.n121 VTAIL.n120 12.8005
R366 VTAIL.n126 VTAIL.n88 12.8005
R367 VTAIL.n298 VTAIL.n260 12.8005
R368 VTAIL.n293 VTAIL.n264 12.8005
R369 VTAIL.n254 VTAIL.n216 12.8005
R370 VTAIL.n249 VTAIL.n220 12.8005
R371 VTAIL.n212 VTAIL.n174 12.8005
R372 VTAIL.n207 VTAIL.n178 12.8005
R373 VTAIL.n168 VTAIL.n130 12.8005
R374 VTAIL.n163 VTAIL.n134 12.8005
R375 VTAIL.n333 VTAIL.n306 12.0247
R376 VTAIL.n33 VTAIL.n6 12.0247
R377 VTAIL.n75 VTAIL.n48 12.0247
R378 VTAIL.n119 VTAIL.n92 12.0247
R379 VTAIL.n292 VTAIL.n265 12.0247
R380 VTAIL.n248 VTAIL.n221 12.0247
R381 VTAIL.n206 VTAIL.n179 12.0247
R382 VTAIL.n162 VTAIL.n135 12.0247
R383 VTAIL.n330 VTAIL.n329 11.249
R384 VTAIL.n30 VTAIL.n29 11.249
R385 VTAIL.n72 VTAIL.n71 11.249
R386 VTAIL.n116 VTAIL.n115 11.249
R387 VTAIL.n289 VTAIL.n288 11.249
R388 VTAIL.n245 VTAIL.n244 11.249
R389 VTAIL.n203 VTAIL.n202 11.249
R390 VTAIL.n159 VTAIL.n158 11.249
R391 VTAIL.n315 VTAIL.n314 10.7238
R392 VTAIL.n15 VTAIL.n14 10.7238
R393 VTAIL.n57 VTAIL.n56 10.7238
R394 VTAIL.n101 VTAIL.n100 10.7238
R395 VTAIL.n274 VTAIL.n273 10.7238
R396 VTAIL.n230 VTAIL.n229 10.7238
R397 VTAIL.n188 VTAIL.n187 10.7238
R398 VTAIL.n144 VTAIL.n143 10.7238
R399 VTAIL.n326 VTAIL.n308 10.4732
R400 VTAIL.n26 VTAIL.n8 10.4732
R401 VTAIL.n68 VTAIL.n50 10.4732
R402 VTAIL.n112 VTAIL.n94 10.4732
R403 VTAIL.n285 VTAIL.n267 10.4732
R404 VTAIL.n241 VTAIL.n223 10.4732
R405 VTAIL.n199 VTAIL.n181 10.4732
R406 VTAIL.n155 VTAIL.n137 10.4732
R407 VTAIL.n325 VTAIL.n310 9.69747
R408 VTAIL.n25 VTAIL.n10 9.69747
R409 VTAIL.n67 VTAIL.n52 9.69747
R410 VTAIL.n111 VTAIL.n96 9.69747
R411 VTAIL.n284 VTAIL.n269 9.69747
R412 VTAIL.n240 VTAIL.n225 9.69747
R413 VTAIL.n198 VTAIL.n183 9.69747
R414 VTAIL.n154 VTAIL.n139 9.69747
R415 VTAIL.n342 VTAIL.n341 9.45567
R416 VTAIL.n42 VTAIL.n41 9.45567
R417 VTAIL.n84 VTAIL.n83 9.45567
R418 VTAIL.n128 VTAIL.n127 9.45567
R419 VTAIL.n300 VTAIL.n299 9.45567
R420 VTAIL.n256 VTAIL.n255 9.45567
R421 VTAIL.n214 VTAIL.n213 9.45567
R422 VTAIL.n170 VTAIL.n169 9.45567
R423 VTAIL.n341 VTAIL.n340 9.3005
R424 VTAIL.n317 VTAIL.n316 9.3005
R425 VTAIL.n312 VTAIL.n311 9.3005
R426 VTAIL.n323 VTAIL.n322 9.3005
R427 VTAIL.n325 VTAIL.n324 9.3005
R428 VTAIL.n308 VTAIL.n307 9.3005
R429 VTAIL.n331 VTAIL.n330 9.3005
R430 VTAIL.n333 VTAIL.n332 9.3005
R431 VTAIL.n334 VTAIL.n303 9.3005
R432 VTAIL.n41 VTAIL.n40 9.3005
R433 VTAIL.n17 VTAIL.n16 9.3005
R434 VTAIL.n12 VTAIL.n11 9.3005
R435 VTAIL.n23 VTAIL.n22 9.3005
R436 VTAIL.n25 VTAIL.n24 9.3005
R437 VTAIL.n8 VTAIL.n7 9.3005
R438 VTAIL.n31 VTAIL.n30 9.3005
R439 VTAIL.n33 VTAIL.n32 9.3005
R440 VTAIL.n34 VTAIL.n3 9.3005
R441 VTAIL.n83 VTAIL.n82 9.3005
R442 VTAIL.n59 VTAIL.n58 9.3005
R443 VTAIL.n54 VTAIL.n53 9.3005
R444 VTAIL.n65 VTAIL.n64 9.3005
R445 VTAIL.n67 VTAIL.n66 9.3005
R446 VTAIL.n50 VTAIL.n49 9.3005
R447 VTAIL.n73 VTAIL.n72 9.3005
R448 VTAIL.n75 VTAIL.n74 9.3005
R449 VTAIL.n76 VTAIL.n45 9.3005
R450 VTAIL.n127 VTAIL.n126 9.3005
R451 VTAIL.n103 VTAIL.n102 9.3005
R452 VTAIL.n98 VTAIL.n97 9.3005
R453 VTAIL.n109 VTAIL.n108 9.3005
R454 VTAIL.n111 VTAIL.n110 9.3005
R455 VTAIL.n94 VTAIL.n93 9.3005
R456 VTAIL.n117 VTAIL.n116 9.3005
R457 VTAIL.n119 VTAIL.n118 9.3005
R458 VTAIL.n120 VTAIL.n89 9.3005
R459 VTAIL.n276 VTAIL.n275 9.3005
R460 VTAIL.n271 VTAIL.n270 9.3005
R461 VTAIL.n282 VTAIL.n281 9.3005
R462 VTAIL.n284 VTAIL.n283 9.3005
R463 VTAIL.n267 VTAIL.n266 9.3005
R464 VTAIL.n290 VTAIL.n289 9.3005
R465 VTAIL.n292 VTAIL.n291 9.3005
R466 VTAIL.n264 VTAIL.n261 9.3005
R467 VTAIL.n299 VTAIL.n298 9.3005
R468 VTAIL.n232 VTAIL.n231 9.3005
R469 VTAIL.n227 VTAIL.n226 9.3005
R470 VTAIL.n238 VTAIL.n237 9.3005
R471 VTAIL.n240 VTAIL.n239 9.3005
R472 VTAIL.n223 VTAIL.n222 9.3005
R473 VTAIL.n246 VTAIL.n245 9.3005
R474 VTAIL.n248 VTAIL.n247 9.3005
R475 VTAIL.n220 VTAIL.n217 9.3005
R476 VTAIL.n255 VTAIL.n254 9.3005
R477 VTAIL.n190 VTAIL.n189 9.3005
R478 VTAIL.n185 VTAIL.n184 9.3005
R479 VTAIL.n196 VTAIL.n195 9.3005
R480 VTAIL.n198 VTAIL.n197 9.3005
R481 VTAIL.n181 VTAIL.n180 9.3005
R482 VTAIL.n204 VTAIL.n203 9.3005
R483 VTAIL.n206 VTAIL.n205 9.3005
R484 VTAIL.n178 VTAIL.n175 9.3005
R485 VTAIL.n213 VTAIL.n212 9.3005
R486 VTAIL.n146 VTAIL.n145 9.3005
R487 VTAIL.n141 VTAIL.n140 9.3005
R488 VTAIL.n152 VTAIL.n151 9.3005
R489 VTAIL.n154 VTAIL.n153 9.3005
R490 VTAIL.n137 VTAIL.n136 9.3005
R491 VTAIL.n160 VTAIL.n159 9.3005
R492 VTAIL.n162 VTAIL.n161 9.3005
R493 VTAIL.n134 VTAIL.n131 9.3005
R494 VTAIL.n169 VTAIL.n168 9.3005
R495 VTAIL.n322 VTAIL.n321 8.92171
R496 VTAIL.n22 VTAIL.n21 8.92171
R497 VTAIL.n64 VTAIL.n63 8.92171
R498 VTAIL.n108 VTAIL.n107 8.92171
R499 VTAIL.n281 VTAIL.n280 8.92171
R500 VTAIL.n237 VTAIL.n236 8.92171
R501 VTAIL.n195 VTAIL.n194 8.92171
R502 VTAIL.n151 VTAIL.n150 8.92171
R503 VTAIL.n318 VTAIL.n312 8.14595
R504 VTAIL.n18 VTAIL.n12 8.14595
R505 VTAIL.n60 VTAIL.n54 8.14595
R506 VTAIL.n104 VTAIL.n98 8.14595
R507 VTAIL.n277 VTAIL.n271 8.14595
R508 VTAIL.n233 VTAIL.n227 8.14595
R509 VTAIL.n191 VTAIL.n185 8.14595
R510 VTAIL.n147 VTAIL.n141 8.14595
R511 VTAIL.n317 VTAIL.n314 7.3702
R512 VTAIL.n17 VTAIL.n14 7.3702
R513 VTAIL.n59 VTAIL.n56 7.3702
R514 VTAIL.n103 VTAIL.n100 7.3702
R515 VTAIL.n276 VTAIL.n273 7.3702
R516 VTAIL.n232 VTAIL.n229 7.3702
R517 VTAIL.n190 VTAIL.n187 7.3702
R518 VTAIL.n146 VTAIL.n143 7.3702
R519 VTAIL.n318 VTAIL.n317 5.81868
R520 VTAIL.n18 VTAIL.n17 5.81868
R521 VTAIL.n60 VTAIL.n59 5.81868
R522 VTAIL.n104 VTAIL.n103 5.81868
R523 VTAIL.n277 VTAIL.n276 5.81868
R524 VTAIL.n233 VTAIL.n232 5.81868
R525 VTAIL.n191 VTAIL.n190 5.81868
R526 VTAIL.n147 VTAIL.n146 5.81868
R527 VTAIL.n321 VTAIL.n312 5.04292
R528 VTAIL.n21 VTAIL.n12 5.04292
R529 VTAIL.n63 VTAIL.n54 5.04292
R530 VTAIL.n107 VTAIL.n98 5.04292
R531 VTAIL.n280 VTAIL.n271 5.04292
R532 VTAIL.n236 VTAIL.n227 5.04292
R533 VTAIL.n194 VTAIL.n185 5.04292
R534 VTAIL.n150 VTAIL.n141 5.04292
R535 VTAIL.n322 VTAIL.n310 4.26717
R536 VTAIL.n22 VTAIL.n10 4.26717
R537 VTAIL.n64 VTAIL.n52 4.26717
R538 VTAIL.n108 VTAIL.n96 4.26717
R539 VTAIL.n281 VTAIL.n269 4.26717
R540 VTAIL.n237 VTAIL.n225 4.26717
R541 VTAIL.n195 VTAIL.n183 4.26717
R542 VTAIL.n151 VTAIL.n139 4.26717
R543 VTAIL.n0 VTAIL.t3 4.05349
R544 VTAIL.n0 VTAIL.t0 4.05349
R545 VTAIL.n86 VTAIL.t9 4.05349
R546 VTAIL.n86 VTAIL.t14 4.05349
R547 VTAIL.n258 VTAIL.t13 4.05349
R548 VTAIL.n258 VTAIL.t15 4.05349
R549 VTAIL.n172 VTAIL.t5 4.05349
R550 VTAIL.n172 VTAIL.t4 4.05349
R551 VTAIL.n173 VTAIL.n171 3.72464
R552 VTAIL.n215 VTAIL.n173 3.72464
R553 VTAIL.n259 VTAIL.n257 3.72464
R554 VTAIL.n301 VTAIL.n259 3.72464
R555 VTAIL.n129 VTAIL.n87 3.72464
R556 VTAIL.n87 VTAIL.n85 3.72464
R557 VTAIL.n43 VTAIL.n1 3.72464
R558 VTAIL VTAIL.n343 3.66645
R559 VTAIL.n326 VTAIL.n325 3.49141
R560 VTAIL.n26 VTAIL.n25 3.49141
R561 VTAIL.n68 VTAIL.n67 3.49141
R562 VTAIL.n112 VTAIL.n111 3.49141
R563 VTAIL.n285 VTAIL.n284 3.49141
R564 VTAIL.n241 VTAIL.n240 3.49141
R565 VTAIL.n199 VTAIL.n198 3.49141
R566 VTAIL.n155 VTAIL.n154 3.49141
R567 VTAIL.n329 VTAIL.n308 2.71565
R568 VTAIL.n29 VTAIL.n8 2.71565
R569 VTAIL.n71 VTAIL.n50 2.71565
R570 VTAIL.n115 VTAIL.n94 2.71565
R571 VTAIL.n288 VTAIL.n267 2.71565
R572 VTAIL.n244 VTAIL.n223 2.71565
R573 VTAIL.n202 VTAIL.n181 2.71565
R574 VTAIL.n158 VTAIL.n137 2.71565
R575 VTAIL.n316 VTAIL.n315 2.4129
R576 VTAIL.n16 VTAIL.n15 2.4129
R577 VTAIL.n58 VTAIL.n57 2.4129
R578 VTAIL.n102 VTAIL.n101 2.4129
R579 VTAIL.n275 VTAIL.n274 2.4129
R580 VTAIL.n231 VTAIL.n230 2.4129
R581 VTAIL.n189 VTAIL.n188 2.4129
R582 VTAIL.n145 VTAIL.n144 2.4129
R583 VTAIL.n330 VTAIL.n306 1.93989
R584 VTAIL.n30 VTAIL.n6 1.93989
R585 VTAIL.n72 VTAIL.n48 1.93989
R586 VTAIL.n116 VTAIL.n92 1.93989
R587 VTAIL.n289 VTAIL.n265 1.93989
R588 VTAIL.n245 VTAIL.n221 1.93989
R589 VTAIL.n203 VTAIL.n179 1.93989
R590 VTAIL.n159 VTAIL.n135 1.93989
R591 VTAIL.n335 VTAIL.n333 1.16414
R592 VTAIL.n342 VTAIL.n302 1.16414
R593 VTAIL.n35 VTAIL.n33 1.16414
R594 VTAIL.n42 VTAIL.n2 1.16414
R595 VTAIL.n77 VTAIL.n75 1.16414
R596 VTAIL.n84 VTAIL.n44 1.16414
R597 VTAIL.n121 VTAIL.n119 1.16414
R598 VTAIL.n128 VTAIL.n88 1.16414
R599 VTAIL.n300 VTAIL.n260 1.16414
R600 VTAIL.n293 VTAIL.n292 1.16414
R601 VTAIL.n256 VTAIL.n216 1.16414
R602 VTAIL.n249 VTAIL.n248 1.16414
R603 VTAIL.n214 VTAIL.n174 1.16414
R604 VTAIL.n207 VTAIL.n206 1.16414
R605 VTAIL.n170 VTAIL.n130 1.16414
R606 VTAIL.n163 VTAIL.n162 1.16414
R607 VTAIL.n257 VTAIL.n215 0.470328
R608 VTAIL.n85 VTAIL.n43 0.470328
R609 VTAIL.n334 VTAIL.n304 0.388379
R610 VTAIL.n340 VTAIL.n339 0.388379
R611 VTAIL.n34 VTAIL.n4 0.388379
R612 VTAIL.n40 VTAIL.n39 0.388379
R613 VTAIL.n76 VTAIL.n46 0.388379
R614 VTAIL.n82 VTAIL.n81 0.388379
R615 VTAIL.n120 VTAIL.n90 0.388379
R616 VTAIL.n126 VTAIL.n125 0.388379
R617 VTAIL.n298 VTAIL.n297 0.388379
R618 VTAIL.n264 VTAIL.n262 0.388379
R619 VTAIL.n254 VTAIL.n253 0.388379
R620 VTAIL.n220 VTAIL.n218 0.388379
R621 VTAIL.n212 VTAIL.n211 0.388379
R622 VTAIL.n178 VTAIL.n176 0.388379
R623 VTAIL.n168 VTAIL.n167 0.388379
R624 VTAIL.n134 VTAIL.n132 0.388379
R625 VTAIL.n316 VTAIL.n311 0.155672
R626 VTAIL.n323 VTAIL.n311 0.155672
R627 VTAIL.n324 VTAIL.n323 0.155672
R628 VTAIL.n324 VTAIL.n307 0.155672
R629 VTAIL.n331 VTAIL.n307 0.155672
R630 VTAIL.n332 VTAIL.n331 0.155672
R631 VTAIL.n332 VTAIL.n303 0.155672
R632 VTAIL.n341 VTAIL.n303 0.155672
R633 VTAIL.n16 VTAIL.n11 0.155672
R634 VTAIL.n23 VTAIL.n11 0.155672
R635 VTAIL.n24 VTAIL.n23 0.155672
R636 VTAIL.n24 VTAIL.n7 0.155672
R637 VTAIL.n31 VTAIL.n7 0.155672
R638 VTAIL.n32 VTAIL.n31 0.155672
R639 VTAIL.n32 VTAIL.n3 0.155672
R640 VTAIL.n41 VTAIL.n3 0.155672
R641 VTAIL.n58 VTAIL.n53 0.155672
R642 VTAIL.n65 VTAIL.n53 0.155672
R643 VTAIL.n66 VTAIL.n65 0.155672
R644 VTAIL.n66 VTAIL.n49 0.155672
R645 VTAIL.n73 VTAIL.n49 0.155672
R646 VTAIL.n74 VTAIL.n73 0.155672
R647 VTAIL.n74 VTAIL.n45 0.155672
R648 VTAIL.n83 VTAIL.n45 0.155672
R649 VTAIL.n102 VTAIL.n97 0.155672
R650 VTAIL.n109 VTAIL.n97 0.155672
R651 VTAIL.n110 VTAIL.n109 0.155672
R652 VTAIL.n110 VTAIL.n93 0.155672
R653 VTAIL.n117 VTAIL.n93 0.155672
R654 VTAIL.n118 VTAIL.n117 0.155672
R655 VTAIL.n118 VTAIL.n89 0.155672
R656 VTAIL.n127 VTAIL.n89 0.155672
R657 VTAIL.n299 VTAIL.n261 0.155672
R658 VTAIL.n291 VTAIL.n261 0.155672
R659 VTAIL.n291 VTAIL.n290 0.155672
R660 VTAIL.n290 VTAIL.n266 0.155672
R661 VTAIL.n283 VTAIL.n266 0.155672
R662 VTAIL.n283 VTAIL.n282 0.155672
R663 VTAIL.n282 VTAIL.n270 0.155672
R664 VTAIL.n275 VTAIL.n270 0.155672
R665 VTAIL.n255 VTAIL.n217 0.155672
R666 VTAIL.n247 VTAIL.n217 0.155672
R667 VTAIL.n247 VTAIL.n246 0.155672
R668 VTAIL.n246 VTAIL.n222 0.155672
R669 VTAIL.n239 VTAIL.n222 0.155672
R670 VTAIL.n239 VTAIL.n238 0.155672
R671 VTAIL.n238 VTAIL.n226 0.155672
R672 VTAIL.n231 VTAIL.n226 0.155672
R673 VTAIL.n213 VTAIL.n175 0.155672
R674 VTAIL.n205 VTAIL.n175 0.155672
R675 VTAIL.n205 VTAIL.n204 0.155672
R676 VTAIL.n204 VTAIL.n180 0.155672
R677 VTAIL.n197 VTAIL.n180 0.155672
R678 VTAIL.n197 VTAIL.n196 0.155672
R679 VTAIL.n196 VTAIL.n184 0.155672
R680 VTAIL.n189 VTAIL.n184 0.155672
R681 VTAIL.n169 VTAIL.n131 0.155672
R682 VTAIL.n161 VTAIL.n131 0.155672
R683 VTAIL.n161 VTAIL.n160 0.155672
R684 VTAIL.n160 VTAIL.n136 0.155672
R685 VTAIL.n153 VTAIL.n136 0.155672
R686 VTAIL.n153 VTAIL.n152 0.155672
R687 VTAIL.n152 VTAIL.n140 0.155672
R688 VTAIL.n145 VTAIL.n140 0.155672
R689 VTAIL VTAIL.n1 0.0586897
R690 VN.n75 VN.n39 161.3
R691 VN.n74 VN.n73 161.3
R692 VN.n72 VN.n40 161.3
R693 VN.n71 VN.n70 161.3
R694 VN.n69 VN.n41 161.3
R695 VN.n68 VN.n67 161.3
R696 VN.n66 VN.n42 161.3
R697 VN.n65 VN.n64 161.3
R698 VN.n62 VN.n43 161.3
R699 VN.n61 VN.n60 161.3
R700 VN.n59 VN.n44 161.3
R701 VN.n58 VN.n57 161.3
R702 VN.n56 VN.n45 161.3
R703 VN.n55 VN.n54 161.3
R704 VN.n53 VN.n46 161.3
R705 VN.n52 VN.n51 161.3
R706 VN.n50 VN.n47 161.3
R707 VN.n36 VN.n0 161.3
R708 VN.n35 VN.n34 161.3
R709 VN.n33 VN.n1 161.3
R710 VN.n32 VN.n31 161.3
R711 VN.n30 VN.n2 161.3
R712 VN.n29 VN.n28 161.3
R713 VN.n27 VN.n3 161.3
R714 VN.n26 VN.n25 161.3
R715 VN.n23 VN.n4 161.3
R716 VN.n22 VN.n21 161.3
R717 VN.n20 VN.n5 161.3
R718 VN.n19 VN.n18 161.3
R719 VN.n17 VN.n6 161.3
R720 VN.n16 VN.n15 161.3
R721 VN.n14 VN.n7 161.3
R722 VN.n13 VN.n12 161.3
R723 VN.n11 VN.n8 161.3
R724 VN.n9 VN.t7 80.5654
R725 VN.n48 VN.t3 80.5654
R726 VN.n10 VN.n9 67.5408
R727 VN.n49 VN.n48 67.5408
R728 VN.n38 VN.n37 58.7717
R729 VN.n77 VN.n76 58.7717
R730 VN.n31 VN.n30 56.5617
R731 VN.n70 VN.n69 56.5617
R732 VN VN.n77 54.7165
R733 VN.n10 VN.t5 48.4421
R734 VN.n24 VN.t1 48.4421
R735 VN.n37 VN.t6 48.4421
R736 VN.n49 VN.t4 48.4421
R737 VN.n63 VN.t2 48.4421
R738 VN.n76 VN.t0 48.4421
R739 VN.n17 VN.n16 40.577
R740 VN.n18 VN.n17 40.577
R741 VN.n56 VN.n55 40.577
R742 VN.n57 VN.n56 40.577
R743 VN.n12 VN.n11 24.5923
R744 VN.n12 VN.n7 24.5923
R745 VN.n16 VN.n7 24.5923
R746 VN.n18 VN.n5 24.5923
R747 VN.n22 VN.n5 24.5923
R748 VN.n23 VN.n22 24.5923
R749 VN.n25 VN.n3 24.5923
R750 VN.n29 VN.n3 24.5923
R751 VN.n30 VN.n29 24.5923
R752 VN.n31 VN.n1 24.5923
R753 VN.n35 VN.n1 24.5923
R754 VN.n36 VN.n35 24.5923
R755 VN.n55 VN.n46 24.5923
R756 VN.n51 VN.n46 24.5923
R757 VN.n51 VN.n50 24.5923
R758 VN.n69 VN.n68 24.5923
R759 VN.n68 VN.n42 24.5923
R760 VN.n64 VN.n42 24.5923
R761 VN.n62 VN.n61 24.5923
R762 VN.n61 VN.n44 24.5923
R763 VN.n57 VN.n44 24.5923
R764 VN.n75 VN.n74 24.5923
R765 VN.n74 VN.n40 24.5923
R766 VN.n70 VN.n40 24.5923
R767 VN.n37 VN.n36 23.6087
R768 VN.n76 VN.n75 23.6087
R769 VN.n25 VN.n24 16.7229
R770 VN.n64 VN.n63 16.7229
R771 VN.n11 VN.n10 7.86989
R772 VN.n24 VN.n23 7.86989
R773 VN.n50 VN.n49 7.86989
R774 VN.n63 VN.n62 7.86989
R775 VN.n48 VN.n47 2.56253
R776 VN.n9 VN.n8 2.56253
R777 VN.n77 VN.n39 0.417304
R778 VN.n38 VN.n0 0.417304
R779 VN VN.n38 0.394524
R780 VN.n73 VN.n39 0.189894
R781 VN.n73 VN.n72 0.189894
R782 VN.n72 VN.n71 0.189894
R783 VN.n71 VN.n41 0.189894
R784 VN.n67 VN.n41 0.189894
R785 VN.n67 VN.n66 0.189894
R786 VN.n66 VN.n65 0.189894
R787 VN.n65 VN.n43 0.189894
R788 VN.n60 VN.n43 0.189894
R789 VN.n60 VN.n59 0.189894
R790 VN.n59 VN.n58 0.189894
R791 VN.n58 VN.n45 0.189894
R792 VN.n54 VN.n45 0.189894
R793 VN.n54 VN.n53 0.189894
R794 VN.n53 VN.n52 0.189894
R795 VN.n52 VN.n47 0.189894
R796 VN.n13 VN.n8 0.189894
R797 VN.n14 VN.n13 0.189894
R798 VN.n15 VN.n14 0.189894
R799 VN.n15 VN.n6 0.189894
R800 VN.n19 VN.n6 0.189894
R801 VN.n20 VN.n19 0.189894
R802 VN.n21 VN.n20 0.189894
R803 VN.n21 VN.n4 0.189894
R804 VN.n26 VN.n4 0.189894
R805 VN.n27 VN.n26 0.189894
R806 VN.n28 VN.n27 0.189894
R807 VN.n28 VN.n2 0.189894
R808 VN.n32 VN.n2 0.189894
R809 VN.n33 VN.n32 0.189894
R810 VN.n34 VN.n33 0.189894
R811 VN.n34 VN.n0 0.189894
R812 VDD2.n2 VDD2.n1 88.4325
R813 VDD2.n2 VDD2.n0 88.4325
R814 VDD2 VDD2.n5 88.4296
R815 VDD2.n4 VDD2.n3 86.6259
R816 VDD2.n4 VDD2.n2 47.3877
R817 VDD2.n5 VDD2.t3 4.05349
R818 VDD2.n5 VDD2.t4 4.05349
R819 VDD2.n3 VDD2.t7 4.05349
R820 VDD2.n3 VDD2.t5 4.05349
R821 VDD2.n1 VDD2.t6 4.05349
R822 VDD2.n1 VDD2.t1 4.05349
R823 VDD2.n0 VDD2.t0 4.05349
R824 VDD2.n0 VDD2.t2 4.05349
R825 VDD2 VDD2.n4 1.92076
R826 B.n432 B.n149 585
R827 B.n431 B.n430 585
R828 B.n429 B.n150 585
R829 B.n428 B.n427 585
R830 B.n426 B.n151 585
R831 B.n425 B.n424 585
R832 B.n423 B.n152 585
R833 B.n422 B.n421 585
R834 B.n420 B.n153 585
R835 B.n419 B.n418 585
R836 B.n417 B.n154 585
R837 B.n416 B.n415 585
R838 B.n414 B.n155 585
R839 B.n413 B.n412 585
R840 B.n411 B.n156 585
R841 B.n410 B.n409 585
R842 B.n408 B.n157 585
R843 B.n407 B.n406 585
R844 B.n405 B.n158 585
R845 B.n404 B.n403 585
R846 B.n402 B.n159 585
R847 B.n401 B.n400 585
R848 B.n399 B.n160 585
R849 B.n398 B.n397 585
R850 B.n396 B.n161 585
R851 B.n395 B.n394 585
R852 B.n393 B.n162 585
R853 B.n392 B.n391 585
R854 B.n390 B.n163 585
R855 B.n389 B.n388 585
R856 B.n386 B.n164 585
R857 B.n385 B.n384 585
R858 B.n383 B.n167 585
R859 B.n382 B.n381 585
R860 B.n380 B.n168 585
R861 B.n379 B.n378 585
R862 B.n377 B.n169 585
R863 B.n376 B.n375 585
R864 B.n374 B.n170 585
R865 B.n372 B.n371 585
R866 B.n370 B.n173 585
R867 B.n369 B.n368 585
R868 B.n367 B.n174 585
R869 B.n366 B.n365 585
R870 B.n364 B.n175 585
R871 B.n363 B.n362 585
R872 B.n361 B.n176 585
R873 B.n360 B.n359 585
R874 B.n358 B.n177 585
R875 B.n357 B.n356 585
R876 B.n355 B.n178 585
R877 B.n354 B.n353 585
R878 B.n352 B.n179 585
R879 B.n351 B.n350 585
R880 B.n349 B.n180 585
R881 B.n348 B.n347 585
R882 B.n346 B.n181 585
R883 B.n345 B.n344 585
R884 B.n343 B.n182 585
R885 B.n342 B.n341 585
R886 B.n340 B.n183 585
R887 B.n339 B.n338 585
R888 B.n337 B.n184 585
R889 B.n336 B.n335 585
R890 B.n334 B.n185 585
R891 B.n333 B.n332 585
R892 B.n331 B.n186 585
R893 B.n330 B.n329 585
R894 B.n328 B.n187 585
R895 B.n434 B.n433 585
R896 B.n435 B.n148 585
R897 B.n437 B.n436 585
R898 B.n438 B.n147 585
R899 B.n440 B.n439 585
R900 B.n441 B.n146 585
R901 B.n443 B.n442 585
R902 B.n444 B.n145 585
R903 B.n446 B.n445 585
R904 B.n447 B.n144 585
R905 B.n449 B.n448 585
R906 B.n450 B.n143 585
R907 B.n452 B.n451 585
R908 B.n453 B.n142 585
R909 B.n455 B.n454 585
R910 B.n456 B.n141 585
R911 B.n458 B.n457 585
R912 B.n459 B.n140 585
R913 B.n461 B.n460 585
R914 B.n462 B.n139 585
R915 B.n464 B.n463 585
R916 B.n465 B.n138 585
R917 B.n467 B.n466 585
R918 B.n468 B.n137 585
R919 B.n470 B.n469 585
R920 B.n471 B.n136 585
R921 B.n473 B.n472 585
R922 B.n474 B.n135 585
R923 B.n476 B.n475 585
R924 B.n477 B.n134 585
R925 B.n479 B.n478 585
R926 B.n480 B.n133 585
R927 B.n482 B.n481 585
R928 B.n483 B.n132 585
R929 B.n485 B.n484 585
R930 B.n486 B.n131 585
R931 B.n488 B.n487 585
R932 B.n489 B.n130 585
R933 B.n491 B.n490 585
R934 B.n492 B.n129 585
R935 B.n494 B.n493 585
R936 B.n495 B.n128 585
R937 B.n497 B.n496 585
R938 B.n498 B.n127 585
R939 B.n500 B.n499 585
R940 B.n501 B.n126 585
R941 B.n503 B.n502 585
R942 B.n504 B.n125 585
R943 B.n506 B.n505 585
R944 B.n507 B.n124 585
R945 B.n509 B.n508 585
R946 B.n510 B.n123 585
R947 B.n512 B.n511 585
R948 B.n513 B.n122 585
R949 B.n515 B.n514 585
R950 B.n516 B.n121 585
R951 B.n518 B.n517 585
R952 B.n519 B.n120 585
R953 B.n521 B.n520 585
R954 B.n522 B.n119 585
R955 B.n524 B.n523 585
R956 B.n525 B.n118 585
R957 B.n527 B.n526 585
R958 B.n528 B.n117 585
R959 B.n530 B.n529 585
R960 B.n531 B.n116 585
R961 B.n533 B.n532 585
R962 B.n534 B.n115 585
R963 B.n536 B.n535 585
R964 B.n537 B.n114 585
R965 B.n539 B.n538 585
R966 B.n540 B.n113 585
R967 B.n542 B.n541 585
R968 B.n543 B.n112 585
R969 B.n545 B.n544 585
R970 B.n546 B.n111 585
R971 B.n548 B.n547 585
R972 B.n549 B.n110 585
R973 B.n551 B.n550 585
R974 B.n552 B.n109 585
R975 B.n554 B.n553 585
R976 B.n555 B.n108 585
R977 B.n557 B.n556 585
R978 B.n558 B.n107 585
R979 B.n560 B.n559 585
R980 B.n561 B.n106 585
R981 B.n563 B.n562 585
R982 B.n564 B.n105 585
R983 B.n566 B.n565 585
R984 B.n567 B.n104 585
R985 B.n569 B.n568 585
R986 B.n570 B.n103 585
R987 B.n572 B.n571 585
R988 B.n573 B.n102 585
R989 B.n575 B.n574 585
R990 B.n576 B.n101 585
R991 B.n578 B.n577 585
R992 B.n579 B.n100 585
R993 B.n581 B.n580 585
R994 B.n582 B.n99 585
R995 B.n584 B.n583 585
R996 B.n585 B.n98 585
R997 B.n587 B.n586 585
R998 B.n588 B.n97 585
R999 B.n590 B.n589 585
R1000 B.n591 B.n96 585
R1001 B.n593 B.n592 585
R1002 B.n594 B.n95 585
R1003 B.n596 B.n595 585
R1004 B.n597 B.n94 585
R1005 B.n599 B.n598 585
R1006 B.n600 B.n93 585
R1007 B.n602 B.n601 585
R1008 B.n603 B.n92 585
R1009 B.n605 B.n604 585
R1010 B.n606 B.n91 585
R1011 B.n608 B.n607 585
R1012 B.n609 B.n90 585
R1013 B.n611 B.n610 585
R1014 B.n612 B.n89 585
R1015 B.n614 B.n613 585
R1016 B.n615 B.n88 585
R1017 B.n617 B.n616 585
R1018 B.n618 B.n87 585
R1019 B.n620 B.n619 585
R1020 B.n621 B.n86 585
R1021 B.n623 B.n622 585
R1022 B.n624 B.n85 585
R1023 B.n626 B.n625 585
R1024 B.n627 B.n84 585
R1025 B.n629 B.n628 585
R1026 B.n630 B.n83 585
R1027 B.n632 B.n631 585
R1028 B.n633 B.n82 585
R1029 B.n635 B.n634 585
R1030 B.n636 B.n81 585
R1031 B.n638 B.n637 585
R1032 B.n639 B.n80 585
R1033 B.n641 B.n640 585
R1034 B.n642 B.n79 585
R1035 B.n644 B.n643 585
R1036 B.n645 B.n78 585
R1037 B.n647 B.n646 585
R1038 B.n648 B.n77 585
R1039 B.n753 B.n752 585
R1040 B.n751 B.n38 585
R1041 B.n750 B.n749 585
R1042 B.n748 B.n39 585
R1043 B.n747 B.n746 585
R1044 B.n745 B.n40 585
R1045 B.n744 B.n743 585
R1046 B.n742 B.n41 585
R1047 B.n741 B.n740 585
R1048 B.n739 B.n42 585
R1049 B.n738 B.n737 585
R1050 B.n736 B.n43 585
R1051 B.n735 B.n734 585
R1052 B.n733 B.n44 585
R1053 B.n732 B.n731 585
R1054 B.n730 B.n45 585
R1055 B.n729 B.n728 585
R1056 B.n727 B.n46 585
R1057 B.n726 B.n725 585
R1058 B.n724 B.n47 585
R1059 B.n723 B.n722 585
R1060 B.n721 B.n48 585
R1061 B.n720 B.n719 585
R1062 B.n718 B.n49 585
R1063 B.n717 B.n716 585
R1064 B.n715 B.n50 585
R1065 B.n714 B.n713 585
R1066 B.n712 B.n51 585
R1067 B.n711 B.n710 585
R1068 B.n709 B.n52 585
R1069 B.n708 B.n707 585
R1070 B.n706 B.n53 585
R1071 B.n705 B.n704 585
R1072 B.n703 B.n57 585
R1073 B.n702 B.n701 585
R1074 B.n700 B.n58 585
R1075 B.n699 B.n698 585
R1076 B.n697 B.n59 585
R1077 B.n696 B.n695 585
R1078 B.n693 B.n60 585
R1079 B.n692 B.n691 585
R1080 B.n690 B.n63 585
R1081 B.n689 B.n688 585
R1082 B.n687 B.n64 585
R1083 B.n686 B.n685 585
R1084 B.n684 B.n65 585
R1085 B.n683 B.n682 585
R1086 B.n681 B.n66 585
R1087 B.n680 B.n679 585
R1088 B.n678 B.n67 585
R1089 B.n677 B.n676 585
R1090 B.n675 B.n68 585
R1091 B.n674 B.n673 585
R1092 B.n672 B.n69 585
R1093 B.n671 B.n670 585
R1094 B.n669 B.n70 585
R1095 B.n668 B.n667 585
R1096 B.n666 B.n71 585
R1097 B.n665 B.n664 585
R1098 B.n663 B.n72 585
R1099 B.n662 B.n661 585
R1100 B.n660 B.n73 585
R1101 B.n659 B.n658 585
R1102 B.n657 B.n74 585
R1103 B.n656 B.n655 585
R1104 B.n654 B.n75 585
R1105 B.n653 B.n652 585
R1106 B.n651 B.n76 585
R1107 B.n650 B.n649 585
R1108 B.n754 B.n37 585
R1109 B.n756 B.n755 585
R1110 B.n757 B.n36 585
R1111 B.n759 B.n758 585
R1112 B.n760 B.n35 585
R1113 B.n762 B.n761 585
R1114 B.n763 B.n34 585
R1115 B.n765 B.n764 585
R1116 B.n766 B.n33 585
R1117 B.n768 B.n767 585
R1118 B.n769 B.n32 585
R1119 B.n771 B.n770 585
R1120 B.n772 B.n31 585
R1121 B.n774 B.n773 585
R1122 B.n775 B.n30 585
R1123 B.n777 B.n776 585
R1124 B.n778 B.n29 585
R1125 B.n780 B.n779 585
R1126 B.n781 B.n28 585
R1127 B.n783 B.n782 585
R1128 B.n784 B.n27 585
R1129 B.n786 B.n785 585
R1130 B.n787 B.n26 585
R1131 B.n789 B.n788 585
R1132 B.n790 B.n25 585
R1133 B.n792 B.n791 585
R1134 B.n793 B.n24 585
R1135 B.n795 B.n794 585
R1136 B.n796 B.n23 585
R1137 B.n798 B.n797 585
R1138 B.n799 B.n22 585
R1139 B.n801 B.n800 585
R1140 B.n802 B.n21 585
R1141 B.n804 B.n803 585
R1142 B.n805 B.n20 585
R1143 B.n807 B.n806 585
R1144 B.n808 B.n19 585
R1145 B.n810 B.n809 585
R1146 B.n811 B.n18 585
R1147 B.n813 B.n812 585
R1148 B.n814 B.n17 585
R1149 B.n816 B.n815 585
R1150 B.n817 B.n16 585
R1151 B.n819 B.n818 585
R1152 B.n820 B.n15 585
R1153 B.n822 B.n821 585
R1154 B.n823 B.n14 585
R1155 B.n825 B.n824 585
R1156 B.n826 B.n13 585
R1157 B.n828 B.n827 585
R1158 B.n829 B.n12 585
R1159 B.n831 B.n830 585
R1160 B.n832 B.n11 585
R1161 B.n834 B.n833 585
R1162 B.n835 B.n10 585
R1163 B.n837 B.n836 585
R1164 B.n838 B.n9 585
R1165 B.n840 B.n839 585
R1166 B.n841 B.n8 585
R1167 B.n843 B.n842 585
R1168 B.n844 B.n7 585
R1169 B.n846 B.n845 585
R1170 B.n847 B.n6 585
R1171 B.n849 B.n848 585
R1172 B.n850 B.n5 585
R1173 B.n852 B.n851 585
R1174 B.n853 B.n4 585
R1175 B.n855 B.n854 585
R1176 B.n856 B.n3 585
R1177 B.n858 B.n857 585
R1178 B.n859 B.n0 585
R1179 B.n2 B.n1 585
R1180 B.n223 B.n222 585
R1181 B.n225 B.n224 585
R1182 B.n226 B.n221 585
R1183 B.n228 B.n227 585
R1184 B.n229 B.n220 585
R1185 B.n231 B.n230 585
R1186 B.n232 B.n219 585
R1187 B.n234 B.n233 585
R1188 B.n235 B.n218 585
R1189 B.n237 B.n236 585
R1190 B.n238 B.n217 585
R1191 B.n240 B.n239 585
R1192 B.n241 B.n216 585
R1193 B.n243 B.n242 585
R1194 B.n244 B.n215 585
R1195 B.n246 B.n245 585
R1196 B.n247 B.n214 585
R1197 B.n249 B.n248 585
R1198 B.n250 B.n213 585
R1199 B.n252 B.n251 585
R1200 B.n253 B.n212 585
R1201 B.n255 B.n254 585
R1202 B.n256 B.n211 585
R1203 B.n258 B.n257 585
R1204 B.n259 B.n210 585
R1205 B.n261 B.n260 585
R1206 B.n262 B.n209 585
R1207 B.n264 B.n263 585
R1208 B.n265 B.n208 585
R1209 B.n267 B.n266 585
R1210 B.n268 B.n207 585
R1211 B.n270 B.n269 585
R1212 B.n271 B.n206 585
R1213 B.n273 B.n272 585
R1214 B.n274 B.n205 585
R1215 B.n276 B.n275 585
R1216 B.n277 B.n204 585
R1217 B.n279 B.n278 585
R1218 B.n280 B.n203 585
R1219 B.n282 B.n281 585
R1220 B.n283 B.n202 585
R1221 B.n285 B.n284 585
R1222 B.n286 B.n201 585
R1223 B.n288 B.n287 585
R1224 B.n289 B.n200 585
R1225 B.n291 B.n290 585
R1226 B.n292 B.n199 585
R1227 B.n294 B.n293 585
R1228 B.n295 B.n198 585
R1229 B.n297 B.n296 585
R1230 B.n298 B.n197 585
R1231 B.n300 B.n299 585
R1232 B.n301 B.n196 585
R1233 B.n303 B.n302 585
R1234 B.n304 B.n195 585
R1235 B.n306 B.n305 585
R1236 B.n307 B.n194 585
R1237 B.n309 B.n308 585
R1238 B.n310 B.n193 585
R1239 B.n312 B.n311 585
R1240 B.n313 B.n192 585
R1241 B.n315 B.n314 585
R1242 B.n316 B.n191 585
R1243 B.n318 B.n317 585
R1244 B.n319 B.n190 585
R1245 B.n321 B.n320 585
R1246 B.n322 B.n189 585
R1247 B.n324 B.n323 585
R1248 B.n325 B.n188 585
R1249 B.n327 B.n326 585
R1250 B.n328 B.n327 554.963
R1251 B.n433 B.n432 554.963
R1252 B.n649 B.n648 554.963
R1253 B.n752 B.n37 554.963
R1254 B.n165 B.t1 387.86
R1255 B.n61 B.t8 387.86
R1256 B.n171 B.t10 387.86
R1257 B.n54 B.t5 387.86
R1258 B.n166 B.t2 304.079
R1259 B.n62 B.t7 304.079
R1260 B.n172 B.t11 304.077
R1261 B.n55 B.t4 304.077
R1262 B.n171 B.t9 257.926
R1263 B.n165 B.t0 257.926
R1264 B.n61 B.t6 257.926
R1265 B.n54 B.t3 257.926
R1266 B.n861 B.n860 256.663
R1267 B.n860 B.n859 235.042
R1268 B.n860 B.n2 235.042
R1269 B.n329 B.n328 163.367
R1270 B.n329 B.n186 163.367
R1271 B.n333 B.n186 163.367
R1272 B.n334 B.n333 163.367
R1273 B.n335 B.n334 163.367
R1274 B.n335 B.n184 163.367
R1275 B.n339 B.n184 163.367
R1276 B.n340 B.n339 163.367
R1277 B.n341 B.n340 163.367
R1278 B.n341 B.n182 163.367
R1279 B.n345 B.n182 163.367
R1280 B.n346 B.n345 163.367
R1281 B.n347 B.n346 163.367
R1282 B.n347 B.n180 163.367
R1283 B.n351 B.n180 163.367
R1284 B.n352 B.n351 163.367
R1285 B.n353 B.n352 163.367
R1286 B.n353 B.n178 163.367
R1287 B.n357 B.n178 163.367
R1288 B.n358 B.n357 163.367
R1289 B.n359 B.n358 163.367
R1290 B.n359 B.n176 163.367
R1291 B.n363 B.n176 163.367
R1292 B.n364 B.n363 163.367
R1293 B.n365 B.n364 163.367
R1294 B.n365 B.n174 163.367
R1295 B.n369 B.n174 163.367
R1296 B.n370 B.n369 163.367
R1297 B.n371 B.n370 163.367
R1298 B.n371 B.n170 163.367
R1299 B.n376 B.n170 163.367
R1300 B.n377 B.n376 163.367
R1301 B.n378 B.n377 163.367
R1302 B.n378 B.n168 163.367
R1303 B.n382 B.n168 163.367
R1304 B.n383 B.n382 163.367
R1305 B.n384 B.n383 163.367
R1306 B.n384 B.n164 163.367
R1307 B.n389 B.n164 163.367
R1308 B.n390 B.n389 163.367
R1309 B.n391 B.n390 163.367
R1310 B.n391 B.n162 163.367
R1311 B.n395 B.n162 163.367
R1312 B.n396 B.n395 163.367
R1313 B.n397 B.n396 163.367
R1314 B.n397 B.n160 163.367
R1315 B.n401 B.n160 163.367
R1316 B.n402 B.n401 163.367
R1317 B.n403 B.n402 163.367
R1318 B.n403 B.n158 163.367
R1319 B.n407 B.n158 163.367
R1320 B.n408 B.n407 163.367
R1321 B.n409 B.n408 163.367
R1322 B.n409 B.n156 163.367
R1323 B.n413 B.n156 163.367
R1324 B.n414 B.n413 163.367
R1325 B.n415 B.n414 163.367
R1326 B.n415 B.n154 163.367
R1327 B.n419 B.n154 163.367
R1328 B.n420 B.n419 163.367
R1329 B.n421 B.n420 163.367
R1330 B.n421 B.n152 163.367
R1331 B.n425 B.n152 163.367
R1332 B.n426 B.n425 163.367
R1333 B.n427 B.n426 163.367
R1334 B.n427 B.n150 163.367
R1335 B.n431 B.n150 163.367
R1336 B.n432 B.n431 163.367
R1337 B.n648 B.n647 163.367
R1338 B.n647 B.n78 163.367
R1339 B.n643 B.n78 163.367
R1340 B.n643 B.n642 163.367
R1341 B.n642 B.n641 163.367
R1342 B.n641 B.n80 163.367
R1343 B.n637 B.n80 163.367
R1344 B.n637 B.n636 163.367
R1345 B.n636 B.n635 163.367
R1346 B.n635 B.n82 163.367
R1347 B.n631 B.n82 163.367
R1348 B.n631 B.n630 163.367
R1349 B.n630 B.n629 163.367
R1350 B.n629 B.n84 163.367
R1351 B.n625 B.n84 163.367
R1352 B.n625 B.n624 163.367
R1353 B.n624 B.n623 163.367
R1354 B.n623 B.n86 163.367
R1355 B.n619 B.n86 163.367
R1356 B.n619 B.n618 163.367
R1357 B.n618 B.n617 163.367
R1358 B.n617 B.n88 163.367
R1359 B.n613 B.n88 163.367
R1360 B.n613 B.n612 163.367
R1361 B.n612 B.n611 163.367
R1362 B.n611 B.n90 163.367
R1363 B.n607 B.n90 163.367
R1364 B.n607 B.n606 163.367
R1365 B.n606 B.n605 163.367
R1366 B.n605 B.n92 163.367
R1367 B.n601 B.n92 163.367
R1368 B.n601 B.n600 163.367
R1369 B.n600 B.n599 163.367
R1370 B.n599 B.n94 163.367
R1371 B.n595 B.n94 163.367
R1372 B.n595 B.n594 163.367
R1373 B.n594 B.n593 163.367
R1374 B.n593 B.n96 163.367
R1375 B.n589 B.n96 163.367
R1376 B.n589 B.n588 163.367
R1377 B.n588 B.n587 163.367
R1378 B.n587 B.n98 163.367
R1379 B.n583 B.n98 163.367
R1380 B.n583 B.n582 163.367
R1381 B.n582 B.n581 163.367
R1382 B.n581 B.n100 163.367
R1383 B.n577 B.n100 163.367
R1384 B.n577 B.n576 163.367
R1385 B.n576 B.n575 163.367
R1386 B.n575 B.n102 163.367
R1387 B.n571 B.n102 163.367
R1388 B.n571 B.n570 163.367
R1389 B.n570 B.n569 163.367
R1390 B.n569 B.n104 163.367
R1391 B.n565 B.n104 163.367
R1392 B.n565 B.n564 163.367
R1393 B.n564 B.n563 163.367
R1394 B.n563 B.n106 163.367
R1395 B.n559 B.n106 163.367
R1396 B.n559 B.n558 163.367
R1397 B.n558 B.n557 163.367
R1398 B.n557 B.n108 163.367
R1399 B.n553 B.n108 163.367
R1400 B.n553 B.n552 163.367
R1401 B.n552 B.n551 163.367
R1402 B.n551 B.n110 163.367
R1403 B.n547 B.n110 163.367
R1404 B.n547 B.n546 163.367
R1405 B.n546 B.n545 163.367
R1406 B.n545 B.n112 163.367
R1407 B.n541 B.n112 163.367
R1408 B.n541 B.n540 163.367
R1409 B.n540 B.n539 163.367
R1410 B.n539 B.n114 163.367
R1411 B.n535 B.n114 163.367
R1412 B.n535 B.n534 163.367
R1413 B.n534 B.n533 163.367
R1414 B.n533 B.n116 163.367
R1415 B.n529 B.n116 163.367
R1416 B.n529 B.n528 163.367
R1417 B.n528 B.n527 163.367
R1418 B.n527 B.n118 163.367
R1419 B.n523 B.n118 163.367
R1420 B.n523 B.n522 163.367
R1421 B.n522 B.n521 163.367
R1422 B.n521 B.n120 163.367
R1423 B.n517 B.n120 163.367
R1424 B.n517 B.n516 163.367
R1425 B.n516 B.n515 163.367
R1426 B.n515 B.n122 163.367
R1427 B.n511 B.n122 163.367
R1428 B.n511 B.n510 163.367
R1429 B.n510 B.n509 163.367
R1430 B.n509 B.n124 163.367
R1431 B.n505 B.n124 163.367
R1432 B.n505 B.n504 163.367
R1433 B.n504 B.n503 163.367
R1434 B.n503 B.n126 163.367
R1435 B.n499 B.n126 163.367
R1436 B.n499 B.n498 163.367
R1437 B.n498 B.n497 163.367
R1438 B.n497 B.n128 163.367
R1439 B.n493 B.n128 163.367
R1440 B.n493 B.n492 163.367
R1441 B.n492 B.n491 163.367
R1442 B.n491 B.n130 163.367
R1443 B.n487 B.n130 163.367
R1444 B.n487 B.n486 163.367
R1445 B.n486 B.n485 163.367
R1446 B.n485 B.n132 163.367
R1447 B.n481 B.n132 163.367
R1448 B.n481 B.n480 163.367
R1449 B.n480 B.n479 163.367
R1450 B.n479 B.n134 163.367
R1451 B.n475 B.n134 163.367
R1452 B.n475 B.n474 163.367
R1453 B.n474 B.n473 163.367
R1454 B.n473 B.n136 163.367
R1455 B.n469 B.n136 163.367
R1456 B.n469 B.n468 163.367
R1457 B.n468 B.n467 163.367
R1458 B.n467 B.n138 163.367
R1459 B.n463 B.n138 163.367
R1460 B.n463 B.n462 163.367
R1461 B.n462 B.n461 163.367
R1462 B.n461 B.n140 163.367
R1463 B.n457 B.n140 163.367
R1464 B.n457 B.n456 163.367
R1465 B.n456 B.n455 163.367
R1466 B.n455 B.n142 163.367
R1467 B.n451 B.n142 163.367
R1468 B.n451 B.n450 163.367
R1469 B.n450 B.n449 163.367
R1470 B.n449 B.n144 163.367
R1471 B.n445 B.n144 163.367
R1472 B.n445 B.n444 163.367
R1473 B.n444 B.n443 163.367
R1474 B.n443 B.n146 163.367
R1475 B.n439 B.n146 163.367
R1476 B.n439 B.n438 163.367
R1477 B.n438 B.n437 163.367
R1478 B.n437 B.n148 163.367
R1479 B.n433 B.n148 163.367
R1480 B.n752 B.n751 163.367
R1481 B.n751 B.n750 163.367
R1482 B.n750 B.n39 163.367
R1483 B.n746 B.n39 163.367
R1484 B.n746 B.n745 163.367
R1485 B.n745 B.n744 163.367
R1486 B.n744 B.n41 163.367
R1487 B.n740 B.n41 163.367
R1488 B.n740 B.n739 163.367
R1489 B.n739 B.n738 163.367
R1490 B.n738 B.n43 163.367
R1491 B.n734 B.n43 163.367
R1492 B.n734 B.n733 163.367
R1493 B.n733 B.n732 163.367
R1494 B.n732 B.n45 163.367
R1495 B.n728 B.n45 163.367
R1496 B.n728 B.n727 163.367
R1497 B.n727 B.n726 163.367
R1498 B.n726 B.n47 163.367
R1499 B.n722 B.n47 163.367
R1500 B.n722 B.n721 163.367
R1501 B.n721 B.n720 163.367
R1502 B.n720 B.n49 163.367
R1503 B.n716 B.n49 163.367
R1504 B.n716 B.n715 163.367
R1505 B.n715 B.n714 163.367
R1506 B.n714 B.n51 163.367
R1507 B.n710 B.n51 163.367
R1508 B.n710 B.n709 163.367
R1509 B.n709 B.n708 163.367
R1510 B.n708 B.n53 163.367
R1511 B.n704 B.n53 163.367
R1512 B.n704 B.n703 163.367
R1513 B.n703 B.n702 163.367
R1514 B.n702 B.n58 163.367
R1515 B.n698 B.n58 163.367
R1516 B.n698 B.n697 163.367
R1517 B.n697 B.n696 163.367
R1518 B.n696 B.n60 163.367
R1519 B.n691 B.n60 163.367
R1520 B.n691 B.n690 163.367
R1521 B.n690 B.n689 163.367
R1522 B.n689 B.n64 163.367
R1523 B.n685 B.n64 163.367
R1524 B.n685 B.n684 163.367
R1525 B.n684 B.n683 163.367
R1526 B.n683 B.n66 163.367
R1527 B.n679 B.n66 163.367
R1528 B.n679 B.n678 163.367
R1529 B.n678 B.n677 163.367
R1530 B.n677 B.n68 163.367
R1531 B.n673 B.n68 163.367
R1532 B.n673 B.n672 163.367
R1533 B.n672 B.n671 163.367
R1534 B.n671 B.n70 163.367
R1535 B.n667 B.n70 163.367
R1536 B.n667 B.n666 163.367
R1537 B.n666 B.n665 163.367
R1538 B.n665 B.n72 163.367
R1539 B.n661 B.n72 163.367
R1540 B.n661 B.n660 163.367
R1541 B.n660 B.n659 163.367
R1542 B.n659 B.n74 163.367
R1543 B.n655 B.n74 163.367
R1544 B.n655 B.n654 163.367
R1545 B.n654 B.n653 163.367
R1546 B.n653 B.n76 163.367
R1547 B.n649 B.n76 163.367
R1548 B.n756 B.n37 163.367
R1549 B.n757 B.n756 163.367
R1550 B.n758 B.n757 163.367
R1551 B.n758 B.n35 163.367
R1552 B.n762 B.n35 163.367
R1553 B.n763 B.n762 163.367
R1554 B.n764 B.n763 163.367
R1555 B.n764 B.n33 163.367
R1556 B.n768 B.n33 163.367
R1557 B.n769 B.n768 163.367
R1558 B.n770 B.n769 163.367
R1559 B.n770 B.n31 163.367
R1560 B.n774 B.n31 163.367
R1561 B.n775 B.n774 163.367
R1562 B.n776 B.n775 163.367
R1563 B.n776 B.n29 163.367
R1564 B.n780 B.n29 163.367
R1565 B.n781 B.n780 163.367
R1566 B.n782 B.n781 163.367
R1567 B.n782 B.n27 163.367
R1568 B.n786 B.n27 163.367
R1569 B.n787 B.n786 163.367
R1570 B.n788 B.n787 163.367
R1571 B.n788 B.n25 163.367
R1572 B.n792 B.n25 163.367
R1573 B.n793 B.n792 163.367
R1574 B.n794 B.n793 163.367
R1575 B.n794 B.n23 163.367
R1576 B.n798 B.n23 163.367
R1577 B.n799 B.n798 163.367
R1578 B.n800 B.n799 163.367
R1579 B.n800 B.n21 163.367
R1580 B.n804 B.n21 163.367
R1581 B.n805 B.n804 163.367
R1582 B.n806 B.n805 163.367
R1583 B.n806 B.n19 163.367
R1584 B.n810 B.n19 163.367
R1585 B.n811 B.n810 163.367
R1586 B.n812 B.n811 163.367
R1587 B.n812 B.n17 163.367
R1588 B.n816 B.n17 163.367
R1589 B.n817 B.n816 163.367
R1590 B.n818 B.n817 163.367
R1591 B.n818 B.n15 163.367
R1592 B.n822 B.n15 163.367
R1593 B.n823 B.n822 163.367
R1594 B.n824 B.n823 163.367
R1595 B.n824 B.n13 163.367
R1596 B.n828 B.n13 163.367
R1597 B.n829 B.n828 163.367
R1598 B.n830 B.n829 163.367
R1599 B.n830 B.n11 163.367
R1600 B.n834 B.n11 163.367
R1601 B.n835 B.n834 163.367
R1602 B.n836 B.n835 163.367
R1603 B.n836 B.n9 163.367
R1604 B.n840 B.n9 163.367
R1605 B.n841 B.n840 163.367
R1606 B.n842 B.n841 163.367
R1607 B.n842 B.n7 163.367
R1608 B.n846 B.n7 163.367
R1609 B.n847 B.n846 163.367
R1610 B.n848 B.n847 163.367
R1611 B.n848 B.n5 163.367
R1612 B.n852 B.n5 163.367
R1613 B.n853 B.n852 163.367
R1614 B.n854 B.n853 163.367
R1615 B.n854 B.n3 163.367
R1616 B.n858 B.n3 163.367
R1617 B.n859 B.n858 163.367
R1618 B.n222 B.n2 163.367
R1619 B.n225 B.n222 163.367
R1620 B.n226 B.n225 163.367
R1621 B.n227 B.n226 163.367
R1622 B.n227 B.n220 163.367
R1623 B.n231 B.n220 163.367
R1624 B.n232 B.n231 163.367
R1625 B.n233 B.n232 163.367
R1626 B.n233 B.n218 163.367
R1627 B.n237 B.n218 163.367
R1628 B.n238 B.n237 163.367
R1629 B.n239 B.n238 163.367
R1630 B.n239 B.n216 163.367
R1631 B.n243 B.n216 163.367
R1632 B.n244 B.n243 163.367
R1633 B.n245 B.n244 163.367
R1634 B.n245 B.n214 163.367
R1635 B.n249 B.n214 163.367
R1636 B.n250 B.n249 163.367
R1637 B.n251 B.n250 163.367
R1638 B.n251 B.n212 163.367
R1639 B.n255 B.n212 163.367
R1640 B.n256 B.n255 163.367
R1641 B.n257 B.n256 163.367
R1642 B.n257 B.n210 163.367
R1643 B.n261 B.n210 163.367
R1644 B.n262 B.n261 163.367
R1645 B.n263 B.n262 163.367
R1646 B.n263 B.n208 163.367
R1647 B.n267 B.n208 163.367
R1648 B.n268 B.n267 163.367
R1649 B.n269 B.n268 163.367
R1650 B.n269 B.n206 163.367
R1651 B.n273 B.n206 163.367
R1652 B.n274 B.n273 163.367
R1653 B.n275 B.n274 163.367
R1654 B.n275 B.n204 163.367
R1655 B.n279 B.n204 163.367
R1656 B.n280 B.n279 163.367
R1657 B.n281 B.n280 163.367
R1658 B.n281 B.n202 163.367
R1659 B.n285 B.n202 163.367
R1660 B.n286 B.n285 163.367
R1661 B.n287 B.n286 163.367
R1662 B.n287 B.n200 163.367
R1663 B.n291 B.n200 163.367
R1664 B.n292 B.n291 163.367
R1665 B.n293 B.n292 163.367
R1666 B.n293 B.n198 163.367
R1667 B.n297 B.n198 163.367
R1668 B.n298 B.n297 163.367
R1669 B.n299 B.n298 163.367
R1670 B.n299 B.n196 163.367
R1671 B.n303 B.n196 163.367
R1672 B.n304 B.n303 163.367
R1673 B.n305 B.n304 163.367
R1674 B.n305 B.n194 163.367
R1675 B.n309 B.n194 163.367
R1676 B.n310 B.n309 163.367
R1677 B.n311 B.n310 163.367
R1678 B.n311 B.n192 163.367
R1679 B.n315 B.n192 163.367
R1680 B.n316 B.n315 163.367
R1681 B.n317 B.n316 163.367
R1682 B.n317 B.n190 163.367
R1683 B.n321 B.n190 163.367
R1684 B.n322 B.n321 163.367
R1685 B.n323 B.n322 163.367
R1686 B.n323 B.n188 163.367
R1687 B.n327 B.n188 163.367
R1688 B.n172 B.n171 83.7823
R1689 B.n166 B.n165 83.7823
R1690 B.n62 B.n61 83.7823
R1691 B.n55 B.n54 83.7823
R1692 B.n373 B.n172 59.5399
R1693 B.n387 B.n166 59.5399
R1694 B.n694 B.n62 59.5399
R1695 B.n56 B.n55 59.5399
R1696 B.n754 B.n753 36.059
R1697 B.n650 B.n77 36.059
R1698 B.n326 B.n187 36.059
R1699 B.n434 B.n149 36.059
R1700 B B.n861 18.0485
R1701 B.n755 B.n754 10.6151
R1702 B.n755 B.n36 10.6151
R1703 B.n759 B.n36 10.6151
R1704 B.n760 B.n759 10.6151
R1705 B.n761 B.n760 10.6151
R1706 B.n761 B.n34 10.6151
R1707 B.n765 B.n34 10.6151
R1708 B.n766 B.n765 10.6151
R1709 B.n767 B.n766 10.6151
R1710 B.n767 B.n32 10.6151
R1711 B.n771 B.n32 10.6151
R1712 B.n772 B.n771 10.6151
R1713 B.n773 B.n772 10.6151
R1714 B.n773 B.n30 10.6151
R1715 B.n777 B.n30 10.6151
R1716 B.n778 B.n777 10.6151
R1717 B.n779 B.n778 10.6151
R1718 B.n779 B.n28 10.6151
R1719 B.n783 B.n28 10.6151
R1720 B.n784 B.n783 10.6151
R1721 B.n785 B.n784 10.6151
R1722 B.n785 B.n26 10.6151
R1723 B.n789 B.n26 10.6151
R1724 B.n790 B.n789 10.6151
R1725 B.n791 B.n790 10.6151
R1726 B.n791 B.n24 10.6151
R1727 B.n795 B.n24 10.6151
R1728 B.n796 B.n795 10.6151
R1729 B.n797 B.n796 10.6151
R1730 B.n797 B.n22 10.6151
R1731 B.n801 B.n22 10.6151
R1732 B.n802 B.n801 10.6151
R1733 B.n803 B.n802 10.6151
R1734 B.n803 B.n20 10.6151
R1735 B.n807 B.n20 10.6151
R1736 B.n808 B.n807 10.6151
R1737 B.n809 B.n808 10.6151
R1738 B.n809 B.n18 10.6151
R1739 B.n813 B.n18 10.6151
R1740 B.n814 B.n813 10.6151
R1741 B.n815 B.n814 10.6151
R1742 B.n815 B.n16 10.6151
R1743 B.n819 B.n16 10.6151
R1744 B.n820 B.n819 10.6151
R1745 B.n821 B.n820 10.6151
R1746 B.n821 B.n14 10.6151
R1747 B.n825 B.n14 10.6151
R1748 B.n826 B.n825 10.6151
R1749 B.n827 B.n826 10.6151
R1750 B.n827 B.n12 10.6151
R1751 B.n831 B.n12 10.6151
R1752 B.n832 B.n831 10.6151
R1753 B.n833 B.n832 10.6151
R1754 B.n833 B.n10 10.6151
R1755 B.n837 B.n10 10.6151
R1756 B.n838 B.n837 10.6151
R1757 B.n839 B.n838 10.6151
R1758 B.n839 B.n8 10.6151
R1759 B.n843 B.n8 10.6151
R1760 B.n844 B.n843 10.6151
R1761 B.n845 B.n844 10.6151
R1762 B.n845 B.n6 10.6151
R1763 B.n849 B.n6 10.6151
R1764 B.n850 B.n849 10.6151
R1765 B.n851 B.n850 10.6151
R1766 B.n851 B.n4 10.6151
R1767 B.n855 B.n4 10.6151
R1768 B.n856 B.n855 10.6151
R1769 B.n857 B.n856 10.6151
R1770 B.n857 B.n0 10.6151
R1771 B.n753 B.n38 10.6151
R1772 B.n749 B.n38 10.6151
R1773 B.n749 B.n748 10.6151
R1774 B.n748 B.n747 10.6151
R1775 B.n747 B.n40 10.6151
R1776 B.n743 B.n40 10.6151
R1777 B.n743 B.n742 10.6151
R1778 B.n742 B.n741 10.6151
R1779 B.n741 B.n42 10.6151
R1780 B.n737 B.n42 10.6151
R1781 B.n737 B.n736 10.6151
R1782 B.n736 B.n735 10.6151
R1783 B.n735 B.n44 10.6151
R1784 B.n731 B.n44 10.6151
R1785 B.n731 B.n730 10.6151
R1786 B.n730 B.n729 10.6151
R1787 B.n729 B.n46 10.6151
R1788 B.n725 B.n46 10.6151
R1789 B.n725 B.n724 10.6151
R1790 B.n724 B.n723 10.6151
R1791 B.n723 B.n48 10.6151
R1792 B.n719 B.n48 10.6151
R1793 B.n719 B.n718 10.6151
R1794 B.n718 B.n717 10.6151
R1795 B.n717 B.n50 10.6151
R1796 B.n713 B.n50 10.6151
R1797 B.n713 B.n712 10.6151
R1798 B.n712 B.n711 10.6151
R1799 B.n711 B.n52 10.6151
R1800 B.n707 B.n706 10.6151
R1801 B.n706 B.n705 10.6151
R1802 B.n705 B.n57 10.6151
R1803 B.n701 B.n57 10.6151
R1804 B.n701 B.n700 10.6151
R1805 B.n700 B.n699 10.6151
R1806 B.n699 B.n59 10.6151
R1807 B.n695 B.n59 10.6151
R1808 B.n693 B.n692 10.6151
R1809 B.n692 B.n63 10.6151
R1810 B.n688 B.n63 10.6151
R1811 B.n688 B.n687 10.6151
R1812 B.n687 B.n686 10.6151
R1813 B.n686 B.n65 10.6151
R1814 B.n682 B.n65 10.6151
R1815 B.n682 B.n681 10.6151
R1816 B.n681 B.n680 10.6151
R1817 B.n680 B.n67 10.6151
R1818 B.n676 B.n67 10.6151
R1819 B.n676 B.n675 10.6151
R1820 B.n675 B.n674 10.6151
R1821 B.n674 B.n69 10.6151
R1822 B.n670 B.n69 10.6151
R1823 B.n670 B.n669 10.6151
R1824 B.n669 B.n668 10.6151
R1825 B.n668 B.n71 10.6151
R1826 B.n664 B.n71 10.6151
R1827 B.n664 B.n663 10.6151
R1828 B.n663 B.n662 10.6151
R1829 B.n662 B.n73 10.6151
R1830 B.n658 B.n73 10.6151
R1831 B.n658 B.n657 10.6151
R1832 B.n657 B.n656 10.6151
R1833 B.n656 B.n75 10.6151
R1834 B.n652 B.n75 10.6151
R1835 B.n652 B.n651 10.6151
R1836 B.n651 B.n650 10.6151
R1837 B.n646 B.n77 10.6151
R1838 B.n646 B.n645 10.6151
R1839 B.n645 B.n644 10.6151
R1840 B.n644 B.n79 10.6151
R1841 B.n640 B.n79 10.6151
R1842 B.n640 B.n639 10.6151
R1843 B.n639 B.n638 10.6151
R1844 B.n638 B.n81 10.6151
R1845 B.n634 B.n81 10.6151
R1846 B.n634 B.n633 10.6151
R1847 B.n633 B.n632 10.6151
R1848 B.n632 B.n83 10.6151
R1849 B.n628 B.n83 10.6151
R1850 B.n628 B.n627 10.6151
R1851 B.n627 B.n626 10.6151
R1852 B.n626 B.n85 10.6151
R1853 B.n622 B.n85 10.6151
R1854 B.n622 B.n621 10.6151
R1855 B.n621 B.n620 10.6151
R1856 B.n620 B.n87 10.6151
R1857 B.n616 B.n87 10.6151
R1858 B.n616 B.n615 10.6151
R1859 B.n615 B.n614 10.6151
R1860 B.n614 B.n89 10.6151
R1861 B.n610 B.n89 10.6151
R1862 B.n610 B.n609 10.6151
R1863 B.n609 B.n608 10.6151
R1864 B.n608 B.n91 10.6151
R1865 B.n604 B.n91 10.6151
R1866 B.n604 B.n603 10.6151
R1867 B.n603 B.n602 10.6151
R1868 B.n602 B.n93 10.6151
R1869 B.n598 B.n93 10.6151
R1870 B.n598 B.n597 10.6151
R1871 B.n597 B.n596 10.6151
R1872 B.n596 B.n95 10.6151
R1873 B.n592 B.n95 10.6151
R1874 B.n592 B.n591 10.6151
R1875 B.n591 B.n590 10.6151
R1876 B.n590 B.n97 10.6151
R1877 B.n586 B.n97 10.6151
R1878 B.n586 B.n585 10.6151
R1879 B.n585 B.n584 10.6151
R1880 B.n584 B.n99 10.6151
R1881 B.n580 B.n99 10.6151
R1882 B.n580 B.n579 10.6151
R1883 B.n579 B.n578 10.6151
R1884 B.n578 B.n101 10.6151
R1885 B.n574 B.n101 10.6151
R1886 B.n574 B.n573 10.6151
R1887 B.n573 B.n572 10.6151
R1888 B.n572 B.n103 10.6151
R1889 B.n568 B.n103 10.6151
R1890 B.n568 B.n567 10.6151
R1891 B.n567 B.n566 10.6151
R1892 B.n566 B.n105 10.6151
R1893 B.n562 B.n105 10.6151
R1894 B.n562 B.n561 10.6151
R1895 B.n561 B.n560 10.6151
R1896 B.n560 B.n107 10.6151
R1897 B.n556 B.n107 10.6151
R1898 B.n556 B.n555 10.6151
R1899 B.n555 B.n554 10.6151
R1900 B.n554 B.n109 10.6151
R1901 B.n550 B.n109 10.6151
R1902 B.n550 B.n549 10.6151
R1903 B.n549 B.n548 10.6151
R1904 B.n548 B.n111 10.6151
R1905 B.n544 B.n111 10.6151
R1906 B.n544 B.n543 10.6151
R1907 B.n543 B.n542 10.6151
R1908 B.n542 B.n113 10.6151
R1909 B.n538 B.n113 10.6151
R1910 B.n538 B.n537 10.6151
R1911 B.n537 B.n536 10.6151
R1912 B.n536 B.n115 10.6151
R1913 B.n532 B.n115 10.6151
R1914 B.n532 B.n531 10.6151
R1915 B.n531 B.n530 10.6151
R1916 B.n530 B.n117 10.6151
R1917 B.n526 B.n117 10.6151
R1918 B.n526 B.n525 10.6151
R1919 B.n525 B.n524 10.6151
R1920 B.n524 B.n119 10.6151
R1921 B.n520 B.n119 10.6151
R1922 B.n520 B.n519 10.6151
R1923 B.n519 B.n518 10.6151
R1924 B.n518 B.n121 10.6151
R1925 B.n514 B.n121 10.6151
R1926 B.n514 B.n513 10.6151
R1927 B.n513 B.n512 10.6151
R1928 B.n512 B.n123 10.6151
R1929 B.n508 B.n123 10.6151
R1930 B.n508 B.n507 10.6151
R1931 B.n507 B.n506 10.6151
R1932 B.n506 B.n125 10.6151
R1933 B.n502 B.n125 10.6151
R1934 B.n502 B.n501 10.6151
R1935 B.n501 B.n500 10.6151
R1936 B.n500 B.n127 10.6151
R1937 B.n496 B.n127 10.6151
R1938 B.n496 B.n495 10.6151
R1939 B.n495 B.n494 10.6151
R1940 B.n494 B.n129 10.6151
R1941 B.n490 B.n129 10.6151
R1942 B.n490 B.n489 10.6151
R1943 B.n489 B.n488 10.6151
R1944 B.n488 B.n131 10.6151
R1945 B.n484 B.n131 10.6151
R1946 B.n484 B.n483 10.6151
R1947 B.n483 B.n482 10.6151
R1948 B.n482 B.n133 10.6151
R1949 B.n478 B.n133 10.6151
R1950 B.n478 B.n477 10.6151
R1951 B.n477 B.n476 10.6151
R1952 B.n476 B.n135 10.6151
R1953 B.n472 B.n135 10.6151
R1954 B.n472 B.n471 10.6151
R1955 B.n471 B.n470 10.6151
R1956 B.n470 B.n137 10.6151
R1957 B.n466 B.n137 10.6151
R1958 B.n466 B.n465 10.6151
R1959 B.n465 B.n464 10.6151
R1960 B.n464 B.n139 10.6151
R1961 B.n460 B.n139 10.6151
R1962 B.n460 B.n459 10.6151
R1963 B.n459 B.n458 10.6151
R1964 B.n458 B.n141 10.6151
R1965 B.n454 B.n141 10.6151
R1966 B.n454 B.n453 10.6151
R1967 B.n453 B.n452 10.6151
R1968 B.n452 B.n143 10.6151
R1969 B.n448 B.n143 10.6151
R1970 B.n448 B.n447 10.6151
R1971 B.n447 B.n446 10.6151
R1972 B.n446 B.n145 10.6151
R1973 B.n442 B.n145 10.6151
R1974 B.n442 B.n441 10.6151
R1975 B.n441 B.n440 10.6151
R1976 B.n440 B.n147 10.6151
R1977 B.n436 B.n147 10.6151
R1978 B.n436 B.n435 10.6151
R1979 B.n435 B.n434 10.6151
R1980 B.n223 B.n1 10.6151
R1981 B.n224 B.n223 10.6151
R1982 B.n224 B.n221 10.6151
R1983 B.n228 B.n221 10.6151
R1984 B.n229 B.n228 10.6151
R1985 B.n230 B.n229 10.6151
R1986 B.n230 B.n219 10.6151
R1987 B.n234 B.n219 10.6151
R1988 B.n235 B.n234 10.6151
R1989 B.n236 B.n235 10.6151
R1990 B.n236 B.n217 10.6151
R1991 B.n240 B.n217 10.6151
R1992 B.n241 B.n240 10.6151
R1993 B.n242 B.n241 10.6151
R1994 B.n242 B.n215 10.6151
R1995 B.n246 B.n215 10.6151
R1996 B.n247 B.n246 10.6151
R1997 B.n248 B.n247 10.6151
R1998 B.n248 B.n213 10.6151
R1999 B.n252 B.n213 10.6151
R2000 B.n253 B.n252 10.6151
R2001 B.n254 B.n253 10.6151
R2002 B.n254 B.n211 10.6151
R2003 B.n258 B.n211 10.6151
R2004 B.n259 B.n258 10.6151
R2005 B.n260 B.n259 10.6151
R2006 B.n260 B.n209 10.6151
R2007 B.n264 B.n209 10.6151
R2008 B.n265 B.n264 10.6151
R2009 B.n266 B.n265 10.6151
R2010 B.n266 B.n207 10.6151
R2011 B.n270 B.n207 10.6151
R2012 B.n271 B.n270 10.6151
R2013 B.n272 B.n271 10.6151
R2014 B.n272 B.n205 10.6151
R2015 B.n276 B.n205 10.6151
R2016 B.n277 B.n276 10.6151
R2017 B.n278 B.n277 10.6151
R2018 B.n278 B.n203 10.6151
R2019 B.n282 B.n203 10.6151
R2020 B.n283 B.n282 10.6151
R2021 B.n284 B.n283 10.6151
R2022 B.n284 B.n201 10.6151
R2023 B.n288 B.n201 10.6151
R2024 B.n289 B.n288 10.6151
R2025 B.n290 B.n289 10.6151
R2026 B.n290 B.n199 10.6151
R2027 B.n294 B.n199 10.6151
R2028 B.n295 B.n294 10.6151
R2029 B.n296 B.n295 10.6151
R2030 B.n296 B.n197 10.6151
R2031 B.n300 B.n197 10.6151
R2032 B.n301 B.n300 10.6151
R2033 B.n302 B.n301 10.6151
R2034 B.n302 B.n195 10.6151
R2035 B.n306 B.n195 10.6151
R2036 B.n307 B.n306 10.6151
R2037 B.n308 B.n307 10.6151
R2038 B.n308 B.n193 10.6151
R2039 B.n312 B.n193 10.6151
R2040 B.n313 B.n312 10.6151
R2041 B.n314 B.n313 10.6151
R2042 B.n314 B.n191 10.6151
R2043 B.n318 B.n191 10.6151
R2044 B.n319 B.n318 10.6151
R2045 B.n320 B.n319 10.6151
R2046 B.n320 B.n189 10.6151
R2047 B.n324 B.n189 10.6151
R2048 B.n325 B.n324 10.6151
R2049 B.n326 B.n325 10.6151
R2050 B.n330 B.n187 10.6151
R2051 B.n331 B.n330 10.6151
R2052 B.n332 B.n331 10.6151
R2053 B.n332 B.n185 10.6151
R2054 B.n336 B.n185 10.6151
R2055 B.n337 B.n336 10.6151
R2056 B.n338 B.n337 10.6151
R2057 B.n338 B.n183 10.6151
R2058 B.n342 B.n183 10.6151
R2059 B.n343 B.n342 10.6151
R2060 B.n344 B.n343 10.6151
R2061 B.n344 B.n181 10.6151
R2062 B.n348 B.n181 10.6151
R2063 B.n349 B.n348 10.6151
R2064 B.n350 B.n349 10.6151
R2065 B.n350 B.n179 10.6151
R2066 B.n354 B.n179 10.6151
R2067 B.n355 B.n354 10.6151
R2068 B.n356 B.n355 10.6151
R2069 B.n356 B.n177 10.6151
R2070 B.n360 B.n177 10.6151
R2071 B.n361 B.n360 10.6151
R2072 B.n362 B.n361 10.6151
R2073 B.n362 B.n175 10.6151
R2074 B.n366 B.n175 10.6151
R2075 B.n367 B.n366 10.6151
R2076 B.n368 B.n367 10.6151
R2077 B.n368 B.n173 10.6151
R2078 B.n372 B.n173 10.6151
R2079 B.n375 B.n374 10.6151
R2080 B.n375 B.n169 10.6151
R2081 B.n379 B.n169 10.6151
R2082 B.n380 B.n379 10.6151
R2083 B.n381 B.n380 10.6151
R2084 B.n381 B.n167 10.6151
R2085 B.n385 B.n167 10.6151
R2086 B.n386 B.n385 10.6151
R2087 B.n388 B.n163 10.6151
R2088 B.n392 B.n163 10.6151
R2089 B.n393 B.n392 10.6151
R2090 B.n394 B.n393 10.6151
R2091 B.n394 B.n161 10.6151
R2092 B.n398 B.n161 10.6151
R2093 B.n399 B.n398 10.6151
R2094 B.n400 B.n399 10.6151
R2095 B.n400 B.n159 10.6151
R2096 B.n404 B.n159 10.6151
R2097 B.n405 B.n404 10.6151
R2098 B.n406 B.n405 10.6151
R2099 B.n406 B.n157 10.6151
R2100 B.n410 B.n157 10.6151
R2101 B.n411 B.n410 10.6151
R2102 B.n412 B.n411 10.6151
R2103 B.n412 B.n155 10.6151
R2104 B.n416 B.n155 10.6151
R2105 B.n417 B.n416 10.6151
R2106 B.n418 B.n417 10.6151
R2107 B.n418 B.n153 10.6151
R2108 B.n422 B.n153 10.6151
R2109 B.n423 B.n422 10.6151
R2110 B.n424 B.n423 10.6151
R2111 B.n424 B.n151 10.6151
R2112 B.n428 B.n151 10.6151
R2113 B.n429 B.n428 10.6151
R2114 B.n430 B.n429 10.6151
R2115 B.n430 B.n149 10.6151
R2116 B.n861 B.n0 8.11757
R2117 B.n861 B.n1 8.11757
R2118 B.n707 B.n56 6.5566
R2119 B.n695 B.n694 6.5566
R2120 B.n374 B.n373 6.5566
R2121 B.n387 B.n386 6.5566
R2122 B.n56 B.n52 4.05904
R2123 B.n694 B.n693 4.05904
R2124 B.n373 B.n372 4.05904
R2125 B.n388 B.n387 4.05904
C0 VDD1 VN 0.154728f
C1 VP VDD2 0.668069f
C2 w_n5290_n2572# B 11.127f
C3 VN VP 8.61824f
C4 VDD2 VTAIL 7.71095f
C5 VN VTAIL 7.44595f
C6 VDD1 w_n5290_n2572# 2.29589f
C7 VN VDD2 6.382f
C8 VP w_n5290_n2572# 11.754701f
C9 VDD1 B 1.967f
C10 w_n5290_n2572# VTAIL 3.46621f
C11 VP B 2.67246f
C12 VTAIL B 4.15291f
C13 w_n5290_n2572# VDD2 2.4689f
C14 VN w_n5290_n2572# 11.0638f
C15 VDD1 VP 6.89324f
C16 VDD2 B 2.10676f
C17 VN B 1.50695f
C18 VDD1 VTAIL 7.64722f
C19 VP VTAIL 7.46006f
C20 VDD1 VDD2 2.5005f
C21 VDD2 VSUBS 2.560182f
C22 VDD1 VSUBS 3.28771f
C23 VTAIL VSUBS 1.450732f
C24 VN VSUBS 8.63107f
C25 VP VSUBS 4.898775f
C26 B VSUBS 6.216903f
C27 w_n5290_n2572# VSUBS 0.168793p
C28 B.n0 VSUBS 0.00809f
C29 B.n1 VSUBS 0.00809f
C30 B.n2 VSUBS 0.011965f
C31 B.n3 VSUBS 0.009169f
C32 B.n4 VSUBS 0.009169f
C33 B.n5 VSUBS 0.009169f
C34 B.n6 VSUBS 0.009169f
C35 B.n7 VSUBS 0.009169f
C36 B.n8 VSUBS 0.009169f
C37 B.n9 VSUBS 0.009169f
C38 B.n10 VSUBS 0.009169f
C39 B.n11 VSUBS 0.009169f
C40 B.n12 VSUBS 0.009169f
C41 B.n13 VSUBS 0.009169f
C42 B.n14 VSUBS 0.009169f
C43 B.n15 VSUBS 0.009169f
C44 B.n16 VSUBS 0.009169f
C45 B.n17 VSUBS 0.009169f
C46 B.n18 VSUBS 0.009169f
C47 B.n19 VSUBS 0.009169f
C48 B.n20 VSUBS 0.009169f
C49 B.n21 VSUBS 0.009169f
C50 B.n22 VSUBS 0.009169f
C51 B.n23 VSUBS 0.009169f
C52 B.n24 VSUBS 0.009169f
C53 B.n25 VSUBS 0.009169f
C54 B.n26 VSUBS 0.009169f
C55 B.n27 VSUBS 0.009169f
C56 B.n28 VSUBS 0.009169f
C57 B.n29 VSUBS 0.009169f
C58 B.n30 VSUBS 0.009169f
C59 B.n31 VSUBS 0.009169f
C60 B.n32 VSUBS 0.009169f
C61 B.n33 VSUBS 0.009169f
C62 B.n34 VSUBS 0.009169f
C63 B.n35 VSUBS 0.009169f
C64 B.n36 VSUBS 0.009169f
C65 B.n37 VSUBS 0.022503f
C66 B.n38 VSUBS 0.009169f
C67 B.n39 VSUBS 0.009169f
C68 B.n40 VSUBS 0.009169f
C69 B.n41 VSUBS 0.009169f
C70 B.n42 VSUBS 0.009169f
C71 B.n43 VSUBS 0.009169f
C72 B.n44 VSUBS 0.009169f
C73 B.n45 VSUBS 0.009169f
C74 B.n46 VSUBS 0.009169f
C75 B.n47 VSUBS 0.009169f
C76 B.n48 VSUBS 0.009169f
C77 B.n49 VSUBS 0.009169f
C78 B.n50 VSUBS 0.009169f
C79 B.n51 VSUBS 0.009169f
C80 B.n52 VSUBS 0.006337f
C81 B.n53 VSUBS 0.009169f
C82 B.t4 VSUBS 0.166441f
C83 B.t5 VSUBS 0.219537f
C84 B.t3 VSUBS 1.99672f
C85 B.n54 VSUBS 0.354724f
C86 B.n55 VSUBS 0.258879f
C87 B.n56 VSUBS 0.021243f
C88 B.n57 VSUBS 0.009169f
C89 B.n58 VSUBS 0.009169f
C90 B.n59 VSUBS 0.009169f
C91 B.n60 VSUBS 0.009169f
C92 B.t7 VSUBS 0.166444f
C93 B.t8 VSUBS 0.219539f
C94 B.t6 VSUBS 1.99672f
C95 B.n61 VSUBS 0.354721f
C96 B.n62 VSUBS 0.258876f
C97 B.n63 VSUBS 0.009169f
C98 B.n64 VSUBS 0.009169f
C99 B.n65 VSUBS 0.009169f
C100 B.n66 VSUBS 0.009169f
C101 B.n67 VSUBS 0.009169f
C102 B.n68 VSUBS 0.009169f
C103 B.n69 VSUBS 0.009169f
C104 B.n70 VSUBS 0.009169f
C105 B.n71 VSUBS 0.009169f
C106 B.n72 VSUBS 0.009169f
C107 B.n73 VSUBS 0.009169f
C108 B.n74 VSUBS 0.009169f
C109 B.n75 VSUBS 0.009169f
C110 B.n76 VSUBS 0.009169f
C111 B.n77 VSUBS 0.022503f
C112 B.n78 VSUBS 0.009169f
C113 B.n79 VSUBS 0.009169f
C114 B.n80 VSUBS 0.009169f
C115 B.n81 VSUBS 0.009169f
C116 B.n82 VSUBS 0.009169f
C117 B.n83 VSUBS 0.009169f
C118 B.n84 VSUBS 0.009169f
C119 B.n85 VSUBS 0.009169f
C120 B.n86 VSUBS 0.009169f
C121 B.n87 VSUBS 0.009169f
C122 B.n88 VSUBS 0.009169f
C123 B.n89 VSUBS 0.009169f
C124 B.n90 VSUBS 0.009169f
C125 B.n91 VSUBS 0.009169f
C126 B.n92 VSUBS 0.009169f
C127 B.n93 VSUBS 0.009169f
C128 B.n94 VSUBS 0.009169f
C129 B.n95 VSUBS 0.009169f
C130 B.n96 VSUBS 0.009169f
C131 B.n97 VSUBS 0.009169f
C132 B.n98 VSUBS 0.009169f
C133 B.n99 VSUBS 0.009169f
C134 B.n100 VSUBS 0.009169f
C135 B.n101 VSUBS 0.009169f
C136 B.n102 VSUBS 0.009169f
C137 B.n103 VSUBS 0.009169f
C138 B.n104 VSUBS 0.009169f
C139 B.n105 VSUBS 0.009169f
C140 B.n106 VSUBS 0.009169f
C141 B.n107 VSUBS 0.009169f
C142 B.n108 VSUBS 0.009169f
C143 B.n109 VSUBS 0.009169f
C144 B.n110 VSUBS 0.009169f
C145 B.n111 VSUBS 0.009169f
C146 B.n112 VSUBS 0.009169f
C147 B.n113 VSUBS 0.009169f
C148 B.n114 VSUBS 0.009169f
C149 B.n115 VSUBS 0.009169f
C150 B.n116 VSUBS 0.009169f
C151 B.n117 VSUBS 0.009169f
C152 B.n118 VSUBS 0.009169f
C153 B.n119 VSUBS 0.009169f
C154 B.n120 VSUBS 0.009169f
C155 B.n121 VSUBS 0.009169f
C156 B.n122 VSUBS 0.009169f
C157 B.n123 VSUBS 0.009169f
C158 B.n124 VSUBS 0.009169f
C159 B.n125 VSUBS 0.009169f
C160 B.n126 VSUBS 0.009169f
C161 B.n127 VSUBS 0.009169f
C162 B.n128 VSUBS 0.009169f
C163 B.n129 VSUBS 0.009169f
C164 B.n130 VSUBS 0.009169f
C165 B.n131 VSUBS 0.009169f
C166 B.n132 VSUBS 0.009169f
C167 B.n133 VSUBS 0.009169f
C168 B.n134 VSUBS 0.009169f
C169 B.n135 VSUBS 0.009169f
C170 B.n136 VSUBS 0.009169f
C171 B.n137 VSUBS 0.009169f
C172 B.n138 VSUBS 0.009169f
C173 B.n139 VSUBS 0.009169f
C174 B.n140 VSUBS 0.009169f
C175 B.n141 VSUBS 0.009169f
C176 B.n142 VSUBS 0.009169f
C177 B.n143 VSUBS 0.009169f
C178 B.n144 VSUBS 0.009169f
C179 B.n145 VSUBS 0.009169f
C180 B.n146 VSUBS 0.009169f
C181 B.n147 VSUBS 0.009169f
C182 B.n148 VSUBS 0.009169f
C183 B.n149 VSUBS 0.022359f
C184 B.n150 VSUBS 0.009169f
C185 B.n151 VSUBS 0.009169f
C186 B.n152 VSUBS 0.009169f
C187 B.n153 VSUBS 0.009169f
C188 B.n154 VSUBS 0.009169f
C189 B.n155 VSUBS 0.009169f
C190 B.n156 VSUBS 0.009169f
C191 B.n157 VSUBS 0.009169f
C192 B.n158 VSUBS 0.009169f
C193 B.n159 VSUBS 0.009169f
C194 B.n160 VSUBS 0.009169f
C195 B.n161 VSUBS 0.009169f
C196 B.n162 VSUBS 0.009169f
C197 B.n163 VSUBS 0.009169f
C198 B.n164 VSUBS 0.009169f
C199 B.t2 VSUBS 0.166444f
C200 B.t1 VSUBS 0.219539f
C201 B.t0 VSUBS 1.99672f
C202 B.n165 VSUBS 0.354721f
C203 B.n166 VSUBS 0.258876f
C204 B.n167 VSUBS 0.009169f
C205 B.n168 VSUBS 0.009169f
C206 B.n169 VSUBS 0.009169f
C207 B.n170 VSUBS 0.009169f
C208 B.t11 VSUBS 0.166441f
C209 B.t10 VSUBS 0.219537f
C210 B.t9 VSUBS 1.99672f
C211 B.n171 VSUBS 0.354724f
C212 B.n172 VSUBS 0.258879f
C213 B.n173 VSUBS 0.009169f
C214 B.n174 VSUBS 0.009169f
C215 B.n175 VSUBS 0.009169f
C216 B.n176 VSUBS 0.009169f
C217 B.n177 VSUBS 0.009169f
C218 B.n178 VSUBS 0.009169f
C219 B.n179 VSUBS 0.009169f
C220 B.n180 VSUBS 0.009169f
C221 B.n181 VSUBS 0.009169f
C222 B.n182 VSUBS 0.009169f
C223 B.n183 VSUBS 0.009169f
C224 B.n184 VSUBS 0.009169f
C225 B.n185 VSUBS 0.009169f
C226 B.n186 VSUBS 0.009169f
C227 B.n187 VSUBS 0.02334f
C228 B.n188 VSUBS 0.009169f
C229 B.n189 VSUBS 0.009169f
C230 B.n190 VSUBS 0.009169f
C231 B.n191 VSUBS 0.009169f
C232 B.n192 VSUBS 0.009169f
C233 B.n193 VSUBS 0.009169f
C234 B.n194 VSUBS 0.009169f
C235 B.n195 VSUBS 0.009169f
C236 B.n196 VSUBS 0.009169f
C237 B.n197 VSUBS 0.009169f
C238 B.n198 VSUBS 0.009169f
C239 B.n199 VSUBS 0.009169f
C240 B.n200 VSUBS 0.009169f
C241 B.n201 VSUBS 0.009169f
C242 B.n202 VSUBS 0.009169f
C243 B.n203 VSUBS 0.009169f
C244 B.n204 VSUBS 0.009169f
C245 B.n205 VSUBS 0.009169f
C246 B.n206 VSUBS 0.009169f
C247 B.n207 VSUBS 0.009169f
C248 B.n208 VSUBS 0.009169f
C249 B.n209 VSUBS 0.009169f
C250 B.n210 VSUBS 0.009169f
C251 B.n211 VSUBS 0.009169f
C252 B.n212 VSUBS 0.009169f
C253 B.n213 VSUBS 0.009169f
C254 B.n214 VSUBS 0.009169f
C255 B.n215 VSUBS 0.009169f
C256 B.n216 VSUBS 0.009169f
C257 B.n217 VSUBS 0.009169f
C258 B.n218 VSUBS 0.009169f
C259 B.n219 VSUBS 0.009169f
C260 B.n220 VSUBS 0.009169f
C261 B.n221 VSUBS 0.009169f
C262 B.n222 VSUBS 0.009169f
C263 B.n223 VSUBS 0.009169f
C264 B.n224 VSUBS 0.009169f
C265 B.n225 VSUBS 0.009169f
C266 B.n226 VSUBS 0.009169f
C267 B.n227 VSUBS 0.009169f
C268 B.n228 VSUBS 0.009169f
C269 B.n229 VSUBS 0.009169f
C270 B.n230 VSUBS 0.009169f
C271 B.n231 VSUBS 0.009169f
C272 B.n232 VSUBS 0.009169f
C273 B.n233 VSUBS 0.009169f
C274 B.n234 VSUBS 0.009169f
C275 B.n235 VSUBS 0.009169f
C276 B.n236 VSUBS 0.009169f
C277 B.n237 VSUBS 0.009169f
C278 B.n238 VSUBS 0.009169f
C279 B.n239 VSUBS 0.009169f
C280 B.n240 VSUBS 0.009169f
C281 B.n241 VSUBS 0.009169f
C282 B.n242 VSUBS 0.009169f
C283 B.n243 VSUBS 0.009169f
C284 B.n244 VSUBS 0.009169f
C285 B.n245 VSUBS 0.009169f
C286 B.n246 VSUBS 0.009169f
C287 B.n247 VSUBS 0.009169f
C288 B.n248 VSUBS 0.009169f
C289 B.n249 VSUBS 0.009169f
C290 B.n250 VSUBS 0.009169f
C291 B.n251 VSUBS 0.009169f
C292 B.n252 VSUBS 0.009169f
C293 B.n253 VSUBS 0.009169f
C294 B.n254 VSUBS 0.009169f
C295 B.n255 VSUBS 0.009169f
C296 B.n256 VSUBS 0.009169f
C297 B.n257 VSUBS 0.009169f
C298 B.n258 VSUBS 0.009169f
C299 B.n259 VSUBS 0.009169f
C300 B.n260 VSUBS 0.009169f
C301 B.n261 VSUBS 0.009169f
C302 B.n262 VSUBS 0.009169f
C303 B.n263 VSUBS 0.009169f
C304 B.n264 VSUBS 0.009169f
C305 B.n265 VSUBS 0.009169f
C306 B.n266 VSUBS 0.009169f
C307 B.n267 VSUBS 0.009169f
C308 B.n268 VSUBS 0.009169f
C309 B.n269 VSUBS 0.009169f
C310 B.n270 VSUBS 0.009169f
C311 B.n271 VSUBS 0.009169f
C312 B.n272 VSUBS 0.009169f
C313 B.n273 VSUBS 0.009169f
C314 B.n274 VSUBS 0.009169f
C315 B.n275 VSUBS 0.009169f
C316 B.n276 VSUBS 0.009169f
C317 B.n277 VSUBS 0.009169f
C318 B.n278 VSUBS 0.009169f
C319 B.n279 VSUBS 0.009169f
C320 B.n280 VSUBS 0.009169f
C321 B.n281 VSUBS 0.009169f
C322 B.n282 VSUBS 0.009169f
C323 B.n283 VSUBS 0.009169f
C324 B.n284 VSUBS 0.009169f
C325 B.n285 VSUBS 0.009169f
C326 B.n286 VSUBS 0.009169f
C327 B.n287 VSUBS 0.009169f
C328 B.n288 VSUBS 0.009169f
C329 B.n289 VSUBS 0.009169f
C330 B.n290 VSUBS 0.009169f
C331 B.n291 VSUBS 0.009169f
C332 B.n292 VSUBS 0.009169f
C333 B.n293 VSUBS 0.009169f
C334 B.n294 VSUBS 0.009169f
C335 B.n295 VSUBS 0.009169f
C336 B.n296 VSUBS 0.009169f
C337 B.n297 VSUBS 0.009169f
C338 B.n298 VSUBS 0.009169f
C339 B.n299 VSUBS 0.009169f
C340 B.n300 VSUBS 0.009169f
C341 B.n301 VSUBS 0.009169f
C342 B.n302 VSUBS 0.009169f
C343 B.n303 VSUBS 0.009169f
C344 B.n304 VSUBS 0.009169f
C345 B.n305 VSUBS 0.009169f
C346 B.n306 VSUBS 0.009169f
C347 B.n307 VSUBS 0.009169f
C348 B.n308 VSUBS 0.009169f
C349 B.n309 VSUBS 0.009169f
C350 B.n310 VSUBS 0.009169f
C351 B.n311 VSUBS 0.009169f
C352 B.n312 VSUBS 0.009169f
C353 B.n313 VSUBS 0.009169f
C354 B.n314 VSUBS 0.009169f
C355 B.n315 VSUBS 0.009169f
C356 B.n316 VSUBS 0.009169f
C357 B.n317 VSUBS 0.009169f
C358 B.n318 VSUBS 0.009169f
C359 B.n319 VSUBS 0.009169f
C360 B.n320 VSUBS 0.009169f
C361 B.n321 VSUBS 0.009169f
C362 B.n322 VSUBS 0.009169f
C363 B.n323 VSUBS 0.009169f
C364 B.n324 VSUBS 0.009169f
C365 B.n325 VSUBS 0.009169f
C366 B.n326 VSUBS 0.022503f
C367 B.n327 VSUBS 0.022503f
C368 B.n328 VSUBS 0.02334f
C369 B.n329 VSUBS 0.009169f
C370 B.n330 VSUBS 0.009169f
C371 B.n331 VSUBS 0.009169f
C372 B.n332 VSUBS 0.009169f
C373 B.n333 VSUBS 0.009169f
C374 B.n334 VSUBS 0.009169f
C375 B.n335 VSUBS 0.009169f
C376 B.n336 VSUBS 0.009169f
C377 B.n337 VSUBS 0.009169f
C378 B.n338 VSUBS 0.009169f
C379 B.n339 VSUBS 0.009169f
C380 B.n340 VSUBS 0.009169f
C381 B.n341 VSUBS 0.009169f
C382 B.n342 VSUBS 0.009169f
C383 B.n343 VSUBS 0.009169f
C384 B.n344 VSUBS 0.009169f
C385 B.n345 VSUBS 0.009169f
C386 B.n346 VSUBS 0.009169f
C387 B.n347 VSUBS 0.009169f
C388 B.n348 VSUBS 0.009169f
C389 B.n349 VSUBS 0.009169f
C390 B.n350 VSUBS 0.009169f
C391 B.n351 VSUBS 0.009169f
C392 B.n352 VSUBS 0.009169f
C393 B.n353 VSUBS 0.009169f
C394 B.n354 VSUBS 0.009169f
C395 B.n355 VSUBS 0.009169f
C396 B.n356 VSUBS 0.009169f
C397 B.n357 VSUBS 0.009169f
C398 B.n358 VSUBS 0.009169f
C399 B.n359 VSUBS 0.009169f
C400 B.n360 VSUBS 0.009169f
C401 B.n361 VSUBS 0.009169f
C402 B.n362 VSUBS 0.009169f
C403 B.n363 VSUBS 0.009169f
C404 B.n364 VSUBS 0.009169f
C405 B.n365 VSUBS 0.009169f
C406 B.n366 VSUBS 0.009169f
C407 B.n367 VSUBS 0.009169f
C408 B.n368 VSUBS 0.009169f
C409 B.n369 VSUBS 0.009169f
C410 B.n370 VSUBS 0.009169f
C411 B.n371 VSUBS 0.009169f
C412 B.n372 VSUBS 0.006337f
C413 B.n373 VSUBS 0.021243f
C414 B.n374 VSUBS 0.007416f
C415 B.n375 VSUBS 0.009169f
C416 B.n376 VSUBS 0.009169f
C417 B.n377 VSUBS 0.009169f
C418 B.n378 VSUBS 0.009169f
C419 B.n379 VSUBS 0.009169f
C420 B.n380 VSUBS 0.009169f
C421 B.n381 VSUBS 0.009169f
C422 B.n382 VSUBS 0.009169f
C423 B.n383 VSUBS 0.009169f
C424 B.n384 VSUBS 0.009169f
C425 B.n385 VSUBS 0.009169f
C426 B.n386 VSUBS 0.007416f
C427 B.n387 VSUBS 0.021243f
C428 B.n388 VSUBS 0.006337f
C429 B.n389 VSUBS 0.009169f
C430 B.n390 VSUBS 0.009169f
C431 B.n391 VSUBS 0.009169f
C432 B.n392 VSUBS 0.009169f
C433 B.n393 VSUBS 0.009169f
C434 B.n394 VSUBS 0.009169f
C435 B.n395 VSUBS 0.009169f
C436 B.n396 VSUBS 0.009169f
C437 B.n397 VSUBS 0.009169f
C438 B.n398 VSUBS 0.009169f
C439 B.n399 VSUBS 0.009169f
C440 B.n400 VSUBS 0.009169f
C441 B.n401 VSUBS 0.009169f
C442 B.n402 VSUBS 0.009169f
C443 B.n403 VSUBS 0.009169f
C444 B.n404 VSUBS 0.009169f
C445 B.n405 VSUBS 0.009169f
C446 B.n406 VSUBS 0.009169f
C447 B.n407 VSUBS 0.009169f
C448 B.n408 VSUBS 0.009169f
C449 B.n409 VSUBS 0.009169f
C450 B.n410 VSUBS 0.009169f
C451 B.n411 VSUBS 0.009169f
C452 B.n412 VSUBS 0.009169f
C453 B.n413 VSUBS 0.009169f
C454 B.n414 VSUBS 0.009169f
C455 B.n415 VSUBS 0.009169f
C456 B.n416 VSUBS 0.009169f
C457 B.n417 VSUBS 0.009169f
C458 B.n418 VSUBS 0.009169f
C459 B.n419 VSUBS 0.009169f
C460 B.n420 VSUBS 0.009169f
C461 B.n421 VSUBS 0.009169f
C462 B.n422 VSUBS 0.009169f
C463 B.n423 VSUBS 0.009169f
C464 B.n424 VSUBS 0.009169f
C465 B.n425 VSUBS 0.009169f
C466 B.n426 VSUBS 0.009169f
C467 B.n427 VSUBS 0.009169f
C468 B.n428 VSUBS 0.009169f
C469 B.n429 VSUBS 0.009169f
C470 B.n430 VSUBS 0.009169f
C471 B.n431 VSUBS 0.009169f
C472 B.n432 VSUBS 0.02334f
C473 B.n433 VSUBS 0.022503f
C474 B.n434 VSUBS 0.023484f
C475 B.n435 VSUBS 0.009169f
C476 B.n436 VSUBS 0.009169f
C477 B.n437 VSUBS 0.009169f
C478 B.n438 VSUBS 0.009169f
C479 B.n439 VSUBS 0.009169f
C480 B.n440 VSUBS 0.009169f
C481 B.n441 VSUBS 0.009169f
C482 B.n442 VSUBS 0.009169f
C483 B.n443 VSUBS 0.009169f
C484 B.n444 VSUBS 0.009169f
C485 B.n445 VSUBS 0.009169f
C486 B.n446 VSUBS 0.009169f
C487 B.n447 VSUBS 0.009169f
C488 B.n448 VSUBS 0.009169f
C489 B.n449 VSUBS 0.009169f
C490 B.n450 VSUBS 0.009169f
C491 B.n451 VSUBS 0.009169f
C492 B.n452 VSUBS 0.009169f
C493 B.n453 VSUBS 0.009169f
C494 B.n454 VSUBS 0.009169f
C495 B.n455 VSUBS 0.009169f
C496 B.n456 VSUBS 0.009169f
C497 B.n457 VSUBS 0.009169f
C498 B.n458 VSUBS 0.009169f
C499 B.n459 VSUBS 0.009169f
C500 B.n460 VSUBS 0.009169f
C501 B.n461 VSUBS 0.009169f
C502 B.n462 VSUBS 0.009169f
C503 B.n463 VSUBS 0.009169f
C504 B.n464 VSUBS 0.009169f
C505 B.n465 VSUBS 0.009169f
C506 B.n466 VSUBS 0.009169f
C507 B.n467 VSUBS 0.009169f
C508 B.n468 VSUBS 0.009169f
C509 B.n469 VSUBS 0.009169f
C510 B.n470 VSUBS 0.009169f
C511 B.n471 VSUBS 0.009169f
C512 B.n472 VSUBS 0.009169f
C513 B.n473 VSUBS 0.009169f
C514 B.n474 VSUBS 0.009169f
C515 B.n475 VSUBS 0.009169f
C516 B.n476 VSUBS 0.009169f
C517 B.n477 VSUBS 0.009169f
C518 B.n478 VSUBS 0.009169f
C519 B.n479 VSUBS 0.009169f
C520 B.n480 VSUBS 0.009169f
C521 B.n481 VSUBS 0.009169f
C522 B.n482 VSUBS 0.009169f
C523 B.n483 VSUBS 0.009169f
C524 B.n484 VSUBS 0.009169f
C525 B.n485 VSUBS 0.009169f
C526 B.n486 VSUBS 0.009169f
C527 B.n487 VSUBS 0.009169f
C528 B.n488 VSUBS 0.009169f
C529 B.n489 VSUBS 0.009169f
C530 B.n490 VSUBS 0.009169f
C531 B.n491 VSUBS 0.009169f
C532 B.n492 VSUBS 0.009169f
C533 B.n493 VSUBS 0.009169f
C534 B.n494 VSUBS 0.009169f
C535 B.n495 VSUBS 0.009169f
C536 B.n496 VSUBS 0.009169f
C537 B.n497 VSUBS 0.009169f
C538 B.n498 VSUBS 0.009169f
C539 B.n499 VSUBS 0.009169f
C540 B.n500 VSUBS 0.009169f
C541 B.n501 VSUBS 0.009169f
C542 B.n502 VSUBS 0.009169f
C543 B.n503 VSUBS 0.009169f
C544 B.n504 VSUBS 0.009169f
C545 B.n505 VSUBS 0.009169f
C546 B.n506 VSUBS 0.009169f
C547 B.n507 VSUBS 0.009169f
C548 B.n508 VSUBS 0.009169f
C549 B.n509 VSUBS 0.009169f
C550 B.n510 VSUBS 0.009169f
C551 B.n511 VSUBS 0.009169f
C552 B.n512 VSUBS 0.009169f
C553 B.n513 VSUBS 0.009169f
C554 B.n514 VSUBS 0.009169f
C555 B.n515 VSUBS 0.009169f
C556 B.n516 VSUBS 0.009169f
C557 B.n517 VSUBS 0.009169f
C558 B.n518 VSUBS 0.009169f
C559 B.n519 VSUBS 0.009169f
C560 B.n520 VSUBS 0.009169f
C561 B.n521 VSUBS 0.009169f
C562 B.n522 VSUBS 0.009169f
C563 B.n523 VSUBS 0.009169f
C564 B.n524 VSUBS 0.009169f
C565 B.n525 VSUBS 0.009169f
C566 B.n526 VSUBS 0.009169f
C567 B.n527 VSUBS 0.009169f
C568 B.n528 VSUBS 0.009169f
C569 B.n529 VSUBS 0.009169f
C570 B.n530 VSUBS 0.009169f
C571 B.n531 VSUBS 0.009169f
C572 B.n532 VSUBS 0.009169f
C573 B.n533 VSUBS 0.009169f
C574 B.n534 VSUBS 0.009169f
C575 B.n535 VSUBS 0.009169f
C576 B.n536 VSUBS 0.009169f
C577 B.n537 VSUBS 0.009169f
C578 B.n538 VSUBS 0.009169f
C579 B.n539 VSUBS 0.009169f
C580 B.n540 VSUBS 0.009169f
C581 B.n541 VSUBS 0.009169f
C582 B.n542 VSUBS 0.009169f
C583 B.n543 VSUBS 0.009169f
C584 B.n544 VSUBS 0.009169f
C585 B.n545 VSUBS 0.009169f
C586 B.n546 VSUBS 0.009169f
C587 B.n547 VSUBS 0.009169f
C588 B.n548 VSUBS 0.009169f
C589 B.n549 VSUBS 0.009169f
C590 B.n550 VSUBS 0.009169f
C591 B.n551 VSUBS 0.009169f
C592 B.n552 VSUBS 0.009169f
C593 B.n553 VSUBS 0.009169f
C594 B.n554 VSUBS 0.009169f
C595 B.n555 VSUBS 0.009169f
C596 B.n556 VSUBS 0.009169f
C597 B.n557 VSUBS 0.009169f
C598 B.n558 VSUBS 0.009169f
C599 B.n559 VSUBS 0.009169f
C600 B.n560 VSUBS 0.009169f
C601 B.n561 VSUBS 0.009169f
C602 B.n562 VSUBS 0.009169f
C603 B.n563 VSUBS 0.009169f
C604 B.n564 VSUBS 0.009169f
C605 B.n565 VSUBS 0.009169f
C606 B.n566 VSUBS 0.009169f
C607 B.n567 VSUBS 0.009169f
C608 B.n568 VSUBS 0.009169f
C609 B.n569 VSUBS 0.009169f
C610 B.n570 VSUBS 0.009169f
C611 B.n571 VSUBS 0.009169f
C612 B.n572 VSUBS 0.009169f
C613 B.n573 VSUBS 0.009169f
C614 B.n574 VSUBS 0.009169f
C615 B.n575 VSUBS 0.009169f
C616 B.n576 VSUBS 0.009169f
C617 B.n577 VSUBS 0.009169f
C618 B.n578 VSUBS 0.009169f
C619 B.n579 VSUBS 0.009169f
C620 B.n580 VSUBS 0.009169f
C621 B.n581 VSUBS 0.009169f
C622 B.n582 VSUBS 0.009169f
C623 B.n583 VSUBS 0.009169f
C624 B.n584 VSUBS 0.009169f
C625 B.n585 VSUBS 0.009169f
C626 B.n586 VSUBS 0.009169f
C627 B.n587 VSUBS 0.009169f
C628 B.n588 VSUBS 0.009169f
C629 B.n589 VSUBS 0.009169f
C630 B.n590 VSUBS 0.009169f
C631 B.n591 VSUBS 0.009169f
C632 B.n592 VSUBS 0.009169f
C633 B.n593 VSUBS 0.009169f
C634 B.n594 VSUBS 0.009169f
C635 B.n595 VSUBS 0.009169f
C636 B.n596 VSUBS 0.009169f
C637 B.n597 VSUBS 0.009169f
C638 B.n598 VSUBS 0.009169f
C639 B.n599 VSUBS 0.009169f
C640 B.n600 VSUBS 0.009169f
C641 B.n601 VSUBS 0.009169f
C642 B.n602 VSUBS 0.009169f
C643 B.n603 VSUBS 0.009169f
C644 B.n604 VSUBS 0.009169f
C645 B.n605 VSUBS 0.009169f
C646 B.n606 VSUBS 0.009169f
C647 B.n607 VSUBS 0.009169f
C648 B.n608 VSUBS 0.009169f
C649 B.n609 VSUBS 0.009169f
C650 B.n610 VSUBS 0.009169f
C651 B.n611 VSUBS 0.009169f
C652 B.n612 VSUBS 0.009169f
C653 B.n613 VSUBS 0.009169f
C654 B.n614 VSUBS 0.009169f
C655 B.n615 VSUBS 0.009169f
C656 B.n616 VSUBS 0.009169f
C657 B.n617 VSUBS 0.009169f
C658 B.n618 VSUBS 0.009169f
C659 B.n619 VSUBS 0.009169f
C660 B.n620 VSUBS 0.009169f
C661 B.n621 VSUBS 0.009169f
C662 B.n622 VSUBS 0.009169f
C663 B.n623 VSUBS 0.009169f
C664 B.n624 VSUBS 0.009169f
C665 B.n625 VSUBS 0.009169f
C666 B.n626 VSUBS 0.009169f
C667 B.n627 VSUBS 0.009169f
C668 B.n628 VSUBS 0.009169f
C669 B.n629 VSUBS 0.009169f
C670 B.n630 VSUBS 0.009169f
C671 B.n631 VSUBS 0.009169f
C672 B.n632 VSUBS 0.009169f
C673 B.n633 VSUBS 0.009169f
C674 B.n634 VSUBS 0.009169f
C675 B.n635 VSUBS 0.009169f
C676 B.n636 VSUBS 0.009169f
C677 B.n637 VSUBS 0.009169f
C678 B.n638 VSUBS 0.009169f
C679 B.n639 VSUBS 0.009169f
C680 B.n640 VSUBS 0.009169f
C681 B.n641 VSUBS 0.009169f
C682 B.n642 VSUBS 0.009169f
C683 B.n643 VSUBS 0.009169f
C684 B.n644 VSUBS 0.009169f
C685 B.n645 VSUBS 0.009169f
C686 B.n646 VSUBS 0.009169f
C687 B.n647 VSUBS 0.009169f
C688 B.n648 VSUBS 0.022503f
C689 B.n649 VSUBS 0.02334f
C690 B.n650 VSUBS 0.02334f
C691 B.n651 VSUBS 0.009169f
C692 B.n652 VSUBS 0.009169f
C693 B.n653 VSUBS 0.009169f
C694 B.n654 VSUBS 0.009169f
C695 B.n655 VSUBS 0.009169f
C696 B.n656 VSUBS 0.009169f
C697 B.n657 VSUBS 0.009169f
C698 B.n658 VSUBS 0.009169f
C699 B.n659 VSUBS 0.009169f
C700 B.n660 VSUBS 0.009169f
C701 B.n661 VSUBS 0.009169f
C702 B.n662 VSUBS 0.009169f
C703 B.n663 VSUBS 0.009169f
C704 B.n664 VSUBS 0.009169f
C705 B.n665 VSUBS 0.009169f
C706 B.n666 VSUBS 0.009169f
C707 B.n667 VSUBS 0.009169f
C708 B.n668 VSUBS 0.009169f
C709 B.n669 VSUBS 0.009169f
C710 B.n670 VSUBS 0.009169f
C711 B.n671 VSUBS 0.009169f
C712 B.n672 VSUBS 0.009169f
C713 B.n673 VSUBS 0.009169f
C714 B.n674 VSUBS 0.009169f
C715 B.n675 VSUBS 0.009169f
C716 B.n676 VSUBS 0.009169f
C717 B.n677 VSUBS 0.009169f
C718 B.n678 VSUBS 0.009169f
C719 B.n679 VSUBS 0.009169f
C720 B.n680 VSUBS 0.009169f
C721 B.n681 VSUBS 0.009169f
C722 B.n682 VSUBS 0.009169f
C723 B.n683 VSUBS 0.009169f
C724 B.n684 VSUBS 0.009169f
C725 B.n685 VSUBS 0.009169f
C726 B.n686 VSUBS 0.009169f
C727 B.n687 VSUBS 0.009169f
C728 B.n688 VSUBS 0.009169f
C729 B.n689 VSUBS 0.009169f
C730 B.n690 VSUBS 0.009169f
C731 B.n691 VSUBS 0.009169f
C732 B.n692 VSUBS 0.009169f
C733 B.n693 VSUBS 0.006337f
C734 B.n694 VSUBS 0.021243f
C735 B.n695 VSUBS 0.007416f
C736 B.n696 VSUBS 0.009169f
C737 B.n697 VSUBS 0.009169f
C738 B.n698 VSUBS 0.009169f
C739 B.n699 VSUBS 0.009169f
C740 B.n700 VSUBS 0.009169f
C741 B.n701 VSUBS 0.009169f
C742 B.n702 VSUBS 0.009169f
C743 B.n703 VSUBS 0.009169f
C744 B.n704 VSUBS 0.009169f
C745 B.n705 VSUBS 0.009169f
C746 B.n706 VSUBS 0.009169f
C747 B.n707 VSUBS 0.007416f
C748 B.n708 VSUBS 0.009169f
C749 B.n709 VSUBS 0.009169f
C750 B.n710 VSUBS 0.009169f
C751 B.n711 VSUBS 0.009169f
C752 B.n712 VSUBS 0.009169f
C753 B.n713 VSUBS 0.009169f
C754 B.n714 VSUBS 0.009169f
C755 B.n715 VSUBS 0.009169f
C756 B.n716 VSUBS 0.009169f
C757 B.n717 VSUBS 0.009169f
C758 B.n718 VSUBS 0.009169f
C759 B.n719 VSUBS 0.009169f
C760 B.n720 VSUBS 0.009169f
C761 B.n721 VSUBS 0.009169f
C762 B.n722 VSUBS 0.009169f
C763 B.n723 VSUBS 0.009169f
C764 B.n724 VSUBS 0.009169f
C765 B.n725 VSUBS 0.009169f
C766 B.n726 VSUBS 0.009169f
C767 B.n727 VSUBS 0.009169f
C768 B.n728 VSUBS 0.009169f
C769 B.n729 VSUBS 0.009169f
C770 B.n730 VSUBS 0.009169f
C771 B.n731 VSUBS 0.009169f
C772 B.n732 VSUBS 0.009169f
C773 B.n733 VSUBS 0.009169f
C774 B.n734 VSUBS 0.009169f
C775 B.n735 VSUBS 0.009169f
C776 B.n736 VSUBS 0.009169f
C777 B.n737 VSUBS 0.009169f
C778 B.n738 VSUBS 0.009169f
C779 B.n739 VSUBS 0.009169f
C780 B.n740 VSUBS 0.009169f
C781 B.n741 VSUBS 0.009169f
C782 B.n742 VSUBS 0.009169f
C783 B.n743 VSUBS 0.009169f
C784 B.n744 VSUBS 0.009169f
C785 B.n745 VSUBS 0.009169f
C786 B.n746 VSUBS 0.009169f
C787 B.n747 VSUBS 0.009169f
C788 B.n748 VSUBS 0.009169f
C789 B.n749 VSUBS 0.009169f
C790 B.n750 VSUBS 0.009169f
C791 B.n751 VSUBS 0.009169f
C792 B.n752 VSUBS 0.02334f
C793 B.n753 VSUBS 0.02334f
C794 B.n754 VSUBS 0.022503f
C795 B.n755 VSUBS 0.009169f
C796 B.n756 VSUBS 0.009169f
C797 B.n757 VSUBS 0.009169f
C798 B.n758 VSUBS 0.009169f
C799 B.n759 VSUBS 0.009169f
C800 B.n760 VSUBS 0.009169f
C801 B.n761 VSUBS 0.009169f
C802 B.n762 VSUBS 0.009169f
C803 B.n763 VSUBS 0.009169f
C804 B.n764 VSUBS 0.009169f
C805 B.n765 VSUBS 0.009169f
C806 B.n766 VSUBS 0.009169f
C807 B.n767 VSUBS 0.009169f
C808 B.n768 VSUBS 0.009169f
C809 B.n769 VSUBS 0.009169f
C810 B.n770 VSUBS 0.009169f
C811 B.n771 VSUBS 0.009169f
C812 B.n772 VSUBS 0.009169f
C813 B.n773 VSUBS 0.009169f
C814 B.n774 VSUBS 0.009169f
C815 B.n775 VSUBS 0.009169f
C816 B.n776 VSUBS 0.009169f
C817 B.n777 VSUBS 0.009169f
C818 B.n778 VSUBS 0.009169f
C819 B.n779 VSUBS 0.009169f
C820 B.n780 VSUBS 0.009169f
C821 B.n781 VSUBS 0.009169f
C822 B.n782 VSUBS 0.009169f
C823 B.n783 VSUBS 0.009169f
C824 B.n784 VSUBS 0.009169f
C825 B.n785 VSUBS 0.009169f
C826 B.n786 VSUBS 0.009169f
C827 B.n787 VSUBS 0.009169f
C828 B.n788 VSUBS 0.009169f
C829 B.n789 VSUBS 0.009169f
C830 B.n790 VSUBS 0.009169f
C831 B.n791 VSUBS 0.009169f
C832 B.n792 VSUBS 0.009169f
C833 B.n793 VSUBS 0.009169f
C834 B.n794 VSUBS 0.009169f
C835 B.n795 VSUBS 0.009169f
C836 B.n796 VSUBS 0.009169f
C837 B.n797 VSUBS 0.009169f
C838 B.n798 VSUBS 0.009169f
C839 B.n799 VSUBS 0.009169f
C840 B.n800 VSUBS 0.009169f
C841 B.n801 VSUBS 0.009169f
C842 B.n802 VSUBS 0.009169f
C843 B.n803 VSUBS 0.009169f
C844 B.n804 VSUBS 0.009169f
C845 B.n805 VSUBS 0.009169f
C846 B.n806 VSUBS 0.009169f
C847 B.n807 VSUBS 0.009169f
C848 B.n808 VSUBS 0.009169f
C849 B.n809 VSUBS 0.009169f
C850 B.n810 VSUBS 0.009169f
C851 B.n811 VSUBS 0.009169f
C852 B.n812 VSUBS 0.009169f
C853 B.n813 VSUBS 0.009169f
C854 B.n814 VSUBS 0.009169f
C855 B.n815 VSUBS 0.009169f
C856 B.n816 VSUBS 0.009169f
C857 B.n817 VSUBS 0.009169f
C858 B.n818 VSUBS 0.009169f
C859 B.n819 VSUBS 0.009169f
C860 B.n820 VSUBS 0.009169f
C861 B.n821 VSUBS 0.009169f
C862 B.n822 VSUBS 0.009169f
C863 B.n823 VSUBS 0.009169f
C864 B.n824 VSUBS 0.009169f
C865 B.n825 VSUBS 0.009169f
C866 B.n826 VSUBS 0.009169f
C867 B.n827 VSUBS 0.009169f
C868 B.n828 VSUBS 0.009169f
C869 B.n829 VSUBS 0.009169f
C870 B.n830 VSUBS 0.009169f
C871 B.n831 VSUBS 0.009169f
C872 B.n832 VSUBS 0.009169f
C873 B.n833 VSUBS 0.009169f
C874 B.n834 VSUBS 0.009169f
C875 B.n835 VSUBS 0.009169f
C876 B.n836 VSUBS 0.009169f
C877 B.n837 VSUBS 0.009169f
C878 B.n838 VSUBS 0.009169f
C879 B.n839 VSUBS 0.009169f
C880 B.n840 VSUBS 0.009169f
C881 B.n841 VSUBS 0.009169f
C882 B.n842 VSUBS 0.009169f
C883 B.n843 VSUBS 0.009169f
C884 B.n844 VSUBS 0.009169f
C885 B.n845 VSUBS 0.009169f
C886 B.n846 VSUBS 0.009169f
C887 B.n847 VSUBS 0.009169f
C888 B.n848 VSUBS 0.009169f
C889 B.n849 VSUBS 0.009169f
C890 B.n850 VSUBS 0.009169f
C891 B.n851 VSUBS 0.009169f
C892 B.n852 VSUBS 0.009169f
C893 B.n853 VSUBS 0.009169f
C894 B.n854 VSUBS 0.009169f
C895 B.n855 VSUBS 0.009169f
C896 B.n856 VSUBS 0.009169f
C897 B.n857 VSUBS 0.009169f
C898 B.n858 VSUBS 0.009169f
C899 B.n859 VSUBS 0.011965f
C900 B.n860 VSUBS 0.012745f
C901 B.n861 VSUBS 0.025345f
C902 VDD2.t0 VSUBS 0.228683f
C903 VDD2.t2 VSUBS 0.228683f
C904 VDD2.n0 VSUBS 1.68887f
C905 VDD2.t6 VSUBS 0.228683f
C906 VDD2.t1 VSUBS 0.228683f
C907 VDD2.n1 VSUBS 1.68887f
C908 VDD2.n2 VSUBS 6.14653f
C909 VDD2.t7 VSUBS 0.228683f
C910 VDD2.t5 VSUBS 0.228683f
C911 VDD2.n3 VSUBS 1.66308f
C912 VDD2.n4 VSUBS 4.82513f
C913 VDD2.t3 VSUBS 0.228683f
C914 VDD2.t4 VSUBS 0.228683f
C915 VDD2.n5 VSUBS 1.68882f
C916 VN.n0 VSUBS 0.050965f
C917 VN.t6 VSUBS 2.32951f
C918 VN.n1 VSUBS 0.050259f
C919 VN.n2 VSUBS 0.027103f
C920 VN.n3 VSUBS 0.050259f
C921 VN.n4 VSUBS 0.027103f
C922 VN.t1 VSUBS 2.32951f
C923 VN.n5 VSUBS 0.050259f
C924 VN.n6 VSUBS 0.027103f
C925 VN.n7 VSUBS 0.050259f
C926 VN.n8 VSUBS 0.35778f
C927 VN.t5 VSUBS 2.32951f
C928 VN.t7 VSUBS 2.74922f
C929 VN.n9 VSUBS 0.894075f
C930 VN.n10 VSUBS 0.929223f
C931 VN.n11 VSUBS 0.033387f
C932 VN.n12 VSUBS 0.050259f
C933 VN.n13 VSUBS 0.027103f
C934 VN.n14 VSUBS 0.027103f
C935 VN.n15 VSUBS 0.027103f
C936 VN.n16 VSUBS 0.053583f
C937 VN.n17 VSUBS 0.02189f
C938 VN.n18 VSUBS 0.053583f
C939 VN.n19 VSUBS 0.027103f
C940 VN.n20 VSUBS 0.027103f
C941 VN.n21 VSUBS 0.027103f
C942 VN.n22 VSUBS 0.050259f
C943 VN.n23 VSUBS 0.033387f
C944 VN.n24 VSUBS 0.834987f
C945 VN.n25 VSUBS 0.04232f
C946 VN.n26 VSUBS 0.027103f
C947 VN.n27 VSUBS 0.027103f
C948 VN.n28 VSUBS 0.027103f
C949 VN.n29 VSUBS 0.050259f
C950 VN.n30 VSUBS 0.044647f
C951 VN.n31 VSUBS 0.034149f
C952 VN.n32 VSUBS 0.027103f
C953 VN.n33 VSUBS 0.027103f
C954 VN.n34 VSUBS 0.027103f
C955 VN.n35 VSUBS 0.050259f
C956 VN.n36 VSUBS 0.049267f
C957 VN.n37 VSUBS 0.959982f
C958 VN.n38 VSUBS 0.08133f
C959 VN.n39 VSUBS 0.050965f
C960 VN.t0 VSUBS 2.32951f
C961 VN.n40 VSUBS 0.050259f
C962 VN.n41 VSUBS 0.027103f
C963 VN.n42 VSUBS 0.050259f
C964 VN.n43 VSUBS 0.027103f
C965 VN.t2 VSUBS 2.32951f
C966 VN.n44 VSUBS 0.050259f
C967 VN.n45 VSUBS 0.027103f
C968 VN.n46 VSUBS 0.050259f
C969 VN.n47 VSUBS 0.35778f
C970 VN.t4 VSUBS 2.32951f
C971 VN.t3 VSUBS 2.74922f
C972 VN.n48 VSUBS 0.894075f
C973 VN.n49 VSUBS 0.929223f
C974 VN.n50 VSUBS 0.033387f
C975 VN.n51 VSUBS 0.050259f
C976 VN.n52 VSUBS 0.027103f
C977 VN.n53 VSUBS 0.027103f
C978 VN.n54 VSUBS 0.027103f
C979 VN.n55 VSUBS 0.053583f
C980 VN.n56 VSUBS 0.02189f
C981 VN.n57 VSUBS 0.053583f
C982 VN.n58 VSUBS 0.027103f
C983 VN.n59 VSUBS 0.027103f
C984 VN.n60 VSUBS 0.027103f
C985 VN.n61 VSUBS 0.050259f
C986 VN.n62 VSUBS 0.033387f
C987 VN.n63 VSUBS 0.834987f
C988 VN.n64 VSUBS 0.04232f
C989 VN.n65 VSUBS 0.027103f
C990 VN.n66 VSUBS 0.027103f
C991 VN.n67 VSUBS 0.027103f
C992 VN.n68 VSUBS 0.050259f
C993 VN.n69 VSUBS 0.044647f
C994 VN.n70 VSUBS 0.034149f
C995 VN.n71 VSUBS 0.027103f
C996 VN.n72 VSUBS 0.027103f
C997 VN.n73 VSUBS 0.027103f
C998 VN.n74 VSUBS 0.050259f
C999 VN.n75 VSUBS 0.049267f
C1000 VN.n76 VSUBS 0.959982f
C1001 VN.n77 VSUBS 1.78904f
C1002 VTAIL.t3 VSUBS 0.182472f
C1003 VTAIL.t0 VSUBS 0.182472f
C1004 VTAIL.n0 VSUBS 1.21326f
C1005 VTAIL.n1 VSUBS 0.908016f
C1006 VTAIL.n2 VSUBS 0.031271f
C1007 VTAIL.n3 VSUBS 0.028792f
C1008 VTAIL.n4 VSUBS 0.015927f
C1009 VTAIL.n5 VSUBS 0.036569f
C1010 VTAIL.n6 VSUBS 0.016382f
C1011 VTAIL.n7 VSUBS 0.028792f
C1012 VTAIL.n8 VSUBS 0.015472f
C1013 VTAIL.n9 VSUBS 0.036569f
C1014 VTAIL.n10 VSUBS 0.016382f
C1015 VTAIL.n11 VSUBS 0.028792f
C1016 VTAIL.n12 VSUBS 0.015472f
C1017 VTAIL.n13 VSUBS 0.027427f
C1018 VTAIL.n14 VSUBS 0.027509f
C1019 VTAIL.t1 VSUBS 0.078573f
C1020 VTAIL.n15 VSUBS 0.175072f
C1021 VTAIL.n16 VSUBS 0.912244f
C1022 VTAIL.n17 VSUBS 0.015472f
C1023 VTAIL.n18 VSUBS 0.016382f
C1024 VTAIL.n19 VSUBS 0.036569f
C1025 VTAIL.n20 VSUBS 0.036569f
C1026 VTAIL.n21 VSUBS 0.016382f
C1027 VTAIL.n22 VSUBS 0.015472f
C1028 VTAIL.n23 VSUBS 0.028792f
C1029 VTAIL.n24 VSUBS 0.028792f
C1030 VTAIL.n25 VSUBS 0.015472f
C1031 VTAIL.n26 VSUBS 0.016382f
C1032 VTAIL.n27 VSUBS 0.036569f
C1033 VTAIL.n28 VSUBS 0.036569f
C1034 VTAIL.n29 VSUBS 0.016382f
C1035 VTAIL.n30 VSUBS 0.015472f
C1036 VTAIL.n31 VSUBS 0.028792f
C1037 VTAIL.n32 VSUBS 0.028792f
C1038 VTAIL.n33 VSUBS 0.015472f
C1039 VTAIL.n34 VSUBS 0.015472f
C1040 VTAIL.n35 VSUBS 0.016382f
C1041 VTAIL.n36 VSUBS 0.036569f
C1042 VTAIL.n37 VSUBS 0.036569f
C1043 VTAIL.n38 VSUBS 0.087288f
C1044 VTAIL.n39 VSUBS 0.015927f
C1045 VTAIL.n40 VSUBS 0.015472f
C1046 VTAIL.n41 VSUBS 0.075204f
C1047 VTAIL.n42 VSUBS 0.044093f
C1048 VTAIL.n43 VSUBS 0.418577f
C1049 VTAIL.n44 VSUBS 0.031271f
C1050 VTAIL.n45 VSUBS 0.028792f
C1051 VTAIL.n46 VSUBS 0.015927f
C1052 VTAIL.n47 VSUBS 0.036569f
C1053 VTAIL.n48 VSUBS 0.016382f
C1054 VTAIL.n49 VSUBS 0.028792f
C1055 VTAIL.n50 VSUBS 0.015472f
C1056 VTAIL.n51 VSUBS 0.036569f
C1057 VTAIL.n52 VSUBS 0.016382f
C1058 VTAIL.n53 VSUBS 0.028792f
C1059 VTAIL.n54 VSUBS 0.015472f
C1060 VTAIL.n55 VSUBS 0.027427f
C1061 VTAIL.n56 VSUBS 0.027509f
C1062 VTAIL.t12 VSUBS 0.078573f
C1063 VTAIL.n57 VSUBS 0.175072f
C1064 VTAIL.n58 VSUBS 0.912244f
C1065 VTAIL.n59 VSUBS 0.015472f
C1066 VTAIL.n60 VSUBS 0.016382f
C1067 VTAIL.n61 VSUBS 0.036569f
C1068 VTAIL.n62 VSUBS 0.036569f
C1069 VTAIL.n63 VSUBS 0.016382f
C1070 VTAIL.n64 VSUBS 0.015472f
C1071 VTAIL.n65 VSUBS 0.028792f
C1072 VTAIL.n66 VSUBS 0.028792f
C1073 VTAIL.n67 VSUBS 0.015472f
C1074 VTAIL.n68 VSUBS 0.016382f
C1075 VTAIL.n69 VSUBS 0.036569f
C1076 VTAIL.n70 VSUBS 0.036569f
C1077 VTAIL.n71 VSUBS 0.016382f
C1078 VTAIL.n72 VSUBS 0.015472f
C1079 VTAIL.n73 VSUBS 0.028792f
C1080 VTAIL.n74 VSUBS 0.028792f
C1081 VTAIL.n75 VSUBS 0.015472f
C1082 VTAIL.n76 VSUBS 0.015472f
C1083 VTAIL.n77 VSUBS 0.016382f
C1084 VTAIL.n78 VSUBS 0.036569f
C1085 VTAIL.n79 VSUBS 0.036569f
C1086 VTAIL.n80 VSUBS 0.087288f
C1087 VTAIL.n81 VSUBS 0.015927f
C1088 VTAIL.n82 VSUBS 0.015472f
C1089 VTAIL.n83 VSUBS 0.075204f
C1090 VTAIL.n84 VSUBS 0.044093f
C1091 VTAIL.n85 VSUBS 0.418577f
C1092 VTAIL.t9 VSUBS 0.182472f
C1093 VTAIL.t14 VSUBS 0.182472f
C1094 VTAIL.n86 VSUBS 1.21326f
C1095 VTAIL.n87 VSUBS 1.24812f
C1096 VTAIL.n88 VSUBS 0.031271f
C1097 VTAIL.n89 VSUBS 0.028792f
C1098 VTAIL.n90 VSUBS 0.015927f
C1099 VTAIL.n91 VSUBS 0.036569f
C1100 VTAIL.n92 VSUBS 0.016382f
C1101 VTAIL.n93 VSUBS 0.028792f
C1102 VTAIL.n94 VSUBS 0.015472f
C1103 VTAIL.n95 VSUBS 0.036569f
C1104 VTAIL.n96 VSUBS 0.016382f
C1105 VTAIL.n97 VSUBS 0.028792f
C1106 VTAIL.n98 VSUBS 0.015472f
C1107 VTAIL.n99 VSUBS 0.027427f
C1108 VTAIL.n100 VSUBS 0.027509f
C1109 VTAIL.t11 VSUBS 0.078573f
C1110 VTAIL.n101 VSUBS 0.175072f
C1111 VTAIL.n102 VSUBS 0.912244f
C1112 VTAIL.n103 VSUBS 0.015472f
C1113 VTAIL.n104 VSUBS 0.016382f
C1114 VTAIL.n105 VSUBS 0.036569f
C1115 VTAIL.n106 VSUBS 0.036569f
C1116 VTAIL.n107 VSUBS 0.016382f
C1117 VTAIL.n108 VSUBS 0.015472f
C1118 VTAIL.n109 VSUBS 0.028792f
C1119 VTAIL.n110 VSUBS 0.028792f
C1120 VTAIL.n111 VSUBS 0.015472f
C1121 VTAIL.n112 VSUBS 0.016382f
C1122 VTAIL.n113 VSUBS 0.036569f
C1123 VTAIL.n114 VSUBS 0.036569f
C1124 VTAIL.n115 VSUBS 0.016382f
C1125 VTAIL.n116 VSUBS 0.015472f
C1126 VTAIL.n117 VSUBS 0.028792f
C1127 VTAIL.n118 VSUBS 0.028792f
C1128 VTAIL.n119 VSUBS 0.015472f
C1129 VTAIL.n120 VSUBS 0.015472f
C1130 VTAIL.n121 VSUBS 0.016382f
C1131 VTAIL.n122 VSUBS 0.036569f
C1132 VTAIL.n123 VSUBS 0.036569f
C1133 VTAIL.n124 VSUBS 0.087288f
C1134 VTAIL.n125 VSUBS 0.015927f
C1135 VTAIL.n126 VSUBS 0.015472f
C1136 VTAIL.n127 VSUBS 0.075204f
C1137 VTAIL.n128 VSUBS 0.044093f
C1138 VTAIL.n129 VSUBS 1.75301f
C1139 VTAIL.n130 VSUBS 0.031271f
C1140 VTAIL.n131 VSUBS 0.028792f
C1141 VTAIL.n132 VSUBS 0.015927f
C1142 VTAIL.n133 VSUBS 0.036569f
C1143 VTAIL.n134 VSUBS 0.015472f
C1144 VTAIL.n135 VSUBS 0.016382f
C1145 VTAIL.n136 VSUBS 0.028792f
C1146 VTAIL.n137 VSUBS 0.015472f
C1147 VTAIL.n138 VSUBS 0.036569f
C1148 VTAIL.n139 VSUBS 0.016382f
C1149 VTAIL.n140 VSUBS 0.028792f
C1150 VTAIL.n141 VSUBS 0.015472f
C1151 VTAIL.n142 VSUBS 0.027427f
C1152 VTAIL.n143 VSUBS 0.027509f
C1153 VTAIL.t6 VSUBS 0.078573f
C1154 VTAIL.n144 VSUBS 0.175072f
C1155 VTAIL.n145 VSUBS 0.912244f
C1156 VTAIL.n146 VSUBS 0.015472f
C1157 VTAIL.n147 VSUBS 0.016382f
C1158 VTAIL.n148 VSUBS 0.036569f
C1159 VTAIL.n149 VSUBS 0.036569f
C1160 VTAIL.n150 VSUBS 0.016382f
C1161 VTAIL.n151 VSUBS 0.015472f
C1162 VTAIL.n152 VSUBS 0.028792f
C1163 VTAIL.n153 VSUBS 0.028792f
C1164 VTAIL.n154 VSUBS 0.015472f
C1165 VTAIL.n155 VSUBS 0.016382f
C1166 VTAIL.n156 VSUBS 0.036569f
C1167 VTAIL.n157 VSUBS 0.036569f
C1168 VTAIL.n158 VSUBS 0.016382f
C1169 VTAIL.n159 VSUBS 0.015472f
C1170 VTAIL.n160 VSUBS 0.028792f
C1171 VTAIL.n161 VSUBS 0.028792f
C1172 VTAIL.n162 VSUBS 0.015472f
C1173 VTAIL.n163 VSUBS 0.016382f
C1174 VTAIL.n164 VSUBS 0.036569f
C1175 VTAIL.n165 VSUBS 0.036569f
C1176 VTAIL.n166 VSUBS 0.087288f
C1177 VTAIL.n167 VSUBS 0.015927f
C1178 VTAIL.n168 VSUBS 0.015472f
C1179 VTAIL.n169 VSUBS 0.075204f
C1180 VTAIL.n170 VSUBS 0.044093f
C1181 VTAIL.n171 VSUBS 1.75301f
C1182 VTAIL.t5 VSUBS 0.182472f
C1183 VTAIL.t4 VSUBS 0.182472f
C1184 VTAIL.n172 VSUBS 1.21327f
C1185 VTAIL.n173 VSUBS 1.24811f
C1186 VTAIL.n174 VSUBS 0.031271f
C1187 VTAIL.n175 VSUBS 0.028792f
C1188 VTAIL.n176 VSUBS 0.015927f
C1189 VTAIL.n177 VSUBS 0.036569f
C1190 VTAIL.n178 VSUBS 0.015472f
C1191 VTAIL.n179 VSUBS 0.016382f
C1192 VTAIL.n180 VSUBS 0.028792f
C1193 VTAIL.n181 VSUBS 0.015472f
C1194 VTAIL.n182 VSUBS 0.036569f
C1195 VTAIL.n183 VSUBS 0.016382f
C1196 VTAIL.n184 VSUBS 0.028792f
C1197 VTAIL.n185 VSUBS 0.015472f
C1198 VTAIL.n186 VSUBS 0.027427f
C1199 VTAIL.n187 VSUBS 0.027509f
C1200 VTAIL.t7 VSUBS 0.078573f
C1201 VTAIL.n188 VSUBS 0.175072f
C1202 VTAIL.n189 VSUBS 0.912244f
C1203 VTAIL.n190 VSUBS 0.015472f
C1204 VTAIL.n191 VSUBS 0.016382f
C1205 VTAIL.n192 VSUBS 0.036569f
C1206 VTAIL.n193 VSUBS 0.036569f
C1207 VTAIL.n194 VSUBS 0.016382f
C1208 VTAIL.n195 VSUBS 0.015472f
C1209 VTAIL.n196 VSUBS 0.028792f
C1210 VTAIL.n197 VSUBS 0.028792f
C1211 VTAIL.n198 VSUBS 0.015472f
C1212 VTAIL.n199 VSUBS 0.016382f
C1213 VTAIL.n200 VSUBS 0.036569f
C1214 VTAIL.n201 VSUBS 0.036569f
C1215 VTAIL.n202 VSUBS 0.016382f
C1216 VTAIL.n203 VSUBS 0.015472f
C1217 VTAIL.n204 VSUBS 0.028792f
C1218 VTAIL.n205 VSUBS 0.028792f
C1219 VTAIL.n206 VSUBS 0.015472f
C1220 VTAIL.n207 VSUBS 0.016382f
C1221 VTAIL.n208 VSUBS 0.036569f
C1222 VTAIL.n209 VSUBS 0.036569f
C1223 VTAIL.n210 VSUBS 0.087288f
C1224 VTAIL.n211 VSUBS 0.015927f
C1225 VTAIL.n212 VSUBS 0.015472f
C1226 VTAIL.n213 VSUBS 0.075204f
C1227 VTAIL.n214 VSUBS 0.044093f
C1228 VTAIL.n215 VSUBS 0.418577f
C1229 VTAIL.n216 VSUBS 0.031271f
C1230 VTAIL.n217 VSUBS 0.028792f
C1231 VTAIL.n218 VSUBS 0.015927f
C1232 VTAIL.n219 VSUBS 0.036569f
C1233 VTAIL.n220 VSUBS 0.015472f
C1234 VTAIL.n221 VSUBS 0.016382f
C1235 VTAIL.n222 VSUBS 0.028792f
C1236 VTAIL.n223 VSUBS 0.015472f
C1237 VTAIL.n224 VSUBS 0.036569f
C1238 VTAIL.n225 VSUBS 0.016382f
C1239 VTAIL.n226 VSUBS 0.028792f
C1240 VTAIL.n227 VSUBS 0.015472f
C1241 VTAIL.n228 VSUBS 0.027427f
C1242 VTAIL.n229 VSUBS 0.027509f
C1243 VTAIL.t10 VSUBS 0.078573f
C1244 VTAIL.n230 VSUBS 0.175072f
C1245 VTAIL.n231 VSUBS 0.912244f
C1246 VTAIL.n232 VSUBS 0.015472f
C1247 VTAIL.n233 VSUBS 0.016382f
C1248 VTAIL.n234 VSUBS 0.036569f
C1249 VTAIL.n235 VSUBS 0.036569f
C1250 VTAIL.n236 VSUBS 0.016382f
C1251 VTAIL.n237 VSUBS 0.015472f
C1252 VTAIL.n238 VSUBS 0.028792f
C1253 VTAIL.n239 VSUBS 0.028792f
C1254 VTAIL.n240 VSUBS 0.015472f
C1255 VTAIL.n241 VSUBS 0.016382f
C1256 VTAIL.n242 VSUBS 0.036569f
C1257 VTAIL.n243 VSUBS 0.036569f
C1258 VTAIL.n244 VSUBS 0.016382f
C1259 VTAIL.n245 VSUBS 0.015472f
C1260 VTAIL.n246 VSUBS 0.028792f
C1261 VTAIL.n247 VSUBS 0.028792f
C1262 VTAIL.n248 VSUBS 0.015472f
C1263 VTAIL.n249 VSUBS 0.016382f
C1264 VTAIL.n250 VSUBS 0.036569f
C1265 VTAIL.n251 VSUBS 0.036569f
C1266 VTAIL.n252 VSUBS 0.087288f
C1267 VTAIL.n253 VSUBS 0.015927f
C1268 VTAIL.n254 VSUBS 0.015472f
C1269 VTAIL.n255 VSUBS 0.075204f
C1270 VTAIL.n256 VSUBS 0.044093f
C1271 VTAIL.n257 VSUBS 0.418577f
C1272 VTAIL.t13 VSUBS 0.182472f
C1273 VTAIL.t15 VSUBS 0.182472f
C1274 VTAIL.n258 VSUBS 1.21327f
C1275 VTAIL.n259 VSUBS 1.24811f
C1276 VTAIL.n260 VSUBS 0.031271f
C1277 VTAIL.n261 VSUBS 0.028792f
C1278 VTAIL.n262 VSUBS 0.015927f
C1279 VTAIL.n263 VSUBS 0.036569f
C1280 VTAIL.n264 VSUBS 0.015472f
C1281 VTAIL.n265 VSUBS 0.016382f
C1282 VTAIL.n266 VSUBS 0.028792f
C1283 VTAIL.n267 VSUBS 0.015472f
C1284 VTAIL.n268 VSUBS 0.036569f
C1285 VTAIL.n269 VSUBS 0.016382f
C1286 VTAIL.n270 VSUBS 0.028792f
C1287 VTAIL.n271 VSUBS 0.015472f
C1288 VTAIL.n272 VSUBS 0.027427f
C1289 VTAIL.n273 VSUBS 0.027509f
C1290 VTAIL.t8 VSUBS 0.078573f
C1291 VTAIL.n274 VSUBS 0.175072f
C1292 VTAIL.n275 VSUBS 0.912244f
C1293 VTAIL.n276 VSUBS 0.015472f
C1294 VTAIL.n277 VSUBS 0.016382f
C1295 VTAIL.n278 VSUBS 0.036569f
C1296 VTAIL.n279 VSUBS 0.036569f
C1297 VTAIL.n280 VSUBS 0.016382f
C1298 VTAIL.n281 VSUBS 0.015472f
C1299 VTAIL.n282 VSUBS 0.028792f
C1300 VTAIL.n283 VSUBS 0.028792f
C1301 VTAIL.n284 VSUBS 0.015472f
C1302 VTAIL.n285 VSUBS 0.016382f
C1303 VTAIL.n286 VSUBS 0.036569f
C1304 VTAIL.n287 VSUBS 0.036569f
C1305 VTAIL.n288 VSUBS 0.016382f
C1306 VTAIL.n289 VSUBS 0.015472f
C1307 VTAIL.n290 VSUBS 0.028792f
C1308 VTAIL.n291 VSUBS 0.028792f
C1309 VTAIL.n292 VSUBS 0.015472f
C1310 VTAIL.n293 VSUBS 0.016382f
C1311 VTAIL.n294 VSUBS 0.036569f
C1312 VTAIL.n295 VSUBS 0.036569f
C1313 VTAIL.n296 VSUBS 0.087288f
C1314 VTAIL.n297 VSUBS 0.015927f
C1315 VTAIL.n298 VSUBS 0.015472f
C1316 VTAIL.n299 VSUBS 0.075204f
C1317 VTAIL.n300 VSUBS 0.044093f
C1318 VTAIL.n301 VSUBS 1.75301f
C1319 VTAIL.n302 VSUBS 0.031271f
C1320 VTAIL.n303 VSUBS 0.028792f
C1321 VTAIL.n304 VSUBS 0.015927f
C1322 VTAIL.n305 VSUBS 0.036569f
C1323 VTAIL.n306 VSUBS 0.016382f
C1324 VTAIL.n307 VSUBS 0.028792f
C1325 VTAIL.n308 VSUBS 0.015472f
C1326 VTAIL.n309 VSUBS 0.036569f
C1327 VTAIL.n310 VSUBS 0.016382f
C1328 VTAIL.n311 VSUBS 0.028792f
C1329 VTAIL.n312 VSUBS 0.015472f
C1330 VTAIL.n313 VSUBS 0.027427f
C1331 VTAIL.n314 VSUBS 0.027509f
C1332 VTAIL.t2 VSUBS 0.078573f
C1333 VTAIL.n315 VSUBS 0.175072f
C1334 VTAIL.n316 VSUBS 0.912244f
C1335 VTAIL.n317 VSUBS 0.015472f
C1336 VTAIL.n318 VSUBS 0.016382f
C1337 VTAIL.n319 VSUBS 0.036569f
C1338 VTAIL.n320 VSUBS 0.036569f
C1339 VTAIL.n321 VSUBS 0.016382f
C1340 VTAIL.n322 VSUBS 0.015472f
C1341 VTAIL.n323 VSUBS 0.028792f
C1342 VTAIL.n324 VSUBS 0.028792f
C1343 VTAIL.n325 VSUBS 0.015472f
C1344 VTAIL.n326 VSUBS 0.016382f
C1345 VTAIL.n327 VSUBS 0.036569f
C1346 VTAIL.n328 VSUBS 0.036569f
C1347 VTAIL.n329 VSUBS 0.016382f
C1348 VTAIL.n330 VSUBS 0.015472f
C1349 VTAIL.n331 VSUBS 0.028792f
C1350 VTAIL.n332 VSUBS 0.028792f
C1351 VTAIL.n333 VSUBS 0.015472f
C1352 VTAIL.n334 VSUBS 0.015472f
C1353 VTAIL.n335 VSUBS 0.016382f
C1354 VTAIL.n336 VSUBS 0.036569f
C1355 VTAIL.n337 VSUBS 0.036569f
C1356 VTAIL.n338 VSUBS 0.087288f
C1357 VTAIL.n339 VSUBS 0.015927f
C1358 VTAIL.n340 VSUBS 0.015472f
C1359 VTAIL.n341 VSUBS 0.075204f
C1360 VTAIL.n342 VSUBS 0.044093f
C1361 VTAIL.n343 VSUBS 1.74761f
C1362 VDD1.t0 VSUBS 0.206888f
C1363 VDD1.t7 VSUBS 0.206888f
C1364 VDD1.n0 VSUBS 1.5296f
C1365 VDD1.t2 VSUBS 0.206888f
C1366 VDD1.t1 VSUBS 0.206888f
C1367 VDD1.n1 VSUBS 1.52791f
C1368 VDD1.t5 VSUBS 0.206888f
C1369 VDD1.t6 VSUBS 0.206888f
C1370 VDD1.n2 VSUBS 1.52791f
C1371 VDD1.n3 VSUBS 5.62792f
C1372 VDD1.t4 VSUBS 0.206888f
C1373 VDD1.t3 VSUBS 0.206888f
C1374 VDD1.n4 VSUBS 1.50457f
C1375 VDD1.n5 VSUBS 4.40637f
C1376 VP.n0 VSUBS 0.057116f
C1377 VP.t3 VSUBS 2.61062f
C1378 VP.n1 VSUBS 0.056325f
C1379 VP.n2 VSUBS 0.030373f
C1380 VP.n3 VSUBS 0.056325f
C1381 VP.n4 VSUBS 0.030373f
C1382 VP.t1 VSUBS 2.61062f
C1383 VP.n5 VSUBS 0.056325f
C1384 VP.n6 VSUBS 0.030373f
C1385 VP.n7 VSUBS 0.056325f
C1386 VP.n8 VSUBS 0.030373f
C1387 VP.t6 VSUBS 2.61062f
C1388 VP.n9 VSUBS 0.056325f
C1389 VP.n10 VSUBS 0.030373f
C1390 VP.n11 VSUBS 0.056325f
C1391 VP.n12 VSUBS 0.057116f
C1392 VP.t4 VSUBS 2.61062f
C1393 VP.n13 VSUBS 0.057116f
C1394 VP.t7 VSUBS 2.61062f
C1395 VP.n14 VSUBS 0.056325f
C1396 VP.n15 VSUBS 0.030373f
C1397 VP.n16 VSUBS 0.056325f
C1398 VP.n17 VSUBS 0.030373f
C1399 VP.t0 VSUBS 2.61062f
C1400 VP.n18 VSUBS 0.056325f
C1401 VP.n19 VSUBS 0.030373f
C1402 VP.n20 VSUBS 0.056325f
C1403 VP.n21 VSUBS 0.400957f
C1404 VP.t2 VSUBS 2.61062f
C1405 VP.t5 VSUBS 3.08099f
C1406 VP.n22 VSUBS 1.00197f
C1407 VP.n23 VSUBS 1.04136f
C1408 VP.n24 VSUBS 0.037416f
C1409 VP.n25 VSUBS 0.056325f
C1410 VP.n26 VSUBS 0.030373f
C1411 VP.n27 VSUBS 0.030373f
C1412 VP.n28 VSUBS 0.030373f
C1413 VP.n29 VSUBS 0.060049f
C1414 VP.n30 VSUBS 0.024532f
C1415 VP.n31 VSUBS 0.060049f
C1416 VP.n32 VSUBS 0.030373f
C1417 VP.n33 VSUBS 0.030373f
C1418 VP.n34 VSUBS 0.030373f
C1419 VP.n35 VSUBS 0.056325f
C1420 VP.n36 VSUBS 0.037416f
C1421 VP.n37 VSUBS 0.935751f
C1422 VP.n38 VSUBS 0.047427f
C1423 VP.n39 VSUBS 0.030373f
C1424 VP.n40 VSUBS 0.030373f
C1425 VP.n41 VSUBS 0.030373f
C1426 VP.n42 VSUBS 0.056325f
C1427 VP.n43 VSUBS 0.050035f
C1428 VP.n44 VSUBS 0.03827f
C1429 VP.n45 VSUBS 0.030373f
C1430 VP.n46 VSUBS 0.030373f
C1431 VP.n47 VSUBS 0.030373f
C1432 VP.n48 VSUBS 0.056325f
C1433 VP.n49 VSUBS 0.055212f
C1434 VP.n50 VSUBS 1.07583f
C1435 VP.n51 VSUBS 1.99754f
C1436 VP.n52 VSUBS 2.01756f
C1437 VP.n53 VSUBS 1.07583f
C1438 VP.n54 VSUBS 0.055212f
C1439 VP.n55 VSUBS 0.056325f
C1440 VP.n56 VSUBS 0.030373f
C1441 VP.n57 VSUBS 0.030373f
C1442 VP.n58 VSUBS 0.030373f
C1443 VP.n59 VSUBS 0.03827f
C1444 VP.n60 VSUBS 0.050035f
C1445 VP.n61 VSUBS 0.056325f
C1446 VP.n62 VSUBS 0.030373f
C1447 VP.n63 VSUBS 0.030373f
C1448 VP.n64 VSUBS 0.030373f
C1449 VP.n65 VSUBS 0.047427f
C1450 VP.n66 VSUBS 0.935751f
C1451 VP.n67 VSUBS 0.037416f
C1452 VP.n68 VSUBS 0.056325f
C1453 VP.n69 VSUBS 0.030373f
C1454 VP.n70 VSUBS 0.030373f
C1455 VP.n71 VSUBS 0.030373f
C1456 VP.n72 VSUBS 0.060049f
C1457 VP.n73 VSUBS 0.024532f
C1458 VP.n74 VSUBS 0.060049f
C1459 VP.n75 VSUBS 0.030373f
C1460 VP.n76 VSUBS 0.030373f
C1461 VP.n77 VSUBS 0.030373f
C1462 VP.n78 VSUBS 0.056325f
C1463 VP.n79 VSUBS 0.037416f
C1464 VP.n80 VSUBS 0.935751f
C1465 VP.n81 VSUBS 0.047427f
C1466 VP.n82 VSUBS 0.030373f
C1467 VP.n83 VSUBS 0.030373f
C1468 VP.n84 VSUBS 0.030373f
C1469 VP.n85 VSUBS 0.056325f
C1470 VP.n86 VSUBS 0.050035f
C1471 VP.n87 VSUBS 0.03827f
C1472 VP.n88 VSUBS 0.030373f
C1473 VP.n89 VSUBS 0.030373f
C1474 VP.n90 VSUBS 0.030373f
C1475 VP.n91 VSUBS 0.056325f
C1476 VP.n92 VSUBS 0.055212f
C1477 VP.n93 VSUBS 1.07583f
C1478 VP.n94 VSUBS 0.091144f
.ends

