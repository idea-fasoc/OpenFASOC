* NGSPICE file created from diff_pair_sample_0857.ext - technology: sky130A

.subckt diff_pair_sample_0857 VTAIL VN VP B VDD2 VDD1
X0 B.t11 B.t9 B.t10 w_n2662_n1594# sky130_fd_pr__pfet_01v8 ad=1.2207 pd=7.04 as=0 ps=0 w=3.13 l=2.49
X1 VDD2.t3 VN.t0 VTAIL.t7 w_n2662_n1594# sky130_fd_pr__pfet_01v8 ad=0.51645 pd=3.46 as=1.2207 ps=7.04 w=3.13 l=2.49
X2 VDD1.t3 VP.t0 VTAIL.t1 w_n2662_n1594# sky130_fd_pr__pfet_01v8 ad=0.51645 pd=3.46 as=1.2207 ps=7.04 w=3.13 l=2.49
X3 VTAIL.t4 VN.t1 VDD2.t2 w_n2662_n1594# sky130_fd_pr__pfet_01v8 ad=1.2207 pd=7.04 as=0.51645 ps=3.46 w=3.13 l=2.49
X4 VTAIL.t5 VN.t2 VDD2.t1 w_n2662_n1594# sky130_fd_pr__pfet_01v8 ad=1.2207 pd=7.04 as=0.51645 ps=3.46 w=3.13 l=2.49
X5 VDD2.t0 VN.t3 VTAIL.t6 w_n2662_n1594# sky130_fd_pr__pfet_01v8 ad=0.51645 pd=3.46 as=1.2207 ps=7.04 w=3.13 l=2.49
X6 VTAIL.t2 VP.t1 VDD1.t2 w_n2662_n1594# sky130_fd_pr__pfet_01v8 ad=1.2207 pd=7.04 as=0.51645 ps=3.46 w=3.13 l=2.49
X7 B.t8 B.t6 B.t7 w_n2662_n1594# sky130_fd_pr__pfet_01v8 ad=1.2207 pd=7.04 as=0 ps=0 w=3.13 l=2.49
X8 B.t5 B.t3 B.t4 w_n2662_n1594# sky130_fd_pr__pfet_01v8 ad=1.2207 pd=7.04 as=0 ps=0 w=3.13 l=2.49
X9 B.t2 B.t0 B.t1 w_n2662_n1594# sky130_fd_pr__pfet_01v8 ad=1.2207 pd=7.04 as=0 ps=0 w=3.13 l=2.49
X10 VDD1.t1 VP.t2 VTAIL.t3 w_n2662_n1594# sky130_fd_pr__pfet_01v8 ad=0.51645 pd=3.46 as=1.2207 ps=7.04 w=3.13 l=2.49
X11 VTAIL.t0 VP.t3 VDD1.t0 w_n2662_n1594# sky130_fd_pr__pfet_01v8 ad=1.2207 pd=7.04 as=0.51645 ps=3.46 w=3.13 l=2.49
R0 B.n331 B.n330 585
R1 B.n332 B.n43 585
R2 B.n334 B.n333 585
R3 B.n335 B.n42 585
R4 B.n337 B.n336 585
R5 B.n338 B.n41 585
R6 B.n340 B.n339 585
R7 B.n341 B.n40 585
R8 B.n343 B.n342 585
R9 B.n344 B.n39 585
R10 B.n346 B.n345 585
R11 B.n347 B.n38 585
R12 B.n349 B.n348 585
R13 B.n350 B.n37 585
R14 B.n352 B.n351 585
R15 B.n353 B.n34 585
R16 B.n356 B.n355 585
R17 B.n357 B.n33 585
R18 B.n359 B.n358 585
R19 B.n360 B.n32 585
R20 B.n362 B.n361 585
R21 B.n363 B.n31 585
R22 B.n365 B.n364 585
R23 B.n366 B.n27 585
R24 B.n368 B.n367 585
R25 B.n369 B.n26 585
R26 B.n371 B.n370 585
R27 B.n372 B.n25 585
R28 B.n374 B.n373 585
R29 B.n375 B.n24 585
R30 B.n377 B.n376 585
R31 B.n378 B.n23 585
R32 B.n380 B.n379 585
R33 B.n381 B.n22 585
R34 B.n383 B.n382 585
R35 B.n384 B.n21 585
R36 B.n386 B.n385 585
R37 B.n387 B.n20 585
R38 B.n389 B.n388 585
R39 B.n390 B.n19 585
R40 B.n392 B.n391 585
R41 B.n329 B.n44 585
R42 B.n328 B.n327 585
R43 B.n326 B.n45 585
R44 B.n325 B.n324 585
R45 B.n323 B.n46 585
R46 B.n322 B.n321 585
R47 B.n320 B.n47 585
R48 B.n319 B.n318 585
R49 B.n317 B.n48 585
R50 B.n316 B.n315 585
R51 B.n314 B.n49 585
R52 B.n313 B.n312 585
R53 B.n311 B.n50 585
R54 B.n310 B.n309 585
R55 B.n308 B.n51 585
R56 B.n307 B.n306 585
R57 B.n305 B.n52 585
R58 B.n304 B.n303 585
R59 B.n302 B.n53 585
R60 B.n301 B.n300 585
R61 B.n299 B.n54 585
R62 B.n298 B.n297 585
R63 B.n296 B.n55 585
R64 B.n295 B.n294 585
R65 B.n293 B.n56 585
R66 B.n292 B.n291 585
R67 B.n290 B.n57 585
R68 B.n289 B.n288 585
R69 B.n287 B.n58 585
R70 B.n286 B.n285 585
R71 B.n284 B.n59 585
R72 B.n283 B.n282 585
R73 B.n281 B.n60 585
R74 B.n280 B.n279 585
R75 B.n278 B.n61 585
R76 B.n277 B.n276 585
R77 B.n275 B.n62 585
R78 B.n274 B.n273 585
R79 B.n272 B.n63 585
R80 B.n271 B.n270 585
R81 B.n269 B.n64 585
R82 B.n268 B.n267 585
R83 B.n266 B.n65 585
R84 B.n265 B.n264 585
R85 B.n263 B.n66 585
R86 B.n262 B.n261 585
R87 B.n260 B.n67 585
R88 B.n259 B.n258 585
R89 B.n257 B.n68 585
R90 B.n256 B.n255 585
R91 B.n254 B.n69 585
R92 B.n253 B.n252 585
R93 B.n251 B.n70 585
R94 B.n250 B.n249 585
R95 B.n248 B.n71 585
R96 B.n247 B.n246 585
R97 B.n245 B.n72 585
R98 B.n244 B.n243 585
R99 B.n242 B.n73 585
R100 B.n241 B.n240 585
R101 B.n239 B.n74 585
R102 B.n238 B.n237 585
R103 B.n236 B.n75 585
R104 B.n235 B.n234 585
R105 B.n233 B.n76 585
R106 B.n232 B.n231 585
R107 B.n230 B.n77 585
R108 B.n165 B.n164 585
R109 B.n166 B.n99 585
R110 B.n168 B.n167 585
R111 B.n169 B.n98 585
R112 B.n171 B.n170 585
R113 B.n172 B.n97 585
R114 B.n174 B.n173 585
R115 B.n175 B.n96 585
R116 B.n177 B.n176 585
R117 B.n178 B.n95 585
R118 B.n180 B.n179 585
R119 B.n181 B.n94 585
R120 B.n183 B.n182 585
R121 B.n184 B.n93 585
R122 B.n186 B.n185 585
R123 B.n187 B.n90 585
R124 B.n190 B.n189 585
R125 B.n191 B.n89 585
R126 B.n193 B.n192 585
R127 B.n194 B.n88 585
R128 B.n196 B.n195 585
R129 B.n197 B.n87 585
R130 B.n199 B.n198 585
R131 B.n200 B.n86 585
R132 B.n205 B.n204 585
R133 B.n206 B.n85 585
R134 B.n208 B.n207 585
R135 B.n209 B.n84 585
R136 B.n211 B.n210 585
R137 B.n212 B.n83 585
R138 B.n214 B.n213 585
R139 B.n215 B.n82 585
R140 B.n217 B.n216 585
R141 B.n218 B.n81 585
R142 B.n220 B.n219 585
R143 B.n221 B.n80 585
R144 B.n223 B.n222 585
R145 B.n224 B.n79 585
R146 B.n226 B.n225 585
R147 B.n227 B.n78 585
R148 B.n229 B.n228 585
R149 B.n163 B.n100 585
R150 B.n162 B.n161 585
R151 B.n160 B.n101 585
R152 B.n159 B.n158 585
R153 B.n157 B.n102 585
R154 B.n156 B.n155 585
R155 B.n154 B.n103 585
R156 B.n153 B.n152 585
R157 B.n151 B.n104 585
R158 B.n150 B.n149 585
R159 B.n148 B.n105 585
R160 B.n147 B.n146 585
R161 B.n145 B.n106 585
R162 B.n144 B.n143 585
R163 B.n142 B.n107 585
R164 B.n141 B.n140 585
R165 B.n139 B.n108 585
R166 B.n138 B.n137 585
R167 B.n136 B.n109 585
R168 B.n135 B.n134 585
R169 B.n133 B.n110 585
R170 B.n132 B.n131 585
R171 B.n130 B.n111 585
R172 B.n129 B.n128 585
R173 B.n127 B.n112 585
R174 B.n126 B.n125 585
R175 B.n124 B.n113 585
R176 B.n123 B.n122 585
R177 B.n121 B.n114 585
R178 B.n120 B.n119 585
R179 B.n118 B.n115 585
R180 B.n117 B.n116 585
R181 B.n2 B.n0 585
R182 B.n441 B.n1 585
R183 B.n440 B.n439 585
R184 B.n438 B.n3 585
R185 B.n437 B.n436 585
R186 B.n435 B.n4 585
R187 B.n434 B.n433 585
R188 B.n432 B.n5 585
R189 B.n431 B.n430 585
R190 B.n429 B.n6 585
R191 B.n428 B.n427 585
R192 B.n426 B.n7 585
R193 B.n425 B.n424 585
R194 B.n423 B.n8 585
R195 B.n422 B.n421 585
R196 B.n420 B.n9 585
R197 B.n419 B.n418 585
R198 B.n417 B.n10 585
R199 B.n416 B.n415 585
R200 B.n414 B.n11 585
R201 B.n413 B.n412 585
R202 B.n411 B.n12 585
R203 B.n410 B.n409 585
R204 B.n408 B.n13 585
R205 B.n407 B.n406 585
R206 B.n405 B.n14 585
R207 B.n404 B.n403 585
R208 B.n402 B.n15 585
R209 B.n401 B.n400 585
R210 B.n399 B.n16 585
R211 B.n398 B.n397 585
R212 B.n396 B.n17 585
R213 B.n395 B.n394 585
R214 B.n393 B.n18 585
R215 B.n443 B.n442 585
R216 B.n165 B.n100 468.476
R217 B.n393 B.n392 468.476
R218 B.n230 B.n229 468.476
R219 B.n331 B.n44 468.476
R220 B.n201 B.t8 278.894
R221 B.n35 B.t10 278.894
R222 B.n91 B.t2 278.894
R223 B.n28 B.t4 278.894
R224 B.n201 B.t6 238.169
R225 B.n91 B.t0 238.169
R226 B.n28 B.t3 238.169
R227 B.n35 B.t9 238.169
R228 B.n202 B.t7 224.203
R229 B.n36 B.t11 224.203
R230 B.n92 B.t1 224.203
R231 B.n29 B.t5 224.203
R232 B.n161 B.n100 163.367
R233 B.n161 B.n160 163.367
R234 B.n160 B.n159 163.367
R235 B.n159 B.n102 163.367
R236 B.n155 B.n102 163.367
R237 B.n155 B.n154 163.367
R238 B.n154 B.n153 163.367
R239 B.n153 B.n104 163.367
R240 B.n149 B.n104 163.367
R241 B.n149 B.n148 163.367
R242 B.n148 B.n147 163.367
R243 B.n147 B.n106 163.367
R244 B.n143 B.n106 163.367
R245 B.n143 B.n142 163.367
R246 B.n142 B.n141 163.367
R247 B.n141 B.n108 163.367
R248 B.n137 B.n108 163.367
R249 B.n137 B.n136 163.367
R250 B.n136 B.n135 163.367
R251 B.n135 B.n110 163.367
R252 B.n131 B.n110 163.367
R253 B.n131 B.n130 163.367
R254 B.n130 B.n129 163.367
R255 B.n129 B.n112 163.367
R256 B.n125 B.n112 163.367
R257 B.n125 B.n124 163.367
R258 B.n124 B.n123 163.367
R259 B.n123 B.n114 163.367
R260 B.n119 B.n114 163.367
R261 B.n119 B.n118 163.367
R262 B.n118 B.n117 163.367
R263 B.n117 B.n2 163.367
R264 B.n442 B.n2 163.367
R265 B.n442 B.n441 163.367
R266 B.n441 B.n440 163.367
R267 B.n440 B.n3 163.367
R268 B.n436 B.n3 163.367
R269 B.n436 B.n435 163.367
R270 B.n435 B.n434 163.367
R271 B.n434 B.n5 163.367
R272 B.n430 B.n5 163.367
R273 B.n430 B.n429 163.367
R274 B.n429 B.n428 163.367
R275 B.n428 B.n7 163.367
R276 B.n424 B.n7 163.367
R277 B.n424 B.n423 163.367
R278 B.n423 B.n422 163.367
R279 B.n422 B.n9 163.367
R280 B.n418 B.n9 163.367
R281 B.n418 B.n417 163.367
R282 B.n417 B.n416 163.367
R283 B.n416 B.n11 163.367
R284 B.n412 B.n11 163.367
R285 B.n412 B.n411 163.367
R286 B.n411 B.n410 163.367
R287 B.n410 B.n13 163.367
R288 B.n406 B.n13 163.367
R289 B.n406 B.n405 163.367
R290 B.n405 B.n404 163.367
R291 B.n404 B.n15 163.367
R292 B.n400 B.n15 163.367
R293 B.n400 B.n399 163.367
R294 B.n399 B.n398 163.367
R295 B.n398 B.n17 163.367
R296 B.n394 B.n17 163.367
R297 B.n394 B.n393 163.367
R298 B.n166 B.n165 163.367
R299 B.n167 B.n166 163.367
R300 B.n167 B.n98 163.367
R301 B.n171 B.n98 163.367
R302 B.n172 B.n171 163.367
R303 B.n173 B.n172 163.367
R304 B.n173 B.n96 163.367
R305 B.n177 B.n96 163.367
R306 B.n178 B.n177 163.367
R307 B.n179 B.n178 163.367
R308 B.n179 B.n94 163.367
R309 B.n183 B.n94 163.367
R310 B.n184 B.n183 163.367
R311 B.n185 B.n184 163.367
R312 B.n185 B.n90 163.367
R313 B.n190 B.n90 163.367
R314 B.n191 B.n190 163.367
R315 B.n192 B.n191 163.367
R316 B.n192 B.n88 163.367
R317 B.n196 B.n88 163.367
R318 B.n197 B.n196 163.367
R319 B.n198 B.n197 163.367
R320 B.n198 B.n86 163.367
R321 B.n205 B.n86 163.367
R322 B.n206 B.n205 163.367
R323 B.n207 B.n206 163.367
R324 B.n207 B.n84 163.367
R325 B.n211 B.n84 163.367
R326 B.n212 B.n211 163.367
R327 B.n213 B.n212 163.367
R328 B.n213 B.n82 163.367
R329 B.n217 B.n82 163.367
R330 B.n218 B.n217 163.367
R331 B.n219 B.n218 163.367
R332 B.n219 B.n80 163.367
R333 B.n223 B.n80 163.367
R334 B.n224 B.n223 163.367
R335 B.n225 B.n224 163.367
R336 B.n225 B.n78 163.367
R337 B.n229 B.n78 163.367
R338 B.n231 B.n230 163.367
R339 B.n231 B.n76 163.367
R340 B.n235 B.n76 163.367
R341 B.n236 B.n235 163.367
R342 B.n237 B.n236 163.367
R343 B.n237 B.n74 163.367
R344 B.n241 B.n74 163.367
R345 B.n242 B.n241 163.367
R346 B.n243 B.n242 163.367
R347 B.n243 B.n72 163.367
R348 B.n247 B.n72 163.367
R349 B.n248 B.n247 163.367
R350 B.n249 B.n248 163.367
R351 B.n249 B.n70 163.367
R352 B.n253 B.n70 163.367
R353 B.n254 B.n253 163.367
R354 B.n255 B.n254 163.367
R355 B.n255 B.n68 163.367
R356 B.n259 B.n68 163.367
R357 B.n260 B.n259 163.367
R358 B.n261 B.n260 163.367
R359 B.n261 B.n66 163.367
R360 B.n265 B.n66 163.367
R361 B.n266 B.n265 163.367
R362 B.n267 B.n266 163.367
R363 B.n267 B.n64 163.367
R364 B.n271 B.n64 163.367
R365 B.n272 B.n271 163.367
R366 B.n273 B.n272 163.367
R367 B.n273 B.n62 163.367
R368 B.n277 B.n62 163.367
R369 B.n278 B.n277 163.367
R370 B.n279 B.n278 163.367
R371 B.n279 B.n60 163.367
R372 B.n283 B.n60 163.367
R373 B.n284 B.n283 163.367
R374 B.n285 B.n284 163.367
R375 B.n285 B.n58 163.367
R376 B.n289 B.n58 163.367
R377 B.n290 B.n289 163.367
R378 B.n291 B.n290 163.367
R379 B.n291 B.n56 163.367
R380 B.n295 B.n56 163.367
R381 B.n296 B.n295 163.367
R382 B.n297 B.n296 163.367
R383 B.n297 B.n54 163.367
R384 B.n301 B.n54 163.367
R385 B.n302 B.n301 163.367
R386 B.n303 B.n302 163.367
R387 B.n303 B.n52 163.367
R388 B.n307 B.n52 163.367
R389 B.n308 B.n307 163.367
R390 B.n309 B.n308 163.367
R391 B.n309 B.n50 163.367
R392 B.n313 B.n50 163.367
R393 B.n314 B.n313 163.367
R394 B.n315 B.n314 163.367
R395 B.n315 B.n48 163.367
R396 B.n319 B.n48 163.367
R397 B.n320 B.n319 163.367
R398 B.n321 B.n320 163.367
R399 B.n321 B.n46 163.367
R400 B.n325 B.n46 163.367
R401 B.n326 B.n325 163.367
R402 B.n327 B.n326 163.367
R403 B.n327 B.n44 163.367
R404 B.n392 B.n19 163.367
R405 B.n388 B.n19 163.367
R406 B.n388 B.n387 163.367
R407 B.n387 B.n386 163.367
R408 B.n386 B.n21 163.367
R409 B.n382 B.n21 163.367
R410 B.n382 B.n381 163.367
R411 B.n381 B.n380 163.367
R412 B.n380 B.n23 163.367
R413 B.n376 B.n23 163.367
R414 B.n376 B.n375 163.367
R415 B.n375 B.n374 163.367
R416 B.n374 B.n25 163.367
R417 B.n370 B.n25 163.367
R418 B.n370 B.n369 163.367
R419 B.n369 B.n368 163.367
R420 B.n368 B.n27 163.367
R421 B.n364 B.n27 163.367
R422 B.n364 B.n363 163.367
R423 B.n363 B.n362 163.367
R424 B.n362 B.n32 163.367
R425 B.n358 B.n32 163.367
R426 B.n358 B.n357 163.367
R427 B.n357 B.n356 163.367
R428 B.n356 B.n34 163.367
R429 B.n351 B.n34 163.367
R430 B.n351 B.n350 163.367
R431 B.n350 B.n349 163.367
R432 B.n349 B.n38 163.367
R433 B.n345 B.n38 163.367
R434 B.n345 B.n344 163.367
R435 B.n344 B.n343 163.367
R436 B.n343 B.n40 163.367
R437 B.n339 B.n40 163.367
R438 B.n339 B.n338 163.367
R439 B.n338 B.n337 163.367
R440 B.n337 B.n42 163.367
R441 B.n333 B.n42 163.367
R442 B.n333 B.n332 163.367
R443 B.n332 B.n331 163.367
R444 B.n203 B.n202 59.5399
R445 B.n188 B.n92 59.5399
R446 B.n30 B.n29 59.5399
R447 B.n354 B.n36 59.5399
R448 B.n202 B.n201 54.6914
R449 B.n92 B.n91 54.6914
R450 B.n29 B.n28 54.6914
R451 B.n36 B.n35 54.6914
R452 B.n391 B.n18 30.4395
R453 B.n330 B.n329 30.4395
R454 B.n228 B.n77 30.4395
R455 B.n164 B.n163 30.4395
R456 B B.n443 18.0485
R457 B.n391 B.n390 10.6151
R458 B.n390 B.n389 10.6151
R459 B.n389 B.n20 10.6151
R460 B.n385 B.n20 10.6151
R461 B.n385 B.n384 10.6151
R462 B.n384 B.n383 10.6151
R463 B.n383 B.n22 10.6151
R464 B.n379 B.n22 10.6151
R465 B.n379 B.n378 10.6151
R466 B.n378 B.n377 10.6151
R467 B.n377 B.n24 10.6151
R468 B.n373 B.n24 10.6151
R469 B.n373 B.n372 10.6151
R470 B.n372 B.n371 10.6151
R471 B.n371 B.n26 10.6151
R472 B.n367 B.n366 10.6151
R473 B.n366 B.n365 10.6151
R474 B.n365 B.n31 10.6151
R475 B.n361 B.n31 10.6151
R476 B.n361 B.n360 10.6151
R477 B.n360 B.n359 10.6151
R478 B.n359 B.n33 10.6151
R479 B.n355 B.n33 10.6151
R480 B.n353 B.n352 10.6151
R481 B.n352 B.n37 10.6151
R482 B.n348 B.n37 10.6151
R483 B.n348 B.n347 10.6151
R484 B.n347 B.n346 10.6151
R485 B.n346 B.n39 10.6151
R486 B.n342 B.n39 10.6151
R487 B.n342 B.n341 10.6151
R488 B.n341 B.n340 10.6151
R489 B.n340 B.n41 10.6151
R490 B.n336 B.n41 10.6151
R491 B.n336 B.n335 10.6151
R492 B.n335 B.n334 10.6151
R493 B.n334 B.n43 10.6151
R494 B.n330 B.n43 10.6151
R495 B.n232 B.n77 10.6151
R496 B.n233 B.n232 10.6151
R497 B.n234 B.n233 10.6151
R498 B.n234 B.n75 10.6151
R499 B.n238 B.n75 10.6151
R500 B.n239 B.n238 10.6151
R501 B.n240 B.n239 10.6151
R502 B.n240 B.n73 10.6151
R503 B.n244 B.n73 10.6151
R504 B.n245 B.n244 10.6151
R505 B.n246 B.n245 10.6151
R506 B.n246 B.n71 10.6151
R507 B.n250 B.n71 10.6151
R508 B.n251 B.n250 10.6151
R509 B.n252 B.n251 10.6151
R510 B.n252 B.n69 10.6151
R511 B.n256 B.n69 10.6151
R512 B.n257 B.n256 10.6151
R513 B.n258 B.n257 10.6151
R514 B.n258 B.n67 10.6151
R515 B.n262 B.n67 10.6151
R516 B.n263 B.n262 10.6151
R517 B.n264 B.n263 10.6151
R518 B.n264 B.n65 10.6151
R519 B.n268 B.n65 10.6151
R520 B.n269 B.n268 10.6151
R521 B.n270 B.n269 10.6151
R522 B.n270 B.n63 10.6151
R523 B.n274 B.n63 10.6151
R524 B.n275 B.n274 10.6151
R525 B.n276 B.n275 10.6151
R526 B.n276 B.n61 10.6151
R527 B.n280 B.n61 10.6151
R528 B.n281 B.n280 10.6151
R529 B.n282 B.n281 10.6151
R530 B.n282 B.n59 10.6151
R531 B.n286 B.n59 10.6151
R532 B.n287 B.n286 10.6151
R533 B.n288 B.n287 10.6151
R534 B.n288 B.n57 10.6151
R535 B.n292 B.n57 10.6151
R536 B.n293 B.n292 10.6151
R537 B.n294 B.n293 10.6151
R538 B.n294 B.n55 10.6151
R539 B.n298 B.n55 10.6151
R540 B.n299 B.n298 10.6151
R541 B.n300 B.n299 10.6151
R542 B.n300 B.n53 10.6151
R543 B.n304 B.n53 10.6151
R544 B.n305 B.n304 10.6151
R545 B.n306 B.n305 10.6151
R546 B.n306 B.n51 10.6151
R547 B.n310 B.n51 10.6151
R548 B.n311 B.n310 10.6151
R549 B.n312 B.n311 10.6151
R550 B.n312 B.n49 10.6151
R551 B.n316 B.n49 10.6151
R552 B.n317 B.n316 10.6151
R553 B.n318 B.n317 10.6151
R554 B.n318 B.n47 10.6151
R555 B.n322 B.n47 10.6151
R556 B.n323 B.n322 10.6151
R557 B.n324 B.n323 10.6151
R558 B.n324 B.n45 10.6151
R559 B.n328 B.n45 10.6151
R560 B.n329 B.n328 10.6151
R561 B.n164 B.n99 10.6151
R562 B.n168 B.n99 10.6151
R563 B.n169 B.n168 10.6151
R564 B.n170 B.n169 10.6151
R565 B.n170 B.n97 10.6151
R566 B.n174 B.n97 10.6151
R567 B.n175 B.n174 10.6151
R568 B.n176 B.n175 10.6151
R569 B.n176 B.n95 10.6151
R570 B.n180 B.n95 10.6151
R571 B.n181 B.n180 10.6151
R572 B.n182 B.n181 10.6151
R573 B.n182 B.n93 10.6151
R574 B.n186 B.n93 10.6151
R575 B.n187 B.n186 10.6151
R576 B.n189 B.n89 10.6151
R577 B.n193 B.n89 10.6151
R578 B.n194 B.n193 10.6151
R579 B.n195 B.n194 10.6151
R580 B.n195 B.n87 10.6151
R581 B.n199 B.n87 10.6151
R582 B.n200 B.n199 10.6151
R583 B.n204 B.n200 10.6151
R584 B.n208 B.n85 10.6151
R585 B.n209 B.n208 10.6151
R586 B.n210 B.n209 10.6151
R587 B.n210 B.n83 10.6151
R588 B.n214 B.n83 10.6151
R589 B.n215 B.n214 10.6151
R590 B.n216 B.n215 10.6151
R591 B.n216 B.n81 10.6151
R592 B.n220 B.n81 10.6151
R593 B.n221 B.n220 10.6151
R594 B.n222 B.n221 10.6151
R595 B.n222 B.n79 10.6151
R596 B.n226 B.n79 10.6151
R597 B.n227 B.n226 10.6151
R598 B.n228 B.n227 10.6151
R599 B.n163 B.n162 10.6151
R600 B.n162 B.n101 10.6151
R601 B.n158 B.n101 10.6151
R602 B.n158 B.n157 10.6151
R603 B.n157 B.n156 10.6151
R604 B.n156 B.n103 10.6151
R605 B.n152 B.n103 10.6151
R606 B.n152 B.n151 10.6151
R607 B.n151 B.n150 10.6151
R608 B.n150 B.n105 10.6151
R609 B.n146 B.n105 10.6151
R610 B.n146 B.n145 10.6151
R611 B.n145 B.n144 10.6151
R612 B.n144 B.n107 10.6151
R613 B.n140 B.n107 10.6151
R614 B.n140 B.n139 10.6151
R615 B.n139 B.n138 10.6151
R616 B.n138 B.n109 10.6151
R617 B.n134 B.n109 10.6151
R618 B.n134 B.n133 10.6151
R619 B.n133 B.n132 10.6151
R620 B.n132 B.n111 10.6151
R621 B.n128 B.n111 10.6151
R622 B.n128 B.n127 10.6151
R623 B.n127 B.n126 10.6151
R624 B.n126 B.n113 10.6151
R625 B.n122 B.n113 10.6151
R626 B.n122 B.n121 10.6151
R627 B.n121 B.n120 10.6151
R628 B.n120 B.n115 10.6151
R629 B.n116 B.n115 10.6151
R630 B.n116 B.n0 10.6151
R631 B.n439 B.n1 10.6151
R632 B.n439 B.n438 10.6151
R633 B.n438 B.n437 10.6151
R634 B.n437 B.n4 10.6151
R635 B.n433 B.n4 10.6151
R636 B.n433 B.n432 10.6151
R637 B.n432 B.n431 10.6151
R638 B.n431 B.n6 10.6151
R639 B.n427 B.n6 10.6151
R640 B.n427 B.n426 10.6151
R641 B.n426 B.n425 10.6151
R642 B.n425 B.n8 10.6151
R643 B.n421 B.n8 10.6151
R644 B.n421 B.n420 10.6151
R645 B.n420 B.n419 10.6151
R646 B.n419 B.n10 10.6151
R647 B.n415 B.n10 10.6151
R648 B.n415 B.n414 10.6151
R649 B.n414 B.n413 10.6151
R650 B.n413 B.n12 10.6151
R651 B.n409 B.n12 10.6151
R652 B.n409 B.n408 10.6151
R653 B.n408 B.n407 10.6151
R654 B.n407 B.n14 10.6151
R655 B.n403 B.n14 10.6151
R656 B.n403 B.n402 10.6151
R657 B.n402 B.n401 10.6151
R658 B.n401 B.n16 10.6151
R659 B.n397 B.n16 10.6151
R660 B.n397 B.n396 10.6151
R661 B.n396 B.n395 10.6151
R662 B.n395 B.n18 10.6151
R663 B.n367 B.n30 6.5566
R664 B.n355 B.n354 6.5566
R665 B.n189 B.n188 6.5566
R666 B.n204 B.n203 6.5566
R667 B.n30 B.n26 4.05904
R668 B.n354 B.n353 4.05904
R669 B.n188 B.n187 4.05904
R670 B.n203 B.n85 4.05904
R671 B.n443 B.n0 2.81026
R672 B.n443 B.n1 2.81026
R673 VN.n0 VN.t1 65.6408
R674 VN.n1 VN.t3 65.6408
R675 VN.n0 VN.t0 64.885
R676 VN.n1 VN.t2 64.885
R677 VN VN.n1 44.0224
R678 VN VN.n0 4.54889
R679 VTAIL.n122 VTAIL.n112 756.745
R680 VTAIL.n10 VTAIL.n0 756.745
R681 VTAIL.n26 VTAIL.n16 756.745
R682 VTAIL.n42 VTAIL.n32 756.745
R683 VTAIL.n106 VTAIL.n96 756.745
R684 VTAIL.n90 VTAIL.n80 756.745
R685 VTAIL.n74 VTAIL.n64 756.745
R686 VTAIL.n58 VTAIL.n48 756.745
R687 VTAIL.n116 VTAIL.n115 585
R688 VTAIL.n121 VTAIL.n120 585
R689 VTAIL.n123 VTAIL.n122 585
R690 VTAIL.n4 VTAIL.n3 585
R691 VTAIL.n9 VTAIL.n8 585
R692 VTAIL.n11 VTAIL.n10 585
R693 VTAIL.n20 VTAIL.n19 585
R694 VTAIL.n25 VTAIL.n24 585
R695 VTAIL.n27 VTAIL.n26 585
R696 VTAIL.n36 VTAIL.n35 585
R697 VTAIL.n41 VTAIL.n40 585
R698 VTAIL.n43 VTAIL.n42 585
R699 VTAIL.n107 VTAIL.n106 585
R700 VTAIL.n105 VTAIL.n104 585
R701 VTAIL.n100 VTAIL.n99 585
R702 VTAIL.n91 VTAIL.n90 585
R703 VTAIL.n89 VTAIL.n88 585
R704 VTAIL.n84 VTAIL.n83 585
R705 VTAIL.n75 VTAIL.n74 585
R706 VTAIL.n73 VTAIL.n72 585
R707 VTAIL.n68 VTAIL.n67 585
R708 VTAIL.n59 VTAIL.n58 585
R709 VTAIL.n57 VTAIL.n56 585
R710 VTAIL.n52 VTAIL.n51 585
R711 VTAIL.n117 VTAIL.t7 336.901
R712 VTAIL.n5 VTAIL.t4 336.901
R713 VTAIL.n21 VTAIL.t3 336.901
R714 VTAIL.n37 VTAIL.t0 336.901
R715 VTAIL.n101 VTAIL.t1 336.901
R716 VTAIL.n85 VTAIL.t2 336.901
R717 VTAIL.n69 VTAIL.t6 336.901
R718 VTAIL.n53 VTAIL.t5 336.901
R719 VTAIL.n121 VTAIL.n115 171.744
R720 VTAIL.n122 VTAIL.n121 171.744
R721 VTAIL.n9 VTAIL.n3 171.744
R722 VTAIL.n10 VTAIL.n9 171.744
R723 VTAIL.n25 VTAIL.n19 171.744
R724 VTAIL.n26 VTAIL.n25 171.744
R725 VTAIL.n41 VTAIL.n35 171.744
R726 VTAIL.n42 VTAIL.n41 171.744
R727 VTAIL.n106 VTAIL.n105 171.744
R728 VTAIL.n105 VTAIL.n99 171.744
R729 VTAIL.n90 VTAIL.n89 171.744
R730 VTAIL.n89 VTAIL.n83 171.744
R731 VTAIL.n74 VTAIL.n73 171.744
R732 VTAIL.n73 VTAIL.n67 171.744
R733 VTAIL.n58 VTAIL.n57 171.744
R734 VTAIL.n57 VTAIL.n51 171.744
R735 VTAIL.t7 VTAIL.n115 85.8723
R736 VTAIL.t4 VTAIL.n3 85.8723
R737 VTAIL.t3 VTAIL.n19 85.8723
R738 VTAIL.t0 VTAIL.n35 85.8723
R739 VTAIL.t1 VTAIL.n99 85.8723
R740 VTAIL.t2 VTAIL.n83 85.8723
R741 VTAIL.t6 VTAIL.n67 85.8723
R742 VTAIL.t5 VTAIL.n51 85.8723
R743 VTAIL.n127 VTAIL.n126 32.3793
R744 VTAIL.n15 VTAIL.n14 32.3793
R745 VTAIL.n31 VTAIL.n30 32.3793
R746 VTAIL.n47 VTAIL.n46 32.3793
R747 VTAIL.n111 VTAIL.n110 32.3793
R748 VTAIL.n95 VTAIL.n94 32.3793
R749 VTAIL.n79 VTAIL.n78 32.3793
R750 VTAIL.n63 VTAIL.n62 32.3793
R751 VTAIL.n127 VTAIL.n111 17.4962
R752 VTAIL.n63 VTAIL.n47 17.4962
R753 VTAIL.n117 VTAIL.n116 16.193
R754 VTAIL.n5 VTAIL.n4 16.193
R755 VTAIL.n21 VTAIL.n20 16.193
R756 VTAIL.n37 VTAIL.n36 16.193
R757 VTAIL.n101 VTAIL.n100 16.193
R758 VTAIL.n85 VTAIL.n84 16.193
R759 VTAIL.n69 VTAIL.n68 16.193
R760 VTAIL.n53 VTAIL.n52 16.193
R761 VTAIL.n120 VTAIL.n119 12.8005
R762 VTAIL.n8 VTAIL.n7 12.8005
R763 VTAIL.n24 VTAIL.n23 12.8005
R764 VTAIL.n40 VTAIL.n39 12.8005
R765 VTAIL.n104 VTAIL.n103 12.8005
R766 VTAIL.n88 VTAIL.n87 12.8005
R767 VTAIL.n72 VTAIL.n71 12.8005
R768 VTAIL.n56 VTAIL.n55 12.8005
R769 VTAIL.n123 VTAIL.n114 12.0247
R770 VTAIL.n11 VTAIL.n2 12.0247
R771 VTAIL.n27 VTAIL.n18 12.0247
R772 VTAIL.n43 VTAIL.n34 12.0247
R773 VTAIL.n107 VTAIL.n98 12.0247
R774 VTAIL.n91 VTAIL.n82 12.0247
R775 VTAIL.n75 VTAIL.n66 12.0247
R776 VTAIL.n59 VTAIL.n50 12.0247
R777 VTAIL.n124 VTAIL.n112 11.249
R778 VTAIL.n12 VTAIL.n0 11.249
R779 VTAIL.n28 VTAIL.n16 11.249
R780 VTAIL.n44 VTAIL.n32 11.249
R781 VTAIL.n108 VTAIL.n96 11.249
R782 VTAIL.n92 VTAIL.n80 11.249
R783 VTAIL.n76 VTAIL.n64 11.249
R784 VTAIL.n60 VTAIL.n48 11.249
R785 VTAIL.n126 VTAIL.n125 9.45567
R786 VTAIL.n14 VTAIL.n13 9.45567
R787 VTAIL.n30 VTAIL.n29 9.45567
R788 VTAIL.n46 VTAIL.n45 9.45567
R789 VTAIL.n110 VTAIL.n109 9.45567
R790 VTAIL.n94 VTAIL.n93 9.45567
R791 VTAIL.n78 VTAIL.n77 9.45567
R792 VTAIL.n62 VTAIL.n61 9.45567
R793 VTAIL.n125 VTAIL.n124 9.3005
R794 VTAIL.n114 VTAIL.n113 9.3005
R795 VTAIL.n119 VTAIL.n118 9.3005
R796 VTAIL.n13 VTAIL.n12 9.3005
R797 VTAIL.n2 VTAIL.n1 9.3005
R798 VTAIL.n7 VTAIL.n6 9.3005
R799 VTAIL.n29 VTAIL.n28 9.3005
R800 VTAIL.n18 VTAIL.n17 9.3005
R801 VTAIL.n23 VTAIL.n22 9.3005
R802 VTAIL.n45 VTAIL.n44 9.3005
R803 VTAIL.n34 VTAIL.n33 9.3005
R804 VTAIL.n39 VTAIL.n38 9.3005
R805 VTAIL.n109 VTAIL.n108 9.3005
R806 VTAIL.n98 VTAIL.n97 9.3005
R807 VTAIL.n103 VTAIL.n102 9.3005
R808 VTAIL.n93 VTAIL.n92 9.3005
R809 VTAIL.n82 VTAIL.n81 9.3005
R810 VTAIL.n87 VTAIL.n86 9.3005
R811 VTAIL.n77 VTAIL.n76 9.3005
R812 VTAIL.n66 VTAIL.n65 9.3005
R813 VTAIL.n71 VTAIL.n70 9.3005
R814 VTAIL.n61 VTAIL.n60 9.3005
R815 VTAIL.n50 VTAIL.n49 9.3005
R816 VTAIL.n55 VTAIL.n54 9.3005
R817 VTAIL.n102 VTAIL.n101 3.91276
R818 VTAIL.n86 VTAIL.n85 3.91276
R819 VTAIL.n70 VTAIL.n69 3.91276
R820 VTAIL.n54 VTAIL.n53 3.91276
R821 VTAIL.n118 VTAIL.n117 3.91276
R822 VTAIL.n6 VTAIL.n5 3.91276
R823 VTAIL.n22 VTAIL.n21 3.91276
R824 VTAIL.n38 VTAIL.n37 3.91276
R825 VTAIL.n126 VTAIL.n112 2.71565
R826 VTAIL.n14 VTAIL.n0 2.71565
R827 VTAIL.n30 VTAIL.n16 2.71565
R828 VTAIL.n46 VTAIL.n32 2.71565
R829 VTAIL.n110 VTAIL.n96 2.71565
R830 VTAIL.n94 VTAIL.n80 2.71565
R831 VTAIL.n78 VTAIL.n64 2.71565
R832 VTAIL.n62 VTAIL.n48 2.71565
R833 VTAIL.n79 VTAIL.n63 2.43153
R834 VTAIL.n111 VTAIL.n95 2.43153
R835 VTAIL.n47 VTAIL.n31 2.43153
R836 VTAIL.n124 VTAIL.n123 1.93989
R837 VTAIL.n12 VTAIL.n11 1.93989
R838 VTAIL.n28 VTAIL.n27 1.93989
R839 VTAIL.n44 VTAIL.n43 1.93989
R840 VTAIL.n108 VTAIL.n107 1.93989
R841 VTAIL.n92 VTAIL.n91 1.93989
R842 VTAIL.n76 VTAIL.n75 1.93989
R843 VTAIL.n60 VTAIL.n59 1.93989
R844 VTAIL VTAIL.n15 1.27421
R845 VTAIL.n120 VTAIL.n114 1.16414
R846 VTAIL.n8 VTAIL.n2 1.16414
R847 VTAIL.n24 VTAIL.n18 1.16414
R848 VTAIL.n40 VTAIL.n34 1.16414
R849 VTAIL.n104 VTAIL.n98 1.16414
R850 VTAIL.n88 VTAIL.n82 1.16414
R851 VTAIL.n72 VTAIL.n66 1.16414
R852 VTAIL.n56 VTAIL.n50 1.16414
R853 VTAIL VTAIL.n127 1.15783
R854 VTAIL.n95 VTAIL.n79 0.470328
R855 VTAIL.n31 VTAIL.n15 0.470328
R856 VTAIL.n119 VTAIL.n116 0.388379
R857 VTAIL.n7 VTAIL.n4 0.388379
R858 VTAIL.n23 VTAIL.n20 0.388379
R859 VTAIL.n39 VTAIL.n36 0.388379
R860 VTAIL.n103 VTAIL.n100 0.388379
R861 VTAIL.n87 VTAIL.n84 0.388379
R862 VTAIL.n71 VTAIL.n68 0.388379
R863 VTAIL.n55 VTAIL.n52 0.388379
R864 VTAIL.n118 VTAIL.n113 0.155672
R865 VTAIL.n125 VTAIL.n113 0.155672
R866 VTAIL.n6 VTAIL.n1 0.155672
R867 VTAIL.n13 VTAIL.n1 0.155672
R868 VTAIL.n22 VTAIL.n17 0.155672
R869 VTAIL.n29 VTAIL.n17 0.155672
R870 VTAIL.n38 VTAIL.n33 0.155672
R871 VTAIL.n45 VTAIL.n33 0.155672
R872 VTAIL.n109 VTAIL.n97 0.155672
R873 VTAIL.n102 VTAIL.n97 0.155672
R874 VTAIL.n93 VTAIL.n81 0.155672
R875 VTAIL.n86 VTAIL.n81 0.155672
R876 VTAIL.n77 VTAIL.n65 0.155672
R877 VTAIL.n70 VTAIL.n65 0.155672
R878 VTAIL.n61 VTAIL.n49 0.155672
R879 VTAIL.n54 VTAIL.n49 0.155672
R880 VDD2.n2 VDD2.n0 161.75
R881 VDD2.n2 VDD2.n1 128.044
R882 VDD2.n1 VDD2.t1 10.3855
R883 VDD2.n1 VDD2.t0 10.3855
R884 VDD2.n0 VDD2.t2 10.3855
R885 VDD2.n0 VDD2.t3 10.3855
R886 VDD2 VDD2.n2 0.0586897
R887 VP.n14 VP.n0 161.3
R888 VP.n13 VP.n12 161.3
R889 VP.n11 VP.n1 161.3
R890 VP.n10 VP.n9 161.3
R891 VP.n8 VP.n2 161.3
R892 VP.n7 VP.n6 161.3
R893 VP.n5 VP.n3 102.927
R894 VP.n16 VP.n15 102.927
R895 VP.n4 VP.t1 65.6408
R896 VP.n4 VP.t0 64.885
R897 VP.n9 VP.n1 56.5193
R898 VP.n5 VP.n4 43.7435
R899 VP.n3 VP.t3 30.2949
R900 VP.n15 VP.t2 30.2949
R901 VP.n8 VP.n7 24.4675
R902 VP.n9 VP.n8 24.4675
R903 VP.n13 VP.n1 24.4675
R904 VP.n14 VP.n13 24.4675
R905 VP.n7 VP.n3 7.82994
R906 VP.n15 VP.n14 7.82994
R907 VP.n6 VP.n5 0.278367
R908 VP.n16 VP.n0 0.278367
R909 VP.n6 VP.n2 0.189894
R910 VP.n10 VP.n2 0.189894
R911 VP.n11 VP.n10 0.189894
R912 VP.n12 VP.n11 0.189894
R913 VP.n12 VP.n0 0.189894
R914 VP VP.n16 0.153454
R915 VDD1 VDD1.n1 162.275
R916 VDD1 VDD1.n0 128.102
R917 VDD1.n0 VDD1.t2 10.3855
R918 VDD1.n0 VDD1.t3 10.3855
R919 VDD1.n1 VDD1.t0 10.3855
R920 VDD1.n1 VDD1.t1 10.3855
C0 VN VTAIL 1.90885f
C1 VDD2 VTAIL 3.29977f
C2 B VTAIL 1.9493f
C3 VDD1 w_n2662_n1594# 1.19427f
C4 VDD1 VP 1.70131f
C5 w_n2662_n1594# VP 4.65797f
C6 VDD1 VN 0.153842f
C7 VDD2 VDD1 1.00702f
C8 w_n2662_n1594# VN 4.31816f
C9 VDD2 w_n2662_n1594# 1.2475f
C10 VN VP 4.47726f
C11 VDD2 VP 0.392837f
C12 B VDD1 1.00165f
C13 B w_n2662_n1594# 6.64433f
C14 B VP 1.54474f
C15 VDD2 VN 1.46369f
C16 VDD1 VTAIL 3.2463f
C17 B VN 0.978219f
C18 w_n2662_n1594# VTAIL 1.94378f
C19 B VDD2 1.05217f
C20 VTAIL VP 1.92296f
C21 VDD2 VSUBS 0.640861f
C22 VDD1 VSUBS 3.193252f
C23 VTAIL VSUBS 0.450404f
C24 VN VSUBS 4.69349f
C25 VP VSUBS 1.724829f
C26 B VSUBS 3.244775f
C27 w_n2662_n1594# VSUBS 53.6979f
C28 VDD1.t2 VSUBS 0.046028f
C29 VDD1.t3 VSUBS 0.046028f
C30 VDD1.n0 VSUBS 0.24683f
C31 VDD1.t0 VSUBS 0.046028f
C32 VDD1.t1 VSUBS 0.046028f
C33 VDD1.n1 VSUBS 0.431649f
C34 VP.n0 VSUBS 0.051044f
C35 VP.t2 VSUBS 0.755584f
C36 VP.n1 VSUBS 0.05652f
C37 VP.n2 VSUBS 0.038717f
C38 VP.t3 VSUBS 0.755584f
C39 VP.n3 VSUBS 0.437048f
C40 VP.t0 VSUBS 1.05018f
C41 VP.t1 VSUBS 1.05655f
C42 VP.n4 VSUBS 2.29294f
C43 VP.n5 VSUBS 1.69691f
C44 VP.n6 VSUBS 0.051044f
C45 VP.n7 VSUBS 0.047934f
C46 VP.n8 VSUBS 0.072159f
C47 VP.n9 VSUBS 0.05652f
C48 VP.n10 VSUBS 0.038717f
C49 VP.n11 VSUBS 0.038717f
C50 VP.n12 VSUBS 0.038717f
C51 VP.n13 VSUBS 0.072159f
C52 VP.n14 VSUBS 0.047934f
C53 VP.n15 VSUBS 0.437048f
C54 VP.n16 VSUBS 0.06362f
C55 VDD2.t2 VSUBS 0.048508f
C56 VDD2.t3 VSUBS 0.048508f
C57 VDD2.n0 VSUBS 0.444264f
C58 VDD2.t1 VSUBS 0.048508f
C59 VDD2.t0 VSUBS 0.048508f
C60 VDD2.n1 VSUBS 0.259942f
C61 VDD2.n2 VSUBS 2.24391f
C62 VTAIL.n0 VSUBS 0.0152f
C63 VTAIL.n1 VSUBS 0.014743f
C64 VTAIL.n2 VSUBS 0.007922f
C65 VTAIL.n3 VSUBS 0.014044f
C66 VTAIL.n4 VSUBS 0.01156f
C67 VTAIL.t4 VSUBS 0.041285f
C68 VTAIL.n5 VSUBS 0.052812f
C69 VTAIL.n6 VSUBS 0.145131f
C70 VTAIL.n7 VSUBS 0.007922f
C71 VTAIL.n8 VSUBS 0.008388f
C72 VTAIL.n9 VSUBS 0.018725f
C73 VTAIL.n10 VSUBS 0.041928f
C74 VTAIL.n11 VSUBS 0.008388f
C75 VTAIL.n12 VSUBS 0.007922f
C76 VTAIL.n13 VSUBS 0.034278f
C77 VTAIL.n14 VSUBS 0.02094f
C78 VTAIL.n15 VSUBS 0.09553f
C79 VTAIL.n16 VSUBS 0.0152f
C80 VTAIL.n17 VSUBS 0.014743f
C81 VTAIL.n18 VSUBS 0.007922f
C82 VTAIL.n19 VSUBS 0.014044f
C83 VTAIL.n20 VSUBS 0.01156f
C84 VTAIL.t3 VSUBS 0.041285f
C85 VTAIL.n21 VSUBS 0.052812f
C86 VTAIL.n22 VSUBS 0.145131f
C87 VTAIL.n23 VSUBS 0.007922f
C88 VTAIL.n24 VSUBS 0.008388f
C89 VTAIL.n25 VSUBS 0.018725f
C90 VTAIL.n26 VSUBS 0.041928f
C91 VTAIL.n27 VSUBS 0.008388f
C92 VTAIL.n28 VSUBS 0.007922f
C93 VTAIL.n29 VSUBS 0.034278f
C94 VTAIL.n30 VSUBS 0.02094f
C95 VTAIL.n31 VSUBS 0.150508f
C96 VTAIL.n32 VSUBS 0.0152f
C97 VTAIL.n33 VSUBS 0.014743f
C98 VTAIL.n34 VSUBS 0.007922f
C99 VTAIL.n35 VSUBS 0.014044f
C100 VTAIL.n36 VSUBS 0.01156f
C101 VTAIL.t0 VSUBS 0.041285f
C102 VTAIL.n37 VSUBS 0.052812f
C103 VTAIL.n38 VSUBS 0.145131f
C104 VTAIL.n39 VSUBS 0.007922f
C105 VTAIL.n40 VSUBS 0.008388f
C106 VTAIL.n41 VSUBS 0.018725f
C107 VTAIL.n42 VSUBS 0.041928f
C108 VTAIL.n43 VSUBS 0.008388f
C109 VTAIL.n44 VSUBS 0.007922f
C110 VTAIL.n45 VSUBS 0.034278f
C111 VTAIL.n46 VSUBS 0.02094f
C112 VTAIL.n47 VSUBS 0.572115f
C113 VTAIL.n48 VSUBS 0.0152f
C114 VTAIL.n49 VSUBS 0.014743f
C115 VTAIL.n50 VSUBS 0.007922f
C116 VTAIL.n51 VSUBS 0.014044f
C117 VTAIL.n52 VSUBS 0.01156f
C118 VTAIL.t5 VSUBS 0.041285f
C119 VTAIL.n53 VSUBS 0.052812f
C120 VTAIL.n54 VSUBS 0.145131f
C121 VTAIL.n55 VSUBS 0.007922f
C122 VTAIL.n56 VSUBS 0.008388f
C123 VTAIL.n57 VSUBS 0.018725f
C124 VTAIL.n58 VSUBS 0.041928f
C125 VTAIL.n59 VSUBS 0.008388f
C126 VTAIL.n60 VSUBS 0.007922f
C127 VTAIL.n61 VSUBS 0.034278f
C128 VTAIL.n62 VSUBS 0.02094f
C129 VTAIL.n63 VSUBS 0.572115f
C130 VTAIL.n64 VSUBS 0.0152f
C131 VTAIL.n65 VSUBS 0.014743f
C132 VTAIL.n66 VSUBS 0.007922f
C133 VTAIL.n67 VSUBS 0.014044f
C134 VTAIL.n68 VSUBS 0.01156f
C135 VTAIL.t6 VSUBS 0.041285f
C136 VTAIL.n69 VSUBS 0.052812f
C137 VTAIL.n70 VSUBS 0.145131f
C138 VTAIL.n71 VSUBS 0.007922f
C139 VTAIL.n72 VSUBS 0.008388f
C140 VTAIL.n73 VSUBS 0.018725f
C141 VTAIL.n74 VSUBS 0.041928f
C142 VTAIL.n75 VSUBS 0.008388f
C143 VTAIL.n76 VSUBS 0.007922f
C144 VTAIL.n77 VSUBS 0.034278f
C145 VTAIL.n78 VSUBS 0.02094f
C146 VTAIL.n79 VSUBS 0.150508f
C147 VTAIL.n80 VSUBS 0.0152f
C148 VTAIL.n81 VSUBS 0.014743f
C149 VTAIL.n82 VSUBS 0.007922f
C150 VTAIL.n83 VSUBS 0.014044f
C151 VTAIL.n84 VSUBS 0.01156f
C152 VTAIL.t2 VSUBS 0.041285f
C153 VTAIL.n85 VSUBS 0.052812f
C154 VTAIL.n86 VSUBS 0.145131f
C155 VTAIL.n87 VSUBS 0.007922f
C156 VTAIL.n88 VSUBS 0.008388f
C157 VTAIL.n89 VSUBS 0.018725f
C158 VTAIL.n90 VSUBS 0.041928f
C159 VTAIL.n91 VSUBS 0.008388f
C160 VTAIL.n92 VSUBS 0.007922f
C161 VTAIL.n93 VSUBS 0.034278f
C162 VTAIL.n94 VSUBS 0.02094f
C163 VTAIL.n95 VSUBS 0.150508f
C164 VTAIL.n96 VSUBS 0.0152f
C165 VTAIL.n97 VSUBS 0.014743f
C166 VTAIL.n98 VSUBS 0.007922f
C167 VTAIL.n99 VSUBS 0.014044f
C168 VTAIL.n100 VSUBS 0.01156f
C169 VTAIL.t1 VSUBS 0.041285f
C170 VTAIL.n101 VSUBS 0.052812f
C171 VTAIL.n102 VSUBS 0.145131f
C172 VTAIL.n103 VSUBS 0.007922f
C173 VTAIL.n104 VSUBS 0.008388f
C174 VTAIL.n105 VSUBS 0.018725f
C175 VTAIL.n106 VSUBS 0.041928f
C176 VTAIL.n107 VSUBS 0.008388f
C177 VTAIL.n108 VSUBS 0.007922f
C178 VTAIL.n109 VSUBS 0.034278f
C179 VTAIL.n110 VSUBS 0.02094f
C180 VTAIL.n111 VSUBS 0.572115f
C181 VTAIL.n112 VSUBS 0.0152f
C182 VTAIL.n113 VSUBS 0.014743f
C183 VTAIL.n114 VSUBS 0.007922f
C184 VTAIL.n115 VSUBS 0.014044f
C185 VTAIL.n116 VSUBS 0.01156f
C186 VTAIL.t7 VSUBS 0.041285f
C187 VTAIL.n117 VSUBS 0.052812f
C188 VTAIL.n118 VSUBS 0.145131f
C189 VTAIL.n119 VSUBS 0.007922f
C190 VTAIL.n120 VSUBS 0.008388f
C191 VTAIL.n121 VSUBS 0.018725f
C192 VTAIL.n122 VSUBS 0.041928f
C193 VTAIL.n123 VSUBS 0.008388f
C194 VTAIL.n124 VSUBS 0.007922f
C195 VTAIL.n125 VSUBS 0.034278f
C196 VTAIL.n126 VSUBS 0.02094f
C197 VTAIL.n127 VSUBS 0.511609f
C198 VN.t1 VSUBS 1.00467f
C199 VN.t0 VSUBS 0.998609f
C200 VN.n0 VSUBS 0.63851f
C201 VN.t3 VSUBS 1.00467f
C202 VN.t2 VSUBS 0.998609f
C203 VN.n1 VSUBS 2.20003f
C204 B.n0 VSUBS 0.004869f
C205 B.n1 VSUBS 0.004869f
C206 B.n2 VSUBS 0.0077f
C207 B.n3 VSUBS 0.0077f
C208 B.n4 VSUBS 0.0077f
C209 B.n5 VSUBS 0.0077f
C210 B.n6 VSUBS 0.0077f
C211 B.n7 VSUBS 0.0077f
C212 B.n8 VSUBS 0.0077f
C213 B.n9 VSUBS 0.0077f
C214 B.n10 VSUBS 0.0077f
C215 B.n11 VSUBS 0.0077f
C216 B.n12 VSUBS 0.0077f
C217 B.n13 VSUBS 0.0077f
C218 B.n14 VSUBS 0.0077f
C219 B.n15 VSUBS 0.0077f
C220 B.n16 VSUBS 0.0077f
C221 B.n17 VSUBS 0.0077f
C222 B.n18 VSUBS 0.016604f
C223 B.n19 VSUBS 0.0077f
C224 B.n20 VSUBS 0.0077f
C225 B.n21 VSUBS 0.0077f
C226 B.n22 VSUBS 0.0077f
C227 B.n23 VSUBS 0.0077f
C228 B.n24 VSUBS 0.0077f
C229 B.n25 VSUBS 0.0077f
C230 B.n26 VSUBS 0.005322f
C231 B.n27 VSUBS 0.0077f
C232 B.t5 VSUBS 0.050554f
C233 B.t4 VSUBS 0.069053f
C234 B.t3 VSUBS 0.415701f
C235 B.n28 VSUBS 0.122328f
C236 B.n29 VSUBS 0.105318f
C237 B.n30 VSUBS 0.017839f
C238 B.n31 VSUBS 0.0077f
C239 B.n32 VSUBS 0.0077f
C240 B.n33 VSUBS 0.0077f
C241 B.n34 VSUBS 0.0077f
C242 B.t11 VSUBS 0.050554f
C243 B.t10 VSUBS 0.069053f
C244 B.t9 VSUBS 0.415701f
C245 B.n35 VSUBS 0.122328f
C246 B.n36 VSUBS 0.105317f
C247 B.n37 VSUBS 0.0077f
C248 B.n38 VSUBS 0.0077f
C249 B.n39 VSUBS 0.0077f
C250 B.n40 VSUBS 0.0077f
C251 B.n41 VSUBS 0.0077f
C252 B.n42 VSUBS 0.0077f
C253 B.n43 VSUBS 0.0077f
C254 B.n44 VSUBS 0.016604f
C255 B.n45 VSUBS 0.0077f
C256 B.n46 VSUBS 0.0077f
C257 B.n47 VSUBS 0.0077f
C258 B.n48 VSUBS 0.0077f
C259 B.n49 VSUBS 0.0077f
C260 B.n50 VSUBS 0.0077f
C261 B.n51 VSUBS 0.0077f
C262 B.n52 VSUBS 0.0077f
C263 B.n53 VSUBS 0.0077f
C264 B.n54 VSUBS 0.0077f
C265 B.n55 VSUBS 0.0077f
C266 B.n56 VSUBS 0.0077f
C267 B.n57 VSUBS 0.0077f
C268 B.n58 VSUBS 0.0077f
C269 B.n59 VSUBS 0.0077f
C270 B.n60 VSUBS 0.0077f
C271 B.n61 VSUBS 0.0077f
C272 B.n62 VSUBS 0.0077f
C273 B.n63 VSUBS 0.0077f
C274 B.n64 VSUBS 0.0077f
C275 B.n65 VSUBS 0.0077f
C276 B.n66 VSUBS 0.0077f
C277 B.n67 VSUBS 0.0077f
C278 B.n68 VSUBS 0.0077f
C279 B.n69 VSUBS 0.0077f
C280 B.n70 VSUBS 0.0077f
C281 B.n71 VSUBS 0.0077f
C282 B.n72 VSUBS 0.0077f
C283 B.n73 VSUBS 0.0077f
C284 B.n74 VSUBS 0.0077f
C285 B.n75 VSUBS 0.0077f
C286 B.n76 VSUBS 0.0077f
C287 B.n77 VSUBS 0.016604f
C288 B.n78 VSUBS 0.0077f
C289 B.n79 VSUBS 0.0077f
C290 B.n80 VSUBS 0.0077f
C291 B.n81 VSUBS 0.0077f
C292 B.n82 VSUBS 0.0077f
C293 B.n83 VSUBS 0.0077f
C294 B.n84 VSUBS 0.0077f
C295 B.n85 VSUBS 0.005322f
C296 B.n86 VSUBS 0.0077f
C297 B.n87 VSUBS 0.0077f
C298 B.n88 VSUBS 0.0077f
C299 B.n89 VSUBS 0.0077f
C300 B.n90 VSUBS 0.0077f
C301 B.t1 VSUBS 0.050554f
C302 B.t2 VSUBS 0.069053f
C303 B.t0 VSUBS 0.415701f
C304 B.n91 VSUBS 0.122328f
C305 B.n92 VSUBS 0.105318f
C306 B.n93 VSUBS 0.0077f
C307 B.n94 VSUBS 0.0077f
C308 B.n95 VSUBS 0.0077f
C309 B.n96 VSUBS 0.0077f
C310 B.n97 VSUBS 0.0077f
C311 B.n98 VSUBS 0.0077f
C312 B.n99 VSUBS 0.0077f
C313 B.n100 VSUBS 0.016604f
C314 B.n101 VSUBS 0.0077f
C315 B.n102 VSUBS 0.0077f
C316 B.n103 VSUBS 0.0077f
C317 B.n104 VSUBS 0.0077f
C318 B.n105 VSUBS 0.0077f
C319 B.n106 VSUBS 0.0077f
C320 B.n107 VSUBS 0.0077f
C321 B.n108 VSUBS 0.0077f
C322 B.n109 VSUBS 0.0077f
C323 B.n110 VSUBS 0.0077f
C324 B.n111 VSUBS 0.0077f
C325 B.n112 VSUBS 0.0077f
C326 B.n113 VSUBS 0.0077f
C327 B.n114 VSUBS 0.0077f
C328 B.n115 VSUBS 0.0077f
C329 B.n116 VSUBS 0.0077f
C330 B.n117 VSUBS 0.0077f
C331 B.n118 VSUBS 0.0077f
C332 B.n119 VSUBS 0.0077f
C333 B.n120 VSUBS 0.0077f
C334 B.n121 VSUBS 0.0077f
C335 B.n122 VSUBS 0.0077f
C336 B.n123 VSUBS 0.0077f
C337 B.n124 VSUBS 0.0077f
C338 B.n125 VSUBS 0.0077f
C339 B.n126 VSUBS 0.0077f
C340 B.n127 VSUBS 0.0077f
C341 B.n128 VSUBS 0.0077f
C342 B.n129 VSUBS 0.0077f
C343 B.n130 VSUBS 0.0077f
C344 B.n131 VSUBS 0.0077f
C345 B.n132 VSUBS 0.0077f
C346 B.n133 VSUBS 0.0077f
C347 B.n134 VSUBS 0.0077f
C348 B.n135 VSUBS 0.0077f
C349 B.n136 VSUBS 0.0077f
C350 B.n137 VSUBS 0.0077f
C351 B.n138 VSUBS 0.0077f
C352 B.n139 VSUBS 0.0077f
C353 B.n140 VSUBS 0.0077f
C354 B.n141 VSUBS 0.0077f
C355 B.n142 VSUBS 0.0077f
C356 B.n143 VSUBS 0.0077f
C357 B.n144 VSUBS 0.0077f
C358 B.n145 VSUBS 0.0077f
C359 B.n146 VSUBS 0.0077f
C360 B.n147 VSUBS 0.0077f
C361 B.n148 VSUBS 0.0077f
C362 B.n149 VSUBS 0.0077f
C363 B.n150 VSUBS 0.0077f
C364 B.n151 VSUBS 0.0077f
C365 B.n152 VSUBS 0.0077f
C366 B.n153 VSUBS 0.0077f
C367 B.n154 VSUBS 0.0077f
C368 B.n155 VSUBS 0.0077f
C369 B.n156 VSUBS 0.0077f
C370 B.n157 VSUBS 0.0077f
C371 B.n158 VSUBS 0.0077f
C372 B.n159 VSUBS 0.0077f
C373 B.n160 VSUBS 0.0077f
C374 B.n161 VSUBS 0.0077f
C375 B.n162 VSUBS 0.0077f
C376 B.n163 VSUBS 0.016604f
C377 B.n164 VSUBS 0.017818f
C378 B.n165 VSUBS 0.017818f
C379 B.n166 VSUBS 0.0077f
C380 B.n167 VSUBS 0.0077f
C381 B.n168 VSUBS 0.0077f
C382 B.n169 VSUBS 0.0077f
C383 B.n170 VSUBS 0.0077f
C384 B.n171 VSUBS 0.0077f
C385 B.n172 VSUBS 0.0077f
C386 B.n173 VSUBS 0.0077f
C387 B.n174 VSUBS 0.0077f
C388 B.n175 VSUBS 0.0077f
C389 B.n176 VSUBS 0.0077f
C390 B.n177 VSUBS 0.0077f
C391 B.n178 VSUBS 0.0077f
C392 B.n179 VSUBS 0.0077f
C393 B.n180 VSUBS 0.0077f
C394 B.n181 VSUBS 0.0077f
C395 B.n182 VSUBS 0.0077f
C396 B.n183 VSUBS 0.0077f
C397 B.n184 VSUBS 0.0077f
C398 B.n185 VSUBS 0.0077f
C399 B.n186 VSUBS 0.0077f
C400 B.n187 VSUBS 0.005322f
C401 B.n188 VSUBS 0.017839f
C402 B.n189 VSUBS 0.006228f
C403 B.n190 VSUBS 0.0077f
C404 B.n191 VSUBS 0.0077f
C405 B.n192 VSUBS 0.0077f
C406 B.n193 VSUBS 0.0077f
C407 B.n194 VSUBS 0.0077f
C408 B.n195 VSUBS 0.0077f
C409 B.n196 VSUBS 0.0077f
C410 B.n197 VSUBS 0.0077f
C411 B.n198 VSUBS 0.0077f
C412 B.n199 VSUBS 0.0077f
C413 B.n200 VSUBS 0.0077f
C414 B.t7 VSUBS 0.050554f
C415 B.t8 VSUBS 0.069053f
C416 B.t6 VSUBS 0.415701f
C417 B.n201 VSUBS 0.122328f
C418 B.n202 VSUBS 0.105317f
C419 B.n203 VSUBS 0.017839f
C420 B.n204 VSUBS 0.006228f
C421 B.n205 VSUBS 0.0077f
C422 B.n206 VSUBS 0.0077f
C423 B.n207 VSUBS 0.0077f
C424 B.n208 VSUBS 0.0077f
C425 B.n209 VSUBS 0.0077f
C426 B.n210 VSUBS 0.0077f
C427 B.n211 VSUBS 0.0077f
C428 B.n212 VSUBS 0.0077f
C429 B.n213 VSUBS 0.0077f
C430 B.n214 VSUBS 0.0077f
C431 B.n215 VSUBS 0.0077f
C432 B.n216 VSUBS 0.0077f
C433 B.n217 VSUBS 0.0077f
C434 B.n218 VSUBS 0.0077f
C435 B.n219 VSUBS 0.0077f
C436 B.n220 VSUBS 0.0077f
C437 B.n221 VSUBS 0.0077f
C438 B.n222 VSUBS 0.0077f
C439 B.n223 VSUBS 0.0077f
C440 B.n224 VSUBS 0.0077f
C441 B.n225 VSUBS 0.0077f
C442 B.n226 VSUBS 0.0077f
C443 B.n227 VSUBS 0.0077f
C444 B.n228 VSUBS 0.017818f
C445 B.n229 VSUBS 0.017818f
C446 B.n230 VSUBS 0.016604f
C447 B.n231 VSUBS 0.0077f
C448 B.n232 VSUBS 0.0077f
C449 B.n233 VSUBS 0.0077f
C450 B.n234 VSUBS 0.0077f
C451 B.n235 VSUBS 0.0077f
C452 B.n236 VSUBS 0.0077f
C453 B.n237 VSUBS 0.0077f
C454 B.n238 VSUBS 0.0077f
C455 B.n239 VSUBS 0.0077f
C456 B.n240 VSUBS 0.0077f
C457 B.n241 VSUBS 0.0077f
C458 B.n242 VSUBS 0.0077f
C459 B.n243 VSUBS 0.0077f
C460 B.n244 VSUBS 0.0077f
C461 B.n245 VSUBS 0.0077f
C462 B.n246 VSUBS 0.0077f
C463 B.n247 VSUBS 0.0077f
C464 B.n248 VSUBS 0.0077f
C465 B.n249 VSUBS 0.0077f
C466 B.n250 VSUBS 0.0077f
C467 B.n251 VSUBS 0.0077f
C468 B.n252 VSUBS 0.0077f
C469 B.n253 VSUBS 0.0077f
C470 B.n254 VSUBS 0.0077f
C471 B.n255 VSUBS 0.0077f
C472 B.n256 VSUBS 0.0077f
C473 B.n257 VSUBS 0.0077f
C474 B.n258 VSUBS 0.0077f
C475 B.n259 VSUBS 0.0077f
C476 B.n260 VSUBS 0.0077f
C477 B.n261 VSUBS 0.0077f
C478 B.n262 VSUBS 0.0077f
C479 B.n263 VSUBS 0.0077f
C480 B.n264 VSUBS 0.0077f
C481 B.n265 VSUBS 0.0077f
C482 B.n266 VSUBS 0.0077f
C483 B.n267 VSUBS 0.0077f
C484 B.n268 VSUBS 0.0077f
C485 B.n269 VSUBS 0.0077f
C486 B.n270 VSUBS 0.0077f
C487 B.n271 VSUBS 0.0077f
C488 B.n272 VSUBS 0.0077f
C489 B.n273 VSUBS 0.0077f
C490 B.n274 VSUBS 0.0077f
C491 B.n275 VSUBS 0.0077f
C492 B.n276 VSUBS 0.0077f
C493 B.n277 VSUBS 0.0077f
C494 B.n278 VSUBS 0.0077f
C495 B.n279 VSUBS 0.0077f
C496 B.n280 VSUBS 0.0077f
C497 B.n281 VSUBS 0.0077f
C498 B.n282 VSUBS 0.0077f
C499 B.n283 VSUBS 0.0077f
C500 B.n284 VSUBS 0.0077f
C501 B.n285 VSUBS 0.0077f
C502 B.n286 VSUBS 0.0077f
C503 B.n287 VSUBS 0.0077f
C504 B.n288 VSUBS 0.0077f
C505 B.n289 VSUBS 0.0077f
C506 B.n290 VSUBS 0.0077f
C507 B.n291 VSUBS 0.0077f
C508 B.n292 VSUBS 0.0077f
C509 B.n293 VSUBS 0.0077f
C510 B.n294 VSUBS 0.0077f
C511 B.n295 VSUBS 0.0077f
C512 B.n296 VSUBS 0.0077f
C513 B.n297 VSUBS 0.0077f
C514 B.n298 VSUBS 0.0077f
C515 B.n299 VSUBS 0.0077f
C516 B.n300 VSUBS 0.0077f
C517 B.n301 VSUBS 0.0077f
C518 B.n302 VSUBS 0.0077f
C519 B.n303 VSUBS 0.0077f
C520 B.n304 VSUBS 0.0077f
C521 B.n305 VSUBS 0.0077f
C522 B.n306 VSUBS 0.0077f
C523 B.n307 VSUBS 0.0077f
C524 B.n308 VSUBS 0.0077f
C525 B.n309 VSUBS 0.0077f
C526 B.n310 VSUBS 0.0077f
C527 B.n311 VSUBS 0.0077f
C528 B.n312 VSUBS 0.0077f
C529 B.n313 VSUBS 0.0077f
C530 B.n314 VSUBS 0.0077f
C531 B.n315 VSUBS 0.0077f
C532 B.n316 VSUBS 0.0077f
C533 B.n317 VSUBS 0.0077f
C534 B.n318 VSUBS 0.0077f
C535 B.n319 VSUBS 0.0077f
C536 B.n320 VSUBS 0.0077f
C537 B.n321 VSUBS 0.0077f
C538 B.n322 VSUBS 0.0077f
C539 B.n323 VSUBS 0.0077f
C540 B.n324 VSUBS 0.0077f
C541 B.n325 VSUBS 0.0077f
C542 B.n326 VSUBS 0.0077f
C543 B.n327 VSUBS 0.0077f
C544 B.n328 VSUBS 0.0077f
C545 B.n329 VSUBS 0.01758f
C546 B.n330 VSUBS 0.016842f
C547 B.n331 VSUBS 0.017818f
C548 B.n332 VSUBS 0.0077f
C549 B.n333 VSUBS 0.0077f
C550 B.n334 VSUBS 0.0077f
C551 B.n335 VSUBS 0.0077f
C552 B.n336 VSUBS 0.0077f
C553 B.n337 VSUBS 0.0077f
C554 B.n338 VSUBS 0.0077f
C555 B.n339 VSUBS 0.0077f
C556 B.n340 VSUBS 0.0077f
C557 B.n341 VSUBS 0.0077f
C558 B.n342 VSUBS 0.0077f
C559 B.n343 VSUBS 0.0077f
C560 B.n344 VSUBS 0.0077f
C561 B.n345 VSUBS 0.0077f
C562 B.n346 VSUBS 0.0077f
C563 B.n347 VSUBS 0.0077f
C564 B.n348 VSUBS 0.0077f
C565 B.n349 VSUBS 0.0077f
C566 B.n350 VSUBS 0.0077f
C567 B.n351 VSUBS 0.0077f
C568 B.n352 VSUBS 0.0077f
C569 B.n353 VSUBS 0.005322f
C570 B.n354 VSUBS 0.017839f
C571 B.n355 VSUBS 0.006228f
C572 B.n356 VSUBS 0.0077f
C573 B.n357 VSUBS 0.0077f
C574 B.n358 VSUBS 0.0077f
C575 B.n359 VSUBS 0.0077f
C576 B.n360 VSUBS 0.0077f
C577 B.n361 VSUBS 0.0077f
C578 B.n362 VSUBS 0.0077f
C579 B.n363 VSUBS 0.0077f
C580 B.n364 VSUBS 0.0077f
C581 B.n365 VSUBS 0.0077f
C582 B.n366 VSUBS 0.0077f
C583 B.n367 VSUBS 0.006228f
C584 B.n368 VSUBS 0.0077f
C585 B.n369 VSUBS 0.0077f
C586 B.n370 VSUBS 0.0077f
C587 B.n371 VSUBS 0.0077f
C588 B.n372 VSUBS 0.0077f
C589 B.n373 VSUBS 0.0077f
C590 B.n374 VSUBS 0.0077f
C591 B.n375 VSUBS 0.0077f
C592 B.n376 VSUBS 0.0077f
C593 B.n377 VSUBS 0.0077f
C594 B.n378 VSUBS 0.0077f
C595 B.n379 VSUBS 0.0077f
C596 B.n380 VSUBS 0.0077f
C597 B.n381 VSUBS 0.0077f
C598 B.n382 VSUBS 0.0077f
C599 B.n383 VSUBS 0.0077f
C600 B.n384 VSUBS 0.0077f
C601 B.n385 VSUBS 0.0077f
C602 B.n386 VSUBS 0.0077f
C603 B.n387 VSUBS 0.0077f
C604 B.n388 VSUBS 0.0077f
C605 B.n389 VSUBS 0.0077f
C606 B.n390 VSUBS 0.0077f
C607 B.n391 VSUBS 0.017818f
C608 B.n392 VSUBS 0.017818f
C609 B.n393 VSUBS 0.016604f
C610 B.n394 VSUBS 0.0077f
C611 B.n395 VSUBS 0.0077f
C612 B.n396 VSUBS 0.0077f
C613 B.n397 VSUBS 0.0077f
C614 B.n398 VSUBS 0.0077f
C615 B.n399 VSUBS 0.0077f
C616 B.n400 VSUBS 0.0077f
C617 B.n401 VSUBS 0.0077f
C618 B.n402 VSUBS 0.0077f
C619 B.n403 VSUBS 0.0077f
C620 B.n404 VSUBS 0.0077f
C621 B.n405 VSUBS 0.0077f
C622 B.n406 VSUBS 0.0077f
C623 B.n407 VSUBS 0.0077f
C624 B.n408 VSUBS 0.0077f
C625 B.n409 VSUBS 0.0077f
C626 B.n410 VSUBS 0.0077f
C627 B.n411 VSUBS 0.0077f
C628 B.n412 VSUBS 0.0077f
C629 B.n413 VSUBS 0.0077f
C630 B.n414 VSUBS 0.0077f
C631 B.n415 VSUBS 0.0077f
C632 B.n416 VSUBS 0.0077f
C633 B.n417 VSUBS 0.0077f
C634 B.n418 VSUBS 0.0077f
C635 B.n419 VSUBS 0.0077f
C636 B.n420 VSUBS 0.0077f
C637 B.n421 VSUBS 0.0077f
C638 B.n422 VSUBS 0.0077f
C639 B.n423 VSUBS 0.0077f
C640 B.n424 VSUBS 0.0077f
C641 B.n425 VSUBS 0.0077f
C642 B.n426 VSUBS 0.0077f
C643 B.n427 VSUBS 0.0077f
C644 B.n428 VSUBS 0.0077f
C645 B.n429 VSUBS 0.0077f
C646 B.n430 VSUBS 0.0077f
C647 B.n431 VSUBS 0.0077f
C648 B.n432 VSUBS 0.0077f
C649 B.n433 VSUBS 0.0077f
C650 B.n434 VSUBS 0.0077f
C651 B.n435 VSUBS 0.0077f
C652 B.n436 VSUBS 0.0077f
C653 B.n437 VSUBS 0.0077f
C654 B.n438 VSUBS 0.0077f
C655 B.n439 VSUBS 0.0077f
C656 B.n440 VSUBS 0.0077f
C657 B.n441 VSUBS 0.0077f
C658 B.n442 VSUBS 0.0077f
C659 B.n443 VSUBS 0.017435f
.ends

