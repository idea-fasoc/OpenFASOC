* NGSPICE file created from diff_pair_sample_0941.ext - technology: sky130A

.subckt diff_pair_sample_0941 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t11 VN.t0 VDD2.t1 B.t5 sky130_fd_pr__nfet_01v8 ad=0.5313 pd=3.55 as=0.5313 ps=3.55 w=3.22 l=2.79
X1 VDD1.t5 VP.t0 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=0.5313 pd=3.55 as=1.2558 ps=7.22 w=3.22 l=2.79
X2 VDD1.t4 VP.t1 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=1.2558 pd=7.22 as=0.5313 ps=3.55 w=3.22 l=2.79
X3 VTAIL.t5 VP.t2 VDD1.t3 B.t5 sky130_fd_pr__nfet_01v8 ad=0.5313 pd=3.55 as=0.5313 ps=3.55 w=3.22 l=2.79
X4 VDD2.t0 VN.t1 VTAIL.t10 B.t0 sky130_fd_pr__nfet_01v8 ad=0.5313 pd=3.55 as=1.2558 ps=7.22 w=3.22 l=2.79
X5 B.t19 B.t17 B.t18 B.t14 sky130_fd_pr__nfet_01v8 ad=1.2558 pd=7.22 as=0 ps=0 w=3.22 l=2.79
X6 VDD2.t4 VN.t2 VTAIL.t9 B.t3 sky130_fd_pr__nfet_01v8 ad=1.2558 pd=7.22 as=0.5313 ps=3.55 w=3.22 l=2.79
X7 VDD1.t2 VP.t3 VTAIL.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=0.5313 pd=3.55 as=1.2558 ps=7.22 w=3.22 l=2.79
X8 B.t16 B.t13 B.t15 B.t14 sky130_fd_pr__nfet_01v8 ad=1.2558 pd=7.22 as=0 ps=0 w=3.22 l=2.79
X9 VTAIL.t8 VN.t3 VDD2.t3 B.t2 sky130_fd_pr__nfet_01v8 ad=0.5313 pd=3.55 as=0.5313 ps=3.55 w=3.22 l=2.79
X10 VDD2.t2 VN.t4 VTAIL.t7 B.t4 sky130_fd_pr__nfet_01v8 ad=0.5313 pd=3.55 as=1.2558 ps=7.22 w=3.22 l=2.79
X11 VDD1.t1 VP.t4 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=1.2558 pd=7.22 as=0.5313 ps=3.55 w=3.22 l=2.79
X12 VTAIL.t2 VP.t5 VDD1.t0 B.t2 sky130_fd_pr__nfet_01v8 ad=0.5313 pd=3.55 as=0.5313 ps=3.55 w=3.22 l=2.79
X13 VDD2.t5 VN.t5 VTAIL.t6 B.t1 sky130_fd_pr__nfet_01v8 ad=1.2558 pd=7.22 as=0.5313 ps=3.55 w=3.22 l=2.79
X14 B.t12 B.t10 B.t11 B.t7 sky130_fd_pr__nfet_01v8 ad=1.2558 pd=7.22 as=0 ps=0 w=3.22 l=2.79
X15 B.t9 B.t6 B.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=1.2558 pd=7.22 as=0 ps=0 w=3.22 l=2.79
R0 VN.n29 VN.n16 161.3
R1 VN.n28 VN.n27 161.3
R2 VN.n26 VN.n17 161.3
R3 VN.n25 VN.n24 161.3
R4 VN.n23 VN.n18 161.3
R5 VN.n22 VN.n21 161.3
R6 VN.n13 VN.n0 161.3
R7 VN.n12 VN.n11 161.3
R8 VN.n10 VN.n1 161.3
R9 VN.n9 VN.n8 161.3
R10 VN.n7 VN.n2 161.3
R11 VN.n6 VN.n5 161.3
R12 VN.n15 VN.n14 104.763
R13 VN.n31 VN.n30 104.763
R14 VN.n4 VN.t5 62.0673
R15 VN.n20 VN.t4 62.0673
R16 VN.n20 VN.n19 48.81
R17 VN.n4 VN.n3 48.81
R18 VN.n8 VN.n1 46.253
R19 VN.n24 VN.n17 46.253
R20 VN VN.n31 43.0511
R21 VN.n8 VN.n7 34.5682
R22 VN.n24 VN.n23 34.5682
R23 VN.n3 VN.t3 27.8148
R24 VN.n14 VN.t1 27.8148
R25 VN.n19 VN.t0 27.8148
R26 VN.n30 VN.t2 27.8148
R27 VN.n6 VN.n3 24.3439
R28 VN.n7 VN.n6 24.3439
R29 VN.n12 VN.n1 24.3439
R30 VN.n13 VN.n12 24.3439
R31 VN.n23 VN.n22 24.3439
R32 VN.n22 VN.n19 24.3439
R33 VN.n29 VN.n28 24.3439
R34 VN.n28 VN.n17 24.3439
R35 VN.n14 VN.n13 5.84292
R36 VN.n30 VN.n29 5.84292
R37 VN.n21 VN.n20 4.95772
R38 VN.n5 VN.n4 4.95772
R39 VN.n31 VN.n16 0.278398
R40 VN.n15 VN.n0 0.278398
R41 VN.n27 VN.n16 0.189894
R42 VN.n27 VN.n26 0.189894
R43 VN.n26 VN.n25 0.189894
R44 VN.n25 VN.n18 0.189894
R45 VN.n21 VN.n18 0.189894
R46 VN.n5 VN.n2 0.189894
R47 VN.n9 VN.n2 0.189894
R48 VN.n10 VN.n9 0.189894
R49 VN.n11 VN.n10 0.189894
R50 VN.n11 VN.n0 0.189894
R51 VN VN.n15 0.153422
R52 VDD2.n27 VDD2.n17 289.615
R53 VDD2.n10 VDD2.n0 289.615
R54 VDD2.n28 VDD2.n27 185
R55 VDD2.n26 VDD2.n25 185
R56 VDD2.n21 VDD2.n20 185
R57 VDD2.n4 VDD2.n3 185
R58 VDD2.n9 VDD2.n8 185
R59 VDD2.n11 VDD2.n10 185
R60 VDD2.n22 VDD2.t4 148.606
R61 VDD2.n5 VDD2.t5 148.606
R62 VDD2.n27 VDD2.n26 104.615
R63 VDD2.n26 VDD2.n20 104.615
R64 VDD2.n9 VDD2.n3 104.615
R65 VDD2.n10 VDD2.n9 104.615
R66 VDD2.n16 VDD2.n15 80.3055
R67 VDD2 VDD2.n33 80.3027
R68 VDD2.n16 VDD2.n14 52.7654
R69 VDD2.t4 VDD2.n20 52.3082
R70 VDD2.t5 VDD2.n3 52.3082
R71 VDD2.n32 VDD2.n31 50.8035
R72 VDD2.n32 VDD2.n16 35.2325
R73 VDD2.n22 VDD2.n21 15.5966
R74 VDD2.n5 VDD2.n4 15.5966
R75 VDD2.n25 VDD2.n24 12.8005
R76 VDD2.n8 VDD2.n7 12.8005
R77 VDD2.n28 VDD2.n19 12.0247
R78 VDD2.n11 VDD2.n2 12.0247
R79 VDD2.n29 VDD2.n17 11.249
R80 VDD2.n12 VDD2.n0 11.249
R81 VDD2.n31 VDD2.n30 9.45567
R82 VDD2.n14 VDD2.n13 9.45567
R83 VDD2.n30 VDD2.n29 9.3005
R84 VDD2.n19 VDD2.n18 9.3005
R85 VDD2.n24 VDD2.n23 9.3005
R86 VDD2.n13 VDD2.n12 9.3005
R87 VDD2.n2 VDD2.n1 9.3005
R88 VDD2.n7 VDD2.n6 9.3005
R89 VDD2.n33 VDD2.t1 6.14957
R90 VDD2.n33 VDD2.t2 6.14957
R91 VDD2.n15 VDD2.t3 6.14957
R92 VDD2.n15 VDD2.t0 6.14957
R93 VDD2.n23 VDD2.n22 4.46457
R94 VDD2.n6 VDD2.n5 4.46457
R95 VDD2.n31 VDD2.n17 2.71565
R96 VDD2.n14 VDD2.n0 2.71565
R97 VDD2 VDD2.n32 2.07593
R98 VDD2.n29 VDD2.n28 1.93989
R99 VDD2.n12 VDD2.n11 1.93989
R100 VDD2.n25 VDD2.n19 1.16414
R101 VDD2.n8 VDD2.n2 1.16414
R102 VDD2.n24 VDD2.n21 0.388379
R103 VDD2.n7 VDD2.n4 0.388379
R104 VDD2.n30 VDD2.n18 0.155672
R105 VDD2.n23 VDD2.n18 0.155672
R106 VDD2.n6 VDD2.n1 0.155672
R107 VDD2.n13 VDD2.n1 0.155672
R108 VTAIL.n66 VTAIL.n56 289.615
R109 VTAIL.n12 VTAIL.n2 289.615
R110 VTAIL.n50 VTAIL.n40 289.615
R111 VTAIL.n32 VTAIL.n22 289.615
R112 VTAIL.n60 VTAIL.n59 185
R113 VTAIL.n65 VTAIL.n64 185
R114 VTAIL.n67 VTAIL.n66 185
R115 VTAIL.n6 VTAIL.n5 185
R116 VTAIL.n11 VTAIL.n10 185
R117 VTAIL.n13 VTAIL.n12 185
R118 VTAIL.n51 VTAIL.n50 185
R119 VTAIL.n49 VTAIL.n48 185
R120 VTAIL.n44 VTAIL.n43 185
R121 VTAIL.n33 VTAIL.n32 185
R122 VTAIL.n31 VTAIL.n30 185
R123 VTAIL.n26 VTAIL.n25 185
R124 VTAIL.n61 VTAIL.t10 148.606
R125 VTAIL.n7 VTAIL.t4 148.606
R126 VTAIL.n45 VTAIL.t0 148.606
R127 VTAIL.n27 VTAIL.t7 148.606
R128 VTAIL.n65 VTAIL.n59 104.615
R129 VTAIL.n66 VTAIL.n65 104.615
R130 VTAIL.n11 VTAIL.n5 104.615
R131 VTAIL.n12 VTAIL.n11 104.615
R132 VTAIL.n50 VTAIL.n49 104.615
R133 VTAIL.n49 VTAIL.n43 104.615
R134 VTAIL.n32 VTAIL.n31 104.615
R135 VTAIL.n31 VTAIL.n25 104.615
R136 VTAIL.n39 VTAIL.n38 63.0098
R137 VTAIL.n21 VTAIL.n20 63.0098
R138 VTAIL.n1 VTAIL.n0 63.0097
R139 VTAIL.n19 VTAIL.n18 63.0097
R140 VTAIL.t10 VTAIL.n59 52.3082
R141 VTAIL.t4 VTAIL.n5 52.3082
R142 VTAIL.t0 VTAIL.n43 52.3082
R143 VTAIL.t7 VTAIL.n25 52.3082
R144 VTAIL.n71 VTAIL.n70 34.1247
R145 VTAIL.n17 VTAIL.n16 34.1247
R146 VTAIL.n55 VTAIL.n54 34.1247
R147 VTAIL.n37 VTAIL.n36 34.1247
R148 VTAIL.n21 VTAIL.n19 20.5221
R149 VTAIL.n71 VTAIL.n55 17.8324
R150 VTAIL.n61 VTAIL.n60 15.5966
R151 VTAIL.n7 VTAIL.n6 15.5966
R152 VTAIL.n45 VTAIL.n44 15.5966
R153 VTAIL.n27 VTAIL.n26 15.5966
R154 VTAIL.n64 VTAIL.n63 12.8005
R155 VTAIL.n10 VTAIL.n9 12.8005
R156 VTAIL.n48 VTAIL.n47 12.8005
R157 VTAIL.n30 VTAIL.n29 12.8005
R158 VTAIL.n67 VTAIL.n58 12.0247
R159 VTAIL.n13 VTAIL.n4 12.0247
R160 VTAIL.n51 VTAIL.n42 12.0247
R161 VTAIL.n33 VTAIL.n24 12.0247
R162 VTAIL.n68 VTAIL.n56 11.249
R163 VTAIL.n14 VTAIL.n2 11.249
R164 VTAIL.n52 VTAIL.n40 11.249
R165 VTAIL.n34 VTAIL.n22 11.249
R166 VTAIL.n70 VTAIL.n69 9.45567
R167 VTAIL.n16 VTAIL.n15 9.45567
R168 VTAIL.n54 VTAIL.n53 9.45567
R169 VTAIL.n36 VTAIL.n35 9.45567
R170 VTAIL.n69 VTAIL.n68 9.3005
R171 VTAIL.n58 VTAIL.n57 9.3005
R172 VTAIL.n63 VTAIL.n62 9.3005
R173 VTAIL.n15 VTAIL.n14 9.3005
R174 VTAIL.n4 VTAIL.n3 9.3005
R175 VTAIL.n9 VTAIL.n8 9.3005
R176 VTAIL.n53 VTAIL.n52 9.3005
R177 VTAIL.n42 VTAIL.n41 9.3005
R178 VTAIL.n47 VTAIL.n46 9.3005
R179 VTAIL.n35 VTAIL.n34 9.3005
R180 VTAIL.n24 VTAIL.n23 9.3005
R181 VTAIL.n29 VTAIL.n28 9.3005
R182 VTAIL.n0 VTAIL.t6 6.14957
R183 VTAIL.n0 VTAIL.t8 6.14957
R184 VTAIL.n18 VTAIL.t3 6.14957
R185 VTAIL.n18 VTAIL.t5 6.14957
R186 VTAIL.n38 VTAIL.t1 6.14957
R187 VTAIL.n38 VTAIL.t2 6.14957
R188 VTAIL.n20 VTAIL.t9 6.14957
R189 VTAIL.n20 VTAIL.t11 6.14957
R190 VTAIL.n62 VTAIL.n61 4.46457
R191 VTAIL.n8 VTAIL.n7 4.46457
R192 VTAIL.n46 VTAIL.n45 4.46457
R193 VTAIL.n28 VTAIL.n27 4.46457
R194 VTAIL.n70 VTAIL.n56 2.71565
R195 VTAIL.n16 VTAIL.n2 2.71565
R196 VTAIL.n54 VTAIL.n40 2.71565
R197 VTAIL.n36 VTAIL.n22 2.71565
R198 VTAIL.n37 VTAIL.n21 2.69016
R199 VTAIL.n55 VTAIL.n39 2.69016
R200 VTAIL.n19 VTAIL.n17 2.69016
R201 VTAIL VTAIL.n71 1.95955
R202 VTAIL.n68 VTAIL.n67 1.93989
R203 VTAIL.n14 VTAIL.n13 1.93989
R204 VTAIL.n52 VTAIL.n51 1.93989
R205 VTAIL.n34 VTAIL.n33 1.93989
R206 VTAIL.n39 VTAIL.n37 1.81516
R207 VTAIL.n17 VTAIL.n1 1.81516
R208 VTAIL.n64 VTAIL.n58 1.16414
R209 VTAIL.n10 VTAIL.n4 1.16414
R210 VTAIL.n48 VTAIL.n42 1.16414
R211 VTAIL.n30 VTAIL.n24 1.16414
R212 VTAIL VTAIL.n1 0.731103
R213 VTAIL.n63 VTAIL.n60 0.388379
R214 VTAIL.n9 VTAIL.n6 0.388379
R215 VTAIL.n47 VTAIL.n44 0.388379
R216 VTAIL.n29 VTAIL.n26 0.388379
R217 VTAIL.n62 VTAIL.n57 0.155672
R218 VTAIL.n69 VTAIL.n57 0.155672
R219 VTAIL.n8 VTAIL.n3 0.155672
R220 VTAIL.n15 VTAIL.n3 0.155672
R221 VTAIL.n53 VTAIL.n41 0.155672
R222 VTAIL.n46 VTAIL.n41 0.155672
R223 VTAIL.n35 VTAIL.n23 0.155672
R224 VTAIL.n28 VTAIL.n23 0.155672
R225 B.n579 B.n578 585
R226 B.n580 B.n579 585
R227 B.n189 B.n104 585
R228 B.n188 B.n187 585
R229 B.n186 B.n185 585
R230 B.n184 B.n183 585
R231 B.n182 B.n181 585
R232 B.n180 B.n179 585
R233 B.n178 B.n177 585
R234 B.n176 B.n175 585
R235 B.n174 B.n173 585
R236 B.n172 B.n171 585
R237 B.n170 B.n169 585
R238 B.n168 B.n167 585
R239 B.n166 B.n165 585
R240 B.n164 B.n163 585
R241 B.n162 B.n161 585
R242 B.n159 B.n158 585
R243 B.n157 B.n156 585
R244 B.n155 B.n154 585
R245 B.n153 B.n152 585
R246 B.n151 B.n150 585
R247 B.n149 B.n148 585
R248 B.n147 B.n146 585
R249 B.n145 B.n144 585
R250 B.n143 B.n142 585
R251 B.n141 B.n140 585
R252 B.n139 B.n138 585
R253 B.n137 B.n136 585
R254 B.n135 B.n134 585
R255 B.n133 B.n132 585
R256 B.n131 B.n130 585
R257 B.n129 B.n128 585
R258 B.n127 B.n126 585
R259 B.n125 B.n124 585
R260 B.n123 B.n122 585
R261 B.n121 B.n120 585
R262 B.n119 B.n118 585
R263 B.n117 B.n116 585
R264 B.n115 B.n114 585
R265 B.n113 B.n112 585
R266 B.n111 B.n110 585
R267 B.n577 B.n83 585
R268 B.n581 B.n83 585
R269 B.n576 B.n82 585
R270 B.n582 B.n82 585
R271 B.n575 B.n574 585
R272 B.n574 B.n78 585
R273 B.n573 B.n77 585
R274 B.n588 B.n77 585
R275 B.n572 B.n76 585
R276 B.n589 B.n76 585
R277 B.n571 B.n75 585
R278 B.n590 B.n75 585
R279 B.n570 B.n569 585
R280 B.n569 B.n71 585
R281 B.n568 B.n70 585
R282 B.n596 B.n70 585
R283 B.n567 B.n69 585
R284 B.n597 B.n69 585
R285 B.n566 B.n68 585
R286 B.n598 B.n68 585
R287 B.n565 B.n564 585
R288 B.n564 B.n64 585
R289 B.n563 B.n63 585
R290 B.n604 B.n63 585
R291 B.n562 B.n62 585
R292 B.n605 B.n62 585
R293 B.n561 B.n61 585
R294 B.n606 B.n61 585
R295 B.n560 B.n559 585
R296 B.n559 B.n57 585
R297 B.n558 B.n56 585
R298 B.n612 B.n56 585
R299 B.n557 B.n55 585
R300 B.n613 B.n55 585
R301 B.n556 B.n54 585
R302 B.n614 B.n54 585
R303 B.n555 B.n554 585
R304 B.n554 B.n50 585
R305 B.n553 B.n49 585
R306 B.n620 B.n49 585
R307 B.n552 B.n48 585
R308 B.n621 B.n48 585
R309 B.n551 B.n47 585
R310 B.n622 B.n47 585
R311 B.n550 B.n549 585
R312 B.n549 B.n43 585
R313 B.n548 B.n42 585
R314 B.n628 B.n42 585
R315 B.n547 B.n41 585
R316 B.n629 B.n41 585
R317 B.n546 B.n40 585
R318 B.n630 B.n40 585
R319 B.n545 B.n544 585
R320 B.n544 B.n36 585
R321 B.n543 B.n35 585
R322 B.n636 B.n35 585
R323 B.n542 B.n34 585
R324 B.n637 B.n34 585
R325 B.n541 B.n33 585
R326 B.n638 B.n33 585
R327 B.n540 B.n539 585
R328 B.n539 B.n29 585
R329 B.n538 B.n28 585
R330 B.n644 B.n28 585
R331 B.n537 B.n27 585
R332 B.n645 B.n27 585
R333 B.n536 B.n26 585
R334 B.n646 B.n26 585
R335 B.n535 B.n534 585
R336 B.n534 B.n22 585
R337 B.n533 B.n21 585
R338 B.n652 B.n21 585
R339 B.n532 B.n20 585
R340 B.n653 B.n20 585
R341 B.n531 B.n19 585
R342 B.n654 B.n19 585
R343 B.n530 B.n529 585
R344 B.n529 B.n18 585
R345 B.n528 B.n14 585
R346 B.n660 B.n14 585
R347 B.n527 B.n13 585
R348 B.n661 B.n13 585
R349 B.n526 B.n12 585
R350 B.n662 B.n12 585
R351 B.n525 B.n524 585
R352 B.n524 B.n8 585
R353 B.n523 B.n7 585
R354 B.n668 B.n7 585
R355 B.n522 B.n6 585
R356 B.n669 B.n6 585
R357 B.n521 B.n5 585
R358 B.n670 B.n5 585
R359 B.n520 B.n519 585
R360 B.n519 B.n4 585
R361 B.n518 B.n190 585
R362 B.n518 B.n517 585
R363 B.n508 B.n191 585
R364 B.n192 B.n191 585
R365 B.n510 B.n509 585
R366 B.n511 B.n510 585
R367 B.n507 B.n197 585
R368 B.n197 B.n196 585
R369 B.n506 B.n505 585
R370 B.n505 B.n504 585
R371 B.n199 B.n198 585
R372 B.n497 B.n199 585
R373 B.n496 B.n495 585
R374 B.n498 B.n496 585
R375 B.n494 B.n204 585
R376 B.n204 B.n203 585
R377 B.n493 B.n492 585
R378 B.n492 B.n491 585
R379 B.n206 B.n205 585
R380 B.n207 B.n206 585
R381 B.n484 B.n483 585
R382 B.n485 B.n484 585
R383 B.n482 B.n212 585
R384 B.n212 B.n211 585
R385 B.n481 B.n480 585
R386 B.n480 B.n479 585
R387 B.n214 B.n213 585
R388 B.n215 B.n214 585
R389 B.n472 B.n471 585
R390 B.n473 B.n472 585
R391 B.n470 B.n220 585
R392 B.n220 B.n219 585
R393 B.n469 B.n468 585
R394 B.n468 B.n467 585
R395 B.n222 B.n221 585
R396 B.n223 B.n222 585
R397 B.n460 B.n459 585
R398 B.n461 B.n460 585
R399 B.n458 B.n228 585
R400 B.n228 B.n227 585
R401 B.n457 B.n456 585
R402 B.n456 B.n455 585
R403 B.n230 B.n229 585
R404 B.n231 B.n230 585
R405 B.n448 B.n447 585
R406 B.n449 B.n448 585
R407 B.n446 B.n235 585
R408 B.n239 B.n235 585
R409 B.n445 B.n444 585
R410 B.n444 B.n443 585
R411 B.n237 B.n236 585
R412 B.n238 B.n237 585
R413 B.n436 B.n435 585
R414 B.n437 B.n436 585
R415 B.n434 B.n244 585
R416 B.n244 B.n243 585
R417 B.n433 B.n432 585
R418 B.n432 B.n431 585
R419 B.n246 B.n245 585
R420 B.n247 B.n246 585
R421 B.n424 B.n423 585
R422 B.n425 B.n424 585
R423 B.n422 B.n252 585
R424 B.n252 B.n251 585
R425 B.n421 B.n420 585
R426 B.n420 B.n419 585
R427 B.n254 B.n253 585
R428 B.n255 B.n254 585
R429 B.n412 B.n411 585
R430 B.n413 B.n412 585
R431 B.n410 B.n259 585
R432 B.n263 B.n259 585
R433 B.n409 B.n408 585
R434 B.n408 B.n407 585
R435 B.n261 B.n260 585
R436 B.n262 B.n261 585
R437 B.n400 B.n399 585
R438 B.n401 B.n400 585
R439 B.n398 B.n268 585
R440 B.n268 B.n267 585
R441 B.n397 B.n396 585
R442 B.n396 B.n395 585
R443 B.n270 B.n269 585
R444 B.n271 B.n270 585
R445 B.n388 B.n387 585
R446 B.n389 B.n388 585
R447 B.n386 B.n276 585
R448 B.n276 B.n275 585
R449 B.n380 B.n379 585
R450 B.n378 B.n298 585
R451 B.n377 B.n297 585
R452 B.n382 B.n297 585
R453 B.n376 B.n375 585
R454 B.n374 B.n373 585
R455 B.n372 B.n371 585
R456 B.n370 B.n369 585
R457 B.n368 B.n367 585
R458 B.n366 B.n365 585
R459 B.n364 B.n363 585
R460 B.n362 B.n361 585
R461 B.n360 B.n359 585
R462 B.n358 B.n357 585
R463 B.n356 B.n355 585
R464 B.n354 B.n353 585
R465 B.n352 B.n351 585
R466 B.n349 B.n348 585
R467 B.n347 B.n346 585
R468 B.n345 B.n344 585
R469 B.n343 B.n342 585
R470 B.n341 B.n340 585
R471 B.n339 B.n338 585
R472 B.n337 B.n336 585
R473 B.n335 B.n334 585
R474 B.n333 B.n332 585
R475 B.n331 B.n330 585
R476 B.n329 B.n328 585
R477 B.n327 B.n326 585
R478 B.n325 B.n324 585
R479 B.n323 B.n322 585
R480 B.n321 B.n320 585
R481 B.n319 B.n318 585
R482 B.n317 B.n316 585
R483 B.n315 B.n314 585
R484 B.n313 B.n312 585
R485 B.n311 B.n310 585
R486 B.n309 B.n308 585
R487 B.n307 B.n306 585
R488 B.n305 B.n304 585
R489 B.n278 B.n277 585
R490 B.n385 B.n384 585
R491 B.n274 B.n273 585
R492 B.n275 B.n274 585
R493 B.n391 B.n390 585
R494 B.n390 B.n389 585
R495 B.n392 B.n272 585
R496 B.n272 B.n271 585
R497 B.n394 B.n393 585
R498 B.n395 B.n394 585
R499 B.n266 B.n265 585
R500 B.n267 B.n266 585
R501 B.n403 B.n402 585
R502 B.n402 B.n401 585
R503 B.n404 B.n264 585
R504 B.n264 B.n262 585
R505 B.n406 B.n405 585
R506 B.n407 B.n406 585
R507 B.n258 B.n257 585
R508 B.n263 B.n258 585
R509 B.n415 B.n414 585
R510 B.n414 B.n413 585
R511 B.n416 B.n256 585
R512 B.n256 B.n255 585
R513 B.n418 B.n417 585
R514 B.n419 B.n418 585
R515 B.n250 B.n249 585
R516 B.n251 B.n250 585
R517 B.n427 B.n426 585
R518 B.n426 B.n425 585
R519 B.n428 B.n248 585
R520 B.n248 B.n247 585
R521 B.n430 B.n429 585
R522 B.n431 B.n430 585
R523 B.n242 B.n241 585
R524 B.n243 B.n242 585
R525 B.n439 B.n438 585
R526 B.n438 B.n437 585
R527 B.n440 B.n240 585
R528 B.n240 B.n238 585
R529 B.n442 B.n441 585
R530 B.n443 B.n442 585
R531 B.n234 B.n233 585
R532 B.n239 B.n234 585
R533 B.n451 B.n450 585
R534 B.n450 B.n449 585
R535 B.n452 B.n232 585
R536 B.n232 B.n231 585
R537 B.n454 B.n453 585
R538 B.n455 B.n454 585
R539 B.n226 B.n225 585
R540 B.n227 B.n226 585
R541 B.n463 B.n462 585
R542 B.n462 B.n461 585
R543 B.n464 B.n224 585
R544 B.n224 B.n223 585
R545 B.n466 B.n465 585
R546 B.n467 B.n466 585
R547 B.n218 B.n217 585
R548 B.n219 B.n218 585
R549 B.n475 B.n474 585
R550 B.n474 B.n473 585
R551 B.n476 B.n216 585
R552 B.n216 B.n215 585
R553 B.n478 B.n477 585
R554 B.n479 B.n478 585
R555 B.n210 B.n209 585
R556 B.n211 B.n210 585
R557 B.n487 B.n486 585
R558 B.n486 B.n485 585
R559 B.n488 B.n208 585
R560 B.n208 B.n207 585
R561 B.n490 B.n489 585
R562 B.n491 B.n490 585
R563 B.n202 B.n201 585
R564 B.n203 B.n202 585
R565 B.n500 B.n499 585
R566 B.n499 B.n498 585
R567 B.n501 B.n200 585
R568 B.n497 B.n200 585
R569 B.n503 B.n502 585
R570 B.n504 B.n503 585
R571 B.n195 B.n194 585
R572 B.n196 B.n195 585
R573 B.n513 B.n512 585
R574 B.n512 B.n511 585
R575 B.n514 B.n193 585
R576 B.n193 B.n192 585
R577 B.n516 B.n515 585
R578 B.n517 B.n516 585
R579 B.n2 B.n0 585
R580 B.n4 B.n2 585
R581 B.n3 B.n1 585
R582 B.n669 B.n3 585
R583 B.n667 B.n666 585
R584 B.n668 B.n667 585
R585 B.n665 B.n9 585
R586 B.n9 B.n8 585
R587 B.n664 B.n663 585
R588 B.n663 B.n662 585
R589 B.n11 B.n10 585
R590 B.n661 B.n11 585
R591 B.n659 B.n658 585
R592 B.n660 B.n659 585
R593 B.n657 B.n15 585
R594 B.n18 B.n15 585
R595 B.n656 B.n655 585
R596 B.n655 B.n654 585
R597 B.n17 B.n16 585
R598 B.n653 B.n17 585
R599 B.n651 B.n650 585
R600 B.n652 B.n651 585
R601 B.n649 B.n23 585
R602 B.n23 B.n22 585
R603 B.n648 B.n647 585
R604 B.n647 B.n646 585
R605 B.n25 B.n24 585
R606 B.n645 B.n25 585
R607 B.n643 B.n642 585
R608 B.n644 B.n643 585
R609 B.n641 B.n30 585
R610 B.n30 B.n29 585
R611 B.n640 B.n639 585
R612 B.n639 B.n638 585
R613 B.n32 B.n31 585
R614 B.n637 B.n32 585
R615 B.n635 B.n634 585
R616 B.n636 B.n635 585
R617 B.n633 B.n37 585
R618 B.n37 B.n36 585
R619 B.n632 B.n631 585
R620 B.n631 B.n630 585
R621 B.n39 B.n38 585
R622 B.n629 B.n39 585
R623 B.n627 B.n626 585
R624 B.n628 B.n627 585
R625 B.n625 B.n44 585
R626 B.n44 B.n43 585
R627 B.n624 B.n623 585
R628 B.n623 B.n622 585
R629 B.n46 B.n45 585
R630 B.n621 B.n46 585
R631 B.n619 B.n618 585
R632 B.n620 B.n619 585
R633 B.n617 B.n51 585
R634 B.n51 B.n50 585
R635 B.n616 B.n615 585
R636 B.n615 B.n614 585
R637 B.n53 B.n52 585
R638 B.n613 B.n53 585
R639 B.n611 B.n610 585
R640 B.n612 B.n611 585
R641 B.n609 B.n58 585
R642 B.n58 B.n57 585
R643 B.n608 B.n607 585
R644 B.n607 B.n606 585
R645 B.n60 B.n59 585
R646 B.n605 B.n60 585
R647 B.n603 B.n602 585
R648 B.n604 B.n603 585
R649 B.n601 B.n65 585
R650 B.n65 B.n64 585
R651 B.n600 B.n599 585
R652 B.n599 B.n598 585
R653 B.n67 B.n66 585
R654 B.n597 B.n67 585
R655 B.n595 B.n594 585
R656 B.n596 B.n595 585
R657 B.n593 B.n72 585
R658 B.n72 B.n71 585
R659 B.n592 B.n591 585
R660 B.n591 B.n590 585
R661 B.n74 B.n73 585
R662 B.n589 B.n74 585
R663 B.n587 B.n586 585
R664 B.n588 B.n587 585
R665 B.n585 B.n79 585
R666 B.n79 B.n78 585
R667 B.n584 B.n583 585
R668 B.n583 B.n582 585
R669 B.n81 B.n80 585
R670 B.n581 B.n81 585
R671 B.n672 B.n671 585
R672 B.n671 B.n670 585
R673 B.n380 B.n274 482.89
R674 B.n110 B.n81 482.89
R675 B.n384 B.n276 482.89
R676 B.n579 B.n83 482.89
R677 B.n580 B.n103 256.663
R678 B.n580 B.n102 256.663
R679 B.n580 B.n101 256.663
R680 B.n580 B.n100 256.663
R681 B.n580 B.n99 256.663
R682 B.n580 B.n98 256.663
R683 B.n580 B.n97 256.663
R684 B.n580 B.n96 256.663
R685 B.n580 B.n95 256.663
R686 B.n580 B.n94 256.663
R687 B.n580 B.n93 256.663
R688 B.n580 B.n92 256.663
R689 B.n580 B.n91 256.663
R690 B.n580 B.n90 256.663
R691 B.n580 B.n89 256.663
R692 B.n580 B.n88 256.663
R693 B.n580 B.n87 256.663
R694 B.n580 B.n86 256.663
R695 B.n580 B.n85 256.663
R696 B.n580 B.n84 256.663
R697 B.n382 B.n381 256.663
R698 B.n382 B.n279 256.663
R699 B.n382 B.n280 256.663
R700 B.n382 B.n281 256.663
R701 B.n382 B.n282 256.663
R702 B.n382 B.n283 256.663
R703 B.n382 B.n284 256.663
R704 B.n382 B.n285 256.663
R705 B.n382 B.n286 256.663
R706 B.n382 B.n287 256.663
R707 B.n382 B.n288 256.663
R708 B.n382 B.n289 256.663
R709 B.n382 B.n290 256.663
R710 B.n382 B.n291 256.663
R711 B.n382 B.n292 256.663
R712 B.n382 B.n293 256.663
R713 B.n382 B.n294 256.663
R714 B.n382 B.n295 256.663
R715 B.n382 B.n296 256.663
R716 B.n383 B.n382 256.663
R717 B.n301 B.t13 236.131
R718 B.n299 B.t17 236.131
R719 B.n107 B.t10 236.131
R720 B.n105 B.t6 236.131
R721 B.n301 B.t16 193.077
R722 B.n105 B.t8 193.077
R723 B.n299 B.t19 193.077
R724 B.n107 B.t11 193.077
R725 B.n390 B.n274 163.367
R726 B.n390 B.n272 163.367
R727 B.n394 B.n272 163.367
R728 B.n394 B.n266 163.367
R729 B.n402 B.n266 163.367
R730 B.n402 B.n264 163.367
R731 B.n406 B.n264 163.367
R732 B.n406 B.n258 163.367
R733 B.n414 B.n258 163.367
R734 B.n414 B.n256 163.367
R735 B.n418 B.n256 163.367
R736 B.n418 B.n250 163.367
R737 B.n426 B.n250 163.367
R738 B.n426 B.n248 163.367
R739 B.n430 B.n248 163.367
R740 B.n430 B.n242 163.367
R741 B.n438 B.n242 163.367
R742 B.n438 B.n240 163.367
R743 B.n442 B.n240 163.367
R744 B.n442 B.n234 163.367
R745 B.n450 B.n234 163.367
R746 B.n450 B.n232 163.367
R747 B.n454 B.n232 163.367
R748 B.n454 B.n226 163.367
R749 B.n462 B.n226 163.367
R750 B.n462 B.n224 163.367
R751 B.n466 B.n224 163.367
R752 B.n466 B.n218 163.367
R753 B.n474 B.n218 163.367
R754 B.n474 B.n216 163.367
R755 B.n478 B.n216 163.367
R756 B.n478 B.n210 163.367
R757 B.n486 B.n210 163.367
R758 B.n486 B.n208 163.367
R759 B.n490 B.n208 163.367
R760 B.n490 B.n202 163.367
R761 B.n499 B.n202 163.367
R762 B.n499 B.n200 163.367
R763 B.n503 B.n200 163.367
R764 B.n503 B.n195 163.367
R765 B.n512 B.n195 163.367
R766 B.n512 B.n193 163.367
R767 B.n516 B.n193 163.367
R768 B.n516 B.n2 163.367
R769 B.n671 B.n2 163.367
R770 B.n671 B.n3 163.367
R771 B.n667 B.n3 163.367
R772 B.n667 B.n9 163.367
R773 B.n663 B.n9 163.367
R774 B.n663 B.n11 163.367
R775 B.n659 B.n11 163.367
R776 B.n659 B.n15 163.367
R777 B.n655 B.n15 163.367
R778 B.n655 B.n17 163.367
R779 B.n651 B.n17 163.367
R780 B.n651 B.n23 163.367
R781 B.n647 B.n23 163.367
R782 B.n647 B.n25 163.367
R783 B.n643 B.n25 163.367
R784 B.n643 B.n30 163.367
R785 B.n639 B.n30 163.367
R786 B.n639 B.n32 163.367
R787 B.n635 B.n32 163.367
R788 B.n635 B.n37 163.367
R789 B.n631 B.n37 163.367
R790 B.n631 B.n39 163.367
R791 B.n627 B.n39 163.367
R792 B.n627 B.n44 163.367
R793 B.n623 B.n44 163.367
R794 B.n623 B.n46 163.367
R795 B.n619 B.n46 163.367
R796 B.n619 B.n51 163.367
R797 B.n615 B.n51 163.367
R798 B.n615 B.n53 163.367
R799 B.n611 B.n53 163.367
R800 B.n611 B.n58 163.367
R801 B.n607 B.n58 163.367
R802 B.n607 B.n60 163.367
R803 B.n603 B.n60 163.367
R804 B.n603 B.n65 163.367
R805 B.n599 B.n65 163.367
R806 B.n599 B.n67 163.367
R807 B.n595 B.n67 163.367
R808 B.n595 B.n72 163.367
R809 B.n591 B.n72 163.367
R810 B.n591 B.n74 163.367
R811 B.n587 B.n74 163.367
R812 B.n587 B.n79 163.367
R813 B.n583 B.n79 163.367
R814 B.n583 B.n81 163.367
R815 B.n298 B.n297 163.367
R816 B.n375 B.n297 163.367
R817 B.n373 B.n372 163.367
R818 B.n369 B.n368 163.367
R819 B.n365 B.n364 163.367
R820 B.n361 B.n360 163.367
R821 B.n357 B.n356 163.367
R822 B.n353 B.n352 163.367
R823 B.n348 B.n347 163.367
R824 B.n344 B.n343 163.367
R825 B.n340 B.n339 163.367
R826 B.n336 B.n335 163.367
R827 B.n332 B.n331 163.367
R828 B.n328 B.n327 163.367
R829 B.n324 B.n323 163.367
R830 B.n320 B.n319 163.367
R831 B.n316 B.n315 163.367
R832 B.n312 B.n311 163.367
R833 B.n308 B.n307 163.367
R834 B.n304 B.n278 163.367
R835 B.n388 B.n276 163.367
R836 B.n388 B.n270 163.367
R837 B.n396 B.n270 163.367
R838 B.n396 B.n268 163.367
R839 B.n400 B.n268 163.367
R840 B.n400 B.n261 163.367
R841 B.n408 B.n261 163.367
R842 B.n408 B.n259 163.367
R843 B.n412 B.n259 163.367
R844 B.n412 B.n254 163.367
R845 B.n420 B.n254 163.367
R846 B.n420 B.n252 163.367
R847 B.n424 B.n252 163.367
R848 B.n424 B.n246 163.367
R849 B.n432 B.n246 163.367
R850 B.n432 B.n244 163.367
R851 B.n436 B.n244 163.367
R852 B.n436 B.n237 163.367
R853 B.n444 B.n237 163.367
R854 B.n444 B.n235 163.367
R855 B.n448 B.n235 163.367
R856 B.n448 B.n230 163.367
R857 B.n456 B.n230 163.367
R858 B.n456 B.n228 163.367
R859 B.n460 B.n228 163.367
R860 B.n460 B.n222 163.367
R861 B.n468 B.n222 163.367
R862 B.n468 B.n220 163.367
R863 B.n472 B.n220 163.367
R864 B.n472 B.n214 163.367
R865 B.n480 B.n214 163.367
R866 B.n480 B.n212 163.367
R867 B.n484 B.n212 163.367
R868 B.n484 B.n206 163.367
R869 B.n492 B.n206 163.367
R870 B.n492 B.n204 163.367
R871 B.n496 B.n204 163.367
R872 B.n496 B.n199 163.367
R873 B.n505 B.n199 163.367
R874 B.n505 B.n197 163.367
R875 B.n510 B.n197 163.367
R876 B.n510 B.n191 163.367
R877 B.n518 B.n191 163.367
R878 B.n519 B.n518 163.367
R879 B.n519 B.n5 163.367
R880 B.n6 B.n5 163.367
R881 B.n7 B.n6 163.367
R882 B.n524 B.n7 163.367
R883 B.n524 B.n12 163.367
R884 B.n13 B.n12 163.367
R885 B.n14 B.n13 163.367
R886 B.n529 B.n14 163.367
R887 B.n529 B.n19 163.367
R888 B.n20 B.n19 163.367
R889 B.n21 B.n20 163.367
R890 B.n534 B.n21 163.367
R891 B.n534 B.n26 163.367
R892 B.n27 B.n26 163.367
R893 B.n28 B.n27 163.367
R894 B.n539 B.n28 163.367
R895 B.n539 B.n33 163.367
R896 B.n34 B.n33 163.367
R897 B.n35 B.n34 163.367
R898 B.n544 B.n35 163.367
R899 B.n544 B.n40 163.367
R900 B.n41 B.n40 163.367
R901 B.n42 B.n41 163.367
R902 B.n549 B.n42 163.367
R903 B.n549 B.n47 163.367
R904 B.n48 B.n47 163.367
R905 B.n49 B.n48 163.367
R906 B.n554 B.n49 163.367
R907 B.n554 B.n54 163.367
R908 B.n55 B.n54 163.367
R909 B.n56 B.n55 163.367
R910 B.n559 B.n56 163.367
R911 B.n559 B.n61 163.367
R912 B.n62 B.n61 163.367
R913 B.n63 B.n62 163.367
R914 B.n564 B.n63 163.367
R915 B.n564 B.n68 163.367
R916 B.n69 B.n68 163.367
R917 B.n70 B.n69 163.367
R918 B.n569 B.n70 163.367
R919 B.n569 B.n75 163.367
R920 B.n76 B.n75 163.367
R921 B.n77 B.n76 163.367
R922 B.n574 B.n77 163.367
R923 B.n574 B.n82 163.367
R924 B.n83 B.n82 163.367
R925 B.n114 B.n113 163.367
R926 B.n118 B.n117 163.367
R927 B.n122 B.n121 163.367
R928 B.n126 B.n125 163.367
R929 B.n130 B.n129 163.367
R930 B.n134 B.n133 163.367
R931 B.n138 B.n137 163.367
R932 B.n142 B.n141 163.367
R933 B.n146 B.n145 163.367
R934 B.n150 B.n149 163.367
R935 B.n154 B.n153 163.367
R936 B.n158 B.n157 163.367
R937 B.n163 B.n162 163.367
R938 B.n167 B.n166 163.367
R939 B.n171 B.n170 163.367
R940 B.n175 B.n174 163.367
R941 B.n179 B.n178 163.367
R942 B.n183 B.n182 163.367
R943 B.n187 B.n186 163.367
R944 B.n579 B.n104 163.367
R945 B.n382 B.n275 143.732
R946 B.n581 B.n580 143.732
R947 B.n302 B.t15 132.567
R948 B.n106 B.t9 132.567
R949 B.n300 B.t18 132.567
R950 B.n108 B.t12 132.567
R951 B.n389 B.n275 88.0523
R952 B.n389 B.n271 88.0523
R953 B.n395 B.n271 88.0523
R954 B.n395 B.n267 88.0523
R955 B.n401 B.n267 88.0523
R956 B.n401 B.n262 88.0523
R957 B.n407 B.n262 88.0523
R958 B.n407 B.n263 88.0523
R959 B.n413 B.n255 88.0523
R960 B.n419 B.n255 88.0523
R961 B.n419 B.n251 88.0523
R962 B.n425 B.n251 88.0523
R963 B.n425 B.n247 88.0523
R964 B.n431 B.n247 88.0523
R965 B.n431 B.n243 88.0523
R966 B.n437 B.n243 88.0523
R967 B.n437 B.n238 88.0523
R968 B.n443 B.n238 88.0523
R969 B.n443 B.n239 88.0523
R970 B.n449 B.n231 88.0523
R971 B.n455 B.n231 88.0523
R972 B.n455 B.n227 88.0523
R973 B.n461 B.n227 88.0523
R974 B.n461 B.n223 88.0523
R975 B.n467 B.n223 88.0523
R976 B.n467 B.n219 88.0523
R977 B.n473 B.n219 88.0523
R978 B.n479 B.n215 88.0523
R979 B.n479 B.n211 88.0523
R980 B.n485 B.n211 88.0523
R981 B.n485 B.n207 88.0523
R982 B.n491 B.n207 88.0523
R983 B.n491 B.n203 88.0523
R984 B.n498 B.n203 88.0523
R985 B.n498 B.n497 88.0523
R986 B.n504 B.n196 88.0523
R987 B.n511 B.n196 88.0523
R988 B.n511 B.n192 88.0523
R989 B.n517 B.n192 88.0523
R990 B.n517 B.n4 88.0523
R991 B.n670 B.n4 88.0523
R992 B.n670 B.n669 88.0523
R993 B.n669 B.n668 88.0523
R994 B.n668 B.n8 88.0523
R995 B.n662 B.n8 88.0523
R996 B.n662 B.n661 88.0523
R997 B.n661 B.n660 88.0523
R998 B.n654 B.n18 88.0523
R999 B.n654 B.n653 88.0523
R1000 B.n653 B.n652 88.0523
R1001 B.n652 B.n22 88.0523
R1002 B.n646 B.n22 88.0523
R1003 B.n646 B.n645 88.0523
R1004 B.n645 B.n644 88.0523
R1005 B.n644 B.n29 88.0523
R1006 B.n638 B.n637 88.0523
R1007 B.n637 B.n636 88.0523
R1008 B.n636 B.n36 88.0523
R1009 B.n630 B.n36 88.0523
R1010 B.n630 B.n629 88.0523
R1011 B.n629 B.n628 88.0523
R1012 B.n628 B.n43 88.0523
R1013 B.n622 B.n43 88.0523
R1014 B.n621 B.n620 88.0523
R1015 B.n620 B.n50 88.0523
R1016 B.n614 B.n50 88.0523
R1017 B.n614 B.n613 88.0523
R1018 B.n613 B.n612 88.0523
R1019 B.n612 B.n57 88.0523
R1020 B.n606 B.n57 88.0523
R1021 B.n606 B.n605 88.0523
R1022 B.n605 B.n604 88.0523
R1023 B.n604 B.n64 88.0523
R1024 B.n598 B.n64 88.0523
R1025 B.n597 B.n596 88.0523
R1026 B.n596 B.n71 88.0523
R1027 B.n590 B.n71 88.0523
R1028 B.n590 B.n589 88.0523
R1029 B.n589 B.n588 88.0523
R1030 B.n588 B.n78 88.0523
R1031 B.n582 B.n78 88.0523
R1032 B.n582 B.n581 88.0523
R1033 B.n413 B.t14 81.5779
R1034 B.n598 B.t7 81.5779
R1035 B.n381 B.n380 71.676
R1036 B.n375 B.n279 71.676
R1037 B.n372 B.n280 71.676
R1038 B.n368 B.n281 71.676
R1039 B.n364 B.n282 71.676
R1040 B.n360 B.n283 71.676
R1041 B.n356 B.n284 71.676
R1042 B.n352 B.n285 71.676
R1043 B.n347 B.n286 71.676
R1044 B.n343 B.n287 71.676
R1045 B.n339 B.n288 71.676
R1046 B.n335 B.n289 71.676
R1047 B.n331 B.n290 71.676
R1048 B.n327 B.n291 71.676
R1049 B.n323 B.n292 71.676
R1050 B.n319 B.n293 71.676
R1051 B.n315 B.n294 71.676
R1052 B.n311 B.n295 71.676
R1053 B.n307 B.n296 71.676
R1054 B.n383 B.n278 71.676
R1055 B.n110 B.n84 71.676
R1056 B.n114 B.n85 71.676
R1057 B.n118 B.n86 71.676
R1058 B.n122 B.n87 71.676
R1059 B.n126 B.n88 71.676
R1060 B.n130 B.n89 71.676
R1061 B.n134 B.n90 71.676
R1062 B.n138 B.n91 71.676
R1063 B.n142 B.n92 71.676
R1064 B.n146 B.n93 71.676
R1065 B.n150 B.n94 71.676
R1066 B.n154 B.n95 71.676
R1067 B.n158 B.n96 71.676
R1068 B.n163 B.n97 71.676
R1069 B.n167 B.n98 71.676
R1070 B.n171 B.n99 71.676
R1071 B.n175 B.n100 71.676
R1072 B.n179 B.n101 71.676
R1073 B.n183 B.n102 71.676
R1074 B.n187 B.n103 71.676
R1075 B.n104 B.n103 71.676
R1076 B.n186 B.n102 71.676
R1077 B.n182 B.n101 71.676
R1078 B.n178 B.n100 71.676
R1079 B.n174 B.n99 71.676
R1080 B.n170 B.n98 71.676
R1081 B.n166 B.n97 71.676
R1082 B.n162 B.n96 71.676
R1083 B.n157 B.n95 71.676
R1084 B.n153 B.n94 71.676
R1085 B.n149 B.n93 71.676
R1086 B.n145 B.n92 71.676
R1087 B.n141 B.n91 71.676
R1088 B.n137 B.n90 71.676
R1089 B.n133 B.n89 71.676
R1090 B.n129 B.n88 71.676
R1091 B.n125 B.n87 71.676
R1092 B.n121 B.n86 71.676
R1093 B.n117 B.n85 71.676
R1094 B.n113 B.n84 71.676
R1095 B.n381 B.n298 71.676
R1096 B.n373 B.n279 71.676
R1097 B.n369 B.n280 71.676
R1098 B.n365 B.n281 71.676
R1099 B.n361 B.n282 71.676
R1100 B.n357 B.n283 71.676
R1101 B.n353 B.n284 71.676
R1102 B.n348 B.n285 71.676
R1103 B.n344 B.n286 71.676
R1104 B.n340 B.n287 71.676
R1105 B.n336 B.n288 71.676
R1106 B.n332 B.n289 71.676
R1107 B.n328 B.n290 71.676
R1108 B.n324 B.n291 71.676
R1109 B.n320 B.n292 71.676
R1110 B.n316 B.n293 71.676
R1111 B.n312 B.n294 71.676
R1112 B.n308 B.n295 71.676
R1113 B.n304 B.n296 71.676
R1114 B.n384 B.n383 71.676
R1115 B.n497 B.t4 71.2189
R1116 B.n18 B.t1 71.2189
R1117 B.n302 B.n301 60.5096
R1118 B.n300 B.n299 60.5096
R1119 B.n108 B.n107 60.5096
R1120 B.n106 B.n105 60.5096
R1121 B.n303 B.n302 59.5399
R1122 B.n350 B.n300 59.5399
R1123 B.n109 B.n108 59.5399
R1124 B.n160 B.n106 59.5399
R1125 B.n473 B.t5 55.6803
R1126 B.n638 B.t2 55.6803
R1127 B.n449 B.t3 47.911
R1128 B.n622 B.t0 47.911
R1129 B.n239 B.t3 40.1418
R1130 B.t0 B.n621 40.1418
R1131 B.t5 B.n215 32.3725
R1132 B.t2 B.n29 32.3725
R1133 B.n111 B.n80 31.3761
R1134 B.n578 B.n577 31.3761
R1135 B.n386 B.n385 31.3761
R1136 B.n379 B.n273 31.3761
R1137 B B.n672 18.0485
R1138 B.n504 B.t4 16.8339
R1139 B.n660 B.t1 16.8339
R1140 B.n112 B.n111 10.6151
R1141 B.n115 B.n112 10.6151
R1142 B.n116 B.n115 10.6151
R1143 B.n119 B.n116 10.6151
R1144 B.n120 B.n119 10.6151
R1145 B.n123 B.n120 10.6151
R1146 B.n124 B.n123 10.6151
R1147 B.n127 B.n124 10.6151
R1148 B.n128 B.n127 10.6151
R1149 B.n131 B.n128 10.6151
R1150 B.n132 B.n131 10.6151
R1151 B.n135 B.n132 10.6151
R1152 B.n136 B.n135 10.6151
R1153 B.n139 B.n136 10.6151
R1154 B.n140 B.n139 10.6151
R1155 B.n144 B.n143 10.6151
R1156 B.n147 B.n144 10.6151
R1157 B.n148 B.n147 10.6151
R1158 B.n151 B.n148 10.6151
R1159 B.n152 B.n151 10.6151
R1160 B.n155 B.n152 10.6151
R1161 B.n156 B.n155 10.6151
R1162 B.n159 B.n156 10.6151
R1163 B.n164 B.n161 10.6151
R1164 B.n165 B.n164 10.6151
R1165 B.n168 B.n165 10.6151
R1166 B.n169 B.n168 10.6151
R1167 B.n172 B.n169 10.6151
R1168 B.n173 B.n172 10.6151
R1169 B.n176 B.n173 10.6151
R1170 B.n177 B.n176 10.6151
R1171 B.n180 B.n177 10.6151
R1172 B.n181 B.n180 10.6151
R1173 B.n184 B.n181 10.6151
R1174 B.n185 B.n184 10.6151
R1175 B.n188 B.n185 10.6151
R1176 B.n189 B.n188 10.6151
R1177 B.n578 B.n189 10.6151
R1178 B.n387 B.n386 10.6151
R1179 B.n387 B.n269 10.6151
R1180 B.n397 B.n269 10.6151
R1181 B.n398 B.n397 10.6151
R1182 B.n399 B.n398 10.6151
R1183 B.n399 B.n260 10.6151
R1184 B.n409 B.n260 10.6151
R1185 B.n410 B.n409 10.6151
R1186 B.n411 B.n410 10.6151
R1187 B.n411 B.n253 10.6151
R1188 B.n421 B.n253 10.6151
R1189 B.n422 B.n421 10.6151
R1190 B.n423 B.n422 10.6151
R1191 B.n423 B.n245 10.6151
R1192 B.n433 B.n245 10.6151
R1193 B.n434 B.n433 10.6151
R1194 B.n435 B.n434 10.6151
R1195 B.n435 B.n236 10.6151
R1196 B.n445 B.n236 10.6151
R1197 B.n446 B.n445 10.6151
R1198 B.n447 B.n446 10.6151
R1199 B.n447 B.n229 10.6151
R1200 B.n457 B.n229 10.6151
R1201 B.n458 B.n457 10.6151
R1202 B.n459 B.n458 10.6151
R1203 B.n459 B.n221 10.6151
R1204 B.n469 B.n221 10.6151
R1205 B.n470 B.n469 10.6151
R1206 B.n471 B.n470 10.6151
R1207 B.n471 B.n213 10.6151
R1208 B.n481 B.n213 10.6151
R1209 B.n482 B.n481 10.6151
R1210 B.n483 B.n482 10.6151
R1211 B.n483 B.n205 10.6151
R1212 B.n493 B.n205 10.6151
R1213 B.n494 B.n493 10.6151
R1214 B.n495 B.n494 10.6151
R1215 B.n495 B.n198 10.6151
R1216 B.n506 B.n198 10.6151
R1217 B.n507 B.n506 10.6151
R1218 B.n509 B.n507 10.6151
R1219 B.n509 B.n508 10.6151
R1220 B.n508 B.n190 10.6151
R1221 B.n520 B.n190 10.6151
R1222 B.n521 B.n520 10.6151
R1223 B.n522 B.n521 10.6151
R1224 B.n523 B.n522 10.6151
R1225 B.n525 B.n523 10.6151
R1226 B.n526 B.n525 10.6151
R1227 B.n527 B.n526 10.6151
R1228 B.n528 B.n527 10.6151
R1229 B.n530 B.n528 10.6151
R1230 B.n531 B.n530 10.6151
R1231 B.n532 B.n531 10.6151
R1232 B.n533 B.n532 10.6151
R1233 B.n535 B.n533 10.6151
R1234 B.n536 B.n535 10.6151
R1235 B.n537 B.n536 10.6151
R1236 B.n538 B.n537 10.6151
R1237 B.n540 B.n538 10.6151
R1238 B.n541 B.n540 10.6151
R1239 B.n542 B.n541 10.6151
R1240 B.n543 B.n542 10.6151
R1241 B.n545 B.n543 10.6151
R1242 B.n546 B.n545 10.6151
R1243 B.n547 B.n546 10.6151
R1244 B.n548 B.n547 10.6151
R1245 B.n550 B.n548 10.6151
R1246 B.n551 B.n550 10.6151
R1247 B.n552 B.n551 10.6151
R1248 B.n553 B.n552 10.6151
R1249 B.n555 B.n553 10.6151
R1250 B.n556 B.n555 10.6151
R1251 B.n557 B.n556 10.6151
R1252 B.n558 B.n557 10.6151
R1253 B.n560 B.n558 10.6151
R1254 B.n561 B.n560 10.6151
R1255 B.n562 B.n561 10.6151
R1256 B.n563 B.n562 10.6151
R1257 B.n565 B.n563 10.6151
R1258 B.n566 B.n565 10.6151
R1259 B.n567 B.n566 10.6151
R1260 B.n568 B.n567 10.6151
R1261 B.n570 B.n568 10.6151
R1262 B.n571 B.n570 10.6151
R1263 B.n572 B.n571 10.6151
R1264 B.n573 B.n572 10.6151
R1265 B.n575 B.n573 10.6151
R1266 B.n576 B.n575 10.6151
R1267 B.n577 B.n576 10.6151
R1268 B.n379 B.n378 10.6151
R1269 B.n378 B.n377 10.6151
R1270 B.n377 B.n376 10.6151
R1271 B.n376 B.n374 10.6151
R1272 B.n374 B.n371 10.6151
R1273 B.n371 B.n370 10.6151
R1274 B.n370 B.n367 10.6151
R1275 B.n367 B.n366 10.6151
R1276 B.n366 B.n363 10.6151
R1277 B.n363 B.n362 10.6151
R1278 B.n362 B.n359 10.6151
R1279 B.n359 B.n358 10.6151
R1280 B.n358 B.n355 10.6151
R1281 B.n355 B.n354 10.6151
R1282 B.n354 B.n351 10.6151
R1283 B.n349 B.n346 10.6151
R1284 B.n346 B.n345 10.6151
R1285 B.n345 B.n342 10.6151
R1286 B.n342 B.n341 10.6151
R1287 B.n341 B.n338 10.6151
R1288 B.n338 B.n337 10.6151
R1289 B.n337 B.n334 10.6151
R1290 B.n334 B.n333 10.6151
R1291 B.n330 B.n329 10.6151
R1292 B.n329 B.n326 10.6151
R1293 B.n326 B.n325 10.6151
R1294 B.n325 B.n322 10.6151
R1295 B.n322 B.n321 10.6151
R1296 B.n321 B.n318 10.6151
R1297 B.n318 B.n317 10.6151
R1298 B.n317 B.n314 10.6151
R1299 B.n314 B.n313 10.6151
R1300 B.n313 B.n310 10.6151
R1301 B.n310 B.n309 10.6151
R1302 B.n309 B.n306 10.6151
R1303 B.n306 B.n305 10.6151
R1304 B.n305 B.n277 10.6151
R1305 B.n385 B.n277 10.6151
R1306 B.n391 B.n273 10.6151
R1307 B.n392 B.n391 10.6151
R1308 B.n393 B.n392 10.6151
R1309 B.n393 B.n265 10.6151
R1310 B.n403 B.n265 10.6151
R1311 B.n404 B.n403 10.6151
R1312 B.n405 B.n404 10.6151
R1313 B.n405 B.n257 10.6151
R1314 B.n415 B.n257 10.6151
R1315 B.n416 B.n415 10.6151
R1316 B.n417 B.n416 10.6151
R1317 B.n417 B.n249 10.6151
R1318 B.n427 B.n249 10.6151
R1319 B.n428 B.n427 10.6151
R1320 B.n429 B.n428 10.6151
R1321 B.n429 B.n241 10.6151
R1322 B.n439 B.n241 10.6151
R1323 B.n440 B.n439 10.6151
R1324 B.n441 B.n440 10.6151
R1325 B.n441 B.n233 10.6151
R1326 B.n451 B.n233 10.6151
R1327 B.n452 B.n451 10.6151
R1328 B.n453 B.n452 10.6151
R1329 B.n453 B.n225 10.6151
R1330 B.n463 B.n225 10.6151
R1331 B.n464 B.n463 10.6151
R1332 B.n465 B.n464 10.6151
R1333 B.n465 B.n217 10.6151
R1334 B.n475 B.n217 10.6151
R1335 B.n476 B.n475 10.6151
R1336 B.n477 B.n476 10.6151
R1337 B.n477 B.n209 10.6151
R1338 B.n487 B.n209 10.6151
R1339 B.n488 B.n487 10.6151
R1340 B.n489 B.n488 10.6151
R1341 B.n489 B.n201 10.6151
R1342 B.n500 B.n201 10.6151
R1343 B.n501 B.n500 10.6151
R1344 B.n502 B.n501 10.6151
R1345 B.n502 B.n194 10.6151
R1346 B.n513 B.n194 10.6151
R1347 B.n514 B.n513 10.6151
R1348 B.n515 B.n514 10.6151
R1349 B.n515 B.n0 10.6151
R1350 B.n666 B.n1 10.6151
R1351 B.n666 B.n665 10.6151
R1352 B.n665 B.n664 10.6151
R1353 B.n664 B.n10 10.6151
R1354 B.n658 B.n10 10.6151
R1355 B.n658 B.n657 10.6151
R1356 B.n657 B.n656 10.6151
R1357 B.n656 B.n16 10.6151
R1358 B.n650 B.n16 10.6151
R1359 B.n650 B.n649 10.6151
R1360 B.n649 B.n648 10.6151
R1361 B.n648 B.n24 10.6151
R1362 B.n642 B.n24 10.6151
R1363 B.n642 B.n641 10.6151
R1364 B.n641 B.n640 10.6151
R1365 B.n640 B.n31 10.6151
R1366 B.n634 B.n31 10.6151
R1367 B.n634 B.n633 10.6151
R1368 B.n633 B.n632 10.6151
R1369 B.n632 B.n38 10.6151
R1370 B.n626 B.n38 10.6151
R1371 B.n626 B.n625 10.6151
R1372 B.n625 B.n624 10.6151
R1373 B.n624 B.n45 10.6151
R1374 B.n618 B.n45 10.6151
R1375 B.n618 B.n617 10.6151
R1376 B.n617 B.n616 10.6151
R1377 B.n616 B.n52 10.6151
R1378 B.n610 B.n52 10.6151
R1379 B.n610 B.n609 10.6151
R1380 B.n609 B.n608 10.6151
R1381 B.n608 B.n59 10.6151
R1382 B.n602 B.n59 10.6151
R1383 B.n602 B.n601 10.6151
R1384 B.n601 B.n600 10.6151
R1385 B.n600 B.n66 10.6151
R1386 B.n594 B.n66 10.6151
R1387 B.n594 B.n593 10.6151
R1388 B.n593 B.n592 10.6151
R1389 B.n592 B.n73 10.6151
R1390 B.n586 B.n73 10.6151
R1391 B.n586 B.n585 10.6151
R1392 B.n585 B.n584 10.6151
R1393 B.n584 B.n80 10.6151
R1394 B.n143 B.n109 6.5566
R1395 B.n160 B.n159 6.5566
R1396 B.n350 B.n349 6.5566
R1397 B.n333 B.n303 6.5566
R1398 B.n263 B.t14 6.4749
R1399 B.t7 B.n597 6.4749
R1400 B.n140 B.n109 4.05904
R1401 B.n161 B.n160 4.05904
R1402 B.n351 B.n350 4.05904
R1403 B.n330 B.n303 4.05904
R1404 B.n672 B.n0 2.81026
R1405 B.n672 B.n1 2.81026
R1406 VP.n13 VP.n12 161.3
R1407 VP.n14 VP.n9 161.3
R1408 VP.n16 VP.n15 161.3
R1409 VP.n17 VP.n8 161.3
R1410 VP.n19 VP.n18 161.3
R1411 VP.n20 VP.n7 161.3
R1412 VP.n43 VP.n0 161.3
R1413 VP.n42 VP.n41 161.3
R1414 VP.n40 VP.n1 161.3
R1415 VP.n39 VP.n38 161.3
R1416 VP.n37 VP.n2 161.3
R1417 VP.n36 VP.n35 161.3
R1418 VP.n34 VP.n3 161.3
R1419 VP.n33 VP.n32 161.3
R1420 VP.n31 VP.n4 161.3
R1421 VP.n30 VP.n29 161.3
R1422 VP.n28 VP.n5 161.3
R1423 VP.n27 VP.n26 161.3
R1424 VP.n25 VP.n6 161.3
R1425 VP.n24 VP.n23 104.763
R1426 VP.n45 VP.n44 104.763
R1427 VP.n22 VP.n21 104.763
R1428 VP.n11 VP.t1 62.0673
R1429 VP.n11 VP.n10 48.81
R1430 VP.n30 VP.n5 46.253
R1431 VP.n38 VP.n1 46.253
R1432 VP.n15 VP.n8 46.253
R1433 VP.n23 VP.n22 42.7723
R1434 VP.n31 VP.n30 34.5682
R1435 VP.n38 VP.n37 34.5682
R1436 VP.n15 VP.n14 34.5682
R1437 VP.n3 VP.t2 27.8148
R1438 VP.n24 VP.t4 27.8148
R1439 VP.n44 VP.t3 27.8148
R1440 VP.n10 VP.t5 27.8148
R1441 VP.n21 VP.t0 27.8148
R1442 VP.n26 VP.n25 24.3439
R1443 VP.n26 VP.n5 24.3439
R1444 VP.n32 VP.n31 24.3439
R1445 VP.n32 VP.n3 24.3439
R1446 VP.n36 VP.n3 24.3439
R1447 VP.n37 VP.n36 24.3439
R1448 VP.n42 VP.n1 24.3439
R1449 VP.n43 VP.n42 24.3439
R1450 VP.n19 VP.n8 24.3439
R1451 VP.n20 VP.n19 24.3439
R1452 VP.n13 VP.n10 24.3439
R1453 VP.n14 VP.n13 24.3439
R1454 VP.n25 VP.n24 5.84292
R1455 VP.n44 VP.n43 5.84292
R1456 VP.n21 VP.n20 5.84292
R1457 VP.n12 VP.n11 4.95772
R1458 VP.n22 VP.n7 0.278398
R1459 VP.n23 VP.n6 0.278398
R1460 VP.n45 VP.n0 0.278398
R1461 VP.n12 VP.n9 0.189894
R1462 VP.n16 VP.n9 0.189894
R1463 VP.n17 VP.n16 0.189894
R1464 VP.n18 VP.n17 0.189894
R1465 VP.n18 VP.n7 0.189894
R1466 VP.n27 VP.n6 0.189894
R1467 VP.n28 VP.n27 0.189894
R1468 VP.n29 VP.n28 0.189894
R1469 VP.n29 VP.n4 0.189894
R1470 VP.n33 VP.n4 0.189894
R1471 VP.n34 VP.n33 0.189894
R1472 VP.n35 VP.n34 0.189894
R1473 VP.n35 VP.n2 0.189894
R1474 VP.n39 VP.n2 0.189894
R1475 VP.n40 VP.n39 0.189894
R1476 VP.n41 VP.n40 0.189894
R1477 VP.n41 VP.n0 0.189894
R1478 VP VP.n45 0.153422
R1479 VDD1.n10 VDD1.n0 289.615
R1480 VDD1.n25 VDD1.n15 289.615
R1481 VDD1.n11 VDD1.n10 185
R1482 VDD1.n9 VDD1.n8 185
R1483 VDD1.n4 VDD1.n3 185
R1484 VDD1.n19 VDD1.n18 185
R1485 VDD1.n24 VDD1.n23 185
R1486 VDD1.n26 VDD1.n25 185
R1487 VDD1.n5 VDD1.t4 148.606
R1488 VDD1.n20 VDD1.t1 148.606
R1489 VDD1.n10 VDD1.n9 104.615
R1490 VDD1.n9 VDD1.n3 104.615
R1491 VDD1.n24 VDD1.n18 104.615
R1492 VDD1.n25 VDD1.n24 104.615
R1493 VDD1.n31 VDD1.n30 80.3055
R1494 VDD1.n33 VDD1.n32 79.6885
R1495 VDD1 VDD1.n14 52.879
R1496 VDD1.n31 VDD1.n29 52.7654
R1497 VDD1.t4 VDD1.n3 52.3082
R1498 VDD1.t1 VDD1.n18 52.3082
R1499 VDD1.n33 VDD1.n31 37.1604
R1500 VDD1.n5 VDD1.n4 15.5966
R1501 VDD1.n20 VDD1.n19 15.5966
R1502 VDD1.n8 VDD1.n7 12.8005
R1503 VDD1.n23 VDD1.n22 12.8005
R1504 VDD1.n11 VDD1.n2 12.0247
R1505 VDD1.n26 VDD1.n17 12.0247
R1506 VDD1.n12 VDD1.n0 11.249
R1507 VDD1.n27 VDD1.n15 11.249
R1508 VDD1.n14 VDD1.n13 9.45567
R1509 VDD1.n29 VDD1.n28 9.45567
R1510 VDD1.n13 VDD1.n12 9.3005
R1511 VDD1.n2 VDD1.n1 9.3005
R1512 VDD1.n7 VDD1.n6 9.3005
R1513 VDD1.n28 VDD1.n27 9.3005
R1514 VDD1.n17 VDD1.n16 9.3005
R1515 VDD1.n22 VDD1.n21 9.3005
R1516 VDD1.n32 VDD1.t0 6.14957
R1517 VDD1.n32 VDD1.t5 6.14957
R1518 VDD1.n30 VDD1.t3 6.14957
R1519 VDD1.n30 VDD1.t2 6.14957
R1520 VDD1.n6 VDD1.n5 4.46457
R1521 VDD1.n21 VDD1.n20 4.46457
R1522 VDD1.n14 VDD1.n0 2.71565
R1523 VDD1.n29 VDD1.n15 2.71565
R1524 VDD1.n12 VDD1.n11 1.93989
R1525 VDD1.n27 VDD1.n26 1.93989
R1526 VDD1.n8 VDD1.n2 1.16414
R1527 VDD1.n23 VDD1.n17 1.16414
R1528 VDD1 VDD1.n33 0.614724
R1529 VDD1.n7 VDD1.n4 0.388379
R1530 VDD1.n22 VDD1.n19 0.388379
R1531 VDD1.n13 VDD1.n1 0.155672
R1532 VDD1.n6 VDD1.n1 0.155672
R1533 VDD1.n21 VDD1.n16 0.155672
R1534 VDD1.n28 VDD1.n16 0.155672
C0 VDD2 VTAIL 4.72118f
C1 VP VTAIL 2.93616f
C2 VDD2 VDD1 1.47933f
C3 VN VTAIL 2.92201f
C4 VDD1 VP 2.43759f
C5 VDD2 VP 0.478912f
C6 VDD1 VN 0.155476f
C7 VDD1 VTAIL 4.66697f
C8 VDD2 VN 2.11665f
C9 VN VP 5.49543f
C10 VDD2 B 4.559636f
C11 VDD1 B 4.709325f
C12 VTAIL B 4.038346f
C13 VN B 12.654891f
C14 VP B 11.268737f
C15 VDD1.n0 B 0.031278f
C16 VDD1.n1 B 0.022912f
C17 VDD1.n2 B 0.012312f
C18 VDD1.n3 B 0.021826f
C19 VDD1.n4 B 0.016969f
C20 VDD1.t4 B 0.049139f
C21 VDD1.n5 B 0.084982f
C22 VDD1.n6 B 0.248645f
C23 VDD1.n7 B 0.012312f
C24 VDD1.n8 B 0.013036f
C25 VDD1.n9 B 0.029101f
C26 VDD1.n10 B 0.061359f
C27 VDD1.n11 B 0.013036f
C28 VDD1.n12 B 0.012312f
C29 VDD1.n13 B 0.056091f
C30 VDD1.n14 B 0.057871f
C31 VDD1.n15 B 0.031278f
C32 VDD1.n16 B 0.022912f
C33 VDD1.n17 B 0.012312f
C34 VDD1.n18 B 0.021826f
C35 VDD1.n19 B 0.016969f
C36 VDD1.t1 B 0.049139f
C37 VDD1.n20 B 0.084982f
C38 VDD1.n21 B 0.248645f
C39 VDD1.n22 B 0.012312f
C40 VDD1.n23 B 0.013036f
C41 VDD1.n24 B 0.029101f
C42 VDD1.n25 B 0.061359f
C43 VDD1.n26 B 0.013036f
C44 VDD1.n27 B 0.012312f
C45 VDD1.n28 B 0.056091f
C46 VDD1.n29 B 0.057158f
C47 VDD1.t3 B 0.058301f
C48 VDD1.t2 B 0.058301f
C49 VDD1.n30 B 0.44248f
C50 VDD1.n31 B 2.14432f
C51 VDD1.t0 B 0.058301f
C52 VDD1.t5 B 0.058301f
C53 VDD1.n32 B 0.439191f
C54 VDD1.n33 B 1.96526f
C55 VP.n0 B 0.03869f
C56 VP.t3 B 0.66232f
C57 VP.n1 B 0.05625f
C58 VP.n2 B 0.029345f
C59 VP.t2 B 0.66232f
C60 VP.n3 B 0.301232f
C61 VP.n4 B 0.029345f
C62 VP.n5 B 0.05625f
C63 VP.n6 B 0.03869f
C64 VP.t4 B 0.66232f
C65 VP.n7 B 0.03869f
C66 VP.t0 B 0.66232f
C67 VP.n8 B 0.05625f
C68 VP.n9 B 0.029345f
C69 VP.t5 B 0.66232f
C70 VP.n10 B 0.378879f
C71 VP.t1 B 0.922491f
C72 VP.n11 B 0.348292f
C73 VP.n12 B 0.307793f
C74 VP.n13 B 0.054965f
C75 VP.n14 B 0.05962f
C76 VP.n15 B 0.025142f
C77 VP.n16 B 0.029345f
C78 VP.n17 B 0.029345f
C79 VP.n18 B 0.029345f
C80 VP.n19 B 0.054965f
C81 VP.n20 B 0.03434f
C82 VP.n21 B 0.373204f
C83 VP.n22 B 1.29106f
C84 VP.n23 B 1.31565f
C85 VP.n24 B 0.373204f
C86 VP.n25 B 0.03434f
C87 VP.n26 B 0.054965f
C88 VP.n27 B 0.029345f
C89 VP.n28 B 0.029345f
C90 VP.n29 B 0.029345f
C91 VP.n30 B 0.025142f
C92 VP.n31 B 0.05962f
C93 VP.n32 B 0.054965f
C94 VP.n33 B 0.029345f
C95 VP.n34 B 0.029345f
C96 VP.n35 B 0.029345f
C97 VP.n36 B 0.054965f
C98 VP.n37 B 0.05962f
C99 VP.n38 B 0.025142f
C100 VP.n39 B 0.029345f
C101 VP.n40 B 0.029345f
C102 VP.n41 B 0.029345f
C103 VP.n42 B 0.054965f
C104 VP.n43 B 0.03434f
C105 VP.n44 B 0.373204f
C106 VP.n45 B 0.052679f
C107 VTAIL.t6 B 0.079562f
C108 VTAIL.t8 B 0.079562f
C109 VTAIL.n0 B 0.538122f
C110 VTAIL.n1 B 0.51242f
C111 VTAIL.n2 B 0.042684f
C112 VTAIL.n3 B 0.031268f
C113 VTAIL.n4 B 0.016802f
C114 VTAIL.n5 B 0.029785f
C115 VTAIL.n6 B 0.023157f
C116 VTAIL.t4 B 0.067058f
C117 VTAIL.n7 B 0.115973f
C118 VTAIL.n8 B 0.339318f
C119 VTAIL.n9 B 0.016802f
C120 VTAIL.n10 B 0.01779f
C121 VTAIL.n11 B 0.039713f
C122 VTAIL.n12 B 0.083734f
C123 VTAIL.n13 B 0.01779f
C124 VTAIL.n14 B 0.016802f
C125 VTAIL.n15 B 0.076545f
C126 VTAIL.n16 B 0.046751f
C127 VTAIL.n17 B 0.482933f
C128 VTAIL.t3 B 0.079562f
C129 VTAIL.t5 B 0.079562f
C130 VTAIL.n18 B 0.538122f
C131 VTAIL.n19 B 1.77334f
C132 VTAIL.t9 B 0.079562f
C133 VTAIL.t11 B 0.079562f
C134 VTAIL.n20 B 0.538125f
C135 VTAIL.n21 B 1.77334f
C136 VTAIL.n22 B 0.042684f
C137 VTAIL.n23 B 0.031268f
C138 VTAIL.n24 B 0.016802f
C139 VTAIL.n25 B 0.029785f
C140 VTAIL.n26 B 0.023157f
C141 VTAIL.t7 B 0.067058f
C142 VTAIL.n27 B 0.115973f
C143 VTAIL.n28 B 0.339318f
C144 VTAIL.n29 B 0.016802f
C145 VTAIL.n30 B 0.01779f
C146 VTAIL.n31 B 0.039713f
C147 VTAIL.n32 B 0.083734f
C148 VTAIL.n33 B 0.01779f
C149 VTAIL.n34 B 0.016802f
C150 VTAIL.n35 B 0.076545f
C151 VTAIL.n36 B 0.046751f
C152 VTAIL.n37 B 0.482933f
C153 VTAIL.t1 B 0.079562f
C154 VTAIL.t2 B 0.079562f
C155 VTAIL.n38 B 0.538125f
C156 VTAIL.n39 B 0.709793f
C157 VTAIL.n40 B 0.042684f
C158 VTAIL.n41 B 0.031268f
C159 VTAIL.n42 B 0.016802f
C160 VTAIL.n43 B 0.029785f
C161 VTAIL.n44 B 0.023157f
C162 VTAIL.t0 B 0.067058f
C163 VTAIL.n45 B 0.115973f
C164 VTAIL.n46 B 0.339318f
C165 VTAIL.n47 B 0.016802f
C166 VTAIL.n48 B 0.01779f
C167 VTAIL.n49 B 0.039713f
C168 VTAIL.n50 B 0.083734f
C169 VTAIL.n51 B 0.01779f
C170 VTAIL.n52 B 0.016802f
C171 VTAIL.n53 B 0.076545f
C172 VTAIL.n54 B 0.046751f
C173 VTAIL.n55 B 1.27549f
C174 VTAIL.n56 B 0.042684f
C175 VTAIL.n57 B 0.031268f
C176 VTAIL.n58 B 0.016802f
C177 VTAIL.n59 B 0.029785f
C178 VTAIL.n60 B 0.023157f
C179 VTAIL.t10 B 0.067058f
C180 VTAIL.n61 B 0.115973f
C181 VTAIL.n62 B 0.339318f
C182 VTAIL.n63 B 0.016802f
C183 VTAIL.n64 B 0.01779f
C184 VTAIL.n65 B 0.039713f
C185 VTAIL.n66 B 0.083734f
C186 VTAIL.n67 B 0.01779f
C187 VTAIL.n68 B 0.016802f
C188 VTAIL.n69 B 0.076545f
C189 VTAIL.n70 B 0.046751f
C190 VTAIL.n71 B 1.20189f
C191 VDD2.n0 B 0.030318f
C192 VDD2.n1 B 0.022209f
C193 VDD2.n2 B 0.011934f
C194 VDD2.n3 B 0.021156f
C195 VDD2.n4 B 0.016448f
C196 VDD2.t5 B 0.04763f
C197 VDD2.n5 B 0.082373f
C198 VDD2.n6 B 0.241012f
C199 VDD2.n7 B 0.011934f
C200 VDD2.n8 B 0.012636f
C201 VDD2.n9 B 0.028208f
C202 VDD2.n10 B 0.059475f
C203 VDD2.n11 B 0.012636f
C204 VDD2.n12 B 0.011934f
C205 VDD2.n13 B 0.054369f
C206 VDD2.n14 B 0.055403f
C207 VDD2.t3 B 0.056511f
C208 VDD2.t0 B 0.056511f
C209 VDD2.n15 B 0.428896f
C210 VDD2.n16 B 1.97205f
C211 VDD2.n17 B 0.030318f
C212 VDD2.n18 B 0.022209f
C213 VDD2.n19 B 0.011934f
C214 VDD2.n20 B 0.021156f
C215 VDD2.n21 B 0.016448f
C216 VDD2.t4 B 0.04763f
C217 VDD2.n22 B 0.082373f
C218 VDD2.n23 B 0.241012f
C219 VDD2.n24 B 0.011934f
C220 VDD2.n25 B 0.012636f
C221 VDD2.n26 B 0.028208f
C222 VDD2.n27 B 0.059475f
C223 VDD2.n28 B 0.012636f
C224 VDD2.n29 B 0.011934f
C225 VDD2.n30 B 0.054369f
C226 VDD2.n31 B 0.048518f
C227 VDD2.n32 B 1.70846f
C228 VDD2.t1 B 0.056511f
C229 VDD2.t2 B 0.056511f
C230 VDD2.n33 B 0.428873f
C231 VN.n0 B 0.037472f
C232 VN.t1 B 0.641472f
C233 VN.n1 B 0.05448f
C234 VN.n2 B 0.028421f
C235 VN.t3 B 0.641472f
C236 VN.n3 B 0.366953f
C237 VN.t5 B 0.893454f
C238 VN.n4 B 0.337329f
C239 VN.n5 B 0.298104f
C240 VN.n6 B 0.053235f
C241 VN.n7 B 0.057744f
C242 VN.n8 B 0.024351f
C243 VN.n9 B 0.028421f
C244 VN.n10 B 0.028421f
C245 VN.n11 B 0.028421f
C246 VN.n12 B 0.053235f
C247 VN.n13 B 0.033259f
C248 VN.n14 B 0.361457f
C249 VN.n15 B 0.051021f
C250 VN.n16 B 0.037472f
C251 VN.t2 B 0.641472f
C252 VN.n17 B 0.05448f
C253 VN.n18 B 0.028421f
C254 VN.t0 B 0.641472f
C255 VN.n19 B 0.366953f
C256 VN.t4 B 0.893454f
C257 VN.n20 B 0.337329f
C258 VN.n21 B 0.298104f
C259 VN.n22 B 0.053235f
C260 VN.n23 B 0.057744f
C261 VN.n24 B 0.024351f
C262 VN.n25 B 0.028421f
C263 VN.n26 B 0.028421f
C264 VN.n27 B 0.028421f
C265 VN.n28 B 0.053235f
C266 VN.n29 B 0.033259f
C267 VN.n30 B 0.361457f
C268 VN.n31 B 1.2661f
.ends

