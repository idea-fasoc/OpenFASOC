* NGSPICE file created from diff_pair_sample_0921.ext - technology: sky130A

.subckt diff_pair_sample_0921 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t7 VP.t0 VTAIL.t12 B.t3 sky130_fd_pr__nfet_01v8 ad=1.6236 pd=10.17 as=1.6236 ps=10.17 w=9.84 l=0.83
X1 VTAIL.t9 VP.t1 VDD1.t6 B.t1 sky130_fd_pr__nfet_01v8 ad=3.8376 pd=20.46 as=1.6236 ps=10.17 w=9.84 l=0.83
X2 VDD2.t7 VN.t0 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=1.6236 pd=10.17 as=1.6236 ps=10.17 w=9.84 l=0.83
X3 VDD1.t5 VP.t2 VTAIL.t8 B.t4 sky130_fd_pr__nfet_01v8 ad=1.6236 pd=10.17 as=3.8376 ps=20.46 w=9.84 l=0.83
X4 VTAIL.t13 VP.t3 VDD1.t4 B.t7 sky130_fd_pr__nfet_01v8 ad=3.8376 pd=20.46 as=1.6236 ps=10.17 w=9.84 l=0.83
X5 VDD2.t6 VN.t1 VTAIL.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=1.6236 pd=10.17 as=3.8376 ps=20.46 w=9.84 l=0.83
X6 VDD1.t3 VP.t4 VTAIL.t11 B.t6 sky130_fd_pr__nfet_01v8 ad=1.6236 pd=10.17 as=3.8376 ps=20.46 w=9.84 l=0.83
X7 VTAIL.t5 VN.t2 VDD2.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=1.6236 pd=10.17 as=1.6236 ps=10.17 w=9.84 l=0.83
X8 B.t21 B.t19 B.t20 B.t16 sky130_fd_pr__nfet_01v8 ad=3.8376 pd=20.46 as=0 ps=0 w=9.84 l=0.83
X9 B.t18 B.t15 B.t17 B.t16 sky130_fd_pr__nfet_01v8 ad=3.8376 pd=20.46 as=0 ps=0 w=9.84 l=0.83
X10 B.t14 B.t12 B.t13 B.t9 sky130_fd_pr__nfet_01v8 ad=3.8376 pd=20.46 as=0 ps=0 w=9.84 l=0.83
X11 VTAIL.t2 VN.t3 VDD2.t4 B.t2 sky130_fd_pr__nfet_01v8 ad=1.6236 pd=10.17 as=1.6236 ps=10.17 w=9.84 l=0.83
X12 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=3.8376 pd=20.46 as=0 ps=0 w=9.84 l=0.83
X13 VDD2.t3 VN.t4 VTAIL.t6 B.t6 sky130_fd_pr__nfet_01v8 ad=1.6236 pd=10.17 as=3.8376 ps=20.46 w=9.84 l=0.83
X14 VTAIL.t1 VN.t5 VDD2.t2 B.t1 sky130_fd_pr__nfet_01v8 ad=3.8376 pd=20.46 as=1.6236 ps=10.17 w=9.84 l=0.83
X15 VDD1.t2 VP.t5 VTAIL.t14 B.t0 sky130_fd_pr__nfet_01v8 ad=1.6236 pd=10.17 as=1.6236 ps=10.17 w=9.84 l=0.83
X16 VTAIL.t15 VP.t6 VDD1.t1 B.t2 sky130_fd_pr__nfet_01v8 ad=1.6236 pd=10.17 as=1.6236 ps=10.17 w=9.84 l=0.83
X17 VDD2.t1 VN.t6 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=1.6236 pd=10.17 as=1.6236 ps=10.17 w=9.84 l=0.83
X18 VTAIL.t7 VN.t7 VDD2.t0 B.t7 sky130_fd_pr__nfet_01v8 ad=3.8376 pd=20.46 as=1.6236 ps=10.17 w=9.84 l=0.83
X19 VTAIL.t10 VP.t7 VDD1.t0 B.t5 sky130_fd_pr__nfet_01v8 ad=1.6236 pd=10.17 as=1.6236 ps=10.17 w=9.84 l=0.83
R0 VP.n7 VP.t1 352.868
R1 VP.n17 VP.t3 333.046
R2 VP.n29 VP.t4 333.046
R3 VP.n15 VP.t2 333.046
R4 VP.n22 VP.t5 285.716
R5 VP.n1 VP.t6 285.716
R6 VP.n5 VP.t7 285.716
R7 VP.n8 VP.t0 285.716
R8 VP.n30 VP.n29 161.3
R9 VP.n9 VP.n6 161.3
R10 VP.n11 VP.n10 161.3
R11 VP.n13 VP.n12 161.3
R12 VP.n14 VP.n4 161.3
R13 VP.n16 VP.n15 161.3
R14 VP.n28 VP.n0 161.3
R15 VP.n27 VP.n26 161.3
R16 VP.n25 VP.n24 161.3
R17 VP.n23 VP.n2 161.3
R18 VP.n21 VP.n20 161.3
R19 VP.n19 VP.n3 161.3
R20 VP.n18 VP.n17 161.3
R21 VP.n24 VP.n23 56.5617
R22 VP.n10 VP.n9 56.5617
R23 VP.n21 VP.n3 49.296
R24 VP.n28 VP.n27 49.296
R25 VP.n14 VP.n13 49.296
R26 VP.n7 VP.n6 43.0963
R27 VP.n18 VP.n16 40.955
R28 VP.n8 VP.n7 38.2995
R29 VP.n23 VP.n22 16.2311
R30 VP.n24 VP.n1 16.2311
R31 VP.n10 VP.n5 16.2311
R32 VP.n9 VP.n8 16.2311
R33 VP.n17 VP.n3 10.955
R34 VP.n29 VP.n28 10.955
R35 VP.n15 VP.n14 10.955
R36 VP.n22 VP.n21 8.36172
R37 VP.n27 VP.n1 8.36172
R38 VP.n13 VP.n5 8.36172
R39 VP.n11 VP.n6 0.189894
R40 VP.n12 VP.n11 0.189894
R41 VP.n12 VP.n4 0.189894
R42 VP.n16 VP.n4 0.189894
R43 VP.n19 VP.n18 0.189894
R44 VP.n20 VP.n19 0.189894
R45 VP.n20 VP.n2 0.189894
R46 VP.n25 VP.n2 0.189894
R47 VP.n26 VP.n25 0.189894
R48 VP.n26 VP.n0 0.189894
R49 VP.n30 VP.n0 0.189894
R50 VP VP.n30 0.0516364
R51 VTAIL.n11 VTAIL.t9 46.2788
R52 VTAIL.n10 VTAIL.t6 46.2788
R53 VTAIL.n7 VTAIL.t7 46.2788
R54 VTAIL.n14 VTAIL.t8 46.2788
R55 VTAIL.n15 VTAIL.t4 46.2786
R56 VTAIL.n2 VTAIL.t1 46.2786
R57 VTAIL.n3 VTAIL.t11 46.2786
R58 VTAIL.n6 VTAIL.t13 46.2786
R59 VTAIL.n13 VTAIL.n12 44.2666
R60 VTAIL.n9 VTAIL.n8 44.2666
R61 VTAIL.n1 VTAIL.n0 44.2664
R62 VTAIL.n5 VTAIL.n4 44.2664
R63 VTAIL.n15 VTAIL.n14 21.8496
R64 VTAIL.n7 VTAIL.n6 21.8496
R65 VTAIL.n0 VTAIL.t3 2.0127
R66 VTAIL.n0 VTAIL.t5 2.0127
R67 VTAIL.n4 VTAIL.t14 2.0127
R68 VTAIL.n4 VTAIL.t15 2.0127
R69 VTAIL.n12 VTAIL.t12 2.0127
R70 VTAIL.n12 VTAIL.t10 2.0127
R71 VTAIL.n8 VTAIL.t0 2.0127
R72 VTAIL.n8 VTAIL.t2 2.0127
R73 VTAIL.n9 VTAIL.n7 1.0005
R74 VTAIL.n10 VTAIL.n9 1.0005
R75 VTAIL.n13 VTAIL.n11 1.0005
R76 VTAIL.n14 VTAIL.n13 1.0005
R77 VTAIL.n6 VTAIL.n5 1.0005
R78 VTAIL.n5 VTAIL.n3 1.0005
R79 VTAIL.n2 VTAIL.n1 1.0005
R80 VTAIL VTAIL.n15 0.94231
R81 VTAIL.n11 VTAIL.n10 0.470328
R82 VTAIL.n3 VTAIL.n2 0.470328
R83 VTAIL VTAIL.n1 0.0586897
R84 VDD1 VDD1.n0 61.5036
R85 VDD1.n3 VDD1.n2 61.3899
R86 VDD1.n3 VDD1.n1 61.3899
R87 VDD1.n5 VDD1.n4 60.9454
R88 VDD1.n5 VDD1.n3 37.2811
R89 VDD1.n4 VDD1.t0 2.0127
R90 VDD1.n4 VDD1.t5 2.0127
R91 VDD1.n0 VDD1.t6 2.0127
R92 VDD1.n0 VDD1.t7 2.0127
R93 VDD1.n2 VDD1.t1 2.0127
R94 VDD1.n2 VDD1.t3 2.0127
R95 VDD1.n1 VDD1.t4 2.0127
R96 VDD1.n1 VDD1.t2 2.0127
R97 VDD1 VDD1.n5 0.44231
R98 B.n613 B.n612 585
R99 B.n251 B.n88 585
R100 B.n250 B.n249 585
R101 B.n248 B.n247 585
R102 B.n246 B.n245 585
R103 B.n244 B.n243 585
R104 B.n242 B.n241 585
R105 B.n240 B.n239 585
R106 B.n238 B.n237 585
R107 B.n236 B.n235 585
R108 B.n234 B.n233 585
R109 B.n232 B.n231 585
R110 B.n230 B.n229 585
R111 B.n228 B.n227 585
R112 B.n226 B.n225 585
R113 B.n224 B.n223 585
R114 B.n222 B.n221 585
R115 B.n220 B.n219 585
R116 B.n218 B.n217 585
R117 B.n216 B.n215 585
R118 B.n214 B.n213 585
R119 B.n212 B.n211 585
R120 B.n210 B.n209 585
R121 B.n208 B.n207 585
R122 B.n206 B.n205 585
R123 B.n204 B.n203 585
R124 B.n202 B.n201 585
R125 B.n200 B.n199 585
R126 B.n198 B.n197 585
R127 B.n196 B.n195 585
R128 B.n194 B.n193 585
R129 B.n192 B.n191 585
R130 B.n190 B.n189 585
R131 B.n188 B.n187 585
R132 B.n186 B.n185 585
R133 B.n183 B.n182 585
R134 B.n181 B.n180 585
R135 B.n179 B.n178 585
R136 B.n177 B.n176 585
R137 B.n175 B.n174 585
R138 B.n173 B.n172 585
R139 B.n171 B.n170 585
R140 B.n169 B.n168 585
R141 B.n167 B.n166 585
R142 B.n165 B.n164 585
R143 B.n162 B.n161 585
R144 B.n160 B.n159 585
R145 B.n158 B.n157 585
R146 B.n156 B.n155 585
R147 B.n154 B.n153 585
R148 B.n152 B.n151 585
R149 B.n150 B.n149 585
R150 B.n148 B.n147 585
R151 B.n146 B.n145 585
R152 B.n144 B.n143 585
R153 B.n142 B.n141 585
R154 B.n140 B.n139 585
R155 B.n138 B.n137 585
R156 B.n136 B.n135 585
R157 B.n134 B.n133 585
R158 B.n132 B.n131 585
R159 B.n130 B.n129 585
R160 B.n128 B.n127 585
R161 B.n126 B.n125 585
R162 B.n124 B.n123 585
R163 B.n122 B.n121 585
R164 B.n120 B.n119 585
R165 B.n118 B.n117 585
R166 B.n116 B.n115 585
R167 B.n114 B.n113 585
R168 B.n112 B.n111 585
R169 B.n110 B.n109 585
R170 B.n108 B.n107 585
R171 B.n106 B.n105 585
R172 B.n104 B.n103 585
R173 B.n102 B.n101 585
R174 B.n100 B.n99 585
R175 B.n98 B.n97 585
R176 B.n96 B.n95 585
R177 B.n94 B.n93 585
R178 B.n611 B.n48 585
R179 B.n616 B.n48 585
R180 B.n610 B.n47 585
R181 B.n617 B.n47 585
R182 B.n609 B.n608 585
R183 B.n608 B.n43 585
R184 B.n607 B.n42 585
R185 B.n623 B.n42 585
R186 B.n606 B.n41 585
R187 B.n624 B.n41 585
R188 B.n605 B.n40 585
R189 B.n625 B.n40 585
R190 B.n604 B.n603 585
R191 B.n603 B.n36 585
R192 B.n602 B.n35 585
R193 B.n631 B.n35 585
R194 B.n601 B.n34 585
R195 B.n632 B.n34 585
R196 B.n600 B.n33 585
R197 B.n633 B.n33 585
R198 B.n599 B.n598 585
R199 B.n598 B.n29 585
R200 B.n597 B.n28 585
R201 B.n639 B.n28 585
R202 B.n596 B.n27 585
R203 B.n640 B.n27 585
R204 B.n595 B.n26 585
R205 B.n641 B.n26 585
R206 B.n594 B.n593 585
R207 B.n593 B.n25 585
R208 B.n592 B.n21 585
R209 B.n647 B.n21 585
R210 B.n591 B.n20 585
R211 B.n648 B.n20 585
R212 B.n590 B.n19 585
R213 B.n649 B.n19 585
R214 B.n589 B.n588 585
R215 B.n588 B.n18 585
R216 B.n587 B.n14 585
R217 B.n655 B.n14 585
R218 B.n586 B.n13 585
R219 B.n656 B.n13 585
R220 B.n585 B.n12 585
R221 B.n657 B.n12 585
R222 B.n584 B.n583 585
R223 B.n583 B.n8 585
R224 B.n582 B.n7 585
R225 B.n663 B.n7 585
R226 B.n581 B.n6 585
R227 B.n664 B.n6 585
R228 B.n580 B.n5 585
R229 B.n665 B.n5 585
R230 B.n579 B.n578 585
R231 B.n578 B.n4 585
R232 B.n577 B.n252 585
R233 B.n577 B.n576 585
R234 B.n567 B.n253 585
R235 B.n254 B.n253 585
R236 B.n569 B.n568 585
R237 B.n570 B.n569 585
R238 B.n566 B.n259 585
R239 B.n259 B.n258 585
R240 B.n565 B.n564 585
R241 B.n564 B.n563 585
R242 B.n261 B.n260 585
R243 B.n556 B.n261 585
R244 B.n555 B.n554 585
R245 B.n557 B.n555 585
R246 B.n553 B.n266 585
R247 B.n266 B.n265 585
R248 B.n552 B.n551 585
R249 B.n551 B.n550 585
R250 B.n268 B.n267 585
R251 B.n543 B.n268 585
R252 B.n542 B.n541 585
R253 B.n544 B.n542 585
R254 B.n540 B.n273 585
R255 B.n273 B.n272 585
R256 B.n539 B.n538 585
R257 B.n538 B.n537 585
R258 B.n275 B.n274 585
R259 B.n276 B.n275 585
R260 B.n530 B.n529 585
R261 B.n531 B.n530 585
R262 B.n528 B.n281 585
R263 B.n281 B.n280 585
R264 B.n527 B.n526 585
R265 B.n526 B.n525 585
R266 B.n283 B.n282 585
R267 B.n284 B.n283 585
R268 B.n518 B.n517 585
R269 B.n519 B.n518 585
R270 B.n516 B.n288 585
R271 B.n292 B.n288 585
R272 B.n515 B.n514 585
R273 B.n514 B.n513 585
R274 B.n290 B.n289 585
R275 B.n291 B.n290 585
R276 B.n506 B.n505 585
R277 B.n507 B.n506 585
R278 B.n504 B.n297 585
R279 B.n297 B.n296 585
R280 B.n499 B.n498 585
R281 B.n497 B.n339 585
R282 B.n496 B.n338 585
R283 B.n501 B.n338 585
R284 B.n495 B.n494 585
R285 B.n493 B.n492 585
R286 B.n491 B.n490 585
R287 B.n489 B.n488 585
R288 B.n487 B.n486 585
R289 B.n485 B.n484 585
R290 B.n483 B.n482 585
R291 B.n481 B.n480 585
R292 B.n479 B.n478 585
R293 B.n477 B.n476 585
R294 B.n475 B.n474 585
R295 B.n473 B.n472 585
R296 B.n471 B.n470 585
R297 B.n469 B.n468 585
R298 B.n467 B.n466 585
R299 B.n465 B.n464 585
R300 B.n463 B.n462 585
R301 B.n461 B.n460 585
R302 B.n459 B.n458 585
R303 B.n457 B.n456 585
R304 B.n455 B.n454 585
R305 B.n453 B.n452 585
R306 B.n451 B.n450 585
R307 B.n449 B.n448 585
R308 B.n447 B.n446 585
R309 B.n445 B.n444 585
R310 B.n443 B.n442 585
R311 B.n441 B.n440 585
R312 B.n439 B.n438 585
R313 B.n437 B.n436 585
R314 B.n435 B.n434 585
R315 B.n433 B.n432 585
R316 B.n431 B.n430 585
R317 B.n429 B.n428 585
R318 B.n427 B.n426 585
R319 B.n425 B.n424 585
R320 B.n423 B.n422 585
R321 B.n421 B.n420 585
R322 B.n419 B.n418 585
R323 B.n417 B.n416 585
R324 B.n415 B.n414 585
R325 B.n413 B.n412 585
R326 B.n411 B.n410 585
R327 B.n409 B.n408 585
R328 B.n407 B.n406 585
R329 B.n405 B.n404 585
R330 B.n403 B.n402 585
R331 B.n401 B.n400 585
R332 B.n399 B.n398 585
R333 B.n397 B.n396 585
R334 B.n395 B.n394 585
R335 B.n393 B.n392 585
R336 B.n391 B.n390 585
R337 B.n389 B.n388 585
R338 B.n387 B.n386 585
R339 B.n385 B.n384 585
R340 B.n383 B.n382 585
R341 B.n381 B.n380 585
R342 B.n379 B.n378 585
R343 B.n377 B.n376 585
R344 B.n375 B.n374 585
R345 B.n373 B.n372 585
R346 B.n371 B.n370 585
R347 B.n369 B.n368 585
R348 B.n367 B.n366 585
R349 B.n365 B.n364 585
R350 B.n363 B.n362 585
R351 B.n361 B.n360 585
R352 B.n359 B.n358 585
R353 B.n357 B.n356 585
R354 B.n355 B.n354 585
R355 B.n353 B.n352 585
R356 B.n351 B.n350 585
R357 B.n349 B.n348 585
R358 B.n347 B.n346 585
R359 B.n299 B.n298 585
R360 B.n503 B.n502 585
R361 B.n502 B.n501 585
R362 B.n295 B.n294 585
R363 B.n296 B.n295 585
R364 B.n509 B.n508 585
R365 B.n508 B.n507 585
R366 B.n510 B.n293 585
R367 B.n293 B.n291 585
R368 B.n512 B.n511 585
R369 B.n513 B.n512 585
R370 B.n287 B.n286 585
R371 B.n292 B.n287 585
R372 B.n521 B.n520 585
R373 B.n520 B.n519 585
R374 B.n522 B.n285 585
R375 B.n285 B.n284 585
R376 B.n524 B.n523 585
R377 B.n525 B.n524 585
R378 B.n279 B.n278 585
R379 B.n280 B.n279 585
R380 B.n533 B.n532 585
R381 B.n532 B.n531 585
R382 B.n534 B.n277 585
R383 B.n277 B.n276 585
R384 B.n536 B.n535 585
R385 B.n537 B.n536 585
R386 B.n271 B.n270 585
R387 B.n272 B.n271 585
R388 B.n546 B.n545 585
R389 B.n545 B.n544 585
R390 B.n547 B.n269 585
R391 B.n543 B.n269 585
R392 B.n549 B.n548 585
R393 B.n550 B.n549 585
R394 B.n264 B.n263 585
R395 B.n265 B.n264 585
R396 B.n559 B.n558 585
R397 B.n558 B.n557 585
R398 B.n560 B.n262 585
R399 B.n556 B.n262 585
R400 B.n562 B.n561 585
R401 B.n563 B.n562 585
R402 B.n257 B.n256 585
R403 B.n258 B.n257 585
R404 B.n572 B.n571 585
R405 B.n571 B.n570 585
R406 B.n573 B.n255 585
R407 B.n255 B.n254 585
R408 B.n575 B.n574 585
R409 B.n576 B.n575 585
R410 B.n2 B.n0 585
R411 B.n4 B.n2 585
R412 B.n3 B.n1 585
R413 B.n664 B.n3 585
R414 B.n662 B.n661 585
R415 B.n663 B.n662 585
R416 B.n660 B.n9 585
R417 B.n9 B.n8 585
R418 B.n659 B.n658 585
R419 B.n658 B.n657 585
R420 B.n11 B.n10 585
R421 B.n656 B.n11 585
R422 B.n654 B.n653 585
R423 B.n655 B.n654 585
R424 B.n652 B.n15 585
R425 B.n18 B.n15 585
R426 B.n651 B.n650 585
R427 B.n650 B.n649 585
R428 B.n17 B.n16 585
R429 B.n648 B.n17 585
R430 B.n646 B.n645 585
R431 B.n647 B.n646 585
R432 B.n644 B.n22 585
R433 B.n25 B.n22 585
R434 B.n643 B.n642 585
R435 B.n642 B.n641 585
R436 B.n24 B.n23 585
R437 B.n640 B.n24 585
R438 B.n638 B.n637 585
R439 B.n639 B.n638 585
R440 B.n636 B.n30 585
R441 B.n30 B.n29 585
R442 B.n635 B.n634 585
R443 B.n634 B.n633 585
R444 B.n32 B.n31 585
R445 B.n632 B.n32 585
R446 B.n630 B.n629 585
R447 B.n631 B.n630 585
R448 B.n628 B.n37 585
R449 B.n37 B.n36 585
R450 B.n627 B.n626 585
R451 B.n626 B.n625 585
R452 B.n39 B.n38 585
R453 B.n624 B.n39 585
R454 B.n622 B.n621 585
R455 B.n623 B.n622 585
R456 B.n620 B.n44 585
R457 B.n44 B.n43 585
R458 B.n619 B.n618 585
R459 B.n618 B.n617 585
R460 B.n46 B.n45 585
R461 B.n616 B.n46 585
R462 B.n667 B.n666 585
R463 B.n666 B.n665 585
R464 B.n499 B.n295 535.745
R465 B.n93 B.n46 535.745
R466 B.n502 B.n297 535.745
R467 B.n613 B.n48 535.745
R468 B.n343 B.t19 487.332
R469 B.n340 B.t15 487.332
R470 B.n91 B.t8 487.332
R471 B.n89 B.t12 487.332
R472 B.n615 B.n614 256.663
R473 B.n615 B.n87 256.663
R474 B.n615 B.n86 256.663
R475 B.n615 B.n85 256.663
R476 B.n615 B.n84 256.663
R477 B.n615 B.n83 256.663
R478 B.n615 B.n82 256.663
R479 B.n615 B.n81 256.663
R480 B.n615 B.n80 256.663
R481 B.n615 B.n79 256.663
R482 B.n615 B.n78 256.663
R483 B.n615 B.n77 256.663
R484 B.n615 B.n76 256.663
R485 B.n615 B.n75 256.663
R486 B.n615 B.n74 256.663
R487 B.n615 B.n73 256.663
R488 B.n615 B.n72 256.663
R489 B.n615 B.n71 256.663
R490 B.n615 B.n70 256.663
R491 B.n615 B.n69 256.663
R492 B.n615 B.n68 256.663
R493 B.n615 B.n67 256.663
R494 B.n615 B.n66 256.663
R495 B.n615 B.n65 256.663
R496 B.n615 B.n64 256.663
R497 B.n615 B.n63 256.663
R498 B.n615 B.n62 256.663
R499 B.n615 B.n61 256.663
R500 B.n615 B.n60 256.663
R501 B.n615 B.n59 256.663
R502 B.n615 B.n58 256.663
R503 B.n615 B.n57 256.663
R504 B.n615 B.n56 256.663
R505 B.n615 B.n55 256.663
R506 B.n615 B.n54 256.663
R507 B.n615 B.n53 256.663
R508 B.n615 B.n52 256.663
R509 B.n615 B.n51 256.663
R510 B.n615 B.n50 256.663
R511 B.n615 B.n49 256.663
R512 B.n501 B.n500 256.663
R513 B.n501 B.n300 256.663
R514 B.n501 B.n301 256.663
R515 B.n501 B.n302 256.663
R516 B.n501 B.n303 256.663
R517 B.n501 B.n304 256.663
R518 B.n501 B.n305 256.663
R519 B.n501 B.n306 256.663
R520 B.n501 B.n307 256.663
R521 B.n501 B.n308 256.663
R522 B.n501 B.n309 256.663
R523 B.n501 B.n310 256.663
R524 B.n501 B.n311 256.663
R525 B.n501 B.n312 256.663
R526 B.n501 B.n313 256.663
R527 B.n501 B.n314 256.663
R528 B.n501 B.n315 256.663
R529 B.n501 B.n316 256.663
R530 B.n501 B.n317 256.663
R531 B.n501 B.n318 256.663
R532 B.n501 B.n319 256.663
R533 B.n501 B.n320 256.663
R534 B.n501 B.n321 256.663
R535 B.n501 B.n322 256.663
R536 B.n501 B.n323 256.663
R537 B.n501 B.n324 256.663
R538 B.n501 B.n325 256.663
R539 B.n501 B.n326 256.663
R540 B.n501 B.n327 256.663
R541 B.n501 B.n328 256.663
R542 B.n501 B.n329 256.663
R543 B.n501 B.n330 256.663
R544 B.n501 B.n331 256.663
R545 B.n501 B.n332 256.663
R546 B.n501 B.n333 256.663
R547 B.n501 B.n334 256.663
R548 B.n501 B.n335 256.663
R549 B.n501 B.n336 256.663
R550 B.n501 B.n337 256.663
R551 B.n508 B.n295 163.367
R552 B.n508 B.n293 163.367
R553 B.n512 B.n293 163.367
R554 B.n512 B.n287 163.367
R555 B.n520 B.n287 163.367
R556 B.n520 B.n285 163.367
R557 B.n524 B.n285 163.367
R558 B.n524 B.n279 163.367
R559 B.n532 B.n279 163.367
R560 B.n532 B.n277 163.367
R561 B.n536 B.n277 163.367
R562 B.n536 B.n271 163.367
R563 B.n545 B.n271 163.367
R564 B.n545 B.n269 163.367
R565 B.n549 B.n269 163.367
R566 B.n549 B.n264 163.367
R567 B.n558 B.n264 163.367
R568 B.n558 B.n262 163.367
R569 B.n562 B.n262 163.367
R570 B.n562 B.n257 163.367
R571 B.n571 B.n257 163.367
R572 B.n571 B.n255 163.367
R573 B.n575 B.n255 163.367
R574 B.n575 B.n2 163.367
R575 B.n666 B.n2 163.367
R576 B.n666 B.n3 163.367
R577 B.n662 B.n3 163.367
R578 B.n662 B.n9 163.367
R579 B.n658 B.n9 163.367
R580 B.n658 B.n11 163.367
R581 B.n654 B.n11 163.367
R582 B.n654 B.n15 163.367
R583 B.n650 B.n15 163.367
R584 B.n650 B.n17 163.367
R585 B.n646 B.n17 163.367
R586 B.n646 B.n22 163.367
R587 B.n642 B.n22 163.367
R588 B.n642 B.n24 163.367
R589 B.n638 B.n24 163.367
R590 B.n638 B.n30 163.367
R591 B.n634 B.n30 163.367
R592 B.n634 B.n32 163.367
R593 B.n630 B.n32 163.367
R594 B.n630 B.n37 163.367
R595 B.n626 B.n37 163.367
R596 B.n626 B.n39 163.367
R597 B.n622 B.n39 163.367
R598 B.n622 B.n44 163.367
R599 B.n618 B.n44 163.367
R600 B.n618 B.n46 163.367
R601 B.n339 B.n338 163.367
R602 B.n494 B.n338 163.367
R603 B.n492 B.n491 163.367
R604 B.n488 B.n487 163.367
R605 B.n484 B.n483 163.367
R606 B.n480 B.n479 163.367
R607 B.n476 B.n475 163.367
R608 B.n472 B.n471 163.367
R609 B.n468 B.n467 163.367
R610 B.n464 B.n463 163.367
R611 B.n460 B.n459 163.367
R612 B.n456 B.n455 163.367
R613 B.n452 B.n451 163.367
R614 B.n448 B.n447 163.367
R615 B.n444 B.n443 163.367
R616 B.n440 B.n439 163.367
R617 B.n436 B.n435 163.367
R618 B.n432 B.n431 163.367
R619 B.n428 B.n427 163.367
R620 B.n424 B.n423 163.367
R621 B.n420 B.n419 163.367
R622 B.n416 B.n415 163.367
R623 B.n412 B.n411 163.367
R624 B.n408 B.n407 163.367
R625 B.n404 B.n403 163.367
R626 B.n400 B.n399 163.367
R627 B.n396 B.n395 163.367
R628 B.n392 B.n391 163.367
R629 B.n388 B.n387 163.367
R630 B.n384 B.n383 163.367
R631 B.n380 B.n379 163.367
R632 B.n376 B.n375 163.367
R633 B.n372 B.n371 163.367
R634 B.n368 B.n367 163.367
R635 B.n364 B.n363 163.367
R636 B.n360 B.n359 163.367
R637 B.n356 B.n355 163.367
R638 B.n352 B.n351 163.367
R639 B.n348 B.n347 163.367
R640 B.n502 B.n299 163.367
R641 B.n506 B.n297 163.367
R642 B.n506 B.n290 163.367
R643 B.n514 B.n290 163.367
R644 B.n514 B.n288 163.367
R645 B.n518 B.n288 163.367
R646 B.n518 B.n283 163.367
R647 B.n526 B.n283 163.367
R648 B.n526 B.n281 163.367
R649 B.n530 B.n281 163.367
R650 B.n530 B.n275 163.367
R651 B.n538 B.n275 163.367
R652 B.n538 B.n273 163.367
R653 B.n542 B.n273 163.367
R654 B.n542 B.n268 163.367
R655 B.n551 B.n268 163.367
R656 B.n551 B.n266 163.367
R657 B.n555 B.n266 163.367
R658 B.n555 B.n261 163.367
R659 B.n564 B.n261 163.367
R660 B.n564 B.n259 163.367
R661 B.n569 B.n259 163.367
R662 B.n569 B.n253 163.367
R663 B.n577 B.n253 163.367
R664 B.n578 B.n577 163.367
R665 B.n578 B.n5 163.367
R666 B.n6 B.n5 163.367
R667 B.n7 B.n6 163.367
R668 B.n583 B.n7 163.367
R669 B.n583 B.n12 163.367
R670 B.n13 B.n12 163.367
R671 B.n14 B.n13 163.367
R672 B.n588 B.n14 163.367
R673 B.n588 B.n19 163.367
R674 B.n20 B.n19 163.367
R675 B.n21 B.n20 163.367
R676 B.n593 B.n21 163.367
R677 B.n593 B.n26 163.367
R678 B.n27 B.n26 163.367
R679 B.n28 B.n27 163.367
R680 B.n598 B.n28 163.367
R681 B.n598 B.n33 163.367
R682 B.n34 B.n33 163.367
R683 B.n35 B.n34 163.367
R684 B.n603 B.n35 163.367
R685 B.n603 B.n40 163.367
R686 B.n41 B.n40 163.367
R687 B.n42 B.n41 163.367
R688 B.n608 B.n42 163.367
R689 B.n608 B.n47 163.367
R690 B.n48 B.n47 163.367
R691 B.n97 B.n96 163.367
R692 B.n101 B.n100 163.367
R693 B.n105 B.n104 163.367
R694 B.n109 B.n108 163.367
R695 B.n113 B.n112 163.367
R696 B.n117 B.n116 163.367
R697 B.n121 B.n120 163.367
R698 B.n125 B.n124 163.367
R699 B.n129 B.n128 163.367
R700 B.n133 B.n132 163.367
R701 B.n137 B.n136 163.367
R702 B.n141 B.n140 163.367
R703 B.n145 B.n144 163.367
R704 B.n149 B.n148 163.367
R705 B.n153 B.n152 163.367
R706 B.n157 B.n156 163.367
R707 B.n161 B.n160 163.367
R708 B.n166 B.n165 163.367
R709 B.n170 B.n169 163.367
R710 B.n174 B.n173 163.367
R711 B.n178 B.n177 163.367
R712 B.n182 B.n181 163.367
R713 B.n187 B.n186 163.367
R714 B.n191 B.n190 163.367
R715 B.n195 B.n194 163.367
R716 B.n199 B.n198 163.367
R717 B.n203 B.n202 163.367
R718 B.n207 B.n206 163.367
R719 B.n211 B.n210 163.367
R720 B.n215 B.n214 163.367
R721 B.n219 B.n218 163.367
R722 B.n223 B.n222 163.367
R723 B.n227 B.n226 163.367
R724 B.n231 B.n230 163.367
R725 B.n235 B.n234 163.367
R726 B.n239 B.n238 163.367
R727 B.n243 B.n242 163.367
R728 B.n247 B.n246 163.367
R729 B.n249 B.n88 163.367
R730 B.n501 B.n296 98.2473
R731 B.n616 B.n615 98.2473
R732 B.n343 B.t21 96.8517
R733 B.n89 B.t13 96.8517
R734 B.n340 B.t18 96.8399
R735 B.n91 B.t10 96.8399
R736 B.n344 B.t20 74.3547
R737 B.n90 B.t14 74.3547
R738 B.n341 B.t17 74.343
R739 B.n92 B.t11 74.343
R740 B.n500 B.n499 71.676
R741 B.n494 B.n300 71.676
R742 B.n491 B.n301 71.676
R743 B.n487 B.n302 71.676
R744 B.n483 B.n303 71.676
R745 B.n479 B.n304 71.676
R746 B.n475 B.n305 71.676
R747 B.n471 B.n306 71.676
R748 B.n467 B.n307 71.676
R749 B.n463 B.n308 71.676
R750 B.n459 B.n309 71.676
R751 B.n455 B.n310 71.676
R752 B.n451 B.n311 71.676
R753 B.n447 B.n312 71.676
R754 B.n443 B.n313 71.676
R755 B.n439 B.n314 71.676
R756 B.n435 B.n315 71.676
R757 B.n431 B.n316 71.676
R758 B.n427 B.n317 71.676
R759 B.n423 B.n318 71.676
R760 B.n419 B.n319 71.676
R761 B.n415 B.n320 71.676
R762 B.n411 B.n321 71.676
R763 B.n407 B.n322 71.676
R764 B.n403 B.n323 71.676
R765 B.n399 B.n324 71.676
R766 B.n395 B.n325 71.676
R767 B.n391 B.n326 71.676
R768 B.n387 B.n327 71.676
R769 B.n383 B.n328 71.676
R770 B.n379 B.n329 71.676
R771 B.n375 B.n330 71.676
R772 B.n371 B.n331 71.676
R773 B.n367 B.n332 71.676
R774 B.n363 B.n333 71.676
R775 B.n359 B.n334 71.676
R776 B.n355 B.n335 71.676
R777 B.n351 B.n336 71.676
R778 B.n347 B.n337 71.676
R779 B.n93 B.n49 71.676
R780 B.n97 B.n50 71.676
R781 B.n101 B.n51 71.676
R782 B.n105 B.n52 71.676
R783 B.n109 B.n53 71.676
R784 B.n113 B.n54 71.676
R785 B.n117 B.n55 71.676
R786 B.n121 B.n56 71.676
R787 B.n125 B.n57 71.676
R788 B.n129 B.n58 71.676
R789 B.n133 B.n59 71.676
R790 B.n137 B.n60 71.676
R791 B.n141 B.n61 71.676
R792 B.n145 B.n62 71.676
R793 B.n149 B.n63 71.676
R794 B.n153 B.n64 71.676
R795 B.n157 B.n65 71.676
R796 B.n161 B.n66 71.676
R797 B.n166 B.n67 71.676
R798 B.n170 B.n68 71.676
R799 B.n174 B.n69 71.676
R800 B.n178 B.n70 71.676
R801 B.n182 B.n71 71.676
R802 B.n187 B.n72 71.676
R803 B.n191 B.n73 71.676
R804 B.n195 B.n74 71.676
R805 B.n199 B.n75 71.676
R806 B.n203 B.n76 71.676
R807 B.n207 B.n77 71.676
R808 B.n211 B.n78 71.676
R809 B.n215 B.n79 71.676
R810 B.n219 B.n80 71.676
R811 B.n223 B.n81 71.676
R812 B.n227 B.n82 71.676
R813 B.n231 B.n83 71.676
R814 B.n235 B.n84 71.676
R815 B.n239 B.n85 71.676
R816 B.n243 B.n86 71.676
R817 B.n247 B.n87 71.676
R818 B.n614 B.n88 71.676
R819 B.n614 B.n613 71.676
R820 B.n249 B.n87 71.676
R821 B.n246 B.n86 71.676
R822 B.n242 B.n85 71.676
R823 B.n238 B.n84 71.676
R824 B.n234 B.n83 71.676
R825 B.n230 B.n82 71.676
R826 B.n226 B.n81 71.676
R827 B.n222 B.n80 71.676
R828 B.n218 B.n79 71.676
R829 B.n214 B.n78 71.676
R830 B.n210 B.n77 71.676
R831 B.n206 B.n76 71.676
R832 B.n202 B.n75 71.676
R833 B.n198 B.n74 71.676
R834 B.n194 B.n73 71.676
R835 B.n190 B.n72 71.676
R836 B.n186 B.n71 71.676
R837 B.n181 B.n70 71.676
R838 B.n177 B.n69 71.676
R839 B.n173 B.n68 71.676
R840 B.n169 B.n67 71.676
R841 B.n165 B.n66 71.676
R842 B.n160 B.n65 71.676
R843 B.n156 B.n64 71.676
R844 B.n152 B.n63 71.676
R845 B.n148 B.n62 71.676
R846 B.n144 B.n61 71.676
R847 B.n140 B.n60 71.676
R848 B.n136 B.n59 71.676
R849 B.n132 B.n58 71.676
R850 B.n128 B.n57 71.676
R851 B.n124 B.n56 71.676
R852 B.n120 B.n55 71.676
R853 B.n116 B.n54 71.676
R854 B.n112 B.n53 71.676
R855 B.n108 B.n52 71.676
R856 B.n104 B.n51 71.676
R857 B.n100 B.n50 71.676
R858 B.n96 B.n49 71.676
R859 B.n500 B.n339 71.676
R860 B.n492 B.n300 71.676
R861 B.n488 B.n301 71.676
R862 B.n484 B.n302 71.676
R863 B.n480 B.n303 71.676
R864 B.n476 B.n304 71.676
R865 B.n472 B.n305 71.676
R866 B.n468 B.n306 71.676
R867 B.n464 B.n307 71.676
R868 B.n460 B.n308 71.676
R869 B.n456 B.n309 71.676
R870 B.n452 B.n310 71.676
R871 B.n448 B.n311 71.676
R872 B.n444 B.n312 71.676
R873 B.n440 B.n313 71.676
R874 B.n436 B.n314 71.676
R875 B.n432 B.n315 71.676
R876 B.n428 B.n316 71.676
R877 B.n424 B.n317 71.676
R878 B.n420 B.n318 71.676
R879 B.n416 B.n319 71.676
R880 B.n412 B.n320 71.676
R881 B.n408 B.n321 71.676
R882 B.n404 B.n322 71.676
R883 B.n400 B.n323 71.676
R884 B.n396 B.n324 71.676
R885 B.n392 B.n325 71.676
R886 B.n388 B.n326 71.676
R887 B.n384 B.n327 71.676
R888 B.n380 B.n328 71.676
R889 B.n376 B.n329 71.676
R890 B.n372 B.n330 71.676
R891 B.n368 B.n331 71.676
R892 B.n364 B.n332 71.676
R893 B.n360 B.n333 71.676
R894 B.n356 B.n334 71.676
R895 B.n352 B.n335 71.676
R896 B.n348 B.n336 71.676
R897 B.n337 B.n299 71.676
R898 B.n345 B.n344 59.5399
R899 B.n342 B.n341 59.5399
R900 B.n163 B.n92 59.5399
R901 B.n184 B.n90 59.5399
R902 B.n507 B.n296 49.4878
R903 B.n507 B.n291 49.4878
R904 B.n513 B.n291 49.4878
R905 B.n513 B.n292 49.4878
R906 B.n519 B.n284 49.4878
R907 B.n525 B.n284 49.4878
R908 B.n525 B.n280 49.4878
R909 B.n531 B.n280 49.4878
R910 B.n531 B.n276 49.4878
R911 B.n537 B.n276 49.4878
R912 B.n544 B.n272 49.4878
R913 B.n544 B.n543 49.4878
R914 B.n550 B.n265 49.4878
R915 B.n557 B.n265 49.4878
R916 B.n557 B.n556 49.4878
R917 B.n563 B.n258 49.4878
R918 B.n570 B.n258 49.4878
R919 B.n576 B.n254 49.4878
R920 B.n576 B.n4 49.4878
R921 B.n665 B.n4 49.4878
R922 B.n665 B.n664 49.4878
R923 B.n664 B.n663 49.4878
R924 B.n663 B.n8 49.4878
R925 B.n657 B.n656 49.4878
R926 B.n656 B.n655 49.4878
R927 B.n649 B.n18 49.4878
R928 B.n649 B.n648 49.4878
R929 B.n648 B.n647 49.4878
R930 B.n641 B.n25 49.4878
R931 B.n641 B.n640 49.4878
R932 B.n639 B.n29 49.4878
R933 B.n633 B.n29 49.4878
R934 B.n633 B.n632 49.4878
R935 B.n632 B.n631 49.4878
R936 B.n631 B.n36 49.4878
R937 B.n625 B.n36 49.4878
R938 B.n624 B.n623 49.4878
R939 B.n623 B.n43 49.4878
R940 B.n617 B.n43 49.4878
R941 B.n617 B.n616 49.4878
R942 B.n543 B.t0 42.938
R943 B.n25 B.t5 42.938
R944 B.n292 B.t16 41.4825
R945 B.t9 B.n624 41.4825
R946 B.n563 B.t2 35.6604
R947 B.n655 B.t3 35.6604
R948 B.n612 B.n611 34.8103
R949 B.n94 B.n45 34.8103
R950 B.n504 B.n503 34.8103
R951 B.n498 B.n294 34.8103
R952 B.n570 B.t6 34.2049
R953 B.n657 B.t1 34.2049
R954 B.t7 B.n272 26.9274
R955 B.n640 B.t4 26.9274
R956 B.n537 B.t7 22.5609
R957 B.t4 B.n639 22.5609
R958 B.n344 B.n343 22.4975
R959 B.n341 B.n340 22.4975
R960 B.n92 B.n91 22.4975
R961 B.n90 B.n89 22.4975
R962 B B.n667 18.0485
R963 B.t6 B.n254 15.2833
R964 B.t1 B.n8 15.2833
R965 B.n556 B.t2 13.8278
R966 B.n18 B.t3 13.8278
R967 B.n95 B.n94 10.6151
R968 B.n98 B.n95 10.6151
R969 B.n99 B.n98 10.6151
R970 B.n102 B.n99 10.6151
R971 B.n103 B.n102 10.6151
R972 B.n106 B.n103 10.6151
R973 B.n107 B.n106 10.6151
R974 B.n110 B.n107 10.6151
R975 B.n111 B.n110 10.6151
R976 B.n114 B.n111 10.6151
R977 B.n115 B.n114 10.6151
R978 B.n118 B.n115 10.6151
R979 B.n119 B.n118 10.6151
R980 B.n122 B.n119 10.6151
R981 B.n123 B.n122 10.6151
R982 B.n126 B.n123 10.6151
R983 B.n127 B.n126 10.6151
R984 B.n130 B.n127 10.6151
R985 B.n131 B.n130 10.6151
R986 B.n134 B.n131 10.6151
R987 B.n135 B.n134 10.6151
R988 B.n138 B.n135 10.6151
R989 B.n139 B.n138 10.6151
R990 B.n142 B.n139 10.6151
R991 B.n143 B.n142 10.6151
R992 B.n146 B.n143 10.6151
R993 B.n147 B.n146 10.6151
R994 B.n150 B.n147 10.6151
R995 B.n151 B.n150 10.6151
R996 B.n154 B.n151 10.6151
R997 B.n155 B.n154 10.6151
R998 B.n158 B.n155 10.6151
R999 B.n159 B.n158 10.6151
R1000 B.n162 B.n159 10.6151
R1001 B.n167 B.n164 10.6151
R1002 B.n168 B.n167 10.6151
R1003 B.n171 B.n168 10.6151
R1004 B.n172 B.n171 10.6151
R1005 B.n175 B.n172 10.6151
R1006 B.n176 B.n175 10.6151
R1007 B.n179 B.n176 10.6151
R1008 B.n180 B.n179 10.6151
R1009 B.n183 B.n180 10.6151
R1010 B.n188 B.n185 10.6151
R1011 B.n189 B.n188 10.6151
R1012 B.n192 B.n189 10.6151
R1013 B.n193 B.n192 10.6151
R1014 B.n196 B.n193 10.6151
R1015 B.n197 B.n196 10.6151
R1016 B.n200 B.n197 10.6151
R1017 B.n201 B.n200 10.6151
R1018 B.n204 B.n201 10.6151
R1019 B.n205 B.n204 10.6151
R1020 B.n208 B.n205 10.6151
R1021 B.n209 B.n208 10.6151
R1022 B.n212 B.n209 10.6151
R1023 B.n213 B.n212 10.6151
R1024 B.n216 B.n213 10.6151
R1025 B.n217 B.n216 10.6151
R1026 B.n220 B.n217 10.6151
R1027 B.n221 B.n220 10.6151
R1028 B.n224 B.n221 10.6151
R1029 B.n225 B.n224 10.6151
R1030 B.n228 B.n225 10.6151
R1031 B.n229 B.n228 10.6151
R1032 B.n232 B.n229 10.6151
R1033 B.n233 B.n232 10.6151
R1034 B.n236 B.n233 10.6151
R1035 B.n237 B.n236 10.6151
R1036 B.n240 B.n237 10.6151
R1037 B.n241 B.n240 10.6151
R1038 B.n244 B.n241 10.6151
R1039 B.n245 B.n244 10.6151
R1040 B.n248 B.n245 10.6151
R1041 B.n250 B.n248 10.6151
R1042 B.n251 B.n250 10.6151
R1043 B.n612 B.n251 10.6151
R1044 B.n505 B.n504 10.6151
R1045 B.n505 B.n289 10.6151
R1046 B.n515 B.n289 10.6151
R1047 B.n516 B.n515 10.6151
R1048 B.n517 B.n516 10.6151
R1049 B.n517 B.n282 10.6151
R1050 B.n527 B.n282 10.6151
R1051 B.n528 B.n527 10.6151
R1052 B.n529 B.n528 10.6151
R1053 B.n529 B.n274 10.6151
R1054 B.n539 B.n274 10.6151
R1055 B.n540 B.n539 10.6151
R1056 B.n541 B.n540 10.6151
R1057 B.n541 B.n267 10.6151
R1058 B.n552 B.n267 10.6151
R1059 B.n553 B.n552 10.6151
R1060 B.n554 B.n553 10.6151
R1061 B.n554 B.n260 10.6151
R1062 B.n565 B.n260 10.6151
R1063 B.n566 B.n565 10.6151
R1064 B.n568 B.n566 10.6151
R1065 B.n568 B.n567 10.6151
R1066 B.n567 B.n252 10.6151
R1067 B.n579 B.n252 10.6151
R1068 B.n580 B.n579 10.6151
R1069 B.n581 B.n580 10.6151
R1070 B.n582 B.n581 10.6151
R1071 B.n584 B.n582 10.6151
R1072 B.n585 B.n584 10.6151
R1073 B.n586 B.n585 10.6151
R1074 B.n587 B.n586 10.6151
R1075 B.n589 B.n587 10.6151
R1076 B.n590 B.n589 10.6151
R1077 B.n591 B.n590 10.6151
R1078 B.n592 B.n591 10.6151
R1079 B.n594 B.n592 10.6151
R1080 B.n595 B.n594 10.6151
R1081 B.n596 B.n595 10.6151
R1082 B.n597 B.n596 10.6151
R1083 B.n599 B.n597 10.6151
R1084 B.n600 B.n599 10.6151
R1085 B.n601 B.n600 10.6151
R1086 B.n602 B.n601 10.6151
R1087 B.n604 B.n602 10.6151
R1088 B.n605 B.n604 10.6151
R1089 B.n606 B.n605 10.6151
R1090 B.n607 B.n606 10.6151
R1091 B.n609 B.n607 10.6151
R1092 B.n610 B.n609 10.6151
R1093 B.n611 B.n610 10.6151
R1094 B.n498 B.n497 10.6151
R1095 B.n497 B.n496 10.6151
R1096 B.n496 B.n495 10.6151
R1097 B.n495 B.n493 10.6151
R1098 B.n493 B.n490 10.6151
R1099 B.n490 B.n489 10.6151
R1100 B.n489 B.n486 10.6151
R1101 B.n486 B.n485 10.6151
R1102 B.n485 B.n482 10.6151
R1103 B.n482 B.n481 10.6151
R1104 B.n481 B.n478 10.6151
R1105 B.n478 B.n477 10.6151
R1106 B.n477 B.n474 10.6151
R1107 B.n474 B.n473 10.6151
R1108 B.n473 B.n470 10.6151
R1109 B.n470 B.n469 10.6151
R1110 B.n469 B.n466 10.6151
R1111 B.n466 B.n465 10.6151
R1112 B.n465 B.n462 10.6151
R1113 B.n462 B.n461 10.6151
R1114 B.n461 B.n458 10.6151
R1115 B.n458 B.n457 10.6151
R1116 B.n457 B.n454 10.6151
R1117 B.n454 B.n453 10.6151
R1118 B.n453 B.n450 10.6151
R1119 B.n450 B.n449 10.6151
R1120 B.n449 B.n446 10.6151
R1121 B.n446 B.n445 10.6151
R1122 B.n445 B.n442 10.6151
R1123 B.n442 B.n441 10.6151
R1124 B.n441 B.n438 10.6151
R1125 B.n438 B.n437 10.6151
R1126 B.n437 B.n434 10.6151
R1127 B.n434 B.n433 10.6151
R1128 B.n430 B.n429 10.6151
R1129 B.n429 B.n426 10.6151
R1130 B.n426 B.n425 10.6151
R1131 B.n425 B.n422 10.6151
R1132 B.n422 B.n421 10.6151
R1133 B.n421 B.n418 10.6151
R1134 B.n418 B.n417 10.6151
R1135 B.n417 B.n414 10.6151
R1136 B.n414 B.n413 10.6151
R1137 B.n410 B.n409 10.6151
R1138 B.n409 B.n406 10.6151
R1139 B.n406 B.n405 10.6151
R1140 B.n405 B.n402 10.6151
R1141 B.n402 B.n401 10.6151
R1142 B.n401 B.n398 10.6151
R1143 B.n398 B.n397 10.6151
R1144 B.n397 B.n394 10.6151
R1145 B.n394 B.n393 10.6151
R1146 B.n393 B.n390 10.6151
R1147 B.n390 B.n389 10.6151
R1148 B.n389 B.n386 10.6151
R1149 B.n386 B.n385 10.6151
R1150 B.n385 B.n382 10.6151
R1151 B.n382 B.n381 10.6151
R1152 B.n381 B.n378 10.6151
R1153 B.n378 B.n377 10.6151
R1154 B.n377 B.n374 10.6151
R1155 B.n374 B.n373 10.6151
R1156 B.n373 B.n370 10.6151
R1157 B.n370 B.n369 10.6151
R1158 B.n369 B.n366 10.6151
R1159 B.n366 B.n365 10.6151
R1160 B.n365 B.n362 10.6151
R1161 B.n362 B.n361 10.6151
R1162 B.n361 B.n358 10.6151
R1163 B.n358 B.n357 10.6151
R1164 B.n357 B.n354 10.6151
R1165 B.n354 B.n353 10.6151
R1166 B.n353 B.n350 10.6151
R1167 B.n350 B.n349 10.6151
R1168 B.n349 B.n346 10.6151
R1169 B.n346 B.n298 10.6151
R1170 B.n503 B.n298 10.6151
R1171 B.n509 B.n294 10.6151
R1172 B.n510 B.n509 10.6151
R1173 B.n511 B.n510 10.6151
R1174 B.n511 B.n286 10.6151
R1175 B.n521 B.n286 10.6151
R1176 B.n522 B.n521 10.6151
R1177 B.n523 B.n522 10.6151
R1178 B.n523 B.n278 10.6151
R1179 B.n533 B.n278 10.6151
R1180 B.n534 B.n533 10.6151
R1181 B.n535 B.n534 10.6151
R1182 B.n535 B.n270 10.6151
R1183 B.n546 B.n270 10.6151
R1184 B.n547 B.n546 10.6151
R1185 B.n548 B.n547 10.6151
R1186 B.n548 B.n263 10.6151
R1187 B.n559 B.n263 10.6151
R1188 B.n560 B.n559 10.6151
R1189 B.n561 B.n560 10.6151
R1190 B.n561 B.n256 10.6151
R1191 B.n572 B.n256 10.6151
R1192 B.n573 B.n572 10.6151
R1193 B.n574 B.n573 10.6151
R1194 B.n574 B.n0 10.6151
R1195 B.n661 B.n1 10.6151
R1196 B.n661 B.n660 10.6151
R1197 B.n660 B.n659 10.6151
R1198 B.n659 B.n10 10.6151
R1199 B.n653 B.n10 10.6151
R1200 B.n653 B.n652 10.6151
R1201 B.n652 B.n651 10.6151
R1202 B.n651 B.n16 10.6151
R1203 B.n645 B.n16 10.6151
R1204 B.n645 B.n644 10.6151
R1205 B.n644 B.n643 10.6151
R1206 B.n643 B.n23 10.6151
R1207 B.n637 B.n23 10.6151
R1208 B.n637 B.n636 10.6151
R1209 B.n636 B.n635 10.6151
R1210 B.n635 B.n31 10.6151
R1211 B.n629 B.n31 10.6151
R1212 B.n629 B.n628 10.6151
R1213 B.n628 B.n627 10.6151
R1214 B.n627 B.n38 10.6151
R1215 B.n621 B.n38 10.6151
R1216 B.n621 B.n620 10.6151
R1217 B.n620 B.n619 10.6151
R1218 B.n619 B.n45 10.6151
R1219 B.n163 B.n162 9.36635
R1220 B.n185 B.n184 9.36635
R1221 B.n433 B.n342 9.36635
R1222 B.n410 B.n345 9.36635
R1223 B.n519 B.t16 8.00579
R1224 B.n625 B.t9 8.00579
R1225 B.n550 B.t0 6.55029
R1226 B.n647 B.t5 6.55029
R1227 B.n667 B.n0 2.81026
R1228 B.n667 B.n1 2.81026
R1229 B.n164 B.n163 1.24928
R1230 B.n184 B.n183 1.24928
R1231 B.n430 B.n342 1.24928
R1232 B.n413 B.n345 1.24928
R1233 VN.n3 VN.t5 352.868
R1234 VN.n16 VN.t4 352.868
R1235 VN.n11 VN.t1 333.046
R1236 VN.n24 VN.t7 333.046
R1237 VN.n4 VN.t0 285.716
R1238 VN.n1 VN.t2 285.716
R1239 VN.n17 VN.t3 285.716
R1240 VN.n14 VN.t6 285.716
R1241 VN.n12 VN.n11 161.3
R1242 VN.n25 VN.n24 161.3
R1243 VN.n23 VN.n13 161.3
R1244 VN.n22 VN.n21 161.3
R1245 VN.n20 VN.n19 161.3
R1246 VN.n18 VN.n15 161.3
R1247 VN.n10 VN.n0 161.3
R1248 VN.n9 VN.n8 161.3
R1249 VN.n7 VN.n6 161.3
R1250 VN.n5 VN.n2 161.3
R1251 VN.n6 VN.n5 56.5617
R1252 VN.n19 VN.n18 56.5617
R1253 VN.n10 VN.n9 49.296
R1254 VN.n23 VN.n22 49.296
R1255 VN.n16 VN.n15 43.0963
R1256 VN.n3 VN.n2 43.0963
R1257 VN VN.n25 41.3357
R1258 VN.n4 VN.n3 38.2995
R1259 VN.n17 VN.n16 38.2995
R1260 VN.n5 VN.n4 16.2311
R1261 VN.n6 VN.n1 16.2311
R1262 VN.n18 VN.n17 16.2311
R1263 VN.n19 VN.n14 16.2311
R1264 VN.n11 VN.n10 10.955
R1265 VN.n24 VN.n23 10.955
R1266 VN.n9 VN.n1 8.36172
R1267 VN.n22 VN.n14 8.36172
R1268 VN.n25 VN.n13 0.189894
R1269 VN.n21 VN.n13 0.189894
R1270 VN.n21 VN.n20 0.189894
R1271 VN.n20 VN.n15 0.189894
R1272 VN.n7 VN.n2 0.189894
R1273 VN.n8 VN.n7 0.189894
R1274 VN.n8 VN.n0 0.189894
R1275 VN.n12 VN.n0 0.189894
R1276 VN VN.n12 0.0516364
R1277 VDD2.n2 VDD2.n1 61.3899
R1278 VDD2.n2 VDD2.n0 61.3899
R1279 VDD2 VDD2.n5 61.3872
R1280 VDD2.n4 VDD2.n3 60.9454
R1281 VDD2.n4 VDD2.n2 36.6981
R1282 VDD2.n5 VDD2.t4 2.0127
R1283 VDD2.n5 VDD2.t3 2.0127
R1284 VDD2.n3 VDD2.t0 2.0127
R1285 VDD2.n3 VDD2.t1 2.0127
R1286 VDD2.n1 VDD2.t5 2.0127
R1287 VDD2.n1 VDD2.t6 2.0127
R1288 VDD2.n0 VDD2.t2 2.0127
R1289 VDD2.n0 VDD2.t7 2.0127
R1290 VDD2 VDD2.n4 0.55869
C0 VP VDD1 5.16782f
C1 VTAIL VDD2 8.8903f
C2 VN VDD2 4.98552f
C3 VTAIL VN 4.87559f
C4 VDD2 VP 0.331421f
C5 VTAIL VP 4.88969f
C6 VDD2 VDD1 0.889127f
C7 VN VP 5.09548f
C8 VTAIL VDD1 8.847751f
C9 VN VDD1 0.148625f
C10 VDD2 B 3.454609f
C11 VDD1 B 3.701661f
C12 VTAIL B 7.837358f
C13 VN B 8.776269f
C14 VP B 6.993078f
C15 VDD2.t2 B 0.206489f
C16 VDD2.t7 B 0.206489f
C17 VDD2.n0 B 1.80804f
C18 VDD2.t5 B 0.206489f
C19 VDD2.t6 B 0.206489f
C20 VDD2.n1 B 1.80804f
C21 VDD2.n2 B 2.2646f
C22 VDD2.t0 B 0.206489f
C23 VDD2.t1 B 0.206489f
C24 VDD2.n3 B 1.80542f
C25 VDD2.n4 B 2.31003f
C26 VDD2.t4 B 0.206489f
C27 VDD2.t3 B 0.206489f
C28 VDD2.n5 B 1.80801f
C29 VN.n0 B 0.041567f
C30 VN.t2 B 0.91916f
C31 VN.n1 B 0.355182f
C32 VN.n2 B 0.173351f
C33 VN.t0 B 0.91916f
C34 VN.t5 B 0.994408f
C35 VN.n3 B 0.397643f
C36 VN.n4 B 0.396688f
C37 VN.n5 B 0.047485f
C38 VN.n6 B 0.047485f
C39 VN.n7 B 0.041567f
C40 VN.n8 B 0.041567f
C41 VN.n9 B 0.051585f
C42 VN.n10 B 0.015588f
C43 VN.t1 B 0.971692f
C44 VN.n11 B 0.39383f
C45 VN.n12 B 0.032212f
C46 VN.n13 B 0.041567f
C47 VN.t6 B 0.91916f
C48 VN.n14 B 0.355182f
C49 VN.n15 B 0.173351f
C50 VN.t3 B 0.91916f
C51 VN.t4 B 0.994408f
C52 VN.n16 B 0.397643f
C53 VN.n17 B 0.396688f
C54 VN.n18 B 0.047485f
C55 VN.n19 B 0.047485f
C56 VN.n20 B 0.041567f
C57 VN.n21 B 0.041567f
C58 VN.n22 B 0.051585f
C59 VN.n23 B 0.015588f
C60 VN.t7 B 0.971692f
C61 VN.n24 B 0.39383f
C62 VN.n25 B 1.67186f
C63 VDD1.t6 B 0.206517f
C64 VDD1.t7 B 0.206517f
C65 VDD1.n0 B 1.80903f
C66 VDD1.t4 B 0.206517f
C67 VDD1.t2 B 0.206517f
C68 VDD1.n1 B 1.80828f
C69 VDD1.t1 B 0.206517f
C70 VDD1.t3 B 0.206517f
C71 VDD1.n2 B 1.80828f
C72 VDD1.n3 B 2.32159f
C73 VDD1.t0 B 0.206517f
C74 VDD1.t5 B 0.206517f
C75 VDD1.n4 B 1.80566f
C76 VDD1.n5 B 2.34181f
C77 VTAIL.t3 B 0.1563f
C78 VTAIL.t5 B 0.1563f
C79 VTAIL.n0 B 1.30331f
C80 VTAIL.n1 B 0.27627f
C81 VTAIL.t1 B 1.66117f
C82 VTAIL.n2 B 0.371338f
C83 VTAIL.t11 B 1.66117f
C84 VTAIL.n3 B 0.371338f
C85 VTAIL.t14 B 0.1563f
C86 VTAIL.t15 B 0.1563f
C87 VTAIL.n4 B 1.30331f
C88 VTAIL.n5 B 0.33727f
C89 VTAIL.t13 B 1.66117f
C90 VTAIL.n6 B 1.22814f
C91 VTAIL.t7 B 1.66118f
C92 VTAIL.n7 B 1.22813f
C93 VTAIL.t0 B 0.1563f
C94 VTAIL.t2 B 0.1563f
C95 VTAIL.n8 B 1.30332f
C96 VTAIL.n9 B 0.337263f
C97 VTAIL.t6 B 1.66118f
C98 VTAIL.n10 B 0.371332f
C99 VTAIL.t9 B 1.66118f
C100 VTAIL.n11 B 0.371332f
C101 VTAIL.t12 B 0.1563f
C102 VTAIL.t10 B 0.1563f
C103 VTAIL.n12 B 1.30332f
C104 VTAIL.n13 B 0.337263f
C105 VTAIL.t8 B 1.66118f
C106 VTAIL.n14 B 1.22813f
C107 VTAIL.t4 B 1.66117f
C108 VTAIL.n15 B 1.22437f
C109 VP.n0 B 0.042285f
C110 VP.t6 B 0.935058f
C111 VP.n1 B 0.361326f
C112 VP.n2 B 0.042285f
C113 VP.t5 B 0.935058f
C114 VP.n3 B 0.015857f
C115 VP.n4 B 0.042285f
C116 VP.t2 B 0.988499f
C117 VP.t7 B 0.935058f
C118 VP.n5 B 0.361326f
C119 VP.n6 B 0.176349f
C120 VP.t0 B 0.935058f
C121 VP.t1 B 1.01161f
C122 VP.n7 B 0.40452f
C123 VP.n8 B 0.403549f
C124 VP.n9 B 0.048307f
C125 VP.n10 B 0.048307f
C126 VP.n11 B 0.042285f
C127 VP.n12 B 0.042285f
C128 VP.n13 B 0.052477f
C129 VP.n14 B 0.015857f
C130 VP.n15 B 0.400642f
C131 VP.n16 B 1.67298f
C132 VP.t3 B 0.988499f
C133 VP.n17 B 0.400642f
C134 VP.n18 B 1.7102f
C135 VP.n19 B 0.042285f
C136 VP.n20 B 0.042285f
C137 VP.n21 B 0.052477f
C138 VP.n22 B 0.361326f
C139 VP.n23 B 0.048307f
C140 VP.n24 B 0.048307f
C141 VP.n25 B 0.042285f
C142 VP.n26 B 0.042285f
C143 VP.n27 B 0.052477f
C144 VP.n28 B 0.015857f
C145 VP.t4 B 0.988499f
C146 VP.n29 B 0.400642f
C147 VP.n30 B 0.03277f
.ends

