* NGSPICE file created from diff_pair_sample_1028.ext - technology: sky130A

.subckt diff_pair_sample_1028 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t3 VN.t0 VTAIL.t4 B.t1 sky130_fd_pr__nfet_01v8 ad=1.584 pd=9.93 as=3.744 ps=19.98 w=9.6 l=1.4
X1 VTAIL.t5 VN.t1 VDD2.t2 B.t0 sky130_fd_pr__nfet_01v8 ad=3.744 pd=19.98 as=1.584 ps=9.93 w=9.6 l=1.4
X2 B.t17 B.t15 B.t16 B.t5 sky130_fd_pr__nfet_01v8 ad=3.744 pd=19.98 as=0 ps=0 w=9.6 l=1.4
X3 VTAIL.t0 VP.t0 VDD1.t3 B.t0 sky130_fd_pr__nfet_01v8 ad=3.744 pd=19.98 as=1.584 ps=9.93 w=9.6 l=1.4
X4 VDD1.t2 VP.t1 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=1.584 pd=9.93 as=3.744 ps=19.98 w=9.6 l=1.4
X5 B.t14 B.t12 B.t13 B.t9 sky130_fd_pr__nfet_01v8 ad=3.744 pd=19.98 as=0 ps=0 w=9.6 l=1.4
X6 VTAIL.t2 VP.t2 VDD1.t1 B.t2 sky130_fd_pr__nfet_01v8 ad=3.744 pd=19.98 as=1.584 ps=9.93 w=9.6 l=1.4
X7 VDD1.t0 VP.t3 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=1.584 pd=9.93 as=3.744 ps=19.98 w=9.6 l=1.4
X8 VDD2.t1 VN.t2 VTAIL.t7 B.t3 sky130_fd_pr__nfet_01v8 ad=1.584 pd=9.93 as=3.744 ps=19.98 w=9.6 l=1.4
X9 VTAIL.t6 VN.t3 VDD2.t0 B.t2 sky130_fd_pr__nfet_01v8 ad=3.744 pd=19.98 as=1.584 ps=9.93 w=9.6 l=1.4
X10 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=3.744 pd=19.98 as=0 ps=0 w=9.6 l=1.4
X11 B.t7 B.t4 B.t6 B.t5 sky130_fd_pr__nfet_01v8 ad=3.744 pd=19.98 as=0 ps=0 w=9.6 l=1.4
R0 VN.n0 VN.t1 200.209
R1 VN.n1 VN.t2 200.209
R2 VN.n0 VN.t0 199.901
R3 VN.n1 VN.t3 199.901
R4 VN VN.n1 54.4041
R5 VN VN.n0 13.4003
R6 VTAIL.n5 VTAIL.t0 48.1958
R7 VTAIL.n4 VTAIL.t7 48.1958
R8 VTAIL.n3 VTAIL.t6 48.1958
R9 VTAIL.n7 VTAIL.t4 48.1957
R10 VTAIL.n0 VTAIL.t5 48.1957
R11 VTAIL.n1 VTAIL.t3 48.1957
R12 VTAIL.n2 VTAIL.t2 48.1957
R13 VTAIL.n6 VTAIL.t1 48.1957
R14 VTAIL.n7 VTAIL.n6 22.1341
R15 VTAIL.n3 VTAIL.n2 22.1341
R16 VTAIL.n4 VTAIL.n3 1.49188
R17 VTAIL.n6 VTAIL.n5 1.49188
R18 VTAIL.n2 VTAIL.n1 1.49188
R19 VTAIL VTAIL.n0 0.804379
R20 VTAIL VTAIL.n7 0.688
R21 VTAIL.n5 VTAIL.n4 0.470328
R22 VTAIL.n1 VTAIL.n0 0.470328
R23 VDD2.n2 VDD2.n0 99.2767
R24 VDD2.n2 VDD2.n1 62.812
R25 VDD2.n1 VDD2.t0 2.063
R26 VDD2.n1 VDD2.t1 2.063
R27 VDD2.n0 VDD2.t2 2.063
R28 VDD2.n0 VDD2.t3 2.063
R29 VDD2 VDD2.n2 0.0586897
R30 B.n593 B.n592 585
R31 B.n594 B.n593 585
R32 B.n243 B.n85 585
R33 B.n242 B.n241 585
R34 B.n240 B.n239 585
R35 B.n238 B.n237 585
R36 B.n236 B.n235 585
R37 B.n234 B.n233 585
R38 B.n232 B.n231 585
R39 B.n230 B.n229 585
R40 B.n228 B.n227 585
R41 B.n226 B.n225 585
R42 B.n224 B.n223 585
R43 B.n222 B.n221 585
R44 B.n220 B.n219 585
R45 B.n218 B.n217 585
R46 B.n216 B.n215 585
R47 B.n214 B.n213 585
R48 B.n212 B.n211 585
R49 B.n210 B.n209 585
R50 B.n208 B.n207 585
R51 B.n206 B.n205 585
R52 B.n204 B.n203 585
R53 B.n202 B.n201 585
R54 B.n200 B.n199 585
R55 B.n198 B.n197 585
R56 B.n196 B.n195 585
R57 B.n194 B.n193 585
R58 B.n192 B.n191 585
R59 B.n190 B.n189 585
R60 B.n188 B.n187 585
R61 B.n186 B.n185 585
R62 B.n184 B.n183 585
R63 B.n182 B.n181 585
R64 B.n180 B.n179 585
R65 B.n178 B.n177 585
R66 B.n176 B.n175 585
R67 B.n174 B.n173 585
R68 B.n172 B.n171 585
R69 B.n170 B.n169 585
R70 B.n168 B.n167 585
R71 B.n166 B.n165 585
R72 B.n164 B.n163 585
R73 B.n162 B.n161 585
R74 B.n160 B.n159 585
R75 B.n157 B.n156 585
R76 B.n155 B.n154 585
R77 B.n153 B.n152 585
R78 B.n151 B.n150 585
R79 B.n149 B.n148 585
R80 B.n147 B.n146 585
R81 B.n145 B.n144 585
R82 B.n143 B.n142 585
R83 B.n141 B.n140 585
R84 B.n139 B.n138 585
R85 B.n137 B.n136 585
R86 B.n135 B.n134 585
R87 B.n133 B.n132 585
R88 B.n131 B.n130 585
R89 B.n129 B.n128 585
R90 B.n127 B.n126 585
R91 B.n125 B.n124 585
R92 B.n123 B.n122 585
R93 B.n121 B.n120 585
R94 B.n119 B.n118 585
R95 B.n117 B.n116 585
R96 B.n115 B.n114 585
R97 B.n113 B.n112 585
R98 B.n111 B.n110 585
R99 B.n109 B.n108 585
R100 B.n107 B.n106 585
R101 B.n105 B.n104 585
R102 B.n103 B.n102 585
R103 B.n101 B.n100 585
R104 B.n99 B.n98 585
R105 B.n97 B.n96 585
R106 B.n95 B.n94 585
R107 B.n93 B.n92 585
R108 B.n46 B.n45 585
R109 B.n597 B.n596 585
R110 B.n591 B.n86 585
R111 B.n86 B.n43 585
R112 B.n590 B.n42 585
R113 B.n601 B.n42 585
R114 B.n589 B.n41 585
R115 B.n602 B.n41 585
R116 B.n588 B.n40 585
R117 B.n603 B.n40 585
R118 B.n587 B.n586 585
R119 B.n586 B.n36 585
R120 B.n585 B.n35 585
R121 B.n609 B.n35 585
R122 B.n584 B.n34 585
R123 B.n610 B.n34 585
R124 B.n583 B.n33 585
R125 B.n611 B.n33 585
R126 B.n582 B.n581 585
R127 B.n581 B.n29 585
R128 B.n580 B.n28 585
R129 B.n617 B.n28 585
R130 B.n579 B.n27 585
R131 B.n618 B.n27 585
R132 B.n578 B.n26 585
R133 B.n619 B.n26 585
R134 B.n577 B.n576 585
R135 B.n576 B.n22 585
R136 B.n575 B.n21 585
R137 B.n625 B.n21 585
R138 B.n574 B.n20 585
R139 B.n626 B.n20 585
R140 B.n573 B.n19 585
R141 B.n627 B.n19 585
R142 B.n572 B.n571 585
R143 B.n571 B.n15 585
R144 B.n570 B.n14 585
R145 B.n633 B.n14 585
R146 B.n569 B.n13 585
R147 B.n634 B.n13 585
R148 B.n568 B.n12 585
R149 B.n635 B.n12 585
R150 B.n567 B.n566 585
R151 B.n566 B.n565 585
R152 B.n564 B.n563 585
R153 B.n564 B.n8 585
R154 B.n562 B.n7 585
R155 B.n642 B.n7 585
R156 B.n561 B.n6 585
R157 B.n643 B.n6 585
R158 B.n560 B.n5 585
R159 B.n644 B.n5 585
R160 B.n559 B.n558 585
R161 B.n558 B.n4 585
R162 B.n557 B.n244 585
R163 B.n557 B.n556 585
R164 B.n547 B.n245 585
R165 B.n246 B.n245 585
R166 B.n549 B.n548 585
R167 B.n550 B.n549 585
R168 B.n546 B.n251 585
R169 B.n251 B.n250 585
R170 B.n545 B.n544 585
R171 B.n544 B.n543 585
R172 B.n253 B.n252 585
R173 B.n254 B.n253 585
R174 B.n536 B.n535 585
R175 B.n537 B.n536 585
R176 B.n534 B.n258 585
R177 B.n262 B.n258 585
R178 B.n533 B.n532 585
R179 B.n532 B.n531 585
R180 B.n260 B.n259 585
R181 B.n261 B.n260 585
R182 B.n524 B.n523 585
R183 B.n525 B.n524 585
R184 B.n522 B.n267 585
R185 B.n267 B.n266 585
R186 B.n521 B.n520 585
R187 B.n520 B.n519 585
R188 B.n269 B.n268 585
R189 B.n270 B.n269 585
R190 B.n512 B.n511 585
R191 B.n513 B.n512 585
R192 B.n510 B.n275 585
R193 B.n275 B.n274 585
R194 B.n509 B.n508 585
R195 B.n508 B.n507 585
R196 B.n277 B.n276 585
R197 B.n278 B.n277 585
R198 B.n500 B.n499 585
R199 B.n501 B.n500 585
R200 B.n498 B.n283 585
R201 B.n283 B.n282 585
R202 B.n497 B.n496 585
R203 B.n496 B.n495 585
R204 B.n285 B.n284 585
R205 B.n286 B.n285 585
R206 B.n491 B.n490 585
R207 B.n289 B.n288 585
R208 B.n487 B.n486 585
R209 B.n488 B.n487 585
R210 B.n485 B.n328 585
R211 B.n484 B.n483 585
R212 B.n482 B.n481 585
R213 B.n480 B.n479 585
R214 B.n478 B.n477 585
R215 B.n476 B.n475 585
R216 B.n474 B.n473 585
R217 B.n472 B.n471 585
R218 B.n470 B.n469 585
R219 B.n468 B.n467 585
R220 B.n466 B.n465 585
R221 B.n464 B.n463 585
R222 B.n462 B.n461 585
R223 B.n460 B.n459 585
R224 B.n458 B.n457 585
R225 B.n456 B.n455 585
R226 B.n454 B.n453 585
R227 B.n452 B.n451 585
R228 B.n450 B.n449 585
R229 B.n448 B.n447 585
R230 B.n446 B.n445 585
R231 B.n444 B.n443 585
R232 B.n442 B.n441 585
R233 B.n440 B.n439 585
R234 B.n438 B.n437 585
R235 B.n436 B.n435 585
R236 B.n434 B.n433 585
R237 B.n432 B.n431 585
R238 B.n430 B.n429 585
R239 B.n428 B.n427 585
R240 B.n426 B.n425 585
R241 B.n424 B.n423 585
R242 B.n422 B.n421 585
R243 B.n420 B.n419 585
R244 B.n418 B.n417 585
R245 B.n416 B.n415 585
R246 B.n414 B.n413 585
R247 B.n412 B.n411 585
R248 B.n410 B.n409 585
R249 B.n408 B.n407 585
R250 B.n406 B.n405 585
R251 B.n403 B.n402 585
R252 B.n401 B.n400 585
R253 B.n399 B.n398 585
R254 B.n397 B.n396 585
R255 B.n395 B.n394 585
R256 B.n393 B.n392 585
R257 B.n391 B.n390 585
R258 B.n389 B.n388 585
R259 B.n387 B.n386 585
R260 B.n385 B.n384 585
R261 B.n383 B.n382 585
R262 B.n381 B.n380 585
R263 B.n379 B.n378 585
R264 B.n377 B.n376 585
R265 B.n375 B.n374 585
R266 B.n373 B.n372 585
R267 B.n371 B.n370 585
R268 B.n369 B.n368 585
R269 B.n367 B.n366 585
R270 B.n365 B.n364 585
R271 B.n363 B.n362 585
R272 B.n361 B.n360 585
R273 B.n359 B.n358 585
R274 B.n357 B.n356 585
R275 B.n355 B.n354 585
R276 B.n353 B.n352 585
R277 B.n351 B.n350 585
R278 B.n349 B.n348 585
R279 B.n347 B.n346 585
R280 B.n345 B.n344 585
R281 B.n343 B.n342 585
R282 B.n341 B.n340 585
R283 B.n339 B.n338 585
R284 B.n337 B.n336 585
R285 B.n335 B.n334 585
R286 B.n492 B.n287 585
R287 B.n287 B.n286 585
R288 B.n494 B.n493 585
R289 B.n495 B.n494 585
R290 B.n281 B.n280 585
R291 B.n282 B.n281 585
R292 B.n503 B.n502 585
R293 B.n502 B.n501 585
R294 B.n504 B.n279 585
R295 B.n279 B.n278 585
R296 B.n506 B.n505 585
R297 B.n507 B.n506 585
R298 B.n273 B.n272 585
R299 B.n274 B.n273 585
R300 B.n515 B.n514 585
R301 B.n514 B.n513 585
R302 B.n516 B.n271 585
R303 B.n271 B.n270 585
R304 B.n518 B.n517 585
R305 B.n519 B.n518 585
R306 B.n265 B.n264 585
R307 B.n266 B.n265 585
R308 B.n527 B.n526 585
R309 B.n526 B.n525 585
R310 B.n528 B.n263 585
R311 B.n263 B.n261 585
R312 B.n530 B.n529 585
R313 B.n531 B.n530 585
R314 B.n257 B.n256 585
R315 B.n262 B.n257 585
R316 B.n539 B.n538 585
R317 B.n538 B.n537 585
R318 B.n540 B.n255 585
R319 B.n255 B.n254 585
R320 B.n542 B.n541 585
R321 B.n543 B.n542 585
R322 B.n249 B.n248 585
R323 B.n250 B.n249 585
R324 B.n552 B.n551 585
R325 B.n551 B.n550 585
R326 B.n553 B.n247 585
R327 B.n247 B.n246 585
R328 B.n555 B.n554 585
R329 B.n556 B.n555 585
R330 B.n3 B.n0 585
R331 B.n4 B.n3 585
R332 B.n641 B.n1 585
R333 B.n642 B.n641 585
R334 B.n640 B.n639 585
R335 B.n640 B.n8 585
R336 B.n638 B.n9 585
R337 B.n565 B.n9 585
R338 B.n637 B.n636 585
R339 B.n636 B.n635 585
R340 B.n11 B.n10 585
R341 B.n634 B.n11 585
R342 B.n632 B.n631 585
R343 B.n633 B.n632 585
R344 B.n630 B.n16 585
R345 B.n16 B.n15 585
R346 B.n629 B.n628 585
R347 B.n628 B.n627 585
R348 B.n18 B.n17 585
R349 B.n626 B.n18 585
R350 B.n624 B.n623 585
R351 B.n625 B.n624 585
R352 B.n622 B.n23 585
R353 B.n23 B.n22 585
R354 B.n621 B.n620 585
R355 B.n620 B.n619 585
R356 B.n25 B.n24 585
R357 B.n618 B.n25 585
R358 B.n616 B.n615 585
R359 B.n617 B.n616 585
R360 B.n614 B.n30 585
R361 B.n30 B.n29 585
R362 B.n613 B.n612 585
R363 B.n612 B.n611 585
R364 B.n32 B.n31 585
R365 B.n610 B.n32 585
R366 B.n608 B.n607 585
R367 B.n609 B.n608 585
R368 B.n606 B.n37 585
R369 B.n37 B.n36 585
R370 B.n605 B.n604 585
R371 B.n604 B.n603 585
R372 B.n39 B.n38 585
R373 B.n602 B.n39 585
R374 B.n600 B.n599 585
R375 B.n601 B.n600 585
R376 B.n598 B.n44 585
R377 B.n44 B.n43 585
R378 B.n645 B.n644 585
R379 B.n643 B.n2 585
R380 B.n596 B.n44 454.062
R381 B.n593 B.n86 454.062
R382 B.n334 B.n285 454.062
R383 B.n490 B.n287 454.062
R384 B.n90 B.t15 370.305
R385 B.n87 B.t4 370.305
R386 B.n332 B.t12 370.305
R387 B.n329 B.t8 370.305
R388 B.n594 B.n84 256.663
R389 B.n594 B.n83 256.663
R390 B.n594 B.n82 256.663
R391 B.n594 B.n81 256.663
R392 B.n594 B.n80 256.663
R393 B.n594 B.n79 256.663
R394 B.n594 B.n78 256.663
R395 B.n594 B.n77 256.663
R396 B.n594 B.n76 256.663
R397 B.n594 B.n75 256.663
R398 B.n594 B.n74 256.663
R399 B.n594 B.n73 256.663
R400 B.n594 B.n72 256.663
R401 B.n594 B.n71 256.663
R402 B.n594 B.n70 256.663
R403 B.n594 B.n69 256.663
R404 B.n594 B.n68 256.663
R405 B.n594 B.n67 256.663
R406 B.n594 B.n66 256.663
R407 B.n594 B.n65 256.663
R408 B.n594 B.n64 256.663
R409 B.n594 B.n63 256.663
R410 B.n594 B.n62 256.663
R411 B.n594 B.n61 256.663
R412 B.n594 B.n60 256.663
R413 B.n594 B.n59 256.663
R414 B.n594 B.n58 256.663
R415 B.n594 B.n57 256.663
R416 B.n594 B.n56 256.663
R417 B.n594 B.n55 256.663
R418 B.n594 B.n54 256.663
R419 B.n594 B.n53 256.663
R420 B.n594 B.n52 256.663
R421 B.n594 B.n51 256.663
R422 B.n594 B.n50 256.663
R423 B.n594 B.n49 256.663
R424 B.n594 B.n48 256.663
R425 B.n594 B.n47 256.663
R426 B.n595 B.n594 256.663
R427 B.n489 B.n488 256.663
R428 B.n488 B.n290 256.663
R429 B.n488 B.n291 256.663
R430 B.n488 B.n292 256.663
R431 B.n488 B.n293 256.663
R432 B.n488 B.n294 256.663
R433 B.n488 B.n295 256.663
R434 B.n488 B.n296 256.663
R435 B.n488 B.n297 256.663
R436 B.n488 B.n298 256.663
R437 B.n488 B.n299 256.663
R438 B.n488 B.n300 256.663
R439 B.n488 B.n301 256.663
R440 B.n488 B.n302 256.663
R441 B.n488 B.n303 256.663
R442 B.n488 B.n304 256.663
R443 B.n488 B.n305 256.663
R444 B.n488 B.n306 256.663
R445 B.n488 B.n307 256.663
R446 B.n488 B.n308 256.663
R447 B.n488 B.n309 256.663
R448 B.n488 B.n310 256.663
R449 B.n488 B.n311 256.663
R450 B.n488 B.n312 256.663
R451 B.n488 B.n313 256.663
R452 B.n488 B.n314 256.663
R453 B.n488 B.n315 256.663
R454 B.n488 B.n316 256.663
R455 B.n488 B.n317 256.663
R456 B.n488 B.n318 256.663
R457 B.n488 B.n319 256.663
R458 B.n488 B.n320 256.663
R459 B.n488 B.n321 256.663
R460 B.n488 B.n322 256.663
R461 B.n488 B.n323 256.663
R462 B.n488 B.n324 256.663
R463 B.n488 B.n325 256.663
R464 B.n488 B.n326 256.663
R465 B.n488 B.n327 256.663
R466 B.n647 B.n646 256.663
R467 B.n92 B.n46 163.367
R468 B.n96 B.n95 163.367
R469 B.n100 B.n99 163.367
R470 B.n104 B.n103 163.367
R471 B.n108 B.n107 163.367
R472 B.n112 B.n111 163.367
R473 B.n116 B.n115 163.367
R474 B.n120 B.n119 163.367
R475 B.n124 B.n123 163.367
R476 B.n128 B.n127 163.367
R477 B.n132 B.n131 163.367
R478 B.n136 B.n135 163.367
R479 B.n140 B.n139 163.367
R480 B.n144 B.n143 163.367
R481 B.n148 B.n147 163.367
R482 B.n152 B.n151 163.367
R483 B.n156 B.n155 163.367
R484 B.n161 B.n160 163.367
R485 B.n165 B.n164 163.367
R486 B.n169 B.n168 163.367
R487 B.n173 B.n172 163.367
R488 B.n177 B.n176 163.367
R489 B.n181 B.n180 163.367
R490 B.n185 B.n184 163.367
R491 B.n189 B.n188 163.367
R492 B.n193 B.n192 163.367
R493 B.n197 B.n196 163.367
R494 B.n201 B.n200 163.367
R495 B.n205 B.n204 163.367
R496 B.n209 B.n208 163.367
R497 B.n213 B.n212 163.367
R498 B.n217 B.n216 163.367
R499 B.n221 B.n220 163.367
R500 B.n225 B.n224 163.367
R501 B.n229 B.n228 163.367
R502 B.n233 B.n232 163.367
R503 B.n237 B.n236 163.367
R504 B.n241 B.n240 163.367
R505 B.n593 B.n85 163.367
R506 B.n496 B.n285 163.367
R507 B.n496 B.n283 163.367
R508 B.n500 B.n283 163.367
R509 B.n500 B.n277 163.367
R510 B.n508 B.n277 163.367
R511 B.n508 B.n275 163.367
R512 B.n512 B.n275 163.367
R513 B.n512 B.n269 163.367
R514 B.n520 B.n269 163.367
R515 B.n520 B.n267 163.367
R516 B.n524 B.n267 163.367
R517 B.n524 B.n260 163.367
R518 B.n532 B.n260 163.367
R519 B.n532 B.n258 163.367
R520 B.n536 B.n258 163.367
R521 B.n536 B.n253 163.367
R522 B.n544 B.n253 163.367
R523 B.n544 B.n251 163.367
R524 B.n549 B.n251 163.367
R525 B.n549 B.n245 163.367
R526 B.n557 B.n245 163.367
R527 B.n558 B.n557 163.367
R528 B.n558 B.n5 163.367
R529 B.n6 B.n5 163.367
R530 B.n7 B.n6 163.367
R531 B.n564 B.n7 163.367
R532 B.n566 B.n564 163.367
R533 B.n566 B.n12 163.367
R534 B.n13 B.n12 163.367
R535 B.n14 B.n13 163.367
R536 B.n571 B.n14 163.367
R537 B.n571 B.n19 163.367
R538 B.n20 B.n19 163.367
R539 B.n21 B.n20 163.367
R540 B.n576 B.n21 163.367
R541 B.n576 B.n26 163.367
R542 B.n27 B.n26 163.367
R543 B.n28 B.n27 163.367
R544 B.n581 B.n28 163.367
R545 B.n581 B.n33 163.367
R546 B.n34 B.n33 163.367
R547 B.n35 B.n34 163.367
R548 B.n586 B.n35 163.367
R549 B.n586 B.n40 163.367
R550 B.n41 B.n40 163.367
R551 B.n42 B.n41 163.367
R552 B.n86 B.n42 163.367
R553 B.n487 B.n289 163.367
R554 B.n487 B.n328 163.367
R555 B.n483 B.n482 163.367
R556 B.n479 B.n478 163.367
R557 B.n475 B.n474 163.367
R558 B.n471 B.n470 163.367
R559 B.n467 B.n466 163.367
R560 B.n463 B.n462 163.367
R561 B.n459 B.n458 163.367
R562 B.n455 B.n454 163.367
R563 B.n451 B.n450 163.367
R564 B.n447 B.n446 163.367
R565 B.n443 B.n442 163.367
R566 B.n439 B.n438 163.367
R567 B.n435 B.n434 163.367
R568 B.n431 B.n430 163.367
R569 B.n427 B.n426 163.367
R570 B.n423 B.n422 163.367
R571 B.n419 B.n418 163.367
R572 B.n415 B.n414 163.367
R573 B.n411 B.n410 163.367
R574 B.n407 B.n406 163.367
R575 B.n402 B.n401 163.367
R576 B.n398 B.n397 163.367
R577 B.n394 B.n393 163.367
R578 B.n390 B.n389 163.367
R579 B.n386 B.n385 163.367
R580 B.n382 B.n381 163.367
R581 B.n378 B.n377 163.367
R582 B.n374 B.n373 163.367
R583 B.n370 B.n369 163.367
R584 B.n366 B.n365 163.367
R585 B.n362 B.n361 163.367
R586 B.n358 B.n357 163.367
R587 B.n354 B.n353 163.367
R588 B.n350 B.n349 163.367
R589 B.n346 B.n345 163.367
R590 B.n342 B.n341 163.367
R591 B.n338 B.n337 163.367
R592 B.n494 B.n287 163.367
R593 B.n494 B.n281 163.367
R594 B.n502 B.n281 163.367
R595 B.n502 B.n279 163.367
R596 B.n506 B.n279 163.367
R597 B.n506 B.n273 163.367
R598 B.n514 B.n273 163.367
R599 B.n514 B.n271 163.367
R600 B.n518 B.n271 163.367
R601 B.n518 B.n265 163.367
R602 B.n526 B.n265 163.367
R603 B.n526 B.n263 163.367
R604 B.n530 B.n263 163.367
R605 B.n530 B.n257 163.367
R606 B.n538 B.n257 163.367
R607 B.n538 B.n255 163.367
R608 B.n542 B.n255 163.367
R609 B.n542 B.n249 163.367
R610 B.n551 B.n249 163.367
R611 B.n551 B.n247 163.367
R612 B.n555 B.n247 163.367
R613 B.n555 B.n3 163.367
R614 B.n645 B.n3 163.367
R615 B.n641 B.n2 163.367
R616 B.n641 B.n640 163.367
R617 B.n640 B.n9 163.367
R618 B.n636 B.n9 163.367
R619 B.n636 B.n11 163.367
R620 B.n632 B.n11 163.367
R621 B.n632 B.n16 163.367
R622 B.n628 B.n16 163.367
R623 B.n628 B.n18 163.367
R624 B.n624 B.n18 163.367
R625 B.n624 B.n23 163.367
R626 B.n620 B.n23 163.367
R627 B.n620 B.n25 163.367
R628 B.n616 B.n25 163.367
R629 B.n616 B.n30 163.367
R630 B.n612 B.n30 163.367
R631 B.n612 B.n32 163.367
R632 B.n608 B.n32 163.367
R633 B.n608 B.n37 163.367
R634 B.n604 B.n37 163.367
R635 B.n604 B.n39 163.367
R636 B.n600 B.n39 163.367
R637 B.n600 B.n44 163.367
R638 B.n87 B.t6 103.302
R639 B.n332 B.t14 103.302
R640 B.n90 B.t16 103.29
R641 B.n329 B.t11 103.29
R642 B.n488 B.n286 85.0425
R643 B.n594 B.n43 85.0425
R644 B.n596 B.n595 71.676
R645 B.n92 B.n47 71.676
R646 B.n96 B.n48 71.676
R647 B.n100 B.n49 71.676
R648 B.n104 B.n50 71.676
R649 B.n108 B.n51 71.676
R650 B.n112 B.n52 71.676
R651 B.n116 B.n53 71.676
R652 B.n120 B.n54 71.676
R653 B.n124 B.n55 71.676
R654 B.n128 B.n56 71.676
R655 B.n132 B.n57 71.676
R656 B.n136 B.n58 71.676
R657 B.n140 B.n59 71.676
R658 B.n144 B.n60 71.676
R659 B.n148 B.n61 71.676
R660 B.n152 B.n62 71.676
R661 B.n156 B.n63 71.676
R662 B.n161 B.n64 71.676
R663 B.n165 B.n65 71.676
R664 B.n169 B.n66 71.676
R665 B.n173 B.n67 71.676
R666 B.n177 B.n68 71.676
R667 B.n181 B.n69 71.676
R668 B.n185 B.n70 71.676
R669 B.n189 B.n71 71.676
R670 B.n193 B.n72 71.676
R671 B.n197 B.n73 71.676
R672 B.n201 B.n74 71.676
R673 B.n205 B.n75 71.676
R674 B.n209 B.n76 71.676
R675 B.n213 B.n77 71.676
R676 B.n217 B.n78 71.676
R677 B.n221 B.n79 71.676
R678 B.n225 B.n80 71.676
R679 B.n229 B.n81 71.676
R680 B.n233 B.n82 71.676
R681 B.n237 B.n83 71.676
R682 B.n241 B.n84 71.676
R683 B.n85 B.n84 71.676
R684 B.n240 B.n83 71.676
R685 B.n236 B.n82 71.676
R686 B.n232 B.n81 71.676
R687 B.n228 B.n80 71.676
R688 B.n224 B.n79 71.676
R689 B.n220 B.n78 71.676
R690 B.n216 B.n77 71.676
R691 B.n212 B.n76 71.676
R692 B.n208 B.n75 71.676
R693 B.n204 B.n74 71.676
R694 B.n200 B.n73 71.676
R695 B.n196 B.n72 71.676
R696 B.n192 B.n71 71.676
R697 B.n188 B.n70 71.676
R698 B.n184 B.n69 71.676
R699 B.n180 B.n68 71.676
R700 B.n176 B.n67 71.676
R701 B.n172 B.n66 71.676
R702 B.n168 B.n65 71.676
R703 B.n164 B.n64 71.676
R704 B.n160 B.n63 71.676
R705 B.n155 B.n62 71.676
R706 B.n151 B.n61 71.676
R707 B.n147 B.n60 71.676
R708 B.n143 B.n59 71.676
R709 B.n139 B.n58 71.676
R710 B.n135 B.n57 71.676
R711 B.n131 B.n56 71.676
R712 B.n127 B.n55 71.676
R713 B.n123 B.n54 71.676
R714 B.n119 B.n53 71.676
R715 B.n115 B.n52 71.676
R716 B.n111 B.n51 71.676
R717 B.n107 B.n50 71.676
R718 B.n103 B.n49 71.676
R719 B.n99 B.n48 71.676
R720 B.n95 B.n47 71.676
R721 B.n595 B.n46 71.676
R722 B.n490 B.n489 71.676
R723 B.n328 B.n290 71.676
R724 B.n482 B.n291 71.676
R725 B.n478 B.n292 71.676
R726 B.n474 B.n293 71.676
R727 B.n470 B.n294 71.676
R728 B.n466 B.n295 71.676
R729 B.n462 B.n296 71.676
R730 B.n458 B.n297 71.676
R731 B.n454 B.n298 71.676
R732 B.n450 B.n299 71.676
R733 B.n446 B.n300 71.676
R734 B.n442 B.n301 71.676
R735 B.n438 B.n302 71.676
R736 B.n434 B.n303 71.676
R737 B.n430 B.n304 71.676
R738 B.n426 B.n305 71.676
R739 B.n422 B.n306 71.676
R740 B.n418 B.n307 71.676
R741 B.n414 B.n308 71.676
R742 B.n410 B.n309 71.676
R743 B.n406 B.n310 71.676
R744 B.n401 B.n311 71.676
R745 B.n397 B.n312 71.676
R746 B.n393 B.n313 71.676
R747 B.n389 B.n314 71.676
R748 B.n385 B.n315 71.676
R749 B.n381 B.n316 71.676
R750 B.n377 B.n317 71.676
R751 B.n373 B.n318 71.676
R752 B.n369 B.n319 71.676
R753 B.n365 B.n320 71.676
R754 B.n361 B.n321 71.676
R755 B.n357 B.n322 71.676
R756 B.n353 B.n323 71.676
R757 B.n349 B.n324 71.676
R758 B.n345 B.n325 71.676
R759 B.n341 B.n326 71.676
R760 B.n337 B.n327 71.676
R761 B.n489 B.n289 71.676
R762 B.n483 B.n290 71.676
R763 B.n479 B.n291 71.676
R764 B.n475 B.n292 71.676
R765 B.n471 B.n293 71.676
R766 B.n467 B.n294 71.676
R767 B.n463 B.n295 71.676
R768 B.n459 B.n296 71.676
R769 B.n455 B.n297 71.676
R770 B.n451 B.n298 71.676
R771 B.n447 B.n299 71.676
R772 B.n443 B.n300 71.676
R773 B.n439 B.n301 71.676
R774 B.n435 B.n302 71.676
R775 B.n431 B.n303 71.676
R776 B.n427 B.n304 71.676
R777 B.n423 B.n305 71.676
R778 B.n419 B.n306 71.676
R779 B.n415 B.n307 71.676
R780 B.n411 B.n308 71.676
R781 B.n407 B.n309 71.676
R782 B.n402 B.n310 71.676
R783 B.n398 B.n311 71.676
R784 B.n394 B.n312 71.676
R785 B.n390 B.n313 71.676
R786 B.n386 B.n314 71.676
R787 B.n382 B.n315 71.676
R788 B.n378 B.n316 71.676
R789 B.n374 B.n317 71.676
R790 B.n370 B.n318 71.676
R791 B.n366 B.n319 71.676
R792 B.n362 B.n320 71.676
R793 B.n358 B.n321 71.676
R794 B.n354 B.n322 71.676
R795 B.n350 B.n323 71.676
R796 B.n346 B.n324 71.676
R797 B.n342 B.n325 71.676
R798 B.n338 B.n326 71.676
R799 B.n334 B.n327 71.676
R800 B.n646 B.n645 71.676
R801 B.n646 B.n2 71.676
R802 B.n88 B.t7 69.7505
R803 B.n333 B.t13 69.7505
R804 B.n91 B.t17 69.7387
R805 B.n330 B.t10 69.7387
R806 B.n158 B.n91 59.5399
R807 B.n89 B.n88 59.5399
R808 B.n404 B.n333 59.5399
R809 B.n331 B.n330 59.5399
R810 B.n495 B.n286 50.2862
R811 B.n495 B.n282 50.2862
R812 B.n501 B.n282 50.2862
R813 B.n501 B.n278 50.2862
R814 B.n507 B.n278 50.2862
R815 B.n513 B.n274 50.2862
R816 B.n513 B.n270 50.2862
R817 B.n519 B.n270 50.2862
R818 B.n519 B.n266 50.2862
R819 B.n525 B.n266 50.2862
R820 B.n525 B.n261 50.2862
R821 B.n531 B.n261 50.2862
R822 B.n531 B.n262 50.2862
R823 B.n537 B.n254 50.2862
R824 B.n543 B.n254 50.2862
R825 B.n543 B.n250 50.2862
R826 B.n550 B.n250 50.2862
R827 B.n556 B.n246 50.2862
R828 B.n556 B.n4 50.2862
R829 B.n644 B.n4 50.2862
R830 B.n644 B.n643 50.2862
R831 B.n643 B.n642 50.2862
R832 B.n642 B.n8 50.2862
R833 B.n565 B.n8 50.2862
R834 B.n635 B.n634 50.2862
R835 B.n634 B.n633 50.2862
R836 B.n633 B.n15 50.2862
R837 B.n627 B.n15 50.2862
R838 B.n626 B.n625 50.2862
R839 B.n625 B.n22 50.2862
R840 B.n619 B.n22 50.2862
R841 B.n619 B.n618 50.2862
R842 B.n618 B.n617 50.2862
R843 B.n617 B.n29 50.2862
R844 B.n611 B.n29 50.2862
R845 B.n611 B.n610 50.2862
R846 B.n609 B.n36 50.2862
R847 B.n603 B.n36 50.2862
R848 B.n603 B.n602 50.2862
R849 B.n602 B.n601 50.2862
R850 B.n601 B.n43 50.2862
R851 B.n507 B.t9 48.8072
R852 B.t5 B.n609 48.8072
R853 B.n537 B.t2 36.9753
R854 B.n627 B.t1 36.9753
R855 B.n91 B.n90 33.552
R856 B.n88 B.n87 33.552
R857 B.n333 B.n332 33.552
R858 B.n330 B.n329 33.552
R859 B.t3 B.n246 32.5383
R860 B.n565 B.t0 32.5383
R861 B.n492 B.n491 29.5029
R862 B.n335 B.n284 29.5029
R863 B.n592 B.n591 29.5029
R864 B.n598 B.n597 29.5029
R865 B B.n647 18.0485
R866 B.n550 B.t3 17.7484
R867 B.n635 B.t0 17.7484
R868 B.n262 B.t2 13.3114
R869 B.t1 B.n626 13.3114
R870 B.n493 B.n492 10.6151
R871 B.n493 B.n280 10.6151
R872 B.n503 B.n280 10.6151
R873 B.n504 B.n503 10.6151
R874 B.n505 B.n504 10.6151
R875 B.n505 B.n272 10.6151
R876 B.n515 B.n272 10.6151
R877 B.n516 B.n515 10.6151
R878 B.n517 B.n516 10.6151
R879 B.n517 B.n264 10.6151
R880 B.n527 B.n264 10.6151
R881 B.n528 B.n527 10.6151
R882 B.n529 B.n528 10.6151
R883 B.n529 B.n256 10.6151
R884 B.n539 B.n256 10.6151
R885 B.n540 B.n539 10.6151
R886 B.n541 B.n540 10.6151
R887 B.n541 B.n248 10.6151
R888 B.n552 B.n248 10.6151
R889 B.n553 B.n552 10.6151
R890 B.n554 B.n553 10.6151
R891 B.n554 B.n0 10.6151
R892 B.n491 B.n288 10.6151
R893 B.n486 B.n288 10.6151
R894 B.n486 B.n485 10.6151
R895 B.n485 B.n484 10.6151
R896 B.n484 B.n481 10.6151
R897 B.n481 B.n480 10.6151
R898 B.n480 B.n477 10.6151
R899 B.n477 B.n476 10.6151
R900 B.n476 B.n473 10.6151
R901 B.n473 B.n472 10.6151
R902 B.n472 B.n469 10.6151
R903 B.n469 B.n468 10.6151
R904 B.n468 B.n465 10.6151
R905 B.n465 B.n464 10.6151
R906 B.n464 B.n461 10.6151
R907 B.n461 B.n460 10.6151
R908 B.n460 B.n457 10.6151
R909 B.n457 B.n456 10.6151
R910 B.n456 B.n453 10.6151
R911 B.n453 B.n452 10.6151
R912 B.n452 B.n449 10.6151
R913 B.n449 B.n448 10.6151
R914 B.n448 B.n445 10.6151
R915 B.n445 B.n444 10.6151
R916 B.n444 B.n441 10.6151
R917 B.n441 B.n440 10.6151
R918 B.n440 B.n437 10.6151
R919 B.n437 B.n436 10.6151
R920 B.n436 B.n433 10.6151
R921 B.n433 B.n432 10.6151
R922 B.n432 B.n429 10.6151
R923 B.n429 B.n428 10.6151
R924 B.n428 B.n425 10.6151
R925 B.n425 B.n424 10.6151
R926 B.n421 B.n420 10.6151
R927 B.n420 B.n417 10.6151
R928 B.n417 B.n416 10.6151
R929 B.n416 B.n413 10.6151
R930 B.n413 B.n412 10.6151
R931 B.n412 B.n409 10.6151
R932 B.n409 B.n408 10.6151
R933 B.n408 B.n405 10.6151
R934 B.n403 B.n400 10.6151
R935 B.n400 B.n399 10.6151
R936 B.n399 B.n396 10.6151
R937 B.n396 B.n395 10.6151
R938 B.n395 B.n392 10.6151
R939 B.n392 B.n391 10.6151
R940 B.n391 B.n388 10.6151
R941 B.n388 B.n387 10.6151
R942 B.n387 B.n384 10.6151
R943 B.n384 B.n383 10.6151
R944 B.n383 B.n380 10.6151
R945 B.n380 B.n379 10.6151
R946 B.n379 B.n376 10.6151
R947 B.n376 B.n375 10.6151
R948 B.n375 B.n372 10.6151
R949 B.n372 B.n371 10.6151
R950 B.n371 B.n368 10.6151
R951 B.n368 B.n367 10.6151
R952 B.n367 B.n364 10.6151
R953 B.n364 B.n363 10.6151
R954 B.n363 B.n360 10.6151
R955 B.n360 B.n359 10.6151
R956 B.n359 B.n356 10.6151
R957 B.n356 B.n355 10.6151
R958 B.n355 B.n352 10.6151
R959 B.n352 B.n351 10.6151
R960 B.n351 B.n348 10.6151
R961 B.n348 B.n347 10.6151
R962 B.n347 B.n344 10.6151
R963 B.n344 B.n343 10.6151
R964 B.n343 B.n340 10.6151
R965 B.n340 B.n339 10.6151
R966 B.n339 B.n336 10.6151
R967 B.n336 B.n335 10.6151
R968 B.n497 B.n284 10.6151
R969 B.n498 B.n497 10.6151
R970 B.n499 B.n498 10.6151
R971 B.n499 B.n276 10.6151
R972 B.n509 B.n276 10.6151
R973 B.n510 B.n509 10.6151
R974 B.n511 B.n510 10.6151
R975 B.n511 B.n268 10.6151
R976 B.n521 B.n268 10.6151
R977 B.n522 B.n521 10.6151
R978 B.n523 B.n522 10.6151
R979 B.n523 B.n259 10.6151
R980 B.n533 B.n259 10.6151
R981 B.n534 B.n533 10.6151
R982 B.n535 B.n534 10.6151
R983 B.n535 B.n252 10.6151
R984 B.n545 B.n252 10.6151
R985 B.n546 B.n545 10.6151
R986 B.n548 B.n546 10.6151
R987 B.n548 B.n547 10.6151
R988 B.n547 B.n244 10.6151
R989 B.n559 B.n244 10.6151
R990 B.n560 B.n559 10.6151
R991 B.n561 B.n560 10.6151
R992 B.n562 B.n561 10.6151
R993 B.n563 B.n562 10.6151
R994 B.n567 B.n563 10.6151
R995 B.n568 B.n567 10.6151
R996 B.n569 B.n568 10.6151
R997 B.n570 B.n569 10.6151
R998 B.n572 B.n570 10.6151
R999 B.n573 B.n572 10.6151
R1000 B.n574 B.n573 10.6151
R1001 B.n575 B.n574 10.6151
R1002 B.n577 B.n575 10.6151
R1003 B.n578 B.n577 10.6151
R1004 B.n579 B.n578 10.6151
R1005 B.n580 B.n579 10.6151
R1006 B.n582 B.n580 10.6151
R1007 B.n583 B.n582 10.6151
R1008 B.n584 B.n583 10.6151
R1009 B.n585 B.n584 10.6151
R1010 B.n587 B.n585 10.6151
R1011 B.n588 B.n587 10.6151
R1012 B.n589 B.n588 10.6151
R1013 B.n590 B.n589 10.6151
R1014 B.n591 B.n590 10.6151
R1015 B.n639 B.n1 10.6151
R1016 B.n639 B.n638 10.6151
R1017 B.n638 B.n637 10.6151
R1018 B.n637 B.n10 10.6151
R1019 B.n631 B.n10 10.6151
R1020 B.n631 B.n630 10.6151
R1021 B.n630 B.n629 10.6151
R1022 B.n629 B.n17 10.6151
R1023 B.n623 B.n17 10.6151
R1024 B.n623 B.n622 10.6151
R1025 B.n622 B.n621 10.6151
R1026 B.n621 B.n24 10.6151
R1027 B.n615 B.n24 10.6151
R1028 B.n615 B.n614 10.6151
R1029 B.n614 B.n613 10.6151
R1030 B.n613 B.n31 10.6151
R1031 B.n607 B.n31 10.6151
R1032 B.n607 B.n606 10.6151
R1033 B.n606 B.n605 10.6151
R1034 B.n605 B.n38 10.6151
R1035 B.n599 B.n38 10.6151
R1036 B.n599 B.n598 10.6151
R1037 B.n597 B.n45 10.6151
R1038 B.n93 B.n45 10.6151
R1039 B.n94 B.n93 10.6151
R1040 B.n97 B.n94 10.6151
R1041 B.n98 B.n97 10.6151
R1042 B.n101 B.n98 10.6151
R1043 B.n102 B.n101 10.6151
R1044 B.n105 B.n102 10.6151
R1045 B.n106 B.n105 10.6151
R1046 B.n109 B.n106 10.6151
R1047 B.n110 B.n109 10.6151
R1048 B.n113 B.n110 10.6151
R1049 B.n114 B.n113 10.6151
R1050 B.n117 B.n114 10.6151
R1051 B.n118 B.n117 10.6151
R1052 B.n121 B.n118 10.6151
R1053 B.n122 B.n121 10.6151
R1054 B.n125 B.n122 10.6151
R1055 B.n126 B.n125 10.6151
R1056 B.n129 B.n126 10.6151
R1057 B.n130 B.n129 10.6151
R1058 B.n133 B.n130 10.6151
R1059 B.n134 B.n133 10.6151
R1060 B.n137 B.n134 10.6151
R1061 B.n138 B.n137 10.6151
R1062 B.n141 B.n138 10.6151
R1063 B.n142 B.n141 10.6151
R1064 B.n145 B.n142 10.6151
R1065 B.n146 B.n145 10.6151
R1066 B.n149 B.n146 10.6151
R1067 B.n150 B.n149 10.6151
R1068 B.n153 B.n150 10.6151
R1069 B.n154 B.n153 10.6151
R1070 B.n157 B.n154 10.6151
R1071 B.n162 B.n159 10.6151
R1072 B.n163 B.n162 10.6151
R1073 B.n166 B.n163 10.6151
R1074 B.n167 B.n166 10.6151
R1075 B.n170 B.n167 10.6151
R1076 B.n171 B.n170 10.6151
R1077 B.n174 B.n171 10.6151
R1078 B.n175 B.n174 10.6151
R1079 B.n179 B.n178 10.6151
R1080 B.n182 B.n179 10.6151
R1081 B.n183 B.n182 10.6151
R1082 B.n186 B.n183 10.6151
R1083 B.n187 B.n186 10.6151
R1084 B.n190 B.n187 10.6151
R1085 B.n191 B.n190 10.6151
R1086 B.n194 B.n191 10.6151
R1087 B.n195 B.n194 10.6151
R1088 B.n198 B.n195 10.6151
R1089 B.n199 B.n198 10.6151
R1090 B.n202 B.n199 10.6151
R1091 B.n203 B.n202 10.6151
R1092 B.n206 B.n203 10.6151
R1093 B.n207 B.n206 10.6151
R1094 B.n210 B.n207 10.6151
R1095 B.n211 B.n210 10.6151
R1096 B.n214 B.n211 10.6151
R1097 B.n215 B.n214 10.6151
R1098 B.n218 B.n215 10.6151
R1099 B.n219 B.n218 10.6151
R1100 B.n222 B.n219 10.6151
R1101 B.n223 B.n222 10.6151
R1102 B.n226 B.n223 10.6151
R1103 B.n227 B.n226 10.6151
R1104 B.n230 B.n227 10.6151
R1105 B.n231 B.n230 10.6151
R1106 B.n234 B.n231 10.6151
R1107 B.n235 B.n234 10.6151
R1108 B.n238 B.n235 10.6151
R1109 B.n239 B.n238 10.6151
R1110 B.n242 B.n239 10.6151
R1111 B.n243 B.n242 10.6151
R1112 B.n592 B.n243 10.6151
R1113 B.n647 B.n0 8.11757
R1114 B.n647 B.n1 8.11757
R1115 B.n421 B.n331 6.5566
R1116 B.n405 B.n404 6.5566
R1117 B.n159 B.n158 6.5566
R1118 B.n175 B.n89 6.5566
R1119 B.n424 B.n331 4.05904
R1120 B.n404 B.n403 4.05904
R1121 B.n158 B.n157 4.05904
R1122 B.n178 B.n89 4.05904
R1123 B.t9 B.n274 1.47949
R1124 B.n610 B.t5 1.47949
R1125 VP.n2 VP.t0 200.209
R1126 VP.n2 VP.t1 199.901
R1127 VP.n4 VP.n3 180.237
R1128 VP.n12 VP.n11 180.237
R1129 VP.n4 VP.t2 165.257
R1130 VP.n11 VP.t3 165.257
R1131 VP.n10 VP.n0 161.3
R1132 VP.n9 VP.n8 161.3
R1133 VP.n7 VP.n1 161.3
R1134 VP.n6 VP.n5 161.3
R1135 VP.n9 VP.n1 56.5617
R1136 VP.n3 VP.n2 54.0234
R1137 VP.n5 VP.n1 24.5923
R1138 VP.n10 VP.n9 24.5923
R1139 VP.n5 VP.n4 5.65662
R1140 VP.n11 VP.n10 5.65662
R1141 VP.n6 VP.n3 0.189894
R1142 VP.n7 VP.n6 0.189894
R1143 VP.n8 VP.n7 0.189894
R1144 VP.n8 VP.n0 0.189894
R1145 VP.n12 VP.n0 0.189894
R1146 VP VP.n12 0.0516364
R1147 VDD1 VDD1.n1 99.8015
R1148 VDD1 VDD1.n0 62.8701
R1149 VDD1.n0 VDD1.t3 2.063
R1150 VDD1.n0 VDD1.t2 2.063
R1151 VDD1.n1 VDD1.t1 2.063
R1152 VDD1.n1 VDD1.t0 2.063
C0 VDD2 VTAIL 4.89551f
C1 VDD2 VDD1 0.735181f
C2 VN VP 4.88294f
C3 VTAIL VP 3.17957f
C4 VDD1 VP 3.50703f
C5 VTAIL VN 3.16546f
C6 VN VDD1 0.148365f
C7 VTAIL VDD1 4.84934f
C8 VDD2 VP 0.318397f
C9 VDD2 VN 3.33743f
C10 VDD2 B 2.907846f
C11 VDD1 B 6.36342f
C12 VTAIL B 7.925405f
C13 VN B 8.43953f
C14 VP B 6.21795f
C15 VDD1.t3 B 0.202779f
C16 VDD1.t2 B 0.202779f
C17 VDD1.n0 B 1.78059f
C18 VDD1.t1 B 0.202779f
C19 VDD1.t0 B 0.202779f
C20 VDD1.n1 B 2.32946f
C21 VP.n0 B 0.037846f
C22 VP.t3 B 1.37597f
C23 VP.n1 B 0.055015f
C24 VP.t0 B 1.48957f
C25 VP.t1 B 1.48852f
C26 VP.n2 B 2.38921f
C27 VP.n3 B 1.9369f
C28 VP.t2 B 1.37597f
C29 VP.n4 B 0.57354f
C30 VP.n5 B 0.043503f
C31 VP.n6 B 0.037846f
C32 VP.n7 B 0.037846f
C33 VP.n8 B 0.037846f
C34 VP.n9 B 0.055015f
C35 VP.n10 B 0.043503f
C36 VP.n11 B 0.57354f
C37 VP.n12 B 0.036812f
C38 VDD2.t2 B 0.202747f
C39 VDD2.t3 B 0.202747f
C40 VDD2.n0 B 2.3043f
C41 VDD2.t0 B 0.202747f
C42 VDD2.t1 B 0.202747f
C43 VDD2.n1 B 1.77998f
C44 VDD2.n2 B 3.17054f
C45 VTAIL.t5 B 1.33674f
C46 VTAIL.n0 B 0.280571f
C47 VTAIL.t3 B 1.33674f
C48 VTAIL.n1 B 0.317069f
C49 VTAIL.t2 B 1.33674f
C50 VTAIL.n2 B 1.03446f
C51 VTAIL.t6 B 1.33675f
C52 VTAIL.n3 B 1.03445f
C53 VTAIL.t7 B 1.33675f
C54 VTAIL.n4 B 0.31706f
C55 VTAIL.t0 B 1.33675f
C56 VTAIL.n5 B 0.31706f
C57 VTAIL.t1 B 1.33674f
C58 VTAIL.n6 B 1.03446f
C59 VTAIL.t4 B 1.33674f
C60 VTAIL.n7 B 0.991781f
C61 VN.t1 B 1.4572f
C62 VN.t0 B 1.45618f
C63 VN.n0 B 1.09831f
C64 VN.t2 B 1.4572f
C65 VN.t3 B 1.45618f
C66 VN.n1 B 2.35852f
.ends

