* NGSPICE file created from diff_pair_sample_1312.ext - technology: sky130A

.subckt diff_pair_sample_1312 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t5 VN.t0 VTAIL.t9 B.t1 sky130_fd_pr__nfet_01v8 ad=5.0856 pd=26.86 as=2.1516 ps=13.37 w=13.04 l=0.32
X1 VDD1.t5 VP.t0 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=2.1516 pd=13.37 as=5.0856 ps=26.86 w=13.04 l=0.32
X2 B.t19 B.t17 B.t18 B.t7 sky130_fd_pr__nfet_01v8 ad=5.0856 pd=26.86 as=0 ps=0 w=13.04 l=0.32
X3 VTAIL.t7 VN.t1 VDD2.t4 B.t0 sky130_fd_pr__nfet_01v8 ad=2.1516 pd=13.37 as=2.1516 ps=13.37 w=13.04 l=0.32
X4 VTAIL.t11 VP.t1 VDD1.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=2.1516 pd=13.37 as=2.1516 ps=13.37 w=13.04 l=0.32
X5 VDD2.t3 VN.t2 VTAIL.t4 B.t5 sky130_fd_pr__nfet_01v8 ad=2.1516 pd=13.37 as=5.0856 ps=26.86 w=13.04 l=0.32
X6 B.t16 B.t14 B.t15 B.t11 sky130_fd_pr__nfet_01v8 ad=5.0856 pd=26.86 as=0 ps=0 w=13.04 l=0.32
X7 VTAIL.t8 VN.t3 VDD2.t2 B.t4 sky130_fd_pr__nfet_01v8 ad=2.1516 pd=13.37 as=2.1516 ps=13.37 w=13.04 l=0.32
X8 VDD2.t1 VN.t4 VTAIL.t5 B.t2 sky130_fd_pr__nfet_01v8 ad=2.1516 pd=13.37 as=5.0856 ps=26.86 w=13.04 l=0.32
X9 VDD2.t0 VN.t5 VTAIL.t6 B.t3 sky130_fd_pr__nfet_01v8 ad=5.0856 pd=26.86 as=2.1516 ps=13.37 w=13.04 l=0.32
X10 VDD1.t3 VP.t2 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=5.0856 pd=26.86 as=2.1516 ps=13.37 w=13.04 l=0.32
X11 VDD1.t2 VP.t3 VTAIL.t10 B.t5 sky130_fd_pr__nfet_01v8 ad=2.1516 pd=13.37 as=5.0856 ps=26.86 w=13.04 l=0.32
X12 B.t13 B.t10 B.t12 B.t11 sky130_fd_pr__nfet_01v8 ad=5.0856 pd=26.86 as=0 ps=0 w=13.04 l=0.32
X13 VTAIL.t0 VP.t4 VDD1.t1 B.t0 sky130_fd_pr__nfet_01v8 ad=2.1516 pd=13.37 as=2.1516 ps=13.37 w=13.04 l=0.32
X14 B.t9 B.t6 B.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=5.0856 pd=26.86 as=0 ps=0 w=13.04 l=0.32
X15 VDD1.t0 VP.t5 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=5.0856 pd=26.86 as=2.1516 ps=13.37 w=13.04 l=0.32
R0 VN.n0 VN.t0 1131.69
R1 VN.n4 VN.t4 1131.69
R2 VN.n2 VN.t2 1101.89
R3 VN.n6 VN.t5 1101.89
R4 VN.n1 VN.t1 1079.98
R5 VN.n5 VN.t3 1079.98
R6 VN.n3 VN.n2 161.3
R7 VN.n7 VN.n6 161.3
R8 VN.n2 VN.n1 73.0308
R9 VN.n6 VN.n5 73.0308
R10 VN.n7 VN.n4 65.9987
R11 VN.n3 VN.n0 65.9987
R12 VN VN.n7 40.8774
R13 VN.n5 VN.n4 29.7615
R14 VN.n1 VN.n0 29.7615
R15 VN VN.n3 0.0516364
R16 VTAIL.n7 VTAIL.t5 49.8953
R17 VTAIL.n11 VTAIL.t4 49.8942
R18 VTAIL.n2 VTAIL.t2 49.8942
R19 VTAIL.n10 VTAIL.t10 49.8942
R20 VTAIL.n9 VTAIL.n8 48.3769
R21 VTAIL.n6 VTAIL.n5 48.3769
R22 VTAIL.n1 VTAIL.n0 48.3758
R23 VTAIL.n4 VTAIL.n3 48.3758
R24 VTAIL.n6 VTAIL.n4 24.7289
R25 VTAIL.n11 VTAIL.n10 24.1686
R26 VTAIL.n0 VTAIL.t9 1.5189
R27 VTAIL.n0 VTAIL.t7 1.5189
R28 VTAIL.n3 VTAIL.t3 1.5189
R29 VTAIL.n3 VTAIL.t11 1.5189
R30 VTAIL.n8 VTAIL.t1 1.5189
R31 VTAIL.n8 VTAIL.t0 1.5189
R32 VTAIL.n5 VTAIL.t6 1.5189
R33 VTAIL.n5 VTAIL.t8 1.5189
R34 VTAIL.n9 VTAIL.n7 0.7505
R35 VTAIL.n2 VTAIL.n1 0.7505
R36 VTAIL.n7 VTAIL.n6 0.560845
R37 VTAIL.n10 VTAIL.n9 0.560845
R38 VTAIL.n4 VTAIL.n2 0.560845
R39 VTAIL VTAIL.n11 0.362569
R40 VTAIL VTAIL.n1 0.198776
R41 VDD2.n1 VDD2.t5 66.9379
R42 VDD2.n2 VDD2.t0 66.5741
R43 VDD2.n1 VDD2.n0 65.1393
R44 VDD2 VDD2.n3 65.1365
R45 VDD2.n2 VDD2.n1 36.7778
R46 VDD2.n3 VDD2.t2 1.5189
R47 VDD2.n3 VDD2.t1 1.5189
R48 VDD2.n0 VDD2.t4 1.5189
R49 VDD2.n0 VDD2.t3 1.5189
R50 VDD2 VDD2.n2 0.478948
R51 B.n85 B.t14 1195.83
R52 B.n82 B.t10 1195.83
R53 B.n359 B.t6 1195.83
R54 B.n356 B.t17 1195.83
R55 B.n627 B.n626 585
R56 B.n628 B.n627 585
R57 B.n278 B.n80 585
R58 B.n277 B.n276 585
R59 B.n275 B.n274 585
R60 B.n273 B.n272 585
R61 B.n271 B.n270 585
R62 B.n269 B.n268 585
R63 B.n267 B.n266 585
R64 B.n265 B.n264 585
R65 B.n263 B.n262 585
R66 B.n261 B.n260 585
R67 B.n259 B.n258 585
R68 B.n257 B.n256 585
R69 B.n255 B.n254 585
R70 B.n253 B.n252 585
R71 B.n251 B.n250 585
R72 B.n249 B.n248 585
R73 B.n247 B.n246 585
R74 B.n245 B.n244 585
R75 B.n243 B.n242 585
R76 B.n241 B.n240 585
R77 B.n239 B.n238 585
R78 B.n237 B.n236 585
R79 B.n235 B.n234 585
R80 B.n233 B.n232 585
R81 B.n231 B.n230 585
R82 B.n229 B.n228 585
R83 B.n227 B.n226 585
R84 B.n225 B.n224 585
R85 B.n223 B.n222 585
R86 B.n221 B.n220 585
R87 B.n219 B.n218 585
R88 B.n217 B.n216 585
R89 B.n215 B.n214 585
R90 B.n213 B.n212 585
R91 B.n211 B.n210 585
R92 B.n209 B.n208 585
R93 B.n207 B.n206 585
R94 B.n205 B.n204 585
R95 B.n203 B.n202 585
R96 B.n201 B.n200 585
R97 B.n199 B.n198 585
R98 B.n197 B.n196 585
R99 B.n195 B.n194 585
R100 B.n193 B.n192 585
R101 B.n191 B.n190 585
R102 B.n189 B.n188 585
R103 B.n187 B.n186 585
R104 B.n185 B.n184 585
R105 B.n183 B.n182 585
R106 B.n181 B.n180 585
R107 B.n179 B.n178 585
R108 B.n177 B.n176 585
R109 B.n175 B.n174 585
R110 B.n172 B.n171 585
R111 B.n170 B.n169 585
R112 B.n168 B.n167 585
R113 B.n166 B.n165 585
R114 B.n164 B.n163 585
R115 B.n162 B.n161 585
R116 B.n160 B.n159 585
R117 B.n158 B.n157 585
R118 B.n156 B.n155 585
R119 B.n154 B.n153 585
R120 B.n152 B.n151 585
R121 B.n150 B.n149 585
R122 B.n148 B.n147 585
R123 B.n146 B.n145 585
R124 B.n144 B.n143 585
R125 B.n142 B.n141 585
R126 B.n140 B.n139 585
R127 B.n138 B.n137 585
R128 B.n136 B.n135 585
R129 B.n134 B.n133 585
R130 B.n132 B.n131 585
R131 B.n130 B.n129 585
R132 B.n128 B.n127 585
R133 B.n126 B.n125 585
R134 B.n124 B.n123 585
R135 B.n122 B.n121 585
R136 B.n120 B.n119 585
R137 B.n118 B.n117 585
R138 B.n116 B.n115 585
R139 B.n114 B.n113 585
R140 B.n112 B.n111 585
R141 B.n110 B.n109 585
R142 B.n108 B.n107 585
R143 B.n106 B.n105 585
R144 B.n104 B.n103 585
R145 B.n102 B.n101 585
R146 B.n100 B.n99 585
R147 B.n98 B.n97 585
R148 B.n96 B.n95 585
R149 B.n94 B.n93 585
R150 B.n92 B.n91 585
R151 B.n90 B.n89 585
R152 B.n88 B.n87 585
R153 B.n31 B.n30 585
R154 B.n631 B.n630 585
R155 B.n625 B.n81 585
R156 B.n81 B.n28 585
R157 B.n624 B.n27 585
R158 B.n635 B.n27 585
R159 B.n623 B.n26 585
R160 B.n636 B.n26 585
R161 B.n622 B.n25 585
R162 B.n637 B.n25 585
R163 B.n621 B.n620 585
R164 B.n620 B.t11 585
R165 B.n619 B.n21 585
R166 B.n643 B.n21 585
R167 B.n618 B.n20 585
R168 B.n644 B.n20 585
R169 B.n617 B.n19 585
R170 B.n645 B.n19 585
R171 B.n616 B.n615 585
R172 B.n615 B.n15 585
R173 B.n614 B.n14 585
R174 B.n651 B.n14 585
R175 B.n613 B.n13 585
R176 B.n652 B.n13 585
R177 B.n612 B.n12 585
R178 B.n653 B.n12 585
R179 B.n611 B.n610 585
R180 B.n610 B.n609 585
R181 B.n608 B.n607 585
R182 B.n608 B.n8 585
R183 B.n606 B.n7 585
R184 B.n660 B.n7 585
R185 B.n605 B.n6 585
R186 B.n661 B.n6 585
R187 B.n604 B.n5 585
R188 B.n662 B.n5 585
R189 B.n603 B.n602 585
R190 B.n602 B.n4 585
R191 B.n601 B.n279 585
R192 B.n601 B.n600 585
R193 B.n590 B.n280 585
R194 B.n593 B.n280 585
R195 B.n592 B.n591 585
R196 B.n594 B.n592 585
R197 B.n589 B.n285 585
R198 B.n285 B.n284 585
R199 B.n588 B.n587 585
R200 B.n587 B.n586 585
R201 B.n287 B.n286 585
R202 B.n288 B.n287 585
R203 B.n579 B.n578 585
R204 B.n580 B.n579 585
R205 B.n577 B.n293 585
R206 B.n293 B.n292 585
R207 B.n576 B.n575 585
R208 B.n575 B.n574 585
R209 B.n295 B.n294 585
R210 B.t7 B.n295 585
R211 B.n567 B.n566 585
R212 B.n568 B.n567 585
R213 B.n565 B.n300 585
R214 B.n300 B.n299 585
R215 B.n564 B.n563 585
R216 B.n563 B.n562 585
R217 B.n302 B.n301 585
R218 B.n303 B.n302 585
R219 B.n558 B.n557 585
R220 B.n306 B.n305 585
R221 B.n554 B.n553 585
R222 B.n555 B.n554 585
R223 B.n552 B.n355 585
R224 B.n551 B.n550 585
R225 B.n549 B.n548 585
R226 B.n547 B.n546 585
R227 B.n545 B.n544 585
R228 B.n543 B.n542 585
R229 B.n541 B.n540 585
R230 B.n539 B.n538 585
R231 B.n537 B.n536 585
R232 B.n535 B.n534 585
R233 B.n533 B.n532 585
R234 B.n531 B.n530 585
R235 B.n529 B.n528 585
R236 B.n527 B.n526 585
R237 B.n525 B.n524 585
R238 B.n523 B.n522 585
R239 B.n521 B.n520 585
R240 B.n519 B.n518 585
R241 B.n517 B.n516 585
R242 B.n515 B.n514 585
R243 B.n513 B.n512 585
R244 B.n511 B.n510 585
R245 B.n509 B.n508 585
R246 B.n507 B.n506 585
R247 B.n505 B.n504 585
R248 B.n503 B.n502 585
R249 B.n501 B.n500 585
R250 B.n499 B.n498 585
R251 B.n497 B.n496 585
R252 B.n495 B.n494 585
R253 B.n493 B.n492 585
R254 B.n491 B.n490 585
R255 B.n489 B.n488 585
R256 B.n487 B.n486 585
R257 B.n485 B.n484 585
R258 B.n483 B.n482 585
R259 B.n481 B.n480 585
R260 B.n479 B.n478 585
R261 B.n477 B.n476 585
R262 B.n475 B.n474 585
R263 B.n473 B.n472 585
R264 B.n471 B.n470 585
R265 B.n469 B.n468 585
R266 B.n467 B.n466 585
R267 B.n465 B.n464 585
R268 B.n463 B.n462 585
R269 B.n461 B.n460 585
R270 B.n459 B.n458 585
R271 B.n457 B.n456 585
R272 B.n455 B.n454 585
R273 B.n453 B.n452 585
R274 B.n450 B.n449 585
R275 B.n448 B.n447 585
R276 B.n446 B.n445 585
R277 B.n444 B.n443 585
R278 B.n442 B.n441 585
R279 B.n440 B.n439 585
R280 B.n438 B.n437 585
R281 B.n436 B.n435 585
R282 B.n434 B.n433 585
R283 B.n432 B.n431 585
R284 B.n430 B.n429 585
R285 B.n428 B.n427 585
R286 B.n426 B.n425 585
R287 B.n424 B.n423 585
R288 B.n422 B.n421 585
R289 B.n420 B.n419 585
R290 B.n418 B.n417 585
R291 B.n416 B.n415 585
R292 B.n414 B.n413 585
R293 B.n412 B.n411 585
R294 B.n410 B.n409 585
R295 B.n408 B.n407 585
R296 B.n406 B.n405 585
R297 B.n404 B.n403 585
R298 B.n402 B.n401 585
R299 B.n400 B.n399 585
R300 B.n398 B.n397 585
R301 B.n396 B.n395 585
R302 B.n394 B.n393 585
R303 B.n392 B.n391 585
R304 B.n390 B.n389 585
R305 B.n388 B.n387 585
R306 B.n386 B.n385 585
R307 B.n384 B.n383 585
R308 B.n382 B.n381 585
R309 B.n380 B.n379 585
R310 B.n378 B.n377 585
R311 B.n376 B.n375 585
R312 B.n374 B.n373 585
R313 B.n372 B.n371 585
R314 B.n370 B.n369 585
R315 B.n368 B.n367 585
R316 B.n366 B.n365 585
R317 B.n364 B.n363 585
R318 B.n362 B.n361 585
R319 B.n559 B.n304 585
R320 B.n304 B.n303 585
R321 B.n561 B.n560 585
R322 B.n562 B.n561 585
R323 B.n298 B.n297 585
R324 B.n299 B.n298 585
R325 B.n570 B.n569 585
R326 B.n569 B.n568 585
R327 B.n571 B.n296 585
R328 B.n296 B.t7 585
R329 B.n573 B.n572 585
R330 B.n574 B.n573 585
R331 B.n291 B.n290 585
R332 B.n292 B.n291 585
R333 B.n582 B.n581 585
R334 B.n581 B.n580 585
R335 B.n583 B.n289 585
R336 B.n289 B.n288 585
R337 B.n585 B.n584 585
R338 B.n586 B.n585 585
R339 B.n283 B.n282 585
R340 B.n284 B.n283 585
R341 B.n596 B.n595 585
R342 B.n595 B.n594 585
R343 B.n597 B.n281 585
R344 B.n593 B.n281 585
R345 B.n599 B.n598 585
R346 B.n600 B.n599 585
R347 B.n3 B.n0 585
R348 B.n4 B.n3 585
R349 B.n659 B.n1 585
R350 B.n660 B.n659 585
R351 B.n658 B.n657 585
R352 B.n658 B.n8 585
R353 B.n656 B.n9 585
R354 B.n609 B.n9 585
R355 B.n655 B.n654 585
R356 B.n654 B.n653 585
R357 B.n11 B.n10 585
R358 B.n652 B.n11 585
R359 B.n650 B.n649 585
R360 B.n651 B.n650 585
R361 B.n648 B.n16 585
R362 B.n16 B.n15 585
R363 B.n647 B.n646 585
R364 B.n646 B.n645 585
R365 B.n18 B.n17 585
R366 B.n644 B.n18 585
R367 B.n642 B.n641 585
R368 B.n643 B.n642 585
R369 B.n640 B.n22 585
R370 B.n22 B.t11 585
R371 B.n639 B.n638 585
R372 B.n638 B.n637 585
R373 B.n24 B.n23 585
R374 B.n636 B.n24 585
R375 B.n634 B.n633 585
R376 B.n635 B.n634 585
R377 B.n632 B.n29 585
R378 B.n29 B.n28 585
R379 B.n663 B.n662 585
R380 B.n661 B.n2 585
R381 B.n630 B.n29 535.745
R382 B.n627 B.n81 535.745
R383 B.n361 B.n302 535.745
R384 B.n557 B.n304 535.745
R385 B.n628 B.n79 256.663
R386 B.n628 B.n78 256.663
R387 B.n628 B.n77 256.663
R388 B.n628 B.n76 256.663
R389 B.n628 B.n75 256.663
R390 B.n628 B.n74 256.663
R391 B.n628 B.n73 256.663
R392 B.n628 B.n72 256.663
R393 B.n628 B.n71 256.663
R394 B.n628 B.n70 256.663
R395 B.n628 B.n69 256.663
R396 B.n628 B.n68 256.663
R397 B.n628 B.n67 256.663
R398 B.n628 B.n66 256.663
R399 B.n628 B.n65 256.663
R400 B.n628 B.n64 256.663
R401 B.n628 B.n63 256.663
R402 B.n628 B.n62 256.663
R403 B.n628 B.n61 256.663
R404 B.n628 B.n60 256.663
R405 B.n628 B.n59 256.663
R406 B.n628 B.n58 256.663
R407 B.n628 B.n57 256.663
R408 B.n628 B.n56 256.663
R409 B.n628 B.n55 256.663
R410 B.n628 B.n54 256.663
R411 B.n628 B.n53 256.663
R412 B.n628 B.n52 256.663
R413 B.n628 B.n51 256.663
R414 B.n628 B.n50 256.663
R415 B.n628 B.n49 256.663
R416 B.n628 B.n48 256.663
R417 B.n628 B.n47 256.663
R418 B.n628 B.n46 256.663
R419 B.n628 B.n45 256.663
R420 B.n628 B.n44 256.663
R421 B.n628 B.n43 256.663
R422 B.n628 B.n42 256.663
R423 B.n628 B.n41 256.663
R424 B.n628 B.n40 256.663
R425 B.n628 B.n39 256.663
R426 B.n628 B.n38 256.663
R427 B.n628 B.n37 256.663
R428 B.n628 B.n36 256.663
R429 B.n628 B.n35 256.663
R430 B.n628 B.n34 256.663
R431 B.n628 B.n33 256.663
R432 B.n628 B.n32 256.663
R433 B.n629 B.n628 256.663
R434 B.n556 B.n555 256.663
R435 B.n555 B.n307 256.663
R436 B.n555 B.n308 256.663
R437 B.n555 B.n309 256.663
R438 B.n555 B.n310 256.663
R439 B.n555 B.n311 256.663
R440 B.n555 B.n312 256.663
R441 B.n555 B.n313 256.663
R442 B.n555 B.n314 256.663
R443 B.n555 B.n315 256.663
R444 B.n555 B.n316 256.663
R445 B.n555 B.n317 256.663
R446 B.n555 B.n318 256.663
R447 B.n555 B.n319 256.663
R448 B.n555 B.n320 256.663
R449 B.n555 B.n321 256.663
R450 B.n555 B.n322 256.663
R451 B.n555 B.n323 256.663
R452 B.n555 B.n324 256.663
R453 B.n555 B.n325 256.663
R454 B.n555 B.n326 256.663
R455 B.n555 B.n327 256.663
R456 B.n555 B.n328 256.663
R457 B.n555 B.n329 256.663
R458 B.n555 B.n330 256.663
R459 B.n555 B.n331 256.663
R460 B.n555 B.n332 256.663
R461 B.n555 B.n333 256.663
R462 B.n555 B.n334 256.663
R463 B.n555 B.n335 256.663
R464 B.n555 B.n336 256.663
R465 B.n555 B.n337 256.663
R466 B.n555 B.n338 256.663
R467 B.n555 B.n339 256.663
R468 B.n555 B.n340 256.663
R469 B.n555 B.n341 256.663
R470 B.n555 B.n342 256.663
R471 B.n555 B.n343 256.663
R472 B.n555 B.n344 256.663
R473 B.n555 B.n345 256.663
R474 B.n555 B.n346 256.663
R475 B.n555 B.n347 256.663
R476 B.n555 B.n348 256.663
R477 B.n555 B.n349 256.663
R478 B.n555 B.n350 256.663
R479 B.n555 B.n351 256.663
R480 B.n555 B.n352 256.663
R481 B.n555 B.n353 256.663
R482 B.n555 B.n354 256.663
R483 B.n665 B.n664 256.663
R484 B.n87 B.n31 163.367
R485 B.n91 B.n90 163.367
R486 B.n95 B.n94 163.367
R487 B.n99 B.n98 163.367
R488 B.n103 B.n102 163.367
R489 B.n107 B.n106 163.367
R490 B.n111 B.n110 163.367
R491 B.n115 B.n114 163.367
R492 B.n119 B.n118 163.367
R493 B.n123 B.n122 163.367
R494 B.n127 B.n126 163.367
R495 B.n131 B.n130 163.367
R496 B.n135 B.n134 163.367
R497 B.n139 B.n138 163.367
R498 B.n143 B.n142 163.367
R499 B.n147 B.n146 163.367
R500 B.n151 B.n150 163.367
R501 B.n155 B.n154 163.367
R502 B.n159 B.n158 163.367
R503 B.n163 B.n162 163.367
R504 B.n167 B.n166 163.367
R505 B.n171 B.n170 163.367
R506 B.n176 B.n175 163.367
R507 B.n180 B.n179 163.367
R508 B.n184 B.n183 163.367
R509 B.n188 B.n187 163.367
R510 B.n192 B.n191 163.367
R511 B.n196 B.n195 163.367
R512 B.n200 B.n199 163.367
R513 B.n204 B.n203 163.367
R514 B.n208 B.n207 163.367
R515 B.n212 B.n211 163.367
R516 B.n216 B.n215 163.367
R517 B.n220 B.n219 163.367
R518 B.n224 B.n223 163.367
R519 B.n228 B.n227 163.367
R520 B.n232 B.n231 163.367
R521 B.n236 B.n235 163.367
R522 B.n240 B.n239 163.367
R523 B.n244 B.n243 163.367
R524 B.n248 B.n247 163.367
R525 B.n252 B.n251 163.367
R526 B.n256 B.n255 163.367
R527 B.n260 B.n259 163.367
R528 B.n264 B.n263 163.367
R529 B.n268 B.n267 163.367
R530 B.n272 B.n271 163.367
R531 B.n276 B.n275 163.367
R532 B.n627 B.n80 163.367
R533 B.n563 B.n302 163.367
R534 B.n563 B.n300 163.367
R535 B.n567 B.n300 163.367
R536 B.n567 B.n295 163.367
R537 B.n575 B.n295 163.367
R538 B.n575 B.n293 163.367
R539 B.n579 B.n293 163.367
R540 B.n579 B.n287 163.367
R541 B.n587 B.n287 163.367
R542 B.n587 B.n285 163.367
R543 B.n592 B.n285 163.367
R544 B.n592 B.n280 163.367
R545 B.n601 B.n280 163.367
R546 B.n602 B.n601 163.367
R547 B.n602 B.n5 163.367
R548 B.n6 B.n5 163.367
R549 B.n7 B.n6 163.367
R550 B.n608 B.n7 163.367
R551 B.n610 B.n608 163.367
R552 B.n610 B.n12 163.367
R553 B.n13 B.n12 163.367
R554 B.n14 B.n13 163.367
R555 B.n615 B.n14 163.367
R556 B.n615 B.n19 163.367
R557 B.n20 B.n19 163.367
R558 B.n21 B.n20 163.367
R559 B.n620 B.n21 163.367
R560 B.n620 B.n25 163.367
R561 B.n26 B.n25 163.367
R562 B.n27 B.n26 163.367
R563 B.n81 B.n27 163.367
R564 B.n554 B.n306 163.367
R565 B.n554 B.n355 163.367
R566 B.n550 B.n549 163.367
R567 B.n546 B.n545 163.367
R568 B.n542 B.n541 163.367
R569 B.n538 B.n537 163.367
R570 B.n534 B.n533 163.367
R571 B.n530 B.n529 163.367
R572 B.n526 B.n525 163.367
R573 B.n522 B.n521 163.367
R574 B.n518 B.n517 163.367
R575 B.n514 B.n513 163.367
R576 B.n510 B.n509 163.367
R577 B.n506 B.n505 163.367
R578 B.n502 B.n501 163.367
R579 B.n498 B.n497 163.367
R580 B.n494 B.n493 163.367
R581 B.n490 B.n489 163.367
R582 B.n486 B.n485 163.367
R583 B.n482 B.n481 163.367
R584 B.n478 B.n477 163.367
R585 B.n474 B.n473 163.367
R586 B.n470 B.n469 163.367
R587 B.n466 B.n465 163.367
R588 B.n462 B.n461 163.367
R589 B.n458 B.n457 163.367
R590 B.n454 B.n453 163.367
R591 B.n449 B.n448 163.367
R592 B.n445 B.n444 163.367
R593 B.n441 B.n440 163.367
R594 B.n437 B.n436 163.367
R595 B.n433 B.n432 163.367
R596 B.n429 B.n428 163.367
R597 B.n425 B.n424 163.367
R598 B.n421 B.n420 163.367
R599 B.n417 B.n416 163.367
R600 B.n413 B.n412 163.367
R601 B.n409 B.n408 163.367
R602 B.n405 B.n404 163.367
R603 B.n401 B.n400 163.367
R604 B.n397 B.n396 163.367
R605 B.n393 B.n392 163.367
R606 B.n389 B.n388 163.367
R607 B.n385 B.n384 163.367
R608 B.n381 B.n380 163.367
R609 B.n377 B.n376 163.367
R610 B.n373 B.n372 163.367
R611 B.n369 B.n368 163.367
R612 B.n365 B.n364 163.367
R613 B.n561 B.n304 163.367
R614 B.n561 B.n298 163.367
R615 B.n569 B.n298 163.367
R616 B.n569 B.n296 163.367
R617 B.n573 B.n296 163.367
R618 B.n573 B.n291 163.367
R619 B.n581 B.n291 163.367
R620 B.n581 B.n289 163.367
R621 B.n585 B.n289 163.367
R622 B.n585 B.n283 163.367
R623 B.n595 B.n283 163.367
R624 B.n595 B.n281 163.367
R625 B.n599 B.n281 163.367
R626 B.n599 B.n3 163.367
R627 B.n663 B.n3 163.367
R628 B.n659 B.n2 163.367
R629 B.n659 B.n658 163.367
R630 B.n658 B.n9 163.367
R631 B.n654 B.n9 163.367
R632 B.n654 B.n11 163.367
R633 B.n650 B.n11 163.367
R634 B.n650 B.n16 163.367
R635 B.n646 B.n16 163.367
R636 B.n646 B.n18 163.367
R637 B.n642 B.n18 163.367
R638 B.n642 B.n22 163.367
R639 B.n638 B.n22 163.367
R640 B.n638 B.n24 163.367
R641 B.n634 B.n24 163.367
R642 B.n634 B.n29 163.367
R643 B.n555 B.n303 84.6852
R644 B.n628 B.n28 84.6852
R645 B.n82 B.t12 82.5931
R646 B.n359 B.t9 82.5931
R647 B.n85 B.t15 82.5764
R648 B.n356 B.t19 82.5764
R649 B.n630 B.n629 71.676
R650 B.n87 B.n32 71.676
R651 B.n91 B.n33 71.676
R652 B.n95 B.n34 71.676
R653 B.n99 B.n35 71.676
R654 B.n103 B.n36 71.676
R655 B.n107 B.n37 71.676
R656 B.n111 B.n38 71.676
R657 B.n115 B.n39 71.676
R658 B.n119 B.n40 71.676
R659 B.n123 B.n41 71.676
R660 B.n127 B.n42 71.676
R661 B.n131 B.n43 71.676
R662 B.n135 B.n44 71.676
R663 B.n139 B.n45 71.676
R664 B.n143 B.n46 71.676
R665 B.n147 B.n47 71.676
R666 B.n151 B.n48 71.676
R667 B.n155 B.n49 71.676
R668 B.n159 B.n50 71.676
R669 B.n163 B.n51 71.676
R670 B.n167 B.n52 71.676
R671 B.n171 B.n53 71.676
R672 B.n176 B.n54 71.676
R673 B.n180 B.n55 71.676
R674 B.n184 B.n56 71.676
R675 B.n188 B.n57 71.676
R676 B.n192 B.n58 71.676
R677 B.n196 B.n59 71.676
R678 B.n200 B.n60 71.676
R679 B.n204 B.n61 71.676
R680 B.n208 B.n62 71.676
R681 B.n212 B.n63 71.676
R682 B.n216 B.n64 71.676
R683 B.n220 B.n65 71.676
R684 B.n224 B.n66 71.676
R685 B.n228 B.n67 71.676
R686 B.n232 B.n68 71.676
R687 B.n236 B.n69 71.676
R688 B.n240 B.n70 71.676
R689 B.n244 B.n71 71.676
R690 B.n248 B.n72 71.676
R691 B.n252 B.n73 71.676
R692 B.n256 B.n74 71.676
R693 B.n260 B.n75 71.676
R694 B.n264 B.n76 71.676
R695 B.n268 B.n77 71.676
R696 B.n272 B.n78 71.676
R697 B.n276 B.n79 71.676
R698 B.n80 B.n79 71.676
R699 B.n275 B.n78 71.676
R700 B.n271 B.n77 71.676
R701 B.n267 B.n76 71.676
R702 B.n263 B.n75 71.676
R703 B.n259 B.n74 71.676
R704 B.n255 B.n73 71.676
R705 B.n251 B.n72 71.676
R706 B.n247 B.n71 71.676
R707 B.n243 B.n70 71.676
R708 B.n239 B.n69 71.676
R709 B.n235 B.n68 71.676
R710 B.n231 B.n67 71.676
R711 B.n227 B.n66 71.676
R712 B.n223 B.n65 71.676
R713 B.n219 B.n64 71.676
R714 B.n215 B.n63 71.676
R715 B.n211 B.n62 71.676
R716 B.n207 B.n61 71.676
R717 B.n203 B.n60 71.676
R718 B.n199 B.n59 71.676
R719 B.n195 B.n58 71.676
R720 B.n191 B.n57 71.676
R721 B.n187 B.n56 71.676
R722 B.n183 B.n55 71.676
R723 B.n179 B.n54 71.676
R724 B.n175 B.n53 71.676
R725 B.n170 B.n52 71.676
R726 B.n166 B.n51 71.676
R727 B.n162 B.n50 71.676
R728 B.n158 B.n49 71.676
R729 B.n154 B.n48 71.676
R730 B.n150 B.n47 71.676
R731 B.n146 B.n46 71.676
R732 B.n142 B.n45 71.676
R733 B.n138 B.n44 71.676
R734 B.n134 B.n43 71.676
R735 B.n130 B.n42 71.676
R736 B.n126 B.n41 71.676
R737 B.n122 B.n40 71.676
R738 B.n118 B.n39 71.676
R739 B.n114 B.n38 71.676
R740 B.n110 B.n37 71.676
R741 B.n106 B.n36 71.676
R742 B.n102 B.n35 71.676
R743 B.n98 B.n34 71.676
R744 B.n94 B.n33 71.676
R745 B.n90 B.n32 71.676
R746 B.n629 B.n31 71.676
R747 B.n557 B.n556 71.676
R748 B.n355 B.n307 71.676
R749 B.n549 B.n308 71.676
R750 B.n545 B.n309 71.676
R751 B.n541 B.n310 71.676
R752 B.n537 B.n311 71.676
R753 B.n533 B.n312 71.676
R754 B.n529 B.n313 71.676
R755 B.n525 B.n314 71.676
R756 B.n521 B.n315 71.676
R757 B.n517 B.n316 71.676
R758 B.n513 B.n317 71.676
R759 B.n509 B.n318 71.676
R760 B.n505 B.n319 71.676
R761 B.n501 B.n320 71.676
R762 B.n497 B.n321 71.676
R763 B.n493 B.n322 71.676
R764 B.n489 B.n323 71.676
R765 B.n485 B.n324 71.676
R766 B.n481 B.n325 71.676
R767 B.n477 B.n326 71.676
R768 B.n473 B.n327 71.676
R769 B.n469 B.n328 71.676
R770 B.n465 B.n329 71.676
R771 B.n461 B.n330 71.676
R772 B.n457 B.n331 71.676
R773 B.n453 B.n332 71.676
R774 B.n448 B.n333 71.676
R775 B.n444 B.n334 71.676
R776 B.n440 B.n335 71.676
R777 B.n436 B.n336 71.676
R778 B.n432 B.n337 71.676
R779 B.n428 B.n338 71.676
R780 B.n424 B.n339 71.676
R781 B.n420 B.n340 71.676
R782 B.n416 B.n341 71.676
R783 B.n412 B.n342 71.676
R784 B.n408 B.n343 71.676
R785 B.n404 B.n344 71.676
R786 B.n400 B.n345 71.676
R787 B.n396 B.n346 71.676
R788 B.n392 B.n347 71.676
R789 B.n388 B.n348 71.676
R790 B.n384 B.n349 71.676
R791 B.n380 B.n350 71.676
R792 B.n376 B.n351 71.676
R793 B.n372 B.n352 71.676
R794 B.n368 B.n353 71.676
R795 B.n364 B.n354 71.676
R796 B.n556 B.n306 71.676
R797 B.n550 B.n307 71.676
R798 B.n546 B.n308 71.676
R799 B.n542 B.n309 71.676
R800 B.n538 B.n310 71.676
R801 B.n534 B.n311 71.676
R802 B.n530 B.n312 71.676
R803 B.n526 B.n313 71.676
R804 B.n522 B.n314 71.676
R805 B.n518 B.n315 71.676
R806 B.n514 B.n316 71.676
R807 B.n510 B.n317 71.676
R808 B.n506 B.n318 71.676
R809 B.n502 B.n319 71.676
R810 B.n498 B.n320 71.676
R811 B.n494 B.n321 71.676
R812 B.n490 B.n322 71.676
R813 B.n486 B.n323 71.676
R814 B.n482 B.n324 71.676
R815 B.n478 B.n325 71.676
R816 B.n474 B.n326 71.676
R817 B.n470 B.n327 71.676
R818 B.n466 B.n328 71.676
R819 B.n462 B.n329 71.676
R820 B.n458 B.n330 71.676
R821 B.n454 B.n331 71.676
R822 B.n449 B.n332 71.676
R823 B.n445 B.n333 71.676
R824 B.n441 B.n334 71.676
R825 B.n437 B.n335 71.676
R826 B.n433 B.n336 71.676
R827 B.n429 B.n337 71.676
R828 B.n425 B.n338 71.676
R829 B.n421 B.n339 71.676
R830 B.n417 B.n340 71.676
R831 B.n413 B.n341 71.676
R832 B.n409 B.n342 71.676
R833 B.n405 B.n343 71.676
R834 B.n401 B.n344 71.676
R835 B.n397 B.n345 71.676
R836 B.n393 B.n346 71.676
R837 B.n389 B.n347 71.676
R838 B.n385 B.n348 71.676
R839 B.n381 B.n349 71.676
R840 B.n377 B.n350 71.676
R841 B.n373 B.n351 71.676
R842 B.n369 B.n352 71.676
R843 B.n365 B.n353 71.676
R844 B.n361 B.n354 71.676
R845 B.n664 B.n663 71.676
R846 B.n664 B.n2 71.676
R847 B.n83 B.t13 69.9871
R848 B.n360 B.t8 69.9871
R849 B.n86 B.t16 69.9703
R850 B.n357 B.t18 69.9703
R851 B.n173 B.n86 59.5399
R852 B.n84 B.n83 59.5399
R853 B.n451 B.n360 59.5399
R854 B.n358 B.n357 59.5399
R855 B.n562 B.n303 40.8413
R856 B.n562 B.n299 40.8413
R857 B.n568 B.n299 40.8413
R858 B.n568 B.t7 40.8413
R859 B.n574 B.t7 40.8413
R860 B.n574 B.n292 40.8413
R861 B.n580 B.n292 40.8413
R862 B.n580 B.n288 40.8413
R863 B.n586 B.n288 40.8413
R864 B.n594 B.n284 40.8413
R865 B.n600 B.n4 40.8413
R866 B.n662 B.n4 40.8413
R867 B.n662 B.n661 40.8413
R868 B.n661 B.n660 40.8413
R869 B.n660 B.n8 40.8413
R870 B.n653 B.n652 40.8413
R871 B.n651 B.n15 40.8413
R872 B.n645 B.n15 40.8413
R873 B.n645 B.n644 40.8413
R874 B.n644 B.n643 40.8413
R875 B.n643 B.t11 40.8413
R876 B.n637 B.t11 40.8413
R877 B.n637 B.n636 40.8413
R878 B.n636 B.n635 40.8413
R879 B.n635 B.n28 40.8413
R880 B.t4 B.n593 39.6401
R881 B.n609 B.t0 39.6401
R882 B.n593 B.t2 38.4389
R883 B.n609 B.t1 38.4389
R884 B.t3 B.n284 36.0365
R885 B.n652 B.t5 36.0365
R886 B.n559 B.n558 34.8103
R887 B.n362 B.n301 34.8103
R888 B.n626 B.n625 34.8103
R889 B.n632 B.n631 34.8103
R890 B B.n665 18.0485
R891 B.n86 B.n85 12.6066
R892 B.n83 B.n82 12.6066
R893 B.n360 B.n359 12.6066
R894 B.n357 B.n356 12.6066
R895 B.n560 B.n559 10.6151
R896 B.n560 B.n297 10.6151
R897 B.n570 B.n297 10.6151
R898 B.n571 B.n570 10.6151
R899 B.n572 B.n571 10.6151
R900 B.n572 B.n290 10.6151
R901 B.n582 B.n290 10.6151
R902 B.n583 B.n582 10.6151
R903 B.n584 B.n583 10.6151
R904 B.n584 B.n282 10.6151
R905 B.n596 B.n282 10.6151
R906 B.n597 B.n596 10.6151
R907 B.n598 B.n597 10.6151
R908 B.n598 B.n0 10.6151
R909 B.n558 B.n305 10.6151
R910 B.n553 B.n305 10.6151
R911 B.n553 B.n552 10.6151
R912 B.n552 B.n551 10.6151
R913 B.n551 B.n548 10.6151
R914 B.n548 B.n547 10.6151
R915 B.n547 B.n544 10.6151
R916 B.n544 B.n543 10.6151
R917 B.n543 B.n540 10.6151
R918 B.n540 B.n539 10.6151
R919 B.n539 B.n536 10.6151
R920 B.n536 B.n535 10.6151
R921 B.n535 B.n532 10.6151
R922 B.n532 B.n531 10.6151
R923 B.n531 B.n528 10.6151
R924 B.n528 B.n527 10.6151
R925 B.n527 B.n524 10.6151
R926 B.n524 B.n523 10.6151
R927 B.n523 B.n520 10.6151
R928 B.n520 B.n519 10.6151
R929 B.n519 B.n516 10.6151
R930 B.n516 B.n515 10.6151
R931 B.n515 B.n512 10.6151
R932 B.n512 B.n511 10.6151
R933 B.n511 B.n508 10.6151
R934 B.n508 B.n507 10.6151
R935 B.n507 B.n504 10.6151
R936 B.n504 B.n503 10.6151
R937 B.n503 B.n500 10.6151
R938 B.n500 B.n499 10.6151
R939 B.n499 B.n496 10.6151
R940 B.n496 B.n495 10.6151
R941 B.n495 B.n492 10.6151
R942 B.n492 B.n491 10.6151
R943 B.n491 B.n488 10.6151
R944 B.n488 B.n487 10.6151
R945 B.n487 B.n484 10.6151
R946 B.n484 B.n483 10.6151
R947 B.n483 B.n480 10.6151
R948 B.n480 B.n479 10.6151
R949 B.n479 B.n476 10.6151
R950 B.n476 B.n475 10.6151
R951 B.n475 B.n472 10.6151
R952 B.n472 B.n471 10.6151
R953 B.n468 B.n467 10.6151
R954 B.n467 B.n464 10.6151
R955 B.n464 B.n463 10.6151
R956 B.n463 B.n460 10.6151
R957 B.n460 B.n459 10.6151
R958 B.n459 B.n456 10.6151
R959 B.n456 B.n455 10.6151
R960 B.n455 B.n452 10.6151
R961 B.n450 B.n447 10.6151
R962 B.n447 B.n446 10.6151
R963 B.n446 B.n443 10.6151
R964 B.n443 B.n442 10.6151
R965 B.n442 B.n439 10.6151
R966 B.n439 B.n438 10.6151
R967 B.n438 B.n435 10.6151
R968 B.n435 B.n434 10.6151
R969 B.n434 B.n431 10.6151
R970 B.n431 B.n430 10.6151
R971 B.n430 B.n427 10.6151
R972 B.n427 B.n426 10.6151
R973 B.n426 B.n423 10.6151
R974 B.n423 B.n422 10.6151
R975 B.n422 B.n419 10.6151
R976 B.n419 B.n418 10.6151
R977 B.n418 B.n415 10.6151
R978 B.n415 B.n414 10.6151
R979 B.n414 B.n411 10.6151
R980 B.n411 B.n410 10.6151
R981 B.n410 B.n407 10.6151
R982 B.n407 B.n406 10.6151
R983 B.n406 B.n403 10.6151
R984 B.n403 B.n402 10.6151
R985 B.n402 B.n399 10.6151
R986 B.n399 B.n398 10.6151
R987 B.n398 B.n395 10.6151
R988 B.n395 B.n394 10.6151
R989 B.n394 B.n391 10.6151
R990 B.n391 B.n390 10.6151
R991 B.n390 B.n387 10.6151
R992 B.n387 B.n386 10.6151
R993 B.n386 B.n383 10.6151
R994 B.n383 B.n382 10.6151
R995 B.n382 B.n379 10.6151
R996 B.n379 B.n378 10.6151
R997 B.n378 B.n375 10.6151
R998 B.n375 B.n374 10.6151
R999 B.n374 B.n371 10.6151
R1000 B.n371 B.n370 10.6151
R1001 B.n370 B.n367 10.6151
R1002 B.n367 B.n366 10.6151
R1003 B.n366 B.n363 10.6151
R1004 B.n363 B.n362 10.6151
R1005 B.n564 B.n301 10.6151
R1006 B.n565 B.n564 10.6151
R1007 B.n566 B.n565 10.6151
R1008 B.n566 B.n294 10.6151
R1009 B.n576 B.n294 10.6151
R1010 B.n577 B.n576 10.6151
R1011 B.n578 B.n577 10.6151
R1012 B.n578 B.n286 10.6151
R1013 B.n588 B.n286 10.6151
R1014 B.n589 B.n588 10.6151
R1015 B.n591 B.n589 10.6151
R1016 B.n591 B.n590 10.6151
R1017 B.n590 B.n279 10.6151
R1018 B.n603 B.n279 10.6151
R1019 B.n604 B.n603 10.6151
R1020 B.n605 B.n604 10.6151
R1021 B.n606 B.n605 10.6151
R1022 B.n607 B.n606 10.6151
R1023 B.n611 B.n607 10.6151
R1024 B.n612 B.n611 10.6151
R1025 B.n613 B.n612 10.6151
R1026 B.n614 B.n613 10.6151
R1027 B.n616 B.n614 10.6151
R1028 B.n617 B.n616 10.6151
R1029 B.n618 B.n617 10.6151
R1030 B.n619 B.n618 10.6151
R1031 B.n621 B.n619 10.6151
R1032 B.n622 B.n621 10.6151
R1033 B.n623 B.n622 10.6151
R1034 B.n624 B.n623 10.6151
R1035 B.n625 B.n624 10.6151
R1036 B.n657 B.n1 10.6151
R1037 B.n657 B.n656 10.6151
R1038 B.n656 B.n655 10.6151
R1039 B.n655 B.n10 10.6151
R1040 B.n649 B.n10 10.6151
R1041 B.n649 B.n648 10.6151
R1042 B.n648 B.n647 10.6151
R1043 B.n647 B.n17 10.6151
R1044 B.n641 B.n17 10.6151
R1045 B.n641 B.n640 10.6151
R1046 B.n640 B.n639 10.6151
R1047 B.n639 B.n23 10.6151
R1048 B.n633 B.n23 10.6151
R1049 B.n633 B.n632 10.6151
R1050 B.n631 B.n30 10.6151
R1051 B.n88 B.n30 10.6151
R1052 B.n89 B.n88 10.6151
R1053 B.n92 B.n89 10.6151
R1054 B.n93 B.n92 10.6151
R1055 B.n96 B.n93 10.6151
R1056 B.n97 B.n96 10.6151
R1057 B.n100 B.n97 10.6151
R1058 B.n101 B.n100 10.6151
R1059 B.n104 B.n101 10.6151
R1060 B.n105 B.n104 10.6151
R1061 B.n108 B.n105 10.6151
R1062 B.n109 B.n108 10.6151
R1063 B.n112 B.n109 10.6151
R1064 B.n113 B.n112 10.6151
R1065 B.n116 B.n113 10.6151
R1066 B.n117 B.n116 10.6151
R1067 B.n120 B.n117 10.6151
R1068 B.n121 B.n120 10.6151
R1069 B.n124 B.n121 10.6151
R1070 B.n125 B.n124 10.6151
R1071 B.n128 B.n125 10.6151
R1072 B.n129 B.n128 10.6151
R1073 B.n132 B.n129 10.6151
R1074 B.n133 B.n132 10.6151
R1075 B.n136 B.n133 10.6151
R1076 B.n137 B.n136 10.6151
R1077 B.n140 B.n137 10.6151
R1078 B.n141 B.n140 10.6151
R1079 B.n144 B.n141 10.6151
R1080 B.n145 B.n144 10.6151
R1081 B.n148 B.n145 10.6151
R1082 B.n149 B.n148 10.6151
R1083 B.n152 B.n149 10.6151
R1084 B.n153 B.n152 10.6151
R1085 B.n156 B.n153 10.6151
R1086 B.n157 B.n156 10.6151
R1087 B.n160 B.n157 10.6151
R1088 B.n161 B.n160 10.6151
R1089 B.n164 B.n161 10.6151
R1090 B.n165 B.n164 10.6151
R1091 B.n168 B.n165 10.6151
R1092 B.n169 B.n168 10.6151
R1093 B.n172 B.n169 10.6151
R1094 B.n177 B.n174 10.6151
R1095 B.n178 B.n177 10.6151
R1096 B.n181 B.n178 10.6151
R1097 B.n182 B.n181 10.6151
R1098 B.n185 B.n182 10.6151
R1099 B.n186 B.n185 10.6151
R1100 B.n189 B.n186 10.6151
R1101 B.n190 B.n189 10.6151
R1102 B.n194 B.n193 10.6151
R1103 B.n197 B.n194 10.6151
R1104 B.n198 B.n197 10.6151
R1105 B.n201 B.n198 10.6151
R1106 B.n202 B.n201 10.6151
R1107 B.n205 B.n202 10.6151
R1108 B.n206 B.n205 10.6151
R1109 B.n209 B.n206 10.6151
R1110 B.n210 B.n209 10.6151
R1111 B.n213 B.n210 10.6151
R1112 B.n214 B.n213 10.6151
R1113 B.n217 B.n214 10.6151
R1114 B.n218 B.n217 10.6151
R1115 B.n221 B.n218 10.6151
R1116 B.n222 B.n221 10.6151
R1117 B.n225 B.n222 10.6151
R1118 B.n226 B.n225 10.6151
R1119 B.n229 B.n226 10.6151
R1120 B.n230 B.n229 10.6151
R1121 B.n233 B.n230 10.6151
R1122 B.n234 B.n233 10.6151
R1123 B.n237 B.n234 10.6151
R1124 B.n238 B.n237 10.6151
R1125 B.n241 B.n238 10.6151
R1126 B.n242 B.n241 10.6151
R1127 B.n245 B.n242 10.6151
R1128 B.n246 B.n245 10.6151
R1129 B.n249 B.n246 10.6151
R1130 B.n250 B.n249 10.6151
R1131 B.n253 B.n250 10.6151
R1132 B.n254 B.n253 10.6151
R1133 B.n257 B.n254 10.6151
R1134 B.n258 B.n257 10.6151
R1135 B.n261 B.n258 10.6151
R1136 B.n262 B.n261 10.6151
R1137 B.n265 B.n262 10.6151
R1138 B.n266 B.n265 10.6151
R1139 B.n269 B.n266 10.6151
R1140 B.n270 B.n269 10.6151
R1141 B.n273 B.n270 10.6151
R1142 B.n274 B.n273 10.6151
R1143 B.n277 B.n274 10.6151
R1144 B.n278 B.n277 10.6151
R1145 B.n626 B.n278 10.6151
R1146 B.n665 B.n0 8.11757
R1147 B.n665 B.n1 8.11757
R1148 B.n468 B.n358 6.5566
R1149 B.n452 B.n451 6.5566
R1150 B.n174 B.n173 6.5566
R1151 B.n190 B.n84 6.5566
R1152 B.n586 B.t3 4.8053
R1153 B.t5 B.n651 4.8053
R1154 B.n471 B.n358 4.05904
R1155 B.n451 B.n450 4.05904
R1156 B.n173 B.n172 4.05904
R1157 B.n193 B.n84 4.05904
R1158 B.n600 B.t2 2.4029
R1159 B.t1 B.n8 2.4029
R1160 B.n594 B.t4 1.2017
R1161 B.n653 B.t0 1.2017
R1162 VP.n1 VP.t5 1131.69
R1163 VP.n8 VP.t0 1101.89
R1164 VP.n6 VP.t2 1101.89
R1165 VP.n3 VP.t3 1101.89
R1166 VP.n7 VP.t1 1079.98
R1167 VP.n2 VP.t4 1079.98
R1168 VP.n9 VP.n8 161.3
R1169 VP.n4 VP.n3 161.3
R1170 VP.n7 VP.n0 161.3
R1171 VP.n6 VP.n5 161.3
R1172 VP.n7 VP.n6 73.0308
R1173 VP.n8 VP.n7 73.0308
R1174 VP.n3 VP.n2 73.0308
R1175 VP.n4 VP.n1 65.9987
R1176 VP.n5 VP.n4 40.4967
R1177 VP.n2 VP.n1 29.7615
R1178 VP.n5 VP.n0 0.189894
R1179 VP.n9 VP.n0 0.189894
R1180 VP VP.n9 0.0516364
R1181 VDD1 VDD1.t0 67.0526
R1182 VDD1.n1 VDD1.t3 66.9379
R1183 VDD1.n1 VDD1.n0 65.1393
R1184 VDD1.n3 VDD1.n2 65.0546
R1185 VDD1.n3 VDD1.n1 37.641
R1186 VDD1.n2 VDD1.t1 1.5189
R1187 VDD1.n2 VDD1.t2 1.5189
R1188 VDD1.n0 VDD1.t4 1.5189
R1189 VDD1.n0 VDD1.t5 1.5189
R1190 VDD1 VDD1.n3 0.0823966
C0 VTAIL VN 2.5312f
C1 VTAIL VDD1 14.6138f
C2 VDD2 VP 0.266198f
C3 VDD2 VN 3.03178f
C4 VDD2 VDD1 0.578066f
C5 VN VP 4.90503f
C6 VDD1 VP 3.14447f
C7 VDD2 VTAIL 14.642799f
C8 VN VDD1 0.148008f
C9 VTAIL VP 2.54601f
C10 VDD2 B 4.396122f
C11 VDD1 B 4.60187f
C12 VTAIL B 6.394814f
C13 VN B 7.00615f
C14 VP B 4.687886f
C15 VDD1.t0 B 3.23523f
C16 VDD1.t3 B 3.2346f
C17 VDD1.t4 B 0.281734f
C18 VDD1.t5 B 0.281734f
C19 VDD1.n0 B 2.5337f
C20 VDD1.n1 B 2.22307f
C21 VDD1.t1 B 0.281734f
C22 VDD1.t2 B 0.281734f
C23 VDD1.n2 B 2.53331f
C24 VDD1.n3 B 2.42718f
C25 VP.n0 B 0.057307f
C26 VP.t1 B 0.675299f
C27 VP.t2 B 0.680513f
C28 VP.t5 B 0.687923f
C29 VP.n1 B 0.274362f
C30 VP.t4 B 0.675299f
C31 VP.n2 B 0.282334f
C32 VP.t3 B 0.680513f
C33 VP.n3 B 0.281359f
C34 VP.n4 B 2.3427f
C35 VP.n5 B 2.27528f
C36 VP.n6 B 0.281359f
C37 VP.n7 B 0.282334f
C38 VP.t0 B 0.680513f
C39 VP.n8 B 0.281359f
C40 VP.n9 B 0.044411f
C41 VDD2.t5 B 3.23478f
C42 VDD2.t4 B 0.281749f
C43 VDD2.t3 B 0.281749f
C44 VDD2.n0 B 2.53384f
C45 VDD2.n1 B 2.14814f
C46 VDD2.t0 B 3.23299f
C47 VDD2.n2 B 2.45583f
C48 VDD2.t2 B 0.281749f
C49 VDD2.t1 B 0.281749f
C50 VDD2.n3 B 2.53381f
C51 VTAIL.t9 B 0.288181f
C52 VTAIL.t7 B 0.288181f
C53 VTAIL.n0 B 2.5166f
C54 VTAIL.n1 B 0.34409f
C55 VTAIL.t2 B 3.21081f
C56 VTAIL.n2 B 0.468456f
C57 VTAIL.t3 B 0.288181f
C58 VTAIL.t11 B 0.288181f
C59 VTAIL.n3 B 2.5166f
C60 VTAIL.n4 B 1.80301f
C61 VTAIL.t6 B 0.288181f
C62 VTAIL.t8 B 0.288181f
C63 VTAIL.n5 B 2.51661f
C64 VTAIL.n6 B 1.803f
C65 VTAIL.t5 B 3.21083f
C66 VTAIL.n7 B 0.468437f
C67 VTAIL.t1 B 0.288181f
C68 VTAIL.t0 B 0.288181f
C69 VTAIL.n8 B 2.51661f
C70 VTAIL.n9 B 0.376706f
C71 VTAIL.t10 B 3.21081f
C72 VTAIL.n10 B 1.84426f
C73 VTAIL.t4 B 3.21081f
C74 VTAIL.n11 B 1.82639f
C75 VN.t0 B 0.676184f
C76 VN.n0 B 0.26968f
C77 VN.t1 B 0.663775f
C78 VN.n1 B 0.277516f
C79 VN.t2 B 0.6689f
C80 VN.n2 B 0.276557f
C81 VN.n3 B 0.160073f
C82 VN.t4 B 0.676184f
C83 VN.n4 B 0.26968f
C84 VN.t5 B 0.6689f
C85 VN.t3 B 0.663775f
C86 VN.n5 B 0.277516f
C87 VN.n6 B 0.276557f
C88 VN.n7 B 2.33979f
.ends

