* NGSPICE file created from diff_pair_sample_0744.ext - technology: sky130A

.subckt diff_pair_sample_0744 VTAIL VN VP B VDD2 VDD1
X0 B.t19 B.t17 B.t18 B.t11 sky130_fd_pr__nfet_01v8 ad=2.652 pd=14.38 as=0 ps=0 w=6.8 l=1.28
X1 VDD1.t5 VP.t0 VTAIL.t10 B.t1 sky130_fd_pr__nfet_01v8 ad=1.122 pd=7.13 as=2.652 ps=14.38 w=6.8 l=1.28
X2 B.t16 B.t14 B.t15 B.t7 sky130_fd_pr__nfet_01v8 ad=2.652 pd=14.38 as=0 ps=0 w=6.8 l=1.28
X3 VTAIL.t1 VN.t0 VDD2.t5 B.t2 sky130_fd_pr__nfet_01v8 ad=1.122 pd=7.13 as=1.122 ps=7.13 w=6.8 l=1.28
X4 B.t13 B.t10 B.t12 B.t11 sky130_fd_pr__nfet_01v8 ad=2.652 pd=14.38 as=0 ps=0 w=6.8 l=1.28
X5 VDD2.t4 VN.t1 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=2.652 pd=14.38 as=1.122 ps=7.13 w=6.8 l=1.28
X6 B.t9 B.t6 B.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=2.652 pd=14.38 as=0 ps=0 w=6.8 l=1.28
X7 VDD1.t4 VP.t1 VTAIL.t6 B.t5 sky130_fd_pr__nfet_01v8 ad=2.652 pd=14.38 as=1.122 ps=7.13 w=6.8 l=1.28
X8 VDD2.t3 VN.t2 VTAIL.t2 B.t5 sky130_fd_pr__nfet_01v8 ad=2.652 pd=14.38 as=1.122 ps=7.13 w=6.8 l=1.28
X9 VTAIL.t3 VN.t3 VDD2.t2 B.t3 sky130_fd_pr__nfet_01v8 ad=1.122 pd=7.13 as=1.122 ps=7.13 w=6.8 l=1.28
X10 VDD2.t1 VN.t4 VTAIL.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=1.122 pd=7.13 as=2.652 ps=14.38 w=6.8 l=1.28
X11 VDD2.t0 VN.t5 VTAIL.t5 B.t1 sky130_fd_pr__nfet_01v8 ad=1.122 pd=7.13 as=2.652 ps=14.38 w=6.8 l=1.28
X12 VDD1.t3 VP.t2 VTAIL.t9 B.t0 sky130_fd_pr__nfet_01v8 ad=2.652 pd=14.38 as=1.122 ps=7.13 w=6.8 l=1.28
X13 VDD1.t2 VP.t3 VTAIL.t11 B.t4 sky130_fd_pr__nfet_01v8 ad=1.122 pd=7.13 as=2.652 ps=14.38 w=6.8 l=1.28
X14 VTAIL.t8 VP.t4 VDD1.t1 B.t3 sky130_fd_pr__nfet_01v8 ad=1.122 pd=7.13 as=1.122 ps=7.13 w=6.8 l=1.28
X15 VTAIL.t7 VP.t5 VDD1.t0 B.t2 sky130_fd_pr__nfet_01v8 ad=1.122 pd=7.13 as=1.122 ps=7.13 w=6.8 l=1.28
R0 B.n536 B.n535 585
R1 B.n207 B.n83 585
R2 B.n206 B.n205 585
R3 B.n204 B.n203 585
R4 B.n202 B.n201 585
R5 B.n200 B.n199 585
R6 B.n198 B.n197 585
R7 B.n196 B.n195 585
R8 B.n194 B.n193 585
R9 B.n192 B.n191 585
R10 B.n190 B.n189 585
R11 B.n188 B.n187 585
R12 B.n186 B.n185 585
R13 B.n184 B.n183 585
R14 B.n182 B.n181 585
R15 B.n180 B.n179 585
R16 B.n178 B.n177 585
R17 B.n176 B.n175 585
R18 B.n174 B.n173 585
R19 B.n172 B.n171 585
R20 B.n170 B.n169 585
R21 B.n168 B.n167 585
R22 B.n166 B.n165 585
R23 B.n164 B.n163 585
R24 B.n162 B.n161 585
R25 B.n160 B.n159 585
R26 B.n158 B.n157 585
R27 B.n156 B.n155 585
R28 B.n154 B.n153 585
R29 B.n152 B.n151 585
R30 B.n150 B.n149 585
R31 B.n148 B.n147 585
R32 B.n146 B.n145 585
R33 B.n144 B.n143 585
R34 B.n142 B.n141 585
R35 B.n140 B.n139 585
R36 B.n138 B.n137 585
R37 B.n136 B.n135 585
R38 B.n134 B.n133 585
R39 B.n132 B.n131 585
R40 B.n130 B.n129 585
R41 B.n128 B.n127 585
R42 B.n126 B.n125 585
R43 B.n124 B.n123 585
R44 B.n122 B.n121 585
R45 B.n120 B.n119 585
R46 B.n118 B.n117 585
R47 B.n116 B.n115 585
R48 B.n114 B.n113 585
R49 B.n112 B.n111 585
R50 B.n110 B.n109 585
R51 B.n108 B.n107 585
R52 B.n106 B.n105 585
R53 B.n104 B.n103 585
R54 B.n102 B.n101 585
R55 B.n100 B.n99 585
R56 B.n98 B.n97 585
R57 B.n96 B.n95 585
R58 B.n94 B.n93 585
R59 B.n92 B.n91 585
R60 B.n53 B.n52 585
R61 B.n541 B.n540 585
R62 B.n534 B.n84 585
R63 B.n84 B.n50 585
R64 B.n533 B.n49 585
R65 B.n545 B.n49 585
R66 B.n532 B.n48 585
R67 B.n546 B.n48 585
R68 B.n531 B.n47 585
R69 B.n547 B.n47 585
R70 B.n530 B.n529 585
R71 B.n529 B.n43 585
R72 B.n528 B.n42 585
R73 B.n553 B.n42 585
R74 B.n527 B.n41 585
R75 B.n554 B.n41 585
R76 B.n526 B.n40 585
R77 B.n555 B.n40 585
R78 B.n525 B.n524 585
R79 B.n524 B.n36 585
R80 B.n523 B.n35 585
R81 B.n561 B.n35 585
R82 B.n522 B.n34 585
R83 B.n562 B.n34 585
R84 B.n521 B.n33 585
R85 B.n563 B.n33 585
R86 B.n520 B.n519 585
R87 B.n519 B.n29 585
R88 B.n518 B.n28 585
R89 B.n569 B.n28 585
R90 B.n517 B.n27 585
R91 B.n570 B.n27 585
R92 B.n516 B.n26 585
R93 B.n571 B.n26 585
R94 B.n515 B.n514 585
R95 B.n514 B.n22 585
R96 B.n513 B.n21 585
R97 B.n577 B.n21 585
R98 B.n512 B.n20 585
R99 B.n578 B.n20 585
R100 B.n511 B.n19 585
R101 B.n579 B.n19 585
R102 B.n510 B.n509 585
R103 B.n509 B.n15 585
R104 B.n508 B.n14 585
R105 B.n585 B.n14 585
R106 B.n507 B.n13 585
R107 B.n586 B.n13 585
R108 B.n506 B.n12 585
R109 B.n587 B.n12 585
R110 B.n505 B.n504 585
R111 B.n504 B.n8 585
R112 B.n503 B.n7 585
R113 B.n593 B.n7 585
R114 B.n502 B.n6 585
R115 B.n594 B.n6 585
R116 B.n501 B.n5 585
R117 B.n595 B.n5 585
R118 B.n500 B.n499 585
R119 B.n499 B.n4 585
R120 B.n498 B.n208 585
R121 B.n498 B.n497 585
R122 B.n488 B.n209 585
R123 B.n210 B.n209 585
R124 B.n490 B.n489 585
R125 B.n491 B.n490 585
R126 B.n487 B.n215 585
R127 B.n215 B.n214 585
R128 B.n486 B.n485 585
R129 B.n485 B.n484 585
R130 B.n217 B.n216 585
R131 B.n218 B.n217 585
R132 B.n477 B.n476 585
R133 B.n478 B.n477 585
R134 B.n475 B.n222 585
R135 B.n226 B.n222 585
R136 B.n474 B.n473 585
R137 B.n473 B.n472 585
R138 B.n224 B.n223 585
R139 B.n225 B.n224 585
R140 B.n465 B.n464 585
R141 B.n466 B.n465 585
R142 B.n463 B.n231 585
R143 B.n231 B.n230 585
R144 B.n462 B.n461 585
R145 B.n461 B.n460 585
R146 B.n233 B.n232 585
R147 B.n234 B.n233 585
R148 B.n453 B.n452 585
R149 B.n454 B.n453 585
R150 B.n451 B.n239 585
R151 B.n239 B.n238 585
R152 B.n450 B.n449 585
R153 B.n449 B.n448 585
R154 B.n241 B.n240 585
R155 B.n242 B.n241 585
R156 B.n441 B.n440 585
R157 B.n442 B.n441 585
R158 B.n439 B.n247 585
R159 B.n247 B.n246 585
R160 B.n438 B.n437 585
R161 B.n437 B.n436 585
R162 B.n249 B.n248 585
R163 B.n250 B.n249 585
R164 B.n429 B.n428 585
R165 B.n430 B.n429 585
R166 B.n427 B.n255 585
R167 B.n255 B.n254 585
R168 B.n426 B.n425 585
R169 B.n425 B.n424 585
R170 B.n257 B.n256 585
R171 B.n258 B.n257 585
R172 B.n420 B.n419 585
R173 B.n261 B.n260 585
R174 B.n416 B.n415 585
R175 B.n417 B.n416 585
R176 B.n414 B.n292 585
R177 B.n413 B.n412 585
R178 B.n411 B.n410 585
R179 B.n409 B.n408 585
R180 B.n407 B.n406 585
R181 B.n405 B.n404 585
R182 B.n403 B.n402 585
R183 B.n401 B.n400 585
R184 B.n399 B.n398 585
R185 B.n397 B.n396 585
R186 B.n395 B.n394 585
R187 B.n393 B.n392 585
R188 B.n391 B.n390 585
R189 B.n389 B.n388 585
R190 B.n387 B.n386 585
R191 B.n385 B.n384 585
R192 B.n383 B.n382 585
R193 B.n381 B.n380 585
R194 B.n379 B.n378 585
R195 B.n377 B.n376 585
R196 B.n375 B.n374 585
R197 B.n373 B.n372 585
R198 B.n371 B.n370 585
R199 B.n368 B.n367 585
R200 B.n366 B.n365 585
R201 B.n364 B.n363 585
R202 B.n362 B.n361 585
R203 B.n360 B.n359 585
R204 B.n358 B.n357 585
R205 B.n356 B.n355 585
R206 B.n354 B.n353 585
R207 B.n352 B.n351 585
R208 B.n350 B.n349 585
R209 B.n347 B.n346 585
R210 B.n345 B.n344 585
R211 B.n343 B.n342 585
R212 B.n341 B.n340 585
R213 B.n339 B.n338 585
R214 B.n337 B.n336 585
R215 B.n335 B.n334 585
R216 B.n333 B.n332 585
R217 B.n331 B.n330 585
R218 B.n329 B.n328 585
R219 B.n327 B.n326 585
R220 B.n325 B.n324 585
R221 B.n323 B.n322 585
R222 B.n321 B.n320 585
R223 B.n319 B.n318 585
R224 B.n317 B.n316 585
R225 B.n315 B.n314 585
R226 B.n313 B.n312 585
R227 B.n311 B.n310 585
R228 B.n309 B.n308 585
R229 B.n307 B.n306 585
R230 B.n305 B.n304 585
R231 B.n303 B.n302 585
R232 B.n301 B.n300 585
R233 B.n299 B.n298 585
R234 B.n297 B.n291 585
R235 B.n417 B.n291 585
R236 B.n421 B.n259 585
R237 B.n259 B.n258 585
R238 B.n423 B.n422 585
R239 B.n424 B.n423 585
R240 B.n253 B.n252 585
R241 B.n254 B.n253 585
R242 B.n432 B.n431 585
R243 B.n431 B.n430 585
R244 B.n433 B.n251 585
R245 B.n251 B.n250 585
R246 B.n435 B.n434 585
R247 B.n436 B.n435 585
R248 B.n245 B.n244 585
R249 B.n246 B.n245 585
R250 B.n444 B.n443 585
R251 B.n443 B.n442 585
R252 B.n445 B.n243 585
R253 B.n243 B.n242 585
R254 B.n447 B.n446 585
R255 B.n448 B.n447 585
R256 B.n237 B.n236 585
R257 B.n238 B.n237 585
R258 B.n456 B.n455 585
R259 B.n455 B.n454 585
R260 B.n457 B.n235 585
R261 B.n235 B.n234 585
R262 B.n459 B.n458 585
R263 B.n460 B.n459 585
R264 B.n229 B.n228 585
R265 B.n230 B.n229 585
R266 B.n468 B.n467 585
R267 B.n467 B.n466 585
R268 B.n469 B.n227 585
R269 B.n227 B.n225 585
R270 B.n471 B.n470 585
R271 B.n472 B.n471 585
R272 B.n221 B.n220 585
R273 B.n226 B.n221 585
R274 B.n480 B.n479 585
R275 B.n479 B.n478 585
R276 B.n481 B.n219 585
R277 B.n219 B.n218 585
R278 B.n483 B.n482 585
R279 B.n484 B.n483 585
R280 B.n213 B.n212 585
R281 B.n214 B.n213 585
R282 B.n493 B.n492 585
R283 B.n492 B.n491 585
R284 B.n494 B.n211 585
R285 B.n211 B.n210 585
R286 B.n496 B.n495 585
R287 B.n497 B.n496 585
R288 B.n2 B.n0 585
R289 B.n4 B.n2 585
R290 B.n3 B.n1 585
R291 B.n594 B.n3 585
R292 B.n592 B.n591 585
R293 B.n593 B.n592 585
R294 B.n590 B.n9 585
R295 B.n9 B.n8 585
R296 B.n589 B.n588 585
R297 B.n588 B.n587 585
R298 B.n11 B.n10 585
R299 B.n586 B.n11 585
R300 B.n584 B.n583 585
R301 B.n585 B.n584 585
R302 B.n582 B.n16 585
R303 B.n16 B.n15 585
R304 B.n581 B.n580 585
R305 B.n580 B.n579 585
R306 B.n18 B.n17 585
R307 B.n578 B.n18 585
R308 B.n576 B.n575 585
R309 B.n577 B.n576 585
R310 B.n574 B.n23 585
R311 B.n23 B.n22 585
R312 B.n573 B.n572 585
R313 B.n572 B.n571 585
R314 B.n25 B.n24 585
R315 B.n570 B.n25 585
R316 B.n568 B.n567 585
R317 B.n569 B.n568 585
R318 B.n566 B.n30 585
R319 B.n30 B.n29 585
R320 B.n565 B.n564 585
R321 B.n564 B.n563 585
R322 B.n32 B.n31 585
R323 B.n562 B.n32 585
R324 B.n560 B.n559 585
R325 B.n561 B.n560 585
R326 B.n558 B.n37 585
R327 B.n37 B.n36 585
R328 B.n557 B.n556 585
R329 B.n556 B.n555 585
R330 B.n39 B.n38 585
R331 B.n554 B.n39 585
R332 B.n552 B.n551 585
R333 B.n553 B.n552 585
R334 B.n550 B.n44 585
R335 B.n44 B.n43 585
R336 B.n549 B.n548 585
R337 B.n548 B.n547 585
R338 B.n46 B.n45 585
R339 B.n546 B.n46 585
R340 B.n544 B.n543 585
R341 B.n545 B.n544 585
R342 B.n542 B.n51 585
R343 B.n51 B.n50 585
R344 B.n597 B.n596 585
R345 B.n596 B.n595 585
R346 B.n419 B.n259 526.135
R347 B.n540 B.n51 526.135
R348 B.n291 B.n257 526.135
R349 B.n536 B.n84 526.135
R350 B.n295 B.t14 332.546
R351 B.n293 B.t6 332.546
R352 B.n88 B.t10 332.546
R353 B.n85 B.t17 332.546
R354 B.n538 B.n537 256.663
R355 B.n538 B.n82 256.663
R356 B.n538 B.n81 256.663
R357 B.n538 B.n80 256.663
R358 B.n538 B.n79 256.663
R359 B.n538 B.n78 256.663
R360 B.n538 B.n77 256.663
R361 B.n538 B.n76 256.663
R362 B.n538 B.n75 256.663
R363 B.n538 B.n74 256.663
R364 B.n538 B.n73 256.663
R365 B.n538 B.n72 256.663
R366 B.n538 B.n71 256.663
R367 B.n538 B.n70 256.663
R368 B.n538 B.n69 256.663
R369 B.n538 B.n68 256.663
R370 B.n538 B.n67 256.663
R371 B.n538 B.n66 256.663
R372 B.n538 B.n65 256.663
R373 B.n538 B.n64 256.663
R374 B.n538 B.n63 256.663
R375 B.n538 B.n62 256.663
R376 B.n538 B.n61 256.663
R377 B.n538 B.n60 256.663
R378 B.n538 B.n59 256.663
R379 B.n538 B.n58 256.663
R380 B.n538 B.n57 256.663
R381 B.n538 B.n56 256.663
R382 B.n538 B.n55 256.663
R383 B.n538 B.n54 256.663
R384 B.n539 B.n538 256.663
R385 B.n418 B.n417 256.663
R386 B.n417 B.n262 256.663
R387 B.n417 B.n263 256.663
R388 B.n417 B.n264 256.663
R389 B.n417 B.n265 256.663
R390 B.n417 B.n266 256.663
R391 B.n417 B.n267 256.663
R392 B.n417 B.n268 256.663
R393 B.n417 B.n269 256.663
R394 B.n417 B.n270 256.663
R395 B.n417 B.n271 256.663
R396 B.n417 B.n272 256.663
R397 B.n417 B.n273 256.663
R398 B.n417 B.n274 256.663
R399 B.n417 B.n275 256.663
R400 B.n417 B.n276 256.663
R401 B.n417 B.n277 256.663
R402 B.n417 B.n278 256.663
R403 B.n417 B.n279 256.663
R404 B.n417 B.n280 256.663
R405 B.n417 B.n281 256.663
R406 B.n417 B.n282 256.663
R407 B.n417 B.n283 256.663
R408 B.n417 B.n284 256.663
R409 B.n417 B.n285 256.663
R410 B.n417 B.n286 256.663
R411 B.n417 B.n287 256.663
R412 B.n417 B.n288 256.663
R413 B.n417 B.n289 256.663
R414 B.n417 B.n290 256.663
R415 B.n295 B.t16 224.216
R416 B.n85 B.t18 224.216
R417 B.n293 B.t9 224.216
R418 B.n88 B.t12 224.216
R419 B.n296 B.t15 192.993
R420 B.n86 B.t19 192.993
R421 B.n294 B.t8 192.993
R422 B.n89 B.t13 192.993
R423 B.n423 B.n259 163.367
R424 B.n423 B.n253 163.367
R425 B.n431 B.n253 163.367
R426 B.n431 B.n251 163.367
R427 B.n435 B.n251 163.367
R428 B.n435 B.n245 163.367
R429 B.n443 B.n245 163.367
R430 B.n443 B.n243 163.367
R431 B.n447 B.n243 163.367
R432 B.n447 B.n237 163.367
R433 B.n455 B.n237 163.367
R434 B.n455 B.n235 163.367
R435 B.n459 B.n235 163.367
R436 B.n459 B.n229 163.367
R437 B.n467 B.n229 163.367
R438 B.n467 B.n227 163.367
R439 B.n471 B.n227 163.367
R440 B.n471 B.n221 163.367
R441 B.n479 B.n221 163.367
R442 B.n479 B.n219 163.367
R443 B.n483 B.n219 163.367
R444 B.n483 B.n213 163.367
R445 B.n492 B.n213 163.367
R446 B.n492 B.n211 163.367
R447 B.n496 B.n211 163.367
R448 B.n496 B.n2 163.367
R449 B.n596 B.n2 163.367
R450 B.n596 B.n3 163.367
R451 B.n592 B.n3 163.367
R452 B.n592 B.n9 163.367
R453 B.n588 B.n9 163.367
R454 B.n588 B.n11 163.367
R455 B.n584 B.n11 163.367
R456 B.n584 B.n16 163.367
R457 B.n580 B.n16 163.367
R458 B.n580 B.n18 163.367
R459 B.n576 B.n18 163.367
R460 B.n576 B.n23 163.367
R461 B.n572 B.n23 163.367
R462 B.n572 B.n25 163.367
R463 B.n568 B.n25 163.367
R464 B.n568 B.n30 163.367
R465 B.n564 B.n30 163.367
R466 B.n564 B.n32 163.367
R467 B.n560 B.n32 163.367
R468 B.n560 B.n37 163.367
R469 B.n556 B.n37 163.367
R470 B.n556 B.n39 163.367
R471 B.n552 B.n39 163.367
R472 B.n552 B.n44 163.367
R473 B.n548 B.n44 163.367
R474 B.n548 B.n46 163.367
R475 B.n544 B.n46 163.367
R476 B.n544 B.n51 163.367
R477 B.n416 B.n261 163.367
R478 B.n416 B.n292 163.367
R479 B.n412 B.n411 163.367
R480 B.n408 B.n407 163.367
R481 B.n404 B.n403 163.367
R482 B.n400 B.n399 163.367
R483 B.n396 B.n395 163.367
R484 B.n392 B.n391 163.367
R485 B.n388 B.n387 163.367
R486 B.n384 B.n383 163.367
R487 B.n380 B.n379 163.367
R488 B.n376 B.n375 163.367
R489 B.n372 B.n371 163.367
R490 B.n367 B.n366 163.367
R491 B.n363 B.n362 163.367
R492 B.n359 B.n358 163.367
R493 B.n355 B.n354 163.367
R494 B.n351 B.n350 163.367
R495 B.n346 B.n345 163.367
R496 B.n342 B.n341 163.367
R497 B.n338 B.n337 163.367
R498 B.n334 B.n333 163.367
R499 B.n330 B.n329 163.367
R500 B.n326 B.n325 163.367
R501 B.n322 B.n321 163.367
R502 B.n318 B.n317 163.367
R503 B.n314 B.n313 163.367
R504 B.n310 B.n309 163.367
R505 B.n306 B.n305 163.367
R506 B.n302 B.n301 163.367
R507 B.n298 B.n291 163.367
R508 B.n425 B.n257 163.367
R509 B.n425 B.n255 163.367
R510 B.n429 B.n255 163.367
R511 B.n429 B.n249 163.367
R512 B.n437 B.n249 163.367
R513 B.n437 B.n247 163.367
R514 B.n441 B.n247 163.367
R515 B.n441 B.n241 163.367
R516 B.n449 B.n241 163.367
R517 B.n449 B.n239 163.367
R518 B.n453 B.n239 163.367
R519 B.n453 B.n233 163.367
R520 B.n461 B.n233 163.367
R521 B.n461 B.n231 163.367
R522 B.n465 B.n231 163.367
R523 B.n465 B.n224 163.367
R524 B.n473 B.n224 163.367
R525 B.n473 B.n222 163.367
R526 B.n477 B.n222 163.367
R527 B.n477 B.n217 163.367
R528 B.n485 B.n217 163.367
R529 B.n485 B.n215 163.367
R530 B.n490 B.n215 163.367
R531 B.n490 B.n209 163.367
R532 B.n498 B.n209 163.367
R533 B.n499 B.n498 163.367
R534 B.n499 B.n5 163.367
R535 B.n6 B.n5 163.367
R536 B.n7 B.n6 163.367
R537 B.n504 B.n7 163.367
R538 B.n504 B.n12 163.367
R539 B.n13 B.n12 163.367
R540 B.n14 B.n13 163.367
R541 B.n509 B.n14 163.367
R542 B.n509 B.n19 163.367
R543 B.n20 B.n19 163.367
R544 B.n21 B.n20 163.367
R545 B.n514 B.n21 163.367
R546 B.n514 B.n26 163.367
R547 B.n27 B.n26 163.367
R548 B.n28 B.n27 163.367
R549 B.n519 B.n28 163.367
R550 B.n519 B.n33 163.367
R551 B.n34 B.n33 163.367
R552 B.n35 B.n34 163.367
R553 B.n524 B.n35 163.367
R554 B.n524 B.n40 163.367
R555 B.n41 B.n40 163.367
R556 B.n42 B.n41 163.367
R557 B.n529 B.n42 163.367
R558 B.n529 B.n47 163.367
R559 B.n48 B.n47 163.367
R560 B.n49 B.n48 163.367
R561 B.n84 B.n49 163.367
R562 B.n91 B.n53 163.367
R563 B.n95 B.n94 163.367
R564 B.n99 B.n98 163.367
R565 B.n103 B.n102 163.367
R566 B.n107 B.n106 163.367
R567 B.n111 B.n110 163.367
R568 B.n115 B.n114 163.367
R569 B.n119 B.n118 163.367
R570 B.n123 B.n122 163.367
R571 B.n127 B.n126 163.367
R572 B.n131 B.n130 163.367
R573 B.n135 B.n134 163.367
R574 B.n139 B.n138 163.367
R575 B.n143 B.n142 163.367
R576 B.n147 B.n146 163.367
R577 B.n151 B.n150 163.367
R578 B.n155 B.n154 163.367
R579 B.n159 B.n158 163.367
R580 B.n163 B.n162 163.367
R581 B.n167 B.n166 163.367
R582 B.n171 B.n170 163.367
R583 B.n175 B.n174 163.367
R584 B.n179 B.n178 163.367
R585 B.n183 B.n182 163.367
R586 B.n187 B.n186 163.367
R587 B.n191 B.n190 163.367
R588 B.n195 B.n194 163.367
R589 B.n199 B.n198 163.367
R590 B.n203 B.n202 163.367
R591 B.n205 B.n83 163.367
R592 B.n417 B.n258 115.695
R593 B.n538 B.n50 115.695
R594 B.n419 B.n418 71.676
R595 B.n292 B.n262 71.676
R596 B.n411 B.n263 71.676
R597 B.n407 B.n264 71.676
R598 B.n403 B.n265 71.676
R599 B.n399 B.n266 71.676
R600 B.n395 B.n267 71.676
R601 B.n391 B.n268 71.676
R602 B.n387 B.n269 71.676
R603 B.n383 B.n270 71.676
R604 B.n379 B.n271 71.676
R605 B.n375 B.n272 71.676
R606 B.n371 B.n273 71.676
R607 B.n366 B.n274 71.676
R608 B.n362 B.n275 71.676
R609 B.n358 B.n276 71.676
R610 B.n354 B.n277 71.676
R611 B.n350 B.n278 71.676
R612 B.n345 B.n279 71.676
R613 B.n341 B.n280 71.676
R614 B.n337 B.n281 71.676
R615 B.n333 B.n282 71.676
R616 B.n329 B.n283 71.676
R617 B.n325 B.n284 71.676
R618 B.n321 B.n285 71.676
R619 B.n317 B.n286 71.676
R620 B.n313 B.n287 71.676
R621 B.n309 B.n288 71.676
R622 B.n305 B.n289 71.676
R623 B.n301 B.n290 71.676
R624 B.n540 B.n539 71.676
R625 B.n91 B.n54 71.676
R626 B.n95 B.n55 71.676
R627 B.n99 B.n56 71.676
R628 B.n103 B.n57 71.676
R629 B.n107 B.n58 71.676
R630 B.n111 B.n59 71.676
R631 B.n115 B.n60 71.676
R632 B.n119 B.n61 71.676
R633 B.n123 B.n62 71.676
R634 B.n127 B.n63 71.676
R635 B.n131 B.n64 71.676
R636 B.n135 B.n65 71.676
R637 B.n139 B.n66 71.676
R638 B.n143 B.n67 71.676
R639 B.n147 B.n68 71.676
R640 B.n151 B.n69 71.676
R641 B.n155 B.n70 71.676
R642 B.n159 B.n71 71.676
R643 B.n163 B.n72 71.676
R644 B.n167 B.n73 71.676
R645 B.n171 B.n74 71.676
R646 B.n175 B.n75 71.676
R647 B.n179 B.n76 71.676
R648 B.n183 B.n77 71.676
R649 B.n187 B.n78 71.676
R650 B.n191 B.n79 71.676
R651 B.n195 B.n80 71.676
R652 B.n199 B.n81 71.676
R653 B.n203 B.n82 71.676
R654 B.n537 B.n83 71.676
R655 B.n537 B.n536 71.676
R656 B.n205 B.n82 71.676
R657 B.n202 B.n81 71.676
R658 B.n198 B.n80 71.676
R659 B.n194 B.n79 71.676
R660 B.n190 B.n78 71.676
R661 B.n186 B.n77 71.676
R662 B.n182 B.n76 71.676
R663 B.n178 B.n75 71.676
R664 B.n174 B.n74 71.676
R665 B.n170 B.n73 71.676
R666 B.n166 B.n72 71.676
R667 B.n162 B.n71 71.676
R668 B.n158 B.n70 71.676
R669 B.n154 B.n69 71.676
R670 B.n150 B.n68 71.676
R671 B.n146 B.n67 71.676
R672 B.n142 B.n66 71.676
R673 B.n138 B.n65 71.676
R674 B.n134 B.n64 71.676
R675 B.n130 B.n63 71.676
R676 B.n126 B.n62 71.676
R677 B.n122 B.n61 71.676
R678 B.n118 B.n60 71.676
R679 B.n114 B.n59 71.676
R680 B.n110 B.n58 71.676
R681 B.n106 B.n57 71.676
R682 B.n102 B.n56 71.676
R683 B.n98 B.n55 71.676
R684 B.n94 B.n54 71.676
R685 B.n539 B.n53 71.676
R686 B.n418 B.n261 71.676
R687 B.n412 B.n262 71.676
R688 B.n408 B.n263 71.676
R689 B.n404 B.n264 71.676
R690 B.n400 B.n265 71.676
R691 B.n396 B.n266 71.676
R692 B.n392 B.n267 71.676
R693 B.n388 B.n268 71.676
R694 B.n384 B.n269 71.676
R695 B.n380 B.n270 71.676
R696 B.n376 B.n271 71.676
R697 B.n372 B.n272 71.676
R698 B.n367 B.n273 71.676
R699 B.n363 B.n274 71.676
R700 B.n359 B.n275 71.676
R701 B.n355 B.n276 71.676
R702 B.n351 B.n277 71.676
R703 B.n346 B.n278 71.676
R704 B.n342 B.n279 71.676
R705 B.n338 B.n280 71.676
R706 B.n334 B.n281 71.676
R707 B.n330 B.n282 71.676
R708 B.n326 B.n283 71.676
R709 B.n322 B.n284 71.676
R710 B.n318 B.n285 71.676
R711 B.n314 B.n286 71.676
R712 B.n310 B.n287 71.676
R713 B.n306 B.n288 71.676
R714 B.n302 B.n289 71.676
R715 B.n298 B.n290 71.676
R716 B.n424 B.n258 61.9467
R717 B.n424 B.n254 61.9467
R718 B.n430 B.n254 61.9467
R719 B.n430 B.n250 61.9467
R720 B.n436 B.n250 61.9467
R721 B.n442 B.n246 61.9467
R722 B.n442 B.n242 61.9467
R723 B.n448 B.n242 61.9467
R724 B.n448 B.n238 61.9467
R725 B.n454 B.n238 61.9467
R726 B.n454 B.n234 61.9467
R727 B.n460 B.n234 61.9467
R728 B.n466 B.n230 61.9467
R729 B.n466 B.n225 61.9467
R730 B.n472 B.n225 61.9467
R731 B.n472 B.n226 61.9467
R732 B.n478 B.n218 61.9467
R733 B.n484 B.n218 61.9467
R734 B.n484 B.n214 61.9467
R735 B.n491 B.n214 61.9467
R736 B.n497 B.n210 61.9467
R737 B.n497 B.n4 61.9467
R738 B.n595 B.n4 61.9467
R739 B.n595 B.n594 61.9467
R740 B.n594 B.n593 61.9467
R741 B.n593 B.n8 61.9467
R742 B.n587 B.n586 61.9467
R743 B.n586 B.n585 61.9467
R744 B.n585 B.n15 61.9467
R745 B.n579 B.n15 61.9467
R746 B.n578 B.n577 61.9467
R747 B.n577 B.n22 61.9467
R748 B.n571 B.n22 61.9467
R749 B.n571 B.n570 61.9467
R750 B.n569 B.n29 61.9467
R751 B.n563 B.n29 61.9467
R752 B.n563 B.n562 61.9467
R753 B.n562 B.n561 61.9467
R754 B.n561 B.n36 61.9467
R755 B.n555 B.n36 61.9467
R756 B.n555 B.n554 61.9467
R757 B.n553 B.n43 61.9467
R758 B.n547 B.n43 61.9467
R759 B.n547 B.n546 61.9467
R760 B.n546 B.n545 61.9467
R761 B.n545 B.n50 61.9467
R762 B.t1 B.n210 60.1247
R763 B.t0 B.n8 60.1247
R764 B.n348 B.n296 59.5399
R765 B.n369 B.n294 59.5399
R766 B.n90 B.n89 59.5399
R767 B.n87 B.n86 59.5399
R768 B.n478 B.t3 43.7272
R769 B.n579 B.t2 43.7272
R770 B.n436 B.t7 38.2614
R771 B.t11 B.n553 38.2614
R772 B.n460 B.t5 34.6175
R773 B.t4 B.n569 34.6175
R774 B.n542 B.n541 34.1859
R775 B.n535 B.n534 34.1859
R776 B.n297 B.n256 34.1859
R777 B.n421 B.n420 34.1859
R778 B.n296 B.n295 31.2247
R779 B.n294 B.n293 31.2247
R780 B.n89 B.n88 31.2247
R781 B.n86 B.n85 31.2247
R782 B.t5 B.n230 27.3297
R783 B.n570 B.t4 27.3297
R784 B.t7 B.n246 23.6858
R785 B.n554 B.t11 23.6858
R786 B.n226 B.t3 18.22
R787 B.t2 B.n578 18.22
R788 B B.n597 18.0485
R789 B.n541 B.n52 10.6151
R790 B.n92 B.n52 10.6151
R791 B.n93 B.n92 10.6151
R792 B.n96 B.n93 10.6151
R793 B.n97 B.n96 10.6151
R794 B.n100 B.n97 10.6151
R795 B.n101 B.n100 10.6151
R796 B.n104 B.n101 10.6151
R797 B.n105 B.n104 10.6151
R798 B.n108 B.n105 10.6151
R799 B.n109 B.n108 10.6151
R800 B.n112 B.n109 10.6151
R801 B.n113 B.n112 10.6151
R802 B.n116 B.n113 10.6151
R803 B.n117 B.n116 10.6151
R804 B.n120 B.n117 10.6151
R805 B.n121 B.n120 10.6151
R806 B.n124 B.n121 10.6151
R807 B.n125 B.n124 10.6151
R808 B.n128 B.n125 10.6151
R809 B.n129 B.n128 10.6151
R810 B.n132 B.n129 10.6151
R811 B.n133 B.n132 10.6151
R812 B.n136 B.n133 10.6151
R813 B.n137 B.n136 10.6151
R814 B.n141 B.n140 10.6151
R815 B.n144 B.n141 10.6151
R816 B.n145 B.n144 10.6151
R817 B.n148 B.n145 10.6151
R818 B.n149 B.n148 10.6151
R819 B.n152 B.n149 10.6151
R820 B.n153 B.n152 10.6151
R821 B.n156 B.n153 10.6151
R822 B.n157 B.n156 10.6151
R823 B.n161 B.n160 10.6151
R824 B.n164 B.n161 10.6151
R825 B.n165 B.n164 10.6151
R826 B.n168 B.n165 10.6151
R827 B.n169 B.n168 10.6151
R828 B.n172 B.n169 10.6151
R829 B.n173 B.n172 10.6151
R830 B.n176 B.n173 10.6151
R831 B.n177 B.n176 10.6151
R832 B.n180 B.n177 10.6151
R833 B.n181 B.n180 10.6151
R834 B.n184 B.n181 10.6151
R835 B.n185 B.n184 10.6151
R836 B.n188 B.n185 10.6151
R837 B.n189 B.n188 10.6151
R838 B.n192 B.n189 10.6151
R839 B.n193 B.n192 10.6151
R840 B.n196 B.n193 10.6151
R841 B.n197 B.n196 10.6151
R842 B.n200 B.n197 10.6151
R843 B.n201 B.n200 10.6151
R844 B.n204 B.n201 10.6151
R845 B.n206 B.n204 10.6151
R846 B.n207 B.n206 10.6151
R847 B.n535 B.n207 10.6151
R848 B.n426 B.n256 10.6151
R849 B.n427 B.n426 10.6151
R850 B.n428 B.n427 10.6151
R851 B.n428 B.n248 10.6151
R852 B.n438 B.n248 10.6151
R853 B.n439 B.n438 10.6151
R854 B.n440 B.n439 10.6151
R855 B.n440 B.n240 10.6151
R856 B.n450 B.n240 10.6151
R857 B.n451 B.n450 10.6151
R858 B.n452 B.n451 10.6151
R859 B.n452 B.n232 10.6151
R860 B.n462 B.n232 10.6151
R861 B.n463 B.n462 10.6151
R862 B.n464 B.n463 10.6151
R863 B.n464 B.n223 10.6151
R864 B.n474 B.n223 10.6151
R865 B.n475 B.n474 10.6151
R866 B.n476 B.n475 10.6151
R867 B.n476 B.n216 10.6151
R868 B.n486 B.n216 10.6151
R869 B.n487 B.n486 10.6151
R870 B.n489 B.n487 10.6151
R871 B.n489 B.n488 10.6151
R872 B.n488 B.n208 10.6151
R873 B.n500 B.n208 10.6151
R874 B.n501 B.n500 10.6151
R875 B.n502 B.n501 10.6151
R876 B.n503 B.n502 10.6151
R877 B.n505 B.n503 10.6151
R878 B.n506 B.n505 10.6151
R879 B.n507 B.n506 10.6151
R880 B.n508 B.n507 10.6151
R881 B.n510 B.n508 10.6151
R882 B.n511 B.n510 10.6151
R883 B.n512 B.n511 10.6151
R884 B.n513 B.n512 10.6151
R885 B.n515 B.n513 10.6151
R886 B.n516 B.n515 10.6151
R887 B.n517 B.n516 10.6151
R888 B.n518 B.n517 10.6151
R889 B.n520 B.n518 10.6151
R890 B.n521 B.n520 10.6151
R891 B.n522 B.n521 10.6151
R892 B.n523 B.n522 10.6151
R893 B.n525 B.n523 10.6151
R894 B.n526 B.n525 10.6151
R895 B.n527 B.n526 10.6151
R896 B.n528 B.n527 10.6151
R897 B.n530 B.n528 10.6151
R898 B.n531 B.n530 10.6151
R899 B.n532 B.n531 10.6151
R900 B.n533 B.n532 10.6151
R901 B.n534 B.n533 10.6151
R902 B.n420 B.n260 10.6151
R903 B.n415 B.n260 10.6151
R904 B.n415 B.n414 10.6151
R905 B.n414 B.n413 10.6151
R906 B.n413 B.n410 10.6151
R907 B.n410 B.n409 10.6151
R908 B.n409 B.n406 10.6151
R909 B.n406 B.n405 10.6151
R910 B.n405 B.n402 10.6151
R911 B.n402 B.n401 10.6151
R912 B.n401 B.n398 10.6151
R913 B.n398 B.n397 10.6151
R914 B.n397 B.n394 10.6151
R915 B.n394 B.n393 10.6151
R916 B.n393 B.n390 10.6151
R917 B.n390 B.n389 10.6151
R918 B.n389 B.n386 10.6151
R919 B.n386 B.n385 10.6151
R920 B.n385 B.n382 10.6151
R921 B.n382 B.n381 10.6151
R922 B.n381 B.n378 10.6151
R923 B.n378 B.n377 10.6151
R924 B.n377 B.n374 10.6151
R925 B.n374 B.n373 10.6151
R926 B.n373 B.n370 10.6151
R927 B.n368 B.n365 10.6151
R928 B.n365 B.n364 10.6151
R929 B.n364 B.n361 10.6151
R930 B.n361 B.n360 10.6151
R931 B.n360 B.n357 10.6151
R932 B.n357 B.n356 10.6151
R933 B.n356 B.n353 10.6151
R934 B.n353 B.n352 10.6151
R935 B.n352 B.n349 10.6151
R936 B.n347 B.n344 10.6151
R937 B.n344 B.n343 10.6151
R938 B.n343 B.n340 10.6151
R939 B.n340 B.n339 10.6151
R940 B.n339 B.n336 10.6151
R941 B.n336 B.n335 10.6151
R942 B.n335 B.n332 10.6151
R943 B.n332 B.n331 10.6151
R944 B.n331 B.n328 10.6151
R945 B.n328 B.n327 10.6151
R946 B.n327 B.n324 10.6151
R947 B.n324 B.n323 10.6151
R948 B.n323 B.n320 10.6151
R949 B.n320 B.n319 10.6151
R950 B.n319 B.n316 10.6151
R951 B.n316 B.n315 10.6151
R952 B.n315 B.n312 10.6151
R953 B.n312 B.n311 10.6151
R954 B.n311 B.n308 10.6151
R955 B.n308 B.n307 10.6151
R956 B.n307 B.n304 10.6151
R957 B.n304 B.n303 10.6151
R958 B.n303 B.n300 10.6151
R959 B.n300 B.n299 10.6151
R960 B.n299 B.n297 10.6151
R961 B.n422 B.n421 10.6151
R962 B.n422 B.n252 10.6151
R963 B.n432 B.n252 10.6151
R964 B.n433 B.n432 10.6151
R965 B.n434 B.n433 10.6151
R966 B.n434 B.n244 10.6151
R967 B.n444 B.n244 10.6151
R968 B.n445 B.n444 10.6151
R969 B.n446 B.n445 10.6151
R970 B.n446 B.n236 10.6151
R971 B.n456 B.n236 10.6151
R972 B.n457 B.n456 10.6151
R973 B.n458 B.n457 10.6151
R974 B.n458 B.n228 10.6151
R975 B.n468 B.n228 10.6151
R976 B.n469 B.n468 10.6151
R977 B.n470 B.n469 10.6151
R978 B.n470 B.n220 10.6151
R979 B.n480 B.n220 10.6151
R980 B.n481 B.n480 10.6151
R981 B.n482 B.n481 10.6151
R982 B.n482 B.n212 10.6151
R983 B.n493 B.n212 10.6151
R984 B.n494 B.n493 10.6151
R985 B.n495 B.n494 10.6151
R986 B.n495 B.n0 10.6151
R987 B.n591 B.n1 10.6151
R988 B.n591 B.n590 10.6151
R989 B.n590 B.n589 10.6151
R990 B.n589 B.n10 10.6151
R991 B.n583 B.n10 10.6151
R992 B.n583 B.n582 10.6151
R993 B.n582 B.n581 10.6151
R994 B.n581 B.n17 10.6151
R995 B.n575 B.n17 10.6151
R996 B.n575 B.n574 10.6151
R997 B.n574 B.n573 10.6151
R998 B.n573 B.n24 10.6151
R999 B.n567 B.n24 10.6151
R1000 B.n567 B.n566 10.6151
R1001 B.n566 B.n565 10.6151
R1002 B.n565 B.n31 10.6151
R1003 B.n559 B.n31 10.6151
R1004 B.n559 B.n558 10.6151
R1005 B.n558 B.n557 10.6151
R1006 B.n557 B.n38 10.6151
R1007 B.n551 B.n38 10.6151
R1008 B.n551 B.n550 10.6151
R1009 B.n550 B.n549 10.6151
R1010 B.n549 B.n45 10.6151
R1011 B.n543 B.n45 10.6151
R1012 B.n543 B.n542 10.6151
R1013 B.n137 B.n90 9.36635
R1014 B.n160 B.n87 9.36635
R1015 B.n370 B.n369 9.36635
R1016 B.n348 B.n347 9.36635
R1017 B.n597 B.n0 2.81026
R1018 B.n597 B.n1 2.81026
R1019 B.n491 B.t1 1.82245
R1020 B.n587 B.t0 1.82245
R1021 B.n140 B.n90 1.24928
R1022 B.n157 B.n87 1.24928
R1023 B.n369 B.n368 1.24928
R1024 B.n349 B.n348 1.24928
R1025 VP.n5 VP.t2 178.02
R1026 VP.n7 VP.n6 161.3
R1027 VP.n8 VP.n3 161.3
R1028 VP.n18 VP.n0 161.3
R1029 VP.n17 VP.n16 161.3
R1030 VP.n15 VP.n14 161.3
R1031 VP.n13 VP.n2 161.3
R1032 VP.n12 VP.t1 158.721
R1033 VP.n19 VP.t0 158.721
R1034 VP.n9 VP.t3 158.721
R1035 VP.n1 VP.t4 128.031
R1036 VP.n4 VP.t5 128.031
R1037 VP.n10 VP.n9 80.6037
R1038 VP.n20 VP.n19 80.6037
R1039 VP.n12 VP.n11 80.6037
R1040 VP.n5 VP.n4 45.4787
R1041 VP.n11 VP.n10 39.74
R1042 VP.n14 VP.n13 35.2488
R1043 VP.n18 VP.n17 35.2488
R1044 VP.n8 VP.n7 35.2488
R1045 VP.n13 VP.n12 32.1338
R1046 VP.n19 VP.n18 32.1338
R1047 VP.n9 VP.n8 32.1338
R1048 VP.n6 VP.n5 29.4552
R1049 VP.n14 VP.n1 12.2964
R1050 VP.n17 VP.n1 12.2964
R1051 VP.n7 VP.n4 12.2964
R1052 VP.n10 VP.n3 0.285035
R1053 VP.n11 VP.n2 0.285035
R1054 VP.n20 VP.n0 0.285035
R1055 VP.n6 VP.n3 0.189894
R1056 VP.n15 VP.n2 0.189894
R1057 VP.n16 VP.n15 0.189894
R1058 VP.n16 VP.n0 0.189894
R1059 VP VP.n20 0.146778
R1060 VTAIL.n146 VTAIL.n116 289.615
R1061 VTAIL.n32 VTAIL.n2 289.615
R1062 VTAIL.n110 VTAIL.n80 289.615
R1063 VTAIL.n72 VTAIL.n42 289.615
R1064 VTAIL.n129 VTAIL.n128 185
R1065 VTAIL.n131 VTAIL.n130 185
R1066 VTAIL.n124 VTAIL.n123 185
R1067 VTAIL.n137 VTAIL.n136 185
R1068 VTAIL.n139 VTAIL.n138 185
R1069 VTAIL.n120 VTAIL.n119 185
R1070 VTAIL.n145 VTAIL.n144 185
R1071 VTAIL.n147 VTAIL.n146 185
R1072 VTAIL.n15 VTAIL.n14 185
R1073 VTAIL.n17 VTAIL.n16 185
R1074 VTAIL.n10 VTAIL.n9 185
R1075 VTAIL.n23 VTAIL.n22 185
R1076 VTAIL.n25 VTAIL.n24 185
R1077 VTAIL.n6 VTAIL.n5 185
R1078 VTAIL.n31 VTAIL.n30 185
R1079 VTAIL.n33 VTAIL.n32 185
R1080 VTAIL.n111 VTAIL.n110 185
R1081 VTAIL.n109 VTAIL.n108 185
R1082 VTAIL.n84 VTAIL.n83 185
R1083 VTAIL.n103 VTAIL.n102 185
R1084 VTAIL.n101 VTAIL.n100 185
R1085 VTAIL.n88 VTAIL.n87 185
R1086 VTAIL.n95 VTAIL.n94 185
R1087 VTAIL.n93 VTAIL.n92 185
R1088 VTAIL.n73 VTAIL.n72 185
R1089 VTAIL.n71 VTAIL.n70 185
R1090 VTAIL.n46 VTAIL.n45 185
R1091 VTAIL.n65 VTAIL.n64 185
R1092 VTAIL.n63 VTAIL.n62 185
R1093 VTAIL.n50 VTAIL.n49 185
R1094 VTAIL.n57 VTAIL.n56 185
R1095 VTAIL.n55 VTAIL.n54 185
R1096 VTAIL.n127 VTAIL.t4 147.659
R1097 VTAIL.n13 VTAIL.t10 147.659
R1098 VTAIL.n91 VTAIL.t11 147.659
R1099 VTAIL.n53 VTAIL.t5 147.659
R1100 VTAIL.n130 VTAIL.n129 104.615
R1101 VTAIL.n130 VTAIL.n123 104.615
R1102 VTAIL.n137 VTAIL.n123 104.615
R1103 VTAIL.n138 VTAIL.n137 104.615
R1104 VTAIL.n138 VTAIL.n119 104.615
R1105 VTAIL.n145 VTAIL.n119 104.615
R1106 VTAIL.n146 VTAIL.n145 104.615
R1107 VTAIL.n16 VTAIL.n15 104.615
R1108 VTAIL.n16 VTAIL.n9 104.615
R1109 VTAIL.n23 VTAIL.n9 104.615
R1110 VTAIL.n24 VTAIL.n23 104.615
R1111 VTAIL.n24 VTAIL.n5 104.615
R1112 VTAIL.n31 VTAIL.n5 104.615
R1113 VTAIL.n32 VTAIL.n31 104.615
R1114 VTAIL.n110 VTAIL.n109 104.615
R1115 VTAIL.n109 VTAIL.n83 104.615
R1116 VTAIL.n102 VTAIL.n83 104.615
R1117 VTAIL.n102 VTAIL.n101 104.615
R1118 VTAIL.n101 VTAIL.n87 104.615
R1119 VTAIL.n94 VTAIL.n87 104.615
R1120 VTAIL.n94 VTAIL.n93 104.615
R1121 VTAIL.n72 VTAIL.n71 104.615
R1122 VTAIL.n71 VTAIL.n45 104.615
R1123 VTAIL.n64 VTAIL.n45 104.615
R1124 VTAIL.n64 VTAIL.n63 104.615
R1125 VTAIL.n63 VTAIL.n49 104.615
R1126 VTAIL.n56 VTAIL.n49 104.615
R1127 VTAIL.n56 VTAIL.n55 104.615
R1128 VTAIL.n129 VTAIL.t4 52.3082
R1129 VTAIL.n15 VTAIL.t10 52.3082
R1130 VTAIL.n93 VTAIL.t11 52.3082
R1131 VTAIL.n55 VTAIL.t5 52.3082
R1132 VTAIL.n79 VTAIL.n78 50.9468
R1133 VTAIL.n41 VTAIL.n40 50.9468
R1134 VTAIL.n1 VTAIL.n0 50.9467
R1135 VTAIL.n39 VTAIL.n38 50.9467
R1136 VTAIL.n151 VTAIL.n150 33.7369
R1137 VTAIL.n37 VTAIL.n36 33.7369
R1138 VTAIL.n115 VTAIL.n114 33.7369
R1139 VTAIL.n77 VTAIL.n76 33.7369
R1140 VTAIL.n41 VTAIL.n39 21.0048
R1141 VTAIL.n151 VTAIL.n115 19.6169
R1142 VTAIL.n128 VTAIL.n127 15.6676
R1143 VTAIL.n14 VTAIL.n13 15.6676
R1144 VTAIL.n92 VTAIL.n91 15.6676
R1145 VTAIL.n54 VTAIL.n53 15.6676
R1146 VTAIL.n131 VTAIL.n126 12.8005
R1147 VTAIL.n17 VTAIL.n12 12.8005
R1148 VTAIL.n95 VTAIL.n90 12.8005
R1149 VTAIL.n57 VTAIL.n52 12.8005
R1150 VTAIL.n132 VTAIL.n124 12.0247
R1151 VTAIL.n18 VTAIL.n10 12.0247
R1152 VTAIL.n96 VTAIL.n88 12.0247
R1153 VTAIL.n58 VTAIL.n50 12.0247
R1154 VTAIL.n136 VTAIL.n135 11.249
R1155 VTAIL.n22 VTAIL.n21 11.249
R1156 VTAIL.n100 VTAIL.n99 11.249
R1157 VTAIL.n62 VTAIL.n61 11.249
R1158 VTAIL.n139 VTAIL.n122 10.4732
R1159 VTAIL.n25 VTAIL.n8 10.4732
R1160 VTAIL.n103 VTAIL.n86 10.4732
R1161 VTAIL.n65 VTAIL.n48 10.4732
R1162 VTAIL.n140 VTAIL.n120 9.69747
R1163 VTAIL.n26 VTAIL.n6 9.69747
R1164 VTAIL.n104 VTAIL.n84 9.69747
R1165 VTAIL.n66 VTAIL.n46 9.69747
R1166 VTAIL.n150 VTAIL.n149 9.45567
R1167 VTAIL.n36 VTAIL.n35 9.45567
R1168 VTAIL.n114 VTAIL.n113 9.45567
R1169 VTAIL.n76 VTAIL.n75 9.45567
R1170 VTAIL.n118 VTAIL.n117 9.3005
R1171 VTAIL.n143 VTAIL.n142 9.3005
R1172 VTAIL.n141 VTAIL.n140 9.3005
R1173 VTAIL.n122 VTAIL.n121 9.3005
R1174 VTAIL.n135 VTAIL.n134 9.3005
R1175 VTAIL.n133 VTAIL.n132 9.3005
R1176 VTAIL.n126 VTAIL.n125 9.3005
R1177 VTAIL.n149 VTAIL.n148 9.3005
R1178 VTAIL.n4 VTAIL.n3 9.3005
R1179 VTAIL.n29 VTAIL.n28 9.3005
R1180 VTAIL.n27 VTAIL.n26 9.3005
R1181 VTAIL.n8 VTAIL.n7 9.3005
R1182 VTAIL.n21 VTAIL.n20 9.3005
R1183 VTAIL.n19 VTAIL.n18 9.3005
R1184 VTAIL.n12 VTAIL.n11 9.3005
R1185 VTAIL.n35 VTAIL.n34 9.3005
R1186 VTAIL.n113 VTAIL.n112 9.3005
R1187 VTAIL.n82 VTAIL.n81 9.3005
R1188 VTAIL.n107 VTAIL.n106 9.3005
R1189 VTAIL.n105 VTAIL.n104 9.3005
R1190 VTAIL.n86 VTAIL.n85 9.3005
R1191 VTAIL.n99 VTAIL.n98 9.3005
R1192 VTAIL.n97 VTAIL.n96 9.3005
R1193 VTAIL.n90 VTAIL.n89 9.3005
R1194 VTAIL.n75 VTAIL.n74 9.3005
R1195 VTAIL.n44 VTAIL.n43 9.3005
R1196 VTAIL.n69 VTAIL.n68 9.3005
R1197 VTAIL.n67 VTAIL.n66 9.3005
R1198 VTAIL.n48 VTAIL.n47 9.3005
R1199 VTAIL.n61 VTAIL.n60 9.3005
R1200 VTAIL.n59 VTAIL.n58 9.3005
R1201 VTAIL.n52 VTAIL.n51 9.3005
R1202 VTAIL.n144 VTAIL.n143 8.92171
R1203 VTAIL.n30 VTAIL.n29 8.92171
R1204 VTAIL.n108 VTAIL.n107 8.92171
R1205 VTAIL.n70 VTAIL.n69 8.92171
R1206 VTAIL.n147 VTAIL.n118 8.14595
R1207 VTAIL.n33 VTAIL.n4 8.14595
R1208 VTAIL.n111 VTAIL.n82 8.14595
R1209 VTAIL.n73 VTAIL.n44 8.14595
R1210 VTAIL.n148 VTAIL.n116 7.3702
R1211 VTAIL.n34 VTAIL.n2 7.3702
R1212 VTAIL.n112 VTAIL.n80 7.3702
R1213 VTAIL.n74 VTAIL.n42 7.3702
R1214 VTAIL.n150 VTAIL.n116 6.59444
R1215 VTAIL.n36 VTAIL.n2 6.59444
R1216 VTAIL.n114 VTAIL.n80 6.59444
R1217 VTAIL.n76 VTAIL.n42 6.59444
R1218 VTAIL.n148 VTAIL.n147 5.81868
R1219 VTAIL.n34 VTAIL.n33 5.81868
R1220 VTAIL.n112 VTAIL.n111 5.81868
R1221 VTAIL.n74 VTAIL.n73 5.81868
R1222 VTAIL.n144 VTAIL.n118 5.04292
R1223 VTAIL.n30 VTAIL.n4 5.04292
R1224 VTAIL.n108 VTAIL.n82 5.04292
R1225 VTAIL.n70 VTAIL.n44 5.04292
R1226 VTAIL.n127 VTAIL.n125 4.38571
R1227 VTAIL.n13 VTAIL.n11 4.38571
R1228 VTAIL.n91 VTAIL.n89 4.38571
R1229 VTAIL.n53 VTAIL.n51 4.38571
R1230 VTAIL.n143 VTAIL.n120 4.26717
R1231 VTAIL.n29 VTAIL.n6 4.26717
R1232 VTAIL.n107 VTAIL.n84 4.26717
R1233 VTAIL.n69 VTAIL.n46 4.26717
R1234 VTAIL.n140 VTAIL.n139 3.49141
R1235 VTAIL.n26 VTAIL.n25 3.49141
R1236 VTAIL.n104 VTAIL.n103 3.49141
R1237 VTAIL.n66 VTAIL.n65 3.49141
R1238 VTAIL.n0 VTAIL.t0 2.91226
R1239 VTAIL.n0 VTAIL.t1 2.91226
R1240 VTAIL.n38 VTAIL.t6 2.91226
R1241 VTAIL.n38 VTAIL.t8 2.91226
R1242 VTAIL.n78 VTAIL.t9 2.91226
R1243 VTAIL.n78 VTAIL.t7 2.91226
R1244 VTAIL.n40 VTAIL.t2 2.91226
R1245 VTAIL.n40 VTAIL.t3 2.91226
R1246 VTAIL.n136 VTAIL.n122 2.71565
R1247 VTAIL.n22 VTAIL.n8 2.71565
R1248 VTAIL.n100 VTAIL.n86 2.71565
R1249 VTAIL.n62 VTAIL.n48 2.71565
R1250 VTAIL.n135 VTAIL.n124 1.93989
R1251 VTAIL.n21 VTAIL.n10 1.93989
R1252 VTAIL.n99 VTAIL.n88 1.93989
R1253 VTAIL.n61 VTAIL.n50 1.93989
R1254 VTAIL.n77 VTAIL.n41 1.38843
R1255 VTAIL.n115 VTAIL.n79 1.38843
R1256 VTAIL.n39 VTAIL.n37 1.38843
R1257 VTAIL.n79 VTAIL.n77 1.16429
R1258 VTAIL.n37 VTAIL.n1 1.16429
R1259 VTAIL.n132 VTAIL.n131 1.16414
R1260 VTAIL.n18 VTAIL.n17 1.16414
R1261 VTAIL.n96 VTAIL.n95 1.16414
R1262 VTAIL.n58 VTAIL.n57 1.16414
R1263 VTAIL VTAIL.n151 0.983259
R1264 VTAIL VTAIL.n1 0.405672
R1265 VTAIL.n128 VTAIL.n126 0.388379
R1266 VTAIL.n14 VTAIL.n12 0.388379
R1267 VTAIL.n92 VTAIL.n90 0.388379
R1268 VTAIL.n54 VTAIL.n52 0.388379
R1269 VTAIL.n133 VTAIL.n125 0.155672
R1270 VTAIL.n134 VTAIL.n133 0.155672
R1271 VTAIL.n134 VTAIL.n121 0.155672
R1272 VTAIL.n141 VTAIL.n121 0.155672
R1273 VTAIL.n142 VTAIL.n141 0.155672
R1274 VTAIL.n142 VTAIL.n117 0.155672
R1275 VTAIL.n149 VTAIL.n117 0.155672
R1276 VTAIL.n19 VTAIL.n11 0.155672
R1277 VTAIL.n20 VTAIL.n19 0.155672
R1278 VTAIL.n20 VTAIL.n7 0.155672
R1279 VTAIL.n27 VTAIL.n7 0.155672
R1280 VTAIL.n28 VTAIL.n27 0.155672
R1281 VTAIL.n28 VTAIL.n3 0.155672
R1282 VTAIL.n35 VTAIL.n3 0.155672
R1283 VTAIL.n113 VTAIL.n81 0.155672
R1284 VTAIL.n106 VTAIL.n81 0.155672
R1285 VTAIL.n106 VTAIL.n105 0.155672
R1286 VTAIL.n105 VTAIL.n85 0.155672
R1287 VTAIL.n98 VTAIL.n85 0.155672
R1288 VTAIL.n98 VTAIL.n97 0.155672
R1289 VTAIL.n97 VTAIL.n89 0.155672
R1290 VTAIL.n75 VTAIL.n43 0.155672
R1291 VTAIL.n68 VTAIL.n43 0.155672
R1292 VTAIL.n68 VTAIL.n67 0.155672
R1293 VTAIL.n67 VTAIL.n47 0.155672
R1294 VTAIL.n60 VTAIL.n47 0.155672
R1295 VTAIL.n60 VTAIL.n59 0.155672
R1296 VTAIL.n59 VTAIL.n51 0.155672
R1297 VDD1.n30 VDD1.n0 289.615
R1298 VDD1.n65 VDD1.n35 289.615
R1299 VDD1.n31 VDD1.n30 185
R1300 VDD1.n29 VDD1.n28 185
R1301 VDD1.n4 VDD1.n3 185
R1302 VDD1.n23 VDD1.n22 185
R1303 VDD1.n21 VDD1.n20 185
R1304 VDD1.n8 VDD1.n7 185
R1305 VDD1.n15 VDD1.n14 185
R1306 VDD1.n13 VDD1.n12 185
R1307 VDD1.n48 VDD1.n47 185
R1308 VDD1.n50 VDD1.n49 185
R1309 VDD1.n43 VDD1.n42 185
R1310 VDD1.n56 VDD1.n55 185
R1311 VDD1.n58 VDD1.n57 185
R1312 VDD1.n39 VDD1.n38 185
R1313 VDD1.n64 VDD1.n63 185
R1314 VDD1.n66 VDD1.n65 185
R1315 VDD1.n11 VDD1.t3 147.659
R1316 VDD1.n46 VDD1.t4 147.659
R1317 VDD1.n30 VDD1.n29 104.615
R1318 VDD1.n29 VDD1.n3 104.615
R1319 VDD1.n22 VDD1.n3 104.615
R1320 VDD1.n22 VDD1.n21 104.615
R1321 VDD1.n21 VDD1.n7 104.615
R1322 VDD1.n14 VDD1.n7 104.615
R1323 VDD1.n14 VDD1.n13 104.615
R1324 VDD1.n49 VDD1.n48 104.615
R1325 VDD1.n49 VDD1.n42 104.615
R1326 VDD1.n56 VDD1.n42 104.615
R1327 VDD1.n57 VDD1.n56 104.615
R1328 VDD1.n57 VDD1.n38 104.615
R1329 VDD1.n64 VDD1.n38 104.615
R1330 VDD1.n65 VDD1.n64 104.615
R1331 VDD1.n71 VDD1.n70 67.9171
R1332 VDD1.n73 VDD1.n72 67.6255
R1333 VDD1.n13 VDD1.t3 52.3082
R1334 VDD1.n48 VDD1.t4 52.3082
R1335 VDD1 VDD1.n34 51.5148
R1336 VDD1.n71 VDD1.n69 51.4013
R1337 VDD1.n73 VDD1.n71 35.3651
R1338 VDD1.n12 VDD1.n11 15.6676
R1339 VDD1.n47 VDD1.n46 15.6676
R1340 VDD1.n15 VDD1.n10 12.8005
R1341 VDD1.n50 VDD1.n45 12.8005
R1342 VDD1.n16 VDD1.n8 12.0247
R1343 VDD1.n51 VDD1.n43 12.0247
R1344 VDD1.n20 VDD1.n19 11.249
R1345 VDD1.n55 VDD1.n54 11.249
R1346 VDD1.n23 VDD1.n6 10.4732
R1347 VDD1.n58 VDD1.n41 10.4732
R1348 VDD1.n24 VDD1.n4 9.69747
R1349 VDD1.n59 VDD1.n39 9.69747
R1350 VDD1.n34 VDD1.n33 9.45567
R1351 VDD1.n69 VDD1.n68 9.45567
R1352 VDD1.n33 VDD1.n32 9.3005
R1353 VDD1.n2 VDD1.n1 9.3005
R1354 VDD1.n27 VDD1.n26 9.3005
R1355 VDD1.n25 VDD1.n24 9.3005
R1356 VDD1.n6 VDD1.n5 9.3005
R1357 VDD1.n19 VDD1.n18 9.3005
R1358 VDD1.n17 VDD1.n16 9.3005
R1359 VDD1.n10 VDD1.n9 9.3005
R1360 VDD1.n37 VDD1.n36 9.3005
R1361 VDD1.n62 VDD1.n61 9.3005
R1362 VDD1.n60 VDD1.n59 9.3005
R1363 VDD1.n41 VDD1.n40 9.3005
R1364 VDD1.n54 VDD1.n53 9.3005
R1365 VDD1.n52 VDD1.n51 9.3005
R1366 VDD1.n45 VDD1.n44 9.3005
R1367 VDD1.n68 VDD1.n67 9.3005
R1368 VDD1.n28 VDD1.n27 8.92171
R1369 VDD1.n63 VDD1.n62 8.92171
R1370 VDD1.n31 VDD1.n2 8.14595
R1371 VDD1.n66 VDD1.n37 8.14595
R1372 VDD1.n32 VDD1.n0 7.3702
R1373 VDD1.n67 VDD1.n35 7.3702
R1374 VDD1.n34 VDD1.n0 6.59444
R1375 VDD1.n69 VDD1.n35 6.59444
R1376 VDD1.n32 VDD1.n31 5.81868
R1377 VDD1.n67 VDD1.n66 5.81868
R1378 VDD1.n28 VDD1.n2 5.04292
R1379 VDD1.n63 VDD1.n37 5.04292
R1380 VDD1.n11 VDD1.n9 4.38571
R1381 VDD1.n46 VDD1.n44 4.38571
R1382 VDD1.n27 VDD1.n4 4.26717
R1383 VDD1.n62 VDD1.n39 4.26717
R1384 VDD1.n24 VDD1.n23 3.49141
R1385 VDD1.n59 VDD1.n58 3.49141
R1386 VDD1.n72 VDD1.t0 2.91226
R1387 VDD1.n72 VDD1.t2 2.91226
R1388 VDD1.n70 VDD1.t1 2.91226
R1389 VDD1.n70 VDD1.t5 2.91226
R1390 VDD1.n20 VDD1.n6 2.71565
R1391 VDD1.n55 VDD1.n41 2.71565
R1392 VDD1.n19 VDD1.n8 1.93989
R1393 VDD1.n54 VDD1.n43 1.93989
R1394 VDD1.n16 VDD1.n15 1.16414
R1395 VDD1.n51 VDD1.n50 1.16414
R1396 VDD1.n12 VDD1.n10 0.388379
R1397 VDD1.n47 VDD1.n45 0.388379
R1398 VDD1 VDD1.n73 0.289293
R1399 VDD1.n33 VDD1.n1 0.155672
R1400 VDD1.n26 VDD1.n1 0.155672
R1401 VDD1.n26 VDD1.n25 0.155672
R1402 VDD1.n25 VDD1.n5 0.155672
R1403 VDD1.n18 VDD1.n5 0.155672
R1404 VDD1.n18 VDD1.n17 0.155672
R1405 VDD1.n17 VDD1.n9 0.155672
R1406 VDD1.n52 VDD1.n44 0.155672
R1407 VDD1.n53 VDD1.n52 0.155672
R1408 VDD1.n53 VDD1.n40 0.155672
R1409 VDD1.n60 VDD1.n40 0.155672
R1410 VDD1.n61 VDD1.n60 0.155672
R1411 VDD1.n61 VDD1.n36 0.155672
R1412 VDD1.n68 VDD1.n36 0.155672
R1413 VN.n2 VN.t1 178.02
R1414 VN.n10 VN.t5 178.02
R1415 VN.n13 VN.n8 161.3
R1416 VN.n12 VN.n11 161.3
R1417 VN.n5 VN.n0 161.3
R1418 VN.n4 VN.n3 161.3
R1419 VN.n6 VN.t4 158.721
R1420 VN.n14 VN.t2 158.721
R1421 VN.n1 VN.t0 128.031
R1422 VN.n9 VN.t3 128.031
R1423 VN.n15 VN.n14 80.6037
R1424 VN.n7 VN.n6 80.6037
R1425 VN.n2 VN.n1 45.4787
R1426 VN.n10 VN.n9 45.4787
R1427 VN VN.n15 40.0256
R1428 VN.n5 VN.n4 35.2488
R1429 VN.n13 VN.n12 35.2488
R1430 VN.n6 VN.n5 32.1338
R1431 VN.n14 VN.n13 32.1338
R1432 VN.n11 VN.n10 29.4552
R1433 VN.n3 VN.n2 29.4552
R1434 VN.n4 VN.n1 12.2964
R1435 VN.n12 VN.n9 12.2964
R1436 VN.n15 VN.n8 0.285035
R1437 VN.n7 VN.n0 0.285035
R1438 VN.n11 VN.n8 0.189894
R1439 VN.n3 VN.n0 0.189894
R1440 VN VN.n7 0.146778
R1441 VDD2.n67 VDD2.n37 289.615
R1442 VDD2.n30 VDD2.n0 289.615
R1443 VDD2.n68 VDD2.n67 185
R1444 VDD2.n66 VDD2.n65 185
R1445 VDD2.n41 VDD2.n40 185
R1446 VDD2.n60 VDD2.n59 185
R1447 VDD2.n58 VDD2.n57 185
R1448 VDD2.n45 VDD2.n44 185
R1449 VDD2.n52 VDD2.n51 185
R1450 VDD2.n50 VDD2.n49 185
R1451 VDD2.n13 VDD2.n12 185
R1452 VDD2.n15 VDD2.n14 185
R1453 VDD2.n8 VDD2.n7 185
R1454 VDD2.n21 VDD2.n20 185
R1455 VDD2.n23 VDD2.n22 185
R1456 VDD2.n4 VDD2.n3 185
R1457 VDD2.n29 VDD2.n28 185
R1458 VDD2.n31 VDD2.n30 185
R1459 VDD2.n48 VDD2.t3 147.659
R1460 VDD2.n11 VDD2.t4 147.659
R1461 VDD2.n67 VDD2.n66 104.615
R1462 VDD2.n66 VDD2.n40 104.615
R1463 VDD2.n59 VDD2.n40 104.615
R1464 VDD2.n59 VDD2.n58 104.615
R1465 VDD2.n58 VDD2.n44 104.615
R1466 VDD2.n51 VDD2.n44 104.615
R1467 VDD2.n51 VDD2.n50 104.615
R1468 VDD2.n14 VDD2.n13 104.615
R1469 VDD2.n14 VDD2.n7 104.615
R1470 VDD2.n21 VDD2.n7 104.615
R1471 VDD2.n22 VDD2.n21 104.615
R1472 VDD2.n22 VDD2.n3 104.615
R1473 VDD2.n29 VDD2.n3 104.615
R1474 VDD2.n30 VDD2.n29 104.615
R1475 VDD2.n36 VDD2.n35 67.9171
R1476 VDD2 VDD2.n73 67.9143
R1477 VDD2.n50 VDD2.t3 52.3082
R1478 VDD2.n13 VDD2.t4 52.3082
R1479 VDD2.n36 VDD2.n34 51.4013
R1480 VDD2.n72 VDD2.n71 50.4157
R1481 VDD2.n72 VDD2.n36 34.0881
R1482 VDD2.n49 VDD2.n48 15.6676
R1483 VDD2.n12 VDD2.n11 15.6676
R1484 VDD2.n52 VDD2.n47 12.8005
R1485 VDD2.n15 VDD2.n10 12.8005
R1486 VDD2.n53 VDD2.n45 12.0247
R1487 VDD2.n16 VDD2.n8 12.0247
R1488 VDD2.n57 VDD2.n56 11.249
R1489 VDD2.n20 VDD2.n19 11.249
R1490 VDD2.n60 VDD2.n43 10.4732
R1491 VDD2.n23 VDD2.n6 10.4732
R1492 VDD2.n61 VDD2.n41 9.69747
R1493 VDD2.n24 VDD2.n4 9.69747
R1494 VDD2.n71 VDD2.n70 9.45567
R1495 VDD2.n34 VDD2.n33 9.45567
R1496 VDD2.n70 VDD2.n69 9.3005
R1497 VDD2.n39 VDD2.n38 9.3005
R1498 VDD2.n64 VDD2.n63 9.3005
R1499 VDD2.n62 VDD2.n61 9.3005
R1500 VDD2.n43 VDD2.n42 9.3005
R1501 VDD2.n56 VDD2.n55 9.3005
R1502 VDD2.n54 VDD2.n53 9.3005
R1503 VDD2.n47 VDD2.n46 9.3005
R1504 VDD2.n2 VDD2.n1 9.3005
R1505 VDD2.n27 VDD2.n26 9.3005
R1506 VDD2.n25 VDD2.n24 9.3005
R1507 VDD2.n6 VDD2.n5 9.3005
R1508 VDD2.n19 VDD2.n18 9.3005
R1509 VDD2.n17 VDD2.n16 9.3005
R1510 VDD2.n10 VDD2.n9 9.3005
R1511 VDD2.n33 VDD2.n32 9.3005
R1512 VDD2.n65 VDD2.n64 8.92171
R1513 VDD2.n28 VDD2.n27 8.92171
R1514 VDD2.n68 VDD2.n39 8.14595
R1515 VDD2.n31 VDD2.n2 8.14595
R1516 VDD2.n69 VDD2.n37 7.3702
R1517 VDD2.n32 VDD2.n0 7.3702
R1518 VDD2.n71 VDD2.n37 6.59444
R1519 VDD2.n34 VDD2.n0 6.59444
R1520 VDD2.n69 VDD2.n68 5.81868
R1521 VDD2.n32 VDD2.n31 5.81868
R1522 VDD2.n65 VDD2.n39 5.04292
R1523 VDD2.n28 VDD2.n2 5.04292
R1524 VDD2.n48 VDD2.n46 4.38571
R1525 VDD2.n11 VDD2.n9 4.38571
R1526 VDD2.n64 VDD2.n41 4.26717
R1527 VDD2.n27 VDD2.n4 4.26717
R1528 VDD2.n61 VDD2.n60 3.49141
R1529 VDD2.n24 VDD2.n23 3.49141
R1530 VDD2.n73 VDD2.t2 2.91226
R1531 VDD2.n73 VDD2.t0 2.91226
R1532 VDD2.n35 VDD2.t5 2.91226
R1533 VDD2.n35 VDD2.t1 2.91226
R1534 VDD2.n57 VDD2.n43 2.71565
R1535 VDD2.n20 VDD2.n6 2.71565
R1536 VDD2.n56 VDD2.n45 1.93989
R1537 VDD2.n19 VDD2.n8 1.93989
R1538 VDD2.n53 VDD2.n52 1.16414
R1539 VDD2.n16 VDD2.n15 1.16414
R1540 VDD2 VDD2.n72 1.09964
R1541 VDD2.n49 VDD2.n47 0.388379
R1542 VDD2.n12 VDD2.n10 0.388379
R1543 VDD2.n70 VDD2.n38 0.155672
R1544 VDD2.n63 VDD2.n38 0.155672
R1545 VDD2.n63 VDD2.n62 0.155672
R1546 VDD2.n62 VDD2.n42 0.155672
R1547 VDD2.n55 VDD2.n42 0.155672
R1548 VDD2.n55 VDD2.n54 0.155672
R1549 VDD2.n54 VDD2.n46 0.155672
R1550 VDD2.n17 VDD2.n9 0.155672
R1551 VDD2.n18 VDD2.n17 0.155672
R1552 VDD2.n18 VDD2.n5 0.155672
R1553 VDD2.n25 VDD2.n5 0.155672
R1554 VDD2.n26 VDD2.n25 0.155672
R1555 VDD2.n26 VDD2.n1 0.155672
R1556 VDD2.n33 VDD2.n1 0.155672
C0 VN VP 4.67564f
C1 VN VDD2 3.31856f
C2 VP VDD1 3.51312f
C3 VN VTAIL 3.4612f
C4 VDD1 VDD2 0.922464f
C5 VTAIL VDD1 5.68171f
C6 VN VDD1 0.149128f
C7 VP VDD2 0.346145f
C8 VP VTAIL 3.4755f
C9 VTAIL VDD2 5.72363f
C10 VDD2 B 4.011139f
C11 VDD1 B 4.071072f
C12 VTAIL B 4.700381f
C13 VN B 8.608259f
C14 VP B 7.083687f
C15 VDD2.n0 B 0.032786f
C16 VDD2.n1 B 0.022055f
C17 VDD2.n2 B 0.011852f
C18 VDD2.n3 B 0.028013f
C19 VDD2.n4 B 0.012549f
C20 VDD2.n5 B 0.022055f
C21 VDD2.n6 B 0.011852f
C22 VDD2.n7 B 0.028013f
C23 VDD2.n8 B 0.012549f
C24 VDD2.n9 B 0.605821f
C25 VDD2.n10 B 0.011852f
C26 VDD2.t4 B 0.04566f
C27 VDD2.n11 B 0.098692f
C28 VDD2.n12 B 0.016548f
C29 VDD2.n13 B 0.02101f
C30 VDD2.n14 B 0.028013f
C31 VDD2.n15 B 0.012549f
C32 VDD2.n16 B 0.011852f
C33 VDD2.n17 B 0.022055f
C34 VDD2.n18 B 0.022055f
C35 VDD2.n19 B 0.011852f
C36 VDD2.n20 B 0.012549f
C37 VDD2.n21 B 0.028013f
C38 VDD2.n22 B 0.028013f
C39 VDD2.n23 B 0.012549f
C40 VDD2.n24 B 0.011852f
C41 VDD2.n25 B 0.022055f
C42 VDD2.n26 B 0.022055f
C43 VDD2.n27 B 0.011852f
C44 VDD2.n28 B 0.012549f
C45 VDD2.n29 B 0.028013f
C46 VDD2.n30 B 0.063801f
C47 VDD2.n31 B 0.012549f
C48 VDD2.n32 B 0.011852f
C49 VDD2.n33 B 0.05339f
C50 VDD2.n34 B 0.053501f
C51 VDD2.t5 B 0.118516f
C52 VDD2.t1 B 0.118516f
C53 VDD2.n35 B 1.00471f
C54 VDD2.n36 B 1.5828f
C55 VDD2.n37 B 0.032786f
C56 VDD2.n38 B 0.022055f
C57 VDD2.n39 B 0.011852f
C58 VDD2.n40 B 0.028013f
C59 VDD2.n41 B 0.012549f
C60 VDD2.n42 B 0.022055f
C61 VDD2.n43 B 0.011852f
C62 VDD2.n44 B 0.028013f
C63 VDD2.n45 B 0.012549f
C64 VDD2.n46 B 0.605821f
C65 VDD2.n47 B 0.011852f
C66 VDD2.t3 B 0.04566f
C67 VDD2.n48 B 0.098692f
C68 VDD2.n49 B 0.016548f
C69 VDD2.n50 B 0.02101f
C70 VDD2.n51 B 0.028013f
C71 VDD2.n52 B 0.012549f
C72 VDD2.n53 B 0.011852f
C73 VDD2.n54 B 0.022055f
C74 VDD2.n55 B 0.022055f
C75 VDD2.n56 B 0.011852f
C76 VDD2.n57 B 0.012549f
C77 VDD2.n58 B 0.028013f
C78 VDD2.n59 B 0.028013f
C79 VDD2.n60 B 0.012549f
C80 VDD2.n61 B 0.011852f
C81 VDD2.n62 B 0.022055f
C82 VDD2.n63 B 0.022055f
C83 VDD2.n64 B 0.011852f
C84 VDD2.n65 B 0.012549f
C85 VDD2.n66 B 0.028013f
C86 VDD2.n67 B 0.063801f
C87 VDD2.n68 B 0.012549f
C88 VDD2.n69 B 0.011852f
C89 VDD2.n70 B 0.05339f
C90 VDD2.n71 B 0.051307f
C91 VDD2.n72 B 1.58158f
C92 VDD2.t2 B 0.118516f
C93 VDD2.t0 B 0.118516f
C94 VDD2.n73 B 1.00469f
C95 VN.n0 B 0.049573f
C96 VN.t0 B 0.861786f
C97 VN.n1 B 0.384311f
C98 VN.t1 B 0.97963f
C99 VN.n2 B 0.400562f
C100 VN.n3 B 0.195438f
C101 VN.n4 B 0.057646f
C102 VN.n5 B 0.024238f
C103 VN.t4 B 0.934194f
C104 VN.n6 B 0.410578f
C105 VN.n7 B 0.034793f
C106 VN.n8 B 0.049573f
C107 VN.t3 B 0.861786f
C108 VN.n9 B 0.384311f
C109 VN.t5 B 0.97963f
C110 VN.n10 B 0.400562f
C111 VN.n11 B 0.195438f
C112 VN.n12 B 0.057646f
C113 VN.n13 B 0.024238f
C114 VN.t2 B 0.934194f
C115 VN.n14 B 0.410578f
C116 VN.n15 B 1.43013f
C117 VDD1.n0 B 0.033214f
C118 VDD1.n1 B 0.022343f
C119 VDD1.n2 B 0.012006f
C120 VDD1.n3 B 0.028378f
C121 VDD1.n4 B 0.012713f
C122 VDD1.n5 B 0.022343f
C123 VDD1.n6 B 0.012006f
C124 VDD1.n7 B 0.028378f
C125 VDD1.n8 B 0.012713f
C126 VDD1.n9 B 0.613729f
C127 VDD1.n10 B 0.012006f
C128 VDD1.t3 B 0.046256f
C129 VDD1.n11 B 0.09998f
C130 VDD1.n12 B 0.016764f
C131 VDD1.n13 B 0.021284f
C132 VDD1.n14 B 0.028378f
C133 VDD1.n15 B 0.012713f
C134 VDD1.n16 B 0.012006f
C135 VDD1.n17 B 0.022343f
C136 VDD1.n18 B 0.022343f
C137 VDD1.n19 B 0.012006f
C138 VDD1.n20 B 0.012713f
C139 VDD1.n21 B 0.028378f
C140 VDD1.n22 B 0.028378f
C141 VDD1.n23 B 0.012713f
C142 VDD1.n24 B 0.012006f
C143 VDD1.n25 B 0.022343f
C144 VDD1.n26 B 0.022343f
C145 VDD1.n27 B 0.012006f
C146 VDD1.n28 B 0.012713f
C147 VDD1.n29 B 0.028378f
C148 VDD1.n30 B 0.064634f
C149 VDD1.n31 B 0.012713f
C150 VDD1.n32 B 0.012006f
C151 VDD1.n33 B 0.054087f
C152 VDD1.n34 B 0.054613f
C153 VDD1.n35 B 0.033214f
C154 VDD1.n36 B 0.022343f
C155 VDD1.n37 B 0.012006f
C156 VDD1.n38 B 0.028378f
C157 VDD1.n39 B 0.012713f
C158 VDD1.n40 B 0.022343f
C159 VDD1.n41 B 0.012006f
C160 VDD1.n42 B 0.028378f
C161 VDD1.n43 B 0.012713f
C162 VDD1.n44 B 0.613729f
C163 VDD1.n45 B 0.012006f
C164 VDD1.t4 B 0.046256f
C165 VDD1.n46 B 0.09998f
C166 VDD1.n47 B 0.016764f
C167 VDD1.n48 B 0.021284f
C168 VDD1.n49 B 0.028378f
C169 VDD1.n50 B 0.012713f
C170 VDD1.n51 B 0.012006f
C171 VDD1.n52 B 0.022343f
C172 VDD1.n53 B 0.022343f
C173 VDD1.n54 B 0.012006f
C174 VDD1.n55 B 0.012713f
C175 VDD1.n56 B 0.028378f
C176 VDD1.n57 B 0.028378f
C177 VDD1.n58 B 0.012713f
C178 VDD1.n59 B 0.012006f
C179 VDD1.n60 B 0.022343f
C180 VDD1.n61 B 0.022343f
C181 VDD1.n62 B 0.012006f
C182 VDD1.n63 B 0.012713f
C183 VDD1.n64 B 0.028378f
C184 VDD1.n65 B 0.064634f
C185 VDD1.n66 B 0.012713f
C186 VDD1.n67 B 0.012006f
C187 VDD1.n68 B 0.054087f
C188 VDD1.n69 B 0.054199f
C189 VDD1.t1 B 0.120063f
C190 VDD1.t5 B 0.120063f
C191 VDD1.n70 B 1.01783f
C192 VDD1.n71 B 1.68192f
C193 VDD1.t0 B 0.120063f
C194 VDD1.t2 B 0.120063f
C195 VDD1.n72 B 1.01647f
C196 VDD1.n73 B 1.79525f
C197 VTAIL.t0 B 0.135883f
C198 VTAIL.t1 B 0.135883f
C199 VTAIL.n0 B 1.08426f
C200 VTAIL.n1 B 0.366507f
C201 VTAIL.n2 B 0.037591f
C202 VTAIL.n3 B 0.025287f
C203 VTAIL.n4 B 0.013588f
C204 VTAIL.n5 B 0.032118f
C205 VTAIL.n6 B 0.014388f
C206 VTAIL.n7 B 0.025287f
C207 VTAIL.n8 B 0.013588f
C208 VTAIL.n9 B 0.032118f
C209 VTAIL.n10 B 0.014388f
C210 VTAIL.n11 B 0.694598f
C211 VTAIL.n12 B 0.013588f
C212 VTAIL.t10 B 0.052351f
C213 VTAIL.n13 B 0.113154f
C214 VTAIL.n14 B 0.018973f
C215 VTAIL.n15 B 0.024088f
C216 VTAIL.n16 B 0.032118f
C217 VTAIL.n17 B 0.014388f
C218 VTAIL.n18 B 0.013588f
C219 VTAIL.n19 B 0.025287f
C220 VTAIL.n20 B 0.025287f
C221 VTAIL.n21 B 0.013588f
C222 VTAIL.n22 B 0.014388f
C223 VTAIL.n23 B 0.032118f
C224 VTAIL.n24 B 0.032118f
C225 VTAIL.n25 B 0.014388f
C226 VTAIL.n26 B 0.013588f
C227 VTAIL.n27 B 0.025287f
C228 VTAIL.n28 B 0.025287f
C229 VTAIL.n29 B 0.013588f
C230 VTAIL.n30 B 0.014388f
C231 VTAIL.n31 B 0.032118f
C232 VTAIL.n32 B 0.07315f
C233 VTAIL.n33 B 0.014388f
C234 VTAIL.n34 B 0.013588f
C235 VTAIL.n35 B 0.061214f
C236 VTAIL.n36 B 0.041386f
C237 VTAIL.n37 B 0.231077f
C238 VTAIL.t6 B 0.135883f
C239 VTAIL.t8 B 0.135883f
C240 VTAIL.n38 B 1.08426f
C241 VTAIL.n39 B 1.39909f
C242 VTAIL.t2 B 0.135883f
C243 VTAIL.t3 B 0.135883f
C244 VTAIL.n40 B 1.08427f
C245 VTAIL.n41 B 1.39908f
C246 VTAIL.n42 B 0.037591f
C247 VTAIL.n43 B 0.025287f
C248 VTAIL.n44 B 0.013588f
C249 VTAIL.n45 B 0.032118f
C250 VTAIL.n46 B 0.014388f
C251 VTAIL.n47 B 0.025287f
C252 VTAIL.n48 B 0.013588f
C253 VTAIL.n49 B 0.032118f
C254 VTAIL.n50 B 0.014388f
C255 VTAIL.n51 B 0.694598f
C256 VTAIL.n52 B 0.013588f
C257 VTAIL.t5 B 0.052351f
C258 VTAIL.n53 B 0.113154f
C259 VTAIL.n54 B 0.018973f
C260 VTAIL.n55 B 0.024088f
C261 VTAIL.n56 B 0.032118f
C262 VTAIL.n57 B 0.014388f
C263 VTAIL.n58 B 0.013588f
C264 VTAIL.n59 B 0.025287f
C265 VTAIL.n60 B 0.025287f
C266 VTAIL.n61 B 0.013588f
C267 VTAIL.n62 B 0.014388f
C268 VTAIL.n63 B 0.032118f
C269 VTAIL.n64 B 0.032118f
C270 VTAIL.n65 B 0.014388f
C271 VTAIL.n66 B 0.013588f
C272 VTAIL.n67 B 0.025287f
C273 VTAIL.n68 B 0.025287f
C274 VTAIL.n69 B 0.013588f
C275 VTAIL.n70 B 0.014388f
C276 VTAIL.n71 B 0.032118f
C277 VTAIL.n72 B 0.07315f
C278 VTAIL.n73 B 0.014388f
C279 VTAIL.n74 B 0.013588f
C280 VTAIL.n75 B 0.061214f
C281 VTAIL.n76 B 0.041386f
C282 VTAIL.n77 B 0.231077f
C283 VTAIL.t9 B 0.135883f
C284 VTAIL.t7 B 0.135883f
C285 VTAIL.n78 B 1.08427f
C286 VTAIL.n79 B 0.446576f
C287 VTAIL.n80 B 0.037591f
C288 VTAIL.n81 B 0.025287f
C289 VTAIL.n82 B 0.013588f
C290 VTAIL.n83 B 0.032118f
C291 VTAIL.n84 B 0.014388f
C292 VTAIL.n85 B 0.025287f
C293 VTAIL.n86 B 0.013588f
C294 VTAIL.n87 B 0.032118f
C295 VTAIL.n88 B 0.014388f
C296 VTAIL.n89 B 0.694598f
C297 VTAIL.n90 B 0.013588f
C298 VTAIL.t11 B 0.052351f
C299 VTAIL.n91 B 0.113154f
C300 VTAIL.n92 B 0.018973f
C301 VTAIL.n93 B 0.024088f
C302 VTAIL.n94 B 0.032118f
C303 VTAIL.n95 B 0.014388f
C304 VTAIL.n96 B 0.013588f
C305 VTAIL.n97 B 0.025287f
C306 VTAIL.n98 B 0.025287f
C307 VTAIL.n99 B 0.013588f
C308 VTAIL.n100 B 0.014388f
C309 VTAIL.n101 B 0.032118f
C310 VTAIL.n102 B 0.032118f
C311 VTAIL.n103 B 0.014388f
C312 VTAIL.n104 B 0.013588f
C313 VTAIL.n105 B 0.025287f
C314 VTAIL.n106 B 0.025287f
C315 VTAIL.n107 B 0.013588f
C316 VTAIL.n108 B 0.014388f
C317 VTAIL.n109 B 0.032118f
C318 VTAIL.n110 B 0.07315f
C319 VTAIL.n111 B 0.014388f
C320 VTAIL.n112 B 0.013588f
C321 VTAIL.n113 B 0.061214f
C322 VTAIL.n114 B 0.041386f
C323 VTAIL.n115 B 1.07049f
C324 VTAIL.n116 B 0.037591f
C325 VTAIL.n117 B 0.025287f
C326 VTAIL.n118 B 0.013588f
C327 VTAIL.n119 B 0.032118f
C328 VTAIL.n120 B 0.014388f
C329 VTAIL.n121 B 0.025287f
C330 VTAIL.n122 B 0.013588f
C331 VTAIL.n123 B 0.032118f
C332 VTAIL.n124 B 0.014388f
C333 VTAIL.n125 B 0.694598f
C334 VTAIL.n126 B 0.013588f
C335 VTAIL.t4 B 0.052351f
C336 VTAIL.n127 B 0.113154f
C337 VTAIL.n128 B 0.018973f
C338 VTAIL.n129 B 0.024088f
C339 VTAIL.n130 B 0.032118f
C340 VTAIL.n131 B 0.014388f
C341 VTAIL.n132 B 0.013588f
C342 VTAIL.n133 B 0.025287f
C343 VTAIL.n134 B 0.025287f
C344 VTAIL.n135 B 0.013588f
C345 VTAIL.n136 B 0.014388f
C346 VTAIL.n137 B 0.032118f
C347 VTAIL.n138 B 0.032118f
C348 VTAIL.n139 B 0.014388f
C349 VTAIL.n140 B 0.013588f
C350 VTAIL.n141 B 0.025287f
C351 VTAIL.n142 B 0.025287f
C352 VTAIL.n143 B 0.013588f
C353 VTAIL.n144 B 0.014388f
C354 VTAIL.n145 B 0.032118f
C355 VTAIL.n146 B 0.07315f
C356 VTAIL.n147 B 0.014388f
C357 VTAIL.n148 B 0.013588f
C358 VTAIL.n149 B 0.061214f
C359 VTAIL.n150 B 0.041386f
C360 VTAIL.n151 B 1.03748f
C361 VP.n0 B 0.050665f
C362 VP.t4 B 0.880773f
C363 VP.n1 B 0.343485f
C364 VP.n2 B 0.050665f
C365 VP.n3 B 0.050665f
C366 VP.t3 B 0.954777f
C367 VP.t5 B 0.880773f
C368 VP.n4 B 0.392779f
C369 VP.t2 B 1.00121f
C370 VP.n5 B 0.409387f
C371 VP.n6 B 0.199744f
C372 VP.n7 B 0.058916f
C373 VP.n8 B 0.024772f
C374 VP.n9 B 0.419624f
C375 VP.n10 B 1.44013f
C376 VP.n11 B 1.47457f
C377 VP.t1 B 0.954777f
C378 VP.n12 B 0.419624f
C379 VP.n13 B 0.024772f
C380 VP.n14 B 0.058916f
C381 VP.n15 B 0.037969f
C382 VP.n16 B 0.037969f
C383 VP.n17 B 0.058916f
C384 VP.n18 B 0.024772f
C385 VP.t0 B 0.954777f
C386 VP.n19 B 0.419624f
C387 VP.n20 B 0.03556f
.ends

