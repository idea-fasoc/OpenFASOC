* NGSPICE file created from diff_pair_sample_1593.ext - technology: sky130A

.subckt diff_pair_sample_1593 VTAIL VN VP B VDD2 VDD1
X0 B.t19 B.t17 B.t18 B.t7 sky130_fd_pr__nfet_01v8 ad=7.1253 pd=37.32 as=0 ps=0 w=18.27 l=2.29
X1 VDD1.t5 VP.t0 VTAIL.t7 B.t0 sky130_fd_pr__nfet_01v8 ad=3.01455 pd=18.6 as=7.1253 ps=37.32 w=18.27 l=2.29
X2 VTAIL.t9 VP.t1 VDD1.t4 B.t5 sky130_fd_pr__nfet_01v8 ad=3.01455 pd=18.6 as=3.01455 ps=18.6 w=18.27 l=2.29
X3 VDD2.t5 VN.t0 VTAIL.t2 B.t3 sky130_fd_pr__nfet_01v8 ad=7.1253 pd=37.32 as=3.01455 ps=18.6 w=18.27 l=2.29
X4 VDD1.t3 VP.t2 VTAIL.t11 B.t1 sky130_fd_pr__nfet_01v8 ad=3.01455 pd=18.6 as=7.1253 ps=37.32 w=18.27 l=2.29
X5 VDD2.t4 VN.t1 VTAIL.t5 B.t0 sky130_fd_pr__nfet_01v8 ad=3.01455 pd=18.6 as=7.1253 ps=37.32 w=18.27 l=2.29
X6 VTAIL.t6 VP.t3 VDD1.t2 B.t4 sky130_fd_pr__nfet_01v8 ad=3.01455 pd=18.6 as=3.01455 ps=18.6 w=18.27 l=2.29
X7 VTAIL.t4 VN.t2 VDD2.t3 B.t5 sky130_fd_pr__nfet_01v8 ad=3.01455 pd=18.6 as=3.01455 ps=18.6 w=18.27 l=2.29
X8 VTAIL.t3 VN.t3 VDD2.t2 B.t4 sky130_fd_pr__nfet_01v8 ad=3.01455 pd=18.6 as=3.01455 ps=18.6 w=18.27 l=2.29
X9 VDD1.t1 VP.t4 VTAIL.t8 B.t3 sky130_fd_pr__nfet_01v8 ad=7.1253 pd=37.32 as=3.01455 ps=18.6 w=18.27 l=2.29
X10 VDD1.t0 VP.t5 VTAIL.t10 B.t2 sky130_fd_pr__nfet_01v8 ad=7.1253 pd=37.32 as=3.01455 ps=18.6 w=18.27 l=2.29
X11 VDD2.t1 VN.t4 VTAIL.t1 B.t2 sky130_fd_pr__nfet_01v8 ad=7.1253 pd=37.32 as=3.01455 ps=18.6 w=18.27 l=2.29
X12 B.t16 B.t14 B.t15 B.t11 sky130_fd_pr__nfet_01v8 ad=7.1253 pd=37.32 as=0 ps=0 w=18.27 l=2.29
X13 B.t13 B.t10 B.t12 B.t11 sky130_fd_pr__nfet_01v8 ad=7.1253 pd=37.32 as=0 ps=0 w=18.27 l=2.29
X14 VDD2.t0 VN.t5 VTAIL.t0 B.t1 sky130_fd_pr__nfet_01v8 ad=3.01455 pd=18.6 as=7.1253 ps=37.32 w=18.27 l=2.29
X15 B.t9 B.t6 B.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=7.1253 pd=37.32 as=0 ps=0 w=18.27 l=2.29
R0 B.n972 B.n971 585
R1 B.n398 B.n138 585
R2 B.n397 B.n396 585
R3 B.n395 B.n394 585
R4 B.n393 B.n392 585
R5 B.n391 B.n390 585
R6 B.n389 B.n388 585
R7 B.n387 B.n386 585
R8 B.n385 B.n384 585
R9 B.n383 B.n382 585
R10 B.n381 B.n380 585
R11 B.n379 B.n378 585
R12 B.n377 B.n376 585
R13 B.n375 B.n374 585
R14 B.n373 B.n372 585
R15 B.n371 B.n370 585
R16 B.n369 B.n368 585
R17 B.n367 B.n366 585
R18 B.n365 B.n364 585
R19 B.n363 B.n362 585
R20 B.n361 B.n360 585
R21 B.n359 B.n358 585
R22 B.n357 B.n356 585
R23 B.n355 B.n354 585
R24 B.n353 B.n352 585
R25 B.n351 B.n350 585
R26 B.n349 B.n348 585
R27 B.n347 B.n346 585
R28 B.n345 B.n344 585
R29 B.n343 B.n342 585
R30 B.n341 B.n340 585
R31 B.n339 B.n338 585
R32 B.n337 B.n336 585
R33 B.n335 B.n334 585
R34 B.n333 B.n332 585
R35 B.n331 B.n330 585
R36 B.n329 B.n328 585
R37 B.n327 B.n326 585
R38 B.n325 B.n324 585
R39 B.n323 B.n322 585
R40 B.n321 B.n320 585
R41 B.n319 B.n318 585
R42 B.n317 B.n316 585
R43 B.n315 B.n314 585
R44 B.n313 B.n312 585
R45 B.n311 B.n310 585
R46 B.n309 B.n308 585
R47 B.n307 B.n306 585
R48 B.n305 B.n304 585
R49 B.n303 B.n302 585
R50 B.n301 B.n300 585
R51 B.n299 B.n298 585
R52 B.n297 B.n296 585
R53 B.n295 B.n294 585
R54 B.n293 B.n292 585
R55 B.n291 B.n290 585
R56 B.n289 B.n288 585
R57 B.n287 B.n286 585
R58 B.n285 B.n284 585
R59 B.n283 B.n282 585
R60 B.n281 B.n280 585
R61 B.n279 B.n278 585
R62 B.n277 B.n276 585
R63 B.n275 B.n274 585
R64 B.n273 B.n272 585
R65 B.n271 B.n270 585
R66 B.n269 B.n268 585
R67 B.n267 B.n266 585
R68 B.n265 B.n264 585
R69 B.n263 B.n262 585
R70 B.n261 B.n260 585
R71 B.n259 B.n258 585
R72 B.n257 B.n256 585
R73 B.n255 B.n254 585
R74 B.n253 B.n252 585
R75 B.n251 B.n250 585
R76 B.n249 B.n248 585
R77 B.n247 B.n246 585
R78 B.n245 B.n244 585
R79 B.n243 B.n242 585
R80 B.n241 B.n240 585
R81 B.n239 B.n238 585
R82 B.n237 B.n236 585
R83 B.n235 B.n234 585
R84 B.n233 B.n232 585
R85 B.n231 B.n230 585
R86 B.n229 B.n228 585
R87 B.n227 B.n226 585
R88 B.n225 B.n224 585
R89 B.n223 B.n222 585
R90 B.n221 B.n220 585
R91 B.n219 B.n218 585
R92 B.n217 B.n216 585
R93 B.n215 B.n214 585
R94 B.n213 B.n212 585
R95 B.n211 B.n210 585
R96 B.n209 B.n208 585
R97 B.n207 B.n206 585
R98 B.n205 B.n204 585
R99 B.n203 B.n202 585
R100 B.n201 B.n200 585
R101 B.n199 B.n198 585
R102 B.n197 B.n196 585
R103 B.n195 B.n194 585
R104 B.n193 B.n192 585
R105 B.n191 B.n190 585
R106 B.n189 B.n188 585
R107 B.n187 B.n186 585
R108 B.n185 B.n184 585
R109 B.n183 B.n182 585
R110 B.n181 B.n180 585
R111 B.n179 B.n178 585
R112 B.n177 B.n176 585
R113 B.n175 B.n174 585
R114 B.n173 B.n172 585
R115 B.n171 B.n170 585
R116 B.n169 B.n168 585
R117 B.n167 B.n166 585
R118 B.n165 B.n164 585
R119 B.n163 B.n162 585
R120 B.n161 B.n160 585
R121 B.n159 B.n158 585
R122 B.n157 B.n156 585
R123 B.n155 B.n154 585
R124 B.n153 B.n152 585
R125 B.n151 B.n150 585
R126 B.n149 B.n148 585
R127 B.n147 B.n146 585
R128 B.n74 B.n73 585
R129 B.n977 B.n976 585
R130 B.n970 B.n139 585
R131 B.n139 B.n71 585
R132 B.n969 B.n70 585
R133 B.n981 B.n70 585
R134 B.n968 B.n69 585
R135 B.n982 B.n69 585
R136 B.n967 B.n68 585
R137 B.n983 B.n68 585
R138 B.n966 B.n965 585
R139 B.n965 B.n64 585
R140 B.n964 B.n63 585
R141 B.n989 B.n63 585
R142 B.n963 B.n62 585
R143 B.n990 B.n62 585
R144 B.n962 B.n61 585
R145 B.n991 B.n61 585
R146 B.n961 B.n960 585
R147 B.n960 B.n57 585
R148 B.n959 B.n56 585
R149 B.n997 B.n56 585
R150 B.n958 B.n55 585
R151 B.n998 B.n55 585
R152 B.n957 B.n54 585
R153 B.n999 B.n54 585
R154 B.n956 B.n955 585
R155 B.n955 B.n50 585
R156 B.n954 B.n49 585
R157 B.n1005 B.n49 585
R158 B.n953 B.n48 585
R159 B.n1006 B.n48 585
R160 B.n952 B.n47 585
R161 B.n1007 B.n47 585
R162 B.n951 B.n950 585
R163 B.n950 B.n43 585
R164 B.n949 B.n42 585
R165 B.n1013 B.n42 585
R166 B.n948 B.n41 585
R167 B.n1014 B.n41 585
R168 B.n947 B.n40 585
R169 B.n1015 B.n40 585
R170 B.n946 B.n945 585
R171 B.n945 B.n36 585
R172 B.n944 B.n35 585
R173 B.n1021 B.n35 585
R174 B.n943 B.n34 585
R175 B.n1022 B.n34 585
R176 B.n942 B.n33 585
R177 B.n1023 B.n33 585
R178 B.n941 B.n940 585
R179 B.n940 B.n29 585
R180 B.n939 B.n28 585
R181 B.n1029 B.n28 585
R182 B.n938 B.n27 585
R183 B.n1030 B.n27 585
R184 B.n937 B.n26 585
R185 B.n1031 B.n26 585
R186 B.n936 B.n935 585
R187 B.n935 B.n22 585
R188 B.n934 B.n21 585
R189 B.n1037 B.n21 585
R190 B.n933 B.n20 585
R191 B.n1038 B.n20 585
R192 B.n932 B.n19 585
R193 B.n1039 B.n19 585
R194 B.n931 B.n930 585
R195 B.n930 B.n15 585
R196 B.n929 B.n14 585
R197 B.n1045 B.n14 585
R198 B.n928 B.n13 585
R199 B.n1046 B.n13 585
R200 B.n927 B.n12 585
R201 B.n1047 B.n12 585
R202 B.n926 B.n925 585
R203 B.n925 B.n8 585
R204 B.n924 B.n7 585
R205 B.n1053 B.n7 585
R206 B.n923 B.n6 585
R207 B.n1054 B.n6 585
R208 B.n922 B.n5 585
R209 B.n1055 B.n5 585
R210 B.n921 B.n920 585
R211 B.n920 B.n4 585
R212 B.n919 B.n399 585
R213 B.n919 B.n918 585
R214 B.n909 B.n400 585
R215 B.n401 B.n400 585
R216 B.n911 B.n910 585
R217 B.n912 B.n911 585
R218 B.n908 B.n406 585
R219 B.n406 B.n405 585
R220 B.n907 B.n906 585
R221 B.n906 B.n905 585
R222 B.n408 B.n407 585
R223 B.n409 B.n408 585
R224 B.n898 B.n897 585
R225 B.n899 B.n898 585
R226 B.n896 B.n414 585
R227 B.n414 B.n413 585
R228 B.n895 B.n894 585
R229 B.n894 B.n893 585
R230 B.n416 B.n415 585
R231 B.n417 B.n416 585
R232 B.n886 B.n885 585
R233 B.n887 B.n886 585
R234 B.n884 B.n422 585
R235 B.n422 B.n421 585
R236 B.n883 B.n882 585
R237 B.n882 B.n881 585
R238 B.n424 B.n423 585
R239 B.n425 B.n424 585
R240 B.n874 B.n873 585
R241 B.n875 B.n874 585
R242 B.n872 B.n430 585
R243 B.n430 B.n429 585
R244 B.n871 B.n870 585
R245 B.n870 B.n869 585
R246 B.n432 B.n431 585
R247 B.n433 B.n432 585
R248 B.n862 B.n861 585
R249 B.n863 B.n862 585
R250 B.n860 B.n437 585
R251 B.n441 B.n437 585
R252 B.n859 B.n858 585
R253 B.n858 B.n857 585
R254 B.n439 B.n438 585
R255 B.n440 B.n439 585
R256 B.n850 B.n849 585
R257 B.n851 B.n850 585
R258 B.n848 B.n446 585
R259 B.n446 B.n445 585
R260 B.n847 B.n846 585
R261 B.n846 B.n845 585
R262 B.n448 B.n447 585
R263 B.n449 B.n448 585
R264 B.n838 B.n837 585
R265 B.n839 B.n838 585
R266 B.n836 B.n454 585
R267 B.n454 B.n453 585
R268 B.n835 B.n834 585
R269 B.n834 B.n833 585
R270 B.n456 B.n455 585
R271 B.n457 B.n456 585
R272 B.n826 B.n825 585
R273 B.n827 B.n826 585
R274 B.n824 B.n462 585
R275 B.n462 B.n461 585
R276 B.n823 B.n822 585
R277 B.n822 B.n821 585
R278 B.n464 B.n463 585
R279 B.n465 B.n464 585
R280 B.n814 B.n813 585
R281 B.n815 B.n814 585
R282 B.n812 B.n470 585
R283 B.n470 B.n469 585
R284 B.n811 B.n810 585
R285 B.n810 B.n809 585
R286 B.n472 B.n471 585
R287 B.n473 B.n472 585
R288 B.n805 B.n804 585
R289 B.n476 B.n475 585
R290 B.n801 B.n800 585
R291 B.n802 B.n801 585
R292 B.n799 B.n541 585
R293 B.n798 B.n797 585
R294 B.n796 B.n795 585
R295 B.n794 B.n793 585
R296 B.n792 B.n791 585
R297 B.n790 B.n789 585
R298 B.n788 B.n787 585
R299 B.n786 B.n785 585
R300 B.n784 B.n783 585
R301 B.n782 B.n781 585
R302 B.n780 B.n779 585
R303 B.n778 B.n777 585
R304 B.n776 B.n775 585
R305 B.n774 B.n773 585
R306 B.n772 B.n771 585
R307 B.n770 B.n769 585
R308 B.n768 B.n767 585
R309 B.n766 B.n765 585
R310 B.n764 B.n763 585
R311 B.n762 B.n761 585
R312 B.n760 B.n759 585
R313 B.n758 B.n757 585
R314 B.n756 B.n755 585
R315 B.n754 B.n753 585
R316 B.n752 B.n751 585
R317 B.n750 B.n749 585
R318 B.n748 B.n747 585
R319 B.n746 B.n745 585
R320 B.n744 B.n743 585
R321 B.n742 B.n741 585
R322 B.n740 B.n739 585
R323 B.n738 B.n737 585
R324 B.n736 B.n735 585
R325 B.n734 B.n733 585
R326 B.n732 B.n731 585
R327 B.n730 B.n729 585
R328 B.n728 B.n727 585
R329 B.n726 B.n725 585
R330 B.n724 B.n723 585
R331 B.n722 B.n721 585
R332 B.n720 B.n719 585
R333 B.n718 B.n717 585
R334 B.n716 B.n715 585
R335 B.n714 B.n713 585
R336 B.n712 B.n711 585
R337 B.n710 B.n709 585
R338 B.n708 B.n707 585
R339 B.n706 B.n705 585
R340 B.n704 B.n703 585
R341 B.n702 B.n701 585
R342 B.n700 B.n699 585
R343 B.n698 B.n697 585
R344 B.n696 B.n695 585
R345 B.n694 B.n693 585
R346 B.n692 B.n691 585
R347 B.n690 B.n689 585
R348 B.n688 B.n687 585
R349 B.n685 B.n684 585
R350 B.n683 B.n682 585
R351 B.n681 B.n680 585
R352 B.n679 B.n678 585
R353 B.n677 B.n676 585
R354 B.n675 B.n674 585
R355 B.n673 B.n672 585
R356 B.n671 B.n670 585
R357 B.n669 B.n668 585
R358 B.n667 B.n666 585
R359 B.n664 B.n663 585
R360 B.n662 B.n661 585
R361 B.n660 B.n659 585
R362 B.n658 B.n657 585
R363 B.n656 B.n655 585
R364 B.n654 B.n653 585
R365 B.n652 B.n651 585
R366 B.n650 B.n649 585
R367 B.n648 B.n647 585
R368 B.n646 B.n645 585
R369 B.n644 B.n643 585
R370 B.n642 B.n641 585
R371 B.n640 B.n639 585
R372 B.n638 B.n637 585
R373 B.n636 B.n635 585
R374 B.n634 B.n633 585
R375 B.n632 B.n631 585
R376 B.n630 B.n629 585
R377 B.n628 B.n627 585
R378 B.n626 B.n625 585
R379 B.n624 B.n623 585
R380 B.n622 B.n621 585
R381 B.n620 B.n619 585
R382 B.n618 B.n617 585
R383 B.n616 B.n615 585
R384 B.n614 B.n613 585
R385 B.n612 B.n611 585
R386 B.n610 B.n609 585
R387 B.n608 B.n607 585
R388 B.n606 B.n605 585
R389 B.n604 B.n603 585
R390 B.n602 B.n601 585
R391 B.n600 B.n599 585
R392 B.n598 B.n597 585
R393 B.n596 B.n595 585
R394 B.n594 B.n593 585
R395 B.n592 B.n591 585
R396 B.n590 B.n589 585
R397 B.n588 B.n587 585
R398 B.n586 B.n585 585
R399 B.n584 B.n583 585
R400 B.n582 B.n581 585
R401 B.n580 B.n579 585
R402 B.n578 B.n577 585
R403 B.n576 B.n575 585
R404 B.n574 B.n573 585
R405 B.n572 B.n571 585
R406 B.n570 B.n569 585
R407 B.n568 B.n567 585
R408 B.n566 B.n565 585
R409 B.n564 B.n563 585
R410 B.n562 B.n561 585
R411 B.n560 B.n559 585
R412 B.n558 B.n557 585
R413 B.n556 B.n555 585
R414 B.n554 B.n553 585
R415 B.n552 B.n551 585
R416 B.n550 B.n549 585
R417 B.n548 B.n547 585
R418 B.n546 B.n540 585
R419 B.n802 B.n540 585
R420 B.n806 B.n474 585
R421 B.n474 B.n473 585
R422 B.n808 B.n807 585
R423 B.n809 B.n808 585
R424 B.n468 B.n467 585
R425 B.n469 B.n468 585
R426 B.n817 B.n816 585
R427 B.n816 B.n815 585
R428 B.n818 B.n466 585
R429 B.n466 B.n465 585
R430 B.n820 B.n819 585
R431 B.n821 B.n820 585
R432 B.n460 B.n459 585
R433 B.n461 B.n460 585
R434 B.n829 B.n828 585
R435 B.n828 B.n827 585
R436 B.n830 B.n458 585
R437 B.n458 B.n457 585
R438 B.n832 B.n831 585
R439 B.n833 B.n832 585
R440 B.n452 B.n451 585
R441 B.n453 B.n452 585
R442 B.n841 B.n840 585
R443 B.n840 B.n839 585
R444 B.n842 B.n450 585
R445 B.n450 B.n449 585
R446 B.n844 B.n843 585
R447 B.n845 B.n844 585
R448 B.n444 B.n443 585
R449 B.n445 B.n444 585
R450 B.n853 B.n852 585
R451 B.n852 B.n851 585
R452 B.n854 B.n442 585
R453 B.n442 B.n440 585
R454 B.n856 B.n855 585
R455 B.n857 B.n856 585
R456 B.n436 B.n435 585
R457 B.n441 B.n436 585
R458 B.n865 B.n864 585
R459 B.n864 B.n863 585
R460 B.n866 B.n434 585
R461 B.n434 B.n433 585
R462 B.n868 B.n867 585
R463 B.n869 B.n868 585
R464 B.n428 B.n427 585
R465 B.n429 B.n428 585
R466 B.n877 B.n876 585
R467 B.n876 B.n875 585
R468 B.n878 B.n426 585
R469 B.n426 B.n425 585
R470 B.n880 B.n879 585
R471 B.n881 B.n880 585
R472 B.n420 B.n419 585
R473 B.n421 B.n420 585
R474 B.n889 B.n888 585
R475 B.n888 B.n887 585
R476 B.n890 B.n418 585
R477 B.n418 B.n417 585
R478 B.n892 B.n891 585
R479 B.n893 B.n892 585
R480 B.n412 B.n411 585
R481 B.n413 B.n412 585
R482 B.n901 B.n900 585
R483 B.n900 B.n899 585
R484 B.n902 B.n410 585
R485 B.n410 B.n409 585
R486 B.n904 B.n903 585
R487 B.n905 B.n904 585
R488 B.n404 B.n403 585
R489 B.n405 B.n404 585
R490 B.n914 B.n913 585
R491 B.n913 B.n912 585
R492 B.n915 B.n402 585
R493 B.n402 B.n401 585
R494 B.n917 B.n916 585
R495 B.n918 B.n917 585
R496 B.n2 B.n0 585
R497 B.n4 B.n2 585
R498 B.n3 B.n1 585
R499 B.n1054 B.n3 585
R500 B.n1052 B.n1051 585
R501 B.n1053 B.n1052 585
R502 B.n1050 B.n9 585
R503 B.n9 B.n8 585
R504 B.n1049 B.n1048 585
R505 B.n1048 B.n1047 585
R506 B.n11 B.n10 585
R507 B.n1046 B.n11 585
R508 B.n1044 B.n1043 585
R509 B.n1045 B.n1044 585
R510 B.n1042 B.n16 585
R511 B.n16 B.n15 585
R512 B.n1041 B.n1040 585
R513 B.n1040 B.n1039 585
R514 B.n18 B.n17 585
R515 B.n1038 B.n18 585
R516 B.n1036 B.n1035 585
R517 B.n1037 B.n1036 585
R518 B.n1034 B.n23 585
R519 B.n23 B.n22 585
R520 B.n1033 B.n1032 585
R521 B.n1032 B.n1031 585
R522 B.n25 B.n24 585
R523 B.n1030 B.n25 585
R524 B.n1028 B.n1027 585
R525 B.n1029 B.n1028 585
R526 B.n1026 B.n30 585
R527 B.n30 B.n29 585
R528 B.n1025 B.n1024 585
R529 B.n1024 B.n1023 585
R530 B.n32 B.n31 585
R531 B.n1022 B.n32 585
R532 B.n1020 B.n1019 585
R533 B.n1021 B.n1020 585
R534 B.n1018 B.n37 585
R535 B.n37 B.n36 585
R536 B.n1017 B.n1016 585
R537 B.n1016 B.n1015 585
R538 B.n39 B.n38 585
R539 B.n1014 B.n39 585
R540 B.n1012 B.n1011 585
R541 B.n1013 B.n1012 585
R542 B.n1010 B.n44 585
R543 B.n44 B.n43 585
R544 B.n1009 B.n1008 585
R545 B.n1008 B.n1007 585
R546 B.n46 B.n45 585
R547 B.n1006 B.n46 585
R548 B.n1004 B.n1003 585
R549 B.n1005 B.n1004 585
R550 B.n1002 B.n51 585
R551 B.n51 B.n50 585
R552 B.n1001 B.n1000 585
R553 B.n1000 B.n999 585
R554 B.n53 B.n52 585
R555 B.n998 B.n53 585
R556 B.n996 B.n995 585
R557 B.n997 B.n996 585
R558 B.n994 B.n58 585
R559 B.n58 B.n57 585
R560 B.n993 B.n992 585
R561 B.n992 B.n991 585
R562 B.n60 B.n59 585
R563 B.n990 B.n60 585
R564 B.n988 B.n987 585
R565 B.n989 B.n988 585
R566 B.n986 B.n65 585
R567 B.n65 B.n64 585
R568 B.n985 B.n984 585
R569 B.n984 B.n983 585
R570 B.n67 B.n66 585
R571 B.n982 B.n67 585
R572 B.n980 B.n979 585
R573 B.n981 B.n980 585
R574 B.n978 B.n72 585
R575 B.n72 B.n71 585
R576 B.n1057 B.n1056 585
R577 B.n1056 B.n1055 585
R578 B.n804 B.n474 463.671
R579 B.n976 B.n72 463.671
R580 B.n540 B.n472 463.671
R581 B.n972 B.n139 463.671
R582 B.n544 B.t16 441.142
R583 B.n542 B.t13 441.142
R584 B.n143 B.t18 441.142
R585 B.n140 B.t8 441.142
R586 B.n544 B.t14 399.8
R587 B.n542 B.t10 399.8
R588 B.n143 B.t17 399.8
R589 B.n140 B.t6 399.8
R590 B.n545 B.t15 390.329
R591 B.n141 B.t9 390.329
R592 B.n543 B.t12 390.329
R593 B.n144 B.t19 390.329
R594 B.n974 B.n973 256.663
R595 B.n974 B.n137 256.663
R596 B.n974 B.n136 256.663
R597 B.n974 B.n135 256.663
R598 B.n974 B.n134 256.663
R599 B.n974 B.n133 256.663
R600 B.n974 B.n132 256.663
R601 B.n974 B.n131 256.663
R602 B.n974 B.n130 256.663
R603 B.n974 B.n129 256.663
R604 B.n974 B.n128 256.663
R605 B.n974 B.n127 256.663
R606 B.n974 B.n126 256.663
R607 B.n974 B.n125 256.663
R608 B.n974 B.n124 256.663
R609 B.n974 B.n123 256.663
R610 B.n974 B.n122 256.663
R611 B.n974 B.n121 256.663
R612 B.n974 B.n120 256.663
R613 B.n974 B.n119 256.663
R614 B.n974 B.n118 256.663
R615 B.n974 B.n117 256.663
R616 B.n974 B.n116 256.663
R617 B.n974 B.n115 256.663
R618 B.n974 B.n114 256.663
R619 B.n974 B.n113 256.663
R620 B.n974 B.n112 256.663
R621 B.n974 B.n111 256.663
R622 B.n974 B.n110 256.663
R623 B.n974 B.n109 256.663
R624 B.n974 B.n108 256.663
R625 B.n974 B.n107 256.663
R626 B.n974 B.n106 256.663
R627 B.n974 B.n105 256.663
R628 B.n974 B.n104 256.663
R629 B.n974 B.n103 256.663
R630 B.n974 B.n102 256.663
R631 B.n974 B.n101 256.663
R632 B.n974 B.n100 256.663
R633 B.n974 B.n99 256.663
R634 B.n974 B.n98 256.663
R635 B.n974 B.n97 256.663
R636 B.n974 B.n96 256.663
R637 B.n974 B.n95 256.663
R638 B.n974 B.n94 256.663
R639 B.n974 B.n93 256.663
R640 B.n974 B.n92 256.663
R641 B.n974 B.n91 256.663
R642 B.n974 B.n90 256.663
R643 B.n974 B.n89 256.663
R644 B.n974 B.n88 256.663
R645 B.n974 B.n87 256.663
R646 B.n974 B.n86 256.663
R647 B.n974 B.n85 256.663
R648 B.n974 B.n84 256.663
R649 B.n974 B.n83 256.663
R650 B.n974 B.n82 256.663
R651 B.n974 B.n81 256.663
R652 B.n974 B.n80 256.663
R653 B.n974 B.n79 256.663
R654 B.n974 B.n78 256.663
R655 B.n974 B.n77 256.663
R656 B.n974 B.n76 256.663
R657 B.n974 B.n75 256.663
R658 B.n975 B.n974 256.663
R659 B.n803 B.n802 256.663
R660 B.n802 B.n477 256.663
R661 B.n802 B.n478 256.663
R662 B.n802 B.n479 256.663
R663 B.n802 B.n480 256.663
R664 B.n802 B.n481 256.663
R665 B.n802 B.n482 256.663
R666 B.n802 B.n483 256.663
R667 B.n802 B.n484 256.663
R668 B.n802 B.n485 256.663
R669 B.n802 B.n486 256.663
R670 B.n802 B.n487 256.663
R671 B.n802 B.n488 256.663
R672 B.n802 B.n489 256.663
R673 B.n802 B.n490 256.663
R674 B.n802 B.n491 256.663
R675 B.n802 B.n492 256.663
R676 B.n802 B.n493 256.663
R677 B.n802 B.n494 256.663
R678 B.n802 B.n495 256.663
R679 B.n802 B.n496 256.663
R680 B.n802 B.n497 256.663
R681 B.n802 B.n498 256.663
R682 B.n802 B.n499 256.663
R683 B.n802 B.n500 256.663
R684 B.n802 B.n501 256.663
R685 B.n802 B.n502 256.663
R686 B.n802 B.n503 256.663
R687 B.n802 B.n504 256.663
R688 B.n802 B.n505 256.663
R689 B.n802 B.n506 256.663
R690 B.n802 B.n507 256.663
R691 B.n802 B.n508 256.663
R692 B.n802 B.n509 256.663
R693 B.n802 B.n510 256.663
R694 B.n802 B.n511 256.663
R695 B.n802 B.n512 256.663
R696 B.n802 B.n513 256.663
R697 B.n802 B.n514 256.663
R698 B.n802 B.n515 256.663
R699 B.n802 B.n516 256.663
R700 B.n802 B.n517 256.663
R701 B.n802 B.n518 256.663
R702 B.n802 B.n519 256.663
R703 B.n802 B.n520 256.663
R704 B.n802 B.n521 256.663
R705 B.n802 B.n522 256.663
R706 B.n802 B.n523 256.663
R707 B.n802 B.n524 256.663
R708 B.n802 B.n525 256.663
R709 B.n802 B.n526 256.663
R710 B.n802 B.n527 256.663
R711 B.n802 B.n528 256.663
R712 B.n802 B.n529 256.663
R713 B.n802 B.n530 256.663
R714 B.n802 B.n531 256.663
R715 B.n802 B.n532 256.663
R716 B.n802 B.n533 256.663
R717 B.n802 B.n534 256.663
R718 B.n802 B.n535 256.663
R719 B.n802 B.n536 256.663
R720 B.n802 B.n537 256.663
R721 B.n802 B.n538 256.663
R722 B.n802 B.n539 256.663
R723 B.n808 B.n474 163.367
R724 B.n808 B.n468 163.367
R725 B.n816 B.n468 163.367
R726 B.n816 B.n466 163.367
R727 B.n820 B.n466 163.367
R728 B.n820 B.n460 163.367
R729 B.n828 B.n460 163.367
R730 B.n828 B.n458 163.367
R731 B.n832 B.n458 163.367
R732 B.n832 B.n452 163.367
R733 B.n840 B.n452 163.367
R734 B.n840 B.n450 163.367
R735 B.n844 B.n450 163.367
R736 B.n844 B.n444 163.367
R737 B.n852 B.n444 163.367
R738 B.n852 B.n442 163.367
R739 B.n856 B.n442 163.367
R740 B.n856 B.n436 163.367
R741 B.n864 B.n436 163.367
R742 B.n864 B.n434 163.367
R743 B.n868 B.n434 163.367
R744 B.n868 B.n428 163.367
R745 B.n876 B.n428 163.367
R746 B.n876 B.n426 163.367
R747 B.n880 B.n426 163.367
R748 B.n880 B.n420 163.367
R749 B.n888 B.n420 163.367
R750 B.n888 B.n418 163.367
R751 B.n892 B.n418 163.367
R752 B.n892 B.n412 163.367
R753 B.n900 B.n412 163.367
R754 B.n900 B.n410 163.367
R755 B.n904 B.n410 163.367
R756 B.n904 B.n404 163.367
R757 B.n913 B.n404 163.367
R758 B.n913 B.n402 163.367
R759 B.n917 B.n402 163.367
R760 B.n917 B.n2 163.367
R761 B.n1056 B.n2 163.367
R762 B.n1056 B.n3 163.367
R763 B.n1052 B.n3 163.367
R764 B.n1052 B.n9 163.367
R765 B.n1048 B.n9 163.367
R766 B.n1048 B.n11 163.367
R767 B.n1044 B.n11 163.367
R768 B.n1044 B.n16 163.367
R769 B.n1040 B.n16 163.367
R770 B.n1040 B.n18 163.367
R771 B.n1036 B.n18 163.367
R772 B.n1036 B.n23 163.367
R773 B.n1032 B.n23 163.367
R774 B.n1032 B.n25 163.367
R775 B.n1028 B.n25 163.367
R776 B.n1028 B.n30 163.367
R777 B.n1024 B.n30 163.367
R778 B.n1024 B.n32 163.367
R779 B.n1020 B.n32 163.367
R780 B.n1020 B.n37 163.367
R781 B.n1016 B.n37 163.367
R782 B.n1016 B.n39 163.367
R783 B.n1012 B.n39 163.367
R784 B.n1012 B.n44 163.367
R785 B.n1008 B.n44 163.367
R786 B.n1008 B.n46 163.367
R787 B.n1004 B.n46 163.367
R788 B.n1004 B.n51 163.367
R789 B.n1000 B.n51 163.367
R790 B.n1000 B.n53 163.367
R791 B.n996 B.n53 163.367
R792 B.n996 B.n58 163.367
R793 B.n992 B.n58 163.367
R794 B.n992 B.n60 163.367
R795 B.n988 B.n60 163.367
R796 B.n988 B.n65 163.367
R797 B.n984 B.n65 163.367
R798 B.n984 B.n67 163.367
R799 B.n980 B.n67 163.367
R800 B.n980 B.n72 163.367
R801 B.n801 B.n476 163.367
R802 B.n801 B.n541 163.367
R803 B.n797 B.n796 163.367
R804 B.n793 B.n792 163.367
R805 B.n789 B.n788 163.367
R806 B.n785 B.n784 163.367
R807 B.n781 B.n780 163.367
R808 B.n777 B.n776 163.367
R809 B.n773 B.n772 163.367
R810 B.n769 B.n768 163.367
R811 B.n765 B.n764 163.367
R812 B.n761 B.n760 163.367
R813 B.n757 B.n756 163.367
R814 B.n753 B.n752 163.367
R815 B.n749 B.n748 163.367
R816 B.n745 B.n744 163.367
R817 B.n741 B.n740 163.367
R818 B.n737 B.n736 163.367
R819 B.n733 B.n732 163.367
R820 B.n729 B.n728 163.367
R821 B.n725 B.n724 163.367
R822 B.n721 B.n720 163.367
R823 B.n717 B.n716 163.367
R824 B.n713 B.n712 163.367
R825 B.n709 B.n708 163.367
R826 B.n705 B.n704 163.367
R827 B.n701 B.n700 163.367
R828 B.n697 B.n696 163.367
R829 B.n693 B.n692 163.367
R830 B.n689 B.n688 163.367
R831 B.n684 B.n683 163.367
R832 B.n680 B.n679 163.367
R833 B.n676 B.n675 163.367
R834 B.n672 B.n671 163.367
R835 B.n668 B.n667 163.367
R836 B.n663 B.n662 163.367
R837 B.n659 B.n658 163.367
R838 B.n655 B.n654 163.367
R839 B.n651 B.n650 163.367
R840 B.n647 B.n646 163.367
R841 B.n643 B.n642 163.367
R842 B.n639 B.n638 163.367
R843 B.n635 B.n634 163.367
R844 B.n631 B.n630 163.367
R845 B.n627 B.n626 163.367
R846 B.n623 B.n622 163.367
R847 B.n619 B.n618 163.367
R848 B.n615 B.n614 163.367
R849 B.n611 B.n610 163.367
R850 B.n607 B.n606 163.367
R851 B.n603 B.n602 163.367
R852 B.n599 B.n598 163.367
R853 B.n595 B.n594 163.367
R854 B.n591 B.n590 163.367
R855 B.n587 B.n586 163.367
R856 B.n583 B.n582 163.367
R857 B.n579 B.n578 163.367
R858 B.n575 B.n574 163.367
R859 B.n571 B.n570 163.367
R860 B.n567 B.n566 163.367
R861 B.n563 B.n562 163.367
R862 B.n559 B.n558 163.367
R863 B.n555 B.n554 163.367
R864 B.n551 B.n550 163.367
R865 B.n547 B.n540 163.367
R866 B.n810 B.n472 163.367
R867 B.n810 B.n470 163.367
R868 B.n814 B.n470 163.367
R869 B.n814 B.n464 163.367
R870 B.n822 B.n464 163.367
R871 B.n822 B.n462 163.367
R872 B.n826 B.n462 163.367
R873 B.n826 B.n456 163.367
R874 B.n834 B.n456 163.367
R875 B.n834 B.n454 163.367
R876 B.n838 B.n454 163.367
R877 B.n838 B.n448 163.367
R878 B.n846 B.n448 163.367
R879 B.n846 B.n446 163.367
R880 B.n850 B.n446 163.367
R881 B.n850 B.n439 163.367
R882 B.n858 B.n439 163.367
R883 B.n858 B.n437 163.367
R884 B.n862 B.n437 163.367
R885 B.n862 B.n432 163.367
R886 B.n870 B.n432 163.367
R887 B.n870 B.n430 163.367
R888 B.n874 B.n430 163.367
R889 B.n874 B.n424 163.367
R890 B.n882 B.n424 163.367
R891 B.n882 B.n422 163.367
R892 B.n886 B.n422 163.367
R893 B.n886 B.n416 163.367
R894 B.n894 B.n416 163.367
R895 B.n894 B.n414 163.367
R896 B.n898 B.n414 163.367
R897 B.n898 B.n408 163.367
R898 B.n906 B.n408 163.367
R899 B.n906 B.n406 163.367
R900 B.n911 B.n406 163.367
R901 B.n911 B.n400 163.367
R902 B.n919 B.n400 163.367
R903 B.n920 B.n919 163.367
R904 B.n920 B.n5 163.367
R905 B.n6 B.n5 163.367
R906 B.n7 B.n6 163.367
R907 B.n925 B.n7 163.367
R908 B.n925 B.n12 163.367
R909 B.n13 B.n12 163.367
R910 B.n14 B.n13 163.367
R911 B.n930 B.n14 163.367
R912 B.n930 B.n19 163.367
R913 B.n20 B.n19 163.367
R914 B.n21 B.n20 163.367
R915 B.n935 B.n21 163.367
R916 B.n935 B.n26 163.367
R917 B.n27 B.n26 163.367
R918 B.n28 B.n27 163.367
R919 B.n940 B.n28 163.367
R920 B.n940 B.n33 163.367
R921 B.n34 B.n33 163.367
R922 B.n35 B.n34 163.367
R923 B.n945 B.n35 163.367
R924 B.n945 B.n40 163.367
R925 B.n41 B.n40 163.367
R926 B.n42 B.n41 163.367
R927 B.n950 B.n42 163.367
R928 B.n950 B.n47 163.367
R929 B.n48 B.n47 163.367
R930 B.n49 B.n48 163.367
R931 B.n955 B.n49 163.367
R932 B.n955 B.n54 163.367
R933 B.n55 B.n54 163.367
R934 B.n56 B.n55 163.367
R935 B.n960 B.n56 163.367
R936 B.n960 B.n61 163.367
R937 B.n62 B.n61 163.367
R938 B.n63 B.n62 163.367
R939 B.n965 B.n63 163.367
R940 B.n965 B.n68 163.367
R941 B.n69 B.n68 163.367
R942 B.n70 B.n69 163.367
R943 B.n139 B.n70 163.367
R944 B.n146 B.n74 163.367
R945 B.n150 B.n149 163.367
R946 B.n154 B.n153 163.367
R947 B.n158 B.n157 163.367
R948 B.n162 B.n161 163.367
R949 B.n166 B.n165 163.367
R950 B.n170 B.n169 163.367
R951 B.n174 B.n173 163.367
R952 B.n178 B.n177 163.367
R953 B.n182 B.n181 163.367
R954 B.n186 B.n185 163.367
R955 B.n190 B.n189 163.367
R956 B.n194 B.n193 163.367
R957 B.n198 B.n197 163.367
R958 B.n202 B.n201 163.367
R959 B.n206 B.n205 163.367
R960 B.n210 B.n209 163.367
R961 B.n214 B.n213 163.367
R962 B.n218 B.n217 163.367
R963 B.n222 B.n221 163.367
R964 B.n226 B.n225 163.367
R965 B.n230 B.n229 163.367
R966 B.n234 B.n233 163.367
R967 B.n238 B.n237 163.367
R968 B.n242 B.n241 163.367
R969 B.n246 B.n245 163.367
R970 B.n250 B.n249 163.367
R971 B.n254 B.n253 163.367
R972 B.n258 B.n257 163.367
R973 B.n262 B.n261 163.367
R974 B.n266 B.n265 163.367
R975 B.n270 B.n269 163.367
R976 B.n274 B.n273 163.367
R977 B.n278 B.n277 163.367
R978 B.n282 B.n281 163.367
R979 B.n286 B.n285 163.367
R980 B.n290 B.n289 163.367
R981 B.n294 B.n293 163.367
R982 B.n298 B.n297 163.367
R983 B.n302 B.n301 163.367
R984 B.n306 B.n305 163.367
R985 B.n310 B.n309 163.367
R986 B.n314 B.n313 163.367
R987 B.n318 B.n317 163.367
R988 B.n322 B.n321 163.367
R989 B.n326 B.n325 163.367
R990 B.n330 B.n329 163.367
R991 B.n334 B.n333 163.367
R992 B.n338 B.n337 163.367
R993 B.n342 B.n341 163.367
R994 B.n346 B.n345 163.367
R995 B.n350 B.n349 163.367
R996 B.n354 B.n353 163.367
R997 B.n358 B.n357 163.367
R998 B.n362 B.n361 163.367
R999 B.n366 B.n365 163.367
R1000 B.n370 B.n369 163.367
R1001 B.n374 B.n373 163.367
R1002 B.n378 B.n377 163.367
R1003 B.n382 B.n381 163.367
R1004 B.n386 B.n385 163.367
R1005 B.n390 B.n389 163.367
R1006 B.n394 B.n393 163.367
R1007 B.n396 B.n138 163.367
R1008 B.n804 B.n803 71.676
R1009 B.n541 B.n477 71.676
R1010 B.n796 B.n478 71.676
R1011 B.n792 B.n479 71.676
R1012 B.n788 B.n480 71.676
R1013 B.n784 B.n481 71.676
R1014 B.n780 B.n482 71.676
R1015 B.n776 B.n483 71.676
R1016 B.n772 B.n484 71.676
R1017 B.n768 B.n485 71.676
R1018 B.n764 B.n486 71.676
R1019 B.n760 B.n487 71.676
R1020 B.n756 B.n488 71.676
R1021 B.n752 B.n489 71.676
R1022 B.n748 B.n490 71.676
R1023 B.n744 B.n491 71.676
R1024 B.n740 B.n492 71.676
R1025 B.n736 B.n493 71.676
R1026 B.n732 B.n494 71.676
R1027 B.n728 B.n495 71.676
R1028 B.n724 B.n496 71.676
R1029 B.n720 B.n497 71.676
R1030 B.n716 B.n498 71.676
R1031 B.n712 B.n499 71.676
R1032 B.n708 B.n500 71.676
R1033 B.n704 B.n501 71.676
R1034 B.n700 B.n502 71.676
R1035 B.n696 B.n503 71.676
R1036 B.n692 B.n504 71.676
R1037 B.n688 B.n505 71.676
R1038 B.n683 B.n506 71.676
R1039 B.n679 B.n507 71.676
R1040 B.n675 B.n508 71.676
R1041 B.n671 B.n509 71.676
R1042 B.n667 B.n510 71.676
R1043 B.n662 B.n511 71.676
R1044 B.n658 B.n512 71.676
R1045 B.n654 B.n513 71.676
R1046 B.n650 B.n514 71.676
R1047 B.n646 B.n515 71.676
R1048 B.n642 B.n516 71.676
R1049 B.n638 B.n517 71.676
R1050 B.n634 B.n518 71.676
R1051 B.n630 B.n519 71.676
R1052 B.n626 B.n520 71.676
R1053 B.n622 B.n521 71.676
R1054 B.n618 B.n522 71.676
R1055 B.n614 B.n523 71.676
R1056 B.n610 B.n524 71.676
R1057 B.n606 B.n525 71.676
R1058 B.n602 B.n526 71.676
R1059 B.n598 B.n527 71.676
R1060 B.n594 B.n528 71.676
R1061 B.n590 B.n529 71.676
R1062 B.n586 B.n530 71.676
R1063 B.n582 B.n531 71.676
R1064 B.n578 B.n532 71.676
R1065 B.n574 B.n533 71.676
R1066 B.n570 B.n534 71.676
R1067 B.n566 B.n535 71.676
R1068 B.n562 B.n536 71.676
R1069 B.n558 B.n537 71.676
R1070 B.n554 B.n538 71.676
R1071 B.n550 B.n539 71.676
R1072 B.n976 B.n975 71.676
R1073 B.n146 B.n75 71.676
R1074 B.n150 B.n76 71.676
R1075 B.n154 B.n77 71.676
R1076 B.n158 B.n78 71.676
R1077 B.n162 B.n79 71.676
R1078 B.n166 B.n80 71.676
R1079 B.n170 B.n81 71.676
R1080 B.n174 B.n82 71.676
R1081 B.n178 B.n83 71.676
R1082 B.n182 B.n84 71.676
R1083 B.n186 B.n85 71.676
R1084 B.n190 B.n86 71.676
R1085 B.n194 B.n87 71.676
R1086 B.n198 B.n88 71.676
R1087 B.n202 B.n89 71.676
R1088 B.n206 B.n90 71.676
R1089 B.n210 B.n91 71.676
R1090 B.n214 B.n92 71.676
R1091 B.n218 B.n93 71.676
R1092 B.n222 B.n94 71.676
R1093 B.n226 B.n95 71.676
R1094 B.n230 B.n96 71.676
R1095 B.n234 B.n97 71.676
R1096 B.n238 B.n98 71.676
R1097 B.n242 B.n99 71.676
R1098 B.n246 B.n100 71.676
R1099 B.n250 B.n101 71.676
R1100 B.n254 B.n102 71.676
R1101 B.n258 B.n103 71.676
R1102 B.n262 B.n104 71.676
R1103 B.n266 B.n105 71.676
R1104 B.n270 B.n106 71.676
R1105 B.n274 B.n107 71.676
R1106 B.n278 B.n108 71.676
R1107 B.n282 B.n109 71.676
R1108 B.n286 B.n110 71.676
R1109 B.n290 B.n111 71.676
R1110 B.n294 B.n112 71.676
R1111 B.n298 B.n113 71.676
R1112 B.n302 B.n114 71.676
R1113 B.n306 B.n115 71.676
R1114 B.n310 B.n116 71.676
R1115 B.n314 B.n117 71.676
R1116 B.n318 B.n118 71.676
R1117 B.n322 B.n119 71.676
R1118 B.n326 B.n120 71.676
R1119 B.n330 B.n121 71.676
R1120 B.n334 B.n122 71.676
R1121 B.n338 B.n123 71.676
R1122 B.n342 B.n124 71.676
R1123 B.n346 B.n125 71.676
R1124 B.n350 B.n126 71.676
R1125 B.n354 B.n127 71.676
R1126 B.n358 B.n128 71.676
R1127 B.n362 B.n129 71.676
R1128 B.n366 B.n130 71.676
R1129 B.n370 B.n131 71.676
R1130 B.n374 B.n132 71.676
R1131 B.n378 B.n133 71.676
R1132 B.n382 B.n134 71.676
R1133 B.n386 B.n135 71.676
R1134 B.n390 B.n136 71.676
R1135 B.n394 B.n137 71.676
R1136 B.n973 B.n138 71.676
R1137 B.n973 B.n972 71.676
R1138 B.n396 B.n137 71.676
R1139 B.n393 B.n136 71.676
R1140 B.n389 B.n135 71.676
R1141 B.n385 B.n134 71.676
R1142 B.n381 B.n133 71.676
R1143 B.n377 B.n132 71.676
R1144 B.n373 B.n131 71.676
R1145 B.n369 B.n130 71.676
R1146 B.n365 B.n129 71.676
R1147 B.n361 B.n128 71.676
R1148 B.n357 B.n127 71.676
R1149 B.n353 B.n126 71.676
R1150 B.n349 B.n125 71.676
R1151 B.n345 B.n124 71.676
R1152 B.n341 B.n123 71.676
R1153 B.n337 B.n122 71.676
R1154 B.n333 B.n121 71.676
R1155 B.n329 B.n120 71.676
R1156 B.n325 B.n119 71.676
R1157 B.n321 B.n118 71.676
R1158 B.n317 B.n117 71.676
R1159 B.n313 B.n116 71.676
R1160 B.n309 B.n115 71.676
R1161 B.n305 B.n114 71.676
R1162 B.n301 B.n113 71.676
R1163 B.n297 B.n112 71.676
R1164 B.n293 B.n111 71.676
R1165 B.n289 B.n110 71.676
R1166 B.n285 B.n109 71.676
R1167 B.n281 B.n108 71.676
R1168 B.n277 B.n107 71.676
R1169 B.n273 B.n106 71.676
R1170 B.n269 B.n105 71.676
R1171 B.n265 B.n104 71.676
R1172 B.n261 B.n103 71.676
R1173 B.n257 B.n102 71.676
R1174 B.n253 B.n101 71.676
R1175 B.n249 B.n100 71.676
R1176 B.n245 B.n99 71.676
R1177 B.n241 B.n98 71.676
R1178 B.n237 B.n97 71.676
R1179 B.n233 B.n96 71.676
R1180 B.n229 B.n95 71.676
R1181 B.n225 B.n94 71.676
R1182 B.n221 B.n93 71.676
R1183 B.n217 B.n92 71.676
R1184 B.n213 B.n91 71.676
R1185 B.n209 B.n90 71.676
R1186 B.n205 B.n89 71.676
R1187 B.n201 B.n88 71.676
R1188 B.n197 B.n87 71.676
R1189 B.n193 B.n86 71.676
R1190 B.n189 B.n85 71.676
R1191 B.n185 B.n84 71.676
R1192 B.n181 B.n83 71.676
R1193 B.n177 B.n82 71.676
R1194 B.n173 B.n81 71.676
R1195 B.n169 B.n80 71.676
R1196 B.n165 B.n79 71.676
R1197 B.n161 B.n78 71.676
R1198 B.n157 B.n77 71.676
R1199 B.n153 B.n76 71.676
R1200 B.n149 B.n75 71.676
R1201 B.n975 B.n74 71.676
R1202 B.n803 B.n476 71.676
R1203 B.n797 B.n477 71.676
R1204 B.n793 B.n478 71.676
R1205 B.n789 B.n479 71.676
R1206 B.n785 B.n480 71.676
R1207 B.n781 B.n481 71.676
R1208 B.n777 B.n482 71.676
R1209 B.n773 B.n483 71.676
R1210 B.n769 B.n484 71.676
R1211 B.n765 B.n485 71.676
R1212 B.n761 B.n486 71.676
R1213 B.n757 B.n487 71.676
R1214 B.n753 B.n488 71.676
R1215 B.n749 B.n489 71.676
R1216 B.n745 B.n490 71.676
R1217 B.n741 B.n491 71.676
R1218 B.n737 B.n492 71.676
R1219 B.n733 B.n493 71.676
R1220 B.n729 B.n494 71.676
R1221 B.n725 B.n495 71.676
R1222 B.n721 B.n496 71.676
R1223 B.n717 B.n497 71.676
R1224 B.n713 B.n498 71.676
R1225 B.n709 B.n499 71.676
R1226 B.n705 B.n500 71.676
R1227 B.n701 B.n501 71.676
R1228 B.n697 B.n502 71.676
R1229 B.n693 B.n503 71.676
R1230 B.n689 B.n504 71.676
R1231 B.n684 B.n505 71.676
R1232 B.n680 B.n506 71.676
R1233 B.n676 B.n507 71.676
R1234 B.n672 B.n508 71.676
R1235 B.n668 B.n509 71.676
R1236 B.n663 B.n510 71.676
R1237 B.n659 B.n511 71.676
R1238 B.n655 B.n512 71.676
R1239 B.n651 B.n513 71.676
R1240 B.n647 B.n514 71.676
R1241 B.n643 B.n515 71.676
R1242 B.n639 B.n516 71.676
R1243 B.n635 B.n517 71.676
R1244 B.n631 B.n518 71.676
R1245 B.n627 B.n519 71.676
R1246 B.n623 B.n520 71.676
R1247 B.n619 B.n521 71.676
R1248 B.n615 B.n522 71.676
R1249 B.n611 B.n523 71.676
R1250 B.n607 B.n524 71.676
R1251 B.n603 B.n525 71.676
R1252 B.n599 B.n526 71.676
R1253 B.n595 B.n527 71.676
R1254 B.n591 B.n528 71.676
R1255 B.n587 B.n529 71.676
R1256 B.n583 B.n530 71.676
R1257 B.n579 B.n531 71.676
R1258 B.n575 B.n532 71.676
R1259 B.n571 B.n533 71.676
R1260 B.n567 B.n534 71.676
R1261 B.n563 B.n535 71.676
R1262 B.n559 B.n536 71.676
R1263 B.n555 B.n537 71.676
R1264 B.n551 B.n538 71.676
R1265 B.n547 B.n539 71.676
R1266 B.n665 B.n545 59.5399
R1267 B.n686 B.n543 59.5399
R1268 B.n145 B.n144 59.5399
R1269 B.n142 B.n141 59.5399
R1270 B.n802 B.n473 55.5962
R1271 B.n974 B.n71 55.5962
R1272 B.n545 B.n544 50.8126
R1273 B.n543 B.n542 50.8126
R1274 B.n144 B.n143 50.8126
R1275 B.n141 B.n140 50.8126
R1276 B.n809 B.n473 31.7695
R1277 B.n809 B.n469 31.7695
R1278 B.n815 B.n469 31.7695
R1279 B.n815 B.n465 31.7695
R1280 B.n821 B.n465 31.7695
R1281 B.n821 B.n461 31.7695
R1282 B.n827 B.n461 31.7695
R1283 B.n833 B.n457 31.7695
R1284 B.n833 B.n453 31.7695
R1285 B.n839 B.n453 31.7695
R1286 B.n839 B.n449 31.7695
R1287 B.n845 B.n449 31.7695
R1288 B.n845 B.n445 31.7695
R1289 B.n851 B.n445 31.7695
R1290 B.n851 B.n440 31.7695
R1291 B.n857 B.n440 31.7695
R1292 B.n857 B.n441 31.7695
R1293 B.n863 B.n433 31.7695
R1294 B.n869 B.n433 31.7695
R1295 B.n869 B.n429 31.7695
R1296 B.n875 B.n429 31.7695
R1297 B.n875 B.n425 31.7695
R1298 B.n881 B.n425 31.7695
R1299 B.n887 B.n421 31.7695
R1300 B.n887 B.n417 31.7695
R1301 B.n893 B.n417 31.7695
R1302 B.n893 B.n413 31.7695
R1303 B.n899 B.n413 31.7695
R1304 B.n899 B.n409 31.7695
R1305 B.n905 B.n409 31.7695
R1306 B.n912 B.n405 31.7695
R1307 B.n912 B.n401 31.7695
R1308 B.n918 B.n401 31.7695
R1309 B.n918 B.n4 31.7695
R1310 B.n1055 B.n4 31.7695
R1311 B.n1055 B.n1054 31.7695
R1312 B.n1054 B.n1053 31.7695
R1313 B.n1053 B.n8 31.7695
R1314 B.n1047 B.n8 31.7695
R1315 B.n1047 B.n1046 31.7695
R1316 B.n1045 B.n15 31.7695
R1317 B.n1039 B.n15 31.7695
R1318 B.n1039 B.n1038 31.7695
R1319 B.n1038 B.n1037 31.7695
R1320 B.n1037 B.n22 31.7695
R1321 B.n1031 B.n22 31.7695
R1322 B.n1031 B.n1030 31.7695
R1323 B.n1029 B.n29 31.7695
R1324 B.n1023 B.n29 31.7695
R1325 B.n1023 B.n1022 31.7695
R1326 B.n1022 B.n1021 31.7695
R1327 B.n1021 B.n36 31.7695
R1328 B.n1015 B.n36 31.7695
R1329 B.n1014 B.n1013 31.7695
R1330 B.n1013 B.n43 31.7695
R1331 B.n1007 B.n43 31.7695
R1332 B.n1007 B.n1006 31.7695
R1333 B.n1006 B.n1005 31.7695
R1334 B.n1005 B.n50 31.7695
R1335 B.n999 B.n50 31.7695
R1336 B.n999 B.n998 31.7695
R1337 B.n998 B.n997 31.7695
R1338 B.n997 B.n57 31.7695
R1339 B.n991 B.n990 31.7695
R1340 B.n990 B.n989 31.7695
R1341 B.n989 B.n64 31.7695
R1342 B.n983 B.n64 31.7695
R1343 B.n983 B.n982 31.7695
R1344 B.n982 B.n981 31.7695
R1345 B.n981 B.n71 31.7695
R1346 B.n978 B.n977 30.1273
R1347 B.n971 B.n970 30.1273
R1348 B.n546 B.n471 30.1273
R1349 B.n806 B.n805 30.1273
R1350 B.n863 B.t3 27.5647
R1351 B.n1015 B.t0 27.5647
R1352 B.n881 B.t5 26.6304
R1353 B.t4 B.n1029 26.6304
R1354 B.t11 B.n457 24.7616
R1355 B.t7 B.n57 24.7616
R1356 B B.n1057 18.0485
R1357 B.n905 B.t1 17.2865
R1358 B.t2 B.n1045 17.2865
R1359 B.t1 B.n405 14.4834
R1360 B.n1046 B.t2 14.4834
R1361 B.n977 B.n73 10.6151
R1362 B.n147 B.n73 10.6151
R1363 B.n148 B.n147 10.6151
R1364 B.n151 B.n148 10.6151
R1365 B.n152 B.n151 10.6151
R1366 B.n155 B.n152 10.6151
R1367 B.n156 B.n155 10.6151
R1368 B.n159 B.n156 10.6151
R1369 B.n160 B.n159 10.6151
R1370 B.n163 B.n160 10.6151
R1371 B.n164 B.n163 10.6151
R1372 B.n167 B.n164 10.6151
R1373 B.n168 B.n167 10.6151
R1374 B.n171 B.n168 10.6151
R1375 B.n172 B.n171 10.6151
R1376 B.n175 B.n172 10.6151
R1377 B.n176 B.n175 10.6151
R1378 B.n179 B.n176 10.6151
R1379 B.n180 B.n179 10.6151
R1380 B.n183 B.n180 10.6151
R1381 B.n184 B.n183 10.6151
R1382 B.n187 B.n184 10.6151
R1383 B.n188 B.n187 10.6151
R1384 B.n191 B.n188 10.6151
R1385 B.n192 B.n191 10.6151
R1386 B.n195 B.n192 10.6151
R1387 B.n196 B.n195 10.6151
R1388 B.n199 B.n196 10.6151
R1389 B.n200 B.n199 10.6151
R1390 B.n203 B.n200 10.6151
R1391 B.n204 B.n203 10.6151
R1392 B.n207 B.n204 10.6151
R1393 B.n208 B.n207 10.6151
R1394 B.n211 B.n208 10.6151
R1395 B.n212 B.n211 10.6151
R1396 B.n215 B.n212 10.6151
R1397 B.n216 B.n215 10.6151
R1398 B.n219 B.n216 10.6151
R1399 B.n220 B.n219 10.6151
R1400 B.n223 B.n220 10.6151
R1401 B.n224 B.n223 10.6151
R1402 B.n227 B.n224 10.6151
R1403 B.n228 B.n227 10.6151
R1404 B.n231 B.n228 10.6151
R1405 B.n232 B.n231 10.6151
R1406 B.n235 B.n232 10.6151
R1407 B.n236 B.n235 10.6151
R1408 B.n239 B.n236 10.6151
R1409 B.n240 B.n239 10.6151
R1410 B.n243 B.n240 10.6151
R1411 B.n244 B.n243 10.6151
R1412 B.n247 B.n244 10.6151
R1413 B.n248 B.n247 10.6151
R1414 B.n251 B.n248 10.6151
R1415 B.n252 B.n251 10.6151
R1416 B.n255 B.n252 10.6151
R1417 B.n256 B.n255 10.6151
R1418 B.n259 B.n256 10.6151
R1419 B.n260 B.n259 10.6151
R1420 B.n264 B.n263 10.6151
R1421 B.n267 B.n264 10.6151
R1422 B.n268 B.n267 10.6151
R1423 B.n271 B.n268 10.6151
R1424 B.n272 B.n271 10.6151
R1425 B.n275 B.n272 10.6151
R1426 B.n276 B.n275 10.6151
R1427 B.n279 B.n276 10.6151
R1428 B.n280 B.n279 10.6151
R1429 B.n284 B.n283 10.6151
R1430 B.n287 B.n284 10.6151
R1431 B.n288 B.n287 10.6151
R1432 B.n291 B.n288 10.6151
R1433 B.n292 B.n291 10.6151
R1434 B.n295 B.n292 10.6151
R1435 B.n296 B.n295 10.6151
R1436 B.n299 B.n296 10.6151
R1437 B.n300 B.n299 10.6151
R1438 B.n303 B.n300 10.6151
R1439 B.n304 B.n303 10.6151
R1440 B.n307 B.n304 10.6151
R1441 B.n308 B.n307 10.6151
R1442 B.n311 B.n308 10.6151
R1443 B.n312 B.n311 10.6151
R1444 B.n315 B.n312 10.6151
R1445 B.n316 B.n315 10.6151
R1446 B.n319 B.n316 10.6151
R1447 B.n320 B.n319 10.6151
R1448 B.n323 B.n320 10.6151
R1449 B.n324 B.n323 10.6151
R1450 B.n327 B.n324 10.6151
R1451 B.n328 B.n327 10.6151
R1452 B.n331 B.n328 10.6151
R1453 B.n332 B.n331 10.6151
R1454 B.n335 B.n332 10.6151
R1455 B.n336 B.n335 10.6151
R1456 B.n339 B.n336 10.6151
R1457 B.n340 B.n339 10.6151
R1458 B.n343 B.n340 10.6151
R1459 B.n344 B.n343 10.6151
R1460 B.n347 B.n344 10.6151
R1461 B.n348 B.n347 10.6151
R1462 B.n351 B.n348 10.6151
R1463 B.n352 B.n351 10.6151
R1464 B.n355 B.n352 10.6151
R1465 B.n356 B.n355 10.6151
R1466 B.n359 B.n356 10.6151
R1467 B.n360 B.n359 10.6151
R1468 B.n363 B.n360 10.6151
R1469 B.n364 B.n363 10.6151
R1470 B.n367 B.n364 10.6151
R1471 B.n368 B.n367 10.6151
R1472 B.n371 B.n368 10.6151
R1473 B.n372 B.n371 10.6151
R1474 B.n375 B.n372 10.6151
R1475 B.n376 B.n375 10.6151
R1476 B.n379 B.n376 10.6151
R1477 B.n380 B.n379 10.6151
R1478 B.n383 B.n380 10.6151
R1479 B.n384 B.n383 10.6151
R1480 B.n387 B.n384 10.6151
R1481 B.n388 B.n387 10.6151
R1482 B.n391 B.n388 10.6151
R1483 B.n392 B.n391 10.6151
R1484 B.n395 B.n392 10.6151
R1485 B.n397 B.n395 10.6151
R1486 B.n398 B.n397 10.6151
R1487 B.n971 B.n398 10.6151
R1488 B.n811 B.n471 10.6151
R1489 B.n812 B.n811 10.6151
R1490 B.n813 B.n812 10.6151
R1491 B.n813 B.n463 10.6151
R1492 B.n823 B.n463 10.6151
R1493 B.n824 B.n823 10.6151
R1494 B.n825 B.n824 10.6151
R1495 B.n825 B.n455 10.6151
R1496 B.n835 B.n455 10.6151
R1497 B.n836 B.n835 10.6151
R1498 B.n837 B.n836 10.6151
R1499 B.n837 B.n447 10.6151
R1500 B.n847 B.n447 10.6151
R1501 B.n848 B.n847 10.6151
R1502 B.n849 B.n848 10.6151
R1503 B.n849 B.n438 10.6151
R1504 B.n859 B.n438 10.6151
R1505 B.n860 B.n859 10.6151
R1506 B.n861 B.n860 10.6151
R1507 B.n861 B.n431 10.6151
R1508 B.n871 B.n431 10.6151
R1509 B.n872 B.n871 10.6151
R1510 B.n873 B.n872 10.6151
R1511 B.n873 B.n423 10.6151
R1512 B.n883 B.n423 10.6151
R1513 B.n884 B.n883 10.6151
R1514 B.n885 B.n884 10.6151
R1515 B.n885 B.n415 10.6151
R1516 B.n895 B.n415 10.6151
R1517 B.n896 B.n895 10.6151
R1518 B.n897 B.n896 10.6151
R1519 B.n897 B.n407 10.6151
R1520 B.n907 B.n407 10.6151
R1521 B.n908 B.n907 10.6151
R1522 B.n910 B.n908 10.6151
R1523 B.n910 B.n909 10.6151
R1524 B.n909 B.n399 10.6151
R1525 B.n921 B.n399 10.6151
R1526 B.n922 B.n921 10.6151
R1527 B.n923 B.n922 10.6151
R1528 B.n924 B.n923 10.6151
R1529 B.n926 B.n924 10.6151
R1530 B.n927 B.n926 10.6151
R1531 B.n928 B.n927 10.6151
R1532 B.n929 B.n928 10.6151
R1533 B.n931 B.n929 10.6151
R1534 B.n932 B.n931 10.6151
R1535 B.n933 B.n932 10.6151
R1536 B.n934 B.n933 10.6151
R1537 B.n936 B.n934 10.6151
R1538 B.n937 B.n936 10.6151
R1539 B.n938 B.n937 10.6151
R1540 B.n939 B.n938 10.6151
R1541 B.n941 B.n939 10.6151
R1542 B.n942 B.n941 10.6151
R1543 B.n943 B.n942 10.6151
R1544 B.n944 B.n943 10.6151
R1545 B.n946 B.n944 10.6151
R1546 B.n947 B.n946 10.6151
R1547 B.n948 B.n947 10.6151
R1548 B.n949 B.n948 10.6151
R1549 B.n951 B.n949 10.6151
R1550 B.n952 B.n951 10.6151
R1551 B.n953 B.n952 10.6151
R1552 B.n954 B.n953 10.6151
R1553 B.n956 B.n954 10.6151
R1554 B.n957 B.n956 10.6151
R1555 B.n958 B.n957 10.6151
R1556 B.n959 B.n958 10.6151
R1557 B.n961 B.n959 10.6151
R1558 B.n962 B.n961 10.6151
R1559 B.n963 B.n962 10.6151
R1560 B.n964 B.n963 10.6151
R1561 B.n966 B.n964 10.6151
R1562 B.n967 B.n966 10.6151
R1563 B.n968 B.n967 10.6151
R1564 B.n969 B.n968 10.6151
R1565 B.n970 B.n969 10.6151
R1566 B.n805 B.n475 10.6151
R1567 B.n800 B.n475 10.6151
R1568 B.n800 B.n799 10.6151
R1569 B.n799 B.n798 10.6151
R1570 B.n798 B.n795 10.6151
R1571 B.n795 B.n794 10.6151
R1572 B.n794 B.n791 10.6151
R1573 B.n791 B.n790 10.6151
R1574 B.n790 B.n787 10.6151
R1575 B.n787 B.n786 10.6151
R1576 B.n786 B.n783 10.6151
R1577 B.n783 B.n782 10.6151
R1578 B.n782 B.n779 10.6151
R1579 B.n779 B.n778 10.6151
R1580 B.n778 B.n775 10.6151
R1581 B.n775 B.n774 10.6151
R1582 B.n774 B.n771 10.6151
R1583 B.n771 B.n770 10.6151
R1584 B.n770 B.n767 10.6151
R1585 B.n767 B.n766 10.6151
R1586 B.n766 B.n763 10.6151
R1587 B.n763 B.n762 10.6151
R1588 B.n762 B.n759 10.6151
R1589 B.n759 B.n758 10.6151
R1590 B.n758 B.n755 10.6151
R1591 B.n755 B.n754 10.6151
R1592 B.n754 B.n751 10.6151
R1593 B.n751 B.n750 10.6151
R1594 B.n750 B.n747 10.6151
R1595 B.n747 B.n746 10.6151
R1596 B.n746 B.n743 10.6151
R1597 B.n743 B.n742 10.6151
R1598 B.n742 B.n739 10.6151
R1599 B.n739 B.n738 10.6151
R1600 B.n738 B.n735 10.6151
R1601 B.n735 B.n734 10.6151
R1602 B.n734 B.n731 10.6151
R1603 B.n731 B.n730 10.6151
R1604 B.n730 B.n727 10.6151
R1605 B.n727 B.n726 10.6151
R1606 B.n726 B.n723 10.6151
R1607 B.n723 B.n722 10.6151
R1608 B.n722 B.n719 10.6151
R1609 B.n719 B.n718 10.6151
R1610 B.n718 B.n715 10.6151
R1611 B.n715 B.n714 10.6151
R1612 B.n714 B.n711 10.6151
R1613 B.n711 B.n710 10.6151
R1614 B.n710 B.n707 10.6151
R1615 B.n707 B.n706 10.6151
R1616 B.n706 B.n703 10.6151
R1617 B.n703 B.n702 10.6151
R1618 B.n702 B.n699 10.6151
R1619 B.n699 B.n698 10.6151
R1620 B.n698 B.n695 10.6151
R1621 B.n695 B.n694 10.6151
R1622 B.n694 B.n691 10.6151
R1623 B.n691 B.n690 10.6151
R1624 B.n690 B.n687 10.6151
R1625 B.n685 B.n682 10.6151
R1626 B.n682 B.n681 10.6151
R1627 B.n681 B.n678 10.6151
R1628 B.n678 B.n677 10.6151
R1629 B.n677 B.n674 10.6151
R1630 B.n674 B.n673 10.6151
R1631 B.n673 B.n670 10.6151
R1632 B.n670 B.n669 10.6151
R1633 B.n669 B.n666 10.6151
R1634 B.n664 B.n661 10.6151
R1635 B.n661 B.n660 10.6151
R1636 B.n660 B.n657 10.6151
R1637 B.n657 B.n656 10.6151
R1638 B.n656 B.n653 10.6151
R1639 B.n653 B.n652 10.6151
R1640 B.n652 B.n649 10.6151
R1641 B.n649 B.n648 10.6151
R1642 B.n648 B.n645 10.6151
R1643 B.n645 B.n644 10.6151
R1644 B.n644 B.n641 10.6151
R1645 B.n641 B.n640 10.6151
R1646 B.n640 B.n637 10.6151
R1647 B.n637 B.n636 10.6151
R1648 B.n636 B.n633 10.6151
R1649 B.n633 B.n632 10.6151
R1650 B.n632 B.n629 10.6151
R1651 B.n629 B.n628 10.6151
R1652 B.n628 B.n625 10.6151
R1653 B.n625 B.n624 10.6151
R1654 B.n624 B.n621 10.6151
R1655 B.n621 B.n620 10.6151
R1656 B.n620 B.n617 10.6151
R1657 B.n617 B.n616 10.6151
R1658 B.n616 B.n613 10.6151
R1659 B.n613 B.n612 10.6151
R1660 B.n612 B.n609 10.6151
R1661 B.n609 B.n608 10.6151
R1662 B.n608 B.n605 10.6151
R1663 B.n605 B.n604 10.6151
R1664 B.n604 B.n601 10.6151
R1665 B.n601 B.n600 10.6151
R1666 B.n600 B.n597 10.6151
R1667 B.n597 B.n596 10.6151
R1668 B.n596 B.n593 10.6151
R1669 B.n593 B.n592 10.6151
R1670 B.n592 B.n589 10.6151
R1671 B.n589 B.n588 10.6151
R1672 B.n588 B.n585 10.6151
R1673 B.n585 B.n584 10.6151
R1674 B.n584 B.n581 10.6151
R1675 B.n581 B.n580 10.6151
R1676 B.n580 B.n577 10.6151
R1677 B.n577 B.n576 10.6151
R1678 B.n576 B.n573 10.6151
R1679 B.n573 B.n572 10.6151
R1680 B.n572 B.n569 10.6151
R1681 B.n569 B.n568 10.6151
R1682 B.n568 B.n565 10.6151
R1683 B.n565 B.n564 10.6151
R1684 B.n564 B.n561 10.6151
R1685 B.n561 B.n560 10.6151
R1686 B.n560 B.n557 10.6151
R1687 B.n557 B.n556 10.6151
R1688 B.n556 B.n553 10.6151
R1689 B.n553 B.n552 10.6151
R1690 B.n552 B.n549 10.6151
R1691 B.n549 B.n548 10.6151
R1692 B.n548 B.n546 10.6151
R1693 B.n807 B.n806 10.6151
R1694 B.n807 B.n467 10.6151
R1695 B.n817 B.n467 10.6151
R1696 B.n818 B.n817 10.6151
R1697 B.n819 B.n818 10.6151
R1698 B.n819 B.n459 10.6151
R1699 B.n829 B.n459 10.6151
R1700 B.n830 B.n829 10.6151
R1701 B.n831 B.n830 10.6151
R1702 B.n831 B.n451 10.6151
R1703 B.n841 B.n451 10.6151
R1704 B.n842 B.n841 10.6151
R1705 B.n843 B.n842 10.6151
R1706 B.n843 B.n443 10.6151
R1707 B.n853 B.n443 10.6151
R1708 B.n854 B.n853 10.6151
R1709 B.n855 B.n854 10.6151
R1710 B.n855 B.n435 10.6151
R1711 B.n865 B.n435 10.6151
R1712 B.n866 B.n865 10.6151
R1713 B.n867 B.n866 10.6151
R1714 B.n867 B.n427 10.6151
R1715 B.n877 B.n427 10.6151
R1716 B.n878 B.n877 10.6151
R1717 B.n879 B.n878 10.6151
R1718 B.n879 B.n419 10.6151
R1719 B.n889 B.n419 10.6151
R1720 B.n890 B.n889 10.6151
R1721 B.n891 B.n890 10.6151
R1722 B.n891 B.n411 10.6151
R1723 B.n901 B.n411 10.6151
R1724 B.n902 B.n901 10.6151
R1725 B.n903 B.n902 10.6151
R1726 B.n903 B.n403 10.6151
R1727 B.n914 B.n403 10.6151
R1728 B.n915 B.n914 10.6151
R1729 B.n916 B.n915 10.6151
R1730 B.n916 B.n0 10.6151
R1731 B.n1051 B.n1 10.6151
R1732 B.n1051 B.n1050 10.6151
R1733 B.n1050 B.n1049 10.6151
R1734 B.n1049 B.n10 10.6151
R1735 B.n1043 B.n10 10.6151
R1736 B.n1043 B.n1042 10.6151
R1737 B.n1042 B.n1041 10.6151
R1738 B.n1041 B.n17 10.6151
R1739 B.n1035 B.n17 10.6151
R1740 B.n1035 B.n1034 10.6151
R1741 B.n1034 B.n1033 10.6151
R1742 B.n1033 B.n24 10.6151
R1743 B.n1027 B.n24 10.6151
R1744 B.n1027 B.n1026 10.6151
R1745 B.n1026 B.n1025 10.6151
R1746 B.n1025 B.n31 10.6151
R1747 B.n1019 B.n31 10.6151
R1748 B.n1019 B.n1018 10.6151
R1749 B.n1018 B.n1017 10.6151
R1750 B.n1017 B.n38 10.6151
R1751 B.n1011 B.n38 10.6151
R1752 B.n1011 B.n1010 10.6151
R1753 B.n1010 B.n1009 10.6151
R1754 B.n1009 B.n45 10.6151
R1755 B.n1003 B.n45 10.6151
R1756 B.n1003 B.n1002 10.6151
R1757 B.n1002 B.n1001 10.6151
R1758 B.n1001 B.n52 10.6151
R1759 B.n995 B.n52 10.6151
R1760 B.n995 B.n994 10.6151
R1761 B.n994 B.n993 10.6151
R1762 B.n993 B.n59 10.6151
R1763 B.n987 B.n59 10.6151
R1764 B.n987 B.n986 10.6151
R1765 B.n986 B.n985 10.6151
R1766 B.n985 B.n66 10.6151
R1767 B.n979 B.n66 10.6151
R1768 B.n979 B.n978 10.6151
R1769 B.n260 B.n145 9.36635
R1770 B.n283 B.n142 9.36635
R1771 B.n687 B.n686 9.36635
R1772 B.n665 B.n664 9.36635
R1773 B.n827 B.t11 7.00836
R1774 B.n991 B.t7 7.00836
R1775 B.t5 B.n421 5.1396
R1776 B.n1030 B.t4 5.1396
R1777 B.n441 B.t3 4.20521
R1778 B.t0 B.n1014 4.20521
R1779 B.n1057 B.n0 2.81026
R1780 B.n1057 B.n1 2.81026
R1781 B.n263 B.n145 1.24928
R1782 B.n280 B.n142 1.24928
R1783 B.n686 B.n685 1.24928
R1784 B.n666 B.n665 1.24928
R1785 VP.n9 VP.t5 225.816
R1786 VP.n5 VP.t4 192.274
R1787 VP.n29 VP.t1 192.274
R1788 VP.n37 VP.t2 192.274
R1789 VP.n18 VP.t0 192.274
R1790 VP.n10 VP.t3 192.274
R1791 VP.n11 VP.n8 161.3
R1792 VP.n13 VP.n12 161.3
R1793 VP.n14 VP.n7 161.3
R1794 VP.n16 VP.n15 161.3
R1795 VP.n17 VP.n6 161.3
R1796 VP.n36 VP.n0 161.3
R1797 VP.n35 VP.n34 161.3
R1798 VP.n33 VP.n1 161.3
R1799 VP.n32 VP.n31 161.3
R1800 VP.n30 VP.n2 161.3
R1801 VP.n28 VP.n27 161.3
R1802 VP.n26 VP.n3 161.3
R1803 VP.n25 VP.n24 161.3
R1804 VP.n23 VP.n4 161.3
R1805 VP.n22 VP.n21 161.3
R1806 VP.n20 VP.n5 92.6509
R1807 VP.n38 VP.n37 92.6509
R1808 VP.n19 VP.n18 92.6509
R1809 VP.n10 VP.n9 59.2423
R1810 VP.n20 VP.n19 52.2799
R1811 VP.n24 VP.n23 46.321
R1812 VP.n35 VP.n1 46.321
R1813 VP.n16 VP.n7 46.321
R1814 VP.n24 VP.n3 34.6658
R1815 VP.n31 VP.n1 34.6658
R1816 VP.n12 VP.n7 34.6658
R1817 VP.n23 VP.n22 24.4675
R1818 VP.n28 VP.n3 24.4675
R1819 VP.n31 VP.n30 24.4675
R1820 VP.n36 VP.n35 24.4675
R1821 VP.n17 VP.n16 24.4675
R1822 VP.n12 VP.n11 24.4675
R1823 VP.n22 VP.n5 18.1061
R1824 VP.n37 VP.n36 18.1061
R1825 VP.n18 VP.n17 18.1061
R1826 VP.n29 VP.n28 12.234
R1827 VP.n30 VP.n29 12.234
R1828 VP.n11 VP.n10 12.234
R1829 VP.n9 VP.n8 9.15515
R1830 VP.n19 VP.n6 0.278367
R1831 VP.n21 VP.n20 0.278367
R1832 VP.n38 VP.n0 0.278367
R1833 VP.n13 VP.n8 0.189894
R1834 VP.n14 VP.n13 0.189894
R1835 VP.n15 VP.n14 0.189894
R1836 VP.n15 VP.n6 0.189894
R1837 VP.n21 VP.n4 0.189894
R1838 VP.n25 VP.n4 0.189894
R1839 VP.n26 VP.n25 0.189894
R1840 VP.n27 VP.n26 0.189894
R1841 VP.n27 VP.n2 0.189894
R1842 VP.n32 VP.n2 0.189894
R1843 VP.n33 VP.n32 0.189894
R1844 VP.n34 VP.n33 0.189894
R1845 VP.n34 VP.n0 0.189894
R1846 VP VP.n38 0.153454
R1847 VTAIL.n410 VTAIL.n314 289.615
R1848 VTAIL.n98 VTAIL.n2 289.615
R1849 VTAIL.n308 VTAIL.n212 289.615
R1850 VTAIL.n204 VTAIL.n108 289.615
R1851 VTAIL.n346 VTAIL.n345 185
R1852 VTAIL.n351 VTAIL.n350 185
R1853 VTAIL.n353 VTAIL.n352 185
R1854 VTAIL.n342 VTAIL.n341 185
R1855 VTAIL.n359 VTAIL.n358 185
R1856 VTAIL.n361 VTAIL.n360 185
R1857 VTAIL.n338 VTAIL.n337 185
R1858 VTAIL.n367 VTAIL.n366 185
R1859 VTAIL.n369 VTAIL.n368 185
R1860 VTAIL.n334 VTAIL.n333 185
R1861 VTAIL.n375 VTAIL.n374 185
R1862 VTAIL.n377 VTAIL.n376 185
R1863 VTAIL.n330 VTAIL.n329 185
R1864 VTAIL.n383 VTAIL.n382 185
R1865 VTAIL.n385 VTAIL.n384 185
R1866 VTAIL.n326 VTAIL.n325 185
R1867 VTAIL.n392 VTAIL.n391 185
R1868 VTAIL.n393 VTAIL.n324 185
R1869 VTAIL.n395 VTAIL.n394 185
R1870 VTAIL.n322 VTAIL.n321 185
R1871 VTAIL.n401 VTAIL.n400 185
R1872 VTAIL.n403 VTAIL.n402 185
R1873 VTAIL.n318 VTAIL.n317 185
R1874 VTAIL.n409 VTAIL.n408 185
R1875 VTAIL.n411 VTAIL.n410 185
R1876 VTAIL.n34 VTAIL.n33 185
R1877 VTAIL.n39 VTAIL.n38 185
R1878 VTAIL.n41 VTAIL.n40 185
R1879 VTAIL.n30 VTAIL.n29 185
R1880 VTAIL.n47 VTAIL.n46 185
R1881 VTAIL.n49 VTAIL.n48 185
R1882 VTAIL.n26 VTAIL.n25 185
R1883 VTAIL.n55 VTAIL.n54 185
R1884 VTAIL.n57 VTAIL.n56 185
R1885 VTAIL.n22 VTAIL.n21 185
R1886 VTAIL.n63 VTAIL.n62 185
R1887 VTAIL.n65 VTAIL.n64 185
R1888 VTAIL.n18 VTAIL.n17 185
R1889 VTAIL.n71 VTAIL.n70 185
R1890 VTAIL.n73 VTAIL.n72 185
R1891 VTAIL.n14 VTAIL.n13 185
R1892 VTAIL.n80 VTAIL.n79 185
R1893 VTAIL.n81 VTAIL.n12 185
R1894 VTAIL.n83 VTAIL.n82 185
R1895 VTAIL.n10 VTAIL.n9 185
R1896 VTAIL.n89 VTAIL.n88 185
R1897 VTAIL.n91 VTAIL.n90 185
R1898 VTAIL.n6 VTAIL.n5 185
R1899 VTAIL.n97 VTAIL.n96 185
R1900 VTAIL.n99 VTAIL.n98 185
R1901 VTAIL.n309 VTAIL.n308 185
R1902 VTAIL.n307 VTAIL.n306 185
R1903 VTAIL.n216 VTAIL.n215 185
R1904 VTAIL.n301 VTAIL.n300 185
R1905 VTAIL.n299 VTAIL.n298 185
R1906 VTAIL.n220 VTAIL.n219 185
R1907 VTAIL.n293 VTAIL.n292 185
R1908 VTAIL.n291 VTAIL.n222 185
R1909 VTAIL.n290 VTAIL.n289 185
R1910 VTAIL.n225 VTAIL.n223 185
R1911 VTAIL.n284 VTAIL.n283 185
R1912 VTAIL.n282 VTAIL.n281 185
R1913 VTAIL.n229 VTAIL.n228 185
R1914 VTAIL.n276 VTAIL.n275 185
R1915 VTAIL.n274 VTAIL.n273 185
R1916 VTAIL.n233 VTAIL.n232 185
R1917 VTAIL.n268 VTAIL.n267 185
R1918 VTAIL.n266 VTAIL.n265 185
R1919 VTAIL.n237 VTAIL.n236 185
R1920 VTAIL.n260 VTAIL.n259 185
R1921 VTAIL.n258 VTAIL.n257 185
R1922 VTAIL.n241 VTAIL.n240 185
R1923 VTAIL.n252 VTAIL.n251 185
R1924 VTAIL.n250 VTAIL.n249 185
R1925 VTAIL.n245 VTAIL.n244 185
R1926 VTAIL.n205 VTAIL.n204 185
R1927 VTAIL.n203 VTAIL.n202 185
R1928 VTAIL.n112 VTAIL.n111 185
R1929 VTAIL.n197 VTAIL.n196 185
R1930 VTAIL.n195 VTAIL.n194 185
R1931 VTAIL.n116 VTAIL.n115 185
R1932 VTAIL.n189 VTAIL.n188 185
R1933 VTAIL.n187 VTAIL.n118 185
R1934 VTAIL.n186 VTAIL.n185 185
R1935 VTAIL.n121 VTAIL.n119 185
R1936 VTAIL.n180 VTAIL.n179 185
R1937 VTAIL.n178 VTAIL.n177 185
R1938 VTAIL.n125 VTAIL.n124 185
R1939 VTAIL.n172 VTAIL.n171 185
R1940 VTAIL.n170 VTAIL.n169 185
R1941 VTAIL.n129 VTAIL.n128 185
R1942 VTAIL.n164 VTAIL.n163 185
R1943 VTAIL.n162 VTAIL.n161 185
R1944 VTAIL.n133 VTAIL.n132 185
R1945 VTAIL.n156 VTAIL.n155 185
R1946 VTAIL.n154 VTAIL.n153 185
R1947 VTAIL.n137 VTAIL.n136 185
R1948 VTAIL.n148 VTAIL.n147 185
R1949 VTAIL.n146 VTAIL.n145 185
R1950 VTAIL.n141 VTAIL.n140 185
R1951 VTAIL.n347 VTAIL.t5 147.659
R1952 VTAIL.n35 VTAIL.t11 147.659
R1953 VTAIL.n246 VTAIL.t7 147.659
R1954 VTAIL.n142 VTAIL.t0 147.659
R1955 VTAIL.n351 VTAIL.n345 104.615
R1956 VTAIL.n352 VTAIL.n351 104.615
R1957 VTAIL.n352 VTAIL.n341 104.615
R1958 VTAIL.n359 VTAIL.n341 104.615
R1959 VTAIL.n360 VTAIL.n359 104.615
R1960 VTAIL.n360 VTAIL.n337 104.615
R1961 VTAIL.n367 VTAIL.n337 104.615
R1962 VTAIL.n368 VTAIL.n367 104.615
R1963 VTAIL.n368 VTAIL.n333 104.615
R1964 VTAIL.n375 VTAIL.n333 104.615
R1965 VTAIL.n376 VTAIL.n375 104.615
R1966 VTAIL.n376 VTAIL.n329 104.615
R1967 VTAIL.n383 VTAIL.n329 104.615
R1968 VTAIL.n384 VTAIL.n383 104.615
R1969 VTAIL.n384 VTAIL.n325 104.615
R1970 VTAIL.n392 VTAIL.n325 104.615
R1971 VTAIL.n393 VTAIL.n392 104.615
R1972 VTAIL.n394 VTAIL.n393 104.615
R1973 VTAIL.n394 VTAIL.n321 104.615
R1974 VTAIL.n401 VTAIL.n321 104.615
R1975 VTAIL.n402 VTAIL.n401 104.615
R1976 VTAIL.n402 VTAIL.n317 104.615
R1977 VTAIL.n409 VTAIL.n317 104.615
R1978 VTAIL.n410 VTAIL.n409 104.615
R1979 VTAIL.n39 VTAIL.n33 104.615
R1980 VTAIL.n40 VTAIL.n39 104.615
R1981 VTAIL.n40 VTAIL.n29 104.615
R1982 VTAIL.n47 VTAIL.n29 104.615
R1983 VTAIL.n48 VTAIL.n47 104.615
R1984 VTAIL.n48 VTAIL.n25 104.615
R1985 VTAIL.n55 VTAIL.n25 104.615
R1986 VTAIL.n56 VTAIL.n55 104.615
R1987 VTAIL.n56 VTAIL.n21 104.615
R1988 VTAIL.n63 VTAIL.n21 104.615
R1989 VTAIL.n64 VTAIL.n63 104.615
R1990 VTAIL.n64 VTAIL.n17 104.615
R1991 VTAIL.n71 VTAIL.n17 104.615
R1992 VTAIL.n72 VTAIL.n71 104.615
R1993 VTAIL.n72 VTAIL.n13 104.615
R1994 VTAIL.n80 VTAIL.n13 104.615
R1995 VTAIL.n81 VTAIL.n80 104.615
R1996 VTAIL.n82 VTAIL.n81 104.615
R1997 VTAIL.n82 VTAIL.n9 104.615
R1998 VTAIL.n89 VTAIL.n9 104.615
R1999 VTAIL.n90 VTAIL.n89 104.615
R2000 VTAIL.n90 VTAIL.n5 104.615
R2001 VTAIL.n97 VTAIL.n5 104.615
R2002 VTAIL.n98 VTAIL.n97 104.615
R2003 VTAIL.n308 VTAIL.n307 104.615
R2004 VTAIL.n307 VTAIL.n215 104.615
R2005 VTAIL.n300 VTAIL.n215 104.615
R2006 VTAIL.n300 VTAIL.n299 104.615
R2007 VTAIL.n299 VTAIL.n219 104.615
R2008 VTAIL.n292 VTAIL.n219 104.615
R2009 VTAIL.n292 VTAIL.n291 104.615
R2010 VTAIL.n291 VTAIL.n290 104.615
R2011 VTAIL.n290 VTAIL.n223 104.615
R2012 VTAIL.n283 VTAIL.n223 104.615
R2013 VTAIL.n283 VTAIL.n282 104.615
R2014 VTAIL.n282 VTAIL.n228 104.615
R2015 VTAIL.n275 VTAIL.n228 104.615
R2016 VTAIL.n275 VTAIL.n274 104.615
R2017 VTAIL.n274 VTAIL.n232 104.615
R2018 VTAIL.n267 VTAIL.n232 104.615
R2019 VTAIL.n267 VTAIL.n266 104.615
R2020 VTAIL.n266 VTAIL.n236 104.615
R2021 VTAIL.n259 VTAIL.n236 104.615
R2022 VTAIL.n259 VTAIL.n258 104.615
R2023 VTAIL.n258 VTAIL.n240 104.615
R2024 VTAIL.n251 VTAIL.n240 104.615
R2025 VTAIL.n251 VTAIL.n250 104.615
R2026 VTAIL.n250 VTAIL.n244 104.615
R2027 VTAIL.n204 VTAIL.n203 104.615
R2028 VTAIL.n203 VTAIL.n111 104.615
R2029 VTAIL.n196 VTAIL.n111 104.615
R2030 VTAIL.n196 VTAIL.n195 104.615
R2031 VTAIL.n195 VTAIL.n115 104.615
R2032 VTAIL.n188 VTAIL.n115 104.615
R2033 VTAIL.n188 VTAIL.n187 104.615
R2034 VTAIL.n187 VTAIL.n186 104.615
R2035 VTAIL.n186 VTAIL.n119 104.615
R2036 VTAIL.n179 VTAIL.n119 104.615
R2037 VTAIL.n179 VTAIL.n178 104.615
R2038 VTAIL.n178 VTAIL.n124 104.615
R2039 VTAIL.n171 VTAIL.n124 104.615
R2040 VTAIL.n171 VTAIL.n170 104.615
R2041 VTAIL.n170 VTAIL.n128 104.615
R2042 VTAIL.n163 VTAIL.n128 104.615
R2043 VTAIL.n163 VTAIL.n162 104.615
R2044 VTAIL.n162 VTAIL.n132 104.615
R2045 VTAIL.n155 VTAIL.n132 104.615
R2046 VTAIL.n155 VTAIL.n154 104.615
R2047 VTAIL.n154 VTAIL.n136 104.615
R2048 VTAIL.n147 VTAIL.n136 104.615
R2049 VTAIL.n147 VTAIL.n146 104.615
R2050 VTAIL.n146 VTAIL.n140 104.615
R2051 VTAIL.t5 VTAIL.n345 52.3082
R2052 VTAIL.t11 VTAIL.n33 52.3082
R2053 VTAIL.t7 VTAIL.n244 52.3082
R2054 VTAIL.t0 VTAIL.n140 52.3082
R2055 VTAIL.n211 VTAIL.n210 44.5513
R2056 VTAIL.n107 VTAIL.n106 44.5513
R2057 VTAIL.n1 VTAIL.n0 44.5511
R2058 VTAIL.n105 VTAIL.n104 44.5511
R2059 VTAIL.n415 VTAIL.n414 32.7672
R2060 VTAIL.n103 VTAIL.n102 32.7672
R2061 VTAIL.n313 VTAIL.n312 32.7672
R2062 VTAIL.n209 VTAIL.n208 32.7672
R2063 VTAIL.n107 VTAIL.n105 32.6341
R2064 VTAIL.n415 VTAIL.n313 30.3755
R2065 VTAIL.n347 VTAIL.n346 15.6677
R2066 VTAIL.n35 VTAIL.n34 15.6677
R2067 VTAIL.n246 VTAIL.n245 15.6677
R2068 VTAIL.n142 VTAIL.n141 15.6677
R2069 VTAIL.n395 VTAIL.n324 13.1884
R2070 VTAIL.n83 VTAIL.n12 13.1884
R2071 VTAIL.n293 VTAIL.n222 13.1884
R2072 VTAIL.n189 VTAIL.n118 13.1884
R2073 VTAIL.n350 VTAIL.n349 12.8005
R2074 VTAIL.n391 VTAIL.n390 12.8005
R2075 VTAIL.n396 VTAIL.n322 12.8005
R2076 VTAIL.n38 VTAIL.n37 12.8005
R2077 VTAIL.n79 VTAIL.n78 12.8005
R2078 VTAIL.n84 VTAIL.n10 12.8005
R2079 VTAIL.n294 VTAIL.n220 12.8005
R2080 VTAIL.n289 VTAIL.n224 12.8005
R2081 VTAIL.n249 VTAIL.n248 12.8005
R2082 VTAIL.n190 VTAIL.n116 12.8005
R2083 VTAIL.n185 VTAIL.n120 12.8005
R2084 VTAIL.n145 VTAIL.n144 12.8005
R2085 VTAIL.n353 VTAIL.n344 12.0247
R2086 VTAIL.n389 VTAIL.n326 12.0247
R2087 VTAIL.n400 VTAIL.n399 12.0247
R2088 VTAIL.n41 VTAIL.n32 12.0247
R2089 VTAIL.n77 VTAIL.n14 12.0247
R2090 VTAIL.n88 VTAIL.n87 12.0247
R2091 VTAIL.n298 VTAIL.n297 12.0247
R2092 VTAIL.n288 VTAIL.n225 12.0247
R2093 VTAIL.n252 VTAIL.n243 12.0247
R2094 VTAIL.n194 VTAIL.n193 12.0247
R2095 VTAIL.n184 VTAIL.n121 12.0247
R2096 VTAIL.n148 VTAIL.n139 12.0247
R2097 VTAIL.n354 VTAIL.n342 11.249
R2098 VTAIL.n386 VTAIL.n385 11.249
R2099 VTAIL.n403 VTAIL.n320 11.249
R2100 VTAIL.n42 VTAIL.n30 11.249
R2101 VTAIL.n74 VTAIL.n73 11.249
R2102 VTAIL.n91 VTAIL.n8 11.249
R2103 VTAIL.n301 VTAIL.n218 11.249
R2104 VTAIL.n285 VTAIL.n284 11.249
R2105 VTAIL.n253 VTAIL.n241 11.249
R2106 VTAIL.n197 VTAIL.n114 11.249
R2107 VTAIL.n181 VTAIL.n180 11.249
R2108 VTAIL.n149 VTAIL.n137 11.249
R2109 VTAIL.n358 VTAIL.n357 10.4732
R2110 VTAIL.n382 VTAIL.n328 10.4732
R2111 VTAIL.n404 VTAIL.n318 10.4732
R2112 VTAIL.n46 VTAIL.n45 10.4732
R2113 VTAIL.n70 VTAIL.n16 10.4732
R2114 VTAIL.n92 VTAIL.n6 10.4732
R2115 VTAIL.n302 VTAIL.n216 10.4732
R2116 VTAIL.n281 VTAIL.n227 10.4732
R2117 VTAIL.n257 VTAIL.n256 10.4732
R2118 VTAIL.n198 VTAIL.n112 10.4732
R2119 VTAIL.n177 VTAIL.n123 10.4732
R2120 VTAIL.n153 VTAIL.n152 10.4732
R2121 VTAIL.n361 VTAIL.n340 9.69747
R2122 VTAIL.n381 VTAIL.n330 9.69747
R2123 VTAIL.n408 VTAIL.n407 9.69747
R2124 VTAIL.n49 VTAIL.n28 9.69747
R2125 VTAIL.n69 VTAIL.n18 9.69747
R2126 VTAIL.n96 VTAIL.n95 9.69747
R2127 VTAIL.n306 VTAIL.n305 9.69747
R2128 VTAIL.n280 VTAIL.n229 9.69747
R2129 VTAIL.n260 VTAIL.n239 9.69747
R2130 VTAIL.n202 VTAIL.n201 9.69747
R2131 VTAIL.n176 VTAIL.n125 9.69747
R2132 VTAIL.n156 VTAIL.n135 9.69747
R2133 VTAIL.n414 VTAIL.n413 9.45567
R2134 VTAIL.n102 VTAIL.n101 9.45567
R2135 VTAIL.n312 VTAIL.n311 9.45567
R2136 VTAIL.n208 VTAIL.n207 9.45567
R2137 VTAIL.n413 VTAIL.n412 9.3005
R2138 VTAIL.n316 VTAIL.n315 9.3005
R2139 VTAIL.n407 VTAIL.n406 9.3005
R2140 VTAIL.n405 VTAIL.n404 9.3005
R2141 VTAIL.n320 VTAIL.n319 9.3005
R2142 VTAIL.n399 VTAIL.n398 9.3005
R2143 VTAIL.n397 VTAIL.n396 9.3005
R2144 VTAIL.n336 VTAIL.n335 9.3005
R2145 VTAIL.n365 VTAIL.n364 9.3005
R2146 VTAIL.n363 VTAIL.n362 9.3005
R2147 VTAIL.n340 VTAIL.n339 9.3005
R2148 VTAIL.n357 VTAIL.n356 9.3005
R2149 VTAIL.n355 VTAIL.n354 9.3005
R2150 VTAIL.n344 VTAIL.n343 9.3005
R2151 VTAIL.n349 VTAIL.n348 9.3005
R2152 VTAIL.n371 VTAIL.n370 9.3005
R2153 VTAIL.n373 VTAIL.n372 9.3005
R2154 VTAIL.n332 VTAIL.n331 9.3005
R2155 VTAIL.n379 VTAIL.n378 9.3005
R2156 VTAIL.n381 VTAIL.n380 9.3005
R2157 VTAIL.n328 VTAIL.n327 9.3005
R2158 VTAIL.n387 VTAIL.n386 9.3005
R2159 VTAIL.n389 VTAIL.n388 9.3005
R2160 VTAIL.n390 VTAIL.n323 9.3005
R2161 VTAIL.n101 VTAIL.n100 9.3005
R2162 VTAIL.n4 VTAIL.n3 9.3005
R2163 VTAIL.n95 VTAIL.n94 9.3005
R2164 VTAIL.n93 VTAIL.n92 9.3005
R2165 VTAIL.n8 VTAIL.n7 9.3005
R2166 VTAIL.n87 VTAIL.n86 9.3005
R2167 VTAIL.n85 VTAIL.n84 9.3005
R2168 VTAIL.n24 VTAIL.n23 9.3005
R2169 VTAIL.n53 VTAIL.n52 9.3005
R2170 VTAIL.n51 VTAIL.n50 9.3005
R2171 VTAIL.n28 VTAIL.n27 9.3005
R2172 VTAIL.n45 VTAIL.n44 9.3005
R2173 VTAIL.n43 VTAIL.n42 9.3005
R2174 VTAIL.n32 VTAIL.n31 9.3005
R2175 VTAIL.n37 VTAIL.n36 9.3005
R2176 VTAIL.n59 VTAIL.n58 9.3005
R2177 VTAIL.n61 VTAIL.n60 9.3005
R2178 VTAIL.n20 VTAIL.n19 9.3005
R2179 VTAIL.n67 VTAIL.n66 9.3005
R2180 VTAIL.n69 VTAIL.n68 9.3005
R2181 VTAIL.n16 VTAIL.n15 9.3005
R2182 VTAIL.n75 VTAIL.n74 9.3005
R2183 VTAIL.n77 VTAIL.n76 9.3005
R2184 VTAIL.n78 VTAIL.n11 9.3005
R2185 VTAIL.n272 VTAIL.n271 9.3005
R2186 VTAIL.n231 VTAIL.n230 9.3005
R2187 VTAIL.n278 VTAIL.n277 9.3005
R2188 VTAIL.n280 VTAIL.n279 9.3005
R2189 VTAIL.n227 VTAIL.n226 9.3005
R2190 VTAIL.n286 VTAIL.n285 9.3005
R2191 VTAIL.n288 VTAIL.n287 9.3005
R2192 VTAIL.n224 VTAIL.n221 9.3005
R2193 VTAIL.n311 VTAIL.n310 9.3005
R2194 VTAIL.n214 VTAIL.n213 9.3005
R2195 VTAIL.n305 VTAIL.n304 9.3005
R2196 VTAIL.n303 VTAIL.n302 9.3005
R2197 VTAIL.n218 VTAIL.n217 9.3005
R2198 VTAIL.n297 VTAIL.n296 9.3005
R2199 VTAIL.n295 VTAIL.n294 9.3005
R2200 VTAIL.n270 VTAIL.n269 9.3005
R2201 VTAIL.n235 VTAIL.n234 9.3005
R2202 VTAIL.n264 VTAIL.n263 9.3005
R2203 VTAIL.n262 VTAIL.n261 9.3005
R2204 VTAIL.n239 VTAIL.n238 9.3005
R2205 VTAIL.n256 VTAIL.n255 9.3005
R2206 VTAIL.n254 VTAIL.n253 9.3005
R2207 VTAIL.n243 VTAIL.n242 9.3005
R2208 VTAIL.n248 VTAIL.n247 9.3005
R2209 VTAIL.n168 VTAIL.n167 9.3005
R2210 VTAIL.n127 VTAIL.n126 9.3005
R2211 VTAIL.n174 VTAIL.n173 9.3005
R2212 VTAIL.n176 VTAIL.n175 9.3005
R2213 VTAIL.n123 VTAIL.n122 9.3005
R2214 VTAIL.n182 VTAIL.n181 9.3005
R2215 VTAIL.n184 VTAIL.n183 9.3005
R2216 VTAIL.n120 VTAIL.n117 9.3005
R2217 VTAIL.n207 VTAIL.n206 9.3005
R2218 VTAIL.n110 VTAIL.n109 9.3005
R2219 VTAIL.n201 VTAIL.n200 9.3005
R2220 VTAIL.n199 VTAIL.n198 9.3005
R2221 VTAIL.n114 VTAIL.n113 9.3005
R2222 VTAIL.n193 VTAIL.n192 9.3005
R2223 VTAIL.n191 VTAIL.n190 9.3005
R2224 VTAIL.n166 VTAIL.n165 9.3005
R2225 VTAIL.n131 VTAIL.n130 9.3005
R2226 VTAIL.n160 VTAIL.n159 9.3005
R2227 VTAIL.n158 VTAIL.n157 9.3005
R2228 VTAIL.n135 VTAIL.n134 9.3005
R2229 VTAIL.n152 VTAIL.n151 9.3005
R2230 VTAIL.n150 VTAIL.n149 9.3005
R2231 VTAIL.n139 VTAIL.n138 9.3005
R2232 VTAIL.n144 VTAIL.n143 9.3005
R2233 VTAIL.n362 VTAIL.n338 8.92171
R2234 VTAIL.n378 VTAIL.n377 8.92171
R2235 VTAIL.n411 VTAIL.n316 8.92171
R2236 VTAIL.n50 VTAIL.n26 8.92171
R2237 VTAIL.n66 VTAIL.n65 8.92171
R2238 VTAIL.n99 VTAIL.n4 8.92171
R2239 VTAIL.n309 VTAIL.n214 8.92171
R2240 VTAIL.n277 VTAIL.n276 8.92171
R2241 VTAIL.n261 VTAIL.n237 8.92171
R2242 VTAIL.n205 VTAIL.n110 8.92171
R2243 VTAIL.n173 VTAIL.n172 8.92171
R2244 VTAIL.n157 VTAIL.n133 8.92171
R2245 VTAIL.n366 VTAIL.n365 8.14595
R2246 VTAIL.n374 VTAIL.n332 8.14595
R2247 VTAIL.n412 VTAIL.n314 8.14595
R2248 VTAIL.n54 VTAIL.n53 8.14595
R2249 VTAIL.n62 VTAIL.n20 8.14595
R2250 VTAIL.n100 VTAIL.n2 8.14595
R2251 VTAIL.n310 VTAIL.n212 8.14595
R2252 VTAIL.n273 VTAIL.n231 8.14595
R2253 VTAIL.n265 VTAIL.n264 8.14595
R2254 VTAIL.n206 VTAIL.n108 8.14595
R2255 VTAIL.n169 VTAIL.n127 8.14595
R2256 VTAIL.n161 VTAIL.n160 8.14595
R2257 VTAIL.n369 VTAIL.n336 7.3702
R2258 VTAIL.n373 VTAIL.n334 7.3702
R2259 VTAIL.n57 VTAIL.n24 7.3702
R2260 VTAIL.n61 VTAIL.n22 7.3702
R2261 VTAIL.n272 VTAIL.n233 7.3702
R2262 VTAIL.n268 VTAIL.n235 7.3702
R2263 VTAIL.n168 VTAIL.n129 7.3702
R2264 VTAIL.n164 VTAIL.n131 7.3702
R2265 VTAIL.n370 VTAIL.n369 6.59444
R2266 VTAIL.n370 VTAIL.n334 6.59444
R2267 VTAIL.n58 VTAIL.n57 6.59444
R2268 VTAIL.n58 VTAIL.n22 6.59444
R2269 VTAIL.n269 VTAIL.n233 6.59444
R2270 VTAIL.n269 VTAIL.n268 6.59444
R2271 VTAIL.n165 VTAIL.n129 6.59444
R2272 VTAIL.n165 VTAIL.n164 6.59444
R2273 VTAIL.n366 VTAIL.n336 5.81868
R2274 VTAIL.n374 VTAIL.n373 5.81868
R2275 VTAIL.n414 VTAIL.n314 5.81868
R2276 VTAIL.n54 VTAIL.n24 5.81868
R2277 VTAIL.n62 VTAIL.n61 5.81868
R2278 VTAIL.n102 VTAIL.n2 5.81868
R2279 VTAIL.n312 VTAIL.n212 5.81868
R2280 VTAIL.n273 VTAIL.n272 5.81868
R2281 VTAIL.n265 VTAIL.n235 5.81868
R2282 VTAIL.n208 VTAIL.n108 5.81868
R2283 VTAIL.n169 VTAIL.n168 5.81868
R2284 VTAIL.n161 VTAIL.n131 5.81868
R2285 VTAIL.n365 VTAIL.n338 5.04292
R2286 VTAIL.n377 VTAIL.n332 5.04292
R2287 VTAIL.n412 VTAIL.n411 5.04292
R2288 VTAIL.n53 VTAIL.n26 5.04292
R2289 VTAIL.n65 VTAIL.n20 5.04292
R2290 VTAIL.n100 VTAIL.n99 5.04292
R2291 VTAIL.n310 VTAIL.n309 5.04292
R2292 VTAIL.n276 VTAIL.n231 5.04292
R2293 VTAIL.n264 VTAIL.n237 5.04292
R2294 VTAIL.n206 VTAIL.n205 5.04292
R2295 VTAIL.n172 VTAIL.n127 5.04292
R2296 VTAIL.n160 VTAIL.n133 5.04292
R2297 VTAIL.n348 VTAIL.n347 4.38563
R2298 VTAIL.n36 VTAIL.n35 4.38563
R2299 VTAIL.n247 VTAIL.n246 4.38563
R2300 VTAIL.n143 VTAIL.n142 4.38563
R2301 VTAIL.n362 VTAIL.n361 4.26717
R2302 VTAIL.n378 VTAIL.n330 4.26717
R2303 VTAIL.n408 VTAIL.n316 4.26717
R2304 VTAIL.n50 VTAIL.n49 4.26717
R2305 VTAIL.n66 VTAIL.n18 4.26717
R2306 VTAIL.n96 VTAIL.n4 4.26717
R2307 VTAIL.n306 VTAIL.n214 4.26717
R2308 VTAIL.n277 VTAIL.n229 4.26717
R2309 VTAIL.n261 VTAIL.n260 4.26717
R2310 VTAIL.n202 VTAIL.n110 4.26717
R2311 VTAIL.n173 VTAIL.n125 4.26717
R2312 VTAIL.n157 VTAIL.n156 4.26717
R2313 VTAIL.n358 VTAIL.n340 3.49141
R2314 VTAIL.n382 VTAIL.n381 3.49141
R2315 VTAIL.n407 VTAIL.n318 3.49141
R2316 VTAIL.n46 VTAIL.n28 3.49141
R2317 VTAIL.n70 VTAIL.n69 3.49141
R2318 VTAIL.n95 VTAIL.n6 3.49141
R2319 VTAIL.n305 VTAIL.n216 3.49141
R2320 VTAIL.n281 VTAIL.n280 3.49141
R2321 VTAIL.n257 VTAIL.n239 3.49141
R2322 VTAIL.n201 VTAIL.n112 3.49141
R2323 VTAIL.n177 VTAIL.n176 3.49141
R2324 VTAIL.n153 VTAIL.n135 3.49141
R2325 VTAIL.n357 VTAIL.n342 2.71565
R2326 VTAIL.n385 VTAIL.n328 2.71565
R2327 VTAIL.n404 VTAIL.n403 2.71565
R2328 VTAIL.n45 VTAIL.n30 2.71565
R2329 VTAIL.n73 VTAIL.n16 2.71565
R2330 VTAIL.n92 VTAIL.n91 2.71565
R2331 VTAIL.n302 VTAIL.n301 2.71565
R2332 VTAIL.n284 VTAIL.n227 2.71565
R2333 VTAIL.n256 VTAIL.n241 2.71565
R2334 VTAIL.n198 VTAIL.n197 2.71565
R2335 VTAIL.n180 VTAIL.n123 2.71565
R2336 VTAIL.n152 VTAIL.n137 2.71565
R2337 VTAIL.n209 VTAIL.n107 2.25912
R2338 VTAIL.n313 VTAIL.n211 2.25912
R2339 VTAIL.n105 VTAIL.n103 2.25912
R2340 VTAIL.n354 VTAIL.n353 1.93989
R2341 VTAIL.n386 VTAIL.n326 1.93989
R2342 VTAIL.n400 VTAIL.n320 1.93989
R2343 VTAIL.n42 VTAIL.n41 1.93989
R2344 VTAIL.n74 VTAIL.n14 1.93989
R2345 VTAIL.n88 VTAIL.n8 1.93989
R2346 VTAIL.n298 VTAIL.n218 1.93989
R2347 VTAIL.n285 VTAIL.n225 1.93989
R2348 VTAIL.n253 VTAIL.n252 1.93989
R2349 VTAIL.n194 VTAIL.n114 1.93989
R2350 VTAIL.n181 VTAIL.n121 1.93989
R2351 VTAIL.n149 VTAIL.n148 1.93989
R2352 VTAIL VTAIL.n415 1.63628
R2353 VTAIL.n211 VTAIL.n209 1.59964
R2354 VTAIL.n103 VTAIL.n1 1.59964
R2355 VTAIL.n350 VTAIL.n344 1.16414
R2356 VTAIL.n391 VTAIL.n389 1.16414
R2357 VTAIL.n399 VTAIL.n322 1.16414
R2358 VTAIL.n38 VTAIL.n32 1.16414
R2359 VTAIL.n79 VTAIL.n77 1.16414
R2360 VTAIL.n87 VTAIL.n10 1.16414
R2361 VTAIL.n297 VTAIL.n220 1.16414
R2362 VTAIL.n289 VTAIL.n288 1.16414
R2363 VTAIL.n249 VTAIL.n243 1.16414
R2364 VTAIL.n193 VTAIL.n116 1.16414
R2365 VTAIL.n185 VTAIL.n184 1.16414
R2366 VTAIL.n145 VTAIL.n139 1.16414
R2367 VTAIL.n0 VTAIL.t1 1.08424
R2368 VTAIL.n0 VTAIL.t3 1.08424
R2369 VTAIL.n104 VTAIL.t8 1.08424
R2370 VTAIL.n104 VTAIL.t9 1.08424
R2371 VTAIL.n210 VTAIL.t10 1.08424
R2372 VTAIL.n210 VTAIL.t6 1.08424
R2373 VTAIL.n106 VTAIL.t2 1.08424
R2374 VTAIL.n106 VTAIL.t4 1.08424
R2375 VTAIL VTAIL.n1 0.623345
R2376 VTAIL.n349 VTAIL.n346 0.388379
R2377 VTAIL.n390 VTAIL.n324 0.388379
R2378 VTAIL.n396 VTAIL.n395 0.388379
R2379 VTAIL.n37 VTAIL.n34 0.388379
R2380 VTAIL.n78 VTAIL.n12 0.388379
R2381 VTAIL.n84 VTAIL.n83 0.388379
R2382 VTAIL.n294 VTAIL.n293 0.388379
R2383 VTAIL.n224 VTAIL.n222 0.388379
R2384 VTAIL.n248 VTAIL.n245 0.388379
R2385 VTAIL.n190 VTAIL.n189 0.388379
R2386 VTAIL.n120 VTAIL.n118 0.388379
R2387 VTAIL.n144 VTAIL.n141 0.388379
R2388 VTAIL.n348 VTAIL.n343 0.155672
R2389 VTAIL.n355 VTAIL.n343 0.155672
R2390 VTAIL.n356 VTAIL.n355 0.155672
R2391 VTAIL.n356 VTAIL.n339 0.155672
R2392 VTAIL.n363 VTAIL.n339 0.155672
R2393 VTAIL.n364 VTAIL.n363 0.155672
R2394 VTAIL.n364 VTAIL.n335 0.155672
R2395 VTAIL.n371 VTAIL.n335 0.155672
R2396 VTAIL.n372 VTAIL.n371 0.155672
R2397 VTAIL.n372 VTAIL.n331 0.155672
R2398 VTAIL.n379 VTAIL.n331 0.155672
R2399 VTAIL.n380 VTAIL.n379 0.155672
R2400 VTAIL.n380 VTAIL.n327 0.155672
R2401 VTAIL.n387 VTAIL.n327 0.155672
R2402 VTAIL.n388 VTAIL.n387 0.155672
R2403 VTAIL.n388 VTAIL.n323 0.155672
R2404 VTAIL.n397 VTAIL.n323 0.155672
R2405 VTAIL.n398 VTAIL.n397 0.155672
R2406 VTAIL.n398 VTAIL.n319 0.155672
R2407 VTAIL.n405 VTAIL.n319 0.155672
R2408 VTAIL.n406 VTAIL.n405 0.155672
R2409 VTAIL.n406 VTAIL.n315 0.155672
R2410 VTAIL.n413 VTAIL.n315 0.155672
R2411 VTAIL.n36 VTAIL.n31 0.155672
R2412 VTAIL.n43 VTAIL.n31 0.155672
R2413 VTAIL.n44 VTAIL.n43 0.155672
R2414 VTAIL.n44 VTAIL.n27 0.155672
R2415 VTAIL.n51 VTAIL.n27 0.155672
R2416 VTAIL.n52 VTAIL.n51 0.155672
R2417 VTAIL.n52 VTAIL.n23 0.155672
R2418 VTAIL.n59 VTAIL.n23 0.155672
R2419 VTAIL.n60 VTAIL.n59 0.155672
R2420 VTAIL.n60 VTAIL.n19 0.155672
R2421 VTAIL.n67 VTAIL.n19 0.155672
R2422 VTAIL.n68 VTAIL.n67 0.155672
R2423 VTAIL.n68 VTAIL.n15 0.155672
R2424 VTAIL.n75 VTAIL.n15 0.155672
R2425 VTAIL.n76 VTAIL.n75 0.155672
R2426 VTAIL.n76 VTAIL.n11 0.155672
R2427 VTAIL.n85 VTAIL.n11 0.155672
R2428 VTAIL.n86 VTAIL.n85 0.155672
R2429 VTAIL.n86 VTAIL.n7 0.155672
R2430 VTAIL.n93 VTAIL.n7 0.155672
R2431 VTAIL.n94 VTAIL.n93 0.155672
R2432 VTAIL.n94 VTAIL.n3 0.155672
R2433 VTAIL.n101 VTAIL.n3 0.155672
R2434 VTAIL.n311 VTAIL.n213 0.155672
R2435 VTAIL.n304 VTAIL.n213 0.155672
R2436 VTAIL.n304 VTAIL.n303 0.155672
R2437 VTAIL.n303 VTAIL.n217 0.155672
R2438 VTAIL.n296 VTAIL.n217 0.155672
R2439 VTAIL.n296 VTAIL.n295 0.155672
R2440 VTAIL.n295 VTAIL.n221 0.155672
R2441 VTAIL.n287 VTAIL.n221 0.155672
R2442 VTAIL.n287 VTAIL.n286 0.155672
R2443 VTAIL.n286 VTAIL.n226 0.155672
R2444 VTAIL.n279 VTAIL.n226 0.155672
R2445 VTAIL.n279 VTAIL.n278 0.155672
R2446 VTAIL.n278 VTAIL.n230 0.155672
R2447 VTAIL.n271 VTAIL.n230 0.155672
R2448 VTAIL.n271 VTAIL.n270 0.155672
R2449 VTAIL.n270 VTAIL.n234 0.155672
R2450 VTAIL.n263 VTAIL.n234 0.155672
R2451 VTAIL.n263 VTAIL.n262 0.155672
R2452 VTAIL.n262 VTAIL.n238 0.155672
R2453 VTAIL.n255 VTAIL.n238 0.155672
R2454 VTAIL.n255 VTAIL.n254 0.155672
R2455 VTAIL.n254 VTAIL.n242 0.155672
R2456 VTAIL.n247 VTAIL.n242 0.155672
R2457 VTAIL.n207 VTAIL.n109 0.155672
R2458 VTAIL.n200 VTAIL.n109 0.155672
R2459 VTAIL.n200 VTAIL.n199 0.155672
R2460 VTAIL.n199 VTAIL.n113 0.155672
R2461 VTAIL.n192 VTAIL.n113 0.155672
R2462 VTAIL.n192 VTAIL.n191 0.155672
R2463 VTAIL.n191 VTAIL.n117 0.155672
R2464 VTAIL.n183 VTAIL.n117 0.155672
R2465 VTAIL.n183 VTAIL.n182 0.155672
R2466 VTAIL.n182 VTAIL.n122 0.155672
R2467 VTAIL.n175 VTAIL.n122 0.155672
R2468 VTAIL.n175 VTAIL.n174 0.155672
R2469 VTAIL.n174 VTAIL.n126 0.155672
R2470 VTAIL.n167 VTAIL.n126 0.155672
R2471 VTAIL.n167 VTAIL.n166 0.155672
R2472 VTAIL.n166 VTAIL.n130 0.155672
R2473 VTAIL.n159 VTAIL.n130 0.155672
R2474 VTAIL.n159 VTAIL.n158 0.155672
R2475 VTAIL.n158 VTAIL.n134 0.155672
R2476 VTAIL.n151 VTAIL.n134 0.155672
R2477 VTAIL.n151 VTAIL.n150 0.155672
R2478 VTAIL.n150 VTAIL.n138 0.155672
R2479 VTAIL.n143 VTAIL.n138 0.155672
R2480 VDD1.n96 VDD1.n0 289.615
R2481 VDD1.n197 VDD1.n101 289.615
R2482 VDD1.n97 VDD1.n96 185
R2483 VDD1.n95 VDD1.n94 185
R2484 VDD1.n4 VDD1.n3 185
R2485 VDD1.n89 VDD1.n88 185
R2486 VDD1.n87 VDD1.n86 185
R2487 VDD1.n8 VDD1.n7 185
R2488 VDD1.n81 VDD1.n80 185
R2489 VDD1.n79 VDD1.n10 185
R2490 VDD1.n78 VDD1.n77 185
R2491 VDD1.n13 VDD1.n11 185
R2492 VDD1.n72 VDD1.n71 185
R2493 VDD1.n70 VDD1.n69 185
R2494 VDD1.n17 VDD1.n16 185
R2495 VDD1.n64 VDD1.n63 185
R2496 VDD1.n62 VDD1.n61 185
R2497 VDD1.n21 VDD1.n20 185
R2498 VDD1.n56 VDD1.n55 185
R2499 VDD1.n54 VDD1.n53 185
R2500 VDD1.n25 VDD1.n24 185
R2501 VDD1.n48 VDD1.n47 185
R2502 VDD1.n46 VDD1.n45 185
R2503 VDD1.n29 VDD1.n28 185
R2504 VDD1.n40 VDD1.n39 185
R2505 VDD1.n38 VDD1.n37 185
R2506 VDD1.n33 VDD1.n32 185
R2507 VDD1.n133 VDD1.n132 185
R2508 VDD1.n138 VDD1.n137 185
R2509 VDD1.n140 VDD1.n139 185
R2510 VDD1.n129 VDD1.n128 185
R2511 VDD1.n146 VDD1.n145 185
R2512 VDD1.n148 VDD1.n147 185
R2513 VDD1.n125 VDD1.n124 185
R2514 VDD1.n154 VDD1.n153 185
R2515 VDD1.n156 VDD1.n155 185
R2516 VDD1.n121 VDD1.n120 185
R2517 VDD1.n162 VDD1.n161 185
R2518 VDD1.n164 VDD1.n163 185
R2519 VDD1.n117 VDD1.n116 185
R2520 VDD1.n170 VDD1.n169 185
R2521 VDD1.n172 VDD1.n171 185
R2522 VDD1.n113 VDD1.n112 185
R2523 VDD1.n179 VDD1.n178 185
R2524 VDD1.n180 VDD1.n111 185
R2525 VDD1.n182 VDD1.n181 185
R2526 VDD1.n109 VDD1.n108 185
R2527 VDD1.n188 VDD1.n187 185
R2528 VDD1.n190 VDD1.n189 185
R2529 VDD1.n105 VDD1.n104 185
R2530 VDD1.n196 VDD1.n195 185
R2531 VDD1.n198 VDD1.n197 185
R2532 VDD1.n34 VDD1.t0 147.659
R2533 VDD1.n134 VDD1.t1 147.659
R2534 VDD1.n96 VDD1.n95 104.615
R2535 VDD1.n95 VDD1.n3 104.615
R2536 VDD1.n88 VDD1.n3 104.615
R2537 VDD1.n88 VDD1.n87 104.615
R2538 VDD1.n87 VDD1.n7 104.615
R2539 VDD1.n80 VDD1.n7 104.615
R2540 VDD1.n80 VDD1.n79 104.615
R2541 VDD1.n79 VDD1.n78 104.615
R2542 VDD1.n78 VDD1.n11 104.615
R2543 VDD1.n71 VDD1.n11 104.615
R2544 VDD1.n71 VDD1.n70 104.615
R2545 VDD1.n70 VDD1.n16 104.615
R2546 VDD1.n63 VDD1.n16 104.615
R2547 VDD1.n63 VDD1.n62 104.615
R2548 VDD1.n62 VDD1.n20 104.615
R2549 VDD1.n55 VDD1.n20 104.615
R2550 VDD1.n55 VDD1.n54 104.615
R2551 VDD1.n54 VDD1.n24 104.615
R2552 VDD1.n47 VDD1.n24 104.615
R2553 VDD1.n47 VDD1.n46 104.615
R2554 VDD1.n46 VDD1.n28 104.615
R2555 VDD1.n39 VDD1.n28 104.615
R2556 VDD1.n39 VDD1.n38 104.615
R2557 VDD1.n38 VDD1.n32 104.615
R2558 VDD1.n138 VDD1.n132 104.615
R2559 VDD1.n139 VDD1.n138 104.615
R2560 VDD1.n139 VDD1.n128 104.615
R2561 VDD1.n146 VDD1.n128 104.615
R2562 VDD1.n147 VDD1.n146 104.615
R2563 VDD1.n147 VDD1.n124 104.615
R2564 VDD1.n154 VDD1.n124 104.615
R2565 VDD1.n155 VDD1.n154 104.615
R2566 VDD1.n155 VDD1.n120 104.615
R2567 VDD1.n162 VDD1.n120 104.615
R2568 VDD1.n163 VDD1.n162 104.615
R2569 VDD1.n163 VDD1.n116 104.615
R2570 VDD1.n170 VDD1.n116 104.615
R2571 VDD1.n171 VDD1.n170 104.615
R2572 VDD1.n171 VDD1.n112 104.615
R2573 VDD1.n179 VDD1.n112 104.615
R2574 VDD1.n180 VDD1.n179 104.615
R2575 VDD1.n181 VDD1.n180 104.615
R2576 VDD1.n181 VDD1.n108 104.615
R2577 VDD1.n188 VDD1.n108 104.615
R2578 VDD1.n189 VDD1.n188 104.615
R2579 VDD1.n189 VDD1.n104 104.615
R2580 VDD1.n196 VDD1.n104 104.615
R2581 VDD1.n197 VDD1.n196 104.615
R2582 VDD1.n203 VDD1.n202 61.7392
R2583 VDD1.n205 VDD1.n204 61.2299
R2584 VDD1.t0 VDD1.n32 52.3082
R2585 VDD1.t1 VDD1.n132 52.3082
R2586 VDD1 VDD1.n100 51.1981
R2587 VDD1.n203 VDD1.n201 51.0846
R2588 VDD1.n205 VDD1.n203 48.5181
R2589 VDD1.n34 VDD1.n33 15.6677
R2590 VDD1.n134 VDD1.n133 15.6677
R2591 VDD1.n81 VDD1.n10 13.1884
R2592 VDD1.n182 VDD1.n111 13.1884
R2593 VDD1.n82 VDD1.n8 12.8005
R2594 VDD1.n77 VDD1.n12 12.8005
R2595 VDD1.n37 VDD1.n36 12.8005
R2596 VDD1.n137 VDD1.n136 12.8005
R2597 VDD1.n178 VDD1.n177 12.8005
R2598 VDD1.n183 VDD1.n109 12.8005
R2599 VDD1.n86 VDD1.n85 12.0247
R2600 VDD1.n76 VDD1.n13 12.0247
R2601 VDD1.n40 VDD1.n31 12.0247
R2602 VDD1.n140 VDD1.n131 12.0247
R2603 VDD1.n176 VDD1.n113 12.0247
R2604 VDD1.n187 VDD1.n186 12.0247
R2605 VDD1.n89 VDD1.n6 11.249
R2606 VDD1.n73 VDD1.n72 11.249
R2607 VDD1.n41 VDD1.n29 11.249
R2608 VDD1.n141 VDD1.n129 11.249
R2609 VDD1.n173 VDD1.n172 11.249
R2610 VDD1.n190 VDD1.n107 11.249
R2611 VDD1.n90 VDD1.n4 10.4732
R2612 VDD1.n69 VDD1.n15 10.4732
R2613 VDD1.n45 VDD1.n44 10.4732
R2614 VDD1.n145 VDD1.n144 10.4732
R2615 VDD1.n169 VDD1.n115 10.4732
R2616 VDD1.n191 VDD1.n105 10.4732
R2617 VDD1.n94 VDD1.n93 9.69747
R2618 VDD1.n68 VDD1.n17 9.69747
R2619 VDD1.n48 VDD1.n27 9.69747
R2620 VDD1.n148 VDD1.n127 9.69747
R2621 VDD1.n168 VDD1.n117 9.69747
R2622 VDD1.n195 VDD1.n194 9.69747
R2623 VDD1.n100 VDD1.n99 9.45567
R2624 VDD1.n201 VDD1.n200 9.45567
R2625 VDD1.n60 VDD1.n59 9.3005
R2626 VDD1.n19 VDD1.n18 9.3005
R2627 VDD1.n66 VDD1.n65 9.3005
R2628 VDD1.n68 VDD1.n67 9.3005
R2629 VDD1.n15 VDD1.n14 9.3005
R2630 VDD1.n74 VDD1.n73 9.3005
R2631 VDD1.n76 VDD1.n75 9.3005
R2632 VDD1.n12 VDD1.n9 9.3005
R2633 VDD1.n99 VDD1.n98 9.3005
R2634 VDD1.n2 VDD1.n1 9.3005
R2635 VDD1.n93 VDD1.n92 9.3005
R2636 VDD1.n91 VDD1.n90 9.3005
R2637 VDD1.n6 VDD1.n5 9.3005
R2638 VDD1.n85 VDD1.n84 9.3005
R2639 VDD1.n83 VDD1.n82 9.3005
R2640 VDD1.n58 VDD1.n57 9.3005
R2641 VDD1.n23 VDD1.n22 9.3005
R2642 VDD1.n52 VDD1.n51 9.3005
R2643 VDD1.n50 VDD1.n49 9.3005
R2644 VDD1.n27 VDD1.n26 9.3005
R2645 VDD1.n44 VDD1.n43 9.3005
R2646 VDD1.n42 VDD1.n41 9.3005
R2647 VDD1.n31 VDD1.n30 9.3005
R2648 VDD1.n36 VDD1.n35 9.3005
R2649 VDD1.n200 VDD1.n199 9.3005
R2650 VDD1.n103 VDD1.n102 9.3005
R2651 VDD1.n194 VDD1.n193 9.3005
R2652 VDD1.n192 VDD1.n191 9.3005
R2653 VDD1.n107 VDD1.n106 9.3005
R2654 VDD1.n186 VDD1.n185 9.3005
R2655 VDD1.n184 VDD1.n183 9.3005
R2656 VDD1.n123 VDD1.n122 9.3005
R2657 VDD1.n152 VDD1.n151 9.3005
R2658 VDD1.n150 VDD1.n149 9.3005
R2659 VDD1.n127 VDD1.n126 9.3005
R2660 VDD1.n144 VDD1.n143 9.3005
R2661 VDD1.n142 VDD1.n141 9.3005
R2662 VDD1.n131 VDD1.n130 9.3005
R2663 VDD1.n136 VDD1.n135 9.3005
R2664 VDD1.n158 VDD1.n157 9.3005
R2665 VDD1.n160 VDD1.n159 9.3005
R2666 VDD1.n119 VDD1.n118 9.3005
R2667 VDD1.n166 VDD1.n165 9.3005
R2668 VDD1.n168 VDD1.n167 9.3005
R2669 VDD1.n115 VDD1.n114 9.3005
R2670 VDD1.n174 VDD1.n173 9.3005
R2671 VDD1.n176 VDD1.n175 9.3005
R2672 VDD1.n177 VDD1.n110 9.3005
R2673 VDD1.n97 VDD1.n2 8.92171
R2674 VDD1.n65 VDD1.n64 8.92171
R2675 VDD1.n49 VDD1.n25 8.92171
R2676 VDD1.n149 VDD1.n125 8.92171
R2677 VDD1.n165 VDD1.n164 8.92171
R2678 VDD1.n198 VDD1.n103 8.92171
R2679 VDD1.n98 VDD1.n0 8.14595
R2680 VDD1.n61 VDD1.n19 8.14595
R2681 VDD1.n53 VDD1.n52 8.14595
R2682 VDD1.n153 VDD1.n152 8.14595
R2683 VDD1.n161 VDD1.n119 8.14595
R2684 VDD1.n199 VDD1.n101 8.14595
R2685 VDD1.n60 VDD1.n21 7.3702
R2686 VDD1.n56 VDD1.n23 7.3702
R2687 VDD1.n156 VDD1.n123 7.3702
R2688 VDD1.n160 VDD1.n121 7.3702
R2689 VDD1.n57 VDD1.n21 6.59444
R2690 VDD1.n57 VDD1.n56 6.59444
R2691 VDD1.n157 VDD1.n156 6.59444
R2692 VDD1.n157 VDD1.n121 6.59444
R2693 VDD1.n100 VDD1.n0 5.81868
R2694 VDD1.n61 VDD1.n60 5.81868
R2695 VDD1.n53 VDD1.n23 5.81868
R2696 VDD1.n153 VDD1.n123 5.81868
R2697 VDD1.n161 VDD1.n160 5.81868
R2698 VDD1.n201 VDD1.n101 5.81868
R2699 VDD1.n98 VDD1.n97 5.04292
R2700 VDD1.n64 VDD1.n19 5.04292
R2701 VDD1.n52 VDD1.n25 5.04292
R2702 VDD1.n152 VDD1.n125 5.04292
R2703 VDD1.n164 VDD1.n119 5.04292
R2704 VDD1.n199 VDD1.n198 5.04292
R2705 VDD1.n35 VDD1.n34 4.38563
R2706 VDD1.n135 VDD1.n134 4.38563
R2707 VDD1.n94 VDD1.n2 4.26717
R2708 VDD1.n65 VDD1.n17 4.26717
R2709 VDD1.n49 VDD1.n48 4.26717
R2710 VDD1.n149 VDD1.n148 4.26717
R2711 VDD1.n165 VDD1.n117 4.26717
R2712 VDD1.n195 VDD1.n103 4.26717
R2713 VDD1.n93 VDD1.n4 3.49141
R2714 VDD1.n69 VDD1.n68 3.49141
R2715 VDD1.n45 VDD1.n27 3.49141
R2716 VDD1.n145 VDD1.n127 3.49141
R2717 VDD1.n169 VDD1.n168 3.49141
R2718 VDD1.n194 VDD1.n105 3.49141
R2719 VDD1.n90 VDD1.n89 2.71565
R2720 VDD1.n72 VDD1.n15 2.71565
R2721 VDD1.n44 VDD1.n29 2.71565
R2722 VDD1.n144 VDD1.n129 2.71565
R2723 VDD1.n172 VDD1.n115 2.71565
R2724 VDD1.n191 VDD1.n190 2.71565
R2725 VDD1.n86 VDD1.n6 1.93989
R2726 VDD1.n73 VDD1.n13 1.93989
R2727 VDD1.n41 VDD1.n40 1.93989
R2728 VDD1.n141 VDD1.n140 1.93989
R2729 VDD1.n173 VDD1.n113 1.93989
R2730 VDD1.n187 VDD1.n107 1.93989
R2731 VDD1.n85 VDD1.n8 1.16414
R2732 VDD1.n77 VDD1.n76 1.16414
R2733 VDD1.n37 VDD1.n31 1.16414
R2734 VDD1.n137 VDD1.n131 1.16414
R2735 VDD1.n178 VDD1.n176 1.16414
R2736 VDD1.n186 VDD1.n109 1.16414
R2737 VDD1.n204 VDD1.t2 1.08424
R2738 VDD1.n204 VDD1.t5 1.08424
R2739 VDD1.n202 VDD1.t4 1.08424
R2740 VDD1.n202 VDD1.t3 1.08424
R2741 VDD1 VDD1.n205 0.506965
R2742 VDD1.n82 VDD1.n81 0.388379
R2743 VDD1.n12 VDD1.n10 0.388379
R2744 VDD1.n36 VDD1.n33 0.388379
R2745 VDD1.n136 VDD1.n133 0.388379
R2746 VDD1.n177 VDD1.n111 0.388379
R2747 VDD1.n183 VDD1.n182 0.388379
R2748 VDD1.n99 VDD1.n1 0.155672
R2749 VDD1.n92 VDD1.n1 0.155672
R2750 VDD1.n92 VDD1.n91 0.155672
R2751 VDD1.n91 VDD1.n5 0.155672
R2752 VDD1.n84 VDD1.n5 0.155672
R2753 VDD1.n84 VDD1.n83 0.155672
R2754 VDD1.n83 VDD1.n9 0.155672
R2755 VDD1.n75 VDD1.n9 0.155672
R2756 VDD1.n75 VDD1.n74 0.155672
R2757 VDD1.n74 VDD1.n14 0.155672
R2758 VDD1.n67 VDD1.n14 0.155672
R2759 VDD1.n67 VDD1.n66 0.155672
R2760 VDD1.n66 VDD1.n18 0.155672
R2761 VDD1.n59 VDD1.n18 0.155672
R2762 VDD1.n59 VDD1.n58 0.155672
R2763 VDD1.n58 VDD1.n22 0.155672
R2764 VDD1.n51 VDD1.n22 0.155672
R2765 VDD1.n51 VDD1.n50 0.155672
R2766 VDD1.n50 VDD1.n26 0.155672
R2767 VDD1.n43 VDD1.n26 0.155672
R2768 VDD1.n43 VDD1.n42 0.155672
R2769 VDD1.n42 VDD1.n30 0.155672
R2770 VDD1.n35 VDD1.n30 0.155672
R2771 VDD1.n135 VDD1.n130 0.155672
R2772 VDD1.n142 VDD1.n130 0.155672
R2773 VDD1.n143 VDD1.n142 0.155672
R2774 VDD1.n143 VDD1.n126 0.155672
R2775 VDD1.n150 VDD1.n126 0.155672
R2776 VDD1.n151 VDD1.n150 0.155672
R2777 VDD1.n151 VDD1.n122 0.155672
R2778 VDD1.n158 VDD1.n122 0.155672
R2779 VDD1.n159 VDD1.n158 0.155672
R2780 VDD1.n159 VDD1.n118 0.155672
R2781 VDD1.n166 VDD1.n118 0.155672
R2782 VDD1.n167 VDD1.n166 0.155672
R2783 VDD1.n167 VDD1.n114 0.155672
R2784 VDD1.n174 VDD1.n114 0.155672
R2785 VDD1.n175 VDD1.n174 0.155672
R2786 VDD1.n175 VDD1.n110 0.155672
R2787 VDD1.n184 VDD1.n110 0.155672
R2788 VDD1.n185 VDD1.n184 0.155672
R2789 VDD1.n185 VDD1.n106 0.155672
R2790 VDD1.n192 VDD1.n106 0.155672
R2791 VDD1.n193 VDD1.n192 0.155672
R2792 VDD1.n193 VDD1.n102 0.155672
R2793 VDD1.n200 VDD1.n102 0.155672
R2794 VN.n3 VN.t4 225.816
R2795 VN.n17 VN.t5 225.816
R2796 VN.n4 VN.t3 192.274
R2797 VN.n12 VN.t1 192.274
R2798 VN.n18 VN.t2 192.274
R2799 VN.n26 VN.t0 192.274
R2800 VN.n25 VN.n14 161.3
R2801 VN.n24 VN.n23 161.3
R2802 VN.n22 VN.n15 161.3
R2803 VN.n21 VN.n20 161.3
R2804 VN.n19 VN.n16 161.3
R2805 VN.n11 VN.n0 161.3
R2806 VN.n10 VN.n9 161.3
R2807 VN.n8 VN.n1 161.3
R2808 VN.n7 VN.n6 161.3
R2809 VN.n5 VN.n2 161.3
R2810 VN.n13 VN.n12 92.6509
R2811 VN.n27 VN.n26 92.6509
R2812 VN.n4 VN.n3 59.2423
R2813 VN.n18 VN.n17 59.2423
R2814 VN VN.n27 52.5588
R2815 VN.n10 VN.n1 46.321
R2816 VN.n24 VN.n15 46.321
R2817 VN.n6 VN.n1 34.6658
R2818 VN.n20 VN.n15 34.6658
R2819 VN.n6 VN.n5 24.4675
R2820 VN.n11 VN.n10 24.4675
R2821 VN.n20 VN.n19 24.4675
R2822 VN.n25 VN.n24 24.4675
R2823 VN.n12 VN.n11 18.1061
R2824 VN.n26 VN.n25 18.1061
R2825 VN.n5 VN.n4 12.234
R2826 VN.n19 VN.n18 12.234
R2827 VN.n17 VN.n16 9.15515
R2828 VN.n3 VN.n2 9.15515
R2829 VN.n27 VN.n14 0.278367
R2830 VN.n13 VN.n0 0.278367
R2831 VN.n23 VN.n14 0.189894
R2832 VN.n23 VN.n22 0.189894
R2833 VN.n22 VN.n21 0.189894
R2834 VN.n21 VN.n16 0.189894
R2835 VN.n7 VN.n2 0.189894
R2836 VN.n8 VN.n7 0.189894
R2837 VN.n9 VN.n8 0.189894
R2838 VN.n9 VN.n0 0.189894
R2839 VN VN.n13 0.153454
R2840 VDD2.n199 VDD2.n103 289.615
R2841 VDD2.n96 VDD2.n0 289.615
R2842 VDD2.n200 VDD2.n199 185
R2843 VDD2.n198 VDD2.n197 185
R2844 VDD2.n107 VDD2.n106 185
R2845 VDD2.n192 VDD2.n191 185
R2846 VDD2.n190 VDD2.n189 185
R2847 VDD2.n111 VDD2.n110 185
R2848 VDD2.n184 VDD2.n183 185
R2849 VDD2.n182 VDD2.n113 185
R2850 VDD2.n181 VDD2.n180 185
R2851 VDD2.n116 VDD2.n114 185
R2852 VDD2.n175 VDD2.n174 185
R2853 VDD2.n173 VDD2.n172 185
R2854 VDD2.n120 VDD2.n119 185
R2855 VDD2.n167 VDD2.n166 185
R2856 VDD2.n165 VDD2.n164 185
R2857 VDD2.n124 VDD2.n123 185
R2858 VDD2.n159 VDD2.n158 185
R2859 VDD2.n157 VDD2.n156 185
R2860 VDD2.n128 VDD2.n127 185
R2861 VDD2.n151 VDD2.n150 185
R2862 VDD2.n149 VDD2.n148 185
R2863 VDD2.n132 VDD2.n131 185
R2864 VDD2.n143 VDD2.n142 185
R2865 VDD2.n141 VDD2.n140 185
R2866 VDD2.n136 VDD2.n135 185
R2867 VDD2.n32 VDD2.n31 185
R2868 VDD2.n37 VDD2.n36 185
R2869 VDD2.n39 VDD2.n38 185
R2870 VDD2.n28 VDD2.n27 185
R2871 VDD2.n45 VDD2.n44 185
R2872 VDD2.n47 VDD2.n46 185
R2873 VDD2.n24 VDD2.n23 185
R2874 VDD2.n53 VDD2.n52 185
R2875 VDD2.n55 VDD2.n54 185
R2876 VDD2.n20 VDD2.n19 185
R2877 VDD2.n61 VDD2.n60 185
R2878 VDD2.n63 VDD2.n62 185
R2879 VDD2.n16 VDD2.n15 185
R2880 VDD2.n69 VDD2.n68 185
R2881 VDD2.n71 VDD2.n70 185
R2882 VDD2.n12 VDD2.n11 185
R2883 VDD2.n78 VDD2.n77 185
R2884 VDD2.n79 VDD2.n10 185
R2885 VDD2.n81 VDD2.n80 185
R2886 VDD2.n8 VDD2.n7 185
R2887 VDD2.n87 VDD2.n86 185
R2888 VDD2.n89 VDD2.n88 185
R2889 VDD2.n4 VDD2.n3 185
R2890 VDD2.n95 VDD2.n94 185
R2891 VDD2.n97 VDD2.n96 185
R2892 VDD2.n137 VDD2.t5 147.659
R2893 VDD2.n33 VDD2.t1 147.659
R2894 VDD2.n199 VDD2.n198 104.615
R2895 VDD2.n198 VDD2.n106 104.615
R2896 VDD2.n191 VDD2.n106 104.615
R2897 VDD2.n191 VDD2.n190 104.615
R2898 VDD2.n190 VDD2.n110 104.615
R2899 VDD2.n183 VDD2.n110 104.615
R2900 VDD2.n183 VDD2.n182 104.615
R2901 VDD2.n182 VDD2.n181 104.615
R2902 VDD2.n181 VDD2.n114 104.615
R2903 VDD2.n174 VDD2.n114 104.615
R2904 VDD2.n174 VDD2.n173 104.615
R2905 VDD2.n173 VDD2.n119 104.615
R2906 VDD2.n166 VDD2.n119 104.615
R2907 VDD2.n166 VDD2.n165 104.615
R2908 VDD2.n165 VDD2.n123 104.615
R2909 VDD2.n158 VDD2.n123 104.615
R2910 VDD2.n158 VDD2.n157 104.615
R2911 VDD2.n157 VDD2.n127 104.615
R2912 VDD2.n150 VDD2.n127 104.615
R2913 VDD2.n150 VDD2.n149 104.615
R2914 VDD2.n149 VDD2.n131 104.615
R2915 VDD2.n142 VDD2.n131 104.615
R2916 VDD2.n142 VDD2.n141 104.615
R2917 VDD2.n141 VDD2.n135 104.615
R2918 VDD2.n37 VDD2.n31 104.615
R2919 VDD2.n38 VDD2.n37 104.615
R2920 VDD2.n38 VDD2.n27 104.615
R2921 VDD2.n45 VDD2.n27 104.615
R2922 VDD2.n46 VDD2.n45 104.615
R2923 VDD2.n46 VDD2.n23 104.615
R2924 VDD2.n53 VDD2.n23 104.615
R2925 VDD2.n54 VDD2.n53 104.615
R2926 VDD2.n54 VDD2.n19 104.615
R2927 VDD2.n61 VDD2.n19 104.615
R2928 VDD2.n62 VDD2.n61 104.615
R2929 VDD2.n62 VDD2.n15 104.615
R2930 VDD2.n69 VDD2.n15 104.615
R2931 VDD2.n70 VDD2.n69 104.615
R2932 VDD2.n70 VDD2.n11 104.615
R2933 VDD2.n78 VDD2.n11 104.615
R2934 VDD2.n79 VDD2.n78 104.615
R2935 VDD2.n80 VDD2.n79 104.615
R2936 VDD2.n80 VDD2.n7 104.615
R2937 VDD2.n87 VDD2.n7 104.615
R2938 VDD2.n88 VDD2.n87 104.615
R2939 VDD2.n88 VDD2.n3 104.615
R2940 VDD2.n95 VDD2.n3 104.615
R2941 VDD2.n96 VDD2.n95 104.615
R2942 VDD2.n102 VDD2.n101 61.7392
R2943 VDD2 VDD2.n205 61.7364
R2944 VDD2.t5 VDD2.n135 52.3082
R2945 VDD2.t1 VDD2.n31 52.3082
R2946 VDD2.n102 VDD2.n100 51.0846
R2947 VDD2.n204 VDD2.n203 49.446
R2948 VDD2.n204 VDD2.n102 46.8058
R2949 VDD2.n137 VDD2.n136 15.6677
R2950 VDD2.n33 VDD2.n32 15.6677
R2951 VDD2.n184 VDD2.n113 13.1884
R2952 VDD2.n81 VDD2.n10 13.1884
R2953 VDD2.n185 VDD2.n111 12.8005
R2954 VDD2.n180 VDD2.n115 12.8005
R2955 VDD2.n140 VDD2.n139 12.8005
R2956 VDD2.n36 VDD2.n35 12.8005
R2957 VDD2.n77 VDD2.n76 12.8005
R2958 VDD2.n82 VDD2.n8 12.8005
R2959 VDD2.n189 VDD2.n188 12.0247
R2960 VDD2.n179 VDD2.n116 12.0247
R2961 VDD2.n143 VDD2.n134 12.0247
R2962 VDD2.n39 VDD2.n30 12.0247
R2963 VDD2.n75 VDD2.n12 12.0247
R2964 VDD2.n86 VDD2.n85 12.0247
R2965 VDD2.n192 VDD2.n109 11.249
R2966 VDD2.n176 VDD2.n175 11.249
R2967 VDD2.n144 VDD2.n132 11.249
R2968 VDD2.n40 VDD2.n28 11.249
R2969 VDD2.n72 VDD2.n71 11.249
R2970 VDD2.n89 VDD2.n6 11.249
R2971 VDD2.n193 VDD2.n107 10.4732
R2972 VDD2.n172 VDD2.n118 10.4732
R2973 VDD2.n148 VDD2.n147 10.4732
R2974 VDD2.n44 VDD2.n43 10.4732
R2975 VDD2.n68 VDD2.n14 10.4732
R2976 VDD2.n90 VDD2.n4 10.4732
R2977 VDD2.n197 VDD2.n196 9.69747
R2978 VDD2.n171 VDD2.n120 9.69747
R2979 VDD2.n151 VDD2.n130 9.69747
R2980 VDD2.n47 VDD2.n26 9.69747
R2981 VDD2.n67 VDD2.n16 9.69747
R2982 VDD2.n94 VDD2.n93 9.69747
R2983 VDD2.n203 VDD2.n202 9.45567
R2984 VDD2.n100 VDD2.n99 9.45567
R2985 VDD2.n163 VDD2.n162 9.3005
R2986 VDD2.n122 VDD2.n121 9.3005
R2987 VDD2.n169 VDD2.n168 9.3005
R2988 VDD2.n171 VDD2.n170 9.3005
R2989 VDD2.n118 VDD2.n117 9.3005
R2990 VDD2.n177 VDD2.n176 9.3005
R2991 VDD2.n179 VDD2.n178 9.3005
R2992 VDD2.n115 VDD2.n112 9.3005
R2993 VDD2.n202 VDD2.n201 9.3005
R2994 VDD2.n105 VDD2.n104 9.3005
R2995 VDD2.n196 VDD2.n195 9.3005
R2996 VDD2.n194 VDD2.n193 9.3005
R2997 VDD2.n109 VDD2.n108 9.3005
R2998 VDD2.n188 VDD2.n187 9.3005
R2999 VDD2.n186 VDD2.n185 9.3005
R3000 VDD2.n161 VDD2.n160 9.3005
R3001 VDD2.n126 VDD2.n125 9.3005
R3002 VDD2.n155 VDD2.n154 9.3005
R3003 VDD2.n153 VDD2.n152 9.3005
R3004 VDD2.n130 VDD2.n129 9.3005
R3005 VDD2.n147 VDD2.n146 9.3005
R3006 VDD2.n145 VDD2.n144 9.3005
R3007 VDD2.n134 VDD2.n133 9.3005
R3008 VDD2.n139 VDD2.n138 9.3005
R3009 VDD2.n99 VDD2.n98 9.3005
R3010 VDD2.n2 VDD2.n1 9.3005
R3011 VDD2.n93 VDD2.n92 9.3005
R3012 VDD2.n91 VDD2.n90 9.3005
R3013 VDD2.n6 VDD2.n5 9.3005
R3014 VDD2.n85 VDD2.n84 9.3005
R3015 VDD2.n83 VDD2.n82 9.3005
R3016 VDD2.n22 VDD2.n21 9.3005
R3017 VDD2.n51 VDD2.n50 9.3005
R3018 VDD2.n49 VDD2.n48 9.3005
R3019 VDD2.n26 VDD2.n25 9.3005
R3020 VDD2.n43 VDD2.n42 9.3005
R3021 VDD2.n41 VDD2.n40 9.3005
R3022 VDD2.n30 VDD2.n29 9.3005
R3023 VDD2.n35 VDD2.n34 9.3005
R3024 VDD2.n57 VDD2.n56 9.3005
R3025 VDD2.n59 VDD2.n58 9.3005
R3026 VDD2.n18 VDD2.n17 9.3005
R3027 VDD2.n65 VDD2.n64 9.3005
R3028 VDD2.n67 VDD2.n66 9.3005
R3029 VDD2.n14 VDD2.n13 9.3005
R3030 VDD2.n73 VDD2.n72 9.3005
R3031 VDD2.n75 VDD2.n74 9.3005
R3032 VDD2.n76 VDD2.n9 9.3005
R3033 VDD2.n200 VDD2.n105 8.92171
R3034 VDD2.n168 VDD2.n167 8.92171
R3035 VDD2.n152 VDD2.n128 8.92171
R3036 VDD2.n48 VDD2.n24 8.92171
R3037 VDD2.n64 VDD2.n63 8.92171
R3038 VDD2.n97 VDD2.n2 8.92171
R3039 VDD2.n201 VDD2.n103 8.14595
R3040 VDD2.n164 VDD2.n122 8.14595
R3041 VDD2.n156 VDD2.n155 8.14595
R3042 VDD2.n52 VDD2.n51 8.14595
R3043 VDD2.n60 VDD2.n18 8.14595
R3044 VDD2.n98 VDD2.n0 8.14595
R3045 VDD2.n163 VDD2.n124 7.3702
R3046 VDD2.n159 VDD2.n126 7.3702
R3047 VDD2.n55 VDD2.n22 7.3702
R3048 VDD2.n59 VDD2.n20 7.3702
R3049 VDD2.n160 VDD2.n124 6.59444
R3050 VDD2.n160 VDD2.n159 6.59444
R3051 VDD2.n56 VDD2.n55 6.59444
R3052 VDD2.n56 VDD2.n20 6.59444
R3053 VDD2.n203 VDD2.n103 5.81868
R3054 VDD2.n164 VDD2.n163 5.81868
R3055 VDD2.n156 VDD2.n126 5.81868
R3056 VDD2.n52 VDD2.n22 5.81868
R3057 VDD2.n60 VDD2.n59 5.81868
R3058 VDD2.n100 VDD2.n0 5.81868
R3059 VDD2.n201 VDD2.n200 5.04292
R3060 VDD2.n167 VDD2.n122 5.04292
R3061 VDD2.n155 VDD2.n128 5.04292
R3062 VDD2.n51 VDD2.n24 5.04292
R3063 VDD2.n63 VDD2.n18 5.04292
R3064 VDD2.n98 VDD2.n97 5.04292
R3065 VDD2.n138 VDD2.n137 4.38563
R3066 VDD2.n34 VDD2.n33 4.38563
R3067 VDD2.n197 VDD2.n105 4.26717
R3068 VDD2.n168 VDD2.n120 4.26717
R3069 VDD2.n152 VDD2.n151 4.26717
R3070 VDD2.n48 VDD2.n47 4.26717
R3071 VDD2.n64 VDD2.n16 4.26717
R3072 VDD2.n94 VDD2.n2 4.26717
R3073 VDD2.n196 VDD2.n107 3.49141
R3074 VDD2.n172 VDD2.n171 3.49141
R3075 VDD2.n148 VDD2.n130 3.49141
R3076 VDD2.n44 VDD2.n26 3.49141
R3077 VDD2.n68 VDD2.n67 3.49141
R3078 VDD2.n93 VDD2.n4 3.49141
R3079 VDD2.n193 VDD2.n192 2.71565
R3080 VDD2.n175 VDD2.n118 2.71565
R3081 VDD2.n147 VDD2.n132 2.71565
R3082 VDD2.n43 VDD2.n28 2.71565
R3083 VDD2.n71 VDD2.n14 2.71565
R3084 VDD2.n90 VDD2.n89 2.71565
R3085 VDD2.n189 VDD2.n109 1.93989
R3086 VDD2.n176 VDD2.n116 1.93989
R3087 VDD2.n144 VDD2.n143 1.93989
R3088 VDD2.n40 VDD2.n39 1.93989
R3089 VDD2.n72 VDD2.n12 1.93989
R3090 VDD2.n86 VDD2.n6 1.93989
R3091 VDD2 VDD2.n204 1.75266
R3092 VDD2.n188 VDD2.n111 1.16414
R3093 VDD2.n180 VDD2.n179 1.16414
R3094 VDD2.n140 VDD2.n134 1.16414
R3095 VDD2.n36 VDD2.n30 1.16414
R3096 VDD2.n77 VDD2.n75 1.16414
R3097 VDD2.n85 VDD2.n8 1.16414
R3098 VDD2.n205 VDD2.t3 1.08424
R3099 VDD2.n205 VDD2.t0 1.08424
R3100 VDD2.n101 VDD2.t2 1.08424
R3101 VDD2.n101 VDD2.t4 1.08424
R3102 VDD2.n185 VDD2.n184 0.388379
R3103 VDD2.n115 VDD2.n113 0.388379
R3104 VDD2.n139 VDD2.n136 0.388379
R3105 VDD2.n35 VDD2.n32 0.388379
R3106 VDD2.n76 VDD2.n10 0.388379
R3107 VDD2.n82 VDD2.n81 0.388379
R3108 VDD2.n202 VDD2.n104 0.155672
R3109 VDD2.n195 VDD2.n104 0.155672
R3110 VDD2.n195 VDD2.n194 0.155672
R3111 VDD2.n194 VDD2.n108 0.155672
R3112 VDD2.n187 VDD2.n108 0.155672
R3113 VDD2.n187 VDD2.n186 0.155672
R3114 VDD2.n186 VDD2.n112 0.155672
R3115 VDD2.n178 VDD2.n112 0.155672
R3116 VDD2.n178 VDD2.n177 0.155672
R3117 VDD2.n177 VDD2.n117 0.155672
R3118 VDD2.n170 VDD2.n117 0.155672
R3119 VDD2.n170 VDD2.n169 0.155672
R3120 VDD2.n169 VDD2.n121 0.155672
R3121 VDD2.n162 VDD2.n121 0.155672
R3122 VDD2.n162 VDD2.n161 0.155672
R3123 VDD2.n161 VDD2.n125 0.155672
R3124 VDD2.n154 VDD2.n125 0.155672
R3125 VDD2.n154 VDD2.n153 0.155672
R3126 VDD2.n153 VDD2.n129 0.155672
R3127 VDD2.n146 VDD2.n129 0.155672
R3128 VDD2.n146 VDD2.n145 0.155672
R3129 VDD2.n145 VDD2.n133 0.155672
R3130 VDD2.n138 VDD2.n133 0.155672
R3131 VDD2.n34 VDD2.n29 0.155672
R3132 VDD2.n41 VDD2.n29 0.155672
R3133 VDD2.n42 VDD2.n41 0.155672
R3134 VDD2.n42 VDD2.n25 0.155672
R3135 VDD2.n49 VDD2.n25 0.155672
R3136 VDD2.n50 VDD2.n49 0.155672
R3137 VDD2.n50 VDD2.n21 0.155672
R3138 VDD2.n57 VDD2.n21 0.155672
R3139 VDD2.n58 VDD2.n57 0.155672
R3140 VDD2.n58 VDD2.n17 0.155672
R3141 VDD2.n65 VDD2.n17 0.155672
R3142 VDD2.n66 VDD2.n65 0.155672
R3143 VDD2.n66 VDD2.n13 0.155672
R3144 VDD2.n73 VDD2.n13 0.155672
R3145 VDD2.n74 VDD2.n73 0.155672
R3146 VDD2.n74 VDD2.n9 0.155672
R3147 VDD2.n83 VDD2.n9 0.155672
R3148 VDD2.n84 VDD2.n83 0.155672
R3149 VDD2.n84 VDD2.n5 0.155672
R3150 VDD2.n91 VDD2.n5 0.155672
R3151 VDD2.n92 VDD2.n91 0.155672
R3152 VDD2.n92 VDD2.n1 0.155672
R3153 VDD2.n99 VDD2.n1 0.155672
C0 VTAIL VP 9.6121f
C1 VTAIL VN 9.597671f
C2 VDD1 VP 10.062901f
C3 VDD1 VN 0.150198f
C4 VP VN 7.7848f
C5 VDD2 VTAIL 10.137f
C6 VDD2 VDD1 1.28627f
C7 VDD2 VP 0.432484f
C8 VDD2 VN 9.78513f
C9 VTAIL VDD1 10.0903f
C10 VDD2 B 6.867476f
C11 VDD1 B 6.97935f
C12 VTAIL B 10.09282f
C13 VN B 12.55378f
C14 VP B 10.998202f
C15 VDD2.n0 B 0.030265f
C16 VDD2.n1 B 0.021226f
C17 VDD2.n2 B 0.011406f
C18 VDD2.n3 B 0.026959f
C19 VDD2.n4 B 0.012077f
C20 VDD2.n5 B 0.021226f
C21 VDD2.n6 B 0.011406f
C22 VDD2.n7 B 0.026959f
C23 VDD2.n8 B 0.012077f
C24 VDD2.n9 B 0.021226f
C25 VDD2.n10 B 0.011741f
C26 VDD2.n11 B 0.026959f
C27 VDD2.n12 B 0.012077f
C28 VDD2.n13 B 0.021226f
C29 VDD2.n14 B 0.011406f
C30 VDD2.n15 B 0.026959f
C31 VDD2.n16 B 0.012077f
C32 VDD2.n17 B 0.021226f
C33 VDD2.n18 B 0.011406f
C34 VDD2.n19 B 0.026959f
C35 VDD2.n20 B 0.012077f
C36 VDD2.n21 B 0.021226f
C37 VDD2.n22 B 0.011406f
C38 VDD2.n23 B 0.026959f
C39 VDD2.n24 B 0.012077f
C40 VDD2.n25 B 0.021226f
C41 VDD2.n26 B 0.011406f
C42 VDD2.n27 B 0.026959f
C43 VDD2.n28 B 0.012077f
C44 VDD2.n29 B 0.021226f
C45 VDD2.n30 B 0.011406f
C46 VDD2.n31 B 0.02022f
C47 VDD2.n32 B 0.015926f
C48 VDD2.t1 B 0.044691f
C49 VDD2.n33 B 0.155843f
C50 VDD2.n34 B 1.6991f
C51 VDD2.n35 B 0.011406f
C52 VDD2.n36 B 0.012077f
C53 VDD2.n37 B 0.026959f
C54 VDD2.n38 B 0.026959f
C55 VDD2.n39 B 0.012077f
C56 VDD2.n40 B 0.011406f
C57 VDD2.n41 B 0.021226f
C58 VDD2.n42 B 0.021226f
C59 VDD2.n43 B 0.011406f
C60 VDD2.n44 B 0.012077f
C61 VDD2.n45 B 0.026959f
C62 VDD2.n46 B 0.026959f
C63 VDD2.n47 B 0.012077f
C64 VDD2.n48 B 0.011406f
C65 VDD2.n49 B 0.021226f
C66 VDD2.n50 B 0.021226f
C67 VDD2.n51 B 0.011406f
C68 VDD2.n52 B 0.012077f
C69 VDD2.n53 B 0.026959f
C70 VDD2.n54 B 0.026959f
C71 VDD2.n55 B 0.012077f
C72 VDD2.n56 B 0.011406f
C73 VDD2.n57 B 0.021226f
C74 VDD2.n58 B 0.021226f
C75 VDD2.n59 B 0.011406f
C76 VDD2.n60 B 0.012077f
C77 VDD2.n61 B 0.026959f
C78 VDD2.n62 B 0.026959f
C79 VDD2.n63 B 0.012077f
C80 VDD2.n64 B 0.011406f
C81 VDD2.n65 B 0.021226f
C82 VDD2.n66 B 0.021226f
C83 VDD2.n67 B 0.011406f
C84 VDD2.n68 B 0.012077f
C85 VDD2.n69 B 0.026959f
C86 VDD2.n70 B 0.026959f
C87 VDD2.n71 B 0.012077f
C88 VDD2.n72 B 0.011406f
C89 VDD2.n73 B 0.021226f
C90 VDD2.n74 B 0.021226f
C91 VDD2.n75 B 0.011406f
C92 VDD2.n76 B 0.011406f
C93 VDD2.n77 B 0.012077f
C94 VDD2.n78 B 0.026959f
C95 VDD2.n79 B 0.026959f
C96 VDD2.n80 B 0.026959f
C97 VDD2.n81 B 0.011741f
C98 VDD2.n82 B 0.011406f
C99 VDD2.n83 B 0.021226f
C100 VDD2.n84 B 0.021226f
C101 VDD2.n85 B 0.011406f
C102 VDD2.n86 B 0.012077f
C103 VDD2.n87 B 0.026959f
C104 VDD2.n88 B 0.026959f
C105 VDD2.n89 B 0.012077f
C106 VDD2.n90 B 0.011406f
C107 VDD2.n91 B 0.021226f
C108 VDD2.n92 B 0.021226f
C109 VDD2.n93 B 0.011406f
C110 VDD2.n94 B 0.012077f
C111 VDD2.n95 B 0.026959f
C112 VDD2.n96 B 0.059122f
C113 VDD2.n97 B 0.012077f
C114 VDD2.n98 B 0.011406f
C115 VDD2.n99 B 0.049933f
C116 VDD2.n100 B 0.052767f
C117 VDD2.t2 B 0.30645f
C118 VDD2.t4 B 0.30645f
C119 VDD2.n101 B 2.79683f
C120 VDD2.n102 B 2.49417f
C121 VDD2.n103 B 0.030265f
C122 VDD2.n104 B 0.021226f
C123 VDD2.n105 B 0.011406f
C124 VDD2.n106 B 0.026959f
C125 VDD2.n107 B 0.012077f
C126 VDD2.n108 B 0.021226f
C127 VDD2.n109 B 0.011406f
C128 VDD2.n110 B 0.026959f
C129 VDD2.n111 B 0.012077f
C130 VDD2.n112 B 0.021226f
C131 VDD2.n113 B 0.011741f
C132 VDD2.n114 B 0.026959f
C133 VDD2.n115 B 0.011406f
C134 VDD2.n116 B 0.012077f
C135 VDD2.n117 B 0.021226f
C136 VDD2.n118 B 0.011406f
C137 VDD2.n119 B 0.026959f
C138 VDD2.n120 B 0.012077f
C139 VDD2.n121 B 0.021226f
C140 VDD2.n122 B 0.011406f
C141 VDD2.n123 B 0.026959f
C142 VDD2.n124 B 0.012077f
C143 VDD2.n125 B 0.021226f
C144 VDD2.n126 B 0.011406f
C145 VDD2.n127 B 0.026959f
C146 VDD2.n128 B 0.012077f
C147 VDD2.n129 B 0.021226f
C148 VDD2.n130 B 0.011406f
C149 VDD2.n131 B 0.026959f
C150 VDD2.n132 B 0.012077f
C151 VDD2.n133 B 0.021226f
C152 VDD2.n134 B 0.011406f
C153 VDD2.n135 B 0.02022f
C154 VDD2.n136 B 0.015926f
C155 VDD2.t5 B 0.044691f
C156 VDD2.n137 B 0.155843f
C157 VDD2.n138 B 1.6991f
C158 VDD2.n139 B 0.011406f
C159 VDD2.n140 B 0.012077f
C160 VDD2.n141 B 0.026959f
C161 VDD2.n142 B 0.026959f
C162 VDD2.n143 B 0.012077f
C163 VDD2.n144 B 0.011406f
C164 VDD2.n145 B 0.021226f
C165 VDD2.n146 B 0.021226f
C166 VDD2.n147 B 0.011406f
C167 VDD2.n148 B 0.012077f
C168 VDD2.n149 B 0.026959f
C169 VDD2.n150 B 0.026959f
C170 VDD2.n151 B 0.012077f
C171 VDD2.n152 B 0.011406f
C172 VDD2.n153 B 0.021226f
C173 VDD2.n154 B 0.021226f
C174 VDD2.n155 B 0.011406f
C175 VDD2.n156 B 0.012077f
C176 VDD2.n157 B 0.026959f
C177 VDD2.n158 B 0.026959f
C178 VDD2.n159 B 0.012077f
C179 VDD2.n160 B 0.011406f
C180 VDD2.n161 B 0.021226f
C181 VDD2.n162 B 0.021226f
C182 VDD2.n163 B 0.011406f
C183 VDD2.n164 B 0.012077f
C184 VDD2.n165 B 0.026959f
C185 VDD2.n166 B 0.026959f
C186 VDD2.n167 B 0.012077f
C187 VDD2.n168 B 0.011406f
C188 VDD2.n169 B 0.021226f
C189 VDD2.n170 B 0.021226f
C190 VDD2.n171 B 0.011406f
C191 VDD2.n172 B 0.012077f
C192 VDD2.n173 B 0.026959f
C193 VDD2.n174 B 0.026959f
C194 VDD2.n175 B 0.012077f
C195 VDD2.n176 B 0.011406f
C196 VDD2.n177 B 0.021226f
C197 VDD2.n178 B 0.021226f
C198 VDD2.n179 B 0.011406f
C199 VDD2.n180 B 0.012077f
C200 VDD2.n181 B 0.026959f
C201 VDD2.n182 B 0.026959f
C202 VDD2.n183 B 0.026959f
C203 VDD2.n184 B 0.011741f
C204 VDD2.n185 B 0.011406f
C205 VDD2.n186 B 0.021226f
C206 VDD2.n187 B 0.021226f
C207 VDD2.n188 B 0.011406f
C208 VDD2.n189 B 0.012077f
C209 VDD2.n190 B 0.026959f
C210 VDD2.n191 B 0.026959f
C211 VDD2.n192 B 0.012077f
C212 VDD2.n193 B 0.011406f
C213 VDD2.n194 B 0.021226f
C214 VDD2.n195 B 0.021226f
C215 VDD2.n196 B 0.011406f
C216 VDD2.n197 B 0.012077f
C217 VDD2.n198 B 0.026959f
C218 VDD2.n199 B 0.059122f
C219 VDD2.n200 B 0.012077f
C220 VDD2.n201 B 0.011406f
C221 VDD2.n202 B 0.049933f
C222 VDD2.n203 B 0.047835f
C223 VDD2.n204 B 2.51043f
C224 VDD2.t3 B 0.30645f
C225 VDD2.t0 B 0.30645f
C226 VDD2.n205 B 2.7968f
C227 VN.n0 B 0.031953f
C228 VN.t1 B 2.78984f
C229 VN.n1 B 0.020737f
C230 VN.n2 B 0.208362f
C231 VN.t3 B 2.78984f
C232 VN.t4 B 2.95429f
C233 VN.n3 B 1.02129f
C234 VN.n4 B 1.03357f
C235 VN.n5 B 0.03402f
C236 VN.n6 B 0.048974f
C237 VN.n7 B 0.024236f
C238 VN.n8 B 0.024236f
C239 VN.n9 B 0.024236f
C240 VN.n10 B 0.04622f
C241 VN.n11 B 0.039372f
C242 VN.n12 B 1.05187f
C243 VN.n13 B 0.031899f
C244 VN.n14 B 0.031953f
C245 VN.t0 B 2.78984f
C246 VN.n15 B 0.020737f
C247 VN.n16 B 0.208362f
C248 VN.t2 B 2.78984f
C249 VN.t5 B 2.95429f
C250 VN.n17 B 1.02129f
C251 VN.n18 B 1.03357f
C252 VN.n19 B 0.03402f
C253 VN.n20 B 0.048974f
C254 VN.n21 B 0.024236f
C255 VN.n22 B 0.024236f
C256 VN.n23 B 0.024236f
C257 VN.n24 B 0.04622f
C258 VN.n25 B 0.039372f
C259 VN.n26 B 1.05187f
C260 VN.n27 B 1.44451f
C261 VDD1.n0 B 0.0306f
C262 VDD1.n1 B 0.021461f
C263 VDD1.n2 B 0.011532f
C264 VDD1.n3 B 0.027259f
C265 VDD1.n4 B 0.012211f
C266 VDD1.n5 B 0.021461f
C267 VDD1.n6 B 0.011532f
C268 VDD1.n7 B 0.027259f
C269 VDD1.n8 B 0.012211f
C270 VDD1.n9 B 0.021461f
C271 VDD1.n10 B 0.011872f
C272 VDD1.n11 B 0.027259f
C273 VDD1.n12 B 0.011532f
C274 VDD1.n13 B 0.012211f
C275 VDD1.n14 B 0.021461f
C276 VDD1.n15 B 0.011532f
C277 VDD1.n16 B 0.027259f
C278 VDD1.n17 B 0.012211f
C279 VDD1.n18 B 0.021461f
C280 VDD1.n19 B 0.011532f
C281 VDD1.n20 B 0.027259f
C282 VDD1.n21 B 0.012211f
C283 VDD1.n22 B 0.021461f
C284 VDD1.n23 B 0.011532f
C285 VDD1.n24 B 0.027259f
C286 VDD1.n25 B 0.012211f
C287 VDD1.n26 B 0.021461f
C288 VDD1.n27 B 0.011532f
C289 VDD1.n28 B 0.027259f
C290 VDD1.n29 B 0.012211f
C291 VDD1.n30 B 0.021461f
C292 VDD1.n31 B 0.011532f
C293 VDD1.n32 B 0.020444f
C294 VDD1.n33 B 0.016102f
C295 VDD1.t0 B 0.045187f
C296 VDD1.n34 B 0.157572f
C297 VDD1.n35 B 1.71794f
C298 VDD1.n36 B 0.011532f
C299 VDD1.n37 B 0.012211f
C300 VDD1.n38 B 0.027259f
C301 VDD1.n39 B 0.027259f
C302 VDD1.n40 B 0.012211f
C303 VDD1.n41 B 0.011532f
C304 VDD1.n42 B 0.021461f
C305 VDD1.n43 B 0.021461f
C306 VDD1.n44 B 0.011532f
C307 VDD1.n45 B 0.012211f
C308 VDD1.n46 B 0.027259f
C309 VDD1.n47 B 0.027259f
C310 VDD1.n48 B 0.012211f
C311 VDD1.n49 B 0.011532f
C312 VDD1.n50 B 0.021461f
C313 VDD1.n51 B 0.021461f
C314 VDD1.n52 B 0.011532f
C315 VDD1.n53 B 0.012211f
C316 VDD1.n54 B 0.027259f
C317 VDD1.n55 B 0.027259f
C318 VDD1.n56 B 0.012211f
C319 VDD1.n57 B 0.011532f
C320 VDD1.n58 B 0.021461f
C321 VDD1.n59 B 0.021461f
C322 VDD1.n60 B 0.011532f
C323 VDD1.n61 B 0.012211f
C324 VDD1.n62 B 0.027259f
C325 VDD1.n63 B 0.027259f
C326 VDD1.n64 B 0.012211f
C327 VDD1.n65 B 0.011532f
C328 VDD1.n66 B 0.021461f
C329 VDD1.n67 B 0.021461f
C330 VDD1.n68 B 0.011532f
C331 VDD1.n69 B 0.012211f
C332 VDD1.n70 B 0.027259f
C333 VDD1.n71 B 0.027259f
C334 VDD1.n72 B 0.012211f
C335 VDD1.n73 B 0.011532f
C336 VDD1.n74 B 0.021461f
C337 VDD1.n75 B 0.021461f
C338 VDD1.n76 B 0.011532f
C339 VDD1.n77 B 0.012211f
C340 VDD1.n78 B 0.027259f
C341 VDD1.n79 B 0.027259f
C342 VDD1.n80 B 0.027259f
C343 VDD1.n81 B 0.011872f
C344 VDD1.n82 B 0.011532f
C345 VDD1.n83 B 0.021461f
C346 VDD1.n84 B 0.021461f
C347 VDD1.n85 B 0.011532f
C348 VDD1.n86 B 0.012211f
C349 VDD1.n87 B 0.027259f
C350 VDD1.n88 B 0.027259f
C351 VDD1.n89 B 0.012211f
C352 VDD1.n90 B 0.011532f
C353 VDD1.n91 B 0.021461f
C354 VDD1.n92 B 0.021461f
C355 VDD1.n93 B 0.011532f
C356 VDD1.n94 B 0.012211f
C357 VDD1.n95 B 0.027259f
C358 VDD1.n96 B 0.059778f
C359 VDD1.n97 B 0.012211f
C360 VDD1.n98 B 0.011532f
C361 VDD1.n99 B 0.050487f
C362 VDD1.n100 B 0.053944f
C363 VDD1.n101 B 0.0306f
C364 VDD1.n102 B 0.021461f
C365 VDD1.n103 B 0.011532f
C366 VDD1.n104 B 0.027259f
C367 VDD1.n105 B 0.012211f
C368 VDD1.n106 B 0.021461f
C369 VDD1.n107 B 0.011532f
C370 VDD1.n108 B 0.027259f
C371 VDD1.n109 B 0.012211f
C372 VDD1.n110 B 0.021461f
C373 VDD1.n111 B 0.011872f
C374 VDD1.n112 B 0.027259f
C375 VDD1.n113 B 0.012211f
C376 VDD1.n114 B 0.021461f
C377 VDD1.n115 B 0.011532f
C378 VDD1.n116 B 0.027259f
C379 VDD1.n117 B 0.012211f
C380 VDD1.n118 B 0.021461f
C381 VDD1.n119 B 0.011532f
C382 VDD1.n120 B 0.027259f
C383 VDD1.n121 B 0.012211f
C384 VDD1.n122 B 0.021461f
C385 VDD1.n123 B 0.011532f
C386 VDD1.n124 B 0.027259f
C387 VDD1.n125 B 0.012211f
C388 VDD1.n126 B 0.021461f
C389 VDD1.n127 B 0.011532f
C390 VDD1.n128 B 0.027259f
C391 VDD1.n129 B 0.012211f
C392 VDD1.n130 B 0.021461f
C393 VDD1.n131 B 0.011532f
C394 VDD1.n132 B 0.020444f
C395 VDD1.n133 B 0.016102f
C396 VDD1.t1 B 0.045187f
C397 VDD1.n134 B 0.157572f
C398 VDD1.n135 B 1.71794f
C399 VDD1.n136 B 0.011532f
C400 VDD1.n137 B 0.012211f
C401 VDD1.n138 B 0.027259f
C402 VDD1.n139 B 0.027259f
C403 VDD1.n140 B 0.012211f
C404 VDD1.n141 B 0.011532f
C405 VDD1.n142 B 0.021461f
C406 VDD1.n143 B 0.021461f
C407 VDD1.n144 B 0.011532f
C408 VDD1.n145 B 0.012211f
C409 VDD1.n146 B 0.027259f
C410 VDD1.n147 B 0.027259f
C411 VDD1.n148 B 0.012211f
C412 VDD1.n149 B 0.011532f
C413 VDD1.n150 B 0.021461f
C414 VDD1.n151 B 0.021461f
C415 VDD1.n152 B 0.011532f
C416 VDD1.n153 B 0.012211f
C417 VDD1.n154 B 0.027259f
C418 VDD1.n155 B 0.027259f
C419 VDD1.n156 B 0.012211f
C420 VDD1.n157 B 0.011532f
C421 VDD1.n158 B 0.021461f
C422 VDD1.n159 B 0.021461f
C423 VDD1.n160 B 0.011532f
C424 VDD1.n161 B 0.012211f
C425 VDD1.n162 B 0.027259f
C426 VDD1.n163 B 0.027259f
C427 VDD1.n164 B 0.012211f
C428 VDD1.n165 B 0.011532f
C429 VDD1.n166 B 0.021461f
C430 VDD1.n167 B 0.021461f
C431 VDD1.n168 B 0.011532f
C432 VDD1.n169 B 0.012211f
C433 VDD1.n170 B 0.027259f
C434 VDD1.n171 B 0.027259f
C435 VDD1.n172 B 0.012211f
C436 VDD1.n173 B 0.011532f
C437 VDD1.n174 B 0.021461f
C438 VDD1.n175 B 0.021461f
C439 VDD1.n176 B 0.011532f
C440 VDD1.n177 B 0.011532f
C441 VDD1.n178 B 0.012211f
C442 VDD1.n179 B 0.027259f
C443 VDD1.n180 B 0.027259f
C444 VDD1.n181 B 0.027259f
C445 VDD1.n182 B 0.011872f
C446 VDD1.n183 B 0.011532f
C447 VDD1.n184 B 0.021461f
C448 VDD1.n185 B 0.021461f
C449 VDD1.n186 B 0.011532f
C450 VDD1.n187 B 0.012211f
C451 VDD1.n188 B 0.027259f
C452 VDD1.n189 B 0.027259f
C453 VDD1.n190 B 0.012211f
C454 VDD1.n191 B 0.011532f
C455 VDD1.n192 B 0.021461f
C456 VDD1.n193 B 0.021461f
C457 VDD1.n194 B 0.011532f
C458 VDD1.n195 B 0.012211f
C459 VDD1.n196 B 0.027259f
C460 VDD1.n197 B 0.059778f
C461 VDD1.n198 B 0.012211f
C462 VDD1.n199 B 0.011532f
C463 VDD1.n200 B 0.050487f
C464 VDD1.n201 B 0.053352f
C465 VDD1.t4 B 0.309849f
C466 VDD1.t3 B 0.309849f
C467 VDD1.n202 B 2.82785f
C468 VDD1.n203 B 2.62477f
C469 VDD1.t2 B 0.309849f
C470 VDD1.t5 B 0.309849f
C471 VDD1.n204 B 2.82472f
C472 VDD1.n205 B 2.72962f
C473 VTAIL.t1 B 0.322961f
C474 VTAIL.t3 B 0.322961f
C475 VTAIL.n0 B 2.87633f
C476 VTAIL.n1 B 0.383371f
C477 VTAIL.n2 B 0.031895f
C478 VTAIL.n3 B 0.02237f
C479 VTAIL.n4 B 0.012021f
C480 VTAIL.n5 B 0.028412f
C481 VTAIL.n6 B 0.012727f
C482 VTAIL.n7 B 0.02237f
C483 VTAIL.n8 B 0.012021f
C484 VTAIL.n9 B 0.028412f
C485 VTAIL.n10 B 0.012727f
C486 VTAIL.n11 B 0.02237f
C487 VTAIL.n12 B 0.012374f
C488 VTAIL.n13 B 0.028412f
C489 VTAIL.n14 B 0.012727f
C490 VTAIL.n15 B 0.02237f
C491 VTAIL.n16 B 0.012021f
C492 VTAIL.n17 B 0.028412f
C493 VTAIL.n18 B 0.012727f
C494 VTAIL.n19 B 0.02237f
C495 VTAIL.n20 B 0.012021f
C496 VTAIL.n21 B 0.028412f
C497 VTAIL.n22 B 0.012727f
C498 VTAIL.n23 B 0.02237f
C499 VTAIL.n24 B 0.012021f
C500 VTAIL.n25 B 0.028412f
C501 VTAIL.n26 B 0.012727f
C502 VTAIL.n27 B 0.02237f
C503 VTAIL.n28 B 0.012021f
C504 VTAIL.n29 B 0.028412f
C505 VTAIL.n30 B 0.012727f
C506 VTAIL.n31 B 0.02237f
C507 VTAIL.n32 B 0.012021f
C508 VTAIL.n33 B 0.021309f
C509 VTAIL.n34 B 0.016784f
C510 VTAIL.t11 B 0.047099f
C511 VTAIL.n35 B 0.164239f
C512 VTAIL.n36 B 1.79064f
C513 VTAIL.n37 B 0.012021f
C514 VTAIL.n38 B 0.012727f
C515 VTAIL.n39 B 0.028412f
C516 VTAIL.n40 B 0.028412f
C517 VTAIL.n41 B 0.012727f
C518 VTAIL.n42 B 0.012021f
C519 VTAIL.n43 B 0.02237f
C520 VTAIL.n44 B 0.02237f
C521 VTAIL.n45 B 0.012021f
C522 VTAIL.n46 B 0.012727f
C523 VTAIL.n47 B 0.028412f
C524 VTAIL.n48 B 0.028412f
C525 VTAIL.n49 B 0.012727f
C526 VTAIL.n50 B 0.012021f
C527 VTAIL.n51 B 0.02237f
C528 VTAIL.n52 B 0.02237f
C529 VTAIL.n53 B 0.012021f
C530 VTAIL.n54 B 0.012727f
C531 VTAIL.n55 B 0.028412f
C532 VTAIL.n56 B 0.028412f
C533 VTAIL.n57 B 0.012727f
C534 VTAIL.n58 B 0.012021f
C535 VTAIL.n59 B 0.02237f
C536 VTAIL.n60 B 0.02237f
C537 VTAIL.n61 B 0.012021f
C538 VTAIL.n62 B 0.012727f
C539 VTAIL.n63 B 0.028412f
C540 VTAIL.n64 B 0.028412f
C541 VTAIL.n65 B 0.012727f
C542 VTAIL.n66 B 0.012021f
C543 VTAIL.n67 B 0.02237f
C544 VTAIL.n68 B 0.02237f
C545 VTAIL.n69 B 0.012021f
C546 VTAIL.n70 B 0.012727f
C547 VTAIL.n71 B 0.028412f
C548 VTAIL.n72 B 0.028412f
C549 VTAIL.n73 B 0.012727f
C550 VTAIL.n74 B 0.012021f
C551 VTAIL.n75 B 0.02237f
C552 VTAIL.n76 B 0.02237f
C553 VTAIL.n77 B 0.012021f
C554 VTAIL.n78 B 0.012021f
C555 VTAIL.n79 B 0.012727f
C556 VTAIL.n80 B 0.028412f
C557 VTAIL.n81 B 0.028412f
C558 VTAIL.n82 B 0.028412f
C559 VTAIL.n83 B 0.012374f
C560 VTAIL.n84 B 0.012021f
C561 VTAIL.n85 B 0.02237f
C562 VTAIL.n86 B 0.02237f
C563 VTAIL.n87 B 0.012021f
C564 VTAIL.n88 B 0.012727f
C565 VTAIL.n89 B 0.028412f
C566 VTAIL.n90 B 0.028412f
C567 VTAIL.n91 B 0.012727f
C568 VTAIL.n92 B 0.012021f
C569 VTAIL.n93 B 0.02237f
C570 VTAIL.n94 B 0.02237f
C571 VTAIL.n95 B 0.012021f
C572 VTAIL.n96 B 0.012727f
C573 VTAIL.n97 B 0.028412f
C574 VTAIL.n98 B 0.062308f
C575 VTAIL.n99 B 0.012727f
C576 VTAIL.n100 B 0.012021f
C577 VTAIL.n101 B 0.052623f
C578 VTAIL.n102 B 0.034974f
C579 VTAIL.n103 B 0.29769f
C580 VTAIL.t8 B 0.322961f
C581 VTAIL.t9 B 0.322961f
C582 VTAIL.n104 B 2.87633f
C583 VTAIL.n105 B 2.15074f
C584 VTAIL.t2 B 0.322961f
C585 VTAIL.t4 B 0.322961f
C586 VTAIL.n106 B 2.87634f
C587 VTAIL.n107 B 2.15072f
C588 VTAIL.n108 B 0.031895f
C589 VTAIL.n109 B 0.02237f
C590 VTAIL.n110 B 0.012021f
C591 VTAIL.n111 B 0.028412f
C592 VTAIL.n112 B 0.012727f
C593 VTAIL.n113 B 0.02237f
C594 VTAIL.n114 B 0.012021f
C595 VTAIL.n115 B 0.028412f
C596 VTAIL.n116 B 0.012727f
C597 VTAIL.n117 B 0.02237f
C598 VTAIL.n118 B 0.012374f
C599 VTAIL.n119 B 0.028412f
C600 VTAIL.n120 B 0.012021f
C601 VTAIL.n121 B 0.012727f
C602 VTAIL.n122 B 0.02237f
C603 VTAIL.n123 B 0.012021f
C604 VTAIL.n124 B 0.028412f
C605 VTAIL.n125 B 0.012727f
C606 VTAIL.n126 B 0.02237f
C607 VTAIL.n127 B 0.012021f
C608 VTAIL.n128 B 0.028412f
C609 VTAIL.n129 B 0.012727f
C610 VTAIL.n130 B 0.02237f
C611 VTAIL.n131 B 0.012021f
C612 VTAIL.n132 B 0.028412f
C613 VTAIL.n133 B 0.012727f
C614 VTAIL.n134 B 0.02237f
C615 VTAIL.n135 B 0.012021f
C616 VTAIL.n136 B 0.028412f
C617 VTAIL.n137 B 0.012727f
C618 VTAIL.n138 B 0.02237f
C619 VTAIL.n139 B 0.012021f
C620 VTAIL.n140 B 0.021309f
C621 VTAIL.n141 B 0.016784f
C622 VTAIL.t0 B 0.047099f
C623 VTAIL.n142 B 0.164239f
C624 VTAIL.n143 B 1.79064f
C625 VTAIL.n144 B 0.012021f
C626 VTAIL.n145 B 0.012727f
C627 VTAIL.n146 B 0.028412f
C628 VTAIL.n147 B 0.028412f
C629 VTAIL.n148 B 0.012727f
C630 VTAIL.n149 B 0.012021f
C631 VTAIL.n150 B 0.02237f
C632 VTAIL.n151 B 0.02237f
C633 VTAIL.n152 B 0.012021f
C634 VTAIL.n153 B 0.012727f
C635 VTAIL.n154 B 0.028412f
C636 VTAIL.n155 B 0.028412f
C637 VTAIL.n156 B 0.012727f
C638 VTAIL.n157 B 0.012021f
C639 VTAIL.n158 B 0.02237f
C640 VTAIL.n159 B 0.02237f
C641 VTAIL.n160 B 0.012021f
C642 VTAIL.n161 B 0.012727f
C643 VTAIL.n162 B 0.028412f
C644 VTAIL.n163 B 0.028412f
C645 VTAIL.n164 B 0.012727f
C646 VTAIL.n165 B 0.012021f
C647 VTAIL.n166 B 0.02237f
C648 VTAIL.n167 B 0.02237f
C649 VTAIL.n168 B 0.012021f
C650 VTAIL.n169 B 0.012727f
C651 VTAIL.n170 B 0.028412f
C652 VTAIL.n171 B 0.028412f
C653 VTAIL.n172 B 0.012727f
C654 VTAIL.n173 B 0.012021f
C655 VTAIL.n174 B 0.02237f
C656 VTAIL.n175 B 0.02237f
C657 VTAIL.n176 B 0.012021f
C658 VTAIL.n177 B 0.012727f
C659 VTAIL.n178 B 0.028412f
C660 VTAIL.n179 B 0.028412f
C661 VTAIL.n180 B 0.012727f
C662 VTAIL.n181 B 0.012021f
C663 VTAIL.n182 B 0.02237f
C664 VTAIL.n183 B 0.02237f
C665 VTAIL.n184 B 0.012021f
C666 VTAIL.n185 B 0.012727f
C667 VTAIL.n186 B 0.028412f
C668 VTAIL.n187 B 0.028412f
C669 VTAIL.n188 B 0.028412f
C670 VTAIL.n189 B 0.012374f
C671 VTAIL.n190 B 0.012021f
C672 VTAIL.n191 B 0.02237f
C673 VTAIL.n192 B 0.02237f
C674 VTAIL.n193 B 0.012021f
C675 VTAIL.n194 B 0.012727f
C676 VTAIL.n195 B 0.028412f
C677 VTAIL.n196 B 0.028412f
C678 VTAIL.n197 B 0.012727f
C679 VTAIL.n198 B 0.012021f
C680 VTAIL.n199 B 0.02237f
C681 VTAIL.n200 B 0.02237f
C682 VTAIL.n201 B 0.012021f
C683 VTAIL.n202 B 0.012727f
C684 VTAIL.n203 B 0.028412f
C685 VTAIL.n204 B 0.062308f
C686 VTAIL.n205 B 0.012727f
C687 VTAIL.n206 B 0.012021f
C688 VTAIL.n207 B 0.052623f
C689 VTAIL.n208 B 0.034974f
C690 VTAIL.n209 B 0.29769f
C691 VTAIL.t10 B 0.322961f
C692 VTAIL.t6 B 0.322961f
C693 VTAIL.n210 B 2.87634f
C694 VTAIL.n211 B 0.501265f
C695 VTAIL.n212 B 0.031895f
C696 VTAIL.n213 B 0.02237f
C697 VTAIL.n214 B 0.012021f
C698 VTAIL.n215 B 0.028412f
C699 VTAIL.n216 B 0.012727f
C700 VTAIL.n217 B 0.02237f
C701 VTAIL.n218 B 0.012021f
C702 VTAIL.n219 B 0.028412f
C703 VTAIL.n220 B 0.012727f
C704 VTAIL.n221 B 0.02237f
C705 VTAIL.n222 B 0.012374f
C706 VTAIL.n223 B 0.028412f
C707 VTAIL.n224 B 0.012021f
C708 VTAIL.n225 B 0.012727f
C709 VTAIL.n226 B 0.02237f
C710 VTAIL.n227 B 0.012021f
C711 VTAIL.n228 B 0.028412f
C712 VTAIL.n229 B 0.012727f
C713 VTAIL.n230 B 0.02237f
C714 VTAIL.n231 B 0.012021f
C715 VTAIL.n232 B 0.028412f
C716 VTAIL.n233 B 0.012727f
C717 VTAIL.n234 B 0.02237f
C718 VTAIL.n235 B 0.012021f
C719 VTAIL.n236 B 0.028412f
C720 VTAIL.n237 B 0.012727f
C721 VTAIL.n238 B 0.02237f
C722 VTAIL.n239 B 0.012021f
C723 VTAIL.n240 B 0.028412f
C724 VTAIL.n241 B 0.012727f
C725 VTAIL.n242 B 0.02237f
C726 VTAIL.n243 B 0.012021f
C727 VTAIL.n244 B 0.021309f
C728 VTAIL.n245 B 0.016784f
C729 VTAIL.t7 B 0.047099f
C730 VTAIL.n246 B 0.164239f
C731 VTAIL.n247 B 1.79064f
C732 VTAIL.n248 B 0.012021f
C733 VTAIL.n249 B 0.012727f
C734 VTAIL.n250 B 0.028412f
C735 VTAIL.n251 B 0.028412f
C736 VTAIL.n252 B 0.012727f
C737 VTAIL.n253 B 0.012021f
C738 VTAIL.n254 B 0.02237f
C739 VTAIL.n255 B 0.02237f
C740 VTAIL.n256 B 0.012021f
C741 VTAIL.n257 B 0.012727f
C742 VTAIL.n258 B 0.028412f
C743 VTAIL.n259 B 0.028412f
C744 VTAIL.n260 B 0.012727f
C745 VTAIL.n261 B 0.012021f
C746 VTAIL.n262 B 0.02237f
C747 VTAIL.n263 B 0.02237f
C748 VTAIL.n264 B 0.012021f
C749 VTAIL.n265 B 0.012727f
C750 VTAIL.n266 B 0.028412f
C751 VTAIL.n267 B 0.028412f
C752 VTAIL.n268 B 0.012727f
C753 VTAIL.n269 B 0.012021f
C754 VTAIL.n270 B 0.02237f
C755 VTAIL.n271 B 0.02237f
C756 VTAIL.n272 B 0.012021f
C757 VTAIL.n273 B 0.012727f
C758 VTAIL.n274 B 0.028412f
C759 VTAIL.n275 B 0.028412f
C760 VTAIL.n276 B 0.012727f
C761 VTAIL.n277 B 0.012021f
C762 VTAIL.n278 B 0.02237f
C763 VTAIL.n279 B 0.02237f
C764 VTAIL.n280 B 0.012021f
C765 VTAIL.n281 B 0.012727f
C766 VTAIL.n282 B 0.028412f
C767 VTAIL.n283 B 0.028412f
C768 VTAIL.n284 B 0.012727f
C769 VTAIL.n285 B 0.012021f
C770 VTAIL.n286 B 0.02237f
C771 VTAIL.n287 B 0.02237f
C772 VTAIL.n288 B 0.012021f
C773 VTAIL.n289 B 0.012727f
C774 VTAIL.n290 B 0.028412f
C775 VTAIL.n291 B 0.028412f
C776 VTAIL.n292 B 0.028412f
C777 VTAIL.n293 B 0.012374f
C778 VTAIL.n294 B 0.012021f
C779 VTAIL.n295 B 0.02237f
C780 VTAIL.n296 B 0.02237f
C781 VTAIL.n297 B 0.012021f
C782 VTAIL.n298 B 0.012727f
C783 VTAIL.n299 B 0.028412f
C784 VTAIL.n300 B 0.028412f
C785 VTAIL.n301 B 0.012727f
C786 VTAIL.n302 B 0.012021f
C787 VTAIL.n303 B 0.02237f
C788 VTAIL.n304 B 0.02237f
C789 VTAIL.n305 B 0.012021f
C790 VTAIL.n306 B 0.012727f
C791 VTAIL.n307 B 0.028412f
C792 VTAIL.n308 B 0.062308f
C793 VTAIL.n309 B 0.012727f
C794 VTAIL.n310 B 0.012021f
C795 VTAIL.n311 B 0.052623f
C796 VTAIL.n312 B 0.034974f
C797 VTAIL.n313 B 1.78435f
C798 VTAIL.n314 B 0.031895f
C799 VTAIL.n315 B 0.02237f
C800 VTAIL.n316 B 0.012021f
C801 VTAIL.n317 B 0.028412f
C802 VTAIL.n318 B 0.012727f
C803 VTAIL.n319 B 0.02237f
C804 VTAIL.n320 B 0.012021f
C805 VTAIL.n321 B 0.028412f
C806 VTAIL.n322 B 0.012727f
C807 VTAIL.n323 B 0.02237f
C808 VTAIL.n324 B 0.012374f
C809 VTAIL.n325 B 0.028412f
C810 VTAIL.n326 B 0.012727f
C811 VTAIL.n327 B 0.02237f
C812 VTAIL.n328 B 0.012021f
C813 VTAIL.n329 B 0.028412f
C814 VTAIL.n330 B 0.012727f
C815 VTAIL.n331 B 0.02237f
C816 VTAIL.n332 B 0.012021f
C817 VTAIL.n333 B 0.028412f
C818 VTAIL.n334 B 0.012727f
C819 VTAIL.n335 B 0.02237f
C820 VTAIL.n336 B 0.012021f
C821 VTAIL.n337 B 0.028412f
C822 VTAIL.n338 B 0.012727f
C823 VTAIL.n339 B 0.02237f
C824 VTAIL.n340 B 0.012021f
C825 VTAIL.n341 B 0.028412f
C826 VTAIL.n342 B 0.012727f
C827 VTAIL.n343 B 0.02237f
C828 VTAIL.n344 B 0.012021f
C829 VTAIL.n345 B 0.021309f
C830 VTAIL.n346 B 0.016784f
C831 VTAIL.t5 B 0.047099f
C832 VTAIL.n347 B 0.164239f
C833 VTAIL.n348 B 1.79064f
C834 VTAIL.n349 B 0.012021f
C835 VTAIL.n350 B 0.012727f
C836 VTAIL.n351 B 0.028412f
C837 VTAIL.n352 B 0.028412f
C838 VTAIL.n353 B 0.012727f
C839 VTAIL.n354 B 0.012021f
C840 VTAIL.n355 B 0.02237f
C841 VTAIL.n356 B 0.02237f
C842 VTAIL.n357 B 0.012021f
C843 VTAIL.n358 B 0.012727f
C844 VTAIL.n359 B 0.028412f
C845 VTAIL.n360 B 0.028412f
C846 VTAIL.n361 B 0.012727f
C847 VTAIL.n362 B 0.012021f
C848 VTAIL.n363 B 0.02237f
C849 VTAIL.n364 B 0.02237f
C850 VTAIL.n365 B 0.012021f
C851 VTAIL.n366 B 0.012727f
C852 VTAIL.n367 B 0.028412f
C853 VTAIL.n368 B 0.028412f
C854 VTAIL.n369 B 0.012727f
C855 VTAIL.n370 B 0.012021f
C856 VTAIL.n371 B 0.02237f
C857 VTAIL.n372 B 0.02237f
C858 VTAIL.n373 B 0.012021f
C859 VTAIL.n374 B 0.012727f
C860 VTAIL.n375 B 0.028412f
C861 VTAIL.n376 B 0.028412f
C862 VTAIL.n377 B 0.012727f
C863 VTAIL.n378 B 0.012021f
C864 VTAIL.n379 B 0.02237f
C865 VTAIL.n380 B 0.02237f
C866 VTAIL.n381 B 0.012021f
C867 VTAIL.n382 B 0.012727f
C868 VTAIL.n383 B 0.028412f
C869 VTAIL.n384 B 0.028412f
C870 VTAIL.n385 B 0.012727f
C871 VTAIL.n386 B 0.012021f
C872 VTAIL.n387 B 0.02237f
C873 VTAIL.n388 B 0.02237f
C874 VTAIL.n389 B 0.012021f
C875 VTAIL.n390 B 0.012021f
C876 VTAIL.n391 B 0.012727f
C877 VTAIL.n392 B 0.028412f
C878 VTAIL.n393 B 0.028412f
C879 VTAIL.n394 B 0.028412f
C880 VTAIL.n395 B 0.012374f
C881 VTAIL.n396 B 0.012021f
C882 VTAIL.n397 B 0.02237f
C883 VTAIL.n398 B 0.02237f
C884 VTAIL.n399 B 0.012021f
C885 VTAIL.n400 B 0.012727f
C886 VTAIL.n401 B 0.028412f
C887 VTAIL.n402 B 0.028412f
C888 VTAIL.n403 B 0.012727f
C889 VTAIL.n404 B 0.012021f
C890 VTAIL.n405 B 0.02237f
C891 VTAIL.n406 B 0.02237f
C892 VTAIL.n407 B 0.012021f
C893 VTAIL.n408 B 0.012727f
C894 VTAIL.n409 B 0.028412f
C895 VTAIL.n410 B 0.062308f
C896 VTAIL.n411 B 0.012727f
C897 VTAIL.n412 B 0.012021f
C898 VTAIL.n413 B 0.052623f
C899 VTAIL.n414 B 0.034974f
C900 VTAIL.n415 B 1.73945f
C901 VP.n0 B 0.032346f
C902 VP.t2 B 2.82415f
C903 VP.n1 B 0.020992f
C904 VP.n2 B 0.024534f
C905 VP.t1 B 2.82415f
C906 VP.n3 B 0.049576f
C907 VP.n4 B 0.024534f
C908 VP.t4 B 2.82415f
C909 VP.n5 B 1.06481f
C910 VP.n6 B 0.032346f
C911 VP.t0 B 2.82415f
C912 VP.n7 B 0.020992f
C913 VP.n8 B 0.210925f
C914 VP.t3 B 2.82415f
C915 VP.t5 B 2.99062f
C916 VP.n9 B 1.03384f
C917 VP.n10 B 1.04629f
C918 VP.n11 B 0.034438f
C919 VP.n12 B 0.049576f
C920 VP.n13 B 0.024534f
C921 VP.n14 B 0.024534f
C922 VP.n15 B 0.024534f
C923 VP.n16 B 0.046789f
C924 VP.n17 B 0.039856f
C925 VP.n18 B 1.06481f
C926 VP.n19 B 1.44918f
C927 VP.n20 B 1.46605f
C928 VP.n21 B 0.032346f
C929 VP.n22 B 0.039856f
C930 VP.n23 B 0.046789f
C931 VP.n24 B 0.020992f
C932 VP.n25 B 0.024534f
C933 VP.n26 B 0.024534f
C934 VP.n27 B 0.024534f
C935 VP.n28 B 0.034438f
C936 VP.n29 B 0.981454f
C937 VP.n30 B 0.034438f
C938 VP.n31 B 0.049576f
C939 VP.n32 B 0.024534f
C940 VP.n33 B 0.024534f
C941 VP.n34 B 0.024534f
C942 VP.n35 B 0.046789f
C943 VP.n36 B 0.039856f
C944 VP.n37 B 1.06481f
C945 VP.n38 B 0.032291f
.ends

