* NGSPICE file created from diff_pair_sample_0379.ext - technology: sky130A

.subckt diff_pair_sample_0379 VTAIL VN VP B VDD2 VDD1
X0 B.t15 B.t13 B.t14 B.t7 sky130_fd_pr__nfet_01v8 ad=6.4428 pd=33.82 as=0 ps=0 w=16.52 l=2.77
X1 VDD1.t1 VP.t0 VTAIL.t3 B.t0 sky130_fd_pr__nfet_01v8 ad=6.4428 pd=33.82 as=6.4428 ps=33.82 w=16.52 l=2.77
X2 B.t12 B.t10 B.t11 B.t3 sky130_fd_pr__nfet_01v8 ad=6.4428 pd=33.82 as=0 ps=0 w=16.52 l=2.77
X3 VDD1.t0 VP.t1 VTAIL.t2 B.t1 sky130_fd_pr__nfet_01v8 ad=6.4428 pd=33.82 as=6.4428 ps=33.82 w=16.52 l=2.77
X4 VDD2.t1 VN.t0 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=6.4428 pd=33.82 as=6.4428 ps=33.82 w=16.52 l=2.77
X5 B.t9 B.t6 B.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=6.4428 pd=33.82 as=0 ps=0 w=16.52 l=2.77
X6 B.t5 B.t2 B.t4 B.t3 sky130_fd_pr__nfet_01v8 ad=6.4428 pd=33.82 as=0 ps=0 w=16.52 l=2.77
X7 VDD2.t0 VN.t1 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=6.4428 pd=33.82 as=6.4428 ps=33.82 w=16.52 l=2.77
R0 B.n583 B.n582 585
R1 B.n583 B.n51 585
R2 B.n586 B.n585 585
R3 B.n587 B.n115 585
R4 B.n589 B.n588 585
R5 B.n591 B.n114 585
R6 B.n594 B.n593 585
R7 B.n595 B.n113 585
R8 B.n597 B.n596 585
R9 B.n599 B.n112 585
R10 B.n602 B.n601 585
R11 B.n603 B.n111 585
R12 B.n605 B.n604 585
R13 B.n607 B.n110 585
R14 B.n610 B.n609 585
R15 B.n611 B.n109 585
R16 B.n613 B.n612 585
R17 B.n615 B.n108 585
R18 B.n618 B.n617 585
R19 B.n619 B.n107 585
R20 B.n621 B.n620 585
R21 B.n623 B.n106 585
R22 B.n626 B.n625 585
R23 B.n627 B.n105 585
R24 B.n629 B.n628 585
R25 B.n631 B.n104 585
R26 B.n634 B.n633 585
R27 B.n635 B.n103 585
R28 B.n637 B.n636 585
R29 B.n639 B.n102 585
R30 B.n642 B.n641 585
R31 B.n643 B.n101 585
R32 B.n645 B.n644 585
R33 B.n647 B.n100 585
R34 B.n650 B.n649 585
R35 B.n651 B.n99 585
R36 B.n653 B.n652 585
R37 B.n655 B.n98 585
R38 B.n658 B.n657 585
R39 B.n659 B.n97 585
R40 B.n661 B.n660 585
R41 B.n663 B.n96 585
R42 B.n666 B.n665 585
R43 B.n667 B.n95 585
R44 B.n669 B.n668 585
R45 B.n671 B.n94 585
R46 B.n674 B.n673 585
R47 B.n675 B.n93 585
R48 B.n677 B.n676 585
R49 B.n679 B.n92 585
R50 B.n682 B.n681 585
R51 B.n683 B.n91 585
R52 B.n685 B.n684 585
R53 B.n687 B.n90 585
R54 B.n690 B.n689 585
R55 B.n691 B.n87 585
R56 B.n694 B.n693 585
R57 B.n696 B.n86 585
R58 B.n699 B.n698 585
R59 B.n700 B.n85 585
R60 B.n702 B.n701 585
R61 B.n704 B.n84 585
R62 B.n707 B.n706 585
R63 B.n708 B.n80 585
R64 B.n710 B.n709 585
R65 B.n712 B.n79 585
R66 B.n715 B.n714 585
R67 B.n716 B.n78 585
R68 B.n718 B.n717 585
R69 B.n720 B.n77 585
R70 B.n723 B.n722 585
R71 B.n724 B.n76 585
R72 B.n726 B.n725 585
R73 B.n728 B.n75 585
R74 B.n731 B.n730 585
R75 B.n732 B.n74 585
R76 B.n734 B.n733 585
R77 B.n736 B.n73 585
R78 B.n739 B.n738 585
R79 B.n740 B.n72 585
R80 B.n742 B.n741 585
R81 B.n744 B.n71 585
R82 B.n747 B.n746 585
R83 B.n748 B.n70 585
R84 B.n750 B.n749 585
R85 B.n752 B.n69 585
R86 B.n755 B.n754 585
R87 B.n756 B.n68 585
R88 B.n758 B.n757 585
R89 B.n760 B.n67 585
R90 B.n763 B.n762 585
R91 B.n764 B.n66 585
R92 B.n766 B.n765 585
R93 B.n768 B.n65 585
R94 B.n771 B.n770 585
R95 B.n772 B.n64 585
R96 B.n774 B.n773 585
R97 B.n776 B.n63 585
R98 B.n779 B.n778 585
R99 B.n780 B.n62 585
R100 B.n782 B.n781 585
R101 B.n784 B.n61 585
R102 B.n787 B.n786 585
R103 B.n788 B.n60 585
R104 B.n790 B.n789 585
R105 B.n792 B.n59 585
R106 B.n795 B.n794 585
R107 B.n796 B.n58 585
R108 B.n798 B.n797 585
R109 B.n800 B.n57 585
R110 B.n803 B.n802 585
R111 B.n804 B.n56 585
R112 B.n806 B.n805 585
R113 B.n808 B.n55 585
R114 B.n811 B.n810 585
R115 B.n812 B.n54 585
R116 B.n814 B.n813 585
R117 B.n816 B.n53 585
R118 B.n819 B.n818 585
R119 B.n820 B.n52 585
R120 B.n581 B.n50 585
R121 B.n823 B.n50 585
R122 B.n580 B.n49 585
R123 B.n824 B.n49 585
R124 B.n579 B.n48 585
R125 B.n825 B.n48 585
R126 B.n578 B.n577 585
R127 B.n577 B.n44 585
R128 B.n576 B.n43 585
R129 B.n831 B.n43 585
R130 B.n575 B.n42 585
R131 B.n832 B.n42 585
R132 B.n574 B.n41 585
R133 B.n833 B.n41 585
R134 B.n573 B.n572 585
R135 B.n572 B.n37 585
R136 B.n571 B.n36 585
R137 B.n839 B.n36 585
R138 B.n570 B.n35 585
R139 B.n840 B.n35 585
R140 B.n569 B.n34 585
R141 B.n841 B.n34 585
R142 B.n568 B.n567 585
R143 B.n567 B.n30 585
R144 B.n566 B.n29 585
R145 B.n847 B.n29 585
R146 B.n565 B.n28 585
R147 B.n848 B.n28 585
R148 B.n564 B.n27 585
R149 B.n849 B.n27 585
R150 B.n563 B.n562 585
R151 B.n562 B.n23 585
R152 B.n561 B.n22 585
R153 B.n855 B.n22 585
R154 B.n560 B.n21 585
R155 B.n856 B.n21 585
R156 B.n559 B.n20 585
R157 B.n857 B.n20 585
R158 B.n558 B.n557 585
R159 B.n557 B.n16 585
R160 B.n556 B.n15 585
R161 B.n863 B.n15 585
R162 B.n555 B.n14 585
R163 B.n864 B.n14 585
R164 B.n554 B.n13 585
R165 B.n865 B.n13 585
R166 B.n553 B.n552 585
R167 B.n552 B.n12 585
R168 B.n551 B.n550 585
R169 B.n551 B.n8 585
R170 B.n549 B.n7 585
R171 B.n872 B.n7 585
R172 B.n548 B.n6 585
R173 B.n873 B.n6 585
R174 B.n547 B.n5 585
R175 B.n874 B.n5 585
R176 B.n546 B.n545 585
R177 B.n545 B.n4 585
R178 B.n544 B.n116 585
R179 B.n544 B.n543 585
R180 B.n534 B.n117 585
R181 B.n118 B.n117 585
R182 B.n536 B.n535 585
R183 B.n537 B.n536 585
R184 B.n533 B.n123 585
R185 B.n123 B.n122 585
R186 B.n532 B.n531 585
R187 B.n531 B.n530 585
R188 B.n125 B.n124 585
R189 B.n126 B.n125 585
R190 B.n523 B.n522 585
R191 B.n524 B.n523 585
R192 B.n521 B.n131 585
R193 B.n131 B.n130 585
R194 B.n520 B.n519 585
R195 B.n519 B.n518 585
R196 B.n133 B.n132 585
R197 B.n134 B.n133 585
R198 B.n511 B.n510 585
R199 B.n512 B.n511 585
R200 B.n509 B.n139 585
R201 B.n139 B.n138 585
R202 B.n508 B.n507 585
R203 B.n507 B.n506 585
R204 B.n141 B.n140 585
R205 B.n142 B.n141 585
R206 B.n499 B.n498 585
R207 B.n500 B.n499 585
R208 B.n497 B.n147 585
R209 B.n147 B.n146 585
R210 B.n496 B.n495 585
R211 B.n495 B.n494 585
R212 B.n149 B.n148 585
R213 B.n150 B.n149 585
R214 B.n487 B.n486 585
R215 B.n488 B.n487 585
R216 B.n485 B.n155 585
R217 B.n155 B.n154 585
R218 B.n484 B.n483 585
R219 B.n483 B.n482 585
R220 B.n157 B.n156 585
R221 B.n158 B.n157 585
R222 B.n475 B.n474 585
R223 B.n476 B.n475 585
R224 B.n473 B.n163 585
R225 B.n163 B.n162 585
R226 B.n472 B.n471 585
R227 B.n471 B.n470 585
R228 B.n467 B.n167 585
R229 B.n466 B.n465 585
R230 B.n463 B.n168 585
R231 B.n463 B.n166 585
R232 B.n462 B.n461 585
R233 B.n460 B.n459 585
R234 B.n458 B.n170 585
R235 B.n456 B.n455 585
R236 B.n454 B.n171 585
R237 B.n453 B.n452 585
R238 B.n450 B.n172 585
R239 B.n448 B.n447 585
R240 B.n446 B.n173 585
R241 B.n445 B.n444 585
R242 B.n442 B.n174 585
R243 B.n440 B.n439 585
R244 B.n438 B.n175 585
R245 B.n437 B.n436 585
R246 B.n434 B.n176 585
R247 B.n432 B.n431 585
R248 B.n430 B.n177 585
R249 B.n429 B.n428 585
R250 B.n426 B.n178 585
R251 B.n424 B.n423 585
R252 B.n422 B.n179 585
R253 B.n421 B.n420 585
R254 B.n418 B.n180 585
R255 B.n416 B.n415 585
R256 B.n414 B.n181 585
R257 B.n413 B.n412 585
R258 B.n410 B.n182 585
R259 B.n408 B.n407 585
R260 B.n406 B.n183 585
R261 B.n405 B.n404 585
R262 B.n402 B.n184 585
R263 B.n400 B.n399 585
R264 B.n398 B.n185 585
R265 B.n397 B.n396 585
R266 B.n394 B.n186 585
R267 B.n392 B.n391 585
R268 B.n390 B.n187 585
R269 B.n389 B.n388 585
R270 B.n386 B.n188 585
R271 B.n384 B.n383 585
R272 B.n382 B.n189 585
R273 B.n381 B.n380 585
R274 B.n378 B.n190 585
R275 B.n376 B.n375 585
R276 B.n374 B.n191 585
R277 B.n373 B.n372 585
R278 B.n370 B.n192 585
R279 B.n368 B.n367 585
R280 B.n366 B.n193 585
R281 B.n365 B.n364 585
R282 B.n362 B.n194 585
R283 B.n360 B.n359 585
R284 B.n357 B.n195 585
R285 B.n356 B.n355 585
R286 B.n353 B.n198 585
R287 B.n351 B.n350 585
R288 B.n349 B.n199 585
R289 B.n348 B.n347 585
R290 B.n345 B.n200 585
R291 B.n343 B.n342 585
R292 B.n341 B.n201 585
R293 B.n339 B.n338 585
R294 B.n336 B.n204 585
R295 B.n334 B.n333 585
R296 B.n332 B.n205 585
R297 B.n331 B.n330 585
R298 B.n328 B.n206 585
R299 B.n326 B.n325 585
R300 B.n324 B.n207 585
R301 B.n323 B.n322 585
R302 B.n320 B.n208 585
R303 B.n318 B.n317 585
R304 B.n316 B.n209 585
R305 B.n315 B.n314 585
R306 B.n312 B.n210 585
R307 B.n310 B.n309 585
R308 B.n308 B.n211 585
R309 B.n307 B.n306 585
R310 B.n304 B.n212 585
R311 B.n302 B.n301 585
R312 B.n300 B.n213 585
R313 B.n299 B.n298 585
R314 B.n296 B.n214 585
R315 B.n294 B.n293 585
R316 B.n292 B.n215 585
R317 B.n291 B.n290 585
R318 B.n288 B.n216 585
R319 B.n286 B.n285 585
R320 B.n284 B.n217 585
R321 B.n283 B.n282 585
R322 B.n280 B.n218 585
R323 B.n278 B.n277 585
R324 B.n276 B.n219 585
R325 B.n275 B.n274 585
R326 B.n272 B.n220 585
R327 B.n270 B.n269 585
R328 B.n268 B.n221 585
R329 B.n267 B.n266 585
R330 B.n264 B.n222 585
R331 B.n262 B.n261 585
R332 B.n260 B.n223 585
R333 B.n259 B.n258 585
R334 B.n256 B.n224 585
R335 B.n254 B.n253 585
R336 B.n252 B.n225 585
R337 B.n251 B.n250 585
R338 B.n248 B.n226 585
R339 B.n246 B.n245 585
R340 B.n244 B.n227 585
R341 B.n243 B.n242 585
R342 B.n240 B.n228 585
R343 B.n238 B.n237 585
R344 B.n236 B.n229 585
R345 B.n235 B.n234 585
R346 B.n232 B.n230 585
R347 B.n165 B.n164 585
R348 B.n469 B.n468 585
R349 B.n470 B.n469 585
R350 B.n161 B.n160 585
R351 B.n162 B.n161 585
R352 B.n478 B.n477 585
R353 B.n477 B.n476 585
R354 B.n479 B.n159 585
R355 B.n159 B.n158 585
R356 B.n481 B.n480 585
R357 B.n482 B.n481 585
R358 B.n153 B.n152 585
R359 B.n154 B.n153 585
R360 B.n490 B.n489 585
R361 B.n489 B.n488 585
R362 B.n491 B.n151 585
R363 B.n151 B.n150 585
R364 B.n493 B.n492 585
R365 B.n494 B.n493 585
R366 B.n145 B.n144 585
R367 B.n146 B.n145 585
R368 B.n502 B.n501 585
R369 B.n501 B.n500 585
R370 B.n503 B.n143 585
R371 B.n143 B.n142 585
R372 B.n505 B.n504 585
R373 B.n506 B.n505 585
R374 B.n137 B.n136 585
R375 B.n138 B.n137 585
R376 B.n514 B.n513 585
R377 B.n513 B.n512 585
R378 B.n515 B.n135 585
R379 B.n135 B.n134 585
R380 B.n517 B.n516 585
R381 B.n518 B.n517 585
R382 B.n129 B.n128 585
R383 B.n130 B.n129 585
R384 B.n526 B.n525 585
R385 B.n525 B.n524 585
R386 B.n527 B.n127 585
R387 B.n127 B.n126 585
R388 B.n529 B.n528 585
R389 B.n530 B.n529 585
R390 B.n121 B.n120 585
R391 B.n122 B.n121 585
R392 B.n539 B.n538 585
R393 B.n538 B.n537 585
R394 B.n540 B.n119 585
R395 B.n119 B.n118 585
R396 B.n542 B.n541 585
R397 B.n543 B.n542 585
R398 B.n3 B.n0 585
R399 B.n4 B.n3 585
R400 B.n871 B.n1 585
R401 B.n872 B.n871 585
R402 B.n870 B.n869 585
R403 B.n870 B.n8 585
R404 B.n868 B.n9 585
R405 B.n12 B.n9 585
R406 B.n867 B.n866 585
R407 B.n866 B.n865 585
R408 B.n11 B.n10 585
R409 B.n864 B.n11 585
R410 B.n862 B.n861 585
R411 B.n863 B.n862 585
R412 B.n860 B.n17 585
R413 B.n17 B.n16 585
R414 B.n859 B.n858 585
R415 B.n858 B.n857 585
R416 B.n19 B.n18 585
R417 B.n856 B.n19 585
R418 B.n854 B.n853 585
R419 B.n855 B.n854 585
R420 B.n852 B.n24 585
R421 B.n24 B.n23 585
R422 B.n851 B.n850 585
R423 B.n850 B.n849 585
R424 B.n26 B.n25 585
R425 B.n848 B.n26 585
R426 B.n846 B.n845 585
R427 B.n847 B.n846 585
R428 B.n844 B.n31 585
R429 B.n31 B.n30 585
R430 B.n843 B.n842 585
R431 B.n842 B.n841 585
R432 B.n33 B.n32 585
R433 B.n840 B.n33 585
R434 B.n838 B.n837 585
R435 B.n839 B.n838 585
R436 B.n836 B.n38 585
R437 B.n38 B.n37 585
R438 B.n835 B.n834 585
R439 B.n834 B.n833 585
R440 B.n40 B.n39 585
R441 B.n832 B.n40 585
R442 B.n830 B.n829 585
R443 B.n831 B.n830 585
R444 B.n828 B.n45 585
R445 B.n45 B.n44 585
R446 B.n827 B.n826 585
R447 B.n826 B.n825 585
R448 B.n47 B.n46 585
R449 B.n824 B.n47 585
R450 B.n822 B.n821 585
R451 B.n823 B.n822 585
R452 B.n875 B.n874 585
R453 B.n873 B.n2 585
R454 B.n822 B.n52 506.916
R455 B.n583 B.n50 506.916
R456 B.n471 B.n165 506.916
R457 B.n469 B.n167 506.916
R458 B.n81 B.t6 352.021
R459 B.n88 B.t13 352.021
R460 B.n202 B.t10 352.021
R461 B.n196 B.t2 352.021
R462 B.n584 B.n51 256.663
R463 B.n590 B.n51 256.663
R464 B.n592 B.n51 256.663
R465 B.n598 B.n51 256.663
R466 B.n600 B.n51 256.663
R467 B.n606 B.n51 256.663
R468 B.n608 B.n51 256.663
R469 B.n614 B.n51 256.663
R470 B.n616 B.n51 256.663
R471 B.n622 B.n51 256.663
R472 B.n624 B.n51 256.663
R473 B.n630 B.n51 256.663
R474 B.n632 B.n51 256.663
R475 B.n638 B.n51 256.663
R476 B.n640 B.n51 256.663
R477 B.n646 B.n51 256.663
R478 B.n648 B.n51 256.663
R479 B.n654 B.n51 256.663
R480 B.n656 B.n51 256.663
R481 B.n662 B.n51 256.663
R482 B.n664 B.n51 256.663
R483 B.n670 B.n51 256.663
R484 B.n672 B.n51 256.663
R485 B.n678 B.n51 256.663
R486 B.n680 B.n51 256.663
R487 B.n686 B.n51 256.663
R488 B.n688 B.n51 256.663
R489 B.n695 B.n51 256.663
R490 B.n697 B.n51 256.663
R491 B.n703 B.n51 256.663
R492 B.n705 B.n51 256.663
R493 B.n711 B.n51 256.663
R494 B.n713 B.n51 256.663
R495 B.n719 B.n51 256.663
R496 B.n721 B.n51 256.663
R497 B.n727 B.n51 256.663
R498 B.n729 B.n51 256.663
R499 B.n735 B.n51 256.663
R500 B.n737 B.n51 256.663
R501 B.n743 B.n51 256.663
R502 B.n745 B.n51 256.663
R503 B.n751 B.n51 256.663
R504 B.n753 B.n51 256.663
R505 B.n759 B.n51 256.663
R506 B.n761 B.n51 256.663
R507 B.n767 B.n51 256.663
R508 B.n769 B.n51 256.663
R509 B.n775 B.n51 256.663
R510 B.n777 B.n51 256.663
R511 B.n783 B.n51 256.663
R512 B.n785 B.n51 256.663
R513 B.n791 B.n51 256.663
R514 B.n793 B.n51 256.663
R515 B.n799 B.n51 256.663
R516 B.n801 B.n51 256.663
R517 B.n807 B.n51 256.663
R518 B.n809 B.n51 256.663
R519 B.n815 B.n51 256.663
R520 B.n817 B.n51 256.663
R521 B.n464 B.n166 256.663
R522 B.n169 B.n166 256.663
R523 B.n457 B.n166 256.663
R524 B.n451 B.n166 256.663
R525 B.n449 B.n166 256.663
R526 B.n443 B.n166 256.663
R527 B.n441 B.n166 256.663
R528 B.n435 B.n166 256.663
R529 B.n433 B.n166 256.663
R530 B.n427 B.n166 256.663
R531 B.n425 B.n166 256.663
R532 B.n419 B.n166 256.663
R533 B.n417 B.n166 256.663
R534 B.n411 B.n166 256.663
R535 B.n409 B.n166 256.663
R536 B.n403 B.n166 256.663
R537 B.n401 B.n166 256.663
R538 B.n395 B.n166 256.663
R539 B.n393 B.n166 256.663
R540 B.n387 B.n166 256.663
R541 B.n385 B.n166 256.663
R542 B.n379 B.n166 256.663
R543 B.n377 B.n166 256.663
R544 B.n371 B.n166 256.663
R545 B.n369 B.n166 256.663
R546 B.n363 B.n166 256.663
R547 B.n361 B.n166 256.663
R548 B.n354 B.n166 256.663
R549 B.n352 B.n166 256.663
R550 B.n346 B.n166 256.663
R551 B.n344 B.n166 256.663
R552 B.n337 B.n166 256.663
R553 B.n335 B.n166 256.663
R554 B.n329 B.n166 256.663
R555 B.n327 B.n166 256.663
R556 B.n321 B.n166 256.663
R557 B.n319 B.n166 256.663
R558 B.n313 B.n166 256.663
R559 B.n311 B.n166 256.663
R560 B.n305 B.n166 256.663
R561 B.n303 B.n166 256.663
R562 B.n297 B.n166 256.663
R563 B.n295 B.n166 256.663
R564 B.n289 B.n166 256.663
R565 B.n287 B.n166 256.663
R566 B.n281 B.n166 256.663
R567 B.n279 B.n166 256.663
R568 B.n273 B.n166 256.663
R569 B.n271 B.n166 256.663
R570 B.n265 B.n166 256.663
R571 B.n263 B.n166 256.663
R572 B.n257 B.n166 256.663
R573 B.n255 B.n166 256.663
R574 B.n249 B.n166 256.663
R575 B.n247 B.n166 256.663
R576 B.n241 B.n166 256.663
R577 B.n239 B.n166 256.663
R578 B.n233 B.n166 256.663
R579 B.n231 B.n166 256.663
R580 B.n877 B.n876 256.663
R581 B.n818 B.n816 163.367
R582 B.n814 B.n54 163.367
R583 B.n810 B.n808 163.367
R584 B.n806 B.n56 163.367
R585 B.n802 B.n800 163.367
R586 B.n798 B.n58 163.367
R587 B.n794 B.n792 163.367
R588 B.n790 B.n60 163.367
R589 B.n786 B.n784 163.367
R590 B.n782 B.n62 163.367
R591 B.n778 B.n776 163.367
R592 B.n774 B.n64 163.367
R593 B.n770 B.n768 163.367
R594 B.n766 B.n66 163.367
R595 B.n762 B.n760 163.367
R596 B.n758 B.n68 163.367
R597 B.n754 B.n752 163.367
R598 B.n750 B.n70 163.367
R599 B.n746 B.n744 163.367
R600 B.n742 B.n72 163.367
R601 B.n738 B.n736 163.367
R602 B.n734 B.n74 163.367
R603 B.n730 B.n728 163.367
R604 B.n726 B.n76 163.367
R605 B.n722 B.n720 163.367
R606 B.n718 B.n78 163.367
R607 B.n714 B.n712 163.367
R608 B.n710 B.n80 163.367
R609 B.n706 B.n704 163.367
R610 B.n702 B.n85 163.367
R611 B.n698 B.n696 163.367
R612 B.n694 B.n87 163.367
R613 B.n689 B.n687 163.367
R614 B.n685 B.n91 163.367
R615 B.n681 B.n679 163.367
R616 B.n677 B.n93 163.367
R617 B.n673 B.n671 163.367
R618 B.n669 B.n95 163.367
R619 B.n665 B.n663 163.367
R620 B.n661 B.n97 163.367
R621 B.n657 B.n655 163.367
R622 B.n653 B.n99 163.367
R623 B.n649 B.n647 163.367
R624 B.n645 B.n101 163.367
R625 B.n641 B.n639 163.367
R626 B.n637 B.n103 163.367
R627 B.n633 B.n631 163.367
R628 B.n629 B.n105 163.367
R629 B.n625 B.n623 163.367
R630 B.n621 B.n107 163.367
R631 B.n617 B.n615 163.367
R632 B.n613 B.n109 163.367
R633 B.n609 B.n607 163.367
R634 B.n605 B.n111 163.367
R635 B.n601 B.n599 163.367
R636 B.n597 B.n113 163.367
R637 B.n593 B.n591 163.367
R638 B.n589 B.n115 163.367
R639 B.n585 B.n583 163.367
R640 B.n471 B.n163 163.367
R641 B.n475 B.n163 163.367
R642 B.n475 B.n157 163.367
R643 B.n483 B.n157 163.367
R644 B.n483 B.n155 163.367
R645 B.n487 B.n155 163.367
R646 B.n487 B.n149 163.367
R647 B.n495 B.n149 163.367
R648 B.n495 B.n147 163.367
R649 B.n499 B.n147 163.367
R650 B.n499 B.n141 163.367
R651 B.n507 B.n141 163.367
R652 B.n507 B.n139 163.367
R653 B.n511 B.n139 163.367
R654 B.n511 B.n133 163.367
R655 B.n519 B.n133 163.367
R656 B.n519 B.n131 163.367
R657 B.n523 B.n131 163.367
R658 B.n523 B.n125 163.367
R659 B.n531 B.n125 163.367
R660 B.n531 B.n123 163.367
R661 B.n536 B.n123 163.367
R662 B.n536 B.n117 163.367
R663 B.n544 B.n117 163.367
R664 B.n545 B.n544 163.367
R665 B.n545 B.n5 163.367
R666 B.n6 B.n5 163.367
R667 B.n7 B.n6 163.367
R668 B.n551 B.n7 163.367
R669 B.n552 B.n551 163.367
R670 B.n552 B.n13 163.367
R671 B.n14 B.n13 163.367
R672 B.n15 B.n14 163.367
R673 B.n557 B.n15 163.367
R674 B.n557 B.n20 163.367
R675 B.n21 B.n20 163.367
R676 B.n22 B.n21 163.367
R677 B.n562 B.n22 163.367
R678 B.n562 B.n27 163.367
R679 B.n28 B.n27 163.367
R680 B.n29 B.n28 163.367
R681 B.n567 B.n29 163.367
R682 B.n567 B.n34 163.367
R683 B.n35 B.n34 163.367
R684 B.n36 B.n35 163.367
R685 B.n572 B.n36 163.367
R686 B.n572 B.n41 163.367
R687 B.n42 B.n41 163.367
R688 B.n43 B.n42 163.367
R689 B.n577 B.n43 163.367
R690 B.n577 B.n48 163.367
R691 B.n49 B.n48 163.367
R692 B.n50 B.n49 163.367
R693 B.n465 B.n463 163.367
R694 B.n463 B.n462 163.367
R695 B.n459 B.n458 163.367
R696 B.n456 B.n171 163.367
R697 B.n452 B.n450 163.367
R698 B.n448 B.n173 163.367
R699 B.n444 B.n442 163.367
R700 B.n440 B.n175 163.367
R701 B.n436 B.n434 163.367
R702 B.n432 B.n177 163.367
R703 B.n428 B.n426 163.367
R704 B.n424 B.n179 163.367
R705 B.n420 B.n418 163.367
R706 B.n416 B.n181 163.367
R707 B.n412 B.n410 163.367
R708 B.n408 B.n183 163.367
R709 B.n404 B.n402 163.367
R710 B.n400 B.n185 163.367
R711 B.n396 B.n394 163.367
R712 B.n392 B.n187 163.367
R713 B.n388 B.n386 163.367
R714 B.n384 B.n189 163.367
R715 B.n380 B.n378 163.367
R716 B.n376 B.n191 163.367
R717 B.n372 B.n370 163.367
R718 B.n368 B.n193 163.367
R719 B.n364 B.n362 163.367
R720 B.n360 B.n195 163.367
R721 B.n355 B.n353 163.367
R722 B.n351 B.n199 163.367
R723 B.n347 B.n345 163.367
R724 B.n343 B.n201 163.367
R725 B.n338 B.n336 163.367
R726 B.n334 B.n205 163.367
R727 B.n330 B.n328 163.367
R728 B.n326 B.n207 163.367
R729 B.n322 B.n320 163.367
R730 B.n318 B.n209 163.367
R731 B.n314 B.n312 163.367
R732 B.n310 B.n211 163.367
R733 B.n306 B.n304 163.367
R734 B.n302 B.n213 163.367
R735 B.n298 B.n296 163.367
R736 B.n294 B.n215 163.367
R737 B.n290 B.n288 163.367
R738 B.n286 B.n217 163.367
R739 B.n282 B.n280 163.367
R740 B.n278 B.n219 163.367
R741 B.n274 B.n272 163.367
R742 B.n270 B.n221 163.367
R743 B.n266 B.n264 163.367
R744 B.n262 B.n223 163.367
R745 B.n258 B.n256 163.367
R746 B.n254 B.n225 163.367
R747 B.n250 B.n248 163.367
R748 B.n246 B.n227 163.367
R749 B.n242 B.n240 163.367
R750 B.n238 B.n229 163.367
R751 B.n234 B.n232 163.367
R752 B.n469 B.n161 163.367
R753 B.n477 B.n161 163.367
R754 B.n477 B.n159 163.367
R755 B.n481 B.n159 163.367
R756 B.n481 B.n153 163.367
R757 B.n489 B.n153 163.367
R758 B.n489 B.n151 163.367
R759 B.n493 B.n151 163.367
R760 B.n493 B.n145 163.367
R761 B.n501 B.n145 163.367
R762 B.n501 B.n143 163.367
R763 B.n505 B.n143 163.367
R764 B.n505 B.n137 163.367
R765 B.n513 B.n137 163.367
R766 B.n513 B.n135 163.367
R767 B.n517 B.n135 163.367
R768 B.n517 B.n129 163.367
R769 B.n525 B.n129 163.367
R770 B.n525 B.n127 163.367
R771 B.n529 B.n127 163.367
R772 B.n529 B.n121 163.367
R773 B.n538 B.n121 163.367
R774 B.n538 B.n119 163.367
R775 B.n542 B.n119 163.367
R776 B.n542 B.n3 163.367
R777 B.n875 B.n3 163.367
R778 B.n871 B.n2 163.367
R779 B.n871 B.n870 163.367
R780 B.n870 B.n9 163.367
R781 B.n866 B.n9 163.367
R782 B.n866 B.n11 163.367
R783 B.n862 B.n11 163.367
R784 B.n862 B.n17 163.367
R785 B.n858 B.n17 163.367
R786 B.n858 B.n19 163.367
R787 B.n854 B.n19 163.367
R788 B.n854 B.n24 163.367
R789 B.n850 B.n24 163.367
R790 B.n850 B.n26 163.367
R791 B.n846 B.n26 163.367
R792 B.n846 B.n31 163.367
R793 B.n842 B.n31 163.367
R794 B.n842 B.n33 163.367
R795 B.n838 B.n33 163.367
R796 B.n838 B.n38 163.367
R797 B.n834 B.n38 163.367
R798 B.n834 B.n40 163.367
R799 B.n830 B.n40 163.367
R800 B.n830 B.n45 163.367
R801 B.n826 B.n45 163.367
R802 B.n826 B.n47 163.367
R803 B.n822 B.n47 163.367
R804 B.n88 B.t14 131.345
R805 B.n202 B.t12 131.345
R806 B.n81 B.t8 131.323
R807 B.n196 B.t5 131.323
R808 B.n817 B.n52 71.676
R809 B.n816 B.n815 71.676
R810 B.n809 B.n54 71.676
R811 B.n808 B.n807 71.676
R812 B.n801 B.n56 71.676
R813 B.n800 B.n799 71.676
R814 B.n793 B.n58 71.676
R815 B.n792 B.n791 71.676
R816 B.n785 B.n60 71.676
R817 B.n784 B.n783 71.676
R818 B.n777 B.n62 71.676
R819 B.n776 B.n775 71.676
R820 B.n769 B.n64 71.676
R821 B.n768 B.n767 71.676
R822 B.n761 B.n66 71.676
R823 B.n760 B.n759 71.676
R824 B.n753 B.n68 71.676
R825 B.n752 B.n751 71.676
R826 B.n745 B.n70 71.676
R827 B.n744 B.n743 71.676
R828 B.n737 B.n72 71.676
R829 B.n736 B.n735 71.676
R830 B.n729 B.n74 71.676
R831 B.n728 B.n727 71.676
R832 B.n721 B.n76 71.676
R833 B.n720 B.n719 71.676
R834 B.n713 B.n78 71.676
R835 B.n712 B.n711 71.676
R836 B.n705 B.n80 71.676
R837 B.n704 B.n703 71.676
R838 B.n697 B.n85 71.676
R839 B.n696 B.n695 71.676
R840 B.n688 B.n87 71.676
R841 B.n687 B.n686 71.676
R842 B.n680 B.n91 71.676
R843 B.n679 B.n678 71.676
R844 B.n672 B.n93 71.676
R845 B.n671 B.n670 71.676
R846 B.n664 B.n95 71.676
R847 B.n663 B.n662 71.676
R848 B.n656 B.n97 71.676
R849 B.n655 B.n654 71.676
R850 B.n648 B.n99 71.676
R851 B.n647 B.n646 71.676
R852 B.n640 B.n101 71.676
R853 B.n639 B.n638 71.676
R854 B.n632 B.n103 71.676
R855 B.n631 B.n630 71.676
R856 B.n624 B.n105 71.676
R857 B.n623 B.n622 71.676
R858 B.n616 B.n107 71.676
R859 B.n615 B.n614 71.676
R860 B.n608 B.n109 71.676
R861 B.n607 B.n606 71.676
R862 B.n600 B.n111 71.676
R863 B.n599 B.n598 71.676
R864 B.n592 B.n113 71.676
R865 B.n591 B.n590 71.676
R866 B.n584 B.n115 71.676
R867 B.n585 B.n584 71.676
R868 B.n590 B.n589 71.676
R869 B.n593 B.n592 71.676
R870 B.n598 B.n597 71.676
R871 B.n601 B.n600 71.676
R872 B.n606 B.n605 71.676
R873 B.n609 B.n608 71.676
R874 B.n614 B.n613 71.676
R875 B.n617 B.n616 71.676
R876 B.n622 B.n621 71.676
R877 B.n625 B.n624 71.676
R878 B.n630 B.n629 71.676
R879 B.n633 B.n632 71.676
R880 B.n638 B.n637 71.676
R881 B.n641 B.n640 71.676
R882 B.n646 B.n645 71.676
R883 B.n649 B.n648 71.676
R884 B.n654 B.n653 71.676
R885 B.n657 B.n656 71.676
R886 B.n662 B.n661 71.676
R887 B.n665 B.n664 71.676
R888 B.n670 B.n669 71.676
R889 B.n673 B.n672 71.676
R890 B.n678 B.n677 71.676
R891 B.n681 B.n680 71.676
R892 B.n686 B.n685 71.676
R893 B.n689 B.n688 71.676
R894 B.n695 B.n694 71.676
R895 B.n698 B.n697 71.676
R896 B.n703 B.n702 71.676
R897 B.n706 B.n705 71.676
R898 B.n711 B.n710 71.676
R899 B.n714 B.n713 71.676
R900 B.n719 B.n718 71.676
R901 B.n722 B.n721 71.676
R902 B.n727 B.n726 71.676
R903 B.n730 B.n729 71.676
R904 B.n735 B.n734 71.676
R905 B.n738 B.n737 71.676
R906 B.n743 B.n742 71.676
R907 B.n746 B.n745 71.676
R908 B.n751 B.n750 71.676
R909 B.n754 B.n753 71.676
R910 B.n759 B.n758 71.676
R911 B.n762 B.n761 71.676
R912 B.n767 B.n766 71.676
R913 B.n770 B.n769 71.676
R914 B.n775 B.n774 71.676
R915 B.n778 B.n777 71.676
R916 B.n783 B.n782 71.676
R917 B.n786 B.n785 71.676
R918 B.n791 B.n790 71.676
R919 B.n794 B.n793 71.676
R920 B.n799 B.n798 71.676
R921 B.n802 B.n801 71.676
R922 B.n807 B.n806 71.676
R923 B.n810 B.n809 71.676
R924 B.n815 B.n814 71.676
R925 B.n818 B.n817 71.676
R926 B.n464 B.n167 71.676
R927 B.n462 B.n169 71.676
R928 B.n458 B.n457 71.676
R929 B.n451 B.n171 71.676
R930 B.n450 B.n449 71.676
R931 B.n443 B.n173 71.676
R932 B.n442 B.n441 71.676
R933 B.n435 B.n175 71.676
R934 B.n434 B.n433 71.676
R935 B.n427 B.n177 71.676
R936 B.n426 B.n425 71.676
R937 B.n419 B.n179 71.676
R938 B.n418 B.n417 71.676
R939 B.n411 B.n181 71.676
R940 B.n410 B.n409 71.676
R941 B.n403 B.n183 71.676
R942 B.n402 B.n401 71.676
R943 B.n395 B.n185 71.676
R944 B.n394 B.n393 71.676
R945 B.n387 B.n187 71.676
R946 B.n386 B.n385 71.676
R947 B.n379 B.n189 71.676
R948 B.n378 B.n377 71.676
R949 B.n371 B.n191 71.676
R950 B.n370 B.n369 71.676
R951 B.n363 B.n193 71.676
R952 B.n362 B.n361 71.676
R953 B.n354 B.n195 71.676
R954 B.n353 B.n352 71.676
R955 B.n346 B.n199 71.676
R956 B.n345 B.n344 71.676
R957 B.n337 B.n201 71.676
R958 B.n336 B.n335 71.676
R959 B.n329 B.n205 71.676
R960 B.n328 B.n327 71.676
R961 B.n321 B.n207 71.676
R962 B.n320 B.n319 71.676
R963 B.n313 B.n209 71.676
R964 B.n312 B.n311 71.676
R965 B.n305 B.n211 71.676
R966 B.n304 B.n303 71.676
R967 B.n297 B.n213 71.676
R968 B.n296 B.n295 71.676
R969 B.n289 B.n215 71.676
R970 B.n288 B.n287 71.676
R971 B.n281 B.n217 71.676
R972 B.n280 B.n279 71.676
R973 B.n273 B.n219 71.676
R974 B.n272 B.n271 71.676
R975 B.n265 B.n221 71.676
R976 B.n264 B.n263 71.676
R977 B.n257 B.n223 71.676
R978 B.n256 B.n255 71.676
R979 B.n249 B.n225 71.676
R980 B.n248 B.n247 71.676
R981 B.n241 B.n227 71.676
R982 B.n240 B.n239 71.676
R983 B.n233 B.n229 71.676
R984 B.n232 B.n231 71.676
R985 B.n465 B.n464 71.676
R986 B.n459 B.n169 71.676
R987 B.n457 B.n456 71.676
R988 B.n452 B.n451 71.676
R989 B.n449 B.n448 71.676
R990 B.n444 B.n443 71.676
R991 B.n441 B.n440 71.676
R992 B.n436 B.n435 71.676
R993 B.n433 B.n432 71.676
R994 B.n428 B.n427 71.676
R995 B.n425 B.n424 71.676
R996 B.n420 B.n419 71.676
R997 B.n417 B.n416 71.676
R998 B.n412 B.n411 71.676
R999 B.n409 B.n408 71.676
R1000 B.n404 B.n403 71.676
R1001 B.n401 B.n400 71.676
R1002 B.n396 B.n395 71.676
R1003 B.n393 B.n392 71.676
R1004 B.n388 B.n387 71.676
R1005 B.n385 B.n384 71.676
R1006 B.n380 B.n379 71.676
R1007 B.n377 B.n376 71.676
R1008 B.n372 B.n371 71.676
R1009 B.n369 B.n368 71.676
R1010 B.n364 B.n363 71.676
R1011 B.n361 B.n360 71.676
R1012 B.n355 B.n354 71.676
R1013 B.n352 B.n351 71.676
R1014 B.n347 B.n346 71.676
R1015 B.n344 B.n343 71.676
R1016 B.n338 B.n337 71.676
R1017 B.n335 B.n334 71.676
R1018 B.n330 B.n329 71.676
R1019 B.n327 B.n326 71.676
R1020 B.n322 B.n321 71.676
R1021 B.n319 B.n318 71.676
R1022 B.n314 B.n313 71.676
R1023 B.n311 B.n310 71.676
R1024 B.n306 B.n305 71.676
R1025 B.n303 B.n302 71.676
R1026 B.n298 B.n297 71.676
R1027 B.n295 B.n294 71.676
R1028 B.n290 B.n289 71.676
R1029 B.n287 B.n286 71.676
R1030 B.n282 B.n281 71.676
R1031 B.n279 B.n278 71.676
R1032 B.n274 B.n273 71.676
R1033 B.n271 B.n270 71.676
R1034 B.n266 B.n265 71.676
R1035 B.n263 B.n262 71.676
R1036 B.n258 B.n257 71.676
R1037 B.n255 B.n254 71.676
R1038 B.n250 B.n249 71.676
R1039 B.n247 B.n246 71.676
R1040 B.n242 B.n241 71.676
R1041 B.n239 B.n238 71.676
R1042 B.n234 B.n233 71.676
R1043 B.n231 B.n165 71.676
R1044 B.n876 B.n875 71.676
R1045 B.n876 B.n2 71.676
R1046 B.n89 B.t15 71.2237
R1047 B.n203 B.t11 71.2237
R1048 B.n82 B.t9 71.202
R1049 B.n197 B.t4 71.202
R1050 B.n82 B.n81 60.1217
R1051 B.n89 B.n88 60.1217
R1052 B.n203 B.n202 60.1217
R1053 B.n197 B.n196 60.1217
R1054 B.n83 B.n82 59.5399
R1055 B.n692 B.n89 59.5399
R1056 B.n340 B.n203 59.5399
R1057 B.n358 B.n197 59.5399
R1058 B.n470 B.n166 57.0319
R1059 B.n823 B.n51 57.0319
R1060 B.n470 B.n162 34.3203
R1061 B.n476 B.n162 34.3203
R1062 B.n476 B.n158 34.3203
R1063 B.n482 B.n158 34.3203
R1064 B.n482 B.n154 34.3203
R1065 B.n488 B.n154 34.3203
R1066 B.n488 B.n150 34.3203
R1067 B.n494 B.n150 34.3203
R1068 B.n500 B.n146 34.3203
R1069 B.n500 B.n142 34.3203
R1070 B.n506 B.n142 34.3203
R1071 B.n506 B.n138 34.3203
R1072 B.n512 B.n138 34.3203
R1073 B.n512 B.n134 34.3203
R1074 B.n518 B.n134 34.3203
R1075 B.n518 B.n130 34.3203
R1076 B.n524 B.n130 34.3203
R1077 B.n524 B.n126 34.3203
R1078 B.n530 B.n126 34.3203
R1079 B.n537 B.n122 34.3203
R1080 B.n537 B.n118 34.3203
R1081 B.n543 B.n118 34.3203
R1082 B.n543 B.n4 34.3203
R1083 B.n874 B.n4 34.3203
R1084 B.n874 B.n873 34.3203
R1085 B.n873 B.n872 34.3203
R1086 B.n872 B.n8 34.3203
R1087 B.n12 B.n8 34.3203
R1088 B.n865 B.n12 34.3203
R1089 B.n865 B.n864 34.3203
R1090 B.n863 B.n16 34.3203
R1091 B.n857 B.n16 34.3203
R1092 B.n857 B.n856 34.3203
R1093 B.n856 B.n855 34.3203
R1094 B.n855 B.n23 34.3203
R1095 B.n849 B.n23 34.3203
R1096 B.n849 B.n848 34.3203
R1097 B.n848 B.n847 34.3203
R1098 B.n847 B.n30 34.3203
R1099 B.n841 B.n30 34.3203
R1100 B.n841 B.n840 34.3203
R1101 B.n839 B.n37 34.3203
R1102 B.n833 B.n37 34.3203
R1103 B.n833 B.n832 34.3203
R1104 B.n832 B.n831 34.3203
R1105 B.n831 B.n44 34.3203
R1106 B.n825 B.n44 34.3203
R1107 B.n825 B.n824 34.3203
R1108 B.n824 B.n823 34.3203
R1109 B.t3 B.n146 33.8156
R1110 B.n840 B.t7 33.8156
R1111 B.n468 B.n467 32.9371
R1112 B.n472 B.n164 32.9371
R1113 B.n582 B.n581 32.9371
R1114 B.n821 B.n820 32.9371
R1115 B.t1 B.n122 22.7121
R1116 B.n864 B.t0 22.7121
R1117 B B.n877 18.0485
R1118 B.n530 B.t1 11.6087
R1119 B.t0 B.n863 11.6087
R1120 B.n468 B.n160 10.6151
R1121 B.n478 B.n160 10.6151
R1122 B.n479 B.n478 10.6151
R1123 B.n480 B.n479 10.6151
R1124 B.n480 B.n152 10.6151
R1125 B.n490 B.n152 10.6151
R1126 B.n491 B.n490 10.6151
R1127 B.n492 B.n491 10.6151
R1128 B.n492 B.n144 10.6151
R1129 B.n502 B.n144 10.6151
R1130 B.n503 B.n502 10.6151
R1131 B.n504 B.n503 10.6151
R1132 B.n504 B.n136 10.6151
R1133 B.n514 B.n136 10.6151
R1134 B.n515 B.n514 10.6151
R1135 B.n516 B.n515 10.6151
R1136 B.n516 B.n128 10.6151
R1137 B.n526 B.n128 10.6151
R1138 B.n527 B.n526 10.6151
R1139 B.n528 B.n527 10.6151
R1140 B.n528 B.n120 10.6151
R1141 B.n539 B.n120 10.6151
R1142 B.n540 B.n539 10.6151
R1143 B.n541 B.n540 10.6151
R1144 B.n541 B.n0 10.6151
R1145 B.n467 B.n466 10.6151
R1146 B.n466 B.n168 10.6151
R1147 B.n461 B.n168 10.6151
R1148 B.n461 B.n460 10.6151
R1149 B.n460 B.n170 10.6151
R1150 B.n455 B.n170 10.6151
R1151 B.n455 B.n454 10.6151
R1152 B.n454 B.n453 10.6151
R1153 B.n453 B.n172 10.6151
R1154 B.n447 B.n172 10.6151
R1155 B.n447 B.n446 10.6151
R1156 B.n446 B.n445 10.6151
R1157 B.n445 B.n174 10.6151
R1158 B.n439 B.n174 10.6151
R1159 B.n439 B.n438 10.6151
R1160 B.n438 B.n437 10.6151
R1161 B.n437 B.n176 10.6151
R1162 B.n431 B.n176 10.6151
R1163 B.n431 B.n430 10.6151
R1164 B.n430 B.n429 10.6151
R1165 B.n429 B.n178 10.6151
R1166 B.n423 B.n178 10.6151
R1167 B.n423 B.n422 10.6151
R1168 B.n422 B.n421 10.6151
R1169 B.n421 B.n180 10.6151
R1170 B.n415 B.n180 10.6151
R1171 B.n415 B.n414 10.6151
R1172 B.n414 B.n413 10.6151
R1173 B.n413 B.n182 10.6151
R1174 B.n407 B.n182 10.6151
R1175 B.n407 B.n406 10.6151
R1176 B.n406 B.n405 10.6151
R1177 B.n405 B.n184 10.6151
R1178 B.n399 B.n184 10.6151
R1179 B.n399 B.n398 10.6151
R1180 B.n398 B.n397 10.6151
R1181 B.n397 B.n186 10.6151
R1182 B.n391 B.n186 10.6151
R1183 B.n391 B.n390 10.6151
R1184 B.n390 B.n389 10.6151
R1185 B.n389 B.n188 10.6151
R1186 B.n383 B.n188 10.6151
R1187 B.n383 B.n382 10.6151
R1188 B.n382 B.n381 10.6151
R1189 B.n381 B.n190 10.6151
R1190 B.n375 B.n190 10.6151
R1191 B.n375 B.n374 10.6151
R1192 B.n374 B.n373 10.6151
R1193 B.n373 B.n192 10.6151
R1194 B.n367 B.n192 10.6151
R1195 B.n367 B.n366 10.6151
R1196 B.n366 B.n365 10.6151
R1197 B.n365 B.n194 10.6151
R1198 B.n359 B.n194 10.6151
R1199 B.n357 B.n356 10.6151
R1200 B.n356 B.n198 10.6151
R1201 B.n350 B.n198 10.6151
R1202 B.n350 B.n349 10.6151
R1203 B.n349 B.n348 10.6151
R1204 B.n348 B.n200 10.6151
R1205 B.n342 B.n200 10.6151
R1206 B.n342 B.n341 10.6151
R1207 B.n339 B.n204 10.6151
R1208 B.n333 B.n204 10.6151
R1209 B.n333 B.n332 10.6151
R1210 B.n332 B.n331 10.6151
R1211 B.n331 B.n206 10.6151
R1212 B.n325 B.n206 10.6151
R1213 B.n325 B.n324 10.6151
R1214 B.n324 B.n323 10.6151
R1215 B.n323 B.n208 10.6151
R1216 B.n317 B.n208 10.6151
R1217 B.n317 B.n316 10.6151
R1218 B.n316 B.n315 10.6151
R1219 B.n315 B.n210 10.6151
R1220 B.n309 B.n210 10.6151
R1221 B.n309 B.n308 10.6151
R1222 B.n308 B.n307 10.6151
R1223 B.n307 B.n212 10.6151
R1224 B.n301 B.n212 10.6151
R1225 B.n301 B.n300 10.6151
R1226 B.n300 B.n299 10.6151
R1227 B.n299 B.n214 10.6151
R1228 B.n293 B.n214 10.6151
R1229 B.n293 B.n292 10.6151
R1230 B.n292 B.n291 10.6151
R1231 B.n291 B.n216 10.6151
R1232 B.n285 B.n216 10.6151
R1233 B.n285 B.n284 10.6151
R1234 B.n284 B.n283 10.6151
R1235 B.n283 B.n218 10.6151
R1236 B.n277 B.n218 10.6151
R1237 B.n277 B.n276 10.6151
R1238 B.n276 B.n275 10.6151
R1239 B.n275 B.n220 10.6151
R1240 B.n269 B.n220 10.6151
R1241 B.n269 B.n268 10.6151
R1242 B.n268 B.n267 10.6151
R1243 B.n267 B.n222 10.6151
R1244 B.n261 B.n222 10.6151
R1245 B.n261 B.n260 10.6151
R1246 B.n260 B.n259 10.6151
R1247 B.n259 B.n224 10.6151
R1248 B.n253 B.n224 10.6151
R1249 B.n253 B.n252 10.6151
R1250 B.n252 B.n251 10.6151
R1251 B.n251 B.n226 10.6151
R1252 B.n245 B.n226 10.6151
R1253 B.n245 B.n244 10.6151
R1254 B.n244 B.n243 10.6151
R1255 B.n243 B.n228 10.6151
R1256 B.n237 B.n228 10.6151
R1257 B.n237 B.n236 10.6151
R1258 B.n236 B.n235 10.6151
R1259 B.n235 B.n230 10.6151
R1260 B.n230 B.n164 10.6151
R1261 B.n473 B.n472 10.6151
R1262 B.n474 B.n473 10.6151
R1263 B.n474 B.n156 10.6151
R1264 B.n484 B.n156 10.6151
R1265 B.n485 B.n484 10.6151
R1266 B.n486 B.n485 10.6151
R1267 B.n486 B.n148 10.6151
R1268 B.n496 B.n148 10.6151
R1269 B.n497 B.n496 10.6151
R1270 B.n498 B.n497 10.6151
R1271 B.n498 B.n140 10.6151
R1272 B.n508 B.n140 10.6151
R1273 B.n509 B.n508 10.6151
R1274 B.n510 B.n509 10.6151
R1275 B.n510 B.n132 10.6151
R1276 B.n520 B.n132 10.6151
R1277 B.n521 B.n520 10.6151
R1278 B.n522 B.n521 10.6151
R1279 B.n522 B.n124 10.6151
R1280 B.n532 B.n124 10.6151
R1281 B.n533 B.n532 10.6151
R1282 B.n535 B.n533 10.6151
R1283 B.n535 B.n534 10.6151
R1284 B.n534 B.n116 10.6151
R1285 B.n546 B.n116 10.6151
R1286 B.n547 B.n546 10.6151
R1287 B.n548 B.n547 10.6151
R1288 B.n549 B.n548 10.6151
R1289 B.n550 B.n549 10.6151
R1290 B.n553 B.n550 10.6151
R1291 B.n554 B.n553 10.6151
R1292 B.n555 B.n554 10.6151
R1293 B.n556 B.n555 10.6151
R1294 B.n558 B.n556 10.6151
R1295 B.n559 B.n558 10.6151
R1296 B.n560 B.n559 10.6151
R1297 B.n561 B.n560 10.6151
R1298 B.n563 B.n561 10.6151
R1299 B.n564 B.n563 10.6151
R1300 B.n565 B.n564 10.6151
R1301 B.n566 B.n565 10.6151
R1302 B.n568 B.n566 10.6151
R1303 B.n569 B.n568 10.6151
R1304 B.n570 B.n569 10.6151
R1305 B.n571 B.n570 10.6151
R1306 B.n573 B.n571 10.6151
R1307 B.n574 B.n573 10.6151
R1308 B.n575 B.n574 10.6151
R1309 B.n576 B.n575 10.6151
R1310 B.n578 B.n576 10.6151
R1311 B.n579 B.n578 10.6151
R1312 B.n580 B.n579 10.6151
R1313 B.n581 B.n580 10.6151
R1314 B.n869 B.n1 10.6151
R1315 B.n869 B.n868 10.6151
R1316 B.n868 B.n867 10.6151
R1317 B.n867 B.n10 10.6151
R1318 B.n861 B.n10 10.6151
R1319 B.n861 B.n860 10.6151
R1320 B.n860 B.n859 10.6151
R1321 B.n859 B.n18 10.6151
R1322 B.n853 B.n18 10.6151
R1323 B.n853 B.n852 10.6151
R1324 B.n852 B.n851 10.6151
R1325 B.n851 B.n25 10.6151
R1326 B.n845 B.n25 10.6151
R1327 B.n845 B.n844 10.6151
R1328 B.n844 B.n843 10.6151
R1329 B.n843 B.n32 10.6151
R1330 B.n837 B.n32 10.6151
R1331 B.n837 B.n836 10.6151
R1332 B.n836 B.n835 10.6151
R1333 B.n835 B.n39 10.6151
R1334 B.n829 B.n39 10.6151
R1335 B.n829 B.n828 10.6151
R1336 B.n828 B.n827 10.6151
R1337 B.n827 B.n46 10.6151
R1338 B.n821 B.n46 10.6151
R1339 B.n820 B.n819 10.6151
R1340 B.n819 B.n53 10.6151
R1341 B.n813 B.n53 10.6151
R1342 B.n813 B.n812 10.6151
R1343 B.n812 B.n811 10.6151
R1344 B.n811 B.n55 10.6151
R1345 B.n805 B.n55 10.6151
R1346 B.n805 B.n804 10.6151
R1347 B.n804 B.n803 10.6151
R1348 B.n803 B.n57 10.6151
R1349 B.n797 B.n57 10.6151
R1350 B.n797 B.n796 10.6151
R1351 B.n796 B.n795 10.6151
R1352 B.n795 B.n59 10.6151
R1353 B.n789 B.n59 10.6151
R1354 B.n789 B.n788 10.6151
R1355 B.n788 B.n787 10.6151
R1356 B.n787 B.n61 10.6151
R1357 B.n781 B.n61 10.6151
R1358 B.n781 B.n780 10.6151
R1359 B.n780 B.n779 10.6151
R1360 B.n779 B.n63 10.6151
R1361 B.n773 B.n63 10.6151
R1362 B.n773 B.n772 10.6151
R1363 B.n772 B.n771 10.6151
R1364 B.n771 B.n65 10.6151
R1365 B.n765 B.n65 10.6151
R1366 B.n765 B.n764 10.6151
R1367 B.n764 B.n763 10.6151
R1368 B.n763 B.n67 10.6151
R1369 B.n757 B.n67 10.6151
R1370 B.n757 B.n756 10.6151
R1371 B.n756 B.n755 10.6151
R1372 B.n755 B.n69 10.6151
R1373 B.n749 B.n69 10.6151
R1374 B.n749 B.n748 10.6151
R1375 B.n748 B.n747 10.6151
R1376 B.n747 B.n71 10.6151
R1377 B.n741 B.n71 10.6151
R1378 B.n741 B.n740 10.6151
R1379 B.n740 B.n739 10.6151
R1380 B.n739 B.n73 10.6151
R1381 B.n733 B.n73 10.6151
R1382 B.n733 B.n732 10.6151
R1383 B.n732 B.n731 10.6151
R1384 B.n731 B.n75 10.6151
R1385 B.n725 B.n75 10.6151
R1386 B.n725 B.n724 10.6151
R1387 B.n724 B.n723 10.6151
R1388 B.n723 B.n77 10.6151
R1389 B.n717 B.n77 10.6151
R1390 B.n717 B.n716 10.6151
R1391 B.n716 B.n715 10.6151
R1392 B.n715 B.n79 10.6151
R1393 B.n709 B.n708 10.6151
R1394 B.n708 B.n707 10.6151
R1395 B.n707 B.n84 10.6151
R1396 B.n701 B.n84 10.6151
R1397 B.n701 B.n700 10.6151
R1398 B.n700 B.n699 10.6151
R1399 B.n699 B.n86 10.6151
R1400 B.n693 B.n86 10.6151
R1401 B.n691 B.n690 10.6151
R1402 B.n690 B.n90 10.6151
R1403 B.n684 B.n90 10.6151
R1404 B.n684 B.n683 10.6151
R1405 B.n683 B.n682 10.6151
R1406 B.n682 B.n92 10.6151
R1407 B.n676 B.n92 10.6151
R1408 B.n676 B.n675 10.6151
R1409 B.n675 B.n674 10.6151
R1410 B.n674 B.n94 10.6151
R1411 B.n668 B.n94 10.6151
R1412 B.n668 B.n667 10.6151
R1413 B.n667 B.n666 10.6151
R1414 B.n666 B.n96 10.6151
R1415 B.n660 B.n96 10.6151
R1416 B.n660 B.n659 10.6151
R1417 B.n659 B.n658 10.6151
R1418 B.n658 B.n98 10.6151
R1419 B.n652 B.n98 10.6151
R1420 B.n652 B.n651 10.6151
R1421 B.n651 B.n650 10.6151
R1422 B.n650 B.n100 10.6151
R1423 B.n644 B.n100 10.6151
R1424 B.n644 B.n643 10.6151
R1425 B.n643 B.n642 10.6151
R1426 B.n642 B.n102 10.6151
R1427 B.n636 B.n102 10.6151
R1428 B.n636 B.n635 10.6151
R1429 B.n635 B.n634 10.6151
R1430 B.n634 B.n104 10.6151
R1431 B.n628 B.n104 10.6151
R1432 B.n628 B.n627 10.6151
R1433 B.n627 B.n626 10.6151
R1434 B.n626 B.n106 10.6151
R1435 B.n620 B.n106 10.6151
R1436 B.n620 B.n619 10.6151
R1437 B.n619 B.n618 10.6151
R1438 B.n618 B.n108 10.6151
R1439 B.n612 B.n108 10.6151
R1440 B.n612 B.n611 10.6151
R1441 B.n611 B.n610 10.6151
R1442 B.n610 B.n110 10.6151
R1443 B.n604 B.n110 10.6151
R1444 B.n604 B.n603 10.6151
R1445 B.n603 B.n602 10.6151
R1446 B.n602 B.n112 10.6151
R1447 B.n596 B.n112 10.6151
R1448 B.n596 B.n595 10.6151
R1449 B.n595 B.n594 10.6151
R1450 B.n594 B.n114 10.6151
R1451 B.n588 B.n114 10.6151
R1452 B.n588 B.n587 10.6151
R1453 B.n587 B.n586 10.6151
R1454 B.n586 B.n582 10.6151
R1455 B.n877 B.n0 8.11757
R1456 B.n877 B.n1 8.11757
R1457 B.n358 B.n357 6.5566
R1458 B.n341 B.n340 6.5566
R1459 B.n709 B.n83 6.5566
R1460 B.n693 B.n692 6.5566
R1461 B.n359 B.n358 4.05904
R1462 B.n340 B.n339 4.05904
R1463 B.n83 B.n79 4.05904
R1464 B.n692 B.n691 4.05904
R1465 B.n494 B.t3 0.505203
R1466 B.t7 B.n839 0.505203
R1467 VP.n0 VP.t0 233.4
R1468 VP.n0 VP.t1 184.869
R1469 VP VP.n0 0.431812
R1470 VTAIL.n1 VTAIL.t1 46.8209
R1471 VTAIL.n2 VTAIL.t3 46.8207
R1472 VTAIL.n3 VTAIL.t0 46.8207
R1473 VTAIL.n0 VTAIL.t2 46.8207
R1474 VTAIL.n1 VTAIL.n0 31.9531
R1475 VTAIL.n3 VTAIL.n2 29.2807
R1476 VTAIL.n2 VTAIL.n1 1.80653
R1477 VTAIL VTAIL.n0 1.19662
R1478 VTAIL VTAIL.n3 0.610414
R1479 VDD1 VDD1.t0 107.939
R1480 VDD1 VDD1.t1 64.2258
R1481 VN VN.t0 233.401
R1482 VN VN.t1 185.299
R1483 VDD2.n0 VDD2.t0 106.746
R1484 VDD2.n0 VDD2.t1 63.4995
R1485 VDD2 VDD2.n0 0.726793
C0 VDD2 VP 0.340881f
C1 VDD2 VN 3.76937f
C2 VTAIL VDD1 6.27314f
C3 VDD1 VP 3.95851f
C4 VTAIL VP 3.26074f
C5 VDD1 VN 0.148534f
C6 VTAIL VN 3.24641f
C7 VDD1 VDD2 0.695643f
C8 VTAIL VDD2 6.32408f
C9 VP VN 6.37145f
C10 VDD2 B 5.300358f
C11 VDD1 B 8.812981f
C12 VTAIL B 9.266233f
C13 VN B 11.967171f
C14 VP B 6.922541f
C15 VDD2.t0 B 3.70166f
C16 VDD2.t1 B 3.03317f
C17 VDD2.n0 B 3.23157f
C18 VN.t1 B 3.91294f
C19 VN.t0 B 4.48513f
C20 VDD1.t1 B 3.07387f
C21 VDD1.t0 B 3.78785f
C22 VTAIL.t2 B 2.94865f
C23 VTAIL.n0 B 1.87306f
C24 VTAIL.t1 B 2.94866f
C25 VTAIL.n1 B 1.91229f
C26 VTAIL.t3 B 2.94865f
C27 VTAIL.n2 B 1.7404f
C28 VTAIL.t0 B 2.94865f
C29 VTAIL.n3 B 1.66347f
C30 VP.t1 B 4.00954f
C31 VP.t0 B 4.59791f
C32 VP.n0 B 5.01239f
.ends

