* NGSPICE file created from diff_pair_sample_1617.ext - technology: sky130A

.subckt diff_pair_sample_1617 VTAIL VN VP B VDD2 VDD1
X0 B.t17 B.t15 B.t16 B.t5 sky130_fd_pr__nfet_01v8 ad=5.8695 pd=30.88 as=0 ps=0 w=15.05 l=3.63
X1 VDD1.t3 VP.t0 VTAIL.t6 B.t0 sky130_fd_pr__nfet_01v8 ad=2.48325 pd=15.38 as=5.8695 ps=30.88 w=15.05 l=3.63
X2 VTAIL.t4 VP.t1 VDD1.t2 B.t3 sky130_fd_pr__nfet_01v8 ad=5.8695 pd=30.88 as=2.48325 ps=15.38 w=15.05 l=3.63
X3 B.t14 B.t12 B.t13 B.t9 sky130_fd_pr__nfet_01v8 ad=5.8695 pd=30.88 as=0 ps=0 w=15.05 l=3.63
X4 VDD1.t1 VP.t2 VTAIL.t7 B.t2 sky130_fd_pr__nfet_01v8 ad=2.48325 pd=15.38 as=5.8695 ps=30.88 w=15.05 l=3.63
X5 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=5.8695 pd=30.88 as=0 ps=0 w=15.05 l=3.63
X6 VDD2.t3 VN.t0 VTAIL.t1 B.t2 sky130_fd_pr__nfet_01v8 ad=2.48325 pd=15.38 as=5.8695 ps=30.88 w=15.05 l=3.63
X7 B.t7 B.t4 B.t6 B.t5 sky130_fd_pr__nfet_01v8 ad=5.8695 pd=30.88 as=0 ps=0 w=15.05 l=3.63
X8 VDD2.t2 VN.t1 VTAIL.t2 B.t0 sky130_fd_pr__nfet_01v8 ad=2.48325 pd=15.38 as=5.8695 ps=30.88 w=15.05 l=3.63
X9 VTAIL.t3 VN.t2 VDD2.t1 B.t3 sky130_fd_pr__nfet_01v8 ad=5.8695 pd=30.88 as=2.48325 ps=15.38 w=15.05 l=3.63
X10 VTAIL.t0 VN.t3 VDD2.t0 B.t1 sky130_fd_pr__nfet_01v8 ad=5.8695 pd=30.88 as=2.48325 ps=15.38 w=15.05 l=3.63
X11 VTAIL.t5 VP.t3 VDD1.t0 B.t1 sky130_fd_pr__nfet_01v8 ad=5.8695 pd=30.88 as=2.48325 ps=15.38 w=15.05 l=3.63
R0 B.n910 B.n909 585
R1 B.n911 B.n910 585
R2 B.n358 B.n136 585
R3 B.n357 B.n356 585
R4 B.n355 B.n354 585
R5 B.n353 B.n352 585
R6 B.n351 B.n350 585
R7 B.n349 B.n348 585
R8 B.n347 B.n346 585
R9 B.n345 B.n344 585
R10 B.n343 B.n342 585
R11 B.n341 B.n340 585
R12 B.n339 B.n338 585
R13 B.n337 B.n336 585
R14 B.n335 B.n334 585
R15 B.n333 B.n332 585
R16 B.n331 B.n330 585
R17 B.n329 B.n328 585
R18 B.n327 B.n326 585
R19 B.n325 B.n324 585
R20 B.n323 B.n322 585
R21 B.n321 B.n320 585
R22 B.n319 B.n318 585
R23 B.n317 B.n316 585
R24 B.n315 B.n314 585
R25 B.n313 B.n312 585
R26 B.n311 B.n310 585
R27 B.n309 B.n308 585
R28 B.n307 B.n306 585
R29 B.n305 B.n304 585
R30 B.n303 B.n302 585
R31 B.n301 B.n300 585
R32 B.n299 B.n298 585
R33 B.n297 B.n296 585
R34 B.n295 B.n294 585
R35 B.n293 B.n292 585
R36 B.n291 B.n290 585
R37 B.n289 B.n288 585
R38 B.n287 B.n286 585
R39 B.n285 B.n284 585
R40 B.n283 B.n282 585
R41 B.n281 B.n280 585
R42 B.n279 B.n278 585
R43 B.n277 B.n276 585
R44 B.n275 B.n274 585
R45 B.n273 B.n272 585
R46 B.n271 B.n270 585
R47 B.n269 B.n268 585
R48 B.n267 B.n266 585
R49 B.n265 B.n264 585
R50 B.n263 B.n262 585
R51 B.n261 B.n260 585
R52 B.n259 B.n258 585
R53 B.n257 B.n256 585
R54 B.n255 B.n254 585
R55 B.n253 B.n252 585
R56 B.n251 B.n250 585
R57 B.n249 B.n248 585
R58 B.n247 B.n246 585
R59 B.n245 B.n244 585
R60 B.n243 B.n242 585
R61 B.n240 B.n239 585
R62 B.n238 B.n237 585
R63 B.n236 B.n235 585
R64 B.n234 B.n233 585
R65 B.n232 B.n231 585
R66 B.n230 B.n229 585
R67 B.n228 B.n227 585
R68 B.n226 B.n225 585
R69 B.n224 B.n223 585
R70 B.n222 B.n221 585
R71 B.n220 B.n219 585
R72 B.n218 B.n217 585
R73 B.n216 B.n215 585
R74 B.n214 B.n213 585
R75 B.n212 B.n211 585
R76 B.n210 B.n209 585
R77 B.n208 B.n207 585
R78 B.n206 B.n205 585
R79 B.n204 B.n203 585
R80 B.n202 B.n201 585
R81 B.n200 B.n199 585
R82 B.n198 B.n197 585
R83 B.n196 B.n195 585
R84 B.n194 B.n193 585
R85 B.n192 B.n191 585
R86 B.n190 B.n189 585
R87 B.n188 B.n187 585
R88 B.n186 B.n185 585
R89 B.n184 B.n183 585
R90 B.n182 B.n181 585
R91 B.n180 B.n179 585
R92 B.n178 B.n177 585
R93 B.n176 B.n175 585
R94 B.n174 B.n173 585
R95 B.n172 B.n171 585
R96 B.n170 B.n169 585
R97 B.n168 B.n167 585
R98 B.n166 B.n165 585
R99 B.n164 B.n163 585
R100 B.n162 B.n161 585
R101 B.n160 B.n159 585
R102 B.n158 B.n157 585
R103 B.n156 B.n155 585
R104 B.n154 B.n153 585
R105 B.n152 B.n151 585
R106 B.n150 B.n149 585
R107 B.n148 B.n147 585
R108 B.n146 B.n145 585
R109 B.n144 B.n143 585
R110 B.n81 B.n80 585
R111 B.n914 B.n913 585
R112 B.n908 B.n137 585
R113 B.n137 B.n78 585
R114 B.n907 B.n77 585
R115 B.n918 B.n77 585
R116 B.n906 B.n76 585
R117 B.n919 B.n76 585
R118 B.n905 B.n75 585
R119 B.n920 B.n75 585
R120 B.n904 B.n903 585
R121 B.n903 B.n71 585
R122 B.n902 B.n70 585
R123 B.n926 B.n70 585
R124 B.n901 B.n69 585
R125 B.n927 B.n69 585
R126 B.n900 B.n68 585
R127 B.n928 B.n68 585
R128 B.n899 B.n898 585
R129 B.n898 B.n64 585
R130 B.n897 B.n63 585
R131 B.n934 B.n63 585
R132 B.n896 B.n62 585
R133 B.n935 B.n62 585
R134 B.n895 B.n61 585
R135 B.n936 B.n61 585
R136 B.n894 B.n893 585
R137 B.n893 B.n57 585
R138 B.n892 B.n56 585
R139 B.n942 B.n56 585
R140 B.n891 B.n55 585
R141 B.n943 B.n55 585
R142 B.n890 B.n54 585
R143 B.n944 B.n54 585
R144 B.n889 B.n888 585
R145 B.n888 B.n50 585
R146 B.n887 B.n49 585
R147 B.n950 B.n49 585
R148 B.n886 B.n48 585
R149 B.n951 B.n48 585
R150 B.n885 B.n47 585
R151 B.n952 B.n47 585
R152 B.n884 B.n883 585
R153 B.n883 B.n43 585
R154 B.n882 B.n42 585
R155 B.n958 B.n42 585
R156 B.n881 B.n41 585
R157 B.n959 B.n41 585
R158 B.n880 B.n40 585
R159 B.n960 B.n40 585
R160 B.n879 B.n878 585
R161 B.n878 B.n36 585
R162 B.n877 B.n35 585
R163 B.n966 B.n35 585
R164 B.n876 B.n34 585
R165 B.n967 B.n34 585
R166 B.n875 B.n33 585
R167 B.n968 B.n33 585
R168 B.n874 B.n873 585
R169 B.n873 B.n29 585
R170 B.n872 B.n28 585
R171 B.n974 B.n28 585
R172 B.n871 B.n27 585
R173 B.n975 B.n27 585
R174 B.n870 B.n26 585
R175 B.n976 B.n26 585
R176 B.n869 B.n868 585
R177 B.n868 B.n22 585
R178 B.n867 B.n21 585
R179 B.n982 B.n21 585
R180 B.n866 B.n20 585
R181 B.n983 B.n20 585
R182 B.n865 B.n19 585
R183 B.n984 B.n19 585
R184 B.n864 B.n863 585
R185 B.n863 B.n15 585
R186 B.n862 B.n14 585
R187 B.n990 B.n14 585
R188 B.n861 B.n13 585
R189 B.n991 B.n13 585
R190 B.n860 B.n12 585
R191 B.n992 B.n12 585
R192 B.n859 B.n858 585
R193 B.n858 B.n8 585
R194 B.n857 B.n7 585
R195 B.n998 B.n7 585
R196 B.n856 B.n6 585
R197 B.n999 B.n6 585
R198 B.n855 B.n5 585
R199 B.n1000 B.n5 585
R200 B.n854 B.n853 585
R201 B.n853 B.n4 585
R202 B.n852 B.n359 585
R203 B.n852 B.n851 585
R204 B.n842 B.n360 585
R205 B.n361 B.n360 585
R206 B.n844 B.n843 585
R207 B.n845 B.n844 585
R208 B.n841 B.n366 585
R209 B.n366 B.n365 585
R210 B.n840 B.n839 585
R211 B.n839 B.n838 585
R212 B.n368 B.n367 585
R213 B.n369 B.n368 585
R214 B.n831 B.n830 585
R215 B.n832 B.n831 585
R216 B.n829 B.n374 585
R217 B.n374 B.n373 585
R218 B.n828 B.n827 585
R219 B.n827 B.n826 585
R220 B.n376 B.n375 585
R221 B.n377 B.n376 585
R222 B.n819 B.n818 585
R223 B.n820 B.n819 585
R224 B.n817 B.n382 585
R225 B.n382 B.n381 585
R226 B.n816 B.n815 585
R227 B.n815 B.n814 585
R228 B.n384 B.n383 585
R229 B.n385 B.n384 585
R230 B.n807 B.n806 585
R231 B.n808 B.n807 585
R232 B.n805 B.n390 585
R233 B.n390 B.n389 585
R234 B.n804 B.n803 585
R235 B.n803 B.n802 585
R236 B.n392 B.n391 585
R237 B.n393 B.n392 585
R238 B.n795 B.n794 585
R239 B.n796 B.n795 585
R240 B.n793 B.n398 585
R241 B.n398 B.n397 585
R242 B.n792 B.n791 585
R243 B.n791 B.n790 585
R244 B.n400 B.n399 585
R245 B.n401 B.n400 585
R246 B.n783 B.n782 585
R247 B.n784 B.n783 585
R248 B.n781 B.n406 585
R249 B.n406 B.n405 585
R250 B.n780 B.n779 585
R251 B.n779 B.n778 585
R252 B.n408 B.n407 585
R253 B.n409 B.n408 585
R254 B.n771 B.n770 585
R255 B.n772 B.n771 585
R256 B.n769 B.n414 585
R257 B.n414 B.n413 585
R258 B.n768 B.n767 585
R259 B.n767 B.n766 585
R260 B.n416 B.n415 585
R261 B.n417 B.n416 585
R262 B.n759 B.n758 585
R263 B.n760 B.n759 585
R264 B.n757 B.n422 585
R265 B.n422 B.n421 585
R266 B.n756 B.n755 585
R267 B.n755 B.n754 585
R268 B.n424 B.n423 585
R269 B.n425 B.n424 585
R270 B.n747 B.n746 585
R271 B.n748 B.n747 585
R272 B.n745 B.n430 585
R273 B.n430 B.n429 585
R274 B.n744 B.n743 585
R275 B.n743 B.n742 585
R276 B.n432 B.n431 585
R277 B.n433 B.n432 585
R278 B.n735 B.n734 585
R279 B.n736 B.n735 585
R280 B.n733 B.n438 585
R281 B.n438 B.n437 585
R282 B.n732 B.n731 585
R283 B.n731 B.n730 585
R284 B.n440 B.n439 585
R285 B.n441 B.n440 585
R286 B.n726 B.n725 585
R287 B.n444 B.n443 585
R288 B.n722 B.n721 585
R289 B.n723 B.n722 585
R290 B.n720 B.n499 585
R291 B.n719 B.n718 585
R292 B.n717 B.n716 585
R293 B.n715 B.n714 585
R294 B.n713 B.n712 585
R295 B.n711 B.n710 585
R296 B.n709 B.n708 585
R297 B.n707 B.n706 585
R298 B.n705 B.n704 585
R299 B.n703 B.n702 585
R300 B.n701 B.n700 585
R301 B.n699 B.n698 585
R302 B.n697 B.n696 585
R303 B.n695 B.n694 585
R304 B.n693 B.n692 585
R305 B.n691 B.n690 585
R306 B.n689 B.n688 585
R307 B.n687 B.n686 585
R308 B.n685 B.n684 585
R309 B.n683 B.n682 585
R310 B.n681 B.n680 585
R311 B.n679 B.n678 585
R312 B.n677 B.n676 585
R313 B.n675 B.n674 585
R314 B.n673 B.n672 585
R315 B.n671 B.n670 585
R316 B.n669 B.n668 585
R317 B.n667 B.n666 585
R318 B.n665 B.n664 585
R319 B.n663 B.n662 585
R320 B.n661 B.n660 585
R321 B.n659 B.n658 585
R322 B.n657 B.n656 585
R323 B.n655 B.n654 585
R324 B.n653 B.n652 585
R325 B.n651 B.n650 585
R326 B.n649 B.n648 585
R327 B.n647 B.n646 585
R328 B.n645 B.n644 585
R329 B.n643 B.n642 585
R330 B.n641 B.n640 585
R331 B.n639 B.n638 585
R332 B.n637 B.n636 585
R333 B.n635 B.n634 585
R334 B.n633 B.n632 585
R335 B.n631 B.n630 585
R336 B.n629 B.n628 585
R337 B.n627 B.n626 585
R338 B.n625 B.n624 585
R339 B.n623 B.n622 585
R340 B.n621 B.n620 585
R341 B.n619 B.n618 585
R342 B.n617 B.n616 585
R343 B.n615 B.n614 585
R344 B.n613 B.n612 585
R345 B.n611 B.n610 585
R346 B.n609 B.n608 585
R347 B.n606 B.n605 585
R348 B.n604 B.n603 585
R349 B.n602 B.n601 585
R350 B.n600 B.n599 585
R351 B.n598 B.n597 585
R352 B.n596 B.n595 585
R353 B.n594 B.n593 585
R354 B.n592 B.n591 585
R355 B.n590 B.n589 585
R356 B.n588 B.n587 585
R357 B.n586 B.n585 585
R358 B.n584 B.n583 585
R359 B.n582 B.n581 585
R360 B.n580 B.n579 585
R361 B.n578 B.n577 585
R362 B.n576 B.n575 585
R363 B.n574 B.n573 585
R364 B.n572 B.n571 585
R365 B.n570 B.n569 585
R366 B.n568 B.n567 585
R367 B.n566 B.n565 585
R368 B.n564 B.n563 585
R369 B.n562 B.n561 585
R370 B.n560 B.n559 585
R371 B.n558 B.n557 585
R372 B.n556 B.n555 585
R373 B.n554 B.n553 585
R374 B.n552 B.n551 585
R375 B.n550 B.n549 585
R376 B.n548 B.n547 585
R377 B.n546 B.n545 585
R378 B.n544 B.n543 585
R379 B.n542 B.n541 585
R380 B.n540 B.n539 585
R381 B.n538 B.n537 585
R382 B.n536 B.n535 585
R383 B.n534 B.n533 585
R384 B.n532 B.n531 585
R385 B.n530 B.n529 585
R386 B.n528 B.n527 585
R387 B.n526 B.n525 585
R388 B.n524 B.n523 585
R389 B.n522 B.n521 585
R390 B.n520 B.n519 585
R391 B.n518 B.n517 585
R392 B.n516 B.n515 585
R393 B.n514 B.n513 585
R394 B.n512 B.n511 585
R395 B.n510 B.n509 585
R396 B.n508 B.n507 585
R397 B.n506 B.n505 585
R398 B.n727 B.n442 585
R399 B.n442 B.n441 585
R400 B.n729 B.n728 585
R401 B.n730 B.n729 585
R402 B.n436 B.n435 585
R403 B.n437 B.n436 585
R404 B.n738 B.n737 585
R405 B.n737 B.n736 585
R406 B.n739 B.n434 585
R407 B.n434 B.n433 585
R408 B.n741 B.n740 585
R409 B.n742 B.n741 585
R410 B.n428 B.n427 585
R411 B.n429 B.n428 585
R412 B.n750 B.n749 585
R413 B.n749 B.n748 585
R414 B.n751 B.n426 585
R415 B.n426 B.n425 585
R416 B.n753 B.n752 585
R417 B.n754 B.n753 585
R418 B.n420 B.n419 585
R419 B.n421 B.n420 585
R420 B.n762 B.n761 585
R421 B.n761 B.n760 585
R422 B.n763 B.n418 585
R423 B.n418 B.n417 585
R424 B.n765 B.n764 585
R425 B.n766 B.n765 585
R426 B.n412 B.n411 585
R427 B.n413 B.n412 585
R428 B.n774 B.n773 585
R429 B.n773 B.n772 585
R430 B.n775 B.n410 585
R431 B.n410 B.n409 585
R432 B.n777 B.n776 585
R433 B.n778 B.n777 585
R434 B.n404 B.n403 585
R435 B.n405 B.n404 585
R436 B.n786 B.n785 585
R437 B.n785 B.n784 585
R438 B.n787 B.n402 585
R439 B.n402 B.n401 585
R440 B.n789 B.n788 585
R441 B.n790 B.n789 585
R442 B.n396 B.n395 585
R443 B.n397 B.n396 585
R444 B.n798 B.n797 585
R445 B.n797 B.n796 585
R446 B.n799 B.n394 585
R447 B.n394 B.n393 585
R448 B.n801 B.n800 585
R449 B.n802 B.n801 585
R450 B.n388 B.n387 585
R451 B.n389 B.n388 585
R452 B.n810 B.n809 585
R453 B.n809 B.n808 585
R454 B.n811 B.n386 585
R455 B.n386 B.n385 585
R456 B.n813 B.n812 585
R457 B.n814 B.n813 585
R458 B.n380 B.n379 585
R459 B.n381 B.n380 585
R460 B.n822 B.n821 585
R461 B.n821 B.n820 585
R462 B.n823 B.n378 585
R463 B.n378 B.n377 585
R464 B.n825 B.n824 585
R465 B.n826 B.n825 585
R466 B.n372 B.n371 585
R467 B.n373 B.n372 585
R468 B.n834 B.n833 585
R469 B.n833 B.n832 585
R470 B.n835 B.n370 585
R471 B.n370 B.n369 585
R472 B.n837 B.n836 585
R473 B.n838 B.n837 585
R474 B.n364 B.n363 585
R475 B.n365 B.n364 585
R476 B.n847 B.n846 585
R477 B.n846 B.n845 585
R478 B.n848 B.n362 585
R479 B.n362 B.n361 585
R480 B.n850 B.n849 585
R481 B.n851 B.n850 585
R482 B.n2 B.n0 585
R483 B.n4 B.n2 585
R484 B.n3 B.n1 585
R485 B.n999 B.n3 585
R486 B.n997 B.n996 585
R487 B.n998 B.n997 585
R488 B.n995 B.n9 585
R489 B.n9 B.n8 585
R490 B.n994 B.n993 585
R491 B.n993 B.n992 585
R492 B.n11 B.n10 585
R493 B.n991 B.n11 585
R494 B.n989 B.n988 585
R495 B.n990 B.n989 585
R496 B.n987 B.n16 585
R497 B.n16 B.n15 585
R498 B.n986 B.n985 585
R499 B.n985 B.n984 585
R500 B.n18 B.n17 585
R501 B.n983 B.n18 585
R502 B.n981 B.n980 585
R503 B.n982 B.n981 585
R504 B.n979 B.n23 585
R505 B.n23 B.n22 585
R506 B.n978 B.n977 585
R507 B.n977 B.n976 585
R508 B.n25 B.n24 585
R509 B.n975 B.n25 585
R510 B.n973 B.n972 585
R511 B.n974 B.n973 585
R512 B.n971 B.n30 585
R513 B.n30 B.n29 585
R514 B.n970 B.n969 585
R515 B.n969 B.n968 585
R516 B.n32 B.n31 585
R517 B.n967 B.n32 585
R518 B.n965 B.n964 585
R519 B.n966 B.n965 585
R520 B.n963 B.n37 585
R521 B.n37 B.n36 585
R522 B.n962 B.n961 585
R523 B.n961 B.n960 585
R524 B.n39 B.n38 585
R525 B.n959 B.n39 585
R526 B.n957 B.n956 585
R527 B.n958 B.n957 585
R528 B.n955 B.n44 585
R529 B.n44 B.n43 585
R530 B.n954 B.n953 585
R531 B.n953 B.n952 585
R532 B.n46 B.n45 585
R533 B.n951 B.n46 585
R534 B.n949 B.n948 585
R535 B.n950 B.n949 585
R536 B.n947 B.n51 585
R537 B.n51 B.n50 585
R538 B.n946 B.n945 585
R539 B.n945 B.n944 585
R540 B.n53 B.n52 585
R541 B.n943 B.n53 585
R542 B.n941 B.n940 585
R543 B.n942 B.n941 585
R544 B.n939 B.n58 585
R545 B.n58 B.n57 585
R546 B.n938 B.n937 585
R547 B.n937 B.n936 585
R548 B.n60 B.n59 585
R549 B.n935 B.n60 585
R550 B.n933 B.n932 585
R551 B.n934 B.n933 585
R552 B.n931 B.n65 585
R553 B.n65 B.n64 585
R554 B.n930 B.n929 585
R555 B.n929 B.n928 585
R556 B.n67 B.n66 585
R557 B.n927 B.n67 585
R558 B.n925 B.n924 585
R559 B.n926 B.n925 585
R560 B.n923 B.n72 585
R561 B.n72 B.n71 585
R562 B.n922 B.n921 585
R563 B.n921 B.n920 585
R564 B.n74 B.n73 585
R565 B.n919 B.n74 585
R566 B.n917 B.n916 585
R567 B.n918 B.n917 585
R568 B.n915 B.n79 585
R569 B.n79 B.n78 585
R570 B.n1002 B.n1001 585
R571 B.n1001 B.n1000 585
R572 B.n725 B.n442 487.695
R573 B.n913 B.n79 487.695
R574 B.n505 B.n440 487.695
R575 B.n910 B.n137 487.695
R576 B.n503 B.t15 309.125
R577 B.n500 B.t4 309.125
R578 B.n141 B.t8 309.125
R579 B.n138 B.t12 309.125
R580 B.n911 B.n135 256.663
R581 B.n911 B.n134 256.663
R582 B.n911 B.n133 256.663
R583 B.n911 B.n132 256.663
R584 B.n911 B.n131 256.663
R585 B.n911 B.n130 256.663
R586 B.n911 B.n129 256.663
R587 B.n911 B.n128 256.663
R588 B.n911 B.n127 256.663
R589 B.n911 B.n126 256.663
R590 B.n911 B.n125 256.663
R591 B.n911 B.n124 256.663
R592 B.n911 B.n123 256.663
R593 B.n911 B.n122 256.663
R594 B.n911 B.n121 256.663
R595 B.n911 B.n120 256.663
R596 B.n911 B.n119 256.663
R597 B.n911 B.n118 256.663
R598 B.n911 B.n117 256.663
R599 B.n911 B.n116 256.663
R600 B.n911 B.n115 256.663
R601 B.n911 B.n114 256.663
R602 B.n911 B.n113 256.663
R603 B.n911 B.n112 256.663
R604 B.n911 B.n111 256.663
R605 B.n911 B.n110 256.663
R606 B.n911 B.n109 256.663
R607 B.n911 B.n108 256.663
R608 B.n911 B.n107 256.663
R609 B.n911 B.n106 256.663
R610 B.n911 B.n105 256.663
R611 B.n911 B.n104 256.663
R612 B.n911 B.n103 256.663
R613 B.n911 B.n102 256.663
R614 B.n911 B.n101 256.663
R615 B.n911 B.n100 256.663
R616 B.n911 B.n99 256.663
R617 B.n911 B.n98 256.663
R618 B.n911 B.n97 256.663
R619 B.n911 B.n96 256.663
R620 B.n911 B.n95 256.663
R621 B.n911 B.n94 256.663
R622 B.n911 B.n93 256.663
R623 B.n911 B.n92 256.663
R624 B.n911 B.n91 256.663
R625 B.n911 B.n90 256.663
R626 B.n911 B.n89 256.663
R627 B.n911 B.n88 256.663
R628 B.n911 B.n87 256.663
R629 B.n911 B.n86 256.663
R630 B.n911 B.n85 256.663
R631 B.n911 B.n84 256.663
R632 B.n911 B.n83 256.663
R633 B.n911 B.n82 256.663
R634 B.n912 B.n911 256.663
R635 B.n724 B.n723 256.663
R636 B.n723 B.n445 256.663
R637 B.n723 B.n446 256.663
R638 B.n723 B.n447 256.663
R639 B.n723 B.n448 256.663
R640 B.n723 B.n449 256.663
R641 B.n723 B.n450 256.663
R642 B.n723 B.n451 256.663
R643 B.n723 B.n452 256.663
R644 B.n723 B.n453 256.663
R645 B.n723 B.n454 256.663
R646 B.n723 B.n455 256.663
R647 B.n723 B.n456 256.663
R648 B.n723 B.n457 256.663
R649 B.n723 B.n458 256.663
R650 B.n723 B.n459 256.663
R651 B.n723 B.n460 256.663
R652 B.n723 B.n461 256.663
R653 B.n723 B.n462 256.663
R654 B.n723 B.n463 256.663
R655 B.n723 B.n464 256.663
R656 B.n723 B.n465 256.663
R657 B.n723 B.n466 256.663
R658 B.n723 B.n467 256.663
R659 B.n723 B.n468 256.663
R660 B.n723 B.n469 256.663
R661 B.n723 B.n470 256.663
R662 B.n723 B.n471 256.663
R663 B.n723 B.n472 256.663
R664 B.n723 B.n473 256.663
R665 B.n723 B.n474 256.663
R666 B.n723 B.n475 256.663
R667 B.n723 B.n476 256.663
R668 B.n723 B.n477 256.663
R669 B.n723 B.n478 256.663
R670 B.n723 B.n479 256.663
R671 B.n723 B.n480 256.663
R672 B.n723 B.n481 256.663
R673 B.n723 B.n482 256.663
R674 B.n723 B.n483 256.663
R675 B.n723 B.n484 256.663
R676 B.n723 B.n485 256.663
R677 B.n723 B.n486 256.663
R678 B.n723 B.n487 256.663
R679 B.n723 B.n488 256.663
R680 B.n723 B.n489 256.663
R681 B.n723 B.n490 256.663
R682 B.n723 B.n491 256.663
R683 B.n723 B.n492 256.663
R684 B.n723 B.n493 256.663
R685 B.n723 B.n494 256.663
R686 B.n723 B.n495 256.663
R687 B.n723 B.n496 256.663
R688 B.n723 B.n497 256.663
R689 B.n723 B.n498 256.663
R690 B.n729 B.n442 163.367
R691 B.n729 B.n436 163.367
R692 B.n737 B.n436 163.367
R693 B.n737 B.n434 163.367
R694 B.n741 B.n434 163.367
R695 B.n741 B.n428 163.367
R696 B.n749 B.n428 163.367
R697 B.n749 B.n426 163.367
R698 B.n753 B.n426 163.367
R699 B.n753 B.n420 163.367
R700 B.n761 B.n420 163.367
R701 B.n761 B.n418 163.367
R702 B.n765 B.n418 163.367
R703 B.n765 B.n412 163.367
R704 B.n773 B.n412 163.367
R705 B.n773 B.n410 163.367
R706 B.n777 B.n410 163.367
R707 B.n777 B.n404 163.367
R708 B.n785 B.n404 163.367
R709 B.n785 B.n402 163.367
R710 B.n789 B.n402 163.367
R711 B.n789 B.n396 163.367
R712 B.n797 B.n396 163.367
R713 B.n797 B.n394 163.367
R714 B.n801 B.n394 163.367
R715 B.n801 B.n388 163.367
R716 B.n809 B.n388 163.367
R717 B.n809 B.n386 163.367
R718 B.n813 B.n386 163.367
R719 B.n813 B.n380 163.367
R720 B.n821 B.n380 163.367
R721 B.n821 B.n378 163.367
R722 B.n825 B.n378 163.367
R723 B.n825 B.n372 163.367
R724 B.n833 B.n372 163.367
R725 B.n833 B.n370 163.367
R726 B.n837 B.n370 163.367
R727 B.n837 B.n364 163.367
R728 B.n846 B.n364 163.367
R729 B.n846 B.n362 163.367
R730 B.n850 B.n362 163.367
R731 B.n850 B.n2 163.367
R732 B.n1001 B.n2 163.367
R733 B.n1001 B.n3 163.367
R734 B.n997 B.n3 163.367
R735 B.n997 B.n9 163.367
R736 B.n993 B.n9 163.367
R737 B.n993 B.n11 163.367
R738 B.n989 B.n11 163.367
R739 B.n989 B.n16 163.367
R740 B.n985 B.n16 163.367
R741 B.n985 B.n18 163.367
R742 B.n981 B.n18 163.367
R743 B.n981 B.n23 163.367
R744 B.n977 B.n23 163.367
R745 B.n977 B.n25 163.367
R746 B.n973 B.n25 163.367
R747 B.n973 B.n30 163.367
R748 B.n969 B.n30 163.367
R749 B.n969 B.n32 163.367
R750 B.n965 B.n32 163.367
R751 B.n965 B.n37 163.367
R752 B.n961 B.n37 163.367
R753 B.n961 B.n39 163.367
R754 B.n957 B.n39 163.367
R755 B.n957 B.n44 163.367
R756 B.n953 B.n44 163.367
R757 B.n953 B.n46 163.367
R758 B.n949 B.n46 163.367
R759 B.n949 B.n51 163.367
R760 B.n945 B.n51 163.367
R761 B.n945 B.n53 163.367
R762 B.n941 B.n53 163.367
R763 B.n941 B.n58 163.367
R764 B.n937 B.n58 163.367
R765 B.n937 B.n60 163.367
R766 B.n933 B.n60 163.367
R767 B.n933 B.n65 163.367
R768 B.n929 B.n65 163.367
R769 B.n929 B.n67 163.367
R770 B.n925 B.n67 163.367
R771 B.n925 B.n72 163.367
R772 B.n921 B.n72 163.367
R773 B.n921 B.n74 163.367
R774 B.n917 B.n74 163.367
R775 B.n917 B.n79 163.367
R776 B.n722 B.n444 163.367
R777 B.n722 B.n499 163.367
R778 B.n718 B.n717 163.367
R779 B.n714 B.n713 163.367
R780 B.n710 B.n709 163.367
R781 B.n706 B.n705 163.367
R782 B.n702 B.n701 163.367
R783 B.n698 B.n697 163.367
R784 B.n694 B.n693 163.367
R785 B.n690 B.n689 163.367
R786 B.n686 B.n685 163.367
R787 B.n682 B.n681 163.367
R788 B.n678 B.n677 163.367
R789 B.n674 B.n673 163.367
R790 B.n670 B.n669 163.367
R791 B.n666 B.n665 163.367
R792 B.n662 B.n661 163.367
R793 B.n658 B.n657 163.367
R794 B.n654 B.n653 163.367
R795 B.n650 B.n649 163.367
R796 B.n646 B.n645 163.367
R797 B.n642 B.n641 163.367
R798 B.n638 B.n637 163.367
R799 B.n634 B.n633 163.367
R800 B.n630 B.n629 163.367
R801 B.n626 B.n625 163.367
R802 B.n622 B.n621 163.367
R803 B.n618 B.n617 163.367
R804 B.n614 B.n613 163.367
R805 B.n610 B.n609 163.367
R806 B.n605 B.n604 163.367
R807 B.n601 B.n600 163.367
R808 B.n597 B.n596 163.367
R809 B.n593 B.n592 163.367
R810 B.n589 B.n588 163.367
R811 B.n585 B.n584 163.367
R812 B.n581 B.n580 163.367
R813 B.n577 B.n576 163.367
R814 B.n573 B.n572 163.367
R815 B.n569 B.n568 163.367
R816 B.n565 B.n564 163.367
R817 B.n561 B.n560 163.367
R818 B.n557 B.n556 163.367
R819 B.n553 B.n552 163.367
R820 B.n549 B.n548 163.367
R821 B.n545 B.n544 163.367
R822 B.n541 B.n540 163.367
R823 B.n537 B.n536 163.367
R824 B.n533 B.n532 163.367
R825 B.n529 B.n528 163.367
R826 B.n525 B.n524 163.367
R827 B.n521 B.n520 163.367
R828 B.n517 B.n516 163.367
R829 B.n513 B.n512 163.367
R830 B.n509 B.n508 163.367
R831 B.n731 B.n440 163.367
R832 B.n731 B.n438 163.367
R833 B.n735 B.n438 163.367
R834 B.n735 B.n432 163.367
R835 B.n743 B.n432 163.367
R836 B.n743 B.n430 163.367
R837 B.n747 B.n430 163.367
R838 B.n747 B.n424 163.367
R839 B.n755 B.n424 163.367
R840 B.n755 B.n422 163.367
R841 B.n759 B.n422 163.367
R842 B.n759 B.n416 163.367
R843 B.n767 B.n416 163.367
R844 B.n767 B.n414 163.367
R845 B.n771 B.n414 163.367
R846 B.n771 B.n408 163.367
R847 B.n779 B.n408 163.367
R848 B.n779 B.n406 163.367
R849 B.n783 B.n406 163.367
R850 B.n783 B.n400 163.367
R851 B.n791 B.n400 163.367
R852 B.n791 B.n398 163.367
R853 B.n795 B.n398 163.367
R854 B.n795 B.n392 163.367
R855 B.n803 B.n392 163.367
R856 B.n803 B.n390 163.367
R857 B.n807 B.n390 163.367
R858 B.n807 B.n384 163.367
R859 B.n815 B.n384 163.367
R860 B.n815 B.n382 163.367
R861 B.n819 B.n382 163.367
R862 B.n819 B.n376 163.367
R863 B.n827 B.n376 163.367
R864 B.n827 B.n374 163.367
R865 B.n831 B.n374 163.367
R866 B.n831 B.n368 163.367
R867 B.n839 B.n368 163.367
R868 B.n839 B.n366 163.367
R869 B.n844 B.n366 163.367
R870 B.n844 B.n360 163.367
R871 B.n852 B.n360 163.367
R872 B.n853 B.n852 163.367
R873 B.n853 B.n5 163.367
R874 B.n6 B.n5 163.367
R875 B.n7 B.n6 163.367
R876 B.n858 B.n7 163.367
R877 B.n858 B.n12 163.367
R878 B.n13 B.n12 163.367
R879 B.n14 B.n13 163.367
R880 B.n863 B.n14 163.367
R881 B.n863 B.n19 163.367
R882 B.n20 B.n19 163.367
R883 B.n21 B.n20 163.367
R884 B.n868 B.n21 163.367
R885 B.n868 B.n26 163.367
R886 B.n27 B.n26 163.367
R887 B.n28 B.n27 163.367
R888 B.n873 B.n28 163.367
R889 B.n873 B.n33 163.367
R890 B.n34 B.n33 163.367
R891 B.n35 B.n34 163.367
R892 B.n878 B.n35 163.367
R893 B.n878 B.n40 163.367
R894 B.n41 B.n40 163.367
R895 B.n42 B.n41 163.367
R896 B.n883 B.n42 163.367
R897 B.n883 B.n47 163.367
R898 B.n48 B.n47 163.367
R899 B.n49 B.n48 163.367
R900 B.n888 B.n49 163.367
R901 B.n888 B.n54 163.367
R902 B.n55 B.n54 163.367
R903 B.n56 B.n55 163.367
R904 B.n893 B.n56 163.367
R905 B.n893 B.n61 163.367
R906 B.n62 B.n61 163.367
R907 B.n63 B.n62 163.367
R908 B.n898 B.n63 163.367
R909 B.n898 B.n68 163.367
R910 B.n69 B.n68 163.367
R911 B.n70 B.n69 163.367
R912 B.n903 B.n70 163.367
R913 B.n903 B.n75 163.367
R914 B.n76 B.n75 163.367
R915 B.n77 B.n76 163.367
R916 B.n137 B.n77 163.367
R917 B.n143 B.n81 163.367
R918 B.n147 B.n146 163.367
R919 B.n151 B.n150 163.367
R920 B.n155 B.n154 163.367
R921 B.n159 B.n158 163.367
R922 B.n163 B.n162 163.367
R923 B.n167 B.n166 163.367
R924 B.n171 B.n170 163.367
R925 B.n175 B.n174 163.367
R926 B.n179 B.n178 163.367
R927 B.n183 B.n182 163.367
R928 B.n187 B.n186 163.367
R929 B.n191 B.n190 163.367
R930 B.n195 B.n194 163.367
R931 B.n199 B.n198 163.367
R932 B.n203 B.n202 163.367
R933 B.n207 B.n206 163.367
R934 B.n211 B.n210 163.367
R935 B.n215 B.n214 163.367
R936 B.n219 B.n218 163.367
R937 B.n223 B.n222 163.367
R938 B.n227 B.n226 163.367
R939 B.n231 B.n230 163.367
R940 B.n235 B.n234 163.367
R941 B.n239 B.n238 163.367
R942 B.n244 B.n243 163.367
R943 B.n248 B.n247 163.367
R944 B.n252 B.n251 163.367
R945 B.n256 B.n255 163.367
R946 B.n260 B.n259 163.367
R947 B.n264 B.n263 163.367
R948 B.n268 B.n267 163.367
R949 B.n272 B.n271 163.367
R950 B.n276 B.n275 163.367
R951 B.n280 B.n279 163.367
R952 B.n284 B.n283 163.367
R953 B.n288 B.n287 163.367
R954 B.n292 B.n291 163.367
R955 B.n296 B.n295 163.367
R956 B.n300 B.n299 163.367
R957 B.n304 B.n303 163.367
R958 B.n308 B.n307 163.367
R959 B.n312 B.n311 163.367
R960 B.n316 B.n315 163.367
R961 B.n320 B.n319 163.367
R962 B.n324 B.n323 163.367
R963 B.n328 B.n327 163.367
R964 B.n332 B.n331 163.367
R965 B.n336 B.n335 163.367
R966 B.n340 B.n339 163.367
R967 B.n344 B.n343 163.367
R968 B.n348 B.n347 163.367
R969 B.n352 B.n351 163.367
R970 B.n356 B.n355 163.367
R971 B.n910 B.n136 163.367
R972 B.n503 B.t17 146.006
R973 B.n138 B.t13 146.006
R974 B.n500 B.t7 145.986
R975 B.n141 B.t10 145.986
R976 B.n504 B.n503 76.8005
R977 B.n501 B.n500 76.8005
R978 B.n142 B.n141 76.8005
R979 B.n139 B.n138 76.8005
R980 B.n725 B.n724 71.676
R981 B.n499 B.n445 71.676
R982 B.n717 B.n446 71.676
R983 B.n713 B.n447 71.676
R984 B.n709 B.n448 71.676
R985 B.n705 B.n449 71.676
R986 B.n701 B.n450 71.676
R987 B.n697 B.n451 71.676
R988 B.n693 B.n452 71.676
R989 B.n689 B.n453 71.676
R990 B.n685 B.n454 71.676
R991 B.n681 B.n455 71.676
R992 B.n677 B.n456 71.676
R993 B.n673 B.n457 71.676
R994 B.n669 B.n458 71.676
R995 B.n665 B.n459 71.676
R996 B.n661 B.n460 71.676
R997 B.n657 B.n461 71.676
R998 B.n653 B.n462 71.676
R999 B.n649 B.n463 71.676
R1000 B.n645 B.n464 71.676
R1001 B.n641 B.n465 71.676
R1002 B.n637 B.n466 71.676
R1003 B.n633 B.n467 71.676
R1004 B.n629 B.n468 71.676
R1005 B.n625 B.n469 71.676
R1006 B.n621 B.n470 71.676
R1007 B.n617 B.n471 71.676
R1008 B.n613 B.n472 71.676
R1009 B.n609 B.n473 71.676
R1010 B.n604 B.n474 71.676
R1011 B.n600 B.n475 71.676
R1012 B.n596 B.n476 71.676
R1013 B.n592 B.n477 71.676
R1014 B.n588 B.n478 71.676
R1015 B.n584 B.n479 71.676
R1016 B.n580 B.n480 71.676
R1017 B.n576 B.n481 71.676
R1018 B.n572 B.n482 71.676
R1019 B.n568 B.n483 71.676
R1020 B.n564 B.n484 71.676
R1021 B.n560 B.n485 71.676
R1022 B.n556 B.n486 71.676
R1023 B.n552 B.n487 71.676
R1024 B.n548 B.n488 71.676
R1025 B.n544 B.n489 71.676
R1026 B.n540 B.n490 71.676
R1027 B.n536 B.n491 71.676
R1028 B.n532 B.n492 71.676
R1029 B.n528 B.n493 71.676
R1030 B.n524 B.n494 71.676
R1031 B.n520 B.n495 71.676
R1032 B.n516 B.n496 71.676
R1033 B.n512 B.n497 71.676
R1034 B.n508 B.n498 71.676
R1035 B.n913 B.n912 71.676
R1036 B.n143 B.n82 71.676
R1037 B.n147 B.n83 71.676
R1038 B.n151 B.n84 71.676
R1039 B.n155 B.n85 71.676
R1040 B.n159 B.n86 71.676
R1041 B.n163 B.n87 71.676
R1042 B.n167 B.n88 71.676
R1043 B.n171 B.n89 71.676
R1044 B.n175 B.n90 71.676
R1045 B.n179 B.n91 71.676
R1046 B.n183 B.n92 71.676
R1047 B.n187 B.n93 71.676
R1048 B.n191 B.n94 71.676
R1049 B.n195 B.n95 71.676
R1050 B.n199 B.n96 71.676
R1051 B.n203 B.n97 71.676
R1052 B.n207 B.n98 71.676
R1053 B.n211 B.n99 71.676
R1054 B.n215 B.n100 71.676
R1055 B.n219 B.n101 71.676
R1056 B.n223 B.n102 71.676
R1057 B.n227 B.n103 71.676
R1058 B.n231 B.n104 71.676
R1059 B.n235 B.n105 71.676
R1060 B.n239 B.n106 71.676
R1061 B.n244 B.n107 71.676
R1062 B.n248 B.n108 71.676
R1063 B.n252 B.n109 71.676
R1064 B.n256 B.n110 71.676
R1065 B.n260 B.n111 71.676
R1066 B.n264 B.n112 71.676
R1067 B.n268 B.n113 71.676
R1068 B.n272 B.n114 71.676
R1069 B.n276 B.n115 71.676
R1070 B.n280 B.n116 71.676
R1071 B.n284 B.n117 71.676
R1072 B.n288 B.n118 71.676
R1073 B.n292 B.n119 71.676
R1074 B.n296 B.n120 71.676
R1075 B.n300 B.n121 71.676
R1076 B.n304 B.n122 71.676
R1077 B.n308 B.n123 71.676
R1078 B.n312 B.n124 71.676
R1079 B.n316 B.n125 71.676
R1080 B.n320 B.n126 71.676
R1081 B.n324 B.n127 71.676
R1082 B.n328 B.n128 71.676
R1083 B.n332 B.n129 71.676
R1084 B.n336 B.n130 71.676
R1085 B.n340 B.n131 71.676
R1086 B.n344 B.n132 71.676
R1087 B.n348 B.n133 71.676
R1088 B.n352 B.n134 71.676
R1089 B.n356 B.n135 71.676
R1090 B.n136 B.n135 71.676
R1091 B.n355 B.n134 71.676
R1092 B.n351 B.n133 71.676
R1093 B.n347 B.n132 71.676
R1094 B.n343 B.n131 71.676
R1095 B.n339 B.n130 71.676
R1096 B.n335 B.n129 71.676
R1097 B.n331 B.n128 71.676
R1098 B.n327 B.n127 71.676
R1099 B.n323 B.n126 71.676
R1100 B.n319 B.n125 71.676
R1101 B.n315 B.n124 71.676
R1102 B.n311 B.n123 71.676
R1103 B.n307 B.n122 71.676
R1104 B.n303 B.n121 71.676
R1105 B.n299 B.n120 71.676
R1106 B.n295 B.n119 71.676
R1107 B.n291 B.n118 71.676
R1108 B.n287 B.n117 71.676
R1109 B.n283 B.n116 71.676
R1110 B.n279 B.n115 71.676
R1111 B.n275 B.n114 71.676
R1112 B.n271 B.n113 71.676
R1113 B.n267 B.n112 71.676
R1114 B.n263 B.n111 71.676
R1115 B.n259 B.n110 71.676
R1116 B.n255 B.n109 71.676
R1117 B.n251 B.n108 71.676
R1118 B.n247 B.n107 71.676
R1119 B.n243 B.n106 71.676
R1120 B.n238 B.n105 71.676
R1121 B.n234 B.n104 71.676
R1122 B.n230 B.n103 71.676
R1123 B.n226 B.n102 71.676
R1124 B.n222 B.n101 71.676
R1125 B.n218 B.n100 71.676
R1126 B.n214 B.n99 71.676
R1127 B.n210 B.n98 71.676
R1128 B.n206 B.n97 71.676
R1129 B.n202 B.n96 71.676
R1130 B.n198 B.n95 71.676
R1131 B.n194 B.n94 71.676
R1132 B.n190 B.n93 71.676
R1133 B.n186 B.n92 71.676
R1134 B.n182 B.n91 71.676
R1135 B.n178 B.n90 71.676
R1136 B.n174 B.n89 71.676
R1137 B.n170 B.n88 71.676
R1138 B.n166 B.n87 71.676
R1139 B.n162 B.n86 71.676
R1140 B.n158 B.n85 71.676
R1141 B.n154 B.n84 71.676
R1142 B.n150 B.n83 71.676
R1143 B.n146 B.n82 71.676
R1144 B.n912 B.n81 71.676
R1145 B.n724 B.n444 71.676
R1146 B.n718 B.n445 71.676
R1147 B.n714 B.n446 71.676
R1148 B.n710 B.n447 71.676
R1149 B.n706 B.n448 71.676
R1150 B.n702 B.n449 71.676
R1151 B.n698 B.n450 71.676
R1152 B.n694 B.n451 71.676
R1153 B.n690 B.n452 71.676
R1154 B.n686 B.n453 71.676
R1155 B.n682 B.n454 71.676
R1156 B.n678 B.n455 71.676
R1157 B.n674 B.n456 71.676
R1158 B.n670 B.n457 71.676
R1159 B.n666 B.n458 71.676
R1160 B.n662 B.n459 71.676
R1161 B.n658 B.n460 71.676
R1162 B.n654 B.n461 71.676
R1163 B.n650 B.n462 71.676
R1164 B.n646 B.n463 71.676
R1165 B.n642 B.n464 71.676
R1166 B.n638 B.n465 71.676
R1167 B.n634 B.n466 71.676
R1168 B.n630 B.n467 71.676
R1169 B.n626 B.n468 71.676
R1170 B.n622 B.n469 71.676
R1171 B.n618 B.n470 71.676
R1172 B.n614 B.n471 71.676
R1173 B.n610 B.n472 71.676
R1174 B.n605 B.n473 71.676
R1175 B.n601 B.n474 71.676
R1176 B.n597 B.n475 71.676
R1177 B.n593 B.n476 71.676
R1178 B.n589 B.n477 71.676
R1179 B.n585 B.n478 71.676
R1180 B.n581 B.n479 71.676
R1181 B.n577 B.n480 71.676
R1182 B.n573 B.n481 71.676
R1183 B.n569 B.n482 71.676
R1184 B.n565 B.n483 71.676
R1185 B.n561 B.n484 71.676
R1186 B.n557 B.n485 71.676
R1187 B.n553 B.n486 71.676
R1188 B.n549 B.n487 71.676
R1189 B.n545 B.n488 71.676
R1190 B.n541 B.n489 71.676
R1191 B.n537 B.n490 71.676
R1192 B.n533 B.n491 71.676
R1193 B.n529 B.n492 71.676
R1194 B.n525 B.n493 71.676
R1195 B.n521 B.n494 71.676
R1196 B.n517 B.n495 71.676
R1197 B.n513 B.n496 71.676
R1198 B.n509 B.n497 71.676
R1199 B.n505 B.n498 71.676
R1200 B.n504 B.t16 69.2055
R1201 B.n139 B.t14 69.2055
R1202 B.n501 B.t6 69.1857
R1203 B.n142 B.t11 69.1857
R1204 B.n723 B.n441 68.7336
R1205 B.n911 B.n78 68.7336
R1206 B.n607 B.n504 59.5399
R1207 B.n502 B.n501 59.5399
R1208 B.n241 B.n142 59.5399
R1209 B.n140 B.n139 59.5399
R1210 B.n730 B.n441 36.8025
R1211 B.n730 B.n437 36.8025
R1212 B.n736 B.n437 36.8025
R1213 B.n736 B.n433 36.8025
R1214 B.n742 B.n433 36.8025
R1215 B.n742 B.n429 36.8025
R1216 B.n748 B.n429 36.8025
R1217 B.n748 B.n425 36.8025
R1218 B.n754 B.n425 36.8025
R1219 B.n760 B.n421 36.8025
R1220 B.n760 B.n417 36.8025
R1221 B.n766 B.n417 36.8025
R1222 B.n766 B.n413 36.8025
R1223 B.n772 B.n413 36.8025
R1224 B.n772 B.n409 36.8025
R1225 B.n778 B.n409 36.8025
R1226 B.n778 B.n405 36.8025
R1227 B.n784 B.n405 36.8025
R1228 B.n784 B.n401 36.8025
R1229 B.n790 B.n401 36.8025
R1230 B.n790 B.n397 36.8025
R1231 B.n796 B.n397 36.8025
R1232 B.n802 B.n393 36.8025
R1233 B.n802 B.n389 36.8025
R1234 B.n808 B.n389 36.8025
R1235 B.n808 B.n385 36.8025
R1236 B.n814 B.n385 36.8025
R1237 B.n814 B.n381 36.8025
R1238 B.n820 B.n381 36.8025
R1239 B.n820 B.n377 36.8025
R1240 B.n826 B.n377 36.8025
R1241 B.n826 B.n373 36.8025
R1242 B.n832 B.n373 36.8025
R1243 B.n838 B.n369 36.8025
R1244 B.n838 B.n365 36.8025
R1245 B.n845 B.n365 36.8025
R1246 B.n845 B.n361 36.8025
R1247 B.n851 B.n361 36.8025
R1248 B.n851 B.n4 36.8025
R1249 B.n1000 B.n4 36.8025
R1250 B.n1000 B.n999 36.8025
R1251 B.n999 B.n998 36.8025
R1252 B.n998 B.n8 36.8025
R1253 B.n992 B.n8 36.8025
R1254 B.n992 B.n991 36.8025
R1255 B.n991 B.n990 36.8025
R1256 B.n990 B.n15 36.8025
R1257 B.n984 B.n983 36.8025
R1258 B.n983 B.n982 36.8025
R1259 B.n982 B.n22 36.8025
R1260 B.n976 B.n22 36.8025
R1261 B.n976 B.n975 36.8025
R1262 B.n975 B.n974 36.8025
R1263 B.n974 B.n29 36.8025
R1264 B.n968 B.n29 36.8025
R1265 B.n968 B.n967 36.8025
R1266 B.n967 B.n966 36.8025
R1267 B.n966 B.n36 36.8025
R1268 B.n960 B.n959 36.8025
R1269 B.n959 B.n958 36.8025
R1270 B.n958 B.n43 36.8025
R1271 B.n952 B.n43 36.8025
R1272 B.n952 B.n951 36.8025
R1273 B.n951 B.n950 36.8025
R1274 B.n950 B.n50 36.8025
R1275 B.n944 B.n50 36.8025
R1276 B.n944 B.n943 36.8025
R1277 B.n943 B.n942 36.8025
R1278 B.n942 B.n57 36.8025
R1279 B.n936 B.n57 36.8025
R1280 B.n936 B.n935 36.8025
R1281 B.n934 B.n64 36.8025
R1282 B.n928 B.n64 36.8025
R1283 B.n928 B.n927 36.8025
R1284 B.n927 B.n926 36.8025
R1285 B.n926 B.n71 36.8025
R1286 B.n920 B.n71 36.8025
R1287 B.n920 B.n919 36.8025
R1288 B.n919 B.n918 36.8025
R1289 B.n918 B.n78 36.8025
R1290 B.t5 B.n421 34.0964
R1291 B.n796 B.t3 34.0964
R1292 B.n960 B.t0 34.0964
R1293 B.n935 B.t9 34.0964
R1294 B.n915 B.n914 31.6883
R1295 B.n909 B.n908 31.6883
R1296 B.n506 B.n439 31.6883
R1297 B.n727 B.n726 31.6883
R1298 B.n832 B.t2 21.1075
R1299 B.n984 B.t1 21.1075
R1300 B B.n1002 18.0485
R1301 B.t2 B.n369 15.6955
R1302 B.t1 B.n15 15.6955
R1303 B.n914 B.n80 10.6151
R1304 B.n144 B.n80 10.6151
R1305 B.n145 B.n144 10.6151
R1306 B.n148 B.n145 10.6151
R1307 B.n149 B.n148 10.6151
R1308 B.n152 B.n149 10.6151
R1309 B.n153 B.n152 10.6151
R1310 B.n156 B.n153 10.6151
R1311 B.n157 B.n156 10.6151
R1312 B.n160 B.n157 10.6151
R1313 B.n161 B.n160 10.6151
R1314 B.n164 B.n161 10.6151
R1315 B.n165 B.n164 10.6151
R1316 B.n168 B.n165 10.6151
R1317 B.n169 B.n168 10.6151
R1318 B.n172 B.n169 10.6151
R1319 B.n173 B.n172 10.6151
R1320 B.n176 B.n173 10.6151
R1321 B.n177 B.n176 10.6151
R1322 B.n180 B.n177 10.6151
R1323 B.n181 B.n180 10.6151
R1324 B.n184 B.n181 10.6151
R1325 B.n185 B.n184 10.6151
R1326 B.n188 B.n185 10.6151
R1327 B.n189 B.n188 10.6151
R1328 B.n192 B.n189 10.6151
R1329 B.n193 B.n192 10.6151
R1330 B.n196 B.n193 10.6151
R1331 B.n197 B.n196 10.6151
R1332 B.n200 B.n197 10.6151
R1333 B.n201 B.n200 10.6151
R1334 B.n204 B.n201 10.6151
R1335 B.n205 B.n204 10.6151
R1336 B.n208 B.n205 10.6151
R1337 B.n209 B.n208 10.6151
R1338 B.n212 B.n209 10.6151
R1339 B.n213 B.n212 10.6151
R1340 B.n216 B.n213 10.6151
R1341 B.n217 B.n216 10.6151
R1342 B.n220 B.n217 10.6151
R1343 B.n221 B.n220 10.6151
R1344 B.n224 B.n221 10.6151
R1345 B.n225 B.n224 10.6151
R1346 B.n228 B.n225 10.6151
R1347 B.n229 B.n228 10.6151
R1348 B.n232 B.n229 10.6151
R1349 B.n233 B.n232 10.6151
R1350 B.n236 B.n233 10.6151
R1351 B.n237 B.n236 10.6151
R1352 B.n240 B.n237 10.6151
R1353 B.n245 B.n242 10.6151
R1354 B.n246 B.n245 10.6151
R1355 B.n249 B.n246 10.6151
R1356 B.n250 B.n249 10.6151
R1357 B.n253 B.n250 10.6151
R1358 B.n254 B.n253 10.6151
R1359 B.n257 B.n254 10.6151
R1360 B.n258 B.n257 10.6151
R1361 B.n262 B.n261 10.6151
R1362 B.n265 B.n262 10.6151
R1363 B.n266 B.n265 10.6151
R1364 B.n269 B.n266 10.6151
R1365 B.n270 B.n269 10.6151
R1366 B.n273 B.n270 10.6151
R1367 B.n274 B.n273 10.6151
R1368 B.n277 B.n274 10.6151
R1369 B.n278 B.n277 10.6151
R1370 B.n281 B.n278 10.6151
R1371 B.n282 B.n281 10.6151
R1372 B.n285 B.n282 10.6151
R1373 B.n286 B.n285 10.6151
R1374 B.n289 B.n286 10.6151
R1375 B.n290 B.n289 10.6151
R1376 B.n293 B.n290 10.6151
R1377 B.n294 B.n293 10.6151
R1378 B.n297 B.n294 10.6151
R1379 B.n298 B.n297 10.6151
R1380 B.n301 B.n298 10.6151
R1381 B.n302 B.n301 10.6151
R1382 B.n305 B.n302 10.6151
R1383 B.n306 B.n305 10.6151
R1384 B.n309 B.n306 10.6151
R1385 B.n310 B.n309 10.6151
R1386 B.n313 B.n310 10.6151
R1387 B.n314 B.n313 10.6151
R1388 B.n317 B.n314 10.6151
R1389 B.n318 B.n317 10.6151
R1390 B.n321 B.n318 10.6151
R1391 B.n322 B.n321 10.6151
R1392 B.n325 B.n322 10.6151
R1393 B.n326 B.n325 10.6151
R1394 B.n329 B.n326 10.6151
R1395 B.n330 B.n329 10.6151
R1396 B.n333 B.n330 10.6151
R1397 B.n334 B.n333 10.6151
R1398 B.n337 B.n334 10.6151
R1399 B.n338 B.n337 10.6151
R1400 B.n341 B.n338 10.6151
R1401 B.n342 B.n341 10.6151
R1402 B.n345 B.n342 10.6151
R1403 B.n346 B.n345 10.6151
R1404 B.n349 B.n346 10.6151
R1405 B.n350 B.n349 10.6151
R1406 B.n353 B.n350 10.6151
R1407 B.n354 B.n353 10.6151
R1408 B.n357 B.n354 10.6151
R1409 B.n358 B.n357 10.6151
R1410 B.n909 B.n358 10.6151
R1411 B.n732 B.n439 10.6151
R1412 B.n733 B.n732 10.6151
R1413 B.n734 B.n733 10.6151
R1414 B.n734 B.n431 10.6151
R1415 B.n744 B.n431 10.6151
R1416 B.n745 B.n744 10.6151
R1417 B.n746 B.n745 10.6151
R1418 B.n746 B.n423 10.6151
R1419 B.n756 B.n423 10.6151
R1420 B.n757 B.n756 10.6151
R1421 B.n758 B.n757 10.6151
R1422 B.n758 B.n415 10.6151
R1423 B.n768 B.n415 10.6151
R1424 B.n769 B.n768 10.6151
R1425 B.n770 B.n769 10.6151
R1426 B.n770 B.n407 10.6151
R1427 B.n780 B.n407 10.6151
R1428 B.n781 B.n780 10.6151
R1429 B.n782 B.n781 10.6151
R1430 B.n782 B.n399 10.6151
R1431 B.n792 B.n399 10.6151
R1432 B.n793 B.n792 10.6151
R1433 B.n794 B.n793 10.6151
R1434 B.n794 B.n391 10.6151
R1435 B.n804 B.n391 10.6151
R1436 B.n805 B.n804 10.6151
R1437 B.n806 B.n805 10.6151
R1438 B.n806 B.n383 10.6151
R1439 B.n816 B.n383 10.6151
R1440 B.n817 B.n816 10.6151
R1441 B.n818 B.n817 10.6151
R1442 B.n818 B.n375 10.6151
R1443 B.n828 B.n375 10.6151
R1444 B.n829 B.n828 10.6151
R1445 B.n830 B.n829 10.6151
R1446 B.n830 B.n367 10.6151
R1447 B.n840 B.n367 10.6151
R1448 B.n841 B.n840 10.6151
R1449 B.n843 B.n841 10.6151
R1450 B.n843 B.n842 10.6151
R1451 B.n842 B.n359 10.6151
R1452 B.n854 B.n359 10.6151
R1453 B.n855 B.n854 10.6151
R1454 B.n856 B.n855 10.6151
R1455 B.n857 B.n856 10.6151
R1456 B.n859 B.n857 10.6151
R1457 B.n860 B.n859 10.6151
R1458 B.n861 B.n860 10.6151
R1459 B.n862 B.n861 10.6151
R1460 B.n864 B.n862 10.6151
R1461 B.n865 B.n864 10.6151
R1462 B.n866 B.n865 10.6151
R1463 B.n867 B.n866 10.6151
R1464 B.n869 B.n867 10.6151
R1465 B.n870 B.n869 10.6151
R1466 B.n871 B.n870 10.6151
R1467 B.n872 B.n871 10.6151
R1468 B.n874 B.n872 10.6151
R1469 B.n875 B.n874 10.6151
R1470 B.n876 B.n875 10.6151
R1471 B.n877 B.n876 10.6151
R1472 B.n879 B.n877 10.6151
R1473 B.n880 B.n879 10.6151
R1474 B.n881 B.n880 10.6151
R1475 B.n882 B.n881 10.6151
R1476 B.n884 B.n882 10.6151
R1477 B.n885 B.n884 10.6151
R1478 B.n886 B.n885 10.6151
R1479 B.n887 B.n886 10.6151
R1480 B.n889 B.n887 10.6151
R1481 B.n890 B.n889 10.6151
R1482 B.n891 B.n890 10.6151
R1483 B.n892 B.n891 10.6151
R1484 B.n894 B.n892 10.6151
R1485 B.n895 B.n894 10.6151
R1486 B.n896 B.n895 10.6151
R1487 B.n897 B.n896 10.6151
R1488 B.n899 B.n897 10.6151
R1489 B.n900 B.n899 10.6151
R1490 B.n901 B.n900 10.6151
R1491 B.n902 B.n901 10.6151
R1492 B.n904 B.n902 10.6151
R1493 B.n905 B.n904 10.6151
R1494 B.n906 B.n905 10.6151
R1495 B.n907 B.n906 10.6151
R1496 B.n908 B.n907 10.6151
R1497 B.n726 B.n443 10.6151
R1498 B.n721 B.n443 10.6151
R1499 B.n721 B.n720 10.6151
R1500 B.n720 B.n719 10.6151
R1501 B.n719 B.n716 10.6151
R1502 B.n716 B.n715 10.6151
R1503 B.n715 B.n712 10.6151
R1504 B.n712 B.n711 10.6151
R1505 B.n711 B.n708 10.6151
R1506 B.n708 B.n707 10.6151
R1507 B.n707 B.n704 10.6151
R1508 B.n704 B.n703 10.6151
R1509 B.n703 B.n700 10.6151
R1510 B.n700 B.n699 10.6151
R1511 B.n699 B.n696 10.6151
R1512 B.n696 B.n695 10.6151
R1513 B.n695 B.n692 10.6151
R1514 B.n692 B.n691 10.6151
R1515 B.n691 B.n688 10.6151
R1516 B.n688 B.n687 10.6151
R1517 B.n687 B.n684 10.6151
R1518 B.n684 B.n683 10.6151
R1519 B.n683 B.n680 10.6151
R1520 B.n680 B.n679 10.6151
R1521 B.n679 B.n676 10.6151
R1522 B.n676 B.n675 10.6151
R1523 B.n675 B.n672 10.6151
R1524 B.n672 B.n671 10.6151
R1525 B.n671 B.n668 10.6151
R1526 B.n668 B.n667 10.6151
R1527 B.n667 B.n664 10.6151
R1528 B.n664 B.n663 10.6151
R1529 B.n663 B.n660 10.6151
R1530 B.n660 B.n659 10.6151
R1531 B.n659 B.n656 10.6151
R1532 B.n656 B.n655 10.6151
R1533 B.n655 B.n652 10.6151
R1534 B.n652 B.n651 10.6151
R1535 B.n651 B.n648 10.6151
R1536 B.n648 B.n647 10.6151
R1537 B.n647 B.n644 10.6151
R1538 B.n644 B.n643 10.6151
R1539 B.n643 B.n640 10.6151
R1540 B.n640 B.n639 10.6151
R1541 B.n639 B.n636 10.6151
R1542 B.n636 B.n635 10.6151
R1543 B.n635 B.n632 10.6151
R1544 B.n632 B.n631 10.6151
R1545 B.n631 B.n628 10.6151
R1546 B.n628 B.n627 10.6151
R1547 B.n624 B.n623 10.6151
R1548 B.n623 B.n620 10.6151
R1549 B.n620 B.n619 10.6151
R1550 B.n619 B.n616 10.6151
R1551 B.n616 B.n615 10.6151
R1552 B.n615 B.n612 10.6151
R1553 B.n612 B.n611 10.6151
R1554 B.n611 B.n608 10.6151
R1555 B.n606 B.n603 10.6151
R1556 B.n603 B.n602 10.6151
R1557 B.n602 B.n599 10.6151
R1558 B.n599 B.n598 10.6151
R1559 B.n598 B.n595 10.6151
R1560 B.n595 B.n594 10.6151
R1561 B.n594 B.n591 10.6151
R1562 B.n591 B.n590 10.6151
R1563 B.n590 B.n587 10.6151
R1564 B.n587 B.n586 10.6151
R1565 B.n586 B.n583 10.6151
R1566 B.n583 B.n582 10.6151
R1567 B.n582 B.n579 10.6151
R1568 B.n579 B.n578 10.6151
R1569 B.n578 B.n575 10.6151
R1570 B.n575 B.n574 10.6151
R1571 B.n574 B.n571 10.6151
R1572 B.n571 B.n570 10.6151
R1573 B.n570 B.n567 10.6151
R1574 B.n567 B.n566 10.6151
R1575 B.n566 B.n563 10.6151
R1576 B.n563 B.n562 10.6151
R1577 B.n562 B.n559 10.6151
R1578 B.n559 B.n558 10.6151
R1579 B.n558 B.n555 10.6151
R1580 B.n555 B.n554 10.6151
R1581 B.n554 B.n551 10.6151
R1582 B.n551 B.n550 10.6151
R1583 B.n550 B.n547 10.6151
R1584 B.n547 B.n546 10.6151
R1585 B.n546 B.n543 10.6151
R1586 B.n543 B.n542 10.6151
R1587 B.n542 B.n539 10.6151
R1588 B.n539 B.n538 10.6151
R1589 B.n538 B.n535 10.6151
R1590 B.n535 B.n534 10.6151
R1591 B.n534 B.n531 10.6151
R1592 B.n531 B.n530 10.6151
R1593 B.n530 B.n527 10.6151
R1594 B.n527 B.n526 10.6151
R1595 B.n526 B.n523 10.6151
R1596 B.n523 B.n522 10.6151
R1597 B.n522 B.n519 10.6151
R1598 B.n519 B.n518 10.6151
R1599 B.n518 B.n515 10.6151
R1600 B.n515 B.n514 10.6151
R1601 B.n514 B.n511 10.6151
R1602 B.n511 B.n510 10.6151
R1603 B.n510 B.n507 10.6151
R1604 B.n507 B.n506 10.6151
R1605 B.n728 B.n727 10.6151
R1606 B.n728 B.n435 10.6151
R1607 B.n738 B.n435 10.6151
R1608 B.n739 B.n738 10.6151
R1609 B.n740 B.n739 10.6151
R1610 B.n740 B.n427 10.6151
R1611 B.n750 B.n427 10.6151
R1612 B.n751 B.n750 10.6151
R1613 B.n752 B.n751 10.6151
R1614 B.n752 B.n419 10.6151
R1615 B.n762 B.n419 10.6151
R1616 B.n763 B.n762 10.6151
R1617 B.n764 B.n763 10.6151
R1618 B.n764 B.n411 10.6151
R1619 B.n774 B.n411 10.6151
R1620 B.n775 B.n774 10.6151
R1621 B.n776 B.n775 10.6151
R1622 B.n776 B.n403 10.6151
R1623 B.n786 B.n403 10.6151
R1624 B.n787 B.n786 10.6151
R1625 B.n788 B.n787 10.6151
R1626 B.n788 B.n395 10.6151
R1627 B.n798 B.n395 10.6151
R1628 B.n799 B.n798 10.6151
R1629 B.n800 B.n799 10.6151
R1630 B.n800 B.n387 10.6151
R1631 B.n810 B.n387 10.6151
R1632 B.n811 B.n810 10.6151
R1633 B.n812 B.n811 10.6151
R1634 B.n812 B.n379 10.6151
R1635 B.n822 B.n379 10.6151
R1636 B.n823 B.n822 10.6151
R1637 B.n824 B.n823 10.6151
R1638 B.n824 B.n371 10.6151
R1639 B.n834 B.n371 10.6151
R1640 B.n835 B.n834 10.6151
R1641 B.n836 B.n835 10.6151
R1642 B.n836 B.n363 10.6151
R1643 B.n847 B.n363 10.6151
R1644 B.n848 B.n847 10.6151
R1645 B.n849 B.n848 10.6151
R1646 B.n849 B.n0 10.6151
R1647 B.n996 B.n1 10.6151
R1648 B.n996 B.n995 10.6151
R1649 B.n995 B.n994 10.6151
R1650 B.n994 B.n10 10.6151
R1651 B.n988 B.n10 10.6151
R1652 B.n988 B.n987 10.6151
R1653 B.n987 B.n986 10.6151
R1654 B.n986 B.n17 10.6151
R1655 B.n980 B.n17 10.6151
R1656 B.n980 B.n979 10.6151
R1657 B.n979 B.n978 10.6151
R1658 B.n978 B.n24 10.6151
R1659 B.n972 B.n24 10.6151
R1660 B.n972 B.n971 10.6151
R1661 B.n971 B.n970 10.6151
R1662 B.n970 B.n31 10.6151
R1663 B.n964 B.n31 10.6151
R1664 B.n964 B.n963 10.6151
R1665 B.n963 B.n962 10.6151
R1666 B.n962 B.n38 10.6151
R1667 B.n956 B.n38 10.6151
R1668 B.n956 B.n955 10.6151
R1669 B.n955 B.n954 10.6151
R1670 B.n954 B.n45 10.6151
R1671 B.n948 B.n45 10.6151
R1672 B.n948 B.n947 10.6151
R1673 B.n947 B.n946 10.6151
R1674 B.n946 B.n52 10.6151
R1675 B.n940 B.n52 10.6151
R1676 B.n940 B.n939 10.6151
R1677 B.n939 B.n938 10.6151
R1678 B.n938 B.n59 10.6151
R1679 B.n932 B.n59 10.6151
R1680 B.n932 B.n931 10.6151
R1681 B.n931 B.n930 10.6151
R1682 B.n930 B.n66 10.6151
R1683 B.n924 B.n66 10.6151
R1684 B.n924 B.n923 10.6151
R1685 B.n923 B.n922 10.6151
R1686 B.n922 B.n73 10.6151
R1687 B.n916 B.n73 10.6151
R1688 B.n916 B.n915 10.6151
R1689 B.n242 B.n241 6.5566
R1690 B.n258 B.n140 6.5566
R1691 B.n624 B.n502 6.5566
R1692 B.n608 B.n607 6.5566
R1693 B.n241 B.n240 4.05904
R1694 B.n261 B.n140 4.05904
R1695 B.n627 B.n502 4.05904
R1696 B.n607 B.n606 4.05904
R1697 B.n1002 B.n0 2.81026
R1698 B.n1002 B.n1 2.81026
R1699 B.n754 B.t5 2.70653
R1700 B.t3 B.n393 2.70653
R1701 B.t0 B.n36 2.70653
R1702 B.t9 B.n934 2.70653
R1703 VP.n19 VP.n18 161.3
R1704 VP.n17 VP.n1 161.3
R1705 VP.n16 VP.n15 161.3
R1706 VP.n14 VP.n2 161.3
R1707 VP.n13 VP.n12 161.3
R1708 VP.n11 VP.n3 161.3
R1709 VP.n10 VP.n9 161.3
R1710 VP.n8 VP.n4 161.3
R1711 VP.n5 VP.t3 134.905
R1712 VP.n5 VP.t0 133.654
R1713 VP.n6 VP.t1 99.9192
R1714 VP.n0 VP.t2 99.9192
R1715 VP.n7 VP.n6 78.8126
R1716 VP.n20 VP.n0 78.8126
R1717 VP.n12 VP.n2 56.5193
R1718 VP.n7 VP.n5 53.968
R1719 VP.n10 VP.n4 24.4675
R1720 VP.n11 VP.n10 24.4675
R1721 VP.n12 VP.n11 24.4675
R1722 VP.n16 VP.n2 24.4675
R1723 VP.n17 VP.n16 24.4675
R1724 VP.n18 VP.n17 24.4675
R1725 VP.n6 VP.n4 11.2553
R1726 VP.n18 VP.n0 11.2553
R1727 VP.n8 VP.n7 0.354971
R1728 VP.n20 VP.n19 0.354971
R1729 VP VP.n20 0.26696
R1730 VP.n9 VP.n8 0.189894
R1731 VP.n9 VP.n3 0.189894
R1732 VP.n13 VP.n3 0.189894
R1733 VP.n14 VP.n13 0.189894
R1734 VP.n15 VP.n14 0.189894
R1735 VP.n15 VP.n1 0.189894
R1736 VP.n19 VP.n1 0.189894
R1737 VTAIL.n5 VTAIL.t5 46.4863
R1738 VTAIL.n4 VTAIL.t1 46.4863
R1739 VTAIL.n3 VTAIL.t3 46.4863
R1740 VTAIL.n7 VTAIL.t2 46.4861
R1741 VTAIL.n0 VTAIL.t0 46.4861
R1742 VTAIL.n1 VTAIL.t7 46.4861
R1743 VTAIL.n2 VTAIL.t4 46.4861
R1744 VTAIL.n6 VTAIL.t6 46.4861
R1745 VTAIL.n7 VTAIL.n6 28.7548
R1746 VTAIL.n3 VTAIL.n2 28.7548
R1747 VTAIL.n4 VTAIL.n3 3.41429
R1748 VTAIL.n6 VTAIL.n5 3.41429
R1749 VTAIL.n2 VTAIL.n1 3.41429
R1750 VTAIL VTAIL.n0 1.76559
R1751 VTAIL VTAIL.n7 1.64921
R1752 VTAIL.n5 VTAIL.n4 0.470328
R1753 VTAIL.n1 VTAIL.n0 0.470328
R1754 VDD1 VDD1.n1 109.305
R1755 VDD1 VDD1.n0 61.9075
R1756 VDD1.n0 VDD1.t0 1.31611
R1757 VDD1.n0 VDD1.t3 1.31611
R1758 VDD1.n1 VDD1.t2 1.31611
R1759 VDD1.n1 VDD1.t1 1.31611
R1760 VN.n1 VN.t0 134.905
R1761 VN.n0 VN.t3 134.905
R1762 VN.n1 VN.t2 133.654
R1763 VN.n0 VN.t1 133.654
R1764 VN VN.n1 54.1333
R1765 VN VN.n0 2.06893
R1766 VDD2.n2 VDD2.n0 108.779
R1767 VDD2.n2 VDD2.n1 61.8493
R1768 VDD2.n1 VDD2.t1 1.31611
R1769 VDD2.n1 VDD2.t3 1.31611
R1770 VDD2.n0 VDD2.t0 1.31611
R1771 VDD2.n0 VDD2.t2 1.31611
R1772 VDD2 VDD2.n2 0.0586897
C0 VTAIL VDD1 6.33019f
C1 VP VTAIL 6.12396f
C2 VN VDD2 6.18797f
C3 VN VDD1 0.150083f
C4 VP VN 7.49583f
C5 VDD2 VDD1 1.27546f
C6 VP VDD2 0.459998f
C7 VN VTAIL 6.10985f
C8 VP VDD1 6.49688f
C9 VTAIL VDD2 6.3913f
C10 VDD2 B 4.591511f
C11 VDD1 B 9.398971f
C12 VTAIL B 12.493767f
C13 VN B 12.91463f
C14 VP B 11.32685f
C15 VDD2.t0 B 0.320705f
C16 VDD2.t2 B 0.320705f
C17 VDD2.n0 B 3.74463f
C18 VDD2.t1 B 0.320705f
C19 VDD2.t3 B 0.320705f
C20 VDD2.n1 B 2.90044f
C21 VDD2.n2 B 4.36967f
C22 VN.t1 B 3.25821f
C23 VN.t3 B 3.26867f
C24 VN.n0 B 1.95986f
C25 VN.t0 B 3.26867f
C26 VN.t2 B 3.25821f
C27 VN.n1 B 3.31255f
C28 VDD1.t0 B 0.323241f
C29 VDD1.t3 B 0.323241f
C30 VDD1.n0 B 2.92388f
C31 VDD1.t2 B 0.323241f
C32 VDD1.t1 B 0.323241f
C33 VDD1.n1 B 3.80275f
C34 VTAIL.t0 B 2.16738f
C35 VTAIL.n0 B 0.332311f
C36 VTAIL.t7 B 2.16738f
C37 VTAIL.n1 B 0.41855f
C38 VTAIL.t4 B 2.16738f
C39 VTAIL.n2 B 1.47169f
C40 VTAIL.t3 B 2.16738f
C41 VTAIL.n3 B 1.47169f
C42 VTAIL.t1 B 2.16738f
C43 VTAIL.n4 B 0.418548f
C44 VTAIL.t5 B 2.16738f
C45 VTAIL.n5 B 0.418548f
C46 VTAIL.t6 B 2.16738f
C47 VTAIL.n6 B 1.47169f
C48 VTAIL.t2 B 2.16738f
C49 VTAIL.n7 B 1.37937f
C50 VP.t2 B 3.01003f
C51 VP.n0 B 1.12637f
C52 VP.n1 B 0.020105f
C53 VP.n2 B 0.02935f
C54 VP.n3 B 0.020105f
C55 VP.n4 B 0.027482f
C56 VP.t3 B 3.32286f
C57 VP.t0 B 3.31223f
C58 VP.n5 B 3.35949f
C59 VP.t1 B 3.01003f
C60 VP.n6 B 1.12637f
C61 VP.n7 B 1.28431f
C62 VP.n8 B 0.03245f
C63 VP.n9 B 0.020105f
C64 VP.n10 B 0.037472f
C65 VP.n11 B 0.037472f
C66 VP.n12 B 0.02935f
C67 VP.n13 B 0.020105f
C68 VP.n14 B 0.020105f
C69 VP.n15 B 0.020105f
C70 VP.n16 B 0.037472f
C71 VP.n17 B 0.037472f
C72 VP.n18 B 0.027482f
C73 VP.n19 B 0.03245f
C74 VP.n20 B 0.054274f
.ends

