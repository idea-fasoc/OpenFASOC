* NGSPICE file created from diff_pair_sample_0058.ext - technology: sky130A

.subckt diff_pair_sample_0058 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t10 VN.t0 VDD2.t1 B.t5 sky130_fd_pr__nfet_01v8 ad=2.06415 pd=12.84 as=2.06415 ps=12.84 w=12.51 l=1.45
X1 VDD1.t5 VP.t0 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=2.06415 pd=12.84 as=4.8789 ps=25.8 w=12.51 l=1.45
X2 B.t19 B.t17 B.t18 B.t11 sky130_fd_pr__nfet_01v8 ad=4.8789 pd=25.8 as=0 ps=0 w=12.51 l=1.45
X3 B.t16 B.t14 B.t15 B.t7 sky130_fd_pr__nfet_01v8 ad=4.8789 pd=25.8 as=0 ps=0 w=12.51 l=1.45
X4 VDD2.t2 VN.t1 VTAIL.t9 B.t4 sky130_fd_pr__nfet_01v8 ad=4.8789 pd=25.8 as=2.06415 ps=12.84 w=12.51 l=1.45
X5 VTAIL.t8 VN.t2 VDD2.t5 B.t0 sky130_fd_pr__nfet_01v8 ad=2.06415 pd=12.84 as=2.06415 ps=12.84 w=12.51 l=1.45
X6 B.t13 B.t10 B.t12 B.t11 sky130_fd_pr__nfet_01v8 ad=4.8789 pd=25.8 as=0 ps=0 w=12.51 l=1.45
X7 VDD2.t3 VN.t3 VTAIL.t7 B.t1 sky130_fd_pr__nfet_01v8 ad=2.06415 pd=12.84 as=4.8789 ps=25.8 w=12.51 l=1.45
X8 VDD2.t4 VN.t4 VTAIL.t6 B.t2 sky130_fd_pr__nfet_01v8 ad=4.8789 pd=25.8 as=2.06415 ps=12.84 w=12.51 l=1.45
X9 VTAIL.t11 VP.t1 VDD1.t4 B.t5 sky130_fd_pr__nfet_01v8 ad=2.06415 pd=12.84 as=2.06415 ps=12.84 w=12.51 l=1.45
X10 VDD1.t3 VP.t2 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=4.8789 pd=25.8 as=2.06415 ps=12.84 w=12.51 l=1.45
X11 VDD1.t2 VP.t3 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=2.06415 pd=12.84 as=4.8789 ps=25.8 w=12.51 l=1.45
X12 VDD1.t1 VP.t4 VTAIL.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=4.8789 pd=25.8 as=2.06415 ps=12.84 w=12.51 l=1.45
X13 VTAIL.t0 VP.t5 VDD1.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=2.06415 pd=12.84 as=2.06415 ps=12.84 w=12.51 l=1.45
X14 B.t9 B.t6 B.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=4.8789 pd=25.8 as=0 ps=0 w=12.51 l=1.45
X15 VDD2.t0 VN.t5 VTAIL.t5 B.t3 sky130_fd_pr__nfet_01v8 ad=2.06415 pd=12.84 as=4.8789 ps=25.8 w=12.51 l=1.45
R0 VN.n3 VN.t1 244.256
R1 VN.n13 VN.t3 244.256
R2 VN.n2 VN.t0 207.925
R3 VN.n8 VN.t5 207.925
R4 VN.n12 VN.t2 207.925
R5 VN.n18 VN.t4 207.925
R6 VN.n9 VN.n8 172.065
R7 VN.n19 VN.n18 172.065
R8 VN.n17 VN.n10 161.3
R9 VN.n16 VN.n15 161.3
R10 VN.n14 VN.n11 161.3
R11 VN.n7 VN.n0 161.3
R12 VN.n6 VN.n5 161.3
R13 VN.n4 VN.n1 161.3
R14 VN.n6 VN.n1 51.1773
R15 VN.n16 VN.n11 51.1773
R16 VN VN.n19 44.9039
R17 VN.n3 VN.n2 41.8525
R18 VN.n13 VN.n12 41.8525
R19 VN.n7 VN.n6 29.8095
R20 VN.n17 VN.n16 29.8095
R21 VN.n2 VN.n1 24.4675
R22 VN.n12 VN.n11 24.4675
R23 VN.n14 VN.n13 17.3787
R24 VN.n4 VN.n3 17.3787
R25 VN.n8 VN.n7 13.702
R26 VN.n18 VN.n17 13.702
R27 VN.n19 VN.n10 0.189894
R28 VN.n15 VN.n10 0.189894
R29 VN.n15 VN.n14 0.189894
R30 VN.n5 VN.n4 0.189894
R31 VN.n5 VN.n0 0.189894
R32 VN.n9 VN.n0 0.189894
R33 VN VN.n9 0.0516364
R34 VDD2.n1 VDD2.t2 65.0474
R35 VDD2.n2 VDD2.t4 63.952
R36 VDD2.n1 VDD2.n0 62.6974
R37 VDD2 VDD2.n3 62.6946
R38 VDD2.n2 VDD2.n1 39.4868
R39 VDD2.n3 VDD2.t5 1.58323
R40 VDD2.n3 VDD2.t3 1.58323
R41 VDD2.n0 VDD2.t1 1.58323
R42 VDD2.n0 VDD2.t0 1.58323
R43 VDD2 VDD2.n2 1.20955
R44 VTAIL.n7 VTAIL.t7 47.2732
R45 VTAIL.n11 VTAIL.t5 47.2731
R46 VTAIL.n2 VTAIL.t1 47.2731
R47 VTAIL.n10 VTAIL.t3 47.2731
R48 VTAIL.n9 VTAIL.n8 45.6906
R49 VTAIL.n6 VTAIL.n5 45.6906
R50 VTAIL.n1 VTAIL.n0 45.6903
R51 VTAIL.n4 VTAIL.n3 45.6903
R52 VTAIL.n6 VTAIL.n4 26.2203
R53 VTAIL.n11 VTAIL.n10 24.6858
R54 VTAIL.n0 VTAIL.t9 1.58323
R55 VTAIL.n0 VTAIL.t10 1.58323
R56 VTAIL.n3 VTAIL.t2 1.58323
R57 VTAIL.n3 VTAIL.t0 1.58323
R58 VTAIL.n8 VTAIL.t4 1.58323
R59 VTAIL.n8 VTAIL.t11 1.58323
R60 VTAIL.n5 VTAIL.t6 1.58323
R61 VTAIL.n5 VTAIL.t8 1.58323
R62 VTAIL.n7 VTAIL.n6 1.53498
R63 VTAIL.n10 VTAIL.n9 1.53498
R64 VTAIL.n4 VTAIL.n2 1.53498
R65 VTAIL.n9 VTAIL.n7 1.23757
R66 VTAIL.n2 VTAIL.n1 1.23757
R67 VTAIL VTAIL.n11 1.09317
R68 VTAIL VTAIL.n1 0.44231
R69 B.n725 B.n724 585
R70 B.n298 B.n103 585
R71 B.n297 B.n296 585
R72 B.n295 B.n294 585
R73 B.n293 B.n292 585
R74 B.n291 B.n290 585
R75 B.n289 B.n288 585
R76 B.n287 B.n286 585
R77 B.n285 B.n284 585
R78 B.n283 B.n282 585
R79 B.n281 B.n280 585
R80 B.n279 B.n278 585
R81 B.n277 B.n276 585
R82 B.n275 B.n274 585
R83 B.n273 B.n272 585
R84 B.n271 B.n270 585
R85 B.n269 B.n268 585
R86 B.n267 B.n266 585
R87 B.n265 B.n264 585
R88 B.n263 B.n262 585
R89 B.n261 B.n260 585
R90 B.n259 B.n258 585
R91 B.n257 B.n256 585
R92 B.n255 B.n254 585
R93 B.n253 B.n252 585
R94 B.n251 B.n250 585
R95 B.n249 B.n248 585
R96 B.n247 B.n246 585
R97 B.n245 B.n244 585
R98 B.n243 B.n242 585
R99 B.n241 B.n240 585
R100 B.n239 B.n238 585
R101 B.n237 B.n236 585
R102 B.n235 B.n234 585
R103 B.n233 B.n232 585
R104 B.n231 B.n230 585
R105 B.n229 B.n228 585
R106 B.n227 B.n226 585
R107 B.n225 B.n224 585
R108 B.n223 B.n222 585
R109 B.n221 B.n220 585
R110 B.n219 B.n218 585
R111 B.n217 B.n216 585
R112 B.n214 B.n213 585
R113 B.n212 B.n211 585
R114 B.n210 B.n209 585
R115 B.n208 B.n207 585
R116 B.n206 B.n205 585
R117 B.n204 B.n203 585
R118 B.n202 B.n201 585
R119 B.n200 B.n199 585
R120 B.n198 B.n197 585
R121 B.n196 B.n195 585
R122 B.n193 B.n192 585
R123 B.n191 B.n190 585
R124 B.n189 B.n188 585
R125 B.n187 B.n186 585
R126 B.n185 B.n184 585
R127 B.n183 B.n182 585
R128 B.n181 B.n180 585
R129 B.n179 B.n178 585
R130 B.n177 B.n176 585
R131 B.n175 B.n174 585
R132 B.n173 B.n172 585
R133 B.n171 B.n170 585
R134 B.n169 B.n168 585
R135 B.n167 B.n166 585
R136 B.n165 B.n164 585
R137 B.n163 B.n162 585
R138 B.n161 B.n160 585
R139 B.n159 B.n158 585
R140 B.n157 B.n156 585
R141 B.n155 B.n154 585
R142 B.n153 B.n152 585
R143 B.n151 B.n150 585
R144 B.n149 B.n148 585
R145 B.n147 B.n146 585
R146 B.n145 B.n144 585
R147 B.n143 B.n142 585
R148 B.n141 B.n140 585
R149 B.n139 B.n138 585
R150 B.n137 B.n136 585
R151 B.n135 B.n134 585
R152 B.n133 B.n132 585
R153 B.n131 B.n130 585
R154 B.n129 B.n128 585
R155 B.n127 B.n126 585
R156 B.n125 B.n124 585
R157 B.n123 B.n122 585
R158 B.n121 B.n120 585
R159 B.n119 B.n118 585
R160 B.n117 B.n116 585
R161 B.n115 B.n114 585
R162 B.n113 B.n112 585
R163 B.n111 B.n110 585
R164 B.n109 B.n108 585
R165 B.n723 B.n55 585
R166 B.n728 B.n55 585
R167 B.n722 B.n54 585
R168 B.n729 B.n54 585
R169 B.n721 B.n720 585
R170 B.n720 B.n50 585
R171 B.n719 B.n49 585
R172 B.n735 B.n49 585
R173 B.n718 B.n48 585
R174 B.n736 B.n48 585
R175 B.n717 B.n47 585
R176 B.n737 B.n47 585
R177 B.n716 B.n715 585
R178 B.n715 B.n43 585
R179 B.n714 B.n42 585
R180 B.n743 B.n42 585
R181 B.n713 B.n41 585
R182 B.n744 B.n41 585
R183 B.n712 B.n40 585
R184 B.n745 B.n40 585
R185 B.n711 B.n710 585
R186 B.n710 B.n36 585
R187 B.n709 B.n35 585
R188 B.n751 B.n35 585
R189 B.n708 B.n34 585
R190 B.n752 B.n34 585
R191 B.n707 B.n33 585
R192 B.n753 B.n33 585
R193 B.n706 B.n705 585
R194 B.n705 B.n32 585
R195 B.n704 B.n28 585
R196 B.n759 B.n28 585
R197 B.n703 B.n27 585
R198 B.n760 B.n27 585
R199 B.n702 B.n26 585
R200 B.n761 B.n26 585
R201 B.n701 B.n700 585
R202 B.n700 B.n22 585
R203 B.n699 B.n21 585
R204 B.n767 B.n21 585
R205 B.n698 B.n20 585
R206 B.n768 B.n20 585
R207 B.n697 B.n19 585
R208 B.n769 B.n19 585
R209 B.n696 B.n695 585
R210 B.n695 B.n15 585
R211 B.n694 B.n14 585
R212 B.n775 B.n14 585
R213 B.n693 B.n13 585
R214 B.n776 B.n13 585
R215 B.n692 B.n12 585
R216 B.n777 B.n12 585
R217 B.n691 B.n690 585
R218 B.n690 B.n8 585
R219 B.n689 B.n7 585
R220 B.n783 B.n7 585
R221 B.n688 B.n6 585
R222 B.n784 B.n6 585
R223 B.n687 B.n5 585
R224 B.n785 B.n5 585
R225 B.n686 B.n685 585
R226 B.n685 B.n4 585
R227 B.n684 B.n299 585
R228 B.n684 B.n683 585
R229 B.n674 B.n300 585
R230 B.n301 B.n300 585
R231 B.n676 B.n675 585
R232 B.n677 B.n676 585
R233 B.n673 B.n305 585
R234 B.n309 B.n305 585
R235 B.n672 B.n671 585
R236 B.n671 B.n670 585
R237 B.n307 B.n306 585
R238 B.n308 B.n307 585
R239 B.n663 B.n662 585
R240 B.n664 B.n663 585
R241 B.n661 B.n314 585
R242 B.n314 B.n313 585
R243 B.n660 B.n659 585
R244 B.n659 B.n658 585
R245 B.n316 B.n315 585
R246 B.n317 B.n316 585
R247 B.n651 B.n650 585
R248 B.n652 B.n651 585
R249 B.n649 B.n322 585
R250 B.n322 B.n321 585
R251 B.n648 B.n647 585
R252 B.n647 B.n646 585
R253 B.n324 B.n323 585
R254 B.n639 B.n324 585
R255 B.n638 B.n637 585
R256 B.n640 B.n638 585
R257 B.n636 B.n329 585
R258 B.n329 B.n328 585
R259 B.n635 B.n634 585
R260 B.n634 B.n633 585
R261 B.n331 B.n330 585
R262 B.n332 B.n331 585
R263 B.n626 B.n625 585
R264 B.n627 B.n626 585
R265 B.n624 B.n337 585
R266 B.n337 B.n336 585
R267 B.n623 B.n622 585
R268 B.n622 B.n621 585
R269 B.n339 B.n338 585
R270 B.n340 B.n339 585
R271 B.n614 B.n613 585
R272 B.n615 B.n614 585
R273 B.n612 B.n345 585
R274 B.n345 B.n344 585
R275 B.n611 B.n610 585
R276 B.n610 B.n609 585
R277 B.n347 B.n346 585
R278 B.n348 B.n347 585
R279 B.n602 B.n601 585
R280 B.n603 B.n602 585
R281 B.n600 B.n353 585
R282 B.n353 B.n352 585
R283 B.n595 B.n594 585
R284 B.n593 B.n403 585
R285 B.n592 B.n402 585
R286 B.n597 B.n402 585
R287 B.n591 B.n590 585
R288 B.n589 B.n588 585
R289 B.n587 B.n586 585
R290 B.n585 B.n584 585
R291 B.n583 B.n582 585
R292 B.n581 B.n580 585
R293 B.n579 B.n578 585
R294 B.n577 B.n576 585
R295 B.n575 B.n574 585
R296 B.n573 B.n572 585
R297 B.n571 B.n570 585
R298 B.n569 B.n568 585
R299 B.n567 B.n566 585
R300 B.n565 B.n564 585
R301 B.n563 B.n562 585
R302 B.n561 B.n560 585
R303 B.n559 B.n558 585
R304 B.n557 B.n556 585
R305 B.n555 B.n554 585
R306 B.n553 B.n552 585
R307 B.n551 B.n550 585
R308 B.n549 B.n548 585
R309 B.n547 B.n546 585
R310 B.n545 B.n544 585
R311 B.n543 B.n542 585
R312 B.n541 B.n540 585
R313 B.n539 B.n538 585
R314 B.n537 B.n536 585
R315 B.n535 B.n534 585
R316 B.n533 B.n532 585
R317 B.n531 B.n530 585
R318 B.n529 B.n528 585
R319 B.n527 B.n526 585
R320 B.n525 B.n524 585
R321 B.n523 B.n522 585
R322 B.n521 B.n520 585
R323 B.n519 B.n518 585
R324 B.n517 B.n516 585
R325 B.n515 B.n514 585
R326 B.n513 B.n512 585
R327 B.n511 B.n510 585
R328 B.n509 B.n508 585
R329 B.n507 B.n506 585
R330 B.n505 B.n504 585
R331 B.n503 B.n502 585
R332 B.n501 B.n500 585
R333 B.n499 B.n498 585
R334 B.n497 B.n496 585
R335 B.n495 B.n494 585
R336 B.n493 B.n492 585
R337 B.n491 B.n490 585
R338 B.n489 B.n488 585
R339 B.n487 B.n486 585
R340 B.n485 B.n484 585
R341 B.n483 B.n482 585
R342 B.n481 B.n480 585
R343 B.n479 B.n478 585
R344 B.n477 B.n476 585
R345 B.n475 B.n474 585
R346 B.n473 B.n472 585
R347 B.n471 B.n470 585
R348 B.n469 B.n468 585
R349 B.n467 B.n466 585
R350 B.n465 B.n464 585
R351 B.n463 B.n462 585
R352 B.n461 B.n460 585
R353 B.n459 B.n458 585
R354 B.n457 B.n456 585
R355 B.n455 B.n454 585
R356 B.n453 B.n452 585
R357 B.n451 B.n450 585
R358 B.n449 B.n448 585
R359 B.n447 B.n446 585
R360 B.n445 B.n444 585
R361 B.n443 B.n442 585
R362 B.n441 B.n440 585
R363 B.n439 B.n438 585
R364 B.n437 B.n436 585
R365 B.n435 B.n434 585
R366 B.n433 B.n432 585
R367 B.n431 B.n430 585
R368 B.n429 B.n428 585
R369 B.n427 B.n426 585
R370 B.n425 B.n424 585
R371 B.n423 B.n422 585
R372 B.n421 B.n420 585
R373 B.n419 B.n418 585
R374 B.n417 B.n416 585
R375 B.n415 B.n414 585
R376 B.n413 B.n412 585
R377 B.n411 B.n410 585
R378 B.n355 B.n354 585
R379 B.n599 B.n598 585
R380 B.n598 B.n597 585
R381 B.n351 B.n350 585
R382 B.n352 B.n351 585
R383 B.n605 B.n604 585
R384 B.n604 B.n603 585
R385 B.n606 B.n349 585
R386 B.n349 B.n348 585
R387 B.n608 B.n607 585
R388 B.n609 B.n608 585
R389 B.n343 B.n342 585
R390 B.n344 B.n343 585
R391 B.n617 B.n616 585
R392 B.n616 B.n615 585
R393 B.n618 B.n341 585
R394 B.n341 B.n340 585
R395 B.n620 B.n619 585
R396 B.n621 B.n620 585
R397 B.n335 B.n334 585
R398 B.n336 B.n335 585
R399 B.n629 B.n628 585
R400 B.n628 B.n627 585
R401 B.n630 B.n333 585
R402 B.n333 B.n332 585
R403 B.n632 B.n631 585
R404 B.n633 B.n632 585
R405 B.n327 B.n326 585
R406 B.n328 B.n327 585
R407 B.n642 B.n641 585
R408 B.n641 B.n640 585
R409 B.n643 B.n325 585
R410 B.n639 B.n325 585
R411 B.n645 B.n644 585
R412 B.n646 B.n645 585
R413 B.n320 B.n319 585
R414 B.n321 B.n320 585
R415 B.n654 B.n653 585
R416 B.n653 B.n652 585
R417 B.n655 B.n318 585
R418 B.n318 B.n317 585
R419 B.n657 B.n656 585
R420 B.n658 B.n657 585
R421 B.n312 B.n311 585
R422 B.n313 B.n312 585
R423 B.n666 B.n665 585
R424 B.n665 B.n664 585
R425 B.n667 B.n310 585
R426 B.n310 B.n308 585
R427 B.n669 B.n668 585
R428 B.n670 B.n669 585
R429 B.n304 B.n303 585
R430 B.n309 B.n304 585
R431 B.n679 B.n678 585
R432 B.n678 B.n677 585
R433 B.n680 B.n302 585
R434 B.n302 B.n301 585
R435 B.n682 B.n681 585
R436 B.n683 B.n682 585
R437 B.n2 B.n0 585
R438 B.n4 B.n2 585
R439 B.n3 B.n1 585
R440 B.n784 B.n3 585
R441 B.n782 B.n781 585
R442 B.n783 B.n782 585
R443 B.n780 B.n9 585
R444 B.n9 B.n8 585
R445 B.n779 B.n778 585
R446 B.n778 B.n777 585
R447 B.n11 B.n10 585
R448 B.n776 B.n11 585
R449 B.n774 B.n773 585
R450 B.n775 B.n774 585
R451 B.n772 B.n16 585
R452 B.n16 B.n15 585
R453 B.n771 B.n770 585
R454 B.n770 B.n769 585
R455 B.n18 B.n17 585
R456 B.n768 B.n18 585
R457 B.n766 B.n765 585
R458 B.n767 B.n766 585
R459 B.n764 B.n23 585
R460 B.n23 B.n22 585
R461 B.n763 B.n762 585
R462 B.n762 B.n761 585
R463 B.n25 B.n24 585
R464 B.n760 B.n25 585
R465 B.n758 B.n757 585
R466 B.n759 B.n758 585
R467 B.n756 B.n29 585
R468 B.n32 B.n29 585
R469 B.n755 B.n754 585
R470 B.n754 B.n753 585
R471 B.n31 B.n30 585
R472 B.n752 B.n31 585
R473 B.n750 B.n749 585
R474 B.n751 B.n750 585
R475 B.n748 B.n37 585
R476 B.n37 B.n36 585
R477 B.n747 B.n746 585
R478 B.n746 B.n745 585
R479 B.n39 B.n38 585
R480 B.n744 B.n39 585
R481 B.n742 B.n741 585
R482 B.n743 B.n742 585
R483 B.n740 B.n44 585
R484 B.n44 B.n43 585
R485 B.n739 B.n738 585
R486 B.n738 B.n737 585
R487 B.n46 B.n45 585
R488 B.n736 B.n46 585
R489 B.n734 B.n733 585
R490 B.n735 B.n734 585
R491 B.n732 B.n51 585
R492 B.n51 B.n50 585
R493 B.n731 B.n730 585
R494 B.n730 B.n729 585
R495 B.n53 B.n52 585
R496 B.n728 B.n53 585
R497 B.n787 B.n786 585
R498 B.n786 B.n785 585
R499 B.n595 B.n351 492.5
R500 B.n108 B.n53 492.5
R501 B.n598 B.n353 492.5
R502 B.n725 B.n55 492.5
R503 B.n407 B.t10 413.173
R504 B.n404 B.t17 413.173
R505 B.n106 B.t14 413.173
R506 B.n104 B.t6 413.173
R507 B.n727 B.n726 256.663
R508 B.n727 B.n102 256.663
R509 B.n727 B.n101 256.663
R510 B.n727 B.n100 256.663
R511 B.n727 B.n99 256.663
R512 B.n727 B.n98 256.663
R513 B.n727 B.n97 256.663
R514 B.n727 B.n96 256.663
R515 B.n727 B.n95 256.663
R516 B.n727 B.n94 256.663
R517 B.n727 B.n93 256.663
R518 B.n727 B.n92 256.663
R519 B.n727 B.n91 256.663
R520 B.n727 B.n90 256.663
R521 B.n727 B.n89 256.663
R522 B.n727 B.n88 256.663
R523 B.n727 B.n87 256.663
R524 B.n727 B.n86 256.663
R525 B.n727 B.n85 256.663
R526 B.n727 B.n84 256.663
R527 B.n727 B.n83 256.663
R528 B.n727 B.n82 256.663
R529 B.n727 B.n81 256.663
R530 B.n727 B.n80 256.663
R531 B.n727 B.n79 256.663
R532 B.n727 B.n78 256.663
R533 B.n727 B.n77 256.663
R534 B.n727 B.n76 256.663
R535 B.n727 B.n75 256.663
R536 B.n727 B.n74 256.663
R537 B.n727 B.n73 256.663
R538 B.n727 B.n72 256.663
R539 B.n727 B.n71 256.663
R540 B.n727 B.n70 256.663
R541 B.n727 B.n69 256.663
R542 B.n727 B.n68 256.663
R543 B.n727 B.n67 256.663
R544 B.n727 B.n66 256.663
R545 B.n727 B.n65 256.663
R546 B.n727 B.n64 256.663
R547 B.n727 B.n63 256.663
R548 B.n727 B.n62 256.663
R549 B.n727 B.n61 256.663
R550 B.n727 B.n60 256.663
R551 B.n727 B.n59 256.663
R552 B.n727 B.n58 256.663
R553 B.n727 B.n57 256.663
R554 B.n727 B.n56 256.663
R555 B.n597 B.n596 256.663
R556 B.n597 B.n356 256.663
R557 B.n597 B.n357 256.663
R558 B.n597 B.n358 256.663
R559 B.n597 B.n359 256.663
R560 B.n597 B.n360 256.663
R561 B.n597 B.n361 256.663
R562 B.n597 B.n362 256.663
R563 B.n597 B.n363 256.663
R564 B.n597 B.n364 256.663
R565 B.n597 B.n365 256.663
R566 B.n597 B.n366 256.663
R567 B.n597 B.n367 256.663
R568 B.n597 B.n368 256.663
R569 B.n597 B.n369 256.663
R570 B.n597 B.n370 256.663
R571 B.n597 B.n371 256.663
R572 B.n597 B.n372 256.663
R573 B.n597 B.n373 256.663
R574 B.n597 B.n374 256.663
R575 B.n597 B.n375 256.663
R576 B.n597 B.n376 256.663
R577 B.n597 B.n377 256.663
R578 B.n597 B.n378 256.663
R579 B.n597 B.n379 256.663
R580 B.n597 B.n380 256.663
R581 B.n597 B.n381 256.663
R582 B.n597 B.n382 256.663
R583 B.n597 B.n383 256.663
R584 B.n597 B.n384 256.663
R585 B.n597 B.n385 256.663
R586 B.n597 B.n386 256.663
R587 B.n597 B.n387 256.663
R588 B.n597 B.n388 256.663
R589 B.n597 B.n389 256.663
R590 B.n597 B.n390 256.663
R591 B.n597 B.n391 256.663
R592 B.n597 B.n392 256.663
R593 B.n597 B.n393 256.663
R594 B.n597 B.n394 256.663
R595 B.n597 B.n395 256.663
R596 B.n597 B.n396 256.663
R597 B.n597 B.n397 256.663
R598 B.n597 B.n398 256.663
R599 B.n597 B.n399 256.663
R600 B.n597 B.n400 256.663
R601 B.n597 B.n401 256.663
R602 B.n604 B.n351 163.367
R603 B.n604 B.n349 163.367
R604 B.n608 B.n349 163.367
R605 B.n608 B.n343 163.367
R606 B.n616 B.n343 163.367
R607 B.n616 B.n341 163.367
R608 B.n620 B.n341 163.367
R609 B.n620 B.n335 163.367
R610 B.n628 B.n335 163.367
R611 B.n628 B.n333 163.367
R612 B.n632 B.n333 163.367
R613 B.n632 B.n327 163.367
R614 B.n641 B.n327 163.367
R615 B.n641 B.n325 163.367
R616 B.n645 B.n325 163.367
R617 B.n645 B.n320 163.367
R618 B.n653 B.n320 163.367
R619 B.n653 B.n318 163.367
R620 B.n657 B.n318 163.367
R621 B.n657 B.n312 163.367
R622 B.n665 B.n312 163.367
R623 B.n665 B.n310 163.367
R624 B.n669 B.n310 163.367
R625 B.n669 B.n304 163.367
R626 B.n678 B.n304 163.367
R627 B.n678 B.n302 163.367
R628 B.n682 B.n302 163.367
R629 B.n682 B.n2 163.367
R630 B.n786 B.n2 163.367
R631 B.n786 B.n3 163.367
R632 B.n782 B.n3 163.367
R633 B.n782 B.n9 163.367
R634 B.n778 B.n9 163.367
R635 B.n778 B.n11 163.367
R636 B.n774 B.n11 163.367
R637 B.n774 B.n16 163.367
R638 B.n770 B.n16 163.367
R639 B.n770 B.n18 163.367
R640 B.n766 B.n18 163.367
R641 B.n766 B.n23 163.367
R642 B.n762 B.n23 163.367
R643 B.n762 B.n25 163.367
R644 B.n758 B.n25 163.367
R645 B.n758 B.n29 163.367
R646 B.n754 B.n29 163.367
R647 B.n754 B.n31 163.367
R648 B.n750 B.n31 163.367
R649 B.n750 B.n37 163.367
R650 B.n746 B.n37 163.367
R651 B.n746 B.n39 163.367
R652 B.n742 B.n39 163.367
R653 B.n742 B.n44 163.367
R654 B.n738 B.n44 163.367
R655 B.n738 B.n46 163.367
R656 B.n734 B.n46 163.367
R657 B.n734 B.n51 163.367
R658 B.n730 B.n51 163.367
R659 B.n730 B.n53 163.367
R660 B.n403 B.n402 163.367
R661 B.n590 B.n402 163.367
R662 B.n588 B.n587 163.367
R663 B.n584 B.n583 163.367
R664 B.n580 B.n579 163.367
R665 B.n576 B.n575 163.367
R666 B.n572 B.n571 163.367
R667 B.n568 B.n567 163.367
R668 B.n564 B.n563 163.367
R669 B.n560 B.n559 163.367
R670 B.n556 B.n555 163.367
R671 B.n552 B.n551 163.367
R672 B.n548 B.n547 163.367
R673 B.n544 B.n543 163.367
R674 B.n540 B.n539 163.367
R675 B.n536 B.n535 163.367
R676 B.n532 B.n531 163.367
R677 B.n528 B.n527 163.367
R678 B.n524 B.n523 163.367
R679 B.n520 B.n519 163.367
R680 B.n516 B.n515 163.367
R681 B.n512 B.n511 163.367
R682 B.n508 B.n507 163.367
R683 B.n504 B.n503 163.367
R684 B.n500 B.n499 163.367
R685 B.n496 B.n495 163.367
R686 B.n492 B.n491 163.367
R687 B.n488 B.n487 163.367
R688 B.n484 B.n483 163.367
R689 B.n480 B.n479 163.367
R690 B.n476 B.n475 163.367
R691 B.n472 B.n471 163.367
R692 B.n468 B.n467 163.367
R693 B.n464 B.n463 163.367
R694 B.n460 B.n459 163.367
R695 B.n456 B.n455 163.367
R696 B.n452 B.n451 163.367
R697 B.n448 B.n447 163.367
R698 B.n444 B.n443 163.367
R699 B.n440 B.n439 163.367
R700 B.n436 B.n435 163.367
R701 B.n432 B.n431 163.367
R702 B.n428 B.n427 163.367
R703 B.n424 B.n423 163.367
R704 B.n420 B.n419 163.367
R705 B.n416 B.n415 163.367
R706 B.n412 B.n411 163.367
R707 B.n598 B.n355 163.367
R708 B.n602 B.n353 163.367
R709 B.n602 B.n347 163.367
R710 B.n610 B.n347 163.367
R711 B.n610 B.n345 163.367
R712 B.n614 B.n345 163.367
R713 B.n614 B.n339 163.367
R714 B.n622 B.n339 163.367
R715 B.n622 B.n337 163.367
R716 B.n626 B.n337 163.367
R717 B.n626 B.n331 163.367
R718 B.n634 B.n331 163.367
R719 B.n634 B.n329 163.367
R720 B.n638 B.n329 163.367
R721 B.n638 B.n324 163.367
R722 B.n647 B.n324 163.367
R723 B.n647 B.n322 163.367
R724 B.n651 B.n322 163.367
R725 B.n651 B.n316 163.367
R726 B.n659 B.n316 163.367
R727 B.n659 B.n314 163.367
R728 B.n663 B.n314 163.367
R729 B.n663 B.n307 163.367
R730 B.n671 B.n307 163.367
R731 B.n671 B.n305 163.367
R732 B.n676 B.n305 163.367
R733 B.n676 B.n300 163.367
R734 B.n684 B.n300 163.367
R735 B.n685 B.n684 163.367
R736 B.n685 B.n5 163.367
R737 B.n6 B.n5 163.367
R738 B.n7 B.n6 163.367
R739 B.n690 B.n7 163.367
R740 B.n690 B.n12 163.367
R741 B.n13 B.n12 163.367
R742 B.n14 B.n13 163.367
R743 B.n695 B.n14 163.367
R744 B.n695 B.n19 163.367
R745 B.n20 B.n19 163.367
R746 B.n21 B.n20 163.367
R747 B.n700 B.n21 163.367
R748 B.n700 B.n26 163.367
R749 B.n27 B.n26 163.367
R750 B.n28 B.n27 163.367
R751 B.n705 B.n28 163.367
R752 B.n705 B.n33 163.367
R753 B.n34 B.n33 163.367
R754 B.n35 B.n34 163.367
R755 B.n710 B.n35 163.367
R756 B.n710 B.n40 163.367
R757 B.n41 B.n40 163.367
R758 B.n42 B.n41 163.367
R759 B.n715 B.n42 163.367
R760 B.n715 B.n47 163.367
R761 B.n48 B.n47 163.367
R762 B.n49 B.n48 163.367
R763 B.n720 B.n49 163.367
R764 B.n720 B.n54 163.367
R765 B.n55 B.n54 163.367
R766 B.n112 B.n111 163.367
R767 B.n116 B.n115 163.367
R768 B.n120 B.n119 163.367
R769 B.n124 B.n123 163.367
R770 B.n128 B.n127 163.367
R771 B.n132 B.n131 163.367
R772 B.n136 B.n135 163.367
R773 B.n140 B.n139 163.367
R774 B.n144 B.n143 163.367
R775 B.n148 B.n147 163.367
R776 B.n152 B.n151 163.367
R777 B.n156 B.n155 163.367
R778 B.n160 B.n159 163.367
R779 B.n164 B.n163 163.367
R780 B.n168 B.n167 163.367
R781 B.n172 B.n171 163.367
R782 B.n176 B.n175 163.367
R783 B.n180 B.n179 163.367
R784 B.n184 B.n183 163.367
R785 B.n188 B.n187 163.367
R786 B.n192 B.n191 163.367
R787 B.n197 B.n196 163.367
R788 B.n201 B.n200 163.367
R789 B.n205 B.n204 163.367
R790 B.n209 B.n208 163.367
R791 B.n213 B.n212 163.367
R792 B.n218 B.n217 163.367
R793 B.n222 B.n221 163.367
R794 B.n226 B.n225 163.367
R795 B.n230 B.n229 163.367
R796 B.n234 B.n233 163.367
R797 B.n238 B.n237 163.367
R798 B.n242 B.n241 163.367
R799 B.n246 B.n245 163.367
R800 B.n250 B.n249 163.367
R801 B.n254 B.n253 163.367
R802 B.n258 B.n257 163.367
R803 B.n262 B.n261 163.367
R804 B.n266 B.n265 163.367
R805 B.n270 B.n269 163.367
R806 B.n274 B.n273 163.367
R807 B.n278 B.n277 163.367
R808 B.n282 B.n281 163.367
R809 B.n286 B.n285 163.367
R810 B.n290 B.n289 163.367
R811 B.n294 B.n293 163.367
R812 B.n296 B.n103 163.367
R813 B.n407 B.t13 107.481
R814 B.n104 B.t8 107.481
R815 B.n404 B.t19 107.465
R816 B.n106 B.t15 107.465
R817 B.n597 B.n352 78.5498
R818 B.n728 B.n727 78.5498
R819 B.n408 B.t12 72.9595
R820 B.n105 B.t9 72.9595
R821 B.n405 B.t18 72.9438
R822 B.n107 B.t16 72.9438
R823 B.n596 B.n595 71.676
R824 B.n590 B.n356 71.676
R825 B.n587 B.n357 71.676
R826 B.n583 B.n358 71.676
R827 B.n579 B.n359 71.676
R828 B.n575 B.n360 71.676
R829 B.n571 B.n361 71.676
R830 B.n567 B.n362 71.676
R831 B.n563 B.n363 71.676
R832 B.n559 B.n364 71.676
R833 B.n555 B.n365 71.676
R834 B.n551 B.n366 71.676
R835 B.n547 B.n367 71.676
R836 B.n543 B.n368 71.676
R837 B.n539 B.n369 71.676
R838 B.n535 B.n370 71.676
R839 B.n531 B.n371 71.676
R840 B.n527 B.n372 71.676
R841 B.n523 B.n373 71.676
R842 B.n519 B.n374 71.676
R843 B.n515 B.n375 71.676
R844 B.n511 B.n376 71.676
R845 B.n507 B.n377 71.676
R846 B.n503 B.n378 71.676
R847 B.n499 B.n379 71.676
R848 B.n495 B.n380 71.676
R849 B.n491 B.n381 71.676
R850 B.n487 B.n382 71.676
R851 B.n483 B.n383 71.676
R852 B.n479 B.n384 71.676
R853 B.n475 B.n385 71.676
R854 B.n471 B.n386 71.676
R855 B.n467 B.n387 71.676
R856 B.n463 B.n388 71.676
R857 B.n459 B.n389 71.676
R858 B.n455 B.n390 71.676
R859 B.n451 B.n391 71.676
R860 B.n447 B.n392 71.676
R861 B.n443 B.n393 71.676
R862 B.n439 B.n394 71.676
R863 B.n435 B.n395 71.676
R864 B.n431 B.n396 71.676
R865 B.n427 B.n397 71.676
R866 B.n423 B.n398 71.676
R867 B.n419 B.n399 71.676
R868 B.n415 B.n400 71.676
R869 B.n411 B.n401 71.676
R870 B.n108 B.n56 71.676
R871 B.n112 B.n57 71.676
R872 B.n116 B.n58 71.676
R873 B.n120 B.n59 71.676
R874 B.n124 B.n60 71.676
R875 B.n128 B.n61 71.676
R876 B.n132 B.n62 71.676
R877 B.n136 B.n63 71.676
R878 B.n140 B.n64 71.676
R879 B.n144 B.n65 71.676
R880 B.n148 B.n66 71.676
R881 B.n152 B.n67 71.676
R882 B.n156 B.n68 71.676
R883 B.n160 B.n69 71.676
R884 B.n164 B.n70 71.676
R885 B.n168 B.n71 71.676
R886 B.n172 B.n72 71.676
R887 B.n176 B.n73 71.676
R888 B.n180 B.n74 71.676
R889 B.n184 B.n75 71.676
R890 B.n188 B.n76 71.676
R891 B.n192 B.n77 71.676
R892 B.n197 B.n78 71.676
R893 B.n201 B.n79 71.676
R894 B.n205 B.n80 71.676
R895 B.n209 B.n81 71.676
R896 B.n213 B.n82 71.676
R897 B.n218 B.n83 71.676
R898 B.n222 B.n84 71.676
R899 B.n226 B.n85 71.676
R900 B.n230 B.n86 71.676
R901 B.n234 B.n87 71.676
R902 B.n238 B.n88 71.676
R903 B.n242 B.n89 71.676
R904 B.n246 B.n90 71.676
R905 B.n250 B.n91 71.676
R906 B.n254 B.n92 71.676
R907 B.n258 B.n93 71.676
R908 B.n262 B.n94 71.676
R909 B.n266 B.n95 71.676
R910 B.n270 B.n96 71.676
R911 B.n274 B.n97 71.676
R912 B.n278 B.n98 71.676
R913 B.n282 B.n99 71.676
R914 B.n286 B.n100 71.676
R915 B.n290 B.n101 71.676
R916 B.n294 B.n102 71.676
R917 B.n726 B.n103 71.676
R918 B.n726 B.n725 71.676
R919 B.n296 B.n102 71.676
R920 B.n293 B.n101 71.676
R921 B.n289 B.n100 71.676
R922 B.n285 B.n99 71.676
R923 B.n281 B.n98 71.676
R924 B.n277 B.n97 71.676
R925 B.n273 B.n96 71.676
R926 B.n269 B.n95 71.676
R927 B.n265 B.n94 71.676
R928 B.n261 B.n93 71.676
R929 B.n257 B.n92 71.676
R930 B.n253 B.n91 71.676
R931 B.n249 B.n90 71.676
R932 B.n245 B.n89 71.676
R933 B.n241 B.n88 71.676
R934 B.n237 B.n87 71.676
R935 B.n233 B.n86 71.676
R936 B.n229 B.n85 71.676
R937 B.n225 B.n84 71.676
R938 B.n221 B.n83 71.676
R939 B.n217 B.n82 71.676
R940 B.n212 B.n81 71.676
R941 B.n208 B.n80 71.676
R942 B.n204 B.n79 71.676
R943 B.n200 B.n78 71.676
R944 B.n196 B.n77 71.676
R945 B.n191 B.n76 71.676
R946 B.n187 B.n75 71.676
R947 B.n183 B.n74 71.676
R948 B.n179 B.n73 71.676
R949 B.n175 B.n72 71.676
R950 B.n171 B.n71 71.676
R951 B.n167 B.n70 71.676
R952 B.n163 B.n69 71.676
R953 B.n159 B.n68 71.676
R954 B.n155 B.n67 71.676
R955 B.n151 B.n66 71.676
R956 B.n147 B.n65 71.676
R957 B.n143 B.n64 71.676
R958 B.n139 B.n63 71.676
R959 B.n135 B.n62 71.676
R960 B.n131 B.n61 71.676
R961 B.n127 B.n60 71.676
R962 B.n123 B.n59 71.676
R963 B.n119 B.n58 71.676
R964 B.n115 B.n57 71.676
R965 B.n111 B.n56 71.676
R966 B.n596 B.n403 71.676
R967 B.n588 B.n356 71.676
R968 B.n584 B.n357 71.676
R969 B.n580 B.n358 71.676
R970 B.n576 B.n359 71.676
R971 B.n572 B.n360 71.676
R972 B.n568 B.n361 71.676
R973 B.n564 B.n362 71.676
R974 B.n560 B.n363 71.676
R975 B.n556 B.n364 71.676
R976 B.n552 B.n365 71.676
R977 B.n548 B.n366 71.676
R978 B.n544 B.n367 71.676
R979 B.n540 B.n368 71.676
R980 B.n536 B.n369 71.676
R981 B.n532 B.n370 71.676
R982 B.n528 B.n371 71.676
R983 B.n524 B.n372 71.676
R984 B.n520 B.n373 71.676
R985 B.n516 B.n374 71.676
R986 B.n512 B.n375 71.676
R987 B.n508 B.n376 71.676
R988 B.n504 B.n377 71.676
R989 B.n500 B.n378 71.676
R990 B.n496 B.n379 71.676
R991 B.n492 B.n380 71.676
R992 B.n488 B.n381 71.676
R993 B.n484 B.n382 71.676
R994 B.n480 B.n383 71.676
R995 B.n476 B.n384 71.676
R996 B.n472 B.n385 71.676
R997 B.n468 B.n386 71.676
R998 B.n464 B.n387 71.676
R999 B.n460 B.n388 71.676
R1000 B.n456 B.n389 71.676
R1001 B.n452 B.n390 71.676
R1002 B.n448 B.n391 71.676
R1003 B.n444 B.n392 71.676
R1004 B.n440 B.n393 71.676
R1005 B.n436 B.n394 71.676
R1006 B.n432 B.n395 71.676
R1007 B.n428 B.n396 71.676
R1008 B.n424 B.n397 71.676
R1009 B.n420 B.n398 71.676
R1010 B.n416 B.n399 71.676
R1011 B.n412 B.n400 71.676
R1012 B.n401 B.n355 71.676
R1013 B.n409 B.n408 59.5399
R1014 B.n406 B.n405 59.5399
R1015 B.n194 B.n107 59.5399
R1016 B.n215 B.n105 59.5399
R1017 B.n603 B.n352 42.0584
R1018 B.n603 B.n348 42.0584
R1019 B.n609 B.n348 42.0584
R1020 B.n609 B.n344 42.0584
R1021 B.n615 B.n344 42.0584
R1022 B.n621 B.n340 42.0584
R1023 B.n621 B.n336 42.0584
R1024 B.n627 B.n336 42.0584
R1025 B.n627 B.n332 42.0584
R1026 B.n633 B.n332 42.0584
R1027 B.n633 B.n328 42.0584
R1028 B.n640 B.n328 42.0584
R1029 B.n640 B.n639 42.0584
R1030 B.n646 B.n321 42.0584
R1031 B.n652 B.n321 42.0584
R1032 B.n652 B.n317 42.0584
R1033 B.n658 B.n317 42.0584
R1034 B.n664 B.n313 42.0584
R1035 B.n664 B.n308 42.0584
R1036 B.n670 B.n308 42.0584
R1037 B.n670 B.n309 42.0584
R1038 B.n677 B.n301 42.0584
R1039 B.n683 B.n301 42.0584
R1040 B.n683 B.n4 42.0584
R1041 B.n785 B.n4 42.0584
R1042 B.n785 B.n784 42.0584
R1043 B.n784 B.n783 42.0584
R1044 B.n783 B.n8 42.0584
R1045 B.n777 B.n8 42.0584
R1046 B.n776 B.n775 42.0584
R1047 B.n775 B.n15 42.0584
R1048 B.n769 B.n15 42.0584
R1049 B.n769 B.n768 42.0584
R1050 B.n767 B.n22 42.0584
R1051 B.n761 B.n22 42.0584
R1052 B.n761 B.n760 42.0584
R1053 B.n760 B.n759 42.0584
R1054 B.n753 B.n32 42.0584
R1055 B.n753 B.n752 42.0584
R1056 B.n752 B.n751 42.0584
R1057 B.n751 B.n36 42.0584
R1058 B.n745 B.n36 42.0584
R1059 B.n745 B.n744 42.0584
R1060 B.n744 B.n743 42.0584
R1061 B.n743 B.n43 42.0584
R1062 B.n737 B.n736 42.0584
R1063 B.n736 B.n735 42.0584
R1064 B.n735 B.n50 42.0584
R1065 B.n729 B.n50 42.0584
R1066 B.n729 B.n728 42.0584
R1067 B.n615 B.t11 36.4919
R1068 B.n737 B.t7 36.4919
R1069 B.n408 B.n407 34.5217
R1070 B.n405 B.n404 34.5217
R1071 B.n107 B.n106 34.5217
R1072 B.n105 B.n104 34.5217
R1073 B.n309 B.t1 32.7809
R1074 B.t4 B.n776 32.7809
R1075 B.n109 B.n52 32.0005
R1076 B.n724 B.n723 32.0005
R1077 B.n600 B.n599 32.0005
R1078 B.n594 B.n350 32.0005
R1079 B.n646 B.t2 29.0699
R1080 B.n759 B.t3 29.0699
R1081 B.n658 B.t0 22.885
R1082 B.t5 B.n767 22.885
R1083 B.t0 B.n313 19.174
R1084 B.n768 B.t5 19.174
R1085 B B.n787 18.0485
R1086 B.n639 B.t2 12.989
R1087 B.n32 B.t3 12.989
R1088 B.n110 B.n109 10.6151
R1089 B.n113 B.n110 10.6151
R1090 B.n114 B.n113 10.6151
R1091 B.n117 B.n114 10.6151
R1092 B.n118 B.n117 10.6151
R1093 B.n121 B.n118 10.6151
R1094 B.n122 B.n121 10.6151
R1095 B.n125 B.n122 10.6151
R1096 B.n126 B.n125 10.6151
R1097 B.n129 B.n126 10.6151
R1098 B.n130 B.n129 10.6151
R1099 B.n133 B.n130 10.6151
R1100 B.n134 B.n133 10.6151
R1101 B.n137 B.n134 10.6151
R1102 B.n138 B.n137 10.6151
R1103 B.n141 B.n138 10.6151
R1104 B.n142 B.n141 10.6151
R1105 B.n145 B.n142 10.6151
R1106 B.n146 B.n145 10.6151
R1107 B.n149 B.n146 10.6151
R1108 B.n150 B.n149 10.6151
R1109 B.n153 B.n150 10.6151
R1110 B.n154 B.n153 10.6151
R1111 B.n157 B.n154 10.6151
R1112 B.n158 B.n157 10.6151
R1113 B.n161 B.n158 10.6151
R1114 B.n162 B.n161 10.6151
R1115 B.n165 B.n162 10.6151
R1116 B.n166 B.n165 10.6151
R1117 B.n169 B.n166 10.6151
R1118 B.n170 B.n169 10.6151
R1119 B.n173 B.n170 10.6151
R1120 B.n174 B.n173 10.6151
R1121 B.n177 B.n174 10.6151
R1122 B.n178 B.n177 10.6151
R1123 B.n181 B.n178 10.6151
R1124 B.n182 B.n181 10.6151
R1125 B.n185 B.n182 10.6151
R1126 B.n186 B.n185 10.6151
R1127 B.n189 B.n186 10.6151
R1128 B.n190 B.n189 10.6151
R1129 B.n193 B.n190 10.6151
R1130 B.n198 B.n195 10.6151
R1131 B.n199 B.n198 10.6151
R1132 B.n202 B.n199 10.6151
R1133 B.n203 B.n202 10.6151
R1134 B.n206 B.n203 10.6151
R1135 B.n207 B.n206 10.6151
R1136 B.n210 B.n207 10.6151
R1137 B.n211 B.n210 10.6151
R1138 B.n214 B.n211 10.6151
R1139 B.n219 B.n216 10.6151
R1140 B.n220 B.n219 10.6151
R1141 B.n223 B.n220 10.6151
R1142 B.n224 B.n223 10.6151
R1143 B.n227 B.n224 10.6151
R1144 B.n228 B.n227 10.6151
R1145 B.n231 B.n228 10.6151
R1146 B.n232 B.n231 10.6151
R1147 B.n235 B.n232 10.6151
R1148 B.n236 B.n235 10.6151
R1149 B.n239 B.n236 10.6151
R1150 B.n240 B.n239 10.6151
R1151 B.n243 B.n240 10.6151
R1152 B.n244 B.n243 10.6151
R1153 B.n247 B.n244 10.6151
R1154 B.n248 B.n247 10.6151
R1155 B.n251 B.n248 10.6151
R1156 B.n252 B.n251 10.6151
R1157 B.n255 B.n252 10.6151
R1158 B.n256 B.n255 10.6151
R1159 B.n259 B.n256 10.6151
R1160 B.n260 B.n259 10.6151
R1161 B.n263 B.n260 10.6151
R1162 B.n264 B.n263 10.6151
R1163 B.n267 B.n264 10.6151
R1164 B.n268 B.n267 10.6151
R1165 B.n271 B.n268 10.6151
R1166 B.n272 B.n271 10.6151
R1167 B.n275 B.n272 10.6151
R1168 B.n276 B.n275 10.6151
R1169 B.n279 B.n276 10.6151
R1170 B.n280 B.n279 10.6151
R1171 B.n283 B.n280 10.6151
R1172 B.n284 B.n283 10.6151
R1173 B.n287 B.n284 10.6151
R1174 B.n288 B.n287 10.6151
R1175 B.n291 B.n288 10.6151
R1176 B.n292 B.n291 10.6151
R1177 B.n295 B.n292 10.6151
R1178 B.n297 B.n295 10.6151
R1179 B.n298 B.n297 10.6151
R1180 B.n724 B.n298 10.6151
R1181 B.n601 B.n600 10.6151
R1182 B.n601 B.n346 10.6151
R1183 B.n611 B.n346 10.6151
R1184 B.n612 B.n611 10.6151
R1185 B.n613 B.n612 10.6151
R1186 B.n613 B.n338 10.6151
R1187 B.n623 B.n338 10.6151
R1188 B.n624 B.n623 10.6151
R1189 B.n625 B.n624 10.6151
R1190 B.n625 B.n330 10.6151
R1191 B.n635 B.n330 10.6151
R1192 B.n636 B.n635 10.6151
R1193 B.n637 B.n636 10.6151
R1194 B.n637 B.n323 10.6151
R1195 B.n648 B.n323 10.6151
R1196 B.n649 B.n648 10.6151
R1197 B.n650 B.n649 10.6151
R1198 B.n650 B.n315 10.6151
R1199 B.n660 B.n315 10.6151
R1200 B.n661 B.n660 10.6151
R1201 B.n662 B.n661 10.6151
R1202 B.n662 B.n306 10.6151
R1203 B.n672 B.n306 10.6151
R1204 B.n673 B.n672 10.6151
R1205 B.n675 B.n673 10.6151
R1206 B.n675 B.n674 10.6151
R1207 B.n674 B.n299 10.6151
R1208 B.n686 B.n299 10.6151
R1209 B.n687 B.n686 10.6151
R1210 B.n688 B.n687 10.6151
R1211 B.n689 B.n688 10.6151
R1212 B.n691 B.n689 10.6151
R1213 B.n692 B.n691 10.6151
R1214 B.n693 B.n692 10.6151
R1215 B.n694 B.n693 10.6151
R1216 B.n696 B.n694 10.6151
R1217 B.n697 B.n696 10.6151
R1218 B.n698 B.n697 10.6151
R1219 B.n699 B.n698 10.6151
R1220 B.n701 B.n699 10.6151
R1221 B.n702 B.n701 10.6151
R1222 B.n703 B.n702 10.6151
R1223 B.n704 B.n703 10.6151
R1224 B.n706 B.n704 10.6151
R1225 B.n707 B.n706 10.6151
R1226 B.n708 B.n707 10.6151
R1227 B.n709 B.n708 10.6151
R1228 B.n711 B.n709 10.6151
R1229 B.n712 B.n711 10.6151
R1230 B.n713 B.n712 10.6151
R1231 B.n714 B.n713 10.6151
R1232 B.n716 B.n714 10.6151
R1233 B.n717 B.n716 10.6151
R1234 B.n718 B.n717 10.6151
R1235 B.n719 B.n718 10.6151
R1236 B.n721 B.n719 10.6151
R1237 B.n722 B.n721 10.6151
R1238 B.n723 B.n722 10.6151
R1239 B.n594 B.n593 10.6151
R1240 B.n593 B.n592 10.6151
R1241 B.n592 B.n591 10.6151
R1242 B.n591 B.n589 10.6151
R1243 B.n589 B.n586 10.6151
R1244 B.n586 B.n585 10.6151
R1245 B.n585 B.n582 10.6151
R1246 B.n582 B.n581 10.6151
R1247 B.n581 B.n578 10.6151
R1248 B.n578 B.n577 10.6151
R1249 B.n577 B.n574 10.6151
R1250 B.n574 B.n573 10.6151
R1251 B.n573 B.n570 10.6151
R1252 B.n570 B.n569 10.6151
R1253 B.n569 B.n566 10.6151
R1254 B.n566 B.n565 10.6151
R1255 B.n565 B.n562 10.6151
R1256 B.n562 B.n561 10.6151
R1257 B.n561 B.n558 10.6151
R1258 B.n558 B.n557 10.6151
R1259 B.n557 B.n554 10.6151
R1260 B.n554 B.n553 10.6151
R1261 B.n553 B.n550 10.6151
R1262 B.n550 B.n549 10.6151
R1263 B.n549 B.n546 10.6151
R1264 B.n546 B.n545 10.6151
R1265 B.n545 B.n542 10.6151
R1266 B.n542 B.n541 10.6151
R1267 B.n541 B.n538 10.6151
R1268 B.n538 B.n537 10.6151
R1269 B.n537 B.n534 10.6151
R1270 B.n534 B.n533 10.6151
R1271 B.n533 B.n530 10.6151
R1272 B.n530 B.n529 10.6151
R1273 B.n529 B.n526 10.6151
R1274 B.n526 B.n525 10.6151
R1275 B.n525 B.n522 10.6151
R1276 B.n522 B.n521 10.6151
R1277 B.n521 B.n518 10.6151
R1278 B.n518 B.n517 10.6151
R1279 B.n517 B.n514 10.6151
R1280 B.n514 B.n513 10.6151
R1281 B.n510 B.n509 10.6151
R1282 B.n509 B.n506 10.6151
R1283 B.n506 B.n505 10.6151
R1284 B.n505 B.n502 10.6151
R1285 B.n502 B.n501 10.6151
R1286 B.n501 B.n498 10.6151
R1287 B.n498 B.n497 10.6151
R1288 B.n497 B.n494 10.6151
R1289 B.n494 B.n493 10.6151
R1290 B.n490 B.n489 10.6151
R1291 B.n489 B.n486 10.6151
R1292 B.n486 B.n485 10.6151
R1293 B.n485 B.n482 10.6151
R1294 B.n482 B.n481 10.6151
R1295 B.n481 B.n478 10.6151
R1296 B.n478 B.n477 10.6151
R1297 B.n477 B.n474 10.6151
R1298 B.n474 B.n473 10.6151
R1299 B.n473 B.n470 10.6151
R1300 B.n470 B.n469 10.6151
R1301 B.n469 B.n466 10.6151
R1302 B.n466 B.n465 10.6151
R1303 B.n465 B.n462 10.6151
R1304 B.n462 B.n461 10.6151
R1305 B.n461 B.n458 10.6151
R1306 B.n458 B.n457 10.6151
R1307 B.n457 B.n454 10.6151
R1308 B.n454 B.n453 10.6151
R1309 B.n453 B.n450 10.6151
R1310 B.n450 B.n449 10.6151
R1311 B.n449 B.n446 10.6151
R1312 B.n446 B.n445 10.6151
R1313 B.n445 B.n442 10.6151
R1314 B.n442 B.n441 10.6151
R1315 B.n441 B.n438 10.6151
R1316 B.n438 B.n437 10.6151
R1317 B.n437 B.n434 10.6151
R1318 B.n434 B.n433 10.6151
R1319 B.n433 B.n430 10.6151
R1320 B.n430 B.n429 10.6151
R1321 B.n429 B.n426 10.6151
R1322 B.n426 B.n425 10.6151
R1323 B.n425 B.n422 10.6151
R1324 B.n422 B.n421 10.6151
R1325 B.n421 B.n418 10.6151
R1326 B.n418 B.n417 10.6151
R1327 B.n417 B.n414 10.6151
R1328 B.n414 B.n413 10.6151
R1329 B.n413 B.n410 10.6151
R1330 B.n410 B.n354 10.6151
R1331 B.n599 B.n354 10.6151
R1332 B.n605 B.n350 10.6151
R1333 B.n606 B.n605 10.6151
R1334 B.n607 B.n606 10.6151
R1335 B.n607 B.n342 10.6151
R1336 B.n617 B.n342 10.6151
R1337 B.n618 B.n617 10.6151
R1338 B.n619 B.n618 10.6151
R1339 B.n619 B.n334 10.6151
R1340 B.n629 B.n334 10.6151
R1341 B.n630 B.n629 10.6151
R1342 B.n631 B.n630 10.6151
R1343 B.n631 B.n326 10.6151
R1344 B.n642 B.n326 10.6151
R1345 B.n643 B.n642 10.6151
R1346 B.n644 B.n643 10.6151
R1347 B.n644 B.n319 10.6151
R1348 B.n654 B.n319 10.6151
R1349 B.n655 B.n654 10.6151
R1350 B.n656 B.n655 10.6151
R1351 B.n656 B.n311 10.6151
R1352 B.n666 B.n311 10.6151
R1353 B.n667 B.n666 10.6151
R1354 B.n668 B.n667 10.6151
R1355 B.n668 B.n303 10.6151
R1356 B.n679 B.n303 10.6151
R1357 B.n680 B.n679 10.6151
R1358 B.n681 B.n680 10.6151
R1359 B.n681 B.n0 10.6151
R1360 B.n781 B.n1 10.6151
R1361 B.n781 B.n780 10.6151
R1362 B.n780 B.n779 10.6151
R1363 B.n779 B.n10 10.6151
R1364 B.n773 B.n10 10.6151
R1365 B.n773 B.n772 10.6151
R1366 B.n772 B.n771 10.6151
R1367 B.n771 B.n17 10.6151
R1368 B.n765 B.n17 10.6151
R1369 B.n765 B.n764 10.6151
R1370 B.n764 B.n763 10.6151
R1371 B.n763 B.n24 10.6151
R1372 B.n757 B.n24 10.6151
R1373 B.n757 B.n756 10.6151
R1374 B.n756 B.n755 10.6151
R1375 B.n755 B.n30 10.6151
R1376 B.n749 B.n30 10.6151
R1377 B.n749 B.n748 10.6151
R1378 B.n748 B.n747 10.6151
R1379 B.n747 B.n38 10.6151
R1380 B.n741 B.n38 10.6151
R1381 B.n741 B.n740 10.6151
R1382 B.n740 B.n739 10.6151
R1383 B.n739 B.n45 10.6151
R1384 B.n733 B.n45 10.6151
R1385 B.n733 B.n732 10.6151
R1386 B.n732 B.n731 10.6151
R1387 B.n731 B.n52 10.6151
R1388 B.n194 B.n193 9.36635
R1389 B.n216 B.n215 9.36635
R1390 B.n513 B.n406 9.36635
R1391 B.n490 B.n409 9.36635
R1392 B.n677 B.t1 9.27798
R1393 B.n777 B.t4 9.27798
R1394 B.t11 B.n340 5.56699
R1395 B.t7 B.n43 5.56699
R1396 B.n787 B.n0 2.81026
R1397 B.n787 B.n1 2.81026
R1398 B.n195 B.n194 1.24928
R1399 B.n215 B.n214 1.24928
R1400 B.n510 B.n406 1.24928
R1401 B.n493 B.n409 1.24928
R1402 VP.n7 VP.t4 244.256
R1403 VP.n20 VP.t5 207.925
R1404 VP.n14 VP.t2 207.925
R1405 VP.n26 VP.t0 207.925
R1406 VP.n6 VP.t1 207.925
R1407 VP.n12 VP.t3 207.925
R1408 VP.n15 VP.n14 172.065
R1409 VP.n27 VP.n26 172.065
R1410 VP.n13 VP.n12 172.065
R1411 VP.n8 VP.n5 161.3
R1412 VP.n10 VP.n9 161.3
R1413 VP.n11 VP.n4 161.3
R1414 VP.n25 VP.n0 161.3
R1415 VP.n24 VP.n23 161.3
R1416 VP.n22 VP.n1 161.3
R1417 VP.n21 VP.n20 161.3
R1418 VP.n19 VP.n2 161.3
R1419 VP.n18 VP.n17 161.3
R1420 VP.n16 VP.n3 161.3
R1421 VP.n19 VP.n18 51.1773
R1422 VP.n24 VP.n1 51.1773
R1423 VP.n10 VP.n5 51.1773
R1424 VP.n15 VP.n13 44.5232
R1425 VP.n7 VP.n6 41.8525
R1426 VP.n18 VP.n3 29.8095
R1427 VP.n25 VP.n24 29.8095
R1428 VP.n11 VP.n10 29.8095
R1429 VP.n20 VP.n19 24.4675
R1430 VP.n20 VP.n1 24.4675
R1431 VP.n6 VP.n5 24.4675
R1432 VP.n8 VP.n7 17.3787
R1433 VP.n14 VP.n3 13.702
R1434 VP.n26 VP.n25 13.702
R1435 VP.n12 VP.n11 13.702
R1436 VP.n9 VP.n8 0.189894
R1437 VP.n9 VP.n4 0.189894
R1438 VP.n13 VP.n4 0.189894
R1439 VP.n16 VP.n15 0.189894
R1440 VP.n17 VP.n16 0.189894
R1441 VP.n17 VP.n2 0.189894
R1442 VP.n21 VP.n2 0.189894
R1443 VP.n22 VP.n21 0.189894
R1444 VP.n23 VP.n22 0.189894
R1445 VP.n23 VP.n0 0.189894
R1446 VP.n27 VP.n0 0.189894
R1447 VP VP.n27 0.0516364
R1448 VDD1 VDD1.t1 65.1611
R1449 VDD1.n1 VDD1.t3 65.0474
R1450 VDD1.n1 VDD1.n0 62.6974
R1451 VDD1.n3 VDD1.n2 62.3692
R1452 VDD1.n3 VDD1.n1 40.8371
R1453 VDD1.n2 VDD1.t4 1.58323
R1454 VDD1.n2 VDD1.t2 1.58323
R1455 VDD1.n0 VDD1.t0 1.58323
R1456 VDD1.n0 VDD1.t5 1.58323
R1457 VDD1 VDD1.n3 0.325931
C0 VDD2 VN 6.048491f
C1 VN VP 5.90163f
C2 VTAIL VDD2 8.32012f
C3 VTAIL VP 5.93517f
C4 VN VDD1 0.149127f
C5 VDD2 VP 0.360974f
C6 VTAIL VDD1 8.27898f
C7 VDD2 VDD1 0.988127f
C8 VDD1 VP 6.25647f
C9 VTAIL VN 5.92073f
C10 VDD2 B 5.165182f
C11 VDD1 B 5.436512f
C12 VTAIL B 7.192953f
C13 VN B 9.68244f
C14 VP B 8.055183f
C15 VDD1.t1 B 2.48452f
C16 VDD1.t3 B 2.48381f
C17 VDD1.t0 B 0.21744f
C18 VDD1.t5 B 0.21744f
C19 VDD1.n0 B 1.94437f
C20 VDD1.n1 B 2.23325f
C21 VDD1.t4 B 0.21744f
C22 VDD1.t2 B 0.21744f
C23 VDD1.n2 B 1.94266f
C24 VDD1.n3 B 2.20489f
C25 VP.n0 B 0.033464f
C26 VP.t0 B 1.65583f
C27 VP.n1 B 0.060759f
C28 VP.n2 B 0.033464f
C29 VP.t5 B 1.65583f
C30 VP.n3 B 0.053122f
C31 VP.n4 B 0.033464f
C32 VP.t3 B 1.65583f
C33 VP.n5 B 0.060759f
C34 VP.t4 B 1.76392f
C35 VP.t1 B 1.65583f
C36 VP.n6 B 0.675353f
C37 VP.n7 B 0.665814f
C38 VP.n8 B 0.212372f
C39 VP.n9 B 0.033464f
C40 VP.n10 B 0.032642f
C41 VP.n11 B 0.053122f
C42 VP.n12 B 0.669589f
C43 VP.n13 B 1.52433f
C44 VP.t2 B 1.65583f
C45 VP.n14 B 0.669589f
C46 VP.n15 B 1.55135f
C47 VP.n16 B 0.033464f
C48 VP.n17 B 0.033464f
C49 VP.n18 B 0.032642f
C50 VP.n19 B 0.060759f
C51 VP.n20 B 0.629421f
C52 VP.n21 B 0.033464f
C53 VP.n22 B 0.033464f
C54 VP.n23 B 0.033464f
C55 VP.n24 B 0.032642f
C56 VP.n25 B 0.053122f
C57 VP.n26 B 0.669589f
C58 VP.n27 B 0.030722f
C59 VTAIL.t9 B 0.228734f
C60 VTAIL.t10 B 0.228734f
C61 VTAIL.n0 B 1.97519f
C62 VTAIL.n1 B 0.353846f
C63 VTAIL.t1 B 2.51965f
C64 VTAIL.n2 B 0.514674f
C65 VTAIL.t2 B 0.228734f
C66 VTAIL.t0 B 0.228734f
C67 VTAIL.n3 B 1.97519f
C68 VTAIL.n4 B 1.69022f
C69 VTAIL.t6 B 0.228734f
C70 VTAIL.t8 B 0.228734f
C71 VTAIL.n5 B 1.9752f
C72 VTAIL.n6 B 1.69021f
C73 VTAIL.t7 B 2.51966f
C74 VTAIL.n7 B 0.514659f
C75 VTAIL.t4 B 0.228734f
C76 VTAIL.t11 B 0.228734f
C77 VTAIL.n8 B 1.9752f
C78 VTAIL.n9 B 0.435304f
C79 VTAIL.t3 B 2.51965f
C80 VTAIL.n10 B 1.65518f
C81 VTAIL.t5 B 2.51965f
C82 VTAIL.n11 B 1.62224f
C83 VDD2.t2 B 2.44638f
C84 VDD2.t1 B 0.214164f
C85 VDD2.t0 B 0.214164f
C86 VDD2.n0 B 1.91507f
C87 VDD2.n1 B 2.11703f
C88 VDD2.t4 B 2.44098f
C89 VDD2.n2 B 2.18529f
C90 VDD2.t5 B 0.214164f
C91 VDD2.t3 B 0.214164f
C92 VDD2.n3 B 1.91504f
C93 VN.n0 B 0.032824f
C94 VN.t5 B 1.62416f
C95 VN.n1 B 0.059597f
C96 VN.t1 B 1.73019f
C97 VN.t0 B 1.62416f
C98 VN.n2 B 0.662438f
C99 VN.n3 B 0.653081f
C100 VN.n4 B 0.20831f
C101 VN.n5 B 0.032824f
C102 VN.n6 B 0.032018f
C103 VN.n7 B 0.052106f
C104 VN.n8 B 0.656784f
C105 VN.n9 B 0.030134f
C106 VN.n10 B 0.032824f
C107 VN.t4 B 1.62416f
C108 VN.n11 B 0.059597f
C109 VN.t3 B 1.73019f
C110 VN.t2 B 1.62416f
C111 VN.n12 B 0.662438f
C112 VN.n13 B 0.653081f
C113 VN.n14 B 0.20831f
C114 VN.n15 B 0.032824f
C115 VN.n16 B 0.032018f
C116 VN.n17 B 0.052106f
C117 VN.n18 B 0.656784f
C118 VN.n19 B 1.51665f
.ends

