* NGSPICE file created from diff_pair_sample_1164.ext - technology: sky130A

.subckt diff_pair_sample_1164 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t5 VP.t0 VTAIL.t7 B.t4 sky130_fd_pr__nfet_01v8 ad=3.3657 pd=18.04 as=1.42395 ps=8.96 w=8.63 l=0.74
X1 B.t19 B.t17 B.t18 B.t11 sky130_fd_pr__nfet_01v8 ad=3.3657 pd=18.04 as=0 ps=0 w=8.63 l=0.74
X2 VDD2.t5 VN.t0 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=1.42395 pd=8.96 as=3.3657 ps=18.04 w=8.63 l=0.74
X3 VDD2.t4 VN.t1 VTAIL.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=3.3657 pd=18.04 as=1.42395 ps=8.96 w=8.63 l=0.74
X4 VDD2.t3 VN.t2 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=3.3657 pd=18.04 as=1.42395 ps=8.96 w=8.63 l=0.74
X5 VTAIL.t1 VN.t3 VDD2.t2 B.t1 sky130_fd_pr__nfet_01v8 ad=1.42395 pd=8.96 as=1.42395 ps=8.96 w=8.63 l=0.74
X6 B.t16 B.t14 B.t15 B.t7 sky130_fd_pr__nfet_01v8 ad=3.3657 pd=18.04 as=0 ps=0 w=8.63 l=0.74
X7 B.t13 B.t10 B.t12 B.t11 sky130_fd_pr__nfet_01v8 ad=3.3657 pd=18.04 as=0 ps=0 w=8.63 l=0.74
X8 VDD1.t4 VP.t1 VTAIL.t6 B.t0 sky130_fd_pr__nfet_01v8 ad=1.42395 pd=8.96 as=3.3657 ps=18.04 w=8.63 l=0.74
X9 VDD1.t3 VP.t2 VTAIL.t8 B.t2 sky130_fd_pr__nfet_01v8 ad=1.42395 pd=8.96 as=3.3657 ps=18.04 w=8.63 l=0.74
X10 VDD1.t2 VP.t3 VTAIL.t5 B.t3 sky130_fd_pr__nfet_01v8 ad=3.3657 pd=18.04 as=1.42395 ps=8.96 w=8.63 l=0.74
X11 VDD2.t1 VN.t4 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=1.42395 pd=8.96 as=3.3657 ps=18.04 w=8.63 l=0.74
X12 VTAIL.t9 VP.t4 VDD1.t1 B.t5 sky130_fd_pr__nfet_01v8 ad=1.42395 pd=8.96 as=1.42395 ps=8.96 w=8.63 l=0.74
X13 VTAIL.t11 VN.t5 VDD2.t0 B.t5 sky130_fd_pr__nfet_01v8 ad=1.42395 pd=8.96 as=1.42395 ps=8.96 w=8.63 l=0.74
X14 B.t9 B.t6 B.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=3.3657 pd=18.04 as=0 ps=0 w=8.63 l=0.74
X15 VTAIL.t10 VP.t5 VDD1.t0 B.t1 sky130_fd_pr__nfet_01v8 ad=1.42395 pd=8.96 as=1.42395 ps=8.96 w=8.63 l=0.74
R0 VP.n3 VP.t3 356.839
R1 VP.n8 VP.t0 334.469
R2 VP.n12 VP.t5 334.469
R3 VP.n14 VP.t1 334.469
R4 VP.n6 VP.t2 334.469
R5 VP.n4 VP.t4 334.469
R6 VP.n15 VP.n14 161.3
R7 VP.n5 VP.n2 161.3
R8 VP.n7 VP.n6 161.3
R9 VP.n13 VP.n0 161.3
R10 VP.n12 VP.n11 161.3
R11 VP.n10 VP.n1 161.3
R12 VP.n9 VP.n8 161.3
R13 VP.n3 VP.n2 44.8655
R14 VP.n9 VP.n7 38.8452
R15 VP.n8 VP.n1 29.2126
R16 VP.n14 VP.n13 29.2126
R17 VP.n6 VP.n5 29.2126
R18 VP.n4 VP.n3 19.4959
R19 VP.n12 VP.n1 18.9884
R20 VP.n13 VP.n12 18.9884
R21 VP.n5 VP.n4 18.9884
R22 VP.n7 VP.n2 0.189894
R23 VP.n10 VP.n9 0.189894
R24 VP.n11 VP.n10 0.189894
R25 VP.n11 VP.n0 0.189894
R26 VP.n15 VP.n0 0.189894
R27 VP VP.n15 0.0516364
R28 VTAIL.n186 VTAIL.n146 289.615
R29 VTAIL.n42 VTAIL.n2 289.615
R30 VTAIL.n140 VTAIL.n100 289.615
R31 VTAIL.n92 VTAIL.n52 289.615
R32 VTAIL.n161 VTAIL.n160 185
R33 VTAIL.n158 VTAIL.n157 185
R34 VTAIL.n167 VTAIL.n166 185
R35 VTAIL.n169 VTAIL.n168 185
R36 VTAIL.n154 VTAIL.n153 185
R37 VTAIL.n175 VTAIL.n174 185
R38 VTAIL.n178 VTAIL.n177 185
R39 VTAIL.n176 VTAIL.n150 185
R40 VTAIL.n183 VTAIL.n149 185
R41 VTAIL.n185 VTAIL.n184 185
R42 VTAIL.n187 VTAIL.n186 185
R43 VTAIL.n17 VTAIL.n16 185
R44 VTAIL.n14 VTAIL.n13 185
R45 VTAIL.n23 VTAIL.n22 185
R46 VTAIL.n25 VTAIL.n24 185
R47 VTAIL.n10 VTAIL.n9 185
R48 VTAIL.n31 VTAIL.n30 185
R49 VTAIL.n34 VTAIL.n33 185
R50 VTAIL.n32 VTAIL.n6 185
R51 VTAIL.n39 VTAIL.n5 185
R52 VTAIL.n41 VTAIL.n40 185
R53 VTAIL.n43 VTAIL.n42 185
R54 VTAIL.n141 VTAIL.n140 185
R55 VTAIL.n139 VTAIL.n138 185
R56 VTAIL.n137 VTAIL.n103 185
R57 VTAIL.n107 VTAIL.n104 185
R58 VTAIL.n132 VTAIL.n131 185
R59 VTAIL.n130 VTAIL.n129 185
R60 VTAIL.n109 VTAIL.n108 185
R61 VTAIL.n124 VTAIL.n123 185
R62 VTAIL.n122 VTAIL.n121 185
R63 VTAIL.n113 VTAIL.n112 185
R64 VTAIL.n116 VTAIL.n115 185
R65 VTAIL.n93 VTAIL.n92 185
R66 VTAIL.n91 VTAIL.n90 185
R67 VTAIL.n89 VTAIL.n55 185
R68 VTAIL.n59 VTAIL.n56 185
R69 VTAIL.n84 VTAIL.n83 185
R70 VTAIL.n82 VTAIL.n81 185
R71 VTAIL.n61 VTAIL.n60 185
R72 VTAIL.n76 VTAIL.n75 185
R73 VTAIL.n74 VTAIL.n73 185
R74 VTAIL.n65 VTAIL.n64 185
R75 VTAIL.n68 VTAIL.n67 185
R76 VTAIL.t2 VTAIL.n159 149.524
R77 VTAIL.t6 VTAIL.n15 149.524
R78 VTAIL.t8 VTAIL.n114 149.524
R79 VTAIL.t0 VTAIL.n66 149.524
R80 VTAIL.n160 VTAIL.n157 104.615
R81 VTAIL.n167 VTAIL.n157 104.615
R82 VTAIL.n168 VTAIL.n167 104.615
R83 VTAIL.n168 VTAIL.n153 104.615
R84 VTAIL.n175 VTAIL.n153 104.615
R85 VTAIL.n177 VTAIL.n175 104.615
R86 VTAIL.n177 VTAIL.n176 104.615
R87 VTAIL.n176 VTAIL.n149 104.615
R88 VTAIL.n185 VTAIL.n149 104.615
R89 VTAIL.n186 VTAIL.n185 104.615
R90 VTAIL.n16 VTAIL.n13 104.615
R91 VTAIL.n23 VTAIL.n13 104.615
R92 VTAIL.n24 VTAIL.n23 104.615
R93 VTAIL.n24 VTAIL.n9 104.615
R94 VTAIL.n31 VTAIL.n9 104.615
R95 VTAIL.n33 VTAIL.n31 104.615
R96 VTAIL.n33 VTAIL.n32 104.615
R97 VTAIL.n32 VTAIL.n5 104.615
R98 VTAIL.n41 VTAIL.n5 104.615
R99 VTAIL.n42 VTAIL.n41 104.615
R100 VTAIL.n140 VTAIL.n139 104.615
R101 VTAIL.n139 VTAIL.n103 104.615
R102 VTAIL.n107 VTAIL.n103 104.615
R103 VTAIL.n131 VTAIL.n107 104.615
R104 VTAIL.n131 VTAIL.n130 104.615
R105 VTAIL.n130 VTAIL.n108 104.615
R106 VTAIL.n123 VTAIL.n108 104.615
R107 VTAIL.n123 VTAIL.n122 104.615
R108 VTAIL.n122 VTAIL.n112 104.615
R109 VTAIL.n115 VTAIL.n112 104.615
R110 VTAIL.n92 VTAIL.n91 104.615
R111 VTAIL.n91 VTAIL.n55 104.615
R112 VTAIL.n59 VTAIL.n55 104.615
R113 VTAIL.n83 VTAIL.n59 104.615
R114 VTAIL.n83 VTAIL.n82 104.615
R115 VTAIL.n82 VTAIL.n60 104.615
R116 VTAIL.n75 VTAIL.n60 104.615
R117 VTAIL.n75 VTAIL.n74 104.615
R118 VTAIL.n74 VTAIL.n64 104.615
R119 VTAIL.n67 VTAIL.n64 104.615
R120 VTAIL.n160 VTAIL.t2 52.3082
R121 VTAIL.n16 VTAIL.t6 52.3082
R122 VTAIL.n115 VTAIL.t8 52.3082
R123 VTAIL.n67 VTAIL.t0 52.3082
R124 VTAIL.n99 VTAIL.n98 48.8957
R125 VTAIL.n51 VTAIL.n50 48.8957
R126 VTAIL.n1 VTAIL.n0 48.8956
R127 VTAIL.n49 VTAIL.n48 48.8956
R128 VTAIL.n191 VTAIL.n190 34.3187
R129 VTAIL.n47 VTAIL.n46 34.3187
R130 VTAIL.n145 VTAIL.n144 34.3187
R131 VTAIL.n97 VTAIL.n96 34.3187
R132 VTAIL.n51 VTAIL.n49 21.6514
R133 VTAIL.n191 VTAIL.n145 20.7289
R134 VTAIL.n184 VTAIL.n183 13.1884
R135 VTAIL.n40 VTAIL.n39 13.1884
R136 VTAIL.n138 VTAIL.n137 13.1884
R137 VTAIL.n90 VTAIL.n89 13.1884
R138 VTAIL.n182 VTAIL.n150 12.8005
R139 VTAIL.n187 VTAIL.n148 12.8005
R140 VTAIL.n38 VTAIL.n6 12.8005
R141 VTAIL.n43 VTAIL.n4 12.8005
R142 VTAIL.n141 VTAIL.n102 12.8005
R143 VTAIL.n136 VTAIL.n104 12.8005
R144 VTAIL.n93 VTAIL.n54 12.8005
R145 VTAIL.n88 VTAIL.n56 12.8005
R146 VTAIL.n179 VTAIL.n178 12.0247
R147 VTAIL.n188 VTAIL.n146 12.0247
R148 VTAIL.n35 VTAIL.n34 12.0247
R149 VTAIL.n44 VTAIL.n2 12.0247
R150 VTAIL.n142 VTAIL.n100 12.0247
R151 VTAIL.n133 VTAIL.n132 12.0247
R152 VTAIL.n94 VTAIL.n52 12.0247
R153 VTAIL.n85 VTAIL.n84 12.0247
R154 VTAIL.n174 VTAIL.n152 11.249
R155 VTAIL.n30 VTAIL.n8 11.249
R156 VTAIL.n129 VTAIL.n106 11.249
R157 VTAIL.n81 VTAIL.n58 11.249
R158 VTAIL.n173 VTAIL.n154 10.4732
R159 VTAIL.n29 VTAIL.n10 10.4732
R160 VTAIL.n128 VTAIL.n109 10.4732
R161 VTAIL.n80 VTAIL.n61 10.4732
R162 VTAIL.n161 VTAIL.n159 10.2747
R163 VTAIL.n17 VTAIL.n15 10.2747
R164 VTAIL.n116 VTAIL.n114 10.2747
R165 VTAIL.n68 VTAIL.n66 10.2747
R166 VTAIL.n170 VTAIL.n169 9.69747
R167 VTAIL.n26 VTAIL.n25 9.69747
R168 VTAIL.n125 VTAIL.n124 9.69747
R169 VTAIL.n77 VTAIL.n76 9.69747
R170 VTAIL.n190 VTAIL.n189 9.45567
R171 VTAIL.n46 VTAIL.n45 9.45567
R172 VTAIL.n144 VTAIL.n143 9.45567
R173 VTAIL.n96 VTAIL.n95 9.45567
R174 VTAIL.n189 VTAIL.n188 9.3005
R175 VTAIL.n148 VTAIL.n147 9.3005
R176 VTAIL.n163 VTAIL.n162 9.3005
R177 VTAIL.n165 VTAIL.n164 9.3005
R178 VTAIL.n156 VTAIL.n155 9.3005
R179 VTAIL.n171 VTAIL.n170 9.3005
R180 VTAIL.n173 VTAIL.n172 9.3005
R181 VTAIL.n152 VTAIL.n151 9.3005
R182 VTAIL.n180 VTAIL.n179 9.3005
R183 VTAIL.n182 VTAIL.n181 9.3005
R184 VTAIL.n45 VTAIL.n44 9.3005
R185 VTAIL.n4 VTAIL.n3 9.3005
R186 VTAIL.n19 VTAIL.n18 9.3005
R187 VTAIL.n21 VTAIL.n20 9.3005
R188 VTAIL.n12 VTAIL.n11 9.3005
R189 VTAIL.n27 VTAIL.n26 9.3005
R190 VTAIL.n29 VTAIL.n28 9.3005
R191 VTAIL.n8 VTAIL.n7 9.3005
R192 VTAIL.n36 VTAIL.n35 9.3005
R193 VTAIL.n38 VTAIL.n37 9.3005
R194 VTAIL.n118 VTAIL.n117 9.3005
R195 VTAIL.n120 VTAIL.n119 9.3005
R196 VTAIL.n111 VTAIL.n110 9.3005
R197 VTAIL.n126 VTAIL.n125 9.3005
R198 VTAIL.n128 VTAIL.n127 9.3005
R199 VTAIL.n106 VTAIL.n105 9.3005
R200 VTAIL.n134 VTAIL.n133 9.3005
R201 VTAIL.n136 VTAIL.n135 9.3005
R202 VTAIL.n143 VTAIL.n142 9.3005
R203 VTAIL.n102 VTAIL.n101 9.3005
R204 VTAIL.n70 VTAIL.n69 9.3005
R205 VTAIL.n72 VTAIL.n71 9.3005
R206 VTAIL.n63 VTAIL.n62 9.3005
R207 VTAIL.n78 VTAIL.n77 9.3005
R208 VTAIL.n80 VTAIL.n79 9.3005
R209 VTAIL.n58 VTAIL.n57 9.3005
R210 VTAIL.n86 VTAIL.n85 9.3005
R211 VTAIL.n88 VTAIL.n87 9.3005
R212 VTAIL.n95 VTAIL.n94 9.3005
R213 VTAIL.n54 VTAIL.n53 9.3005
R214 VTAIL.n166 VTAIL.n156 8.92171
R215 VTAIL.n22 VTAIL.n12 8.92171
R216 VTAIL.n121 VTAIL.n111 8.92171
R217 VTAIL.n73 VTAIL.n63 8.92171
R218 VTAIL.n165 VTAIL.n158 8.14595
R219 VTAIL.n21 VTAIL.n14 8.14595
R220 VTAIL.n120 VTAIL.n113 8.14595
R221 VTAIL.n72 VTAIL.n65 8.14595
R222 VTAIL.n162 VTAIL.n161 7.3702
R223 VTAIL.n18 VTAIL.n17 7.3702
R224 VTAIL.n117 VTAIL.n116 7.3702
R225 VTAIL.n69 VTAIL.n68 7.3702
R226 VTAIL.n162 VTAIL.n158 5.81868
R227 VTAIL.n18 VTAIL.n14 5.81868
R228 VTAIL.n117 VTAIL.n113 5.81868
R229 VTAIL.n69 VTAIL.n65 5.81868
R230 VTAIL.n166 VTAIL.n165 5.04292
R231 VTAIL.n22 VTAIL.n21 5.04292
R232 VTAIL.n121 VTAIL.n120 5.04292
R233 VTAIL.n73 VTAIL.n72 5.04292
R234 VTAIL.n169 VTAIL.n156 4.26717
R235 VTAIL.n25 VTAIL.n12 4.26717
R236 VTAIL.n124 VTAIL.n111 4.26717
R237 VTAIL.n76 VTAIL.n63 4.26717
R238 VTAIL.n170 VTAIL.n154 3.49141
R239 VTAIL.n26 VTAIL.n10 3.49141
R240 VTAIL.n125 VTAIL.n109 3.49141
R241 VTAIL.n77 VTAIL.n61 3.49141
R242 VTAIL.n163 VTAIL.n159 2.84303
R243 VTAIL.n19 VTAIL.n15 2.84303
R244 VTAIL.n118 VTAIL.n114 2.84303
R245 VTAIL.n70 VTAIL.n66 2.84303
R246 VTAIL.n174 VTAIL.n173 2.71565
R247 VTAIL.n30 VTAIL.n29 2.71565
R248 VTAIL.n129 VTAIL.n128 2.71565
R249 VTAIL.n81 VTAIL.n80 2.71565
R250 VTAIL.n0 VTAIL.t3 2.29482
R251 VTAIL.n0 VTAIL.t11 2.29482
R252 VTAIL.n48 VTAIL.t7 2.29482
R253 VTAIL.n48 VTAIL.t10 2.29482
R254 VTAIL.n98 VTAIL.t5 2.29482
R255 VTAIL.n98 VTAIL.t9 2.29482
R256 VTAIL.n50 VTAIL.t4 2.29482
R257 VTAIL.n50 VTAIL.t1 2.29482
R258 VTAIL.n178 VTAIL.n152 1.93989
R259 VTAIL.n190 VTAIL.n146 1.93989
R260 VTAIL.n34 VTAIL.n8 1.93989
R261 VTAIL.n46 VTAIL.n2 1.93989
R262 VTAIL.n144 VTAIL.n100 1.93989
R263 VTAIL.n132 VTAIL.n106 1.93989
R264 VTAIL.n96 VTAIL.n52 1.93989
R265 VTAIL.n84 VTAIL.n58 1.93989
R266 VTAIL.n179 VTAIL.n150 1.16414
R267 VTAIL.n188 VTAIL.n187 1.16414
R268 VTAIL.n35 VTAIL.n6 1.16414
R269 VTAIL.n44 VTAIL.n43 1.16414
R270 VTAIL.n142 VTAIL.n141 1.16414
R271 VTAIL.n133 VTAIL.n104 1.16414
R272 VTAIL.n94 VTAIL.n93 1.16414
R273 VTAIL.n85 VTAIL.n56 1.16414
R274 VTAIL.n99 VTAIL.n97 0.931535
R275 VTAIL.n47 VTAIL.n1 0.931535
R276 VTAIL.n97 VTAIL.n51 0.922914
R277 VTAIL.n145 VTAIL.n99 0.922914
R278 VTAIL.n49 VTAIL.n47 0.922914
R279 VTAIL VTAIL.n191 0.634121
R280 VTAIL.n183 VTAIL.n182 0.388379
R281 VTAIL.n184 VTAIL.n148 0.388379
R282 VTAIL.n39 VTAIL.n38 0.388379
R283 VTAIL.n40 VTAIL.n4 0.388379
R284 VTAIL.n138 VTAIL.n102 0.388379
R285 VTAIL.n137 VTAIL.n136 0.388379
R286 VTAIL.n90 VTAIL.n54 0.388379
R287 VTAIL.n89 VTAIL.n88 0.388379
R288 VTAIL VTAIL.n1 0.289293
R289 VTAIL.n164 VTAIL.n163 0.155672
R290 VTAIL.n164 VTAIL.n155 0.155672
R291 VTAIL.n171 VTAIL.n155 0.155672
R292 VTAIL.n172 VTAIL.n171 0.155672
R293 VTAIL.n172 VTAIL.n151 0.155672
R294 VTAIL.n180 VTAIL.n151 0.155672
R295 VTAIL.n181 VTAIL.n180 0.155672
R296 VTAIL.n181 VTAIL.n147 0.155672
R297 VTAIL.n189 VTAIL.n147 0.155672
R298 VTAIL.n20 VTAIL.n19 0.155672
R299 VTAIL.n20 VTAIL.n11 0.155672
R300 VTAIL.n27 VTAIL.n11 0.155672
R301 VTAIL.n28 VTAIL.n27 0.155672
R302 VTAIL.n28 VTAIL.n7 0.155672
R303 VTAIL.n36 VTAIL.n7 0.155672
R304 VTAIL.n37 VTAIL.n36 0.155672
R305 VTAIL.n37 VTAIL.n3 0.155672
R306 VTAIL.n45 VTAIL.n3 0.155672
R307 VTAIL.n143 VTAIL.n101 0.155672
R308 VTAIL.n135 VTAIL.n101 0.155672
R309 VTAIL.n135 VTAIL.n134 0.155672
R310 VTAIL.n134 VTAIL.n105 0.155672
R311 VTAIL.n127 VTAIL.n105 0.155672
R312 VTAIL.n127 VTAIL.n126 0.155672
R313 VTAIL.n126 VTAIL.n110 0.155672
R314 VTAIL.n119 VTAIL.n110 0.155672
R315 VTAIL.n119 VTAIL.n118 0.155672
R316 VTAIL.n95 VTAIL.n53 0.155672
R317 VTAIL.n87 VTAIL.n53 0.155672
R318 VTAIL.n87 VTAIL.n86 0.155672
R319 VTAIL.n86 VTAIL.n57 0.155672
R320 VTAIL.n79 VTAIL.n57 0.155672
R321 VTAIL.n79 VTAIL.n78 0.155672
R322 VTAIL.n78 VTAIL.n62 0.155672
R323 VTAIL.n71 VTAIL.n62 0.155672
R324 VTAIL.n71 VTAIL.n70 0.155672
R325 VDD1.n40 VDD1.n0 289.615
R326 VDD1.n85 VDD1.n45 289.615
R327 VDD1.n41 VDD1.n40 185
R328 VDD1.n39 VDD1.n38 185
R329 VDD1.n37 VDD1.n3 185
R330 VDD1.n7 VDD1.n4 185
R331 VDD1.n32 VDD1.n31 185
R332 VDD1.n30 VDD1.n29 185
R333 VDD1.n9 VDD1.n8 185
R334 VDD1.n24 VDD1.n23 185
R335 VDD1.n22 VDD1.n21 185
R336 VDD1.n13 VDD1.n12 185
R337 VDD1.n16 VDD1.n15 185
R338 VDD1.n60 VDD1.n59 185
R339 VDD1.n57 VDD1.n56 185
R340 VDD1.n66 VDD1.n65 185
R341 VDD1.n68 VDD1.n67 185
R342 VDD1.n53 VDD1.n52 185
R343 VDD1.n74 VDD1.n73 185
R344 VDD1.n77 VDD1.n76 185
R345 VDD1.n75 VDD1.n49 185
R346 VDD1.n82 VDD1.n48 185
R347 VDD1.n84 VDD1.n83 185
R348 VDD1.n86 VDD1.n85 185
R349 VDD1.t2 VDD1.n14 149.524
R350 VDD1.t5 VDD1.n58 149.524
R351 VDD1.n40 VDD1.n39 104.615
R352 VDD1.n39 VDD1.n3 104.615
R353 VDD1.n7 VDD1.n3 104.615
R354 VDD1.n31 VDD1.n7 104.615
R355 VDD1.n31 VDD1.n30 104.615
R356 VDD1.n30 VDD1.n8 104.615
R357 VDD1.n23 VDD1.n8 104.615
R358 VDD1.n23 VDD1.n22 104.615
R359 VDD1.n22 VDD1.n12 104.615
R360 VDD1.n15 VDD1.n12 104.615
R361 VDD1.n59 VDD1.n56 104.615
R362 VDD1.n66 VDD1.n56 104.615
R363 VDD1.n67 VDD1.n66 104.615
R364 VDD1.n67 VDD1.n52 104.615
R365 VDD1.n74 VDD1.n52 104.615
R366 VDD1.n76 VDD1.n74 104.615
R367 VDD1.n76 VDD1.n75 104.615
R368 VDD1.n75 VDD1.n48 104.615
R369 VDD1.n84 VDD1.n48 104.615
R370 VDD1.n85 VDD1.n84 104.615
R371 VDD1.n91 VDD1.n90 65.7496
R372 VDD1.n93 VDD1.n92 65.5743
R373 VDD1.n15 VDD1.t2 52.3082
R374 VDD1.n59 VDD1.t5 52.3082
R375 VDD1 VDD1.n44 51.7475
R376 VDD1.n91 VDD1.n89 51.6339
R377 VDD1.n93 VDD1.n91 35.197
R378 VDD1.n38 VDD1.n37 13.1884
R379 VDD1.n83 VDD1.n82 13.1884
R380 VDD1.n41 VDD1.n2 12.8005
R381 VDD1.n36 VDD1.n4 12.8005
R382 VDD1.n81 VDD1.n49 12.8005
R383 VDD1.n86 VDD1.n47 12.8005
R384 VDD1.n42 VDD1.n0 12.0247
R385 VDD1.n33 VDD1.n32 12.0247
R386 VDD1.n78 VDD1.n77 12.0247
R387 VDD1.n87 VDD1.n45 12.0247
R388 VDD1.n29 VDD1.n6 11.249
R389 VDD1.n73 VDD1.n51 11.249
R390 VDD1.n28 VDD1.n9 10.4732
R391 VDD1.n72 VDD1.n53 10.4732
R392 VDD1.n16 VDD1.n14 10.2747
R393 VDD1.n60 VDD1.n58 10.2747
R394 VDD1.n25 VDD1.n24 9.69747
R395 VDD1.n69 VDD1.n68 9.69747
R396 VDD1.n44 VDD1.n43 9.45567
R397 VDD1.n89 VDD1.n88 9.45567
R398 VDD1.n18 VDD1.n17 9.3005
R399 VDD1.n20 VDD1.n19 9.3005
R400 VDD1.n11 VDD1.n10 9.3005
R401 VDD1.n26 VDD1.n25 9.3005
R402 VDD1.n28 VDD1.n27 9.3005
R403 VDD1.n6 VDD1.n5 9.3005
R404 VDD1.n34 VDD1.n33 9.3005
R405 VDD1.n36 VDD1.n35 9.3005
R406 VDD1.n43 VDD1.n42 9.3005
R407 VDD1.n2 VDD1.n1 9.3005
R408 VDD1.n88 VDD1.n87 9.3005
R409 VDD1.n47 VDD1.n46 9.3005
R410 VDD1.n62 VDD1.n61 9.3005
R411 VDD1.n64 VDD1.n63 9.3005
R412 VDD1.n55 VDD1.n54 9.3005
R413 VDD1.n70 VDD1.n69 9.3005
R414 VDD1.n72 VDD1.n71 9.3005
R415 VDD1.n51 VDD1.n50 9.3005
R416 VDD1.n79 VDD1.n78 9.3005
R417 VDD1.n81 VDD1.n80 9.3005
R418 VDD1.n21 VDD1.n11 8.92171
R419 VDD1.n65 VDD1.n55 8.92171
R420 VDD1.n20 VDD1.n13 8.14595
R421 VDD1.n64 VDD1.n57 8.14595
R422 VDD1.n17 VDD1.n16 7.3702
R423 VDD1.n61 VDD1.n60 7.3702
R424 VDD1.n17 VDD1.n13 5.81868
R425 VDD1.n61 VDD1.n57 5.81868
R426 VDD1.n21 VDD1.n20 5.04292
R427 VDD1.n65 VDD1.n64 5.04292
R428 VDD1.n24 VDD1.n11 4.26717
R429 VDD1.n68 VDD1.n55 4.26717
R430 VDD1.n25 VDD1.n9 3.49141
R431 VDD1.n69 VDD1.n53 3.49141
R432 VDD1.n62 VDD1.n58 2.84303
R433 VDD1.n18 VDD1.n14 2.84303
R434 VDD1.n29 VDD1.n28 2.71565
R435 VDD1.n73 VDD1.n72 2.71565
R436 VDD1.n92 VDD1.t1 2.29482
R437 VDD1.n92 VDD1.t3 2.29482
R438 VDD1.n90 VDD1.t0 2.29482
R439 VDD1.n90 VDD1.t4 2.29482
R440 VDD1.n44 VDD1.n0 1.93989
R441 VDD1.n32 VDD1.n6 1.93989
R442 VDD1.n77 VDD1.n51 1.93989
R443 VDD1.n89 VDD1.n45 1.93989
R444 VDD1.n42 VDD1.n41 1.16414
R445 VDD1.n33 VDD1.n4 1.16414
R446 VDD1.n78 VDD1.n49 1.16414
R447 VDD1.n87 VDD1.n86 1.16414
R448 VDD1.n38 VDD1.n2 0.388379
R449 VDD1.n37 VDD1.n36 0.388379
R450 VDD1.n82 VDD1.n81 0.388379
R451 VDD1.n83 VDD1.n47 0.388379
R452 VDD1 VDD1.n93 0.172914
R453 VDD1.n43 VDD1.n1 0.155672
R454 VDD1.n35 VDD1.n1 0.155672
R455 VDD1.n35 VDD1.n34 0.155672
R456 VDD1.n34 VDD1.n5 0.155672
R457 VDD1.n27 VDD1.n5 0.155672
R458 VDD1.n27 VDD1.n26 0.155672
R459 VDD1.n26 VDD1.n10 0.155672
R460 VDD1.n19 VDD1.n10 0.155672
R461 VDD1.n19 VDD1.n18 0.155672
R462 VDD1.n63 VDD1.n62 0.155672
R463 VDD1.n63 VDD1.n54 0.155672
R464 VDD1.n70 VDD1.n54 0.155672
R465 VDD1.n71 VDD1.n70 0.155672
R466 VDD1.n71 VDD1.n50 0.155672
R467 VDD1.n79 VDD1.n50 0.155672
R468 VDD1.n80 VDD1.n79 0.155672
R469 VDD1.n80 VDD1.n46 0.155672
R470 VDD1.n88 VDD1.n46 0.155672
R471 B.n541 B.n540 585
R472 B.n542 B.n541 585
R473 B.n225 B.n78 585
R474 B.n224 B.n223 585
R475 B.n222 B.n221 585
R476 B.n220 B.n219 585
R477 B.n218 B.n217 585
R478 B.n216 B.n215 585
R479 B.n214 B.n213 585
R480 B.n212 B.n211 585
R481 B.n210 B.n209 585
R482 B.n208 B.n207 585
R483 B.n206 B.n205 585
R484 B.n204 B.n203 585
R485 B.n202 B.n201 585
R486 B.n200 B.n199 585
R487 B.n198 B.n197 585
R488 B.n196 B.n195 585
R489 B.n194 B.n193 585
R490 B.n192 B.n191 585
R491 B.n190 B.n189 585
R492 B.n188 B.n187 585
R493 B.n186 B.n185 585
R494 B.n184 B.n183 585
R495 B.n182 B.n181 585
R496 B.n180 B.n179 585
R497 B.n178 B.n177 585
R498 B.n176 B.n175 585
R499 B.n174 B.n173 585
R500 B.n172 B.n171 585
R501 B.n170 B.n169 585
R502 B.n168 B.n167 585
R503 B.n166 B.n165 585
R504 B.n163 B.n162 585
R505 B.n161 B.n160 585
R506 B.n159 B.n158 585
R507 B.n157 B.n156 585
R508 B.n155 B.n154 585
R509 B.n153 B.n152 585
R510 B.n151 B.n150 585
R511 B.n149 B.n148 585
R512 B.n147 B.n146 585
R513 B.n145 B.n144 585
R514 B.n143 B.n142 585
R515 B.n141 B.n140 585
R516 B.n139 B.n138 585
R517 B.n137 B.n136 585
R518 B.n135 B.n134 585
R519 B.n133 B.n132 585
R520 B.n131 B.n130 585
R521 B.n129 B.n128 585
R522 B.n127 B.n126 585
R523 B.n125 B.n124 585
R524 B.n123 B.n122 585
R525 B.n121 B.n120 585
R526 B.n119 B.n118 585
R527 B.n117 B.n116 585
R528 B.n115 B.n114 585
R529 B.n113 B.n112 585
R530 B.n111 B.n110 585
R531 B.n109 B.n108 585
R532 B.n107 B.n106 585
R533 B.n105 B.n104 585
R534 B.n103 B.n102 585
R535 B.n101 B.n100 585
R536 B.n99 B.n98 585
R537 B.n97 B.n96 585
R538 B.n95 B.n94 585
R539 B.n93 B.n92 585
R540 B.n91 B.n90 585
R541 B.n89 B.n88 585
R542 B.n87 B.n86 585
R543 B.n85 B.n84 585
R544 B.n40 B.n39 585
R545 B.n539 B.n41 585
R546 B.n543 B.n41 585
R547 B.n538 B.n537 585
R548 B.n537 B.n37 585
R549 B.n536 B.n36 585
R550 B.n549 B.n36 585
R551 B.n535 B.n35 585
R552 B.n550 B.n35 585
R553 B.n534 B.n34 585
R554 B.n551 B.n34 585
R555 B.n533 B.n532 585
R556 B.n532 B.n30 585
R557 B.n531 B.n29 585
R558 B.n557 B.n29 585
R559 B.n530 B.n28 585
R560 B.n558 B.n28 585
R561 B.n529 B.n27 585
R562 B.n559 B.n27 585
R563 B.n528 B.n527 585
R564 B.n527 B.n23 585
R565 B.n526 B.n22 585
R566 B.n565 B.n22 585
R567 B.n525 B.n21 585
R568 B.n566 B.n21 585
R569 B.n524 B.n20 585
R570 B.n567 B.n20 585
R571 B.n523 B.n522 585
R572 B.n522 B.n16 585
R573 B.n521 B.n15 585
R574 B.n573 B.n15 585
R575 B.n520 B.n14 585
R576 B.n574 B.n14 585
R577 B.n519 B.n13 585
R578 B.n575 B.n13 585
R579 B.n518 B.n517 585
R580 B.n517 B.n12 585
R581 B.n516 B.n515 585
R582 B.n516 B.n8 585
R583 B.n514 B.n7 585
R584 B.n582 B.n7 585
R585 B.n513 B.n6 585
R586 B.n583 B.n6 585
R587 B.n512 B.n5 585
R588 B.n584 B.n5 585
R589 B.n511 B.n510 585
R590 B.n510 B.n4 585
R591 B.n509 B.n226 585
R592 B.n509 B.n508 585
R593 B.n498 B.n227 585
R594 B.n501 B.n227 585
R595 B.n500 B.n499 585
R596 B.n502 B.n500 585
R597 B.n497 B.n232 585
R598 B.n232 B.n231 585
R599 B.n496 B.n495 585
R600 B.n495 B.n494 585
R601 B.n234 B.n233 585
R602 B.n235 B.n234 585
R603 B.n487 B.n486 585
R604 B.n488 B.n487 585
R605 B.n485 B.n239 585
R606 B.n243 B.n239 585
R607 B.n484 B.n483 585
R608 B.n483 B.n482 585
R609 B.n241 B.n240 585
R610 B.n242 B.n241 585
R611 B.n475 B.n474 585
R612 B.n476 B.n475 585
R613 B.n473 B.n248 585
R614 B.n248 B.n247 585
R615 B.n472 B.n471 585
R616 B.n471 B.n470 585
R617 B.n250 B.n249 585
R618 B.n251 B.n250 585
R619 B.n463 B.n462 585
R620 B.n464 B.n463 585
R621 B.n461 B.n256 585
R622 B.n256 B.n255 585
R623 B.n460 B.n459 585
R624 B.n459 B.n458 585
R625 B.n258 B.n257 585
R626 B.n259 B.n258 585
R627 B.n451 B.n450 585
R628 B.n452 B.n451 585
R629 B.n262 B.n261 585
R630 B.n306 B.n304 585
R631 B.n307 B.n303 585
R632 B.n307 B.n263 585
R633 B.n310 B.n309 585
R634 B.n311 B.n302 585
R635 B.n313 B.n312 585
R636 B.n315 B.n301 585
R637 B.n318 B.n317 585
R638 B.n319 B.n300 585
R639 B.n321 B.n320 585
R640 B.n323 B.n299 585
R641 B.n326 B.n325 585
R642 B.n327 B.n298 585
R643 B.n329 B.n328 585
R644 B.n331 B.n297 585
R645 B.n334 B.n333 585
R646 B.n335 B.n296 585
R647 B.n337 B.n336 585
R648 B.n339 B.n295 585
R649 B.n342 B.n341 585
R650 B.n343 B.n294 585
R651 B.n345 B.n344 585
R652 B.n347 B.n293 585
R653 B.n350 B.n349 585
R654 B.n351 B.n292 585
R655 B.n353 B.n352 585
R656 B.n355 B.n291 585
R657 B.n358 B.n357 585
R658 B.n359 B.n290 585
R659 B.n361 B.n360 585
R660 B.n363 B.n289 585
R661 B.n366 B.n365 585
R662 B.n368 B.n286 585
R663 B.n370 B.n369 585
R664 B.n372 B.n285 585
R665 B.n375 B.n374 585
R666 B.n376 B.n284 585
R667 B.n378 B.n377 585
R668 B.n380 B.n283 585
R669 B.n383 B.n382 585
R670 B.n384 B.n280 585
R671 B.n387 B.n386 585
R672 B.n389 B.n279 585
R673 B.n392 B.n391 585
R674 B.n393 B.n278 585
R675 B.n395 B.n394 585
R676 B.n397 B.n277 585
R677 B.n400 B.n399 585
R678 B.n401 B.n276 585
R679 B.n403 B.n402 585
R680 B.n405 B.n275 585
R681 B.n408 B.n407 585
R682 B.n409 B.n274 585
R683 B.n411 B.n410 585
R684 B.n413 B.n273 585
R685 B.n416 B.n415 585
R686 B.n417 B.n272 585
R687 B.n419 B.n418 585
R688 B.n421 B.n271 585
R689 B.n424 B.n423 585
R690 B.n425 B.n270 585
R691 B.n427 B.n426 585
R692 B.n429 B.n269 585
R693 B.n432 B.n431 585
R694 B.n433 B.n268 585
R695 B.n435 B.n434 585
R696 B.n437 B.n267 585
R697 B.n440 B.n439 585
R698 B.n441 B.n266 585
R699 B.n443 B.n442 585
R700 B.n445 B.n265 585
R701 B.n448 B.n447 585
R702 B.n449 B.n264 585
R703 B.n454 B.n453 585
R704 B.n453 B.n452 585
R705 B.n455 B.n260 585
R706 B.n260 B.n259 585
R707 B.n457 B.n456 585
R708 B.n458 B.n457 585
R709 B.n254 B.n253 585
R710 B.n255 B.n254 585
R711 B.n466 B.n465 585
R712 B.n465 B.n464 585
R713 B.n467 B.n252 585
R714 B.n252 B.n251 585
R715 B.n469 B.n468 585
R716 B.n470 B.n469 585
R717 B.n246 B.n245 585
R718 B.n247 B.n246 585
R719 B.n478 B.n477 585
R720 B.n477 B.n476 585
R721 B.n479 B.n244 585
R722 B.n244 B.n242 585
R723 B.n481 B.n480 585
R724 B.n482 B.n481 585
R725 B.n238 B.n237 585
R726 B.n243 B.n238 585
R727 B.n490 B.n489 585
R728 B.n489 B.n488 585
R729 B.n491 B.n236 585
R730 B.n236 B.n235 585
R731 B.n493 B.n492 585
R732 B.n494 B.n493 585
R733 B.n230 B.n229 585
R734 B.n231 B.n230 585
R735 B.n504 B.n503 585
R736 B.n503 B.n502 585
R737 B.n505 B.n228 585
R738 B.n501 B.n228 585
R739 B.n507 B.n506 585
R740 B.n508 B.n507 585
R741 B.n3 B.n0 585
R742 B.n4 B.n3 585
R743 B.n581 B.n1 585
R744 B.n582 B.n581 585
R745 B.n580 B.n579 585
R746 B.n580 B.n8 585
R747 B.n578 B.n9 585
R748 B.n12 B.n9 585
R749 B.n577 B.n576 585
R750 B.n576 B.n575 585
R751 B.n11 B.n10 585
R752 B.n574 B.n11 585
R753 B.n572 B.n571 585
R754 B.n573 B.n572 585
R755 B.n570 B.n17 585
R756 B.n17 B.n16 585
R757 B.n569 B.n568 585
R758 B.n568 B.n567 585
R759 B.n19 B.n18 585
R760 B.n566 B.n19 585
R761 B.n564 B.n563 585
R762 B.n565 B.n564 585
R763 B.n562 B.n24 585
R764 B.n24 B.n23 585
R765 B.n561 B.n560 585
R766 B.n560 B.n559 585
R767 B.n26 B.n25 585
R768 B.n558 B.n26 585
R769 B.n556 B.n555 585
R770 B.n557 B.n556 585
R771 B.n554 B.n31 585
R772 B.n31 B.n30 585
R773 B.n553 B.n552 585
R774 B.n552 B.n551 585
R775 B.n33 B.n32 585
R776 B.n550 B.n33 585
R777 B.n548 B.n547 585
R778 B.n549 B.n548 585
R779 B.n546 B.n38 585
R780 B.n38 B.n37 585
R781 B.n545 B.n544 585
R782 B.n544 B.n543 585
R783 B.n585 B.n584 585
R784 B.n583 B.n2 585
R785 B.n544 B.n40 530.939
R786 B.n541 B.n41 530.939
R787 B.n451 B.n264 530.939
R788 B.n453 B.n262 530.939
R789 B.n81 B.t6 483.558
R790 B.n79 B.t14 483.558
R791 B.n281 B.t10 483.558
R792 B.n287 B.t17 483.558
R793 B.n542 B.n77 256.663
R794 B.n542 B.n76 256.663
R795 B.n542 B.n75 256.663
R796 B.n542 B.n74 256.663
R797 B.n542 B.n73 256.663
R798 B.n542 B.n72 256.663
R799 B.n542 B.n71 256.663
R800 B.n542 B.n70 256.663
R801 B.n542 B.n69 256.663
R802 B.n542 B.n68 256.663
R803 B.n542 B.n67 256.663
R804 B.n542 B.n66 256.663
R805 B.n542 B.n65 256.663
R806 B.n542 B.n64 256.663
R807 B.n542 B.n63 256.663
R808 B.n542 B.n62 256.663
R809 B.n542 B.n61 256.663
R810 B.n542 B.n60 256.663
R811 B.n542 B.n59 256.663
R812 B.n542 B.n58 256.663
R813 B.n542 B.n57 256.663
R814 B.n542 B.n56 256.663
R815 B.n542 B.n55 256.663
R816 B.n542 B.n54 256.663
R817 B.n542 B.n53 256.663
R818 B.n542 B.n52 256.663
R819 B.n542 B.n51 256.663
R820 B.n542 B.n50 256.663
R821 B.n542 B.n49 256.663
R822 B.n542 B.n48 256.663
R823 B.n542 B.n47 256.663
R824 B.n542 B.n46 256.663
R825 B.n542 B.n45 256.663
R826 B.n542 B.n44 256.663
R827 B.n542 B.n43 256.663
R828 B.n542 B.n42 256.663
R829 B.n305 B.n263 256.663
R830 B.n308 B.n263 256.663
R831 B.n314 B.n263 256.663
R832 B.n316 B.n263 256.663
R833 B.n322 B.n263 256.663
R834 B.n324 B.n263 256.663
R835 B.n330 B.n263 256.663
R836 B.n332 B.n263 256.663
R837 B.n338 B.n263 256.663
R838 B.n340 B.n263 256.663
R839 B.n346 B.n263 256.663
R840 B.n348 B.n263 256.663
R841 B.n354 B.n263 256.663
R842 B.n356 B.n263 256.663
R843 B.n362 B.n263 256.663
R844 B.n364 B.n263 256.663
R845 B.n371 B.n263 256.663
R846 B.n373 B.n263 256.663
R847 B.n379 B.n263 256.663
R848 B.n381 B.n263 256.663
R849 B.n388 B.n263 256.663
R850 B.n390 B.n263 256.663
R851 B.n396 B.n263 256.663
R852 B.n398 B.n263 256.663
R853 B.n404 B.n263 256.663
R854 B.n406 B.n263 256.663
R855 B.n412 B.n263 256.663
R856 B.n414 B.n263 256.663
R857 B.n420 B.n263 256.663
R858 B.n422 B.n263 256.663
R859 B.n428 B.n263 256.663
R860 B.n430 B.n263 256.663
R861 B.n436 B.n263 256.663
R862 B.n438 B.n263 256.663
R863 B.n444 B.n263 256.663
R864 B.n446 B.n263 256.663
R865 B.n587 B.n586 256.663
R866 B.n79 B.t15 244.782
R867 B.n281 B.t13 244.782
R868 B.n81 B.t8 244.782
R869 B.n287 B.t19 244.782
R870 B.n80 B.t16 224.03
R871 B.n282 B.t12 224.03
R872 B.n82 B.t9 224.03
R873 B.n288 B.t18 224.03
R874 B.n86 B.n85 163.367
R875 B.n90 B.n89 163.367
R876 B.n94 B.n93 163.367
R877 B.n98 B.n97 163.367
R878 B.n102 B.n101 163.367
R879 B.n106 B.n105 163.367
R880 B.n110 B.n109 163.367
R881 B.n114 B.n113 163.367
R882 B.n118 B.n117 163.367
R883 B.n122 B.n121 163.367
R884 B.n126 B.n125 163.367
R885 B.n130 B.n129 163.367
R886 B.n134 B.n133 163.367
R887 B.n138 B.n137 163.367
R888 B.n142 B.n141 163.367
R889 B.n146 B.n145 163.367
R890 B.n150 B.n149 163.367
R891 B.n154 B.n153 163.367
R892 B.n158 B.n157 163.367
R893 B.n162 B.n161 163.367
R894 B.n167 B.n166 163.367
R895 B.n171 B.n170 163.367
R896 B.n175 B.n174 163.367
R897 B.n179 B.n178 163.367
R898 B.n183 B.n182 163.367
R899 B.n187 B.n186 163.367
R900 B.n191 B.n190 163.367
R901 B.n195 B.n194 163.367
R902 B.n199 B.n198 163.367
R903 B.n203 B.n202 163.367
R904 B.n207 B.n206 163.367
R905 B.n211 B.n210 163.367
R906 B.n215 B.n214 163.367
R907 B.n219 B.n218 163.367
R908 B.n223 B.n222 163.367
R909 B.n541 B.n78 163.367
R910 B.n451 B.n258 163.367
R911 B.n459 B.n258 163.367
R912 B.n459 B.n256 163.367
R913 B.n463 B.n256 163.367
R914 B.n463 B.n250 163.367
R915 B.n471 B.n250 163.367
R916 B.n471 B.n248 163.367
R917 B.n475 B.n248 163.367
R918 B.n475 B.n241 163.367
R919 B.n483 B.n241 163.367
R920 B.n483 B.n239 163.367
R921 B.n487 B.n239 163.367
R922 B.n487 B.n234 163.367
R923 B.n495 B.n234 163.367
R924 B.n495 B.n232 163.367
R925 B.n500 B.n232 163.367
R926 B.n500 B.n227 163.367
R927 B.n509 B.n227 163.367
R928 B.n510 B.n509 163.367
R929 B.n510 B.n5 163.367
R930 B.n6 B.n5 163.367
R931 B.n7 B.n6 163.367
R932 B.n516 B.n7 163.367
R933 B.n517 B.n516 163.367
R934 B.n517 B.n13 163.367
R935 B.n14 B.n13 163.367
R936 B.n15 B.n14 163.367
R937 B.n522 B.n15 163.367
R938 B.n522 B.n20 163.367
R939 B.n21 B.n20 163.367
R940 B.n22 B.n21 163.367
R941 B.n527 B.n22 163.367
R942 B.n527 B.n27 163.367
R943 B.n28 B.n27 163.367
R944 B.n29 B.n28 163.367
R945 B.n532 B.n29 163.367
R946 B.n532 B.n34 163.367
R947 B.n35 B.n34 163.367
R948 B.n36 B.n35 163.367
R949 B.n537 B.n36 163.367
R950 B.n537 B.n41 163.367
R951 B.n307 B.n306 163.367
R952 B.n309 B.n307 163.367
R953 B.n313 B.n302 163.367
R954 B.n317 B.n315 163.367
R955 B.n321 B.n300 163.367
R956 B.n325 B.n323 163.367
R957 B.n329 B.n298 163.367
R958 B.n333 B.n331 163.367
R959 B.n337 B.n296 163.367
R960 B.n341 B.n339 163.367
R961 B.n345 B.n294 163.367
R962 B.n349 B.n347 163.367
R963 B.n353 B.n292 163.367
R964 B.n357 B.n355 163.367
R965 B.n361 B.n290 163.367
R966 B.n365 B.n363 163.367
R967 B.n370 B.n286 163.367
R968 B.n374 B.n372 163.367
R969 B.n378 B.n284 163.367
R970 B.n382 B.n380 163.367
R971 B.n387 B.n280 163.367
R972 B.n391 B.n389 163.367
R973 B.n395 B.n278 163.367
R974 B.n399 B.n397 163.367
R975 B.n403 B.n276 163.367
R976 B.n407 B.n405 163.367
R977 B.n411 B.n274 163.367
R978 B.n415 B.n413 163.367
R979 B.n419 B.n272 163.367
R980 B.n423 B.n421 163.367
R981 B.n427 B.n270 163.367
R982 B.n431 B.n429 163.367
R983 B.n435 B.n268 163.367
R984 B.n439 B.n437 163.367
R985 B.n443 B.n266 163.367
R986 B.n447 B.n445 163.367
R987 B.n453 B.n260 163.367
R988 B.n457 B.n260 163.367
R989 B.n457 B.n254 163.367
R990 B.n465 B.n254 163.367
R991 B.n465 B.n252 163.367
R992 B.n469 B.n252 163.367
R993 B.n469 B.n246 163.367
R994 B.n477 B.n246 163.367
R995 B.n477 B.n244 163.367
R996 B.n481 B.n244 163.367
R997 B.n481 B.n238 163.367
R998 B.n489 B.n238 163.367
R999 B.n489 B.n236 163.367
R1000 B.n493 B.n236 163.367
R1001 B.n493 B.n230 163.367
R1002 B.n503 B.n230 163.367
R1003 B.n503 B.n228 163.367
R1004 B.n507 B.n228 163.367
R1005 B.n507 B.n3 163.367
R1006 B.n585 B.n3 163.367
R1007 B.n581 B.n2 163.367
R1008 B.n581 B.n580 163.367
R1009 B.n580 B.n9 163.367
R1010 B.n576 B.n9 163.367
R1011 B.n576 B.n11 163.367
R1012 B.n572 B.n11 163.367
R1013 B.n572 B.n17 163.367
R1014 B.n568 B.n17 163.367
R1015 B.n568 B.n19 163.367
R1016 B.n564 B.n19 163.367
R1017 B.n564 B.n24 163.367
R1018 B.n560 B.n24 163.367
R1019 B.n560 B.n26 163.367
R1020 B.n556 B.n26 163.367
R1021 B.n556 B.n31 163.367
R1022 B.n552 B.n31 163.367
R1023 B.n552 B.n33 163.367
R1024 B.n548 B.n33 163.367
R1025 B.n548 B.n38 163.367
R1026 B.n544 B.n38 163.367
R1027 B.n452 B.n263 108.379
R1028 B.n543 B.n542 108.379
R1029 B.n42 B.n40 71.676
R1030 B.n86 B.n43 71.676
R1031 B.n90 B.n44 71.676
R1032 B.n94 B.n45 71.676
R1033 B.n98 B.n46 71.676
R1034 B.n102 B.n47 71.676
R1035 B.n106 B.n48 71.676
R1036 B.n110 B.n49 71.676
R1037 B.n114 B.n50 71.676
R1038 B.n118 B.n51 71.676
R1039 B.n122 B.n52 71.676
R1040 B.n126 B.n53 71.676
R1041 B.n130 B.n54 71.676
R1042 B.n134 B.n55 71.676
R1043 B.n138 B.n56 71.676
R1044 B.n142 B.n57 71.676
R1045 B.n146 B.n58 71.676
R1046 B.n150 B.n59 71.676
R1047 B.n154 B.n60 71.676
R1048 B.n158 B.n61 71.676
R1049 B.n162 B.n62 71.676
R1050 B.n167 B.n63 71.676
R1051 B.n171 B.n64 71.676
R1052 B.n175 B.n65 71.676
R1053 B.n179 B.n66 71.676
R1054 B.n183 B.n67 71.676
R1055 B.n187 B.n68 71.676
R1056 B.n191 B.n69 71.676
R1057 B.n195 B.n70 71.676
R1058 B.n199 B.n71 71.676
R1059 B.n203 B.n72 71.676
R1060 B.n207 B.n73 71.676
R1061 B.n211 B.n74 71.676
R1062 B.n215 B.n75 71.676
R1063 B.n219 B.n76 71.676
R1064 B.n223 B.n77 71.676
R1065 B.n78 B.n77 71.676
R1066 B.n222 B.n76 71.676
R1067 B.n218 B.n75 71.676
R1068 B.n214 B.n74 71.676
R1069 B.n210 B.n73 71.676
R1070 B.n206 B.n72 71.676
R1071 B.n202 B.n71 71.676
R1072 B.n198 B.n70 71.676
R1073 B.n194 B.n69 71.676
R1074 B.n190 B.n68 71.676
R1075 B.n186 B.n67 71.676
R1076 B.n182 B.n66 71.676
R1077 B.n178 B.n65 71.676
R1078 B.n174 B.n64 71.676
R1079 B.n170 B.n63 71.676
R1080 B.n166 B.n62 71.676
R1081 B.n161 B.n61 71.676
R1082 B.n157 B.n60 71.676
R1083 B.n153 B.n59 71.676
R1084 B.n149 B.n58 71.676
R1085 B.n145 B.n57 71.676
R1086 B.n141 B.n56 71.676
R1087 B.n137 B.n55 71.676
R1088 B.n133 B.n54 71.676
R1089 B.n129 B.n53 71.676
R1090 B.n125 B.n52 71.676
R1091 B.n121 B.n51 71.676
R1092 B.n117 B.n50 71.676
R1093 B.n113 B.n49 71.676
R1094 B.n109 B.n48 71.676
R1095 B.n105 B.n47 71.676
R1096 B.n101 B.n46 71.676
R1097 B.n97 B.n45 71.676
R1098 B.n93 B.n44 71.676
R1099 B.n89 B.n43 71.676
R1100 B.n85 B.n42 71.676
R1101 B.n305 B.n262 71.676
R1102 B.n309 B.n308 71.676
R1103 B.n314 B.n313 71.676
R1104 B.n317 B.n316 71.676
R1105 B.n322 B.n321 71.676
R1106 B.n325 B.n324 71.676
R1107 B.n330 B.n329 71.676
R1108 B.n333 B.n332 71.676
R1109 B.n338 B.n337 71.676
R1110 B.n341 B.n340 71.676
R1111 B.n346 B.n345 71.676
R1112 B.n349 B.n348 71.676
R1113 B.n354 B.n353 71.676
R1114 B.n357 B.n356 71.676
R1115 B.n362 B.n361 71.676
R1116 B.n365 B.n364 71.676
R1117 B.n371 B.n370 71.676
R1118 B.n374 B.n373 71.676
R1119 B.n379 B.n378 71.676
R1120 B.n382 B.n381 71.676
R1121 B.n388 B.n387 71.676
R1122 B.n391 B.n390 71.676
R1123 B.n396 B.n395 71.676
R1124 B.n399 B.n398 71.676
R1125 B.n404 B.n403 71.676
R1126 B.n407 B.n406 71.676
R1127 B.n412 B.n411 71.676
R1128 B.n415 B.n414 71.676
R1129 B.n420 B.n419 71.676
R1130 B.n423 B.n422 71.676
R1131 B.n428 B.n427 71.676
R1132 B.n431 B.n430 71.676
R1133 B.n436 B.n435 71.676
R1134 B.n439 B.n438 71.676
R1135 B.n444 B.n443 71.676
R1136 B.n447 B.n446 71.676
R1137 B.n306 B.n305 71.676
R1138 B.n308 B.n302 71.676
R1139 B.n315 B.n314 71.676
R1140 B.n316 B.n300 71.676
R1141 B.n323 B.n322 71.676
R1142 B.n324 B.n298 71.676
R1143 B.n331 B.n330 71.676
R1144 B.n332 B.n296 71.676
R1145 B.n339 B.n338 71.676
R1146 B.n340 B.n294 71.676
R1147 B.n347 B.n346 71.676
R1148 B.n348 B.n292 71.676
R1149 B.n355 B.n354 71.676
R1150 B.n356 B.n290 71.676
R1151 B.n363 B.n362 71.676
R1152 B.n364 B.n286 71.676
R1153 B.n372 B.n371 71.676
R1154 B.n373 B.n284 71.676
R1155 B.n380 B.n379 71.676
R1156 B.n381 B.n280 71.676
R1157 B.n389 B.n388 71.676
R1158 B.n390 B.n278 71.676
R1159 B.n397 B.n396 71.676
R1160 B.n398 B.n276 71.676
R1161 B.n405 B.n404 71.676
R1162 B.n406 B.n274 71.676
R1163 B.n413 B.n412 71.676
R1164 B.n414 B.n272 71.676
R1165 B.n421 B.n420 71.676
R1166 B.n422 B.n270 71.676
R1167 B.n429 B.n428 71.676
R1168 B.n430 B.n268 71.676
R1169 B.n437 B.n436 71.676
R1170 B.n438 B.n266 71.676
R1171 B.n445 B.n444 71.676
R1172 B.n446 B.n264 71.676
R1173 B.n586 B.n585 71.676
R1174 B.n586 B.n2 71.676
R1175 B.n83 B.n82 59.5399
R1176 B.n164 B.n80 59.5399
R1177 B.n385 B.n282 59.5399
R1178 B.n367 B.n288 59.5399
R1179 B.n452 B.n259 53.7941
R1180 B.n458 B.n259 53.7941
R1181 B.n458 B.n255 53.7941
R1182 B.n464 B.n255 53.7941
R1183 B.n470 B.n251 53.7941
R1184 B.n470 B.n247 53.7941
R1185 B.n476 B.n247 53.7941
R1186 B.n476 B.n242 53.7941
R1187 B.n482 B.n242 53.7941
R1188 B.n482 B.n243 53.7941
R1189 B.n488 B.n235 53.7941
R1190 B.n494 B.n235 53.7941
R1191 B.n502 B.n231 53.7941
R1192 B.n502 B.n501 53.7941
R1193 B.n508 B.n4 53.7941
R1194 B.n584 B.n4 53.7941
R1195 B.n584 B.n583 53.7941
R1196 B.n583 B.n582 53.7941
R1197 B.n582 B.n8 53.7941
R1198 B.n575 B.n12 53.7941
R1199 B.n575 B.n574 53.7941
R1200 B.n573 B.n16 53.7941
R1201 B.n567 B.n16 53.7941
R1202 B.n566 B.n565 53.7941
R1203 B.n565 B.n23 53.7941
R1204 B.n559 B.n23 53.7941
R1205 B.n559 B.n558 53.7941
R1206 B.n558 B.n557 53.7941
R1207 B.n557 B.n30 53.7941
R1208 B.n551 B.n550 53.7941
R1209 B.n550 B.n549 53.7941
R1210 B.n549 B.n37 53.7941
R1211 B.n543 B.n37 53.7941
R1212 B.n488 B.t4 52.2119
R1213 B.n567 B.t2 52.2119
R1214 B.t1 B.n231 44.3011
R1215 B.n574 B.t5 44.3011
R1216 B.n464 B.t11 36.3903
R1217 B.n508 B.t0 36.3903
R1218 B.t3 B.n8 36.3903
R1219 B.n551 B.t7 36.3903
R1220 B.n454 B.n261 34.4981
R1221 B.n450 B.n449 34.4981
R1222 B.n540 B.n539 34.4981
R1223 B.n545 B.n39 34.4981
R1224 B.n82 B.n81 20.752
R1225 B.n80 B.n79 20.752
R1226 B.n282 B.n281 20.752
R1227 B.n288 B.n287 20.752
R1228 B B.n587 18.0485
R1229 B.t11 B.n251 17.4043
R1230 B.n501 B.t0 17.4043
R1231 B.n12 B.t3 17.4043
R1232 B.t7 B.n30 17.4043
R1233 B.n455 B.n454 10.6151
R1234 B.n456 B.n455 10.6151
R1235 B.n456 B.n253 10.6151
R1236 B.n466 B.n253 10.6151
R1237 B.n467 B.n466 10.6151
R1238 B.n468 B.n467 10.6151
R1239 B.n468 B.n245 10.6151
R1240 B.n478 B.n245 10.6151
R1241 B.n479 B.n478 10.6151
R1242 B.n480 B.n479 10.6151
R1243 B.n480 B.n237 10.6151
R1244 B.n490 B.n237 10.6151
R1245 B.n491 B.n490 10.6151
R1246 B.n492 B.n491 10.6151
R1247 B.n492 B.n229 10.6151
R1248 B.n504 B.n229 10.6151
R1249 B.n505 B.n504 10.6151
R1250 B.n506 B.n505 10.6151
R1251 B.n506 B.n0 10.6151
R1252 B.n304 B.n261 10.6151
R1253 B.n304 B.n303 10.6151
R1254 B.n310 B.n303 10.6151
R1255 B.n311 B.n310 10.6151
R1256 B.n312 B.n311 10.6151
R1257 B.n312 B.n301 10.6151
R1258 B.n318 B.n301 10.6151
R1259 B.n319 B.n318 10.6151
R1260 B.n320 B.n319 10.6151
R1261 B.n320 B.n299 10.6151
R1262 B.n326 B.n299 10.6151
R1263 B.n327 B.n326 10.6151
R1264 B.n328 B.n327 10.6151
R1265 B.n328 B.n297 10.6151
R1266 B.n334 B.n297 10.6151
R1267 B.n335 B.n334 10.6151
R1268 B.n336 B.n335 10.6151
R1269 B.n336 B.n295 10.6151
R1270 B.n342 B.n295 10.6151
R1271 B.n343 B.n342 10.6151
R1272 B.n344 B.n343 10.6151
R1273 B.n344 B.n293 10.6151
R1274 B.n350 B.n293 10.6151
R1275 B.n351 B.n350 10.6151
R1276 B.n352 B.n351 10.6151
R1277 B.n352 B.n291 10.6151
R1278 B.n358 B.n291 10.6151
R1279 B.n359 B.n358 10.6151
R1280 B.n360 B.n359 10.6151
R1281 B.n360 B.n289 10.6151
R1282 B.n366 B.n289 10.6151
R1283 B.n369 B.n368 10.6151
R1284 B.n369 B.n285 10.6151
R1285 B.n375 B.n285 10.6151
R1286 B.n376 B.n375 10.6151
R1287 B.n377 B.n376 10.6151
R1288 B.n377 B.n283 10.6151
R1289 B.n383 B.n283 10.6151
R1290 B.n384 B.n383 10.6151
R1291 B.n386 B.n279 10.6151
R1292 B.n392 B.n279 10.6151
R1293 B.n393 B.n392 10.6151
R1294 B.n394 B.n393 10.6151
R1295 B.n394 B.n277 10.6151
R1296 B.n400 B.n277 10.6151
R1297 B.n401 B.n400 10.6151
R1298 B.n402 B.n401 10.6151
R1299 B.n402 B.n275 10.6151
R1300 B.n408 B.n275 10.6151
R1301 B.n409 B.n408 10.6151
R1302 B.n410 B.n409 10.6151
R1303 B.n410 B.n273 10.6151
R1304 B.n416 B.n273 10.6151
R1305 B.n417 B.n416 10.6151
R1306 B.n418 B.n417 10.6151
R1307 B.n418 B.n271 10.6151
R1308 B.n424 B.n271 10.6151
R1309 B.n425 B.n424 10.6151
R1310 B.n426 B.n425 10.6151
R1311 B.n426 B.n269 10.6151
R1312 B.n432 B.n269 10.6151
R1313 B.n433 B.n432 10.6151
R1314 B.n434 B.n433 10.6151
R1315 B.n434 B.n267 10.6151
R1316 B.n440 B.n267 10.6151
R1317 B.n441 B.n440 10.6151
R1318 B.n442 B.n441 10.6151
R1319 B.n442 B.n265 10.6151
R1320 B.n448 B.n265 10.6151
R1321 B.n449 B.n448 10.6151
R1322 B.n450 B.n257 10.6151
R1323 B.n460 B.n257 10.6151
R1324 B.n461 B.n460 10.6151
R1325 B.n462 B.n461 10.6151
R1326 B.n462 B.n249 10.6151
R1327 B.n472 B.n249 10.6151
R1328 B.n473 B.n472 10.6151
R1329 B.n474 B.n473 10.6151
R1330 B.n474 B.n240 10.6151
R1331 B.n484 B.n240 10.6151
R1332 B.n485 B.n484 10.6151
R1333 B.n486 B.n485 10.6151
R1334 B.n486 B.n233 10.6151
R1335 B.n496 B.n233 10.6151
R1336 B.n497 B.n496 10.6151
R1337 B.n499 B.n497 10.6151
R1338 B.n499 B.n498 10.6151
R1339 B.n498 B.n226 10.6151
R1340 B.n511 B.n226 10.6151
R1341 B.n512 B.n511 10.6151
R1342 B.n513 B.n512 10.6151
R1343 B.n514 B.n513 10.6151
R1344 B.n515 B.n514 10.6151
R1345 B.n518 B.n515 10.6151
R1346 B.n519 B.n518 10.6151
R1347 B.n520 B.n519 10.6151
R1348 B.n521 B.n520 10.6151
R1349 B.n523 B.n521 10.6151
R1350 B.n524 B.n523 10.6151
R1351 B.n525 B.n524 10.6151
R1352 B.n526 B.n525 10.6151
R1353 B.n528 B.n526 10.6151
R1354 B.n529 B.n528 10.6151
R1355 B.n530 B.n529 10.6151
R1356 B.n531 B.n530 10.6151
R1357 B.n533 B.n531 10.6151
R1358 B.n534 B.n533 10.6151
R1359 B.n535 B.n534 10.6151
R1360 B.n536 B.n535 10.6151
R1361 B.n538 B.n536 10.6151
R1362 B.n539 B.n538 10.6151
R1363 B.n579 B.n1 10.6151
R1364 B.n579 B.n578 10.6151
R1365 B.n578 B.n577 10.6151
R1366 B.n577 B.n10 10.6151
R1367 B.n571 B.n10 10.6151
R1368 B.n571 B.n570 10.6151
R1369 B.n570 B.n569 10.6151
R1370 B.n569 B.n18 10.6151
R1371 B.n563 B.n18 10.6151
R1372 B.n563 B.n562 10.6151
R1373 B.n562 B.n561 10.6151
R1374 B.n561 B.n25 10.6151
R1375 B.n555 B.n25 10.6151
R1376 B.n555 B.n554 10.6151
R1377 B.n554 B.n553 10.6151
R1378 B.n553 B.n32 10.6151
R1379 B.n547 B.n32 10.6151
R1380 B.n547 B.n546 10.6151
R1381 B.n546 B.n545 10.6151
R1382 B.n84 B.n39 10.6151
R1383 B.n87 B.n84 10.6151
R1384 B.n88 B.n87 10.6151
R1385 B.n91 B.n88 10.6151
R1386 B.n92 B.n91 10.6151
R1387 B.n95 B.n92 10.6151
R1388 B.n96 B.n95 10.6151
R1389 B.n99 B.n96 10.6151
R1390 B.n100 B.n99 10.6151
R1391 B.n103 B.n100 10.6151
R1392 B.n104 B.n103 10.6151
R1393 B.n107 B.n104 10.6151
R1394 B.n108 B.n107 10.6151
R1395 B.n111 B.n108 10.6151
R1396 B.n112 B.n111 10.6151
R1397 B.n115 B.n112 10.6151
R1398 B.n116 B.n115 10.6151
R1399 B.n119 B.n116 10.6151
R1400 B.n120 B.n119 10.6151
R1401 B.n123 B.n120 10.6151
R1402 B.n124 B.n123 10.6151
R1403 B.n127 B.n124 10.6151
R1404 B.n128 B.n127 10.6151
R1405 B.n131 B.n128 10.6151
R1406 B.n132 B.n131 10.6151
R1407 B.n135 B.n132 10.6151
R1408 B.n136 B.n135 10.6151
R1409 B.n139 B.n136 10.6151
R1410 B.n140 B.n139 10.6151
R1411 B.n143 B.n140 10.6151
R1412 B.n144 B.n143 10.6151
R1413 B.n148 B.n147 10.6151
R1414 B.n151 B.n148 10.6151
R1415 B.n152 B.n151 10.6151
R1416 B.n155 B.n152 10.6151
R1417 B.n156 B.n155 10.6151
R1418 B.n159 B.n156 10.6151
R1419 B.n160 B.n159 10.6151
R1420 B.n163 B.n160 10.6151
R1421 B.n168 B.n165 10.6151
R1422 B.n169 B.n168 10.6151
R1423 B.n172 B.n169 10.6151
R1424 B.n173 B.n172 10.6151
R1425 B.n176 B.n173 10.6151
R1426 B.n177 B.n176 10.6151
R1427 B.n180 B.n177 10.6151
R1428 B.n181 B.n180 10.6151
R1429 B.n184 B.n181 10.6151
R1430 B.n185 B.n184 10.6151
R1431 B.n188 B.n185 10.6151
R1432 B.n189 B.n188 10.6151
R1433 B.n192 B.n189 10.6151
R1434 B.n193 B.n192 10.6151
R1435 B.n196 B.n193 10.6151
R1436 B.n197 B.n196 10.6151
R1437 B.n200 B.n197 10.6151
R1438 B.n201 B.n200 10.6151
R1439 B.n204 B.n201 10.6151
R1440 B.n205 B.n204 10.6151
R1441 B.n208 B.n205 10.6151
R1442 B.n209 B.n208 10.6151
R1443 B.n212 B.n209 10.6151
R1444 B.n213 B.n212 10.6151
R1445 B.n216 B.n213 10.6151
R1446 B.n217 B.n216 10.6151
R1447 B.n220 B.n217 10.6151
R1448 B.n221 B.n220 10.6151
R1449 B.n224 B.n221 10.6151
R1450 B.n225 B.n224 10.6151
R1451 B.n540 B.n225 10.6151
R1452 B.n494 B.t1 9.49349
R1453 B.t5 B.n573 9.49349
R1454 B.n587 B.n0 8.11757
R1455 B.n587 B.n1 8.11757
R1456 B.n368 B.n367 6.5566
R1457 B.n385 B.n384 6.5566
R1458 B.n147 B.n83 6.5566
R1459 B.n164 B.n163 6.5566
R1460 B.n367 B.n366 4.05904
R1461 B.n386 B.n385 4.05904
R1462 B.n144 B.n83 4.05904
R1463 B.n165 B.n164 4.05904
R1464 B.n243 B.t4 1.58266
R1465 B.t2 B.n566 1.58266
R1466 VN.n1 VN.t2 356.839
R1467 VN.n7 VN.t4 356.839
R1468 VN.n2 VN.t5 334.469
R1469 VN.n4 VN.t0 334.469
R1470 VN.n8 VN.t3 334.469
R1471 VN.n10 VN.t1 334.469
R1472 VN.n5 VN.n4 161.3
R1473 VN.n11 VN.n10 161.3
R1474 VN.n9 VN.n6 161.3
R1475 VN.n3 VN.n0 161.3
R1476 VN.n7 VN.n6 44.8655
R1477 VN.n1 VN.n0 44.8655
R1478 VN VN.n11 39.2259
R1479 VN.n4 VN.n3 29.2126
R1480 VN.n10 VN.n9 29.2126
R1481 VN.n2 VN.n1 19.4959
R1482 VN.n8 VN.n7 19.4959
R1483 VN.n3 VN.n2 18.9884
R1484 VN.n9 VN.n8 18.9884
R1485 VN.n11 VN.n6 0.189894
R1486 VN.n5 VN.n0 0.189894
R1487 VN VN.n5 0.0516364
R1488 VDD2.n87 VDD2.n47 289.615
R1489 VDD2.n40 VDD2.n0 289.615
R1490 VDD2.n88 VDD2.n87 185
R1491 VDD2.n86 VDD2.n85 185
R1492 VDD2.n84 VDD2.n50 185
R1493 VDD2.n54 VDD2.n51 185
R1494 VDD2.n79 VDD2.n78 185
R1495 VDD2.n77 VDD2.n76 185
R1496 VDD2.n56 VDD2.n55 185
R1497 VDD2.n71 VDD2.n70 185
R1498 VDD2.n69 VDD2.n68 185
R1499 VDD2.n60 VDD2.n59 185
R1500 VDD2.n63 VDD2.n62 185
R1501 VDD2.n15 VDD2.n14 185
R1502 VDD2.n12 VDD2.n11 185
R1503 VDD2.n21 VDD2.n20 185
R1504 VDD2.n23 VDD2.n22 185
R1505 VDD2.n8 VDD2.n7 185
R1506 VDD2.n29 VDD2.n28 185
R1507 VDD2.n32 VDD2.n31 185
R1508 VDD2.n30 VDD2.n4 185
R1509 VDD2.n37 VDD2.n3 185
R1510 VDD2.n39 VDD2.n38 185
R1511 VDD2.n41 VDD2.n40 185
R1512 VDD2.t4 VDD2.n61 149.524
R1513 VDD2.t3 VDD2.n13 149.524
R1514 VDD2.n87 VDD2.n86 104.615
R1515 VDD2.n86 VDD2.n50 104.615
R1516 VDD2.n54 VDD2.n50 104.615
R1517 VDD2.n78 VDD2.n54 104.615
R1518 VDD2.n78 VDD2.n77 104.615
R1519 VDD2.n77 VDD2.n55 104.615
R1520 VDD2.n70 VDD2.n55 104.615
R1521 VDD2.n70 VDD2.n69 104.615
R1522 VDD2.n69 VDD2.n59 104.615
R1523 VDD2.n62 VDD2.n59 104.615
R1524 VDD2.n14 VDD2.n11 104.615
R1525 VDD2.n21 VDD2.n11 104.615
R1526 VDD2.n22 VDD2.n21 104.615
R1527 VDD2.n22 VDD2.n7 104.615
R1528 VDD2.n29 VDD2.n7 104.615
R1529 VDD2.n31 VDD2.n29 104.615
R1530 VDD2.n31 VDD2.n30 104.615
R1531 VDD2.n30 VDD2.n3 104.615
R1532 VDD2.n39 VDD2.n3 104.615
R1533 VDD2.n40 VDD2.n39 104.615
R1534 VDD2.n46 VDD2.n45 65.7496
R1535 VDD2 VDD2.n93 65.7468
R1536 VDD2.n62 VDD2.t4 52.3082
R1537 VDD2.n14 VDD2.t3 52.3082
R1538 VDD2.n46 VDD2.n44 51.6339
R1539 VDD2.n92 VDD2.n91 50.9975
R1540 VDD2.n92 VDD2.n46 34.1528
R1541 VDD2.n85 VDD2.n84 13.1884
R1542 VDD2.n38 VDD2.n37 13.1884
R1543 VDD2.n88 VDD2.n49 12.8005
R1544 VDD2.n83 VDD2.n51 12.8005
R1545 VDD2.n36 VDD2.n4 12.8005
R1546 VDD2.n41 VDD2.n2 12.8005
R1547 VDD2.n89 VDD2.n47 12.0247
R1548 VDD2.n80 VDD2.n79 12.0247
R1549 VDD2.n33 VDD2.n32 12.0247
R1550 VDD2.n42 VDD2.n0 12.0247
R1551 VDD2.n76 VDD2.n53 11.249
R1552 VDD2.n28 VDD2.n6 11.249
R1553 VDD2.n75 VDD2.n56 10.4732
R1554 VDD2.n27 VDD2.n8 10.4732
R1555 VDD2.n63 VDD2.n61 10.2747
R1556 VDD2.n15 VDD2.n13 10.2747
R1557 VDD2.n72 VDD2.n71 9.69747
R1558 VDD2.n24 VDD2.n23 9.69747
R1559 VDD2.n91 VDD2.n90 9.45567
R1560 VDD2.n44 VDD2.n43 9.45567
R1561 VDD2.n65 VDD2.n64 9.3005
R1562 VDD2.n67 VDD2.n66 9.3005
R1563 VDD2.n58 VDD2.n57 9.3005
R1564 VDD2.n73 VDD2.n72 9.3005
R1565 VDD2.n75 VDD2.n74 9.3005
R1566 VDD2.n53 VDD2.n52 9.3005
R1567 VDD2.n81 VDD2.n80 9.3005
R1568 VDD2.n83 VDD2.n82 9.3005
R1569 VDD2.n90 VDD2.n89 9.3005
R1570 VDD2.n49 VDD2.n48 9.3005
R1571 VDD2.n43 VDD2.n42 9.3005
R1572 VDD2.n2 VDD2.n1 9.3005
R1573 VDD2.n17 VDD2.n16 9.3005
R1574 VDD2.n19 VDD2.n18 9.3005
R1575 VDD2.n10 VDD2.n9 9.3005
R1576 VDD2.n25 VDD2.n24 9.3005
R1577 VDD2.n27 VDD2.n26 9.3005
R1578 VDD2.n6 VDD2.n5 9.3005
R1579 VDD2.n34 VDD2.n33 9.3005
R1580 VDD2.n36 VDD2.n35 9.3005
R1581 VDD2.n68 VDD2.n58 8.92171
R1582 VDD2.n20 VDD2.n10 8.92171
R1583 VDD2.n67 VDD2.n60 8.14595
R1584 VDD2.n19 VDD2.n12 8.14595
R1585 VDD2.n64 VDD2.n63 7.3702
R1586 VDD2.n16 VDD2.n15 7.3702
R1587 VDD2.n64 VDD2.n60 5.81868
R1588 VDD2.n16 VDD2.n12 5.81868
R1589 VDD2.n68 VDD2.n67 5.04292
R1590 VDD2.n20 VDD2.n19 5.04292
R1591 VDD2.n71 VDD2.n58 4.26717
R1592 VDD2.n23 VDD2.n10 4.26717
R1593 VDD2.n72 VDD2.n56 3.49141
R1594 VDD2.n24 VDD2.n8 3.49141
R1595 VDD2.n17 VDD2.n13 2.84303
R1596 VDD2.n65 VDD2.n61 2.84303
R1597 VDD2.n76 VDD2.n75 2.71565
R1598 VDD2.n28 VDD2.n27 2.71565
R1599 VDD2.n93 VDD2.t2 2.29482
R1600 VDD2.n93 VDD2.t1 2.29482
R1601 VDD2.n45 VDD2.t0 2.29482
R1602 VDD2.n45 VDD2.t5 2.29482
R1603 VDD2.n91 VDD2.n47 1.93989
R1604 VDD2.n79 VDD2.n53 1.93989
R1605 VDD2.n32 VDD2.n6 1.93989
R1606 VDD2.n44 VDD2.n0 1.93989
R1607 VDD2.n89 VDD2.n88 1.16414
R1608 VDD2.n80 VDD2.n51 1.16414
R1609 VDD2.n33 VDD2.n4 1.16414
R1610 VDD2.n42 VDD2.n41 1.16414
R1611 VDD2 VDD2.n92 0.7505
R1612 VDD2.n85 VDD2.n49 0.388379
R1613 VDD2.n84 VDD2.n83 0.388379
R1614 VDD2.n37 VDD2.n36 0.388379
R1615 VDD2.n38 VDD2.n2 0.388379
R1616 VDD2.n90 VDD2.n48 0.155672
R1617 VDD2.n82 VDD2.n48 0.155672
R1618 VDD2.n82 VDD2.n81 0.155672
R1619 VDD2.n81 VDD2.n52 0.155672
R1620 VDD2.n74 VDD2.n52 0.155672
R1621 VDD2.n74 VDD2.n73 0.155672
R1622 VDD2.n73 VDD2.n57 0.155672
R1623 VDD2.n66 VDD2.n57 0.155672
R1624 VDD2.n66 VDD2.n65 0.155672
R1625 VDD2.n18 VDD2.n17 0.155672
R1626 VDD2.n18 VDD2.n9 0.155672
R1627 VDD2.n25 VDD2.n9 0.155672
R1628 VDD2.n26 VDD2.n25 0.155672
R1629 VDD2.n26 VDD2.n5 0.155672
R1630 VDD2.n34 VDD2.n5 0.155672
R1631 VDD2.n35 VDD2.n34 0.155672
R1632 VDD2.n35 VDD2.n1 0.155672
R1633 VDD2.n43 VDD2.n1 0.155672
C0 VN VTAIL 3.13368f
C1 VP VTAIL 3.14814f
C2 VDD1 VTAIL 7.53467f
C3 VP VN 4.49487f
C4 VN VDD1 0.148015f
C5 VDD2 VTAIL 7.571f
C6 VP VDD1 3.4495f
C7 VN VDD2 3.30052f
C8 VP VDD2 0.300313f
C9 VDD2 VDD1 0.723108f
C10 VDD2 B 3.914121f
C11 VDD1 B 3.9405f
C12 VTAIL B 5.185055f
C13 VN B 7.42609f
C14 VP B 5.657275f
C15 VDD2.n0 B 0.03131f
C16 VDD2.n1 B 0.023281f
C17 VDD2.n2 B 0.01251f
C18 VDD2.n3 B 0.029569f
C19 VDD2.n4 B 0.013246f
C20 VDD2.n5 B 0.023281f
C21 VDD2.n6 B 0.01251f
C22 VDD2.n7 B 0.029569f
C23 VDD2.n8 B 0.013246f
C24 VDD2.n9 B 0.023281f
C25 VDD2.n10 B 0.01251f
C26 VDD2.n11 B 0.029569f
C27 VDD2.n12 B 0.013246f
C28 VDD2.n13 B 0.137746f
C29 VDD2.t3 B 0.049526f
C30 VDD2.n14 B 0.022177f
C31 VDD2.n15 B 0.020903f
C32 VDD2.n16 B 0.01251f
C33 VDD2.n17 B 0.825498f
C34 VDD2.n18 B 0.023281f
C35 VDD2.n19 B 0.01251f
C36 VDD2.n20 B 0.013246f
C37 VDD2.n21 B 0.029569f
C38 VDD2.n22 B 0.029569f
C39 VDD2.n23 B 0.013246f
C40 VDD2.n24 B 0.01251f
C41 VDD2.n25 B 0.023281f
C42 VDD2.n26 B 0.023281f
C43 VDD2.n27 B 0.01251f
C44 VDD2.n28 B 0.013246f
C45 VDD2.n29 B 0.029569f
C46 VDD2.n30 B 0.029569f
C47 VDD2.n31 B 0.029569f
C48 VDD2.n32 B 0.013246f
C49 VDD2.n33 B 0.01251f
C50 VDD2.n34 B 0.023281f
C51 VDD2.n35 B 0.023281f
C52 VDD2.n36 B 0.01251f
C53 VDD2.n37 B 0.012878f
C54 VDD2.n38 B 0.012878f
C55 VDD2.n39 B 0.029569f
C56 VDD2.n40 B 0.061513f
C57 VDD2.n41 B 0.013246f
C58 VDD2.n42 B 0.01251f
C59 VDD2.n43 B 0.057311f
C60 VDD2.n44 B 0.051492f
C61 VDD2.t0 B 0.158769f
C62 VDD2.t5 B 0.158769f
C63 VDD2.n45 B 1.38474f
C64 VDD2.n46 B 1.54917f
C65 VDD2.n47 B 0.03131f
C66 VDD2.n48 B 0.023281f
C67 VDD2.n49 B 0.01251f
C68 VDD2.n50 B 0.029569f
C69 VDD2.n51 B 0.013246f
C70 VDD2.n52 B 0.023281f
C71 VDD2.n53 B 0.01251f
C72 VDD2.n54 B 0.029569f
C73 VDD2.n55 B 0.029569f
C74 VDD2.n56 B 0.013246f
C75 VDD2.n57 B 0.023281f
C76 VDD2.n58 B 0.01251f
C77 VDD2.n59 B 0.029569f
C78 VDD2.n60 B 0.013246f
C79 VDD2.n61 B 0.137746f
C80 VDD2.t4 B 0.049526f
C81 VDD2.n62 B 0.022177f
C82 VDD2.n63 B 0.020903f
C83 VDD2.n64 B 0.01251f
C84 VDD2.n65 B 0.825498f
C85 VDD2.n66 B 0.023281f
C86 VDD2.n67 B 0.01251f
C87 VDD2.n68 B 0.013246f
C88 VDD2.n69 B 0.029569f
C89 VDD2.n70 B 0.029569f
C90 VDD2.n71 B 0.013246f
C91 VDD2.n72 B 0.01251f
C92 VDD2.n73 B 0.023281f
C93 VDD2.n74 B 0.023281f
C94 VDD2.n75 B 0.01251f
C95 VDD2.n76 B 0.013246f
C96 VDD2.n77 B 0.029569f
C97 VDD2.n78 B 0.029569f
C98 VDD2.n79 B 0.013246f
C99 VDD2.n80 B 0.01251f
C100 VDD2.n81 B 0.023281f
C101 VDD2.n82 B 0.023281f
C102 VDD2.n83 B 0.01251f
C103 VDD2.n84 B 0.012878f
C104 VDD2.n85 B 0.012878f
C105 VDD2.n86 B 0.029569f
C106 VDD2.n87 B 0.061513f
C107 VDD2.n88 B 0.013246f
C108 VDD2.n89 B 0.01251f
C109 VDD2.n90 B 0.057311f
C110 VDD2.n91 B 0.050316f
C111 VDD2.n92 B 1.66817f
C112 VDD2.t2 B 0.158769f
C113 VDD2.t1 B 0.158769f
C114 VDD2.n93 B 1.38472f
C115 VN.n0 B 0.191167f
C116 VN.t2 B 0.854132f
C117 VN.n1 B 0.334369f
C118 VN.t5 B 0.832063f
C119 VN.n2 B 0.355393f
C120 VN.n3 B 0.010295f
C121 VN.t0 B 0.832063f
C122 VN.n4 B 0.349458f
C123 VN.n5 B 0.03516f
C124 VN.n6 B 0.191167f
C125 VN.t4 B 0.854132f
C126 VN.n7 B 0.334369f
C127 VN.t3 B 0.832063f
C128 VN.n8 B 0.355393f
C129 VN.n9 B 0.010295f
C130 VN.t1 B 0.832063f
C131 VN.n10 B 0.349458f
C132 VN.n11 B 1.66811f
C133 VDD1.n0 B 0.031065f
C134 VDD1.n1 B 0.023099f
C135 VDD1.n2 B 0.012412f
C136 VDD1.n3 B 0.029338f
C137 VDD1.n4 B 0.013142f
C138 VDD1.n5 B 0.023099f
C139 VDD1.n6 B 0.012412f
C140 VDD1.n7 B 0.029338f
C141 VDD1.n8 B 0.029338f
C142 VDD1.n9 B 0.013142f
C143 VDD1.n10 B 0.023099f
C144 VDD1.n11 B 0.012412f
C145 VDD1.n12 B 0.029338f
C146 VDD1.n13 B 0.013142f
C147 VDD1.n14 B 0.136668f
C148 VDD1.t2 B 0.049139f
C149 VDD1.n15 B 0.022004f
C150 VDD1.n16 B 0.02074f
C151 VDD1.n17 B 0.012412f
C152 VDD1.n18 B 0.819037f
C153 VDD1.n19 B 0.023099f
C154 VDD1.n20 B 0.012412f
C155 VDD1.n21 B 0.013142f
C156 VDD1.n22 B 0.029338f
C157 VDD1.n23 B 0.029338f
C158 VDD1.n24 B 0.013142f
C159 VDD1.n25 B 0.012412f
C160 VDD1.n26 B 0.023099f
C161 VDD1.n27 B 0.023099f
C162 VDD1.n28 B 0.012412f
C163 VDD1.n29 B 0.013142f
C164 VDD1.n30 B 0.029338f
C165 VDD1.n31 B 0.029338f
C166 VDD1.n32 B 0.013142f
C167 VDD1.n33 B 0.012412f
C168 VDD1.n34 B 0.023099f
C169 VDD1.n35 B 0.023099f
C170 VDD1.n36 B 0.012412f
C171 VDD1.n37 B 0.012777f
C172 VDD1.n38 B 0.012777f
C173 VDD1.n39 B 0.029338f
C174 VDD1.n40 B 0.061032f
C175 VDD1.n41 B 0.013142f
C176 VDD1.n42 B 0.012412f
C177 VDD1.n43 B 0.056863f
C178 VDD1.n44 B 0.051405f
C179 VDD1.n45 B 0.031065f
C180 VDD1.n46 B 0.023099f
C181 VDD1.n47 B 0.012412f
C182 VDD1.n48 B 0.029338f
C183 VDD1.n49 B 0.013142f
C184 VDD1.n50 B 0.023099f
C185 VDD1.n51 B 0.012412f
C186 VDD1.n52 B 0.029338f
C187 VDD1.n53 B 0.013142f
C188 VDD1.n54 B 0.023099f
C189 VDD1.n55 B 0.012412f
C190 VDD1.n56 B 0.029338f
C191 VDD1.n57 B 0.013142f
C192 VDD1.n58 B 0.136668f
C193 VDD1.t5 B 0.049139f
C194 VDD1.n59 B 0.022004f
C195 VDD1.n60 B 0.02074f
C196 VDD1.n61 B 0.012412f
C197 VDD1.n62 B 0.819037f
C198 VDD1.n63 B 0.023099f
C199 VDD1.n64 B 0.012412f
C200 VDD1.n65 B 0.013142f
C201 VDD1.n66 B 0.029338f
C202 VDD1.n67 B 0.029338f
C203 VDD1.n68 B 0.013142f
C204 VDD1.n69 B 0.012412f
C205 VDD1.n70 B 0.023099f
C206 VDD1.n71 B 0.023099f
C207 VDD1.n72 B 0.012412f
C208 VDD1.n73 B 0.013142f
C209 VDD1.n74 B 0.029338f
C210 VDD1.n75 B 0.029338f
C211 VDD1.n76 B 0.029338f
C212 VDD1.n77 B 0.013142f
C213 VDD1.n78 B 0.012412f
C214 VDD1.n79 B 0.023099f
C215 VDD1.n80 B 0.023099f
C216 VDD1.n81 B 0.012412f
C217 VDD1.n82 B 0.012777f
C218 VDD1.n83 B 0.012777f
C219 VDD1.n84 B 0.029338f
C220 VDD1.n85 B 0.061032f
C221 VDD1.n86 B 0.013142f
C222 VDD1.n87 B 0.012412f
C223 VDD1.n88 B 0.056863f
C224 VDD1.n89 B 0.051089f
C225 VDD1.t0 B 0.157526f
C226 VDD1.t4 B 0.157526f
C227 VDD1.n90 B 1.37391f
C228 VDD1.n91 B 1.60795f
C229 VDD1.t1 B 0.157526f
C230 VDD1.t3 B 0.157526f
C231 VDD1.n92 B 1.37316f
C232 VDD1.n93 B 1.84253f
C233 VTAIL.t3 B 0.168633f
C234 VTAIL.t11 B 0.168633f
C235 VTAIL.n0 B 1.40421f
C236 VTAIL.n1 B 0.326857f
C237 VTAIL.n2 B 0.033255f
C238 VTAIL.n3 B 0.024727f
C239 VTAIL.n4 B 0.013287f
C240 VTAIL.n5 B 0.031407f
C241 VTAIL.n6 B 0.014069f
C242 VTAIL.n7 B 0.024727f
C243 VTAIL.n8 B 0.013287f
C244 VTAIL.n9 B 0.031407f
C245 VTAIL.n10 B 0.014069f
C246 VTAIL.n11 B 0.024727f
C247 VTAIL.n12 B 0.013287f
C248 VTAIL.n13 B 0.031407f
C249 VTAIL.n14 B 0.014069f
C250 VTAIL.n15 B 0.146304f
C251 VTAIL.t6 B 0.052603f
C252 VTAIL.n16 B 0.023555f
C253 VTAIL.n17 B 0.022202f
C254 VTAIL.n18 B 0.013287f
C255 VTAIL.n19 B 0.876783f
C256 VTAIL.n20 B 0.024727f
C257 VTAIL.n21 B 0.013287f
C258 VTAIL.n22 B 0.014069f
C259 VTAIL.n23 B 0.031407f
C260 VTAIL.n24 B 0.031407f
C261 VTAIL.n25 B 0.014069f
C262 VTAIL.n26 B 0.013287f
C263 VTAIL.n27 B 0.024727f
C264 VTAIL.n28 B 0.024727f
C265 VTAIL.n29 B 0.013287f
C266 VTAIL.n30 B 0.014069f
C267 VTAIL.n31 B 0.031407f
C268 VTAIL.n32 B 0.031407f
C269 VTAIL.n33 B 0.031407f
C270 VTAIL.n34 B 0.014069f
C271 VTAIL.n35 B 0.013287f
C272 VTAIL.n36 B 0.024727f
C273 VTAIL.n37 B 0.024727f
C274 VTAIL.n38 B 0.013287f
C275 VTAIL.n39 B 0.013678f
C276 VTAIL.n40 B 0.013678f
C277 VTAIL.n41 B 0.031407f
C278 VTAIL.n42 B 0.065335f
C279 VTAIL.n43 B 0.014069f
C280 VTAIL.n44 B 0.013287f
C281 VTAIL.n45 B 0.060872f
C282 VTAIL.n46 B 0.036395f
C283 VTAIL.n47 B 0.170897f
C284 VTAIL.t7 B 0.168633f
C285 VTAIL.t10 B 0.168633f
C286 VTAIL.n48 B 1.40421f
C287 VTAIL.n49 B 1.37881f
C288 VTAIL.t4 B 0.168633f
C289 VTAIL.t1 B 0.168633f
C290 VTAIL.n50 B 1.40422f
C291 VTAIL.n51 B 1.3788f
C292 VTAIL.n52 B 0.033255f
C293 VTAIL.n53 B 0.024727f
C294 VTAIL.n54 B 0.013287f
C295 VTAIL.n55 B 0.031407f
C296 VTAIL.n56 B 0.014069f
C297 VTAIL.n57 B 0.024727f
C298 VTAIL.n58 B 0.013287f
C299 VTAIL.n59 B 0.031407f
C300 VTAIL.n60 B 0.031407f
C301 VTAIL.n61 B 0.014069f
C302 VTAIL.n62 B 0.024727f
C303 VTAIL.n63 B 0.013287f
C304 VTAIL.n64 B 0.031407f
C305 VTAIL.n65 B 0.014069f
C306 VTAIL.n66 B 0.146304f
C307 VTAIL.t0 B 0.052603f
C308 VTAIL.n67 B 0.023555f
C309 VTAIL.n68 B 0.022202f
C310 VTAIL.n69 B 0.013287f
C311 VTAIL.n70 B 0.876783f
C312 VTAIL.n71 B 0.024727f
C313 VTAIL.n72 B 0.013287f
C314 VTAIL.n73 B 0.014069f
C315 VTAIL.n74 B 0.031407f
C316 VTAIL.n75 B 0.031407f
C317 VTAIL.n76 B 0.014069f
C318 VTAIL.n77 B 0.013287f
C319 VTAIL.n78 B 0.024727f
C320 VTAIL.n79 B 0.024727f
C321 VTAIL.n80 B 0.013287f
C322 VTAIL.n81 B 0.014069f
C323 VTAIL.n82 B 0.031407f
C324 VTAIL.n83 B 0.031407f
C325 VTAIL.n84 B 0.014069f
C326 VTAIL.n85 B 0.013287f
C327 VTAIL.n86 B 0.024727f
C328 VTAIL.n87 B 0.024727f
C329 VTAIL.n88 B 0.013287f
C330 VTAIL.n89 B 0.013678f
C331 VTAIL.n90 B 0.013678f
C332 VTAIL.n91 B 0.031407f
C333 VTAIL.n92 B 0.065335f
C334 VTAIL.n93 B 0.014069f
C335 VTAIL.n94 B 0.013287f
C336 VTAIL.n95 B 0.060872f
C337 VTAIL.n96 B 0.036395f
C338 VTAIL.n97 B 0.170897f
C339 VTAIL.t5 B 0.168633f
C340 VTAIL.t9 B 0.168633f
C341 VTAIL.n98 B 1.40422f
C342 VTAIL.n99 B 0.377333f
C343 VTAIL.n100 B 0.033255f
C344 VTAIL.n101 B 0.024727f
C345 VTAIL.n102 B 0.013287f
C346 VTAIL.n103 B 0.031407f
C347 VTAIL.n104 B 0.014069f
C348 VTAIL.n105 B 0.024727f
C349 VTAIL.n106 B 0.013287f
C350 VTAIL.n107 B 0.031407f
C351 VTAIL.n108 B 0.031407f
C352 VTAIL.n109 B 0.014069f
C353 VTAIL.n110 B 0.024727f
C354 VTAIL.n111 B 0.013287f
C355 VTAIL.n112 B 0.031407f
C356 VTAIL.n113 B 0.014069f
C357 VTAIL.n114 B 0.146304f
C358 VTAIL.t8 B 0.052603f
C359 VTAIL.n115 B 0.023555f
C360 VTAIL.n116 B 0.022202f
C361 VTAIL.n117 B 0.013287f
C362 VTAIL.n118 B 0.876783f
C363 VTAIL.n119 B 0.024727f
C364 VTAIL.n120 B 0.013287f
C365 VTAIL.n121 B 0.014069f
C366 VTAIL.n122 B 0.031407f
C367 VTAIL.n123 B 0.031407f
C368 VTAIL.n124 B 0.014069f
C369 VTAIL.n125 B 0.013287f
C370 VTAIL.n126 B 0.024727f
C371 VTAIL.n127 B 0.024727f
C372 VTAIL.n128 B 0.013287f
C373 VTAIL.n129 B 0.014069f
C374 VTAIL.n130 B 0.031407f
C375 VTAIL.n131 B 0.031407f
C376 VTAIL.n132 B 0.014069f
C377 VTAIL.n133 B 0.013287f
C378 VTAIL.n134 B 0.024727f
C379 VTAIL.n135 B 0.024727f
C380 VTAIL.n136 B 0.013287f
C381 VTAIL.n137 B 0.013678f
C382 VTAIL.n138 B 0.013678f
C383 VTAIL.n139 B 0.031407f
C384 VTAIL.n140 B 0.065335f
C385 VTAIL.n141 B 0.014069f
C386 VTAIL.n142 B 0.013287f
C387 VTAIL.n143 B 0.060872f
C388 VTAIL.n144 B 0.036395f
C389 VTAIL.n145 B 1.09887f
C390 VTAIL.n146 B 0.033255f
C391 VTAIL.n147 B 0.024727f
C392 VTAIL.n148 B 0.013287f
C393 VTAIL.n149 B 0.031407f
C394 VTAIL.n150 B 0.014069f
C395 VTAIL.n151 B 0.024727f
C396 VTAIL.n152 B 0.013287f
C397 VTAIL.n153 B 0.031407f
C398 VTAIL.n154 B 0.014069f
C399 VTAIL.n155 B 0.024727f
C400 VTAIL.n156 B 0.013287f
C401 VTAIL.n157 B 0.031407f
C402 VTAIL.n158 B 0.014069f
C403 VTAIL.n159 B 0.146304f
C404 VTAIL.t2 B 0.052603f
C405 VTAIL.n160 B 0.023555f
C406 VTAIL.n161 B 0.022202f
C407 VTAIL.n162 B 0.013287f
C408 VTAIL.n163 B 0.876783f
C409 VTAIL.n164 B 0.024727f
C410 VTAIL.n165 B 0.013287f
C411 VTAIL.n166 B 0.014069f
C412 VTAIL.n167 B 0.031407f
C413 VTAIL.n168 B 0.031407f
C414 VTAIL.n169 B 0.014069f
C415 VTAIL.n170 B 0.013287f
C416 VTAIL.n171 B 0.024727f
C417 VTAIL.n172 B 0.024727f
C418 VTAIL.n173 B 0.013287f
C419 VTAIL.n174 B 0.014069f
C420 VTAIL.n175 B 0.031407f
C421 VTAIL.n176 B 0.031407f
C422 VTAIL.n177 B 0.031407f
C423 VTAIL.n178 B 0.014069f
C424 VTAIL.n179 B 0.013287f
C425 VTAIL.n180 B 0.024727f
C426 VTAIL.n181 B 0.024727f
C427 VTAIL.n182 B 0.013287f
C428 VTAIL.n183 B 0.013678f
C429 VTAIL.n184 B 0.013678f
C430 VTAIL.n185 B 0.031407f
C431 VTAIL.n186 B 0.065335f
C432 VTAIL.n187 B 0.014069f
C433 VTAIL.n188 B 0.013287f
C434 VTAIL.n189 B 0.060872f
C435 VTAIL.n190 B 0.036395f
C436 VTAIL.n191 B 1.07586f
C437 VP.n0 B 0.046056f
C438 VP.n1 B 0.010451f
C439 VP.n2 B 0.194056f
C440 VP.t2 B 0.844639f
C441 VP.t4 B 0.844639f
C442 VP.t3 B 0.867042f
C443 VP.n3 B 0.339423f
C444 VP.n4 B 0.360764f
C445 VP.n5 B 0.010451f
C446 VP.n6 B 0.354739f
C447 VP.n7 B 1.66294f
C448 VP.t0 B 0.844639f
C449 VP.n8 B 0.354739f
C450 VP.n9 B 1.70556f
C451 VP.n10 B 0.046056f
C452 VP.n11 B 0.046056f
C453 VP.t5 B 0.844639f
C454 VP.n12 B 0.356443f
C455 VP.n13 B 0.010451f
C456 VP.t1 B 0.844639f
C457 VP.n14 B 0.354739f
C458 VP.n15 B 0.035691f
.ends

