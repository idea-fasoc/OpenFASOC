* NGSPICE file created from diff_pair_sample_1310.ext - technology: sky130A

.subckt diff_pair_sample_1310 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t13 VP.t0 VDD1.t6 w_n4942_n2748# sky130_fd_pr__pfet_01v8 ad=1.4685 pd=9.23 as=1.4685 ps=9.23 w=8.9 l=2.98
X1 VDD2.t9 VN.t0 VTAIL.t1 w_n4942_n2748# sky130_fd_pr__pfet_01v8 ad=1.4685 pd=9.23 as=1.4685 ps=9.23 w=8.9 l=2.98
X2 VDD1.t5 VP.t1 VTAIL.t12 w_n4942_n2748# sky130_fd_pr__pfet_01v8 ad=1.4685 pd=9.23 as=1.4685 ps=9.23 w=8.9 l=2.98
X3 VDD2.t8 VN.t1 VTAIL.t0 w_n4942_n2748# sky130_fd_pr__pfet_01v8 ad=1.4685 pd=9.23 as=3.471 ps=18.58 w=8.9 l=2.98
X4 VDD1.t8 VP.t2 VTAIL.t11 w_n4942_n2748# sky130_fd_pr__pfet_01v8 ad=1.4685 pd=9.23 as=3.471 ps=18.58 w=8.9 l=2.98
X5 VDD2.t7 VN.t2 VTAIL.t16 w_n4942_n2748# sky130_fd_pr__pfet_01v8 ad=3.471 pd=18.58 as=1.4685 ps=9.23 w=8.9 l=2.98
X6 B.t11 B.t9 B.t10 w_n4942_n2748# sky130_fd_pr__pfet_01v8 ad=3.471 pd=18.58 as=0 ps=0 w=8.9 l=2.98
X7 VDD2.t6 VN.t3 VTAIL.t3 w_n4942_n2748# sky130_fd_pr__pfet_01v8 ad=1.4685 pd=9.23 as=3.471 ps=18.58 w=8.9 l=2.98
X8 B.t8 B.t6 B.t7 w_n4942_n2748# sky130_fd_pr__pfet_01v8 ad=3.471 pd=18.58 as=0 ps=0 w=8.9 l=2.98
X9 B.t5 B.t3 B.t4 w_n4942_n2748# sky130_fd_pr__pfet_01v8 ad=3.471 pd=18.58 as=0 ps=0 w=8.9 l=2.98
X10 B.t2 B.t0 B.t1 w_n4942_n2748# sky130_fd_pr__pfet_01v8 ad=3.471 pd=18.58 as=0 ps=0 w=8.9 l=2.98
X11 VTAIL.t2 VN.t4 VDD2.t5 w_n4942_n2748# sky130_fd_pr__pfet_01v8 ad=1.4685 pd=9.23 as=1.4685 ps=9.23 w=8.9 l=2.98
X12 VTAIL.t10 VP.t3 VDD1.t9 w_n4942_n2748# sky130_fd_pr__pfet_01v8 ad=1.4685 pd=9.23 as=1.4685 ps=9.23 w=8.9 l=2.98
X13 VTAIL.t14 VN.t5 VDD2.t4 w_n4942_n2748# sky130_fd_pr__pfet_01v8 ad=1.4685 pd=9.23 as=1.4685 ps=9.23 w=8.9 l=2.98
X14 VDD1.t1 VP.t4 VTAIL.t9 w_n4942_n2748# sky130_fd_pr__pfet_01v8 ad=1.4685 pd=9.23 as=1.4685 ps=9.23 w=8.9 l=2.98
X15 VTAIL.t8 VP.t5 VDD1.t2 w_n4942_n2748# sky130_fd_pr__pfet_01v8 ad=1.4685 pd=9.23 as=1.4685 ps=9.23 w=8.9 l=2.98
X16 VDD2.t3 VN.t6 VTAIL.t18 w_n4942_n2748# sky130_fd_pr__pfet_01v8 ad=1.4685 pd=9.23 as=1.4685 ps=9.23 w=8.9 l=2.98
X17 VTAIL.t15 VN.t7 VDD2.t2 w_n4942_n2748# sky130_fd_pr__pfet_01v8 ad=1.4685 pd=9.23 as=1.4685 ps=9.23 w=8.9 l=2.98
X18 VDD1.t0 VP.t6 VTAIL.t7 w_n4942_n2748# sky130_fd_pr__pfet_01v8 ad=1.4685 pd=9.23 as=3.471 ps=18.58 w=8.9 l=2.98
X19 VDD1.t7 VP.t7 VTAIL.t6 w_n4942_n2748# sky130_fd_pr__pfet_01v8 ad=3.471 pd=18.58 as=1.4685 ps=9.23 w=8.9 l=2.98
X20 VTAIL.t19 VN.t8 VDD2.t1 w_n4942_n2748# sky130_fd_pr__pfet_01v8 ad=1.4685 pd=9.23 as=1.4685 ps=9.23 w=8.9 l=2.98
X21 VDD2.t0 VN.t9 VTAIL.t17 w_n4942_n2748# sky130_fd_pr__pfet_01v8 ad=3.471 pd=18.58 as=1.4685 ps=9.23 w=8.9 l=2.98
X22 VTAIL.t5 VP.t8 VDD1.t3 w_n4942_n2748# sky130_fd_pr__pfet_01v8 ad=1.4685 pd=9.23 as=1.4685 ps=9.23 w=8.9 l=2.98
X23 VDD1.t4 VP.t9 VTAIL.t4 w_n4942_n2748# sky130_fd_pr__pfet_01v8 ad=3.471 pd=18.58 as=1.4685 ps=9.23 w=8.9 l=2.98
R0 VP.n27 VP.n24 161.3
R1 VP.n29 VP.n28 161.3
R2 VP.n30 VP.n23 161.3
R3 VP.n32 VP.n31 161.3
R4 VP.n33 VP.n22 161.3
R5 VP.n35 VP.n34 161.3
R6 VP.n36 VP.n21 161.3
R7 VP.n39 VP.n38 161.3
R8 VP.n40 VP.n20 161.3
R9 VP.n42 VP.n41 161.3
R10 VP.n43 VP.n19 161.3
R11 VP.n45 VP.n44 161.3
R12 VP.n46 VP.n18 161.3
R13 VP.n48 VP.n47 161.3
R14 VP.n50 VP.n17 161.3
R15 VP.n52 VP.n51 161.3
R16 VP.n53 VP.n16 161.3
R17 VP.n55 VP.n54 161.3
R18 VP.n56 VP.n15 161.3
R19 VP.n58 VP.n57 161.3
R20 VP.n103 VP.n102 161.3
R21 VP.n101 VP.n1 161.3
R22 VP.n100 VP.n99 161.3
R23 VP.n98 VP.n2 161.3
R24 VP.n97 VP.n96 161.3
R25 VP.n95 VP.n3 161.3
R26 VP.n93 VP.n92 161.3
R27 VP.n91 VP.n4 161.3
R28 VP.n90 VP.n89 161.3
R29 VP.n88 VP.n5 161.3
R30 VP.n87 VP.n86 161.3
R31 VP.n85 VP.n6 161.3
R32 VP.n84 VP.n83 161.3
R33 VP.n81 VP.n7 161.3
R34 VP.n80 VP.n79 161.3
R35 VP.n78 VP.n8 161.3
R36 VP.n77 VP.n76 161.3
R37 VP.n75 VP.n9 161.3
R38 VP.n74 VP.n73 161.3
R39 VP.n72 VP.n10 161.3
R40 VP.n71 VP.n70 161.3
R41 VP.n68 VP.n11 161.3
R42 VP.n67 VP.n66 161.3
R43 VP.n65 VP.n12 161.3
R44 VP.n64 VP.n63 161.3
R45 VP.n62 VP.n13 161.3
R46 VP.n26 VP.t7 103.49
R47 VP.n61 VP.t9 71.977
R48 VP.n69 VP.t3 71.977
R49 VP.n82 VP.t1 71.977
R50 VP.n94 VP.t8 71.977
R51 VP.n0 VP.t2 71.977
R52 VP.n14 VP.t6 71.977
R53 VP.n49 VP.t0 71.977
R54 VP.n37 VP.t4 71.977
R55 VP.n25 VP.t5 71.977
R56 VP.n61 VP.n60 71.8769
R57 VP.n104 VP.n0 71.8769
R58 VP.n59 VP.n14 71.8769
R59 VP.n26 VP.n25 70.3732
R60 VP.n67 VP.n12 56.4773
R61 VP.n100 VP.n2 56.4773
R62 VP.n55 VP.n16 56.4773
R63 VP.n60 VP.n59 52.9196
R64 VP.n76 VP.n8 49.6611
R65 VP.n88 VP.n87 49.6611
R66 VP.n43 VP.n42 49.6611
R67 VP.n31 VP.n22 49.6611
R68 VP.n76 VP.n75 31.1601
R69 VP.n89 VP.n88 31.1601
R70 VP.n44 VP.n43 31.1601
R71 VP.n31 VP.n30 31.1601
R72 VP.n63 VP.n62 24.3439
R73 VP.n63 VP.n12 24.3439
R74 VP.n68 VP.n67 24.3439
R75 VP.n70 VP.n68 24.3439
R76 VP.n74 VP.n10 24.3439
R77 VP.n75 VP.n74 24.3439
R78 VP.n80 VP.n8 24.3439
R79 VP.n81 VP.n80 24.3439
R80 VP.n83 VP.n6 24.3439
R81 VP.n87 VP.n6 24.3439
R82 VP.n89 VP.n4 24.3439
R83 VP.n93 VP.n4 24.3439
R84 VP.n96 VP.n95 24.3439
R85 VP.n96 VP.n2 24.3439
R86 VP.n101 VP.n100 24.3439
R87 VP.n102 VP.n101 24.3439
R88 VP.n56 VP.n55 24.3439
R89 VP.n57 VP.n56 24.3439
R90 VP.n44 VP.n18 24.3439
R91 VP.n48 VP.n18 24.3439
R92 VP.n51 VP.n50 24.3439
R93 VP.n51 VP.n16 24.3439
R94 VP.n35 VP.n22 24.3439
R95 VP.n36 VP.n35 24.3439
R96 VP.n38 VP.n20 24.3439
R97 VP.n42 VP.n20 24.3439
R98 VP.n29 VP.n24 24.3439
R99 VP.n30 VP.n29 24.3439
R100 VP.n70 VP.n69 21.4227
R101 VP.n95 VP.n94 21.4227
R102 VP.n50 VP.n49 21.4227
R103 VP.n62 VP.n61 18.0146
R104 VP.n102 VP.n0 18.0146
R105 VP.n57 VP.n14 18.0146
R106 VP.n82 VP.n81 12.1722
R107 VP.n83 VP.n82 12.1722
R108 VP.n37 VP.n36 12.1722
R109 VP.n38 VP.n37 12.1722
R110 VP.n27 VP.n26 5.7067
R111 VP.n69 VP.n10 2.92171
R112 VP.n94 VP.n93 2.92171
R113 VP.n49 VP.n48 2.92171
R114 VP.n25 VP.n24 2.92171
R115 VP.n59 VP.n58 0.355081
R116 VP.n60 VP.n13 0.355081
R117 VP.n104 VP.n103 0.355081
R118 VP VP.n104 0.26685
R119 VP.n28 VP.n27 0.189894
R120 VP.n28 VP.n23 0.189894
R121 VP.n32 VP.n23 0.189894
R122 VP.n33 VP.n32 0.189894
R123 VP.n34 VP.n33 0.189894
R124 VP.n34 VP.n21 0.189894
R125 VP.n39 VP.n21 0.189894
R126 VP.n40 VP.n39 0.189894
R127 VP.n41 VP.n40 0.189894
R128 VP.n41 VP.n19 0.189894
R129 VP.n45 VP.n19 0.189894
R130 VP.n46 VP.n45 0.189894
R131 VP.n47 VP.n46 0.189894
R132 VP.n47 VP.n17 0.189894
R133 VP.n52 VP.n17 0.189894
R134 VP.n53 VP.n52 0.189894
R135 VP.n54 VP.n53 0.189894
R136 VP.n54 VP.n15 0.189894
R137 VP.n58 VP.n15 0.189894
R138 VP.n64 VP.n13 0.189894
R139 VP.n65 VP.n64 0.189894
R140 VP.n66 VP.n65 0.189894
R141 VP.n66 VP.n11 0.189894
R142 VP.n71 VP.n11 0.189894
R143 VP.n72 VP.n71 0.189894
R144 VP.n73 VP.n72 0.189894
R145 VP.n73 VP.n9 0.189894
R146 VP.n77 VP.n9 0.189894
R147 VP.n78 VP.n77 0.189894
R148 VP.n79 VP.n78 0.189894
R149 VP.n79 VP.n7 0.189894
R150 VP.n84 VP.n7 0.189894
R151 VP.n85 VP.n84 0.189894
R152 VP.n86 VP.n85 0.189894
R153 VP.n86 VP.n5 0.189894
R154 VP.n90 VP.n5 0.189894
R155 VP.n91 VP.n90 0.189894
R156 VP.n92 VP.n91 0.189894
R157 VP.n92 VP.n3 0.189894
R158 VP.n97 VP.n3 0.189894
R159 VP.n98 VP.n97 0.189894
R160 VP.n99 VP.n98 0.189894
R161 VP.n99 VP.n1 0.189894
R162 VP.n103 VP.n1 0.189894
R163 VDD1.n1 VDD1.t7 86.2991
R164 VDD1.n3 VDD1.t4 86.2988
R165 VDD1.n5 VDD1.n4 81.8779
R166 VDD1.n1 VDD1.n0 79.7934
R167 VDD1.n7 VDD1.n6 79.7932
R168 VDD1.n3 VDD1.n2 79.7931
R169 VDD1.n7 VDD1.n5 46.9513
R170 VDD1.n6 VDD1.t6 3.65275
R171 VDD1.n6 VDD1.t0 3.65275
R172 VDD1.n0 VDD1.t2 3.65275
R173 VDD1.n0 VDD1.t1 3.65275
R174 VDD1.n4 VDD1.t3 3.65275
R175 VDD1.n4 VDD1.t8 3.65275
R176 VDD1.n2 VDD1.t9 3.65275
R177 VDD1.n2 VDD1.t5 3.65275
R178 VDD1 VDD1.n7 2.0824
R179 VDD1 VDD1.n1 0.772052
R180 VDD1.n5 VDD1.n3 0.658516
R181 VTAIL.n11 VTAIL.t3 66.7669
R182 VTAIL.n16 VTAIL.t7 66.7666
R183 VTAIL.n17 VTAIL.t0 66.7666
R184 VTAIL.n2 VTAIL.t11 66.7666
R185 VTAIL.n15 VTAIL.n14 63.1146
R186 VTAIL.n13 VTAIL.n12 63.1146
R187 VTAIL.n10 VTAIL.n9 63.1146
R188 VTAIL.n8 VTAIL.n7 63.1146
R189 VTAIL.n19 VTAIL.n18 63.1144
R190 VTAIL.n1 VTAIL.n0 63.1144
R191 VTAIL.n4 VTAIL.n3 63.1144
R192 VTAIL.n6 VTAIL.n5 63.1144
R193 VTAIL.n8 VTAIL.n6 25.7462
R194 VTAIL.n17 VTAIL.n16 22.8927
R195 VTAIL.n18 VTAIL.t1 3.65275
R196 VTAIL.n18 VTAIL.t15 3.65275
R197 VTAIL.n0 VTAIL.t16 3.65275
R198 VTAIL.n0 VTAIL.t2 3.65275
R199 VTAIL.n3 VTAIL.t12 3.65275
R200 VTAIL.n3 VTAIL.t5 3.65275
R201 VTAIL.n5 VTAIL.t4 3.65275
R202 VTAIL.n5 VTAIL.t10 3.65275
R203 VTAIL.n14 VTAIL.t9 3.65275
R204 VTAIL.n14 VTAIL.t13 3.65275
R205 VTAIL.n12 VTAIL.t6 3.65275
R206 VTAIL.n12 VTAIL.t8 3.65275
R207 VTAIL.n9 VTAIL.t18 3.65275
R208 VTAIL.n9 VTAIL.t14 3.65275
R209 VTAIL.n7 VTAIL.t17 3.65275
R210 VTAIL.n7 VTAIL.t19 3.65275
R211 VTAIL.n10 VTAIL.n8 2.85395
R212 VTAIL.n11 VTAIL.n10 2.85395
R213 VTAIL.n15 VTAIL.n13 2.85395
R214 VTAIL.n16 VTAIL.n15 2.85395
R215 VTAIL.n6 VTAIL.n4 2.85395
R216 VTAIL.n4 VTAIL.n2 2.85395
R217 VTAIL.n19 VTAIL.n17 2.85395
R218 VTAIL VTAIL.n1 2.19878
R219 VTAIL.n13 VTAIL.n11 1.89705
R220 VTAIL.n2 VTAIL.n1 1.89705
R221 VTAIL VTAIL.n19 0.655672
R222 VN.n90 VN.n89 161.3
R223 VN.n88 VN.n47 161.3
R224 VN.n87 VN.n86 161.3
R225 VN.n85 VN.n48 161.3
R226 VN.n84 VN.n83 161.3
R227 VN.n82 VN.n49 161.3
R228 VN.n80 VN.n79 161.3
R229 VN.n78 VN.n50 161.3
R230 VN.n77 VN.n76 161.3
R231 VN.n75 VN.n51 161.3
R232 VN.n74 VN.n73 161.3
R233 VN.n72 VN.n52 161.3
R234 VN.n71 VN.n70 161.3
R235 VN.n68 VN.n53 161.3
R236 VN.n67 VN.n66 161.3
R237 VN.n65 VN.n54 161.3
R238 VN.n64 VN.n63 161.3
R239 VN.n62 VN.n55 161.3
R240 VN.n61 VN.n60 161.3
R241 VN.n59 VN.n56 161.3
R242 VN.n44 VN.n43 161.3
R243 VN.n42 VN.n1 161.3
R244 VN.n41 VN.n40 161.3
R245 VN.n39 VN.n2 161.3
R246 VN.n38 VN.n37 161.3
R247 VN.n36 VN.n3 161.3
R248 VN.n34 VN.n33 161.3
R249 VN.n32 VN.n4 161.3
R250 VN.n31 VN.n30 161.3
R251 VN.n29 VN.n5 161.3
R252 VN.n28 VN.n27 161.3
R253 VN.n26 VN.n6 161.3
R254 VN.n25 VN.n24 161.3
R255 VN.n22 VN.n7 161.3
R256 VN.n21 VN.n20 161.3
R257 VN.n19 VN.n8 161.3
R258 VN.n18 VN.n17 161.3
R259 VN.n16 VN.n9 161.3
R260 VN.n15 VN.n14 161.3
R261 VN.n13 VN.n10 161.3
R262 VN.n58 VN.t3 103.49
R263 VN.n12 VN.t2 103.49
R264 VN.n11 VN.t4 71.977
R265 VN.n23 VN.t0 71.977
R266 VN.n35 VN.t7 71.977
R267 VN.n0 VN.t1 71.977
R268 VN.n57 VN.t5 71.977
R269 VN.n69 VN.t6 71.977
R270 VN.n81 VN.t8 71.977
R271 VN.n46 VN.t9 71.977
R272 VN.n45 VN.n0 71.8769
R273 VN.n91 VN.n46 71.8769
R274 VN.n12 VN.n11 70.3732
R275 VN.n58 VN.n57 70.3732
R276 VN.n41 VN.n2 56.4773
R277 VN.n87 VN.n48 56.4773
R278 VN VN.n91 53.085
R279 VN.n17 VN.n8 49.6611
R280 VN.n29 VN.n28 49.6611
R281 VN.n63 VN.n54 49.6611
R282 VN.n75 VN.n74 49.6611
R283 VN.n17 VN.n16 31.1601
R284 VN.n30 VN.n29 31.1601
R285 VN.n63 VN.n62 31.1601
R286 VN.n76 VN.n75 31.1601
R287 VN.n15 VN.n10 24.3439
R288 VN.n16 VN.n15 24.3439
R289 VN.n21 VN.n8 24.3439
R290 VN.n22 VN.n21 24.3439
R291 VN.n24 VN.n6 24.3439
R292 VN.n28 VN.n6 24.3439
R293 VN.n30 VN.n4 24.3439
R294 VN.n34 VN.n4 24.3439
R295 VN.n37 VN.n36 24.3439
R296 VN.n37 VN.n2 24.3439
R297 VN.n42 VN.n41 24.3439
R298 VN.n43 VN.n42 24.3439
R299 VN.n62 VN.n61 24.3439
R300 VN.n61 VN.n56 24.3439
R301 VN.n74 VN.n52 24.3439
R302 VN.n70 VN.n52 24.3439
R303 VN.n68 VN.n67 24.3439
R304 VN.n67 VN.n54 24.3439
R305 VN.n83 VN.n48 24.3439
R306 VN.n83 VN.n82 24.3439
R307 VN.n80 VN.n50 24.3439
R308 VN.n76 VN.n50 24.3439
R309 VN.n89 VN.n88 24.3439
R310 VN.n88 VN.n87 24.3439
R311 VN.n36 VN.n35 21.4227
R312 VN.n82 VN.n81 21.4227
R313 VN.n43 VN.n0 18.0146
R314 VN.n89 VN.n46 18.0146
R315 VN.n23 VN.n22 12.1722
R316 VN.n24 VN.n23 12.1722
R317 VN.n70 VN.n69 12.1722
R318 VN.n69 VN.n68 12.1722
R319 VN.n59 VN.n58 5.70674
R320 VN.n13 VN.n12 5.70674
R321 VN.n11 VN.n10 2.92171
R322 VN.n35 VN.n34 2.92171
R323 VN.n57 VN.n56 2.92171
R324 VN.n81 VN.n80 2.92171
R325 VN.n91 VN.n90 0.355081
R326 VN.n45 VN.n44 0.355081
R327 VN VN.n45 0.26685
R328 VN.n90 VN.n47 0.189894
R329 VN.n86 VN.n47 0.189894
R330 VN.n86 VN.n85 0.189894
R331 VN.n85 VN.n84 0.189894
R332 VN.n84 VN.n49 0.189894
R333 VN.n79 VN.n49 0.189894
R334 VN.n79 VN.n78 0.189894
R335 VN.n78 VN.n77 0.189894
R336 VN.n77 VN.n51 0.189894
R337 VN.n73 VN.n51 0.189894
R338 VN.n73 VN.n72 0.189894
R339 VN.n72 VN.n71 0.189894
R340 VN.n71 VN.n53 0.189894
R341 VN.n66 VN.n53 0.189894
R342 VN.n66 VN.n65 0.189894
R343 VN.n65 VN.n64 0.189894
R344 VN.n64 VN.n55 0.189894
R345 VN.n60 VN.n55 0.189894
R346 VN.n60 VN.n59 0.189894
R347 VN.n14 VN.n13 0.189894
R348 VN.n14 VN.n9 0.189894
R349 VN.n18 VN.n9 0.189894
R350 VN.n19 VN.n18 0.189894
R351 VN.n20 VN.n19 0.189894
R352 VN.n20 VN.n7 0.189894
R353 VN.n25 VN.n7 0.189894
R354 VN.n26 VN.n25 0.189894
R355 VN.n27 VN.n26 0.189894
R356 VN.n27 VN.n5 0.189894
R357 VN.n31 VN.n5 0.189894
R358 VN.n32 VN.n31 0.189894
R359 VN.n33 VN.n32 0.189894
R360 VN.n33 VN.n3 0.189894
R361 VN.n38 VN.n3 0.189894
R362 VN.n39 VN.n38 0.189894
R363 VN.n40 VN.n39 0.189894
R364 VN.n40 VN.n1 0.189894
R365 VN.n44 VN.n1 0.189894
R366 VDD2.n1 VDD2.t7 86.2988
R367 VDD2.n4 VDD2.t0 83.4457
R368 VDD2.n3 VDD2.n2 81.8779
R369 VDD2 VDD2.n7 81.8751
R370 VDD2.n6 VDD2.n5 79.7934
R371 VDD2.n1 VDD2.n0 79.7931
R372 VDD2.n4 VDD2.n3 44.9416
R373 VDD2.n7 VDD2.t4 3.65275
R374 VDD2.n7 VDD2.t6 3.65275
R375 VDD2.n5 VDD2.t1 3.65275
R376 VDD2.n5 VDD2.t3 3.65275
R377 VDD2.n2 VDD2.t2 3.65275
R378 VDD2.n2 VDD2.t8 3.65275
R379 VDD2.n0 VDD2.t5 3.65275
R380 VDD2.n0 VDD2.t9 3.65275
R381 VDD2.n6 VDD2.n4 2.85395
R382 VDD2 VDD2.n6 0.772052
R383 VDD2.n3 VDD2.n1 0.658516
R384 B.n429 B.n144 585
R385 B.n428 B.n427 585
R386 B.n426 B.n145 585
R387 B.n425 B.n424 585
R388 B.n423 B.n146 585
R389 B.n422 B.n421 585
R390 B.n420 B.n147 585
R391 B.n419 B.n418 585
R392 B.n417 B.n148 585
R393 B.n416 B.n415 585
R394 B.n414 B.n149 585
R395 B.n413 B.n412 585
R396 B.n411 B.n150 585
R397 B.n410 B.n409 585
R398 B.n408 B.n151 585
R399 B.n407 B.n406 585
R400 B.n405 B.n152 585
R401 B.n404 B.n403 585
R402 B.n402 B.n153 585
R403 B.n401 B.n400 585
R404 B.n399 B.n154 585
R405 B.n398 B.n397 585
R406 B.n396 B.n155 585
R407 B.n395 B.n394 585
R408 B.n393 B.n156 585
R409 B.n392 B.n391 585
R410 B.n390 B.n157 585
R411 B.n389 B.n388 585
R412 B.n387 B.n158 585
R413 B.n386 B.n385 585
R414 B.n384 B.n159 585
R415 B.n383 B.n382 585
R416 B.n381 B.n160 585
R417 B.n380 B.n379 585
R418 B.n375 B.n161 585
R419 B.n374 B.n373 585
R420 B.n372 B.n162 585
R421 B.n371 B.n370 585
R422 B.n369 B.n163 585
R423 B.n368 B.n367 585
R424 B.n366 B.n164 585
R425 B.n365 B.n364 585
R426 B.n362 B.n165 585
R427 B.n361 B.n360 585
R428 B.n359 B.n168 585
R429 B.n358 B.n357 585
R430 B.n356 B.n169 585
R431 B.n355 B.n354 585
R432 B.n353 B.n170 585
R433 B.n352 B.n351 585
R434 B.n350 B.n171 585
R435 B.n349 B.n348 585
R436 B.n347 B.n172 585
R437 B.n346 B.n345 585
R438 B.n344 B.n173 585
R439 B.n343 B.n342 585
R440 B.n341 B.n174 585
R441 B.n340 B.n339 585
R442 B.n338 B.n175 585
R443 B.n337 B.n336 585
R444 B.n335 B.n176 585
R445 B.n334 B.n333 585
R446 B.n332 B.n177 585
R447 B.n331 B.n330 585
R448 B.n329 B.n178 585
R449 B.n328 B.n327 585
R450 B.n326 B.n179 585
R451 B.n325 B.n324 585
R452 B.n323 B.n180 585
R453 B.n322 B.n321 585
R454 B.n320 B.n181 585
R455 B.n319 B.n318 585
R456 B.n317 B.n182 585
R457 B.n316 B.n315 585
R458 B.n314 B.n183 585
R459 B.n431 B.n430 585
R460 B.n432 B.n143 585
R461 B.n434 B.n433 585
R462 B.n435 B.n142 585
R463 B.n437 B.n436 585
R464 B.n438 B.n141 585
R465 B.n440 B.n439 585
R466 B.n441 B.n140 585
R467 B.n443 B.n442 585
R468 B.n444 B.n139 585
R469 B.n446 B.n445 585
R470 B.n447 B.n138 585
R471 B.n449 B.n448 585
R472 B.n450 B.n137 585
R473 B.n452 B.n451 585
R474 B.n453 B.n136 585
R475 B.n455 B.n454 585
R476 B.n456 B.n135 585
R477 B.n458 B.n457 585
R478 B.n459 B.n134 585
R479 B.n461 B.n460 585
R480 B.n462 B.n133 585
R481 B.n464 B.n463 585
R482 B.n465 B.n132 585
R483 B.n467 B.n466 585
R484 B.n468 B.n131 585
R485 B.n470 B.n469 585
R486 B.n471 B.n130 585
R487 B.n473 B.n472 585
R488 B.n474 B.n129 585
R489 B.n476 B.n475 585
R490 B.n477 B.n128 585
R491 B.n479 B.n478 585
R492 B.n480 B.n127 585
R493 B.n482 B.n481 585
R494 B.n483 B.n126 585
R495 B.n485 B.n484 585
R496 B.n486 B.n125 585
R497 B.n488 B.n487 585
R498 B.n489 B.n124 585
R499 B.n491 B.n490 585
R500 B.n492 B.n123 585
R501 B.n494 B.n493 585
R502 B.n495 B.n122 585
R503 B.n497 B.n496 585
R504 B.n498 B.n121 585
R505 B.n500 B.n499 585
R506 B.n501 B.n120 585
R507 B.n503 B.n502 585
R508 B.n504 B.n119 585
R509 B.n506 B.n505 585
R510 B.n507 B.n118 585
R511 B.n509 B.n508 585
R512 B.n510 B.n117 585
R513 B.n512 B.n511 585
R514 B.n513 B.n116 585
R515 B.n515 B.n514 585
R516 B.n516 B.n115 585
R517 B.n518 B.n517 585
R518 B.n519 B.n114 585
R519 B.n521 B.n520 585
R520 B.n522 B.n113 585
R521 B.n524 B.n523 585
R522 B.n525 B.n112 585
R523 B.n527 B.n526 585
R524 B.n528 B.n111 585
R525 B.n530 B.n529 585
R526 B.n531 B.n110 585
R527 B.n533 B.n532 585
R528 B.n534 B.n109 585
R529 B.n536 B.n535 585
R530 B.n537 B.n108 585
R531 B.n539 B.n538 585
R532 B.n540 B.n107 585
R533 B.n542 B.n541 585
R534 B.n543 B.n106 585
R535 B.n545 B.n544 585
R536 B.n546 B.n105 585
R537 B.n548 B.n547 585
R538 B.n549 B.n104 585
R539 B.n551 B.n550 585
R540 B.n552 B.n103 585
R541 B.n554 B.n553 585
R542 B.n555 B.n102 585
R543 B.n557 B.n556 585
R544 B.n558 B.n101 585
R545 B.n560 B.n559 585
R546 B.n561 B.n100 585
R547 B.n563 B.n562 585
R548 B.n564 B.n99 585
R549 B.n566 B.n565 585
R550 B.n567 B.n98 585
R551 B.n569 B.n568 585
R552 B.n570 B.n97 585
R553 B.n572 B.n571 585
R554 B.n573 B.n96 585
R555 B.n575 B.n574 585
R556 B.n576 B.n95 585
R557 B.n578 B.n577 585
R558 B.n579 B.n94 585
R559 B.n581 B.n580 585
R560 B.n582 B.n93 585
R561 B.n584 B.n583 585
R562 B.n585 B.n92 585
R563 B.n587 B.n586 585
R564 B.n588 B.n91 585
R565 B.n590 B.n589 585
R566 B.n591 B.n90 585
R567 B.n593 B.n592 585
R568 B.n594 B.n89 585
R569 B.n596 B.n595 585
R570 B.n597 B.n88 585
R571 B.n599 B.n598 585
R572 B.n600 B.n87 585
R573 B.n602 B.n601 585
R574 B.n603 B.n86 585
R575 B.n605 B.n604 585
R576 B.n606 B.n85 585
R577 B.n608 B.n607 585
R578 B.n609 B.n84 585
R579 B.n611 B.n610 585
R580 B.n612 B.n83 585
R581 B.n614 B.n613 585
R582 B.n615 B.n82 585
R583 B.n617 B.n616 585
R584 B.n618 B.n81 585
R585 B.n620 B.n619 585
R586 B.n621 B.n80 585
R587 B.n623 B.n622 585
R588 B.n624 B.n79 585
R589 B.n626 B.n625 585
R590 B.n627 B.n78 585
R591 B.n629 B.n628 585
R592 B.n630 B.n77 585
R593 B.n744 B.n35 585
R594 B.n743 B.n742 585
R595 B.n741 B.n36 585
R596 B.n740 B.n739 585
R597 B.n738 B.n37 585
R598 B.n737 B.n736 585
R599 B.n735 B.n38 585
R600 B.n734 B.n733 585
R601 B.n732 B.n39 585
R602 B.n731 B.n730 585
R603 B.n729 B.n40 585
R604 B.n728 B.n727 585
R605 B.n726 B.n41 585
R606 B.n725 B.n724 585
R607 B.n723 B.n42 585
R608 B.n722 B.n721 585
R609 B.n720 B.n43 585
R610 B.n719 B.n718 585
R611 B.n717 B.n44 585
R612 B.n716 B.n715 585
R613 B.n714 B.n45 585
R614 B.n713 B.n712 585
R615 B.n711 B.n46 585
R616 B.n710 B.n709 585
R617 B.n708 B.n47 585
R618 B.n707 B.n706 585
R619 B.n705 B.n48 585
R620 B.n704 B.n703 585
R621 B.n702 B.n49 585
R622 B.n701 B.n700 585
R623 B.n699 B.n50 585
R624 B.n698 B.n697 585
R625 B.n696 B.n51 585
R626 B.n694 B.n693 585
R627 B.n692 B.n54 585
R628 B.n691 B.n690 585
R629 B.n689 B.n55 585
R630 B.n688 B.n687 585
R631 B.n686 B.n56 585
R632 B.n685 B.n684 585
R633 B.n683 B.n57 585
R634 B.n682 B.n681 585
R635 B.n680 B.n679 585
R636 B.n678 B.n61 585
R637 B.n677 B.n676 585
R638 B.n675 B.n62 585
R639 B.n674 B.n673 585
R640 B.n672 B.n63 585
R641 B.n671 B.n670 585
R642 B.n669 B.n64 585
R643 B.n668 B.n667 585
R644 B.n666 B.n65 585
R645 B.n665 B.n664 585
R646 B.n663 B.n66 585
R647 B.n662 B.n661 585
R648 B.n660 B.n67 585
R649 B.n659 B.n658 585
R650 B.n657 B.n68 585
R651 B.n656 B.n655 585
R652 B.n654 B.n69 585
R653 B.n653 B.n652 585
R654 B.n651 B.n70 585
R655 B.n650 B.n649 585
R656 B.n648 B.n71 585
R657 B.n647 B.n646 585
R658 B.n645 B.n72 585
R659 B.n644 B.n643 585
R660 B.n642 B.n73 585
R661 B.n641 B.n640 585
R662 B.n639 B.n74 585
R663 B.n638 B.n637 585
R664 B.n636 B.n75 585
R665 B.n635 B.n634 585
R666 B.n633 B.n76 585
R667 B.n632 B.n631 585
R668 B.n746 B.n745 585
R669 B.n747 B.n34 585
R670 B.n749 B.n748 585
R671 B.n750 B.n33 585
R672 B.n752 B.n751 585
R673 B.n753 B.n32 585
R674 B.n755 B.n754 585
R675 B.n756 B.n31 585
R676 B.n758 B.n757 585
R677 B.n759 B.n30 585
R678 B.n761 B.n760 585
R679 B.n762 B.n29 585
R680 B.n764 B.n763 585
R681 B.n765 B.n28 585
R682 B.n767 B.n766 585
R683 B.n768 B.n27 585
R684 B.n770 B.n769 585
R685 B.n771 B.n26 585
R686 B.n773 B.n772 585
R687 B.n774 B.n25 585
R688 B.n776 B.n775 585
R689 B.n777 B.n24 585
R690 B.n779 B.n778 585
R691 B.n780 B.n23 585
R692 B.n782 B.n781 585
R693 B.n783 B.n22 585
R694 B.n785 B.n784 585
R695 B.n786 B.n21 585
R696 B.n788 B.n787 585
R697 B.n789 B.n20 585
R698 B.n791 B.n790 585
R699 B.n792 B.n19 585
R700 B.n794 B.n793 585
R701 B.n795 B.n18 585
R702 B.n797 B.n796 585
R703 B.n798 B.n17 585
R704 B.n800 B.n799 585
R705 B.n801 B.n16 585
R706 B.n803 B.n802 585
R707 B.n804 B.n15 585
R708 B.n806 B.n805 585
R709 B.n807 B.n14 585
R710 B.n809 B.n808 585
R711 B.n810 B.n13 585
R712 B.n812 B.n811 585
R713 B.n813 B.n12 585
R714 B.n815 B.n814 585
R715 B.n816 B.n11 585
R716 B.n818 B.n817 585
R717 B.n819 B.n10 585
R718 B.n821 B.n820 585
R719 B.n822 B.n9 585
R720 B.n824 B.n823 585
R721 B.n825 B.n8 585
R722 B.n827 B.n826 585
R723 B.n828 B.n7 585
R724 B.n830 B.n829 585
R725 B.n831 B.n6 585
R726 B.n833 B.n832 585
R727 B.n834 B.n5 585
R728 B.n836 B.n835 585
R729 B.n837 B.n4 585
R730 B.n839 B.n838 585
R731 B.n840 B.n3 585
R732 B.n842 B.n841 585
R733 B.n843 B.n0 585
R734 B.n2 B.n1 585
R735 B.n217 B.n216 585
R736 B.n218 B.n215 585
R737 B.n220 B.n219 585
R738 B.n221 B.n214 585
R739 B.n223 B.n222 585
R740 B.n224 B.n213 585
R741 B.n226 B.n225 585
R742 B.n227 B.n212 585
R743 B.n229 B.n228 585
R744 B.n230 B.n211 585
R745 B.n232 B.n231 585
R746 B.n233 B.n210 585
R747 B.n235 B.n234 585
R748 B.n236 B.n209 585
R749 B.n238 B.n237 585
R750 B.n239 B.n208 585
R751 B.n241 B.n240 585
R752 B.n242 B.n207 585
R753 B.n244 B.n243 585
R754 B.n245 B.n206 585
R755 B.n247 B.n246 585
R756 B.n248 B.n205 585
R757 B.n250 B.n249 585
R758 B.n251 B.n204 585
R759 B.n253 B.n252 585
R760 B.n254 B.n203 585
R761 B.n256 B.n255 585
R762 B.n257 B.n202 585
R763 B.n259 B.n258 585
R764 B.n260 B.n201 585
R765 B.n262 B.n261 585
R766 B.n263 B.n200 585
R767 B.n265 B.n264 585
R768 B.n266 B.n199 585
R769 B.n268 B.n267 585
R770 B.n269 B.n198 585
R771 B.n271 B.n270 585
R772 B.n272 B.n197 585
R773 B.n274 B.n273 585
R774 B.n275 B.n196 585
R775 B.n277 B.n276 585
R776 B.n278 B.n195 585
R777 B.n280 B.n279 585
R778 B.n281 B.n194 585
R779 B.n283 B.n282 585
R780 B.n284 B.n193 585
R781 B.n286 B.n285 585
R782 B.n287 B.n192 585
R783 B.n289 B.n288 585
R784 B.n290 B.n191 585
R785 B.n292 B.n291 585
R786 B.n293 B.n190 585
R787 B.n295 B.n294 585
R788 B.n296 B.n189 585
R789 B.n298 B.n297 585
R790 B.n299 B.n188 585
R791 B.n301 B.n300 585
R792 B.n302 B.n187 585
R793 B.n304 B.n303 585
R794 B.n305 B.n186 585
R795 B.n307 B.n306 585
R796 B.n308 B.n185 585
R797 B.n310 B.n309 585
R798 B.n311 B.n184 585
R799 B.n313 B.n312 585
R800 B.n312 B.n183 468.476
R801 B.n430 B.n429 468.476
R802 B.n632 B.n77 468.476
R803 B.n746 B.n35 468.476
R804 B.n166 B.t9 280.534
R805 B.n376 B.t0 280.534
R806 B.n58 B.t3 280.534
R807 B.n52 B.t6 280.534
R808 B.n845 B.n844 256.663
R809 B.n844 B.n843 235.042
R810 B.n844 B.n2 235.042
R811 B.n376 B.t1 173.493
R812 B.n58 B.t5 173.493
R813 B.n166 B.t10 173.482
R814 B.n52 B.t8 173.482
R815 B.n316 B.n183 163.367
R816 B.n317 B.n316 163.367
R817 B.n318 B.n317 163.367
R818 B.n318 B.n181 163.367
R819 B.n322 B.n181 163.367
R820 B.n323 B.n322 163.367
R821 B.n324 B.n323 163.367
R822 B.n324 B.n179 163.367
R823 B.n328 B.n179 163.367
R824 B.n329 B.n328 163.367
R825 B.n330 B.n329 163.367
R826 B.n330 B.n177 163.367
R827 B.n334 B.n177 163.367
R828 B.n335 B.n334 163.367
R829 B.n336 B.n335 163.367
R830 B.n336 B.n175 163.367
R831 B.n340 B.n175 163.367
R832 B.n341 B.n340 163.367
R833 B.n342 B.n341 163.367
R834 B.n342 B.n173 163.367
R835 B.n346 B.n173 163.367
R836 B.n347 B.n346 163.367
R837 B.n348 B.n347 163.367
R838 B.n348 B.n171 163.367
R839 B.n352 B.n171 163.367
R840 B.n353 B.n352 163.367
R841 B.n354 B.n353 163.367
R842 B.n354 B.n169 163.367
R843 B.n358 B.n169 163.367
R844 B.n359 B.n358 163.367
R845 B.n360 B.n359 163.367
R846 B.n360 B.n165 163.367
R847 B.n365 B.n165 163.367
R848 B.n366 B.n365 163.367
R849 B.n367 B.n366 163.367
R850 B.n367 B.n163 163.367
R851 B.n371 B.n163 163.367
R852 B.n372 B.n371 163.367
R853 B.n373 B.n372 163.367
R854 B.n373 B.n161 163.367
R855 B.n380 B.n161 163.367
R856 B.n381 B.n380 163.367
R857 B.n382 B.n381 163.367
R858 B.n382 B.n159 163.367
R859 B.n386 B.n159 163.367
R860 B.n387 B.n386 163.367
R861 B.n388 B.n387 163.367
R862 B.n388 B.n157 163.367
R863 B.n392 B.n157 163.367
R864 B.n393 B.n392 163.367
R865 B.n394 B.n393 163.367
R866 B.n394 B.n155 163.367
R867 B.n398 B.n155 163.367
R868 B.n399 B.n398 163.367
R869 B.n400 B.n399 163.367
R870 B.n400 B.n153 163.367
R871 B.n404 B.n153 163.367
R872 B.n405 B.n404 163.367
R873 B.n406 B.n405 163.367
R874 B.n406 B.n151 163.367
R875 B.n410 B.n151 163.367
R876 B.n411 B.n410 163.367
R877 B.n412 B.n411 163.367
R878 B.n412 B.n149 163.367
R879 B.n416 B.n149 163.367
R880 B.n417 B.n416 163.367
R881 B.n418 B.n417 163.367
R882 B.n418 B.n147 163.367
R883 B.n422 B.n147 163.367
R884 B.n423 B.n422 163.367
R885 B.n424 B.n423 163.367
R886 B.n424 B.n145 163.367
R887 B.n428 B.n145 163.367
R888 B.n429 B.n428 163.367
R889 B.n628 B.n77 163.367
R890 B.n628 B.n627 163.367
R891 B.n627 B.n626 163.367
R892 B.n626 B.n79 163.367
R893 B.n622 B.n79 163.367
R894 B.n622 B.n621 163.367
R895 B.n621 B.n620 163.367
R896 B.n620 B.n81 163.367
R897 B.n616 B.n81 163.367
R898 B.n616 B.n615 163.367
R899 B.n615 B.n614 163.367
R900 B.n614 B.n83 163.367
R901 B.n610 B.n83 163.367
R902 B.n610 B.n609 163.367
R903 B.n609 B.n608 163.367
R904 B.n608 B.n85 163.367
R905 B.n604 B.n85 163.367
R906 B.n604 B.n603 163.367
R907 B.n603 B.n602 163.367
R908 B.n602 B.n87 163.367
R909 B.n598 B.n87 163.367
R910 B.n598 B.n597 163.367
R911 B.n597 B.n596 163.367
R912 B.n596 B.n89 163.367
R913 B.n592 B.n89 163.367
R914 B.n592 B.n591 163.367
R915 B.n591 B.n590 163.367
R916 B.n590 B.n91 163.367
R917 B.n586 B.n91 163.367
R918 B.n586 B.n585 163.367
R919 B.n585 B.n584 163.367
R920 B.n584 B.n93 163.367
R921 B.n580 B.n93 163.367
R922 B.n580 B.n579 163.367
R923 B.n579 B.n578 163.367
R924 B.n578 B.n95 163.367
R925 B.n574 B.n95 163.367
R926 B.n574 B.n573 163.367
R927 B.n573 B.n572 163.367
R928 B.n572 B.n97 163.367
R929 B.n568 B.n97 163.367
R930 B.n568 B.n567 163.367
R931 B.n567 B.n566 163.367
R932 B.n566 B.n99 163.367
R933 B.n562 B.n99 163.367
R934 B.n562 B.n561 163.367
R935 B.n561 B.n560 163.367
R936 B.n560 B.n101 163.367
R937 B.n556 B.n101 163.367
R938 B.n556 B.n555 163.367
R939 B.n555 B.n554 163.367
R940 B.n554 B.n103 163.367
R941 B.n550 B.n103 163.367
R942 B.n550 B.n549 163.367
R943 B.n549 B.n548 163.367
R944 B.n548 B.n105 163.367
R945 B.n544 B.n105 163.367
R946 B.n544 B.n543 163.367
R947 B.n543 B.n542 163.367
R948 B.n542 B.n107 163.367
R949 B.n538 B.n107 163.367
R950 B.n538 B.n537 163.367
R951 B.n537 B.n536 163.367
R952 B.n536 B.n109 163.367
R953 B.n532 B.n109 163.367
R954 B.n532 B.n531 163.367
R955 B.n531 B.n530 163.367
R956 B.n530 B.n111 163.367
R957 B.n526 B.n111 163.367
R958 B.n526 B.n525 163.367
R959 B.n525 B.n524 163.367
R960 B.n524 B.n113 163.367
R961 B.n520 B.n113 163.367
R962 B.n520 B.n519 163.367
R963 B.n519 B.n518 163.367
R964 B.n518 B.n115 163.367
R965 B.n514 B.n115 163.367
R966 B.n514 B.n513 163.367
R967 B.n513 B.n512 163.367
R968 B.n512 B.n117 163.367
R969 B.n508 B.n117 163.367
R970 B.n508 B.n507 163.367
R971 B.n507 B.n506 163.367
R972 B.n506 B.n119 163.367
R973 B.n502 B.n119 163.367
R974 B.n502 B.n501 163.367
R975 B.n501 B.n500 163.367
R976 B.n500 B.n121 163.367
R977 B.n496 B.n121 163.367
R978 B.n496 B.n495 163.367
R979 B.n495 B.n494 163.367
R980 B.n494 B.n123 163.367
R981 B.n490 B.n123 163.367
R982 B.n490 B.n489 163.367
R983 B.n489 B.n488 163.367
R984 B.n488 B.n125 163.367
R985 B.n484 B.n125 163.367
R986 B.n484 B.n483 163.367
R987 B.n483 B.n482 163.367
R988 B.n482 B.n127 163.367
R989 B.n478 B.n127 163.367
R990 B.n478 B.n477 163.367
R991 B.n477 B.n476 163.367
R992 B.n476 B.n129 163.367
R993 B.n472 B.n129 163.367
R994 B.n472 B.n471 163.367
R995 B.n471 B.n470 163.367
R996 B.n470 B.n131 163.367
R997 B.n466 B.n131 163.367
R998 B.n466 B.n465 163.367
R999 B.n465 B.n464 163.367
R1000 B.n464 B.n133 163.367
R1001 B.n460 B.n133 163.367
R1002 B.n460 B.n459 163.367
R1003 B.n459 B.n458 163.367
R1004 B.n458 B.n135 163.367
R1005 B.n454 B.n135 163.367
R1006 B.n454 B.n453 163.367
R1007 B.n453 B.n452 163.367
R1008 B.n452 B.n137 163.367
R1009 B.n448 B.n137 163.367
R1010 B.n448 B.n447 163.367
R1011 B.n447 B.n446 163.367
R1012 B.n446 B.n139 163.367
R1013 B.n442 B.n139 163.367
R1014 B.n442 B.n441 163.367
R1015 B.n441 B.n440 163.367
R1016 B.n440 B.n141 163.367
R1017 B.n436 B.n141 163.367
R1018 B.n436 B.n435 163.367
R1019 B.n435 B.n434 163.367
R1020 B.n434 B.n143 163.367
R1021 B.n430 B.n143 163.367
R1022 B.n742 B.n35 163.367
R1023 B.n742 B.n741 163.367
R1024 B.n741 B.n740 163.367
R1025 B.n740 B.n37 163.367
R1026 B.n736 B.n37 163.367
R1027 B.n736 B.n735 163.367
R1028 B.n735 B.n734 163.367
R1029 B.n734 B.n39 163.367
R1030 B.n730 B.n39 163.367
R1031 B.n730 B.n729 163.367
R1032 B.n729 B.n728 163.367
R1033 B.n728 B.n41 163.367
R1034 B.n724 B.n41 163.367
R1035 B.n724 B.n723 163.367
R1036 B.n723 B.n722 163.367
R1037 B.n722 B.n43 163.367
R1038 B.n718 B.n43 163.367
R1039 B.n718 B.n717 163.367
R1040 B.n717 B.n716 163.367
R1041 B.n716 B.n45 163.367
R1042 B.n712 B.n45 163.367
R1043 B.n712 B.n711 163.367
R1044 B.n711 B.n710 163.367
R1045 B.n710 B.n47 163.367
R1046 B.n706 B.n47 163.367
R1047 B.n706 B.n705 163.367
R1048 B.n705 B.n704 163.367
R1049 B.n704 B.n49 163.367
R1050 B.n700 B.n49 163.367
R1051 B.n700 B.n699 163.367
R1052 B.n699 B.n698 163.367
R1053 B.n698 B.n51 163.367
R1054 B.n693 B.n51 163.367
R1055 B.n693 B.n692 163.367
R1056 B.n692 B.n691 163.367
R1057 B.n691 B.n55 163.367
R1058 B.n687 B.n55 163.367
R1059 B.n687 B.n686 163.367
R1060 B.n686 B.n685 163.367
R1061 B.n685 B.n57 163.367
R1062 B.n681 B.n57 163.367
R1063 B.n681 B.n680 163.367
R1064 B.n680 B.n61 163.367
R1065 B.n676 B.n61 163.367
R1066 B.n676 B.n675 163.367
R1067 B.n675 B.n674 163.367
R1068 B.n674 B.n63 163.367
R1069 B.n670 B.n63 163.367
R1070 B.n670 B.n669 163.367
R1071 B.n669 B.n668 163.367
R1072 B.n668 B.n65 163.367
R1073 B.n664 B.n65 163.367
R1074 B.n664 B.n663 163.367
R1075 B.n663 B.n662 163.367
R1076 B.n662 B.n67 163.367
R1077 B.n658 B.n67 163.367
R1078 B.n658 B.n657 163.367
R1079 B.n657 B.n656 163.367
R1080 B.n656 B.n69 163.367
R1081 B.n652 B.n69 163.367
R1082 B.n652 B.n651 163.367
R1083 B.n651 B.n650 163.367
R1084 B.n650 B.n71 163.367
R1085 B.n646 B.n71 163.367
R1086 B.n646 B.n645 163.367
R1087 B.n645 B.n644 163.367
R1088 B.n644 B.n73 163.367
R1089 B.n640 B.n73 163.367
R1090 B.n640 B.n639 163.367
R1091 B.n639 B.n638 163.367
R1092 B.n638 B.n75 163.367
R1093 B.n634 B.n75 163.367
R1094 B.n634 B.n633 163.367
R1095 B.n633 B.n632 163.367
R1096 B.n747 B.n746 163.367
R1097 B.n748 B.n747 163.367
R1098 B.n748 B.n33 163.367
R1099 B.n752 B.n33 163.367
R1100 B.n753 B.n752 163.367
R1101 B.n754 B.n753 163.367
R1102 B.n754 B.n31 163.367
R1103 B.n758 B.n31 163.367
R1104 B.n759 B.n758 163.367
R1105 B.n760 B.n759 163.367
R1106 B.n760 B.n29 163.367
R1107 B.n764 B.n29 163.367
R1108 B.n765 B.n764 163.367
R1109 B.n766 B.n765 163.367
R1110 B.n766 B.n27 163.367
R1111 B.n770 B.n27 163.367
R1112 B.n771 B.n770 163.367
R1113 B.n772 B.n771 163.367
R1114 B.n772 B.n25 163.367
R1115 B.n776 B.n25 163.367
R1116 B.n777 B.n776 163.367
R1117 B.n778 B.n777 163.367
R1118 B.n778 B.n23 163.367
R1119 B.n782 B.n23 163.367
R1120 B.n783 B.n782 163.367
R1121 B.n784 B.n783 163.367
R1122 B.n784 B.n21 163.367
R1123 B.n788 B.n21 163.367
R1124 B.n789 B.n788 163.367
R1125 B.n790 B.n789 163.367
R1126 B.n790 B.n19 163.367
R1127 B.n794 B.n19 163.367
R1128 B.n795 B.n794 163.367
R1129 B.n796 B.n795 163.367
R1130 B.n796 B.n17 163.367
R1131 B.n800 B.n17 163.367
R1132 B.n801 B.n800 163.367
R1133 B.n802 B.n801 163.367
R1134 B.n802 B.n15 163.367
R1135 B.n806 B.n15 163.367
R1136 B.n807 B.n806 163.367
R1137 B.n808 B.n807 163.367
R1138 B.n808 B.n13 163.367
R1139 B.n812 B.n13 163.367
R1140 B.n813 B.n812 163.367
R1141 B.n814 B.n813 163.367
R1142 B.n814 B.n11 163.367
R1143 B.n818 B.n11 163.367
R1144 B.n819 B.n818 163.367
R1145 B.n820 B.n819 163.367
R1146 B.n820 B.n9 163.367
R1147 B.n824 B.n9 163.367
R1148 B.n825 B.n824 163.367
R1149 B.n826 B.n825 163.367
R1150 B.n826 B.n7 163.367
R1151 B.n830 B.n7 163.367
R1152 B.n831 B.n830 163.367
R1153 B.n832 B.n831 163.367
R1154 B.n832 B.n5 163.367
R1155 B.n836 B.n5 163.367
R1156 B.n837 B.n836 163.367
R1157 B.n838 B.n837 163.367
R1158 B.n838 B.n3 163.367
R1159 B.n842 B.n3 163.367
R1160 B.n843 B.n842 163.367
R1161 B.n216 B.n2 163.367
R1162 B.n216 B.n215 163.367
R1163 B.n220 B.n215 163.367
R1164 B.n221 B.n220 163.367
R1165 B.n222 B.n221 163.367
R1166 B.n222 B.n213 163.367
R1167 B.n226 B.n213 163.367
R1168 B.n227 B.n226 163.367
R1169 B.n228 B.n227 163.367
R1170 B.n228 B.n211 163.367
R1171 B.n232 B.n211 163.367
R1172 B.n233 B.n232 163.367
R1173 B.n234 B.n233 163.367
R1174 B.n234 B.n209 163.367
R1175 B.n238 B.n209 163.367
R1176 B.n239 B.n238 163.367
R1177 B.n240 B.n239 163.367
R1178 B.n240 B.n207 163.367
R1179 B.n244 B.n207 163.367
R1180 B.n245 B.n244 163.367
R1181 B.n246 B.n245 163.367
R1182 B.n246 B.n205 163.367
R1183 B.n250 B.n205 163.367
R1184 B.n251 B.n250 163.367
R1185 B.n252 B.n251 163.367
R1186 B.n252 B.n203 163.367
R1187 B.n256 B.n203 163.367
R1188 B.n257 B.n256 163.367
R1189 B.n258 B.n257 163.367
R1190 B.n258 B.n201 163.367
R1191 B.n262 B.n201 163.367
R1192 B.n263 B.n262 163.367
R1193 B.n264 B.n263 163.367
R1194 B.n264 B.n199 163.367
R1195 B.n268 B.n199 163.367
R1196 B.n269 B.n268 163.367
R1197 B.n270 B.n269 163.367
R1198 B.n270 B.n197 163.367
R1199 B.n274 B.n197 163.367
R1200 B.n275 B.n274 163.367
R1201 B.n276 B.n275 163.367
R1202 B.n276 B.n195 163.367
R1203 B.n280 B.n195 163.367
R1204 B.n281 B.n280 163.367
R1205 B.n282 B.n281 163.367
R1206 B.n282 B.n193 163.367
R1207 B.n286 B.n193 163.367
R1208 B.n287 B.n286 163.367
R1209 B.n288 B.n287 163.367
R1210 B.n288 B.n191 163.367
R1211 B.n292 B.n191 163.367
R1212 B.n293 B.n292 163.367
R1213 B.n294 B.n293 163.367
R1214 B.n294 B.n189 163.367
R1215 B.n298 B.n189 163.367
R1216 B.n299 B.n298 163.367
R1217 B.n300 B.n299 163.367
R1218 B.n300 B.n187 163.367
R1219 B.n304 B.n187 163.367
R1220 B.n305 B.n304 163.367
R1221 B.n306 B.n305 163.367
R1222 B.n306 B.n185 163.367
R1223 B.n310 B.n185 163.367
R1224 B.n311 B.n310 163.367
R1225 B.n312 B.n311 163.367
R1226 B.n377 B.t2 109.299
R1227 B.n59 B.t4 109.299
R1228 B.n167 B.t11 109.288
R1229 B.n53 B.t7 109.288
R1230 B.n167 B.n166 64.1944
R1231 B.n377 B.n376 64.1944
R1232 B.n59 B.n58 64.1944
R1233 B.n53 B.n52 64.1944
R1234 B.n363 B.n167 59.5399
R1235 B.n378 B.n377 59.5399
R1236 B.n60 B.n59 59.5399
R1237 B.n695 B.n53 59.5399
R1238 B.n431 B.n144 30.4395
R1239 B.n745 B.n744 30.4395
R1240 B.n631 B.n630 30.4395
R1241 B.n314 B.n313 30.4395
R1242 B B.n845 18.0485
R1243 B.n745 B.n34 10.6151
R1244 B.n749 B.n34 10.6151
R1245 B.n750 B.n749 10.6151
R1246 B.n751 B.n750 10.6151
R1247 B.n751 B.n32 10.6151
R1248 B.n755 B.n32 10.6151
R1249 B.n756 B.n755 10.6151
R1250 B.n757 B.n756 10.6151
R1251 B.n757 B.n30 10.6151
R1252 B.n761 B.n30 10.6151
R1253 B.n762 B.n761 10.6151
R1254 B.n763 B.n762 10.6151
R1255 B.n763 B.n28 10.6151
R1256 B.n767 B.n28 10.6151
R1257 B.n768 B.n767 10.6151
R1258 B.n769 B.n768 10.6151
R1259 B.n769 B.n26 10.6151
R1260 B.n773 B.n26 10.6151
R1261 B.n774 B.n773 10.6151
R1262 B.n775 B.n774 10.6151
R1263 B.n775 B.n24 10.6151
R1264 B.n779 B.n24 10.6151
R1265 B.n780 B.n779 10.6151
R1266 B.n781 B.n780 10.6151
R1267 B.n781 B.n22 10.6151
R1268 B.n785 B.n22 10.6151
R1269 B.n786 B.n785 10.6151
R1270 B.n787 B.n786 10.6151
R1271 B.n787 B.n20 10.6151
R1272 B.n791 B.n20 10.6151
R1273 B.n792 B.n791 10.6151
R1274 B.n793 B.n792 10.6151
R1275 B.n793 B.n18 10.6151
R1276 B.n797 B.n18 10.6151
R1277 B.n798 B.n797 10.6151
R1278 B.n799 B.n798 10.6151
R1279 B.n799 B.n16 10.6151
R1280 B.n803 B.n16 10.6151
R1281 B.n804 B.n803 10.6151
R1282 B.n805 B.n804 10.6151
R1283 B.n805 B.n14 10.6151
R1284 B.n809 B.n14 10.6151
R1285 B.n810 B.n809 10.6151
R1286 B.n811 B.n810 10.6151
R1287 B.n811 B.n12 10.6151
R1288 B.n815 B.n12 10.6151
R1289 B.n816 B.n815 10.6151
R1290 B.n817 B.n816 10.6151
R1291 B.n817 B.n10 10.6151
R1292 B.n821 B.n10 10.6151
R1293 B.n822 B.n821 10.6151
R1294 B.n823 B.n822 10.6151
R1295 B.n823 B.n8 10.6151
R1296 B.n827 B.n8 10.6151
R1297 B.n828 B.n827 10.6151
R1298 B.n829 B.n828 10.6151
R1299 B.n829 B.n6 10.6151
R1300 B.n833 B.n6 10.6151
R1301 B.n834 B.n833 10.6151
R1302 B.n835 B.n834 10.6151
R1303 B.n835 B.n4 10.6151
R1304 B.n839 B.n4 10.6151
R1305 B.n840 B.n839 10.6151
R1306 B.n841 B.n840 10.6151
R1307 B.n841 B.n0 10.6151
R1308 B.n744 B.n743 10.6151
R1309 B.n743 B.n36 10.6151
R1310 B.n739 B.n36 10.6151
R1311 B.n739 B.n738 10.6151
R1312 B.n738 B.n737 10.6151
R1313 B.n737 B.n38 10.6151
R1314 B.n733 B.n38 10.6151
R1315 B.n733 B.n732 10.6151
R1316 B.n732 B.n731 10.6151
R1317 B.n731 B.n40 10.6151
R1318 B.n727 B.n40 10.6151
R1319 B.n727 B.n726 10.6151
R1320 B.n726 B.n725 10.6151
R1321 B.n725 B.n42 10.6151
R1322 B.n721 B.n42 10.6151
R1323 B.n721 B.n720 10.6151
R1324 B.n720 B.n719 10.6151
R1325 B.n719 B.n44 10.6151
R1326 B.n715 B.n44 10.6151
R1327 B.n715 B.n714 10.6151
R1328 B.n714 B.n713 10.6151
R1329 B.n713 B.n46 10.6151
R1330 B.n709 B.n46 10.6151
R1331 B.n709 B.n708 10.6151
R1332 B.n708 B.n707 10.6151
R1333 B.n707 B.n48 10.6151
R1334 B.n703 B.n48 10.6151
R1335 B.n703 B.n702 10.6151
R1336 B.n702 B.n701 10.6151
R1337 B.n701 B.n50 10.6151
R1338 B.n697 B.n50 10.6151
R1339 B.n697 B.n696 10.6151
R1340 B.n694 B.n54 10.6151
R1341 B.n690 B.n54 10.6151
R1342 B.n690 B.n689 10.6151
R1343 B.n689 B.n688 10.6151
R1344 B.n688 B.n56 10.6151
R1345 B.n684 B.n56 10.6151
R1346 B.n684 B.n683 10.6151
R1347 B.n683 B.n682 10.6151
R1348 B.n679 B.n678 10.6151
R1349 B.n678 B.n677 10.6151
R1350 B.n677 B.n62 10.6151
R1351 B.n673 B.n62 10.6151
R1352 B.n673 B.n672 10.6151
R1353 B.n672 B.n671 10.6151
R1354 B.n671 B.n64 10.6151
R1355 B.n667 B.n64 10.6151
R1356 B.n667 B.n666 10.6151
R1357 B.n666 B.n665 10.6151
R1358 B.n665 B.n66 10.6151
R1359 B.n661 B.n66 10.6151
R1360 B.n661 B.n660 10.6151
R1361 B.n660 B.n659 10.6151
R1362 B.n659 B.n68 10.6151
R1363 B.n655 B.n68 10.6151
R1364 B.n655 B.n654 10.6151
R1365 B.n654 B.n653 10.6151
R1366 B.n653 B.n70 10.6151
R1367 B.n649 B.n70 10.6151
R1368 B.n649 B.n648 10.6151
R1369 B.n648 B.n647 10.6151
R1370 B.n647 B.n72 10.6151
R1371 B.n643 B.n72 10.6151
R1372 B.n643 B.n642 10.6151
R1373 B.n642 B.n641 10.6151
R1374 B.n641 B.n74 10.6151
R1375 B.n637 B.n74 10.6151
R1376 B.n637 B.n636 10.6151
R1377 B.n636 B.n635 10.6151
R1378 B.n635 B.n76 10.6151
R1379 B.n631 B.n76 10.6151
R1380 B.n630 B.n629 10.6151
R1381 B.n629 B.n78 10.6151
R1382 B.n625 B.n78 10.6151
R1383 B.n625 B.n624 10.6151
R1384 B.n624 B.n623 10.6151
R1385 B.n623 B.n80 10.6151
R1386 B.n619 B.n80 10.6151
R1387 B.n619 B.n618 10.6151
R1388 B.n618 B.n617 10.6151
R1389 B.n617 B.n82 10.6151
R1390 B.n613 B.n82 10.6151
R1391 B.n613 B.n612 10.6151
R1392 B.n612 B.n611 10.6151
R1393 B.n611 B.n84 10.6151
R1394 B.n607 B.n84 10.6151
R1395 B.n607 B.n606 10.6151
R1396 B.n606 B.n605 10.6151
R1397 B.n605 B.n86 10.6151
R1398 B.n601 B.n86 10.6151
R1399 B.n601 B.n600 10.6151
R1400 B.n600 B.n599 10.6151
R1401 B.n599 B.n88 10.6151
R1402 B.n595 B.n88 10.6151
R1403 B.n595 B.n594 10.6151
R1404 B.n594 B.n593 10.6151
R1405 B.n593 B.n90 10.6151
R1406 B.n589 B.n90 10.6151
R1407 B.n589 B.n588 10.6151
R1408 B.n588 B.n587 10.6151
R1409 B.n587 B.n92 10.6151
R1410 B.n583 B.n92 10.6151
R1411 B.n583 B.n582 10.6151
R1412 B.n582 B.n581 10.6151
R1413 B.n581 B.n94 10.6151
R1414 B.n577 B.n94 10.6151
R1415 B.n577 B.n576 10.6151
R1416 B.n576 B.n575 10.6151
R1417 B.n575 B.n96 10.6151
R1418 B.n571 B.n96 10.6151
R1419 B.n571 B.n570 10.6151
R1420 B.n570 B.n569 10.6151
R1421 B.n569 B.n98 10.6151
R1422 B.n565 B.n98 10.6151
R1423 B.n565 B.n564 10.6151
R1424 B.n564 B.n563 10.6151
R1425 B.n563 B.n100 10.6151
R1426 B.n559 B.n100 10.6151
R1427 B.n559 B.n558 10.6151
R1428 B.n558 B.n557 10.6151
R1429 B.n557 B.n102 10.6151
R1430 B.n553 B.n102 10.6151
R1431 B.n553 B.n552 10.6151
R1432 B.n552 B.n551 10.6151
R1433 B.n551 B.n104 10.6151
R1434 B.n547 B.n104 10.6151
R1435 B.n547 B.n546 10.6151
R1436 B.n546 B.n545 10.6151
R1437 B.n545 B.n106 10.6151
R1438 B.n541 B.n106 10.6151
R1439 B.n541 B.n540 10.6151
R1440 B.n540 B.n539 10.6151
R1441 B.n539 B.n108 10.6151
R1442 B.n535 B.n108 10.6151
R1443 B.n535 B.n534 10.6151
R1444 B.n534 B.n533 10.6151
R1445 B.n533 B.n110 10.6151
R1446 B.n529 B.n110 10.6151
R1447 B.n529 B.n528 10.6151
R1448 B.n528 B.n527 10.6151
R1449 B.n527 B.n112 10.6151
R1450 B.n523 B.n112 10.6151
R1451 B.n523 B.n522 10.6151
R1452 B.n522 B.n521 10.6151
R1453 B.n521 B.n114 10.6151
R1454 B.n517 B.n114 10.6151
R1455 B.n517 B.n516 10.6151
R1456 B.n516 B.n515 10.6151
R1457 B.n515 B.n116 10.6151
R1458 B.n511 B.n116 10.6151
R1459 B.n511 B.n510 10.6151
R1460 B.n510 B.n509 10.6151
R1461 B.n509 B.n118 10.6151
R1462 B.n505 B.n118 10.6151
R1463 B.n505 B.n504 10.6151
R1464 B.n504 B.n503 10.6151
R1465 B.n503 B.n120 10.6151
R1466 B.n499 B.n120 10.6151
R1467 B.n499 B.n498 10.6151
R1468 B.n498 B.n497 10.6151
R1469 B.n497 B.n122 10.6151
R1470 B.n493 B.n122 10.6151
R1471 B.n493 B.n492 10.6151
R1472 B.n492 B.n491 10.6151
R1473 B.n491 B.n124 10.6151
R1474 B.n487 B.n124 10.6151
R1475 B.n487 B.n486 10.6151
R1476 B.n486 B.n485 10.6151
R1477 B.n485 B.n126 10.6151
R1478 B.n481 B.n126 10.6151
R1479 B.n481 B.n480 10.6151
R1480 B.n480 B.n479 10.6151
R1481 B.n479 B.n128 10.6151
R1482 B.n475 B.n128 10.6151
R1483 B.n475 B.n474 10.6151
R1484 B.n474 B.n473 10.6151
R1485 B.n473 B.n130 10.6151
R1486 B.n469 B.n130 10.6151
R1487 B.n469 B.n468 10.6151
R1488 B.n468 B.n467 10.6151
R1489 B.n467 B.n132 10.6151
R1490 B.n463 B.n132 10.6151
R1491 B.n463 B.n462 10.6151
R1492 B.n462 B.n461 10.6151
R1493 B.n461 B.n134 10.6151
R1494 B.n457 B.n134 10.6151
R1495 B.n457 B.n456 10.6151
R1496 B.n456 B.n455 10.6151
R1497 B.n455 B.n136 10.6151
R1498 B.n451 B.n136 10.6151
R1499 B.n451 B.n450 10.6151
R1500 B.n450 B.n449 10.6151
R1501 B.n449 B.n138 10.6151
R1502 B.n445 B.n138 10.6151
R1503 B.n445 B.n444 10.6151
R1504 B.n444 B.n443 10.6151
R1505 B.n443 B.n140 10.6151
R1506 B.n439 B.n140 10.6151
R1507 B.n439 B.n438 10.6151
R1508 B.n438 B.n437 10.6151
R1509 B.n437 B.n142 10.6151
R1510 B.n433 B.n142 10.6151
R1511 B.n433 B.n432 10.6151
R1512 B.n432 B.n431 10.6151
R1513 B.n217 B.n1 10.6151
R1514 B.n218 B.n217 10.6151
R1515 B.n219 B.n218 10.6151
R1516 B.n219 B.n214 10.6151
R1517 B.n223 B.n214 10.6151
R1518 B.n224 B.n223 10.6151
R1519 B.n225 B.n224 10.6151
R1520 B.n225 B.n212 10.6151
R1521 B.n229 B.n212 10.6151
R1522 B.n230 B.n229 10.6151
R1523 B.n231 B.n230 10.6151
R1524 B.n231 B.n210 10.6151
R1525 B.n235 B.n210 10.6151
R1526 B.n236 B.n235 10.6151
R1527 B.n237 B.n236 10.6151
R1528 B.n237 B.n208 10.6151
R1529 B.n241 B.n208 10.6151
R1530 B.n242 B.n241 10.6151
R1531 B.n243 B.n242 10.6151
R1532 B.n243 B.n206 10.6151
R1533 B.n247 B.n206 10.6151
R1534 B.n248 B.n247 10.6151
R1535 B.n249 B.n248 10.6151
R1536 B.n249 B.n204 10.6151
R1537 B.n253 B.n204 10.6151
R1538 B.n254 B.n253 10.6151
R1539 B.n255 B.n254 10.6151
R1540 B.n255 B.n202 10.6151
R1541 B.n259 B.n202 10.6151
R1542 B.n260 B.n259 10.6151
R1543 B.n261 B.n260 10.6151
R1544 B.n261 B.n200 10.6151
R1545 B.n265 B.n200 10.6151
R1546 B.n266 B.n265 10.6151
R1547 B.n267 B.n266 10.6151
R1548 B.n267 B.n198 10.6151
R1549 B.n271 B.n198 10.6151
R1550 B.n272 B.n271 10.6151
R1551 B.n273 B.n272 10.6151
R1552 B.n273 B.n196 10.6151
R1553 B.n277 B.n196 10.6151
R1554 B.n278 B.n277 10.6151
R1555 B.n279 B.n278 10.6151
R1556 B.n279 B.n194 10.6151
R1557 B.n283 B.n194 10.6151
R1558 B.n284 B.n283 10.6151
R1559 B.n285 B.n284 10.6151
R1560 B.n285 B.n192 10.6151
R1561 B.n289 B.n192 10.6151
R1562 B.n290 B.n289 10.6151
R1563 B.n291 B.n290 10.6151
R1564 B.n291 B.n190 10.6151
R1565 B.n295 B.n190 10.6151
R1566 B.n296 B.n295 10.6151
R1567 B.n297 B.n296 10.6151
R1568 B.n297 B.n188 10.6151
R1569 B.n301 B.n188 10.6151
R1570 B.n302 B.n301 10.6151
R1571 B.n303 B.n302 10.6151
R1572 B.n303 B.n186 10.6151
R1573 B.n307 B.n186 10.6151
R1574 B.n308 B.n307 10.6151
R1575 B.n309 B.n308 10.6151
R1576 B.n309 B.n184 10.6151
R1577 B.n313 B.n184 10.6151
R1578 B.n315 B.n314 10.6151
R1579 B.n315 B.n182 10.6151
R1580 B.n319 B.n182 10.6151
R1581 B.n320 B.n319 10.6151
R1582 B.n321 B.n320 10.6151
R1583 B.n321 B.n180 10.6151
R1584 B.n325 B.n180 10.6151
R1585 B.n326 B.n325 10.6151
R1586 B.n327 B.n326 10.6151
R1587 B.n327 B.n178 10.6151
R1588 B.n331 B.n178 10.6151
R1589 B.n332 B.n331 10.6151
R1590 B.n333 B.n332 10.6151
R1591 B.n333 B.n176 10.6151
R1592 B.n337 B.n176 10.6151
R1593 B.n338 B.n337 10.6151
R1594 B.n339 B.n338 10.6151
R1595 B.n339 B.n174 10.6151
R1596 B.n343 B.n174 10.6151
R1597 B.n344 B.n343 10.6151
R1598 B.n345 B.n344 10.6151
R1599 B.n345 B.n172 10.6151
R1600 B.n349 B.n172 10.6151
R1601 B.n350 B.n349 10.6151
R1602 B.n351 B.n350 10.6151
R1603 B.n351 B.n170 10.6151
R1604 B.n355 B.n170 10.6151
R1605 B.n356 B.n355 10.6151
R1606 B.n357 B.n356 10.6151
R1607 B.n357 B.n168 10.6151
R1608 B.n361 B.n168 10.6151
R1609 B.n362 B.n361 10.6151
R1610 B.n364 B.n164 10.6151
R1611 B.n368 B.n164 10.6151
R1612 B.n369 B.n368 10.6151
R1613 B.n370 B.n369 10.6151
R1614 B.n370 B.n162 10.6151
R1615 B.n374 B.n162 10.6151
R1616 B.n375 B.n374 10.6151
R1617 B.n379 B.n375 10.6151
R1618 B.n383 B.n160 10.6151
R1619 B.n384 B.n383 10.6151
R1620 B.n385 B.n384 10.6151
R1621 B.n385 B.n158 10.6151
R1622 B.n389 B.n158 10.6151
R1623 B.n390 B.n389 10.6151
R1624 B.n391 B.n390 10.6151
R1625 B.n391 B.n156 10.6151
R1626 B.n395 B.n156 10.6151
R1627 B.n396 B.n395 10.6151
R1628 B.n397 B.n396 10.6151
R1629 B.n397 B.n154 10.6151
R1630 B.n401 B.n154 10.6151
R1631 B.n402 B.n401 10.6151
R1632 B.n403 B.n402 10.6151
R1633 B.n403 B.n152 10.6151
R1634 B.n407 B.n152 10.6151
R1635 B.n408 B.n407 10.6151
R1636 B.n409 B.n408 10.6151
R1637 B.n409 B.n150 10.6151
R1638 B.n413 B.n150 10.6151
R1639 B.n414 B.n413 10.6151
R1640 B.n415 B.n414 10.6151
R1641 B.n415 B.n148 10.6151
R1642 B.n419 B.n148 10.6151
R1643 B.n420 B.n419 10.6151
R1644 B.n421 B.n420 10.6151
R1645 B.n421 B.n146 10.6151
R1646 B.n425 B.n146 10.6151
R1647 B.n426 B.n425 10.6151
R1648 B.n427 B.n426 10.6151
R1649 B.n427 B.n144 10.6151
R1650 B.n845 B.n0 8.11757
R1651 B.n845 B.n1 8.11757
R1652 B.n695 B.n694 6.5566
R1653 B.n682 B.n60 6.5566
R1654 B.n364 B.n363 6.5566
R1655 B.n379 B.n378 6.5566
R1656 B.n696 B.n695 4.05904
R1657 B.n679 B.n60 4.05904
R1658 B.n363 B.n362 4.05904
R1659 B.n378 B.n160 4.05904
C0 w_n4942_n2748# VTAIL 2.83858f
C1 VDD2 VTAIL 9.23178f
C2 B VP 2.42548f
C3 VN VP 8.39608f
C4 w_n4942_n2748# VP 11.293599f
C5 VDD1 B 2.38191f
C6 VDD2 VP 0.631534f
C7 VDD1 VN 0.153929f
C8 VDD1 w_n4942_n2748# 2.72029f
C9 VDD1 VDD2 2.42178f
C10 B VN 1.33946f
C11 w_n4942_n2748# B 10.3169f
C12 w_n4942_n2748# VN 10.649f
C13 VDD2 B 2.51463f
C14 VTAIL VP 9.21278f
C15 VDD2 VN 8.25064f
C16 w_n4942_n2748# VDD2 2.88359f
C17 VDD1 VTAIL 9.17728f
C18 VDD1 VP 8.72486f
C19 VTAIL B 3.17193f
C20 VTAIL VN 9.198559f
C21 VDD2 VSUBS 2.261767f
C22 VDD1 VSUBS 2.041982f
C23 VTAIL VSUBS 1.29775f
C24 VN VSUBS 8.26688f
C25 VP VSUBS 4.621844f
C26 B VSUBS 5.577731f
C27 w_n4942_n2748# VSUBS 0.168127p
C28 B.n0 VSUBS 0.008989f
C29 B.n1 VSUBS 0.008989f
C30 B.n2 VSUBS 0.013295f
C31 B.n3 VSUBS 0.010188f
C32 B.n4 VSUBS 0.010188f
C33 B.n5 VSUBS 0.010188f
C34 B.n6 VSUBS 0.010188f
C35 B.n7 VSUBS 0.010188f
C36 B.n8 VSUBS 0.010188f
C37 B.n9 VSUBS 0.010188f
C38 B.n10 VSUBS 0.010188f
C39 B.n11 VSUBS 0.010188f
C40 B.n12 VSUBS 0.010188f
C41 B.n13 VSUBS 0.010188f
C42 B.n14 VSUBS 0.010188f
C43 B.n15 VSUBS 0.010188f
C44 B.n16 VSUBS 0.010188f
C45 B.n17 VSUBS 0.010188f
C46 B.n18 VSUBS 0.010188f
C47 B.n19 VSUBS 0.010188f
C48 B.n20 VSUBS 0.010188f
C49 B.n21 VSUBS 0.010188f
C50 B.n22 VSUBS 0.010188f
C51 B.n23 VSUBS 0.010188f
C52 B.n24 VSUBS 0.010188f
C53 B.n25 VSUBS 0.010188f
C54 B.n26 VSUBS 0.010188f
C55 B.n27 VSUBS 0.010188f
C56 B.n28 VSUBS 0.010188f
C57 B.n29 VSUBS 0.010188f
C58 B.n30 VSUBS 0.010188f
C59 B.n31 VSUBS 0.010188f
C60 B.n32 VSUBS 0.010188f
C61 B.n33 VSUBS 0.010188f
C62 B.n34 VSUBS 0.010188f
C63 B.n35 VSUBS 0.023639f
C64 B.n36 VSUBS 0.010188f
C65 B.n37 VSUBS 0.010188f
C66 B.n38 VSUBS 0.010188f
C67 B.n39 VSUBS 0.010188f
C68 B.n40 VSUBS 0.010188f
C69 B.n41 VSUBS 0.010188f
C70 B.n42 VSUBS 0.010188f
C71 B.n43 VSUBS 0.010188f
C72 B.n44 VSUBS 0.010188f
C73 B.n45 VSUBS 0.010188f
C74 B.n46 VSUBS 0.010188f
C75 B.n47 VSUBS 0.010188f
C76 B.n48 VSUBS 0.010188f
C77 B.n49 VSUBS 0.010188f
C78 B.n50 VSUBS 0.010188f
C79 B.n51 VSUBS 0.010188f
C80 B.t7 VSUBS 0.406469f
C81 B.t8 VSUBS 0.440445f
C82 B.t6 VSUBS 1.80358f
C83 B.n52 VSUBS 0.240473f
C84 B.n53 VSUBS 0.10635f
C85 B.n54 VSUBS 0.010188f
C86 B.n55 VSUBS 0.010188f
C87 B.n56 VSUBS 0.010188f
C88 B.n57 VSUBS 0.010188f
C89 B.t4 VSUBS 0.406464f
C90 B.t5 VSUBS 0.44044f
C91 B.t3 VSUBS 1.80358f
C92 B.n58 VSUBS 0.240477f
C93 B.n59 VSUBS 0.106355f
C94 B.n60 VSUBS 0.023604f
C95 B.n61 VSUBS 0.010188f
C96 B.n62 VSUBS 0.010188f
C97 B.n63 VSUBS 0.010188f
C98 B.n64 VSUBS 0.010188f
C99 B.n65 VSUBS 0.010188f
C100 B.n66 VSUBS 0.010188f
C101 B.n67 VSUBS 0.010188f
C102 B.n68 VSUBS 0.010188f
C103 B.n69 VSUBS 0.010188f
C104 B.n70 VSUBS 0.010188f
C105 B.n71 VSUBS 0.010188f
C106 B.n72 VSUBS 0.010188f
C107 B.n73 VSUBS 0.010188f
C108 B.n74 VSUBS 0.010188f
C109 B.n75 VSUBS 0.010188f
C110 B.n76 VSUBS 0.010188f
C111 B.n77 VSUBS 0.021907f
C112 B.n78 VSUBS 0.010188f
C113 B.n79 VSUBS 0.010188f
C114 B.n80 VSUBS 0.010188f
C115 B.n81 VSUBS 0.010188f
C116 B.n82 VSUBS 0.010188f
C117 B.n83 VSUBS 0.010188f
C118 B.n84 VSUBS 0.010188f
C119 B.n85 VSUBS 0.010188f
C120 B.n86 VSUBS 0.010188f
C121 B.n87 VSUBS 0.010188f
C122 B.n88 VSUBS 0.010188f
C123 B.n89 VSUBS 0.010188f
C124 B.n90 VSUBS 0.010188f
C125 B.n91 VSUBS 0.010188f
C126 B.n92 VSUBS 0.010188f
C127 B.n93 VSUBS 0.010188f
C128 B.n94 VSUBS 0.010188f
C129 B.n95 VSUBS 0.010188f
C130 B.n96 VSUBS 0.010188f
C131 B.n97 VSUBS 0.010188f
C132 B.n98 VSUBS 0.010188f
C133 B.n99 VSUBS 0.010188f
C134 B.n100 VSUBS 0.010188f
C135 B.n101 VSUBS 0.010188f
C136 B.n102 VSUBS 0.010188f
C137 B.n103 VSUBS 0.010188f
C138 B.n104 VSUBS 0.010188f
C139 B.n105 VSUBS 0.010188f
C140 B.n106 VSUBS 0.010188f
C141 B.n107 VSUBS 0.010188f
C142 B.n108 VSUBS 0.010188f
C143 B.n109 VSUBS 0.010188f
C144 B.n110 VSUBS 0.010188f
C145 B.n111 VSUBS 0.010188f
C146 B.n112 VSUBS 0.010188f
C147 B.n113 VSUBS 0.010188f
C148 B.n114 VSUBS 0.010188f
C149 B.n115 VSUBS 0.010188f
C150 B.n116 VSUBS 0.010188f
C151 B.n117 VSUBS 0.010188f
C152 B.n118 VSUBS 0.010188f
C153 B.n119 VSUBS 0.010188f
C154 B.n120 VSUBS 0.010188f
C155 B.n121 VSUBS 0.010188f
C156 B.n122 VSUBS 0.010188f
C157 B.n123 VSUBS 0.010188f
C158 B.n124 VSUBS 0.010188f
C159 B.n125 VSUBS 0.010188f
C160 B.n126 VSUBS 0.010188f
C161 B.n127 VSUBS 0.010188f
C162 B.n128 VSUBS 0.010188f
C163 B.n129 VSUBS 0.010188f
C164 B.n130 VSUBS 0.010188f
C165 B.n131 VSUBS 0.010188f
C166 B.n132 VSUBS 0.010188f
C167 B.n133 VSUBS 0.010188f
C168 B.n134 VSUBS 0.010188f
C169 B.n135 VSUBS 0.010188f
C170 B.n136 VSUBS 0.010188f
C171 B.n137 VSUBS 0.010188f
C172 B.n138 VSUBS 0.010188f
C173 B.n139 VSUBS 0.010188f
C174 B.n140 VSUBS 0.010188f
C175 B.n141 VSUBS 0.010188f
C176 B.n142 VSUBS 0.010188f
C177 B.n143 VSUBS 0.010188f
C178 B.n144 VSUBS 0.022348f
C179 B.n145 VSUBS 0.010188f
C180 B.n146 VSUBS 0.010188f
C181 B.n147 VSUBS 0.010188f
C182 B.n148 VSUBS 0.010188f
C183 B.n149 VSUBS 0.010188f
C184 B.n150 VSUBS 0.010188f
C185 B.n151 VSUBS 0.010188f
C186 B.n152 VSUBS 0.010188f
C187 B.n153 VSUBS 0.010188f
C188 B.n154 VSUBS 0.010188f
C189 B.n155 VSUBS 0.010188f
C190 B.n156 VSUBS 0.010188f
C191 B.n157 VSUBS 0.010188f
C192 B.n158 VSUBS 0.010188f
C193 B.n159 VSUBS 0.010188f
C194 B.n160 VSUBS 0.007042f
C195 B.n161 VSUBS 0.010188f
C196 B.n162 VSUBS 0.010188f
C197 B.n163 VSUBS 0.010188f
C198 B.n164 VSUBS 0.010188f
C199 B.n165 VSUBS 0.010188f
C200 B.t11 VSUBS 0.406469f
C201 B.t10 VSUBS 0.440445f
C202 B.t9 VSUBS 1.80358f
C203 B.n166 VSUBS 0.240473f
C204 B.n167 VSUBS 0.10635f
C205 B.n168 VSUBS 0.010188f
C206 B.n169 VSUBS 0.010188f
C207 B.n170 VSUBS 0.010188f
C208 B.n171 VSUBS 0.010188f
C209 B.n172 VSUBS 0.010188f
C210 B.n173 VSUBS 0.010188f
C211 B.n174 VSUBS 0.010188f
C212 B.n175 VSUBS 0.010188f
C213 B.n176 VSUBS 0.010188f
C214 B.n177 VSUBS 0.010188f
C215 B.n178 VSUBS 0.010188f
C216 B.n179 VSUBS 0.010188f
C217 B.n180 VSUBS 0.010188f
C218 B.n181 VSUBS 0.010188f
C219 B.n182 VSUBS 0.010188f
C220 B.n183 VSUBS 0.023639f
C221 B.n184 VSUBS 0.010188f
C222 B.n185 VSUBS 0.010188f
C223 B.n186 VSUBS 0.010188f
C224 B.n187 VSUBS 0.010188f
C225 B.n188 VSUBS 0.010188f
C226 B.n189 VSUBS 0.010188f
C227 B.n190 VSUBS 0.010188f
C228 B.n191 VSUBS 0.010188f
C229 B.n192 VSUBS 0.010188f
C230 B.n193 VSUBS 0.010188f
C231 B.n194 VSUBS 0.010188f
C232 B.n195 VSUBS 0.010188f
C233 B.n196 VSUBS 0.010188f
C234 B.n197 VSUBS 0.010188f
C235 B.n198 VSUBS 0.010188f
C236 B.n199 VSUBS 0.010188f
C237 B.n200 VSUBS 0.010188f
C238 B.n201 VSUBS 0.010188f
C239 B.n202 VSUBS 0.010188f
C240 B.n203 VSUBS 0.010188f
C241 B.n204 VSUBS 0.010188f
C242 B.n205 VSUBS 0.010188f
C243 B.n206 VSUBS 0.010188f
C244 B.n207 VSUBS 0.010188f
C245 B.n208 VSUBS 0.010188f
C246 B.n209 VSUBS 0.010188f
C247 B.n210 VSUBS 0.010188f
C248 B.n211 VSUBS 0.010188f
C249 B.n212 VSUBS 0.010188f
C250 B.n213 VSUBS 0.010188f
C251 B.n214 VSUBS 0.010188f
C252 B.n215 VSUBS 0.010188f
C253 B.n216 VSUBS 0.010188f
C254 B.n217 VSUBS 0.010188f
C255 B.n218 VSUBS 0.010188f
C256 B.n219 VSUBS 0.010188f
C257 B.n220 VSUBS 0.010188f
C258 B.n221 VSUBS 0.010188f
C259 B.n222 VSUBS 0.010188f
C260 B.n223 VSUBS 0.010188f
C261 B.n224 VSUBS 0.010188f
C262 B.n225 VSUBS 0.010188f
C263 B.n226 VSUBS 0.010188f
C264 B.n227 VSUBS 0.010188f
C265 B.n228 VSUBS 0.010188f
C266 B.n229 VSUBS 0.010188f
C267 B.n230 VSUBS 0.010188f
C268 B.n231 VSUBS 0.010188f
C269 B.n232 VSUBS 0.010188f
C270 B.n233 VSUBS 0.010188f
C271 B.n234 VSUBS 0.010188f
C272 B.n235 VSUBS 0.010188f
C273 B.n236 VSUBS 0.010188f
C274 B.n237 VSUBS 0.010188f
C275 B.n238 VSUBS 0.010188f
C276 B.n239 VSUBS 0.010188f
C277 B.n240 VSUBS 0.010188f
C278 B.n241 VSUBS 0.010188f
C279 B.n242 VSUBS 0.010188f
C280 B.n243 VSUBS 0.010188f
C281 B.n244 VSUBS 0.010188f
C282 B.n245 VSUBS 0.010188f
C283 B.n246 VSUBS 0.010188f
C284 B.n247 VSUBS 0.010188f
C285 B.n248 VSUBS 0.010188f
C286 B.n249 VSUBS 0.010188f
C287 B.n250 VSUBS 0.010188f
C288 B.n251 VSUBS 0.010188f
C289 B.n252 VSUBS 0.010188f
C290 B.n253 VSUBS 0.010188f
C291 B.n254 VSUBS 0.010188f
C292 B.n255 VSUBS 0.010188f
C293 B.n256 VSUBS 0.010188f
C294 B.n257 VSUBS 0.010188f
C295 B.n258 VSUBS 0.010188f
C296 B.n259 VSUBS 0.010188f
C297 B.n260 VSUBS 0.010188f
C298 B.n261 VSUBS 0.010188f
C299 B.n262 VSUBS 0.010188f
C300 B.n263 VSUBS 0.010188f
C301 B.n264 VSUBS 0.010188f
C302 B.n265 VSUBS 0.010188f
C303 B.n266 VSUBS 0.010188f
C304 B.n267 VSUBS 0.010188f
C305 B.n268 VSUBS 0.010188f
C306 B.n269 VSUBS 0.010188f
C307 B.n270 VSUBS 0.010188f
C308 B.n271 VSUBS 0.010188f
C309 B.n272 VSUBS 0.010188f
C310 B.n273 VSUBS 0.010188f
C311 B.n274 VSUBS 0.010188f
C312 B.n275 VSUBS 0.010188f
C313 B.n276 VSUBS 0.010188f
C314 B.n277 VSUBS 0.010188f
C315 B.n278 VSUBS 0.010188f
C316 B.n279 VSUBS 0.010188f
C317 B.n280 VSUBS 0.010188f
C318 B.n281 VSUBS 0.010188f
C319 B.n282 VSUBS 0.010188f
C320 B.n283 VSUBS 0.010188f
C321 B.n284 VSUBS 0.010188f
C322 B.n285 VSUBS 0.010188f
C323 B.n286 VSUBS 0.010188f
C324 B.n287 VSUBS 0.010188f
C325 B.n288 VSUBS 0.010188f
C326 B.n289 VSUBS 0.010188f
C327 B.n290 VSUBS 0.010188f
C328 B.n291 VSUBS 0.010188f
C329 B.n292 VSUBS 0.010188f
C330 B.n293 VSUBS 0.010188f
C331 B.n294 VSUBS 0.010188f
C332 B.n295 VSUBS 0.010188f
C333 B.n296 VSUBS 0.010188f
C334 B.n297 VSUBS 0.010188f
C335 B.n298 VSUBS 0.010188f
C336 B.n299 VSUBS 0.010188f
C337 B.n300 VSUBS 0.010188f
C338 B.n301 VSUBS 0.010188f
C339 B.n302 VSUBS 0.010188f
C340 B.n303 VSUBS 0.010188f
C341 B.n304 VSUBS 0.010188f
C342 B.n305 VSUBS 0.010188f
C343 B.n306 VSUBS 0.010188f
C344 B.n307 VSUBS 0.010188f
C345 B.n308 VSUBS 0.010188f
C346 B.n309 VSUBS 0.010188f
C347 B.n310 VSUBS 0.010188f
C348 B.n311 VSUBS 0.010188f
C349 B.n312 VSUBS 0.021907f
C350 B.n313 VSUBS 0.021907f
C351 B.n314 VSUBS 0.023639f
C352 B.n315 VSUBS 0.010188f
C353 B.n316 VSUBS 0.010188f
C354 B.n317 VSUBS 0.010188f
C355 B.n318 VSUBS 0.010188f
C356 B.n319 VSUBS 0.010188f
C357 B.n320 VSUBS 0.010188f
C358 B.n321 VSUBS 0.010188f
C359 B.n322 VSUBS 0.010188f
C360 B.n323 VSUBS 0.010188f
C361 B.n324 VSUBS 0.010188f
C362 B.n325 VSUBS 0.010188f
C363 B.n326 VSUBS 0.010188f
C364 B.n327 VSUBS 0.010188f
C365 B.n328 VSUBS 0.010188f
C366 B.n329 VSUBS 0.010188f
C367 B.n330 VSUBS 0.010188f
C368 B.n331 VSUBS 0.010188f
C369 B.n332 VSUBS 0.010188f
C370 B.n333 VSUBS 0.010188f
C371 B.n334 VSUBS 0.010188f
C372 B.n335 VSUBS 0.010188f
C373 B.n336 VSUBS 0.010188f
C374 B.n337 VSUBS 0.010188f
C375 B.n338 VSUBS 0.010188f
C376 B.n339 VSUBS 0.010188f
C377 B.n340 VSUBS 0.010188f
C378 B.n341 VSUBS 0.010188f
C379 B.n342 VSUBS 0.010188f
C380 B.n343 VSUBS 0.010188f
C381 B.n344 VSUBS 0.010188f
C382 B.n345 VSUBS 0.010188f
C383 B.n346 VSUBS 0.010188f
C384 B.n347 VSUBS 0.010188f
C385 B.n348 VSUBS 0.010188f
C386 B.n349 VSUBS 0.010188f
C387 B.n350 VSUBS 0.010188f
C388 B.n351 VSUBS 0.010188f
C389 B.n352 VSUBS 0.010188f
C390 B.n353 VSUBS 0.010188f
C391 B.n354 VSUBS 0.010188f
C392 B.n355 VSUBS 0.010188f
C393 B.n356 VSUBS 0.010188f
C394 B.n357 VSUBS 0.010188f
C395 B.n358 VSUBS 0.010188f
C396 B.n359 VSUBS 0.010188f
C397 B.n360 VSUBS 0.010188f
C398 B.n361 VSUBS 0.010188f
C399 B.n362 VSUBS 0.007042f
C400 B.n363 VSUBS 0.023604f
C401 B.n364 VSUBS 0.00824f
C402 B.n365 VSUBS 0.010188f
C403 B.n366 VSUBS 0.010188f
C404 B.n367 VSUBS 0.010188f
C405 B.n368 VSUBS 0.010188f
C406 B.n369 VSUBS 0.010188f
C407 B.n370 VSUBS 0.010188f
C408 B.n371 VSUBS 0.010188f
C409 B.n372 VSUBS 0.010188f
C410 B.n373 VSUBS 0.010188f
C411 B.n374 VSUBS 0.010188f
C412 B.n375 VSUBS 0.010188f
C413 B.t2 VSUBS 0.406464f
C414 B.t1 VSUBS 0.44044f
C415 B.t0 VSUBS 1.80358f
C416 B.n376 VSUBS 0.240477f
C417 B.n377 VSUBS 0.106355f
C418 B.n378 VSUBS 0.023604f
C419 B.n379 VSUBS 0.00824f
C420 B.n380 VSUBS 0.010188f
C421 B.n381 VSUBS 0.010188f
C422 B.n382 VSUBS 0.010188f
C423 B.n383 VSUBS 0.010188f
C424 B.n384 VSUBS 0.010188f
C425 B.n385 VSUBS 0.010188f
C426 B.n386 VSUBS 0.010188f
C427 B.n387 VSUBS 0.010188f
C428 B.n388 VSUBS 0.010188f
C429 B.n389 VSUBS 0.010188f
C430 B.n390 VSUBS 0.010188f
C431 B.n391 VSUBS 0.010188f
C432 B.n392 VSUBS 0.010188f
C433 B.n393 VSUBS 0.010188f
C434 B.n394 VSUBS 0.010188f
C435 B.n395 VSUBS 0.010188f
C436 B.n396 VSUBS 0.010188f
C437 B.n397 VSUBS 0.010188f
C438 B.n398 VSUBS 0.010188f
C439 B.n399 VSUBS 0.010188f
C440 B.n400 VSUBS 0.010188f
C441 B.n401 VSUBS 0.010188f
C442 B.n402 VSUBS 0.010188f
C443 B.n403 VSUBS 0.010188f
C444 B.n404 VSUBS 0.010188f
C445 B.n405 VSUBS 0.010188f
C446 B.n406 VSUBS 0.010188f
C447 B.n407 VSUBS 0.010188f
C448 B.n408 VSUBS 0.010188f
C449 B.n409 VSUBS 0.010188f
C450 B.n410 VSUBS 0.010188f
C451 B.n411 VSUBS 0.010188f
C452 B.n412 VSUBS 0.010188f
C453 B.n413 VSUBS 0.010188f
C454 B.n414 VSUBS 0.010188f
C455 B.n415 VSUBS 0.010188f
C456 B.n416 VSUBS 0.010188f
C457 B.n417 VSUBS 0.010188f
C458 B.n418 VSUBS 0.010188f
C459 B.n419 VSUBS 0.010188f
C460 B.n420 VSUBS 0.010188f
C461 B.n421 VSUBS 0.010188f
C462 B.n422 VSUBS 0.010188f
C463 B.n423 VSUBS 0.010188f
C464 B.n424 VSUBS 0.010188f
C465 B.n425 VSUBS 0.010188f
C466 B.n426 VSUBS 0.010188f
C467 B.n427 VSUBS 0.010188f
C468 B.n428 VSUBS 0.010188f
C469 B.n429 VSUBS 0.023639f
C470 B.n430 VSUBS 0.021907f
C471 B.n431 VSUBS 0.023198f
C472 B.n432 VSUBS 0.010188f
C473 B.n433 VSUBS 0.010188f
C474 B.n434 VSUBS 0.010188f
C475 B.n435 VSUBS 0.010188f
C476 B.n436 VSUBS 0.010188f
C477 B.n437 VSUBS 0.010188f
C478 B.n438 VSUBS 0.010188f
C479 B.n439 VSUBS 0.010188f
C480 B.n440 VSUBS 0.010188f
C481 B.n441 VSUBS 0.010188f
C482 B.n442 VSUBS 0.010188f
C483 B.n443 VSUBS 0.010188f
C484 B.n444 VSUBS 0.010188f
C485 B.n445 VSUBS 0.010188f
C486 B.n446 VSUBS 0.010188f
C487 B.n447 VSUBS 0.010188f
C488 B.n448 VSUBS 0.010188f
C489 B.n449 VSUBS 0.010188f
C490 B.n450 VSUBS 0.010188f
C491 B.n451 VSUBS 0.010188f
C492 B.n452 VSUBS 0.010188f
C493 B.n453 VSUBS 0.010188f
C494 B.n454 VSUBS 0.010188f
C495 B.n455 VSUBS 0.010188f
C496 B.n456 VSUBS 0.010188f
C497 B.n457 VSUBS 0.010188f
C498 B.n458 VSUBS 0.010188f
C499 B.n459 VSUBS 0.010188f
C500 B.n460 VSUBS 0.010188f
C501 B.n461 VSUBS 0.010188f
C502 B.n462 VSUBS 0.010188f
C503 B.n463 VSUBS 0.010188f
C504 B.n464 VSUBS 0.010188f
C505 B.n465 VSUBS 0.010188f
C506 B.n466 VSUBS 0.010188f
C507 B.n467 VSUBS 0.010188f
C508 B.n468 VSUBS 0.010188f
C509 B.n469 VSUBS 0.010188f
C510 B.n470 VSUBS 0.010188f
C511 B.n471 VSUBS 0.010188f
C512 B.n472 VSUBS 0.010188f
C513 B.n473 VSUBS 0.010188f
C514 B.n474 VSUBS 0.010188f
C515 B.n475 VSUBS 0.010188f
C516 B.n476 VSUBS 0.010188f
C517 B.n477 VSUBS 0.010188f
C518 B.n478 VSUBS 0.010188f
C519 B.n479 VSUBS 0.010188f
C520 B.n480 VSUBS 0.010188f
C521 B.n481 VSUBS 0.010188f
C522 B.n482 VSUBS 0.010188f
C523 B.n483 VSUBS 0.010188f
C524 B.n484 VSUBS 0.010188f
C525 B.n485 VSUBS 0.010188f
C526 B.n486 VSUBS 0.010188f
C527 B.n487 VSUBS 0.010188f
C528 B.n488 VSUBS 0.010188f
C529 B.n489 VSUBS 0.010188f
C530 B.n490 VSUBS 0.010188f
C531 B.n491 VSUBS 0.010188f
C532 B.n492 VSUBS 0.010188f
C533 B.n493 VSUBS 0.010188f
C534 B.n494 VSUBS 0.010188f
C535 B.n495 VSUBS 0.010188f
C536 B.n496 VSUBS 0.010188f
C537 B.n497 VSUBS 0.010188f
C538 B.n498 VSUBS 0.010188f
C539 B.n499 VSUBS 0.010188f
C540 B.n500 VSUBS 0.010188f
C541 B.n501 VSUBS 0.010188f
C542 B.n502 VSUBS 0.010188f
C543 B.n503 VSUBS 0.010188f
C544 B.n504 VSUBS 0.010188f
C545 B.n505 VSUBS 0.010188f
C546 B.n506 VSUBS 0.010188f
C547 B.n507 VSUBS 0.010188f
C548 B.n508 VSUBS 0.010188f
C549 B.n509 VSUBS 0.010188f
C550 B.n510 VSUBS 0.010188f
C551 B.n511 VSUBS 0.010188f
C552 B.n512 VSUBS 0.010188f
C553 B.n513 VSUBS 0.010188f
C554 B.n514 VSUBS 0.010188f
C555 B.n515 VSUBS 0.010188f
C556 B.n516 VSUBS 0.010188f
C557 B.n517 VSUBS 0.010188f
C558 B.n518 VSUBS 0.010188f
C559 B.n519 VSUBS 0.010188f
C560 B.n520 VSUBS 0.010188f
C561 B.n521 VSUBS 0.010188f
C562 B.n522 VSUBS 0.010188f
C563 B.n523 VSUBS 0.010188f
C564 B.n524 VSUBS 0.010188f
C565 B.n525 VSUBS 0.010188f
C566 B.n526 VSUBS 0.010188f
C567 B.n527 VSUBS 0.010188f
C568 B.n528 VSUBS 0.010188f
C569 B.n529 VSUBS 0.010188f
C570 B.n530 VSUBS 0.010188f
C571 B.n531 VSUBS 0.010188f
C572 B.n532 VSUBS 0.010188f
C573 B.n533 VSUBS 0.010188f
C574 B.n534 VSUBS 0.010188f
C575 B.n535 VSUBS 0.010188f
C576 B.n536 VSUBS 0.010188f
C577 B.n537 VSUBS 0.010188f
C578 B.n538 VSUBS 0.010188f
C579 B.n539 VSUBS 0.010188f
C580 B.n540 VSUBS 0.010188f
C581 B.n541 VSUBS 0.010188f
C582 B.n542 VSUBS 0.010188f
C583 B.n543 VSUBS 0.010188f
C584 B.n544 VSUBS 0.010188f
C585 B.n545 VSUBS 0.010188f
C586 B.n546 VSUBS 0.010188f
C587 B.n547 VSUBS 0.010188f
C588 B.n548 VSUBS 0.010188f
C589 B.n549 VSUBS 0.010188f
C590 B.n550 VSUBS 0.010188f
C591 B.n551 VSUBS 0.010188f
C592 B.n552 VSUBS 0.010188f
C593 B.n553 VSUBS 0.010188f
C594 B.n554 VSUBS 0.010188f
C595 B.n555 VSUBS 0.010188f
C596 B.n556 VSUBS 0.010188f
C597 B.n557 VSUBS 0.010188f
C598 B.n558 VSUBS 0.010188f
C599 B.n559 VSUBS 0.010188f
C600 B.n560 VSUBS 0.010188f
C601 B.n561 VSUBS 0.010188f
C602 B.n562 VSUBS 0.010188f
C603 B.n563 VSUBS 0.010188f
C604 B.n564 VSUBS 0.010188f
C605 B.n565 VSUBS 0.010188f
C606 B.n566 VSUBS 0.010188f
C607 B.n567 VSUBS 0.010188f
C608 B.n568 VSUBS 0.010188f
C609 B.n569 VSUBS 0.010188f
C610 B.n570 VSUBS 0.010188f
C611 B.n571 VSUBS 0.010188f
C612 B.n572 VSUBS 0.010188f
C613 B.n573 VSUBS 0.010188f
C614 B.n574 VSUBS 0.010188f
C615 B.n575 VSUBS 0.010188f
C616 B.n576 VSUBS 0.010188f
C617 B.n577 VSUBS 0.010188f
C618 B.n578 VSUBS 0.010188f
C619 B.n579 VSUBS 0.010188f
C620 B.n580 VSUBS 0.010188f
C621 B.n581 VSUBS 0.010188f
C622 B.n582 VSUBS 0.010188f
C623 B.n583 VSUBS 0.010188f
C624 B.n584 VSUBS 0.010188f
C625 B.n585 VSUBS 0.010188f
C626 B.n586 VSUBS 0.010188f
C627 B.n587 VSUBS 0.010188f
C628 B.n588 VSUBS 0.010188f
C629 B.n589 VSUBS 0.010188f
C630 B.n590 VSUBS 0.010188f
C631 B.n591 VSUBS 0.010188f
C632 B.n592 VSUBS 0.010188f
C633 B.n593 VSUBS 0.010188f
C634 B.n594 VSUBS 0.010188f
C635 B.n595 VSUBS 0.010188f
C636 B.n596 VSUBS 0.010188f
C637 B.n597 VSUBS 0.010188f
C638 B.n598 VSUBS 0.010188f
C639 B.n599 VSUBS 0.010188f
C640 B.n600 VSUBS 0.010188f
C641 B.n601 VSUBS 0.010188f
C642 B.n602 VSUBS 0.010188f
C643 B.n603 VSUBS 0.010188f
C644 B.n604 VSUBS 0.010188f
C645 B.n605 VSUBS 0.010188f
C646 B.n606 VSUBS 0.010188f
C647 B.n607 VSUBS 0.010188f
C648 B.n608 VSUBS 0.010188f
C649 B.n609 VSUBS 0.010188f
C650 B.n610 VSUBS 0.010188f
C651 B.n611 VSUBS 0.010188f
C652 B.n612 VSUBS 0.010188f
C653 B.n613 VSUBS 0.010188f
C654 B.n614 VSUBS 0.010188f
C655 B.n615 VSUBS 0.010188f
C656 B.n616 VSUBS 0.010188f
C657 B.n617 VSUBS 0.010188f
C658 B.n618 VSUBS 0.010188f
C659 B.n619 VSUBS 0.010188f
C660 B.n620 VSUBS 0.010188f
C661 B.n621 VSUBS 0.010188f
C662 B.n622 VSUBS 0.010188f
C663 B.n623 VSUBS 0.010188f
C664 B.n624 VSUBS 0.010188f
C665 B.n625 VSUBS 0.010188f
C666 B.n626 VSUBS 0.010188f
C667 B.n627 VSUBS 0.010188f
C668 B.n628 VSUBS 0.010188f
C669 B.n629 VSUBS 0.010188f
C670 B.n630 VSUBS 0.021907f
C671 B.n631 VSUBS 0.023639f
C672 B.n632 VSUBS 0.023639f
C673 B.n633 VSUBS 0.010188f
C674 B.n634 VSUBS 0.010188f
C675 B.n635 VSUBS 0.010188f
C676 B.n636 VSUBS 0.010188f
C677 B.n637 VSUBS 0.010188f
C678 B.n638 VSUBS 0.010188f
C679 B.n639 VSUBS 0.010188f
C680 B.n640 VSUBS 0.010188f
C681 B.n641 VSUBS 0.010188f
C682 B.n642 VSUBS 0.010188f
C683 B.n643 VSUBS 0.010188f
C684 B.n644 VSUBS 0.010188f
C685 B.n645 VSUBS 0.010188f
C686 B.n646 VSUBS 0.010188f
C687 B.n647 VSUBS 0.010188f
C688 B.n648 VSUBS 0.010188f
C689 B.n649 VSUBS 0.010188f
C690 B.n650 VSUBS 0.010188f
C691 B.n651 VSUBS 0.010188f
C692 B.n652 VSUBS 0.010188f
C693 B.n653 VSUBS 0.010188f
C694 B.n654 VSUBS 0.010188f
C695 B.n655 VSUBS 0.010188f
C696 B.n656 VSUBS 0.010188f
C697 B.n657 VSUBS 0.010188f
C698 B.n658 VSUBS 0.010188f
C699 B.n659 VSUBS 0.010188f
C700 B.n660 VSUBS 0.010188f
C701 B.n661 VSUBS 0.010188f
C702 B.n662 VSUBS 0.010188f
C703 B.n663 VSUBS 0.010188f
C704 B.n664 VSUBS 0.010188f
C705 B.n665 VSUBS 0.010188f
C706 B.n666 VSUBS 0.010188f
C707 B.n667 VSUBS 0.010188f
C708 B.n668 VSUBS 0.010188f
C709 B.n669 VSUBS 0.010188f
C710 B.n670 VSUBS 0.010188f
C711 B.n671 VSUBS 0.010188f
C712 B.n672 VSUBS 0.010188f
C713 B.n673 VSUBS 0.010188f
C714 B.n674 VSUBS 0.010188f
C715 B.n675 VSUBS 0.010188f
C716 B.n676 VSUBS 0.010188f
C717 B.n677 VSUBS 0.010188f
C718 B.n678 VSUBS 0.010188f
C719 B.n679 VSUBS 0.007042f
C720 B.n680 VSUBS 0.010188f
C721 B.n681 VSUBS 0.010188f
C722 B.n682 VSUBS 0.00824f
C723 B.n683 VSUBS 0.010188f
C724 B.n684 VSUBS 0.010188f
C725 B.n685 VSUBS 0.010188f
C726 B.n686 VSUBS 0.010188f
C727 B.n687 VSUBS 0.010188f
C728 B.n688 VSUBS 0.010188f
C729 B.n689 VSUBS 0.010188f
C730 B.n690 VSUBS 0.010188f
C731 B.n691 VSUBS 0.010188f
C732 B.n692 VSUBS 0.010188f
C733 B.n693 VSUBS 0.010188f
C734 B.n694 VSUBS 0.00824f
C735 B.n695 VSUBS 0.023604f
C736 B.n696 VSUBS 0.007042f
C737 B.n697 VSUBS 0.010188f
C738 B.n698 VSUBS 0.010188f
C739 B.n699 VSUBS 0.010188f
C740 B.n700 VSUBS 0.010188f
C741 B.n701 VSUBS 0.010188f
C742 B.n702 VSUBS 0.010188f
C743 B.n703 VSUBS 0.010188f
C744 B.n704 VSUBS 0.010188f
C745 B.n705 VSUBS 0.010188f
C746 B.n706 VSUBS 0.010188f
C747 B.n707 VSUBS 0.010188f
C748 B.n708 VSUBS 0.010188f
C749 B.n709 VSUBS 0.010188f
C750 B.n710 VSUBS 0.010188f
C751 B.n711 VSUBS 0.010188f
C752 B.n712 VSUBS 0.010188f
C753 B.n713 VSUBS 0.010188f
C754 B.n714 VSUBS 0.010188f
C755 B.n715 VSUBS 0.010188f
C756 B.n716 VSUBS 0.010188f
C757 B.n717 VSUBS 0.010188f
C758 B.n718 VSUBS 0.010188f
C759 B.n719 VSUBS 0.010188f
C760 B.n720 VSUBS 0.010188f
C761 B.n721 VSUBS 0.010188f
C762 B.n722 VSUBS 0.010188f
C763 B.n723 VSUBS 0.010188f
C764 B.n724 VSUBS 0.010188f
C765 B.n725 VSUBS 0.010188f
C766 B.n726 VSUBS 0.010188f
C767 B.n727 VSUBS 0.010188f
C768 B.n728 VSUBS 0.010188f
C769 B.n729 VSUBS 0.010188f
C770 B.n730 VSUBS 0.010188f
C771 B.n731 VSUBS 0.010188f
C772 B.n732 VSUBS 0.010188f
C773 B.n733 VSUBS 0.010188f
C774 B.n734 VSUBS 0.010188f
C775 B.n735 VSUBS 0.010188f
C776 B.n736 VSUBS 0.010188f
C777 B.n737 VSUBS 0.010188f
C778 B.n738 VSUBS 0.010188f
C779 B.n739 VSUBS 0.010188f
C780 B.n740 VSUBS 0.010188f
C781 B.n741 VSUBS 0.010188f
C782 B.n742 VSUBS 0.010188f
C783 B.n743 VSUBS 0.010188f
C784 B.n744 VSUBS 0.023639f
C785 B.n745 VSUBS 0.021907f
C786 B.n746 VSUBS 0.021907f
C787 B.n747 VSUBS 0.010188f
C788 B.n748 VSUBS 0.010188f
C789 B.n749 VSUBS 0.010188f
C790 B.n750 VSUBS 0.010188f
C791 B.n751 VSUBS 0.010188f
C792 B.n752 VSUBS 0.010188f
C793 B.n753 VSUBS 0.010188f
C794 B.n754 VSUBS 0.010188f
C795 B.n755 VSUBS 0.010188f
C796 B.n756 VSUBS 0.010188f
C797 B.n757 VSUBS 0.010188f
C798 B.n758 VSUBS 0.010188f
C799 B.n759 VSUBS 0.010188f
C800 B.n760 VSUBS 0.010188f
C801 B.n761 VSUBS 0.010188f
C802 B.n762 VSUBS 0.010188f
C803 B.n763 VSUBS 0.010188f
C804 B.n764 VSUBS 0.010188f
C805 B.n765 VSUBS 0.010188f
C806 B.n766 VSUBS 0.010188f
C807 B.n767 VSUBS 0.010188f
C808 B.n768 VSUBS 0.010188f
C809 B.n769 VSUBS 0.010188f
C810 B.n770 VSUBS 0.010188f
C811 B.n771 VSUBS 0.010188f
C812 B.n772 VSUBS 0.010188f
C813 B.n773 VSUBS 0.010188f
C814 B.n774 VSUBS 0.010188f
C815 B.n775 VSUBS 0.010188f
C816 B.n776 VSUBS 0.010188f
C817 B.n777 VSUBS 0.010188f
C818 B.n778 VSUBS 0.010188f
C819 B.n779 VSUBS 0.010188f
C820 B.n780 VSUBS 0.010188f
C821 B.n781 VSUBS 0.010188f
C822 B.n782 VSUBS 0.010188f
C823 B.n783 VSUBS 0.010188f
C824 B.n784 VSUBS 0.010188f
C825 B.n785 VSUBS 0.010188f
C826 B.n786 VSUBS 0.010188f
C827 B.n787 VSUBS 0.010188f
C828 B.n788 VSUBS 0.010188f
C829 B.n789 VSUBS 0.010188f
C830 B.n790 VSUBS 0.010188f
C831 B.n791 VSUBS 0.010188f
C832 B.n792 VSUBS 0.010188f
C833 B.n793 VSUBS 0.010188f
C834 B.n794 VSUBS 0.010188f
C835 B.n795 VSUBS 0.010188f
C836 B.n796 VSUBS 0.010188f
C837 B.n797 VSUBS 0.010188f
C838 B.n798 VSUBS 0.010188f
C839 B.n799 VSUBS 0.010188f
C840 B.n800 VSUBS 0.010188f
C841 B.n801 VSUBS 0.010188f
C842 B.n802 VSUBS 0.010188f
C843 B.n803 VSUBS 0.010188f
C844 B.n804 VSUBS 0.010188f
C845 B.n805 VSUBS 0.010188f
C846 B.n806 VSUBS 0.010188f
C847 B.n807 VSUBS 0.010188f
C848 B.n808 VSUBS 0.010188f
C849 B.n809 VSUBS 0.010188f
C850 B.n810 VSUBS 0.010188f
C851 B.n811 VSUBS 0.010188f
C852 B.n812 VSUBS 0.010188f
C853 B.n813 VSUBS 0.010188f
C854 B.n814 VSUBS 0.010188f
C855 B.n815 VSUBS 0.010188f
C856 B.n816 VSUBS 0.010188f
C857 B.n817 VSUBS 0.010188f
C858 B.n818 VSUBS 0.010188f
C859 B.n819 VSUBS 0.010188f
C860 B.n820 VSUBS 0.010188f
C861 B.n821 VSUBS 0.010188f
C862 B.n822 VSUBS 0.010188f
C863 B.n823 VSUBS 0.010188f
C864 B.n824 VSUBS 0.010188f
C865 B.n825 VSUBS 0.010188f
C866 B.n826 VSUBS 0.010188f
C867 B.n827 VSUBS 0.010188f
C868 B.n828 VSUBS 0.010188f
C869 B.n829 VSUBS 0.010188f
C870 B.n830 VSUBS 0.010188f
C871 B.n831 VSUBS 0.010188f
C872 B.n832 VSUBS 0.010188f
C873 B.n833 VSUBS 0.010188f
C874 B.n834 VSUBS 0.010188f
C875 B.n835 VSUBS 0.010188f
C876 B.n836 VSUBS 0.010188f
C877 B.n837 VSUBS 0.010188f
C878 B.n838 VSUBS 0.010188f
C879 B.n839 VSUBS 0.010188f
C880 B.n840 VSUBS 0.010188f
C881 B.n841 VSUBS 0.010188f
C882 B.n842 VSUBS 0.010188f
C883 B.n843 VSUBS 0.013295f
C884 B.n844 VSUBS 0.014162f
C885 B.n845 VSUBS 0.028163f
C886 VDD2.t7 VSUBS 2.2218f
C887 VDD2.t5 VSUBS 0.225512f
C888 VDD2.t9 VSUBS 0.225512f
C889 VDD2.n0 VSUBS 1.66495f
C890 VDD2.n1 VSUBS 1.85468f
C891 VDD2.t2 VSUBS 0.225512f
C892 VDD2.t8 VSUBS 0.225512f
C893 VDD2.n2 VSUBS 1.6926f
C894 VDD2.n3 VSUBS 4.03185f
C895 VDD2.t0 VSUBS 2.19006f
C896 VDD2.n4 VSUBS 4.19305f
C897 VDD2.t1 VSUBS 0.225512f
C898 VDD2.t3 VSUBS 0.225512f
C899 VDD2.n5 VSUBS 1.66495f
C900 VDD2.n6 VSUBS 0.936949f
C901 VDD2.t4 VSUBS 0.225512f
C902 VDD2.t6 VSUBS 0.225512f
C903 VDD2.n7 VSUBS 1.69254f
C904 VN.t1 VSUBS 2.07344f
C905 VN.n0 VSUBS 0.855705f
C906 VN.n1 VSUBS 0.028982f
C907 VN.n2 VSUBS 0.039646f
C908 VN.n3 VSUBS 0.028982f
C909 VN.t7 VSUBS 2.07344f
C910 VN.n4 VSUBS 0.054285f
C911 VN.n5 VSUBS 0.028982f
C912 VN.n6 VSUBS 0.054285f
C913 VN.n7 VSUBS 0.028982f
C914 VN.t0 VSUBS 2.07344f
C915 VN.n8 VSUBS 0.053739f
C916 VN.n9 VSUBS 0.028982f
C917 VN.n10 VSUBS 0.030699f
C918 VN.t4 VSUBS 2.07344f
C919 VN.n11 VSUBS 0.827601f
C920 VN.t2 VSUBS 2.35867f
C921 VN.n12 VSUBS 0.803687f
C922 VN.n13 VSUBS 0.313676f
C923 VN.n14 VSUBS 0.028982f
C924 VN.n15 VSUBS 0.054285f
C925 VN.n16 VSUBS 0.058507f
C926 VN.n17 VSUBS 0.027024f
C927 VN.n18 VSUBS 0.028982f
C928 VN.n19 VSUBS 0.028982f
C929 VN.n20 VSUBS 0.028982f
C930 VN.n21 VSUBS 0.054285f
C931 VN.n22 VSUBS 0.040884f
C932 VN.n23 VSUBS 0.744843f
C933 VN.n24 VSUBS 0.040884f
C934 VN.n25 VSUBS 0.028982f
C935 VN.n26 VSUBS 0.028982f
C936 VN.n27 VSUBS 0.028982f
C937 VN.n28 VSUBS 0.053739f
C938 VN.n29 VSUBS 0.027024f
C939 VN.n30 VSUBS 0.058507f
C940 VN.n31 VSUBS 0.028982f
C941 VN.n32 VSUBS 0.028982f
C942 VN.n33 VSUBS 0.028982f
C943 VN.n34 VSUBS 0.030699f
C944 VN.n35 VSUBS 0.744843f
C945 VN.n36 VSUBS 0.051069f
C946 VN.n37 VSUBS 0.054285f
C947 VN.n38 VSUBS 0.028982f
C948 VN.n39 VSUBS 0.028982f
C949 VN.n40 VSUBS 0.028982f
C950 VN.n41 VSUBS 0.045339f
C951 VN.n42 VSUBS 0.054285f
C952 VN.n43 VSUBS 0.047317f
C953 VN.n44 VSUBS 0.046783f
C954 VN.n45 VSUBS 0.062546f
C955 VN.t9 VSUBS 2.07344f
C956 VN.n46 VSUBS 0.855705f
C957 VN.n47 VSUBS 0.028982f
C958 VN.n48 VSUBS 0.039646f
C959 VN.n49 VSUBS 0.028982f
C960 VN.t8 VSUBS 2.07344f
C961 VN.n50 VSUBS 0.054285f
C962 VN.n51 VSUBS 0.028982f
C963 VN.n52 VSUBS 0.054285f
C964 VN.n53 VSUBS 0.028982f
C965 VN.t6 VSUBS 2.07344f
C966 VN.n54 VSUBS 0.053739f
C967 VN.n55 VSUBS 0.028982f
C968 VN.n56 VSUBS 0.030699f
C969 VN.t3 VSUBS 2.35867f
C970 VN.t5 VSUBS 2.07344f
C971 VN.n57 VSUBS 0.827601f
C972 VN.n58 VSUBS 0.803687f
C973 VN.n59 VSUBS 0.313676f
C974 VN.n60 VSUBS 0.028982f
C975 VN.n61 VSUBS 0.054285f
C976 VN.n62 VSUBS 0.058507f
C977 VN.n63 VSUBS 0.027024f
C978 VN.n64 VSUBS 0.028982f
C979 VN.n65 VSUBS 0.028982f
C980 VN.n66 VSUBS 0.028982f
C981 VN.n67 VSUBS 0.054285f
C982 VN.n68 VSUBS 0.040884f
C983 VN.n69 VSUBS 0.744843f
C984 VN.n70 VSUBS 0.040884f
C985 VN.n71 VSUBS 0.028982f
C986 VN.n72 VSUBS 0.028982f
C987 VN.n73 VSUBS 0.028982f
C988 VN.n74 VSUBS 0.053739f
C989 VN.n75 VSUBS 0.027024f
C990 VN.n76 VSUBS 0.058507f
C991 VN.n77 VSUBS 0.028982f
C992 VN.n78 VSUBS 0.028982f
C993 VN.n79 VSUBS 0.028982f
C994 VN.n80 VSUBS 0.030699f
C995 VN.n81 VSUBS 0.744843f
C996 VN.n82 VSUBS 0.051069f
C997 VN.n83 VSUBS 0.054285f
C998 VN.n84 VSUBS 0.028982f
C999 VN.n85 VSUBS 0.028982f
C1000 VN.n86 VSUBS 0.028982f
C1001 VN.n87 VSUBS 0.045339f
C1002 VN.n88 VSUBS 0.054285f
C1003 VN.n89 VSUBS 0.047317f
C1004 VN.n90 VSUBS 0.046783f
C1005 VN.n91 VSUBS 1.78942f
C1006 VTAIL.t16 VSUBS 0.217109f
C1007 VTAIL.t2 VSUBS 0.217109f
C1008 VTAIL.n0 VSUBS 1.46137f
C1009 VTAIL.n1 VSUBS 1.04835f
C1010 VTAIL.t11 VSUBS 1.95303f
C1011 VTAIL.n2 VSUBS 1.21397f
C1012 VTAIL.t12 VSUBS 0.217109f
C1013 VTAIL.t5 VSUBS 0.217109f
C1014 VTAIL.n3 VSUBS 1.46137f
C1015 VTAIL.n4 VSUBS 1.2087f
C1016 VTAIL.t4 VSUBS 0.217109f
C1017 VTAIL.t10 VSUBS 0.217109f
C1018 VTAIL.n5 VSUBS 1.46137f
C1019 VTAIL.n6 VSUBS 2.67503f
C1020 VTAIL.t17 VSUBS 0.217109f
C1021 VTAIL.t19 VSUBS 0.217109f
C1022 VTAIL.n7 VSUBS 1.46138f
C1023 VTAIL.n8 VSUBS 2.67503f
C1024 VTAIL.t18 VSUBS 0.217109f
C1025 VTAIL.t14 VSUBS 0.217109f
C1026 VTAIL.n9 VSUBS 1.46138f
C1027 VTAIL.n10 VSUBS 1.2087f
C1028 VTAIL.t3 VSUBS 1.95304f
C1029 VTAIL.n11 VSUBS 1.21397f
C1030 VTAIL.t6 VSUBS 0.217109f
C1031 VTAIL.t8 VSUBS 0.217109f
C1032 VTAIL.n12 VSUBS 1.46138f
C1033 VTAIL.n13 VSUBS 1.11352f
C1034 VTAIL.t9 VSUBS 0.217109f
C1035 VTAIL.t13 VSUBS 0.217109f
C1036 VTAIL.n14 VSUBS 1.46138f
C1037 VTAIL.n15 VSUBS 1.2087f
C1038 VTAIL.t7 VSUBS 1.95303f
C1039 VTAIL.n16 VSUBS 2.49166f
C1040 VTAIL.t0 VSUBS 1.95303f
C1041 VTAIL.n17 VSUBS 2.49166f
C1042 VTAIL.t1 VSUBS 0.217109f
C1043 VTAIL.t15 VSUBS 0.217109f
C1044 VTAIL.n18 VSUBS 1.46137f
C1045 VTAIL.n19 VSUBS 0.990042f
C1046 VDD1.t7 VSUBS 2.2202f
C1047 VDD1.t2 VSUBS 0.225348f
C1048 VDD1.t1 VSUBS 0.225348f
C1049 VDD1.n0 VSUBS 1.66374f
C1050 VDD1.n1 VSUBS 1.86392f
C1051 VDD1.t4 VSUBS 2.22019f
C1052 VDD1.t9 VSUBS 0.225348f
C1053 VDD1.t5 VSUBS 0.225348f
C1054 VDD1.n2 VSUBS 1.66374f
C1055 VDD1.n3 VSUBS 1.85334f
C1056 VDD1.t3 VSUBS 0.225348f
C1057 VDD1.t8 VSUBS 0.225348f
C1058 VDD1.n4 VSUBS 1.69137f
C1059 VDD1.n5 VSUBS 4.19927f
C1060 VDD1.t6 VSUBS 0.225348f
C1061 VDD1.t0 VSUBS 0.225348f
C1062 VDD1.n6 VSUBS 1.66374f
C1063 VDD1.n7 VSUBS 4.2631f
C1064 VP.t2 VSUBS 2.27481f
C1065 VP.n0 VSUBS 0.938806f
C1066 VP.n1 VSUBS 0.031796f
C1067 VP.n2 VSUBS 0.043496f
C1068 VP.n3 VSUBS 0.031796f
C1069 VP.t8 VSUBS 2.27481f
C1070 VP.n4 VSUBS 0.059557f
C1071 VP.n5 VSUBS 0.031796f
C1072 VP.n6 VSUBS 0.059557f
C1073 VP.n7 VSUBS 0.031796f
C1074 VP.t1 VSUBS 2.27481f
C1075 VP.n8 VSUBS 0.058958f
C1076 VP.n9 VSUBS 0.031796f
C1077 VP.n10 VSUBS 0.03368f
C1078 VP.n11 VSUBS 0.031796f
C1079 VP.n12 VSUBS 0.049742f
C1080 VP.n13 VSUBS 0.051327f
C1081 VP.t9 VSUBS 2.27481f
C1082 VP.t6 VSUBS 2.27481f
C1083 VP.n14 VSUBS 0.938806f
C1084 VP.n15 VSUBS 0.031796f
C1085 VP.n16 VSUBS 0.043496f
C1086 VP.n17 VSUBS 0.031796f
C1087 VP.t0 VSUBS 2.27481f
C1088 VP.n18 VSUBS 0.059557f
C1089 VP.n19 VSUBS 0.031796f
C1090 VP.n20 VSUBS 0.059557f
C1091 VP.n21 VSUBS 0.031796f
C1092 VP.t4 VSUBS 2.27481f
C1093 VP.n22 VSUBS 0.058958f
C1094 VP.n23 VSUBS 0.031796f
C1095 VP.n24 VSUBS 0.03368f
C1096 VP.t7 VSUBS 2.58773f
C1097 VP.t5 VSUBS 2.27481f
C1098 VP.n25 VSUBS 0.907973f
C1099 VP.n26 VSUBS 0.881738f
C1100 VP.n27 VSUBS 0.34414f
C1101 VP.n28 VSUBS 0.031796f
C1102 VP.n29 VSUBS 0.059557f
C1103 VP.n30 VSUBS 0.064189f
C1104 VP.n31 VSUBS 0.029648f
C1105 VP.n32 VSUBS 0.031796f
C1106 VP.n33 VSUBS 0.031796f
C1107 VP.n34 VSUBS 0.031796f
C1108 VP.n35 VSUBS 0.059557f
C1109 VP.n36 VSUBS 0.044854f
C1110 VP.n37 VSUBS 0.817179f
C1111 VP.n38 VSUBS 0.044854f
C1112 VP.n39 VSUBS 0.031796f
C1113 VP.n40 VSUBS 0.031796f
C1114 VP.n41 VSUBS 0.031796f
C1115 VP.n42 VSUBS 0.058958f
C1116 VP.n43 VSUBS 0.029648f
C1117 VP.n44 VSUBS 0.064189f
C1118 VP.n45 VSUBS 0.031796f
C1119 VP.n46 VSUBS 0.031796f
C1120 VP.n47 VSUBS 0.031796f
C1121 VP.n48 VSUBS 0.03368f
C1122 VP.n49 VSUBS 0.817179f
C1123 VP.n50 VSUBS 0.056028f
C1124 VP.n51 VSUBS 0.059557f
C1125 VP.n52 VSUBS 0.031796f
C1126 VP.n53 VSUBS 0.031796f
C1127 VP.n54 VSUBS 0.031796f
C1128 VP.n55 VSUBS 0.049742f
C1129 VP.n56 VSUBS 0.059557f
C1130 VP.n57 VSUBS 0.051912f
C1131 VP.n58 VSUBS 0.051327f
C1132 VP.n59 VSUBS 1.95043f
C1133 VP.n60 VSUBS 1.97196f
C1134 VP.n61 VSUBS 0.938806f
C1135 VP.n62 VSUBS 0.051912f
C1136 VP.n63 VSUBS 0.059557f
C1137 VP.n64 VSUBS 0.031796f
C1138 VP.n65 VSUBS 0.031796f
C1139 VP.n66 VSUBS 0.031796f
C1140 VP.n67 VSUBS 0.043496f
C1141 VP.n68 VSUBS 0.059557f
C1142 VP.t3 VSUBS 2.27481f
C1143 VP.n69 VSUBS 0.817179f
C1144 VP.n70 VSUBS 0.056028f
C1145 VP.n71 VSUBS 0.031796f
C1146 VP.n72 VSUBS 0.031796f
C1147 VP.n73 VSUBS 0.031796f
C1148 VP.n74 VSUBS 0.059557f
C1149 VP.n75 VSUBS 0.064189f
C1150 VP.n76 VSUBS 0.029648f
C1151 VP.n77 VSUBS 0.031796f
C1152 VP.n78 VSUBS 0.031796f
C1153 VP.n79 VSUBS 0.031796f
C1154 VP.n80 VSUBS 0.059557f
C1155 VP.n81 VSUBS 0.044854f
C1156 VP.n82 VSUBS 0.817179f
C1157 VP.n83 VSUBS 0.044854f
C1158 VP.n84 VSUBS 0.031796f
C1159 VP.n85 VSUBS 0.031796f
C1160 VP.n86 VSUBS 0.031796f
C1161 VP.n87 VSUBS 0.058958f
C1162 VP.n88 VSUBS 0.029648f
C1163 VP.n89 VSUBS 0.064189f
C1164 VP.n90 VSUBS 0.031796f
C1165 VP.n91 VSUBS 0.031796f
C1166 VP.n92 VSUBS 0.031796f
C1167 VP.n93 VSUBS 0.03368f
C1168 VP.n94 VSUBS 0.817179f
C1169 VP.n95 VSUBS 0.056028f
C1170 VP.n96 VSUBS 0.059557f
C1171 VP.n97 VSUBS 0.031796f
C1172 VP.n98 VSUBS 0.031796f
C1173 VP.n99 VSUBS 0.031796f
C1174 VP.n100 VSUBS 0.049742f
C1175 VP.n101 VSUBS 0.059557f
C1176 VP.n102 VSUBS 0.051912f
C1177 VP.n103 VSUBS 0.051327f
C1178 VP.n104 VSUBS 0.06862f
.ends

