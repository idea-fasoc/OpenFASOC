* NGSPICE file created from diff_pair_sample_0962.ext - technology: sky130A

.subckt diff_pair_sample_0962 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t1 VN.t0 VTAIL.t3 w_n2166_n4924# sky130_fd_pr__pfet_01v8 ad=7.7142 pd=40.34 as=7.7142 ps=40.34 w=19.78 l=2.66
X1 VDD1.t1 VP.t0 VTAIL.t0 w_n2166_n4924# sky130_fd_pr__pfet_01v8 ad=7.7142 pd=40.34 as=7.7142 ps=40.34 w=19.78 l=2.66
X2 VDD2.t0 VN.t1 VTAIL.t2 w_n2166_n4924# sky130_fd_pr__pfet_01v8 ad=7.7142 pd=40.34 as=7.7142 ps=40.34 w=19.78 l=2.66
X3 B.t11 B.t9 B.t10 w_n2166_n4924# sky130_fd_pr__pfet_01v8 ad=7.7142 pd=40.34 as=0 ps=0 w=19.78 l=2.66
X4 VDD1.t0 VP.t1 VTAIL.t1 w_n2166_n4924# sky130_fd_pr__pfet_01v8 ad=7.7142 pd=40.34 as=7.7142 ps=40.34 w=19.78 l=2.66
X5 B.t8 B.t6 B.t7 w_n2166_n4924# sky130_fd_pr__pfet_01v8 ad=7.7142 pd=40.34 as=0 ps=0 w=19.78 l=2.66
X6 B.t5 B.t3 B.t4 w_n2166_n4924# sky130_fd_pr__pfet_01v8 ad=7.7142 pd=40.34 as=0 ps=0 w=19.78 l=2.66
X7 B.t2 B.t0 B.t1 w_n2166_n4924# sky130_fd_pr__pfet_01v8 ad=7.7142 pd=40.34 as=0 ps=0 w=19.78 l=2.66
R0 VN VN.t1 270.976
R1 VN VN.t0 220.696
R2 VTAIL.n1 VTAIL.t2 54.6261
R3 VTAIL.n3 VTAIL.t3 54.6259
R4 VTAIL.n0 VTAIL.t1 54.6259
R5 VTAIL.n2 VTAIL.t0 54.6259
R6 VTAIL.n1 VTAIL.n0 34.5738
R7 VTAIL.n3 VTAIL.n2 31.9962
R8 VTAIL.n2 VTAIL.n1 1.75912
R9 VTAIL VTAIL.n0 1.17291
R10 VTAIL VTAIL.n3 0.586707
R11 VDD2.n0 VDD2.t1 117.171
R12 VDD2.n0 VDD2.t0 71.3047
R13 VDD2 VDD2.n0 0.703086
R14 VP.n0 VP.t0 270.974
R15 VP.n0 VP.t1 220.264
R16 VP VP.n0 0.43181
R17 VDD1 VDD1.t0 118.341
R18 VDD1 VDD1.t1 72.0073
R19 B.n445 B.n114 585
R20 B.n444 B.n443 585
R21 B.n442 B.n115 585
R22 B.n441 B.n440 585
R23 B.n439 B.n116 585
R24 B.n438 B.n437 585
R25 B.n436 B.n117 585
R26 B.n435 B.n434 585
R27 B.n433 B.n118 585
R28 B.n432 B.n431 585
R29 B.n430 B.n119 585
R30 B.n429 B.n428 585
R31 B.n427 B.n120 585
R32 B.n426 B.n425 585
R33 B.n424 B.n121 585
R34 B.n423 B.n422 585
R35 B.n421 B.n122 585
R36 B.n420 B.n419 585
R37 B.n418 B.n123 585
R38 B.n417 B.n416 585
R39 B.n415 B.n124 585
R40 B.n414 B.n413 585
R41 B.n412 B.n125 585
R42 B.n411 B.n410 585
R43 B.n409 B.n126 585
R44 B.n408 B.n407 585
R45 B.n406 B.n127 585
R46 B.n405 B.n404 585
R47 B.n403 B.n128 585
R48 B.n402 B.n401 585
R49 B.n400 B.n129 585
R50 B.n399 B.n398 585
R51 B.n397 B.n130 585
R52 B.n396 B.n395 585
R53 B.n394 B.n131 585
R54 B.n393 B.n392 585
R55 B.n391 B.n132 585
R56 B.n390 B.n389 585
R57 B.n388 B.n133 585
R58 B.n387 B.n386 585
R59 B.n385 B.n134 585
R60 B.n384 B.n383 585
R61 B.n382 B.n135 585
R62 B.n381 B.n380 585
R63 B.n379 B.n136 585
R64 B.n378 B.n377 585
R65 B.n376 B.n137 585
R66 B.n375 B.n374 585
R67 B.n373 B.n138 585
R68 B.n372 B.n371 585
R69 B.n370 B.n139 585
R70 B.n369 B.n368 585
R71 B.n367 B.n140 585
R72 B.n366 B.n365 585
R73 B.n364 B.n141 585
R74 B.n363 B.n362 585
R75 B.n361 B.n142 585
R76 B.n360 B.n359 585
R77 B.n358 B.n143 585
R78 B.n357 B.n356 585
R79 B.n355 B.n144 585
R80 B.n354 B.n353 585
R81 B.n352 B.n145 585
R82 B.n351 B.n350 585
R83 B.n349 B.n146 585
R84 B.n348 B.n347 585
R85 B.n343 B.n147 585
R86 B.n342 B.n341 585
R87 B.n340 B.n148 585
R88 B.n339 B.n338 585
R89 B.n337 B.n149 585
R90 B.n336 B.n335 585
R91 B.n334 B.n150 585
R92 B.n333 B.n332 585
R93 B.n330 B.n151 585
R94 B.n329 B.n328 585
R95 B.n327 B.n154 585
R96 B.n326 B.n325 585
R97 B.n324 B.n155 585
R98 B.n323 B.n322 585
R99 B.n321 B.n156 585
R100 B.n320 B.n319 585
R101 B.n318 B.n157 585
R102 B.n317 B.n316 585
R103 B.n315 B.n158 585
R104 B.n314 B.n313 585
R105 B.n312 B.n159 585
R106 B.n311 B.n310 585
R107 B.n309 B.n160 585
R108 B.n308 B.n307 585
R109 B.n306 B.n161 585
R110 B.n305 B.n304 585
R111 B.n303 B.n162 585
R112 B.n302 B.n301 585
R113 B.n300 B.n163 585
R114 B.n299 B.n298 585
R115 B.n297 B.n164 585
R116 B.n296 B.n295 585
R117 B.n294 B.n165 585
R118 B.n293 B.n292 585
R119 B.n291 B.n166 585
R120 B.n290 B.n289 585
R121 B.n288 B.n167 585
R122 B.n287 B.n286 585
R123 B.n285 B.n168 585
R124 B.n284 B.n283 585
R125 B.n282 B.n169 585
R126 B.n281 B.n280 585
R127 B.n279 B.n170 585
R128 B.n278 B.n277 585
R129 B.n276 B.n171 585
R130 B.n275 B.n274 585
R131 B.n273 B.n172 585
R132 B.n272 B.n271 585
R133 B.n270 B.n173 585
R134 B.n269 B.n268 585
R135 B.n267 B.n174 585
R136 B.n266 B.n265 585
R137 B.n264 B.n175 585
R138 B.n263 B.n262 585
R139 B.n261 B.n176 585
R140 B.n260 B.n259 585
R141 B.n258 B.n177 585
R142 B.n257 B.n256 585
R143 B.n255 B.n178 585
R144 B.n254 B.n253 585
R145 B.n252 B.n179 585
R146 B.n251 B.n250 585
R147 B.n249 B.n180 585
R148 B.n248 B.n247 585
R149 B.n246 B.n181 585
R150 B.n245 B.n244 585
R151 B.n243 B.n182 585
R152 B.n242 B.n241 585
R153 B.n240 B.n183 585
R154 B.n239 B.n238 585
R155 B.n237 B.n184 585
R156 B.n236 B.n235 585
R157 B.n234 B.n185 585
R158 B.n447 B.n446 585
R159 B.n448 B.n113 585
R160 B.n450 B.n449 585
R161 B.n451 B.n112 585
R162 B.n453 B.n452 585
R163 B.n454 B.n111 585
R164 B.n456 B.n455 585
R165 B.n457 B.n110 585
R166 B.n459 B.n458 585
R167 B.n460 B.n109 585
R168 B.n462 B.n461 585
R169 B.n463 B.n108 585
R170 B.n465 B.n464 585
R171 B.n466 B.n107 585
R172 B.n468 B.n467 585
R173 B.n469 B.n106 585
R174 B.n471 B.n470 585
R175 B.n472 B.n105 585
R176 B.n474 B.n473 585
R177 B.n475 B.n104 585
R178 B.n477 B.n476 585
R179 B.n478 B.n103 585
R180 B.n480 B.n479 585
R181 B.n481 B.n102 585
R182 B.n483 B.n482 585
R183 B.n484 B.n101 585
R184 B.n486 B.n485 585
R185 B.n487 B.n100 585
R186 B.n489 B.n488 585
R187 B.n490 B.n99 585
R188 B.n492 B.n491 585
R189 B.n493 B.n98 585
R190 B.n495 B.n494 585
R191 B.n496 B.n97 585
R192 B.n498 B.n497 585
R193 B.n499 B.n96 585
R194 B.n501 B.n500 585
R195 B.n502 B.n95 585
R196 B.n504 B.n503 585
R197 B.n505 B.n94 585
R198 B.n507 B.n506 585
R199 B.n508 B.n93 585
R200 B.n510 B.n509 585
R201 B.n511 B.n92 585
R202 B.n513 B.n512 585
R203 B.n514 B.n91 585
R204 B.n516 B.n515 585
R205 B.n517 B.n90 585
R206 B.n519 B.n518 585
R207 B.n520 B.n89 585
R208 B.n522 B.n521 585
R209 B.n523 B.n88 585
R210 B.n734 B.n733 585
R211 B.n732 B.n15 585
R212 B.n731 B.n730 585
R213 B.n729 B.n16 585
R214 B.n728 B.n727 585
R215 B.n726 B.n17 585
R216 B.n725 B.n724 585
R217 B.n723 B.n18 585
R218 B.n722 B.n721 585
R219 B.n720 B.n19 585
R220 B.n719 B.n718 585
R221 B.n717 B.n20 585
R222 B.n716 B.n715 585
R223 B.n714 B.n21 585
R224 B.n713 B.n712 585
R225 B.n711 B.n22 585
R226 B.n710 B.n709 585
R227 B.n708 B.n23 585
R228 B.n707 B.n706 585
R229 B.n705 B.n24 585
R230 B.n704 B.n703 585
R231 B.n702 B.n25 585
R232 B.n701 B.n700 585
R233 B.n699 B.n26 585
R234 B.n698 B.n697 585
R235 B.n696 B.n27 585
R236 B.n695 B.n694 585
R237 B.n693 B.n28 585
R238 B.n692 B.n691 585
R239 B.n690 B.n29 585
R240 B.n689 B.n688 585
R241 B.n687 B.n30 585
R242 B.n686 B.n685 585
R243 B.n684 B.n31 585
R244 B.n683 B.n682 585
R245 B.n681 B.n32 585
R246 B.n680 B.n679 585
R247 B.n678 B.n33 585
R248 B.n677 B.n676 585
R249 B.n675 B.n34 585
R250 B.n674 B.n673 585
R251 B.n672 B.n35 585
R252 B.n671 B.n670 585
R253 B.n669 B.n36 585
R254 B.n668 B.n667 585
R255 B.n666 B.n37 585
R256 B.n665 B.n664 585
R257 B.n663 B.n38 585
R258 B.n662 B.n661 585
R259 B.n660 B.n39 585
R260 B.n659 B.n658 585
R261 B.n657 B.n40 585
R262 B.n656 B.n655 585
R263 B.n654 B.n41 585
R264 B.n653 B.n652 585
R265 B.n651 B.n42 585
R266 B.n650 B.n649 585
R267 B.n648 B.n43 585
R268 B.n647 B.n646 585
R269 B.n645 B.n44 585
R270 B.n644 B.n643 585
R271 B.n642 B.n45 585
R272 B.n641 B.n640 585
R273 B.n639 B.n46 585
R274 B.n638 B.n637 585
R275 B.n635 B.n47 585
R276 B.n634 B.n633 585
R277 B.n632 B.n50 585
R278 B.n631 B.n630 585
R279 B.n629 B.n51 585
R280 B.n628 B.n627 585
R281 B.n626 B.n52 585
R282 B.n625 B.n624 585
R283 B.n623 B.n53 585
R284 B.n621 B.n620 585
R285 B.n619 B.n56 585
R286 B.n618 B.n617 585
R287 B.n616 B.n57 585
R288 B.n615 B.n614 585
R289 B.n613 B.n58 585
R290 B.n612 B.n611 585
R291 B.n610 B.n59 585
R292 B.n609 B.n608 585
R293 B.n607 B.n60 585
R294 B.n606 B.n605 585
R295 B.n604 B.n61 585
R296 B.n603 B.n602 585
R297 B.n601 B.n62 585
R298 B.n600 B.n599 585
R299 B.n598 B.n63 585
R300 B.n597 B.n596 585
R301 B.n595 B.n64 585
R302 B.n594 B.n593 585
R303 B.n592 B.n65 585
R304 B.n591 B.n590 585
R305 B.n589 B.n66 585
R306 B.n588 B.n587 585
R307 B.n586 B.n67 585
R308 B.n585 B.n584 585
R309 B.n583 B.n68 585
R310 B.n582 B.n581 585
R311 B.n580 B.n69 585
R312 B.n579 B.n578 585
R313 B.n577 B.n70 585
R314 B.n576 B.n575 585
R315 B.n574 B.n71 585
R316 B.n573 B.n572 585
R317 B.n571 B.n72 585
R318 B.n570 B.n569 585
R319 B.n568 B.n73 585
R320 B.n567 B.n566 585
R321 B.n565 B.n74 585
R322 B.n564 B.n563 585
R323 B.n562 B.n75 585
R324 B.n561 B.n560 585
R325 B.n559 B.n76 585
R326 B.n558 B.n557 585
R327 B.n556 B.n77 585
R328 B.n555 B.n554 585
R329 B.n553 B.n78 585
R330 B.n552 B.n551 585
R331 B.n550 B.n79 585
R332 B.n549 B.n548 585
R333 B.n547 B.n80 585
R334 B.n546 B.n545 585
R335 B.n544 B.n81 585
R336 B.n543 B.n542 585
R337 B.n541 B.n82 585
R338 B.n540 B.n539 585
R339 B.n538 B.n83 585
R340 B.n537 B.n536 585
R341 B.n535 B.n84 585
R342 B.n534 B.n533 585
R343 B.n532 B.n85 585
R344 B.n531 B.n530 585
R345 B.n529 B.n86 585
R346 B.n528 B.n527 585
R347 B.n526 B.n87 585
R348 B.n525 B.n524 585
R349 B.n735 B.n14 585
R350 B.n737 B.n736 585
R351 B.n738 B.n13 585
R352 B.n740 B.n739 585
R353 B.n741 B.n12 585
R354 B.n743 B.n742 585
R355 B.n744 B.n11 585
R356 B.n746 B.n745 585
R357 B.n747 B.n10 585
R358 B.n749 B.n748 585
R359 B.n750 B.n9 585
R360 B.n752 B.n751 585
R361 B.n753 B.n8 585
R362 B.n755 B.n754 585
R363 B.n756 B.n7 585
R364 B.n758 B.n757 585
R365 B.n759 B.n6 585
R366 B.n761 B.n760 585
R367 B.n762 B.n5 585
R368 B.n764 B.n763 585
R369 B.n765 B.n4 585
R370 B.n767 B.n766 585
R371 B.n768 B.n3 585
R372 B.n770 B.n769 585
R373 B.n771 B.n0 585
R374 B.n2 B.n1 585
R375 B.n198 B.n197 585
R376 B.n200 B.n199 585
R377 B.n201 B.n196 585
R378 B.n203 B.n202 585
R379 B.n204 B.n195 585
R380 B.n206 B.n205 585
R381 B.n207 B.n194 585
R382 B.n209 B.n208 585
R383 B.n210 B.n193 585
R384 B.n212 B.n211 585
R385 B.n213 B.n192 585
R386 B.n215 B.n214 585
R387 B.n216 B.n191 585
R388 B.n218 B.n217 585
R389 B.n219 B.n190 585
R390 B.n221 B.n220 585
R391 B.n222 B.n189 585
R392 B.n224 B.n223 585
R393 B.n225 B.n188 585
R394 B.n227 B.n226 585
R395 B.n228 B.n187 585
R396 B.n230 B.n229 585
R397 B.n231 B.n186 585
R398 B.n233 B.n232 585
R399 B.n232 B.n185 497.305
R400 B.n446 B.n445 497.305
R401 B.n524 B.n523 497.305
R402 B.n735 B.n734 497.305
R403 B.n152 B.t6 387.346
R404 B.n344 B.t9 387.346
R405 B.n54 B.t0 387.346
R406 B.n48 B.t3 387.346
R407 B.n773 B.n772 256.663
R408 B.n772 B.n771 235.042
R409 B.n772 B.n2 235.042
R410 B.n344 B.t10 165.196
R411 B.n54 B.t2 165.196
R412 B.n152 B.t7 165.169
R413 B.n48 B.t5 165.169
R414 B.n236 B.n185 163.367
R415 B.n237 B.n236 163.367
R416 B.n238 B.n237 163.367
R417 B.n238 B.n183 163.367
R418 B.n242 B.n183 163.367
R419 B.n243 B.n242 163.367
R420 B.n244 B.n243 163.367
R421 B.n244 B.n181 163.367
R422 B.n248 B.n181 163.367
R423 B.n249 B.n248 163.367
R424 B.n250 B.n249 163.367
R425 B.n250 B.n179 163.367
R426 B.n254 B.n179 163.367
R427 B.n255 B.n254 163.367
R428 B.n256 B.n255 163.367
R429 B.n256 B.n177 163.367
R430 B.n260 B.n177 163.367
R431 B.n261 B.n260 163.367
R432 B.n262 B.n261 163.367
R433 B.n262 B.n175 163.367
R434 B.n266 B.n175 163.367
R435 B.n267 B.n266 163.367
R436 B.n268 B.n267 163.367
R437 B.n268 B.n173 163.367
R438 B.n272 B.n173 163.367
R439 B.n273 B.n272 163.367
R440 B.n274 B.n273 163.367
R441 B.n274 B.n171 163.367
R442 B.n278 B.n171 163.367
R443 B.n279 B.n278 163.367
R444 B.n280 B.n279 163.367
R445 B.n280 B.n169 163.367
R446 B.n284 B.n169 163.367
R447 B.n285 B.n284 163.367
R448 B.n286 B.n285 163.367
R449 B.n286 B.n167 163.367
R450 B.n290 B.n167 163.367
R451 B.n291 B.n290 163.367
R452 B.n292 B.n291 163.367
R453 B.n292 B.n165 163.367
R454 B.n296 B.n165 163.367
R455 B.n297 B.n296 163.367
R456 B.n298 B.n297 163.367
R457 B.n298 B.n163 163.367
R458 B.n302 B.n163 163.367
R459 B.n303 B.n302 163.367
R460 B.n304 B.n303 163.367
R461 B.n304 B.n161 163.367
R462 B.n308 B.n161 163.367
R463 B.n309 B.n308 163.367
R464 B.n310 B.n309 163.367
R465 B.n310 B.n159 163.367
R466 B.n314 B.n159 163.367
R467 B.n315 B.n314 163.367
R468 B.n316 B.n315 163.367
R469 B.n316 B.n157 163.367
R470 B.n320 B.n157 163.367
R471 B.n321 B.n320 163.367
R472 B.n322 B.n321 163.367
R473 B.n322 B.n155 163.367
R474 B.n326 B.n155 163.367
R475 B.n327 B.n326 163.367
R476 B.n328 B.n327 163.367
R477 B.n328 B.n151 163.367
R478 B.n333 B.n151 163.367
R479 B.n334 B.n333 163.367
R480 B.n335 B.n334 163.367
R481 B.n335 B.n149 163.367
R482 B.n339 B.n149 163.367
R483 B.n340 B.n339 163.367
R484 B.n341 B.n340 163.367
R485 B.n341 B.n147 163.367
R486 B.n348 B.n147 163.367
R487 B.n349 B.n348 163.367
R488 B.n350 B.n349 163.367
R489 B.n350 B.n145 163.367
R490 B.n354 B.n145 163.367
R491 B.n355 B.n354 163.367
R492 B.n356 B.n355 163.367
R493 B.n356 B.n143 163.367
R494 B.n360 B.n143 163.367
R495 B.n361 B.n360 163.367
R496 B.n362 B.n361 163.367
R497 B.n362 B.n141 163.367
R498 B.n366 B.n141 163.367
R499 B.n367 B.n366 163.367
R500 B.n368 B.n367 163.367
R501 B.n368 B.n139 163.367
R502 B.n372 B.n139 163.367
R503 B.n373 B.n372 163.367
R504 B.n374 B.n373 163.367
R505 B.n374 B.n137 163.367
R506 B.n378 B.n137 163.367
R507 B.n379 B.n378 163.367
R508 B.n380 B.n379 163.367
R509 B.n380 B.n135 163.367
R510 B.n384 B.n135 163.367
R511 B.n385 B.n384 163.367
R512 B.n386 B.n385 163.367
R513 B.n386 B.n133 163.367
R514 B.n390 B.n133 163.367
R515 B.n391 B.n390 163.367
R516 B.n392 B.n391 163.367
R517 B.n392 B.n131 163.367
R518 B.n396 B.n131 163.367
R519 B.n397 B.n396 163.367
R520 B.n398 B.n397 163.367
R521 B.n398 B.n129 163.367
R522 B.n402 B.n129 163.367
R523 B.n403 B.n402 163.367
R524 B.n404 B.n403 163.367
R525 B.n404 B.n127 163.367
R526 B.n408 B.n127 163.367
R527 B.n409 B.n408 163.367
R528 B.n410 B.n409 163.367
R529 B.n410 B.n125 163.367
R530 B.n414 B.n125 163.367
R531 B.n415 B.n414 163.367
R532 B.n416 B.n415 163.367
R533 B.n416 B.n123 163.367
R534 B.n420 B.n123 163.367
R535 B.n421 B.n420 163.367
R536 B.n422 B.n421 163.367
R537 B.n422 B.n121 163.367
R538 B.n426 B.n121 163.367
R539 B.n427 B.n426 163.367
R540 B.n428 B.n427 163.367
R541 B.n428 B.n119 163.367
R542 B.n432 B.n119 163.367
R543 B.n433 B.n432 163.367
R544 B.n434 B.n433 163.367
R545 B.n434 B.n117 163.367
R546 B.n438 B.n117 163.367
R547 B.n439 B.n438 163.367
R548 B.n440 B.n439 163.367
R549 B.n440 B.n115 163.367
R550 B.n444 B.n115 163.367
R551 B.n445 B.n444 163.367
R552 B.n523 B.n522 163.367
R553 B.n522 B.n89 163.367
R554 B.n518 B.n89 163.367
R555 B.n518 B.n517 163.367
R556 B.n517 B.n516 163.367
R557 B.n516 B.n91 163.367
R558 B.n512 B.n91 163.367
R559 B.n512 B.n511 163.367
R560 B.n511 B.n510 163.367
R561 B.n510 B.n93 163.367
R562 B.n506 B.n93 163.367
R563 B.n506 B.n505 163.367
R564 B.n505 B.n504 163.367
R565 B.n504 B.n95 163.367
R566 B.n500 B.n95 163.367
R567 B.n500 B.n499 163.367
R568 B.n499 B.n498 163.367
R569 B.n498 B.n97 163.367
R570 B.n494 B.n97 163.367
R571 B.n494 B.n493 163.367
R572 B.n493 B.n492 163.367
R573 B.n492 B.n99 163.367
R574 B.n488 B.n99 163.367
R575 B.n488 B.n487 163.367
R576 B.n487 B.n486 163.367
R577 B.n486 B.n101 163.367
R578 B.n482 B.n101 163.367
R579 B.n482 B.n481 163.367
R580 B.n481 B.n480 163.367
R581 B.n480 B.n103 163.367
R582 B.n476 B.n103 163.367
R583 B.n476 B.n475 163.367
R584 B.n475 B.n474 163.367
R585 B.n474 B.n105 163.367
R586 B.n470 B.n105 163.367
R587 B.n470 B.n469 163.367
R588 B.n469 B.n468 163.367
R589 B.n468 B.n107 163.367
R590 B.n464 B.n107 163.367
R591 B.n464 B.n463 163.367
R592 B.n463 B.n462 163.367
R593 B.n462 B.n109 163.367
R594 B.n458 B.n109 163.367
R595 B.n458 B.n457 163.367
R596 B.n457 B.n456 163.367
R597 B.n456 B.n111 163.367
R598 B.n452 B.n111 163.367
R599 B.n452 B.n451 163.367
R600 B.n451 B.n450 163.367
R601 B.n450 B.n113 163.367
R602 B.n446 B.n113 163.367
R603 B.n734 B.n15 163.367
R604 B.n730 B.n15 163.367
R605 B.n730 B.n729 163.367
R606 B.n729 B.n728 163.367
R607 B.n728 B.n17 163.367
R608 B.n724 B.n17 163.367
R609 B.n724 B.n723 163.367
R610 B.n723 B.n722 163.367
R611 B.n722 B.n19 163.367
R612 B.n718 B.n19 163.367
R613 B.n718 B.n717 163.367
R614 B.n717 B.n716 163.367
R615 B.n716 B.n21 163.367
R616 B.n712 B.n21 163.367
R617 B.n712 B.n711 163.367
R618 B.n711 B.n710 163.367
R619 B.n710 B.n23 163.367
R620 B.n706 B.n23 163.367
R621 B.n706 B.n705 163.367
R622 B.n705 B.n704 163.367
R623 B.n704 B.n25 163.367
R624 B.n700 B.n25 163.367
R625 B.n700 B.n699 163.367
R626 B.n699 B.n698 163.367
R627 B.n698 B.n27 163.367
R628 B.n694 B.n27 163.367
R629 B.n694 B.n693 163.367
R630 B.n693 B.n692 163.367
R631 B.n692 B.n29 163.367
R632 B.n688 B.n29 163.367
R633 B.n688 B.n687 163.367
R634 B.n687 B.n686 163.367
R635 B.n686 B.n31 163.367
R636 B.n682 B.n31 163.367
R637 B.n682 B.n681 163.367
R638 B.n681 B.n680 163.367
R639 B.n680 B.n33 163.367
R640 B.n676 B.n33 163.367
R641 B.n676 B.n675 163.367
R642 B.n675 B.n674 163.367
R643 B.n674 B.n35 163.367
R644 B.n670 B.n35 163.367
R645 B.n670 B.n669 163.367
R646 B.n669 B.n668 163.367
R647 B.n668 B.n37 163.367
R648 B.n664 B.n37 163.367
R649 B.n664 B.n663 163.367
R650 B.n663 B.n662 163.367
R651 B.n662 B.n39 163.367
R652 B.n658 B.n39 163.367
R653 B.n658 B.n657 163.367
R654 B.n657 B.n656 163.367
R655 B.n656 B.n41 163.367
R656 B.n652 B.n41 163.367
R657 B.n652 B.n651 163.367
R658 B.n651 B.n650 163.367
R659 B.n650 B.n43 163.367
R660 B.n646 B.n43 163.367
R661 B.n646 B.n645 163.367
R662 B.n645 B.n644 163.367
R663 B.n644 B.n45 163.367
R664 B.n640 B.n45 163.367
R665 B.n640 B.n639 163.367
R666 B.n639 B.n638 163.367
R667 B.n638 B.n47 163.367
R668 B.n633 B.n47 163.367
R669 B.n633 B.n632 163.367
R670 B.n632 B.n631 163.367
R671 B.n631 B.n51 163.367
R672 B.n627 B.n51 163.367
R673 B.n627 B.n626 163.367
R674 B.n626 B.n625 163.367
R675 B.n625 B.n53 163.367
R676 B.n620 B.n53 163.367
R677 B.n620 B.n619 163.367
R678 B.n619 B.n618 163.367
R679 B.n618 B.n57 163.367
R680 B.n614 B.n57 163.367
R681 B.n614 B.n613 163.367
R682 B.n613 B.n612 163.367
R683 B.n612 B.n59 163.367
R684 B.n608 B.n59 163.367
R685 B.n608 B.n607 163.367
R686 B.n607 B.n606 163.367
R687 B.n606 B.n61 163.367
R688 B.n602 B.n61 163.367
R689 B.n602 B.n601 163.367
R690 B.n601 B.n600 163.367
R691 B.n600 B.n63 163.367
R692 B.n596 B.n63 163.367
R693 B.n596 B.n595 163.367
R694 B.n595 B.n594 163.367
R695 B.n594 B.n65 163.367
R696 B.n590 B.n65 163.367
R697 B.n590 B.n589 163.367
R698 B.n589 B.n588 163.367
R699 B.n588 B.n67 163.367
R700 B.n584 B.n67 163.367
R701 B.n584 B.n583 163.367
R702 B.n583 B.n582 163.367
R703 B.n582 B.n69 163.367
R704 B.n578 B.n69 163.367
R705 B.n578 B.n577 163.367
R706 B.n577 B.n576 163.367
R707 B.n576 B.n71 163.367
R708 B.n572 B.n71 163.367
R709 B.n572 B.n571 163.367
R710 B.n571 B.n570 163.367
R711 B.n570 B.n73 163.367
R712 B.n566 B.n73 163.367
R713 B.n566 B.n565 163.367
R714 B.n565 B.n564 163.367
R715 B.n564 B.n75 163.367
R716 B.n560 B.n75 163.367
R717 B.n560 B.n559 163.367
R718 B.n559 B.n558 163.367
R719 B.n558 B.n77 163.367
R720 B.n554 B.n77 163.367
R721 B.n554 B.n553 163.367
R722 B.n553 B.n552 163.367
R723 B.n552 B.n79 163.367
R724 B.n548 B.n79 163.367
R725 B.n548 B.n547 163.367
R726 B.n547 B.n546 163.367
R727 B.n546 B.n81 163.367
R728 B.n542 B.n81 163.367
R729 B.n542 B.n541 163.367
R730 B.n541 B.n540 163.367
R731 B.n540 B.n83 163.367
R732 B.n536 B.n83 163.367
R733 B.n536 B.n535 163.367
R734 B.n535 B.n534 163.367
R735 B.n534 B.n85 163.367
R736 B.n530 B.n85 163.367
R737 B.n530 B.n529 163.367
R738 B.n529 B.n528 163.367
R739 B.n528 B.n87 163.367
R740 B.n524 B.n87 163.367
R741 B.n736 B.n735 163.367
R742 B.n736 B.n13 163.367
R743 B.n740 B.n13 163.367
R744 B.n741 B.n740 163.367
R745 B.n742 B.n741 163.367
R746 B.n742 B.n11 163.367
R747 B.n746 B.n11 163.367
R748 B.n747 B.n746 163.367
R749 B.n748 B.n747 163.367
R750 B.n748 B.n9 163.367
R751 B.n752 B.n9 163.367
R752 B.n753 B.n752 163.367
R753 B.n754 B.n753 163.367
R754 B.n754 B.n7 163.367
R755 B.n758 B.n7 163.367
R756 B.n759 B.n758 163.367
R757 B.n760 B.n759 163.367
R758 B.n760 B.n5 163.367
R759 B.n764 B.n5 163.367
R760 B.n765 B.n764 163.367
R761 B.n766 B.n765 163.367
R762 B.n766 B.n3 163.367
R763 B.n770 B.n3 163.367
R764 B.n771 B.n770 163.367
R765 B.n197 B.n2 163.367
R766 B.n200 B.n197 163.367
R767 B.n201 B.n200 163.367
R768 B.n202 B.n201 163.367
R769 B.n202 B.n195 163.367
R770 B.n206 B.n195 163.367
R771 B.n207 B.n206 163.367
R772 B.n208 B.n207 163.367
R773 B.n208 B.n193 163.367
R774 B.n212 B.n193 163.367
R775 B.n213 B.n212 163.367
R776 B.n214 B.n213 163.367
R777 B.n214 B.n191 163.367
R778 B.n218 B.n191 163.367
R779 B.n219 B.n218 163.367
R780 B.n220 B.n219 163.367
R781 B.n220 B.n189 163.367
R782 B.n224 B.n189 163.367
R783 B.n225 B.n224 163.367
R784 B.n226 B.n225 163.367
R785 B.n226 B.n187 163.367
R786 B.n230 B.n187 163.367
R787 B.n231 B.n230 163.367
R788 B.n232 B.n231 163.367
R789 B.n345 B.t11 107.207
R790 B.n55 B.t1 107.207
R791 B.n153 B.t8 107.181
R792 B.n49 B.t4 107.181
R793 B.n331 B.n153 59.5399
R794 B.n346 B.n345 59.5399
R795 B.n622 B.n55 59.5399
R796 B.n636 B.n49 59.5399
R797 B.n153 B.n152 57.9884
R798 B.n345 B.n344 57.9884
R799 B.n55 B.n54 57.9884
R800 B.n49 B.n48 57.9884
R801 B.n733 B.n14 32.3127
R802 B.n525 B.n88 32.3127
R803 B.n447 B.n114 32.3127
R804 B.n234 B.n233 32.3127
R805 B B.n773 18.0485
R806 B.n737 B.n14 10.6151
R807 B.n738 B.n737 10.6151
R808 B.n739 B.n738 10.6151
R809 B.n739 B.n12 10.6151
R810 B.n743 B.n12 10.6151
R811 B.n744 B.n743 10.6151
R812 B.n745 B.n744 10.6151
R813 B.n745 B.n10 10.6151
R814 B.n749 B.n10 10.6151
R815 B.n750 B.n749 10.6151
R816 B.n751 B.n750 10.6151
R817 B.n751 B.n8 10.6151
R818 B.n755 B.n8 10.6151
R819 B.n756 B.n755 10.6151
R820 B.n757 B.n756 10.6151
R821 B.n757 B.n6 10.6151
R822 B.n761 B.n6 10.6151
R823 B.n762 B.n761 10.6151
R824 B.n763 B.n762 10.6151
R825 B.n763 B.n4 10.6151
R826 B.n767 B.n4 10.6151
R827 B.n768 B.n767 10.6151
R828 B.n769 B.n768 10.6151
R829 B.n769 B.n0 10.6151
R830 B.n733 B.n732 10.6151
R831 B.n732 B.n731 10.6151
R832 B.n731 B.n16 10.6151
R833 B.n727 B.n16 10.6151
R834 B.n727 B.n726 10.6151
R835 B.n726 B.n725 10.6151
R836 B.n725 B.n18 10.6151
R837 B.n721 B.n18 10.6151
R838 B.n721 B.n720 10.6151
R839 B.n720 B.n719 10.6151
R840 B.n719 B.n20 10.6151
R841 B.n715 B.n20 10.6151
R842 B.n715 B.n714 10.6151
R843 B.n714 B.n713 10.6151
R844 B.n713 B.n22 10.6151
R845 B.n709 B.n22 10.6151
R846 B.n709 B.n708 10.6151
R847 B.n708 B.n707 10.6151
R848 B.n707 B.n24 10.6151
R849 B.n703 B.n24 10.6151
R850 B.n703 B.n702 10.6151
R851 B.n702 B.n701 10.6151
R852 B.n701 B.n26 10.6151
R853 B.n697 B.n26 10.6151
R854 B.n697 B.n696 10.6151
R855 B.n696 B.n695 10.6151
R856 B.n695 B.n28 10.6151
R857 B.n691 B.n28 10.6151
R858 B.n691 B.n690 10.6151
R859 B.n690 B.n689 10.6151
R860 B.n689 B.n30 10.6151
R861 B.n685 B.n30 10.6151
R862 B.n685 B.n684 10.6151
R863 B.n684 B.n683 10.6151
R864 B.n683 B.n32 10.6151
R865 B.n679 B.n32 10.6151
R866 B.n679 B.n678 10.6151
R867 B.n678 B.n677 10.6151
R868 B.n677 B.n34 10.6151
R869 B.n673 B.n34 10.6151
R870 B.n673 B.n672 10.6151
R871 B.n672 B.n671 10.6151
R872 B.n671 B.n36 10.6151
R873 B.n667 B.n36 10.6151
R874 B.n667 B.n666 10.6151
R875 B.n666 B.n665 10.6151
R876 B.n665 B.n38 10.6151
R877 B.n661 B.n38 10.6151
R878 B.n661 B.n660 10.6151
R879 B.n660 B.n659 10.6151
R880 B.n659 B.n40 10.6151
R881 B.n655 B.n40 10.6151
R882 B.n655 B.n654 10.6151
R883 B.n654 B.n653 10.6151
R884 B.n653 B.n42 10.6151
R885 B.n649 B.n42 10.6151
R886 B.n649 B.n648 10.6151
R887 B.n648 B.n647 10.6151
R888 B.n647 B.n44 10.6151
R889 B.n643 B.n44 10.6151
R890 B.n643 B.n642 10.6151
R891 B.n642 B.n641 10.6151
R892 B.n641 B.n46 10.6151
R893 B.n637 B.n46 10.6151
R894 B.n635 B.n634 10.6151
R895 B.n634 B.n50 10.6151
R896 B.n630 B.n50 10.6151
R897 B.n630 B.n629 10.6151
R898 B.n629 B.n628 10.6151
R899 B.n628 B.n52 10.6151
R900 B.n624 B.n52 10.6151
R901 B.n624 B.n623 10.6151
R902 B.n621 B.n56 10.6151
R903 B.n617 B.n56 10.6151
R904 B.n617 B.n616 10.6151
R905 B.n616 B.n615 10.6151
R906 B.n615 B.n58 10.6151
R907 B.n611 B.n58 10.6151
R908 B.n611 B.n610 10.6151
R909 B.n610 B.n609 10.6151
R910 B.n609 B.n60 10.6151
R911 B.n605 B.n60 10.6151
R912 B.n605 B.n604 10.6151
R913 B.n604 B.n603 10.6151
R914 B.n603 B.n62 10.6151
R915 B.n599 B.n62 10.6151
R916 B.n599 B.n598 10.6151
R917 B.n598 B.n597 10.6151
R918 B.n597 B.n64 10.6151
R919 B.n593 B.n64 10.6151
R920 B.n593 B.n592 10.6151
R921 B.n592 B.n591 10.6151
R922 B.n591 B.n66 10.6151
R923 B.n587 B.n66 10.6151
R924 B.n587 B.n586 10.6151
R925 B.n586 B.n585 10.6151
R926 B.n585 B.n68 10.6151
R927 B.n581 B.n68 10.6151
R928 B.n581 B.n580 10.6151
R929 B.n580 B.n579 10.6151
R930 B.n579 B.n70 10.6151
R931 B.n575 B.n70 10.6151
R932 B.n575 B.n574 10.6151
R933 B.n574 B.n573 10.6151
R934 B.n573 B.n72 10.6151
R935 B.n569 B.n72 10.6151
R936 B.n569 B.n568 10.6151
R937 B.n568 B.n567 10.6151
R938 B.n567 B.n74 10.6151
R939 B.n563 B.n74 10.6151
R940 B.n563 B.n562 10.6151
R941 B.n562 B.n561 10.6151
R942 B.n561 B.n76 10.6151
R943 B.n557 B.n76 10.6151
R944 B.n557 B.n556 10.6151
R945 B.n556 B.n555 10.6151
R946 B.n555 B.n78 10.6151
R947 B.n551 B.n78 10.6151
R948 B.n551 B.n550 10.6151
R949 B.n550 B.n549 10.6151
R950 B.n549 B.n80 10.6151
R951 B.n545 B.n80 10.6151
R952 B.n545 B.n544 10.6151
R953 B.n544 B.n543 10.6151
R954 B.n543 B.n82 10.6151
R955 B.n539 B.n82 10.6151
R956 B.n539 B.n538 10.6151
R957 B.n538 B.n537 10.6151
R958 B.n537 B.n84 10.6151
R959 B.n533 B.n84 10.6151
R960 B.n533 B.n532 10.6151
R961 B.n532 B.n531 10.6151
R962 B.n531 B.n86 10.6151
R963 B.n527 B.n86 10.6151
R964 B.n527 B.n526 10.6151
R965 B.n526 B.n525 10.6151
R966 B.n521 B.n88 10.6151
R967 B.n521 B.n520 10.6151
R968 B.n520 B.n519 10.6151
R969 B.n519 B.n90 10.6151
R970 B.n515 B.n90 10.6151
R971 B.n515 B.n514 10.6151
R972 B.n514 B.n513 10.6151
R973 B.n513 B.n92 10.6151
R974 B.n509 B.n92 10.6151
R975 B.n509 B.n508 10.6151
R976 B.n508 B.n507 10.6151
R977 B.n507 B.n94 10.6151
R978 B.n503 B.n94 10.6151
R979 B.n503 B.n502 10.6151
R980 B.n502 B.n501 10.6151
R981 B.n501 B.n96 10.6151
R982 B.n497 B.n96 10.6151
R983 B.n497 B.n496 10.6151
R984 B.n496 B.n495 10.6151
R985 B.n495 B.n98 10.6151
R986 B.n491 B.n98 10.6151
R987 B.n491 B.n490 10.6151
R988 B.n490 B.n489 10.6151
R989 B.n489 B.n100 10.6151
R990 B.n485 B.n100 10.6151
R991 B.n485 B.n484 10.6151
R992 B.n484 B.n483 10.6151
R993 B.n483 B.n102 10.6151
R994 B.n479 B.n102 10.6151
R995 B.n479 B.n478 10.6151
R996 B.n478 B.n477 10.6151
R997 B.n477 B.n104 10.6151
R998 B.n473 B.n104 10.6151
R999 B.n473 B.n472 10.6151
R1000 B.n472 B.n471 10.6151
R1001 B.n471 B.n106 10.6151
R1002 B.n467 B.n106 10.6151
R1003 B.n467 B.n466 10.6151
R1004 B.n466 B.n465 10.6151
R1005 B.n465 B.n108 10.6151
R1006 B.n461 B.n108 10.6151
R1007 B.n461 B.n460 10.6151
R1008 B.n460 B.n459 10.6151
R1009 B.n459 B.n110 10.6151
R1010 B.n455 B.n110 10.6151
R1011 B.n455 B.n454 10.6151
R1012 B.n454 B.n453 10.6151
R1013 B.n453 B.n112 10.6151
R1014 B.n449 B.n112 10.6151
R1015 B.n449 B.n448 10.6151
R1016 B.n448 B.n447 10.6151
R1017 B.n198 B.n1 10.6151
R1018 B.n199 B.n198 10.6151
R1019 B.n199 B.n196 10.6151
R1020 B.n203 B.n196 10.6151
R1021 B.n204 B.n203 10.6151
R1022 B.n205 B.n204 10.6151
R1023 B.n205 B.n194 10.6151
R1024 B.n209 B.n194 10.6151
R1025 B.n210 B.n209 10.6151
R1026 B.n211 B.n210 10.6151
R1027 B.n211 B.n192 10.6151
R1028 B.n215 B.n192 10.6151
R1029 B.n216 B.n215 10.6151
R1030 B.n217 B.n216 10.6151
R1031 B.n217 B.n190 10.6151
R1032 B.n221 B.n190 10.6151
R1033 B.n222 B.n221 10.6151
R1034 B.n223 B.n222 10.6151
R1035 B.n223 B.n188 10.6151
R1036 B.n227 B.n188 10.6151
R1037 B.n228 B.n227 10.6151
R1038 B.n229 B.n228 10.6151
R1039 B.n229 B.n186 10.6151
R1040 B.n233 B.n186 10.6151
R1041 B.n235 B.n234 10.6151
R1042 B.n235 B.n184 10.6151
R1043 B.n239 B.n184 10.6151
R1044 B.n240 B.n239 10.6151
R1045 B.n241 B.n240 10.6151
R1046 B.n241 B.n182 10.6151
R1047 B.n245 B.n182 10.6151
R1048 B.n246 B.n245 10.6151
R1049 B.n247 B.n246 10.6151
R1050 B.n247 B.n180 10.6151
R1051 B.n251 B.n180 10.6151
R1052 B.n252 B.n251 10.6151
R1053 B.n253 B.n252 10.6151
R1054 B.n253 B.n178 10.6151
R1055 B.n257 B.n178 10.6151
R1056 B.n258 B.n257 10.6151
R1057 B.n259 B.n258 10.6151
R1058 B.n259 B.n176 10.6151
R1059 B.n263 B.n176 10.6151
R1060 B.n264 B.n263 10.6151
R1061 B.n265 B.n264 10.6151
R1062 B.n265 B.n174 10.6151
R1063 B.n269 B.n174 10.6151
R1064 B.n270 B.n269 10.6151
R1065 B.n271 B.n270 10.6151
R1066 B.n271 B.n172 10.6151
R1067 B.n275 B.n172 10.6151
R1068 B.n276 B.n275 10.6151
R1069 B.n277 B.n276 10.6151
R1070 B.n277 B.n170 10.6151
R1071 B.n281 B.n170 10.6151
R1072 B.n282 B.n281 10.6151
R1073 B.n283 B.n282 10.6151
R1074 B.n283 B.n168 10.6151
R1075 B.n287 B.n168 10.6151
R1076 B.n288 B.n287 10.6151
R1077 B.n289 B.n288 10.6151
R1078 B.n289 B.n166 10.6151
R1079 B.n293 B.n166 10.6151
R1080 B.n294 B.n293 10.6151
R1081 B.n295 B.n294 10.6151
R1082 B.n295 B.n164 10.6151
R1083 B.n299 B.n164 10.6151
R1084 B.n300 B.n299 10.6151
R1085 B.n301 B.n300 10.6151
R1086 B.n301 B.n162 10.6151
R1087 B.n305 B.n162 10.6151
R1088 B.n306 B.n305 10.6151
R1089 B.n307 B.n306 10.6151
R1090 B.n307 B.n160 10.6151
R1091 B.n311 B.n160 10.6151
R1092 B.n312 B.n311 10.6151
R1093 B.n313 B.n312 10.6151
R1094 B.n313 B.n158 10.6151
R1095 B.n317 B.n158 10.6151
R1096 B.n318 B.n317 10.6151
R1097 B.n319 B.n318 10.6151
R1098 B.n319 B.n156 10.6151
R1099 B.n323 B.n156 10.6151
R1100 B.n324 B.n323 10.6151
R1101 B.n325 B.n324 10.6151
R1102 B.n325 B.n154 10.6151
R1103 B.n329 B.n154 10.6151
R1104 B.n330 B.n329 10.6151
R1105 B.n332 B.n150 10.6151
R1106 B.n336 B.n150 10.6151
R1107 B.n337 B.n336 10.6151
R1108 B.n338 B.n337 10.6151
R1109 B.n338 B.n148 10.6151
R1110 B.n342 B.n148 10.6151
R1111 B.n343 B.n342 10.6151
R1112 B.n347 B.n343 10.6151
R1113 B.n351 B.n146 10.6151
R1114 B.n352 B.n351 10.6151
R1115 B.n353 B.n352 10.6151
R1116 B.n353 B.n144 10.6151
R1117 B.n357 B.n144 10.6151
R1118 B.n358 B.n357 10.6151
R1119 B.n359 B.n358 10.6151
R1120 B.n359 B.n142 10.6151
R1121 B.n363 B.n142 10.6151
R1122 B.n364 B.n363 10.6151
R1123 B.n365 B.n364 10.6151
R1124 B.n365 B.n140 10.6151
R1125 B.n369 B.n140 10.6151
R1126 B.n370 B.n369 10.6151
R1127 B.n371 B.n370 10.6151
R1128 B.n371 B.n138 10.6151
R1129 B.n375 B.n138 10.6151
R1130 B.n376 B.n375 10.6151
R1131 B.n377 B.n376 10.6151
R1132 B.n377 B.n136 10.6151
R1133 B.n381 B.n136 10.6151
R1134 B.n382 B.n381 10.6151
R1135 B.n383 B.n382 10.6151
R1136 B.n383 B.n134 10.6151
R1137 B.n387 B.n134 10.6151
R1138 B.n388 B.n387 10.6151
R1139 B.n389 B.n388 10.6151
R1140 B.n389 B.n132 10.6151
R1141 B.n393 B.n132 10.6151
R1142 B.n394 B.n393 10.6151
R1143 B.n395 B.n394 10.6151
R1144 B.n395 B.n130 10.6151
R1145 B.n399 B.n130 10.6151
R1146 B.n400 B.n399 10.6151
R1147 B.n401 B.n400 10.6151
R1148 B.n401 B.n128 10.6151
R1149 B.n405 B.n128 10.6151
R1150 B.n406 B.n405 10.6151
R1151 B.n407 B.n406 10.6151
R1152 B.n407 B.n126 10.6151
R1153 B.n411 B.n126 10.6151
R1154 B.n412 B.n411 10.6151
R1155 B.n413 B.n412 10.6151
R1156 B.n413 B.n124 10.6151
R1157 B.n417 B.n124 10.6151
R1158 B.n418 B.n417 10.6151
R1159 B.n419 B.n418 10.6151
R1160 B.n419 B.n122 10.6151
R1161 B.n423 B.n122 10.6151
R1162 B.n424 B.n423 10.6151
R1163 B.n425 B.n424 10.6151
R1164 B.n425 B.n120 10.6151
R1165 B.n429 B.n120 10.6151
R1166 B.n430 B.n429 10.6151
R1167 B.n431 B.n430 10.6151
R1168 B.n431 B.n118 10.6151
R1169 B.n435 B.n118 10.6151
R1170 B.n436 B.n435 10.6151
R1171 B.n437 B.n436 10.6151
R1172 B.n437 B.n116 10.6151
R1173 B.n441 B.n116 10.6151
R1174 B.n442 B.n441 10.6151
R1175 B.n443 B.n442 10.6151
R1176 B.n443 B.n114 10.6151
R1177 B.n773 B.n0 8.11757
R1178 B.n773 B.n1 8.11757
R1179 B.n636 B.n635 6.5566
R1180 B.n623 B.n622 6.5566
R1181 B.n332 B.n331 6.5566
R1182 B.n347 B.n346 6.5566
R1183 B.n637 B.n636 4.05904
R1184 B.n622 B.n621 4.05904
R1185 B.n331 B.n330 4.05904
R1186 B.n346 B.n146 4.05904
C0 w_n2166_n4924# VN 3.15931f
C1 VDD2 VN 4.43726f
C2 w_n2166_n4924# VP 3.43535f
C3 w_n2166_n4924# B 11.0549f
C4 w_n2166_n4924# VTAIL 3.83128f
C5 VDD2 VP 0.335861f
C6 VN VDD1 0.147815f
C7 VDD2 B 2.35992f
C8 VDD2 VTAIL 7.17229f
C9 VP VDD1 4.62147f
C10 B VDD1 2.3293f
C11 VDD1 VTAIL 7.12298f
C12 VDD2 w_n2166_n4924# 2.3541f
C13 w_n2166_n4924# VDD1 2.32748f
C14 VDD2 VDD1 0.682727f
C15 VN VP 6.93152f
C16 VN B 1.14754f
C17 VN VTAIL 3.75713f
C18 B VP 1.60159f
C19 VP VTAIL 3.77153f
C20 B VTAIL 5.43166f
C21 VDD2 VSUBS 1.18629f
C22 VDD1 VSUBS 6.9201f
C23 VTAIL VSUBS 1.313434f
C24 VN VSUBS 9.54378f
C25 VP VSUBS 1.988365f
C26 B VSUBS 4.611975f
C27 w_n2166_n4924# VSUBS 0.130246p
C28 B.n0 VSUBS 0.005908f
C29 B.n1 VSUBS 0.005908f
C30 B.n2 VSUBS 0.008737f
C31 B.n3 VSUBS 0.006696f
C32 B.n4 VSUBS 0.006696f
C33 B.n5 VSUBS 0.006696f
C34 B.n6 VSUBS 0.006696f
C35 B.n7 VSUBS 0.006696f
C36 B.n8 VSUBS 0.006696f
C37 B.n9 VSUBS 0.006696f
C38 B.n10 VSUBS 0.006696f
C39 B.n11 VSUBS 0.006696f
C40 B.n12 VSUBS 0.006696f
C41 B.n13 VSUBS 0.006696f
C42 B.n14 VSUBS 0.014904f
C43 B.n15 VSUBS 0.006696f
C44 B.n16 VSUBS 0.006696f
C45 B.n17 VSUBS 0.006696f
C46 B.n18 VSUBS 0.006696f
C47 B.n19 VSUBS 0.006696f
C48 B.n20 VSUBS 0.006696f
C49 B.n21 VSUBS 0.006696f
C50 B.n22 VSUBS 0.006696f
C51 B.n23 VSUBS 0.006696f
C52 B.n24 VSUBS 0.006696f
C53 B.n25 VSUBS 0.006696f
C54 B.n26 VSUBS 0.006696f
C55 B.n27 VSUBS 0.006696f
C56 B.n28 VSUBS 0.006696f
C57 B.n29 VSUBS 0.006696f
C58 B.n30 VSUBS 0.006696f
C59 B.n31 VSUBS 0.006696f
C60 B.n32 VSUBS 0.006696f
C61 B.n33 VSUBS 0.006696f
C62 B.n34 VSUBS 0.006696f
C63 B.n35 VSUBS 0.006696f
C64 B.n36 VSUBS 0.006696f
C65 B.n37 VSUBS 0.006696f
C66 B.n38 VSUBS 0.006696f
C67 B.n39 VSUBS 0.006696f
C68 B.n40 VSUBS 0.006696f
C69 B.n41 VSUBS 0.006696f
C70 B.n42 VSUBS 0.006696f
C71 B.n43 VSUBS 0.006696f
C72 B.n44 VSUBS 0.006696f
C73 B.n45 VSUBS 0.006696f
C74 B.n46 VSUBS 0.006696f
C75 B.n47 VSUBS 0.006696f
C76 B.t4 VSUBS 0.642713f
C77 B.t5 VSUBS 0.66369f
C78 B.t3 VSUBS 2.22179f
C79 B.n48 VSUBS 0.373047f
C80 B.n49 VSUBS 0.0693f
C81 B.n50 VSUBS 0.006696f
C82 B.n51 VSUBS 0.006696f
C83 B.n52 VSUBS 0.006696f
C84 B.n53 VSUBS 0.006696f
C85 B.t1 VSUBS 0.642685f
C86 B.t2 VSUBS 0.663669f
C87 B.t0 VSUBS 2.22179f
C88 B.n54 VSUBS 0.373069f
C89 B.n55 VSUBS 0.069328f
C90 B.n56 VSUBS 0.006696f
C91 B.n57 VSUBS 0.006696f
C92 B.n58 VSUBS 0.006696f
C93 B.n59 VSUBS 0.006696f
C94 B.n60 VSUBS 0.006696f
C95 B.n61 VSUBS 0.006696f
C96 B.n62 VSUBS 0.006696f
C97 B.n63 VSUBS 0.006696f
C98 B.n64 VSUBS 0.006696f
C99 B.n65 VSUBS 0.006696f
C100 B.n66 VSUBS 0.006696f
C101 B.n67 VSUBS 0.006696f
C102 B.n68 VSUBS 0.006696f
C103 B.n69 VSUBS 0.006696f
C104 B.n70 VSUBS 0.006696f
C105 B.n71 VSUBS 0.006696f
C106 B.n72 VSUBS 0.006696f
C107 B.n73 VSUBS 0.006696f
C108 B.n74 VSUBS 0.006696f
C109 B.n75 VSUBS 0.006696f
C110 B.n76 VSUBS 0.006696f
C111 B.n77 VSUBS 0.006696f
C112 B.n78 VSUBS 0.006696f
C113 B.n79 VSUBS 0.006696f
C114 B.n80 VSUBS 0.006696f
C115 B.n81 VSUBS 0.006696f
C116 B.n82 VSUBS 0.006696f
C117 B.n83 VSUBS 0.006696f
C118 B.n84 VSUBS 0.006696f
C119 B.n85 VSUBS 0.006696f
C120 B.n86 VSUBS 0.006696f
C121 B.n87 VSUBS 0.006696f
C122 B.n88 VSUBS 0.014904f
C123 B.n89 VSUBS 0.006696f
C124 B.n90 VSUBS 0.006696f
C125 B.n91 VSUBS 0.006696f
C126 B.n92 VSUBS 0.006696f
C127 B.n93 VSUBS 0.006696f
C128 B.n94 VSUBS 0.006696f
C129 B.n95 VSUBS 0.006696f
C130 B.n96 VSUBS 0.006696f
C131 B.n97 VSUBS 0.006696f
C132 B.n98 VSUBS 0.006696f
C133 B.n99 VSUBS 0.006696f
C134 B.n100 VSUBS 0.006696f
C135 B.n101 VSUBS 0.006696f
C136 B.n102 VSUBS 0.006696f
C137 B.n103 VSUBS 0.006696f
C138 B.n104 VSUBS 0.006696f
C139 B.n105 VSUBS 0.006696f
C140 B.n106 VSUBS 0.006696f
C141 B.n107 VSUBS 0.006696f
C142 B.n108 VSUBS 0.006696f
C143 B.n109 VSUBS 0.006696f
C144 B.n110 VSUBS 0.006696f
C145 B.n111 VSUBS 0.006696f
C146 B.n112 VSUBS 0.006696f
C147 B.n113 VSUBS 0.006696f
C148 B.n114 VSUBS 0.015411f
C149 B.n115 VSUBS 0.006696f
C150 B.n116 VSUBS 0.006696f
C151 B.n117 VSUBS 0.006696f
C152 B.n118 VSUBS 0.006696f
C153 B.n119 VSUBS 0.006696f
C154 B.n120 VSUBS 0.006696f
C155 B.n121 VSUBS 0.006696f
C156 B.n122 VSUBS 0.006696f
C157 B.n123 VSUBS 0.006696f
C158 B.n124 VSUBS 0.006696f
C159 B.n125 VSUBS 0.006696f
C160 B.n126 VSUBS 0.006696f
C161 B.n127 VSUBS 0.006696f
C162 B.n128 VSUBS 0.006696f
C163 B.n129 VSUBS 0.006696f
C164 B.n130 VSUBS 0.006696f
C165 B.n131 VSUBS 0.006696f
C166 B.n132 VSUBS 0.006696f
C167 B.n133 VSUBS 0.006696f
C168 B.n134 VSUBS 0.006696f
C169 B.n135 VSUBS 0.006696f
C170 B.n136 VSUBS 0.006696f
C171 B.n137 VSUBS 0.006696f
C172 B.n138 VSUBS 0.006696f
C173 B.n139 VSUBS 0.006696f
C174 B.n140 VSUBS 0.006696f
C175 B.n141 VSUBS 0.006696f
C176 B.n142 VSUBS 0.006696f
C177 B.n143 VSUBS 0.006696f
C178 B.n144 VSUBS 0.006696f
C179 B.n145 VSUBS 0.006696f
C180 B.n146 VSUBS 0.004628f
C181 B.n147 VSUBS 0.006696f
C182 B.n148 VSUBS 0.006696f
C183 B.n149 VSUBS 0.006696f
C184 B.n150 VSUBS 0.006696f
C185 B.n151 VSUBS 0.006696f
C186 B.t8 VSUBS 0.642713f
C187 B.t7 VSUBS 0.66369f
C188 B.t6 VSUBS 2.22179f
C189 B.n152 VSUBS 0.373047f
C190 B.n153 VSUBS 0.0693f
C191 B.n154 VSUBS 0.006696f
C192 B.n155 VSUBS 0.006696f
C193 B.n156 VSUBS 0.006696f
C194 B.n157 VSUBS 0.006696f
C195 B.n158 VSUBS 0.006696f
C196 B.n159 VSUBS 0.006696f
C197 B.n160 VSUBS 0.006696f
C198 B.n161 VSUBS 0.006696f
C199 B.n162 VSUBS 0.006696f
C200 B.n163 VSUBS 0.006696f
C201 B.n164 VSUBS 0.006696f
C202 B.n165 VSUBS 0.006696f
C203 B.n166 VSUBS 0.006696f
C204 B.n167 VSUBS 0.006696f
C205 B.n168 VSUBS 0.006696f
C206 B.n169 VSUBS 0.006696f
C207 B.n170 VSUBS 0.006696f
C208 B.n171 VSUBS 0.006696f
C209 B.n172 VSUBS 0.006696f
C210 B.n173 VSUBS 0.006696f
C211 B.n174 VSUBS 0.006696f
C212 B.n175 VSUBS 0.006696f
C213 B.n176 VSUBS 0.006696f
C214 B.n177 VSUBS 0.006696f
C215 B.n178 VSUBS 0.006696f
C216 B.n179 VSUBS 0.006696f
C217 B.n180 VSUBS 0.006696f
C218 B.n181 VSUBS 0.006696f
C219 B.n182 VSUBS 0.006696f
C220 B.n183 VSUBS 0.006696f
C221 B.n184 VSUBS 0.006696f
C222 B.n185 VSUBS 0.016211f
C223 B.n186 VSUBS 0.006696f
C224 B.n187 VSUBS 0.006696f
C225 B.n188 VSUBS 0.006696f
C226 B.n189 VSUBS 0.006696f
C227 B.n190 VSUBS 0.006696f
C228 B.n191 VSUBS 0.006696f
C229 B.n192 VSUBS 0.006696f
C230 B.n193 VSUBS 0.006696f
C231 B.n194 VSUBS 0.006696f
C232 B.n195 VSUBS 0.006696f
C233 B.n196 VSUBS 0.006696f
C234 B.n197 VSUBS 0.006696f
C235 B.n198 VSUBS 0.006696f
C236 B.n199 VSUBS 0.006696f
C237 B.n200 VSUBS 0.006696f
C238 B.n201 VSUBS 0.006696f
C239 B.n202 VSUBS 0.006696f
C240 B.n203 VSUBS 0.006696f
C241 B.n204 VSUBS 0.006696f
C242 B.n205 VSUBS 0.006696f
C243 B.n206 VSUBS 0.006696f
C244 B.n207 VSUBS 0.006696f
C245 B.n208 VSUBS 0.006696f
C246 B.n209 VSUBS 0.006696f
C247 B.n210 VSUBS 0.006696f
C248 B.n211 VSUBS 0.006696f
C249 B.n212 VSUBS 0.006696f
C250 B.n213 VSUBS 0.006696f
C251 B.n214 VSUBS 0.006696f
C252 B.n215 VSUBS 0.006696f
C253 B.n216 VSUBS 0.006696f
C254 B.n217 VSUBS 0.006696f
C255 B.n218 VSUBS 0.006696f
C256 B.n219 VSUBS 0.006696f
C257 B.n220 VSUBS 0.006696f
C258 B.n221 VSUBS 0.006696f
C259 B.n222 VSUBS 0.006696f
C260 B.n223 VSUBS 0.006696f
C261 B.n224 VSUBS 0.006696f
C262 B.n225 VSUBS 0.006696f
C263 B.n226 VSUBS 0.006696f
C264 B.n227 VSUBS 0.006696f
C265 B.n228 VSUBS 0.006696f
C266 B.n229 VSUBS 0.006696f
C267 B.n230 VSUBS 0.006696f
C268 B.n231 VSUBS 0.006696f
C269 B.n232 VSUBS 0.014904f
C270 B.n233 VSUBS 0.014904f
C271 B.n234 VSUBS 0.016211f
C272 B.n235 VSUBS 0.006696f
C273 B.n236 VSUBS 0.006696f
C274 B.n237 VSUBS 0.006696f
C275 B.n238 VSUBS 0.006696f
C276 B.n239 VSUBS 0.006696f
C277 B.n240 VSUBS 0.006696f
C278 B.n241 VSUBS 0.006696f
C279 B.n242 VSUBS 0.006696f
C280 B.n243 VSUBS 0.006696f
C281 B.n244 VSUBS 0.006696f
C282 B.n245 VSUBS 0.006696f
C283 B.n246 VSUBS 0.006696f
C284 B.n247 VSUBS 0.006696f
C285 B.n248 VSUBS 0.006696f
C286 B.n249 VSUBS 0.006696f
C287 B.n250 VSUBS 0.006696f
C288 B.n251 VSUBS 0.006696f
C289 B.n252 VSUBS 0.006696f
C290 B.n253 VSUBS 0.006696f
C291 B.n254 VSUBS 0.006696f
C292 B.n255 VSUBS 0.006696f
C293 B.n256 VSUBS 0.006696f
C294 B.n257 VSUBS 0.006696f
C295 B.n258 VSUBS 0.006696f
C296 B.n259 VSUBS 0.006696f
C297 B.n260 VSUBS 0.006696f
C298 B.n261 VSUBS 0.006696f
C299 B.n262 VSUBS 0.006696f
C300 B.n263 VSUBS 0.006696f
C301 B.n264 VSUBS 0.006696f
C302 B.n265 VSUBS 0.006696f
C303 B.n266 VSUBS 0.006696f
C304 B.n267 VSUBS 0.006696f
C305 B.n268 VSUBS 0.006696f
C306 B.n269 VSUBS 0.006696f
C307 B.n270 VSUBS 0.006696f
C308 B.n271 VSUBS 0.006696f
C309 B.n272 VSUBS 0.006696f
C310 B.n273 VSUBS 0.006696f
C311 B.n274 VSUBS 0.006696f
C312 B.n275 VSUBS 0.006696f
C313 B.n276 VSUBS 0.006696f
C314 B.n277 VSUBS 0.006696f
C315 B.n278 VSUBS 0.006696f
C316 B.n279 VSUBS 0.006696f
C317 B.n280 VSUBS 0.006696f
C318 B.n281 VSUBS 0.006696f
C319 B.n282 VSUBS 0.006696f
C320 B.n283 VSUBS 0.006696f
C321 B.n284 VSUBS 0.006696f
C322 B.n285 VSUBS 0.006696f
C323 B.n286 VSUBS 0.006696f
C324 B.n287 VSUBS 0.006696f
C325 B.n288 VSUBS 0.006696f
C326 B.n289 VSUBS 0.006696f
C327 B.n290 VSUBS 0.006696f
C328 B.n291 VSUBS 0.006696f
C329 B.n292 VSUBS 0.006696f
C330 B.n293 VSUBS 0.006696f
C331 B.n294 VSUBS 0.006696f
C332 B.n295 VSUBS 0.006696f
C333 B.n296 VSUBS 0.006696f
C334 B.n297 VSUBS 0.006696f
C335 B.n298 VSUBS 0.006696f
C336 B.n299 VSUBS 0.006696f
C337 B.n300 VSUBS 0.006696f
C338 B.n301 VSUBS 0.006696f
C339 B.n302 VSUBS 0.006696f
C340 B.n303 VSUBS 0.006696f
C341 B.n304 VSUBS 0.006696f
C342 B.n305 VSUBS 0.006696f
C343 B.n306 VSUBS 0.006696f
C344 B.n307 VSUBS 0.006696f
C345 B.n308 VSUBS 0.006696f
C346 B.n309 VSUBS 0.006696f
C347 B.n310 VSUBS 0.006696f
C348 B.n311 VSUBS 0.006696f
C349 B.n312 VSUBS 0.006696f
C350 B.n313 VSUBS 0.006696f
C351 B.n314 VSUBS 0.006696f
C352 B.n315 VSUBS 0.006696f
C353 B.n316 VSUBS 0.006696f
C354 B.n317 VSUBS 0.006696f
C355 B.n318 VSUBS 0.006696f
C356 B.n319 VSUBS 0.006696f
C357 B.n320 VSUBS 0.006696f
C358 B.n321 VSUBS 0.006696f
C359 B.n322 VSUBS 0.006696f
C360 B.n323 VSUBS 0.006696f
C361 B.n324 VSUBS 0.006696f
C362 B.n325 VSUBS 0.006696f
C363 B.n326 VSUBS 0.006696f
C364 B.n327 VSUBS 0.006696f
C365 B.n328 VSUBS 0.006696f
C366 B.n329 VSUBS 0.006696f
C367 B.n330 VSUBS 0.004628f
C368 B.n331 VSUBS 0.015513f
C369 B.n332 VSUBS 0.005415f
C370 B.n333 VSUBS 0.006696f
C371 B.n334 VSUBS 0.006696f
C372 B.n335 VSUBS 0.006696f
C373 B.n336 VSUBS 0.006696f
C374 B.n337 VSUBS 0.006696f
C375 B.n338 VSUBS 0.006696f
C376 B.n339 VSUBS 0.006696f
C377 B.n340 VSUBS 0.006696f
C378 B.n341 VSUBS 0.006696f
C379 B.n342 VSUBS 0.006696f
C380 B.n343 VSUBS 0.006696f
C381 B.t11 VSUBS 0.642685f
C382 B.t10 VSUBS 0.663669f
C383 B.t9 VSUBS 2.22179f
C384 B.n344 VSUBS 0.373069f
C385 B.n345 VSUBS 0.069328f
C386 B.n346 VSUBS 0.015513f
C387 B.n347 VSUBS 0.005415f
C388 B.n348 VSUBS 0.006696f
C389 B.n349 VSUBS 0.006696f
C390 B.n350 VSUBS 0.006696f
C391 B.n351 VSUBS 0.006696f
C392 B.n352 VSUBS 0.006696f
C393 B.n353 VSUBS 0.006696f
C394 B.n354 VSUBS 0.006696f
C395 B.n355 VSUBS 0.006696f
C396 B.n356 VSUBS 0.006696f
C397 B.n357 VSUBS 0.006696f
C398 B.n358 VSUBS 0.006696f
C399 B.n359 VSUBS 0.006696f
C400 B.n360 VSUBS 0.006696f
C401 B.n361 VSUBS 0.006696f
C402 B.n362 VSUBS 0.006696f
C403 B.n363 VSUBS 0.006696f
C404 B.n364 VSUBS 0.006696f
C405 B.n365 VSUBS 0.006696f
C406 B.n366 VSUBS 0.006696f
C407 B.n367 VSUBS 0.006696f
C408 B.n368 VSUBS 0.006696f
C409 B.n369 VSUBS 0.006696f
C410 B.n370 VSUBS 0.006696f
C411 B.n371 VSUBS 0.006696f
C412 B.n372 VSUBS 0.006696f
C413 B.n373 VSUBS 0.006696f
C414 B.n374 VSUBS 0.006696f
C415 B.n375 VSUBS 0.006696f
C416 B.n376 VSUBS 0.006696f
C417 B.n377 VSUBS 0.006696f
C418 B.n378 VSUBS 0.006696f
C419 B.n379 VSUBS 0.006696f
C420 B.n380 VSUBS 0.006696f
C421 B.n381 VSUBS 0.006696f
C422 B.n382 VSUBS 0.006696f
C423 B.n383 VSUBS 0.006696f
C424 B.n384 VSUBS 0.006696f
C425 B.n385 VSUBS 0.006696f
C426 B.n386 VSUBS 0.006696f
C427 B.n387 VSUBS 0.006696f
C428 B.n388 VSUBS 0.006696f
C429 B.n389 VSUBS 0.006696f
C430 B.n390 VSUBS 0.006696f
C431 B.n391 VSUBS 0.006696f
C432 B.n392 VSUBS 0.006696f
C433 B.n393 VSUBS 0.006696f
C434 B.n394 VSUBS 0.006696f
C435 B.n395 VSUBS 0.006696f
C436 B.n396 VSUBS 0.006696f
C437 B.n397 VSUBS 0.006696f
C438 B.n398 VSUBS 0.006696f
C439 B.n399 VSUBS 0.006696f
C440 B.n400 VSUBS 0.006696f
C441 B.n401 VSUBS 0.006696f
C442 B.n402 VSUBS 0.006696f
C443 B.n403 VSUBS 0.006696f
C444 B.n404 VSUBS 0.006696f
C445 B.n405 VSUBS 0.006696f
C446 B.n406 VSUBS 0.006696f
C447 B.n407 VSUBS 0.006696f
C448 B.n408 VSUBS 0.006696f
C449 B.n409 VSUBS 0.006696f
C450 B.n410 VSUBS 0.006696f
C451 B.n411 VSUBS 0.006696f
C452 B.n412 VSUBS 0.006696f
C453 B.n413 VSUBS 0.006696f
C454 B.n414 VSUBS 0.006696f
C455 B.n415 VSUBS 0.006696f
C456 B.n416 VSUBS 0.006696f
C457 B.n417 VSUBS 0.006696f
C458 B.n418 VSUBS 0.006696f
C459 B.n419 VSUBS 0.006696f
C460 B.n420 VSUBS 0.006696f
C461 B.n421 VSUBS 0.006696f
C462 B.n422 VSUBS 0.006696f
C463 B.n423 VSUBS 0.006696f
C464 B.n424 VSUBS 0.006696f
C465 B.n425 VSUBS 0.006696f
C466 B.n426 VSUBS 0.006696f
C467 B.n427 VSUBS 0.006696f
C468 B.n428 VSUBS 0.006696f
C469 B.n429 VSUBS 0.006696f
C470 B.n430 VSUBS 0.006696f
C471 B.n431 VSUBS 0.006696f
C472 B.n432 VSUBS 0.006696f
C473 B.n433 VSUBS 0.006696f
C474 B.n434 VSUBS 0.006696f
C475 B.n435 VSUBS 0.006696f
C476 B.n436 VSUBS 0.006696f
C477 B.n437 VSUBS 0.006696f
C478 B.n438 VSUBS 0.006696f
C479 B.n439 VSUBS 0.006696f
C480 B.n440 VSUBS 0.006696f
C481 B.n441 VSUBS 0.006696f
C482 B.n442 VSUBS 0.006696f
C483 B.n443 VSUBS 0.006696f
C484 B.n444 VSUBS 0.006696f
C485 B.n445 VSUBS 0.016211f
C486 B.n446 VSUBS 0.014904f
C487 B.n447 VSUBS 0.015703f
C488 B.n448 VSUBS 0.006696f
C489 B.n449 VSUBS 0.006696f
C490 B.n450 VSUBS 0.006696f
C491 B.n451 VSUBS 0.006696f
C492 B.n452 VSUBS 0.006696f
C493 B.n453 VSUBS 0.006696f
C494 B.n454 VSUBS 0.006696f
C495 B.n455 VSUBS 0.006696f
C496 B.n456 VSUBS 0.006696f
C497 B.n457 VSUBS 0.006696f
C498 B.n458 VSUBS 0.006696f
C499 B.n459 VSUBS 0.006696f
C500 B.n460 VSUBS 0.006696f
C501 B.n461 VSUBS 0.006696f
C502 B.n462 VSUBS 0.006696f
C503 B.n463 VSUBS 0.006696f
C504 B.n464 VSUBS 0.006696f
C505 B.n465 VSUBS 0.006696f
C506 B.n466 VSUBS 0.006696f
C507 B.n467 VSUBS 0.006696f
C508 B.n468 VSUBS 0.006696f
C509 B.n469 VSUBS 0.006696f
C510 B.n470 VSUBS 0.006696f
C511 B.n471 VSUBS 0.006696f
C512 B.n472 VSUBS 0.006696f
C513 B.n473 VSUBS 0.006696f
C514 B.n474 VSUBS 0.006696f
C515 B.n475 VSUBS 0.006696f
C516 B.n476 VSUBS 0.006696f
C517 B.n477 VSUBS 0.006696f
C518 B.n478 VSUBS 0.006696f
C519 B.n479 VSUBS 0.006696f
C520 B.n480 VSUBS 0.006696f
C521 B.n481 VSUBS 0.006696f
C522 B.n482 VSUBS 0.006696f
C523 B.n483 VSUBS 0.006696f
C524 B.n484 VSUBS 0.006696f
C525 B.n485 VSUBS 0.006696f
C526 B.n486 VSUBS 0.006696f
C527 B.n487 VSUBS 0.006696f
C528 B.n488 VSUBS 0.006696f
C529 B.n489 VSUBS 0.006696f
C530 B.n490 VSUBS 0.006696f
C531 B.n491 VSUBS 0.006696f
C532 B.n492 VSUBS 0.006696f
C533 B.n493 VSUBS 0.006696f
C534 B.n494 VSUBS 0.006696f
C535 B.n495 VSUBS 0.006696f
C536 B.n496 VSUBS 0.006696f
C537 B.n497 VSUBS 0.006696f
C538 B.n498 VSUBS 0.006696f
C539 B.n499 VSUBS 0.006696f
C540 B.n500 VSUBS 0.006696f
C541 B.n501 VSUBS 0.006696f
C542 B.n502 VSUBS 0.006696f
C543 B.n503 VSUBS 0.006696f
C544 B.n504 VSUBS 0.006696f
C545 B.n505 VSUBS 0.006696f
C546 B.n506 VSUBS 0.006696f
C547 B.n507 VSUBS 0.006696f
C548 B.n508 VSUBS 0.006696f
C549 B.n509 VSUBS 0.006696f
C550 B.n510 VSUBS 0.006696f
C551 B.n511 VSUBS 0.006696f
C552 B.n512 VSUBS 0.006696f
C553 B.n513 VSUBS 0.006696f
C554 B.n514 VSUBS 0.006696f
C555 B.n515 VSUBS 0.006696f
C556 B.n516 VSUBS 0.006696f
C557 B.n517 VSUBS 0.006696f
C558 B.n518 VSUBS 0.006696f
C559 B.n519 VSUBS 0.006696f
C560 B.n520 VSUBS 0.006696f
C561 B.n521 VSUBS 0.006696f
C562 B.n522 VSUBS 0.006696f
C563 B.n523 VSUBS 0.014904f
C564 B.n524 VSUBS 0.016211f
C565 B.n525 VSUBS 0.016211f
C566 B.n526 VSUBS 0.006696f
C567 B.n527 VSUBS 0.006696f
C568 B.n528 VSUBS 0.006696f
C569 B.n529 VSUBS 0.006696f
C570 B.n530 VSUBS 0.006696f
C571 B.n531 VSUBS 0.006696f
C572 B.n532 VSUBS 0.006696f
C573 B.n533 VSUBS 0.006696f
C574 B.n534 VSUBS 0.006696f
C575 B.n535 VSUBS 0.006696f
C576 B.n536 VSUBS 0.006696f
C577 B.n537 VSUBS 0.006696f
C578 B.n538 VSUBS 0.006696f
C579 B.n539 VSUBS 0.006696f
C580 B.n540 VSUBS 0.006696f
C581 B.n541 VSUBS 0.006696f
C582 B.n542 VSUBS 0.006696f
C583 B.n543 VSUBS 0.006696f
C584 B.n544 VSUBS 0.006696f
C585 B.n545 VSUBS 0.006696f
C586 B.n546 VSUBS 0.006696f
C587 B.n547 VSUBS 0.006696f
C588 B.n548 VSUBS 0.006696f
C589 B.n549 VSUBS 0.006696f
C590 B.n550 VSUBS 0.006696f
C591 B.n551 VSUBS 0.006696f
C592 B.n552 VSUBS 0.006696f
C593 B.n553 VSUBS 0.006696f
C594 B.n554 VSUBS 0.006696f
C595 B.n555 VSUBS 0.006696f
C596 B.n556 VSUBS 0.006696f
C597 B.n557 VSUBS 0.006696f
C598 B.n558 VSUBS 0.006696f
C599 B.n559 VSUBS 0.006696f
C600 B.n560 VSUBS 0.006696f
C601 B.n561 VSUBS 0.006696f
C602 B.n562 VSUBS 0.006696f
C603 B.n563 VSUBS 0.006696f
C604 B.n564 VSUBS 0.006696f
C605 B.n565 VSUBS 0.006696f
C606 B.n566 VSUBS 0.006696f
C607 B.n567 VSUBS 0.006696f
C608 B.n568 VSUBS 0.006696f
C609 B.n569 VSUBS 0.006696f
C610 B.n570 VSUBS 0.006696f
C611 B.n571 VSUBS 0.006696f
C612 B.n572 VSUBS 0.006696f
C613 B.n573 VSUBS 0.006696f
C614 B.n574 VSUBS 0.006696f
C615 B.n575 VSUBS 0.006696f
C616 B.n576 VSUBS 0.006696f
C617 B.n577 VSUBS 0.006696f
C618 B.n578 VSUBS 0.006696f
C619 B.n579 VSUBS 0.006696f
C620 B.n580 VSUBS 0.006696f
C621 B.n581 VSUBS 0.006696f
C622 B.n582 VSUBS 0.006696f
C623 B.n583 VSUBS 0.006696f
C624 B.n584 VSUBS 0.006696f
C625 B.n585 VSUBS 0.006696f
C626 B.n586 VSUBS 0.006696f
C627 B.n587 VSUBS 0.006696f
C628 B.n588 VSUBS 0.006696f
C629 B.n589 VSUBS 0.006696f
C630 B.n590 VSUBS 0.006696f
C631 B.n591 VSUBS 0.006696f
C632 B.n592 VSUBS 0.006696f
C633 B.n593 VSUBS 0.006696f
C634 B.n594 VSUBS 0.006696f
C635 B.n595 VSUBS 0.006696f
C636 B.n596 VSUBS 0.006696f
C637 B.n597 VSUBS 0.006696f
C638 B.n598 VSUBS 0.006696f
C639 B.n599 VSUBS 0.006696f
C640 B.n600 VSUBS 0.006696f
C641 B.n601 VSUBS 0.006696f
C642 B.n602 VSUBS 0.006696f
C643 B.n603 VSUBS 0.006696f
C644 B.n604 VSUBS 0.006696f
C645 B.n605 VSUBS 0.006696f
C646 B.n606 VSUBS 0.006696f
C647 B.n607 VSUBS 0.006696f
C648 B.n608 VSUBS 0.006696f
C649 B.n609 VSUBS 0.006696f
C650 B.n610 VSUBS 0.006696f
C651 B.n611 VSUBS 0.006696f
C652 B.n612 VSUBS 0.006696f
C653 B.n613 VSUBS 0.006696f
C654 B.n614 VSUBS 0.006696f
C655 B.n615 VSUBS 0.006696f
C656 B.n616 VSUBS 0.006696f
C657 B.n617 VSUBS 0.006696f
C658 B.n618 VSUBS 0.006696f
C659 B.n619 VSUBS 0.006696f
C660 B.n620 VSUBS 0.006696f
C661 B.n621 VSUBS 0.004628f
C662 B.n622 VSUBS 0.015513f
C663 B.n623 VSUBS 0.005415f
C664 B.n624 VSUBS 0.006696f
C665 B.n625 VSUBS 0.006696f
C666 B.n626 VSUBS 0.006696f
C667 B.n627 VSUBS 0.006696f
C668 B.n628 VSUBS 0.006696f
C669 B.n629 VSUBS 0.006696f
C670 B.n630 VSUBS 0.006696f
C671 B.n631 VSUBS 0.006696f
C672 B.n632 VSUBS 0.006696f
C673 B.n633 VSUBS 0.006696f
C674 B.n634 VSUBS 0.006696f
C675 B.n635 VSUBS 0.005415f
C676 B.n636 VSUBS 0.015513f
C677 B.n637 VSUBS 0.004628f
C678 B.n638 VSUBS 0.006696f
C679 B.n639 VSUBS 0.006696f
C680 B.n640 VSUBS 0.006696f
C681 B.n641 VSUBS 0.006696f
C682 B.n642 VSUBS 0.006696f
C683 B.n643 VSUBS 0.006696f
C684 B.n644 VSUBS 0.006696f
C685 B.n645 VSUBS 0.006696f
C686 B.n646 VSUBS 0.006696f
C687 B.n647 VSUBS 0.006696f
C688 B.n648 VSUBS 0.006696f
C689 B.n649 VSUBS 0.006696f
C690 B.n650 VSUBS 0.006696f
C691 B.n651 VSUBS 0.006696f
C692 B.n652 VSUBS 0.006696f
C693 B.n653 VSUBS 0.006696f
C694 B.n654 VSUBS 0.006696f
C695 B.n655 VSUBS 0.006696f
C696 B.n656 VSUBS 0.006696f
C697 B.n657 VSUBS 0.006696f
C698 B.n658 VSUBS 0.006696f
C699 B.n659 VSUBS 0.006696f
C700 B.n660 VSUBS 0.006696f
C701 B.n661 VSUBS 0.006696f
C702 B.n662 VSUBS 0.006696f
C703 B.n663 VSUBS 0.006696f
C704 B.n664 VSUBS 0.006696f
C705 B.n665 VSUBS 0.006696f
C706 B.n666 VSUBS 0.006696f
C707 B.n667 VSUBS 0.006696f
C708 B.n668 VSUBS 0.006696f
C709 B.n669 VSUBS 0.006696f
C710 B.n670 VSUBS 0.006696f
C711 B.n671 VSUBS 0.006696f
C712 B.n672 VSUBS 0.006696f
C713 B.n673 VSUBS 0.006696f
C714 B.n674 VSUBS 0.006696f
C715 B.n675 VSUBS 0.006696f
C716 B.n676 VSUBS 0.006696f
C717 B.n677 VSUBS 0.006696f
C718 B.n678 VSUBS 0.006696f
C719 B.n679 VSUBS 0.006696f
C720 B.n680 VSUBS 0.006696f
C721 B.n681 VSUBS 0.006696f
C722 B.n682 VSUBS 0.006696f
C723 B.n683 VSUBS 0.006696f
C724 B.n684 VSUBS 0.006696f
C725 B.n685 VSUBS 0.006696f
C726 B.n686 VSUBS 0.006696f
C727 B.n687 VSUBS 0.006696f
C728 B.n688 VSUBS 0.006696f
C729 B.n689 VSUBS 0.006696f
C730 B.n690 VSUBS 0.006696f
C731 B.n691 VSUBS 0.006696f
C732 B.n692 VSUBS 0.006696f
C733 B.n693 VSUBS 0.006696f
C734 B.n694 VSUBS 0.006696f
C735 B.n695 VSUBS 0.006696f
C736 B.n696 VSUBS 0.006696f
C737 B.n697 VSUBS 0.006696f
C738 B.n698 VSUBS 0.006696f
C739 B.n699 VSUBS 0.006696f
C740 B.n700 VSUBS 0.006696f
C741 B.n701 VSUBS 0.006696f
C742 B.n702 VSUBS 0.006696f
C743 B.n703 VSUBS 0.006696f
C744 B.n704 VSUBS 0.006696f
C745 B.n705 VSUBS 0.006696f
C746 B.n706 VSUBS 0.006696f
C747 B.n707 VSUBS 0.006696f
C748 B.n708 VSUBS 0.006696f
C749 B.n709 VSUBS 0.006696f
C750 B.n710 VSUBS 0.006696f
C751 B.n711 VSUBS 0.006696f
C752 B.n712 VSUBS 0.006696f
C753 B.n713 VSUBS 0.006696f
C754 B.n714 VSUBS 0.006696f
C755 B.n715 VSUBS 0.006696f
C756 B.n716 VSUBS 0.006696f
C757 B.n717 VSUBS 0.006696f
C758 B.n718 VSUBS 0.006696f
C759 B.n719 VSUBS 0.006696f
C760 B.n720 VSUBS 0.006696f
C761 B.n721 VSUBS 0.006696f
C762 B.n722 VSUBS 0.006696f
C763 B.n723 VSUBS 0.006696f
C764 B.n724 VSUBS 0.006696f
C765 B.n725 VSUBS 0.006696f
C766 B.n726 VSUBS 0.006696f
C767 B.n727 VSUBS 0.006696f
C768 B.n728 VSUBS 0.006696f
C769 B.n729 VSUBS 0.006696f
C770 B.n730 VSUBS 0.006696f
C771 B.n731 VSUBS 0.006696f
C772 B.n732 VSUBS 0.006696f
C773 B.n733 VSUBS 0.016211f
C774 B.n734 VSUBS 0.016211f
C775 B.n735 VSUBS 0.014904f
C776 B.n736 VSUBS 0.006696f
C777 B.n737 VSUBS 0.006696f
C778 B.n738 VSUBS 0.006696f
C779 B.n739 VSUBS 0.006696f
C780 B.n740 VSUBS 0.006696f
C781 B.n741 VSUBS 0.006696f
C782 B.n742 VSUBS 0.006696f
C783 B.n743 VSUBS 0.006696f
C784 B.n744 VSUBS 0.006696f
C785 B.n745 VSUBS 0.006696f
C786 B.n746 VSUBS 0.006696f
C787 B.n747 VSUBS 0.006696f
C788 B.n748 VSUBS 0.006696f
C789 B.n749 VSUBS 0.006696f
C790 B.n750 VSUBS 0.006696f
C791 B.n751 VSUBS 0.006696f
C792 B.n752 VSUBS 0.006696f
C793 B.n753 VSUBS 0.006696f
C794 B.n754 VSUBS 0.006696f
C795 B.n755 VSUBS 0.006696f
C796 B.n756 VSUBS 0.006696f
C797 B.n757 VSUBS 0.006696f
C798 B.n758 VSUBS 0.006696f
C799 B.n759 VSUBS 0.006696f
C800 B.n760 VSUBS 0.006696f
C801 B.n761 VSUBS 0.006696f
C802 B.n762 VSUBS 0.006696f
C803 B.n763 VSUBS 0.006696f
C804 B.n764 VSUBS 0.006696f
C805 B.n765 VSUBS 0.006696f
C806 B.n766 VSUBS 0.006696f
C807 B.n767 VSUBS 0.006696f
C808 B.n768 VSUBS 0.006696f
C809 B.n769 VSUBS 0.006696f
C810 B.n770 VSUBS 0.006696f
C811 B.n771 VSUBS 0.008737f
C812 B.n772 VSUBS 0.009307f
C813 B.n773 VSUBS 0.018509f
C814 VDD1.t1 VSUBS 4.74441f
C815 VDD1.t0 VSUBS 5.90299f
C816 VP.t1 VSUBS 5.53448f
C817 VP.t0 VSUBS 6.246161f
C818 VP.n0 VSUBS 6.82602f
C819 VDD2.t1 VSUBS 5.92047f
C820 VDD2.t0 VSUBS 4.79666f
C821 VDD2.n0 VSUBS 5.50199f
C822 VTAIL.t1 VSUBS 4.56545f
C823 VTAIL.n0 VSUBS 3.27259f
C824 VTAIL.t2 VSUBS 4.56545f
C825 VTAIL.n1 VSUBS 3.32519f
C826 VTAIL.t0 VSUBS 4.56545f
C827 VTAIL.n2 VSUBS 3.0939f
C828 VTAIL.t3 VSUBS 4.56545f
C829 VTAIL.n3 VSUBS 2.9887f
C830 VN.t0 VSUBS 5.40511f
C831 VN.t1 VSUBS 6.09769f
.ends

