* NGSPICE file created from diff_pair_sample_0424.ext - technology: sky130A

.subckt diff_pair_sample_0424 VTAIL VN VP B VDD2 VDD1
X0 B.t14 B.t12 B.t13 B.t2 sky130_fd_pr__nfet_01v8 ad=5.3235 pd=28.08 as=0 ps=0 w=13.65 l=3.48
X1 B.t11 B.t9 B.t10 B.t6 sky130_fd_pr__nfet_01v8 ad=5.3235 pd=28.08 as=0 ps=0 w=13.65 l=3.48
X2 B.t8 B.t5 B.t7 B.t6 sky130_fd_pr__nfet_01v8 ad=5.3235 pd=28.08 as=0 ps=0 w=13.65 l=3.48
X3 B.t4 B.t1 B.t3 B.t2 sky130_fd_pr__nfet_01v8 ad=5.3235 pd=28.08 as=0 ps=0 w=13.65 l=3.48
X4 VDD2.t1 VN.t0 VTAIL.t2 B.t0 sky130_fd_pr__nfet_01v8 ad=5.3235 pd=28.08 as=5.3235 ps=28.08 w=13.65 l=3.48
X5 VDD1.t1 VP.t0 VTAIL.t1 B.t15 sky130_fd_pr__nfet_01v8 ad=5.3235 pd=28.08 as=5.3235 ps=28.08 w=13.65 l=3.48
X6 VDD1.t0 VP.t1 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=5.3235 pd=28.08 as=5.3235 ps=28.08 w=13.65 l=3.48
X7 VDD2.t0 VN.t1 VTAIL.t3 B.t15 sky130_fd_pr__nfet_01v8 ad=5.3235 pd=28.08 as=5.3235 ps=28.08 w=13.65 l=3.48
R0 B.n566 B.n565 585
R1 B.n567 B.n115 585
R2 B.n569 B.n568 585
R3 B.n571 B.n114 585
R4 B.n574 B.n573 585
R5 B.n575 B.n113 585
R6 B.n577 B.n576 585
R7 B.n579 B.n112 585
R8 B.n582 B.n581 585
R9 B.n583 B.n111 585
R10 B.n585 B.n584 585
R11 B.n587 B.n110 585
R12 B.n590 B.n589 585
R13 B.n591 B.n109 585
R14 B.n593 B.n592 585
R15 B.n595 B.n108 585
R16 B.n598 B.n597 585
R17 B.n599 B.n107 585
R18 B.n601 B.n600 585
R19 B.n603 B.n106 585
R20 B.n606 B.n605 585
R21 B.n607 B.n105 585
R22 B.n609 B.n608 585
R23 B.n611 B.n104 585
R24 B.n614 B.n613 585
R25 B.n615 B.n103 585
R26 B.n617 B.n616 585
R27 B.n619 B.n102 585
R28 B.n622 B.n621 585
R29 B.n623 B.n101 585
R30 B.n625 B.n624 585
R31 B.n627 B.n100 585
R32 B.n630 B.n629 585
R33 B.n631 B.n99 585
R34 B.n633 B.n632 585
R35 B.n635 B.n98 585
R36 B.n638 B.n637 585
R37 B.n639 B.n97 585
R38 B.n641 B.n640 585
R39 B.n643 B.n96 585
R40 B.n646 B.n645 585
R41 B.n647 B.n95 585
R42 B.n649 B.n648 585
R43 B.n651 B.n94 585
R44 B.n653 B.n652 585
R45 B.n655 B.n654 585
R46 B.n658 B.n657 585
R47 B.n659 B.n89 585
R48 B.n661 B.n660 585
R49 B.n663 B.n88 585
R50 B.n666 B.n665 585
R51 B.n667 B.n87 585
R52 B.n669 B.n668 585
R53 B.n671 B.n86 585
R54 B.n673 B.n672 585
R55 B.n675 B.n674 585
R56 B.n678 B.n677 585
R57 B.n679 B.n81 585
R58 B.n681 B.n680 585
R59 B.n683 B.n80 585
R60 B.n686 B.n685 585
R61 B.n687 B.n79 585
R62 B.n689 B.n688 585
R63 B.n691 B.n78 585
R64 B.n694 B.n693 585
R65 B.n695 B.n77 585
R66 B.n697 B.n696 585
R67 B.n699 B.n76 585
R68 B.n702 B.n701 585
R69 B.n703 B.n75 585
R70 B.n705 B.n704 585
R71 B.n707 B.n74 585
R72 B.n710 B.n709 585
R73 B.n711 B.n73 585
R74 B.n713 B.n712 585
R75 B.n715 B.n72 585
R76 B.n718 B.n717 585
R77 B.n719 B.n71 585
R78 B.n721 B.n720 585
R79 B.n723 B.n70 585
R80 B.n726 B.n725 585
R81 B.n727 B.n69 585
R82 B.n729 B.n728 585
R83 B.n731 B.n68 585
R84 B.n734 B.n733 585
R85 B.n735 B.n67 585
R86 B.n737 B.n736 585
R87 B.n739 B.n66 585
R88 B.n742 B.n741 585
R89 B.n743 B.n65 585
R90 B.n745 B.n744 585
R91 B.n747 B.n64 585
R92 B.n750 B.n749 585
R93 B.n751 B.n63 585
R94 B.n753 B.n752 585
R95 B.n755 B.n62 585
R96 B.n758 B.n757 585
R97 B.n759 B.n61 585
R98 B.n761 B.n760 585
R99 B.n763 B.n60 585
R100 B.n766 B.n765 585
R101 B.n767 B.n59 585
R102 B.n563 B.n57 585
R103 B.n770 B.n57 585
R104 B.n562 B.n56 585
R105 B.n771 B.n56 585
R106 B.n561 B.n55 585
R107 B.n772 B.n55 585
R108 B.n560 B.n559 585
R109 B.n559 B.n51 585
R110 B.n558 B.n50 585
R111 B.n778 B.n50 585
R112 B.n557 B.n49 585
R113 B.n779 B.n49 585
R114 B.n556 B.n48 585
R115 B.n780 B.n48 585
R116 B.n555 B.n554 585
R117 B.n554 B.n44 585
R118 B.n553 B.n43 585
R119 B.n786 B.n43 585
R120 B.n552 B.n42 585
R121 B.n787 B.n42 585
R122 B.n551 B.n41 585
R123 B.n788 B.n41 585
R124 B.n550 B.n549 585
R125 B.n549 B.n37 585
R126 B.n548 B.n36 585
R127 B.n794 B.n36 585
R128 B.n547 B.n35 585
R129 B.n795 B.n35 585
R130 B.n546 B.n34 585
R131 B.n796 B.n34 585
R132 B.n545 B.n544 585
R133 B.n544 B.n30 585
R134 B.n543 B.n29 585
R135 B.n802 B.n29 585
R136 B.n542 B.n28 585
R137 B.n803 B.n28 585
R138 B.n541 B.n27 585
R139 B.n804 B.n27 585
R140 B.n540 B.n539 585
R141 B.n539 B.n23 585
R142 B.n538 B.n22 585
R143 B.n810 B.n22 585
R144 B.n537 B.n21 585
R145 B.n811 B.n21 585
R146 B.n536 B.n20 585
R147 B.n812 B.n20 585
R148 B.n535 B.n534 585
R149 B.n534 B.n19 585
R150 B.n533 B.n15 585
R151 B.n818 B.n15 585
R152 B.n532 B.n14 585
R153 B.n819 B.n14 585
R154 B.n531 B.n13 585
R155 B.n820 B.n13 585
R156 B.n530 B.n529 585
R157 B.n529 B.n12 585
R158 B.n528 B.n527 585
R159 B.n528 B.n8 585
R160 B.n526 B.n7 585
R161 B.n827 B.n7 585
R162 B.n525 B.n6 585
R163 B.n828 B.n6 585
R164 B.n524 B.n5 585
R165 B.n829 B.n5 585
R166 B.n523 B.n522 585
R167 B.n522 B.n4 585
R168 B.n521 B.n116 585
R169 B.n521 B.n520 585
R170 B.n511 B.n117 585
R171 B.n118 B.n117 585
R172 B.n513 B.n512 585
R173 B.n514 B.n513 585
R174 B.n510 B.n123 585
R175 B.n123 B.n122 585
R176 B.n509 B.n508 585
R177 B.n508 B.n507 585
R178 B.n125 B.n124 585
R179 B.n500 B.n125 585
R180 B.n499 B.n498 585
R181 B.n501 B.n499 585
R182 B.n497 B.n130 585
R183 B.n130 B.n129 585
R184 B.n496 B.n495 585
R185 B.n495 B.n494 585
R186 B.n132 B.n131 585
R187 B.n133 B.n132 585
R188 B.n487 B.n486 585
R189 B.n488 B.n487 585
R190 B.n485 B.n138 585
R191 B.n138 B.n137 585
R192 B.n484 B.n483 585
R193 B.n483 B.n482 585
R194 B.n140 B.n139 585
R195 B.n141 B.n140 585
R196 B.n475 B.n474 585
R197 B.n476 B.n475 585
R198 B.n473 B.n146 585
R199 B.n146 B.n145 585
R200 B.n472 B.n471 585
R201 B.n471 B.n470 585
R202 B.n148 B.n147 585
R203 B.n149 B.n148 585
R204 B.n463 B.n462 585
R205 B.n464 B.n463 585
R206 B.n461 B.n154 585
R207 B.n154 B.n153 585
R208 B.n460 B.n459 585
R209 B.n459 B.n458 585
R210 B.n156 B.n155 585
R211 B.n157 B.n156 585
R212 B.n451 B.n450 585
R213 B.n452 B.n451 585
R214 B.n449 B.n162 585
R215 B.n162 B.n161 585
R216 B.n448 B.n447 585
R217 B.n447 B.n446 585
R218 B.n164 B.n163 585
R219 B.n165 B.n164 585
R220 B.n439 B.n438 585
R221 B.n440 B.n439 585
R222 B.n437 B.n170 585
R223 B.n170 B.n169 585
R224 B.n436 B.n435 585
R225 B.n435 B.n434 585
R226 B.n431 B.n174 585
R227 B.n430 B.n429 585
R228 B.n427 B.n175 585
R229 B.n427 B.n173 585
R230 B.n426 B.n425 585
R231 B.n424 B.n423 585
R232 B.n422 B.n177 585
R233 B.n420 B.n419 585
R234 B.n418 B.n178 585
R235 B.n417 B.n416 585
R236 B.n414 B.n179 585
R237 B.n412 B.n411 585
R238 B.n410 B.n180 585
R239 B.n409 B.n408 585
R240 B.n406 B.n181 585
R241 B.n404 B.n403 585
R242 B.n402 B.n182 585
R243 B.n401 B.n400 585
R244 B.n398 B.n183 585
R245 B.n396 B.n395 585
R246 B.n394 B.n184 585
R247 B.n393 B.n392 585
R248 B.n390 B.n185 585
R249 B.n388 B.n387 585
R250 B.n386 B.n186 585
R251 B.n385 B.n384 585
R252 B.n382 B.n187 585
R253 B.n380 B.n379 585
R254 B.n378 B.n188 585
R255 B.n377 B.n376 585
R256 B.n374 B.n189 585
R257 B.n372 B.n371 585
R258 B.n370 B.n190 585
R259 B.n369 B.n368 585
R260 B.n366 B.n191 585
R261 B.n364 B.n363 585
R262 B.n362 B.n192 585
R263 B.n361 B.n360 585
R264 B.n358 B.n193 585
R265 B.n356 B.n355 585
R266 B.n354 B.n194 585
R267 B.n353 B.n352 585
R268 B.n350 B.n195 585
R269 B.n348 B.n347 585
R270 B.n346 B.n196 585
R271 B.n345 B.n344 585
R272 B.n342 B.n197 585
R273 B.n340 B.n339 585
R274 B.n338 B.n198 585
R275 B.n337 B.n336 585
R276 B.n334 B.n202 585
R277 B.n332 B.n331 585
R278 B.n330 B.n203 585
R279 B.n329 B.n328 585
R280 B.n326 B.n204 585
R281 B.n324 B.n323 585
R282 B.n322 B.n205 585
R283 B.n320 B.n319 585
R284 B.n317 B.n208 585
R285 B.n315 B.n314 585
R286 B.n313 B.n209 585
R287 B.n312 B.n311 585
R288 B.n309 B.n210 585
R289 B.n307 B.n306 585
R290 B.n305 B.n211 585
R291 B.n304 B.n303 585
R292 B.n301 B.n212 585
R293 B.n299 B.n298 585
R294 B.n297 B.n213 585
R295 B.n296 B.n295 585
R296 B.n293 B.n214 585
R297 B.n291 B.n290 585
R298 B.n289 B.n215 585
R299 B.n288 B.n287 585
R300 B.n285 B.n216 585
R301 B.n283 B.n282 585
R302 B.n281 B.n217 585
R303 B.n280 B.n279 585
R304 B.n277 B.n218 585
R305 B.n275 B.n274 585
R306 B.n273 B.n219 585
R307 B.n272 B.n271 585
R308 B.n269 B.n220 585
R309 B.n267 B.n266 585
R310 B.n265 B.n221 585
R311 B.n264 B.n263 585
R312 B.n261 B.n222 585
R313 B.n259 B.n258 585
R314 B.n257 B.n223 585
R315 B.n256 B.n255 585
R316 B.n253 B.n224 585
R317 B.n251 B.n250 585
R318 B.n249 B.n225 585
R319 B.n248 B.n247 585
R320 B.n245 B.n226 585
R321 B.n243 B.n242 585
R322 B.n241 B.n227 585
R323 B.n240 B.n239 585
R324 B.n237 B.n228 585
R325 B.n235 B.n234 585
R326 B.n233 B.n229 585
R327 B.n232 B.n231 585
R328 B.n172 B.n171 585
R329 B.n173 B.n172 585
R330 B.n433 B.n432 585
R331 B.n434 B.n433 585
R332 B.n168 B.n167 585
R333 B.n169 B.n168 585
R334 B.n442 B.n441 585
R335 B.n441 B.n440 585
R336 B.n443 B.n166 585
R337 B.n166 B.n165 585
R338 B.n445 B.n444 585
R339 B.n446 B.n445 585
R340 B.n160 B.n159 585
R341 B.n161 B.n160 585
R342 B.n454 B.n453 585
R343 B.n453 B.n452 585
R344 B.n455 B.n158 585
R345 B.n158 B.n157 585
R346 B.n457 B.n456 585
R347 B.n458 B.n457 585
R348 B.n152 B.n151 585
R349 B.n153 B.n152 585
R350 B.n466 B.n465 585
R351 B.n465 B.n464 585
R352 B.n467 B.n150 585
R353 B.n150 B.n149 585
R354 B.n469 B.n468 585
R355 B.n470 B.n469 585
R356 B.n144 B.n143 585
R357 B.n145 B.n144 585
R358 B.n478 B.n477 585
R359 B.n477 B.n476 585
R360 B.n479 B.n142 585
R361 B.n142 B.n141 585
R362 B.n481 B.n480 585
R363 B.n482 B.n481 585
R364 B.n136 B.n135 585
R365 B.n137 B.n136 585
R366 B.n490 B.n489 585
R367 B.n489 B.n488 585
R368 B.n491 B.n134 585
R369 B.n134 B.n133 585
R370 B.n493 B.n492 585
R371 B.n494 B.n493 585
R372 B.n128 B.n127 585
R373 B.n129 B.n128 585
R374 B.n503 B.n502 585
R375 B.n502 B.n501 585
R376 B.n504 B.n126 585
R377 B.n500 B.n126 585
R378 B.n506 B.n505 585
R379 B.n507 B.n506 585
R380 B.n121 B.n120 585
R381 B.n122 B.n121 585
R382 B.n516 B.n515 585
R383 B.n515 B.n514 585
R384 B.n517 B.n119 585
R385 B.n119 B.n118 585
R386 B.n519 B.n518 585
R387 B.n520 B.n519 585
R388 B.n3 B.n0 585
R389 B.n4 B.n3 585
R390 B.n826 B.n1 585
R391 B.n827 B.n826 585
R392 B.n825 B.n824 585
R393 B.n825 B.n8 585
R394 B.n823 B.n9 585
R395 B.n12 B.n9 585
R396 B.n822 B.n821 585
R397 B.n821 B.n820 585
R398 B.n11 B.n10 585
R399 B.n819 B.n11 585
R400 B.n817 B.n816 585
R401 B.n818 B.n817 585
R402 B.n815 B.n16 585
R403 B.n19 B.n16 585
R404 B.n814 B.n813 585
R405 B.n813 B.n812 585
R406 B.n18 B.n17 585
R407 B.n811 B.n18 585
R408 B.n809 B.n808 585
R409 B.n810 B.n809 585
R410 B.n807 B.n24 585
R411 B.n24 B.n23 585
R412 B.n806 B.n805 585
R413 B.n805 B.n804 585
R414 B.n26 B.n25 585
R415 B.n803 B.n26 585
R416 B.n801 B.n800 585
R417 B.n802 B.n801 585
R418 B.n799 B.n31 585
R419 B.n31 B.n30 585
R420 B.n798 B.n797 585
R421 B.n797 B.n796 585
R422 B.n33 B.n32 585
R423 B.n795 B.n33 585
R424 B.n793 B.n792 585
R425 B.n794 B.n793 585
R426 B.n791 B.n38 585
R427 B.n38 B.n37 585
R428 B.n790 B.n789 585
R429 B.n789 B.n788 585
R430 B.n40 B.n39 585
R431 B.n787 B.n40 585
R432 B.n785 B.n784 585
R433 B.n786 B.n785 585
R434 B.n783 B.n45 585
R435 B.n45 B.n44 585
R436 B.n782 B.n781 585
R437 B.n781 B.n780 585
R438 B.n47 B.n46 585
R439 B.n779 B.n47 585
R440 B.n777 B.n776 585
R441 B.n778 B.n777 585
R442 B.n775 B.n52 585
R443 B.n52 B.n51 585
R444 B.n774 B.n773 585
R445 B.n773 B.n772 585
R446 B.n54 B.n53 585
R447 B.n771 B.n54 585
R448 B.n769 B.n768 585
R449 B.n770 B.n769 585
R450 B.n830 B.n829 585
R451 B.n828 B.n2 585
R452 B.n769 B.n59 545.355
R453 B.n565 B.n57 545.355
R454 B.n435 B.n172 545.355
R455 B.n433 B.n174 545.355
R456 B.n82 B.t12 303.606
R457 B.n90 B.t1 303.606
R458 B.n206 B.t9 303.606
R459 B.n199 B.t5 303.606
R460 B.n564 B.n58 256.663
R461 B.n570 B.n58 256.663
R462 B.n572 B.n58 256.663
R463 B.n578 B.n58 256.663
R464 B.n580 B.n58 256.663
R465 B.n586 B.n58 256.663
R466 B.n588 B.n58 256.663
R467 B.n594 B.n58 256.663
R468 B.n596 B.n58 256.663
R469 B.n602 B.n58 256.663
R470 B.n604 B.n58 256.663
R471 B.n610 B.n58 256.663
R472 B.n612 B.n58 256.663
R473 B.n618 B.n58 256.663
R474 B.n620 B.n58 256.663
R475 B.n626 B.n58 256.663
R476 B.n628 B.n58 256.663
R477 B.n634 B.n58 256.663
R478 B.n636 B.n58 256.663
R479 B.n642 B.n58 256.663
R480 B.n644 B.n58 256.663
R481 B.n650 B.n58 256.663
R482 B.n93 B.n58 256.663
R483 B.n656 B.n58 256.663
R484 B.n662 B.n58 256.663
R485 B.n664 B.n58 256.663
R486 B.n670 B.n58 256.663
R487 B.n85 B.n58 256.663
R488 B.n676 B.n58 256.663
R489 B.n682 B.n58 256.663
R490 B.n684 B.n58 256.663
R491 B.n690 B.n58 256.663
R492 B.n692 B.n58 256.663
R493 B.n698 B.n58 256.663
R494 B.n700 B.n58 256.663
R495 B.n706 B.n58 256.663
R496 B.n708 B.n58 256.663
R497 B.n714 B.n58 256.663
R498 B.n716 B.n58 256.663
R499 B.n722 B.n58 256.663
R500 B.n724 B.n58 256.663
R501 B.n730 B.n58 256.663
R502 B.n732 B.n58 256.663
R503 B.n738 B.n58 256.663
R504 B.n740 B.n58 256.663
R505 B.n746 B.n58 256.663
R506 B.n748 B.n58 256.663
R507 B.n754 B.n58 256.663
R508 B.n756 B.n58 256.663
R509 B.n762 B.n58 256.663
R510 B.n764 B.n58 256.663
R511 B.n428 B.n173 256.663
R512 B.n176 B.n173 256.663
R513 B.n421 B.n173 256.663
R514 B.n415 B.n173 256.663
R515 B.n413 B.n173 256.663
R516 B.n407 B.n173 256.663
R517 B.n405 B.n173 256.663
R518 B.n399 B.n173 256.663
R519 B.n397 B.n173 256.663
R520 B.n391 B.n173 256.663
R521 B.n389 B.n173 256.663
R522 B.n383 B.n173 256.663
R523 B.n381 B.n173 256.663
R524 B.n375 B.n173 256.663
R525 B.n373 B.n173 256.663
R526 B.n367 B.n173 256.663
R527 B.n365 B.n173 256.663
R528 B.n359 B.n173 256.663
R529 B.n357 B.n173 256.663
R530 B.n351 B.n173 256.663
R531 B.n349 B.n173 256.663
R532 B.n343 B.n173 256.663
R533 B.n341 B.n173 256.663
R534 B.n335 B.n173 256.663
R535 B.n333 B.n173 256.663
R536 B.n327 B.n173 256.663
R537 B.n325 B.n173 256.663
R538 B.n318 B.n173 256.663
R539 B.n316 B.n173 256.663
R540 B.n310 B.n173 256.663
R541 B.n308 B.n173 256.663
R542 B.n302 B.n173 256.663
R543 B.n300 B.n173 256.663
R544 B.n294 B.n173 256.663
R545 B.n292 B.n173 256.663
R546 B.n286 B.n173 256.663
R547 B.n284 B.n173 256.663
R548 B.n278 B.n173 256.663
R549 B.n276 B.n173 256.663
R550 B.n270 B.n173 256.663
R551 B.n268 B.n173 256.663
R552 B.n262 B.n173 256.663
R553 B.n260 B.n173 256.663
R554 B.n254 B.n173 256.663
R555 B.n252 B.n173 256.663
R556 B.n246 B.n173 256.663
R557 B.n244 B.n173 256.663
R558 B.n238 B.n173 256.663
R559 B.n236 B.n173 256.663
R560 B.n230 B.n173 256.663
R561 B.n832 B.n831 256.663
R562 B.n765 B.n763 163.367
R563 B.n761 B.n61 163.367
R564 B.n757 B.n755 163.367
R565 B.n753 B.n63 163.367
R566 B.n749 B.n747 163.367
R567 B.n745 B.n65 163.367
R568 B.n741 B.n739 163.367
R569 B.n737 B.n67 163.367
R570 B.n733 B.n731 163.367
R571 B.n729 B.n69 163.367
R572 B.n725 B.n723 163.367
R573 B.n721 B.n71 163.367
R574 B.n717 B.n715 163.367
R575 B.n713 B.n73 163.367
R576 B.n709 B.n707 163.367
R577 B.n705 B.n75 163.367
R578 B.n701 B.n699 163.367
R579 B.n697 B.n77 163.367
R580 B.n693 B.n691 163.367
R581 B.n689 B.n79 163.367
R582 B.n685 B.n683 163.367
R583 B.n681 B.n81 163.367
R584 B.n677 B.n675 163.367
R585 B.n672 B.n671 163.367
R586 B.n669 B.n87 163.367
R587 B.n665 B.n663 163.367
R588 B.n661 B.n89 163.367
R589 B.n657 B.n655 163.367
R590 B.n652 B.n651 163.367
R591 B.n649 B.n95 163.367
R592 B.n645 B.n643 163.367
R593 B.n641 B.n97 163.367
R594 B.n637 B.n635 163.367
R595 B.n633 B.n99 163.367
R596 B.n629 B.n627 163.367
R597 B.n625 B.n101 163.367
R598 B.n621 B.n619 163.367
R599 B.n617 B.n103 163.367
R600 B.n613 B.n611 163.367
R601 B.n609 B.n105 163.367
R602 B.n605 B.n603 163.367
R603 B.n601 B.n107 163.367
R604 B.n597 B.n595 163.367
R605 B.n593 B.n109 163.367
R606 B.n589 B.n587 163.367
R607 B.n585 B.n111 163.367
R608 B.n581 B.n579 163.367
R609 B.n577 B.n113 163.367
R610 B.n573 B.n571 163.367
R611 B.n569 B.n115 163.367
R612 B.n435 B.n170 163.367
R613 B.n439 B.n170 163.367
R614 B.n439 B.n164 163.367
R615 B.n447 B.n164 163.367
R616 B.n447 B.n162 163.367
R617 B.n451 B.n162 163.367
R618 B.n451 B.n156 163.367
R619 B.n459 B.n156 163.367
R620 B.n459 B.n154 163.367
R621 B.n463 B.n154 163.367
R622 B.n463 B.n148 163.367
R623 B.n471 B.n148 163.367
R624 B.n471 B.n146 163.367
R625 B.n475 B.n146 163.367
R626 B.n475 B.n140 163.367
R627 B.n483 B.n140 163.367
R628 B.n483 B.n138 163.367
R629 B.n487 B.n138 163.367
R630 B.n487 B.n132 163.367
R631 B.n495 B.n132 163.367
R632 B.n495 B.n130 163.367
R633 B.n499 B.n130 163.367
R634 B.n499 B.n125 163.367
R635 B.n508 B.n125 163.367
R636 B.n508 B.n123 163.367
R637 B.n513 B.n123 163.367
R638 B.n513 B.n117 163.367
R639 B.n521 B.n117 163.367
R640 B.n522 B.n521 163.367
R641 B.n522 B.n5 163.367
R642 B.n6 B.n5 163.367
R643 B.n7 B.n6 163.367
R644 B.n528 B.n7 163.367
R645 B.n529 B.n528 163.367
R646 B.n529 B.n13 163.367
R647 B.n14 B.n13 163.367
R648 B.n15 B.n14 163.367
R649 B.n534 B.n15 163.367
R650 B.n534 B.n20 163.367
R651 B.n21 B.n20 163.367
R652 B.n22 B.n21 163.367
R653 B.n539 B.n22 163.367
R654 B.n539 B.n27 163.367
R655 B.n28 B.n27 163.367
R656 B.n29 B.n28 163.367
R657 B.n544 B.n29 163.367
R658 B.n544 B.n34 163.367
R659 B.n35 B.n34 163.367
R660 B.n36 B.n35 163.367
R661 B.n549 B.n36 163.367
R662 B.n549 B.n41 163.367
R663 B.n42 B.n41 163.367
R664 B.n43 B.n42 163.367
R665 B.n554 B.n43 163.367
R666 B.n554 B.n48 163.367
R667 B.n49 B.n48 163.367
R668 B.n50 B.n49 163.367
R669 B.n559 B.n50 163.367
R670 B.n559 B.n55 163.367
R671 B.n56 B.n55 163.367
R672 B.n57 B.n56 163.367
R673 B.n429 B.n427 163.367
R674 B.n427 B.n426 163.367
R675 B.n423 B.n422 163.367
R676 B.n420 B.n178 163.367
R677 B.n416 B.n414 163.367
R678 B.n412 B.n180 163.367
R679 B.n408 B.n406 163.367
R680 B.n404 B.n182 163.367
R681 B.n400 B.n398 163.367
R682 B.n396 B.n184 163.367
R683 B.n392 B.n390 163.367
R684 B.n388 B.n186 163.367
R685 B.n384 B.n382 163.367
R686 B.n380 B.n188 163.367
R687 B.n376 B.n374 163.367
R688 B.n372 B.n190 163.367
R689 B.n368 B.n366 163.367
R690 B.n364 B.n192 163.367
R691 B.n360 B.n358 163.367
R692 B.n356 B.n194 163.367
R693 B.n352 B.n350 163.367
R694 B.n348 B.n196 163.367
R695 B.n344 B.n342 163.367
R696 B.n340 B.n198 163.367
R697 B.n336 B.n334 163.367
R698 B.n332 B.n203 163.367
R699 B.n328 B.n326 163.367
R700 B.n324 B.n205 163.367
R701 B.n319 B.n317 163.367
R702 B.n315 B.n209 163.367
R703 B.n311 B.n309 163.367
R704 B.n307 B.n211 163.367
R705 B.n303 B.n301 163.367
R706 B.n299 B.n213 163.367
R707 B.n295 B.n293 163.367
R708 B.n291 B.n215 163.367
R709 B.n287 B.n285 163.367
R710 B.n283 B.n217 163.367
R711 B.n279 B.n277 163.367
R712 B.n275 B.n219 163.367
R713 B.n271 B.n269 163.367
R714 B.n267 B.n221 163.367
R715 B.n263 B.n261 163.367
R716 B.n259 B.n223 163.367
R717 B.n255 B.n253 163.367
R718 B.n251 B.n225 163.367
R719 B.n247 B.n245 163.367
R720 B.n243 B.n227 163.367
R721 B.n239 B.n237 163.367
R722 B.n235 B.n229 163.367
R723 B.n231 B.n172 163.367
R724 B.n433 B.n168 163.367
R725 B.n441 B.n168 163.367
R726 B.n441 B.n166 163.367
R727 B.n445 B.n166 163.367
R728 B.n445 B.n160 163.367
R729 B.n453 B.n160 163.367
R730 B.n453 B.n158 163.367
R731 B.n457 B.n158 163.367
R732 B.n457 B.n152 163.367
R733 B.n465 B.n152 163.367
R734 B.n465 B.n150 163.367
R735 B.n469 B.n150 163.367
R736 B.n469 B.n144 163.367
R737 B.n477 B.n144 163.367
R738 B.n477 B.n142 163.367
R739 B.n481 B.n142 163.367
R740 B.n481 B.n136 163.367
R741 B.n489 B.n136 163.367
R742 B.n489 B.n134 163.367
R743 B.n493 B.n134 163.367
R744 B.n493 B.n128 163.367
R745 B.n502 B.n128 163.367
R746 B.n502 B.n126 163.367
R747 B.n506 B.n126 163.367
R748 B.n506 B.n121 163.367
R749 B.n515 B.n121 163.367
R750 B.n515 B.n119 163.367
R751 B.n519 B.n119 163.367
R752 B.n519 B.n3 163.367
R753 B.n830 B.n3 163.367
R754 B.n826 B.n2 163.367
R755 B.n826 B.n825 163.367
R756 B.n825 B.n9 163.367
R757 B.n821 B.n9 163.367
R758 B.n821 B.n11 163.367
R759 B.n817 B.n11 163.367
R760 B.n817 B.n16 163.367
R761 B.n813 B.n16 163.367
R762 B.n813 B.n18 163.367
R763 B.n809 B.n18 163.367
R764 B.n809 B.n24 163.367
R765 B.n805 B.n24 163.367
R766 B.n805 B.n26 163.367
R767 B.n801 B.n26 163.367
R768 B.n801 B.n31 163.367
R769 B.n797 B.n31 163.367
R770 B.n797 B.n33 163.367
R771 B.n793 B.n33 163.367
R772 B.n793 B.n38 163.367
R773 B.n789 B.n38 163.367
R774 B.n789 B.n40 163.367
R775 B.n785 B.n40 163.367
R776 B.n785 B.n45 163.367
R777 B.n781 B.n45 163.367
R778 B.n781 B.n47 163.367
R779 B.n777 B.n47 163.367
R780 B.n777 B.n52 163.367
R781 B.n773 B.n52 163.367
R782 B.n773 B.n54 163.367
R783 B.n769 B.n54 163.367
R784 B.n90 B.t3 142.453
R785 B.n206 B.t11 142.453
R786 B.n82 B.t13 142.435
R787 B.n199 B.t8 142.435
R788 B.n83 B.n82 73.8914
R789 B.n91 B.n90 73.8914
R790 B.n207 B.n206 73.8914
R791 B.n200 B.n199 73.8914
R792 B.n434 B.n173 72.6557
R793 B.n770 B.n58 72.6557
R794 B.n764 B.n59 71.676
R795 B.n763 B.n762 71.676
R796 B.n756 B.n61 71.676
R797 B.n755 B.n754 71.676
R798 B.n748 B.n63 71.676
R799 B.n747 B.n746 71.676
R800 B.n740 B.n65 71.676
R801 B.n739 B.n738 71.676
R802 B.n732 B.n67 71.676
R803 B.n731 B.n730 71.676
R804 B.n724 B.n69 71.676
R805 B.n723 B.n722 71.676
R806 B.n716 B.n71 71.676
R807 B.n715 B.n714 71.676
R808 B.n708 B.n73 71.676
R809 B.n707 B.n706 71.676
R810 B.n700 B.n75 71.676
R811 B.n699 B.n698 71.676
R812 B.n692 B.n77 71.676
R813 B.n691 B.n690 71.676
R814 B.n684 B.n79 71.676
R815 B.n683 B.n682 71.676
R816 B.n676 B.n81 71.676
R817 B.n675 B.n85 71.676
R818 B.n671 B.n670 71.676
R819 B.n664 B.n87 71.676
R820 B.n663 B.n662 71.676
R821 B.n656 B.n89 71.676
R822 B.n655 B.n93 71.676
R823 B.n651 B.n650 71.676
R824 B.n644 B.n95 71.676
R825 B.n643 B.n642 71.676
R826 B.n636 B.n97 71.676
R827 B.n635 B.n634 71.676
R828 B.n628 B.n99 71.676
R829 B.n627 B.n626 71.676
R830 B.n620 B.n101 71.676
R831 B.n619 B.n618 71.676
R832 B.n612 B.n103 71.676
R833 B.n611 B.n610 71.676
R834 B.n604 B.n105 71.676
R835 B.n603 B.n602 71.676
R836 B.n596 B.n107 71.676
R837 B.n595 B.n594 71.676
R838 B.n588 B.n109 71.676
R839 B.n587 B.n586 71.676
R840 B.n580 B.n111 71.676
R841 B.n579 B.n578 71.676
R842 B.n572 B.n113 71.676
R843 B.n571 B.n570 71.676
R844 B.n564 B.n115 71.676
R845 B.n565 B.n564 71.676
R846 B.n570 B.n569 71.676
R847 B.n573 B.n572 71.676
R848 B.n578 B.n577 71.676
R849 B.n581 B.n580 71.676
R850 B.n586 B.n585 71.676
R851 B.n589 B.n588 71.676
R852 B.n594 B.n593 71.676
R853 B.n597 B.n596 71.676
R854 B.n602 B.n601 71.676
R855 B.n605 B.n604 71.676
R856 B.n610 B.n609 71.676
R857 B.n613 B.n612 71.676
R858 B.n618 B.n617 71.676
R859 B.n621 B.n620 71.676
R860 B.n626 B.n625 71.676
R861 B.n629 B.n628 71.676
R862 B.n634 B.n633 71.676
R863 B.n637 B.n636 71.676
R864 B.n642 B.n641 71.676
R865 B.n645 B.n644 71.676
R866 B.n650 B.n649 71.676
R867 B.n652 B.n93 71.676
R868 B.n657 B.n656 71.676
R869 B.n662 B.n661 71.676
R870 B.n665 B.n664 71.676
R871 B.n670 B.n669 71.676
R872 B.n672 B.n85 71.676
R873 B.n677 B.n676 71.676
R874 B.n682 B.n681 71.676
R875 B.n685 B.n684 71.676
R876 B.n690 B.n689 71.676
R877 B.n693 B.n692 71.676
R878 B.n698 B.n697 71.676
R879 B.n701 B.n700 71.676
R880 B.n706 B.n705 71.676
R881 B.n709 B.n708 71.676
R882 B.n714 B.n713 71.676
R883 B.n717 B.n716 71.676
R884 B.n722 B.n721 71.676
R885 B.n725 B.n724 71.676
R886 B.n730 B.n729 71.676
R887 B.n733 B.n732 71.676
R888 B.n738 B.n737 71.676
R889 B.n741 B.n740 71.676
R890 B.n746 B.n745 71.676
R891 B.n749 B.n748 71.676
R892 B.n754 B.n753 71.676
R893 B.n757 B.n756 71.676
R894 B.n762 B.n761 71.676
R895 B.n765 B.n764 71.676
R896 B.n428 B.n174 71.676
R897 B.n426 B.n176 71.676
R898 B.n422 B.n421 71.676
R899 B.n415 B.n178 71.676
R900 B.n414 B.n413 71.676
R901 B.n407 B.n180 71.676
R902 B.n406 B.n405 71.676
R903 B.n399 B.n182 71.676
R904 B.n398 B.n397 71.676
R905 B.n391 B.n184 71.676
R906 B.n390 B.n389 71.676
R907 B.n383 B.n186 71.676
R908 B.n382 B.n381 71.676
R909 B.n375 B.n188 71.676
R910 B.n374 B.n373 71.676
R911 B.n367 B.n190 71.676
R912 B.n366 B.n365 71.676
R913 B.n359 B.n192 71.676
R914 B.n358 B.n357 71.676
R915 B.n351 B.n194 71.676
R916 B.n350 B.n349 71.676
R917 B.n343 B.n196 71.676
R918 B.n342 B.n341 71.676
R919 B.n335 B.n198 71.676
R920 B.n334 B.n333 71.676
R921 B.n327 B.n203 71.676
R922 B.n326 B.n325 71.676
R923 B.n318 B.n205 71.676
R924 B.n317 B.n316 71.676
R925 B.n310 B.n209 71.676
R926 B.n309 B.n308 71.676
R927 B.n302 B.n211 71.676
R928 B.n301 B.n300 71.676
R929 B.n294 B.n213 71.676
R930 B.n293 B.n292 71.676
R931 B.n286 B.n215 71.676
R932 B.n285 B.n284 71.676
R933 B.n278 B.n217 71.676
R934 B.n277 B.n276 71.676
R935 B.n270 B.n219 71.676
R936 B.n269 B.n268 71.676
R937 B.n262 B.n221 71.676
R938 B.n261 B.n260 71.676
R939 B.n254 B.n223 71.676
R940 B.n253 B.n252 71.676
R941 B.n246 B.n225 71.676
R942 B.n245 B.n244 71.676
R943 B.n238 B.n227 71.676
R944 B.n237 B.n236 71.676
R945 B.n230 B.n229 71.676
R946 B.n429 B.n428 71.676
R947 B.n423 B.n176 71.676
R948 B.n421 B.n420 71.676
R949 B.n416 B.n415 71.676
R950 B.n413 B.n412 71.676
R951 B.n408 B.n407 71.676
R952 B.n405 B.n404 71.676
R953 B.n400 B.n399 71.676
R954 B.n397 B.n396 71.676
R955 B.n392 B.n391 71.676
R956 B.n389 B.n388 71.676
R957 B.n384 B.n383 71.676
R958 B.n381 B.n380 71.676
R959 B.n376 B.n375 71.676
R960 B.n373 B.n372 71.676
R961 B.n368 B.n367 71.676
R962 B.n365 B.n364 71.676
R963 B.n360 B.n359 71.676
R964 B.n357 B.n356 71.676
R965 B.n352 B.n351 71.676
R966 B.n349 B.n348 71.676
R967 B.n344 B.n343 71.676
R968 B.n341 B.n340 71.676
R969 B.n336 B.n335 71.676
R970 B.n333 B.n332 71.676
R971 B.n328 B.n327 71.676
R972 B.n325 B.n324 71.676
R973 B.n319 B.n318 71.676
R974 B.n316 B.n315 71.676
R975 B.n311 B.n310 71.676
R976 B.n308 B.n307 71.676
R977 B.n303 B.n302 71.676
R978 B.n300 B.n299 71.676
R979 B.n295 B.n294 71.676
R980 B.n292 B.n291 71.676
R981 B.n287 B.n286 71.676
R982 B.n284 B.n283 71.676
R983 B.n279 B.n278 71.676
R984 B.n276 B.n275 71.676
R985 B.n271 B.n270 71.676
R986 B.n268 B.n267 71.676
R987 B.n263 B.n262 71.676
R988 B.n260 B.n259 71.676
R989 B.n255 B.n254 71.676
R990 B.n252 B.n251 71.676
R991 B.n247 B.n246 71.676
R992 B.n244 B.n243 71.676
R993 B.n239 B.n238 71.676
R994 B.n236 B.n235 71.676
R995 B.n231 B.n230 71.676
R996 B.n831 B.n830 71.676
R997 B.n831 B.n2 71.676
R998 B.n91 B.t4 68.5626
R999 B.n207 B.t10 68.5626
R1000 B.n83 B.t14 68.5449
R1001 B.n200 B.t7 68.5449
R1002 B.n84 B.n83 59.5399
R1003 B.n92 B.n91 59.5399
R1004 B.n321 B.n207 59.5399
R1005 B.n201 B.n200 59.5399
R1006 B.n434 B.n169 39.5249
R1007 B.n440 B.n169 39.5249
R1008 B.n440 B.n165 39.5249
R1009 B.n446 B.n165 39.5249
R1010 B.n446 B.n161 39.5249
R1011 B.n452 B.n161 39.5249
R1012 B.n452 B.n157 39.5249
R1013 B.n458 B.n157 39.5249
R1014 B.n464 B.n153 39.5249
R1015 B.n464 B.n149 39.5249
R1016 B.n470 B.n149 39.5249
R1017 B.n470 B.n145 39.5249
R1018 B.n476 B.n145 39.5249
R1019 B.n476 B.n141 39.5249
R1020 B.n482 B.n141 39.5249
R1021 B.n482 B.n137 39.5249
R1022 B.n488 B.n137 39.5249
R1023 B.n488 B.n133 39.5249
R1024 B.n494 B.n133 39.5249
R1025 B.n494 B.n129 39.5249
R1026 B.n501 B.n129 39.5249
R1027 B.n501 B.n500 39.5249
R1028 B.n507 B.n122 39.5249
R1029 B.n514 B.n122 39.5249
R1030 B.n514 B.n118 39.5249
R1031 B.n520 B.n118 39.5249
R1032 B.n520 B.n4 39.5249
R1033 B.n829 B.n4 39.5249
R1034 B.n829 B.n828 39.5249
R1035 B.n828 B.n827 39.5249
R1036 B.n827 B.n8 39.5249
R1037 B.n12 B.n8 39.5249
R1038 B.n820 B.n12 39.5249
R1039 B.n820 B.n819 39.5249
R1040 B.n819 B.n818 39.5249
R1041 B.n812 B.n19 39.5249
R1042 B.n812 B.n811 39.5249
R1043 B.n811 B.n810 39.5249
R1044 B.n810 B.n23 39.5249
R1045 B.n804 B.n23 39.5249
R1046 B.n804 B.n803 39.5249
R1047 B.n803 B.n802 39.5249
R1048 B.n802 B.n30 39.5249
R1049 B.n796 B.n30 39.5249
R1050 B.n796 B.n795 39.5249
R1051 B.n795 B.n794 39.5249
R1052 B.n794 B.n37 39.5249
R1053 B.n788 B.n37 39.5249
R1054 B.n788 B.n787 39.5249
R1055 B.n786 B.n44 39.5249
R1056 B.n780 B.n44 39.5249
R1057 B.n780 B.n779 39.5249
R1058 B.n779 B.n778 39.5249
R1059 B.n778 B.n51 39.5249
R1060 B.n772 B.n51 39.5249
R1061 B.n772 B.n771 39.5249
R1062 B.n771 B.n770 39.5249
R1063 B.n432 B.n431 35.4346
R1064 B.n436 B.n171 35.4346
R1065 B.n566 B.n563 35.4346
R1066 B.n768 B.n767 35.4346
R1067 B.n458 B.t6 34.875
R1068 B.t2 B.n786 34.875
R1069 B.n507 B.t0 27.9001
R1070 B.n818 B.t15 27.9001
R1071 B B.n832 18.0485
R1072 B.n500 B.t0 11.6253
R1073 B.n19 B.t15 11.6253
R1074 B.n432 B.n167 10.6151
R1075 B.n442 B.n167 10.6151
R1076 B.n443 B.n442 10.6151
R1077 B.n444 B.n443 10.6151
R1078 B.n444 B.n159 10.6151
R1079 B.n454 B.n159 10.6151
R1080 B.n455 B.n454 10.6151
R1081 B.n456 B.n455 10.6151
R1082 B.n456 B.n151 10.6151
R1083 B.n466 B.n151 10.6151
R1084 B.n467 B.n466 10.6151
R1085 B.n468 B.n467 10.6151
R1086 B.n468 B.n143 10.6151
R1087 B.n478 B.n143 10.6151
R1088 B.n479 B.n478 10.6151
R1089 B.n480 B.n479 10.6151
R1090 B.n480 B.n135 10.6151
R1091 B.n490 B.n135 10.6151
R1092 B.n491 B.n490 10.6151
R1093 B.n492 B.n491 10.6151
R1094 B.n492 B.n127 10.6151
R1095 B.n503 B.n127 10.6151
R1096 B.n504 B.n503 10.6151
R1097 B.n505 B.n504 10.6151
R1098 B.n505 B.n120 10.6151
R1099 B.n516 B.n120 10.6151
R1100 B.n517 B.n516 10.6151
R1101 B.n518 B.n517 10.6151
R1102 B.n518 B.n0 10.6151
R1103 B.n431 B.n430 10.6151
R1104 B.n430 B.n175 10.6151
R1105 B.n425 B.n175 10.6151
R1106 B.n425 B.n424 10.6151
R1107 B.n424 B.n177 10.6151
R1108 B.n419 B.n177 10.6151
R1109 B.n419 B.n418 10.6151
R1110 B.n418 B.n417 10.6151
R1111 B.n417 B.n179 10.6151
R1112 B.n411 B.n179 10.6151
R1113 B.n411 B.n410 10.6151
R1114 B.n410 B.n409 10.6151
R1115 B.n409 B.n181 10.6151
R1116 B.n403 B.n181 10.6151
R1117 B.n403 B.n402 10.6151
R1118 B.n402 B.n401 10.6151
R1119 B.n401 B.n183 10.6151
R1120 B.n395 B.n183 10.6151
R1121 B.n395 B.n394 10.6151
R1122 B.n394 B.n393 10.6151
R1123 B.n393 B.n185 10.6151
R1124 B.n387 B.n185 10.6151
R1125 B.n387 B.n386 10.6151
R1126 B.n386 B.n385 10.6151
R1127 B.n385 B.n187 10.6151
R1128 B.n379 B.n187 10.6151
R1129 B.n379 B.n378 10.6151
R1130 B.n378 B.n377 10.6151
R1131 B.n377 B.n189 10.6151
R1132 B.n371 B.n189 10.6151
R1133 B.n371 B.n370 10.6151
R1134 B.n370 B.n369 10.6151
R1135 B.n369 B.n191 10.6151
R1136 B.n363 B.n191 10.6151
R1137 B.n363 B.n362 10.6151
R1138 B.n362 B.n361 10.6151
R1139 B.n361 B.n193 10.6151
R1140 B.n355 B.n193 10.6151
R1141 B.n355 B.n354 10.6151
R1142 B.n354 B.n353 10.6151
R1143 B.n353 B.n195 10.6151
R1144 B.n347 B.n195 10.6151
R1145 B.n347 B.n346 10.6151
R1146 B.n346 B.n345 10.6151
R1147 B.n345 B.n197 10.6151
R1148 B.n339 B.n338 10.6151
R1149 B.n338 B.n337 10.6151
R1150 B.n337 B.n202 10.6151
R1151 B.n331 B.n202 10.6151
R1152 B.n331 B.n330 10.6151
R1153 B.n330 B.n329 10.6151
R1154 B.n329 B.n204 10.6151
R1155 B.n323 B.n204 10.6151
R1156 B.n323 B.n322 10.6151
R1157 B.n320 B.n208 10.6151
R1158 B.n314 B.n208 10.6151
R1159 B.n314 B.n313 10.6151
R1160 B.n313 B.n312 10.6151
R1161 B.n312 B.n210 10.6151
R1162 B.n306 B.n210 10.6151
R1163 B.n306 B.n305 10.6151
R1164 B.n305 B.n304 10.6151
R1165 B.n304 B.n212 10.6151
R1166 B.n298 B.n212 10.6151
R1167 B.n298 B.n297 10.6151
R1168 B.n297 B.n296 10.6151
R1169 B.n296 B.n214 10.6151
R1170 B.n290 B.n214 10.6151
R1171 B.n290 B.n289 10.6151
R1172 B.n289 B.n288 10.6151
R1173 B.n288 B.n216 10.6151
R1174 B.n282 B.n216 10.6151
R1175 B.n282 B.n281 10.6151
R1176 B.n281 B.n280 10.6151
R1177 B.n280 B.n218 10.6151
R1178 B.n274 B.n218 10.6151
R1179 B.n274 B.n273 10.6151
R1180 B.n273 B.n272 10.6151
R1181 B.n272 B.n220 10.6151
R1182 B.n266 B.n220 10.6151
R1183 B.n266 B.n265 10.6151
R1184 B.n265 B.n264 10.6151
R1185 B.n264 B.n222 10.6151
R1186 B.n258 B.n222 10.6151
R1187 B.n258 B.n257 10.6151
R1188 B.n257 B.n256 10.6151
R1189 B.n256 B.n224 10.6151
R1190 B.n250 B.n224 10.6151
R1191 B.n250 B.n249 10.6151
R1192 B.n249 B.n248 10.6151
R1193 B.n248 B.n226 10.6151
R1194 B.n242 B.n226 10.6151
R1195 B.n242 B.n241 10.6151
R1196 B.n241 B.n240 10.6151
R1197 B.n240 B.n228 10.6151
R1198 B.n234 B.n228 10.6151
R1199 B.n234 B.n233 10.6151
R1200 B.n233 B.n232 10.6151
R1201 B.n232 B.n171 10.6151
R1202 B.n437 B.n436 10.6151
R1203 B.n438 B.n437 10.6151
R1204 B.n438 B.n163 10.6151
R1205 B.n448 B.n163 10.6151
R1206 B.n449 B.n448 10.6151
R1207 B.n450 B.n449 10.6151
R1208 B.n450 B.n155 10.6151
R1209 B.n460 B.n155 10.6151
R1210 B.n461 B.n460 10.6151
R1211 B.n462 B.n461 10.6151
R1212 B.n462 B.n147 10.6151
R1213 B.n472 B.n147 10.6151
R1214 B.n473 B.n472 10.6151
R1215 B.n474 B.n473 10.6151
R1216 B.n474 B.n139 10.6151
R1217 B.n484 B.n139 10.6151
R1218 B.n485 B.n484 10.6151
R1219 B.n486 B.n485 10.6151
R1220 B.n486 B.n131 10.6151
R1221 B.n496 B.n131 10.6151
R1222 B.n497 B.n496 10.6151
R1223 B.n498 B.n497 10.6151
R1224 B.n498 B.n124 10.6151
R1225 B.n509 B.n124 10.6151
R1226 B.n510 B.n509 10.6151
R1227 B.n512 B.n510 10.6151
R1228 B.n512 B.n511 10.6151
R1229 B.n511 B.n116 10.6151
R1230 B.n523 B.n116 10.6151
R1231 B.n524 B.n523 10.6151
R1232 B.n525 B.n524 10.6151
R1233 B.n526 B.n525 10.6151
R1234 B.n527 B.n526 10.6151
R1235 B.n530 B.n527 10.6151
R1236 B.n531 B.n530 10.6151
R1237 B.n532 B.n531 10.6151
R1238 B.n533 B.n532 10.6151
R1239 B.n535 B.n533 10.6151
R1240 B.n536 B.n535 10.6151
R1241 B.n537 B.n536 10.6151
R1242 B.n538 B.n537 10.6151
R1243 B.n540 B.n538 10.6151
R1244 B.n541 B.n540 10.6151
R1245 B.n542 B.n541 10.6151
R1246 B.n543 B.n542 10.6151
R1247 B.n545 B.n543 10.6151
R1248 B.n546 B.n545 10.6151
R1249 B.n547 B.n546 10.6151
R1250 B.n548 B.n547 10.6151
R1251 B.n550 B.n548 10.6151
R1252 B.n551 B.n550 10.6151
R1253 B.n552 B.n551 10.6151
R1254 B.n553 B.n552 10.6151
R1255 B.n555 B.n553 10.6151
R1256 B.n556 B.n555 10.6151
R1257 B.n557 B.n556 10.6151
R1258 B.n558 B.n557 10.6151
R1259 B.n560 B.n558 10.6151
R1260 B.n561 B.n560 10.6151
R1261 B.n562 B.n561 10.6151
R1262 B.n563 B.n562 10.6151
R1263 B.n824 B.n1 10.6151
R1264 B.n824 B.n823 10.6151
R1265 B.n823 B.n822 10.6151
R1266 B.n822 B.n10 10.6151
R1267 B.n816 B.n10 10.6151
R1268 B.n816 B.n815 10.6151
R1269 B.n815 B.n814 10.6151
R1270 B.n814 B.n17 10.6151
R1271 B.n808 B.n17 10.6151
R1272 B.n808 B.n807 10.6151
R1273 B.n807 B.n806 10.6151
R1274 B.n806 B.n25 10.6151
R1275 B.n800 B.n25 10.6151
R1276 B.n800 B.n799 10.6151
R1277 B.n799 B.n798 10.6151
R1278 B.n798 B.n32 10.6151
R1279 B.n792 B.n32 10.6151
R1280 B.n792 B.n791 10.6151
R1281 B.n791 B.n790 10.6151
R1282 B.n790 B.n39 10.6151
R1283 B.n784 B.n39 10.6151
R1284 B.n784 B.n783 10.6151
R1285 B.n783 B.n782 10.6151
R1286 B.n782 B.n46 10.6151
R1287 B.n776 B.n46 10.6151
R1288 B.n776 B.n775 10.6151
R1289 B.n775 B.n774 10.6151
R1290 B.n774 B.n53 10.6151
R1291 B.n768 B.n53 10.6151
R1292 B.n767 B.n766 10.6151
R1293 B.n766 B.n60 10.6151
R1294 B.n760 B.n60 10.6151
R1295 B.n760 B.n759 10.6151
R1296 B.n759 B.n758 10.6151
R1297 B.n758 B.n62 10.6151
R1298 B.n752 B.n62 10.6151
R1299 B.n752 B.n751 10.6151
R1300 B.n751 B.n750 10.6151
R1301 B.n750 B.n64 10.6151
R1302 B.n744 B.n64 10.6151
R1303 B.n744 B.n743 10.6151
R1304 B.n743 B.n742 10.6151
R1305 B.n742 B.n66 10.6151
R1306 B.n736 B.n66 10.6151
R1307 B.n736 B.n735 10.6151
R1308 B.n735 B.n734 10.6151
R1309 B.n734 B.n68 10.6151
R1310 B.n728 B.n68 10.6151
R1311 B.n728 B.n727 10.6151
R1312 B.n727 B.n726 10.6151
R1313 B.n726 B.n70 10.6151
R1314 B.n720 B.n70 10.6151
R1315 B.n720 B.n719 10.6151
R1316 B.n719 B.n718 10.6151
R1317 B.n718 B.n72 10.6151
R1318 B.n712 B.n72 10.6151
R1319 B.n712 B.n711 10.6151
R1320 B.n711 B.n710 10.6151
R1321 B.n710 B.n74 10.6151
R1322 B.n704 B.n74 10.6151
R1323 B.n704 B.n703 10.6151
R1324 B.n703 B.n702 10.6151
R1325 B.n702 B.n76 10.6151
R1326 B.n696 B.n76 10.6151
R1327 B.n696 B.n695 10.6151
R1328 B.n695 B.n694 10.6151
R1329 B.n694 B.n78 10.6151
R1330 B.n688 B.n78 10.6151
R1331 B.n688 B.n687 10.6151
R1332 B.n687 B.n686 10.6151
R1333 B.n686 B.n80 10.6151
R1334 B.n680 B.n80 10.6151
R1335 B.n680 B.n679 10.6151
R1336 B.n679 B.n678 10.6151
R1337 B.n674 B.n673 10.6151
R1338 B.n673 B.n86 10.6151
R1339 B.n668 B.n86 10.6151
R1340 B.n668 B.n667 10.6151
R1341 B.n667 B.n666 10.6151
R1342 B.n666 B.n88 10.6151
R1343 B.n660 B.n88 10.6151
R1344 B.n660 B.n659 10.6151
R1345 B.n659 B.n658 10.6151
R1346 B.n654 B.n653 10.6151
R1347 B.n653 B.n94 10.6151
R1348 B.n648 B.n94 10.6151
R1349 B.n648 B.n647 10.6151
R1350 B.n647 B.n646 10.6151
R1351 B.n646 B.n96 10.6151
R1352 B.n640 B.n96 10.6151
R1353 B.n640 B.n639 10.6151
R1354 B.n639 B.n638 10.6151
R1355 B.n638 B.n98 10.6151
R1356 B.n632 B.n98 10.6151
R1357 B.n632 B.n631 10.6151
R1358 B.n631 B.n630 10.6151
R1359 B.n630 B.n100 10.6151
R1360 B.n624 B.n100 10.6151
R1361 B.n624 B.n623 10.6151
R1362 B.n623 B.n622 10.6151
R1363 B.n622 B.n102 10.6151
R1364 B.n616 B.n102 10.6151
R1365 B.n616 B.n615 10.6151
R1366 B.n615 B.n614 10.6151
R1367 B.n614 B.n104 10.6151
R1368 B.n608 B.n104 10.6151
R1369 B.n608 B.n607 10.6151
R1370 B.n607 B.n606 10.6151
R1371 B.n606 B.n106 10.6151
R1372 B.n600 B.n106 10.6151
R1373 B.n600 B.n599 10.6151
R1374 B.n599 B.n598 10.6151
R1375 B.n598 B.n108 10.6151
R1376 B.n592 B.n108 10.6151
R1377 B.n592 B.n591 10.6151
R1378 B.n591 B.n590 10.6151
R1379 B.n590 B.n110 10.6151
R1380 B.n584 B.n110 10.6151
R1381 B.n584 B.n583 10.6151
R1382 B.n583 B.n582 10.6151
R1383 B.n582 B.n112 10.6151
R1384 B.n576 B.n112 10.6151
R1385 B.n576 B.n575 10.6151
R1386 B.n575 B.n574 10.6151
R1387 B.n574 B.n114 10.6151
R1388 B.n568 B.n114 10.6151
R1389 B.n568 B.n567 10.6151
R1390 B.n567 B.n566 10.6151
R1391 B.n201 B.n197 9.36635
R1392 B.n321 B.n320 9.36635
R1393 B.n678 B.n84 9.36635
R1394 B.n654 B.n92 9.36635
R1395 B.n832 B.n0 8.11757
R1396 B.n832 B.n1 8.11757
R1397 B.t6 B.n153 4.65043
R1398 B.n787 B.t2 4.65043
R1399 B.n339 B.n201 1.24928
R1400 B.n322 B.n321 1.24928
R1401 B.n674 B.n84 1.24928
R1402 B.n658 B.n92 1.24928
R1403 VN VN.t0 181.465
R1404 VN VN.t1 133.845
R1405 VTAIL.n1 VTAIL.t2 47.5843
R1406 VTAIL.n3 VTAIL.t3 47.5841
R1407 VTAIL.n0 VTAIL.t0 47.5841
R1408 VTAIL.n2 VTAIL.t1 47.5841
R1409 VTAIL.n1 VTAIL.n0 30.7031
R1410 VTAIL.n3 VTAIL.n2 27.4186
R1411 VTAIL.n2 VTAIL.n1 2.11257
R1412 VTAIL VTAIL.n0 1.34964
R1413 VTAIL VTAIL.n3 0.763431
R1414 VDD2.n0 VDD2.t0 106.258
R1415 VDD2.n0 VDD2.t1 64.2629
R1416 VDD2 VDD2.n0 0.87981
R1417 VP.n0 VP.t0 181.559
R1418 VP.n0 VP.t1 133.319
R1419 VP VP.n0 0.52637
R1420 VDD1 VDD1.t0 107.605
R1421 VDD1 VDD1.t1 65.1422
C0 VTAIL VDD1 5.65159f
C1 VP VDD2 0.370145f
C2 VP VN 6.17326f
C3 VDD2 VN 3.25436f
C4 VP VDD1 3.47358f
C5 VDD1 VDD2 0.782243f
C6 VDD1 VN 0.148526f
C7 VP VTAIL 2.9134f
C8 VTAIL VDD2 5.70858f
C9 VTAIL VN 2.89915f
C10 VDD2 B 5.032715f
C11 VDD1 B 8.49076f
C12 VTAIL B 8.460104f
C13 VN B 11.97076f
C14 VP B 7.598394f
C15 VDD1.t1 B 2.56263f
C16 VDD1.t0 B 3.24124f
C17 VP.t0 B 4.44083f
C18 VP.t1 B 3.77159f
C19 VP.n0 B 4.29127f
C20 VDD2.t0 B 3.1538f
C21 VDD2.t1 B 2.52405f
C22 VDD2.n0 B 3.15611f
C23 VTAIL.t0 B 2.49324f
C24 VTAIL.n0 B 1.8655f
C25 VTAIL.t2 B 2.49324f
C26 VTAIL.n1 B 1.91646f
C27 VTAIL.t1 B 2.49324f
C28 VTAIL.n2 B 1.69706f
C29 VTAIL.t3 B 2.49324f
C30 VTAIL.n3 B 1.60694f
C31 VN.t1 B 3.70548f
C32 VN.t0 B 4.35759f
.ends

