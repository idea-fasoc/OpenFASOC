* NGSPICE file created from diff_pair_sample_0544.ext - technology: sky130A

.subckt diff_pair_sample_0544 VTAIL VN VP B VDD2 VDD1
X0 B.t11 B.t9 B.t10 w_n2308_n4336# sky130_fd_pr__pfet_01v8 ad=6.5676 pd=34.46 as=0 ps=0 w=16.84 l=1.9
X1 B.t8 B.t6 B.t7 w_n2308_n4336# sky130_fd_pr__pfet_01v8 ad=6.5676 pd=34.46 as=0 ps=0 w=16.84 l=1.9
X2 VDD2.t3 VN.t0 VTAIL.t7 w_n2308_n4336# sky130_fd_pr__pfet_01v8 ad=2.7786 pd=17.17 as=6.5676 ps=34.46 w=16.84 l=1.9
X3 VTAIL.t6 VN.t1 VDD2.t2 w_n2308_n4336# sky130_fd_pr__pfet_01v8 ad=6.5676 pd=34.46 as=2.7786 ps=17.17 w=16.84 l=1.9
X4 VTAIL.t5 VN.t2 VDD2.t1 w_n2308_n4336# sky130_fd_pr__pfet_01v8 ad=6.5676 pd=34.46 as=2.7786 ps=17.17 w=16.84 l=1.9
X5 VDD2.t0 VN.t3 VTAIL.t4 w_n2308_n4336# sky130_fd_pr__pfet_01v8 ad=2.7786 pd=17.17 as=6.5676 ps=34.46 w=16.84 l=1.9
X6 B.t5 B.t3 B.t4 w_n2308_n4336# sky130_fd_pr__pfet_01v8 ad=6.5676 pd=34.46 as=0 ps=0 w=16.84 l=1.9
X7 VDD1.t3 VP.t0 VTAIL.t1 w_n2308_n4336# sky130_fd_pr__pfet_01v8 ad=2.7786 pd=17.17 as=6.5676 ps=34.46 w=16.84 l=1.9
X8 VTAIL.t2 VP.t1 VDD1.t2 w_n2308_n4336# sky130_fd_pr__pfet_01v8 ad=6.5676 pd=34.46 as=2.7786 ps=17.17 w=16.84 l=1.9
X9 VTAIL.t3 VP.t2 VDD1.t1 w_n2308_n4336# sky130_fd_pr__pfet_01v8 ad=6.5676 pd=34.46 as=2.7786 ps=17.17 w=16.84 l=1.9
X10 VDD1.t0 VP.t3 VTAIL.t0 w_n2308_n4336# sky130_fd_pr__pfet_01v8 ad=2.7786 pd=17.17 as=6.5676 ps=34.46 w=16.84 l=1.9
X11 B.t2 B.t0 B.t1 w_n2308_n4336# sky130_fd_pr__pfet_01v8 ad=6.5676 pd=34.46 as=0 ps=0 w=16.84 l=1.9
R0 B.n408 B.n407 585
R1 B.n406 B.n109 585
R2 B.n405 B.n404 585
R3 B.n403 B.n110 585
R4 B.n402 B.n401 585
R5 B.n400 B.n111 585
R6 B.n399 B.n398 585
R7 B.n397 B.n112 585
R8 B.n396 B.n395 585
R9 B.n394 B.n113 585
R10 B.n393 B.n392 585
R11 B.n391 B.n114 585
R12 B.n390 B.n389 585
R13 B.n388 B.n115 585
R14 B.n387 B.n386 585
R15 B.n385 B.n116 585
R16 B.n384 B.n383 585
R17 B.n382 B.n117 585
R18 B.n381 B.n380 585
R19 B.n379 B.n118 585
R20 B.n378 B.n377 585
R21 B.n376 B.n119 585
R22 B.n375 B.n374 585
R23 B.n373 B.n120 585
R24 B.n372 B.n371 585
R25 B.n370 B.n121 585
R26 B.n369 B.n368 585
R27 B.n367 B.n122 585
R28 B.n366 B.n365 585
R29 B.n364 B.n123 585
R30 B.n363 B.n362 585
R31 B.n361 B.n124 585
R32 B.n360 B.n359 585
R33 B.n358 B.n125 585
R34 B.n357 B.n356 585
R35 B.n355 B.n126 585
R36 B.n354 B.n353 585
R37 B.n352 B.n127 585
R38 B.n351 B.n350 585
R39 B.n349 B.n128 585
R40 B.n348 B.n347 585
R41 B.n346 B.n129 585
R42 B.n345 B.n344 585
R43 B.n343 B.n130 585
R44 B.n342 B.n341 585
R45 B.n340 B.n131 585
R46 B.n339 B.n338 585
R47 B.n337 B.n132 585
R48 B.n336 B.n335 585
R49 B.n334 B.n133 585
R50 B.n333 B.n332 585
R51 B.n331 B.n134 585
R52 B.n330 B.n329 585
R53 B.n328 B.n135 585
R54 B.n327 B.n326 585
R55 B.n325 B.n136 585
R56 B.n324 B.n323 585
R57 B.n319 B.n137 585
R58 B.n318 B.n317 585
R59 B.n316 B.n138 585
R60 B.n315 B.n314 585
R61 B.n313 B.n139 585
R62 B.n312 B.n311 585
R63 B.n310 B.n140 585
R64 B.n309 B.n308 585
R65 B.n306 B.n141 585
R66 B.n305 B.n304 585
R67 B.n303 B.n144 585
R68 B.n302 B.n301 585
R69 B.n300 B.n145 585
R70 B.n299 B.n298 585
R71 B.n297 B.n146 585
R72 B.n296 B.n295 585
R73 B.n294 B.n147 585
R74 B.n293 B.n292 585
R75 B.n291 B.n148 585
R76 B.n290 B.n289 585
R77 B.n288 B.n149 585
R78 B.n287 B.n286 585
R79 B.n285 B.n150 585
R80 B.n284 B.n283 585
R81 B.n282 B.n151 585
R82 B.n281 B.n280 585
R83 B.n279 B.n152 585
R84 B.n278 B.n277 585
R85 B.n276 B.n153 585
R86 B.n275 B.n274 585
R87 B.n273 B.n154 585
R88 B.n272 B.n271 585
R89 B.n270 B.n155 585
R90 B.n269 B.n268 585
R91 B.n267 B.n156 585
R92 B.n266 B.n265 585
R93 B.n264 B.n157 585
R94 B.n263 B.n262 585
R95 B.n261 B.n158 585
R96 B.n260 B.n259 585
R97 B.n258 B.n159 585
R98 B.n257 B.n256 585
R99 B.n255 B.n160 585
R100 B.n254 B.n253 585
R101 B.n252 B.n161 585
R102 B.n251 B.n250 585
R103 B.n249 B.n162 585
R104 B.n248 B.n247 585
R105 B.n246 B.n163 585
R106 B.n245 B.n244 585
R107 B.n243 B.n164 585
R108 B.n242 B.n241 585
R109 B.n240 B.n165 585
R110 B.n239 B.n238 585
R111 B.n237 B.n166 585
R112 B.n236 B.n235 585
R113 B.n234 B.n167 585
R114 B.n233 B.n232 585
R115 B.n231 B.n168 585
R116 B.n230 B.n229 585
R117 B.n228 B.n169 585
R118 B.n227 B.n226 585
R119 B.n225 B.n170 585
R120 B.n224 B.n223 585
R121 B.n409 B.n108 585
R122 B.n411 B.n410 585
R123 B.n412 B.n107 585
R124 B.n414 B.n413 585
R125 B.n415 B.n106 585
R126 B.n417 B.n416 585
R127 B.n418 B.n105 585
R128 B.n420 B.n419 585
R129 B.n421 B.n104 585
R130 B.n423 B.n422 585
R131 B.n424 B.n103 585
R132 B.n426 B.n425 585
R133 B.n427 B.n102 585
R134 B.n429 B.n428 585
R135 B.n430 B.n101 585
R136 B.n432 B.n431 585
R137 B.n433 B.n100 585
R138 B.n435 B.n434 585
R139 B.n436 B.n99 585
R140 B.n438 B.n437 585
R141 B.n439 B.n98 585
R142 B.n441 B.n440 585
R143 B.n442 B.n97 585
R144 B.n444 B.n443 585
R145 B.n445 B.n96 585
R146 B.n447 B.n446 585
R147 B.n448 B.n95 585
R148 B.n450 B.n449 585
R149 B.n451 B.n94 585
R150 B.n453 B.n452 585
R151 B.n454 B.n93 585
R152 B.n456 B.n455 585
R153 B.n457 B.n92 585
R154 B.n459 B.n458 585
R155 B.n460 B.n91 585
R156 B.n462 B.n461 585
R157 B.n463 B.n90 585
R158 B.n465 B.n464 585
R159 B.n466 B.n89 585
R160 B.n468 B.n467 585
R161 B.n469 B.n88 585
R162 B.n471 B.n470 585
R163 B.n472 B.n87 585
R164 B.n474 B.n473 585
R165 B.n475 B.n86 585
R166 B.n477 B.n476 585
R167 B.n478 B.n85 585
R168 B.n480 B.n479 585
R169 B.n481 B.n84 585
R170 B.n483 B.n482 585
R171 B.n484 B.n83 585
R172 B.n486 B.n485 585
R173 B.n487 B.n82 585
R174 B.n489 B.n488 585
R175 B.n490 B.n81 585
R176 B.n492 B.n491 585
R177 B.n675 B.n674 585
R178 B.n673 B.n16 585
R179 B.n672 B.n671 585
R180 B.n670 B.n17 585
R181 B.n669 B.n668 585
R182 B.n667 B.n18 585
R183 B.n666 B.n665 585
R184 B.n664 B.n19 585
R185 B.n663 B.n662 585
R186 B.n661 B.n20 585
R187 B.n660 B.n659 585
R188 B.n658 B.n21 585
R189 B.n657 B.n656 585
R190 B.n655 B.n22 585
R191 B.n654 B.n653 585
R192 B.n652 B.n23 585
R193 B.n651 B.n650 585
R194 B.n649 B.n24 585
R195 B.n648 B.n647 585
R196 B.n646 B.n25 585
R197 B.n645 B.n644 585
R198 B.n643 B.n26 585
R199 B.n642 B.n641 585
R200 B.n640 B.n27 585
R201 B.n639 B.n638 585
R202 B.n637 B.n28 585
R203 B.n636 B.n635 585
R204 B.n634 B.n29 585
R205 B.n633 B.n632 585
R206 B.n631 B.n30 585
R207 B.n630 B.n629 585
R208 B.n628 B.n31 585
R209 B.n627 B.n626 585
R210 B.n625 B.n32 585
R211 B.n624 B.n623 585
R212 B.n622 B.n33 585
R213 B.n621 B.n620 585
R214 B.n619 B.n34 585
R215 B.n618 B.n617 585
R216 B.n616 B.n35 585
R217 B.n615 B.n614 585
R218 B.n613 B.n36 585
R219 B.n612 B.n611 585
R220 B.n610 B.n37 585
R221 B.n609 B.n608 585
R222 B.n607 B.n38 585
R223 B.n606 B.n605 585
R224 B.n604 B.n39 585
R225 B.n603 B.n602 585
R226 B.n601 B.n40 585
R227 B.n600 B.n599 585
R228 B.n598 B.n41 585
R229 B.n597 B.n596 585
R230 B.n595 B.n42 585
R231 B.n594 B.n593 585
R232 B.n592 B.n43 585
R233 B.n590 B.n589 585
R234 B.n588 B.n46 585
R235 B.n587 B.n586 585
R236 B.n585 B.n47 585
R237 B.n584 B.n583 585
R238 B.n582 B.n48 585
R239 B.n581 B.n580 585
R240 B.n579 B.n49 585
R241 B.n578 B.n577 585
R242 B.n576 B.n575 585
R243 B.n574 B.n53 585
R244 B.n573 B.n572 585
R245 B.n571 B.n54 585
R246 B.n570 B.n569 585
R247 B.n568 B.n55 585
R248 B.n567 B.n566 585
R249 B.n565 B.n56 585
R250 B.n564 B.n563 585
R251 B.n562 B.n57 585
R252 B.n561 B.n560 585
R253 B.n559 B.n58 585
R254 B.n558 B.n557 585
R255 B.n556 B.n59 585
R256 B.n555 B.n554 585
R257 B.n553 B.n60 585
R258 B.n552 B.n551 585
R259 B.n550 B.n61 585
R260 B.n549 B.n548 585
R261 B.n547 B.n62 585
R262 B.n546 B.n545 585
R263 B.n544 B.n63 585
R264 B.n543 B.n542 585
R265 B.n541 B.n64 585
R266 B.n540 B.n539 585
R267 B.n538 B.n65 585
R268 B.n537 B.n536 585
R269 B.n535 B.n66 585
R270 B.n534 B.n533 585
R271 B.n532 B.n67 585
R272 B.n531 B.n530 585
R273 B.n529 B.n68 585
R274 B.n528 B.n527 585
R275 B.n526 B.n69 585
R276 B.n525 B.n524 585
R277 B.n523 B.n70 585
R278 B.n522 B.n521 585
R279 B.n520 B.n71 585
R280 B.n519 B.n518 585
R281 B.n517 B.n72 585
R282 B.n516 B.n515 585
R283 B.n514 B.n73 585
R284 B.n513 B.n512 585
R285 B.n511 B.n74 585
R286 B.n510 B.n509 585
R287 B.n508 B.n75 585
R288 B.n507 B.n506 585
R289 B.n505 B.n76 585
R290 B.n504 B.n503 585
R291 B.n502 B.n77 585
R292 B.n501 B.n500 585
R293 B.n499 B.n78 585
R294 B.n498 B.n497 585
R295 B.n496 B.n79 585
R296 B.n495 B.n494 585
R297 B.n493 B.n80 585
R298 B.n676 B.n15 585
R299 B.n678 B.n677 585
R300 B.n679 B.n14 585
R301 B.n681 B.n680 585
R302 B.n682 B.n13 585
R303 B.n684 B.n683 585
R304 B.n685 B.n12 585
R305 B.n687 B.n686 585
R306 B.n688 B.n11 585
R307 B.n690 B.n689 585
R308 B.n691 B.n10 585
R309 B.n693 B.n692 585
R310 B.n694 B.n9 585
R311 B.n696 B.n695 585
R312 B.n697 B.n8 585
R313 B.n699 B.n698 585
R314 B.n700 B.n7 585
R315 B.n702 B.n701 585
R316 B.n703 B.n6 585
R317 B.n705 B.n704 585
R318 B.n706 B.n5 585
R319 B.n708 B.n707 585
R320 B.n709 B.n4 585
R321 B.n711 B.n710 585
R322 B.n712 B.n3 585
R323 B.n714 B.n713 585
R324 B.n715 B.n0 585
R325 B.n2 B.n1 585
R326 B.n185 B.n184 585
R327 B.n186 B.n183 585
R328 B.n188 B.n187 585
R329 B.n189 B.n182 585
R330 B.n191 B.n190 585
R331 B.n192 B.n181 585
R332 B.n194 B.n193 585
R333 B.n195 B.n180 585
R334 B.n197 B.n196 585
R335 B.n198 B.n179 585
R336 B.n200 B.n199 585
R337 B.n201 B.n178 585
R338 B.n203 B.n202 585
R339 B.n204 B.n177 585
R340 B.n206 B.n205 585
R341 B.n207 B.n176 585
R342 B.n209 B.n208 585
R343 B.n210 B.n175 585
R344 B.n212 B.n211 585
R345 B.n213 B.n174 585
R346 B.n215 B.n214 585
R347 B.n216 B.n173 585
R348 B.n218 B.n217 585
R349 B.n219 B.n172 585
R350 B.n221 B.n220 585
R351 B.n222 B.n171 585
R352 B.n224 B.n171 569.379
R353 B.n409 B.n408 569.379
R354 B.n493 B.n492 569.379
R355 B.n674 B.n15 569.379
R356 B.n320 B.t7 506.065
R357 B.n50 B.t5 506.065
R358 B.n142 B.t10 506.065
R359 B.n44 B.t2 506.065
R360 B.n321 B.t8 462.817
R361 B.n51 B.t4 462.817
R362 B.n143 B.t11 462.817
R363 B.n45 B.t1 462.817
R364 B.n142 B.t9 420.276
R365 B.n320 B.t6 420.276
R366 B.n50 B.t3 420.276
R367 B.n44 B.t0 420.276
R368 B.n717 B.n716 256.663
R369 B.n716 B.n715 235.042
R370 B.n716 B.n2 235.042
R371 B.n225 B.n224 163.367
R372 B.n226 B.n225 163.367
R373 B.n226 B.n169 163.367
R374 B.n230 B.n169 163.367
R375 B.n231 B.n230 163.367
R376 B.n232 B.n231 163.367
R377 B.n232 B.n167 163.367
R378 B.n236 B.n167 163.367
R379 B.n237 B.n236 163.367
R380 B.n238 B.n237 163.367
R381 B.n238 B.n165 163.367
R382 B.n242 B.n165 163.367
R383 B.n243 B.n242 163.367
R384 B.n244 B.n243 163.367
R385 B.n244 B.n163 163.367
R386 B.n248 B.n163 163.367
R387 B.n249 B.n248 163.367
R388 B.n250 B.n249 163.367
R389 B.n250 B.n161 163.367
R390 B.n254 B.n161 163.367
R391 B.n255 B.n254 163.367
R392 B.n256 B.n255 163.367
R393 B.n256 B.n159 163.367
R394 B.n260 B.n159 163.367
R395 B.n261 B.n260 163.367
R396 B.n262 B.n261 163.367
R397 B.n262 B.n157 163.367
R398 B.n266 B.n157 163.367
R399 B.n267 B.n266 163.367
R400 B.n268 B.n267 163.367
R401 B.n268 B.n155 163.367
R402 B.n272 B.n155 163.367
R403 B.n273 B.n272 163.367
R404 B.n274 B.n273 163.367
R405 B.n274 B.n153 163.367
R406 B.n278 B.n153 163.367
R407 B.n279 B.n278 163.367
R408 B.n280 B.n279 163.367
R409 B.n280 B.n151 163.367
R410 B.n284 B.n151 163.367
R411 B.n285 B.n284 163.367
R412 B.n286 B.n285 163.367
R413 B.n286 B.n149 163.367
R414 B.n290 B.n149 163.367
R415 B.n291 B.n290 163.367
R416 B.n292 B.n291 163.367
R417 B.n292 B.n147 163.367
R418 B.n296 B.n147 163.367
R419 B.n297 B.n296 163.367
R420 B.n298 B.n297 163.367
R421 B.n298 B.n145 163.367
R422 B.n302 B.n145 163.367
R423 B.n303 B.n302 163.367
R424 B.n304 B.n303 163.367
R425 B.n304 B.n141 163.367
R426 B.n309 B.n141 163.367
R427 B.n310 B.n309 163.367
R428 B.n311 B.n310 163.367
R429 B.n311 B.n139 163.367
R430 B.n315 B.n139 163.367
R431 B.n316 B.n315 163.367
R432 B.n317 B.n316 163.367
R433 B.n317 B.n137 163.367
R434 B.n324 B.n137 163.367
R435 B.n325 B.n324 163.367
R436 B.n326 B.n325 163.367
R437 B.n326 B.n135 163.367
R438 B.n330 B.n135 163.367
R439 B.n331 B.n330 163.367
R440 B.n332 B.n331 163.367
R441 B.n332 B.n133 163.367
R442 B.n336 B.n133 163.367
R443 B.n337 B.n336 163.367
R444 B.n338 B.n337 163.367
R445 B.n338 B.n131 163.367
R446 B.n342 B.n131 163.367
R447 B.n343 B.n342 163.367
R448 B.n344 B.n343 163.367
R449 B.n344 B.n129 163.367
R450 B.n348 B.n129 163.367
R451 B.n349 B.n348 163.367
R452 B.n350 B.n349 163.367
R453 B.n350 B.n127 163.367
R454 B.n354 B.n127 163.367
R455 B.n355 B.n354 163.367
R456 B.n356 B.n355 163.367
R457 B.n356 B.n125 163.367
R458 B.n360 B.n125 163.367
R459 B.n361 B.n360 163.367
R460 B.n362 B.n361 163.367
R461 B.n362 B.n123 163.367
R462 B.n366 B.n123 163.367
R463 B.n367 B.n366 163.367
R464 B.n368 B.n367 163.367
R465 B.n368 B.n121 163.367
R466 B.n372 B.n121 163.367
R467 B.n373 B.n372 163.367
R468 B.n374 B.n373 163.367
R469 B.n374 B.n119 163.367
R470 B.n378 B.n119 163.367
R471 B.n379 B.n378 163.367
R472 B.n380 B.n379 163.367
R473 B.n380 B.n117 163.367
R474 B.n384 B.n117 163.367
R475 B.n385 B.n384 163.367
R476 B.n386 B.n385 163.367
R477 B.n386 B.n115 163.367
R478 B.n390 B.n115 163.367
R479 B.n391 B.n390 163.367
R480 B.n392 B.n391 163.367
R481 B.n392 B.n113 163.367
R482 B.n396 B.n113 163.367
R483 B.n397 B.n396 163.367
R484 B.n398 B.n397 163.367
R485 B.n398 B.n111 163.367
R486 B.n402 B.n111 163.367
R487 B.n403 B.n402 163.367
R488 B.n404 B.n403 163.367
R489 B.n404 B.n109 163.367
R490 B.n408 B.n109 163.367
R491 B.n492 B.n81 163.367
R492 B.n488 B.n81 163.367
R493 B.n488 B.n487 163.367
R494 B.n487 B.n486 163.367
R495 B.n486 B.n83 163.367
R496 B.n482 B.n83 163.367
R497 B.n482 B.n481 163.367
R498 B.n481 B.n480 163.367
R499 B.n480 B.n85 163.367
R500 B.n476 B.n85 163.367
R501 B.n476 B.n475 163.367
R502 B.n475 B.n474 163.367
R503 B.n474 B.n87 163.367
R504 B.n470 B.n87 163.367
R505 B.n470 B.n469 163.367
R506 B.n469 B.n468 163.367
R507 B.n468 B.n89 163.367
R508 B.n464 B.n89 163.367
R509 B.n464 B.n463 163.367
R510 B.n463 B.n462 163.367
R511 B.n462 B.n91 163.367
R512 B.n458 B.n91 163.367
R513 B.n458 B.n457 163.367
R514 B.n457 B.n456 163.367
R515 B.n456 B.n93 163.367
R516 B.n452 B.n93 163.367
R517 B.n452 B.n451 163.367
R518 B.n451 B.n450 163.367
R519 B.n450 B.n95 163.367
R520 B.n446 B.n95 163.367
R521 B.n446 B.n445 163.367
R522 B.n445 B.n444 163.367
R523 B.n444 B.n97 163.367
R524 B.n440 B.n97 163.367
R525 B.n440 B.n439 163.367
R526 B.n439 B.n438 163.367
R527 B.n438 B.n99 163.367
R528 B.n434 B.n99 163.367
R529 B.n434 B.n433 163.367
R530 B.n433 B.n432 163.367
R531 B.n432 B.n101 163.367
R532 B.n428 B.n101 163.367
R533 B.n428 B.n427 163.367
R534 B.n427 B.n426 163.367
R535 B.n426 B.n103 163.367
R536 B.n422 B.n103 163.367
R537 B.n422 B.n421 163.367
R538 B.n421 B.n420 163.367
R539 B.n420 B.n105 163.367
R540 B.n416 B.n105 163.367
R541 B.n416 B.n415 163.367
R542 B.n415 B.n414 163.367
R543 B.n414 B.n107 163.367
R544 B.n410 B.n107 163.367
R545 B.n410 B.n409 163.367
R546 B.n674 B.n673 163.367
R547 B.n673 B.n672 163.367
R548 B.n672 B.n17 163.367
R549 B.n668 B.n17 163.367
R550 B.n668 B.n667 163.367
R551 B.n667 B.n666 163.367
R552 B.n666 B.n19 163.367
R553 B.n662 B.n19 163.367
R554 B.n662 B.n661 163.367
R555 B.n661 B.n660 163.367
R556 B.n660 B.n21 163.367
R557 B.n656 B.n21 163.367
R558 B.n656 B.n655 163.367
R559 B.n655 B.n654 163.367
R560 B.n654 B.n23 163.367
R561 B.n650 B.n23 163.367
R562 B.n650 B.n649 163.367
R563 B.n649 B.n648 163.367
R564 B.n648 B.n25 163.367
R565 B.n644 B.n25 163.367
R566 B.n644 B.n643 163.367
R567 B.n643 B.n642 163.367
R568 B.n642 B.n27 163.367
R569 B.n638 B.n27 163.367
R570 B.n638 B.n637 163.367
R571 B.n637 B.n636 163.367
R572 B.n636 B.n29 163.367
R573 B.n632 B.n29 163.367
R574 B.n632 B.n631 163.367
R575 B.n631 B.n630 163.367
R576 B.n630 B.n31 163.367
R577 B.n626 B.n31 163.367
R578 B.n626 B.n625 163.367
R579 B.n625 B.n624 163.367
R580 B.n624 B.n33 163.367
R581 B.n620 B.n33 163.367
R582 B.n620 B.n619 163.367
R583 B.n619 B.n618 163.367
R584 B.n618 B.n35 163.367
R585 B.n614 B.n35 163.367
R586 B.n614 B.n613 163.367
R587 B.n613 B.n612 163.367
R588 B.n612 B.n37 163.367
R589 B.n608 B.n37 163.367
R590 B.n608 B.n607 163.367
R591 B.n607 B.n606 163.367
R592 B.n606 B.n39 163.367
R593 B.n602 B.n39 163.367
R594 B.n602 B.n601 163.367
R595 B.n601 B.n600 163.367
R596 B.n600 B.n41 163.367
R597 B.n596 B.n41 163.367
R598 B.n596 B.n595 163.367
R599 B.n595 B.n594 163.367
R600 B.n594 B.n43 163.367
R601 B.n589 B.n43 163.367
R602 B.n589 B.n588 163.367
R603 B.n588 B.n587 163.367
R604 B.n587 B.n47 163.367
R605 B.n583 B.n47 163.367
R606 B.n583 B.n582 163.367
R607 B.n582 B.n581 163.367
R608 B.n581 B.n49 163.367
R609 B.n577 B.n49 163.367
R610 B.n577 B.n576 163.367
R611 B.n576 B.n53 163.367
R612 B.n572 B.n53 163.367
R613 B.n572 B.n571 163.367
R614 B.n571 B.n570 163.367
R615 B.n570 B.n55 163.367
R616 B.n566 B.n55 163.367
R617 B.n566 B.n565 163.367
R618 B.n565 B.n564 163.367
R619 B.n564 B.n57 163.367
R620 B.n560 B.n57 163.367
R621 B.n560 B.n559 163.367
R622 B.n559 B.n558 163.367
R623 B.n558 B.n59 163.367
R624 B.n554 B.n59 163.367
R625 B.n554 B.n553 163.367
R626 B.n553 B.n552 163.367
R627 B.n552 B.n61 163.367
R628 B.n548 B.n61 163.367
R629 B.n548 B.n547 163.367
R630 B.n547 B.n546 163.367
R631 B.n546 B.n63 163.367
R632 B.n542 B.n63 163.367
R633 B.n542 B.n541 163.367
R634 B.n541 B.n540 163.367
R635 B.n540 B.n65 163.367
R636 B.n536 B.n65 163.367
R637 B.n536 B.n535 163.367
R638 B.n535 B.n534 163.367
R639 B.n534 B.n67 163.367
R640 B.n530 B.n67 163.367
R641 B.n530 B.n529 163.367
R642 B.n529 B.n528 163.367
R643 B.n528 B.n69 163.367
R644 B.n524 B.n69 163.367
R645 B.n524 B.n523 163.367
R646 B.n523 B.n522 163.367
R647 B.n522 B.n71 163.367
R648 B.n518 B.n71 163.367
R649 B.n518 B.n517 163.367
R650 B.n517 B.n516 163.367
R651 B.n516 B.n73 163.367
R652 B.n512 B.n73 163.367
R653 B.n512 B.n511 163.367
R654 B.n511 B.n510 163.367
R655 B.n510 B.n75 163.367
R656 B.n506 B.n75 163.367
R657 B.n506 B.n505 163.367
R658 B.n505 B.n504 163.367
R659 B.n504 B.n77 163.367
R660 B.n500 B.n77 163.367
R661 B.n500 B.n499 163.367
R662 B.n499 B.n498 163.367
R663 B.n498 B.n79 163.367
R664 B.n494 B.n79 163.367
R665 B.n494 B.n493 163.367
R666 B.n678 B.n15 163.367
R667 B.n679 B.n678 163.367
R668 B.n680 B.n679 163.367
R669 B.n680 B.n13 163.367
R670 B.n684 B.n13 163.367
R671 B.n685 B.n684 163.367
R672 B.n686 B.n685 163.367
R673 B.n686 B.n11 163.367
R674 B.n690 B.n11 163.367
R675 B.n691 B.n690 163.367
R676 B.n692 B.n691 163.367
R677 B.n692 B.n9 163.367
R678 B.n696 B.n9 163.367
R679 B.n697 B.n696 163.367
R680 B.n698 B.n697 163.367
R681 B.n698 B.n7 163.367
R682 B.n702 B.n7 163.367
R683 B.n703 B.n702 163.367
R684 B.n704 B.n703 163.367
R685 B.n704 B.n5 163.367
R686 B.n708 B.n5 163.367
R687 B.n709 B.n708 163.367
R688 B.n710 B.n709 163.367
R689 B.n710 B.n3 163.367
R690 B.n714 B.n3 163.367
R691 B.n715 B.n714 163.367
R692 B.n184 B.n2 163.367
R693 B.n184 B.n183 163.367
R694 B.n188 B.n183 163.367
R695 B.n189 B.n188 163.367
R696 B.n190 B.n189 163.367
R697 B.n190 B.n181 163.367
R698 B.n194 B.n181 163.367
R699 B.n195 B.n194 163.367
R700 B.n196 B.n195 163.367
R701 B.n196 B.n179 163.367
R702 B.n200 B.n179 163.367
R703 B.n201 B.n200 163.367
R704 B.n202 B.n201 163.367
R705 B.n202 B.n177 163.367
R706 B.n206 B.n177 163.367
R707 B.n207 B.n206 163.367
R708 B.n208 B.n207 163.367
R709 B.n208 B.n175 163.367
R710 B.n212 B.n175 163.367
R711 B.n213 B.n212 163.367
R712 B.n214 B.n213 163.367
R713 B.n214 B.n173 163.367
R714 B.n218 B.n173 163.367
R715 B.n219 B.n218 163.367
R716 B.n220 B.n219 163.367
R717 B.n220 B.n171 163.367
R718 B.n307 B.n143 59.5399
R719 B.n322 B.n321 59.5399
R720 B.n52 B.n51 59.5399
R721 B.n591 B.n45 59.5399
R722 B.n143 B.n142 43.249
R723 B.n321 B.n320 43.249
R724 B.n51 B.n50 43.249
R725 B.n45 B.n44 43.249
R726 B.n676 B.n675 36.9956
R727 B.n491 B.n80 36.9956
R728 B.n407 B.n108 36.9956
R729 B.n223 B.n222 36.9956
R730 B B.n717 18.0485
R731 B.n677 B.n676 10.6151
R732 B.n677 B.n14 10.6151
R733 B.n681 B.n14 10.6151
R734 B.n682 B.n681 10.6151
R735 B.n683 B.n682 10.6151
R736 B.n683 B.n12 10.6151
R737 B.n687 B.n12 10.6151
R738 B.n688 B.n687 10.6151
R739 B.n689 B.n688 10.6151
R740 B.n689 B.n10 10.6151
R741 B.n693 B.n10 10.6151
R742 B.n694 B.n693 10.6151
R743 B.n695 B.n694 10.6151
R744 B.n695 B.n8 10.6151
R745 B.n699 B.n8 10.6151
R746 B.n700 B.n699 10.6151
R747 B.n701 B.n700 10.6151
R748 B.n701 B.n6 10.6151
R749 B.n705 B.n6 10.6151
R750 B.n706 B.n705 10.6151
R751 B.n707 B.n706 10.6151
R752 B.n707 B.n4 10.6151
R753 B.n711 B.n4 10.6151
R754 B.n712 B.n711 10.6151
R755 B.n713 B.n712 10.6151
R756 B.n713 B.n0 10.6151
R757 B.n675 B.n16 10.6151
R758 B.n671 B.n16 10.6151
R759 B.n671 B.n670 10.6151
R760 B.n670 B.n669 10.6151
R761 B.n669 B.n18 10.6151
R762 B.n665 B.n18 10.6151
R763 B.n665 B.n664 10.6151
R764 B.n664 B.n663 10.6151
R765 B.n663 B.n20 10.6151
R766 B.n659 B.n20 10.6151
R767 B.n659 B.n658 10.6151
R768 B.n658 B.n657 10.6151
R769 B.n657 B.n22 10.6151
R770 B.n653 B.n22 10.6151
R771 B.n653 B.n652 10.6151
R772 B.n652 B.n651 10.6151
R773 B.n651 B.n24 10.6151
R774 B.n647 B.n24 10.6151
R775 B.n647 B.n646 10.6151
R776 B.n646 B.n645 10.6151
R777 B.n645 B.n26 10.6151
R778 B.n641 B.n26 10.6151
R779 B.n641 B.n640 10.6151
R780 B.n640 B.n639 10.6151
R781 B.n639 B.n28 10.6151
R782 B.n635 B.n28 10.6151
R783 B.n635 B.n634 10.6151
R784 B.n634 B.n633 10.6151
R785 B.n633 B.n30 10.6151
R786 B.n629 B.n30 10.6151
R787 B.n629 B.n628 10.6151
R788 B.n628 B.n627 10.6151
R789 B.n627 B.n32 10.6151
R790 B.n623 B.n32 10.6151
R791 B.n623 B.n622 10.6151
R792 B.n622 B.n621 10.6151
R793 B.n621 B.n34 10.6151
R794 B.n617 B.n34 10.6151
R795 B.n617 B.n616 10.6151
R796 B.n616 B.n615 10.6151
R797 B.n615 B.n36 10.6151
R798 B.n611 B.n36 10.6151
R799 B.n611 B.n610 10.6151
R800 B.n610 B.n609 10.6151
R801 B.n609 B.n38 10.6151
R802 B.n605 B.n38 10.6151
R803 B.n605 B.n604 10.6151
R804 B.n604 B.n603 10.6151
R805 B.n603 B.n40 10.6151
R806 B.n599 B.n40 10.6151
R807 B.n599 B.n598 10.6151
R808 B.n598 B.n597 10.6151
R809 B.n597 B.n42 10.6151
R810 B.n593 B.n42 10.6151
R811 B.n593 B.n592 10.6151
R812 B.n590 B.n46 10.6151
R813 B.n586 B.n46 10.6151
R814 B.n586 B.n585 10.6151
R815 B.n585 B.n584 10.6151
R816 B.n584 B.n48 10.6151
R817 B.n580 B.n48 10.6151
R818 B.n580 B.n579 10.6151
R819 B.n579 B.n578 10.6151
R820 B.n575 B.n574 10.6151
R821 B.n574 B.n573 10.6151
R822 B.n573 B.n54 10.6151
R823 B.n569 B.n54 10.6151
R824 B.n569 B.n568 10.6151
R825 B.n568 B.n567 10.6151
R826 B.n567 B.n56 10.6151
R827 B.n563 B.n56 10.6151
R828 B.n563 B.n562 10.6151
R829 B.n562 B.n561 10.6151
R830 B.n561 B.n58 10.6151
R831 B.n557 B.n58 10.6151
R832 B.n557 B.n556 10.6151
R833 B.n556 B.n555 10.6151
R834 B.n555 B.n60 10.6151
R835 B.n551 B.n60 10.6151
R836 B.n551 B.n550 10.6151
R837 B.n550 B.n549 10.6151
R838 B.n549 B.n62 10.6151
R839 B.n545 B.n62 10.6151
R840 B.n545 B.n544 10.6151
R841 B.n544 B.n543 10.6151
R842 B.n543 B.n64 10.6151
R843 B.n539 B.n64 10.6151
R844 B.n539 B.n538 10.6151
R845 B.n538 B.n537 10.6151
R846 B.n537 B.n66 10.6151
R847 B.n533 B.n66 10.6151
R848 B.n533 B.n532 10.6151
R849 B.n532 B.n531 10.6151
R850 B.n531 B.n68 10.6151
R851 B.n527 B.n68 10.6151
R852 B.n527 B.n526 10.6151
R853 B.n526 B.n525 10.6151
R854 B.n525 B.n70 10.6151
R855 B.n521 B.n70 10.6151
R856 B.n521 B.n520 10.6151
R857 B.n520 B.n519 10.6151
R858 B.n519 B.n72 10.6151
R859 B.n515 B.n72 10.6151
R860 B.n515 B.n514 10.6151
R861 B.n514 B.n513 10.6151
R862 B.n513 B.n74 10.6151
R863 B.n509 B.n74 10.6151
R864 B.n509 B.n508 10.6151
R865 B.n508 B.n507 10.6151
R866 B.n507 B.n76 10.6151
R867 B.n503 B.n76 10.6151
R868 B.n503 B.n502 10.6151
R869 B.n502 B.n501 10.6151
R870 B.n501 B.n78 10.6151
R871 B.n497 B.n78 10.6151
R872 B.n497 B.n496 10.6151
R873 B.n496 B.n495 10.6151
R874 B.n495 B.n80 10.6151
R875 B.n491 B.n490 10.6151
R876 B.n490 B.n489 10.6151
R877 B.n489 B.n82 10.6151
R878 B.n485 B.n82 10.6151
R879 B.n485 B.n484 10.6151
R880 B.n484 B.n483 10.6151
R881 B.n483 B.n84 10.6151
R882 B.n479 B.n84 10.6151
R883 B.n479 B.n478 10.6151
R884 B.n478 B.n477 10.6151
R885 B.n477 B.n86 10.6151
R886 B.n473 B.n86 10.6151
R887 B.n473 B.n472 10.6151
R888 B.n472 B.n471 10.6151
R889 B.n471 B.n88 10.6151
R890 B.n467 B.n88 10.6151
R891 B.n467 B.n466 10.6151
R892 B.n466 B.n465 10.6151
R893 B.n465 B.n90 10.6151
R894 B.n461 B.n90 10.6151
R895 B.n461 B.n460 10.6151
R896 B.n460 B.n459 10.6151
R897 B.n459 B.n92 10.6151
R898 B.n455 B.n92 10.6151
R899 B.n455 B.n454 10.6151
R900 B.n454 B.n453 10.6151
R901 B.n453 B.n94 10.6151
R902 B.n449 B.n94 10.6151
R903 B.n449 B.n448 10.6151
R904 B.n448 B.n447 10.6151
R905 B.n447 B.n96 10.6151
R906 B.n443 B.n96 10.6151
R907 B.n443 B.n442 10.6151
R908 B.n442 B.n441 10.6151
R909 B.n441 B.n98 10.6151
R910 B.n437 B.n98 10.6151
R911 B.n437 B.n436 10.6151
R912 B.n436 B.n435 10.6151
R913 B.n435 B.n100 10.6151
R914 B.n431 B.n100 10.6151
R915 B.n431 B.n430 10.6151
R916 B.n430 B.n429 10.6151
R917 B.n429 B.n102 10.6151
R918 B.n425 B.n102 10.6151
R919 B.n425 B.n424 10.6151
R920 B.n424 B.n423 10.6151
R921 B.n423 B.n104 10.6151
R922 B.n419 B.n104 10.6151
R923 B.n419 B.n418 10.6151
R924 B.n418 B.n417 10.6151
R925 B.n417 B.n106 10.6151
R926 B.n413 B.n106 10.6151
R927 B.n413 B.n412 10.6151
R928 B.n412 B.n411 10.6151
R929 B.n411 B.n108 10.6151
R930 B.n185 B.n1 10.6151
R931 B.n186 B.n185 10.6151
R932 B.n187 B.n186 10.6151
R933 B.n187 B.n182 10.6151
R934 B.n191 B.n182 10.6151
R935 B.n192 B.n191 10.6151
R936 B.n193 B.n192 10.6151
R937 B.n193 B.n180 10.6151
R938 B.n197 B.n180 10.6151
R939 B.n198 B.n197 10.6151
R940 B.n199 B.n198 10.6151
R941 B.n199 B.n178 10.6151
R942 B.n203 B.n178 10.6151
R943 B.n204 B.n203 10.6151
R944 B.n205 B.n204 10.6151
R945 B.n205 B.n176 10.6151
R946 B.n209 B.n176 10.6151
R947 B.n210 B.n209 10.6151
R948 B.n211 B.n210 10.6151
R949 B.n211 B.n174 10.6151
R950 B.n215 B.n174 10.6151
R951 B.n216 B.n215 10.6151
R952 B.n217 B.n216 10.6151
R953 B.n217 B.n172 10.6151
R954 B.n221 B.n172 10.6151
R955 B.n222 B.n221 10.6151
R956 B.n223 B.n170 10.6151
R957 B.n227 B.n170 10.6151
R958 B.n228 B.n227 10.6151
R959 B.n229 B.n228 10.6151
R960 B.n229 B.n168 10.6151
R961 B.n233 B.n168 10.6151
R962 B.n234 B.n233 10.6151
R963 B.n235 B.n234 10.6151
R964 B.n235 B.n166 10.6151
R965 B.n239 B.n166 10.6151
R966 B.n240 B.n239 10.6151
R967 B.n241 B.n240 10.6151
R968 B.n241 B.n164 10.6151
R969 B.n245 B.n164 10.6151
R970 B.n246 B.n245 10.6151
R971 B.n247 B.n246 10.6151
R972 B.n247 B.n162 10.6151
R973 B.n251 B.n162 10.6151
R974 B.n252 B.n251 10.6151
R975 B.n253 B.n252 10.6151
R976 B.n253 B.n160 10.6151
R977 B.n257 B.n160 10.6151
R978 B.n258 B.n257 10.6151
R979 B.n259 B.n258 10.6151
R980 B.n259 B.n158 10.6151
R981 B.n263 B.n158 10.6151
R982 B.n264 B.n263 10.6151
R983 B.n265 B.n264 10.6151
R984 B.n265 B.n156 10.6151
R985 B.n269 B.n156 10.6151
R986 B.n270 B.n269 10.6151
R987 B.n271 B.n270 10.6151
R988 B.n271 B.n154 10.6151
R989 B.n275 B.n154 10.6151
R990 B.n276 B.n275 10.6151
R991 B.n277 B.n276 10.6151
R992 B.n277 B.n152 10.6151
R993 B.n281 B.n152 10.6151
R994 B.n282 B.n281 10.6151
R995 B.n283 B.n282 10.6151
R996 B.n283 B.n150 10.6151
R997 B.n287 B.n150 10.6151
R998 B.n288 B.n287 10.6151
R999 B.n289 B.n288 10.6151
R1000 B.n289 B.n148 10.6151
R1001 B.n293 B.n148 10.6151
R1002 B.n294 B.n293 10.6151
R1003 B.n295 B.n294 10.6151
R1004 B.n295 B.n146 10.6151
R1005 B.n299 B.n146 10.6151
R1006 B.n300 B.n299 10.6151
R1007 B.n301 B.n300 10.6151
R1008 B.n301 B.n144 10.6151
R1009 B.n305 B.n144 10.6151
R1010 B.n306 B.n305 10.6151
R1011 B.n308 B.n140 10.6151
R1012 B.n312 B.n140 10.6151
R1013 B.n313 B.n312 10.6151
R1014 B.n314 B.n313 10.6151
R1015 B.n314 B.n138 10.6151
R1016 B.n318 B.n138 10.6151
R1017 B.n319 B.n318 10.6151
R1018 B.n323 B.n319 10.6151
R1019 B.n327 B.n136 10.6151
R1020 B.n328 B.n327 10.6151
R1021 B.n329 B.n328 10.6151
R1022 B.n329 B.n134 10.6151
R1023 B.n333 B.n134 10.6151
R1024 B.n334 B.n333 10.6151
R1025 B.n335 B.n334 10.6151
R1026 B.n335 B.n132 10.6151
R1027 B.n339 B.n132 10.6151
R1028 B.n340 B.n339 10.6151
R1029 B.n341 B.n340 10.6151
R1030 B.n341 B.n130 10.6151
R1031 B.n345 B.n130 10.6151
R1032 B.n346 B.n345 10.6151
R1033 B.n347 B.n346 10.6151
R1034 B.n347 B.n128 10.6151
R1035 B.n351 B.n128 10.6151
R1036 B.n352 B.n351 10.6151
R1037 B.n353 B.n352 10.6151
R1038 B.n353 B.n126 10.6151
R1039 B.n357 B.n126 10.6151
R1040 B.n358 B.n357 10.6151
R1041 B.n359 B.n358 10.6151
R1042 B.n359 B.n124 10.6151
R1043 B.n363 B.n124 10.6151
R1044 B.n364 B.n363 10.6151
R1045 B.n365 B.n364 10.6151
R1046 B.n365 B.n122 10.6151
R1047 B.n369 B.n122 10.6151
R1048 B.n370 B.n369 10.6151
R1049 B.n371 B.n370 10.6151
R1050 B.n371 B.n120 10.6151
R1051 B.n375 B.n120 10.6151
R1052 B.n376 B.n375 10.6151
R1053 B.n377 B.n376 10.6151
R1054 B.n377 B.n118 10.6151
R1055 B.n381 B.n118 10.6151
R1056 B.n382 B.n381 10.6151
R1057 B.n383 B.n382 10.6151
R1058 B.n383 B.n116 10.6151
R1059 B.n387 B.n116 10.6151
R1060 B.n388 B.n387 10.6151
R1061 B.n389 B.n388 10.6151
R1062 B.n389 B.n114 10.6151
R1063 B.n393 B.n114 10.6151
R1064 B.n394 B.n393 10.6151
R1065 B.n395 B.n394 10.6151
R1066 B.n395 B.n112 10.6151
R1067 B.n399 B.n112 10.6151
R1068 B.n400 B.n399 10.6151
R1069 B.n401 B.n400 10.6151
R1070 B.n401 B.n110 10.6151
R1071 B.n405 B.n110 10.6151
R1072 B.n406 B.n405 10.6151
R1073 B.n407 B.n406 10.6151
R1074 B.n717 B.n0 8.11757
R1075 B.n717 B.n1 8.11757
R1076 B.n591 B.n590 6.5566
R1077 B.n578 B.n52 6.5566
R1078 B.n308 B.n307 6.5566
R1079 B.n323 B.n322 6.5566
R1080 B.n592 B.n591 4.05904
R1081 B.n575 B.n52 4.05904
R1082 B.n307 B.n306 4.05904
R1083 B.n322 B.n136 4.05904
R1084 VN.n0 VN.t2 248.671
R1085 VN.n1 VN.t3 248.671
R1086 VN.n0 VN.t0 248.154
R1087 VN.n1 VN.t1 248.154
R1088 VN VN.n1 55.647
R1089 VN VN.n0 7.64316
R1090 VTAIL.n746 VTAIL.n658 756.745
R1091 VTAIL.n88 VTAIL.n0 756.745
R1092 VTAIL.n182 VTAIL.n94 756.745
R1093 VTAIL.n276 VTAIL.n188 756.745
R1094 VTAIL.n652 VTAIL.n564 756.745
R1095 VTAIL.n558 VTAIL.n470 756.745
R1096 VTAIL.n464 VTAIL.n376 756.745
R1097 VTAIL.n370 VTAIL.n282 756.745
R1098 VTAIL.n689 VTAIL.n688 585
R1099 VTAIL.n686 VTAIL.n685 585
R1100 VTAIL.n695 VTAIL.n694 585
R1101 VTAIL.n697 VTAIL.n696 585
R1102 VTAIL.n682 VTAIL.n681 585
R1103 VTAIL.n703 VTAIL.n702 585
R1104 VTAIL.n705 VTAIL.n704 585
R1105 VTAIL.n678 VTAIL.n677 585
R1106 VTAIL.n711 VTAIL.n710 585
R1107 VTAIL.n713 VTAIL.n712 585
R1108 VTAIL.n674 VTAIL.n673 585
R1109 VTAIL.n719 VTAIL.n718 585
R1110 VTAIL.n721 VTAIL.n720 585
R1111 VTAIL.n670 VTAIL.n669 585
R1112 VTAIL.n727 VTAIL.n726 585
R1113 VTAIL.n730 VTAIL.n729 585
R1114 VTAIL.n728 VTAIL.n666 585
R1115 VTAIL.n735 VTAIL.n665 585
R1116 VTAIL.n737 VTAIL.n736 585
R1117 VTAIL.n739 VTAIL.n738 585
R1118 VTAIL.n662 VTAIL.n661 585
R1119 VTAIL.n745 VTAIL.n744 585
R1120 VTAIL.n747 VTAIL.n746 585
R1121 VTAIL.n31 VTAIL.n30 585
R1122 VTAIL.n28 VTAIL.n27 585
R1123 VTAIL.n37 VTAIL.n36 585
R1124 VTAIL.n39 VTAIL.n38 585
R1125 VTAIL.n24 VTAIL.n23 585
R1126 VTAIL.n45 VTAIL.n44 585
R1127 VTAIL.n47 VTAIL.n46 585
R1128 VTAIL.n20 VTAIL.n19 585
R1129 VTAIL.n53 VTAIL.n52 585
R1130 VTAIL.n55 VTAIL.n54 585
R1131 VTAIL.n16 VTAIL.n15 585
R1132 VTAIL.n61 VTAIL.n60 585
R1133 VTAIL.n63 VTAIL.n62 585
R1134 VTAIL.n12 VTAIL.n11 585
R1135 VTAIL.n69 VTAIL.n68 585
R1136 VTAIL.n72 VTAIL.n71 585
R1137 VTAIL.n70 VTAIL.n8 585
R1138 VTAIL.n77 VTAIL.n7 585
R1139 VTAIL.n79 VTAIL.n78 585
R1140 VTAIL.n81 VTAIL.n80 585
R1141 VTAIL.n4 VTAIL.n3 585
R1142 VTAIL.n87 VTAIL.n86 585
R1143 VTAIL.n89 VTAIL.n88 585
R1144 VTAIL.n125 VTAIL.n124 585
R1145 VTAIL.n122 VTAIL.n121 585
R1146 VTAIL.n131 VTAIL.n130 585
R1147 VTAIL.n133 VTAIL.n132 585
R1148 VTAIL.n118 VTAIL.n117 585
R1149 VTAIL.n139 VTAIL.n138 585
R1150 VTAIL.n141 VTAIL.n140 585
R1151 VTAIL.n114 VTAIL.n113 585
R1152 VTAIL.n147 VTAIL.n146 585
R1153 VTAIL.n149 VTAIL.n148 585
R1154 VTAIL.n110 VTAIL.n109 585
R1155 VTAIL.n155 VTAIL.n154 585
R1156 VTAIL.n157 VTAIL.n156 585
R1157 VTAIL.n106 VTAIL.n105 585
R1158 VTAIL.n163 VTAIL.n162 585
R1159 VTAIL.n166 VTAIL.n165 585
R1160 VTAIL.n164 VTAIL.n102 585
R1161 VTAIL.n171 VTAIL.n101 585
R1162 VTAIL.n173 VTAIL.n172 585
R1163 VTAIL.n175 VTAIL.n174 585
R1164 VTAIL.n98 VTAIL.n97 585
R1165 VTAIL.n181 VTAIL.n180 585
R1166 VTAIL.n183 VTAIL.n182 585
R1167 VTAIL.n219 VTAIL.n218 585
R1168 VTAIL.n216 VTAIL.n215 585
R1169 VTAIL.n225 VTAIL.n224 585
R1170 VTAIL.n227 VTAIL.n226 585
R1171 VTAIL.n212 VTAIL.n211 585
R1172 VTAIL.n233 VTAIL.n232 585
R1173 VTAIL.n235 VTAIL.n234 585
R1174 VTAIL.n208 VTAIL.n207 585
R1175 VTAIL.n241 VTAIL.n240 585
R1176 VTAIL.n243 VTAIL.n242 585
R1177 VTAIL.n204 VTAIL.n203 585
R1178 VTAIL.n249 VTAIL.n248 585
R1179 VTAIL.n251 VTAIL.n250 585
R1180 VTAIL.n200 VTAIL.n199 585
R1181 VTAIL.n257 VTAIL.n256 585
R1182 VTAIL.n260 VTAIL.n259 585
R1183 VTAIL.n258 VTAIL.n196 585
R1184 VTAIL.n265 VTAIL.n195 585
R1185 VTAIL.n267 VTAIL.n266 585
R1186 VTAIL.n269 VTAIL.n268 585
R1187 VTAIL.n192 VTAIL.n191 585
R1188 VTAIL.n275 VTAIL.n274 585
R1189 VTAIL.n277 VTAIL.n276 585
R1190 VTAIL.n653 VTAIL.n652 585
R1191 VTAIL.n651 VTAIL.n650 585
R1192 VTAIL.n568 VTAIL.n567 585
R1193 VTAIL.n645 VTAIL.n644 585
R1194 VTAIL.n643 VTAIL.n642 585
R1195 VTAIL.n641 VTAIL.n571 585
R1196 VTAIL.n575 VTAIL.n572 585
R1197 VTAIL.n636 VTAIL.n635 585
R1198 VTAIL.n634 VTAIL.n633 585
R1199 VTAIL.n577 VTAIL.n576 585
R1200 VTAIL.n628 VTAIL.n627 585
R1201 VTAIL.n626 VTAIL.n625 585
R1202 VTAIL.n581 VTAIL.n580 585
R1203 VTAIL.n620 VTAIL.n619 585
R1204 VTAIL.n618 VTAIL.n617 585
R1205 VTAIL.n585 VTAIL.n584 585
R1206 VTAIL.n612 VTAIL.n611 585
R1207 VTAIL.n610 VTAIL.n609 585
R1208 VTAIL.n589 VTAIL.n588 585
R1209 VTAIL.n604 VTAIL.n603 585
R1210 VTAIL.n602 VTAIL.n601 585
R1211 VTAIL.n593 VTAIL.n592 585
R1212 VTAIL.n596 VTAIL.n595 585
R1213 VTAIL.n559 VTAIL.n558 585
R1214 VTAIL.n557 VTAIL.n556 585
R1215 VTAIL.n474 VTAIL.n473 585
R1216 VTAIL.n551 VTAIL.n550 585
R1217 VTAIL.n549 VTAIL.n548 585
R1218 VTAIL.n547 VTAIL.n477 585
R1219 VTAIL.n481 VTAIL.n478 585
R1220 VTAIL.n542 VTAIL.n541 585
R1221 VTAIL.n540 VTAIL.n539 585
R1222 VTAIL.n483 VTAIL.n482 585
R1223 VTAIL.n534 VTAIL.n533 585
R1224 VTAIL.n532 VTAIL.n531 585
R1225 VTAIL.n487 VTAIL.n486 585
R1226 VTAIL.n526 VTAIL.n525 585
R1227 VTAIL.n524 VTAIL.n523 585
R1228 VTAIL.n491 VTAIL.n490 585
R1229 VTAIL.n518 VTAIL.n517 585
R1230 VTAIL.n516 VTAIL.n515 585
R1231 VTAIL.n495 VTAIL.n494 585
R1232 VTAIL.n510 VTAIL.n509 585
R1233 VTAIL.n508 VTAIL.n507 585
R1234 VTAIL.n499 VTAIL.n498 585
R1235 VTAIL.n502 VTAIL.n501 585
R1236 VTAIL.n465 VTAIL.n464 585
R1237 VTAIL.n463 VTAIL.n462 585
R1238 VTAIL.n380 VTAIL.n379 585
R1239 VTAIL.n457 VTAIL.n456 585
R1240 VTAIL.n455 VTAIL.n454 585
R1241 VTAIL.n453 VTAIL.n383 585
R1242 VTAIL.n387 VTAIL.n384 585
R1243 VTAIL.n448 VTAIL.n447 585
R1244 VTAIL.n446 VTAIL.n445 585
R1245 VTAIL.n389 VTAIL.n388 585
R1246 VTAIL.n440 VTAIL.n439 585
R1247 VTAIL.n438 VTAIL.n437 585
R1248 VTAIL.n393 VTAIL.n392 585
R1249 VTAIL.n432 VTAIL.n431 585
R1250 VTAIL.n430 VTAIL.n429 585
R1251 VTAIL.n397 VTAIL.n396 585
R1252 VTAIL.n424 VTAIL.n423 585
R1253 VTAIL.n422 VTAIL.n421 585
R1254 VTAIL.n401 VTAIL.n400 585
R1255 VTAIL.n416 VTAIL.n415 585
R1256 VTAIL.n414 VTAIL.n413 585
R1257 VTAIL.n405 VTAIL.n404 585
R1258 VTAIL.n408 VTAIL.n407 585
R1259 VTAIL.n371 VTAIL.n370 585
R1260 VTAIL.n369 VTAIL.n368 585
R1261 VTAIL.n286 VTAIL.n285 585
R1262 VTAIL.n363 VTAIL.n362 585
R1263 VTAIL.n361 VTAIL.n360 585
R1264 VTAIL.n359 VTAIL.n289 585
R1265 VTAIL.n293 VTAIL.n290 585
R1266 VTAIL.n354 VTAIL.n353 585
R1267 VTAIL.n352 VTAIL.n351 585
R1268 VTAIL.n295 VTAIL.n294 585
R1269 VTAIL.n346 VTAIL.n345 585
R1270 VTAIL.n344 VTAIL.n343 585
R1271 VTAIL.n299 VTAIL.n298 585
R1272 VTAIL.n338 VTAIL.n337 585
R1273 VTAIL.n336 VTAIL.n335 585
R1274 VTAIL.n303 VTAIL.n302 585
R1275 VTAIL.n330 VTAIL.n329 585
R1276 VTAIL.n328 VTAIL.n327 585
R1277 VTAIL.n307 VTAIL.n306 585
R1278 VTAIL.n322 VTAIL.n321 585
R1279 VTAIL.n320 VTAIL.n319 585
R1280 VTAIL.n311 VTAIL.n310 585
R1281 VTAIL.n314 VTAIL.n313 585
R1282 VTAIL.t1 VTAIL.n594 327.466
R1283 VTAIL.t2 VTAIL.n500 327.466
R1284 VTAIL.t4 VTAIL.n406 327.466
R1285 VTAIL.t6 VTAIL.n312 327.466
R1286 VTAIL.t7 VTAIL.n687 327.466
R1287 VTAIL.t5 VTAIL.n29 327.466
R1288 VTAIL.t0 VTAIL.n123 327.466
R1289 VTAIL.t3 VTAIL.n217 327.466
R1290 VTAIL.n688 VTAIL.n685 171.744
R1291 VTAIL.n695 VTAIL.n685 171.744
R1292 VTAIL.n696 VTAIL.n695 171.744
R1293 VTAIL.n696 VTAIL.n681 171.744
R1294 VTAIL.n703 VTAIL.n681 171.744
R1295 VTAIL.n704 VTAIL.n703 171.744
R1296 VTAIL.n704 VTAIL.n677 171.744
R1297 VTAIL.n711 VTAIL.n677 171.744
R1298 VTAIL.n712 VTAIL.n711 171.744
R1299 VTAIL.n712 VTAIL.n673 171.744
R1300 VTAIL.n719 VTAIL.n673 171.744
R1301 VTAIL.n720 VTAIL.n719 171.744
R1302 VTAIL.n720 VTAIL.n669 171.744
R1303 VTAIL.n727 VTAIL.n669 171.744
R1304 VTAIL.n729 VTAIL.n727 171.744
R1305 VTAIL.n729 VTAIL.n728 171.744
R1306 VTAIL.n728 VTAIL.n665 171.744
R1307 VTAIL.n737 VTAIL.n665 171.744
R1308 VTAIL.n738 VTAIL.n737 171.744
R1309 VTAIL.n738 VTAIL.n661 171.744
R1310 VTAIL.n745 VTAIL.n661 171.744
R1311 VTAIL.n746 VTAIL.n745 171.744
R1312 VTAIL.n30 VTAIL.n27 171.744
R1313 VTAIL.n37 VTAIL.n27 171.744
R1314 VTAIL.n38 VTAIL.n37 171.744
R1315 VTAIL.n38 VTAIL.n23 171.744
R1316 VTAIL.n45 VTAIL.n23 171.744
R1317 VTAIL.n46 VTAIL.n45 171.744
R1318 VTAIL.n46 VTAIL.n19 171.744
R1319 VTAIL.n53 VTAIL.n19 171.744
R1320 VTAIL.n54 VTAIL.n53 171.744
R1321 VTAIL.n54 VTAIL.n15 171.744
R1322 VTAIL.n61 VTAIL.n15 171.744
R1323 VTAIL.n62 VTAIL.n61 171.744
R1324 VTAIL.n62 VTAIL.n11 171.744
R1325 VTAIL.n69 VTAIL.n11 171.744
R1326 VTAIL.n71 VTAIL.n69 171.744
R1327 VTAIL.n71 VTAIL.n70 171.744
R1328 VTAIL.n70 VTAIL.n7 171.744
R1329 VTAIL.n79 VTAIL.n7 171.744
R1330 VTAIL.n80 VTAIL.n79 171.744
R1331 VTAIL.n80 VTAIL.n3 171.744
R1332 VTAIL.n87 VTAIL.n3 171.744
R1333 VTAIL.n88 VTAIL.n87 171.744
R1334 VTAIL.n124 VTAIL.n121 171.744
R1335 VTAIL.n131 VTAIL.n121 171.744
R1336 VTAIL.n132 VTAIL.n131 171.744
R1337 VTAIL.n132 VTAIL.n117 171.744
R1338 VTAIL.n139 VTAIL.n117 171.744
R1339 VTAIL.n140 VTAIL.n139 171.744
R1340 VTAIL.n140 VTAIL.n113 171.744
R1341 VTAIL.n147 VTAIL.n113 171.744
R1342 VTAIL.n148 VTAIL.n147 171.744
R1343 VTAIL.n148 VTAIL.n109 171.744
R1344 VTAIL.n155 VTAIL.n109 171.744
R1345 VTAIL.n156 VTAIL.n155 171.744
R1346 VTAIL.n156 VTAIL.n105 171.744
R1347 VTAIL.n163 VTAIL.n105 171.744
R1348 VTAIL.n165 VTAIL.n163 171.744
R1349 VTAIL.n165 VTAIL.n164 171.744
R1350 VTAIL.n164 VTAIL.n101 171.744
R1351 VTAIL.n173 VTAIL.n101 171.744
R1352 VTAIL.n174 VTAIL.n173 171.744
R1353 VTAIL.n174 VTAIL.n97 171.744
R1354 VTAIL.n181 VTAIL.n97 171.744
R1355 VTAIL.n182 VTAIL.n181 171.744
R1356 VTAIL.n218 VTAIL.n215 171.744
R1357 VTAIL.n225 VTAIL.n215 171.744
R1358 VTAIL.n226 VTAIL.n225 171.744
R1359 VTAIL.n226 VTAIL.n211 171.744
R1360 VTAIL.n233 VTAIL.n211 171.744
R1361 VTAIL.n234 VTAIL.n233 171.744
R1362 VTAIL.n234 VTAIL.n207 171.744
R1363 VTAIL.n241 VTAIL.n207 171.744
R1364 VTAIL.n242 VTAIL.n241 171.744
R1365 VTAIL.n242 VTAIL.n203 171.744
R1366 VTAIL.n249 VTAIL.n203 171.744
R1367 VTAIL.n250 VTAIL.n249 171.744
R1368 VTAIL.n250 VTAIL.n199 171.744
R1369 VTAIL.n257 VTAIL.n199 171.744
R1370 VTAIL.n259 VTAIL.n257 171.744
R1371 VTAIL.n259 VTAIL.n258 171.744
R1372 VTAIL.n258 VTAIL.n195 171.744
R1373 VTAIL.n267 VTAIL.n195 171.744
R1374 VTAIL.n268 VTAIL.n267 171.744
R1375 VTAIL.n268 VTAIL.n191 171.744
R1376 VTAIL.n275 VTAIL.n191 171.744
R1377 VTAIL.n276 VTAIL.n275 171.744
R1378 VTAIL.n652 VTAIL.n651 171.744
R1379 VTAIL.n651 VTAIL.n567 171.744
R1380 VTAIL.n644 VTAIL.n567 171.744
R1381 VTAIL.n644 VTAIL.n643 171.744
R1382 VTAIL.n643 VTAIL.n571 171.744
R1383 VTAIL.n575 VTAIL.n571 171.744
R1384 VTAIL.n635 VTAIL.n575 171.744
R1385 VTAIL.n635 VTAIL.n634 171.744
R1386 VTAIL.n634 VTAIL.n576 171.744
R1387 VTAIL.n627 VTAIL.n576 171.744
R1388 VTAIL.n627 VTAIL.n626 171.744
R1389 VTAIL.n626 VTAIL.n580 171.744
R1390 VTAIL.n619 VTAIL.n580 171.744
R1391 VTAIL.n619 VTAIL.n618 171.744
R1392 VTAIL.n618 VTAIL.n584 171.744
R1393 VTAIL.n611 VTAIL.n584 171.744
R1394 VTAIL.n611 VTAIL.n610 171.744
R1395 VTAIL.n610 VTAIL.n588 171.744
R1396 VTAIL.n603 VTAIL.n588 171.744
R1397 VTAIL.n603 VTAIL.n602 171.744
R1398 VTAIL.n602 VTAIL.n592 171.744
R1399 VTAIL.n595 VTAIL.n592 171.744
R1400 VTAIL.n558 VTAIL.n557 171.744
R1401 VTAIL.n557 VTAIL.n473 171.744
R1402 VTAIL.n550 VTAIL.n473 171.744
R1403 VTAIL.n550 VTAIL.n549 171.744
R1404 VTAIL.n549 VTAIL.n477 171.744
R1405 VTAIL.n481 VTAIL.n477 171.744
R1406 VTAIL.n541 VTAIL.n481 171.744
R1407 VTAIL.n541 VTAIL.n540 171.744
R1408 VTAIL.n540 VTAIL.n482 171.744
R1409 VTAIL.n533 VTAIL.n482 171.744
R1410 VTAIL.n533 VTAIL.n532 171.744
R1411 VTAIL.n532 VTAIL.n486 171.744
R1412 VTAIL.n525 VTAIL.n486 171.744
R1413 VTAIL.n525 VTAIL.n524 171.744
R1414 VTAIL.n524 VTAIL.n490 171.744
R1415 VTAIL.n517 VTAIL.n490 171.744
R1416 VTAIL.n517 VTAIL.n516 171.744
R1417 VTAIL.n516 VTAIL.n494 171.744
R1418 VTAIL.n509 VTAIL.n494 171.744
R1419 VTAIL.n509 VTAIL.n508 171.744
R1420 VTAIL.n508 VTAIL.n498 171.744
R1421 VTAIL.n501 VTAIL.n498 171.744
R1422 VTAIL.n464 VTAIL.n463 171.744
R1423 VTAIL.n463 VTAIL.n379 171.744
R1424 VTAIL.n456 VTAIL.n379 171.744
R1425 VTAIL.n456 VTAIL.n455 171.744
R1426 VTAIL.n455 VTAIL.n383 171.744
R1427 VTAIL.n387 VTAIL.n383 171.744
R1428 VTAIL.n447 VTAIL.n387 171.744
R1429 VTAIL.n447 VTAIL.n446 171.744
R1430 VTAIL.n446 VTAIL.n388 171.744
R1431 VTAIL.n439 VTAIL.n388 171.744
R1432 VTAIL.n439 VTAIL.n438 171.744
R1433 VTAIL.n438 VTAIL.n392 171.744
R1434 VTAIL.n431 VTAIL.n392 171.744
R1435 VTAIL.n431 VTAIL.n430 171.744
R1436 VTAIL.n430 VTAIL.n396 171.744
R1437 VTAIL.n423 VTAIL.n396 171.744
R1438 VTAIL.n423 VTAIL.n422 171.744
R1439 VTAIL.n422 VTAIL.n400 171.744
R1440 VTAIL.n415 VTAIL.n400 171.744
R1441 VTAIL.n415 VTAIL.n414 171.744
R1442 VTAIL.n414 VTAIL.n404 171.744
R1443 VTAIL.n407 VTAIL.n404 171.744
R1444 VTAIL.n370 VTAIL.n369 171.744
R1445 VTAIL.n369 VTAIL.n285 171.744
R1446 VTAIL.n362 VTAIL.n285 171.744
R1447 VTAIL.n362 VTAIL.n361 171.744
R1448 VTAIL.n361 VTAIL.n289 171.744
R1449 VTAIL.n293 VTAIL.n289 171.744
R1450 VTAIL.n353 VTAIL.n293 171.744
R1451 VTAIL.n353 VTAIL.n352 171.744
R1452 VTAIL.n352 VTAIL.n294 171.744
R1453 VTAIL.n345 VTAIL.n294 171.744
R1454 VTAIL.n345 VTAIL.n344 171.744
R1455 VTAIL.n344 VTAIL.n298 171.744
R1456 VTAIL.n337 VTAIL.n298 171.744
R1457 VTAIL.n337 VTAIL.n336 171.744
R1458 VTAIL.n336 VTAIL.n302 171.744
R1459 VTAIL.n329 VTAIL.n302 171.744
R1460 VTAIL.n329 VTAIL.n328 171.744
R1461 VTAIL.n328 VTAIL.n306 171.744
R1462 VTAIL.n321 VTAIL.n306 171.744
R1463 VTAIL.n321 VTAIL.n320 171.744
R1464 VTAIL.n320 VTAIL.n310 171.744
R1465 VTAIL.n313 VTAIL.n310 171.744
R1466 VTAIL.n688 VTAIL.t7 85.8723
R1467 VTAIL.n30 VTAIL.t5 85.8723
R1468 VTAIL.n124 VTAIL.t0 85.8723
R1469 VTAIL.n218 VTAIL.t3 85.8723
R1470 VTAIL.n595 VTAIL.t1 85.8723
R1471 VTAIL.n501 VTAIL.t2 85.8723
R1472 VTAIL.n407 VTAIL.t4 85.8723
R1473 VTAIL.n313 VTAIL.t6 85.8723
R1474 VTAIL.n751 VTAIL.n750 32.9611
R1475 VTAIL.n93 VTAIL.n92 32.9611
R1476 VTAIL.n187 VTAIL.n186 32.9611
R1477 VTAIL.n281 VTAIL.n280 32.9611
R1478 VTAIL.n657 VTAIL.n656 32.9611
R1479 VTAIL.n563 VTAIL.n562 32.9611
R1480 VTAIL.n469 VTAIL.n468 32.9611
R1481 VTAIL.n375 VTAIL.n374 32.9611
R1482 VTAIL.n751 VTAIL.n657 28.8065
R1483 VTAIL.n375 VTAIL.n281 28.8065
R1484 VTAIL.n689 VTAIL.n687 16.3895
R1485 VTAIL.n31 VTAIL.n29 16.3895
R1486 VTAIL.n125 VTAIL.n123 16.3895
R1487 VTAIL.n219 VTAIL.n217 16.3895
R1488 VTAIL.n596 VTAIL.n594 16.3895
R1489 VTAIL.n502 VTAIL.n500 16.3895
R1490 VTAIL.n408 VTAIL.n406 16.3895
R1491 VTAIL.n314 VTAIL.n312 16.3895
R1492 VTAIL.n736 VTAIL.n735 13.1884
R1493 VTAIL.n78 VTAIL.n77 13.1884
R1494 VTAIL.n172 VTAIL.n171 13.1884
R1495 VTAIL.n266 VTAIL.n265 13.1884
R1496 VTAIL.n642 VTAIL.n641 13.1884
R1497 VTAIL.n548 VTAIL.n547 13.1884
R1498 VTAIL.n454 VTAIL.n453 13.1884
R1499 VTAIL.n360 VTAIL.n359 13.1884
R1500 VTAIL.n690 VTAIL.n686 12.8005
R1501 VTAIL.n734 VTAIL.n666 12.8005
R1502 VTAIL.n739 VTAIL.n664 12.8005
R1503 VTAIL.n32 VTAIL.n28 12.8005
R1504 VTAIL.n76 VTAIL.n8 12.8005
R1505 VTAIL.n81 VTAIL.n6 12.8005
R1506 VTAIL.n126 VTAIL.n122 12.8005
R1507 VTAIL.n170 VTAIL.n102 12.8005
R1508 VTAIL.n175 VTAIL.n100 12.8005
R1509 VTAIL.n220 VTAIL.n216 12.8005
R1510 VTAIL.n264 VTAIL.n196 12.8005
R1511 VTAIL.n269 VTAIL.n194 12.8005
R1512 VTAIL.n645 VTAIL.n570 12.8005
R1513 VTAIL.n640 VTAIL.n572 12.8005
R1514 VTAIL.n597 VTAIL.n593 12.8005
R1515 VTAIL.n551 VTAIL.n476 12.8005
R1516 VTAIL.n546 VTAIL.n478 12.8005
R1517 VTAIL.n503 VTAIL.n499 12.8005
R1518 VTAIL.n457 VTAIL.n382 12.8005
R1519 VTAIL.n452 VTAIL.n384 12.8005
R1520 VTAIL.n409 VTAIL.n405 12.8005
R1521 VTAIL.n363 VTAIL.n288 12.8005
R1522 VTAIL.n358 VTAIL.n290 12.8005
R1523 VTAIL.n315 VTAIL.n311 12.8005
R1524 VTAIL.n694 VTAIL.n693 12.0247
R1525 VTAIL.n731 VTAIL.n730 12.0247
R1526 VTAIL.n740 VTAIL.n662 12.0247
R1527 VTAIL.n36 VTAIL.n35 12.0247
R1528 VTAIL.n73 VTAIL.n72 12.0247
R1529 VTAIL.n82 VTAIL.n4 12.0247
R1530 VTAIL.n130 VTAIL.n129 12.0247
R1531 VTAIL.n167 VTAIL.n166 12.0247
R1532 VTAIL.n176 VTAIL.n98 12.0247
R1533 VTAIL.n224 VTAIL.n223 12.0247
R1534 VTAIL.n261 VTAIL.n260 12.0247
R1535 VTAIL.n270 VTAIL.n192 12.0247
R1536 VTAIL.n646 VTAIL.n568 12.0247
R1537 VTAIL.n637 VTAIL.n636 12.0247
R1538 VTAIL.n601 VTAIL.n600 12.0247
R1539 VTAIL.n552 VTAIL.n474 12.0247
R1540 VTAIL.n543 VTAIL.n542 12.0247
R1541 VTAIL.n507 VTAIL.n506 12.0247
R1542 VTAIL.n458 VTAIL.n380 12.0247
R1543 VTAIL.n449 VTAIL.n448 12.0247
R1544 VTAIL.n413 VTAIL.n412 12.0247
R1545 VTAIL.n364 VTAIL.n286 12.0247
R1546 VTAIL.n355 VTAIL.n354 12.0247
R1547 VTAIL.n319 VTAIL.n318 12.0247
R1548 VTAIL.n697 VTAIL.n684 11.249
R1549 VTAIL.n726 VTAIL.n668 11.249
R1550 VTAIL.n744 VTAIL.n743 11.249
R1551 VTAIL.n39 VTAIL.n26 11.249
R1552 VTAIL.n68 VTAIL.n10 11.249
R1553 VTAIL.n86 VTAIL.n85 11.249
R1554 VTAIL.n133 VTAIL.n120 11.249
R1555 VTAIL.n162 VTAIL.n104 11.249
R1556 VTAIL.n180 VTAIL.n179 11.249
R1557 VTAIL.n227 VTAIL.n214 11.249
R1558 VTAIL.n256 VTAIL.n198 11.249
R1559 VTAIL.n274 VTAIL.n273 11.249
R1560 VTAIL.n650 VTAIL.n649 11.249
R1561 VTAIL.n633 VTAIL.n574 11.249
R1562 VTAIL.n604 VTAIL.n591 11.249
R1563 VTAIL.n556 VTAIL.n555 11.249
R1564 VTAIL.n539 VTAIL.n480 11.249
R1565 VTAIL.n510 VTAIL.n497 11.249
R1566 VTAIL.n462 VTAIL.n461 11.249
R1567 VTAIL.n445 VTAIL.n386 11.249
R1568 VTAIL.n416 VTAIL.n403 11.249
R1569 VTAIL.n368 VTAIL.n367 11.249
R1570 VTAIL.n351 VTAIL.n292 11.249
R1571 VTAIL.n322 VTAIL.n309 11.249
R1572 VTAIL.n698 VTAIL.n682 10.4732
R1573 VTAIL.n725 VTAIL.n670 10.4732
R1574 VTAIL.n747 VTAIL.n660 10.4732
R1575 VTAIL.n40 VTAIL.n24 10.4732
R1576 VTAIL.n67 VTAIL.n12 10.4732
R1577 VTAIL.n89 VTAIL.n2 10.4732
R1578 VTAIL.n134 VTAIL.n118 10.4732
R1579 VTAIL.n161 VTAIL.n106 10.4732
R1580 VTAIL.n183 VTAIL.n96 10.4732
R1581 VTAIL.n228 VTAIL.n212 10.4732
R1582 VTAIL.n255 VTAIL.n200 10.4732
R1583 VTAIL.n277 VTAIL.n190 10.4732
R1584 VTAIL.n653 VTAIL.n566 10.4732
R1585 VTAIL.n632 VTAIL.n577 10.4732
R1586 VTAIL.n605 VTAIL.n589 10.4732
R1587 VTAIL.n559 VTAIL.n472 10.4732
R1588 VTAIL.n538 VTAIL.n483 10.4732
R1589 VTAIL.n511 VTAIL.n495 10.4732
R1590 VTAIL.n465 VTAIL.n378 10.4732
R1591 VTAIL.n444 VTAIL.n389 10.4732
R1592 VTAIL.n417 VTAIL.n401 10.4732
R1593 VTAIL.n371 VTAIL.n284 10.4732
R1594 VTAIL.n350 VTAIL.n295 10.4732
R1595 VTAIL.n323 VTAIL.n307 10.4732
R1596 VTAIL.n702 VTAIL.n701 9.69747
R1597 VTAIL.n722 VTAIL.n721 9.69747
R1598 VTAIL.n748 VTAIL.n658 9.69747
R1599 VTAIL.n44 VTAIL.n43 9.69747
R1600 VTAIL.n64 VTAIL.n63 9.69747
R1601 VTAIL.n90 VTAIL.n0 9.69747
R1602 VTAIL.n138 VTAIL.n137 9.69747
R1603 VTAIL.n158 VTAIL.n157 9.69747
R1604 VTAIL.n184 VTAIL.n94 9.69747
R1605 VTAIL.n232 VTAIL.n231 9.69747
R1606 VTAIL.n252 VTAIL.n251 9.69747
R1607 VTAIL.n278 VTAIL.n188 9.69747
R1608 VTAIL.n654 VTAIL.n564 9.69747
R1609 VTAIL.n629 VTAIL.n628 9.69747
R1610 VTAIL.n609 VTAIL.n608 9.69747
R1611 VTAIL.n560 VTAIL.n470 9.69747
R1612 VTAIL.n535 VTAIL.n534 9.69747
R1613 VTAIL.n515 VTAIL.n514 9.69747
R1614 VTAIL.n466 VTAIL.n376 9.69747
R1615 VTAIL.n441 VTAIL.n440 9.69747
R1616 VTAIL.n421 VTAIL.n420 9.69747
R1617 VTAIL.n372 VTAIL.n282 9.69747
R1618 VTAIL.n347 VTAIL.n346 9.69747
R1619 VTAIL.n327 VTAIL.n326 9.69747
R1620 VTAIL.n750 VTAIL.n749 9.45567
R1621 VTAIL.n92 VTAIL.n91 9.45567
R1622 VTAIL.n186 VTAIL.n185 9.45567
R1623 VTAIL.n280 VTAIL.n279 9.45567
R1624 VTAIL.n656 VTAIL.n655 9.45567
R1625 VTAIL.n562 VTAIL.n561 9.45567
R1626 VTAIL.n468 VTAIL.n467 9.45567
R1627 VTAIL.n374 VTAIL.n373 9.45567
R1628 VTAIL.n749 VTAIL.n748 9.3005
R1629 VTAIL.n660 VTAIL.n659 9.3005
R1630 VTAIL.n743 VTAIL.n742 9.3005
R1631 VTAIL.n741 VTAIL.n740 9.3005
R1632 VTAIL.n664 VTAIL.n663 9.3005
R1633 VTAIL.n709 VTAIL.n708 9.3005
R1634 VTAIL.n707 VTAIL.n706 9.3005
R1635 VTAIL.n680 VTAIL.n679 9.3005
R1636 VTAIL.n701 VTAIL.n700 9.3005
R1637 VTAIL.n699 VTAIL.n698 9.3005
R1638 VTAIL.n684 VTAIL.n683 9.3005
R1639 VTAIL.n693 VTAIL.n692 9.3005
R1640 VTAIL.n691 VTAIL.n690 9.3005
R1641 VTAIL.n676 VTAIL.n675 9.3005
R1642 VTAIL.n715 VTAIL.n714 9.3005
R1643 VTAIL.n717 VTAIL.n716 9.3005
R1644 VTAIL.n672 VTAIL.n671 9.3005
R1645 VTAIL.n723 VTAIL.n722 9.3005
R1646 VTAIL.n725 VTAIL.n724 9.3005
R1647 VTAIL.n668 VTAIL.n667 9.3005
R1648 VTAIL.n732 VTAIL.n731 9.3005
R1649 VTAIL.n734 VTAIL.n733 9.3005
R1650 VTAIL.n91 VTAIL.n90 9.3005
R1651 VTAIL.n2 VTAIL.n1 9.3005
R1652 VTAIL.n85 VTAIL.n84 9.3005
R1653 VTAIL.n83 VTAIL.n82 9.3005
R1654 VTAIL.n6 VTAIL.n5 9.3005
R1655 VTAIL.n51 VTAIL.n50 9.3005
R1656 VTAIL.n49 VTAIL.n48 9.3005
R1657 VTAIL.n22 VTAIL.n21 9.3005
R1658 VTAIL.n43 VTAIL.n42 9.3005
R1659 VTAIL.n41 VTAIL.n40 9.3005
R1660 VTAIL.n26 VTAIL.n25 9.3005
R1661 VTAIL.n35 VTAIL.n34 9.3005
R1662 VTAIL.n33 VTAIL.n32 9.3005
R1663 VTAIL.n18 VTAIL.n17 9.3005
R1664 VTAIL.n57 VTAIL.n56 9.3005
R1665 VTAIL.n59 VTAIL.n58 9.3005
R1666 VTAIL.n14 VTAIL.n13 9.3005
R1667 VTAIL.n65 VTAIL.n64 9.3005
R1668 VTAIL.n67 VTAIL.n66 9.3005
R1669 VTAIL.n10 VTAIL.n9 9.3005
R1670 VTAIL.n74 VTAIL.n73 9.3005
R1671 VTAIL.n76 VTAIL.n75 9.3005
R1672 VTAIL.n185 VTAIL.n184 9.3005
R1673 VTAIL.n96 VTAIL.n95 9.3005
R1674 VTAIL.n179 VTAIL.n178 9.3005
R1675 VTAIL.n177 VTAIL.n176 9.3005
R1676 VTAIL.n100 VTAIL.n99 9.3005
R1677 VTAIL.n145 VTAIL.n144 9.3005
R1678 VTAIL.n143 VTAIL.n142 9.3005
R1679 VTAIL.n116 VTAIL.n115 9.3005
R1680 VTAIL.n137 VTAIL.n136 9.3005
R1681 VTAIL.n135 VTAIL.n134 9.3005
R1682 VTAIL.n120 VTAIL.n119 9.3005
R1683 VTAIL.n129 VTAIL.n128 9.3005
R1684 VTAIL.n127 VTAIL.n126 9.3005
R1685 VTAIL.n112 VTAIL.n111 9.3005
R1686 VTAIL.n151 VTAIL.n150 9.3005
R1687 VTAIL.n153 VTAIL.n152 9.3005
R1688 VTAIL.n108 VTAIL.n107 9.3005
R1689 VTAIL.n159 VTAIL.n158 9.3005
R1690 VTAIL.n161 VTAIL.n160 9.3005
R1691 VTAIL.n104 VTAIL.n103 9.3005
R1692 VTAIL.n168 VTAIL.n167 9.3005
R1693 VTAIL.n170 VTAIL.n169 9.3005
R1694 VTAIL.n279 VTAIL.n278 9.3005
R1695 VTAIL.n190 VTAIL.n189 9.3005
R1696 VTAIL.n273 VTAIL.n272 9.3005
R1697 VTAIL.n271 VTAIL.n270 9.3005
R1698 VTAIL.n194 VTAIL.n193 9.3005
R1699 VTAIL.n239 VTAIL.n238 9.3005
R1700 VTAIL.n237 VTAIL.n236 9.3005
R1701 VTAIL.n210 VTAIL.n209 9.3005
R1702 VTAIL.n231 VTAIL.n230 9.3005
R1703 VTAIL.n229 VTAIL.n228 9.3005
R1704 VTAIL.n214 VTAIL.n213 9.3005
R1705 VTAIL.n223 VTAIL.n222 9.3005
R1706 VTAIL.n221 VTAIL.n220 9.3005
R1707 VTAIL.n206 VTAIL.n205 9.3005
R1708 VTAIL.n245 VTAIL.n244 9.3005
R1709 VTAIL.n247 VTAIL.n246 9.3005
R1710 VTAIL.n202 VTAIL.n201 9.3005
R1711 VTAIL.n253 VTAIL.n252 9.3005
R1712 VTAIL.n255 VTAIL.n254 9.3005
R1713 VTAIL.n198 VTAIL.n197 9.3005
R1714 VTAIL.n262 VTAIL.n261 9.3005
R1715 VTAIL.n264 VTAIL.n263 9.3005
R1716 VTAIL.n622 VTAIL.n621 9.3005
R1717 VTAIL.n624 VTAIL.n623 9.3005
R1718 VTAIL.n579 VTAIL.n578 9.3005
R1719 VTAIL.n630 VTAIL.n629 9.3005
R1720 VTAIL.n632 VTAIL.n631 9.3005
R1721 VTAIL.n574 VTAIL.n573 9.3005
R1722 VTAIL.n638 VTAIL.n637 9.3005
R1723 VTAIL.n640 VTAIL.n639 9.3005
R1724 VTAIL.n655 VTAIL.n654 9.3005
R1725 VTAIL.n566 VTAIL.n565 9.3005
R1726 VTAIL.n649 VTAIL.n648 9.3005
R1727 VTAIL.n647 VTAIL.n646 9.3005
R1728 VTAIL.n570 VTAIL.n569 9.3005
R1729 VTAIL.n583 VTAIL.n582 9.3005
R1730 VTAIL.n616 VTAIL.n615 9.3005
R1731 VTAIL.n614 VTAIL.n613 9.3005
R1732 VTAIL.n587 VTAIL.n586 9.3005
R1733 VTAIL.n608 VTAIL.n607 9.3005
R1734 VTAIL.n606 VTAIL.n605 9.3005
R1735 VTAIL.n591 VTAIL.n590 9.3005
R1736 VTAIL.n600 VTAIL.n599 9.3005
R1737 VTAIL.n598 VTAIL.n597 9.3005
R1738 VTAIL.n528 VTAIL.n527 9.3005
R1739 VTAIL.n530 VTAIL.n529 9.3005
R1740 VTAIL.n485 VTAIL.n484 9.3005
R1741 VTAIL.n536 VTAIL.n535 9.3005
R1742 VTAIL.n538 VTAIL.n537 9.3005
R1743 VTAIL.n480 VTAIL.n479 9.3005
R1744 VTAIL.n544 VTAIL.n543 9.3005
R1745 VTAIL.n546 VTAIL.n545 9.3005
R1746 VTAIL.n561 VTAIL.n560 9.3005
R1747 VTAIL.n472 VTAIL.n471 9.3005
R1748 VTAIL.n555 VTAIL.n554 9.3005
R1749 VTAIL.n553 VTAIL.n552 9.3005
R1750 VTAIL.n476 VTAIL.n475 9.3005
R1751 VTAIL.n489 VTAIL.n488 9.3005
R1752 VTAIL.n522 VTAIL.n521 9.3005
R1753 VTAIL.n520 VTAIL.n519 9.3005
R1754 VTAIL.n493 VTAIL.n492 9.3005
R1755 VTAIL.n514 VTAIL.n513 9.3005
R1756 VTAIL.n512 VTAIL.n511 9.3005
R1757 VTAIL.n497 VTAIL.n496 9.3005
R1758 VTAIL.n506 VTAIL.n505 9.3005
R1759 VTAIL.n504 VTAIL.n503 9.3005
R1760 VTAIL.n434 VTAIL.n433 9.3005
R1761 VTAIL.n436 VTAIL.n435 9.3005
R1762 VTAIL.n391 VTAIL.n390 9.3005
R1763 VTAIL.n442 VTAIL.n441 9.3005
R1764 VTAIL.n444 VTAIL.n443 9.3005
R1765 VTAIL.n386 VTAIL.n385 9.3005
R1766 VTAIL.n450 VTAIL.n449 9.3005
R1767 VTAIL.n452 VTAIL.n451 9.3005
R1768 VTAIL.n467 VTAIL.n466 9.3005
R1769 VTAIL.n378 VTAIL.n377 9.3005
R1770 VTAIL.n461 VTAIL.n460 9.3005
R1771 VTAIL.n459 VTAIL.n458 9.3005
R1772 VTAIL.n382 VTAIL.n381 9.3005
R1773 VTAIL.n395 VTAIL.n394 9.3005
R1774 VTAIL.n428 VTAIL.n427 9.3005
R1775 VTAIL.n426 VTAIL.n425 9.3005
R1776 VTAIL.n399 VTAIL.n398 9.3005
R1777 VTAIL.n420 VTAIL.n419 9.3005
R1778 VTAIL.n418 VTAIL.n417 9.3005
R1779 VTAIL.n403 VTAIL.n402 9.3005
R1780 VTAIL.n412 VTAIL.n411 9.3005
R1781 VTAIL.n410 VTAIL.n409 9.3005
R1782 VTAIL.n340 VTAIL.n339 9.3005
R1783 VTAIL.n342 VTAIL.n341 9.3005
R1784 VTAIL.n297 VTAIL.n296 9.3005
R1785 VTAIL.n348 VTAIL.n347 9.3005
R1786 VTAIL.n350 VTAIL.n349 9.3005
R1787 VTAIL.n292 VTAIL.n291 9.3005
R1788 VTAIL.n356 VTAIL.n355 9.3005
R1789 VTAIL.n358 VTAIL.n357 9.3005
R1790 VTAIL.n373 VTAIL.n372 9.3005
R1791 VTAIL.n284 VTAIL.n283 9.3005
R1792 VTAIL.n367 VTAIL.n366 9.3005
R1793 VTAIL.n365 VTAIL.n364 9.3005
R1794 VTAIL.n288 VTAIL.n287 9.3005
R1795 VTAIL.n301 VTAIL.n300 9.3005
R1796 VTAIL.n334 VTAIL.n333 9.3005
R1797 VTAIL.n332 VTAIL.n331 9.3005
R1798 VTAIL.n305 VTAIL.n304 9.3005
R1799 VTAIL.n326 VTAIL.n325 9.3005
R1800 VTAIL.n324 VTAIL.n323 9.3005
R1801 VTAIL.n309 VTAIL.n308 9.3005
R1802 VTAIL.n318 VTAIL.n317 9.3005
R1803 VTAIL.n316 VTAIL.n315 9.3005
R1804 VTAIL.n705 VTAIL.n680 8.92171
R1805 VTAIL.n718 VTAIL.n672 8.92171
R1806 VTAIL.n47 VTAIL.n22 8.92171
R1807 VTAIL.n60 VTAIL.n14 8.92171
R1808 VTAIL.n141 VTAIL.n116 8.92171
R1809 VTAIL.n154 VTAIL.n108 8.92171
R1810 VTAIL.n235 VTAIL.n210 8.92171
R1811 VTAIL.n248 VTAIL.n202 8.92171
R1812 VTAIL.n625 VTAIL.n579 8.92171
R1813 VTAIL.n612 VTAIL.n587 8.92171
R1814 VTAIL.n531 VTAIL.n485 8.92171
R1815 VTAIL.n518 VTAIL.n493 8.92171
R1816 VTAIL.n437 VTAIL.n391 8.92171
R1817 VTAIL.n424 VTAIL.n399 8.92171
R1818 VTAIL.n343 VTAIL.n297 8.92171
R1819 VTAIL.n330 VTAIL.n305 8.92171
R1820 VTAIL.n706 VTAIL.n678 8.14595
R1821 VTAIL.n717 VTAIL.n674 8.14595
R1822 VTAIL.n48 VTAIL.n20 8.14595
R1823 VTAIL.n59 VTAIL.n16 8.14595
R1824 VTAIL.n142 VTAIL.n114 8.14595
R1825 VTAIL.n153 VTAIL.n110 8.14595
R1826 VTAIL.n236 VTAIL.n208 8.14595
R1827 VTAIL.n247 VTAIL.n204 8.14595
R1828 VTAIL.n624 VTAIL.n581 8.14595
R1829 VTAIL.n613 VTAIL.n585 8.14595
R1830 VTAIL.n530 VTAIL.n487 8.14595
R1831 VTAIL.n519 VTAIL.n491 8.14595
R1832 VTAIL.n436 VTAIL.n393 8.14595
R1833 VTAIL.n425 VTAIL.n397 8.14595
R1834 VTAIL.n342 VTAIL.n299 8.14595
R1835 VTAIL.n331 VTAIL.n303 8.14595
R1836 VTAIL.n710 VTAIL.n709 7.3702
R1837 VTAIL.n714 VTAIL.n713 7.3702
R1838 VTAIL.n52 VTAIL.n51 7.3702
R1839 VTAIL.n56 VTAIL.n55 7.3702
R1840 VTAIL.n146 VTAIL.n145 7.3702
R1841 VTAIL.n150 VTAIL.n149 7.3702
R1842 VTAIL.n240 VTAIL.n239 7.3702
R1843 VTAIL.n244 VTAIL.n243 7.3702
R1844 VTAIL.n621 VTAIL.n620 7.3702
R1845 VTAIL.n617 VTAIL.n616 7.3702
R1846 VTAIL.n527 VTAIL.n526 7.3702
R1847 VTAIL.n523 VTAIL.n522 7.3702
R1848 VTAIL.n433 VTAIL.n432 7.3702
R1849 VTAIL.n429 VTAIL.n428 7.3702
R1850 VTAIL.n339 VTAIL.n338 7.3702
R1851 VTAIL.n335 VTAIL.n334 7.3702
R1852 VTAIL.n710 VTAIL.n676 6.59444
R1853 VTAIL.n713 VTAIL.n676 6.59444
R1854 VTAIL.n52 VTAIL.n18 6.59444
R1855 VTAIL.n55 VTAIL.n18 6.59444
R1856 VTAIL.n146 VTAIL.n112 6.59444
R1857 VTAIL.n149 VTAIL.n112 6.59444
R1858 VTAIL.n240 VTAIL.n206 6.59444
R1859 VTAIL.n243 VTAIL.n206 6.59444
R1860 VTAIL.n620 VTAIL.n583 6.59444
R1861 VTAIL.n617 VTAIL.n583 6.59444
R1862 VTAIL.n526 VTAIL.n489 6.59444
R1863 VTAIL.n523 VTAIL.n489 6.59444
R1864 VTAIL.n432 VTAIL.n395 6.59444
R1865 VTAIL.n429 VTAIL.n395 6.59444
R1866 VTAIL.n338 VTAIL.n301 6.59444
R1867 VTAIL.n335 VTAIL.n301 6.59444
R1868 VTAIL.n709 VTAIL.n678 5.81868
R1869 VTAIL.n714 VTAIL.n674 5.81868
R1870 VTAIL.n51 VTAIL.n20 5.81868
R1871 VTAIL.n56 VTAIL.n16 5.81868
R1872 VTAIL.n145 VTAIL.n114 5.81868
R1873 VTAIL.n150 VTAIL.n110 5.81868
R1874 VTAIL.n239 VTAIL.n208 5.81868
R1875 VTAIL.n244 VTAIL.n204 5.81868
R1876 VTAIL.n621 VTAIL.n581 5.81868
R1877 VTAIL.n616 VTAIL.n585 5.81868
R1878 VTAIL.n527 VTAIL.n487 5.81868
R1879 VTAIL.n522 VTAIL.n491 5.81868
R1880 VTAIL.n433 VTAIL.n393 5.81868
R1881 VTAIL.n428 VTAIL.n397 5.81868
R1882 VTAIL.n339 VTAIL.n299 5.81868
R1883 VTAIL.n334 VTAIL.n303 5.81868
R1884 VTAIL.n706 VTAIL.n705 5.04292
R1885 VTAIL.n718 VTAIL.n717 5.04292
R1886 VTAIL.n48 VTAIL.n47 5.04292
R1887 VTAIL.n60 VTAIL.n59 5.04292
R1888 VTAIL.n142 VTAIL.n141 5.04292
R1889 VTAIL.n154 VTAIL.n153 5.04292
R1890 VTAIL.n236 VTAIL.n235 5.04292
R1891 VTAIL.n248 VTAIL.n247 5.04292
R1892 VTAIL.n625 VTAIL.n624 5.04292
R1893 VTAIL.n613 VTAIL.n612 5.04292
R1894 VTAIL.n531 VTAIL.n530 5.04292
R1895 VTAIL.n519 VTAIL.n518 5.04292
R1896 VTAIL.n437 VTAIL.n436 5.04292
R1897 VTAIL.n425 VTAIL.n424 5.04292
R1898 VTAIL.n343 VTAIL.n342 5.04292
R1899 VTAIL.n331 VTAIL.n330 5.04292
R1900 VTAIL.n702 VTAIL.n680 4.26717
R1901 VTAIL.n721 VTAIL.n672 4.26717
R1902 VTAIL.n750 VTAIL.n658 4.26717
R1903 VTAIL.n44 VTAIL.n22 4.26717
R1904 VTAIL.n63 VTAIL.n14 4.26717
R1905 VTAIL.n92 VTAIL.n0 4.26717
R1906 VTAIL.n138 VTAIL.n116 4.26717
R1907 VTAIL.n157 VTAIL.n108 4.26717
R1908 VTAIL.n186 VTAIL.n94 4.26717
R1909 VTAIL.n232 VTAIL.n210 4.26717
R1910 VTAIL.n251 VTAIL.n202 4.26717
R1911 VTAIL.n280 VTAIL.n188 4.26717
R1912 VTAIL.n656 VTAIL.n564 4.26717
R1913 VTAIL.n628 VTAIL.n579 4.26717
R1914 VTAIL.n609 VTAIL.n587 4.26717
R1915 VTAIL.n562 VTAIL.n470 4.26717
R1916 VTAIL.n534 VTAIL.n485 4.26717
R1917 VTAIL.n515 VTAIL.n493 4.26717
R1918 VTAIL.n468 VTAIL.n376 4.26717
R1919 VTAIL.n440 VTAIL.n391 4.26717
R1920 VTAIL.n421 VTAIL.n399 4.26717
R1921 VTAIL.n374 VTAIL.n282 4.26717
R1922 VTAIL.n346 VTAIL.n297 4.26717
R1923 VTAIL.n327 VTAIL.n305 4.26717
R1924 VTAIL.n691 VTAIL.n687 3.70982
R1925 VTAIL.n33 VTAIL.n29 3.70982
R1926 VTAIL.n127 VTAIL.n123 3.70982
R1927 VTAIL.n221 VTAIL.n217 3.70982
R1928 VTAIL.n598 VTAIL.n594 3.70982
R1929 VTAIL.n504 VTAIL.n500 3.70982
R1930 VTAIL.n410 VTAIL.n406 3.70982
R1931 VTAIL.n316 VTAIL.n312 3.70982
R1932 VTAIL.n701 VTAIL.n682 3.49141
R1933 VTAIL.n722 VTAIL.n670 3.49141
R1934 VTAIL.n748 VTAIL.n747 3.49141
R1935 VTAIL.n43 VTAIL.n24 3.49141
R1936 VTAIL.n64 VTAIL.n12 3.49141
R1937 VTAIL.n90 VTAIL.n89 3.49141
R1938 VTAIL.n137 VTAIL.n118 3.49141
R1939 VTAIL.n158 VTAIL.n106 3.49141
R1940 VTAIL.n184 VTAIL.n183 3.49141
R1941 VTAIL.n231 VTAIL.n212 3.49141
R1942 VTAIL.n252 VTAIL.n200 3.49141
R1943 VTAIL.n278 VTAIL.n277 3.49141
R1944 VTAIL.n654 VTAIL.n653 3.49141
R1945 VTAIL.n629 VTAIL.n577 3.49141
R1946 VTAIL.n608 VTAIL.n589 3.49141
R1947 VTAIL.n560 VTAIL.n559 3.49141
R1948 VTAIL.n535 VTAIL.n483 3.49141
R1949 VTAIL.n514 VTAIL.n495 3.49141
R1950 VTAIL.n466 VTAIL.n465 3.49141
R1951 VTAIL.n441 VTAIL.n389 3.49141
R1952 VTAIL.n420 VTAIL.n401 3.49141
R1953 VTAIL.n372 VTAIL.n371 3.49141
R1954 VTAIL.n347 VTAIL.n295 3.49141
R1955 VTAIL.n326 VTAIL.n307 3.49141
R1956 VTAIL.n698 VTAIL.n697 2.71565
R1957 VTAIL.n726 VTAIL.n725 2.71565
R1958 VTAIL.n744 VTAIL.n660 2.71565
R1959 VTAIL.n40 VTAIL.n39 2.71565
R1960 VTAIL.n68 VTAIL.n67 2.71565
R1961 VTAIL.n86 VTAIL.n2 2.71565
R1962 VTAIL.n134 VTAIL.n133 2.71565
R1963 VTAIL.n162 VTAIL.n161 2.71565
R1964 VTAIL.n180 VTAIL.n96 2.71565
R1965 VTAIL.n228 VTAIL.n227 2.71565
R1966 VTAIL.n256 VTAIL.n255 2.71565
R1967 VTAIL.n274 VTAIL.n190 2.71565
R1968 VTAIL.n650 VTAIL.n566 2.71565
R1969 VTAIL.n633 VTAIL.n632 2.71565
R1970 VTAIL.n605 VTAIL.n604 2.71565
R1971 VTAIL.n556 VTAIL.n472 2.71565
R1972 VTAIL.n539 VTAIL.n538 2.71565
R1973 VTAIL.n511 VTAIL.n510 2.71565
R1974 VTAIL.n462 VTAIL.n378 2.71565
R1975 VTAIL.n445 VTAIL.n444 2.71565
R1976 VTAIL.n417 VTAIL.n416 2.71565
R1977 VTAIL.n368 VTAIL.n284 2.71565
R1978 VTAIL.n351 VTAIL.n350 2.71565
R1979 VTAIL.n323 VTAIL.n322 2.71565
R1980 VTAIL.n694 VTAIL.n684 1.93989
R1981 VTAIL.n730 VTAIL.n668 1.93989
R1982 VTAIL.n743 VTAIL.n662 1.93989
R1983 VTAIL.n36 VTAIL.n26 1.93989
R1984 VTAIL.n72 VTAIL.n10 1.93989
R1985 VTAIL.n85 VTAIL.n4 1.93989
R1986 VTAIL.n130 VTAIL.n120 1.93989
R1987 VTAIL.n166 VTAIL.n104 1.93989
R1988 VTAIL.n179 VTAIL.n98 1.93989
R1989 VTAIL.n224 VTAIL.n214 1.93989
R1990 VTAIL.n260 VTAIL.n198 1.93989
R1991 VTAIL.n273 VTAIL.n192 1.93989
R1992 VTAIL.n649 VTAIL.n568 1.93989
R1993 VTAIL.n636 VTAIL.n574 1.93989
R1994 VTAIL.n601 VTAIL.n591 1.93989
R1995 VTAIL.n555 VTAIL.n474 1.93989
R1996 VTAIL.n542 VTAIL.n480 1.93989
R1997 VTAIL.n507 VTAIL.n497 1.93989
R1998 VTAIL.n461 VTAIL.n380 1.93989
R1999 VTAIL.n448 VTAIL.n386 1.93989
R2000 VTAIL.n413 VTAIL.n403 1.93989
R2001 VTAIL.n367 VTAIL.n286 1.93989
R2002 VTAIL.n354 VTAIL.n292 1.93989
R2003 VTAIL.n319 VTAIL.n309 1.93989
R2004 VTAIL.n469 VTAIL.n375 1.92291
R2005 VTAIL.n657 VTAIL.n563 1.92291
R2006 VTAIL.n281 VTAIL.n187 1.92291
R2007 VTAIL.n693 VTAIL.n686 1.16414
R2008 VTAIL.n731 VTAIL.n666 1.16414
R2009 VTAIL.n740 VTAIL.n739 1.16414
R2010 VTAIL.n35 VTAIL.n28 1.16414
R2011 VTAIL.n73 VTAIL.n8 1.16414
R2012 VTAIL.n82 VTAIL.n81 1.16414
R2013 VTAIL.n129 VTAIL.n122 1.16414
R2014 VTAIL.n167 VTAIL.n102 1.16414
R2015 VTAIL.n176 VTAIL.n175 1.16414
R2016 VTAIL.n223 VTAIL.n216 1.16414
R2017 VTAIL.n261 VTAIL.n196 1.16414
R2018 VTAIL.n270 VTAIL.n269 1.16414
R2019 VTAIL.n646 VTAIL.n645 1.16414
R2020 VTAIL.n637 VTAIL.n572 1.16414
R2021 VTAIL.n600 VTAIL.n593 1.16414
R2022 VTAIL.n552 VTAIL.n551 1.16414
R2023 VTAIL.n543 VTAIL.n478 1.16414
R2024 VTAIL.n506 VTAIL.n499 1.16414
R2025 VTAIL.n458 VTAIL.n457 1.16414
R2026 VTAIL.n449 VTAIL.n384 1.16414
R2027 VTAIL.n412 VTAIL.n405 1.16414
R2028 VTAIL.n364 VTAIL.n363 1.16414
R2029 VTAIL.n355 VTAIL.n290 1.16414
R2030 VTAIL.n318 VTAIL.n311 1.16414
R2031 VTAIL VTAIL.n93 1.0199
R2032 VTAIL VTAIL.n751 0.903517
R2033 VTAIL.n563 VTAIL.n469 0.470328
R2034 VTAIL.n187 VTAIL.n93 0.470328
R2035 VTAIL.n690 VTAIL.n689 0.388379
R2036 VTAIL.n735 VTAIL.n734 0.388379
R2037 VTAIL.n736 VTAIL.n664 0.388379
R2038 VTAIL.n32 VTAIL.n31 0.388379
R2039 VTAIL.n77 VTAIL.n76 0.388379
R2040 VTAIL.n78 VTAIL.n6 0.388379
R2041 VTAIL.n126 VTAIL.n125 0.388379
R2042 VTAIL.n171 VTAIL.n170 0.388379
R2043 VTAIL.n172 VTAIL.n100 0.388379
R2044 VTAIL.n220 VTAIL.n219 0.388379
R2045 VTAIL.n265 VTAIL.n264 0.388379
R2046 VTAIL.n266 VTAIL.n194 0.388379
R2047 VTAIL.n642 VTAIL.n570 0.388379
R2048 VTAIL.n641 VTAIL.n640 0.388379
R2049 VTAIL.n597 VTAIL.n596 0.388379
R2050 VTAIL.n548 VTAIL.n476 0.388379
R2051 VTAIL.n547 VTAIL.n546 0.388379
R2052 VTAIL.n503 VTAIL.n502 0.388379
R2053 VTAIL.n454 VTAIL.n382 0.388379
R2054 VTAIL.n453 VTAIL.n452 0.388379
R2055 VTAIL.n409 VTAIL.n408 0.388379
R2056 VTAIL.n360 VTAIL.n288 0.388379
R2057 VTAIL.n359 VTAIL.n358 0.388379
R2058 VTAIL.n315 VTAIL.n314 0.388379
R2059 VTAIL.n692 VTAIL.n691 0.155672
R2060 VTAIL.n692 VTAIL.n683 0.155672
R2061 VTAIL.n699 VTAIL.n683 0.155672
R2062 VTAIL.n700 VTAIL.n699 0.155672
R2063 VTAIL.n700 VTAIL.n679 0.155672
R2064 VTAIL.n707 VTAIL.n679 0.155672
R2065 VTAIL.n708 VTAIL.n707 0.155672
R2066 VTAIL.n708 VTAIL.n675 0.155672
R2067 VTAIL.n715 VTAIL.n675 0.155672
R2068 VTAIL.n716 VTAIL.n715 0.155672
R2069 VTAIL.n716 VTAIL.n671 0.155672
R2070 VTAIL.n723 VTAIL.n671 0.155672
R2071 VTAIL.n724 VTAIL.n723 0.155672
R2072 VTAIL.n724 VTAIL.n667 0.155672
R2073 VTAIL.n732 VTAIL.n667 0.155672
R2074 VTAIL.n733 VTAIL.n732 0.155672
R2075 VTAIL.n733 VTAIL.n663 0.155672
R2076 VTAIL.n741 VTAIL.n663 0.155672
R2077 VTAIL.n742 VTAIL.n741 0.155672
R2078 VTAIL.n742 VTAIL.n659 0.155672
R2079 VTAIL.n749 VTAIL.n659 0.155672
R2080 VTAIL.n34 VTAIL.n33 0.155672
R2081 VTAIL.n34 VTAIL.n25 0.155672
R2082 VTAIL.n41 VTAIL.n25 0.155672
R2083 VTAIL.n42 VTAIL.n41 0.155672
R2084 VTAIL.n42 VTAIL.n21 0.155672
R2085 VTAIL.n49 VTAIL.n21 0.155672
R2086 VTAIL.n50 VTAIL.n49 0.155672
R2087 VTAIL.n50 VTAIL.n17 0.155672
R2088 VTAIL.n57 VTAIL.n17 0.155672
R2089 VTAIL.n58 VTAIL.n57 0.155672
R2090 VTAIL.n58 VTAIL.n13 0.155672
R2091 VTAIL.n65 VTAIL.n13 0.155672
R2092 VTAIL.n66 VTAIL.n65 0.155672
R2093 VTAIL.n66 VTAIL.n9 0.155672
R2094 VTAIL.n74 VTAIL.n9 0.155672
R2095 VTAIL.n75 VTAIL.n74 0.155672
R2096 VTAIL.n75 VTAIL.n5 0.155672
R2097 VTAIL.n83 VTAIL.n5 0.155672
R2098 VTAIL.n84 VTAIL.n83 0.155672
R2099 VTAIL.n84 VTAIL.n1 0.155672
R2100 VTAIL.n91 VTAIL.n1 0.155672
R2101 VTAIL.n128 VTAIL.n127 0.155672
R2102 VTAIL.n128 VTAIL.n119 0.155672
R2103 VTAIL.n135 VTAIL.n119 0.155672
R2104 VTAIL.n136 VTAIL.n135 0.155672
R2105 VTAIL.n136 VTAIL.n115 0.155672
R2106 VTAIL.n143 VTAIL.n115 0.155672
R2107 VTAIL.n144 VTAIL.n143 0.155672
R2108 VTAIL.n144 VTAIL.n111 0.155672
R2109 VTAIL.n151 VTAIL.n111 0.155672
R2110 VTAIL.n152 VTAIL.n151 0.155672
R2111 VTAIL.n152 VTAIL.n107 0.155672
R2112 VTAIL.n159 VTAIL.n107 0.155672
R2113 VTAIL.n160 VTAIL.n159 0.155672
R2114 VTAIL.n160 VTAIL.n103 0.155672
R2115 VTAIL.n168 VTAIL.n103 0.155672
R2116 VTAIL.n169 VTAIL.n168 0.155672
R2117 VTAIL.n169 VTAIL.n99 0.155672
R2118 VTAIL.n177 VTAIL.n99 0.155672
R2119 VTAIL.n178 VTAIL.n177 0.155672
R2120 VTAIL.n178 VTAIL.n95 0.155672
R2121 VTAIL.n185 VTAIL.n95 0.155672
R2122 VTAIL.n222 VTAIL.n221 0.155672
R2123 VTAIL.n222 VTAIL.n213 0.155672
R2124 VTAIL.n229 VTAIL.n213 0.155672
R2125 VTAIL.n230 VTAIL.n229 0.155672
R2126 VTAIL.n230 VTAIL.n209 0.155672
R2127 VTAIL.n237 VTAIL.n209 0.155672
R2128 VTAIL.n238 VTAIL.n237 0.155672
R2129 VTAIL.n238 VTAIL.n205 0.155672
R2130 VTAIL.n245 VTAIL.n205 0.155672
R2131 VTAIL.n246 VTAIL.n245 0.155672
R2132 VTAIL.n246 VTAIL.n201 0.155672
R2133 VTAIL.n253 VTAIL.n201 0.155672
R2134 VTAIL.n254 VTAIL.n253 0.155672
R2135 VTAIL.n254 VTAIL.n197 0.155672
R2136 VTAIL.n262 VTAIL.n197 0.155672
R2137 VTAIL.n263 VTAIL.n262 0.155672
R2138 VTAIL.n263 VTAIL.n193 0.155672
R2139 VTAIL.n271 VTAIL.n193 0.155672
R2140 VTAIL.n272 VTAIL.n271 0.155672
R2141 VTAIL.n272 VTAIL.n189 0.155672
R2142 VTAIL.n279 VTAIL.n189 0.155672
R2143 VTAIL.n655 VTAIL.n565 0.155672
R2144 VTAIL.n648 VTAIL.n565 0.155672
R2145 VTAIL.n648 VTAIL.n647 0.155672
R2146 VTAIL.n647 VTAIL.n569 0.155672
R2147 VTAIL.n639 VTAIL.n569 0.155672
R2148 VTAIL.n639 VTAIL.n638 0.155672
R2149 VTAIL.n638 VTAIL.n573 0.155672
R2150 VTAIL.n631 VTAIL.n573 0.155672
R2151 VTAIL.n631 VTAIL.n630 0.155672
R2152 VTAIL.n630 VTAIL.n578 0.155672
R2153 VTAIL.n623 VTAIL.n578 0.155672
R2154 VTAIL.n623 VTAIL.n622 0.155672
R2155 VTAIL.n622 VTAIL.n582 0.155672
R2156 VTAIL.n615 VTAIL.n582 0.155672
R2157 VTAIL.n615 VTAIL.n614 0.155672
R2158 VTAIL.n614 VTAIL.n586 0.155672
R2159 VTAIL.n607 VTAIL.n586 0.155672
R2160 VTAIL.n607 VTAIL.n606 0.155672
R2161 VTAIL.n606 VTAIL.n590 0.155672
R2162 VTAIL.n599 VTAIL.n590 0.155672
R2163 VTAIL.n599 VTAIL.n598 0.155672
R2164 VTAIL.n561 VTAIL.n471 0.155672
R2165 VTAIL.n554 VTAIL.n471 0.155672
R2166 VTAIL.n554 VTAIL.n553 0.155672
R2167 VTAIL.n553 VTAIL.n475 0.155672
R2168 VTAIL.n545 VTAIL.n475 0.155672
R2169 VTAIL.n545 VTAIL.n544 0.155672
R2170 VTAIL.n544 VTAIL.n479 0.155672
R2171 VTAIL.n537 VTAIL.n479 0.155672
R2172 VTAIL.n537 VTAIL.n536 0.155672
R2173 VTAIL.n536 VTAIL.n484 0.155672
R2174 VTAIL.n529 VTAIL.n484 0.155672
R2175 VTAIL.n529 VTAIL.n528 0.155672
R2176 VTAIL.n528 VTAIL.n488 0.155672
R2177 VTAIL.n521 VTAIL.n488 0.155672
R2178 VTAIL.n521 VTAIL.n520 0.155672
R2179 VTAIL.n520 VTAIL.n492 0.155672
R2180 VTAIL.n513 VTAIL.n492 0.155672
R2181 VTAIL.n513 VTAIL.n512 0.155672
R2182 VTAIL.n512 VTAIL.n496 0.155672
R2183 VTAIL.n505 VTAIL.n496 0.155672
R2184 VTAIL.n505 VTAIL.n504 0.155672
R2185 VTAIL.n467 VTAIL.n377 0.155672
R2186 VTAIL.n460 VTAIL.n377 0.155672
R2187 VTAIL.n460 VTAIL.n459 0.155672
R2188 VTAIL.n459 VTAIL.n381 0.155672
R2189 VTAIL.n451 VTAIL.n381 0.155672
R2190 VTAIL.n451 VTAIL.n450 0.155672
R2191 VTAIL.n450 VTAIL.n385 0.155672
R2192 VTAIL.n443 VTAIL.n385 0.155672
R2193 VTAIL.n443 VTAIL.n442 0.155672
R2194 VTAIL.n442 VTAIL.n390 0.155672
R2195 VTAIL.n435 VTAIL.n390 0.155672
R2196 VTAIL.n435 VTAIL.n434 0.155672
R2197 VTAIL.n434 VTAIL.n394 0.155672
R2198 VTAIL.n427 VTAIL.n394 0.155672
R2199 VTAIL.n427 VTAIL.n426 0.155672
R2200 VTAIL.n426 VTAIL.n398 0.155672
R2201 VTAIL.n419 VTAIL.n398 0.155672
R2202 VTAIL.n419 VTAIL.n418 0.155672
R2203 VTAIL.n418 VTAIL.n402 0.155672
R2204 VTAIL.n411 VTAIL.n402 0.155672
R2205 VTAIL.n411 VTAIL.n410 0.155672
R2206 VTAIL.n373 VTAIL.n283 0.155672
R2207 VTAIL.n366 VTAIL.n283 0.155672
R2208 VTAIL.n366 VTAIL.n365 0.155672
R2209 VTAIL.n365 VTAIL.n287 0.155672
R2210 VTAIL.n357 VTAIL.n287 0.155672
R2211 VTAIL.n357 VTAIL.n356 0.155672
R2212 VTAIL.n356 VTAIL.n291 0.155672
R2213 VTAIL.n349 VTAIL.n291 0.155672
R2214 VTAIL.n349 VTAIL.n348 0.155672
R2215 VTAIL.n348 VTAIL.n296 0.155672
R2216 VTAIL.n341 VTAIL.n296 0.155672
R2217 VTAIL.n341 VTAIL.n340 0.155672
R2218 VTAIL.n340 VTAIL.n300 0.155672
R2219 VTAIL.n333 VTAIL.n300 0.155672
R2220 VTAIL.n333 VTAIL.n332 0.155672
R2221 VTAIL.n332 VTAIL.n304 0.155672
R2222 VTAIL.n325 VTAIL.n304 0.155672
R2223 VTAIL.n325 VTAIL.n324 0.155672
R2224 VTAIL.n324 VTAIL.n308 0.155672
R2225 VTAIL.n317 VTAIL.n308 0.155672
R2226 VTAIL.n317 VTAIL.n316 0.155672
R2227 VDD2.n2 VDD2.n0 114.166
R2228 VDD2.n2 VDD2.n1 70.1676
R2229 VDD2.n1 VDD2.t2 1.93073
R2230 VDD2.n1 VDD2.t0 1.93073
R2231 VDD2.n0 VDD2.t1 1.93073
R2232 VDD2.n0 VDD2.t3 1.93073
R2233 VDD2 VDD2.n2 0.0586897
R2234 VP.n2 VP.t1 248.671
R2235 VP.n2 VP.t0 248.154
R2236 VP.n4 VP.t2 213.602
R2237 VP.n11 VP.t3 213.602
R2238 VP.n10 VP.n0 161.3
R2239 VP.n9 VP.n8 161.3
R2240 VP.n7 VP.n1 161.3
R2241 VP.n6 VP.n5 161.3
R2242 VP.n4 VP.n3 92.9562
R2243 VP.n12 VP.n11 92.9562
R2244 VP.n9 VP.n1 56.5617
R2245 VP.n3 VP.n2 55.3681
R2246 VP.n5 VP.n1 24.5923
R2247 VP.n10 VP.n9 24.5923
R2248 VP.n5 VP.n4 17.9525
R2249 VP.n11 VP.n10 17.9525
R2250 VP.n6 VP.n3 0.278335
R2251 VP.n12 VP.n0 0.278335
R2252 VP.n7 VP.n6 0.189894
R2253 VP.n8 VP.n7 0.189894
R2254 VP.n8 VP.n0 0.189894
R2255 VP VP.n12 0.153485
R2256 VDD1 VDD1.n1 114.692
R2257 VDD1 VDD1.n0 70.2258
R2258 VDD1.n0 VDD1.t2 1.93073
R2259 VDD1.n0 VDD1.t3 1.93073
R2260 VDD1.n1 VDD1.t1 1.93073
R2261 VDD1.n1 VDD1.t0 1.93073
C0 VTAIL VDD1 6.70452f
C1 VTAIL B 6.11488f
C2 VTAIL VDD2 6.75403f
C3 VN VDD1 0.148825f
C4 VTAIL VP 5.753779f
C5 VN B 1.03593f
C6 VTAIL w_n2308_n4336# 5.09205f
C7 VN VDD2 6.12103f
C8 VN VP 6.58385f
C9 VN w_n2308_n4336# 3.87606f
C10 VDD1 B 1.26953f
C11 VDD1 VDD2 0.858804f
C12 VDD2 B 1.31022f
C13 VDD1 VP 6.32186f
C14 B VP 1.5221f
C15 VDD1 w_n2308_n4336# 1.4483f
C16 VDD2 VP 0.350221f
C17 w_n2308_n4336# B 9.74149f
C18 VDD2 w_n2308_n4336# 1.48877f
C19 w_n2308_n4336# VP 4.171f
C20 VN VTAIL 5.73967f
C21 VDD2 VSUBS 0.950965f
C22 VDD1 VSUBS 5.96899f
C23 VTAIL VSUBS 1.369509f
C24 VN VSUBS 5.41908f
C25 VP VSUBS 2.101485f
C26 B VSUBS 4.077576f
C27 w_n2308_n4336# VSUBS 0.122499p
C28 VDD1.t2 VSUBS 0.353457f
C29 VDD1.t3 VSUBS 0.353457f
C30 VDD1.n0 VSUBS 2.91559f
C31 VDD1.t1 VSUBS 0.353457f
C32 VDD1.t0 VSUBS 0.353457f
C33 VDD1.n1 VSUBS 3.801f
C34 VP.n0 VSUBS 0.048994f
C35 VP.t3 VSUBS 3.26643f
C36 VP.n1 VSUBS 0.054023f
C37 VP.t0 VSUBS 3.45105f
C38 VP.t1 VSUBS 3.45384f
C39 VP.n2 VSUBS 4.23755f
C40 VP.n3 VSUBS 2.24433f
C41 VP.t2 VSUBS 3.26643f
C42 VP.n4 VSUBS 1.24841f
C43 VP.n5 VSUBS 0.059731f
C44 VP.n6 VSUBS 0.048994f
C45 VP.n7 VSUBS 0.037164f
C46 VP.n8 VSUBS 0.037164f
C47 VP.n9 VSUBS 0.054023f
C48 VP.n10 VSUBS 0.059731f
C49 VP.n11 VSUBS 1.24841f
C50 VP.n12 VSUBS 0.046367f
C51 VDD2.t1 VSUBS 0.353405f
C52 VDD2.t3 VSUBS 0.353405f
C53 VDD2.n0 VSUBS 3.77372f
C54 VDD2.t2 VSUBS 0.353405f
C55 VDD2.t0 VSUBS 0.353405f
C56 VDD2.n1 VSUBS 2.91458f
C57 VDD2.n2 VSUBS 4.62785f
C58 VTAIL.n0 VSUBS 0.023865f
C59 VTAIL.n1 VSUBS 0.022145f
C60 VTAIL.n2 VSUBS 0.0119f
C61 VTAIL.n3 VSUBS 0.028127f
C62 VTAIL.n4 VSUBS 0.0126f
C63 VTAIL.n5 VSUBS 0.022145f
C64 VTAIL.n6 VSUBS 0.0119f
C65 VTAIL.n7 VSUBS 0.028127f
C66 VTAIL.n8 VSUBS 0.0126f
C67 VTAIL.n9 VSUBS 0.022145f
C68 VTAIL.n10 VSUBS 0.0119f
C69 VTAIL.n11 VSUBS 0.028127f
C70 VTAIL.n12 VSUBS 0.0126f
C71 VTAIL.n13 VSUBS 0.022145f
C72 VTAIL.n14 VSUBS 0.0119f
C73 VTAIL.n15 VSUBS 0.028127f
C74 VTAIL.n16 VSUBS 0.0126f
C75 VTAIL.n17 VSUBS 0.022145f
C76 VTAIL.n18 VSUBS 0.0119f
C77 VTAIL.n19 VSUBS 0.028127f
C78 VTAIL.n20 VSUBS 0.0126f
C79 VTAIL.n21 VSUBS 0.022145f
C80 VTAIL.n22 VSUBS 0.0119f
C81 VTAIL.n23 VSUBS 0.028127f
C82 VTAIL.n24 VSUBS 0.0126f
C83 VTAIL.n25 VSUBS 0.022145f
C84 VTAIL.n26 VSUBS 0.0119f
C85 VTAIL.n27 VSUBS 0.028127f
C86 VTAIL.n28 VSUBS 0.0126f
C87 VTAIL.n29 VSUBS 0.168125f
C88 VTAIL.t5 VSUBS 0.060316f
C89 VTAIL.n30 VSUBS 0.021096f
C90 VTAIL.n31 VSUBS 0.017893f
C91 VTAIL.n32 VSUBS 0.0119f
C92 VTAIL.n33 VSUBS 1.59902f
C93 VTAIL.n34 VSUBS 0.022145f
C94 VTAIL.n35 VSUBS 0.0119f
C95 VTAIL.n36 VSUBS 0.0126f
C96 VTAIL.n37 VSUBS 0.028127f
C97 VTAIL.n38 VSUBS 0.028127f
C98 VTAIL.n39 VSUBS 0.0126f
C99 VTAIL.n40 VSUBS 0.0119f
C100 VTAIL.n41 VSUBS 0.022145f
C101 VTAIL.n42 VSUBS 0.022145f
C102 VTAIL.n43 VSUBS 0.0119f
C103 VTAIL.n44 VSUBS 0.0126f
C104 VTAIL.n45 VSUBS 0.028127f
C105 VTAIL.n46 VSUBS 0.028127f
C106 VTAIL.n47 VSUBS 0.0126f
C107 VTAIL.n48 VSUBS 0.0119f
C108 VTAIL.n49 VSUBS 0.022145f
C109 VTAIL.n50 VSUBS 0.022145f
C110 VTAIL.n51 VSUBS 0.0119f
C111 VTAIL.n52 VSUBS 0.0126f
C112 VTAIL.n53 VSUBS 0.028127f
C113 VTAIL.n54 VSUBS 0.028127f
C114 VTAIL.n55 VSUBS 0.0126f
C115 VTAIL.n56 VSUBS 0.0119f
C116 VTAIL.n57 VSUBS 0.022145f
C117 VTAIL.n58 VSUBS 0.022145f
C118 VTAIL.n59 VSUBS 0.0119f
C119 VTAIL.n60 VSUBS 0.0126f
C120 VTAIL.n61 VSUBS 0.028127f
C121 VTAIL.n62 VSUBS 0.028127f
C122 VTAIL.n63 VSUBS 0.0126f
C123 VTAIL.n64 VSUBS 0.0119f
C124 VTAIL.n65 VSUBS 0.022145f
C125 VTAIL.n66 VSUBS 0.022145f
C126 VTAIL.n67 VSUBS 0.0119f
C127 VTAIL.n68 VSUBS 0.0126f
C128 VTAIL.n69 VSUBS 0.028127f
C129 VTAIL.n70 VSUBS 0.028127f
C130 VTAIL.n71 VSUBS 0.028127f
C131 VTAIL.n72 VSUBS 0.0126f
C132 VTAIL.n73 VSUBS 0.0119f
C133 VTAIL.n74 VSUBS 0.022145f
C134 VTAIL.n75 VSUBS 0.022145f
C135 VTAIL.n76 VSUBS 0.0119f
C136 VTAIL.n77 VSUBS 0.01225f
C137 VTAIL.n78 VSUBS 0.01225f
C138 VTAIL.n79 VSUBS 0.028127f
C139 VTAIL.n80 VSUBS 0.028127f
C140 VTAIL.n81 VSUBS 0.0126f
C141 VTAIL.n82 VSUBS 0.0119f
C142 VTAIL.n83 VSUBS 0.022145f
C143 VTAIL.n84 VSUBS 0.022145f
C144 VTAIL.n85 VSUBS 0.0119f
C145 VTAIL.n86 VSUBS 0.0126f
C146 VTAIL.n87 VSUBS 0.028127f
C147 VTAIL.n88 VSUBS 0.066499f
C148 VTAIL.n89 VSUBS 0.0126f
C149 VTAIL.n90 VSUBS 0.0119f
C150 VTAIL.n91 VSUBS 0.052398f
C151 VTAIL.n92 VSUBS 0.033408f
C152 VTAIL.n93 VSUBS 0.125865f
C153 VTAIL.n94 VSUBS 0.023865f
C154 VTAIL.n95 VSUBS 0.022145f
C155 VTAIL.n96 VSUBS 0.0119f
C156 VTAIL.n97 VSUBS 0.028127f
C157 VTAIL.n98 VSUBS 0.0126f
C158 VTAIL.n99 VSUBS 0.022145f
C159 VTAIL.n100 VSUBS 0.0119f
C160 VTAIL.n101 VSUBS 0.028127f
C161 VTAIL.n102 VSUBS 0.0126f
C162 VTAIL.n103 VSUBS 0.022145f
C163 VTAIL.n104 VSUBS 0.0119f
C164 VTAIL.n105 VSUBS 0.028127f
C165 VTAIL.n106 VSUBS 0.0126f
C166 VTAIL.n107 VSUBS 0.022145f
C167 VTAIL.n108 VSUBS 0.0119f
C168 VTAIL.n109 VSUBS 0.028127f
C169 VTAIL.n110 VSUBS 0.0126f
C170 VTAIL.n111 VSUBS 0.022145f
C171 VTAIL.n112 VSUBS 0.0119f
C172 VTAIL.n113 VSUBS 0.028127f
C173 VTAIL.n114 VSUBS 0.0126f
C174 VTAIL.n115 VSUBS 0.022145f
C175 VTAIL.n116 VSUBS 0.0119f
C176 VTAIL.n117 VSUBS 0.028127f
C177 VTAIL.n118 VSUBS 0.0126f
C178 VTAIL.n119 VSUBS 0.022145f
C179 VTAIL.n120 VSUBS 0.0119f
C180 VTAIL.n121 VSUBS 0.028127f
C181 VTAIL.n122 VSUBS 0.0126f
C182 VTAIL.n123 VSUBS 0.168125f
C183 VTAIL.t0 VSUBS 0.060316f
C184 VTAIL.n124 VSUBS 0.021096f
C185 VTAIL.n125 VSUBS 0.017893f
C186 VTAIL.n126 VSUBS 0.0119f
C187 VTAIL.n127 VSUBS 1.59902f
C188 VTAIL.n128 VSUBS 0.022145f
C189 VTAIL.n129 VSUBS 0.0119f
C190 VTAIL.n130 VSUBS 0.0126f
C191 VTAIL.n131 VSUBS 0.028127f
C192 VTAIL.n132 VSUBS 0.028127f
C193 VTAIL.n133 VSUBS 0.0126f
C194 VTAIL.n134 VSUBS 0.0119f
C195 VTAIL.n135 VSUBS 0.022145f
C196 VTAIL.n136 VSUBS 0.022145f
C197 VTAIL.n137 VSUBS 0.0119f
C198 VTAIL.n138 VSUBS 0.0126f
C199 VTAIL.n139 VSUBS 0.028127f
C200 VTAIL.n140 VSUBS 0.028127f
C201 VTAIL.n141 VSUBS 0.0126f
C202 VTAIL.n142 VSUBS 0.0119f
C203 VTAIL.n143 VSUBS 0.022145f
C204 VTAIL.n144 VSUBS 0.022145f
C205 VTAIL.n145 VSUBS 0.0119f
C206 VTAIL.n146 VSUBS 0.0126f
C207 VTAIL.n147 VSUBS 0.028127f
C208 VTAIL.n148 VSUBS 0.028127f
C209 VTAIL.n149 VSUBS 0.0126f
C210 VTAIL.n150 VSUBS 0.0119f
C211 VTAIL.n151 VSUBS 0.022145f
C212 VTAIL.n152 VSUBS 0.022145f
C213 VTAIL.n153 VSUBS 0.0119f
C214 VTAIL.n154 VSUBS 0.0126f
C215 VTAIL.n155 VSUBS 0.028127f
C216 VTAIL.n156 VSUBS 0.028127f
C217 VTAIL.n157 VSUBS 0.0126f
C218 VTAIL.n158 VSUBS 0.0119f
C219 VTAIL.n159 VSUBS 0.022145f
C220 VTAIL.n160 VSUBS 0.022145f
C221 VTAIL.n161 VSUBS 0.0119f
C222 VTAIL.n162 VSUBS 0.0126f
C223 VTAIL.n163 VSUBS 0.028127f
C224 VTAIL.n164 VSUBS 0.028127f
C225 VTAIL.n165 VSUBS 0.028127f
C226 VTAIL.n166 VSUBS 0.0126f
C227 VTAIL.n167 VSUBS 0.0119f
C228 VTAIL.n168 VSUBS 0.022145f
C229 VTAIL.n169 VSUBS 0.022145f
C230 VTAIL.n170 VSUBS 0.0119f
C231 VTAIL.n171 VSUBS 0.01225f
C232 VTAIL.n172 VSUBS 0.01225f
C233 VTAIL.n173 VSUBS 0.028127f
C234 VTAIL.n174 VSUBS 0.028127f
C235 VTAIL.n175 VSUBS 0.0126f
C236 VTAIL.n176 VSUBS 0.0119f
C237 VTAIL.n177 VSUBS 0.022145f
C238 VTAIL.n178 VSUBS 0.022145f
C239 VTAIL.n179 VSUBS 0.0119f
C240 VTAIL.n180 VSUBS 0.0126f
C241 VTAIL.n181 VSUBS 0.028127f
C242 VTAIL.n182 VSUBS 0.066499f
C243 VTAIL.n183 VSUBS 0.0126f
C244 VTAIL.n184 VSUBS 0.0119f
C245 VTAIL.n185 VSUBS 0.052398f
C246 VTAIL.n186 VSUBS 0.033408f
C247 VTAIL.n187 VSUBS 0.190302f
C248 VTAIL.n188 VSUBS 0.023865f
C249 VTAIL.n189 VSUBS 0.022145f
C250 VTAIL.n190 VSUBS 0.0119f
C251 VTAIL.n191 VSUBS 0.028127f
C252 VTAIL.n192 VSUBS 0.0126f
C253 VTAIL.n193 VSUBS 0.022145f
C254 VTAIL.n194 VSUBS 0.0119f
C255 VTAIL.n195 VSUBS 0.028127f
C256 VTAIL.n196 VSUBS 0.0126f
C257 VTAIL.n197 VSUBS 0.022145f
C258 VTAIL.n198 VSUBS 0.0119f
C259 VTAIL.n199 VSUBS 0.028127f
C260 VTAIL.n200 VSUBS 0.0126f
C261 VTAIL.n201 VSUBS 0.022145f
C262 VTAIL.n202 VSUBS 0.0119f
C263 VTAIL.n203 VSUBS 0.028127f
C264 VTAIL.n204 VSUBS 0.0126f
C265 VTAIL.n205 VSUBS 0.022145f
C266 VTAIL.n206 VSUBS 0.0119f
C267 VTAIL.n207 VSUBS 0.028127f
C268 VTAIL.n208 VSUBS 0.0126f
C269 VTAIL.n209 VSUBS 0.022145f
C270 VTAIL.n210 VSUBS 0.0119f
C271 VTAIL.n211 VSUBS 0.028127f
C272 VTAIL.n212 VSUBS 0.0126f
C273 VTAIL.n213 VSUBS 0.022145f
C274 VTAIL.n214 VSUBS 0.0119f
C275 VTAIL.n215 VSUBS 0.028127f
C276 VTAIL.n216 VSUBS 0.0126f
C277 VTAIL.n217 VSUBS 0.168125f
C278 VTAIL.t3 VSUBS 0.060316f
C279 VTAIL.n218 VSUBS 0.021096f
C280 VTAIL.n219 VSUBS 0.017893f
C281 VTAIL.n220 VSUBS 0.0119f
C282 VTAIL.n221 VSUBS 1.59902f
C283 VTAIL.n222 VSUBS 0.022145f
C284 VTAIL.n223 VSUBS 0.0119f
C285 VTAIL.n224 VSUBS 0.0126f
C286 VTAIL.n225 VSUBS 0.028127f
C287 VTAIL.n226 VSUBS 0.028127f
C288 VTAIL.n227 VSUBS 0.0126f
C289 VTAIL.n228 VSUBS 0.0119f
C290 VTAIL.n229 VSUBS 0.022145f
C291 VTAIL.n230 VSUBS 0.022145f
C292 VTAIL.n231 VSUBS 0.0119f
C293 VTAIL.n232 VSUBS 0.0126f
C294 VTAIL.n233 VSUBS 0.028127f
C295 VTAIL.n234 VSUBS 0.028127f
C296 VTAIL.n235 VSUBS 0.0126f
C297 VTAIL.n236 VSUBS 0.0119f
C298 VTAIL.n237 VSUBS 0.022145f
C299 VTAIL.n238 VSUBS 0.022145f
C300 VTAIL.n239 VSUBS 0.0119f
C301 VTAIL.n240 VSUBS 0.0126f
C302 VTAIL.n241 VSUBS 0.028127f
C303 VTAIL.n242 VSUBS 0.028127f
C304 VTAIL.n243 VSUBS 0.0126f
C305 VTAIL.n244 VSUBS 0.0119f
C306 VTAIL.n245 VSUBS 0.022145f
C307 VTAIL.n246 VSUBS 0.022145f
C308 VTAIL.n247 VSUBS 0.0119f
C309 VTAIL.n248 VSUBS 0.0126f
C310 VTAIL.n249 VSUBS 0.028127f
C311 VTAIL.n250 VSUBS 0.028127f
C312 VTAIL.n251 VSUBS 0.0126f
C313 VTAIL.n252 VSUBS 0.0119f
C314 VTAIL.n253 VSUBS 0.022145f
C315 VTAIL.n254 VSUBS 0.022145f
C316 VTAIL.n255 VSUBS 0.0119f
C317 VTAIL.n256 VSUBS 0.0126f
C318 VTAIL.n257 VSUBS 0.028127f
C319 VTAIL.n258 VSUBS 0.028127f
C320 VTAIL.n259 VSUBS 0.028127f
C321 VTAIL.n260 VSUBS 0.0126f
C322 VTAIL.n261 VSUBS 0.0119f
C323 VTAIL.n262 VSUBS 0.022145f
C324 VTAIL.n263 VSUBS 0.022145f
C325 VTAIL.n264 VSUBS 0.0119f
C326 VTAIL.n265 VSUBS 0.01225f
C327 VTAIL.n266 VSUBS 0.01225f
C328 VTAIL.n267 VSUBS 0.028127f
C329 VTAIL.n268 VSUBS 0.028127f
C330 VTAIL.n269 VSUBS 0.0126f
C331 VTAIL.n270 VSUBS 0.0119f
C332 VTAIL.n271 VSUBS 0.022145f
C333 VTAIL.n272 VSUBS 0.022145f
C334 VTAIL.n273 VSUBS 0.0119f
C335 VTAIL.n274 VSUBS 0.0126f
C336 VTAIL.n275 VSUBS 0.028127f
C337 VTAIL.n276 VSUBS 0.066499f
C338 VTAIL.n277 VSUBS 0.0126f
C339 VTAIL.n278 VSUBS 0.0119f
C340 VTAIL.n279 VSUBS 0.052398f
C341 VTAIL.n280 VSUBS 0.033408f
C342 VTAIL.n281 VSUBS 1.63069f
C343 VTAIL.n282 VSUBS 0.023865f
C344 VTAIL.n283 VSUBS 0.022145f
C345 VTAIL.n284 VSUBS 0.0119f
C346 VTAIL.n285 VSUBS 0.028127f
C347 VTAIL.n286 VSUBS 0.0126f
C348 VTAIL.n287 VSUBS 0.022145f
C349 VTAIL.n288 VSUBS 0.0119f
C350 VTAIL.n289 VSUBS 0.028127f
C351 VTAIL.n290 VSUBS 0.0126f
C352 VTAIL.n291 VSUBS 0.022145f
C353 VTAIL.n292 VSUBS 0.0119f
C354 VTAIL.n293 VSUBS 0.028127f
C355 VTAIL.n294 VSUBS 0.028127f
C356 VTAIL.n295 VSUBS 0.0126f
C357 VTAIL.n296 VSUBS 0.022145f
C358 VTAIL.n297 VSUBS 0.0119f
C359 VTAIL.n298 VSUBS 0.028127f
C360 VTAIL.n299 VSUBS 0.0126f
C361 VTAIL.n300 VSUBS 0.022145f
C362 VTAIL.n301 VSUBS 0.0119f
C363 VTAIL.n302 VSUBS 0.028127f
C364 VTAIL.n303 VSUBS 0.0126f
C365 VTAIL.n304 VSUBS 0.022145f
C366 VTAIL.n305 VSUBS 0.0119f
C367 VTAIL.n306 VSUBS 0.028127f
C368 VTAIL.n307 VSUBS 0.0126f
C369 VTAIL.n308 VSUBS 0.022145f
C370 VTAIL.n309 VSUBS 0.0119f
C371 VTAIL.n310 VSUBS 0.028127f
C372 VTAIL.n311 VSUBS 0.0126f
C373 VTAIL.n312 VSUBS 0.168125f
C374 VTAIL.t6 VSUBS 0.060316f
C375 VTAIL.n313 VSUBS 0.021096f
C376 VTAIL.n314 VSUBS 0.017893f
C377 VTAIL.n315 VSUBS 0.0119f
C378 VTAIL.n316 VSUBS 1.59902f
C379 VTAIL.n317 VSUBS 0.022145f
C380 VTAIL.n318 VSUBS 0.0119f
C381 VTAIL.n319 VSUBS 0.0126f
C382 VTAIL.n320 VSUBS 0.028127f
C383 VTAIL.n321 VSUBS 0.028127f
C384 VTAIL.n322 VSUBS 0.0126f
C385 VTAIL.n323 VSUBS 0.0119f
C386 VTAIL.n324 VSUBS 0.022145f
C387 VTAIL.n325 VSUBS 0.022145f
C388 VTAIL.n326 VSUBS 0.0119f
C389 VTAIL.n327 VSUBS 0.0126f
C390 VTAIL.n328 VSUBS 0.028127f
C391 VTAIL.n329 VSUBS 0.028127f
C392 VTAIL.n330 VSUBS 0.0126f
C393 VTAIL.n331 VSUBS 0.0119f
C394 VTAIL.n332 VSUBS 0.022145f
C395 VTAIL.n333 VSUBS 0.022145f
C396 VTAIL.n334 VSUBS 0.0119f
C397 VTAIL.n335 VSUBS 0.0126f
C398 VTAIL.n336 VSUBS 0.028127f
C399 VTAIL.n337 VSUBS 0.028127f
C400 VTAIL.n338 VSUBS 0.0126f
C401 VTAIL.n339 VSUBS 0.0119f
C402 VTAIL.n340 VSUBS 0.022145f
C403 VTAIL.n341 VSUBS 0.022145f
C404 VTAIL.n342 VSUBS 0.0119f
C405 VTAIL.n343 VSUBS 0.0126f
C406 VTAIL.n344 VSUBS 0.028127f
C407 VTAIL.n345 VSUBS 0.028127f
C408 VTAIL.n346 VSUBS 0.0126f
C409 VTAIL.n347 VSUBS 0.0119f
C410 VTAIL.n348 VSUBS 0.022145f
C411 VTAIL.n349 VSUBS 0.022145f
C412 VTAIL.n350 VSUBS 0.0119f
C413 VTAIL.n351 VSUBS 0.0126f
C414 VTAIL.n352 VSUBS 0.028127f
C415 VTAIL.n353 VSUBS 0.028127f
C416 VTAIL.n354 VSUBS 0.0126f
C417 VTAIL.n355 VSUBS 0.0119f
C418 VTAIL.n356 VSUBS 0.022145f
C419 VTAIL.n357 VSUBS 0.022145f
C420 VTAIL.n358 VSUBS 0.0119f
C421 VTAIL.n359 VSUBS 0.01225f
C422 VTAIL.n360 VSUBS 0.01225f
C423 VTAIL.n361 VSUBS 0.028127f
C424 VTAIL.n362 VSUBS 0.028127f
C425 VTAIL.n363 VSUBS 0.0126f
C426 VTAIL.n364 VSUBS 0.0119f
C427 VTAIL.n365 VSUBS 0.022145f
C428 VTAIL.n366 VSUBS 0.022145f
C429 VTAIL.n367 VSUBS 0.0119f
C430 VTAIL.n368 VSUBS 0.0126f
C431 VTAIL.n369 VSUBS 0.028127f
C432 VTAIL.n370 VSUBS 0.066499f
C433 VTAIL.n371 VSUBS 0.0126f
C434 VTAIL.n372 VSUBS 0.0119f
C435 VTAIL.n373 VSUBS 0.052398f
C436 VTAIL.n374 VSUBS 0.033408f
C437 VTAIL.n375 VSUBS 1.63069f
C438 VTAIL.n376 VSUBS 0.023865f
C439 VTAIL.n377 VSUBS 0.022145f
C440 VTAIL.n378 VSUBS 0.0119f
C441 VTAIL.n379 VSUBS 0.028127f
C442 VTAIL.n380 VSUBS 0.0126f
C443 VTAIL.n381 VSUBS 0.022145f
C444 VTAIL.n382 VSUBS 0.0119f
C445 VTAIL.n383 VSUBS 0.028127f
C446 VTAIL.n384 VSUBS 0.0126f
C447 VTAIL.n385 VSUBS 0.022145f
C448 VTAIL.n386 VSUBS 0.0119f
C449 VTAIL.n387 VSUBS 0.028127f
C450 VTAIL.n388 VSUBS 0.028127f
C451 VTAIL.n389 VSUBS 0.0126f
C452 VTAIL.n390 VSUBS 0.022145f
C453 VTAIL.n391 VSUBS 0.0119f
C454 VTAIL.n392 VSUBS 0.028127f
C455 VTAIL.n393 VSUBS 0.0126f
C456 VTAIL.n394 VSUBS 0.022145f
C457 VTAIL.n395 VSUBS 0.0119f
C458 VTAIL.n396 VSUBS 0.028127f
C459 VTAIL.n397 VSUBS 0.0126f
C460 VTAIL.n398 VSUBS 0.022145f
C461 VTAIL.n399 VSUBS 0.0119f
C462 VTAIL.n400 VSUBS 0.028127f
C463 VTAIL.n401 VSUBS 0.0126f
C464 VTAIL.n402 VSUBS 0.022145f
C465 VTAIL.n403 VSUBS 0.0119f
C466 VTAIL.n404 VSUBS 0.028127f
C467 VTAIL.n405 VSUBS 0.0126f
C468 VTAIL.n406 VSUBS 0.168125f
C469 VTAIL.t4 VSUBS 0.060316f
C470 VTAIL.n407 VSUBS 0.021096f
C471 VTAIL.n408 VSUBS 0.017893f
C472 VTAIL.n409 VSUBS 0.0119f
C473 VTAIL.n410 VSUBS 1.59902f
C474 VTAIL.n411 VSUBS 0.022145f
C475 VTAIL.n412 VSUBS 0.0119f
C476 VTAIL.n413 VSUBS 0.0126f
C477 VTAIL.n414 VSUBS 0.028127f
C478 VTAIL.n415 VSUBS 0.028127f
C479 VTAIL.n416 VSUBS 0.0126f
C480 VTAIL.n417 VSUBS 0.0119f
C481 VTAIL.n418 VSUBS 0.022145f
C482 VTAIL.n419 VSUBS 0.022145f
C483 VTAIL.n420 VSUBS 0.0119f
C484 VTAIL.n421 VSUBS 0.0126f
C485 VTAIL.n422 VSUBS 0.028127f
C486 VTAIL.n423 VSUBS 0.028127f
C487 VTAIL.n424 VSUBS 0.0126f
C488 VTAIL.n425 VSUBS 0.0119f
C489 VTAIL.n426 VSUBS 0.022145f
C490 VTAIL.n427 VSUBS 0.022145f
C491 VTAIL.n428 VSUBS 0.0119f
C492 VTAIL.n429 VSUBS 0.0126f
C493 VTAIL.n430 VSUBS 0.028127f
C494 VTAIL.n431 VSUBS 0.028127f
C495 VTAIL.n432 VSUBS 0.0126f
C496 VTAIL.n433 VSUBS 0.0119f
C497 VTAIL.n434 VSUBS 0.022145f
C498 VTAIL.n435 VSUBS 0.022145f
C499 VTAIL.n436 VSUBS 0.0119f
C500 VTAIL.n437 VSUBS 0.0126f
C501 VTAIL.n438 VSUBS 0.028127f
C502 VTAIL.n439 VSUBS 0.028127f
C503 VTAIL.n440 VSUBS 0.0126f
C504 VTAIL.n441 VSUBS 0.0119f
C505 VTAIL.n442 VSUBS 0.022145f
C506 VTAIL.n443 VSUBS 0.022145f
C507 VTAIL.n444 VSUBS 0.0119f
C508 VTAIL.n445 VSUBS 0.0126f
C509 VTAIL.n446 VSUBS 0.028127f
C510 VTAIL.n447 VSUBS 0.028127f
C511 VTAIL.n448 VSUBS 0.0126f
C512 VTAIL.n449 VSUBS 0.0119f
C513 VTAIL.n450 VSUBS 0.022145f
C514 VTAIL.n451 VSUBS 0.022145f
C515 VTAIL.n452 VSUBS 0.0119f
C516 VTAIL.n453 VSUBS 0.01225f
C517 VTAIL.n454 VSUBS 0.01225f
C518 VTAIL.n455 VSUBS 0.028127f
C519 VTAIL.n456 VSUBS 0.028127f
C520 VTAIL.n457 VSUBS 0.0126f
C521 VTAIL.n458 VSUBS 0.0119f
C522 VTAIL.n459 VSUBS 0.022145f
C523 VTAIL.n460 VSUBS 0.022145f
C524 VTAIL.n461 VSUBS 0.0119f
C525 VTAIL.n462 VSUBS 0.0126f
C526 VTAIL.n463 VSUBS 0.028127f
C527 VTAIL.n464 VSUBS 0.066499f
C528 VTAIL.n465 VSUBS 0.0126f
C529 VTAIL.n466 VSUBS 0.0119f
C530 VTAIL.n467 VSUBS 0.052398f
C531 VTAIL.n468 VSUBS 0.033408f
C532 VTAIL.n469 VSUBS 0.190302f
C533 VTAIL.n470 VSUBS 0.023865f
C534 VTAIL.n471 VSUBS 0.022145f
C535 VTAIL.n472 VSUBS 0.0119f
C536 VTAIL.n473 VSUBS 0.028127f
C537 VTAIL.n474 VSUBS 0.0126f
C538 VTAIL.n475 VSUBS 0.022145f
C539 VTAIL.n476 VSUBS 0.0119f
C540 VTAIL.n477 VSUBS 0.028127f
C541 VTAIL.n478 VSUBS 0.0126f
C542 VTAIL.n479 VSUBS 0.022145f
C543 VTAIL.n480 VSUBS 0.0119f
C544 VTAIL.n481 VSUBS 0.028127f
C545 VTAIL.n482 VSUBS 0.028127f
C546 VTAIL.n483 VSUBS 0.0126f
C547 VTAIL.n484 VSUBS 0.022145f
C548 VTAIL.n485 VSUBS 0.0119f
C549 VTAIL.n486 VSUBS 0.028127f
C550 VTAIL.n487 VSUBS 0.0126f
C551 VTAIL.n488 VSUBS 0.022145f
C552 VTAIL.n489 VSUBS 0.0119f
C553 VTAIL.n490 VSUBS 0.028127f
C554 VTAIL.n491 VSUBS 0.0126f
C555 VTAIL.n492 VSUBS 0.022145f
C556 VTAIL.n493 VSUBS 0.0119f
C557 VTAIL.n494 VSUBS 0.028127f
C558 VTAIL.n495 VSUBS 0.0126f
C559 VTAIL.n496 VSUBS 0.022145f
C560 VTAIL.n497 VSUBS 0.0119f
C561 VTAIL.n498 VSUBS 0.028127f
C562 VTAIL.n499 VSUBS 0.0126f
C563 VTAIL.n500 VSUBS 0.168125f
C564 VTAIL.t2 VSUBS 0.060316f
C565 VTAIL.n501 VSUBS 0.021096f
C566 VTAIL.n502 VSUBS 0.017893f
C567 VTAIL.n503 VSUBS 0.0119f
C568 VTAIL.n504 VSUBS 1.59902f
C569 VTAIL.n505 VSUBS 0.022145f
C570 VTAIL.n506 VSUBS 0.0119f
C571 VTAIL.n507 VSUBS 0.0126f
C572 VTAIL.n508 VSUBS 0.028127f
C573 VTAIL.n509 VSUBS 0.028127f
C574 VTAIL.n510 VSUBS 0.0126f
C575 VTAIL.n511 VSUBS 0.0119f
C576 VTAIL.n512 VSUBS 0.022145f
C577 VTAIL.n513 VSUBS 0.022145f
C578 VTAIL.n514 VSUBS 0.0119f
C579 VTAIL.n515 VSUBS 0.0126f
C580 VTAIL.n516 VSUBS 0.028127f
C581 VTAIL.n517 VSUBS 0.028127f
C582 VTAIL.n518 VSUBS 0.0126f
C583 VTAIL.n519 VSUBS 0.0119f
C584 VTAIL.n520 VSUBS 0.022145f
C585 VTAIL.n521 VSUBS 0.022145f
C586 VTAIL.n522 VSUBS 0.0119f
C587 VTAIL.n523 VSUBS 0.0126f
C588 VTAIL.n524 VSUBS 0.028127f
C589 VTAIL.n525 VSUBS 0.028127f
C590 VTAIL.n526 VSUBS 0.0126f
C591 VTAIL.n527 VSUBS 0.0119f
C592 VTAIL.n528 VSUBS 0.022145f
C593 VTAIL.n529 VSUBS 0.022145f
C594 VTAIL.n530 VSUBS 0.0119f
C595 VTAIL.n531 VSUBS 0.0126f
C596 VTAIL.n532 VSUBS 0.028127f
C597 VTAIL.n533 VSUBS 0.028127f
C598 VTAIL.n534 VSUBS 0.0126f
C599 VTAIL.n535 VSUBS 0.0119f
C600 VTAIL.n536 VSUBS 0.022145f
C601 VTAIL.n537 VSUBS 0.022145f
C602 VTAIL.n538 VSUBS 0.0119f
C603 VTAIL.n539 VSUBS 0.0126f
C604 VTAIL.n540 VSUBS 0.028127f
C605 VTAIL.n541 VSUBS 0.028127f
C606 VTAIL.n542 VSUBS 0.0126f
C607 VTAIL.n543 VSUBS 0.0119f
C608 VTAIL.n544 VSUBS 0.022145f
C609 VTAIL.n545 VSUBS 0.022145f
C610 VTAIL.n546 VSUBS 0.0119f
C611 VTAIL.n547 VSUBS 0.01225f
C612 VTAIL.n548 VSUBS 0.01225f
C613 VTAIL.n549 VSUBS 0.028127f
C614 VTAIL.n550 VSUBS 0.028127f
C615 VTAIL.n551 VSUBS 0.0126f
C616 VTAIL.n552 VSUBS 0.0119f
C617 VTAIL.n553 VSUBS 0.022145f
C618 VTAIL.n554 VSUBS 0.022145f
C619 VTAIL.n555 VSUBS 0.0119f
C620 VTAIL.n556 VSUBS 0.0126f
C621 VTAIL.n557 VSUBS 0.028127f
C622 VTAIL.n558 VSUBS 0.066499f
C623 VTAIL.n559 VSUBS 0.0126f
C624 VTAIL.n560 VSUBS 0.0119f
C625 VTAIL.n561 VSUBS 0.052398f
C626 VTAIL.n562 VSUBS 0.033408f
C627 VTAIL.n563 VSUBS 0.190302f
C628 VTAIL.n564 VSUBS 0.023865f
C629 VTAIL.n565 VSUBS 0.022145f
C630 VTAIL.n566 VSUBS 0.0119f
C631 VTAIL.n567 VSUBS 0.028127f
C632 VTAIL.n568 VSUBS 0.0126f
C633 VTAIL.n569 VSUBS 0.022145f
C634 VTAIL.n570 VSUBS 0.0119f
C635 VTAIL.n571 VSUBS 0.028127f
C636 VTAIL.n572 VSUBS 0.0126f
C637 VTAIL.n573 VSUBS 0.022145f
C638 VTAIL.n574 VSUBS 0.0119f
C639 VTAIL.n575 VSUBS 0.028127f
C640 VTAIL.n576 VSUBS 0.028127f
C641 VTAIL.n577 VSUBS 0.0126f
C642 VTAIL.n578 VSUBS 0.022145f
C643 VTAIL.n579 VSUBS 0.0119f
C644 VTAIL.n580 VSUBS 0.028127f
C645 VTAIL.n581 VSUBS 0.0126f
C646 VTAIL.n582 VSUBS 0.022145f
C647 VTAIL.n583 VSUBS 0.0119f
C648 VTAIL.n584 VSUBS 0.028127f
C649 VTAIL.n585 VSUBS 0.0126f
C650 VTAIL.n586 VSUBS 0.022145f
C651 VTAIL.n587 VSUBS 0.0119f
C652 VTAIL.n588 VSUBS 0.028127f
C653 VTAIL.n589 VSUBS 0.0126f
C654 VTAIL.n590 VSUBS 0.022145f
C655 VTAIL.n591 VSUBS 0.0119f
C656 VTAIL.n592 VSUBS 0.028127f
C657 VTAIL.n593 VSUBS 0.0126f
C658 VTAIL.n594 VSUBS 0.168125f
C659 VTAIL.t1 VSUBS 0.060316f
C660 VTAIL.n595 VSUBS 0.021096f
C661 VTAIL.n596 VSUBS 0.017893f
C662 VTAIL.n597 VSUBS 0.0119f
C663 VTAIL.n598 VSUBS 1.59902f
C664 VTAIL.n599 VSUBS 0.022145f
C665 VTAIL.n600 VSUBS 0.0119f
C666 VTAIL.n601 VSUBS 0.0126f
C667 VTAIL.n602 VSUBS 0.028127f
C668 VTAIL.n603 VSUBS 0.028127f
C669 VTAIL.n604 VSUBS 0.0126f
C670 VTAIL.n605 VSUBS 0.0119f
C671 VTAIL.n606 VSUBS 0.022145f
C672 VTAIL.n607 VSUBS 0.022145f
C673 VTAIL.n608 VSUBS 0.0119f
C674 VTAIL.n609 VSUBS 0.0126f
C675 VTAIL.n610 VSUBS 0.028127f
C676 VTAIL.n611 VSUBS 0.028127f
C677 VTAIL.n612 VSUBS 0.0126f
C678 VTAIL.n613 VSUBS 0.0119f
C679 VTAIL.n614 VSUBS 0.022145f
C680 VTAIL.n615 VSUBS 0.022145f
C681 VTAIL.n616 VSUBS 0.0119f
C682 VTAIL.n617 VSUBS 0.0126f
C683 VTAIL.n618 VSUBS 0.028127f
C684 VTAIL.n619 VSUBS 0.028127f
C685 VTAIL.n620 VSUBS 0.0126f
C686 VTAIL.n621 VSUBS 0.0119f
C687 VTAIL.n622 VSUBS 0.022145f
C688 VTAIL.n623 VSUBS 0.022145f
C689 VTAIL.n624 VSUBS 0.0119f
C690 VTAIL.n625 VSUBS 0.0126f
C691 VTAIL.n626 VSUBS 0.028127f
C692 VTAIL.n627 VSUBS 0.028127f
C693 VTAIL.n628 VSUBS 0.0126f
C694 VTAIL.n629 VSUBS 0.0119f
C695 VTAIL.n630 VSUBS 0.022145f
C696 VTAIL.n631 VSUBS 0.022145f
C697 VTAIL.n632 VSUBS 0.0119f
C698 VTAIL.n633 VSUBS 0.0126f
C699 VTAIL.n634 VSUBS 0.028127f
C700 VTAIL.n635 VSUBS 0.028127f
C701 VTAIL.n636 VSUBS 0.0126f
C702 VTAIL.n637 VSUBS 0.0119f
C703 VTAIL.n638 VSUBS 0.022145f
C704 VTAIL.n639 VSUBS 0.022145f
C705 VTAIL.n640 VSUBS 0.0119f
C706 VTAIL.n641 VSUBS 0.01225f
C707 VTAIL.n642 VSUBS 0.01225f
C708 VTAIL.n643 VSUBS 0.028127f
C709 VTAIL.n644 VSUBS 0.028127f
C710 VTAIL.n645 VSUBS 0.0126f
C711 VTAIL.n646 VSUBS 0.0119f
C712 VTAIL.n647 VSUBS 0.022145f
C713 VTAIL.n648 VSUBS 0.022145f
C714 VTAIL.n649 VSUBS 0.0119f
C715 VTAIL.n650 VSUBS 0.0126f
C716 VTAIL.n651 VSUBS 0.028127f
C717 VTAIL.n652 VSUBS 0.066499f
C718 VTAIL.n653 VSUBS 0.0126f
C719 VTAIL.n654 VSUBS 0.0119f
C720 VTAIL.n655 VSUBS 0.052398f
C721 VTAIL.n656 VSUBS 0.033408f
C722 VTAIL.n657 VSUBS 1.63069f
C723 VTAIL.n658 VSUBS 0.023865f
C724 VTAIL.n659 VSUBS 0.022145f
C725 VTAIL.n660 VSUBS 0.0119f
C726 VTAIL.n661 VSUBS 0.028127f
C727 VTAIL.n662 VSUBS 0.0126f
C728 VTAIL.n663 VSUBS 0.022145f
C729 VTAIL.n664 VSUBS 0.0119f
C730 VTAIL.n665 VSUBS 0.028127f
C731 VTAIL.n666 VSUBS 0.0126f
C732 VTAIL.n667 VSUBS 0.022145f
C733 VTAIL.n668 VSUBS 0.0119f
C734 VTAIL.n669 VSUBS 0.028127f
C735 VTAIL.n670 VSUBS 0.0126f
C736 VTAIL.n671 VSUBS 0.022145f
C737 VTAIL.n672 VSUBS 0.0119f
C738 VTAIL.n673 VSUBS 0.028127f
C739 VTAIL.n674 VSUBS 0.0126f
C740 VTAIL.n675 VSUBS 0.022145f
C741 VTAIL.n676 VSUBS 0.0119f
C742 VTAIL.n677 VSUBS 0.028127f
C743 VTAIL.n678 VSUBS 0.0126f
C744 VTAIL.n679 VSUBS 0.022145f
C745 VTAIL.n680 VSUBS 0.0119f
C746 VTAIL.n681 VSUBS 0.028127f
C747 VTAIL.n682 VSUBS 0.0126f
C748 VTAIL.n683 VSUBS 0.022145f
C749 VTAIL.n684 VSUBS 0.0119f
C750 VTAIL.n685 VSUBS 0.028127f
C751 VTAIL.n686 VSUBS 0.0126f
C752 VTAIL.n687 VSUBS 0.168125f
C753 VTAIL.t7 VSUBS 0.060316f
C754 VTAIL.n688 VSUBS 0.021096f
C755 VTAIL.n689 VSUBS 0.017893f
C756 VTAIL.n690 VSUBS 0.0119f
C757 VTAIL.n691 VSUBS 1.59902f
C758 VTAIL.n692 VSUBS 0.022145f
C759 VTAIL.n693 VSUBS 0.0119f
C760 VTAIL.n694 VSUBS 0.0126f
C761 VTAIL.n695 VSUBS 0.028127f
C762 VTAIL.n696 VSUBS 0.028127f
C763 VTAIL.n697 VSUBS 0.0126f
C764 VTAIL.n698 VSUBS 0.0119f
C765 VTAIL.n699 VSUBS 0.022145f
C766 VTAIL.n700 VSUBS 0.022145f
C767 VTAIL.n701 VSUBS 0.0119f
C768 VTAIL.n702 VSUBS 0.0126f
C769 VTAIL.n703 VSUBS 0.028127f
C770 VTAIL.n704 VSUBS 0.028127f
C771 VTAIL.n705 VSUBS 0.0126f
C772 VTAIL.n706 VSUBS 0.0119f
C773 VTAIL.n707 VSUBS 0.022145f
C774 VTAIL.n708 VSUBS 0.022145f
C775 VTAIL.n709 VSUBS 0.0119f
C776 VTAIL.n710 VSUBS 0.0126f
C777 VTAIL.n711 VSUBS 0.028127f
C778 VTAIL.n712 VSUBS 0.028127f
C779 VTAIL.n713 VSUBS 0.0126f
C780 VTAIL.n714 VSUBS 0.0119f
C781 VTAIL.n715 VSUBS 0.022145f
C782 VTAIL.n716 VSUBS 0.022145f
C783 VTAIL.n717 VSUBS 0.0119f
C784 VTAIL.n718 VSUBS 0.0126f
C785 VTAIL.n719 VSUBS 0.028127f
C786 VTAIL.n720 VSUBS 0.028127f
C787 VTAIL.n721 VSUBS 0.0126f
C788 VTAIL.n722 VSUBS 0.0119f
C789 VTAIL.n723 VSUBS 0.022145f
C790 VTAIL.n724 VSUBS 0.022145f
C791 VTAIL.n725 VSUBS 0.0119f
C792 VTAIL.n726 VSUBS 0.0126f
C793 VTAIL.n727 VSUBS 0.028127f
C794 VTAIL.n728 VSUBS 0.028127f
C795 VTAIL.n729 VSUBS 0.028127f
C796 VTAIL.n730 VSUBS 0.0126f
C797 VTAIL.n731 VSUBS 0.0119f
C798 VTAIL.n732 VSUBS 0.022145f
C799 VTAIL.n733 VSUBS 0.022145f
C800 VTAIL.n734 VSUBS 0.0119f
C801 VTAIL.n735 VSUBS 0.01225f
C802 VTAIL.n736 VSUBS 0.01225f
C803 VTAIL.n737 VSUBS 0.028127f
C804 VTAIL.n738 VSUBS 0.028127f
C805 VTAIL.n739 VSUBS 0.0126f
C806 VTAIL.n740 VSUBS 0.0119f
C807 VTAIL.n741 VSUBS 0.022145f
C808 VTAIL.n742 VSUBS 0.022145f
C809 VTAIL.n743 VSUBS 0.0119f
C810 VTAIL.n744 VSUBS 0.0126f
C811 VTAIL.n745 VSUBS 0.028127f
C812 VTAIL.n746 VSUBS 0.066499f
C813 VTAIL.n747 VSUBS 0.0126f
C814 VTAIL.n748 VSUBS 0.0119f
C815 VTAIL.n749 VSUBS 0.052398f
C816 VTAIL.n750 VSUBS 0.033408f
C817 VTAIL.n751 VSUBS 1.55795f
C818 VN.t2 VSUBS 3.3557f
C819 VN.t0 VSUBS 3.35298f
C820 VN.n0 VSUBS 2.2995f
C821 VN.t3 VSUBS 3.3557f
C822 VN.t1 VSUBS 3.35298f
C823 VN.n1 VSUBS 4.13547f
C824 B.n0 VSUBS 0.005825f
C825 B.n1 VSUBS 0.005825f
C826 B.n2 VSUBS 0.008614f
C827 B.n3 VSUBS 0.006601f
C828 B.n4 VSUBS 0.006601f
C829 B.n5 VSUBS 0.006601f
C830 B.n6 VSUBS 0.006601f
C831 B.n7 VSUBS 0.006601f
C832 B.n8 VSUBS 0.006601f
C833 B.n9 VSUBS 0.006601f
C834 B.n10 VSUBS 0.006601f
C835 B.n11 VSUBS 0.006601f
C836 B.n12 VSUBS 0.006601f
C837 B.n13 VSUBS 0.006601f
C838 B.n14 VSUBS 0.006601f
C839 B.n15 VSUBS 0.016383f
C840 B.n16 VSUBS 0.006601f
C841 B.n17 VSUBS 0.006601f
C842 B.n18 VSUBS 0.006601f
C843 B.n19 VSUBS 0.006601f
C844 B.n20 VSUBS 0.006601f
C845 B.n21 VSUBS 0.006601f
C846 B.n22 VSUBS 0.006601f
C847 B.n23 VSUBS 0.006601f
C848 B.n24 VSUBS 0.006601f
C849 B.n25 VSUBS 0.006601f
C850 B.n26 VSUBS 0.006601f
C851 B.n27 VSUBS 0.006601f
C852 B.n28 VSUBS 0.006601f
C853 B.n29 VSUBS 0.006601f
C854 B.n30 VSUBS 0.006601f
C855 B.n31 VSUBS 0.006601f
C856 B.n32 VSUBS 0.006601f
C857 B.n33 VSUBS 0.006601f
C858 B.n34 VSUBS 0.006601f
C859 B.n35 VSUBS 0.006601f
C860 B.n36 VSUBS 0.006601f
C861 B.n37 VSUBS 0.006601f
C862 B.n38 VSUBS 0.006601f
C863 B.n39 VSUBS 0.006601f
C864 B.n40 VSUBS 0.006601f
C865 B.n41 VSUBS 0.006601f
C866 B.n42 VSUBS 0.006601f
C867 B.n43 VSUBS 0.006601f
C868 B.t1 VSUBS 0.30477f
C869 B.t2 VSUBS 0.329091f
C870 B.t0 VSUBS 1.31288f
C871 B.n44 VSUBS 0.485122f
C872 B.n45 VSUBS 0.294004f
C873 B.n46 VSUBS 0.006601f
C874 B.n47 VSUBS 0.006601f
C875 B.n48 VSUBS 0.006601f
C876 B.n49 VSUBS 0.006601f
C877 B.t4 VSUBS 0.304774f
C878 B.t5 VSUBS 0.329094f
C879 B.t3 VSUBS 1.31288f
C880 B.n50 VSUBS 0.485119f
C881 B.n51 VSUBS 0.294001f
C882 B.n52 VSUBS 0.015294f
C883 B.n53 VSUBS 0.006601f
C884 B.n54 VSUBS 0.006601f
C885 B.n55 VSUBS 0.006601f
C886 B.n56 VSUBS 0.006601f
C887 B.n57 VSUBS 0.006601f
C888 B.n58 VSUBS 0.006601f
C889 B.n59 VSUBS 0.006601f
C890 B.n60 VSUBS 0.006601f
C891 B.n61 VSUBS 0.006601f
C892 B.n62 VSUBS 0.006601f
C893 B.n63 VSUBS 0.006601f
C894 B.n64 VSUBS 0.006601f
C895 B.n65 VSUBS 0.006601f
C896 B.n66 VSUBS 0.006601f
C897 B.n67 VSUBS 0.006601f
C898 B.n68 VSUBS 0.006601f
C899 B.n69 VSUBS 0.006601f
C900 B.n70 VSUBS 0.006601f
C901 B.n71 VSUBS 0.006601f
C902 B.n72 VSUBS 0.006601f
C903 B.n73 VSUBS 0.006601f
C904 B.n74 VSUBS 0.006601f
C905 B.n75 VSUBS 0.006601f
C906 B.n76 VSUBS 0.006601f
C907 B.n77 VSUBS 0.006601f
C908 B.n78 VSUBS 0.006601f
C909 B.n79 VSUBS 0.006601f
C910 B.n80 VSUBS 0.017206f
C911 B.n81 VSUBS 0.006601f
C912 B.n82 VSUBS 0.006601f
C913 B.n83 VSUBS 0.006601f
C914 B.n84 VSUBS 0.006601f
C915 B.n85 VSUBS 0.006601f
C916 B.n86 VSUBS 0.006601f
C917 B.n87 VSUBS 0.006601f
C918 B.n88 VSUBS 0.006601f
C919 B.n89 VSUBS 0.006601f
C920 B.n90 VSUBS 0.006601f
C921 B.n91 VSUBS 0.006601f
C922 B.n92 VSUBS 0.006601f
C923 B.n93 VSUBS 0.006601f
C924 B.n94 VSUBS 0.006601f
C925 B.n95 VSUBS 0.006601f
C926 B.n96 VSUBS 0.006601f
C927 B.n97 VSUBS 0.006601f
C928 B.n98 VSUBS 0.006601f
C929 B.n99 VSUBS 0.006601f
C930 B.n100 VSUBS 0.006601f
C931 B.n101 VSUBS 0.006601f
C932 B.n102 VSUBS 0.006601f
C933 B.n103 VSUBS 0.006601f
C934 B.n104 VSUBS 0.006601f
C935 B.n105 VSUBS 0.006601f
C936 B.n106 VSUBS 0.006601f
C937 B.n107 VSUBS 0.006601f
C938 B.n108 VSUBS 0.017071f
C939 B.n109 VSUBS 0.006601f
C940 B.n110 VSUBS 0.006601f
C941 B.n111 VSUBS 0.006601f
C942 B.n112 VSUBS 0.006601f
C943 B.n113 VSUBS 0.006601f
C944 B.n114 VSUBS 0.006601f
C945 B.n115 VSUBS 0.006601f
C946 B.n116 VSUBS 0.006601f
C947 B.n117 VSUBS 0.006601f
C948 B.n118 VSUBS 0.006601f
C949 B.n119 VSUBS 0.006601f
C950 B.n120 VSUBS 0.006601f
C951 B.n121 VSUBS 0.006601f
C952 B.n122 VSUBS 0.006601f
C953 B.n123 VSUBS 0.006601f
C954 B.n124 VSUBS 0.006601f
C955 B.n125 VSUBS 0.006601f
C956 B.n126 VSUBS 0.006601f
C957 B.n127 VSUBS 0.006601f
C958 B.n128 VSUBS 0.006601f
C959 B.n129 VSUBS 0.006601f
C960 B.n130 VSUBS 0.006601f
C961 B.n131 VSUBS 0.006601f
C962 B.n132 VSUBS 0.006601f
C963 B.n133 VSUBS 0.006601f
C964 B.n134 VSUBS 0.006601f
C965 B.n135 VSUBS 0.006601f
C966 B.n136 VSUBS 0.004563f
C967 B.n137 VSUBS 0.006601f
C968 B.n138 VSUBS 0.006601f
C969 B.n139 VSUBS 0.006601f
C970 B.n140 VSUBS 0.006601f
C971 B.n141 VSUBS 0.006601f
C972 B.t11 VSUBS 0.30477f
C973 B.t10 VSUBS 0.329091f
C974 B.t9 VSUBS 1.31288f
C975 B.n142 VSUBS 0.485122f
C976 B.n143 VSUBS 0.294004f
C977 B.n144 VSUBS 0.006601f
C978 B.n145 VSUBS 0.006601f
C979 B.n146 VSUBS 0.006601f
C980 B.n147 VSUBS 0.006601f
C981 B.n148 VSUBS 0.006601f
C982 B.n149 VSUBS 0.006601f
C983 B.n150 VSUBS 0.006601f
C984 B.n151 VSUBS 0.006601f
C985 B.n152 VSUBS 0.006601f
C986 B.n153 VSUBS 0.006601f
C987 B.n154 VSUBS 0.006601f
C988 B.n155 VSUBS 0.006601f
C989 B.n156 VSUBS 0.006601f
C990 B.n157 VSUBS 0.006601f
C991 B.n158 VSUBS 0.006601f
C992 B.n159 VSUBS 0.006601f
C993 B.n160 VSUBS 0.006601f
C994 B.n161 VSUBS 0.006601f
C995 B.n162 VSUBS 0.006601f
C996 B.n163 VSUBS 0.006601f
C997 B.n164 VSUBS 0.006601f
C998 B.n165 VSUBS 0.006601f
C999 B.n166 VSUBS 0.006601f
C1000 B.n167 VSUBS 0.006601f
C1001 B.n168 VSUBS 0.006601f
C1002 B.n169 VSUBS 0.006601f
C1003 B.n170 VSUBS 0.006601f
C1004 B.n171 VSUBS 0.016383f
C1005 B.n172 VSUBS 0.006601f
C1006 B.n173 VSUBS 0.006601f
C1007 B.n174 VSUBS 0.006601f
C1008 B.n175 VSUBS 0.006601f
C1009 B.n176 VSUBS 0.006601f
C1010 B.n177 VSUBS 0.006601f
C1011 B.n178 VSUBS 0.006601f
C1012 B.n179 VSUBS 0.006601f
C1013 B.n180 VSUBS 0.006601f
C1014 B.n181 VSUBS 0.006601f
C1015 B.n182 VSUBS 0.006601f
C1016 B.n183 VSUBS 0.006601f
C1017 B.n184 VSUBS 0.006601f
C1018 B.n185 VSUBS 0.006601f
C1019 B.n186 VSUBS 0.006601f
C1020 B.n187 VSUBS 0.006601f
C1021 B.n188 VSUBS 0.006601f
C1022 B.n189 VSUBS 0.006601f
C1023 B.n190 VSUBS 0.006601f
C1024 B.n191 VSUBS 0.006601f
C1025 B.n192 VSUBS 0.006601f
C1026 B.n193 VSUBS 0.006601f
C1027 B.n194 VSUBS 0.006601f
C1028 B.n195 VSUBS 0.006601f
C1029 B.n196 VSUBS 0.006601f
C1030 B.n197 VSUBS 0.006601f
C1031 B.n198 VSUBS 0.006601f
C1032 B.n199 VSUBS 0.006601f
C1033 B.n200 VSUBS 0.006601f
C1034 B.n201 VSUBS 0.006601f
C1035 B.n202 VSUBS 0.006601f
C1036 B.n203 VSUBS 0.006601f
C1037 B.n204 VSUBS 0.006601f
C1038 B.n205 VSUBS 0.006601f
C1039 B.n206 VSUBS 0.006601f
C1040 B.n207 VSUBS 0.006601f
C1041 B.n208 VSUBS 0.006601f
C1042 B.n209 VSUBS 0.006601f
C1043 B.n210 VSUBS 0.006601f
C1044 B.n211 VSUBS 0.006601f
C1045 B.n212 VSUBS 0.006601f
C1046 B.n213 VSUBS 0.006601f
C1047 B.n214 VSUBS 0.006601f
C1048 B.n215 VSUBS 0.006601f
C1049 B.n216 VSUBS 0.006601f
C1050 B.n217 VSUBS 0.006601f
C1051 B.n218 VSUBS 0.006601f
C1052 B.n219 VSUBS 0.006601f
C1053 B.n220 VSUBS 0.006601f
C1054 B.n221 VSUBS 0.006601f
C1055 B.n222 VSUBS 0.016383f
C1056 B.n223 VSUBS 0.017206f
C1057 B.n224 VSUBS 0.017206f
C1058 B.n225 VSUBS 0.006601f
C1059 B.n226 VSUBS 0.006601f
C1060 B.n227 VSUBS 0.006601f
C1061 B.n228 VSUBS 0.006601f
C1062 B.n229 VSUBS 0.006601f
C1063 B.n230 VSUBS 0.006601f
C1064 B.n231 VSUBS 0.006601f
C1065 B.n232 VSUBS 0.006601f
C1066 B.n233 VSUBS 0.006601f
C1067 B.n234 VSUBS 0.006601f
C1068 B.n235 VSUBS 0.006601f
C1069 B.n236 VSUBS 0.006601f
C1070 B.n237 VSUBS 0.006601f
C1071 B.n238 VSUBS 0.006601f
C1072 B.n239 VSUBS 0.006601f
C1073 B.n240 VSUBS 0.006601f
C1074 B.n241 VSUBS 0.006601f
C1075 B.n242 VSUBS 0.006601f
C1076 B.n243 VSUBS 0.006601f
C1077 B.n244 VSUBS 0.006601f
C1078 B.n245 VSUBS 0.006601f
C1079 B.n246 VSUBS 0.006601f
C1080 B.n247 VSUBS 0.006601f
C1081 B.n248 VSUBS 0.006601f
C1082 B.n249 VSUBS 0.006601f
C1083 B.n250 VSUBS 0.006601f
C1084 B.n251 VSUBS 0.006601f
C1085 B.n252 VSUBS 0.006601f
C1086 B.n253 VSUBS 0.006601f
C1087 B.n254 VSUBS 0.006601f
C1088 B.n255 VSUBS 0.006601f
C1089 B.n256 VSUBS 0.006601f
C1090 B.n257 VSUBS 0.006601f
C1091 B.n258 VSUBS 0.006601f
C1092 B.n259 VSUBS 0.006601f
C1093 B.n260 VSUBS 0.006601f
C1094 B.n261 VSUBS 0.006601f
C1095 B.n262 VSUBS 0.006601f
C1096 B.n263 VSUBS 0.006601f
C1097 B.n264 VSUBS 0.006601f
C1098 B.n265 VSUBS 0.006601f
C1099 B.n266 VSUBS 0.006601f
C1100 B.n267 VSUBS 0.006601f
C1101 B.n268 VSUBS 0.006601f
C1102 B.n269 VSUBS 0.006601f
C1103 B.n270 VSUBS 0.006601f
C1104 B.n271 VSUBS 0.006601f
C1105 B.n272 VSUBS 0.006601f
C1106 B.n273 VSUBS 0.006601f
C1107 B.n274 VSUBS 0.006601f
C1108 B.n275 VSUBS 0.006601f
C1109 B.n276 VSUBS 0.006601f
C1110 B.n277 VSUBS 0.006601f
C1111 B.n278 VSUBS 0.006601f
C1112 B.n279 VSUBS 0.006601f
C1113 B.n280 VSUBS 0.006601f
C1114 B.n281 VSUBS 0.006601f
C1115 B.n282 VSUBS 0.006601f
C1116 B.n283 VSUBS 0.006601f
C1117 B.n284 VSUBS 0.006601f
C1118 B.n285 VSUBS 0.006601f
C1119 B.n286 VSUBS 0.006601f
C1120 B.n287 VSUBS 0.006601f
C1121 B.n288 VSUBS 0.006601f
C1122 B.n289 VSUBS 0.006601f
C1123 B.n290 VSUBS 0.006601f
C1124 B.n291 VSUBS 0.006601f
C1125 B.n292 VSUBS 0.006601f
C1126 B.n293 VSUBS 0.006601f
C1127 B.n294 VSUBS 0.006601f
C1128 B.n295 VSUBS 0.006601f
C1129 B.n296 VSUBS 0.006601f
C1130 B.n297 VSUBS 0.006601f
C1131 B.n298 VSUBS 0.006601f
C1132 B.n299 VSUBS 0.006601f
C1133 B.n300 VSUBS 0.006601f
C1134 B.n301 VSUBS 0.006601f
C1135 B.n302 VSUBS 0.006601f
C1136 B.n303 VSUBS 0.006601f
C1137 B.n304 VSUBS 0.006601f
C1138 B.n305 VSUBS 0.006601f
C1139 B.n306 VSUBS 0.004563f
C1140 B.n307 VSUBS 0.015294f
C1141 B.n308 VSUBS 0.005339f
C1142 B.n309 VSUBS 0.006601f
C1143 B.n310 VSUBS 0.006601f
C1144 B.n311 VSUBS 0.006601f
C1145 B.n312 VSUBS 0.006601f
C1146 B.n313 VSUBS 0.006601f
C1147 B.n314 VSUBS 0.006601f
C1148 B.n315 VSUBS 0.006601f
C1149 B.n316 VSUBS 0.006601f
C1150 B.n317 VSUBS 0.006601f
C1151 B.n318 VSUBS 0.006601f
C1152 B.n319 VSUBS 0.006601f
C1153 B.t8 VSUBS 0.304774f
C1154 B.t7 VSUBS 0.329094f
C1155 B.t6 VSUBS 1.31288f
C1156 B.n320 VSUBS 0.485119f
C1157 B.n321 VSUBS 0.294001f
C1158 B.n322 VSUBS 0.015294f
C1159 B.n323 VSUBS 0.005339f
C1160 B.n324 VSUBS 0.006601f
C1161 B.n325 VSUBS 0.006601f
C1162 B.n326 VSUBS 0.006601f
C1163 B.n327 VSUBS 0.006601f
C1164 B.n328 VSUBS 0.006601f
C1165 B.n329 VSUBS 0.006601f
C1166 B.n330 VSUBS 0.006601f
C1167 B.n331 VSUBS 0.006601f
C1168 B.n332 VSUBS 0.006601f
C1169 B.n333 VSUBS 0.006601f
C1170 B.n334 VSUBS 0.006601f
C1171 B.n335 VSUBS 0.006601f
C1172 B.n336 VSUBS 0.006601f
C1173 B.n337 VSUBS 0.006601f
C1174 B.n338 VSUBS 0.006601f
C1175 B.n339 VSUBS 0.006601f
C1176 B.n340 VSUBS 0.006601f
C1177 B.n341 VSUBS 0.006601f
C1178 B.n342 VSUBS 0.006601f
C1179 B.n343 VSUBS 0.006601f
C1180 B.n344 VSUBS 0.006601f
C1181 B.n345 VSUBS 0.006601f
C1182 B.n346 VSUBS 0.006601f
C1183 B.n347 VSUBS 0.006601f
C1184 B.n348 VSUBS 0.006601f
C1185 B.n349 VSUBS 0.006601f
C1186 B.n350 VSUBS 0.006601f
C1187 B.n351 VSUBS 0.006601f
C1188 B.n352 VSUBS 0.006601f
C1189 B.n353 VSUBS 0.006601f
C1190 B.n354 VSUBS 0.006601f
C1191 B.n355 VSUBS 0.006601f
C1192 B.n356 VSUBS 0.006601f
C1193 B.n357 VSUBS 0.006601f
C1194 B.n358 VSUBS 0.006601f
C1195 B.n359 VSUBS 0.006601f
C1196 B.n360 VSUBS 0.006601f
C1197 B.n361 VSUBS 0.006601f
C1198 B.n362 VSUBS 0.006601f
C1199 B.n363 VSUBS 0.006601f
C1200 B.n364 VSUBS 0.006601f
C1201 B.n365 VSUBS 0.006601f
C1202 B.n366 VSUBS 0.006601f
C1203 B.n367 VSUBS 0.006601f
C1204 B.n368 VSUBS 0.006601f
C1205 B.n369 VSUBS 0.006601f
C1206 B.n370 VSUBS 0.006601f
C1207 B.n371 VSUBS 0.006601f
C1208 B.n372 VSUBS 0.006601f
C1209 B.n373 VSUBS 0.006601f
C1210 B.n374 VSUBS 0.006601f
C1211 B.n375 VSUBS 0.006601f
C1212 B.n376 VSUBS 0.006601f
C1213 B.n377 VSUBS 0.006601f
C1214 B.n378 VSUBS 0.006601f
C1215 B.n379 VSUBS 0.006601f
C1216 B.n380 VSUBS 0.006601f
C1217 B.n381 VSUBS 0.006601f
C1218 B.n382 VSUBS 0.006601f
C1219 B.n383 VSUBS 0.006601f
C1220 B.n384 VSUBS 0.006601f
C1221 B.n385 VSUBS 0.006601f
C1222 B.n386 VSUBS 0.006601f
C1223 B.n387 VSUBS 0.006601f
C1224 B.n388 VSUBS 0.006601f
C1225 B.n389 VSUBS 0.006601f
C1226 B.n390 VSUBS 0.006601f
C1227 B.n391 VSUBS 0.006601f
C1228 B.n392 VSUBS 0.006601f
C1229 B.n393 VSUBS 0.006601f
C1230 B.n394 VSUBS 0.006601f
C1231 B.n395 VSUBS 0.006601f
C1232 B.n396 VSUBS 0.006601f
C1233 B.n397 VSUBS 0.006601f
C1234 B.n398 VSUBS 0.006601f
C1235 B.n399 VSUBS 0.006601f
C1236 B.n400 VSUBS 0.006601f
C1237 B.n401 VSUBS 0.006601f
C1238 B.n402 VSUBS 0.006601f
C1239 B.n403 VSUBS 0.006601f
C1240 B.n404 VSUBS 0.006601f
C1241 B.n405 VSUBS 0.006601f
C1242 B.n406 VSUBS 0.006601f
C1243 B.n407 VSUBS 0.016517f
C1244 B.n408 VSUBS 0.017206f
C1245 B.n409 VSUBS 0.016383f
C1246 B.n410 VSUBS 0.006601f
C1247 B.n411 VSUBS 0.006601f
C1248 B.n412 VSUBS 0.006601f
C1249 B.n413 VSUBS 0.006601f
C1250 B.n414 VSUBS 0.006601f
C1251 B.n415 VSUBS 0.006601f
C1252 B.n416 VSUBS 0.006601f
C1253 B.n417 VSUBS 0.006601f
C1254 B.n418 VSUBS 0.006601f
C1255 B.n419 VSUBS 0.006601f
C1256 B.n420 VSUBS 0.006601f
C1257 B.n421 VSUBS 0.006601f
C1258 B.n422 VSUBS 0.006601f
C1259 B.n423 VSUBS 0.006601f
C1260 B.n424 VSUBS 0.006601f
C1261 B.n425 VSUBS 0.006601f
C1262 B.n426 VSUBS 0.006601f
C1263 B.n427 VSUBS 0.006601f
C1264 B.n428 VSUBS 0.006601f
C1265 B.n429 VSUBS 0.006601f
C1266 B.n430 VSUBS 0.006601f
C1267 B.n431 VSUBS 0.006601f
C1268 B.n432 VSUBS 0.006601f
C1269 B.n433 VSUBS 0.006601f
C1270 B.n434 VSUBS 0.006601f
C1271 B.n435 VSUBS 0.006601f
C1272 B.n436 VSUBS 0.006601f
C1273 B.n437 VSUBS 0.006601f
C1274 B.n438 VSUBS 0.006601f
C1275 B.n439 VSUBS 0.006601f
C1276 B.n440 VSUBS 0.006601f
C1277 B.n441 VSUBS 0.006601f
C1278 B.n442 VSUBS 0.006601f
C1279 B.n443 VSUBS 0.006601f
C1280 B.n444 VSUBS 0.006601f
C1281 B.n445 VSUBS 0.006601f
C1282 B.n446 VSUBS 0.006601f
C1283 B.n447 VSUBS 0.006601f
C1284 B.n448 VSUBS 0.006601f
C1285 B.n449 VSUBS 0.006601f
C1286 B.n450 VSUBS 0.006601f
C1287 B.n451 VSUBS 0.006601f
C1288 B.n452 VSUBS 0.006601f
C1289 B.n453 VSUBS 0.006601f
C1290 B.n454 VSUBS 0.006601f
C1291 B.n455 VSUBS 0.006601f
C1292 B.n456 VSUBS 0.006601f
C1293 B.n457 VSUBS 0.006601f
C1294 B.n458 VSUBS 0.006601f
C1295 B.n459 VSUBS 0.006601f
C1296 B.n460 VSUBS 0.006601f
C1297 B.n461 VSUBS 0.006601f
C1298 B.n462 VSUBS 0.006601f
C1299 B.n463 VSUBS 0.006601f
C1300 B.n464 VSUBS 0.006601f
C1301 B.n465 VSUBS 0.006601f
C1302 B.n466 VSUBS 0.006601f
C1303 B.n467 VSUBS 0.006601f
C1304 B.n468 VSUBS 0.006601f
C1305 B.n469 VSUBS 0.006601f
C1306 B.n470 VSUBS 0.006601f
C1307 B.n471 VSUBS 0.006601f
C1308 B.n472 VSUBS 0.006601f
C1309 B.n473 VSUBS 0.006601f
C1310 B.n474 VSUBS 0.006601f
C1311 B.n475 VSUBS 0.006601f
C1312 B.n476 VSUBS 0.006601f
C1313 B.n477 VSUBS 0.006601f
C1314 B.n478 VSUBS 0.006601f
C1315 B.n479 VSUBS 0.006601f
C1316 B.n480 VSUBS 0.006601f
C1317 B.n481 VSUBS 0.006601f
C1318 B.n482 VSUBS 0.006601f
C1319 B.n483 VSUBS 0.006601f
C1320 B.n484 VSUBS 0.006601f
C1321 B.n485 VSUBS 0.006601f
C1322 B.n486 VSUBS 0.006601f
C1323 B.n487 VSUBS 0.006601f
C1324 B.n488 VSUBS 0.006601f
C1325 B.n489 VSUBS 0.006601f
C1326 B.n490 VSUBS 0.006601f
C1327 B.n491 VSUBS 0.016383f
C1328 B.n492 VSUBS 0.016383f
C1329 B.n493 VSUBS 0.017206f
C1330 B.n494 VSUBS 0.006601f
C1331 B.n495 VSUBS 0.006601f
C1332 B.n496 VSUBS 0.006601f
C1333 B.n497 VSUBS 0.006601f
C1334 B.n498 VSUBS 0.006601f
C1335 B.n499 VSUBS 0.006601f
C1336 B.n500 VSUBS 0.006601f
C1337 B.n501 VSUBS 0.006601f
C1338 B.n502 VSUBS 0.006601f
C1339 B.n503 VSUBS 0.006601f
C1340 B.n504 VSUBS 0.006601f
C1341 B.n505 VSUBS 0.006601f
C1342 B.n506 VSUBS 0.006601f
C1343 B.n507 VSUBS 0.006601f
C1344 B.n508 VSUBS 0.006601f
C1345 B.n509 VSUBS 0.006601f
C1346 B.n510 VSUBS 0.006601f
C1347 B.n511 VSUBS 0.006601f
C1348 B.n512 VSUBS 0.006601f
C1349 B.n513 VSUBS 0.006601f
C1350 B.n514 VSUBS 0.006601f
C1351 B.n515 VSUBS 0.006601f
C1352 B.n516 VSUBS 0.006601f
C1353 B.n517 VSUBS 0.006601f
C1354 B.n518 VSUBS 0.006601f
C1355 B.n519 VSUBS 0.006601f
C1356 B.n520 VSUBS 0.006601f
C1357 B.n521 VSUBS 0.006601f
C1358 B.n522 VSUBS 0.006601f
C1359 B.n523 VSUBS 0.006601f
C1360 B.n524 VSUBS 0.006601f
C1361 B.n525 VSUBS 0.006601f
C1362 B.n526 VSUBS 0.006601f
C1363 B.n527 VSUBS 0.006601f
C1364 B.n528 VSUBS 0.006601f
C1365 B.n529 VSUBS 0.006601f
C1366 B.n530 VSUBS 0.006601f
C1367 B.n531 VSUBS 0.006601f
C1368 B.n532 VSUBS 0.006601f
C1369 B.n533 VSUBS 0.006601f
C1370 B.n534 VSUBS 0.006601f
C1371 B.n535 VSUBS 0.006601f
C1372 B.n536 VSUBS 0.006601f
C1373 B.n537 VSUBS 0.006601f
C1374 B.n538 VSUBS 0.006601f
C1375 B.n539 VSUBS 0.006601f
C1376 B.n540 VSUBS 0.006601f
C1377 B.n541 VSUBS 0.006601f
C1378 B.n542 VSUBS 0.006601f
C1379 B.n543 VSUBS 0.006601f
C1380 B.n544 VSUBS 0.006601f
C1381 B.n545 VSUBS 0.006601f
C1382 B.n546 VSUBS 0.006601f
C1383 B.n547 VSUBS 0.006601f
C1384 B.n548 VSUBS 0.006601f
C1385 B.n549 VSUBS 0.006601f
C1386 B.n550 VSUBS 0.006601f
C1387 B.n551 VSUBS 0.006601f
C1388 B.n552 VSUBS 0.006601f
C1389 B.n553 VSUBS 0.006601f
C1390 B.n554 VSUBS 0.006601f
C1391 B.n555 VSUBS 0.006601f
C1392 B.n556 VSUBS 0.006601f
C1393 B.n557 VSUBS 0.006601f
C1394 B.n558 VSUBS 0.006601f
C1395 B.n559 VSUBS 0.006601f
C1396 B.n560 VSUBS 0.006601f
C1397 B.n561 VSUBS 0.006601f
C1398 B.n562 VSUBS 0.006601f
C1399 B.n563 VSUBS 0.006601f
C1400 B.n564 VSUBS 0.006601f
C1401 B.n565 VSUBS 0.006601f
C1402 B.n566 VSUBS 0.006601f
C1403 B.n567 VSUBS 0.006601f
C1404 B.n568 VSUBS 0.006601f
C1405 B.n569 VSUBS 0.006601f
C1406 B.n570 VSUBS 0.006601f
C1407 B.n571 VSUBS 0.006601f
C1408 B.n572 VSUBS 0.006601f
C1409 B.n573 VSUBS 0.006601f
C1410 B.n574 VSUBS 0.006601f
C1411 B.n575 VSUBS 0.004563f
C1412 B.n576 VSUBS 0.006601f
C1413 B.n577 VSUBS 0.006601f
C1414 B.n578 VSUBS 0.005339f
C1415 B.n579 VSUBS 0.006601f
C1416 B.n580 VSUBS 0.006601f
C1417 B.n581 VSUBS 0.006601f
C1418 B.n582 VSUBS 0.006601f
C1419 B.n583 VSUBS 0.006601f
C1420 B.n584 VSUBS 0.006601f
C1421 B.n585 VSUBS 0.006601f
C1422 B.n586 VSUBS 0.006601f
C1423 B.n587 VSUBS 0.006601f
C1424 B.n588 VSUBS 0.006601f
C1425 B.n589 VSUBS 0.006601f
C1426 B.n590 VSUBS 0.005339f
C1427 B.n591 VSUBS 0.015294f
C1428 B.n592 VSUBS 0.004563f
C1429 B.n593 VSUBS 0.006601f
C1430 B.n594 VSUBS 0.006601f
C1431 B.n595 VSUBS 0.006601f
C1432 B.n596 VSUBS 0.006601f
C1433 B.n597 VSUBS 0.006601f
C1434 B.n598 VSUBS 0.006601f
C1435 B.n599 VSUBS 0.006601f
C1436 B.n600 VSUBS 0.006601f
C1437 B.n601 VSUBS 0.006601f
C1438 B.n602 VSUBS 0.006601f
C1439 B.n603 VSUBS 0.006601f
C1440 B.n604 VSUBS 0.006601f
C1441 B.n605 VSUBS 0.006601f
C1442 B.n606 VSUBS 0.006601f
C1443 B.n607 VSUBS 0.006601f
C1444 B.n608 VSUBS 0.006601f
C1445 B.n609 VSUBS 0.006601f
C1446 B.n610 VSUBS 0.006601f
C1447 B.n611 VSUBS 0.006601f
C1448 B.n612 VSUBS 0.006601f
C1449 B.n613 VSUBS 0.006601f
C1450 B.n614 VSUBS 0.006601f
C1451 B.n615 VSUBS 0.006601f
C1452 B.n616 VSUBS 0.006601f
C1453 B.n617 VSUBS 0.006601f
C1454 B.n618 VSUBS 0.006601f
C1455 B.n619 VSUBS 0.006601f
C1456 B.n620 VSUBS 0.006601f
C1457 B.n621 VSUBS 0.006601f
C1458 B.n622 VSUBS 0.006601f
C1459 B.n623 VSUBS 0.006601f
C1460 B.n624 VSUBS 0.006601f
C1461 B.n625 VSUBS 0.006601f
C1462 B.n626 VSUBS 0.006601f
C1463 B.n627 VSUBS 0.006601f
C1464 B.n628 VSUBS 0.006601f
C1465 B.n629 VSUBS 0.006601f
C1466 B.n630 VSUBS 0.006601f
C1467 B.n631 VSUBS 0.006601f
C1468 B.n632 VSUBS 0.006601f
C1469 B.n633 VSUBS 0.006601f
C1470 B.n634 VSUBS 0.006601f
C1471 B.n635 VSUBS 0.006601f
C1472 B.n636 VSUBS 0.006601f
C1473 B.n637 VSUBS 0.006601f
C1474 B.n638 VSUBS 0.006601f
C1475 B.n639 VSUBS 0.006601f
C1476 B.n640 VSUBS 0.006601f
C1477 B.n641 VSUBS 0.006601f
C1478 B.n642 VSUBS 0.006601f
C1479 B.n643 VSUBS 0.006601f
C1480 B.n644 VSUBS 0.006601f
C1481 B.n645 VSUBS 0.006601f
C1482 B.n646 VSUBS 0.006601f
C1483 B.n647 VSUBS 0.006601f
C1484 B.n648 VSUBS 0.006601f
C1485 B.n649 VSUBS 0.006601f
C1486 B.n650 VSUBS 0.006601f
C1487 B.n651 VSUBS 0.006601f
C1488 B.n652 VSUBS 0.006601f
C1489 B.n653 VSUBS 0.006601f
C1490 B.n654 VSUBS 0.006601f
C1491 B.n655 VSUBS 0.006601f
C1492 B.n656 VSUBS 0.006601f
C1493 B.n657 VSUBS 0.006601f
C1494 B.n658 VSUBS 0.006601f
C1495 B.n659 VSUBS 0.006601f
C1496 B.n660 VSUBS 0.006601f
C1497 B.n661 VSUBS 0.006601f
C1498 B.n662 VSUBS 0.006601f
C1499 B.n663 VSUBS 0.006601f
C1500 B.n664 VSUBS 0.006601f
C1501 B.n665 VSUBS 0.006601f
C1502 B.n666 VSUBS 0.006601f
C1503 B.n667 VSUBS 0.006601f
C1504 B.n668 VSUBS 0.006601f
C1505 B.n669 VSUBS 0.006601f
C1506 B.n670 VSUBS 0.006601f
C1507 B.n671 VSUBS 0.006601f
C1508 B.n672 VSUBS 0.006601f
C1509 B.n673 VSUBS 0.006601f
C1510 B.n674 VSUBS 0.017206f
C1511 B.n675 VSUBS 0.017206f
C1512 B.n676 VSUBS 0.016383f
C1513 B.n677 VSUBS 0.006601f
C1514 B.n678 VSUBS 0.006601f
C1515 B.n679 VSUBS 0.006601f
C1516 B.n680 VSUBS 0.006601f
C1517 B.n681 VSUBS 0.006601f
C1518 B.n682 VSUBS 0.006601f
C1519 B.n683 VSUBS 0.006601f
C1520 B.n684 VSUBS 0.006601f
C1521 B.n685 VSUBS 0.006601f
C1522 B.n686 VSUBS 0.006601f
C1523 B.n687 VSUBS 0.006601f
C1524 B.n688 VSUBS 0.006601f
C1525 B.n689 VSUBS 0.006601f
C1526 B.n690 VSUBS 0.006601f
C1527 B.n691 VSUBS 0.006601f
C1528 B.n692 VSUBS 0.006601f
C1529 B.n693 VSUBS 0.006601f
C1530 B.n694 VSUBS 0.006601f
C1531 B.n695 VSUBS 0.006601f
C1532 B.n696 VSUBS 0.006601f
C1533 B.n697 VSUBS 0.006601f
C1534 B.n698 VSUBS 0.006601f
C1535 B.n699 VSUBS 0.006601f
C1536 B.n700 VSUBS 0.006601f
C1537 B.n701 VSUBS 0.006601f
C1538 B.n702 VSUBS 0.006601f
C1539 B.n703 VSUBS 0.006601f
C1540 B.n704 VSUBS 0.006601f
C1541 B.n705 VSUBS 0.006601f
C1542 B.n706 VSUBS 0.006601f
C1543 B.n707 VSUBS 0.006601f
C1544 B.n708 VSUBS 0.006601f
C1545 B.n709 VSUBS 0.006601f
C1546 B.n710 VSUBS 0.006601f
C1547 B.n711 VSUBS 0.006601f
C1548 B.n712 VSUBS 0.006601f
C1549 B.n713 VSUBS 0.006601f
C1550 B.n714 VSUBS 0.006601f
C1551 B.n715 VSUBS 0.008614f
C1552 B.n716 VSUBS 0.009176f
C1553 B.n717 VSUBS 0.018248f
.ends

