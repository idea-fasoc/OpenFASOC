* NGSPICE file created from diff_pair_sample_0831.ext - technology: sky130A

.subckt diff_pair_sample_0831 VTAIL VN VP B VDD2 VDD1
X0 B.t11 B.t9 B.t10 w_n2030_n4172# sky130_fd_pr__pfet_01v8 ad=6.2478 pd=32.82 as=0 ps=0 w=16.02 l=0.73
X1 VTAIL.t14 VP.t0 VDD1.t1 w_n2030_n4172# sky130_fd_pr__pfet_01v8 ad=6.2478 pd=32.82 as=2.6433 ps=16.35 w=16.02 l=0.73
X2 VDD2.t7 VN.t0 VTAIL.t2 w_n2030_n4172# sky130_fd_pr__pfet_01v8 ad=2.6433 pd=16.35 as=2.6433 ps=16.35 w=16.02 l=0.73
X3 VDD2.t6 VN.t1 VTAIL.t5 w_n2030_n4172# sky130_fd_pr__pfet_01v8 ad=2.6433 pd=16.35 as=6.2478 ps=32.82 w=16.02 l=0.73
X4 VTAIL.t4 VN.t2 VDD2.t5 w_n2030_n4172# sky130_fd_pr__pfet_01v8 ad=6.2478 pd=32.82 as=2.6433 ps=16.35 w=16.02 l=0.73
X5 VTAIL.t3 VN.t3 VDD2.t4 w_n2030_n4172# sky130_fd_pr__pfet_01v8 ad=2.6433 pd=16.35 as=2.6433 ps=16.35 w=16.02 l=0.73
X6 VTAIL.t13 VP.t1 VDD1.t0 w_n2030_n4172# sky130_fd_pr__pfet_01v8 ad=2.6433 pd=16.35 as=2.6433 ps=16.35 w=16.02 l=0.73
X7 B.t8 B.t6 B.t7 w_n2030_n4172# sky130_fd_pr__pfet_01v8 ad=6.2478 pd=32.82 as=0 ps=0 w=16.02 l=0.73
X8 VDD2.t3 VN.t4 VTAIL.t0 w_n2030_n4172# sky130_fd_pr__pfet_01v8 ad=2.6433 pd=16.35 as=6.2478 ps=32.82 w=16.02 l=0.73
X9 VDD2.t2 VN.t5 VTAIL.t1 w_n2030_n4172# sky130_fd_pr__pfet_01v8 ad=2.6433 pd=16.35 as=2.6433 ps=16.35 w=16.02 l=0.73
X10 VDD1.t2 VP.t2 VTAIL.t12 w_n2030_n4172# sky130_fd_pr__pfet_01v8 ad=2.6433 pd=16.35 as=2.6433 ps=16.35 w=16.02 l=0.73
X11 VDD1.t5 VP.t3 VTAIL.t11 w_n2030_n4172# sky130_fd_pr__pfet_01v8 ad=2.6433 pd=16.35 as=2.6433 ps=16.35 w=16.02 l=0.73
X12 VTAIL.t10 VP.t4 VDD1.t4 w_n2030_n4172# sky130_fd_pr__pfet_01v8 ad=6.2478 pd=32.82 as=2.6433 ps=16.35 w=16.02 l=0.73
X13 VTAIL.t9 VP.t5 VDD1.t3 w_n2030_n4172# sky130_fd_pr__pfet_01v8 ad=2.6433 pd=16.35 as=2.6433 ps=16.35 w=16.02 l=0.73
X14 VDD1.t7 VP.t6 VTAIL.t8 w_n2030_n4172# sky130_fd_pr__pfet_01v8 ad=2.6433 pd=16.35 as=6.2478 ps=32.82 w=16.02 l=0.73
X15 B.t5 B.t3 B.t4 w_n2030_n4172# sky130_fd_pr__pfet_01v8 ad=6.2478 pd=32.82 as=0 ps=0 w=16.02 l=0.73
X16 B.t2 B.t0 B.t1 w_n2030_n4172# sky130_fd_pr__pfet_01v8 ad=6.2478 pd=32.82 as=0 ps=0 w=16.02 l=0.73
X17 VDD1.t6 VP.t7 VTAIL.t7 w_n2030_n4172# sky130_fd_pr__pfet_01v8 ad=2.6433 pd=16.35 as=6.2478 ps=32.82 w=16.02 l=0.73
X18 VTAIL.t6 VN.t6 VDD2.t1 w_n2030_n4172# sky130_fd_pr__pfet_01v8 ad=2.6433 pd=16.35 as=2.6433 ps=16.35 w=16.02 l=0.73
X19 VTAIL.t15 VN.t7 VDD2.t0 w_n2030_n4172# sky130_fd_pr__pfet_01v8 ad=6.2478 pd=32.82 as=2.6433 ps=16.35 w=16.02 l=0.73
R0 B.n132 B.t0 731.49
R1 B.n298 B.t9 731.49
R2 B.n48 B.t3 731.49
R3 B.n40 B.t6 731.49
R4 B.n381 B.n100 585
R5 B.n380 B.n379 585
R6 B.n378 B.n101 585
R7 B.n377 B.n376 585
R8 B.n375 B.n102 585
R9 B.n374 B.n373 585
R10 B.n372 B.n103 585
R11 B.n371 B.n370 585
R12 B.n369 B.n104 585
R13 B.n368 B.n367 585
R14 B.n366 B.n105 585
R15 B.n365 B.n364 585
R16 B.n363 B.n106 585
R17 B.n362 B.n361 585
R18 B.n360 B.n107 585
R19 B.n359 B.n358 585
R20 B.n357 B.n108 585
R21 B.n356 B.n355 585
R22 B.n354 B.n109 585
R23 B.n353 B.n352 585
R24 B.n351 B.n110 585
R25 B.n350 B.n349 585
R26 B.n348 B.n111 585
R27 B.n347 B.n346 585
R28 B.n345 B.n112 585
R29 B.n344 B.n343 585
R30 B.n342 B.n113 585
R31 B.n341 B.n340 585
R32 B.n339 B.n114 585
R33 B.n338 B.n337 585
R34 B.n336 B.n115 585
R35 B.n335 B.n334 585
R36 B.n333 B.n116 585
R37 B.n332 B.n331 585
R38 B.n330 B.n117 585
R39 B.n329 B.n328 585
R40 B.n327 B.n118 585
R41 B.n326 B.n325 585
R42 B.n324 B.n119 585
R43 B.n323 B.n322 585
R44 B.n321 B.n120 585
R45 B.n320 B.n319 585
R46 B.n318 B.n121 585
R47 B.n317 B.n316 585
R48 B.n315 B.n122 585
R49 B.n314 B.n313 585
R50 B.n312 B.n123 585
R51 B.n311 B.n310 585
R52 B.n309 B.n124 585
R53 B.n308 B.n307 585
R54 B.n306 B.n125 585
R55 B.n305 B.n304 585
R56 B.n303 B.n126 585
R57 B.n302 B.n301 585
R58 B.n297 B.n127 585
R59 B.n296 B.n295 585
R60 B.n294 B.n128 585
R61 B.n293 B.n292 585
R62 B.n291 B.n129 585
R63 B.n290 B.n289 585
R64 B.n288 B.n130 585
R65 B.n287 B.n286 585
R66 B.n285 B.n131 585
R67 B.n283 B.n282 585
R68 B.n281 B.n134 585
R69 B.n280 B.n279 585
R70 B.n278 B.n135 585
R71 B.n277 B.n276 585
R72 B.n275 B.n136 585
R73 B.n274 B.n273 585
R74 B.n272 B.n137 585
R75 B.n271 B.n270 585
R76 B.n269 B.n138 585
R77 B.n268 B.n267 585
R78 B.n266 B.n139 585
R79 B.n265 B.n264 585
R80 B.n263 B.n140 585
R81 B.n262 B.n261 585
R82 B.n260 B.n141 585
R83 B.n259 B.n258 585
R84 B.n257 B.n142 585
R85 B.n256 B.n255 585
R86 B.n254 B.n143 585
R87 B.n253 B.n252 585
R88 B.n251 B.n144 585
R89 B.n250 B.n249 585
R90 B.n248 B.n145 585
R91 B.n247 B.n246 585
R92 B.n245 B.n146 585
R93 B.n244 B.n243 585
R94 B.n242 B.n147 585
R95 B.n241 B.n240 585
R96 B.n239 B.n148 585
R97 B.n238 B.n237 585
R98 B.n236 B.n149 585
R99 B.n235 B.n234 585
R100 B.n233 B.n150 585
R101 B.n232 B.n231 585
R102 B.n230 B.n151 585
R103 B.n229 B.n228 585
R104 B.n227 B.n152 585
R105 B.n226 B.n225 585
R106 B.n224 B.n153 585
R107 B.n223 B.n222 585
R108 B.n221 B.n154 585
R109 B.n220 B.n219 585
R110 B.n218 B.n155 585
R111 B.n217 B.n216 585
R112 B.n215 B.n156 585
R113 B.n214 B.n213 585
R114 B.n212 B.n157 585
R115 B.n211 B.n210 585
R116 B.n209 B.n158 585
R117 B.n208 B.n207 585
R118 B.n206 B.n159 585
R119 B.n205 B.n204 585
R120 B.n383 B.n382 585
R121 B.n384 B.n99 585
R122 B.n386 B.n385 585
R123 B.n387 B.n98 585
R124 B.n389 B.n388 585
R125 B.n390 B.n97 585
R126 B.n392 B.n391 585
R127 B.n393 B.n96 585
R128 B.n395 B.n394 585
R129 B.n396 B.n95 585
R130 B.n398 B.n397 585
R131 B.n399 B.n94 585
R132 B.n401 B.n400 585
R133 B.n402 B.n93 585
R134 B.n404 B.n403 585
R135 B.n405 B.n92 585
R136 B.n407 B.n406 585
R137 B.n408 B.n91 585
R138 B.n410 B.n409 585
R139 B.n411 B.n90 585
R140 B.n413 B.n412 585
R141 B.n414 B.n89 585
R142 B.n416 B.n415 585
R143 B.n417 B.n88 585
R144 B.n419 B.n418 585
R145 B.n420 B.n87 585
R146 B.n422 B.n421 585
R147 B.n423 B.n86 585
R148 B.n425 B.n424 585
R149 B.n426 B.n85 585
R150 B.n428 B.n427 585
R151 B.n429 B.n84 585
R152 B.n431 B.n430 585
R153 B.n432 B.n83 585
R154 B.n434 B.n433 585
R155 B.n435 B.n82 585
R156 B.n437 B.n436 585
R157 B.n438 B.n81 585
R158 B.n440 B.n439 585
R159 B.n441 B.n80 585
R160 B.n443 B.n442 585
R161 B.n444 B.n79 585
R162 B.n446 B.n445 585
R163 B.n447 B.n78 585
R164 B.n449 B.n448 585
R165 B.n450 B.n77 585
R166 B.n452 B.n451 585
R167 B.n453 B.n76 585
R168 B.n629 B.n628 585
R169 B.n627 B.n14 585
R170 B.n626 B.n625 585
R171 B.n624 B.n15 585
R172 B.n623 B.n622 585
R173 B.n621 B.n16 585
R174 B.n620 B.n619 585
R175 B.n618 B.n17 585
R176 B.n617 B.n616 585
R177 B.n615 B.n18 585
R178 B.n614 B.n613 585
R179 B.n612 B.n19 585
R180 B.n611 B.n610 585
R181 B.n609 B.n20 585
R182 B.n608 B.n607 585
R183 B.n606 B.n21 585
R184 B.n605 B.n604 585
R185 B.n603 B.n22 585
R186 B.n602 B.n601 585
R187 B.n600 B.n23 585
R188 B.n599 B.n598 585
R189 B.n597 B.n24 585
R190 B.n596 B.n595 585
R191 B.n594 B.n25 585
R192 B.n593 B.n592 585
R193 B.n591 B.n26 585
R194 B.n590 B.n589 585
R195 B.n588 B.n27 585
R196 B.n587 B.n586 585
R197 B.n585 B.n28 585
R198 B.n584 B.n583 585
R199 B.n582 B.n29 585
R200 B.n581 B.n580 585
R201 B.n579 B.n30 585
R202 B.n578 B.n577 585
R203 B.n576 B.n31 585
R204 B.n575 B.n574 585
R205 B.n573 B.n32 585
R206 B.n572 B.n571 585
R207 B.n570 B.n33 585
R208 B.n569 B.n568 585
R209 B.n567 B.n34 585
R210 B.n566 B.n565 585
R211 B.n564 B.n35 585
R212 B.n563 B.n562 585
R213 B.n561 B.n36 585
R214 B.n560 B.n559 585
R215 B.n558 B.n37 585
R216 B.n557 B.n556 585
R217 B.n555 B.n38 585
R218 B.n554 B.n553 585
R219 B.n552 B.n39 585
R220 B.n551 B.n550 585
R221 B.n549 B.n548 585
R222 B.n547 B.n43 585
R223 B.n546 B.n545 585
R224 B.n544 B.n44 585
R225 B.n543 B.n542 585
R226 B.n541 B.n45 585
R227 B.n540 B.n539 585
R228 B.n538 B.n46 585
R229 B.n537 B.n536 585
R230 B.n535 B.n47 585
R231 B.n533 B.n532 585
R232 B.n531 B.n50 585
R233 B.n530 B.n529 585
R234 B.n528 B.n51 585
R235 B.n527 B.n526 585
R236 B.n525 B.n52 585
R237 B.n524 B.n523 585
R238 B.n522 B.n53 585
R239 B.n521 B.n520 585
R240 B.n519 B.n54 585
R241 B.n518 B.n517 585
R242 B.n516 B.n55 585
R243 B.n515 B.n514 585
R244 B.n513 B.n56 585
R245 B.n512 B.n511 585
R246 B.n510 B.n57 585
R247 B.n509 B.n508 585
R248 B.n507 B.n58 585
R249 B.n506 B.n505 585
R250 B.n504 B.n59 585
R251 B.n503 B.n502 585
R252 B.n501 B.n60 585
R253 B.n500 B.n499 585
R254 B.n498 B.n61 585
R255 B.n497 B.n496 585
R256 B.n495 B.n62 585
R257 B.n494 B.n493 585
R258 B.n492 B.n63 585
R259 B.n491 B.n490 585
R260 B.n489 B.n64 585
R261 B.n488 B.n487 585
R262 B.n486 B.n65 585
R263 B.n485 B.n484 585
R264 B.n483 B.n66 585
R265 B.n482 B.n481 585
R266 B.n480 B.n67 585
R267 B.n479 B.n478 585
R268 B.n477 B.n68 585
R269 B.n476 B.n475 585
R270 B.n474 B.n69 585
R271 B.n473 B.n472 585
R272 B.n471 B.n70 585
R273 B.n470 B.n469 585
R274 B.n468 B.n71 585
R275 B.n467 B.n466 585
R276 B.n465 B.n72 585
R277 B.n464 B.n463 585
R278 B.n462 B.n73 585
R279 B.n461 B.n460 585
R280 B.n459 B.n74 585
R281 B.n458 B.n457 585
R282 B.n456 B.n75 585
R283 B.n455 B.n454 585
R284 B.n630 B.n13 585
R285 B.n632 B.n631 585
R286 B.n633 B.n12 585
R287 B.n635 B.n634 585
R288 B.n636 B.n11 585
R289 B.n638 B.n637 585
R290 B.n639 B.n10 585
R291 B.n641 B.n640 585
R292 B.n642 B.n9 585
R293 B.n644 B.n643 585
R294 B.n645 B.n8 585
R295 B.n647 B.n646 585
R296 B.n648 B.n7 585
R297 B.n650 B.n649 585
R298 B.n651 B.n6 585
R299 B.n653 B.n652 585
R300 B.n654 B.n5 585
R301 B.n656 B.n655 585
R302 B.n657 B.n4 585
R303 B.n659 B.n658 585
R304 B.n660 B.n3 585
R305 B.n662 B.n661 585
R306 B.n663 B.n0 585
R307 B.n2 B.n1 585
R308 B.n172 B.n171 585
R309 B.n173 B.n170 585
R310 B.n175 B.n174 585
R311 B.n176 B.n169 585
R312 B.n178 B.n177 585
R313 B.n179 B.n168 585
R314 B.n181 B.n180 585
R315 B.n182 B.n167 585
R316 B.n184 B.n183 585
R317 B.n185 B.n166 585
R318 B.n187 B.n186 585
R319 B.n188 B.n165 585
R320 B.n190 B.n189 585
R321 B.n191 B.n164 585
R322 B.n193 B.n192 585
R323 B.n194 B.n163 585
R324 B.n196 B.n195 585
R325 B.n197 B.n162 585
R326 B.n199 B.n198 585
R327 B.n200 B.n161 585
R328 B.n202 B.n201 585
R329 B.n203 B.n160 585
R330 B.n204 B.n203 569.379
R331 B.n382 B.n381 569.379
R332 B.n454 B.n453 569.379
R333 B.n628 B.n13 569.379
R334 B.n298 B.t10 468.411
R335 B.n48 B.t5 468.411
R336 B.n132 B.t1 468.411
R337 B.n40 B.t8 468.411
R338 B.n299 B.t11 447.853
R339 B.n49 B.t4 447.853
R340 B.n133 B.t2 447.853
R341 B.n41 B.t7 447.853
R342 B.n665 B.n664 256.663
R343 B.n664 B.n663 235.042
R344 B.n664 B.n2 235.042
R345 B.n204 B.n159 163.367
R346 B.n208 B.n159 163.367
R347 B.n209 B.n208 163.367
R348 B.n210 B.n209 163.367
R349 B.n210 B.n157 163.367
R350 B.n214 B.n157 163.367
R351 B.n215 B.n214 163.367
R352 B.n216 B.n215 163.367
R353 B.n216 B.n155 163.367
R354 B.n220 B.n155 163.367
R355 B.n221 B.n220 163.367
R356 B.n222 B.n221 163.367
R357 B.n222 B.n153 163.367
R358 B.n226 B.n153 163.367
R359 B.n227 B.n226 163.367
R360 B.n228 B.n227 163.367
R361 B.n228 B.n151 163.367
R362 B.n232 B.n151 163.367
R363 B.n233 B.n232 163.367
R364 B.n234 B.n233 163.367
R365 B.n234 B.n149 163.367
R366 B.n238 B.n149 163.367
R367 B.n239 B.n238 163.367
R368 B.n240 B.n239 163.367
R369 B.n240 B.n147 163.367
R370 B.n244 B.n147 163.367
R371 B.n245 B.n244 163.367
R372 B.n246 B.n245 163.367
R373 B.n246 B.n145 163.367
R374 B.n250 B.n145 163.367
R375 B.n251 B.n250 163.367
R376 B.n252 B.n251 163.367
R377 B.n252 B.n143 163.367
R378 B.n256 B.n143 163.367
R379 B.n257 B.n256 163.367
R380 B.n258 B.n257 163.367
R381 B.n258 B.n141 163.367
R382 B.n262 B.n141 163.367
R383 B.n263 B.n262 163.367
R384 B.n264 B.n263 163.367
R385 B.n264 B.n139 163.367
R386 B.n268 B.n139 163.367
R387 B.n269 B.n268 163.367
R388 B.n270 B.n269 163.367
R389 B.n270 B.n137 163.367
R390 B.n274 B.n137 163.367
R391 B.n275 B.n274 163.367
R392 B.n276 B.n275 163.367
R393 B.n276 B.n135 163.367
R394 B.n280 B.n135 163.367
R395 B.n281 B.n280 163.367
R396 B.n282 B.n281 163.367
R397 B.n282 B.n131 163.367
R398 B.n287 B.n131 163.367
R399 B.n288 B.n287 163.367
R400 B.n289 B.n288 163.367
R401 B.n289 B.n129 163.367
R402 B.n293 B.n129 163.367
R403 B.n294 B.n293 163.367
R404 B.n295 B.n294 163.367
R405 B.n295 B.n127 163.367
R406 B.n302 B.n127 163.367
R407 B.n303 B.n302 163.367
R408 B.n304 B.n303 163.367
R409 B.n304 B.n125 163.367
R410 B.n308 B.n125 163.367
R411 B.n309 B.n308 163.367
R412 B.n310 B.n309 163.367
R413 B.n310 B.n123 163.367
R414 B.n314 B.n123 163.367
R415 B.n315 B.n314 163.367
R416 B.n316 B.n315 163.367
R417 B.n316 B.n121 163.367
R418 B.n320 B.n121 163.367
R419 B.n321 B.n320 163.367
R420 B.n322 B.n321 163.367
R421 B.n322 B.n119 163.367
R422 B.n326 B.n119 163.367
R423 B.n327 B.n326 163.367
R424 B.n328 B.n327 163.367
R425 B.n328 B.n117 163.367
R426 B.n332 B.n117 163.367
R427 B.n333 B.n332 163.367
R428 B.n334 B.n333 163.367
R429 B.n334 B.n115 163.367
R430 B.n338 B.n115 163.367
R431 B.n339 B.n338 163.367
R432 B.n340 B.n339 163.367
R433 B.n340 B.n113 163.367
R434 B.n344 B.n113 163.367
R435 B.n345 B.n344 163.367
R436 B.n346 B.n345 163.367
R437 B.n346 B.n111 163.367
R438 B.n350 B.n111 163.367
R439 B.n351 B.n350 163.367
R440 B.n352 B.n351 163.367
R441 B.n352 B.n109 163.367
R442 B.n356 B.n109 163.367
R443 B.n357 B.n356 163.367
R444 B.n358 B.n357 163.367
R445 B.n358 B.n107 163.367
R446 B.n362 B.n107 163.367
R447 B.n363 B.n362 163.367
R448 B.n364 B.n363 163.367
R449 B.n364 B.n105 163.367
R450 B.n368 B.n105 163.367
R451 B.n369 B.n368 163.367
R452 B.n370 B.n369 163.367
R453 B.n370 B.n103 163.367
R454 B.n374 B.n103 163.367
R455 B.n375 B.n374 163.367
R456 B.n376 B.n375 163.367
R457 B.n376 B.n101 163.367
R458 B.n380 B.n101 163.367
R459 B.n381 B.n380 163.367
R460 B.n453 B.n452 163.367
R461 B.n452 B.n77 163.367
R462 B.n448 B.n77 163.367
R463 B.n448 B.n447 163.367
R464 B.n447 B.n446 163.367
R465 B.n446 B.n79 163.367
R466 B.n442 B.n79 163.367
R467 B.n442 B.n441 163.367
R468 B.n441 B.n440 163.367
R469 B.n440 B.n81 163.367
R470 B.n436 B.n81 163.367
R471 B.n436 B.n435 163.367
R472 B.n435 B.n434 163.367
R473 B.n434 B.n83 163.367
R474 B.n430 B.n83 163.367
R475 B.n430 B.n429 163.367
R476 B.n429 B.n428 163.367
R477 B.n428 B.n85 163.367
R478 B.n424 B.n85 163.367
R479 B.n424 B.n423 163.367
R480 B.n423 B.n422 163.367
R481 B.n422 B.n87 163.367
R482 B.n418 B.n87 163.367
R483 B.n418 B.n417 163.367
R484 B.n417 B.n416 163.367
R485 B.n416 B.n89 163.367
R486 B.n412 B.n89 163.367
R487 B.n412 B.n411 163.367
R488 B.n411 B.n410 163.367
R489 B.n410 B.n91 163.367
R490 B.n406 B.n91 163.367
R491 B.n406 B.n405 163.367
R492 B.n405 B.n404 163.367
R493 B.n404 B.n93 163.367
R494 B.n400 B.n93 163.367
R495 B.n400 B.n399 163.367
R496 B.n399 B.n398 163.367
R497 B.n398 B.n95 163.367
R498 B.n394 B.n95 163.367
R499 B.n394 B.n393 163.367
R500 B.n393 B.n392 163.367
R501 B.n392 B.n97 163.367
R502 B.n388 B.n97 163.367
R503 B.n388 B.n387 163.367
R504 B.n387 B.n386 163.367
R505 B.n386 B.n99 163.367
R506 B.n382 B.n99 163.367
R507 B.n628 B.n627 163.367
R508 B.n627 B.n626 163.367
R509 B.n626 B.n15 163.367
R510 B.n622 B.n15 163.367
R511 B.n622 B.n621 163.367
R512 B.n621 B.n620 163.367
R513 B.n620 B.n17 163.367
R514 B.n616 B.n17 163.367
R515 B.n616 B.n615 163.367
R516 B.n615 B.n614 163.367
R517 B.n614 B.n19 163.367
R518 B.n610 B.n19 163.367
R519 B.n610 B.n609 163.367
R520 B.n609 B.n608 163.367
R521 B.n608 B.n21 163.367
R522 B.n604 B.n21 163.367
R523 B.n604 B.n603 163.367
R524 B.n603 B.n602 163.367
R525 B.n602 B.n23 163.367
R526 B.n598 B.n23 163.367
R527 B.n598 B.n597 163.367
R528 B.n597 B.n596 163.367
R529 B.n596 B.n25 163.367
R530 B.n592 B.n25 163.367
R531 B.n592 B.n591 163.367
R532 B.n591 B.n590 163.367
R533 B.n590 B.n27 163.367
R534 B.n586 B.n27 163.367
R535 B.n586 B.n585 163.367
R536 B.n585 B.n584 163.367
R537 B.n584 B.n29 163.367
R538 B.n580 B.n29 163.367
R539 B.n580 B.n579 163.367
R540 B.n579 B.n578 163.367
R541 B.n578 B.n31 163.367
R542 B.n574 B.n31 163.367
R543 B.n574 B.n573 163.367
R544 B.n573 B.n572 163.367
R545 B.n572 B.n33 163.367
R546 B.n568 B.n33 163.367
R547 B.n568 B.n567 163.367
R548 B.n567 B.n566 163.367
R549 B.n566 B.n35 163.367
R550 B.n562 B.n35 163.367
R551 B.n562 B.n561 163.367
R552 B.n561 B.n560 163.367
R553 B.n560 B.n37 163.367
R554 B.n556 B.n37 163.367
R555 B.n556 B.n555 163.367
R556 B.n555 B.n554 163.367
R557 B.n554 B.n39 163.367
R558 B.n550 B.n39 163.367
R559 B.n550 B.n549 163.367
R560 B.n549 B.n43 163.367
R561 B.n545 B.n43 163.367
R562 B.n545 B.n544 163.367
R563 B.n544 B.n543 163.367
R564 B.n543 B.n45 163.367
R565 B.n539 B.n45 163.367
R566 B.n539 B.n538 163.367
R567 B.n538 B.n537 163.367
R568 B.n537 B.n47 163.367
R569 B.n532 B.n47 163.367
R570 B.n532 B.n531 163.367
R571 B.n531 B.n530 163.367
R572 B.n530 B.n51 163.367
R573 B.n526 B.n51 163.367
R574 B.n526 B.n525 163.367
R575 B.n525 B.n524 163.367
R576 B.n524 B.n53 163.367
R577 B.n520 B.n53 163.367
R578 B.n520 B.n519 163.367
R579 B.n519 B.n518 163.367
R580 B.n518 B.n55 163.367
R581 B.n514 B.n55 163.367
R582 B.n514 B.n513 163.367
R583 B.n513 B.n512 163.367
R584 B.n512 B.n57 163.367
R585 B.n508 B.n57 163.367
R586 B.n508 B.n507 163.367
R587 B.n507 B.n506 163.367
R588 B.n506 B.n59 163.367
R589 B.n502 B.n59 163.367
R590 B.n502 B.n501 163.367
R591 B.n501 B.n500 163.367
R592 B.n500 B.n61 163.367
R593 B.n496 B.n61 163.367
R594 B.n496 B.n495 163.367
R595 B.n495 B.n494 163.367
R596 B.n494 B.n63 163.367
R597 B.n490 B.n63 163.367
R598 B.n490 B.n489 163.367
R599 B.n489 B.n488 163.367
R600 B.n488 B.n65 163.367
R601 B.n484 B.n65 163.367
R602 B.n484 B.n483 163.367
R603 B.n483 B.n482 163.367
R604 B.n482 B.n67 163.367
R605 B.n478 B.n67 163.367
R606 B.n478 B.n477 163.367
R607 B.n477 B.n476 163.367
R608 B.n476 B.n69 163.367
R609 B.n472 B.n69 163.367
R610 B.n472 B.n471 163.367
R611 B.n471 B.n470 163.367
R612 B.n470 B.n71 163.367
R613 B.n466 B.n71 163.367
R614 B.n466 B.n465 163.367
R615 B.n465 B.n464 163.367
R616 B.n464 B.n73 163.367
R617 B.n460 B.n73 163.367
R618 B.n460 B.n459 163.367
R619 B.n459 B.n458 163.367
R620 B.n458 B.n75 163.367
R621 B.n454 B.n75 163.367
R622 B.n632 B.n13 163.367
R623 B.n633 B.n632 163.367
R624 B.n634 B.n633 163.367
R625 B.n634 B.n11 163.367
R626 B.n638 B.n11 163.367
R627 B.n639 B.n638 163.367
R628 B.n640 B.n639 163.367
R629 B.n640 B.n9 163.367
R630 B.n644 B.n9 163.367
R631 B.n645 B.n644 163.367
R632 B.n646 B.n645 163.367
R633 B.n646 B.n7 163.367
R634 B.n650 B.n7 163.367
R635 B.n651 B.n650 163.367
R636 B.n652 B.n651 163.367
R637 B.n652 B.n5 163.367
R638 B.n656 B.n5 163.367
R639 B.n657 B.n656 163.367
R640 B.n658 B.n657 163.367
R641 B.n658 B.n3 163.367
R642 B.n662 B.n3 163.367
R643 B.n663 B.n662 163.367
R644 B.n172 B.n2 163.367
R645 B.n173 B.n172 163.367
R646 B.n174 B.n173 163.367
R647 B.n174 B.n169 163.367
R648 B.n178 B.n169 163.367
R649 B.n179 B.n178 163.367
R650 B.n180 B.n179 163.367
R651 B.n180 B.n167 163.367
R652 B.n184 B.n167 163.367
R653 B.n185 B.n184 163.367
R654 B.n186 B.n185 163.367
R655 B.n186 B.n165 163.367
R656 B.n190 B.n165 163.367
R657 B.n191 B.n190 163.367
R658 B.n192 B.n191 163.367
R659 B.n192 B.n163 163.367
R660 B.n196 B.n163 163.367
R661 B.n197 B.n196 163.367
R662 B.n198 B.n197 163.367
R663 B.n198 B.n161 163.367
R664 B.n202 B.n161 163.367
R665 B.n203 B.n202 163.367
R666 B.n284 B.n133 59.5399
R667 B.n300 B.n299 59.5399
R668 B.n534 B.n49 59.5399
R669 B.n42 B.n41 59.5399
R670 B.n630 B.n629 36.9956
R671 B.n455 B.n76 36.9956
R672 B.n383 B.n100 36.9956
R673 B.n205 B.n160 36.9956
R674 B.n133 B.n132 20.5581
R675 B.n299 B.n298 20.5581
R676 B.n49 B.n48 20.5581
R677 B.n41 B.n40 20.5581
R678 B B.n665 18.0485
R679 B.n631 B.n630 10.6151
R680 B.n631 B.n12 10.6151
R681 B.n635 B.n12 10.6151
R682 B.n636 B.n635 10.6151
R683 B.n637 B.n636 10.6151
R684 B.n637 B.n10 10.6151
R685 B.n641 B.n10 10.6151
R686 B.n642 B.n641 10.6151
R687 B.n643 B.n642 10.6151
R688 B.n643 B.n8 10.6151
R689 B.n647 B.n8 10.6151
R690 B.n648 B.n647 10.6151
R691 B.n649 B.n648 10.6151
R692 B.n649 B.n6 10.6151
R693 B.n653 B.n6 10.6151
R694 B.n654 B.n653 10.6151
R695 B.n655 B.n654 10.6151
R696 B.n655 B.n4 10.6151
R697 B.n659 B.n4 10.6151
R698 B.n660 B.n659 10.6151
R699 B.n661 B.n660 10.6151
R700 B.n661 B.n0 10.6151
R701 B.n629 B.n14 10.6151
R702 B.n625 B.n14 10.6151
R703 B.n625 B.n624 10.6151
R704 B.n624 B.n623 10.6151
R705 B.n623 B.n16 10.6151
R706 B.n619 B.n16 10.6151
R707 B.n619 B.n618 10.6151
R708 B.n618 B.n617 10.6151
R709 B.n617 B.n18 10.6151
R710 B.n613 B.n18 10.6151
R711 B.n613 B.n612 10.6151
R712 B.n612 B.n611 10.6151
R713 B.n611 B.n20 10.6151
R714 B.n607 B.n20 10.6151
R715 B.n607 B.n606 10.6151
R716 B.n606 B.n605 10.6151
R717 B.n605 B.n22 10.6151
R718 B.n601 B.n22 10.6151
R719 B.n601 B.n600 10.6151
R720 B.n600 B.n599 10.6151
R721 B.n599 B.n24 10.6151
R722 B.n595 B.n24 10.6151
R723 B.n595 B.n594 10.6151
R724 B.n594 B.n593 10.6151
R725 B.n593 B.n26 10.6151
R726 B.n589 B.n26 10.6151
R727 B.n589 B.n588 10.6151
R728 B.n588 B.n587 10.6151
R729 B.n587 B.n28 10.6151
R730 B.n583 B.n28 10.6151
R731 B.n583 B.n582 10.6151
R732 B.n582 B.n581 10.6151
R733 B.n581 B.n30 10.6151
R734 B.n577 B.n30 10.6151
R735 B.n577 B.n576 10.6151
R736 B.n576 B.n575 10.6151
R737 B.n575 B.n32 10.6151
R738 B.n571 B.n32 10.6151
R739 B.n571 B.n570 10.6151
R740 B.n570 B.n569 10.6151
R741 B.n569 B.n34 10.6151
R742 B.n565 B.n34 10.6151
R743 B.n565 B.n564 10.6151
R744 B.n564 B.n563 10.6151
R745 B.n563 B.n36 10.6151
R746 B.n559 B.n36 10.6151
R747 B.n559 B.n558 10.6151
R748 B.n558 B.n557 10.6151
R749 B.n557 B.n38 10.6151
R750 B.n553 B.n38 10.6151
R751 B.n553 B.n552 10.6151
R752 B.n552 B.n551 10.6151
R753 B.n548 B.n547 10.6151
R754 B.n547 B.n546 10.6151
R755 B.n546 B.n44 10.6151
R756 B.n542 B.n44 10.6151
R757 B.n542 B.n541 10.6151
R758 B.n541 B.n540 10.6151
R759 B.n540 B.n46 10.6151
R760 B.n536 B.n46 10.6151
R761 B.n536 B.n535 10.6151
R762 B.n533 B.n50 10.6151
R763 B.n529 B.n50 10.6151
R764 B.n529 B.n528 10.6151
R765 B.n528 B.n527 10.6151
R766 B.n527 B.n52 10.6151
R767 B.n523 B.n52 10.6151
R768 B.n523 B.n522 10.6151
R769 B.n522 B.n521 10.6151
R770 B.n521 B.n54 10.6151
R771 B.n517 B.n54 10.6151
R772 B.n517 B.n516 10.6151
R773 B.n516 B.n515 10.6151
R774 B.n515 B.n56 10.6151
R775 B.n511 B.n56 10.6151
R776 B.n511 B.n510 10.6151
R777 B.n510 B.n509 10.6151
R778 B.n509 B.n58 10.6151
R779 B.n505 B.n58 10.6151
R780 B.n505 B.n504 10.6151
R781 B.n504 B.n503 10.6151
R782 B.n503 B.n60 10.6151
R783 B.n499 B.n60 10.6151
R784 B.n499 B.n498 10.6151
R785 B.n498 B.n497 10.6151
R786 B.n497 B.n62 10.6151
R787 B.n493 B.n62 10.6151
R788 B.n493 B.n492 10.6151
R789 B.n492 B.n491 10.6151
R790 B.n491 B.n64 10.6151
R791 B.n487 B.n64 10.6151
R792 B.n487 B.n486 10.6151
R793 B.n486 B.n485 10.6151
R794 B.n485 B.n66 10.6151
R795 B.n481 B.n66 10.6151
R796 B.n481 B.n480 10.6151
R797 B.n480 B.n479 10.6151
R798 B.n479 B.n68 10.6151
R799 B.n475 B.n68 10.6151
R800 B.n475 B.n474 10.6151
R801 B.n474 B.n473 10.6151
R802 B.n473 B.n70 10.6151
R803 B.n469 B.n70 10.6151
R804 B.n469 B.n468 10.6151
R805 B.n468 B.n467 10.6151
R806 B.n467 B.n72 10.6151
R807 B.n463 B.n72 10.6151
R808 B.n463 B.n462 10.6151
R809 B.n462 B.n461 10.6151
R810 B.n461 B.n74 10.6151
R811 B.n457 B.n74 10.6151
R812 B.n457 B.n456 10.6151
R813 B.n456 B.n455 10.6151
R814 B.n451 B.n76 10.6151
R815 B.n451 B.n450 10.6151
R816 B.n450 B.n449 10.6151
R817 B.n449 B.n78 10.6151
R818 B.n445 B.n78 10.6151
R819 B.n445 B.n444 10.6151
R820 B.n444 B.n443 10.6151
R821 B.n443 B.n80 10.6151
R822 B.n439 B.n80 10.6151
R823 B.n439 B.n438 10.6151
R824 B.n438 B.n437 10.6151
R825 B.n437 B.n82 10.6151
R826 B.n433 B.n82 10.6151
R827 B.n433 B.n432 10.6151
R828 B.n432 B.n431 10.6151
R829 B.n431 B.n84 10.6151
R830 B.n427 B.n84 10.6151
R831 B.n427 B.n426 10.6151
R832 B.n426 B.n425 10.6151
R833 B.n425 B.n86 10.6151
R834 B.n421 B.n86 10.6151
R835 B.n421 B.n420 10.6151
R836 B.n420 B.n419 10.6151
R837 B.n419 B.n88 10.6151
R838 B.n415 B.n88 10.6151
R839 B.n415 B.n414 10.6151
R840 B.n414 B.n413 10.6151
R841 B.n413 B.n90 10.6151
R842 B.n409 B.n90 10.6151
R843 B.n409 B.n408 10.6151
R844 B.n408 B.n407 10.6151
R845 B.n407 B.n92 10.6151
R846 B.n403 B.n92 10.6151
R847 B.n403 B.n402 10.6151
R848 B.n402 B.n401 10.6151
R849 B.n401 B.n94 10.6151
R850 B.n397 B.n94 10.6151
R851 B.n397 B.n396 10.6151
R852 B.n396 B.n395 10.6151
R853 B.n395 B.n96 10.6151
R854 B.n391 B.n96 10.6151
R855 B.n391 B.n390 10.6151
R856 B.n390 B.n389 10.6151
R857 B.n389 B.n98 10.6151
R858 B.n385 B.n98 10.6151
R859 B.n385 B.n384 10.6151
R860 B.n384 B.n383 10.6151
R861 B.n171 B.n1 10.6151
R862 B.n171 B.n170 10.6151
R863 B.n175 B.n170 10.6151
R864 B.n176 B.n175 10.6151
R865 B.n177 B.n176 10.6151
R866 B.n177 B.n168 10.6151
R867 B.n181 B.n168 10.6151
R868 B.n182 B.n181 10.6151
R869 B.n183 B.n182 10.6151
R870 B.n183 B.n166 10.6151
R871 B.n187 B.n166 10.6151
R872 B.n188 B.n187 10.6151
R873 B.n189 B.n188 10.6151
R874 B.n189 B.n164 10.6151
R875 B.n193 B.n164 10.6151
R876 B.n194 B.n193 10.6151
R877 B.n195 B.n194 10.6151
R878 B.n195 B.n162 10.6151
R879 B.n199 B.n162 10.6151
R880 B.n200 B.n199 10.6151
R881 B.n201 B.n200 10.6151
R882 B.n201 B.n160 10.6151
R883 B.n206 B.n205 10.6151
R884 B.n207 B.n206 10.6151
R885 B.n207 B.n158 10.6151
R886 B.n211 B.n158 10.6151
R887 B.n212 B.n211 10.6151
R888 B.n213 B.n212 10.6151
R889 B.n213 B.n156 10.6151
R890 B.n217 B.n156 10.6151
R891 B.n218 B.n217 10.6151
R892 B.n219 B.n218 10.6151
R893 B.n219 B.n154 10.6151
R894 B.n223 B.n154 10.6151
R895 B.n224 B.n223 10.6151
R896 B.n225 B.n224 10.6151
R897 B.n225 B.n152 10.6151
R898 B.n229 B.n152 10.6151
R899 B.n230 B.n229 10.6151
R900 B.n231 B.n230 10.6151
R901 B.n231 B.n150 10.6151
R902 B.n235 B.n150 10.6151
R903 B.n236 B.n235 10.6151
R904 B.n237 B.n236 10.6151
R905 B.n237 B.n148 10.6151
R906 B.n241 B.n148 10.6151
R907 B.n242 B.n241 10.6151
R908 B.n243 B.n242 10.6151
R909 B.n243 B.n146 10.6151
R910 B.n247 B.n146 10.6151
R911 B.n248 B.n247 10.6151
R912 B.n249 B.n248 10.6151
R913 B.n249 B.n144 10.6151
R914 B.n253 B.n144 10.6151
R915 B.n254 B.n253 10.6151
R916 B.n255 B.n254 10.6151
R917 B.n255 B.n142 10.6151
R918 B.n259 B.n142 10.6151
R919 B.n260 B.n259 10.6151
R920 B.n261 B.n260 10.6151
R921 B.n261 B.n140 10.6151
R922 B.n265 B.n140 10.6151
R923 B.n266 B.n265 10.6151
R924 B.n267 B.n266 10.6151
R925 B.n267 B.n138 10.6151
R926 B.n271 B.n138 10.6151
R927 B.n272 B.n271 10.6151
R928 B.n273 B.n272 10.6151
R929 B.n273 B.n136 10.6151
R930 B.n277 B.n136 10.6151
R931 B.n278 B.n277 10.6151
R932 B.n279 B.n278 10.6151
R933 B.n279 B.n134 10.6151
R934 B.n283 B.n134 10.6151
R935 B.n286 B.n285 10.6151
R936 B.n286 B.n130 10.6151
R937 B.n290 B.n130 10.6151
R938 B.n291 B.n290 10.6151
R939 B.n292 B.n291 10.6151
R940 B.n292 B.n128 10.6151
R941 B.n296 B.n128 10.6151
R942 B.n297 B.n296 10.6151
R943 B.n301 B.n297 10.6151
R944 B.n305 B.n126 10.6151
R945 B.n306 B.n305 10.6151
R946 B.n307 B.n306 10.6151
R947 B.n307 B.n124 10.6151
R948 B.n311 B.n124 10.6151
R949 B.n312 B.n311 10.6151
R950 B.n313 B.n312 10.6151
R951 B.n313 B.n122 10.6151
R952 B.n317 B.n122 10.6151
R953 B.n318 B.n317 10.6151
R954 B.n319 B.n318 10.6151
R955 B.n319 B.n120 10.6151
R956 B.n323 B.n120 10.6151
R957 B.n324 B.n323 10.6151
R958 B.n325 B.n324 10.6151
R959 B.n325 B.n118 10.6151
R960 B.n329 B.n118 10.6151
R961 B.n330 B.n329 10.6151
R962 B.n331 B.n330 10.6151
R963 B.n331 B.n116 10.6151
R964 B.n335 B.n116 10.6151
R965 B.n336 B.n335 10.6151
R966 B.n337 B.n336 10.6151
R967 B.n337 B.n114 10.6151
R968 B.n341 B.n114 10.6151
R969 B.n342 B.n341 10.6151
R970 B.n343 B.n342 10.6151
R971 B.n343 B.n112 10.6151
R972 B.n347 B.n112 10.6151
R973 B.n348 B.n347 10.6151
R974 B.n349 B.n348 10.6151
R975 B.n349 B.n110 10.6151
R976 B.n353 B.n110 10.6151
R977 B.n354 B.n353 10.6151
R978 B.n355 B.n354 10.6151
R979 B.n355 B.n108 10.6151
R980 B.n359 B.n108 10.6151
R981 B.n360 B.n359 10.6151
R982 B.n361 B.n360 10.6151
R983 B.n361 B.n106 10.6151
R984 B.n365 B.n106 10.6151
R985 B.n366 B.n365 10.6151
R986 B.n367 B.n366 10.6151
R987 B.n367 B.n104 10.6151
R988 B.n371 B.n104 10.6151
R989 B.n372 B.n371 10.6151
R990 B.n373 B.n372 10.6151
R991 B.n373 B.n102 10.6151
R992 B.n377 B.n102 10.6151
R993 B.n378 B.n377 10.6151
R994 B.n379 B.n378 10.6151
R995 B.n379 B.n100 10.6151
R996 B.n551 B.n42 9.36635
R997 B.n534 B.n533 9.36635
R998 B.n284 B.n283 9.36635
R999 B.n300 B.n126 9.36635
R1000 B.n665 B.n0 8.11757
R1001 B.n665 B.n1 8.11757
R1002 B.n548 B.n42 1.24928
R1003 B.n535 B.n534 1.24928
R1004 B.n285 B.n284 1.24928
R1005 B.n301 B.n300 1.24928
R1006 VP.n6 VP.t0 605.996
R1007 VP.n14 VP.t4 582.692
R1008 VP.n16 VP.t3 582.692
R1009 VP.n20 VP.t5 582.692
R1010 VP.n22 VP.t6 582.692
R1011 VP.n11 VP.t7 582.692
R1012 VP.n9 VP.t1 582.692
R1013 VP.n5 VP.t2 582.692
R1014 VP.n23 VP.n22 161.3
R1015 VP.n8 VP.n7 161.3
R1016 VP.n9 VP.n4 161.3
R1017 VP.n10 VP.n3 161.3
R1018 VP.n12 VP.n11 161.3
R1019 VP.n21 VP.n0 161.3
R1020 VP.n20 VP.n19 161.3
R1021 VP.n18 VP.n1 161.3
R1022 VP.n17 VP.n16 161.3
R1023 VP.n15 VP.n2 161.3
R1024 VP.n14 VP.n13 161.3
R1025 VP.n13 VP.n12 45.2202
R1026 VP.n7 VP.n6 44.8907
R1027 VP.n15 VP.n14 32.8641
R1028 VP.n22 VP.n21 32.8641
R1029 VP.n11 VP.n10 32.8641
R1030 VP.n16 VP.n1 24.1005
R1031 VP.n20 VP.n1 24.1005
R1032 VP.n8 VP.n5 24.1005
R1033 VP.n9 VP.n8 24.1005
R1034 VP.n6 VP.n5 18.4104
R1035 VP.n16 VP.n15 15.3369
R1036 VP.n21 VP.n20 15.3369
R1037 VP.n10 VP.n9 15.3369
R1038 VP.n7 VP.n4 0.189894
R1039 VP.n4 VP.n3 0.189894
R1040 VP.n12 VP.n3 0.189894
R1041 VP.n13 VP.n2 0.189894
R1042 VP.n17 VP.n2 0.189894
R1043 VP.n18 VP.n17 0.189894
R1044 VP.n19 VP.n18 0.189894
R1045 VP.n19 VP.n0 0.189894
R1046 VP.n23 VP.n0 0.189894
R1047 VP VP.n23 0.0516364
R1048 VDD1 VDD1.n0 69.1536
R1049 VDD1.n3 VDD1.n2 69.0399
R1050 VDD1.n3 VDD1.n1 69.0399
R1051 VDD1.n5 VDD1.n4 68.6383
R1052 VDD1.n5 VDD1.n3 42.2207
R1053 VDD1.n4 VDD1.t0 2.02953
R1054 VDD1.n4 VDD1.t6 2.02953
R1055 VDD1.n0 VDD1.t1 2.02953
R1056 VDD1.n0 VDD1.t2 2.02953
R1057 VDD1.n2 VDD1.t3 2.02953
R1058 VDD1.n2 VDD1.t7 2.02953
R1059 VDD1.n1 VDD1.t4 2.02953
R1060 VDD1.n1 VDD1.t5 2.02953
R1061 VDD1 VDD1.n5 0.399207
R1062 VTAIL.n722 VTAIL.n638 756.745
R1063 VTAIL.n86 VTAIL.n2 756.745
R1064 VTAIL.n176 VTAIL.n92 756.745
R1065 VTAIL.n268 VTAIL.n184 756.745
R1066 VTAIL.n632 VTAIL.n548 756.745
R1067 VTAIL.n540 VTAIL.n456 756.745
R1068 VTAIL.n450 VTAIL.n366 756.745
R1069 VTAIL.n358 VTAIL.n274 756.745
R1070 VTAIL.n666 VTAIL.n665 585
R1071 VTAIL.n671 VTAIL.n670 585
R1072 VTAIL.n673 VTAIL.n672 585
R1073 VTAIL.n662 VTAIL.n661 585
R1074 VTAIL.n679 VTAIL.n678 585
R1075 VTAIL.n681 VTAIL.n680 585
R1076 VTAIL.n658 VTAIL.n657 585
R1077 VTAIL.n687 VTAIL.n686 585
R1078 VTAIL.n689 VTAIL.n688 585
R1079 VTAIL.n654 VTAIL.n653 585
R1080 VTAIL.n695 VTAIL.n694 585
R1081 VTAIL.n697 VTAIL.n696 585
R1082 VTAIL.n650 VTAIL.n649 585
R1083 VTAIL.n703 VTAIL.n702 585
R1084 VTAIL.n705 VTAIL.n704 585
R1085 VTAIL.n646 VTAIL.n645 585
R1086 VTAIL.n712 VTAIL.n711 585
R1087 VTAIL.n713 VTAIL.n644 585
R1088 VTAIL.n715 VTAIL.n714 585
R1089 VTAIL.n642 VTAIL.n641 585
R1090 VTAIL.n721 VTAIL.n720 585
R1091 VTAIL.n723 VTAIL.n722 585
R1092 VTAIL.n30 VTAIL.n29 585
R1093 VTAIL.n35 VTAIL.n34 585
R1094 VTAIL.n37 VTAIL.n36 585
R1095 VTAIL.n26 VTAIL.n25 585
R1096 VTAIL.n43 VTAIL.n42 585
R1097 VTAIL.n45 VTAIL.n44 585
R1098 VTAIL.n22 VTAIL.n21 585
R1099 VTAIL.n51 VTAIL.n50 585
R1100 VTAIL.n53 VTAIL.n52 585
R1101 VTAIL.n18 VTAIL.n17 585
R1102 VTAIL.n59 VTAIL.n58 585
R1103 VTAIL.n61 VTAIL.n60 585
R1104 VTAIL.n14 VTAIL.n13 585
R1105 VTAIL.n67 VTAIL.n66 585
R1106 VTAIL.n69 VTAIL.n68 585
R1107 VTAIL.n10 VTAIL.n9 585
R1108 VTAIL.n76 VTAIL.n75 585
R1109 VTAIL.n77 VTAIL.n8 585
R1110 VTAIL.n79 VTAIL.n78 585
R1111 VTAIL.n6 VTAIL.n5 585
R1112 VTAIL.n85 VTAIL.n84 585
R1113 VTAIL.n87 VTAIL.n86 585
R1114 VTAIL.n120 VTAIL.n119 585
R1115 VTAIL.n125 VTAIL.n124 585
R1116 VTAIL.n127 VTAIL.n126 585
R1117 VTAIL.n116 VTAIL.n115 585
R1118 VTAIL.n133 VTAIL.n132 585
R1119 VTAIL.n135 VTAIL.n134 585
R1120 VTAIL.n112 VTAIL.n111 585
R1121 VTAIL.n141 VTAIL.n140 585
R1122 VTAIL.n143 VTAIL.n142 585
R1123 VTAIL.n108 VTAIL.n107 585
R1124 VTAIL.n149 VTAIL.n148 585
R1125 VTAIL.n151 VTAIL.n150 585
R1126 VTAIL.n104 VTAIL.n103 585
R1127 VTAIL.n157 VTAIL.n156 585
R1128 VTAIL.n159 VTAIL.n158 585
R1129 VTAIL.n100 VTAIL.n99 585
R1130 VTAIL.n166 VTAIL.n165 585
R1131 VTAIL.n167 VTAIL.n98 585
R1132 VTAIL.n169 VTAIL.n168 585
R1133 VTAIL.n96 VTAIL.n95 585
R1134 VTAIL.n175 VTAIL.n174 585
R1135 VTAIL.n177 VTAIL.n176 585
R1136 VTAIL.n212 VTAIL.n211 585
R1137 VTAIL.n217 VTAIL.n216 585
R1138 VTAIL.n219 VTAIL.n218 585
R1139 VTAIL.n208 VTAIL.n207 585
R1140 VTAIL.n225 VTAIL.n224 585
R1141 VTAIL.n227 VTAIL.n226 585
R1142 VTAIL.n204 VTAIL.n203 585
R1143 VTAIL.n233 VTAIL.n232 585
R1144 VTAIL.n235 VTAIL.n234 585
R1145 VTAIL.n200 VTAIL.n199 585
R1146 VTAIL.n241 VTAIL.n240 585
R1147 VTAIL.n243 VTAIL.n242 585
R1148 VTAIL.n196 VTAIL.n195 585
R1149 VTAIL.n249 VTAIL.n248 585
R1150 VTAIL.n251 VTAIL.n250 585
R1151 VTAIL.n192 VTAIL.n191 585
R1152 VTAIL.n258 VTAIL.n257 585
R1153 VTAIL.n259 VTAIL.n190 585
R1154 VTAIL.n261 VTAIL.n260 585
R1155 VTAIL.n188 VTAIL.n187 585
R1156 VTAIL.n267 VTAIL.n266 585
R1157 VTAIL.n269 VTAIL.n268 585
R1158 VTAIL.n633 VTAIL.n632 585
R1159 VTAIL.n631 VTAIL.n630 585
R1160 VTAIL.n552 VTAIL.n551 585
R1161 VTAIL.n625 VTAIL.n624 585
R1162 VTAIL.n623 VTAIL.n554 585
R1163 VTAIL.n622 VTAIL.n621 585
R1164 VTAIL.n557 VTAIL.n555 585
R1165 VTAIL.n616 VTAIL.n615 585
R1166 VTAIL.n614 VTAIL.n613 585
R1167 VTAIL.n561 VTAIL.n560 585
R1168 VTAIL.n608 VTAIL.n607 585
R1169 VTAIL.n606 VTAIL.n605 585
R1170 VTAIL.n565 VTAIL.n564 585
R1171 VTAIL.n600 VTAIL.n599 585
R1172 VTAIL.n598 VTAIL.n597 585
R1173 VTAIL.n569 VTAIL.n568 585
R1174 VTAIL.n592 VTAIL.n591 585
R1175 VTAIL.n590 VTAIL.n589 585
R1176 VTAIL.n573 VTAIL.n572 585
R1177 VTAIL.n584 VTAIL.n583 585
R1178 VTAIL.n582 VTAIL.n581 585
R1179 VTAIL.n577 VTAIL.n576 585
R1180 VTAIL.n541 VTAIL.n540 585
R1181 VTAIL.n539 VTAIL.n538 585
R1182 VTAIL.n460 VTAIL.n459 585
R1183 VTAIL.n533 VTAIL.n532 585
R1184 VTAIL.n531 VTAIL.n462 585
R1185 VTAIL.n530 VTAIL.n529 585
R1186 VTAIL.n465 VTAIL.n463 585
R1187 VTAIL.n524 VTAIL.n523 585
R1188 VTAIL.n522 VTAIL.n521 585
R1189 VTAIL.n469 VTAIL.n468 585
R1190 VTAIL.n516 VTAIL.n515 585
R1191 VTAIL.n514 VTAIL.n513 585
R1192 VTAIL.n473 VTAIL.n472 585
R1193 VTAIL.n508 VTAIL.n507 585
R1194 VTAIL.n506 VTAIL.n505 585
R1195 VTAIL.n477 VTAIL.n476 585
R1196 VTAIL.n500 VTAIL.n499 585
R1197 VTAIL.n498 VTAIL.n497 585
R1198 VTAIL.n481 VTAIL.n480 585
R1199 VTAIL.n492 VTAIL.n491 585
R1200 VTAIL.n490 VTAIL.n489 585
R1201 VTAIL.n485 VTAIL.n484 585
R1202 VTAIL.n451 VTAIL.n450 585
R1203 VTAIL.n449 VTAIL.n448 585
R1204 VTAIL.n370 VTAIL.n369 585
R1205 VTAIL.n443 VTAIL.n442 585
R1206 VTAIL.n441 VTAIL.n372 585
R1207 VTAIL.n440 VTAIL.n439 585
R1208 VTAIL.n375 VTAIL.n373 585
R1209 VTAIL.n434 VTAIL.n433 585
R1210 VTAIL.n432 VTAIL.n431 585
R1211 VTAIL.n379 VTAIL.n378 585
R1212 VTAIL.n426 VTAIL.n425 585
R1213 VTAIL.n424 VTAIL.n423 585
R1214 VTAIL.n383 VTAIL.n382 585
R1215 VTAIL.n418 VTAIL.n417 585
R1216 VTAIL.n416 VTAIL.n415 585
R1217 VTAIL.n387 VTAIL.n386 585
R1218 VTAIL.n410 VTAIL.n409 585
R1219 VTAIL.n408 VTAIL.n407 585
R1220 VTAIL.n391 VTAIL.n390 585
R1221 VTAIL.n402 VTAIL.n401 585
R1222 VTAIL.n400 VTAIL.n399 585
R1223 VTAIL.n395 VTAIL.n394 585
R1224 VTAIL.n359 VTAIL.n358 585
R1225 VTAIL.n357 VTAIL.n356 585
R1226 VTAIL.n278 VTAIL.n277 585
R1227 VTAIL.n351 VTAIL.n350 585
R1228 VTAIL.n349 VTAIL.n280 585
R1229 VTAIL.n348 VTAIL.n347 585
R1230 VTAIL.n283 VTAIL.n281 585
R1231 VTAIL.n342 VTAIL.n341 585
R1232 VTAIL.n340 VTAIL.n339 585
R1233 VTAIL.n287 VTAIL.n286 585
R1234 VTAIL.n334 VTAIL.n333 585
R1235 VTAIL.n332 VTAIL.n331 585
R1236 VTAIL.n291 VTAIL.n290 585
R1237 VTAIL.n326 VTAIL.n325 585
R1238 VTAIL.n324 VTAIL.n323 585
R1239 VTAIL.n295 VTAIL.n294 585
R1240 VTAIL.n318 VTAIL.n317 585
R1241 VTAIL.n316 VTAIL.n315 585
R1242 VTAIL.n299 VTAIL.n298 585
R1243 VTAIL.n310 VTAIL.n309 585
R1244 VTAIL.n308 VTAIL.n307 585
R1245 VTAIL.n303 VTAIL.n302 585
R1246 VTAIL.n667 VTAIL.t5 327.466
R1247 VTAIL.n31 VTAIL.t4 327.466
R1248 VTAIL.n121 VTAIL.t8 327.466
R1249 VTAIL.n213 VTAIL.t10 327.466
R1250 VTAIL.n578 VTAIL.t7 327.466
R1251 VTAIL.n486 VTAIL.t14 327.466
R1252 VTAIL.n396 VTAIL.t0 327.466
R1253 VTAIL.n304 VTAIL.t15 327.466
R1254 VTAIL.n671 VTAIL.n665 171.744
R1255 VTAIL.n672 VTAIL.n671 171.744
R1256 VTAIL.n672 VTAIL.n661 171.744
R1257 VTAIL.n679 VTAIL.n661 171.744
R1258 VTAIL.n680 VTAIL.n679 171.744
R1259 VTAIL.n680 VTAIL.n657 171.744
R1260 VTAIL.n687 VTAIL.n657 171.744
R1261 VTAIL.n688 VTAIL.n687 171.744
R1262 VTAIL.n688 VTAIL.n653 171.744
R1263 VTAIL.n695 VTAIL.n653 171.744
R1264 VTAIL.n696 VTAIL.n695 171.744
R1265 VTAIL.n696 VTAIL.n649 171.744
R1266 VTAIL.n703 VTAIL.n649 171.744
R1267 VTAIL.n704 VTAIL.n703 171.744
R1268 VTAIL.n704 VTAIL.n645 171.744
R1269 VTAIL.n712 VTAIL.n645 171.744
R1270 VTAIL.n713 VTAIL.n712 171.744
R1271 VTAIL.n714 VTAIL.n713 171.744
R1272 VTAIL.n714 VTAIL.n641 171.744
R1273 VTAIL.n721 VTAIL.n641 171.744
R1274 VTAIL.n722 VTAIL.n721 171.744
R1275 VTAIL.n35 VTAIL.n29 171.744
R1276 VTAIL.n36 VTAIL.n35 171.744
R1277 VTAIL.n36 VTAIL.n25 171.744
R1278 VTAIL.n43 VTAIL.n25 171.744
R1279 VTAIL.n44 VTAIL.n43 171.744
R1280 VTAIL.n44 VTAIL.n21 171.744
R1281 VTAIL.n51 VTAIL.n21 171.744
R1282 VTAIL.n52 VTAIL.n51 171.744
R1283 VTAIL.n52 VTAIL.n17 171.744
R1284 VTAIL.n59 VTAIL.n17 171.744
R1285 VTAIL.n60 VTAIL.n59 171.744
R1286 VTAIL.n60 VTAIL.n13 171.744
R1287 VTAIL.n67 VTAIL.n13 171.744
R1288 VTAIL.n68 VTAIL.n67 171.744
R1289 VTAIL.n68 VTAIL.n9 171.744
R1290 VTAIL.n76 VTAIL.n9 171.744
R1291 VTAIL.n77 VTAIL.n76 171.744
R1292 VTAIL.n78 VTAIL.n77 171.744
R1293 VTAIL.n78 VTAIL.n5 171.744
R1294 VTAIL.n85 VTAIL.n5 171.744
R1295 VTAIL.n86 VTAIL.n85 171.744
R1296 VTAIL.n125 VTAIL.n119 171.744
R1297 VTAIL.n126 VTAIL.n125 171.744
R1298 VTAIL.n126 VTAIL.n115 171.744
R1299 VTAIL.n133 VTAIL.n115 171.744
R1300 VTAIL.n134 VTAIL.n133 171.744
R1301 VTAIL.n134 VTAIL.n111 171.744
R1302 VTAIL.n141 VTAIL.n111 171.744
R1303 VTAIL.n142 VTAIL.n141 171.744
R1304 VTAIL.n142 VTAIL.n107 171.744
R1305 VTAIL.n149 VTAIL.n107 171.744
R1306 VTAIL.n150 VTAIL.n149 171.744
R1307 VTAIL.n150 VTAIL.n103 171.744
R1308 VTAIL.n157 VTAIL.n103 171.744
R1309 VTAIL.n158 VTAIL.n157 171.744
R1310 VTAIL.n158 VTAIL.n99 171.744
R1311 VTAIL.n166 VTAIL.n99 171.744
R1312 VTAIL.n167 VTAIL.n166 171.744
R1313 VTAIL.n168 VTAIL.n167 171.744
R1314 VTAIL.n168 VTAIL.n95 171.744
R1315 VTAIL.n175 VTAIL.n95 171.744
R1316 VTAIL.n176 VTAIL.n175 171.744
R1317 VTAIL.n217 VTAIL.n211 171.744
R1318 VTAIL.n218 VTAIL.n217 171.744
R1319 VTAIL.n218 VTAIL.n207 171.744
R1320 VTAIL.n225 VTAIL.n207 171.744
R1321 VTAIL.n226 VTAIL.n225 171.744
R1322 VTAIL.n226 VTAIL.n203 171.744
R1323 VTAIL.n233 VTAIL.n203 171.744
R1324 VTAIL.n234 VTAIL.n233 171.744
R1325 VTAIL.n234 VTAIL.n199 171.744
R1326 VTAIL.n241 VTAIL.n199 171.744
R1327 VTAIL.n242 VTAIL.n241 171.744
R1328 VTAIL.n242 VTAIL.n195 171.744
R1329 VTAIL.n249 VTAIL.n195 171.744
R1330 VTAIL.n250 VTAIL.n249 171.744
R1331 VTAIL.n250 VTAIL.n191 171.744
R1332 VTAIL.n258 VTAIL.n191 171.744
R1333 VTAIL.n259 VTAIL.n258 171.744
R1334 VTAIL.n260 VTAIL.n259 171.744
R1335 VTAIL.n260 VTAIL.n187 171.744
R1336 VTAIL.n267 VTAIL.n187 171.744
R1337 VTAIL.n268 VTAIL.n267 171.744
R1338 VTAIL.n632 VTAIL.n631 171.744
R1339 VTAIL.n631 VTAIL.n551 171.744
R1340 VTAIL.n624 VTAIL.n551 171.744
R1341 VTAIL.n624 VTAIL.n623 171.744
R1342 VTAIL.n623 VTAIL.n622 171.744
R1343 VTAIL.n622 VTAIL.n555 171.744
R1344 VTAIL.n615 VTAIL.n555 171.744
R1345 VTAIL.n615 VTAIL.n614 171.744
R1346 VTAIL.n614 VTAIL.n560 171.744
R1347 VTAIL.n607 VTAIL.n560 171.744
R1348 VTAIL.n607 VTAIL.n606 171.744
R1349 VTAIL.n606 VTAIL.n564 171.744
R1350 VTAIL.n599 VTAIL.n564 171.744
R1351 VTAIL.n599 VTAIL.n598 171.744
R1352 VTAIL.n598 VTAIL.n568 171.744
R1353 VTAIL.n591 VTAIL.n568 171.744
R1354 VTAIL.n591 VTAIL.n590 171.744
R1355 VTAIL.n590 VTAIL.n572 171.744
R1356 VTAIL.n583 VTAIL.n572 171.744
R1357 VTAIL.n583 VTAIL.n582 171.744
R1358 VTAIL.n582 VTAIL.n576 171.744
R1359 VTAIL.n540 VTAIL.n539 171.744
R1360 VTAIL.n539 VTAIL.n459 171.744
R1361 VTAIL.n532 VTAIL.n459 171.744
R1362 VTAIL.n532 VTAIL.n531 171.744
R1363 VTAIL.n531 VTAIL.n530 171.744
R1364 VTAIL.n530 VTAIL.n463 171.744
R1365 VTAIL.n523 VTAIL.n463 171.744
R1366 VTAIL.n523 VTAIL.n522 171.744
R1367 VTAIL.n522 VTAIL.n468 171.744
R1368 VTAIL.n515 VTAIL.n468 171.744
R1369 VTAIL.n515 VTAIL.n514 171.744
R1370 VTAIL.n514 VTAIL.n472 171.744
R1371 VTAIL.n507 VTAIL.n472 171.744
R1372 VTAIL.n507 VTAIL.n506 171.744
R1373 VTAIL.n506 VTAIL.n476 171.744
R1374 VTAIL.n499 VTAIL.n476 171.744
R1375 VTAIL.n499 VTAIL.n498 171.744
R1376 VTAIL.n498 VTAIL.n480 171.744
R1377 VTAIL.n491 VTAIL.n480 171.744
R1378 VTAIL.n491 VTAIL.n490 171.744
R1379 VTAIL.n490 VTAIL.n484 171.744
R1380 VTAIL.n450 VTAIL.n449 171.744
R1381 VTAIL.n449 VTAIL.n369 171.744
R1382 VTAIL.n442 VTAIL.n369 171.744
R1383 VTAIL.n442 VTAIL.n441 171.744
R1384 VTAIL.n441 VTAIL.n440 171.744
R1385 VTAIL.n440 VTAIL.n373 171.744
R1386 VTAIL.n433 VTAIL.n373 171.744
R1387 VTAIL.n433 VTAIL.n432 171.744
R1388 VTAIL.n432 VTAIL.n378 171.744
R1389 VTAIL.n425 VTAIL.n378 171.744
R1390 VTAIL.n425 VTAIL.n424 171.744
R1391 VTAIL.n424 VTAIL.n382 171.744
R1392 VTAIL.n417 VTAIL.n382 171.744
R1393 VTAIL.n417 VTAIL.n416 171.744
R1394 VTAIL.n416 VTAIL.n386 171.744
R1395 VTAIL.n409 VTAIL.n386 171.744
R1396 VTAIL.n409 VTAIL.n408 171.744
R1397 VTAIL.n408 VTAIL.n390 171.744
R1398 VTAIL.n401 VTAIL.n390 171.744
R1399 VTAIL.n401 VTAIL.n400 171.744
R1400 VTAIL.n400 VTAIL.n394 171.744
R1401 VTAIL.n358 VTAIL.n357 171.744
R1402 VTAIL.n357 VTAIL.n277 171.744
R1403 VTAIL.n350 VTAIL.n277 171.744
R1404 VTAIL.n350 VTAIL.n349 171.744
R1405 VTAIL.n349 VTAIL.n348 171.744
R1406 VTAIL.n348 VTAIL.n281 171.744
R1407 VTAIL.n341 VTAIL.n281 171.744
R1408 VTAIL.n341 VTAIL.n340 171.744
R1409 VTAIL.n340 VTAIL.n286 171.744
R1410 VTAIL.n333 VTAIL.n286 171.744
R1411 VTAIL.n333 VTAIL.n332 171.744
R1412 VTAIL.n332 VTAIL.n290 171.744
R1413 VTAIL.n325 VTAIL.n290 171.744
R1414 VTAIL.n325 VTAIL.n324 171.744
R1415 VTAIL.n324 VTAIL.n294 171.744
R1416 VTAIL.n317 VTAIL.n294 171.744
R1417 VTAIL.n317 VTAIL.n316 171.744
R1418 VTAIL.n316 VTAIL.n298 171.744
R1419 VTAIL.n309 VTAIL.n298 171.744
R1420 VTAIL.n309 VTAIL.n308 171.744
R1421 VTAIL.n308 VTAIL.n302 171.744
R1422 VTAIL.t5 VTAIL.n665 85.8723
R1423 VTAIL.t4 VTAIL.n29 85.8723
R1424 VTAIL.t8 VTAIL.n119 85.8723
R1425 VTAIL.t10 VTAIL.n211 85.8723
R1426 VTAIL.t7 VTAIL.n576 85.8723
R1427 VTAIL.t14 VTAIL.n484 85.8723
R1428 VTAIL.t0 VTAIL.n394 85.8723
R1429 VTAIL.t15 VTAIL.n302 85.8723
R1430 VTAIL.n547 VTAIL.n546 51.9597
R1431 VTAIL.n365 VTAIL.n364 51.9597
R1432 VTAIL.n1 VTAIL.n0 51.9595
R1433 VTAIL.n183 VTAIL.n182 51.9595
R1434 VTAIL.n727 VTAIL.n726 31.0217
R1435 VTAIL.n91 VTAIL.n90 31.0217
R1436 VTAIL.n181 VTAIL.n180 31.0217
R1437 VTAIL.n273 VTAIL.n272 31.0217
R1438 VTAIL.n637 VTAIL.n636 31.0217
R1439 VTAIL.n545 VTAIL.n544 31.0217
R1440 VTAIL.n455 VTAIL.n454 31.0217
R1441 VTAIL.n363 VTAIL.n362 31.0217
R1442 VTAIL.n727 VTAIL.n637 27.091
R1443 VTAIL.n363 VTAIL.n273 27.091
R1444 VTAIL.n667 VTAIL.n666 16.3895
R1445 VTAIL.n31 VTAIL.n30 16.3895
R1446 VTAIL.n121 VTAIL.n120 16.3895
R1447 VTAIL.n213 VTAIL.n212 16.3895
R1448 VTAIL.n578 VTAIL.n577 16.3895
R1449 VTAIL.n486 VTAIL.n485 16.3895
R1450 VTAIL.n396 VTAIL.n395 16.3895
R1451 VTAIL.n304 VTAIL.n303 16.3895
R1452 VTAIL.n715 VTAIL.n644 13.1884
R1453 VTAIL.n79 VTAIL.n8 13.1884
R1454 VTAIL.n169 VTAIL.n98 13.1884
R1455 VTAIL.n261 VTAIL.n190 13.1884
R1456 VTAIL.n625 VTAIL.n554 13.1884
R1457 VTAIL.n533 VTAIL.n462 13.1884
R1458 VTAIL.n443 VTAIL.n372 13.1884
R1459 VTAIL.n351 VTAIL.n280 13.1884
R1460 VTAIL.n670 VTAIL.n669 12.8005
R1461 VTAIL.n711 VTAIL.n710 12.8005
R1462 VTAIL.n716 VTAIL.n642 12.8005
R1463 VTAIL.n34 VTAIL.n33 12.8005
R1464 VTAIL.n75 VTAIL.n74 12.8005
R1465 VTAIL.n80 VTAIL.n6 12.8005
R1466 VTAIL.n124 VTAIL.n123 12.8005
R1467 VTAIL.n165 VTAIL.n164 12.8005
R1468 VTAIL.n170 VTAIL.n96 12.8005
R1469 VTAIL.n216 VTAIL.n215 12.8005
R1470 VTAIL.n257 VTAIL.n256 12.8005
R1471 VTAIL.n262 VTAIL.n188 12.8005
R1472 VTAIL.n626 VTAIL.n552 12.8005
R1473 VTAIL.n621 VTAIL.n556 12.8005
R1474 VTAIL.n581 VTAIL.n580 12.8005
R1475 VTAIL.n534 VTAIL.n460 12.8005
R1476 VTAIL.n529 VTAIL.n464 12.8005
R1477 VTAIL.n489 VTAIL.n488 12.8005
R1478 VTAIL.n444 VTAIL.n370 12.8005
R1479 VTAIL.n439 VTAIL.n374 12.8005
R1480 VTAIL.n399 VTAIL.n398 12.8005
R1481 VTAIL.n352 VTAIL.n278 12.8005
R1482 VTAIL.n347 VTAIL.n282 12.8005
R1483 VTAIL.n307 VTAIL.n306 12.8005
R1484 VTAIL.n673 VTAIL.n664 12.0247
R1485 VTAIL.n709 VTAIL.n646 12.0247
R1486 VTAIL.n720 VTAIL.n719 12.0247
R1487 VTAIL.n37 VTAIL.n28 12.0247
R1488 VTAIL.n73 VTAIL.n10 12.0247
R1489 VTAIL.n84 VTAIL.n83 12.0247
R1490 VTAIL.n127 VTAIL.n118 12.0247
R1491 VTAIL.n163 VTAIL.n100 12.0247
R1492 VTAIL.n174 VTAIL.n173 12.0247
R1493 VTAIL.n219 VTAIL.n210 12.0247
R1494 VTAIL.n255 VTAIL.n192 12.0247
R1495 VTAIL.n266 VTAIL.n265 12.0247
R1496 VTAIL.n630 VTAIL.n629 12.0247
R1497 VTAIL.n620 VTAIL.n557 12.0247
R1498 VTAIL.n584 VTAIL.n575 12.0247
R1499 VTAIL.n538 VTAIL.n537 12.0247
R1500 VTAIL.n528 VTAIL.n465 12.0247
R1501 VTAIL.n492 VTAIL.n483 12.0247
R1502 VTAIL.n448 VTAIL.n447 12.0247
R1503 VTAIL.n438 VTAIL.n375 12.0247
R1504 VTAIL.n402 VTAIL.n393 12.0247
R1505 VTAIL.n356 VTAIL.n355 12.0247
R1506 VTAIL.n346 VTAIL.n283 12.0247
R1507 VTAIL.n310 VTAIL.n301 12.0247
R1508 VTAIL.n674 VTAIL.n662 11.249
R1509 VTAIL.n706 VTAIL.n705 11.249
R1510 VTAIL.n723 VTAIL.n640 11.249
R1511 VTAIL.n38 VTAIL.n26 11.249
R1512 VTAIL.n70 VTAIL.n69 11.249
R1513 VTAIL.n87 VTAIL.n4 11.249
R1514 VTAIL.n128 VTAIL.n116 11.249
R1515 VTAIL.n160 VTAIL.n159 11.249
R1516 VTAIL.n177 VTAIL.n94 11.249
R1517 VTAIL.n220 VTAIL.n208 11.249
R1518 VTAIL.n252 VTAIL.n251 11.249
R1519 VTAIL.n269 VTAIL.n186 11.249
R1520 VTAIL.n633 VTAIL.n550 11.249
R1521 VTAIL.n617 VTAIL.n616 11.249
R1522 VTAIL.n585 VTAIL.n573 11.249
R1523 VTAIL.n541 VTAIL.n458 11.249
R1524 VTAIL.n525 VTAIL.n524 11.249
R1525 VTAIL.n493 VTAIL.n481 11.249
R1526 VTAIL.n451 VTAIL.n368 11.249
R1527 VTAIL.n435 VTAIL.n434 11.249
R1528 VTAIL.n403 VTAIL.n391 11.249
R1529 VTAIL.n359 VTAIL.n276 11.249
R1530 VTAIL.n343 VTAIL.n342 11.249
R1531 VTAIL.n311 VTAIL.n299 11.249
R1532 VTAIL.n678 VTAIL.n677 10.4732
R1533 VTAIL.n702 VTAIL.n648 10.4732
R1534 VTAIL.n724 VTAIL.n638 10.4732
R1535 VTAIL.n42 VTAIL.n41 10.4732
R1536 VTAIL.n66 VTAIL.n12 10.4732
R1537 VTAIL.n88 VTAIL.n2 10.4732
R1538 VTAIL.n132 VTAIL.n131 10.4732
R1539 VTAIL.n156 VTAIL.n102 10.4732
R1540 VTAIL.n178 VTAIL.n92 10.4732
R1541 VTAIL.n224 VTAIL.n223 10.4732
R1542 VTAIL.n248 VTAIL.n194 10.4732
R1543 VTAIL.n270 VTAIL.n184 10.4732
R1544 VTAIL.n634 VTAIL.n548 10.4732
R1545 VTAIL.n613 VTAIL.n559 10.4732
R1546 VTAIL.n589 VTAIL.n588 10.4732
R1547 VTAIL.n542 VTAIL.n456 10.4732
R1548 VTAIL.n521 VTAIL.n467 10.4732
R1549 VTAIL.n497 VTAIL.n496 10.4732
R1550 VTAIL.n452 VTAIL.n366 10.4732
R1551 VTAIL.n431 VTAIL.n377 10.4732
R1552 VTAIL.n407 VTAIL.n406 10.4732
R1553 VTAIL.n360 VTAIL.n274 10.4732
R1554 VTAIL.n339 VTAIL.n285 10.4732
R1555 VTAIL.n315 VTAIL.n314 10.4732
R1556 VTAIL.n681 VTAIL.n660 9.69747
R1557 VTAIL.n701 VTAIL.n650 9.69747
R1558 VTAIL.n45 VTAIL.n24 9.69747
R1559 VTAIL.n65 VTAIL.n14 9.69747
R1560 VTAIL.n135 VTAIL.n114 9.69747
R1561 VTAIL.n155 VTAIL.n104 9.69747
R1562 VTAIL.n227 VTAIL.n206 9.69747
R1563 VTAIL.n247 VTAIL.n196 9.69747
R1564 VTAIL.n612 VTAIL.n561 9.69747
R1565 VTAIL.n592 VTAIL.n571 9.69747
R1566 VTAIL.n520 VTAIL.n469 9.69747
R1567 VTAIL.n500 VTAIL.n479 9.69747
R1568 VTAIL.n430 VTAIL.n379 9.69747
R1569 VTAIL.n410 VTAIL.n389 9.69747
R1570 VTAIL.n338 VTAIL.n287 9.69747
R1571 VTAIL.n318 VTAIL.n297 9.69747
R1572 VTAIL.n726 VTAIL.n725 9.45567
R1573 VTAIL.n90 VTAIL.n89 9.45567
R1574 VTAIL.n180 VTAIL.n179 9.45567
R1575 VTAIL.n272 VTAIL.n271 9.45567
R1576 VTAIL.n636 VTAIL.n635 9.45567
R1577 VTAIL.n544 VTAIL.n543 9.45567
R1578 VTAIL.n454 VTAIL.n453 9.45567
R1579 VTAIL.n362 VTAIL.n361 9.45567
R1580 VTAIL.n725 VTAIL.n724 9.3005
R1581 VTAIL.n640 VTAIL.n639 9.3005
R1582 VTAIL.n719 VTAIL.n718 9.3005
R1583 VTAIL.n717 VTAIL.n716 9.3005
R1584 VTAIL.n656 VTAIL.n655 9.3005
R1585 VTAIL.n685 VTAIL.n684 9.3005
R1586 VTAIL.n683 VTAIL.n682 9.3005
R1587 VTAIL.n660 VTAIL.n659 9.3005
R1588 VTAIL.n677 VTAIL.n676 9.3005
R1589 VTAIL.n675 VTAIL.n674 9.3005
R1590 VTAIL.n664 VTAIL.n663 9.3005
R1591 VTAIL.n669 VTAIL.n668 9.3005
R1592 VTAIL.n691 VTAIL.n690 9.3005
R1593 VTAIL.n693 VTAIL.n692 9.3005
R1594 VTAIL.n652 VTAIL.n651 9.3005
R1595 VTAIL.n699 VTAIL.n698 9.3005
R1596 VTAIL.n701 VTAIL.n700 9.3005
R1597 VTAIL.n648 VTAIL.n647 9.3005
R1598 VTAIL.n707 VTAIL.n706 9.3005
R1599 VTAIL.n709 VTAIL.n708 9.3005
R1600 VTAIL.n710 VTAIL.n643 9.3005
R1601 VTAIL.n89 VTAIL.n88 9.3005
R1602 VTAIL.n4 VTAIL.n3 9.3005
R1603 VTAIL.n83 VTAIL.n82 9.3005
R1604 VTAIL.n81 VTAIL.n80 9.3005
R1605 VTAIL.n20 VTAIL.n19 9.3005
R1606 VTAIL.n49 VTAIL.n48 9.3005
R1607 VTAIL.n47 VTAIL.n46 9.3005
R1608 VTAIL.n24 VTAIL.n23 9.3005
R1609 VTAIL.n41 VTAIL.n40 9.3005
R1610 VTAIL.n39 VTAIL.n38 9.3005
R1611 VTAIL.n28 VTAIL.n27 9.3005
R1612 VTAIL.n33 VTAIL.n32 9.3005
R1613 VTAIL.n55 VTAIL.n54 9.3005
R1614 VTAIL.n57 VTAIL.n56 9.3005
R1615 VTAIL.n16 VTAIL.n15 9.3005
R1616 VTAIL.n63 VTAIL.n62 9.3005
R1617 VTAIL.n65 VTAIL.n64 9.3005
R1618 VTAIL.n12 VTAIL.n11 9.3005
R1619 VTAIL.n71 VTAIL.n70 9.3005
R1620 VTAIL.n73 VTAIL.n72 9.3005
R1621 VTAIL.n74 VTAIL.n7 9.3005
R1622 VTAIL.n179 VTAIL.n178 9.3005
R1623 VTAIL.n94 VTAIL.n93 9.3005
R1624 VTAIL.n173 VTAIL.n172 9.3005
R1625 VTAIL.n171 VTAIL.n170 9.3005
R1626 VTAIL.n110 VTAIL.n109 9.3005
R1627 VTAIL.n139 VTAIL.n138 9.3005
R1628 VTAIL.n137 VTAIL.n136 9.3005
R1629 VTAIL.n114 VTAIL.n113 9.3005
R1630 VTAIL.n131 VTAIL.n130 9.3005
R1631 VTAIL.n129 VTAIL.n128 9.3005
R1632 VTAIL.n118 VTAIL.n117 9.3005
R1633 VTAIL.n123 VTAIL.n122 9.3005
R1634 VTAIL.n145 VTAIL.n144 9.3005
R1635 VTAIL.n147 VTAIL.n146 9.3005
R1636 VTAIL.n106 VTAIL.n105 9.3005
R1637 VTAIL.n153 VTAIL.n152 9.3005
R1638 VTAIL.n155 VTAIL.n154 9.3005
R1639 VTAIL.n102 VTAIL.n101 9.3005
R1640 VTAIL.n161 VTAIL.n160 9.3005
R1641 VTAIL.n163 VTAIL.n162 9.3005
R1642 VTAIL.n164 VTAIL.n97 9.3005
R1643 VTAIL.n271 VTAIL.n270 9.3005
R1644 VTAIL.n186 VTAIL.n185 9.3005
R1645 VTAIL.n265 VTAIL.n264 9.3005
R1646 VTAIL.n263 VTAIL.n262 9.3005
R1647 VTAIL.n202 VTAIL.n201 9.3005
R1648 VTAIL.n231 VTAIL.n230 9.3005
R1649 VTAIL.n229 VTAIL.n228 9.3005
R1650 VTAIL.n206 VTAIL.n205 9.3005
R1651 VTAIL.n223 VTAIL.n222 9.3005
R1652 VTAIL.n221 VTAIL.n220 9.3005
R1653 VTAIL.n210 VTAIL.n209 9.3005
R1654 VTAIL.n215 VTAIL.n214 9.3005
R1655 VTAIL.n237 VTAIL.n236 9.3005
R1656 VTAIL.n239 VTAIL.n238 9.3005
R1657 VTAIL.n198 VTAIL.n197 9.3005
R1658 VTAIL.n245 VTAIL.n244 9.3005
R1659 VTAIL.n247 VTAIL.n246 9.3005
R1660 VTAIL.n194 VTAIL.n193 9.3005
R1661 VTAIL.n253 VTAIL.n252 9.3005
R1662 VTAIL.n255 VTAIL.n254 9.3005
R1663 VTAIL.n256 VTAIL.n189 9.3005
R1664 VTAIL.n604 VTAIL.n603 9.3005
R1665 VTAIL.n563 VTAIL.n562 9.3005
R1666 VTAIL.n610 VTAIL.n609 9.3005
R1667 VTAIL.n612 VTAIL.n611 9.3005
R1668 VTAIL.n559 VTAIL.n558 9.3005
R1669 VTAIL.n618 VTAIL.n617 9.3005
R1670 VTAIL.n620 VTAIL.n619 9.3005
R1671 VTAIL.n556 VTAIL.n553 9.3005
R1672 VTAIL.n635 VTAIL.n634 9.3005
R1673 VTAIL.n550 VTAIL.n549 9.3005
R1674 VTAIL.n629 VTAIL.n628 9.3005
R1675 VTAIL.n627 VTAIL.n626 9.3005
R1676 VTAIL.n602 VTAIL.n601 9.3005
R1677 VTAIL.n567 VTAIL.n566 9.3005
R1678 VTAIL.n596 VTAIL.n595 9.3005
R1679 VTAIL.n594 VTAIL.n593 9.3005
R1680 VTAIL.n571 VTAIL.n570 9.3005
R1681 VTAIL.n588 VTAIL.n587 9.3005
R1682 VTAIL.n586 VTAIL.n585 9.3005
R1683 VTAIL.n575 VTAIL.n574 9.3005
R1684 VTAIL.n580 VTAIL.n579 9.3005
R1685 VTAIL.n512 VTAIL.n511 9.3005
R1686 VTAIL.n471 VTAIL.n470 9.3005
R1687 VTAIL.n518 VTAIL.n517 9.3005
R1688 VTAIL.n520 VTAIL.n519 9.3005
R1689 VTAIL.n467 VTAIL.n466 9.3005
R1690 VTAIL.n526 VTAIL.n525 9.3005
R1691 VTAIL.n528 VTAIL.n527 9.3005
R1692 VTAIL.n464 VTAIL.n461 9.3005
R1693 VTAIL.n543 VTAIL.n542 9.3005
R1694 VTAIL.n458 VTAIL.n457 9.3005
R1695 VTAIL.n537 VTAIL.n536 9.3005
R1696 VTAIL.n535 VTAIL.n534 9.3005
R1697 VTAIL.n510 VTAIL.n509 9.3005
R1698 VTAIL.n475 VTAIL.n474 9.3005
R1699 VTAIL.n504 VTAIL.n503 9.3005
R1700 VTAIL.n502 VTAIL.n501 9.3005
R1701 VTAIL.n479 VTAIL.n478 9.3005
R1702 VTAIL.n496 VTAIL.n495 9.3005
R1703 VTAIL.n494 VTAIL.n493 9.3005
R1704 VTAIL.n483 VTAIL.n482 9.3005
R1705 VTAIL.n488 VTAIL.n487 9.3005
R1706 VTAIL.n422 VTAIL.n421 9.3005
R1707 VTAIL.n381 VTAIL.n380 9.3005
R1708 VTAIL.n428 VTAIL.n427 9.3005
R1709 VTAIL.n430 VTAIL.n429 9.3005
R1710 VTAIL.n377 VTAIL.n376 9.3005
R1711 VTAIL.n436 VTAIL.n435 9.3005
R1712 VTAIL.n438 VTAIL.n437 9.3005
R1713 VTAIL.n374 VTAIL.n371 9.3005
R1714 VTAIL.n453 VTAIL.n452 9.3005
R1715 VTAIL.n368 VTAIL.n367 9.3005
R1716 VTAIL.n447 VTAIL.n446 9.3005
R1717 VTAIL.n445 VTAIL.n444 9.3005
R1718 VTAIL.n420 VTAIL.n419 9.3005
R1719 VTAIL.n385 VTAIL.n384 9.3005
R1720 VTAIL.n414 VTAIL.n413 9.3005
R1721 VTAIL.n412 VTAIL.n411 9.3005
R1722 VTAIL.n389 VTAIL.n388 9.3005
R1723 VTAIL.n406 VTAIL.n405 9.3005
R1724 VTAIL.n404 VTAIL.n403 9.3005
R1725 VTAIL.n393 VTAIL.n392 9.3005
R1726 VTAIL.n398 VTAIL.n397 9.3005
R1727 VTAIL.n330 VTAIL.n329 9.3005
R1728 VTAIL.n289 VTAIL.n288 9.3005
R1729 VTAIL.n336 VTAIL.n335 9.3005
R1730 VTAIL.n338 VTAIL.n337 9.3005
R1731 VTAIL.n285 VTAIL.n284 9.3005
R1732 VTAIL.n344 VTAIL.n343 9.3005
R1733 VTAIL.n346 VTAIL.n345 9.3005
R1734 VTAIL.n282 VTAIL.n279 9.3005
R1735 VTAIL.n361 VTAIL.n360 9.3005
R1736 VTAIL.n276 VTAIL.n275 9.3005
R1737 VTAIL.n355 VTAIL.n354 9.3005
R1738 VTAIL.n353 VTAIL.n352 9.3005
R1739 VTAIL.n328 VTAIL.n327 9.3005
R1740 VTAIL.n293 VTAIL.n292 9.3005
R1741 VTAIL.n322 VTAIL.n321 9.3005
R1742 VTAIL.n320 VTAIL.n319 9.3005
R1743 VTAIL.n297 VTAIL.n296 9.3005
R1744 VTAIL.n314 VTAIL.n313 9.3005
R1745 VTAIL.n312 VTAIL.n311 9.3005
R1746 VTAIL.n301 VTAIL.n300 9.3005
R1747 VTAIL.n306 VTAIL.n305 9.3005
R1748 VTAIL.n682 VTAIL.n658 8.92171
R1749 VTAIL.n698 VTAIL.n697 8.92171
R1750 VTAIL.n46 VTAIL.n22 8.92171
R1751 VTAIL.n62 VTAIL.n61 8.92171
R1752 VTAIL.n136 VTAIL.n112 8.92171
R1753 VTAIL.n152 VTAIL.n151 8.92171
R1754 VTAIL.n228 VTAIL.n204 8.92171
R1755 VTAIL.n244 VTAIL.n243 8.92171
R1756 VTAIL.n609 VTAIL.n608 8.92171
R1757 VTAIL.n593 VTAIL.n569 8.92171
R1758 VTAIL.n517 VTAIL.n516 8.92171
R1759 VTAIL.n501 VTAIL.n477 8.92171
R1760 VTAIL.n427 VTAIL.n426 8.92171
R1761 VTAIL.n411 VTAIL.n387 8.92171
R1762 VTAIL.n335 VTAIL.n334 8.92171
R1763 VTAIL.n319 VTAIL.n295 8.92171
R1764 VTAIL.n686 VTAIL.n685 8.14595
R1765 VTAIL.n694 VTAIL.n652 8.14595
R1766 VTAIL.n50 VTAIL.n49 8.14595
R1767 VTAIL.n58 VTAIL.n16 8.14595
R1768 VTAIL.n140 VTAIL.n139 8.14595
R1769 VTAIL.n148 VTAIL.n106 8.14595
R1770 VTAIL.n232 VTAIL.n231 8.14595
R1771 VTAIL.n240 VTAIL.n198 8.14595
R1772 VTAIL.n605 VTAIL.n563 8.14595
R1773 VTAIL.n597 VTAIL.n596 8.14595
R1774 VTAIL.n513 VTAIL.n471 8.14595
R1775 VTAIL.n505 VTAIL.n504 8.14595
R1776 VTAIL.n423 VTAIL.n381 8.14595
R1777 VTAIL.n415 VTAIL.n414 8.14595
R1778 VTAIL.n331 VTAIL.n289 8.14595
R1779 VTAIL.n323 VTAIL.n322 8.14595
R1780 VTAIL.n689 VTAIL.n656 7.3702
R1781 VTAIL.n693 VTAIL.n654 7.3702
R1782 VTAIL.n53 VTAIL.n20 7.3702
R1783 VTAIL.n57 VTAIL.n18 7.3702
R1784 VTAIL.n143 VTAIL.n110 7.3702
R1785 VTAIL.n147 VTAIL.n108 7.3702
R1786 VTAIL.n235 VTAIL.n202 7.3702
R1787 VTAIL.n239 VTAIL.n200 7.3702
R1788 VTAIL.n604 VTAIL.n565 7.3702
R1789 VTAIL.n600 VTAIL.n567 7.3702
R1790 VTAIL.n512 VTAIL.n473 7.3702
R1791 VTAIL.n508 VTAIL.n475 7.3702
R1792 VTAIL.n422 VTAIL.n383 7.3702
R1793 VTAIL.n418 VTAIL.n385 7.3702
R1794 VTAIL.n330 VTAIL.n291 7.3702
R1795 VTAIL.n326 VTAIL.n293 7.3702
R1796 VTAIL.n690 VTAIL.n689 6.59444
R1797 VTAIL.n690 VTAIL.n654 6.59444
R1798 VTAIL.n54 VTAIL.n53 6.59444
R1799 VTAIL.n54 VTAIL.n18 6.59444
R1800 VTAIL.n144 VTAIL.n143 6.59444
R1801 VTAIL.n144 VTAIL.n108 6.59444
R1802 VTAIL.n236 VTAIL.n235 6.59444
R1803 VTAIL.n236 VTAIL.n200 6.59444
R1804 VTAIL.n601 VTAIL.n565 6.59444
R1805 VTAIL.n601 VTAIL.n600 6.59444
R1806 VTAIL.n509 VTAIL.n473 6.59444
R1807 VTAIL.n509 VTAIL.n508 6.59444
R1808 VTAIL.n419 VTAIL.n383 6.59444
R1809 VTAIL.n419 VTAIL.n418 6.59444
R1810 VTAIL.n327 VTAIL.n291 6.59444
R1811 VTAIL.n327 VTAIL.n326 6.59444
R1812 VTAIL.n686 VTAIL.n656 5.81868
R1813 VTAIL.n694 VTAIL.n693 5.81868
R1814 VTAIL.n50 VTAIL.n20 5.81868
R1815 VTAIL.n58 VTAIL.n57 5.81868
R1816 VTAIL.n140 VTAIL.n110 5.81868
R1817 VTAIL.n148 VTAIL.n147 5.81868
R1818 VTAIL.n232 VTAIL.n202 5.81868
R1819 VTAIL.n240 VTAIL.n239 5.81868
R1820 VTAIL.n605 VTAIL.n604 5.81868
R1821 VTAIL.n597 VTAIL.n567 5.81868
R1822 VTAIL.n513 VTAIL.n512 5.81868
R1823 VTAIL.n505 VTAIL.n475 5.81868
R1824 VTAIL.n423 VTAIL.n422 5.81868
R1825 VTAIL.n415 VTAIL.n385 5.81868
R1826 VTAIL.n331 VTAIL.n330 5.81868
R1827 VTAIL.n323 VTAIL.n293 5.81868
R1828 VTAIL.n685 VTAIL.n658 5.04292
R1829 VTAIL.n697 VTAIL.n652 5.04292
R1830 VTAIL.n49 VTAIL.n22 5.04292
R1831 VTAIL.n61 VTAIL.n16 5.04292
R1832 VTAIL.n139 VTAIL.n112 5.04292
R1833 VTAIL.n151 VTAIL.n106 5.04292
R1834 VTAIL.n231 VTAIL.n204 5.04292
R1835 VTAIL.n243 VTAIL.n198 5.04292
R1836 VTAIL.n608 VTAIL.n563 5.04292
R1837 VTAIL.n596 VTAIL.n569 5.04292
R1838 VTAIL.n516 VTAIL.n471 5.04292
R1839 VTAIL.n504 VTAIL.n477 5.04292
R1840 VTAIL.n426 VTAIL.n381 5.04292
R1841 VTAIL.n414 VTAIL.n387 5.04292
R1842 VTAIL.n334 VTAIL.n289 5.04292
R1843 VTAIL.n322 VTAIL.n295 5.04292
R1844 VTAIL.n682 VTAIL.n681 4.26717
R1845 VTAIL.n698 VTAIL.n650 4.26717
R1846 VTAIL.n46 VTAIL.n45 4.26717
R1847 VTAIL.n62 VTAIL.n14 4.26717
R1848 VTAIL.n136 VTAIL.n135 4.26717
R1849 VTAIL.n152 VTAIL.n104 4.26717
R1850 VTAIL.n228 VTAIL.n227 4.26717
R1851 VTAIL.n244 VTAIL.n196 4.26717
R1852 VTAIL.n609 VTAIL.n561 4.26717
R1853 VTAIL.n593 VTAIL.n592 4.26717
R1854 VTAIL.n517 VTAIL.n469 4.26717
R1855 VTAIL.n501 VTAIL.n500 4.26717
R1856 VTAIL.n427 VTAIL.n379 4.26717
R1857 VTAIL.n411 VTAIL.n410 4.26717
R1858 VTAIL.n335 VTAIL.n287 4.26717
R1859 VTAIL.n319 VTAIL.n318 4.26717
R1860 VTAIL.n668 VTAIL.n667 3.70982
R1861 VTAIL.n32 VTAIL.n31 3.70982
R1862 VTAIL.n122 VTAIL.n121 3.70982
R1863 VTAIL.n214 VTAIL.n213 3.70982
R1864 VTAIL.n579 VTAIL.n578 3.70982
R1865 VTAIL.n487 VTAIL.n486 3.70982
R1866 VTAIL.n397 VTAIL.n396 3.70982
R1867 VTAIL.n305 VTAIL.n304 3.70982
R1868 VTAIL.n678 VTAIL.n660 3.49141
R1869 VTAIL.n702 VTAIL.n701 3.49141
R1870 VTAIL.n726 VTAIL.n638 3.49141
R1871 VTAIL.n42 VTAIL.n24 3.49141
R1872 VTAIL.n66 VTAIL.n65 3.49141
R1873 VTAIL.n90 VTAIL.n2 3.49141
R1874 VTAIL.n132 VTAIL.n114 3.49141
R1875 VTAIL.n156 VTAIL.n155 3.49141
R1876 VTAIL.n180 VTAIL.n92 3.49141
R1877 VTAIL.n224 VTAIL.n206 3.49141
R1878 VTAIL.n248 VTAIL.n247 3.49141
R1879 VTAIL.n272 VTAIL.n184 3.49141
R1880 VTAIL.n636 VTAIL.n548 3.49141
R1881 VTAIL.n613 VTAIL.n612 3.49141
R1882 VTAIL.n589 VTAIL.n571 3.49141
R1883 VTAIL.n544 VTAIL.n456 3.49141
R1884 VTAIL.n521 VTAIL.n520 3.49141
R1885 VTAIL.n497 VTAIL.n479 3.49141
R1886 VTAIL.n454 VTAIL.n366 3.49141
R1887 VTAIL.n431 VTAIL.n430 3.49141
R1888 VTAIL.n407 VTAIL.n389 3.49141
R1889 VTAIL.n362 VTAIL.n274 3.49141
R1890 VTAIL.n339 VTAIL.n338 3.49141
R1891 VTAIL.n315 VTAIL.n297 3.49141
R1892 VTAIL.n677 VTAIL.n662 2.71565
R1893 VTAIL.n705 VTAIL.n648 2.71565
R1894 VTAIL.n724 VTAIL.n723 2.71565
R1895 VTAIL.n41 VTAIL.n26 2.71565
R1896 VTAIL.n69 VTAIL.n12 2.71565
R1897 VTAIL.n88 VTAIL.n87 2.71565
R1898 VTAIL.n131 VTAIL.n116 2.71565
R1899 VTAIL.n159 VTAIL.n102 2.71565
R1900 VTAIL.n178 VTAIL.n177 2.71565
R1901 VTAIL.n223 VTAIL.n208 2.71565
R1902 VTAIL.n251 VTAIL.n194 2.71565
R1903 VTAIL.n270 VTAIL.n269 2.71565
R1904 VTAIL.n634 VTAIL.n633 2.71565
R1905 VTAIL.n616 VTAIL.n559 2.71565
R1906 VTAIL.n588 VTAIL.n573 2.71565
R1907 VTAIL.n542 VTAIL.n541 2.71565
R1908 VTAIL.n524 VTAIL.n467 2.71565
R1909 VTAIL.n496 VTAIL.n481 2.71565
R1910 VTAIL.n452 VTAIL.n451 2.71565
R1911 VTAIL.n434 VTAIL.n377 2.71565
R1912 VTAIL.n406 VTAIL.n391 2.71565
R1913 VTAIL.n360 VTAIL.n359 2.71565
R1914 VTAIL.n342 VTAIL.n285 2.71565
R1915 VTAIL.n314 VTAIL.n299 2.71565
R1916 VTAIL.n0 VTAIL.t2 2.02953
R1917 VTAIL.n0 VTAIL.t3 2.02953
R1918 VTAIL.n182 VTAIL.t11 2.02953
R1919 VTAIL.n182 VTAIL.t9 2.02953
R1920 VTAIL.n546 VTAIL.t12 2.02953
R1921 VTAIL.n546 VTAIL.t13 2.02953
R1922 VTAIL.n364 VTAIL.t1 2.02953
R1923 VTAIL.n364 VTAIL.t6 2.02953
R1924 VTAIL.n674 VTAIL.n673 1.93989
R1925 VTAIL.n706 VTAIL.n646 1.93989
R1926 VTAIL.n720 VTAIL.n640 1.93989
R1927 VTAIL.n38 VTAIL.n37 1.93989
R1928 VTAIL.n70 VTAIL.n10 1.93989
R1929 VTAIL.n84 VTAIL.n4 1.93989
R1930 VTAIL.n128 VTAIL.n127 1.93989
R1931 VTAIL.n160 VTAIL.n100 1.93989
R1932 VTAIL.n174 VTAIL.n94 1.93989
R1933 VTAIL.n220 VTAIL.n219 1.93989
R1934 VTAIL.n252 VTAIL.n192 1.93989
R1935 VTAIL.n266 VTAIL.n186 1.93989
R1936 VTAIL.n630 VTAIL.n550 1.93989
R1937 VTAIL.n617 VTAIL.n557 1.93989
R1938 VTAIL.n585 VTAIL.n584 1.93989
R1939 VTAIL.n538 VTAIL.n458 1.93989
R1940 VTAIL.n525 VTAIL.n465 1.93989
R1941 VTAIL.n493 VTAIL.n492 1.93989
R1942 VTAIL.n448 VTAIL.n368 1.93989
R1943 VTAIL.n435 VTAIL.n375 1.93989
R1944 VTAIL.n403 VTAIL.n402 1.93989
R1945 VTAIL.n356 VTAIL.n276 1.93989
R1946 VTAIL.n343 VTAIL.n283 1.93989
R1947 VTAIL.n311 VTAIL.n310 1.93989
R1948 VTAIL.n670 VTAIL.n664 1.16414
R1949 VTAIL.n711 VTAIL.n709 1.16414
R1950 VTAIL.n719 VTAIL.n642 1.16414
R1951 VTAIL.n34 VTAIL.n28 1.16414
R1952 VTAIL.n75 VTAIL.n73 1.16414
R1953 VTAIL.n83 VTAIL.n6 1.16414
R1954 VTAIL.n124 VTAIL.n118 1.16414
R1955 VTAIL.n165 VTAIL.n163 1.16414
R1956 VTAIL.n173 VTAIL.n96 1.16414
R1957 VTAIL.n216 VTAIL.n210 1.16414
R1958 VTAIL.n257 VTAIL.n255 1.16414
R1959 VTAIL.n265 VTAIL.n188 1.16414
R1960 VTAIL.n629 VTAIL.n552 1.16414
R1961 VTAIL.n621 VTAIL.n620 1.16414
R1962 VTAIL.n581 VTAIL.n575 1.16414
R1963 VTAIL.n537 VTAIL.n460 1.16414
R1964 VTAIL.n529 VTAIL.n528 1.16414
R1965 VTAIL.n489 VTAIL.n483 1.16414
R1966 VTAIL.n447 VTAIL.n370 1.16414
R1967 VTAIL.n439 VTAIL.n438 1.16414
R1968 VTAIL.n399 VTAIL.n393 1.16414
R1969 VTAIL.n355 VTAIL.n278 1.16414
R1970 VTAIL.n347 VTAIL.n346 1.16414
R1971 VTAIL.n307 VTAIL.n301 1.16414
R1972 VTAIL.n365 VTAIL.n363 0.914293
R1973 VTAIL.n455 VTAIL.n365 0.914293
R1974 VTAIL.n547 VTAIL.n545 0.914293
R1975 VTAIL.n637 VTAIL.n547 0.914293
R1976 VTAIL.n273 VTAIL.n183 0.914293
R1977 VTAIL.n183 VTAIL.n181 0.914293
R1978 VTAIL.n91 VTAIL.n1 0.914293
R1979 VTAIL VTAIL.n727 0.856103
R1980 VTAIL.n545 VTAIL.n455 0.470328
R1981 VTAIL.n181 VTAIL.n91 0.470328
R1982 VTAIL.n669 VTAIL.n666 0.388379
R1983 VTAIL.n710 VTAIL.n644 0.388379
R1984 VTAIL.n716 VTAIL.n715 0.388379
R1985 VTAIL.n33 VTAIL.n30 0.388379
R1986 VTAIL.n74 VTAIL.n8 0.388379
R1987 VTAIL.n80 VTAIL.n79 0.388379
R1988 VTAIL.n123 VTAIL.n120 0.388379
R1989 VTAIL.n164 VTAIL.n98 0.388379
R1990 VTAIL.n170 VTAIL.n169 0.388379
R1991 VTAIL.n215 VTAIL.n212 0.388379
R1992 VTAIL.n256 VTAIL.n190 0.388379
R1993 VTAIL.n262 VTAIL.n261 0.388379
R1994 VTAIL.n626 VTAIL.n625 0.388379
R1995 VTAIL.n556 VTAIL.n554 0.388379
R1996 VTAIL.n580 VTAIL.n577 0.388379
R1997 VTAIL.n534 VTAIL.n533 0.388379
R1998 VTAIL.n464 VTAIL.n462 0.388379
R1999 VTAIL.n488 VTAIL.n485 0.388379
R2000 VTAIL.n444 VTAIL.n443 0.388379
R2001 VTAIL.n374 VTAIL.n372 0.388379
R2002 VTAIL.n398 VTAIL.n395 0.388379
R2003 VTAIL.n352 VTAIL.n351 0.388379
R2004 VTAIL.n282 VTAIL.n280 0.388379
R2005 VTAIL.n306 VTAIL.n303 0.388379
R2006 VTAIL.n668 VTAIL.n663 0.155672
R2007 VTAIL.n675 VTAIL.n663 0.155672
R2008 VTAIL.n676 VTAIL.n675 0.155672
R2009 VTAIL.n676 VTAIL.n659 0.155672
R2010 VTAIL.n683 VTAIL.n659 0.155672
R2011 VTAIL.n684 VTAIL.n683 0.155672
R2012 VTAIL.n684 VTAIL.n655 0.155672
R2013 VTAIL.n691 VTAIL.n655 0.155672
R2014 VTAIL.n692 VTAIL.n691 0.155672
R2015 VTAIL.n692 VTAIL.n651 0.155672
R2016 VTAIL.n699 VTAIL.n651 0.155672
R2017 VTAIL.n700 VTAIL.n699 0.155672
R2018 VTAIL.n700 VTAIL.n647 0.155672
R2019 VTAIL.n707 VTAIL.n647 0.155672
R2020 VTAIL.n708 VTAIL.n707 0.155672
R2021 VTAIL.n708 VTAIL.n643 0.155672
R2022 VTAIL.n717 VTAIL.n643 0.155672
R2023 VTAIL.n718 VTAIL.n717 0.155672
R2024 VTAIL.n718 VTAIL.n639 0.155672
R2025 VTAIL.n725 VTAIL.n639 0.155672
R2026 VTAIL.n32 VTAIL.n27 0.155672
R2027 VTAIL.n39 VTAIL.n27 0.155672
R2028 VTAIL.n40 VTAIL.n39 0.155672
R2029 VTAIL.n40 VTAIL.n23 0.155672
R2030 VTAIL.n47 VTAIL.n23 0.155672
R2031 VTAIL.n48 VTAIL.n47 0.155672
R2032 VTAIL.n48 VTAIL.n19 0.155672
R2033 VTAIL.n55 VTAIL.n19 0.155672
R2034 VTAIL.n56 VTAIL.n55 0.155672
R2035 VTAIL.n56 VTAIL.n15 0.155672
R2036 VTAIL.n63 VTAIL.n15 0.155672
R2037 VTAIL.n64 VTAIL.n63 0.155672
R2038 VTAIL.n64 VTAIL.n11 0.155672
R2039 VTAIL.n71 VTAIL.n11 0.155672
R2040 VTAIL.n72 VTAIL.n71 0.155672
R2041 VTAIL.n72 VTAIL.n7 0.155672
R2042 VTAIL.n81 VTAIL.n7 0.155672
R2043 VTAIL.n82 VTAIL.n81 0.155672
R2044 VTAIL.n82 VTAIL.n3 0.155672
R2045 VTAIL.n89 VTAIL.n3 0.155672
R2046 VTAIL.n122 VTAIL.n117 0.155672
R2047 VTAIL.n129 VTAIL.n117 0.155672
R2048 VTAIL.n130 VTAIL.n129 0.155672
R2049 VTAIL.n130 VTAIL.n113 0.155672
R2050 VTAIL.n137 VTAIL.n113 0.155672
R2051 VTAIL.n138 VTAIL.n137 0.155672
R2052 VTAIL.n138 VTAIL.n109 0.155672
R2053 VTAIL.n145 VTAIL.n109 0.155672
R2054 VTAIL.n146 VTAIL.n145 0.155672
R2055 VTAIL.n146 VTAIL.n105 0.155672
R2056 VTAIL.n153 VTAIL.n105 0.155672
R2057 VTAIL.n154 VTAIL.n153 0.155672
R2058 VTAIL.n154 VTAIL.n101 0.155672
R2059 VTAIL.n161 VTAIL.n101 0.155672
R2060 VTAIL.n162 VTAIL.n161 0.155672
R2061 VTAIL.n162 VTAIL.n97 0.155672
R2062 VTAIL.n171 VTAIL.n97 0.155672
R2063 VTAIL.n172 VTAIL.n171 0.155672
R2064 VTAIL.n172 VTAIL.n93 0.155672
R2065 VTAIL.n179 VTAIL.n93 0.155672
R2066 VTAIL.n214 VTAIL.n209 0.155672
R2067 VTAIL.n221 VTAIL.n209 0.155672
R2068 VTAIL.n222 VTAIL.n221 0.155672
R2069 VTAIL.n222 VTAIL.n205 0.155672
R2070 VTAIL.n229 VTAIL.n205 0.155672
R2071 VTAIL.n230 VTAIL.n229 0.155672
R2072 VTAIL.n230 VTAIL.n201 0.155672
R2073 VTAIL.n237 VTAIL.n201 0.155672
R2074 VTAIL.n238 VTAIL.n237 0.155672
R2075 VTAIL.n238 VTAIL.n197 0.155672
R2076 VTAIL.n245 VTAIL.n197 0.155672
R2077 VTAIL.n246 VTAIL.n245 0.155672
R2078 VTAIL.n246 VTAIL.n193 0.155672
R2079 VTAIL.n253 VTAIL.n193 0.155672
R2080 VTAIL.n254 VTAIL.n253 0.155672
R2081 VTAIL.n254 VTAIL.n189 0.155672
R2082 VTAIL.n263 VTAIL.n189 0.155672
R2083 VTAIL.n264 VTAIL.n263 0.155672
R2084 VTAIL.n264 VTAIL.n185 0.155672
R2085 VTAIL.n271 VTAIL.n185 0.155672
R2086 VTAIL.n635 VTAIL.n549 0.155672
R2087 VTAIL.n628 VTAIL.n549 0.155672
R2088 VTAIL.n628 VTAIL.n627 0.155672
R2089 VTAIL.n627 VTAIL.n553 0.155672
R2090 VTAIL.n619 VTAIL.n553 0.155672
R2091 VTAIL.n619 VTAIL.n618 0.155672
R2092 VTAIL.n618 VTAIL.n558 0.155672
R2093 VTAIL.n611 VTAIL.n558 0.155672
R2094 VTAIL.n611 VTAIL.n610 0.155672
R2095 VTAIL.n610 VTAIL.n562 0.155672
R2096 VTAIL.n603 VTAIL.n562 0.155672
R2097 VTAIL.n603 VTAIL.n602 0.155672
R2098 VTAIL.n602 VTAIL.n566 0.155672
R2099 VTAIL.n595 VTAIL.n566 0.155672
R2100 VTAIL.n595 VTAIL.n594 0.155672
R2101 VTAIL.n594 VTAIL.n570 0.155672
R2102 VTAIL.n587 VTAIL.n570 0.155672
R2103 VTAIL.n587 VTAIL.n586 0.155672
R2104 VTAIL.n586 VTAIL.n574 0.155672
R2105 VTAIL.n579 VTAIL.n574 0.155672
R2106 VTAIL.n543 VTAIL.n457 0.155672
R2107 VTAIL.n536 VTAIL.n457 0.155672
R2108 VTAIL.n536 VTAIL.n535 0.155672
R2109 VTAIL.n535 VTAIL.n461 0.155672
R2110 VTAIL.n527 VTAIL.n461 0.155672
R2111 VTAIL.n527 VTAIL.n526 0.155672
R2112 VTAIL.n526 VTAIL.n466 0.155672
R2113 VTAIL.n519 VTAIL.n466 0.155672
R2114 VTAIL.n519 VTAIL.n518 0.155672
R2115 VTAIL.n518 VTAIL.n470 0.155672
R2116 VTAIL.n511 VTAIL.n470 0.155672
R2117 VTAIL.n511 VTAIL.n510 0.155672
R2118 VTAIL.n510 VTAIL.n474 0.155672
R2119 VTAIL.n503 VTAIL.n474 0.155672
R2120 VTAIL.n503 VTAIL.n502 0.155672
R2121 VTAIL.n502 VTAIL.n478 0.155672
R2122 VTAIL.n495 VTAIL.n478 0.155672
R2123 VTAIL.n495 VTAIL.n494 0.155672
R2124 VTAIL.n494 VTAIL.n482 0.155672
R2125 VTAIL.n487 VTAIL.n482 0.155672
R2126 VTAIL.n453 VTAIL.n367 0.155672
R2127 VTAIL.n446 VTAIL.n367 0.155672
R2128 VTAIL.n446 VTAIL.n445 0.155672
R2129 VTAIL.n445 VTAIL.n371 0.155672
R2130 VTAIL.n437 VTAIL.n371 0.155672
R2131 VTAIL.n437 VTAIL.n436 0.155672
R2132 VTAIL.n436 VTAIL.n376 0.155672
R2133 VTAIL.n429 VTAIL.n376 0.155672
R2134 VTAIL.n429 VTAIL.n428 0.155672
R2135 VTAIL.n428 VTAIL.n380 0.155672
R2136 VTAIL.n421 VTAIL.n380 0.155672
R2137 VTAIL.n421 VTAIL.n420 0.155672
R2138 VTAIL.n420 VTAIL.n384 0.155672
R2139 VTAIL.n413 VTAIL.n384 0.155672
R2140 VTAIL.n413 VTAIL.n412 0.155672
R2141 VTAIL.n412 VTAIL.n388 0.155672
R2142 VTAIL.n405 VTAIL.n388 0.155672
R2143 VTAIL.n405 VTAIL.n404 0.155672
R2144 VTAIL.n404 VTAIL.n392 0.155672
R2145 VTAIL.n397 VTAIL.n392 0.155672
R2146 VTAIL.n361 VTAIL.n275 0.155672
R2147 VTAIL.n354 VTAIL.n275 0.155672
R2148 VTAIL.n354 VTAIL.n353 0.155672
R2149 VTAIL.n353 VTAIL.n279 0.155672
R2150 VTAIL.n345 VTAIL.n279 0.155672
R2151 VTAIL.n345 VTAIL.n344 0.155672
R2152 VTAIL.n344 VTAIL.n284 0.155672
R2153 VTAIL.n337 VTAIL.n284 0.155672
R2154 VTAIL.n337 VTAIL.n336 0.155672
R2155 VTAIL.n336 VTAIL.n288 0.155672
R2156 VTAIL.n329 VTAIL.n288 0.155672
R2157 VTAIL.n329 VTAIL.n328 0.155672
R2158 VTAIL.n328 VTAIL.n292 0.155672
R2159 VTAIL.n321 VTAIL.n292 0.155672
R2160 VTAIL.n321 VTAIL.n320 0.155672
R2161 VTAIL.n320 VTAIL.n296 0.155672
R2162 VTAIL.n313 VTAIL.n296 0.155672
R2163 VTAIL.n313 VTAIL.n312 0.155672
R2164 VTAIL.n312 VTAIL.n300 0.155672
R2165 VTAIL.n305 VTAIL.n300 0.155672
R2166 VTAIL VTAIL.n1 0.0586897
R2167 VN.n3 VN.t2 605.996
R2168 VN.n13 VN.t4 605.996
R2169 VN.n2 VN.t0 582.692
R2170 VN.n6 VN.t3 582.692
R2171 VN.n8 VN.t1 582.692
R2172 VN.n12 VN.t6 582.692
R2173 VN.n16 VN.t5 582.692
R2174 VN.n18 VN.t7 582.692
R2175 VN.n9 VN.n8 161.3
R2176 VN.n19 VN.n18 161.3
R2177 VN.n17 VN.n10 161.3
R2178 VN.n16 VN.n15 161.3
R2179 VN.n14 VN.n11 161.3
R2180 VN.n7 VN.n0 161.3
R2181 VN.n6 VN.n5 161.3
R2182 VN.n4 VN.n1 161.3
R2183 VN VN.n19 45.6009
R2184 VN.n14 VN.n13 44.8907
R2185 VN.n4 VN.n3 44.8907
R2186 VN.n8 VN.n7 32.8641
R2187 VN.n18 VN.n17 32.8641
R2188 VN.n2 VN.n1 24.1005
R2189 VN.n6 VN.n1 24.1005
R2190 VN.n16 VN.n11 24.1005
R2191 VN.n12 VN.n11 24.1005
R2192 VN.n3 VN.n2 18.4104
R2193 VN.n13 VN.n12 18.4104
R2194 VN.n7 VN.n6 15.3369
R2195 VN.n17 VN.n16 15.3369
R2196 VN.n19 VN.n10 0.189894
R2197 VN.n15 VN.n10 0.189894
R2198 VN.n15 VN.n14 0.189894
R2199 VN.n5 VN.n4 0.189894
R2200 VN.n5 VN.n0 0.189894
R2201 VN.n9 VN.n0 0.189894
R2202 VN VN.n9 0.0516364
R2203 VDD2.n2 VDD2.n1 69.0399
R2204 VDD2.n2 VDD2.n0 69.0399
R2205 VDD2 VDD2.n5 69.037
R2206 VDD2.n4 VDD2.n3 68.6385
R2207 VDD2.n4 VDD2.n2 41.6377
R2208 VDD2.n5 VDD2.t1 2.02953
R2209 VDD2.n5 VDD2.t3 2.02953
R2210 VDD2.n3 VDD2.t0 2.02953
R2211 VDD2.n3 VDD2.t2 2.02953
R2212 VDD2.n1 VDD2.t4 2.02953
R2213 VDD2.n1 VDD2.t6 2.02953
R2214 VDD2.n0 VDD2.t5 2.02953
R2215 VDD2.n0 VDD2.t7 2.02953
R2216 VDD2 VDD2.n4 0.515586
C0 w_n2030_n4172# VDD1 1.4142f
C1 w_n2030_n4172# VDD2 1.45029f
C2 VDD1 VDD2 0.838674f
C3 B VTAIL 4.95454f
C4 VP VTAIL 7.01596f
C5 VN VTAIL 7.00185f
C6 B VP 1.26043f
C7 B VN 0.837859f
C8 VP VN 6.11606f
C9 w_n2030_n4172# VTAIL 5.20898f
C10 w_n2030_n4172# B 8.38118f
C11 VTAIL VDD1 13.7987f
C12 B VDD1 1.18748f
C13 w_n2030_n4172# VP 3.94091f
C14 w_n2030_n4172# VN 3.68288f
C15 VTAIL VDD2 13.8406f
C16 B VDD2 1.22507f
C17 VP VDD1 7.56314f
C18 VN VDD1 0.148335f
C19 VP VDD2 0.320671f
C20 VN VDD2 7.39126f
C21 VDD2 VSUBS 1.46088f
C22 VDD1 VSUBS 1.77458f
C23 VTAIL VSUBS 1.086827f
C24 VN VSUBS 5.00276f
C25 VP VSUBS 1.823913f
C26 B VSUBS 3.260284f
C27 w_n2030_n4172# VSUBS 0.103749p
C28 VDD2.t5 VSUBS 0.344842f
C29 VDD2.t7 VSUBS 0.344842f
C30 VDD2.n0 VSUBS 2.82043f
C31 VDD2.t4 VSUBS 0.344842f
C32 VDD2.t6 VSUBS 0.344842f
C33 VDD2.n1 VSUBS 2.82043f
C34 VDD2.n2 VSUBS 3.27307f
C35 VDD2.t0 VSUBS 0.344842f
C36 VDD2.t2 VSUBS 0.344842f
C37 VDD2.n3 VSUBS 2.81659f
C38 VDD2.n4 VSUBS 3.15383f
C39 VDD2.t1 VSUBS 0.344842f
C40 VDD2.t3 VSUBS 0.344842f
C41 VDD2.n5 VSUBS 2.82039f
C42 VN.n0 VSUBS 0.050831f
C43 VN.n1 VSUBS 0.011534f
C44 VN.t2 VSUBS 1.71256f
C45 VN.t0 VSUBS 1.68775f
C46 VN.n2 VSUBS 0.650022f
C47 VN.n3 VSUBS 0.62503f
C48 VN.n4 VSUBS 0.215106f
C49 VN.n5 VSUBS 0.050831f
C50 VN.t3 VSUBS 1.68775f
C51 VN.n6 VSUBS 0.644337f
C52 VN.n7 VSUBS 0.011534f
C53 VN.t1 VSUBS 1.68775f
C54 VN.n8 VSUBS 0.642927f
C55 VN.n9 VSUBS 0.039392f
C56 VN.n10 VSUBS 0.050831f
C57 VN.n11 VSUBS 0.011534f
C58 VN.t5 VSUBS 1.68775f
C59 VN.t4 VSUBS 1.71256f
C60 VN.t6 VSUBS 1.68775f
C61 VN.n12 VSUBS 0.650022f
C62 VN.n13 VSUBS 0.62503f
C63 VN.n14 VSUBS 0.215106f
C64 VN.n15 VSUBS 0.050831f
C65 VN.n16 VSUBS 0.644337f
C66 VN.n17 VSUBS 0.011534f
C67 VN.t7 VSUBS 1.68775f
C68 VN.n18 VSUBS 0.642927f
C69 VN.n19 VSUBS 2.39927f
C70 VTAIL.t2 VSUBS 0.307224f
C71 VTAIL.t3 VSUBS 0.307224f
C72 VTAIL.n0 VSUBS 2.35811f
C73 VTAIL.n1 VSUBS 0.669956f
C74 VTAIL.n2 VSUBS 0.024712f
C75 VTAIL.n3 VSUBS 0.024268f
C76 VTAIL.n4 VSUBS 0.013041f
C77 VTAIL.n5 VSUBS 0.030824f
C78 VTAIL.n6 VSUBS 0.013808f
C79 VTAIL.n7 VSUBS 0.024268f
C80 VTAIL.n8 VSUBS 0.013424f
C81 VTAIL.n9 VSUBS 0.030824f
C82 VTAIL.n10 VSUBS 0.013808f
C83 VTAIL.n11 VSUBS 0.024268f
C84 VTAIL.n12 VSUBS 0.013041f
C85 VTAIL.n13 VSUBS 0.030824f
C86 VTAIL.n14 VSUBS 0.013808f
C87 VTAIL.n15 VSUBS 0.024268f
C88 VTAIL.n16 VSUBS 0.013041f
C89 VTAIL.n17 VSUBS 0.030824f
C90 VTAIL.n18 VSUBS 0.013808f
C91 VTAIL.n19 VSUBS 0.024268f
C92 VTAIL.n20 VSUBS 0.013041f
C93 VTAIL.n21 VSUBS 0.030824f
C94 VTAIL.n22 VSUBS 0.013808f
C95 VTAIL.n23 VSUBS 0.024268f
C96 VTAIL.n24 VSUBS 0.013041f
C97 VTAIL.n25 VSUBS 0.030824f
C98 VTAIL.n26 VSUBS 0.013808f
C99 VTAIL.n27 VSUBS 0.024268f
C100 VTAIL.n28 VSUBS 0.013041f
C101 VTAIL.n29 VSUBS 0.023118f
C102 VTAIL.n30 VSUBS 0.019608f
C103 VTAIL.t4 VSUBS 0.066048f
C104 VTAIL.n31 VSUBS 0.178372f
C105 VTAIL.n32 VSUBS 1.66196f
C106 VTAIL.n33 VSUBS 0.013041f
C107 VTAIL.n34 VSUBS 0.013808f
C108 VTAIL.n35 VSUBS 0.030824f
C109 VTAIL.n36 VSUBS 0.030824f
C110 VTAIL.n37 VSUBS 0.013808f
C111 VTAIL.n38 VSUBS 0.013041f
C112 VTAIL.n39 VSUBS 0.024268f
C113 VTAIL.n40 VSUBS 0.024268f
C114 VTAIL.n41 VSUBS 0.013041f
C115 VTAIL.n42 VSUBS 0.013808f
C116 VTAIL.n43 VSUBS 0.030824f
C117 VTAIL.n44 VSUBS 0.030824f
C118 VTAIL.n45 VSUBS 0.013808f
C119 VTAIL.n46 VSUBS 0.013041f
C120 VTAIL.n47 VSUBS 0.024268f
C121 VTAIL.n48 VSUBS 0.024268f
C122 VTAIL.n49 VSUBS 0.013041f
C123 VTAIL.n50 VSUBS 0.013808f
C124 VTAIL.n51 VSUBS 0.030824f
C125 VTAIL.n52 VSUBS 0.030824f
C126 VTAIL.n53 VSUBS 0.013808f
C127 VTAIL.n54 VSUBS 0.013041f
C128 VTAIL.n55 VSUBS 0.024268f
C129 VTAIL.n56 VSUBS 0.024268f
C130 VTAIL.n57 VSUBS 0.013041f
C131 VTAIL.n58 VSUBS 0.013808f
C132 VTAIL.n59 VSUBS 0.030824f
C133 VTAIL.n60 VSUBS 0.030824f
C134 VTAIL.n61 VSUBS 0.013808f
C135 VTAIL.n62 VSUBS 0.013041f
C136 VTAIL.n63 VSUBS 0.024268f
C137 VTAIL.n64 VSUBS 0.024268f
C138 VTAIL.n65 VSUBS 0.013041f
C139 VTAIL.n66 VSUBS 0.013808f
C140 VTAIL.n67 VSUBS 0.030824f
C141 VTAIL.n68 VSUBS 0.030824f
C142 VTAIL.n69 VSUBS 0.013808f
C143 VTAIL.n70 VSUBS 0.013041f
C144 VTAIL.n71 VSUBS 0.024268f
C145 VTAIL.n72 VSUBS 0.024268f
C146 VTAIL.n73 VSUBS 0.013041f
C147 VTAIL.n74 VSUBS 0.013041f
C148 VTAIL.n75 VSUBS 0.013808f
C149 VTAIL.n76 VSUBS 0.030824f
C150 VTAIL.n77 VSUBS 0.030824f
C151 VTAIL.n78 VSUBS 0.030824f
C152 VTAIL.n79 VSUBS 0.013424f
C153 VTAIL.n80 VSUBS 0.013041f
C154 VTAIL.n81 VSUBS 0.024268f
C155 VTAIL.n82 VSUBS 0.024268f
C156 VTAIL.n83 VSUBS 0.013041f
C157 VTAIL.n84 VSUBS 0.013808f
C158 VTAIL.n85 VSUBS 0.030824f
C159 VTAIL.n86 VSUBS 0.067967f
C160 VTAIL.n87 VSUBS 0.013808f
C161 VTAIL.n88 VSUBS 0.013041f
C162 VTAIL.n89 VSUBS 0.054106f
C163 VTAIL.n90 VSUBS 0.033823f
C164 VTAIL.n91 VSUBS 0.127801f
C165 VTAIL.n92 VSUBS 0.024712f
C166 VTAIL.n93 VSUBS 0.024268f
C167 VTAIL.n94 VSUBS 0.013041f
C168 VTAIL.n95 VSUBS 0.030824f
C169 VTAIL.n96 VSUBS 0.013808f
C170 VTAIL.n97 VSUBS 0.024268f
C171 VTAIL.n98 VSUBS 0.013424f
C172 VTAIL.n99 VSUBS 0.030824f
C173 VTAIL.n100 VSUBS 0.013808f
C174 VTAIL.n101 VSUBS 0.024268f
C175 VTAIL.n102 VSUBS 0.013041f
C176 VTAIL.n103 VSUBS 0.030824f
C177 VTAIL.n104 VSUBS 0.013808f
C178 VTAIL.n105 VSUBS 0.024268f
C179 VTAIL.n106 VSUBS 0.013041f
C180 VTAIL.n107 VSUBS 0.030824f
C181 VTAIL.n108 VSUBS 0.013808f
C182 VTAIL.n109 VSUBS 0.024268f
C183 VTAIL.n110 VSUBS 0.013041f
C184 VTAIL.n111 VSUBS 0.030824f
C185 VTAIL.n112 VSUBS 0.013808f
C186 VTAIL.n113 VSUBS 0.024268f
C187 VTAIL.n114 VSUBS 0.013041f
C188 VTAIL.n115 VSUBS 0.030824f
C189 VTAIL.n116 VSUBS 0.013808f
C190 VTAIL.n117 VSUBS 0.024268f
C191 VTAIL.n118 VSUBS 0.013041f
C192 VTAIL.n119 VSUBS 0.023118f
C193 VTAIL.n120 VSUBS 0.019608f
C194 VTAIL.t8 VSUBS 0.066048f
C195 VTAIL.n121 VSUBS 0.178372f
C196 VTAIL.n122 VSUBS 1.66196f
C197 VTAIL.n123 VSUBS 0.013041f
C198 VTAIL.n124 VSUBS 0.013808f
C199 VTAIL.n125 VSUBS 0.030824f
C200 VTAIL.n126 VSUBS 0.030824f
C201 VTAIL.n127 VSUBS 0.013808f
C202 VTAIL.n128 VSUBS 0.013041f
C203 VTAIL.n129 VSUBS 0.024268f
C204 VTAIL.n130 VSUBS 0.024268f
C205 VTAIL.n131 VSUBS 0.013041f
C206 VTAIL.n132 VSUBS 0.013808f
C207 VTAIL.n133 VSUBS 0.030824f
C208 VTAIL.n134 VSUBS 0.030824f
C209 VTAIL.n135 VSUBS 0.013808f
C210 VTAIL.n136 VSUBS 0.013041f
C211 VTAIL.n137 VSUBS 0.024268f
C212 VTAIL.n138 VSUBS 0.024268f
C213 VTAIL.n139 VSUBS 0.013041f
C214 VTAIL.n140 VSUBS 0.013808f
C215 VTAIL.n141 VSUBS 0.030824f
C216 VTAIL.n142 VSUBS 0.030824f
C217 VTAIL.n143 VSUBS 0.013808f
C218 VTAIL.n144 VSUBS 0.013041f
C219 VTAIL.n145 VSUBS 0.024268f
C220 VTAIL.n146 VSUBS 0.024268f
C221 VTAIL.n147 VSUBS 0.013041f
C222 VTAIL.n148 VSUBS 0.013808f
C223 VTAIL.n149 VSUBS 0.030824f
C224 VTAIL.n150 VSUBS 0.030824f
C225 VTAIL.n151 VSUBS 0.013808f
C226 VTAIL.n152 VSUBS 0.013041f
C227 VTAIL.n153 VSUBS 0.024268f
C228 VTAIL.n154 VSUBS 0.024268f
C229 VTAIL.n155 VSUBS 0.013041f
C230 VTAIL.n156 VSUBS 0.013808f
C231 VTAIL.n157 VSUBS 0.030824f
C232 VTAIL.n158 VSUBS 0.030824f
C233 VTAIL.n159 VSUBS 0.013808f
C234 VTAIL.n160 VSUBS 0.013041f
C235 VTAIL.n161 VSUBS 0.024268f
C236 VTAIL.n162 VSUBS 0.024268f
C237 VTAIL.n163 VSUBS 0.013041f
C238 VTAIL.n164 VSUBS 0.013041f
C239 VTAIL.n165 VSUBS 0.013808f
C240 VTAIL.n166 VSUBS 0.030824f
C241 VTAIL.n167 VSUBS 0.030824f
C242 VTAIL.n168 VSUBS 0.030824f
C243 VTAIL.n169 VSUBS 0.013424f
C244 VTAIL.n170 VSUBS 0.013041f
C245 VTAIL.n171 VSUBS 0.024268f
C246 VTAIL.n172 VSUBS 0.024268f
C247 VTAIL.n173 VSUBS 0.013041f
C248 VTAIL.n174 VSUBS 0.013808f
C249 VTAIL.n175 VSUBS 0.030824f
C250 VTAIL.n176 VSUBS 0.067967f
C251 VTAIL.n177 VSUBS 0.013808f
C252 VTAIL.n178 VSUBS 0.013041f
C253 VTAIL.n179 VSUBS 0.054106f
C254 VTAIL.n180 VSUBS 0.033823f
C255 VTAIL.n181 VSUBS 0.127801f
C256 VTAIL.t11 VSUBS 0.307224f
C257 VTAIL.t9 VSUBS 0.307224f
C258 VTAIL.n182 VSUBS 2.35811f
C259 VTAIL.n183 VSUBS 0.736862f
C260 VTAIL.n184 VSUBS 0.024712f
C261 VTAIL.n185 VSUBS 0.024268f
C262 VTAIL.n186 VSUBS 0.013041f
C263 VTAIL.n187 VSUBS 0.030824f
C264 VTAIL.n188 VSUBS 0.013808f
C265 VTAIL.n189 VSUBS 0.024268f
C266 VTAIL.n190 VSUBS 0.013424f
C267 VTAIL.n191 VSUBS 0.030824f
C268 VTAIL.n192 VSUBS 0.013808f
C269 VTAIL.n193 VSUBS 0.024268f
C270 VTAIL.n194 VSUBS 0.013041f
C271 VTAIL.n195 VSUBS 0.030824f
C272 VTAIL.n196 VSUBS 0.013808f
C273 VTAIL.n197 VSUBS 0.024268f
C274 VTAIL.n198 VSUBS 0.013041f
C275 VTAIL.n199 VSUBS 0.030824f
C276 VTAIL.n200 VSUBS 0.013808f
C277 VTAIL.n201 VSUBS 0.024268f
C278 VTAIL.n202 VSUBS 0.013041f
C279 VTAIL.n203 VSUBS 0.030824f
C280 VTAIL.n204 VSUBS 0.013808f
C281 VTAIL.n205 VSUBS 0.024268f
C282 VTAIL.n206 VSUBS 0.013041f
C283 VTAIL.n207 VSUBS 0.030824f
C284 VTAIL.n208 VSUBS 0.013808f
C285 VTAIL.n209 VSUBS 0.024268f
C286 VTAIL.n210 VSUBS 0.013041f
C287 VTAIL.n211 VSUBS 0.023118f
C288 VTAIL.n212 VSUBS 0.019608f
C289 VTAIL.t10 VSUBS 0.066048f
C290 VTAIL.n213 VSUBS 0.178372f
C291 VTAIL.n214 VSUBS 1.66196f
C292 VTAIL.n215 VSUBS 0.013041f
C293 VTAIL.n216 VSUBS 0.013808f
C294 VTAIL.n217 VSUBS 0.030824f
C295 VTAIL.n218 VSUBS 0.030824f
C296 VTAIL.n219 VSUBS 0.013808f
C297 VTAIL.n220 VSUBS 0.013041f
C298 VTAIL.n221 VSUBS 0.024268f
C299 VTAIL.n222 VSUBS 0.024268f
C300 VTAIL.n223 VSUBS 0.013041f
C301 VTAIL.n224 VSUBS 0.013808f
C302 VTAIL.n225 VSUBS 0.030824f
C303 VTAIL.n226 VSUBS 0.030824f
C304 VTAIL.n227 VSUBS 0.013808f
C305 VTAIL.n228 VSUBS 0.013041f
C306 VTAIL.n229 VSUBS 0.024268f
C307 VTAIL.n230 VSUBS 0.024268f
C308 VTAIL.n231 VSUBS 0.013041f
C309 VTAIL.n232 VSUBS 0.013808f
C310 VTAIL.n233 VSUBS 0.030824f
C311 VTAIL.n234 VSUBS 0.030824f
C312 VTAIL.n235 VSUBS 0.013808f
C313 VTAIL.n236 VSUBS 0.013041f
C314 VTAIL.n237 VSUBS 0.024268f
C315 VTAIL.n238 VSUBS 0.024268f
C316 VTAIL.n239 VSUBS 0.013041f
C317 VTAIL.n240 VSUBS 0.013808f
C318 VTAIL.n241 VSUBS 0.030824f
C319 VTAIL.n242 VSUBS 0.030824f
C320 VTAIL.n243 VSUBS 0.013808f
C321 VTAIL.n244 VSUBS 0.013041f
C322 VTAIL.n245 VSUBS 0.024268f
C323 VTAIL.n246 VSUBS 0.024268f
C324 VTAIL.n247 VSUBS 0.013041f
C325 VTAIL.n248 VSUBS 0.013808f
C326 VTAIL.n249 VSUBS 0.030824f
C327 VTAIL.n250 VSUBS 0.030824f
C328 VTAIL.n251 VSUBS 0.013808f
C329 VTAIL.n252 VSUBS 0.013041f
C330 VTAIL.n253 VSUBS 0.024268f
C331 VTAIL.n254 VSUBS 0.024268f
C332 VTAIL.n255 VSUBS 0.013041f
C333 VTAIL.n256 VSUBS 0.013041f
C334 VTAIL.n257 VSUBS 0.013808f
C335 VTAIL.n258 VSUBS 0.030824f
C336 VTAIL.n259 VSUBS 0.030824f
C337 VTAIL.n260 VSUBS 0.030824f
C338 VTAIL.n261 VSUBS 0.013424f
C339 VTAIL.n262 VSUBS 0.013041f
C340 VTAIL.n263 VSUBS 0.024268f
C341 VTAIL.n264 VSUBS 0.024268f
C342 VTAIL.n265 VSUBS 0.013041f
C343 VTAIL.n266 VSUBS 0.013808f
C344 VTAIL.n267 VSUBS 0.030824f
C345 VTAIL.n268 VSUBS 0.067967f
C346 VTAIL.n269 VSUBS 0.013808f
C347 VTAIL.n270 VSUBS 0.013041f
C348 VTAIL.n271 VSUBS 0.054106f
C349 VTAIL.n272 VSUBS 0.033823f
C350 VTAIL.n273 VSUBS 1.57212f
C351 VTAIL.n274 VSUBS 0.024712f
C352 VTAIL.n275 VSUBS 0.024268f
C353 VTAIL.n276 VSUBS 0.013041f
C354 VTAIL.n277 VSUBS 0.030824f
C355 VTAIL.n278 VSUBS 0.013808f
C356 VTAIL.n279 VSUBS 0.024268f
C357 VTAIL.n280 VSUBS 0.013424f
C358 VTAIL.n281 VSUBS 0.030824f
C359 VTAIL.n282 VSUBS 0.013041f
C360 VTAIL.n283 VSUBS 0.013808f
C361 VTAIL.n284 VSUBS 0.024268f
C362 VTAIL.n285 VSUBS 0.013041f
C363 VTAIL.n286 VSUBS 0.030824f
C364 VTAIL.n287 VSUBS 0.013808f
C365 VTAIL.n288 VSUBS 0.024268f
C366 VTAIL.n289 VSUBS 0.013041f
C367 VTAIL.n290 VSUBS 0.030824f
C368 VTAIL.n291 VSUBS 0.013808f
C369 VTAIL.n292 VSUBS 0.024268f
C370 VTAIL.n293 VSUBS 0.013041f
C371 VTAIL.n294 VSUBS 0.030824f
C372 VTAIL.n295 VSUBS 0.013808f
C373 VTAIL.n296 VSUBS 0.024268f
C374 VTAIL.n297 VSUBS 0.013041f
C375 VTAIL.n298 VSUBS 0.030824f
C376 VTAIL.n299 VSUBS 0.013808f
C377 VTAIL.n300 VSUBS 0.024268f
C378 VTAIL.n301 VSUBS 0.013041f
C379 VTAIL.n302 VSUBS 0.023118f
C380 VTAIL.n303 VSUBS 0.019608f
C381 VTAIL.t15 VSUBS 0.066048f
C382 VTAIL.n304 VSUBS 0.178372f
C383 VTAIL.n305 VSUBS 1.66196f
C384 VTAIL.n306 VSUBS 0.013041f
C385 VTAIL.n307 VSUBS 0.013808f
C386 VTAIL.n308 VSUBS 0.030824f
C387 VTAIL.n309 VSUBS 0.030824f
C388 VTAIL.n310 VSUBS 0.013808f
C389 VTAIL.n311 VSUBS 0.013041f
C390 VTAIL.n312 VSUBS 0.024268f
C391 VTAIL.n313 VSUBS 0.024268f
C392 VTAIL.n314 VSUBS 0.013041f
C393 VTAIL.n315 VSUBS 0.013808f
C394 VTAIL.n316 VSUBS 0.030824f
C395 VTAIL.n317 VSUBS 0.030824f
C396 VTAIL.n318 VSUBS 0.013808f
C397 VTAIL.n319 VSUBS 0.013041f
C398 VTAIL.n320 VSUBS 0.024268f
C399 VTAIL.n321 VSUBS 0.024268f
C400 VTAIL.n322 VSUBS 0.013041f
C401 VTAIL.n323 VSUBS 0.013808f
C402 VTAIL.n324 VSUBS 0.030824f
C403 VTAIL.n325 VSUBS 0.030824f
C404 VTAIL.n326 VSUBS 0.013808f
C405 VTAIL.n327 VSUBS 0.013041f
C406 VTAIL.n328 VSUBS 0.024268f
C407 VTAIL.n329 VSUBS 0.024268f
C408 VTAIL.n330 VSUBS 0.013041f
C409 VTAIL.n331 VSUBS 0.013808f
C410 VTAIL.n332 VSUBS 0.030824f
C411 VTAIL.n333 VSUBS 0.030824f
C412 VTAIL.n334 VSUBS 0.013808f
C413 VTAIL.n335 VSUBS 0.013041f
C414 VTAIL.n336 VSUBS 0.024268f
C415 VTAIL.n337 VSUBS 0.024268f
C416 VTAIL.n338 VSUBS 0.013041f
C417 VTAIL.n339 VSUBS 0.013808f
C418 VTAIL.n340 VSUBS 0.030824f
C419 VTAIL.n341 VSUBS 0.030824f
C420 VTAIL.n342 VSUBS 0.013808f
C421 VTAIL.n343 VSUBS 0.013041f
C422 VTAIL.n344 VSUBS 0.024268f
C423 VTAIL.n345 VSUBS 0.024268f
C424 VTAIL.n346 VSUBS 0.013041f
C425 VTAIL.n347 VSUBS 0.013808f
C426 VTAIL.n348 VSUBS 0.030824f
C427 VTAIL.n349 VSUBS 0.030824f
C428 VTAIL.n350 VSUBS 0.030824f
C429 VTAIL.n351 VSUBS 0.013424f
C430 VTAIL.n352 VSUBS 0.013041f
C431 VTAIL.n353 VSUBS 0.024268f
C432 VTAIL.n354 VSUBS 0.024268f
C433 VTAIL.n355 VSUBS 0.013041f
C434 VTAIL.n356 VSUBS 0.013808f
C435 VTAIL.n357 VSUBS 0.030824f
C436 VTAIL.n358 VSUBS 0.067967f
C437 VTAIL.n359 VSUBS 0.013808f
C438 VTAIL.n360 VSUBS 0.013041f
C439 VTAIL.n361 VSUBS 0.054106f
C440 VTAIL.n362 VSUBS 0.033823f
C441 VTAIL.n363 VSUBS 1.57212f
C442 VTAIL.t1 VSUBS 0.307224f
C443 VTAIL.t6 VSUBS 0.307224f
C444 VTAIL.n364 VSUBS 2.35812f
C445 VTAIL.n365 VSUBS 0.736847f
C446 VTAIL.n366 VSUBS 0.024712f
C447 VTAIL.n367 VSUBS 0.024268f
C448 VTAIL.n368 VSUBS 0.013041f
C449 VTAIL.n369 VSUBS 0.030824f
C450 VTAIL.n370 VSUBS 0.013808f
C451 VTAIL.n371 VSUBS 0.024268f
C452 VTAIL.n372 VSUBS 0.013424f
C453 VTAIL.n373 VSUBS 0.030824f
C454 VTAIL.n374 VSUBS 0.013041f
C455 VTAIL.n375 VSUBS 0.013808f
C456 VTAIL.n376 VSUBS 0.024268f
C457 VTAIL.n377 VSUBS 0.013041f
C458 VTAIL.n378 VSUBS 0.030824f
C459 VTAIL.n379 VSUBS 0.013808f
C460 VTAIL.n380 VSUBS 0.024268f
C461 VTAIL.n381 VSUBS 0.013041f
C462 VTAIL.n382 VSUBS 0.030824f
C463 VTAIL.n383 VSUBS 0.013808f
C464 VTAIL.n384 VSUBS 0.024268f
C465 VTAIL.n385 VSUBS 0.013041f
C466 VTAIL.n386 VSUBS 0.030824f
C467 VTAIL.n387 VSUBS 0.013808f
C468 VTAIL.n388 VSUBS 0.024268f
C469 VTAIL.n389 VSUBS 0.013041f
C470 VTAIL.n390 VSUBS 0.030824f
C471 VTAIL.n391 VSUBS 0.013808f
C472 VTAIL.n392 VSUBS 0.024268f
C473 VTAIL.n393 VSUBS 0.013041f
C474 VTAIL.n394 VSUBS 0.023118f
C475 VTAIL.n395 VSUBS 0.019608f
C476 VTAIL.t0 VSUBS 0.066048f
C477 VTAIL.n396 VSUBS 0.178372f
C478 VTAIL.n397 VSUBS 1.66196f
C479 VTAIL.n398 VSUBS 0.013041f
C480 VTAIL.n399 VSUBS 0.013808f
C481 VTAIL.n400 VSUBS 0.030824f
C482 VTAIL.n401 VSUBS 0.030824f
C483 VTAIL.n402 VSUBS 0.013808f
C484 VTAIL.n403 VSUBS 0.013041f
C485 VTAIL.n404 VSUBS 0.024268f
C486 VTAIL.n405 VSUBS 0.024268f
C487 VTAIL.n406 VSUBS 0.013041f
C488 VTAIL.n407 VSUBS 0.013808f
C489 VTAIL.n408 VSUBS 0.030824f
C490 VTAIL.n409 VSUBS 0.030824f
C491 VTAIL.n410 VSUBS 0.013808f
C492 VTAIL.n411 VSUBS 0.013041f
C493 VTAIL.n412 VSUBS 0.024268f
C494 VTAIL.n413 VSUBS 0.024268f
C495 VTAIL.n414 VSUBS 0.013041f
C496 VTAIL.n415 VSUBS 0.013808f
C497 VTAIL.n416 VSUBS 0.030824f
C498 VTAIL.n417 VSUBS 0.030824f
C499 VTAIL.n418 VSUBS 0.013808f
C500 VTAIL.n419 VSUBS 0.013041f
C501 VTAIL.n420 VSUBS 0.024268f
C502 VTAIL.n421 VSUBS 0.024268f
C503 VTAIL.n422 VSUBS 0.013041f
C504 VTAIL.n423 VSUBS 0.013808f
C505 VTAIL.n424 VSUBS 0.030824f
C506 VTAIL.n425 VSUBS 0.030824f
C507 VTAIL.n426 VSUBS 0.013808f
C508 VTAIL.n427 VSUBS 0.013041f
C509 VTAIL.n428 VSUBS 0.024268f
C510 VTAIL.n429 VSUBS 0.024268f
C511 VTAIL.n430 VSUBS 0.013041f
C512 VTAIL.n431 VSUBS 0.013808f
C513 VTAIL.n432 VSUBS 0.030824f
C514 VTAIL.n433 VSUBS 0.030824f
C515 VTAIL.n434 VSUBS 0.013808f
C516 VTAIL.n435 VSUBS 0.013041f
C517 VTAIL.n436 VSUBS 0.024268f
C518 VTAIL.n437 VSUBS 0.024268f
C519 VTAIL.n438 VSUBS 0.013041f
C520 VTAIL.n439 VSUBS 0.013808f
C521 VTAIL.n440 VSUBS 0.030824f
C522 VTAIL.n441 VSUBS 0.030824f
C523 VTAIL.n442 VSUBS 0.030824f
C524 VTAIL.n443 VSUBS 0.013424f
C525 VTAIL.n444 VSUBS 0.013041f
C526 VTAIL.n445 VSUBS 0.024268f
C527 VTAIL.n446 VSUBS 0.024268f
C528 VTAIL.n447 VSUBS 0.013041f
C529 VTAIL.n448 VSUBS 0.013808f
C530 VTAIL.n449 VSUBS 0.030824f
C531 VTAIL.n450 VSUBS 0.067967f
C532 VTAIL.n451 VSUBS 0.013808f
C533 VTAIL.n452 VSUBS 0.013041f
C534 VTAIL.n453 VSUBS 0.054106f
C535 VTAIL.n454 VSUBS 0.033823f
C536 VTAIL.n455 VSUBS 0.127801f
C537 VTAIL.n456 VSUBS 0.024712f
C538 VTAIL.n457 VSUBS 0.024268f
C539 VTAIL.n458 VSUBS 0.013041f
C540 VTAIL.n459 VSUBS 0.030824f
C541 VTAIL.n460 VSUBS 0.013808f
C542 VTAIL.n461 VSUBS 0.024268f
C543 VTAIL.n462 VSUBS 0.013424f
C544 VTAIL.n463 VSUBS 0.030824f
C545 VTAIL.n464 VSUBS 0.013041f
C546 VTAIL.n465 VSUBS 0.013808f
C547 VTAIL.n466 VSUBS 0.024268f
C548 VTAIL.n467 VSUBS 0.013041f
C549 VTAIL.n468 VSUBS 0.030824f
C550 VTAIL.n469 VSUBS 0.013808f
C551 VTAIL.n470 VSUBS 0.024268f
C552 VTAIL.n471 VSUBS 0.013041f
C553 VTAIL.n472 VSUBS 0.030824f
C554 VTAIL.n473 VSUBS 0.013808f
C555 VTAIL.n474 VSUBS 0.024268f
C556 VTAIL.n475 VSUBS 0.013041f
C557 VTAIL.n476 VSUBS 0.030824f
C558 VTAIL.n477 VSUBS 0.013808f
C559 VTAIL.n478 VSUBS 0.024268f
C560 VTAIL.n479 VSUBS 0.013041f
C561 VTAIL.n480 VSUBS 0.030824f
C562 VTAIL.n481 VSUBS 0.013808f
C563 VTAIL.n482 VSUBS 0.024268f
C564 VTAIL.n483 VSUBS 0.013041f
C565 VTAIL.n484 VSUBS 0.023118f
C566 VTAIL.n485 VSUBS 0.019608f
C567 VTAIL.t14 VSUBS 0.066048f
C568 VTAIL.n486 VSUBS 0.178372f
C569 VTAIL.n487 VSUBS 1.66196f
C570 VTAIL.n488 VSUBS 0.013041f
C571 VTAIL.n489 VSUBS 0.013808f
C572 VTAIL.n490 VSUBS 0.030824f
C573 VTAIL.n491 VSUBS 0.030824f
C574 VTAIL.n492 VSUBS 0.013808f
C575 VTAIL.n493 VSUBS 0.013041f
C576 VTAIL.n494 VSUBS 0.024268f
C577 VTAIL.n495 VSUBS 0.024268f
C578 VTAIL.n496 VSUBS 0.013041f
C579 VTAIL.n497 VSUBS 0.013808f
C580 VTAIL.n498 VSUBS 0.030824f
C581 VTAIL.n499 VSUBS 0.030824f
C582 VTAIL.n500 VSUBS 0.013808f
C583 VTAIL.n501 VSUBS 0.013041f
C584 VTAIL.n502 VSUBS 0.024268f
C585 VTAIL.n503 VSUBS 0.024268f
C586 VTAIL.n504 VSUBS 0.013041f
C587 VTAIL.n505 VSUBS 0.013808f
C588 VTAIL.n506 VSUBS 0.030824f
C589 VTAIL.n507 VSUBS 0.030824f
C590 VTAIL.n508 VSUBS 0.013808f
C591 VTAIL.n509 VSUBS 0.013041f
C592 VTAIL.n510 VSUBS 0.024268f
C593 VTAIL.n511 VSUBS 0.024268f
C594 VTAIL.n512 VSUBS 0.013041f
C595 VTAIL.n513 VSUBS 0.013808f
C596 VTAIL.n514 VSUBS 0.030824f
C597 VTAIL.n515 VSUBS 0.030824f
C598 VTAIL.n516 VSUBS 0.013808f
C599 VTAIL.n517 VSUBS 0.013041f
C600 VTAIL.n518 VSUBS 0.024268f
C601 VTAIL.n519 VSUBS 0.024268f
C602 VTAIL.n520 VSUBS 0.013041f
C603 VTAIL.n521 VSUBS 0.013808f
C604 VTAIL.n522 VSUBS 0.030824f
C605 VTAIL.n523 VSUBS 0.030824f
C606 VTAIL.n524 VSUBS 0.013808f
C607 VTAIL.n525 VSUBS 0.013041f
C608 VTAIL.n526 VSUBS 0.024268f
C609 VTAIL.n527 VSUBS 0.024268f
C610 VTAIL.n528 VSUBS 0.013041f
C611 VTAIL.n529 VSUBS 0.013808f
C612 VTAIL.n530 VSUBS 0.030824f
C613 VTAIL.n531 VSUBS 0.030824f
C614 VTAIL.n532 VSUBS 0.030824f
C615 VTAIL.n533 VSUBS 0.013424f
C616 VTAIL.n534 VSUBS 0.013041f
C617 VTAIL.n535 VSUBS 0.024268f
C618 VTAIL.n536 VSUBS 0.024268f
C619 VTAIL.n537 VSUBS 0.013041f
C620 VTAIL.n538 VSUBS 0.013808f
C621 VTAIL.n539 VSUBS 0.030824f
C622 VTAIL.n540 VSUBS 0.067967f
C623 VTAIL.n541 VSUBS 0.013808f
C624 VTAIL.n542 VSUBS 0.013041f
C625 VTAIL.n543 VSUBS 0.054106f
C626 VTAIL.n544 VSUBS 0.033823f
C627 VTAIL.n545 VSUBS 0.127801f
C628 VTAIL.t12 VSUBS 0.307224f
C629 VTAIL.t13 VSUBS 0.307224f
C630 VTAIL.n546 VSUBS 2.35812f
C631 VTAIL.n547 VSUBS 0.736847f
C632 VTAIL.n548 VSUBS 0.024712f
C633 VTAIL.n549 VSUBS 0.024268f
C634 VTAIL.n550 VSUBS 0.013041f
C635 VTAIL.n551 VSUBS 0.030824f
C636 VTAIL.n552 VSUBS 0.013808f
C637 VTAIL.n553 VSUBS 0.024268f
C638 VTAIL.n554 VSUBS 0.013424f
C639 VTAIL.n555 VSUBS 0.030824f
C640 VTAIL.n556 VSUBS 0.013041f
C641 VTAIL.n557 VSUBS 0.013808f
C642 VTAIL.n558 VSUBS 0.024268f
C643 VTAIL.n559 VSUBS 0.013041f
C644 VTAIL.n560 VSUBS 0.030824f
C645 VTAIL.n561 VSUBS 0.013808f
C646 VTAIL.n562 VSUBS 0.024268f
C647 VTAIL.n563 VSUBS 0.013041f
C648 VTAIL.n564 VSUBS 0.030824f
C649 VTAIL.n565 VSUBS 0.013808f
C650 VTAIL.n566 VSUBS 0.024268f
C651 VTAIL.n567 VSUBS 0.013041f
C652 VTAIL.n568 VSUBS 0.030824f
C653 VTAIL.n569 VSUBS 0.013808f
C654 VTAIL.n570 VSUBS 0.024268f
C655 VTAIL.n571 VSUBS 0.013041f
C656 VTAIL.n572 VSUBS 0.030824f
C657 VTAIL.n573 VSUBS 0.013808f
C658 VTAIL.n574 VSUBS 0.024268f
C659 VTAIL.n575 VSUBS 0.013041f
C660 VTAIL.n576 VSUBS 0.023118f
C661 VTAIL.n577 VSUBS 0.019608f
C662 VTAIL.t7 VSUBS 0.066048f
C663 VTAIL.n578 VSUBS 0.178372f
C664 VTAIL.n579 VSUBS 1.66196f
C665 VTAIL.n580 VSUBS 0.013041f
C666 VTAIL.n581 VSUBS 0.013808f
C667 VTAIL.n582 VSUBS 0.030824f
C668 VTAIL.n583 VSUBS 0.030824f
C669 VTAIL.n584 VSUBS 0.013808f
C670 VTAIL.n585 VSUBS 0.013041f
C671 VTAIL.n586 VSUBS 0.024268f
C672 VTAIL.n587 VSUBS 0.024268f
C673 VTAIL.n588 VSUBS 0.013041f
C674 VTAIL.n589 VSUBS 0.013808f
C675 VTAIL.n590 VSUBS 0.030824f
C676 VTAIL.n591 VSUBS 0.030824f
C677 VTAIL.n592 VSUBS 0.013808f
C678 VTAIL.n593 VSUBS 0.013041f
C679 VTAIL.n594 VSUBS 0.024268f
C680 VTAIL.n595 VSUBS 0.024268f
C681 VTAIL.n596 VSUBS 0.013041f
C682 VTAIL.n597 VSUBS 0.013808f
C683 VTAIL.n598 VSUBS 0.030824f
C684 VTAIL.n599 VSUBS 0.030824f
C685 VTAIL.n600 VSUBS 0.013808f
C686 VTAIL.n601 VSUBS 0.013041f
C687 VTAIL.n602 VSUBS 0.024268f
C688 VTAIL.n603 VSUBS 0.024268f
C689 VTAIL.n604 VSUBS 0.013041f
C690 VTAIL.n605 VSUBS 0.013808f
C691 VTAIL.n606 VSUBS 0.030824f
C692 VTAIL.n607 VSUBS 0.030824f
C693 VTAIL.n608 VSUBS 0.013808f
C694 VTAIL.n609 VSUBS 0.013041f
C695 VTAIL.n610 VSUBS 0.024268f
C696 VTAIL.n611 VSUBS 0.024268f
C697 VTAIL.n612 VSUBS 0.013041f
C698 VTAIL.n613 VSUBS 0.013808f
C699 VTAIL.n614 VSUBS 0.030824f
C700 VTAIL.n615 VSUBS 0.030824f
C701 VTAIL.n616 VSUBS 0.013808f
C702 VTAIL.n617 VSUBS 0.013041f
C703 VTAIL.n618 VSUBS 0.024268f
C704 VTAIL.n619 VSUBS 0.024268f
C705 VTAIL.n620 VSUBS 0.013041f
C706 VTAIL.n621 VSUBS 0.013808f
C707 VTAIL.n622 VSUBS 0.030824f
C708 VTAIL.n623 VSUBS 0.030824f
C709 VTAIL.n624 VSUBS 0.030824f
C710 VTAIL.n625 VSUBS 0.013424f
C711 VTAIL.n626 VSUBS 0.013041f
C712 VTAIL.n627 VSUBS 0.024268f
C713 VTAIL.n628 VSUBS 0.024268f
C714 VTAIL.n629 VSUBS 0.013041f
C715 VTAIL.n630 VSUBS 0.013808f
C716 VTAIL.n631 VSUBS 0.030824f
C717 VTAIL.n632 VSUBS 0.067967f
C718 VTAIL.n633 VSUBS 0.013808f
C719 VTAIL.n634 VSUBS 0.013041f
C720 VTAIL.n635 VSUBS 0.054106f
C721 VTAIL.n636 VSUBS 0.033823f
C722 VTAIL.n637 VSUBS 1.57212f
C723 VTAIL.n638 VSUBS 0.024712f
C724 VTAIL.n639 VSUBS 0.024268f
C725 VTAIL.n640 VSUBS 0.013041f
C726 VTAIL.n641 VSUBS 0.030824f
C727 VTAIL.n642 VSUBS 0.013808f
C728 VTAIL.n643 VSUBS 0.024268f
C729 VTAIL.n644 VSUBS 0.013424f
C730 VTAIL.n645 VSUBS 0.030824f
C731 VTAIL.n646 VSUBS 0.013808f
C732 VTAIL.n647 VSUBS 0.024268f
C733 VTAIL.n648 VSUBS 0.013041f
C734 VTAIL.n649 VSUBS 0.030824f
C735 VTAIL.n650 VSUBS 0.013808f
C736 VTAIL.n651 VSUBS 0.024268f
C737 VTAIL.n652 VSUBS 0.013041f
C738 VTAIL.n653 VSUBS 0.030824f
C739 VTAIL.n654 VSUBS 0.013808f
C740 VTAIL.n655 VSUBS 0.024268f
C741 VTAIL.n656 VSUBS 0.013041f
C742 VTAIL.n657 VSUBS 0.030824f
C743 VTAIL.n658 VSUBS 0.013808f
C744 VTAIL.n659 VSUBS 0.024268f
C745 VTAIL.n660 VSUBS 0.013041f
C746 VTAIL.n661 VSUBS 0.030824f
C747 VTAIL.n662 VSUBS 0.013808f
C748 VTAIL.n663 VSUBS 0.024268f
C749 VTAIL.n664 VSUBS 0.013041f
C750 VTAIL.n665 VSUBS 0.023118f
C751 VTAIL.n666 VSUBS 0.019608f
C752 VTAIL.t5 VSUBS 0.066048f
C753 VTAIL.n667 VSUBS 0.178372f
C754 VTAIL.n668 VSUBS 1.66196f
C755 VTAIL.n669 VSUBS 0.013041f
C756 VTAIL.n670 VSUBS 0.013808f
C757 VTAIL.n671 VSUBS 0.030824f
C758 VTAIL.n672 VSUBS 0.030824f
C759 VTAIL.n673 VSUBS 0.013808f
C760 VTAIL.n674 VSUBS 0.013041f
C761 VTAIL.n675 VSUBS 0.024268f
C762 VTAIL.n676 VSUBS 0.024268f
C763 VTAIL.n677 VSUBS 0.013041f
C764 VTAIL.n678 VSUBS 0.013808f
C765 VTAIL.n679 VSUBS 0.030824f
C766 VTAIL.n680 VSUBS 0.030824f
C767 VTAIL.n681 VSUBS 0.013808f
C768 VTAIL.n682 VSUBS 0.013041f
C769 VTAIL.n683 VSUBS 0.024268f
C770 VTAIL.n684 VSUBS 0.024268f
C771 VTAIL.n685 VSUBS 0.013041f
C772 VTAIL.n686 VSUBS 0.013808f
C773 VTAIL.n687 VSUBS 0.030824f
C774 VTAIL.n688 VSUBS 0.030824f
C775 VTAIL.n689 VSUBS 0.013808f
C776 VTAIL.n690 VSUBS 0.013041f
C777 VTAIL.n691 VSUBS 0.024268f
C778 VTAIL.n692 VSUBS 0.024268f
C779 VTAIL.n693 VSUBS 0.013041f
C780 VTAIL.n694 VSUBS 0.013808f
C781 VTAIL.n695 VSUBS 0.030824f
C782 VTAIL.n696 VSUBS 0.030824f
C783 VTAIL.n697 VSUBS 0.013808f
C784 VTAIL.n698 VSUBS 0.013041f
C785 VTAIL.n699 VSUBS 0.024268f
C786 VTAIL.n700 VSUBS 0.024268f
C787 VTAIL.n701 VSUBS 0.013041f
C788 VTAIL.n702 VSUBS 0.013808f
C789 VTAIL.n703 VSUBS 0.030824f
C790 VTAIL.n704 VSUBS 0.030824f
C791 VTAIL.n705 VSUBS 0.013808f
C792 VTAIL.n706 VSUBS 0.013041f
C793 VTAIL.n707 VSUBS 0.024268f
C794 VTAIL.n708 VSUBS 0.024268f
C795 VTAIL.n709 VSUBS 0.013041f
C796 VTAIL.n710 VSUBS 0.013041f
C797 VTAIL.n711 VSUBS 0.013808f
C798 VTAIL.n712 VSUBS 0.030824f
C799 VTAIL.n713 VSUBS 0.030824f
C800 VTAIL.n714 VSUBS 0.030824f
C801 VTAIL.n715 VSUBS 0.013424f
C802 VTAIL.n716 VSUBS 0.013041f
C803 VTAIL.n717 VSUBS 0.024268f
C804 VTAIL.n718 VSUBS 0.024268f
C805 VTAIL.n719 VSUBS 0.013041f
C806 VTAIL.n720 VSUBS 0.013808f
C807 VTAIL.n721 VSUBS 0.030824f
C808 VTAIL.n722 VSUBS 0.067967f
C809 VTAIL.n723 VSUBS 0.013808f
C810 VTAIL.n724 VSUBS 0.013041f
C811 VTAIL.n725 VSUBS 0.054106f
C812 VTAIL.n726 VSUBS 0.033823f
C813 VTAIL.n727 VSUBS 1.56757f
C814 VDD1.t1 VSUBS 0.346451f
C815 VDD1.t2 VSUBS 0.346451f
C816 VDD1.n0 VSUBS 2.83475f
C817 VDD1.t4 VSUBS 0.346451f
C818 VDD1.t5 VSUBS 0.346451f
C819 VDD1.n1 VSUBS 2.83359f
C820 VDD1.t3 VSUBS 0.346451f
C821 VDD1.t7 VSUBS 0.346451f
C822 VDD1.n2 VSUBS 2.83359f
C823 VDD1.n3 VSUBS 3.34646f
C824 VDD1.t0 VSUBS 0.346451f
C825 VDD1.t6 VSUBS 0.346451f
C826 VDD1.n4 VSUBS 2.82972f
C827 VDD1.n5 VSUBS 3.20126f
C828 VP.n0 VSUBS 0.051824f
C829 VP.n1 VSUBS 0.01176f
C830 VP.n2 VSUBS 0.051824f
C831 VP.n3 VSUBS 0.051824f
C832 VP.t7 VSUBS 1.72073f
C833 VP.t1 VSUBS 1.72073f
C834 VP.n4 VSUBS 0.051824f
C835 VP.t2 VSUBS 1.72073f
C836 VP.n5 VSUBS 0.662723f
C837 VP.t0 VSUBS 1.74602f
C838 VP.n6 VSUBS 0.637242f
C839 VP.n7 VSUBS 0.219309f
C840 VP.n8 VSUBS 0.01176f
C841 VP.n9 VSUBS 0.656927f
C842 VP.n10 VSUBS 0.01176f
C843 VP.n11 VSUBS 0.655489f
C844 VP.n12 VSUBS 2.41228f
C845 VP.n13 VSUBS 2.4536f
C846 VP.t4 VSUBS 1.72073f
C847 VP.n14 VSUBS 0.655489f
C848 VP.n15 VSUBS 0.01176f
C849 VP.t3 VSUBS 1.72073f
C850 VP.n16 VSUBS 0.656927f
C851 VP.n17 VSUBS 0.051824f
C852 VP.n18 VSUBS 0.051824f
C853 VP.n19 VSUBS 0.051824f
C854 VP.t5 VSUBS 1.72073f
C855 VP.n20 VSUBS 0.656927f
C856 VP.n21 VSUBS 0.01176f
C857 VP.t6 VSUBS 1.72073f
C858 VP.n22 VSUBS 0.655489f
C859 VP.n23 VSUBS 0.040161f
C860 B.n0 VSUBS 0.006898f
C861 B.n1 VSUBS 0.006898f
C862 B.n2 VSUBS 0.010202f
C863 B.n3 VSUBS 0.007818f
C864 B.n4 VSUBS 0.007818f
C865 B.n5 VSUBS 0.007818f
C866 B.n6 VSUBS 0.007818f
C867 B.n7 VSUBS 0.007818f
C868 B.n8 VSUBS 0.007818f
C869 B.n9 VSUBS 0.007818f
C870 B.n10 VSUBS 0.007818f
C871 B.n11 VSUBS 0.007818f
C872 B.n12 VSUBS 0.007818f
C873 B.n13 VSUBS 0.019522f
C874 B.n14 VSUBS 0.007818f
C875 B.n15 VSUBS 0.007818f
C876 B.n16 VSUBS 0.007818f
C877 B.n17 VSUBS 0.007818f
C878 B.n18 VSUBS 0.007818f
C879 B.n19 VSUBS 0.007818f
C880 B.n20 VSUBS 0.007818f
C881 B.n21 VSUBS 0.007818f
C882 B.n22 VSUBS 0.007818f
C883 B.n23 VSUBS 0.007818f
C884 B.n24 VSUBS 0.007818f
C885 B.n25 VSUBS 0.007818f
C886 B.n26 VSUBS 0.007818f
C887 B.n27 VSUBS 0.007818f
C888 B.n28 VSUBS 0.007818f
C889 B.n29 VSUBS 0.007818f
C890 B.n30 VSUBS 0.007818f
C891 B.n31 VSUBS 0.007818f
C892 B.n32 VSUBS 0.007818f
C893 B.n33 VSUBS 0.007818f
C894 B.n34 VSUBS 0.007818f
C895 B.n35 VSUBS 0.007818f
C896 B.n36 VSUBS 0.007818f
C897 B.n37 VSUBS 0.007818f
C898 B.n38 VSUBS 0.007818f
C899 B.n39 VSUBS 0.007818f
C900 B.t7 VSUBS 0.33891f
C901 B.t8 VSUBS 0.352978f
C902 B.t6 VSUBS 0.531118f
C903 B.n40 VSUBS 0.44715f
C904 B.n41 VSUBS 0.331706f
C905 B.n42 VSUBS 0.018113f
C906 B.n43 VSUBS 0.007818f
C907 B.n44 VSUBS 0.007818f
C908 B.n45 VSUBS 0.007818f
C909 B.n46 VSUBS 0.007818f
C910 B.n47 VSUBS 0.007818f
C911 B.t4 VSUBS 0.338914f
C912 B.t5 VSUBS 0.352982f
C913 B.t3 VSUBS 0.531118f
C914 B.n48 VSUBS 0.447146f
C915 B.n49 VSUBS 0.331702f
C916 B.n50 VSUBS 0.007818f
C917 B.n51 VSUBS 0.007818f
C918 B.n52 VSUBS 0.007818f
C919 B.n53 VSUBS 0.007818f
C920 B.n54 VSUBS 0.007818f
C921 B.n55 VSUBS 0.007818f
C922 B.n56 VSUBS 0.007818f
C923 B.n57 VSUBS 0.007818f
C924 B.n58 VSUBS 0.007818f
C925 B.n59 VSUBS 0.007818f
C926 B.n60 VSUBS 0.007818f
C927 B.n61 VSUBS 0.007818f
C928 B.n62 VSUBS 0.007818f
C929 B.n63 VSUBS 0.007818f
C930 B.n64 VSUBS 0.007818f
C931 B.n65 VSUBS 0.007818f
C932 B.n66 VSUBS 0.007818f
C933 B.n67 VSUBS 0.007818f
C934 B.n68 VSUBS 0.007818f
C935 B.n69 VSUBS 0.007818f
C936 B.n70 VSUBS 0.007818f
C937 B.n71 VSUBS 0.007818f
C938 B.n72 VSUBS 0.007818f
C939 B.n73 VSUBS 0.007818f
C940 B.n74 VSUBS 0.007818f
C941 B.n75 VSUBS 0.007818f
C942 B.n76 VSUBS 0.019522f
C943 B.n77 VSUBS 0.007818f
C944 B.n78 VSUBS 0.007818f
C945 B.n79 VSUBS 0.007818f
C946 B.n80 VSUBS 0.007818f
C947 B.n81 VSUBS 0.007818f
C948 B.n82 VSUBS 0.007818f
C949 B.n83 VSUBS 0.007818f
C950 B.n84 VSUBS 0.007818f
C951 B.n85 VSUBS 0.007818f
C952 B.n86 VSUBS 0.007818f
C953 B.n87 VSUBS 0.007818f
C954 B.n88 VSUBS 0.007818f
C955 B.n89 VSUBS 0.007818f
C956 B.n90 VSUBS 0.007818f
C957 B.n91 VSUBS 0.007818f
C958 B.n92 VSUBS 0.007818f
C959 B.n93 VSUBS 0.007818f
C960 B.n94 VSUBS 0.007818f
C961 B.n95 VSUBS 0.007818f
C962 B.n96 VSUBS 0.007818f
C963 B.n97 VSUBS 0.007818f
C964 B.n98 VSUBS 0.007818f
C965 B.n99 VSUBS 0.007818f
C966 B.n100 VSUBS 0.019442f
C967 B.n101 VSUBS 0.007818f
C968 B.n102 VSUBS 0.007818f
C969 B.n103 VSUBS 0.007818f
C970 B.n104 VSUBS 0.007818f
C971 B.n105 VSUBS 0.007818f
C972 B.n106 VSUBS 0.007818f
C973 B.n107 VSUBS 0.007818f
C974 B.n108 VSUBS 0.007818f
C975 B.n109 VSUBS 0.007818f
C976 B.n110 VSUBS 0.007818f
C977 B.n111 VSUBS 0.007818f
C978 B.n112 VSUBS 0.007818f
C979 B.n113 VSUBS 0.007818f
C980 B.n114 VSUBS 0.007818f
C981 B.n115 VSUBS 0.007818f
C982 B.n116 VSUBS 0.007818f
C983 B.n117 VSUBS 0.007818f
C984 B.n118 VSUBS 0.007818f
C985 B.n119 VSUBS 0.007818f
C986 B.n120 VSUBS 0.007818f
C987 B.n121 VSUBS 0.007818f
C988 B.n122 VSUBS 0.007818f
C989 B.n123 VSUBS 0.007818f
C990 B.n124 VSUBS 0.007818f
C991 B.n125 VSUBS 0.007818f
C992 B.n126 VSUBS 0.007358f
C993 B.n127 VSUBS 0.007818f
C994 B.n128 VSUBS 0.007818f
C995 B.n129 VSUBS 0.007818f
C996 B.n130 VSUBS 0.007818f
C997 B.n131 VSUBS 0.007818f
C998 B.t2 VSUBS 0.33891f
C999 B.t1 VSUBS 0.352978f
C1000 B.t0 VSUBS 0.531118f
C1001 B.n132 VSUBS 0.44715f
C1002 B.n133 VSUBS 0.331706f
C1003 B.n134 VSUBS 0.007818f
C1004 B.n135 VSUBS 0.007818f
C1005 B.n136 VSUBS 0.007818f
C1006 B.n137 VSUBS 0.007818f
C1007 B.n138 VSUBS 0.007818f
C1008 B.n139 VSUBS 0.007818f
C1009 B.n140 VSUBS 0.007818f
C1010 B.n141 VSUBS 0.007818f
C1011 B.n142 VSUBS 0.007818f
C1012 B.n143 VSUBS 0.007818f
C1013 B.n144 VSUBS 0.007818f
C1014 B.n145 VSUBS 0.007818f
C1015 B.n146 VSUBS 0.007818f
C1016 B.n147 VSUBS 0.007818f
C1017 B.n148 VSUBS 0.007818f
C1018 B.n149 VSUBS 0.007818f
C1019 B.n150 VSUBS 0.007818f
C1020 B.n151 VSUBS 0.007818f
C1021 B.n152 VSUBS 0.007818f
C1022 B.n153 VSUBS 0.007818f
C1023 B.n154 VSUBS 0.007818f
C1024 B.n155 VSUBS 0.007818f
C1025 B.n156 VSUBS 0.007818f
C1026 B.n157 VSUBS 0.007818f
C1027 B.n158 VSUBS 0.007818f
C1028 B.n159 VSUBS 0.007818f
C1029 B.n160 VSUBS 0.019522f
C1030 B.n161 VSUBS 0.007818f
C1031 B.n162 VSUBS 0.007818f
C1032 B.n163 VSUBS 0.007818f
C1033 B.n164 VSUBS 0.007818f
C1034 B.n165 VSUBS 0.007818f
C1035 B.n166 VSUBS 0.007818f
C1036 B.n167 VSUBS 0.007818f
C1037 B.n168 VSUBS 0.007818f
C1038 B.n169 VSUBS 0.007818f
C1039 B.n170 VSUBS 0.007818f
C1040 B.n171 VSUBS 0.007818f
C1041 B.n172 VSUBS 0.007818f
C1042 B.n173 VSUBS 0.007818f
C1043 B.n174 VSUBS 0.007818f
C1044 B.n175 VSUBS 0.007818f
C1045 B.n176 VSUBS 0.007818f
C1046 B.n177 VSUBS 0.007818f
C1047 B.n178 VSUBS 0.007818f
C1048 B.n179 VSUBS 0.007818f
C1049 B.n180 VSUBS 0.007818f
C1050 B.n181 VSUBS 0.007818f
C1051 B.n182 VSUBS 0.007818f
C1052 B.n183 VSUBS 0.007818f
C1053 B.n184 VSUBS 0.007818f
C1054 B.n185 VSUBS 0.007818f
C1055 B.n186 VSUBS 0.007818f
C1056 B.n187 VSUBS 0.007818f
C1057 B.n188 VSUBS 0.007818f
C1058 B.n189 VSUBS 0.007818f
C1059 B.n190 VSUBS 0.007818f
C1060 B.n191 VSUBS 0.007818f
C1061 B.n192 VSUBS 0.007818f
C1062 B.n193 VSUBS 0.007818f
C1063 B.n194 VSUBS 0.007818f
C1064 B.n195 VSUBS 0.007818f
C1065 B.n196 VSUBS 0.007818f
C1066 B.n197 VSUBS 0.007818f
C1067 B.n198 VSUBS 0.007818f
C1068 B.n199 VSUBS 0.007818f
C1069 B.n200 VSUBS 0.007818f
C1070 B.n201 VSUBS 0.007818f
C1071 B.n202 VSUBS 0.007818f
C1072 B.n203 VSUBS 0.019522f
C1073 B.n204 VSUBS 0.020258f
C1074 B.n205 VSUBS 0.020258f
C1075 B.n206 VSUBS 0.007818f
C1076 B.n207 VSUBS 0.007818f
C1077 B.n208 VSUBS 0.007818f
C1078 B.n209 VSUBS 0.007818f
C1079 B.n210 VSUBS 0.007818f
C1080 B.n211 VSUBS 0.007818f
C1081 B.n212 VSUBS 0.007818f
C1082 B.n213 VSUBS 0.007818f
C1083 B.n214 VSUBS 0.007818f
C1084 B.n215 VSUBS 0.007818f
C1085 B.n216 VSUBS 0.007818f
C1086 B.n217 VSUBS 0.007818f
C1087 B.n218 VSUBS 0.007818f
C1088 B.n219 VSUBS 0.007818f
C1089 B.n220 VSUBS 0.007818f
C1090 B.n221 VSUBS 0.007818f
C1091 B.n222 VSUBS 0.007818f
C1092 B.n223 VSUBS 0.007818f
C1093 B.n224 VSUBS 0.007818f
C1094 B.n225 VSUBS 0.007818f
C1095 B.n226 VSUBS 0.007818f
C1096 B.n227 VSUBS 0.007818f
C1097 B.n228 VSUBS 0.007818f
C1098 B.n229 VSUBS 0.007818f
C1099 B.n230 VSUBS 0.007818f
C1100 B.n231 VSUBS 0.007818f
C1101 B.n232 VSUBS 0.007818f
C1102 B.n233 VSUBS 0.007818f
C1103 B.n234 VSUBS 0.007818f
C1104 B.n235 VSUBS 0.007818f
C1105 B.n236 VSUBS 0.007818f
C1106 B.n237 VSUBS 0.007818f
C1107 B.n238 VSUBS 0.007818f
C1108 B.n239 VSUBS 0.007818f
C1109 B.n240 VSUBS 0.007818f
C1110 B.n241 VSUBS 0.007818f
C1111 B.n242 VSUBS 0.007818f
C1112 B.n243 VSUBS 0.007818f
C1113 B.n244 VSUBS 0.007818f
C1114 B.n245 VSUBS 0.007818f
C1115 B.n246 VSUBS 0.007818f
C1116 B.n247 VSUBS 0.007818f
C1117 B.n248 VSUBS 0.007818f
C1118 B.n249 VSUBS 0.007818f
C1119 B.n250 VSUBS 0.007818f
C1120 B.n251 VSUBS 0.007818f
C1121 B.n252 VSUBS 0.007818f
C1122 B.n253 VSUBS 0.007818f
C1123 B.n254 VSUBS 0.007818f
C1124 B.n255 VSUBS 0.007818f
C1125 B.n256 VSUBS 0.007818f
C1126 B.n257 VSUBS 0.007818f
C1127 B.n258 VSUBS 0.007818f
C1128 B.n259 VSUBS 0.007818f
C1129 B.n260 VSUBS 0.007818f
C1130 B.n261 VSUBS 0.007818f
C1131 B.n262 VSUBS 0.007818f
C1132 B.n263 VSUBS 0.007818f
C1133 B.n264 VSUBS 0.007818f
C1134 B.n265 VSUBS 0.007818f
C1135 B.n266 VSUBS 0.007818f
C1136 B.n267 VSUBS 0.007818f
C1137 B.n268 VSUBS 0.007818f
C1138 B.n269 VSUBS 0.007818f
C1139 B.n270 VSUBS 0.007818f
C1140 B.n271 VSUBS 0.007818f
C1141 B.n272 VSUBS 0.007818f
C1142 B.n273 VSUBS 0.007818f
C1143 B.n274 VSUBS 0.007818f
C1144 B.n275 VSUBS 0.007818f
C1145 B.n276 VSUBS 0.007818f
C1146 B.n277 VSUBS 0.007818f
C1147 B.n278 VSUBS 0.007818f
C1148 B.n279 VSUBS 0.007818f
C1149 B.n280 VSUBS 0.007818f
C1150 B.n281 VSUBS 0.007818f
C1151 B.n282 VSUBS 0.007818f
C1152 B.n283 VSUBS 0.007358f
C1153 B.n284 VSUBS 0.018113f
C1154 B.n285 VSUBS 0.004369f
C1155 B.n286 VSUBS 0.007818f
C1156 B.n287 VSUBS 0.007818f
C1157 B.n288 VSUBS 0.007818f
C1158 B.n289 VSUBS 0.007818f
C1159 B.n290 VSUBS 0.007818f
C1160 B.n291 VSUBS 0.007818f
C1161 B.n292 VSUBS 0.007818f
C1162 B.n293 VSUBS 0.007818f
C1163 B.n294 VSUBS 0.007818f
C1164 B.n295 VSUBS 0.007818f
C1165 B.n296 VSUBS 0.007818f
C1166 B.n297 VSUBS 0.007818f
C1167 B.t11 VSUBS 0.338914f
C1168 B.t10 VSUBS 0.352982f
C1169 B.t9 VSUBS 0.531118f
C1170 B.n298 VSUBS 0.447146f
C1171 B.n299 VSUBS 0.331702f
C1172 B.n300 VSUBS 0.018113f
C1173 B.n301 VSUBS 0.004369f
C1174 B.n302 VSUBS 0.007818f
C1175 B.n303 VSUBS 0.007818f
C1176 B.n304 VSUBS 0.007818f
C1177 B.n305 VSUBS 0.007818f
C1178 B.n306 VSUBS 0.007818f
C1179 B.n307 VSUBS 0.007818f
C1180 B.n308 VSUBS 0.007818f
C1181 B.n309 VSUBS 0.007818f
C1182 B.n310 VSUBS 0.007818f
C1183 B.n311 VSUBS 0.007818f
C1184 B.n312 VSUBS 0.007818f
C1185 B.n313 VSUBS 0.007818f
C1186 B.n314 VSUBS 0.007818f
C1187 B.n315 VSUBS 0.007818f
C1188 B.n316 VSUBS 0.007818f
C1189 B.n317 VSUBS 0.007818f
C1190 B.n318 VSUBS 0.007818f
C1191 B.n319 VSUBS 0.007818f
C1192 B.n320 VSUBS 0.007818f
C1193 B.n321 VSUBS 0.007818f
C1194 B.n322 VSUBS 0.007818f
C1195 B.n323 VSUBS 0.007818f
C1196 B.n324 VSUBS 0.007818f
C1197 B.n325 VSUBS 0.007818f
C1198 B.n326 VSUBS 0.007818f
C1199 B.n327 VSUBS 0.007818f
C1200 B.n328 VSUBS 0.007818f
C1201 B.n329 VSUBS 0.007818f
C1202 B.n330 VSUBS 0.007818f
C1203 B.n331 VSUBS 0.007818f
C1204 B.n332 VSUBS 0.007818f
C1205 B.n333 VSUBS 0.007818f
C1206 B.n334 VSUBS 0.007818f
C1207 B.n335 VSUBS 0.007818f
C1208 B.n336 VSUBS 0.007818f
C1209 B.n337 VSUBS 0.007818f
C1210 B.n338 VSUBS 0.007818f
C1211 B.n339 VSUBS 0.007818f
C1212 B.n340 VSUBS 0.007818f
C1213 B.n341 VSUBS 0.007818f
C1214 B.n342 VSUBS 0.007818f
C1215 B.n343 VSUBS 0.007818f
C1216 B.n344 VSUBS 0.007818f
C1217 B.n345 VSUBS 0.007818f
C1218 B.n346 VSUBS 0.007818f
C1219 B.n347 VSUBS 0.007818f
C1220 B.n348 VSUBS 0.007818f
C1221 B.n349 VSUBS 0.007818f
C1222 B.n350 VSUBS 0.007818f
C1223 B.n351 VSUBS 0.007818f
C1224 B.n352 VSUBS 0.007818f
C1225 B.n353 VSUBS 0.007818f
C1226 B.n354 VSUBS 0.007818f
C1227 B.n355 VSUBS 0.007818f
C1228 B.n356 VSUBS 0.007818f
C1229 B.n357 VSUBS 0.007818f
C1230 B.n358 VSUBS 0.007818f
C1231 B.n359 VSUBS 0.007818f
C1232 B.n360 VSUBS 0.007818f
C1233 B.n361 VSUBS 0.007818f
C1234 B.n362 VSUBS 0.007818f
C1235 B.n363 VSUBS 0.007818f
C1236 B.n364 VSUBS 0.007818f
C1237 B.n365 VSUBS 0.007818f
C1238 B.n366 VSUBS 0.007818f
C1239 B.n367 VSUBS 0.007818f
C1240 B.n368 VSUBS 0.007818f
C1241 B.n369 VSUBS 0.007818f
C1242 B.n370 VSUBS 0.007818f
C1243 B.n371 VSUBS 0.007818f
C1244 B.n372 VSUBS 0.007818f
C1245 B.n373 VSUBS 0.007818f
C1246 B.n374 VSUBS 0.007818f
C1247 B.n375 VSUBS 0.007818f
C1248 B.n376 VSUBS 0.007818f
C1249 B.n377 VSUBS 0.007818f
C1250 B.n378 VSUBS 0.007818f
C1251 B.n379 VSUBS 0.007818f
C1252 B.n380 VSUBS 0.007818f
C1253 B.n381 VSUBS 0.020258f
C1254 B.n382 VSUBS 0.019522f
C1255 B.n383 VSUBS 0.020337f
C1256 B.n384 VSUBS 0.007818f
C1257 B.n385 VSUBS 0.007818f
C1258 B.n386 VSUBS 0.007818f
C1259 B.n387 VSUBS 0.007818f
C1260 B.n388 VSUBS 0.007818f
C1261 B.n389 VSUBS 0.007818f
C1262 B.n390 VSUBS 0.007818f
C1263 B.n391 VSUBS 0.007818f
C1264 B.n392 VSUBS 0.007818f
C1265 B.n393 VSUBS 0.007818f
C1266 B.n394 VSUBS 0.007818f
C1267 B.n395 VSUBS 0.007818f
C1268 B.n396 VSUBS 0.007818f
C1269 B.n397 VSUBS 0.007818f
C1270 B.n398 VSUBS 0.007818f
C1271 B.n399 VSUBS 0.007818f
C1272 B.n400 VSUBS 0.007818f
C1273 B.n401 VSUBS 0.007818f
C1274 B.n402 VSUBS 0.007818f
C1275 B.n403 VSUBS 0.007818f
C1276 B.n404 VSUBS 0.007818f
C1277 B.n405 VSUBS 0.007818f
C1278 B.n406 VSUBS 0.007818f
C1279 B.n407 VSUBS 0.007818f
C1280 B.n408 VSUBS 0.007818f
C1281 B.n409 VSUBS 0.007818f
C1282 B.n410 VSUBS 0.007818f
C1283 B.n411 VSUBS 0.007818f
C1284 B.n412 VSUBS 0.007818f
C1285 B.n413 VSUBS 0.007818f
C1286 B.n414 VSUBS 0.007818f
C1287 B.n415 VSUBS 0.007818f
C1288 B.n416 VSUBS 0.007818f
C1289 B.n417 VSUBS 0.007818f
C1290 B.n418 VSUBS 0.007818f
C1291 B.n419 VSUBS 0.007818f
C1292 B.n420 VSUBS 0.007818f
C1293 B.n421 VSUBS 0.007818f
C1294 B.n422 VSUBS 0.007818f
C1295 B.n423 VSUBS 0.007818f
C1296 B.n424 VSUBS 0.007818f
C1297 B.n425 VSUBS 0.007818f
C1298 B.n426 VSUBS 0.007818f
C1299 B.n427 VSUBS 0.007818f
C1300 B.n428 VSUBS 0.007818f
C1301 B.n429 VSUBS 0.007818f
C1302 B.n430 VSUBS 0.007818f
C1303 B.n431 VSUBS 0.007818f
C1304 B.n432 VSUBS 0.007818f
C1305 B.n433 VSUBS 0.007818f
C1306 B.n434 VSUBS 0.007818f
C1307 B.n435 VSUBS 0.007818f
C1308 B.n436 VSUBS 0.007818f
C1309 B.n437 VSUBS 0.007818f
C1310 B.n438 VSUBS 0.007818f
C1311 B.n439 VSUBS 0.007818f
C1312 B.n440 VSUBS 0.007818f
C1313 B.n441 VSUBS 0.007818f
C1314 B.n442 VSUBS 0.007818f
C1315 B.n443 VSUBS 0.007818f
C1316 B.n444 VSUBS 0.007818f
C1317 B.n445 VSUBS 0.007818f
C1318 B.n446 VSUBS 0.007818f
C1319 B.n447 VSUBS 0.007818f
C1320 B.n448 VSUBS 0.007818f
C1321 B.n449 VSUBS 0.007818f
C1322 B.n450 VSUBS 0.007818f
C1323 B.n451 VSUBS 0.007818f
C1324 B.n452 VSUBS 0.007818f
C1325 B.n453 VSUBS 0.019522f
C1326 B.n454 VSUBS 0.020258f
C1327 B.n455 VSUBS 0.020258f
C1328 B.n456 VSUBS 0.007818f
C1329 B.n457 VSUBS 0.007818f
C1330 B.n458 VSUBS 0.007818f
C1331 B.n459 VSUBS 0.007818f
C1332 B.n460 VSUBS 0.007818f
C1333 B.n461 VSUBS 0.007818f
C1334 B.n462 VSUBS 0.007818f
C1335 B.n463 VSUBS 0.007818f
C1336 B.n464 VSUBS 0.007818f
C1337 B.n465 VSUBS 0.007818f
C1338 B.n466 VSUBS 0.007818f
C1339 B.n467 VSUBS 0.007818f
C1340 B.n468 VSUBS 0.007818f
C1341 B.n469 VSUBS 0.007818f
C1342 B.n470 VSUBS 0.007818f
C1343 B.n471 VSUBS 0.007818f
C1344 B.n472 VSUBS 0.007818f
C1345 B.n473 VSUBS 0.007818f
C1346 B.n474 VSUBS 0.007818f
C1347 B.n475 VSUBS 0.007818f
C1348 B.n476 VSUBS 0.007818f
C1349 B.n477 VSUBS 0.007818f
C1350 B.n478 VSUBS 0.007818f
C1351 B.n479 VSUBS 0.007818f
C1352 B.n480 VSUBS 0.007818f
C1353 B.n481 VSUBS 0.007818f
C1354 B.n482 VSUBS 0.007818f
C1355 B.n483 VSUBS 0.007818f
C1356 B.n484 VSUBS 0.007818f
C1357 B.n485 VSUBS 0.007818f
C1358 B.n486 VSUBS 0.007818f
C1359 B.n487 VSUBS 0.007818f
C1360 B.n488 VSUBS 0.007818f
C1361 B.n489 VSUBS 0.007818f
C1362 B.n490 VSUBS 0.007818f
C1363 B.n491 VSUBS 0.007818f
C1364 B.n492 VSUBS 0.007818f
C1365 B.n493 VSUBS 0.007818f
C1366 B.n494 VSUBS 0.007818f
C1367 B.n495 VSUBS 0.007818f
C1368 B.n496 VSUBS 0.007818f
C1369 B.n497 VSUBS 0.007818f
C1370 B.n498 VSUBS 0.007818f
C1371 B.n499 VSUBS 0.007818f
C1372 B.n500 VSUBS 0.007818f
C1373 B.n501 VSUBS 0.007818f
C1374 B.n502 VSUBS 0.007818f
C1375 B.n503 VSUBS 0.007818f
C1376 B.n504 VSUBS 0.007818f
C1377 B.n505 VSUBS 0.007818f
C1378 B.n506 VSUBS 0.007818f
C1379 B.n507 VSUBS 0.007818f
C1380 B.n508 VSUBS 0.007818f
C1381 B.n509 VSUBS 0.007818f
C1382 B.n510 VSUBS 0.007818f
C1383 B.n511 VSUBS 0.007818f
C1384 B.n512 VSUBS 0.007818f
C1385 B.n513 VSUBS 0.007818f
C1386 B.n514 VSUBS 0.007818f
C1387 B.n515 VSUBS 0.007818f
C1388 B.n516 VSUBS 0.007818f
C1389 B.n517 VSUBS 0.007818f
C1390 B.n518 VSUBS 0.007818f
C1391 B.n519 VSUBS 0.007818f
C1392 B.n520 VSUBS 0.007818f
C1393 B.n521 VSUBS 0.007818f
C1394 B.n522 VSUBS 0.007818f
C1395 B.n523 VSUBS 0.007818f
C1396 B.n524 VSUBS 0.007818f
C1397 B.n525 VSUBS 0.007818f
C1398 B.n526 VSUBS 0.007818f
C1399 B.n527 VSUBS 0.007818f
C1400 B.n528 VSUBS 0.007818f
C1401 B.n529 VSUBS 0.007818f
C1402 B.n530 VSUBS 0.007818f
C1403 B.n531 VSUBS 0.007818f
C1404 B.n532 VSUBS 0.007818f
C1405 B.n533 VSUBS 0.007358f
C1406 B.n534 VSUBS 0.018113f
C1407 B.n535 VSUBS 0.004369f
C1408 B.n536 VSUBS 0.007818f
C1409 B.n537 VSUBS 0.007818f
C1410 B.n538 VSUBS 0.007818f
C1411 B.n539 VSUBS 0.007818f
C1412 B.n540 VSUBS 0.007818f
C1413 B.n541 VSUBS 0.007818f
C1414 B.n542 VSUBS 0.007818f
C1415 B.n543 VSUBS 0.007818f
C1416 B.n544 VSUBS 0.007818f
C1417 B.n545 VSUBS 0.007818f
C1418 B.n546 VSUBS 0.007818f
C1419 B.n547 VSUBS 0.007818f
C1420 B.n548 VSUBS 0.004369f
C1421 B.n549 VSUBS 0.007818f
C1422 B.n550 VSUBS 0.007818f
C1423 B.n551 VSUBS 0.007358f
C1424 B.n552 VSUBS 0.007818f
C1425 B.n553 VSUBS 0.007818f
C1426 B.n554 VSUBS 0.007818f
C1427 B.n555 VSUBS 0.007818f
C1428 B.n556 VSUBS 0.007818f
C1429 B.n557 VSUBS 0.007818f
C1430 B.n558 VSUBS 0.007818f
C1431 B.n559 VSUBS 0.007818f
C1432 B.n560 VSUBS 0.007818f
C1433 B.n561 VSUBS 0.007818f
C1434 B.n562 VSUBS 0.007818f
C1435 B.n563 VSUBS 0.007818f
C1436 B.n564 VSUBS 0.007818f
C1437 B.n565 VSUBS 0.007818f
C1438 B.n566 VSUBS 0.007818f
C1439 B.n567 VSUBS 0.007818f
C1440 B.n568 VSUBS 0.007818f
C1441 B.n569 VSUBS 0.007818f
C1442 B.n570 VSUBS 0.007818f
C1443 B.n571 VSUBS 0.007818f
C1444 B.n572 VSUBS 0.007818f
C1445 B.n573 VSUBS 0.007818f
C1446 B.n574 VSUBS 0.007818f
C1447 B.n575 VSUBS 0.007818f
C1448 B.n576 VSUBS 0.007818f
C1449 B.n577 VSUBS 0.007818f
C1450 B.n578 VSUBS 0.007818f
C1451 B.n579 VSUBS 0.007818f
C1452 B.n580 VSUBS 0.007818f
C1453 B.n581 VSUBS 0.007818f
C1454 B.n582 VSUBS 0.007818f
C1455 B.n583 VSUBS 0.007818f
C1456 B.n584 VSUBS 0.007818f
C1457 B.n585 VSUBS 0.007818f
C1458 B.n586 VSUBS 0.007818f
C1459 B.n587 VSUBS 0.007818f
C1460 B.n588 VSUBS 0.007818f
C1461 B.n589 VSUBS 0.007818f
C1462 B.n590 VSUBS 0.007818f
C1463 B.n591 VSUBS 0.007818f
C1464 B.n592 VSUBS 0.007818f
C1465 B.n593 VSUBS 0.007818f
C1466 B.n594 VSUBS 0.007818f
C1467 B.n595 VSUBS 0.007818f
C1468 B.n596 VSUBS 0.007818f
C1469 B.n597 VSUBS 0.007818f
C1470 B.n598 VSUBS 0.007818f
C1471 B.n599 VSUBS 0.007818f
C1472 B.n600 VSUBS 0.007818f
C1473 B.n601 VSUBS 0.007818f
C1474 B.n602 VSUBS 0.007818f
C1475 B.n603 VSUBS 0.007818f
C1476 B.n604 VSUBS 0.007818f
C1477 B.n605 VSUBS 0.007818f
C1478 B.n606 VSUBS 0.007818f
C1479 B.n607 VSUBS 0.007818f
C1480 B.n608 VSUBS 0.007818f
C1481 B.n609 VSUBS 0.007818f
C1482 B.n610 VSUBS 0.007818f
C1483 B.n611 VSUBS 0.007818f
C1484 B.n612 VSUBS 0.007818f
C1485 B.n613 VSUBS 0.007818f
C1486 B.n614 VSUBS 0.007818f
C1487 B.n615 VSUBS 0.007818f
C1488 B.n616 VSUBS 0.007818f
C1489 B.n617 VSUBS 0.007818f
C1490 B.n618 VSUBS 0.007818f
C1491 B.n619 VSUBS 0.007818f
C1492 B.n620 VSUBS 0.007818f
C1493 B.n621 VSUBS 0.007818f
C1494 B.n622 VSUBS 0.007818f
C1495 B.n623 VSUBS 0.007818f
C1496 B.n624 VSUBS 0.007818f
C1497 B.n625 VSUBS 0.007818f
C1498 B.n626 VSUBS 0.007818f
C1499 B.n627 VSUBS 0.007818f
C1500 B.n628 VSUBS 0.020258f
C1501 B.n629 VSUBS 0.020258f
C1502 B.n630 VSUBS 0.019522f
C1503 B.n631 VSUBS 0.007818f
C1504 B.n632 VSUBS 0.007818f
C1505 B.n633 VSUBS 0.007818f
C1506 B.n634 VSUBS 0.007818f
C1507 B.n635 VSUBS 0.007818f
C1508 B.n636 VSUBS 0.007818f
C1509 B.n637 VSUBS 0.007818f
C1510 B.n638 VSUBS 0.007818f
C1511 B.n639 VSUBS 0.007818f
C1512 B.n640 VSUBS 0.007818f
C1513 B.n641 VSUBS 0.007818f
C1514 B.n642 VSUBS 0.007818f
C1515 B.n643 VSUBS 0.007818f
C1516 B.n644 VSUBS 0.007818f
C1517 B.n645 VSUBS 0.007818f
C1518 B.n646 VSUBS 0.007818f
C1519 B.n647 VSUBS 0.007818f
C1520 B.n648 VSUBS 0.007818f
C1521 B.n649 VSUBS 0.007818f
C1522 B.n650 VSUBS 0.007818f
C1523 B.n651 VSUBS 0.007818f
C1524 B.n652 VSUBS 0.007818f
C1525 B.n653 VSUBS 0.007818f
C1526 B.n654 VSUBS 0.007818f
C1527 B.n655 VSUBS 0.007818f
C1528 B.n656 VSUBS 0.007818f
C1529 B.n657 VSUBS 0.007818f
C1530 B.n658 VSUBS 0.007818f
C1531 B.n659 VSUBS 0.007818f
C1532 B.n660 VSUBS 0.007818f
C1533 B.n661 VSUBS 0.007818f
C1534 B.n662 VSUBS 0.007818f
C1535 B.n663 VSUBS 0.010202f
C1536 B.n664 VSUBS 0.010868f
C1537 B.n665 VSUBS 0.021612f
.ends

