* NGSPICE file created from diff_pair_sample_0192.ext - technology: sky130A

.subckt diff_pair_sample_0192 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t7 VN.t0 VTAIL.t10 B.t4 sky130_fd_pr__nfet_01v8 ad=2.7489 pd=16.99 as=2.7489 ps=16.99 w=16.66 l=3.22
X1 B.t20 B.t18 B.t19 B.t12 sky130_fd_pr__nfet_01v8 ad=6.4974 pd=34.1 as=0 ps=0 w=16.66 l=3.22
X2 VTAIL.t14 VN.t1 VDD2.t6 B.t5 sky130_fd_pr__nfet_01v8 ad=6.4974 pd=34.1 as=2.7489 ps=16.99 w=16.66 l=3.22
X3 VTAIL.t13 VN.t2 VDD2.t5 B.t21 sky130_fd_pr__nfet_01v8 ad=2.7489 pd=16.99 as=2.7489 ps=16.99 w=16.66 l=3.22
X4 VDD1.t7 VP.t0 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=2.7489 pd=16.99 as=6.4974 ps=34.1 w=16.66 l=3.22
X5 VDD2.t4 VN.t3 VTAIL.t7 B.t2 sky130_fd_pr__nfet_01v8 ad=2.7489 pd=16.99 as=2.7489 ps=16.99 w=16.66 l=3.22
X6 VTAIL.t5 VP.t1 VDD1.t6 B.t5 sky130_fd_pr__nfet_01v8 ad=6.4974 pd=34.1 as=2.7489 ps=16.99 w=16.66 l=3.22
X7 VTAIL.t12 VN.t4 VDD2.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=6.4974 pd=34.1 as=2.7489 ps=16.99 w=16.66 l=3.22
X8 B.t17 B.t15 B.t16 B.t8 sky130_fd_pr__nfet_01v8 ad=6.4974 pd=34.1 as=0 ps=0 w=16.66 l=3.22
X9 VTAIL.t0 VP.t2 VDD1.t5 B.t0 sky130_fd_pr__nfet_01v8 ad=2.7489 pd=16.99 as=2.7489 ps=16.99 w=16.66 l=3.22
X10 VDD2.t2 VN.t5 VTAIL.t9 B.t6 sky130_fd_pr__nfet_01v8 ad=2.7489 pd=16.99 as=6.4974 ps=34.1 w=16.66 l=3.22
X11 VTAIL.t11 VN.t6 VDD2.t1 B.t0 sky130_fd_pr__nfet_01v8 ad=2.7489 pd=16.99 as=2.7489 ps=16.99 w=16.66 l=3.22
X12 VDD1.t4 VP.t3 VTAIL.t6 B.t6 sky130_fd_pr__nfet_01v8 ad=2.7489 pd=16.99 as=6.4974 ps=34.1 w=16.66 l=3.22
X13 VDD1.t3 VP.t4 VTAIL.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=2.7489 pd=16.99 as=2.7489 ps=16.99 w=16.66 l=3.22
X14 VTAIL.t3 VP.t5 VDD1.t2 B.t3 sky130_fd_pr__nfet_01v8 ad=6.4974 pd=34.1 as=2.7489 ps=16.99 w=16.66 l=3.22
X15 B.t14 B.t11 B.t13 B.t12 sky130_fd_pr__nfet_01v8 ad=6.4974 pd=34.1 as=0 ps=0 w=16.66 l=3.22
X16 VTAIL.t15 VP.t6 VDD1.t1 B.t21 sky130_fd_pr__nfet_01v8 ad=2.7489 pd=16.99 as=2.7489 ps=16.99 w=16.66 l=3.22
X17 VDD2.t0 VN.t7 VTAIL.t8 B.t1 sky130_fd_pr__nfet_01v8 ad=2.7489 pd=16.99 as=6.4974 ps=34.1 w=16.66 l=3.22
X18 VDD1.t0 VP.t7 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=2.7489 pd=16.99 as=2.7489 ps=16.99 w=16.66 l=3.22
X19 B.t10 B.t7 B.t9 B.t8 sky130_fd_pr__nfet_01v8 ad=6.4974 pd=34.1 as=0 ps=0 w=16.66 l=3.22
R0 VN.n64 VN.n63 161.3
R1 VN.n62 VN.n34 161.3
R2 VN.n61 VN.n60 161.3
R3 VN.n59 VN.n35 161.3
R4 VN.n58 VN.n57 161.3
R5 VN.n56 VN.n36 161.3
R6 VN.n55 VN.n54 161.3
R7 VN.n53 VN.n52 161.3
R8 VN.n51 VN.n38 161.3
R9 VN.n50 VN.n49 161.3
R10 VN.n48 VN.n39 161.3
R11 VN.n47 VN.n46 161.3
R12 VN.n45 VN.n40 161.3
R13 VN.n44 VN.n43 161.3
R14 VN.n31 VN.n30 161.3
R15 VN.n29 VN.n1 161.3
R16 VN.n28 VN.n27 161.3
R17 VN.n26 VN.n2 161.3
R18 VN.n25 VN.n24 161.3
R19 VN.n23 VN.n3 161.3
R20 VN.n22 VN.n21 161.3
R21 VN.n20 VN.n19 161.3
R22 VN.n18 VN.n5 161.3
R23 VN.n17 VN.n16 161.3
R24 VN.n15 VN.n6 161.3
R25 VN.n14 VN.n13 161.3
R26 VN.n12 VN.n7 161.3
R27 VN.n11 VN.n10 161.3
R28 VN.n42 VN.t5 157.864
R29 VN.n9 VN.t1 157.864
R30 VN.n8 VN.t3 124.692
R31 VN.n4 VN.t6 124.692
R32 VN.n0 VN.t7 124.692
R33 VN.n41 VN.t2 124.692
R34 VN.n37 VN.t0 124.692
R35 VN.n33 VN.t4 124.692
R36 VN.n32 VN.n0 74.2609
R37 VN.n65 VN.n33 74.2609
R38 VN.n9 VN.n8 60.9336
R39 VN.n42 VN.n41 60.9336
R40 VN VN.n65 57.6042
R41 VN.n28 VN.n2 45.4209
R42 VN.n61 VN.n35 45.4209
R43 VN.n13 VN.n6 40.577
R44 VN.n17 VN.n6 40.577
R45 VN.n46 VN.n39 40.577
R46 VN.n50 VN.n39 40.577
R47 VN.n24 VN.n2 35.7332
R48 VN.n57 VN.n35 35.7332
R49 VN.n12 VN.n11 24.5923
R50 VN.n13 VN.n12 24.5923
R51 VN.n18 VN.n17 24.5923
R52 VN.n19 VN.n18 24.5923
R53 VN.n23 VN.n22 24.5923
R54 VN.n24 VN.n23 24.5923
R55 VN.n29 VN.n28 24.5923
R56 VN.n30 VN.n29 24.5923
R57 VN.n46 VN.n45 24.5923
R58 VN.n45 VN.n44 24.5923
R59 VN.n57 VN.n56 24.5923
R60 VN.n56 VN.n55 24.5923
R61 VN.n52 VN.n51 24.5923
R62 VN.n51 VN.n50 24.5923
R63 VN.n63 VN.n62 24.5923
R64 VN.n62 VN.n61 24.5923
R65 VN.n30 VN.n0 15.9852
R66 VN.n63 VN.n33 15.9852
R67 VN.n11 VN.n8 13.526
R68 VN.n19 VN.n4 13.526
R69 VN.n44 VN.n41 13.526
R70 VN.n52 VN.n37 13.526
R71 VN.n22 VN.n4 11.0668
R72 VN.n55 VN.n37 11.0668
R73 VN.n43 VN.n42 4.08484
R74 VN.n10 VN.n9 4.08484
R75 VN.n65 VN.n64 0.354861
R76 VN.n32 VN.n31 0.354861
R77 VN VN.n32 0.267071
R78 VN.n64 VN.n34 0.189894
R79 VN.n60 VN.n34 0.189894
R80 VN.n60 VN.n59 0.189894
R81 VN.n59 VN.n58 0.189894
R82 VN.n58 VN.n36 0.189894
R83 VN.n54 VN.n36 0.189894
R84 VN.n54 VN.n53 0.189894
R85 VN.n53 VN.n38 0.189894
R86 VN.n49 VN.n38 0.189894
R87 VN.n49 VN.n48 0.189894
R88 VN.n48 VN.n47 0.189894
R89 VN.n47 VN.n40 0.189894
R90 VN.n43 VN.n40 0.189894
R91 VN.n10 VN.n7 0.189894
R92 VN.n14 VN.n7 0.189894
R93 VN.n15 VN.n14 0.189894
R94 VN.n16 VN.n15 0.189894
R95 VN.n16 VN.n5 0.189894
R96 VN.n20 VN.n5 0.189894
R97 VN.n21 VN.n20 0.189894
R98 VN.n21 VN.n3 0.189894
R99 VN.n25 VN.n3 0.189894
R100 VN.n26 VN.n25 0.189894
R101 VN.n27 VN.n26 0.189894
R102 VN.n27 VN.n1 0.189894
R103 VN.n31 VN.n1 0.189894
R104 VTAIL.n742 VTAIL.n741 289.615
R105 VTAIL.n92 VTAIL.n91 289.615
R106 VTAIL.n184 VTAIL.n183 289.615
R107 VTAIL.n278 VTAIL.n277 289.615
R108 VTAIL.n650 VTAIL.n649 289.615
R109 VTAIL.n556 VTAIL.n555 289.615
R110 VTAIL.n464 VTAIL.n463 289.615
R111 VTAIL.n370 VTAIL.n369 289.615
R112 VTAIL.n683 VTAIL.n682 185
R113 VTAIL.n685 VTAIL.n684 185
R114 VTAIL.n678 VTAIL.n677 185
R115 VTAIL.n691 VTAIL.n690 185
R116 VTAIL.n693 VTAIL.n692 185
R117 VTAIL.n674 VTAIL.n673 185
R118 VTAIL.n700 VTAIL.n699 185
R119 VTAIL.n701 VTAIL.n672 185
R120 VTAIL.n703 VTAIL.n702 185
R121 VTAIL.n670 VTAIL.n669 185
R122 VTAIL.n709 VTAIL.n708 185
R123 VTAIL.n711 VTAIL.n710 185
R124 VTAIL.n666 VTAIL.n665 185
R125 VTAIL.n717 VTAIL.n716 185
R126 VTAIL.n719 VTAIL.n718 185
R127 VTAIL.n662 VTAIL.n661 185
R128 VTAIL.n725 VTAIL.n724 185
R129 VTAIL.n727 VTAIL.n726 185
R130 VTAIL.n658 VTAIL.n657 185
R131 VTAIL.n733 VTAIL.n732 185
R132 VTAIL.n735 VTAIL.n734 185
R133 VTAIL.n654 VTAIL.n653 185
R134 VTAIL.n741 VTAIL.n740 185
R135 VTAIL.n33 VTAIL.n32 185
R136 VTAIL.n35 VTAIL.n34 185
R137 VTAIL.n28 VTAIL.n27 185
R138 VTAIL.n41 VTAIL.n40 185
R139 VTAIL.n43 VTAIL.n42 185
R140 VTAIL.n24 VTAIL.n23 185
R141 VTAIL.n50 VTAIL.n49 185
R142 VTAIL.n51 VTAIL.n22 185
R143 VTAIL.n53 VTAIL.n52 185
R144 VTAIL.n20 VTAIL.n19 185
R145 VTAIL.n59 VTAIL.n58 185
R146 VTAIL.n61 VTAIL.n60 185
R147 VTAIL.n16 VTAIL.n15 185
R148 VTAIL.n67 VTAIL.n66 185
R149 VTAIL.n69 VTAIL.n68 185
R150 VTAIL.n12 VTAIL.n11 185
R151 VTAIL.n75 VTAIL.n74 185
R152 VTAIL.n77 VTAIL.n76 185
R153 VTAIL.n8 VTAIL.n7 185
R154 VTAIL.n83 VTAIL.n82 185
R155 VTAIL.n85 VTAIL.n84 185
R156 VTAIL.n4 VTAIL.n3 185
R157 VTAIL.n91 VTAIL.n90 185
R158 VTAIL.n125 VTAIL.n124 185
R159 VTAIL.n127 VTAIL.n126 185
R160 VTAIL.n120 VTAIL.n119 185
R161 VTAIL.n133 VTAIL.n132 185
R162 VTAIL.n135 VTAIL.n134 185
R163 VTAIL.n116 VTAIL.n115 185
R164 VTAIL.n142 VTAIL.n141 185
R165 VTAIL.n143 VTAIL.n114 185
R166 VTAIL.n145 VTAIL.n144 185
R167 VTAIL.n112 VTAIL.n111 185
R168 VTAIL.n151 VTAIL.n150 185
R169 VTAIL.n153 VTAIL.n152 185
R170 VTAIL.n108 VTAIL.n107 185
R171 VTAIL.n159 VTAIL.n158 185
R172 VTAIL.n161 VTAIL.n160 185
R173 VTAIL.n104 VTAIL.n103 185
R174 VTAIL.n167 VTAIL.n166 185
R175 VTAIL.n169 VTAIL.n168 185
R176 VTAIL.n100 VTAIL.n99 185
R177 VTAIL.n175 VTAIL.n174 185
R178 VTAIL.n177 VTAIL.n176 185
R179 VTAIL.n96 VTAIL.n95 185
R180 VTAIL.n183 VTAIL.n182 185
R181 VTAIL.n219 VTAIL.n218 185
R182 VTAIL.n221 VTAIL.n220 185
R183 VTAIL.n214 VTAIL.n213 185
R184 VTAIL.n227 VTAIL.n226 185
R185 VTAIL.n229 VTAIL.n228 185
R186 VTAIL.n210 VTAIL.n209 185
R187 VTAIL.n236 VTAIL.n235 185
R188 VTAIL.n237 VTAIL.n208 185
R189 VTAIL.n239 VTAIL.n238 185
R190 VTAIL.n206 VTAIL.n205 185
R191 VTAIL.n245 VTAIL.n244 185
R192 VTAIL.n247 VTAIL.n246 185
R193 VTAIL.n202 VTAIL.n201 185
R194 VTAIL.n253 VTAIL.n252 185
R195 VTAIL.n255 VTAIL.n254 185
R196 VTAIL.n198 VTAIL.n197 185
R197 VTAIL.n261 VTAIL.n260 185
R198 VTAIL.n263 VTAIL.n262 185
R199 VTAIL.n194 VTAIL.n193 185
R200 VTAIL.n269 VTAIL.n268 185
R201 VTAIL.n271 VTAIL.n270 185
R202 VTAIL.n190 VTAIL.n189 185
R203 VTAIL.n277 VTAIL.n276 185
R204 VTAIL.n649 VTAIL.n648 185
R205 VTAIL.n562 VTAIL.n561 185
R206 VTAIL.n643 VTAIL.n642 185
R207 VTAIL.n641 VTAIL.n640 185
R208 VTAIL.n566 VTAIL.n565 185
R209 VTAIL.n635 VTAIL.n634 185
R210 VTAIL.n633 VTAIL.n632 185
R211 VTAIL.n570 VTAIL.n569 185
R212 VTAIL.n627 VTAIL.n626 185
R213 VTAIL.n625 VTAIL.n624 185
R214 VTAIL.n574 VTAIL.n573 185
R215 VTAIL.n619 VTAIL.n618 185
R216 VTAIL.n617 VTAIL.n616 185
R217 VTAIL.n578 VTAIL.n577 185
R218 VTAIL.n582 VTAIL.n580 185
R219 VTAIL.n611 VTAIL.n610 185
R220 VTAIL.n609 VTAIL.n608 185
R221 VTAIL.n584 VTAIL.n583 185
R222 VTAIL.n603 VTAIL.n602 185
R223 VTAIL.n601 VTAIL.n600 185
R224 VTAIL.n588 VTAIL.n587 185
R225 VTAIL.n595 VTAIL.n594 185
R226 VTAIL.n593 VTAIL.n592 185
R227 VTAIL.n555 VTAIL.n554 185
R228 VTAIL.n468 VTAIL.n467 185
R229 VTAIL.n549 VTAIL.n548 185
R230 VTAIL.n547 VTAIL.n546 185
R231 VTAIL.n472 VTAIL.n471 185
R232 VTAIL.n541 VTAIL.n540 185
R233 VTAIL.n539 VTAIL.n538 185
R234 VTAIL.n476 VTAIL.n475 185
R235 VTAIL.n533 VTAIL.n532 185
R236 VTAIL.n531 VTAIL.n530 185
R237 VTAIL.n480 VTAIL.n479 185
R238 VTAIL.n525 VTAIL.n524 185
R239 VTAIL.n523 VTAIL.n522 185
R240 VTAIL.n484 VTAIL.n483 185
R241 VTAIL.n488 VTAIL.n486 185
R242 VTAIL.n517 VTAIL.n516 185
R243 VTAIL.n515 VTAIL.n514 185
R244 VTAIL.n490 VTAIL.n489 185
R245 VTAIL.n509 VTAIL.n508 185
R246 VTAIL.n507 VTAIL.n506 185
R247 VTAIL.n494 VTAIL.n493 185
R248 VTAIL.n501 VTAIL.n500 185
R249 VTAIL.n499 VTAIL.n498 185
R250 VTAIL.n463 VTAIL.n462 185
R251 VTAIL.n376 VTAIL.n375 185
R252 VTAIL.n457 VTAIL.n456 185
R253 VTAIL.n455 VTAIL.n454 185
R254 VTAIL.n380 VTAIL.n379 185
R255 VTAIL.n449 VTAIL.n448 185
R256 VTAIL.n447 VTAIL.n446 185
R257 VTAIL.n384 VTAIL.n383 185
R258 VTAIL.n441 VTAIL.n440 185
R259 VTAIL.n439 VTAIL.n438 185
R260 VTAIL.n388 VTAIL.n387 185
R261 VTAIL.n433 VTAIL.n432 185
R262 VTAIL.n431 VTAIL.n430 185
R263 VTAIL.n392 VTAIL.n391 185
R264 VTAIL.n396 VTAIL.n394 185
R265 VTAIL.n425 VTAIL.n424 185
R266 VTAIL.n423 VTAIL.n422 185
R267 VTAIL.n398 VTAIL.n397 185
R268 VTAIL.n417 VTAIL.n416 185
R269 VTAIL.n415 VTAIL.n414 185
R270 VTAIL.n402 VTAIL.n401 185
R271 VTAIL.n409 VTAIL.n408 185
R272 VTAIL.n407 VTAIL.n406 185
R273 VTAIL.n369 VTAIL.n368 185
R274 VTAIL.n282 VTAIL.n281 185
R275 VTAIL.n363 VTAIL.n362 185
R276 VTAIL.n361 VTAIL.n360 185
R277 VTAIL.n286 VTAIL.n285 185
R278 VTAIL.n355 VTAIL.n354 185
R279 VTAIL.n353 VTAIL.n352 185
R280 VTAIL.n290 VTAIL.n289 185
R281 VTAIL.n347 VTAIL.n346 185
R282 VTAIL.n345 VTAIL.n344 185
R283 VTAIL.n294 VTAIL.n293 185
R284 VTAIL.n339 VTAIL.n338 185
R285 VTAIL.n337 VTAIL.n336 185
R286 VTAIL.n298 VTAIL.n297 185
R287 VTAIL.n302 VTAIL.n300 185
R288 VTAIL.n331 VTAIL.n330 185
R289 VTAIL.n329 VTAIL.n328 185
R290 VTAIL.n304 VTAIL.n303 185
R291 VTAIL.n323 VTAIL.n322 185
R292 VTAIL.n321 VTAIL.n320 185
R293 VTAIL.n308 VTAIL.n307 185
R294 VTAIL.n315 VTAIL.n314 185
R295 VTAIL.n313 VTAIL.n312 185
R296 VTAIL.n681 VTAIL.t8 149.524
R297 VTAIL.n31 VTAIL.t14 149.524
R298 VTAIL.n123 VTAIL.t6 149.524
R299 VTAIL.n217 VTAIL.t3 149.524
R300 VTAIL.n591 VTAIL.t1 149.524
R301 VTAIL.n497 VTAIL.t5 149.524
R302 VTAIL.n405 VTAIL.t9 149.524
R303 VTAIL.n311 VTAIL.t12 149.524
R304 VTAIL.n684 VTAIL.n683 104.615
R305 VTAIL.n684 VTAIL.n677 104.615
R306 VTAIL.n691 VTAIL.n677 104.615
R307 VTAIL.n692 VTAIL.n691 104.615
R308 VTAIL.n692 VTAIL.n673 104.615
R309 VTAIL.n700 VTAIL.n673 104.615
R310 VTAIL.n701 VTAIL.n700 104.615
R311 VTAIL.n702 VTAIL.n701 104.615
R312 VTAIL.n702 VTAIL.n669 104.615
R313 VTAIL.n709 VTAIL.n669 104.615
R314 VTAIL.n710 VTAIL.n709 104.615
R315 VTAIL.n710 VTAIL.n665 104.615
R316 VTAIL.n717 VTAIL.n665 104.615
R317 VTAIL.n718 VTAIL.n717 104.615
R318 VTAIL.n718 VTAIL.n661 104.615
R319 VTAIL.n725 VTAIL.n661 104.615
R320 VTAIL.n726 VTAIL.n725 104.615
R321 VTAIL.n726 VTAIL.n657 104.615
R322 VTAIL.n733 VTAIL.n657 104.615
R323 VTAIL.n734 VTAIL.n733 104.615
R324 VTAIL.n734 VTAIL.n653 104.615
R325 VTAIL.n741 VTAIL.n653 104.615
R326 VTAIL.n34 VTAIL.n33 104.615
R327 VTAIL.n34 VTAIL.n27 104.615
R328 VTAIL.n41 VTAIL.n27 104.615
R329 VTAIL.n42 VTAIL.n41 104.615
R330 VTAIL.n42 VTAIL.n23 104.615
R331 VTAIL.n50 VTAIL.n23 104.615
R332 VTAIL.n51 VTAIL.n50 104.615
R333 VTAIL.n52 VTAIL.n51 104.615
R334 VTAIL.n52 VTAIL.n19 104.615
R335 VTAIL.n59 VTAIL.n19 104.615
R336 VTAIL.n60 VTAIL.n59 104.615
R337 VTAIL.n60 VTAIL.n15 104.615
R338 VTAIL.n67 VTAIL.n15 104.615
R339 VTAIL.n68 VTAIL.n67 104.615
R340 VTAIL.n68 VTAIL.n11 104.615
R341 VTAIL.n75 VTAIL.n11 104.615
R342 VTAIL.n76 VTAIL.n75 104.615
R343 VTAIL.n76 VTAIL.n7 104.615
R344 VTAIL.n83 VTAIL.n7 104.615
R345 VTAIL.n84 VTAIL.n83 104.615
R346 VTAIL.n84 VTAIL.n3 104.615
R347 VTAIL.n91 VTAIL.n3 104.615
R348 VTAIL.n126 VTAIL.n125 104.615
R349 VTAIL.n126 VTAIL.n119 104.615
R350 VTAIL.n133 VTAIL.n119 104.615
R351 VTAIL.n134 VTAIL.n133 104.615
R352 VTAIL.n134 VTAIL.n115 104.615
R353 VTAIL.n142 VTAIL.n115 104.615
R354 VTAIL.n143 VTAIL.n142 104.615
R355 VTAIL.n144 VTAIL.n143 104.615
R356 VTAIL.n144 VTAIL.n111 104.615
R357 VTAIL.n151 VTAIL.n111 104.615
R358 VTAIL.n152 VTAIL.n151 104.615
R359 VTAIL.n152 VTAIL.n107 104.615
R360 VTAIL.n159 VTAIL.n107 104.615
R361 VTAIL.n160 VTAIL.n159 104.615
R362 VTAIL.n160 VTAIL.n103 104.615
R363 VTAIL.n167 VTAIL.n103 104.615
R364 VTAIL.n168 VTAIL.n167 104.615
R365 VTAIL.n168 VTAIL.n99 104.615
R366 VTAIL.n175 VTAIL.n99 104.615
R367 VTAIL.n176 VTAIL.n175 104.615
R368 VTAIL.n176 VTAIL.n95 104.615
R369 VTAIL.n183 VTAIL.n95 104.615
R370 VTAIL.n220 VTAIL.n219 104.615
R371 VTAIL.n220 VTAIL.n213 104.615
R372 VTAIL.n227 VTAIL.n213 104.615
R373 VTAIL.n228 VTAIL.n227 104.615
R374 VTAIL.n228 VTAIL.n209 104.615
R375 VTAIL.n236 VTAIL.n209 104.615
R376 VTAIL.n237 VTAIL.n236 104.615
R377 VTAIL.n238 VTAIL.n237 104.615
R378 VTAIL.n238 VTAIL.n205 104.615
R379 VTAIL.n245 VTAIL.n205 104.615
R380 VTAIL.n246 VTAIL.n245 104.615
R381 VTAIL.n246 VTAIL.n201 104.615
R382 VTAIL.n253 VTAIL.n201 104.615
R383 VTAIL.n254 VTAIL.n253 104.615
R384 VTAIL.n254 VTAIL.n197 104.615
R385 VTAIL.n261 VTAIL.n197 104.615
R386 VTAIL.n262 VTAIL.n261 104.615
R387 VTAIL.n262 VTAIL.n193 104.615
R388 VTAIL.n269 VTAIL.n193 104.615
R389 VTAIL.n270 VTAIL.n269 104.615
R390 VTAIL.n270 VTAIL.n189 104.615
R391 VTAIL.n277 VTAIL.n189 104.615
R392 VTAIL.n649 VTAIL.n561 104.615
R393 VTAIL.n642 VTAIL.n561 104.615
R394 VTAIL.n642 VTAIL.n641 104.615
R395 VTAIL.n641 VTAIL.n565 104.615
R396 VTAIL.n634 VTAIL.n565 104.615
R397 VTAIL.n634 VTAIL.n633 104.615
R398 VTAIL.n633 VTAIL.n569 104.615
R399 VTAIL.n626 VTAIL.n569 104.615
R400 VTAIL.n626 VTAIL.n625 104.615
R401 VTAIL.n625 VTAIL.n573 104.615
R402 VTAIL.n618 VTAIL.n573 104.615
R403 VTAIL.n618 VTAIL.n617 104.615
R404 VTAIL.n617 VTAIL.n577 104.615
R405 VTAIL.n582 VTAIL.n577 104.615
R406 VTAIL.n610 VTAIL.n582 104.615
R407 VTAIL.n610 VTAIL.n609 104.615
R408 VTAIL.n609 VTAIL.n583 104.615
R409 VTAIL.n602 VTAIL.n583 104.615
R410 VTAIL.n602 VTAIL.n601 104.615
R411 VTAIL.n601 VTAIL.n587 104.615
R412 VTAIL.n594 VTAIL.n587 104.615
R413 VTAIL.n594 VTAIL.n593 104.615
R414 VTAIL.n555 VTAIL.n467 104.615
R415 VTAIL.n548 VTAIL.n467 104.615
R416 VTAIL.n548 VTAIL.n547 104.615
R417 VTAIL.n547 VTAIL.n471 104.615
R418 VTAIL.n540 VTAIL.n471 104.615
R419 VTAIL.n540 VTAIL.n539 104.615
R420 VTAIL.n539 VTAIL.n475 104.615
R421 VTAIL.n532 VTAIL.n475 104.615
R422 VTAIL.n532 VTAIL.n531 104.615
R423 VTAIL.n531 VTAIL.n479 104.615
R424 VTAIL.n524 VTAIL.n479 104.615
R425 VTAIL.n524 VTAIL.n523 104.615
R426 VTAIL.n523 VTAIL.n483 104.615
R427 VTAIL.n488 VTAIL.n483 104.615
R428 VTAIL.n516 VTAIL.n488 104.615
R429 VTAIL.n516 VTAIL.n515 104.615
R430 VTAIL.n515 VTAIL.n489 104.615
R431 VTAIL.n508 VTAIL.n489 104.615
R432 VTAIL.n508 VTAIL.n507 104.615
R433 VTAIL.n507 VTAIL.n493 104.615
R434 VTAIL.n500 VTAIL.n493 104.615
R435 VTAIL.n500 VTAIL.n499 104.615
R436 VTAIL.n463 VTAIL.n375 104.615
R437 VTAIL.n456 VTAIL.n375 104.615
R438 VTAIL.n456 VTAIL.n455 104.615
R439 VTAIL.n455 VTAIL.n379 104.615
R440 VTAIL.n448 VTAIL.n379 104.615
R441 VTAIL.n448 VTAIL.n447 104.615
R442 VTAIL.n447 VTAIL.n383 104.615
R443 VTAIL.n440 VTAIL.n383 104.615
R444 VTAIL.n440 VTAIL.n439 104.615
R445 VTAIL.n439 VTAIL.n387 104.615
R446 VTAIL.n432 VTAIL.n387 104.615
R447 VTAIL.n432 VTAIL.n431 104.615
R448 VTAIL.n431 VTAIL.n391 104.615
R449 VTAIL.n396 VTAIL.n391 104.615
R450 VTAIL.n424 VTAIL.n396 104.615
R451 VTAIL.n424 VTAIL.n423 104.615
R452 VTAIL.n423 VTAIL.n397 104.615
R453 VTAIL.n416 VTAIL.n397 104.615
R454 VTAIL.n416 VTAIL.n415 104.615
R455 VTAIL.n415 VTAIL.n401 104.615
R456 VTAIL.n408 VTAIL.n401 104.615
R457 VTAIL.n408 VTAIL.n407 104.615
R458 VTAIL.n369 VTAIL.n281 104.615
R459 VTAIL.n362 VTAIL.n281 104.615
R460 VTAIL.n362 VTAIL.n361 104.615
R461 VTAIL.n361 VTAIL.n285 104.615
R462 VTAIL.n354 VTAIL.n285 104.615
R463 VTAIL.n354 VTAIL.n353 104.615
R464 VTAIL.n353 VTAIL.n289 104.615
R465 VTAIL.n346 VTAIL.n289 104.615
R466 VTAIL.n346 VTAIL.n345 104.615
R467 VTAIL.n345 VTAIL.n293 104.615
R468 VTAIL.n338 VTAIL.n293 104.615
R469 VTAIL.n338 VTAIL.n337 104.615
R470 VTAIL.n337 VTAIL.n297 104.615
R471 VTAIL.n302 VTAIL.n297 104.615
R472 VTAIL.n330 VTAIL.n302 104.615
R473 VTAIL.n330 VTAIL.n329 104.615
R474 VTAIL.n329 VTAIL.n303 104.615
R475 VTAIL.n322 VTAIL.n303 104.615
R476 VTAIL.n322 VTAIL.n321 104.615
R477 VTAIL.n321 VTAIL.n307 104.615
R478 VTAIL.n314 VTAIL.n307 104.615
R479 VTAIL.n314 VTAIL.n313 104.615
R480 VTAIL.n683 VTAIL.t8 52.3082
R481 VTAIL.n33 VTAIL.t14 52.3082
R482 VTAIL.n125 VTAIL.t6 52.3082
R483 VTAIL.n219 VTAIL.t3 52.3082
R484 VTAIL.n593 VTAIL.t1 52.3082
R485 VTAIL.n499 VTAIL.t5 52.3082
R486 VTAIL.n407 VTAIL.t9 52.3082
R487 VTAIL.n313 VTAIL.t12 52.3082
R488 VTAIL.n559 VTAIL.n558 47.5752
R489 VTAIL.n373 VTAIL.n372 47.5752
R490 VTAIL.n1 VTAIL.n0 47.5751
R491 VTAIL.n187 VTAIL.n186 47.5751
R492 VTAIL.n743 VTAIL.n742 33.7369
R493 VTAIL.n93 VTAIL.n92 33.7369
R494 VTAIL.n185 VTAIL.n184 33.7369
R495 VTAIL.n279 VTAIL.n278 33.7369
R496 VTAIL.n651 VTAIL.n650 33.7369
R497 VTAIL.n557 VTAIL.n556 33.7369
R498 VTAIL.n465 VTAIL.n464 33.7369
R499 VTAIL.n371 VTAIL.n370 33.7369
R500 VTAIL.n743 VTAIL.n651 29.7893
R501 VTAIL.n371 VTAIL.n279 29.7893
R502 VTAIL.n703 VTAIL.n670 13.1884
R503 VTAIL.n53 VTAIL.n20 13.1884
R504 VTAIL.n145 VTAIL.n112 13.1884
R505 VTAIL.n239 VTAIL.n206 13.1884
R506 VTAIL.n580 VTAIL.n578 13.1884
R507 VTAIL.n486 VTAIL.n484 13.1884
R508 VTAIL.n394 VTAIL.n392 13.1884
R509 VTAIL.n300 VTAIL.n298 13.1884
R510 VTAIL.n704 VTAIL.n672 12.8005
R511 VTAIL.n708 VTAIL.n707 12.8005
R512 VTAIL.n54 VTAIL.n22 12.8005
R513 VTAIL.n58 VTAIL.n57 12.8005
R514 VTAIL.n146 VTAIL.n114 12.8005
R515 VTAIL.n150 VTAIL.n149 12.8005
R516 VTAIL.n240 VTAIL.n208 12.8005
R517 VTAIL.n244 VTAIL.n243 12.8005
R518 VTAIL.n616 VTAIL.n615 12.8005
R519 VTAIL.n612 VTAIL.n611 12.8005
R520 VTAIL.n522 VTAIL.n521 12.8005
R521 VTAIL.n518 VTAIL.n517 12.8005
R522 VTAIL.n430 VTAIL.n429 12.8005
R523 VTAIL.n426 VTAIL.n425 12.8005
R524 VTAIL.n336 VTAIL.n335 12.8005
R525 VTAIL.n332 VTAIL.n331 12.8005
R526 VTAIL.n699 VTAIL.n698 12.0247
R527 VTAIL.n711 VTAIL.n668 12.0247
R528 VTAIL.n49 VTAIL.n48 12.0247
R529 VTAIL.n61 VTAIL.n18 12.0247
R530 VTAIL.n141 VTAIL.n140 12.0247
R531 VTAIL.n153 VTAIL.n110 12.0247
R532 VTAIL.n235 VTAIL.n234 12.0247
R533 VTAIL.n247 VTAIL.n204 12.0247
R534 VTAIL.n619 VTAIL.n576 12.0247
R535 VTAIL.n608 VTAIL.n581 12.0247
R536 VTAIL.n525 VTAIL.n482 12.0247
R537 VTAIL.n514 VTAIL.n487 12.0247
R538 VTAIL.n433 VTAIL.n390 12.0247
R539 VTAIL.n422 VTAIL.n395 12.0247
R540 VTAIL.n339 VTAIL.n296 12.0247
R541 VTAIL.n328 VTAIL.n301 12.0247
R542 VTAIL.n697 VTAIL.n674 11.249
R543 VTAIL.n712 VTAIL.n666 11.249
R544 VTAIL.n47 VTAIL.n24 11.249
R545 VTAIL.n62 VTAIL.n16 11.249
R546 VTAIL.n139 VTAIL.n116 11.249
R547 VTAIL.n154 VTAIL.n108 11.249
R548 VTAIL.n233 VTAIL.n210 11.249
R549 VTAIL.n248 VTAIL.n202 11.249
R550 VTAIL.n620 VTAIL.n574 11.249
R551 VTAIL.n607 VTAIL.n584 11.249
R552 VTAIL.n526 VTAIL.n480 11.249
R553 VTAIL.n513 VTAIL.n490 11.249
R554 VTAIL.n434 VTAIL.n388 11.249
R555 VTAIL.n421 VTAIL.n398 11.249
R556 VTAIL.n340 VTAIL.n294 11.249
R557 VTAIL.n327 VTAIL.n304 11.249
R558 VTAIL.n694 VTAIL.n693 10.4732
R559 VTAIL.n716 VTAIL.n715 10.4732
R560 VTAIL.n740 VTAIL.n652 10.4732
R561 VTAIL.n44 VTAIL.n43 10.4732
R562 VTAIL.n66 VTAIL.n65 10.4732
R563 VTAIL.n90 VTAIL.n2 10.4732
R564 VTAIL.n136 VTAIL.n135 10.4732
R565 VTAIL.n158 VTAIL.n157 10.4732
R566 VTAIL.n182 VTAIL.n94 10.4732
R567 VTAIL.n230 VTAIL.n229 10.4732
R568 VTAIL.n252 VTAIL.n251 10.4732
R569 VTAIL.n276 VTAIL.n188 10.4732
R570 VTAIL.n648 VTAIL.n560 10.4732
R571 VTAIL.n624 VTAIL.n623 10.4732
R572 VTAIL.n604 VTAIL.n603 10.4732
R573 VTAIL.n554 VTAIL.n466 10.4732
R574 VTAIL.n530 VTAIL.n529 10.4732
R575 VTAIL.n510 VTAIL.n509 10.4732
R576 VTAIL.n462 VTAIL.n374 10.4732
R577 VTAIL.n438 VTAIL.n437 10.4732
R578 VTAIL.n418 VTAIL.n417 10.4732
R579 VTAIL.n368 VTAIL.n280 10.4732
R580 VTAIL.n344 VTAIL.n343 10.4732
R581 VTAIL.n324 VTAIL.n323 10.4732
R582 VTAIL.n682 VTAIL.n681 10.2747
R583 VTAIL.n32 VTAIL.n31 10.2747
R584 VTAIL.n124 VTAIL.n123 10.2747
R585 VTAIL.n218 VTAIL.n217 10.2747
R586 VTAIL.n592 VTAIL.n591 10.2747
R587 VTAIL.n498 VTAIL.n497 10.2747
R588 VTAIL.n406 VTAIL.n405 10.2747
R589 VTAIL.n312 VTAIL.n311 10.2747
R590 VTAIL.n690 VTAIL.n676 9.69747
R591 VTAIL.n719 VTAIL.n664 9.69747
R592 VTAIL.n739 VTAIL.n654 9.69747
R593 VTAIL.n40 VTAIL.n26 9.69747
R594 VTAIL.n69 VTAIL.n14 9.69747
R595 VTAIL.n89 VTAIL.n4 9.69747
R596 VTAIL.n132 VTAIL.n118 9.69747
R597 VTAIL.n161 VTAIL.n106 9.69747
R598 VTAIL.n181 VTAIL.n96 9.69747
R599 VTAIL.n226 VTAIL.n212 9.69747
R600 VTAIL.n255 VTAIL.n200 9.69747
R601 VTAIL.n275 VTAIL.n190 9.69747
R602 VTAIL.n647 VTAIL.n562 9.69747
R603 VTAIL.n627 VTAIL.n572 9.69747
R604 VTAIL.n600 VTAIL.n586 9.69747
R605 VTAIL.n553 VTAIL.n468 9.69747
R606 VTAIL.n533 VTAIL.n478 9.69747
R607 VTAIL.n506 VTAIL.n492 9.69747
R608 VTAIL.n461 VTAIL.n376 9.69747
R609 VTAIL.n441 VTAIL.n386 9.69747
R610 VTAIL.n414 VTAIL.n400 9.69747
R611 VTAIL.n367 VTAIL.n282 9.69747
R612 VTAIL.n347 VTAIL.n292 9.69747
R613 VTAIL.n320 VTAIL.n306 9.69747
R614 VTAIL.n738 VTAIL.n652 9.45567
R615 VTAIL.n88 VTAIL.n2 9.45567
R616 VTAIL.n180 VTAIL.n94 9.45567
R617 VTAIL.n274 VTAIL.n188 9.45567
R618 VTAIL.n646 VTAIL.n560 9.45567
R619 VTAIL.n552 VTAIL.n466 9.45567
R620 VTAIL.n460 VTAIL.n374 9.45567
R621 VTAIL.n366 VTAIL.n280 9.45567
R622 VTAIL.n729 VTAIL.n728 9.3005
R623 VTAIL.n731 VTAIL.n730 9.3005
R624 VTAIL.n656 VTAIL.n655 9.3005
R625 VTAIL.n737 VTAIL.n736 9.3005
R626 VTAIL.n739 VTAIL.n738 9.3005
R627 VTAIL.n723 VTAIL.n722 9.3005
R628 VTAIL.n721 VTAIL.n720 9.3005
R629 VTAIL.n664 VTAIL.n663 9.3005
R630 VTAIL.n715 VTAIL.n714 9.3005
R631 VTAIL.n713 VTAIL.n712 9.3005
R632 VTAIL.n668 VTAIL.n667 9.3005
R633 VTAIL.n707 VTAIL.n706 9.3005
R634 VTAIL.n680 VTAIL.n679 9.3005
R635 VTAIL.n687 VTAIL.n686 9.3005
R636 VTAIL.n689 VTAIL.n688 9.3005
R637 VTAIL.n676 VTAIL.n675 9.3005
R638 VTAIL.n695 VTAIL.n694 9.3005
R639 VTAIL.n697 VTAIL.n696 9.3005
R640 VTAIL.n698 VTAIL.n671 9.3005
R641 VTAIL.n705 VTAIL.n704 9.3005
R642 VTAIL.n660 VTAIL.n659 9.3005
R643 VTAIL.n79 VTAIL.n78 9.3005
R644 VTAIL.n81 VTAIL.n80 9.3005
R645 VTAIL.n6 VTAIL.n5 9.3005
R646 VTAIL.n87 VTAIL.n86 9.3005
R647 VTAIL.n89 VTAIL.n88 9.3005
R648 VTAIL.n73 VTAIL.n72 9.3005
R649 VTAIL.n71 VTAIL.n70 9.3005
R650 VTAIL.n14 VTAIL.n13 9.3005
R651 VTAIL.n65 VTAIL.n64 9.3005
R652 VTAIL.n63 VTAIL.n62 9.3005
R653 VTAIL.n18 VTAIL.n17 9.3005
R654 VTAIL.n57 VTAIL.n56 9.3005
R655 VTAIL.n30 VTAIL.n29 9.3005
R656 VTAIL.n37 VTAIL.n36 9.3005
R657 VTAIL.n39 VTAIL.n38 9.3005
R658 VTAIL.n26 VTAIL.n25 9.3005
R659 VTAIL.n45 VTAIL.n44 9.3005
R660 VTAIL.n47 VTAIL.n46 9.3005
R661 VTAIL.n48 VTAIL.n21 9.3005
R662 VTAIL.n55 VTAIL.n54 9.3005
R663 VTAIL.n10 VTAIL.n9 9.3005
R664 VTAIL.n171 VTAIL.n170 9.3005
R665 VTAIL.n173 VTAIL.n172 9.3005
R666 VTAIL.n98 VTAIL.n97 9.3005
R667 VTAIL.n179 VTAIL.n178 9.3005
R668 VTAIL.n181 VTAIL.n180 9.3005
R669 VTAIL.n165 VTAIL.n164 9.3005
R670 VTAIL.n163 VTAIL.n162 9.3005
R671 VTAIL.n106 VTAIL.n105 9.3005
R672 VTAIL.n157 VTAIL.n156 9.3005
R673 VTAIL.n155 VTAIL.n154 9.3005
R674 VTAIL.n110 VTAIL.n109 9.3005
R675 VTAIL.n149 VTAIL.n148 9.3005
R676 VTAIL.n122 VTAIL.n121 9.3005
R677 VTAIL.n129 VTAIL.n128 9.3005
R678 VTAIL.n131 VTAIL.n130 9.3005
R679 VTAIL.n118 VTAIL.n117 9.3005
R680 VTAIL.n137 VTAIL.n136 9.3005
R681 VTAIL.n139 VTAIL.n138 9.3005
R682 VTAIL.n140 VTAIL.n113 9.3005
R683 VTAIL.n147 VTAIL.n146 9.3005
R684 VTAIL.n102 VTAIL.n101 9.3005
R685 VTAIL.n265 VTAIL.n264 9.3005
R686 VTAIL.n267 VTAIL.n266 9.3005
R687 VTAIL.n192 VTAIL.n191 9.3005
R688 VTAIL.n273 VTAIL.n272 9.3005
R689 VTAIL.n275 VTAIL.n274 9.3005
R690 VTAIL.n259 VTAIL.n258 9.3005
R691 VTAIL.n257 VTAIL.n256 9.3005
R692 VTAIL.n200 VTAIL.n199 9.3005
R693 VTAIL.n251 VTAIL.n250 9.3005
R694 VTAIL.n249 VTAIL.n248 9.3005
R695 VTAIL.n204 VTAIL.n203 9.3005
R696 VTAIL.n243 VTAIL.n242 9.3005
R697 VTAIL.n216 VTAIL.n215 9.3005
R698 VTAIL.n223 VTAIL.n222 9.3005
R699 VTAIL.n225 VTAIL.n224 9.3005
R700 VTAIL.n212 VTAIL.n211 9.3005
R701 VTAIL.n231 VTAIL.n230 9.3005
R702 VTAIL.n233 VTAIL.n232 9.3005
R703 VTAIL.n234 VTAIL.n207 9.3005
R704 VTAIL.n241 VTAIL.n240 9.3005
R705 VTAIL.n196 VTAIL.n195 9.3005
R706 VTAIL.n647 VTAIL.n646 9.3005
R707 VTAIL.n645 VTAIL.n644 9.3005
R708 VTAIL.n564 VTAIL.n563 9.3005
R709 VTAIL.n639 VTAIL.n638 9.3005
R710 VTAIL.n637 VTAIL.n636 9.3005
R711 VTAIL.n568 VTAIL.n567 9.3005
R712 VTAIL.n631 VTAIL.n630 9.3005
R713 VTAIL.n629 VTAIL.n628 9.3005
R714 VTAIL.n572 VTAIL.n571 9.3005
R715 VTAIL.n623 VTAIL.n622 9.3005
R716 VTAIL.n621 VTAIL.n620 9.3005
R717 VTAIL.n576 VTAIL.n575 9.3005
R718 VTAIL.n615 VTAIL.n614 9.3005
R719 VTAIL.n613 VTAIL.n612 9.3005
R720 VTAIL.n581 VTAIL.n579 9.3005
R721 VTAIL.n607 VTAIL.n606 9.3005
R722 VTAIL.n605 VTAIL.n604 9.3005
R723 VTAIL.n586 VTAIL.n585 9.3005
R724 VTAIL.n599 VTAIL.n598 9.3005
R725 VTAIL.n597 VTAIL.n596 9.3005
R726 VTAIL.n590 VTAIL.n589 9.3005
R727 VTAIL.n496 VTAIL.n495 9.3005
R728 VTAIL.n503 VTAIL.n502 9.3005
R729 VTAIL.n505 VTAIL.n504 9.3005
R730 VTAIL.n492 VTAIL.n491 9.3005
R731 VTAIL.n511 VTAIL.n510 9.3005
R732 VTAIL.n513 VTAIL.n512 9.3005
R733 VTAIL.n487 VTAIL.n485 9.3005
R734 VTAIL.n519 VTAIL.n518 9.3005
R735 VTAIL.n545 VTAIL.n544 9.3005
R736 VTAIL.n470 VTAIL.n469 9.3005
R737 VTAIL.n551 VTAIL.n550 9.3005
R738 VTAIL.n553 VTAIL.n552 9.3005
R739 VTAIL.n543 VTAIL.n542 9.3005
R740 VTAIL.n474 VTAIL.n473 9.3005
R741 VTAIL.n537 VTAIL.n536 9.3005
R742 VTAIL.n535 VTAIL.n534 9.3005
R743 VTAIL.n478 VTAIL.n477 9.3005
R744 VTAIL.n529 VTAIL.n528 9.3005
R745 VTAIL.n527 VTAIL.n526 9.3005
R746 VTAIL.n482 VTAIL.n481 9.3005
R747 VTAIL.n521 VTAIL.n520 9.3005
R748 VTAIL.n404 VTAIL.n403 9.3005
R749 VTAIL.n411 VTAIL.n410 9.3005
R750 VTAIL.n413 VTAIL.n412 9.3005
R751 VTAIL.n400 VTAIL.n399 9.3005
R752 VTAIL.n419 VTAIL.n418 9.3005
R753 VTAIL.n421 VTAIL.n420 9.3005
R754 VTAIL.n395 VTAIL.n393 9.3005
R755 VTAIL.n427 VTAIL.n426 9.3005
R756 VTAIL.n453 VTAIL.n452 9.3005
R757 VTAIL.n378 VTAIL.n377 9.3005
R758 VTAIL.n459 VTAIL.n458 9.3005
R759 VTAIL.n461 VTAIL.n460 9.3005
R760 VTAIL.n451 VTAIL.n450 9.3005
R761 VTAIL.n382 VTAIL.n381 9.3005
R762 VTAIL.n445 VTAIL.n444 9.3005
R763 VTAIL.n443 VTAIL.n442 9.3005
R764 VTAIL.n386 VTAIL.n385 9.3005
R765 VTAIL.n437 VTAIL.n436 9.3005
R766 VTAIL.n435 VTAIL.n434 9.3005
R767 VTAIL.n390 VTAIL.n389 9.3005
R768 VTAIL.n429 VTAIL.n428 9.3005
R769 VTAIL.n310 VTAIL.n309 9.3005
R770 VTAIL.n317 VTAIL.n316 9.3005
R771 VTAIL.n319 VTAIL.n318 9.3005
R772 VTAIL.n306 VTAIL.n305 9.3005
R773 VTAIL.n325 VTAIL.n324 9.3005
R774 VTAIL.n327 VTAIL.n326 9.3005
R775 VTAIL.n301 VTAIL.n299 9.3005
R776 VTAIL.n333 VTAIL.n332 9.3005
R777 VTAIL.n359 VTAIL.n358 9.3005
R778 VTAIL.n284 VTAIL.n283 9.3005
R779 VTAIL.n365 VTAIL.n364 9.3005
R780 VTAIL.n367 VTAIL.n366 9.3005
R781 VTAIL.n357 VTAIL.n356 9.3005
R782 VTAIL.n288 VTAIL.n287 9.3005
R783 VTAIL.n351 VTAIL.n350 9.3005
R784 VTAIL.n349 VTAIL.n348 9.3005
R785 VTAIL.n292 VTAIL.n291 9.3005
R786 VTAIL.n343 VTAIL.n342 9.3005
R787 VTAIL.n341 VTAIL.n340 9.3005
R788 VTAIL.n296 VTAIL.n295 9.3005
R789 VTAIL.n335 VTAIL.n334 9.3005
R790 VTAIL.n689 VTAIL.n678 8.92171
R791 VTAIL.n720 VTAIL.n662 8.92171
R792 VTAIL.n736 VTAIL.n735 8.92171
R793 VTAIL.n39 VTAIL.n28 8.92171
R794 VTAIL.n70 VTAIL.n12 8.92171
R795 VTAIL.n86 VTAIL.n85 8.92171
R796 VTAIL.n131 VTAIL.n120 8.92171
R797 VTAIL.n162 VTAIL.n104 8.92171
R798 VTAIL.n178 VTAIL.n177 8.92171
R799 VTAIL.n225 VTAIL.n214 8.92171
R800 VTAIL.n256 VTAIL.n198 8.92171
R801 VTAIL.n272 VTAIL.n271 8.92171
R802 VTAIL.n644 VTAIL.n643 8.92171
R803 VTAIL.n628 VTAIL.n570 8.92171
R804 VTAIL.n599 VTAIL.n588 8.92171
R805 VTAIL.n550 VTAIL.n549 8.92171
R806 VTAIL.n534 VTAIL.n476 8.92171
R807 VTAIL.n505 VTAIL.n494 8.92171
R808 VTAIL.n458 VTAIL.n457 8.92171
R809 VTAIL.n442 VTAIL.n384 8.92171
R810 VTAIL.n413 VTAIL.n402 8.92171
R811 VTAIL.n364 VTAIL.n363 8.92171
R812 VTAIL.n348 VTAIL.n290 8.92171
R813 VTAIL.n319 VTAIL.n308 8.92171
R814 VTAIL.n686 VTAIL.n685 8.14595
R815 VTAIL.n724 VTAIL.n723 8.14595
R816 VTAIL.n732 VTAIL.n656 8.14595
R817 VTAIL.n36 VTAIL.n35 8.14595
R818 VTAIL.n74 VTAIL.n73 8.14595
R819 VTAIL.n82 VTAIL.n6 8.14595
R820 VTAIL.n128 VTAIL.n127 8.14595
R821 VTAIL.n166 VTAIL.n165 8.14595
R822 VTAIL.n174 VTAIL.n98 8.14595
R823 VTAIL.n222 VTAIL.n221 8.14595
R824 VTAIL.n260 VTAIL.n259 8.14595
R825 VTAIL.n268 VTAIL.n192 8.14595
R826 VTAIL.n640 VTAIL.n564 8.14595
R827 VTAIL.n632 VTAIL.n631 8.14595
R828 VTAIL.n596 VTAIL.n595 8.14595
R829 VTAIL.n546 VTAIL.n470 8.14595
R830 VTAIL.n538 VTAIL.n537 8.14595
R831 VTAIL.n502 VTAIL.n501 8.14595
R832 VTAIL.n454 VTAIL.n378 8.14595
R833 VTAIL.n446 VTAIL.n445 8.14595
R834 VTAIL.n410 VTAIL.n409 8.14595
R835 VTAIL.n360 VTAIL.n284 8.14595
R836 VTAIL.n352 VTAIL.n351 8.14595
R837 VTAIL.n316 VTAIL.n315 8.14595
R838 VTAIL.n682 VTAIL.n680 7.3702
R839 VTAIL.n727 VTAIL.n660 7.3702
R840 VTAIL.n731 VTAIL.n658 7.3702
R841 VTAIL.n32 VTAIL.n30 7.3702
R842 VTAIL.n77 VTAIL.n10 7.3702
R843 VTAIL.n81 VTAIL.n8 7.3702
R844 VTAIL.n124 VTAIL.n122 7.3702
R845 VTAIL.n169 VTAIL.n102 7.3702
R846 VTAIL.n173 VTAIL.n100 7.3702
R847 VTAIL.n218 VTAIL.n216 7.3702
R848 VTAIL.n263 VTAIL.n196 7.3702
R849 VTAIL.n267 VTAIL.n194 7.3702
R850 VTAIL.n639 VTAIL.n566 7.3702
R851 VTAIL.n635 VTAIL.n568 7.3702
R852 VTAIL.n592 VTAIL.n590 7.3702
R853 VTAIL.n545 VTAIL.n472 7.3702
R854 VTAIL.n541 VTAIL.n474 7.3702
R855 VTAIL.n498 VTAIL.n496 7.3702
R856 VTAIL.n453 VTAIL.n380 7.3702
R857 VTAIL.n449 VTAIL.n382 7.3702
R858 VTAIL.n406 VTAIL.n404 7.3702
R859 VTAIL.n359 VTAIL.n286 7.3702
R860 VTAIL.n355 VTAIL.n288 7.3702
R861 VTAIL.n312 VTAIL.n310 7.3702
R862 VTAIL.n728 VTAIL.n727 6.59444
R863 VTAIL.n728 VTAIL.n658 6.59444
R864 VTAIL.n78 VTAIL.n77 6.59444
R865 VTAIL.n78 VTAIL.n8 6.59444
R866 VTAIL.n170 VTAIL.n169 6.59444
R867 VTAIL.n170 VTAIL.n100 6.59444
R868 VTAIL.n264 VTAIL.n263 6.59444
R869 VTAIL.n264 VTAIL.n194 6.59444
R870 VTAIL.n636 VTAIL.n566 6.59444
R871 VTAIL.n636 VTAIL.n635 6.59444
R872 VTAIL.n542 VTAIL.n472 6.59444
R873 VTAIL.n542 VTAIL.n541 6.59444
R874 VTAIL.n450 VTAIL.n380 6.59444
R875 VTAIL.n450 VTAIL.n449 6.59444
R876 VTAIL.n356 VTAIL.n286 6.59444
R877 VTAIL.n356 VTAIL.n355 6.59444
R878 VTAIL.n685 VTAIL.n680 5.81868
R879 VTAIL.n724 VTAIL.n660 5.81868
R880 VTAIL.n732 VTAIL.n731 5.81868
R881 VTAIL.n35 VTAIL.n30 5.81868
R882 VTAIL.n74 VTAIL.n10 5.81868
R883 VTAIL.n82 VTAIL.n81 5.81868
R884 VTAIL.n127 VTAIL.n122 5.81868
R885 VTAIL.n166 VTAIL.n102 5.81868
R886 VTAIL.n174 VTAIL.n173 5.81868
R887 VTAIL.n221 VTAIL.n216 5.81868
R888 VTAIL.n260 VTAIL.n196 5.81868
R889 VTAIL.n268 VTAIL.n267 5.81868
R890 VTAIL.n640 VTAIL.n639 5.81868
R891 VTAIL.n632 VTAIL.n568 5.81868
R892 VTAIL.n595 VTAIL.n590 5.81868
R893 VTAIL.n546 VTAIL.n545 5.81868
R894 VTAIL.n538 VTAIL.n474 5.81868
R895 VTAIL.n501 VTAIL.n496 5.81868
R896 VTAIL.n454 VTAIL.n453 5.81868
R897 VTAIL.n446 VTAIL.n382 5.81868
R898 VTAIL.n409 VTAIL.n404 5.81868
R899 VTAIL.n360 VTAIL.n359 5.81868
R900 VTAIL.n352 VTAIL.n288 5.81868
R901 VTAIL.n315 VTAIL.n310 5.81868
R902 VTAIL.n686 VTAIL.n678 5.04292
R903 VTAIL.n723 VTAIL.n662 5.04292
R904 VTAIL.n735 VTAIL.n656 5.04292
R905 VTAIL.n36 VTAIL.n28 5.04292
R906 VTAIL.n73 VTAIL.n12 5.04292
R907 VTAIL.n85 VTAIL.n6 5.04292
R908 VTAIL.n128 VTAIL.n120 5.04292
R909 VTAIL.n165 VTAIL.n104 5.04292
R910 VTAIL.n177 VTAIL.n98 5.04292
R911 VTAIL.n222 VTAIL.n214 5.04292
R912 VTAIL.n259 VTAIL.n198 5.04292
R913 VTAIL.n271 VTAIL.n192 5.04292
R914 VTAIL.n643 VTAIL.n564 5.04292
R915 VTAIL.n631 VTAIL.n570 5.04292
R916 VTAIL.n596 VTAIL.n588 5.04292
R917 VTAIL.n549 VTAIL.n470 5.04292
R918 VTAIL.n537 VTAIL.n476 5.04292
R919 VTAIL.n502 VTAIL.n494 5.04292
R920 VTAIL.n457 VTAIL.n378 5.04292
R921 VTAIL.n445 VTAIL.n384 5.04292
R922 VTAIL.n410 VTAIL.n402 5.04292
R923 VTAIL.n363 VTAIL.n284 5.04292
R924 VTAIL.n351 VTAIL.n290 5.04292
R925 VTAIL.n316 VTAIL.n308 5.04292
R926 VTAIL.n690 VTAIL.n689 4.26717
R927 VTAIL.n720 VTAIL.n719 4.26717
R928 VTAIL.n736 VTAIL.n654 4.26717
R929 VTAIL.n40 VTAIL.n39 4.26717
R930 VTAIL.n70 VTAIL.n69 4.26717
R931 VTAIL.n86 VTAIL.n4 4.26717
R932 VTAIL.n132 VTAIL.n131 4.26717
R933 VTAIL.n162 VTAIL.n161 4.26717
R934 VTAIL.n178 VTAIL.n96 4.26717
R935 VTAIL.n226 VTAIL.n225 4.26717
R936 VTAIL.n256 VTAIL.n255 4.26717
R937 VTAIL.n272 VTAIL.n190 4.26717
R938 VTAIL.n644 VTAIL.n562 4.26717
R939 VTAIL.n628 VTAIL.n627 4.26717
R940 VTAIL.n600 VTAIL.n599 4.26717
R941 VTAIL.n550 VTAIL.n468 4.26717
R942 VTAIL.n534 VTAIL.n533 4.26717
R943 VTAIL.n506 VTAIL.n505 4.26717
R944 VTAIL.n458 VTAIL.n376 4.26717
R945 VTAIL.n442 VTAIL.n441 4.26717
R946 VTAIL.n414 VTAIL.n413 4.26717
R947 VTAIL.n364 VTAIL.n282 4.26717
R948 VTAIL.n348 VTAIL.n347 4.26717
R949 VTAIL.n320 VTAIL.n319 4.26717
R950 VTAIL.n693 VTAIL.n676 3.49141
R951 VTAIL.n716 VTAIL.n664 3.49141
R952 VTAIL.n740 VTAIL.n739 3.49141
R953 VTAIL.n43 VTAIL.n26 3.49141
R954 VTAIL.n66 VTAIL.n14 3.49141
R955 VTAIL.n90 VTAIL.n89 3.49141
R956 VTAIL.n135 VTAIL.n118 3.49141
R957 VTAIL.n158 VTAIL.n106 3.49141
R958 VTAIL.n182 VTAIL.n181 3.49141
R959 VTAIL.n229 VTAIL.n212 3.49141
R960 VTAIL.n252 VTAIL.n200 3.49141
R961 VTAIL.n276 VTAIL.n275 3.49141
R962 VTAIL.n648 VTAIL.n647 3.49141
R963 VTAIL.n624 VTAIL.n572 3.49141
R964 VTAIL.n603 VTAIL.n586 3.49141
R965 VTAIL.n554 VTAIL.n553 3.49141
R966 VTAIL.n530 VTAIL.n478 3.49141
R967 VTAIL.n509 VTAIL.n492 3.49141
R968 VTAIL.n462 VTAIL.n461 3.49141
R969 VTAIL.n438 VTAIL.n386 3.49141
R970 VTAIL.n417 VTAIL.n400 3.49141
R971 VTAIL.n368 VTAIL.n367 3.49141
R972 VTAIL.n344 VTAIL.n292 3.49141
R973 VTAIL.n323 VTAIL.n306 3.49141
R974 VTAIL.n373 VTAIL.n371 3.06084
R975 VTAIL.n465 VTAIL.n373 3.06084
R976 VTAIL.n559 VTAIL.n557 3.06084
R977 VTAIL.n651 VTAIL.n559 3.06084
R978 VTAIL.n279 VTAIL.n187 3.06084
R979 VTAIL.n187 VTAIL.n185 3.06084
R980 VTAIL.n93 VTAIL.n1 3.06084
R981 VTAIL VTAIL.n743 3.00266
R982 VTAIL.n681 VTAIL.n679 2.84303
R983 VTAIL.n31 VTAIL.n29 2.84303
R984 VTAIL.n123 VTAIL.n121 2.84303
R985 VTAIL.n217 VTAIL.n215 2.84303
R986 VTAIL.n591 VTAIL.n589 2.84303
R987 VTAIL.n497 VTAIL.n495 2.84303
R988 VTAIL.n405 VTAIL.n403 2.84303
R989 VTAIL.n311 VTAIL.n309 2.84303
R990 VTAIL.n694 VTAIL.n674 2.71565
R991 VTAIL.n715 VTAIL.n666 2.71565
R992 VTAIL.n742 VTAIL.n652 2.71565
R993 VTAIL.n44 VTAIL.n24 2.71565
R994 VTAIL.n65 VTAIL.n16 2.71565
R995 VTAIL.n92 VTAIL.n2 2.71565
R996 VTAIL.n136 VTAIL.n116 2.71565
R997 VTAIL.n157 VTAIL.n108 2.71565
R998 VTAIL.n184 VTAIL.n94 2.71565
R999 VTAIL.n230 VTAIL.n210 2.71565
R1000 VTAIL.n251 VTAIL.n202 2.71565
R1001 VTAIL.n278 VTAIL.n188 2.71565
R1002 VTAIL.n650 VTAIL.n560 2.71565
R1003 VTAIL.n623 VTAIL.n574 2.71565
R1004 VTAIL.n604 VTAIL.n584 2.71565
R1005 VTAIL.n556 VTAIL.n466 2.71565
R1006 VTAIL.n529 VTAIL.n480 2.71565
R1007 VTAIL.n510 VTAIL.n490 2.71565
R1008 VTAIL.n464 VTAIL.n374 2.71565
R1009 VTAIL.n437 VTAIL.n388 2.71565
R1010 VTAIL.n418 VTAIL.n398 2.71565
R1011 VTAIL.n370 VTAIL.n280 2.71565
R1012 VTAIL.n343 VTAIL.n294 2.71565
R1013 VTAIL.n324 VTAIL.n304 2.71565
R1014 VTAIL.n699 VTAIL.n697 1.93989
R1015 VTAIL.n712 VTAIL.n711 1.93989
R1016 VTAIL.n49 VTAIL.n47 1.93989
R1017 VTAIL.n62 VTAIL.n61 1.93989
R1018 VTAIL.n141 VTAIL.n139 1.93989
R1019 VTAIL.n154 VTAIL.n153 1.93989
R1020 VTAIL.n235 VTAIL.n233 1.93989
R1021 VTAIL.n248 VTAIL.n247 1.93989
R1022 VTAIL.n620 VTAIL.n619 1.93989
R1023 VTAIL.n608 VTAIL.n607 1.93989
R1024 VTAIL.n526 VTAIL.n525 1.93989
R1025 VTAIL.n514 VTAIL.n513 1.93989
R1026 VTAIL.n434 VTAIL.n433 1.93989
R1027 VTAIL.n422 VTAIL.n421 1.93989
R1028 VTAIL.n340 VTAIL.n339 1.93989
R1029 VTAIL.n328 VTAIL.n327 1.93989
R1030 VTAIL.n0 VTAIL.t7 1.18898
R1031 VTAIL.n0 VTAIL.t11 1.18898
R1032 VTAIL.n186 VTAIL.t4 1.18898
R1033 VTAIL.n186 VTAIL.t15 1.18898
R1034 VTAIL.n558 VTAIL.t2 1.18898
R1035 VTAIL.n558 VTAIL.t0 1.18898
R1036 VTAIL.n372 VTAIL.t10 1.18898
R1037 VTAIL.n372 VTAIL.t13 1.18898
R1038 VTAIL.n698 VTAIL.n672 1.16414
R1039 VTAIL.n708 VTAIL.n668 1.16414
R1040 VTAIL.n48 VTAIL.n22 1.16414
R1041 VTAIL.n58 VTAIL.n18 1.16414
R1042 VTAIL.n140 VTAIL.n114 1.16414
R1043 VTAIL.n150 VTAIL.n110 1.16414
R1044 VTAIL.n234 VTAIL.n208 1.16414
R1045 VTAIL.n244 VTAIL.n204 1.16414
R1046 VTAIL.n616 VTAIL.n576 1.16414
R1047 VTAIL.n611 VTAIL.n581 1.16414
R1048 VTAIL.n522 VTAIL.n482 1.16414
R1049 VTAIL.n517 VTAIL.n487 1.16414
R1050 VTAIL.n430 VTAIL.n390 1.16414
R1051 VTAIL.n425 VTAIL.n395 1.16414
R1052 VTAIL.n336 VTAIL.n296 1.16414
R1053 VTAIL.n331 VTAIL.n301 1.16414
R1054 VTAIL.n557 VTAIL.n465 0.470328
R1055 VTAIL.n185 VTAIL.n93 0.470328
R1056 VTAIL.n704 VTAIL.n703 0.388379
R1057 VTAIL.n707 VTAIL.n670 0.388379
R1058 VTAIL.n54 VTAIL.n53 0.388379
R1059 VTAIL.n57 VTAIL.n20 0.388379
R1060 VTAIL.n146 VTAIL.n145 0.388379
R1061 VTAIL.n149 VTAIL.n112 0.388379
R1062 VTAIL.n240 VTAIL.n239 0.388379
R1063 VTAIL.n243 VTAIL.n206 0.388379
R1064 VTAIL.n615 VTAIL.n578 0.388379
R1065 VTAIL.n612 VTAIL.n580 0.388379
R1066 VTAIL.n521 VTAIL.n484 0.388379
R1067 VTAIL.n518 VTAIL.n486 0.388379
R1068 VTAIL.n429 VTAIL.n392 0.388379
R1069 VTAIL.n426 VTAIL.n394 0.388379
R1070 VTAIL.n335 VTAIL.n298 0.388379
R1071 VTAIL.n332 VTAIL.n300 0.388379
R1072 VTAIL.n687 VTAIL.n679 0.155672
R1073 VTAIL.n688 VTAIL.n687 0.155672
R1074 VTAIL.n688 VTAIL.n675 0.155672
R1075 VTAIL.n695 VTAIL.n675 0.155672
R1076 VTAIL.n696 VTAIL.n695 0.155672
R1077 VTAIL.n696 VTAIL.n671 0.155672
R1078 VTAIL.n705 VTAIL.n671 0.155672
R1079 VTAIL.n706 VTAIL.n705 0.155672
R1080 VTAIL.n706 VTAIL.n667 0.155672
R1081 VTAIL.n713 VTAIL.n667 0.155672
R1082 VTAIL.n714 VTAIL.n713 0.155672
R1083 VTAIL.n714 VTAIL.n663 0.155672
R1084 VTAIL.n721 VTAIL.n663 0.155672
R1085 VTAIL.n722 VTAIL.n721 0.155672
R1086 VTAIL.n722 VTAIL.n659 0.155672
R1087 VTAIL.n729 VTAIL.n659 0.155672
R1088 VTAIL.n730 VTAIL.n729 0.155672
R1089 VTAIL.n730 VTAIL.n655 0.155672
R1090 VTAIL.n737 VTAIL.n655 0.155672
R1091 VTAIL.n738 VTAIL.n737 0.155672
R1092 VTAIL.n37 VTAIL.n29 0.155672
R1093 VTAIL.n38 VTAIL.n37 0.155672
R1094 VTAIL.n38 VTAIL.n25 0.155672
R1095 VTAIL.n45 VTAIL.n25 0.155672
R1096 VTAIL.n46 VTAIL.n45 0.155672
R1097 VTAIL.n46 VTAIL.n21 0.155672
R1098 VTAIL.n55 VTAIL.n21 0.155672
R1099 VTAIL.n56 VTAIL.n55 0.155672
R1100 VTAIL.n56 VTAIL.n17 0.155672
R1101 VTAIL.n63 VTAIL.n17 0.155672
R1102 VTAIL.n64 VTAIL.n63 0.155672
R1103 VTAIL.n64 VTAIL.n13 0.155672
R1104 VTAIL.n71 VTAIL.n13 0.155672
R1105 VTAIL.n72 VTAIL.n71 0.155672
R1106 VTAIL.n72 VTAIL.n9 0.155672
R1107 VTAIL.n79 VTAIL.n9 0.155672
R1108 VTAIL.n80 VTAIL.n79 0.155672
R1109 VTAIL.n80 VTAIL.n5 0.155672
R1110 VTAIL.n87 VTAIL.n5 0.155672
R1111 VTAIL.n88 VTAIL.n87 0.155672
R1112 VTAIL.n129 VTAIL.n121 0.155672
R1113 VTAIL.n130 VTAIL.n129 0.155672
R1114 VTAIL.n130 VTAIL.n117 0.155672
R1115 VTAIL.n137 VTAIL.n117 0.155672
R1116 VTAIL.n138 VTAIL.n137 0.155672
R1117 VTAIL.n138 VTAIL.n113 0.155672
R1118 VTAIL.n147 VTAIL.n113 0.155672
R1119 VTAIL.n148 VTAIL.n147 0.155672
R1120 VTAIL.n148 VTAIL.n109 0.155672
R1121 VTAIL.n155 VTAIL.n109 0.155672
R1122 VTAIL.n156 VTAIL.n155 0.155672
R1123 VTAIL.n156 VTAIL.n105 0.155672
R1124 VTAIL.n163 VTAIL.n105 0.155672
R1125 VTAIL.n164 VTAIL.n163 0.155672
R1126 VTAIL.n164 VTAIL.n101 0.155672
R1127 VTAIL.n171 VTAIL.n101 0.155672
R1128 VTAIL.n172 VTAIL.n171 0.155672
R1129 VTAIL.n172 VTAIL.n97 0.155672
R1130 VTAIL.n179 VTAIL.n97 0.155672
R1131 VTAIL.n180 VTAIL.n179 0.155672
R1132 VTAIL.n223 VTAIL.n215 0.155672
R1133 VTAIL.n224 VTAIL.n223 0.155672
R1134 VTAIL.n224 VTAIL.n211 0.155672
R1135 VTAIL.n231 VTAIL.n211 0.155672
R1136 VTAIL.n232 VTAIL.n231 0.155672
R1137 VTAIL.n232 VTAIL.n207 0.155672
R1138 VTAIL.n241 VTAIL.n207 0.155672
R1139 VTAIL.n242 VTAIL.n241 0.155672
R1140 VTAIL.n242 VTAIL.n203 0.155672
R1141 VTAIL.n249 VTAIL.n203 0.155672
R1142 VTAIL.n250 VTAIL.n249 0.155672
R1143 VTAIL.n250 VTAIL.n199 0.155672
R1144 VTAIL.n257 VTAIL.n199 0.155672
R1145 VTAIL.n258 VTAIL.n257 0.155672
R1146 VTAIL.n258 VTAIL.n195 0.155672
R1147 VTAIL.n265 VTAIL.n195 0.155672
R1148 VTAIL.n266 VTAIL.n265 0.155672
R1149 VTAIL.n266 VTAIL.n191 0.155672
R1150 VTAIL.n273 VTAIL.n191 0.155672
R1151 VTAIL.n274 VTAIL.n273 0.155672
R1152 VTAIL.n646 VTAIL.n645 0.155672
R1153 VTAIL.n645 VTAIL.n563 0.155672
R1154 VTAIL.n638 VTAIL.n563 0.155672
R1155 VTAIL.n638 VTAIL.n637 0.155672
R1156 VTAIL.n637 VTAIL.n567 0.155672
R1157 VTAIL.n630 VTAIL.n567 0.155672
R1158 VTAIL.n630 VTAIL.n629 0.155672
R1159 VTAIL.n629 VTAIL.n571 0.155672
R1160 VTAIL.n622 VTAIL.n571 0.155672
R1161 VTAIL.n622 VTAIL.n621 0.155672
R1162 VTAIL.n621 VTAIL.n575 0.155672
R1163 VTAIL.n614 VTAIL.n575 0.155672
R1164 VTAIL.n614 VTAIL.n613 0.155672
R1165 VTAIL.n613 VTAIL.n579 0.155672
R1166 VTAIL.n606 VTAIL.n579 0.155672
R1167 VTAIL.n606 VTAIL.n605 0.155672
R1168 VTAIL.n605 VTAIL.n585 0.155672
R1169 VTAIL.n598 VTAIL.n585 0.155672
R1170 VTAIL.n598 VTAIL.n597 0.155672
R1171 VTAIL.n597 VTAIL.n589 0.155672
R1172 VTAIL.n552 VTAIL.n551 0.155672
R1173 VTAIL.n551 VTAIL.n469 0.155672
R1174 VTAIL.n544 VTAIL.n469 0.155672
R1175 VTAIL.n544 VTAIL.n543 0.155672
R1176 VTAIL.n543 VTAIL.n473 0.155672
R1177 VTAIL.n536 VTAIL.n473 0.155672
R1178 VTAIL.n536 VTAIL.n535 0.155672
R1179 VTAIL.n535 VTAIL.n477 0.155672
R1180 VTAIL.n528 VTAIL.n477 0.155672
R1181 VTAIL.n528 VTAIL.n527 0.155672
R1182 VTAIL.n527 VTAIL.n481 0.155672
R1183 VTAIL.n520 VTAIL.n481 0.155672
R1184 VTAIL.n520 VTAIL.n519 0.155672
R1185 VTAIL.n519 VTAIL.n485 0.155672
R1186 VTAIL.n512 VTAIL.n485 0.155672
R1187 VTAIL.n512 VTAIL.n511 0.155672
R1188 VTAIL.n511 VTAIL.n491 0.155672
R1189 VTAIL.n504 VTAIL.n491 0.155672
R1190 VTAIL.n504 VTAIL.n503 0.155672
R1191 VTAIL.n503 VTAIL.n495 0.155672
R1192 VTAIL.n460 VTAIL.n459 0.155672
R1193 VTAIL.n459 VTAIL.n377 0.155672
R1194 VTAIL.n452 VTAIL.n377 0.155672
R1195 VTAIL.n452 VTAIL.n451 0.155672
R1196 VTAIL.n451 VTAIL.n381 0.155672
R1197 VTAIL.n444 VTAIL.n381 0.155672
R1198 VTAIL.n444 VTAIL.n443 0.155672
R1199 VTAIL.n443 VTAIL.n385 0.155672
R1200 VTAIL.n436 VTAIL.n385 0.155672
R1201 VTAIL.n436 VTAIL.n435 0.155672
R1202 VTAIL.n435 VTAIL.n389 0.155672
R1203 VTAIL.n428 VTAIL.n389 0.155672
R1204 VTAIL.n428 VTAIL.n427 0.155672
R1205 VTAIL.n427 VTAIL.n393 0.155672
R1206 VTAIL.n420 VTAIL.n393 0.155672
R1207 VTAIL.n420 VTAIL.n419 0.155672
R1208 VTAIL.n419 VTAIL.n399 0.155672
R1209 VTAIL.n412 VTAIL.n399 0.155672
R1210 VTAIL.n412 VTAIL.n411 0.155672
R1211 VTAIL.n411 VTAIL.n403 0.155672
R1212 VTAIL.n366 VTAIL.n365 0.155672
R1213 VTAIL.n365 VTAIL.n283 0.155672
R1214 VTAIL.n358 VTAIL.n283 0.155672
R1215 VTAIL.n358 VTAIL.n357 0.155672
R1216 VTAIL.n357 VTAIL.n287 0.155672
R1217 VTAIL.n350 VTAIL.n287 0.155672
R1218 VTAIL.n350 VTAIL.n349 0.155672
R1219 VTAIL.n349 VTAIL.n291 0.155672
R1220 VTAIL.n342 VTAIL.n291 0.155672
R1221 VTAIL.n342 VTAIL.n341 0.155672
R1222 VTAIL.n341 VTAIL.n295 0.155672
R1223 VTAIL.n334 VTAIL.n295 0.155672
R1224 VTAIL.n334 VTAIL.n333 0.155672
R1225 VTAIL.n333 VTAIL.n299 0.155672
R1226 VTAIL.n326 VTAIL.n299 0.155672
R1227 VTAIL.n326 VTAIL.n325 0.155672
R1228 VTAIL.n325 VTAIL.n305 0.155672
R1229 VTAIL.n318 VTAIL.n305 0.155672
R1230 VTAIL.n318 VTAIL.n317 0.155672
R1231 VTAIL.n317 VTAIL.n309 0.155672
R1232 VTAIL VTAIL.n1 0.0586897
R1233 VDD2.n2 VDD2.n1 65.7287
R1234 VDD2.n2 VDD2.n0 65.7287
R1235 VDD2 VDD2.n5 65.7248
R1236 VDD2.n4 VDD2.n3 64.254
R1237 VDD2.n4 VDD2.n2 51.8489
R1238 VDD2 VDD2.n4 1.58886
R1239 VDD2.n5 VDD2.t5 1.18898
R1240 VDD2.n5 VDD2.t2 1.18898
R1241 VDD2.n3 VDD2.t3 1.18898
R1242 VDD2.n3 VDD2.t7 1.18898
R1243 VDD2.n1 VDD2.t1 1.18898
R1244 VDD2.n1 VDD2.t0 1.18898
R1245 VDD2.n0 VDD2.t6 1.18898
R1246 VDD2.n0 VDD2.t4 1.18898
R1247 B.n1095 B.n1094 585
R1248 B.n412 B.n171 585
R1249 B.n411 B.n410 585
R1250 B.n409 B.n408 585
R1251 B.n407 B.n406 585
R1252 B.n405 B.n404 585
R1253 B.n403 B.n402 585
R1254 B.n401 B.n400 585
R1255 B.n399 B.n398 585
R1256 B.n397 B.n396 585
R1257 B.n395 B.n394 585
R1258 B.n393 B.n392 585
R1259 B.n391 B.n390 585
R1260 B.n389 B.n388 585
R1261 B.n387 B.n386 585
R1262 B.n385 B.n384 585
R1263 B.n383 B.n382 585
R1264 B.n381 B.n380 585
R1265 B.n379 B.n378 585
R1266 B.n377 B.n376 585
R1267 B.n375 B.n374 585
R1268 B.n373 B.n372 585
R1269 B.n371 B.n370 585
R1270 B.n369 B.n368 585
R1271 B.n367 B.n366 585
R1272 B.n365 B.n364 585
R1273 B.n363 B.n362 585
R1274 B.n361 B.n360 585
R1275 B.n359 B.n358 585
R1276 B.n357 B.n356 585
R1277 B.n355 B.n354 585
R1278 B.n353 B.n352 585
R1279 B.n351 B.n350 585
R1280 B.n349 B.n348 585
R1281 B.n347 B.n346 585
R1282 B.n345 B.n344 585
R1283 B.n343 B.n342 585
R1284 B.n341 B.n340 585
R1285 B.n339 B.n338 585
R1286 B.n337 B.n336 585
R1287 B.n335 B.n334 585
R1288 B.n333 B.n332 585
R1289 B.n331 B.n330 585
R1290 B.n329 B.n328 585
R1291 B.n327 B.n326 585
R1292 B.n325 B.n324 585
R1293 B.n323 B.n322 585
R1294 B.n321 B.n320 585
R1295 B.n319 B.n318 585
R1296 B.n317 B.n316 585
R1297 B.n315 B.n314 585
R1298 B.n313 B.n312 585
R1299 B.n311 B.n310 585
R1300 B.n309 B.n308 585
R1301 B.n307 B.n306 585
R1302 B.n304 B.n303 585
R1303 B.n302 B.n301 585
R1304 B.n300 B.n299 585
R1305 B.n298 B.n297 585
R1306 B.n296 B.n295 585
R1307 B.n294 B.n293 585
R1308 B.n292 B.n291 585
R1309 B.n290 B.n289 585
R1310 B.n288 B.n287 585
R1311 B.n286 B.n285 585
R1312 B.n283 B.n282 585
R1313 B.n281 B.n280 585
R1314 B.n279 B.n278 585
R1315 B.n277 B.n276 585
R1316 B.n275 B.n274 585
R1317 B.n273 B.n272 585
R1318 B.n271 B.n270 585
R1319 B.n269 B.n268 585
R1320 B.n267 B.n266 585
R1321 B.n265 B.n264 585
R1322 B.n263 B.n262 585
R1323 B.n261 B.n260 585
R1324 B.n259 B.n258 585
R1325 B.n257 B.n256 585
R1326 B.n255 B.n254 585
R1327 B.n253 B.n252 585
R1328 B.n251 B.n250 585
R1329 B.n249 B.n248 585
R1330 B.n247 B.n246 585
R1331 B.n245 B.n244 585
R1332 B.n243 B.n242 585
R1333 B.n241 B.n240 585
R1334 B.n239 B.n238 585
R1335 B.n237 B.n236 585
R1336 B.n235 B.n234 585
R1337 B.n233 B.n232 585
R1338 B.n231 B.n230 585
R1339 B.n229 B.n228 585
R1340 B.n227 B.n226 585
R1341 B.n225 B.n224 585
R1342 B.n223 B.n222 585
R1343 B.n221 B.n220 585
R1344 B.n219 B.n218 585
R1345 B.n217 B.n216 585
R1346 B.n215 B.n214 585
R1347 B.n213 B.n212 585
R1348 B.n211 B.n210 585
R1349 B.n209 B.n208 585
R1350 B.n207 B.n206 585
R1351 B.n205 B.n204 585
R1352 B.n203 B.n202 585
R1353 B.n201 B.n200 585
R1354 B.n199 B.n198 585
R1355 B.n197 B.n196 585
R1356 B.n195 B.n194 585
R1357 B.n193 B.n192 585
R1358 B.n191 B.n190 585
R1359 B.n189 B.n188 585
R1360 B.n187 B.n186 585
R1361 B.n185 B.n184 585
R1362 B.n183 B.n182 585
R1363 B.n181 B.n180 585
R1364 B.n179 B.n178 585
R1365 B.n177 B.n176 585
R1366 B.n110 B.n109 585
R1367 B.n1093 B.n111 585
R1368 B.n1098 B.n111 585
R1369 B.n1092 B.n1091 585
R1370 B.n1091 B.n107 585
R1371 B.n1090 B.n106 585
R1372 B.n1104 B.n106 585
R1373 B.n1089 B.n105 585
R1374 B.n1105 B.n105 585
R1375 B.n1088 B.n104 585
R1376 B.n1106 B.n104 585
R1377 B.n1087 B.n1086 585
R1378 B.n1086 B.n100 585
R1379 B.n1085 B.n99 585
R1380 B.n1112 B.n99 585
R1381 B.n1084 B.n98 585
R1382 B.n1113 B.n98 585
R1383 B.n1083 B.n97 585
R1384 B.n1114 B.n97 585
R1385 B.n1082 B.n1081 585
R1386 B.n1081 B.n93 585
R1387 B.n1080 B.n92 585
R1388 B.n1120 B.n92 585
R1389 B.n1079 B.n91 585
R1390 B.n1121 B.n91 585
R1391 B.n1078 B.n90 585
R1392 B.n1122 B.n90 585
R1393 B.n1077 B.n1076 585
R1394 B.n1076 B.n86 585
R1395 B.n1075 B.n85 585
R1396 B.n1128 B.n85 585
R1397 B.n1074 B.n84 585
R1398 B.n1129 B.n84 585
R1399 B.n1073 B.n83 585
R1400 B.n1130 B.n83 585
R1401 B.n1072 B.n1071 585
R1402 B.n1071 B.n79 585
R1403 B.n1070 B.n78 585
R1404 B.n1136 B.n78 585
R1405 B.n1069 B.n77 585
R1406 B.n1137 B.n77 585
R1407 B.n1068 B.n76 585
R1408 B.n1138 B.n76 585
R1409 B.n1067 B.n1066 585
R1410 B.n1066 B.n72 585
R1411 B.n1065 B.n71 585
R1412 B.n1144 B.n71 585
R1413 B.n1064 B.n70 585
R1414 B.n1145 B.n70 585
R1415 B.n1063 B.n69 585
R1416 B.n1146 B.n69 585
R1417 B.n1062 B.n1061 585
R1418 B.n1061 B.n65 585
R1419 B.n1060 B.n64 585
R1420 B.n1152 B.n64 585
R1421 B.n1059 B.n63 585
R1422 B.n1153 B.n63 585
R1423 B.n1058 B.n62 585
R1424 B.n1154 B.n62 585
R1425 B.n1057 B.n1056 585
R1426 B.n1056 B.n58 585
R1427 B.n1055 B.n57 585
R1428 B.n1160 B.n57 585
R1429 B.n1054 B.n56 585
R1430 B.n1161 B.n56 585
R1431 B.n1053 B.n55 585
R1432 B.n1162 B.n55 585
R1433 B.n1052 B.n1051 585
R1434 B.n1051 B.n51 585
R1435 B.n1050 B.n50 585
R1436 B.n1168 B.n50 585
R1437 B.n1049 B.n49 585
R1438 B.n1169 B.n49 585
R1439 B.n1048 B.n48 585
R1440 B.n1170 B.n48 585
R1441 B.n1047 B.n1046 585
R1442 B.n1046 B.n44 585
R1443 B.n1045 B.n43 585
R1444 B.n1176 B.n43 585
R1445 B.n1044 B.n42 585
R1446 B.n1177 B.n42 585
R1447 B.n1043 B.n41 585
R1448 B.n1178 B.n41 585
R1449 B.n1042 B.n1041 585
R1450 B.n1041 B.n37 585
R1451 B.n1040 B.n36 585
R1452 B.n1184 B.n36 585
R1453 B.n1039 B.n35 585
R1454 B.n1185 B.n35 585
R1455 B.n1038 B.n34 585
R1456 B.n1186 B.n34 585
R1457 B.n1037 B.n1036 585
R1458 B.n1036 B.n30 585
R1459 B.n1035 B.n29 585
R1460 B.n1192 B.n29 585
R1461 B.n1034 B.n28 585
R1462 B.n1193 B.n28 585
R1463 B.n1033 B.n27 585
R1464 B.n1194 B.n27 585
R1465 B.n1032 B.n1031 585
R1466 B.n1031 B.n23 585
R1467 B.n1030 B.n22 585
R1468 B.n1200 B.n22 585
R1469 B.n1029 B.n21 585
R1470 B.n1201 B.n21 585
R1471 B.n1028 B.n20 585
R1472 B.n1202 B.n20 585
R1473 B.n1027 B.n1026 585
R1474 B.n1026 B.n19 585
R1475 B.n1025 B.n15 585
R1476 B.n1208 B.n15 585
R1477 B.n1024 B.n14 585
R1478 B.n1209 B.n14 585
R1479 B.n1023 B.n13 585
R1480 B.n1210 B.n13 585
R1481 B.n1022 B.n1021 585
R1482 B.n1021 B.n12 585
R1483 B.n1020 B.n1019 585
R1484 B.n1020 B.n8 585
R1485 B.n1018 B.n7 585
R1486 B.n1217 B.n7 585
R1487 B.n1017 B.n6 585
R1488 B.n1218 B.n6 585
R1489 B.n1016 B.n5 585
R1490 B.n1219 B.n5 585
R1491 B.n1015 B.n1014 585
R1492 B.n1014 B.n4 585
R1493 B.n1013 B.n413 585
R1494 B.n1013 B.n1012 585
R1495 B.n1003 B.n414 585
R1496 B.n415 B.n414 585
R1497 B.n1005 B.n1004 585
R1498 B.n1006 B.n1005 585
R1499 B.n1002 B.n420 585
R1500 B.n420 B.n419 585
R1501 B.n1001 B.n1000 585
R1502 B.n1000 B.n999 585
R1503 B.n422 B.n421 585
R1504 B.n992 B.n422 585
R1505 B.n991 B.n990 585
R1506 B.n993 B.n991 585
R1507 B.n989 B.n427 585
R1508 B.n427 B.n426 585
R1509 B.n988 B.n987 585
R1510 B.n987 B.n986 585
R1511 B.n429 B.n428 585
R1512 B.n430 B.n429 585
R1513 B.n979 B.n978 585
R1514 B.n980 B.n979 585
R1515 B.n977 B.n435 585
R1516 B.n435 B.n434 585
R1517 B.n976 B.n975 585
R1518 B.n975 B.n974 585
R1519 B.n437 B.n436 585
R1520 B.n438 B.n437 585
R1521 B.n967 B.n966 585
R1522 B.n968 B.n967 585
R1523 B.n965 B.n442 585
R1524 B.n446 B.n442 585
R1525 B.n964 B.n963 585
R1526 B.n963 B.n962 585
R1527 B.n444 B.n443 585
R1528 B.n445 B.n444 585
R1529 B.n955 B.n954 585
R1530 B.n956 B.n955 585
R1531 B.n953 B.n451 585
R1532 B.n451 B.n450 585
R1533 B.n952 B.n951 585
R1534 B.n951 B.n950 585
R1535 B.n453 B.n452 585
R1536 B.n454 B.n453 585
R1537 B.n943 B.n942 585
R1538 B.n944 B.n943 585
R1539 B.n941 B.n459 585
R1540 B.n459 B.n458 585
R1541 B.n940 B.n939 585
R1542 B.n939 B.n938 585
R1543 B.n461 B.n460 585
R1544 B.n462 B.n461 585
R1545 B.n931 B.n930 585
R1546 B.n932 B.n931 585
R1547 B.n929 B.n467 585
R1548 B.n467 B.n466 585
R1549 B.n928 B.n927 585
R1550 B.n927 B.n926 585
R1551 B.n469 B.n468 585
R1552 B.n470 B.n469 585
R1553 B.n919 B.n918 585
R1554 B.n920 B.n919 585
R1555 B.n917 B.n475 585
R1556 B.n475 B.n474 585
R1557 B.n916 B.n915 585
R1558 B.n915 B.n914 585
R1559 B.n477 B.n476 585
R1560 B.n478 B.n477 585
R1561 B.n907 B.n906 585
R1562 B.n908 B.n907 585
R1563 B.n905 B.n483 585
R1564 B.n483 B.n482 585
R1565 B.n904 B.n903 585
R1566 B.n903 B.n902 585
R1567 B.n485 B.n484 585
R1568 B.n486 B.n485 585
R1569 B.n895 B.n894 585
R1570 B.n896 B.n895 585
R1571 B.n893 B.n491 585
R1572 B.n491 B.n490 585
R1573 B.n892 B.n891 585
R1574 B.n891 B.n890 585
R1575 B.n493 B.n492 585
R1576 B.n494 B.n493 585
R1577 B.n883 B.n882 585
R1578 B.n884 B.n883 585
R1579 B.n881 B.n499 585
R1580 B.n499 B.n498 585
R1581 B.n880 B.n879 585
R1582 B.n879 B.n878 585
R1583 B.n501 B.n500 585
R1584 B.n502 B.n501 585
R1585 B.n871 B.n870 585
R1586 B.n872 B.n871 585
R1587 B.n869 B.n507 585
R1588 B.n507 B.n506 585
R1589 B.n868 B.n867 585
R1590 B.n867 B.n866 585
R1591 B.n509 B.n508 585
R1592 B.n510 B.n509 585
R1593 B.n859 B.n858 585
R1594 B.n860 B.n859 585
R1595 B.n857 B.n515 585
R1596 B.n515 B.n514 585
R1597 B.n856 B.n855 585
R1598 B.n855 B.n854 585
R1599 B.n517 B.n516 585
R1600 B.n518 B.n517 585
R1601 B.n847 B.n846 585
R1602 B.n848 B.n847 585
R1603 B.n845 B.n523 585
R1604 B.n523 B.n522 585
R1605 B.n844 B.n843 585
R1606 B.n843 B.n842 585
R1607 B.n525 B.n524 585
R1608 B.n526 B.n525 585
R1609 B.n835 B.n834 585
R1610 B.n836 B.n835 585
R1611 B.n529 B.n528 585
R1612 B.n598 B.n597 585
R1613 B.n599 B.n595 585
R1614 B.n595 B.n530 585
R1615 B.n601 B.n600 585
R1616 B.n603 B.n594 585
R1617 B.n606 B.n605 585
R1618 B.n607 B.n593 585
R1619 B.n609 B.n608 585
R1620 B.n611 B.n592 585
R1621 B.n614 B.n613 585
R1622 B.n615 B.n591 585
R1623 B.n617 B.n616 585
R1624 B.n619 B.n590 585
R1625 B.n622 B.n621 585
R1626 B.n623 B.n589 585
R1627 B.n625 B.n624 585
R1628 B.n627 B.n588 585
R1629 B.n630 B.n629 585
R1630 B.n631 B.n587 585
R1631 B.n633 B.n632 585
R1632 B.n635 B.n586 585
R1633 B.n638 B.n637 585
R1634 B.n639 B.n585 585
R1635 B.n641 B.n640 585
R1636 B.n643 B.n584 585
R1637 B.n646 B.n645 585
R1638 B.n647 B.n583 585
R1639 B.n649 B.n648 585
R1640 B.n651 B.n582 585
R1641 B.n654 B.n653 585
R1642 B.n655 B.n581 585
R1643 B.n657 B.n656 585
R1644 B.n659 B.n580 585
R1645 B.n662 B.n661 585
R1646 B.n663 B.n579 585
R1647 B.n665 B.n664 585
R1648 B.n667 B.n578 585
R1649 B.n670 B.n669 585
R1650 B.n671 B.n577 585
R1651 B.n673 B.n672 585
R1652 B.n675 B.n576 585
R1653 B.n678 B.n677 585
R1654 B.n679 B.n575 585
R1655 B.n681 B.n680 585
R1656 B.n683 B.n574 585
R1657 B.n686 B.n685 585
R1658 B.n687 B.n573 585
R1659 B.n689 B.n688 585
R1660 B.n691 B.n572 585
R1661 B.n694 B.n693 585
R1662 B.n695 B.n571 585
R1663 B.n697 B.n696 585
R1664 B.n699 B.n570 585
R1665 B.n702 B.n701 585
R1666 B.n703 B.n567 585
R1667 B.n706 B.n705 585
R1668 B.n708 B.n566 585
R1669 B.n711 B.n710 585
R1670 B.n712 B.n565 585
R1671 B.n714 B.n713 585
R1672 B.n716 B.n564 585
R1673 B.n719 B.n718 585
R1674 B.n720 B.n563 585
R1675 B.n722 B.n721 585
R1676 B.n724 B.n562 585
R1677 B.n727 B.n726 585
R1678 B.n728 B.n558 585
R1679 B.n730 B.n729 585
R1680 B.n732 B.n557 585
R1681 B.n735 B.n734 585
R1682 B.n736 B.n556 585
R1683 B.n738 B.n737 585
R1684 B.n740 B.n555 585
R1685 B.n743 B.n742 585
R1686 B.n744 B.n554 585
R1687 B.n746 B.n745 585
R1688 B.n748 B.n553 585
R1689 B.n751 B.n750 585
R1690 B.n752 B.n552 585
R1691 B.n754 B.n753 585
R1692 B.n756 B.n551 585
R1693 B.n759 B.n758 585
R1694 B.n760 B.n550 585
R1695 B.n762 B.n761 585
R1696 B.n764 B.n549 585
R1697 B.n767 B.n766 585
R1698 B.n768 B.n548 585
R1699 B.n770 B.n769 585
R1700 B.n772 B.n547 585
R1701 B.n775 B.n774 585
R1702 B.n776 B.n546 585
R1703 B.n778 B.n777 585
R1704 B.n780 B.n545 585
R1705 B.n783 B.n782 585
R1706 B.n784 B.n544 585
R1707 B.n786 B.n785 585
R1708 B.n788 B.n543 585
R1709 B.n791 B.n790 585
R1710 B.n792 B.n542 585
R1711 B.n794 B.n793 585
R1712 B.n796 B.n541 585
R1713 B.n799 B.n798 585
R1714 B.n800 B.n540 585
R1715 B.n802 B.n801 585
R1716 B.n804 B.n539 585
R1717 B.n807 B.n806 585
R1718 B.n808 B.n538 585
R1719 B.n810 B.n809 585
R1720 B.n812 B.n537 585
R1721 B.n815 B.n814 585
R1722 B.n816 B.n536 585
R1723 B.n818 B.n817 585
R1724 B.n820 B.n535 585
R1725 B.n823 B.n822 585
R1726 B.n824 B.n534 585
R1727 B.n826 B.n825 585
R1728 B.n828 B.n533 585
R1729 B.n829 B.n532 585
R1730 B.n832 B.n831 585
R1731 B.n833 B.n531 585
R1732 B.n531 B.n530 585
R1733 B.n838 B.n837 585
R1734 B.n837 B.n836 585
R1735 B.n839 B.n527 585
R1736 B.n527 B.n526 585
R1737 B.n841 B.n840 585
R1738 B.n842 B.n841 585
R1739 B.n521 B.n520 585
R1740 B.n522 B.n521 585
R1741 B.n850 B.n849 585
R1742 B.n849 B.n848 585
R1743 B.n851 B.n519 585
R1744 B.n519 B.n518 585
R1745 B.n853 B.n852 585
R1746 B.n854 B.n853 585
R1747 B.n513 B.n512 585
R1748 B.n514 B.n513 585
R1749 B.n862 B.n861 585
R1750 B.n861 B.n860 585
R1751 B.n863 B.n511 585
R1752 B.n511 B.n510 585
R1753 B.n865 B.n864 585
R1754 B.n866 B.n865 585
R1755 B.n505 B.n504 585
R1756 B.n506 B.n505 585
R1757 B.n874 B.n873 585
R1758 B.n873 B.n872 585
R1759 B.n875 B.n503 585
R1760 B.n503 B.n502 585
R1761 B.n877 B.n876 585
R1762 B.n878 B.n877 585
R1763 B.n497 B.n496 585
R1764 B.n498 B.n497 585
R1765 B.n886 B.n885 585
R1766 B.n885 B.n884 585
R1767 B.n887 B.n495 585
R1768 B.n495 B.n494 585
R1769 B.n889 B.n888 585
R1770 B.n890 B.n889 585
R1771 B.n489 B.n488 585
R1772 B.n490 B.n489 585
R1773 B.n898 B.n897 585
R1774 B.n897 B.n896 585
R1775 B.n899 B.n487 585
R1776 B.n487 B.n486 585
R1777 B.n901 B.n900 585
R1778 B.n902 B.n901 585
R1779 B.n481 B.n480 585
R1780 B.n482 B.n481 585
R1781 B.n910 B.n909 585
R1782 B.n909 B.n908 585
R1783 B.n911 B.n479 585
R1784 B.n479 B.n478 585
R1785 B.n913 B.n912 585
R1786 B.n914 B.n913 585
R1787 B.n473 B.n472 585
R1788 B.n474 B.n473 585
R1789 B.n922 B.n921 585
R1790 B.n921 B.n920 585
R1791 B.n923 B.n471 585
R1792 B.n471 B.n470 585
R1793 B.n925 B.n924 585
R1794 B.n926 B.n925 585
R1795 B.n465 B.n464 585
R1796 B.n466 B.n465 585
R1797 B.n934 B.n933 585
R1798 B.n933 B.n932 585
R1799 B.n935 B.n463 585
R1800 B.n463 B.n462 585
R1801 B.n937 B.n936 585
R1802 B.n938 B.n937 585
R1803 B.n457 B.n456 585
R1804 B.n458 B.n457 585
R1805 B.n946 B.n945 585
R1806 B.n945 B.n944 585
R1807 B.n947 B.n455 585
R1808 B.n455 B.n454 585
R1809 B.n949 B.n948 585
R1810 B.n950 B.n949 585
R1811 B.n449 B.n448 585
R1812 B.n450 B.n449 585
R1813 B.n958 B.n957 585
R1814 B.n957 B.n956 585
R1815 B.n959 B.n447 585
R1816 B.n447 B.n445 585
R1817 B.n961 B.n960 585
R1818 B.n962 B.n961 585
R1819 B.n441 B.n440 585
R1820 B.n446 B.n441 585
R1821 B.n970 B.n969 585
R1822 B.n969 B.n968 585
R1823 B.n971 B.n439 585
R1824 B.n439 B.n438 585
R1825 B.n973 B.n972 585
R1826 B.n974 B.n973 585
R1827 B.n433 B.n432 585
R1828 B.n434 B.n433 585
R1829 B.n982 B.n981 585
R1830 B.n981 B.n980 585
R1831 B.n983 B.n431 585
R1832 B.n431 B.n430 585
R1833 B.n985 B.n984 585
R1834 B.n986 B.n985 585
R1835 B.n425 B.n424 585
R1836 B.n426 B.n425 585
R1837 B.n995 B.n994 585
R1838 B.n994 B.n993 585
R1839 B.n996 B.n423 585
R1840 B.n992 B.n423 585
R1841 B.n998 B.n997 585
R1842 B.n999 B.n998 585
R1843 B.n418 B.n417 585
R1844 B.n419 B.n418 585
R1845 B.n1008 B.n1007 585
R1846 B.n1007 B.n1006 585
R1847 B.n1009 B.n416 585
R1848 B.n416 B.n415 585
R1849 B.n1011 B.n1010 585
R1850 B.n1012 B.n1011 585
R1851 B.n3 B.n0 585
R1852 B.n4 B.n3 585
R1853 B.n1216 B.n1 585
R1854 B.n1217 B.n1216 585
R1855 B.n1215 B.n1214 585
R1856 B.n1215 B.n8 585
R1857 B.n1213 B.n9 585
R1858 B.n12 B.n9 585
R1859 B.n1212 B.n1211 585
R1860 B.n1211 B.n1210 585
R1861 B.n11 B.n10 585
R1862 B.n1209 B.n11 585
R1863 B.n1207 B.n1206 585
R1864 B.n1208 B.n1207 585
R1865 B.n1205 B.n16 585
R1866 B.n19 B.n16 585
R1867 B.n1204 B.n1203 585
R1868 B.n1203 B.n1202 585
R1869 B.n18 B.n17 585
R1870 B.n1201 B.n18 585
R1871 B.n1199 B.n1198 585
R1872 B.n1200 B.n1199 585
R1873 B.n1197 B.n24 585
R1874 B.n24 B.n23 585
R1875 B.n1196 B.n1195 585
R1876 B.n1195 B.n1194 585
R1877 B.n26 B.n25 585
R1878 B.n1193 B.n26 585
R1879 B.n1191 B.n1190 585
R1880 B.n1192 B.n1191 585
R1881 B.n1189 B.n31 585
R1882 B.n31 B.n30 585
R1883 B.n1188 B.n1187 585
R1884 B.n1187 B.n1186 585
R1885 B.n33 B.n32 585
R1886 B.n1185 B.n33 585
R1887 B.n1183 B.n1182 585
R1888 B.n1184 B.n1183 585
R1889 B.n1181 B.n38 585
R1890 B.n38 B.n37 585
R1891 B.n1180 B.n1179 585
R1892 B.n1179 B.n1178 585
R1893 B.n40 B.n39 585
R1894 B.n1177 B.n40 585
R1895 B.n1175 B.n1174 585
R1896 B.n1176 B.n1175 585
R1897 B.n1173 B.n45 585
R1898 B.n45 B.n44 585
R1899 B.n1172 B.n1171 585
R1900 B.n1171 B.n1170 585
R1901 B.n47 B.n46 585
R1902 B.n1169 B.n47 585
R1903 B.n1167 B.n1166 585
R1904 B.n1168 B.n1167 585
R1905 B.n1165 B.n52 585
R1906 B.n52 B.n51 585
R1907 B.n1164 B.n1163 585
R1908 B.n1163 B.n1162 585
R1909 B.n54 B.n53 585
R1910 B.n1161 B.n54 585
R1911 B.n1159 B.n1158 585
R1912 B.n1160 B.n1159 585
R1913 B.n1157 B.n59 585
R1914 B.n59 B.n58 585
R1915 B.n1156 B.n1155 585
R1916 B.n1155 B.n1154 585
R1917 B.n61 B.n60 585
R1918 B.n1153 B.n61 585
R1919 B.n1151 B.n1150 585
R1920 B.n1152 B.n1151 585
R1921 B.n1149 B.n66 585
R1922 B.n66 B.n65 585
R1923 B.n1148 B.n1147 585
R1924 B.n1147 B.n1146 585
R1925 B.n68 B.n67 585
R1926 B.n1145 B.n68 585
R1927 B.n1143 B.n1142 585
R1928 B.n1144 B.n1143 585
R1929 B.n1141 B.n73 585
R1930 B.n73 B.n72 585
R1931 B.n1140 B.n1139 585
R1932 B.n1139 B.n1138 585
R1933 B.n75 B.n74 585
R1934 B.n1137 B.n75 585
R1935 B.n1135 B.n1134 585
R1936 B.n1136 B.n1135 585
R1937 B.n1133 B.n80 585
R1938 B.n80 B.n79 585
R1939 B.n1132 B.n1131 585
R1940 B.n1131 B.n1130 585
R1941 B.n82 B.n81 585
R1942 B.n1129 B.n82 585
R1943 B.n1127 B.n1126 585
R1944 B.n1128 B.n1127 585
R1945 B.n1125 B.n87 585
R1946 B.n87 B.n86 585
R1947 B.n1124 B.n1123 585
R1948 B.n1123 B.n1122 585
R1949 B.n89 B.n88 585
R1950 B.n1121 B.n89 585
R1951 B.n1119 B.n1118 585
R1952 B.n1120 B.n1119 585
R1953 B.n1117 B.n94 585
R1954 B.n94 B.n93 585
R1955 B.n1116 B.n1115 585
R1956 B.n1115 B.n1114 585
R1957 B.n96 B.n95 585
R1958 B.n1113 B.n96 585
R1959 B.n1111 B.n1110 585
R1960 B.n1112 B.n1111 585
R1961 B.n1109 B.n101 585
R1962 B.n101 B.n100 585
R1963 B.n1108 B.n1107 585
R1964 B.n1107 B.n1106 585
R1965 B.n103 B.n102 585
R1966 B.n1105 B.n103 585
R1967 B.n1103 B.n1102 585
R1968 B.n1104 B.n1103 585
R1969 B.n1101 B.n108 585
R1970 B.n108 B.n107 585
R1971 B.n1100 B.n1099 585
R1972 B.n1099 B.n1098 585
R1973 B.n1220 B.n1219 585
R1974 B.n1218 B.n2 585
R1975 B.n1099 B.n110 487.695
R1976 B.n1095 B.n111 487.695
R1977 B.n835 B.n531 487.695
R1978 B.n837 B.n529 487.695
R1979 B.n174 B.t19 430.904
R1980 B.n172 B.t13 430.904
R1981 B.n559 B.t10 430.904
R1982 B.n568 B.t17 430.904
R1983 B.n173 B.t14 362.055
R1984 B.n560 B.t9 362.055
R1985 B.n175 B.t20 362.055
R1986 B.n569 B.t16 362.055
R1987 B.n174 B.t18 333.514
R1988 B.n172 B.t11 333.514
R1989 B.n559 B.t7 333.514
R1990 B.n568 B.t15 333.514
R1991 B.n1097 B.n1096 256.663
R1992 B.n1097 B.n170 256.663
R1993 B.n1097 B.n169 256.663
R1994 B.n1097 B.n168 256.663
R1995 B.n1097 B.n167 256.663
R1996 B.n1097 B.n166 256.663
R1997 B.n1097 B.n165 256.663
R1998 B.n1097 B.n164 256.663
R1999 B.n1097 B.n163 256.663
R2000 B.n1097 B.n162 256.663
R2001 B.n1097 B.n161 256.663
R2002 B.n1097 B.n160 256.663
R2003 B.n1097 B.n159 256.663
R2004 B.n1097 B.n158 256.663
R2005 B.n1097 B.n157 256.663
R2006 B.n1097 B.n156 256.663
R2007 B.n1097 B.n155 256.663
R2008 B.n1097 B.n154 256.663
R2009 B.n1097 B.n153 256.663
R2010 B.n1097 B.n152 256.663
R2011 B.n1097 B.n151 256.663
R2012 B.n1097 B.n150 256.663
R2013 B.n1097 B.n149 256.663
R2014 B.n1097 B.n148 256.663
R2015 B.n1097 B.n147 256.663
R2016 B.n1097 B.n146 256.663
R2017 B.n1097 B.n145 256.663
R2018 B.n1097 B.n144 256.663
R2019 B.n1097 B.n143 256.663
R2020 B.n1097 B.n142 256.663
R2021 B.n1097 B.n141 256.663
R2022 B.n1097 B.n140 256.663
R2023 B.n1097 B.n139 256.663
R2024 B.n1097 B.n138 256.663
R2025 B.n1097 B.n137 256.663
R2026 B.n1097 B.n136 256.663
R2027 B.n1097 B.n135 256.663
R2028 B.n1097 B.n134 256.663
R2029 B.n1097 B.n133 256.663
R2030 B.n1097 B.n132 256.663
R2031 B.n1097 B.n131 256.663
R2032 B.n1097 B.n130 256.663
R2033 B.n1097 B.n129 256.663
R2034 B.n1097 B.n128 256.663
R2035 B.n1097 B.n127 256.663
R2036 B.n1097 B.n126 256.663
R2037 B.n1097 B.n125 256.663
R2038 B.n1097 B.n124 256.663
R2039 B.n1097 B.n123 256.663
R2040 B.n1097 B.n122 256.663
R2041 B.n1097 B.n121 256.663
R2042 B.n1097 B.n120 256.663
R2043 B.n1097 B.n119 256.663
R2044 B.n1097 B.n118 256.663
R2045 B.n1097 B.n117 256.663
R2046 B.n1097 B.n116 256.663
R2047 B.n1097 B.n115 256.663
R2048 B.n1097 B.n114 256.663
R2049 B.n1097 B.n113 256.663
R2050 B.n1097 B.n112 256.663
R2051 B.n596 B.n530 256.663
R2052 B.n602 B.n530 256.663
R2053 B.n604 B.n530 256.663
R2054 B.n610 B.n530 256.663
R2055 B.n612 B.n530 256.663
R2056 B.n618 B.n530 256.663
R2057 B.n620 B.n530 256.663
R2058 B.n626 B.n530 256.663
R2059 B.n628 B.n530 256.663
R2060 B.n634 B.n530 256.663
R2061 B.n636 B.n530 256.663
R2062 B.n642 B.n530 256.663
R2063 B.n644 B.n530 256.663
R2064 B.n650 B.n530 256.663
R2065 B.n652 B.n530 256.663
R2066 B.n658 B.n530 256.663
R2067 B.n660 B.n530 256.663
R2068 B.n666 B.n530 256.663
R2069 B.n668 B.n530 256.663
R2070 B.n674 B.n530 256.663
R2071 B.n676 B.n530 256.663
R2072 B.n682 B.n530 256.663
R2073 B.n684 B.n530 256.663
R2074 B.n690 B.n530 256.663
R2075 B.n692 B.n530 256.663
R2076 B.n698 B.n530 256.663
R2077 B.n700 B.n530 256.663
R2078 B.n707 B.n530 256.663
R2079 B.n709 B.n530 256.663
R2080 B.n715 B.n530 256.663
R2081 B.n717 B.n530 256.663
R2082 B.n723 B.n530 256.663
R2083 B.n725 B.n530 256.663
R2084 B.n731 B.n530 256.663
R2085 B.n733 B.n530 256.663
R2086 B.n739 B.n530 256.663
R2087 B.n741 B.n530 256.663
R2088 B.n747 B.n530 256.663
R2089 B.n749 B.n530 256.663
R2090 B.n755 B.n530 256.663
R2091 B.n757 B.n530 256.663
R2092 B.n763 B.n530 256.663
R2093 B.n765 B.n530 256.663
R2094 B.n771 B.n530 256.663
R2095 B.n773 B.n530 256.663
R2096 B.n779 B.n530 256.663
R2097 B.n781 B.n530 256.663
R2098 B.n787 B.n530 256.663
R2099 B.n789 B.n530 256.663
R2100 B.n795 B.n530 256.663
R2101 B.n797 B.n530 256.663
R2102 B.n803 B.n530 256.663
R2103 B.n805 B.n530 256.663
R2104 B.n811 B.n530 256.663
R2105 B.n813 B.n530 256.663
R2106 B.n819 B.n530 256.663
R2107 B.n821 B.n530 256.663
R2108 B.n827 B.n530 256.663
R2109 B.n830 B.n530 256.663
R2110 B.n1222 B.n1221 256.663
R2111 B.n178 B.n177 163.367
R2112 B.n182 B.n181 163.367
R2113 B.n186 B.n185 163.367
R2114 B.n190 B.n189 163.367
R2115 B.n194 B.n193 163.367
R2116 B.n198 B.n197 163.367
R2117 B.n202 B.n201 163.367
R2118 B.n206 B.n205 163.367
R2119 B.n210 B.n209 163.367
R2120 B.n214 B.n213 163.367
R2121 B.n218 B.n217 163.367
R2122 B.n222 B.n221 163.367
R2123 B.n226 B.n225 163.367
R2124 B.n230 B.n229 163.367
R2125 B.n234 B.n233 163.367
R2126 B.n238 B.n237 163.367
R2127 B.n242 B.n241 163.367
R2128 B.n246 B.n245 163.367
R2129 B.n250 B.n249 163.367
R2130 B.n254 B.n253 163.367
R2131 B.n258 B.n257 163.367
R2132 B.n262 B.n261 163.367
R2133 B.n266 B.n265 163.367
R2134 B.n270 B.n269 163.367
R2135 B.n274 B.n273 163.367
R2136 B.n278 B.n277 163.367
R2137 B.n282 B.n281 163.367
R2138 B.n287 B.n286 163.367
R2139 B.n291 B.n290 163.367
R2140 B.n295 B.n294 163.367
R2141 B.n299 B.n298 163.367
R2142 B.n303 B.n302 163.367
R2143 B.n308 B.n307 163.367
R2144 B.n312 B.n311 163.367
R2145 B.n316 B.n315 163.367
R2146 B.n320 B.n319 163.367
R2147 B.n324 B.n323 163.367
R2148 B.n328 B.n327 163.367
R2149 B.n332 B.n331 163.367
R2150 B.n336 B.n335 163.367
R2151 B.n340 B.n339 163.367
R2152 B.n344 B.n343 163.367
R2153 B.n348 B.n347 163.367
R2154 B.n352 B.n351 163.367
R2155 B.n356 B.n355 163.367
R2156 B.n360 B.n359 163.367
R2157 B.n364 B.n363 163.367
R2158 B.n368 B.n367 163.367
R2159 B.n372 B.n371 163.367
R2160 B.n376 B.n375 163.367
R2161 B.n380 B.n379 163.367
R2162 B.n384 B.n383 163.367
R2163 B.n388 B.n387 163.367
R2164 B.n392 B.n391 163.367
R2165 B.n396 B.n395 163.367
R2166 B.n400 B.n399 163.367
R2167 B.n404 B.n403 163.367
R2168 B.n408 B.n407 163.367
R2169 B.n410 B.n171 163.367
R2170 B.n835 B.n525 163.367
R2171 B.n843 B.n525 163.367
R2172 B.n843 B.n523 163.367
R2173 B.n847 B.n523 163.367
R2174 B.n847 B.n517 163.367
R2175 B.n855 B.n517 163.367
R2176 B.n855 B.n515 163.367
R2177 B.n859 B.n515 163.367
R2178 B.n859 B.n509 163.367
R2179 B.n867 B.n509 163.367
R2180 B.n867 B.n507 163.367
R2181 B.n871 B.n507 163.367
R2182 B.n871 B.n501 163.367
R2183 B.n879 B.n501 163.367
R2184 B.n879 B.n499 163.367
R2185 B.n883 B.n499 163.367
R2186 B.n883 B.n493 163.367
R2187 B.n891 B.n493 163.367
R2188 B.n891 B.n491 163.367
R2189 B.n895 B.n491 163.367
R2190 B.n895 B.n485 163.367
R2191 B.n903 B.n485 163.367
R2192 B.n903 B.n483 163.367
R2193 B.n907 B.n483 163.367
R2194 B.n907 B.n477 163.367
R2195 B.n915 B.n477 163.367
R2196 B.n915 B.n475 163.367
R2197 B.n919 B.n475 163.367
R2198 B.n919 B.n469 163.367
R2199 B.n927 B.n469 163.367
R2200 B.n927 B.n467 163.367
R2201 B.n931 B.n467 163.367
R2202 B.n931 B.n461 163.367
R2203 B.n939 B.n461 163.367
R2204 B.n939 B.n459 163.367
R2205 B.n943 B.n459 163.367
R2206 B.n943 B.n453 163.367
R2207 B.n951 B.n453 163.367
R2208 B.n951 B.n451 163.367
R2209 B.n955 B.n451 163.367
R2210 B.n955 B.n444 163.367
R2211 B.n963 B.n444 163.367
R2212 B.n963 B.n442 163.367
R2213 B.n967 B.n442 163.367
R2214 B.n967 B.n437 163.367
R2215 B.n975 B.n437 163.367
R2216 B.n975 B.n435 163.367
R2217 B.n979 B.n435 163.367
R2218 B.n979 B.n429 163.367
R2219 B.n987 B.n429 163.367
R2220 B.n987 B.n427 163.367
R2221 B.n991 B.n427 163.367
R2222 B.n991 B.n422 163.367
R2223 B.n1000 B.n422 163.367
R2224 B.n1000 B.n420 163.367
R2225 B.n1005 B.n420 163.367
R2226 B.n1005 B.n414 163.367
R2227 B.n1013 B.n414 163.367
R2228 B.n1014 B.n1013 163.367
R2229 B.n1014 B.n5 163.367
R2230 B.n6 B.n5 163.367
R2231 B.n7 B.n6 163.367
R2232 B.n1020 B.n7 163.367
R2233 B.n1021 B.n1020 163.367
R2234 B.n1021 B.n13 163.367
R2235 B.n14 B.n13 163.367
R2236 B.n15 B.n14 163.367
R2237 B.n1026 B.n15 163.367
R2238 B.n1026 B.n20 163.367
R2239 B.n21 B.n20 163.367
R2240 B.n22 B.n21 163.367
R2241 B.n1031 B.n22 163.367
R2242 B.n1031 B.n27 163.367
R2243 B.n28 B.n27 163.367
R2244 B.n29 B.n28 163.367
R2245 B.n1036 B.n29 163.367
R2246 B.n1036 B.n34 163.367
R2247 B.n35 B.n34 163.367
R2248 B.n36 B.n35 163.367
R2249 B.n1041 B.n36 163.367
R2250 B.n1041 B.n41 163.367
R2251 B.n42 B.n41 163.367
R2252 B.n43 B.n42 163.367
R2253 B.n1046 B.n43 163.367
R2254 B.n1046 B.n48 163.367
R2255 B.n49 B.n48 163.367
R2256 B.n50 B.n49 163.367
R2257 B.n1051 B.n50 163.367
R2258 B.n1051 B.n55 163.367
R2259 B.n56 B.n55 163.367
R2260 B.n57 B.n56 163.367
R2261 B.n1056 B.n57 163.367
R2262 B.n1056 B.n62 163.367
R2263 B.n63 B.n62 163.367
R2264 B.n64 B.n63 163.367
R2265 B.n1061 B.n64 163.367
R2266 B.n1061 B.n69 163.367
R2267 B.n70 B.n69 163.367
R2268 B.n71 B.n70 163.367
R2269 B.n1066 B.n71 163.367
R2270 B.n1066 B.n76 163.367
R2271 B.n77 B.n76 163.367
R2272 B.n78 B.n77 163.367
R2273 B.n1071 B.n78 163.367
R2274 B.n1071 B.n83 163.367
R2275 B.n84 B.n83 163.367
R2276 B.n85 B.n84 163.367
R2277 B.n1076 B.n85 163.367
R2278 B.n1076 B.n90 163.367
R2279 B.n91 B.n90 163.367
R2280 B.n92 B.n91 163.367
R2281 B.n1081 B.n92 163.367
R2282 B.n1081 B.n97 163.367
R2283 B.n98 B.n97 163.367
R2284 B.n99 B.n98 163.367
R2285 B.n1086 B.n99 163.367
R2286 B.n1086 B.n104 163.367
R2287 B.n105 B.n104 163.367
R2288 B.n106 B.n105 163.367
R2289 B.n1091 B.n106 163.367
R2290 B.n1091 B.n111 163.367
R2291 B.n597 B.n595 163.367
R2292 B.n601 B.n595 163.367
R2293 B.n605 B.n603 163.367
R2294 B.n609 B.n593 163.367
R2295 B.n613 B.n611 163.367
R2296 B.n617 B.n591 163.367
R2297 B.n621 B.n619 163.367
R2298 B.n625 B.n589 163.367
R2299 B.n629 B.n627 163.367
R2300 B.n633 B.n587 163.367
R2301 B.n637 B.n635 163.367
R2302 B.n641 B.n585 163.367
R2303 B.n645 B.n643 163.367
R2304 B.n649 B.n583 163.367
R2305 B.n653 B.n651 163.367
R2306 B.n657 B.n581 163.367
R2307 B.n661 B.n659 163.367
R2308 B.n665 B.n579 163.367
R2309 B.n669 B.n667 163.367
R2310 B.n673 B.n577 163.367
R2311 B.n677 B.n675 163.367
R2312 B.n681 B.n575 163.367
R2313 B.n685 B.n683 163.367
R2314 B.n689 B.n573 163.367
R2315 B.n693 B.n691 163.367
R2316 B.n697 B.n571 163.367
R2317 B.n701 B.n699 163.367
R2318 B.n706 B.n567 163.367
R2319 B.n710 B.n708 163.367
R2320 B.n714 B.n565 163.367
R2321 B.n718 B.n716 163.367
R2322 B.n722 B.n563 163.367
R2323 B.n726 B.n724 163.367
R2324 B.n730 B.n558 163.367
R2325 B.n734 B.n732 163.367
R2326 B.n738 B.n556 163.367
R2327 B.n742 B.n740 163.367
R2328 B.n746 B.n554 163.367
R2329 B.n750 B.n748 163.367
R2330 B.n754 B.n552 163.367
R2331 B.n758 B.n756 163.367
R2332 B.n762 B.n550 163.367
R2333 B.n766 B.n764 163.367
R2334 B.n770 B.n548 163.367
R2335 B.n774 B.n772 163.367
R2336 B.n778 B.n546 163.367
R2337 B.n782 B.n780 163.367
R2338 B.n786 B.n544 163.367
R2339 B.n790 B.n788 163.367
R2340 B.n794 B.n542 163.367
R2341 B.n798 B.n796 163.367
R2342 B.n802 B.n540 163.367
R2343 B.n806 B.n804 163.367
R2344 B.n810 B.n538 163.367
R2345 B.n814 B.n812 163.367
R2346 B.n818 B.n536 163.367
R2347 B.n822 B.n820 163.367
R2348 B.n826 B.n534 163.367
R2349 B.n829 B.n828 163.367
R2350 B.n831 B.n531 163.367
R2351 B.n837 B.n527 163.367
R2352 B.n841 B.n527 163.367
R2353 B.n841 B.n521 163.367
R2354 B.n849 B.n521 163.367
R2355 B.n849 B.n519 163.367
R2356 B.n853 B.n519 163.367
R2357 B.n853 B.n513 163.367
R2358 B.n861 B.n513 163.367
R2359 B.n861 B.n511 163.367
R2360 B.n865 B.n511 163.367
R2361 B.n865 B.n505 163.367
R2362 B.n873 B.n505 163.367
R2363 B.n873 B.n503 163.367
R2364 B.n877 B.n503 163.367
R2365 B.n877 B.n497 163.367
R2366 B.n885 B.n497 163.367
R2367 B.n885 B.n495 163.367
R2368 B.n889 B.n495 163.367
R2369 B.n889 B.n489 163.367
R2370 B.n897 B.n489 163.367
R2371 B.n897 B.n487 163.367
R2372 B.n901 B.n487 163.367
R2373 B.n901 B.n481 163.367
R2374 B.n909 B.n481 163.367
R2375 B.n909 B.n479 163.367
R2376 B.n913 B.n479 163.367
R2377 B.n913 B.n473 163.367
R2378 B.n921 B.n473 163.367
R2379 B.n921 B.n471 163.367
R2380 B.n925 B.n471 163.367
R2381 B.n925 B.n465 163.367
R2382 B.n933 B.n465 163.367
R2383 B.n933 B.n463 163.367
R2384 B.n937 B.n463 163.367
R2385 B.n937 B.n457 163.367
R2386 B.n945 B.n457 163.367
R2387 B.n945 B.n455 163.367
R2388 B.n949 B.n455 163.367
R2389 B.n949 B.n449 163.367
R2390 B.n957 B.n449 163.367
R2391 B.n957 B.n447 163.367
R2392 B.n961 B.n447 163.367
R2393 B.n961 B.n441 163.367
R2394 B.n969 B.n441 163.367
R2395 B.n969 B.n439 163.367
R2396 B.n973 B.n439 163.367
R2397 B.n973 B.n433 163.367
R2398 B.n981 B.n433 163.367
R2399 B.n981 B.n431 163.367
R2400 B.n985 B.n431 163.367
R2401 B.n985 B.n425 163.367
R2402 B.n994 B.n425 163.367
R2403 B.n994 B.n423 163.367
R2404 B.n998 B.n423 163.367
R2405 B.n998 B.n418 163.367
R2406 B.n1007 B.n418 163.367
R2407 B.n1007 B.n416 163.367
R2408 B.n1011 B.n416 163.367
R2409 B.n1011 B.n3 163.367
R2410 B.n1220 B.n3 163.367
R2411 B.n1216 B.n2 163.367
R2412 B.n1216 B.n1215 163.367
R2413 B.n1215 B.n9 163.367
R2414 B.n1211 B.n9 163.367
R2415 B.n1211 B.n11 163.367
R2416 B.n1207 B.n11 163.367
R2417 B.n1207 B.n16 163.367
R2418 B.n1203 B.n16 163.367
R2419 B.n1203 B.n18 163.367
R2420 B.n1199 B.n18 163.367
R2421 B.n1199 B.n24 163.367
R2422 B.n1195 B.n24 163.367
R2423 B.n1195 B.n26 163.367
R2424 B.n1191 B.n26 163.367
R2425 B.n1191 B.n31 163.367
R2426 B.n1187 B.n31 163.367
R2427 B.n1187 B.n33 163.367
R2428 B.n1183 B.n33 163.367
R2429 B.n1183 B.n38 163.367
R2430 B.n1179 B.n38 163.367
R2431 B.n1179 B.n40 163.367
R2432 B.n1175 B.n40 163.367
R2433 B.n1175 B.n45 163.367
R2434 B.n1171 B.n45 163.367
R2435 B.n1171 B.n47 163.367
R2436 B.n1167 B.n47 163.367
R2437 B.n1167 B.n52 163.367
R2438 B.n1163 B.n52 163.367
R2439 B.n1163 B.n54 163.367
R2440 B.n1159 B.n54 163.367
R2441 B.n1159 B.n59 163.367
R2442 B.n1155 B.n59 163.367
R2443 B.n1155 B.n61 163.367
R2444 B.n1151 B.n61 163.367
R2445 B.n1151 B.n66 163.367
R2446 B.n1147 B.n66 163.367
R2447 B.n1147 B.n68 163.367
R2448 B.n1143 B.n68 163.367
R2449 B.n1143 B.n73 163.367
R2450 B.n1139 B.n73 163.367
R2451 B.n1139 B.n75 163.367
R2452 B.n1135 B.n75 163.367
R2453 B.n1135 B.n80 163.367
R2454 B.n1131 B.n80 163.367
R2455 B.n1131 B.n82 163.367
R2456 B.n1127 B.n82 163.367
R2457 B.n1127 B.n87 163.367
R2458 B.n1123 B.n87 163.367
R2459 B.n1123 B.n89 163.367
R2460 B.n1119 B.n89 163.367
R2461 B.n1119 B.n94 163.367
R2462 B.n1115 B.n94 163.367
R2463 B.n1115 B.n96 163.367
R2464 B.n1111 B.n96 163.367
R2465 B.n1111 B.n101 163.367
R2466 B.n1107 B.n101 163.367
R2467 B.n1107 B.n103 163.367
R2468 B.n1103 B.n103 163.367
R2469 B.n1103 B.n108 163.367
R2470 B.n1099 B.n108 163.367
R2471 B.n112 B.n110 71.676
R2472 B.n178 B.n113 71.676
R2473 B.n182 B.n114 71.676
R2474 B.n186 B.n115 71.676
R2475 B.n190 B.n116 71.676
R2476 B.n194 B.n117 71.676
R2477 B.n198 B.n118 71.676
R2478 B.n202 B.n119 71.676
R2479 B.n206 B.n120 71.676
R2480 B.n210 B.n121 71.676
R2481 B.n214 B.n122 71.676
R2482 B.n218 B.n123 71.676
R2483 B.n222 B.n124 71.676
R2484 B.n226 B.n125 71.676
R2485 B.n230 B.n126 71.676
R2486 B.n234 B.n127 71.676
R2487 B.n238 B.n128 71.676
R2488 B.n242 B.n129 71.676
R2489 B.n246 B.n130 71.676
R2490 B.n250 B.n131 71.676
R2491 B.n254 B.n132 71.676
R2492 B.n258 B.n133 71.676
R2493 B.n262 B.n134 71.676
R2494 B.n266 B.n135 71.676
R2495 B.n270 B.n136 71.676
R2496 B.n274 B.n137 71.676
R2497 B.n278 B.n138 71.676
R2498 B.n282 B.n139 71.676
R2499 B.n287 B.n140 71.676
R2500 B.n291 B.n141 71.676
R2501 B.n295 B.n142 71.676
R2502 B.n299 B.n143 71.676
R2503 B.n303 B.n144 71.676
R2504 B.n308 B.n145 71.676
R2505 B.n312 B.n146 71.676
R2506 B.n316 B.n147 71.676
R2507 B.n320 B.n148 71.676
R2508 B.n324 B.n149 71.676
R2509 B.n328 B.n150 71.676
R2510 B.n332 B.n151 71.676
R2511 B.n336 B.n152 71.676
R2512 B.n340 B.n153 71.676
R2513 B.n344 B.n154 71.676
R2514 B.n348 B.n155 71.676
R2515 B.n352 B.n156 71.676
R2516 B.n356 B.n157 71.676
R2517 B.n360 B.n158 71.676
R2518 B.n364 B.n159 71.676
R2519 B.n368 B.n160 71.676
R2520 B.n372 B.n161 71.676
R2521 B.n376 B.n162 71.676
R2522 B.n380 B.n163 71.676
R2523 B.n384 B.n164 71.676
R2524 B.n388 B.n165 71.676
R2525 B.n392 B.n166 71.676
R2526 B.n396 B.n167 71.676
R2527 B.n400 B.n168 71.676
R2528 B.n404 B.n169 71.676
R2529 B.n408 B.n170 71.676
R2530 B.n1096 B.n171 71.676
R2531 B.n1096 B.n1095 71.676
R2532 B.n410 B.n170 71.676
R2533 B.n407 B.n169 71.676
R2534 B.n403 B.n168 71.676
R2535 B.n399 B.n167 71.676
R2536 B.n395 B.n166 71.676
R2537 B.n391 B.n165 71.676
R2538 B.n387 B.n164 71.676
R2539 B.n383 B.n163 71.676
R2540 B.n379 B.n162 71.676
R2541 B.n375 B.n161 71.676
R2542 B.n371 B.n160 71.676
R2543 B.n367 B.n159 71.676
R2544 B.n363 B.n158 71.676
R2545 B.n359 B.n157 71.676
R2546 B.n355 B.n156 71.676
R2547 B.n351 B.n155 71.676
R2548 B.n347 B.n154 71.676
R2549 B.n343 B.n153 71.676
R2550 B.n339 B.n152 71.676
R2551 B.n335 B.n151 71.676
R2552 B.n331 B.n150 71.676
R2553 B.n327 B.n149 71.676
R2554 B.n323 B.n148 71.676
R2555 B.n319 B.n147 71.676
R2556 B.n315 B.n146 71.676
R2557 B.n311 B.n145 71.676
R2558 B.n307 B.n144 71.676
R2559 B.n302 B.n143 71.676
R2560 B.n298 B.n142 71.676
R2561 B.n294 B.n141 71.676
R2562 B.n290 B.n140 71.676
R2563 B.n286 B.n139 71.676
R2564 B.n281 B.n138 71.676
R2565 B.n277 B.n137 71.676
R2566 B.n273 B.n136 71.676
R2567 B.n269 B.n135 71.676
R2568 B.n265 B.n134 71.676
R2569 B.n261 B.n133 71.676
R2570 B.n257 B.n132 71.676
R2571 B.n253 B.n131 71.676
R2572 B.n249 B.n130 71.676
R2573 B.n245 B.n129 71.676
R2574 B.n241 B.n128 71.676
R2575 B.n237 B.n127 71.676
R2576 B.n233 B.n126 71.676
R2577 B.n229 B.n125 71.676
R2578 B.n225 B.n124 71.676
R2579 B.n221 B.n123 71.676
R2580 B.n217 B.n122 71.676
R2581 B.n213 B.n121 71.676
R2582 B.n209 B.n120 71.676
R2583 B.n205 B.n119 71.676
R2584 B.n201 B.n118 71.676
R2585 B.n197 B.n117 71.676
R2586 B.n193 B.n116 71.676
R2587 B.n189 B.n115 71.676
R2588 B.n185 B.n114 71.676
R2589 B.n181 B.n113 71.676
R2590 B.n177 B.n112 71.676
R2591 B.n596 B.n529 71.676
R2592 B.n602 B.n601 71.676
R2593 B.n605 B.n604 71.676
R2594 B.n610 B.n609 71.676
R2595 B.n613 B.n612 71.676
R2596 B.n618 B.n617 71.676
R2597 B.n621 B.n620 71.676
R2598 B.n626 B.n625 71.676
R2599 B.n629 B.n628 71.676
R2600 B.n634 B.n633 71.676
R2601 B.n637 B.n636 71.676
R2602 B.n642 B.n641 71.676
R2603 B.n645 B.n644 71.676
R2604 B.n650 B.n649 71.676
R2605 B.n653 B.n652 71.676
R2606 B.n658 B.n657 71.676
R2607 B.n661 B.n660 71.676
R2608 B.n666 B.n665 71.676
R2609 B.n669 B.n668 71.676
R2610 B.n674 B.n673 71.676
R2611 B.n677 B.n676 71.676
R2612 B.n682 B.n681 71.676
R2613 B.n685 B.n684 71.676
R2614 B.n690 B.n689 71.676
R2615 B.n693 B.n692 71.676
R2616 B.n698 B.n697 71.676
R2617 B.n701 B.n700 71.676
R2618 B.n707 B.n706 71.676
R2619 B.n710 B.n709 71.676
R2620 B.n715 B.n714 71.676
R2621 B.n718 B.n717 71.676
R2622 B.n723 B.n722 71.676
R2623 B.n726 B.n725 71.676
R2624 B.n731 B.n730 71.676
R2625 B.n734 B.n733 71.676
R2626 B.n739 B.n738 71.676
R2627 B.n742 B.n741 71.676
R2628 B.n747 B.n746 71.676
R2629 B.n750 B.n749 71.676
R2630 B.n755 B.n754 71.676
R2631 B.n758 B.n757 71.676
R2632 B.n763 B.n762 71.676
R2633 B.n766 B.n765 71.676
R2634 B.n771 B.n770 71.676
R2635 B.n774 B.n773 71.676
R2636 B.n779 B.n778 71.676
R2637 B.n782 B.n781 71.676
R2638 B.n787 B.n786 71.676
R2639 B.n790 B.n789 71.676
R2640 B.n795 B.n794 71.676
R2641 B.n798 B.n797 71.676
R2642 B.n803 B.n802 71.676
R2643 B.n806 B.n805 71.676
R2644 B.n811 B.n810 71.676
R2645 B.n814 B.n813 71.676
R2646 B.n819 B.n818 71.676
R2647 B.n822 B.n821 71.676
R2648 B.n827 B.n826 71.676
R2649 B.n830 B.n829 71.676
R2650 B.n597 B.n596 71.676
R2651 B.n603 B.n602 71.676
R2652 B.n604 B.n593 71.676
R2653 B.n611 B.n610 71.676
R2654 B.n612 B.n591 71.676
R2655 B.n619 B.n618 71.676
R2656 B.n620 B.n589 71.676
R2657 B.n627 B.n626 71.676
R2658 B.n628 B.n587 71.676
R2659 B.n635 B.n634 71.676
R2660 B.n636 B.n585 71.676
R2661 B.n643 B.n642 71.676
R2662 B.n644 B.n583 71.676
R2663 B.n651 B.n650 71.676
R2664 B.n652 B.n581 71.676
R2665 B.n659 B.n658 71.676
R2666 B.n660 B.n579 71.676
R2667 B.n667 B.n666 71.676
R2668 B.n668 B.n577 71.676
R2669 B.n675 B.n674 71.676
R2670 B.n676 B.n575 71.676
R2671 B.n683 B.n682 71.676
R2672 B.n684 B.n573 71.676
R2673 B.n691 B.n690 71.676
R2674 B.n692 B.n571 71.676
R2675 B.n699 B.n698 71.676
R2676 B.n700 B.n567 71.676
R2677 B.n708 B.n707 71.676
R2678 B.n709 B.n565 71.676
R2679 B.n716 B.n715 71.676
R2680 B.n717 B.n563 71.676
R2681 B.n724 B.n723 71.676
R2682 B.n725 B.n558 71.676
R2683 B.n732 B.n731 71.676
R2684 B.n733 B.n556 71.676
R2685 B.n740 B.n739 71.676
R2686 B.n741 B.n554 71.676
R2687 B.n748 B.n747 71.676
R2688 B.n749 B.n552 71.676
R2689 B.n756 B.n755 71.676
R2690 B.n757 B.n550 71.676
R2691 B.n764 B.n763 71.676
R2692 B.n765 B.n548 71.676
R2693 B.n772 B.n771 71.676
R2694 B.n773 B.n546 71.676
R2695 B.n780 B.n779 71.676
R2696 B.n781 B.n544 71.676
R2697 B.n788 B.n787 71.676
R2698 B.n789 B.n542 71.676
R2699 B.n796 B.n795 71.676
R2700 B.n797 B.n540 71.676
R2701 B.n804 B.n803 71.676
R2702 B.n805 B.n538 71.676
R2703 B.n812 B.n811 71.676
R2704 B.n813 B.n536 71.676
R2705 B.n820 B.n819 71.676
R2706 B.n821 B.n534 71.676
R2707 B.n828 B.n827 71.676
R2708 B.n831 B.n830 71.676
R2709 B.n1221 B.n1220 71.676
R2710 B.n1221 B.n2 71.676
R2711 B.n175 B.n174 68.849
R2712 B.n173 B.n172 68.849
R2713 B.n560 B.n559 68.849
R2714 B.n569 B.n568 68.849
R2715 B.n284 B.n175 59.5399
R2716 B.n305 B.n173 59.5399
R2717 B.n561 B.n560 59.5399
R2718 B.n704 B.n569 59.5399
R2719 B.n836 B.n530 55.665
R2720 B.n1098 B.n1097 55.665
R2721 B.n836 B.n526 34.1013
R2722 B.n842 B.n526 34.1013
R2723 B.n842 B.n522 34.1013
R2724 B.n848 B.n522 34.1013
R2725 B.n848 B.n518 34.1013
R2726 B.n854 B.n518 34.1013
R2727 B.n854 B.n514 34.1013
R2728 B.n860 B.n514 34.1013
R2729 B.n866 B.n510 34.1013
R2730 B.n866 B.n506 34.1013
R2731 B.n872 B.n506 34.1013
R2732 B.n872 B.n502 34.1013
R2733 B.n878 B.n502 34.1013
R2734 B.n878 B.n498 34.1013
R2735 B.n884 B.n498 34.1013
R2736 B.n884 B.n494 34.1013
R2737 B.n890 B.n494 34.1013
R2738 B.n890 B.n490 34.1013
R2739 B.n896 B.n490 34.1013
R2740 B.n896 B.n486 34.1013
R2741 B.n902 B.n486 34.1013
R2742 B.n908 B.n482 34.1013
R2743 B.n908 B.n478 34.1013
R2744 B.n914 B.n478 34.1013
R2745 B.n914 B.n474 34.1013
R2746 B.n920 B.n474 34.1013
R2747 B.n920 B.n470 34.1013
R2748 B.n926 B.n470 34.1013
R2749 B.n926 B.n466 34.1013
R2750 B.n932 B.n466 34.1013
R2751 B.n938 B.n462 34.1013
R2752 B.n938 B.n458 34.1013
R2753 B.n944 B.n458 34.1013
R2754 B.n944 B.n454 34.1013
R2755 B.n950 B.n454 34.1013
R2756 B.n950 B.n450 34.1013
R2757 B.n956 B.n450 34.1013
R2758 B.n956 B.n445 34.1013
R2759 B.n962 B.n445 34.1013
R2760 B.n962 B.n446 34.1013
R2761 B.n968 B.n438 34.1013
R2762 B.n974 B.n438 34.1013
R2763 B.n974 B.n434 34.1013
R2764 B.n980 B.n434 34.1013
R2765 B.n980 B.n430 34.1013
R2766 B.n986 B.n430 34.1013
R2767 B.n986 B.n426 34.1013
R2768 B.n993 B.n426 34.1013
R2769 B.n993 B.n992 34.1013
R2770 B.n999 B.n419 34.1013
R2771 B.n1006 B.n419 34.1013
R2772 B.n1006 B.n415 34.1013
R2773 B.n1012 B.n415 34.1013
R2774 B.n1012 B.n4 34.1013
R2775 B.n1219 B.n4 34.1013
R2776 B.n1219 B.n1218 34.1013
R2777 B.n1218 B.n1217 34.1013
R2778 B.n1217 B.n8 34.1013
R2779 B.n12 B.n8 34.1013
R2780 B.n1210 B.n12 34.1013
R2781 B.n1210 B.n1209 34.1013
R2782 B.n1209 B.n1208 34.1013
R2783 B.n1202 B.n19 34.1013
R2784 B.n1202 B.n1201 34.1013
R2785 B.n1201 B.n1200 34.1013
R2786 B.n1200 B.n23 34.1013
R2787 B.n1194 B.n23 34.1013
R2788 B.n1194 B.n1193 34.1013
R2789 B.n1193 B.n1192 34.1013
R2790 B.n1192 B.n30 34.1013
R2791 B.n1186 B.n30 34.1013
R2792 B.n1185 B.n1184 34.1013
R2793 B.n1184 B.n37 34.1013
R2794 B.n1178 B.n37 34.1013
R2795 B.n1178 B.n1177 34.1013
R2796 B.n1177 B.n1176 34.1013
R2797 B.n1176 B.n44 34.1013
R2798 B.n1170 B.n44 34.1013
R2799 B.n1170 B.n1169 34.1013
R2800 B.n1169 B.n1168 34.1013
R2801 B.n1168 B.n51 34.1013
R2802 B.n1162 B.n1161 34.1013
R2803 B.n1161 B.n1160 34.1013
R2804 B.n1160 B.n58 34.1013
R2805 B.n1154 B.n58 34.1013
R2806 B.n1154 B.n1153 34.1013
R2807 B.n1153 B.n1152 34.1013
R2808 B.n1152 B.n65 34.1013
R2809 B.n1146 B.n65 34.1013
R2810 B.n1146 B.n1145 34.1013
R2811 B.n1144 B.n72 34.1013
R2812 B.n1138 B.n72 34.1013
R2813 B.n1138 B.n1137 34.1013
R2814 B.n1137 B.n1136 34.1013
R2815 B.n1136 B.n79 34.1013
R2816 B.n1130 B.n79 34.1013
R2817 B.n1130 B.n1129 34.1013
R2818 B.n1129 B.n1128 34.1013
R2819 B.n1128 B.n86 34.1013
R2820 B.n1122 B.n86 34.1013
R2821 B.n1122 B.n1121 34.1013
R2822 B.n1121 B.n1120 34.1013
R2823 B.n1120 B.n93 34.1013
R2824 B.n1114 B.n1113 34.1013
R2825 B.n1113 B.n1112 34.1013
R2826 B.n1112 B.n100 34.1013
R2827 B.n1106 B.n100 34.1013
R2828 B.n1106 B.n1105 34.1013
R2829 B.n1105 B.n1104 34.1013
R2830 B.n1104 B.n107 34.1013
R2831 B.n1098 B.n107 34.1013
R2832 B.n838 B.n528 31.6883
R2833 B.n834 B.n833 31.6883
R2834 B.n1094 B.n1093 31.6883
R2835 B.n1100 B.n109 31.6883
R2836 B.n932 B.t4 27.0805
R2837 B.n1162 B.t0 27.0805
R2838 B.n968 B.t21 26.0775
R2839 B.n1186 B.t2 26.0775
R2840 B.n860 B.t8 24.0716
R2841 B.n1114 B.t12 24.0716
R2842 B.n992 B.t6 23.0687
R2843 B.n19 B.t5 23.0687
R2844 B.t3 B.n482 22.0657
R2845 B.n1145 B.t1 22.0657
R2846 B B.n1222 18.0485
R2847 B.n902 B.t3 12.0361
R2848 B.t1 B.n1144 12.0361
R2849 B.n999 B.t6 11.0331
R2850 B.n1208 B.t5 11.0331
R2851 B.n839 B.n838 10.6151
R2852 B.n840 B.n839 10.6151
R2853 B.n840 B.n520 10.6151
R2854 B.n850 B.n520 10.6151
R2855 B.n851 B.n850 10.6151
R2856 B.n852 B.n851 10.6151
R2857 B.n852 B.n512 10.6151
R2858 B.n862 B.n512 10.6151
R2859 B.n863 B.n862 10.6151
R2860 B.n864 B.n863 10.6151
R2861 B.n864 B.n504 10.6151
R2862 B.n874 B.n504 10.6151
R2863 B.n875 B.n874 10.6151
R2864 B.n876 B.n875 10.6151
R2865 B.n876 B.n496 10.6151
R2866 B.n886 B.n496 10.6151
R2867 B.n887 B.n886 10.6151
R2868 B.n888 B.n887 10.6151
R2869 B.n888 B.n488 10.6151
R2870 B.n898 B.n488 10.6151
R2871 B.n899 B.n898 10.6151
R2872 B.n900 B.n899 10.6151
R2873 B.n900 B.n480 10.6151
R2874 B.n910 B.n480 10.6151
R2875 B.n911 B.n910 10.6151
R2876 B.n912 B.n911 10.6151
R2877 B.n912 B.n472 10.6151
R2878 B.n922 B.n472 10.6151
R2879 B.n923 B.n922 10.6151
R2880 B.n924 B.n923 10.6151
R2881 B.n924 B.n464 10.6151
R2882 B.n934 B.n464 10.6151
R2883 B.n935 B.n934 10.6151
R2884 B.n936 B.n935 10.6151
R2885 B.n936 B.n456 10.6151
R2886 B.n946 B.n456 10.6151
R2887 B.n947 B.n946 10.6151
R2888 B.n948 B.n947 10.6151
R2889 B.n948 B.n448 10.6151
R2890 B.n958 B.n448 10.6151
R2891 B.n959 B.n958 10.6151
R2892 B.n960 B.n959 10.6151
R2893 B.n960 B.n440 10.6151
R2894 B.n970 B.n440 10.6151
R2895 B.n971 B.n970 10.6151
R2896 B.n972 B.n971 10.6151
R2897 B.n972 B.n432 10.6151
R2898 B.n982 B.n432 10.6151
R2899 B.n983 B.n982 10.6151
R2900 B.n984 B.n983 10.6151
R2901 B.n984 B.n424 10.6151
R2902 B.n995 B.n424 10.6151
R2903 B.n996 B.n995 10.6151
R2904 B.n997 B.n996 10.6151
R2905 B.n997 B.n417 10.6151
R2906 B.n1008 B.n417 10.6151
R2907 B.n1009 B.n1008 10.6151
R2908 B.n1010 B.n1009 10.6151
R2909 B.n1010 B.n0 10.6151
R2910 B.n598 B.n528 10.6151
R2911 B.n599 B.n598 10.6151
R2912 B.n600 B.n599 10.6151
R2913 B.n600 B.n594 10.6151
R2914 B.n606 B.n594 10.6151
R2915 B.n607 B.n606 10.6151
R2916 B.n608 B.n607 10.6151
R2917 B.n608 B.n592 10.6151
R2918 B.n614 B.n592 10.6151
R2919 B.n615 B.n614 10.6151
R2920 B.n616 B.n615 10.6151
R2921 B.n616 B.n590 10.6151
R2922 B.n622 B.n590 10.6151
R2923 B.n623 B.n622 10.6151
R2924 B.n624 B.n623 10.6151
R2925 B.n624 B.n588 10.6151
R2926 B.n630 B.n588 10.6151
R2927 B.n631 B.n630 10.6151
R2928 B.n632 B.n631 10.6151
R2929 B.n632 B.n586 10.6151
R2930 B.n638 B.n586 10.6151
R2931 B.n639 B.n638 10.6151
R2932 B.n640 B.n639 10.6151
R2933 B.n640 B.n584 10.6151
R2934 B.n646 B.n584 10.6151
R2935 B.n647 B.n646 10.6151
R2936 B.n648 B.n647 10.6151
R2937 B.n648 B.n582 10.6151
R2938 B.n654 B.n582 10.6151
R2939 B.n655 B.n654 10.6151
R2940 B.n656 B.n655 10.6151
R2941 B.n656 B.n580 10.6151
R2942 B.n662 B.n580 10.6151
R2943 B.n663 B.n662 10.6151
R2944 B.n664 B.n663 10.6151
R2945 B.n664 B.n578 10.6151
R2946 B.n670 B.n578 10.6151
R2947 B.n671 B.n670 10.6151
R2948 B.n672 B.n671 10.6151
R2949 B.n672 B.n576 10.6151
R2950 B.n678 B.n576 10.6151
R2951 B.n679 B.n678 10.6151
R2952 B.n680 B.n679 10.6151
R2953 B.n680 B.n574 10.6151
R2954 B.n686 B.n574 10.6151
R2955 B.n687 B.n686 10.6151
R2956 B.n688 B.n687 10.6151
R2957 B.n688 B.n572 10.6151
R2958 B.n694 B.n572 10.6151
R2959 B.n695 B.n694 10.6151
R2960 B.n696 B.n695 10.6151
R2961 B.n696 B.n570 10.6151
R2962 B.n702 B.n570 10.6151
R2963 B.n703 B.n702 10.6151
R2964 B.n705 B.n566 10.6151
R2965 B.n711 B.n566 10.6151
R2966 B.n712 B.n711 10.6151
R2967 B.n713 B.n712 10.6151
R2968 B.n713 B.n564 10.6151
R2969 B.n719 B.n564 10.6151
R2970 B.n720 B.n719 10.6151
R2971 B.n721 B.n720 10.6151
R2972 B.n721 B.n562 10.6151
R2973 B.n728 B.n727 10.6151
R2974 B.n729 B.n728 10.6151
R2975 B.n729 B.n557 10.6151
R2976 B.n735 B.n557 10.6151
R2977 B.n736 B.n735 10.6151
R2978 B.n737 B.n736 10.6151
R2979 B.n737 B.n555 10.6151
R2980 B.n743 B.n555 10.6151
R2981 B.n744 B.n743 10.6151
R2982 B.n745 B.n744 10.6151
R2983 B.n745 B.n553 10.6151
R2984 B.n751 B.n553 10.6151
R2985 B.n752 B.n751 10.6151
R2986 B.n753 B.n752 10.6151
R2987 B.n753 B.n551 10.6151
R2988 B.n759 B.n551 10.6151
R2989 B.n760 B.n759 10.6151
R2990 B.n761 B.n760 10.6151
R2991 B.n761 B.n549 10.6151
R2992 B.n767 B.n549 10.6151
R2993 B.n768 B.n767 10.6151
R2994 B.n769 B.n768 10.6151
R2995 B.n769 B.n547 10.6151
R2996 B.n775 B.n547 10.6151
R2997 B.n776 B.n775 10.6151
R2998 B.n777 B.n776 10.6151
R2999 B.n777 B.n545 10.6151
R3000 B.n783 B.n545 10.6151
R3001 B.n784 B.n783 10.6151
R3002 B.n785 B.n784 10.6151
R3003 B.n785 B.n543 10.6151
R3004 B.n791 B.n543 10.6151
R3005 B.n792 B.n791 10.6151
R3006 B.n793 B.n792 10.6151
R3007 B.n793 B.n541 10.6151
R3008 B.n799 B.n541 10.6151
R3009 B.n800 B.n799 10.6151
R3010 B.n801 B.n800 10.6151
R3011 B.n801 B.n539 10.6151
R3012 B.n807 B.n539 10.6151
R3013 B.n808 B.n807 10.6151
R3014 B.n809 B.n808 10.6151
R3015 B.n809 B.n537 10.6151
R3016 B.n815 B.n537 10.6151
R3017 B.n816 B.n815 10.6151
R3018 B.n817 B.n816 10.6151
R3019 B.n817 B.n535 10.6151
R3020 B.n823 B.n535 10.6151
R3021 B.n824 B.n823 10.6151
R3022 B.n825 B.n824 10.6151
R3023 B.n825 B.n533 10.6151
R3024 B.n533 B.n532 10.6151
R3025 B.n832 B.n532 10.6151
R3026 B.n833 B.n832 10.6151
R3027 B.n834 B.n524 10.6151
R3028 B.n844 B.n524 10.6151
R3029 B.n845 B.n844 10.6151
R3030 B.n846 B.n845 10.6151
R3031 B.n846 B.n516 10.6151
R3032 B.n856 B.n516 10.6151
R3033 B.n857 B.n856 10.6151
R3034 B.n858 B.n857 10.6151
R3035 B.n858 B.n508 10.6151
R3036 B.n868 B.n508 10.6151
R3037 B.n869 B.n868 10.6151
R3038 B.n870 B.n869 10.6151
R3039 B.n870 B.n500 10.6151
R3040 B.n880 B.n500 10.6151
R3041 B.n881 B.n880 10.6151
R3042 B.n882 B.n881 10.6151
R3043 B.n882 B.n492 10.6151
R3044 B.n892 B.n492 10.6151
R3045 B.n893 B.n892 10.6151
R3046 B.n894 B.n893 10.6151
R3047 B.n894 B.n484 10.6151
R3048 B.n904 B.n484 10.6151
R3049 B.n905 B.n904 10.6151
R3050 B.n906 B.n905 10.6151
R3051 B.n906 B.n476 10.6151
R3052 B.n916 B.n476 10.6151
R3053 B.n917 B.n916 10.6151
R3054 B.n918 B.n917 10.6151
R3055 B.n918 B.n468 10.6151
R3056 B.n928 B.n468 10.6151
R3057 B.n929 B.n928 10.6151
R3058 B.n930 B.n929 10.6151
R3059 B.n930 B.n460 10.6151
R3060 B.n940 B.n460 10.6151
R3061 B.n941 B.n940 10.6151
R3062 B.n942 B.n941 10.6151
R3063 B.n942 B.n452 10.6151
R3064 B.n952 B.n452 10.6151
R3065 B.n953 B.n952 10.6151
R3066 B.n954 B.n953 10.6151
R3067 B.n954 B.n443 10.6151
R3068 B.n964 B.n443 10.6151
R3069 B.n965 B.n964 10.6151
R3070 B.n966 B.n965 10.6151
R3071 B.n966 B.n436 10.6151
R3072 B.n976 B.n436 10.6151
R3073 B.n977 B.n976 10.6151
R3074 B.n978 B.n977 10.6151
R3075 B.n978 B.n428 10.6151
R3076 B.n988 B.n428 10.6151
R3077 B.n989 B.n988 10.6151
R3078 B.n990 B.n989 10.6151
R3079 B.n990 B.n421 10.6151
R3080 B.n1001 B.n421 10.6151
R3081 B.n1002 B.n1001 10.6151
R3082 B.n1004 B.n1002 10.6151
R3083 B.n1004 B.n1003 10.6151
R3084 B.n1003 B.n413 10.6151
R3085 B.n1015 B.n413 10.6151
R3086 B.n1016 B.n1015 10.6151
R3087 B.n1017 B.n1016 10.6151
R3088 B.n1018 B.n1017 10.6151
R3089 B.n1019 B.n1018 10.6151
R3090 B.n1022 B.n1019 10.6151
R3091 B.n1023 B.n1022 10.6151
R3092 B.n1024 B.n1023 10.6151
R3093 B.n1025 B.n1024 10.6151
R3094 B.n1027 B.n1025 10.6151
R3095 B.n1028 B.n1027 10.6151
R3096 B.n1029 B.n1028 10.6151
R3097 B.n1030 B.n1029 10.6151
R3098 B.n1032 B.n1030 10.6151
R3099 B.n1033 B.n1032 10.6151
R3100 B.n1034 B.n1033 10.6151
R3101 B.n1035 B.n1034 10.6151
R3102 B.n1037 B.n1035 10.6151
R3103 B.n1038 B.n1037 10.6151
R3104 B.n1039 B.n1038 10.6151
R3105 B.n1040 B.n1039 10.6151
R3106 B.n1042 B.n1040 10.6151
R3107 B.n1043 B.n1042 10.6151
R3108 B.n1044 B.n1043 10.6151
R3109 B.n1045 B.n1044 10.6151
R3110 B.n1047 B.n1045 10.6151
R3111 B.n1048 B.n1047 10.6151
R3112 B.n1049 B.n1048 10.6151
R3113 B.n1050 B.n1049 10.6151
R3114 B.n1052 B.n1050 10.6151
R3115 B.n1053 B.n1052 10.6151
R3116 B.n1054 B.n1053 10.6151
R3117 B.n1055 B.n1054 10.6151
R3118 B.n1057 B.n1055 10.6151
R3119 B.n1058 B.n1057 10.6151
R3120 B.n1059 B.n1058 10.6151
R3121 B.n1060 B.n1059 10.6151
R3122 B.n1062 B.n1060 10.6151
R3123 B.n1063 B.n1062 10.6151
R3124 B.n1064 B.n1063 10.6151
R3125 B.n1065 B.n1064 10.6151
R3126 B.n1067 B.n1065 10.6151
R3127 B.n1068 B.n1067 10.6151
R3128 B.n1069 B.n1068 10.6151
R3129 B.n1070 B.n1069 10.6151
R3130 B.n1072 B.n1070 10.6151
R3131 B.n1073 B.n1072 10.6151
R3132 B.n1074 B.n1073 10.6151
R3133 B.n1075 B.n1074 10.6151
R3134 B.n1077 B.n1075 10.6151
R3135 B.n1078 B.n1077 10.6151
R3136 B.n1079 B.n1078 10.6151
R3137 B.n1080 B.n1079 10.6151
R3138 B.n1082 B.n1080 10.6151
R3139 B.n1083 B.n1082 10.6151
R3140 B.n1084 B.n1083 10.6151
R3141 B.n1085 B.n1084 10.6151
R3142 B.n1087 B.n1085 10.6151
R3143 B.n1088 B.n1087 10.6151
R3144 B.n1089 B.n1088 10.6151
R3145 B.n1090 B.n1089 10.6151
R3146 B.n1092 B.n1090 10.6151
R3147 B.n1093 B.n1092 10.6151
R3148 B.n1214 B.n1 10.6151
R3149 B.n1214 B.n1213 10.6151
R3150 B.n1213 B.n1212 10.6151
R3151 B.n1212 B.n10 10.6151
R3152 B.n1206 B.n10 10.6151
R3153 B.n1206 B.n1205 10.6151
R3154 B.n1205 B.n1204 10.6151
R3155 B.n1204 B.n17 10.6151
R3156 B.n1198 B.n17 10.6151
R3157 B.n1198 B.n1197 10.6151
R3158 B.n1197 B.n1196 10.6151
R3159 B.n1196 B.n25 10.6151
R3160 B.n1190 B.n25 10.6151
R3161 B.n1190 B.n1189 10.6151
R3162 B.n1189 B.n1188 10.6151
R3163 B.n1188 B.n32 10.6151
R3164 B.n1182 B.n32 10.6151
R3165 B.n1182 B.n1181 10.6151
R3166 B.n1181 B.n1180 10.6151
R3167 B.n1180 B.n39 10.6151
R3168 B.n1174 B.n39 10.6151
R3169 B.n1174 B.n1173 10.6151
R3170 B.n1173 B.n1172 10.6151
R3171 B.n1172 B.n46 10.6151
R3172 B.n1166 B.n46 10.6151
R3173 B.n1166 B.n1165 10.6151
R3174 B.n1165 B.n1164 10.6151
R3175 B.n1164 B.n53 10.6151
R3176 B.n1158 B.n53 10.6151
R3177 B.n1158 B.n1157 10.6151
R3178 B.n1157 B.n1156 10.6151
R3179 B.n1156 B.n60 10.6151
R3180 B.n1150 B.n60 10.6151
R3181 B.n1150 B.n1149 10.6151
R3182 B.n1149 B.n1148 10.6151
R3183 B.n1148 B.n67 10.6151
R3184 B.n1142 B.n67 10.6151
R3185 B.n1142 B.n1141 10.6151
R3186 B.n1141 B.n1140 10.6151
R3187 B.n1140 B.n74 10.6151
R3188 B.n1134 B.n74 10.6151
R3189 B.n1134 B.n1133 10.6151
R3190 B.n1133 B.n1132 10.6151
R3191 B.n1132 B.n81 10.6151
R3192 B.n1126 B.n81 10.6151
R3193 B.n1126 B.n1125 10.6151
R3194 B.n1125 B.n1124 10.6151
R3195 B.n1124 B.n88 10.6151
R3196 B.n1118 B.n88 10.6151
R3197 B.n1118 B.n1117 10.6151
R3198 B.n1117 B.n1116 10.6151
R3199 B.n1116 B.n95 10.6151
R3200 B.n1110 B.n95 10.6151
R3201 B.n1110 B.n1109 10.6151
R3202 B.n1109 B.n1108 10.6151
R3203 B.n1108 B.n102 10.6151
R3204 B.n1102 B.n102 10.6151
R3205 B.n1102 B.n1101 10.6151
R3206 B.n1101 B.n1100 10.6151
R3207 B.n176 B.n109 10.6151
R3208 B.n179 B.n176 10.6151
R3209 B.n180 B.n179 10.6151
R3210 B.n183 B.n180 10.6151
R3211 B.n184 B.n183 10.6151
R3212 B.n187 B.n184 10.6151
R3213 B.n188 B.n187 10.6151
R3214 B.n191 B.n188 10.6151
R3215 B.n192 B.n191 10.6151
R3216 B.n195 B.n192 10.6151
R3217 B.n196 B.n195 10.6151
R3218 B.n199 B.n196 10.6151
R3219 B.n200 B.n199 10.6151
R3220 B.n203 B.n200 10.6151
R3221 B.n204 B.n203 10.6151
R3222 B.n207 B.n204 10.6151
R3223 B.n208 B.n207 10.6151
R3224 B.n211 B.n208 10.6151
R3225 B.n212 B.n211 10.6151
R3226 B.n215 B.n212 10.6151
R3227 B.n216 B.n215 10.6151
R3228 B.n219 B.n216 10.6151
R3229 B.n220 B.n219 10.6151
R3230 B.n223 B.n220 10.6151
R3231 B.n224 B.n223 10.6151
R3232 B.n227 B.n224 10.6151
R3233 B.n228 B.n227 10.6151
R3234 B.n231 B.n228 10.6151
R3235 B.n232 B.n231 10.6151
R3236 B.n235 B.n232 10.6151
R3237 B.n236 B.n235 10.6151
R3238 B.n239 B.n236 10.6151
R3239 B.n240 B.n239 10.6151
R3240 B.n243 B.n240 10.6151
R3241 B.n244 B.n243 10.6151
R3242 B.n247 B.n244 10.6151
R3243 B.n248 B.n247 10.6151
R3244 B.n251 B.n248 10.6151
R3245 B.n252 B.n251 10.6151
R3246 B.n255 B.n252 10.6151
R3247 B.n256 B.n255 10.6151
R3248 B.n259 B.n256 10.6151
R3249 B.n260 B.n259 10.6151
R3250 B.n263 B.n260 10.6151
R3251 B.n264 B.n263 10.6151
R3252 B.n267 B.n264 10.6151
R3253 B.n268 B.n267 10.6151
R3254 B.n271 B.n268 10.6151
R3255 B.n272 B.n271 10.6151
R3256 B.n275 B.n272 10.6151
R3257 B.n276 B.n275 10.6151
R3258 B.n279 B.n276 10.6151
R3259 B.n280 B.n279 10.6151
R3260 B.n283 B.n280 10.6151
R3261 B.n288 B.n285 10.6151
R3262 B.n289 B.n288 10.6151
R3263 B.n292 B.n289 10.6151
R3264 B.n293 B.n292 10.6151
R3265 B.n296 B.n293 10.6151
R3266 B.n297 B.n296 10.6151
R3267 B.n300 B.n297 10.6151
R3268 B.n301 B.n300 10.6151
R3269 B.n304 B.n301 10.6151
R3270 B.n309 B.n306 10.6151
R3271 B.n310 B.n309 10.6151
R3272 B.n313 B.n310 10.6151
R3273 B.n314 B.n313 10.6151
R3274 B.n317 B.n314 10.6151
R3275 B.n318 B.n317 10.6151
R3276 B.n321 B.n318 10.6151
R3277 B.n322 B.n321 10.6151
R3278 B.n325 B.n322 10.6151
R3279 B.n326 B.n325 10.6151
R3280 B.n329 B.n326 10.6151
R3281 B.n330 B.n329 10.6151
R3282 B.n333 B.n330 10.6151
R3283 B.n334 B.n333 10.6151
R3284 B.n337 B.n334 10.6151
R3285 B.n338 B.n337 10.6151
R3286 B.n341 B.n338 10.6151
R3287 B.n342 B.n341 10.6151
R3288 B.n345 B.n342 10.6151
R3289 B.n346 B.n345 10.6151
R3290 B.n349 B.n346 10.6151
R3291 B.n350 B.n349 10.6151
R3292 B.n353 B.n350 10.6151
R3293 B.n354 B.n353 10.6151
R3294 B.n357 B.n354 10.6151
R3295 B.n358 B.n357 10.6151
R3296 B.n361 B.n358 10.6151
R3297 B.n362 B.n361 10.6151
R3298 B.n365 B.n362 10.6151
R3299 B.n366 B.n365 10.6151
R3300 B.n369 B.n366 10.6151
R3301 B.n370 B.n369 10.6151
R3302 B.n373 B.n370 10.6151
R3303 B.n374 B.n373 10.6151
R3304 B.n377 B.n374 10.6151
R3305 B.n378 B.n377 10.6151
R3306 B.n381 B.n378 10.6151
R3307 B.n382 B.n381 10.6151
R3308 B.n385 B.n382 10.6151
R3309 B.n386 B.n385 10.6151
R3310 B.n389 B.n386 10.6151
R3311 B.n390 B.n389 10.6151
R3312 B.n393 B.n390 10.6151
R3313 B.n394 B.n393 10.6151
R3314 B.n397 B.n394 10.6151
R3315 B.n398 B.n397 10.6151
R3316 B.n401 B.n398 10.6151
R3317 B.n402 B.n401 10.6151
R3318 B.n405 B.n402 10.6151
R3319 B.n406 B.n405 10.6151
R3320 B.n409 B.n406 10.6151
R3321 B.n411 B.n409 10.6151
R3322 B.n412 B.n411 10.6151
R3323 B.n1094 B.n412 10.6151
R3324 B.t8 B.n510 10.0301
R3325 B.t12 B.n93 10.0301
R3326 B.n704 B.n703 9.36635
R3327 B.n727 B.n561 9.36635
R3328 B.n284 B.n283 9.36635
R3329 B.n306 B.n305 9.36635
R3330 B.n1222 B.n0 8.11757
R3331 B.n1222 B.n1 8.11757
R3332 B.n446 B.t21 8.02421
R3333 B.t2 B.n1185 8.02421
R3334 B.t4 B.n462 7.02124
R3335 B.t0 B.n51 7.02124
R3336 B.n705 B.n704 1.24928
R3337 B.n562 B.n561 1.24928
R3338 B.n285 B.n284 1.24928
R3339 B.n305 B.n304 1.24928
R3340 VP.n24 VP.n23 161.3
R3341 VP.n25 VP.n20 161.3
R3342 VP.n27 VP.n26 161.3
R3343 VP.n28 VP.n19 161.3
R3344 VP.n30 VP.n29 161.3
R3345 VP.n31 VP.n18 161.3
R3346 VP.n33 VP.n32 161.3
R3347 VP.n35 VP.n34 161.3
R3348 VP.n36 VP.n16 161.3
R3349 VP.n38 VP.n37 161.3
R3350 VP.n39 VP.n15 161.3
R3351 VP.n41 VP.n40 161.3
R3352 VP.n42 VP.n14 161.3
R3353 VP.n44 VP.n43 161.3
R3354 VP.n79 VP.n78 161.3
R3355 VP.n77 VP.n1 161.3
R3356 VP.n76 VP.n75 161.3
R3357 VP.n74 VP.n2 161.3
R3358 VP.n73 VP.n72 161.3
R3359 VP.n71 VP.n3 161.3
R3360 VP.n70 VP.n69 161.3
R3361 VP.n68 VP.n67 161.3
R3362 VP.n66 VP.n5 161.3
R3363 VP.n65 VP.n64 161.3
R3364 VP.n63 VP.n6 161.3
R3365 VP.n62 VP.n61 161.3
R3366 VP.n60 VP.n7 161.3
R3367 VP.n59 VP.n58 161.3
R3368 VP.n57 VP.n56 161.3
R3369 VP.n55 VP.n9 161.3
R3370 VP.n54 VP.n53 161.3
R3371 VP.n52 VP.n10 161.3
R3372 VP.n51 VP.n50 161.3
R3373 VP.n49 VP.n11 161.3
R3374 VP.n48 VP.n47 161.3
R3375 VP.n22 VP.t1 157.864
R3376 VP.n12 VP.t5 124.692
R3377 VP.n8 VP.t4 124.692
R3378 VP.n4 VP.t6 124.692
R3379 VP.n0 VP.t3 124.692
R3380 VP.n13 VP.t0 124.692
R3381 VP.n17 VP.t2 124.692
R3382 VP.n21 VP.t7 124.692
R3383 VP.n46 VP.n12 74.2609
R3384 VP.n80 VP.n0 74.2609
R3385 VP.n45 VP.n13 74.2609
R3386 VP.n22 VP.n21 60.9336
R3387 VP.n46 VP.n45 57.4389
R3388 VP.n50 VP.n10 45.4209
R3389 VP.n76 VP.n2 45.4209
R3390 VP.n41 VP.n15 45.4209
R3391 VP.n61 VP.n6 40.577
R3392 VP.n65 VP.n6 40.577
R3393 VP.n30 VP.n19 40.577
R3394 VP.n26 VP.n19 40.577
R3395 VP.n54 VP.n10 35.7332
R3396 VP.n72 VP.n2 35.7332
R3397 VP.n37 VP.n15 35.7332
R3398 VP.n49 VP.n48 24.5923
R3399 VP.n50 VP.n49 24.5923
R3400 VP.n55 VP.n54 24.5923
R3401 VP.n56 VP.n55 24.5923
R3402 VP.n60 VP.n59 24.5923
R3403 VP.n61 VP.n60 24.5923
R3404 VP.n66 VP.n65 24.5923
R3405 VP.n67 VP.n66 24.5923
R3406 VP.n71 VP.n70 24.5923
R3407 VP.n72 VP.n71 24.5923
R3408 VP.n77 VP.n76 24.5923
R3409 VP.n78 VP.n77 24.5923
R3410 VP.n42 VP.n41 24.5923
R3411 VP.n43 VP.n42 24.5923
R3412 VP.n31 VP.n30 24.5923
R3413 VP.n32 VP.n31 24.5923
R3414 VP.n36 VP.n35 24.5923
R3415 VP.n37 VP.n36 24.5923
R3416 VP.n25 VP.n24 24.5923
R3417 VP.n26 VP.n25 24.5923
R3418 VP.n48 VP.n12 15.9852
R3419 VP.n78 VP.n0 15.9852
R3420 VP.n43 VP.n13 15.9852
R3421 VP.n59 VP.n8 13.526
R3422 VP.n67 VP.n4 13.526
R3423 VP.n32 VP.n17 13.526
R3424 VP.n24 VP.n21 13.526
R3425 VP.n56 VP.n8 11.0668
R3426 VP.n70 VP.n4 11.0668
R3427 VP.n35 VP.n17 11.0668
R3428 VP.n23 VP.n22 4.08481
R3429 VP.n45 VP.n44 0.354861
R3430 VP.n47 VP.n46 0.354861
R3431 VP.n80 VP.n79 0.354861
R3432 VP VP.n80 0.267071
R3433 VP.n23 VP.n20 0.189894
R3434 VP.n27 VP.n20 0.189894
R3435 VP.n28 VP.n27 0.189894
R3436 VP.n29 VP.n28 0.189894
R3437 VP.n29 VP.n18 0.189894
R3438 VP.n33 VP.n18 0.189894
R3439 VP.n34 VP.n33 0.189894
R3440 VP.n34 VP.n16 0.189894
R3441 VP.n38 VP.n16 0.189894
R3442 VP.n39 VP.n38 0.189894
R3443 VP.n40 VP.n39 0.189894
R3444 VP.n40 VP.n14 0.189894
R3445 VP.n44 VP.n14 0.189894
R3446 VP.n47 VP.n11 0.189894
R3447 VP.n51 VP.n11 0.189894
R3448 VP.n52 VP.n51 0.189894
R3449 VP.n53 VP.n52 0.189894
R3450 VP.n53 VP.n9 0.189894
R3451 VP.n57 VP.n9 0.189894
R3452 VP.n58 VP.n57 0.189894
R3453 VP.n58 VP.n7 0.189894
R3454 VP.n62 VP.n7 0.189894
R3455 VP.n63 VP.n62 0.189894
R3456 VP.n64 VP.n63 0.189894
R3457 VP.n64 VP.n5 0.189894
R3458 VP.n68 VP.n5 0.189894
R3459 VP.n69 VP.n68 0.189894
R3460 VP.n69 VP.n3 0.189894
R3461 VP.n73 VP.n3 0.189894
R3462 VP.n74 VP.n73 0.189894
R3463 VP.n75 VP.n74 0.189894
R3464 VP.n75 VP.n1 0.189894
R3465 VP.n79 VP.n1 0.189894
R3466 VDD1 VDD1.n0 65.8424
R3467 VDD1.n3 VDD1.n2 65.7287
R3468 VDD1.n3 VDD1.n1 65.7287
R3469 VDD1.n5 VDD1.n4 64.2529
R3470 VDD1.n5 VDD1.n3 52.4319
R3471 VDD1 VDD1.n5 1.47248
R3472 VDD1.n4 VDD1.t5 1.18898
R3473 VDD1.n4 VDD1.t7 1.18898
R3474 VDD1.n0 VDD1.t6 1.18898
R3475 VDD1.n0 VDD1.t0 1.18898
R3476 VDD1.n2 VDD1.t1 1.18898
R3477 VDD1.n2 VDD1.t4 1.18898
R3478 VDD1.n1 VDD1.t2 1.18898
R3479 VDD1.n1 VDD1.t3 1.18898
C0 VP VN 9.27851f
C1 VDD2 VTAIL 9.746039f
C2 VDD2 VDD1 2.09833f
C3 VTAIL VDD1 9.68747f
C4 VDD2 VP 0.585682f
C5 VDD2 VN 12.3658f
C6 VP VTAIL 12.768099f
C7 VP VDD1 12.7969f
C8 VN VTAIL 12.754001f
C9 VN VDD1 0.152886f
C10 VDD2 B 6.35346f
C11 VDD1 B 6.856782f
C12 VTAIL B 13.71251f
C13 VN B 18.26633f
C14 VP B 16.844118f
C15 VDD1.t6 B 0.352225f
C16 VDD1.t0 B 0.352225f
C17 VDD1.n0 B 3.22546f
C18 VDD1.t2 B 0.352225f
C19 VDD1.t3 B 0.352225f
C20 VDD1.n1 B 3.2242f
C21 VDD1.t1 B 0.352225f
C22 VDD1.t4 B 0.352225f
C23 VDD1.n2 B 3.2242f
C24 VDD1.n3 B 4.24197f
C25 VDD1.t5 B 0.352225f
C26 VDD1.t7 B 0.352225f
C27 VDD1.n4 B 3.21049f
C28 VDD1.n5 B 3.78643f
C29 VP.t3 B 2.761f
C30 VP.n0 B 1.02938f
C31 VP.n1 B 0.01874f
C32 VP.n2 B 0.015742f
C33 VP.n3 B 0.01874f
C34 VP.t6 B 2.761f
C35 VP.n4 B 0.95628f
C36 VP.n5 B 0.01874f
C37 VP.n6 B 0.015136f
C38 VP.n7 B 0.01874f
C39 VP.t4 B 2.761f
C40 VP.n8 B 0.95628f
C41 VP.n9 B 0.01874f
C42 VP.n10 B 0.015742f
C43 VP.n11 B 0.01874f
C44 VP.t5 B 2.761f
C45 VP.n12 B 1.02938f
C46 VP.t0 B 2.761f
C47 VP.n13 B 1.02938f
C48 VP.n14 B 0.01874f
C49 VP.n15 B 0.015742f
C50 VP.n16 B 0.01874f
C51 VP.t2 B 2.761f
C52 VP.n17 B 0.95628f
C53 VP.n18 B 0.01874f
C54 VP.n19 B 0.015136f
C55 VP.n20 B 0.01874f
C56 VP.t7 B 2.761f
C57 VP.n21 B 1.01852f
C58 VP.t1 B 2.98973f
C59 VP.n22 B 0.976461f
C60 VP.n23 B 0.217871f
C61 VP.n24 B 0.027032f
C62 VP.n25 B 0.034752f
C63 VP.n26 B 0.03705f
C64 VP.n27 B 0.01874f
C65 VP.n28 B 0.01874f
C66 VP.n29 B 0.01874f
C67 VP.n30 B 0.03705f
C68 VP.n31 B 0.034752f
C69 VP.n32 B 0.027032f
C70 VP.n33 B 0.01874f
C71 VP.n34 B 0.01874f
C72 VP.n35 B 0.025316f
C73 VP.n36 B 0.034752f
C74 VP.n37 B 0.03764f
C75 VP.n38 B 0.01874f
C76 VP.n39 B 0.01874f
C77 VP.n40 B 0.01874f
C78 VP.n41 B 0.035853f
C79 VP.n42 B 0.034752f
C80 VP.n43 B 0.028747f
C81 VP.n44 B 0.030241f
C82 VP.n45 B 1.29214f
C83 VP.n46 B 1.3039f
C84 VP.n47 B 0.030241f
C85 VP.n48 B 0.028747f
C86 VP.n49 B 0.034752f
C87 VP.n50 B 0.035853f
C88 VP.n51 B 0.01874f
C89 VP.n52 B 0.01874f
C90 VP.n53 B 0.01874f
C91 VP.n54 B 0.03764f
C92 VP.n55 B 0.034752f
C93 VP.n56 B 0.025316f
C94 VP.n57 B 0.01874f
C95 VP.n58 B 0.01874f
C96 VP.n59 B 0.027032f
C97 VP.n60 B 0.034752f
C98 VP.n61 B 0.03705f
C99 VP.n62 B 0.01874f
C100 VP.n63 B 0.01874f
C101 VP.n64 B 0.01874f
C102 VP.n65 B 0.03705f
C103 VP.n66 B 0.034752f
C104 VP.n67 B 0.027032f
C105 VP.n68 B 0.01874f
C106 VP.n69 B 0.01874f
C107 VP.n70 B 0.025316f
C108 VP.n71 B 0.034752f
C109 VP.n72 B 0.03764f
C110 VP.n73 B 0.01874f
C111 VP.n74 B 0.01874f
C112 VP.n75 B 0.01874f
C113 VP.n76 B 0.035853f
C114 VP.n77 B 0.034752f
C115 VP.n78 B 0.028747f
C116 VP.n79 B 0.030241f
C117 VP.n80 B 0.043771f
C118 VDD2.t6 B 0.347895f
C119 VDD2.t4 B 0.347895f
C120 VDD2.n0 B 3.18457f
C121 VDD2.t1 B 0.347895f
C122 VDD2.t0 B 0.347895f
C123 VDD2.n1 B 3.18457f
C124 VDD2.n2 B 4.13532f
C125 VDD2.t3 B 0.347895f
C126 VDD2.t7 B 0.347895f
C127 VDD2.n3 B 3.17103f
C128 VDD2.n4 B 3.70669f
C129 VDD2.t5 B 0.347895f
C130 VDD2.t2 B 0.347895f
C131 VDD2.n5 B 3.18453f
C132 VTAIL.t7 B 0.251806f
C133 VTAIL.t11 B 0.251806f
C134 VTAIL.n0 B 2.24407f
C135 VTAIL.n1 B 0.366779f
C136 VTAIL.n2 B 0.010792f
C137 VTAIL.n3 B 0.024293f
C138 VTAIL.n4 B 0.010882f
C139 VTAIL.n5 B 0.019127f
C140 VTAIL.n6 B 0.010278f
C141 VTAIL.n7 B 0.024293f
C142 VTAIL.n8 B 0.010882f
C143 VTAIL.n9 B 0.019127f
C144 VTAIL.n10 B 0.010278f
C145 VTAIL.n11 B 0.024293f
C146 VTAIL.n12 B 0.010882f
C147 VTAIL.n13 B 0.019127f
C148 VTAIL.n14 B 0.010278f
C149 VTAIL.n15 B 0.024293f
C150 VTAIL.n16 B 0.010882f
C151 VTAIL.n17 B 0.019127f
C152 VTAIL.n18 B 0.010278f
C153 VTAIL.n19 B 0.024293f
C154 VTAIL.n20 B 0.01058f
C155 VTAIL.n21 B 0.019127f
C156 VTAIL.n22 B 0.010882f
C157 VTAIL.n23 B 0.024293f
C158 VTAIL.n24 B 0.010882f
C159 VTAIL.n25 B 0.019127f
C160 VTAIL.n26 B 0.010278f
C161 VTAIL.n27 B 0.024293f
C162 VTAIL.n28 B 0.010882f
C163 VTAIL.n29 B 1.36134f
C164 VTAIL.n30 B 0.010278f
C165 VTAIL.t14 B 0.041509f
C166 VTAIL.n31 B 0.172119f
C167 VTAIL.n32 B 0.017173f
C168 VTAIL.n33 B 0.01822f
C169 VTAIL.n34 B 0.024293f
C170 VTAIL.n35 B 0.010882f
C171 VTAIL.n36 B 0.010278f
C172 VTAIL.n37 B 0.019127f
C173 VTAIL.n38 B 0.019127f
C174 VTAIL.n39 B 0.010278f
C175 VTAIL.n40 B 0.010882f
C176 VTAIL.n41 B 0.024293f
C177 VTAIL.n42 B 0.024293f
C178 VTAIL.n43 B 0.010882f
C179 VTAIL.n44 B 0.010278f
C180 VTAIL.n45 B 0.019127f
C181 VTAIL.n46 B 0.019127f
C182 VTAIL.n47 B 0.010278f
C183 VTAIL.n48 B 0.010278f
C184 VTAIL.n49 B 0.010882f
C185 VTAIL.n50 B 0.024293f
C186 VTAIL.n51 B 0.024293f
C187 VTAIL.n52 B 0.024293f
C188 VTAIL.n53 B 0.01058f
C189 VTAIL.n54 B 0.010278f
C190 VTAIL.n55 B 0.019127f
C191 VTAIL.n56 B 0.019127f
C192 VTAIL.n57 B 0.010278f
C193 VTAIL.n58 B 0.010882f
C194 VTAIL.n59 B 0.024293f
C195 VTAIL.n60 B 0.024293f
C196 VTAIL.n61 B 0.010882f
C197 VTAIL.n62 B 0.010278f
C198 VTAIL.n63 B 0.019127f
C199 VTAIL.n64 B 0.019127f
C200 VTAIL.n65 B 0.010278f
C201 VTAIL.n66 B 0.010882f
C202 VTAIL.n67 B 0.024293f
C203 VTAIL.n68 B 0.024293f
C204 VTAIL.n69 B 0.010882f
C205 VTAIL.n70 B 0.010278f
C206 VTAIL.n71 B 0.019127f
C207 VTAIL.n72 B 0.019127f
C208 VTAIL.n73 B 0.010278f
C209 VTAIL.n74 B 0.010882f
C210 VTAIL.n75 B 0.024293f
C211 VTAIL.n76 B 0.024293f
C212 VTAIL.n77 B 0.010882f
C213 VTAIL.n78 B 0.010278f
C214 VTAIL.n79 B 0.019127f
C215 VTAIL.n80 B 0.019127f
C216 VTAIL.n81 B 0.010278f
C217 VTAIL.n82 B 0.010882f
C218 VTAIL.n83 B 0.024293f
C219 VTAIL.n84 B 0.024293f
C220 VTAIL.n85 B 0.010882f
C221 VTAIL.n86 B 0.010278f
C222 VTAIL.n87 B 0.019127f
C223 VTAIL.n88 B 0.049959f
C224 VTAIL.n89 B 0.010278f
C225 VTAIL.n90 B 0.010882f
C226 VTAIL.n91 B 0.04757f
C227 VTAIL.n92 B 0.040989f
C228 VTAIL.n93 B 0.235082f
C229 VTAIL.n94 B 0.010792f
C230 VTAIL.n95 B 0.024293f
C231 VTAIL.n96 B 0.010882f
C232 VTAIL.n97 B 0.019127f
C233 VTAIL.n98 B 0.010278f
C234 VTAIL.n99 B 0.024293f
C235 VTAIL.n100 B 0.010882f
C236 VTAIL.n101 B 0.019127f
C237 VTAIL.n102 B 0.010278f
C238 VTAIL.n103 B 0.024293f
C239 VTAIL.n104 B 0.010882f
C240 VTAIL.n105 B 0.019127f
C241 VTAIL.n106 B 0.010278f
C242 VTAIL.n107 B 0.024293f
C243 VTAIL.n108 B 0.010882f
C244 VTAIL.n109 B 0.019127f
C245 VTAIL.n110 B 0.010278f
C246 VTAIL.n111 B 0.024293f
C247 VTAIL.n112 B 0.01058f
C248 VTAIL.n113 B 0.019127f
C249 VTAIL.n114 B 0.010882f
C250 VTAIL.n115 B 0.024293f
C251 VTAIL.n116 B 0.010882f
C252 VTAIL.n117 B 0.019127f
C253 VTAIL.n118 B 0.010278f
C254 VTAIL.n119 B 0.024293f
C255 VTAIL.n120 B 0.010882f
C256 VTAIL.n121 B 1.36134f
C257 VTAIL.n122 B 0.010278f
C258 VTAIL.t6 B 0.041509f
C259 VTAIL.n123 B 0.172119f
C260 VTAIL.n124 B 0.017173f
C261 VTAIL.n125 B 0.01822f
C262 VTAIL.n126 B 0.024293f
C263 VTAIL.n127 B 0.010882f
C264 VTAIL.n128 B 0.010278f
C265 VTAIL.n129 B 0.019127f
C266 VTAIL.n130 B 0.019127f
C267 VTAIL.n131 B 0.010278f
C268 VTAIL.n132 B 0.010882f
C269 VTAIL.n133 B 0.024293f
C270 VTAIL.n134 B 0.024293f
C271 VTAIL.n135 B 0.010882f
C272 VTAIL.n136 B 0.010278f
C273 VTAIL.n137 B 0.019127f
C274 VTAIL.n138 B 0.019127f
C275 VTAIL.n139 B 0.010278f
C276 VTAIL.n140 B 0.010278f
C277 VTAIL.n141 B 0.010882f
C278 VTAIL.n142 B 0.024293f
C279 VTAIL.n143 B 0.024293f
C280 VTAIL.n144 B 0.024293f
C281 VTAIL.n145 B 0.01058f
C282 VTAIL.n146 B 0.010278f
C283 VTAIL.n147 B 0.019127f
C284 VTAIL.n148 B 0.019127f
C285 VTAIL.n149 B 0.010278f
C286 VTAIL.n150 B 0.010882f
C287 VTAIL.n151 B 0.024293f
C288 VTAIL.n152 B 0.024293f
C289 VTAIL.n153 B 0.010882f
C290 VTAIL.n154 B 0.010278f
C291 VTAIL.n155 B 0.019127f
C292 VTAIL.n156 B 0.019127f
C293 VTAIL.n157 B 0.010278f
C294 VTAIL.n158 B 0.010882f
C295 VTAIL.n159 B 0.024293f
C296 VTAIL.n160 B 0.024293f
C297 VTAIL.n161 B 0.010882f
C298 VTAIL.n162 B 0.010278f
C299 VTAIL.n163 B 0.019127f
C300 VTAIL.n164 B 0.019127f
C301 VTAIL.n165 B 0.010278f
C302 VTAIL.n166 B 0.010882f
C303 VTAIL.n167 B 0.024293f
C304 VTAIL.n168 B 0.024293f
C305 VTAIL.n169 B 0.010882f
C306 VTAIL.n170 B 0.010278f
C307 VTAIL.n171 B 0.019127f
C308 VTAIL.n172 B 0.019127f
C309 VTAIL.n173 B 0.010278f
C310 VTAIL.n174 B 0.010882f
C311 VTAIL.n175 B 0.024293f
C312 VTAIL.n176 B 0.024293f
C313 VTAIL.n177 B 0.010882f
C314 VTAIL.n178 B 0.010278f
C315 VTAIL.n179 B 0.019127f
C316 VTAIL.n180 B 0.049959f
C317 VTAIL.n181 B 0.010278f
C318 VTAIL.n182 B 0.010882f
C319 VTAIL.n183 B 0.04757f
C320 VTAIL.n184 B 0.040989f
C321 VTAIL.n185 B 0.235082f
C322 VTAIL.t4 B 0.251806f
C323 VTAIL.t15 B 0.251806f
C324 VTAIL.n186 B 2.24407f
C325 VTAIL.n187 B 0.551802f
C326 VTAIL.n188 B 0.010792f
C327 VTAIL.n189 B 0.024293f
C328 VTAIL.n190 B 0.010882f
C329 VTAIL.n191 B 0.019127f
C330 VTAIL.n192 B 0.010278f
C331 VTAIL.n193 B 0.024293f
C332 VTAIL.n194 B 0.010882f
C333 VTAIL.n195 B 0.019127f
C334 VTAIL.n196 B 0.010278f
C335 VTAIL.n197 B 0.024293f
C336 VTAIL.n198 B 0.010882f
C337 VTAIL.n199 B 0.019127f
C338 VTAIL.n200 B 0.010278f
C339 VTAIL.n201 B 0.024293f
C340 VTAIL.n202 B 0.010882f
C341 VTAIL.n203 B 0.019127f
C342 VTAIL.n204 B 0.010278f
C343 VTAIL.n205 B 0.024293f
C344 VTAIL.n206 B 0.01058f
C345 VTAIL.n207 B 0.019127f
C346 VTAIL.n208 B 0.010882f
C347 VTAIL.n209 B 0.024293f
C348 VTAIL.n210 B 0.010882f
C349 VTAIL.n211 B 0.019127f
C350 VTAIL.n212 B 0.010278f
C351 VTAIL.n213 B 0.024293f
C352 VTAIL.n214 B 0.010882f
C353 VTAIL.n215 B 1.36134f
C354 VTAIL.n216 B 0.010278f
C355 VTAIL.t3 B 0.041509f
C356 VTAIL.n217 B 0.172119f
C357 VTAIL.n218 B 0.017173f
C358 VTAIL.n219 B 0.01822f
C359 VTAIL.n220 B 0.024293f
C360 VTAIL.n221 B 0.010882f
C361 VTAIL.n222 B 0.010278f
C362 VTAIL.n223 B 0.019127f
C363 VTAIL.n224 B 0.019127f
C364 VTAIL.n225 B 0.010278f
C365 VTAIL.n226 B 0.010882f
C366 VTAIL.n227 B 0.024293f
C367 VTAIL.n228 B 0.024293f
C368 VTAIL.n229 B 0.010882f
C369 VTAIL.n230 B 0.010278f
C370 VTAIL.n231 B 0.019127f
C371 VTAIL.n232 B 0.019127f
C372 VTAIL.n233 B 0.010278f
C373 VTAIL.n234 B 0.010278f
C374 VTAIL.n235 B 0.010882f
C375 VTAIL.n236 B 0.024293f
C376 VTAIL.n237 B 0.024293f
C377 VTAIL.n238 B 0.024293f
C378 VTAIL.n239 B 0.01058f
C379 VTAIL.n240 B 0.010278f
C380 VTAIL.n241 B 0.019127f
C381 VTAIL.n242 B 0.019127f
C382 VTAIL.n243 B 0.010278f
C383 VTAIL.n244 B 0.010882f
C384 VTAIL.n245 B 0.024293f
C385 VTAIL.n246 B 0.024293f
C386 VTAIL.n247 B 0.010882f
C387 VTAIL.n248 B 0.010278f
C388 VTAIL.n249 B 0.019127f
C389 VTAIL.n250 B 0.019127f
C390 VTAIL.n251 B 0.010278f
C391 VTAIL.n252 B 0.010882f
C392 VTAIL.n253 B 0.024293f
C393 VTAIL.n254 B 0.024293f
C394 VTAIL.n255 B 0.010882f
C395 VTAIL.n256 B 0.010278f
C396 VTAIL.n257 B 0.019127f
C397 VTAIL.n258 B 0.019127f
C398 VTAIL.n259 B 0.010278f
C399 VTAIL.n260 B 0.010882f
C400 VTAIL.n261 B 0.024293f
C401 VTAIL.n262 B 0.024293f
C402 VTAIL.n263 B 0.010882f
C403 VTAIL.n264 B 0.010278f
C404 VTAIL.n265 B 0.019127f
C405 VTAIL.n266 B 0.019127f
C406 VTAIL.n267 B 0.010278f
C407 VTAIL.n268 B 0.010882f
C408 VTAIL.n269 B 0.024293f
C409 VTAIL.n270 B 0.024293f
C410 VTAIL.n271 B 0.010882f
C411 VTAIL.n272 B 0.010278f
C412 VTAIL.n273 B 0.019127f
C413 VTAIL.n274 B 0.049959f
C414 VTAIL.n275 B 0.010278f
C415 VTAIL.n276 B 0.010882f
C416 VTAIL.n277 B 0.04757f
C417 VTAIL.n278 B 0.040989f
C418 VTAIL.n279 B 1.53969f
C419 VTAIL.n280 B 0.010792f
C420 VTAIL.n281 B 0.024293f
C421 VTAIL.n282 B 0.010882f
C422 VTAIL.n283 B 0.019127f
C423 VTAIL.n284 B 0.010278f
C424 VTAIL.n285 B 0.024293f
C425 VTAIL.n286 B 0.010882f
C426 VTAIL.n287 B 0.019127f
C427 VTAIL.n288 B 0.010278f
C428 VTAIL.n289 B 0.024293f
C429 VTAIL.n290 B 0.010882f
C430 VTAIL.n291 B 0.019127f
C431 VTAIL.n292 B 0.010278f
C432 VTAIL.n293 B 0.024293f
C433 VTAIL.n294 B 0.010882f
C434 VTAIL.n295 B 0.019127f
C435 VTAIL.n296 B 0.010278f
C436 VTAIL.n297 B 0.024293f
C437 VTAIL.n298 B 0.01058f
C438 VTAIL.n299 B 0.019127f
C439 VTAIL.n300 B 0.01058f
C440 VTAIL.n301 B 0.010278f
C441 VTAIL.n302 B 0.024293f
C442 VTAIL.n303 B 0.024293f
C443 VTAIL.n304 B 0.010882f
C444 VTAIL.n305 B 0.019127f
C445 VTAIL.n306 B 0.010278f
C446 VTAIL.n307 B 0.024293f
C447 VTAIL.n308 B 0.010882f
C448 VTAIL.n309 B 1.36134f
C449 VTAIL.n310 B 0.010278f
C450 VTAIL.t12 B 0.041509f
C451 VTAIL.n311 B 0.172119f
C452 VTAIL.n312 B 0.017173f
C453 VTAIL.n313 B 0.01822f
C454 VTAIL.n314 B 0.024293f
C455 VTAIL.n315 B 0.010882f
C456 VTAIL.n316 B 0.010278f
C457 VTAIL.n317 B 0.019127f
C458 VTAIL.n318 B 0.019127f
C459 VTAIL.n319 B 0.010278f
C460 VTAIL.n320 B 0.010882f
C461 VTAIL.n321 B 0.024293f
C462 VTAIL.n322 B 0.024293f
C463 VTAIL.n323 B 0.010882f
C464 VTAIL.n324 B 0.010278f
C465 VTAIL.n325 B 0.019127f
C466 VTAIL.n326 B 0.019127f
C467 VTAIL.n327 B 0.010278f
C468 VTAIL.n328 B 0.010882f
C469 VTAIL.n329 B 0.024293f
C470 VTAIL.n330 B 0.024293f
C471 VTAIL.n331 B 0.010882f
C472 VTAIL.n332 B 0.010278f
C473 VTAIL.n333 B 0.019127f
C474 VTAIL.n334 B 0.019127f
C475 VTAIL.n335 B 0.010278f
C476 VTAIL.n336 B 0.010882f
C477 VTAIL.n337 B 0.024293f
C478 VTAIL.n338 B 0.024293f
C479 VTAIL.n339 B 0.010882f
C480 VTAIL.n340 B 0.010278f
C481 VTAIL.n341 B 0.019127f
C482 VTAIL.n342 B 0.019127f
C483 VTAIL.n343 B 0.010278f
C484 VTAIL.n344 B 0.010882f
C485 VTAIL.n345 B 0.024293f
C486 VTAIL.n346 B 0.024293f
C487 VTAIL.n347 B 0.010882f
C488 VTAIL.n348 B 0.010278f
C489 VTAIL.n349 B 0.019127f
C490 VTAIL.n350 B 0.019127f
C491 VTAIL.n351 B 0.010278f
C492 VTAIL.n352 B 0.010882f
C493 VTAIL.n353 B 0.024293f
C494 VTAIL.n354 B 0.024293f
C495 VTAIL.n355 B 0.010882f
C496 VTAIL.n356 B 0.010278f
C497 VTAIL.n357 B 0.019127f
C498 VTAIL.n358 B 0.019127f
C499 VTAIL.n359 B 0.010278f
C500 VTAIL.n360 B 0.010882f
C501 VTAIL.n361 B 0.024293f
C502 VTAIL.n362 B 0.024293f
C503 VTAIL.n363 B 0.010882f
C504 VTAIL.n364 B 0.010278f
C505 VTAIL.n365 B 0.019127f
C506 VTAIL.n366 B 0.049959f
C507 VTAIL.n367 B 0.010278f
C508 VTAIL.n368 B 0.010882f
C509 VTAIL.n369 B 0.04757f
C510 VTAIL.n370 B 0.040989f
C511 VTAIL.n371 B 1.53969f
C512 VTAIL.t10 B 0.251806f
C513 VTAIL.t13 B 0.251806f
C514 VTAIL.n372 B 2.24407f
C515 VTAIL.n373 B 0.551797f
C516 VTAIL.n374 B 0.010792f
C517 VTAIL.n375 B 0.024293f
C518 VTAIL.n376 B 0.010882f
C519 VTAIL.n377 B 0.019127f
C520 VTAIL.n378 B 0.010278f
C521 VTAIL.n379 B 0.024293f
C522 VTAIL.n380 B 0.010882f
C523 VTAIL.n381 B 0.019127f
C524 VTAIL.n382 B 0.010278f
C525 VTAIL.n383 B 0.024293f
C526 VTAIL.n384 B 0.010882f
C527 VTAIL.n385 B 0.019127f
C528 VTAIL.n386 B 0.010278f
C529 VTAIL.n387 B 0.024293f
C530 VTAIL.n388 B 0.010882f
C531 VTAIL.n389 B 0.019127f
C532 VTAIL.n390 B 0.010278f
C533 VTAIL.n391 B 0.024293f
C534 VTAIL.n392 B 0.01058f
C535 VTAIL.n393 B 0.019127f
C536 VTAIL.n394 B 0.01058f
C537 VTAIL.n395 B 0.010278f
C538 VTAIL.n396 B 0.024293f
C539 VTAIL.n397 B 0.024293f
C540 VTAIL.n398 B 0.010882f
C541 VTAIL.n399 B 0.019127f
C542 VTAIL.n400 B 0.010278f
C543 VTAIL.n401 B 0.024293f
C544 VTAIL.n402 B 0.010882f
C545 VTAIL.n403 B 1.36134f
C546 VTAIL.n404 B 0.010278f
C547 VTAIL.t9 B 0.041509f
C548 VTAIL.n405 B 0.172119f
C549 VTAIL.n406 B 0.017173f
C550 VTAIL.n407 B 0.01822f
C551 VTAIL.n408 B 0.024293f
C552 VTAIL.n409 B 0.010882f
C553 VTAIL.n410 B 0.010278f
C554 VTAIL.n411 B 0.019127f
C555 VTAIL.n412 B 0.019127f
C556 VTAIL.n413 B 0.010278f
C557 VTAIL.n414 B 0.010882f
C558 VTAIL.n415 B 0.024293f
C559 VTAIL.n416 B 0.024293f
C560 VTAIL.n417 B 0.010882f
C561 VTAIL.n418 B 0.010278f
C562 VTAIL.n419 B 0.019127f
C563 VTAIL.n420 B 0.019127f
C564 VTAIL.n421 B 0.010278f
C565 VTAIL.n422 B 0.010882f
C566 VTAIL.n423 B 0.024293f
C567 VTAIL.n424 B 0.024293f
C568 VTAIL.n425 B 0.010882f
C569 VTAIL.n426 B 0.010278f
C570 VTAIL.n427 B 0.019127f
C571 VTAIL.n428 B 0.019127f
C572 VTAIL.n429 B 0.010278f
C573 VTAIL.n430 B 0.010882f
C574 VTAIL.n431 B 0.024293f
C575 VTAIL.n432 B 0.024293f
C576 VTAIL.n433 B 0.010882f
C577 VTAIL.n434 B 0.010278f
C578 VTAIL.n435 B 0.019127f
C579 VTAIL.n436 B 0.019127f
C580 VTAIL.n437 B 0.010278f
C581 VTAIL.n438 B 0.010882f
C582 VTAIL.n439 B 0.024293f
C583 VTAIL.n440 B 0.024293f
C584 VTAIL.n441 B 0.010882f
C585 VTAIL.n442 B 0.010278f
C586 VTAIL.n443 B 0.019127f
C587 VTAIL.n444 B 0.019127f
C588 VTAIL.n445 B 0.010278f
C589 VTAIL.n446 B 0.010882f
C590 VTAIL.n447 B 0.024293f
C591 VTAIL.n448 B 0.024293f
C592 VTAIL.n449 B 0.010882f
C593 VTAIL.n450 B 0.010278f
C594 VTAIL.n451 B 0.019127f
C595 VTAIL.n452 B 0.019127f
C596 VTAIL.n453 B 0.010278f
C597 VTAIL.n454 B 0.010882f
C598 VTAIL.n455 B 0.024293f
C599 VTAIL.n456 B 0.024293f
C600 VTAIL.n457 B 0.010882f
C601 VTAIL.n458 B 0.010278f
C602 VTAIL.n459 B 0.019127f
C603 VTAIL.n460 B 0.049959f
C604 VTAIL.n461 B 0.010278f
C605 VTAIL.n462 B 0.010882f
C606 VTAIL.n463 B 0.04757f
C607 VTAIL.n464 B 0.040989f
C608 VTAIL.n465 B 0.235082f
C609 VTAIL.n466 B 0.010792f
C610 VTAIL.n467 B 0.024293f
C611 VTAIL.n468 B 0.010882f
C612 VTAIL.n469 B 0.019127f
C613 VTAIL.n470 B 0.010278f
C614 VTAIL.n471 B 0.024293f
C615 VTAIL.n472 B 0.010882f
C616 VTAIL.n473 B 0.019127f
C617 VTAIL.n474 B 0.010278f
C618 VTAIL.n475 B 0.024293f
C619 VTAIL.n476 B 0.010882f
C620 VTAIL.n477 B 0.019127f
C621 VTAIL.n478 B 0.010278f
C622 VTAIL.n479 B 0.024293f
C623 VTAIL.n480 B 0.010882f
C624 VTAIL.n481 B 0.019127f
C625 VTAIL.n482 B 0.010278f
C626 VTAIL.n483 B 0.024293f
C627 VTAIL.n484 B 0.01058f
C628 VTAIL.n485 B 0.019127f
C629 VTAIL.n486 B 0.01058f
C630 VTAIL.n487 B 0.010278f
C631 VTAIL.n488 B 0.024293f
C632 VTAIL.n489 B 0.024293f
C633 VTAIL.n490 B 0.010882f
C634 VTAIL.n491 B 0.019127f
C635 VTAIL.n492 B 0.010278f
C636 VTAIL.n493 B 0.024293f
C637 VTAIL.n494 B 0.010882f
C638 VTAIL.n495 B 1.36134f
C639 VTAIL.n496 B 0.010278f
C640 VTAIL.t5 B 0.041509f
C641 VTAIL.n497 B 0.172119f
C642 VTAIL.n498 B 0.017173f
C643 VTAIL.n499 B 0.01822f
C644 VTAIL.n500 B 0.024293f
C645 VTAIL.n501 B 0.010882f
C646 VTAIL.n502 B 0.010278f
C647 VTAIL.n503 B 0.019127f
C648 VTAIL.n504 B 0.019127f
C649 VTAIL.n505 B 0.010278f
C650 VTAIL.n506 B 0.010882f
C651 VTAIL.n507 B 0.024293f
C652 VTAIL.n508 B 0.024293f
C653 VTAIL.n509 B 0.010882f
C654 VTAIL.n510 B 0.010278f
C655 VTAIL.n511 B 0.019127f
C656 VTAIL.n512 B 0.019127f
C657 VTAIL.n513 B 0.010278f
C658 VTAIL.n514 B 0.010882f
C659 VTAIL.n515 B 0.024293f
C660 VTAIL.n516 B 0.024293f
C661 VTAIL.n517 B 0.010882f
C662 VTAIL.n518 B 0.010278f
C663 VTAIL.n519 B 0.019127f
C664 VTAIL.n520 B 0.019127f
C665 VTAIL.n521 B 0.010278f
C666 VTAIL.n522 B 0.010882f
C667 VTAIL.n523 B 0.024293f
C668 VTAIL.n524 B 0.024293f
C669 VTAIL.n525 B 0.010882f
C670 VTAIL.n526 B 0.010278f
C671 VTAIL.n527 B 0.019127f
C672 VTAIL.n528 B 0.019127f
C673 VTAIL.n529 B 0.010278f
C674 VTAIL.n530 B 0.010882f
C675 VTAIL.n531 B 0.024293f
C676 VTAIL.n532 B 0.024293f
C677 VTAIL.n533 B 0.010882f
C678 VTAIL.n534 B 0.010278f
C679 VTAIL.n535 B 0.019127f
C680 VTAIL.n536 B 0.019127f
C681 VTAIL.n537 B 0.010278f
C682 VTAIL.n538 B 0.010882f
C683 VTAIL.n539 B 0.024293f
C684 VTAIL.n540 B 0.024293f
C685 VTAIL.n541 B 0.010882f
C686 VTAIL.n542 B 0.010278f
C687 VTAIL.n543 B 0.019127f
C688 VTAIL.n544 B 0.019127f
C689 VTAIL.n545 B 0.010278f
C690 VTAIL.n546 B 0.010882f
C691 VTAIL.n547 B 0.024293f
C692 VTAIL.n548 B 0.024293f
C693 VTAIL.n549 B 0.010882f
C694 VTAIL.n550 B 0.010278f
C695 VTAIL.n551 B 0.019127f
C696 VTAIL.n552 B 0.049959f
C697 VTAIL.n553 B 0.010278f
C698 VTAIL.n554 B 0.010882f
C699 VTAIL.n555 B 0.04757f
C700 VTAIL.n556 B 0.040989f
C701 VTAIL.n557 B 0.235082f
C702 VTAIL.t2 B 0.251806f
C703 VTAIL.t0 B 0.251806f
C704 VTAIL.n558 B 2.24407f
C705 VTAIL.n559 B 0.551797f
C706 VTAIL.n560 B 0.010792f
C707 VTAIL.n561 B 0.024293f
C708 VTAIL.n562 B 0.010882f
C709 VTAIL.n563 B 0.019127f
C710 VTAIL.n564 B 0.010278f
C711 VTAIL.n565 B 0.024293f
C712 VTAIL.n566 B 0.010882f
C713 VTAIL.n567 B 0.019127f
C714 VTAIL.n568 B 0.010278f
C715 VTAIL.n569 B 0.024293f
C716 VTAIL.n570 B 0.010882f
C717 VTAIL.n571 B 0.019127f
C718 VTAIL.n572 B 0.010278f
C719 VTAIL.n573 B 0.024293f
C720 VTAIL.n574 B 0.010882f
C721 VTAIL.n575 B 0.019127f
C722 VTAIL.n576 B 0.010278f
C723 VTAIL.n577 B 0.024293f
C724 VTAIL.n578 B 0.01058f
C725 VTAIL.n579 B 0.019127f
C726 VTAIL.n580 B 0.01058f
C727 VTAIL.n581 B 0.010278f
C728 VTAIL.n582 B 0.024293f
C729 VTAIL.n583 B 0.024293f
C730 VTAIL.n584 B 0.010882f
C731 VTAIL.n585 B 0.019127f
C732 VTAIL.n586 B 0.010278f
C733 VTAIL.n587 B 0.024293f
C734 VTAIL.n588 B 0.010882f
C735 VTAIL.n589 B 1.36134f
C736 VTAIL.n590 B 0.010278f
C737 VTAIL.t1 B 0.041509f
C738 VTAIL.n591 B 0.172119f
C739 VTAIL.n592 B 0.017173f
C740 VTAIL.n593 B 0.01822f
C741 VTAIL.n594 B 0.024293f
C742 VTAIL.n595 B 0.010882f
C743 VTAIL.n596 B 0.010278f
C744 VTAIL.n597 B 0.019127f
C745 VTAIL.n598 B 0.019127f
C746 VTAIL.n599 B 0.010278f
C747 VTAIL.n600 B 0.010882f
C748 VTAIL.n601 B 0.024293f
C749 VTAIL.n602 B 0.024293f
C750 VTAIL.n603 B 0.010882f
C751 VTAIL.n604 B 0.010278f
C752 VTAIL.n605 B 0.019127f
C753 VTAIL.n606 B 0.019127f
C754 VTAIL.n607 B 0.010278f
C755 VTAIL.n608 B 0.010882f
C756 VTAIL.n609 B 0.024293f
C757 VTAIL.n610 B 0.024293f
C758 VTAIL.n611 B 0.010882f
C759 VTAIL.n612 B 0.010278f
C760 VTAIL.n613 B 0.019127f
C761 VTAIL.n614 B 0.019127f
C762 VTAIL.n615 B 0.010278f
C763 VTAIL.n616 B 0.010882f
C764 VTAIL.n617 B 0.024293f
C765 VTAIL.n618 B 0.024293f
C766 VTAIL.n619 B 0.010882f
C767 VTAIL.n620 B 0.010278f
C768 VTAIL.n621 B 0.019127f
C769 VTAIL.n622 B 0.019127f
C770 VTAIL.n623 B 0.010278f
C771 VTAIL.n624 B 0.010882f
C772 VTAIL.n625 B 0.024293f
C773 VTAIL.n626 B 0.024293f
C774 VTAIL.n627 B 0.010882f
C775 VTAIL.n628 B 0.010278f
C776 VTAIL.n629 B 0.019127f
C777 VTAIL.n630 B 0.019127f
C778 VTAIL.n631 B 0.010278f
C779 VTAIL.n632 B 0.010882f
C780 VTAIL.n633 B 0.024293f
C781 VTAIL.n634 B 0.024293f
C782 VTAIL.n635 B 0.010882f
C783 VTAIL.n636 B 0.010278f
C784 VTAIL.n637 B 0.019127f
C785 VTAIL.n638 B 0.019127f
C786 VTAIL.n639 B 0.010278f
C787 VTAIL.n640 B 0.010882f
C788 VTAIL.n641 B 0.024293f
C789 VTAIL.n642 B 0.024293f
C790 VTAIL.n643 B 0.010882f
C791 VTAIL.n644 B 0.010278f
C792 VTAIL.n645 B 0.019127f
C793 VTAIL.n646 B 0.049959f
C794 VTAIL.n647 B 0.010278f
C795 VTAIL.n648 B 0.010882f
C796 VTAIL.n649 B 0.04757f
C797 VTAIL.n650 B 0.040989f
C798 VTAIL.n651 B 1.53969f
C799 VTAIL.n652 B 0.010792f
C800 VTAIL.n653 B 0.024293f
C801 VTAIL.n654 B 0.010882f
C802 VTAIL.n655 B 0.019127f
C803 VTAIL.n656 B 0.010278f
C804 VTAIL.n657 B 0.024293f
C805 VTAIL.n658 B 0.010882f
C806 VTAIL.n659 B 0.019127f
C807 VTAIL.n660 B 0.010278f
C808 VTAIL.n661 B 0.024293f
C809 VTAIL.n662 B 0.010882f
C810 VTAIL.n663 B 0.019127f
C811 VTAIL.n664 B 0.010278f
C812 VTAIL.n665 B 0.024293f
C813 VTAIL.n666 B 0.010882f
C814 VTAIL.n667 B 0.019127f
C815 VTAIL.n668 B 0.010278f
C816 VTAIL.n669 B 0.024293f
C817 VTAIL.n670 B 0.01058f
C818 VTAIL.n671 B 0.019127f
C819 VTAIL.n672 B 0.010882f
C820 VTAIL.n673 B 0.024293f
C821 VTAIL.n674 B 0.010882f
C822 VTAIL.n675 B 0.019127f
C823 VTAIL.n676 B 0.010278f
C824 VTAIL.n677 B 0.024293f
C825 VTAIL.n678 B 0.010882f
C826 VTAIL.n679 B 1.36134f
C827 VTAIL.n680 B 0.010278f
C828 VTAIL.t8 B 0.041509f
C829 VTAIL.n681 B 0.172119f
C830 VTAIL.n682 B 0.017173f
C831 VTAIL.n683 B 0.01822f
C832 VTAIL.n684 B 0.024293f
C833 VTAIL.n685 B 0.010882f
C834 VTAIL.n686 B 0.010278f
C835 VTAIL.n687 B 0.019127f
C836 VTAIL.n688 B 0.019127f
C837 VTAIL.n689 B 0.010278f
C838 VTAIL.n690 B 0.010882f
C839 VTAIL.n691 B 0.024293f
C840 VTAIL.n692 B 0.024293f
C841 VTAIL.n693 B 0.010882f
C842 VTAIL.n694 B 0.010278f
C843 VTAIL.n695 B 0.019127f
C844 VTAIL.n696 B 0.019127f
C845 VTAIL.n697 B 0.010278f
C846 VTAIL.n698 B 0.010278f
C847 VTAIL.n699 B 0.010882f
C848 VTAIL.n700 B 0.024293f
C849 VTAIL.n701 B 0.024293f
C850 VTAIL.n702 B 0.024293f
C851 VTAIL.n703 B 0.01058f
C852 VTAIL.n704 B 0.010278f
C853 VTAIL.n705 B 0.019127f
C854 VTAIL.n706 B 0.019127f
C855 VTAIL.n707 B 0.010278f
C856 VTAIL.n708 B 0.010882f
C857 VTAIL.n709 B 0.024293f
C858 VTAIL.n710 B 0.024293f
C859 VTAIL.n711 B 0.010882f
C860 VTAIL.n712 B 0.010278f
C861 VTAIL.n713 B 0.019127f
C862 VTAIL.n714 B 0.019127f
C863 VTAIL.n715 B 0.010278f
C864 VTAIL.n716 B 0.010882f
C865 VTAIL.n717 B 0.024293f
C866 VTAIL.n718 B 0.024293f
C867 VTAIL.n719 B 0.010882f
C868 VTAIL.n720 B 0.010278f
C869 VTAIL.n721 B 0.019127f
C870 VTAIL.n722 B 0.019127f
C871 VTAIL.n723 B 0.010278f
C872 VTAIL.n724 B 0.010882f
C873 VTAIL.n725 B 0.024293f
C874 VTAIL.n726 B 0.024293f
C875 VTAIL.n727 B 0.010882f
C876 VTAIL.n728 B 0.010278f
C877 VTAIL.n729 B 0.019127f
C878 VTAIL.n730 B 0.019127f
C879 VTAIL.n731 B 0.010278f
C880 VTAIL.n732 B 0.010882f
C881 VTAIL.n733 B 0.024293f
C882 VTAIL.n734 B 0.024293f
C883 VTAIL.n735 B 0.010882f
C884 VTAIL.n736 B 0.010278f
C885 VTAIL.n737 B 0.019127f
C886 VTAIL.n738 B 0.049959f
C887 VTAIL.n739 B 0.010278f
C888 VTAIL.n740 B 0.010882f
C889 VTAIL.n741 B 0.04757f
C890 VTAIL.n742 B 0.040989f
C891 VTAIL.n743 B 1.5361f
C892 VN.t7 B 2.7273f
C893 VN.n0 B 1.01682f
C894 VN.n1 B 0.018511f
C895 VN.n2 B 0.015549f
C896 VN.n3 B 0.018511f
C897 VN.t6 B 2.7273f
C898 VN.n4 B 0.944607f
C899 VN.n5 B 0.018511f
C900 VN.n6 B 0.014951f
C901 VN.n7 B 0.018511f
C902 VN.t3 B 2.7273f
C903 VN.n8 B 1.00608f
C904 VN.t1 B 2.95324f
C905 VN.n9 B 0.96454f
C906 VN.n10 B 0.215212f
C907 VN.n11 B 0.026702f
C908 VN.n12 B 0.034328f
C909 VN.n13 B 0.036598f
C910 VN.n14 B 0.018511f
C911 VN.n15 B 0.018511f
C912 VN.n16 B 0.018511f
C913 VN.n17 B 0.036598f
C914 VN.n18 B 0.034328f
C915 VN.n19 B 0.026702f
C916 VN.n20 B 0.018511f
C917 VN.n21 B 0.018511f
C918 VN.n22 B 0.025007f
C919 VN.n23 B 0.034328f
C920 VN.n24 B 0.037181f
C921 VN.n25 B 0.018511f
C922 VN.n26 B 0.018511f
C923 VN.n27 B 0.018511f
C924 VN.n28 B 0.035416f
C925 VN.n29 B 0.034328f
C926 VN.n30 B 0.028396f
C927 VN.n31 B 0.029872f
C928 VN.n32 B 0.043237f
C929 VN.t4 B 2.7273f
C930 VN.n33 B 1.01682f
C931 VN.n34 B 0.018511f
C932 VN.n35 B 0.015549f
C933 VN.n36 B 0.018511f
C934 VN.t0 B 2.7273f
C935 VN.n37 B 0.944607f
C936 VN.n38 B 0.018511f
C937 VN.n39 B 0.014951f
C938 VN.n40 B 0.018511f
C939 VN.t2 B 2.7273f
C940 VN.n41 B 1.00608f
C941 VN.t5 B 2.95324f
C942 VN.n42 B 0.96454f
C943 VN.n43 B 0.215212f
C944 VN.n44 B 0.026702f
C945 VN.n45 B 0.034328f
C946 VN.n46 B 0.036598f
C947 VN.n47 B 0.018511f
C948 VN.n48 B 0.018511f
C949 VN.n49 B 0.018511f
C950 VN.n50 B 0.036598f
C951 VN.n51 B 0.034328f
C952 VN.n52 B 0.026702f
C953 VN.n53 B 0.018511f
C954 VN.n54 B 0.018511f
C955 VN.n55 B 0.025007f
C956 VN.n56 B 0.034328f
C957 VN.n57 B 0.037181f
C958 VN.n58 B 0.018511f
C959 VN.n59 B 0.018511f
C960 VN.n60 B 0.018511f
C961 VN.n61 B 0.035416f
C962 VN.n62 B 0.034328f
C963 VN.n63 B 0.028396f
C964 VN.n64 B 0.029872f
C965 VN.n65 B 1.2836f
.ends

