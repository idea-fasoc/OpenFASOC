* NGSPICE file created from diff_pair_sample_0108.ext - technology: sky130A

.subckt diff_pair_sample_0108 VTAIL VN VP B VDD2 VDD1
X0 B.t11 B.t9 B.t10 w_n4582_n2676# sky130_fd_pr__pfet_01v8 ad=3.3306 pd=17.86 as=0 ps=0 w=8.54 l=2.68
X1 VTAIL.t19 VN.t0 VDD2.t5 w_n4582_n2676# sky130_fd_pr__pfet_01v8 ad=1.4091 pd=8.87 as=1.4091 ps=8.87 w=8.54 l=2.68
X2 VDD1.t9 VP.t0 VTAIL.t2 w_n4582_n2676# sky130_fd_pr__pfet_01v8 ad=1.4091 pd=8.87 as=1.4091 ps=8.87 w=8.54 l=2.68
X3 VDD1.t8 VP.t1 VTAIL.t4 w_n4582_n2676# sky130_fd_pr__pfet_01v8 ad=3.3306 pd=17.86 as=1.4091 ps=8.87 w=8.54 l=2.68
X4 VDD1.t7 VP.t2 VTAIL.t3 w_n4582_n2676# sky130_fd_pr__pfet_01v8 ad=1.4091 pd=8.87 as=1.4091 ps=8.87 w=8.54 l=2.68
X5 B.t8 B.t6 B.t7 w_n4582_n2676# sky130_fd_pr__pfet_01v8 ad=3.3306 pd=17.86 as=0 ps=0 w=8.54 l=2.68
X6 VTAIL.t18 VN.t1 VDD2.t9 w_n4582_n2676# sky130_fd_pr__pfet_01v8 ad=1.4091 pd=8.87 as=1.4091 ps=8.87 w=8.54 l=2.68
X7 B.t5 B.t3 B.t4 w_n4582_n2676# sky130_fd_pr__pfet_01v8 ad=3.3306 pd=17.86 as=0 ps=0 w=8.54 l=2.68
X8 VDD2.t7 VN.t2 VTAIL.t17 w_n4582_n2676# sky130_fd_pr__pfet_01v8 ad=1.4091 pd=8.87 as=1.4091 ps=8.87 w=8.54 l=2.68
X9 VDD2.t1 VN.t3 VTAIL.t16 w_n4582_n2676# sky130_fd_pr__pfet_01v8 ad=1.4091 pd=8.87 as=3.3306 ps=17.86 w=8.54 l=2.68
X10 VTAIL.t0 VP.t3 VDD1.t6 w_n4582_n2676# sky130_fd_pr__pfet_01v8 ad=1.4091 pd=8.87 as=1.4091 ps=8.87 w=8.54 l=2.68
X11 VTAIL.t5 VP.t4 VDD1.t5 w_n4582_n2676# sky130_fd_pr__pfet_01v8 ad=1.4091 pd=8.87 as=1.4091 ps=8.87 w=8.54 l=2.68
X12 VDD2.t6 VN.t4 VTAIL.t15 w_n4582_n2676# sky130_fd_pr__pfet_01v8 ad=3.3306 pd=17.86 as=1.4091 ps=8.87 w=8.54 l=2.68
X13 VDD1.t4 VP.t5 VTAIL.t8 w_n4582_n2676# sky130_fd_pr__pfet_01v8 ad=3.3306 pd=17.86 as=1.4091 ps=8.87 w=8.54 l=2.68
X14 VTAIL.t9 VP.t6 VDD1.t3 w_n4582_n2676# sky130_fd_pr__pfet_01v8 ad=1.4091 pd=8.87 as=1.4091 ps=8.87 w=8.54 l=2.68
X15 VDD1.t2 VP.t7 VTAIL.t6 w_n4582_n2676# sky130_fd_pr__pfet_01v8 ad=1.4091 pd=8.87 as=3.3306 ps=17.86 w=8.54 l=2.68
X16 VDD2.t3 VN.t5 VTAIL.t14 w_n4582_n2676# sky130_fd_pr__pfet_01v8 ad=1.4091 pd=8.87 as=1.4091 ps=8.87 w=8.54 l=2.68
X17 VDD1.t1 VP.t8 VTAIL.t1 w_n4582_n2676# sky130_fd_pr__pfet_01v8 ad=1.4091 pd=8.87 as=3.3306 ps=17.86 w=8.54 l=2.68
X18 VTAIL.t13 VN.t6 VDD2.t0 w_n4582_n2676# sky130_fd_pr__pfet_01v8 ad=1.4091 pd=8.87 as=1.4091 ps=8.87 w=8.54 l=2.68
X19 VDD2.t8 VN.t7 VTAIL.t12 w_n4582_n2676# sky130_fd_pr__pfet_01v8 ad=1.4091 pd=8.87 as=3.3306 ps=17.86 w=8.54 l=2.68
X20 VDD2.t4 VN.t8 VTAIL.t11 w_n4582_n2676# sky130_fd_pr__pfet_01v8 ad=3.3306 pd=17.86 as=1.4091 ps=8.87 w=8.54 l=2.68
X21 B.t2 B.t0 B.t1 w_n4582_n2676# sky130_fd_pr__pfet_01v8 ad=3.3306 pd=17.86 as=0 ps=0 w=8.54 l=2.68
X22 VTAIL.t10 VN.t9 VDD2.t2 w_n4582_n2676# sky130_fd_pr__pfet_01v8 ad=1.4091 pd=8.87 as=1.4091 ps=8.87 w=8.54 l=2.68
X23 VTAIL.t7 VP.t9 VDD1.t0 w_n4582_n2676# sky130_fd_pr__pfet_01v8 ad=1.4091 pd=8.87 as=1.4091 ps=8.87 w=8.54 l=2.68
R0 B.n590 B.n589 585
R1 B.n591 B.n72 585
R2 B.n593 B.n592 585
R3 B.n594 B.n71 585
R4 B.n596 B.n595 585
R5 B.n597 B.n70 585
R6 B.n599 B.n598 585
R7 B.n600 B.n69 585
R8 B.n602 B.n601 585
R9 B.n603 B.n68 585
R10 B.n605 B.n604 585
R11 B.n606 B.n67 585
R12 B.n608 B.n607 585
R13 B.n609 B.n66 585
R14 B.n611 B.n610 585
R15 B.n612 B.n65 585
R16 B.n614 B.n613 585
R17 B.n615 B.n64 585
R18 B.n617 B.n616 585
R19 B.n618 B.n63 585
R20 B.n620 B.n619 585
R21 B.n621 B.n62 585
R22 B.n623 B.n622 585
R23 B.n624 B.n61 585
R24 B.n626 B.n625 585
R25 B.n627 B.n60 585
R26 B.n629 B.n628 585
R27 B.n630 B.n59 585
R28 B.n632 B.n631 585
R29 B.n633 B.n58 585
R30 B.n635 B.n634 585
R31 B.n637 B.n55 585
R32 B.n639 B.n638 585
R33 B.n640 B.n54 585
R34 B.n642 B.n641 585
R35 B.n643 B.n53 585
R36 B.n645 B.n644 585
R37 B.n646 B.n52 585
R38 B.n648 B.n647 585
R39 B.n649 B.n51 585
R40 B.n651 B.n650 585
R41 B.n653 B.n652 585
R42 B.n654 B.n47 585
R43 B.n656 B.n655 585
R44 B.n657 B.n46 585
R45 B.n659 B.n658 585
R46 B.n660 B.n45 585
R47 B.n662 B.n661 585
R48 B.n663 B.n44 585
R49 B.n665 B.n664 585
R50 B.n666 B.n43 585
R51 B.n668 B.n667 585
R52 B.n669 B.n42 585
R53 B.n671 B.n670 585
R54 B.n672 B.n41 585
R55 B.n674 B.n673 585
R56 B.n675 B.n40 585
R57 B.n677 B.n676 585
R58 B.n678 B.n39 585
R59 B.n680 B.n679 585
R60 B.n681 B.n38 585
R61 B.n683 B.n682 585
R62 B.n684 B.n37 585
R63 B.n686 B.n685 585
R64 B.n687 B.n36 585
R65 B.n689 B.n688 585
R66 B.n690 B.n35 585
R67 B.n692 B.n691 585
R68 B.n693 B.n34 585
R69 B.n695 B.n694 585
R70 B.n696 B.n33 585
R71 B.n698 B.n697 585
R72 B.n588 B.n73 585
R73 B.n587 B.n586 585
R74 B.n585 B.n74 585
R75 B.n584 B.n583 585
R76 B.n582 B.n75 585
R77 B.n581 B.n580 585
R78 B.n579 B.n76 585
R79 B.n578 B.n577 585
R80 B.n576 B.n77 585
R81 B.n575 B.n574 585
R82 B.n573 B.n78 585
R83 B.n572 B.n571 585
R84 B.n570 B.n79 585
R85 B.n569 B.n568 585
R86 B.n567 B.n80 585
R87 B.n566 B.n565 585
R88 B.n564 B.n81 585
R89 B.n563 B.n562 585
R90 B.n561 B.n82 585
R91 B.n560 B.n559 585
R92 B.n558 B.n83 585
R93 B.n557 B.n556 585
R94 B.n555 B.n84 585
R95 B.n554 B.n553 585
R96 B.n552 B.n85 585
R97 B.n551 B.n550 585
R98 B.n549 B.n86 585
R99 B.n548 B.n547 585
R100 B.n546 B.n87 585
R101 B.n545 B.n544 585
R102 B.n543 B.n88 585
R103 B.n542 B.n541 585
R104 B.n540 B.n89 585
R105 B.n539 B.n538 585
R106 B.n537 B.n90 585
R107 B.n536 B.n535 585
R108 B.n534 B.n91 585
R109 B.n533 B.n532 585
R110 B.n531 B.n92 585
R111 B.n530 B.n529 585
R112 B.n528 B.n93 585
R113 B.n527 B.n526 585
R114 B.n525 B.n94 585
R115 B.n524 B.n523 585
R116 B.n522 B.n95 585
R117 B.n521 B.n520 585
R118 B.n519 B.n96 585
R119 B.n518 B.n517 585
R120 B.n516 B.n97 585
R121 B.n515 B.n514 585
R122 B.n513 B.n98 585
R123 B.n512 B.n511 585
R124 B.n510 B.n99 585
R125 B.n509 B.n508 585
R126 B.n507 B.n100 585
R127 B.n506 B.n505 585
R128 B.n504 B.n101 585
R129 B.n503 B.n502 585
R130 B.n501 B.n102 585
R131 B.n500 B.n499 585
R132 B.n498 B.n103 585
R133 B.n497 B.n496 585
R134 B.n495 B.n104 585
R135 B.n494 B.n493 585
R136 B.n492 B.n105 585
R137 B.n491 B.n490 585
R138 B.n489 B.n106 585
R139 B.n488 B.n487 585
R140 B.n486 B.n107 585
R141 B.n485 B.n484 585
R142 B.n483 B.n108 585
R143 B.n482 B.n481 585
R144 B.n480 B.n109 585
R145 B.n479 B.n478 585
R146 B.n477 B.n110 585
R147 B.n476 B.n475 585
R148 B.n474 B.n111 585
R149 B.n473 B.n472 585
R150 B.n471 B.n112 585
R151 B.n470 B.n469 585
R152 B.n468 B.n113 585
R153 B.n467 B.n466 585
R154 B.n465 B.n114 585
R155 B.n464 B.n463 585
R156 B.n462 B.n115 585
R157 B.n461 B.n460 585
R158 B.n459 B.n116 585
R159 B.n458 B.n457 585
R160 B.n456 B.n117 585
R161 B.n455 B.n454 585
R162 B.n453 B.n118 585
R163 B.n452 B.n451 585
R164 B.n450 B.n119 585
R165 B.n449 B.n448 585
R166 B.n447 B.n120 585
R167 B.n446 B.n445 585
R168 B.n444 B.n121 585
R169 B.n443 B.n442 585
R170 B.n441 B.n122 585
R171 B.n440 B.n439 585
R172 B.n438 B.n123 585
R173 B.n437 B.n436 585
R174 B.n435 B.n124 585
R175 B.n434 B.n433 585
R176 B.n432 B.n125 585
R177 B.n431 B.n430 585
R178 B.n429 B.n126 585
R179 B.n428 B.n427 585
R180 B.n426 B.n127 585
R181 B.n425 B.n424 585
R182 B.n423 B.n128 585
R183 B.n422 B.n421 585
R184 B.n420 B.n129 585
R185 B.n419 B.n418 585
R186 B.n417 B.n130 585
R187 B.n416 B.n415 585
R188 B.n414 B.n131 585
R189 B.n413 B.n412 585
R190 B.n411 B.n132 585
R191 B.n410 B.n409 585
R192 B.n408 B.n133 585
R193 B.n407 B.n406 585
R194 B.n405 B.n134 585
R195 B.n296 B.n295 585
R196 B.n297 B.n174 585
R197 B.n299 B.n298 585
R198 B.n300 B.n173 585
R199 B.n302 B.n301 585
R200 B.n303 B.n172 585
R201 B.n305 B.n304 585
R202 B.n306 B.n171 585
R203 B.n308 B.n307 585
R204 B.n309 B.n170 585
R205 B.n311 B.n310 585
R206 B.n312 B.n169 585
R207 B.n314 B.n313 585
R208 B.n315 B.n168 585
R209 B.n317 B.n316 585
R210 B.n318 B.n167 585
R211 B.n320 B.n319 585
R212 B.n321 B.n166 585
R213 B.n323 B.n322 585
R214 B.n324 B.n165 585
R215 B.n326 B.n325 585
R216 B.n327 B.n164 585
R217 B.n329 B.n328 585
R218 B.n330 B.n163 585
R219 B.n332 B.n331 585
R220 B.n333 B.n162 585
R221 B.n335 B.n334 585
R222 B.n336 B.n161 585
R223 B.n338 B.n337 585
R224 B.n339 B.n160 585
R225 B.n341 B.n340 585
R226 B.n343 B.n157 585
R227 B.n345 B.n344 585
R228 B.n346 B.n156 585
R229 B.n348 B.n347 585
R230 B.n349 B.n155 585
R231 B.n351 B.n350 585
R232 B.n352 B.n154 585
R233 B.n354 B.n353 585
R234 B.n355 B.n153 585
R235 B.n357 B.n356 585
R236 B.n359 B.n358 585
R237 B.n360 B.n149 585
R238 B.n362 B.n361 585
R239 B.n363 B.n148 585
R240 B.n365 B.n364 585
R241 B.n366 B.n147 585
R242 B.n368 B.n367 585
R243 B.n369 B.n146 585
R244 B.n371 B.n370 585
R245 B.n372 B.n145 585
R246 B.n374 B.n373 585
R247 B.n375 B.n144 585
R248 B.n377 B.n376 585
R249 B.n378 B.n143 585
R250 B.n380 B.n379 585
R251 B.n381 B.n142 585
R252 B.n383 B.n382 585
R253 B.n384 B.n141 585
R254 B.n386 B.n385 585
R255 B.n387 B.n140 585
R256 B.n389 B.n388 585
R257 B.n390 B.n139 585
R258 B.n392 B.n391 585
R259 B.n393 B.n138 585
R260 B.n395 B.n394 585
R261 B.n396 B.n137 585
R262 B.n398 B.n397 585
R263 B.n399 B.n136 585
R264 B.n401 B.n400 585
R265 B.n402 B.n135 585
R266 B.n404 B.n403 585
R267 B.n294 B.n175 585
R268 B.n293 B.n292 585
R269 B.n291 B.n176 585
R270 B.n290 B.n289 585
R271 B.n288 B.n177 585
R272 B.n287 B.n286 585
R273 B.n285 B.n178 585
R274 B.n284 B.n283 585
R275 B.n282 B.n179 585
R276 B.n281 B.n280 585
R277 B.n279 B.n180 585
R278 B.n278 B.n277 585
R279 B.n276 B.n181 585
R280 B.n275 B.n274 585
R281 B.n273 B.n182 585
R282 B.n272 B.n271 585
R283 B.n270 B.n183 585
R284 B.n269 B.n268 585
R285 B.n267 B.n184 585
R286 B.n266 B.n265 585
R287 B.n264 B.n185 585
R288 B.n263 B.n262 585
R289 B.n261 B.n186 585
R290 B.n260 B.n259 585
R291 B.n258 B.n187 585
R292 B.n257 B.n256 585
R293 B.n255 B.n188 585
R294 B.n254 B.n253 585
R295 B.n252 B.n189 585
R296 B.n251 B.n250 585
R297 B.n249 B.n190 585
R298 B.n248 B.n247 585
R299 B.n246 B.n191 585
R300 B.n245 B.n244 585
R301 B.n243 B.n192 585
R302 B.n242 B.n241 585
R303 B.n240 B.n193 585
R304 B.n239 B.n238 585
R305 B.n237 B.n194 585
R306 B.n236 B.n235 585
R307 B.n234 B.n195 585
R308 B.n233 B.n232 585
R309 B.n231 B.n196 585
R310 B.n230 B.n229 585
R311 B.n228 B.n197 585
R312 B.n227 B.n226 585
R313 B.n225 B.n198 585
R314 B.n224 B.n223 585
R315 B.n222 B.n199 585
R316 B.n221 B.n220 585
R317 B.n219 B.n200 585
R318 B.n218 B.n217 585
R319 B.n216 B.n201 585
R320 B.n215 B.n214 585
R321 B.n213 B.n202 585
R322 B.n212 B.n211 585
R323 B.n210 B.n203 585
R324 B.n209 B.n208 585
R325 B.n207 B.n204 585
R326 B.n206 B.n205 585
R327 B.n2 B.n0 585
R328 B.n789 B.n1 585
R329 B.n788 B.n787 585
R330 B.n786 B.n3 585
R331 B.n785 B.n784 585
R332 B.n783 B.n4 585
R333 B.n782 B.n781 585
R334 B.n780 B.n5 585
R335 B.n779 B.n778 585
R336 B.n777 B.n6 585
R337 B.n776 B.n775 585
R338 B.n774 B.n7 585
R339 B.n773 B.n772 585
R340 B.n771 B.n8 585
R341 B.n770 B.n769 585
R342 B.n768 B.n9 585
R343 B.n767 B.n766 585
R344 B.n765 B.n10 585
R345 B.n764 B.n763 585
R346 B.n762 B.n11 585
R347 B.n761 B.n760 585
R348 B.n759 B.n12 585
R349 B.n758 B.n757 585
R350 B.n756 B.n13 585
R351 B.n755 B.n754 585
R352 B.n753 B.n14 585
R353 B.n752 B.n751 585
R354 B.n750 B.n15 585
R355 B.n749 B.n748 585
R356 B.n747 B.n16 585
R357 B.n746 B.n745 585
R358 B.n744 B.n17 585
R359 B.n743 B.n742 585
R360 B.n741 B.n18 585
R361 B.n740 B.n739 585
R362 B.n738 B.n19 585
R363 B.n737 B.n736 585
R364 B.n735 B.n20 585
R365 B.n734 B.n733 585
R366 B.n732 B.n21 585
R367 B.n731 B.n730 585
R368 B.n729 B.n22 585
R369 B.n728 B.n727 585
R370 B.n726 B.n23 585
R371 B.n725 B.n724 585
R372 B.n723 B.n24 585
R373 B.n722 B.n721 585
R374 B.n720 B.n25 585
R375 B.n719 B.n718 585
R376 B.n717 B.n26 585
R377 B.n716 B.n715 585
R378 B.n714 B.n27 585
R379 B.n713 B.n712 585
R380 B.n711 B.n28 585
R381 B.n710 B.n709 585
R382 B.n708 B.n29 585
R383 B.n707 B.n706 585
R384 B.n705 B.n30 585
R385 B.n704 B.n703 585
R386 B.n702 B.n31 585
R387 B.n701 B.n700 585
R388 B.n699 B.n32 585
R389 B.n791 B.n790 585
R390 B.n296 B.n175 574.183
R391 B.n699 B.n698 574.183
R392 B.n405 B.n404 574.183
R393 B.n590 B.n73 574.183
R394 B.n150 B.t8 371.555
R395 B.n56 B.t1 371.555
R396 B.n158 B.t5 371.555
R397 B.n48 B.t10 371.555
R398 B.n151 B.t7 313.18
R399 B.n57 B.t2 313.18
R400 B.n159 B.t4 313.18
R401 B.n49 B.t11 313.18
R402 B.n150 B.t6 284.961
R403 B.n158 B.t3 284.961
R404 B.n48 B.t9 284.961
R405 B.n56 B.t0 284.961
R406 B.n292 B.n175 163.367
R407 B.n292 B.n291 163.367
R408 B.n291 B.n290 163.367
R409 B.n290 B.n177 163.367
R410 B.n286 B.n177 163.367
R411 B.n286 B.n285 163.367
R412 B.n285 B.n284 163.367
R413 B.n284 B.n179 163.367
R414 B.n280 B.n179 163.367
R415 B.n280 B.n279 163.367
R416 B.n279 B.n278 163.367
R417 B.n278 B.n181 163.367
R418 B.n274 B.n181 163.367
R419 B.n274 B.n273 163.367
R420 B.n273 B.n272 163.367
R421 B.n272 B.n183 163.367
R422 B.n268 B.n183 163.367
R423 B.n268 B.n267 163.367
R424 B.n267 B.n266 163.367
R425 B.n266 B.n185 163.367
R426 B.n262 B.n185 163.367
R427 B.n262 B.n261 163.367
R428 B.n261 B.n260 163.367
R429 B.n260 B.n187 163.367
R430 B.n256 B.n187 163.367
R431 B.n256 B.n255 163.367
R432 B.n255 B.n254 163.367
R433 B.n254 B.n189 163.367
R434 B.n250 B.n189 163.367
R435 B.n250 B.n249 163.367
R436 B.n249 B.n248 163.367
R437 B.n248 B.n191 163.367
R438 B.n244 B.n191 163.367
R439 B.n244 B.n243 163.367
R440 B.n243 B.n242 163.367
R441 B.n242 B.n193 163.367
R442 B.n238 B.n193 163.367
R443 B.n238 B.n237 163.367
R444 B.n237 B.n236 163.367
R445 B.n236 B.n195 163.367
R446 B.n232 B.n195 163.367
R447 B.n232 B.n231 163.367
R448 B.n231 B.n230 163.367
R449 B.n230 B.n197 163.367
R450 B.n226 B.n197 163.367
R451 B.n226 B.n225 163.367
R452 B.n225 B.n224 163.367
R453 B.n224 B.n199 163.367
R454 B.n220 B.n199 163.367
R455 B.n220 B.n219 163.367
R456 B.n219 B.n218 163.367
R457 B.n218 B.n201 163.367
R458 B.n214 B.n201 163.367
R459 B.n214 B.n213 163.367
R460 B.n213 B.n212 163.367
R461 B.n212 B.n203 163.367
R462 B.n208 B.n203 163.367
R463 B.n208 B.n207 163.367
R464 B.n207 B.n206 163.367
R465 B.n206 B.n2 163.367
R466 B.n790 B.n2 163.367
R467 B.n790 B.n789 163.367
R468 B.n789 B.n788 163.367
R469 B.n788 B.n3 163.367
R470 B.n784 B.n3 163.367
R471 B.n784 B.n783 163.367
R472 B.n783 B.n782 163.367
R473 B.n782 B.n5 163.367
R474 B.n778 B.n5 163.367
R475 B.n778 B.n777 163.367
R476 B.n777 B.n776 163.367
R477 B.n776 B.n7 163.367
R478 B.n772 B.n7 163.367
R479 B.n772 B.n771 163.367
R480 B.n771 B.n770 163.367
R481 B.n770 B.n9 163.367
R482 B.n766 B.n9 163.367
R483 B.n766 B.n765 163.367
R484 B.n765 B.n764 163.367
R485 B.n764 B.n11 163.367
R486 B.n760 B.n11 163.367
R487 B.n760 B.n759 163.367
R488 B.n759 B.n758 163.367
R489 B.n758 B.n13 163.367
R490 B.n754 B.n13 163.367
R491 B.n754 B.n753 163.367
R492 B.n753 B.n752 163.367
R493 B.n752 B.n15 163.367
R494 B.n748 B.n15 163.367
R495 B.n748 B.n747 163.367
R496 B.n747 B.n746 163.367
R497 B.n746 B.n17 163.367
R498 B.n742 B.n17 163.367
R499 B.n742 B.n741 163.367
R500 B.n741 B.n740 163.367
R501 B.n740 B.n19 163.367
R502 B.n736 B.n19 163.367
R503 B.n736 B.n735 163.367
R504 B.n735 B.n734 163.367
R505 B.n734 B.n21 163.367
R506 B.n730 B.n21 163.367
R507 B.n730 B.n729 163.367
R508 B.n729 B.n728 163.367
R509 B.n728 B.n23 163.367
R510 B.n724 B.n23 163.367
R511 B.n724 B.n723 163.367
R512 B.n723 B.n722 163.367
R513 B.n722 B.n25 163.367
R514 B.n718 B.n25 163.367
R515 B.n718 B.n717 163.367
R516 B.n717 B.n716 163.367
R517 B.n716 B.n27 163.367
R518 B.n712 B.n27 163.367
R519 B.n712 B.n711 163.367
R520 B.n711 B.n710 163.367
R521 B.n710 B.n29 163.367
R522 B.n706 B.n29 163.367
R523 B.n706 B.n705 163.367
R524 B.n705 B.n704 163.367
R525 B.n704 B.n31 163.367
R526 B.n700 B.n31 163.367
R527 B.n700 B.n699 163.367
R528 B.n297 B.n296 163.367
R529 B.n298 B.n297 163.367
R530 B.n298 B.n173 163.367
R531 B.n302 B.n173 163.367
R532 B.n303 B.n302 163.367
R533 B.n304 B.n303 163.367
R534 B.n304 B.n171 163.367
R535 B.n308 B.n171 163.367
R536 B.n309 B.n308 163.367
R537 B.n310 B.n309 163.367
R538 B.n310 B.n169 163.367
R539 B.n314 B.n169 163.367
R540 B.n315 B.n314 163.367
R541 B.n316 B.n315 163.367
R542 B.n316 B.n167 163.367
R543 B.n320 B.n167 163.367
R544 B.n321 B.n320 163.367
R545 B.n322 B.n321 163.367
R546 B.n322 B.n165 163.367
R547 B.n326 B.n165 163.367
R548 B.n327 B.n326 163.367
R549 B.n328 B.n327 163.367
R550 B.n328 B.n163 163.367
R551 B.n332 B.n163 163.367
R552 B.n333 B.n332 163.367
R553 B.n334 B.n333 163.367
R554 B.n334 B.n161 163.367
R555 B.n338 B.n161 163.367
R556 B.n339 B.n338 163.367
R557 B.n340 B.n339 163.367
R558 B.n340 B.n157 163.367
R559 B.n345 B.n157 163.367
R560 B.n346 B.n345 163.367
R561 B.n347 B.n346 163.367
R562 B.n347 B.n155 163.367
R563 B.n351 B.n155 163.367
R564 B.n352 B.n351 163.367
R565 B.n353 B.n352 163.367
R566 B.n353 B.n153 163.367
R567 B.n357 B.n153 163.367
R568 B.n358 B.n357 163.367
R569 B.n358 B.n149 163.367
R570 B.n362 B.n149 163.367
R571 B.n363 B.n362 163.367
R572 B.n364 B.n363 163.367
R573 B.n364 B.n147 163.367
R574 B.n368 B.n147 163.367
R575 B.n369 B.n368 163.367
R576 B.n370 B.n369 163.367
R577 B.n370 B.n145 163.367
R578 B.n374 B.n145 163.367
R579 B.n375 B.n374 163.367
R580 B.n376 B.n375 163.367
R581 B.n376 B.n143 163.367
R582 B.n380 B.n143 163.367
R583 B.n381 B.n380 163.367
R584 B.n382 B.n381 163.367
R585 B.n382 B.n141 163.367
R586 B.n386 B.n141 163.367
R587 B.n387 B.n386 163.367
R588 B.n388 B.n387 163.367
R589 B.n388 B.n139 163.367
R590 B.n392 B.n139 163.367
R591 B.n393 B.n392 163.367
R592 B.n394 B.n393 163.367
R593 B.n394 B.n137 163.367
R594 B.n398 B.n137 163.367
R595 B.n399 B.n398 163.367
R596 B.n400 B.n399 163.367
R597 B.n400 B.n135 163.367
R598 B.n404 B.n135 163.367
R599 B.n406 B.n405 163.367
R600 B.n406 B.n133 163.367
R601 B.n410 B.n133 163.367
R602 B.n411 B.n410 163.367
R603 B.n412 B.n411 163.367
R604 B.n412 B.n131 163.367
R605 B.n416 B.n131 163.367
R606 B.n417 B.n416 163.367
R607 B.n418 B.n417 163.367
R608 B.n418 B.n129 163.367
R609 B.n422 B.n129 163.367
R610 B.n423 B.n422 163.367
R611 B.n424 B.n423 163.367
R612 B.n424 B.n127 163.367
R613 B.n428 B.n127 163.367
R614 B.n429 B.n428 163.367
R615 B.n430 B.n429 163.367
R616 B.n430 B.n125 163.367
R617 B.n434 B.n125 163.367
R618 B.n435 B.n434 163.367
R619 B.n436 B.n435 163.367
R620 B.n436 B.n123 163.367
R621 B.n440 B.n123 163.367
R622 B.n441 B.n440 163.367
R623 B.n442 B.n441 163.367
R624 B.n442 B.n121 163.367
R625 B.n446 B.n121 163.367
R626 B.n447 B.n446 163.367
R627 B.n448 B.n447 163.367
R628 B.n448 B.n119 163.367
R629 B.n452 B.n119 163.367
R630 B.n453 B.n452 163.367
R631 B.n454 B.n453 163.367
R632 B.n454 B.n117 163.367
R633 B.n458 B.n117 163.367
R634 B.n459 B.n458 163.367
R635 B.n460 B.n459 163.367
R636 B.n460 B.n115 163.367
R637 B.n464 B.n115 163.367
R638 B.n465 B.n464 163.367
R639 B.n466 B.n465 163.367
R640 B.n466 B.n113 163.367
R641 B.n470 B.n113 163.367
R642 B.n471 B.n470 163.367
R643 B.n472 B.n471 163.367
R644 B.n472 B.n111 163.367
R645 B.n476 B.n111 163.367
R646 B.n477 B.n476 163.367
R647 B.n478 B.n477 163.367
R648 B.n478 B.n109 163.367
R649 B.n482 B.n109 163.367
R650 B.n483 B.n482 163.367
R651 B.n484 B.n483 163.367
R652 B.n484 B.n107 163.367
R653 B.n488 B.n107 163.367
R654 B.n489 B.n488 163.367
R655 B.n490 B.n489 163.367
R656 B.n490 B.n105 163.367
R657 B.n494 B.n105 163.367
R658 B.n495 B.n494 163.367
R659 B.n496 B.n495 163.367
R660 B.n496 B.n103 163.367
R661 B.n500 B.n103 163.367
R662 B.n501 B.n500 163.367
R663 B.n502 B.n501 163.367
R664 B.n502 B.n101 163.367
R665 B.n506 B.n101 163.367
R666 B.n507 B.n506 163.367
R667 B.n508 B.n507 163.367
R668 B.n508 B.n99 163.367
R669 B.n512 B.n99 163.367
R670 B.n513 B.n512 163.367
R671 B.n514 B.n513 163.367
R672 B.n514 B.n97 163.367
R673 B.n518 B.n97 163.367
R674 B.n519 B.n518 163.367
R675 B.n520 B.n519 163.367
R676 B.n520 B.n95 163.367
R677 B.n524 B.n95 163.367
R678 B.n525 B.n524 163.367
R679 B.n526 B.n525 163.367
R680 B.n526 B.n93 163.367
R681 B.n530 B.n93 163.367
R682 B.n531 B.n530 163.367
R683 B.n532 B.n531 163.367
R684 B.n532 B.n91 163.367
R685 B.n536 B.n91 163.367
R686 B.n537 B.n536 163.367
R687 B.n538 B.n537 163.367
R688 B.n538 B.n89 163.367
R689 B.n542 B.n89 163.367
R690 B.n543 B.n542 163.367
R691 B.n544 B.n543 163.367
R692 B.n544 B.n87 163.367
R693 B.n548 B.n87 163.367
R694 B.n549 B.n548 163.367
R695 B.n550 B.n549 163.367
R696 B.n550 B.n85 163.367
R697 B.n554 B.n85 163.367
R698 B.n555 B.n554 163.367
R699 B.n556 B.n555 163.367
R700 B.n556 B.n83 163.367
R701 B.n560 B.n83 163.367
R702 B.n561 B.n560 163.367
R703 B.n562 B.n561 163.367
R704 B.n562 B.n81 163.367
R705 B.n566 B.n81 163.367
R706 B.n567 B.n566 163.367
R707 B.n568 B.n567 163.367
R708 B.n568 B.n79 163.367
R709 B.n572 B.n79 163.367
R710 B.n573 B.n572 163.367
R711 B.n574 B.n573 163.367
R712 B.n574 B.n77 163.367
R713 B.n578 B.n77 163.367
R714 B.n579 B.n578 163.367
R715 B.n580 B.n579 163.367
R716 B.n580 B.n75 163.367
R717 B.n584 B.n75 163.367
R718 B.n585 B.n584 163.367
R719 B.n586 B.n585 163.367
R720 B.n586 B.n73 163.367
R721 B.n698 B.n33 163.367
R722 B.n694 B.n33 163.367
R723 B.n694 B.n693 163.367
R724 B.n693 B.n692 163.367
R725 B.n692 B.n35 163.367
R726 B.n688 B.n35 163.367
R727 B.n688 B.n687 163.367
R728 B.n687 B.n686 163.367
R729 B.n686 B.n37 163.367
R730 B.n682 B.n37 163.367
R731 B.n682 B.n681 163.367
R732 B.n681 B.n680 163.367
R733 B.n680 B.n39 163.367
R734 B.n676 B.n39 163.367
R735 B.n676 B.n675 163.367
R736 B.n675 B.n674 163.367
R737 B.n674 B.n41 163.367
R738 B.n670 B.n41 163.367
R739 B.n670 B.n669 163.367
R740 B.n669 B.n668 163.367
R741 B.n668 B.n43 163.367
R742 B.n664 B.n43 163.367
R743 B.n664 B.n663 163.367
R744 B.n663 B.n662 163.367
R745 B.n662 B.n45 163.367
R746 B.n658 B.n45 163.367
R747 B.n658 B.n657 163.367
R748 B.n657 B.n656 163.367
R749 B.n656 B.n47 163.367
R750 B.n652 B.n47 163.367
R751 B.n652 B.n651 163.367
R752 B.n651 B.n51 163.367
R753 B.n647 B.n51 163.367
R754 B.n647 B.n646 163.367
R755 B.n646 B.n645 163.367
R756 B.n645 B.n53 163.367
R757 B.n641 B.n53 163.367
R758 B.n641 B.n640 163.367
R759 B.n640 B.n639 163.367
R760 B.n639 B.n55 163.367
R761 B.n634 B.n55 163.367
R762 B.n634 B.n633 163.367
R763 B.n633 B.n632 163.367
R764 B.n632 B.n59 163.367
R765 B.n628 B.n59 163.367
R766 B.n628 B.n627 163.367
R767 B.n627 B.n626 163.367
R768 B.n626 B.n61 163.367
R769 B.n622 B.n61 163.367
R770 B.n622 B.n621 163.367
R771 B.n621 B.n620 163.367
R772 B.n620 B.n63 163.367
R773 B.n616 B.n63 163.367
R774 B.n616 B.n615 163.367
R775 B.n615 B.n614 163.367
R776 B.n614 B.n65 163.367
R777 B.n610 B.n65 163.367
R778 B.n610 B.n609 163.367
R779 B.n609 B.n608 163.367
R780 B.n608 B.n67 163.367
R781 B.n604 B.n67 163.367
R782 B.n604 B.n603 163.367
R783 B.n603 B.n602 163.367
R784 B.n602 B.n69 163.367
R785 B.n598 B.n69 163.367
R786 B.n598 B.n597 163.367
R787 B.n597 B.n596 163.367
R788 B.n596 B.n71 163.367
R789 B.n592 B.n71 163.367
R790 B.n592 B.n591 163.367
R791 B.n591 B.n590 163.367
R792 B.n152 B.n151 59.5399
R793 B.n342 B.n159 59.5399
R794 B.n50 B.n49 59.5399
R795 B.n636 B.n57 59.5399
R796 B.n151 B.n150 58.3763
R797 B.n159 B.n158 58.3763
R798 B.n49 B.n48 58.3763
R799 B.n57 B.n56 58.3763
R800 B.n697 B.n32 37.3078
R801 B.n589 B.n588 37.3078
R802 B.n403 B.n134 37.3078
R803 B.n295 B.n294 37.3078
R804 B B.n791 18.0485
R805 B.n697 B.n696 10.6151
R806 B.n696 B.n695 10.6151
R807 B.n695 B.n34 10.6151
R808 B.n691 B.n34 10.6151
R809 B.n691 B.n690 10.6151
R810 B.n690 B.n689 10.6151
R811 B.n689 B.n36 10.6151
R812 B.n685 B.n36 10.6151
R813 B.n685 B.n684 10.6151
R814 B.n684 B.n683 10.6151
R815 B.n683 B.n38 10.6151
R816 B.n679 B.n38 10.6151
R817 B.n679 B.n678 10.6151
R818 B.n678 B.n677 10.6151
R819 B.n677 B.n40 10.6151
R820 B.n673 B.n40 10.6151
R821 B.n673 B.n672 10.6151
R822 B.n672 B.n671 10.6151
R823 B.n671 B.n42 10.6151
R824 B.n667 B.n42 10.6151
R825 B.n667 B.n666 10.6151
R826 B.n666 B.n665 10.6151
R827 B.n665 B.n44 10.6151
R828 B.n661 B.n44 10.6151
R829 B.n661 B.n660 10.6151
R830 B.n660 B.n659 10.6151
R831 B.n659 B.n46 10.6151
R832 B.n655 B.n46 10.6151
R833 B.n655 B.n654 10.6151
R834 B.n654 B.n653 10.6151
R835 B.n650 B.n649 10.6151
R836 B.n649 B.n648 10.6151
R837 B.n648 B.n52 10.6151
R838 B.n644 B.n52 10.6151
R839 B.n644 B.n643 10.6151
R840 B.n643 B.n642 10.6151
R841 B.n642 B.n54 10.6151
R842 B.n638 B.n54 10.6151
R843 B.n638 B.n637 10.6151
R844 B.n635 B.n58 10.6151
R845 B.n631 B.n58 10.6151
R846 B.n631 B.n630 10.6151
R847 B.n630 B.n629 10.6151
R848 B.n629 B.n60 10.6151
R849 B.n625 B.n60 10.6151
R850 B.n625 B.n624 10.6151
R851 B.n624 B.n623 10.6151
R852 B.n623 B.n62 10.6151
R853 B.n619 B.n62 10.6151
R854 B.n619 B.n618 10.6151
R855 B.n618 B.n617 10.6151
R856 B.n617 B.n64 10.6151
R857 B.n613 B.n64 10.6151
R858 B.n613 B.n612 10.6151
R859 B.n612 B.n611 10.6151
R860 B.n611 B.n66 10.6151
R861 B.n607 B.n66 10.6151
R862 B.n607 B.n606 10.6151
R863 B.n606 B.n605 10.6151
R864 B.n605 B.n68 10.6151
R865 B.n601 B.n68 10.6151
R866 B.n601 B.n600 10.6151
R867 B.n600 B.n599 10.6151
R868 B.n599 B.n70 10.6151
R869 B.n595 B.n70 10.6151
R870 B.n595 B.n594 10.6151
R871 B.n594 B.n593 10.6151
R872 B.n593 B.n72 10.6151
R873 B.n589 B.n72 10.6151
R874 B.n407 B.n134 10.6151
R875 B.n408 B.n407 10.6151
R876 B.n409 B.n408 10.6151
R877 B.n409 B.n132 10.6151
R878 B.n413 B.n132 10.6151
R879 B.n414 B.n413 10.6151
R880 B.n415 B.n414 10.6151
R881 B.n415 B.n130 10.6151
R882 B.n419 B.n130 10.6151
R883 B.n420 B.n419 10.6151
R884 B.n421 B.n420 10.6151
R885 B.n421 B.n128 10.6151
R886 B.n425 B.n128 10.6151
R887 B.n426 B.n425 10.6151
R888 B.n427 B.n426 10.6151
R889 B.n427 B.n126 10.6151
R890 B.n431 B.n126 10.6151
R891 B.n432 B.n431 10.6151
R892 B.n433 B.n432 10.6151
R893 B.n433 B.n124 10.6151
R894 B.n437 B.n124 10.6151
R895 B.n438 B.n437 10.6151
R896 B.n439 B.n438 10.6151
R897 B.n439 B.n122 10.6151
R898 B.n443 B.n122 10.6151
R899 B.n444 B.n443 10.6151
R900 B.n445 B.n444 10.6151
R901 B.n445 B.n120 10.6151
R902 B.n449 B.n120 10.6151
R903 B.n450 B.n449 10.6151
R904 B.n451 B.n450 10.6151
R905 B.n451 B.n118 10.6151
R906 B.n455 B.n118 10.6151
R907 B.n456 B.n455 10.6151
R908 B.n457 B.n456 10.6151
R909 B.n457 B.n116 10.6151
R910 B.n461 B.n116 10.6151
R911 B.n462 B.n461 10.6151
R912 B.n463 B.n462 10.6151
R913 B.n463 B.n114 10.6151
R914 B.n467 B.n114 10.6151
R915 B.n468 B.n467 10.6151
R916 B.n469 B.n468 10.6151
R917 B.n469 B.n112 10.6151
R918 B.n473 B.n112 10.6151
R919 B.n474 B.n473 10.6151
R920 B.n475 B.n474 10.6151
R921 B.n475 B.n110 10.6151
R922 B.n479 B.n110 10.6151
R923 B.n480 B.n479 10.6151
R924 B.n481 B.n480 10.6151
R925 B.n481 B.n108 10.6151
R926 B.n485 B.n108 10.6151
R927 B.n486 B.n485 10.6151
R928 B.n487 B.n486 10.6151
R929 B.n487 B.n106 10.6151
R930 B.n491 B.n106 10.6151
R931 B.n492 B.n491 10.6151
R932 B.n493 B.n492 10.6151
R933 B.n493 B.n104 10.6151
R934 B.n497 B.n104 10.6151
R935 B.n498 B.n497 10.6151
R936 B.n499 B.n498 10.6151
R937 B.n499 B.n102 10.6151
R938 B.n503 B.n102 10.6151
R939 B.n504 B.n503 10.6151
R940 B.n505 B.n504 10.6151
R941 B.n505 B.n100 10.6151
R942 B.n509 B.n100 10.6151
R943 B.n510 B.n509 10.6151
R944 B.n511 B.n510 10.6151
R945 B.n511 B.n98 10.6151
R946 B.n515 B.n98 10.6151
R947 B.n516 B.n515 10.6151
R948 B.n517 B.n516 10.6151
R949 B.n517 B.n96 10.6151
R950 B.n521 B.n96 10.6151
R951 B.n522 B.n521 10.6151
R952 B.n523 B.n522 10.6151
R953 B.n523 B.n94 10.6151
R954 B.n527 B.n94 10.6151
R955 B.n528 B.n527 10.6151
R956 B.n529 B.n528 10.6151
R957 B.n529 B.n92 10.6151
R958 B.n533 B.n92 10.6151
R959 B.n534 B.n533 10.6151
R960 B.n535 B.n534 10.6151
R961 B.n535 B.n90 10.6151
R962 B.n539 B.n90 10.6151
R963 B.n540 B.n539 10.6151
R964 B.n541 B.n540 10.6151
R965 B.n541 B.n88 10.6151
R966 B.n545 B.n88 10.6151
R967 B.n546 B.n545 10.6151
R968 B.n547 B.n546 10.6151
R969 B.n547 B.n86 10.6151
R970 B.n551 B.n86 10.6151
R971 B.n552 B.n551 10.6151
R972 B.n553 B.n552 10.6151
R973 B.n553 B.n84 10.6151
R974 B.n557 B.n84 10.6151
R975 B.n558 B.n557 10.6151
R976 B.n559 B.n558 10.6151
R977 B.n559 B.n82 10.6151
R978 B.n563 B.n82 10.6151
R979 B.n564 B.n563 10.6151
R980 B.n565 B.n564 10.6151
R981 B.n565 B.n80 10.6151
R982 B.n569 B.n80 10.6151
R983 B.n570 B.n569 10.6151
R984 B.n571 B.n570 10.6151
R985 B.n571 B.n78 10.6151
R986 B.n575 B.n78 10.6151
R987 B.n576 B.n575 10.6151
R988 B.n577 B.n576 10.6151
R989 B.n577 B.n76 10.6151
R990 B.n581 B.n76 10.6151
R991 B.n582 B.n581 10.6151
R992 B.n583 B.n582 10.6151
R993 B.n583 B.n74 10.6151
R994 B.n587 B.n74 10.6151
R995 B.n588 B.n587 10.6151
R996 B.n295 B.n174 10.6151
R997 B.n299 B.n174 10.6151
R998 B.n300 B.n299 10.6151
R999 B.n301 B.n300 10.6151
R1000 B.n301 B.n172 10.6151
R1001 B.n305 B.n172 10.6151
R1002 B.n306 B.n305 10.6151
R1003 B.n307 B.n306 10.6151
R1004 B.n307 B.n170 10.6151
R1005 B.n311 B.n170 10.6151
R1006 B.n312 B.n311 10.6151
R1007 B.n313 B.n312 10.6151
R1008 B.n313 B.n168 10.6151
R1009 B.n317 B.n168 10.6151
R1010 B.n318 B.n317 10.6151
R1011 B.n319 B.n318 10.6151
R1012 B.n319 B.n166 10.6151
R1013 B.n323 B.n166 10.6151
R1014 B.n324 B.n323 10.6151
R1015 B.n325 B.n324 10.6151
R1016 B.n325 B.n164 10.6151
R1017 B.n329 B.n164 10.6151
R1018 B.n330 B.n329 10.6151
R1019 B.n331 B.n330 10.6151
R1020 B.n331 B.n162 10.6151
R1021 B.n335 B.n162 10.6151
R1022 B.n336 B.n335 10.6151
R1023 B.n337 B.n336 10.6151
R1024 B.n337 B.n160 10.6151
R1025 B.n341 B.n160 10.6151
R1026 B.n344 B.n343 10.6151
R1027 B.n344 B.n156 10.6151
R1028 B.n348 B.n156 10.6151
R1029 B.n349 B.n348 10.6151
R1030 B.n350 B.n349 10.6151
R1031 B.n350 B.n154 10.6151
R1032 B.n354 B.n154 10.6151
R1033 B.n355 B.n354 10.6151
R1034 B.n356 B.n355 10.6151
R1035 B.n360 B.n359 10.6151
R1036 B.n361 B.n360 10.6151
R1037 B.n361 B.n148 10.6151
R1038 B.n365 B.n148 10.6151
R1039 B.n366 B.n365 10.6151
R1040 B.n367 B.n366 10.6151
R1041 B.n367 B.n146 10.6151
R1042 B.n371 B.n146 10.6151
R1043 B.n372 B.n371 10.6151
R1044 B.n373 B.n372 10.6151
R1045 B.n373 B.n144 10.6151
R1046 B.n377 B.n144 10.6151
R1047 B.n378 B.n377 10.6151
R1048 B.n379 B.n378 10.6151
R1049 B.n379 B.n142 10.6151
R1050 B.n383 B.n142 10.6151
R1051 B.n384 B.n383 10.6151
R1052 B.n385 B.n384 10.6151
R1053 B.n385 B.n140 10.6151
R1054 B.n389 B.n140 10.6151
R1055 B.n390 B.n389 10.6151
R1056 B.n391 B.n390 10.6151
R1057 B.n391 B.n138 10.6151
R1058 B.n395 B.n138 10.6151
R1059 B.n396 B.n395 10.6151
R1060 B.n397 B.n396 10.6151
R1061 B.n397 B.n136 10.6151
R1062 B.n401 B.n136 10.6151
R1063 B.n402 B.n401 10.6151
R1064 B.n403 B.n402 10.6151
R1065 B.n294 B.n293 10.6151
R1066 B.n293 B.n176 10.6151
R1067 B.n289 B.n176 10.6151
R1068 B.n289 B.n288 10.6151
R1069 B.n288 B.n287 10.6151
R1070 B.n287 B.n178 10.6151
R1071 B.n283 B.n178 10.6151
R1072 B.n283 B.n282 10.6151
R1073 B.n282 B.n281 10.6151
R1074 B.n281 B.n180 10.6151
R1075 B.n277 B.n180 10.6151
R1076 B.n277 B.n276 10.6151
R1077 B.n276 B.n275 10.6151
R1078 B.n275 B.n182 10.6151
R1079 B.n271 B.n182 10.6151
R1080 B.n271 B.n270 10.6151
R1081 B.n270 B.n269 10.6151
R1082 B.n269 B.n184 10.6151
R1083 B.n265 B.n184 10.6151
R1084 B.n265 B.n264 10.6151
R1085 B.n264 B.n263 10.6151
R1086 B.n263 B.n186 10.6151
R1087 B.n259 B.n186 10.6151
R1088 B.n259 B.n258 10.6151
R1089 B.n258 B.n257 10.6151
R1090 B.n257 B.n188 10.6151
R1091 B.n253 B.n188 10.6151
R1092 B.n253 B.n252 10.6151
R1093 B.n252 B.n251 10.6151
R1094 B.n251 B.n190 10.6151
R1095 B.n247 B.n190 10.6151
R1096 B.n247 B.n246 10.6151
R1097 B.n246 B.n245 10.6151
R1098 B.n245 B.n192 10.6151
R1099 B.n241 B.n192 10.6151
R1100 B.n241 B.n240 10.6151
R1101 B.n240 B.n239 10.6151
R1102 B.n239 B.n194 10.6151
R1103 B.n235 B.n194 10.6151
R1104 B.n235 B.n234 10.6151
R1105 B.n234 B.n233 10.6151
R1106 B.n233 B.n196 10.6151
R1107 B.n229 B.n196 10.6151
R1108 B.n229 B.n228 10.6151
R1109 B.n228 B.n227 10.6151
R1110 B.n227 B.n198 10.6151
R1111 B.n223 B.n198 10.6151
R1112 B.n223 B.n222 10.6151
R1113 B.n222 B.n221 10.6151
R1114 B.n221 B.n200 10.6151
R1115 B.n217 B.n200 10.6151
R1116 B.n217 B.n216 10.6151
R1117 B.n216 B.n215 10.6151
R1118 B.n215 B.n202 10.6151
R1119 B.n211 B.n202 10.6151
R1120 B.n211 B.n210 10.6151
R1121 B.n210 B.n209 10.6151
R1122 B.n209 B.n204 10.6151
R1123 B.n205 B.n204 10.6151
R1124 B.n205 B.n0 10.6151
R1125 B.n787 B.n1 10.6151
R1126 B.n787 B.n786 10.6151
R1127 B.n786 B.n785 10.6151
R1128 B.n785 B.n4 10.6151
R1129 B.n781 B.n4 10.6151
R1130 B.n781 B.n780 10.6151
R1131 B.n780 B.n779 10.6151
R1132 B.n779 B.n6 10.6151
R1133 B.n775 B.n6 10.6151
R1134 B.n775 B.n774 10.6151
R1135 B.n774 B.n773 10.6151
R1136 B.n773 B.n8 10.6151
R1137 B.n769 B.n8 10.6151
R1138 B.n769 B.n768 10.6151
R1139 B.n768 B.n767 10.6151
R1140 B.n767 B.n10 10.6151
R1141 B.n763 B.n10 10.6151
R1142 B.n763 B.n762 10.6151
R1143 B.n762 B.n761 10.6151
R1144 B.n761 B.n12 10.6151
R1145 B.n757 B.n12 10.6151
R1146 B.n757 B.n756 10.6151
R1147 B.n756 B.n755 10.6151
R1148 B.n755 B.n14 10.6151
R1149 B.n751 B.n14 10.6151
R1150 B.n751 B.n750 10.6151
R1151 B.n750 B.n749 10.6151
R1152 B.n749 B.n16 10.6151
R1153 B.n745 B.n16 10.6151
R1154 B.n745 B.n744 10.6151
R1155 B.n744 B.n743 10.6151
R1156 B.n743 B.n18 10.6151
R1157 B.n739 B.n18 10.6151
R1158 B.n739 B.n738 10.6151
R1159 B.n738 B.n737 10.6151
R1160 B.n737 B.n20 10.6151
R1161 B.n733 B.n20 10.6151
R1162 B.n733 B.n732 10.6151
R1163 B.n732 B.n731 10.6151
R1164 B.n731 B.n22 10.6151
R1165 B.n727 B.n22 10.6151
R1166 B.n727 B.n726 10.6151
R1167 B.n726 B.n725 10.6151
R1168 B.n725 B.n24 10.6151
R1169 B.n721 B.n24 10.6151
R1170 B.n721 B.n720 10.6151
R1171 B.n720 B.n719 10.6151
R1172 B.n719 B.n26 10.6151
R1173 B.n715 B.n26 10.6151
R1174 B.n715 B.n714 10.6151
R1175 B.n714 B.n713 10.6151
R1176 B.n713 B.n28 10.6151
R1177 B.n709 B.n28 10.6151
R1178 B.n709 B.n708 10.6151
R1179 B.n708 B.n707 10.6151
R1180 B.n707 B.n30 10.6151
R1181 B.n703 B.n30 10.6151
R1182 B.n703 B.n702 10.6151
R1183 B.n702 B.n701 10.6151
R1184 B.n701 B.n32 10.6151
R1185 B.n653 B.n50 9.36635
R1186 B.n636 B.n635 9.36635
R1187 B.n342 B.n341 9.36635
R1188 B.n359 B.n152 9.36635
R1189 B.n791 B.n0 2.81026
R1190 B.n791 B.n1 2.81026
R1191 B.n650 B.n50 1.24928
R1192 B.n637 B.n636 1.24928
R1193 B.n343 B.n342 1.24928
R1194 B.n356 B.n152 1.24928
R1195 VN.n83 VN.n43 161.3
R1196 VN.n82 VN.n81 161.3
R1197 VN.n80 VN.n44 161.3
R1198 VN.n79 VN.n78 161.3
R1199 VN.n77 VN.n45 161.3
R1200 VN.n76 VN.n75 161.3
R1201 VN.n74 VN.n73 161.3
R1202 VN.n72 VN.n47 161.3
R1203 VN.n71 VN.n70 161.3
R1204 VN.n69 VN.n48 161.3
R1205 VN.n68 VN.n67 161.3
R1206 VN.n66 VN.n49 161.3
R1207 VN.n65 VN.n64 161.3
R1208 VN.n63 VN.n50 161.3
R1209 VN.n62 VN.n61 161.3
R1210 VN.n60 VN.n51 161.3
R1211 VN.n59 VN.n58 161.3
R1212 VN.n57 VN.n52 161.3
R1213 VN.n56 VN.n55 161.3
R1214 VN.n40 VN.n0 161.3
R1215 VN.n39 VN.n38 161.3
R1216 VN.n37 VN.n1 161.3
R1217 VN.n36 VN.n35 161.3
R1218 VN.n34 VN.n2 161.3
R1219 VN.n33 VN.n32 161.3
R1220 VN.n31 VN.n30 161.3
R1221 VN.n29 VN.n4 161.3
R1222 VN.n28 VN.n27 161.3
R1223 VN.n26 VN.n5 161.3
R1224 VN.n25 VN.n24 161.3
R1225 VN.n23 VN.n6 161.3
R1226 VN.n22 VN.n21 161.3
R1227 VN.n20 VN.n7 161.3
R1228 VN.n19 VN.n18 161.3
R1229 VN.n17 VN.n8 161.3
R1230 VN.n16 VN.n15 161.3
R1231 VN.n14 VN.n9 161.3
R1232 VN.n13 VN.n12 161.3
R1233 VN.n42 VN.n41 109.924
R1234 VN.n85 VN.n84 109.924
R1235 VN.n10 VN.t8 107.171
R1236 VN.n53 VN.t3 107.171
R1237 VN.n22 VN.t2 76.7968
R1238 VN.n11 VN.t6 76.7968
R1239 VN.n3 VN.t0 76.7968
R1240 VN.n41 VN.t7 76.7968
R1241 VN.n65 VN.t5 76.7968
R1242 VN.n54 VN.t9 76.7968
R1243 VN.n46 VN.t1 76.7968
R1244 VN.n84 VN.t4 76.7968
R1245 VN.n11 VN.n10 73.1566
R1246 VN.n54 VN.n53 73.1566
R1247 VN VN.n85 51.108
R1248 VN.n35 VN.n1 42.0302
R1249 VN.n78 VN.n44 42.0302
R1250 VN.n17 VN.n16 41.0614
R1251 VN.n28 VN.n5 41.0614
R1252 VN.n60 VN.n59 41.0614
R1253 VN.n71 VN.n48 41.0614
R1254 VN.n18 VN.n17 40.0926
R1255 VN.n24 VN.n5 40.0926
R1256 VN.n61 VN.n60 40.0926
R1257 VN.n67 VN.n48 40.0926
R1258 VN.n35 VN.n34 39.1239
R1259 VN.n78 VN.n77 39.1239
R1260 VN.n12 VN.n9 24.5923
R1261 VN.n16 VN.n9 24.5923
R1262 VN.n18 VN.n7 24.5923
R1263 VN.n22 VN.n7 24.5923
R1264 VN.n23 VN.n22 24.5923
R1265 VN.n24 VN.n23 24.5923
R1266 VN.n29 VN.n28 24.5923
R1267 VN.n30 VN.n29 24.5923
R1268 VN.n34 VN.n33 24.5923
R1269 VN.n39 VN.n1 24.5923
R1270 VN.n40 VN.n39 24.5923
R1271 VN.n59 VN.n52 24.5923
R1272 VN.n55 VN.n52 24.5923
R1273 VN.n67 VN.n66 24.5923
R1274 VN.n66 VN.n65 24.5923
R1275 VN.n65 VN.n50 24.5923
R1276 VN.n61 VN.n50 24.5923
R1277 VN.n77 VN.n76 24.5923
R1278 VN.n73 VN.n72 24.5923
R1279 VN.n72 VN.n71 24.5923
R1280 VN.n83 VN.n82 24.5923
R1281 VN.n82 VN.n44 24.5923
R1282 VN.n33 VN.n3 24.1005
R1283 VN.n76 VN.n46 24.1005
R1284 VN.n56 VN.n53 7.42269
R1285 VN.n13 VN.n10 7.42269
R1286 VN.n41 VN.n40 0.984173
R1287 VN.n84 VN.n83 0.984173
R1288 VN.n12 VN.n11 0.492337
R1289 VN.n30 VN.n3 0.492337
R1290 VN.n55 VN.n54 0.492337
R1291 VN.n73 VN.n46 0.492337
R1292 VN.n85 VN.n43 0.278335
R1293 VN.n42 VN.n0 0.278335
R1294 VN.n81 VN.n43 0.189894
R1295 VN.n81 VN.n80 0.189894
R1296 VN.n80 VN.n79 0.189894
R1297 VN.n79 VN.n45 0.189894
R1298 VN.n75 VN.n45 0.189894
R1299 VN.n75 VN.n74 0.189894
R1300 VN.n74 VN.n47 0.189894
R1301 VN.n70 VN.n47 0.189894
R1302 VN.n70 VN.n69 0.189894
R1303 VN.n69 VN.n68 0.189894
R1304 VN.n68 VN.n49 0.189894
R1305 VN.n64 VN.n49 0.189894
R1306 VN.n64 VN.n63 0.189894
R1307 VN.n63 VN.n62 0.189894
R1308 VN.n62 VN.n51 0.189894
R1309 VN.n58 VN.n51 0.189894
R1310 VN.n58 VN.n57 0.189894
R1311 VN.n57 VN.n56 0.189894
R1312 VN.n14 VN.n13 0.189894
R1313 VN.n15 VN.n14 0.189894
R1314 VN.n15 VN.n8 0.189894
R1315 VN.n19 VN.n8 0.189894
R1316 VN.n20 VN.n19 0.189894
R1317 VN.n21 VN.n20 0.189894
R1318 VN.n21 VN.n6 0.189894
R1319 VN.n25 VN.n6 0.189894
R1320 VN.n26 VN.n25 0.189894
R1321 VN.n27 VN.n26 0.189894
R1322 VN.n27 VN.n4 0.189894
R1323 VN.n31 VN.n4 0.189894
R1324 VN.n32 VN.n31 0.189894
R1325 VN.n32 VN.n2 0.189894
R1326 VN.n36 VN.n2 0.189894
R1327 VN.n37 VN.n36 0.189894
R1328 VN.n38 VN.n37 0.189894
R1329 VN.n38 VN.n0 0.189894
R1330 VN VN.n42 0.153485
R1331 VDD2.n89 VDD2.n49 756.745
R1332 VDD2.n40 VDD2.n0 756.745
R1333 VDD2.n90 VDD2.n89 585
R1334 VDD2.n88 VDD2.n87 585
R1335 VDD2.n86 VDD2.n52 585
R1336 VDD2.n56 VDD2.n53 585
R1337 VDD2.n81 VDD2.n80 585
R1338 VDD2.n79 VDD2.n78 585
R1339 VDD2.n58 VDD2.n57 585
R1340 VDD2.n73 VDD2.n72 585
R1341 VDD2.n71 VDD2.n70 585
R1342 VDD2.n62 VDD2.n61 585
R1343 VDD2.n65 VDD2.n64 585
R1344 VDD2.n15 VDD2.n14 585
R1345 VDD2.n12 VDD2.n11 585
R1346 VDD2.n21 VDD2.n20 585
R1347 VDD2.n23 VDD2.n22 585
R1348 VDD2.n8 VDD2.n7 585
R1349 VDD2.n29 VDD2.n28 585
R1350 VDD2.n32 VDD2.n31 585
R1351 VDD2.n30 VDD2.n4 585
R1352 VDD2.n37 VDD2.n3 585
R1353 VDD2.n39 VDD2.n38 585
R1354 VDD2.n41 VDD2.n40 585
R1355 VDD2.t6 VDD2.n63 329.039
R1356 VDD2.t4 VDD2.n13 329.038
R1357 VDD2.n89 VDD2.n88 171.744
R1358 VDD2.n88 VDD2.n52 171.744
R1359 VDD2.n56 VDD2.n52 171.744
R1360 VDD2.n80 VDD2.n56 171.744
R1361 VDD2.n80 VDD2.n79 171.744
R1362 VDD2.n79 VDD2.n57 171.744
R1363 VDD2.n72 VDD2.n57 171.744
R1364 VDD2.n72 VDD2.n71 171.744
R1365 VDD2.n71 VDD2.n61 171.744
R1366 VDD2.n64 VDD2.n61 171.744
R1367 VDD2.n14 VDD2.n11 171.744
R1368 VDD2.n21 VDD2.n11 171.744
R1369 VDD2.n22 VDD2.n21 171.744
R1370 VDD2.n22 VDD2.n7 171.744
R1371 VDD2.n29 VDD2.n7 171.744
R1372 VDD2.n31 VDD2.n29 171.744
R1373 VDD2.n31 VDD2.n30 171.744
R1374 VDD2.n30 VDD2.n3 171.744
R1375 VDD2.n39 VDD2.n3 171.744
R1376 VDD2.n40 VDD2.n39 171.744
R1377 VDD2.n64 VDD2.t6 85.8723
R1378 VDD2.n14 VDD2.t4 85.8723
R1379 VDD2.n48 VDD2.n47 82.5828
R1380 VDD2 VDD2.n97 82.5799
R1381 VDD2.n96 VDD2.n95 80.6922
R1382 VDD2.n46 VDD2.n45 80.692
R1383 VDD2.n46 VDD2.n44 51.8468
R1384 VDD2.n94 VDD2.n93 49.252
R1385 VDD2.n94 VDD2.n48 43.4028
R1386 VDD2.n87 VDD2.n86 13.1884
R1387 VDD2.n38 VDD2.n37 13.1884
R1388 VDD2.n90 VDD2.n51 12.8005
R1389 VDD2.n85 VDD2.n53 12.8005
R1390 VDD2.n36 VDD2.n4 12.8005
R1391 VDD2.n41 VDD2.n2 12.8005
R1392 VDD2.n91 VDD2.n49 12.0247
R1393 VDD2.n82 VDD2.n81 12.0247
R1394 VDD2.n33 VDD2.n32 12.0247
R1395 VDD2.n42 VDD2.n0 12.0247
R1396 VDD2.n78 VDD2.n55 11.249
R1397 VDD2.n28 VDD2.n6 11.249
R1398 VDD2.n65 VDD2.n63 10.7239
R1399 VDD2.n15 VDD2.n13 10.7239
R1400 VDD2.n77 VDD2.n58 10.4732
R1401 VDD2.n27 VDD2.n8 10.4732
R1402 VDD2.n74 VDD2.n73 9.69747
R1403 VDD2.n24 VDD2.n23 9.69747
R1404 VDD2.n93 VDD2.n92 9.45567
R1405 VDD2.n44 VDD2.n43 9.45567
R1406 VDD2.n67 VDD2.n66 9.3005
R1407 VDD2.n69 VDD2.n68 9.3005
R1408 VDD2.n60 VDD2.n59 9.3005
R1409 VDD2.n75 VDD2.n74 9.3005
R1410 VDD2.n77 VDD2.n76 9.3005
R1411 VDD2.n55 VDD2.n54 9.3005
R1412 VDD2.n83 VDD2.n82 9.3005
R1413 VDD2.n85 VDD2.n84 9.3005
R1414 VDD2.n92 VDD2.n91 9.3005
R1415 VDD2.n51 VDD2.n50 9.3005
R1416 VDD2.n43 VDD2.n42 9.3005
R1417 VDD2.n2 VDD2.n1 9.3005
R1418 VDD2.n17 VDD2.n16 9.3005
R1419 VDD2.n19 VDD2.n18 9.3005
R1420 VDD2.n10 VDD2.n9 9.3005
R1421 VDD2.n25 VDD2.n24 9.3005
R1422 VDD2.n27 VDD2.n26 9.3005
R1423 VDD2.n6 VDD2.n5 9.3005
R1424 VDD2.n34 VDD2.n33 9.3005
R1425 VDD2.n36 VDD2.n35 9.3005
R1426 VDD2.n70 VDD2.n60 8.92171
R1427 VDD2.n20 VDD2.n10 8.92171
R1428 VDD2.n69 VDD2.n62 8.14595
R1429 VDD2.n19 VDD2.n12 8.14595
R1430 VDD2.n66 VDD2.n65 7.3702
R1431 VDD2.n16 VDD2.n15 7.3702
R1432 VDD2.n66 VDD2.n62 5.81868
R1433 VDD2.n16 VDD2.n12 5.81868
R1434 VDD2.n70 VDD2.n69 5.04292
R1435 VDD2.n20 VDD2.n19 5.04292
R1436 VDD2.n73 VDD2.n60 4.26717
R1437 VDD2.n23 VDD2.n10 4.26717
R1438 VDD2.n97 VDD2.t2 3.80671
R1439 VDD2.n97 VDD2.t1 3.80671
R1440 VDD2.n95 VDD2.t9 3.80671
R1441 VDD2.n95 VDD2.t3 3.80671
R1442 VDD2.n47 VDD2.t5 3.80671
R1443 VDD2.n47 VDD2.t8 3.80671
R1444 VDD2.n45 VDD2.t0 3.80671
R1445 VDD2.n45 VDD2.t7 3.80671
R1446 VDD2.n74 VDD2.n58 3.49141
R1447 VDD2.n24 VDD2.n8 3.49141
R1448 VDD2.n78 VDD2.n77 2.71565
R1449 VDD2.n28 VDD2.n27 2.71565
R1450 VDD2.n96 VDD2.n94 2.59533
R1451 VDD2.n67 VDD2.n63 2.41285
R1452 VDD2.n17 VDD2.n13 2.41285
R1453 VDD2.n93 VDD2.n49 1.93989
R1454 VDD2.n81 VDD2.n55 1.93989
R1455 VDD2.n32 VDD2.n6 1.93989
R1456 VDD2.n44 VDD2.n0 1.93989
R1457 VDD2.n91 VDD2.n90 1.16414
R1458 VDD2.n82 VDD2.n53 1.16414
R1459 VDD2.n33 VDD2.n4 1.16414
R1460 VDD2.n42 VDD2.n41 1.16414
R1461 VDD2 VDD2.n96 0.707397
R1462 VDD2.n48 VDD2.n46 0.593861
R1463 VDD2.n87 VDD2.n51 0.388379
R1464 VDD2.n86 VDD2.n85 0.388379
R1465 VDD2.n37 VDD2.n36 0.388379
R1466 VDD2.n38 VDD2.n2 0.388379
R1467 VDD2.n92 VDD2.n50 0.155672
R1468 VDD2.n84 VDD2.n50 0.155672
R1469 VDD2.n84 VDD2.n83 0.155672
R1470 VDD2.n83 VDD2.n54 0.155672
R1471 VDD2.n76 VDD2.n54 0.155672
R1472 VDD2.n76 VDD2.n75 0.155672
R1473 VDD2.n75 VDD2.n59 0.155672
R1474 VDD2.n68 VDD2.n59 0.155672
R1475 VDD2.n68 VDD2.n67 0.155672
R1476 VDD2.n18 VDD2.n17 0.155672
R1477 VDD2.n18 VDD2.n9 0.155672
R1478 VDD2.n25 VDD2.n9 0.155672
R1479 VDD2.n26 VDD2.n25 0.155672
R1480 VDD2.n26 VDD2.n5 0.155672
R1481 VDD2.n34 VDD2.n5 0.155672
R1482 VDD2.n35 VDD2.n34 0.155672
R1483 VDD2.n35 VDD2.n1 0.155672
R1484 VDD2.n43 VDD2.n1 0.155672
R1485 VTAIL.n192 VTAIL.n152 756.745
R1486 VTAIL.n42 VTAIL.n2 756.745
R1487 VTAIL.n146 VTAIL.n106 756.745
R1488 VTAIL.n96 VTAIL.n56 756.745
R1489 VTAIL.n167 VTAIL.n166 585
R1490 VTAIL.n164 VTAIL.n163 585
R1491 VTAIL.n173 VTAIL.n172 585
R1492 VTAIL.n175 VTAIL.n174 585
R1493 VTAIL.n160 VTAIL.n159 585
R1494 VTAIL.n181 VTAIL.n180 585
R1495 VTAIL.n184 VTAIL.n183 585
R1496 VTAIL.n182 VTAIL.n156 585
R1497 VTAIL.n189 VTAIL.n155 585
R1498 VTAIL.n191 VTAIL.n190 585
R1499 VTAIL.n193 VTAIL.n192 585
R1500 VTAIL.n17 VTAIL.n16 585
R1501 VTAIL.n14 VTAIL.n13 585
R1502 VTAIL.n23 VTAIL.n22 585
R1503 VTAIL.n25 VTAIL.n24 585
R1504 VTAIL.n10 VTAIL.n9 585
R1505 VTAIL.n31 VTAIL.n30 585
R1506 VTAIL.n34 VTAIL.n33 585
R1507 VTAIL.n32 VTAIL.n6 585
R1508 VTAIL.n39 VTAIL.n5 585
R1509 VTAIL.n41 VTAIL.n40 585
R1510 VTAIL.n43 VTAIL.n42 585
R1511 VTAIL.n147 VTAIL.n146 585
R1512 VTAIL.n145 VTAIL.n144 585
R1513 VTAIL.n143 VTAIL.n109 585
R1514 VTAIL.n113 VTAIL.n110 585
R1515 VTAIL.n138 VTAIL.n137 585
R1516 VTAIL.n136 VTAIL.n135 585
R1517 VTAIL.n115 VTAIL.n114 585
R1518 VTAIL.n130 VTAIL.n129 585
R1519 VTAIL.n128 VTAIL.n127 585
R1520 VTAIL.n119 VTAIL.n118 585
R1521 VTAIL.n122 VTAIL.n121 585
R1522 VTAIL.n97 VTAIL.n96 585
R1523 VTAIL.n95 VTAIL.n94 585
R1524 VTAIL.n93 VTAIL.n59 585
R1525 VTAIL.n63 VTAIL.n60 585
R1526 VTAIL.n88 VTAIL.n87 585
R1527 VTAIL.n86 VTAIL.n85 585
R1528 VTAIL.n65 VTAIL.n64 585
R1529 VTAIL.n80 VTAIL.n79 585
R1530 VTAIL.n78 VTAIL.n77 585
R1531 VTAIL.n69 VTAIL.n68 585
R1532 VTAIL.n72 VTAIL.n71 585
R1533 VTAIL.t1 VTAIL.n120 329.039
R1534 VTAIL.t16 VTAIL.n70 329.039
R1535 VTAIL.t12 VTAIL.n165 329.038
R1536 VTAIL.t6 VTAIL.n15 329.038
R1537 VTAIL.n166 VTAIL.n163 171.744
R1538 VTAIL.n173 VTAIL.n163 171.744
R1539 VTAIL.n174 VTAIL.n173 171.744
R1540 VTAIL.n174 VTAIL.n159 171.744
R1541 VTAIL.n181 VTAIL.n159 171.744
R1542 VTAIL.n183 VTAIL.n181 171.744
R1543 VTAIL.n183 VTAIL.n182 171.744
R1544 VTAIL.n182 VTAIL.n155 171.744
R1545 VTAIL.n191 VTAIL.n155 171.744
R1546 VTAIL.n192 VTAIL.n191 171.744
R1547 VTAIL.n16 VTAIL.n13 171.744
R1548 VTAIL.n23 VTAIL.n13 171.744
R1549 VTAIL.n24 VTAIL.n23 171.744
R1550 VTAIL.n24 VTAIL.n9 171.744
R1551 VTAIL.n31 VTAIL.n9 171.744
R1552 VTAIL.n33 VTAIL.n31 171.744
R1553 VTAIL.n33 VTAIL.n32 171.744
R1554 VTAIL.n32 VTAIL.n5 171.744
R1555 VTAIL.n41 VTAIL.n5 171.744
R1556 VTAIL.n42 VTAIL.n41 171.744
R1557 VTAIL.n146 VTAIL.n145 171.744
R1558 VTAIL.n145 VTAIL.n109 171.744
R1559 VTAIL.n113 VTAIL.n109 171.744
R1560 VTAIL.n137 VTAIL.n113 171.744
R1561 VTAIL.n137 VTAIL.n136 171.744
R1562 VTAIL.n136 VTAIL.n114 171.744
R1563 VTAIL.n129 VTAIL.n114 171.744
R1564 VTAIL.n129 VTAIL.n128 171.744
R1565 VTAIL.n128 VTAIL.n118 171.744
R1566 VTAIL.n121 VTAIL.n118 171.744
R1567 VTAIL.n96 VTAIL.n95 171.744
R1568 VTAIL.n95 VTAIL.n59 171.744
R1569 VTAIL.n63 VTAIL.n59 171.744
R1570 VTAIL.n87 VTAIL.n63 171.744
R1571 VTAIL.n87 VTAIL.n86 171.744
R1572 VTAIL.n86 VTAIL.n64 171.744
R1573 VTAIL.n79 VTAIL.n64 171.744
R1574 VTAIL.n79 VTAIL.n78 171.744
R1575 VTAIL.n78 VTAIL.n68 171.744
R1576 VTAIL.n71 VTAIL.n68 171.744
R1577 VTAIL.n166 VTAIL.t12 85.8723
R1578 VTAIL.n16 VTAIL.t6 85.8723
R1579 VTAIL.n121 VTAIL.t1 85.8723
R1580 VTAIL.n71 VTAIL.t16 85.8723
R1581 VTAIL.n105 VTAIL.n104 64.0134
R1582 VTAIL.n103 VTAIL.n102 64.0134
R1583 VTAIL.n55 VTAIL.n54 64.0134
R1584 VTAIL.n53 VTAIL.n52 64.0134
R1585 VTAIL.n199 VTAIL.n198 64.0132
R1586 VTAIL.n1 VTAIL.n0 64.0132
R1587 VTAIL.n49 VTAIL.n48 64.0132
R1588 VTAIL.n51 VTAIL.n50 64.0132
R1589 VTAIL.n197 VTAIL.n196 32.5732
R1590 VTAIL.n47 VTAIL.n46 32.5732
R1591 VTAIL.n151 VTAIL.n150 32.5732
R1592 VTAIL.n101 VTAIL.n100 32.5732
R1593 VTAIL.n53 VTAIL.n51 24.9186
R1594 VTAIL.n197 VTAIL.n151 22.3238
R1595 VTAIL.n190 VTAIL.n189 13.1884
R1596 VTAIL.n40 VTAIL.n39 13.1884
R1597 VTAIL.n144 VTAIL.n143 13.1884
R1598 VTAIL.n94 VTAIL.n93 13.1884
R1599 VTAIL.n188 VTAIL.n156 12.8005
R1600 VTAIL.n193 VTAIL.n154 12.8005
R1601 VTAIL.n38 VTAIL.n6 12.8005
R1602 VTAIL.n43 VTAIL.n4 12.8005
R1603 VTAIL.n147 VTAIL.n108 12.8005
R1604 VTAIL.n142 VTAIL.n110 12.8005
R1605 VTAIL.n97 VTAIL.n58 12.8005
R1606 VTAIL.n92 VTAIL.n60 12.8005
R1607 VTAIL.n185 VTAIL.n184 12.0247
R1608 VTAIL.n194 VTAIL.n152 12.0247
R1609 VTAIL.n35 VTAIL.n34 12.0247
R1610 VTAIL.n44 VTAIL.n2 12.0247
R1611 VTAIL.n148 VTAIL.n106 12.0247
R1612 VTAIL.n139 VTAIL.n138 12.0247
R1613 VTAIL.n98 VTAIL.n56 12.0247
R1614 VTAIL.n89 VTAIL.n88 12.0247
R1615 VTAIL.n180 VTAIL.n158 11.249
R1616 VTAIL.n30 VTAIL.n8 11.249
R1617 VTAIL.n135 VTAIL.n112 11.249
R1618 VTAIL.n85 VTAIL.n62 11.249
R1619 VTAIL.n167 VTAIL.n165 10.7239
R1620 VTAIL.n17 VTAIL.n15 10.7239
R1621 VTAIL.n122 VTAIL.n120 10.7239
R1622 VTAIL.n72 VTAIL.n70 10.7239
R1623 VTAIL.n179 VTAIL.n160 10.4732
R1624 VTAIL.n29 VTAIL.n10 10.4732
R1625 VTAIL.n134 VTAIL.n115 10.4732
R1626 VTAIL.n84 VTAIL.n65 10.4732
R1627 VTAIL.n176 VTAIL.n175 9.69747
R1628 VTAIL.n26 VTAIL.n25 9.69747
R1629 VTAIL.n131 VTAIL.n130 9.69747
R1630 VTAIL.n81 VTAIL.n80 9.69747
R1631 VTAIL.n196 VTAIL.n195 9.45567
R1632 VTAIL.n46 VTAIL.n45 9.45567
R1633 VTAIL.n150 VTAIL.n149 9.45567
R1634 VTAIL.n100 VTAIL.n99 9.45567
R1635 VTAIL.n195 VTAIL.n194 9.3005
R1636 VTAIL.n154 VTAIL.n153 9.3005
R1637 VTAIL.n169 VTAIL.n168 9.3005
R1638 VTAIL.n171 VTAIL.n170 9.3005
R1639 VTAIL.n162 VTAIL.n161 9.3005
R1640 VTAIL.n177 VTAIL.n176 9.3005
R1641 VTAIL.n179 VTAIL.n178 9.3005
R1642 VTAIL.n158 VTAIL.n157 9.3005
R1643 VTAIL.n186 VTAIL.n185 9.3005
R1644 VTAIL.n188 VTAIL.n187 9.3005
R1645 VTAIL.n45 VTAIL.n44 9.3005
R1646 VTAIL.n4 VTAIL.n3 9.3005
R1647 VTAIL.n19 VTAIL.n18 9.3005
R1648 VTAIL.n21 VTAIL.n20 9.3005
R1649 VTAIL.n12 VTAIL.n11 9.3005
R1650 VTAIL.n27 VTAIL.n26 9.3005
R1651 VTAIL.n29 VTAIL.n28 9.3005
R1652 VTAIL.n8 VTAIL.n7 9.3005
R1653 VTAIL.n36 VTAIL.n35 9.3005
R1654 VTAIL.n38 VTAIL.n37 9.3005
R1655 VTAIL.n124 VTAIL.n123 9.3005
R1656 VTAIL.n126 VTAIL.n125 9.3005
R1657 VTAIL.n117 VTAIL.n116 9.3005
R1658 VTAIL.n132 VTAIL.n131 9.3005
R1659 VTAIL.n134 VTAIL.n133 9.3005
R1660 VTAIL.n112 VTAIL.n111 9.3005
R1661 VTAIL.n140 VTAIL.n139 9.3005
R1662 VTAIL.n142 VTAIL.n141 9.3005
R1663 VTAIL.n149 VTAIL.n148 9.3005
R1664 VTAIL.n108 VTAIL.n107 9.3005
R1665 VTAIL.n74 VTAIL.n73 9.3005
R1666 VTAIL.n76 VTAIL.n75 9.3005
R1667 VTAIL.n67 VTAIL.n66 9.3005
R1668 VTAIL.n82 VTAIL.n81 9.3005
R1669 VTAIL.n84 VTAIL.n83 9.3005
R1670 VTAIL.n62 VTAIL.n61 9.3005
R1671 VTAIL.n90 VTAIL.n89 9.3005
R1672 VTAIL.n92 VTAIL.n91 9.3005
R1673 VTAIL.n99 VTAIL.n98 9.3005
R1674 VTAIL.n58 VTAIL.n57 9.3005
R1675 VTAIL.n172 VTAIL.n162 8.92171
R1676 VTAIL.n22 VTAIL.n12 8.92171
R1677 VTAIL.n127 VTAIL.n117 8.92171
R1678 VTAIL.n77 VTAIL.n67 8.92171
R1679 VTAIL.n171 VTAIL.n164 8.14595
R1680 VTAIL.n21 VTAIL.n14 8.14595
R1681 VTAIL.n126 VTAIL.n119 8.14595
R1682 VTAIL.n76 VTAIL.n69 8.14595
R1683 VTAIL.n168 VTAIL.n167 7.3702
R1684 VTAIL.n18 VTAIL.n17 7.3702
R1685 VTAIL.n123 VTAIL.n122 7.3702
R1686 VTAIL.n73 VTAIL.n72 7.3702
R1687 VTAIL.n168 VTAIL.n164 5.81868
R1688 VTAIL.n18 VTAIL.n14 5.81868
R1689 VTAIL.n123 VTAIL.n119 5.81868
R1690 VTAIL.n73 VTAIL.n69 5.81868
R1691 VTAIL.n172 VTAIL.n171 5.04292
R1692 VTAIL.n22 VTAIL.n21 5.04292
R1693 VTAIL.n127 VTAIL.n126 5.04292
R1694 VTAIL.n77 VTAIL.n76 5.04292
R1695 VTAIL.n175 VTAIL.n162 4.26717
R1696 VTAIL.n25 VTAIL.n12 4.26717
R1697 VTAIL.n130 VTAIL.n117 4.26717
R1698 VTAIL.n80 VTAIL.n67 4.26717
R1699 VTAIL.n198 VTAIL.t17 3.80671
R1700 VTAIL.n198 VTAIL.t19 3.80671
R1701 VTAIL.n0 VTAIL.t11 3.80671
R1702 VTAIL.n0 VTAIL.t13 3.80671
R1703 VTAIL.n48 VTAIL.t3 3.80671
R1704 VTAIL.n48 VTAIL.t5 3.80671
R1705 VTAIL.n50 VTAIL.t8 3.80671
R1706 VTAIL.n50 VTAIL.t7 3.80671
R1707 VTAIL.n104 VTAIL.t2 3.80671
R1708 VTAIL.n104 VTAIL.t0 3.80671
R1709 VTAIL.n102 VTAIL.t4 3.80671
R1710 VTAIL.n102 VTAIL.t9 3.80671
R1711 VTAIL.n54 VTAIL.t14 3.80671
R1712 VTAIL.n54 VTAIL.t10 3.80671
R1713 VTAIL.n52 VTAIL.t15 3.80671
R1714 VTAIL.n52 VTAIL.t18 3.80671
R1715 VTAIL.n176 VTAIL.n160 3.49141
R1716 VTAIL.n26 VTAIL.n10 3.49141
R1717 VTAIL.n131 VTAIL.n115 3.49141
R1718 VTAIL.n81 VTAIL.n65 3.49141
R1719 VTAIL.n180 VTAIL.n179 2.71565
R1720 VTAIL.n30 VTAIL.n29 2.71565
R1721 VTAIL.n135 VTAIL.n134 2.71565
R1722 VTAIL.n85 VTAIL.n84 2.71565
R1723 VTAIL.n55 VTAIL.n53 2.59533
R1724 VTAIL.n101 VTAIL.n55 2.59533
R1725 VTAIL.n105 VTAIL.n103 2.59533
R1726 VTAIL.n151 VTAIL.n105 2.59533
R1727 VTAIL.n51 VTAIL.n49 2.59533
R1728 VTAIL.n49 VTAIL.n47 2.59533
R1729 VTAIL.n199 VTAIL.n197 2.59533
R1730 VTAIL.n169 VTAIL.n165 2.41285
R1731 VTAIL.n19 VTAIL.n15 2.41285
R1732 VTAIL.n124 VTAIL.n120 2.41285
R1733 VTAIL.n74 VTAIL.n70 2.41285
R1734 VTAIL VTAIL.n1 2.00481
R1735 VTAIL.n184 VTAIL.n158 1.93989
R1736 VTAIL.n196 VTAIL.n152 1.93989
R1737 VTAIL.n34 VTAIL.n8 1.93989
R1738 VTAIL.n46 VTAIL.n2 1.93989
R1739 VTAIL.n150 VTAIL.n106 1.93989
R1740 VTAIL.n138 VTAIL.n112 1.93989
R1741 VTAIL.n100 VTAIL.n56 1.93989
R1742 VTAIL.n88 VTAIL.n62 1.93989
R1743 VTAIL.n103 VTAIL.n101 1.76774
R1744 VTAIL.n47 VTAIL.n1 1.76774
R1745 VTAIL.n185 VTAIL.n156 1.16414
R1746 VTAIL.n194 VTAIL.n193 1.16414
R1747 VTAIL.n35 VTAIL.n6 1.16414
R1748 VTAIL.n44 VTAIL.n43 1.16414
R1749 VTAIL.n148 VTAIL.n147 1.16414
R1750 VTAIL.n139 VTAIL.n110 1.16414
R1751 VTAIL.n98 VTAIL.n97 1.16414
R1752 VTAIL.n89 VTAIL.n60 1.16414
R1753 VTAIL VTAIL.n199 0.591017
R1754 VTAIL.n189 VTAIL.n188 0.388379
R1755 VTAIL.n190 VTAIL.n154 0.388379
R1756 VTAIL.n39 VTAIL.n38 0.388379
R1757 VTAIL.n40 VTAIL.n4 0.388379
R1758 VTAIL.n144 VTAIL.n108 0.388379
R1759 VTAIL.n143 VTAIL.n142 0.388379
R1760 VTAIL.n94 VTAIL.n58 0.388379
R1761 VTAIL.n93 VTAIL.n92 0.388379
R1762 VTAIL.n170 VTAIL.n169 0.155672
R1763 VTAIL.n170 VTAIL.n161 0.155672
R1764 VTAIL.n177 VTAIL.n161 0.155672
R1765 VTAIL.n178 VTAIL.n177 0.155672
R1766 VTAIL.n178 VTAIL.n157 0.155672
R1767 VTAIL.n186 VTAIL.n157 0.155672
R1768 VTAIL.n187 VTAIL.n186 0.155672
R1769 VTAIL.n187 VTAIL.n153 0.155672
R1770 VTAIL.n195 VTAIL.n153 0.155672
R1771 VTAIL.n20 VTAIL.n19 0.155672
R1772 VTAIL.n20 VTAIL.n11 0.155672
R1773 VTAIL.n27 VTAIL.n11 0.155672
R1774 VTAIL.n28 VTAIL.n27 0.155672
R1775 VTAIL.n28 VTAIL.n7 0.155672
R1776 VTAIL.n36 VTAIL.n7 0.155672
R1777 VTAIL.n37 VTAIL.n36 0.155672
R1778 VTAIL.n37 VTAIL.n3 0.155672
R1779 VTAIL.n45 VTAIL.n3 0.155672
R1780 VTAIL.n149 VTAIL.n107 0.155672
R1781 VTAIL.n141 VTAIL.n107 0.155672
R1782 VTAIL.n141 VTAIL.n140 0.155672
R1783 VTAIL.n140 VTAIL.n111 0.155672
R1784 VTAIL.n133 VTAIL.n111 0.155672
R1785 VTAIL.n133 VTAIL.n132 0.155672
R1786 VTAIL.n132 VTAIL.n116 0.155672
R1787 VTAIL.n125 VTAIL.n116 0.155672
R1788 VTAIL.n125 VTAIL.n124 0.155672
R1789 VTAIL.n99 VTAIL.n57 0.155672
R1790 VTAIL.n91 VTAIL.n57 0.155672
R1791 VTAIL.n91 VTAIL.n90 0.155672
R1792 VTAIL.n90 VTAIL.n61 0.155672
R1793 VTAIL.n83 VTAIL.n61 0.155672
R1794 VTAIL.n83 VTAIL.n82 0.155672
R1795 VTAIL.n82 VTAIL.n66 0.155672
R1796 VTAIL.n75 VTAIL.n66 0.155672
R1797 VTAIL.n75 VTAIL.n74 0.155672
R1798 VP.n27 VP.n26 161.3
R1799 VP.n28 VP.n23 161.3
R1800 VP.n30 VP.n29 161.3
R1801 VP.n31 VP.n22 161.3
R1802 VP.n33 VP.n32 161.3
R1803 VP.n34 VP.n21 161.3
R1804 VP.n36 VP.n35 161.3
R1805 VP.n37 VP.n20 161.3
R1806 VP.n39 VP.n38 161.3
R1807 VP.n40 VP.n19 161.3
R1808 VP.n42 VP.n41 161.3
R1809 VP.n43 VP.n18 161.3
R1810 VP.n45 VP.n44 161.3
R1811 VP.n47 VP.n46 161.3
R1812 VP.n48 VP.n16 161.3
R1813 VP.n50 VP.n49 161.3
R1814 VP.n51 VP.n15 161.3
R1815 VP.n53 VP.n52 161.3
R1816 VP.n54 VP.n14 161.3
R1817 VP.n96 VP.n0 161.3
R1818 VP.n95 VP.n94 161.3
R1819 VP.n93 VP.n1 161.3
R1820 VP.n92 VP.n91 161.3
R1821 VP.n90 VP.n2 161.3
R1822 VP.n89 VP.n88 161.3
R1823 VP.n87 VP.n86 161.3
R1824 VP.n85 VP.n4 161.3
R1825 VP.n84 VP.n83 161.3
R1826 VP.n82 VP.n5 161.3
R1827 VP.n81 VP.n80 161.3
R1828 VP.n79 VP.n6 161.3
R1829 VP.n78 VP.n77 161.3
R1830 VP.n76 VP.n7 161.3
R1831 VP.n75 VP.n74 161.3
R1832 VP.n73 VP.n8 161.3
R1833 VP.n72 VP.n71 161.3
R1834 VP.n70 VP.n9 161.3
R1835 VP.n69 VP.n68 161.3
R1836 VP.n66 VP.n10 161.3
R1837 VP.n65 VP.n64 161.3
R1838 VP.n63 VP.n11 161.3
R1839 VP.n62 VP.n61 161.3
R1840 VP.n60 VP.n12 161.3
R1841 VP.n59 VP.n58 161.3
R1842 VP.n57 VP.n13 109.924
R1843 VP.n98 VP.n97 109.924
R1844 VP.n56 VP.n55 109.924
R1845 VP.n24 VP.t1 107.171
R1846 VP.n78 VP.t2 76.7968
R1847 VP.n13 VP.t5 76.7968
R1848 VP.n67 VP.t9 76.7968
R1849 VP.n3 VP.t4 76.7968
R1850 VP.n97 VP.t7 76.7968
R1851 VP.n36 VP.t0 76.7968
R1852 VP.n55 VP.t8 76.7968
R1853 VP.n17 VP.t3 76.7968
R1854 VP.n25 VP.t6 76.7968
R1855 VP.n25 VP.n24 73.1566
R1856 VP.n57 VP.n56 50.8292
R1857 VP.n61 VP.n11 42.0302
R1858 VP.n91 VP.n1 42.0302
R1859 VP.n49 VP.n15 42.0302
R1860 VP.n73 VP.n72 41.0614
R1861 VP.n84 VP.n5 41.0614
R1862 VP.n42 VP.n19 41.0614
R1863 VP.n31 VP.n30 41.0614
R1864 VP.n74 VP.n73 40.0926
R1865 VP.n80 VP.n5 40.0926
R1866 VP.n38 VP.n19 40.0926
R1867 VP.n32 VP.n31 40.0926
R1868 VP.n65 VP.n11 39.1239
R1869 VP.n91 VP.n90 39.1239
R1870 VP.n49 VP.n48 39.1239
R1871 VP.n60 VP.n59 24.5923
R1872 VP.n61 VP.n60 24.5923
R1873 VP.n66 VP.n65 24.5923
R1874 VP.n68 VP.n9 24.5923
R1875 VP.n72 VP.n9 24.5923
R1876 VP.n74 VP.n7 24.5923
R1877 VP.n78 VP.n7 24.5923
R1878 VP.n79 VP.n78 24.5923
R1879 VP.n80 VP.n79 24.5923
R1880 VP.n85 VP.n84 24.5923
R1881 VP.n86 VP.n85 24.5923
R1882 VP.n90 VP.n89 24.5923
R1883 VP.n95 VP.n1 24.5923
R1884 VP.n96 VP.n95 24.5923
R1885 VP.n53 VP.n15 24.5923
R1886 VP.n54 VP.n53 24.5923
R1887 VP.n43 VP.n42 24.5923
R1888 VP.n44 VP.n43 24.5923
R1889 VP.n48 VP.n47 24.5923
R1890 VP.n32 VP.n21 24.5923
R1891 VP.n36 VP.n21 24.5923
R1892 VP.n37 VP.n36 24.5923
R1893 VP.n38 VP.n37 24.5923
R1894 VP.n26 VP.n23 24.5923
R1895 VP.n30 VP.n23 24.5923
R1896 VP.n67 VP.n66 24.1005
R1897 VP.n89 VP.n3 24.1005
R1898 VP.n47 VP.n17 24.1005
R1899 VP.n27 VP.n24 7.42269
R1900 VP.n59 VP.n13 0.984173
R1901 VP.n97 VP.n96 0.984173
R1902 VP.n55 VP.n54 0.984173
R1903 VP.n68 VP.n67 0.492337
R1904 VP.n86 VP.n3 0.492337
R1905 VP.n44 VP.n17 0.492337
R1906 VP.n26 VP.n25 0.492337
R1907 VP.n56 VP.n14 0.278335
R1908 VP.n58 VP.n57 0.278335
R1909 VP.n98 VP.n0 0.278335
R1910 VP.n28 VP.n27 0.189894
R1911 VP.n29 VP.n28 0.189894
R1912 VP.n29 VP.n22 0.189894
R1913 VP.n33 VP.n22 0.189894
R1914 VP.n34 VP.n33 0.189894
R1915 VP.n35 VP.n34 0.189894
R1916 VP.n35 VP.n20 0.189894
R1917 VP.n39 VP.n20 0.189894
R1918 VP.n40 VP.n39 0.189894
R1919 VP.n41 VP.n40 0.189894
R1920 VP.n41 VP.n18 0.189894
R1921 VP.n45 VP.n18 0.189894
R1922 VP.n46 VP.n45 0.189894
R1923 VP.n46 VP.n16 0.189894
R1924 VP.n50 VP.n16 0.189894
R1925 VP.n51 VP.n50 0.189894
R1926 VP.n52 VP.n51 0.189894
R1927 VP.n52 VP.n14 0.189894
R1928 VP.n58 VP.n12 0.189894
R1929 VP.n62 VP.n12 0.189894
R1930 VP.n63 VP.n62 0.189894
R1931 VP.n64 VP.n63 0.189894
R1932 VP.n64 VP.n10 0.189894
R1933 VP.n69 VP.n10 0.189894
R1934 VP.n70 VP.n69 0.189894
R1935 VP.n71 VP.n70 0.189894
R1936 VP.n71 VP.n8 0.189894
R1937 VP.n75 VP.n8 0.189894
R1938 VP.n76 VP.n75 0.189894
R1939 VP.n77 VP.n76 0.189894
R1940 VP.n77 VP.n6 0.189894
R1941 VP.n81 VP.n6 0.189894
R1942 VP.n82 VP.n81 0.189894
R1943 VP.n83 VP.n82 0.189894
R1944 VP.n83 VP.n4 0.189894
R1945 VP.n87 VP.n4 0.189894
R1946 VP.n88 VP.n87 0.189894
R1947 VP.n88 VP.n2 0.189894
R1948 VP.n92 VP.n2 0.189894
R1949 VP.n93 VP.n92 0.189894
R1950 VP.n94 VP.n93 0.189894
R1951 VP.n94 VP.n0 0.189894
R1952 VP VP.n98 0.153485
R1953 VDD1.n40 VDD1.n0 756.745
R1954 VDD1.n87 VDD1.n47 756.745
R1955 VDD1.n41 VDD1.n40 585
R1956 VDD1.n39 VDD1.n38 585
R1957 VDD1.n37 VDD1.n3 585
R1958 VDD1.n7 VDD1.n4 585
R1959 VDD1.n32 VDD1.n31 585
R1960 VDD1.n30 VDD1.n29 585
R1961 VDD1.n9 VDD1.n8 585
R1962 VDD1.n24 VDD1.n23 585
R1963 VDD1.n22 VDD1.n21 585
R1964 VDD1.n13 VDD1.n12 585
R1965 VDD1.n16 VDD1.n15 585
R1966 VDD1.n62 VDD1.n61 585
R1967 VDD1.n59 VDD1.n58 585
R1968 VDD1.n68 VDD1.n67 585
R1969 VDD1.n70 VDD1.n69 585
R1970 VDD1.n55 VDD1.n54 585
R1971 VDD1.n76 VDD1.n75 585
R1972 VDD1.n79 VDD1.n78 585
R1973 VDD1.n77 VDD1.n51 585
R1974 VDD1.n84 VDD1.n50 585
R1975 VDD1.n86 VDD1.n85 585
R1976 VDD1.n88 VDD1.n87 585
R1977 VDD1.t8 VDD1.n14 329.039
R1978 VDD1.t4 VDD1.n60 329.038
R1979 VDD1.n40 VDD1.n39 171.744
R1980 VDD1.n39 VDD1.n3 171.744
R1981 VDD1.n7 VDD1.n3 171.744
R1982 VDD1.n31 VDD1.n7 171.744
R1983 VDD1.n31 VDD1.n30 171.744
R1984 VDD1.n30 VDD1.n8 171.744
R1985 VDD1.n23 VDD1.n8 171.744
R1986 VDD1.n23 VDD1.n22 171.744
R1987 VDD1.n22 VDD1.n12 171.744
R1988 VDD1.n15 VDD1.n12 171.744
R1989 VDD1.n61 VDD1.n58 171.744
R1990 VDD1.n68 VDD1.n58 171.744
R1991 VDD1.n69 VDD1.n68 171.744
R1992 VDD1.n69 VDD1.n54 171.744
R1993 VDD1.n76 VDD1.n54 171.744
R1994 VDD1.n78 VDD1.n76 171.744
R1995 VDD1.n78 VDD1.n77 171.744
R1996 VDD1.n77 VDD1.n50 171.744
R1997 VDD1.n86 VDD1.n50 171.744
R1998 VDD1.n87 VDD1.n86 171.744
R1999 VDD1.n15 VDD1.t8 85.8723
R2000 VDD1.n61 VDD1.t4 85.8723
R2001 VDD1.n95 VDD1.n94 82.5828
R2002 VDD1.n46 VDD1.n45 80.6922
R2003 VDD1.n97 VDD1.n96 80.692
R2004 VDD1.n93 VDD1.n92 80.692
R2005 VDD1.n46 VDD1.n44 51.8468
R2006 VDD1.n93 VDD1.n91 51.8468
R2007 VDD1.n97 VDD1.n95 45.2832
R2008 VDD1.n38 VDD1.n37 13.1884
R2009 VDD1.n85 VDD1.n84 13.1884
R2010 VDD1.n41 VDD1.n2 12.8005
R2011 VDD1.n36 VDD1.n4 12.8005
R2012 VDD1.n83 VDD1.n51 12.8005
R2013 VDD1.n88 VDD1.n49 12.8005
R2014 VDD1.n42 VDD1.n0 12.0247
R2015 VDD1.n33 VDD1.n32 12.0247
R2016 VDD1.n80 VDD1.n79 12.0247
R2017 VDD1.n89 VDD1.n47 12.0247
R2018 VDD1.n29 VDD1.n6 11.249
R2019 VDD1.n75 VDD1.n53 11.249
R2020 VDD1.n16 VDD1.n14 10.7239
R2021 VDD1.n62 VDD1.n60 10.7239
R2022 VDD1.n28 VDD1.n9 10.4732
R2023 VDD1.n74 VDD1.n55 10.4732
R2024 VDD1.n25 VDD1.n24 9.69747
R2025 VDD1.n71 VDD1.n70 9.69747
R2026 VDD1.n44 VDD1.n43 9.45567
R2027 VDD1.n91 VDD1.n90 9.45567
R2028 VDD1.n18 VDD1.n17 9.3005
R2029 VDD1.n20 VDD1.n19 9.3005
R2030 VDD1.n11 VDD1.n10 9.3005
R2031 VDD1.n26 VDD1.n25 9.3005
R2032 VDD1.n28 VDD1.n27 9.3005
R2033 VDD1.n6 VDD1.n5 9.3005
R2034 VDD1.n34 VDD1.n33 9.3005
R2035 VDD1.n36 VDD1.n35 9.3005
R2036 VDD1.n43 VDD1.n42 9.3005
R2037 VDD1.n2 VDD1.n1 9.3005
R2038 VDD1.n90 VDD1.n89 9.3005
R2039 VDD1.n49 VDD1.n48 9.3005
R2040 VDD1.n64 VDD1.n63 9.3005
R2041 VDD1.n66 VDD1.n65 9.3005
R2042 VDD1.n57 VDD1.n56 9.3005
R2043 VDD1.n72 VDD1.n71 9.3005
R2044 VDD1.n74 VDD1.n73 9.3005
R2045 VDD1.n53 VDD1.n52 9.3005
R2046 VDD1.n81 VDD1.n80 9.3005
R2047 VDD1.n83 VDD1.n82 9.3005
R2048 VDD1.n21 VDD1.n11 8.92171
R2049 VDD1.n67 VDD1.n57 8.92171
R2050 VDD1.n20 VDD1.n13 8.14595
R2051 VDD1.n66 VDD1.n59 8.14595
R2052 VDD1.n17 VDD1.n16 7.3702
R2053 VDD1.n63 VDD1.n62 7.3702
R2054 VDD1.n17 VDD1.n13 5.81868
R2055 VDD1.n63 VDD1.n59 5.81868
R2056 VDD1.n21 VDD1.n20 5.04292
R2057 VDD1.n67 VDD1.n66 5.04292
R2058 VDD1.n24 VDD1.n11 4.26717
R2059 VDD1.n70 VDD1.n57 4.26717
R2060 VDD1.n96 VDD1.t6 3.80671
R2061 VDD1.n96 VDD1.t1 3.80671
R2062 VDD1.n45 VDD1.t3 3.80671
R2063 VDD1.n45 VDD1.t9 3.80671
R2064 VDD1.n94 VDD1.t5 3.80671
R2065 VDD1.n94 VDD1.t2 3.80671
R2066 VDD1.n92 VDD1.t0 3.80671
R2067 VDD1.n92 VDD1.t7 3.80671
R2068 VDD1.n25 VDD1.n9 3.49141
R2069 VDD1.n71 VDD1.n55 3.49141
R2070 VDD1.n29 VDD1.n28 2.71565
R2071 VDD1.n75 VDD1.n74 2.71565
R2072 VDD1.n18 VDD1.n14 2.41285
R2073 VDD1.n64 VDD1.n60 2.41285
R2074 VDD1.n44 VDD1.n0 1.93989
R2075 VDD1.n32 VDD1.n6 1.93989
R2076 VDD1.n79 VDD1.n53 1.93989
R2077 VDD1.n91 VDD1.n47 1.93989
R2078 VDD1 VDD1.n97 1.88843
R2079 VDD1.n42 VDD1.n41 1.16414
R2080 VDD1.n33 VDD1.n4 1.16414
R2081 VDD1.n80 VDD1.n51 1.16414
R2082 VDD1.n89 VDD1.n88 1.16414
R2083 VDD1 VDD1.n46 0.707397
R2084 VDD1.n95 VDD1.n93 0.593861
R2085 VDD1.n38 VDD1.n2 0.388379
R2086 VDD1.n37 VDD1.n36 0.388379
R2087 VDD1.n84 VDD1.n83 0.388379
R2088 VDD1.n85 VDD1.n49 0.388379
R2089 VDD1.n43 VDD1.n1 0.155672
R2090 VDD1.n35 VDD1.n1 0.155672
R2091 VDD1.n35 VDD1.n34 0.155672
R2092 VDD1.n34 VDD1.n5 0.155672
R2093 VDD1.n27 VDD1.n5 0.155672
R2094 VDD1.n27 VDD1.n26 0.155672
R2095 VDD1.n26 VDD1.n10 0.155672
R2096 VDD1.n19 VDD1.n10 0.155672
R2097 VDD1.n19 VDD1.n18 0.155672
R2098 VDD1.n65 VDD1.n64 0.155672
R2099 VDD1.n65 VDD1.n56 0.155672
R2100 VDD1.n72 VDD1.n56 0.155672
R2101 VDD1.n73 VDD1.n72 0.155672
R2102 VDD1.n73 VDD1.n52 0.155672
R2103 VDD1.n81 VDD1.n52 0.155672
R2104 VDD1.n82 VDD1.n81 0.155672
R2105 VDD1.n82 VDD1.n48 0.155672
R2106 VDD1.n90 VDD1.n48 0.155672
C0 w_n4582_n2676# VDD1 2.57272f
C1 VTAIL VDD1 8.83939f
C2 B VDD1 2.23774f
C3 VP VDD1 8.232361f
C4 VDD2 VDD1 2.22325f
C5 VN VDD1 0.153471f
C6 w_n4582_n2676# VTAIL 2.72758f
C7 w_n4582_n2676# B 9.71158f
C8 VTAIL B 2.98465f
C9 VP w_n4582_n2676# 10.3625f
C10 VP VTAIL 8.63958f
C11 w_n4582_n2676# VDD2 2.72043f
C12 VTAIL VDD2 8.89173f
C13 VP B 2.27089f
C14 w_n4582_n2676# VN 9.76566f
C15 VDD2 B 2.35877f
C16 VTAIL VN 8.625349f
C17 VN B 1.2669f
C18 VP VDD2 0.593442f
C19 VP VN 7.87227f
C20 VDD2 VN 7.79565f
C21 VDD2 VSUBS 2.141299f
C22 VDD1 VSUBS 1.906363f
C23 VTAIL VSUBS 1.204452f
C24 VN VSUBS 7.726281f
C25 VP VSUBS 4.202421f
C26 B VSUBS 5.176231f
C27 w_n4582_n2676# VSUBS 0.151921p
C28 VDD1.n0 VSUBS 0.032395f
C29 VDD1.n1 VSUBS 0.031813f
C30 VDD1.n2 VSUBS 0.017095f
C31 VDD1.n3 VSUBS 0.040406f
C32 VDD1.n4 VSUBS 0.018101f
C33 VDD1.n5 VSUBS 0.031813f
C34 VDD1.n6 VSUBS 0.017095f
C35 VDD1.n7 VSUBS 0.040406f
C36 VDD1.n8 VSUBS 0.040406f
C37 VDD1.n9 VSUBS 0.018101f
C38 VDD1.n10 VSUBS 0.031813f
C39 VDD1.n11 VSUBS 0.017095f
C40 VDD1.n12 VSUBS 0.040406f
C41 VDD1.n13 VSUBS 0.018101f
C42 VDD1.n14 VSUBS 0.200831f
C43 VDD1.t8 VSUBS 0.086765f
C44 VDD1.n15 VSUBS 0.030305f
C45 VDD1.n16 VSUBS 0.030396f
C46 VDD1.n17 VSUBS 0.017095f
C47 VDD1.n18 VSUBS 1.08066f
C48 VDD1.n19 VSUBS 0.031813f
C49 VDD1.n20 VSUBS 0.017095f
C50 VDD1.n21 VSUBS 0.018101f
C51 VDD1.n22 VSUBS 0.040406f
C52 VDD1.n23 VSUBS 0.040406f
C53 VDD1.n24 VSUBS 0.018101f
C54 VDD1.n25 VSUBS 0.017095f
C55 VDD1.n26 VSUBS 0.031813f
C56 VDD1.n27 VSUBS 0.031813f
C57 VDD1.n28 VSUBS 0.017095f
C58 VDD1.n29 VSUBS 0.018101f
C59 VDD1.n30 VSUBS 0.040406f
C60 VDD1.n31 VSUBS 0.040406f
C61 VDD1.n32 VSUBS 0.018101f
C62 VDD1.n33 VSUBS 0.017095f
C63 VDD1.n34 VSUBS 0.031813f
C64 VDD1.n35 VSUBS 0.031813f
C65 VDD1.n36 VSUBS 0.017095f
C66 VDD1.n37 VSUBS 0.017598f
C67 VDD1.n38 VSUBS 0.017598f
C68 VDD1.n39 VSUBS 0.040406f
C69 VDD1.n40 VSUBS 0.089098f
C70 VDD1.n41 VSUBS 0.018101f
C71 VDD1.n42 VSUBS 0.017095f
C72 VDD1.n43 VSUBS 0.074404f
C73 VDD1.n44 VSUBS 0.082809f
C74 VDD1.t3 VSUBS 0.214693f
C75 VDD1.t9 VSUBS 0.214693f
C76 VDD1.n45 VSUBS 1.57151f
C77 VDD1.n46 VSUBS 1.20207f
C78 VDD1.n47 VSUBS 0.032395f
C79 VDD1.n48 VSUBS 0.031813f
C80 VDD1.n49 VSUBS 0.017095f
C81 VDD1.n50 VSUBS 0.040406f
C82 VDD1.n51 VSUBS 0.018101f
C83 VDD1.n52 VSUBS 0.031813f
C84 VDD1.n53 VSUBS 0.017095f
C85 VDD1.n54 VSUBS 0.040406f
C86 VDD1.n55 VSUBS 0.018101f
C87 VDD1.n56 VSUBS 0.031813f
C88 VDD1.n57 VSUBS 0.017095f
C89 VDD1.n58 VSUBS 0.040406f
C90 VDD1.n59 VSUBS 0.018101f
C91 VDD1.n60 VSUBS 0.200831f
C92 VDD1.t4 VSUBS 0.086765f
C93 VDD1.n61 VSUBS 0.030305f
C94 VDD1.n62 VSUBS 0.030396f
C95 VDD1.n63 VSUBS 0.017095f
C96 VDD1.n64 VSUBS 1.08066f
C97 VDD1.n65 VSUBS 0.031813f
C98 VDD1.n66 VSUBS 0.017095f
C99 VDD1.n67 VSUBS 0.018101f
C100 VDD1.n68 VSUBS 0.040406f
C101 VDD1.n69 VSUBS 0.040406f
C102 VDD1.n70 VSUBS 0.018101f
C103 VDD1.n71 VSUBS 0.017095f
C104 VDD1.n72 VSUBS 0.031813f
C105 VDD1.n73 VSUBS 0.031813f
C106 VDD1.n74 VSUBS 0.017095f
C107 VDD1.n75 VSUBS 0.018101f
C108 VDD1.n76 VSUBS 0.040406f
C109 VDD1.n77 VSUBS 0.040406f
C110 VDD1.n78 VSUBS 0.040406f
C111 VDD1.n79 VSUBS 0.018101f
C112 VDD1.n80 VSUBS 0.017095f
C113 VDD1.n81 VSUBS 0.031813f
C114 VDD1.n82 VSUBS 0.031813f
C115 VDD1.n83 VSUBS 0.017095f
C116 VDD1.n84 VSUBS 0.017598f
C117 VDD1.n85 VSUBS 0.017598f
C118 VDD1.n86 VSUBS 0.040406f
C119 VDD1.n87 VSUBS 0.089098f
C120 VDD1.n88 VSUBS 0.018101f
C121 VDD1.n89 VSUBS 0.017095f
C122 VDD1.n90 VSUBS 0.074404f
C123 VDD1.n91 VSUBS 0.082809f
C124 VDD1.t0 VSUBS 0.214693f
C125 VDD1.t7 VSUBS 0.214693f
C126 VDD1.n92 VSUBS 1.57151f
C127 VDD1.n93 VSUBS 1.19168f
C128 VDD1.t5 VSUBS 0.214693f
C129 VDD1.t2 VSUBS 0.214693f
C130 VDD1.n94 VSUBS 1.59498f
C131 VDD1.n95 VSUBS 3.92706f
C132 VDD1.t6 VSUBS 0.214693f
C133 VDD1.t1 VSUBS 0.214693f
C134 VDD1.n96 VSUBS 1.57151f
C135 VDD1.n97 VSUBS 4.03261f
C136 VP.n0 VSUBS 0.044795f
C137 VP.t7 VSUBS 2.09435f
C138 VP.n1 VSUBS 0.066624f
C139 VP.n2 VSUBS 0.033979f
C140 VP.t4 VSUBS 2.09435f
C141 VP.n3 VSUBS 0.757579f
C142 VP.n4 VSUBS 0.033979f
C143 VP.n5 VSUBS 0.027454f
C144 VP.n6 VSUBS 0.033979f
C145 VP.t2 VSUBS 2.09435f
C146 VP.n7 VSUBS 0.06301f
C147 VP.n8 VSUBS 0.033979f
C148 VP.n9 VSUBS 0.06301f
C149 VP.n10 VSUBS 0.033979f
C150 VP.t9 VSUBS 2.09435f
C151 VP.n11 VSUBS 0.027541f
C152 VP.n12 VSUBS 0.033979f
C153 VP.t5 VSUBS 2.09435f
C154 VP.n13 VSUBS 0.858338f
C155 VP.n14 VSUBS 0.044795f
C156 VP.t8 VSUBS 2.09435f
C157 VP.n15 VSUBS 0.066624f
C158 VP.n16 VSUBS 0.033979f
C159 VP.t3 VSUBS 2.09435f
C160 VP.n17 VSUBS 0.757579f
C161 VP.n18 VSUBS 0.033979f
C162 VP.n19 VSUBS 0.027454f
C163 VP.n20 VSUBS 0.033979f
C164 VP.t0 VSUBS 2.09435f
C165 VP.n21 VSUBS 0.06301f
C166 VP.n22 VSUBS 0.033979f
C167 VP.n23 VSUBS 0.06301f
C168 VP.t1 VSUBS 2.36819f
C169 VP.n24 VSUBS 0.835393f
C170 VP.t6 VSUBS 2.09435f
C171 VP.n25 VSUBS 0.84497f
C172 VP.n26 VSUBS 0.032526f
C173 VP.n27 VSUBS 0.330185f
C174 VP.n28 VSUBS 0.033979f
C175 VP.n29 VSUBS 0.033979f
C176 VP.n30 VSUBS 0.067003f
C177 VP.n31 VSUBS 0.027454f
C178 VP.n32 VSUBS 0.06734f
C179 VP.n33 VSUBS 0.033979f
C180 VP.n34 VSUBS 0.033979f
C181 VP.n35 VSUBS 0.033979f
C182 VP.n36 VSUBS 0.789483f
C183 VP.n37 VSUBS 0.06301f
C184 VP.n38 VSUBS 0.06734f
C185 VP.n39 VSUBS 0.033979f
C186 VP.n40 VSUBS 0.033979f
C187 VP.n41 VSUBS 0.033979f
C188 VP.n42 VSUBS 0.067003f
C189 VP.n43 VSUBS 0.06301f
C190 VP.n44 VSUBS 0.032526f
C191 VP.n45 VSUBS 0.033979f
C192 VP.n46 VSUBS 0.033979f
C193 VP.n47 VSUBS 0.062388f
C194 VP.n48 VSUBS 0.067632f
C195 VP.n49 VSUBS 0.027541f
C196 VP.n50 VSUBS 0.033979f
C197 VP.n51 VSUBS 0.033979f
C198 VP.n52 VSUBS 0.033979f
C199 VP.n53 VSUBS 0.06301f
C200 VP.n54 VSUBS 0.033148f
C201 VP.n55 VSUBS 0.858338f
C202 VP.n56 VSUBS 1.94294f
C203 VP.n57 VSUBS 1.96704f
C204 VP.n58 VSUBS 0.044795f
C205 VP.n59 VSUBS 0.033148f
C206 VP.n60 VSUBS 0.06301f
C207 VP.n61 VSUBS 0.066624f
C208 VP.n62 VSUBS 0.033979f
C209 VP.n63 VSUBS 0.033979f
C210 VP.n64 VSUBS 0.033979f
C211 VP.n65 VSUBS 0.067632f
C212 VP.n66 VSUBS 0.062388f
C213 VP.n67 VSUBS 0.757579f
C214 VP.n68 VSUBS 0.032526f
C215 VP.n69 VSUBS 0.033979f
C216 VP.n70 VSUBS 0.033979f
C217 VP.n71 VSUBS 0.033979f
C218 VP.n72 VSUBS 0.067003f
C219 VP.n73 VSUBS 0.027454f
C220 VP.n74 VSUBS 0.06734f
C221 VP.n75 VSUBS 0.033979f
C222 VP.n76 VSUBS 0.033979f
C223 VP.n77 VSUBS 0.033979f
C224 VP.n78 VSUBS 0.789483f
C225 VP.n79 VSUBS 0.06301f
C226 VP.n80 VSUBS 0.06734f
C227 VP.n81 VSUBS 0.033979f
C228 VP.n82 VSUBS 0.033979f
C229 VP.n83 VSUBS 0.033979f
C230 VP.n84 VSUBS 0.067003f
C231 VP.n85 VSUBS 0.06301f
C232 VP.n86 VSUBS 0.032526f
C233 VP.n87 VSUBS 0.033979f
C234 VP.n88 VSUBS 0.033979f
C235 VP.n89 VSUBS 0.062388f
C236 VP.n90 VSUBS 0.067632f
C237 VP.n91 VSUBS 0.027541f
C238 VP.n92 VSUBS 0.033979f
C239 VP.n93 VSUBS 0.033979f
C240 VP.n94 VSUBS 0.033979f
C241 VP.n95 VSUBS 0.06301f
C242 VP.n96 VSUBS 0.033148f
C243 VP.n97 VSUBS 0.858338f
C244 VP.n98 VSUBS 0.062914f
C245 VTAIL.t11 VSUBS 0.207204f
C246 VTAIL.t13 VSUBS 0.207204f
C247 VTAIL.n0 VSUBS 1.37933f
C248 VTAIL.n1 VSUBS 1.00176f
C249 VTAIL.n2 VSUBS 0.031265f
C250 VTAIL.n3 VSUBS 0.030703f
C251 VTAIL.n4 VSUBS 0.016499f
C252 VTAIL.n5 VSUBS 0.038997f
C253 VTAIL.n6 VSUBS 0.017469f
C254 VTAIL.n7 VSUBS 0.030703f
C255 VTAIL.n8 VSUBS 0.016499f
C256 VTAIL.n9 VSUBS 0.038997f
C257 VTAIL.n10 VSUBS 0.017469f
C258 VTAIL.n11 VSUBS 0.030703f
C259 VTAIL.n12 VSUBS 0.016499f
C260 VTAIL.n13 VSUBS 0.038997f
C261 VTAIL.n14 VSUBS 0.017469f
C262 VTAIL.n15 VSUBS 0.193826f
C263 VTAIL.t6 VSUBS 0.083738f
C264 VTAIL.n16 VSUBS 0.029248f
C265 VTAIL.n17 VSUBS 0.029335f
C266 VTAIL.n18 VSUBS 0.016499f
C267 VTAIL.n19 VSUBS 1.04296f
C268 VTAIL.n20 VSUBS 0.030703f
C269 VTAIL.n21 VSUBS 0.016499f
C270 VTAIL.n22 VSUBS 0.017469f
C271 VTAIL.n23 VSUBS 0.038997f
C272 VTAIL.n24 VSUBS 0.038997f
C273 VTAIL.n25 VSUBS 0.017469f
C274 VTAIL.n26 VSUBS 0.016499f
C275 VTAIL.n27 VSUBS 0.030703f
C276 VTAIL.n28 VSUBS 0.030703f
C277 VTAIL.n29 VSUBS 0.016499f
C278 VTAIL.n30 VSUBS 0.017469f
C279 VTAIL.n31 VSUBS 0.038997f
C280 VTAIL.n32 VSUBS 0.038997f
C281 VTAIL.n33 VSUBS 0.038997f
C282 VTAIL.n34 VSUBS 0.017469f
C283 VTAIL.n35 VSUBS 0.016499f
C284 VTAIL.n36 VSUBS 0.030703f
C285 VTAIL.n37 VSUBS 0.030703f
C286 VTAIL.n38 VSUBS 0.016499f
C287 VTAIL.n39 VSUBS 0.016984f
C288 VTAIL.n40 VSUBS 0.016984f
C289 VTAIL.n41 VSUBS 0.038997f
C290 VTAIL.n42 VSUBS 0.08599f
C291 VTAIL.n43 VSUBS 0.017469f
C292 VTAIL.n44 VSUBS 0.016499f
C293 VTAIL.n45 VSUBS 0.071808f
C294 VTAIL.n46 VSUBS 0.042895f
C295 VTAIL.n47 VSUBS 0.458249f
C296 VTAIL.t3 VSUBS 0.207204f
C297 VTAIL.t5 VSUBS 0.207204f
C298 VTAIL.n48 VSUBS 1.37933f
C299 VTAIL.n49 VSUBS 1.14206f
C300 VTAIL.t8 VSUBS 0.207204f
C301 VTAIL.t7 VSUBS 0.207204f
C302 VTAIL.n50 VSUBS 1.37933f
C303 VTAIL.n51 VSUBS 2.5442f
C304 VTAIL.t15 VSUBS 0.207204f
C305 VTAIL.t18 VSUBS 0.207204f
C306 VTAIL.n52 VSUBS 1.37934f
C307 VTAIL.n53 VSUBS 2.54419f
C308 VTAIL.t14 VSUBS 0.207204f
C309 VTAIL.t10 VSUBS 0.207204f
C310 VTAIL.n54 VSUBS 1.37934f
C311 VTAIL.n55 VSUBS 1.14205f
C312 VTAIL.n56 VSUBS 0.031265f
C313 VTAIL.n57 VSUBS 0.030703f
C314 VTAIL.n58 VSUBS 0.016499f
C315 VTAIL.n59 VSUBS 0.038997f
C316 VTAIL.n60 VSUBS 0.017469f
C317 VTAIL.n61 VSUBS 0.030703f
C318 VTAIL.n62 VSUBS 0.016499f
C319 VTAIL.n63 VSUBS 0.038997f
C320 VTAIL.n64 VSUBS 0.038997f
C321 VTAIL.n65 VSUBS 0.017469f
C322 VTAIL.n66 VSUBS 0.030703f
C323 VTAIL.n67 VSUBS 0.016499f
C324 VTAIL.n68 VSUBS 0.038997f
C325 VTAIL.n69 VSUBS 0.017469f
C326 VTAIL.n70 VSUBS 0.193826f
C327 VTAIL.t16 VSUBS 0.083738f
C328 VTAIL.n71 VSUBS 0.029248f
C329 VTAIL.n72 VSUBS 0.029335f
C330 VTAIL.n73 VSUBS 0.016499f
C331 VTAIL.n74 VSUBS 1.04296f
C332 VTAIL.n75 VSUBS 0.030703f
C333 VTAIL.n76 VSUBS 0.016499f
C334 VTAIL.n77 VSUBS 0.017469f
C335 VTAIL.n78 VSUBS 0.038997f
C336 VTAIL.n79 VSUBS 0.038997f
C337 VTAIL.n80 VSUBS 0.017469f
C338 VTAIL.n81 VSUBS 0.016499f
C339 VTAIL.n82 VSUBS 0.030703f
C340 VTAIL.n83 VSUBS 0.030703f
C341 VTAIL.n84 VSUBS 0.016499f
C342 VTAIL.n85 VSUBS 0.017469f
C343 VTAIL.n86 VSUBS 0.038997f
C344 VTAIL.n87 VSUBS 0.038997f
C345 VTAIL.n88 VSUBS 0.017469f
C346 VTAIL.n89 VSUBS 0.016499f
C347 VTAIL.n90 VSUBS 0.030703f
C348 VTAIL.n91 VSUBS 0.030703f
C349 VTAIL.n92 VSUBS 0.016499f
C350 VTAIL.n93 VSUBS 0.016984f
C351 VTAIL.n94 VSUBS 0.016984f
C352 VTAIL.n95 VSUBS 0.038997f
C353 VTAIL.n96 VSUBS 0.08599f
C354 VTAIL.n97 VSUBS 0.017469f
C355 VTAIL.n98 VSUBS 0.016499f
C356 VTAIL.n99 VSUBS 0.071808f
C357 VTAIL.n100 VSUBS 0.042895f
C358 VTAIL.n101 VSUBS 0.458249f
C359 VTAIL.t4 VSUBS 0.207204f
C360 VTAIL.t9 VSUBS 0.207204f
C361 VTAIL.n102 VSUBS 1.37934f
C362 VTAIL.n103 VSUBS 1.06018f
C363 VTAIL.t2 VSUBS 0.207204f
C364 VTAIL.t0 VSUBS 0.207204f
C365 VTAIL.n104 VSUBS 1.37934f
C366 VTAIL.n105 VSUBS 1.14205f
C367 VTAIL.n106 VSUBS 0.031265f
C368 VTAIL.n107 VSUBS 0.030703f
C369 VTAIL.n108 VSUBS 0.016499f
C370 VTAIL.n109 VSUBS 0.038997f
C371 VTAIL.n110 VSUBS 0.017469f
C372 VTAIL.n111 VSUBS 0.030703f
C373 VTAIL.n112 VSUBS 0.016499f
C374 VTAIL.n113 VSUBS 0.038997f
C375 VTAIL.n114 VSUBS 0.038997f
C376 VTAIL.n115 VSUBS 0.017469f
C377 VTAIL.n116 VSUBS 0.030703f
C378 VTAIL.n117 VSUBS 0.016499f
C379 VTAIL.n118 VSUBS 0.038997f
C380 VTAIL.n119 VSUBS 0.017469f
C381 VTAIL.n120 VSUBS 0.193826f
C382 VTAIL.t1 VSUBS 0.083738f
C383 VTAIL.n121 VSUBS 0.029248f
C384 VTAIL.n122 VSUBS 0.029335f
C385 VTAIL.n123 VSUBS 0.016499f
C386 VTAIL.n124 VSUBS 1.04296f
C387 VTAIL.n125 VSUBS 0.030703f
C388 VTAIL.n126 VSUBS 0.016499f
C389 VTAIL.n127 VSUBS 0.017469f
C390 VTAIL.n128 VSUBS 0.038997f
C391 VTAIL.n129 VSUBS 0.038997f
C392 VTAIL.n130 VSUBS 0.017469f
C393 VTAIL.n131 VSUBS 0.016499f
C394 VTAIL.n132 VSUBS 0.030703f
C395 VTAIL.n133 VSUBS 0.030703f
C396 VTAIL.n134 VSUBS 0.016499f
C397 VTAIL.n135 VSUBS 0.017469f
C398 VTAIL.n136 VSUBS 0.038997f
C399 VTAIL.n137 VSUBS 0.038997f
C400 VTAIL.n138 VSUBS 0.017469f
C401 VTAIL.n139 VSUBS 0.016499f
C402 VTAIL.n140 VSUBS 0.030703f
C403 VTAIL.n141 VSUBS 0.030703f
C404 VTAIL.n142 VSUBS 0.016499f
C405 VTAIL.n143 VSUBS 0.016984f
C406 VTAIL.n144 VSUBS 0.016984f
C407 VTAIL.n145 VSUBS 0.038997f
C408 VTAIL.n146 VSUBS 0.08599f
C409 VTAIL.n147 VSUBS 0.017469f
C410 VTAIL.n148 VSUBS 0.016499f
C411 VTAIL.n149 VSUBS 0.071808f
C412 VTAIL.n150 VSUBS 0.042895f
C413 VTAIL.n151 VSUBS 1.68555f
C414 VTAIL.n152 VSUBS 0.031265f
C415 VTAIL.n153 VSUBS 0.030703f
C416 VTAIL.n154 VSUBS 0.016499f
C417 VTAIL.n155 VSUBS 0.038997f
C418 VTAIL.n156 VSUBS 0.017469f
C419 VTAIL.n157 VSUBS 0.030703f
C420 VTAIL.n158 VSUBS 0.016499f
C421 VTAIL.n159 VSUBS 0.038997f
C422 VTAIL.n160 VSUBS 0.017469f
C423 VTAIL.n161 VSUBS 0.030703f
C424 VTAIL.n162 VSUBS 0.016499f
C425 VTAIL.n163 VSUBS 0.038997f
C426 VTAIL.n164 VSUBS 0.017469f
C427 VTAIL.n165 VSUBS 0.193826f
C428 VTAIL.t12 VSUBS 0.083738f
C429 VTAIL.n166 VSUBS 0.029248f
C430 VTAIL.n167 VSUBS 0.029335f
C431 VTAIL.n168 VSUBS 0.016499f
C432 VTAIL.n169 VSUBS 1.04296f
C433 VTAIL.n170 VSUBS 0.030703f
C434 VTAIL.n171 VSUBS 0.016499f
C435 VTAIL.n172 VSUBS 0.017469f
C436 VTAIL.n173 VSUBS 0.038997f
C437 VTAIL.n174 VSUBS 0.038997f
C438 VTAIL.n175 VSUBS 0.017469f
C439 VTAIL.n176 VSUBS 0.016499f
C440 VTAIL.n177 VSUBS 0.030703f
C441 VTAIL.n178 VSUBS 0.030703f
C442 VTAIL.n179 VSUBS 0.016499f
C443 VTAIL.n180 VSUBS 0.017469f
C444 VTAIL.n181 VSUBS 0.038997f
C445 VTAIL.n182 VSUBS 0.038997f
C446 VTAIL.n183 VSUBS 0.038997f
C447 VTAIL.n184 VSUBS 0.017469f
C448 VTAIL.n185 VSUBS 0.016499f
C449 VTAIL.n186 VSUBS 0.030703f
C450 VTAIL.n187 VSUBS 0.030703f
C451 VTAIL.n188 VSUBS 0.016499f
C452 VTAIL.n189 VSUBS 0.016984f
C453 VTAIL.n190 VSUBS 0.016984f
C454 VTAIL.n191 VSUBS 0.038997f
C455 VTAIL.n192 VSUBS 0.08599f
C456 VTAIL.n193 VSUBS 0.017469f
C457 VTAIL.n194 VSUBS 0.016499f
C458 VTAIL.n195 VSUBS 0.071808f
C459 VTAIL.n196 VSUBS 0.042895f
C460 VTAIL.n197 VSUBS 1.68554f
C461 VTAIL.t17 VSUBS 0.207204f
C462 VTAIL.t19 VSUBS 0.207204f
C463 VTAIL.n198 VSUBS 1.37933f
C464 VTAIL.n199 VSUBS 0.943769f
C465 VDD2.n0 VSUBS 0.032555f
C466 VDD2.n1 VSUBS 0.03197f
C467 VDD2.n2 VSUBS 0.017179f
C468 VDD2.n3 VSUBS 0.040605f
C469 VDD2.n4 VSUBS 0.01819f
C470 VDD2.n5 VSUBS 0.03197f
C471 VDD2.n6 VSUBS 0.017179f
C472 VDD2.n7 VSUBS 0.040605f
C473 VDD2.n8 VSUBS 0.01819f
C474 VDD2.n9 VSUBS 0.03197f
C475 VDD2.n10 VSUBS 0.017179f
C476 VDD2.n11 VSUBS 0.040605f
C477 VDD2.n12 VSUBS 0.01819f
C478 VDD2.n13 VSUBS 0.201819f
C479 VDD2.t4 VSUBS 0.087191f
C480 VDD2.n14 VSUBS 0.030454f
C481 VDD2.n15 VSUBS 0.030545f
C482 VDD2.n16 VSUBS 0.017179f
C483 VDD2.n17 VSUBS 1.08597f
C484 VDD2.n18 VSUBS 0.03197f
C485 VDD2.n19 VSUBS 0.017179f
C486 VDD2.n20 VSUBS 0.01819f
C487 VDD2.n21 VSUBS 0.040605f
C488 VDD2.n22 VSUBS 0.040605f
C489 VDD2.n23 VSUBS 0.01819f
C490 VDD2.n24 VSUBS 0.017179f
C491 VDD2.n25 VSUBS 0.03197f
C492 VDD2.n26 VSUBS 0.03197f
C493 VDD2.n27 VSUBS 0.017179f
C494 VDD2.n28 VSUBS 0.01819f
C495 VDD2.n29 VSUBS 0.040605f
C496 VDD2.n30 VSUBS 0.040605f
C497 VDD2.n31 VSUBS 0.040605f
C498 VDD2.n32 VSUBS 0.01819f
C499 VDD2.n33 VSUBS 0.017179f
C500 VDD2.n34 VSUBS 0.03197f
C501 VDD2.n35 VSUBS 0.03197f
C502 VDD2.n36 VSUBS 0.017179f
C503 VDD2.n37 VSUBS 0.017684f
C504 VDD2.n38 VSUBS 0.017684f
C505 VDD2.n39 VSUBS 0.040605f
C506 VDD2.n40 VSUBS 0.089536f
C507 VDD2.n41 VSUBS 0.01819f
C508 VDD2.n42 VSUBS 0.017179f
C509 VDD2.n43 VSUBS 0.07477f
C510 VDD2.n44 VSUBS 0.083216f
C511 VDD2.t0 VSUBS 0.215749f
C512 VDD2.t7 VSUBS 0.215749f
C513 VDD2.n45 VSUBS 1.57924f
C514 VDD2.n46 VSUBS 1.19754f
C515 VDD2.t5 VSUBS 0.215749f
C516 VDD2.t8 VSUBS 0.215749f
C517 VDD2.n47 VSUBS 1.60283f
C518 VDD2.n48 VSUBS 3.78708f
C519 VDD2.n49 VSUBS 0.032555f
C520 VDD2.n50 VSUBS 0.03197f
C521 VDD2.n51 VSUBS 0.017179f
C522 VDD2.n52 VSUBS 0.040605f
C523 VDD2.n53 VSUBS 0.01819f
C524 VDD2.n54 VSUBS 0.03197f
C525 VDD2.n55 VSUBS 0.017179f
C526 VDD2.n56 VSUBS 0.040605f
C527 VDD2.n57 VSUBS 0.040605f
C528 VDD2.n58 VSUBS 0.01819f
C529 VDD2.n59 VSUBS 0.03197f
C530 VDD2.n60 VSUBS 0.017179f
C531 VDD2.n61 VSUBS 0.040605f
C532 VDD2.n62 VSUBS 0.01819f
C533 VDD2.n63 VSUBS 0.201819f
C534 VDD2.t6 VSUBS 0.087191f
C535 VDD2.n64 VSUBS 0.030454f
C536 VDD2.n65 VSUBS 0.030545f
C537 VDD2.n66 VSUBS 0.017179f
C538 VDD2.n67 VSUBS 1.08597f
C539 VDD2.n68 VSUBS 0.03197f
C540 VDD2.n69 VSUBS 0.017179f
C541 VDD2.n70 VSUBS 0.01819f
C542 VDD2.n71 VSUBS 0.040605f
C543 VDD2.n72 VSUBS 0.040605f
C544 VDD2.n73 VSUBS 0.01819f
C545 VDD2.n74 VSUBS 0.017179f
C546 VDD2.n75 VSUBS 0.03197f
C547 VDD2.n76 VSUBS 0.03197f
C548 VDD2.n77 VSUBS 0.017179f
C549 VDD2.n78 VSUBS 0.01819f
C550 VDD2.n79 VSUBS 0.040605f
C551 VDD2.n80 VSUBS 0.040605f
C552 VDD2.n81 VSUBS 0.01819f
C553 VDD2.n82 VSUBS 0.017179f
C554 VDD2.n83 VSUBS 0.03197f
C555 VDD2.n84 VSUBS 0.03197f
C556 VDD2.n85 VSUBS 0.017179f
C557 VDD2.n86 VSUBS 0.017684f
C558 VDD2.n87 VSUBS 0.017684f
C559 VDD2.n88 VSUBS 0.040605f
C560 VDD2.n89 VSUBS 0.089536f
C561 VDD2.n90 VSUBS 0.01819f
C562 VDD2.n91 VSUBS 0.017179f
C563 VDD2.n92 VSUBS 0.07477f
C564 VDD2.n93 VSUBS 0.066732f
C565 VDD2.n94 VSUBS 3.39338f
C566 VDD2.t9 VSUBS 0.215749f
C567 VDD2.t3 VSUBS 0.215749f
C568 VDD2.n95 VSUBS 1.57925f
C569 VDD2.n96 VSUBS 0.895106f
C570 VDD2.t2 VSUBS 0.215749f
C571 VDD2.t1 VSUBS 0.215749f
C572 VDD2.n97 VSUBS 1.60278f
C573 VN.n0 VSUBS 0.04079f
C574 VN.t7 VSUBS 1.90712f
C575 VN.n1 VSUBS 0.060668f
C576 VN.n2 VSUBS 0.030941f
C577 VN.t0 VSUBS 1.90712f
C578 VN.n3 VSUBS 0.689853f
C579 VN.n4 VSUBS 0.030941f
C580 VN.n5 VSUBS 0.025f
C581 VN.n6 VSUBS 0.030941f
C582 VN.t2 VSUBS 1.90712f
C583 VN.n7 VSUBS 0.057377f
C584 VN.n8 VSUBS 0.030941f
C585 VN.n9 VSUBS 0.057377f
C586 VN.t8 VSUBS 2.15648f
C587 VN.n10 VSUBS 0.760711f
C588 VN.t6 VSUBS 1.90712f
C589 VN.n11 VSUBS 0.769432f
C590 VN.n12 VSUBS 0.029618f
C591 VN.n13 VSUBS 0.300667f
C592 VN.n14 VSUBS 0.030941f
C593 VN.n15 VSUBS 0.030941f
C594 VN.n16 VSUBS 0.061013f
C595 VN.n17 VSUBS 0.025f
C596 VN.n18 VSUBS 0.06132f
C597 VN.n19 VSUBS 0.030941f
C598 VN.n20 VSUBS 0.030941f
C599 VN.n21 VSUBS 0.030941f
C600 VN.n22 VSUBS 0.718905f
C601 VN.n23 VSUBS 0.057377f
C602 VN.n24 VSUBS 0.06132f
C603 VN.n25 VSUBS 0.030941f
C604 VN.n26 VSUBS 0.030941f
C605 VN.n27 VSUBS 0.030941f
C606 VN.n28 VSUBS 0.061013f
C607 VN.n29 VSUBS 0.057377f
C608 VN.n30 VSUBS 0.029618f
C609 VN.n31 VSUBS 0.030941f
C610 VN.n32 VSUBS 0.030941f
C611 VN.n33 VSUBS 0.056811f
C612 VN.n34 VSUBS 0.061586f
C613 VN.n35 VSUBS 0.025079f
C614 VN.n36 VSUBS 0.030941f
C615 VN.n37 VSUBS 0.030941f
C616 VN.n38 VSUBS 0.030941f
C617 VN.n39 VSUBS 0.057377f
C618 VN.n40 VSUBS 0.030185f
C619 VN.n41 VSUBS 0.781604f
C620 VN.n42 VSUBS 0.05729f
C621 VN.n43 VSUBS 0.04079f
C622 VN.t4 VSUBS 1.90712f
C623 VN.n44 VSUBS 0.060668f
C624 VN.n45 VSUBS 0.030941f
C625 VN.t1 VSUBS 1.90712f
C626 VN.n46 VSUBS 0.689853f
C627 VN.n47 VSUBS 0.030941f
C628 VN.n48 VSUBS 0.025f
C629 VN.n49 VSUBS 0.030941f
C630 VN.t5 VSUBS 1.90712f
C631 VN.n50 VSUBS 0.057377f
C632 VN.n51 VSUBS 0.030941f
C633 VN.n52 VSUBS 0.057377f
C634 VN.t3 VSUBS 2.15648f
C635 VN.n53 VSUBS 0.760711f
C636 VN.t9 VSUBS 1.90712f
C637 VN.n54 VSUBS 0.769432f
C638 VN.n55 VSUBS 0.029618f
C639 VN.n56 VSUBS 0.300667f
C640 VN.n57 VSUBS 0.030941f
C641 VN.n58 VSUBS 0.030941f
C642 VN.n59 VSUBS 0.061013f
C643 VN.n60 VSUBS 0.025f
C644 VN.n61 VSUBS 0.06132f
C645 VN.n62 VSUBS 0.030941f
C646 VN.n63 VSUBS 0.030941f
C647 VN.n64 VSUBS 0.030941f
C648 VN.n65 VSUBS 0.718905f
C649 VN.n66 VSUBS 0.057377f
C650 VN.n67 VSUBS 0.06132f
C651 VN.n68 VSUBS 0.030941f
C652 VN.n69 VSUBS 0.030941f
C653 VN.n70 VSUBS 0.030941f
C654 VN.n71 VSUBS 0.061013f
C655 VN.n72 VSUBS 0.057377f
C656 VN.n73 VSUBS 0.029618f
C657 VN.n74 VSUBS 0.030941f
C658 VN.n75 VSUBS 0.030941f
C659 VN.n76 VSUBS 0.056811f
C660 VN.n77 VSUBS 0.061586f
C661 VN.n78 VSUBS 0.025079f
C662 VN.n79 VSUBS 0.030941f
C663 VN.n80 VSUBS 0.030941f
C664 VN.n81 VSUBS 0.030941f
C665 VN.n82 VSUBS 0.057377f
C666 VN.n83 VSUBS 0.030185f
C667 VN.n84 VSUBS 0.781604f
C668 VN.n85 VSUBS 1.78583f
C669 B.n0 VSUBS 0.006632f
C670 B.n1 VSUBS 0.006632f
C671 B.n2 VSUBS 0.010488f
C672 B.n3 VSUBS 0.010488f
C673 B.n4 VSUBS 0.010488f
C674 B.n5 VSUBS 0.010488f
C675 B.n6 VSUBS 0.010488f
C676 B.n7 VSUBS 0.010488f
C677 B.n8 VSUBS 0.010488f
C678 B.n9 VSUBS 0.010488f
C679 B.n10 VSUBS 0.010488f
C680 B.n11 VSUBS 0.010488f
C681 B.n12 VSUBS 0.010488f
C682 B.n13 VSUBS 0.010488f
C683 B.n14 VSUBS 0.010488f
C684 B.n15 VSUBS 0.010488f
C685 B.n16 VSUBS 0.010488f
C686 B.n17 VSUBS 0.010488f
C687 B.n18 VSUBS 0.010488f
C688 B.n19 VSUBS 0.010488f
C689 B.n20 VSUBS 0.010488f
C690 B.n21 VSUBS 0.010488f
C691 B.n22 VSUBS 0.010488f
C692 B.n23 VSUBS 0.010488f
C693 B.n24 VSUBS 0.010488f
C694 B.n25 VSUBS 0.010488f
C695 B.n26 VSUBS 0.010488f
C696 B.n27 VSUBS 0.010488f
C697 B.n28 VSUBS 0.010488f
C698 B.n29 VSUBS 0.010488f
C699 B.n30 VSUBS 0.010488f
C700 B.n31 VSUBS 0.010488f
C701 B.n32 VSUBS 0.026321f
C702 B.n33 VSUBS 0.010488f
C703 B.n34 VSUBS 0.010488f
C704 B.n35 VSUBS 0.010488f
C705 B.n36 VSUBS 0.010488f
C706 B.n37 VSUBS 0.010488f
C707 B.n38 VSUBS 0.010488f
C708 B.n39 VSUBS 0.010488f
C709 B.n40 VSUBS 0.010488f
C710 B.n41 VSUBS 0.010488f
C711 B.n42 VSUBS 0.010488f
C712 B.n43 VSUBS 0.010488f
C713 B.n44 VSUBS 0.010488f
C714 B.n45 VSUBS 0.010488f
C715 B.n46 VSUBS 0.010488f
C716 B.n47 VSUBS 0.010488f
C717 B.t11 VSUBS 0.205487f
C718 B.t10 VSUBS 0.250439f
C719 B.t9 VSUBS 1.59604f
C720 B.n48 VSUBS 0.412641f
C721 B.n49 VSUBS 0.301075f
C722 B.n50 VSUBS 0.0243f
C723 B.n51 VSUBS 0.010488f
C724 B.n52 VSUBS 0.010488f
C725 B.n53 VSUBS 0.010488f
C726 B.n54 VSUBS 0.010488f
C727 B.n55 VSUBS 0.010488f
C728 B.t2 VSUBS 0.205491f
C729 B.t1 VSUBS 0.250442f
C730 B.t0 VSUBS 1.59604f
C731 B.n56 VSUBS 0.412638f
C732 B.n57 VSUBS 0.301071f
C733 B.n58 VSUBS 0.010488f
C734 B.n59 VSUBS 0.010488f
C735 B.n60 VSUBS 0.010488f
C736 B.n61 VSUBS 0.010488f
C737 B.n62 VSUBS 0.010488f
C738 B.n63 VSUBS 0.010488f
C739 B.n64 VSUBS 0.010488f
C740 B.n65 VSUBS 0.010488f
C741 B.n66 VSUBS 0.010488f
C742 B.n67 VSUBS 0.010488f
C743 B.n68 VSUBS 0.010488f
C744 B.n69 VSUBS 0.010488f
C745 B.n70 VSUBS 0.010488f
C746 B.n71 VSUBS 0.010488f
C747 B.n72 VSUBS 0.010488f
C748 B.n73 VSUBS 0.026321f
C749 B.n74 VSUBS 0.010488f
C750 B.n75 VSUBS 0.010488f
C751 B.n76 VSUBS 0.010488f
C752 B.n77 VSUBS 0.010488f
C753 B.n78 VSUBS 0.010488f
C754 B.n79 VSUBS 0.010488f
C755 B.n80 VSUBS 0.010488f
C756 B.n81 VSUBS 0.010488f
C757 B.n82 VSUBS 0.010488f
C758 B.n83 VSUBS 0.010488f
C759 B.n84 VSUBS 0.010488f
C760 B.n85 VSUBS 0.010488f
C761 B.n86 VSUBS 0.010488f
C762 B.n87 VSUBS 0.010488f
C763 B.n88 VSUBS 0.010488f
C764 B.n89 VSUBS 0.010488f
C765 B.n90 VSUBS 0.010488f
C766 B.n91 VSUBS 0.010488f
C767 B.n92 VSUBS 0.010488f
C768 B.n93 VSUBS 0.010488f
C769 B.n94 VSUBS 0.010488f
C770 B.n95 VSUBS 0.010488f
C771 B.n96 VSUBS 0.010488f
C772 B.n97 VSUBS 0.010488f
C773 B.n98 VSUBS 0.010488f
C774 B.n99 VSUBS 0.010488f
C775 B.n100 VSUBS 0.010488f
C776 B.n101 VSUBS 0.010488f
C777 B.n102 VSUBS 0.010488f
C778 B.n103 VSUBS 0.010488f
C779 B.n104 VSUBS 0.010488f
C780 B.n105 VSUBS 0.010488f
C781 B.n106 VSUBS 0.010488f
C782 B.n107 VSUBS 0.010488f
C783 B.n108 VSUBS 0.010488f
C784 B.n109 VSUBS 0.010488f
C785 B.n110 VSUBS 0.010488f
C786 B.n111 VSUBS 0.010488f
C787 B.n112 VSUBS 0.010488f
C788 B.n113 VSUBS 0.010488f
C789 B.n114 VSUBS 0.010488f
C790 B.n115 VSUBS 0.010488f
C791 B.n116 VSUBS 0.010488f
C792 B.n117 VSUBS 0.010488f
C793 B.n118 VSUBS 0.010488f
C794 B.n119 VSUBS 0.010488f
C795 B.n120 VSUBS 0.010488f
C796 B.n121 VSUBS 0.010488f
C797 B.n122 VSUBS 0.010488f
C798 B.n123 VSUBS 0.010488f
C799 B.n124 VSUBS 0.010488f
C800 B.n125 VSUBS 0.010488f
C801 B.n126 VSUBS 0.010488f
C802 B.n127 VSUBS 0.010488f
C803 B.n128 VSUBS 0.010488f
C804 B.n129 VSUBS 0.010488f
C805 B.n130 VSUBS 0.010488f
C806 B.n131 VSUBS 0.010488f
C807 B.n132 VSUBS 0.010488f
C808 B.n133 VSUBS 0.010488f
C809 B.n134 VSUBS 0.026321f
C810 B.n135 VSUBS 0.010488f
C811 B.n136 VSUBS 0.010488f
C812 B.n137 VSUBS 0.010488f
C813 B.n138 VSUBS 0.010488f
C814 B.n139 VSUBS 0.010488f
C815 B.n140 VSUBS 0.010488f
C816 B.n141 VSUBS 0.010488f
C817 B.n142 VSUBS 0.010488f
C818 B.n143 VSUBS 0.010488f
C819 B.n144 VSUBS 0.010488f
C820 B.n145 VSUBS 0.010488f
C821 B.n146 VSUBS 0.010488f
C822 B.n147 VSUBS 0.010488f
C823 B.n148 VSUBS 0.010488f
C824 B.n149 VSUBS 0.010488f
C825 B.t7 VSUBS 0.205491f
C826 B.t8 VSUBS 0.250442f
C827 B.t6 VSUBS 1.59604f
C828 B.n150 VSUBS 0.412638f
C829 B.n151 VSUBS 0.301071f
C830 B.n152 VSUBS 0.0243f
C831 B.n153 VSUBS 0.010488f
C832 B.n154 VSUBS 0.010488f
C833 B.n155 VSUBS 0.010488f
C834 B.n156 VSUBS 0.010488f
C835 B.n157 VSUBS 0.010488f
C836 B.t4 VSUBS 0.205487f
C837 B.t5 VSUBS 0.250439f
C838 B.t3 VSUBS 1.59604f
C839 B.n158 VSUBS 0.412641f
C840 B.n159 VSUBS 0.301075f
C841 B.n160 VSUBS 0.010488f
C842 B.n161 VSUBS 0.010488f
C843 B.n162 VSUBS 0.010488f
C844 B.n163 VSUBS 0.010488f
C845 B.n164 VSUBS 0.010488f
C846 B.n165 VSUBS 0.010488f
C847 B.n166 VSUBS 0.010488f
C848 B.n167 VSUBS 0.010488f
C849 B.n168 VSUBS 0.010488f
C850 B.n169 VSUBS 0.010488f
C851 B.n170 VSUBS 0.010488f
C852 B.n171 VSUBS 0.010488f
C853 B.n172 VSUBS 0.010488f
C854 B.n173 VSUBS 0.010488f
C855 B.n174 VSUBS 0.010488f
C856 B.n175 VSUBS 0.026321f
C857 B.n176 VSUBS 0.010488f
C858 B.n177 VSUBS 0.010488f
C859 B.n178 VSUBS 0.010488f
C860 B.n179 VSUBS 0.010488f
C861 B.n180 VSUBS 0.010488f
C862 B.n181 VSUBS 0.010488f
C863 B.n182 VSUBS 0.010488f
C864 B.n183 VSUBS 0.010488f
C865 B.n184 VSUBS 0.010488f
C866 B.n185 VSUBS 0.010488f
C867 B.n186 VSUBS 0.010488f
C868 B.n187 VSUBS 0.010488f
C869 B.n188 VSUBS 0.010488f
C870 B.n189 VSUBS 0.010488f
C871 B.n190 VSUBS 0.010488f
C872 B.n191 VSUBS 0.010488f
C873 B.n192 VSUBS 0.010488f
C874 B.n193 VSUBS 0.010488f
C875 B.n194 VSUBS 0.010488f
C876 B.n195 VSUBS 0.010488f
C877 B.n196 VSUBS 0.010488f
C878 B.n197 VSUBS 0.010488f
C879 B.n198 VSUBS 0.010488f
C880 B.n199 VSUBS 0.010488f
C881 B.n200 VSUBS 0.010488f
C882 B.n201 VSUBS 0.010488f
C883 B.n202 VSUBS 0.010488f
C884 B.n203 VSUBS 0.010488f
C885 B.n204 VSUBS 0.010488f
C886 B.n205 VSUBS 0.010488f
C887 B.n206 VSUBS 0.010488f
C888 B.n207 VSUBS 0.010488f
C889 B.n208 VSUBS 0.010488f
C890 B.n209 VSUBS 0.010488f
C891 B.n210 VSUBS 0.010488f
C892 B.n211 VSUBS 0.010488f
C893 B.n212 VSUBS 0.010488f
C894 B.n213 VSUBS 0.010488f
C895 B.n214 VSUBS 0.010488f
C896 B.n215 VSUBS 0.010488f
C897 B.n216 VSUBS 0.010488f
C898 B.n217 VSUBS 0.010488f
C899 B.n218 VSUBS 0.010488f
C900 B.n219 VSUBS 0.010488f
C901 B.n220 VSUBS 0.010488f
C902 B.n221 VSUBS 0.010488f
C903 B.n222 VSUBS 0.010488f
C904 B.n223 VSUBS 0.010488f
C905 B.n224 VSUBS 0.010488f
C906 B.n225 VSUBS 0.010488f
C907 B.n226 VSUBS 0.010488f
C908 B.n227 VSUBS 0.010488f
C909 B.n228 VSUBS 0.010488f
C910 B.n229 VSUBS 0.010488f
C911 B.n230 VSUBS 0.010488f
C912 B.n231 VSUBS 0.010488f
C913 B.n232 VSUBS 0.010488f
C914 B.n233 VSUBS 0.010488f
C915 B.n234 VSUBS 0.010488f
C916 B.n235 VSUBS 0.010488f
C917 B.n236 VSUBS 0.010488f
C918 B.n237 VSUBS 0.010488f
C919 B.n238 VSUBS 0.010488f
C920 B.n239 VSUBS 0.010488f
C921 B.n240 VSUBS 0.010488f
C922 B.n241 VSUBS 0.010488f
C923 B.n242 VSUBS 0.010488f
C924 B.n243 VSUBS 0.010488f
C925 B.n244 VSUBS 0.010488f
C926 B.n245 VSUBS 0.010488f
C927 B.n246 VSUBS 0.010488f
C928 B.n247 VSUBS 0.010488f
C929 B.n248 VSUBS 0.010488f
C930 B.n249 VSUBS 0.010488f
C931 B.n250 VSUBS 0.010488f
C932 B.n251 VSUBS 0.010488f
C933 B.n252 VSUBS 0.010488f
C934 B.n253 VSUBS 0.010488f
C935 B.n254 VSUBS 0.010488f
C936 B.n255 VSUBS 0.010488f
C937 B.n256 VSUBS 0.010488f
C938 B.n257 VSUBS 0.010488f
C939 B.n258 VSUBS 0.010488f
C940 B.n259 VSUBS 0.010488f
C941 B.n260 VSUBS 0.010488f
C942 B.n261 VSUBS 0.010488f
C943 B.n262 VSUBS 0.010488f
C944 B.n263 VSUBS 0.010488f
C945 B.n264 VSUBS 0.010488f
C946 B.n265 VSUBS 0.010488f
C947 B.n266 VSUBS 0.010488f
C948 B.n267 VSUBS 0.010488f
C949 B.n268 VSUBS 0.010488f
C950 B.n269 VSUBS 0.010488f
C951 B.n270 VSUBS 0.010488f
C952 B.n271 VSUBS 0.010488f
C953 B.n272 VSUBS 0.010488f
C954 B.n273 VSUBS 0.010488f
C955 B.n274 VSUBS 0.010488f
C956 B.n275 VSUBS 0.010488f
C957 B.n276 VSUBS 0.010488f
C958 B.n277 VSUBS 0.010488f
C959 B.n278 VSUBS 0.010488f
C960 B.n279 VSUBS 0.010488f
C961 B.n280 VSUBS 0.010488f
C962 B.n281 VSUBS 0.010488f
C963 B.n282 VSUBS 0.010488f
C964 B.n283 VSUBS 0.010488f
C965 B.n284 VSUBS 0.010488f
C966 B.n285 VSUBS 0.010488f
C967 B.n286 VSUBS 0.010488f
C968 B.n287 VSUBS 0.010488f
C969 B.n288 VSUBS 0.010488f
C970 B.n289 VSUBS 0.010488f
C971 B.n290 VSUBS 0.010488f
C972 B.n291 VSUBS 0.010488f
C973 B.n292 VSUBS 0.010488f
C974 B.n293 VSUBS 0.010488f
C975 B.n294 VSUBS 0.026321f
C976 B.n295 VSUBS 0.027353f
C977 B.n296 VSUBS 0.027353f
C978 B.n297 VSUBS 0.010488f
C979 B.n298 VSUBS 0.010488f
C980 B.n299 VSUBS 0.010488f
C981 B.n300 VSUBS 0.010488f
C982 B.n301 VSUBS 0.010488f
C983 B.n302 VSUBS 0.010488f
C984 B.n303 VSUBS 0.010488f
C985 B.n304 VSUBS 0.010488f
C986 B.n305 VSUBS 0.010488f
C987 B.n306 VSUBS 0.010488f
C988 B.n307 VSUBS 0.010488f
C989 B.n308 VSUBS 0.010488f
C990 B.n309 VSUBS 0.010488f
C991 B.n310 VSUBS 0.010488f
C992 B.n311 VSUBS 0.010488f
C993 B.n312 VSUBS 0.010488f
C994 B.n313 VSUBS 0.010488f
C995 B.n314 VSUBS 0.010488f
C996 B.n315 VSUBS 0.010488f
C997 B.n316 VSUBS 0.010488f
C998 B.n317 VSUBS 0.010488f
C999 B.n318 VSUBS 0.010488f
C1000 B.n319 VSUBS 0.010488f
C1001 B.n320 VSUBS 0.010488f
C1002 B.n321 VSUBS 0.010488f
C1003 B.n322 VSUBS 0.010488f
C1004 B.n323 VSUBS 0.010488f
C1005 B.n324 VSUBS 0.010488f
C1006 B.n325 VSUBS 0.010488f
C1007 B.n326 VSUBS 0.010488f
C1008 B.n327 VSUBS 0.010488f
C1009 B.n328 VSUBS 0.010488f
C1010 B.n329 VSUBS 0.010488f
C1011 B.n330 VSUBS 0.010488f
C1012 B.n331 VSUBS 0.010488f
C1013 B.n332 VSUBS 0.010488f
C1014 B.n333 VSUBS 0.010488f
C1015 B.n334 VSUBS 0.010488f
C1016 B.n335 VSUBS 0.010488f
C1017 B.n336 VSUBS 0.010488f
C1018 B.n337 VSUBS 0.010488f
C1019 B.n338 VSUBS 0.010488f
C1020 B.n339 VSUBS 0.010488f
C1021 B.n340 VSUBS 0.010488f
C1022 B.n341 VSUBS 0.009871f
C1023 B.n342 VSUBS 0.0243f
C1024 B.n343 VSUBS 0.005861f
C1025 B.n344 VSUBS 0.010488f
C1026 B.n345 VSUBS 0.010488f
C1027 B.n346 VSUBS 0.010488f
C1028 B.n347 VSUBS 0.010488f
C1029 B.n348 VSUBS 0.010488f
C1030 B.n349 VSUBS 0.010488f
C1031 B.n350 VSUBS 0.010488f
C1032 B.n351 VSUBS 0.010488f
C1033 B.n352 VSUBS 0.010488f
C1034 B.n353 VSUBS 0.010488f
C1035 B.n354 VSUBS 0.010488f
C1036 B.n355 VSUBS 0.010488f
C1037 B.n356 VSUBS 0.005861f
C1038 B.n357 VSUBS 0.010488f
C1039 B.n358 VSUBS 0.010488f
C1040 B.n359 VSUBS 0.009871f
C1041 B.n360 VSUBS 0.010488f
C1042 B.n361 VSUBS 0.010488f
C1043 B.n362 VSUBS 0.010488f
C1044 B.n363 VSUBS 0.010488f
C1045 B.n364 VSUBS 0.010488f
C1046 B.n365 VSUBS 0.010488f
C1047 B.n366 VSUBS 0.010488f
C1048 B.n367 VSUBS 0.010488f
C1049 B.n368 VSUBS 0.010488f
C1050 B.n369 VSUBS 0.010488f
C1051 B.n370 VSUBS 0.010488f
C1052 B.n371 VSUBS 0.010488f
C1053 B.n372 VSUBS 0.010488f
C1054 B.n373 VSUBS 0.010488f
C1055 B.n374 VSUBS 0.010488f
C1056 B.n375 VSUBS 0.010488f
C1057 B.n376 VSUBS 0.010488f
C1058 B.n377 VSUBS 0.010488f
C1059 B.n378 VSUBS 0.010488f
C1060 B.n379 VSUBS 0.010488f
C1061 B.n380 VSUBS 0.010488f
C1062 B.n381 VSUBS 0.010488f
C1063 B.n382 VSUBS 0.010488f
C1064 B.n383 VSUBS 0.010488f
C1065 B.n384 VSUBS 0.010488f
C1066 B.n385 VSUBS 0.010488f
C1067 B.n386 VSUBS 0.010488f
C1068 B.n387 VSUBS 0.010488f
C1069 B.n388 VSUBS 0.010488f
C1070 B.n389 VSUBS 0.010488f
C1071 B.n390 VSUBS 0.010488f
C1072 B.n391 VSUBS 0.010488f
C1073 B.n392 VSUBS 0.010488f
C1074 B.n393 VSUBS 0.010488f
C1075 B.n394 VSUBS 0.010488f
C1076 B.n395 VSUBS 0.010488f
C1077 B.n396 VSUBS 0.010488f
C1078 B.n397 VSUBS 0.010488f
C1079 B.n398 VSUBS 0.010488f
C1080 B.n399 VSUBS 0.010488f
C1081 B.n400 VSUBS 0.010488f
C1082 B.n401 VSUBS 0.010488f
C1083 B.n402 VSUBS 0.010488f
C1084 B.n403 VSUBS 0.027353f
C1085 B.n404 VSUBS 0.027353f
C1086 B.n405 VSUBS 0.026321f
C1087 B.n406 VSUBS 0.010488f
C1088 B.n407 VSUBS 0.010488f
C1089 B.n408 VSUBS 0.010488f
C1090 B.n409 VSUBS 0.010488f
C1091 B.n410 VSUBS 0.010488f
C1092 B.n411 VSUBS 0.010488f
C1093 B.n412 VSUBS 0.010488f
C1094 B.n413 VSUBS 0.010488f
C1095 B.n414 VSUBS 0.010488f
C1096 B.n415 VSUBS 0.010488f
C1097 B.n416 VSUBS 0.010488f
C1098 B.n417 VSUBS 0.010488f
C1099 B.n418 VSUBS 0.010488f
C1100 B.n419 VSUBS 0.010488f
C1101 B.n420 VSUBS 0.010488f
C1102 B.n421 VSUBS 0.010488f
C1103 B.n422 VSUBS 0.010488f
C1104 B.n423 VSUBS 0.010488f
C1105 B.n424 VSUBS 0.010488f
C1106 B.n425 VSUBS 0.010488f
C1107 B.n426 VSUBS 0.010488f
C1108 B.n427 VSUBS 0.010488f
C1109 B.n428 VSUBS 0.010488f
C1110 B.n429 VSUBS 0.010488f
C1111 B.n430 VSUBS 0.010488f
C1112 B.n431 VSUBS 0.010488f
C1113 B.n432 VSUBS 0.010488f
C1114 B.n433 VSUBS 0.010488f
C1115 B.n434 VSUBS 0.010488f
C1116 B.n435 VSUBS 0.010488f
C1117 B.n436 VSUBS 0.010488f
C1118 B.n437 VSUBS 0.010488f
C1119 B.n438 VSUBS 0.010488f
C1120 B.n439 VSUBS 0.010488f
C1121 B.n440 VSUBS 0.010488f
C1122 B.n441 VSUBS 0.010488f
C1123 B.n442 VSUBS 0.010488f
C1124 B.n443 VSUBS 0.010488f
C1125 B.n444 VSUBS 0.010488f
C1126 B.n445 VSUBS 0.010488f
C1127 B.n446 VSUBS 0.010488f
C1128 B.n447 VSUBS 0.010488f
C1129 B.n448 VSUBS 0.010488f
C1130 B.n449 VSUBS 0.010488f
C1131 B.n450 VSUBS 0.010488f
C1132 B.n451 VSUBS 0.010488f
C1133 B.n452 VSUBS 0.010488f
C1134 B.n453 VSUBS 0.010488f
C1135 B.n454 VSUBS 0.010488f
C1136 B.n455 VSUBS 0.010488f
C1137 B.n456 VSUBS 0.010488f
C1138 B.n457 VSUBS 0.010488f
C1139 B.n458 VSUBS 0.010488f
C1140 B.n459 VSUBS 0.010488f
C1141 B.n460 VSUBS 0.010488f
C1142 B.n461 VSUBS 0.010488f
C1143 B.n462 VSUBS 0.010488f
C1144 B.n463 VSUBS 0.010488f
C1145 B.n464 VSUBS 0.010488f
C1146 B.n465 VSUBS 0.010488f
C1147 B.n466 VSUBS 0.010488f
C1148 B.n467 VSUBS 0.010488f
C1149 B.n468 VSUBS 0.010488f
C1150 B.n469 VSUBS 0.010488f
C1151 B.n470 VSUBS 0.010488f
C1152 B.n471 VSUBS 0.010488f
C1153 B.n472 VSUBS 0.010488f
C1154 B.n473 VSUBS 0.010488f
C1155 B.n474 VSUBS 0.010488f
C1156 B.n475 VSUBS 0.010488f
C1157 B.n476 VSUBS 0.010488f
C1158 B.n477 VSUBS 0.010488f
C1159 B.n478 VSUBS 0.010488f
C1160 B.n479 VSUBS 0.010488f
C1161 B.n480 VSUBS 0.010488f
C1162 B.n481 VSUBS 0.010488f
C1163 B.n482 VSUBS 0.010488f
C1164 B.n483 VSUBS 0.010488f
C1165 B.n484 VSUBS 0.010488f
C1166 B.n485 VSUBS 0.010488f
C1167 B.n486 VSUBS 0.010488f
C1168 B.n487 VSUBS 0.010488f
C1169 B.n488 VSUBS 0.010488f
C1170 B.n489 VSUBS 0.010488f
C1171 B.n490 VSUBS 0.010488f
C1172 B.n491 VSUBS 0.010488f
C1173 B.n492 VSUBS 0.010488f
C1174 B.n493 VSUBS 0.010488f
C1175 B.n494 VSUBS 0.010488f
C1176 B.n495 VSUBS 0.010488f
C1177 B.n496 VSUBS 0.010488f
C1178 B.n497 VSUBS 0.010488f
C1179 B.n498 VSUBS 0.010488f
C1180 B.n499 VSUBS 0.010488f
C1181 B.n500 VSUBS 0.010488f
C1182 B.n501 VSUBS 0.010488f
C1183 B.n502 VSUBS 0.010488f
C1184 B.n503 VSUBS 0.010488f
C1185 B.n504 VSUBS 0.010488f
C1186 B.n505 VSUBS 0.010488f
C1187 B.n506 VSUBS 0.010488f
C1188 B.n507 VSUBS 0.010488f
C1189 B.n508 VSUBS 0.010488f
C1190 B.n509 VSUBS 0.010488f
C1191 B.n510 VSUBS 0.010488f
C1192 B.n511 VSUBS 0.010488f
C1193 B.n512 VSUBS 0.010488f
C1194 B.n513 VSUBS 0.010488f
C1195 B.n514 VSUBS 0.010488f
C1196 B.n515 VSUBS 0.010488f
C1197 B.n516 VSUBS 0.010488f
C1198 B.n517 VSUBS 0.010488f
C1199 B.n518 VSUBS 0.010488f
C1200 B.n519 VSUBS 0.010488f
C1201 B.n520 VSUBS 0.010488f
C1202 B.n521 VSUBS 0.010488f
C1203 B.n522 VSUBS 0.010488f
C1204 B.n523 VSUBS 0.010488f
C1205 B.n524 VSUBS 0.010488f
C1206 B.n525 VSUBS 0.010488f
C1207 B.n526 VSUBS 0.010488f
C1208 B.n527 VSUBS 0.010488f
C1209 B.n528 VSUBS 0.010488f
C1210 B.n529 VSUBS 0.010488f
C1211 B.n530 VSUBS 0.010488f
C1212 B.n531 VSUBS 0.010488f
C1213 B.n532 VSUBS 0.010488f
C1214 B.n533 VSUBS 0.010488f
C1215 B.n534 VSUBS 0.010488f
C1216 B.n535 VSUBS 0.010488f
C1217 B.n536 VSUBS 0.010488f
C1218 B.n537 VSUBS 0.010488f
C1219 B.n538 VSUBS 0.010488f
C1220 B.n539 VSUBS 0.010488f
C1221 B.n540 VSUBS 0.010488f
C1222 B.n541 VSUBS 0.010488f
C1223 B.n542 VSUBS 0.010488f
C1224 B.n543 VSUBS 0.010488f
C1225 B.n544 VSUBS 0.010488f
C1226 B.n545 VSUBS 0.010488f
C1227 B.n546 VSUBS 0.010488f
C1228 B.n547 VSUBS 0.010488f
C1229 B.n548 VSUBS 0.010488f
C1230 B.n549 VSUBS 0.010488f
C1231 B.n550 VSUBS 0.010488f
C1232 B.n551 VSUBS 0.010488f
C1233 B.n552 VSUBS 0.010488f
C1234 B.n553 VSUBS 0.010488f
C1235 B.n554 VSUBS 0.010488f
C1236 B.n555 VSUBS 0.010488f
C1237 B.n556 VSUBS 0.010488f
C1238 B.n557 VSUBS 0.010488f
C1239 B.n558 VSUBS 0.010488f
C1240 B.n559 VSUBS 0.010488f
C1241 B.n560 VSUBS 0.010488f
C1242 B.n561 VSUBS 0.010488f
C1243 B.n562 VSUBS 0.010488f
C1244 B.n563 VSUBS 0.010488f
C1245 B.n564 VSUBS 0.010488f
C1246 B.n565 VSUBS 0.010488f
C1247 B.n566 VSUBS 0.010488f
C1248 B.n567 VSUBS 0.010488f
C1249 B.n568 VSUBS 0.010488f
C1250 B.n569 VSUBS 0.010488f
C1251 B.n570 VSUBS 0.010488f
C1252 B.n571 VSUBS 0.010488f
C1253 B.n572 VSUBS 0.010488f
C1254 B.n573 VSUBS 0.010488f
C1255 B.n574 VSUBS 0.010488f
C1256 B.n575 VSUBS 0.010488f
C1257 B.n576 VSUBS 0.010488f
C1258 B.n577 VSUBS 0.010488f
C1259 B.n578 VSUBS 0.010488f
C1260 B.n579 VSUBS 0.010488f
C1261 B.n580 VSUBS 0.010488f
C1262 B.n581 VSUBS 0.010488f
C1263 B.n582 VSUBS 0.010488f
C1264 B.n583 VSUBS 0.010488f
C1265 B.n584 VSUBS 0.010488f
C1266 B.n585 VSUBS 0.010488f
C1267 B.n586 VSUBS 0.010488f
C1268 B.n587 VSUBS 0.010488f
C1269 B.n588 VSUBS 0.027406f
C1270 B.n589 VSUBS 0.026268f
C1271 B.n590 VSUBS 0.027353f
C1272 B.n591 VSUBS 0.010488f
C1273 B.n592 VSUBS 0.010488f
C1274 B.n593 VSUBS 0.010488f
C1275 B.n594 VSUBS 0.010488f
C1276 B.n595 VSUBS 0.010488f
C1277 B.n596 VSUBS 0.010488f
C1278 B.n597 VSUBS 0.010488f
C1279 B.n598 VSUBS 0.010488f
C1280 B.n599 VSUBS 0.010488f
C1281 B.n600 VSUBS 0.010488f
C1282 B.n601 VSUBS 0.010488f
C1283 B.n602 VSUBS 0.010488f
C1284 B.n603 VSUBS 0.010488f
C1285 B.n604 VSUBS 0.010488f
C1286 B.n605 VSUBS 0.010488f
C1287 B.n606 VSUBS 0.010488f
C1288 B.n607 VSUBS 0.010488f
C1289 B.n608 VSUBS 0.010488f
C1290 B.n609 VSUBS 0.010488f
C1291 B.n610 VSUBS 0.010488f
C1292 B.n611 VSUBS 0.010488f
C1293 B.n612 VSUBS 0.010488f
C1294 B.n613 VSUBS 0.010488f
C1295 B.n614 VSUBS 0.010488f
C1296 B.n615 VSUBS 0.010488f
C1297 B.n616 VSUBS 0.010488f
C1298 B.n617 VSUBS 0.010488f
C1299 B.n618 VSUBS 0.010488f
C1300 B.n619 VSUBS 0.010488f
C1301 B.n620 VSUBS 0.010488f
C1302 B.n621 VSUBS 0.010488f
C1303 B.n622 VSUBS 0.010488f
C1304 B.n623 VSUBS 0.010488f
C1305 B.n624 VSUBS 0.010488f
C1306 B.n625 VSUBS 0.010488f
C1307 B.n626 VSUBS 0.010488f
C1308 B.n627 VSUBS 0.010488f
C1309 B.n628 VSUBS 0.010488f
C1310 B.n629 VSUBS 0.010488f
C1311 B.n630 VSUBS 0.010488f
C1312 B.n631 VSUBS 0.010488f
C1313 B.n632 VSUBS 0.010488f
C1314 B.n633 VSUBS 0.010488f
C1315 B.n634 VSUBS 0.010488f
C1316 B.n635 VSUBS 0.009871f
C1317 B.n636 VSUBS 0.0243f
C1318 B.n637 VSUBS 0.005861f
C1319 B.n638 VSUBS 0.010488f
C1320 B.n639 VSUBS 0.010488f
C1321 B.n640 VSUBS 0.010488f
C1322 B.n641 VSUBS 0.010488f
C1323 B.n642 VSUBS 0.010488f
C1324 B.n643 VSUBS 0.010488f
C1325 B.n644 VSUBS 0.010488f
C1326 B.n645 VSUBS 0.010488f
C1327 B.n646 VSUBS 0.010488f
C1328 B.n647 VSUBS 0.010488f
C1329 B.n648 VSUBS 0.010488f
C1330 B.n649 VSUBS 0.010488f
C1331 B.n650 VSUBS 0.005861f
C1332 B.n651 VSUBS 0.010488f
C1333 B.n652 VSUBS 0.010488f
C1334 B.n653 VSUBS 0.009871f
C1335 B.n654 VSUBS 0.010488f
C1336 B.n655 VSUBS 0.010488f
C1337 B.n656 VSUBS 0.010488f
C1338 B.n657 VSUBS 0.010488f
C1339 B.n658 VSUBS 0.010488f
C1340 B.n659 VSUBS 0.010488f
C1341 B.n660 VSUBS 0.010488f
C1342 B.n661 VSUBS 0.010488f
C1343 B.n662 VSUBS 0.010488f
C1344 B.n663 VSUBS 0.010488f
C1345 B.n664 VSUBS 0.010488f
C1346 B.n665 VSUBS 0.010488f
C1347 B.n666 VSUBS 0.010488f
C1348 B.n667 VSUBS 0.010488f
C1349 B.n668 VSUBS 0.010488f
C1350 B.n669 VSUBS 0.010488f
C1351 B.n670 VSUBS 0.010488f
C1352 B.n671 VSUBS 0.010488f
C1353 B.n672 VSUBS 0.010488f
C1354 B.n673 VSUBS 0.010488f
C1355 B.n674 VSUBS 0.010488f
C1356 B.n675 VSUBS 0.010488f
C1357 B.n676 VSUBS 0.010488f
C1358 B.n677 VSUBS 0.010488f
C1359 B.n678 VSUBS 0.010488f
C1360 B.n679 VSUBS 0.010488f
C1361 B.n680 VSUBS 0.010488f
C1362 B.n681 VSUBS 0.010488f
C1363 B.n682 VSUBS 0.010488f
C1364 B.n683 VSUBS 0.010488f
C1365 B.n684 VSUBS 0.010488f
C1366 B.n685 VSUBS 0.010488f
C1367 B.n686 VSUBS 0.010488f
C1368 B.n687 VSUBS 0.010488f
C1369 B.n688 VSUBS 0.010488f
C1370 B.n689 VSUBS 0.010488f
C1371 B.n690 VSUBS 0.010488f
C1372 B.n691 VSUBS 0.010488f
C1373 B.n692 VSUBS 0.010488f
C1374 B.n693 VSUBS 0.010488f
C1375 B.n694 VSUBS 0.010488f
C1376 B.n695 VSUBS 0.010488f
C1377 B.n696 VSUBS 0.010488f
C1378 B.n697 VSUBS 0.027353f
C1379 B.n698 VSUBS 0.027353f
C1380 B.n699 VSUBS 0.026321f
C1381 B.n700 VSUBS 0.010488f
C1382 B.n701 VSUBS 0.010488f
C1383 B.n702 VSUBS 0.010488f
C1384 B.n703 VSUBS 0.010488f
C1385 B.n704 VSUBS 0.010488f
C1386 B.n705 VSUBS 0.010488f
C1387 B.n706 VSUBS 0.010488f
C1388 B.n707 VSUBS 0.010488f
C1389 B.n708 VSUBS 0.010488f
C1390 B.n709 VSUBS 0.010488f
C1391 B.n710 VSUBS 0.010488f
C1392 B.n711 VSUBS 0.010488f
C1393 B.n712 VSUBS 0.010488f
C1394 B.n713 VSUBS 0.010488f
C1395 B.n714 VSUBS 0.010488f
C1396 B.n715 VSUBS 0.010488f
C1397 B.n716 VSUBS 0.010488f
C1398 B.n717 VSUBS 0.010488f
C1399 B.n718 VSUBS 0.010488f
C1400 B.n719 VSUBS 0.010488f
C1401 B.n720 VSUBS 0.010488f
C1402 B.n721 VSUBS 0.010488f
C1403 B.n722 VSUBS 0.010488f
C1404 B.n723 VSUBS 0.010488f
C1405 B.n724 VSUBS 0.010488f
C1406 B.n725 VSUBS 0.010488f
C1407 B.n726 VSUBS 0.010488f
C1408 B.n727 VSUBS 0.010488f
C1409 B.n728 VSUBS 0.010488f
C1410 B.n729 VSUBS 0.010488f
C1411 B.n730 VSUBS 0.010488f
C1412 B.n731 VSUBS 0.010488f
C1413 B.n732 VSUBS 0.010488f
C1414 B.n733 VSUBS 0.010488f
C1415 B.n734 VSUBS 0.010488f
C1416 B.n735 VSUBS 0.010488f
C1417 B.n736 VSUBS 0.010488f
C1418 B.n737 VSUBS 0.010488f
C1419 B.n738 VSUBS 0.010488f
C1420 B.n739 VSUBS 0.010488f
C1421 B.n740 VSUBS 0.010488f
C1422 B.n741 VSUBS 0.010488f
C1423 B.n742 VSUBS 0.010488f
C1424 B.n743 VSUBS 0.010488f
C1425 B.n744 VSUBS 0.010488f
C1426 B.n745 VSUBS 0.010488f
C1427 B.n746 VSUBS 0.010488f
C1428 B.n747 VSUBS 0.010488f
C1429 B.n748 VSUBS 0.010488f
C1430 B.n749 VSUBS 0.010488f
C1431 B.n750 VSUBS 0.010488f
C1432 B.n751 VSUBS 0.010488f
C1433 B.n752 VSUBS 0.010488f
C1434 B.n753 VSUBS 0.010488f
C1435 B.n754 VSUBS 0.010488f
C1436 B.n755 VSUBS 0.010488f
C1437 B.n756 VSUBS 0.010488f
C1438 B.n757 VSUBS 0.010488f
C1439 B.n758 VSUBS 0.010488f
C1440 B.n759 VSUBS 0.010488f
C1441 B.n760 VSUBS 0.010488f
C1442 B.n761 VSUBS 0.010488f
C1443 B.n762 VSUBS 0.010488f
C1444 B.n763 VSUBS 0.010488f
C1445 B.n764 VSUBS 0.010488f
C1446 B.n765 VSUBS 0.010488f
C1447 B.n766 VSUBS 0.010488f
C1448 B.n767 VSUBS 0.010488f
C1449 B.n768 VSUBS 0.010488f
C1450 B.n769 VSUBS 0.010488f
C1451 B.n770 VSUBS 0.010488f
C1452 B.n771 VSUBS 0.010488f
C1453 B.n772 VSUBS 0.010488f
C1454 B.n773 VSUBS 0.010488f
C1455 B.n774 VSUBS 0.010488f
C1456 B.n775 VSUBS 0.010488f
C1457 B.n776 VSUBS 0.010488f
C1458 B.n777 VSUBS 0.010488f
C1459 B.n778 VSUBS 0.010488f
C1460 B.n779 VSUBS 0.010488f
C1461 B.n780 VSUBS 0.010488f
C1462 B.n781 VSUBS 0.010488f
C1463 B.n782 VSUBS 0.010488f
C1464 B.n783 VSUBS 0.010488f
C1465 B.n784 VSUBS 0.010488f
C1466 B.n785 VSUBS 0.010488f
C1467 B.n786 VSUBS 0.010488f
C1468 B.n787 VSUBS 0.010488f
C1469 B.n788 VSUBS 0.010488f
C1470 B.n789 VSUBS 0.010488f
C1471 B.n790 VSUBS 0.010488f
C1472 B.n791 VSUBS 0.023749f
.ends

