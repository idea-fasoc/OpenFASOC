* NGSPICE file created from diff_pair_sample_1031.ext - technology: sky130A

.subckt diff_pair_sample_1031 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t1 VP.t0 VTAIL.t2 w_n2030_n1898# sky130_fd_pr__pfet_01v8 ad=1.8135 pd=10.08 as=1.8135 ps=10.08 w=4.65 l=2.32
X1 VDD2.t1 VN.t0 VTAIL.t0 w_n2030_n1898# sky130_fd_pr__pfet_01v8 ad=1.8135 pd=10.08 as=1.8135 ps=10.08 w=4.65 l=2.32
X2 B.t11 B.t9 B.t10 w_n2030_n1898# sky130_fd_pr__pfet_01v8 ad=1.8135 pd=10.08 as=0 ps=0 w=4.65 l=2.32
X3 VDD1.t0 VP.t1 VTAIL.t3 w_n2030_n1898# sky130_fd_pr__pfet_01v8 ad=1.8135 pd=10.08 as=1.8135 ps=10.08 w=4.65 l=2.32
X4 B.t8 B.t6 B.t7 w_n2030_n1898# sky130_fd_pr__pfet_01v8 ad=1.8135 pd=10.08 as=0 ps=0 w=4.65 l=2.32
X5 VDD2.t0 VN.t1 VTAIL.t1 w_n2030_n1898# sky130_fd_pr__pfet_01v8 ad=1.8135 pd=10.08 as=1.8135 ps=10.08 w=4.65 l=2.32
X6 B.t5 B.t3 B.t4 w_n2030_n1898# sky130_fd_pr__pfet_01v8 ad=1.8135 pd=10.08 as=0 ps=0 w=4.65 l=2.32
X7 B.t2 B.t0 B.t1 w_n2030_n1898# sky130_fd_pr__pfet_01v8 ad=1.8135 pd=10.08 as=0 ps=0 w=4.65 l=2.32
R0 VP.n0 VP.t1 135.821
R1 VP.n0 VP.t0 97.4747
R2 VP VP.n0 0.336784
R3 VTAIL.n90 VTAIL.n72 756.745
R4 VTAIL.n18 VTAIL.n0 756.745
R5 VTAIL.n66 VTAIL.n48 756.745
R6 VTAIL.n42 VTAIL.n24 756.745
R7 VTAIL.n81 VTAIL.n80 585
R8 VTAIL.n83 VTAIL.n82 585
R9 VTAIL.n76 VTAIL.n75 585
R10 VTAIL.n89 VTAIL.n88 585
R11 VTAIL.n91 VTAIL.n90 585
R12 VTAIL.n9 VTAIL.n8 585
R13 VTAIL.n11 VTAIL.n10 585
R14 VTAIL.n4 VTAIL.n3 585
R15 VTAIL.n17 VTAIL.n16 585
R16 VTAIL.n19 VTAIL.n18 585
R17 VTAIL.n67 VTAIL.n66 585
R18 VTAIL.n65 VTAIL.n64 585
R19 VTAIL.n52 VTAIL.n51 585
R20 VTAIL.n59 VTAIL.n58 585
R21 VTAIL.n57 VTAIL.n56 585
R22 VTAIL.n43 VTAIL.n42 585
R23 VTAIL.n41 VTAIL.n40 585
R24 VTAIL.n28 VTAIL.n27 585
R25 VTAIL.n35 VTAIL.n34 585
R26 VTAIL.n33 VTAIL.n32 585
R27 VTAIL.n79 VTAIL.t1 328.587
R28 VTAIL.n7 VTAIL.t2 328.587
R29 VTAIL.n55 VTAIL.t3 328.587
R30 VTAIL.n31 VTAIL.t0 328.587
R31 VTAIL.n82 VTAIL.n81 171.744
R32 VTAIL.n82 VTAIL.n75 171.744
R33 VTAIL.n89 VTAIL.n75 171.744
R34 VTAIL.n90 VTAIL.n89 171.744
R35 VTAIL.n10 VTAIL.n9 171.744
R36 VTAIL.n10 VTAIL.n3 171.744
R37 VTAIL.n17 VTAIL.n3 171.744
R38 VTAIL.n18 VTAIL.n17 171.744
R39 VTAIL.n66 VTAIL.n65 171.744
R40 VTAIL.n65 VTAIL.n51 171.744
R41 VTAIL.n58 VTAIL.n51 171.744
R42 VTAIL.n58 VTAIL.n57 171.744
R43 VTAIL.n42 VTAIL.n41 171.744
R44 VTAIL.n41 VTAIL.n27 171.744
R45 VTAIL.n34 VTAIL.n27 171.744
R46 VTAIL.n34 VTAIL.n33 171.744
R47 VTAIL.n81 VTAIL.t1 85.8723
R48 VTAIL.n9 VTAIL.t2 85.8723
R49 VTAIL.n57 VTAIL.t3 85.8723
R50 VTAIL.n33 VTAIL.t0 85.8723
R51 VTAIL.n95 VTAIL.n94 33.9308
R52 VTAIL.n23 VTAIL.n22 33.9308
R53 VTAIL.n71 VTAIL.n70 33.9308
R54 VTAIL.n47 VTAIL.n46 33.9308
R55 VTAIL.n47 VTAIL.n23 20.9445
R56 VTAIL.n95 VTAIL.n71 18.66
R57 VTAIL.n80 VTAIL.n79 16.3651
R58 VTAIL.n8 VTAIL.n7 16.3651
R59 VTAIL.n56 VTAIL.n55 16.3651
R60 VTAIL.n32 VTAIL.n31 16.3651
R61 VTAIL.n83 VTAIL.n78 12.8005
R62 VTAIL.n11 VTAIL.n6 12.8005
R63 VTAIL.n59 VTAIL.n54 12.8005
R64 VTAIL.n35 VTAIL.n30 12.8005
R65 VTAIL.n84 VTAIL.n76 12.0247
R66 VTAIL.n12 VTAIL.n4 12.0247
R67 VTAIL.n60 VTAIL.n52 12.0247
R68 VTAIL.n36 VTAIL.n28 12.0247
R69 VTAIL.n88 VTAIL.n87 11.249
R70 VTAIL.n16 VTAIL.n15 11.249
R71 VTAIL.n64 VTAIL.n63 11.249
R72 VTAIL.n40 VTAIL.n39 11.249
R73 VTAIL.n91 VTAIL.n74 10.4732
R74 VTAIL.n19 VTAIL.n2 10.4732
R75 VTAIL.n67 VTAIL.n50 10.4732
R76 VTAIL.n43 VTAIL.n26 10.4732
R77 VTAIL.n92 VTAIL.n72 9.69747
R78 VTAIL.n20 VTAIL.n0 9.69747
R79 VTAIL.n68 VTAIL.n48 9.69747
R80 VTAIL.n44 VTAIL.n24 9.69747
R81 VTAIL.n94 VTAIL.n93 9.45567
R82 VTAIL.n22 VTAIL.n21 9.45567
R83 VTAIL.n70 VTAIL.n69 9.45567
R84 VTAIL.n46 VTAIL.n45 9.45567
R85 VTAIL.n93 VTAIL.n92 9.3005
R86 VTAIL.n74 VTAIL.n73 9.3005
R87 VTAIL.n87 VTAIL.n86 9.3005
R88 VTAIL.n85 VTAIL.n84 9.3005
R89 VTAIL.n78 VTAIL.n77 9.3005
R90 VTAIL.n21 VTAIL.n20 9.3005
R91 VTAIL.n2 VTAIL.n1 9.3005
R92 VTAIL.n15 VTAIL.n14 9.3005
R93 VTAIL.n13 VTAIL.n12 9.3005
R94 VTAIL.n6 VTAIL.n5 9.3005
R95 VTAIL.n69 VTAIL.n68 9.3005
R96 VTAIL.n50 VTAIL.n49 9.3005
R97 VTAIL.n63 VTAIL.n62 9.3005
R98 VTAIL.n61 VTAIL.n60 9.3005
R99 VTAIL.n54 VTAIL.n53 9.3005
R100 VTAIL.n45 VTAIL.n44 9.3005
R101 VTAIL.n26 VTAIL.n25 9.3005
R102 VTAIL.n39 VTAIL.n38 9.3005
R103 VTAIL.n37 VTAIL.n36 9.3005
R104 VTAIL.n30 VTAIL.n29 9.3005
R105 VTAIL.n94 VTAIL.n72 4.26717
R106 VTAIL.n22 VTAIL.n0 4.26717
R107 VTAIL.n70 VTAIL.n48 4.26717
R108 VTAIL.n46 VTAIL.n24 4.26717
R109 VTAIL.n79 VTAIL.n77 3.73474
R110 VTAIL.n7 VTAIL.n5 3.73474
R111 VTAIL.n55 VTAIL.n53 3.73474
R112 VTAIL.n31 VTAIL.n29 3.73474
R113 VTAIL.n92 VTAIL.n91 3.49141
R114 VTAIL.n20 VTAIL.n19 3.49141
R115 VTAIL.n68 VTAIL.n67 3.49141
R116 VTAIL.n44 VTAIL.n43 3.49141
R117 VTAIL.n88 VTAIL.n74 2.71565
R118 VTAIL.n16 VTAIL.n2 2.71565
R119 VTAIL.n64 VTAIL.n50 2.71565
R120 VTAIL.n40 VTAIL.n26 2.71565
R121 VTAIL.n87 VTAIL.n76 1.93989
R122 VTAIL.n15 VTAIL.n4 1.93989
R123 VTAIL.n63 VTAIL.n52 1.93989
R124 VTAIL.n39 VTAIL.n28 1.93989
R125 VTAIL.n71 VTAIL.n47 1.61257
R126 VTAIL.n84 VTAIL.n83 1.16414
R127 VTAIL.n12 VTAIL.n11 1.16414
R128 VTAIL.n60 VTAIL.n59 1.16414
R129 VTAIL.n36 VTAIL.n35 1.16414
R130 VTAIL VTAIL.n23 1.09964
R131 VTAIL VTAIL.n95 0.513431
R132 VTAIL.n80 VTAIL.n78 0.388379
R133 VTAIL.n8 VTAIL.n6 0.388379
R134 VTAIL.n56 VTAIL.n54 0.388379
R135 VTAIL.n32 VTAIL.n30 0.388379
R136 VTAIL.n85 VTAIL.n77 0.155672
R137 VTAIL.n86 VTAIL.n85 0.155672
R138 VTAIL.n86 VTAIL.n73 0.155672
R139 VTAIL.n93 VTAIL.n73 0.155672
R140 VTAIL.n13 VTAIL.n5 0.155672
R141 VTAIL.n14 VTAIL.n13 0.155672
R142 VTAIL.n14 VTAIL.n1 0.155672
R143 VTAIL.n21 VTAIL.n1 0.155672
R144 VTAIL.n69 VTAIL.n49 0.155672
R145 VTAIL.n62 VTAIL.n49 0.155672
R146 VTAIL.n62 VTAIL.n61 0.155672
R147 VTAIL.n61 VTAIL.n53 0.155672
R148 VTAIL.n45 VTAIL.n25 0.155672
R149 VTAIL.n38 VTAIL.n25 0.155672
R150 VTAIL.n38 VTAIL.n37 0.155672
R151 VTAIL.n37 VTAIL.n29 0.155672
R152 VDD1.n18 VDD1.n0 756.745
R153 VDD1.n41 VDD1.n23 756.745
R154 VDD1.n19 VDD1.n18 585
R155 VDD1.n17 VDD1.n16 585
R156 VDD1.n4 VDD1.n3 585
R157 VDD1.n11 VDD1.n10 585
R158 VDD1.n9 VDD1.n8 585
R159 VDD1.n32 VDD1.n31 585
R160 VDD1.n34 VDD1.n33 585
R161 VDD1.n27 VDD1.n26 585
R162 VDD1.n40 VDD1.n39 585
R163 VDD1.n42 VDD1.n41 585
R164 VDD1.n7 VDD1.t0 328.587
R165 VDD1.n30 VDD1.t1 328.587
R166 VDD1.n18 VDD1.n17 171.744
R167 VDD1.n17 VDD1.n3 171.744
R168 VDD1.n10 VDD1.n3 171.744
R169 VDD1.n10 VDD1.n9 171.744
R170 VDD1.n33 VDD1.n32 171.744
R171 VDD1.n33 VDD1.n26 171.744
R172 VDD1.n40 VDD1.n26 171.744
R173 VDD1.n41 VDD1.n40 171.744
R174 VDD1.n9 VDD1.t0 85.8723
R175 VDD1.n32 VDD1.t1 85.8723
R176 VDD1 VDD1.n45 83.9426
R177 VDD1 VDD1.n22 51.2389
R178 VDD1.n8 VDD1.n7 16.3651
R179 VDD1.n31 VDD1.n30 16.3651
R180 VDD1.n11 VDD1.n6 12.8005
R181 VDD1.n34 VDD1.n29 12.8005
R182 VDD1.n12 VDD1.n4 12.0247
R183 VDD1.n35 VDD1.n27 12.0247
R184 VDD1.n16 VDD1.n15 11.249
R185 VDD1.n39 VDD1.n38 11.249
R186 VDD1.n19 VDD1.n2 10.4732
R187 VDD1.n42 VDD1.n25 10.4732
R188 VDD1.n20 VDD1.n0 9.69747
R189 VDD1.n43 VDD1.n23 9.69747
R190 VDD1.n22 VDD1.n21 9.45567
R191 VDD1.n45 VDD1.n44 9.45567
R192 VDD1.n21 VDD1.n20 9.3005
R193 VDD1.n2 VDD1.n1 9.3005
R194 VDD1.n15 VDD1.n14 9.3005
R195 VDD1.n13 VDD1.n12 9.3005
R196 VDD1.n6 VDD1.n5 9.3005
R197 VDD1.n44 VDD1.n43 9.3005
R198 VDD1.n25 VDD1.n24 9.3005
R199 VDD1.n38 VDD1.n37 9.3005
R200 VDD1.n36 VDD1.n35 9.3005
R201 VDD1.n29 VDD1.n28 9.3005
R202 VDD1.n22 VDD1.n0 4.26717
R203 VDD1.n45 VDD1.n23 4.26717
R204 VDD1.n7 VDD1.n5 3.73474
R205 VDD1.n30 VDD1.n28 3.73474
R206 VDD1.n20 VDD1.n19 3.49141
R207 VDD1.n43 VDD1.n42 3.49141
R208 VDD1.n16 VDD1.n2 2.71565
R209 VDD1.n39 VDD1.n25 2.71565
R210 VDD1.n15 VDD1.n4 1.93989
R211 VDD1.n38 VDD1.n27 1.93989
R212 VDD1.n12 VDD1.n11 1.16414
R213 VDD1.n35 VDD1.n34 1.16414
R214 VDD1.n8 VDD1.n6 0.388379
R215 VDD1.n31 VDD1.n29 0.388379
R216 VDD1.n21 VDD1.n1 0.155672
R217 VDD1.n14 VDD1.n1 0.155672
R218 VDD1.n14 VDD1.n13 0.155672
R219 VDD1.n13 VDD1.n5 0.155672
R220 VDD1.n36 VDD1.n28 0.155672
R221 VDD1.n37 VDD1.n36 0.155672
R222 VDD1.n37 VDD1.n24 0.155672
R223 VDD1.n44 VDD1.n24 0.155672
R224 VN VN.t0 135.917
R225 VN VN.t1 97.811
R226 VDD2.n41 VDD2.n23 756.745
R227 VDD2.n18 VDD2.n0 756.745
R228 VDD2.n42 VDD2.n41 585
R229 VDD2.n40 VDD2.n39 585
R230 VDD2.n27 VDD2.n26 585
R231 VDD2.n34 VDD2.n33 585
R232 VDD2.n32 VDD2.n31 585
R233 VDD2.n9 VDD2.n8 585
R234 VDD2.n11 VDD2.n10 585
R235 VDD2.n4 VDD2.n3 585
R236 VDD2.n17 VDD2.n16 585
R237 VDD2.n19 VDD2.n18 585
R238 VDD2.n30 VDD2.t1 328.587
R239 VDD2.n7 VDD2.t0 328.587
R240 VDD2.n41 VDD2.n40 171.744
R241 VDD2.n40 VDD2.n26 171.744
R242 VDD2.n33 VDD2.n26 171.744
R243 VDD2.n33 VDD2.n32 171.744
R244 VDD2.n10 VDD2.n9 171.744
R245 VDD2.n10 VDD2.n3 171.744
R246 VDD2.n17 VDD2.n3 171.744
R247 VDD2.n18 VDD2.n17 171.744
R248 VDD2.n32 VDD2.t1 85.8723
R249 VDD2.n9 VDD2.t0 85.8723
R250 VDD2.n46 VDD2.n22 82.8466
R251 VDD2.n46 VDD2.n45 50.6096
R252 VDD2.n31 VDD2.n30 16.3651
R253 VDD2.n8 VDD2.n7 16.3651
R254 VDD2.n34 VDD2.n29 12.8005
R255 VDD2.n11 VDD2.n6 12.8005
R256 VDD2.n35 VDD2.n27 12.0247
R257 VDD2.n12 VDD2.n4 12.0247
R258 VDD2.n39 VDD2.n38 11.249
R259 VDD2.n16 VDD2.n15 11.249
R260 VDD2.n42 VDD2.n25 10.4732
R261 VDD2.n19 VDD2.n2 10.4732
R262 VDD2.n43 VDD2.n23 9.69747
R263 VDD2.n20 VDD2.n0 9.69747
R264 VDD2.n45 VDD2.n44 9.45567
R265 VDD2.n22 VDD2.n21 9.45567
R266 VDD2.n44 VDD2.n43 9.3005
R267 VDD2.n25 VDD2.n24 9.3005
R268 VDD2.n38 VDD2.n37 9.3005
R269 VDD2.n36 VDD2.n35 9.3005
R270 VDD2.n29 VDD2.n28 9.3005
R271 VDD2.n21 VDD2.n20 9.3005
R272 VDD2.n2 VDD2.n1 9.3005
R273 VDD2.n15 VDD2.n14 9.3005
R274 VDD2.n13 VDD2.n12 9.3005
R275 VDD2.n6 VDD2.n5 9.3005
R276 VDD2.n45 VDD2.n23 4.26717
R277 VDD2.n22 VDD2.n0 4.26717
R278 VDD2.n30 VDD2.n28 3.73474
R279 VDD2.n7 VDD2.n5 3.73474
R280 VDD2.n43 VDD2.n42 3.49141
R281 VDD2.n20 VDD2.n19 3.49141
R282 VDD2.n39 VDD2.n25 2.71565
R283 VDD2.n16 VDD2.n2 2.71565
R284 VDD2.n38 VDD2.n27 1.93989
R285 VDD2.n15 VDD2.n4 1.93989
R286 VDD2.n35 VDD2.n34 1.16414
R287 VDD2.n12 VDD2.n11 1.16414
R288 VDD2 VDD2.n46 0.62981
R289 VDD2.n31 VDD2.n29 0.388379
R290 VDD2.n8 VDD2.n6 0.388379
R291 VDD2.n44 VDD2.n24 0.155672
R292 VDD2.n37 VDD2.n24 0.155672
R293 VDD2.n37 VDD2.n36 0.155672
R294 VDD2.n36 VDD2.n28 0.155672
R295 VDD2.n13 VDD2.n5 0.155672
R296 VDD2.n14 VDD2.n13 0.155672
R297 VDD2.n14 VDD2.n1 0.155672
R298 VDD2.n21 VDD2.n1 0.155672
R299 B.n217 B.n216 585
R300 B.n215 B.n68 585
R301 B.n214 B.n213 585
R302 B.n212 B.n69 585
R303 B.n211 B.n210 585
R304 B.n209 B.n70 585
R305 B.n208 B.n207 585
R306 B.n206 B.n71 585
R307 B.n205 B.n204 585
R308 B.n203 B.n72 585
R309 B.n202 B.n201 585
R310 B.n200 B.n73 585
R311 B.n199 B.n198 585
R312 B.n197 B.n74 585
R313 B.n196 B.n195 585
R314 B.n194 B.n75 585
R315 B.n193 B.n192 585
R316 B.n191 B.n76 585
R317 B.n190 B.n189 585
R318 B.n188 B.n77 585
R319 B.n187 B.n186 585
R320 B.n182 B.n78 585
R321 B.n181 B.n180 585
R322 B.n179 B.n79 585
R323 B.n178 B.n177 585
R324 B.n176 B.n80 585
R325 B.n175 B.n174 585
R326 B.n173 B.n81 585
R327 B.n172 B.n171 585
R328 B.n170 B.n82 585
R329 B.n168 B.n167 585
R330 B.n166 B.n85 585
R331 B.n165 B.n164 585
R332 B.n163 B.n86 585
R333 B.n162 B.n161 585
R334 B.n160 B.n87 585
R335 B.n159 B.n158 585
R336 B.n157 B.n88 585
R337 B.n156 B.n155 585
R338 B.n154 B.n89 585
R339 B.n153 B.n152 585
R340 B.n151 B.n90 585
R341 B.n150 B.n149 585
R342 B.n148 B.n91 585
R343 B.n147 B.n146 585
R344 B.n145 B.n92 585
R345 B.n144 B.n143 585
R346 B.n142 B.n93 585
R347 B.n141 B.n140 585
R348 B.n139 B.n94 585
R349 B.n218 B.n67 585
R350 B.n220 B.n219 585
R351 B.n221 B.n66 585
R352 B.n223 B.n222 585
R353 B.n224 B.n65 585
R354 B.n226 B.n225 585
R355 B.n227 B.n64 585
R356 B.n229 B.n228 585
R357 B.n230 B.n63 585
R358 B.n232 B.n231 585
R359 B.n233 B.n62 585
R360 B.n235 B.n234 585
R361 B.n236 B.n61 585
R362 B.n238 B.n237 585
R363 B.n239 B.n60 585
R364 B.n241 B.n240 585
R365 B.n242 B.n59 585
R366 B.n244 B.n243 585
R367 B.n245 B.n58 585
R368 B.n247 B.n246 585
R369 B.n248 B.n57 585
R370 B.n250 B.n249 585
R371 B.n251 B.n56 585
R372 B.n253 B.n252 585
R373 B.n254 B.n55 585
R374 B.n256 B.n255 585
R375 B.n257 B.n54 585
R376 B.n259 B.n258 585
R377 B.n260 B.n53 585
R378 B.n262 B.n261 585
R379 B.n263 B.n52 585
R380 B.n265 B.n264 585
R381 B.n266 B.n51 585
R382 B.n268 B.n267 585
R383 B.n269 B.n50 585
R384 B.n271 B.n270 585
R385 B.n272 B.n49 585
R386 B.n274 B.n273 585
R387 B.n275 B.n48 585
R388 B.n277 B.n276 585
R389 B.n278 B.n47 585
R390 B.n280 B.n279 585
R391 B.n281 B.n46 585
R392 B.n283 B.n282 585
R393 B.n284 B.n45 585
R394 B.n286 B.n285 585
R395 B.n287 B.n44 585
R396 B.n289 B.n288 585
R397 B.n365 B.n364 585
R398 B.n363 B.n14 585
R399 B.n362 B.n361 585
R400 B.n360 B.n15 585
R401 B.n359 B.n358 585
R402 B.n357 B.n16 585
R403 B.n356 B.n355 585
R404 B.n354 B.n17 585
R405 B.n353 B.n352 585
R406 B.n351 B.n18 585
R407 B.n350 B.n349 585
R408 B.n348 B.n19 585
R409 B.n347 B.n346 585
R410 B.n345 B.n20 585
R411 B.n344 B.n343 585
R412 B.n342 B.n21 585
R413 B.n341 B.n340 585
R414 B.n339 B.n22 585
R415 B.n338 B.n337 585
R416 B.n336 B.n23 585
R417 B.n334 B.n333 585
R418 B.n332 B.n26 585
R419 B.n331 B.n330 585
R420 B.n329 B.n27 585
R421 B.n328 B.n327 585
R422 B.n326 B.n28 585
R423 B.n325 B.n324 585
R424 B.n323 B.n29 585
R425 B.n322 B.n321 585
R426 B.n320 B.n30 585
R427 B.n319 B.n318 585
R428 B.n317 B.n31 585
R429 B.n316 B.n315 585
R430 B.n314 B.n35 585
R431 B.n313 B.n312 585
R432 B.n311 B.n36 585
R433 B.n310 B.n309 585
R434 B.n308 B.n37 585
R435 B.n307 B.n306 585
R436 B.n305 B.n38 585
R437 B.n304 B.n303 585
R438 B.n302 B.n39 585
R439 B.n301 B.n300 585
R440 B.n299 B.n40 585
R441 B.n298 B.n297 585
R442 B.n296 B.n41 585
R443 B.n295 B.n294 585
R444 B.n293 B.n42 585
R445 B.n292 B.n291 585
R446 B.n290 B.n43 585
R447 B.n366 B.n13 585
R448 B.n368 B.n367 585
R449 B.n369 B.n12 585
R450 B.n371 B.n370 585
R451 B.n372 B.n11 585
R452 B.n374 B.n373 585
R453 B.n375 B.n10 585
R454 B.n377 B.n376 585
R455 B.n378 B.n9 585
R456 B.n380 B.n379 585
R457 B.n381 B.n8 585
R458 B.n383 B.n382 585
R459 B.n384 B.n7 585
R460 B.n386 B.n385 585
R461 B.n387 B.n6 585
R462 B.n389 B.n388 585
R463 B.n390 B.n5 585
R464 B.n392 B.n391 585
R465 B.n393 B.n4 585
R466 B.n395 B.n394 585
R467 B.n396 B.n3 585
R468 B.n398 B.n397 585
R469 B.n399 B.n0 585
R470 B.n2 B.n1 585
R471 B.n106 B.n105 585
R472 B.n108 B.n107 585
R473 B.n109 B.n104 585
R474 B.n111 B.n110 585
R475 B.n112 B.n103 585
R476 B.n114 B.n113 585
R477 B.n115 B.n102 585
R478 B.n117 B.n116 585
R479 B.n118 B.n101 585
R480 B.n120 B.n119 585
R481 B.n121 B.n100 585
R482 B.n123 B.n122 585
R483 B.n124 B.n99 585
R484 B.n126 B.n125 585
R485 B.n127 B.n98 585
R486 B.n129 B.n128 585
R487 B.n130 B.n97 585
R488 B.n132 B.n131 585
R489 B.n133 B.n96 585
R490 B.n135 B.n134 585
R491 B.n136 B.n95 585
R492 B.n138 B.n137 585
R493 B.n137 B.n94 497.305
R494 B.n218 B.n217 497.305
R495 B.n290 B.n289 497.305
R496 B.n364 B.n13 497.305
R497 B.n183 B.t10 296.709
R498 B.n32 B.t2 296.709
R499 B.n83 B.t4 296.709
R500 B.n24 B.t8 296.709
R501 B.n401 B.n400 256.663
R502 B.n83 B.t3 255.886
R503 B.n183 B.t9 255.886
R504 B.n32 B.t0 255.886
R505 B.n24 B.t6 255.886
R506 B.n184 B.t11 245.315
R507 B.n33 B.t1 245.315
R508 B.n84 B.t5 245.315
R509 B.n25 B.t7 245.315
R510 B.n400 B.n399 235.042
R511 B.n400 B.n2 235.042
R512 B.n141 B.n94 163.367
R513 B.n142 B.n141 163.367
R514 B.n143 B.n142 163.367
R515 B.n143 B.n92 163.367
R516 B.n147 B.n92 163.367
R517 B.n148 B.n147 163.367
R518 B.n149 B.n148 163.367
R519 B.n149 B.n90 163.367
R520 B.n153 B.n90 163.367
R521 B.n154 B.n153 163.367
R522 B.n155 B.n154 163.367
R523 B.n155 B.n88 163.367
R524 B.n159 B.n88 163.367
R525 B.n160 B.n159 163.367
R526 B.n161 B.n160 163.367
R527 B.n161 B.n86 163.367
R528 B.n165 B.n86 163.367
R529 B.n166 B.n165 163.367
R530 B.n167 B.n166 163.367
R531 B.n167 B.n82 163.367
R532 B.n172 B.n82 163.367
R533 B.n173 B.n172 163.367
R534 B.n174 B.n173 163.367
R535 B.n174 B.n80 163.367
R536 B.n178 B.n80 163.367
R537 B.n179 B.n178 163.367
R538 B.n180 B.n179 163.367
R539 B.n180 B.n78 163.367
R540 B.n187 B.n78 163.367
R541 B.n188 B.n187 163.367
R542 B.n189 B.n188 163.367
R543 B.n189 B.n76 163.367
R544 B.n193 B.n76 163.367
R545 B.n194 B.n193 163.367
R546 B.n195 B.n194 163.367
R547 B.n195 B.n74 163.367
R548 B.n199 B.n74 163.367
R549 B.n200 B.n199 163.367
R550 B.n201 B.n200 163.367
R551 B.n201 B.n72 163.367
R552 B.n205 B.n72 163.367
R553 B.n206 B.n205 163.367
R554 B.n207 B.n206 163.367
R555 B.n207 B.n70 163.367
R556 B.n211 B.n70 163.367
R557 B.n212 B.n211 163.367
R558 B.n213 B.n212 163.367
R559 B.n213 B.n68 163.367
R560 B.n217 B.n68 163.367
R561 B.n289 B.n44 163.367
R562 B.n285 B.n44 163.367
R563 B.n285 B.n284 163.367
R564 B.n284 B.n283 163.367
R565 B.n283 B.n46 163.367
R566 B.n279 B.n46 163.367
R567 B.n279 B.n278 163.367
R568 B.n278 B.n277 163.367
R569 B.n277 B.n48 163.367
R570 B.n273 B.n48 163.367
R571 B.n273 B.n272 163.367
R572 B.n272 B.n271 163.367
R573 B.n271 B.n50 163.367
R574 B.n267 B.n50 163.367
R575 B.n267 B.n266 163.367
R576 B.n266 B.n265 163.367
R577 B.n265 B.n52 163.367
R578 B.n261 B.n52 163.367
R579 B.n261 B.n260 163.367
R580 B.n260 B.n259 163.367
R581 B.n259 B.n54 163.367
R582 B.n255 B.n54 163.367
R583 B.n255 B.n254 163.367
R584 B.n254 B.n253 163.367
R585 B.n253 B.n56 163.367
R586 B.n249 B.n56 163.367
R587 B.n249 B.n248 163.367
R588 B.n248 B.n247 163.367
R589 B.n247 B.n58 163.367
R590 B.n243 B.n58 163.367
R591 B.n243 B.n242 163.367
R592 B.n242 B.n241 163.367
R593 B.n241 B.n60 163.367
R594 B.n237 B.n60 163.367
R595 B.n237 B.n236 163.367
R596 B.n236 B.n235 163.367
R597 B.n235 B.n62 163.367
R598 B.n231 B.n62 163.367
R599 B.n231 B.n230 163.367
R600 B.n230 B.n229 163.367
R601 B.n229 B.n64 163.367
R602 B.n225 B.n64 163.367
R603 B.n225 B.n224 163.367
R604 B.n224 B.n223 163.367
R605 B.n223 B.n66 163.367
R606 B.n219 B.n66 163.367
R607 B.n219 B.n218 163.367
R608 B.n364 B.n363 163.367
R609 B.n363 B.n362 163.367
R610 B.n362 B.n15 163.367
R611 B.n358 B.n15 163.367
R612 B.n358 B.n357 163.367
R613 B.n357 B.n356 163.367
R614 B.n356 B.n17 163.367
R615 B.n352 B.n17 163.367
R616 B.n352 B.n351 163.367
R617 B.n351 B.n350 163.367
R618 B.n350 B.n19 163.367
R619 B.n346 B.n19 163.367
R620 B.n346 B.n345 163.367
R621 B.n345 B.n344 163.367
R622 B.n344 B.n21 163.367
R623 B.n340 B.n21 163.367
R624 B.n340 B.n339 163.367
R625 B.n339 B.n338 163.367
R626 B.n338 B.n23 163.367
R627 B.n333 B.n23 163.367
R628 B.n333 B.n332 163.367
R629 B.n332 B.n331 163.367
R630 B.n331 B.n27 163.367
R631 B.n327 B.n27 163.367
R632 B.n327 B.n326 163.367
R633 B.n326 B.n325 163.367
R634 B.n325 B.n29 163.367
R635 B.n321 B.n29 163.367
R636 B.n321 B.n320 163.367
R637 B.n320 B.n319 163.367
R638 B.n319 B.n31 163.367
R639 B.n315 B.n31 163.367
R640 B.n315 B.n314 163.367
R641 B.n314 B.n313 163.367
R642 B.n313 B.n36 163.367
R643 B.n309 B.n36 163.367
R644 B.n309 B.n308 163.367
R645 B.n308 B.n307 163.367
R646 B.n307 B.n38 163.367
R647 B.n303 B.n38 163.367
R648 B.n303 B.n302 163.367
R649 B.n302 B.n301 163.367
R650 B.n301 B.n40 163.367
R651 B.n297 B.n40 163.367
R652 B.n297 B.n296 163.367
R653 B.n296 B.n295 163.367
R654 B.n295 B.n42 163.367
R655 B.n291 B.n42 163.367
R656 B.n291 B.n290 163.367
R657 B.n368 B.n13 163.367
R658 B.n369 B.n368 163.367
R659 B.n370 B.n369 163.367
R660 B.n370 B.n11 163.367
R661 B.n374 B.n11 163.367
R662 B.n375 B.n374 163.367
R663 B.n376 B.n375 163.367
R664 B.n376 B.n9 163.367
R665 B.n380 B.n9 163.367
R666 B.n381 B.n380 163.367
R667 B.n382 B.n381 163.367
R668 B.n382 B.n7 163.367
R669 B.n386 B.n7 163.367
R670 B.n387 B.n386 163.367
R671 B.n388 B.n387 163.367
R672 B.n388 B.n5 163.367
R673 B.n392 B.n5 163.367
R674 B.n393 B.n392 163.367
R675 B.n394 B.n393 163.367
R676 B.n394 B.n3 163.367
R677 B.n398 B.n3 163.367
R678 B.n399 B.n398 163.367
R679 B.n106 B.n2 163.367
R680 B.n107 B.n106 163.367
R681 B.n107 B.n104 163.367
R682 B.n111 B.n104 163.367
R683 B.n112 B.n111 163.367
R684 B.n113 B.n112 163.367
R685 B.n113 B.n102 163.367
R686 B.n117 B.n102 163.367
R687 B.n118 B.n117 163.367
R688 B.n119 B.n118 163.367
R689 B.n119 B.n100 163.367
R690 B.n123 B.n100 163.367
R691 B.n124 B.n123 163.367
R692 B.n125 B.n124 163.367
R693 B.n125 B.n98 163.367
R694 B.n129 B.n98 163.367
R695 B.n130 B.n129 163.367
R696 B.n131 B.n130 163.367
R697 B.n131 B.n96 163.367
R698 B.n135 B.n96 163.367
R699 B.n136 B.n135 163.367
R700 B.n137 B.n136 163.367
R701 B.n169 B.n84 59.5399
R702 B.n185 B.n184 59.5399
R703 B.n34 B.n33 59.5399
R704 B.n335 B.n25 59.5399
R705 B.n84 B.n83 51.3944
R706 B.n184 B.n183 51.3944
R707 B.n33 B.n32 51.3944
R708 B.n25 B.n24 51.3944
R709 B.n366 B.n365 32.3127
R710 B.n288 B.n43 32.3127
R711 B.n216 B.n67 32.3127
R712 B.n139 B.n138 32.3127
R713 B B.n401 18.0485
R714 B.n367 B.n366 10.6151
R715 B.n367 B.n12 10.6151
R716 B.n371 B.n12 10.6151
R717 B.n372 B.n371 10.6151
R718 B.n373 B.n372 10.6151
R719 B.n373 B.n10 10.6151
R720 B.n377 B.n10 10.6151
R721 B.n378 B.n377 10.6151
R722 B.n379 B.n378 10.6151
R723 B.n379 B.n8 10.6151
R724 B.n383 B.n8 10.6151
R725 B.n384 B.n383 10.6151
R726 B.n385 B.n384 10.6151
R727 B.n385 B.n6 10.6151
R728 B.n389 B.n6 10.6151
R729 B.n390 B.n389 10.6151
R730 B.n391 B.n390 10.6151
R731 B.n391 B.n4 10.6151
R732 B.n395 B.n4 10.6151
R733 B.n396 B.n395 10.6151
R734 B.n397 B.n396 10.6151
R735 B.n397 B.n0 10.6151
R736 B.n365 B.n14 10.6151
R737 B.n361 B.n14 10.6151
R738 B.n361 B.n360 10.6151
R739 B.n360 B.n359 10.6151
R740 B.n359 B.n16 10.6151
R741 B.n355 B.n16 10.6151
R742 B.n355 B.n354 10.6151
R743 B.n354 B.n353 10.6151
R744 B.n353 B.n18 10.6151
R745 B.n349 B.n18 10.6151
R746 B.n349 B.n348 10.6151
R747 B.n348 B.n347 10.6151
R748 B.n347 B.n20 10.6151
R749 B.n343 B.n20 10.6151
R750 B.n343 B.n342 10.6151
R751 B.n342 B.n341 10.6151
R752 B.n341 B.n22 10.6151
R753 B.n337 B.n22 10.6151
R754 B.n337 B.n336 10.6151
R755 B.n334 B.n26 10.6151
R756 B.n330 B.n26 10.6151
R757 B.n330 B.n329 10.6151
R758 B.n329 B.n328 10.6151
R759 B.n328 B.n28 10.6151
R760 B.n324 B.n28 10.6151
R761 B.n324 B.n323 10.6151
R762 B.n323 B.n322 10.6151
R763 B.n322 B.n30 10.6151
R764 B.n318 B.n317 10.6151
R765 B.n317 B.n316 10.6151
R766 B.n316 B.n35 10.6151
R767 B.n312 B.n35 10.6151
R768 B.n312 B.n311 10.6151
R769 B.n311 B.n310 10.6151
R770 B.n310 B.n37 10.6151
R771 B.n306 B.n37 10.6151
R772 B.n306 B.n305 10.6151
R773 B.n305 B.n304 10.6151
R774 B.n304 B.n39 10.6151
R775 B.n300 B.n39 10.6151
R776 B.n300 B.n299 10.6151
R777 B.n299 B.n298 10.6151
R778 B.n298 B.n41 10.6151
R779 B.n294 B.n41 10.6151
R780 B.n294 B.n293 10.6151
R781 B.n293 B.n292 10.6151
R782 B.n292 B.n43 10.6151
R783 B.n288 B.n287 10.6151
R784 B.n287 B.n286 10.6151
R785 B.n286 B.n45 10.6151
R786 B.n282 B.n45 10.6151
R787 B.n282 B.n281 10.6151
R788 B.n281 B.n280 10.6151
R789 B.n280 B.n47 10.6151
R790 B.n276 B.n47 10.6151
R791 B.n276 B.n275 10.6151
R792 B.n275 B.n274 10.6151
R793 B.n274 B.n49 10.6151
R794 B.n270 B.n49 10.6151
R795 B.n270 B.n269 10.6151
R796 B.n269 B.n268 10.6151
R797 B.n268 B.n51 10.6151
R798 B.n264 B.n51 10.6151
R799 B.n264 B.n263 10.6151
R800 B.n263 B.n262 10.6151
R801 B.n262 B.n53 10.6151
R802 B.n258 B.n53 10.6151
R803 B.n258 B.n257 10.6151
R804 B.n257 B.n256 10.6151
R805 B.n256 B.n55 10.6151
R806 B.n252 B.n55 10.6151
R807 B.n252 B.n251 10.6151
R808 B.n251 B.n250 10.6151
R809 B.n250 B.n57 10.6151
R810 B.n246 B.n57 10.6151
R811 B.n246 B.n245 10.6151
R812 B.n245 B.n244 10.6151
R813 B.n244 B.n59 10.6151
R814 B.n240 B.n59 10.6151
R815 B.n240 B.n239 10.6151
R816 B.n239 B.n238 10.6151
R817 B.n238 B.n61 10.6151
R818 B.n234 B.n61 10.6151
R819 B.n234 B.n233 10.6151
R820 B.n233 B.n232 10.6151
R821 B.n232 B.n63 10.6151
R822 B.n228 B.n63 10.6151
R823 B.n228 B.n227 10.6151
R824 B.n227 B.n226 10.6151
R825 B.n226 B.n65 10.6151
R826 B.n222 B.n65 10.6151
R827 B.n222 B.n221 10.6151
R828 B.n221 B.n220 10.6151
R829 B.n220 B.n67 10.6151
R830 B.n105 B.n1 10.6151
R831 B.n108 B.n105 10.6151
R832 B.n109 B.n108 10.6151
R833 B.n110 B.n109 10.6151
R834 B.n110 B.n103 10.6151
R835 B.n114 B.n103 10.6151
R836 B.n115 B.n114 10.6151
R837 B.n116 B.n115 10.6151
R838 B.n116 B.n101 10.6151
R839 B.n120 B.n101 10.6151
R840 B.n121 B.n120 10.6151
R841 B.n122 B.n121 10.6151
R842 B.n122 B.n99 10.6151
R843 B.n126 B.n99 10.6151
R844 B.n127 B.n126 10.6151
R845 B.n128 B.n127 10.6151
R846 B.n128 B.n97 10.6151
R847 B.n132 B.n97 10.6151
R848 B.n133 B.n132 10.6151
R849 B.n134 B.n133 10.6151
R850 B.n134 B.n95 10.6151
R851 B.n138 B.n95 10.6151
R852 B.n140 B.n139 10.6151
R853 B.n140 B.n93 10.6151
R854 B.n144 B.n93 10.6151
R855 B.n145 B.n144 10.6151
R856 B.n146 B.n145 10.6151
R857 B.n146 B.n91 10.6151
R858 B.n150 B.n91 10.6151
R859 B.n151 B.n150 10.6151
R860 B.n152 B.n151 10.6151
R861 B.n152 B.n89 10.6151
R862 B.n156 B.n89 10.6151
R863 B.n157 B.n156 10.6151
R864 B.n158 B.n157 10.6151
R865 B.n158 B.n87 10.6151
R866 B.n162 B.n87 10.6151
R867 B.n163 B.n162 10.6151
R868 B.n164 B.n163 10.6151
R869 B.n164 B.n85 10.6151
R870 B.n168 B.n85 10.6151
R871 B.n171 B.n170 10.6151
R872 B.n171 B.n81 10.6151
R873 B.n175 B.n81 10.6151
R874 B.n176 B.n175 10.6151
R875 B.n177 B.n176 10.6151
R876 B.n177 B.n79 10.6151
R877 B.n181 B.n79 10.6151
R878 B.n182 B.n181 10.6151
R879 B.n186 B.n182 10.6151
R880 B.n190 B.n77 10.6151
R881 B.n191 B.n190 10.6151
R882 B.n192 B.n191 10.6151
R883 B.n192 B.n75 10.6151
R884 B.n196 B.n75 10.6151
R885 B.n197 B.n196 10.6151
R886 B.n198 B.n197 10.6151
R887 B.n198 B.n73 10.6151
R888 B.n202 B.n73 10.6151
R889 B.n203 B.n202 10.6151
R890 B.n204 B.n203 10.6151
R891 B.n204 B.n71 10.6151
R892 B.n208 B.n71 10.6151
R893 B.n209 B.n208 10.6151
R894 B.n210 B.n209 10.6151
R895 B.n210 B.n69 10.6151
R896 B.n214 B.n69 10.6151
R897 B.n215 B.n214 10.6151
R898 B.n216 B.n215 10.6151
R899 B.n336 B.n335 9.36635
R900 B.n318 B.n34 9.36635
R901 B.n169 B.n168 9.36635
R902 B.n185 B.n77 9.36635
R903 B.n401 B.n0 8.11757
R904 B.n401 B.n1 8.11757
R905 B.n335 B.n334 1.24928
R906 B.n34 B.n30 1.24928
R907 B.n170 B.n169 1.24928
R908 B.n186 B.n185 1.24928
C0 VTAIL VN 1.2775f
C1 w_n2030_n1898# VDD1 1.23519f
C2 VP B 1.33694f
C3 w_n2030_n1898# VTAIL 1.70153f
C4 VP VN 3.96417f
C5 VP w_n2030_n1898# 2.90095f
C6 VTAIL VDD1 3.05113f
C7 B VDD2 1.11913f
C8 VDD2 VN 1.21295f
C9 VP VDD1 1.38432f
C10 VP VTAIL 1.29169f
C11 w_n2030_n1898# VDD2 1.25741f
C12 B VN 0.91402f
C13 w_n2030_n1898# B 6.45704f
C14 VDD2 VDD1 0.640184f
C15 w_n2030_n1898# VN 2.64307f
C16 VDD2 VTAIL 3.10144f
C17 VP VDD2 0.324909f
C18 B VDD1 1.09142f
C19 VDD1 VN 0.151904f
C20 B VTAIL 1.9049f
C21 VDD2 VSUBS 0.595609f
C22 VDD1 VSUBS 2.204989f
C23 VTAIL VSUBS 0.447732f
C24 VN VSUBS 5.17252f
C25 VP VSUBS 1.222185f
C26 B VSUBS 2.9275f
C27 w_n2030_n1898# VSUBS 48.3546f
C28 B.n0 VSUBS 0.005939f
C29 B.n1 VSUBS 0.005939f
C30 B.n2 VSUBS 0.008783f
C31 B.n3 VSUBS 0.006731f
C32 B.n4 VSUBS 0.006731f
C33 B.n5 VSUBS 0.006731f
C34 B.n6 VSUBS 0.006731f
C35 B.n7 VSUBS 0.006731f
C36 B.n8 VSUBS 0.006731f
C37 B.n9 VSUBS 0.006731f
C38 B.n10 VSUBS 0.006731f
C39 B.n11 VSUBS 0.006731f
C40 B.n12 VSUBS 0.006731f
C41 B.n13 VSUBS 0.014982f
C42 B.n14 VSUBS 0.006731f
C43 B.n15 VSUBS 0.006731f
C44 B.n16 VSUBS 0.006731f
C45 B.n17 VSUBS 0.006731f
C46 B.n18 VSUBS 0.006731f
C47 B.n19 VSUBS 0.006731f
C48 B.n20 VSUBS 0.006731f
C49 B.n21 VSUBS 0.006731f
C50 B.n22 VSUBS 0.006731f
C51 B.n23 VSUBS 0.006731f
C52 B.t7 VSUBS 0.064843f
C53 B.t8 VSUBS 0.084586f
C54 B.t6 VSUBS 0.49373f
C55 B.n24 VSUBS 0.147765f
C56 B.n25 VSUBS 0.12358f
C57 B.n26 VSUBS 0.006731f
C58 B.n27 VSUBS 0.006731f
C59 B.n28 VSUBS 0.006731f
C60 B.n29 VSUBS 0.006731f
C61 B.n30 VSUBS 0.003761f
C62 B.n31 VSUBS 0.006731f
C63 B.t1 VSUBS 0.064844f
C64 B.t2 VSUBS 0.084587f
C65 B.t0 VSUBS 0.49373f
C66 B.n32 VSUBS 0.147764f
C67 B.n33 VSUBS 0.123579f
C68 B.n34 VSUBS 0.015595f
C69 B.n35 VSUBS 0.006731f
C70 B.n36 VSUBS 0.006731f
C71 B.n37 VSUBS 0.006731f
C72 B.n38 VSUBS 0.006731f
C73 B.n39 VSUBS 0.006731f
C74 B.n40 VSUBS 0.006731f
C75 B.n41 VSUBS 0.006731f
C76 B.n42 VSUBS 0.006731f
C77 B.n43 VSUBS 0.016296f
C78 B.n44 VSUBS 0.006731f
C79 B.n45 VSUBS 0.006731f
C80 B.n46 VSUBS 0.006731f
C81 B.n47 VSUBS 0.006731f
C82 B.n48 VSUBS 0.006731f
C83 B.n49 VSUBS 0.006731f
C84 B.n50 VSUBS 0.006731f
C85 B.n51 VSUBS 0.006731f
C86 B.n52 VSUBS 0.006731f
C87 B.n53 VSUBS 0.006731f
C88 B.n54 VSUBS 0.006731f
C89 B.n55 VSUBS 0.006731f
C90 B.n56 VSUBS 0.006731f
C91 B.n57 VSUBS 0.006731f
C92 B.n58 VSUBS 0.006731f
C93 B.n59 VSUBS 0.006731f
C94 B.n60 VSUBS 0.006731f
C95 B.n61 VSUBS 0.006731f
C96 B.n62 VSUBS 0.006731f
C97 B.n63 VSUBS 0.006731f
C98 B.n64 VSUBS 0.006731f
C99 B.n65 VSUBS 0.006731f
C100 B.n66 VSUBS 0.006731f
C101 B.n67 VSUBS 0.015786f
C102 B.n68 VSUBS 0.006731f
C103 B.n69 VSUBS 0.006731f
C104 B.n70 VSUBS 0.006731f
C105 B.n71 VSUBS 0.006731f
C106 B.n72 VSUBS 0.006731f
C107 B.n73 VSUBS 0.006731f
C108 B.n74 VSUBS 0.006731f
C109 B.n75 VSUBS 0.006731f
C110 B.n76 VSUBS 0.006731f
C111 B.n77 VSUBS 0.006335f
C112 B.n78 VSUBS 0.006731f
C113 B.n79 VSUBS 0.006731f
C114 B.n80 VSUBS 0.006731f
C115 B.n81 VSUBS 0.006731f
C116 B.n82 VSUBS 0.006731f
C117 B.t5 VSUBS 0.064843f
C118 B.t4 VSUBS 0.084586f
C119 B.t3 VSUBS 0.49373f
C120 B.n83 VSUBS 0.147765f
C121 B.n84 VSUBS 0.12358f
C122 B.n85 VSUBS 0.006731f
C123 B.n86 VSUBS 0.006731f
C124 B.n87 VSUBS 0.006731f
C125 B.n88 VSUBS 0.006731f
C126 B.n89 VSUBS 0.006731f
C127 B.n90 VSUBS 0.006731f
C128 B.n91 VSUBS 0.006731f
C129 B.n92 VSUBS 0.006731f
C130 B.n93 VSUBS 0.006731f
C131 B.n94 VSUBS 0.016296f
C132 B.n95 VSUBS 0.006731f
C133 B.n96 VSUBS 0.006731f
C134 B.n97 VSUBS 0.006731f
C135 B.n98 VSUBS 0.006731f
C136 B.n99 VSUBS 0.006731f
C137 B.n100 VSUBS 0.006731f
C138 B.n101 VSUBS 0.006731f
C139 B.n102 VSUBS 0.006731f
C140 B.n103 VSUBS 0.006731f
C141 B.n104 VSUBS 0.006731f
C142 B.n105 VSUBS 0.006731f
C143 B.n106 VSUBS 0.006731f
C144 B.n107 VSUBS 0.006731f
C145 B.n108 VSUBS 0.006731f
C146 B.n109 VSUBS 0.006731f
C147 B.n110 VSUBS 0.006731f
C148 B.n111 VSUBS 0.006731f
C149 B.n112 VSUBS 0.006731f
C150 B.n113 VSUBS 0.006731f
C151 B.n114 VSUBS 0.006731f
C152 B.n115 VSUBS 0.006731f
C153 B.n116 VSUBS 0.006731f
C154 B.n117 VSUBS 0.006731f
C155 B.n118 VSUBS 0.006731f
C156 B.n119 VSUBS 0.006731f
C157 B.n120 VSUBS 0.006731f
C158 B.n121 VSUBS 0.006731f
C159 B.n122 VSUBS 0.006731f
C160 B.n123 VSUBS 0.006731f
C161 B.n124 VSUBS 0.006731f
C162 B.n125 VSUBS 0.006731f
C163 B.n126 VSUBS 0.006731f
C164 B.n127 VSUBS 0.006731f
C165 B.n128 VSUBS 0.006731f
C166 B.n129 VSUBS 0.006731f
C167 B.n130 VSUBS 0.006731f
C168 B.n131 VSUBS 0.006731f
C169 B.n132 VSUBS 0.006731f
C170 B.n133 VSUBS 0.006731f
C171 B.n134 VSUBS 0.006731f
C172 B.n135 VSUBS 0.006731f
C173 B.n136 VSUBS 0.006731f
C174 B.n137 VSUBS 0.014982f
C175 B.n138 VSUBS 0.014982f
C176 B.n139 VSUBS 0.016296f
C177 B.n140 VSUBS 0.006731f
C178 B.n141 VSUBS 0.006731f
C179 B.n142 VSUBS 0.006731f
C180 B.n143 VSUBS 0.006731f
C181 B.n144 VSUBS 0.006731f
C182 B.n145 VSUBS 0.006731f
C183 B.n146 VSUBS 0.006731f
C184 B.n147 VSUBS 0.006731f
C185 B.n148 VSUBS 0.006731f
C186 B.n149 VSUBS 0.006731f
C187 B.n150 VSUBS 0.006731f
C188 B.n151 VSUBS 0.006731f
C189 B.n152 VSUBS 0.006731f
C190 B.n153 VSUBS 0.006731f
C191 B.n154 VSUBS 0.006731f
C192 B.n155 VSUBS 0.006731f
C193 B.n156 VSUBS 0.006731f
C194 B.n157 VSUBS 0.006731f
C195 B.n158 VSUBS 0.006731f
C196 B.n159 VSUBS 0.006731f
C197 B.n160 VSUBS 0.006731f
C198 B.n161 VSUBS 0.006731f
C199 B.n162 VSUBS 0.006731f
C200 B.n163 VSUBS 0.006731f
C201 B.n164 VSUBS 0.006731f
C202 B.n165 VSUBS 0.006731f
C203 B.n166 VSUBS 0.006731f
C204 B.n167 VSUBS 0.006731f
C205 B.n168 VSUBS 0.006335f
C206 B.n169 VSUBS 0.015595f
C207 B.n170 VSUBS 0.003761f
C208 B.n171 VSUBS 0.006731f
C209 B.n172 VSUBS 0.006731f
C210 B.n173 VSUBS 0.006731f
C211 B.n174 VSUBS 0.006731f
C212 B.n175 VSUBS 0.006731f
C213 B.n176 VSUBS 0.006731f
C214 B.n177 VSUBS 0.006731f
C215 B.n178 VSUBS 0.006731f
C216 B.n179 VSUBS 0.006731f
C217 B.n180 VSUBS 0.006731f
C218 B.n181 VSUBS 0.006731f
C219 B.n182 VSUBS 0.006731f
C220 B.t11 VSUBS 0.064844f
C221 B.t10 VSUBS 0.084587f
C222 B.t9 VSUBS 0.49373f
C223 B.n183 VSUBS 0.147764f
C224 B.n184 VSUBS 0.123579f
C225 B.n185 VSUBS 0.015595f
C226 B.n186 VSUBS 0.003761f
C227 B.n187 VSUBS 0.006731f
C228 B.n188 VSUBS 0.006731f
C229 B.n189 VSUBS 0.006731f
C230 B.n190 VSUBS 0.006731f
C231 B.n191 VSUBS 0.006731f
C232 B.n192 VSUBS 0.006731f
C233 B.n193 VSUBS 0.006731f
C234 B.n194 VSUBS 0.006731f
C235 B.n195 VSUBS 0.006731f
C236 B.n196 VSUBS 0.006731f
C237 B.n197 VSUBS 0.006731f
C238 B.n198 VSUBS 0.006731f
C239 B.n199 VSUBS 0.006731f
C240 B.n200 VSUBS 0.006731f
C241 B.n201 VSUBS 0.006731f
C242 B.n202 VSUBS 0.006731f
C243 B.n203 VSUBS 0.006731f
C244 B.n204 VSUBS 0.006731f
C245 B.n205 VSUBS 0.006731f
C246 B.n206 VSUBS 0.006731f
C247 B.n207 VSUBS 0.006731f
C248 B.n208 VSUBS 0.006731f
C249 B.n209 VSUBS 0.006731f
C250 B.n210 VSUBS 0.006731f
C251 B.n211 VSUBS 0.006731f
C252 B.n212 VSUBS 0.006731f
C253 B.n213 VSUBS 0.006731f
C254 B.n214 VSUBS 0.006731f
C255 B.n215 VSUBS 0.006731f
C256 B.n216 VSUBS 0.015492f
C257 B.n217 VSUBS 0.016296f
C258 B.n218 VSUBS 0.014982f
C259 B.n219 VSUBS 0.006731f
C260 B.n220 VSUBS 0.006731f
C261 B.n221 VSUBS 0.006731f
C262 B.n222 VSUBS 0.006731f
C263 B.n223 VSUBS 0.006731f
C264 B.n224 VSUBS 0.006731f
C265 B.n225 VSUBS 0.006731f
C266 B.n226 VSUBS 0.006731f
C267 B.n227 VSUBS 0.006731f
C268 B.n228 VSUBS 0.006731f
C269 B.n229 VSUBS 0.006731f
C270 B.n230 VSUBS 0.006731f
C271 B.n231 VSUBS 0.006731f
C272 B.n232 VSUBS 0.006731f
C273 B.n233 VSUBS 0.006731f
C274 B.n234 VSUBS 0.006731f
C275 B.n235 VSUBS 0.006731f
C276 B.n236 VSUBS 0.006731f
C277 B.n237 VSUBS 0.006731f
C278 B.n238 VSUBS 0.006731f
C279 B.n239 VSUBS 0.006731f
C280 B.n240 VSUBS 0.006731f
C281 B.n241 VSUBS 0.006731f
C282 B.n242 VSUBS 0.006731f
C283 B.n243 VSUBS 0.006731f
C284 B.n244 VSUBS 0.006731f
C285 B.n245 VSUBS 0.006731f
C286 B.n246 VSUBS 0.006731f
C287 B.n247 VSUBS 0.006731f
C288 B.n248 VSUBS 0.006731f
C289 B.n249 VSUBS 0.006731f
C290 B.n250 VSUBS 0.006731f
C291 B.n251 VSUBS 0.006731f
C292 B.n252 VSUBS 0.006731f
C293 B.n253 VSUBS 0.006731f
C294 B.n254 VSUBS 0.006731f
C295 B.n255 VSUBS 0.006731f
C296 B.n256 VSUBS 0.006731f
C297 B.n257 VSUBS 0.006731f
C298 B.n258 VSUBS 0.006731f
C299 B.n259 VSUBS 0.006731f
C300 B.n260 VSUBS 0.006731f
C301 B.n261 VSUBS 0.006731f
C302 B.n262 VSUBS 0.006731f
C303 B.n263 VSUBS 0.006731f
C304 B.n264 VSUBS 0.006731f
C305 B.n265 VSUBS 0.006731f
C306 B.n266 VSUBS 0.006731f
C307 B.n267 VSUBS 0.006731f
C308 B.n268 VSUBS 0.006731f
C309 B.n269 VSUBS 0.006731f
C310 B.n270 VSUBS 0.006731f
C311 B.n271 VSUBS 0.006731f
C312 B.n272 VSUBS 0.006731f
C313 B.n273 VSUBS 0.006731f
C314 B.n274 VSUBS 0.006731f
C315 B.n275 VSUBS 0.006731f
C316 B.n276 VSUBS 0.006731f
C317 B.n277 VSUBS 0.006731f
C318 B.n278 VSUBS 0.006731f
C319 B.n279 VSUBS 0.006731f
C320 B.n280 VSUBS 0.006731f
C321 B.n281 VSUBS 0.006731f
C322 B.n282 VSUBS 0.006731f
C323 B.n283 VSUBS 0.006731f
C324 B.n284 VSUBS 0.006731f
C325 B.n285 VSUBS 0.006731f
C326 B.n286 VSUBS 0.006731f
C327 B.n287 VSUBS 0.006731f
C328 B.n288 VSUBS 0.014982f
C329 B.n289 VSUBS 0.014982f
C330 B.n290 VSUBS 0.016296f
C331 B.n291 VSUBS 0.006731f
C332 B.n292 VSUBS 0.006731f
C333 B.n293 VSUBS 0.006731f
C334 B.n294 VSUBS 0.006731f
C335 B.n295 VSUBS 0.006731f
C336 B.n296 VSUBS 0.006731f
C337 B.n297 VSUBS 0.006731f
C338 B.n298 VSUBS 0.006731f
C339 B.n299 VSUBS 0.006731f
C340 B.n300 VSUBS 0.006731f
C341 B.n301 VSUBS 0.006731f
C342 B.n302 VSUBS 0.006731f
C343 B.n303 VSUBS 0.006731f
C344 B.n304 VSUBS 0.006731f
C345 B.n305 VSUBS 0.006731f
C346 B.n306 VSUBS 0.006731f
C347 B.n307 VSUBS 0.006731f
C348 B.n308 VSUBS 0.006731f
C349 B.n309 VSUBS 0.006731f
C350 B.n310 VSUBS 0.006731f
C351 B.n311 VSUBS 0.006731f
C352 B.n312 VSUBS 0.006731f
C353 B.n313 VSUBS 0.006731f
C354 B.n314 VSUBS 0.006731f
C355 B.n315 VSUBS 0.006731f
C356 B.n316 VSUBS 0.006731f
C357 B.n317 VSUBS 0.006731f
C358 B.n318 VSUBS 0.006335f
C359 B.n319 VSUBS 0.006731f
C360 B.n320 VSUBS 0.006731f
C361 B.n321 VSUBS 0.006731f
C362 B.n322 VSUBS 0.006731f
C363 B.n323 VSUBS 0.006731f
C364 B.n324 VSUBS 0.006731f
C365 B.n325 VSUBS 0.006731f
C366 B.n326 VSUBS 0.006731f
C367 B.n327 VSUBS 0.006731f
C368 B.n328 VSUBS 0.006731f
C369 B.n329 VSUBS 0.006731f
C370 B.n330 VSUBS 0.006731f
C371 B.n331 VSUBS 0.006731f
C372 B.n332 VSUBS 0.006731f
C373 B.n333 VSUBS 0.006731f
C374 B.n334 VSUBS 0.003761f
C375 B.n335 VSUBS 0.015595f
C376 B.n336 VSUBS 0.006335f
C377 B.n337 VSUBS 0.006731f
C378 B.n338 VSUBS 0.006731f
C379 B.n339 VSUBS 0.006731f
C380 B.n340 VSUBS 0.006731f
C381 B.n341 VSUBS 0.006731f
C382 B.n342 VSUBS 0.006731f
C383 B.n343 VSUBS 0.006731f
C384 B.n344 VSUBS 0.006731f
C385 B.n345 VSUBS 0.006731f
C386 B.n346 VSUBS 0.006731f
C387 B.n347 VSUBS 0.006731f
C388 B.n348 VSUBS 0.006731f
C389 B.n349 VSUBS 0.006731f
C390 B.n350 VSUBS 0.006731f
C391 B.n351 VSUBS 0.006731f
C392 B.n352 VSUBS 0.006731f
C393 B.n353 VSUBS 0.006731f
C394 B.n354 VSUBS 0.006731f
C395 B.n355 VSUBS 0.006731f
C396 B.n356 VSUBS 0.006731f
C397 B.n357 VSUBS 0.006731f
C398 B.n358 VSUBS 0.006731f
C399 B.n359 VSUBS 0.006731f
C400 B.n360 VSUBS 0.006731f
C401 B.n361 VSUBS 0.006731f
C402 B.n362 VSUBS 0.006731f
C403 B.n363 VSUBS 0.006731f
C404 B.n364 VSUBS 0.016296f
C405 B.n365 VSUBS 0.016296f
C406 B.n366 VSUBS 0.014982f
C407 B.n367 VSUBS 0.006731f
C408 B.n368 VSUBS 0.006731f
C409 B.n369 VSUBS 0.006731f
C410 B.n370 VSUBS 0.006731f
C411 B.n371 VSUBS 0.006731f
C412 B.n372 VSUBS 0.006731f
C413 B.n373 VSUBS 0.006731f
C414 B.n374 VSUBS 0.006731f
C415 B.n375 VSUBS 0.006731f
C416 B.n376 VSUBS 0.006731f
C417 B.n377 VSUBS 0.006731f
C418 B.n378 VSUBS 0.006731f
C419 B.n379 VSUBS 0.006731f
C420 B.n380 VSUBS 0.006731f
C421 B.n381 VSUBS 0.006731f
C422 B.n382 VSUBS 0.006731f
C423 B.n383 VSUBS 0.006731f
C424 B.n384 VSUBS 0.006731f
C425 B.n385 VSUBS 0.006731f
C426 B.n386 VSUBS 0.006731f
C427 B.n387 VSUBS 0.006731f
C428 B.n388 VSUBS 0.006731f
C429 B.n389 VSUBS 0.006731f
C430 B.n390 VSUBS 0.006731f
C431 B.n391 VSUBS 0.006731f
C432 B.n392 VSUBS 0.006731f
C433 B.n393 VSUBS 0.006731f
C434 B.n394 VSUBS 0.006731f
C435 B.n395 VSUBS 0.006731f
C436 B.n396 VSUBS 0.006731f
C437 B.n397 VSUBS 0.006731f
C438 B.n398 VSUBS 0.006731f
C439 B.n399 VSUBS 0.008783f
C440 B.n400 VSUBS 0.009356f
C441 B.n401 VSUBS 0.018606f
C442 VDD2.n0 VSUBS 0.016757f
C443 VDD2.n1 VSUBS 0.015249f
C444 VDD2.n2 VSUBS 0.008194f
C445 VDD2.n3 VSUBS 0.019368f
C446 VDD2.n4 VSUBS 0.008676f
C447 VDD2.n5 VSUBS 0.255019f
C448 VDD2.n6 VSUBS 0.008194f
C449 VDD2.t0 VSUBS 0.042274f
C450 VDD2.n7 VSUBS 0.061965f
C451 VDD2.n8 VSUBS 0.01227f
C452 VDD2.n9 VSUBS 0.014526f
C453 VDD2.n10 VSUBS 0.019368f
C454 VDD2.n11 VSUBS 0.008676f
C455 VDD2.n12 VSUBS 0.008194f
C456 VDD2.n13 VSUBS 0.015249f
C457 VDD2.n14 VSUBS 0.015249f
C458 VDD2.n15 VSUBS 0.008194f
C459 VDD2.n16 VSUBS 0.008676f
C460 VDD2.n17 VSUBS 0.019368f
C461 VDD2.n18 VSUBS 0.046892f
C462 VDD2.n19 VSUBS 0.008676f
C463 VDD2.n20 VSUBS 0.008194f
C464 VDD2.n21 VSUBS 0.037123f
C465 VDD2.n22 VSUBS 0.28674f
C466 VDD2.n23 VSUBS 0.016757f
C467 VDD2.n24 VSUBS 0.015249f
C468 VDD2.n25 VSUBS 0.008194f
C469 VDD2.n26 VSUBS 0.019368f
C470 VDD2.n27 VSUBS 0.008676f
C471 VDD2.n28 VSUBS 0.255019f
C472 VDD2.n29 VSUBS 0.008194f
C473 VDD2.t1 VSUBS 0.042274f
C474 VDD2.n30 VSUBS 0.061965f
C475 VDD2.n31 VSUBS 0.01227f
C476 VDD2.n32 VSUBS 0.014526f
C477 VDD2.n33 VSUBS 0.019368f
C478 VDD2.n34 VSUBS 0.008676f
C479 VDD2.n35 VSUBS 0.008194f
C480 VDD2.n36 VSUBS 0.015249f
C481 VDD2.n37 VSUBS 0.015249f
C482 VDD2.n38 VSUBS 0.008194f
C483 VDD2.n39 VSUBS 0.008676f
C484 VDD2.n40 VSUBS 0.019368f
C485 VDD2.n41 VSUBS 0.046892f
C486 VDD2.n42 VSUBS 0.008676f
C487 VDD2.n43 VSUBS 0.008194f
C488 VDD2.n44 VSUBS 0.037123f
C489 VDD2.n45 VSUBS 0.034153f
C490 VDD2.n46 VSUBS 1.35892f
C491 VN.t1 VSUBS 1.41937f
C492 VN.t0 VSUBS 1.94153f
C493 VDD1.n0 VSUBS 0.016458f
C494 VDD1.n1 VSUBS 0.014977f
C495 VDD1.n2 VSUBS 0.008048f
C496 VDD1.n3 VSUBS 0.019023f
C497 VDD1.n4 VSUBS 0.008522f
C498 VDD1.n5 VSUBS 0.250468f
C499 VDD1.n6 VSUBS 0.008048f
C500 VDD1.t0 VSUBS 0.04152f
C501 VDD1.n7 VSUBS 0.06086f
C502 VDD1.n8 VSUBS 0.012051f
C503 VDD1.n9 VSUBS 0.014267f
C504 VDD1.n10 VSUBS 0.019023f
C505 VDD1.n11 VSUBS 0.008522f
C506 VDD1.n12 VSUBS 0.008048f
C507 VDD1.n13 VSUBS 0.014977f
C508 VDD1.n14 VSUBS 0.014977f
C509 VDD1.n15 VSUBS 0.008048f
C510 VDD1.n16 VSUBS 0.008522f
C511 VDD1.n17 VSUBS 0.019023f
C512 VDD1.n18 VSUBS 0.046055f
C513 VDD1.n19 VSUBS 0.008522f
C514 VDD1.n20 VSUBS 0.008048f
C515 VDD1.n21 VSUBS 0.036461f
C516 VDD1.n22 VSUBS 0.034284f
C517 VDD1.n23 VSUBS 0.016458f
C518 VDD1.n24 VSUBS 0.014977f
C519 VDD1.n25 VSUBS 0.008048f
C520 VDD1.n26 VSUBS 0.019023f
C521 VDD1.n27 VSUBS 0.008522f
C522 VDD1.n28 VSUBS 0.250468f
C523 VDD1.n29 VSUBS 0.008048f
C524 VDD1.t1 VSUBS 0.04152f
C525 VDD1.n30 VSUBS 0.06086f
C526 VDD1.n31 VSUBS 0.012051f
C527 VDD1.n32 VSUBS 0.014267f
C528 VDD1.n33 VSUBS 0.019023f
C529 VDD1.n34 VSUBS 0.008522f
C530 VDD1.n35 VSUBS 0.008048f
C531 VDD1.n36 VSUBS 0.014977f
C532 VDD1.n37 VSUBS 0.014977f
C533 VDD1.n38 VSUBS 0.008048f
C534 VDD1.n39 VSUBS 0.008522f
C535 VDD1.n40 VSUBS 0.019023f
C536 VDD1.n41 VSUBS 0.046055f
C537 VDD1.n42 VSUBS 0.008522f
C538 VDD1.n43 VSUBS 0.008048f
C539 VDD1.n44 VSUBS 0.036461f
C540 VDD1.n45 VSUBS 0.305108f
C541 VTAIL.n0 VSUBS 0.019157f
C542 VTAIL.n1 VSUBS 0.017434f
C543 VTAIL.n2 VSUBS 0.009368f
C544 VTAIL.n3 VSUBS 0.022143f
C545 VTAIL.n4 VSUBS 0.009919f
C546 VTAIL.n5 VSUBS 0.29155f
C547 VTAIL.n6 VSUBS 0.009368f
C548 VTAIL.t2 VSUBS 0.04833f
C549 VTAIL.n7 VSUBS 0.070842f
C550 VTAIL.n8 VSUBS 0.014028f
C551 VTAIL.n9 VSUBS 0.016607f
C552 VTAIL.n10 VSUBS 0.022143f
C553 VTAIL.n11 VSUBS 0.009919f
C554 VTAIL.n12 VSUBS 0.009368f
C555 VTAIL.n13 VSUBS 0.017434f
C556 VTAIL.n14 VSUBS 0.017434f
C557 VTAIL.n15 VSUBS 0.009368f
C558 VTAIL.n16 VSUBS 0.009919f
C559 VTAIL.n17 VSUBS 0.022143f
C560 VTAIL.n18 VSUBS 0.053609f
C561 VTAIL.n19 VSUBS 0.009919f
C562 VTAIL.n20 VSUBS 0.009368f
C563 VTAIL.n21 VSUBS 0.042441f
C564 VTAIL.n22 VSUBS 0.027024f
C565 VTAIL.n23 VSUBS 0.796516f
C566 VTAIL.n24 VSUBS 0.019157f
C567 VTAIL.n25 VSUBS 0.017434f
C568 VTAIL.n26 VSUBS 0.009368f
C569 VTAIL.n27 VSUBS 0.022143f
C570 VTAIL.n28 VSUBS 0.009919f
C571 VTAIL.n29 VSUBS 0.29155f
C572 VTAIL.n30 VSUBS 0.009368f
C573 VTAIL.t0 VSUBS 0.04833f
C574 VTAIL.n31 VSUBS 0.070842f
C575 VTAIL.n32 VSUBS 0.014028f
C576 VTAIL.n33 VSUBS 0.016607f
C577 VTAIL.n34 VSUBS 0.022143f
C578 VTAIL.n35 VSUBS 0.009919f
C579 VTAIL.n36 VSUBS 0.009368f
C580 VTAIL.n37 VSUBS 0.017434f
C581 VTAIL.n38 VSUBS 0.017434f
C582 VTAIL.n39 VSUBS 0.009368f
C583 VTAIL.n40 VSUBS 0.009919f
C584 VTAIL.n41 VSUBS 0.022143f
C585 VTAIL.n42 VSUBS 0.053609f
C586 VTAIL.n43 VSUBS 0.009919f
C587 VTAIL.n44 VSUBS 0.009368f
C588 VTAIL.n45 VSUBS 0.042441f
C589 VTAIL.n46 VSUBS 0.027024f
C590 VTAIL.n47 VSUBS 0.82533f
C591 VTAIL.n48 VSUBS 0.019157f
C592 VTAIL.n49 VSUBS 0.017434f
C593 VTAIL.n50 VSUBS 0.009368f
C594 VTAIL.n51 VSUBS 0.022143f
C595 VTAIL.n52 VSUBS 0.009919f
C596 VTAIL.n53 VSUBS 0.29155f
C597 VTAIL.n54 VSUBS 0.009368f
C598 VTAIL.t3 VSUBS 0.04833f
C599 VTAIL.n55 VSUBS 0.070842f
C600 VTAIL.n56 VSUBS 0.014028f
C601 VTAIL.n57 VSUBS 0.016607f
C602 VTAIL.n58 VSUBS 0.022143f
C603 VTAIL.n59 VSUBS 0.009919f
C604 VTAIL.n60 VSUBS 0.009368f
C605 VTAIL.n61 VSUBS 0.017434f
C606 VTAIL.n62 VSUBS 0.017434f
C607 VTAIL.n63 VSUBS 0.009368f
C608 VTAIL.n64 VSUBS 0.009919f
C609 VTAIL.n65 VSUBS 0.022143f
C610 VTAIL.n66 VSUBS 0.053609f
C611 VTAIL.n67 VSUBS 0.009919f
C612 VTAIL.n68 VSUBS 0.009368f
C613 VTAIL.n69 VSUBS 0.042441f
C614 VTAIL.n70 VSUBS 0.027024f
C615 VTAIL.n71 VSUBS 0.696998f
C616 VTAIL.n72 VSUBS 0.019157f
C617 VTAIL.n73 VSUBS 0.017434f
C618 VTAIL.n74 VSUBS 0.009368f
C619 VTAIL.n75 VSUBS 0.022143f
C620 VTAIL.n76 VSUBS 0.009919f
C621 VTAIL.n77 VSUBS 0.29155f
C622 VTAIL.n78 VSUBS 0.009368f
C623 VTAIL.t1 VSUBS 0.04833f
C624 VTAIL.n79 VSUBS 0.070842f
C625 VTAIL.n80 VSUBS 0.014028f
C626 VTAIL.n81 VSUBS 0.016607f
C627 VTAIL.n82 VSUBS 0.022143f
C628 VTAIL.n83 VSUBS 0.009919f
C629 VTAIL.n84 VSUBS 0.009368f
C630 VTAIL.n85 VSUBS 0.017434f
C631 VTAIL.n86 VSUBS 0.017434f
C632 VTAIL.n87 VSUBS 0.009368f
C633 VTAIL.n88 VSUBS 0.009919f
C634 VTAIL.n89 VSUBS 0.022143f
C635 VTAIL.n90 VSUBS 0.053609f
C636 VTAIL.n91 VSUBS 0.009919f
C637 VTAIL.n92 VSUBS 0.009368f
C638 VTAIL.n93 VSUBS 0.042441f
C639 VTAIL.n94 VSUBS 0.027024f
C640 VTAIL.n95 VSUBS 0.635253f
C641 VP.t1 VSUBS 2.0412f
C642 VP.t0 VSUBS 1.49447f
C643 VP.n0 VSUBS 3.27737f
.ends

