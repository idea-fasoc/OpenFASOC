* NGSPICE file created from diff_pair_sample_0208.ext - technology: sky130A

.subckt diff_pair_sample_0208 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t3 VN.t0 VTAIL.t7 B.t0 sky130_fd_pr__nfet_01v8 ad=0.8019 pd=5.19 as=1.8954 ps=10.5 w=4.86 l=3.77
X1 VDD1.t3 VP.t0 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=0.8019 pd=5.19 as=1.8954 ps=10.5 w=4.86 l=3.77
X2 B.t17 B.t15 B.t16 B.t12 sky130_fd_pr__nfet_01v8 ad=1.8954 pd=10.5 as=0 ps=0 w=4.86 l=3.77
X3 B.t14 B.t11 B.t13 B.t12 sky130_fd_pr__nfet_01v8 ad=1.8954 pd=10.5 as=0 ps=0 w=4.86 l=3.77
X4 B.t10 B.t8 B.t9 B.t5 sky130_fd_pr__nfet_01v8 ad=1.8954 pd=10.5 as=0 ps=0 w=4.86 l=3.77
X5 VTAIL.t1 VP.t1 VDD1.t2 B.t1 sky130_fd_pr__nfet_01v8 ad=1.8954 pd=10.5 as=0.8019 ps=5.19 w=4.86 l=3.77
X6 VDD2.t2 VN.t1 VTAIL.t5 B.t2 sky130_fd_pr__nfet_01v8 ad=0.8019 pd=5.19 as=1.8954 ps=10.5 w=4.86 l=3.77
X7 B.t7 B.t4 B.t6 B.t5 sky130_fd_pr__nfet_01v8 ad=1.8954 pd=10.5 as=0 ps=0 w=4.86 l=3.77
X8 VTAIL.t6 VN.t2 VDD2.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=1.8954 pd=10.5 as=0.8019 ps=5.19 w=4.86 l=3.77
X9 VDD1.t1 VP.t2 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=0.8019 pd=5.19 as=1.8954 ps=10.5 w=4.86 l=3.77
X10 VTAIL.t3 VP.t3 VDD1.t0 B.t3 sky130_fd_pr__nfet_01v8 ad=1.8954 pd=10.5 as=0.8019 ps=5.19 w=4.86 l=3.77
X11 VTAIL.t4 VN.t3 VDD2.t0 B.t3 sky130_fd_pr__nfet_01v8 ad=1.8954 pd=10.5 as=0.8019 ps=5.19 w=4.86 l=3.77
R0 VN.n1 VN.t1 64.8929
R1 VN.n0 VN.t3 64.8929
R2 VN.n0 VN.t0 63.5492
R3 VN.n1 VN.t2 63.5492
R4 VN VN.n1 46.5598
R5 VN VN.n0 1.87422
R6 VTAIL.n5 VTAIL.t3 55.7987
R7 VTAIL.n4 VTAIL.t5 55.7987
R8 VTAIL.n3 VTAIL.t6 55.7987
R9 VTAIL.n7 VTAIL.t7 55.7986
R10 VTAIL.n0 VTAIL.t4 55.7986
R11 VTAIL.n1 VTAIL.t2 55.7986
R12 VTAIL.n2 VTAIL.t1 55.7986
R13 VTAIL.n6 VTAIL.t0 55.7986
R14 VTAIL.n7 VTAIL.n6 20.091
R15 VTAIL.n3 VTAIL.n2 20.091
R16 VTAIL.n4 VTAIL.n3 3.53498
R17 VTAIL.n6 VTAIL.n5 3.53498
R18 VTAIL.n2 VTAIL.n1 3.53498
R19 VTAIL VTAIL.n0 1.82593
R20 VTAIL VTAIL.n7 1.70955
R21 VTAIL.n5 VTAIL.n4 0.470328
R22 VTAIL.n1 VTAIL.n0 0.470328
R23 VDD2.n2 VDD2.n0 106.912
R24 VDD2.n2 VDD2.n1 68.4033
R25 VDD2.n1 VDD2.t1 4.07457
R26 VDD2.n1 VDD2.t2 4.07457
R27 VDD2.n0 VDD2.t0 4.07457
R28 VDD2.n0 VDD2.t3 4.07457
R29 VDD2 VDD2.n2 0.0586897
R30 B.n623 B.n622 585
R31 B.n624 B.n623 585
R32 B.n212 B.n109 585
R33 B.n211 B.n210 585
R34 B.n209 B.n208 585
R35 B.n207 B.n206 585
R36 B.n205 B.n204 585
R37 B.n203 B.n202 585
R38 B.n201 B.n200 585
R39 B.n199 B.n198 585
R40 B.n197 B.n196 585
R41 B.n195 B.n194 585
R42 B.n193 B.n192 585
R43 B.n191 B.n190 585
R44 B.n189 B.n188 585
R45 B.n187 B.n186 585
R46 B.n185 B.n184 585
R47 B.n183 B.n182 585
R48 B.n181 B.n180 585
R49 B.n179 B.n178 585
R50 B.n177 B.n176 585
R51 B.n175 B.n174 585
R52 B.n173 B.n172 585
R53 B.n171 B.n170 585
R54 B.n169 B.n168 585
R55 B.n167 B.n166 585
R56 B.n165 B.n164 585
R57 B.n163 B.n162 585
R58 B.n161 B.n160 585
R59 B.n159 B.n158 585
R60 B.n157 B.n156 585
R61 B.n154 B.n153 585
R62 B.n152 B.n151 585
R63 B.n150 B.n149 585
R64 B.n148 B.n147 585
R65 B.n146 B.n145 585
R66 B.n144 B.n143 585
R67 B.n142 B.n141 585
R68 B.n140 B.n139 585
R69 B.n138 B.n137 585
R70 B.n136 B.n135 585
R71 B.n134 B.n133 585
R72 B.n132 B.n131 585
R73 B.n130 B.n129 585
R74 B.n128 B.n127 585
R75 B.n126 B.n125 585
R76 B.n124 B.n123 585
R77 B.n122 B.n121 585
R78 B.n120 B.n119 585
R79 B.n118 B.n117 585
R80 B.n116 B.n115 585
R81 B.n82 B.n81 585
R82 B.n621 B.n83 585
R83 B.n625 B.n83 585
R84 B.n620 B.n619 585
R85 B.n619 B.n79 585
R86 B.n618 B.n78 585
R87 B.n631 B.n78 585
R88 B.n617 B.n77 585
R89 B.n632 B.n77 585
R90 B.n616 B.n76 585
R91 B.n633 B.n76 585
R92 B.n615 B.n614 585
R93 B.n614 B.n72 585
R94 B.n613 B.n71 585
R95 B.n639 B.n71 585
R96 B.n612 B.n70 585
R97 B.n640 B.n70 585
R98 B.n611 B.n69 585
R99 B.n641 B.n69 585
R100 B.n610 B.n609 585
R101 B.n609 B.n68 585
R102 B.n608 B.n64 585
R103 B.n647 B.n64 585
R104 B.n607 B.n63 585
R105 B.n648 B.n63 585
R106 B.n606 B.n62 585
R107 B.n649 B.n62 585
R108 B.n605 B.n604 585
R109 B.n604 B.n58 585
R110 B.n603 B.n57 585
R111 B.n655 B.n57 585
R112 B.n602 B.n56 585
R113 B.n656 B.n56 585
R114 B.n601 B.n55 585
R115 B.n657 B.n55 585
R116 B.n600 B.n599 585
R117 B.n599 B.n51 585
R118 B.n598 B.n50 585
R119 B.n663 B.n50 585
R120 B.n597 B.n49 585
R121 B.n664 B.n49 585
R122 B.n596 B.n48 585
R123 B.n665 B.n48 585
R124 B.n595 B.n594 585
R125 B.n594 B.n44 585
R126 B.n593 B.n43 585
R127 B.n671 B.n43 585
R128 B.n592 B.n42 585
R129 B.n672 B.n42 585
R130 B.n591 B.n41 585
R131 B.n673 B.n41 585
R132 B.n590 B.n589 585
R133 B.n589 B.n37 585
R134 B.n588 B.n36 585
R135 B.n679 B.n36 585
R136 B.n587 B.n35 585
R137 B.n680 B.n35 585
R138 B.n586 B.n34 585
R139 B.n681 B.n34 585
R140 B.n585 B.n584 585
R141 B.n584 B.n30 585
R142 B.n583 B.n29 585
R143 B.n687 B.n29 585
R144 B.n582 B.n28 585
R145 B.n688 B.n28 585
R146 B.n581 B.n27 585
R147 B.n689 B.n27 585
R148 B.n580 B.n579 585
R149 B.n579 B.n23 585
R150 B.n578 B.n22 585
R151 B.n695 B.n22 585
R152 B.n577 B.n21 585
R153 B.n696 B.n21 585
R154 B.n576 B.n20 585
R155 B.n697 B.n20 585
R156 B.n575 B.n574 585
R157 B.n574 B.n16 585
R158 B.n573 B.n15 585
R159 B.n703 B.n15 585
R160 B.n572 B.n14 585
R161 B.n704 B.n14 585
R162 B.n571 B.n13 585
R163 B.n705 B.n13 585
R164 B.n570 B.n569 585
R165 B.n569 B.n12 585
R166 B.n568 B.n567 585
R167 B.n568 B.n8 585
R168 B.n566 B.n7 585
R169 B.n712 B.n7 585
R170 B.n565 B.n6 585
R171 B.n713 B.n6 585
R172 B.n564 B.n5 585
R173 B.n714 B.n5 585
R174 B.n563 B.n562 585
R175 B.n562 B.n4 585
R176 B.n561 B.n213 585
R177 B.n561 B.n560 585
R178 B.n551 B.n214 585
R179 B.n215 B.n214 585
R180 B.n553 B.n552 585
R181 B.n554 B.n553 585
R182 B.n550 B.n220 585
R183 B.n220 B.n219 585
R184 B.n549 B.n548 585
R185 B.n548 B.n547 585
R186 B.n222 B.n221 585
R187 B.n223 B.n222 585
R188 B.n540 B.n539 585
R189 B.n541 B.n540 585
R190 B.n538 B.n228 585
R191 B.n228 B.n227 585
R192 B.n537 B.n536 585
R193 B.n536 B.n535 585
R194 B.n230 B.n229 585
R195 B.n231 B.n230 585
R196 B.n528 B.n527 585
R197 B.n529 B.n528 585
R198 B.n526 B.n236 585
R199 B.n236 B.n235 585
R200 B.n525 B.n524 585
R201 B.n524 B.n523 585
R202 B.n238 B.n237 585
R203 B.n239 B.n238 585
R204 B.n516 B.n515 585
R205 B.n517 B.n516 585
R206 B.n514 B.n244 585
R207 B.n244 B.n243 585
R208 B.n513 B.n512 585
R209 B.n512 B.n511 585
R210 B.n246 B.n245 585
R211 B.n247 B.n246 585
R212 B.n504 B.n503 585
R213 B.n505 B.n504 585
R214 B.n502 B.n252 585
R215 B.n252 B.n251 585
R216 B.n501 B.n500 585
R217 B.n500 B.n499 585
R218 B.n254 B.n253 585
R219 B.n255 B.n254 585
R220 B.n492 B.n491 585
R221 B.n493 B.n492 585
R222 B.n490 B.n260 585
R223 B.n260 B.n259 585
R224 B.n489 B.n488 585
R225 B.n488 B.n487 585
R226 B.n262 B.n261 585
R227 B.n263 B.n262 585
R228 B.n480 B.n479 585
R229 B.n481 B.n480 585
R230 B.n478 B.n268 585
R231 B.n268 B.n267 585
R232 B.n477 B.n476 585
R233 B.n476 B.n475 585
R234 B.n270 B.n269 585
R235 B.n271 B.n270 585
R236 B.n468 B.n467 585
R237 B.n469 B.n468 585
R238 B.n466 B.n276 585
R239 B.n276 B.n275 585
R240 B.n465 B.n464 585
R241 B.n464 B.n463 585
R242 B.n278 B.n277 585
R243 B.n456 B.n278 585
R244 B.n455 B.n454 585
R245 B.n457 B.n455 585
R246 B.n453 B.n283 585
R247 B.n283 B.n282 585
R248 B.n452 B.n451 585
R249 B.n451 B.n450 585
R250 B.n285 B.n284 585
R251 B.n286 B.n285 585
R252 B.n443 B.n442 585
R253 B.n444 B.n443 585
R254 B.n441 B.n291 585
R255 B.n291 B.n290 585
R256 B.n440 B.n439 585
R257 B.n439 B.n438 585
R258 B.n293 B.n292 585
R259 B.n294 B.n293 585
R260 B.n431 B.n430 585
R261 B.n432 B.n431 585
R262 B.n297 B.n296 585
R263 B.n331 B.n330 585
R264 B.n332 B.n328 585
R265 B.n328 B.n298 585
R266 B.n334 B.n333 585
R267 B.n336 B.n327 585
R268 B.n339 B.n338 585
R269 B.n340 B.n326 585
R270 B.n342 B.n341 585
R271 B.n344 B.n325 585
R272 B.n347 B.n346 585
R273 B.n348 B.n324 585
R274 B.n350 B.n349 585
R275 B.n352 B.n323 585
R276 B.n355 B.n354 585
R277 B.n356 B.n322 585
R278 B.n358 B.n357 585
R279 B.n360 B.n321 585
R280 B.n363 B.n362 585
R281 B.n364 B.n320 585
R282 B.n366 B.n365 585
R283 B.n368 B.n319 585
R284 B.n371 B.n370 585
R285 B.n372 B.n315 585
R286 B.n374 B.n373 585
R287 B.n376 B.n314 585
R288 B.n379 B.n378 585
R289 B.n380 B.n313 585
R290 B.n382 B.n381 585
R291 B.n384 B.n312 585
R292 B.n387 B.n386 585
R293 B.n389 B.n309 585
R294 B.n391 B.n390 585
R295 B.n393 B.n308 585
R296 B.n396 B.n395 585
R297 B.n397 B.n307 585
R298 B.n399 B.n398 585
R299 B.n401 B.n306 585
R300 B.n404 B.n403 585
R301 B.n405 B.n305 585
R302 B.n407 B.n406 585
R303 B.n409 B.n304 585
R304 B.n412 B.n411 585
R305 B.n413 B.n303 585
R306 B.n415 B.n414 585
R307 B.n417 B.n302 585
R308 B.n420 B.n419 585
R309 B.n421 B.n301 585
R310 B.n423 B.n422 585
R311 B.n425 B.n300 585
R312 B.n428 B.n427 585
R313 B.n429 B.n299 585
R314 B.n434 B.n433 585
R315 B.n433 B.n432 585
R316 B.n435 B.n295 585
R317 B.n295 B.n294 585
R318 B.n437 B.n436 585
R319 B.n438 B.n437 585
R320 B.n289 B.n288 585
R321 B.n290 B.n289 585
R322 B.n446 B.n445 585
R323 B.n445 B.n444 585
R324 B.n447 B.n287 585
R325 B.n287 B.n286 585
R326 B.n449 B.n448 585
R327 B.n450 B.n449 585
R328 B.n281 B.n280 585
R329 B.n282 B.n281 585
R330 B.n459 B.n458 585
R331 B.n458 B.n457 585
R332 B.n460 B.n279 585
R333 B.n456 B.n279 585
R334 B.n462 B.n461 585
R335 B.n463 B.n462 585
R336 B.n274 B.n273 585
R337 B.n275 B.n274 585
R338 B.n471 B.n470 585
R339 B.n470 B.n469 585
R340 B.n472 B.n272 585
R341 B.n272 B.n271 585
R342 B.n474 B.n473 585
R343 B.n475 B.n474 585
R344 B.n266 B.n265 585
R345 B.n267 B.n266 585
R346 B.n483 B.n482 585
R347 B.n482 B.n481 585
R348 B.n484 B.n264 585
R349 B.n264 B.n263 585
R350 B.n486 B.n485 585
R351 B.n487 B.n486 585
R352 B.n258 B.n257 585
R353 B.n259 B.n258 585
R354 B.n495 B.n494 585
R355 B.n494 B.n493 585
R356 B.n496 B.n256 585
R357 B.n256 B.n255 585
R358 B.n498 B.n497 585
R359 B.n499 B.n498 585
R360 B.n250 B.n249 585
R361 B.n251 B.n250 585
R362 B.n507 B.n506 585
R363 B.n506 B.n505 585
R364 B.n508 B.n248 585
R365 B.n248 B.n247 585
R366 B.n510 B.n509 585
R367 B.n511 B.n510 585
R368 B.n242 B.n241 585
R369 B.n243 B.n242 585
R370 B.n519 B.n518 585
R371 B.n518 B.n517 585
R372 B.n520 B.n240 585
R373 B.n240 B.n239 585
R374 B.n522 B.n521 585
R375 B.n523 B.n522 585
R376 B.n234 B.n233 585
R377 B.n235 B.n234 585
R378 B.n531 B.n530 585
R379 B.n530 B.n529 585
R380 B.n532 B.n232 585
R381 B.n232 B.n231 585
R382 B.n534 B.n533 585
R383 B.n535 B.n534 585
R384 B.n226 B.n225 585
R385 B.n227 B.n226 585
R386 B.n543 B.n542 585
R387 B.n542 B.n541 585
R388 B.n544 B.n224 585
R389 B.n224 B.n223 585
R390 B.n546 B.n545 585
R391 B.n547 B.n546 585
R392 B.n218 B.n217 585
R393 B.n219 B.n218 585
R394 B.n556 B.n555 585
R395 B.n555 B.n554 585
R396 B.n557 B.n216 585
R397 B.n216 B.n215 585
R398 B.n559 B.n558 585
R399 B.n560 B.n559 585
R400 B.n3 B.n0 585
R401 B.n4 B.n3 585
R402 B.n711 B.n1 585
R403 B.n712 B.n711 585
R404 B.n710 B.n709 585
R405 B.n710 B.n8 585
R406 B.n708 B.n9 585
R407 B.n12 B.n9 585
R408 B.n707 B.n706 585
R409 B.n706 B.n705 585
R410 B.n11 B.n10 585
R411 B.n704 B.n11 585
R412 B.n702 B.n701 585
R413 B.n703 B.n702 585
R414 B.n700 B.n17 585
R415 B.n17 B.n16 585
R416 B.n699 B.n698 585
R417 B.n698 B.n697 585
R418 B.n19 B.n18 585
R419 B.n696 B.n19 585
R420 B.n694 B.n693 585
R421 B.n695 B.n694 585
R422 B.n692 B.n24 585
R423 B.n24 B.n23 585
R424 B.n691 B.n690 585
R425 B.n690 B.n689 585
R426 B.n26 B.n25 585
R427 B.n688 B.n26 585
R428 B.n686 B.n685 585
R429 B.n687 B.n686 585
R430 B.n684 B.n31 585
R431 B.n31 B.n30 585
R432 B.n683 B.n682 585
R433 B.n682 B.n681 585
R434 B.n33 B.n32 585
R435 B.n680 B.n33 585
R436 B.n678 B.n677 585
R437 B.n679 B.n678 585
R438 B.n676 B.n38 585
R439 B.n38 B.n37 585
R440 B.n675 B.n674 585
R441 B.n674 B.n673 585
R442 B.n40 B.n39 585
R443 B.n672 B.n40 585
R444 B.n670 B.n669 585
R445 B.n671 B.n670 585
R446 B.n668 B.n45 585
R447 B.n45 B.n44 585
R448 B.n667 B.n666 585
R449 B.n666 B.n665 585
R450 B.n47 B.n46 585
R451 B.n664 B.n47 585
R452 B.n662 B.n661 585
R453 B.n663 B.n662 585
R454 B.n660 B.n52 585
R455 B.n52 B.n51 585
R456 B.n659 B.n658 585
R457 B.n658 B.n657 585
R458 B.n54 B.n53 585
R459 B.n656 B.n54 585
R460 B.n654 B.n653 585
R461 B.n655 B.n654 585
R462 B.n652 B.n59 585
R463 B.n59 B.n58 585
R464 B.n651 B.n650 585
R465 B.n650 B.n649 585
R466 B.n61 B.n60 585
R467 B.n648 B.n61 585
R468 B.n646 B.n645 585
R469 B.n647 B.n646 585
R470 B.n644 B.n65 585
R471 B.n68 B.n65 585
R472 B.n643 B.n642 585
R473 B.n642 B.n641 585
R474 B.n67 B.n66 585
R475 B.n640 B.n67 585
R476 B.n638 B.n637 585
R477 B.n639 B.n638 585
R478 B.n636 B.n73 585
R479 B.n73 B.n72 585
R480 B.n635 B.n634 585
R481 B.n634 B.n633 585
R482 B.n75 B.n74 585
R483 B.n632 B.n75 585
R484 B.n630 B.n629 585
R485 B.n631 B.n630 585
R486 B.n628 B.n80 585
R487 B.n80 B.n79 585
R488 B.n627 B.n626 585
R489 B.n626 B.n625 585
R490 B.n715 B.n714 585
R491 B.n713 B.n2 585
R492 B.n626 B.n82 449.257
R493 B.n623 B.n83 449.257
R494 B.n431 B.n299 449.257
R495 B.n433 B.n297 449.257
R496 B.n624 B.n108 256.663
R497 B.n624 B.n107 256.663
R498 B.n624 B.n106 256.663
R499 B.n624 B.n105 256.663
R500 B.n624 B.n104 256.663
R501 B.n624 B.n103 256.663
R502 B.n624 B.n102 256.663
R503 B.n624 B.n101 256.663
R504 B.n624 B.n100 256.663
R505 B.n624 B.n99 256.663
R506 B.n624 B.n98 256.663
R507 B.n624 B.n97 256.663
R508 B.n624 B.n96 256.663
R509 B.n624 B.n95 256.663
R510 B.n624 B.n94 256.663
R511 B.n624 B.n93 256.663
R512 B.n624 B.n92 256.663
R513 B.n624 B.n91 256.663
R514 B.n624 B.n90 256.663
R515 B.n624 B.n89 256.663
R516 B.n624 B.n88 256.663
R517 B.n624 B.n87 256.663
R518 B.n624 B.n86 256.663
R519 B.n624 B.n85 256.663
R520 B.n624 B.n84 256.663
R521 B.n329 B.n298 256.663
R522 B.n335 B.n298 256.663
R523 B.n337 B.n298 256.663
R524 B.n343 B.n298 256.663
R525 B.n345 B.n298 256.663
R526 B.n351 B.n298 256.663
R527 B.n353 B.n298 256.663
R528 B.n359 B.n298 256.663
R529 B.n361 B.n298 256.663
R530 B.n367 B.n298 256.663
R531 B.n369 B.n298 256.663
R532 B.n375 B.n298 256.663
R533 B.n377 B.n298 256.663
R534 B.n383 B.n298 256.663
R535 B.n385 B.n298 256.663
R536 B.n392 B.n298 256.663
R537 B.n394 B.n298 256.663
R538 B.n400 B.n298 256.663
R539 B.n402 B.n298 256.663
R540 B.n408 B.n298 256.663
R541 B.n410 B.n298 256.663
R542 B.n416 B.n298 256.663
R543 B.n418 B.n298 256.663
R544 B.n424 B.n298 256.663
R545 B.n426 B.n298 256.663
R546 B.n717 B.n716 256.663
R547 B.n113 B.t8 240.388
R548 B.n110 B.t4 240.388
R549 B.n310 B.t15 240.388
R550 B.n316 B.t11 240.388
R551 B.n117 B.n116 163.367
R552 B.n121 B.n120 163.367
R553 B.n125 B.n124 163.367
R554 B.n129 B.n128 163.367
R555 B.n133 B.n132 163.367
R556 B.n137 B.n136 163.367
R557 B.n141 B.n140 163.367
R558 B.n145 B.n144 163.367
R559 B.n149 B.n148 163.367
R560 B.n153 B.n152 163.367
R561 B.n158 B.n157 163.367
R562 B.n162 B.n161 163.367
R563 B.n166 B.n165 163.367
R564 B.n170 B.n169 163.367
R565 B.n174 B.n173 163.367
R566 B.n178 B.n177 163.367
R567 B.n182 B.n181 163.367
R568 B.n186 B.n185 163.367
R569 B.n190 B.n189 163.367
R570 B.n194 B.n193 163.367
R571 B.n198 B.n197 163.367
R572 B.n202 B.n201 163.367
R573 B.n206 B.n205 163.367
R574 B.n210 B.n209 163.367
R575 B.n623 B.n109 163.367
R576 B.n431 B.n293 163.367
R577 B.n439 B.n293 163.367
R578 B.n439 B.n291 163.367
R579 B.n443 B.n291 163.367
R580 B.n443 B.n285 163.367
R581 B.n451 B.n285 163.367
R582 B.n451 B.n283 163.367
R583 B.n455 B.n283 163.367
R584 B.n455 B.n278 163.367
R585 B.n464 B.n278 163.367
R586 B.n464 B.n276 163.367
R587 B.n468 B.n276 163.367
R588 B.n468 B.n270 163.367
R589 B.n476 B.n270 163.367
R590 B.n476 B.n268 163.367
R591 B.n480 B.n268 163.367
R592 B.n480 B.n262 163.367
R593 B.n488 B.n262 163.367
R594 B.n488 B.n260 163.367
R595 B.n492 B.n260 163.367
R596 B.n492 B.n254 163.367
R597 B.n500 B.n254 163.367
R598 B.n500 B.n252 163.367
R599 B.n504 B.n252 163.367
R600 B.n504 B.n246 163.367
R601 B.n512 B.n246 163.367
R602 B.n512 B.n244 163.367
R603 B.n516 B.n244 163.367
R604 B.n516 B.n238 163.367
R605 B.n524 B.n238 163.367
R606 B.n524 B.n236 163.367
R607 B.n528 B.n236 163.367
R608 B.n528 B.n230 163.367
R609 B.n536 B.n230 163.367
R610 B.n536 B.n228 163.367
R611 B.n540 B.n228 163.367
R612 B.n540 B.n222 163.367
R613 B.n548 B.n222 163.367
R614 B.n548 B.n220 163.367
R615 B.n553 B.n220 163.367
R616 B.n553 B.n214 163.367
R617 B.n561 B.n214 163.367
R618 B.n562 B.n561 163.367
R619 B.n562 B.n5 163.367
R620 B.n6 B.n5 163.367
R621 B.n7 B.n6 163.367
R622 B.n568 B.n7 163.367
R623 B.n569 B.n568 163.367
R624 B.n569 B.n13 163.367
R625 B.n14 B.n13 163.367
R626 B.n15 B.n14 163.367
R627 B.n574 B.n15 163.367
R628 B.n574 B.n20 163.367
R629 B.n21 B.n20 163.367
R630 B.n22 B.n21 163.367
R631 B.n579 B.n22 163.367
R632 B.n579 B.n27 163.367
R633 B.n28 B.n27 163.367
R634 B.n29 B.n28 163.367
R635 B.n584 B.n29 163.367
R636 B.n584 B.n34 163.367
R637 B.n35 B.n34 163.367
R638 B.n36 B.n35 163.367
R639 B.n589 B.n36 163.367
R640 B.n589 B.n41 163.367
R641 B.n42 B.n41 163.367
R642 B.n43 B.n42 163.367
R643 B.n594 B.n43 163.367
R644 B.n594 B.n48 163.367
R645 B.n49 B.n48 163.367
R646 B.n50 B.n49 163.367
R647 B.n599 B.n50 163.367
R648 B.n599 B.n55 163.367
R649 B.n56 B.n55 163.367
R650 B.n57 B.n56 163.367
R651 B.n604 B.n57 163.367
R652 B.n604 B.n62 163.367
R653 B.n63 B.n62 163.367
R654 B.n64 B.n63 163.367
R655 B.n609 B.n64 163.367
R656 B.n609 B.n69 163.367
R657 B.n70 B.n69 163.367
R658 B.n71 B.n70 163.367
R659 B.n614 B.n71 163.367
R660 B.n614 B.n76 163.367
R661 B.n77 B.n76 163.367
R662 B.n78 B.n77 163.367
R663 B.n619 B.n78 163.367
R664 B.n619 B.n83 163.367
R665 B.n330 B.n328 163.367
R666 B.n334 B.n328 163.367
R667 B.n338 B.n336 163.367
R668 B.n342 B.n326 163.367
R669 B.n346 B.n344 163.367
R670 B.n350 B.n324 163.367
R671 B.n354 B.n352 163.367
R672 B.n358 B.n322 163.367
R673 B.n362 B.n360 163.367
R674 B.n366 B.n320 163.367
R675 B.n370 B.n368 163.367
R676 B.n374 B.n315 163.367
R677 B.n378 B.n376 163.367
R678 B.n382 B.n313 163.367
R679 B.n386 B.n384 163.367
R680 B.n391 B.n309 163.367
R681 B.n395 B.n393 163.367
R682 B.n399 B.n307 163.367
R683 B.n403 B.n401 163.367
R684 B.n407 B.n305 163.367
R685 B.n411 B.n409 163.367
R686 B.n415 B.n303 163.367
R687 B.n419 B.n417 163.367
R688 B.n423 B.n301 163.367
R689 B.n427 B.n425 163.367
R690 B.n433 B.n295 163.367
R691 B.n437 B.n295 163.367
R692 B.n437 B.n289 163.367
R693 B.n445 B.n289 163.367
R694 B.n445 B.n287 163.367
R695 B.n449 B.n287 163.367
R696 B.n449 B.n281 163.367
R697 B.n458 B.n281 163.367
R698 B.n458 B.n279 163.367
R699 B.n462 B.n279 163.367
R700 B.n462 B.n274 163.367
R701 B.n470 B.n274 163.367
R702 B.n470 B.n272 163.367
R703 B.n474 B.n272 163.367
R704 B.n474 B.n266 163.367
R705 B.n482 B.n266 163.367
R706 B.n482 B.n264 163.367
R707 B.n486 B.n264 163.367
R708 B.n486 B.n258 163.367
R709 B.n494 B.n258 163.367
R710 B.n494 B.n256 163.367
R711 B.n498 B.n256 163.367
R712 B.n498 B.n250 163.367
R713 B.n506 B.n250 163.367
R714 B.n506 B.n248 163.367
R715 B.n510 B.n248 163.367
R716 B.n510 B.n242 163.367
R717 B.n518 B.n242 163.367
R718 B.n518 B.n240 163.367
R719 B.n522 B.n240 163.367
R720 B.n522 B.n234 163.367
R721 B.n530 B.n234 163.367
R722 B.n530 B.n232 163.367
R723 B.n534 B.n232 163.367
R724 B.n534 B.n226 163.367
R725 B.n542 B.n226 163.367
R726 B.n542 B.n224 163.367
R727 B.n546 B.n224 163.367
R728 B.n546 B.n218 163.367
R729 B.n555 B.n218 163.367
R730 B.n555 B.n216 163.367
R731 B.n559 B.n216 163.367
R732 B.n559 B.n3 163.367
R733 B.n715 B.n3 163.367
R734 B.n711 B.n2 163.367
R735 B.n711 B.n710 163.367
R736 B.n710 B.n9 163.367
R737 B.n706 B.n9 163.367
R738 B.n706 B.n11 163.367
R739 B.n702 B.n11 163.367
R740 B.n702 B.n17 163.367
R741 B.n698 B.n17 163.367
R742 B.n698 B.n19 163.367
R743 B.n694 B.n19 163.367
R744 B.n694 B.n24 163.367
R745 B.n690 B.n24 163.367
R746 B.n690 B.n26 163.367
R747 B.n686 B.n26 163.367
R748 B.n686 B.n31 163.367
R749 B.n682 B.n31 163.367
R750 B.n682 B.n33 163.367
R751 B.n678 B.n33 163.367
R752 B.n678 B.n38 163.367
R753 B.n674 B.n38 163.367
R754 B.n674 B.n40 163.367
R755 B.n670 B.n40 163.367
R756 B.n670 B.n45 163.367
R757 B.n666 B.n45 163.367
R758 B.n666 B.n47 163.367
R759 B.n662 B.n47 163.367
R760 B.n662 B.n52 163.367
R761 B.n658 B.n52 163.367
R762 B.n658 B.n54 163.367
R763 B.n654 B.n54 163.367
R764 B.n654 B.n59 163.367
R765 B.n650 B.n59 163.367
R766 B.n650 B.n61 163.367
R767 B.n646 B.n61 163.367
R768 B.n646 B.n65 163.367
R769 B.n642 B.n65 163.367
R770 B.n642 B.n67 163.367
R771 B.n638 B.n67 163.367
R772 B.n638 B.n73 163.367
R773 B.n634 B.n73 163.367
R774 B.n634 B.n75 163.367
R775 B.n630 B.n75 163.367
R776 B.n630 B.n80 163.367
R777 B.n626 B.n80 163.367
R778 B.n110 B.t6 151.756
R779 B.n310 B.t17 151.756
R780 B.n113 B.t9 151.751
R781 B.n316 B.t14 151.751
R782 B.n432 B.n298 118.303
R783 B.n625 B.n624 118.303
R784 B.n114 B.n113 79.5157
R785 B.n111 B.n110 79.5157
R786 B.n311 B.n310 79.5157
R787 B.n317 B.n316 79.5157
R788 B.n432 B.n294 73.8041
R789 B.n438 B.n294 73.8041
R790 B.n438 B.n290 73.8041
R791 B.n444 B.n290 73.8041
R792 B.n444 B.n286 73.8041
R793 B.n450 B.n286 73.8041
R794 B.n450 B.n282 73.8041
R795 B.n457 B.n282 73.8041
R796 B.n457 B.n456 73.8041
R797 B.n463 B.n275 73.8041
R798 B.n469 B.n275 73.8041
R799 B.n469 B.n271 73.8041
R800 B.n475 B.n271 73.8041
R801 B.n475 B.n267 73.8041
R802 B.n481 B.n267 73.8041
R803 B.n481 B.n263 73.8041
R804 B.n487 B.n263 73.8041
R805 B.n487 B.n259 73.8041
R806 B.n493 B.n259 73.8041
R807 B.n493 B.n255 73.8041
R808 B.n499 B.n255 73.8041
R809 B.n499 B.n251 73.8041
R810 B.n505 B.n251 73.8041
R811 B.n511 B.n247 73.8041
R812 B.n511 B.n243 73.8041
R813 B.n517 B.n243 73.8041
R814 B.n517 B.n239 73.8041
R815 B.n523 B.n239 73.8041
R816 B.n523 B.n235 73.8041
R817 B.n529 B.n235 73.8041
R818 B.n529 B.n231 73.8041
R819 B.n535 B.n231 73.8041
R820 B.n535 B.n227 73.8041
R821 B.n541 B.n227 73.8041
R822 B.n547 B.n223 73.8041
R823 B.n547 B.n219 73.8041
R824 B.n554 B.n219 73.8041
R825 B.n554 B.n215 73.8041
R826 B.n560 B.n215 73.8041
R827 B.n560 B.n4 73.8041
R828 B.n714 B.n4 73.8041
R829 B.n714 B.n713 73.8041
R830 B.n713 B.n712 73.8041
R831 B.n712 B.n8 73.8041
R832 B.n12 B.n8 73.8041
R833 B.n705 B.n12 73.8041
R834 B.n705 B.n704 73.8041
R835 B.n704 B.n703 73.8041
R836 B.n703 B.n16 73.8041
R837 B.n697 B.n696 73.8041
R838 B.n696 B.n695 73.8041
R839 B.n695 B.n23 73.8041
R840 B.n689 B.n23 73.8041
R841 B.n689 B.n688 73.8041
R842 B.n688 B.n687 73.8041
R843 B.n687 B.n30 73.8041
R844 B.n681 B.n30 73.8041
R845 B.n681 B.n680 73.8041
R846 B.n680 B.n679 73.8041
R847 B.n679 B.n37 73.8041
R848 B.n673 B.n672 73.8041
R849 B.n672 B.n671 73.8041
R850 B.n671 B.n44 73.8041
R851 B.n665 B.n44 73.8041
R852 B.n665 B.n664 73.8041
R853 B.n664 B.n663 73.8041
R854 B.n663 B.n51 73.8041
R855 B.n657 B.n51 73.8041
R856 B.n657 B.n656 73.8041
R857 B.n656 B.n655 73.8041
R858 B.n655 B.n58 73.8041
R859 B.n649 B.n58 73.8041
R860 B.n649 B.n648 73.8041
R861 B.n648 B.n647 73.8041
R862 B.n641 B.n68 73.8041
R863 B.n641 B.n640 73.8041
R864 B.n640 B.n639 73.8041
R865 B.n639 B.n72 73.8041
R866 B.n633 B.n72 73.8041
R867 B.n633 B.n632 73.8041
R868 B.n632 B.n631 73.8041
R869 B.n631 B.n79 73.8041
R870 B.n625 B.n79 73.8041
R871 B.n111 B.t7 72.2414
R872 B.n311 B.t16 72.2414
R873 B.n114 B.t10 72.2365
R874 B.n317 B.t13 72.2365
R875 B.n84 B.n82 71.676
R876 B.n117 B.n85 71.676
R877 B.n121 B.n86 71.676
R878 B.n125 B.n87 71.676
R879 B.n129 B.n88 71.676
R880 B.n133 B.n89 71.676
R881 B.n137 B.n90 71.676
R882 B.n141 B.n91 71.676
R883 B.n145 B.n92 71.676
R884 B.n149 B.n93 71.676
R885 B.n153 B.n94 71.676
R886 B.n158 B.n95 71.676
R887 B.n162 B.n96 71.676
R888 B.n166 B.n97 71.676
R889 B.n170 B.n98 71.676
R890 B.n174 B.n99 71.676
R891 B.n178 B.n100 71.676
R892 B.n182 B.n101 71.676
R893 B.n186 B.n102 71.676
R894 B.n190 B.n103 71.676
R895 B.n194 B.n104 71.676
R896 B.n198 B.n105 71.676
R897 B.n202 B.n106 71.676
R898 B.n206 B.n107 71.676
R899 B.n210 B.n108 71.676
R900 B.n109 B.n108 71.676
R901 B.n209 B.n107 71.676
R902 B.n205 B.n106 71.676
R903 B.n201 B.n105 71.676
R904 B.n197 B.n104 71.676
R905 B.n193 B.n103 71.676
R906 B.n189 B.n102 71.676
R907 B.n185 B.n101 71.676
R908 B.n181 B.n100 71.676
R909 B.n177 B.n99 71.676
R910 B.n173 B.n98 71.676
R911 B.n169 B.n97 71.676
R912 B.n165 B.n96 71.676
R913 B.n161 B.n95 71.676
R914 B.n157 B.n94 71.676
R915 B.n152 B.n93 71.676
R916 B.n148 B.n92 71.676
R917 B.n144 B.n91 71.676
R918 B.n140 B.n90 71.676
R919 B.n136 B.n89 71.676
R920 B.n132 B.n88 71.676
R921 B.n128 B.n87 71.676
R922 B.n124 B.n86 71.676
R923 B.n120 B.n85 71.676
R924 B.n116 B.n84 71.676
R925 B.n329 B.n297 71.676
R926 B.n335 B.n334 71.676
R927 B.n338 B.n337 71.676
R928 B.n343 B.n342 71.676
R929 B.n346 B.n345 71.676
R930 B.n351 B.n350 71.676
R931 B.n354 B.n353 71.676
R932 B.n359 B.n358 71.676
R933 B.n362 B.n361 71.676
R934 B.n367 B.n366 71.676
R935 B.n370 B.n369 71.676
R936 B.n375 B.n374 71.676
R937 B.n378 B.n377 71.676
R938 B.n383 B.n382 71.676
R939 B.n386 B.n385 71.676
R940 B.n392 B.n391 71.676
R941 B.n395 B.n394 71.676
R942 B.n400 B.n399 71.676
R943 B.n403 B.n402 71.676
R944 B.n408 B.n407 71.676
R945 B.n411 B.n410 71.676
R946 B.n416 B.n415 71.676
R947 B.n419 B.n418 71.676
R948 B.n424 B.n423 71.676
R949 B.n427 B.n426 71.676
R950 B.n330 B.n329 71.676
R951 B.n336 B.n335 71.676
R952 B.n337 B.n326 71.676
R953 B.n344 B.n343 71.676
R954 B.n345 B.n324 71.676
R955 B.n352 B.n351 71.676
R956 B.n353 B.n322 71.676
R957 B.n360 B.n359 71.676
R958 B.n361 B.n320 71.676
R959 B.n368 B.n367 71.676
R960 B.n369 B.n315 71.676
R961 B.n376 B.n375 71.676
R962 B.n377 B.n313 71.676
R963 B.n384 B.n383 71.676
R964 B.n385 B.n309 71.676
R965 B.n393 B.n392 71.676
R966 B.n394 B.n307 71.676
R967 B.n401 B.n400 71.676
R968 B.n402 B.n305 71.676
R969 B.n409 B.n408 71.676
R970 B.n410 B.n303 71.676
R971 B.n417 B.n416 71.676
R972 B.n418 B.n301 71.676
R973 B.n425 B.n424 71.676
R974 B.n426 B.n299 71.676
R975 B.n716 B.n715 71.676
R976 B.n716 B.n2 71.676
R977 B.n541 B.t2 64.036
R978 B.n697 B.t3 64.036
R979 B.n505 B.t1 59.6946
R980 B.n673 B.t0 59.6946
R981 B.n155 B.n114 59.5399
R982 B.n112 B.n111 59.5399
R983 B.n388 B.n311 59.5399
R984 B.n318 B.n317 59.5399
R985 B.n456 B.t12 40.1584
R986 B.n68 B.t5 40.1584
R987 B.n463 B.t12 33.6463
R988 B.n647 B.t5 33.6463
R989 B.n434 B.n296 29.1907
R990 B.n430 B.n429 29.1907
R991 B.n627 B.n81 29.1907
R992 B.n622 B.n621 29.1907
R993 B B.n717 18.0485
R994 B.t1 B.n247 14.11
R995 B.t0 B.n37 14.11
R996 B.n435 B.n434 10.6151
R997 B.n436 B.n435 10.6151
R998 B.n436 B.n288 10.6151
R999 B.n446 B.n288 10.6151
R1000 B.n447 B.n446 10.6151
R1001 B.n448 B.n447 10.6151
R1002 B.n448 B.n280 10.6151
R1003 B.n459 B.n280 10.6151
R1004 B.n460 B.n459 10.6151
R1005 B.n461 B.n460 10.6151
R1006 B.n461 B.n273 10.6151
R1007 B.n471 B.n273 10.6151
R1008 B.n472 B.n471 10.6151
R1009 B.n473 B.n472 10.6151
R1010 B.n473 B.n265 10.6151
R1011 B.n483 B.n265 10.6151
R1012 B.n484 B.n483 10.6151
R1013 B.n485 B.n484 10.6151
R1014 B.n485 B.n257 10.6151
R1015 B.n495 B.n257 10.6151
R1016 B.n496 B.n495 10.6151
R1017 B.n497 B.n496 10.6151
R1018 B.n497 B.n249 10.6151
R1019 B.n507 B.n249 10.6151
R1020 B.n508 B.n507 10.6151
R1021 B.n509 B.n508 10.6151
R1022 B.n509 B.n241 10.6151
R1023 B.n519 B.n241 10.6151
R1024 B.n520 B.n519 10.6151
R1025 B.n521 B.n520 10.6151
R1026 B.n521 B.n233 10.6151
R1027 B.n531 B.n233 10.6151
R1028 B.n532 B.n531 10.6151
R1029 B.n533 B.n532 10.6151
R1030 B.n533 B.n225 10.6151
R1031 B.n543 B.n225 10.6151
R1032 B.n544 B.n543 10.6151
R1033 B.n545 B.n544 10.6151
R1034 B.n545 B.n217 10.6151
R1035 B.n556 B.n217 10.6151
R1036 B.n557 B.n556 10.6151
R1037 B.n558 B.n557 10.6151
R1038 B.n558 B.n0 10.6151
R1039 B.n331 B.n296 10.6151
R1040 B.n332 B.n331 10.6151
R1041 B.n333 B.n332 10.6151
R1042 B.n333 B.n327 10.6151
R1043 B.n339 B.n327 10.6151
R1044 B.n340 B.n339 10.6151
R1045 B.n341 B.n340 10.6151
R1046 B.n341 B.n325 10.6151
R1047 B.n347 B.n325 10.6151
R1048 B.n348 B.n347 10.6151
R1049 B.n349 B.n348 10.6151
R1050 B.n349 B.n323 10.6151
R1051 B.n355 B.n323 10.6151
R1052 B.n356 B.n355 10.6151
R1053 B.n357 B.n356 10.6151
R1054 B.n357 B.n321 10.6151
R1055 B.n363 B.n321 10.6151
R1056 B.n364 B.n363 10.6151
R1057 B.n365 B.n364 10.6151
R1058 B.n365 B.n319 10.6151
R1059 B.n372 B.n371 10.6151
R1060 B.n373 B.n372 10.6151
R1061 B.n373 B.n314 10.6151
R1062 B.n379 B.n314 10.6151
R1063 B.n380 B.n379 10.6151
R1064 B.n381 B.n380 10.6151
R1065 B.n381 B.n312 10.6151
R1066 B.n387 B.n312 10.6151
R1067 B.n390 B.n389 10.6151
R1068 B.n390 B.n308 10.6151
R1069 B.n396 B.n308 10.6151
R1070 B.n397 B.n396 10.6151
R1071 B.n398 B.n397 10.6151
R1072 B.n398 B.n306 10.6151
R1073 B.n404 B.n306 10.6151
R1074 B.n405 B.n404 10.6151
R1075 B.n406 B.n405 10.6151
R1076 B.n406 B.n304 10.6151
R1077 B.n412 B.n304 10.6151
R1078 B.n413 B.n412 10.6151
R1079 B.n414 B.n413 10.6151
R1080 B.n414 B.n302 10.6151
R1081 B.n420 B.n302 10.6151
R1082 B.n421 B.n420 10.6151
R1083 B.n422 B.n421 10.6151
R1084 B.n422 B.n300 10.6151
R1085 B.n428 B.n300 10.6151
R1086 B.n429 B.n428 10.6151
R1087 B.n430 B.n292 10.6151
R1088 B.n440 B.n292 10.6151
R1089 B.n441 B.n440 10.6151
R1090 B.n442 B.n441 10.6151
R1091 B.n442 B.n284 10.6151
R1092 B.n452 B.n284 10.6151
R1093 B.n453 B.n452 10.6151
R1094 B.n454 B.n453 10.6151
R1095 B.n454 B.n277 10.6151
R1096 B.n465 B.n277 10.6151
R1097 B.n466 B.n465 10.6151
R1098 B.n467 B.n466 10.6151
R1099 B.n467 B.n269 10.6151
R1100 B.n477 B.n269 10.6151
R1101 B.n478 B.n477 10.6151
R1102 B.n479 B.n478 10.6151
R1103 B.n479 B.n261 10.6151
R1104 B.n489 B.n261 10.6151
R1105 B.n490 B.n489 10.6151
R1106 B.n491 B.n490 10.6151
R1107 B.n491 B.n253 10.6151
R1108 B.n501 B.n253 10.6151
R1109 B.n502 B.n501 10.6151
R1110 B.n503 B.n502 10.6151
R1111 B.n503 B.n245 10.6151
R1112 B.n513 B.n245 10.6151
R1113 B.n514 B.n513 10.6151
R1114 B.n515 B.n514 10.6151
R1115 B.n515 B.n237 10.6151
R1116 B.n525 B.n237 10.6151
R1117 B.n526 B.n525 10.6151
R1118 B.n527 B.n526 10.6151
R1119 B.n527 B.n229 10.6151
R1120 B.n537 B.n229 10.6151
R1121 B.n538 B.n537 10.6151
R1122 B.n539 B.n538 10.6151
R1123 B.n539 B.n221 10.6151
R1124 B.n549 B.n221 10.6151
R1125 B.n550 B.n549 10.6151
R1126 B.n552 B.n550 10.6151
R1127 B.n552 B.n551 10.6151
R1128 B.n551 B.n213 10.6151
R1129 B.n563 B.n213 10.6151
R1130 B.n564 B.n563 10.6151
R1131 B.n565 B.n564 10.6151
R1132 B.n566 B.n565 10.6151
R1133 B.n567 B.n566 10.6151
R1134 B.n570 B.n567 10.6151
R1135 B.n571 B.n570 10.6151
R1136 B.n572 B.n571 10.6151
R1137 B.n573 B.n572 10.6151
R1138 B.n575 B.n573 10.6151
R1139 B.n576 B.n575 10.6151
R1140 B.n577 B.n576 10.6151
R1141 B.n578 B.n577 10.6151
R1142 B.n580 B.n578 10.6151
R1143 B.n581 B.n580 10.6151
R1144 B.n582 B.n581 10.6151
R1145 B.n583 B.n582 10.6151
R1146 B.n585 B.n583 10.6151
R1147 B.n586 B.n585 10.6151
R1148 B.n587 B.n586 10.6151
R1149 B.n588 B.n587 10.6151
R1150 B.n590 B.n588 10.6151
R1151 B.n591 B.n590 10.6151
R1152 B.n592 B.n591 10.6151
R1153 B.n593 B.n592 10.6151
R1154 B.n595 B.n593 10.6151
R1155 B.n596 B.n595 10.6151
R1156 B.n597 B.n596 10.6151
R1157 B.n598 B.n597 10.6151
R1158 B.n600 B.n598 10.6151
R1159 B.n601 B.n600 10.6151
R1160 B.n602 B.n601 10.6151
R1161 B.n603 B.n602 10.6151
R1162 B.n605 B.n603 10.6151
R1163 B.n606 B.n605 10.6151
R1164 B.n607 B.n606 10.6151
R1165 B.n608 B.n607 10.6151
R1166 B.n610 B.n608 10.6151
R1167 B.n611 B.n610 10.6151
R1168 B.n612 B.n611 10.6151
R1169 B.n613 B.n612 10.6151
R1170 B.n615 B.n613 10.6151
R1171 B.n616 B.n615 10.6151
R1172 B.n617 B.n616 10.6151
R1173 B.n618 B.n617 10.6151
R1174 B.n620 B.n618 10.6151
R1175 B.n621 B.n620 10.6151
R1176 B.n709 B.n1 10.6151
R1177 B.n709 B.n708 10.6151
R1178 B.n708 B.n707 10.6151
R1179 B.n707 B.n10 10.6151
R1180 B.n701 B.n10 10.6151
R1181 B.n701 B.n700 10.6151
R1182 B.n700 B.n699 10.6151
R1183 B.n699 B.n18 10.6151
R1184 B.n693 B.n18 10.6151
R1185 B.n693 B.n692 10.6151
R1186 B.n692 B.n691 10.6151
R1187 B.n691 B.n25 10.6151
R1188 B.n685 B.n25 10.6151
R1189 B.n685 B.n684 10.6151
R1190 B.n684 B.n683 10.6151
R1191 B.n683 B.n32 10.6151
R1192 B.n677 B.n32 10.6151
R1193 B.n677 B.n676 10.6151
R1194 B.n676 B.n675 10.6151
R1195 B.n675 B.n39 10.6151
R1196 B.n669 B.n39 10.6151
R1197 B.n669 B.n668 10.6151
R1198 B.n668 B.n667 10.6151
R1199 B.n667 B.n46 10.6151
R1200 B.n661 B.n46 10.6151
R1201 B.n661 B.n660 10.6151
R1202 B.n660 B.n659 10.6151
R1203 B.n659 B.n53 10.6151
R1204 B.n653 B.n53 10.6151
R1205 B.n653 B.n652 10.6151
R1206 B.n652 B.n651 10.6151
R1207 B.n651 B.n60 10.6151
R1208 B.n645 B.n60 10.6151
R1209 B.n645 B.n644 10.6151
R1210 B.n644 B.n643 10.6151
R1211 B.n643 B.n66 10.6151
R1212 B.n637 B.n66 10.6151
R1213 B.n637 B.n636 10.6151
R1214 B.n636 B.n635 10.6151
R1215 B.n635 B.n74 10.6151
R1216 B.n629 B.n74 10.6151
R1217 B.n629 B.n628 10.6151
R1218 B.n628 B.n627 10.6151
R1219 B.n115 B.n81 10.6151
R1220 B.n118 B.n115 10.6151
R1221 B.n119 B.n118 10.6151
R1222 B.n122 B.n119 10.6151
R1223 B.n123 B.n122 10.6151
R1224 B.n126 B.n123 10.6151
R1225 B.n127 B.n126 10.6151
R1226 B.n130 B.n127 10.6151
R1227 B.n131 B.n130 10.6151
R1228 B.n134 B.n131 10.6151
R1229 B.n135 B.n134 10.6151
R1230 B.n138 B.n135 10.6151
R1231 B.n139 B.n138 10.6151
R1232 B.n142 B.n139 10.6151
R1233 B.n143 B.n142 10.6151
R1234 B.n146 B.n143 10.6151
R1235 B.n147 B.n146 10.6151
R1236 B.n150 B.n147 10.6151
R1237 B.n151 B.n150 10.6151
R1238 B.n154 B.n151 10.6151
R1239 B.n159 B.n156 10.6151
R1240 B.n160 B.n159 10.6151
R1241 B.n163 B.n160 10.6151
R1242 B.n164 B.n163 10.6151
R1243 B.n167 B.n164 10.6151
R1244 B.n168 B.n167 10.6151
R1245 B.n171 B.n168 10.6151
R1246 B.n172 B.n171 10.6151
R1247 B.n176 B.n175 10.6151
R1248 B.n179 B.n176 10.6151
R1249 B.n180 B.n179 10.6151
R1250 B.n183 B.n180 10.6151
R1251 B.n184 B.n183 10.6151
R1252 B.n187 B.n184 10.6151
R1253 B.n188 B.n187 10.6151
R1254 B.n191 B.n188 10.6151
R1255 B.n192 B.n191 10.6151
R1256 B.n195 B.n192 10.6151
R1257 B.n196 B.n195 10.6151
R1258 B.n199 B.n196 10.6151
R1259 B.n200 B.n199 10.6151
R1260 B.n203 B.n200 10.6151
R1261 B.n204 B.n203 10.6151
R1262 B.n207 B.n204 10.6151
R1263 B.n208 B.n207 10.6151
R1264 B.n211 B.n208 10.6151
R1265 B.n212 B.n211 10.6151
R1266 B.n622 B.n212 10.6151
R1267 B.t2 B.n223 9.76863
R1268 B.t3 B.n16 9.76863
R1269 B.n717 B.n0 8.11757
R1270 B.n717 B.n1 8.11757
R1271 B.n371 B.n318 6.5566
R1272 B.n388 B.n387 6.5566
R1273 B.n156 B.n155 6.5566
R1274 B.n172 B.n112 6.5566
R1275 B.n319 B.n318 4.05904
R1276 B.n389 B.n388 4.05904
R1277 B.n155 B.n154 4.05904
R1278 B.n175 B.n112 4.05904
R1279 VP.n21 VP.n20 161.3
R1280 VP.n19 VP.n1 161.3
R1281 VP.n18 VP.n17 161.3
R1282 VP.n16 VP.n2 161.3
R1283 VP.n15 VP.n14 161.3
R1284 VP.n13 VP.n3 161.3
R1285 VP.n12 VP.n11 161.3
R1286 VP.n10 VP.n4 161.3
R1287 VP.n9 VP.n8 161.3
R1288 VP.n7 VP.n6 87.7864
R1289 VP.n22 VP.n0 87.7864
R1290 VP.n5 VP.t3 64.8928
R1291 VP.n5 VP.t0 63.5492
R1292 VP.n6 VP.n5 46.3946
R1293 VP.n14 VP.n13 40.577
R1294 VP.n14 VP.n2 40.577
R1295 VP.n7 VP.t1 31.0684
R1296 VP.n0 VP.t2 31.0684
R1297 VP.n8 VP.n4 24.5923
R1298 VP.n12 VP.n4 24.5923
R1299 VP.n13 VP.n12 24.5923
R1300 VP.n18 VP.n2 24.5923
R1301 VP.n19 VP.n18 24.5923
R1302 VP.n20 VP.n19 24.5923
R1303 VP.n8 VP.n7 2.45968
R1304 VP.n20 VP.n0 2.45968
R1305 VP.n9 VP.n6 0.354861
R1306 VP.n22 VP.n21 0.354861
R1307 VP VP.n22 0.267071
R1308 VP.n10 VP.n9 0.189894
R1309 VP.n11 VP.n10 0.189894
R1310 VP.n11 VP.n3 0.189894
R1311 VP.n15 VP.n3 0.189894
R1312 VP.n16 VP.n15 0.189894
R1313 VP.n17 VP.n16 0.189894
R1314 VP.n17 VP.n1 0.189894
R1315 VP.n21 VP.n1 0.189894
R1316 VDD1 VDD1.n1 107.436
R1317 VDD1 VDD1.n0 68.4615
R1318 VDD1.n0 VDD1.t0 4.07457
R1319 VDD1.n0 VDD1.t3 4.07457
R1320 VDD1.n1 VDD1.t2 4.07457
R1321 VDD1.n1 VDD1.t1 4.07457
C0 VDD2 VTAIL 4.30912f
C1 VN VP 5.70846f
C2 VDD1 VN 0.154064f
C3 VDD1 VP 2.55808f
C4 VN VTAIL 2.83384f
C5 VN VDD2 2.2405f
C6 VTAIL VP 2.84795f
C7 VDD2 VP 0.473188f
C8 VDD1 VTAIL 4.24706f
C9 VDD1 VDD2 1.30985f
C10 VDD2 B 3.876895f
C11 VDD1 B 7.86691f
C12 VTAIL B 6.027842f
C13 VN B 12.391621f
C14 VP B 10.754909f
C15 VDD1.t0 B 0.113136f
C16 VDD1.t3 B 0.113136f
C17 VDD1.n0 B 0.91791f
C18 VDD1.t2 B 0.113136f
C19 VDD1.t1 B 0.113136f
C20 VDD1.n1 B 1.44457f
C21 VP.t2 B 1.21746f
C22 VP.n0 B 0.552598f
C23 VP.n1 B 0.025456f
C24 VP.n2 B 0.050328f
C25 VP.n3 B 0.025456f
C26 VP.n4 B 0.047206f
C27 VP.t3 B 1.56512f
C28 VP.t0 B 1.55149f
C29 VP.n5 B 2.36971f
C30 VP.n6 B 1.32121f
C31 VP.t1 B 1.21746f
C32 VP.n7 B 0.552598f
C33 VP.n8 B 0.026232f
C34 VP.n9 B 0.041079f
C35 VP.n10 B 0.025456f
C36 VP.n11 B 0.025456f
C37 VP.n12 B 0.047206f
C38 VP.n13 B 0.050328f
C39 VP.n14 B 0.02056f
C40 VP.n15 B 0.025456f
C41 VP.n16 B 0.025456f
C42 VP.n17 B 0.025456f
C43 VP.n18 B 0.047206f
C44 VP.n19 B 0.047206f
C45 VP.n20 B 0.026232f
C46 VP.n21 B 0.041079f
C47 VP.n22 B 0.077989f
C48 VDD2.t0 B 0.109904f
C49 VDD2.t3 B 0.109904f
C50 VDD2.n0 B 1.37833f
C51 VDD2.t1 B 0.109904f
C52 VDD2.t2 B 0.109904f
C53 VDD2.n1 B 0.891197f
C54 VDD2.n2 B 3.45879f
C55 VTAIL.t4 B 0.809229f
C56 VTAIL.n0 B 0.422065f
C57 VTAIL.t2 B 0.809229f
C58 VTAIL.n1 B 0.544023f
C59 VTAIL.t1 B 0.809229f
C60 VTAIL.n2 B 1.36252f
C61 VTAIL.t6 B 0.809234f
C62 VTAIL.n3 B 1.36251f
C63 VTAIL.t5 B 0.809234f
C64 VTAIL.n4 B 0.544017f
C65 VTAIL.t3 B 0.809234f
C66 VTAIL.n5 B 0.544017f
C67 VTAIL.t0 B 0.809229f
C68 VTAIL.n6 B 1.36252f
C69 VTAIL.t7 B 0.809229f
C70 VTAIL.n7 B 1.23226f
C71 VN.t0 B 1.49078f
C72 VN.t3 B 1.50387f
C73 VN.n0 B 0.897091f
C74 VN.t2 B 1.49078f
C75 VN.t1 B 1.50387f
C76 VN.n1 B 2.2872f
.ends

