* NGSPICE file created from diff_pair_sample_0965.ext - technology: sky130A

.subckt diff_pair_sample_0965 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t1 VN.t0 VTAIL.t3 B.t0 sky130_fd_pr__nfet_01v8 ad=3.5841 pd=19.16 as=3.5841 ps=19.16 w=9.19 l=1.21
X1 VDD1.t1 VP.t0 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=3.5841 pd=19.16 as=3.5841 ps=19.16 w=9.19 l=1.21
X2 B.t15 B.t13 B.t14 B.t7 sky130_fd_pr__nfet_01v8 ad=3.5841 pd=19.16 as=0 ps=0 w=9.19 l=1.21
X3 VDD1.t0 VP.t1 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=3.5841 pd=19.16 as=3.5841 ps=19.16 w=9.19 l=1.21
X4 VDD2.t0 VN.t1 VTAIL.t2 B.t1 sky130_fd_pr__nfet_01v8 ad=3.5841 pd=19.16 as=3.5841 ps=19.16 w=9.19 l=1.21
X5 B.t12 B.t10 B.t11 B.t3 sky130_fd_pr__nfet_01v8 ad=3.5841 pd=19.16 as=0 ps=0 w=9.19 l=1.21
X6 B.t9 B.t6 B.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=3.5841 pd=19.16 as=0 ps=0 w=9.19 l=1.21
X7 B.t5 B.t2 B.t4 B.t3 sky130_fd_pr__nfet_01v8 ad=3.5841 pd=19.16 as=0 ps=0 w=9.19 l=1.21
R0 VN VN.t1 335.435
R1 VN VN.t0 296.454
R2 VTAIL.n194 VTAIL.n150 289.615
R3 VTAIL.n44 VTAIL.n0 289.615
R4 VTAIL.n144 VTAIL.n100 289.615
R5 VTAIL.n94 VTAIL.n50 289.615
R6 VTAIL.n167 VTAIL.n166 185
R7 VTAIL.n169 VTAIL.n168 185
R8 VTAIL.n162 VTAIL.n161 185
R9 VTAIL.n175 VTAIL.n174 185
R10 VTAIL.n177 VTAIL.n176 185
R11 VTAIL.n158 VTAIL.n157 185
R12 VTAIL.n184 VTAIL.n183 185
R13 VTAIL.n185 VTAIL.n156 185
R14 VTAIL.n187 VTAIL.n186 185
R15 VTAIL.n154 VTAIL.n153 185
R16 VTAIL.n193 VTAIL.n192 185
R17 VTAIL.n195 VTAIL.n194 185
R18 VTAIL.n17 VTAIL.n16 185
R19 VTAIL.n19 VTAIL.n18 185
R20 VTAIL.n12 VTAIL.n11 185
R21 VTAIL.n25 VTAIL.n24 185
R22 VTAIL.n27 VTAIL.n26 185
R23 VTAIL.n8 VTAIL.n7 185
R24 VTAIL.n34 VTAIL.n33 185
R25 VTAIL.n35 VTAIL.n6 185
R26 VTAIL.n37 VTAIL.n36 185
R27 VTAIL.n4 VTAIL.n3 185
R28 VTAIL.n43 VTAIL.n42 185
R29 VTAIL.n45 VTAIL.n44 185
R30 VTAIL.n145 VTAIL.n144 185
R31 VTAIL.n143 VTAIL.n142 185
R32 VTAIL.n104 VTAIL.n103 185
R33 VTAIL.n108 VTAIL.n106 185
R34 VTAIL.n137 VTAIL.n136 185
R35 VTAIL.n135 VTAIL.n134 185
R36 VTAIL.n110 VTAIL.n109 185
R37 VTAIL.n129 VTAIL.n128 185
R38 VTAIL.n127 VTAIL.n126 185
R39 VTAIL.n114 VTAIL.n113 185
R40 VTAIL.n121 VTAIL.n120 185
R41 VTAIL.n119 VTAIL.n118 185
R42 VTAIL.n95 VTAIL.n94 185
R43 VTAIL.n93 VTAIL.n92 185
R44 VTAIL.n54 VTAIL.n53 185
R45 VTAIL.n58 VTAIL.n56 185
R46 VTAIL.n87 VTAIL.n86 185
R47 VTAIL.n85 VTAIL.n84 185
R48 VTAIL.n60 VTAIL.n59 185
R49 VTAIL.n79 VTAIL.n78 185
R50 VTAIL.n77 VTAIL.n76 185
R51 VTAIL.n64 VTAIL.n63 185
R52 VTAIL.n71 VTAIL.n70 185
R53 VTAIL.n69 VTAIL.n68 185
R54 VTAIL.n165 VTAIL.t3 149.524
R55 VTAIL.n15 VTAIL.t1 149.524
R56 VTAIL.n117 VTAIL.t0 149.524
R57 VTAIL.n67 VTAIL.t2 149.524
R58 VTAIL.n168 VTAIL.n167 104.615
R59 VTAIL.n168 VTAIL.n161 104.615
R60 VTAIL.n175 VTAIL.n161 104.615
R61 VTAIL.n176 VTAIL.n175 104.615
R62 VTAIL.n176 VTAIL.n157 104.615
R63 VTAIL.n184 VTAIL.n157 104.615
R64 VTAIL.n185 VTAIL.n184 104.615
R65 VTAIL.n186 VTAIL.n185 104.615
R66 VTAIL.n186 VTAIL.n153 104.615
R67 VTAIL.n193 VTAIL.n153 104.615
R68 VTAIL.n194 VTAIL.n193 104.615
R69 VTAIL.n18 VTAIL.n17 104.615
R70 VTAIL.n18 VTAIL.n11 104.615
R71 VTAIL.n25 VTAIL.n11 104.615
R72 VTAIL.n26 VTAIL.n25 104.615
R73 VTAIL.n26 VTAIL.n7 104.615
R74 VTAIL.n34 VTAIL.n7 104.615
R75 VTAIL.n35 VTAIL.n34 104.615
R76 VTAIL.n36 VTAIL.n35 104.615
R77 VTAIL.n36 VTAIL.n3 104.615
R78 VTAIL.n43 VTAIL.n3 104.615
R79 VTAIL.n44 VTAIL.n43 104.615
R80 VTAIL.n144 VTAIL.n143 104.615
R81 VTAIL.n143 VTAIL.n103 104.615
R82 VTAIL.n108 VTAIL.n103 104.615
R83 VTAIL.n136 VTAIL.n108 104.615
R84 VTAIL.n136 VTAIL.n135 104.615
R85 VTAIL.n135 VTAIL.n109 104.615
R86 VTAIL.n128 VTAIL.n109 104.615
R87 VTAIL.n128 VTAIL.n127 104.615
R88 VTAIL.n127 VTAIL.n113 104.615
R89 VTAIL.n120 VTAIL.n113 104.615
R90 VTAIL.n120 VTAIL.n119 104.615
R91 VTAIL.n94 VTAIL.n93 104.615
R92 VTAIL.n93 VTAIL.n53 104.615
R93 VTAIL.n58 VTAIL.n53 104.615
R94 VTAIL.n86 VTAIL.n58 104.615
R95 VTAIL.n86 VTAIL.n85 104.615
R96 VTAIL.n85 VTAIL.n59 104.615
R97 VTAIL.n78 VTAIL.n59 104.615
R98 VTAIL.n78 VTAIL.n77 104.615
R99 VTAIL.n77 VTAIL.n63 104.615
R100 VTAIL.n70 VTAIL.n63 104.615
R101 VTAIL.n70 VTAIL.n69 104.615
R102 VTAIL.n167 VTAIL.t3 52.3082
R103 VTAIL.n17 VTAIL.t1 52.3082
R104 VTAIL.n119 VTAIL.t0 52.3082
R105 VTAIL.n69 VTAIL.t2 52.3082
R106 VTAIL.n199 VTAIL.n198 31.2157
R107 VTAIL.n49 VTAIL.n48 31.2157
R108 VTAIL.n149 VTAIL.n148 31.2157
R109 VTAIL.n99 VTAIL.n98 31.2157
R110 VTAIL.n99 VTAIL.n49 22.9445
R111 VTAIL.n199 VTAIL.n149 21.6169
R112 VTAIL.n187 VTAIL.n154 13.1884
R113 VTAIL.n37 VTAIL.n4 13.1884
R114 VTAIL.n106 VTAIL.n104 13.1884
R115 VTAIL.n56 VTAIL.n54 13.1884
R116 VTAIL.n188 VTAIL.n156 12.8005
R117 VTAIL.n192 VTAIL.n191 12.8005
R118 VTAIL.n38 VTAIL.n6 12.8005
R119 VTAIL.n42 VTAIL.n41 12.8005
R120 VTAIL.n142 VTAIL.n141 12.8005
R121 VTAIL.n138 VTAIL.n137 12.8005
R122 VTAIL.n92 VTAIL.n91 12.8005
R123 VTAIL.n88 VTAIL.n87 12.8005
R124 VTAIL.n183 VTAIL.n182 12.0247
R125 VTAIL.n195 VTAIL.n152 12.0247
R126 VTAIL.n33 VTAIL.n32 12.0247
R127 VTAIL.n45 VTAIL.n2 12.0247
R128 VTAIL.n145 VTAIL.n102 12.0247
R129 VTAIL.n134 VTAIL.n107 12.0247
R130 VTAIL.n95 VTAIL.n52 12.0247
R131 VTAIL.n84 VTAIL.n57 12.0247
R132 VTAIL.n181 VTAIL.n158 11.249
R133 VTAIL.n196 VTAIL.n150 11.249
R134 VTAIL.n31 VTAIL.n8 11.249
R135 VTAIL.n46 VTAIL.n0 11.249
R136 VTAIL.n146 VTAIL.n100 11.249
R137 VTAIL.n133 VTAIL.n110 11.249
R138 VTAIL.n96 VTAIL.n50 11.249
R139 VTAIL.n83 VTAIL.n60 11.249
R140 VTAIL.n178 VTAIL.n177 10.4732
R141 VTAIL.n28 VTAIL.n27 10.4732
R142 VTAIL.n130 VTAIL.n129 10.4732
R143 VTAIL.n80 VTAIL.n79 10.4732
R144 VTAIL.n166 VTAIL.n165 10.2747
R145 VTAIL.n16 VTAIL.n15 10.2747
R146 VTAIL.n118 VTAIL.n117 10.2747
R147 VTAIL.n68 VTAIL.n67 10.2747
R148 VTAIL.n174 VTAIL.n160 9.69747
R149 VTAIL.n24 VTAIL.n10 9.69747
R150 VTAIL.n126 VTAIL.n112 9.69747
R151 VTAIL.n76 VTAIL.n62 9.69747
R152 VTAIL.n198 VTAIL.n197 9.45567
R153 VTAIL.n48 VTAIL.n47 9.45567
R154 VTAIL.n148 VTAIL.n147 9.45567
R155 VTAIL.n98 VTAIL.n97 9.45567
R156 VTAIL.n197 VTAIL.n196 9.3005
R157 VTAIL.n152 VTAIL.n151 9.3005
R158 VTAIL.n191 VTAIL.n190 9.3005
R159 VTAIL.n164 VTAIL.n163 9.3005
R160 VTAIL.n171 VTAIL.n170 9.3005
R161 VTAIL.n173 VTAIL.n172 9.3005
R162 VTAIL.n160 VTAIL.n159 9.3005
R163 VTAIL.n179 VTAIL.n178 9.3005
R164 VTAIL.n181 VTAIL.n180 9.3005
R165 VTAIL.n182 VTAIL.n155 9.3005
R166 VTAIL.n189 VTAIL.n188 9.3005
R167 VTAIL.n47 VTAIL.n46 9.3005
R168 VTAIL.n2 VTAIL.n1 9.3005
R169 VTAIL.n41 VTAIL.n40 9.3005
R170 VTAIL.n14 VTAIL.n13 9.3005
R171 VTAIL.n21 VTAIL.n20 9.3005
R172 VTAIL.n23 VTAIL.n22 9.3005
R173 VTAIL.n10 VTAIL.n9 9.3005
R174 VTAIL.n29 VTAIL.n28 9.3005
R175 VTAIL.n31 VTAIL.n30 9.3005
R176 VTAIL.n32 VTAIL.n5 9.3005
R177 VTAIL.n39 VTAIL.n38 9.3005
R178 VTAIL.n116 VTAIL.n115 9.3005
R179 VTAIL.n123 VTAIL.n122 9.3005
R180 VTAIL.n125 VTAIL.n124 9.3005
R181 VTAIL.n112 VTAIL.n111 9.3005
R182 VTAIL.n131 VTAIL.n130 9.3005
R183 VTAIL.n133 VTAIL.n132 9.3005
R184 VTAIL.n107 VTAIL.n105 9.3005
R185 VTAIL.n139 VTAIL.n138 9.3005
R186 VTAIL.n147 VTAIL.n146 9.3005
R187 VTAIL.n102 VTAIL.n101 9.3005
R188 VTAIL.n141 VTAIL.n140 9.3005
R189 VTAIL.n66 VTAIL.n65 9.3005
R190 VTAIL.n73 VTAIL.n72 9.3005
R191 VTAIL.n75 VTAIL.n74 9.3005
R192 VTAIL.n62 VTAIL.n61 9.3005
R193 VTAIL.n81 VTAIL.n80 9.3005
R194 VTAIL.n83 VTAIL.n82 9.3005
R195 VTAIL.n57 VTAIL.n55 9.3005
R196 VTAIL.n89 VTAIL.n88 9.3005
R197 VTAIL.n97 VTAIL.n96 9.3005
R198 VTAIL.n52 VTAIL.n51 9.3005
R199 VTAIL.n91 VTAIL.n90 9.3005
R200 VTAIL.n173 VTAIL.n162 8.92171
R201 VTAIL.n23 VTAIL.n12 8.92171
R202 VTAIL.n125 VTAIL.n114 8.92171
R203 VTAIL.n75 VTAIL.n64 8.92171
R204 VTAIL.n170 VTAIL.n169 8.14595
R205 VTAIL.n20 VTAIL.n19 8.14595
R206 VTAIL.n122 VTAIL.n121 8.14595
R207 VTAIL.n72 VTAIL.n71 8.14595
R208 VTAIL.n166 VTAIL.n164 7.3702
R209 VTAIL.n16 VTAIL.n14 7.3702
R210 VTAIL.n118 VTAIL.n116 7.3702
R211 VTAIL.n68 VTAIL.n66 7.3702
R212 VTAIL.n169 VTAIL.n164 5.81868
R213 VTAIL.n19 VTAIL.n14 5.81868
R214 VTAIL.n121 VTAIL.n116 5.81868
R215 VTAIL.n71 VTAIL.n66 5.81868
R216 VTAIL.n170 VTAIL.n162 5.04292
R217 VTAIL.n20 VTAIL.n12 5.04292
R218 VTAIL.n122 VTAIL.n114 5.04292
R219 VTAIL.n72 VTAIL.n64 5.04292
R220 VTAIL.n174 VTAIL.n173 4.26717
R221 VTAIL.n24 VTAIL.n23 4.26717
R222 VTAIL.n126 VTAIL.n125 4.26717
R223 VTAIL.n76 VTAIL.n75 4.26717
R224 VTAIL.n177 VTAIL.n160 3.49141
R225 VTAIL.n27 VTAIL.n10 3.49141
R226 VTAIL.n129 VTAIL.n112 3.49141
R227 VTAIL.n79 VTAIL.n62 3.49141
R228 VTAIL.n165 VTAIL.n163 2.84303
R229 VTAIL.n15 VTAIL.n13 2.84303
R230 VTAIL.n117 VTAIL.n115 2.84303
R231 VTAIL.n67 VTAIL.n65 2.84303
R232 VTAIL.n178 VTAIL.n158 2.71565
R233 VTAIL.n198 VTAIL.n150 2.71565
R234 VTAIL.n28 VTAIL.n8 2.71565
R235 VTAIL.n48 VTAIL.n0 2.71565
R236 VTAIL.n148 VTAIL.n100 2.71565
R237 VTAIL.n130 VTAIL.n110 2.71565
R238 VTAIL.n98 VTAIL.n50 2.71565
R239 VTAIL.n80 VTAIL.n60 2.71565
R240 VTAIL.n183 VTAIL.n181 1.93989
R241 VTAIL.n196 VTAIL.n195 1.93989
R242 VTAIL.n33 VTAIL.n31 1.93989
R243 VTAIL.n46 VTAIL.n45 1.93989
R244 VTAIL.n146 VTAIL.n145 1.93989
R245 VTAIL.n134 VTAIL.n133 1.93989
R246 VTAIL.n96 VTAIL.n95 1.93989
R247 VTAIL.n84 VTAIL.n83 1.93989
R248 VTAIL.n182 VTAIL.n156 1.16414
R249 VTAIL.n192 VTAIL.n152 1.16414
R250 VTAIL.n32 VTAIL.n6 1.16414
R251 VTAIL.n42 VTAIL.n2 1.16414
R252 VTAIL.n142 VTAIL.n102 1.16414
R253 VTAIL.n137 VTAIL.n107 1.16414
R254 VTAIL.n92 VTAIL.n52 1.16414
R255 VTAIL.n87 VTAIL.n57 1.16414
R256 VTAIL.n149 VTAIL.n99 1.13412
R257 VTAIL VTAIL.n49 0.860414
R258 VTAIL.n188 VTAIL.n187 0.388379
R259 VTAIL.n191 VTAIL.n154 0.388379
R260 VTAIL.n38 VTAIL.n37 0.388379
R261 VTAIL.n41 VTAIL.n4 0.388379
R262 VTAIL.n141 VTAIL.n104 0.388379
R263 VTAIL.n138 VTAIL.n106 0.388379
R264 VTAIL.n91 VTAIL.n54 0.388379
R265 VTAIL.n88 VTAIL.n56 0.388379
R266 VTAIL VTAIL.n199 0.274207
R267 VTAIL.n171 VTAIL.n163 0.155672
R268 VTAIL.n172 VTAIL.n171 0.155672
R269 VTAIL.n172 VTAIL.n159 0.155672
R270 VTAIL.n179 VTAIL.n159 0.155672
R271 VTAIL.n180 VTAIL.n179 0.155672
R272 VTAIL.n180 VTAIL.n155 0.155672
R273 VTAIL.n189 VTAIL.n155 0.155672
R274 VTAIL.n190 VTAIL.n189 0.155672
R275 VTAIL.n190 VTAIL.n151 0.155672
R276 VTAIL.n197 VTAIL.n151 0.155672
R277 VTAIL.n21 VTAIL.n13 0.155672
R278 VTAIL.n22 VTAIL.n21 0.155672
R279 VTAIL.n22 VTAIL.n9 0.155672
R280 VTAIL.n29 VTAIL.n9 0.155672
R281 VTAIL.n30 VTAIL.n29 0.155672
R282 VTAIL.n30 VTAIL.n5 0.155672
R283 VTAIL.n39 VTAIL.n5 0.155672
R284 VTAIL.n40 VTAIL.n39 0.155672
R285 VTAIL.n40 VTAIL.n1 0.155672
R286 VTAIL.n47 VTAIL.n1 0.155672
R287 VTAIL.n147 VTAIL.n101 0.155672
R288 VTAIL.n140 VTAIL.n101 0.155672
R289 VTAIL.n140 VTAIL.n139 0.155672
R290 VTAIL.n139 VTAIL.n105 0.155672
R291 VTAIL.n132 VTAIL.n105 0.155672
R292 VTAIL.n132 VTAIL.n131 0.155672
R293 VTAIL.n131 VTAIL.n111 0.155672
R294 VTAIL.n124 VTAIL.n111 0.155672
R295 VTAIL.n124 VTAIL.n123 0.155672
R296 VTAIL.n123 VTAIL.n115 0.155672
R297 VTAIL.n97 VTAIL.n51 0.155672
R298 VTAIL.n90 VTAIL.n51 0.155672
R299 VTAIL.n90 VTAIL.n89 0.155672
R300 VTAIL.n89 VTAIL.n55 0.155672
R301 VTAIL.n82 VTAIL.n55 0.155672
R302 VTAIL.n82 VTAIL.n81 0.155672
R303 VTAIL.n81 VTAIL.n61 0.155672
R304 VTAIL.n74 VTAIL.n61 0.155672
R305 VTAIL.n74 VTAIL.n73 0.155672
R306 VTAIL.n73 VTAIL.n65 0.155672
R307 VDD2.n93 VDD2.n49 289.615
R308 VDD2.n44 VDD2.n0 289.615
R309 VDD2.n94 VDD2.n93 185
R310 VDD2.n92 VDD2.n91 185
R311 VDD2.n53 VDD2.n52 185
R312 VDD2.n57 VDD2.n55 185
R313 VDD2.n86 VDD2.n85 185
R314 VDD2.n84 VDD2.n83 185
R315 VDD2.n59 VDD2.n58 185
R316 VDD2.n78 VDD2.n77 185
R317 VDD2.n76 VDD2.n75 185
R318 VDD2.n63 VDD2.n62 185
R319 VDD2.n70 VDD2.n69 185
R320 VDD2.n68 VDD2.n67 185
R321 VDD2.n17 VDD2.n16 185
R322 VDD2.n19 VDD2.n18 185
R323 VDD2.n12 VDD2.n11 185
R324 VDD2.n25 VDD2.n24 185
R325 VDD2.n27 VDD2.n26 185
R326 VDD2.n8 VDD2.n7 185
R327 VDD2.n34 VDD2.n33 185
R328 VDD2.n35 VDD2.n6 185
R329 VDD2.n37 VDD2.n36 185
R330 VDD2.n4 VDD2.n3 185
R331 VDD2.n43 VDD2.n42 185
R332 VDD2.n45 VDD2.n44 185
R333 VDD2.n66 VDD2.t0 149.524
R334 VDD2.n15 VDD2.t1 149.524
R335 VDD2.n93 VDD2.n92 104.615
R336 VDD2.n92 VDD2.n52 104.615
R337 VDD2.n57 VDD2.n52 104.615
R338 VDD2.n85 VDD2.n57 104.615
R339 VDD2.n85 VDD2.n84 104.615
R340 VDD2.n84 VDD2.n58 104.615
R341 VDD2.n77 VDD2.n58 104.615
R342 VDD2.n77 VDD2.n76 104.615
R343 VDD2.n76 VDD2.n62 104.615
R344 VDD2.n69 VDD2.n62 104.615
R345 VDD2.n69 VDD2.n68 104.615
R346 VDD2.n18 VDD2.n17 104.615
R347 VDD2.n18 VDD2.n11 104.615
R348 VDD2.n25 VDD2.n11 104.615
R349 VDD2.n26 VDD2.n25 104.615
R350 VDD2.n26 VDD2.n7 104.615
R351 VDD2.n34 VDD2.n7 104.615
R352 VDD2.n35 VDD2.n34 104.615
R353 VDD2.n36 VDD2.n35 104.615
R354 VDD2.n36 VDD2.n3 104.615
R355 VDD2.n43 VDD2.n3 104.615
R356 VDD2.n44 VDD2.n43 104.615
R357 VDD2.n98 VDD2.n48 82.1315
R358 VDD2.n68 VDD2.t0 52.3082
R359 VDD2.n17 VDD2.t1 52.3082
R360 VDD2.n98 VDD2.n97 47.8944
R361 VDD2.n55 VDD2.n53 13.1884
R362 VDD2.n37 VDD2.n4 13.1884
R363 VDD2.n91 VDD2.n90 12.8005
R364 VDD2.n87 VDD2.n86 12.8005
R365 VDD2.n38 VDD2.n6 12.8005
R366 VDD2.n42 VDD2.n41 12.8005
R367 VDD2.n94 VDD2.n51 12.0247
R368 VDD2.n83 VDD2.n56 12.0247
R369 VDD2.n33 VDD2.n32 12.0247
R370 VDD2.n45 VDD2.n2 12.0247
R371 VDD2.n95 VDD2.n49 11.249
R372 VDD2.n82 VDD2.n59 11.249
R373 VDD2.n31 VDD2.n8 11.249
R374 VDD2.n46 VDD2.n0 11.249
R375 VDD2.n79 VDD2.n78 10.4732
R376 VDD2.n28 VDD2.n27 10.4732
R377 VDD2.n67 VDD2.n66 10.2747
R378 VDD2.n16 VDD2.n15 10.2747
R379 VDD2.n75 VDD2.n61 9.69747
R380 VDD2.n24 VDD2.n10 9.69747
R381 VDD2.n97 VDD2.n96 9.45567
R382 VDD2.n48 VDD2.n47 9.45567
R383 VDD2.n65 VDD2.n64 9.3005
R384 VDD2.n72 VDD2.n71 9.3005
R385 VDD2.n74 VDD2.n73 9.3005
R386 VDD2.n61 VDD2.n60 9.3005
R387 VDD2.n80 VDD2.n79 9.3005
R388 VDD2.n82 VDD2.n81 9.3005
R389 VDD2.n56 VDD2.n54 9.3005
R390 VDD2.n88 VDD2.n87 9.3005
R391 VDD2.n96 VDD2.n95 9.3005
R392 VDD2.n51 VDD2.n50 9.3005
R393 VDD2.n90 VDD2.n89 9.3005
R394 VDD2.n47 VDD2.n46 9.3005
R395 VDD2.n2 VDD2.n1 9.3005
R396 VDD2.n41 VDD2.n40 9.3005
R397 VDD2.n14 VDD2.n13 9.3005
R398 VDD2.n21 VDD2.n20 9.3005
R399 VDD2.n23 VDD2.n22 9.3005
R400 VDD2.n10 VDD2.n9 9.3005
R401 VDD2.n29 VDD2.n28 9.3005
R402 VDD2.n31 VDD2.n30 9.3005
R403 VDD2.n32 VDD2.n5 9.3005
R404 VDD2.n39 VDD2.n38 9.3005
R405 VDD2.n74 VDD2.n63 8.92171
R406 VDD2.n23 VDD2.n12 8.92171
R407 VDD2.n71 VDD2.n70 8.14595
R408 VDD2.n20 VDD2.n19 8.14595
R409 VDD2.n67 VDD2.n65 7.3702
R410 VDD2.n16 VDD2.n14 7.3702
R411 VDD2.n70 VDD2.n65 5.81868
R412 VDD2.n19 VDD2.n14 5.81868
R413 VDD2.n71 VDD2.n63 5.04292
R414 VDD2.n20 VDD2.n12 5.04292
R415 VDD2.n75 VDD2.n74 4.26717
R416 VDD2.n24 VDD2.n23 4.26717
R417 VDD2.n78 VDD2.n61 3.49141
R418 VDD2.n27 VDD2.n10 3.49141
R419 VDD2.n66 VDD2.n64 2.84303
R420 VDD2.n15 VDD2.n13 2.84303
R421 VDD2.n97 VDD2.n49 2.71565
R422 VDD2.n79 VDD2.n59 2.71565
R423 VDD2.n28 VDD2.n8 2.71565
R424 VDD2.n48 VDD2.n0 2.71565
R425 VDD2.n95 VDD2.n94 1.93989
R426 VDD2.n83 VDD2.n82 1.93989
R427 VDD2.n33 VDD2.n31 1.93989
R428 VDD2.n46 VDD2.n45 1.93989
R429 VDD2.n91 VDD2.n51 1.16414
R430 VDD2.n86 VDD2.n56 1.16414
R431 VDD2.n32 VDD2.n6 1.16414
R432 VDD2.n42 VDD2.n2 1.16414
R433 VDD2 VDD2.n98 0.390586
R434 VDD2.n90 VDD2.n53 0.388379
R435 VDD2.n87 VDD2.n55 0.388379
R436 VDD2.n38 VDD2.n37 0.388379
R437 VDD2.n41 VDD2.n4 0.388379
R438 VDD2.n96 VDD2.n50 0.155672
R439 VDD2.n89 VDD2.n50 0.155672
R440 VDD2.n89 VDD2.n88 0.155672
R441 VDD2.n88 VDD2.n54 0.155672
R442 VDD2.n81 VDD2.n54 0.155672
R443 VDD2.n81 VDD2.n80 0.155672
R444 VDD2.n80 VDD2.n60 0.155672
R445 VDD2.n73 VDD2.n60 0.155672
R446 VDD2.n73 VDD2.n72 0.155672
R447 VDD2.n72 VDD2.n64 0.155672
R448 VDD2.n21 VDD2.n13 0.155672
R449 VDD2.n22 VDD2.n21 0.155672
R450 VDD2.n22 VDD2.n9 0.155672
R451 VDD2.n29 VDD2.n9 0.155672
R452 VDD2.n30 VDD2.n29 0.155672
R453 VDD2.n30 VDD2.n5 0.155672
R454 VDD2.n39 VDD2.n5 0.155672
R455 VDD2.n40 VDD2.n39 0.155672
R456 VDD2.n40 VDD2.n1 0.155672
R457 VDD2.n47 VDD2.n1 0.155672
R458 B.n529 B.n528 585
R459 B.n227 B.n72 585
R460 B.n226 B.n225 585
R461 B.n224 B.n223 585
R462 B.n222 B.n221 585
R463 B.n220 B.n219 585
R464 B.n218 B.n217 585
R465 B.n216 B.n215 585
R466 B.n214 B.n213 585
R467 B.n212 B.n211 585
R468 B.n210 B.n209 585
R469 B.n208 B.n207 585
R470 B.n206 B.n205 585
R471 B.n204 B.n203 585
R472 B.n202 B.n201 585
R473 B.n200 B.n199 585
R474 B.n198 B.n197 585
R475 B.n196 B.n195 585
R476 B.n194 B.n193 585
R477 B.n192 B.n191 585
R478 B.n190 B.n189 585
R479 B.n188 B.n187 585
R480 B.n186 B.n185 585
R481 B.n184 B.n183 585
R482 B.n182 B.n181 585
R483 B.n180 B.n179 585
R484 B.n178 B.n177 585
R485 B.n176 B.n175 585
R486 B.n174 B.n173 585
R487 B.n172 B.n171 585
R488 B.n170 B.n169 585
R489 B.n168 B.n167 585
R490 B.n166 B.n165 585
R491 B.n163 B.n162 585
R492 B.n161 B.n160 585
R493 B.n159 B.n158 585
R494 B.n157 B.n156 585
R495 B.n155 B.n154 585
R496 B.n153 B.n152 585
R497 B.n151 B.n150 585
R498 B.n149 B.n148 585
R499 B.n147 B.n146 585
R500 B.n145 B.n144 585
R501 B.n142 B.n141 585
R502 B.n140 B.n139 585
R503 B.n138 B.n137 585
R504 B.n136 B.n135 585
R505 B.n134 B.n133 585
R506 B.n132 B.n131 585
R507 B.n130 B.n129 585
R508 B.n128 B.n127 585
R509 B.n126 B.n125 585
R510 B.n124 B.n123 585
R511 B.n122 B.n121 585
R512 B.n120 B.n119 585
R513 B.n118 B.n117 585
R514 B.n116 B.n115 585
R515 B.n114 B.n113 585
R516 B.n112 B.n111 585
R517 B.n110 B.n109 585
R518 B.n108 B.n107 585
R519 B.n106 B.n105 585
R520 B.n104 B.n103 585
R521 B.n102 B.n101 585
R522 B.n100 B.n99 585
R523 B.n98 B.n97 585
R524 B.n96 B.n95 585
R525 B.n94 B.n93 585
R526 B.n92 B.n91 585
R527 B.n90 B.n89 585
R528 B.n88 B.n87 585
R529 B.n86 B.n85 585
R530 B.n84 B.n83 585
R531 B.n82 B.n81 585
R532 B.n80 B.n79 585
R533 B.n78 B.n77 585
R534 B.n527 B.n34 585
R535 B.n532 B.n34 585
R536 B.n526 B.n33 585
R537 B.n533 B.n33 585
R538 B.n525 B.n524 585
R539 B.n524 B.n29 585
R540 B.n523 B.n28 585
R541 B.n539 B.n28 585
R542 B.n522 B.n27 585
R543 B.n540 B.n27 585
R544 B.n521 B.n26 585
R545 B.n541 B.n26 585
R546 B.n520 B.n519 585
R547 B.n519 B.n22 585
R548 B.n518 B.n21 585
R549 B.n547 B.n21 585
R550 B.n517 B.n20 585
R551 B.n548 B.n20 585
R552 B.n516 B.n19 585
R553 B.n549 B.n19 585
R554 B.n515 B.n514 585
R555 B.n514 B.n15 585
R556 B.n513 B.n14 585
R557 B.n555 B.n14 585
R558 B.n512 B.n13 585
R559 B.n556 B.n13 585
R560 B.n511 B.n12 585
R561 B.n557 B.n12 585
R562 B.n510 B.n509 585
R563 B.n509 B.n8 585
R564 B.n508 B.n7 585
R565 B.n563 B.n7 585
R566 B.n507 B.n6 585
R567 B.n564 B.n6 585
R568 B.n506 B.n5 585
R569 B.n565 B.n5 585
R570 B.n505 B.n504 585
R571 B.n504 B.n4 585
R572 B.n503 B.n228 585
R573 B.n503 B.n502 585
R574 B.n493 B.n229 585
R575 B.n230 B.n229 585
R576 B.n495 B.n494 585
R577 B.n496 B.n495 585
R578 B.n492 B.n235 585
R579 B.n235 B.n234 585
R580 B.n491 B.n490 585
R581 B.n490 B.n489 585
R582 B.n237 B.n236 585
R583 B.n238 B.n237 585
R584 B.n482 B.n481 585
R585 B.n483 B.n482 585
R586 B.n480 B.n243 585
R587 B.n243 B.n242 585
R588 B.n479 B.n478 585
R589 B.n478 B.n477 585
R590 B.n245 B.n244 585
R591 B.n246 B.n245 585
R592 B.n470 B.n469 585
R593 B.n471 B.n470 585
R594 B.n468 B.n251 585
R595 B.n251 B.n250 585
R596 B.n467 B.n466 585
R597 B.n466 B.n465 585
R598 B.n253 B.n252 585
R599 B.n254 B.n253 585
R600 B.n458 B.n457 585
R601 B.n459 B.n458 585
R602 B.n456 B.n259 585
R603 B.n259 B.n258 585
R604 B.n451 B.n450 585
R605 B.n449 B.n299 585
R606 B.n448 B.n298 585
R607 B.n453 B.n298 585
R608 B.n447 B.n446 585
R609 B.n445 B.n444 585
R610 B.n443 B.n442 585
R611 B.n441 B.n440 585
R612 B.n439 B.n438 585
R613 B.n437 B.n436 585
R614 B.n435 B.n434 585
R615 B.n433 B.n432 585
R616 B.n431 B.n430 585
R617 B.n429 B.n428 585
R618 B.n427 B.n426 585
R619 B.n425 B.n424 585
R620 B.n423 B.n422 585
R621 B.n421 B.n420 585
R622 B.n419 B.n418 585
R623 B.n417 B.n416 585
R624 B.n415 B.n414 585
R625 B.n413 B.n412 585
R626 B.n411 B.n410 585
R627 B.n409 B.n408 585
R628 B.n407 B.n406 585
R629 B.n405 B.n404 585
R630 B.n403 B.n402 585
R631 B.n401 B.n400 585
R632 B.n399 B.n398 585
R633 B.n397 B.n396 585
R634 B.n395 B.n394 585
R635 B.n393 B.n392 585
R636 B.n391 B.n390 585
R637 B.n389 B.n388 585
R638 B.n387 B.n386 585
R639 B.n385 B.n384 585
R640 B.n383 B.n382 585
R641 B.n381 B.n380 585
R642 B.n379 B.n378 585
R643 B.n377 B.n376 585
R644 B.n375 B.n374 585
R645 B.n373 B.n372 585
R646 B.n371 B.n370 585
R647 B.n369 B.n368 585
R648 B.n367 B.n366 585
R649 B.n365 B.n364 585
R650 B.n363 B.n362 585
R651 B.n361 B.n360 585
R652 B.n359 B.n358 585
R653 B.n357 B.n356 585
R654 B.n355 B.n354 585
R655 B.n353 B.n352 585
R656 B.n351 B.n350 585
R657 B.n349 B.n348 585
R658 B.n347 B.n346 585
R659 B.n345 B.n344 585
R660 B.n343 B.n342 585
R661 B.n341 B.n340 585
R662 B.n339 B.n338 585
R663 B.n337 B.n336 585
R664 B.n335 B.n334 585
R665 B.n333 B.n332 585
R666 B.n331 B.n330 585
R667 B.n329 B.n328 585
R668 B.n327 B.n326 585
R669 B.n325 B.n324 585
R670 B.n323 B.n322 585
R671 B.n321 B.n320 585
R672 B.n319 B.n318 585
R673 B.n317 B.n316 585
R674 B.n315 B.n314 585
R675 B.n313 B.n312 585
R676 B.n311 B.n310 585
R677 B.n309 B.n308 585
R678 B.n307 B.n306 585
R679 B.n261 B.n260 585
R680 B.n455 B.n454 585
R681 B.n454 B.n453 585
R682 B.n257 B.n256 585
R683 B.n258 B.n257 585
R684 B.n461 B.n460 585
R685 B.n460 B.n459 585
R686 B.n462 B.n255 585
R687 B.n255 B.n254 585
R688 B.n464 B.n463 585
R689 B.n465 B.n464 585
R690 B.n249 B.n248 585
R691 B.n250 B.n249 585
R692 B.n473 B.n472 585
R693 B.n472 B.n471 585
R694 B.n474 B.n247 585
R695 B.n247 B.n246 585
R696 B.n476 B.n475 585
R697 B.n477 B.n476 585
R698 B.n241 B.n240 585
R699 B.n242 B.n241 585
R700 B.n485 B.n484 585
R701 B.n484 B.n483 585
R702 B.n486 B.n239 585
R703 B.n239 B.n238 585
R704 B.n488 B.n487 585
R705 B.n489 B.n488 585
R706 B.n233 B.n232 585
R707 B.n234 B.n233 585
R708 B.n498 B.n497 585
R709 B.n497 B.n496 585
R710 B.n499 B.n231 585
R711 B.n231 B.n230 585
R712 B.n501 B.n500 585
R713 B.n502 B.n501 585
R714 B.n2 B.n0 585
R715 B.n4 B.n2 585
R716 B.n3 B.n1 585
R717 B.n564 B.n3 585
R718 B.n562 B.n561 585
R719 B.n563 B.n562 585
R720 B.n560 B.n9 585
R721 B.n9 B.n8 585
R722 B.n559 B.n558 585
R723 B.n558 B.n557 585
R724 B.n11 B.n10 585
R725 B.n556 B.n11 585
R726 B.n554 B.n553 585
R727 B.n555 B.n554 585
R728 B.n552 B.n16 585
R729 B.n16 B.n15 585
R730 B.n551 B.n550 585
R731 B.n550 B.n549 585
R732 B.n18 B.n17 585
R733 B.n548 B.n18 585
R734 B.n546 B.n545 585
R735 B.n547 B.n546 585
R736 B.n544 B.n23 585
R737 B.n23 B.n22 585
R738 B.n543 B.n542 585
R739 B.n542 B.n541 585
R740 B.n25 B.n24 585
R741 B.n540 B.n25 585
R742 B.n538 B.n537 585
R743 B.n539 B.n538 585
R744 B.n536 B.n30 585
R745 B.n30 B.n29 585
R746 B.n535 B.n534 585
R747 B.n534 B.n533 585
R748 B.n32 B.n31 585
R749 B.n532 B.n32 585
R750 B.n567 B.n566 585
R751 B.n566 B.n565 585
R752 B.n451 B.n257 550.159
R753 B.n77 B.n32 550.159
R754 B.n454 B.n259 550.159
R755 B.n529 B.n34 550.159
R756 B.n303 B.t2 387.209
R757 B.n300 B.t10 387.209
R758 B.n75 B.t13 387.209
R759 B.n73 B.t6 387.209
R760 B.n303 B.t5 263.281
R761 B.n73 B.t8 263.281
R762 B.n300 B.t12 263.281
R763 B.n75 B.t14 263.281
R764 B.n531 B.n530 256.663
R765 B.n531 B.n71 256.663
R766 B.n531 B.n70 256.663
R767 B.n531 B.n69 256.663
R768 B.n531 B.n68 256.663
R769 B.n531 B.n67 256.663
R770 B.n531 B.n66 256.663
R771 B.n531 B.n65 256.663
R772 B.n531 B.n64 256.663
R773 B.n531 B.n63 256.663
R774 B.n531 B.n62 256.663
R775 B.n531 B.n61 256.663
R776 B.n531 B.n60 256.663
R777 B.n531 B.n59 256.663
R778 B.n531 B.n58 256.663
R779 B.n531 B.n57 256.663
R780 B.n531 B.n56 256.663
R781 B.n531 B.n55 256.663
R782 B.n531 B.n54 256.663
R783 B.n531 B.n53 256.663
R784 B.n531 B.n52 256.663
R785 B.n531 B.n51 256.663
R786 B.n531 B.n50 256.663
R787 B.n531 B.n49 256.663
R788 B.n531 B.n48 256.663
R789 B.n531 B.n47 256.663
R790 B.n531 B.n46 256.663
R791 B.n531 B.n45 256.663
R792 B.n531 B.n44 256.663
R793 B.n531 B.n43 256.663
R794 B.n531 B.n42 256.663
R795 B.n531 B.n41 256.663
R796 B.n531 B.n40 256.663
R797 B.n531 B.n39 256.663
R798 B.n531 B.n38 256.663
R799 B.n531 B.n37 256.663
R800 B.n531 B.n36 256.663
R801 B.n531 B.n35 256.663
R802 B.n453 B.n452 256.663
R803 B.n453 B.n262 256.663
R804 B.n453 B.n263 256.663
R805 B.n453 B.n264 256.663
R806 B.n453 B.n265 256.663
R807 B.n453 B.n266 256.663
R808 B.n453 B.n267 256.663
R809 B.n453 B.n268 256.663
R810 B.n453 B.n269 256.663
R811 B.n453 B.n270 256.663
R812 B.n453 B.n271 256.663
R813 B.n453 B.n272 256.663
R814 B.n453 B.n273 256.663
R815 B.n453 B.n274 256.663
R816 B.n453 B.n275 256.663
R817 B.n453 B.n276 256.663
R818 B.n453 B.n277 256.663
R819 B.n453 B.n278 256.663
R820 B.n453 B.n279 256.663
R821 B.n453 B.n280 256.663
R822 B.n453 B.n281 256.663
R823 B.n453 B.n282 256.663
R824 B.n453 B.n283 256.663
R825 B.n453 B.n284 256.663
R826 B.n453 B.n285 256.663
R827 B.n453 B.n286 256.663
R828 B.n453 B.n287 256.663
R829 B.n453 B.n288 256.663
R830 B.n453 B.n289 256.663
R831 B.n453 B.n290 256.663
R832 B.n453 B.n291 256.663
R833 B.n453 B.n292 256.663
R834 B.n453 B.n293 256.663
R835 B.n453 B.n294 256.663
R836 B.n453 B.n295 256.663
R837 B.n453 B.n296 256.663
R838 B.n453 B.n297 256.663
R839 B.n304 B.t4 233.415
R840 B.n74 B.t9 233.415
R841 B.n301 B.t11 233.415
R842 B.n76 B.t15 233.415
R843 B.n460 B.n257 163.367
R844 B.n460 B.n255 163.367
R845 B.n464 B.n255 163.367
R846 B.n464 B.n249 163.367
R847 B.n472 B.n249 163.367
R848 B.n472 B.n247 163.367
R849 B.n476 B.n247 163.367
R850 B.n476 B.n241 163.367
R851 B.n484 B.n241 163.367
R852 B.n484 B.n239 163.367
R853 B.n488 B.n239 163.367
R854 B.n488 B.n233 163.367
R855 B.n497 B.n233 163.367
R856 B.n497 B.n231 163.367
R857 B.n501 B.n231 163.367
R858 B.n501 B.n2 163.367
R859 B.n566 B.n2 163.367
R860 B.n566 B.n3 163.367
R861 B.n562 B.n3 163.367
R862 B.n562 B.n9 163.367
R863 B.n558 B.n9 163.367
R864 B.n558 B.n11 163.367
R865 B.n554 B.n11 163.367
R866 B.n554 B.n16 163.367
R867 B.n550 B.n16 163.367
R868 B.n550 B.n18 163.367
R869 B.n546 B.n18 163.367
R870 B.n546 B.n23 163.367
R871 B.n542 B.n23 163.367
R872 B.n542 B.n25 163.367
R873 B.n538 B.n25 163.367
R874 B.n538 B.n30 163.367
R875 B.n534 B.n30 163.367
R876 B.n534 B.n32 163.367
R877 B.n299 B.n298 163.367
R878 B.n446 B.n298 163.367
R879 B.n444 B.n443 163.367
R880 B.n440 B.n439 163.367
R881 B.n436 B.n435 163.367
R882 B.n432 B.n431 163.367
R883 B.n428 B.n427 163.367
R884 B.n424 B.n423 163.367
R885 B.n420 B.n419 163.367
R886 B.n416 B.n415 163.367
R887 B.n412 B.n411 163.367
R888 B.n408 B.n407 163.367
R889 B.n404 B.n403 163.367
R890 B.n400 B.n399 163.367
R891 B.n396 B.n395 163.367
R892 B.n392 B.n391 163.367
R893 B.n388 B.n387 163.367
R894 B.n384 B.n383 163.367
R895 B.n380 B.n379 163.367
R896 B.n376 B.n375 163.367
R897 B.n372 B.n371 163.367
R898 B.n368 B.n367 163.367
R899 B.n364 B.n363 163.367
R900 B.n360 B.n359 163.367
R901 B.n356 B.n355 163.367
R902 B.n352 B.n351 163.367
R903 B.n348 B.n347 163.367
R904 B.n344 B.n343 163.367
R905 B.n340 B.n339 163.367
R906 B.n336 B.n335 163.367
R907 B.n332 B.n331 163.367
R908 B.n328 B.n327 163.367
R909 B.n324 B.n323 163.367
R910 B.n320 B.n319 163.367
R911 B.n316 B.n315 163.367
R912 B.n312 B.n311 163.367
R913 B.n308 B.n307 163.367
R914 B.n454 B.n261 163.367
R915 B.n458 B.n259 163.367
R916 B.n458 B.n253 163.367
R917 B.n466 B.n253 163.367
R918 B.n466 B.n251 163.367
R919 B.n470 B.n251 163.367
R920 B.n470 B.n245 163.367
R921 B.n478 B.n245 163.367
R922 B.n478 B.n243 163.367
R923 B.n482 B.n243 163.367
R924 B.n482 B.n237 163.367
R925 B.n490 B.n237 163.367
R926 B.n490 B.n235 163.367
R927 B.n495 B.n235 163.367
R928 B.n495 B.n229 163.367
R929 B.n503 B.n229 163.367
R930 B.n504 B.n503 163.367
R931 B.n504 B.n5 163.367
R932 B.n6 B.n5 163.367
R933 B.n7 B.n6 163.367
R934 B.n509 B.n7 163.367
R935 B.n509 B.n12 163.367
R936 B.n13 B.n12 163.367
R937 B.n14 B.n13 163.367
R938 B.n514 B.n14 163.367
R939 B.n514 B.n19 163.367
R940 B.n20 B.n19 163.367
R941 B.n21 B.n20 163.367
R942 B.n519 B.n21 163.367
R943 B.n519 B.n26 163.367
R944 B.n27 B.n26 163.367
R945 B.n28 B.n27 163.367
R946 B.n524 B.n28 163.367
R947 B.n524 B.n33 163.367
R948 B.n34 B.n33 163.367
R949 B.n81 B.n80 163.367
R950 B.n85 B.n84 163.367
R951 B.n89 B.n88 163.367
R952 B.n93 B.n92 163.367
R953 B.n97 B.n96 163.367
R954 B.n101 B.n100 163.367
R955 B.n105 B.n104 163.367
R956 B.n109 B.n108 163.367
R957 B.n113 B.n112 163.367
R958 B.n117 B.n116 163.367
R959 B.n121 B.n120 163.367
R960 B.n125 B.n124 163.367
R961 B.n129 B.n128 163.367
R962 B.n133 B.n132 163.367
R963 B.n137 B.n136 163.367
R964 B.n141 B.n140 163.367
R965 B.n146 B.n145 163.367
R966 B.n150 B.n149 163.367
R967 B.n154 B.n153 163.367
R968 B.n158 B.n157 163.367
R969 B.n162 B.n161 163.367
R970 B.n167 B.n166 163.367
R971 B.n171 B.n170 163.367
R972 B.n175 B.n174 163.367
R973 B.n179 B.n178 163.367
R974 B.n183 B.n182 163.367
R975 B.n187 B.n186 163.367
R976 B.n191 B.n190 163.367
R977 B.n195 B.n194 163.367
R978 B.n199 B.n198 163.367
R979 B.n203 B.n202 163.367
R980 B.n207 B.n206 163.367
R981 B.n211 B.n210 163.367
R982 B.n215 B.n214 163.367
R983 B.n219 B.n218 163.367
R984 B.n223 B.n222 163.367
R985 B.n225 B.n72 163.367
R986 B.n453 B.n258 102.662
R987 B.n532 B.n531 102.662
R988 B.n452 B.n451 71.676
R989 B.n446 B.n262 71.676
R990 B.n443 B.n263 71.676
R991 B.n439 B.n264 71.676
R992 B.n435 B.n265 71.676
R993 B.n431 B.n266 71.676
R994 B.n427 B.n267 71.676
R995 B.n423 B.n268 71.676
R996 B.n419 B.n269 71.676
R997 B.n415 B.n270 71.676
R998 B.n411 B.n271 71.676
R999 B.n407 B.n272 71.676
R1000 B.n403 B.n273 71.676
R1001 B.n399 B.n274 71.676
R1002 B.n395 B.n275 71.676
R1003 B.n391 B.n276 71.676
R1004 B.n387 B.n277 71.676
R1005 B.n383 B.n278 71.676
R1006 B.n379 B.n279 71.676
R1007 B.n375 B.n280 71.676
R1008 B.n371 B.n281 71.676
R1009 B.n367 B.n282 71.676
R1010 B.n363 B.n283 71.676
R1011 B.n359 B.n284 71.676
R1012 B.n355 B.n285 71.676
R1013 B.n351 B.n286 71.676
R1014 B.n347 B.n287 71.676
R1015 B.n343 B.n288 71.676
R1016 B.n339 B.n289 71.676
R1017 B.n335 B.n290 71.676
R1018 B.n331 B.n291 71.676
R1019 B.n327 B.n292 71.676
R1020 B.n323 B.n293 71.676
R1021 B.n319 B.n294 71.676
R1022 B.n315 B.n295 71.676
R1023 B.n311 B.n296 71.676
R1024 B.n307 B.n297 71.676
R1025 B.n77 B.n35 71.676
R1026 B.n81 B.n36 71.676
R1027 B.n85 B.n37 71.676
R1028 B.n89 B.n38 71.676
R1029 B.n93 B.n39 71.676
R1030 B.n97 B.n40 71.676
R1031 B.n101 B.n41 71.676
R1032 B.n105 B.n42 71.676
R1033 B.n109 B.n43 71.676
R1034 B.n113 B.n44 71.676
R1035 B.n117 B.n45 71.676
R1036 B.n121 B.n46 71.676
R1037 B.n125 B.n47 71.676
R1038 B.n129 B.n48 71.676
R1039 B.n133 B.n49 71.676
R1040 B.n137 B.n50 71.676
R1041 B.n141 B.n51 71.676
R1042 B.n146 B.n52 71.676
R1043 B.n150 B.n53 71.676
R1044 B.n154 B.n54 71.676
R1045 B.n158 B.n55 71.676
R1046 B.n162 B.n56 71.676
R1047 B.n167 B.n57 71.676
R1048 B.n171 B.n58 71.676
R1049 B.n175 B.n59 71.676
R1050 B.n179 B.n60 71.676
R1051 B.n183 B.n61 71.676
R1052 B.n187 B.n62 71.676
R1053 B.n191 B.n63 71.676
R1054 B.n195 B.n64 71.676
R1055 B.n199 B.n65 71.676
R1056 B.n203 B.n66 71.676
R1057 B.n207 B.n67 71.676
R1058 B.n211 B.n68 71.676
R1059 B.n215 B.n69 71.676
R1060 B.n219 B.n70 71.676
R1061 B.n223 B.n71 71.676
R1062 B.n530 B.n72 71.676
R1063 B.n530 B.n529 71.676
R1064 B.n225 B.n71 71.676
R1065 B.n222 B.n70 71.676
R1066 B.n218 B.n69 71.676
R1067 B.n214 B.n68 71.676
R1068 B.n210 B.n67 71.676
R1069 B.n206 B.n66 71.676
R1070 B.n202 B.n65 71.676
R1071 B.n198 B.n64 71.676
R1072 B.n194 B.n63 71.676
R1073 B.n190 B.n62 71.676
R1074 B.n186 B.n61 71.676
R1075 B.n182 B.n60 71.676
R1076 B.n178 B.n59 71.676
R1077 B.n174 B.n58 71.676
R1078 B.n170 B.n57 71.676
R1079 B.n166 B.n56 71.676
R1080 B.n161 B.n55 71.676
R1081 B.n157 B.n54 71.676
R1082 B.n153 B.n53 71.676
R1083 B.n149 B.n52 71.676
R1084 B.n145 B.n51 71.676
R1085 B.n140 B.n50 71.676
R1086 B.n136 B.n49 71.676
R1087 B.n132 B.n48 71.676
R1088 B.n128 B.n47 71.676
R1089 B.n124 B.n46 71.676
R1090 B.n120 B.n45 71.676
R1091 B.n116 B.n44 71.676
R1092 B.n112 B.n43 71.676
R1093 B.n108 B.n42 71.676
R1094 B.n104 B.n41 71.676
R1095 B.n100 B.n40 71.676
R1096 B.n96 B.n39 71.676
R1097 B.n92 B.n38 71.676
R1098 B.n88 B.n37 71.676
R1099 B.n84 B.n36 71.676
R1100 B.n80 B.n35 71.676
R1101 B.n452 B.n299 71.676
R1102 B.n444 B.n262 71.676
R1103 B.n440 B.n263 71.676
R1104 B.n436 B.n264 71.676
R1105 B.n432 B.n265 71.676
R1106 B.n428 B.n266 71.676
R1107 B.n424 B.n267 71.676
R1108 B.n420 B.n268 71.676
R1109 B.n416 B.n269 71.676
R1110 B.n412 B.n270 71.676
R1111 B.n408 B.n271 71.676
R1112 B.n404 B.n272 71.676
R1113 B.n400 B.n273 71.676
R1114 B.n396 B.n274 71.676
R1115 B.n392 B.n275 71.676
R1116 B.n388 B.n276 71.676
R1117 B.n384 B.n277 71.676
R1118 B.n380 B.n278 71.676
R1119 B.n376 B.n279 71.676
R1120 B.n372 B.n280 71.676
R1121 B.n368 B.n281 71.676
R1122 B.n364 B.n282 71.676
R1123 B.n360 B.n283 71.676
R1124 B.n356 B.n284 71.676
R1125 B.n352 B.n285 71.676
R1126 B.n348 B.n286 71.676
R1127 B.n344 B.n287 71.676
R1128 B.n340 B.n288 71.676
R1129 B.n336 B.n289 71.676
R1130 B.n332 B.n290 71.676
R1131 B.n328 B.n291 71.676
R1132 B.n324 B.n292 71.676
R1133 B.n320 B.n293 71.676
R1134 B.n316 B.n294 71.676
R1135 B.n312 B.n295 71.676
R1136 B.n308 B.n296 71.676
R1137 B.n297 B.n261 71.676
R1138 B.n305 B.n304 59.5399
R1139 B.n302 B.n301 59.5399
R1140 B.n143 B.n76 59.5399
R1141 B.n164 B.n74 59.5399
R1142 B.n459 B.n258 51.7115
R1143 B.n459 B.n254 51.7115
R1144 B.n465 B.n254 51.7115
R1145 B.n465 B.n250 51.7115
R1146 B.n471 B.n250 51.7115
R1147 B.n477 B.n246 51.7115
R1148 B.n477 B.n242 51.7115
R1149 B.n483 B.n242 51.7115
R1150 B.n483 B.n238 51.7115
R1151 B.n489 B.n238 51.7115
R1152 B.n489 B.n234 51.7115
R1153 B.n496 B.n234 51.7115
R1154 B.n502 B.n230 51.7115
R1155 B.n502 B.n4 51.7115
R1156 B.n565 B.n4 51.7115
R1157 B.n565 B.n564 51.7115
R1158 B.n564 B.n563 51.7115
R1159 B.n563 B.n8 51.7115
R1160 B.n557 B.n556 51.7115
R1161 B.n556 B.n555 51.7115
R1162 B.n555 B.n15 51.7115
R1163 B.n549 B.n15 51.7115
R1164 B.n549 B.n548 51.7115
R1165 B.n548 B.n547 51.7115
R1166 B.n547 B.n22 51.7115
R1167 B.n541 B.n540 51.7115
R1168 B.n540 B.n539 51.7115
R1169 B.n539 B.n29 51.7115
R1170 B.n533 B.n29 51.7115
R1171 B.n533 B.n532 51.7115
R1172 B.t1 B.n230 44.8674
R1173 B.t0 B.n8 44.8674
R1174 B.n78 B.n31 35.7468
R1175 B.n528 B.n527 35.7468
R1176 B.n456 B.n455 35.7468
R1177 B.n450 B.n256 35.7468
R1178 B.t3 B.n246 31.1792
R1179 B.t7 B.n22 31.1792
R1180 B.n304 B.n303 29.8672
R1181 B.n301 B.n300 29.8672
R1182 B.n76 B.n75 29.8672
R1183 B.n74 B.n73 29.8672
R1184 B.n471 B.t3 20.5328
R1185 B.n541 B.t7 20.5328
R1186 B B.n567 18.0485
R1187 B.n79 B.n78 10.6151
R1188 B.n82 B.n79 10.6151
R1189 B.n83 B.n82 10.6151
R1190 B.n86 B.n83 10.6151
R1191 B.n87 B.n86 10.6151
R1192 B.n90 B.n87 10.6151
R1193 B.n91 B.n90 10.6151
R1194 B.n94 B.n91 10.6151
R1195 B.n95 B.n94 10.6151
R1196 B.n98 B.n95 10.6151
R1197 B.n99 B.n98 10.6151
R1198 B.n102 B.n99 10.6151
R1199 B.n103 B.n102 10.6151
R1200 B.n106 B.n103 10.6151
R1201 B.n107 B.n106 10.6151
R1202 B.n110 B.n107 10.6151
R1203 B.n111 B.n110 10.6151
R1204 B.n114 B.n111 10.6151
R1205 B.n115 B.n114 10.6151
R1206 B.n118 B.n115 10.6151
R1207 B.n119 B.n118 10.6151
R1208 B.n122 B.n119 10.6151
R1209 B.n123 B.n122 10.6151
R1210 B.n126 B.n123 10.6151
R1211 B.n127 B.n126 10.6151
R1212 B.n130 B.n127 10.6151
R1213 B.n131 B.n130 10.6151
R1214 B.n134 B.n131 10.6151
R1215 B.n135 B.n134 10.6151
R1216 B.n138 B.n135 10.6151
R1217 B.n139 B.n138 10.6151
R1218 B.n142 B.n139 10.6151
R1219 B.n147 B.n144 10.6151
R1220 B.n148 B.n147 10.6151
R1221 B.n151 B.n148 10.6151
R1222 B.n152 B.n151 10.6151
R1223 B.n155 B.n152 10.6151
R1224 B.n156 B.n155 10.6151
R1225 B.n159 B.n156 10.6151
R1226 B.n160 B.n159 10.6151
R1227 B.n163 B.n160 10.6151
R1228 B.n168 B.n165 10.6151
R1229 B.n169 B.n168 10.6151
R1230 B.n172 B.n169 10.6151
R1231 B.n173 B.n172 10.6151
R1232 B.n176 B.n173 10.6151
R1233 B.n177 B.n176 10.6151
R1234 B.n180 B.n177 10.6151
R1235 B.n181 B.n180 10.6151
R1236 B.n184 B.n181 10.6151
R1237 B.n185 B.n184 10.6151
R1238 B.n188 B.n185 10.6151
R1239 B.n189 B.n188 10.6151
R1240 B.n192 B.n189 10.6151
R1241 B.n193 B.n192 10.6151
R1242 B.n196 B.n193 10.6151
R1243 B.n197 B.n196 10.6151
R1244 B.n200 B.n197 10.6151
R1245 B.n201 B.n200 10.6151
R1246 B.n204 B.n201 10.6151
R1247 B.n205 B.n204 10.6151
R1248 B.n208 B.n205 10.6151
R1249 B.n209 B.n208 10.6151
R1250 B.n212 B.n209 10.6151
R1251 B.n213 B.n212 10.6151
R1252 B.n216 B.n213 10.6151
R1253 B.n217 B.n216 10.6151
R1254 B.n220 B.n217 10.6151
R1255 B.n221 B.n220 10.6151
R1256 B.n224 B.n221 10.6151
R1257 B.n226 B.n224 10.6151
R1258 B.n227 B.n226 10.6151
R1259 B.n528 B.n227 10.6151
R1260 B.n457 B.n456 10.6151
R1261 B.n457 B.n252 10.6151
R1262 B.n467 B.n252 10.6151
R1263 B.n468 B.n467 10.6151
R1264 B.n469 B.n468 10.6151
R1265 B.n469 B.n244 10.6151
R1266 B.n479 B.n244 10.6151
R1267 B.n480 B.n479 10.6151
R1268 B.n481 B.n480 10.6151
R1269 B.n481 B.n236 10.6151
R1270 B.n491 B.n236 10.6151
R1271 B.n492 B.n491 10.6151
R1272 B.n494 B.n492 10.6151
R1273 B.n494 B.n493 10.6151
R1274 B.n493 B.n228 10.6151
R1275 B.n505 B.n228 10.6151
R1276 B.n506 B.n505 10.6151
R1277 B.n507 B.n506 10.6151
R1278 B.n508 B.n507 10.6151
R1279 B.n510 B.n508 10.6151
R1280 B.n511 B.n510 10.6151
R1281 B.n512 B.n511 10.6151
R1282 B.n513 B.n512 10.6151
R1283 B.n515 B.n513 10.6151
R1284 B.n516 B.n515 10.6151
R1285 B.n517 B.n516 10.6151
R1286 B.n518 B.n517 10.6151
R1287 B.n520 B.n518 10.6151
R1288 B.n521 B.n520 10.6151
R1289 B.n522 B.n521 10.6151
R1290 B.n523 B.n522 10.6151
R1291 B.n525 B.n523 10.6151
R1292 B.n526 B.n525 10.6151
R1293 B.n527 B.n526 10.6151
R1294 B.n450 B.n449 10.6151
R1295 B.n449 B.n448 10.6151
R1296 B.n448 B.n447 10.6151
R1297 B.n447 B.n445 10.6151
R1298 B.n445 B.n442 10.6151
R1299 B.n442 B.n441 10.6151
R1300 B.n441 B.n438 10.6151
R1301 B.n438 B.n437 10.6151
R1302 B.n437 B.n434 10.6151
R1303 B.n434 B.n433 10.6151
R1304 B.n433 B.n430 10.6151
R1305 B.n430 B.n429 10.6151
R1306 B.n429 B.n426 10.6151
R1307 B.n426 B.n425 10.6151
R1308 B.n425 B.n422 10.6151
R1309 B.n422 B.n421 10.6151
R1310 B.n421 B.n418 10.6151
R1311 B.n418 B.n417 10.6151
R1312 B.n417 B.n414 10.6151
R1313 B.n414 B.n413 10.6151
R1314 B.n413 B.n410 10.6151
R1315 B.n410 B.n409 10.6151
R1316 B.n409 B.n406 10.6151
R1317 B.n406 B.n405 10.6151
R1318 B.n405 B.n402 10.6151
R1319 B.n402 B.n401 10.6151
R1320 B.n401 B.n398 10.6151
R1321 B.n398 B.n397 10.6151
R1322 B.n397 B.n394 10.6151
R1323 B.n394 B.n393 10.6151
R1324 B.n393 B.n390 10.6151
R1325 B.n390 B.n389 10.6151
R1326 B.n386 B.n385 10.6151
R1327 B.n385 B.n382 10.6151
R1328 B.n382 B.n381 10.6151
R1329 B.n381 B.n378 10.6151
R1330 B.n378 B.n377 10.6151
R1331 B.n377 B.n374 10.6151
R1332 B.n374 B.n373 10.6151
R1333 B.n373 B.n370 10.6151
R1334 B.n370 B.n369 10.6151
R1335 B.n366 B.n365 10.6151
R1336 B.n365 B.n362 10.6151
R1337 B.n362 B.n361 10.6151
R1338 B.n361 B.n358 10.6151
R1339 B.n358 B.n357 10.6151
R1340 B.n357 B.n354 10.6151
R1341 B.n354 B.n353 10.6151
R1342 B.n353 B.n350 10.6151
R1343 B.n350 B.n349 10.6151
R1344 B.n349 B.n346 10.6151
R1345 B.n346 B.n345 10.6151
R1346 B.n345 B.n342 10.6151
R1347 B.n342 B.n341 10.6151
R1348 B.n341 B.n338 10.6151
R1349 B.n338 B.n337 10.6151
R1350 B.n337 B.n334 10.6151
R1351 B.n334 B.n333 10.6151
R1352 B.n333 B.n330 10.6151
R1353 B.n330 B.n329 10.6151
R1354 B.n329 B.n326 10.6151
R1355 B.n326 B.n325 10.6151
R1356 B.n325 B.n322 10.6151
R1357 B.n322 B.n321 10.6151
R1358 B.n321 B.n318 10.6151
R1359 B.n318 B.n317 10.6151
R1360 B.n317 B.n314 10.6151
R1361 B.n314 B.n313 10.6151
R1362 B.n313 B.n310 10.6151
R1363 B.n310 B.n309 10.6151
R1364 B.n309 B.n306 10.6151
R1365 B.n306 B.n260 10.6151
R1366 B.n455 B.n260 10.6151
R1367 B.n461 B.n256 10.6151
R1368 B.n462 B.n461 10.6151
R1369 B.n463 B.n462 10.6151
R1370 B.n463 B.n248 10.6151
R1371 B.n473 B.n248 10.6151
R1372 B.n474 B.n473 10.6151
R1373 B.n475 B.n474 10.6151
R1374 B.n475 B.n240 10.6151
R1375 B.n485 B.n240 10.6151
R1376 B.n486 B.n485 10.6151
R1377 B.n487 B.n486 10.6151
R1378 B.n487 B.n232 10.6151
R1379 B.n498 B.n232 10.6151
R1380 B.n499 B.n498 10.6151
R1381 B.n500 B.n499 10.6151
R1382 B.n500 B.n0 10.6151
R1383 B.n561 B.n1 10.6151
R1384 B.n561 B.n560 10.6151
R1385 B.n560 B.n559 10.6151
R1386 B.n559 B.n10 10.6151
R1387 B.n553 B.n10 10.6151
R1388 B.n553 B.n552 10.6151
R1389 B.n552 B.n551 10.6151
R1390 B.n551 B.n17 10.6151
R1391 B.n545 B.n17 10.6151
R1392 B.n545 B.n544 10.6151
R1393 B.n544 B.n543 10.6151
R1394 B.n543 B.n24 10.6151
R1395 B.n537 B.n24 10.6151
R1396 B.n537 B.n536 10.6151
R1397 B.n536 B.n535 10.6151
R1398 B.n535 B.n31 10.6151
R1399 B.n143 B.n142 9.36635
R1400 B.n165 B.n164 9.36635
R1401 B.n389 B.n302 9.36635
R1402 B.n366 B.n305 9.36635
R1403 B.n496 B.t1 6.84461
R1404 B.n557 B.t0 6.84461
R1405 B.n567 B.n0 2.81026
R1406 B.n567 B.n1 2.81026
R1407 B.n144 B.n143 1.24928
R1408 B.n164 B.n163 1.24928
R1409 B.n386 B.n302 1.24928
R1410 B.n369 B.n305 1.24928
R1411 VP.n0 VP.t0 335.151
R1412 VP.n0 VP.t1 296.308
R1413 VP VP.n0 0.146778
R1414 VDD1.n44 VDD1.n0 289.615
R1415 VDD1.n93 VDD1.n49 289.615
R1416 VDD1.n45 VDD1.n44 185
R1417 VDD1.n43 VDD1.n42 185
R1418 VDD1.n4 VDD1.n3 185
R1419 VDD1.n8 VDD1.n6 185
R1420 VDD1.n37 VDD1.n36 185
R1421 VDD1.n35 VDD1.n34 185
R1422 VDD1.n10 VDD1.n9 185
R1423 VDD1.n29 VDD1.n28 185
R1424 VDD1.n27 VDD1.n26 185
R1425 VDD1.n14 VDD1.n13 185
R1426 VDD1.n21 VDD1.n20 185
R1427 VDD1.n19 VDD1.n18 185
R1428 VDD1.n66 VDD1.n65 185
R1429 VDD1.n68 VDD1.n67 185
R1430 VDD1.n61 VDD1.n60 185
R1431 VDD1.n74 VDD1.n73 185
R1432 VDD1.n76 VDD1.n75 185
R1433 VDD1.n57 VDD1.n56 185
R1434 VDD1.n83 VDD1.n82 185
R1435 VDD1.n84 VDD1.n55 185
R1436 VDD1.n86 VDD1.n85 185
R1437 VDD1.n53 VDD1.n52 185
R1438 VDD1.n92 VDD1.n91 185
R1439 VDD1.n94 VDD1.n93 185
R1440 VDD1.n17 VDD1.t1 149.524
R1441 VDD1.n64 VDD1.t0 149.524
R1442 VDD1.n44 VDD1.n43 104.615
R1443 VDD1.n43 VDD1.n3 104.615
R1444 VDD1.n8 VDD1.n3 104.615
R1445 VDD1.n36 VDD1.n8 104.615
R1446 VDD1.n36 VDD1.n35 104.615
R1447 VDD1.n35 VDD1.n9 104.615
R1448 VDD1.n28 VDD1.n9 104.615
R1449 VDD1.n28 VDD1.n27 104.615
R1450 VDD1.n27 VDD1.n13 104.615
R1451 VDD1.n20 VDD1.n13 104.615
R1452 VDD1.n20 VDD1.n19 104.615
R1453 VDD1.n67 VDD1.n66 104.615
R1454 VDD1.n67 VDD1.n60 104.615
R1455 VDD1.n74 VDD1.n60 104.615
R1456 VDD1.n75 VDD1.n74 104.615
R1457 VDD1.n75 VDD1.n56 104.615
R1458 VDD1.n83 VDD1.n56 104.615
R1459 VDD1.n84 VDD1.n83 104.615
R1460 VDD1.n85 VDD1.n84 104.615
R1461 VDD1.n85 VDD1.n52 104.615
R1462 VDD1.n92 VDD1.n52 104.615
R1463 VDD1.n93 VDD1.n92 104.615
R1464 VDD1 VDD1.n97 82.9882
R1465 VDD1.n19 VDD1.t1 52.3082
R1466 VDD1.n66 VDD1.t0 52.3082
R1467 VDD1 VDD1.n48 48.2845
R1468 VDD1.n6 VDD1.n4 13.1884
R1469 VDD1.n86 VDD1.n53 13.1884
R1470 VDD1.n42 VDD1.n41 12.8005
R1471 VDD1.n38 VDD1.n37 12.8005
R1472 VDD1.n87 VDD1.n55 12.8005
R1473 VDD1.n91 VDD1.n90 12.8005
R1474 VDD1.n45 VDD1.n2 12.0247
R1475 VDD1.n34 VDD1.n7 12.0247
R1476 VDD1.n82 VDD1.n81 12.0247
R1477 VDD1.n94 VDD1.n51 12.0247
R1478 VDD1.n46 VDD1.n0 11.249
R1479 VDD1.n33 VDD1.n10 11.249
R1480 VDD1.n80 VDD1.n57 11.249
R1481 VDD1.n95 VDD1.n49 11.249
R1482 VDD1.n30 VDD1.n29 10.4732
R1483 VDD1.n77 VDD1.n76 10.4732
R1484 VDD1.n18 VDD1.n17 10.2747
R1485 VDD1.n65 VDD1.n64 10.2747
R1486 VDD1.n26 VDD1.n12 9.69747
R1487 VDD1.n73 VDD1.n59 9.69747
R1488 VDD1.n48 VDD1.n47 9.45567
R1489 VDD1.n97 VDD1.n96 9.45567
R1490 VDD1.n16 VDD1.n15 9.3005
R1491 VDD1.n23 VDD1.n22 9.3005
R1492 VDD1.n25 VDD1.n24 9.3005
R1493 VDD1.n12 VDD1.n11 9.3005
R1494 VDD1.n31 VDD1.n30 9.3005
R1495 VDD1.n33 VDD1.n32 9.3005
R1496 VDD1.n7 VDD1.n5 9.3005
R1497 VDD1.n39 VDD1.n38 9.3005
R1498 VDD1.n47 VDD1.n46 9.3005
R1499 VDD1.n2 VDD1.n1 9.3005
R1500 VDD1.n41 VDD1.n40 9.3005
R1501 VDD1.n96 VDD1.n95 9.3005
R1502 VDD1.n51 VDD1.n50 9.3005
R1503 VDD1.n90 VDD1.n89 9.3005
R1504 VDD1.n63 VDD1.n62 9.3005
R1505 VDD1.n70 VDD1.n69 9.3005
R1506 VDD1.n72 VDD1.n71 9.3005
R1507 VDD1.n59 VDD1.n58 9.3005
R1508 VDD1.n78 VDD1.n77 9.3005
R1509 VDD1.n80 VDD1.n79 9.3005
R1510 VDD1.n81 VDD1.n54 9.3005
R1511 VDD1.n88 VDD1.n87 9.3005
R1512 VDD1.n25 VDD1.n14 8.92171
R1513 VDD1.n72 VDD1.n61 8.92171
R1514 VDD1.n22 VDD1.n21 8.14595
R1515 VDD1.n69 VDD1.n68 8.14595
R1516 VDD1.n18 VDD1.n16 7.3702
R1517 VDD1.n65 VDD1.n63 7.3702
R1518 VDD1.n21 VDD1.n16 5.81868
R1519 VDD1.n68 VDD1.n63 5.81868
R1520 VDD1.n22 VDD1.n14 5.04292
R1521 VDD1.n69 VDD1.n61 5.04292
R1522 VDD1.n26 VDD1.n25 4.26717
R1523 VDD1.n73 VDD1.n72 4.26717
R1524 VDD1.n29 VDD1.n12 3.49141
R1525 VDD1.n76 VDD1.n59 3.49141
R1526 VDD1.n17 VDD1.n15 2.84303
R1527 VDD1.n64 VDD1.n62 2.84303
R1528 VDD1.n48 VDD1.n0 2.71565
R1529 VDD1.n30 VDD1.n10 2.71565
R1530 VDD1.n77 VDD1.n57 2.71565
R1531 VDD1.n97 VDD1.n49 2.71565
R1532 VDD1.n46 VDD1.n45 1.93989
R1533 VDD1.n34 VDD1.n33 1.93989
R1534 VDD1.n82 VDD1.n80 1.93989
R1535 VDD1.n95 VDD1.n94 1.93989
R1536 VDD1.n42 VDD1.n2 1.16414
R1537 VDD1.n37 VDD1.n7 1.16414
R1538 VDD1.n81 VDD1.n55 1.16414
R1539 VDD1.n91 VDD1.n51 1.16414
R1540 VDD1.n41 VDD1.n4 0.388379
R1541 VDD1.n38 VDD1.n6 0.388379
R1542 VDD1.n87 VDD1.n86 0.388379
R1543 VDD1.n90 VDD1.n53 0.388379
R1544 VDD1.n47 VDD1.n1 0.155672
R1545 VDD1.n40 VDD1.n1 0.155672
R1546 VDD1.n40 VDD1.n39 0.155672
R1547 VDD1.n39 VDD1.n5 0.155672
R1548 VDD1.n32 VDD1.n5 0.155672
R1549 VDD1.n32 VDD1.n31 0.155672
R1550 VDD1.n31 VDD1.n11 0.155672
R1551 VDD1.n24 VDD1.n11 0.155672
R1552 VDD1.n24 VDD1.n23 0.155672
R1553 VDD1.n23 VDD1.n15 0.155672
R1554 VDD1.n70 VDD1.n62 0.155672
R1555 VDD1.n71 VDD1.n70 0.155672
R1556 VDD1.n71 VDD1.n58 0.155672
R1557 VDD1.n78 VDD1.n58 0.155672
R1558 VDD1.n79 VDD1.n78 0.155672
R1559 VDD1.n79 VDD1.n54 0.155672
R1560 VDD1.n88 VDD1.n54 0.155672
R1561 VDD1.n89 VDD1.n88 0.155672
R1562 VDD1.n89 VDD1.n50 0.155672
R1563 VDD1.n96 VDD1.n50 0.155672
C0 VDD1 VTAIL 4.2857f
C1 VDD2 VTAIL 4.32581f
C2 VTAIL VN 1.5507f
C3 VDD1 VP 1.99007f
C4 VDD2 VP 0.274534f
C5 VP VN 4.285089f
C6 VDD2 VDD1 0.513749f
C7 VDD1 VN 0.147485f
C8 VDD2 VN 1.86586f
C9 VP VTAIL 1.56508f
C10 VDD2 B 3.41281f
C11 VDD1 B 4.98144f
C12 VTAIL B 5.525799f
C13 VN B 6.86806f
C14 VP B 4.464707f
C15 VDD1.n0 B 0.017751f
C16 VDD1.n1 B 0.014045f
C17 VDD1.n2 B 0.007547f
C18 VDD1.n3 B 0.017838f
C19 VDD1.n4 B 0.007769f
C20 VDD1.n5 B 0.014045f
C21 VDD1.n6 B 0.007769f
C22 VDD1.n7 B 0.007547f
C23 VDD1.n8 B 0.017838f
C24 VDD1.n9 B 0.017838f
C25 VDD1.n10 B 0.007991f
C26 VDD1.n11 B 0.014045f
C27 VDD1.n12 B 0.007547f
C28 VDD1.n13 B 0.017838f
C29 VDD1.n14 B 0.007991f
C30 VDD1.n15 B 0.53298f
C31 VDD1.n16 B 0.007547f
C32 VDD1.t1 B 0.029916f
C33 VDD1.n17 B 0.08611f
C34 VDD1.n18 B 0.01261f
C35 VDD1.n19 B 0.013379f
C36 VDD1.n20 B 0.017838f
C37 VDD1.n21 B 0.007991f
C38 VDD1.n22 B 0.007547f
C39 VDD1.n23 B 0.014045f
C40 VDD1.n24 B 0.014045f
C41 VDD1.n25 B 0.007547f
C42 VDD1.n26 B 0.007991f
C43 VDD1.n27 B 0.017838f
C44 VDD1.n28 B 0.017838f
C45 VDD1.n29 B 0.007991f
C46 VDD1.n30 B 0.007547f
C47 VDD1.n31 B 0.014045f
C48 VDD1.n32 B 0.014045f
C49 VDD1.n33 B 0.007547f
C50 VDD1.n34 B 0.007991f
C51 VDD1.n35 B 0.017838f
C52 VDD1.n36 B 0.017838f
C53 VDD1.n37 B 0.007991f
C54 VDD1.n38 B 0.007547f
C55 VDD1.n39 B 0.014045f
C56 VDD1.n40 B 0.014045f
C57 VDD1.n41 B 0.007547f
C58 VDD1.n42 B 0.007991f
C59 VDD1.n43 B 0.017838f
C60 VDD1.n44 B 0.035097f
C61 VDD1.n45 B 0.007991f
C62 VDD1.n46 B 0.007547f
C63 VDD1.n47 B 0.031504f
C64 VDD1.n48 B 0.029309f
C65 VDD1.n49 B 0.017751f
C66 VDD1.n50 B 0.014045f
C67 VDD1.n51 B 0.007547f
C68 VDD1.n52 B 0.017838f
C69 VDD1.n53 B 0.007769f
C70 VDD1.n54 B 0.014045f
C71 VDD1.n55 B 0.007991f
C72 VDD1.n56 B 0.017838f
C73 VDD1.n57 B 0.007991f
C74 VDD1.n58 B 0.014045f
C75 VDD1.n59 B 0.007547f
C76 VDD1.n60 B 0.017838f
C77 VDD1.n61 B 0.007991f
C78 VDD1.n62 B 0.53298f
C79 VDD1.n63 B 0.007547f
C80 VDD1.t0 B 0.029916f
C81 VDD1.n64 B 0.08611f
C82 VDD1.n65 B 0.01261f
C83 VDD1.n66 B 0.013379f
C84 VDD1.n67 B 0.017838f
C85 VDD1.n68 B 0.007991f
C86 VDD1.n69 B 0.007547f
C87 VDD1.n70 B 0.014045f
C88 VDD1.n71 B 0.014045f
C89 VDD1.n72 B 0.007547f
C90 VDD1.n73 B 0.007991f
C91 VDD1.n74 B 0.017838f
C92 VDD1.n75 B 0.017838f
C93 VDD1.n76 B 0.007991f
C94 VDD1.n77 B 0.007547f
C95 VDD1.n78 B 0.014045f
C96 VDD1.n79 B 0.014045f
C97 VDD1.n80 B 0.007547f
C98 VDD1.n81 B 0.007547f
C99 VDD1.n82 B 0.007991f
C100 VDD1.n83 B 0.017838f
C101 VDD1.n84 B 0.017838f
C102 VDD1.n85 B 0.017838f
C103 VDD1.n86 B 0.007769f
C104 VDD1.n87 B 0.007547f
C105 VDD1.n88 B 0.014045f
C106 VDD1.n89 B 0.014045f
C107 VDD1.n90 B 0.007547f
C108 VDD1.n91 B 0.007991f
C109 VDD1.n92 B 0.017838f
C110 VDD1.n93 B 0.035097f
C111 VDD1.n94 B 0.007991f
C112 VDD1.n95 B 0.007547f
C113 VDD1.n96 B 0.031504f
C114 VDD1.n97 B 0.331553f
C115 VP.t0 B 1.06607f
C116 VP.t1 B 0.925564f
C117 VP.n0 B 2.28594f
C118 VDD2.n0 B 0.017968f
C119 VDD2.n1 B 0.014216f
C120 VDD2.n2 B 0.007639f
C121 VDD2.n3 B 0.018056f
C122 VDD2.n4 B 0.007864f
C123 VDD2.n5 B 0.014216f
C124 VDD2.n6 B 0.008088f
C125 VDD2.n7 B 0.018056f
C126 VDD2.n8 B 0.008088f
C127 VDD2.n9 B 0.014216f
C128 VDD2.n10 B 0.007639f
C129 VDD2.n11 B 0.018056f
C130 VDD2.n12 B 0.008088f
C131 VDD2.n13 B 0.539488f
C132 VDD2.n14 B 0.007639f
C133 VDD2.t1 B 0.030282f
C134 VDD2.n15 B 0.087162f
C135 VDD2.n16 B 0.012764f
C136 VDD2.n17 B 0.013542f
C137 VDD2.n18 B 0.018056f
C138 VDD2.n19 B 0.008088f
C139 VDD2.n20 B 0.007639f
C140 VDD2.n21 B 0.014216f
C141 VDD2.n22 B 0.014216f
C142 VDD2.n23 B 0.007639f
C143 VDD2.n24 B 0.008088f
C144 VDD2.n25 B 0.018056f
C145 VDD2.n26 B 0.018056f
C146 VDD2.n27 B 0.008088f
C147 VDD2.n28 B 0.007639f
C148 VDD2.n29 B 0.014216f
C149 VDD2.n30 B 0.014216f
C150 VDD2.n31 B 0.007639f
C151 VDD2.n32 B 0.007639f
C152 VDD2.n33 B 0.008088f
C153 VDD2.n34 B 0.018056f
C154 VDD2.n35 B 0.018056f
C155 VDD2.n36 B 0.018056f
C156 VDD2.n37 B 0.007864f
C157 VDD2.n38 B 0.007639f
C158 VDD2.n39 B 0.014216f
C159 VDD2.n40 B 0.014216f
C160 VDD2.n41 B 0.007639f
C161 VDD2.n42 B 0.008088f
C162 VDD2.n43 B 0.018056f
C163 VDD2.n44 B 0.035526f
C164 VDD2.n45 B 0.008088f
C165 VDD2.n46 B 0.007639f
C166 VDD2.n47 B 0.031888f
C167 VDD2.n48 B 0.315257f
C168 VDD2.n49 B 0.017968f
C169 VDD2.n50 B 0.014216f
C170 VDD2.n51 B 0.007639f
C171 VDD2.n52 B 0.018056f
C172 VDD2.n53 B 0.007864f
C173 VDD2.n54 B 0.014216f
C174 VDD2.n55 B 0.007864f
C175 VDD2.n56 B 0.007639f
C176 VDD2.n57 B 0.018056f
C177 VDD2.n58 B 0.018056f
C178 VDD2.n59 B 0.008088f
C179 VDD2.n60 B 0.014216f
C180 VDD2.n61 B 0.007639f
C181 VDD2.n62 B 0.018056f
C182 VDD2.n63 B 0.008088f
C183 VDD2.n64 B 0.539488f
C184 VDD2.n65 B 0.007639f
C185 VDD2.t0 B 0.030282f
C186 VDD2.n66 B 0.087162f
C187 VDD2.n67 B 0.012764f
C188 VDD2.n68 B 0.013542f
C189 VDD2.n69 B 0.018056f
C190 VDD2.n70 B 0.008088f
C191 VDD2.n71 B 0.007639f
C192 VDD2.n72 B 0.014216f
C193 VDD2.n73 B 0.014216f
C194 VDD2.n74 B 0.007639f
C195 VDD2.n75 B 0.008088f
C196 VDD2.n76 B 0.018056f
C197 VDD2.n77 B 0.018056f
C198 VDD2.n78 B 0.008088f
C199 VDD2.n79 B 0.007639f
C200 VDD2.n80 B 0.014216f
C201 VDD2.n81 B 0.014216f
C202 VDD2.n82 B 0.007639f
C203 VDD2.n83 B 0.008088f
C204 VDD2.n84 B 0.018056f
C205 VDD2.n85 B 0.018056f
C206 VDD2.n86 B 0.008088f
C207 VDD2.n87 B 0.007639f
C208 VDD2.n88 B 0.014216f
C209 VDD2.n89 B 0.014216f
C210 VDD2.n90 B 0.007639f
C211 VDD2.n91 B 0.008088f
C212 VDD2.n92 B 0.018056f
C213 VDD2.n93 B 0.035526f
C214 VDD2.n94 B 0.008088f
C215 VDD2.n95 B 0.007639f
C216 VDD2.n96 B 0.031888f
C217 VDD2.n97 B 0.029306f
C218 VDD2.n98 B 1.40742f
C219 VTAIL.n0 B 0.019511f
C220 VTAIL.n1 B 0.015437f
C221 VTAIL.n2 B 0.008295f
C222 VTAIL.n3 B 0.019607f
C223 VTAIL.n4 B 0.008539f
C224 VTAIL.n5 B 0.015437f
C225 VTAIL.n6 B 0.008783f
C226 VTAIL.n7 B 0.019607f
C227 VTAIL.n8 B 0.008783f
C228 VTAIL.n9 B 0.015437f
C229 VTAIL.n10 B 0.008295f
C230 VTAIL.n11 B 0.019607f
C231 VTAIL.n12 B 0.008783f
C232 VTAIL.n13 B 0.585835f
C233 VTAIL.n14 B 0.008295f
C234 VTAIL.t1 B 0.032883f
C235 VTAIL.n15 B 0.09465f
C236 VTAIL.n16 B 0.013861f
C237 VTAIL.n17 B 0.014705f
C238 VTAIL.n18 B 0.019607f
C239 VTAIL.n19 B 0.008783f
C240 VTAIL.n20 B 0.008295f
C241 VTAIL.n21 B 0.015437f
C242 VTAIL.n22 B 0.015437f
C243 VTAIL.n23 B 0.008295f
C244 VTAIL.n24 B 0.008783f
C245 VTAIL.n25 B 0.019607f
C246 VTAIL.n26 B 0.019607f
C247 VTAIL.n27 B 0.008783f
C248 VTAIL.n28 B 0.008295f
C249 VTAIL.n29 B 0.015437f
C250 VTAIL.n30 B 0.015437f
C251 VTAIL.n31 B 0.008295f
C252 VTAIL.n32 B 0.008295f
C253 VTAIL.n33 B 0.008783f
C254 VTAIL.n34 B 0.019607f
C255 VTAIL.n35 B 0.019607f
C256 VTAIL.n36 B 0.019607f
C257 VTAIL.n37 B 0.008539f
C258 VTAIL.n38 B 0.008295f
C259 VTAIL.n39 B 0.015437f
C260 VTAIL.n40 B 0.015437f
C261 VTAIL.n41 B 0.008295f
C262 VTAIL.n42 B 0.008783f
C263 VTAIL.n43 B 0.019607f
C264 VTAIL.n44 B 0.038578f
C265 VTAIL.n45 B 0.008783f
C266 VTAIL.n46 B 0.008295f
C267 VTAIL.n47 B 0.034628f
C268 VTAIL.n48 B 0.021156f
C269 VTAIL.n49 B 0.791214f
C270 VTAIL.n50 B 0.019511f
C271 VTAIL.n51 B 0.015437f
C272 VTAIL.n52 B 0.008295f
C273 VTAIL.n53 B 0.019607f
C274 VTAIL.n54 B 0.008539f
C275 VTAIL.n55 B 0.015437f
C276 VTAIL.n56 B 0.008539f
C277 VTAIL.n57 B 0.008295f
C278 VTAIL.n58 B 0.019607f
C279 VTAIL.n59 B 0.019607f
C280 VTAIL.n60 B 0.008783f
C281 VTAIL.n61 B 0.015437f
C282 VTAIL.n62 B 0.008295f
C283 VTAIL.n63 B 0.019607f
C284 VTAIL.n64 B 0.008783f
C285 VTAIL.n65 B 0.585835f
C286 VTAIL.n66 B 0.008295f
C287 VTAIL.t2 B 0.032883f
C288 VTAIL.n67 B 0.09465f
C289 VTAIL.n68 B 0.013861f
C290 VTAIL.n69 B 0.014705f
C291 VTAIL.n70 B 0.019607f
C292 VTAIL.n71 B 0.008783f
C293 VTAIL.n72 B 0.008295f
C294 VTAIL.n73 B 0.015437f
C295 VTAIL.n74 B 0.015437f
C296 VTAIL.n75 B 0.008295f
C297 VTAIL.n76 B 0.008783f
C298 VTAIL.n77 B 0.019607f
C299 VTAIL.n78 B 0.019607f
C300 VTAIL.n79 B 0.008783f
C301 VTAIL.n80 B 0.008295f
C302 VTAIL.n81 B 0.015437f
C303 VTAIL.n82 B 0.015437f
C304 VTAIL.n83 B 0.008295f
C305 VTAIL.n84 B 0.008783f
C306 VTAIL.n85 B 0.019607f
C307 VTAIL.n86 B 0.019607f
C308 VTAIL.n87 B 0.008783f
C309 VTAIL.n88 B 0.008295f
C310 VTAIL.n89 B 0.015437f
C311 VTAIL.n90 B 0.015437f
C312 VTAIL.n91 B 0.008295f
C313 VTAIL.n92 B 0.008783f
C314 VTAIL.n93 B 0.019607f
C315 VTAIL.n94 B 0.038578f
C316 VTAIL.n95 B 0.008783f
C317 VTAIL.n96 B 0.008295f
C318 VTAIL.n97 B 0.034628f
C319 VTAIL.n98 B 0.021156f
C320 VTAIL.n99 B 0.804829f
C321 VTAIL.n100 B 0.019511f
C322 VTAIL.n101 B 0.015437f
C323 VTAIL.n102 B 0.008295f
C324 VTAIL.n103 B 0.019607f
C325 VTAIL.n104 B 0.008539f
C326 VTAIL.n105 B 0.015437f
C327 VTAIL.n106 B 0.008539f
C328 VTAIL.n107 B 0.008295f
C329 VTAIL.n108 B 0.019607f
C330 VTAIL.n109 B 0.019607f
C331 VTAIL.n110 B 0.008783f
C332 VTAIL.n111 B 0.015437f
C333 VTAIL.n112 B 0.008295f
C334 VTAIL.n113 B 0.019607f
C335 VTAIL.n114 B 0.008783f
C336 VTAIL.n115 B 0.585835f
C337 VTAIL.n116 B 0.008295f
C338 VTAIL.t0 B 0.032883f
C339 VTAIL.n117 B 0.09465f
C340 VTAIL.n118 B 0.013861f
C341 VTAIL.n119 B 0.014705f
C342 VTAIL.n120 B 0.019607f
C343 VTAIL.n121 B 0.008783f
C344 VTAIL.n122 B 0.008295f
C345 VTAIL.n123 B 0.015437f
C346 VTAIL.n124 B 0.015437f
C347 VTAIL.n125 B 0.008295f
C348 VTAIL.n126 B 0.008783f
C349 VTAIL.n127 B 0.019607f
C350 VTAIL.n128 B 0.019607f
C351 VTAIL.n129 B 0.008783f
C352 VTAIL.n130 B 0.008295f
C353 VTAIL.n131 B 0.015437f
C354 VTAIL.n132 B 0.015437f
C355 VTAIL.n133 B 0.008295f
C356 VTAIL.n134 B 0.008783f
C357 VTAIL.n135 B 0.019607f
C358 VTAIL.n136 B 0.019607f
C359 VTAIL.n137 B 0.008783f
C360 VTAIL.n138 B 0.008295f
C361 VTAIL.n139 B 0.015437f
C362 VTAIL.n140 B 0.015437f
C363 VTAIL.n141 B 0.008295f
C364 VTAIL.n142 B 0.008783f
C365 VTAIL.n143 B 0.019607f
C366 VTAIL.n144 B 0.038578f
C367 VTAIL.n145 B 0.008783f
C368 VTAIL.n146 B 0.008295f
C369 VTAIL.n147 B 0.034628f
C370 VTAIL.n148 B 0.021156f
C371 VTAIL.n149 B 0.738792f
C372 VTAIL.n150 B 0.019511f
C373 VTAIL.n151 B 0.015437f
C374 VTAIL.n152 B 0.008295f
C375 VTAIL.n153 B 0.019607f
C376 VTAIL.n154 B 0.008539f
C377 VTAIL.n155 B 0.015437f
C378 VTAIL.n156 B 0.008783f
C379 VTAIL.n157 B 0.019607f
C380 VTAIL.n158 B 0.008783f
C381 VTAIL.n159 B 0.015437f
C382 VTAIL.n160 B 0.008295f
C383 VTAIL.n161 B 0.019607f
C384 VTAIL.n162 B 0.008783f
C385 VTAIL.n163 B 0.585835f
C386 VTAIL.n164 B 0.008295f
C387 VTAIL.t3 B 0.032883f
C388 VTAIL.n165 B 0.09465f
C389 VTAIL.n166 B 0.013861f
C390 VTAIL.n167 B 0.014705f
C391 VTAIL.n168 B 0.019607f
C392 VTAIL.n169 B 0.008783f
C393 VTAIL.n170 B 0.008295f
C394 VTAIL.n171 B 0.015437f
C395 VTAIL.n172 B 0.015437f
C396 VTAIL.n173 B 0.008295f
C397 VTAIL.n174 B 0.008783f
C398 VTAIL.n175 B 0.019607f
C399 VTAIL.n176 B 0.019607f
C400 VTAIL.n177 B 0.008783f
C401 VTAIL.n178 B 0.008295f
C402 VTAIL.n179 B 0.015437f
C403 VTAIL.n180 B 0.015437f
C404 VTAIL.n181 B 0.008295f
C405 VTAIL.n182 B 0.008295f
C406 VTAIL.n183 B 0.008783f
C407 VTAIL.n184 B 0.019607f
C408 VTAIL.n185 B 0.019607f
C409 VTAIL.n186 B 0.019607f
C410 VTAIL.n187 B 0.008539f
C411 VTAIL.n188 B 0.008295f
C412 VTAIL.n189 B 0.015437f
C413 VTAIL.n190 B 0.015437f
C414 VTAIL.n191 B 0.008295f
C415 VTAIL.n192 B 0.008783f
C416 VTAIL.n193 B 0.019607f
C417 VTAIL.n194 B 0.038578f
C418 VTAIL.n195 B 0.008783f
C419 VTAIL.n196 B 0.008295f
C420 VTAIL.n197 B 0.034628f
C421 VTAIL.n198 B 0.021156f
C422 VTAIL.n199 B 0.696017f
C423 VN.t0 B 0.917866f
C424 VN.t1 B 1.05966f
.ends

