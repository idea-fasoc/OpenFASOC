* NGSPICE file created from diff_pair_sample_0825.ext - technology: sky130A

.subckt diff_pair_sample_0825 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t16 VP.t0 VDD1.t5 w_n3874_n1526# sky130_fd_pr__pfet_01v8 ad=0.46035 pd=3.12 as=0.46035 ps=3.12 w=2.79 l=2.09
X1 VTAIL.t15 VP.t1 VDD1.t4 w_n3874_n1526# sky130_fd_pr__pfet_01v8 ad=0.46035 pd=3.12 as=0.46035 ps=3.12 w=2.79 l=2.09
X2 B.t11 B.t9 B.t10 w_n3874_n1526# sky130_fd_pr__pfet_01v8 ad=1.0881 pd=6.36 as=0 ps=0 w=2.79 l=2.09
X3 VDD2.t9 VN.t0 VTAIL.t17 w_n3874_n1526# sky130_fd_pr__pfet_01v8 ad=0.46035 pd=3.12 as=1.0881 ps=6.36 w=2.79 l=2.09
X4 VTAIL.t19 VN.t1 VDD2.t8 w_n3874_n1526# sky130_fd_pr__pfet_01v8 ad=0.46035 pd=3.12 as=0.46035 ps=3.12 w=2.79 l=2.09
X5 VTAIL.t18 VN.t2 VDD2.t7 w_n3874_n1526# sky130_fd_pr__pfet_01v8 ad=0.46035 pd=3.12 as=0.46035 ps=3.12 w=2.79 l=2.09
X6 B.t8 B.t6 B.t7 w_n3874_n1526# sky130_fd_pr__pfet_01v8 ad=1.0881 pd=6.36 as=0 ps=0 w=2.79 l=2.09
X7 VTAIL.t14 VP.t2 VDD1.t8 w_n3874_n1526# sky130_fd_pr__pfet_01v8 ad=0.46035 pd=3.12 as=0.46035 ps=3.12 w=2.79 l=2.09
X8 VDD1.t7 VP.t3 VTAIL.t13 w_n3874_n1526# sky130_fd_pr__pfet_01v8 ad=1.0881 pd=6.36 as=0.46035 ps=3.12 w=2.79 l=2.09
X9 VDD2.t6 VN.t3 VTAIL.t6 w_n3874_n1526# sky130_fd_pr__pfet_01v8 ad=0.46035 pd=3.12 as=1.0881 ps=6.36 w=2.79 l=2.09
X10 VTAIL.t4 VN.t4 VDD2.t5 w_n3874_n1526# sky130_fd_pr__pfet_01v8 ad=0.46035 pd=3.12 as=0.46035 ps=3.12 w=2.79 l=2.09
X11 VTAIL.t5 VN.t5 VDD2.t4 w_n3874_n1526# sky130_fd_pr__pfet_01v8 ad=0.46035 pd=3.12 as=0.46035 ps=3.12 w=2.79 l=2.09
X12 VDD2.t3 VN.t6 VTAIL.t0 w_n3874_n1526# sky130_fd_pr__pfet_01v8 ad=1.0881 pd=6.36 as=0.46035 ps=3.12 w=2.79 l=2.09
X13 VDD1.t2 VP.t4 VTAIL.t12 w_n3874_n1526# sky130_fd_pr__pfet_01v8 ad=0.46035 pd=3.12 as=1.0881 ps=6.36 w=2.79 l=2.09
X14 VDD2.t2 VN.t7 VTAIL.t1 w_n3874_n1526# sky130_fd_pr__pfet_01v8 ad=0.46035 pd=3.12 as=0.46035 ps=3.12 w=2.79 l=2.09
X15 B.t5 B.t3 B.t4 w_n3874_n1526# sky130_fd_pr__pfet_01v8 ad=1.0881 pd=6.36 as=0 ps=0 w=2.79 l=2.09
X16 VDD1.t0 VP.t5 VTAIL.t11 w_n3874_n1526# sky130_fd_pr__pfet_01v8 ad=0.46035 pd=3.12 as=0.46035 ps=3.12 w=2.79 l=2.09
X17 VDD1.t3 VP.t6 VTAIL.t10 w_n3874_n1526# sky130_fd_pr__pfet_01v8 ad=0.46035 pd=3.12 as=0.46035 ps=3.12 w=2.79 l=2.09
X18 VDD1.t1 VP.t7 VTAIL.t9 w_n3874_n1526# sky130_fd_pr__pfet_01v8 ad=0.46035 pd=3.12 as=1.0881 ps=6.36 w=2.79 l=2.09
X19 VDD2.t1 VN.t8 VTAIL.t3 w_n3874_n1526# sky130_fd_pr__pfet_01v8 ad=1.0881 pd=6.36 as=0.46035 ps=3.12 w=2.79 l=2.09
X20 VTAIL.t8 VP.t8 VDD1.t6 w_n3874_n1526# sky130_fd_pr__pfet_01v8 ad=0.46035 pd=3.12 as=0.46035 ps=3.12 w=2.79 l=2.09
X21 VDD1.t9 VP.t9 VTAIL.t7 w_n3874_n1526# sky130_fd_pr__pfet_01v8 ad=1.0881 pd=6.36 as=0.46035 ps=3.12 w=2.79 l=2.09
X22 VDD2.t0 VN.t9 VTAIL.t2 w_n3874_n1526# sky130_fd_pr__pfet_01v8 ad=0.46035 pd=3.12 as=0.46035 ps=3.12 w=2.79 l=2.09
X23 B.t2 B.t0 B.t1 w_n3874_n1526# sky130_fd_pr__pfet_01v8 ad=1.0881 pd=6.36 as=0 ps=0 w=2.79 l=2.09
R0 VP.n20 VP.n19 161.3
R1 VP.n21 VP.n16 161.3
R2 VP.n23 VP.n22 161.3
R3 VP.n24 VP.n15 161.3
R4 VP.n26 VP.n25 161.3
R5 VP.n27 VP.n14 161.3
R6 VP.n29 VP.n28 161.3
R7 VP.n30 VP.n13 161.3
R8 VP.n32 VP.n31 161.3
R9 VP.n34 VP.n12 161.3
R10 VP.n36 VP.n35 161.3
R11 VP.n37 VP.n11 161.3
R12 VP.n39 VP.n38 161.3
R13 VP.n40 VP.n10 161.3
R14 VP.n74 VP.n0 161.3
R15 VP.n73 VP.n72 161.3
R16 VP.n71 VP.n1 161.3
R17 VP.n70 VP.n69 161.3
R18 VP.n68 VP.n2 161.3
R19 VP.n66 VP.n65 161.3
R20 VP.n64 VP.n3 161.3
R21 VP.n63 VP.n62 161.3
R22 VP.n61 VP.n4 161.3
R23 VP.n60 VP.n59 161.3
R24 VP.n58 VP.n5 161.3
R25 VP.n57 VP.n56 161.3
R26 VP.n55 VP.n6 161.3
R27 VP.n54 VP.n53 161.3
R28 VP.n52 VP.n51 161.3
R29 VP.n50 VP.n8 161.3
R30 VP.n49 VP.n48 161.3
R31 VP.n47 VP.n9 161.3
R32 VP.n46 VP.n45 161.3
R33 VP.n44 VP.n43 94.1189
R34 VP.n76 VP.n75 94.1189
R35 VP.n42 VP.n41 94.1189
R36 VP.n18 VP.t3 65.6206
R37 VP.n56 VP.n55 56.5193
R38 VP.n62 VP.n3 56.5193
R39 VP.n28 VP.n13 56.5193
R40 VP.n22 VP.n21 56.5193
R41 VP.n49 VP.n9 53.1199
R42 VP.n73 VP.n1 53.1199
R43 VP.n39 VP.n11 53.1199
R44 VP.n18 VP.n17 50.0611
R45 VP.n43 VP.n42 43.3632
R46 VP.n60 VP.t5 32.1723
R47 VP.n44 VP.t9 32.1723
R48 VP.n7 VP.t2 32.1723
R49 VP.n67 VP.t0 32.1723
R50 VP.n75 VP.t7 32.1723
R51 VP.n26 VP.t6 32.1723
R52 VP.n41 VP.t4 32.1723
R53 VP.n33 VP.t1 32.1723
R54 VP.n17 VP.t8 32.1723
R55 VP.n50 VP.n49 27.8669
R56 VP.n69 VP.n1 27.8669
R57 VP.n35 VP.n11 27.8669
R58 VP.n45 VP.n9 24.4675
R59 VP.n51 VP.n50 24.4675
R60 VP.n55 VP.n54 24.4675
R61 VP.n56 VP.n5 24.4675
R62 VP.n60 VP.n5 24.4675
R63 VP.n61 VP.n60 24.4675
R64 VP.n62 VP.n61 24.4675
R65 VP.n66 VP.n3 24.4675
R66 VP.n69 VP.n68 24.4675
R67 VP.n74 VP.n73 24.4675
R68 VP.n40 VP.n39 24.4675
R69 VP.n32 VP.n13 24.4675
R70 VP.n35 VP.n34 24.4675
R71 VP.n22 VP.n15 24.4675
R72 VP.n26 VP.n15 24.4675
R73 VP.n27 VP.n26 24.4675
R74 VP.n28 VP.n27 24.4675
R75 VP.n21 VP.n20 24.4675
R76 VP.n54 VP.n7 20.5528
R77 VP.n67 VP.n66 20.5528
R78 VP.n33 VP.n32 20.5528
R79 VP.n20 VP.n17 20.5528
R80 VP.n45 VP.n44 16.6381
R81 VP.n75 VP.n74 16.6381
R82 VP.n41 VP.n40 16.6381
R83 VP.n19 VP.n18 9.28282
R84 VP.n51 VP.n7 3.91522
R85 VP.n68 VP.n67 3.91522
R86 VP.n34 VP.n33 3.91522
R87 VP.n42 VP.n10 0.278367
R88 VP.n46 VP.n43 0.278367
R89 VP.n76 VP.n0 0.278367
R90 VP.n19 VP.n16 0.189894
R91 VP.n23 VP.n16 0.189894
R92 VP.n24 VP.n23 0.189894
R93 VP.n25 VP.n24 0.189894
R94 VP.n25 VP.n14 0.189894
R95 VP.n29 VP.n14 0.189894
R96 VP.n30 VP.n29 0.189894
R97 VP.n31 VP.n30 0.189894
R98 VP.n31 VP.n12 0.189894
R99 VP.n36 VP.n12 0.189894
R100 VP.n37 VP.n36 0.189894
R101 VP.n38 VP.n37 0.189894
R102 VP.n38 VP.n10 0.189894
R103 VP.n47 VP.n46 0.189894
R104 VP.n48 VP.n47 0.189894
R105 VP.n48 VP.n8 0.189894
R106 VP.n52 VP.n8 0.189894
R107 VP.n53 VP.n52 0.189894
R108 VP.n53 VP.n6 0.189894
R109 VP.n57 VP.n6 0.189894
R110 VP.n58 VP.n57 0.189894
R111 VP.n59 VP.n58 0.189894
R112 VP.n59 VP.n4 0.189894
R113 VP.n63 VP.n4 0.189894
R114 VP.n64 VP.n63 0.189894
R115 VP.n65 VP.n64 0.189894
R116 VP.n65 VP.n2 0.189894
R117 VP.n70 VP.n2 0.189894
R118 VP.n71 VP.n70 0.189894
R119 VP.n72 VP.n71 0.189894
R120 VP.n72 VP.n0 0.189894
R121 VP VP.n76 0.153454
R122 VDD1.n1 VDD1.t7 152.388
R123 VDD1.n3 VDD1.t9 152.388
R124 VDD1.n5 VDD1.n4 140.161
R125 VDD1.n1 VDD1.n0 138.653
R126 VDD1.n7 VDD1.n6 138.651
R127 VDD1.n3 VDD1.n2 138.651
R128 VDD1.n7 VDD1.n5 37.6561
R129 VDD1.n6 VDD1.t4 11.651
R130 VDD1.n6 VDD1.t2 11.651
R131 VDD1.n0 VDD1.t6 11.651
R132 VDD1.n0 VDD1.t3 11.651
R133 VDD1.n4 VDD1.t5 11.651
R134 VDD1.n4 VDD1.t1 11.651
R135 VDD1.n2 VDD1.t8 11.651
R136 VDD1.n2 VDD1.t0 11.651
R137 VDD1 VDD1.n7 1.50697
R138 VDD1 VDD1.n1 0.580241
R139 VDD1.n5 VDD1.n3 0.466706
R140 VTAIL.n11 VTAIL.t6 133.624
R141 VTAIL.n17 VTAIL.t17 133.624
R142 VTAIL.n2 VTAIL.t9 133.624
R143 VTAIL.n16 VTAIL.t12 133.624
R144 VTAIL.n15 VTAIL.n14 121.974
R145 VTAIL.n13 VTAIL.n12 121.974
R146 VTAIL.n10 VTAIL.n9 121.974
R147 VTAIL.n8 VTAIL.n7 121.974
R148 VTAIL.n19 VTAIL.n18 121.972
R149 VTAIL.n1 VTAIL.n0 121.972
R150 VTAIL.n4 VTAIL.n3 121.972
R151 VTAIL.n6 VTAIL.n5 121.972
R152 VTAIL.n8 VTAIL.n6 18.9445
R153 VTAIL.n17 VTAIL.n16 16.8583
R154 VTAIL.n18 VTAIL.t1 11.651
R155 VTAIL.n18 VTAIL.t5 11.651
R156 VTAIL.n0 VTAIL.t0 11.651
R157 VTAIL.n0 VTAIL.t18 11.651
R158 VTAIL.n3 VTAIL.t11 11.651
R159 VTAIL.n3 VTAIL.t16 11.651
R160 VTAIL.n5 VTAIL.t7 11.651
R161 VTAIL.n5 VTAIL.t14 11.651
R162 VTAIL.n14 VTAIL.t10 11.651
R163 VTAIL.n14 VTAIL.t15 11.651
R164 VTAIL.n12 VTAIL.t13 11.651
R165 VTAIL.n12 VTAIL.t8 11.651
R166 VTAIL.n9 VTAIL.t2 11.651
R167 VTAIL.n9 VTAIL.t19 11.651
R168 VTAIL.n7 VTAIL.t3 11.651
R169 VTAIL.n7 VTAIL.t4 11.651
R170 VTAIL.n10 VTAIL.n8 2.08671
R171 VTAIL.n11 VTAIL.n10 2.08671
R172 VTAIL.n15 VTAIL.n13 2.08671
R173 VTAIL.n16 VTAIL.n15 2.08671
R174 VTAIL.n6 VTAIL.n4 2.08671
R175 VTAIL.n4 VTAIL.n2 2.08671
R176 VTAIL.n19 VTAIL.n17 2.08671
R177 VTAIL VTAIL.n1 1.62334
R178 VTAIL.n13 VTAIL.n11 1.51343
R179 VTAIL.n2 VTAIL.n1 1.51343
R180 VTAIL VTAIL.n19 0.463862
R181 B.n442 B.n441 585
R182 B.n443 B.n50 585
R183 B.n445 B.n444 585
R184 B.n446 B.n49 585
R185 B.n448 B.n447 585
R186 B.n449 B.n48 585
R187 B.n451 B.n450 585
R188 B.n452 B.n47 585
R189 B.n454 B.n453 585
R190 B.n455 B.n46 585
R191 B.n457 B.n456 585
R192 B.n458 B.n45 585
R193 B.n460 B.n459 585
R194 B.n461 B.n44 585
R195 B.n463 B.n462 585
R196 B.n465 B.n41 585
R197 B.n467 B.n466 585
R198 B.n468 B.n40 585
R199 B.n470 B.n469 585
R200 B.n471 B.n39 585
R201 B.n473 B.n472 585
R202 B.n474 B.n38 585
R203 B.n476 B.n475 585
R204 B.n477 B.n35 585
R205 B.n480 B.n479 585
R206 B.n481 B.n34 585
R207 B.n483 B.n482 585
R208 B.n484 B.n33 585
R209 B.n486 B.n485 585
R210 B.n487 B.n32 585
R211 B.n489 B.n488 585
R212 B.n490 B.n31 585
R213 B.n492 B.n491 585
R214 B.n493 B.n30 585
R215 B.n495 B.n494 585
R216 B.n496 B.n29 585
R217 B.n498 B.n497 585
R218 B.n499 B.n28 585
R219 B.n501 B.n500 585
R220 B.n440 B.n51 585
R221 B.n439 B.n438 585
R222 B.n437 B.n52 585
R223 B.n436 B.n435 585
R224 B.n434 B.n53 585
R225 B.n433 B.n432 585
R226 B.n431 B.n54 585
R227 B.n430 B.n429 585
R228 B.n428 B.n55 585
R229 B.n427 B.n426 585
R230 B.n425 B.n56 585
R231 B.n424 B.n423 585
R232 B.n422 B.n57 585
R233 B.n421 B.n420 585
R234 B.n419 B.n58 585
R235 B.n418 B.n417 585
R236 B.n416 B.n59 585
R237 B.n415 B.n414 585
R238 B.n413 B.n60 585
R239 B.n412 B.n411 585
R240 B.n410 B.n61 585
R241 B.n409 B.n408 585
R242 B.n407 B.n62 585
R243 B.n406 B.n405 585
R244 B.n404 B.n63 585
R245 B.n403 B.n402 585
R246 B.n401 B.n64 585
R247 B.n400 B.n399 585
R248 B.n398 B.n65 585
R249 B.n397 B.n396 585
R250 B.n395 B.n66 585
R251 B.n394 B.n393 585
R252 B.n392 B.n67 585
R253 B.n391 B.n390 585
R254 B.n389 B.n68 585
R255 B.n388 B.n387 585
R256 B.n386 B.n69 585
R257 B.n385 B.n384 585
R258 B.n383 B.n70 585
R259 B.n382 B.n381 585
R260 B.n380 B.n71 585
R261 B.n379 B.n378 585
R262 B.n377 B.n72 585
R263 B.n376 B.n375 585
R264 B.n374 B.n73 585
R265 B.n373 B.n372 585
R266 B.n371 B.n74 585
R267 B.n370 B.n369 585
R268 B.n368 B.n75 585
R269 B.n367 B.n366 585
R270 B.n365 B.n76 585
R271 B.n364 B.n363 585
R272 B.n362 B.n77 585
R273 B.n361 B.n360 585
R274 B.n359 B.n78 585
R275 B.n358 B.n357 585
R276 B.n356 B.n79 585
R277 B.n355 B.n354 585
R278 B.n353 B.n80 585
R279 B.n352 B.n351 585
R280 B.n350 B.n81 585
R281 B.n349 B.n348 585
R282 B.n347 B.n82 585
R283 B.n346 B.n345 585
R284 B.n344 B.n83 585
R285 B.n343 B.n342 585
R286 B.n341 B.n84 585
R287 B.n340 B.n339 585
R288 B.n338 B.n85 585
R289 B.n337 B.n336 585
R290 B.n335 B.n86 585
R291 B.n334 B.n333 585
R292 B.n332 B.n87 585
R293 B.n331 B.n330 585
R294 B.n329 B.n88 585
R295 B.n328 B.n327 585
R296 B.n326 B.n89 585
R297 B.n325 B.n324 585
R298 B.n323 B.n90 585
R299 B.n322 B.n321 585
R300 B.n320 B.n91 585
R301 B.n319 B.n318 585
R302 B.n317 B.n92 585
R303 B.n316 B.n315 585
R304 B.n314 B.n93 585
R305 B.n313 B.n312 585
R306 B.n311 B.n94 585
R307 B.n310 B.n309 585
R308 B.n308 B.n95 585
R309 B.n307 B.n306 585
R310 B.n305 B.n96 585
R311 B.n304 B.n303 585
R312 B.n302 B.n97 585
R313 B.n301 B.n300 585
R314 B.n299 B.n98 585
R315 B.n298 B.n297 585
R316 B.n296 B.n99 585
R317 B.n295 B.n294 585
R318 B.n293 B.n100 585
R319 B.n292 B.n291 585
R320 B.n290 B.n101 585
R321 B.n289 B.n288 585
R322 B.n287 B.n102 585
R323 B.n227 B.n126 585
R324 B.n229 B.n228 585
R325 B.n230 B.n125 585
R326 B.n232 B.n231 585
R327 B.n233 B.n124 585
R328 B.n235 B.n234 585
R329 B.n236 B.n123 585
R330 B.n238 B.n237 585
R331 B.n239 B.n122 585
R332 B.n241 B.n240 585
R333 B.n242 B.n121 585
R334 B.n244 B.n243 585
R335 B.n245 B.n120 585
R336 B.n247 B.n246 585
R337 B.n248 B.n117 585
R338 B.n251 B.n250 585
R339 B.n252 B.n116 585
R340 B.n254 B.n253 585
R341 B.n255 B.n115 585
R342 B.n257 B.n256 585
R343 B.n258 B.n114 585
R344 B.n260 B.n259 585
R345 B.n261 B.n113 585
R346 B.n263 B.n262 585
R347 B.n265 B.n264 585
R348 B.n266 B.n109 585
R349 B.n268 B.n267 585
R350 B.n269 B.n108 585
R351 B.n271 B.n270 585
R352 B.n272 B.n107 585
R353 B.n274 B.n273 585
R354 B.n275 B.n106 585
R355 B.n277 B.n276 585
R356 B.n278 B.n105 585
R357 B.n280 B.n279 585
R358 B.n281 B.n104 585
R359 B.n283 B.n282 585
R360 B.n284 B.n103 585
R361 B.n286 B.n285 585
R362 B.n226 B.n225 585
R363 B.n224 B.n127 585
R364 B.n223 B.n222 585
R365 B.n221 B.n128 585
R366 B.n220 B.n219 585
R367 B.n218 B.n129 585
R368 B.n217 B.n216 585
R369 B.n215 B.n130 585
R370 B.n214 B.n213 585
R371 B.n212 B.n131 585
R372 B.n211 B.n210 585
R373 B.n209 B.n132 585
R374 B.n208 B.n207 585
R375 B.n206 B.n133 585
R376 B.n205 B.n204 585
R377 B.n203 B.n134 585
R378 B.n202 B.n201 585
R379 B.n200 B.n135 585
R380 B.n199 B.n198 585
R381 B.n197 B.n136 585
R382 B.n196 B.n195 585
R383 B.n194 B.n137 585
R384 B.n193 B.n192 585
R385 B.n191 B.n138 585
R386 B.n190 B.n189 585
R387 B.n188 B.n139 585
R388 B.n187 B.n186 585
R389 B.n185 B.n140 585
R390 B.n184 B.n183 585
R391 B.n182 B.n141 585
R392 B.n181 B.n180 585
R393 B.n179 B.n142 585
R394 B.n178 B.n177 585
R395 B.n176 B.n143 585
R396 B.n175 B.n174 585
R397 B.n173 B.n144 585
R398 B.n172 B.n171 585
R399 B.n170 B.n145 585
R400 B.n169 B.n168 585
R401 B.n167 B.n146 585
R402 B.n166 B.n165 585
R403 B.n164 B.n147 585
R404 B.n163 B.n162 585
R405 B.n161 B.n148 585
R406 B.n160 B.n159 585
R407 B.n158 B.n149 585
R408 B.n157 B.n156 585
R409 B.n155 B.n150 585
R410 B.n154 B.n153 585
R411 B.n152 B.n151 585
R412 B.n2 B.n0 585
R413 B.n577 B.n1 585
R414 B.n576 B.n575 585
R415 B.n574 B.n3 585
R416 B.n573 B.n572 585
R417 B.n571 B.n4 585
R418 B.n570 B.n569 585
R419 B.n568 B.n5 585
R420 B.n567 B.n566 585
R421 B.n565 B.n6 585
R422 B.n564 B.n563 585
R423 B.n562 B.n7 585
R424 B.n561 B.n560 585
R425 B.n559 B.n8 585
R426 B.n558 B.n557 585
R427 B.n556 B.n9 585
R428 B.n555 B.n554 585
R429 B.n553 B.n10 585
R430 B.n552 B.n551 585
R431 B.n550 B.n11 585
R432 B.n549 B.n548 585
R433 B.n547 B.n12 585
R434 B.n546 B.n545 585
R435 B.n544 B.n13 585
R436 B.n543 B.n542 585
R437 B.n541 B.n14 585
R438 B.n540 B.n539 585
R439 B.n538 B.n15 585
R440 B.n537 B.n536 585
R441 B.n535 B.n16 585
R442 B.n534 B.n533 585
R443 B.n532 B.n17 585
R444 B.n531 B.n530 585
R445 B.n529 B.n18 585
R446 B.n528 B.n527 585
R447 B.n526 B.n19 585
R448 B.n525 B.n524 585
R449 B.n523 B.n20 585
R450 B.n522 B.n521 585
R451 B.n520 B.n21 585
R452 B.n519 B.n518 585
R453 B.n517 B.n22 585
R454 B.n516 B.n515 585
R455 B.n514 B.n23 585
R456 B.n513 B.n512 585
R457 B.n511 B.n24 585
R458 B.n510 B.n509 585
R459 B.n508 B.n25 585
R460 B.n507 B.n506 585
R461 B.n505 B.n26 585
R462 B.n504 B.n503 585
R463 B.n502 B.n27 585
R464 B.n579 B.n578 585
R465 B.n227 B.n226 439.647
R466 B.n500 B.n27 439.647
R467 B.n287 B.n286 439.647
R468 B.n442 B.n51 439.647
R469 B.n110 B.t0 239.293
R470 B.n118 B.t9 239.293
R471 B.n36 B.t3 239.293
R472 B.n42 B.t6 239.293
R473 B.n110 B.t2 188.899
R474 B.n42 B.t7 188.899
R475 B.n118 B.t11 188.898
R476 B.n36 B.t4 188.898
R477 B.n226 B.n127 163.367
R478 B.n222 B.n127 163.367
R479 B.n222 B.n221 163.367
R480 B.n221 B.n220 163.367
R481 B.n220 B.n129 163.367
R482 B.n216 B.n129 163.367
R483 B.n216 B.n215 163.367
R484 B.n215 B.n214 163.367
R485 B.n214 B.n131 163.367
R486 B.n210 B.n131 163.367
R487 B.n210 B.n209 163.367
R488 B.n209 B.n208 163.367
R489 B.n208 B.n133 163.367
R490 B.n204 B.n133 163.367
R491 B.n204 B.n203 163.367
R492 B.n203 B.n202 163.367
R493 B.n202 B.n135 163.367
R494 B.n198 B.n135 163.367
R495 B.n198 B.n197 163.367
R496 B.n197 B.n196 163.367
R497 B.n196 B.n137 163.367
R498 B.n192 B.n137 163.367
R499 B.n192 B.n191 163.367
R500 B.n191 B.n190 163.367
R501 B.n190 B.n139 163.367
R502 B.n186 B.n139 163.367
R503 B.n186 B.n185 163.367
R504 B.n185 B.n184 163.367
R505 B.n184 B.n141 163.367
R506 B.n180 B.n141 163.367
R507 B.n180 B.n179 163.367
R508 B.n179 B.n178 163.367
R509 B.n178 B.n143 163.367
R510 B.n174 B.n143 163.367
R511 B.n174 B.n173 163.367
R512 B.n173 B.n172 163.367
R513 B.n172 B.n145 163.367
R514 B.n168 B.n145 163.367
R515 B.n168 B.n167 163.367
R516 B.n167 B.n166 163.367
R517 B.n166 B.n147 163.367
R518 B.n162 B.n147 163.367
R519 B.n162 B.n161 163.367
R520 B.n161 B.n160 163.367
R521 B.n160 B.n149 163.367
R522 B.n156 B.n149 163.367
R523 B.n156 B.n155 163.367
R524 B.n155 B.n154 163.367
R525 B.n154 B.n151 163.367
R526 B.n151 B.n2 163.367
R527 B.n578 B.n2 163.367
R528 B.n578 B.n577 163.367
R529 B.n577 B.n576 163.367
R530 B.n576 B.n3 163.367
R531 B.n572 B.n3 163.367
R532 B.n572 B.n571 163.367
R533 B.n571 B.n570 163.367
R534 B.n570 B.n5 163.367
R535 B.n566 B.n5 163.367
R536 B.n566 B.n565 163.367
R537 B.n565 B.n564 163.367
R538 B.n564 B.n7 163.367
R539 B.n560 B.n7 163.367
R540 B.n560 B.n559 163.367
R541 B.n559 B.n558 163.367
R542 B.n558 B.n9 163.367
R543 B.n554 B.n9 163.367
R544 B.n554 B.n553 163.367
R545 B.n553 B.n552 163.367
R546 B.n552 B.n11 163.367
R547 B.n548 B.n11 163.367
R548 B.n548 B.n547 163.367
R549 B.n547 B.n546 163.367
R550 B.n546 B.n13 163.367
R551 B.n542 B.n13 163.367
R552 B.n542 B.n541 163.367
R553 B.n541 B.n540 163.367
R554 B.n540 B.n15 163.367
R555 B.n536 B.n15 163.367
R556 B.n536 B.n535 163.367
R557 B.n535 B.n534 163.367
R558 B.n534 B.n17 163.367
R559 B.n530 B.n17 163.367
R560 B.n530 B.n529 163.367
R561 B.n529 B.n528 163.367
R562 B.n528 B.n19 163.367
R563 B.n524 B.n19 163.367
R564 B.n524 B.n523 163.367
R565 B.n523 B.n522 163.367
R566 B.n522 B.n21 163.367
R567 B.n518 B.n21 163.367
R568 B.n518 B.n517 163.367
R569 B.n517 B.n516 163.367
R570 B.n516 B.n23 163.367
R571 B.n512 B.n23 163.367
R572 B.n512 B.n511 163.367
R573 B.n511 B.n510 163.367
R574 B.n510 B.n25 163.367
R575 B.n506 B.n25 163.367
R576 B.n506 B.n505 163.367
R577 B.n505 B.n504 163.367
R578 B.n504 B.n27 163.367
R579 B.n228 B.n227 163.367
R580 B.n228 B.n125 163.367
R581 B.n232 B.n125 163.367
R582 B.n233 B.n232 163.367
R583 B.n234 B.n233 163.367
R584 B.n234 B.n123 163.367
R585 B.n238 B.n123 163.367
R586 B.n239 B.n238 163.367
R587 B.n240 B.n239 163.367
R588 B.n240 B.n121 163.367
R589 B.n244 B.n121 163.367
R590 B.n245 B.n244 163.367
R591 B.n246 B.n245 163.367
R592 B.n246 B.n117 163.367
R593 B.n251 B.n117 163.367
R594 B.n252 B.n251 163.367
R595 B.n253 B.n252 163.367
R596 B.n253 B.n115 163.367
R597 B.n257 B.n115 163.367
R598 B.n258 B.n257 163.367
R599 B.n259 B.n258 163.367
R600 B.n259 B.n113 163.367
R601 B.n263 B.n113 163.367
R602 B.n264 B.n263 163.367
R603 B.n264 B.n109 163.367
R604 B.n268 B.n109 163.367
R605 B.n269 B.n268 163.367
R606 B.n270 B.n269 163.367
R607 B.n270 B.n107 163.367
R608 B.n274 B.n107 163.367
R609 B.n275 B.n274 163.367
R610 B.n276 B.n275 163.367
R611 B.n276 B.n105 163.367
R612 B.n280 B.n105 163.367
R613 B.n281 B.n280 163.367
R614 B.n282 B.n281 163.367
R615 B.n282 B.n103 163.367
R616 B.n286 B.n103 163.367
R617 B.n288 B.n287 163.367
R618 B.n288 B.n101 163.367
R619 B.n292 B.n101 163.367
R620 B.n293 B.n292 163.367
R621 B.n294 B.n293 163.367
R622 B.n294 B.n99 163.367
R623 B.n298 B.n99 163.367
R624 B.n299 B.n298 163.367
R625 B.n300 B.n299 163.367
R626 B.n300 B.n97 163.367
R627 B.n304 B.n97 163.367
R628 B.n305 B.n304 163.367
R629 B.n306 B.n305 163.367
R630 B.n306 B.n95 163.367
R631 B.n310 B.n95 163.367
R632 B.n311 B.n310 163.367
R633 B.n312 B.n311 163.367
R634 B.n312 B.n93 163.367
R635 B.n316 B.n93 163.367
R636 B.n317 B.n316 163.367
R637 B.n318 B.n317 163.367
R638 B.n318 B.n91 163.367
R639 B.n322 B.n91 163.367
R640 B.n323 B.n322 163.367
R641 B.n324 B.n323 163.367
R642 B.n324 B.n89 163.367
R643 B.n328 B.n89 163.367
R644 B.n329 B.n328 163.367
R645 B.n330 B.n329 163.367
R646 B.n330 B.n87 163.367
R647 B.n334 B.n87 163.367
R648 B.n335 B.n334 163.367
R649 B.n336 B.n335 163.367
R650 B.n336 B.n85 163.367
R651 B.n340 B.n85 163.367
R652 B.n341 B.n340 163.367
R653 B.n342 B.n341 163.367
R654 B.n342 B.n83 163.367
R655 B.n346 B.n83 163.367
R656 B.n347 B.n346 163.367
R657 B.n348 B.n347 163.367
R658 B.n348 B.n81 163.367
R659 B.n352 B.n81 163.367
R660 B.n353 B.n352 163.367
R661 B.n354 B.n353 163.367
R662 B.n354 B.n79 163.367
R663 B.n358 B.n79 163.367
R664 B.n359 B.n358 163.367
R665 B.n360 B.n359 163.367
R666 B.n360 B.n77 163.367
R667 B.n364 B.n77 163.367
R668 B.n365 B.n364 163.367
R669 B.n366 B.n365 163.367
R670 B.n366 B.n75 163.367
R671 B.n370 B.n75 163.367
R672 B.n371 B.n370 163.367
R673 B.n372 B.n371 163.367
R674 B.n372 B.n73 163.367
R675 B.n376 B.n73 163.367
R676 B.n377 B.n376 163.367
R677 B.n378 B.n377 163.367
R678 B.n378 B.n71 163.367
R679 B.n382 B.n71 163.367
R680 B.n383 B.n382 163.367
R681 B.n384 B.n383 163.367
R682 B.n384 B.n69 163.367
R683 B.n388 B.n69 163.367
R684 B.n389 B.n388 163.367
R685 B.n390 B.n389 163.367
R686 B.n390 B.n67 163.367
R687 B.n394 B.n67 163.367
R688 B.n395 B.n394 163.367
R689 B.n396 B.n395 163.367
R690 B.n396 B.n65 163.367
R691 B.n400 B.n65 163.367
R692 B.n401 B.n400 163.367
R693 B.n402 B.n401 163.367
R694 B.n402 B.n63 163.367
R695 B.n406 B.n63 163.367
R696 B.n407 B.n406 163.367
R697 B.n408 B.n407 163.367
R698 B.n408 B.n61 163.367
R699 B.n412 B.n61 163.367
R700 B.n413 B.n412 163.367
R701 B.n414 B.n413 163.367
R702 B.n414 B.n59 163.367
R703 B.n418 B.n59 163.367
R704 B.n419 B.n418 163.367
R705 B.n420 B.n419 163.367
R706 B.n420 B.n57 163.367
R707 B.n424 B.n57 163.367
R708 B.n425 B.n424 163.367
R709 B.n426 B.n425 163.367
R710 B.n426 B.n55 163.367
R711 B.n430 B.n55 163.367
R712 B.n431 B.n430 163.367
R713 B.n432 B.n431 163.367
R714 B.n432 B.n53 163.367
R715 B.n436 B.n53 163.367
R716 B.n437 B.n436 163.367
R717 B.n438 B.n437 163.367
R718 B.n438 B.n51 163.367
R719 B.n500 B.n499 163.367
R720 B.n499 B.n498 163.367
R721 B.n498 B.n29 163.367
R722 B.n494 B.n29 163.367
R723 B.n494 B.n493 163.367
R724 B.n493 B.n492 163.367
R725 B.n492 B.n31 163.367
R726 B.n488 B.n31 163.367
R727 B.n488 B.n487 163.367
R728 B.n487 B.n486 163.367
R729 B.n486 B.n33 163.367
R730 B.n482 B.n33 163.367
R731 B.n482 B.n481 163.367
R732 B.n481 B.n480 163.367
R733 B.n480 B.n35 163.367
R734 B.n475 B.n35 163.367
R735 B.n475 B.n474 163.367
R736 B.n474 B.n473 163.367
R737 B.n473 B.n39 163.367
R738 B.n469 B.n39 163.367
R739 B.n469 B.n468 163.367
R740 B.n468 B.n467 163.367
R741 B.n467 B.n41 163.367
R742 B.n462 B.n41 163.367
R743 B.n462 B.n461 163.367
R744 B.n461 B.n460 163.367
R745 B.n460 B.n45 163.367
R746 B.n456 B.n45 163.367
R747 B.n456 B.n455 163.367
R748 B.n455 B.n454 163.367
R749 B.n454 B.n47 163.367
R750 B.n450 B.n47 163.367
R751 B.n450 B.n449 163.367
R752 B.n449 B.n448 163.367
R753 B.n448 B.n49 163.367
R754 B.n444 B.n49 163.367
R755 B.n444 B.n443 163.367
R756 B.n443 B.n442 163.367
R757 B.n111 B.t1 141.965
R758 B.n43 B.t8 141.965
R759 B.n119 B.t10 141.964
R760 B.n37 B.t5 141.964
R761 B.n112 B.n111 59.5399
R762 B.n249 B.n119 59.5399
R763 B.n478 B.n37 59.5399
R764 B.n464 B.n43 59.5399
R765 B.n111 B.n110 46.9338
R766 B.n119 B.n118 46.9338
R767 B.n37 B.n36 46.9338
R768 B.n43 B.n42 46.9338
R769 B.n502 B.n501 28.5664
R770 B.n285 B.n102 28.5664
R771 B.n225 B.n126 28.5664
R772 B.n441 B.n440 28.5664
R773 B B.n579 18.0485
R774 B.n501 B.n28 10.6151
R775 B.n497 B.n28 10.6151
R776 B.n497 B.n496 10.6151
R777 B.n496 B.n495 10.6151
R778 B.n495 B.n30 10.6151
R779 B.n491 B.n30 10.6151
R780 B.n491 B.n490 10.6151
R781 B.n490 B.n489 10.6151
R782 B.n489 B.n32 10.6151
R783 B.n485 B.n32 10.6151
R784 B.n485 B.n484 10.6151
R785 B.n484 B.n483 10.6151
R786 B.n483 B.n34 10.6151
R787 B.n479 B.n34 10.6151
R788 B.n477 B.n476 10.6151
R789 B.n476 B.n38 10.6151
R790 B.n472 B.n38 10.6151
R791 B.n472 B.n471 10.6151
R792 B.n471 B.n470 10.6151
R793 B.n470 B.n40 10.6151
R794 B.n466 B.n40 10.6151
R795 B.n466 B.n465 10.6151
R796 B.n463 B.n44 10.6151
R797 B.n459 B.n44 10.6151
R798 B.n459 B.n458 10.6151
R799 B.n458 B.n457 10.6151
R800 B.n457 B.n46 10.6151
R801 B.n453 B.n46 10.6151
R802 B.n453 B.n452 10.6151
R803 B.n452 B.n451 10.6151
R804 B.n451 B.n48 10.6151
R805 B.n447 B.n48 10.6151
R806 B.n447 B.n446 10.6151
R807 B.n446 B.n445 10.6151
R808 B.n445 B.n50 10.6151
R809 B.n441 B.n50 10.6151
R810 B.n289 B.n102 10.6151
R811 B.n290 B.n289 10.6151
R812 B.n291 B.n290 10.6151
R813 B.n291 B.n100 10.6151
R814 B.n295 B.n100 10.6151
R815 B.n296 B.n295 10.6151
R816 B.n297 B.n296 10.6151
R817 B.n297 B.n98 10.6151
R818 B.n301 B.n98 10.6151
R819 B.n302 B.n301 10.6151
R820 B.n303 B.n302 10.6151
R821 B.n303 B.n96 10.6151
R822 B.n307 B.n96 10.6151
R823 B.n308 B.n307 10.6151
R824 B.n309 B.n308 10.6151
R825 B.n309 B.n94 10.6151
R826 B.n313 B.n94 10.6151
R827 B.n314 B.n313 10.6151
R828 B.n315 B.n314 10.6151
R829 B.n315 B.n92 10.6151
R830 B.n319 B.n92 10.6151
R831 B.n320 B.n319 10.6151
R832 B.n321 B.n320 10.6151
R833 B.n321 B.n90 10.6151
R834 B.n325 B.n90 10.6151
R835 B.n326 B.n325 10.6151
R836 B.n327 B.n326 10.6151
R837 B.n327 B.n88 10.6151
R838 B.n331 B.n88 10.6151
R839 B.n332 B.n331 10.6151
R840 B.n333 B.n332 10.6151
R841 B.n333 B.n86 10.6151
R842 B.n337 B.n86 10.6151
R843 B.n338 B.n337 10.6151
R844 B.n339 B.n338 10.6151
R845 B.n339 B.n84 10.6151
R846 B.n343 B.n84 10.6151
R847 B.n344 B.n343 10.6151
R848 B.n345 B.n344 10.6151
R849 B.n345 B.n82 10.6151
R850 B.n349 B.n82 10.6151
R851 B.n350 B.n349 10.6151
R852 B.n351 B.n350 10.6151
R853 B.n351 B.n80 10.6151
R854 B.n355 B.n80 10.6151
R855 B.n356 B.n355 10.6151
R856 B.n357 B.n356 10.6151
R857 B.n357 B.n78 10.6151
R858 B.n361 B.n78 10.6151
R859 B.n362 B.n361 10.6151
R860 B.n363 B.n362 10.6151
R861 B.n363 B.n76 10.6151
R862 B.n367 B.n76 10.6151
R863 B.n368 B.n367 10.6151
R864 B.n369 B.n368 10.6151
R865 B.n369 B.n74 10.6151
R866 B.n373 B.n74 10.6151
R867 B.n374 B.n373 10.6151
R868 B.n375 B.n374 10.6151
R869 B.n375 B.n72 10.6151
R870 B.n379 B.n72 10.6151
R871 B.n380 B.n379 10.6151
R872 B.n381 B.n380 10.6151
R873 B.n381 B.n70 10.6151
R874 B.n385 B.n70 10.6151
R875 B.n386 B.n385 10.6151
R876 B.n387 B.n386 10.6151
R877 B.n387 B.n68 10.6151
R878 B.n391 B.n68 10.6151
R879 B.n392 B.n391 10.6151
R880 B.n393 B.n392 10.6151
R881 B.n393 B.n66 10.6151
R882 B.n397 B.n66 10.6151
R883 B.n398 B.n397 10.6151
R884 B.n399 B.n398 10.6151
R885 B.n399 B.n64 10.6151
R886 B.n403 B.n64 10.6151
R887 B.n404 B.n403 10.6151
R888 B.n405 B.n404 10.6151
R889 B.n405 B.n62 10.6151
R890 B.n409 B.n62 10.6151
R891 B.n410 B.n409 10.6151
R892 B.n411 B.n410 10.6151
R893 B.n411 B.n60 10.6151
R894 B.n415 B.n60 10.6151
R895 B.n416 B.n415 10.6151
R896 B.n417 B.n416 10.6151
R897 B.n417 B.n58 10.6151
R898 B.n421 B.n58 10.6151
R899 B.n422 B.n421 10.6151
R900 B.n423 B.n422 10.6151
R901 B.n423 B.n56 10.6151
R902 B.n427 B.n56 10.6151
R903 B.n428 B.n427 10.6151
R904 B.n429 B.n428 10.6151
R905 B.n429 B.n54 10.6151
R906 B.n433 B.n54 10.6151
R907 B.n434 B.n433 10.6151
R908 B.n435 B.n434 10.6151
R909 B.n435 B.n52 10.6151
R910 B.n439 B.n52 10.6151
R911 B.n440 B.n439 10.6151
R912 B.n229 B.n126 10.6151
R913 B.n230 B.n229 10.6151
R914 B.n231 B.n230 10.6151
R915 B.n231 B.n124 10.6151
R916 B.n235 B.n124 10.6151
R917 B.n236 B.n235 10.6151
R918 B.n237 B.n236 10.6151
R919 B.n237 B.n122 10.6151
R920 B.n241 B.n122 10.6151
R921 B.n242 B.n241 10.6151
R922 B.n243 B.n242 10.6151
R923 B.n243 B.n120 10.6151
R924 B.n247 B.n120 10.6151
R925 B.n248 B.n247 10.6151
R926 B.n250 B.n116 10.6151
R927 B.n254 B.n116 10.6151
R928 B.n255 B.n254 10.6151
R929 B.n256 B.n255 10.6151
R930 B.n256 B.n114 10.6151
R931 B.n260 B.n114 10.6151
R932 B.n261 B.n260 10.6151
R933 B.n262 B.n261 10.6151
R934 B.n266 B.n265 10.6151
R935 B.n267 B.n266 10.6151
R936 B.n267 B.n108 10.6151
R937 B.n271 B.n108 10.6151
R938 B.n272 B.n271 10.6151
R939 B.n273 B.n272 10.6151
R940 B.n273 B.n106 10.6151
R941 B.n277 B.n106 10.6151
R942 B.n278 B.n277 10.6151
R943 B.n279 B.n278 10.6151
R944 B.n279 B.n104 10.6151
R945 B.n283 B.n104 10.6151
R946 B.n284 B.n283 10.6151
R947 B.n285 B.n284 10.6151
R948 B.n225 B.n224 10.6151
R949 B.n224 B.n223 10.6151
R950 B.n223 B.n128 10.6151
R951 B.n219 B.n128 10.6151
R952 B.n219 B.n218 10.6151
R953 B.n218 B.n217 10.6151
R954 B.n217 B.n130 10.6151
R955 B.n213 B.n130 10.6151
R956 B.n213 B.n212 10.6151
R957 B.n212 B.n211 10.6151
R958 B.n211 B.n132 10.6151
R959 B.n207 B.n132 10.6151
R960 B.n207 B.n206 10.6151
R961 B.n206 B.n205 10.6151
R962 B.n205 B.n134 10.6151
R963 B.n201 B.n134 10.6151
R964 B.n201 B.n200 10.6151
R965 B.n200 B.n199 10.6151
R966 B.n199 B.n136 10.6151
R967 B.n195 B.n136 10.6151
R968 B.n195 B.n194 10.6151
R969 B.n194 B.n193 10.6151
R970 B.n193 B.n138 10.6151
R971 B.n189 B.n138 10.6151
R972 B.n189 B.n188 10.6151
R973 B.n188 B.n187 10.6151
R974 B.n187 B.n140 10.6151
R975 B.n183 B.n140 10.6151
R976 B.n183 B.n182 10.6151
R977 B.n182 B.n181 10.6151
R978 B.n181 B.n142 10.6151
R979 B.n177 B.n142 10.6151
R980 B.n177 B.n176 10.6151
R981 B.n176 B.n175 10.6151
R982 B.n175 B.n144 10.6151
R983 B.n171 B.n144 10.6151
R984 B.n171 B.n170 10.6151
R985 B.n170 B.n169 10.6151
R986 B.n169 B.n146 10.6151
R987 B.n165 B.n146 10.6151
R988 B.n165 B.n164 10.6151
R989 B.n164 B.n163 10.6151
R990 B.n163 B.n148 10.6151
R991 B.n159 B.n148 10.6151
R992 B.n159 B.n158 10.6151
R993 B.n158 B.n157 10.6151
R994 B.n157 B.n150 10.6151
R995 B.n153 B.n150 10.6151
R996 B.n153 B.n152 10.6151
R997 B.n152 B.n0 10.6151
R998 B.n575 B.n1 10.6151
R999 B.n575 B.n574 10.6151
R1000 B.n574 B.n573 10.6151
R1001 B.n573 B.n4 10.6151
R1002 B.n569 B.n4 10.6151
R1003 B.n569 B.n568 10.6151
R1004 B.n568 B.n567 10.6151
R1005 B.n567 B.n6 10.6151
R1006 B.n563 B.n6 10.6151
R1007 B.n563 B.n562 10.6151
R1008 B.n562 B.n561 10.6151
R1009 B.n561 B.n8 10.6151
R1010 B.n557 B.n8 10.6151
R1011 B.n557 B.n556 10.6151
R1012 B.n556 B.n555 10.6151
R1013 B.n555 B.n10 10.6151
R1014 B.n551 B.n10 10.6151
R1015 B.n551 B.n550 10.6151
R1016 B.n550 B.n549 10.6151
R1017 B.n549 B.n12 10.6151
R1018 B.n545 B.n12 10.6151
R1019 B.n545 B.n544 10.6151
R1020 B.n544 B.n543 10.6151
R1021 B.n543 B.n14 10.6151
R1022 B.n539 B.n14 10.6151
R1023 B.n539 B.n538 10.6151
R1024 B.n538 B.n537 10.6151
R1025 B.n537 B.n16 10.6151
R1026 B.n533 B.n16 10.6151
R1027 B.n533 B.n532 10.6151
R1028 B.n532 B.n531 10.6151
R1029 B.n531 B.n18 10.6151
R1030 B.n527 B.n18 10.6151
R1031 B.n527 B.n526 10.6151
R1032 B.n526 B.n525 10.6151
R1033 B.n525 B.n20 10.6151
R1034 B.n521 B.n20 10.6151
R1035 B.n521 B.n520 10.6151
R1036 B.n520 B.n519 10.6151
R1037 B.n519 B.n22 10.6151
R1038 B.n515 B.n22 10.6151
R1039 B.n515 B.n514 10.6151
R1040 B.n514 B.n513 10.6151
R1041 B.n513 B.n24 10.6151
R1042 B.n509 B.n24 10.6151
R1043 B.n509 B.n508 10.6151
R1044 B.n508 B.n507 10.6151
R1045 B.n507 B.n26 10.6151
R1046 B.n503 B.n26 10.6151
R1047 B.n503 B.n502 10.6151
R1048 B.n478 B.n477 6.5566
R1049 B.n465 B.n464 6.5566
R1050 B.n250 B.n249 6.5566
R1051 B.n262 B.n112 6.5566
R1052 B.n479 B.n478 4.05904
R1053 B.n464 B.n463 4.05904
R1054 B.n249 B.n248 4.05904
R1055 B.n265 B.n112 4.05904
R1056 B.n579 B.n0 2.81026
R1057 B.n579 B.n1 2.81026
R1058 VN.n63 VN.n33 161.3
R1059 VN.n62 VN.n61 161.3
R1060 VN.n60 VN.n34 161.3
R1061 VN.n59 VN.n58 161.3
R1062 VN.n57 VN.n35 161.3
R1063 VN.n55 VN.n54 161.3
R1064 VN.n53 VN.n36 161.3
R1065 VN.n52 VN.n51 161.3
R1066 VN.n50 VN.n37 161.3
R1067 VN.n49 VN.n48 161.3
R1068 VN.n47 VN.n38 161.3
R1069 VN.n46 VN.n45 161.3
R1070 VN.n44 VN.n39 161.3
R1071 VN.n43 VN.n42 161.3
R1072 VN.n30 VN.n0 161.3
R1073 VN.n29 VN.n28 161.3
R1074 VN.n27 VN.n1 161.3
R1075 VN.n26 VN.n25 161.3
R1076 VN.n24 VN.n2 161.3
R1077 VN.n22 VN.n21 161.3
R1078 VN.n20 VN.n3 161.3
R1079 VN.n19 VN.n18 161.3
R1080 VN.n17 VN.n4 161.3
R1081 VN.n16 VN.n15 161.3
R1082 VN.n14 VN.n5 161.3
R1083 VN.n13 VN.n12 161.3
R1084 VN.n11 VN.n6 161.3
R1085 VN.n10 VN.n9 161.3
R1086 VN.n32 VN.n31 94.1189
R1087 VN.n65 VN.n64 94.1189
R1088 VN.n8 VN.t6 65.6206
R1089 VN.n41 VN.t3 65.6206
R1090 VN.n12 VN.n11 56.5193
R1091 VN.n18 VN.n3 56.5193
R1092 VN.n45 VN.n44 56.5193
R1093 VN.n51 VN.n36 56.5193
R1094 VN.n29 VN.n1 53.1199
R1095 VN.n62 VN.n34 53.1199
R1096 VN.n8 VN.n7 50.0611
R1097 VN.n41 VN.n40 50.0611
R1098 VN VN.n65 43.6421
R1099 VN.n16 VN.t7 32.1723
R1100 VN.n7 VN.t2 32.1723
R1101 VN.n23 VN.t5 32.1723
R1102 VN.n31 VN.t0 32.1723
R1103 VN.n49 VN.t9 32.1723
R1104 VN.n40 VN.t1 32.1723
R1105 VN.n56 VN.t4 32.1723
R1106 VN.n64 VN.t8 32.1723
R1107 VN.n25 VN.n1 27.8669
R1108 VN.n58 VN.n34 27.8669
R1109 VN.n11 VN.n10 24.4675
R1110 VN.n12 VN.n5 24.4675
R1111 VN.n16 VN.n5 24.4675
R1112 VN.n17 VN.n16 24.4675
R1113 VN.n18 VN.n17 24.4675
R1114 VN.n22 VN.n3 24.4675
R1115 VN.n25 VN.n24 24.4675
R1116 VN.n30 VN.n29 24.4675
R1117 VN.n44 VN.n43 24.4675
R1118 VN.n51 VN.n50 24.4675
R1119 VN.n50 VN.n49 24.4675
R1120 VN.n49 VN.n38 24.4675
R1121 VN.n45 VN.n38 24.4675
R1122 VN.n58 VN.n57 24.4675
R1123 VN.n55 VN.n36 24.4675
R1124 VN.n63 VN.n62 24.4675
R1125 VN.n10 VN.n7 20.5528
R1126 VN.n23 VN.n22 20.5528
R1127 VN.n43 VN.n40 20.5528
R1128 VN.n56 VN.n55 20.5528
R1129 VN.n31 VN.n30 16.6381
R1130 VN.n64 VN.n63 16.6381
R1131 VN.n42 VN.n41 9.28282
R1132 VN.n9 VN.n8 9.28282
R1133 VN.n24 VN.n23 3.91522
R1134 VN.n57 VN.n56 3.91522
R1135 VN.n65 VN.n33 0.278367
R1136 VN.n32 VN.n0 0.278367
R1137 VN.n61 VN.n33 0.189894
R1138 VN.n61 VN.n60 0.189894
R1139 VN.n60 VN.n59 0.189894
R1140 VN.n59 VN.n35 0.189894
R1141 VN.n54 VN.n35 0.189894
R1142 VN.n54 VN.n53 0.189894
R1143 VN.n53 VN.n52 0.189894
R1144 VN.n52 VN.n37 0.189894
R1145 VN.n48 VN.n37 0.189894
R1146 VN.n48 VN.n47 0.189894
R1147 VN.n47 VN.n46 0.189894
R1148 VN.n46 VN.n39 0.189894
R1149 VN.n42 VN.n39 0.189894
R1150 VN.n9 VN.n6 0.189894
R1151 VN.n13 VN.n6 0.189894
R1152 VN.n14 VN.n13 0.189894
R1153 VN.n15 VN.n14 0.189894
R1154 VN.n15 VN.n4 0.189894
R1155 VN.n19 VN.n4 0.189894
R1156 VN.n20 VN.n19 0.189894
R1157 VN.n21 VN.n20 0.189894
R1158 VN.n21 VN.n2 0.189894
R1159 VN.n26 VN.n2 0.189894
R1160 VN.n27 VN.n26 0.189894
R1161 VN.n28 VN.n27 0.189894
R1162 VN.n28 VN.n0 0.189894
R1163 VN VN.n32 0.153454
R1164 VDD2.n1 VDD2.t3 152.388
R1165 VDD2.n4 VDD2.t1 150.303
R1166 VDD2.n3 VDD2.n2 140.161
R1167 VDD2 VDD2.n7 140.159
R1168 VDD2.n6 VDD2.n5 138.653
R1169 VDD2.n1 VDD2.n0 138.651
R1170 VDD2.n4 VDD2.n3 36.03
R1171 VDD2.n7 VDD2.t8 11.651
R1172 VDD2.n7 VDD2.t6 11.651
R1173 VDD2.n5 VDD2.t5 11.651
R1174 VDD2.n5 VDD2.t0 11.651
R1175 VDD2.n2 VDD2.t4 11.651
R1176 VDD2.n2 VDD2.t9 11.651
R1177 VDD2.n0 VDD2.t7 11.651
R1178 VDD2.n0 VDD2.t2 11.651
R1179 VDD2.n6 VDD2.n4 2.08671
R1180 VDD2 VDD2.n6 0.580241
R1181 VDD2.n3 VDD2.n1 0.466706
C0 VDD2 VN 2.74706f
C1 w_n3874_n1526# VN 7.972471f
C2 VDD1 VTAIL 5.65942f
C3 VP VN 5.95022f
C4 B VN 1.06399f
C5 VDD2 VTAIL 5.70892f
C6 VDD2 VDD1 1.84184f
C7 w_n3874_n1526# VTAIL 1.80411f
C8 w_n3874_n1526# VDD1 1.94554f
C9 VP VTAIL 3.81863f
C10 VP VDD1 3.11035f
C11 B VTAIL 1.46915f
C12 B VDD1 1.56101f
C13 w_n3874_n1526# VDD2 2.06212f
C14 VDD2 VP 0.524082f
C15 VDD2 B 1.65926f
C16 w_n3874_n1526# VP 8.47259f
C17 w_n3874_n1526# B 7.13423f
C18 B VP 1.90618f
C19 VN VTAIL 3.80447f
C20 VN VDD1 0.157698f
C21 VDD2 VSUBS 1.506056f
C22 VDD1 VSUBS 1.430318f
C23 VTAIL VSUBS 0.510584f
C24 VN VSUBS 6.70373f
C25 VP VSUBS 3.001343f
C26 B VSUBS 3.712683f
C27 w_n3874_n1526# VSUBS 74.9851f
C28 VDD2.t3 VSUBS 0.470886f
C29 VDD2.t7 VSUBS 0.063205f
C30 VDD2.t2 VSUBS 0.063205f
C31 VDD2.n0 VSUBS 0.324036f
C32 VDD2.n1 VSUBS 1.16762f
C33 VDD2.t4 VSUBS 0.063205f
C34 VDD2.t9 VSUBS 0.063205f
C35 VDD2.n2 VSUBS 0.331514f
C36 VDD2.n3 VSUBS 2.51359f
C37 VDD2.t1 VSUBS 0.462835f
C38 VDD2.n4 VSUBS 2.59278f
C39 VDD2.t5 VSUBS 0.063205f
C40 VDD2.t0 VSUBS 0.063205f
C41 VDD2.n5 VSUBS 0.324037f
C42 VDD2.n6 VSUBS 0.59658f
C43 VDD2.t8 VSUBS 0.063205f
C44 VDD2.t6 VSUBS 0.063205f
C45 VDD2.n7 VSUBS 0.331492f
C46 VN.n0 VSUBS 0.065514f
C47 VN.t0 VSUBS 0.71502f
C48 VN.n1 VSUBS 0.052118f
C49 VN.n2 VSUBS 0.049692f
C50 VN.t5 VSUBS 0.71502f
C51 VN.n3 VSUBS 0.07808f
C52 VN.n4 VSUBS 0.049692f
C53 VN.t7 VSUBS 0.71502f
C54 VN.n5 VSUBS 0.092613f
C55 VN.n6 VSUBS 0.049692f
C56 VN.t2 VSUBS 0.71502f
C57 VN.n7 VSUBS 0.456038f
C58 VN.t6 VSUBS 1.00958f
C59 VN.n8 VSUBS 0.41878f
C60 VN.n9 VSUBS 0.417942f
C61 VN.n10 VSUBS 0.085297f
C62 VN.n11 VSUBS 0.07808f
C63 VN.n12 VSUBS 0.067002f
C64 VN.n13 VSUBS 0.049692f
C65 VN.n14 VSUBS 0.049692f
C66 VN.n15 VSUBS 0.049692f
C67 VN.n16 VSUBS 0.363292f
C68 VN.n17 VSUBS 0.092613f
C69 VN.n18 VSUBS 0.067002f
C70 VN.n19 VSUBS 0.049692f
C71 VN.n20 VSUBS 0.049692f
C72 VN.n21 VSUBS 0.049692f
C73 VN.n22 VSUBS 0.085297f
C74 VN.n23 VSUBS 0.316403f
C75 VN.n24 VSUBS 0.054205f
C76 VN.n25 VSUBS 0.097407f
C77 VN.n26 VSUBS 0.049692f
C78 VN.n27 VSUBS 0.049692f
C79 VN.n28 VSUBS 0.049692f
C80 VN.n29 VSUBS 0.08817f
C81 VN.n30 VSUBS 0.077982f
C82 VN.n31 VSUBS 0.466187f
C83 VN.n32 VSUBS 0.065501f
C84 VN.n33 VSUBS 0.065514f
C85 VN.t8 VSUBS 0.71502f
C86 VN.n34 VSUBS 0.052118f
C87 VN.n35 VSUBS 0.049692f
C88 VN.t4 VSUBS 0.71502f
C89 VN.n36 VSUBS 0.07808f
C90 VN.n37 VSUBS 0.049692f
C91 VN.t9 VSUBS 0.71502f
C92 VN.n38 VSUBS 0.092613f
C93 VN.n39 VSUBS 0.049692f
C94 VN.t1 VSUBS 0.71502f
C95 VN.n40 VSUBS 0.456038f
C96 VN.t3 VSUBS 1.00958f
C97 VN.n41 VSUBS 0.41878f
C98 VN.n42 VSUBS 0.417942f
C99 VN.n43 VSUBS 0.085297f
C100 VN.n44 VSUBS 0.07808f
C101 VN.n45 VSUBS 0.067002f
C102 VN.n46 VSUBS 0.049692f
C103 VN.n47 VSUBS 0.049692f
C104 VN.n48 VSUBS 0.049692f
C105 VN.n49 VSUBS 0.363292f
C106 VN.n50 VSUBS 0.092613f
C107 VN.n51 VSUBS 0.067002f
C108 VN.n52 VSUBS 0.049692f
C109 VN.n53 VSUBS 0.049692f
C110 VN.n54 VSUBS 0.049692f
C111 VN.n55 VSUBS 0.085297f
C112 VN.n56 VSUBS 0.316403f
C113 VN.n57 VSUBS 0.054205f
C114 VN.n58 VSUBS 0.097407f
C115 VN.n59 VSUBS 0.049692f
C116 VN.n60 VSUBS 0.049692f
C117 VN.n61 VSUBS 0.049692f
C118 VN.n62 VSUBS 0.08817f
C119 VN.n63 VSUBS 0.077982f
C120 VN.n64 VSUBS 0.466187f
C121 VN.n65 VSUBS 2.23585f
C122 B.n0 VSUBS 0.004893f
C123 B.n1 VSUBS 0.004893f
C124 B.n2 VSUBS 0.007737f
C125 B.n3 VSUBS 0.007737f
C126 B.n4 VSUBS 0.007737f
C127 B.n5 VSUBS 0.007737f
C128 B.n6 VSUBS 0.007737f
C129 B.n7 VSUBS 0.007737f
C130 B.n8 VSUBS 0.007737f
C131 B.n9 VSUBS 0.007737f
C132 B.n10 VSUBS 0.007737f
C133 B.n11 VSUBS 0.007737f
C134 B.n12 VSUBS 0.007737f
C135 B.n13 VSUBS 0.007737f
C136 B.n14 VSUBS 0.007737f
C137 B.n15 VSUBS 0.007737f
C138 B.n16 VSUBS 0.007737f
C139 B.n17 VSUBS 0.007737f
C140 B.n18 VSUBS 0.007737f
C141 B.n19 VSUBS 0.007737f
C142 B.n20 VSUBS 0.007737f
C143 B.n21 VSUBS 0.007737f
C144 B.n22 VSUBS 0.007737f
C145 B.n23 VSUBS 0.007737f
C146 B.n24 VSUBS 0.007737f
C147 B.n25 VSUBS 0.007737f
C148 B.n26 VSUBS 0.007737f
C149 B.n27 VSUBS 0.016115f
C150 B.n28 VSUBS 0.007737f
C151 B.n29 VSUBS 0.007737f
C152 B.n30 VSUBS 0.007737f
C153 B.n31 VSUBS 0.007737f
C154 B.n32 VSUBS 0.007737f
C155 B.n33 VSUBS 0.007737f
C156 B.n34 VSUBS 0.007737f
C157 B.n35 VSUBS 0.007737f
C158 B.t5 VSUBS 0.072875f
C159 B.t4 VSUBS 0.087113f
C160 B.t3 VSUBS 0.312273f
C161 B.n36 VSUBS 0.082658f
C162 B.n37 VSUBS 0.068343f
C163 B.n38 VSUBS 0.007737f
C164 B.n39 VSUBS 0.007737f
C165 B.n40 VSUBS 0.007737f
C166 B.n41 VSUBS 0.007737f
C167 B.t8 VSUBS 0.072875f
C168 B.t7 VSUBS 0.087113f
C169 B.t6 VSUBS 0.312273f
C170 B.n42 VSUBS 0.082658f
C171 B.n43 VSUBS 0.068342f
C172 B.n44 VSUBS 0.007737f
C173 B.n45 VSUBS 0.007737f
C174 B.n46 VSUBS 0.007737f
C175 B.n47 VSUBS 0.007737f
C176 B.n48 VSUBS 0.007737f
C177 B.n49 VSUBS 0.007737f
C178 B.n50 VSUBS 0.007737f
C179 B.n51 VSUBS 0.016115f
C180 B.n52 VSUBS 0.007737f
C181 B.n53 VSUBS 0.007737f
C182 B.n54 VSUBS 0.007737f
C183 B.n55 VSUBS 0.007737f
C184 B.n56 VSUBS 0.007737f
C185 B.n57 VSUBS 0.007737f
C186 B.n58 VSUBS 0.007737f
C187 B.n59 VSUBS 0.007737f
C188 B.n60 VSUBS 0.007737f
C189 B.n61 VSUBS 0.007737f
C190 B.n62 VSUBS 0.007737f
C191 B.n63 VSUBS 0.007737f
C192 B.n64 VSUBS 0.007737f
C193 B.n65 VSUBS 0.007737f
C194 B.n66 VSUBS 0.007737f
C195 B.n67 VSUBS 0.007737f
C196 B.n68 VSUBS 0.007737f
C197 B.n69 VSUBS 0.007737f
C198 B.n70 VSUBS 0.007737f
C199 B.n71 VSUBS 0.007737f
C200 B.n72 VSUBS 0.007737f
C201 B.n73 VSUBS 0.007737f
C202 B.n74 VSUBS 0.007737f
C203 B.n75 VSUBS 0.007737f
C204 B.n76 VSUBS 0.007737f
C205 B.n77 VSUBS 0.007737f
C206 B.n78 VSUBS 0.007737f
C207 B.n79 VSUBS 0.007737f
C208 B.n80 VSUBS 0.007737f
C209 B.n81 VSUBS 0.007737f
C210 B.n82 VSUBS 0.007737f
C211 B.n83 VSUBS 0.007737f
C212 B.n84 VSUBS 0.007737f
C213 B.n85 VSUBS 0.007737f
C214 B.n86 VSUBS 0.007737f
C215 B.n87 VSUBS 0.007737f
C216 B.n88 VSUBS 0.007737f
C217 B.n89 VSUBS 0.007737f
C218 B.n90 VSUBS 0.007737f
C219 B.n91 VSUBS 0.007737f
C220 B.n92 VSUBS 0.007737f
C221 B.n93 VSUBS 0.007737f
C222 B.n94 VSUBS 0.007737f
C223 B.n95 VSUBS 0.007737f
C224 B.n96 VSUBS 0.007737f
C225 B.n97 VSUBS 0.007737f
C226 B.n98 VSUBS 0.007737f
C227 B.n99 VSUBS 0.007737f
C228 B.n100 VSUBS 0.007737f
C229 B.n101 VSUBS 0.007737f
C230 B.n102 VSUBS 0.016115f
C231 B.n103 VSUBS 0.007737f
C232 B.n104 VSUBS 0.007737f
C233 B.n105 VSUBS 0.007737f
C234 B.n106 VSUBS 0.007737f
C235 B.n107 VSUBS 0.007737f
C236 B.n108 VSUBS 0.007737f
C237 B.n109 VSUBS 0.007737f
C238 B.t1 VSUBS 0.072875f
C239 B.t2 VSUBS 0.087113f
C240 B.t0 VSUBS 0.312273f
C241 B.n110 VSUBS 0.082658f
C242 B.n111 VSUBS 0.068342f
C243 B.n112 VSUBS 0.017927f
C244 B.n113 VSUBS 0.007737f
C245 B.n114 VSUBS 0.007737f
C246 B.n115 VSUBS 0.007737f
C247 B.n116 VSUBS 0.007737f
C248 B.n117 VSUBS 0.007737f
C249 B.t10 VSUBS 0.072875f
C250 B.t11 VSUBS 0.087113f
C251 B.t9 VSUBS 0.312273f
C252 B.n118 VSUBS 0.082658f
C253 B.n119 VSUBS 0.068343f
C254 B.n120 VSUBS 0.007737f
C255 B.n121 VSUBS 0.007737f
C256 B.n122 VSUBS 0.007737f
C257 B.n123 VSUBS 0.007737f
C258 B.n124 VSUBS 0.007737f
C259 B.n125 VSUBS 0.007737f
C260 B.n126 VSUBS 0.01711f
C261 B.n127 VSUBS 0.007737f
C262 B.n128 VSUBS 0.007737f
C263 B.n129 VSUBS 0.007737f
C264 B.n130 VSUBS 0.007737f
C265 B.n131 VSUBS 0.007737f
C266 B.n132 VSUBS 0.007737f
C267 B.n133 VSUBS 0.007737f
C268 B.n134 VSUBS 0.007737f
C269 B.n135 VSUBS 0.007737f
C270 B.n136 VSUBS 0.007737f
C271 B.n137 VSUBS 0.007737f
C272 B.n138 VSUBS 0.007737f
C273 B.n139 VSUBS 0.007737f
C274 B.n140 VSUBS 0.007737f
C275 B.n141 VSUBS 0.007737f
C276 B.n142 VSUBS 0.007737f
C277 B.n143 VSUBS 0.007737f
C278 B.n144 VSUBS 0.007737f
C279 B.n145 VSUBS 0.007737f
C280 B.n146 VSUBS 0.007737f
C281 B.n147 VSUBS 0.007737f
C282 B.n148 VSUBS 0.007737f
C283 B.n149 VSUBS 0.007737f
C284 B.n150 VSUBS 0.007737f
C285 B.n151 VSUBS 0.007737f
C286 B.n152 VSUBS 0.007737f
C287 B.n153 VSUBS 0.007737f
C288 B.n154 VSUBS 0.007737f
C289 B.n155 VSUBS 0.007737f
C290 B.n156 VSUBS 0.007737f
C291 B.n157 VSUBS 0.007737f
C292 B.n158 VSUBS 0.007737f
C293 B.n159 VSUBS 0.007737f
C294 B.n160 VSUBS 0.007737f
C295 B.n161 VSUBS 0.007737f
C296 B.n162 VSUBS 0.007737f
C297 B.n163 VSUBS 0.007737f
C298 B.n164 VSUBS 0.007737f
C299 B.n165 VSUBS 0.007737f
C300 B.n166 VSUBS 0.007737f
C301 B.n167 VSUBS 0.007737f
C302 B.n168 VSUBS 0.007737f
C303 B.n169 VSUBS 0.007737f
C304 B.n170 VSUBS 0.007737f
C305 B.n171 VSUBS 0.007737f
C306 B.n172 VSUBS 0.007737f
C307 B.n173 VSUBS 0.007737f
C308 B.n174 VSUBS 0.007737f
C309 B.n175 VSUBS 0.007737f
C310 B.n176 VSUBS 0.007737f
C311 B.n177 VSUBS 0.007737f
C312 B.n178 VSUBS 0.007737f
C313 B.n179 VSUBS 0.007737f
C314 B.n180 VSUBS 0.007737f
C315 B.n181 VSUBS 0.007737f
C316 B.n182 VSUBS 0.007737f
C317 B.n183 VSUBS 0.007737f
C318 B.n184 VSUBS 0.007737f
C319 B.n185 VSUBS 0.007737f
C320 B.n186 VSUBS 0.007737f
C321 B.n187 VSUBS 0.007737f
C322 B.n188 VSUBS 0.007737f
C323 B.n189 VSUBS 0.007737f
C324 B.n190 VSUBS 0.007737f
C325 B.n191 VSUBS 0.007737f
C326 B.n192 VSUBS 0.007737f
C327 B.n193 VSUBS 0.007737f
C328 B.n194 VSUBS 0.007737f
C329 B.n195 VSUBS 0.007737f
C330 B.n196 VSUBS 0.007737f
C331 B.n197 VSUBS 0.007737f
C332 B.n198 VSUBS 0.007737f
C333 B.n199 VSUBS 0.007737f
C334 B.n200 VSUBS 0.007737f
C335 B.n201 VSUBS 0.007737f
C336 B.n202 VSUBS 0.007737f
C337 B.n203 VSUBS 0.007737f
C338 B.n204 VSUBS 0.007737f
C339 B.n205 VSUBS 0.007737f
C340 B.n206 VSUBS 0.007737f
C341 B.n207 VSUBS 0.007737f
C342 B.n208 VSUBS 0.007737f
C343 B.n209 VSUBS 0.007737f
C344 B.n210 VSUBS 0.007737f
C345 B.n211 VSUBS 0.007737f
C346 B.n212 VSUBS 0.007737f
C347 B.n213 VSUBS 0.007737f
C348 B.n214 VSUBS 0.007737f
C349 B.n215 VSUBS 0.007737f
C350 B.n216 VSUBS 0.007737f
C351 B.n217 VSUBS 0.007737f
C352 B.n218 VSUBS 0.007737f
C353 B.n219 VSUBS 0.007737f
C354 B.n220 VSUBS 0.007737f
C355 B.n221 VSUBS 0.007737f
C356 B.n222 VSUBS 0.007737f
C357 B.n223 VSUBS 0.007737f
C358 B.n224 VSUBS 0.007737f
C359 B.n225 VSUBS 0.016115f
C360 B.n226 VSUBS 0.016115f
C361 B.n227 VSUBS 0.01711f
C362 B.n228 VSUBS 0.007737f
C363 B.n229 VSUBS 0.007737f
C364 B.n230 VSUBS 0.007737f
C365 B.n231 VSUBS 0.007737f
C366 B.n232 VSUBS 0.007737f
C367 B.n233 VSUBS 0.007737f
C368 B.n234 VSUBS 0.007737f
C369 B.n235 VSUBS 0.007737f
C370 B.n236 VSUBS 0.007737f
C371 B.n237 VSUBS 0.007737f
C372 B.n238 VSUBS 0.007737f
C373 B.n239 VSUBS 0.007737f
C374 B.n240 VSUBS 0.007737f
C375 B.n241 VSUBS 0.007737f
C376 B.n242 VSUBS 0.007737f
C377 B.n243 VSUBS 0.007737f
C378 B.n244 VSUBS 0.007737f
C379 B.n245 VSUBS 0.007737f
C380 B.n246 VSUBS 0.007737f
C381 B.n247 VSUBS 0.007737f
C382 B.n248 VSUBS 0.005348f
C383 B.n249 VSUBS 0.017927f
C384 B.n250 VSUBS 0.006258f
C385 B.n251 VSUBS 0.007737f
C386 B.n252 VSUBS 0.007737f
C387 B.n253 VSUBS 0.007737f
C388 B.n254 VSUBS 0.007737f
C389 B.n255 VSUBS 0.007737f
C390 B.n256 VSUBS 0.007737f
C391 B.n257 VSUBS 0.007737f
C392 B.n258 VSUBS 0.007737f
C393 B.n259 VSUBS 0.007737f
C394 B.n260 VSUBS 0.007737f
C395 B.n261 VSUBS 0.007737f
C396 B.n262 VSUBS 0.006258f
C397 B.n263 VSUBS 0.007737f
C398 B.n264 VSUBS 0.007737f
C399 B.n265 VSUBS 0.005348f
C400 B.n266 VSUBS 0.007737f
C401 B.n267 VSUBS 0.007737f
C402 B.n268 VSUBS 0.007737f
C403 B.n269 VSUBS 0.007737f
C404 B.n270 VSUBS 0.007737f
C405 B.n271 VSUBS 0.007737f
C406 B.n272 VSUBS 0.007737f
C407 B.n273 VSUBS 0.007737f
C408 B.n274 VSUBS 0.007737f
C409 B.n275 VSUBS 0.007737f
C410 B.n276 VSUBS 0.007737f
C411 B.n277 VSUBS 0.007737f
C412 B.n278 VSUBS 0.007737f
C413 B.n279 VSUBS 0.007737f
C414 B.n280 VSUBS 0.007737f
C415 B.n281 VSUBS 0.007737f
C416 B.n282 VSUBS 0.007737f
C417 B.n283 VSUBS 0.007737f
C418 B.n284 VSUBS 0.007737f
C419 B.n285 VSUBS 0.01711f
C420 B.n286 VSUBS 0.01711f
C421 B.n287 VSUBS 0.016115f
C422 B.n288 VSUBS 0.007737f
C423 B.n289 VSUBS 0.007737f
C424 B.n290 VSUBS 0.007737f
C425 B.n291 VSUBS 0.007737f
C426 B.n292 VSUBS 0.007737f
C427 B.n293 VSUBS 0.007737f
C428 B.n294 VSUBS 0.007737f
C429 B.n295 VSUBS 0.007737f
C430 B.n296 VSUBS 0.007737f
C431 B.n297 VSUBS 0.007737f
C432 B.n298 VSUBS 0.007737f
C433 B.n299 VSUBS 0.007737f
C434 B.n300 VSUBS 0.007737f
C435 B.n301 VSUBS 0.007737f
C436 B.n302 VSUBS 0.007737f
C437 B.n303 VSUBS 0.007737f
C438 B.n304 VSUBS 0.007737f
C439 B.n305 VSUBS 0.007737f
C440 B.n306 VSUBS 0.007737f
C441 B.n307 VSUBS 0.007737f
C442 B.n308 VSUBS 0.007737f
C443 B.n309 VSUBS 0.007737f
C444 B.n310 VSUBS 0.007737f
C445 B.n311 VSUBS 0.007737f
C446 B.n312 VSUBS 0.007737f
C447 B.n313 VSUBS 0.007737f
C448 B.n314 VSUBS 0.007737f
C449 B.n315 VSUBS 0.007737f
C450 B.n316 VSUBS 0.007737f
C451 B.n317 VSUBS 0.007737f
C452 B.n318 VSUBS 0.007737f
C453 B.n319 VSUBS 0.007737f
C454 B.n320 VSUBS 0.007737f
C455 B.n321 VSUBS 0.007737f
C456 B.n322 VSUBS 0.007737f
C457 B.n323 VSUBS 0.007737f
C458 B.n324 VSUBS 0.007737f
C459 B.n325 VSUBS 0.007737f
C460 B.n326 VSUBS 0.007737f
C461 B.n327 VSUBS 0.007737f
C462 B.n328 VSUBS 0.007737f
C463 B.n329 VSUBS 0.007737f
C464 B.n330 VSUBS 0.007737f
C465 B.n331 VSUBS 0.007737f
C466 B.n332 VSUBS 0.007737f
C467 B.n333 VSUBS 0.007737f
C468 B.n334 VSUBS 0.007737f
C469 B.n335 VSUBS 0.007737f
C470 B.n336 VSUBS 0.007737f
C471 B.n337 VSUBS 0.007737f
C472 B.n338 VSUBS 0.007737f
C473 B.n339 VSUBS 0.007737f
C474 B.n340 VSUBS 0.007737f
C475 B.n341 VSUBS 0.007737f
C476 B.n342 VSUBS 0.007737f
C477 B.n343 VSUBS 0.007737f
C478 B.n344 VSUBS 0.007737f
C479 B.n345 VSUBS 0.007737f
C480 B.n346 VSUBS 0.007737f
C481 B.n347 VSUBS 0.007737f
C482 B.n348 VSUBS 0.007737f
C483 B.n349 VSUBS 0.007737f
C484 B.n350 VSUBS 0.007737f
C485 B.n351 VSUBS 0.007737f
C486 B.n352 VSUBS 0.007737f
C487 B.n353 VSUBS 0.007737f
C488 B.n354 VSUBS 0.007737f
C489 B.n355 VSUBS 0.007737f
C490 B.n356 VSUBS 0.007737f
C491 B.n357 VSUBS 0.007737f
C492 B.n358 VSUBS 0.007737f
C493 B.n359 VSUBS 0.007737f
C494 B.n360 VSUBS 0.007737f
C495 B.n361 VSUBS 0.007737f
C496 B.n362 VSUBS 0.007737f
C497 B.n363 VSUBS 0.007737f
C498 B.n364 VSUBS 0.007737f
C499 B.n365 VSUBS 0.007737f
C500 B.n366 VSUBS 0.007737f
C501 B.n367 VSUBS 0.007737f
C502 B.n368 VSUBS 0.007737f
C503 B.n369 VSUBS 0.007737f
C504 B.n370 VSUBS 0.007737f
C505 B.n371 VSUBS 0.007737f
C506 B.n372 VSUBS 0.007737f
C507 B.n373 VSUBS 0.007737f
C508 B.n374 VSUBS 0.007737f
C509 B.n375 VSUBS 0.007737f
C510 B.n376 VSUBS 0.007737f
C511 B.n377 VSUBS 0.007737f
C512 B.n378 VSUBS 0.007737f
C513 B.n379 VSUBS 0.007737f
C514 B.n380 VSUBS 0.007737f
C515 B.n381 VSUBS 0.007737f
C516 B.n382 VSUBS 0.007737f
C517 B.n383 VSUBS 0.007737f
C518 B.n384 VSUBS 0.007737f
C519 B.n385 VSUBS 0.007737f
C520 B.n386 VSUBS 0.007737f
C521 B.n387 VSUBS 0.007737f
C522 B.n388 VSUBS 0.007737f
C523 B.n389 VSUBS 0.007737f
C524 B.n390 VSUBS 0.007737f
C525 B.n391 VSUBS 0.007737f
C526 B.n392 VSUBS 0.007737f
C527 B.n393 VSUBS 0.007737f
C528 B.n394 VSUBS 0.007737f
C529 B.n395 VSUBS 0.007737f
C530 B.n396 VSUBS 0.007737f
C531 B.n397 VSUBS 0.007737f
C532 B.n398 VSUBS 0.007737f
C533 B.n399 VSUBS 0.007737f
C534 B.n400 VSUBS 0.007737f
C535 B.n401 VSUBS 0.007737f
C536 B.n402 VSUBS 0.007737f
C537 B.n403 VSUBS 0.007737f
C538 B.n404 VSUBS 0.007737f
C539 B.n405 VSUBS 0.007737f
C540 B.n406 VSUBS 0.007737f
C541 B.n407 VSUBS 0.007737f
C542 B.n408 VSUBS 0.007737f
C543 B.n409 VSUBS 0.007737f
C544 B.n410 VSUBS 0.007737f
C545 B.n411 VSUBS 0.007737f
C546 B.n412 VSUBS 0.007737f
C547 B.n413 VSUBS 0.007737f
C548 B.n414 VSUBS 0.007737f
C549 B.n415 VSUBS 0.007737f
C550 B.n416 VSUBS 0.007737f
C551 B.n417 VSUBS 0.007737f
C552 B.n418 VSUBS 0.007737f
C553 B.n419 VSUBS 0.007737f
C554 B.n420 VSUBS 0.007737f
C555 B.n421 VSUBS 0.007737f
C556 B.n422 VSUBS 0.007737f
C557 B.n423 VSUBS 0.007737f
C558 B.n424 VSUBS 0.007737f
C559 B.n425 VSUBS 0.007737f
C560 B.n426 VSUBS 0.007737f
C561 B.n427 VSUBS 0.007737f
C562 B.n428 VSUBS 0.007737f
C563 B.n429 VSUBS 0.007737f
C564 B.n430 VSUBS 0.007737f
C565 B.n431 VSUBS 0.007737f
C566 B.n432 VSUBS 0.007737f
C567 B.n433 VSUBS 0.007737f
C568 B.n434 VSUBS 0.007737f
C569 B.n435 VSUBS 0.007737f
C570 B.n436 VSUBS 0.007737f
C571 B.n437 VSUBS 0.007737f
C572 B.n438 VSUBS 0.007737f
C573 B.n439 VSUBS 0.007737f
C574 B.n440 VSUBS 0.017161f
C575 B.n441 VSUBS 0.016065f
C576 B.n442 VSUBS 0.01711f
C577 B.n443 VSUBS 0.007737f
C578 B.n444 VSUBS 0.007737f
C579 B.n445 VSUBS 0.007737f
C580 B.n446 VSUBS 0.007737f
C581 B.n447 VSUBS 0.007737f
C582 B.n448 VSUBS 0.007737f
C583 B.n449 VSUBS 0.007737f
C584 B.n450 VSUBS 0.007737f
C585 B.n451 VSUBS 0.007737f
C586 B.n452 VSUBS 0.007737f
C587 B.n453 VSUBS 0.007737f
C588 B.n454 VSUBS 0.007737f
C589 B.n455 VSUBS 0.007737f
C590 B.n456 VSUBS 0.007737f
C591 B.n457 VSUBS 0.007737f
C592 B.n458 VSUBS 0.007737f
C593 B.n459 VSUBS 0.007737f
C594 B.n460 VSUBS 0.007737f
C595 B.n461 VSUBS 0.007737f
C596 B.n462 VSUBS 0.007737f
C597 B.n463 VSUBS 0.005348f
C598 B.n464 VSUBS 0.017927f
C599 B.n465 VSUBS 0.006258f
C600 B.n466 VSUBS 0.007737f
C601 B.n467 VSUBS 0.007737f
C602 B.n468 VSUBS 0.007737f
C603 B.n469 VSUBS 0.007737f
C604 B.n470 VSUBS 0.007737f
C605 B.n471 VSUBS 0.007737f
C606 B.n472 VSUBS 0.007737f
C607 B.n473 VSUBS 0.007737f
C608 B.n474 VSUBS 0.007737f
C609 B.n475 VSUBS 0.007737f
C610 B.n476 VSUBS 0.007737f
C611 B.n477 VSUBS 0.006258f
C612 B.n478 VSUBS 0.017927f
C613 B.n479 VSUBS 0.005348f
C614 B.n480 VSUBS 0.007737f
C615 B.n481 VSUBS 0.007737f
C616 B.n482 VSUBS 0.007737f
C617 B.n483 VSUBS 0.007737f
C618 B.n484 VSUBS 0.007737f
C619 B.n485 VSUBS 0.007737f
C620 B.n486 VSUBS 0.007737f
C621 B.n487 VSUBS 0.007737f
C622 B.n488 VSUBS 0.007737f
C623 B.n489 VSUBS 0.007737f
C624 B.n490 VSUBS 0.007737f
C625 B.n491 VSUBS 0.007737f
C626 B.n492 VSUBS 0.007737f
C627 B.n493 VSUBS 0.007737f
C628 B.n494 VSUBS 0.007737f
C629 B.n495 VSUBS 0.007737f
C630 B.n496 VSUBS 0.007737f
C631 B.n497 VSUBS 0.007737f
C632 B.n498 VSUBS 0.007737f
C633 B.n499 VSUBS 0.007737f
C634 B.n500 VSUBS 0.01711f
C635 B.n501 VSUBS 0.01711f
C636 B.n502 VSUBS 0.016115f
C637 B.n503 VSUBS 0.007737f
C638 B.n504 VSUBS 0.007737f
C639 B.n505 VSUBS 0.007737f
C640 B.n506 VSUBS 0.007737f
C641 B.n507 VSUBS 0.007737f
C642 B.n508 VSUBS 0.007737f
C643 B.n509 VSUBS 0.007737f
C644 B.n510 VSUBS 0.007737f
C645 B.n511 VSUBS 0.007737f
C646 B.n512 VSUBS 0.007737f
C647 B.n513 VSUBS 0.007737f
C648 B.n514 VSUBS 0.007737f
C649 B.n515 VSUBS 0.007737f
C650 B.n516 VSUBS 0.007737f
C651 B.n517 VSUBS 0.007737f
C652 B.n518 VSUBS 0.007737f
C653 B.n519 VSUBS 0.007737f
C654 B.n520 VSUBS 0.007737f
C655 B.n521 VSUBS 0.007737f
C656 B.n522 VSUBS 0.007737f
C657 B.n523 VSUBS 0.007737f
C658 B.n524 VSUBS 0.007737f
C659 B.n525 VSUBS 0.007737f
C660 B.n526 VSUBS 0.007737f
C661 B.n527 VSUBS 0.007737f
C662 B.n528 VSUBS 0.007737f
C663 B.n529 VSUBS 0.007737f
C664 B.n530 VSUBS 0.007737f
C665 B.n531 VSUBS 0.007737f
C666 B.n532 VSUBS 0.007737f
C667 B.n533 VSUBS 0.007737f
C668 B.n534 VSUBS 0.007737f
C669 B.n535 VSUBS 0.007737f
C670 B.n536 VSUBS 0.007737f
C671 B.n537 VSUBS 0.007737f
C672 B.n538 VSUBS 0.007737f
C673 B.n539 VSUBS 0.007737f
C674 B.n540 VSUBS 0.007737f
C675 B.n541 VSUBS 0.007737f
C676 B.n542 VSUBS 0.007737f
C677 B.n543 VSUBS 0.007737f
C678 B.n544 VSUBS 0.007737f
C679 B.n545 VSUBS 0.007737f
C680 B.n546 VSUBS 0.007737f
C681 B.n547 VSUBS 0.007737f
C682 B.n548 VSUBS 0.007737f
C683 B.n549 VSUBS 0.007737f
C684 B.n550 VSUBS 0.007737f
C685 B.n551 VSUBS 0.007737f
C686 B.n552 VSUBS 0.007737f
C687 B.n553 VSUBS 0.007737f
C688 B.n554 VSUBS 0.007737f
C689 B.n555 VSUBS 0.007737f
C690 B.n556 VSUBS 0.007737f
C691 B.n557 VSUBS 0.007737f
C692 B.n558 VSUBS 0.007737f
C693 B.n559 VSUBS 0.007737f
C694 B.n560 VSUBS 0.007737f
C695 B.n561 VSUBS 0.007737f
C696 B.n562 VSUBS 0.007737f
C697 B.n563 VSUBS 0.007737f
C698 B.n564 VSUBS 0.007737f
C699 B.n565 VSUBS 0.007737f
C700 B.n566 VSUBS 0.007737f
C701 B.n567 VSUBS 0.007737f
C702 B.n568 VSUBS 0.007737f
C703 B.n569 VSUBS 0.007737f
C704 B.n570 VSUBS 0.007737f
C705 B.n571 VSUBS 0.007737f
C706 B.n572 VSUBS 0.007737f
C707 B.n573 VSUBS 0.007737f
C708 B.n574 VSUBS 0.007737f
C709 B.n575 VSUBS 0.007737f
C710 B.n576 VSUBS 0.007737f
C711 B.n577 VSUBS 0.007737f
C712 B.n578 VSUBS 0.007737f
C713 B.n579 VSUBS 0.01752f
C714 VTAIL.t0 VSUBS 0.072472f
C715 VTAIL.t18 VSUBS 0.072472f
C716 VTAIL.n0 VSUBS 0.317475f
C717 VTAIL.n1 VSUBS 0.743205f
C718 VTAIL.t9 VSUBS 0.476531f
C719 VTAIL.n2 VSUBS 0.830878f
C720 VTAIL.t11 VSUBS 0.072472f
C721 VTAIL.t16 VSUBS 0.072472f
C722 VTAIL.n3 VSUBS 0.317475f
C723 VTAIL.n4 VSUBS 0.853004f
C724 VTAIL.t7 VSUBS 0.072472f
C725 VTAIL.t14 VSUBS 0.072472f
C726 VTAIL.n5 VSUBS 0.317475f
C727 VTAIL.n6 VSUBS 1.77523f
C728 VTAIL.t3 VSUBS 0.072472f
C729 VTAIL.t4 VSUBS 0.072472f
C730 VTAIL.n7 VSUBS 0.317476f
C731 VTAIL.n8 VSUBS 1.77523f
C732 VTAIL.t2 VSUBS 0.072472f
C733 VTAIL.t19 VSUBS 0.072472f
C734 VTAIL.n9 VSUBS 0.317476f
C735 VTAIL.n10 VSUBS 0.853002f
C736 VTAIL.t6 VSUBS 0.476532f
C737 VTAIL.n11 VSUBS 0.830877f
C738 VTAIL.t13 VSUBS 0.072472f
C739 VTAIL.t8 VSUBS 0.072472f
C740 VTAIL.n12 VSUBS 0.317476f
C741 VTAIL.n13 VSUBS 0.792282f
C742 VTAIL.t10 VSUBS 0.072472f
C743 VTAIL.t15 VSUBS 0.072472f
C744 VTAIL.n14 VSUBS 0.317476f
C745 VTAIL.n15 VSUBS 0.853002f
C746 VTAIL.t12 VSUBS 0.476531f
C747 VTAIL.n16 VSUBS 1.59286f
C748 VTAIL.t17 VSUBS 0.476531f
C749 VTAIL.n17 VSUBS 1.59286f
C750 VTAIL.t1 VSUBS 0.072472f
C751 VTAIL.t5 VSUBS 0.072472f
C752 VTAIL.n18 VSUBS 0.317475f
C753 VTAIL.n19 VSUBS 0.681116f
C754 VDD1.t7 VSUBS 0.390708f
C755 VDD1.t6 VSUBS 0.052443f
C756 VDD1.t3 VSUBS 0.052443f
C757 VDD1.n0 VSUBS 0.268863f
C758 VDD1.n1 VSUBS 0.976326f
C759 VDD1.t9 VSUBS 0.390707f
C760 VDD1.t8 VSUBS 0.052443f
C761 VDD1.t0 VSUBS 0.052443f
C762 VDD1.n2 VSUBS 0.268862f
C763 VDD1.n3 VSUBS 0.968809f
C764 VDD1.t5 VSUBS 0.052443f
C765 VDD1.t1 VSUBS 0.052443f
C766 VDD1.n4 VSUBS 0.275067f
C767 VDD1.n5 VSUBS 2.18454f
C768 VDD1.t4 VSUBS 0.052443f
C769 VDD1.t2 VSUBS 0.052443f
C770 VDD1.n6 VSUBS 0.268862f
C771 VDD1.n7 VSUBS 2.22781f
C772 VP.n0 VSUBS 0.068624f
C773 VP.t7 VSUBS 0.748963f
C774 VP.n1 VSUBS 0.054593f
C775 VP.n2 VSUBS 0.052051f
C776 VP.t0 VSUBS 0.748963f
C777 VP.n3 VSUBS 0.081787f
C778 VP.n4 VSUBS 0.052051f
C779 VP.t5 VSUBS 0.748963f
C780 VP.n5 VSUBS 0.09701f
C781 VP.n6 VSUBS 0.052051f
C782 VP.t2 VSUBS 0.748963f
C783 VP.n7 VSUBS 0.331423f
C784 VP.n8 VSUBS 0.052051f
C785 VP.n9 VSUBS 0.092355f
C786 VP.n10 VSUBS 0.068624f
C787 VP.t4 VSUBS 0.748963f
C788 VP.n11 VSUBS 0.054593f
C789 VP.n12 VSUBS 0.052051f
C790 VP.t1 VSUBS 0.748963f
C791 VP.n13 VSUBS 0.081787f
C792 VP.n14 VSUBS 0.052051f
C793 VP.t6 VSUBS 0.748963f
C794 VP.n15 VSUBS 0.09701f
C795 VP.n16 VSUBS 0.052051f
C796 VP.t8 VSUBS 0.748963f
C797 VP.n17 VSUBS 0.477687f
C798 VP.t3 VSUBS 1.05751f
C799 VP.n18 VSUBS 0.43866f
C800 VP.n19 VSUBS 0.437782f
C801 VP.n20 VSUBS 0.089346f
C802 VP.n21 VSUBS 0.081787f
C803 VP.n22 VSUBS 0.070183f
C804 VP.n23 VSUBS 0.052051f
C805 VP.n24 VSUBS 0.052051f
C806 VP.n25 VSUBS 0.052051f
C807 VP.n26 VSUBS 0.380538f
C808 VP.n27 VSUBS 0.09701f
C809 VP.n28 VSUBS 0.070183f
C810 VP.n29 VSUBS 0.052051f
C811 VP.n30 VSUBS 0.052051f
C812 VP.n31 VSUBS 0.052051f
C813 VP.n32 VSUBS 0.089346f
C814 VP.n33 VSUBS 0.331423f
C815 VP.n34 VSUBS 0.056778f
C816 VP.n35 VSUBS 0.102031f
C817 VP.n36 VSUBS 0.052051f
C818 VP.n37 VSUBS 0.052051f
C819 VP.n38 VSUBS 0.052051f
C820 VP.n39 VSUBS 0.092355f
C821 VP.n40 VSUBS 0.081683f
C822 VP.n41 VSUBS 0.488318f
C823 VP.n42 VSUBS 2.31334f
C824 VP.n43 VSUBS 2.35648f
C825 VP.t9 VSUBS 0.748963f
C826 VP.n44 VSUBS 0.488318f
C827 VP.n45 VSUBS 0.081683f
C828 VP.n46 VSUBS 0.068624f
C829 VP.n47 VSUBS 0.052051f
C830 VP.n48 VSUBS 0.052051f
C831 VP.n49 VSUBS 0.054593f
C832 VP.n50 VSUBS 0.102031f
C833 VP.n51 VSUBS 0.056778f
C834 VP.n52 VSUBS 0.052051f
C835 VP.n53 VSUBS 0.052051f
C836 VP.n54 VSUBS 0.089346f
C837 VP.n55 VSUBS 0.081787f
C838 VP.n56 VSUBS 0.070183f
C839 VP.n57 VSUBS 0.052051f
C840 VP.n58 VSUBS 0.052051f
C841 VP.n59 VSUBS 0.052051f
C842 VP.n60 VSUBS 0.380538f
C843 VP.n61 VSUBS 0.09701f
C844 VP.n62 VSUBS 0.070183f
C845 VP.n63 VSUBS 0.052051f
C846 VP.n64 VSUBS 0.052051f
C847 VP.n65 VSUBS 0.052051f
C848 VP.n66 VSUBS 0.089346f
C849 VP.n67 VSUBS 0.331423f
C850 VP.n68 VSUBS 0.056778f
C851 VP.n69 VSUBS 0.102031f
C852 VP.n70 VSUBS 0.052051f
C853 VP.n71 VSUBS 0.052051f
C854 VP.n72 VSUBS 0.052051f
C855 VP.n73 VSUBS 0.092355f
C856 VP.n74 VSUBS 0.081683f
C857 VP.n75 VSUBS 0.488318f
C858 VP.n76 VSUBS 0.06861f
.ends

