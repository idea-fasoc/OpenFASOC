* NGSPICE file created from diff_pair_sample_1269.ext - technology: sky130A

.subckt diff_pair_sample_1269 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t11 VP.t0 VDD1.t2 B.t3 sky130_fd_pr__nfet_01v8 ad=2.40075 pd=14.88 as=2.40075 ps=14.88 w=14.55 l=3.08
X1 VDD1.t4 VP.t1 VTAIL.t10 B.t0 sky130_fd_pr__nfet_01v8 ad=5.6745 pd=29.88 as=2.40075 ps=14.88 w=14.55 l=3.08
X2 B.t19 B.t17 B.t18 B.t14 sky130_fd_pr__nfet_01v8 ad=5.6745 pd=29.88 as=0 ps=0 w=14.55 l=3.08
X3 VTAIL.t9 VP.t2 VDD1.t1 B.t5 sky130_fd_pr__nfet_01v8 ad=2.40075 pd=14.88 as=2.40075 ps=14.88 w=14.55 l=3.08
X4 VDD2.t5 VN.t0 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=5.6745 pd=29.88 as=2.40075 ps=14.88 w=14.55 l=3.08
X5 B.t16 B.t13 B.t15 B.t14 sky130_fd_pr__nfet_01v8 ad=5.6745 pd=29.88 as=0 ps=0 w=14.55 l=3.08
X6 VTAIL.t3 VN.t1 VDD2.t4 B.t3 sky130_fd_pr__nfet_01v8 ad=2.40075 pd=14.88 as=2.40075 ps=14.88 w=14.55 l=3.08
X7 VDD1.t0 VP.t3 VTAIL.t8 B.t2 sky130_fd_pr__nfet_01v8 ad=5.6745 pd=29.88 as=2.40075 ps=14.88 w=14.55 l=3.08
X8 VDD2.t3 VN.t2 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=5.6745 pd=29.88 as=2.40075 ps=14.88 w=14.55 l=3.08
X9 VDD2.t2 VN.t3 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=2.40075 pd=14.88 as=5.6745 ps=29.88 w=14.55 l=3.08
X10 VDD2.t1 VN.t4 VTAIL.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=2.40075 pd=14.88 as=5.6745 ps=29.88 w=14.55 l=3.08
X11 B.t12 B.t10 B.t11 B.t7 sky130_fd_pr__nfet_01v8 ad=5.6745 pd=29.88 as=0 ps=0 w=14.55 l=3.08
X12 VDD1.t5 VP.t4 VTAIL.t7 B.t4 sky130_fd_pr__nfet_01v8 ad=2.40075 pd=14.88 as=5.6745 ps=29.88 w=14.55 l=3.08
X13 B.t9 B.t6 B.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=5.6745 pd=29.88 as=0 ps=0 w=14.55 l=3.08
X14 VTAIL.t5 VN.t5 VDD2.t0 B.t5 sky130_fd_pr__nfet_01v8 ad=2.40075 pd=14.88 as=2.40075 ps=14.88 w=14.55 l=3.08
X15 VDD1.t3 VP.t5 VTAIL.t6 B.t1 sky130_fd_pr__nfet_01v8 ad=2.40075 pd=14.88 as=5.6745 ps=29.88 w=14.55 l=3.08
R0 VP.n13 VP.n10 161.3
R1 VP.n15 VP.n14 161.3
R2 VP.n16 VP.n9 161.3
R3 VP.n18 VP.n17 161.3
R4 VP.n19 VP.n8 161.3
R5 VP.n21 VP.n20 161.3
R6 VP.n44 VP.n43 161.3
R7 VP.n42 VP.n1 161.3
R8 VP.n41 VP.n40 161.3
R9 VP.n39 VP.n2 161.3
R10 VP.n38 VP.n37 161.3
R11 VP.n36 VP.n3 161.3
R12 VP.n35 VP.n34 161.3
R13 VP.n33 VP.n4 161.3
R14 VP.n32 VP.n31 161.3
R15 VP.n30 VP.n5 161.3
R16 VP.n29 VP.n28 161.3
R17 VP.n27 VP.n6 161.3
R18 VP.n26 VP.n25 161.3
R19 VP.n11 VP.t3 147.25
R20 VP.n35 VP.t0 113.85
R21 VP.n24 VP.t1 113.85
R22 VP.n0 VP.t5 113.85
R23 VP.n12 VP.t2 113.85
R24 VP.n7 VP.t4 113.85
R25 VP.n24 VP.n23 70.0045
R26 VP.n45 VP.n0 70.0045
R27 VP.n22 VP.n7 70.0045
R28 VP.n30 VP.n29 56.5193
R29 VP.n41 VP.n2 56.5193
R30 VP.n18 VP.n9 56.5193
R31 VP.n23 VP.n22 52.6319
R32 VP.n12 VP.n11 49.4021
R33 VP.n25 VP.n6 24.4675
R34 VP.n29 VP.n6 24.4675
R35 VP.n31 VP.n30 24.4675
R36 VP.n31 VP.n4 24.4675
R37 VP.n35 VP.n4 24.4675
R38 VP.n36 VP.n35 24.4675
R39 VP.n37 VP.n36 24.4675
R40 VP.n37 VP.n2 24.4675
R41 VP.n42 VP.n41 24.4675
R42 VP.n43 VP.n42 24.4675
R43 VP.n19 VP.n18 24.4675
R44 VP.n20 VP.n19 24.4675
R45 VP.n13 VP.n12 24.4675
R46 VP.n14 VP.n13 24.4675
R47 VP.n14 VP.n9 24.4675
R48 VP.n25 VP.n24 20.0634
R49 VP.n43 VP.n0 20.0634
R50 VP.n20 VP.n7 20.0634
R51 VP.n11 VP.n10 3.91165
R52 VP.n22 VP.n21 0.354971
R53 VP.n26 VP.n23 0.354971
R54 VP.n45 VP.n44 0.354971
R55 VP VP.n45 0.26696
R56 VP.n15 VP.n10 0.189894
R57 VP.n16 VP.n15 0.189894
R58 VP.n17 VP.n16 0.189894
R59 VP.n17 VP.n8 0.189894
R60 VP.n21 VP.n8 0.189894
R61 VP.n27 VP.n26 0.189894
R62 VP.n28 VP.n27 0.189894
R63 VP.n28 VP.n5 0.189894
R64 VP.n32 VP.n5 0.189894
R65 VP.n33 VP.n32 0.189894
R66 VP.n34 VP.n33 0.189894
R67 VP.n34 VP.n3 0.189894
R68 VP.n38 VP.n3 0.189894
R69 VP.n39 VP.n38 0.189894
R70 VP.n40 VP.n39 0.189894
R71 VP.n40 VP.n1 0.189894
R72 VP.n44 VP.n1 0.189894
R73 VDD1 VDD1.t0 63.2508
R74 VDD1.n1 VDD1.t4 63.137
R75 VDD1.n1 VDD1.n0 60.3065
R76 VDD1.n3 VDD1.n2 59.627
R77 VDD1.n3 VDD1.n1 47.8651
R78 VDD1.n2 VDD1.t1 1.36132
R79 VDD1.n2 VDD1.t5 1.36132
R80 VDD1.n0 VDD1.t2 1.36132
R81 VDD1.n0 VDD1.t3 1.36132
R82 VDD1 VDD1.n3 0.677224
R83 VTAIL.n7 VTAIL.t1 44.3091
R84 VTAIL.n10 VTAIL.t7 44.309
R85 VTAIL.n11 VTAIL.t4 44.3088
R86 VTAIL.n2 VTAIL.t6 44.3088
R87 VTAIL.n9 VTAIL.n8 42.9482
R88 VTAIL.n6 VTAIL.n5 42.9482
R89 VTAIL.n1 VTAIL.n0 42.9482
R90 VTAIL.n4 VTAIL.n3 42.9482
R91 VTAIL.n6 VTAIL.n4 30.7893
R92 VTAIL.n11 VTAIL.n10 27.8496
R93 VTAIL.n7 VTAIL.n6 2.94016
R94 VTAIL.n10 VTAIL.n9 2.94016
R95 VTAIL.n4 VTAIL.n2 2.94016
R96 VTAIL VTAIL.n11 2.14705
R97 VTAIL.n9 VTAIL.n7 1.94016
R98 VTAIL.n2 VTAIL.n1 1.94016
R99 VTAIL.n0 VTAIL.t2 1.36132
R100 VTAIL.n0 VTAIL.t5 1.36132
R101 VTAIL.n3 VTAIL.t10 1.36132
R102 VTAIL.n3 VTAIL.t11 1.36132
R103 VTAIL.n8 VTAIL.t8 1.36132
R104 VTAIL.n8 VTAIL.t9 1.36132
R105 VTAIL.n5 VTAIL.t0 1.36132
R106 VTAIL.n5 VTAIL.t3 1.36132
R107 VTAIL VTAIL.n1 0.793603
R108 B.n936 B.n935 585
R109 B.n360 B.n143 585
R110 B.n359 B.n358 585
R111 B.n357 B.n356 585
R112 B.n355 B.n354 585
R113 B.n353 B.n352 585
R114 B.n351 B.n350 585
R115 B.n349 B.n348 585
R116 B.n347 B.n346 585
R117 B.n345 B.n344 585
R118 B.n343 B.n342 585
R119 B.n341 B.n340 585
R120 B.n339 B.n338 585
R121 B.n337 B.n336 585
R122 B.n335 B.n334 585
R123 B.n333 B.n332 585
R124 B.n331 B.n330 585
R125 B.n329 B.n328 585
R126 B.n327 B.n326 585
R127 B.n325 B.n324 585
R128 B.n323 B.n322 585
R129 B.n321 B.n320 585
R130 B.n319 B.n318 585
R131 B.n317 B.n316 585
R132 B.n315 B.n314 585
R133 B.n313 B.n312 585
R134 B.n311 B.n310 585
R135 B.n309 B.n308 585
R136 B.n307 B.n306 585
R137 B.n305 B.n304 585
R138 B.n303 B.n302 585
R139 B.n301 B.n300 585
R140 B.n299 B.n298 585
R141 B.n297 B.n296 585
R142 B.n295 B.n294 585
R143 B.n293 B.n292 585
R144 B.n291 B.n290 585
R145 B.n289 B.n288 585
R146 B.n287 B.n286 585
R147 B.n285 B.n284 585
R148 B.n283 B.n282 585
R149 B.n281 B.n280 585
R150 B.n279 B.n278 585
R151 B.n277 B.n276 585
R152 B.n275 B.n274 585
R153 B.n273 B.n272 585
R154 B.n271 B.n270 585
R155 B.n269 B.n268 585
R156 B.n267 B.n266 585
R157 B.n264 B.n263 585
R158 B.n262 B.n261 585
R159 B.n260 B.n259 585
R160 B.n258 B.n257 585
R161 B.n256 B.n255 585
R162 B.n254 B.n253 585
R163 B.n252 B.n251 585
R164 B.n250 B.n249 585
R165 B.n248 B.n247 585
R166 B.n246 B.n245 585
R167 B.n243 B.n242 585
R168 B.n241 B.n240 585
R169 B.n239 B.n238 585
R170 B.n237 B.n236 585
R171 B.n235 B.n234 585
R172 B.n233 B.n232 585
R173 B.n231 B.n230 585
R174 B.n229 B.n228 585
R175 B.n227 B.n226 585
R176 B.n225 B.n224 585
R177 B.n223 B.n222 585
R178 B.n221 B.n220 585
R179 B.n219 B.n218 585
R180 B.n217 B.n216 585
R181 B.n215 B.n214 585
R182 B.n213 B.n212 585
R183 B.n211 B.n210 585
R184 B.n209 B.n208 585
R185 B.n207 B.n206 585
R186 B.n205 B.n204 585
R187 B.n203 B.n202 585
R188 B.n201 B.n200 585
R189 B.n199 B.n198 585
R190 B.n197 B.n196 585
R191 B.n195 B.n194 585
R192 B.n193 B.n192 585
R193 B.n191 B.n190 585
R194 B.n189 B.n188 585
R195 B.n187 B.n186 585
R196 B.n185 B.n184 585
R197 B.n183 B.n182 585
R198 B.n181 B.n180 585
R199 B.n179 B.n178 585
R200 B.n177 B.n176 585
R201 B.n175 B.n174 585
R202 B.n173 B.n172 585
R203 B.n171 B.n170 585
R204 B.n169 B.n168 585
R205 B.n167 B.n166 585
R206 B.n165 B.n164 585
R207 B.n163 B.n162 585
R208 B.n161 B.n160 585
R209 B.n159 B.n158 585
R210 B.n157 B.n156 585
R211 B.n155 B.n154 585
R212 B.n153 B.n152 585
R213 B.n151 B.n150 585
R214 B.n149 B.n148 585
R215 B.n88 B.n87 585
R216 B.n934 B.n89 585
R217 B.n939 B.n89 585
R218 B.n933 B.n932 585
R219 B.n932 B.n85 585
R220 B.n931 B.n84 585
R221 B.n945 B.n84 585
R222 B.n930 B.n83 585
R223 B.n946 B.n83 585
R224 B.n929 B.n82 585
R225 B.n947 B.n82 585
R226 B.n928 B.n927 585
R227 B.n927 B.n78 585
R228 B.n926 B.n77 585
R229 B.n953 B.n77 585
R230 B.n925 B.n76 585
R231 B.n954 B.n76 585
R232 B.n924 B.n75 585
R233 B.n955 B.n75 585
R234 B.n923 B.n922 585
R235 B.n922 B.n71 585
R236 B.n921 B.n70 585
R237 B.n961 B.n70 585
R238 B.n920 B.n69 585
R239 B.n962 B.n69 585
R240 B.n919 B.n68 585
R241 B.n963 B.n68 585
R242 B.n918 B.n917 585
R243 B.n917 B.n64 585
R244 B.n916 B.n63 585
R245 B.n969 B.n63 585
R246 B.n915 B.n62 585
R247 B.n970 B.n62 585
R248 B.n914 B.n61 585
R249 B.n971 B.n61 585
R250 B.n913 B.n912 585
R251 B.n912 B.n57 585
R252 B.n911 B.n56 585
R253 B.n977 B.n56 585
R254 B.n910 B.n55 585
R255 B.n978 B.n55 585
R256 B.n909 B.n54 585
R257 B.n979 B.n54 585
R258 B.n908 B.n907 585
R259 B.n907 B.n53 585
R260 B.n906 B.n49 585
R261 B.n985 B.n49 585
R262 B.n905 B.n48 585
R263 B.n986 B.n48 585
R264 B.n904 B.n47 585
R265 B.n987 B.n47 585
R266 B.n903 B.n902 585
R267 B.n902 B.n43 585
R268 B.n901 B.n42 585
R269 B.n993 B.n42 585
R270 B.n900 B.n41 585
R271 B.n994 B.n41 585
R272 B.n899 B.n40 585
R273 B.n995 B.n40 585
R274 B.n898 B.n897 585
R275 B.n897 B.n36 585
R276 B.n896 B.n35 585
R277 B.n1001 B.n35 585
R278 B.n895 B.n34 585
R279 B.n1002 B.n34 585
R280 B.n894 B.n33 585
R281 B.n1003 B.n33 585
R282 B.n893 B.n892 585
R283 B.n892 B.n29 585
R284 B.n891 B.n28 585
R285 B.n1009 B.n28 585
R286 B.n890 B.n27 585
R287 B.n1010 B.n27 585
R288 B.n889 B.n26 585
R289 B.n1011 B.n26 585
R290 B.n888 B.n887 585
R291 B.n887 B.n22 585
R292 B.n886 B.n21 585
R293 B.n1017 B.n21 585
R294 B.n885 B.n20 585
R295 B.n1018 B.n20 585
R296 B.n884 B.n19 585
R297 B.n1019 B.n19 585
R298 B.n883 B.n882 585
R299 B.n882 B.n18 585
R300 B.n881 B.n14 585
R301 B.n1025 B.n14 585
R302 B.n880 B.n13 585
R303 B.n1026 B.n13 585
R304 B.n879 B.n12 585
R305 B.n1027 B.n12 585
R306 B.n878 B.n877 585
R307 B.n877 B.n8 585
R308 B.n876 B.n7 585
R309 B.n1033 B.n7 585
R310 B.n875 B.n6 585
R311 B.n1034 B.n6 585
R312 B.n874 B.n5 585
R313 B.n1035 B.n5 585
R314 B.n873 B.n872 585
R315 B.n872 B.n4 585
R316 B.n871 B.n361 585
R317 B.n871 B.n870 585
R318 B.n861 B.n362 585
R319 B.n363 B.n362 585
R320 B.n863 B.n862 585
R321 B.n864 B.n863 585
R322 B.n860 B.n368 585
R323 B.n368 B.n367 585
R324 B.n859 B.n858 585
R325 B.n858 B.n857 585
R326 B.n370 B.n369 585
R327 B.n850 B.n370 585
R328 B.n849 B.n848 585
R329 B.n851 B.n849 585
R330 B.n847 B.n375 585
R331 B.n375 B.n374 585
R332 B.n846 B.n845 585
R333 B.n845 B.n844 585
R334 B.n377 B.n376 585
R335 B.n378 B.n377 585
R336 B.n837 B.n836 585
R337 B.n838 B.n837 585
R338 B.n835 B.n383 585
R339 B.n383 B.n382 585
R340 B.n834 B.n833 585
R341 B.n833 B.n832 585
R342 B.n385 B.n384 585
R343 B.n386 B.n385 585
R344 B.n825 B.n824 585
R345 B.n826 B.n825 585
R346 B.n823 B.n390 585
R347 B.n394 B.n390 585
R348 B.n822 B.n821 585
R349 B.n821 B.n820 585
R350 B.n392 B.n391 585
R351 B.n393 B.n392 585
R352 B.n813 B.n812 585
R353 B.n814 B.n813 585
R354 B.n811 B.n399 585
R355 B.n399 B.n398 585
R356 B.n810 B.n809 585
R357 B.n809 B.n808 585
R358 B.n401 B.n400 585
R359 B.n402 B.n401 585
R360 B.n801 B.n800 585
R361 B.n802 B.n801 585
R362 B.n799 B.n407 585
R363 B.n407 B.n406 585
R364 B.n798 B.n797 585
R365 B.n797 B.n796 585
R366 B.n409 B.n408 585
R367 B.n789 B.n409 585
R368 B.n788 B.n787 585
R369 B.n790 B.n788 585
R370 B.n786 B.n414 585
R371 B.n414 B.n413 585
R372 B.n785 B.n784 585
R373 B.n784 B.n783 585
R374 B.n416 B.n415 585
R375 B.n417 B.n416 585
R376 B.n776 B.n775 585
R377 B.n777 B.n776 585
R378 B.n774 B.n422 585
R379 B.n422 B.n421 585
R380 B.n773 B.n772 585
R381 B.n772 B.n771 585
R382 B.n424 B.n423 585
R383 B.n425 B.n424 585
R384 B.n764 B.n763 585
R385 B.n765 B.n764 585
R386 B.n762 B.n430 585
R387 B.n430 B.n429 585
R388 B.n761 B.n760 585
R389 B.n760 B.n759 585
R390 B.n432 B.n431 585
R391 B.n433 B.n432 585
R392 B.n752 B.n751 585
R393 B.n753 B.n752 585
R394 B.n750 B.n438 585
R395 B.n438 B.n437 585
R396 B.n749 B.n748 585
R397 B.n748 B.n747 585
R398 B.n440 B.n439 585
R399 B.n441 B.n440 585
R400 B.n740 B.n739 585
R401 B.n741 B.n740 585
R402 B.n738 B.n446 585
R403 B.n446 B.n445 585
R404 B.n737 B.n736 585
R405 B.n736 B.n735 585
R406 B.n448 B.n447 585
R407 B.n449 B.n448 585
R408 B.n728 B.n727 585
R409 B.n729 B.n728 585
R410 B.n452 B.n451 585
R411 B.n515 B.n514 585
R412 B.n516 B.n512 585
R413 B.n512 B.n453 585
R414 B.n518 B.n517 585
R415 B.n520 B.n511 585
R416 B.n523 B.n522 585
R417 B.n524 B.n510 585
R418 B.n526 B.n525 585
R419 B.n528 B.n509 585
R420 B.n531 B.n530 585
R421 B.n532 B.n508 585
R422 B.n534 B.n533 585
R423 B.n536 B.n507 585
R424 B.n539 B.n538 585
R425 B.n540 B.n506 585
R426 B.n542 B.n541 585
R427 B.n544 B.n505 585
R428 B.n547 B.n546 585
R429 B.n548 B.n504 585
R430 B.n550 B.n549 585
R431 B.n552 B.n503 585
R432 B.n555 B.n554 585
R433 B.n556 B.n502 585
R434 B.n558 B.n557 585
R435 B.n560 B.n501 585
R436 B.n563 B.n562 585
R437 B.n564 B.n500 585
R438 B.n566 B.n565 585
R439 B.n568 B.n499 585
R440 B.n571 B.n570 585
R441 B.n572 B.n498 585
R442 B.n574 B.n573 585
R443 B.n576 B.n497 585
R444 B.n579 B.n578 585
R445 B.n580 B.n496 585
R446 B.n582 B.n581 585
R447 B.n584 B.n495 585
R448 B.n587 B.n586 585
R449 B.n588 B.n494 585
R450 B.n590 B.n589 585
R451 B.n592 B.n493 585
R452 B.n595 B.n594 585
R453 B.n596 B.n492 585
R454 B.n598 B.n597 585
R455 B.n600 B.n491 585
R456 B.n603 B.n602 585
R457 B.n604 B.n490 585
R458 B.n606 B.n605 585
R459 B.n608 B.n489 585
R460 B.n611 B.n610 585
R461 B.n612 B.n485 585
R462 B.n614 B.n613 585
R463 B.n616 B.n484 585
R464 B.n619 B.n618 585
R465 B.n620 B.n483 585
R466 B.n622 B.n621 585
R467 B.n624 B.n482 585
R468 B.n627 B.n626 585
R469 B.n628 B.n479 585
R470 B.n631 B.n630 585
R471 B.n633 B.n478 585
R472 B.n636 B.n635 585
R473 B.n637 B.n477 585
R474 B.n639 B.n638 585
R475 B.n641 B.n476 585
R476 B.n644 B.n643 585
R477 B.n645 B.n475 585
R478 B.n647 B.n646 585
R479 B.n649 B.n474 585
R480 B.n652 B.n651 585
R481 B.n653 B.n473 585
R482 B.n655 B.n654 585
R483 B.n657 B.n472 585
R484 B.n660 B.n659 585
R485 B.n661 B.n471 585
R486 B.n663 B.n662 585
R487 B.n665 B.n470 585
R488 B.n668 B.n667 585
R489 B.n669 B.n469 585
R490 B.n671 B.n670 585
R491 B.n673 B.n468 585
R492 B.n676 B.n675 585
R493 B.n677 B.n467 585
R494 B.n679 B.n678 585
R495 B.n681 B.n466 585
R496 B.n684 B.n683 585
R497 B.n685 B.n465 585
R498 B.n687 B.n686 585
R499 B.n689 B.n464 585
R500 B.n692 B.n691 585
R501 B.n693 B.n463 585
R502 B.n695 B.n694 585
R503 B.n697 B.n462 585
R504 B.n700 B.n699 585
R505 B.n701 B.n461 585
R506 B.n703 B.n702 585
R507 B.n705 B.n460 585
R508 B.n708 B.n707 585
R509 B.n709 B.n459 585
R510 B.n711 B.n710 585
R511 B.n713 B.n458 585
R512 B.n716 B.n715 585
R513 B.n717 B.n457 585
R514 B.n719 B.n718 585
R515 B.n721 B.n456 585
R516 B.n722 B.n455 585
R517 B.n725 B.n724 585
R518 B.n726 B.n454 585
R519 B.n454 B.n453 585
R520 B.n731 B.n730 585
R521 B.n730 B.n729 585
R522 B.n732 B.n450 585
R523 B.n450 B.n449 585
R524 B.n734 B.n733 585
R525 B.n735 B.n734 585
R526 B.n444 B.n443 585
R527 B.n445 B.n444 585
R528 B.n743 B.n742 585
R529 B.n742 B.n741 585
R530 B.n744 B.n442 585
R531 B.n442 B.n441 585
R532 B.n746 B.n745 585
R533 B.n747 B.n746 585
R534 B.n436 B.n435 585
R535 B.n437 B.n436 585
R536 B.n755 B.n754 585
R537 B.n754 B.n753 585
R538 B.n756 B.n434 585
R539 B.n434 B.n433 585
R540 B.n758 B.n757 585
R541 B.n759 B.n758 585
R542 B.n428 B.n427 585
R543 B.n429 B.n428 585
R544 B.n767 B.n766 585
R545 B.n766 B.n765 585
R546 B.n768 B.n426 585
R547 B.n426 B.n425 585
R548 B.n770 B.n769 585
R549 B.n771 B.n770 585
R550 B.n420 B.n419 585
R551 B.n421 B.n420 585
R552 B.n779 B.n778 585
R553 B.n778 B.n777 585
R554 B.n780 B.n418 585
R555 B.n418 B.n417 585
R556 B.n782 B.n781 585
R557 B.n783 B.n782 585
R558 B.n412 B.n411 585
R559 B.n413 B.n412 585
R560 B.n792 B.n791 585
R561 B.n791 B.n790 585
R562 B.n793 B.n410 585
R563 B.n789 B.n410 585
R564 B.n795 B.n794 585
R565 B.n796 B.n795 585
R566 B.n405 B.n404 585
R567 B.n406 B.n405 585
R568 B.n804 B.n803 585
R569 B.n803 B.n802 585
R570 B.n805 B.n403 585
R571 B.n403 B.n402 585
R572 B.n807 B.n806 585
R573 B.n808 B.n807 585
R574 B.n397 B.n396 585
R575 B.n398 B.n397 585
R576 B.n816 B.n815 585
R577 B.n815 B.n814 585
R578 B.n817 B.n395 585
R579 B.n395 B.n393 585
R580 B.n819 B.n818 585
R581 B.n820 B.n819 585
R582 B.n389 B.n388 585
R583 B.n394 B.n389 585
R584 B.n828 B.n827 585
R585 B.n827 B.n826 585
R586 B.n829 B.n387 585
R587 B.n387 B.n386 585
R588 B.n831 B.n830 585
R589 B.n832 B.n831 585
R590 B.n381 B.n380 585
R591 B.n382 B.n381 585
R592 B.n840 B.n839 585
R593 B.n839 B.n838 585
R594 B.n841 B.n379 585
R595 B.n379 B.n378 585
R596 B.n843 B.n842 585
R597 B.n844 B.n843 585
R598 B.n373 B.n372 585
R599 B.n374 B.n373 585
R600 B.n853 B.n852 585
R601 B.n852 B.n851 585
R602 B.n854 B.n371 585
R603 B.n850 B.n371 585
R604 B.n856 B.n855 585
R605 B.n857 B.n856 585
R606 B.n366 B.n365 585
R607 B.n367 B.n366 585
R608 B.n866 B.n865 585
R609 B.n865 B.n864 585
R610 B.n867 B.n364 585
R611 B.n364 B.n363 585
R612 B.n869 B.n868 585
R613 B.n870 B.n869 585
R614 B.n2 B.n0 585
R615 B.n4 B.n2 585
R616 B.n3 B.n1 585
R617 B.n1034 B.n3 585
R618 B.n1032 B.n1031 585
R619 B.n1033 B.n1032 585
R620 B.n1030 B.n9 585
R621 B.n9 B.n8 585
R622 B.n1029 B.n1028 585
R623 B.n1028 B.n1027 585
R624 B.n11 B.n10 585
R625 B.n1026 B.n11 585
R626 B.n1024 B.n1023 585
R627 B.n1025 B.n1024 585
R628 B.n1022 B.n15 585
R629 B.n18 B.n15 585
R630 B.n1021 B.n1020 585
R631 B.n1020 B.n1019 585
R632 B.n17 B.n16 585
R633 B.n1018 B.n17 585
R634 B.n1016 B.n1015 585
R635 B.n1017 B.n1016 585
R636 B.n1014 B.n23 585
R637 B.n23 B.n22 585
R638 B.n1013 B.n1012 585
R639 B.n1012 B.n1011 585
R640 B.n25 B.n24 585
R641 B.n1010 B.n25 585
R642 B.n1008 B.n1007 585
R643 B.n1009 B.n1008 585
R644 B.n1006 B.n30 585
R645 B.n30 B.n29 585
R646 B.n1005 B.n1004 585
R647 B.n1004 B.n1003 585
R648 B.n32 B.n31 585
R649 B.n1002 B.n32 585
R650 B.n1000 B.n999 585
R651 B.n1001 B.n1000 585
R652 B.n998 B.n37 585
R653 B.n37 B.n36 585
R654 B.n997 B.n996 585
R655 B.n996 B.n995 585
R656 B.n39 B.n38 585
R657 B.n994 B.n39 585
R658 B.n992 B.n991 585
R659 B.n993 B.n992 585
R660 B.n990 B.n44 585
R661 B.n44 B.n43 585
R662 B.n989 B.n988 585
R663 B.n988 B.n987 585
R664 B.n46 B.n45 585
R665 B.n986 B.n46 585
R666 B.n984 B.n983 585
R667 B.n985 B.n984 585
R668 B.n982 B.n50 585
R669 B.n53 B.n50 585
R670 B.n981 B.n980 585
R671 B.n980 B.n979 585
R672 B.n52 B.n51 585
R673 B.n978 B.n52 585
R674 B.n976 B.n975 585
R675 B.n977 B.n976 585
R676 B.n974 B.n58 585
R677 B.n58 B.n57 585
R678 B.n973 B.n972 585
R679 B.n972 B.n971 585
R680 B.n60 B.n59 585
R681 B.n970 B.n60 585
R682 B.n968 B.n967 585
R683 B.n969 B.n968 585
R684 B.n966 B.n65 585
R685 B.n65 B.n64 585
R686 B.n965 B.n964 585
R687 B.n964 B.n963 585
R688 B.n67 B.n66 585
R689 B.n962 B.n67 585
R690 B.n960 B.n959 585
R691 B.n961 B.n960 585
R692 B.n958 B.n72 585
R693 B.n72 B.n71 585
R694 B.n957 B.n956 585
R695 B.n956 B.n955 585
R696 B.n74 B.n73 585
R697 B.n954 B.n74 585
R698 B.n952 B.n951 585
R699 B.n953 B.n952 585
R700 B.n950 B.n79 585
R701 B.n79 B.n78 585
R702 B.n949 B.n948 585
R703 B.n948 B.n947 585
R704 B.n81 B.n80 585
R705 B.n946 B.n81 585
R706 B.n944 B.n943 585
R707 B.n945 B.n944 585
R708 B.n942 B.n86 585
R709 B.n86 B.n85 585
R710 B.n941 B.n940 585
R711 B.n940 B.n939 585
R712 B.n1037 B.n1036 585
R713 B.n1036 B.n1035 585
R714 B.n730 B.n452 521.33
R715 B.n940 B.n88 521.33
R716 B.n728 B.n454 521.33
R717 B.n936 B.n89 521.33
R718 B.n480 B.t17 322.522
R719 B.n486 B.t13 322.522
R720 B.n146 B.t6 322.522
R721 B.n144 B.t10 322.522
R722 B.n938 B.n937 256.663
R723 B.n938 B.n142 256.663
R724 B.n938 B.n141 256.663
R725 B.n938 B.n140 256.663
R726 B.n938 B.n139 256.663
R727 B.n938 B.n138 256.663
R728 B.n938 B.n137 256.663
R729 B.n938 B.n136 256.663
R730 B.n938 B.n135 256.663
R731 B.n938 B.n134 256.663
R732 B.n938 B.n133 256.663
R733 B.n938 B.n132 256.663
R734 B.n938 B.n131 256.663
R735 B.n938 B.n130 256.663
R736 B.n938 B.n129 256.663
R737 B.n938 B.n128 256.663
R738 B.n938 B.n127 256.663
R739 B.n938 B.n126 256.663
R740 B.n938 B.n125 256.663
R741 B.n938 B.n124 256.663
R742 B.n938 B.n123 256.663
R743 B.n938 B.n122 256.663
R744 B.n938 B.n121 256.663
R745 B.n938 B.n120 256.663
R746 B.n938 B.n119 256.663
R747 B.n938 B.n118 256.663
R748 B.n938 B.n117 256.663
R749 B.n938 B.n116 256.663
R750 B.n938 B.n115 256.663
R751 B.n938 B.n114 256.663
R752 B.n938 B.n113 256.663
R753 B.n938 B.n112 256.663
R754 B.n938 B.n111 256.663
R755 B.n938 B.n110 256.663
R756 B.n938 B.n109 256.663
R757 B.n938 B.n108 256.663
R758 B.n938 B.n107 256.663
R759 B.n938 B.n106 256.663
R760 B.n938 B.n105 256.663
R761 B.n938 B.n104 256.663
R762 B.n938 B.n103 256.663
R763 B.n938 B.n102 256.663
R764 B.n938 B.n101 256.663
R765 B.n938 B.n100 256.663
R766 B.n938 B.n99 256.663
R767 B.n938 B.n98 256.663
R768 B.n938 B.n97 256.663
R769 B.n938 B.n96 256.663
R770 B.n938 B.n95 256.663
R771 B.n938 B.n94 256.663
R772 B.n938 B.n93 256.663
R773 B.n938 B.n92 256.663
R774 B.n938 B.n91 256.663
R775 B.n938 B.n90 256.663
R776 B.n513 B.n453 256.663
R777 B.n519 B.n453 256.663
R778 B.n521 B.n453 256.663
R779 B.n527 B.n453 256.663
R780 B.n529 B.n453 256.663
R781 B.n535 B.n453 256.663
R782 B.n537 B.n453 256.663
R783 B.n543 B.n453 256.663
R784 B.n545 B.n453 256.663
R785 B.n551 B.n453 256.663
R786 B.n553 B.n453 256.663
R787 B.n559 B.n453 256.663
R788 B.n561 B.n453 256.663
R789 B.n567 B.n453 256.663
R790 B.n569 B.n453 256.663
R791 B.n575 B.n453 256.663
R792 B.n577 B.n453 256.663
R793 B.n583 B.n453 256.663
R794 B.n585 B.n453 256.663
R795 B.n591 B.n453 256.663
R796 B.n593 B.n453 256.663
R797 B.n599 B.n453 256.663
R798 B.n601 B.n453 256.663
R799 B.n607 B.n453 256.663
R800 B.n609 B.n453 256.663
R801 B.n615 B.n453 256.663
R802 B.n617 B.n453 256.663
R803 B.n623 B.n453 256.663
R804 B.n625 B.n453 256.663
R805 B.n632 B.n453 256.663
R806 B.n634 B.n453 256.663
R807 B.n640 B.n453 256.663
R808 B.n642 B.n453 256.663
R809 B.n648 B.n453 256.663
R810 B.n650 B.n453 256.663
R811 B.n656 B.n453 256.663
R812 B.n658 B.n453 256.663
R813 B.n664 B.n453 256.663
R814 B.n666 B.n453 256.663
R815 B.n672 B.n453 256.663
R816 B.n674 B.n453 256.663
R817 B.n680 B.n453 256.663
R818 B.n682 B.n453 256.663
R819 B.n688 B.n453 256.663
R820 B.n690 B.n453 256.663
R821 B.n696 B.n453 256.663
R822 B.n698 B.n453 256.663
R823 B.n704 B.n453 256.663
R824 B.n706 B.n453 256.663
R825 B.n712 B.n453 256.663
R826 B.n714 B.n453 256.663
R827 B.n720 B.n453 256.663
R828 B.n723 B.n453 256.663
R829 B.n730 B.n450 163.367
R830 B.n734 B.n450 163.367
R831 B.n734 B.n444 163.367
R832 B.n742 B.n444 163.367
R833 B.n742 B.n442 163.367
R834 B.n746 B.n442 163.367
R835 B.n746 B.n436 163.367
R836 B.n754 B.n436 163.367
R837 B.n754 B.n434 163.367
R838 B.n758 B.n434 163.367
R839 B.n758 B.n428 163.367
R840 B.n766 B.n428 163.367
R841 B.n766 B.n426 163.367
R842 B.n770 B.n426 163.367
R843 B.n770 B.n420 163.367
R844 B.n778 B.n420 163.367
R845 B.n778 B.n418 163.367
R846 B.n782 B.n418 163.367
R847 B.n782 B.n412 163.367
R848 B.n791 B.n412 163.367
R849 B.n791 B.n410 163.367
R850 B.n795 B.n410 163.367
R851 B.n795 B.n405 163.367
R852 B.n803 B.n405 163.367
R853 B.n803 B.n403 163.367
R854 B.n807 B.n403 163.367
R855 B.n807 B.n397 163.367
R856 B.n815 B.n397 163.367
R857 B.n815 B.n395 163.367
R858 B.n819 B.n395 163.367
R859 B.n819 B.n389 163.367
R860 B.n827 B.n389 163.367
R861 B.n827 B.n387 163.367
R862 B.n831 B.n387 163.367
R863 B.n831 B.n381 163.367
R864 B.n839 B.n381 163.367
R865 B.n839 B.n379 163.367
R866 B.n843 B.n379 163.367
R867 B.n843 B.n373 163.367
R868 B.n852 B.n373 163.367
R869 B.n852 B.n371 163.367
R870 B.n856 B.n371 163.367
R871 B.n856 B.n366 163.367
R872 B.n865 B.n366 163.367
R873 B.n865 B.n364 163.367
R874 B.n869 B.n364 163.367
R875 B.n869 B.n2 163.367
R876 B.n1036 B.n2 163.367
R877 B.n1036 B.n3 163.367
R878 B.n1032 B.n3 163.367
R879 B.n1032 B.n9 163.367
R880 B.n1028 B.n9 163.367
R881 B.n1028 B.n11 163.367
R882 B.n1024 B.n11 163.367
R883 B.n1024 B.n15 163.367
R884 B.n1020 B.n15 163.367
R885 B.n1020 B.n17 163.367
R886 B.n1016 B.n17 163.367
R887 B.n1016 B.n23 163.367
R888 B.n1012 B.n23 163.367
R889 B.n1012 B.n25 163.367
R890 B.n1008 B.n25 163.367
R891 B.n1008 B.n30 163.367
R892 B.n1004 B.n30 163.367
R893 B.n1004 B.n32 163.367
R894 B.n1000 B.n32 163.367
R895 B.n1000 B.n37 163.367
R896 B.n996 B.n37 163.367
R897 B.n996 B.n39 163.367
R898 B.n992 B.n39 163.367
R899 B.n992 B.n44 163.367
R900 B.n988 B.n44 163.367
R901 B.n988 B.n46 163.367
R902 B.n984 B.n46 163.367
R903 B.n984 B.n50 163.367
R904 B.n980 B.n50 163.367
R905 B.n980 B.n52 163.367
R906 B.n976 B.n52 163.367
R907 B.n976 B.n58 163.367
R908 B.n972 B.n58 163.367
R909 B.n972 B.n60 163.367
R910 B.n968 B.n60 163.367
R911 B.n968 B.n65 163.367
R912 B.n964 B.n65 163.367
R913 B.n964 B.n67 163.367
R914 B.n960 B.n67 163.367
R915 B.n960 B.n72 163.367
R916 B.n956 B.n72 163.367
R917 B.n956 B.n74 163.367
R918 B.n952 B.n74 163.367
R919 B.n952 B.n79 163.367
R920 B.n948 B.n79 163.367
R921 B.n948 B.n81 163.367
R922 B.n944 B.n81 163.367
R923 B.n944 B.n86 163.367
R924 B.n940 B.n86 163.367
R925 B.n514 B.n512 163.367
R926 B.n518 B.n512 163.367
R927 B.n522 B.n520 163.367
R928 B.n526 B.n510 163.367
R929 B.n530 B.n528 163.367
R930 B.n534 B.n508 163.367
R931 B.n538 B.n536 163.367
R932 B.n542 B.n506 163.367
R933 B.n546 B.n544 163.367
R934 B.n550 B.n504 163.367
R935 B.n554 B.n552 163.367
R936 B.n558 B.n502 163.367
R937 B.n562 B.n560 163.367
R938 B.n566 B.n500 163.367
R939 B.n570 B.n568 163.367
R940 B.n574 B.n498 163.367
R941 B.n578 B.n576 163.367
R942 B.n582 B.n496 163.367
R943 B.n586 B.n584 163.367
R944 B.n590 B.n494 163.367
R945 B.n594 B.n592 163.367
R946 B.n598 B.n492 163.367
R947 B.n602 B.n600 163.367
R948 B.n606 B.n490 163.367
R949 B.n610 B.n608 163.367
R950 B.n614 B.n485 163.367
R951 B.n618 B.n616 163.367
R952 B.n622 B.n483 163.367
R953 B.n626 B.n624 163.367
R954 B.n631 B.n479 163.367
R955 B.n635 B.n633 163.367
R956 B.n639 B.n477 163.367
R957 B.n643 B.n641 163.367
R958 B.n647 B.n475 163.367
R959 B.n651 B.n649 163.367
R960 B.n655 B.n473 163.367
R961 B.n659 B.n657 163.367
R962 B.n663 B.n471 163.367
R963 B.n667 B.n665 163.367
R964 B.n671 B.n469 163.367
R965 B.n675 B.n673 163.367
R966 B.n679 B.n467 163.367
R967 B.n683 B.n681 163.367
R968 B.n687 B.n465 163.367
R969 B.n691 B.n689 163.367
R970 B.n695 B.n463 163.367
R971 B.n699 B.n697 163.367
R972 B.n703 B.n461 163.367
R973 B.n707 B.n705 163.367
R974 B.n711 B.n459 163.367
R975 B.n715 B.n713 163.367
R976 B.n719 B.n457 163.367
R977 B.n722 B.n721 163.367
R978 B.n724 B.n454 163.367
R979 B.n728 B.n448 163.367
R980 B.n736 B.n448 163.367
R981 B.n736 B.n446 163.367
R982 B.n740 B.n446 163.367
R983 B.n740 B.n440 163.367
R984 B.n748 B.n440 163.367
R985 B.n748 B.n438 163.367
R986 B.n752 B.n438 163.367
R987 B.n752 B.n432 163.367
R988 B.n760 B.n432 163.367
R989 B.n760 B.n430 163.367
R990 B.n764 B.n430 163.367
R991 B.n764 B.n424 163.367
R992 B.n772 B.n424 163.367
R993 B.n772 B.n422 163.367
R994 B.n776 B.n422 163.367
R995 B.n776 B.n416 163.367
R996 B.n784 B.n416 163.367
R997 B.n784 B.n414 163.367
R998 B.n788 B.n414 163.367
R999 B.n788 B.n409 163.367
R1000 B.n797 B.n409 163.367
R1001 B.n797 B.n407 163.367
R1002 B.n801 B.n407 163.367
R1003 B.n801 B.n401 163.367
R1004 B.n809 B.n401 163.367
R1005 B.n809 B.n399 163.367
R1006 B.n813 B.n399 163.367
R1007 B.n813 B.n392 163.367
R1008 B.n821 B.n392 163.367
R1009 B.n821 B.n390 163.367
R1010 B.n825 B.n390 163.367
R1011 B.n825 B.n385 163.367
R1012 B.n833 B.n385 163.367
R1013 B.n833 B.n383 163.367
R1014 B.n837 B.n383 163.367
R1015 B.n837 B.n377 163.367
R1016 B.n845 B.n377 163.367
R1017 B.n845 B.n375 163.367
R1018 B.n849 B.n375 163.367
R1019 B.n849 B.n370 163.367
R1020 B.n858 B.n370 163.367
R1021 B.n858 B.n368 163.367
R1022 B.n863 B.n368 163.367
R1023 B.n863 B.n362 163.367
R1024 B.n871 B.n362 163.367
R1025 B.n872 B.n871 163.367
R1026 B.n872 B.n5 163.367
R1027 B.n6 B.n5 163.367
R1028 B.n7 B.n6 163.367
R1029 B.n877 B.n7 163.367
R1030 B.n877 B.n12 163.367
R1031 B.n13 B.n12 163.367
R1032 B.n14 B.n13 163.367
R1033 B.n882 B.n14 163.367
R1034 B.n882 B.n19 163.367
R1035 B.n20 B.n19 163.367
R1036 B.n21 B.n20 163.367
R1037 B.n887 B.n21 163.367
R1038 B.n887 B.n26 163.367
R1039 B.n27 B.n26 163.367
R1040 B.n28 B.n27 163.367
R1041 B.n892 B.n28 163.367
R1042 B.n892 B.n33 163.367
R1043 B.n34 B.n33 163.367
R1044 B.n35 B.n34 163.367
R1045 B.n897 B.n35 163.367
R1046 B.n897 B.n40 163.367
R1047 B.n41 B.n40 163.367
R1048 B.n42 B.n41 163.367
R1049 B.n902 B.n42 163.367
R1050 B.n902 B.n47 163.367
R1051 B.n48 B.n47 163.367
R1052 B.n49 B.n48 163.367
R1053 B.n907 B.n49 163.367
R1054 B.n907 B.n54 163.367
R1055 B.n55 B.n54 163.367
R1056 B.n56 B.n55 163.367
R1057 B.n912 B.n56 163.367
R1058 B.n912 B.n61 163.367
R1059 B.n62 B.n61 163.367
R1060 B.n63 B.n62 163.367
R1061 B.n917 B.n63 163.367
R1062 B.n917 B.n68 163.367
R1063 B.n69 B.n68 163.367
R1064 B.n70 B.n69 163.367
R1065 B.n922 B.n70 163.367
R1066 B.n922 B.n75 163.367
R1067 B.n76 B.n75 163.367
R1068 B.n77 B.n76 163.367
R1069 B.n927 B.n77 163.367
R1070 B.n927 B.n82 163.367
R1071 B.n83 B.n82 163.367
R1072 B.n84 B.n83 163.367
R1073 B.n932 B.n84 163.367
R1074 B.n932 B.n89 163.367
R1075 B.n150 B.n149 163.367
R1076 B.n154 B.n153 163.367
R1077 B.n158 B.n157 163.367
R1078 B.n162 B.n161 163.367
R1079 B.n166 B.n165 163.367
R1080 B.n170 B.n169 163.367
R1081 B.n174 B.n173 163.367
R1082 B.n178 B.n177 163.367
R1083 B.n182 B.n181 163.367
R1084 B.n186 B.n185 163.367
R1085 B.n190 B.n189 163.367
R1086 B.n194 B.n193 163.367
R1087 B.n198 B.n197 163.367
R1088 B.n202 B.n201 163.367
R1089 B.n206 B.n205 163.367
R1090 B.n210 B.n209 163.367
R1091 B.n214 B.n213 163.367
R1092 B.n218 B.n217 163.367
R1093 B.n222 B.n221 163.367
R1094 B.n226 B.n225 163.367
R1095 B.n230 B.n229 163.367
R1096 B.n234 B.n233 163.367
R1097 B.n238 B.n237 163.367
R1098 B.n242 B.n241 163.367
R1099 B.n247 B.n246 163.367
R1100 B.n251 B.n250 163.367
R1101 B.n255 B.n254 163.367
R1102 B.n259 B.n258 163.367
R1103 B.n263 B.n262 163.367
R1104 B.n268 B.n267 163.367
R1105 B.n272 B.n271 163.367
R1106 B.n276 B.n275 163.367
R1107 B.n280 B.n279 163.367
R1108 B.n284 B.n283 163.367
R1109 B.n288 B.n287 163.367
R1110 B.n292 B.n291 163.367
R1111 B.n296 B.n295 163.367
R1112 B.n300 B.n299 163.367
R1113 B.n304 B.n303 163.367
R1114 B.n308 B.n307 163.367
R1115 B.n312 B.n311 163.367
R1116 B.n316 B.n315 163.367
R1117 B.n320 B.n319 163.367
R1118 B.n324 B.n323 163.367
R1119 B.n328 B.n327 163.367
R1120 B.n332 B.n331 163.367
R1121 B.n336 B.n335 163.367
R1122 B.n340 B.n339 163.367
R1123 B.n344 B.n343 163.367
R1124 B.n348 B.n347 163.367
R1125 B.n352 B.n351 163.367
R1126 B.n356 B.n355 163.367
R1127 B.n358 B.n143 163.367
R1128 B.n480 B.t19 138.874
R1129 B.n144 B.t11 138.874
R1130 B.n486 B.t16 138.856
R1131 B.n146 B.t8 138.856
R1132 B.n729 B.n453 77.1253
R1133 B.n939 B.n938 77.1253
R1134 B.n481 B.t18 72.7406
R1135 B.n145 B.t12 72.7406
R1136 B.n487 B.t15 72.7219
R1137 B.n147 B.t9 72.7219
R1138 B.n513 B.n452 71.676
R1139 B.n519 B.n518 71.676
R1140 B.n522 B.n521 71.676
R1141 B.n527 B.n526 71.676
R1142 B.n530 B.n529 71.676
R1143 B.n535 B.n534 71.676
R1144 B.n538 B.n537 71.676
R1145 B.n543 B.n542 71.676
R1146 B.n546 B.n545 71.676
R1147 B.n551 B.n550 71.676
R1148 B.n554 B.n553 71.676
R1149 B.n559 B.n558 71.676
R1150 B.n562 B.n561 71.676
R1151 B.n567 B.n566 71.676
R1152 B.n570 B.n569 71.676
R1153 B.n575 B.n574 71.676
R1154 B.n578 B.n577 71.676
R1155 B.n583 B.n582 71.676
R1156 B.n586 B.n585 71.676
R1157 B.n591 B.n590 71.676
R1158 B.n594 B.n593 71.676
R1159 B.n599 B.n598 71.676
R1160 B.n602 B.n601 71.676
R1161 B.n607 B.n606 71.676
R1162 B.n610 B.n609 71.676
R1163 B.n615 B.n614 71.676
R1164 B.n618 B.n617 71.676
R1165 B.n623 B.n622 71.676
R1166 B.n626 B.n625 71.676
R1167 B.n632 B.n631 71.676
R1168 B.n635 B.n634 71.676
R1169 B.n640 B.n639 71.676
R1170 B.n643 B.n642 71.676
R1171 B.n648 B.n647 71.676
R1172 B.n651 B.n650 71.676
R1173 B.n656 B.n655 71.676
R1174 B.n659 B.n658 71.676
R1175 B.n664 B.n663 71.676
R1176 B.n667 B.n666 71.676
R1177 B.n672 B.n671 71.676
R1178 B.n675 B.n674 71.676
R1179 B.n680 B.n679 71.676
R1180 B.n683 B.n682 71.676
R1181 B.n688 B.n687 71.676
R1182 B.n691 B.n690 71.676
R1183 B.n696 B.n695 71.676
R1184 B.n699 B.n698 71.676
R1185 B.n704 B.n703 71.676
R1186 B.n707 B.n706 71.676
R1187 B.n712 B.n711 71.676
R1188 B.n715 B.n714 71.676
R1189 B.n720 B.n719 71.676
R1190 B.n723 B.n722 71.676
R1191 B.n90 B.n88 71.676
R1192 B.n150 B.n91 71.676
R1193 B.n154 B.n92 71.676
R1194 B.n158 B.n93 71.676
R1195 B.n162 B.n94 71.676
R1196 B.n166 B.n95 71.676
R1197 B.n170 B.n96 71.676
R1198 B.n174 B.n97 71.676
R1199 B.n178 B.n98 71.676
R1200 B.n182 B.n99 71.676
R1201 B.n186 B.n100 71.676
R1202 B.n190 B.n101 71.676
R1203 B.n194 B.n102 71.676
R1204 B.n198 B.n103 71.676
R1205 B.n202 B.n104 71.676
R1206 B.n206 B.n105 71.676
R1207 B.n210 B.n106 71.676
R1208 B.n214 B.n107 71.676
R1209 B.n218 B.n108 71.676
R1210 B.n222 B.n109 71.676
R1211 B.n226 B.n110 71.676
R1212 B.n230 B.n111 71.676
R1213 B.n234 B.n112 71.676
R1214 B.n238 B.n113 71.676
R1215 B.n242 B.n114 71.676
R1216 B.n247 B.n115 71.676
R1217 B.n251 B.n116 71.676
R1218 B.n255 B.n117 71.676
R1219 B.n259 B.n118 71.676
R1220 B.n263 B.n119 71.676
R1221 B.n268 B.n120 71.676
R1222 B.n272 B.n121 71.676
R1223 B.n276 B.n122 71.676
R1224 B.n280 B.n123 71.676
R1225 B.n284 B.n124 71.676
R1226 B.n288 B.n125 71.676
R1227 B.n292 B.n126 71.676
R1228 B.n296 B.n127 71.676
R1229 B.n300 B.n128 71.676
R1230 B.n304 B.n129 71.676
R1231 B.n308 B.n130 71.676
R1232 B.n312 B.n131 71.676
R1233 B.n316 B.n132 71.676
R1234 B.n320 B.n133 71.676
R1235 B.n324 B.n134 71.676
R1236 B.n328 B.n135 71.676
R1237 B.n332 B.n136 71.676
R1238 B.n336 B.n137 71.676
R1239 B.n340 B.n138 71.676
R1240 B.n344 B.n139 71.676
R1241 B.n348 B.n140 71.676
R1242 B.n352 B.n141 71.676
R1243 B.n356 B.n142 71.676
R1244 B.n937 B.n143 71.676
R1245 B.n937 B.n936 71.676
R1246 B.n358 B.n142 71.676
R1247 B.n355 B.n141 71.676
R1248 B.n351 B.n140 71.676
R1249 B.n347 B.n139 71.676
R1250 B.n343 B.n138 71.676
R1251 B.n339 B.n137 71.676
R1252 B.n335 B.n136 71.676
R1253 B.n331 B.n135 71.676
R1254 B.n327 B.n134 71.676
R1255 B.n323 B.n133 71.676
R1256 B.n319 B.n132 71.676
R1257 B.n315 B.n131 71.676
R1258 B.n311 B.n130 71.676
R1259 B.n307 B.n129 71.676
R1260 B.n303 B.n128 71.676
R1261 B.n299 B.n127 71.676
R1262 B.n295 B.n126 71.676
R1263 B.n291 B.n125 71.676
R1264 B.n287 B.n124 71.676
R1265 B.n283 B.n123 71.676
R1266 B.n279 B.n122 71.676
R1267 B.n275 B.n121 71.676
R1268 B.n271 B.n120 71.676
R1269 B.n267 B.n119 71.676
R1270 B.n262 B.n118 71.676
R1271 B.n258 B.n117 71.676
R1272 B.n254 B.n116 71.676
R1273 B.n250 B.n115 71.676
R1274 B.n246 B.n114 71.676
R1275 B.n241 B.n113 71.676
R1276 B.n237 B.n112 71.676
R1277 B.n233 B.n111 71.676
R1278 B.n229 B.n110 71.676
R1279 B.n225 B.n109 71.676
R1280 B.n221 B.n108 71.676
R1281 B.n217 B.n107 71.676
R1282 B.n213 B.n106 71.676
R1283 B.n209 B.n105 71.676
R1284 B.n205 B.n104 71.676
R1285 B.n201 B.n103 71.676
R1286 B.n197 B.n102 71.676
R1287 B.n193 B.n101 71.676
R1288 B.n189 B.n100 71.676
R1289 B.n185 B.n99 71.676
R1290 B.n181 B.n98 71.676
R1291 B.n177 B.n97 71.676
R1292 B.n173 B.n96 71.676
R1293 B.n169 B.n95 71.676
R1294 B.n165 B.n94 71.676
R1295 B.n161 B.n93 71.676
R1296 B.n157 B.n92 71.676
R1297 B.n153 B.n91 71.676
R1298 B.n149 B.n90 71.676
R1299 B.n514 B.n513 71.676
R1300 B.n520 B.n519 71.676
R1301 B.n521 B.n510 71.676
R1302 B.n528 B.n527 71.676
R1303 B.n529 B.n508 71.676
R1304 B.n536 B.n535 71.676
R1305 B.n537 B.n506 71.676
R1306 B.n544 B.n543 71.676
R1307 B.n545 B.n504 71.676
R1308 B.n552 B.n551 71.676
R1309 B.n553 B.n502 71.676
R1310 B.n560 B.n559 71.676
R1311 B.n561 B.n500 71.676
R1312 B.n568 B.n567 71.676
R1313 B.n569 B.n498 71.676
R1314 B.n576 B.n575 71.676
R1315 B.n577 B.n496 71.676
R1316 B.n584 B.n583 71.676
R1317 B.n585 B.n494 71.676
R1318 B.n592 B.n591 71.676
R1319 B.n593 B.n492 71.676
R1320 B.n600 B.n599 71.676
R1321 B.n601 B.n490 71.676
R1322 B.n608 B.n607 71.676
R1323 B.n609 B.n485 71.676
R1324 B.n616 B.n615 71.676
R1325 B.n617 B.n483 71.676
R1326 B.n624 B.n623 71.676
R1327 B.n625 B.n479 71.676
R1328 B.n633 B.n632 71.676
R1329 B.n634 B.n477 71.676
R1330 B.n641 B.n640 71.676
R1331 B.n642 B.n475 71.676
R1332 B.n649 B.n648 71.676
R1333 B.n650 B.n473 71.676
R1334 B.n657 B.n656 71.676
R1335 B.n658 B.n471 71.676
R1336 B.n665 B.n664 71.676
R1337 B.n666 B.n469 71.676
R1338 B.n673 B.n672 71.676
R1339 B.n674 B.n467 71.676
R1340 B.n681 B.n680 71.676
R1341 B.n682 B.n465 71.676
R1342 B.n689 B.n688 71.676
R1343 B.n690 B.n463 71.676
R1344 B.n697 B.n696 71.676
R1345 B.n698 B.n461 71.676
R1346 B.n705 B.n704 71.676
R1347 B.n706 B.n459 71.676
R1348 B.n713 B.n712 71.676
R1349 B.n714 B.n457 71.676
R1350 B.n721 B.n720 71.676
R1351 B.n724 B.n723 71.676
R1352 B.n481 B.n480 66.1338
R1353 B.n487 B.n486 66.1338
R1354 B.n147 B.n146 66.1338
R1355 B.n145 B.n144 66.1338
R1356 B.n629 B.n481 59.5399
R1357 B.n488 B.n487 59.5399
R1358 B.n244 B.n147 59.5399
R1359 B.n265 B.n145 59.5399
R1360 B.n729 B.n449 37.7306
R1361 B.n735 B.n449 37.7306
R1362 B.n735 B.n445 37.7306
R1363 B.n741 B.n445 37.7306
R1364 B.n741 B.n441 37.7306
R1365 B.n747 B.n441 37.7306
R1366 B.n747 B.n437 37.7306
R1367 B.n753 B.n437 37.7306
R1368 B.n759 B.n433 37.7306
R1369 B.n759 B.n429 37.7306
R1370 B.n765 B.n429 37.7306
R1371 B.n765 B.n425 37.7306
R1372 B.n771 B.n425 37.7306
R1373 B.n771 B.n421 37.7306
R1374 B.n777 B.n421 37.7306
R1375 B.n777 B.n417 37.7306
R1376 B.n783 B.n417 37.7306
R1377 B.n783 B.n413 37.7306
R1378 B.n790 B.n413 37.7306
R1379 B.n790 B.n789 37.7306
R1380 B.n796 B.n406 37.7306
R1381 B.n802 B.n406 37.7306
R1382 B.n802 B.n402 37.7306
R1383 B.n808 B.n402 37.7306
R1384 B.n808 B.n398 37.7306
R1385 B.n814 B.n398 37.7306
R1386 B.n814 B.n393 37.7306
R1387 B.n820 B.n393 37.7306
R1388 B.n820 B.n394 37.7306
R1389 B.n826 B.n386 37.7306
R1390 B.n832 B.n386 37.7306
R1391 B.n832 B.n382 37.7306
R1392 B.n838 B.n382 37.7306
R1393 B.n838 B.n378 37.7306
R1394 B.n844 B.n378 37.7306
R1395 B.n844 B.n374 37.7306
R1396 B.n851 B.n374 37.7306
R1397 B.n851 B.n850 37.7306
R1398 B.n857 B.n367 37.7306
R1399 B.n864 B.n367 37.7306
R1400 B.n864 B.n363 37.7306
R1401 B.n870 B.n363 37.7306
R1402 B.n870 B.n4 37.7306
R1403 B.n1035 B.n4 37.7306
R1404 B.n1035 B.n1034 37.7306
R1405 B.n1034 B.n1033 37.7306
R1406 B.n1033 B.n8 37.7306
R1407 B.n1027 B.n8 37.7306
R1408 B.n1027 B.n1026 37.7306
R1409 B.n1026 B.n1025 37.7306
R1410 B.n1019 B.n18 37.7306
R1411 B.n1019 B.n1018 37.7306
R1412 B.n1018 B.n1017 37.7306
R1413 B.n1017 B.n22 37.7306
R1414 B.n1011 B.n22 37.7306
R1415 B.n1011 B.n1010 37.7306
R1416 B.n1010 B.n1009 37.7306
R1417 B.n1009 B.n29 37.7306
R1418 B.n1003 B.n29 37.7306
R1419 B.n1002 B.n1001 37.7306
R1420 B.n1001 B.n36 37.7306
R1421 B.n995 B.n36 37.7306
R1422 B.n995 B.n994 37.7306
R1423 B.n994 B.n993 37.7306
R1424 B.n993 B.n43 37.7306
R1425 B.n987 B.n43 37.7306
R1426 B.n987 B.n986 37.7306
R1427 B.n986 B.n985 37.7306
R1428 B.n979 B.n53 37.7306
R1429 B.n979 B.n978 37.7306
R1430 B.n978 B.n977 37.7306
R1431 B.n977 B.n57 37.7306
R1432 B.n971 B.n57 37.7306
R1433 B.n971 B.n970 37.7306
R1434 B.n970 B.n969 37.7306
R1435 B.n969 B.n64 37.7306
R1436 B.n963 B.n64 37.7306
R1437 B.n963 B.n962 37.7306
R1438 B.n962 B.n961 37.7306
R1439 B.n961 B.n71 37.7306
R1440 B.n955 B.n954 37.7306
R1441 B.n954 B.n953 37.7306
R1442 B.n953 B.n78 37.7306
R1443 B.n947 B.n78 37.7306
R1444 B.n947 B.n946 37.7306
R1445 B.n946 B.n945 37.7306
R1446 B.n945 B.n85 37.7306
R1447 B.n939 B.n85 37.7306
R1448 B.t14 B.n433 34.4015
R1449 B.t7 B.n71 34.4015
R1450 B.n941 B.n87 33.8737
R1451 B.n935 B.n934 33.8737
R1452 B.n727 B.n726 33.8737
R1453 B.n731 B.n451 33.8737
R1454 B.n796 B.t0 25.5238
R1455 B.n985 B.t4 25.5238
R1456 B.n826 B.t3 24.4141
R1457 B.n1003 B.t5 24.4141
R1458 B.n857 B.t1 23.3044
R1459 B.n1025 B.t2 23.3044
R1460 B B.n1037 18.0485
R1461 B.n850 B.t1 14.4267
R1462 B.n18 B.t2 14.4267
R1463 B.n394 B.t3 13.317
R1464 B.t5 B.n1002 13.317
R1465 B.n789 B.t0 12.2073
R1466 B.n53 B.t4 12.2073
R1467 B.n148 B.n87 10.6151
R1468 B.n151 B.n148 10.6151
R1469 B.n152 B.n151 10.6151
R1470 B.n155 B.n152 10.6151
R1471 B.n156 B.n155 10.6151
R1472 B.n159 B.n156 10.6151
R1473 B.n160 B.n159 10.6151
R1474 B.n163 B.n160 10.6151
R1475 B.n164 B.n163 10.6151
R1476 B.n167 B.n164 10.6151
R1477 B.n168 B.n167 10.6151
R1478 B.n171 B.n168 10.6151
R1479 B.n172 B.n171 10.6151
R1480 B.n175 B.n172 10.6151
R1481 B.n176 B.n175 10.6151
R1482 B.n179 B.n176 10.6151
R1483 B.n180 B.n179 10.6151
R1484 B.n183 B.n180 10.6151
R1485 B.n184 B.n183 10.6151
R1486 B.n187 B.n184 10.6151
R1487 B.n188 B.n187 10.6151
R1488 B.n191 B.n188 10.6151
R1489 B.n192 B.n191 10.6151
R1490 B.n195 B.n192 10.6151
R1491 B.n196 B.n195 10.6151
R1492 B.n199 B.n196 10.6151
R1493 B.n200 B.n199 10.6151
R1494 B.n203 B.n200 10.6151
R1495 B.n204 B.n203 10.6151
R1496 B.n207 B.n204 10.6151
R1497 B.n208 B.n207 10.6151
R1498 B.n211 B.n208 10.6151
R1499 B.n212 B.n211 10.6151
R1500 B.n215 B.n212 10.6151
R1501 B.n216 B.n215 10.6151
R1502 B.n219 B.n216 10.6151
R1503 B.n220 B.n219 10.6151
R1504 B.n223 B.n220 10.6151
R1505 B.n224 B.n223 10.6151
R1506 B.n227 B.n224 10.6151
R1507 B.n228 B.n227 10.6151
R1508 B.n231 B.n228 10.6151
R1509 B.n232 B.n231 10.6151
R1510 B.n235 B.n232 10.6151
R1511 B.n236 B.n235 10.6151
R1512 B.n239 B.n236 10.6151
R1513 B.n240 B.n239 10.6151
R1514 B.n243 B.n240 10.6151
R1515 B.n248 B.n245 10.6151
R1516 B.n249 B.n248 10.6151
R1517 B.n252 B.n249 10.6151
R1518 B.n253 B.n252 10.6151
R1519 B.n256 B.n253 10.6151
R1520 B.n257 B.n256 10.6151
R1521 B.n260 B.n257 10.6151
R1522 B.n261 B.n260 10.6151
R1523 B.n264 B.n261 10.6151
R1524 B.n269 B.n266 10.6151
R1525 B.n270 B.n269 10.6151
R1526 B.n273 B.n270 10.6151
R1527 B.n274 B.n273 10.6151
R1528 B.n277 B.n274 10.6151
R1529 B.n278 B.n277 10.6151
R1530 B.n281 B.n278 10.6151
R1531 B.n282 B.n281 10.6151
R1532 B.n285 B.n282 10.6151
R1533 B.n286 B.n285 10.6151
R1534 B.n289 B.n286 10.6151
R1535 B.n290 B.n289 10.6151
R1536 B.n293 B.n290 10.6151
R1537 B.n294 B.n293 10.6151
R1538 B.n297 B.n294 10.6151
R1539 B.n298 B.n297 10.6151
R1540 B.n301 B.n298 10.6151
R1541 B.n302 B.n301 10.6151
R1542 B.n305 B.n302 10.6151
R1543 B.n306 B.n305 10.6151
R1544 B.n309 B.n306 10.6151
R1545 B.n310 B.n309 10.6151
R1546 B.n313 B.n310 10.6151
R1547 B.n314 B.n313 10.6151
R1548 B.n317 B.n314 10.6151
R1549 B.n318 B.n317 10.6151
R1550 B.n321 B.n318 10.6151
R1551 B.n322 B.n321 10.6151
R1552 B.n325 B.n322 10.6151
R1553 B.n326 B.n325 10.6151
R1554 B.n329 B.n326 10.6151
R1555 B.n330 B.n329 10.6151
R1556 B.n333 B.n330 10.6151
R1557 B.n334 B.n333 10.6151
R1558 B.n337 B.n334 10.6151
R1559 B.n338 B.n337 10.6151
R1560 B.n341 B.n338 10.6151
R1561 B.n342 B.n341 10.6151
R1562 B.n345 B.n342 10.6151
R1563 B.n346 B.n345 10.6151
R1564 B.n349 B.n346 10.6151
R1565 B.n350 B.n349 10.6151
R1566 B.n353 B.n350 10.6151
R1567 B.n354 B.n353 10.6151
R1568 B.n357 B.n354 10.6151
R1569 B.n359 B.n357 10.6151
R1570 B.n360 B.n359 10.6151
R1571 B.n935 B.n360 10.6151
R1572 B.n727 B.n447 10.6151
R1573 B.n737 B.n447 10.6151
R1574 B.n738 B.n737 10.6151
R1575 B.n739 B.n738 10.6151
R1576 B.n739 B.n439 10.6151
R1577 B.n749 B.n439 10.6151
R1578 B.n750 B.n749 10.6151
R1579 B.n751 B.n750 10.6151
R1580 B.n751 B.n431 10.6151
R1581 B.n761 B.n431 10.6151
R1582 B.n762 B.n761 10.6151
R1583 B.n763 B.n762 10.6151
R1584 B.n763 B.n423 10.6151
R1585 B.n773 B.n423 10.6151
R1586 B.n774 B.n773 10.6151
R1587 B.n775 B.n774 10.6151
R1588 B.n775 B.n415 10.6151
R1589 B.n785 B.n415 10.6151
R1590 B.n786 B.n785 10.6151
R1591 B.n787 B.n786 10.6151
R1592 B.n787 B.n408 10.6151
R1593 B.n798 B.n408 10.6151
R1594 B.n799 B.n798 10.6151
R1595 B.n800 B.n799 10.6151
R1596 B.n800 B.n400 10.6151
R1597 B.n810 B.n400 10.6151
R1598 B.n811 B.n810 10.6151
R1599 B.n812 B.n811 10.6151
R1600 B.n812 B.n391 10.6151
R1601 B.n822 B.n391 10.6151
R1602 B.n823 B.n822 10.6151
R1603 B.n824 B.n823 10.6151
R1604 B.n824 B.n384 10.6151
R1605 B.n834 B.n384 10.6151
R1606 B.n835 B.n834 10.6151
R1607 B.n836 B.n835 10.6151
R1608 B.n836 B.n376 10.6151
R1609 B.n846 B.n376 10.6151
R1610 B.n847 B.n846 10.6151
R1611 B.n848 B.n847 10.6151
R1612 B.n848 B.n369 10.6151
R1613 B.n859 B.n369 10.6151
R1614 B.n860 B.n859 10.6151
R1615 B.n862 B.n860 10.6151
R1616 B.n862 B.n861 10.6151
R1617 B.n861 B.n361 10.6151
R1618 B.n873 B.n361 10.6151
R1619 B.n874 B.n873 10.6151
R1620 B.n875 B.n874 10.6151
R1621 B.n876 B.n875 10.6151
R1622 B.n878 B.n876 10.6151
R1623 B.n879 B.n878 10.6151
R1624 B.n880 B.n879 10.6151
R1625 B.n881 B.n880 10.6151
R1626 B.n883 B.n881 10.6151
R1627 B.n884 B.n883 10.6151
R1628 B.n885 B.n884 10.6151
R1629 B.n886 B.n885 10.6151
R1630 B.n888 B.n886 10.6151
R1631 B.n889 B.n888 10.6151
R1632 B.n890 B.n889 10.6151
R1633 B.n891 B.n890 10.6151
R1634 B.n893 B.n891 10.6151
R1635 B.n894 B.n893 10.6151
R1636 B.n895 B.n894 10.6151
R1637 B.n896 B.n895 10.6151
R1638 B.n898 B.n896 10.6151
R1639 B.n899 B.n898 10.6151
R1640 B.n900 B.n899 10.6151
R1641 B.n901 B.n900 10.6151
R1642 B.n903 B.n901 10.6151
R1643 B.n904 B.n903 10.6151
R1644 B.n905 B.n904 10.6151
R1645 B.n906 B.n905 10.6151
R1646 B.n908 B.n906 10.6151
R1647 B.n909 B.n908 10.6151
R1648 B.n910 B.n909 10.6151
R1649 B.n911 B.n910 10.6151
R1650 B.n913 B.n911 10.6151
R1651 B.n914 B.n913 10.6151
R1652 B.n915 B.n914 10.6151
R1653 B.n916 B.n915 10.6151
R1654 B.n918 B.n916 10.6151
R1655 B.n919 B.n918 10.6151
R1656 B.n920 B.n919 10.6151
R1657 B.n921 B.n920 10.6151
R1658 B.n923 B.n921 10.6151
R1659 B.n924 B.n923 10.6151
R1660 B.n925 B.n924 10.6151
R1661 B.n926 B.n925 10.6151
R1662 B.n928 B.n926 10.6151
R1663 B.n929 B.n928 10.6151
R1664 B.n930 B.n929 10.6151
R1665 B.n931 B.n930 10.6151
R1666 B.n933 B.n931 10.6151
R1667 B.n934 B.n933 10.6151
R1668 B.n515 B.n451 10.6151
R1669 B.n516 B.n515 10.6151
R1670 B.n517 B.n516 10.6151
R1671 B.n517 B.n511 10.6151
R1672 B.n523 B.n511 10.6151
R1673 B.n524 B.n523 10.6151
R1674 B.n525 B.n524 10.6151
R1675 B.n525 B.n509 10.6151
R1676 B.n531 B.n509 10.6151
R1677 B.n532 B.n531 10.6151
R1678 B.n533 B.n532 10.6151
R1679 B.n533 B.n507 10.6151
R1680 B.n539 B.n507 10.6151
R1681 B.n540 B.n539 10.6151
R1682 B.n541 B.n540 10.6151
R1683 B.n541 B.n505 10.6151
R1684 B.n547 B.n505 10.6151
R1685 B.n548 B.n547 10.6151
R1686 B.n549 B.n548 10.6151
R1687 B.n549 B.n503 10.6151
R1688 B.n555 B.n503 10.6151
R1689 B.n556 B.n555 10.6151
R1690 B.n557 B.n556 10.6151
R1691 B.n557 B.n501 10.6151
R1692 B.n563 B.n501 10.6151
R1693 B.n564 B.n563 10.6151
R1694 B.n565 B.n564 10.6151
R1695 B.n565 B.n499 10.6151
R1696 B.n571 B.n499 10.6151
R1697 B.n572 B.n571 10.6151
R1698 B.n573 B.n572 10.6151
R1699 B.n573 B.n497 10.6151
R1700 B.n579 B.n497 10.6151
R1701 B.n580 B.n579 10.6151
R1702 B.n581 B.n580 10.6151
R1703 B.n581 B.n495 10.6151
R1704 B.n587 B.n495 10.6151
R1705 B.n588 B.n587 10.6151
R1706 B.n589 B.n588 10.6151
R1707 B.n589 B.n493 10.6151
R1708 B.n595 B.n493 10.6151
R1709 B.n596 B.n595 10.6151
R1710 B.n597 B.n596 10.6151
R1711 B.n597 B.n491 10.6151
R1712 B.n603 B.n491 10.6151
R1713 B.n604 B.n603 10.6151
R1714 B.n605 B.n604 10.6151
R1715 B.n605 B.n489 10.6151
R1716 B.n612 B.n611 10.6151
R1717 B.n613 B.n612 10.6151
R1718 B.n613 B.n484 10.6151
R1719 B.n619 B.n484 10.6151
R1720 B.n620 B.n619 10.6151
R1721 B.n621 B.n620 10.6151
R1722 B.n621 B.n482 10.6151
R1723 B.n627 B.n482 10.6151
R1724 B.n628 B.n627 10.6151
R1725 B.n630 B.n478 10.6151
R1726 B.n636 B.n478 10.6151
R1727 B.n637 B.n636 10.6151
R1728 B.n638 B.n637 10.6151
R1729 B.n638 B.n476 10.6151
R1730 B.n644 B.n476 10.6151
R1731 B.n645 B.n644 10.6151
R1732 B.n646 B.n645 10.6151
R1733 B.n646 B.n474 10.6151
R1734 B.n652 B.n474 10.6151
R1735 B.n653 B.n652 10.6151
R1736 B.n654 B.n653 10.6151
R1737 B.n654 B.n472 10.6151
R1738 B.n660 B.n472 10.6151
R1739 B.n661 B.n660 10.6151
R1740 B.n662 B.n661 10.6151
R1741 B.n662 B.n470 10.6151
R1742 B.n668 B.n470 10.6151
R1743 B.n669 B.n668 10.6151
R1744 B.n670 B.n669 10.6151
R1745 B.n670 B.n468 10.6151
R1746 B.n676 B.n468 10.6151
R1747 B.n677 B.n676 10.6151
R1748 B.n678 B.n677 10.6151
R1749 B.n678 B.n466 10.6151
R1750 B.n684 B.n466 10.6151
R1751 B.n685 B.n684 10.6151
R1752 B.n686 B.n685 10.6151
R1753 B.n686 B.n464 10.6151
R1754 B.n692 B.n464 10.6151
R1755 B.n693 B.n692 10.6151
R1756 B.n694 B.n693 10.6151
R1757 B.n694 B.n462 10.6151
R1758 B.n700 B.n462 10.6151
R1759 B.n701 B.n700 10.6151
R1760 B.n702 B.n701 10.6151
R1761 B.n702 B.n460 10.6151
R1762 B.n708 B.n460 10.6151
R1763 B.n709 B.n708 10.6151
R1764 B.n710 B.n709 10.6151
R1765 B.n710 B.n458 10.6151
R1766 B.n716 B.n458 10.6151
R1767 B.n717 B.n716 10.6151
R1768 B.n718 B.n717 10.6151
R1769 B.n718 B.n456 10.6151
R1770 B.n456 B.n455 10.6151
R1771 B.n725 B.n455 10.6151
R1772 B.n726 B.n725 10.6151
R1773 B.n732 B.n731 10.6151
R1774 B.n733 B.n732 10.6151
R1775 B.n733 B.n443 10.6151
R1776 B.n743 B.n443 10.6151
R1777 B.n744 B.n743 10.6151
R1778 B.n745 B.n744 10.6151
R1779 B.n745 B.n435 10.6151
R1780 B.n755 B.n435 10.6151
R1781 B.n756 B.n755 10.6151
R1782 B.n757 B.n756 10.6151
R1783 B.n757 B.n427 10.6151
R1784 B.n767 B.n427 10.6151
R1785 B.n768 B.n767 10.6151
R1786 B.n769 B.n768 10.6151
R1787 B.n769 B.n419 10.6151
R1788 B.n779 B.n419 10.6151
R1789 B.n780 B.n779 10.6151
R1790 B.n781 B.n780 10.6151
R1791 B.n781 B.n411 10.6151
R1792 B.n792 B.n411 10.6151
R1793 B.n793 B.n792 10.6151
R1794 B.n794 B.n793 10.6151
R1795 B.n794 B.n404 10.6151
R1796 B.n804 B.n404 10.6151
R1797 B.n805 B.n804 10.6151
R1798 B.n806 B.n805 10.6151
R1799 B.n806 B.n396 10.6151
R1800 B.n816 B.n396 10.6151
R1801 B.n817 B.n816 10.6151
R1802 B.n818 B.n817 10.6151
R1803 B.n818 B.n388 10.6151
R1804 B.n828 B.n388 10.6151
R1805 B.n829 B.n828 10.6151
R1806 B.n830 B.n829 10.6151
R1807 B.n830 B.n380 10.6151
R1808 B.n840 B.n380 10.6151
R1809 B.n841 B.n840 10.6151
R1810 B.n842 B.n841 10.6151
R1811 B.n842 B.n372 10.6151
R1812 B.n853 B.n372 10.6151
R1813 B.n854 B.n853 10.6151
R1814 B.n855 B.n854 10.6151
R1815 B.n855 B.n365 10.6151
R1816 B.n866 B.n365 10.6151
R1817 B.n867 B.n866 10.6151
R1818 B.n868 B.n867 10.6151
R1819 B.n868 B.n0 10.6151
R1820 B.n1031 B.n1 10.6151
R1821 B.n1031 B.n1030 10.6151
R1822 B.n1030 B.n1029 10.6151
R1823 B.n1029 B.n10 10.6151
R1824 B.n1023 B.n10 10.6151
R1825 B.n1023 B.n1022 10.6151
R1826 B.n1022 B.n1021 10.6151
R1827 B.n1021 B.n16 10.6151
R1828 B.n1015 B.n16 10.6151
R1829 B.n1015 B.n1014 10.6151
R1830 B.n1014 B.n1013 10.6151
R1831 B.n1013 B.n24 10.6151
R1832 B.n1007 B.n24 10.6151
R1833 B.n1007 B.n1006 10.6151
R1834 B.n1006 B.n1005 10.6151
R1835 B.n1005 B.n31 10.6151
R1836 B.n999 B.n31 10.6151
R1837 B.n999 B.n998 10.6151
R1838 B.n998 B.n997 10.6151
R1839 B.n997 B.n38 10.6151
R1840 B.n991 B.n38 10.6151
R1841 B.n991 B.n990 10.6151
R1842 B.n990 B.n989 10.6151
R1843 B.n989 B.n45 10.6151
R1844 B.n983 B.n45 10.6151
R1845 B.n983 B.n982 10.6151
R1846 B.n982 B.n981 10.6151
R1847 B.n981 B.n51 10.6151
R1848 B.n975 B.n51 10.6151
R1849 B.n975 B.n974 10.6151
R1850 B.n974 B.n973 10.6151
R1851 B.n973 B.n59 10.6151
R1852 B.n967 B.n59 10.6151
R1853 B.n967 B.n966 10.6151
R1854 B.n966 B.n965 10.6151
R1855 B.n965 B.n66 10.6151
R1856 B.n959 B.n66 10.6151
R1857 B.n959 B.n958 10.6151
R1858 B.n958 B.n957 10.6151
R1859 B.n957 B.n73 10.6151
R1860 B.n951 B.n73 10.6151
R1861 B.n951 B.n950 10.6151
R1862 B.n950 B.n949 10.6151
R1863 B.n949 B.n80 10.6151
R1864 B.n943 B.n80 10.6151
R1865 B.n943 B.n942 10.6151
R1866 B.n942 B.n941 10.6151
R1867 B.n244 B.n243 9.36635
R1868 B.n266 B.n265 9.36635
R1869 B.n489 B.n488 9.36635
R1870 B.n630 B.n629 9.36635
R1871 B.n753 B.t14 3.32963
R1872 B.n955 B.t7 3.32963
R1873 B.n1037 B.n0 2.81026
R1874 B.n1037 B.n1 2.81026
R1875 B.n245 B.n244 1.24928
R1876 B.n265 B.n264 1.24928
R1877 B.n611 B.n488 1.24928
R1878 B.n629 B.n628 1.24928
R1879 VN.n30 VN.n29 161.3
R1880 VN.n28 VN.n17 161.3
R1881 VN.n27 VN.n26 161.3
R1882 VN.n25 VN.n18 161.3
R1883 VN.n24 VN.n23 161.3
R1884 VN.n22 VN.n19 161.3
R1885 VN.n14 VN.n13 161.3
R1886 VN.n12 VN.n1 161.3
R1887 VN.n11 VN.n10 161.3
R1888 VN.n9 VN.n2 161.3
R1889 VN.n8 VN.n7 161.3
R1890 VN.n6 VN.n3 161.3
R1891 VN.n20 VN.t3 147.251
R1892 VN.n4 VN.t2 147.251
R1893 VN.n5 VN.t5 113.85
R1894 VN.n0 VN.t4 113.85
R1895 VN.n21 VN.t1 113.85
R1896 VN.n16 VN.t0 113.85
R1897 VN.n15 VN.n0 70.0045
R1898 VN.n31 VN.n16 70.0045
R1899 VN.n11 VN.n2 56.5193
R1900 VN.n27 VN.n18 56.5193
R1901 VN VN.n31 52.7973
R1902 VN.n5 VN.n4 49.4021
R1903 VN.n21 VN.n20 49.4021
R1904 VN.n6 VN.n5 24.4675
R1905 VN.n7 VN.n6 24.4675
R1906 VN.n7 VN.n2 24.4675
R1907 VN.n12 VN.n11 24.4675
R1908 VN.n13 VN.n12 24.4675
R1909 VN.n23 VN.n18 24.4675
R1910 VN.n23 VN.n22 24.4675
R1911 VN.n22 VN.n21 24.4675
R1912 VN.n29 VN.n28 24.4675
R1913 VN.n28 VN.n27 24.4675
R1914 VN.n13 VN.n0 20.0634
R1915 VN.n29 VN.n16 20.0634
R1916 VN.n20 VN.n19 3.91167
R1917 VN.n4 VN.n3 3.91167
R1918 VN.n31 VN.n30 0.354971
R1919 VN.n15 VN.n14 0.354971
R1920 VN VN.n15 0.26696
R1921 VN.n30 VN.n17 0.189894
R1922 VN.n26 VN.n17 0.189894
R1923 VN.n26 VN.n25 0.189894
R1924 VN.n25 VN.n24 0.189894
R1925 VN.n24 VN.n19 0.189894
R1926 VN.n8 VN.n3 0.189894
R1927 VN.n9 VN.n8 0.189894
R1928 VN.n10 VN.n9 0.189894
R1929 VN.n10 VN.n1 0.189894
R1930 VN.n14 VN.n1 0.189894
R1931 VDD2.n1 VDD2.t3 63.137
R1932 VDD2.n2 VDD2.t5 60.9879
R1933 VDD2.n1 VDD2.n0 60.3065
R1934 VDD2 VDD2.n3 60.3038
R1935 VDD2.n2 VDD2.n1 45.8123
R1936 VDD2 VDD2.n2 2.26343
R1937 VDD2.n3 VDD2.t4 1.36132
R1938 VDD2.n3 VDD2.t2 1.36132
R1939 VDD2.n0 VDD2.t0 1.36132
R1940 VDD2.n0 VDD2.t1 1.36132
C0 VDD1 VTAIL 8.72438f
C1 VDD1 VDD2 1.59504f
C2 VN VTAIL 8.47336f
C3 VP VDD1 8.65905f
C4 VN VDD2 8.314731f
C5 VP VN 7.8663f
C6 VN VDD1 0.151484f
C7 VDD2 VTAIL 8.778389f
C8 VP VTAIL 8.487639f
C9 VP VDD2 0.499282f
C10 VDD2 B 6.811173f
C11 VDD1 B 7.160471f
C12 VTAIL B 9.167163f
C13 VN B 14.50484f
C14 VP B 13.145343f
C15 VDD2.t3 B 2.8199f
C16 VDD2.t0 B 0.244357f
C17 VDD2.t1 B 0.244357f
C18 VDD2.n0 B 2.20343f
C19 VDD2.n1 B 2.79421f
C20 VDD2.t5 B 2.80645f
C21 VDD2.n2 B 2.66189f
C22 VDD2.t4 B 0.244357f
C23 VDD2.t2 B 0.244357f
C24 VDD2.n3 B 2.2034f
C25 VN.t4 B 2.49978f
C26 VN.n0 B 0.954007f
C27 VN.n1 B 0.020371f
C28 VN.n2 B 0.027185f
C29 VN.n3 B 0.231823f
C30 VN.t5 B 2.49978f
C31 VN.t2 B 2.73022f
C32 VN.n4 B 0.90268f
C33 VN.n5 B 0.947954f
C34 VN.n6 B 0.037966f
C35 VN.n7 B 0.037966f
C36 VN.n8 B 0.020371f
C37 VN.n9 B 0.020371f
C38 VN.n10 B 0.020371f
C39 VN.n11 B 0.032294f
C40 VN.n12 B 0.037966f
C41 VN.n13 B 0.034592f
C42 VN.n14 B 0.032878f
C43 VN.n15 B 0.04287f
C44 VN.t0 B 2.49978f
C45 VN.n16 B 0.954007f
C46 VN.n17 B 0.020371f
C47 VN.n18 B 0.027185f
C48 VN.n19 B 0.231823f
C49 VN.t1 B 2.49978f
C50 VN.t3 B 2.73022f
C51 VN.n20 B 0.90268f
C52 VN.n21 B 0.947954f
C53 VN.n22 B 0.037966f
C54 VN.n23 B 0.037966f
C55 VN.n24 B 0.020371f
C56 VN.n25 B 0.020371f
C57 VN.n26 B 0.020371f
C58 VN.n27 B 0.032294f
C59 VN.n28 B 0.037966f
C60 VN.n29 B 0.034592f
C61 VN.n30 B 0.032878f
C62 VN.n31 B 1.24834f
C63 VTAIL.t2 B 0.268798f
C64 VTAIL.t5 B 0.268798f
C65 VTAIL.n0 B 2.34295f
C66 VTAIL.n1 B 0.448273f
C67 VTAIL.t6 B 2.98981f
C68 VTAIL.n2 B 0.696197f
C69 VTAIL.t10 B 0.268798f
C70 VTAIL.t11 B 0.268798f
C71 VTAIL.n3 B 2.34295f
C72 VTAIL.n4 B 2.16917f
C73 VTAIL.t0 B 0.268798f
C74 VTAIL.t3 B 0.268798f
C75 VTAIL.n5 B 2.34295f
C76 VTAIL.n6 B 2.16917f
C77 VTAIL.t1 B 2.98981f
C78 VTAIL.n7 B 0.69619f
C79 VTAIL.t8 B 0.268798f
C80 VTAIL.t9 B 0.268798f
C81 VTAIL.n8 B 2.34295f
C82 VTAIL.n9 B 0.609973f
C83 VTAIL.t7 B 2.98982f
C84 VTAIL.n10 B 2.03394f
C85 VTAIL.t4 B 2.98981f
C86 VTAIL.n11 B 1.97421f
C87 VDD1.t0 B 2.85723f
C88 VDD1.t4 B 2.85626f
C89 VDD1.t2 B 0.247507f
C90 VDD1.t3 B 0.247507f
C91 VDD1.n0 B 2.23185f
C92 VDD1.n1 B 2.94975f
C93 VDD1.t1 B 0.247507f
C94 VDD1.t5 B 0.247507f
C95 VDD1.n2 B 2.22685f
C96 VDD1.n3 B 2.69086f
C97 VP.t5 B 2.54321f
C98 VP.n0 B 0.970581f
C99 VP.n1 B 0.020725f
C100 VP.n2 B 0.027658f
C101 VP.n3 B 0.020725f
C102 VP.t0 B 2.54321f
C103 VP.n4 B 0.038626f
C104 VP.n5 B 0.020725f
C105 VP.n6 B 0.038626f
C106 VP.t4 B 2.54321f
C107 VP.n7 B 0.970581f
C108 VP.n8 B 0.020725f
C109 VP.n9 B 0.027658f
C110 VP.n10 B 0.235851f
C111 VP.t2 B 2.54321f
C112 VP.t3 B 2.77766f
C113 VP.n11 B 0.918364f
C114 VP.n12 B 0.964423f
C115 VP.n13 B 0.038626f
C116 VP.n14 B 0.038626f
C117 VP.n15 B 0.020725f
C118 VP.n16 B 0.020725f
C119 VP.n17 B 0.020725f
C120 VP.n18 B 0.032855f
C121 VP.n19 B 0.038626f
C122 VP.n20 B 0.035193f
C123 VP.n21 B 0.03345f
C124 VP.n22 B 1.2617f
C125 VP.n23 B 1.27585f
C126 VP.t1 B 2.54321f
C127 VP.n24 B 0.970581f
C128 VP.n25 B 0.035193f
C129 VP.n26 B 0.03345f
C130 VP.n27 B 0.020725f
C131 VP.n28 B 0.020725f
C132 VP.n29 B 0.032855f
C133 VP.n30 B 0.027658f
C134 VP.n31 B 0.038626f
C135 VP.n32 B 0.020725f
C136 VP.n33 B 0.020725f
C137 VP.n34 B 0.020725f
C138 VP.n35 B 0.906238f
C139 VP.n36 B 0.038626f
C140 VP.n37 B 0.038626f
C141 VP.n38 B 0.020725f
C142 VP.n39 B 0.020725f
C143 VP.n40 B 0.020725f
C144 VP.n41 B 0.032855f
C145 VP.n42 B 0.038626f
C146 VP.n43 B 0.035193f
C147 VP.n44 B 0.03345f
C148 VP.n45 B 0.043615f
.ends

