* NGSPICE file created from diff_pair_sample_1103.ext - technology: sky130A

.subckt diff_pair_sample_1103 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t9 VN.t0 VTAIL.t18 B.t0 sky130_fd_pr__nfet_01v8 ad=0.16005 pd=1.3 as=0.16005 ps=1.3 w=0.97 l=1.71
X1 VDD2.t8 VN.t1 VTAIL.t16 B.t7 sky130_fd_pr__nfet_01v8 ad=0.16005 pd=1.3 as=0.3783 ps=2.72 w=0.97 l=1.71
X2 VTAIL.t9 VP.t0 VDD1.t9 B.t9 sky130_fd_pr__nfet_01v8 ad=0.16005 pd=1.3 as=0.16005 ps=1.3 w=0.97 l=1.71
X3 VDD1.t8 VP.t1 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=0.3783 pd=2.72 as=0.16005 ps=1.3 w=0.97 l=1.71
X4 B.t23 B.t21 B.t22 B.t11 sky130_fd_pr__nfet_01v8 ad=0.3783 pd=2.72 as=0 ps=0 w=0.97 l=1.71
X5 VDD2.t7 VN.t2 VTAIL.t19 B.t6 sky130_fd_pr__nfet_01v8 ad=0.3783 pd=2.72 as=0.16005 ps=1.3 w=0.97 l=1.71
X6 VDD1.t7 VP.t2 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=0.16005 pd=1.3 as=0.16005 ps=1.3 w=0.97 l=1.71
X7 VTAIL.t13 VN.t3 VDD2.t6 B.t4 sky130_fd_pr__nfet_01v8 ad=0.16005 pd=1.3 as=0.16005 ps=1.3 w=0.97 l=1.71
X8 B.t20 B.t18 B.t19 B.t15 sky130_fd_pr__nfet_01v8 ad=0.3783 pd=2.72 as=0 ps=0 w=0.97 l=1.71
X9 VTAIL.t10 VN.t4 VDD2.t5 B.t9 sky130_fd_pr__nfet_01v8 ad=0.16005 pd=1.3 as=0.16005 ps=1.3 w=0.97 l=1.71
X10 VTAIL.t11 VN.t5 VDD2.t4 B.t1 sky130_fd_pr__nfet_01v8 ad=0.16005 pd=1.3 as=0.16005 ps=1.3 w=0.97 l=1.71
X11 VDD2.t3 VN.t6 VTAIL.t14 B.t2 sky130_fd_pr__nfet_01v8 ad=0.3783 pd=2.72 as=0.16005 ps=1.3 w=0.97 l=1.71
X12 VDD2.t2 VN.t7 VTAIL.t17 B.t3 sky130_fd_pr__nfet_01v8 ad=0.16005 pd=1.3 as=0.16005 ps=1.3 w=0.97 l=1.71
X13 VDD1.t6 VP.t3 VTAIL.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=0.16005 pd=1.3 as=0.3783 ps=2.72 w=0.97 l=1.71
X14 VDD2.t1 VN.t8 VTAIL.t15 B.t5 sky130_fd_pr__nfet_01v8 ad=0.16005 pd=1.3 as=0.3783 ps=2.72 w=0.97 l=1.71
X15 VDD1.t5 VP.t4 VTAIL.t7 B.t7 sky130_fd_pr__nfet_01v8 ad=0.16005 pd=1.3 as=0.3783 ps=2.72 w=0.97 l=1.71
X16 B.t17 B.t14 B.t16 B.t15 sky130_fd_pr__nfet_01v8 ad=0.3783 pd=2.72 as=0 ps=0 w=0.97 l=1.71
X17 VTAIL.t8 VP.t5 VDD1.t4 B.t8 sky130_fd_pr__nfet_01v8 ad=0.16005 pd=1.3 as=0.16005 ps=1.3 w=0.97 l=1.71
X18 VDD1.t3 VP.t6 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=0.16005 pd=1.3 as=0.16005 ps=1.3 w=0.97 l=1.71
X19 VTAIL.t1 VP.t7 VDD1.t2 B.t1 sky130_fd_pr__nfet_01v8 ad=0.16005 pd=1.3 as=0.16005 ps=1.3 w=0.97 l=1.71
X20 VTAIL.t12 VN.t9 VDD2.t0 B.t8 sky130_fd_pr__nfet_01v8 ad=0.16005 pd=1.3 as=0.16005 ps=1.3 w=0.97 l=1.71
X21 VTAIL.t4 VP.t8 VDD1.t1 B.t4 sky130_fd_pr__nfet_01v8 ad=0.16005 pd=1.3 as=0.16005 ps=1.3 w=0.97 l=1.71
X22 B.t13 B.t10 B.t12 B.t11 sky130_fd_pr__nfet_01v8 ad=0.3783 pd=2.72 as=0 ps=0 w=0.97 l=1.71
X23 VDD1.t0 VP.t9 VTAIL.t6 B.t6 sky130_fd_pr__nfet_01v8 ad=0.3783 pd=2.72 as=0.16005 ps=1.3 w=0.97 l=1.71
R0 VN.n30 VN.n29 181.852
R1 VN.n61 VN.n60 181.852
R2 VN.n59 VN.n31 161.3
R3 VN.n58 VN.n57 161.3
R4 VN.n56 VN.n32 161.3
R5 VN.n55 VN.n54 161.3
R6 VN.n52 VN.n33 161.3
R7 VN.n51 VN.n50 161.3
R8 VN.n49 VN.n34 161.3
R9 VN.n48 VN.n47 161.3
R10 VN.n46 VN.n35 161.3
R11 VN.n45 VN.n44 161.3
R12 VN.n43 VN.n36 161.3
R13 VN.n42 VN.n41 161.3
R14 VN.n40 VN.n37 161.3
R15 VN.n28 VN.n0 161.3
R16 VN.n27 VN.n26 161.3
R17 VN.n25 VN.n1 161.3
R18 VN.n24 VN.n23 161.3
R19 VN.n21 VN.n2 161.3
R20 VN.n20 VN.n19 161.3
R21 VN.n18 VN.n3 161.3
R22 VN.n17 VN.n16 161.3
R23 VN.n15 VN.n4 161.3
R24 VN.n14 VN.n13 161.3
R25 VN.n12 VN.n5 161.3
R26 VN.n11 VN.n10 161.3
R27 VN.n9 VN.n6 161.3
R28 VN.n8 VN.n7 66.2588
R29 VN.n39 VN.n38 66.2588
R30 VN.n27 VN.n1 46.321
R31 VN.n58 VN.n32 46.321
R32 VN.n7 VN.t2 43.4126
R33 VN.n38 VN.t8 43.4126
R34 VN.n10 VN.n5 42.4359
R35 VN.n20 VN.n3 42.4359
R36 VN.n41 VN.n36 42.4359
R37 VN.n51 VN.n34 42.4359
R38 VN VN.n61 40.1842
R39 VN.n14 VN.n5 38.5509
R40 VN.n16 VN.n3 38.5509
R41 VN.n45 VN.n36 38.5509
R42 VN.n47 VN.n34 38.5509
R43 VN.n23 VN.n1 34.6658
R44 VN.n54 VN.n32 34.6658
R45 VN.n10 VN.n9 24.4675
R46 VN.n15 VN.n14 24.4675
R47 VN.n16 VN.n15 24.4675
R48 VN.n21 VN.n20 24.4675
R49 VN.n28 VN.n27 24.4675
R50 VN.n41 VN.n40 24.4675
R51 VN.n47 VN.n46 24.4675
R52 VN.n46 VN.n45 24.4675
R53 VN.n52 VN.n51 24.4675
R54 VN.n59 VN.n58 24.4675
R55 VN.n23 VN.n22 22.5101
R56 VN.n54 VN.n53 22.5101
R57 VN.n38 VN.n37 18.5717
R58 VN.n7 VN.n6 18.5717
R59 VN.n15 VN.t7 13.6713
R60 VN.n8 VN.t4 13.6713
R61 VN.n22 VN.t5 13.6713
R62 VN.n29 VN.t1 13.6713
R63 VN.n46 VN.t0 13.6713
R64 VN.n39 VN.t9 13.6713
R65 VN.n53 VN.t3 13.6713
R66 VN.n60 VN.t6 13.6713
R67 VN.n29 VN.n28 3.91522
R68 VN.n60 VN.n59 3.91522
R69 VN.n9 VN.n8 1.95786
R70 VN.n22 VN.n21 1.95786
R71 VN.n40 VN.n39 1.95786
R72 VN.n53 VN.n52 1.95786
R73 VN.n61 VN.n31 0.189894
R74 VN.n57 VN.n31 0.189894
R75 VN.n57 VN.n56 0.189894
R76 VN.n56 VN.n55 0.189894
R77 VN.n55 VN.n33 0.189894
R78 VN.n50 VN.n33 0.189894
R79 VN.n50 VN.n49 0.189894
R80 VN.n49 VN.n48 0.189894
R81 VN.n48 VN.n35 0.189894
R82 VN.n44 VN.n35 0.189894
R83 VN.n44 VN.n43 0.189894
R84 VN.n43 VN.n42 0.189894
R85 VN.n42 VN.n37 0.189894
R86 VN.n11 VN.n6 0.189894
R87 VN.n12 VN.n11 0.189894
R88 VN.n13 VN.n12 0.189894
R89 VN.n13 VN.n4 0.189894
R90 VN.n17 VN.n4 0.189894
R91 VN.n18 VN.n17 0.189894
R92 VN.n19 VN.n18 0.189894
R93 VN.n19 VN.n2 0.189894
R94 VN.n24 VN.n2 0.189894
R95 VN.n25 VN.n24 0.189894
R96 VN.n26 VN.n25 0.189894
R97 VN.n26 VN.n0 0.189894
R98 VN.n30 VN.n0 0.189894
R99 VN VN.n30 0.0516364
R100 VTAIL.n16 VTAIL.t7 243.285
R101 VTAIL.n11 VTAIL.t15 243.285
R102 VTAIL.n17 VTAIL.t16 243.284
R103 VTAIL.n2 VTAIL.t5 243.284
R104 VTAIL.n15 VTAIL.n14 222.873
R105 VTAIL.n13 VTAIL.n12 222.873
R106 VTAIL.n10 VTAIL.n9 222.873
R107 VTAIL.n8 VTAIL.n7 222.873
R108 VTAIL.n19 VTAIL.n18 222.871
R109 VTAIL.n1 VTAIL.n0 222.871
R110 VTAIL.n4 VTAIL.n3 222.871
R111 VTAIL.n6 VTAIL.n5 222.871
R112 VTAIL.n18 VTAIL.t17 20.4129
R113 VTAIL.n18 VTAIL.t11 20.4129
R114 VTAIL.n0 VTAIL.t19 20.4129
R115 VTAIL.n0 VTAIL.t10 20.4129
R116 VTAIL.n3 VTAIL.t0 20.4129
R117 VTAIL.n3 VTAIL.t8 20.4129
R118 VTAIL.n5 VTAIL.t2 20.4129
R119 VTAIL.n5 VTAIL.t4 20.4129
R120 VTAIL.n14 VTAIL.t3 20.4129
R121 VTAIL.n14 VTAIL.t1 20.4129
R122 VTAIL.n12 VTAIL.t6 20.4129
R123 VTAIL.n12 VTAIL.t9 20.4129
R124 VTAIL.n9 VTAIL.t18 20.4129
R125 VTAIL.n9 VTAIL.t12 20.4129
R126 VTAIL.n7 VTAIL.t14 20.4129
R127 VTAIL.n7 VTAIL.t13 20.4129
R128 VTAIL.n8 VTAIL.n6 16.7203
R129 VTAIL.n17 VTAIL.n16 14.9617
R130 VTAIL.n10 VTAIL.n8 1.75912
R131 VTAIL.n11 VTAIL.n10 1.75912
R132 VTAIL.n15 VTAIL.n13 1.75912
R133 VTAIL.n16 VTAIL.n15 1.75912
R134 VTAIL.n6 VTAIL.n4 1.75912
R135 VTAIL.n4 VTAIL.n2 1.75912
R136 VTAIL.n19 VTAIL.n17 1.75912
R137 VTAIL VTAIL.n1 1.37766
R138 VTAIL.n13 VTAIL.n11 1.34964
R139 VTAIL.n2 VTAIL.n1 1.34964
R140 VTAIL VTAIL.n19 0.381966
R141 VDD2.n1 VDD2.t7 261.721
R142 VDD2.n4 VDD2.t3 259.964
R143 VDD2.n3 VDD2.n2 240.814
R144 VDD2 VDD2.n7 240.811
R145 VDD2.n6 VDD2.n5 239.552
R146 VDD2.n1 VDD2.n0 239.55
R147 VDD2.n4 VDD2.n3 32.9049
R148 VDD2.n7 VDD2.t0 20.4129
R149 VDD2.n7 VDD2.t1 20.4129
R150 VDD2.n5 VDD2.t6 20.4129
R151 VDD2.n5 VDD2.t9 20.4129
R152 VDD2.n2 VDD2.t4 20.4129
R153 VDD2.n2 VDD2.t8 20.4129
R154 VDD2.n0 VDD2.t5 20.4129
R155 VDD2.n0 VDD2.t2 20.4129
R156 VDD2.n6 VDD2.n4 1.75912
R157 VDD2 VDD2.n6 0.498345
R158 VDD2.n3 VDD2.n1 0.384809
R159 B.n504 B.n503 585
R160 B.n153 B.n96 585
R161 B.n152 B.n151 585
R162 B.n150 B.n149 585
R163 B.n148 B.n147 585
R164 B.n146 B.n145 585
R165 B.n144 B.n143 585
R166 B.n142 B.n141 585
R167 B.n140 B.n139 585
R168 B.n137 B.n136 585
R169 B.n135 B.n134 585
R170 B.n133 B.n132 585
R171 B.n131 B.n130 585
R172 B.n129 B.n128 585
R173 B.n127 B.n126 585
R174 B.n125 B.n124 585
R175 B.n123 B.n122 585
R176 B.n121 B.n120 585
R177 B.n119 B.n118 585
R178 B.n116 B.n115 585
R179 B.n114 B.n113 585
R180 B.n112 B.n111 585
R181 B.n110 B.n109 585
R182 B.n108 B.n107 585
R183 B.n106 B.n105 585
R184 B.n104 B.n103 585
R185 B.n102 B.n101 585
R186 B.n81 B.n80 585
R187 B.n502 B.n82 585
R188 B.n507 B.n82 585
R189 B.n501 B.n500 585
R190 B.n500 B.n78 585
R191 B.n499 B.n77 585
R192 B.n513 B.n77 585
R193 B.n498 B.n76 585
R194 B.n514 B.n76 585
R195 B.n497 B.n75 585
R196 B.n515 B.n75 585
R197 B.n496 B.n495 585
R198 B.n495 B.n71 585
R199 B.n494 B.n70 585
R200 B.n521 B.n70 585
R201 B.n493 B.n69 585
R202 B.n522 B.n69 585
R203 B.n492 B.n68 585
R204 B.n523 B.n68 585
R205 B.n491 B.n490 585
R206 B.n490 B.n64 585
R207 B.n489 B.n63 585
R208 B.n529 B.n63 585
R209 B.n488 B.n62 585
R210 B.n530 B.n62 585
R211 B.n487 B.n61 585
R212 B.n531 B.n61 585
R213 B.n486 B.n485 585
R214 B.n485 B.n57 585
R215 B.n484 B.n56 585
R216 B.n537 B.n56 585
R217 B.n483 B.n55 585
R218 B.n538 B.n55 585
R219 B.n482 B.n54 585
R220 B.n539 B.n54 585
R221 B.n481 B.n480 585
R222 B.n480 B.n50 585
R223 B.n479 B.n49 585
R224 B.n545 B.n49 585
R225 B.n478 B.n48 585
R226 B.n546 B.n48 585
R227 B.n477 B.n47 585
R228 B.n547 B.n47 585
R229 B.n476 B.n475 585
R230 B.n475 B.n46 585
R231 B.n474 B.n42 585
R232 B.n553 B.n42 585
R233 B.n473 B.n41 585
R234 B.n554 B.n41 585
R235 B.n472 B.n40 585
R236 B.n555 B.n40 585
R237 B.n471 B.n470 585
R238 B.n470 B.n36 585
R239 B.n469 B.n35 585
R240 B.n561 B.n35 585
R241 B.n468 B.n34 585
R242 B.n562 B.n34 585
R243 B.n467 B.n33 585
R244 B.n563 B.n33 585
R245 B.n466 B.n465 585
R246 B.n465 B.n29 585
R247 B.n464 B.n28 585
R248 B.n569 B.n28 585
R249 B.n463 B.n27 585
R250 B.n570 B.n27 585
R251 B.n462 B.n26 585
R252 B.n571 B.n26 585
R253 B.n461 B.n460 585
R254 B.n460 B.n25 585
R255 B.n459 B.n21 585
R256 B.n577 B.n21 585
R257 B.n458 B.n20 585
R258 B.n578 B.n20 585
R259 B.n457 B.n19 585
R260 B.n579 B.n19 585
R261 B.n456 B.n455 585
R262 B.n455 B.n15 585
R263 B.n454 B.n14 585
R264 B.n585 B.n14 585
R265 B.n453 B.n13 585
R266 B.n586 B.n13 585
R267 B.n452 B.n12 585
R268 B.n587 B.n12 585
R269 B.n451 B.n450 585
R270 B.n450 B.n8 585
R271 B.n449 B.n7 585
R272 B.n593 B.n7 585
R273 B.n448 B.n6 585
R274 B.n594 B.n6 585
R275 B.n447 B.n5 585
R276 B.n595 B.n5 585
R277 B.n446 B.n445 585
R278 B.n445 B.n4 585
R279 B.n444 B.n154 585
R280 B.n444 B.n443 585
R281 B.n434 B.n155 585
R282 B.n156 B.n155 585
R283 B.n436 B.n435 585
R284 B.n437 B.n436 585
R285 B.n433 B.n160 585
R286 B.n164 B.n160 585
R287 B.n432 B.n431 585
R288 B.n431 B.n430 585
R289 B.n162 B.n161 585
R290 B.n163 B.n162 585
R291 B.n423 B.n422 585
R292 B.n424 B.n423 585
R293 B.n421 B.n169 585
R294 B.n169 B.n168 585
R295 B.n420 B.n419 585
R296 B.n419 B.n418 585
R297 B.n171 B.n170 585
R298 B.n411 B.n171 585
R299 B.n410 B.n409 585
R300 B.n412 B.n410 585
R301 B.n408 B.n176 585
R302 B.n176 B.n175 585
R303 B.n407 B.n406 585
R304 B.n406 B.n405 585
R305 B.n178 B.n177 585
R306 B.n179 B.n178 585
R307 B.n398 B.n397 585
R308 B.n399 B.n398 585
R309 B.n396 B.n183 585
R310 B.n187 B.n183 585
R311 B.n395 B.n394 585
R312 B.n394 B.n393 585
R313 B.n185 B.n184 585
R314 B.n186 B.n185 585
R315 B.n386 B.n385 585
R316 B.n387 B.n386 585
R317 B.n384 B.n192 585
R318 B.n192 B.n191 585
R319 B.n383 B.n382 585
R320 B.n382 B.n381 585
R321 B.n194 B.n193 585
R322 B.n374 B.n194 585
R323 B.n373 B.n372 585
R324 B.n375 B.n373 585
R325 B.n371 B.n199 585
R326 B.n199 B.n198 585
R327 B.n370 B.n369 585
R328 B.n369 B.n368 585
R329 B.n201 B.n200 585
R330 B.n202 B.n201 585
R331 B.n361 B.n360 585
R332 B.n362 B.n361 585
R333 B.n359 B.n206 585
R334 B.n210 B.n206 585
R335 B.n358 B.n357 585
R336 B.n357 B.n356 585
R337 B.n208 B.n207 585
R338 B.n209 B.n208 585
R339 B.n349 B.n348 585
R340 B.n350 B.n349 585
R341 B.n347 B.n215 585
R342 B.n215 B.n214 585
R343 B.n346 B.n345 585
R344 B.n345 B.n344 585
R345 B.n217 B.n216 585
R346 B.n218 B.n217 585
R347 B.n337 B.n336 585
R348 B.n338 B.n337 585
R349 B.n335 B.n223 585
R350 B.n223 B.n222 585
R351 B.n334 B.n333 585
R352 B.n333 B.n332 585
R353 B.n225 B.n224 585
R354 B.n226 B.n225 585
R355 B.n325 B.n324 585
R356 B.n326 B.n325 585
R357 B.n323 B.n231 585
R358 B.n231 B.n230 585
R359 B.n322 B.n321 585
R360 B.n321 B.n320 585
R361 B.n233 B.n232 585
R362 B.n234 B.n233 585
R363 B.n313 B.n312 585
R364 B.n314 B.n313 585
R365 B.n237 B.n236 585
R366 B.n260 B.n259 585
R367 B.n261 B.n257 585
R368 B.n257 B.n238 585
R369 B.n263 B.n262 585
R370 B.n265 B.n256 585
R371 B.n268 B.n267 585
R372 B.n269 B.n255 585
R373 B.n271 B.n270 585
R374 B.n273 B.n254 585
R375 B.n276 B.n275 585
R376 B.n277 B.n250 585
R377 B.n279 B.n278 585
R378 B.n281 B.n249 585
R379 B.n284 B.n283 585
R380 B.n285 B.n248 585
R381 B.n287 B.n286 585
R382 B.n289 B.n247 585
R383 B.n292 B.n291 585
R384 B.n293 B.n244 585
R385 B.n296 B.n295 585
R386 B.n298 B.n243 585
R387 B.n301 B.n300 585
R388 B.n302 B.n242 585
R389 B.n304 B.n303 585
R390 B.n306 B.n241 585
R391 B.n307 B.n240 585
R392 B.n310 B.n309 585
R393 B.n311 B.n239 585
R394 B.n239 B.n238 585
R395 B.n316 B.n315 585
R396 B.n315 B.n314 585
R397 B.n317 B.n235 585
R398 B.n235 B.n234 585
R399 B.n319 B.n318 585
R400 B.n320 B.n319 585
R401 B.n229 B.n228 585
R402 B.n230 B.n229 585
R403 B.n328 B.n327 585
R404 B.n327 B.n326 585
R405 B.n329 B.n227 585
R406 B.n227 B.n226 585
R407 B.n331 B.n330 585
R408 B.n332 B.n331 585
R409 B.n221 B.n220 585
R410 B.n222 B.n221 585
R411 B.n340 B.n339 585
R412 B.n339 B.n338 585
R413 B.n341 B.n219 585
R414 B.n219 B.n218 585
R415 B.n343 B.n342 585
R416 B.n344 B.n343 585
R417 B.n213 B.n212 585
R418 B.n214 B.n213 585
R419 B.n352 B.n351 585
R420 B.n351 B.n350 585
R421 B.n353 B.n211 585
R422 B.n211 B.n209 585
R423 B.n355 B.n354 585
R424 B.n356 B.n355 585
R425 B.n205 B.n204 585
R426 B.n210 B.n205 585
R427 B.n364 B.n363 585
R428 B.n363 B.n362 585
R429 B.n365 B.n203 585
R430 B.n203 B.n202 585
R431 B.n367 B.n366 585
R432 B.n368 B.n367 585
R433 B.n197 B.n196 585
R434 B.n198 B.n197 585
R435 B.n377 B.n376 585
R436 B.n376 B.n375 585
R437 B.n378 B.n195 585
R438 B.n374 B.n195 585
R439 B.n380 B.n379 585
R440 B.n381 B.n380 585
R441 B.n190 B.n189 585
R442 B.n191 B.n190 585
R443 B.n389 B.n388 585
R444 B.n388 B.n387 585
R445 B.n390 B.n188 585
R446 B.n188 B.n186 585
R447 B.n392 B.n391 585
R448 B.n393 B.n392 585
R449 B.n182 B.n181 585
R450 B.n187 B.n182 585
R451 B.n401 B.n400 585
R452 B.n400 B.n399 585
R453 B.n402 B.n180 585
R454 B.n180 B.n179 585
R455 B.n404 B.n403 585
R456 B.n405 B.n404 585
R457 B.n174 B.n173 585
R458 B.n175 B.n174 585
R459 B.n414 B.n413 585
R460 B.n413 B.n412 585
R461 B.n415 B.n172 585
R462 B.n411 B.n172 585
R463 B.n417 B.n416 585
R464 B.n418 B.n417 585
R465 B.n167 B.n166 585
R466 B.n168 B.n167 585
R467 B.n426 B.n425 585
R468 B.n425 B.n424 585
R469 B.n427 B.n165 585
R470 B.n165 B.n163 585
R471 B.n429 B.n428 585
R472 B.n430 B.n429 585
R473 B.n159 B.n158 585
R474 B.n164 B.n159 585
R475 B.n439 B.n438 585
R476 B.n438 B.n437 585
R477 B.n440 B.n157 585
R478 B.n157 B.n156 585
R479 B.n442 B.n441 585
R480 B.n443 B.n442 585
R481 B.n2 B.n0 585
R482 B.n4 B.n2 585
R483 B.n3 B.n1 585
R484 B.n594 B.n3 585
R485 B.n592 B.n591 585
R486 B.n593 B.n592 585
R487 B.n590 B.n9 585
R488 B.n9 B.n8 585
R489 B.n589 B.n588 585
R490 B.n588 B.n587 585
R491 B.n11 B.n10 585
R492 B.n586 B.n11 585
R493 B.n584 B.n583 585
R494 B.n585 B.n584 585
R495 B.n582 B.n16 585
R496 B.n16 B.n15 585
R497 B.n581 B.n580 585
R498 B.n580 B.n579 585
R499 B.n18 B.n17 585
R500 B.n578 B.n18 585
R501 B.n576 B.n575 585
R502 B.n577 B.n576 585
R503 B.n574 B.n22 585
R504 B.n25 B.n22 585
R505 B.n573 B.n572 585
R506 B.n572 B.n571 585
R507 B.n24 B.n23 585
R508 B.n570 B.n24 585
R509 B.n568 B.n567 585
R510 B.n569 B.n568 585
R511 B.n566 B.n30 585
R512 B.n30 B.n29 585
R513 B.n565 B.n564 585
R514 B.n564 B.n563 585
R515 B.n32 B.n31 585
R516 B.n562 B.n32 585
R517 B.n560 B.n559 585
R518 B.n561 B.n560 585
R519 B.n558 B.n37 585
R520 B.n37 B.n36 585
R521 B.n557 B.n556 585
R522 B.n556 B.n555 585
R523 B.n39 B.n38 585
R524 B.n554 B.n39 585
R525 B.n552 B.n551 585
R526 B.n553 B.n552 585
R527 B.n550 B.n43 585
R528 B.n46 B.n43 585
R529 B.n549 B.n548 585
R530 B.n548 B.n547 585
R531 B.n45 B.n44 585
R532 B.n546 B.n45 585
R533 B.n544 B.n543 585
R534 B.n545 B.n544 585
R535 B.n542 B.n51 585
R536 B.n51 B.n50 585
R537 B.n541 B.n540 585
R538 B.n540 B.n539 585
R539 B.n53 B.n52 585
R540 B.n538 B.n53 585
R541 B.n536 B.n535 585
R542 B.n537 B.n536 585
R543 B.n534 B.n58 585
R544 B.n58 B.n57 585
R545 B.n533 B.n532 585
R546 B.n532 B.n531 585
R547 B.n60 B.n59 585
R548 B.n530 B.n60 585
R549 B.n528 B.n527 585
R550 B.n529 B.n528 585
R551 B.n526 B.n65 585
R552 B.n65 B.n64 585
R553 B.n525 B.n524 585
R554 B.n524 B.n523 585
R555 B.n67 B.n66 585
R556 B.n522 B.n67 585
R557 B.n520 B.n519 585
R558 B.n521 B.n520 585
R559 B.n518 B.n72 585
R560 B.n72 B.n71 585
R561 B.n517 B.n516 585
R562 B.n516 B.n515 585
R563 B.n74 B.n73 585
R564 B.n514 B.n74 585
R565 B.n512 B.n511 585
R566 B.n513 B.n512 585
R567 B.n510 B.n79 585
R568 B.n79 B.n78 585
R569 B.n509 B.n508 585
R570 B.n508 B.n507 585
R571 B.n597 B.n596 585
R572 B.n596 B.n595 585
R573 B.n315 B.n237 511.721
R574 B.n508 B.n81 511.721
R575 B.n313 B.n239 511.721
R576 B.n504 B.n82 511.721
R577 B.n245 B.t13 273.486
R578 B.n251 B.t23 273.486
R579 B.n99 B.t19 273.486
R580 B.n97 B.t16 273.486
R581 B.n506 B.n505 256.663
R582 B.n506 B.n95 256.663
R583 B.n506 B.n94 256.663
R584 B.n506 B.n93 256.663
R585 B.n506 B.n92 256.663
R586 B.n506 B.n91 256.663
R587 B.n506 B.n90 256.663
R588 B.n506 B.n89 256.663
R589 B.n506 B.n88 256.663
R590 B.n506 B.n87 256.663
R591 B.n506 B.n86 256.663
R592 B.n506 B.n85 256.663
R593 B.n506 B.n84 256.663
R594 B.n506 B.n83 256.663
R595 B.n258 B.n238 256.663
R596 B.n264 B.n238 256.663
R597 B.n266 B.n238 256.663
R598 B.n272 B.n238 256.663
R599 B.n274 B.n238 256.663
R600 B.n280 B.n238 256.663
R601 B.n282 B.n238 256.663
R602 B.n288 B.n238 256.663
R603 B.n290 B.n238 256.663
R604 B.n297 B.n238 256.663
R605 B.n299 B.n238 256.663
R606 B.n305 B.n238 256.663
R607 B.n308 B.n238 256.663
R608 B.n246 B.t12 233.922
R609 B.n252 B.t22 233.922
R610 B.n100 B.t20 233.922
R611 B.n98 B.t17 233.922
R612 B.n314 B.n238 230.745
R613 B.n507 B.n506 230.745
R614 B.n245 B.t10 207.423
R615 B.n251 B.t21 207.423
R616 B.n99 B.t18 207.423
R617 B.n97 B.t14 207.423
R618 B.n315 B.n235 163.367
R619 B.n319 B.n235 163.367
R620 B.n319 B.n229 163.367
R621 B.n327 B.n229 163.367
R622 B.n327 B.n227 163.367
R623 B.n331 B.n227 163.367
R624 B.n331 B.n221 163.367
R625 B.n339 B.n221 163.367
R626 B.n339 B.n219 163.367
R627 B.n343 B.n219 163.367
R628 B.n343 B.n213 163.367
R629 B.n351 B.n213 163.367
R630 B.n351 B.n211 163.367
R631 B.n355 B.n211 163.367
R632 B.n355 B.n205 163.367
R633 B.n363 B.n205 163.367
R634 B.n363 B.n203 163.367
R635 B.n367 B.n203 163.367
R636 B.n367 B.n197 163.367
R637 B.n376 B.n197 163.367
R638 B.n376 B.n195 163.367
R639 B.n380 B.n195 163.367
R640 B.n380 B.n190 163.367
R641 B.n388 B.n190 163.367
R642 B.n388 B.n188 163.367
R643 B.n392 B.n188 163.367
R644 B.n392 B.n182 163.367
R645 B.n400 B.n182 163.367
R646 B.n400 B.n180 163.367
R647 B.n404 B.n180 163.367
R648 B.n404 B.n174 163.367
R649 B.n413 B.n174 163.367
R650 B.n413 B.n172 163.367
R651 B.n417 B.n172 163.367
R652 B.n417 B.n167 163.367
R653 B.n425 B.n167 163.367
R654 B.n425 B.n165 163.367
R655 B.n429 B.n165 163.367
R656 B.n429 B.n159 163.367
R657 B.n438 B.n159 163.367
R658 B.n438 B.n157 163.367
R659 B.n442 B.n157 163.367
R660 B.n442 B.n2 163.367
R661 B.n596 B.n2 163.367
R662 B.n596 B.n3 163.367
R663 B.n592 B.n3 163.367
R664 B.n592 B.n9 163.367
R665 B.n588 B.n9 163.367
R666 B.n588 B.n11 163.367
R667 B.n584 B.n11 163.367
R668 B.n584 B.n16 163.367
R669 B.n580 B.n16 163.367
R670 B.n580 B.n18 163.367
R671 B.n576 B.n18 163.367
R672 B.n576 B.n22 163.367
R673 B.n572 B.n22 163.367
R674 B.n572 B.n24 163.367
R675 B.n568 B.n24 163.367
R676 B.n568 B.n30 163.367
R677 B.n564 B.n30 163.367
R678 B.n564 B.n32 163.367
R679 B.n560 B.n32 163.367
R680 B.n560 B.n37 163.367
R681 B.n556 B.n37 163.367
R682 B.n556 B.n39 163.367
R683 B.n552 B.n39 163.367
R684 B.n552 B.n43 163.367
R685 B.n548 B.n43 163.367
R686 B.n548 B.n45 163.367
R687 B.n544 B.n45 163.367
R688 B.n544 B.n51 163.367
R689 B.n540 B.n51 163.367
R690 B.n540 B.n53 163.367
R691 B.n536 B.n53 163.367
R692 B.n536 B.n58 163.367
R693 B.n532 B.n58 163.367
R694 B.n532 B.n60 163.367
R695 B.n528 B.n60 163.367
R696 B.n528 B.n65 163.367
R697 B.n524 B.n65 163.367
R698 B.n524 B.n67 163.367
R699 B.n520 B.n67 163.367
R700 B.n520 B.n72 163.367
R701 B.n516 B.n72 163.367
R702 B.n516 B.n74 163.367
R703 B.n512 B.n74 163.367
R704 B.n512 B.n79 163.367
R705 B.n508 B.n79 163.367
R706 B.n259 B.n257 163.367
R707 B.n263 B.n257 163.367
R708 B.n267 B.n265 163.367
R709 B.n271 B.n255 163.367
R710 B.n275 B.n273 163.367
R711 B.n279 B.n250 163.367
R712 B.n283 B.n281 163.367
R713 B.n287 B.n248 163.367
R714 B.n291 B.n289 163.367
R715 B.n296 B.n244 163.367
R716 B.n300 B.n298 163.367
R717 B.n304 B.n242 163.367
R718 B.n307 B.n306 163.367
R719 B.n309 B.n239 163.367
R720 B.n313 B.n233 163.367
R721 B.n321 B.n233 163.367
R722 B.n321 B.n231 163.367
R723 B.n325 B.n231 163.367
R724 B.n325 B.n225 163.367
R725 B.n333 B.n225 163.367
R726 B.n333 B.n223 163.367
R727 B.n337 B.n223 163.367
R728 B.n337 B.n217 163.367
R729 B.n345 B.n217 163.367
R730 B.n345 B.n215 163.367
R731 B.n349 B.n215 163.367
R732 B.n349 B.n208 163.367
R733 B.n357 B.n208 163.367
R734 B.n357 B.n206 163.367
R735 B.n361 B.n206 163.367
R736 B.n361 B.n201 163.367
R737 B.n369 B.n201 163.367
R738 B.n369 B.n199 163.367
R739 B.n373 B.n199 163.367
R740 B.n373 B.n194 163.367
R741 B.n382 B.n194 163.367
R742 B.n382 B.n192 163.367
R743 B.n386 B.n192 163.367
R744 B.n386 B.n185 163.367
R745 B.n394 B.n185 163.367
R746 B.n394 B.n183 163.367
R747 B.n398 B.n183 163.367
R748 B.n398 B.n178 163.367
R749 B.n406 B.n178 163.367
R750 B.n406 B.n176 163.367
R751 B.n410 B.n176 163.367
R752 B.n410 B.n171 163.367
R753 B.n419 B.n171 163.367
R754 B.n419 B.n169 163.367
R755 B.n423 B.n169 163.367
R756 B.n423 B.n162 163.367
R757 B.n431 B.n162 163.367
R758 B.n431 B.n160 163.367
R759 B.n436 B.n160 163.367
R760 B.n436 B.n155 163.367
R761 B.n444 B.n155 163.367
R762 B.n445 B.n444 163.367
R763 B.n445 B.n5 163.367
R764 B.n6 B.n5 163.367
R765 B.n7 B.n6 163.367
R766 B.n450 B.n7 163.367
R767 B.n450 B.n12 163.367
R768 B.n13 B.n12 163.367
R769 B.n14 B.n13 163.367
R770 B.n455 B.n14 163.367
R771 B.n455 B.n19 163.367
R772 B.n20 B.n19 163.367
R773 B.n21 B.n20 163.367
R774 B.n460 B.n21 163.367
R775 B.n460 B.n26 163.367
R776 B.n27 B.n26 163.367
R777 B.n28 B.n27 163.367
R778 B.n465 B.n28 163.367
R779 B.n465 B.n33 163.367
R780 B.n34 B.n33 163.367
R781 B.n35 B.n34 163.367
R782 B.n470 B.n35 163.367
R783 B.n470 B.n40 163.367
R784 B.n41 B.n40 163.367
R785 B.n42 B.n41 163.367
R786 B.n475 B.n42 163.367
R787 B.n475 B.n47 163.367
R788 B.n48 B.n47 163.367
R789 B.n49 B.n48 163.367
R790 B.n480 B.n49 163.367
R791 B.n480 B.n54 163.367
R792 B.n55 B.n54 163.367
R793 B.n56 B.n55 163.367
R794 B.n485 B.n56 163.367
R795 B.n485 B.n61 163.367
R796 B.n62 B.n61 163.367
R797 B.n63 B.n62 163.367
R798 B.n490 B.n63 163.367
R799 B.n490 B.n68 163.367
R800 B.n69 B.n68 163.367
R801 B.n70 B.n69 163.367
R802 B.n495 B.n70 163.367
R803 B.n495 B.n75 163.367
R804 B.n76 B.n75 163.367
R805 B.n77 B.n76 163.367
R806 B.n500 B.n77 163.367
R807 B.n500 B.n82 163.367
R808 B.n103 B.n102 163.367
R809 B.n107 B.n106 163.367
R810 B.n111 B.n110 163.367
R811 B.n115 B.n114 163.367
R812 B.n120 B.n119 163.367
R813 B.n124 B.n123 163.367
R814 B.n128 B.n127 163.367
R815 B.n132 B.n131 163.367
R816 B.n136 B.n135 163.367
R817 B.n141 B.n140 163.367
R818 B.n145 B.n144 163.367
R819 B.n149 B.n148 163.367
R820 B.n151 B.n96 163.367
R821 B.n314 B.n234 119.776
R822 B.n320 B.n234 119.776
R823 B.n320 B.n230 119.776
R824 B.n326 B.n230 119.776
R825 B.n326 B.n226 119.776
R826 B.n332 B.n226 119.776
R827 B.n338 B.n222 119.776
R828 B.n338 B.n218 119.776
R829 B.n344 B.n218 119.776
R830 B.n344 B.n214 119.776
R831 B.n350 B.n214 119.776
R832 B.n350 B.n209 119.776
R833 B.n356 B.n209 119.776
R834 B.n356 B.n210 119.776
R835 B.n362 B.n202 119.776
R836 B.n368 B.n202 119.776
R837 B.n368 B.n198 119.776
R838 B.n375 B.n198 119.776
R839 B.n375 B.n374 119.776
R840 B.n381 B.n191 119.776
R841 B.n387 B.n191 119.776
R842 B.n387 B.n186 119.776
R843 B.n393 B.n186 119.776
R844 B.n393 B.n187 119.776
R845 B.n399 B.n179 119.776
R846 B.n405 B.n179 119.776
R847 B.n405 B.n175 119.776
R848 B.n412 B.n175 119.776
R849 B.n412 B.n411 119.776
R850 B.n418 B.n168 119.776
R851 B.n424 B.n168 119.776
R852 B.n424 B.n163 119.776
R853 B.n430 B.n163 119.776
R854 B.n430 B.n164 119.776
R855 B.n437 B.n156 119.776
R856 B.n443 B.n156 119.776
R857 B.n443 B.n4 119.776
R858 B.n595 B.n4 119.776
R859 B.n595 B.n594 119.776
R860 B.n594 B.n593 119.776
R861 B.n593 B.n8 119.776
R862 B.n587 B.n8 119.776
R863 B.n586 B.n585 119.776
R864 B.n585 B.n15 119.776
R865 B.n579 B.n15 119.776
R866 B.n579 B.n578 119.776
R867 B.n578 B.n577 119.776
R868 B.n571 B.n25 119.776
R869 B.n571 B.n570 119.776
R870 B.n570 B.n569 119.776
R871 B.n569 B.n29 119.776
R872 B.n563 B.n29 119.776
R873 B.n562 B.n561 119.776
R874 B.n561 B.n36 119.776
R875 B.n555 B.n36 119.776
R876 B.n555 B.n554 119.776
R877 B.n554 B.n553 119.776
R878 B.n547 B.n46 119.776
R879 B.n547 B.n546 119.776
R880 B.n546 B.n545 119.776
R881 B.n545 B.n50 119.776
R882 B.n539 B.n50 119.776
R883 B.n538 B.n537 119.776
R884 B.n537 B.n57 119.776
R885 B.n531 B.n57 119.776
R886 B.n531 B.n530 119.776
R887 B.n530 B.n529 119.776
R888 B.n529 B.n64 119.776
R889 B.n523 B.n64 119.776
R890 B.n523 B.n522 119.776
R891 B.n521 B.n71 119.776
R892 B.n515 B.n71 119.776
R893 B.n515 B.n514 119.776
R894 B.n514 B.n513 119.776
R895 B.n513 B.n78 119.776
R896 B.n507 B.n78 119.776
R897 B.t11 B.n222 96.878
R898 B.n522 B.t15 96.878
R899 B.n362 B.t2 72.2183
R900 B.n381 B.t4 72.2183
R901 B.n399 B.t0 72.2183
R902 B.n418 B.t8 72.2183
R903 B.n437 B.t5 72.2183
R904 B.n587 B.t6 72.2183
R905 B.n577 B.t9 72.2183
R906 B.n563 B.t3 72.2183
R907 B.n553 B.t1 72.2183
R908 B.n539 B.t7 72.2183
R909 B.n258 B.n237 71.676
R910 B.n264 B.n263 71.676
R911 B.n267 B.n266 71.676
R912 B.n272 B.n271 71.676
R913 B.n275 B.n274 71.676
R914 B.n280 B.n279 71.676
R915 B.n283 B.n282 71.676
R916 B.n288 B.n287 71.676
R917 B.n291 B.n290 71.676
R918 B.n297 B.n296 71.676
R919 B.n300 B.n299 71.676
R920 B.n305 B.n304 71.676
R921 B.n308 B.n307 71.676
R922 B.n83 B.n81 71.676
R923 B.n103 B.n84 71.676
R924 B.n107 B.n85 71.676
R925 B.n111 B.n86 71.676
R926 B.n115 B.n87 71.676
R927 B.n120 B.n88 71.676
R928 B.n124 B.n89 71.676
R929 B.n128 B.n90 71.676
R930 B.n132 B.n91 71.676
R931 B.n136 B.n92 71.676
R932 B.n141 B.n93 71.676
R933 B.n145 B.n94 71.676
R934 B.n149 B.n95 71.676
R935 B.n505 B.n96 71.676
R936 B.n505 B.n504 71.676
R937 B.n151 B.n95 71.676
R938 B.n148 B.n94 71.676
R939 B.n144 B.n93 71.676
R940 B.n140 B.n92 71.676
R941 B.n135 B.n91 71.676
R942 B.n131 B.n90 71.676
R943 B.n127 B.n89 71.676
R944 B.n123 B.n88 71.676
R945 B.n119 B.n87 71.676
R946 B.n114 B.n86 71.676
R947 B.n110 B.n85 71.676
R948 B.n106 B.n84 71.676
R949 B.n102 B.n83 71.676
R950 B.n259 B.n258 71.676
R951 B.n265 B.n264 71.676
R952 B.n266 B.n255 71.676
R953 B.n273 B.n272 71.676
R954 B.n274 B.n250 71.676
R955 B.n281 B.n280 71.676
R956 B.n282 B.n248 71.676
R957 B.n289 B.n288 71.676
R958 B.n290 B.n244 71.676
R959 B.n298 B.n297 71.676
R960 B.n299 B.n242 71.676
R961 B.n306 B.n305 71.676
R962 B.n309 B.n308 71.676
R963 B.n294 B.n246 59.5399
R964 B.n253 B.n252 59.5399
R965 B.n117 B.n100 59.5399
R966 B.n138 B.n98 59.5399
R967 B.n210 B.t2 47.5585
R968 B.n374 B.t4 47.5585
R969 B.n187 B.t0 47.5585
R970 B.n411 B.t8 47.5585
R971 B.n164 B.t5 47.5585
R972 B.t6 B.n586 47.5585
R973 B.n25 B.t9 47.5585
R974 B.t3 B.n562 47.5585
R975 B.n46 B.t1 47.5585
R976 B.t7 B.n538 47.5585
R977 B.n246 B.n245 39.5641
R978 B.n252 B.n251 39.5641
R979 B.n100 B.n99 39.5641
R980 B.n98 B.n97 39.5641
R981 B.n509 B.n80 33.2493
R982 B.n503 B.n502 33.2493
R983 B.n312 B.n311 33.2493
R984 B.n316 B.n236 33.2493
R985 B.n332 B.t11 22.8988
R986 B.t15 B.n521 22.8988
R987 B B.n597 18.0485
R988 B.n101 B.n80 10.6151
R989 B.n104 B.n101 10.6151
R990 B.n105 B.n104 10.6151
R991 B.n108 B.n105 10.6151
R992 B.n109 B.n108 10.6151
R993 B.n112 B.n109 10.6151
R994 B.n113 B.n112 10.6151
R995 B.n116 B.n113 10.6151
R996 B.n121 B.n118 10.6151
R997 B.n122 B.n121 10.6151
R998 B.n125 B.n122 10.6151
R999 B.n126 B.n125 10.6151
R1000 B.n129 B.n126 10.6151
R1001 B.n130 B.n129 10.6151
R1002 B.n133 B.n130 10.6151
R1003 B.n134 B.n133 10.6151
R1004 B.n137 B.n134 10.6151
R1005 B.n142 B.n139 10.6151
R1006 B.n143 B.n142 10.6151
R1007 B.n146 B.n143 10.6151
R1008 B.n147 B.n146 10.6151
R1009 B.n150 B.n147 10.6151
R1010 B.n152 B.n150 10.6151
R1011 B.n153 B.n152 10.6151
R1012 B.n503 B.n153 10.6151
R1013 B.n312 B.n232 10.6151
R1014 B.n322 B.n232 10.6151
R1015 B.n323 B.n322 10.6151
R1016 B.n324 B.n323 10.6151
R1017 B.n324 B.n224 10.6151
R1018 B.n334 B.n224 10.6151
R1019 B.n335 B.n334 10.6151
R1020 B.n336 B.n335 10.6151
R1021 B.n336 B.n216 10.6151
R1022 B.n346 B.n216 10.6151
R1023 B.n347 B.n346 10.6151
R1024 B.n348 B.n347 10.6151
R1025 B.n348 B.n207 10.6151
R1026 B.n358 B.n207 10.6151
R1027 B.n359 B.n358 10.6151
R1028 B.n360 B.n359 10.6151
R1029 B.n360 B.n200 10.6151
R1030 B.n370 B.n200 10.6151
R1031 B.n371 B.n370 10.6151
R1032 B.n372 B.n371 10.6151
R1033 B.n372 B.n193 10.6151
R1034 B.n383 B.n193 10.6151
R1035 B.n384 B.n383 10.6151
R1036 B.n385 B.n384 10.6151
R1037 B.n385 B.n184 10.6151
R1038 B.n395 B.n184 10.6151
R1039 B.n396 B.n395 10.6151
R1040 B.n397 B.n396 10.6151
R1041 B.n397 B.n177 10.6151
R1042 B.n407 B.n177 10.6151
R1043 B.n408 B.n407 10.6151
R1044 B.n409 B.n408 10.6151
R1045 B.n409 B.n170 10.6151
R1046 B.n420 B.n170 10.6151
R1047 B.n421 B.n420 10.6151
R1048 B.n422 B.n421 10.6151
R1049 B.n422 B.n161 10.6151
R1050 B.n432 B.n161 10.6151
R1051 B.n433 B.n432 10.6151
R1052 B.n435 B.n433 10.6151
R1053 B.n435 B.n434 10.6151
R1054 B.n434 B.n154 10.6151
R1055 B.n446 B.n154 10.6151
R1056 B.n447 B.n446 10.6151
R1057 B.n448 B.n447 10.6151
R1058 B.n449 B.n448 10.6151
R1059 B.n451 B.n449 10.6151
R1060 B.n452 B.n451 10.6151
R1061 B.n453 B.n452 10.6151
R1062 B.n454 B.n453 10.6151
R1063 B.n456 B.n454 10.6151
R1064 B.n457 B.n456 10.6151
R1065 B.n458 B.n457 10.6151
R1066 B.n459 B.n458 10.6151
R1067 B.n461 B.n459 10.6151
R1068 B.n462 B.n461 10.6151
R1069 B.n463 B.n462 10.6151
R1070 B.n464 B.n463 10.6151
R1071 B.n466 B.n464 10.6151
R1072 B.n467 B.n466 10.6151
R1073 B.n468 B.n467 10.6151
R1074 B.n469 B.n468 10.6151
R1075 B.n471 B.n469 10.6151
R1076 B.n472 B.n471 10.6151
R1077 B.n473 B.n472 10.6151
R1078 B.n474 B.n473 10.6151
R1079 B.n476 B.n474 10.6151
R1080 B.n477 B.n476 10.6151
R1081 B.n478 B.n477 10.6151
R1082 B.n479 B.n478 10.6151
R1083 B.n481 B.n479 10.6151
R1084 B.n482 B.n481 10.6151
R1085 B.n483 B.n482 10.6151
R1086 B.n484 B.n483 10.6151
R1087 B.n486 B.n484 10.6151
R1088 B.n487 B.n486 10.6151
R1089 B.n488 B.n487 10.6151
R1090 B.n489 B.n488 10.6151
R1091 B.n491 B.n489 10.6151
R1092 B.n492 B.n491 10.6151
R1093 B.n493 B.n492 10.6151
R1094 B.n494 B.n493 10.6151
R1095 B.n496 B.n494 10.6151
R1096 B.n497 B.n496 10.6151
R1097 B.n498 B.n497 10.6151
R1098 B.n499 B.n498 10.6151
R1099 B.n501 B.n499 10.6151
R1100 B.n502 B.n501 10.6151
R1101 B.n260 B.n236 10.6151
R1102 B.n261 B.n260 10.6151
R1103 B.n262 B.n261 10.6151
R1104 B.n262 B.n256 10.6151
R1105 B.n268 B.n256 10.6151
R1106 B.n269 B.n268 10.6151
R1107 B.n270 B.n269 10.6151
R1108 B.n270 B.n254 10.6151
R1109 B.n277 B.n276 10.6151
R1110 B.n278 B.n277 10.6151
R1111 B.n278 B.n249 10.6151
R1112 B.n284 B.n249 10.6151
R1113 B.n285 B.n284 10.6151
R1114 B.n286 B.n285 10.6151
R1115 B.n286 B.n247 10.6151
R1116 B.n292 B.n247 10.6151
R1117 B.n293 B.n292 10.6151
R1118 B.n295 B.n243 10.6151
R1119 B.n301 B.n243 10.6151
R1120 B.n302 B.n301 10.6151
R1121 B.n303 B.n302 10.6151
R1122 B.n303 B.n241 10.6151
R1123 B.n241 B.n240 10.6151
R1124 B.n310 B.n240 10.6151
R1125 B.n311 B.n310 10.6151
R1126 B.n317 B.n316 10.6151
R1127 B.n318 B.n317 10.6151
R1128 B.n318 B.n228 10.6151
R1129 B.n328 B.n228 10.6151
R1130 B.n329 B.n328 10.6151
R1131 B.n330 B.n329 10.6151
R1132 B.n330 B.n220 10.6151
R1133 B.n340 B.n220 10.6151
R1134 B.n341 B.n340 10.6151
R1135 B.n342 B.n341 10.6151
R1136 B.n342 B.n212 10.6151
R1137 B.n352 B.n212 10.6151
R1138 B.n353 B.n352 10.6151
R1139 B.n354 B.n353 10.6151
R1140 B.n354 B.n204 10.6151
R1141 B.n364 B.n204 10.6151
R1142 B.n365 B.n364 10.6151
R1143 B.n366 B.n365 10.6151
R1144 B.n366 B.n196 10.6151
R1145 B.n377 B.n196 10.6151
R1146 B.n378 B.n377 10.6151
R1147 B.n379 B.n378 10.6151
R1148 B.n379 B.n189 10.6151
R1149 B.n389 B.n189 10.6151
R1150 B.n390 B.n389 10.6151
R1151 B.n391 B.n390 10.6151
R1152 B.n391 B.n181 10.6151
R1153 B.n401 B.n181 10.6151
R1154 B.n402 B.n401 10.6151
R1155 B.n403 B.n402 10.6151
R1156 B.n403 B.n173 10.6151
R1157 B.n414 B.n173 10.6151
R1158 B.n415 B.n414 10.6151
R1159 B.n416 B.n415 10.6151
R1160 B.n416 B.n166 10.6151
R1161 B.n426 B.n166 10.6151
R1162 B.n427 B.n426 10.6151
R1163 B.n428 B.n427 10.6151
R1164 B.n428 B.n158 10.6151
R1165 B.n439 B.n158 10.6151
R1166 B.n440 B.n439 10.6151
R1167 B.n441 B.n440 10.6151
R1168 B.n441 B.n0 10.6151
R1169 B.n591 B.n1 10.6151
R1170 B.n591 B.n590 10.6151
R1171 B.n590 B.n589 10.6151
R1172 B.n589 B.n10 10.6151
R1173 B.n583 B.n10 10.6151
R1174 B.n583 B.n582 10.6151
R1175 B.n582 B.n581 10.6151
R1176 B.n581 B.n17 10.6151
R1177 B.n575 B.n17 10.6151
R1178 B.n575 B.n574 10.6151
R1179 B.n574 B.n573 10.6151
R1180 B.n573 B.n23 10.6151
R1181 B.n567 B.n23 10.6151
R1182 B.n567 B.n566 10.6151
R1183 B.n566 B.n565 10.6151
R1184 B.n565 B.n31 10.6151
R1185 B.n559 B.n31 10.6151
R1186 B.n559 B.n558 10.6151
R1187 B.n558 B.n557 10.6151
R1188 B.n557 B.n38 10.6151
R1189 B.n551 B.n38 10.6151
R1190 B.n551 B.n550 10.6151
R1191 B.n550 B.n549 10.6151
R1192 B.n549 B.n44 10.6151
R1193 B.n543 B.n44 10.6151
R1194 B.n543 B.n542 10.6151
R1195 B.n542 B.n541 10.6151
R1196 B.n541 B.n52 10.6151
R1197 B.n535 B.n52 10.6151
R1198 B.n535 B.n534 10.6151
R1199 B.n534 B.n533 10.6151
R1200 B.n533 B.n59 10.6151
R1201 B.n527 B.n59 10.6151
R1202 B.n527 B.n526 10.6151
R1203 B.n526 B.n525 10.6151
R1204 B.n525 B.n66 10.6151
R1205 B.n519 B.n66 10.6151
R1206 B.n519 B.n518 10.6151
R1207 B.n518 B.n517 10.6151
R1208 B.n517 B.n73 10.6151
R1209 B.n511 B.n73 10.6151
R1210 B.n511 B.n510 10.6151
R1211 B.n510 B.n509 10.6151
R1212 B.n117 B.n116 9.36635
R1213 B.n139 B.n138 9.36635
R1214 B.n254 B.n253 9.36635
R1215 B.n295 B.n294 9.36635
R1216 B.n597 B.n0 2.81026
R1217 B.n597 B.n1 2.81026
R1218 B.n118 B.n117 1.24928
R1219 B.n138 B.n137 1.24928
R1220 B.n276 B.n253 1.24928
R1221 B.n294 B.n293 1.24928
R1222 VP.n41 VP.n40 181.852
R1223 VP.n70 VP.n69 181.852
R1224 VP.n39 VP.n38 181.852
R1225 VP.n18 VP.n15 161.3
R1226 VP.n20 VP.n19 161.3
R1227 VP.n21 VP.n14 161.3
R1228 VP.n23 VP.n22 161.3
R1229 VP.n24 VP.n13 161.3
R1230 VP.n26 VP.n25 161.3
R1231 VP.n27 VP.n12 161.3
R1232 VP.n29 VP.n28 161.3
R1233 VP.n30 VP.n11 161.3
R1234 VP.n33 VP.n32 161.3
R1235 VP.n34 VP.n10 161.3
R1236 VP.n36 VP.n35 161.3
R1237 VP.n37 VP.n9 161.3
R1238 VP.n68 VP.n0 161.3
R1239 VP.n67 VP.n66 161.3
R1240 VP.n65 VP.n1 161.3
R1241 VP.n64 VP.n63 161.3
R1242 VP.n61 VP.n2 161.3
R1243 VP.n60 VP.n59 161.3
R1244 VP.n58 VP.n3 161.3
R1245 VP.n57 VP.n56 161.3
R1246 VP.n55 VP.n4 161.3
R1247 VP.n54 VP.n53 161.3
R1248 VP.n52 VP.n5 161.3
R1249 VP.n51 VP.n50 161.3
R1250 VP.n49 VP.n6 161.3
R1251 VP.n47 VP.n46 161.3
R1252 VP.n45 VP.n7 161.3
R1253 VP.n44 VP.n43 161.3
R1254 VP.n42 VP.n8 161.3
R1255 VP.n17 VP.n16 66.2588
R1256 VP.n43 VP.n7 46.321
R1257 VP.n67 VP.n1 46.321
R1258 VP.n36 VP.n10 46.321
R1259 VP.n16 VP.t9 43.4126
R1260 VP.n50 VP.n5 42.4359
R1261 VP.n60 VP.n3 42.4359
R1262 VP.n29 VP.n12 42.4359
R1263 VP.n19 VP.n14 42.4359
R1264 VP.n40 VP.n39 39.8035
R1265 VP.n54 VP.n5 38.5509
R1266 VP.n56 VP.n3 38.5509
R1267 VP.n25 VP.n12 38.5509
R1268 VP.n23 VP.n14 38.5509
R1269 VP.n47 VP.n7 34.6658
R1270 VP.n63 VP.n1 34.6658
R1271 VP.n32 VP.n10 34.6658
R1272 VP.n43 VP.n42 24.4675
R1273 VP.n50 VP.n49 24.4675
R1274 VP.n55 VP.n54 24.4675
R1275 VP.n56 VP.n55 24.4675
R1276 VP.n61 VP.n60 24.4675
R1277 VP.n68 VP.n67 24.4675
R1278 VP.n37 VP.n36 24.4675
R1279 VP.n30 VP.n29 24.4675
R1280 VP.n24 VP.n23 24.4675
R1281 VP.n25 VP.n24 24.4675
R1282 VP.n19 VP.n18 24.4675
R1283 VP.n48 VP.n47 22.5101
R1284 VP.n63 VP.n62 22.5101
R1285 VP.n32 VP.n31 22.5101
R1286 VP.n16 VP.n15 18.5717
R1287 VP.n55 VP.t6 13.6713
R1288 VP.n41 VP.t1 13.6713
R1289 VP.n48 VP.t8 13.6713
R1290 VP.n62 VP.t5 13.6713
R1291 VP.n69 VP.t3 13.6713
R1292 VP.n24 VP.t2 13.6713
R1293 VP.n38 VP.t4 13.6713
R1294 VP.n31 VP.t7 13.6713
R1295 VP.n17 VP.t0 13.6713
R1296 VP.n42 VP.n41 3.91522
R1297 VP.n69 VP.n68 3.91522
R1298 VP.n38 VP.n37 3.91522
R1299 VP.n49 VP.n48 1.95786
R1300 VP.n62 VP.n61 1.95786
R1301 VP.n31 VP.n30 1.95786
R1302 VP.n18 VP.n17 1.95786
R1303 VP.n20 VP.n15 0.189894
R1304 VP.n21 VP.n20 0.189894
R1305 VP.n22 VP.n21 0.189894
R1306 VP.n22 VP.n13 0.189894
R1307 VP.n26 VP.n13 0.189894
R1308 VP.n27 VP.n26 0.189894
R1309 VP.n28 VP.n27 0.189894
R1310 VP.n28 VP.n11 0.189894
R1311 VP.n33 VP.n11 0.189894
R1312 VP.n34 VP.n33 0.189894
R1313 VP.n35 VP.n34 0.189894
R1314 VP.n35 VP.n9 0.189894
R1315 VP.n39 VP.n9 0.189894
R1316 VP.n40 VP.n8 0.189894
R1317 VP.n44 VP.n8 0.189894
R1318 VP.n45 VP.n44 0.189894
R1319 VP.n46 VP.n45 0.189894
R1320 VP.n46 VP.n6 0.189894
R1321 VP.n51 VP.n6 0.189894
R1322 VP.n52 VP.n51 0.189894
R1323 VP.n53 VP.n52 0.189894
R1324 VP.n53 VP.n4 0.189894
R1325 VP.n57 VP.n4 0.189894
R1326 VP.n58 VP.n57 0.189894
R1327 VP.n59 VP.n58 0.189894
R1328 VP.n59 VP.n2 0.189894
R1329 VP.n64 VP.n2 0.189894
R1330 VP.n65 VP.n64 0.189894
R1331 VP.n66 VP.n65 0.189894
R1332 VP.n66 VP.n0 0.189894
R1333 VP.n70 VP.n0 0.189894
R1334 VP VP.n70 0.0516364
R1335 VDD1.n1 VDD1.t0 261.723
R1336 VDD1.n3 VDD1.t8 261.721
R1337 VDD1.n5 VDD1.n4 240.814
R1338 VDD1.n7 VDD1.n6 239.552
R1339 VDD1.n1 VDD1.n0 239.552
R1340 VDD1.n3 VDD1.n2 239.55
R1341 VDD1.n7 VDD1.n5 34.3673
R1342 VDD1.n6 VDD1.t2 20.4129
R1343 VDD1.n6 VDD1.t5 20.4129
R1344 VDD1.n0 VDD1.t9 20.4129
R1345 VDD1.n0 VDD1.t7 20.4129
R1346 VDD1.n4 VDD1.t4 20.4129
R1347 VDD1.n4 VDD1.t6 20.4129
R1348 VDD1.n2 VDD1.t1 20.4129
R1349 VDD1.n2 VDD1.t3 20.4129
R1350 VDD1 VDD1.n7 1.26128
R1351 VDD1 VDD1.n1 0.498345
R1352 VDD1.n5 VDD1.n3 0.384809
C0 VDD2 VN 1.23838f
C1 VTAIL VN 2.29018f
C2 VDD2 VDD1 1.59159f
C3 VN VP 5.05365f
C4 VDD1 VTAIL 4.30235f
C5 VDD2 VTAIL 4.34975f
C6 VDD1 VP 1.55426f
C7 VDD2 VP 0.478347f
C8 VDD1 VN 0.159001f
C9 VTAIL VP 2.30431f
C10 VDD2 B 4.05478f
C11 VDD1 B 4.122865f
C12 VTAIL B 2.770452f
C13 VN B 12.79394f
C14 VP B 11.370351f
C15 VDD1.t0 B 0.087134f
C16 VDD1.t9 B 0.01386f
C17 VDD1.t7 B 0.01386f
C18 VDD1.n0 B 0.053827f
C19 VDD1.n1 B 0.49385f
C20 VDD1.t8 B 0.087134f
C21 VDD1.t1 B 0.01386f
C22 VDD1.t3 B 0.01386f
C23 VDD1.n2 B 0.053827f
C24 VDD1.n3 B 0.488325f
C25 VDD1.t4 B 0.01386f
C26 VDD1.t6 B 0.01386f
C27 VDD1.n4 B 0.055442f
C28 VDD1.n5 B 1.33984f
C29 VDD1.t2 B 0.01386f
C30 VDD1.t5 B 0.01386f
C31 VDD1.n6 B 0.053827f
C32 VDD1.n7 B 1.37344f
C33 VP.n0 B 0.032772f
C34 VP.t3 B 0.099988f
C35 VP.n1 B 0.02804f
C36 VP.n2 B 0.032772f
C37 VP.t5 B 0.099988f
C38 VP.n3 B 0.026662f
C39 VP.n4 B 0.032772f
C40 VP.t6 B 0.099988f
C41 VP.n5 B 0.026662f
C42 VP.n6 B 0.032772f
C43 VP.t8 B 0.099988f
C44 VP.n7 B 0.02804f
C45 VP.n8 B 0.032772f
C46 VP.t1 B 0.099988f
C47 VP.n9 B 0.032772f
C48 VP.t4 B 0.099988f
C49 VP.n10 B 0.02804f
C50 VP.n11 B 0.032772f
C51 VP.t7 B 0.099988f
C52 VP.n12 B 0.026662f
C53 VP.n13 B 0.032772f
C54 VP.t2 B 0.099988f
C55 VP.n14 B 0.026662f
C56 VP.n15 B 0.20957f
C57 VP.t0 B 0.099988f
C58 VP.t9 B 0.250811f
C59 VP.n16 B 0.136151f
C60 VP.n17 B 0.138095f
C61 VP.n18 B 0.033336f
C62 VP.n19 B 0.064396f
C63 VP.n20 B 0.032772f
C64 VP.n21 B 0.032772f
C65 VP.n22 B 0.032772f
C66 VP.n23 B 0.065703f
C67 VP.n24 B 0.111858f
C68 VP.n25 B 0.065703f
C69 VP.n26 B 0.032772f
C70 VP.n27 B 0.032772f
C71 VP.n28 B 0.032772f
C72 VP.n29 B 0.064396f
C73 VP.n30 B 0.033336f
C74 VP.n31 B 0.080934f
C75 VP.n32 B 0.063809f
C76 VP.n33 B 0.032772f
C77 VP.n34 B 0.032772f
C78 VP.n35 B 0.032772f
C79 VP.n36 B 0.062498f
C80 VP.n37 B 0.035748f
C81 VP.n38 B 0.150623f
C82 VP.n39 B 1.24366f
C83 VP.n40 B 1.27326f
C84 VP.n41 B 0.150623f
C85 VP.n42 B 0.035748f
C86 VP.n43 B 0.062498f
C87 VP.n44 B 0.032772f
C88 VP.n45 B 0.032772f
C89 VP.n46 B 0.032772f
C90 VP.n47 B 0.063809f
C91 VP.n48 B 0.080934f
C92 VP.n49 B 0.033336f
C93 VP.n50 B 0.064396f
C94 VP.n51 B 0.032772f
C95 VP.n52 B 0.032772f
C96 VP.n53 B 0.032772f
C97 VP.n54 B 0.065703f
C98 VP.n55 B 0.111858f
C99 VP.n56 B 0.065703f
C100 VP.n57 B 0.032772f
C101 VP.n58 B 0.032772f
C102 VP.n59 B 0.032772f
C103 VP.n60 B 0.064396f
C104 VP.n61 B 0.033336f
C105 VP.n62 B 0.080934f
C106 VP.n63 B 0.063809f
C107 VP.n64 B 0.032772f
C108 VP.n65 B 0.032772f
C109 VP.n66 B 0.032772f
C110 VP.n67 B 0.062498f
C111 VP.n68 B 0.035748f
C112 VP.n69 B 0.150623f
C113 VP.n70 B 0.034276f
C114 VDD2.t7 B 0.088508f
C115 VDD2.t5 B 0.014079f
C116 VDD2.t2 B 0.014079f
C117 VDD2.n0 B 0.054676f
C118 VDD2.n1 B 0.496029f
C119 VDD2.t4 B 0.014079f
C120 VDD2.t8 B 0.014079f
C121 VDD2.n2 B 0.056317f
C122 VDD2.n3 B 1.29273f
C123 VDD2.t3 B 0.086871f
C124 VDD2.n4 B 1.32711f
C125 VDD2.t6 B 0.014079f
C126 VDD2.t9 B 0.014079f
C127 VDD2.n5 B 0.054676f
C128 VDD2.n6 B 0.259571f
C129 VDD2.t0 B 0.014079f
C130 VDD2.t1 B 0.014079f
C131 VDD2.n7 B 0.05631f
C132 VTAIL.t19 B 0.030704f
C133 VTAIL.t10 B 0.030704f
C134 VTAIL.n0 B 0.099241f
C135 VTAIL.n1 B 0.592265f
C136 VTAIL.t5 B 0.170201f
C137 VTAIL.n2 B 0.654276f
C138 VTAIL.t0 B 0.030704f
C139 VTAIL.t8 B 0.030704f
C140 VTAIL.n3 B 0.099241f
C141 VTAIL.n4 B 0.694351f
C142 VTAIL.t2 B 0.030704f
C143 VTAIL.t4 B 0.030704f
C144 VTAIL.n5 B 0.099241f
C145 VTAIL.n6 B 1.57337f
C146 VTAIL.t14 B 0.030704f
C147 VTAIL.t13 B 0.030704f
C148 VTAIL.n7 B 0.099241f
C149 VTAIL.n8 B 1.57337f
C150 VTAIL.t18 B 0.030704f
C151 VTAIL.t12 B 0.030704f
C152 VTAIL.n9 B 0.099241f
C153 VTAIL.n10 B 0.694351f
C154 VTAIL.t15 B 0.170202f
C155 VTAIL.n11 B 0.654276f
C156 VTAIL.t6 B 0.030704f
C157 VTAIL.t9 B 0.030704f
C158 VTAIL.n12 B 0.099241f
C159 VTAIL.n13 B 0.641499f
C160 VTAIL.t3 B 0.030704f
C161 VTAIL.t1 B 0.030704f
C162 VTAIL.n14 B 0.099241f
C163 VTAIL.n15 B 0.694351f
C164 VTAIL.t7 B 0.170202f
C165 VTAIL.n16 B 1.35916f
C166 VTAIL.t16 B 0.170201f
C167 VTAIL.n17 B 1.35916f
C168 VTAIL.t17 B 0.030704f
C169 VTAIL.t11 B 0.030704f
C170 VTAIL.n18 B 0.099241f
C171 VTAIL.n19 B 0.516604f
C172 VN.n0 B 0.032569f
C173 VN.t1 B 0.099369f
C174 VN.n1 B 0.027867f
C175 VN.n2 B 0.032569f
C176 VN.t5 B 0.099369f
C177 VN.n3 B 0.026497f
C178 VN.n4 B 0.032569f
C179 VN.t7 B 0.099369f
C180 VN.n5 B 0.026497f
C181 VN.n6 B 0.208274f
C182 VN.t4 B 0.099369f
C183 VN.t2 B 0.249259f
C184 VN.n7 B 0.135308f
C185 VN.n8 B 0.13724f
C186 VN.n9 B 0.03313f
C187 VN.n10 B 0.063997f
C188 VN.n11 B 0.032569f
C189 VN.n12 B 0.032569f
C190 VN.n13 B 0.032569f
C191 VN.n14 B 0.065296f
C192 VN.n15 B 0.111166f
C193 VN.n16 B 0.065296f
C194 VN.n17 B 0.032569f
C195 VN.n18 B 0.032569f
C196 VN.n19 B 0.032569f
C197 VN.n20 B 0.063997f
C198 VN.n21 B 0.03313f
C199 VN.n22 B 0.080433f
C200 VN.n23 B 0.063414f
C201 VN.n24 B 0.032569f
C202 VN.n25 B 0.032569f
C203 VN.n26 B 0.032569f
C204 VN.n27 B 0.062112f
C205 VN.n28 B 0.035527f
C206 VN.n29 B 0.149691f
C207 VN.n30 B 0.034064f
C208 VN.n31 B 0.032569f
C209 VN.t6 B 0.099369f
C210 VN.n32 B 0.027867f
C211 VN.n33 B 0.032569f
C212 VN.t3 B 0.099369f
C213 VN.n34 B 0.026497f
C214 VN.n35 B 0.032569f
C215 VN.t0 B 0.099369f
C216 VN.n36 B 0.026497f
C217 VN.n37 B 0.208274f
C218 VN.t9 B 0.099369f
C219 VN.t8 B 0.249259f
C220 VN.n38 B 0.135308f
C221 VN.n39 B 0.13724f
C222 VN.n40 B 0.03313f
C223 VN.n41 B 0.063997f
C224 VN.n42 B 0.032569f
C225 VN.n43 B 0.032569f
C226 VN.n44 B 0.032569f
C227 VN.n45 B 0.065296f
C228 VN.n46 B 0.111166f
C229 VN.n47 B 0.065296f
C230 VN.n48 B 0.032569f
C231 VN.n49 B 0.032569f
C232 VN.n50 B 0.032569f
C233 VN.n51 B 0.063997f
C234 VN.n52 B 0.03313f
C235 VN.n53 B 0.080433f
C236 VN.n54 B 0.063414f
C237 VN.n55 B 0.032569f
C238 VN.n56 B 0.032569f
C239 VN.n57 B 0.032569f
C240 VN.n58 B 0.062112f
C241 VN.n59 B 0.035527f
C242 VN.n60 B 0.149691f
C243 VN.n61 B 1.25742f
.ends

