* NGSPICE file created from diff_pair_sample_1637.ext - technology: sky130A

.subckt diff_pair_sample_1637 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t1 VP.t0 VTAIL.t3 w_n1778_n3210# sky130_fd_pr__pfet_01v8 ad=4.3719 pd=23.2 as=4.3719 ps=23.2 w=11.21 l=1.69
X1 B.t11 B.t9 B.t10 w_n1778_n3210# sky130_fd_pr__pfet_01v8 ad=4.3719 pd=23.2 as=0 ps=0 w=11.21 l=1.69
X2 VDD2.t1 VN.t0 VTAIL.t0 w_n1778_n3210# sky130_fd_pr__pfet_01v8 ad=4.3719 pd=23.2 as=4.3719 ps=23.2 w=11.21 l=1.69
X3 VDD2.t0 VN.t1 VTAIL.t1 w_n1778_n3210# sky130_fd_pr__pfet_01v8 ad=4.3719 pd=23.2 as=4.3719 ps=23.2 w=11.21 l=1.69
X4 B.t8 B.t6 B.t7 w_n1778_n3210# sky130_fd_pr__pfet_01v8 ad=4.3719 pd=23.2 as=0 ps=0 w=11.21 l=1.69
X5 VDD1.t0 VP.t1 VTAIL.t2 w_n1778_n3210# sky130_fd_pr__pfet_01v8 ad=4.3719 pd=23.2 as=4.3719 ps=23.2 w=11.21 l=1.69
X6 B.t5 B.t3 B.t4 w_n1778_n3210# sky130_fd_pr__pfet_01v8 ad=4.3719 pd=23.2 as=0 ps=0 w=11.21 l=1.69
X7 B.t2 B.t0 B.t1 w_n1778_n3210# sky130_fd_pr__pfet_01v8 ad=4.3719 pd=23.2 as=0 ps=0 w=11.21 l=1.69
R0 VP.n0 VP.t0 260.365
R1 VP.n0 VP.t1 218.72
R2 VP VP.n0 0.241678
R3 VTAIL.n1 VTAIL.t1 64.8228
R4 VTAIL.n3 VTAIL.t0 64.8227
R5 VTAIL.n0 VTAIL.t2 64.8227
R6 VTAIL.n2 VTAIL.t3 64.8227
R7 VTAIL.n1 VTAIL.n0 25.5134
R8 VTAIL.n3 VTAIL.n2 23.7721
R9 VTAIL.n2 VTAIL.n1 1.34102
R10 VTAIL VTAIL.n0 0.963862
R11 VTAIL VTAIL.n3 0.377655
R12 VDD1 VDD1.t0 119.267
R13 VDD1 VDD1.t1 81.995
R14 B.n364 B.n363 585
R15 B.n365 B.n60 585
R16 B.n367 B.n366 585
R17 B.n368 B.n59 585
R18 B.n370 B.n369 585
R19 B.n371 B.n58 585
R20 B.n373 B.n372 585
R21 B.n374 B.n57 585
R22 B.n376 B.n375 585
R23 B.n377 B.n56 585
R24 B.n379 B.n378 585
R25 B.n380 B.n55 585
R26 B.n382 B.n381 585
R27 B.n383 B.n54 585
R28 B.n385 B.n384 585
R29 B.n386 B.n53 585
R30 B.n388 B.n387 585
R31 B.n389 B.n52 585
R32 B.n391 B.n390 585
R33 B.n392 B.n51 585
R34 B.n394 B.n393 585
R35 B.n395 B.n50 585
R36 B.n397 B.n396 585
R37 B.n398 B.n49 585
R38 B.n400 B.n399 585
R39 B.n401 B.n48 585
R40 B.n403 B.n402 585
R41 B.n404 B.n47 585
R42 B.n406 B.n405 585
R43 B.n407 B.n46 585
R44 B.n409 B.n408 585
R45 B.n410 B.n45 585
R46 B.n412 B.n411 585
R47 B.n413 B.n44 585
R48 B.n415 B.n414 585
R49 B.n416 B.n43 585
R50 B.n418 B.n417 585
R51 B.n419 B.n39 585
R52 B.n421 B.n420 585
R53 B.n422 B.n38 585
R54 B.n424 B.n423 585
R55 B.n425 B.n37 585
R56 B.n427 B.n426 585
R57 B.n428 B.n36 585
R58 B.n430 B.n429 585
R59 B.n431 B.n35 585
R60 B.n433 B.n432 585
R61 B.n434 B.n34 585
R62 B.n436 B.n435 585
R63 B.n438 B.n31 585
R64 B.n440 B.n439 585
R65 B.n441 B.n30 585
R66 B.n443 B.n442 585
R67 B.n444 B.n29 585
R68 B.n446 B.n445 585
R69 B.n447 B.n28 585
R70 B.n449 B.n448 585
R71 B.n450 B.n27 585
R72 B.n452 B.n451 585
R73 B.n453 B.n26 585
R74 B.n455 B.n454 585
R75 B.n456 B.n25 585
R76 B.n458 B.n457 585
R77 B.n459 B.n24 585
R78 B.n461 B.n460 585
R79 B.n462 B.n23 585
R80 B.n464 B.n463 585
R81 B.n465 B.n22 585
R82 B.n467 B.n466 585
R83 B.n468 B.n21 585
R84 B.n470 B.n469 585
R85 B.n471 B.n20 585
R86 B.n473 B.n472 585
R87 B.n474 B.n19 585
R88 B.n476 B.n475 585
R89 B.n477 B.n18 585
R90 B.n479 B.n478 585
R91 B.n480 B.n17 585
R92 B.n482 B.n481 585
R93 B.n483 B.n16 585
R94 B.n485 B.n484 585
R95 B.n486 B.n15 585
R96 B.n488 B.n487 585
R97 B.n489 B.n14 585
R98 B.n491 B.n490 585
R99 B.n492 B.n13 585
R100 B.n494 B.n493 585
R101 B.n495 B.n12 585
R102 B.n362 B.n61 585
R103 B.n361 B.n360 585
R104 B.n359 B.n62 585
R105 B.n358 B.n357 585
R106 B.n356 B.n63 585
R107 B.n355 B.n354 585
R108 B.n353 B.n64 585
R109 B.n352 B.n351 585
R110 B.n350 B.n65 585
R111 B.n349 B.n348 585
R112 B.n347 B.n66 585
R113 B.n346 B.n345 585
R114 B.n344 B.n67 585
R115 B.n343 B.n342 585
R116 B.n341 B.n68 585
R117 B.n340 B.n339 585
R118 B.n338 B.n69 585
R119 B.n337 B.n336 585
R120 B.n335 B.n70 585
R121 B.n334 B.n333 585
R122 B.n332 B.n71 585
R123 B.n331 B.n330 585
R124 B.n329 B.n72 585
R125 B.n328 B.n327 585
R126 B.n326 B.n73 585
R127 B.n325 B.n324 585
R128 B.n323 B.n74 585
R129 B.n322 B.n321 585
R130 B.n320 B.n75 585
R131 B.n319 B.n318 585
R132 B.n317 B.n76 585
R133 B.n316 B.n315 585
R134 B.n314 B.n77 585
R135 B.n313 B.n312 585
R136 B.n311 B.n78 585
R137 B.n310 B.n309 585
R138 B.n308 B.n79 585
R139 B.n307 B.n306 585
R140 B.n305 B.n80 585
R141 B.n304 B.n303 585
R142 B.n302 B.n81 585
R143 B.n169 B.n168 585
R144 B.n170 B.n129 585
R145 B.n172 B.n171 585
R146 B.n173 B.n128 585
R147 B.n175 B.n174 585
R148 B.n176 B.n127 585
R149 B.n178 B.n177 585
R150 B.n179 B.n126 585
R151 B.n181 B.n180 585
R152 B.n182 B.n125 585
R153 B.n184 B.n183 585
R154 B.n185 B.n124 585
R155 B.n187 B.n186 585
R156 B.n188 B.n123 585
R157 B.n190 B.n189 585
R158 B.n191 B.n122 585
R159 B.n193 B.n192 585
R160 B.n194 B.n121 585
R161 B.n196 B.n195 585
R162 B.n197 B.n120 585
R163 B.n199 B.n198 585
R164 B.n200 B.n119 585
R165 B.n202 B.n201 585
R166 B.n203 B.n118 585
R167 B.n205 B.n204 585
R168 B.n206 B.n117 585
R169 B.n208 B.n207 585
R170 B.n209 B.n116 585
R171 B.n211 B.n210 585
R172 B.n212 B.n115 585
R173 B.n214 B.n213 585
R174 B.n215 B.n114 585
R175 B.n217 B.n216 585
R176 B.n218 B.n113 585
R177 B.n220 B.n219 585
R178 B.n221 B.n112 585
R179 B.n223 B.n222 585
R180 B.n224 B.n111 585
R181 B.n226 B.n225 585
R182 B.n228 B.n108 585
R183 B.n230 B.n229 585
R184 B.n231 B.n107 585
R185 B.n233 B.n232 585
R186 B.n234 B.n106 585
R187 B.n236 B.n235 585
R188 B.n237 B.n105 585
R189 B.n239 B.n238 585
R190 B.n240 B.n104 585
R191 B.n242 B.n241 585
R192 B.n244 B.n243 585
R193 B.n245 B.n100 585
R194 B.n247 B.n246 585
R195 B.n248 B.n99 585
R196 B.n250 B.n249 585
R197 B.n251 B.n98 585
R198 B.n253 B.n252 585
R199 B.n254 B.n97 585
R200 B.n256 B.n255 585
R201 B.n257 B.n96 585
R202 B.n259 B.n258 585
R203 B.n260 B.n95 585
R204 B.n262 B.n261 585
R205 B.n263 B.n94 585
R206 B.n265 B.n264 585
R207 B.n266 B.n93 585
R208 B.n268 B.n267 585
R209 B.n269 B.n92 585
R210 B.n271 B.n270 585
R211 B.n272 B.n91 585
R212 B.n274 B.n273 585
R213 B.n275 B.n90 585
R214 B.n277 B.n276 585
R215 B.n278 B.n89 585
R216 B.n280 B.n279 585
R217 B.n281 B.n88 585
R218 B.n283 B.n282 585
R219 B.n284 B.n87 585
R220 B.n286 B.n285 585
R221 B.n287 B.n86 585
R222 B.n289 B.n288 585
R223 B.n290 B.n85 585
R224 B.n292 B.n291 585
R225 B.n293 B.n84 585
R226 B.n295 B.n294 585
R227 B.n296 B.n83 585
R228 B.n298 B.n297 585
R229 B.n299 B.n82 585
R230 B.n301 B.n300 585
R231 B.n167 B.n130 585
R232 B.n166 B.n165 585
R233 B.n164 B.n131 585
R234 B.n163 B.n162 585
R235 B.n161 B.n132 585
R236 B.n160 B.n159 585
R237 B.n158 B.n133 585
R238 B.n157 B.n156 585
R239 B.n155 B.n134 585
R240 B.n154 B.n153 585
R241 B.n152 B.n135 585
R242 B.n151 B.n150 585
R243 B.n149 B.n136 585
R244 B.n148 B.n147 585
R245 B.n146 B.n137 585
R246 B.n145 B.n144 585
R247 B.n143 B.n138 585
R248 B.n142 B.n141 585
R249 B.n140 B.n139 585
R250 B.n2 B.n0 585
R251 B.n525 B.n1 585
R252 B.n524 B.n523 585
R253 B.n522 B.n3 585
R254 B.n521 B.n520 585
R255 B.n519 B.n4 585
R256 B.n518 B.n517 585
R257 B.n516 B.n5 585
R258 B.n515 B.n514 585
R259 B.n513 B.n6 585
R260 B.n512 B.n511 585
R261 B.n510 B.n7 585
R262 B.n509 B.n508 585
R263 B.n507 B.n8 585
R264 B.n506 B.n505 585
R265 B.n504 B.n9 585
R266 B.n503 B.n502 585
R267 B.n501 B.n10 585
R268 B.n500 B.n499 585
R269 B.n498 B.n11 585
R270 B.n497 B.n496 585
R271 B.n527 B.n526 585
R272 B.n169 B.n130 511.721
R273 B.n496 B.n495 511.721
R274 B.n302 B.n301 511.721
R275 B.n363 B.n362 511.721
R276 B.n101 B.t0 365.942
R277 B.n109 B.t6 365.942
R278 B.n32 B.t9 365.942
R279 B.n40 B.t3 365.942
R280 B.n165 B.n130 163.367
R281 B.n165 B.n164 163.367
R282 B.n164 B.n163 163.367
R283 B.n163 B.n132 163.367
R284 B.n159 B.n132 163.367
R285 B.n159 B.n158 163.367
R286 B.n158 B.n157 163.367
R287 B.n157 B.n134 163.367
R288 B.n153 B.n134 163.367
R289 B.n153 B.n152 163.367
R290 B.n152 B.n151 163.367
R291 B.n151 B.n136 163.367
R292 B.n147 B.n136 163.367
R293 B.n147 B.n146 163.367
R294 B.n146 B.n145 163.367
R295 B.n145 B.n138 163.367
R296 B.n141 B.n138 163.367
R297 B.n141 B.n140 163.367
R298 B.n140 B.n2 163.367
R299 B.n526 B.n2 163.367
R300 B.n526 B.n525 163.367
R301 B.n525 B.n524 163.367
R302 B.n524 B.n3 163.367
R303 B.n520 B.n3 163.367
R304 B.n520 B.n519 163.367
R305 B.n519 B.n518 163.367
R306 B.n518 B.n5 163.367
R307 B.n514 B.n5 163.367
R308 B.n514 B.n513 163.367
R309 B.n513 B.n512 163.367
R310 B.n512 B.n7 163.367
R311 B.n508 B.n7 163.367
R312 B.n508 B.n507 163.367
R313 B.n507 B.n506 163.367
R314 B.n506 B.n9 163.367
R315 B.n502 B.n9 163.367
R316 B.n502 B.n501 163.367
R317 B.n501 B.n500 163.367
R318 B.n500 B.n11 163.367
R319 B.n496 B.n11 163.367
R320 B.n170 B.n169 163.367
R321 B.n171 B.n170 163.367
R322 B.n171 B.n128 163.367
R323 B.n175 B.n128 163.367
R324 B.n176 B.n175 163.367
R325 B.n177 B.n176 163.367
R326 B.n177 B.n126 163.367
R327 B.n181 B.n126 163.367
R328 B.n182 B.n181 163.367
R329 B.n183 B.n182 163.367
R330 B.n183 B.n124 163.367
R331 B.n187 B.n124 163.367
R332 B.n188 B.n187 163.367
R333 B.n189 B.n188 163.367
R334 B.n189 B.n122 163.367
R335 B.n193 B.n122 163.367
R336 B.n194 B.n193 163.367
R337 B.n195 B.n194 163.367
R338 B.n195 B.n120 163.367
R339 B.n199 B.n120 163.367
R340 B.n200 B.n199 163.367
R341 B.n201 B.n200 163.367
R342 B.n201 B.n118 163.367
R343 B.n205 B.n118 163.367
R344 B.n206 B.n205 163.367
R345 B.n207 B.n206 163.367
R346 B.n207 B.n116 163.367
R347 B.n211 B.n116 163.367
R348 B.n212 B.n211 163.367
R349 B.n213 B.n212 163.367
R350 B.n213 B.n114 163.367
R351 B.n217 B.n114 163.367
R352 B.n218 B.n217 163.367
R353 B.n219 B.n218 163.367
R354 B.n219 B.n112 163.367
R355 B.n223 B.n112 163.367
R356 B.n224 B.n223 163.367
R357 B.n225 B.n224 163.367
R358 B.n225 B.n108 163.367
R359 B.n230 B.n108 163.367
R360 B.n231 B.n230 163.367
R361 B.n232 B.n231 163.367
R362 B.n232 B.n106 163.367
R363 B.n236 B.n106 163.367
R364 B.n237 B.n236 163.367
R365 B.n238 B.n237 163.367
R366 B.n238 B.n104 163.367
R367 B.n242 B.n104 163.367
R368 B.n243 B.n242 163.367
R369 B.n243 B.n100 163.367
R370 B.n247 B.n100 163.367
R371 B.n248 B.n247 163.367
R372 B.n249 B.n248 163.367
R373 B.n249 B.n98 163.367
R374 B.n253 B.n98 163.367
R375 B.n254 B.n253 163.367
R376 B.n255 B.n254 163.367
R377 B.n255 B.n96 163.367
R378 B.n259 B.n96 163.367
R379 B.n260 B.n259 163.367
R380 B.n261 B.n260 163.367
R381 B.n261 B.n94 163.367
R382 B.n265 B.n94 163.367
R383 B.n266 B.n265 163.367
R384 B.n267 B.n266 163.367
R385 B.n267 B.n92 163.367
R386 B.n271 B.n92 163.367
R387 B.n272 B.n271 163.367
R388 B.n273 B.n272 163.367
R389 B.n273 B.n90 163.367
R390 B.n277 B.n90 163.367
R391 B.n278 B.n277 163.367
R392 B.n279 B.n278 163.367
R393 B.n279 B.n88 163.367
R394 B.n283 B.n88 163.367
R395 B.n284 B.n283 163.367
R396 B.n285 B.n284 163.367
R397 B.n285 B.n86 163.367
R398 B.n289 B.n86 163.367
R399 B.n290 B.n289 163.367
R400 B.n291 B.n290 163.367
R401 B.n291 B.n84 163.367
R402 B.n295 B.n84 163.367
R403 B.n296 B.n295 163.367
R404 B.n297 B.n296 163.367
R405 B.n297 B.n82 163.367
R406 B.n301 B.n82 163.367
R407 B.n303 B.n302 163.367
R408 B.n303 B.n80 163.367
R409 B.n307 B.n80 163.367
R410 B.n308 B.n307 163.367
R411 B.n309 B.n308 163.367
R412 B.n309 B.n78 163.367
R413 B.n313 B.n78 163.367
R414 B.n314 B.n313 163.367
R415 B.n315 B.n314 163.367
R416 B.n315 B.n76 163.367
R417 B.n319 B.n76 163.367
R418 B.n320 B.n319 163.367
R419 B.n321 B.n320 163.367
R420 B.n321 B.n74 163.367
R421 B.n325 B.n74 163.367
R422 B.n326 B.n325 163.367
R423 B.n327 B.n326 163.367
R424 B.n327 B.n72 163.367
R425 B.n331 B.n72 163.367
R426 B.n332 B.n331 163.367
R427 B.n333 B.n332 163.367
R428 B.n333 B.n70 163.367
R429 B.n337 B.n70 163.367
R430 B.n338 B.n337 163.367
R431 B.n339 B.n338 163.367
R432 B.n339 B.n68 163.367
R433 B.n343 B.n68 163.367
R434 B.n344 B.n343 163.367
R435 B.n345 B.n344 163.367
R436 B.n345 B.n66 163.367
R437 B.n349 B.n66 163.367
R438 B.n350 B.n349 163.367
R439 B.n351 B.n350 163.367
R440 B.n351 B.n64 163.367
R441 B.n355 B.n64 163.367
R442 B.n356 B.n355 163.367
R443 B.n357 B.n356 163.367
R444 B.n357 B.n62 163.367
R445 B.n361 B.n62 163.367
R446 B.n362 B.n361 163.367
R447 B.n495 B.n494 163.367
R448 B.n494 B.n13 163.367
R449 B.n490 B.n13 163.367
R450 B.n490 B.n489 163.367
R451 B.n489 B.n488 163.367
R452 B.n488 B.n15 163.367
R453 B.n484 B.n15 163.367
R454 B.n484 B.n483 163.367
R455 B.n483 B.n482 163.367
R456 B.n482 B.n17 163.367
R457 B.n478 B.n17 163.367
R458 B.n478 B.n477 163.367
R459 B.n477 B.n476 163.367
R460 B.n476 B.n19 163.367
R461 B.n472 B.n19 163.367
R462 B.n472 B.n471 163.367
R463 B.n471 B.n470 163.367
R464 B.n470 B.n21 163.367
R465 B.n466 B.n21 163.367
R466 B.n466 B.n465 163.367
R467 B.n465 B.n464 163.367
R468 B.n464 B.n23 163.367
R469 B.n460 B.n23 163.367
R470 B.n460 B.n459 163.367
R471 B.n459 B.n458 163.367
R472 B.n458 B.n25 163.367
R473 B.n454 B.n25 163.367
R474 B.n454 B.n453 163.367
R475 B.n453 B.n452 163.367
R476 B.n452 B.n27 163.367
R477 B.n448 B.n27 163.367
R478 B.n448 B.n447 163.367
R479 B.n447 B.n446 163.367
R480 B.n446 B.n29 163.367
R481 B.n442 B.n29 163.367
R482 B.n442 B.n441 163.367
R483 B.n441 B.n440 163.367
R484 B.n440 B.n31 163.367
R485 B.n435 B.n31 163.367
R486 B.n435 B.n434 163.367
R487 B.n434 B.n433 163.367
R488 B.n433 B.n35 163.367
R489 B.n429 B.n35 163.367
R490 B.n429 B.n428 163.367
R491 B.n428 B.n427 163.367
R492 B.n427 B.n37 163.367
R493 B.n423 B.n37 163.367
R494 B.n423 B.n422 163.367
R495 B.n422 B.n421 163.367
R496 B.n421 B.n39 163.367
R497 B.n417 B.n39 163.367
R498 B.n417 B.n416 163.367
R499 B.n416 B.n415 163.367
R500 B.n415 B.n44 163.367
R501 B.n411 B.n44 163.367
R502 B.n411 B.n410 163.367
R503 B.n410 B.n409 163.367
R504 B.n409 B.n46 163.367
R505 B.n405 B.n46 163.367
R506 B.n405 B.n404 163.367
R507 B.n404 B.n403 163.367
R508 B.n403 B.n48 163.367
R509 B.n399 B.n48 163.367
R510 B.n399 B.n398 163.367
R511 B.n398 B.n397 163.367
R512 B.n397 B.n50 163.367
R513 B.n393 B.n50 163.367
R514 B.n393 B.n392 163.367
R515 B.n392 B.n391 163.367
R516 B.n391 B.n52 163.367
R517 B.n387 B.n52 163.367
R518 B.n387 B.n386 163.367
R519 B.n386 B.n385 163.367
R520 B.n385 B.n54 163.367
R521 B.n381 B.n54 163.367
R522 B.n381 B.n380 163.367
R523 B.n380 B.n379 163.367
R524 B.n379 B.n56 163.367
R525 B.n375 B.n56 163.367
R526 B.n375 B.n374 163.367
R527 B.n374 B.n373 163.367
R528 B.n373 B.n58 163.367
R529 B.n369 B.n58 163.367
R530 B.n369 B.n368 163.367
R531 B.n368 B.n367 163.367
R532 B.n367 B.n60 163.367
R533 B.n363 B.n60 163.367
R534 B.n101 B.t2 152.88
R535 B.n40 B.t4 152.88
R536 B.n109 B.t8 152.867
R537 B.n32 B.t10 152.867
R538 B.n102 B.t1 113.704
R539 B.n41 B.t5 113.704
R540 B.n110 B.t7 113.691
R541 B.n33 B.t11 113.691
R542 B.n103 B.n102 59.5399
R543 B.n227 B.n110 59.5399
R544 B.n437 B.n33 59.5399
R545 B.n42 B.n41 59.5399
R546 B.n102 B.n101 39.1763
R547 B.n110 B.n109 39.1763
R548 B.n33 B.n32 39.1763
R549 B.n41 B.n40 39.1763
R550 B.n497 B.n12 33.2493
R551 B.n364 B.n61 33.2493
R552 B.n300 B.n81 33.2493
R553 B.n168 B.n167 33.2493
R554 B B.n527 18.0485
R555 B.n493 B.n12 10.6151
R556 B.n493 B.n492 10.6151
R557 B.n492 B.n491 10.6151
R558 B.n491 B.n14 10.6151
R559 B.n487 B.n14 10.6151
R560 B.n487 B.n486 10.6151
R561 B.n486 B.n485 10.6151
R562 B.n485 B.n16 10.6151
R563 B.n481 B.n16 10.6151
R564 B.n481 B.n480 10.6151
R565 B.n480 B.n479 10.6151
R566 B.n479 B.n18 10.6151
R567 B.n475 B.n18 10.6151
R568 B.n475 B.n474 10.6151
R569 B.n474 B.n473 10.6151
R570 B.n473 B.n20 10.6151
R571 B.n469 B.n20 10.6151
R572 B.n469 B.n468 10.6151
R573 B.n468 B.n467 10.6151
R574 B.n467 B.n22 10.6151
R575 B.n463 B.n22 10.6151
R576 B.n463 B.n462 10.6151
R577 B.n462 B.n461 10.6151
R578 B.n461 B.n24 10.6151
R579 B.n457 B.n24 10.6151
R580 B.n457 B.n456 10.6151
R581 B.n456 B.n455 10.6151
R582 B.n455 B.n26 10.6151
R583 B.n451 B.n26 10.6151
R584 B.n451 B.n450 10.6151
R585 B.n450 B.n449 10.6151
R586 B.n449 B.n28 10.6151
R587 B.n445 B.n28 10.6151
R588 B.n445 B.n444 10.6151
R589 B.n444 B.n443 10.6151
R590 B.n443 B.n30 10.6151
R591 B.n439 B.n30 10.6151
R592 B.n439 B.n438 10.6151
R593 B.n436 B.n34 10.6151
R594 B.n432 B.n34 10.6151
R595 B.n432 B.n431 10.6151
R596 B.n431 B.n430 10.6151
R597 B.n430 B.n36 10.6151
R598 B.n426 B.n36 10.6151
R599 B.n426 B.n425 10.6151
R600 B.n425 B.n424 10.6151
R601 B.n424 B.n38 10.6151
R602 B.n420 B.n419 10.6151
R603 B.n419 B.n418 10.6151
R604 B.n418 B.n43 10.6151
R605 B.n414 B.n43 10.6151
R606 B.n414 B.n413 10.6151
R607 B.n413 B.n412 10.6151
R608 B.n412 B.n45 10.6151
R609 B.n408 B.n45 10.6151
R610 B.n408 B.n407 10.6151
R611 B.n407 B.n406 10.6151
R612 B.n406 B.n47 10.6151
R613 B.n402 B.n47 10.6151
R614 B.n402 B.n401 10.6151
R615 B.n401 B.n400 10.6151
R616 B.n400 B.n49 10.6151
R617 B.n396 B.n49 10.6151
R618 B.n396 B.n395 10.6151
R619 B.n395 B.n394 10.6151
R620 B.n394 B.n51 10.6151
R621 B.n390 B.n51 10.6151
R622 B.n390 B.n389 10.6151
R623 B.n389 B.n388 10.6151
R624 B.n388 B.n53 10.6151
R625 B.n384 B.n53 10.6151
R626 B.n384 B.n383 10.6151
R627 B.n383 B.n382 10.6151
R628 B.n382 B.n55 10.6151
R629 B.n378 B.n55 10.6151
R630 B.n378 B.n377 10.6151
R631 B.n377 B.n376 10.6151
R632 B.n376 B.n57 10.6151
R633 B.n372 B.n57 10.6151
R634 B.n372 B.n371 10.6151
R635 B.n371 B.n370 10.6151
R636 B.n370 B.n59 10.6151
R637 B.n366 B.n59 10.6151
R638 B.n366 B.n365 10.6151
R639 B.n365 B.n364 10.6151
R640 B.n304 B.n81 10.6151
R641 B.n305 B.n304 10.6151
R642 B.n306 B.n305 10.6151
R643 B.n306 B.n79 10.6151
R644 B.n310 B.n79 10.6151
R645 B.n311 B.n310 10.6151
R646 B.n312 B.n311 10.6151
R647 B.n312 B.n77 10.6151
R648 B.n316 B.n77 10.6151
R649 B.n317 B.n316 10.6151
R650 B.n318 B.n317 10.6151
R651 B.n318 B.n75 10.6151
R652 B.n322 B.n75 10.6151
R653 B.n323 B.n322 10.6151
R654 B.n324 B.n323 10.6151
R655 B.n324 B.n73 10.6151
R656 B.n328 B.n73 10.6151
R657 B.n329 B.n328 10.6151
R658 B.n330 B.n329 10.6151
R659 B.n330 B.n71 10.6151
R660 B.n334 B.n71 10.6151
R661 B.n335 B.n334 10.6151
R662 B.n336 B.n335 10.6151
R663 B.n336 B.n69 10.6151
R664 B.n340 B.n69 10.6151
R665 B.n341 B.n340 10.6151
R666 B.n342 B.n341 10.6151
R667 B.n342 B.n67 10.6151
R668 B.n346 B.n67 10.6151
R669 B.n347 B.n346 10.6151
R670 B.n348 B.n347 10.6151
R671 B.n348 B.n65 10.6151
R672 B.n352 B.n65 10.6151
R673 B.n353 B.n352 10.6151
R674 B.n354 B.n353 10.6151
R675 B.n354 B.n63 10.6151
R676 B.n358 B.n63 10.6151
R677 B.n359 B.n358 10.6151
R678 B.n360 B.n359 10.6151
R679 B.n360 B.n61 10.6151
R680 B.n168 B.n129 10.6151
R681 B.n172 B.n129 10.6151
R682 B.n173 B.n172 10.6151
R683 B.n174 B.n173 10.6151
R684 B.n174 B.n127 10.6151
R685 B.n178 B.n127 10.6151
R686 B.n179 B.n178 10.6151
R687 B.n180 B.n179 10.6151
R688 B.n180 B.n125 10.6151
R689 B.n184 B.n125 10.6151
R690 B.n185 B.n184 10.6151
R691 B.n186 B.n185 10.6151
R692 B.n186 B.n123 10.6151
R693 B.n190 B.n123 10.6151
R694 B.n191 B.n190 10.6151
R695 B.n192 B.n191 10.6151
R696 B.n192 B.n121 10.6151
R697 B.n196 B.n121 10.6151
R698 B.n197 B.n196 10.6151
R699 B.n198 B.n197 10.6151
R700 B.n198 B.n119 10.6151
R701 B.n202 B.n119 10.6151
R702 B.n203 B.n202 10.6151
R703 B.n204 B.n203 10.6151
R704 B.n204 B.n117 10.6151
R705 B.n208 B.n117 10.6151
R706 B.n209 B.n208 10.6151
R707 B.n210 B.n209 10.6151
R708 B.n210 B.n115 10.6151
R709 B.n214 B.n115 10.6151
R710 B.n215 B.n214 10.6151
R711 B.n216 B.n215 10.6151
R712 B.n216 B.n113 10.6151
R713 B.n220 B.n113 10.6151
R714 B.n221 B.n220 10.6151
R715 B.n222 B.n221 10.6151
R716 B.n222 B.n111 10.6151
R717 B.n226 B.n111 10.6151
R718 B.n229 B.n228 10.6151
R719 B.n229 B.n107 10.6151
R720 B.n233 B.n107 10.6151
R721 B.n234 B.n233 10.6151
R722 B.n235 B.n234 10.6151
R723 B.n235 B.n105 10.6151
R724 B.n239 B.n105 10.6151
R725 B.n240 B.n239 10.6151
R726 B.n241 B.n240 10.6151
R727 B.n245 B.n244 10.6151
R728 B.n246 B.n245 10.6151
R729 B.n246 B.n99 10.6151
R730 B.n250 B.n99 10.6151
R731 B.n251 B.n250 10.6151
R732 B.n252 B.n251 10.6151
R733 B.n252 B.n97 10.6151
R734 B.n256 B.n97 10.6151
R735 B.n257 B.n256 10.6151
R736 B.n258 B.n257 10.6151
R737 B.n258 B.n95 10.6151
R738 B.n262 B.n95 10.6151
R739 B.n263 B.n262 10.6151
R740 B.n264 B.n263 10.6151
R741 B.n264 B.n93 10.6151
R742 B.n268 B.n93 10.6151
R743 B.n269 B.n268 10.6151
R744 B.n270 B.n269 10.6151
R745 B.n270 B.n91 10.6151
R746 B.n274 B.n91 10.6151
R747 B.n275 B.n274 10.6151
R748 B.n276 B.n275 10.6151
R749 B.n276 B.n89 10.6151
R750 B.n280 B.n89 10.6151
R751 B.n281 B.n280 10.6151
R752 B.n282 B.n281 10.6151
R753 B.n282 B.n87 10.6151
R754 B.n286 B.n87 10.6151
R755 B.n287 B.n286 10.6151
R756 B.n288 B.n287 10.6151
R757 B.n288 B.n85 10.6151
R758 B.n292 B.n85 10.6151
R759 B.n293 B.n292 10.6151
R760 B.n294 B.n293 10.6151
R761 B.n294 B.n83 10.6151
R762 B.n298 B.n83 10.6151
R763 B.n299 B.n298 10.6151
R764 B.n300 B.n299 10.6151
R765 B.n167 B.n166 10.6151
R766 B.n166 B.n131 10.6151
R767 B.n162 B.n131 10.6151
R768 B.n162 B.n161 10.6151
R769 B.n161 B.n160 10.6151
R770 B.n160 B.n133 10.6151
R771 B.n156 B.n133 10.6151
R772 B.n156 B.n155 10.6151
R773 B.n155 B.n154 10.6151
R774 B.n154 B.n135 10.6151
R775 B.n150 B.n135 10.6151
R776 B.n150 B.n149 10.6151
R777 B.n149 B.n148 10.6151
R778 B.n148 B.n137 10.6151
R779 B.n144 B.n137 10.6151
R780 B.n144 B.n143 10.6151
R781 B.n143 B.n142 10.6151
R782 B.n142 B.n139 10.6151
R783 B.n139 B.n0 10.6151
R784 B.n523 B.n1 10.6151
R785 B.n523 B.n522 10.6151
R786 B.n522 B.n521 10.6151
R787 B.n521 B.n4 10.6151
R788 B.n517 B.n4 10.6151
R789 B.n517 B.n516 10.6151
R790 B.n516 B.n515 10.6151
R791 B.n515 B.n6 10.6151
R792 B.n511 B.n6 10.6151
R793 B.n511 B.n510 10.6151
R794 B.n510 B.n509 10.6151
R795 B.n509 B.n8 10.6151
R796 B.n505 B.n8 10.6151
R797 B.n505 B.n504 10.6151
R798 B.n504 B.n503 10.6151
R799 B.n503 B.n10 10.6151
R800 B.n499 B.n10 10.6151
R801 B.n499 B.n498 10.6151
R802 B.n498 B.n497 10.6151
R803 B.n438 B.n437 9.36635
R804 B.n420 B.n42 9.36635
R805 B.n227 B.n226 9.36635
R806 B.n244 B.n103 9.36635
R807 B.n527 B.n0 2.81026
R808 B.n527 B.n1 2.81026
R809 B.n437 B.n436 1.24928
R810 B.n42 B.n38 1.24928
R811 B.n228 B.n227 1.24928
R812 B.n241 B.n103 1.24928
R813 VN VN.t1 260.555
R814 VN VN.t0 218.962
R815 VDD2.n0 VDD2.t1 118.308
R816 VDD2.n0 VDD2.t0 81.5015
R817 VDD2 VDD2.n0 0.494034
C0 VN B 0.886826f
C1 B VTAIL 3.08919f
C2 VN VDD2 2.41416f
C3 VP w_n1778_n3210# 2.59377f
C4 VTAIL VDD2 4.84962f
C5 B VDD2 1.53863f
C6 VDD1 w_n1778_n3210# 1.62355f
C7 VN VP 4.88505f
C8 VTAIL VP 2.06646f
C9 VN VDD1 0.147705f
C10 B VP 1.2523f
C11 VTAIL VDD1 4.80614f
C12 VP VDD2 0.29485f
C13 B VDD1 1.51659f
C14 VN w_n1778_n3210# 2.36925f
C15 VDD1 VDD2 0.567491f
C16 VTAIL w_n1778_n3210# 2.66667f
C17 B w_n1778_n3210# 7.60403f
C18 w_n1778_n3210# VDD2 1.63851f
C19 VDD1 VP 2.55834f
C20 VN VTAIL 2.05209f
C21 VDD2 VSUBS 0.791205f
C22 VDD1 VSUBS 4.141376f
C23 VTAIL VSUBS 0.872073f
C24 VN VSUBS 7.59708f
C25 VP VSUBS 1.394751f
C26 B VSUBS 3.152931f
C27 w_n1778_n3210# VSUBS 70.344795f
C28 VDD2.t1 VSUBS 2.27095f
C29 VDD2.t0 VSUBS 1.80376f
C30 VDD2.n0 VSUBS 3.03652f
C31 VN.t0 VSUBS 2.87146f
C32 VN.t1 VSUBS 3.35151f
C33 B.n0 VSUBS 0.004257f
C34 B.n1 VSUBS 0.004257f
C35 B.n2 VSUBS 0.006731f
C36 B.n3 VSUBS 0.006731f
C37 B.n4 VSUBS 0.006731f
C38 B.n5 VSUBS 0.006731f
C39 B.n6 VSUBS 0.006731f
C40 B.n7 VSUBS 0.006731f
C41 B.n8 VSUBS 0.006731f
C42 B.n9 VSUBS 0.006731f
C43 B.n10 VSUBS 0.006731f
C44 B.n11 VSUBS 0.006731f
C45 B.n12 VSUBS 0.016252f
C46 B.n13 VSUBS 0.006731f
C47 B.n14 VSUBS 0.006731f
C48 B.n15 VSUBS 0.006731f
C49 B.n16 VSUBS 0.006731f
C50 B.n17 VSUBS 0.006731f
C51 B.n18 VSUBS 0.006731f
C52 B.n19 VSUBS 0.006731f
C53 B.n20 VSUBS 0.006731f
C54 B.n21 VSUBS 0.006731f
C55 B.n22 VSUBS 0.006731f
C56 B.n23 VSUBS 0.006731f
C57 B.n24 VSUBS 0.006731f
C58 B.n25 VSUBS 0.006731f
C59 B.n26 VSUBS 0.006731f
C60 B.n27 VSUBS 0.006731f
C61 B.n28 VSUBS 0.006731f
C62 B.n29 VSUBS 0.006731f
C63 B.n30 VSUBS 0.006731f
C64 B.n31 VSUBS 0.006731f
C65 B.t11 VSUBS 0.348635f
C66 B.t10 VSUBS 0.362927f
C67 B.t9 VSUBS 0.80799f
C68 B.n32 VSUBS 0.169656f
C69 B.n33 VSUBS 0.06537f
C70 B.n34 VSUBS 0.006731f
C71 B.n35 VSUBS 0.006731f
C72 B.n36 VSUBS 0.006731f
C73 B.n37 VSUBS 0.006731f
C74 B.n38 VSUBS 0.003762f
C75 B.n39 VSUBS 0.006731f
C76 B.t5 VSUBS 0.348629f
C77 B.t4 VSUBS 0.362922f
C78 B.t3 VSUBS 0.80799f
C79 B.n40 VSUBS 0.169662f
C80 B.n41 VSUBS 0.065376f
C81 B.n42 VSUBS 0.015596f
C82 B.n43 VSUBS 0.006731f
C83 B.n44 VSUBS 0.006731f
C84 B.n45 VSUBS 0.006731f
C85 B.n46 VSUBS 0.006731f
C86 B.n47 VSUBS 0.006731f
C87 B.n48 VSUBS 0.006731f
C88 B.n49 VSUBS 0.006731f
C89 B.n50 VSUBS 0.006731f
C90 B.n51 VSUBS 0.006731f
C91 B.n52 VSUBS 0.006731f
C92 B.n53 VSUBS 0.006731f
C93 B.n54 VSUBS 0.006731f
C94 B.n55 VSUBS 0.006731f
C95 B.n56 VSUBS 0.006731f
C96 B.n57 VSUBS 0.006731f
C97 B.n58 VSUBS 0.006731f
C98 B.n59 VSUBS 0.006731f
C99 B.n60 VSUBS 0.006731f
C100 B.n61 VSUBS 0.016404f
C101 B.n62 VSUBS 0.006731f
C102 B.n63 VSUBS 0.006731f
C103 B.n64 VSUBS 0.006731f
C104 B.n65 VSUBS 0.006731f
C105 B.n66 VSUBS 0.006731f
C106 B.n67 VSUBS 0.006731f
C107 B.n68 VSUBS 0.006731f
C108 B.n69 VSUBS 0.006731f
C109 B.n70 VSUBS 0.006731f
C110 B.n71 VSUBS 0.006731f
C111 B.n72 VSUBS 0.006731f
C112 B.n73 VSUBS 0.006731f
C113 B.n74 VSUBS 0.006731f
C114 B.n75 VSUBS 0.006731f
C115 B.n76 VSUBS 0.006731f
C116 B.n77 VSUBS 0.006731f
C117 B.n78 VSUBS 0.006731f
C118 B.n79 VSUBS 0.006731f
C119 B.n80 VSUBS 0.006731f
C120 B.n81 VSUBS 0.015623f
C121 B.n82 VSUBS 0.006731f
C122 B.n83 VSUBS 0.006731f
C123 B.n84 VSUBS 0.006731f
C124 B.n85 VSUBS 0.006731f
C125 B.n86 VSUBS 0.006731f
C126 B.n87 VSUBS 0.006731f
C127 B.n88 VSUBS 0.006731f
C128 B.n89 VSUBS 0.006731f
C129 B.n90 VSUBS 0.006731f
C130 B.n91 VSUBS 0.006731f
C131 B.n92 VSUBS 0.006731f
C132 B.n93 VSUBS 0.006731f
C133 B.n94 VSUBS 0.006731f
C134 B.n95 VSUBS 0.006731f
C135 B.n96 VSUBS 0.006731f
C136 B.n97 VSUBS 0.006731f
C137 B.n98 VSUBS 0.006731f
C138 B.n99 VSUBS 0.006731f
C139 B.n100 VSUBS 0.006731f
C140 B.t1 VSUBS 0.348629f
C141 B.t2 VSUBS 0.362922f
C142 B.t0 VSUBS 0.80799f
C143 B.n101 VSUBS 0.169662f
C144 B.n102 VSUBS 0.065376f
C145 B.n103 VSUBS 0.015596f
C146 B.n104 VSUBS 0.006731f
C147 B.n105 VSUBS 0.006731f
C148 B.n106 VSUBS 0.006731f
C149 B.n107 VSUBS 0.006731f
C150 B.n108 VSUBS 0.006731f
C151 B.t7 VSUBS 0.348635f
C152 B.t8 VSUBS 0.362927f
C153 B.t6 VSUBS 0.80799f
C154 B.n109 VSUBS 0.169656f
C155 B.n110 VSUBS 0.06537f
C156 B.n111 VSUBS 0.006731f
C157 B.n112 VSUBS 0.006731f
C158 B.n113 VSUBS 0.006731f
C159 B.n114 VSUBS 0.006731f
C160 B.n115 VSUBS 0.006731f
C161 B.n116 VSUBS 0.006731f
C162 B.n117 VSUBS 0.006731f
C163 B.n118 VSUBS 0.006731f
C164 B.n119 VSUBS 0.006731f
C165 B.n120 VSUBS 0.006731f
C166 B.n121 VSUBS 0.006731f
C167 B.n122 VSUBS 0.006731f
C168 B.n123 VSUBS 0.006731f
C169 B.n124 VSUBS 0.006731f
C170 B.n125 VSUBS 0.006731f
C171 B.n126 VSUBS 0.006731f
C172 B.n127 VSUBS 0.006731f
C173 B.n128 VSUBS 0.006731f
C174 B.n129 VSUBS 0.006731f
C175 B.n130 VSUBS 0.015623f
C176 B.n131 VSUBS 0.006731f
C177 B.n132 VSUBS 0.006731f
C178 B.n133 VSUBS 0.006731f
C179 B.n134 VSUBS 0.006731f
C180 B.n135 VSUBS 0.006731f
C181 B.n136 VSUBS 0.006731f
C182 B.n137 VSUBS 0.006731f
C183 B.n138 VSUBS 0.006731f
C184 B.n139 VSUBS 0.006731f
C185 B.n140 VSUBS 0.006731f
C186 B.n141 VSUBS 0.006731f
C187 B.n142 VSUBS 0.006731f
C188 B.n143 VSUBS 0.006731f
C189 B.n144 VSUBS 0.006731f
C190 B.n145 VSUBS 0.006731f
C191 B.n146 VSUBS 0.006731f
C192 B.n147 VSUBS 0.006731f
C193 B.n148 VSUBS 0.006731f
C194 B.n149 VSUBS 0.006731f
C195 B.n150 VSUBS 0.006731f
C196 B.n151 VSUBS 0.006731f
C197 B.n152 VSUBS 0.006731f
C198 B.n153 VSUBS 0.006731f
C199 B.n154 VSUBS 0.006731f
C200 B.n155 VSUBS 0.006731f
C201 B.n156 VSUBS 0.006731f
C202 B.n157 VSUBS 0.006731f
C203 B.n158 VSUBS 0.006731f
C204 B.n159 VSUBS 0.006731f
C205 B.n160 VSUBS 0.006731f
C206 B.n161 VSUBS 0.006731f
C207 B.n162 VSUBS 0.006731f
C208 B.n163 VSUBS 0.006731f
C209 B.n164 VSUBS 0.006731f
C210 B.n165 VSUBS 0.006731f
C211 B.n166 VSUBS 0.006731f
C212 B.n167 VSUBS 0.015623f
C213 B.n168 VSUBS 0.016252f
C214 B.n169 VSUBS 0.016252f
C215 B.n170 VSUBS 0.006731f
C216 B.n171 VSUBS 0.006731f
C217 B.n172 VSUBS 0.006731f
C218 B.n173 VSUBS 0.006731f
C219 B.n174 VSUBS 0.006731f
C220 B.n175 VSUBS 0.006731f
C221 B.n176 VSUBS 0.006731f
C222 B.n177 VSUBS 0.006731f
C223 B.n178 VSUBS 0.006731f
C224 B.n179 VSUBS 0.006731f
C225 B.n180 VSUBS 0.006731f
C226 B.n181 VSUBS 0.006731f
C227 B.n182 VSUBS 0.006731f
C228 B.n183 VSUBS 0.006731f
C229 B.n184 VSUBS 0.006731f
C230 B.n185 VSUBS 0.006731f
C231 B.n186 VSUBS 0.006731f
C232 B.n187 VSUBS 0.006731f
C233 B.n188 VSUBS 0.006731f
C234 B.n189 VSUBS 0.006731f
C235 B.n190 VSUBS 0.006731f
C236 B.n191 VSUBS 0.006731f
C237 B.n192 VSUBS 0.006731f
C238 B.n193 VSUBS 0.006731f
C239 B.n194 VSUBS 0.006731f
C240 B.n195 VSUBS 0.006731f
C241 B.n196 VSUBS 0.006731f
C242 B.n197 VSUBS 0.006731f
C243 B.n198 VSUBS 0.006731f
C244 B.n199 VSUBS 0.006731f
C245 B.n200 VSUBS 0.006731f
C246 B.n201 VSUBS 0.006731f
C247 B.n202 VSUBS 0.006731f
C248 B.n203 VSUBS 0.006731f
C249 B.n204 VSUBS 0.006731f
C250 B.n205 VSUBS 0.006731f
C251 B.n206 VSUBS 0.006731f
C252 B.n207 VSUBS 0.006731f
C253 B.n208 VSUBS 0.006731f
C254 B.n209 VSUBS 0.006731f
C255 B.n210 VSUBS 0.006731f
C256 B.n211 VSUBS 0.006731f
C257 B.n212 VSUBS 0.006731f
C258 B.n213 VSUBS 0.006731f
C259 B.n214 VSUBS 0.006731f
C260 B.n215 VSUBS 0.006731f
C261 B.n216 VSUBS 0.006731f
C262 B.n217 VSUBS 0.006731f
C263 B.n218 VSUBS 0.006731f
C264 B.n219 VSUBS 0.006731f
C265 B.n220 VSUBS 0.006731f
C266 B.n221 VSUBS 0.006731f
C267 B.n222 VSUBS 0.006731f
C268 B.n223 VSUBS 0.006731f
C269 B.n224 VSUBS 0.006731f
C270 B.n225 VSUBS 0.006731f
C271 B.n226 VSUBS 0.006335f
C272 B.n227 VSUBS 0.015596f
C273 B.n228 VSUBS 0.003762f
C274 B.n229 VSUBS 0.006731f
C275 B.n230 VSUBS 0.006731f
C276 B.n231 VSUBS 0.006731f
C277 B.n232 VSUBS 0.006731f
C278 B.n233 VSUBS 0.006731f
C279 B.n234 VSUBS 0.006731f
C280 B.n235 VSUBS 0.006731f
C281 B.n236 VSUBS 0.006731f
C282 B.n237 VSUBS 0.006731f
C283 B.n238 VSUBS 0.006731f
C284 B.n239 VSUBS 0.006731f
C285 B.n240 VSUBS 0.006731f
C286 B.n241 VSUBS 0.003762f
C287 B.n242 VSUBS 0.006731f
C288 B.n243 VSUBS 0.006731f
C289 B.n244 VSUBS 0.006335f
C290 B.n245 VSUBS 0.006731f
C291 B.n246 VSUBS 0.006731f
C292 B.n247 VSUBS 0.006731f
C293 B.n248 VSUBS 0.006731f
C294 B.n249 VSUBS 0.006731f
C295 B.n250 VSUBS 0.006731f
C296 B.n251 VSUBS 0.006731f
C297 B.n252 VSUBS 0.006731f
C298 B.n253 VSUBS 0.006731f
C299 B.n254 VSUBS 0.006731f
C300 B.n255 VSUBS 0.006731f
C301 B.n256 VSUBS 0.006731f
C302 B.n257 VSUBS 0.006731f
C303 B.n258 VSUBS 0.006731f
C304 B.n259 VSUBS 0.006731f
C305 B.n260 VSUBS 0.006731f
C306 B.n261 VSUBS 0.006731f
C307 B.n262 VSUBS 0.006731f
C308 B.n263 VSUBS 0.006731f
C309 B.n264 VSUBS 0.006731f
C310 B.n265 VSUBS 0.006731f
C311 B.n266 VSUBS 0.006731f
C312 B.n267 VSUBS 0.006731f
C313 B.n268 VSUBS 0.006731f
C314 B.n269 VSUBS 0.006731f
C315 B.n270 VSUBS 0.006731f
C316 B.n271 VSUBS 0.006731f
C317 B.n272 VSUBS 0.006731f
C318 B.n273 VSUBS 0.006731f
C319 B.n274 VSUBS 0.006731f
C320 B.n275 VSUBS 0.006731f
C321 B.n276 VSUBS 0.006731f
C322 B.n277 VSUBS 0.006731f
C323 B.n278 VSUBS 0.006731f
C324 B.n279 VSUBS 0.006731f
C325 B.n280 VSUBS 0.006731f
C326 B.n281 VSUBS 0.006731f
C327 B.n282 VSUBS 0.006731f
C328 B.n283 VSUBS 0.006731f
C329 B.n284 VSUBS 0.006731f
C330 B.n285 VSUBS 0.006731f
C331 B.n286 VSUBS 0.006731f
C332 B.n287 VSUBS 0.006731f
C333 B.n288 VSUBS 0.006731f
C334 B.n289 VSUBS 0.006731f
C335 B.n290 VSUBS 0.006731f
C336 B.n291 VSUBS 0.006731f
C337 B.n292 VSUBS 0.006731f
C338 B.n293 VSUBS 0.006731f
C339 B.n294 VSUBS 0.006731f
C340 B.n295 VSUBS 0.006731f
C341 B.n296 VSUBS 0.006731f
C342 B.n297 VSUBS 0.006731f
C343 B.n298 VSUBS 0.006731f
C344 B.n299 VSUBS 0.006731f
C345 B.n300 VSUBS 0.016252f
C346 B.n301 VSUBS 0.016252f
C347 B.n302 VSUBS 0.015623f
C348 B.n303 VSUBS 0.006731f
C349 B.n304 VSUBS 0.006731f
C350 B.n305 VSUBS 0.006731f
C351 B.n306 VSUBS 0.006731f
C352 B.n307 VSUBS 0.006731f
C353 B.n308 VSUBS 0.006731f
C354 B.n309 VSUBS 0.006731f
C355 B.n310 VSUBS 0.006731f
C356 B.n311 VSUBS 0.006731f
C357 B.n312 VSUBS 0.006731f
C358 B.n313 VSUBS 0.006731f
C359 B.n314 VSUBS 0.006731f
C360 B.n315 VSUBS 0.006731f
C361 B.n316 VSUBS 0.006731f
C362 B.n317 VSUBS 0.006731f
C363 B.n318 VSUBS 0.006731f
C364 B.n319 VSUBS 0.006731f
C365 B.n320 VSUBS 0.006731f
C366 B.n321 VSUBS 0.006731f
C367 B.n322 VSUBS 0.006731f
C368 B.n323 VSUBS 0.006731f
C369 B.n324 VSUBS 0.006731f
C370 B.n325 VSUBS 0.006731f
C371 B.n326 VSUBS 0.006731f
C372 B.n327 VSUBS 0.006731f
C373 B.n328 VSUBS 0.006731f
C374 B.n329 VSUBS 0.006731f
C375 B.n330 VSUBS 0.006731f
C376 B.n331 VSUBS 0.006731f
C377 B.n332 VSUBS 0.006731f
C378 B.n333 VSUBS 0.006731f
C379 B.n334 VSUBS 0.006731f
C380 B.n335 VSUBS 0.006731f
C381 B.n336 VSUBS 0.006731f
C382 B.n337 VSUBS 0.006731f
C383 B.n338 VSUBS 0.006731f
C384 B.n339 VSUBS 0.006731f
C385 B.n340 VSUBS 0.006731f
C386 B.n341 VSUBS 0.006731f
C387 B.n342 VSUBS 0.006731f
C388 B.n343 VSUBS 0.006731f
C389 B.n344 VSUBS 0.006731f
C390 B.n345 VSUBS 0.006731f
C391 B.n346 VSUBS 0.006731f
C392 B.n347 VSUBS 0.006731f
C393 B.n348 VSUBS 0.006731f
C394 B.n349 VSUBS 0.006731f
C395 B.n350 VSUBS 0.006731f
C396 B.n351 VSUBS 0.006731f
C397 B.n352 VSUBS 0.006731f
C398 B.n353 VSUBS 0.006731f
C399 B.n354 VSUBS 0.006731f
C400 B.n355 VSUBS 0.006731f
C401 B.n356 VSUBS 0.006731f
C402 B.n357 VSUBS 0.006731f
C403 B.n358 VSUBS 0.006731f
C404 B.n359 VSUBS 0.006731f
C405 B.n360 VSUBS 0.006731f
C406 B.n361 VSUBS 0.006731f
C407 B.n362 VSUBS 0.015623f
C408 B.n363 VSUBS 0.016252f
C409 B.n364 VSUBS 0.015471f
C410 B.n365 VSUBS 0.006731f
C411 B.n366 VSUBS 0.006731f
C412 B.n367 VSUBS 0.006731f
C413 B.n368 VSUBS 0.006731f
C414 B.n369 VSUBS 0.006731f
C415 B.n370 VSUBS 0.006731f
C416 B.n371 VSUBS 0.006731f
C417 B.n372 VSUBS 0.006731f
C418 B.n373 VSUBS 0.006731f
C419 B.n374 VSUBS 0.006731f
C420 B.n375 VSUBS 0.006731f
C421 B.n376 VSUBS 0.006731f
C422 B.n377 VSUBS 0.006731f
C423 B.n378 VSUBS 0.006731f
C424 B.n379 VSUBS 0.006731f
C425 B.n380 VSUBS 0.006731f
C426 B.n381 VSUBS 0.006731f
C427 B.n382 VSUBS 0.006731f
C428 B.n383 VSUBS 0.006731f
C429 B.n384 VSUBS 0.006731f
C430 B.n385 VSUBS 0.006731f
C431 B.n386 VSUBS 0.006731f
C432 B.n387 VSUBS 0.006731f
C433 B.n388 VSUBS 0.006731f
C434 B.n389 VSUBS 0.006731f
C435 B.n390 VSUBS 0.006731f
C436 B.n391 VSUBS 0.006731f
C437 B.n392 VSUBS 0.006731f
C438 B.n393 VSUBS 0.006731f
C439 B.n394 VSUBS 0.006731f
C440 B.n395 VSUBS 0.006731f
C441 B.n396 VSUBS 0.006731f
C442 B.n397 VSUBS 0.006731f
C443 B.n398 VSUBS 0.006731f
C444 B.n399 VSUBS 0.006731f
C445 B.n400 VSUBS 0.006731f
C446 B.n401 VSUBS 0.006731f
C447 B.n402 VSUBS 0.006731f
C448 B.n403 VSUBS 0.006731f
C449 B.n404 VSUBS 0.006731f
C450 B.n405 VSUBS 0.006731f
C451 B.n406 VSUBS 0.006731f
C452 B.n407 VSUBS 0.006731f
C453 B.n408 VSUBS 0.006731f
C454 B.n409 VSUBS 0.006731f
C455 B.n410 VSUBS 0.006731f
C456 B.n411 VSUBS 0.006731f
C457 B.n412 VSUBS 0.006731f
C458 B.n413 VSUBS 0.006731f
C459 B.n414 VSUBS 0.006731f
C460 B.n415 VSUBS 0.006731f
C461 B.n416 VSUBS 0.006731f
C462 B.n417 VSUBS 0.006731f
C463 B.n418 VSUBS 0.006731f
C464 B.n419 VSUBS 0.006731f
C465 B.n420 VSUBS 0.006335f
C466 B.n421 VSUBS 0.006731f
C467 B.n422 VSUBS 0.006731f
C468 B.n423 VSUBS 0.006731f
C469 B.n424 VSUBS 0.006731f
C470 B.n425 VSUBS 0.006731f
C471 B.n426 VSUBS 0.006731f
C472 B.n427 VSUBS 0.006731f
C473 B.n428 VSUBS 0.006731f
C474 B.n429 VSUBS 0.006731f
C475 B.n430 VSUBS 0.006731f
C476 B.n431 VSUBS 0.006731f
C477 B.n432 VSUBS 0.006731f
C478 B.n433 VSUBS 0.006731f
C479 B.n434 VSUBS 0.006731f
C480 B.n435 VSUBS 0.006731f
C481 B.n436 VSUBS 0.003762f
C482 B.n437 VSUBS 0.015596f
C483 B.n438 VSUBS 0.006335f
C484 B.n439 VSUBS 0.006731f
C485 B.n440 VSUBS 0.006731f
C486 B.n441 VSUBS 0.006731f
C487 B.n442 VSUBS 0.006731f
C488 B.n443 VSUBS 0.006731f
C489 B.n444 VSUBS 0.006731f
C490 B.n445 VSUBS 0.006731f
C491 B.n446 VSUBS 0.006731f
C492 B.n447 VSUBS 0.006731f
C493 B.n448 VSUBS 0.006731f
C494 B.n449 VSUBS 0.006731f
C495 B.n450 VSUBS 0.006731f
C496 B.n451 VSUBS 0.006731f
C497 B.n452 VSUBS 0.006731f
C498 B.n453 VSUBS 0.006731f
C499 B.n454 VSUBS 0.006731f
C500 B.n455 VSUBS 0.006731f
C501 B.n456 VSUBS 0.006731f
C502 B.n457 VSUBS 0.006731f
C503 B.n458 VSUBS 0.006731f
C504 B.n459 VSUBS 0.006731f
C505 B.n460 VSUBS 0.006731f
C506 B.n461 VSUBS 0.006731f
C507 B.n462 VSUBS 0.006731f
C508 B.n463 VSUBS 0.006731f
C509 B.n464 VSUBS 0.006731f
C510 B.n465 VSUBS 0.006731f
C511 B.n466 VSUBS 0.006731f
C512 B.n467 VSUBS 0.006731f
C513 B.n468 VSUBS 0.006731f
C514 B.n469 VSUBS 0.006731f
C515 B.n470 VSUBS 0.006731f
C516 B.n471 VSUBS 0.006731f
C517 B.n472 VSUBS 0.006731f
C518 B.n473 VSUBS 0.006731f
C519 B.n474 VSUBS 0.006731f
C520 B.n475 VSUBS 0.006731f
C521 B.n476 VSUBS 0.006731f
C522 B.n477 VSUBS 0.006731f
C523 B.n478 VSUBS 0.006731f
C524 B.n479 VSUBS 0.006731f
C525 B.n480 VSUBS 0.006731f
C526 B.n481 VSUBS 0.006731f
C527 B.n482 VSUBS 0.006731f
C528 B.n483 VSUBS 0.006731f
C529 B.n484 VSUBS 0.006731f
C530 B.n485 VSUBS 0.006731f
C531 B.n486 VSUBS 0.006731f
C532 B.n487 VSUBS 0.006731f
C533 B.n488 VSUBS 0.006731f
C534 B.n489 VSUBS 0.006731f
C535 B.n490 VSUBS 0.006731f
C536 B.n491 VSUBS 0.006731f
C537 B.n492 VSUBS 0.006731f
C538 B.n493 VSUBS 0.006731f
C539 B.n494 VSUBS 0.006731f
C540 B.n495 VSUBS 0.016252f
C541 B.n496 VSUBS 0.015623f
C542 B.n497 VSUBS 0.015623f
C543 B.n498 VSUBS 0.006731f
C544 B.n499 VSUBS 0.006731f
C545 B.n500 VSUBS 0.006731f
C546 B.n501 VSUBS 0.006731f
C547 B.n502 VSUBS 0.006731f
C548 B.n503 VSUBS 0.006731f
C549 B.n504 VSUBS 0.006731f
C550 B.n505 VSUBS 0.006731f
C551 B.n506 VSUBS 0.006731f
C552 B.n507 VSUBS 0.006731f
C553 B.n508 VSUBS 0.006731f
C554 B.n509 VSUBS 0.006731f
C555 B.n510 VSUBS 0.006731f
C556 B.n511 VSUBS 0.006731f
C557 B.n512 VSUBS 0.006731f
C558 B.n513 VSUBS 0.006731f
C559 B.n514 VSUBS 0.006731f
C560 B.n515 VSUBS 0.006731f
C561 B.n516 VSUBS 0.006731f
C562 B.n517 VSUBS 0.006731f
C563 B.n518 VSUBS 0.006731f
C564 B.n519 VSUBS 0.006731f
C565 B.n520 VSUBS 0.006731f
C566 B.n521 VSUBS 0.006731f
C567 B.n522 VSUBS 0.006731f
C568 B.n523 VSUBS 0.006731f
C569 B.n524 VSUBS 0.006731f
C570 B.n525 VSUBS 0.006731f
C571 B.n526 VSUBS 0.006731f
C572 B.n527 VSUBS 0.015242f
C573 VDD1.t1 VSUBS 1.83781f
C574 VDD1.t0 VSUBS 2.33768f
C575 VTAIL.t2 VSUBS 2.47796f
C576 VTAIL.n0 VSUBS 2.46867f
C577 VTAIL.t1 VSUBS 2.47798f
C578 VTAIL.n1 VSUBS 2.50429f
C579 VTAIL.t3 VSUBS 2.47796f
C580 VTAIL.n2 VSUBS 2.33977f
C581 VTAIL.t0 VSUBS 2.47796f
C582 VTAIL.n3 VSUBS 2.24874f
C583 VP.t0 VSUBS 3.47998f
C584 VP.t1 VSUBS 2.98536f
C585 VP.n0 VSUBS 5.66064f
.ends

