* NGSPICE file created from diff_pair_sample_0199.ext - technology: sky130A

.subckt diff_pair_sample_0199 VTAIL VN VP B VDD2 VDD1
X0 B.t17 B.t15 B.t16 B.t5 sky130_fd_pr__nfet_01v8 ad=0.5616 pd=3.66 as=0 ps=0 w=1.44 l=3.89
X1 VDD2.t3 VN.t0 VTAIL.t7 B.t3 sky130_fd_pr__nfet_01v8 ad=0.2376 pd=1.77 as=0.5616 ps=3.66 w=1.44 l=3.89
X2 B.t14 B.t12 B.t13 B.t9 sky130_fd_pr__nfet_01v8 ad=0.5616 pd=3.66 as=0 ps=0 w=1.44 l=3.89
X3 VTAIL.t1 VP.t0 VDD1.t3 B.t2 sky130_fd_pr__nfet_01v8 ad=0.5616 pd=3.66 as=0.2376 ps=1.77 w=1.44 l=3.89
X4 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=0.5616 pd=3.66 as=0 ps=0 w=1.44 l=3.89
X5 VDD1.t2 VP.t1 VTAIL.t2 B.t3 sky130_fd_pr__nfet_01v8 ad=0.2376 pd=1.77 as=0.5616 ps=3.66 w=1.44 l=3.89
X6 VDD2.t2 VN.t1 VTAIL.t6 B.t0 sky130_fd_pr__nfet_01v8 ad=0.2376 pd=1.77 as=0.5616 ps=3.66 w=1.44 l=3.89
X7 VTAIL.t3 VP.t2 VDD1.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=0.5616 pd=3.66 as=0.2376 ps=1.77 w=1.44 l=3.89
X8 B.t7 B.t4 B.t6 B.t5 sky130_fd_pr__nfet_01v8 ad=0.5616 pd=3.66 as=0 ps=0 w=1.44 l=3.89
X9 VDD1.t0 VP.t3 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=0.2376 pd=1.77 as=0.5616 ps=3.66 w=1.44 l=3.89
X10 VTAIL.t5 VN.t2 VDD2.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=0.5616 pd=3.66 as=0.2376 ps=1.77 w=1.44 l=3.89
X11 VTAIL.t4 VN.t3 VDD2.t0 B.t2 sky130_fd_pr__nfet_01v8 ad=0.5616 pd=3.66 as=0.2376 ps=1.77 w=1.44 l=3.89
R0 B.n532 B.n531 585
R1 B.n533 B.n532 585
R2 B.n165 B.n100 585
R3 B.n164 B.n163 585
R4 B.n162 B.n161 585
R5 B.n160 B.n159 585
R6 B.n158 B.n157 585
R7 B.n156 B.n155 585
R8 B.n154 B.n153 585
R9 B.n152 B.n151 585
R10 B.n150 B.n149 585
R11 B.n148 B.n147 585
R12 B.n146 B.n145 585
R13 B.n144 B.n143 585
R14 B.n142 B.n141 585
R15 B.n140 B.n139 585
R16 B.n138 B.n137 585
R17 B.n136 B.n135 585
R18 B.n134 B.n133 585
R19 B.n132 B.n131 585
R20 B.n130 B.n129 585
R21 B.n127 B.n126 585
R22 B.n125 B.n124 585
R23 B.n123 B.n122 585
R24 B.n121 B.n120 585
R25 B.n119 B.n118 585
R26 B.n117 B.n116 585
R27 B.n115 B.n114 585
R28 B.n113 B.n112 585
R29 B.n111 B.n110 585
R30 B.n109 B.n108 585
R31 B.n107 B.n106 585
R32 B.n530 B.n84 585
R33 B.n534 B.n84 585
R34 B.n529 B.n83 585
R35 B.n535 B.n83 585
R36 B.n528 B.n527 585
R37 B.n527 B.n79 585
R38 B.n526 B.n78 585
R39 B.n541 B.n78 585
R40 B.n525 B.n77 585
R41 B.n542 B.n77 585
R42 B.n524 B.n76 585
R43 B.n543 B.n76 585
R44 B.n523 B.n522 585
R45 B.n522 B.n72 585
R46 B.n521 B.n71 585
R47 B.n549 B.n71 585
R48 B.n520 B.n70 585
R49 B.n550 B.n70 585
R50 B.n519 B.n69 585
R51 B.n551 B.n69 585
R52 B.n518 B.n517 585
R53 B.n517 B.n65 585
R54 B.n516 B.n64 585
R55 B.n557 B.n64 585
R56 B.n515 B.n63 585
R57 B.n558 B.n63 585
R58 B.n514 B.n62 585
R59 B.n559 B.n62 585
R60 B.n513 B.n512 585
R61 B.n512 B.n58 585
R62 B.n511 B.n57 585
R63 B.n565 B.n57 585
R64 B.n510 B.n56 585
R65 B.n566 B.n56 585
R66 B.n509 B.n55 585
R67 B.n567 B.n55 585
R68 B.n508 B.n507 585
R69 B.n507 B.n51 585
R70 B.n506 B.n50 585
R71 B.n573 B.n50 585
R72 B.n505 B.n49 585
R73 B.n574 B.n49 585
R74 B.n504 B.n48 585
R75 B.n575 B.n48 585
R76 B.n503 B.n502 585
R77 B.n502 B.n44 585
R78 B.n501 B.n43 585
R79 B.n581 B.n43 585
R80 B.n500 B.n42 585
R81 B.n582 B.n42 585
R82 B.n499 B.n41 585
R83 B.n583 B.n41 585
R84 B.n498 B.n497 585
R85 B.n497 B.n37 585
R86 B.n496 B.n36 585
R87 B.n589 B.n36 585
R88 B.n495 B.n35 585
R89 B.n590 B.n35 585
R90 B.n494 B.n34 585
R91 B.n591 B.n34 585
R92 B.n493 B.n492 585
R93 B.n492 B.n30 585
R94 B.n491 B.n29 585
R95 B.n597 B.n29 585
R96 B.n490 B.n28 585
R97 B.n598 B.n28 585
R98 B.n489 B.n27 585
R99 B.n599 B.n27 585
R100 B.n488 B.n487 585
R101 B.n487 B.n23 585
R102 B.n486 B.n22 585
R103 B.n605 B.n22 585
R104 B.n485 B.n21 585
R105 B.n606 B.n21 585
R106 B.n484 B.n20 585
R107 B.n607 B.n20 585
R108 B.n483 B.n482 585
R109 B.n482 B.n16 585
R110 B.n481 B.n15 585
R111 B.n613 B.n15 585
R112 B.n480 B.n14 585
R113 B.n614 B.n14 585
R114 B.n479 B.n13 585
R115 B.n615 B.n13 585
R116 B.n478 B.n477 585
R117 B.n477 B.n12 585
R118 B.n476 B.n475 585
R119 B.n476 B.n8 585
R120 B.n474 B.n7 585
R121 B.n622 B.n7 585
R122 B.n473 B.n6 585
R123 B.n623 B.n6 585
R124 B.n472 B.n5 585
R125 B.n624 B.n5 585
R126 B.n471 B.n470 585
R127 B.n470 B.n4 585
R128 B.n469 B.n166 585
R129 B.n469 B.n468 585
R130 B.n459 B.n167 585
R131 B.n168 B.n167 585
R132 B.n461 B.n460 585
R133 B.n462 B.n461 585
R134 B.n458 B.n173 585
R135 B.n173 B.n172 585
R136 B.n457 B.n456 585
R137 B.n456 B.n455 585
R138 B.n175 B.n174 585
R139 B.n176 B.n175 585
R140 B.n448 B.n447 585
R141 B.n449 B.n448 585
R142 B.n446 B.n181 585
R143 B.n181 B.n180 585
R144 B.n445 B.n444 585
R145 B.n444 B.n443 585
R146 B.n183 B.n182 585
R147 B.n184 B.n183 585
R148 B.n436 B.n435 585
R149 B.n437 B.n436 585
R150 B.n434 B.n189 585
R151 B.n189 B.n188 585
R152 B.n433 B.n432 585
R153 B.n432 B.n431 585
R154 B.n191 B.n190 585
R155 B.n192 B.n191 585
R156 B.n424 B.n423 585
R157 B.n425 B.n424 585
R158 B.n422 B.n197 585
R159 B.n197 B.n196 585
R160 B.n421 B.n420 585
R161 B.n420 B.n419 585
R162 B.n199 B.n198 585
R163 B.n200 B.n199 585
R164 B.n412 B.n411 585
R165 B.n413 B.n412 585
R166 B.n410 B.n205 585
R167 B.n205 B.n204 585
R168 B.n409 B.n408 585
R169 B.n408 B.n407 585
R170 B.n207 B.n206 585
R171 B.n208 B.n207 585
R172 B.n400 B.n399 585
R173 B.n401 B.n400 585
R174 B.n398 B.n213 585
R175 B.n213 B.n212 585
R176 B.n397 B.n396 585
R177 B.n396 B.n395 585
R178 B.n215 B.n214 585
R179 B.n216 B.n215 585
R180 B.n388 B.n387 585
R181 B.n389 B.n388 585
R182 B.n386 B.n221 585
R183 B.n221 B.n220 585
R184 B.n385 B.n384 585
R185 B.n384 B.n383 585
R186 B.n223 B.n222 585
R187 B.n224 B.n223 585
R188 B.n376 B.n375 585
R189 B.n377 B.n376 585
R190 B.n374 B.n229 585
R191 B.n229 B.n228 585
R192 B.n373 B.n372 585
R193 B.n372 B.n371 585
R194 B.n231 B.n230 585
R195 B.n232 B.n231 585
R196 B.n364 B.n363 585
R197 B.n365 B.n364 585
R198 B.n362 B.n237 585
R199 B.n237 B.n236 585
R200 B.n361 B.n360 585
R201 B.n360 B.n359 585
R202 B.n239 B.n238 585
R203 B.n240 B.n239 585
R204 B.n352 B.n351 585
R205 B.n353 B.n352 585
R206 B.n350 B.n245 585
R207 B.n245 B.n244 585
R208 B.n349 B.n348 585
R209 B.n348 B.n347 585
R210 B.n247 B.n246 585
R211 B.n248 B.n247 585
R212 B.n340 B.n339 585
R213 B.n341 B.n340 585
R214 B.n338 B.n253 585
R215 B.n253 B.n252 585
R216 B.n332 B.n331 585
R217 B.n330 B.n270 585
R218 B.n329 B.n269 585
R219 B.n334 B.n269 585
R220 B.n328 B.n327 585
R221 B.n326 B.n325 585
R222 B.n324 B.n323 585
R223 B.n322 B.n321 585
R224 B.n320 B.n319 585
R225 B.n318 B.n317 585
R226 B.n316 B.n315 585
R227 B.n314 B.n313 585
R228 B.n312 B.n311 585
R229 B.n310 B.n309 585
R230 B.n308 B.n307 585
R231 B.n306 B.n305 585
R232 B.n304 B.n303 585
R233 B.n302 B.n301 585
R234 B.n300 B.n299 585
R235 B.n298 B.n297 585
R236 B.n296 B.n295 585
R237 B.n293 B.n292 585
R238 B.n291 B.n290 585
R239 B.n289 B.n288 585
R240 B.n287 B.n286 585
R241 B.n285 B.n284 585
R242 B.n283 B.n282 585
R243 B.n281 B.n280 585
R244 B.n279 B.n278 585
R245 B.n277 B.n276 585
R246 B.n255 B.n254 585
R247 B.n337 B.n336 585
R248 B.n251 B.n250 585
R249 B.n252 B.n251 585
R250 B.n343 B.n342 585
R251 B.n342 B.n341 585
R252 B.n344 B.n249 585
R253 B.n249 B.n248 585
R254 B.n346 B.n345 585
R255 B.n347 B.n346 585
R256 B.n243 B.n242 585
R257 B.n244 B.n243 585
R258 B.n355 B.n354 585
R259 B.n354 B.n353 585
R260 B.n356 B.n241 585
R261 B.n241 B.n240 585
R262 B.n358 B.n357 585
R263 B.n359 B.n358 585
R264 B.n235 B.n234 585
R265 B.n236 B.n235 585
R266 B.n367 B.n366 585
R267 B.n366 B.n365 585
R268 B.n368 B.n233 585
R269 B.n233 B.n232 585
R270 B.n370 B.n369 585
R271 B.n371 B.n370 585
R272 B.n227 B.n226 585
R273 B.n228 B.n227 585
R274 B.n379 B.n378 585
R275 B.n378 B.n377 585
R276 B.n380 B.n225 585
R277 B.n225 B.n224 585
R278 B.n382 B.n381 585
R279 B.n383 B.n382 585
R280 B.n219 B.n218 585
R281 B.n220 B.n219 585
R282 B.n391 B.n390 585
R283 B.n390 B.n389 585
R284 B.n392 B.n217 585
R285 B.n217 B.n216 585
R286 B.n394 B.n393 585
R287 B.n395 B.n394 585
R288 B.n211 B.n210 585
R289 B.n212 B.n211 585
R290 B.n403 B.n402 585
R291 B.n402 B.n401 585
R292 B.n404 B.n209 585
R293 B.n209 B.n208 585
R294 B.n406 B.n405 585
R295 B.n407 B.n406 585
R296 B.n203 B.n202 585
R297 B.n204 B.n203 585
R298 B.n415 B.n414 585
R299 B.n414 B.n413 585
R300 B.n416 B.n201 585
R301 B.n201 B.n200 585
R302 B.n418 B.n417 585
R303 B.n419 B.n418 585
R304 B.n195 B.n194 585
R305 B.n196 B.n195 585
R306 B.n427 B.n426 585
R307 B.n426 B.n425 585
R308 B.n428 B.n193 585
R309 B.n193 B.n192 585
R310 B.n430 B.n429 585
R311 B.n431 B.n430 585
R312 B.n187 B.n186 585
R313 B.n188 B.n187 585
R314 B.n439 B.n438 585
R315 B.n438 B.n437 585
R316 B.n440 B.n185 585
R317 B.n185 B.n184 585
R318 B.n442 B.n441 585
R319 B.n443 B.n442 585
R320 B.n179 B.n178 585
R321 B.n180 B.n179 585
R322 B.n451 B.n450 585
R323 B.n450 B.n449 585
R324 B.n452 B.n177 585
R325 B.n177 B.n176 585
R326 B.n454 B.n453 585
R327 B.n455 B.n454 585
R328 B.n171 B.n170 585
R329 B.n172 B.n171 585
R330 B.n464 B.n463 585
R331 B.n463 B.n462 585
R332 B.n465 B.n169 585
R333 B.n169 B.n168 585
R334 B.n467 B.n466 585
R335 B.n468 B.n467 585
R336 B.n3 B.n0 585
R337 B.n4 B.n3 585
R338 B.n621 B.n1 585
R339 B.n622 B.n621 585
R340 B.n620 B.n619 585
R341 B.n620 B.n8 585
R342 B.n618 B.n9 585
R343 B.n12 B.n9 585
R344 B.n617 B.n616 585
R345 B.n616 B.n615 585
R346 B.n11 B.n10 585
R347 B.n614 B.n11 585
R348 B.n612 B.n611 585
R349 B.n613 B.n612 585
R350 B.n610 B.n17 585
R351 B.n17 B.n16 585
R352 B.n609 B.n608 585
R353 B.n608 B.n607 585
R354 B.n19 B.n18 585
R355 B.n606 B.n19 585
R356 B.n604 B.n603 585
R357 B.n605 B.n604 585
R358 B.n602 B.n24 585
R359 B.n24 B.n23 585
R360 B.n601 B.n600 585
R361 B.n600 B.n599 585
R362 B.n26 B.n25 585
R363 B.n598 B.n26 585
R364 B.n596 B.n595 585
R365 B.n597 B.n596 585
R366 B.n594 B.n31 585
R367 B.n31 B.n30 585
R368 B.n593 B.n592 585
R369 B.n592 B.n591 585
R370 B.n33 B.n32 585
R371 B.n590 B.n33 585
R372 B.n588 B.n587 585
R373 B.n589 B.n588 585
R374 B.n586 B.n38 585
R375 B.n38 B.n37 585
R376 B.n585 B.n584 585
R377 B.n584 B.n583 585
R378 B.n40 B.n39 585
R379 B.n582 B.n40 585
R380 B.n580 B.n579 585
R381 B.n581 B.n580 585
R382 B.n578 B.n45 585
R383 B.n45 B.n44 585
R384 B.n577 B.n576 585
R385 B.n576 B.n575 585
R386 B.n47 B.n46 585
R387 B.n574 B.n47 585
R388 B.n572 B.n571 585
R389 B.n573 B.n572 585
R390 B.n570 B.n52 585
R391 B.n52 B.n51 585
R392 B.n569 B.n568 585
R393 B.n568 B.n567 585
R394 B.n54 B.n53 585
R395 B.n566 B.n54 585
R396 B.n564 B.n563 585
R397 B.n565 B.n564 585
R398 B.n562 B.n59 585
R399 B.n59 B.n58 585
R400 B.n561 B.n560 585
R401 B.n560 B.n559 585
R402 B.n61 B.n60 585
R403 B.n558 B.n61 585
R404 B.n556 B.n555 585
R405 B.n557 B.n556 585
R406 B.n554 B.n66 585
R407 B.n66 B.n65 585
R408 B.n553 B.n552 585
R409 B.n552 B.n551 585
R410 B.n68 B.n67 585
R411 B.n550 B.n68 585
R412 B.n548 B.n547 585
R413 B.n549 B.n548 585
R414 B.n546 B.n73 585
R415 B.n73 B.n72 585
R416 B.n545 B.n544 585
R417 B.n544 B.n543 585
R418 B.n75 B.n74 585
R419 B.n542 B.n75 585
R420 B.n540 B.n539 585
R421 B.n541 B.n540 585
R422 B.n538 B.n80 585
R423 B.n80 B.n79 585
R424 B.n537 B.n536 585
R425 B.n536 B.n535 585
R426 B.n82 B.n81 585
R427 B.n534 B.n82 585
R428 B.n625 B.n624 585
R429 B.n623 B.n2 585
R430 B.n106 B.n82 449.257
R431 B.n532 B.n84 449.257
R432 B.n336 B.n253 449.257
R433 B.n332 B.n251 449.257
R434 B.n533 B.n99 256.663
R435 B.n533 B.n98 256.663
R436 B.n533 B.n97 256.663
R437 B.n533 B.n96 256.663
R438 B.n533 B.n95 256.663
R439 B.n533 B.n94 256.663
R440 B.n533 B.n93 256.663
R441 B.n533 B.n92 256.663
R442 B.n533 B.n91 256.663
R443 B.n533 B.n90 256.663
R444 B.n533 B.n89 256.663
R445 B.n533 B.n88 256.663
R446 B.n533 B.n87 256.663
R447 B.n533 B.n86 256.663
R448 B.n533 B.n85 256.663
R449 B.n334 B.n333 256.663
R450 B.n334 B.n256 256.663
R451 B.n334 B.n257 256.663
R452 B.n334 B.n258 256.663
R453 B.n334 B.n259 256.663
R454 B.n334 B.n260 256.663
R455 B.n334 B.n261 256.663
R456 B.n334 B.n262 256.663
R457 B.n334 B.n263 256.663
R458 B.n334 B.n264 256.663
R459 B.n334 B.n265 256.663
R460 B.n334 B.n266 256.663
R461 B.n334 B.n267 256.663
R462 B.n334 B.n268 256.663
R463 B.n335 B.n334 256.663
R464 B.n627 B.n626 256.663
R465 B.n104 B.t12 209.876
R466 B.n101 B.t8 209.876
R467 B.n274 B.t15 209.876
R468 B.n271 B.t4 209.876
R469 B.n101 B.t10 188.569
R470 B.n274 B.t17 188.569
R471 B.n104 B.t13 188.567
R472 B.n271 B.t7 188.567
R473 B.n334 B.n252 185.108
R474 B.n534 B.n533 185.108
R475 B.n110 B.n109 163.367
R476 B.n114 B.n113 163.367
R477 B.n118 B.n117 163.367
R478 B.n122 B.n121 163.367
R479 B.n126 B.n125 163.367
R480 B.n131 B.n130 163.367
R481 B.n135 B.n134 163.367
R482 B.n139 B.n138 163.367
R483 B.n143 B.n142 163.367
R484 B.n147 B.n146 163.367
R485 B.n151 B.n150 163.367
R486 B.n155 B.n154 163.367
R487 B.n159 B.n158 163.367
R488 B.n163 B.n162 163.367
R489 B.n532 B.n100 163.367
R490 B.n340 B.n253 163.367
R491 B.n340 B.n247 163.367
R492 B.n348 B.n247 163.367
R493 B.n348 B.n245 163.367
R494 B.n352 B.n245 163.367
R495 B.n352 B.n239 163.367
R496 B.n360 B.n239 163.367
R497 B.n360 B.n237 163.367
R498 B.n364 B.n237 163.367
R499 B.n364 B.n231 163.367
R500 B.n372 B.n231 163.367
R501 B.n372 B.n229 163.367
R502 B.n376 B.n229 163.367
R503 B.n376 B.n223 163.367
R504 B.n384 B.n223 163.367
R505 B.n384 B.n221 163.367
R506 B.n388 B.n221 163.367
R507 B.n388 B.n215 163.367
R508 B.n396 B.n215 163.367
R509 B.n396 B.n213 163.367
R510 B.n400 B.n213 163.367
R511 B.n400 B.n207 163.367
R512 B.n408 B.n207 163.367
R513 B.n408 B.n205 163.367
R514 B.n412 B.n205 163.367
R515 B.n412 B.n199 163.367
R516 B.n420 B.n199 163.367
R517 B.n420 B.n197 163.367
R518 B.n424 B.n197 163.367
R519 B.n424 B.n191 163.367
R520 B.n432 B.n191 163.367
R521 B.n432 B.n189 163.367
R522 B.n436 B.n189 163.367
R523 B.n436 B.n183 163.367
R524 B.n444 B.n183 163.367
R525 B.n444 B.n181 163.367
R526 B.n448 B.n181 163.367
R527 B.n448 B.n175 163.367
R528 B.n456 B.n175 163.367
R529 B.n456 B.n173 163.367
R530 B.n461 B.n173 163.367
R531 B.n461 B.n167 163.367
R532 B.n469 B.n167 163.367
R533 B.n470 B.n469 163.367
R534 B.n470 B.n5 163.367
R535 B.n6 B.n5 163.367
R536 B.n7 B.n6 163.367
R537 B.n476 B.n7 163.367
R538 B.n477 B.n476 163.367
R539 B.n477 B.n13 163.367
R540 B.n14 B.n13 163.367
R541 B.n15 B.n14 163.367
R542 B.n482 B.n15 163.367
R543 B.n482 B.n20 163.367
R544 B.n21 B.n20 163.367
R545 B.n22 B.n21 163.367
R546 B.n487 B.n22 163.367
R547 B.n487 B.n27 163.367
R548 B.n28 B.n27 163.367
R549 B.n29 B.n28 163.367
R550 B.n492 B.n29 163.367
R551 B.n492 B.n34 163.367
R552 B.n35 B.n34 163.367
R553 B.n36 B.n35 163.367
R554 B.n497 B.n36 163.367
R555 B.n497 B.n41 163.367
R556 B.n42 B.n41 163.367
R557 B.n43 B.n42 163.367
R558 B.n502 B.n43 163.367
R559 B.n502 B.n48 163.367
R560 B.n49 B.n48 163.367
R561 B.n50 B.n49 163.367
R562 B.n507 B.n50 163.367
R563 B.n507 B.n55 163.367
R564 B.n56 B.n55 163.367
R565 B.n57 B.n56 163.367
R566 B.n512 B.n57 163.367
R567 B.n512 B.n62 163.367
R568 B.n63 B.n62 163.367
R569 B.n64 B.n63 163.367
R570 B.n517 B.n64 163.367
R571 B.n517 B.n69 163.367
R572 B.n70 B.n69 163.367
R573 B.n71 B.n70 163.367
R574 B.n522 B.n71 163.367
R575 B.n522 B.n76 163.367
R576 B.n77 B.n76 163.367
R577 B.n78 B.n77 163.367
R578 B.n527 B.n78 163.367
R579 B.n527 B.n83 163.367
R580 B.n84 B.n83 163.367
R581 B.n270 B.n269 163.367
R582 B.n327 B.n269 163.367
R583 B.n325 B.n324 163.367
R584 B.n321 B.n320 163.367
R585 B.n317 B.n316 163.367
R586 B.n313 B.n312 163.367
R587 B.n309 B.n308 163.367
R588 B.n305 B.n304 163.367
R589 B.n301 B.n300 163.367
R590 B.n297 B.n296 163.367
R591 B.n292 B.n291 163.367
R592 B.n288 B.n287 163.367
R593 B.n284 B.n283 163.367
R594 B.n280 B.n279 163.367
R595 B.n276 B.n255 163.367
R596 B.n342 B.n251 163.367
R597 B.n342 B.n249 163.367
R598 B.n346 B.n249 163.367
R599 B.n346 B.n243 163.367
R600 B.n354 B.n243 163.367
R601 B.n354 B.n241 163.367
R602 B.n358 B.n241 163.367
R603 B.n358 B.n235 163.367
R604 B.n366 B.n235 163.367
R605 B.n366 B.n233 163.367
R606 B.n370 B.n233 163.367
R607 B.n370 B.n227 163.367
R608 B.n378 B.n227 163.367
R609 B.n378 B.n225 163.367
R610 B.n382 B.n225 163.367
R611 B.n382 B.n219 163.367
R612 B.n390 B.n219 163.367
R613 B.n390 B.n217 163.367
R614 B.n394 B.n217 163.367
R615 B.n394 B.n211 163.367
R616 B.n402 B.n211 163.367
R617 B.n402 B.n209 163.367
R618 B.n406 B.n209 163.367
R619 B.n406 B.n203 163.367
R620 B.n414 B.n203 163.367
R621 B.n414 B.n201 163.367
R622 B.n418 B.n201 163.367
R623 B.n418 B.n195 163.367
R624 B.n426 B.n195 163.367
R625 B.n426 B.n193 163.367
R626 B.n430 B.n193 163.367
R627 B.n430 B.n187 163.367
R628 B.n438 B.n187 163.367
R629 B.n438 B.n185 163.367
R630 B.n442 B.n185 163.367
R631 B.n442 B.n179 163.367
R632 B.n450 B.n179 163.367
R633 B.n450 B.n177 163.367
R634 B.n454 B.n177 163.367
R635 B.n454 B.n171 163.367
R636 B.n463 B.n171 163.367
R637 B.n463 B.n169 163.367
R638 B.n467 B.n169 163.367
R639 B.n467 B.n3 163.367
R640 B.n625 B.n3 163.367
R641 B.n621 B.n2 163.367
R642 B.n621 B.n620 163.367
R643 B.n620 B.n9 163.367
R644 B.n616 B.n9 163.367
R645 B.n616 B.n11 163.367
R646 B.n612 B.n11 163.367
R647 B.n612 B.n17 163.367
R648 B.n608 B.n17 163.367
R649 B.n608 B.n19 163.367
R650 B.n604 B.n19 163.367
R651 B.n604 B.n24 163.367
R652 B.n600 B.n24 163.367
R653 B.n600 B.n26 163.367
R654 B.n596 B.n26 163.367
R655 B.n596 B.n31 163.367
R656 B.n592 B.n31 163.367
R657 B.n592 B.n33 163.367
R658 B.n588 B.n33 163.367
R659 B.n588 B.n38 163.367
R660 B.n584 B.n38 163.367
R661 B.n584 B.n40 163.367
R662 B.n580 B.n40 163.367
R663 B.n580 B.n45 163.367
R664 B.n576 B.n45 163.367
R665 B.n576 B.n47 163.367
R666 B.n572 B.n47 163.367
R667 B.n572 B.n52 163.367
R668 B.n568 B.n52 163.367
R669 B.n568 B.n54 163.367
R670 B.n564 B.n54 163.367
R671 B.n564 B.n59 163.367
R672 B.n560 B.n59 163.367
R673 B.n560 B.n61 163.367
R674 B.n556 B.n61 163.367
R675 B.n556 B.n66 163.367
R676 B.n552 B.n66 163.367
R677 B.n552 B.n68 163.367
R678 B.n548 B.n68 163.367
R679 B.n548 B.n73 163.367
R680 B.n544 B.n73 163.367
R681 B.n544 B.n75 163.367
R682 B.n540 B.n75 163.367
R683 B.n540 B.n80 163.367
R684 B.n536 B.n80 163.367
R685 B.n536 B.n82 163.367
R686 B.n341 B.n252 111.392
R687 B.n341 B.n248 111.392
R688 B.n347 B.n248 111.392
R689 B.n347 B.n244 111.392
R690 B.n353 B.n244 111.392
R691 B.n353 B.n240 111.392
R692 B.n359 B.n240 111.392
R693 B.n359 B.n236 111.392
R694 B.n365 B.n236 111.392
R695 B.n371 B.n232 111.392
R696 B.n371 B.n228 111.392
R697 B.n377 B.n228 111.392
R698 B.n377 B.n224 111.392
R699 B.n383 B.n224 111.392
R700 B.n383 B.n220 111.392
R701 B.n389 B.n220 111.392
R702 B.n389 B.n216 111.392
R703 B.n395 B.n216 111.392
R704 B.n395 B.n212 111.392
R705 B.n401 B.n212 111.392
R706 B.n401 B.n208 111.392
R707 B.n407 B.n208 111.392
R708 B.n407 B.n204 111.392
R709 B.n413 B.n204 111.392
R710 B.n419 B.n200 111.392
R711 B.n419 B.n196 111.392
R712 B.n425 B.n196 111.392
R713 B.n425 B.n192 111.392
R714 B.n431 B.n192 111.392
R715 B.n431 B.n188 111.392
R716 B.n437 B.n188 111.392
R717 B.n437 B.n184 111.392
R718 B.n443 B.n184 111.392
R719 B.n443 B.n180 111.392
R720 B.n449 B.n180 111.392
R721 B.n455 B.n176 111.392
R722 B.n455 B.n172 111.392
R723 B.n462 B.n172 111.392
R724 B.n462 B.n168 111.392
R725 B.n468 B.n168 111.392
R726 B.n468 B.n4 111.392
R727 B.n624 B.n4 111.392
R728 B.n624 B.n623 111.392
R729 B.n623 B.n622 111.392
R730 B.n622 B.n8 111.392
R731 B.n12 B.n8 111.392
R732 B.n615 B.n12 111.392
R733 B.n615 B.n614 111.392
R734 B.n614 B.n613 111.392
R735 B.n613 B.n16 111.392
R736 B.n607 B.n606 111.392
R737 B.n606 B.n605 111.392
R738 B.n605 B.n23 111.392
R739 B.n599 B.n23 111.392
R740 B.n599 B.n598 111.392
R741 B.n598 B.n597 111.392
R742 B.n597 B.n30 111.392
R743 B.n591 B.n30 111.392
R744 B.n591 B.n590 111.392
R745 B.n590 B.n589 111.392
R746 B.n589 B.n37 111.392
R747 B.n583 B.n582 111.392
R748 B.n582 B.n581 111.392
R749 B.n581 B.n44 111.392
R750 B.n575 B.n44 111.392
R751 B.n575 B.n574 111.392
R752 B.n574 B.n573 111.392
R753 B.n573 B.n51 111.392
R754 B.n567 B.n51 111.392
R755 B.n567 B.n566 111.392
R756 B.n566 B.n565 111.392
R757 B.n565 B.n58 111.392
R758 B.n559 B.n58 111.392
R759 B.n559 B.n558 111.392
R760 B.n558 B.n557 111.392
R761 B.n557 B.n65 111.392
R762 B.n551 B.n550 111.392
R763 B.n550 B.n549 111.392
R764 B.n549 B.n72 111.392
R765 B.n543 B.n72 111.392
R766 B.n543 B.n542 111.392
R767 B.n542 B.n541 111.392
R768 B.n541 B.n79 111.392
R769 B.n535 B.n79 111.392
R770 B.n535 B.n534 111.392
R771 B.n102 B.t11 106.725
R772 B.n275 B.t16 106.725
R773 B.n105 B.t14 106.725
R774 B.n272 B.t6 106.725
R775 B.n105 B.n104 81.8429
R776 B.n102 B.n101 81.8429
R777 B.n275 B.n274 81.8429
R778 B.n272 B.n271 81.8429
R779 B.t1 B.n200 80.2686
R780 B.t3 B.n37 80.2686
R781 B.n449 B.t0 76.9923
R782 B.n607 B.t2 76.9923
R783 B.n365 B.t5 73.7161
R784 B.n551 B.t9 73.7161
R785 B.n106 B.n85 71.676
R786 B.n110 B.n86 71.676
R787 B.n114 B.n87 71.676
R788 B.n118 B.n88 71.676
R789 B.n122 B.n89 71.676
R790 B.n126 B.n90 71.676
R791 B.n131 B.n91 71.676
R792 B.n135 B.n92 71.676
R793 B.n139 B.n93 71.676
R794 B.n143 B.n94 71.676
R795 B.n147 B.n95 71.676
R796 B.n151 B.n96 71.676
R797 B.n155 B.n97 71.676
R798 B.n159 B.n98 71.676
R799 B.n163 B.n99 71.676
R800 B.n100 B.n99 71.676
R801 B.n162 B.n98 71.676
R802 B.n158 B.n97 71.676
R803 B.n154 B.n96 71.676
R804 B.n150 B.n95 71.676
R805 B.n146 B.n94 71.676
R806 B.n142 B.n93 71.676
R807 B.n138 B.n92 71.676
R808 B.n134 B.n91 71.676
R809 B.n130 B.n90 71.676
R810 B.n125 B.n89 71.676
R811 B.n121 B.n88 71.676
R812 B.n117 B.n87 71.676
R813 B.n113 B.n86 71.676
R814 B.n109 B.n85 71.676
R815 B.n333 B.n332 71.676
R816 B.n327 B.n256 71.676
R817 B.n324 B.n257 71.676
R818 B.n320 B.n258 71.676
R819 B.n316 B.n259 71.676
R820 B.n312 B.n260 71.676
R821 B.n308 B.n261 71.676
R822 B.n304 B.n262 71.676
R823 B.n300 B.n263 71.676
R824 B.n296 B.n264 71.676
R825 B.n291 B.n265 71.676
R826 B.n287 B.n266 71.676
R827 B.n283 B.n267 71.676
R828 B.n279 B.n268 71.676
R829 B.n335 B.n255 71.676
R830 B.n333 B.n270 71.676
R831 B.n325 B.n256 71.676
R832 B.n321 B.n257 71.676
R833 B.n317 B.n258 71.676
R834 B.n313 B.n259 71.676
R835 B.n309 B.n260 71.676
R836 B.n305 B.n261 71.676
R837 B.n301 B.n262 71.676
R838 B.n297 B.n263 71.676
R839 B.n292 B.n264 71.676
R840 B.n288 B.n265 71.676
R841 B.n284 B.n266 71.676
R842 B.n280 B.n267 71.676
R843 B.n276 B.n268 71.676
R844 B.n336 B.n335 71.676
R845 B.n626 B.n625 71.676
R846 B.n626 B.n2 71.676
R847 B.n128 B.n105 59.5399
R848 B.n103 B.n102 59.5399
R849 B.n294 B.n275 59.5399
R850 B.n273 B.n272 59.5399
R851 B.t5 B.n232 37.6773
R852 B.t9 B.n65 37.6773
R853 B.t0 B.n176 34.4011
R854 B.t2 B.n16 34.4011
R855 B.n413 B.t1 31.1248
R856 B.n583 B.t3 31.1248
R857 B.n331 B.n250 29.1907
R858 B.n338 B.n337 29.1907
R859 B.n531 B.n530 29.1907
R860 B.n107 B.n81 29.1907
R861 B B.n627 18.0485
R862 B.n343 B.n250 10.6151
R863 B.n344 B.n343 10.6151
R864 B.n345 B.n344 10.6151
R865 B.n345 B.n242 10.6151
R866 B.n355 B.n242 10.6151
R867 B.n356 B.n355 10.6151
R868 B.n357 B.n356 10.6151
R869 B.n357 B.n234 10.6151
R870 B.n367 B.n234 10.6151
R871 B.n368 B.n367 10.6151
R872 B.n369 B.n368 10.6151
R873 B.n369 B.n226 10.6151
R874 B.n379 B.n226 10.6151
R875 B.n380 B.n379 10.6151
R876 B.n381 B.n380 10.6151
R877 B.n381 B.n218 10.6151
R878 B.n391 B.n218 10.6151
R879 B.n392 B.n391 10.6151
R880 B.n393 B.n392 10.6151
R881 B.n393 B.n210 10.6151
R882 B.n403 B.n210 10.6151
R883 B.n404 B.n403 10.6151
R884 B.n405 B.n404 10.6151
R885 B.n405 B.n202 10.6151
R886 B.n415 B.n202 10.6151
R887 B.n416 B.n415 10.6151
R888 B.n417 B.n416 10.6151
R889 B.n417 B.n194 10.6151
R890 B.n427 B.n194 10.6151
R891 B.n428 B.n427 10.6151
R892 B.n429 B.n428 10.6151
R893 B.n429 B.n186 10.6151
R894 B.n439 B.n186 10.6151
R895 B.n440 B.n439 10.6151
R896 B.n441 B.n440 10.6151
R897 B.n441 B.n178 10.6151
R898 B.n451 B.n178 10.6151
R899 B.n452 B.n451 10.6151
R900 B.n453 B.n452 10.6151
R901 B.n453 B.n170 10.6151
R902 B.n464 B.n170 10.6151
R903 B.n465 B.n464 10.6151
R904 B.n466 B.n465 10.6151
R905 B.n466 B.n0 10.6151
R906 B.n331 B.n330 10.6151
R907 B.n330 B.n329 10.6151
R908 B.n329 B.n328 10.6151
R909 B.n328 B.n326 10.6151
R910 B.n326 B.n323 10.6151
R911 B.n323 B.n322 10.6151
R912 B.n322 B.n319 10.6151
R913 B.n319 B.n318 10.6151
R914 B.n318 B.n315 10.6151
R915 B.n315 B.n314 10.6151
R916 B.n311 B.n310 10.6151
R917 B.n310 B.n307 10.6151
R918 B.n307 B.n306 10.6151
R919 B.n306 B.n303 10.6151
R920 B.n303 B.n302 10.6151
R921 B.n302 B.n299 10.6151
R922 B.n299 B.n298 10.6151
R923 B.n298 B.n295 10.6151
R924 B.n293 B.n290 10.6151
R925 B.n290 B.n289 10.6151
R926 B.n289 B.n286 10.6151
R927 B.n286 B.n285 10.6151
R928 B.n285 B.n282 10.6151
R929 B.n282 B.n281 10.6151
R930 B.n281 B.n278 10.6151
R931 B.n278 B.n277 10.6151
R932 B.n277 B.n254 10.6151
R933 B.n337 B.n254 10.6151
R934 B.n339 B.n338 10.6151
R935 B.n339 B.n246 10.6151
R936 B.n349 B.n246 10.6151
R937 B.n350 B.n349 10.6151
R938 B.n351 B.n350 10.6151
R939 B.n351 B.n238 10.6151
R940 B.n361 B.n238 10.6151
R941 B.n362 B.n361 10.6151
R942 B.n363 B.n362 10.6151
R943 B.n363 B.n230 10.6151
R944 B.n373 B.n230 10.6151
R945 B.n374 B.n373 10.6151
R946 B.n375 B.n374 10.6151
R947 B.n375 B.n222 10.6151
R948 B.n385 B.n222 10.6151
R949 B.n386 B.n385 10.6151
R950 B.n387 B.n386 10.6151
R951 B.n387 B.n214 10.6151
R952 B.n397 B.n214 10.6151
R953 B.n398 B.n397 10.6151
R954 B.n399 B.n398 10.6151
R955 B.n399 B.n206 10.6151
R956 B.n409 B.n206 10.6151
R957 B.n410 B.n409 10.6151
R958 B.n411 B.n410 10.6151
R959 B.n411 B.n198 10.6151
R960 B.n421 B.n198 10.6151
R961 B.n422 B.n421 10.6151
R962 B.n423 B.n422 10.6151
R963 B.n423 B.n190 10.6151
R964 B.n433 B.n190 10.6151
R965 B.n434 B.n433 10.6151
R966 B.n435 B.n434 10.6151
R967 B.n435 B.n182 10.6151
R968 B.n445 B.n182 10.6151
R969 B.n446 B.n445 10.6151
R970 B.n447 B.n446 10.6151
R971 B.n447 B.n174 10.6151
R972 B.n457 B.n174 10.6151
R973 B.n458 B.n457 10.6151
R974 B.n460 B.n458 10.6151
R975 B.n460 B.n459 10.6151
R976 B.n459 B.n166 10.6151
R977 B.n471 B.n166 10.6151
R978 B.n472 B.n471 10.6151
R979 B.n473 B.n472 10.6151
R980 B.n474 B.n473 10.6151
R981 B.n475 B.n474 10.6151
R982 B.n478 B.n475 10.6151
R983 B.n479 B.n478 10.6151
R984 B.n480 B.n479 10.6151
R985 B.n481 B.n480 10.6151
R986 B.n483 B.n481 10.6151
R987 B.n484 B.n483 10.6151
R988 B.n485 B.n484 10.6151
R989 B.n486 B.n485 10.6151
R990 B.n488 B.n486 10.6151
R991 B.n489 B.n488 10.6151
R992 B.n490 B.n489 10.6151
R993 B.n491 B.n490 10.6151
R994 B.n493 B.n491 10.6151
R995 B.n494 B.n493 10.6151
R996 B.n495 B.n494 10.6151
R997 B.n496 B.n495 10.6151
R998 B.n498 B.n496 10.6151
R999 B.n499 B.n498 10.6151
R1000 B.n500 B.n499 10.6151
R1001 B.n501 B.n500 10.6151
R1002 B.n503 B.n501 10.6151
R1003 B.n504 B.n503 10.6151
R1004 B.n505 B.n504 10.6151
R1005 B.n506 B.n505 10.6151
R1006 B.n508 B.n506 10.6151
R1007 B.n509 B.n508 10.6151
R1008 B.n510 B.n509 10.6151
R1009 B.n511 B.n510 10.6151
R1010 B.n513 B.n511 10.6151
R1011 B.n514 B.n513 10.6151
R1012 B.n515 B.n514 10.6151
R1013 B.n516 B.n515 10.6151
R1014 B.n518 B.n516 10.6151
R1015 B.n519 B.n518 10.6151
R1016 B.n520 B.n519 10.6151
R1017 B.n521 B.n520 10.6151
R1018 B.n523 B.n521 10.6151
R1019 B.n524 B.n523 10.6151
R1020 B.n525 B.n524 10.6151
R1021 B.n526 B.n525 10.6151
R1022 B.n528 B.n526 10.6151
R1023 B.n529 B.n528 10.6151
R1024 B.n530 B.n529 10.6151
R1025 B.n619 B.n1 10.6151
R1026 B.n619 B.n618 10.6151
R1027 B.n618 B.n617 10.6151
R1028 B.n617 B.n10 10.6151
R1029 B.n611 B.n10 10.6151
R1030 B.n611 B.n610 10.6151
R1031 B.n610 B.n609 10.6151
R1032 B.n609 B.n18 10.6151
R1033 B.n603 B.n18 10.6151
R1034 B.n603 B.n602 10.6151
R1035 B.n602 B.n601 10.6151
R1036 B.n601 B.n25 10.6151
R1037 B.n595 B.n25 10.6151
R1038 B.n595 B.n594 10.6151
R1039 B.n594 B.n593 10.6151
R1040 B.n593 B.n32 10.6151
R1041 B.n587 B.n32 10.6151
R1042 B.n587 B.n586 10.6151
R1043 B.n586 B.n585 10.6151
R1044 B.n585 B.n39 10.6151
R1045 B.n579 B.n39 10.6151
R1046 B.n579 B.n578 10.6151
R1047 B.n578 B.n577 10.6151
R1048 B.n577 B.n46 10.6151
R1049 B.n571 B.n46 10.6151
R1050 B.n571 B.n570 10.6151
R1051 B.n570 B.n569 10.6151
R1052 B.n569 B.n53 10.6151
R1053 B.n563 B.n53 10.6151
R1054 B.n563 B.n562 10.6151
R1055 B.n562 B.n561 10.6151
R1056 B.n561 B.n60 10.6151
R1057 B.n555 B.n60 10.6151
R1058 B.n555 B.n554 10.6151
R1059 B.n554 B.n553 10.6151
R1060 B.n553 B.n67 10.6151
R1061 B.n547 B.n67 10.6151
R1062 B.n547 B.n546 10.6151
R1063 B.n546 B.n545 10.6151
R1064 B.n545 B.n74 10.6151
R1065 B.n539 B.n74 10.6151
R1066 B.n539 B.n538 10.6151
R1067 B.n538 B.n537 10.6151
R1068 B.n537 B.n81 10.6151
R1069 B.n108 B.n107 10.6151
R1070 B.n111 B.n108 10.6151
R1071 B.n112 B.n111 10.6151
R1072 B.n115 B.n112 10.6151
R1073 B.n116 B.n115 10.6151
R1074 B.n119 B.n116 10.6151
R1075 B.n120 B.n119 10.6151
R1076 B.n123 B.n120 10.6151
R1077 B.n124 B.n123 10.6151
R1078 B.n127 B.n124 10.6151
R1079 B.n132 B.n129 10.6151
R1080 B.n133 B.n132 10.6151
R1081 B.n136 B.n133 10.6151
R1082 B.n137 B.n136 10.6151
R1083 B.n140 B.n137 10.6151
R1084 B.n141 B.n140 10.6151
R1085 B.n144 B.n141 10.6151
R1086 B.n145 B.n144 10.6151
R1087 B.n149 B.n148 10.6151
R1088 B.n152 B.n149 10.6151
R1089 B.n153 B.n152 10.6151
R1090 B.n156 B.n153 10.6151
R1091 B.n157 B.n156 10.6151
R1092 B.n160 B.n157 10.6151
R1093 B.n161 B.n160 10.6151
R1094 B.n164 B.n161 10.6151
R1095 B.n165 B.n164 10.6151
R1096 B.n531 B.n165 10.6151
R1097 B.n627 B.n0 8.11757
R1098 B.n627 B.n1 8.11757
R1099 B.n311 B.n273 6.5566
R1100 B.n295 B.n294 6.5566
R1101 B.n129 B.n128 6.5566
R1102 B.n145 B.n103 6.5566
R1103 B.n314 B.n273 4.05904
R1104 B.n294 B.n293 4.05904
R1105 B.n128 B.n127 4.05904
R1106 B.n148 B.n103 4.05904
R1107 VN VN.n1 44.3315
R1108 VN.n1 VN.t1 43.4664
R1109 VN.n0 VN.t3 43.4664
R1110 VN.n0 VN.t0 42.0932
R1111 VN.n1 VN.t2 42.0932
R1112 VN VN.n0 1.78227
R1113 VTAIL.n5 VTAIL.t1 113.472
R1114 VTAIL.n4 VTAIL.t6 113.472
R1115 VTAIL.n3 VTAIL.t5 113.472
R1116 VTAIL.n7 VTAIL.t7 113.472
R1117 VTAIL.n0 VTAIL.t4 113.472
R1118 VTAIL.n1 VTAIL.t0 113.472
R1119 VTAIL.n2 VTAIL.t3 113.472
R1120 VTAIL.n6 VTAIL.t2 113.472
R1121 VTAIL.n7 VTAIL.n6 17.2462
R1122 VTAIL.n3 VTAIL.n2 17.2462
R1123 VTAIL.n4 VTAIL.n3 3.63843
R1124 VTAIL.n6 VTAIL.n5 3.63843
R1125 VTAIL.n2 VTAIL.n1 3.63843
R1126 VTAIL VTAIL.n0 1.87766
R1127 VTAIL VTAIL.n7 1.76128
R1128 VTAIL.n5 VTAIL.n4 0.470328
R1129 VTAIL.n1 VTAIL.n0 0.470328
R1130 VDD2.n2 VDD2.n0 152.27
R1131 VDD2.n2 VDD2.n1 116.4
R1132 VDD2.n1 VDD2.t1 13.7505
R1133 VDD2.n1 VDD2.t2 13.7505
R1134 VDD2.n0 VDD2.t0 13.7505
R1135 VDD2.n0 VDD2.t3 13.7505
R1136 VDD2 VDD2.n2 0.0586897
R1137 VP.n21 VP.n20 161.3
R1138 VP.n19 VP.n1 161.3
R1139 VP.n18 VP.n17 161.3
R1140 VP.n16 VP.n2 161.3
R1141 VP.n15 VP.n14 161.3
R1142 VP.n13 VP.n3 161.3
R1143 VP.n12 VP.n11 161.3
R1144 VP.n10 VP.n4 161.3
R1145 VP.n9 VP.n8 161.3
R1146 VP.n7 VP.n6 84.8354
R1147 VP.n22 VP.n0 84.8354
R1148 VP.n6 VP.n5 44.1663
R1149 VP.n5 VP.t0 43.4663
R1150 VP.n5 VP.t1 42.0932
R1151 VP.n14 VP.n13 40.577
R1152 VP.n14 VP.n2 40.577
R1153 VP.n8 VP.n4 24.5923
R1154 VP.n12 VP.n4 24.5923
R1155 VP.n13 VP.n12 24.5923
R1156 VP.n18 VP.n2 24.5923
R1157 VP.n19 VP.n18 24.5923
R1158 VP.n20 VP.n19 24.5923
R1159 VP.n7 VP.t2 8.92184
R1160 VP.n0 VP.t3 8.92184
R1161 VP.n8 VP.n7 5.4107
R1162 VP.n20 VP.n0 5.4107
R1163 VP.n9 VP.n6 0.354861
R1164 VP.n22 VP.n21 0.354861
R1165 VP VP.n22 0.267071
R1166 VP.n10 VP.n9 0.189894
R1167 VP.n11 VP.n10 0.189894
R1168 VP.n11 VP.n3 0.189894
R1169 VP.n15 VP.n3 0.189894
R1170 VP.n16 VP.n15 0.189894
R1171 VP.n17 VP.n16 0.189894
R1172 VP.n17 VP.n1 0.189894
R1173 VP.n21 VP.n1 0.189894
R1174 VDD1 VDD1.n1 152.796
R1175 VDD1 VDD1.n0 116.459
R1176 VDD1.n0 VDD1.t3 13.7505
R1177 VDD1.n0 VDD1.t2 13.7505
R1178 VDD1.n1 VDD1.t1 13.7505
R1179 VDD1.n1 VDD1.t0 13.7505
C0 VN VDD1 0.156755f
C1 VP VDD2 0.484288f
C2 VTAIL VDD1 3.59978f
C3 VP VN 5.1658f
C4 VN VDD2 0.911461f
C5 VP VTAIL 1.8652f
C6 VDD2 VTAIL 3.66264f
C7 VP VDD1 1.23639f
C8 VN VTAIL 1.85109f
C9 VDD2 VDD1 1.34155f
C10 VDD2 B 3.632029f
C11 VDD1 B 6.62252f
C12 VTAIL B 3.763691f
C13 VN B 12.05001f
C14 VP B 10.65193f
C15 VDD1.t3 B 0.027083f
C16 VDD1.t2 B 0.027083f
C17 VDD1.n0 B 0.159334f
C18 VDD1.t1 B 0.027083f
C19 VDD1.t0 B 0.027083f
C20 VDD1.n1 B 0.386108f
C21 VP.t3 B 0.260783f
C22 VP.n0 B 0.21826f
C23 VP.n1 B 0.021616f
C24 VP.n2 B 0.042735f
C25 VP.n3 B 0.021616f
C26 VP.n4 B 0.040085f
C27 VP.t0 B 0.510052f
C28 VP.t1 B 0.49867f
C29 VP.n5 B 1.53971f
C30 VP.n6 B 1.04544f
C31 VP.t2 B 0.260783f
C32 VP.n7 B 0.21826f
C33 VP.n8 B 0.024649f
C34 VP.n9 B 0.034882f
C35 VP.n10 B 0.021616f
C36 VP.n11 B 0.021616f
C37 VP.n12 B 0.040085f
C38 VP.n13 B 0.042735f
C39 VP.n14 B 0.017458f
C40 VP.n15 B 0.021616f
C41 VP.n16 B 0.021616f
C42 VP.n17 B 0.021616f
C43 VP.n18 B 0.040085f
C44 VP.n19 B 0.040085f
C45 VP.n20 B 0.024649f
C46 VP.n21 B 0.034882f
C47 VP.n22 B 0.065663f
C48 VDD2.t0 B 0.028532f
C49 VDD2.t3 B 0.028532f
C50 VDD2.n0 B 0.392295f
C51 VDD2.t1 B 0.028532f
C52 VDD2.t2 B 0.028532f
C53 VDD2.n1 B 0.167621f
C54 VDD2.n2 B 2.72664f
C55 VTAIL.t4 B 0.168152f
C56 VTAIL.n0 B 0.321675f
C57 VTAIL.t0 B 0.168152f
C58 VTAIL.n1 B 0.444216f
C59 VTAIL.t3 B 0.168152f
C60 VTAIL.n2 B 1.04448f
C61 VTAIL.t5 B 0.168152f
C62 VTAIL.n3 B 1.04448f
C63 VTAIL.t6 B 0.168152f
C64 VTAIL.n4 B 0.444216f
C65 VTAIL.t1 B 0.168152f
C66 VTAIL.n5 B 0.444216f
C67 VTAIL.t2 B 0.168152f
C68 VTAIL.n6 B 1.04448f
C69 VTAIL.t7 B 0.168152f
C70 VTAIL.n7 B 0.913841f
C71 VN.t0 B 0.495773f
C72 VN.t3 B 0.50709f
C73 VN.n0 B 0.390661f
C74 VN.t2 B 0.495773f
C75 VN.t1 B 0.50709f
C76 VN.n1 B 1.53991f
.ends

