* NGSPICE file created from diff_pair_sample_1354.ext - technology: sky130A

.subckt diff_pair_sample_1354 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t5 VN.t0 VTAIL.t5 B.t1 sky130_fd_pr__nfet_01v8 ad=4.4031 pd=23.36 as=1.86285 ps=11.62 w=11.29 l=0.28
X1 B.t19 B.t17 B.t18 B.t14 sky130_fd_pr__nfet_01v8 ad=4.4031 pd=23.36 as=0 ps=0 w=11.29 l=0.28
X2 VTAIL.t9 VP.t0 VDD1.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=1.86285 pd=11.62 as=1.86285 ps=11.62 w=11.29 l=0.28
X3 VTAIL.t3 VN.t1 VDD2.t4 B.t0 sky130_fd_pr__nfet_01v8 ad=1.86285 pd=11.62 as=1.86285 ps=11.62 w=11.29 l=0.28
X4 VTAIL.t7 VN.t2 VDD2.t3 B.t5 sky130_fd_pr__nfet_01v8 ad=1.86285 pd=11.62 as=1.86285 ps=11.62 w=11.29 l=0.28
X5 VDD1.t4 VP.t1 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=4.4031 pd=23.36 as=1.86285 ps=11.62 w=11.29 l=0.28
X6 VDD1.t3 VP.t2 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=4.4031 pd=23.36 as=1.86285 ps=11.62 w=11.29 l=0.28
X7 B.t16 B.t13 B.t15 B.t14 sky130_fd_pr__nfet_01v8 ad=4.4031 pd=23.36 as=0 ps=0 w=11.29 l=0.28
X8 B.t12 B.t10 B.t11 B.t7 sky130_fd_pr__nfet_01v8 ad=4.4031 pd=23.36 as=0 ps=0 w=11.29 l=0.28
X9 VTAIL.t0 VP.t3 VDD1.t2 B.t0 sky130_fd_pr__nfet_01v8 ad=1.86285 pd=11.62 as=1.86285 ps=11.62 w=11.29 l=0.28
X10 VDD1.t1 VP.t4 VTAIL.t11 B.t3 sky130_fd_pr__nfet_01v8 ad=1.86285 pd=11.62 as=4.4031 ps=23.36 w=11.29 l=0.28
X11 VDD2.t2 VN.t3 VTAIL.t6 B.t4 sky130_fd_pr__nfet_01v8 ad=1.86285 pd=11.62 as=4.4031 ps=23.36 w=11.29 l=0.28
X12 B.t9 B.t6 B.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=4.4031 pd=23.36 as=0 ps=0 w=11.29 l=0.28
X13 VDD2.t1 VN.t4 VTAIL.t8 B.t2 sky130_fd_pr__nfet_01v8 ad=4.4031 pd=23.36 as=1.86285 ps=11.62 w=11.29 l=0.28
X14 VDD2.t0 VN.t5 VTAIL.t4 B.t3 sky130_fd_pr__nfet_01v8 ad=1.86285 pd=11.62 as=4.4031 ps=23.36 w=11.29 l=0.28
X15 VDD1.t0 VP.t5 VTAIL.t10 B.t4 sky130_fd_pr__nfet_01v8 ad=1.86285 pd=11.62 as=4.4031 ps=23.36 w=11.29 l=0.28
R0 VN.n2 VN.t5 1137.08
R1 VN.n0 VN.t0 1137.08
R2 VN.n6 VN.t4 1137.08
R3 VN.n4 VN.t3 1137.08
R4 VN.n1 VN.t2 1084.5
R5 VN.n5 VN.t1 1084.5
R6 VN.n7 VN.n4 161.489
R7 VN.n3 VN.n0 161.489
R8 VN.n3 VN.n2 161.3
R9 VN.n7 VN.n6 161.3
R10 VN VN.n7 39.5441
R11 VN.n1 VN.n0 36.5157
R12 VN.n2 VN.n1 36.5157
R13 VN.n6 VN.n5 36.5157
R14 VN.n5 VN.n4 36.5157
R15 VN VN.n3 0.0516364
R16 VTAIL.n250 VTAIL.n194 289.615
R17 VTAIL.n58 VTAIL.n2 289.615
R18 VTAIL.n188 VTAIL.n132 289.615
R19 VTAIL.n124 VTAIL.n68 289.615
R20 VTAIL.n215 VTAIL.n214 185
R21 VTAIL.n217 VTAIL.n216 185
R22 VTAIL.n210 VTAIL.n209 185
R23 VTAIL.n223 VTAIL.n222 185
R24 VTAIL.n225 VTAIL.n224 185
R25 VTAIL.n206 VTAIL.n205 185
R26 VTAIL.n232 VTAIL.n231 185
R27 VTAIL.n233 VTAIL.n204 185
R28 VTAIL.n235 VTAIL.n234 185
R29 VTAIL.n202 VTAIL.n201 185
R30 VTAIL.n241 VTAIL.n240 185
R31 VTAIL.n243 VTAIL.n242 185
R32 VTAIL.n198 VTAIL.n197 185
R33 VTAIL.n249 VTAIL.n248 185
R34 VTAIL.n251 VTAIL.n250 185
R35 VTAIL.n23 VTAIL.n22 185
R36 VTAIL.n25 VTAIL.n24 185
R37 VTAIL.n18 VTAIL.n17 185
R38 VTAIL.n31 VTAIL.n30 185
R39 VTAIL.n33 VTAIL.n32 185
R40 VTAIL.n14 VTAIL.n13 185
R41 VTAIL.n40 VTAIL.n39 185
R42 VTAIL.n41 VTAIL.n12 185
R43 VTAIL.n43 VTAIL.n42 185
R44 VTAIL.n10 VTAIL.n9 185
R45 VTAIL.n49 VTAIL.n48 185
R46 VTAIL.n51 VTAIL.n50 185
R47 VTAIL.n6 VTAIL.n5 185
R48 VTAIL.n57 VTAIL.n56 185
R49 VTAIL.n59 VTAIL.n58 185
R50 VTAIL.n189 VTAIL.n188 185
R51 VTAIL.n187 VTAIL.n186 185
R52 VTAIL.n136 VTAIL.n135 185
R53 VTAIL.n181 VTAIL.n180 185
R54 VTAIL.n179 VTAIL.n178 185
R55 VTAIL.n140 VTAIL.n139 185
R56 VTAIL.n144 VTAIL.n142 185
R57 VTAIL.n173 VTAIL.n172 185
R58 VTAIL.n171 VTAIL.n170 185
R59 VTAIL.n146 VTAIL.n145 185
R60 VTAIL.n165 VTAIL.n164 185
R61 VTAIL.n163 VTAIL.n162 185
R62 VTAIL.n150 VTAIL.n149 185
R63 VTAIL.n157 VTAIL.n156 185
R64 VTAIL.n155 VTAIL.n154 185
R65 VTAIL.n125 VTAIL.n124 185
R66 VTAIL.n123 VTAIL.n122 185
R67 VTAIL.n72 VTAIL.n71 185
R68 VTAIL.n117 VTAIL.n116 185
R69 VTAIL.n115 VTAIL.n114 185
R70 VTAIL.n76 VTAIL.n75 185
R71 VTAIL.n80 VTAIL.n78 185
R72 VTAIL.n109 VTAIL.n108 185
R73 VTAIL.n107 VTAIL.n106 185
R74 VTAIL.n82 VTAIL.n81 185
R75 VTAIL.n101 VTAIL.n100 185
R76 VTAIL.n99 VTAIL.n98 185
R77 VTAIL.n86 VTAIL.n85 185
R78 VTAIL.n93 VTAIL.n92 185
R79 VTAIL.n91 VTAIL.n90 185
R80 VTAIL.n213 VTAIL.t4 149.524
R81 VTAIL.n21 VTAIL.t10 149.524
R82 VTAIL.n153 VTAIL.t11 149.524
R83 VTAIL.n89 VTAIL.t6 149.524
R84 VTAIL.n216 VTAIL.n215 104.615
R85 VTAIL.n216 VTAIL.n209 104.615
R86 VTAIL.n223 VTAIL.n209 104.615
R87 VTAIL.n224 VTAIL.n223 104.615
R88 VTAIL.n224 VTAIL.n205 104.615
R89 VTAIL.n232 VTAIL.n205 104.615
R90 VTAIL.n233 VTAIL.n232 104.615
R91 VTAIL.n234 VTAIL.n233 104.615
R92 VTAIL.n234 VTAIL.n201 104.615
R93 VTAIL.n241 VTAIL.n201 104.615
R94 VTAIL.n242 VTAIL.n241 104.615
R95 VTAIL.n242 VTAIL.n197 104.615
R96 VTAIL.n249 VTAIL.n197 104.615
R97 VTAIL.n250 VTAIL.n249 104.615
R98 VTAIL.n24 VTAIL.n23 104.615
R99 VTAIL.n24 VTAIL.n17 104.615
R100 VTAIL.n31 VTAIL.n17 104.615
R101 VTAIL.n32 VTAIL.n31 104.615
R102 VTAIL.n32 VTAIL.n13 104.615
R103 VTAIL.n40 VTAIL.n13 104.615
R104 VTAIL.n41 VTAIL.n40 104.615
R105 VTAIL.n42 VTAIL.n41 104.615
R106 VTAIL.n42 VTAIL.n9 104.615
R107 VTAIL.n49 VTAIL.n9 104.615
R108 VTAIL.n50 VTAIL.n49 104.615
R109 VTAIL.n50 VTAIL.n5 104.615
R110 VTAIL.n57 VTAIL.n5 104.615
R111 VTAIL.n58 VTAIL.n57 104.615
R112 VTAIL.n188 VTAIL.n187 104.615
R113 VTAIL.n187 VTAIL.n135 104.615
R114 VTAIL.n180 VTAIL.n135 104.615
R115 VTAIL.n180 VTAIL.n179 104.615
R116 VTAIL.n179 VTAIL.n139 104.615
R117 VTAIL.n144 VTAIL.n139 104.615
R118 VTAIL.n172 VTAIL.n144 104.615
R119 VTAIL.n172 VTAIL.n171 104.615
R120 VTAIL.n171 VTAIL.n145 104.615
R121 VTAIL.n164 VTAIL.n145 104.615
R122 VTAIL.n164 VTAIL.n163 104.615
R123 VTAIL.n163 VTAIL.n149 104.615
R124 VTAIL.n156 VTAIL.n149 104.615
R125 VTAIL.n156 VTAIL.n155 104.615
R126 VTAIL.n124 VTAIL.n123 104.615
R127 VTAIL.n123 VTAIL.n71 104.615
R128 VTAIL.n116 VTAIL.n71 104.615
R129 VTAIL.n116 VTAIL.n115 104.615
R130 VTAIL.n115 VTAIL.n75 104.615
R131 VTAIL.n80 VTAIL.n75 104.615
R132 VTAIL.n108 VTAIL.n80 104.615
R133 VTAIL.n108 VTAIL.n107 104.615
R134 VTAIL.n107 VTAIL.n81 104.615
R135 VTAIL.n100 VTAIL.n81 104.615
R136 VTAIL.n100 VTAIL.n99 104.615
R137 VTAIL.n99 VTAIL.n85 104.615
R138 VTAIL.n92 VTAIL.n85 104.615
R139 VTAIL.n92 VTAIL.n91 104.615
R140 VTAIL.n215 VTAIL.t4 52.3082
R141 VTAIL.n23 VTAIL.t10 52.3082
R142 VTAIL.n155 VTAIL.t11 52.3082
R143 VTAIL.n91 VTAIL.t6 52.3082
R144 VTAIL.n131 VTAIL.n130 43.2778
R145 VTAIL.n67 VTAIL.n66 43.2778
R146 VTAIL.n1 VTAIL.n0 43.2776
R147 VTAIL.n65 VTAIL.n64 43.2776
R148 VTAIL.n255 VTAIL.n254 30.052
R149 VTAIL.n63 VTAIL.n62 30.052
R150 VTAIL.n193 VTAIL.n192 30.052
R151 VTAIL.n129 VTAIL.n128 30.052
R152 VTAIL.n67 VTAIL.n65 23.1514
R153 VTAIL.n255 VTAIL.n193 22.6255
R154 VTAIL.n235 VTAIL.n202 13.1884
R155 VTAIL.n43 VTAIL.n10 13.1884
R156 VTAIL.n142 VTAIL.n140 13.1884
R157 VTAIL.n78 VTAIL.n76 13.1884
R158 VTAIL.n236 VTAIL.n204 12.8005
R159 VTAIL.n240 VTAIL.n239 12.8005
R160 VTAIL.n44 VTAIL.n12 12.8005
R161 VTAIL.n48 VTAIL.n47 12.8005
R162 VTAIL.n178 VTAIL.n177 12.8005
R163 VTAIL.n174 VTAIL.n173 12.8005
R164 VTAIL.n114 VTAIL.n113 12.8005
R165 VTAIL.n110 VTAIL.n109 12.8005
R166 VTAIL.n231 VTAIL.n230 12.0247
R167 VTAIL.n243 VTAIL.n200 12.0247
R168 VTAIL.n39 VTAIL.n38 12.0247
R169 VTAIL.n51 VTAIL.n8 12.0247
R170 VTAIL.n181 VTAIL.n138 12.0247
R171 VTAIL.n170 VTAIL.n143 12.0247
R172 VTAIL.n117 VTAIL.n74 12.0247
R173 VTAIL.n106 VTAIL.n79 12.0247
R174 VTAIL.n229 VTAIL.n206 11.249
R175 VTAIL.n244 VTAIL.n198 11.249
R176 VTAIL.n37 VTAIL.n14 11.249
R177 VTAIL.n52 VTAIL.n6 11.249
R178 VTAIL.n182 VTAIL.n136 11.249
R179 VTAIL.n169 VTAIL.n146 11.249
R180 VTAIL.n118 VTAIL.n72 11.249
R181 VTAIL.n105 VTAIL.n82 11.249
R182 VTAIL.n226 VTAIL.n225 10.4732
R183 VTAIL.n248 VTAIL.n247 10.4732
R184 VTAIL.n34 VTAIL.n33 10.4732
R185 VTAIL.n56 VTAIL.n55 10.4732
R186 VTAIL.n186 VTAIL.n185 10.4732
R187 VTAIL.n166 VTAIL.n165 10.4732
R188 VTAIL.n122 VTAIL.n121 10.4732
R189 VTAIL.n102 VTAIL.n101 10.4732
R190 VTAIL.n214 VTAIL.n213 10.2747
R191 VTAIL.n22 VTAIL.n21 10.2747
R192 VTAIL.n154 VTAIL.n153 10.2747
R193 VTAIL.n90 VTAIL.n89 10.2747
R194 VTAIL.n222 VTAIL.n208 9.69747
R195 VTAIL.n251 VTAIL.n196 9.69747
R196 VTAIL.n30 VTAIL.n16 9.69747
R197 VTAIL.n59 VTAIL.n4 9.69747
R198 VTAIL.n189 VTAIL.n134 9.69747
R199 VTAIL.n162 VTAIL.n148 9.69747
R200 VTAIL.n125 VTAIL.n70 9.69747
R201 VTAIL.n98 VTAIL.n84 9.69747
R202 VTAIL.n254 VTAIL.n253 9.45567
R203 VTAIL.n62 VTAIL.n61 9.45567
R204 VTAIL.n192 VTAIL.n191 9.45567
R205 VTAIL.n128 VTAIL.n127 9.45567
R206 VTAIL.n253 VTAIL.n252 9.3005
R207 VTAIL.n196 VTAIL.n195 9.3005
R208 VTAIL.n247 VTAIL.n246 9.3005
R209 VTAIL.n245 VTAIL.n244 9.3005
R210 VTAIL.n200 VTAIL.n199 9.3005
R211 VTAIL.n239 VTAIL.n238 9.3005
R212 VTAIL.n212 VTAIL.n211 9.3005
R213 VTAIL.n219 VTAIL.n218 9.3005
R214 VTAIL.n221 VTAIL.n220 9.3005
R215 VTAIL.n208 VTAIL.n207 9.3005
R216 VTAIL.n227 VTAIL.n226 9.3005
R217 VTAIL.n229 VTAIL.n228 9.3005
R218 VTAIL.n230 VTAIL.n203 9.3005
R219 VTAIL.n237 VTAIL.n236 9.3005
R220 VTAIL.n61 VTAIL.n60 9.3005
R221 VTAIL.n4 VTAIL.n3 9.3005
R222 VTAIL.n55 VTAIL.n54 9.3005
R223 VTAIL.n53 VTAIL.n52 9.3005
R224 VTAIL.n8 VTAIL.n7 9.3005
R225 VTAIL.n47 VTAIL.n46 9.3005
R226 VTAIL.n20 VTAIL.n19 9.3005
R227 VTAIL.n27 VTAIL.n26 9.3005
R228 VTAIL.n29 VTAIL.n28 9.3005
R229 VTAIL.n16 VTAIL.n15 9.3005
R230 VTAIL.n35 VTAIL.n34 9.3005
R231 VTAIL.n37 VTAIL.n36 9.3005
R232 VTAIL.n38 VTAIL.n11 9.3005
R233 VTAIL.n45 VTAIL.n44 9.3005
R234 VTAIL.n152 VTAIL.n151 9.3005
R235 VTAIL.n159 VTAIL.n158 9.3005
R236 VTAIL.n161 VTAIL.n160 9.3005
R237 VTAIL.n148 VTAIL.n147 9.3005
R238 VTAIL.n167 VTAIL.n166 9.3005
R239 VTAIL.n169 VTAIL.n168 9.3005
R240 VTAIL.n143 VTAIL.n141 9.3005
R241 VTAIL.n175 VTAIL.n174 9.3005
R242 VTAIL.n191 VTAIL.n190 9.3005
R243 VTAIL.n134 VTAIL.n133 9.3005
R244 VTAIL.n185 VTAIL.n184 9.3005
R245 VTAIL.n183 VTAIL.n182 9.3005
R246 VTAIL.n138 VTAIL.n137 9.3005
R247 VTAIL.n177 VTAIL.n176 9.3005
R248 VTAIL.n88 VTAIL.n87 9.3005
R249 VTAIL.n95 VTAIL.n94 9.3005
R250 VTAIL.n97 VTAIL.n96 9.3005
R251 VTAIL.n84 VTAIL.n83 9.3005
R252 VTAIL.n103 VTAIL.n102 9.3005
R253 VTAIL.n105 VTAIL.n104 9.3005
R254 VTAIL.n79 VTAIL.n77 9.3005
R255 VTAIL.n111 VTAIL.n110 9.3005
R256 VTAIL.n127 VTAIL.n126 9.3005
R257 VTAIL.n70 VTAIL.n69 9.3005
R258 VTAIL.n121 VTAIL.n120 9.3005
R259 VTAIL.n119 VTAIL.n118 9.3005
R260 VTAIL.n74 VTAIL.n73 9.3005
R261 VTAIL.n113 VTAIL.n112 9.3005
R262 VTAIL.n221 VTAIL.n210 8.92171
R263 VTAIL.n252 VTAIL.n194 8.92171
R264 VTAIL.n29 VTAIL.n18 8.92171
R265 VTAIL.n60 VTAIL.n2 8.92171
R266 VTAIL.n190 VTAIL.n132 8.92171
R267 VTAIL.n161 VTAIL.n150 8.92171
R268 VTAIL.n126 VTAIL.n68 8.92171
R269 VTAIL.n97 VTAIL.n86 8.92171
R270 VTAIL.n218 VTAIL.n217 8.14595
R271 VTAIL.n26 VTAIL.n25 8.14595
R272 VTAIL.n158 VTAIL.n157 8.14595
R273 VTAIL.n94 VTAIL.n93 8.14595
R274 VTAIL.n214 VTAIL.n212 7.3702
R275 VTAIL.n22 VTAIL.n20 7.3702
R276 VTAIL.n154 VTAIL.n152 7.3702
R277 VTAIL.n90 VTAIL.n88 7.3702
R278 VTAIL.n217 VTAIL.n212 5.81868
R279 VTAIL.n25 VTAIL.n20 5.81868
R280 VTAIL.n157 VTAIL.n152 5.81868
R281 VTAIL.n93 VTAIL.n88 5.81868
R282 VTAIL.n218 VTAIL.n210 5.04292
R283 VTAIL.n254 VTAIL.n194 5.04292
R284 VTAIL.n26 VTAIL.n18 5.04292
R285 VTAIL.n62 VTAIL.n2 5.04292
R286 VTAIL.n192 VTAIL.n132 5.04292
R287 VTAIL.n158 VTAIL.n150 5.04292
R288 VTAIL.n128 VTAIL.n68 5.04292
R289 VTAIL.n94 VTAIL.n86 5.04292
R290 VTAIL.n222 VTAIL.n221 4.26717
R291 VTAIL.n252 VTAIL.n251 4.26717
R292 VTAIL.n30 VTAIL.n29 4.26717
R293 VTAIL.n60 VTAIL.n59 4.26717
R294 VTAIL.n190 VTAIL.n189 4.26717
R295 VTAIL.n162 VTAIL.n161 4.26717
R296 VTAIL.n126 VTAIL.n125 4.26717
R297 VTAIL.n98 VTAIL.n97 4.26717
R298 VTAIL.n225 VTAIL.n208 3.49141
R299 VTAIL.n248 VTAIL.n196 3.49141
R300 VTAIL.n33 VTAIL.n16 3.49141
R301 VTAIL.n56 VTAIL.n4 3.49141
R302 VTAIL.n186 VTAIL.n134 3.49141
R303 VTAIL.n165 VTAIL.n148 3.49141
R304 VTAIL.n122 VTAIL.n70 3.49141
R305 VTAIL.n101 VTAIL.n84 3.49141
R306 VTAIL.n213 VTAIL.n211 2.84303
R307 VTAIL.n21 VTAIL.n19 2.84303
R308 VTAIL.n153 VTAIL.n151 2.84303
R309 VTAIL.n89 VTAIL.n87 2.84303
R310 VTAIL.n226 VTAIL.n206 2.71565
R311 VTAIL.n247 VTAIL.n198 2.71565
R312 VTAIL.n34 VTAIL.n14 2.71565
R313 VTAIL.n55 VTAIL.n6 2.71565
R314 VTAIL.n185 VTAIL.n136 2.71565
R315 VTAIL.n166 VTAIL.n146 2.71565
R316 VTAIL.n121 VTAIL.n72 2.71565
R317 VTAIL.n102 VTAIL.n82 2.71565
R318 VTAIL.n231 VTAIL.n229 1.93989
R319 VTAIL.n244 VTAIL.n243 1.93989
R320 VTAIL.n39 VTAIL.n37 1.93989
R321 VTAIL.n52 VTAIL.n51 1.93989
R322 VTAIL.n182 VTAIL.n181 1.93989
R323 VTAIL.n170 VTAIL.n169 1.93989
R324 VTAIL.n118 VTAIL.n117 1.93989
R325 VTAIL.n106 VTAIL.n105 1.93989
R326 VTAIL.n0 VTAIL.t5 1.75426
R327 VTAIL.n0 VTAIL.t7 1.75426
R328 VTAIL.n64 VTAIL.t2 1.75426
R329 VTAIL.n64 VTAIL.t0 1.75426
R330 VTAIL.n130 VTAIL.t1 1.75426
R331 VTAIL.n130 VTAIL.t9 1.75426
R332 VTAIL.n66 VTAIL.t8 1.75426
R333 VTAIL.n66 VTAIL.t3 1.75426
R334 VTAIL.n230 VTAIL.n204 1.16414
R335 VTAIL.n240 VTAIL.n200 1.16414
R336 VTAIL.n38 VTAIL.n12 1.16414
R337 VTAIL.n48 VTAIL.n8 1.16414
R338 VTAIL.n178 VTAIL.n138 1.16414
R339 VTAIL.n173 VTAIL.n143 1.16414
R340 VTAIL.n114 VTAIL.n74 1.16414
R341 VTAIL.n109 VTAIL.n79 1.16414
R342 VTAIL.n131 VTAIL.n129 0.733259
R343 VTAIL.n63 VTAIL.n1 0.733259
R344 VTAIL.n129 VTAIL.n67 0.526362
R345 VTAIL.n193 VTAIL.n131 0.526362
R346 VTAIL.n65 VTAIL.n63 0.526362
R347 VTAIL.n236 VTAIL.n235 0.388379
R348 VTAIL.n239 VTAIL.n202 0.388379
R349 VTAIL.n44 VTAIL.n43 0.388379
R350 VTAIL.n47 VTAIL.n10 0.388379
R351 VTAIL.n177 VTAIL.n140 0.388379
R352 VTAIL.n174 VTAIL.n142 0.388379
R353 VTAIL.n113 VTAIL.n76 0.388379
R354 VTAIL.n110 VTAIL.n78 0.388379
R355 VTAIL VTAIL.n255 0.336707
R356 VTAIL VTAIL.n1 0.190155
R357 VTAIL.n219 VTAIL.n211 0.155672
R358 VTAIL.n220 VTAIL.n219 0.155672
R359 VTAIL.n220 VTAIL.n207 0.155672
R360 VTAIL.n227 VTAIL.n207 0.155672
R361 VTAIL.n228 VTAIL.n227 0.155672
R362 VTAIL.n228 VTAIL.n203 0.155672
R363 VTAIL.n237 VTAIL.n203 0.155672
R364 VTAIL.n238 VTAIL.n237 0.155672
R365 VTAIL.n238 VTAIL.n199 0.155672
R366 VTAIL.n245 VTAIL.n199 0.155672
R367 VTAIL.n246 VTAIL.n245 0.155672
R368 VTAIL.n246 VTAIL.n195 0.155672
R369 VTAIL.n253 VTAIL.n195 0.155672
R370 VTAIL.n27 VTAIL.n19 0.155672
R371 VTAIL.n28 VTAIL.n27 0.155672
R372 VTAIL.n28 VTAIL.n15 0.155672
R373 VTAIL.n35 VTAIL.n15 0.155672
R374 VTAIL.n36 VTAIL.n35 0.155672
R375 VTAIL.n36 VTAIL.n11 0.155672
R376 VTAIL.n45 VTAIL.n11 0.155672
R377 VTAIL.n46 VTAIL.n45 0.155672
R378 VTAIL.n46 VTAIL.n7 0.155672
R379 VTAIL.n53 VTAIL.n7 0.155672
R380 VTAIL.n54 VTAIL.n53 0.155672
R381 VTAIL.n54 VTAIL.n3 0.155672
R382 VTAIL.n61 VTAIL.n3 0.155672
R383 VTAIL.n191 VTAIL.n133 0.155672
R384 VTAIL.n184 VTAIL.n133 0.155672
R385 VTAIL.n184 VTAIL.n183 0.155672
R386 VTAIL.n183 VTAIL.n137 0.155672
R387 VTAIL.n176 VTAIL.n137 0.155672
R388 VTAIL.n176 VTAIL.n175 0.155672
R389 VTAIL.n175 VTAIL.n141 0.155672
R390 VTAIL.n168 VTAIL.n141 0.155672
R391 VTAIL.n168 VTAIL.n167 0.155672
R392 VTAIL.n167 VTAIL.n147 0.155672
R393 VTAIL.n160 VTAIL.n147 0.155672
R394 VTAIL.n160 VTAIL.n159 0.155672
R395 VTAIL.n159 VTAIL.n151 0.155672
R396 VTAIL.n127 VTAIL.n69 0.155672
R397 VTAIL.n120 VTAIL.n69 0.155672
R398 VTAIL.n120 VTAIL.n119 0.155672
R399 VTAIL.n119 VTAIL.n73 0.155672
R400 VTAIL.n112 VTAIL.n73 0.155672
R401 VTAIL.n112 VTAIL.n111 0.155672
R402 VTAIL.n111 VTAIL.n77 0.155672
R403 VTAIL.n104 VTAIL.n77 0.155672
R404 VTAIL.n104 VTAIL.n103 0.155672
R405 VTAIL.n103 VTAIL.n83 0.155672
R406 VTAIL.n96 VTAIL.n83 0.155672
R407 VTAIL.n96 VTAIL.n95 0.155672
R408 VTAIL.n95 VTAIL.n87 0.155672
R409 VDD2.n119 VDD2.n63 289.615
R410 VDD2.n56 VDD2.n0 289.615
R411 VDD2.n120 VDD2.n119 185
R412 VDD2.n118 VDD2.n117 185
R413 VDD2.n67 VDD2.n66 185
R414 VDD2.n112 VDD2.n111 185
R415 VDD2.n110 VDD2.n109 185
R416 VDD2.n71 VDD2.n70 185
R417 VDD2.n75 VDD2.n73 185
R418 VDD2.n104 VDD2.n103 185
R419 VDD2.n102 VDD2.n101 185
R420 VDD2.n77 VDD2.n76 185
R421 VDD2.n96 VDD2.n95 185
R422 VDD2.n94 VDD2.n93 185
R423 VDD2.n81 VDD2.n80 185
R424 VDD2.n88 VDD2.n87 185
R425 VDD2.n86 VDD2.n85 185
R426 VDD2.n21 VDD2.n20 185
R427 VDD2.n23 VDD2.n22 185
R428 VDD2.n16 VDD2.n15 185
R429 VDD2.n29 VDD2.n28 185
R430 VDD2.n31 VDD2.n30 185
R431 VDD2.n12 VDD2.n11 185
R432 VDD2.n38 VDD2.n37 185
R433 VDD2.n39 VDD2.n10 185
R434 VDD2.n41 VDD2.n40 185
R435 VDD2.n8 VDD2.n7 185
R436 VDD2.n47 VDD2.n46 185
R437 VDD2.n49 VDD2.n48 185
R438 VDD2.n4 VDD2.n3 185
R439 VDD2.n55 VDD2.n54 185
R440 VDD2.n57 VDD2.n56 185
R441 VDD2.n84 VDD2.t1 149.524
R442 VDD2.n19 VDD2.t5 149.524
R443 VDD2.n119 VDD2.n118 104.615
R444 VDD2.n118 VDD2.n66 104.615
R445 VDD2.n111 VDD2.n66 104.615
R446 VDD2.n111 VDD2.n110 104.615
R447 VDD2.n110 VDD2.n70 104.615
R448 VDD2.n75 VDD2.n70 104.615
R449 VDD2.n103 VDD2.n75 104.615
R450 VDD2.n103 VDD2.n102 104.615
R451 VDD2.n102 VDD2.n76 104.615
R452 VDD2.n95 VDD2.n76 104.615
R453 VDD2.n95 VDD2.n94 104.615
R454 VDD2.n94 VDD2.n80 104.615
R455 VDD2.n87 VDD2.n80 104.615
R456 VDD2.n87 VDD2.n86 104.615
R457 VDD2.n22 VDD2.n21 104.615
R458 VDD2.n22 VDD2.n15 104.615
R459 VDD2.n29 VDD2.n15 104.615
R460 VDD2.n30 VDD2.n29 104.615
R461 VDD2.n30 VDD2.n11 104.615
R462 VDD2.n38 VDD2.n11 104.615
R463 VDD2.n39 VDD2.n38 104.615
R464 VDD2.n40 VDD2.n39 104.615
R465 VDD2.n40 VDD2.n7 104.615
R466 VDD2.n47 VDD2.n7 104.615
R467 VDD2.n48 VDD2.n47 104.615
R468 VDD2.n48 VDD2.n3 104.615
R469 VDD2.n55 VDD2.n3 104.615
R470 VDD2.n56 VDD2.n55 104.615
R471 VDD2.n62 VDD2.n61 60.0325
R472 VDD2 VDD2.n125 60.0297
R473 VDD2.n86 VDD2.t1 52.3082
R474 VDD2.n21 VDD2.t5 52.3082
R475 VDD2.n62 VDD2.n60 47.0699
R476 VDD2.n124 VDD2.n123 46.7308
R477 VDD2.n124 VDD2.n62 35.1571
R478 VDD2.n73 VDD2.n71 13.1884
R479 VDD2.n41 VDD2.n8 13.1884
R480 VDD2.n109 VDD2.n108 12.8005
R481 VDD2.n105 VDD2.n104 12.8005
R482 VDD2.n42 VDD2.n10 12.8005
R483 VDD2.n46 VDD2.n45 12.8005
R484 VDD2.n112 VDD2.n69 12.0247
R485 VDD2.n101 VDD2.n74 12.0247
R486 VDD2.n37 VDD2.n36 12.0247
R487 VDD2.n49 VDD2.n6 12.0247
R488 VDD2.n113 VDD2.n67 11.249
R489 VDD2.n100 VDD2.n77 11.249
R490 VDD2.n35 VDD2.n12 11.249
R491 VDD2.n50 VDD2.n4 11.249
R492 VDD2.n117 VDD2.n116 10.4732
R493 VDD2.n97 VDD2.n96 10.4732
R494 VDD2.n32 VDD2.n31 10.4732
R495 VDD2.n54 VDD2.n53 10.4732
R496 VDD2.n85 VDD2.n84 10.2747
R497 VDD2.n20 VDD2.n19 10.2747
R498 VDD2.n120 VDD2.n65 9.69747
R499 VDD2.n93 VDD2.n79 9.69747
R500 VDD2.n28 VDD2.n14 9.69747
R501 VDD2.n57 VDD2.n2 9.69747
R502 VDD2.n123 VDD2.n122 9.45567
R503 VDD2.n60 VDD2.n59 9.45567
R504 VDD2.n83 VDD2.n82 9.3005
R505 VDD2.n90 VDD2.n89 9.3005
R506 VDD2.n92 VDD2.n91 9.3005
R507 VDD2.n79 VDD2.n78 9.3005
R508 VDD2.n98 VDD2.n97 9.3005
R509 VDD2.n100 VDD2.n99 9.3005
R510 VDD2.n74 VDD2.n72 9.3005
R511 VDD2.n106 VDD2.n105 9.3005
R512 VDD2.n122 VDD2.n121 9.3005
R513 VDD2.n65 VDD2.n64 9.3005
R514 VDD2.n116 VDD2.n115 9.3005
R515 VDD2.n114 VDD2.n113 9.3005
R516 VDD2.n69 VDD2.n68 9.3005
R517 VDD2.n108 VDD2.n107 9.3005
R518 VDD2.n59 VDD2.n58 9.3005
R519 VDD2.n2 VDD2.n1 9.3005
R520 VDD2.n53 VDD2.n52 9.3005
R521 VDD2.n51 VDD2.n50 9.3005
R522 VDD2.n6 VDD2.n5 9.3005
R523 VDD2.n45 VDD2.n44 9.3005
R524 VDD2.n18 VDD2.n17 9.3005
R525 VDD2.n25 VDD2.n24 9.3005
R526 VDD2.n27 VDD2.n26 9.3005
R527 VDD2.n14 VDD2.n13 9.3005
R528 VDD2.n33 VDD2.n32 9.3005
R529 VDD2.n35 VDD2.n34 9.3005
R530 VDD2.n36 VDD2.n9 9.3005
R531 VDD2.n43 VDD2.n42 9.3005
R532 VDD2.n121 VDD2.n63 8.92171
R533 VDD2.n92 VDD2.n81 8.92171
R534 VDD2.n27 VDD2.n16 8.92171
R535 VDD2.n58 VDD2.n0 8.92171
R536 VDD2.n89 VDD2.n88 8.14595
R537 VDD2.n24 VDD2.n23 8.14595
R538 VDD2.n85 VDD2.n83 7.3702
R539 VDD2.n20 VDD2.n18 7.3702
R540 VDD2.n88 VDD2.n83 5.81868
R541 VDD2.n23 VDD2.n18 5.81868
R542 VDD2.n123 VDD2.n63 5.04292
R543 VDD2.n89 VDD2.n81 5.04292
R544 VDD2.n24 VDD2.n16 5.04292
R545 VDD2.n60 VDD2.n0 5.04292
R546 VDD2.n121 VDD2.n120 4.26717
R547 VDD2.n93 VDD2.n92 4.26717
R548 VDD2.n28 VDD2.n27 4.26717
R549 VDD2.n58 VDD2.n57 4.26717
R550 VDD2.n117 VDD2.n65 3.49141
R551 VDD2.n96 VDD2.n79 3.49141
R552 VDD2.n31 VDD2.n14 3.49141
R553 VDD2.n54 VDD2.n2 3.49141
R554 VDD2.n84 VDD2.n82 2.84303
R555 VDD2.n19 VDD2.n17 2.84303
R556 VDD2.n116 VDD2.n67 2.71565
R557 VDD2.n97 VDD2.n77 2.71565
R558 VDD2.n32 VDD2.n12 2.71565
R559 VDD2.n53 VDD2.n4 2.71565
R560 VDD2.n113 VDD2.n112 1.93989
R561 VDD2.n101 VDD2.n100 1.93989
R562 VDD2.n37 VDD2.n35 1.93989
R563 VDD2.n50 VDD2.n49 1.93989
R564 VDD2.n125 VDD2.t4 1.75426
R565 VDD2.n125 VDD2.t2 1.75426
R566 VDD2.n61 VDD2.t3 1.75426
R567 VDD2.n61 VDD2.t0 1.75426
R568 VDD2.n109 VDD2.n69 1.16414
R569 VDD2.n104 VDD2.n74 1.16414
R570 VDD2.n36 VDD2.n10 1.16414
R571 VDD2.n46 VDD2.n6 1.16414
R572 VDD2 VDD2.n124 0.453086
R573 VDD2.n108 VDD2.n71 0.388379
R574 VDD2.n105 VDD2.n73 0.388379
R575 VDD2.n42 VDD2.n41 0.388379
R576 VDD2.n45 VDD2.n8 0.388379
R577 VDD2.n122 VDD2.n64 0.155672
R578 VDD2.n115 VDD2.n64 0.155672
R579 VDD2.n115 VDD2.n114 0.155672
R580 VDD2.n114 VDD2.n68 0.155672
R581 VDD2.n107 VDD2.n68 0.155672
R582 VDD2.n107 VDD2.n106 0.155672
R583 VDD2.n106 VDD2.n72 0.155672
R584 VDD2.n99 VDD2.n72 0.155672
R585 VDD2.n99 VDD2.n98 0.155672
R586 VDD2.n98 VDD2.n78 0.155672
R587 VDD2.n91 VDD2.n78 0.155672
R588 VDD2.n91 VDD2.n90 0.155672
R589 VDD2.n90 VDD2.n82 0.155672
R590 VDD2.n25 VDD2.n17 0.155672
R591 VDD2.n26 VDD2.n25 0.155672
R592 VDD2.n26 VDD2.n13 0.155672
R593 VDD2.n33 VDD2.n13 0.155672
R594 VDD2.n34 VDD2.n33 0.155672
R595 VDD2.n34 VDD2.n9 0.155672
R596 VDD2.n43 VDD2.n9 0.155672
R597 VDD2.n44 VDD2.n43 0.155672
R598 VDD2.n44 VDD2.n5 0.155672
R599 VDD2.n51 VDD2.n5 0.155672
R600 VDD2.n52 VDD2.n51 0.155672
R601 VDD2.n52 VDD2.n1 0.155672
R602 VDD2.n59 VDD2.n1 0.155672
R603 B.n79 B.t6 1190.88
R604 B.n77 B.t10 1190.88
R605 B.n329 B.t13 1190.88
R606 B.n327 B.t17 1190.88
R607 B.n577 B.n576 585
R608 B.n578 B.n577 585
R609 B.n253 B.n75 585
R610 B.n252 B.n251 585
R611 B.n250 B.n249 585
R612 B.n248 B.n247 585
R613 B.n246 B.n245 585
R614 B.n244 B.n243 585
R615 B.n242 B.n241 585
R616 B.n240 B.n239 585
R617 B.n238 B.n237 585
R618 B.n236 B.n235 585
R619 B.n234 B.n233 585
R620 B.n232 B.n231 585
R621 B.n230 B.n229 585
R622 B.n228 B.n227 585
R623 B.n226 B.n225 585
R624 B.n224 B.n223 585
R625 B.n222 B.n221 585
R626 B.n220 B.n219 585
R627 B.n218 B.n217 585
R628 B.n216 B.n215 585
R629 B.n214 B.n213 585
R630 B.n212 B.n211 585
R631 B.n210 B.n209 585
R632 B.n208 B.n207 585
R633 B.n206 B.n205 585
R634 B.n204 B.n203 585
R635 B.n202 B.n201 585
R636 B.n200 B.n199 585
R637 B.n198 B.n197 585
R638 B.n196 B.n195 585
R639 B.n194 B.n193 585
R640 B.n192 B.n191 585
R641 B.n190 B.n189 585
R642 B.n188 B.n187 585
R643 B.n186 B.n185 585
R644 B.n184 B.n183 585
R645 B.n182 B.n181 585
R646 B.n180 B.n179 585
R647 B.n178 B.n177 585
R648 B.n175 B.n174 585
R649 B.n173 B.n172 585
R650 B.n171 B.n170 585
R651 B.n169 B.n168 585
R652 B.n167 B.n166 585
R653 B.n165 B.n164 585
R654 B.n163 B.n162 585
R655 B.n161 B.n160 585
R656 B.n159 B.n158 585
R657 B.n157 B.n156 585
R658 B.n155 B.n154 585
R659 B.n153 B.n152 585
R660 B.n151 B.n150 585
R661 B.n149 B.n148 585
R662 B.n147 B.n146 585
R663 B.n145 B.n144 585
R664 B.n143 B.n142 585
R665 B.n141 B.n140 585
R666 B.n139 B.n138 585
R667 B.n137 B.n136 585
R668 B.n135 B.n134 585
R669 B.n133 B.n132 585
R670 B.n131 B.n130 585
R671 B.n129 B.n128 585
R672 B.n127 B.n126 585
R673 B.n125 B.n124 585
R674 B.n123 B.n122 585
R675 B.n121 B.n120 585
R676 B.n119 B.n118 585
R677 B.n117 B.n116 585
R678 B.n115 B.n114 585
R679 B.n113 B.n112 585
R680 B.n111 B.n110 585
R681 B.n109 B.n108 585
R682 B.n107 B.n106 585
R683 B.n105 B.n104 585
R684 B.n103 B.n102 585
R685 B.n101 B.n100 585
R686 B.n99 B.n98 585
R687 B.n97 B.n96 585
R688 B.n95 B.n94 585
R689 B.n93 B.n92 585
R690 B.n91 B.n90 585
R691 B.n89 B.n88 585
R692 B.n87 B.n86 585
R693 B.n85 B.n84 585
R694 B.n83 B.n82 585
R695 B.n31 B.n30 585
R696 B.n581 B.n580 585
R697 B.n575 B.n76 585
R698 B.n76 B.n28 585
R699 B.n574 B.n27 585
R700 B.n585 B.n27 585
R701 B.n573 B.n26 585
R702 B.n586 B.n26 585
R703 B.n572 B.n25 585
R704 B.n587 B.n25 585
R705 B.n571 B.n570 585
R706 B.n570 B.n24 585
R707 B.n569 B.n20 585
R708 B.n593 B.n20 585
R709 B.n568 B.n19 585
R710 B.n594 B.n19 585
R711 B.n567 B.n18 585
R712 B.n595 B.n18 585
R713 B.n566 B.n565 585
R714 B.n565 B.n14 585
R715 B.n564 B.n13 585
R716 B.n601 B.n13 585
R717 B.n563 B.n12 585
R718 B.n602 B.n12 585
R719 B.n562 B.n11 585
R720 B.n603 B.n11 585
R721 B.n561 B.n560 585
R722 B.n560 B.n559 585
R723 B.n558 B.n557 585
R724 B.n558 B.t1 585
R725 B.n556 B.n7 585
R726 B.n610 B.n7 585
R727 B.n555 B.n6 585
R728 B.n611 B.n6 585
R729 B.n554 B.n5 585
R730 B.n612 B.n5 585
R731 B.n553 B.n552 585
R732 B.n552 B.n4 585
R733 B.n551 B.n254 585
R734 B.n551 B.t4 585
R735 B.n542 B.n255 585
R736 B.n256 B.n255 585
R737 B.n544 B.n543 585
R738 B.n545 B.n544 585
R739 B.n541 B.n261 585
R740 B.n261 B.n260 585
R741 B.n540 B.n539 585
R742 B.n539 B.n538 585
R743 B.n263 B.n262 585
R744 B.n264 B.n263 585
R745 B.n531 B.n530 585
R746 B.n532 B.n531 585
R747 B.n529 B.n269 585
R748 B.n269 B.n268 585
R749 B.n528 B.n527 585
R750 B.n527 B.n526 585
R751 B.n271 B.n270 585
R752 B.n519 B.n271 585
R753 B.n518 B.n517 585
R754 B.n520 B.n518 585
R755 B.n516 B.n276 585
R756 B.n276 B.n275 585
R757 B.n515 B.n514 585
R758 B.n514 B.n513 585
R759 B.n278 B.n277 585
R760 B.n279 B.n278 585
R761 B.n509 B.n508 585
R762 B.n282 B.n281 585
R763 B.n505 B.n504 585
R764 B.n506 B.n505 585
R765 B.n503 B.n326 585
R766 B.n502 B.n501 585
R767 B.n500 B.n499 585
R768 B.n498 B.n497 585
R769 B.n496 B.n495 585
R770 B.n494 B.n493 585
R771 B.n492 B.n491 585
R772 B.n490 B.n489 585
R773 B.n488 B.n487 585
R774 B.n486 B.n485 585
R775 B.n484 B.n483 585
R776 B.n482 B.n481 585
R777 B.n480 B.n479 585
R778 B.n478 B.n477 585
R779 B.n476 B.n475 585
R780 B.n474 B.n473 585
R781 B.n472 B.n471 585
R782 B.n470 B.n469 585
R783 B.n468 B.n467 585
R784 B.n466 B.n465 585
R785 B.n464 B.n463 585
R786 B.n462 B.n461 585
R787 B.n460 B.n459 585
R788 B.n458 B.n457 585
R789 B.n456 B.n455 585
R790 B.n454 B.n453 585
R791 B.n452 B.n451 585
R792 B.n450 B.n449 585
R793 B.n448 B.n447 585
R794 B.n446 B.n445 585
R795 B.n444 B.n443 585
R796 B.n442 B.n441 585
R797 B.n440 B.n439 585
R798 B.n438 B.n437 585
R799 B.n436 B.n435 585
R800 B.n434 B.n433 585
R801 B.n432 B.n431 585
R802 B.n429 B.n428 585
R803 B.n427 B.n426 585
R804 B.n425 B.n424 585
R805 B.n423 B.n422 585
R806 B.n421 B.n420 585
R807 B.n419 B.n418 585
R808 B.n417 B.n416 585
R809 B.n415 B.n414 585
R810 B.n413 B.n412 585
R811 B.n411 B.n410 585
R812 B.n409 B.n408 585
R813 B.n407 B.n406 585
R814 B.n405 B.n404 585
R815 B.n403 B.n402 585
R816 B.n401 B.n400 585
R817 B.n399 B.n398 585
R818 B.n397 B.n396 585
R819 B.n395 B.n394 585
R820 B.n393 B.n392 585
R821 B.n391 B.n390 585
R822 B.n389 B.n388 585
R823 B.n387 B.n386 585
R824 B.n385 B.n384 585
R825 B.n383 B.n382 585
R826 B.n381 B.n380 585
R827 B.n379 B.n378 585
R828 B.n377 B.n376 585
R829 B.n375 B.n374 585
R830 B.n373 B.n372 585
R831 B.n371 B.n370 585
R832 B.n369 B.n368 585
R833 B.n367 B.n366 585
R834 B.n365 B.n364 585
R835 B.n363 B.n362 585
R836 B.n361 B.n360 585
R837 B.n359 B.n358 585
R838 B.n357 B.n356 585
R839 B.n355 B.n354 585
R840 B.n353 B.n352 585
R841 B.n351 B.n350 585
R842 B.n349 B.n348 585
R843 B.n347 B.n346 585
R844 B.n345 B.n344 585
R845 B.n343 B.n342 585
R846 B.n341 B.n340 585
R847 B.n339 B.n338 585
R848 B.n337 B.n336 585
R849 B.n335 B.n334 585
R850 B.n333 B.n332 585
R851 B.n510 B.n280 585
R852 B.n280 B.n279 585
R853 B.n512 B.n511 585
R854 B.n513 B.n512 585
R855 B.n274 B.n273 585
R856 B.n275 B.n274 585
R857 B.n522 B.n521 585
R858 B.n521 B.n520 585
R859 B.n523 B.n272 585
R860 B.n519 B.n272 585
R861 B.n525 B.n524 585
R862 B.n526 B.n525 585
R863 B.n267 B.n266 585
R864 B.n268 B.n267 585
R865 B.n534 B.n533 585
R866 B.n533 B.n532 585
R867 B.n535 B.n265 585
R868 B.n265 B.n264 585
R869 B.n537 B.n536 585
R870 B.n538 B.n537 585
R871 B.n259 B.n258 585
R872 B.n260 B.n259 585
R873 B.n547 B.n546 585
R874 B.n546 B.n545 585
R875 B.n548 B.n257 585
R876 B.n257 B.n256 585
R877 B.n550 B.n549 585
R878 B.t4 B.n550 585
R879 B.n3 B.n0 585
R880 B.n4 B.n3 585
R881 B.n609 B.n1 585
R882 B.n610 B.n609 585
R883 B.n608 B.n607 585
R884 B.n608 B.t1 585
R885 B.n606 B.n8 585
R886 B.n559 B.n8 585
R887 B.n605 B.n604 585
R888 B.n604 B.n603 585
R889 B.n10 B.n9 585
R890 B.n602 B.n10 585
R891 B.n600 B.n599 585
R892 B.n601 B.n600 585
R893 B.n598 B.n15 585
R894 B.n15 B.n14 585
R895 B.n597 B.n596 585
R896 B.n596 B.n595 585
R897 B.n17 B.n16 585
R898 B.n594 B.n17 585
R899 B.n592 B.n591 585
R900 B.n593 B.n592 585
R901 B.n590 B.n21 585
R902 B.n24 B.n21 585
R903 B.n589 B.n588 585
R904 B.n588 B.n587 585
R905 B.n23 B.n22 585
R906 B.n586 B.n23 585
R907 B.n584 B.n583 585
R908 B.n585 B.n584 585
R909 B.n582 B.n29 585
R910 B.n29 B.n28 585
R911 B.n613 B.n612 585
R912 B.n611 B.n2 585
R913 B.n580 B.n29 434.841
R914 B.n577 B.n76 434.841
R915 B.n332 B.n278 434.841
R916 B.n508 B.n280 434.841
R917 B.n77 B.t11 281.545
R918 B.n329 B.t16 281.545
R919 B.n79 B.t8 281.545
R920 B.n327 B.t19 281.545
R921 B.n78 B.t12 269.714
R922 B.n330 B.t15 269.714
R923 B.n80 B.t9 269.714
R924 B.n328 B.t18 269.714
R925 B.n578 B.n74 256.663
R926 B.n578 B.n73 256.663
R927 B.n578 B.n72 256.663
R928 B.n578 B.n71 256.663
R929 B.n578 B.n70 256.663
R930 B.n578 B.n69 256.663
R931 B.n578 B.n68 256.663
R932 B.n578 B.n67 256.663
R933 B.n578 B.n66 256.663
R934 B.n578 B.n65 256.663
R935 B.n578 B.n64 256.663
R936 B.n578 B.n63 256.663
R937 B.n578 B.n62 256.663
R938 B.n578 B.n61 256.663
R939 B.n578 B.n60 256.663
R940 B.n578 B.n59 256.663
R941 B.n578 B.n58 256.663
R942 B.n578 B.n57 256.663
R943 B.n578 B.n56 256.663
R944 B.n578 B.n55 256.663
R945 B.n578 B.n54 256.663
R946 B.n578 B.n53 256.663
R947 B.n578 B.n52 256.663
R948 B.n578 B.n51 256.663
R949 B.n578 B.n50 256.663
R950 B.n578 B.n49 256.663
R951 B.n578 B.n48 256.663
R952 B.n578 B.n47 256.663
R953 B.n578 B.n46 256.663
R954 B.n578 B.n45 256.663
R955 B.n578 B.n44 256.663
R956 B.n578 B.n43 256.663
R957 B.n578 B.n42 256.663
R958 B.n578 B.n41 256.663
R959 B.n578 B.n40 256.663
R960 B.n578 B.n39 256.663
R961 B.n578 B.n38 256.663
R962 B.n578 B.n37 256.663
R963 B.n578 B.n36 256.663
R964 B.n578 B.n35 256.663
R965 B.n578 B.n34 256.663
R966 B.n578 B.n33 256.663
R967 B.n578 B.n32 256.663
R968 B.n579 B.n578 256.663
R969 B.n507 B.n506 256.663
R970 B.n506 B.n283 256.663
R971 B.n506 B.n284 256.663
R972 B.n506 B.n285 256.663
R973 B.n506 B.n286 256.663
R974 B.n506 B.n287 256.663
R975 B.n506 B.n288 256.663
R976 B.n506 B.n289 256.663
R977 B.n506 B.n290 256.663
R978 B.n506 B.n291 256.663
R979 B.n506 B.n292 256.663
R980 B.n506 B.n293 256.663
R981 B.n506 B.n294 256.663
R982 B.n506 B.n295 256.663
R983 B.n506 B.n296 256.663
R984 B.n506 B.n297 256.663
R985 B.n506 B.n298 256.663
R986 B.n506 B.n299 256.663
R987 B.n506 B.n300 256.663
R988 B.n506 B.n301 256.663
R989 B.n506 B.n302 256.663
R990 B.n506 B.n303 256.663
R991 B.n506 B.n304 256.663
R992 B.n506 B.n305 256.663
R993 B.n506 B.n306 256.663
R994 B.n506 B.n307 256.663
R995 B.n506 B.n308 256.663
R996 B.n506 B.n309 256.663
R997 B.n506 B.n310 256.663
R998 B.n506 B.n311 256.663
R999 B.n506 B.n312 256.663
R1000 B.n506 B.n313 256.663
R1001 B.n506 B.n314 256.663
R1002 B.n506 B.n315 256.663
R1003 B.n506 B.n316 256.663
R1004 B.n506 B.n317 256.663
R1005 B.n506 B.n318 256.663
R1006 B.n506 B.n319 256.663
R1007 B.n506 B.n320 256.663
R1008 B.n506 B.n321 256.663
R1009 B.n506 B.n322 256.663
R1010 B.n506 B.n323 256.663
R1011 B.n506 B.n324 256.663
R1012 B.n506 B.n325 256.663
R1013 B.n615 B.n614 256.663
R1014 B.n82 B.n31 163.367
R1015 B.n86 B.n85 163.367
R1016 B.n90 B.n89 163.367
R1017 B.n94 B.n93 163.367
R1018 B.n98 B.n97 163.367
R1019 B.n102 B.n101 163.367
R1020 B.n106 B.n105 163.367
R1021 B.n110 B.n109 163.367
R1022 B.n114 B.n113 163.367
R1023 B.n118 B.n117 163.367
R1024 B.n122 B.n121 163.367
R1025 B.n126 B.n125 163.367
R1026 B.n130 B.n129 163.367
R1027 B.n134 B.n133 163.367
R1028 B.n138 B.n137 163.367
R1029 B.n142 B.n141 163.367
R1030 B.n146 B.n145 163.367
R1031 B.n150 B.n149 163.367
R1032 B.n154 B.n153 163.367
R1033 B.n158 B.n157 163.367
R1034 B.n162 B.n161 163.367
R1035 B.n166 B.n165 163.367
R1036 B.n170 B.n169 163.367
R1037 B.n174 B.n173 163.367
R1038 B.n179 B.n178 163.367
R1039 B.n183 B.n182 163.367
R1040 B.n187 B.n186 163.367
R1041 B.n191 B.n190 163.367
R1042 B.n195 B.n194 163.367
R1043 B.n199 B.n198 163.367
R1044 B.n203 B.n202 163.367
R1045 B.n207 B.n206 163.367
R1046 B.n211 B.n210 163.367
R1047 B.n215 B.n214 163.367
R1048 B.n219 B.n218 163.367
R1049 B.n223 B.n222 163.367
R1050 B.n227 B.n226 163.367
R1051 B.n231 B.n230 163.367
R1052 B.n235 B.n234 163.367
R1053 B.n239 B.n238 163.367
R1054 B.n243 B.n242 163.367
R1055 B.n247 B.n246 163.367
R1056 B.n251 B.n250 163.367
R1057 B.n577 B.n75 163.367
R1058 B.n514 B.n278 163.367
R1059 B.n514 B.n276 163.367
R1060 B.n518 B.n276 163.367
R1061 B.n518 B.n271 163.367
R1062 B.n527 B.n271 163.367
R1063 B.n527 B.n269 163.367
R1064 B.n531 B.n269 163.367
R1065 B.n531 B.n263 163.367
R1066 B.n539 B.n263 163.367
R1067 B.n539 B.n261 163.367
R1068 B.n544 B.n261 163.367
R1069 B.n544 B.n255 163.367
R1070 B.n551 B.n255 163.367
R1071 B.n552 B.n551 163.367
R1072 B.n552 B.n5 163.367
R1073 B.n6 B.n5 163.367
R1074 B.n7 B.n6 163.367
R1075 B.n558 B.n7 163.367
R1076 B.n560 B.n558 163.367
R1077 B.n560 B.n11 163.367
R1078 B.n12 B.n11 163.367
R1079 B.n13 B.n12 163.367
R1080 B.n565 B.n13 163.367
R1081 B.n565 B.n18 163.367
R1082 B.n19 B.n18 163.367
R1083 B.n20 B.n19 163.367
R1084 B.n570 B.n20 163.367
R1085 B.n570 B.n25 163.367
R1086 B.n26 B.n25 163.367
R1087 B.n27 B.n26 163.367
R1088 B.n76 B.n27 163.367
R1089 B.n505 B.n282 163.367
R1090 B.n505 B.n326 163.367
R1091 B.n501 B.n500 163.367
R1092 B.n497 B.n496 163.367
R1093 B.n493 B.n492 163.367
R1094 B.n489 B.n488 163.367
R1095 B.n485 B.n484 163.367
R1096 B.n481 B.n480 163.367
R1097 B.n477 B.n476 163.367
R1098 B.n473 B.n472 163.367
R1099 B.n469 B.n468 163.367
R1100 B.n465 B.n464 163.367
R1101 B.n461 B.n460 163.367
R1102 B.n457 B.n456 163.367
R1103 B.n453 B.n452 163.367
R1104 B.n449 B.n448 163.367
R1105 B.n445 B.n444 163.367
R1106 B.n441 B.n440 163.367
R1107 B.n437 B.n436 163.367
R1108 B.n433 B.n432 163.367
R1109 B.n428 B.n427 163.367
R1110 B.n424 B.n423 163.367
R1111 B.n420 B.n419 163.367
R1112 B.n416 B.n415 163.367
R1113 B.n412 B.n411 163.367
R1114 B.n408 B.n407 163.367
R1115 B.n404 B.n403 163.367
R1116 B.n400 B.n399 163.367
R1117 B.n396 B.n395 163.367
R1118 B.n392 B.n391 163.367
R1119 B.n388 B.n387 163.367
R1120 B.n384 B.n383 163.367
R1121 B.n380 B.n379 163.367
R1122 B.n376 B.n375 163.367
R1123 B.n372 B.n371 163.367
R1124 B.n368 B.n367 163.367
R1125 B.n364 B.n363 163.367
R1126 B.n360 B.n359 163.367
R1127 B.n356 B.n355 163.367
R1128 B.n352 B.n351 163.367
R1129 B.n348 B.n347 163.367
R1130 B.n344 B.n343 163.367
R1131 B.n340 B.n339 163.367
R1132 B.n336 B.n335 163.367
R1133 B.n512 B.n280 163.367
R1134 B.n512 B.n274 163.367
R1135 B.n521 B.n274 163.367
R1136 B.n521 B.n272 163.367
R1137 B.n525 B.n272 163.367
R1138 B.n525 B.n267 163.367
R1139 B.n533 B.n267 163.367
R1140 B.n533 B.n265 163.367
R1141 B.n537 B.n265 163.367
R1142 B.n537 B.n259 163.367
R1143 B.n546 B.n259 163.367
R1144 B.n546 B.n257 163.367
R1145 B.n550 B.n257 163.367
R1146 B.n550 B.n3 163.367
R1147 B.n613 B.n3 163.367
R1148 B.n609 B.n2 163.367
R1149 B.n609 B.n608 163.367
R1150 B.n608 B.n8 163.367
R1151 B.n604 B.n8 163.367
R1152 B.n604 B.n10 163.367
R1153 B.n600 B.n10 163.367
R1154 B.n600 B.n15 163.367
R1155 B.n596 B.n15 163.367
R1156 B.n596 B.n17 163.367
R1157 B.n592 B.n17 163.367
R1158 B.n592 B.n21 163.367
R1159 B.n588 B.n21 163.367
R1160 B.n588 B.n23 163.367
R1161 B.n584 B.n23 163.367
R1162 B.n584 B.n29 163.367
R1163 B.n506 B.n279 72.382
R1164 B.n578 B.n28 72.382
R1165 B.n580 B.n579 71.676
R1166 B.n82 B.n32 71.676
R1167 B.n86 B.n33 71.676
R1168 B.n90 B.n34 71.676
R1169 B.n94 B.n35 71.676
R1170 B.n98 B.n36 71.676
R1171 B.n102 B.n37 71.676
R1172 B.n106 B.n38 71.676
R1173 B.n110 B.n39 71.676
R1174 B.n114 B.n40 71.676
R1175 B.n118 B.n41 71.676
R1176 B.n122 B.n42 71.676
R1177 B.n126 B.n43 71.676
R1178 B.n130 B.n44 71.676
R1179 B.n134 B.n45 71.676
R1180 B.n138 B.n46 71.676
R1181 B.n142 B.n47 71.676
R1182 B.n146 B.n48 71.676
R1183 B.n150 B.n49 71.676
R1184 B.n154 B.n50 71.676
R1185 B.n158 B.n51 71.676
R1186 B.n162 B.n52 71.676
R1187 B.n166 B.n53 71.676
R1188 B.n170 B.n54 71.676
R1189 B.n174 B.n55 71.676
R1190 B.n179 B.n56 71.676
R1191 B.n183 B.n57 71.676
R1192 B.n187 B.n58 71.676
R1193 B.n191 B.n59 71.676
R1194 B.n195 B.n60 71.676
R1195 B.n199 B.n61 71.676
R1196 B.n203 B.n62 71.676
R1197 B.n207 B.n63 71.676
R1198 B.n211 B.n64 71.676
R1199 B.n215 B.n65 71.676
R1200 B.n219 B.n66 71.676
R1201 B.n223 B.n67 71.676
R1202 B.n227 B.n68 71.676
R1203 B.n231 B.n69 71.676
R1204 B.n235 B.n70 71.676
R1205 B.n239 B.n71 71.676
R1206 B.n243 B.n72 71.676
R1207 B.n247 B.n73 71.676
R1208 B.n251 B.n74 71.676
R1209 B.n75 B.n74 71.676
R1210 B.n250 B.n73 71.676
R1211 B.n246 B.n72 71.676
R1212 B.n242 B.n71 71.676
R1213 B.n238 B.n70 71.676
R1214 B.n234 B.n69 71.676
R1215 B.n230 B.n68 71.676
R1216 B.n226 B.n67 71.676
R1217 B.n222 B.n66 71.676
R1218 B.n218 B.n65 71.676
R1219 B.n214 B.n64 71.676
R1220 B.n210 B.n63 71.676
R1221 B.n206 B.n62 71.676
R1222 B.n202 B.n61 71.676
R1223 B.n198 B.n60 71.676
R1224 B.n194 B.n59 71.676
R1225 B.n190 B.n58 71.676
R1226 B.n186 B.n57 71.676
R1227 B.n182 B.n56 71.676
R1228 B.n178 B.n55 71.676
R1229 B.n173 B.n54 71.676
R1230 B.n169 B.n53 71.676
R1231 B.n165 B.n52 71.676
R1232 B.n161 B.n51 71.676
R1233 B.n157 B.n50 71.676
R1234 B.n153 B.n49 71.676
R1235 B.n149 B.n48 71.676
R1236 B.n145 B.n47 71.676
R1237 B.n141 B.n46 71.676
R1238 B.n137 B.n45 71.676
R1239 B.n133 B.n44 71.676
R1240 B.n129 B.n43 71.676
R1241 B.n125 B.n42 71.676
R1242 B.n121 B.n41 71.676
R1243 B.n117 B.n40 71.676
R1244 B.n113 B.n39 71.676
R1245 B.n109 B.n38 71.676
R1246 B.n105 B.n37 71.676
R1247 B.n101 B.n36 71.676
R1248 B.n97 B.n35 71.676
R1249 B.n93 B.n34 71.676
R1250 B.n89 B.n33 71.676
R1251 B.n85 B.n32 71.676
R1252 B.n579 B.n31 71.676
R1253 B.n508 B.n507 71.676
R1254 B.n326 B.n283 71.676
R1255 B.n500 B.n284 71.676
R1256 B.n496 B.n285 71.676
R1257 B.n492 B.n286 71.676
R1258 B.n488 B.n287 71.676
R1259 B.n484 B.n288 71.676
R1260 B.n480 B.n289 71.676
R1261 B.n476 B.n290 71.676
R1262 B.n472 B.n291 71.676
R1263 B.n468 B.n292 71.676
R1264 B.n464 B.n293 71.676
R1265 B.n460 B.n294 71.676
R1266 B.n456 B.n295 71.676
R1267 B.n452 B.n296 71.676
R1268 B.n448 B.n297 71.676
R1269 B.n444 B.n298 71.676
R1270 B.n440 B.n299 71.676
R1271 B.n436 B.n300 71.676
R1272 B.n432 B.n301 71.676
R1273 B.n427 B.n302 71.676
R1274 B.n423 B.n303 71.676
R1275 B.n419 B.n304 71.676
R1276 B.n415 B.n305 71.676
R1277 B.n411 B.n306 71.676
R1278 B.n407 B.n307 71.676
R1279 B.n403 B.n308 71.676
R1280 B.n399 B.n309 71.676
R1281 B.n395 B.n310 71.676
R1282 B.n391 B.n311 71.676
R1283 B.n387 B.n312 71.676
R1284 B.n383 B.n313 71.676
R1285 B.n379 B.n314 71.676
R1286 B.n375 B.n315 71.676
R1287 B.n371 B.n316 71.676
R1288 B.n367 B.n317 71.676
R1289 B.n363 B.n318 71.676
R1290 B.n359 B.n319 71.676
R1291 B.n355 B.n320 71.676
R1292 B.n351 B.n321 71.676
R1293 B.n347 B.n322 71.676
R1294 B.n343 B.n323 71.676
R1295 B.n339 B.n324 71.676
R1296 B.n335 B.n325 71.676
R1297 B.n507 B.n282 71.676
R1298 B.n501 B.n283 71.676
R1299 B.n497 B.n284 71.676
R1300 B.n493 B.n285 71.676
R1301 B.n489 B.n286 71.676
R1302 B.n485 B.n287 71.676
R1303 B.n481 B.n288 71.676
R1304 B.n477 B.n289 71.676
R1305 B.n473 B.n290 71.676
R1306 B.n469 B.n291 71.676
R1307 B.n465 B.n292 71.676
R1308 B.n461 B.n293 71.676
R1309 B.n457 B.n294 71.676
R1310 B.n453 B.n295 71.676
R1311 B.n449 B.n296 71.676
R1312 B.n445 B.n297 71.676
R1313 B.n441 B.n298 71.676
R1314 B.n437 B.n299 71.676
R1315 B.n433 B.n300 71.676
R1316 B.n428 B.n301 71.676
R1317 B.n424 B.n302 71.676
R1318 B.n420 B.n303 71.676
R1319 B.n416 B.n304 71.676
R1320 B.n412 B.n305 71.676
R1321 B.n408 B.n306 71.676
R1322 B.n404 B.n307 71.676
R1323 B.n400 B.n308 71.676
R1324 B.n396 B.n309 71.676
R1325 B.n392 B.n310 71.676
R1326 B.n388 B.n311 71.676
R1327 B.n384 B.n312 71.676
R1328 B.n380 B.n313 71.676
R1329 B.n376 B.n314 71.676
R1330 B.n372 B.n315 71.676
R1331 B.n368 B.n316 71.676
R1332 B.n364 B.n317 71.676
R1333 B.n360 B.n318 71.676
R1334 B.n356 B.n319 71.676
R1335 B.n352 B.n320 71.676
R1336 B.n348 B.n321 71.676
R1337 B.n344 B.n322 71.676
R1338 B.n340 B.n323 71.676
R1339 B.n336 B.n324 71.676
R1340 B.n332 B.n325 71.676
R1341 B.n614 B.n613 71.676
R1342 B.n614 B.n2 71.676
R1343 B.n81 B.n80 59.5399
R1344 B.n176 B.n78 59.5399
R1345 B.n331 B.n330 59.5399
R1346 B.n430 B.n328 59.5399
R1347 B.n513 B.n279 45.1559
R1348 B.n513 B.n275 45.1559
R1349 B.n520 B.n275 45.1559
R1350 B.n520 B.n519 45.1559
R1351 B.n526 B.n268 45.1559
R1352 B.n532 B.n268 45.1559
R1353 B.n532 B.n264 45.1559
R1354 B.n538 B.n264 45.1559
R1355 B.n545 B.n260 45.1559
R1356 B.t4 B.n256 45.1559
R1357 B.t4 B.n4 45.1559
R1358 B.n612 B.n4 45.1559
R1359 B.n612 B.n611 45.1559
R1360 B.n611 B.n610 45.1559
R1361 B.n610 B.t1 45.1559
R1362 B.n559 B.t1 45.1559
R1363 B.n603 B.n602 45.1559
R1364 B.n601 B.n14 45.1559
R1365 B.n595 B.n14 45.1559
R1366 B.n595 B.n594 45.1559
R1367 B.n594 B.n593 45.1559
R1368 B.n587 B.n24 45.1559
R1369 B.n587 B.n586 45.1559
R1370 B.n586 B.n585 45.1559
R1371 B.n585 B.n28 45.1559
R1372 B.t0 B.n256 35.8592
R1373 B.n559 B.t5 35.8592
R1374 B.n510 B.n509 28.2542
R1375 B.n333 B.n277 28.2542
R1376 B.n582 B.n581 28.2542
R1377 B.n576 B.n575 28.2542
R1378 B.n526 B.t14 26.5625
R1379 B.t2 B.n260 26.5625
R1380 B.n602 B.t3 26.5625
R1381 B.n593 B.t7 26.5625
R1382 B.n519 B.t14 18.5939
R1383 B.n538 B.t2 18.5939
R1384 B.t3 B.n601 18.5939
R1385 B.n24 B.t7 18.5939
R1386 B B.n615 18.0485
R1387 B.n80 B.n79 11.8308
R1388 B.n78 B.n77 11.8308
R1389 B.n330 B.n329 11.8308
R1390 B.n328 B.n327 11.8308
R1391 B.n511 B.n510 10.6151
R1392 B.n511 B.n273 10.6151
R1393 B.n522 B.n273 10.6151
R1394 B.n523 B.n522 10.6151
R1395 B.n524 B.n523 10.6151
R1396 B.n524 B.n266 10.6151
R1397 B.n534 B.n266 10.6151
R1398 B.n535 B.n534 10.6151
R1399 B.n536 B.n535 10.6151
R1400 B.n536 B.n258 10.6151
R1401 B.n547 B.n258 10.6151
R1402 B.n548 B.n547 10.6151
R1403 B.n549 B.n548 10.6151
R1404 B.n549 B.n0 10.6151
R1405 B.n509 B.n281 10.6151
R1406 B.n504 B.n281 10.6151
R1407 B.n504 B.n503 10.6151
R1408 B.n503 B.n502 10.6151
R1409 B.n502 B.n499 10.6151
R1410 B.n499 B.n498 10.6151
R1411 B.n498 B.n495 10.6151
R1412 B.n495 B.n494 10.6151
R1413 B.n494 B.n491 10.6151
R1414 B.n491 B.n490 10.6151
R1415 B.n490 B.n487 10.6151
R1416 B.n487 B.n486 10.6151
R1417 B.n486 B.n483 10.6151
R1418 B.n483 B.n482 10.6151
R1419 B.n482 B.n479 10.6151
R1420 B.n479 B.n478 10.6151
R1421 B.n478 B.n475 10.6151
R1422 B.n475 B.n474 10.6151
R1423 B.n474 B.n471 10.6151
R1424 B.n471 B.n470 10.6151
R1425 B.n470 B.n467 10.6151
R1426 B.n467 B.n466 10.6151
R1427 B.n466 B.n463 10.6151
R1428 B.n463 B.n462 10.6151
R1429 B.n462 B.n459 10.6151
R1430 B.n459 B.n458 10.6151
R1431 B.n458 B.n455 10.6151
R1432 B.n455 B.n454 10.6151
R1433 B.n454 B.n451 10.6151
R1434 B.n451 B.n450 10.6151
R1435 B.n450 B.n447 10.6151
R1436 B.n447 B.n446 10.6151
R1437 B.n446 B.n443 10.6151
R1438 B.n443 B.n442 10.6151
R1439 B.n442 B.n439 10.6151
R1440 B.n439 B.n438 10.6151
R1441 B.n438 B.n435 10.6151
R1442 B.n435 B.n434 10.6151
R1443 B.n434 B.n431 10.6151
R1444 B.n429 B.n426 10.6151
R1445 B.n426 B.n425 10.6151
R1446 B.n425 B.n422 10.6151
R1447 B.n422 B.n421 10.6151
R1448 B.n421 B.n418 10.6151
R1449 B.n418 B.n417 10.6151
R1450 B.n417 B.n414 10.6151
R1451 B.n414 B.n413 10.6151
R1452 B.n410 B.n409 10.6151
R1453 B.n409 B.n406 10.6151
R1454 B.n406 B.n405 10.6151
R1455 B.n405 B.n402 10.6151
R1456 B.n402 B.n401 10.6151
R1457 B.n401 B.n398 10.6151
R1458 B.n398 B.n397 10.6151
R1459 B.n397 B.n394 10.6151
R1460 B.n394 B.n393 10.6151
R1461 B.n393 B.n390 10.6151
R1462 B.n390 B.n389 10.6151
R1463 B.n389 B.n386 10.6151
R1464 B.n386 B.n385 10.6151
R1465 B.n385 B.n382 10.6151
R1466 B.n382 B.n381 10.6151
R1467 B.n381 B.n378 10.6151
R1468 B.n378 B.n377 10.6151
R1469 B.n377 B.n374 10.6151
R1470 B.n374 B.n373 10.6151
R1471 B.n373 B.n370 10.6151
R1472 B.n370 B.n369 10.6151
R1473 B.n369 B.n366 10.6151
R1474 B.n366 B.n365 10.6151
R1475 B.n365 B.n362 10.6151
R1476 B.n362 B.n361 10.6151
R1477 B.n361 B.n358 10.6151
R1478 B.n358 B.n357 10.6151
R1479 B.n357 B.n354 10.6151
R1480 B.n354 B.n353 10.6151
R1481 B.n353 B.n350 10.6151
R1482 B.n350 B.n349 10.6151
R1483 B.n349 B.n346 10.6151
R1484 B.n346 B.n345 10.6151
R1485 B.n345 B.n342 10.6151
R1486 B.n342 B.n341 10.6151
R1487 B.n341 B.n338 10.6151
R1488 B.n338 B.n337 10.6151
R1489 B.n337 B.n334 10.6151
R1490 B.n334 B.n333 10.6151
R1491 B.n515 B.n277 10.6151
R1492 B.n516 B.n515 10.6151
R1493 B.n517 B.n516 10.6151
R1494 B.n517 B.n270 10.6151
R1495 B.n528 B.n270 10.6151
R1496 B.n529 B.n528 10.6151
R1497 B.n530 B.n529 10.6151
R1498 B.n530 B.n262 10.6151
R1499 B.n540 B.n262 10.6151
R1500 B.n541 B.n540 10.6151
R1501 B.n543 B.n541 10.6151
R1502 B.n543 B.n542 10.6151
R1503 B.n542 B.n254 10.6151
R1504 B.n553 B.n254 10.6151
R1505 B.n554 B.n553 10.6151
R1506 B.n555 B.n554 10.6151
R1507 B.n556 B.n555 10.6151
R1508 B.n557 B.n556 10.6151
R1509 B.n561 B.n557 10.6151
R1510 B.n562 B.n561 10.6151
R1511 B.n563 B.n562 10.6151
R1512 B.n564 B.n563 10.6151
R1513 B.n566 B.n564 10.6151
R1514 B.n567 B.n566 10.6151
R1515 B.n568 B.n567 10.6151
R1516 B.n569 B.n568 10.6151
R1517 B.n571 B.n569 10.6151
R1518 B.n572 B.n571 10.6151
R1519 B.n573 B.n572 10.6151
R1520 B.n574 B.n573 10.6151
R1521 B.n575 B.n574 10.6151
R1522 B.n607 B.n1 10.6151
R1523 B.n607 B.n606 10.6151
R1524 B.n606 B.n605 10.6151
R1525 B.n605 B.n9 10.6151
R1526 B.n599 B.n9 10.6151
R1527 B.n599 B.n598 10.6151
R1528 B.n598 B.n597 10.6151
R1529 B.n597 B.n16 10.6151
R1530 B.n591 B.n16 10.6151
R1531 B.n591 B.n590 10.6151
R1532 B.n590 B.n589 10.6151
R1533 B.n589 B.n22 10.6151
R1534 B.n583 B.n22 10.6151
R1535 B.n583 B.n582 10.6151
R1536 B.n581 B.n30 10.6151
R1537 B.n83 B.n30 10.6151
R1538 B.n84 B.n83 10.6151
R1539 B.n87 B.n84 10.6151
R1540 B.n88 B.n87 10.6151
R1541 B.n91 B.n88 10.6151
R1542 B.n92 B.n91 10.6151
R1543 B.n95 B.n92 10.6151
R1544 B.n96 B.n95 10.6151
R1545 B.n99 B.n96 10.6151
R1546 B.n100 B.n99 10.6151
R1547 B.n103 B.n100 10.6151
R1548 B.n104 B.n103 10.6151
R1549 B.n107 B.n104 10.6151
R1550 B.n108 B.n107 10.6151
R1551 B.n111 B.n108 10.6151
R1552 B.n112 B.n111 10.6151
R1553 B.n115 B.n112 10.6151
R1554 B.n116 B.n115 10.6151
R1555 B.n119 B.n116 10.6151
R1556 B.n120 B.n119 10.6151
R1557 B.n123 B.n120 10.6151
R1558 B.n124 B.n123 10.6151
R1559 B.n127 B.n124 10.6151
R1560 B.n128 B.n127 10.6151
R1561 B.n131 B.n128 10.6151
R1562 B.n132 B.n131 10.6151
R1563 B.n135 B.n132 10.6151
R1564 B.n136 B.n135 10.6151
R1565 B.n139 B.n136 10.6151
R1566 B.n140 B.n139 10.6151
R1567 B.n143 B.n140 10.6151
R1568 B.n144 B.n143 10.6151
R1569 B.n147 B.n144 10.6151
R1570 B.n148 B.n147 10.6151
R1571 B.n151 B.n148 10.6151
R1572 B.n152 B.n151 10.6151
R1573 B.n155 B.n152 10.6151
R1574 B.n156 B.n155 10.6151
R1575 B.n160 B.n159 10.6151
R1576 B.n163 B.n160 10.6151
R1577 B.n164 B.n163 10.6151
R1578 B.n167 B.n164 10.6151
R1579 B.n168 B.n167 10.6151
R1580 B.n171 B.n168 10.6151
R1581 B.n172 B.n171 10.6151
R1582 B.n175 B.n172 10.6151
R1583 B.n180 B.n177 10.6151
R1584 B.n181 B.n180 10.6151
R1585 B.n184 B.n181 10.6151
R1586 B.n185 B.n184 10.6151
R1587 B.n188 B.n185 10.6151
R1588 B.n189 B.n188 10.6151
R1589 B.n192 B.n189 10.6151
R1590 B.n193 B.n192 10.6151
R1591 B.n196 B.n193 10.6151
R1592 B.n197 B.n196 10.6151
R1593 B.n200 B.n197 10.6151
R1594 B.n201 B.n200 10.6151
R1595 B.n204 B.n201 10.6151
R1596 B.n205 B.n204 10.6151
R1597 B.n208 B.n205 10.6151
R1598 B.n209 B.n208 10.6151
R1599 B.n212 B.n209 10.6151
R1600 B.n213 B.n212 10.6151
R1601 B.n216 B.n213 10.6151
R1602 B.n217 B.n216 10.6151
R1603 B.n220 B.n217 10.6151
R1604 B.n221 B.n220 10.6151
R1605 B.n224 B.n221 10.6151
R1606 B.n225 B.n224 10.6151
R1607 B.n228 B.n225 10.6151
R1608 B.n229 B.n228 10.6151
R1609 B.n232 B.n229 10.6151
R1610 B.n233 B.n232 10.6151
R1611 B.n236 B.n233 10.6151
R1612 B.n237 B.n236 10.6151
R1613 B.n240 B.n237 10.6151
R1614 B.n241 B.n240 10.6151
R1615 B.n244 B.n241 10.6151
R1616 B.n245 B.n244 10.6151
R1617 B.n248 B.n245 10.6151
R1618 B.n249 B.n248 10.6151
R1619 B.n252 B.n249 10.6151
R1620 B.n253 B.n252 10.6151
R1621 B.n576 B.n253 10.6151
R1622 B.n545 B.t0 9.29721
R1623 B.n603 B.t5 9.29721
R1624 B.n615 B.n0 8.11757
R1625 B.n615 B.n1 8.11757
R1626 B.n430 B.n429 6.5566
R1627 B.n413 B.n331 6.5566
R1628 B.n159 B.n81 6.5566
R1629 B.n176 B.n175 6.5566
R1630 B.n431 B.n430 4.05904
R1631 B.n410 B.n331 4.05904
R1632 B.n156 B.n81 4.05904
R1633 B.n177 B.n176 4.05904
R1634 VP.n7 VP.t5 1137.08
R1635 VP.n5 VP.t2 1137.08
R1636 VP.n0 VP.t1 1137.08
R1637 VP.n2 VP.t4 1137.08
R1638 VP.n6 VP.t3 1084.5
R1639 VP.n1 VP.t0 1084.5
R1640 VP.n3 VP.n0 161.489
R1641 VP.n8 VP.n7 161.3
R1642 VP.n3 VP.n2 161.3
R1643 VP.n5 VP.n4 161.3
R1644 VP.n4 VP.n3 39.1634
R1645 VP.n6 VP.n5 36.5157
R1646 VP.n7 VP.n6 36.5157
R1647 VP.n1 VP.n0 36.5157
R1648 VP.n2 VP.n1 36.5157
R1649 VP.n8 VP.n4 0.189894
R1650 VP VP.n8 0.0516364
R1651 VDD1.n56 VDD1.n0 289.615
R1652 VDD1.n117 VDD1.n61 289.615
R1653 VDD1.n57 VDD1.n56 185
R1654 VDD1.n55 VDD1.n54 185
R1655 VDD1.n4 VDD1.n3 185
R1656 VDD1.n49 VDD1.n48 185
R1657 VDD1.n47 VDD1.n46 185
R1658 VDD1.n8 VDD1.n7 185
R1659 VDD1.n12 VDD1.n10 185
R1660 VDD1.n41 VDD1.n40 185
R1661 VDD1.n39 VDD1.n38 185
R1662 VDD1.n14 VDD1.n13 185
R1663 VDD1.n33 VDD1.n32 185
R1664 VDD1.n31 VDD1.n30 185
R1665 VDD1.n18 VDD1.n17 185
R1666 VDD1.n25 VDD1.n24 185
R1667 VDD1.n23 VDD1.n22 185
R1668 VDD1.n82 VDD1.n81 185
R1669 VDD1.n84 VDD1.n83 185
R1670 VDD1.n77 VDD1.n76 185
R1671 VDD1.n90 VDD1.n89 185
R1672 VDD1.n92 VDD1.n91 185
R1673 VDD1.n73 VDD1.n72 185
R1674 VDD1.n99 VDD1.n98 185
R1675 VDD1.n100 VDD1.n71 185
R1676 VDD1.n102 VDD1.n101 185
R1677 VDD1.n69 VDD1.n68 185
R1678 VDD1.n108 VDD1.n107 185
R1679 VDD1.n110 VDD1.n109 185
R1680 VDD1.n65 VDD1.n64 185
R1681 VDD1.n116 VDD1.n115 185
R1682 VDD1.n118 VDD1.n117 185
R1683 VDD1.n21 VDD1.t4 149.524
R1684 VDD1.n80 VDD1.t3 149.524
R1685 VDD1.n56 VDD1.n55 104.615
R1686 VDD1.n55 VDD1.n3 104.615
R1687 VDD1.n48 VDD1.n3 104.615
R1688 VDD1.n48 VDD1.n47 104.615
R1689 VDD1.n47 VDD1.n7 104.615
R1690 VDD1.n12 VDD1.n7 104.615
R1691 VDD1.n40 VDD1.n12 104.615
R1692 VDD1.n40 VDD1.n39 104.615
R1693 VDD1.n39 VDD1.n13 104.615
R1694 VDD1.n32 VDD1.n13 104.615
R1695 VDD1.n32 VDD1.n31 104.615
R1696 VDD1.n31 VDD1.n17 104.615
R1697 VDD1.n24 VDD1.n17 104.615
R1698 VDD1.n24 VDD1.n23 104.615
R1699 VDD1.n83 VDD1.n82 104.615
R1700 VDD1.n83 VDD1.n76 104.615
R1701 VDD1.n90 VDD1.n76 104.615
R1702 VDD1.n91 VDD1.n90 104.615
R1703 VDD1.n91 VDD1.n72 104.615
R1704 VDD1.n99 VDD1.n72 104.615
R1705 VDD1.n100 VDD1.n99 104.615
R1706 VDD1.n101 VDD1.n100 104.615
R1707 VDD1.n101 VDD1.n68 104.615
R1708 VDD1.n108 VDD1.n68 104.615
R1709 VDD1.n109 VDD1.n108 104.615
R1710 VDD1.n109 VDD1.n64 104.615
R1711 VDD1.n116 VDD1.n64 104.615
R1712 VDD1.n117 VDD1.n116 104.615
R1713 VDD1.n123 VDD1.n122 60.0325
R1714 VDD1.n125 VDD1.n124 59.9564
R1715 VDD1.n23 VDD1.t4 52.3082
R1716 VDD1.n82 VDD1.t3 52.3082
R1717 VDD1 VDD1.n60 47.1834
R1718 VDD1.n123 VDD1.n121 47.0699
R1719 VDD1.n125 VDD1.n123 36.0031
R1720 VDD1.n10 VDD1.n8 13.1884
R1721 VDD1.n102 VDD1.n69 13.1884
R1722 VDD1.n46 VDD1.n45 12.8005
R1723 VDD1.n42 VDD1.n41 12.8005
R1724 VDD1.n103 VDD1.n71 12.8005
R1725 VDD1.n107 VDD1.n106 12.8005
R1726 VDD1.n49 VDD1.n6 12.0247
R1727 VDD1.n38 VDD1.n11 12.0247
R1728 VDD1.n98 VDD1.n97 12.0247
R1729 VDD1.n110 VDD1.n67 12.0247
R1730 VDD1.n50 VDD1.n4 11.249
R1731 VDD1.n37 VDD1.n14 11.249
R1732 VDD1.n96 VDD1.n73 11.249
R1733 VDD1.n111 VDD1.n65 11.249
R1734 VDD1.n54 VDD1.n53 10.4732
R1735 VDD1.n34 VDD1.n33 10.4732
R1736 VDD1.n93 VDD1.n92 10.4732
R1737 VDD1.n115 VDD1.n114 10.4732
R1738 VDD1.n22 VDD1.n21 10.2747
R1739 VDD1.n81 VDD1.n80 10.2747
R1740 VDD1.n57 VDD1.n2 9.69747
R1741 VDD1.n30 VDD1.n16 9.69747
R1742 VDD1.n89 VDD1.n75 9.69747
R1743 VDD1.n118 VDD1.n63 9.69747
R1744 VDD1.n60 VDD1.n59 9.45567
R1745 VDD1.n121 VDD1.n120 9.45567
R1746 VDD1.n20 VDD1.n19 9.3005
R1747 VDD1.n27 VDD1.n26 9.3005
R1748 VDD1.n29 VDD1.n28 9.3005
R1749 VDD1.n16 VDD1.n15 9.3005
R1750 VDD1.n35 VDD1.n34 9.3005
R1751 VDD1.n37 VDD1.n36 9.3005
R1752 VDD1.n11 VDD1.n9 9.3005
R1753 VDD1.n43 VDD1.n42 9.3005
R1754 VDD1.n59 VDD1.n58 9.3005
R1755 VDD1.n2 VDD1.n1 9.3005
R1756 VDD1.n53 VDD1.n52 9.3005
R1757 VDD1.n51 VDD1.n50 9.3005
R1758 VDD1.n6 VDD1.n5 9.3005
R1759 VDD1.n45 VDD1.n44 9.3005
R1760 VDD1.n120 VDD1.n119 9.3005
R1761 VDD1.n63 VDD1.n62 9.3005
R1762 VDD1.n114 VDD1.n113 9.3005
R1763 VDD1.n112 VDD1.n111 9.3005
R1764 VDD1.n67 VDD1.n66 9.3005
R1765 VDD1.n106 VDD1.n105 9.3005
R1766 VDD1.n79 VDD1.n78 9.3005
R1767 VDD1.n86 VDD1.n85 9.3005
R1768 VDD1.n88 VDD1.n87 9.3005
R1769 VDD1.n75 VDD1.n74 9.3005
R1770 VDD1.n94 VDD1.n93 9.3005
R1771 VDD1.n96 VDD1.n95 9.3005
R1772 VDD1.n97 VDD1.n70 9.3005
R1773 VDD1.n104 VDD1.n103 9.3005
R1774 VDD1.n58 VDD1.n0 8.92171
R1775 VDD1.n29 VDD1.n18 8.92171
R1776 VDD1.n88 VDD1.n77 8.92171
R1777 VDD1.n119 VDD1.n61 8.92171
R1778 VDD1.n26 VDD1.n25 8.14595
R1779 VDD1.n85 VDD1.n84 8.14595
R1780 VDD1.n22 VDD1.n20 7.3702
R1781 VDD1.n81 VDD1.n79 7.3702
R1782 VDD1.n25 VDD1.n20 5.81868
R1783 VDD1.n84 VDD1.n79 5.81868
R1784 VDD1.n60 VDD1.n0 5.04292
R1785 VDD1.n26 VDD1.n18 5.04292
R1786 VDD1.n85 VDD1.n77 5.04292
R1787 VDD1.n121 VDD1.n61 5.04292
R1788 VDD1.n58 VDD1.n57 4.26717
R1789 VDD1.n30 VDD1.n29 4.26717
R1790 VDD1.n89 VDD1.n88 4.26717
R1791 VDD1.n119 VDD1.n118 4.26717
R1792 VDD1.n54 VDD1.n2 3.49141
R1793 VDD1.n33 VDD1.n16 3.49141
R1794 VDD1.n92 VDD1.n75 3.49141
R1795 VDD1.n115 VDD1.n63 3.49141
R1796 VDD1.n21 VDD1.n19 2.84303
R1797 VDD1.n80 VDD1.n78 2.84303
R1798 VDD1.n53 VDD1.n4 2.71565
R1799 VDD1.n34 VDD1.n14 2.71565
R1800 VDD1.n93 VDD1.n73 2.71565
R1801 VDD1.n114 VDD1.n65 2.71565
R1802 VDD1.n50 VDD1.n49 1.93989
R1803 VDD1.n38 VDD1.n37 1.93989
R1804 VDD1.n98 VDD1.n96 1.93989
R1805 VDD1.n111 VDD1.n110 1.93989
R1806 VDD1.n124 VDD1.t5 1.75426
R1807 VDD1.n124 VDD1.t1 1.75426
R1808 VDD1.n122 VDD1.t2 1.75426
R1809 VDD1.n122 VDD1.t0 1.75426
R1810 VDD1.n46 VDD1.n6 1.16414
R1811 VDD1.n41 VDD1.n11 1.16414
R1812 VDD1.n97 VDD1.n71 1.16414
R1813 VDD1.n107 VDD1.n67 1.16414
R1814 VDD1.n45 VDD1.n8 0.388379
R1815 VDD1.n42 VDD1.n10 0.388379
R1816 VDD1.n103 VDD1.n102 0.388379
R1817 VDD1.n106 VDD1.n69 0.388379
R1818 VDD1.n59 VDD1.n1 0.155672
R1819 VDD1.n52 VDD1.n1 0.155672
R1820 VDD1.n52 VDD1.n51 0.155672
R1821 VDD1.n51 VDD1.n5 0.155672
R1822 VDD1.n44 VDD1.n5 0.155672
R1823 VDD1.n44 VDD1.n43 0.155672
R1824 VDD1.n43 VDD1.n9 0.155672
R1825 VDD1.n36 VDD1.n9 0.155672
R1826 VDD1.n36 VDD1.n35 0.155672
R1827 VDD1.n35 VDD1.n15 0.155672
R1828 VDD1.n28 VDD1.n15 0.155672
R1829 VDD1.n28 VDD1.n27 0.155672
R1830 VDD1.n27 VDD1.n19 0.155672
R1831 VDD1.n86 VDD1.n78 0.155672
R1832 VDD1.n87 VDD1.n86 0.155672
R1833 VDD1.n87 VDD1.n74 0.155672
R1834 VDD1.n94 VDD1.n74 0.155672
R1835 VDD1.n95 VDD1.n94 0.155672
R1836 VDD1.n95 VDD1.n70 0.155672
R1837 VDD1.n104 VDD1.n70 0.155672
R1838 VDD1.n105 VDD1.n104 0.155672
R1839 VDD1.n105 VDD1.n66 0.155672
R1840 VDD1.n112 VDD1.n66 0.155672
R1841 VDD1.n113 VDD1.n112 0.155672
R1842 VDD1.n113 VDD1.n62 0.155672
R1843 VDD1.n120 VDD1.n62 0.155672
R1844 VDD1 VDD1.n125 0.0737759
C0 VDD1 VTAIL 13.563201f
C1 VDD2 VP 0.261984f
C2 VN VTAIL 2.02568f
C3 VDD1 VDD2 0.562509f
C4 VDD1 VP 2.58119f
C5 VDD2 VN 2.47146f
C6 VN VP 4.53818f
C7 VDD2 VTAIL 13.593f
C8 VTAIL VP 2.04041f
C9 VDD1 VN 0.147417f
C10 VDD2 B 4.066954f
C11 VDD1 B 4.006949f
C12 VTAIL B 5.745026f
C13 VN B 6.688529f
C14 VP B 4.447804f
C15 VDD1.n0 B 0.037035f
C16 VDD1.n1 B 0.028393f
C17 VDD1.n2 B 0.015257f
C18 VDD1.n3 B 0.036062f
C19 VDD1.n4 B 0.016154f
C20 VDD1.n5 B 0.028393f
C21 VDD1.n6 B 0.015257f
C22 VDD1.n7 B 0.036062f
C23 VDD1.n8 B 0.015706f
C24 VDD1.n9 B 0.028393f
C25 VDD1.n10 B 0.015706f
C26 VDD1.n11 B 0.015257f
C27 VDD1.n12 B 0.036062f
C28 VDD1.n13 B 0.036062f
C29 VDD1.n14 B 0.016154f
C30 VDD1.n15 B 0.028393f
C31 VDD1.n16 B 0.015257f
C32 VDD1.n17 B 0.036062f
C33 VDD1.n18 B 0.016154f
C34 VDD1.n19 B 1.3427f
C35 VDD1.n20 B 0.015257f
C36 VDD1.t4 B 0.060798f
C37 VDD1.n21 B 0.196969f
C38 VDD1.n22 B 0.025493f
C39 VDD1.n23 B 0.027046f
C40 VDD1.n24 B 0.036062f
C41 VDD1.n25 B 0.016154f
C42 VDD1.n26 B 0.015257f
C43 VDD1.n27 B 0.028393f
C44 VDD1.n28 B 0.028393f
C45 VDD1.n29 B 0.015257f
C46 VDD1.n30 B 0.016154f
C47 VDD1.n31 B 0.036062f
C48 VDD1.n32 B 0.036062f
C49 VDD1.n33 B 0.016154f
C50 VDD1.n34 B 0.015257f
C51 VDD1.n35 B 0.028393f
C52 VDD1.n36 B 0.028393f
C53 VDD1.n37 B 0.015257f
C54 VDD1.n38 B 0.016154f
C55 VDD1.n39 B 0.036062f
C56 VDD1.n40 B 0.036062f
C57 VDD1.n41 B 0.016154f
C58 VDD1.n42 B 0.015257f
C59 VDD1.n43 B 0.028393f
C60 VDD1.n44 B 0.028393f
C61 VDD1.n45 B 0.015257f
C62 VDD1.n46 B 0.016154f
C63 VDD1.n47 B 0.036062f
C64 VDD1.n48 B 0.036062f
C65 VDD1.n49 B 0.016154f
C66 VDD1.n50 B 0.015257f
C67 VDD1.n51 B 0.028393f
C68 VDD1.n52 B 0.028393f
C69 VDD1.n53 B 0.015257f
C70 VDD1.n54 B 0.016154f
C71 VDD1.n55 B 0.036062f
C72 VDD1.n56 B 0.072987f
C73 VDD1.n57 B 0.016154f
C74 VDD1.n58 B 0.015257f
C75 VDD1.n59 B 0.061362f
C76 VDD1.n60 B 0.060721f
C77 VDD1.n61 B 0.037035f
C78 VDD1.n62 B 0.028393f
C79 VDD1.n63 B 0.015257f
C80 VDD1.n64 B 0.036062f
C81 VDD1.n65 B 0.016154f
C82 VDD1.n66 B 0.028393f
C83 VDD1.n67 B 0.015257f
C84 VDD1.n68 B 0.036062f
C85 VDD1.n69 B 0.015706f
C86 VDD1.n70 B 0.028393f
C87 VDD1.n71 B 0.016154f
C88 VDD1.n72 B 0.036062f
C89 VDD1.n73 B 0.016154f
C90 VDD1.n74 B 0.028393f
C91 VDD1.n75 B 0.015257f
C92 VDD1.n76 B 0.036062f
C93 VDD1.n77 B 0.016154f
C94 VDD1.n78 B 1.3427f
C95 VDD1.n79 B 0.015257f
C96 VDD1.t3 B 0.060798f
C97 VDD1.n80 B 0.196969f
C98 VDD1.n81 B 0.025493f
C99 VDD1.n82 B 0.027046f
C100 VDD1.n83 B 0.036062f
C101 VDD1.n84 B 0.016154f
C102 VDD1.n85 B 0.015257f
C103 VDD1.n86 B 0.028393f
C104 VDD1.n87 B 0.028393f
C105 VDD1.n88 B 0.015257f
C106 VDD1.n89 B 0.016154f
C107 VDD1.n90 B 0.036062f
C108 VDD1.n91 B 0.036062f
C109 VDD1.n92 B 0.016154f
C110 VDD1.n93 B 0.015257f
C111 VDD1.n94 B 0.028393f
C112 VDD1.n95 B 0.028393f
C113 VDD1.n96 B 0.015257f
C114 VDD1.n97 B 0.015257f
C115 VDD1.n98 B 0.016154f
C116 VDD1.n99 B 0.036062f
C117 VDD1.n100 B 0.036062f
C118 VDD1.n101 B 0.036062f
C119 VDD1.n102 B 0.015706f
C120 VDD1.n103 B 0.015257f
C121 VDD1.n104 B 0.028393f
C122 VDD1.n105 B 0.028393f
C123 VDD1.n106 B 0.015257f
C124 VDD1.n107 B 0.016154f
C125 VDD1.n108 B 0.036062f
C126 VDD1.n109 B 0.036062f
C127 VDD1.n110 B 0.016154f
C128 VDD1.n111 B 0.015257f
C129 VDD1.n112 B 0.028393f
C130 VDD1.n113 B 0.028393f
C131 VDD1.n114 B 0.015257f
C132 VDD1.n115 B 0.016154f
C133 VDD1.n116 B 0.036062f
C134 VDD1.n117 B 0.072987f
C135 VDD1.n118 B 0.016154f
C136 VDD1.n119 B 0.015257f
C137 VDD1.n120 B 0.061362f
C138 VDD1.n121 B 0.060436f
C139 VDD1.t2 B 0.253311f
C140 VDD1.t0 B 0.253311f
C141 VDD1.n122 B 2.24624f
C142 VDD1.n123 B 1.92325f
C143 VDD1.t5 B 0.253311f
C144 VDD1.t1 B 0.253311f
C145 VDD1.n124 B 2.24584f
C146 VDD1.n125 B 2.36389f
C147 VP.t1 B 0.538368f
C148 VP.n0 B 0.231678f
C149 VP.t0 B 0.528284f
C150 VP.n1 B 0.212961f
C151 VP.t4 B 0.538368f
C152 VP.n2 B 0.231587f
C153 VP.n3 B 2.24163f
C154 VP.n4 B 2.21866f
C155 VP.t3 B 0.528284f
C156 VP.t2 B 0.538368f
C157 VP.n5 B 0.231587f
C158 VP.n6 B 0.212961f
C159 VP.t5 B 0.538368f
C160 VP.n7 B 0.231587f
C161 VP.n8 B 0.045793f
C162 VDD2.n0 B 0.037046f
C163 VDD2.n1 B 0.028401f
C164 VDD2.n2 B 0.015262f
C165 VDD2.n3 B 0.036073f
C166 VDD2.n4 B 0.016159f
C167 VDD2.n5 B 0.028401f
C168 VDD2.n6 B 0.015262f
C169 VDD2.n7 B 0.036073f
C170 VDD2.n8 B 0.01571f
C171 VDD2.n9 B 0.028401f
C172 VDD2.n10 B 0.016159f
C173 VDD2.n11 B 0.036073f
C174 VDD2.n12 B 0.016159f
C175 VDD2.n13 B 0.028401f
C176 VDD2.n14 B 0.015262f
C177 VDD2.n15 B 0.036073f
C178 VDD2.n16 B 0.016159f
C179 VDD2.n17 B 1.3431f
C180 VDD2.n18 B 0.015262f
C181 VDD2.t5 B 0.060816f
C182 VDD2.n19 B 0.197028f
C183 VDD2.n20 B 0.025501f
C184 VDD2.n21 B 0.027055f
C185 VDD2.n22 B 0.036073f
C186 VDD2.n23 B 0.016159f
C187 VDD2.n24 B 0.015262f
C188 VDD2.n25 B 0.028401f
C189 VDD2.n26 B 0.028401f
C190 VDD2.n27 B 0.015262f
C191 VDD2.n28 B 0.016159f
C192 VDD2.n29 B 0.036073f
C193 VDD2.n30 B 0.036073f
C194 VDD2.n31 B 0.016159f
C195 VDD2.n32 B 0.015262f
C196 VDD2.n33 B 0.028401f
C197 VDD2.n34 B 0.028401f
C198 VDD2.n35 B 0.015262f
C199 VDD2.n36 B 0.015262f
C200 VDD2.n37 B 0.016159f
C201 VDD2.n38 B 0.036073f
C202 VDD2.n39 B 0.036073f
C203 VDD2.n40 B 0.036073f
C204 VDD2.n41 B 0.01571f
C205 VDD2.n42 B 0.015262f
C206 VDD2.n43 B 0.028401f
C207 VDD2.n44 B 0.028401f
C208 VDD2.n45 B 0.015262f
C209 VDD2.n46 B 0.016159f
C210 VDD2.n47 B 0.036073f
C211 VDD2.n48 B 0.036073f
C212 VDD2.n49 B 0.016159f
C213 VDD2.n50 B 0.015262f
C214 VDD2.n51 B 0.028401f
C215 VDD2.n52 B 0.028401f
C216 VDD2.n53 B 0.015262f
C217 VDD2.n54 B 0.016159f
C218 VDD2.n55 B 0.036073f
C219 VDD2.n56 B 0.073009f
C220 VDD2.n57 B 0.016159f
C221 VDD2.n58 B 0.015262f
C222 VDD2.n59 B 0.06138f
C223 VDD2.n60 B 0.060455f
C224 VDD2.t3 B 0.253388f
C225 VDD2.t0 B 0.253388f
C226 VDD2.n61 B 2.24691f
C227 VDD2.n62 B 1.84726f
C228 VDD2.n63 B 0.037046f
C229 VDD2.n64 B 0.028401f
C230 VDD2.n65 B 0.015262f
C231 VDD2.n66 B 0.036073f
C232 VDD2.n67 B 0.016159f
C233 VDD2.n68 B 0.028401f
C234 VDD2.n69 B 0.015262f
C235 VDD2.n70 B 0.036073f
C236 VDD2.n71 B 0.01571f
C237 VDD2.n72 B 0.028401f
C238 VDD2.n73 B 0.01571f
C239 VDD2.n74 B 0.015262f
C240 VDD2.n75 B 0.036073f
C241 VDD2.n76 B 0.036073f
C242 VDD2.n77 B 0.016159f
C243 VDD2.n78 B 0.028401f
C244 VDD2.n79 B 0.015262f
C245 VDD2.n80 B 0.036073f
C246 VDD2.n81 B 0.016159f
C247 VDD2.n82 B 1.3431f
C248 VDD2.n83 B 0.015262f
C249 VDD2.t1 B 0.060816f
C250 VDD2.n84 B 0.197028f
C251 VDD2.n85 B 0.025501f
C252 VDD2.n86 B 0.027055f
C253 VDD2.n87 B 0.036073f
C254 VDD2.n88 B 0.016159f
C255 VDD2.n89 B 0.015262f
C256 VDD2.n90 B 0.028401f
C257 VDD2.n91 B 0.028401f
C258 VDD2.n92 B 0.015262f
C259 VDD2.n93 B 0.016159f
C260 VDD2.n94 B 0.036073f
C261 VDD2.n95 B 0.036073f
C262 VDD2.n96 B 0.016159f
C263 VDD2.n97 B 0.015262f
C264 VDD2.n98 B 0.028401f
C265 VDD2.n99 B 0.028401f
C266 VDD2.n100 B 0.015262f
C267 VDD2.n101 B 0.016159f
C268 VDD2.n102 B 0.036073f
C269 VDD2.n103 B 0.036073f
C270 VDD2.n104 B 0.016159f
C271 VDD2.n105 B 0.015262f
C272 VDD2.n106 B 0.028401f
C273 VDD2.n107 B 0.028401f
C274 VDD2.n108 B 0.015262f
C275 VDD2.n109 B 0.016159f
C276 VDD2.n110 B 0.036073f
C277 VDD2.n111 B 0.036073f
C278 VDD2.n112 B 0.016159f
C279 VDD2.n113 B 0.015262f
C280 VDD2.n114 B 0.028401f
C281 VDD2.n115 B 0.028401f
C282 VDD2.n116 B 0.015262f
C283 VDD2.n117 B 0.016159f
C284 VDD2.n118 B 0.036073f
C285 VDD2.n119 B 0.073009f
C286 VDD2.n120 B 0.016159f
C287 VDD2.n121 B 0.015262f
C288 VDD2.n122 B 0.06138f
C289 VDD2.n123 B 0.059841f
C290 VDD2.n124 B 2.1269f
C291 VDD2.t4 B 0.253388f
C292 VDD2.t2 B 0.253388f
C293 VDD2.n125 B 2.24689f
C294 VTAIL.t5 B 0.260083f
C295 VTAIL.t7 B 0.260083f
C296 VTAIL.n0 B 2.21436f
C297 VTAIL.n1 B 0.381571f
C298 VTAIL.n2 B 0.038025f
C299 VTAIL.n3 B 0.029152f
C300 VTAIL.n4 B 0.015665f
C301 VTAIL.n5 B 0.037026f
C302 VTAIL.n6 B 0.016586f
C303 VTAIL.n7 B 0.029152f
C304 VTAIL.n8 B 0.015665f
C305 VTAIL.n9 B 0.037026f
C306 VTAIL.n10 B 0.016126f
C307 VTAIL.n11 B 0.029152f
C308 VTAIL.n12 B 0.016586f
C309 VTAIL.n13 B 0.037026f
C310 VTAIL.n14 B 0.016586f
C311 VTAIL.n15 B 0.029152f
C312 VTAIL.n16 B 0.015665f
C313 VTAIL.n17 B 0.037026f
C314 VTAIL.n18 B 0.016586f
C315 VTAIL.n19 B 1.3786f
C316 VTAIL.n20 B 0.015665f
C317 VTAIL.t10 B 0.062423f
C318 VTAIL.n21 B 0.202235f
C319 VTAIL.n22 B 0.026175f
C320 VTAIL.n23 B 0.02777f
C321 VTAIL.n24 B 0.037026f
C322 VTAIL.n25 B 0.016586f
C323 VTAIL.n26 B 0.015665f
C324 VTAIL.n27 B 0.029152f
C325 VTAIL.n28 B 0.029152f
C326 VTAIL.n29 B 0.015665f
C327 VTAIL.n30 B 0.016586f
C328 VTAIL.n31 B 0.037026f
C329 VTAIL.n32 B 0.037026f
C330 VTAIL.n33 B 0.016586f
C331 VTAIL.n34 B 0.015665f
C332 VTAIL.n35 B 0.029152f
C333 VTAIL.n36 B 0.029152f
C334 VTAIL.n37 B 0.015665f
C335 VTAIL.n38 B 0.015665f
C336 VTAIL.n39 B 0.016586f
C337 VTAIL.n40 B 0.037026f
C338 VTAIL.n41 B 0.037026f
C339 VTAIL.n42 B 0.037026f
C340 VTAIL.n43 B 0.016126f
C341 VTAIL.n44 B 0.015665f
C342 VTAIL.n45 B 0.029152f
C343 VTAIL.n46 B 0.029152f
C344 VTAIL.n47 B 0.015665f
C345 VTAIL.n48 B 0.016586f
C346 VTAIL.n49 B 0.037026f
C347 VTAIL.n50 B 0.037026f
C348 VTAIL.n51 B 0.016586f
C349 VTAIL.n52 B 0.015665f
C350 VTAIL.n53 B 0.029152f
C351 VTAIL.n54 B 0.029152f
C352 VTAIL.n55 B 0.015665f
C353 VTAIL.n56 B 0.016586f
C354 VTAIL.n57 B 0.037026f
C355 VTAIL.n58 B 0.074938f
C356 VTAIL.n59 B 0.016586f
C357 VTAIL.n60 B 0.015665f
C358 VTAIL.n61 B 0.063002f
C359 VTAIL.n62 B 0.041256f
C360 VTAIL.n63 B 0.140656f
C361 VTAIL.t2 B 0.260083f
C362 VTAIL.t0 B 0.260083f
C363 VTAIL.n64 B 2.21436f
C364 VTAIL.n65 B 1.75334f
C365 VTAIL.t8 B 0.260083f
C366 VTAIL.t3 B 0.260083f
C367 VTAIL.n66 B 2.21438f
C368 VTAIL.n67 B 1.75332f
C369 VTAIL.n68 B 0.038025f
C370 VTAIL.n69 B 0.029152f
C371 VTAIL.n70 B 0.015665f
C372 VTAIL.n71 B 0.037026f
C373 VTAIL.n72 B 0.016586f
C374 VTAIL.n73 B 0.029152f
C375 VTAIL.n74 B 0.015665f
C376 VTAIL.n75 B 0.037026f
C377 VTAIL.n76 B 0.016126f
C378 VTAIL.n77 B 0.029152f
C379 VTAIL.n78 B 0.016126f
C380 VTAIL.n79 B 0.015665f
C381 VTAIL.n80 B 0.037026f
C382 VTAIL.n81 B 0.037026f
C383 VTAIL.n82 B 0.016586f
C384 VTAIL.n83 B 0.029152f
C385 VTAIL.n84 B 0.015665f
C386 VTAIL.n85 B 0.037026f
C387 VTAIL.n86 B 0.016586f
C388 VTAIL.n87 B 1.3786f
C389 VTAIL.n88 B 0.015665f
C390 VTAIL.t6 B 0.062423f
C391 VTAIL.n89 B 0.202235f
C392 VTAIL.n90 B 0.026175f
C393 VTAIL.n91 B 0.02777f
C394 VTAIL.n92 B 0.037026f
C395 VTAIL.n93 B 0.016586f
C396 VTAIL.n94 B 0.015665f
C397 VTAIL.n95 B 0.029152f
C398 VTAIL.n96 B 0.029152f
C399 VTAIL.n97 B 0.015665f
C400 VTAIL.n98 B 0.016586f
C401 VTAIL.n99 B 0.037026f
C402 VTAIL.n100 B 0.037026f
C403 VTAIL.n101 B 0.016586f
C404 VTAIL.n102 B 0.015665f
C405 VTAIL.n103 B 0.029152f
C406 VTAIL.n104 B 0.029152f
C407 VTAIL.n105 B 0.015665f
C408 VTAIL.n106 B 0.016586f
C409 VTAIL.n107 B 0.037026f
C410 VTAIL.n108 B 0.037026f
C411 VTAIL.n109 B 0.016586f
C412 VTAIL.n110 B 0.015665f
C413 VTAIL.n111 B 0.029152f
C414 VTAIL.n112 B 0.029152f
C415 VTAIL.n113 B 0.015665f
C416 VTAIL.n114 B 0.016586f
C417 VTAIL.n115 B 0.037026f
C418 VTAIL.n116 B 0.037026f
C419 VTAIL.n117 B 0.016586f
C420 VTAIL.n118 B 0.015665f
C421 VTAIL.n119 B 0.029152f
C422 VTAIL.n120 B 0.029152f
C423 VTAIL.n121 B 0.015665f
C424 VTAIL.n122 B 0.016586f
C425 VTAIL.n123 B 0.037026f
C426 VTAIL.n124 B 0.074938f
C427 VTAIL.n125 B 0.016586f
C428 VTAIL.n126 B 0.015665f
C429 VTAIL.n127 B 0.063002f
C430 VTAIL.n128 B 0.041256f
C431 VTAIL.n129 B 0.140656f
C432 VTAIL.t1 B 0.260083f
C433 VTAIL.t9 B 0.260083f
C434 VTAIL.n130 B 2.21438f
C435 VTAIL.n131 B 0.413138f
C436 VTAIL.n132 B 0.038025f
C437 VTAIL.n133 B 0.029152f
C438 VTAIL.n134 B 0.015665f
C439 VTAIL.n135 B 0.037026f
C440 VTAIL.n136 B 0.016586f
C441 VTAIL.n137 B 0.029152f
C442 VTAIL.n138 B 0.015665f
C443 VTAIL.n139 B 0.037026f
C444 VTAIL.n140 B 0.016126f
C445 VTAIL.n141 B 0.029152f
C446 VTAIL.n142 B 0.016126f
C447 VTAIL.n143 B 0.015665f
C448 VTAIL.n144 B 0.037026f
C449 VTAIL.n145 B 0.037026f
C450 VTAIL.n146 B 0.016586f
C451 VTAIL.n147 B 0.029152f
C452 VTAIL.n148 B 0.015665f
C453 VTAIL.n149 B 0.037026f
C454 VTAIL.n150 B 0.016586f
C455 VTAIL.n151 B 1.3786f
C456 VTAIL.n152 B 0.015665f
C457 VTAIL.t11 B 0.062423f
C458 VTAIL.n153 B 0.202235f
C459 VTAIL.n154 B 0.026175f
C460 VTAIL.n155 B 0.02777f
C461 VTAIL.n156 B 0.037026f
C462 VTAIL.n157 B 0.016586f
C463 VTAIL.n158 B 0.015665f
C464 VTAIL.n159 B 0.029152f
C465 VTAIL.n160 B 0.029152f
C466 VTAIL.n161 B 0.015665f
C467 VTAIL.n162 B 0.016586f
C468 VTAIL.n163 B 0.037026f
C469 VTAIL.n164 B 0.037026f
C470 VTAIL.n165 B 0.016586f
C471 VTAIL.n166 B 0.015665f
C472 VTAIL.n167 B 0.029152f
C473 VTAIL.n168 B 0.029152f
C474 VTAIL.n169 B 0.015665f
C475 VTAIL.n170 B 0.016586f
C476 VTAIL.n171 B 0.037026f
C477 VTAIL.n172 B 0.037026f
C478 VTAIL.n173 B 0.016586f
C479 VTAIL.n174 B 0.015665f
C480 VTAIL.n175 B 0.029152f
C481 VTAIL.n176 B 0.029152f
C482 VTAIL.n177 B 0.015665f
C483 VTAIL.n178 B 0.016586f
C484 VTAIL.n179 B 0.037026f
C485 VTAIL.n180 B 0.037026f
C486 VTAIL.n181 B 0.016586f
C487 VTAIL.n182 B 0.015665f
C488 VTAIL.n183 B 0.029152f
C489 VTAIL.n184 B 0.029152f
C490 VTAIL.n185 B 0.015665f
C491 VTAIL.n186 B 0.016586f
C492 VTAIL.n187 B 0.037026f
C493 VTAIL.n188 B 0.074938f
C494 VTAIL.n189 B 0.016586f
C495 VTAIL.n190 B 0.015665f
C496 VTAIL.n191 B 0.063002f
C497 VTAIL.n192 B 0.041256f
C498 VTAIL.n193 B 1.43145f
C499 VTAIL.n194 B 0.038025f
C500 VTAIL.n195 B 0.029152f
C501 VTAIL.n196 B 0.015665f
C502 VTAIL.n197 B 0.037026f
C503 VTAIL.n198 B 0.016586f
C504 VTAIL.n199 B 0.029152f
C505 VTAIL.n200 B 0.015665f
C506 VTAIL.n201 B 0.037026f
C507 VTAIL.n202 B 0.016126f
C508 VTAIL.n203 B 0.029152f
C509 VTAIL.n204 B 0.016586f
C510 VTAIL.n205 B 0.037026f
C511 VTAIL.n206 B 0.016586f
C512 VTAIL.n207 B 0.029152f
C513 VTAIL.n208 B 0.015665f
C514 VTAIL.n209 B 0.037026f
C515 VTAIL.n210 B 0.016586f
C516 VTAIL.n211 B 1.3786f
C517 VTAIL.n212 B 0.015665f
C518 VTAIL.t4 B 0.062423f
C519 VTAIL.n213 B 0.202235f
C520 VTAIL.n214 B 0.026175f
C521 VTAIL.n215 B 0.02777f
C522 VTAIL.n216 B 0.037026f
C523 VTAIL.n217 B 0.016586f
C524 VTAIL.n218 B 0.015665f
C525 VTAIL.n219 B 0.029152f
C526 VTAIL.n220 B 0.029152f
C527 VTAIL.n221 B 0.015665f
C528 VTAIL.n222 B 0.016586f
C529 VTAIL.n223 B 0.037026f
C530 VTAIL.n224 B 0.037026f
C531 VTAIL.n225 B 0.016586f
C532 VTAIL.n226 B 0.015665f
C533 VTAIL.n227 B 0.029152f
C534 VTAIL.n228 B 0.029152f
C535 VTAIL.n229 B 0.015665f
C536 VTAIL.n230 B 0.015665f
C537 VTAIL.n231 B 0.016586f
C538 VTAIL.n232 B 0.037026f
C539 VTAIL.n233 B 0.037026f
C540 VTAIL.n234 B 0.037026f
C541 VTAIL.n235 B 0.016126f
C542 VTAIL.n236 B 0.015665f
C543 VTAIL.n237 B 0.029152f
C544 VTAIL.n238 B 0.029152f
C545 VTAIL.n239 B 0.015665f
C546 VTAIL.n240 B 0.016586f
C547 VTAIL.n241 B 0.037026f
C548 VTAIL.n242 B 0.037026f
C549 VTAIL.n243 B 0.016586f
C550 VTAIL.n244 B 0.015665f
C551 VTAIL.n245 B 0.029152f
C552 VTAIL.n246 B 0.029152f
C553 VTAIL.n247 B 0.015665f
C554 VTAIL.n248 B 0.016586f
C555 VTAIL.n249 B 0.037026f
C556 VTAIL.n250 B 0.074938f
C557 VTAIL.n251 B 0.016586f
C558 VTAIL.n252 B 0.015665f
C559 VTAIL.n253 B 0.063002f
C560 VTAIL.n254 B 0.041256f
C561 VTAIL.n255 B 1.41363f
C562 VN.t0 B 0.527636f
C563 VN.n0 B 0.22706f
C564 VN.t2 B 0.517753f
C565 VN.n1 B 0.208716f
C566 VN.t5 B 0.527636f
C567 VN.n2 B 0.226971f
C568 VN.n3 B 0.120557f
C569 VN.t3 B 0.527636f
C570 VN.n4 B 0.22706f
C571 VN.t4 B 0.527636f
C572 VN.t1 B 0.517753f
C573 VN.n5 B 0.208716f
C574 VN.n6 B 0.226971f
C575 VN.n7 B 2.23514f
.ends

