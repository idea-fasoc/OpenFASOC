* NGSPICE file created from diff_pair_sample_0288.ext - technology: sky130A

.subckt diff_pair_sample_0288 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t15 VN.t0 VDD2.t7 w_n3510_n1422# sky130_fd_pr__pfet_01v8 ad=0.8853 pd=5.32 as=0.37455 ps=2.6 w=2.27 l=2.21
X1 B.t11 B.t9 B.t10 w_n3510_n1422# sky130_fd_pr__pfet_01v8 ad=0.8853 pd=5.32 as=0 ps=0 w=2.27 l=2.21
X2 VDD1.t7 VP.t0 VTAIL.t6 w_n3510_n1422# sky130_fd_pr__pfet_01v8 ad=0.37455 pd=2.6 as=0.8853 ps=5.32 w=2.27 l=2.21
X3 VDD2.t6 VN.t1 VTAIL.t14 w_n3510_n1422# sky130_fd_pr__pfet_01v8 ad=0.37455 pd=2.6 as=0.37455 ps=2.6 w=2.27 l=2.21
X4 VTAIL.t7 VP.t1 VDD1.t6 w_n3510_n1422# sky130_fd_pr__pfet_01v8 ad=0.37455 pd=2.6 as=0.37455 ps=2.6 w=2.27 l=2.21
X5 VTAIL.t13 VN.t2 VDD2.t4 w_n3510_n1422# sky130_fd_pr__pfet_01v8 ad=0.8853 pd=5.32 as=0.37455 ps=2.6 w=2.27 l=2.21
X6 VDD1.t5 VP.t2 VTAIL.t5 w_n3510_n1422# sky130_fd_pr__pfet_01v8 ad=0.37455 pd=2.6 as=0.37455 ps=2.6 w=2.27 l=2.21
X7 VTAIL.t12 VN.t3 VDD2.t0 w_n3510_n1422# sky130_fd_pr__pfet_01v8 ad=0.37455 pd=2.6 as=0.37455 ps=2.6 w=2.27 l=2.21
X8 VDD1.t4 VP.t3 VTAIL.t0 w_n3510_n1422# sky130_fd_pr__pfet_01v8 ad=0.37455 pd=2.6 as=0.37455 ps=2.6 w=2.27 l=2.21
X9 VTAIL.t1 VP.t4 VDD1.t3 w_n3510_n1422# sky130_fd_pr__pfet_01v8 ad=0.8853 pd=5.32 as=0.37455 ps=2.6 w=2.27 l=2.21
X10 VDD2.t5 VN.t4 VTAIL.t11 w_n3510_n1422# sky130_fd_pr__pfet_01v8 ad=0.37455 pd=2.6 as=0.37455 ps=2.6 w=2.27 l=2.21
X11 B.t8 B.t6 B.t7 w_n3510_n1422# sky130_fd_pr__pfet_01v8 ad=0.8853 pd=5.32 as=0 ps=0 w=2.27 l=2.21
X12 VDD2.t3 VN.t5 VTAIL.t10 w_n3510_n1422# sky130_fd_pr__pfet_01v8 ad=0.37455 pd=2.6 as=0.8853 ps=5.32 w=2.27 l=2.21
X13 B.t5 B.t3 B.t4 w_n3510_n1422# sky130_fd_pr__pfet_01v8 ad=0.8853 pd=5.32 as=0 ps=0 w=2.27 l=2.21
X14 VTAIL.t2 VP.t5 VDD1.t2 w_n3510_n1422# sky130_fd_pr__pfet_01v8 ad=0.8853 pd=5.32 as=0.37455 ps=2.6 w=2.27 l=2.21
X15 B.t2 B.t0 B.t1 w_n3510_n1422# sky130_fd_pr__pfet_01v8 ad=0.8853 pd=5.32 as=0 ps=0 w=2.27 l=2.21
X16 VDD1.t1 VP.t6 VTAIL.t3 w_n3510_n1422# sky130_fd_pr__pfet_01v8 ad=0.37455 pd=2.6 as=0.8853 ps=5.32 w=2.27 l=2.21
X17 VTAIL.t4 VP.t7 VDD1.t0 w_n3510_n1422# sky130_fd_pr__pfet_01v8 ad=0.37455 pd=2.6 as=0.37455 ps=2.6 w=2.27 l=2.21
X18 VTAIL.t9 VN.t6 VDD2.t2 w_n3510_n1422# sky130_fd_pr__pfet_01v8 ad=0.37455 pd=2.6 as=0.37455 ps=2.6 w=2.27 l=2.21
X19 VDD2.t1 VN.t7 VTAIL.t8 w_n3510_n1422# sky130_fd_pr__pfet_01v8 ad=0.37455 pd=2.6 as=0.8853 ps=5.32 w=2.27 l=2.21
R0 VN.n47 VN.n25 161.3
R1 VN.n46 VN.n45 161.3
R2 VN.n44 VN.n26 161.3
R3 VN.n43 VN.n42 161.3
R4 VN.n41 VN.n27 161.3
R5 VN.n39 VN.n38 161.3
R6 VN.n37 VN.n28 161.3
R7 VN.n36 VN.n35 161.3
R8 VN.n34 VN.n29 161.3
R9 VN.n33 VN.n32 161.3
R10 VN.n22 VN.n0 161.3
R11 VN.n21 VN.n20 161.3
R12 VN.n19 VN.n1 161.3
R13 VN.n18 VN.n17 161.3
R14 VN.n16 VN.n2 161.3
R15 VN.n14 VN.n13 161.3
R16 VN.n12 VN.n3 161.3
R17 VN.n11 VN.n10 161.3
R18 VN.n9 VN.n4 161.3
R19 VN.n8 VN.n7 161.3
R20 VN.n24 VN.n23 95.5869
R21 VN.n49 VN.n48 95.5869
R22 VN.n6 VN.n5 58.1831
R23 VN.n31 VN.n30 58.1831
R24 VN.n6 VN.t0 57.6172
R25 VN.n31 VN.t5 57.6172
R26 VN.n21 VN.n1 44.3785
R27 VN.n46 VN.n26 44.3785
R28 VN VN.n49 41.983
R29 VN.n10 VN.n9 40.4934
R30 VN.n10 VN.n3 40.4934
R31 VN.n35 VN.n34 40.4934
R32 VN.n35 VN.n28 40.4934
R33 VN.n17 VN.n1 36.6083
R34 VN.n42 VN.n26 36.6083
R35 VN.n5 VN.t1 24.7548
R36 VN.n15 VN.t6 24.7548
R37 VN.n23 VN.t7 24.7548
R38 VN.n30 VN.t3 24.7548
R39 VN.n40 VN.t4 24.7548
R40 VN.n48 VN.t2 24.7548
R41 VN.n9 VN.n8 24.4675
R42 VN.n14 VN.n3 24.4675
R43 VN.n17 VN.n16 24.4675
R44 VN.n22 VN.n21 24.4675
R45 VN.n34 VN.n33 24.4675
R46 VN.n42 VN.n41 24.4675
R47 VN.n39 VN.n28 24.4675
R48 VN.n47 VN.n46 24.4675
R49 VN.n23 VN.n22 15.17
R50 VN.n48 VN.n47 15.17
R51 VN.n8 VN.n5 13.2127
R52 VN.n15 VN.n14 13.2127
R53 VN.n33 VN.n30 13.2127
R54 VN.n40 VN.n39 13.2127
R55 VN.n16 VN.n15 11.2553
R56 VN.n41 VN.n40 11.2553
R57 VN.n32 VN.n31 9.43557
R58 VN.n7 VN.n6 9.43557
R59 VN.n49 VN.n25 0.278367
R60 VN.n24 VN.n0 0.278367
R61 VN.n45 VN.n25 0.189894
R62 VN.n45 VN.n44 0.189894
R63 VN.n44 VN.n43 0.189894
R64 VN.n43 VN.n27 0.189894
R65 VN.n38 VN.n27 0.189894
R66 VN.n38 VN.n37 0.189894
R67 VN.n37 VN.n36 0.189894
R68 VN.n36 VN.n29 0.189894
R69 VN.n32 VN.n29 0.189894
R70 VN.n7 VN.n4 0.189894
R71 VN.n11 VN.n4 0.189894
R72 VN.n12 VN.n11 0.189894
R73 VN.n13 VN.n12 0.189894
R74 VN.n13 VN.n2 0.189894
R75 VN.n18 VN.n2 0.189894
R76 VN.n19 VN.n18 0.189894
R77 VN.n20 VN.n19 0.189894
R78 VN.n20 VN.n0 0.189894
R79 VN VN.n24 0.153454
R80 VDD2.n2 VDD2.n1 176.339
R81 VDD2.n2 VDD2.n0 176.339
R82 VDD2 VDD2.n5 176.337
R83 VDD2.n4 VDD2.n3 175.299
R84 VDD2.n4 VDD2.n2 35.5256
R85 VDD2.n5 VDD2.t0 14.3199
R86 VDD2.n5 VDD2.t3 14.3199
R87 VDD2.n3 VDD2.t4 14.3199
R88 VDD2.n3 VDD2.t5 14.3199
R89 VDD2.n1 VDD2.t2 14.3199
R90 VDD2.n1 VDD2.t1 14.3199
R91 VDD2.n0 VDD2.t7 14.3199
R92 VDD2.n0 VDD2.t6 14.3199
R93 VDD2 VDD2.n4 1.15352
R94 VTAIL.n15 VTAIL.t8 172.94
R95 VTAIL.n2 VTAIL.t15 172.94
R96 VTAIL.n3 VTAIL.t3 172.94
R97 VTAIL.n6 VTAIL.t1 172.94
R98 VTAIL.n14 VTAIL.t6 172.94
R99 VTAIL.n11 VTAIL.t2 172.94
R100 VTAIL.n10 VTAIL.t10 172.94
R101 VTAIL.n7 VTAIL.t13 172.94
R102 VTAIL.n13 VTAIL.n12 158.621
R103 VTAIL.n9 VTAIL.n8 158.621
R104 VTAIL.n1 VTAIL.n0 158.62
R105 VTAIL.n5 VTAIL.n4 158.62
R106 VTAIL.n15 VTAIL.n14 16.5134
R107 VTAIL.n7 VTAIL.n6 16.5134
R108 VTAIL.n0 VTAIL.t14 14.3199
R109 VTAIL.n0 VTAIL.t9 14.3199
R110 VTAIL.n4 VTAIL.t0 14.3199
R111 VTAIL.n4 VTAIL.t4 14.3199
R112 VTAIL.n12 VTAIL.t5 14.3199
R113 VTAIL.n12 VTAIL.t7 14.3199
R114 VTAIL.n8 VTAIL.t11 14.3199
R115 VTAIL.n8 VTAIL.t12 14.3199
R116 VTAIL.n9 VTAIL.n7 2.19016
R117 VTAIL.n10 VTAIL.n9 2.19016
R118 VTAIL.n13 VTAIL.n11 2.19016
R119 VTAIL.n14 VTAIL.n13 2.19016
R120 VTAIL.n6 VTAIL.n5 2.19016
R121 VTAIL.n5 VTAIL.n3 2.19016
R122 VTAIL.n2 VTAIL.n1 2.19016
R123 VTAIL VTAIL.n15 2.13197
R124 VTAIL.n11 VTAIL.n10 0.470328
R125 VTAIL.n3 VTAIL.n2 0.470328
R126 VTAIL VTAIL.n1 0.0586897
R127 B.n258 B.n93 585
R128 B.n257 B.n256 585
R129 B.n255 B.n94 585
R130 B.n254 B.n253 585
R131 B.n252 B.n95 585
R132 B.n251 B.n250 585
R133 B.n249 B.n96 585
R134 B.n248 B.n247 585
R135 B.n246 B.n97 585
R136 B.n245 B.n244 585
R137 B.n243 B.n98 585
R138 B.n242 B.n241 585
R139 B.n240 B.n99 585
R140 B.n238 B.n237 585
R141 B.n236 B.n102 585
R142 B.n235 B.n234 585
R143 B.n233 B.n103 585
R144 B.n232 B.n231 585
R145 B.n230 B.n104 585
R146 B.n229 B.n228 585
R147 B.n227 B.n105 585
R148 B.n226 B.n225 585
R149 B.n224 B.n106 585
R150 B.n223 B.n222 585
R151 B.n218 B.n107 585
R152 B.n217 B.n216 585
R153 B.n215 B.n108 585
R154 B.n214 B.n213 585
R155 B.n212 B.n109 585
R156 B.n211 B.n210 585
R157 B.n209 B.n110 585
R158 B.n208 B.n207 585
R159 B.n206 B.n111 585
R160 B.n205 B.n204 585
R161 B.n203 B.n112 585
R162 B.n202 B.n201 585
R163 B.n260 B.n259 585
R164 B.n261 B.n92 585
R165 B.n263 B.n262 585
R166 B.n264 B.n91 585
R167 B.n266 B.n265 585
R168 B.n267 B.n90 585
R169 B.n269 B.n268 585
R170 B.n270 B.n89 585
R171 B.n272 B.n271 585
R172 B.n273 B.n88 585
R173 B.n275 B.n274 585
R174 B.n276 B.n87 585
R175 B.n278 B.n277 585
R176 B.n279 B.n86 585
R177 B.n281 B.n280 585
R178 B.n282 B.n85 585
R179 B.n284 B.n283 585
R180 B.n285 B.n84 585
R181 B.n287 B.n286 585
R182 B.n288 B.n83 585
R183 B.n290 B.n289 585
R184 B.n291 B.n82 585
R185 B.n293 B.n292 585
R186 B.n294 B.n81 585
R187 B.n296 B.n295 585
R188 B.n297 B.n80 585
R189 B.n299 B.n298 585
R190 B.n300 B.n79 585
R191 B.n302 B.n301 585
R192 B.n303 B.n78 585
R193 B.n305 B.n304 585
R194 B.n306 B.n77 585
R195 B.n308 B.n307 585
R196 B.n309 B.n76 585
R197 B.n311 B.n310 585
R198 B.n312 B.n75 585
R199 B.n314 B.n313 585
R200 B.n315 B.n74 585
R201 B.n317 B.n316 585
R202 B.n318 B.n73 585
R203 B.n320 B.n319 585
R204 B.n321 B.n72 585
R205 B.n323 B.n322 585
R206 B.n324 B.n71 585
R207 B.n326 B.n325 585
R208 B.n327 B.n70 585
R209 B.n329 B.n328 585
R210 B.n330 B.n69 585
R211 B.n332 B.n331 585
R212 B.n333 B.n68 585
R213 B.n335 B.n334 585
R214 B.n336 B.n67 585
R215 B.n338 B.n337 585
R216 B.n339 B.n66 585
R217 B.n341 B.n340 585
R218 B.n342 B.n65 585
R219 B.n344 B.n343 585
R220 B.n345 B.n64 585
R221 B.n347 B.n346 585
R222 B.n348 B.n63 585
R223 B.n350 B.n349 585
R224 B.n351 B.n62 585
R225 B.n353 B.n352 585
R226 B.n354 B.n61 585
R227 B.n356 B.n355 585
R228 B.n357 B.n60 585
R229 B.n359 B.n358 585
R230 B.n360 B.n59 585
R231 B.n362 B.n361 585
R232 B.n363 B.n58 585
R233 B.n365 B.n364 585
R234 B.n366 B.n57 585
R235 B.n368 B.n367 585
R236 B.n369 B.n56 585
R237 B.n371 B.n370 585
R238 B.n372 B.n55 585
R239 B.n374 B.n373 585
R240 B.n375 B.n54 585
R241 B.n377 B.n376 585
R242 B.n378 B.n53 585
R243 B.n380 B.n379 585
R244 B.n381 B.n52 585
R245 B.n383 B.n382 585
R246 B.n384 B.n51 585
R247 B.n386 B.n385 585
R248 B.n387 B.n50 585
R249 B.n389 B.n388 585
R250 B.n390 B.n49 585
R251 B.n392 B.n391 585
R252 B.n393 B.n48 585
R253 B.n395 B.n394 585
R254 B.n396 B.n47 585
R255 B.n452 B.n451 585
R256 B.n450 B.n25 585
R257 B.n449 B.n448 585
R258 B.n447 B.n26 585
R259 B.n446 B.n445 585
R260 B.n444 B.n27 585
R261 B.n443 B.n442 585
R262 B.n441 B.n28 585
R263 B.n440 B.n439 585
R264 B.n438 B.n29 585
R265 B.n437 B.n436 585
R266 B.n435 B.n30 585
R267 B.n434 B.n433 585
R268 B.n431 B.n31 585
R269 B.n430 B.n429 585
R270 B.n428 B.n34 585
R271 B.n427 B.n426 585
R272 B.n425 B.n35 585
R273 B.n424 B.n423 585
R274 B.n422 B.n36 585
R275 B.n421 B.n420 585
R276 B.n419 B.n37 585
R277 B.n418 B.n417 585
R278 B.n416 B.n415 585
R279 B.n414 B.n41 585
R280 B.n413 B.n412 585
R281 B.n411 B.n42 585
R282 B.n410 B.n409 585
R283 B.n408 B.n43 585
R284 B.n407 B.n406 585
R285 B.n405 B.n44 585
R286 B.n404 B.n403 585
R287 B.n402 B.n45 585
R288 B.n401 B.n400 585
R289 B.n399 B.n46 585
R290 B.n398 B.n397 585
R291 B.n453 B.n24 585
R292 B.n455 B.n454 585
R293 B.n456 B.n23 585
R294 B.n458 B.n457 585
R295 B.n459 B.n22 585
R296 B.n461 B.n460 585
R297 B.n462 B.n21 585
R298 B.n464 B.n463 585
R299 B.n465 B.n20 585
R300 B.n467 B.n466 585
R301 B.n468 B.n19 585
R302 B.n470 B.n469 585
R303 B.n471 B.n18 585
R304 B.n473 B.n472 585
R305 B.n474 B.n17 585
R306 B.n476 B.n475 585
R307 B.n477 B.n16 585
R308 B.n479 B.n478 585
R309 B.n480 B.n15 585
R310 B.n482 B.n481 585
R311 B.n483 B.n14 585
R312 B.n485 B.n484 585
R313 B.n486 B.n13 585
R314 B.n488 B.n487 585
R315 B.n489 B.n12 585
R316 B.n491 B.n490 585
R317 B.n492 B.n11 585
R318 B.n494 B.n493 585
R319 B.n495 B.n10 585
R320 B.n497 B.n496 585
R321 B.n498 B.n9 585
R322 B.n500 B.n499 585
R323 B.n501 B.n8 585
R324 B.n503 B.n502 585
R325 B.n504 B.n7 585
R326 B.n506 B.n505 585
R327 B.n507 B.n6 585
R328 B.n509 B.n508 585
R329 B.n510 B.n5 585
R330 B.n512 B.n511 585
R331 B.n513 B.n4 585
R332 B.n515 B.n514 585
R333 B.n516 B.n3 585
R334 B.n518 B.n517 585
R335 B.n519 B.n0 585
R336 B.n2 B.n1 585
R337 B.n136 B.n135 585
R338 B.n137 B.n134 585
R339 B.n139 B.n138 585
R340 B.n140 B.n133 585
R341 B.n142 B.n141 585
R342 B.n143 B.n132 585
R343 B.n145 B.n144 585
R344 B.n146 B.n131 585
R345 B.n148 B.n147 585
R346 B.n149 B.n130 585
R347 B.n151 B.n150 585
R348 B.n152 B.n129 585
R349 B.n154 B.n153 585
R350 B.n155 B.n128 585
R351 B.n157 B.n156 585
R352 B.n158 B.n127 585
R353 B.n160 B.n159 585
R354 B.n161 B.n126 585
R355 B.n163 B.n162 585
R356 B.n164 B.n125 585
R357 B.n166 B.n165 585
R358 B.n167 B.n124 585
R359 B.n169 B.n168 585
R360 B.n170 B.n123 585
R361 B.n172 B.n171 585
R362 B.n173 B.n122 585
R363 B.n175 B.n174 585
R364 B.n176 B.n121 585
R365 B.n178 B.n177 585
R366 B.n179 B.n120 585
R367 B.n181 B.n180 585
R368 B.n182 B.n119 585
R369 B.n184 B.n183 585
R370 B.n185 B.n118 585
R371 B.n187 B.n186 585
R372 B.n188 B.n117 585
R373 B.n190 B.n189 585
R374 B.n191 B.n116 585
R375 B.n193 B.n192 585
R376 B.n194 B.n115 585
R377 B.n196 B.n195 585
R378 B.n197 B.n114 585
R379 B.n199 B.n198 585
R380 B.n200 B.n113 585
R381 B.n202 B.n113 458.866
R382 B.n260 B.n93 458.866
R383 B.n398 B.n47 458.866
R384 B.n453 B.n452 458.866
R385 B.n521 B.n520 256.663
R386 B.n520 B.n519 235.042
R387 B.n520 B.n2 235.042
R388 B.n219 B.t0 232.125
R389 B.n100 B.t6 232.125
R390 B.n38 B.t9 232.125
R391 B.n32 B.t3 232.125
R392 B.n100 B.t7 223.011
R393 B.n38 B.t11 223.011
R394 B.n219 B.t1 223.011
R395 B.n32 B.t5 223.011
R396 B.n101 B.t8 173.75
R397 B.n39 B.t10 173.75
R398 B.n220 B.t2 173.75
R399 B.n33 B.t4 173.75
R400 B.n203 B.n202 163.367
R401 B.n204 B.n203 163.367
R402 B.n204 B.n111 163.367
R403 B.n208 B.n111 163.367
R404 B.n209 B.n208 163.367
R405 B.n210 B.n209 163.367
R406 B.n210 B.n109 163.367
R407 B.n214 B.n109 163.367
R408 B.n215 B.n214 163.367
R409 B.n216 B.n215 163.367
R410 B.n216 B.n107 163.367
R411 B.n223 B.n107 163.367
R412 B.n224 B.n223 163.367
R413 B.n225 B.n224 163.367
R414 B.n225 B.n105 163.367
R415 B.n229 B.n105 163.367
R416 B.n230 B.n229 163.367
R417 B.n231 B.n230 163.367
R418 B.n231 B.n103 163.367
R419 B.n235 B.n103 163.367
R420 B.n236 B.n235 163.367
R421 B.n237 B.n236 163.367
R422 B.n237 B.n99 163.367
R423 B.n242 B.n99 163.367
R424 B.n243 B.n242 163.367
R425 B.n244 B.n243 163.367
R426 B.n244 B.n97 163.367
R427 B.n248 B.n97 163.367
R428 B.n249 B.n248 163.367
R429 B.n250 B.n249 163.367
R430 B.n250 B.n95 163.367
R431 B.n254 B.n95 163.367
R432 B.n255 B.n254 163.367
R433 B.n256 B.n255 163.367
R434 B.n256 B.n93 163.367
R435 B.n394 B.n47 163.367
R436 B.n394 B.n393 163.367
R437 B.n393 B.n392 163.367
R438 B.n392 B.n49 163.367
R439 B.n388 B.n49 163.367
R440 B.n388 B.n387 163.367
R441 B.n387 B.n386 163.367
R442 B.n386 B.n51 163.367
R443 B.n382 B.n51 163.367
R444 B.n382 B.n381 163.367
R445 B.n381 B.n380 163.367
R446 B.n380 B.n53 163.367
R447 B.n376 B.n53 163.367
R448 B.n376 B.n375 163.367
R449 B.n375 B.n374 163.367
R450 B.n374 B.n55 163.367
R451 B.n370 B.n55 163.367
R452 B.n370 B.n369 163.367
R453 B.n369 B.n368 163.367
R454 B.n368 B.n57 163.367
R455 B.n364 B.n57 163.367
R456 B.n364 B.n363 163.367
R457 B.n363 B.n362 163.367
R458 B.n362 B.n59 163.367
R459 B.n358 B.n59 163.367
R460 B.n358 B.n357 163.367
R461 B.n357 B.n356 163.367
R462 B.n356 B.n61 163.367
R463 B.n352 B.n61 163.367
R464 B.n352 B.n351 163.367
R465 B.n351 B.n350 163.367
R466 B.n350 B.n63 163.367
R467 B.n346 B.n63 163.367
R468 B.n346 B.n345 163.367
R469 B.n345 B.n344 163.367
R470 B.n344 B.n65 163.367
R471 B.n340 B.n65 163.367
R472 B.n340 B.n339 163.367
R473 B.n339 B.n338 163.367
R474 B.n338 B.n67 163.367
R475 B.n334 B.n67 163.367
R476 B.n334 B.n333 163.367
R477 B.n333 B.n332 163.367
R478 B.n332 B.n69 163.367
R479 B.n328 B.n69 163.367
R480 B.n328 B.n327 163.367
R481 B.n327 B.n326 163.367
R482 B.n326 B.n71 163.367
R483 B.n322 B.n71 163.367
R484 B.n322 B.n321 163.367
R485 B.n321 B.n320 163.367
R486 B.n320 B.n73 163.367
R487 B.n316 B.n73 163.367
R488 B.n316 B.n315 163.367
R489 B.n315 B.n314 163.367
R490 B.n314 B.n75 163.367
R491 B.n310 B.n75 163.367
R492 B.n310 B.n309 163.367
R493 B.n309 B.n308 163.367
R494 B.n308 B.n77 163.367
R495 B.n304 B.n77 163.367
R496 B.n304 B.n303 163.367
R497 B.n303 B.n302 163.367
R498 B.n302 B.n79 163.367
R499 B.n298 B.n79 163.367
R500 B.n298 B.n297 163.367
R501 B.n297 B.n296 163.367
R502 B.n296 B.n81 163.367
R503 B.n292 B.n81 163.367
R504 B.n292 B.n291 163.367
R505 B.n291 B.n290 163.367
R506 B.n290 B.n83 163.367
R507 B.n286 B.n83 163.367
R508 B.n286 B.n285 163.367
R509 B.n285 B.n284 163.367
R510 B.n284 B.n85 163.367
R511 B.n280 B.n85 163.367
R512 B.n280 B.n279 163.367
R513 B.n279 B.n278 163.367
R514 B.n278 B.n87 163.367
R515 B.n274 B.n87 163.367
R516 B.n274 B.n273 163.367
R517 B.n273 B.n272 163.367
R518 B.n272 B.n89 163.367
R519 B.n268 B.n89 163.367
R520 B.n268 B.n267 163.367
R521 B.n267 B.n266 163.367
R522 B.n266 B.n91 163.367
R523 B.n262 B.n91 163.367
R524 B.n262 B.n261 163.367
R525 B.n261 B.n260 163.367
R526 B.n452 B.n25 163.367
R527 B.n448 B.n25 163.367
R528 B.n448 B.n447 163.367
R529 B.n447 B.n446 163.367
R530 B.n446 B.n27 163.367
R531 B.n442 B.n27 163.367
R532 B.n442 B.n441 163.367
R533 B.n441 B.n440 163.367
R534 B.n440 B.n29 163.367
R535 B.n436 B.n29 163.367
R536 B.n436 B.n435 163.367
R537 B.n435 B.n434 163.367
R538 B.n434 B.n31 163.367
R539 B.n429 B.n31 163.367
R540 B.n429 B.n428 163.367
R541 B.n428 B.n427 163.367
R542 B.n427 B.n35 163.367
R543 B.n423 B.n35 163.367
R544 B.n423 B.n422 163.367
R545 B.n422 B.n421 163.367
R546 B.n421 B.n37 163.367
R547 B.n417 B.n37 163.367
R548 B.n417 B.n416 163.367
R549 B.n416 B.n41 163.367
R550 B.n412 B.n41 163.367
R551 B.n412 B.n411 163.367
R552 B.n411 B.n410 163.367
R553 B.n410 B.n43 163.367
R554 B.n406 B.n43 163.367
R555 B.n406 B.n405 163.367
R556 B.n405 B.n404 163.367
R557 B.n404 B.n45 163.367
R558 B.n400 B.n45 163.367
R559 B.n400 B.n399 163.367
R560 B.n399 B.n398 163.367
R561 B.n454 B.n453 163.367
R562 B.n454 B.n23 163.367
R563 B.n458 B.n23 163.367
R564 B.n459 B.n458 163.367
R565 B.n460 B.n459 163.367
R566 B.n460 B.n21 163.367
R567 B.n464 B.n21 163.367
R568 B.n465 B.n464 163.367
R569 B.n466 B.n465 163.367
R570 B.n466 B.n19 163.367
R571 B.n470 B.n19 163.367
R572 B.n471 B.n470 163.367
R573 B.n472 B.n471 163.367
R574 B.n472 B.n17 163.367
R575 B.n476 B.n17 163.367
R576 B.n477 B.n476 163.367
R577 B.n478 B.n477 163.367
R578 B.n478 B.n15 163.367
R579 B.n482 B.n15 163.367
R580 B.n483 B.n482 163.367
R581 B.n484 B.n483 163.367
R582 B.n484 B.n13 163.367
R583 B.n488 B.n13 163.367
R584 B.n489 B.n488 163.367
R585 B.n490 B.n489 163.367
R586 B.n490 B.n11 163.367
R587 B.n494 B.n11 163.367
R588 B.n495 B.n494 163.367
R589 B.n496 B.n495 163.367
R590 B.n496 B.n9 163.367
R591 B.n500 B.n9 163.367
R592 B.n501 B.n500 163.367
R593 B.n502 B.n501 163.367
R594 B.n502 B.n7 163.367
R595 B.n506 B.n7 163.367
R596 B.n507 B.n506 163.367
R597 B.n508 B.n507 163.367
R598 B.n508 B.n5 163.367
R599 B.n512 B.n5 163.367
R600 B.n513 B.n512 163.367
R601 B.n514 B.n513 163.367
R602 B.n514 B.n3 163.367
R603 B.n518 B.n3 163.367
R604 B.n519 B.n518 163.367
R605 B.n136 B.n2 163.367
R606 B.n137 B.n136 163.367
R607 B.n138 B.n137 163.367
R608 B.n138 B.n133 163.367
R609 B.n142 B.n133 163.367
R610 B.n143 B.n142 163.367
R611 B.n144 B.n143 163.367
R612 B.n144 B.n131 163.367
R613 B.n148 B.n131 163.367
R614 B.n149 B.n148 163.367
R615 B.n150 B.n149 163.367
R616 B.n150 B.n129 163.367
R617 B.n154 B.n129 163.367
R618 B.n155 B.n154 163.367
R619 B.n156 B.n155 163.367
R620 B.n156 B.n127 163.367
R621 B.n160 B.n127 163.367
R622 B.n161 B.n160 163.367
R623 B.n162 B.n161 163.367
R624 B.n162 B.n125 163.367
R625 B.n166 B.n125 163.367
R626 B.n167 B.n166 163.367
R627 B.n168 B.n167 163.367
R628 B.n168 B.n123 163.367
R629 B.n172 B.n123 163.367
R630 B.n173 B.n172 163.367
R631 B.n174 B.n173 163.367
R632 B.n174 B.n121 163.367
R633 B.n178 B.n121 163.367
R634 B.n179 B.n178 163.367
R635 B.n180 B.n179 163.367
R636 B.n180 B.n119 163.367
R637 B.n184 B.n119 163.367
R638 B.n185 B.n184 163.367
R639 B.n186 B.n185 163.367
R640 B.n186 B.n117 163.367
R641 B.n190 B.n117 163.367
R642 B.n191 B.n190 163.367
R643 B.n192 B.n191 163.367
R644 B.n192 B.n115 163.367
R645 B.n196 B.n115 163.367
R646 B.n197 B.n196 163.367
R647 B.n198 B.n197 163.367
R648 B.n198 B.n113 163.367
R649 B.n221 B.n220 59.5399
R650 B.n239 B.n101 59.5399
R651 B.n40 B.n39 59.5399
R652 B.n432 B.n33 59.5399
R653 B.n220 B.n219 49.2611
R654 B.n101 B.n100 49.2611
R655 B.n39 B.n38 49.2611
R656 B.n33 B.n32 49.2611
R657 B.n259 B.n258 29.8151
R658 B.n451 B.n24 29.8151
R659 B.n397 B.n396 29.8151
R660 B.n201 B.n200 29.8151
R661 B B.n521 18.0485
R662 B.n455 B.n24 10.6151
R663 B.n456 B.n455 10.6151
R664 B.n457 B.n456 10.6151
R665 B.n457 B.n22 10.6151
R666 B.n461 B.n22 10.6151
R667 B.n462 B.n461 10.6151
R668 B.n463 B.n462 10.6151
R669 B.n463 B.n20 10.6151
R670 B.n467 B.n20 10.6151
R671 B.n468 B.n467 10.6151
R672 B.n469 B.n468 10.6151
R673 B.n469 B.n18 10.6151
R674 B.n473 B.n18 10.6151
R675 B.n474 B.n473 10.6151
R676 B.n475 B.n474 10.6151
R677 B.n475 B.n16 10.6151
R678 B.n479 B.n16 10.6151
R679 B.n480 B.n479 10.6151
R680 B.n481 B.n480 10.6151
R681 B.n481 B.n14 10.6151
R682 B.n485 B.n14 10.6151
R683 B.n486 B.n485 10.6151
R684 B.n487 B.n486 10.6151
R685 B.n487 B.n12 10.6151
R686 B.n491 B.n12 10.6151
R687 B.n492 B.n491 10.6151
R688 B.n493 B.n492 10.6151
R689 B.n493 B.n10 10.6151
R690 B.n497 B.n10 10.6151
R691 B.n498 B.n497 10.6151
R692 B.n499 B.n498 10.6151
R693 B.n499 B.n8 10.6151
R694 B.n503 B.n8 10.6151
R695 B.n504 B.n503 10.6151
R696 B.n505 B.n504 10.6151
R697 B.n505 B.n6 10.6151
R698 B.n509 B.n6 10.6151
R699 B.n510 B.n509 10.6151
R700 B.n511 B.n510 10.6151
R701 B.n511 B.n4 10.6151
R702 B.n515 B.n4 10.6151
R703 B.n516 B.n515 10.6151
R704 B.n517 B.n516 10.6151
R705 B.n517 B.n0 10.6151
R706 B.n451 B.n450 10.6151
R707 B.n450 B.n449 10.6151
R708 B.n449 B.n26 10.6151
R709 B.n445 B.n26 10.6151
R710 B.n445 B.n444 10.6151
R711 B.n444 B.n443 10.6151
R712 B.n443 B.n28 10.6151
R713 B.n439 B.n28 10.6151
R714 B.n439 B.n438 10.6151
R715 B.n438 B.n437 10.6151
R716 B.n437 B.n30 10.6151
R717 B.n433 B.n30 10.6151
R718 B.n431 B.n430 10.6151
R719 B.n430 B.n34 10.6151
R720 B.n426 B.n34 10.6151
R721 B.n426 B.n425 10.6151
R722 B.n425 B.n424 10.6151
R723 B.n424 B.n36 10.6151
R724 B.n420 B.n36 10.6151
R725 B.n420 B.n419 10.6151
R726 B.n419 B.n418 10.6151
R727 B.n415 B.n414 10.6151
R728 B.n414 B.n413 10.6151
R729 B.n413 B.n42 10.6151
R730 B.n409 B.n42 10.6151
R731 B.n409 B.n408 10.6151
R732 B.n408 B.n407 10.6151
R733 B.n407 B.n44 10.6151
R734 B.n403 B.n44 10.6151
R735 B.n403 B.n402 10.6151
R736 B.n402 B.n401 10.6151
R737 B.n401 B.n46 10.6151
R738 B.n397 B.n46 10.6151
R739 B.n396 B.n395 10.6151
R740 B.n395 B.n48 10.6151
R741 B.n391 B.n48 10.6151
R742 B.n391 B.n390 10.6151
R743 B.n390 B.n389 10.6151
R744 B.n389 B.n50 10.6151
R745 B.n385 B.n50 10.6151
R746 B.n385 B.n384 10.6151
R747 B.n384 B.n383 10.6151
R748 B.n383 B.n52 10.6151
R749 B.n379 B.n52 10.6151
R750 B.n379 B.n378 10.6151
R751 B.n378 B.n377 10.6151
R752 B.n377 B.n54 10.6151
R753 B.n373 B.n54 10.6151
R754 B.n373 B.n372 10.6151
R755 B.n372 B.n371 10.6151
R756 B.n371 B.n56 10.6151
R757 B.n367 B.n56 10.6151
R758 B.n367 B.n366 10.6151
R759 B.n366 B.n365 10.6151
R760 B.n365 B.n58 10.6151
R761 B.n361 B.n58 10.6151
R762 B.n361 B.n360 10.6151
R763 B.n360 B.n359 10.6151
R764 B.n359 B.n60 10.6151
R765 B.n355 B.n60 10.6151
R766 B.n355 B.n354 10.6151
R767 B.n354 B.n353 10.6151
R768 B.n353 B.n62 10.6151
R769 B.n349 B.n62 10.6151
R770 B.n349 B.n348 10.6151
R771 B.n348 B.n347 10.6151
R772 B.n347 B.n64 10.6151
R773 B.n343 B.n64 10.6151
R774 B.n343 B.n342 10.6151
R775 B.n342 B.n341 10.6151
R776 B.n341 B.n66 10.6151
R777 B.n337 B.n66 10.6151
R778 B.n337 B.n336 10.6151
R779 B.n336 B.n335 10.6151
R780 B.n335 B.n68 10.6151
R781 B.n331 B.n68 10.6151
R782 B.n331 B.n330 10.6151
R783 B.n330 B.n329 10.6151
R784 B.n329 B.n70 10.6151
R785 B.n325 B.n70 10.6151
R786 B.n325 B.n324 10.6151
R787 B.n324 B.n323 10.6151
R788 B.n323 B.n72 10.6151
R789 B.n319 B.n72 10.6151
R790 B.n319 B.n318 10.6151
R791 B.n318 B.n317 10.6151
R792 B.n317 B.n74 10.6151
R793 B.n313 B.n74 10.6151
R794 B.n313 B.n312 10.6151
R795 B.n312 B.n311 10.6151
R796 B.n311 B.n76 10.6151
R797 B.n307 B.n76 10.6151
R798 B.n307 B.n306 10.6151
R799 B.n306 B.n305 10.6151
R800 B.n305 B.n78 10.6151
R801 B.n301 B.n78 10.6151
R802 B.n301 B.n300 10.6151
R803 B.n300 B.n299 10.6151
R804 B.n299 B.n80 10.6151
R805 B.n295 B.n80 10.6151
R806 B.n295 B.n294 10.6151
R807 B.n294 B.n293 10.6151
R808 B.n293 B.n82 10.6151
R809 B.n289 B.n82 10.6151
R810 B.n289 B.n288 10.6151
R811 B.n288 B.n287 10.6151
R812 B.n287 B.n84 10.6151
R813 B.n283 B.n84 10.6151
R814 B.n283 B.n282 10.6151
R815 B.n282 B.n281 10.6151
R816 B.n281 B.n86 10.6151
R817 B.n277 B.n86 10.6151
R818 B.n277 B.n276 10.6151
R819 B.n276 B.n275 10.6151
R820 B.n275 B.n88 10.6151
R821 B.n271 B.n88 10.6151
R822 B.n271 B.n270 10.6151
R823 B.n270 B.n269 10.6151
R824 B.n269 B.n90 10.6151
R825 B.n265 B.n90 10.6151
R826 B.n265 B.n264 10.6151
R827 B.n264 B.n263 10.6151
R828 B.n263 B.n92 10.6151
R829 B.n259 B.n92 10.6151
R830 B.n135 B.n1 10.6151
R831 B.n135 B.n134 10.6151
R832 B.n139 B.n134 10.6151
R833 B.n140 B.n139 10.6151
R834 B.n141 B.n140 10.6151
R835 B.n141 B.n132 10.6151
R836 B.n145 B.n132 10.6151
R837 B.n146 B.n145 10.6151
R838 B.n147 B.n146 10.6151
R839 B.n147 B.n130 10.6151
R840 B.n151 B.n130 10.6151
R841 B.n152 B.n151 10.6151
R842 B.n153 B.n152 10.6151
R843 B.n153 B.n128 10.6151
R844 B.n157 B.n128 10.6151
R845 B.n158 B.n157 10.6151
R846 B.n159 B.n158 10.6151
R847 B.n159 B.n126 10.6151
R848 B.n163 B.n126 10.6151
R849 B.n164 B.n163 10.6151
R850 B.n165 B.n164 10.6151
R851 B.n165 B.n124 10.6151
R852 B.n169 B.n124 10.6151
R853 B.n170 B.n169 10.6151
R854 B.n171 B.n170 10.6151
R855 B.n171 B.n122 10.6151
R856 B.n175 B.n122 10.6151
R857 B.n176 B.n175 10.6151
R858 B.n177 B.n176 10.6151
R859 B.n177 B.n120 10.6151
R860 B.n181 B.n120 10.6151
R861 B.n182 B.n181 10.6151
R862 B.n183 B.n182 10.6151
R863 B.n183 B.n118 10.6151
R864 B.n187 B.n118 10.6151
R865 B.n188 B.n187 10.6151
R866 B.n189 B.n188 10.6151
R867 B.n189 B.n116 10.6151
R868 B.n193 B.n116 10.6151
R869 B.n194 B.n193 10.6151
R870 B.n195 B.n194 10.6151
R871 B.n195 B.n114 10.6151
R872 B.n199 B.n114 10.6151
R873 B.n200 B.n199 10.6151
R874 B.n201 B.n112 10.6151
R875 B.n205 B.n112 10.6151
R876 B.n206 B.n205 10.6151
R877 B.n207 B.n206 10.6151
R878 B.n207 B.n110 10.6151
R879 B.n211 B.n110 10.6151
R880 B.n212 B.n211 10.6151
R881 B.n213 B.n212 10.6151
R882 B.n213 B.n108 10.6151
R883 B.n217 B.n108 10.6151
R884 B.n218 B.n217 10.6151
R885 B.n222 B.n218 10.6151
R886 B.n226 B.n106 10.6151
R887 B.n227 B.n226 10.6151
R888 B.n228 B.n227 10.6151
R889 B.n228 B.n104 10.6151
R890 B.n232 B.n104 10.6151
R891 B.n233 B.n232 10.6151
R892 B.n234 B.n233 10.6151
R893 B.n234 B.n102 10.6151
R894 B.n238 B.n102 10.6151
R895 B.n241 B.n240 10.6151
R896 B.n241 B.n98 10.6151
R897 B.n245 B.n98 10.6151
R898 B.n246 B.n245 10.6151
R899 B.n247 B.n246 10.6151
R900 B.n247 B.n96 10.6151
R901 B.n251 B.n96 10.6151
R902 B.n252 B.n251 10.6151
R903 B.n253 B.n252 10.6151
R904 B.n253 B.n94 10.6151
R905 B.n257 B.n94 10.6151
R906 B.n258 B.n257 10.6151
R907 B.n433 B.n432 9.36635
R908 B.n415 B.n40 9.36635
R909 B.n222 B.n221 9.36635
R910 B.n240 B.n239 9.36635
R911 B.n521 B.n0 8.11757
R912 B.n521 B.n1 8.11757
R913 B.n432 B.n431 1.24928
R914 B.n418 B.n40 1.24928
R915 B.n221 B.n106 1.24928
R916 B.n239 B.n238 1.24928
R917 VP.n16 VP.n15 161.3
R918 VP.n17 VP.n12 161.3
R919 VP.n19 VP.n18 161.3
R920 VP.n20 VP.n11 161.3
R921 VP.n22 VP.n21 161.3
R922 VP.n24 VP.n10 161.3
R923 VP.n26 VP.n25 161.3
R924 VP.n27 VP.n9 161.3
R925 VP.n29 VP.n28 161.3
R926 VP.n30 VP.n8 161.3
R927 VP.n58 VP.n0 161.3
R928 VP.n57 VP.n56 161.3
R929 VP.n55 VP.n1 161.3
R930 VP.n54 VP.n53 161.3
R931 VP.n52 VP.n2 161.3
R932 VP.n50 VP.n49 161.3
R933 VP.n48 VP.n3 161.3
R934 VP.n47 VP.n46 161.3
R935 VP.n45 VP.n4 161.3
R936 VP.n44 VP.n43 161.3
R937 VP.n42 VP.n41 161.3
R938 VP.n40 VP.n6 161.3
R939 VP.n39 VP.n38 161.3
R940 VP.n37 VP.n7 161.3
R941 VP.n36 VP.n35 161.3
R942 VP.n34 VP.n33 95.5869
R943 VP.n60 VP.n59 95.5869
R944 VP.n32 VP.n31 95.5869
R945 VP.n14 VP.n13 58.1831
R946 VP.n14 VP.t5 57.6172
R947 VP.n39 VP.n7 44.3785
R948 VP.n57 VP.n1 44.3785
R949 VP.n29 VP.n9 44.3785
R950 VP.n33 VP.n32 41.7041
R951 VP.n46 VP.n45 40.4934
R952 VP.n46 VP.n3 40.4934
R953 VP.n18 VP.n11 40.4934
R954 VP.n18 VP.n17 40.4934
R955 VP.n40 VP.n39 36.6083
R956 VP.n53 VP.n1 36.6083
R957 VP.n25 VP.n9 36.6083
R958 VP.n34 VP.t4 24.7548
R959 VP.n5 VP.t3 24.7548
R960 VP.n51 VP.t7 24.7548
R961 VP.n59 VP.t6 24.7548
R962 VP.n31 VP.t0 24.7548
R963 VP.n23 VP.t1 24.7548
R964 VP.n13 VP.t2 24.7548
R965 VP.n35 VP.n7 24.4675
R966 VP.n41 VP.n40 24.4675
R967 VP.n45 VP.n44 24.4675
R968 VP.n50 VP.n3 24.4675
R969 VP.n53 VP.n52 24.4675
R970 VP.n58 VP.n57 24.4675
R971 VP.n30 VP.n29 24.4675
R972 VP.n22 VP.n11 24.4675
R973 VP.n25 VP.n24 24.4675
R974 VP.n17 VP.n16 24.4675
R975 VP.n35 VP.n34 15.17
R976 VP.n59 VP.n58 15.17
R977 VP.n31 VP.n30 15.17
R978 VP.n44 VP.n5 13.2127
R979 VP.n51 VP.n50 13.2127
R980 VP.n23 VP.n22 13.2127
R981 VP.n16 VP.n13 13.2127
R982 VP.n41 VP.n5 11.2553
R983 VP.n52 VP.n51 11.2553
R984 VP.n24 VP.n23 11.2553
R985 VP.n15 VP.n14 9.43557
R986 VP.n32 VP.n8 0.278367
R987 VP.n36 VP.n33 0.278367
R988 VP.n60 VP.n0 0.278367
R989 VP.n15 VP.n12 0.189894
R990 VP.n19 VP.n12 0.189894
R991 VP.n20 VP.n19 0.189894
R992 VP.n21 VP.n20 0.189894
R993 VP.n21 VP.n10 0.189894
R994 VP.n26 VP.n10 0.189894
R995 VP.n27 VP.n26 0.189894
R996 VP.n28 VP.n27 0.189894
R997 VP.n28 VP.n8 0.189894
R998 VP.n37 VP.n36 0.189894
R999 VP.n38 VP.n37 0.189894
R1000 VP.n38 VP.n6 0.189894
R1001 VP.n42 VP.n6 0.189894
R1002 VP.n43 VP.n42 0.189894
R1003 VP.n43 VP.n4 0.189894
R1004 VP.n47 VP.n4 0.189894
R1005 VP.n48 VP.n47 0.189894
R1006 VP.n49 VP.n48 0.189894
R1007 VP.n49 VP.n2 0.189894
R1008 VP.n54 VP.n2 0.189894
R1009 VP.n55 VP.n54 0.189894
R1010 VP.n56 VP.n55 0.189894
R1011 VP.n56 VP.n0 0.189894
R1012 VP VP.n60 0.153454
R1013 VDD1 VDD1.n0 176.453
R1014 VDD1.n3 VDD1.n2 176.339
R1015 VDD1.n3 VDD1.n1 176.339
R1016 VDD1.n5 VDD1.n4 175.299
R1017 VDD1.n5 VDD1.n3 36.1087
R1018 VDD1.n4 VDD1.t6 14.3199
R1019 VDD1.n4 VDD1.t7 14.3199
R1020 VDD1.n0 VDD1.t2 14.3199
R1021 VDD1.n0 VDD1.t5 14.3199
R1022 VDD1.n2 VDD1.t0 14.3199
R1023 VDD1.n2 VDD1.t1 14.3199
R1024 VDD1.n1 VDD1.t3 14.3199
R1025 VDD1.n1 VDD1.t4 14.3199
R1026 VDD1 VDD1.n5 1.03714
C0 VN B 1.01992f
C1 VTAIL B 1.60679f
C2 B w_n3510_n1422# 6.82386f
C3 VTAIL VN 2.87803f
C4 VN w_n3510_n1422# 6.86415f
C5 VDD2 VP 0.484329f
C6 VTAIL w_n3510_n1422# 1.91739f
C7 VDD1 VP 2.28272f
C8 VDD1 VDD2 1.57186f
C9 B VP 1.77912f
C10 VN VP 5.39253f
C11 VTAIL VP 2.89213f
C12 VP w_n3510_n1422# 7.31498f
C13 VDD2 B 1.3525f
C14 VN VDD2 1.95695f
C15 VTAIL VDD2 4.52736f
C16 VDD2 w_n3510_n1422# 1.65471f
C17 VDD1 B 1.26846f
C18 VDD1 VN 0.156213f
C19 VDD1 VTAIL 4.47556f
C20 VDD1 w_n3510_n1422# 1.55703f
C21 VDD2 VSUBS 1.054638f
C22 VDD1 VSUBS 1.865603f
C23 VTAIL VSUBS 0.50777f
C24 VN VSUBS 5.93342f
C25 VP VSUBS 2.606605f
C26 B VSUBS 3.52527f
C27 w_n3510_n1422# VSUBS 63.5591f
C28 VDD1.t2 VSUBS 0.045032f
C29 VDD1.t5 VSUBS 0.045032f
C30 VDD1.n0 VSUBS 0.21193f
C31 VDD1.t3 VSUBS 0.045032f
C32 VDD1.t4 VSUBS 0.045032f
C33 VDD1.n1 VSUBS 0.211517f
C34 VDD1.t0 VSUBS 0.045032f
C35 VDD1.t1 VSUBS 0.045032f
C36 VDD1.n2 VSUBS 0.211517f
C37 VDD1.n3 VSUBS 2.68916f
C38 VDD1.t6 VSUBS 0.045032f
C39 VDD1.t7 VSUBS 0.045032f
C40 VDD1.n4 VSUBS 0.20824f
C41 VDD1.n5 VSUBS 2.16933f
C42 VP.n0 VSUBS 0.073738f
C43 VP.t6 VSUBS 0.67086f
C44 VP.n1 VSUBS 0.046374f
C45 VP.n2 VSUBS 0.05593f
C46 VP.t7 VSUBS 0.67086f
C47 VP.n3 VSUBS 0.11116f
C48 VP.n4 VSUBS 0.05593f
C49 VP.t3 VSUBS 0.67086f
C50 VP.n5 VSUBS 0.313572f
C51 VP.n6 VSUBS 0.05593f
C52 VP.n7 VSUBS 0.108391f
C53 VP.n8 VSUBS 0.073738f
C54 VP.t0 VSUBS 0.67086f
C55 VP.n9 VSUBS 0.046374f
C56 VP.n10 VSUBS 0.05593f
C57 VP.t1 VSUBS 0.67086f
C58 VP.n11 VSUBS 0.11116f
C59 VP.n12 VSUBS 0.05593f
C60 VP.t2 VSUBS 0.67086f
C61 VP.n13 VSUBS 0.460121f
C62 VP.t5 VSUBS 1.02271f
C63 VP.n14 VSUBS 0.436394f
C64 VP.n15 VSUBS 0.476801f
C65 VP.n16 VSUBS 0.080566f
C66 VP.n17 VSUBS 0.11116f
C67 VP.n18 VSUBS 0.045214f
C68 VP.n19 VSUBS 0.05593f
C69 VP.n20 VSUBS 0.05593f
C70 VP.n21 VSUBS 0.05593f
C71 VP.n22 VSUBS 0.080566f
C72 VP.n23 VSUBS 0.313572f
C73 VP.n24 VSUBS 0.076449f
C74 VP.n25 VSUBS 0.112769f
C75 VP.n26 VSUBS 0.05593f
C76 VP.n27 VSUBS 0.05593f
C77 VP.n28 VSUBS 0.05593f
C78 VP.n29 VSUBS 0.108391f
C79 VP.n30 VSUBS 0.084683f
C80 VP.n31 VSUBS 0.487199f
C81 VP.n32 VSUBS 2.338f
C82 VP.n33 VSUBS 2.38621f
C83 VP.t4 VSUBS 0.67086f
C84 VP.n34 VSUBS 0.487199f
C85 VP.n35 VSUBS 0.084683f
C86 VP.n36 VSUBS 0.073738f
C87 VP.n37 VSUBS 0.05593f
C88 VP.n38 VSUBS 0.05593f
C89 VP.n39 VSUBS 0.046374f
C90 VP.n40 VSUBS 0.112769f
C91 VP.n41 VSUBS 0.076449f
C92 VP.n42 VSUBS 0.05593f
C93 VP.n43 VSUBS 0.05593f
C94 VP.n44 VSUBS 0.080566f
C95 VP.n45 VSUBS 0.11116f
C96 VP.n46 VSUBS 0.045214f
C97 VP.n47 VSUBS 0.05593f
C98 VP.n48 VSUBS 0.05593f
C99 VP.n49 VSUBS 0.05593f
C100 VP.n50 VSUBS 0.080566f
C101 VP.n51 VSUBS 0.313572f
C102 VP.n52 VSUBS 0.076449f
C103 VP.n53 VSUBS 0.112769f
C104 VP.n54 VSUBS 0.05593f
C105 VP.n55 VSUBS 0.05593f
C106 VP.n56 VSUBS 0.05593f
C107 VP.n57 VSUBS 0.108391f
C108 VP.n58 VSUBS 0.084683f
C109 VP.n59 VSUBS 0.487199f
C110 VP.n60 VSUBS 0.077406f
C111 B.n0 VSUBS 0.007327f
C112 B.n1 VSUBS 0.007327f
C113 B.n2 VSUBS 0.010837f
C114 B.n3 VSUBS 0.008304f
C115 B.n4 VSUBS 0.008304f
C116 B.n5 VSUBS 0.008304f
C117 B.n6 VSUBS 0.008304f
C118 B.n7 VSUBS 0.008304f
C119 B.n8 VSUBS 0.008304f
C120 B.n9 VSUBS 0.008304f
C121 B.n10 VSUBS 0.008304f
C122 B.n11 VSUBS 0.008304f
C123 B.n12 VSUBS 0.008304f
C124 B.n13 VSUBS 0.008304f
C125 B.n14 VSUBS 0.008304f
C126 B.n15 VSUBS 0.008304f
C127 B.n16 VSUBS 0.008304f
C128 B.n17 VSUBS 0.008304f
C129 B.n18 VSUBS 0.008304f
C130 B.n19 VSUBS 0.008304f
C131 B.n20 VSUBS 0.008304f
C132 B.n21 VSUBS 0.008304f
C133 B.n22 VSUBS 0.008304f
C134 B.n23 VSUBS 0.008304f
C135 B.n24 VSUBS 0.01765f
C136 B.n25 VSUBS 0.008304f
C137 B.n26 VSUBS 0.008304f
C138 B.n27 VSUBS 0.008304f
C139 B.n28 VSUBS 0.008304f
C140 B.n29 VSUBS 0.008304f
C141 B.n30 VSUBS 0.008304f
C142 B.n31 VSUBS 0.008304f
C143 B.t4 VSUBS 0.059725f
C144 B.t5 VSUBS 0.072599f
C145 B.t3 VSUBS 0.2911f
C146 B.n32 VSUBS 0.084619f
C147 B.n33 VSUBS 0.070126f
C148 B.n34 VSUBS 0.008304f
C149 B.n35 VSUBS 0.008304f
C150 B.n36 VSUBS 0.008304f
C151 B.n37 VSUBS 0.008304f
C152 B.t10 VSUBS 0.059725f
C153 B.t11 VSUBS 0.072599f
C154 B.t9 VSUBS 0.2911f
C155 B.n38 VSUBS 0.084619f
C156 B.n39 VSUBS 0.070126f
C157 B.n40 VSUBS 0.01924f
C158 B.n41 VSUBS 0.008304f
C159 B.n42 VSUBS 0.008304f
C160 B.n43 VSUBS 0.008304f
C161 B.n44 VSUBS 0.008304f
C162 B.n45 VSUBS 0.008304f
C163 B.n46 VSUBS 0.008304f
C164 B.n47 VSUBS 0.01765f
C165 B.n48 VSUBS 0.008304f
C166 B.n49 VSUBS 0.008304f
C167 B.n50 VSUBS 0.008304f
C168 B.n51 VSUBS 0.008304f
C169 B.n52 VSUBS 0.008304f
C170 B.n53 VSUBS 0.008304f
C171 B.n54 VSUBS 0.008304f
C172 B.n55 VSUBS 0.008304f
C173 B.n56 VSUBS 0.008304f
C174 B.n57 VSUBS 0.008304f
C175 B.n58 VSUBS 0.008304f
C176 B.n59 VSUBS 0.008304f
C177 B.n60 VSUBS 0.008304f
C178 B.n61 VSUBS 0.008304f
C179 B.n62 VSUBS 0.008304f
C180 B.n63 VSUBS 0.008304f
C181 B.n64 VSUBS 0.008304f
C182 B.n65 VSUBS 0.008304f
C183 B.n66 VSUBS 0.008304f
C184 B.n67 VSUBS 0.008304f
C185 B.n68 VSUBS 0.008304f
C186 B.n69 VSUBS 0.008304f
C187 B.n70 VSUBS 0.008304f
C188 B.n71 VSUBS 0.008304f
C189 B.n72 VSUBS 0.008304f
C190 B.n73 VSUBS 0.008304f
C191 B.n74 VSUBS 0.008304f
C192 B.n75 VSUBS 0.008304f
C193 B.n76 VSUBS 0.008304f
C194 B.n77 VSUBS 0.008304f
C195 B.n78 VSUBS 0.008304f
C196 B.n79 VSUBS 0.008304f
C197 B.n80 VSUBS 0.008304f
C198 B.n81 VSUBS 0.008304f
C199 B.n82 VSUBS 0.008304f
C200 B.n83 VSUBS 0.008304f
C201 B.n84 VSUBS 0.008304f
C202 B.n85 VSUBS 0.008304f
C203 B.n86 VSUBS 0.008304f
C204 B.n87 VSUBS 0.008304f
C205 B.n88 VSUBS 0.008304f
C206 B.n89 VSUBS 0.008304f
C207 B.n90 VSUBS 0.008304f
C208 B.n91 VSUBS 0.008304f
C209 B.n92 VSUBS 0.008304f
C210 B.n93 VSUBS 0.018987f
C211 B.n94 VSUBS 0.008304f
C212 B.n95 VSUBS 0.008304f
C213 B.n96 VSUBS 0.008304f
C214 B.n97 VSUBS 0.008304f
C215 B.n98 VSUBS 0.008304f
C216 B.n99 VSUBS 0.008304f
C217 B.t8 VSUBS 0.059725f
C218 B.t7 VSUBS 0.072599f
C219 B.t6 VSUBS 0.2911f
C220 B.n100 VSUBS 0.084619f
C221 B.n101 VSUBS 0.070126f
C222 B.n102 VSUBS 0.008304f
C223 B.n103 VSUBS 0.008304f
C224 B.n104 VSUBS 0.008304f
C225 B.n105 VSUBS 0.008304f
C226 B.n106 VSUBS 0.004641f
C227 B.n107 VSUBS 0.008304f
C228 B.n108 VSUBS 0.008304f
C229 B.n109 VSUBS 0.008304f
C230 B.n110 VSUBS 0.008304f
C231 B.n111 VSUBS 0.008304f
C232 B.n112 VSUBS 0.008304f
C233 B.n113 VSUBS 0.01765f
C234 B.n114 VSUBS 0.008304f
C235 B.n115 VSUBS 0.008304f
C236 B.n116 VSUBS 0.008304f
C237 B.n117 VSUBS 0.008304f
C238 B.n118 VSUBS 0.008304f
C239 B.n119 VSUBS 0.008304f
C240 B.n120 VSUBS 0.008304f
C241 B.n121 VSUBS 0.008304f
C242 B.n122 VSUBS 0.008304f
C243 B.n123 VSUBS 0.008304f
C244 B.n124 VSUBS 0.008304f
C245 B.n125 VSUBS 0.008304f
C246 B.n126 VSUBS 0.008304f
C247 B.n127 VSUBS 0.008304f
C248 B.n128 VSUBS 0.008304f
C249 B.n129 VSUBS 0.008304f
C250 B.n130 VSUBS 0.008304f
C251 B.n131 VSUBS 0.008304f
C252 B.n132 VSUBS 0.008304f
C253 B.n133 VSUBS 0.008304f
C254 B.n134 VSUBS 0.008304f
C255 B.n135 VSUBS 0.008304f
C256 B.n136 VSUBS 0.008304f
C257 B.n137 VSUBS 0.008304f
C258 B.n138 VSUBS 0.008304f
C259 B.n139 VSUBS 0.008304f
C260 B.n140 VSUBS 0.008304f
C261 B.n141 VSUBS 0.008304f
C262 B.n142 VSUBS 0.008304f
C263 B.n143 VSUBS 0.008304f
C264 B.n144 VSUBS 0.008304f
C265 B.n145 VSUBS 0.008304f
C266 B.n146 VSUBS 0.008304f
C267 B.n147 VSUBS 0.008304f
C268 B.n148 VSUBS 0.008304f
C269 B.n149 VSUBS 0.008304f
C270 B.n150 VSUBS 0.008304f
C271 B.n151 VSUBS 0.008304f
C272 B.n152 VSUBS 0.008304f
C273 B.n153 VSUBS 0.008304f
C274 B.n154 VSUBS 0.008304f
C275 B.n155 VSUBS 0.008304f
C276 B.n156 VSUBS 0.008304f
C277 B.n157 VSUBS 0.008304f
C278 B.n158 VSUBS 0.008304f
C279 B.n159 VSUBS 0.008304f
C280 B.n160 VSUBS 0.008304f
C281 B.n161 VSUBS 0.008304f
C282 B.n162 VSUBS 0.008304f
C283 B.n163 VSUBS 0.008304f
C284 B.n164 VSUBS 0.008304f
C285 B.n165 VSUBS 0.008304f
C286 B.n166 VSUBS 0.008304f
C287 B.n167 VSUBS 0.008304f
C288 B.n168 VSUBS 0.008304f
C289 B.n169 VSUBS 0.008304f
C290 B.n170 VSUBS 0.008304f
C291 B.n171 VSUBS 0.008304f
C292 B.n172 VSUBS 0.008304f
C293 B.n173 VSUBS 0.008304f
C294 B.n174 VSUBS 0.008304f
C295 B.n175 VSUBS 0.008304f
C296 B.n176 VSUBS 0.008304f
C297 B.n177 VSUBS 0.008304f
C298 B.n178 VSUBS 0.008304f
C299 B.n179 VSUBS 0.008304f
C300 B.n180 VSUBS 0.008304f
C301 B.n181 VSUBS 0.008304f
C302 B.n182 VSUBS 0.008304f
C303 B.n183 VSUBS 0.008304f
C304 B.n184 VSUBS 0.008304f
C305 B.n185 VSUBS 0.008304f
C306 B.n186 VSUBS 0.008304f
C307 B.n187 VSUBS 0.008304f
C308 B.n188 VSUBS 0.008304f
C309 B.n189 VSUBS 0.008304f
C310 B.n190 VSUBS 0.008304f
C311 B.n191 VSUBS 0.008304f
C312 B.n192 VSUBS 0.008304f
C313 B.n193 VSUBS 0.008304f
C314 B.n194 VSUBS 0.008304f
C315 B.n195 VSUBS 0.008304f
C316 B.n196 VSUBS 0.008304f
C317 B.n197 VSUBS 0.008304f
C318 B.n198 VSUBS 0.008304f
C319 B.n199 VSUBS 0.008304f
C320 B.n200 VSUBS 0.01765f
C321 B.n201 VSUBS 0.018987f
C322 B.n202 VSUBS 0.018987f
C323 B.n203 VSUBS 0.008304f
C324 B.n204 VSUBS 0.008304f
C325 B.n205 VSUBS 0.008304f
C326 B.n206 VSUBS 0.008304f
C327 B.n207 VSUBS 0.008304f
C328 B.n208 VSUBS 0.008304f
C329 B.n209 VSUBS 0.008304f
C330 B.n210 VSUBS 0.008304f
C331 B.n211 VSUBS 0.008304f
C332 B.n212 VSUBS 0.008304f
C333 B.n213 VSUBS 0.008304f
C334 B.n214 VSUBS 0.008304f
C335 B.n215 VSUBS 0.008304f
C336 B.n216 VSUBS 0.008304f
C337 B.n217 VSUBS 0.008304f
C338 B.n218 VSUBS 0.008304f
C339 B.t2 VSUBS 0.059725f
C340 B.t1 VSUBS 0.072599f
C341 B.t0 VSUBS 0.2911f
C342 B.n219 VSUBS 0.084619f
C343 B.n220 VSUBS 0.070126f
C344 B.n221 VSUBS 0.01924f
C345 B.n222 VSUBS 0.007816f
C346 B.n223 VSUBS 0.008304f
C347 B.n224 VSUBS 0.008304f
C348 B.n225 VSUBS 0.008304f
C349 B.n226 VSUBS 0.008304f
C350 B.n227 VSUBS 0.008304f
C351 B.n228 VSUBS 0.008304f
C352 B.n229 VSUBS 0.008304f
C353 B.n230 VSUBS 0.008304f
C354 B.n231 VSUBS 0.008304f
C355 B.n232 VSUBS 0.008304f
C356 B.n233 VSUBS 0.008304f
C357 B.n234 VSUBS 0.008304f
C358 B.n235 VSUBS 0.008304f
C359 B.n236 VSUBS 0.008304f
C360 B.n237 VSUBS 0.008304f
C361 B.n238 VSUBS 0.004641f
C362 B.n239 VSUBS 0.01924f
C363 B.n240 VSUBS 0.007816f
C364 B.n241 VSUBS 0.008304f
C365 B.n242 VSUBS 0.008304f
C366 B.n243 VSUBS 0.008304f
C367 B.n244 VSUBS 0.008304f
C368 B.n245 VSUBS 0.008304f
C369 B.n246 VSUBS 0.008304f
C370 B.n247 VSUBS 0.008304f
C371 B.n248 VSUBS 0.008304f
C372 B.n249 VSUBS 0.008304f
C373 B.n250 VSUBS 0.008304f
C374 B.n251 VSUBS 0.008304f
C375 B.n252 VSUBS 0.008304f
C376 B.n253 VSUBS 0.008304f
C377 B.n254 VSUBS 0.008304f
C378 B.n255 VSUBS 0.008304f
C379 B.n256 VSUBS 0.008304f
C380 B.n257 VSUBS 0.008304f
C381 B.n258 VSUBS 0.017912f
C382 B.n259 VSUBS 0.018725f
C383 B.n260 VSUBS 0.01765f
C384 B.n261 VSUBS 0.008304f
C385 B.n262 VSUBS 0.008304f
C386 B.n263 VSUBS 0.008304f
C387 B.n264 VSUBS 0.008304f
C388 B.n265 VSUBS 0.008304f
C389 B.n266 VSUBS 0.008304f
C390 B.n267 VSUBS 0.008304f
C391 B.n268 VSUBS 0.008304f
C392 B.n269 VSUBS 0.008304f
C393 B.n270 VSUBS 0.008304f
C394 B.n271 VSUBS 0.008304f
C395 B.n272 VSUBS 0.008304f
C396 B.n273 VSUBS 0.008304f
C397 B.n274 VSUBS 0.008304f
C398 B.n275 VSUBS 0.008304f
C399 B.n276 VSUBS 0.008304f
C400 B.n277 VSUBS 0.008304f
C401 B.n278 VSUBS 0.008304f
C402 B.n279 VSUBS 0.008304f
C403 B.n280 VSUBS 0.008304f
C404 B.n281 VSUBS 0.008304f
C405 B.n282 VSUBS 0.008304f
C406 B.n283 VSUBS 0.008304f
C407 B.n284 VSUBS 0.008304f
C408 B.n285 VSUBS 0.008304f
C409 B.n286 VSUBS 0.008304f
C410 B.n287 VSUBS 0.008304f
C411 B.n288 VSUBS 0.008304f
C412 B.n289 VSUBS 0.008304f
C413 B.n290 VSUBS 0.008304f
C414 B.n291 VSUBS 0.008304f
C415 B.n292 VSUBS 0.008304f
C416 B.n293 VSUBS 0.008304f
C417 B.n294 VSUBS 0.008304f
C418 B.n295 VSUBS 0.008304f
C419 B.n296 VSUBS 0.008304f
C420 B.n297 VSUBS 0.008304f
C421 B.n298 VSUBS 0.008304f
C422 B.n299 VSUBS 0.008304f
C423 B.n300 VSUBS 0.008304f
C424 B.n301 VSUBS 0.008304f
C425 B.n302 VSUBS 0.008304f
C426 B.n303 VSUBS 0.008304f
C427 B.n304 VSUBS 0.008304f
C428 B.n305 VSUBS 0.008304f
C429 B.n306 VSUBS 0.008304f
C430 B.n307 VSUBS 0.008304f
C431 B.n308 VSUBS 0.008304f
C432 B.n309 VSUBS 0.008304f
C433 B.n310 VSUBS 0.008304f
C434 B.n311 VSUBS 0.008304f
C435 B.n312 VSUBS 0.008304f
C436 B.n313 VSUBS 0.008304f
C437 B.n314 VSUBS 0.008304f
C438 B.n315 VSUBS 0.008304f
C439 B.n316 VSUBS 0.008304f
C440 B.n317 VSUBS 0.008304f
C441 B.n318 VSUBS 0.008304f
C442 B.n319 VSUBS 0.008304f
C443 B.n320 VSUBS 0.008304f
C444 B.n321 VSUBS 0.008304f
C445 B.n322 VSUBS 0.008304f
C446 B.n323 VSUBS 0.008304f
C447 B.n324 VSUBS 0.008304f
C448 B.n325 VSUBS 0.008304f
C449 B.n326 VSUBS 0.008304f
C450 B.n327 VSUBS 0.008304f
C451 B.n328 VSUBS 0.008304f
C452 B.n329 VSUBS 0.008304f
C453 B.n330 VSUBS 0.008304f
C454 B.n331 VSUBS 0.008304f
C455 B.n332 VSUBS 0.008304f
C456 B.n333 VSUBS 0.008304f
C457 B.n334 VSUBS 0.008304f
C458 B.n335 VSUBS 0.008304f
C459 B.n336 VSUBS 0.008304f
C460 B.n337 VSUBS 0.008304f
C461 B.n338 VSUBS 0.008304f
C462 B.n339 VSUBS 0.008304f
C463 B.n340 VSUBS 0.008304f
C464 B.n341 VSUBS 0.008304f
C465 B.n342 VSUBS 0.008304f
C466 B.n343 VSUBS 0.008304f
C467 B.n344 VSUBS 0.008304f
C468 B.n345 VSUBS 0.008304f
C469 B.n346 VSUBS 0.008304f
C470 B.n347 VSUBS 0.008304f
C471 B.n348 VSUBS 0.008304f
C472 B.n349 VSUBS 0.008304f
C473 B.n350 VSUBS 0.008304f
C474 B.n351 VSUBS 0.008304f
C475 B.n352 VSUBS 0.008304f
C476 B.n353 VSUBS 0.008304f
C477 B.n354 VSUBS 0.008304f
C478 B.n355 VSUBS 0.008304f
C479 B.n356 VSUBS 0.008304f
C480 B.n357 VSUBS 0.008304f
C481 B.n358 VSUBS 0.008304f
C482 B.n359 VSUBS 0.008304f
C483 B.n360 VSUBS 0.008304f
C484 B.n361 VSUBS 0.008304f
C485 B.n362 VSUBS 0.008304f
C486 B.n363 VSUBS 0.008304f
C487 B.n364 VSUBS 0.008304f
C488 B.n365 VSUBS 0.008304f
C489 B.n366 VSUBS 0.008304f
C490 B.n367 VSUBS 0.008304f
C491 B.n368 VSUBS 0.008304f
C492 B.n369 VSUBS 0.008304f
C493 B.n370 VSUBS 0.008304f
C494 B.n371 VSUBS 0.008304f
C495 B.n372 VSUBS 0.008304f
C496 B.n373 VSUBS 0.008304f
C497 B.n374 VSUBS 0.008304f
C498 B.n375 VSUBS 0.008304f
C499 B.n376 VSUBS 0.008304f
C500 B.n377 VSUBS 0.008304f
C501 B.n378 VSUBS 0.008304f
C502 B.n379 VSUBS 0.008304f
C503 B.n380 VSUBS 0.008304f
C504 B.n381 VSUBS 0.008304f
C505 B.n382 VSUBS 0.008304f
C506 B.n383 VSUBS 0.008304f
C507 B.n384 VSUBS 0.008304f
C508 B.n385 VSUBS 0.008304f
C509 B.n386 VSUBS 0.008304f
C510 B.n387 VSUBS 0.008304f
C511 B.n388 VSUBS 0.008304f
C512 B.n389 VSUBS 0.008304f
C513 B.n390 VSUBS 0.008304f
C514 B.n391 VSUBS 0.008304f
C515 B.n392 VSUBS 0.008304f
C516 B.n393 VSUBS 0.008304f
C517 B.n394 VSUBS 0.008304f
C518 B.n395 VSUBS 0.008304f
C519 B.n396 VSUBS 0.01765f
C520 B.n397 VSUBS 0.018987f
C521 B.n398 VSUBS 0.018987f
C522 B.n399 VSUBS 0.008304f
C523 B.n400 VSUBS 0.008304f
C524 B.n401 VSUBS 0.008304f
C525 B.n402 VSUBS 0.008304f
C526 B.n403 VSUBS 0.008304f
C527 B.n404 VSUBS 0.008304f
C528 B.n405 VSUBS 0.008304f
C529 B.n406 VSUBS 0.008304f
C530 B.n407 VSUBS 0.008304f
C531 B.n408 VSUBS 0.008304f
C532 B.n409 VSUBS 0.008304f
C533 B.n410 VSUBS 0.008304f
C534 B.n411 VSUBS 0.008304f
C535 B.n412 VSUBS 0.008304f
C536 B.n413 VSUBS 0.008304f
C537 B.n414 VSUBS 0.008304f
C538 B.n415 VSUBS 0.007816f
C539 B.n416 VSUBS 0.008304f
C540 B.n417 VSUBS 0.008304f
C541 B.n418 VSUBS 0.004641f
C542 B.n419 VSUBS 0.008304f
C543 B.n420 VSUBS 0.008304f
C544 B.n421 VSUBS 0.008304f
C545 B.n422 VSUBS 0.008304f
C546 B.n423 VSUBS 0.008304f
C547 B.n424 VSUBS 0.008304f
C548 B.n425 VSUBS 0.008304f
C549 B.n426 VSUBS 0.008304f
C550 B.n427 VSUBS 0.008304f
C551 B.n428 VSUBS 0.008304f
C552 B.n429 VSUBS 0.008304f
C553 B.n430 VSUBS 0.008304f
C554 B.n431 VSUBS 0.004641f
C555 B.n432 VSUBS 0.01924f
C556 B.n433 VSUBS 0.007816f
C557 B.n434 VSUBS 0.008304f
C558 B.n435 VSUBS 0.008304f
C559 B.n436 VSUBS 0.008304f
C560 B.n437 VSUBS 0.008304f
C561 B.n438 VSUBS 0.008304f
C562 B.n439 VSUBS 0.008304f
C563 B.n440 VSUBS 0.008304f
C564 B.n441 VSUBS 0.008304f
C565 B.n442 VSUBS 0.008304f
C566 B.n443 VSUBS 0.008304f
C567 B.n444 VSUBS 0.008304f
C568 B.n445 VSUBS 0.008304f
C569 B.n446 VSUBS 0.008304f
C570 B.n447 VSUBS 0.008304f
C571 B.n448 VSUBS 0.008304f
C572 B.n449 VSUBS 0.008304f
C573 B.n450 VSUBS 0.008304f
C574 B.n451 VSUBS 0.018987f
C575 B.n452 VSUBS 0.018987f
C576 B.n453 VSUBS 0.01765f
C577 B.n454 VSUBS 0.008304f
C578 B.n455 VSUBS 0.008304f
C579 B.n456 VSUBS 0.008304f
C580 B.n457 VSUBS 0.008304f
C581 B.n458 VSUBS 0.008304f
C582 B.n459 VSUBS 0.008304f
C583 B.n460 VSUBS 0.008304f
C584 B.n461 VSUBS 0.008304f
C585 B.n462 VSUBS 0.008304f
C586 B.n463 VSUBS 0.008304f
C587 B.n464 VSUBS 0.008304f
C588 B.n465 VSUBS 0.008304f
C589 B.n466 VSUBS 0.008304f
C590 B.n467 VSUBS 0.008304f
C591 B.n468 VSUBS 0.008304f
C592 B.n469 VSUBS 0.008304f
C593 B.n470 VSUBS 0.008304f
C594 B.n471 VSUBS 0.008304f
C595 B.n472 VSUBS 0.008304f
C596 B.n473 VSUBS 0.008304f
C597 B.n474 VSUBS 0.008304f
C598 B.n475 VSUBS 0.008304f
C599 B.n476 VSUBS 0.008304f
C600 B.n477 VSUBS 0.008304f
C601 B.n478 VSUBS 0.008304f
C602 B.n479 VSUBS 0.008304f
C603 B.n480 VSUBS 0.008304f
C604 B.n481 VSUBS 0.008304f
C605 B.n482 VSUBS 0.008304f
C606 B.n483 VSUBS 0.008304f
C607 B.n484 VSUBS 0.008304f
C608 B.n485 VSUBS 0.008304f
C609 B.n486 VSUBS 0.008304f
C610 B.n487 VSUBS 0.008304f
C611 B.n488 VSUBS 0.008304f
C612 B.n489 VSUBS 0.008304f
C613 B.n490 VSUBS 0.008304f
C614 B.n491 VSUBS 0.008304f
C615 B.n492 VSUBS 0.008304f
C616 B.n493 VSUBS 0.008304f
C617 B.n494 VSUBS 0.008304f
C618 B.n495 VSUBS 0.008304f
C619 B.n496 VSUBS 0.008304f
C620 B.n497 VSUBS 0.008304f
C621 B.n498 VSUBS 0.008304f
C622 B.n499 VSUBS 0.008304f
C623 B.n500 VSUBS 0.008304f
C624 B.n501 VSUBS 0.008304f
C625 B.n502 VSUBS 0.008304f
C626 B.n503 VSUBS 0.008304f
C627 B.n504 VSUBS 0.008304f
C628 B.n505 VSUBS 0.008304f
C629 B.n506 VSUBS 0.008304f
C630 B.n507 VSUBS 0.008304f
C631 B.n508 VSUBS 0.008304f
C632 B.n509 VSUBS 0.008304f
C633 B.n510 VSUBS 0.008304f
C634 B.n511 VSUBS 0.008304f
C635 B.n512 VSUBS 0.008304f
C636 B.n513 VSUBS 0.008304f
C637 B.n514 VSUBS 0.008304f
C638 B.n515 VSUBS 0.008304f
C639 B.n516 VSUBS 0.008304f
C640 B.n517 VSUBS 0.008304f
C641 B.n518 VSUBS 0.008304f
C642 B.n519 VSUBS 0.010837f
C643 B.n520 VSUBS 0.011544f
C644 B.n521 VSUBS 0.022956f
C645 VTAIL.t14 VSUBS 0.053176f
C646 VTAIL.t9 VSUBS 0.053176f
C647 VTAIL.n0 VSUBS 0.211217f
C648 VTAIL.n1 VSUBS 0.544612f
C649 VTAIL.t15 VSUBS 0.331148f
C650 VTAIL.n2 VSUBS 0.609025f
C651 VTAIL.t3 VSUBS 0.331148f
C652 VTAIL.n3 VSUBS 0.609025f
C653 VTAIL.t0 VSUBS 0.053176f
C654 VTAIL.t4 VSUBS 0.053176f
C655 VTAIL.n4 VSUBS 0.211217f
C656 VTAIL.n5 VSUBS 0.748208f
C657 VTAIL.t1 VSUBS 0.331148f
C658 VTAIL.n6 VSUBS 1.3629f
C659 VTAIL.t13 VSUBS 0.331149f
C660 VTAIL.n7 VSUBS 1.3629f
C661 VTAIL.t11 VSUBS 0.053176f
C662 VTAIL.t12 VSUBS 0.053176f
C663 VTAIL.n8 VSUBS 0.211217f
C664 VTAIL.n9 VSUBS 0.748207f
C665 VTAIL.t10 VSUBS 0.331149f
C666 VTAIL.n10 VSUBS 0.609024f
C667 VTAIL.t2 VSUBS 0.331149f
C668 VTAIL.n11 VSUBS 0.609024f
C669 VTAIL.t5 VSUBS 0.053176f
C670 VTAIL.t7 VSUBS 0.053176f
C671 VTAIL.n12 VSUBS 0.211217f
C672 VTAIL.n13 VSUBS 0.748207f
C673 VTAIL.t6 VSUBS 0.331148f
C674 VTAIL.n14 VSUBS 1.3629f
C675 VTAIL.t8 VSUBS 0.331148f
C676 VTAIL.n15 VSUBS 1.35734f
C677 VDD2.t7 VSUBS 0.030212f
C678 VDD2.t6 VSUBS 0.030212f
C679 VDD2.n0 VSUBS 0.14191f
C680 VDD2.t2 VSUBS 0.030212f
C681 VDD2.t1 VSUBS 0.030212f
C682 VDD2.n1 VSUBS 0.14191f
C683 VDD2.n2 VSUBS 1.76881f
C684 VDD2.t4 VSUBS 0.030212f
C685 VDD2.t5 VSUBS 0.030212f
C686 VDD2.n3 VSUBS 0.139711f
C687 VDD2.n4 VSUBS 1.43492f
C688 VDD2.t0 VSUBS 0.030212f
C689 VDD2.t3 VSUBS 0.030212f
C690 VDD2.n5 VSUBS 0.1419f
C691 VN.n0 VSUBS 0.062342f
C692 VN.t7 VSUBS 0.567178f
C693 VN.n1 VSUBS 0.039207f
C694 VN.n2 VSUBS 0.047286f
C695 VN.t6 VSUBS 0.567178f
C696 VN.n3 VSUBS 0.09398f
C697 VN.n4 VSUBS 0.047286f
C698 VN.t1 VSUBS 0.567178f
C699 VN.n5 VSUBS 0.389008f
C700 VN.t0 VSUBS 0.86465f
C701 VN.n6 VSUBS 0.368949f
C702 VN.n7 VSUBS 0.403111f
C703 VN.n8 VSUBS 0.068115f
C704 VN.n9 VSUBS 0.09398f
C705 VN.n10 VSUBS 0.038226f
C706 VN.n11 VSUBS 0.047286f
C707 VN.n12 VSUBS 0.047286f
C708 VN.n13 VSUBS 0.047286f
C709 VN.n14 VSUBS 0.068115f
C710 VN.n15 VSUBS 0.265109f
C711 VN.n16 VSUBS 0.064634f
C712 VN.n17 VSUBS 0.095341f
C713 VN.n18 VSUBS 0.047286f
C714 VN.n19 VSUBS 0.047286f
C715 VN.n20 VSUBS 0.047286f
C716 VN.n21 VSUBS 0.091639f
C717 VN.n22 VSUBS 0.071595f
C718 VN.n23 VSUBS 0.411902f
C719 VN.n24 VSUBS 0.065443f
C720 VN.n25 VSUBS 0.062342f
C721 VN.t2 VSUBS 0.567178f
C722 VN.n26 VSUBS 0.039207f
C723 VN.n27 VSUBS 0.047286f
C724 VN.t4 VSUBS 0.567178f
C725 VN.n28 VSUBS 0.09398f
C726 VN.n29 VSUBS 0.047286f
C727 VN.t3 VSUBS 0.567178f
C728 VN.n30 VSUBS 0.389008f
C729 VN.t5 VSUBS 0.86465f
C730 VN.n31 VSUBS 0.368949f
C731 VN.n32 VSUBS 0.403111f
C732 VN.n33 VSUBS 0.068115f
C733 VN.n34 VSUBS 0.09398f
C734 VN.n35 VSUBS 0.038226f
C735 VN.n36 VSUBS 0.047286f
C736 VN.n37 VSUBS 0.047286f
C737 VN.n38 VSUBS 0.047286f
C738 VN.n39 VSUBS 0.068115f
C739 VN.n40 VSUBS 0.265109f
C740 VN.n41 VSUBS 0.064634f
C741 VN.n42 VSUBS 0.095341f
C742 VN.n43 VSUBS 0.047286f
C743 VN.n44 VSUBS 0.047286f
C744 VN.n45 VSUBS 0.047286f
C745 VN.n46 VSUBS 0.091639f
C746 VN.n47 VSUBS 0.071595f
C747 VN.n48 VSUBS 0.411902f
C748 VN.n49 VSUBS 2.00287f
.ends

