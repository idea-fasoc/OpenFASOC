* NGSPICE file created from diff_pair_sample_0485.ext - technology: sky130A

.subckt diff_pair_sample_0485 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t19 VP.t0 VDD1.t1 B.t6 sky130_fd_pr__nfet_01v8 ad=2.9007 pd=17.91 as=2.9007 ps=17.91 w=17.58 l=3.12
X1 VDD2.t9 VN.t0 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=2.9007 pd=17.91 as=2.9007 ps=17.91 w=17.58 l=3.12
X2 VTAIL.t4 VN.t1 VDD2.t8 B.t4 sky130_fd_pr__nfet_01v8 ad=2.9007 pd=17.91 as=2.9007 ps=17.91 w=17.58 l=3.12
X3 VTAIL.t18 VP.t1 VDD1.t0 B.t4 sky130_fd_pr__nfet_01v8 ad=2.9007 pd=17.91 as=2.9007 ps=17.91 w=17.58 l=3.12
X4 VDD2.t7 VN.t2 VTAIL.t8 B.t8 sky130_fd_pr__nfet_01v8 ad=6.8562 pd=35.94 as=2.9007 ps=17.91 w=17.58 l=3.12
X5 VDD1.t3 VP.t2 VTAIL.t17 B.t1 sky130_fd_pr__nfet_01v8 ad=2.9007 pd=17.91 as=6.8562 ps=35.94 w=17.58 l=3.12
X6 VDD1.t2 VP.t3 VTAIL.t16 B.t0 sky130_fd_pr__nfet_01v8 ad=2.9007 pd=17.91 as=2.9007 ps=17.91 w=17.58 l=3.12
X7 VDD2.t6 VN.t3 VTAIL.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=6.8562 pd=35.94 as=2.9007 ps=17.91 w=17.58 l=3.12
X8 VDD1.t9 VP.t4 VTAIL.t15 B.t8 sky130_fd_pr__nfet_01v8 ad=6.8562 pd=35.94 as=2.9007 ps=17.91 w=17.58 l=3.12
X9 B.t23 B.t21 B.t22 B.t11 sky130_fd_pr__nfet_01v8 ad=6.8562 pd=35.94 as=0 ps=0 w=17.58 l=3.12
X10 VDD2.t5 VN.t4 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=2.9007 pd=17.91 as=2.9007 ps=17.91 w=17.58 l=3.12
X11 B.t20 B.t18 B.t19 B.t15 sky130_fd_pr__nfet_01v8 ad=6.8562 pd=35.94 as=0 ps=0 w=17.58 l=3.12
X12 VDD2.t4 VN.t5 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=2.9007 pd=17.91 as=6.8562 ps=35.94 w=17.58 l=3.12
X13 VDD2.t3 VN.t6 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=2.9007 pd=17.91 as=6.8562 ps=35.94 w=17.58 l=3.12
X14 VTAIL.t9 VN.t7 VDD2.t2 B.t9 sky130_fd_pr__nfet_01v8 ad=2.9007 pd=17.91 as=2.9007 ps=17.91 w=17.58 l=3.12
X15 VTAIL.t14 VP.t5 VDD1.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=2.9007 pd=17.91 as=2.9007 ps=17.91 w=17.58 l=3.12
X16 B.t17 B.t14 B.t16 B.t15 sky130_fd_pr__nfet_01v8 ad=6.8562 pd=35.94 as=0 ps=0 w=17.58 l=3.12
X17 VDD1.t7 VP.t6 VTAIL.t13 B.t3 sky130_fd_pr__nfet_01v8 ad=2.9007 pd=17.91 as=2.9007 ps=17.91 w=17.58 l=3.12
X18 VDD1.t6 VP.t7 VTAIL.t12 B.t5 sky130_fd_pr__nfet_01v8 ad=6.8562 pd=35.94 as=2.9007 ps=17.91 w=17.58 l=3.12
X19 VTAIL.t11 VP.t8 VDD1.t5 B.t9 sky130_fd_pr__nfet_01v8 ad=2.9007 pd=17.91 as=2.9007 ps=17.91 w=17.58 l=3.12
X20 VTAIL.t7 VN.t8 VDD2.t1 B.t7 sky130_fd_pr__nfet_01v8 ad=2.9007 pd=17.91 as=2.9007 ps=17.91 w=17.58 l=3.12
X21 VTAIL.t6 VN.t9 VDD2.t0 B.t6 sky130_fd_pr__nfet_01v8 ad=2.9007 pd=17.91 as=2.9007 ps=17.91 w=17.58 l=3.12
X22 VDD1.t4 VP.t9 VTAIL.t10 B.t2 sky130_fd_pr__nfet_01v8 ad=2.9007 pd=17.91 as=6.8562 ps=35.94 w=17.58 l=3.12
X23 B.t13 B.t10 B.t12 B.t11 sky130_fd_pr__nfet_01v8 ad=6.8562 pd=35.94 as=0 ps=0 w=17.58 l=3.12
R0 VP.n26 VP.t7 169.263
R1 VP.n29 VP.n28 161.3
R2 VP.n30 VP.n25 161.3
R3 VP.n32 VP.n31 161.3
R4 VP.n33 VP.n24 161.3
R5 VP.n35 VP.n34 161.3
R6 VP.n36 VP.n23 161.3
R7 VP.n38 VP.n37 161.3
R8 VP.n39 VP.n22 161.3
R9 VP.n41 VP.n40 161.3
R10 VP.n42 VP.n21 161.3
R11 VP.n44 VP.n43 161.3
R12 VP.n45 VP.n20 161.3
R13 VP.n47 VP.n46 161.3
R14 VP.n49 VP.n48 161.3
R15 VP.n50 VP.n18 161.3
R16 VP.n52 VP.n51 161.3
R17 VP.n53 VP.n17 161.3
R18 VP.n55 VP.n54 161.3
R19 VP.n56 VP.n16 161.3
R20 VP.n58 VP.n57 161.3
R21 VP.n103 VP.n102 161.3
R22 VP.n101 VP.n1 161.3
R23 VP.n100 VP.n99 161.3
R24 VP.n98 VP.n2 161.3
R25 VP.n97 VP.n96 161.3
R26 VP.n95 VP.n3 161.3
R27 VP.n94 VP.n93 161.3
R28 VP.n92 VP.n91 161.3
R29 VP.n90 VP.n5 161.3
R30 VP.n89 VP.n88 161.3
R31 VP.n87 VP.n6 161.3
R32 VP.n86 VP.n85 161.3
R33 VP.n84 VP.n7 161.3
R34 VP.n83 VP.n82 161.3
R35 VP.n81 VP.n8 161.3
R36 VP.n80 VP.n79 161.3
R37 VP.n78 VP.n9 161.3
R38 VP.n77 VP.n76 161.3
R39 VP.n75 VP.n10 161.3
R40 VP.n74 VP.n73 161.3
R41 VP.n71 VP.n11 161.3
R42 VP.n70 VP.n69 161.3
R43 VP.n68 VP.n12 161.3
R44 VP.n67 VP.n66 161.3
R45 VP.n65 VP.n13 161.3
R46 VP.n64 VP.n63 161.3
R47 VP.n62 VP.n14 161.3
R48 VP.n83 VP.t3 135.794
R49 VP.n60 VP.t4 135.794
R50 VP.n72 VP.t5 135.794
R51 VP.n4 VP.t8 135.794
R52 VP.n0 VP.t2 135.794
R53 VP.n38 VP.t6 135.794
R54 VP.n15 VP.t9 135.794
R55 VP.n19 VP.t1 135.794
R56 VP.n27 VP.t0 135.794
R57 VP.n61 VP.n60 70.5721
R58 VP.n104 VP.n0 70.5721
R59 VP.n59 VP.n15 70.5721
R60 VP.n61 VP.n59 60.3139
R61 VP.n66 VP.n65 56.5617
R62 VP.n78 VP.n77 56.5617
R63 VP.n89 VP.n6 56.5617
R64 VP.n100 VP.n2 56.5617
R65 VP.n55 VP.n17 56.5617
R66 VP.n44 VP.n21 56.5617
R67 VP.n33 VP.n32 56.5617
R68 VP.n27 VP.n26 51.9472
R69 VP.n64 VP.n14 24.5923
R70 VP.n65 VP.n64 24.5923
R71 VP.n66 VP.n12 24.5923
R72 VP.n70 VP.n12 24.5923
R73 VP.n71 VP.n70 24.5923
R74 VP.n73 VP.n10 24.5923
R75 VP.n77 VP.n10 24.5923
R76 VP.n79 VP.n78 24.5923
R77 VP.n79 VP.n8 24.5923
R78 VP.n83 VP.n8 24.5923
R79 VP.n84 VP.n83 24.5923
R80 VP.n85 VP.n84 24.5923
R81 VP.n85 VP.n6 24.5923
R82 VP.n90 VP.n89 24.5923
R83 VP.n91 VP.n90 24.5923
R84 VP.n95 VP.n94 24.5923
R85 VP.n96 VP.n95 24.5923
R86 VP.n96 VP.n2 24.5923
R87 VP.n101 VP.n100 24.5923
R88 VP.n102 VP.n101 24.5923
R89 VP.n56 VP.n55 24.5923
R90 VP.n57 VP.n56 24.5923
R91 VP.n45 VP.n44 24.5923
R92 VP.n46 VP.n45 24.5923
R93 VP.n50 VP.n49 24.5923
R94 VP.n51 VP.n50 24.5923
R95 VP.n51 VP.n17 24.5923
R96 VP.n34 VP.n33 24.5923
R97 VP.n34 VP.n23 24.5923
R98 VP.n38 VP.n23 24.5923
R99 VP.n39 VP.n38 24.5923
R100 VP.n40 VP.n39 24.5923
R101 VP.n40 VP.n21 24.5923
R102 VP.n28 VP.n25 24.5923
R103 VP.n32 VP.n25 24.5923
R104 VP.n73 VP.n72 22.1332
R105 VP.n91 VP.n4 22.1332
R106 VP.n46 VP.n19 22.1332
R107 VP.n28 VP.n27 22.1332
R108 VP.n60 VP.n14 19.674
R109 VP.n102 VP.n0 19.674
R110 VP.n57 VP.n15 19.674
R111 VP.n29 VP.n26 3.92039
R112 VP.n72 VP.n71 2.45968
R113 VP.n94 VP.n4 2.45968
R114 VP.n49 VP.n19 2.45968
R115 VP.n59 VP.n58 0.354861
R116 VP.n62 VP.n61 0.354861
R117 VP.n104 VP.n103 0.354861
R118 VP VP.n104 0.267071
R119 VP.n30 VP.n29 0.189894
R120 VP.n31 VP.n30 0.189894
R121 VP.n31 VP.n24 0.189894
R122 VP.n35 VP.n24 0.189894
R123 VP.n36 VP.n35 0.189894
R124 VP.n37 VP.n36 0.189894
R125 VP.n37 VP.n22 0.189894
R126 VP.n41 VP.n22 0.189894
R127 VP.n42 VP.n41 0.189894
R128 VP.n43 VP.n42 0.189894
R129 VP.n43 VP.n20 0.189894
R130 VP.n47 VP.n20 0.189894
R131 VP.n48 VP.n47 0.189894
R132 VP.n48 VP.n18 0.189894
R133 VP.n52 VP.n18 0.189894
R134 VP.n53 VP.n52 0.189894
R135 VP.n54 VP.n53 0.189894
R136 VP.n54 VP.n16 0.189894
R137 VP.n58 VP.n16 0.189894
R138 VP.n63 VP.n62 0.189894
R139 VP.n63 VP.n13 0.189894
R140 VP.n67 VP.n13 0.189894
R141 VP.n68 VP.n67 0.189894
R142 VP.n69 VP.n68 0.189894
R143 VP.n69 VP.n11 0.189894
R144 VP.n74 VP.n11 0.189894
R145 VP.n75 VP.n74 0.189894
R146 VP.n76 VP.n75 0.189894
R147 VP.n76 VP.n9 0.189894
R148 VP.n80 VP.n9 0.189894
R149 VP.n81 VP.n80 0.189894
R150 VP.n82 VP.n81 0.189894
R151 VP.n82 VP.n7 0.189894
R152 VP.n86 VP.n7 0.189894
R153 VP.n87 VP.n86 0.189894
R154 VP.n88 VP.n87 0.189894
R155 VP.n88 VP.n5 0.189894
R156 VP.n92 VP.n5 0.189894
R157 VP.n93 VP.n92 0.189894
R158 VP.n93 VP.n3 0.189894
R159 VP.n97 VP.n3 0.189894
R160 VP.n98 VP.n97 0.189894
R161 VP.n99 VP.n98 0.189894
R162 VP.n99 VP.n1 0.189894
R163 VP.n103 VP.n1 0.189894
R164 VDD1.n92 VDD1.n0 289.615
R165 VDD1.n191 VDD1.n99 289.615
R166 VDD1.n93 VDD1.n92 185
R167 VDD1.n91 VDD1.n90 185
R168 VDD1.n4 VDD1.n3 185
R169 VDD1.n85 VDD1.n84 185
R170 VDD1.n83 VDD1.n82 185
R171 VDD1.n8 VDD1.n7 185
R172 VDD1.n12 VDD1.n10 185
R173 VDD1.n77 VDD1.n76 185
R174 VDD1.n75 VDD1.n74 185
R175 VDD1.n14 VDD1.n13 185
R176 VDD1.n69 VDD1.n68 185
R177 VDD1.n67 VDD1.n66 185
R178 VDD1.n18 VDD1.n17 185
R179 VDD1.n61 VDD1.n60 185
R180 VDD1.n59 VDD1.n58 185
R181 VDD1.n22 VDD1.n21 185
R182 VDD1.n53 VDD1.n52 185
R183 VDD1.n51 VDD1.n50 185
R184 VDD1.n26 VDD1.n25 185
R185 VDD1.n45 VDD1.n44 185
R186 VDD1.n43 VDD1.n42 185
R187 VDD1.n30 VDD1.n29 185
R188 VDD1.n37 VDD1.n36 185
R189 VDD1.n35 VDD1.n34 185
R190 VDD1.n132 VDD1.n131 185
R191 VDD1.n134 VDD1.n133 185
R192 VDD1.n127 VDD1.n126 185
R193 VDD1.n140 VDD1.n139 185
R194 VDD1.n142 VDD1.n141 185
R195 VDD1.n123 VDD1.n122 185
R196 VDD1.n148 VDD1.n147 185
R197 VDD1.n150 VDD1.n149 185
R198 VDD1.n119 VDD1.n118 185
R199 VDD1.n156 VDD1.n155 185
R200 VDD1.n158 VDD1.n157 185
R201 VDD1.n115 VDD1.n114 185
R202 VDD1.n164 VDD1.n163 185
R203 VDD1.n166 VDD1.n165 185
R204 VDD1.n111 VDD1.n110 185
R205 VDD1.n173 VDD1.n172 185
R206 VDD1.n174 VDD1.n109 185
R207 VDD1.n176 VDD1.n175 185
R208 VDD1.n107 VDD1.n106 185
R209 VDD1.n182 VDD1.n181 185
R210 VDD1.n184 VDD1.n183 185
R211 VDD1.n103 VDD1.n102 185
R212 VDD1.n190 VDD1.n189 185
R213 VDD1.n192 VDD1.n191 185
R214 VDD1.n33 VDD1.t6 147.659
R215 VDD1.n130 VDD1.t9 147.659
R216 VDD1.n92 VDD1.n91 104.615
R217 VDD1.n91 VDD1.n3 104.615
R218 VDD1.n84 VDD1.n3 104.615
R219 VDD1.n84 VDD1.n83 104.615
R220 VDD1.n83 VDD1.n7 104.615
R221 VDD1.n12 VDD1.n7 104.615
R222 VDD1.n76 VDD1.n12 104.615
R223 VDD1.n76 VDD1.n75 104.615
R224 VDD1.n75 VDD1.n13 104.615
R225 VDD1.n68 VDD1.n13 104.615
R226 VDD1.n68 VDD1.n67 104.615
R227 VDD1.n67 VDD1.n17 104.615
R228 VDD1.n60 VDD1.n17 104.615
R229 VDD1.n60 VDD1.n59 104.615
R230 VDD1.n59 VDD1.n21 104.615
R231 VDD1.n52 VDD1.n21 104.615
R232 VDD1.n52 VDD1.n51 104.615
R233 VDD1.n51 VDD1.n25 104.615
R234 VDD1.n44 VDD1.n25 104.615
R235 VDD1.n44 VDD1.n43 104.615
R236 VDD1.n43 VDD1.n29 104.615
R237 VDD1.n36 VDD1.n29 104.615
R238 VDD1.n36 VDD1.n35 104.615
R239 VDD1.n133 VDD1.n132 104.615
R240 VDD1.n133 VDD1.n126 104.615
R241 VDD1.n140 VDD1.n126 104.615
R242 VDD1.n141 VDD1.n140 104.615
R243 VDD1.n141 VDD1.n122 104.615
R244 VDD1.n148 VDD1.n122 104.615
R245 VDD1.n149 VDD1.n148 104.615
R246 VDD1.n149 VDD1.n118 104.615
R247 VDD1.n156 VDD1.n118 104.615
R248 VDD1.n157 VDD1.n156 104.615
R249 VDD1.n157 VDD1.n114 104.615
R250 VDD1.n164 VDD1.n114 104.615
R251 VDD1.n165 VDD1.n164 104.615
R252 VDD1.n165 VDD1.n110 104.615
R253 VDD1.n173 VDD1.n110 104.615
R254 VDD1.n174 VDD1.n173 104.615
R255 VDD1.n175 VDD1.n174 104.615
R256 VDD1.n175 VDD1.n106 104.615
R257 VDD1.n182 VDD1.n106 104.615
R258 VDD1.n183 VDD1.n182 104.615
R259 VDD1.n183 VDD1.n102 104.615
R260 VDD1.n190 VDD1.n102 104.615
R261 VDD1.n191 VDD1.n190 104.615
R262 VDD1.n199 VDD1.n198 64.0209
R263 VDD1.n98 VDD1.n97 61.8458
R264 VDD1.n197 VDD1.n196 61.8456
R265 VDD1.n201 VDD1.n200 61.8456
R266 VDD1.n201 VDD1.n199 55.0677
R267 VDD1.n98 VDD1.n96 53.0019
R268 VDD1.n197 VDD1.n195 53.0019
R269 VDD1.n35 VDD1.t6 52.3082
R270 VDD1.n132 VDD1.t9 52.3082
R271 VDD1.n34 VDD1.n33 15.6677
R272 VDD1.n131 VDD1.n130 15.6677
R273 VDD1.n10 VDD1.n8 13.1884
R274 VDD1.n176 VDD1.n107 13.1884
R275 VDD1.n82 VDD1.n81 12.8005
R276 VDD1.n78 VDD1.n77 12.8005
R277 VDD1.n37 VDD1.n32 12.8005
R278 VDD1.n134 VDD1.n129 12.8005
R279 VDD1.n177 VDD1.n109 12.8005
R280 VDD1.n181 VDD1.n180 12.8005
R281 VDD1.n85 VDD1.n6 12.0247
R282 VDD1.n74 VDD1.n11 12.0247
R283 VDD1.n38 VDD1.n30 12.0247
R284 VDD1.n135 VDD1.n127 12.0247
R285 VDD1.n172 VDD1.n171 12.0247
R286 VDD1.n184 VDD1.n105 12.0247
R287 VDD1.n86 VDD1.n4 11.249
R288 VDD1.n73 VDD1.n14 11.249
R289 VDD1.n42 VDD1.n41 11.249
R290 VDD1.n139 VDD1.n138 11.249
R291 VDD1.n170 VDD1.n111 11.249
R292 VDD1.n185 VDD1.n103 11.249
R293 VDD1.n90 VDD1.n89 10.4732
R294 VDD1.n70 VDD1.n69 10.4732
R295 VDD1.n45 VDD1.n28 10.4732
R296 VDD1.n142 VDD1.n125 10.4732
R297 VDD1.n167 VDD1.n166 10.4732
R298 VDD1.n189 VDD1.n188 10.4732
R299 VDD1.n93 VDD1.n2 9.69747
R300 VDD1.n66 VDD1.n16 9.69747
R301 VDD1.n46 VDD1.n26 9.69747
R302 VDD1.n143 VDD1.n123 9.69747
R303 VDD1.n163 VDD1.n113 9.69747
R304 VDD1.n192 VDD1.n101 9.69747
R305 VDD1.n96 VDD1.n95 9.45567
R306 VDD1.n195 VDD1.n194 9.45567
R307 VDD1.n20 VDD1.n19 9.3005
R308 VDD1.n63 VDD1.n62 9.3005
R309 VDD1.n65 VDD1.n64 9.3005
R310 VDD1.n16 VDD1.n15 9.3005
R311 VDD1.n71 VDD1.n70 9.3005
R312 VDD1.n73 VDD1.n72 9.3005
R313 VDD1.n11 VDD1.n9 9.3005
R314 VDD1.n79 VDD1.n78 9.3005
R315 VDD1.n95 VDD1.n94 9.3005
R316 VDD1.n2 VDD1.n1 9.3005
R317 VDD1.n89 VDD1.n88 9.3005
R318 VDD1.n87 VDD1.n86 9.3005
R319 VDD1.n6 VDD1.n5 9.3005
R320 VDD1.n81 VDD1.n80 9.3005
R321 VDD1.n57 VDD1.n56 9.3005
R322 VDD1.n55 VDD1.n54 9.3005
R323 VDD1.n24 VDD1.n23 9.3005
R324 VDD1.n49 VDD1.n48 9.3005
R325 VDD1.n47 VDD1.n46 9.3005
R326 VDD1.n28 VDD1.n27 9.3005
R327 VDD1.n41 VDD1.n40 9.3005
R328 VDD1.n39 VDD1.n38 9.3005
R329 VDD1.n32 VDD1.n31 9.3005
R330 VDD1.n194 VDD1.n193 9.3005
R331 VDD1.n101 VDD1.n100 9.3005
R332 VDD1.n188 VDD1.n187 9.3005
R333 VDD1.n186 VDD1.n185 9.3005
R334 VDD1.n105 VDD1.n104 9.3005
R335 VDD1.n180 VDD1.n179 9.3005
R336 VDD1.n152 VDD1.n151 9.3005
R337 VDD1.n121 VDD1.n120 9.3005
R338 VDD1.n146 VDD1.n145 9.3005
R339 VDD1.n144 VDD1.n143 9.3005
R340 VDD1.n125 VDD1.n124 9.3005
R341 VDD1.n138 VDD1.n137 9.3005
R342 VDD1.n136 VDD1.n135 9.3005
R343 VDD1.n129 VDD1.n128 9.3005
R344 VDD1.n154 VDD1.n153 9.3005
R345 VDD1.n117 VDD1.n116 9.3005
R346 VDD1.n160 VDD1.n159 9.3005
R347 VDD1.n162 VDD1.n161 9.3005
R348 VDD1.n113 VDD1.n112 9.3005
R349 VDD1.n168 VDD1.n167 9.3005
R350 VDD1.n170 VDD1.n169 9.3005
R351 VDD1.n171 VDD1.n108 9.3005
R352 VDD1.n178 VDD1.n177 9.3005
R353 VDD1.n94 VDD1.n0 8.92171
R354 VDD1.n65 VDD1.n18 8.92171
R355 VDD1.n50 VDD1.n49 8.92171
R356 VDD1.n147 VDD1.n146 8.92171
R357 VDD1.n162 VDD1.n115 8.92171
R358 VDD1.n193 VDD1.n99 8.92171
R359 VDD1.n62 VDD1.n61 8.14595
R360 VDD1.n53 VDD1.n24 8.14595
R361 VDD1.n150 VDD1.n121 8.14595
R362 VDD1.n159 VDD1.n158 8.14595
R363 VDD1.n58 VDD1.n20 7.3702
R364 VDD1.n54 VDD1.n22 7.3702
R365 VDD1.n151 VDD1.n119 7.3702
R366 VDD1.n155 VDD1.n117 7.3702
R367 VDD1.n58 VDD1.n57 6.59444
R368 VDD1.n57 VDD1.n22 6.59444
R369 VDD1.n154 VDD1.n119 6.59444
R370 VDD1.n155 VDD1.n154 6.59444
R371 VDD1.n61 VDD1.n20 5.81868
R372 VDD1.n54 VDD1.n53 5.81868
R373 VDD1.n151 VDD1.n150 5.81868
R374 VDD1.n158 VDD1.n117 5.81868
R375 VDD1.n96 VDD1.n0 5.04292
R376 VDD1.n62 VDD1.n18 5.04292
R377 VDD1.n50 VDD1.n24 5.04292
R378 VDD1.n147 VDD1.n121 5.04292
R379 VDD1.n159 VDD1.n115 5.04292
R380 VDD1.n195 VDD1.n99 5.04292
R381 VDD1.n33 VDD1.n31 4.38563
R382 VDD1.n130 VDD1.n128 4.38563
R383 VDD1.n94 VDD1.n93 4.26717
R384 VDD1.n66 VDD1.n65 4.26717
R385 VDD1.n49 VDD1.n26 4.26717
R386 VDD1.n146 VDD1.n123 4.26717
R387 VDD1.n163 VDD1.n162 4.26717
R388 VDD1.n193 VDD1.n192 4.26717
R389 VDD1.n90 VDD1.n2 3.49141
R390 VDD1.n69 VDD1.n16 3.49141
R391 VDD1.n46 VDD1.n45 3.49141
R392 VDD1.n143 VDD1.n142 3.49141
R393 VDD1.n166 VDD1.n113 3.49141
R394 VDD1.n189 VDD1.n101 3.49141
R395 VDD1.n89 VDD1.n4 2.71565
R396 VDD1.n70 VDD1.n14 2.71565
R397 VDD1.n42 VDD1.n28 2.71565
R398 VDD1.n139 VDD1.n125 2.71565
R399 VDD1.n167 VDD1.n111 2.71565
R400 VDD1.n188 VDD1.n103 2.71565
R401 VDD1 VDD1.n201 2.17291
R402 VDD1.n86 VDD1.n85 1.93989
R403 VDD1.n74 VDD1.n73 1.93989
R404 VDD1.n41 VDD1.n30 1.93989
R405 VDD1.n138 VDD1.n127 1.93989
R406 VDD1.n172 VDD1.n170 1.93989
R407 VDD1.n185 VDD1.n184 1.93989
R408 VDD1.n82 VDD1.n6 1.16414
R409 VDD1.n77 VDD1.n11 1.16414
R410 VDD1.n38 VDD1.n37 1.16414
R411 VDD1.n135 VDD1.n134 1.16414
R412 VDD1.n171 VDD1.n109 1.16414
R413 VDD1.n181 VDD1.n105 1.16414
R414 VDD1.n200 VDD1.t0 1.12678
R415 VDD1.n200 VDD1.t4 1.12678
R416 VDD1.n97 VDD1.t1 1.12678
R417 VDD1.n97 VDD1.t7 1.12678
R418 VDD1.n198 VDD1.t5 1.12678
R419 VDD1.n198 VDD1.t3 1.12678
R420 VDD1.n196 VDD1.t8 1.12678
R421 VDD1.n196 VDD1.t2 1.12678
R422 VDD1 VDD1.n98 0.802224
R423 VDD1.n199 VDD1.n197 0.688688
R424 VDD1.n81 VDD1.n8 0.388379
R425 VDD1.n78 VDD1.n10 0.388379
R426 VDD1.n34 VDD1.n32 0.388379
R427 VDD1.n131 VDD1.n129 0.388379
R428 VDD1.n177 VDD1.n176 0.388379
R429 VDD1.n180 VDD1.n107 0.388379
R430 VDD1.n95 VDD1.n1 0.155672
R431 VDD1.n88 VDD1.n1 0.155672
R432 VDD1.n88 VDD1.n87 0.155672
R433 VDD1.n87 VDD1.n5 0.155672
R434 VDD1.n80 VDD1.n5 0.155672
R435 VDD1.n80 VDD1.n79 0.155672
R436 VDD1.n79 VDD1.n9 0.155672
R437 VDD1.n72 VDD1.n9 0.155672
R438 VDD1.n72 VDD1.n71 0.155672
R439 VDD1.n71 VDD1.n15 0.155672
R440 VDD1.n64 VDD1.n15 0.155672
R441 VDD1.n64 VDD1.n63 0.155672
R442 VDD1.n63 VDD1.n19 0.155672
R443 VDD1.n56 VDD1.n19 0.155672
R444 VDD1.n56 VDD1.n55 0.155672
R445 VDD1.n55 VDD1.n23 0.155672
R446 VDD1.n48 VDD1.n23 0.155672
R447 VDD1.n48 VDD1.n47 0.155672
R448 VDD1.n47 VDD1.n27 0.155672
R449 VDD1.n40 VDD1.n27 0.155672
R450 VDD1.n40 VDD1.n39 0.155672
R451 VDD1.n39 VDD1.n31 0.155672
R452 VDD1.n136 VDD1.n128 0.155672
R453 VDD1.n137 VDD1.n136 0.155672
R454 VDD1.n137 VDD1.n124 0.155672
R455 VDD1.n144 VDD1.n124 0.155672
R456 VDD1.n145 VDD1.n144 0.155672
R457 VDD1.n145 VDD1.n120 0.155672
R458 VDD1.n152 VDD1.n120 0.155672
R459 VDD1.n153 VDD1.n152 0.155672
R460 VDD1.n153 VDD1.n116 0.155672
R461 VDD1.n160 VDD1.n116 0.155672
R462 VDD1.n161 VDD1.n160 0.155672
R463 VDD1.n161 VDD1.n112 0.155672
R464 VDD1.n168 VDD1.n112 0.155672
R465 VDD1.n169 VDD1.n168 0.155672
R466 VDD1.n169 VDD1.n108 0.155672
R467 VDD1.n178 VDD1.n108 0.155672
R468 VDD1.n179 VDD1.n178 0.155672
R469 VDD1.n179 VDD1.n104 0.155672
R470 VDD1.n186 VDD1.n104 0.155672
R471 VDD1.n187 VDD1.n186 0.155672
R472 VDD1.n187 VDD1.n100 0.155672
R473 VDD1.n194 VDD1.n100 0.155672
R474 VTAIL.n400 VTAIL.n308 289.615
R475 VTAIL.n94 VTAIL.n2 289.615
R476 VTAIL.n302 VTAIL.n210 289.615
R477 VTAIL.n200 VTAIL.n108 289.615
R478 VTAIL.n341 VTAIL.n340 185
R479 VTAIL.n343 VTAIL.n342 185
R480 VTAIL.n336 VTAIL.n335 185
R481 VTAIL.n349 VTAIL.n348 185
R482 VTAIL.n351 VTAIL.n350 185
R483 VTAIL.n332 VTAIL.n331 185
R484 VTAIL.n357 VTAIL.n356 185
R485 VTAIL.n359 VTAIL.n358 185
R486 VTAIL.n328 VTAIL.n327 185
R487 VTAIL.n365 VTAIL.n364 185
R488 VTAIL.n367 VTAIL.n366 185
R489 VTAIL.n324 VTAIL.n323 185
R490 VTAIL.n373 VTAIL.n372 185
R491 VTAIL.n375 VTAIL.n374 185
R492 VTAIL.n320 VTAIL.n319 185
R493 VTAIL.n382 VTAIL.n381 185
R494 VTAIL.n383 VTAIL.n318 185
R495 VTAIL.n385 VTAIL.n384 185
R496 VTAIL.n316 VTAIL.n315 185
R497 VTAIL.n391 VTAIL.n390 185
R498 VTAIL.n393 VTAIL.n392 185
R499 VTAIL.n312 VTAIL.n311 185
R500 VTAIL.n399 VTAIL.n398 185
R501 VTAIL.n401 VTAIL.n400 185
R502 VTAIL.n35 VTAIL.n34 185
R503 VTAIL.n37 VTAIL.n36 185
R504 VTAIL.n30 VTAIL.n29 185
R505 VTAIL.n43 VTAIL.n42 185
R506 VTAIL.n45 VTAIL.n44 185
R507 VTAIL.n26 VTAIL.n25 185
R508 VTAIL.n51 VTAIL.n50 185
R509 VTAIL.n53 VTAIL.n52 185
R510 VTAIL.n22 VTAIL.n21 185
R511 VTAIL.n59 VTAIL.n58 185
R512 VTAIL.n61 VTAIL.n60 185
R513 VTAIL.n18 VTAIL.n17 185
R514 VTAIL.n67 VTAIL.n66 185
R515 VTAIL.n69 VTAIL.n68 185
R516 VTAIL.n14 VTAIL.n13 185
R517 VTAIL.n76 VTAIL.n75 185
R518 VTAIL.n77 VTAIL.n12 185
R519 VTAIL.n79 VTAIL.n78 185
R520 VTAIL.n10 VTAIL.n9 185
R521 VTAIL.n85 VTAIL.n84 185
R522 VTAIL.n87 VTAIL.n86 185
R523 VTAIL.n6 VTAIL.n5 185
R524 VTAIL.n93 VTAIL.n92 185
R525 VTAIL.n95 VTAIL.n94 185
R526 VTAIL.n303 VTAIL.n302 185
R527 VTAIL.n301 VTAIL.n300 185
R528 VTAIL.n214 VTAIL.n213 185
R529 VTAIL.n295 VTAIL.n294 185
R530 VTAIL.n293 VTAIL.n292 185
R531 VTAIL.n218 VTAIL.n217 185
R532 VTAIL.n222 VTAIL.n220 185
R533 VTAIL.n287 VTAIL.n286 185
R534 VTAIL.n285 VTAIL.n284 185
R535 VTAIL.n224 VTAIL.n223 185
R536 VTAIL.n279 VTAIL.n278 185
R537 VTAIL.n277 VTAIL.n276 185
R538 VTAIL.n228 VTAIL.n227 185
R539 VTAIL.n271 VTAIL.n270 185
R540 VTAIL.n269 VTAIL.n268 185
R541 VTAIL.n232 VTAIL.n231 185
R542 VTAIL.n263 VTAIL.n262 185
R543 VTAIL.n261 VTAIL.n260 185
R544 VTAIL.n236 VTAIL.n235 185
R545 VTAIL.n255 VTAIL.n254 185
R546 VTAIL.n253 VTAIL.n252 185
R547 VTAIL.n240 VTAIL.n239 185
R548 VTAIL.n247 VTAIL.n246 185
R549 VTAIL.n245 VTAIL.n244 185
R550 VTAIL.n201 VTAIL.n200 185
R551 VTAIL.n199 VTAIL.n198 185
R552 VTAIL.n112 VTAIL.n111 185
R553 VTAIL.n193 VTAIL.n192 185
R554 VTAIL.n191 VTAIL.n190 185
R555 VTAIL.n116 VTAIL.n115 185
R556 VTAIL.n120 VTAIL.n118 185
R557 VTAIL.n185 VTAIL.n184 185
R558 VTAIL.n183 VTAIL.n182 185
R559 VTAIL.n122 VTAIL.n121 185
R560 VTAIL.n177 VTAIL.n176 185
R561 VTAIL.n175 VTAIL.n174 185
R562 VTAIL.n126 VTAIL.n125 185
R563 VTAIL.n169 VTAIL.n168 185
R564 VTAIL.n167 VTAIL.n166 185
R565 VTAIL.n130 VTAIL.n129 185
R566 VTAIL.n161 VTAIL.n160 185
R567 VTAIL.n159 VTAIL.n158 185
R568 VTAIL.n134 VTAIL.n133 185
R569 VTAIL.n153 VTAIL.n152 185
R570 VTAIL.n151 VTAIL.n150 185
R571 VTAIL.n138 VTAIL.n137 185
R572 VTAIL.n145 VTAIL.n144 185
R573 VTAIL.n143 VTAIL.n142 185
R574 VTAIL.n339 VTAIL.t2 147.659
R575 VTAIL.n33 VTAIL.t17 147.659
R576 VTAIL.n243 VTAIL.t10 147.659
R577 VTAIL.n141 VTAIL.t1 147.659
R578 VTAIL.n342 VTAIL.n341 104.615
R579 VTAIL.n342 VTAIL.n335 104.615
R580 VTAIL.n349 VTAIL.n335 104.615
R581 VTAIL.n350 VTAIL.n349 104.615
R582 VTAIL.n350 VTAIL.n331 104.615
R583 VTAIL.n357 VTAIL.n331 104.615
R584 VTAIL.n358 VTAIL.n357 104.615
R585 VTAIL.n358 VTAIL.n327 104.615
R586 VTAIL.n365 VTAIL.n327 104.615
R587 VTAIL.n366 VTAIL.n365 104.615
R588 VTAIL.n366 VTAIL.n323 104.615
R589 VTAIL.n373 VTAIL.n323 104.615
R590 VTAIL.n374 VTAIL.n373 104.615
R591 VTAIL.n374 VTAIL.n319 104.615
R592 VTAIL.n382 VTAIL.n319 104.615
R593 VTAIL.n383 VTAIL.n382 104.615
R594 VTAIL.n384 VTAIL.n383 104.615
R595 VTAIL.n384 VTAIL.n315 104.615
R596 VTAIL.n391 VTAIL.n315 104.615
R597 VTAIL.n392 VTAIL.n391 104.615
R598 VTAIL.n392 VTAIL.n311 104.615
R599 VTAIL.n399 VTAIL.n311 104.615
R600 VTAIL.n400 VTAIL.n399 104.615
R601 VTAIL.n36 VTAIL.n35 104.615
R602 VTAIL.n36 VTAIL.n29 104.615
R603 VTAIL.n43 VTAIL.n29 104.615
R604 VTAIL.n44 VTAIL.n43 104.615
R605 VTAIL.n44 VTAIL.n25 104.615
R606 VTAIL.n51 VTAIL.n25 104.615
R607 VTAIL.n52 VTAIL.n51 104.615
R608 VTAIL.n52 VTAIL.n21 104.615
R609 VTAIL.n59 VTAIL.n21 104.615
R610 VTAIL.n60 VTAIL.n59 104.615
R611 VTAIL.n60 VTAIL.n17 104.615
R612 VTAIL.n67 VTAIL.n17 104.615
R613 VTAIL.n68 VTAIL.n67 104.615
R614 VTAIL.n68 VTAIL.n13 104.615
R615 VTAIL.n76 VTAIL.n13 104.615
R616 VTAIL.n77 VTAIL.n76 104.615
R617 VTAIL.n78 VTAIL.n77 104.615
R618 VTAIL.n78 VTAIL.n9 104.615
R619 VTAIL.n85 VTAIL.n9 104.615
R620 VTAIL.n86 VTAIL.n85 104.615
R621 VTAIL.n86 VTAIL.n5 104.615
R622 VTAIL.n93 VTAIL.n5 104.615
R623 VTAIL.n94 VTAIL.n93 104.615
R624 VTAIL.n302 VTAIL.n301 104.615
R625 VTAIL.n301 VTAIL.n213 104.615
R626 VTAIL.n294 VTAIL.n213 104.615
R627 VTAIL.n294 VTAIL.n293 104.615
R628 VTAIL.n293 VTAIL.n217 104.615
R629 VTAIL.n222 VTAIL.n217 104.615
R630 VTAIL.n286 VTAIL.n222 104.615
R631 VTAIL.n286 VTAIL.n285 104.615
R632 VTAIL.n285 VTAIL.n223 104.615
R633 VTAIL.n278 VTAIL.n223 104.615
R634 VTAIL.n278 VTAIL.n277 104.615
R635 VTAIL.n277 VTAIL.n227 104.615
R636 VTAIL.n270 VTAIL.n227 104.615
R637 VTAIL.n270 VTAIL.n269 104.615
R638 VTAIL.n269 VTAIL.n231 104.615
R639 VTAIL.n262 VTAIL.n231 104.615
R640 VTAIL.n262 VTAIL.n261 104.615
R641 VTAIL.n261 VTAIL.n235 104.615
R642 VTAIL.n254 VTAIL.n235 104.615
R643 VTAIL.n254 VTAIL.n253 104.615
R644 VTAIL.n253 VTAIL.n239 104.615
R645 VTAIL.n246 VTAIL.n239 104.615
R646 VTAIL.n246 VTAIL.n245 104.615
R647 VTAIL.n200 VTAIL.n199 104.615
R648 VTAIL.n199 VTAIL.n111 104.615
R649 VTAIL.n192 VTAIL.n111 104.615
R650 VTAIL.n192 VTAIL.n191 104.615
R651 VTAIL.n191 VTAIL.n115 104.615
R652 VTAIL.n120 VTAIL.n115 104.615
R653 VTAIL.n184 VTAIL.n120 104.615
R654 VTAIL.n184 VTAIL.n183 104.615
R655 VTAIL.n183 VTAIL.n121 104.615
R656 VTAIL.n176 VTAIL.n121 104.615
R657 VTAIL.n176 VTAIL.n175 104.615
R658 VTAIL.n175 VTAIL.n125 104.615
R659 VTAIL.n168 VTAIL.n125 104.615
R660 VTAIL.n168 VTAIL.n167 104.615
R661 VTAIL.n167 VTAIL.n129 104.615
R662 VTAIL.n160 VTAIL.n129 104.615
R663 VTAIL.n160 VTAIL.n159 104.615
R664 VTAIL.n159 VTAIL.n133 104.615
R665 VTAIL.n152 VTAIL.n133 104.615
R666 VTAIL.n152 VTAIL.n151 104.615
R667 VTAIL.n151 VTAIL.n137 104.615
R668 VTAIL.n144 VTAIL.n137 104.615
R669 VTAIL.n144 VTAIL.n143 104.615
R670 VTAIL.n341 VTAIL.t2 52.3082
R671 VTAIL.n35 VTAIL.t17 52.3082
R672 VTAIL.n245 VTAIL.t10 52.3082
R673 VTAIL.n143 VTAIL.t1 52.3082
R674 VTAIL.n209 VTAIL.n208 45.167
R675 VTAIL.n207 VTAIL.n206 45.167
R676 VTAIL.n107 VTAIL.n106 45.167
R677 VTAIL.n105 VTAIL.n104 45.167
R678 VTAIL.n407 VTAIL.n406 45.1668
R679 VTAIL.n1 VTAIL.n0 45.1668
R680 VTAIL.n101 VTAIL.n100 45.1668
R681 VTAIL.n103 VTAIL.n102 45.1668
R682 VTAIL.n105 VTAIL.n103 33.4703
R683 VTAIL.n405 VTAIL.n404 33.349
R684 VTAIL.n99 VTAIL.n98 33.349
R685 VTAIL.n307 VTAIL.n306 33.349
R686 VTAIL.n205 VTAIL.n204 33.349
R687 VTAIL.n405 VTAIL.n307 30.4962
R688 VTAIL.n340 VTAIL.n339 15.6677
R689 VTAIL.n34 VTAIL.n33 15.6677
R690 VTAIL.n244 VTAIL.n243 15.6677
R691 VTAIL.n142 VTAIL.n141 15.6677
R692 VTAIL.n385 VTAIL.n316 13.1884
R693 VTAIL.n79 VTAIL.n10 13.1884
R694 VTAIL.n220 VTAIL.n218 13.1884
R695 VTAIL.n118 VTAIL.n116 13.1884
R696 VTAIL.n343 VTAIL.n338 12.8005
R697 VTAIL.n386 VTAIL.n318 12.8005
R698 VTAIL.n390 VTAIL.n389 12.8005
R699 VTAIL.n37 VTAIL.n32 12.8005
R700 VTAIL.n80 VTAIL.n12 12.8005
R701 VTAIL.n84 VTAIL.n83 12.8005
R702 VTAIL.n292 VTAIL.n291 12.8005
R703 VTAIL.n288 VTAIL.n287 12.8005
R704 VTAIL.n247 VTAIL.n242 12.8005
R705 VTAIL.n190 VTAIL.n189 12.8005
R706 VTAIL.n186 VTAIL.n185 12.8005
R707 VTAIL.n145 VTAIL.n140 12.8005
R708 VTAIL.n344 VTAIL.n336 12.0247
R709 VTAIL.n381 VTAIL.n380 12.0247
R710 VTAIL.n393 VTAIL.n314 12.0247
R711 VTAIL.n38 VTAIL.n30 12.0247
R712 VTAIL.n75 VTAIL.n74 12.0247
R713 VTAIL.n87 VTAIL.n8 12.0247
R714 VTAIL.n295 VTAIL.n216 12.0247
R715 VTAIL.n284 VTAIL.n221 12.0247
R716 VTAIL.n248 VTAIL.n240 12.0247
R717 VTAIL.n193 VTAIL.n114 12.0247
R718 VTAIL.n182 VTAIL.n119 12.0247
R719 VTAIL.n146 VTAIL.n138 12.0247
R720 VTAIL.n348 VTAIL.n347 11.249
R721 VTAIL.n379 VTAIL.n320 11.249
R722 VTAIL.n394 VTAIL.n312 11.249
R723 VTAIL.n42 VTAIL.n41 11.249
R724 VTAIL.n73 VTAIL.n14 11.249
R725 VTAIL.n88 VTAIL.n6 11.249
R726 VTAIL.n296 VTAIL.n214 11.249
R727 VTAIL.n283 VTAIL.n224 11.249
R728 VTAIL.n252 VTAIL.n251 11.249
R729 VTAIL.n194 VTAIL.n112 11.249
R730 VTAIL.n181 VTAIL.n122 11.249
R731 VTAIL.n150 VTAIL.n149 11.249
R732 VTAIL.n351 VTAIL.n334 10.4732
R733 VTAIL.n376 VTAIL.n375 10.4732
R734 VTAIL.n398 VTAIL.n397 10.4732
R735 VTAIL.n45 VTAIL.n28 10.4732
R736 VTAIL.n70 VTAIL.n69 10.4732
R737 VTAIL.n92 VTAIL.n91 10.4732
R738 VTAIL.n300 VTAIL.n299 10.4732
R739 VTAIL.n280 VTAIL.n279 10.4732
R740 VTAIL.n255 VTAIL.n238 10.4732
R741 VTAIL.n198 VTAIL.n197 10.4732
R742 VTAIL.n178 VTAIL.n177 10.4732
R743 VTAIL.n153 VTAIL.n136 10.4732
R744 VTAIL.n352 VTAIL.n332 9.69747
R745 VTAIL.n372 VTAIL.n322 9.69747
R746 VTAIL.n401 VTAIL.n310 9.69747
R747 VTAIL.n46 VTAIL.n26 9.69747
R748 VTAIL.n66 VTAIL.n16 9.69747
R749 VTAIL.n95 VTAIL.n4 9.69747
R750 VTAIL.n303 VTAIL.n212 9.69747
R751 VTAIL.n276 VTAIL.n226 9.69747
R752 VTAIL.n256 VTAIL.n236 9.69747
R753 VTAIL.n201 VTAIL.n110 9.69747
R754 VTAIL.n174 VTAIL.n124 9.69747
R755 VTAIL.n154 VTAIL.n134 9.69747
R756 VTAIL.n404 VTAIL.n403 9.45567
R757 VTAIL.n98 VTAIL.n97 9.45567
R758 VTAIL.n306 VTAIL.n305 9.45567
R759 VTAIL.n204 VTAIL.n203 9.45567
R760 VTAIL.n403 VTAIL.n402 9.3005
R761 VTAIL.n310 VTAIL.n309 9.3005
R762 VTAIL.n397 VTAIL.n396 9.3005
R763 VTAIL.n395 VTAIL.n394 9.3005
R764 VTAIL.n314 VTAIL.n313 9.3005
R765 VTAIL.n389 VTAIL.n388 9.3005
R766 VTAIL.n361 VTAIL.n360 9.3005
R767 VTAIL.n330 VTAIL.n329 9.3005
R768 VTAIL.n355 VTAIL.n354 9.3005
R769 VTAIL.n353 VTAIL.n352 9.3005
R770 VTAIL.n334 VTAIL.n333 9.3005
R771 VTAIL.n347 VTAIL.n346 9.3005
R772 VTAIL.n345 VTAIL.n344 9.3005
R773 VTAIL.n338 VTAIL.n337 9.3005
R774 VTAIL.n363 VTAIL.n362 9.3005
R775 VTAIL.n326 VTAIL.n325 9.3005
R776 VTAIL.n369 VTAIL.n368 9.3005
R777 VTAIL.n371 VTAIL.n370 9.3005
R778 VTAIL.n322 VTAIL.n321 9.3005
R779 VTAIL.n377 VTAIL.n376 9.3005
R780 VTAIL.n379 VTAIL.n378 9.3005
R781 VTAIL.n380 VTAIL.n317 9.3005
R782 VTAIL.n387 VTAIL.n386 9.3005
R783 VTAIL.n97 VTAIL.n96 9.3005
R784 VTAIL.n4 VTAIL.n3 9.3005
R785 VTAIL.n91 VTAIL.n90 9.3005
R786 VTAIL.n89 VTAIL.n88 9.3005
R787 VTAIL.n8 VTAIL.n7 9.3005
R788 VTAIL.n83 VTAIL.n82 9.3005
R789 VTAIL.n55 VTAIL.n54 9.3005
R790 VTAIL.n24 VTAIL.n23 9.3005
R791 VTAIL.n49 VTAIL.n48 9.3005
R792 VTAIL.n47 VTAIL.n46 9.3005
R793 VTAIL.n28 VTAIL.n27 9.3005
R794 VTAIL.n41 VTAIL.n40 9.3005
R795 VTAIL.n39 VTAIL.n38 9.3005
R796 VTAIL.n32 VTAIL.n31 9.3005
R797 VTAIL.n57 VTAIL.n56 9.3005
R798 VTAIL.n20 VTAIL.n19 9.3005
R799 VTAIL.n63 VTAIL.n62 9.3005
R800 VTAIL.n65 VTAIL.n64 9.3005
R801 VTAIL.n16 VTAIL.n15 9.3005
R802 VTAIL.n71 VTAIL.n70 9.3005
R803 VTAIL.n73 VTAIL.n72 9.3005
R804 VTAIL.n74 VTAIL.n11 9.3005
R805 VTAIL.n81 VTAIL.n80 9.3005
R806 VTAIL.n230 VTAIL.n229 9.3005
R807 VTAIL.n273 VTAIL.n272 9.3005
R808 VTAIL.n275 VTAIL.n274 9.3005
R809 VTAIL.n226 VTAIL.n225 9.3005
R810 VTAIL.n281 VTAIL.n280 9.3005
R811 VTAIL.n283 VTAIL.n282 9.3005
R812 VTAIL.n221 VTAIL.n219 9.3005
R813 VTAIL.n289 VTAIL.n288 9.3005
R814 VTAIL.n305 VTAIL.n304 9.3005
R815 VTAIL.n212 VTAIL.n211 9.3005
R816 VTAIL.n299 VTAIL.n298 9.3005
R817 VTAIL.n297 VTAIL.n296 9.3005
R818 VTAIL.n216 VTAIL.n215 9.3005
R819 VTAIL.n291 VTAIL.n290 9.3005
R820 VTAIL.n267 VTAIL.n266 9.3005
R821 VTAIL.n265 VTAIL.n264 9.3005
R822 VTAIL.n234 VTAIL.n233 9.3005
R823 VTAIL.n259 VTAIL.n258 9.3005
R824 VTAIL.n257 VTAIL.n256 9.3005
R825 VTAIL.n238 VTAIL.n237 9.3005
R826 VTAIL.n251 VTAIL.n250 9.3005
R827 VTAIL.n249 VTAIL.n248 9.3005
R828 VTAIL.n242 VTAIL.n241 9.3005
R829 VTAIL.n128 VTAIL.n127 9.3005
R830 VTAIL.n171 VTAIL.n170 9.3005
R831 VTAIL.n173 VTAIL.n172 9.3005
R832 VTAIL.n124 VTAIL.n123 9.3005
R833 VTAIL.n179 VTAIL.n178 9.3005
R834 VTAIL.n181 VTAIL.n180 9.3005
R835 VTAIL.n119 VTAIL.n117 9.3005
R836 VTAIL.n187 VTAIL.n186 9.3005
R837 VTAIL.n203 VTAIL.n202 9.3005
R838 VTAIL.n110 VTAIL.n109 9.3005
R839 VTAIL.n197 VTAIL.n196 9.3005
R840 VTAIL.n195 VTAIL.n194 9.3005
R841 VTAIL.n114 VTAIL.n113 9.3005
R842 VTAIL.n189 VTAIL.n188 9.3005
R843 VTAIL.n165 VTAIL.n164 9.3005
R844 VTAIL.n163 VTAIL.n162 9.3005
R845 VTAIL.n132 VTAIL.n131 9.3005
R846 VTAIL.n157 VTAIL.n156 9.3005
R847 VTAIL.n155 VTAIL.n154 9.3005
R848 VTAIL.n136 VTAIL.n135 9.3005
R849 VTAIL.n149 VTAIL.n148 9.3005
R850 VTAIL.n147 VTAIL.n146 9.3005
R851 VTAIL.n140 VTAIL.n139 9.3005
R852 VTAIL.n356 VTAIL.n355 8.92171
R853 VTAIL.n371 VTAIL.n324 8.92171
R854 VTAIL.n402 VTAIL.n308 8.92171
R855 VTAIL.n50 VTAIL.n49 8.92171
R856 VTAIL.n65 VTAIL.n18 8.92171
R857 VTAIL.n96 VTAIL.n2 8.92171
R858 VTAIL.n304 VTAIL.n210 8.92171
R859 VTAIL.n275 VTAIL.n228 8.92171
R860 VTAIL.n260 VTAIL.n259 8.92171
R861 VTAIL.n202 VTAIL.n108 8.92171
R862 VTAIL.n173 VTAIL.n126 8.92171
R863 VTAIL.n158 VTAIL.n157 8.92171
R864 VTAIL.n359 VTAIL.n330 8.14595
R865 VTAIL.n368 VTAIL.n367 8.14595
R866 VTAIL.n53 VTAIL.n24 8.14595
R867 VTAIL.n62 VTAIL.n61 8.14595
R868 VTAIL.n272 VTAIL.n271 8.14595
R869 VTAIL.n263 VTAIL.n234 8.14595
R870 VTAIL.n170 VTAIL.n169 8.14595
R871 VTAIL.n161 VTAIL.n132 8.14595
R872 VTAIL.n360 VTAIL.n328 7.3702
R873 VTAIL.n364 VTAIL.n326 7.3702
R874 VTAIL.n54 VTAIL.n22 7.3702
R875 VTAIL.n58 VTAIL.n20 7.3702
R876 VTAIL.n268 VTAIL.n230 7.3702
R877 VTAIL.n264 VTAIL.n232 7.3702
R878 VTAIL.n166 VTAIL.n128 7.3702
R879 VTAIL.n162 VTAIL.n130 7.3702
R880 VTAIL.n363 VTAIL.n328 6.59444
R881 VTAIL.n364 VTAIL.n363 6.59444
R882 VTAIL.n57 VTAIL.n22 6.59444
R883 VTAIL.n58 VTAIL.n57 6.59444
R884 VTAIL.n268 VTAIL.n267 6.59444
R885 VTAIL.n267 VTAIL.n232 6.59444
R886 VTAIL.n166 VTAIL.n165 6.59444
R887 VTAIL.n165 VTAIL.n130 6.59444
R888 VTAIL.n360 VTAIL.n359 5.81868
R889 VTAIL.n367 VTAIL.n326 5.81868
R890 VTAIL.n54 VTAIL.n53 5.81868
R891 VTAIL.n61 VTAIL.n20 5.81868
R892 VTAIL.n271 VTAIL.n230 5.81868
R893 VTAIL.n264 VTAIL.n263 5.81868
R894 VTAIL.n169 VTAIL.n128 5.81868
R895 VTAIL.n162 VTAIL.n161 5.81868
R896 VTAIL.n356 VTAIL.n330 5.04292
R897 VTAIL.n368 VTAIL.n324 5.04292
R898 VTAIL.n404 VTAIL.n308 5.04292
R899 VTAIL.n50 VTAIL.n24 5.04292
R900 VTAIL.n62 VTAIL.n18 5.04292
R901 VTAIL.n98 VTAIL.n2 5.04292
R902 VTAIL.n306 VTAIL.n210 5.04292
R903 VTAIL.n272 VTAIL.n228 5.04292
R904 VTAIL.n260 VTAIL.n234 5.04292
R905 VTAIL.n204 VTAIL.n108 5.04292
R906 VTAIL.n170 VTAIL.n126 5.04292
R907 VTAIL.n158 VTAIL.n132 5.04292
R908 VTAIL.n339 VTAIL.n337 4.38563
R909 VTAIL.n33 VTAIL.n31 4.38563
R910 VTAIL.n243 VTAIL.n241 4.38563
R911 VTAIL.n141 VTAIL.n139 4.38563
R912 VTAIL.n355 VTAIL.n332 4.26717
R913 VTAIL.n372 VTAIL.n371 4.26717
R914 VTAIL.n402 VTAIL.n401 4.26717
R915 VTAIL.n49 VTAIL.n26 4.26717
R916 VTAIL.n66 VTAIL.n65 4.26717
R917 VTAIL.n96 VTAIL.n95 4.26717
R918 VTAIL.n304 VTAIL.n303 4.26717
R919 VTAIL.n276 VTAIL.n275 4.26717
R920 VTAIL.n259 VTAIL.n236 4.26717
R921 VTAIL.n202 VTAIL.n201 4.26717
R922 VTAIL.n174 VTAIL.n173 4.26717
R923 VTAIL.n157 VTAIL.n134 4.26717
R924 VTAIL.n352 VTAIL.n351 3.49141
R925 VTAIL.n375 VTAIL.n322 3.49141
R926 VTAIL.n398 VTAIL.n310 3.49141
R927 VTAIL.n46 VTAIL.n45 3.49141
R928 VTAIL.n69 VTAIL.n16 3.49141
R929 VTAIL.n92 VTAIL.n4 3.49141
R930 VTAIL.n300 VTAIL.n212 3.49141
R931 VTAIL.n279 VTAIL.n226 3.49141
R932 VTAIL.n256 VTAIL.n255 3.49141
R933 VTAIL.n198 VTAIL.n110 3.49141
R934 VTAIL.n177 VTAIL.n124 3.49141
R935 VTAIL.n154 VTAIL.n153 3.49141
R936 VTAIL.n107 VTAIL.n105 2.97464
R937 VTAIL.n205 VTAIL.n107 2.97464
R938 VTAIL.n209 VTAIL.n207 2.97464
R939 VTAIL.n307 VTAIL.n209 2.97464
R940 VTAIL.n103 VTAIL.n101 2.97464
R941 VTAIL.n101 VTAIL.n99 2.97464
R942 VTAIL.n407 VTAIL.n405 2.97464
R943 VTAIL.n348 VTAIL.n334 2.71565
R944 VTAIL.n376 VTAIL.n320 2.71565
R945 VTAIL.n397 VTAIL.n312 2.71565
R946 VTAIL.n42 VTAIL.n28 2.71565
R947 VTAIL.n70 VTAIL.n14 2.71565
R948 VTAIL.n91 VTAIL.n6 2.71565
R949 VTAIL.n299 VTAIL.n214 2.71565
R950 VTAIL.n280 VTAIL.n224 2.71565
R951 VTAIL.n252 VTAIL.n238 2.71565
R952 VTAIL.n197 VTAIL.n112 2.71565
R953 VTAIL.n178 VTAIL.n122 2.71565
R954 VTAIL.n150 VTAIL.n136 2.71565
R955 VTAIL VTAIL.n1 2.28929
R956 VTAIL.n207 VTAIL.n205 1.9574
R957 VTAIL.n99 VTAIL.n1 1.9574
R958 VTAIL.n347 VTAIL.n336 1.93989
R959 VTAIL.n381 VTAIL.n379 1.93989
R960 VTAIL.n394 VTAIL.n393 1.93989
R961 VTAIL.n41 VTAIL.n30 1.93989
R962 VTAIL.n75 VTAIL.n73 1.93989
R963 VTAIL.n88 VTAIL.n87 1.93989
R964 VTAIL.n296 VTAIL.n295 1.93989
R965 VTAIL.n284 VTAIL.n283 1.93989
R966 VTAIL.n251 VTAIL.n240 1.93989
R967 VTAIL.n194 VTAIL.n193 1.93989
R968 VTAIL.n182 VTAIL.n181 1.93989
R969 VTAIL.n149 VTAIL.n138 1.93989
R970 VTAIL.n344 VTAIL.n343 1.16414
R971 VTAIL.n380 VTAIL.n318 1.16414
R972 VTAIL.n390 VTAIL.n314 1.16414
R973 VTAIL.n38 VTAIL.n37 1.16414
R974 VTAIL.n74 VTAIL.n12 1.16414
R975 VTAIL.n84 VTAIL.n8 1.16414
R976 VTAIL.n292 VTAIL.n216 1.16414
R977 VTAIL.n287 VTAIL.n221 1.16414
R978 VTAIL.n248 VTAIL.n247 1.16414
R979 VTAIL.n190 VTAIL.n114 1.16414
R980 VTAIL.n185 VTAIL.n119 1.16414
R981 VTAIL.n146 VTAIL.n145 1.16414
R982 VTAIL.n406 VTAIL.t3 1.12678
R983 VTAIL.n406 VTAIL.t4 1.12678
R984 VTAIL.n0 VTAIL.t5 1.12678
R985 VTAIL.n0 VTAIL.t6 1.12678
R986 VTAIL.n100 VTAIL.t16 1.12678
R987 VTAIL.n100 VTAIL.t11 1.12678
R988 VTAIL.n102 VTAIL.t15 1.12678
R989 VTAIL.n102 VTAIL.t14 1.12678
R990 VTAIL.n208 VTAIL.t13 1.12678
R991 VTAIL.n208 VTAIL.t18 1.12678
R992 VTAIL.n206 VTAIL.t12 1.12678
R993 VTAIL.n206 VTAIL.t19 1.12678
R994 VTAIL.n106 VTAIL.t0 1.12678
R995 VTAIL.n106 VTAIL.t9 1.12678
R996 VTAIL.n104 VTAIL.t8 1.12678
R997 VTAIL.n104 VTAIL.t7 1.12678
R998 VTAIL VTAIL.n407 0.685845
R999 VTAIL.n340 VTAIL.n338 0.388379
R1000 VTAIL.n386 VTAIL.n385 0.388379
R1001 VTAIL.n389 VTAIL.n316 0.388379
R1002 VTAIL.n34 VTAIL.n32 0.388379
R1003 VTAIL.n80 VTAIL.n79 0.388379
R1004 VTAIL.n83 VTAIL.n10 0.388379
R1005 VTAIL.n291 VTAIL.n218 0.388379
R1006 VTAIL.n288 VTAIL.n220 0.388379
R1007 VTAIL.n244 VTAIL.n242 0.388379
R1008 VTAIL.n189 VTAIL.n116 0.388379
R1009 VTAIL.n186 VTAIL.n118 0.388379
R1010 VTAIL.n142 VTAIL.n140 0.388379
R1011 VTAIL.n345 VTAIL.n337 0.155672
R1012 VTAIL.n346 VTAIL.n345 0.155672
R1013 VTAIL.n346 VTAIL.n333 0.155672
R1014 VTAIL.n353 VTAIL.n333 0.155672
R1015 VTAIL.n354 VTAIL.n353 0.155672
R1016 VTAIL.n354 VTAIL.n329 0.155672
R1017 VTAIL.n361 VTAIL.n329 0.155672
R1018 VTAIL.n362 VTAIL.n361 0.155672
R1019 VTAIL.n362 VTAIL.n325 0.155672
R1020 VTAIL.n369 VTAIL.n325 0.155672
R1021 VTAIL.n370 VTAIL.n369 0.155672
R1022 VTAIL.n370 VTAIL.n321 0.155672
R1023 VTAIL.n377 VTAIL.n321 0.155672
R1024 VTAIL.n378 VTAIL.n377 0.155672
R1025 VTAIL.n378 VTAIL.n317 0.155672
R1026 VTAIL.n387 VTAIL.n317 0.155672
R1027 VTAIL.n388 VTAIL.n387 0.155672
R1028 VTAIL.n388 VTAIL.n313 0.155672
R1029 VTAIL.n395 VTAIL.n313 0.155672
R1030 VTAIL.n396 VTAIL.n395 0.155672
R1031 VTAIL.n396 VTAIL.n309 0.155672
R1032 VTAIL.n403 VTAIL.n309 0.155672
R1033 VTAIL.n39 VTAIL.n31 0.155672
R1034 VTAIL.n40 VTAIL.n39 0.155672
R1035 VTAIL.n40 VTAIL.n27 0.155672
R1036 VTAIL.n47 VTAIL.n27 0.155672
R1037 VTAIL.n48 VTAIL.n47 0.155672
R1038 VTAIL.n48 VTAIL.n23 0.155672
R1039 VTAIL.n55 VTAIL.n23 0.155672
R1040 VTAIL.n56 VTAIL.n55 0.155672
R1041 VTAIL.n56 VTAIL.n19 0.155672
R1042 VTAIL.n63 VTAIL.n19 0.155672
R1043 VTAIL.n64 VTAIL.n63 0.155672
R1044 VTAIL.n64 VTAIL.n15 0.155672
R1045 VTAIL.n71 VTAIL.n15 0.155672
R1046 VTAIL.n72 VTAIL.n71 0.155672
R1047 VTAIL.n72 VTAIL.n11 0.155672
R1048 VTAIL.n81 VTAIL.n11 0.155672
R1049 VTAIL.n82 VTAIL.n81 0.155672
R1050 VTAIL.n82 VTAIL.n7 0.155672
R1051 VTAIL.n89 VTAIL.n7 0.155672
R1052 VTAIL.n90 VTAIL.n89 0.155672
R1053 VTAIL.n90 VTAIL.n3 0.155672
R1054 VTAIL.n97 VTAIL.n3 0.155672
R1055 VTAIL.n305 VTAIL.n211 0.155672
R1056 VTAIL.n298 VTAIL.n211 0.155672
R1057 VTAIL.n298 VTAIL.n297 0.155672
R1058 VTAIL.n297 VTAIL.n215 0.155672
R1059 VTAIL.n290 VTAIL.n215 0.155672
R1060 VTAIL.n290 VTAIL.n289 0.155672
R1061 VTAIL.n289 VTAIL.n219 0.155672
R1062 VTAIL.n282 VTAIL.n219 0.155672
R1063 VTAIL.n282 VTAIL.n281 0.155672
R1064 VTAIL.n281 VTAIL.n225 0.155672
R1065 VTAIL.n274 VTAIL.n225 0.155672
R1066 VTAIL.n274 VTAIL.n273 0.155672
R1067 VTAIL.n273 VTAIL.n229 0.155672
R1068 VTAIL.n266 VTAIL.n229 0.155672
R1069 VTAIL.n266 VTAIL.n265 0.155672
R1070 VTAIL.n265 VTAIL.n233 0.155672
R1071 VTAIL.n258 VTAIL.n233 0.155672
R1072 VTAIL.n258 VTAIL.n257 0.155672
R1073 VTAIL.n257 VTAIL.n237 0.155672
R1074 VTAIL.n250 VTAIL.n237 0.155672
R1075 VTAIL.n250 VTAIL.n249 0.155672
R1076 VTAIL.n249 VTAIL.n241 0.155672
R1077 VTAIL.n203 VTAIL.n109 0.155672
R1078 VTAIL.n196 VTAIL.n109 0.155672
R1079 VTAIL.n196 VTAIL.n195 0.155672
R1080 VTAIL.n195 VTAIL.n113 0.155672
R1081 VTAIL.n188 VTAIL.n113 0.155672
R1082 VTAIL.n188 VTAIL.n187 0.155672
R1083 VTAIL.n187 VTAIL.n117 0.155672
R1084 VTAIL.n180 VTAIL.n117 0.155672
R1085 VTAIL.n180 VTAIL.n179 0.155672
R1086 VTAIL.n179 VTAIL.n123 0.155672
R1087 VTAIL.n172 VTAIL.n123 0.155672
R1088 VTAIL.n172 VTAIL.n171 0.155672
R1089 VTAIL.n171 VTAIL.n127 0.155672
R1090 VTAIL.n164 VTAIL.n127 0.155672
R1091 VTAIL.n164 VTAIL.n163 0.155672
R1092 VTAIL.n163 VTAIL.n131 0.155672
R1093 VTAIL.n156 VTAIL.n131 0.155672
R1094 VTAIL.n156 VTAIL.n155 0.155672
R1095 VTAIL.n155 VTAIL.n135 0.155672
R1096 VTAIL.n148 VTAIL.n135 0.155672
R1097 VTAIL.n148 VTAIL.n147 0.155672
R1098 VTAIL.n147 VTAIL.n139 0.155672
R1099 B.n1195 B.n1194 585
R1100 B.n443 B.n188 585
R1101 B.n442 B.n441 585
R1102 B.n440 B.n439 585
R1103 B.n438 B.n437 585
R1104 B.n436 B.n435 585
R1105 B.n434 B.n433 585
R1106 B.n432 B.n431 585
R1107 B.n430 B.n429 585
R1108 B.n428 B.n427 585
R1109 B.n426 B.n425 585
R1110 B.n424 B.n423 585
R1111 B.n422 B.n421 585
R1112 B.n420 B.n419 585
R1113 B.n418 B.n417 585
R1114 B.n416 B.n415 585
R1115 B.n414 B.n413 585
R1116 B.n412 B.n411 585
R1117 B.n410 B.n409 585
R1118 B.n408 B.n407 585
R1119 B.n406 B.n405 585
R1120 B.n404 B.n403 585
R1121 B.n402 B.n401 585
R1122 B.n400 B.n399 585
R1123 B.n398 B.n397 585
R1124 B.n396 B.n395 585
R1125 B.n394 B.n393 585
R1126 B.n392 B.n391 585
R1127 B.n390 B.n389 585
R1128 B.n388 B.n387 585
R1129 B.n386 B.n385 585
R1130 B.n384 B.n383 585
R1131 B.n382 B.n381 585
R1132 B.n380 B.n379 585
R1133 B.n378 B.n377 585
R1134 B.n376 B.n375 585
R1135 B.n374 B.n373 585
R1136 B.n372 B.n371 585
R1137 B.n370 B.n369 585
R1138 B.n368 B.n367 585
R1139 B.n366 B.n365 585
R1140 B.n364 B.n363 585
R1141 B.n362 B.n361 585
R1142 B.n360 B.n359 585
R1143 B.n358 B.n357 585
R1144 B.n356 B.n355 585
R1145 B.n354 B.n353 585
R1146 B.n352 B.n351 585
R1147 B.n350 B.n349 585
R1148 B.n348 B.n347 585
R1149 B.n346 B.n345 585
R1150 B.n344 B.n343 585
R1151 B.n342 B.n341 585
R1152 B.n340 B.n339 585
R1153 B.n338 B.n337 585
R1154 B.n336 B.n335 585
R1155 B.n334 B.n333 585
R1156 B.n332 B.n331 585
R1157 B.n330 B.n329 585
R1158 B.n328 B.n327 585
R1159 B.n326 B.n325 585
R1160 B.n324 B.n323 585
R1161 B.n322 B.n321 585
R1162 B.n320 B.n319 585
R1163 B.n318 B.n317 585
R1164 B.n316 B.n315 585
R1165 B.n314 B.n313 585
R1166 B.n312 B.n311 585
R1167 B.n310 B.n309 585
R1168 B.n308 B.n307 585
R1169 B.n306 B.n305 585
R1170 B.n304 B.n303 585
R1171 B.n302 B.n301 585
R1172 B.n300 B.n299 585
R1173 B.n298 B.n297 585
R1174 B.n296 B.n295 585
R1175 B.n294 B.n293 585
R1176 B.n292 B.n291 585
R1177 B.n290 B.n289 585
R1178 B.n288 B.n287 585
R1179 B.n286 B.n285 585
R1180 B.n284 B.n283 585
R1181 B.n282 B.n281 585
R1182 B.n280 B.n279 585
R1183 B.n278 B.n277 585
R1184 B.n276 B.n275 585
R1185 B.n274 B.n273 585
R1186 B.n272 B.n271 585
R1187 B.n270 B.n269 585
R1188 B.n268 B.n267 585
R1189 B.n266 B.n265 585
R1190 B.n264 B.n263 585
R1191 B.n262 B.n261 585
R1192 B.n260 B.n259 585
R1193 B.n258 B.n257 585
R1194 B.n256 B.n255 585
R1195 B.n254 B.n253 585
R1196 B.n252 B.n251 585
R1197 B.n250 B.n249 585
R1198 B.n248 B.n247 585
R1199 B.n246 B.n245 585
R1200 B.n244 B.n243 585
R1201 B.n242 B.n241 585
R1202 B.n240 B.n239 585
R1203 B.n238 B.n237 585
R1204 B.n236 B.n235 585
R1205 B.n234 B.n233 585
R1206 B.n232 B.n231 585
R1207 B.n230 B.n229 585
R1208 B.n228 B.n227 585
R1209 B.n226 B.n225 585
R1210 B.n224 B.n223 585
R1211 B.n222 B.n221 585
R1212 B.n220 B.n219 585
R1213 B.n218 B.n217 585
R1214 B.n216 B.n215 585
R1215 B.n214 B.n213 585
R1216 B.n212 B.n211 585
R1217 B.n210 B.n209 585
R1218 B.n208 B.n207 585
R1219 B.n206 B.n205 585
R1220 B.n204 B.n203 585
R1221 B.n202 B.n201 585
R1222 B.n200 B.n199 585
R1223 B.n198 B.n197 585
R1224 B.n196 B.n195 585
R1225 B.n1193 B.n125 585
R1226 B.n1198 B.n125 585
R1227 B.n1192 B.n124 585
R1228 B.n1199 B.n124 585
R1229 B.n1191 B.n1190 585
R1230 B.n1190 B.n120 585
R1231 B.n1189 B.n119 585
R1232 B.n1205 B.n119 585
R1233 B.n1188 B.n118 585
R1234 B.n1206 B.n118 585
R1235 B.n1187 B.n117 585
R1236 B.n1207 B.n117 585
R1237 B.n1186 B.n1185 585
R1238 B.n1185 B.n113 585
R1239 B.n1184 B.n112 585
R1240 B.n1213 B.n112 585
R1241 B.n1183 B.n111 585
R1242 B.n1214 B.n111 585
R1243 B.n1182 B.n110 585
R1244 B.n1215 B.n110 585
R1245 B.n1181 B.n1180 585
R1246 B.n1180 B.n106 585
R1247 B.n1179 B.n105 585
R1248 B.n1221 B.n105 585
R1249 B.n1178 B.n104 585
R1250 B.n1222 B.n104 585
R1251 B.n1177 B.n103 585
R1252 B.n1223 B.n103 585
R1253 B.n1176 B.n1175 585
R1254 B.n1175 B.n99 585
R1255 B.n1174 B.n98 585
R1256 B.n1229 B.n98 585
R1257 B.n1173 B.n97 585
R1258 B.n1230 B.n97 585
R1259 B.n1172 B.n96 585
R1260 B.n1231 B.n96 585
R1261 B.n1171 B.n1170 585
R1262 B.n1170 B.n92 585
R1263 B.n1169 B.n91 585
R1264 B.n1237 B.n91 585
R1265 B.n1168 B.n90 585
R1266 B.n1238 B.n90 585
R1267 B.n1167 B.n89 585
R1268 B.n1239 B.n89 585
R1269 B.n1166 B.n1165 585
R1270 B.n1165 B.n85 585
R1271 B.n1164 B.n84 585
R1272 B.n1245 B.n84 585
R1273 B.n1163 B.n83 585
R1274 B.n1246 B.n83 585
R1275 B.n1162 B.n82 585
R1276 B.n1247 B.n82 585
R1277 B.n1161 B.n1160 585
R1278 B.n1160 B.n78 585
R1279 B.n1159 B.n77 585
R1280 B.n1253 B.n77 585
R1281 B.n1158 B.n76 585
R1282 B.n1254 B.n76 585
R1283 B.n1157 B.n75 585
R1284 B.n1255 B.n75 585
R1285 B.n1156 B.n1155 585
R1286 B.n1155 B.n71 585
R1287 B.n1154 B.n70 585
R1288 B.n1261 B.n70 585
R1289 B.n1153 B.n69 585
R1290 B.n1262 B.n69 585
R1291 B.n1152 B.n68 585
R1292 B.n1263 B.n68 585
R1293 B.n1151 B.n1150 585
R1294 B.n1150 B.n64 585
R1295 B.n1149 B.n63 585
R1296 B.n1269 B.n63 585
R1297 B.n1148 B.n62 585
R1298 B.n1270 B.n62 585
R1299 B.n1147 B.n61 585
R1300 B.n1271 B.n61 585
R1301 B.n1146 B.n1145 585
R1302 B.n1145 B.n57 585
R1303 B.n1144 B.n56 585
R1304 B.n1277 B.n56 585
R1305 B.n1143 B.n55 585
R1306 B.n1278 B.n55 585
R1307 B.n1142 B.n54 585
R1308 B.n1279 B.n54 585
R1309 B.n1141 B.n1140 585
R1310 B.n1140 B.n53 585
R1311 B.n1139 B.n49 585
R1312 B.n1285 B.n49 585
R1313 B.n1138 B.n48 585
R1314 B.n1286 B.n48 585
R1315 B.n1137 B.n47 585
R1316 B.n1287 B.n47 585
R1317 B.n1136 B.n1135 585
R1318 B.n1135 B.n43 585
R1319 B.n1134 B.n42 585
R1320 B.n1293 B.n42 585
R1321 B.n1133 B.n41 585
R1322 B.n1294 B.n41 585
R1323 B.n1132 B.n40 585
R1324 B.n1295 B.n40 585
R1325 B.n1131 B.n1130 585
R1326 B.n1130 B.n36 585
R1327 B.n1129 B.n35 585
R1328 B.n1301 B.n35 585
R1329 B.n1128 B.n34 585
R1330 B.n1302 B.n34 585
R1331 B.n1127 B.n33 585
R1332 B.n1303 B.n33 585
R1333 B.n1126 B.n1125 585
R1334 B.n1125 B.n29 585
R1335 B.n1124 B.n28 585
R1336 B.n1309 B.n28 585
R1337 B.n1123 B.n27 585
R1338 B.n1310 B.n27 585
R1339 B.n1122 B.n26 585
R1340 B.n1311 B.n26 585
R1341 B.n1121 B.n1120 585
R1342 B.n1120 B.n22 585
R1343 B.n1119 B.n21 585
R1344 B.n1317 B.n21 585
R1345 B.n1118 B.n20 585
R1346 B.n1318 B.n20 585
R1347 B.n1117 B.n19 585
R1348 B.n1319 B.n19 585
R1349 B.n1116 B.n1115 585
R1350 B.n1115 B.n18 585
R1351 B.n1114 B.n14 585
R1352 B.n1325 B.n14 585
R1353 B.n1113 B.n13 585
R1354 B.n1326 B.n13 585
R1355 B.n1112 B.n12 585
R1356 B.n1327 B.n12 585
R1357 B.n1111 B.n1110 585
R1358 B.n1110 B.n8 585
R1359 B.n1109 B.n7 585
R1360 B.n1333 B.n7 585
R1361 B.n1108 B.n6 585
R1362 B.n1334 B.n6 585
R1363 B.n1107 B.n5 585
R1364 B.n1335 B.n5 585
R1365 B.n1106 B.n1105 585
R1366 B.n1105 B.n4 585
R1367 B.n1104 B.n444 585
R1368 B.n1104 B.n1103 585
R1369 B.n1094 B.n445 585
R1370 B.n446 B.n445 585
R1371 B.n1096 B.n1095 585
R1372 B.n1097 B.n1096 585
R1373 B.n1093 B.n451 585
R1374 B.n451 B.n450 585
R1375 B.n1092 B.n1091 585
R1376 B.n1091 B.n1090 585
R1377 B.n453 B.n452 585
R1378 B.n1083 B.n453 585
R1379 B.n1082 B.n1081 585
R1380 B.n1084 B.n1082 585
R1381 B.n1080 B.n458 585
R1382 B.n458 B.n457 585
R1383 B.n1079 B.n1078 585
R1384 B.n1078 B.n1077 585
R1385 B.n460 B.n459 585
R1386 B.n461 B.n460 585
R1387 B.n1070 B.n1069 585
R1388 B.n1071 B.n1070 585
R1389 B.n1068 B.n466 585
R1390 B.n466 B.n465 585
R1391 B.n1067 B.n1066 585
R1392 B.n1066 B.n1065 585
R1393 B.n468 B.n467 585
R1394 B.n469 B.n468 585
R1395 B.n1058 B.n1057 585
R1396 B.n1059 B.n1058 585
R1397 B.n1056 B.n473 585
R1398 B.n477 B.n473 585
R1399 B.n1055 B.n1054 585
R1400 B.n1054 B.n1053 585
R1401 B.n475 B.n474 585
R1402 B.n476 B.n475 585
R1403 B.n1046 B.n1045 585
R1404 B.n1047 B.n1046 585
R1405 B.n1044 B.n482 585
R1406 B.n482 B.n481 585
R1407 B.n1043 B.n1042 585
R1408 B.n1042 B.n1041 585
R1409 B.n484 B.n483 585
R1410 B.n485 B.n484 585
R1411 B.n1034 B.n1033 585
R1412 B.n1035 B.n1034 585
R1413 B.n1032 B.n490 585
R1414 B.n490 B.n489 585
R1415 B.n1031 B.n1030 585
R1416 B.n1030 B.n1029 585
R1417 B.n492 B.n491 585
R1418 B.n1022 B.n492 585
R1419 B.n1021 B.n1020 585
R1420 B.n1023 B.n1021 585
R1421 B.n1019 B.n497 585
R1422 B.n497 B.n496 585
R1423 B.n1018 B.n1017 585
R1424 B.n1017 B.n1016 585
R1425 B.n499 B.n498 585
R1426 B.n500 B.n499 585
R1427 B.n1009 B.n1008 585
R1428 B.n1010 B.n1009 585
R1429 B.n1007 B.n505 585
R1430 B.n505 B.n504 585
R1431 B.n1006 B.n1005 585
R1432 B.n1005 B.n1004 585
R1433 B.n507 B.n506 585
R1434 B.n508 B.n507 585
R1435 B.n997 B.n996 585
R1436 B.n998 B.n997 585
R1437 B.n995 B.n513 585
R1438 B.n513 B.n512 585
R1439 B.n994 B.n993 585
R1440 B.n993 B.n992 585
R1441 B.n515 B.n514 585
R1442 B.n516 B.n515 585
R1443 B.n985 B.n984 585
R1444 B.n986 B.n985 585
R1445 B.n983 B.n521 585
R1446 B.n521 B.n520 585
R1447 B.n982 B.n981 585
R1448 B.n981 B.n980 585
R1449 B.n523 B.n522 585
R1450 B.n524 B.n523 585
R1451 B.n973 B.n972 585
R1452 B.n974 B.n973 585
R1453 B.n971 B.n529 585
R1454 B.n529 B.n528 585
R1455 B.n970 B.n969 585
R1456 B.n969 B.n968 585
R1457 B.n531 B.n530 585
R1458 B.n532 B.n531 585
R1459 B.n961 B.n960 585
R1460 B.n962 B.n961 585
R1461 B.n959 B.n537 585
R1462 B.n537 B.n536 585
R1463 B.n958 B.n957 585
R1464 B.n957 B.n956 585
R1465 B.n539 B.n538 585
R1466 B.n540 B.n539 585
R1467 B.n949 B.n948 585
R1468 B.n950 B.n949 585
R1469 B.n947 B.n545 585
R1470 B.n545 B.n544 585
R1471 B.n946 B.n945 585
R1472 B.n945 B.n944 585
R1473 B.n547 B.n546 585
R1474 B.n548 B.n547 585
R1475 B.n937 B.n936 585
R1476 B.n938 B.n937 585
R1477 B.n935 B.n553 585
R1478 B.n553 B.n552 585
R1479 B.n934 B.n933 585
R1480 B.n933 B.n932 585
R1481 B.n555 B.n554 585
R1482 B.n556 B.n555 585
R1483 B.n925 B.n924 585
R1484 B.n926 B.n925 585
R1485 B.n923 B.n560 585
R1486 B.n564 B.n560 585
R1487 B.n922 B.n921 585
R1488 B.n921 B.n920 585
R1489 B.n562 B.n561 585
R1490 B.n563 B.n562 585
R1491 B.n913 B.n912 585
R1492 B.n914 B.n913 585
R1493 B.n911 B.n569 585
R1494 B.n569 B.n568 585
R1495 B.n910 B.n909 585
R1496 B.n909 B.n908 585
R1497 B.n571 B.n570 585
R1498 B.n572 B.n571 585
R1499 B.n901 B.n900 585
R1500 B.n902 B.n901 585
R1501 B.n899 B.n577 585
R1502 B.n577 B.n576 585
R1503 B.n894 B.n893 585
R1504 B.n892 B.n642 585
R1505 B.n891 B.n641 585
R1506 B.n896 B.n641 585
R1507 B.n890 B.n889 585
R1508 B.n888 B.n887 585
R1509 B.n886 B.n885 585
R1510 B.n884 B.n883 585
R1511 B.n882 B.n881 585
R1512 B.n880 B.n879 585
R1513 B.n878 B.n877 585
R1514 B.n876 B.n875 585
R1515 B.n874 B.n873 585
R1516 B.n872 B.n871 585
R1517 B.n870 B.n869 585
R1518 B.n868 B.n867 585
R1519 B.n866 B.n865 585
R1520 B.n864 B.n863 585
R1521 B.n862 B.n861 585
R1522 B.n860 B.n859 585
R1523 B.n858 B.n857 585
R1524 B.n856 B.n855 585
R1525 B.n854 B.n853 585
R1526 B.n852 B.n851 585
R1527 B.n850 B.n849 585
R1528 B.n848 B.n847 585
R1529 B.n846 B.n845 585
R1530 B.n844 B.n843 585
R1531 B.n842 B.n841 585
R1532 B.n840 B.n839 585
R1533 B.n838 B.n837 585
R1534 B.n836 B.n835 585
R1535 B.n834 B.n833 585
R1536 B.n832 B.n831 585
R1537 B.n830 B.n829 585
R1538 B.n828 B.n827 585
R1539 B.n826 B.n825 585
R1540 B.n824 B.n823 585
R1541 B.n822 B.n821 585
R1542 B.n820 B.n819 585
R1543 B.n818 B.n817 585
R1544 B.n816 B.n815 585
R1545 B.n814 B.n813 585
R1546 B.n812 B.n811 585
R1547 B.n810 B.n809 585
R1548 B.n808 B.n807 585
R1549 B.n806 B.n805 585
R1550 B.n804 B.n803 585
R1551 B.n802 B.n801 585
R1552 B.n800 B.n799 585
R1553 B.n798 B.n797 585
R1554 B.n796 B.n795 585
R1555 B.n794 B.n793 585
R1556 B.n792 B.n791 585
R1557 B.n790 B.n789 585
R1558 B.n788 B.n787 585
R1559 B.n786 B.n785 585
R1560 B.n784 B.n783 585
R1561 B.n782 B.n781 585
R1562 B.n779 B.n778 585
R1563 B.n777 B.n776 585
R1564 B.n775 B.n774 585
R1565 B.n773 B.n772 585
R1566 B.n771 B.n770 585
R1567 B.n769 B.n768 585
R1568 B.n767 B.n766 585
R1569 B.n765 B.n764 585
R1570 B.n763 B.n762 585
R1571 B.n761 B.n760 585
R1572 B.n758 B.n757 585
R1573 B.n756 B.n755 585
R1574 B.n754 B.n753 585
R1575 B.n752 B.n751 585
R1576 B.n750 B.n749 585
R1577 B.n748 B.n747 585
R1578 B.n746 B.n745 585
R1579 B.n744 B.n743 585
R1580 B.n742 B.n741 585
R1581 B.n740 B.n739 585
R1582 B.n738 B.n737 585
R1583 B.n736 B.n735 585
R1584 B.n734 B.n733 585
R1585 B.n732 B.n731 585
R1586 B.n730 B.n729 585
R1587 B.n728 B.n727 585
R1588 B.n726 B.n725 585
R1589 B.n724 B.n723 585
R1590 B.n722 B.n721 585
R1591 B.n720 B.n719 585
R1592 B.n718 B.n717 585
R1593 B.n716 B.n715 585
R1594 B.n714 B.n713 585
R1595 B.n712 B.n711 585
R1596 B.n710 B.n709 585
R1597 B.n708 B.n707 585
R1598 B.n706 B.n705 585
R1599 B.n704 B.n703 585
R1600 B.n702 B.n701 585
R1601 B.n700 B.n699 585
R1602 B.n698 B.n697 585
R1603 B.n696 B.n695 585
R1604 B.n694 B.n693 585
R1605 B.n692 B.n691 585
R1606 B.n690 B.n689 585
R1607 B.n688 B.n687 585
R1608 B.n686 B.n685 585
R1609 B.n684 B.n683 585
R1610 B.n682 B.n681 585
R1611 B.n680 B.n679 585
R1612 B.n678 B.n677 585
R1613 B.n676 B.n675 585
R1614 B.n674 B.n673 585
R1615 B.n672 B.n671 585
R1616 B.n670 B.n669 585
R1617 B.n668 B.n667 585
R1618 B.n666 B.n665 585
R1619 B.n664 B.n663 585
R1620 B.n662 B.n661 585
R1621 B.n660 B.n659 585
R1622 B.n658 B.n657 585
R1623 B.n656 B.n655 585
R1624 B.n654 B.n653 585
R1625 B.n652 B.n651 585
R1626 B.n650 B.n649 585
R1627 B.n648 B.n647 585
R1628 B.n579 B.n578 585
R1629 B.n898 B.n897 585
R1630 B.n897 B.n896 585
R1631 B.n575 B.n574 585
R1632 B.n576 B.n575 585
R1633 B.n904 B.n903 585
R1634 B.n903 B.n902 585
R1635 B.n905 B.n573 585
R1636 B.n573 B.n572 585
R1637 B.n907 B.n906 585
R1638 B.n908 B.n907 585
R1639 B.n567 B.n566 585
R1640 B.n568 B.n567 585
R1641 B.n916 B.n915 585
R1642 B.n915 B.n914 585
R1643 B.n917 B.n565 585
R1644 B.n565 B.n563 585
R1645 B.n919 B.n918 585
R1646 B.n920 B.n919 585
R1647 B.n559 B.n558 585
R1648 B.n564 B.n559 585
R1649 B.n928 B.n927 585
R1650 B.n927 B.n926 585
R1651 B.n929 B.n557 585
R1652 B.n557 B.n556 585
R1653 B.n931 B.n930 585
R1654 B.n932 B.n931 585
R1655 B.n551 B.n550 585
R1656 B.n552 B.n551 585
R1657 B.n940 B.n939 585
R1658 B.n939 B.n938 585
R1659 B.n941 B.n549 585
R1660 B.n549 B.n548 585
R1661 B.n943 B.n942 585
R1662 B.n944 B.n943 585
R1663 B.n543 B.n542 585
R1664 B.n544 B.n543 585
R1665 B.n952 B.n951 585
R1666 B.n951 B.n950 585
R1667 B.n953 B.n541 585
R1668 B.n541 B.n540 585
R1669 B.n955 B.n954 585
R1670 B.n956 B.n955 585
R1671 B.n535 B.n534 585
R1672 B.n536 B.n535 585
R1673 B.n964 B.n963 585
R1674 B.n963 B.n962 585
R1675 B.n965 B.n533 585
R1676 B.n533 B.n532 585
R1677 B.n967 B.n966 585
R1678 B.n968 B.n967 585
R1679 B.n527 B.n526 585
R1680 B.n528 B.n527 585
R1681 B.n976 B.n975 585
R1682 B.n975 B.n974 585
R1683 B.n977 B.n525 585
R1684 B.n525 B.n524 585
R1685 B.n979 B.n978 585
R1686 B.n980 B.n979 585
R1687 B.n519 B.n518 585
R1688 B.n520 B.n519 585
R1689 B.n988 B.n987 585
R1690 B.n987 B.n986 585
R1691 B.n989 B.n517 585
R1692 B.n517 B.n516 585
R1693 B.n991 B.n990 585
R1694 B.n992 B.n991 585
R1695 B.n511 B.n510 585
R1696 B.n512 B.n511 585
R1697 B.n1000 B.n999 585
R1698 B.n999 B.n998 585
R1699 B.n1001 B.n509 585
R1700 B.n509 B.n508 585
R1701 B.n1003 B.n1002 585
R1702 B.n1004 B.n1003 585
R1703 B.n503 B.n502 585
R1704 B.n504 B.n503 585
R1705 B.n1012 B.n1011 585
R1706 B.n1011 B.n1010 585
R1707 B.n1013 B.n501 585
R1708 B.n501 B.n500 585
R1709 B.n1015 B.n1014 585
R1710 B.n1016 B.n1015 585
R1711 B.n495 B.n494 585
R1712 B.n496 B.n495 585
R1713 B.n1025 B.n1024 585
R1714 B.n1024 B.n1023 585
R1715 B.n1026 B.n493 585
R1716 B.n1022 B.n493 585
R1717 B.n1028 B.n1027 585
R1718 B.n1029 B.n1028 585
R1719 B.n488 B.n487 585
R1720 B.n489 B.n488 585
R1721 B.n1037 B.n1036 585
R1722 B.n1036 B.n1035 585
R1723 B.n1038 B.n486 585
R1724 B.n486 B.n485 585
R1725 B.n1040 B.n1039 585
R1726 B.n1041 B.n1040 585
R1727 B.n480 B.n479 585
R1728 B.n481 B.n480 585
R1729 B.n1049 B.n1048 585
R1730 B.n1048 B.n1047 585
R1731 B.n1050 B.n478 585
R1732 B.n478 B.n476 585
R1733 B.n1052 B.n1051 585
R1734 B.n1053 B.n1052 585
R1735 B.n472 B.n471 585
R1736 B.n477 B.n472 585
R1737 B.n1061 B.n1060 585
R1738 B.n1060 B.n1059 585
R1739 B.n1062 B.n470 585
R1740 B.n470 B.n469 585
R1741 B.n1064 B.n1063 585
R1742 B.n1065 B.n1064 585
R1743 B.n464 B.n463 585
R1744 B.n465 B.n464 585
R1745 B.n1073 B.n1072 585
R1746 B.n1072 B.n1071 585
R1747 B.n1074 B.n462 585
R1748 B.n462 B.n461 585
R1749 B.n1076 B.n1075 585
R1750 B.n1077 B.n1076 585
R1751 B.n456 B.n455 585
R1752 B.n457 B.n456 585
R1753 B.n1086 B.n1085 585
R1754 B.n1085 B.n1084 585
R1755 B.n1087 B.n454 585
R1756 B.n1083 B.n454 585
R1757 B.n1089 B.n1088 585
R1758 B.n1090 B.n1089 585
R1759 B.n449 B.n448 585
R1760 B.n450 B.n449 585
R1761 B.n1099 B.n1098 585
R1762 B.n1098 B.n1097 585
R1763 B.n1100 B.n447 585
R1764 B.n447 B.n446 585
R1765 B.n1102 B.n1101 585
R1766 B.n1103 B.n1102 585
R1767 B.n2 B.n0 585
R1768 B.n4 B.n2 585
R1769 B.n3 B.n1 585
R1770 B.n1334 B.n3 585
R1771 B.n1332 B.n1331 585
R1772 B.n1333 B.n1332 585
R1773 B.n1330 B.n9 585
R1774 B.n9 B.n8 585
R1775 B.n1329 B.n1328 585
R1776 B.n1328 B.n1327 585
R1777 B.n11 B.n10 585
R1778 B.n1326 B.n11 585
R1779 B.n1324 B.n1323 585
R1780 B.n1325 B.n1324 585
R1781 B.n1322 B.n15 585
R1782 B.n18 B.n15 585
R1783 B.n1321 B.n1320 585
R1784 B.n1320 B.n1319 585
R1785 B.n17 B.n16 585
R1786 B.n1318 B.n17 585
R1787 B.n1316 B.n1315 585
R1788 B.n1317 B.n1316 585
R1789 B.n1314 B.n23 585
R1790 B.n23 B.n22 585
R1791 B.n1313 B.n1312 585
R1792 B.n1312 B.n1311 585
R1793 B.n25 B.n24 585
R1794 B.n1310 B.n25 585
R1795 B.n1308 B.n1307 585
R1796 B.n1309 B.n1308 585
R1797 B.n1306 B.n30 585
R1798 B.n30 B.n29 585
R1799 B.n1305 B.n1304 585
R1800 B.n1304 B.n1303 585
R1801 B.n32 B.n31 585
R1802 B.n1302 B.n32 585
R1803 B.n1300 B.n1299 585
R1804 B.n1301 B.n1300 585
R1805 B.n1298 B.n37 585
R1806 B.n37 B.n36 585
R1807 B.n1297 B.n1296 585
R1808 B.n1296 B.n1295 585
R1809 B.n39 B.n38 585
R1810 B.n1294 B.n39 585
R1811 B.n1292 B.n1291 585
R1812 B.n1293 B.n1292 585
R1813 B.n1290 B.n44 585
R1814 B.n44 B.n43 585
R1815 B.n1289 B.n1288 585
R1816 B.n1288 B.n1287 585
R1817 B.n46 B.n45 585
R1818 B.n1286 B.n46 585
R1819 B.n1284 B.n1283 585
R1820 B.n1285 B.n1284 585
R1821 B.n1282 B.n50 585
R1822 B.n53 B.n50 585
R1823 B.n1281 B.n1280 585
R1824 B.n1280 B.n1279 585
R1825 B.n52 B.n51 585
R1826 B.n1278 B.n52 585
R1827 B.n1276 B.n1275 585
R1828 B.n1277 B.n1276 585
R1829 B.n1274 B.n58 585
R1830 B.n58 B.n57 585
R1831 B.n1273 B.n1272 585
R1832 B.n1272 B.n1271 585
R1833 B.n60 B.n59 585
R1834 B.n1270 B.n60 585
R1835 B.n1268 B.n1267 585
R1836 B.n1269 B.n1268 585
R1837 B.n1266 B.n65 585
R1838 B.n65 B.n64 585
R1839 B.n1265 B.n1264 585
R1840 B.n1264 B.n1263 585
R1841 B.n67 B.n66 585
R1842 B.n1262 B.n67 585
R1843 B.n1260 B.n1259 585
R1844 B.n1261 B.n1260 585
R1845 B.n1258 B.n72 585
R1846 B.n72 B.n71 585
R1847 B.n1257 B.n1256 585
R1848 B.n1256 B.n1255 585
R1849 B.n74 B.n73 585
R1850 B.n1254 B.n74 585
R1851 B.n1252 B.n1251 585
R1852 B.n1253 B.n1252 585
R1853 B.n1250 B.n79 585
R1854 B.n79 B.n78 585
R1855 B.n1249 B.n1248 585
R1856 B.n1248 B.n1247 585
R1857 B.n81 B.n80 585
R1858 B.n1246 B.n81 585
R1859 B.n1244 B.n1243 585
R1860 B.n1245 B.n1244 585
R1861 B.n1242 B.n86 585
R1862 B.n86 B.n85 585
R1863 B.n1241 B.n1240 585
R1864 B.n1240 B.n1239 585
R1865 B.n88 B.n87 585
R1866 B.n1238 B.n88 585
R1867 B.n1236 B.n1235 585
R1868 B.n1237 B.n1236 585
R1869 B.n1234 B.n93 585
R1870 B.n93 B.n92 585
R1871 B.n1233 B.n1232 585
R1872 B.n1232 B.n1231 585
R1873 B.n95 B.n94 585
R1874 B.n1230 B.n95 585
R1875 B.n1228 B.n1227 585
R1876 B.n1229 B.n1228 585
R1877 B.n1226 B.n100 585
R1878 B.n100 B.n99 585
R1879 B.n1225 B.n1224 585
R1880 B.n1224 B.n1223 585
R1881 B.n102 B.n101 585
R1882 B.n1222 B.n102 585
R1883 B.n1220 B.n1219 585
R1884 B.n1221 B.n1220 585
R1885 B.n1218 B.n107 585
R1886 B.n107 B.n106 585
R1887 B.n1217 B.n1216 585
R1888 B.n1216 B.n1215 585
R1889 B.n109 B.n108 585
R1890 B.n1214 B.n109 585
R1891 B.n1212 B.n1211 585
R1892 B.n1213 B.n1212 585
R1893 B.n1210 B.n114 585
R1894 B.n114 B.n113 585
R1895 B.n1209 B.n1208 585
R1896 B.n1208 B.n1207 585
R1897 B.n116 B.n115 585
R1898 B.n1206 B.n116 585
R1899 B.n1204 B.n1203 585
R1900 B.n1205 B.n1204 585
R1901 B.n1202 B.n121 585
R1902 B.n121 B.n120 585
R1903 B.n1201 B.n1200 585
R1904 B.n1200 B.n1199 585
R1905 B.n123 B.n122 585
R1906 B.n1198 B.n123 585
R1907 B.n1337 B.n1336 585
R1908 B.n1336 B.n1335 585
R1909 B.n894 B.n575 468.476
R1910 B.n195 B.n123 468.476
R1911 B.n897 B.n577 468.476
R1912 B.n1195 B.n125 468.476
R1913 B.n645 B.t17 445.332
R1914 B.n189 B.t12 445.332
R1915 B.n643 B.t20 445.332
R1916 B.n192 B.t22 445.332
R1917 B.n646 B.t16 378.423
R1918 B.n190 B.t13 378.423
R1919 B.n644 B.t19 378.423
R1920 B.n193 B.t23 378.423
R1921 B.n645 B.t14 344.51
R1922 B.n643 B.t18 344.51
R1923 B.n192 B.t21 344.51
R1924 B.n189 B.t10 344.51
R1925 B.n1197 B.n1196 256.663
R1926 B.n1197 B.n187 256.663
R1927 B.n1197 B.n186 256.663
R1928 B.n1197 B.n185 256.663
R1929 B.n1197 B.n184 256.663
R1930 B.n1197 B.n183 256.663
R1931 B.n1197 B.n182 256.663
R1932 B.n1197 B.n181 256.663
R1933 B.n1197 B.n180 256.663
R1934 B.n1197 B.n179 256.663
R1935 B.n1197 B.n178 256.663
R1936 B.n1197 B.n177 256.663
R1937 B.n1197 B.n176 256.663
R1938 B.n1197 B.n175 256.663
R1939 B.n1197 B.n174 256.663
R1940 B.n1197 B.n173 256.663
R1941 B.n1197 B.n172 256.663
R1942 B.n1197 B.n171 256.663
R1943 B.n1197 B.n170 256.663
R1944 B.n1197 B.n169 256.663
R1945 B.n1197 B.n168 256.663
R1946 B.n1197 B.n167 256.663
R1947 B.n1197 B.n166 256.663
R1948 B.n1197 B.n165 256.663
R1949 B.n1197 B.n164 256.663
R1950 B.n1197 B.n163 256.663
R1951 B.n1197 B.n162 256.663
R1952 B.n1197 B.n161 256.663
R1953 B.n1197 B.n160 256.663
R1954 B.n1197 B.n159 256.663
R1955 B.n1197 B.n158 256.663
R1956 B.n1197 B.n157 256.663
R1957 B.n1197 B.n156 256.663
R1958 B.n1197 B.n155 256.663
R1959 B.n1197 B.n154 256.663
R1960 B.n1197 B.n153 256.663
R1961 B.n1197 B.n152 256.663
R1962 B.n1197 B.n151 256.663
R1963 B.n1197 B.n150 256.663
R1964 B.n1197 B.n149 256.663
R1965 B.n1197 B.n148 256.663
R1966 B.n1197 B.n147 256.663
R1967 B.n1197 B.n146 256.663
R1968 B.n1197 B.n145 256.663
R1969 B.n1197 B.n144 256.663
R1970 B.n1197 B.n143 256.663
R1971 B.n1197 B.n142 256.663
R1972 B.n1197 B.n141 256.663
R1973 B.n1197 B.n140 256.663
R1974 B.n1197 B.n139 256.663
R1975 B.n1197 B.n138 256.663
R1976 B.n1197 B.n137 256.663
R1977 B.n1197 B.n136 256.663
R1978 B.n1197 B.n135 256.663
R1979 B.n1197 B.n134 256.663
R1980 B.n1197 B.n133 256.663
R1981 B.n1197 B.n132 256.663
R1982 B.n1197 B.n131 256.663
R1983 B.n1197 B.n130 256.663
R1984 B.n1197 B.n129 256.663
R1985 B.n1197 B.n128 256.663
R1986 B.n1197 B.n127 256.663
R1987 B.n1197 B.n126 256.663
R1988 B.n896 B.n895 256.663
R1989 B.n896 B.n580 256.663
R1990 B.n896 B.n581 256.663
R1991 B.n896 B.n582 256.663
R1992 B.n896 B.n583 256.663
R1993 B.n896 B.n584 256.663
R1994 B.n896 B.n585 256.663
R1995 B.n896 B.n586 256.663
R1996 B.n896 B.n587 256.663
R1997 B.n896 B.n588 256.663
R1998 B.n896 B.n589 256.663
R1999 B.n896 B.n590 256.663
R2000 B.n896 B.n591 256.663
R2001 B.n896 B.n592 256.663
R2002 B.n896 B.n593 256.663
R2003 B.n896 B.n594 256.663
R2004 B.n896 B.n595 256.663
R2005 B.n896 B.n596 256.663
R2006 B.n896 B.n597 256.663
R2007 B.n896 B.n598 256.663
R2008 B.n896 B.n599 256.663
R2009 B.n896 B.n600 256.663
R2010 B.n896 B.n601 256.663
R2011 B.n896 B.n602 256.663
R2012 B.n896 B.n603 256.663
R2013 B.n896 B.n604 256.663
R2014 B.n896 B.n605 256.663
R2015 B.n896 B.n606 256.663
R2016 B.n896 B.n607 256.663
R2017 B.n896 B.n608 256.663
R2018 B.n896 B.n609 256.663
R2019 B.n896 B.n610 256.663
R2020 B.n896 B.n611 256.663
R2021 B.n896 B.n612 256.663
R2022 B.n896 B.n613 256.663
R2023 B.n896 B.n614 256.663
R2024 B.n896 B.n615 256.663
R2025 B.n896 B.n616 256.663
R2026 B.n896 B.n617 256.663
R2027 B.n896 B.n618 256.663
R2028 B.n896 B.n619 256.663
R2029 B.n896 B.n620 256.663
R2030 B.n896 B.n621 256.663
R2031 B.n896 B.n622 256.663
R2032 B.n896 B.n623 256.663
R2033 B.n896 B.n624 256.663
R2034 B.n896 B.n625 256.663
R2035 B.n896 B.n626 256.663
R2036 B.n896 B.n627 256.663
R2037 B.n896 B.n628 256.663
R2038 B.n896 B.n629 256.663
R2039 B.n896 B.n630 256.663
R2040 B.n896 B.n631 256.663
R2041 B.n896 B.n632 256.663
R2042 B.n896 B.n633 256.663
R2043 B.n896 B.n634 256.663
R2044 B.n896 B.n635 256.663
R2045 B.n896 B.n636 256.663
R2046 B.n896 B.n637 256.663
R2047 B.n896 B.n638 256.663
R2048 B.n896 B.n639 256.663
R2049 B.n896 B.n640 256.663
R2050 B.n903 B.n575 163.367
R2051 B.n903 B.n573 163.367
R2052 B.n907 B.n573 163.367
R2053 B.n907 B.n567 163.367
R2054 B.n915 B.n567 163.367
R2055 B.n915 B.n565 163.367
R2056 B.n919 B.n565 163.367
R2057 B.n919 B.n559 163.367
R2058 B.n927 B.n559 163.367
R2059 B.n927 B.n557 163.367
R2060 B.n931 B.n557 163.367
R2061 B.n931 B.n551 163.367
R2062 B.n939 B.n551 163.367
R2063 B.n939 B.n549 163.367
R2064 B.n943 B.n549 163.367
R2065 B.n943 B.n543 163.367
R2066 B.n951 B.n543 163.367
R2067 B.n951 B.n541 163.367
R2068 B.n955 B.n541 163.367
R2069 B.n955 B.n535 163.367
R2070 B.n963 B.n535 163.367
R2071 B.n963 B.n533 163.367
R2072 B.n967 B.n533 163.367
R2073 B.n967 B.n527 163.367
R2074 B.n975 B.n527 163.367
R2075 B.n975 B.n525 163.367
R2076 B.n979 B.n525 163.367
R2077 B.n979 B.n519 163.367
R2078 B.n987 B.n519 163.367
R2079 B.n987 B.n517 163.367
R2080 B.n991 B.n517 163.367
R2081 B.n991 B.n511 163.367
R2082 B.n999 B.n511 163.367
R2083 B.n999 B.n509 163.367
R2084 B.n1003 B.n509 163.367
R2085 B.n1003 B.n503 163.367
R2086 B.n1011 B.n503 163.367
R2087 B.n1011 B.n501 163.367
R2088 B.n1015 B.n501 163.367
R2089 B.n1015 B.n495 163.367
R2090 B.n1024 B.n495 163.367
R2091 B.n1024 B.n493 163.367
R2092 B.n1028 B.n493 163.367
R2093 B.n1028 B.n488 163.367
R2094 B.n1036 B.n488 163.367
R2095 B.n1036 B.n486 163.367
R2096 B.n1040 B.n486 163.367
R2097 B.n1040 B.n480 163.367
R2098 B.n1048 B.n480 163.367
R2099 B.n1048 B.n478 163.367
R2100 B.n1052 B.n478 163.367
R2101 B.n1052 B.n472 163.367
R2102 B.n1060 B.n472 163.367
R2103 B.n1060 B.n470 163.367
R2104 B.n1064 B.n470 163.367
R2105 B.n1064 B.n464 163.367
R2106 B.n1072 B.n464 163.367
R2107 B.n1072 B.n462 163.367
R2108 B.n1076 B.n462 163.367
R2109 B.n1076 B.n456 163.367
R2110 B.n1085 B.n456 163.367
R2111 B.n1085 B.n454 163.367
R2112 B.n1089 B.n454 163.367
R2113 B.n1089 B.n449 163.367
R2114 B.n1098 B.n449 163.367
R2115 B.n1098 B.n447 163.367
R2116 B.n1102 B.n447 163.367
R2117 B.n1102 B.n2 163.367
R2118 B.n1336 B.n2 163.367
R2119 B.n1336 B.n3 163.367
R2120 B.n1332 B.n3 163.367
R2121 B.n1332 B.n9 163.367
R2122 B.n1328 B.n9 163.367
R2123 B.n1328 B.n11 163.367
R2124 B.n1324 B.n11 163.367
R2125 B.n1324 B.n15 163.367
R2126 B.n1320 B.n15 163.367
R2127 B.n1320 B.n17 163.367
R2128 B.n1316 B.n17 163.367
R2129 B.n1316 B.n23 163.367
R2130 B.n1312 B.n23 163.367
R2131 B.n1312 B.n25 163.367
R2132 B.n1308 B.n25 163.367
R2133 B.n1308 B.n30 163.367
R2134 B.n1304 B.n30 163.367
R2135 B.n1304 B.n32 163.367
R2136 B.n1300 B.n32 163.367
R2137 B.n1300 B.n37 163.367
R2138 B.n1296 B.n37 163.367
R2139 B.n1296 B.n39 163.367
R2140 B.n1292 B.n39 163.367
R2141 B.n1292 B.n44 163.367
R2142 B.n1288 B.n44 163.367
R2143 B.n1288 B.n46 163.367
R2144 B.n1284 B.n46 163.367
R2145 B.n1284 B.n50 163.367
R2146 B.n1280 B.n50 163.367
R2147 B.n1280 B.n52 163.367
R2148 B.n1276 B.n52 163.367
R2149 B.n1276 B.n58 163.367
R2150 B.n1272 B.n58 163.367
R2151 B.n1272 B.n60 163.367
R2152 B.n1268 B.n60 163.367
R2153 B.n1268 B.n65 163.367
R2154 B.n1264 B.n65 163.367
R2155 B.n1264 B.n67 163.367
R2156 B.n1260 B.n67 163.367
R2157 B.n1260 B.n72 163.367
R2158 B.n1256 B.n72 163.367
R2159 B.n1256 B.n74 163.367
R2160 B.n1252 B.n74 163.367
R2161 B.n1252 B.n79 163.367
R2162 B.n1248 B.n79 163.367
R2163 B.n1248 B.n81 163.367
R2164 B.n1244 B.n81 163.367
R2165 B.n1244 B.n86 163.367
R2166 B.n1240 B.n86 163.367
R2167 B.n1240 B.n88 163.367
R2168 B.n1236 B.n88 163.367
R2169 B.n1236 B.n93 163.367
R2170 B.n1232 B.n93 163.367
R2171 B.n1232 B.n95 163.367
R2172 B.n1228 B.n95 163.367
R2173 B.n1228 B.n100 163.367
R2174 B.n1224 B.n100 163.367
R2175 B.n1224 B.n102 163.367
R2176 B.n1220 B.n102 163.367
R2177 B.n1220 B.n107 163.367
R2178 B.n1216 B.n107 163.367
R2179 B.n1216 B.n109 163.367
R2180 B.n1212 B.n109 163.367
R2181 B.n1212 B.n114 163.367
R2182 B.n1208 B.n114 163.367
R2183 B.n1208 B.n116 163.367
R2184 B.n1204 B.n116 163.367
R2185 B.n1204 B.n121 163.367
R2186 B.n1200 B.n121 163.367
R2187 B.n1200 B.n123 163.367
R2188 B.n642 B.n641 163.367
R2189 B.n889 B.n641 163.367
R2190 B.n887 B.n886 163.367
R2191 B.n883 B.n882 163.367
R2192 B.n879 B.n878 163.367
R2193 B.n875 B.n874 163.367
R2194 B.n871 B.n870 163.367
R2195 B.n867 B.n866 163.367
R2196 B.n863 B.n862 163.367
R2197 B.n859 B.n858 163.367
R2198 B.n855 B.n854 163.367
R2199 B.n851 B.n850 163.367
R2200 B.n847 B.n846 163.367
R2201 B.n843 B.n842 163.367
R2202 B.n839 B.n838 163.367
R2203 B.n835 B.n834 163.367
R2204 B.n831 B.n830 163.367
R2205 B.n827 B.n826 163.367
R2206 B.n823 B.n822 163.367
R2207 B.n819 B.n818 163.367
R2208 B.n815 B.n814 163.367
R2209 B.n811 B.n810 163.367
R2210 B.n807 B.n806 163.367
R2211 B.n803 B.n802 163.367
R2212 B.n799 B.n798 163.367
R2213 B.n795 B.n794 163.367
R2214 B.n791 B.n790 163.367
R2215 B.n787 B.n786 163.367
R2216 B.n783 B.n782 163.367
R2217 B.n778 B.n777 163.367
R2218 B.n774 B.n773 163.367
R2219 B.n770 B.n769 163.367
R2220 B.n766 B.n765 163.367
R2221 B.n762 B.n761 163.367
R2222 B.n757 B.n756 163.367
R2223 B.n753 B.n752 163.367
R2224 B.n749 B.n748 163.367
R2225 B.n745 B.n744 163.367
R2226 B.n741 B.n740 163.367
R2227 B.n737 B.n736 163.367
R2228 B.n733 B.n732 163.367
R2229 B.n729 B.n728 163.367
R2230 B.n725 B.n724 163.367
R2231 B.n721 B.n720 163.367
R2232 B.n717 B.n716 163.367
R2233 B.n713 B.n712 163.367
R2234 B.n709 B.n708 163.367
R2235 B.n705 B.n704 163.367
R2236 B.n701 B.n700 163.367
R2237 B.n697 B.n696 163.367
R2238 B.n693 B.n692 163.367
R2239 B.n689 B.n688 163.367
R2240 B.n685 B.n684 163.367
R2241 B.n681 B.n680 163.367
R2242 B.n677 B.n676 163.367
R2243 B.n673 B.n672 163.367
R2244 B.n669 B.n668 163.367
R2245 B.n665 B.n664 163.367
R2246 B.n661 B.n660 163.367
R2247 B.n657 B.n656 163.367
R2248 B.n653 B.n652 163.367
R2249 B.n649 B.n648 163.367
R2250 B.n897 B.n579 163.367
R2251 B.n901 B.n577 163.367
R2252 B.n901 B.n571 163.367
R2253 B.n909 B.n571 163.367
R2254 B.n909 B.n569 163.367
R2255 B.n913 B.n569 163.367
R2256 B.n913 B.n562 163.367
R2257 B.n921 B.n562 163.367
R2258 B.n921 B.n560 163.367
R2259 B.n925 B.n560 163.367
R2260 B.n925 B.n555 163.367
R2261 B.n933 B.n555 163.367
R2262 B.n933 B.n553 163.367
R2263 B.n937 B.n553 163.367
R2264 B.n937 B.n547 163.367
R2265 B.n945 B.n547 163.367
R2266 B.n945 B.n545 163.367
R2267 B.n949 B.n545 163.367
R2268 B.n949 B.n539 163.367
R2269 B.n957 B.n539 163.367
R2270 B.n957 B.n537 163.367
R2271 B.n961 B.n537 163.367
R2272 B.n961 B.n531 163.367
R2273 B.n969 B.n531 163.367
R2274 B.n969 B.n529 163.367
R2275 B.n973 B.n529 163.367
R2276 B.n973 B.n523 163.367
R2277 B.n981 B.n523 163.367
R2278 B.n981 B.n521 163.367
R2279 B.n985 B.n521 163.367
R2280 B.n985 B.n515 163.367
R2281 B.n993 B.n515 163.367
R2282 B.n993 B.n513 163.367
R2283 B.n997 B.n513 163.367
R2284 B.n997 B.n507 163.367
R2285 B.n1005 B.n507 163.367
R2286 B.n1005 B.n505 163.367
R2287 B.n1009 B.n505 163.367
R2288 B.n1009 B.n499 163.367
R2289 B.n1017 B.n499 163.367
R2290 B.n1017 B.n497 163.367
R2291 B.n1021 B.n497 163.367
R2292 B.n1021 B.n492 163.367
R2293 B.n1030 B.n492 163.367
R2294 B.n1030 B.n490 163.367
R2295 B.n1034 B.n490 163.367
R2296 B.n1034 B.n484 163.367
R2297 B.n1042 B.n484 163.367
R2298 B.n1042 B.n482 163.367
R2299 B.n1046 B.n482 163.367
R2300 B.n1046 B.n475 163.367
R2301 B.n1054 B.n475 163.367
R2302 B.n1054 B.n473 163.367
R2303 B.n1058 B.n473 163.367
R2304 B.n1058 B.n468 163.367
R2305 B.n1066 B.n468 163.367
R2306 B.n1066 B.n466 163.367
R2307 B.n1070 B.n466 163.367
R2308 B.n1070 B.n460 163.367
R2309 B.n1078 B.n460 163.367
R2310 B.n1078 B.n458 163.367
R2311 B.n1082 B.n458 163.367
R2312 B.n1082 B.n453 163.367
R2313 B.n1091 B.n453 163.367
R2314 B.n1091 B.n451 163.367
R2315 B.n1096 B.n451 163.367
R2316 B.n1096 B.n445 163.367
R2317 B.n1104 B.n445 163.367
R2318 B.n1105 B.n1104 163.367
R2319 B.n1105 B.n5 163.367
R2320 B.n6 B.n5 163.367
R2321 B.n7 B.n6 163.367
R2322 B.n1110 B.n7 163.367
R2323 B.n1110 B.n12 163.367
R2324 B.n13 B.n12 163.367
R2325 B.n14 B.n13 163.367
R2326 B.n1115 B.n14 163.367
R2327 B.n1115 B.n19 163.367
R2328 B.n20 B.n19 163.367
R2329 B.n21 B.n20 163.367
R2330 B.n1120 B.n21 163.367
R2331 B.n1120 B.n26 163.367
R2332 B.n27 B.n26 163.367
R2333 B.n28 B.n27 163.367
R2334 B.n1125 B.n28 163.367
R2335 B.n1125 B.n33 163.367
R2336 B.n34 B.n33 163.367
R2337 B.n35 B.n34 163.367
R2338 B.n1130 B.n35 163.367
R2339 B.n1130 B.n40 163.367
R2340 B.n41 B.n40 163.367
R2341 B.n42 B.n41 163.367
R2342 B.n1135 B.n42 163.367
R2343 B.n1135 B.n47 163.367
R2344 B.n48 B.n47 163.367
R2345 B.n49 B.n48 163.367
R2346 B.n1140 B.n49 163.367
R2347 B.n1140 B.n54 163.367
R2348 B.n55 B.n54 163.367
R2349 B.n56 B.n55 163.367
R2350 B.n1145 B.n56 163.367
R2351 B.n1145 B.n61 163.367
R2352 B.n62 B.n61 163.367
R2353 B.n63 B.n62 163.367
R2354 B.n1150 B.n63 163.367
R2355 B.n1150 B.n68 163.367
R2356 B.n69 B.n68 163.367
R2357 B.n70 B.n69 163.367
R2358 B.n1155 B.n70 163.367
R2359 B.n1155 B.n75 163.367
R2360 B.n76 B.n75 163.367
R2361 B.n77 B.n76 163.367
R2362 B.n1160 B.n77 163.367
R2363 B.n1160 B.n82 163.367
R2364 B.n83 B.n82 163.367
R2365 B.n84 B.n83 163.367
R2366 B.n1165 B.n84 163.367
R2367 B.n1165 B.n89 163.367
R2368 B.n90 B.n89 163.367
R2369 B.n91 B.n90 163.367
R2370 B.n1170 B.n91 163.367
R2371 B.n1170 B.n96 163.367
R2372 B.n97 B.n96 163.367
R2373 B.n98 B.n97 163.367
R2374 B.n1175 B.n98 163.367
R2375 B.n1175 B.n103 163.367
R2376 B.n104 B.n103 163.367
R2377 B.n105 B.n104 163.367
R2378 B.n1180 B.n105 163.367
R2379 B.n1180 B.n110 163.367
R2380 B.n111 B.n110 163.367
R2381 B.n112 B.n111 163.367
R2382 B.n1185 B.n112 163.367
R2383 B.n1185 B.n117 163.367
R2384 B.n118 B.n117 163.367
R2385 B.n119 B.n118 163.367
R2386 B.n1190 B.n119 163.367
R2387 B.n1190 B.n124 163.367
R2388 B.n125 B.n124 163.367
R2389 B.n199 B.n198 163.367
R2390 B.n203 B.n202 163.367
R2391 B.n207 B.n206 163.367
R2392 B.n211 B.n210 163.367
R2393 B.n215 B.n214 163.367
R2394 B.n219 B.n218 163.367
R2395 B.n223 B.n222 163.367
R2396 B.n227 B.n226 163.367
R2397 B.n231 B.n230 163.367
R2398 B.n235 B.n234 163.367
R2399 B.n239 B.n238 163.367
R2400 B.n243 B.n242 163.367
R2401 B.n247 B.n246 163.367
R2402 B.n251 B.n250 163.367
R2403 B.n255 B.n254 163.367
R2404 B.n259 B.n258 163.367
R2405 B.n263 B.n262 163.367
R2406 B.n267 B.n266 163.367
R2407 B.n271 B.n270 163.367
R2408 B.n275 B.n274 163.367
R2409 B.n279 B.n278 163.367
R2410 B.n283 B.n282 163.367
R2411 B.n287 B.n286 163.367
R2412 B.n291 B.n290 163.367
R2413 B.n295 B.n294 163.367
R2414 B.n299 B.n298 163.367
R2415 B.n303 B.n302 163.367
R2416 B.n307 B.n306 163.367
R2417 B.n311 B.n310 163.367
R2418 B.n315 B.n314 163.367
R2419 B.n319 B.n318 163.367
R2420 B.n323 B.n322 163.367
R2421 B.n327 B.n326 163.367
R2422 B.n331 B.n330 163.367
R2423 B.n335 B.n334 163.367
R2424 B.n339 B.n338 163.367
R2425 B.n343 B.n342 163.367
R2426 B.n347 B.n346 163.367
R2427 B.n351 B.n350 163.367
R2428 B.n355 B.n354 163.367
R2429 B.n359 B.n358 163.367
R2430 B.n363 B.n362 163.367
R2431 B.n367 B.n366 163.367
R2432 B.n371 B.n370 163.367
R2433 B.n375 B.n374 163.367
R2434 B.n379 B.n378 163.367
R2435 B.n383 B.n382 163.367
R2436 B.n387 B.n386 163.367
R2437 B.n391 B.n390 163.367
R2438 B.n395 B.n394 163.367
R2439 B.n399 B.n398 163.367
R2440 B.n403 B.n402 163.367
R2441 B.n407 B.n406 163.367
R2442 B.n411 B.n410 163.367
R2443 B.n415 B.n414 163.367
R2444 B.n419 B.n418 163.367
R2445 B.n423 B.n422 163.367
R2446 B.n427 B.n426 163.367
R2447 B.n431 B.n430 163.367
R2448 B.n435 B.n434 163.367
R2449 B.n439 B.n438 163.367
R2450 B.n441 B.n188 163.367
R2451 B.n895 B.n894 71.676
R2452 B.n889 B.n580 71.676
R2453 B.n886 B.n581 71.676
R2454 B.n882 B.n582 71.676
R2455 B.n878 B.n583 71.676
R2456 B.n874 B.n584 71.676
R2457 B.n870 B.n585 71.676
R2458 B.n866 B.n586 71.676
R2459 B.n862 B.n587 71.676
R2460 B.n858 B.n588 71.676
R2461 B.n854 B.n589 71.676
R2462 B.n850 B.n590 71.676
R2463 B.n846 B.n591 71.676
R2464 B.n842 B.n592 71.676
R2465 B.n838 B.n593 71.676
R2466 B.n834 B.n594 71.676
R2467 B.n830 B.n595 71.676
R2468 B.n826 B.n596 71.676
R2469 B.n822 B.n597 71.676
R2470 B.n818 B.n598 71.676
R2471 B.n814 B.n599 71.676
R2472 B.n810 B.n600 71.676
R2473 B.n806 B.n601 71.676
R2474 B.n802 B.n602 71.676
R2475 B.n798 B.n603 71.676
R2476 B.n794 B.n604 71.676
R2477 B.n790 B.n605 71.676
R2478 B.n786 B.n606 71.676
R2479 B.n782 B.n607 71.676
R2480 B.n777 B.n608 71.676
R2481 B.n773 B.n609 71.676
R2482 B.n769 B.n610 71.676
R2483 B.n765 B.n611 71.676
R2484 B.n761 B.n612 71.676
R2485 B.n756 B.n613 71.676
R2486 B.n752 B.n614 71.676
R2487 B.n748 B.n615 71.676
R2488 B.n744 B.n616 71.676
R2489 B.n740 B.n617 71.676
R2490 B.n736 B.n618 71.676
R2491 B.n732 B.n619 71.676
R2492 B.n728 B.n620 71.676
R2493 B.n724 B.n621 71.676
R2494 B.n720 B.n622 71.676
R2495 B.n716 B.n623 71.676
R2496 B.n712 B.n624 71.676
R2497 B.n708 B.n625 71.676
R2498 B.n704 B.n626 71.676
R2499 B.n700 B.n627 71.676
R2500 B.n696 B.n628 71.676
R2501 B.n692 B.n629 71.676
R2502 B.n688 B.n630 71.676
R2503 B.n684 B.n631 71.676
R2504 B.n680 B.n632 71.676
R2505 B.n676 B.n633 71.676
R2506 B.n672 B.n634 71.676
R2507 B.n668 B.n635 71.676
R2508 B.n664 B.n636 71.676
R2509 B.n660 B.n637 71.676
R2510 B.n656 B.n638 71.676
R2511 B.n652 B.n639 71.676
R2512 B.n648 B.n640 71.676
R2513 B.n195 B.n126 71.676
R2514 B.n199 B.n127 71.676
R2515 B.n203 B.n128 71.676
R2516 B.n207 B.n129 71.676
R2517 B.n211 B.n130 71.676
R2518 B.n215 B.n131 71.676
R2519 B.n219 B.n132 71.676
R2520 B.n223 B.n133 71.676
R2521 B.n227 B.n134 71.676
R2522 B.n231 B.n135 71.676
R2523 B.n235 B.n136 71.676
R2524 B.n239 B.n137 71.676
R2525 B.n243 B.n138 71.676
R2526 B.n247 B.n139 71.676
R2527 B.n251 B.n140 71.676
R2528 B.n255 B.n141 71.676
R2529 B.n259 B.n142 71.676
R2530 B.n263 B.n143 71.676
R2531 B.n267 B.n144 71.676
R2532 B.n271 B.n145 71.676
R2533 B.n275 B.n146 71.676
R2534 B.n279 B.n147 71.676
R2535 B.n283 B.n148 71.676
R2536 B.n287 B.n149 71.676
R2537 B.n291 B.n150 71.676
R2538 B.n295 B.n151 71.676
R2539 B.n299 B.n152 71.676
R2540 B.n303 B.n153 71.676
R2541 B.n307 B.n154 71.676
R2542 B.n311 B.n155 71.676
R2543 B.n315 B.n156 71.676
R2544 B.n319 B.n157 71.676
R2545 B.n323 B.n158 71.676
R2546 B.n327 B.n159 71.676
R2547 B.n331 B.n160 71.676
R2548 B.n335 B.n161 71.676
R2549 B.n339 B.n162 71.676
R2550 B.n343 B.n163 71.676
R2551 B.n347 B.n164 71.676
R2552 B.n351 B.n165 71.676
R2553 B.n355 B.n166 71.676
R2554 B.n359 B.n167 71.676
R2555 B.n363 B.n168 71.676
R2556 B.n367 B.n169 71.676
R2557 B.n371 B.n170 71.676
R2558 B.n375 B.n171 71.676
R2559 B.n379 B.n172 71.676
R2560 B.n383 B.n173 71.676
R2561 B.n387 B.n174 71.676
R2562 B.n391 B.n175 71.676
R2563 B.n395 B.n176 71.676
R2564 B.n399 B.n177 71.676
R2565 B.n403 B.n178 71.676
R2566 B.n407 B.n179 71.676
R2567 B.n411 B.n180 71.676
R2568 B.n415 B.n181 71.676
R2569 B.n419 B.n182 71.676
R2570 B.n423 B.n183 71.676
R2571 B.n427 B.n184 71.676
R2572 B.n431 B.n185 71.676
R2573 B.n435 B.n186 71.676
R2574 B.n439 B.n187 71.676
R2575 B.n1196 B.n188 71.676
R2576 B.n1196 B.n1195 71.676
R2577 B.n441 B.n187 71.676
R2578 B.n438 B.n186 71.676
R2579 B.n434 B.n185 71.676
R2580 B.n430 B.n184 71.676
R2581 B.n426 B.n183 71.676
R2582 B.n422 B.n182 71.676
R2583 B.n418 B.n181 71.676
R2584 B.n414 B.n180 71.676
R2585 B.n410 B.n179 71.676
R2586 B.n406 B.n178 71.676
R2587 B.n402 B.n177 71.676
R2588 B.n398 B.n176 71.676
R2589 B.n394 B.n175 71.676
R2590 B.n390 B.n174 71.676
R2591 B.n386 B.n173 71.676
R2592 B.n382 B.n172 71.676
R2593 B.n378 B.n171 71.676
R2594 B.n374 B.n170 71.676
R2595 B.n370 B.n169 71.676
R2596 B.n366 B.n168 71.676
R2597 B.n362 B.n167 71.676
R2598 B.n358 B.n166 71.676
R2599 B.n354 B.n165 71.676
R2600 B.n350 B.n164 71.676
R2601 B.n346 B.n163 71.676
R2602 B.n342 B.n162 71.676
R2603 B.n338 B.n161 71.676
R2604 B.n334 B.n160 71.676
R2605 B.n330 B.n159 71.676
R2606 B.n326 B.n158 71.676
R2607 B.n322 B.n157 71.676
R2608 B.n318 B.n156 71.676
R2609 B.n314 B.n155 71.676
R2610 B.n310 B.n154 71.676
R2611 B.n306 B.n153 71.676
R2612 B.n302 B.n152 71.676
R2613 B.n298 B.n151 71.676
R2614 B.n294 B.n150 71.676
R2615 B.n290 B.n149 71.676
R2616 B.n286 B.n148 71.676
R2617 B.n282 B.n147 71.676
R2618 B.n278 B.n146 71.676
R2619 B.n274 B.n145 71.676
R2620 B.n270 B.n144 71.676
R2621 B.n266 B.n143 71.676
R2622 B.n262 B.n142 71.676
R2623 B.n258 B.n141 71.676
R2624 B.n254 B.n140 71.676
R2625 B.n250 B.n139 71.676
R2626 B.n246 B.n138 71.676
R2627 B.n242 B.n137 71.676
R2628 B.n238 B.n136 71.676
R2629 B.n234 B.n135 71.676
R2630 B.n230 B.n134 71.676
R2631 B.n226 B.n133 71.676
R2632 B.n222 B.n132 71.676
R2633 B.n218 B.n131 71.676
R2634 B.n214 B.n130 71.676
R2635 B.n210 B.n129 71.676
R2636 B.n206 B.n128 71.676
R2637 B.n202 B.n127 71.676
R2638 B.n198 B.n126 71.676
R2639 B.n895 B.n642 71.676
R2640 B.n887 B.n580 71.676
R2641 B.n883 B.n581 71.676
R2642 B.n879 B.n582 71.676
R2643 B.n875 B.n583 71.676
R2644 B.n871 B.n584 71.676
R2645 B.n867 B.n585 71.676
R2646 B.n863 B.n586 71.676
R2647 B.n859 B.n587 71.676
R2648 B.n855 B.n588 71.676
R2649 B.n851 B.n589 71.676
R2650 B.n847 B.n590 71.676
R2651 B.n843 B.n591 71.676
R2652 B.n839 B.n592 71.676
R2653 B.n835 B.n593 71.676
R2654 B.n831 B.n594 71.676
R2655 B.n827 B.n595 71.676
R2656 B.n823 B.n596 71.676
R2657 B.n819 B.n597 71.676
R2658 B.n815 B.n598 71.676
R2659 B.n811 B.n599 71.676
R2660 B.n807 B.n600 71.676
R2661 B.n803 B.n601 71.676
R2662 B.n799 B.n602 71.676
R2663 B.n795 B.n603 71.676
R2664 B.n791 B.n604 71.676
R2665 B.n787 B.n605 71.676
R2666 B.n783 B.n606 71.676
R2667 B.n778 B.n607 71.676
R2668 B.n774 B.n608 71.676
R2669 B.n770 B.n609 71.676
R2670 B.n766 B.n610 71.676
R2671 B.n762 B.n611 71.676
R2672 B.n757 B.n612 71.676
R2673 B.n753 B.n613 71.676
R2674 B.n749 B.n614 71.676
R2675 B.n745 B.n615 71.676
R2676 B.n741 B.n616 71.676
R2677 B.n737 B.n617 71.676
R2678 B.n733 B.n618 71.676
R2679 B.n729 B.n619 71.676
R2680 B.n725 B.n620 71.676
R2681 B.n721 B.n621 71.676
R2682 B.n717 B.n622 71.676
R2683 B.n713 B.n623 71.676
R2684 B.n709 B.n624 71.676
R2685 B.n705 B.n625 71.676
R2686 B.n701 B.n626 71.676
R2687 B.n697 B.n627 71.676
R2688 B.n693 B.n628 71.676
R2689 B.n689 B.n629 71.676
R2690 B.n685 B.n630 71.676
R2691 B.n681 B.n631 71.676
R2692 B.n677 B.n632 71.676
R2693 B.n673 B.n633 71.676
R2694 B.n669 B.n634 71.676
R2695 B.n665 B.n635 71.676
R2696 B.n661 B.n636 71.676
R2697 B.n657 B.n637 71.676
R2698 B.n653 B.n638 71.676
R2699 B.n649 B.n639 71.676
R2700 B.n640 B.n579 71.676
R2701 B.n646 B.n645 66.9096
R2702 B.n644 B.n643 66.9096
R2703 B.n193 B.n192 66.9096
R2704 B.n190 B.n189 66.9096
R2705 B.n759 B.n646 59.5399
R2706 B.n780 B.n644 59.5399
R2707 B.n194 B.n193 59.5399
R2708 B.n191 B.n190 59.5399
R2709 B.n896 B.n576 59.1998
R2710 B.n1198 B.n1197 59.1998
R2711 B.n902 B.n576 32.7286
R2712 B.n902 B.n572 32.7286
R2713 B.n908 B.n572 32.7286
R2714 B.n908 B.n568 32.7286
R2715 B.n914 B.n568 32.7286
R2716 B.n914 B.n563 32.7286
R2717 B.n920 B.n563 32.7286
R2718 B.n920 B.n564 32.7286
R2719 B.n926 B.n556 32.7286
R2720 B.n932 B.n556 32.7286
R2721 B.n932 B.n552 32.7286
R2722 B.n938 B.n552 32.7286
R2723 B.n938 B.n548 32.7286
R2724 B.n944 B.n548 32.7286
R2725 B.n944 B.n544 32.7286
R2726 B.n950 B.n544 32.7286
R2727 B.n950 B.n540 32.7286
R2728 B.n956 B.n540 32.7286
R2729 B.n956 B.n536 32.7286
R2730 B.n962 B.n536 32.7286
R2731 B.n968 B.n532 32.7286
R2732 B.n968 B.n528 32.7286
R2733 B.n974 B.n528 32.7286
R2734 B.n974 B.n524 32.7286
R2735 B.n980 B.n524 32.7286
R2736 B.n980 B.n520 32.7286
R2737 B.n986 B.n520 32.7286
R2738 B.n986 B.n516 32.7286
R2739 B.n992 B.n516 32.7286
R2740 B.n998 B.n512 32.7286
R2741 B.n998 B.n508 32.7286
R2742 B.n1004 B.n508 32.7286
R2743 B.n1004 B.n504 32.7286
R2744 B.n1010 B.n504 32.7286
R2745 B.n1010 B.n500 32.7286
R2746 B.n1016 B.n500 32.7286
R2747 B.n1016 B.n496 32.7286
R2748 B.n1023 B.n496 32.7286
R2749 B.n1023 B.n1022 32.7286
R2750 B.n1029 B.n489 32.7286
R2751 B.n1035 B.n489 32.7286
R2752 B.n1035 B.n485 32.7286
R2753 B.n1041 B.n485 32.7286
R2754 B.n1041 B.n481 32.7286
R2755 B.n1047 B.n481 32.7286
R2756 B.n1047 B.n476 32.7286
R2757 B.n1053 B.n476 32.7286
R2758 B.n1053 B.n477 32.7286
R2759 B.n1059 B.n469 32.7286
R2760 B.n1065 B.n469 32.7286
R2761 B.n1065 B.n465 32.7286
R2762 B.n1071 B.n465 32.7286
R2763 B.n1071 B.n461 32.7286
R2764 B.n1077 B.n461 32.7286
R2765 B.n1077 B.n457 32.7286
R2766 B.n1084 B.n457 32.7286
R2767 B.n1084 B.n1083 32.7286
R2768 B.n1090 B.n450 32.7286
R2769 B.n1097 B.n450 32.7286
R2770 B.n1097 B.n446 32.7286
R2771 B.n1103 B.n446 32.7286
R2772 B.n1103 B.n4 32.7286
R2773 B.n1335 B.n4 32.7286
R2774 B.n1335 B.n1334 32.7286
R2775 B.n1334 B.n1333 32.7286
R2776 B.n1333 B.n8 32.7286
R2777 B.n1327 B.n8 32.7286
R2778 B.n1327 B.n1326 32.7286
R2779 B.n1326 B.n1325 32.7286
R2780 B.n1319 B.n18 32.7286
R2781 B.n1319 B.n1318 32.7286
R2782 B.n1318 B.n1317 32.7286
R2783 B.n1317 B.n22 32.7286
R2784 B.n1311 B.n22 32.7286
R2785 B.n1311 B.n1310 32.7286
R2786 B.n1310 B.n1309 32.7286
R2787 B.n1309 B.n29 32.7286
R2788 B.n1303 B.n29 32.7286
R2789 B.n1302 B.n1301 32.7286
R2790 B.n1301 B.n36 32.7286
R2791 B.n1295 B.n36 32.7286
R2792 B.n1295 B.n1294 32.7286
R2793 B.n1294 B.n1293 32.7286
R2794 B.n1293 B.n43 32.7286
R2795 B.n1287 B.n43 32.7286
R2796 B.n1287 B.n1286 32.7286
R2797 B.n1286 B.n1285 32.7286
R2798 B.n1279 B.n53 32.7286
R2799 B.n1279 B.n1278 32.7286
R2800 B.n1278 B.n1277 32.7286
R2801 B.n1277 B.n57 32.7286
R2802 B.n1271 B.n57 32.7286
R2803 B.n1271 B.n1270 32.7286
R2804 B.n1270 B.n1269 32.7286
R2805 B.n1269 B.n64 32.7286
R2806 B.n1263 B.n64 32.7286
R2807 B.n1263 B.n1262 32.7286
R2808 B.n1261 B.n71 32.7286
R2809 B.n1255 B.n71 32.7286
R2810 B.n1255 B.n1254 32.7286
R2811 B.n1254 B.n1253 32.7286
R2812 B.n1253 B.n78 32.7286
R2813 B.n1247 B.n78 32.7286
R2814 B.n1247 B.n1246 32.7286
R2815 B.n1246 B.n1245 32.7286
R2816 B.n1245 B.n85 32.7286
R2817 B.n1239 B.n1238 32.7286
R2818 B.n1238 B.n1237 32.7286
R2819 B.n1237 B.n92 32.7286
R2820 B.n1231 B.n92 32.7286
R2821 B.n1231 B.n1230 32.7286
R2822 B.n1230 B.n1229 32.7286
R2823 B.n1229 B.n99 32.7286
R2824 B.n1223 B.n99 32.7286
R2825 B.n1223 B.n1222 32.7286
R2826 B.n1222 B.n1221 32.7286
R2827 B.n1221 B.n106 32.7286
R2828 B.n1215 B.n106 32.7286
R2829 B.n1214 B.n1213 32.7286
R2830 B.n1213 B.n113 32.7286
R2831 B.n1207 B.n113 32.7286
R2832 B.n1207 B.n1206 32.7286
R2833 B.n1206 B.n1205 32.7286
R2834 B.n1205 B.n120 32.7286
R2835 B.n1199 B.n120 32.7286
R2836 B.n1199 B.n1198 32.7286
R2837 B.n1029 B.t0 31.766
R2838 B.n1285 B.t3 31.766
R2839 B.n196 B.n122 30.4395
R2840 B.n1194 B.n1193 30.4395
R2841 B.n899 B.n898 30.4395
R2842 B.n893 B.n574 30.4395
R2843 B.n992 B.t7 28.8782
R2844 B.t4 B.n1261 28.8782
R2845 B.n1059 B.t9 26.953
R2846 B.n1303 B.t6 26.953
R2847 B.n962 B.t8 24.0653
R2848 B.n1239 B.t2 24.0653
R2849 B.n1090 B.t1 22.1401
R2850 B.n1325 B.t5 22.1401
R2851 B.n926 B.t15 20.2149
R2852 B.n1215 B.t11 20.2149
R2853 B B.n1337 18.0485
R2854 B.n564 B.t15 12.5142
R2855 B.t11 B.n1214 12.5142
R2856 B.n197 B.n196 10.6151
R2857 B.n200 B.n197 10.6151
R2858 B.n201 B.n200 10.6151
R2859 B.n204 B.n201 10.6151
R2860 B.n205 B.n204 10.6151
R2861 B.n208 B.n205 10.6151
R2862 B.n209 B.n208 10.6151
R2863 B.n212 B.n209 10.6151
R2864 B.n213 B.n212 10.6151
R2865 B.n216 B.n213 10.6151
R2866 B.n217 B.n216 10.6151
R2867 B.n220 B.n217 10.6151
R2868 B.n221 B.n220 10.6151
R2869 B.n224 B.n221 10.6151
R2870 B.n225 B.n224 10.6151
R2871 B.n228 B.n225 10.6151
R2872 B.n229 B.n228 10.6151
R2873 B.n232 B.n229 10.6151
R2874 B.n233 B.n232 10.6151
R2875 B.n236 B.n233 10.6151
R2876 B.n237 B.n236 10.6151
R2877 B.n240 B.n237 10.6151
R2878 B.n241 B.n240 10.6151
R2879 B.n244 B.n241 10.6151
R2880 B.n245 B.n244 10.6151
R2881 B.n248 B.n245 10.6151
R2882 B.n249 B.n248 10.6151
R2883 B.n252 B.n249 10.6151
R2884 B.n253 B.n252 10.6151
R2885 B.n256 B.n253 10.6151
R2886 B.n257 B.n256 10.6151
R2887 B.n260 B.n257 10.6151
R2888 B.n261 B.n260 10.6151
R2889 B.n264 B.n261 10.6151
R2890 B.n265 B.n264 10.6151
R2891 B.n268 B.n265 10.6151
R2892 B.n269 B.n268 10.6151
R2893 B.n272 B.n269 10.6151
R2894 B.n273 B.n272 10.6151
R2895 B.n276 B.n273 10.6151
R2896 B.n277 B.n276 10.6151
R2897 B.n280 B.n277 10.6151
R2898 B.n281 B.n280 10.6151
R2899 B.n284 B.n281 10.6151
R2900 B.n285 B.n284 10.6151
R2901 B.n288 B.n285 10.6151
R2902 B.n289 B.n288 10.6151
R2903 B.n292 B.n289 10.6151
R2904 B.n293 B.n292 10.6151
R2905 B.n296 B.n293 10.6151
R2906 B.n297 B.n296 10.6151
R2907 B.n300 B.n297 10.6151
R2908 B.n301 B.n300 10.6151
R2909 B.n304 B.n301 10.6151
R2910 B.n305 B.n304 10.6151
R2911 B.n308 B.n305 10.6151
R2912 B.n309 B.n308 10.6151
R2913 B.n313 B.n312 10.6151
R2914 B.n316 B.n313 10.6151
R2915 B.n317 B.n316 10.6151
R2916 B.n320 B.n317 10.6151
R2917 B.n321 B.n320 10.6151
R2918 B.n324 B.n321 10.6151
R2919 B.n325 B.n324 10.6151
R2920 B.n328 B.n325 10.6151
R2921 B.n329 B.n328 10.6151
R2922 B.n333 B.n332 10.6151
R2923 B.n336 B.n333 10.6151
R2924 B.n337 B.n336 10.6151
R2925 B.n340 B.n337 10.6151
R2926 B.n341 B.n340 10.6151
R2927 B.n344 B.n341 10.6151
R2928 B.n345 B.n344 10.6151
R2929 B.n348 B.n345 10.6151
R2930 B.n349 B.n348 10.6151
R2931 B.n352 B.n349 10.6151
R2932 B.n353 B.n352 10.6151
R2933 B.n356 B.n353 10.6151
R2934 B.n357 B.n356 10.6151
R2935 B.n360 B.n357 10.6151
R2936 B.n361 B.n360 10.6151
R2937 B.n364 B.n361 10.6151
R2938 B.n365 B.n364 10.6151
R2939 B.n368 B.n365 10.6151
R2940 B.n369 B.n368 10.6151
R2941 B.n372 B.n369 10.6151
R2942 B.n373 B.n372 10.6151
R2943 B.n376 B.n373 10.6151
R2944 B.n377 B.n376 10.6151
R2945 B.n380 B.n377 10.6151
R2946 B.n381 B.n380 10.6151
R2947 B.n384 B.n381 10.6151
R2948 B.n385 B.n384 10.6151
R2949 B.n388 B.n385 10.6151
R2950 B.n389 B.n388 10.6151
R2951 B.n392 B.n389 10.6151
R2952 B.n393 B.n392 10.6151
R2953 B.n396 B.n393 10.6151
R2954 B.n397 B.n396 10.6151
R2955 B.n400 B.n397 10.6151
R2956 B.n401 B.n400 10.6151
R2957 B.n404 B.n401 10.6151
R2958 B.n405 B.n404 10.6151
R2959 B.n408 B.n405 10.6151
R2960 B.n409 B.n408 10.6151
R2961 B.n412 B.n409 10.6151
R2962 B.n413 B.n412 10.6151
R2963 B.n416 B.n413 10.6151
R2964 B.n417 B.n416 10.6151
R2965 B.n420 B.n417 10.6151
R2966 B.n421 B.n420 10.6151
R2967 B.n424 B.n421 10.6151
R2968 B.n425 B.n424 10.6151
R2969 B.n428 B.n425 10.6151
R2970 B.n429 B.n428 10.6151
R2971 B.n432 B.n429 10.6151
R2972 B.n433 B.n432 10.6151
R2973 B.n436 B.n433 10.6151
R2974 B.n437 B.n436 10.6151
R2975 B.n440 B.n437 10.6151
R2976 B.n442 B.n440 10.6151
R2977 B.n443 B.n442 10.6151
R2978 B.n1194 B.n443 10.6151
R2979 B.n900 B.n899 10.6151
R2980 B.n900 B.n570 10.6151
R2981 B.n910 B.n570 10.6151
R2982 B.n911 B.n910 10.6151
R2983 B.n912 B.n911 10.6151
R2984 B.n912 B.n561 10.6151
R2985 B.n922 B.n561 10.6151
R2986 B.n923 B.n922 10.6151
R2987 B.n924 B.n923 10.6151
R2988 B.n924 B.n554 10.6151
R2989 B.n934 B.n554 10.6151
R2990 B.n935 B.n934 10.6151
R2991 B.n936 B.n935 10.6151
R2992 B.n936 B.n546 10.6151
R2993 B.n946 B.n546 10.6151
R2994 B.n947 B.n946 10.6151
R2995 B.n948 B.n947 10.6151
R2996 B.n948 B.n538 10.6151
R2997 B.n958 B.n538 10.6151
R2998 B.n959 B.n958 10.6151
R2999 B.n960 B.n959 10.6151
R3000 B.n960 B.n530 10.6151
R3001 B.n970 B.n530 10.6151
R3002 B.n971 B.n970 10.6151
R3003 B.n972 B.n971 10.6151
R3004 B.n972 B.n522 10.6151
R3005 B.n982 B.n522 10.6151
R3006 B.n983 B.n982 10.6151
R3007 B.n984 B.n983 10.6151
R3008 B.n984 B.n514 10.6151
R3009 B.n994 B.n514 10.6151
R3010 B.n995 B.n994 10.6151
R3011 B.n996 B.n995 10.6151
R3012 B.n996 B.n506 10.6151
R3013 B.n1006 B.n506 10.6151
R3014 B.n1007 B.n1006 10.6151
R3015 B.n1008 B.n1007 10.6151
R3016 B.n1008 B.n498 10.6151
R3017 B.n1018 B.n498 10.6151
R3018 B.n1019 B.n1018 10.6151
R3019 B.n1020 B.n1019 10.6151
R3020 B.n1020 B.n491 10.6151
R3021 B.n1031 B.n491 10.6151
R3022 B.n1032 B.n1031 10.6151
R3023 B.n1033 B.n1032 10.6151
R3024 B.n1033 B.n483 10.6151
R3025 B.n1043 B.n483 10.6151
R3026 B.n1044 B.n1043 10.6151
R3027 B.n1045 B.n1044 10.6151
R3028 B.n1045 B.n474 10.6151
R3029 B.n1055 B.n474 10.6151
R3030 B.n1056 B.n1055 10.6151
R3031 B.n1057 B.n1056 10.6151
R3032 B.n1057 B.n467 10.6151
R3033 B.n1067 B.n467 10.6151
R3034 B.n1068 B.n1067 10.6151
R3035 B.n1069 B.n1068 10.6151
R3036 B.n1069 B.n459 10.6151
R3037 B.n1079 B.n459 10.6151
R3038 B.n1080 B.n1079 10.6151
R3039 B.n1081 B.n1080 10.6151
R3040 B.n1081 B.n452 10.6151
R3041 B.n1092 B.n452 10.6151
R3042 B.n1093 B.n1092 10.6151
R3043 B.n1095 B.n1093 10.6151
R3044 B.n1095 B.n1094 10.6151
R3045 B.n1094 B.n444 10.6151
R3046 B.n1106 B.n444 10.6151
R3047 B.n1107 B.n1106 10.6151
R3048 B.n1108 B.n1107 10.6151
R3049 B.n1109 B.n1108 10.6151
R3050 B.n1111 B.n1109 10.6151
R3051 B.n1112 B.n1111 10.6151
R3052 B.n1113 B.n1112 10.6151
R3053 B.n1114 B.n1113 10.6151
R3054 B.n1116 B.n1114 10.6151
R3055 B.n1117 B.n1116 10.6151
R3056 B.n1118 B.n1117 10.6151
R3057 B.n1119 B.n1118 10.6151
R3058 B.n1121 B.n1119 10.6151
R3059 B.n1122 B.n1121 10.6151
R3060 B.n1123 B.n1122 10.6151
R3061 B.n1124 B.n1123 10.6151
R3062 B.n1126 B.n1124 10.6151
R3063 B.n1127 B.n1126 10.6151
R3064 B.n1128 B.n1127 10.6151
R3065 B.n1129 B.n1128 10.6151
R3066 B.n1131 B.n1129 10.6151
R3067 B.n1132 B.n1131 10.6151
R3068 B.n1133 B.n1132 10.6151
R3069 B.n1134 B.n1133 10.6151
R3070 B.n1136 B.n1134 10.6151
R3071 B.n1137 B.n1136 10.6151
R3072 B.n1138 B.n1137 10.6151
R3073 B.n1139 B.n1138 10.6151
R3074 B.n1141 B.n1139 10.6151
R3075 B.n1142 B.n1141 10.6151
R3076 B.n1143 B.n1142 10.6151
R3077 B.n1144 B.n1143 10.6151
R3078 B.n1146 B.n1144 10.6151
R3079 B.n1147 B.n1146 10.6151
R3080 B.n1148 B.n1147 10.6151
R3081 B.n1149 B.n1148 10.6151
R3082 B.n1151 B.n1149 10.6151
R3083 B.n1152 B.n1151 10.6151
R3084 B.n1153 B.n1152 10.6151
R3085 B.n1154 B.n1153 10.6151
R3086 B.n1156 B.n1154 10.6151
R3087 B.n1157 B.n1156 10.6151
R3088 B.n1158 B.n1157 10.6151
R3089 B.n1159 B.n1158 10.6151
R3090 B.n1161 B.n1159 10.6151
R3091 B.n1162 B.n1161 10.6151
R3092 B.n1163 B.n1162 10.6151
R3093 B.n1164 B.n1163 10.6151
R3094 B.n1166 B.n1164 10.6151
R3095 B.n1167 B.n1166 10.6151
R3096 B.n1168 B.n1167 10.6151
R3097 B.n1169 B.n1168 10.6151
R3098 B.n1171 B.n1169 10.6151
R3099 B.n1172 B.n1171 10.6151
R3100 B.n1173 B.n1172 10.6151
R3101 B.n1174 B.n1173 10.6151
R3102 B.n1176 B.n1174 10.6151
R3103 B.n1177 B.n1176 10.6151
R3104 B.n1178 B.n1177 10.6151
R3105 B.n1179 B.n1178 10.6151
R3106 B.n1181 B.n1179 10.6151
R3107 B.n1182 B.n1181 10.6151
R3108 B.n1183 B.n1182 10.6151
R3109 B.n1184 B.n1183 10.6151
R3110 B.n1186 B.n1184 10.6151
R3111 B.n1187 B.n1186 10.6151
R3112 B.n1188 B.n1187 10.6151
R3113 B.n1189 B.n1188 10.6151
R3114 B.n1191 B.n1189 10.6151
R3115 B.n1192 B.n1191 10.6151
R3116 B.n1193 B.n1192 10.6151
R3117 B.n893 B.n892 10.6151
R3118 B.n892 B.n891 10.6151
R3119 B.n891 B.n890 10.6151
R3120 B.n890 B.n888 10.6151
R3121 B.n888 B.n885 10.6151
R3122 B.n885 B.n884 10.6151
R3123 B.n884 B.n881 10.6151
R3124 B.n881 B.n880 10.6151
R3125 B.n880 B.n877 10.6151
R3126 B.n877 B.n876 10.6151
R3127 B.n876 B.n873 10.6151
R3128 B.n873 B.n872 10.6151
R3129 B.n872 B.n869 10.6151
R3130 B.n869 B.n868 10.6151
R3131 B.n868 B.n865 10.6151
R3132 B.n865 B.n864 10.6151
R3133 B.n864 B.n861 10.6151
R3134 B.n861 B.n860 10.6151
R3135 B.n860 B.n857 10.6151
R3136 B.n857 B.n856 10.6151
R3137 B.n856 B.n853 10.6151
R3138 B.n853 B.n852 10.6151
R3139 B.n852 B.n849 10.6151
R3140 B.n849 B.n848 10.6151
R3141 B.n848 B.n845 10.6151
R3142 B.n845 B.n844 10.6151
R3143 B.n844 B.n841 10.6151
R3144 B.n841 B.n840 10.6151
R3145 B.n840 B.n837 10.6151
R3146 B.n837 B.n836 10.6151
R3147 B.n836 B.n833 10.6151
R3148 B.n833 B.n832 10.6151
R3149 B.n832 B.n829 10.6151
R3150 B.n829 B.n828 10.6151
R3151 B.n828 B.n825 10.6151
R3152 B.n825 B.n824 10.6151
R3153 B.n824 B.n821 10.6151
R3154 B.n821 B.n820 10.6151
R3155 B.n820 B.n817 10.6151
R3156 B.n817 B.n816 10.6151
R3157 B.n816 B.n813 10.6151
R3158 B.n813 B.n812 10.6151
R3159 B.n812 B.n809 10.6151
R3160 B.n809 B.n808 10.6151
R3161 B.n808 B.n805 10.6151
R3162 B.n805 B.n804 10.6151
R3163 B.n804 B.n801 10.6151
R3164 B.n801 B.n800 10.6151
R3165 B.n800 B.n797 10.6151
R3166 B.n797 B.n796 10.6151
R3167 B.n796 B.n793 10.6151
R3168 B.n793 B.n792 10.6151
R3169 B.n792 B.n789 10.6151
R3170 B.n789 B.n788 10.6151
R3171 B.n788 B.n785 10.6151
R3172 B.n785 B.n784 10.6151
R3173 B.n784 B.n781 10.6151
R3174 B.n779 B.n776 10.6151
R3175 B.n776 B.n775 10.6151
R3176 B.n775 B.n772 10.6151
R3177 B.n772 B.n771 10.6151
R3178 B.n771 B.n768 10.6151
R3179 B.n768 B.n767 10.6151
R3180 B.n767 B.n764 10.6151
R3181 B.n764 B.n763 10.6151
R3182 B.n763 B.n760 10.6151
R3183 B.n758 B.n755 10.6151
R3184 B.n755 B.n754 10.6151
R3185 B.n754 B.n751 10.6151
R3186 B.n751 B.n750 10.6151
R3187 B.n750 B.n747 10.6151
R3188 B.n747 B.n746 10.6151
R3189 B.n746 B.n743 10.6151
R3190 B.n743 B.n742 10.6151
R3191 B.n742 B.n739 10.6151
R3192 B.n739 B.n738 10.6151
R3193 B.n738 B.n735 10.6151
R3194 B.n735 B.n734 10.6151
R3195 B.n734 B.n731 10.6151
R3196 B.n731 B.n730 10.6151
R3197 B.n730 B.n727 10.6151
R3198 B.n727 B.n726 10.6151
R3199 B.n726 B.n723 10.6151
R3200 B.n723 B.n722 10.6151
R3201 B.n722 B.n719 10.6151
R3202 B.n719 B.n718 10.6151
R3203 B.n718 B.n715 10.6151
R3204 B.n715 B.n714 10.6151
R3205 B.n714 B.n711 10.6151
R3206 B.n711 B.n710 10.6151
R3207 B.n710 B.n707 10.6151
R3208 B.n707 B.n706 10.6151
R3209 B.n706 B.n703 10.6151
R3210 B.n703 B.n702 10.6151
R3211 B.n702 B.n699 10.6151
R3212 B.n699 B.n698 10.6151
R3213 B.n698 B.n695 10.6151
R3214 B.n695 B.n694 10.6151
R3215 B.n694 B.n691 10.6151
R3216 B.n691 B.n690 10.6151
R3217 B.n690 B.n687 10.6151
R3218 B.n687 B.n686 10.6151
R3219 B.n686 B.n683 10.6151
R3220 B.n683 B.n682 10.6151
R3221 B.n682 B.n679 10.6151
R3222 B.n679 B.n678 10.6151
R3223 B.n678 B.n675 10.6151
R3224 B.n675 B.n674 10.6151
R3225 B.n674 B.n671 10.6151
R3226 B.n671 B.n670 10.6151
R3227 B.n670 B.n667 10.6151
R3228 B.n667 B.n666 10.6151
R3229 B.n666 B.n663 10.6151
R3230 B.n663 B.n662 10.6151
R3231 B.n662 B.n659 10.6151
R3232 B.n659 B.n658 10.6151
R3233 B.n658 B.n655 10.6151
R3234 B.n655 B.n654 10.6151
R3235 B.n654 B.n651 10.6151
R3236 B.n651 B.n650 10.6151
R3237 B.n650 B.n647 10.6151
R3238 B.n647 B.n578 10.6151
R3239 B.n898 B.n578 10.6151
R3240 B.n904 B.n574 10.6151
R3241 B.n905 B.n904 10.6151
R3242 B.n906 B.n905 10.6151
R3243 B.n906 B.n566 10.6151
R3244 B.n916 B.n566 10.6151
R3245 B.n917 B.n916 10.6151
R3246 B.n918 B.n917 10.6151
R3247 B.n918 B.n558 10.6151
R3248 B.n928 B.n558 10.6151
R3249 B.n929 B.n928 10.6151
R3250 B.n930 B.n929 10.6151
R3251 B.n930 B.n550 10.6151
R3252 B.n940 B.n550 10.6151
R3253 B.n941 B.n940 10.6151
R3254 B.n942 B.n941 10.6151
R3255 B.n942 B.n542 10.6151
R3256 B.n952 B.n542 10.6151
R3257 B.n953 B.n952 10.6151
R3258 B.n954 B.n953 10.6151
R3259 B.n954 B.n534 10.6151
R3260 B.n964 B.n534 10.6151
R3261 B.n965 B.n964 10.6151
R3262 B.n966 B.n965 10.6151
R3263 B.n966 B.n526 10.6151
R3264 B.n976 B.n526 10.6151
R3265 B.n977 B.n976 10.6151
R3266 B.n978 B.n977 10.6151
R3267 B.n978 B.n518 10.6151
R3268 B.n988 B.n518 10.6151
R3269 B.n989 B.n988 10.6151
R3270 B.n990 B.n989 10.6151
R3271 B.n990 B.n510 10.6151
R3272 B.n1000 B.n510 10.6151
R3273 B.n1001 B.n1000 10.6151
R3274 B.n1002 B.n1001 10.6151
R3275 B.n1002 B.n502 10.6151
R3276 B.n1012 B.n502 10.6151
R3277 B.n1013 B.n1012 10.6151
R3278 B.n1014 B.n1013 10.6151
R3279 B.n1014 B.n494 10.6151
R3280 B.n1025 B.n494 10.6151
R3281 B.n1026 B.n1025 10.6151
R3282 B.n1027 B.n1026 10.6151
R3283 B.n1027 B.n487 10.6151
R3284 B.n1037 B.n487 10.6151
R3285 B.n1038 B.n1037 10.6151
R3286 B.n1039 B.n1038 10.6151
R3287 B.n1039 B.n479 10.6151
R3288 B.n1049 B.n479 10.6151
R3289 B.n1050 B.n1049 10.6151
R3290 B.n1051 B.n1050 10.6151
R3291 B.n1051 B.n471 10.6151
R3292 B.n1061 B.n471 10.6151
R3293 B.n1062 B.n1061 10.6151
R3294 B.n1063 B.n1062 10.6151
R3295 B.n1063 B.n463 10.6151
R3296 B.n1073 B.n463 10.6151
R3297 B.n1074 B.n1073 10.6151
R3298 B.n1075 B.n1074 10.6151
R3299 B.n1075 B.n455 10.6151
R3300 B.n1086 B.n455 10.6151
R3301 B.n1087 B.n1086 10.6151
R3302 B.n1088 B.n1087 10.6151
R3303 B.n1088 B.n448 10.6151
R3304 B.n1099 B.n448 10.6151
R3305 B.n1100 B.n1099 10.6151
R3306 B.n1101 B.n1100 10.6151
R3307 B.n1101 B.n0 10.6151
R3308 B.n1331 B.n1 10.6151
R3309 B.n1331 B.n1330 10.6151
R3310 B.n1330 B.n1329 10.6151
R3311 B.n1329 B.n10 10.6151
R3312 B.n1323 B.n10 10.6151
R3313 B.n1323 B.n1322 10.6151
R3314 B.n1322 B.n1321 10.6151
R3315 B.n1321 B.n16 10.6151
R3316 B.n1315 B.n16 10.6151
R3317 B.n1315 B.n1314 10.6151
R3318 B.n1314 B.n1313 10.6151
R3319 B.n1313 B.n24 10.6151
R3320 B.n1307 B.n24 10.6151
R3321 B.n1307 B.n1306 10.6151
R3322 B.n1306 B.n1305 10.6151
R3323 B.n1305 B.n31 10.6151
R3324 B.n1299 B.n31 10.6151
R3325 B.n1299 B.n1298 10.6151
R3326 B.n1298 B.n1297 10.6151
R3327 B.n1297 B.n38 10.6151
R3328 B.n1291 B.n38 10.6151
R3329 B.n1291 B.n1290 10.6151
R3330 B.n1290 B.n1289 10.6151
R3331 B.n1289 B.n45 10.6151
R3332 B.n1283 B.n45 10.6151
R3333 B.n1283 B.n1282 10.6151
R3334 B.n1282 B.n1281 10.6151
R3335 B.n1281 B.n51 10.6151
R3336 B.n1275 B.n51 10.6151
R3337 B.n1275 B.n1274 10.6151
R3338 B.n1274 B.n1273 10.6151
R3339 B.n1273 B.n59 10.6151
R3340 B.n1267 B.n59 10.6151
R3341 B.n1267 B.n1266 10.6151
R3342 B.n1266 B.n1265 10.6151
R3343 B.n1265 B.n66 10.6151
R3344 B.n1259 B.n66 10.6151
R3345 B.n1259 B.n1258 10.6151
R3346 B.n1258 B.n1257 10.6151
R3347 B.n1257 B.n73 10.6151
R3348 B.n1251 B.n73 10.6151
R3349 B.n1251 B.n1250 10.6151
R3350 B.n1250 B.n1249 10.6151
R3351 B.n1249 B.n80 10.6151
R3352 B.n1243 B.n80 10.6151
R3353 B.n1243 B.n1242 10.6151
R3354 B.n1242 B.n1241 10.6151
R3355 B.n1241 B.n87 10.6151
R3356 B.n1235 B.n87 10.6151
R3357 B.n1235 B.n1234 10.6151
R3358 B.n1234 B.n1233 10.6151
R3359 B.n1233 B.n94 10.6151
R3360 B.n1227 B.n94 10.6151
R3361 B.n1227 B.n1226 10.6151
R3362 B.n1226 B.n1225 10.6151
R3363 B.n1225 B.n101 10.6151
R3364 B.n1219 B.n101 10.6151
R3365 B.n1219 B.n1218 10.6151
R3366 B.n1218 B.n1217 10.6151
R3367 B.n1217 B.n108 10.6151
R3368 B.n1211 B.n108 10.6151
R3369 B.n1211 B.n1210 10.6151
R3370 B.n1210 B.n1209 10.6151
R3371 B.n1209 B.n115 10.6151
R3372 B.n1203 B.n115 10.6151
R3373 B.n1203 B.n1202 10.6151
R3374 B.n1202 B.n1201 10.6151
R3375 B.n1201 B.n122 10.6151
R3376 B.n1083 B.t1 10.589
R3377 B.n18 B.t5 10.589
R3378 B.n309 B.n194 9.36635
R3379 B.n332 B.n191 9.36635
R3380 B.n781 B.n780 9.36635
R3381 B.n759 B.n758 9.36635
R3382 B.t8 B.n532 8.66381
R3383 B.t2 B.n85 8.66381
R3384 B.n477 B.t9 5.77604
R3385 B.t6 B.n1302 5.77604
R3386 B.t7 B.n512 3.85086
R3387 B.n1262 B.t4 3.85086
R3388 B.n1337 B.n0 2.81026
R3389 B.n1337 B.n1 2.81026
R3390 B.n312 B.n194 1.24928
R3391 B.n329 B.n191 1.24928
R3392 B.n780 B.n779 1.24928
R3393 B.n760 B.n759 1.24928
R3394 B.n1022 B.t0 0.96309
R3395 B.n53 B.t3 0.96309
R3396 VN.n56 VN.t6 169.263
R3397 VN.n11 VN.t3 169.263
R3398 VN.n88 VN.n87 161.3
R3399 VN.n86 VN.n46 161.3
R3400 VN.n85 VN.n84 161.3
R3401 VN.n83 VN.n47 161.3
R3402 VN.n82 VN.n81 161.3
R3403 VN.n80 VN.n48 161.3
R3404 VN.n79 VN.n78 161.3
R3405 VN.n77 VN.n76 161.3
R3406 VN.n75 VN.n50 161.3
R3407 VN.n74 VN.n73 161.3
R3408 VN.n72 VN.n51 161.3
R3409 VN.n71 VN.n70 161.3
R3410 VN.n69 VN.n52 161.3
R3411 VN.n68 VN.n67 161.3
R3412 VN.n66 VN.n53 161.3
R3413 VN.n65 VN.n64 161.3
R3414 VN.n63 VN.n54 161.3
R3415 VN.n62 VN.n61 161.3
R3416 VN.n60 VN.n55 161.3
R3417 VN.n59 VN.n58 161.3
R3418 VN.n43 VN.n42 161.3
R3419 VN.n41 VN.n1 161.3
R3420 VN.n40 VN.n39 161.3
R3421 VN.n38 VN.n2 161.3
R3422 VN.n37 VN.n36 161.3
R3423 VN.n35 VN.n3 161.3
R3424 VN.n34 VN.n33 161.3
R3425 VN.n32 VN.n31 161.3
R3426 VN.n30 VN.n5 161.3
R3427 VN.n29 VN.n28 161.3
R3428 VN.n27 VN.n6 161.3
R3429 VN.n26 VN.n25 161.3
R3430 VN.n24 VN.n7 161.3
R3431 VN.n23 VN.n22 161.3
R3432 VN.n21 VN.n8 161.3
R3433 VN.n20 VN.n19 161.3
R3434 VN.n18 VN.n9 161.3
R3435 VN.n17 VN.n16 161.3
R3436 VN.n15 VN.n10 161.3
R3437 VN.n14 VN.n13 161.3
R3438 VN.n23 VN.t4 135.794
R3439 VN.n12 VN.t9 135.794
R3440 VN.n4 VN.t1 135.794
R3441 VN.n0 VN.t5 135.794
R3442 VN.n68 VN.t0 135.794
R3443 VN.n57 VN.t7 135.794
R3444 VN.n49 VN.t8 135.794
R3445 VN.n45 VN.t2 135.794
R3446 VN.n44 VN.n0 70.5721
R3447 VN.n89 VN.n45 70.5721
R3448 VN VN.n89 60.4792
R3449 VN.n18 VN.n17 56.5617
R3450 VN.n29 VN.n6 56.5617
R3451 VN.n40 VN.n2 56.5617
R3452 VN.n63 VN.n62 56.5617
R3453 VN.n74 VN.n51 56.5617
R3454 VN.n85 VN.n47 56.5617
R3455 VN.n12 VN.n11 51.9472
R3456 VN.n57 VN.n56 51.9472
R3457 VN.n13 VN.n10 24.5923
R3458 VN.n17 VN.n10 24.5923
R3459 VN.n19 VN.n18 24.5923
R3460 VN.n19 VN.n8 24.5923
R3461 VN.n23 VN.n8 24.5923
R3462 VN.n24 VN.n23 24.5923
R3463 VN.n25 VN.n24 24.5923
R3464 VN.n25 VN.n6 24.5923
R3465 VN.n30 VN.n29 24.5923
R3466 VN.n31 VN.n30 24.5923
R3467 VN.n35 VN.n34 24.5923
R3468 VN.n36 VN.n35 24.5923
R3469 VN.n36 VN.n2 24.5923
R3470 VN.n41 VN.n40 24.5923
R3471 VN.n42 VN.n41 24.5923
R3472 VN.n62 VN.n55 24.5923
R3473 VN.n58 VN.n55 24.5923
R3474 VN.n70 VN.n51 24.5923
R3475 VN.n70 VN.n69 24.5923
R3476 VN.n69 VN.n68 24.5923
R3477 VN.n68 VN.n53 24.5923
R3478 VN.n64 VN.n53 24.5923
R3479 VN.n64 VN.n63 24.5923
R3480 VN.n81 VN.n47 24.5923
R3481 VN.n81 VN.n80 24.5923
R3482 VN.n80 VN.n79 24.5923
R3483 VN.n76 VN.n75 24.5923
R3484 VN.n75 VN.n74 24.5923
R3485 VN.n87 VN.n86 24.5923
R3486 VN.n86 VN.n85 24.5923
R3487 VN.n13 VN.n12 22.1332
R3488 VN.n31 VN.n4 22.1332
R3489 VN.n58 VN.n57 22.1332
R3490 VN.n76 VN.n49 22.1332
R3491 VN.n42 VN.n0 19.674
R3492 VN.n87 VN.n45 19.674
R3493 VN.n59 VN.n56 3.92042
R3494 VN.n14 VN.n11 3.92042
R3495 VN.n34 VN.n4 2.45968
R3496 VN.n79 VN.n49 2.45968
R3497 VN.n89 VN.n88 0.354861
R3498 VN.n44 VN.n43 0.354861
R3499 VN VN.n44 0.267071
R3500 VN.n88 VN.n46 0.189894
R3501 VN.n84 VN.n46 0.189894
R3502 VN.n84 VN.n83 0.189894
R3503 VN.n83 VN.n82 0.189894
R3504 VN.n82 VN.n48 0.189894
R3505 VN.n78 VN.n48 0.189894
R3506 VN.n78 VN.n77 0.189894
R3507 VN.n77 VN.n50 0.189894
R3508 VN.n73 VN.n50 0.189894
R3509 VN.n73 VN.n72 0.189894
R3510 VN.n72 VN.n71 0.189894
R3511 VN.n71 VN.n52 0.189894
R3512 VN.n67 VN.n52 0.189894
R3513 VN.n67 VN.n66 0.189894
R3514 VN.n66 VN.n65 0.189894
R3515 VN.n65 VN.n54 0.189894
R3516 VN.n61 VN.n54 0.189894
R3517 VN.n61 VN.n60 0.189894
R3518 VN.n60 VN.n59 0.189894
R3519 VN.n15 VN.n14 0.189894
R3520 VN.n16 VN.n15 0.189894
R3521 VN.n16 VN.n9 0.189894
R3522 VN.n20 VN.n9 0.189894
R3523 VN.n21 VN.n20 0.189894
R3524 VN.n22 VN.n21 0.189894
R3525 VN.n22 VN.n7 0.189894
R3526 VN.n26 VN.n7 0.189894
R3527 VN.n27 VN.n26 0.189894
R3528 VN.n28 VN.n27 0.189894
R3529 VN.n28 VN.n5 0.189894
R3530 VN.n32 VN.n5 0.189894
R3531 VN.n33 VN.n32 0.189894
R3532 VN.n33 VN.n3 0.189894
R3533 VN.n37 VN.n3 0.189894
R3534 VN.n38 VN.n37 0.189894
R3535 VN.n39 VN.n38 0.189894
R3536 VN.n39 VN.n1 0.189894
R3537 VN.n43 VN.n1 0.189894
R3538 VDD2.n193 VDD2.n101 289.615
R3539 VDD2.n92 VDD2.n0 289.615
R3540 VDD2.n194 VDD2.n193 185
R3541 VDD2.n192 VDD2.n191 185
R3542 VDD2.n105 VDD2.n104 185
R3543 VDD2.n186 VDD2.n185 185
R3544 VDD2.n184 VDD2.n183 185
R3545 VDD2.n109 VDD2.n108 185
R3546 VDD2.n113 VDD2.n111 185
R3547 VDD2.n178 VDD2.n177 185
R3548 VDD2.n176 VDD2.n175 185
R3549 VDD2.n115 VDD2.n114 185
R3550 VDD2.n170 VDD2.n169 185
R3551 VDD2.n168 VDD2.n167 185
R3552 VDD2.n119 VDD2.n118 185
R3553 VDD2.n162 VDD2.n161 185
R3554 VDD2.n160 VDD2.n159 185
R3555 VDD2.n123 VDD2.n122 185
R3556 VDD2.n154 VDD2.n153 185
R3557 VDD2.n152 VDD2.n151 185
R3558 VDD2.n127 VDD2.n126 185
R3559 VDD2.n146 VDD2.n145 185
R3560 VDD2.n144 VDD2.n143 185
R3561 VDD2.n131 VDD2.n130 185
R3562 VDD2.n138 VDD2.n137 185
R3563 VDD2.n136 VDD2.n135 185
R3564 VDD2.n33 VDD2.n32 185
R3565 VDD2.n35 VDD2.n34 185
R3566 VDD2.n28 VDD2.n27 185
R3567 VDD2.n41 VDD2.n40 185
R3568 VDD2.n43 VDD2.n42 185
R3569 VDD2.n24 VDD2.n23 185
R3570 VDD2.n49 VDD2.n48 185
R3571 VDD2.n51 VDD2.n50 185
R3572 VDD2.n20 VDD2.n19 185
R3573 VDD2.n57 VDD2.n56 185
R3574 VDD2.n59 VDD2.n58 185
R3575 VDD2.n16 VDD2.n15 185
R3576 VDD2.n65 VDD2.n64 185
R3577 VDD2.n67 VDD2.n66 185
R3578 VDD2.n12 VDD2.n11 185
R3579 VDD2.n74 VDD2.n73 185
R3580 VDD2.n75 VDD2.n10 185
R3581 VDD2.n77 VDD2.n76 185
R3582 VDD2.n8 VDD2.n7 185
R3583 VDD2.n83 VDD2.n82 185
R3584 VDD2.n85 VDD2.n84 185
R3585 VDD2.n4 VDD2.n3 185
R3586 VDD2.n91 VDD2.n90 185
R3587 VDD2.n93 VDD2.n92 185
R3588 VDD2.n134 VDD2.t7 147.659
R3589 VDD2.n31 VDD2.t6 147.659
R3590 VDD2.n193 VDD2.n192 104.615
R3591 VDD2.n192 VDD2.n104 104.615
R3592 VDD2.n185 VDD2.n104 104.615
R3593 VDD2.n185 VDD2.n184 104.615
R3594 VDD2.n184 VDD2.n108 104.615
R3595 VDD2.n113 VDD2.n108 104.615
R3596 VDD2.n177 VDD2.n113 104.615
R3597 VDD2.n177 VDD2.n176 104.615
R3598 VDD2.n176 VDD2.n114 104.615
R3599 VDD2.n169 VDD2.n114 104.615
R3600 VDD2.n169 VDD2.n168 104.615
R3601 VDD2.n168 VDD2.n118 104.615
R3602 VDD2.n161 VDD2.n118 104.615
R3603 VDD2.n161 VDD2.n160 104.615
R3604 VDD2.n160 VDD2.n122 104.615
R3605 VDD2.n153 VDD2.n122 104.615
R3606 VDD2.n153 VDD2.n152 104.615
R3607 VDD2.n152 VDD2.n126 104.615
R3608 VDD2.n145 VDD2.n126 104.615
R3609 VDD2.n145 VDD2.n144 104.615
R3610 VDD2.n144 VDD2.n130 104.615
R3611 VDD2.n137 VDD2.n130 104.615
R3612 VDD2.n137 VDD2.n136 104.615
R3613 VDD2.n34 VDD2.n33 104.615
R3614 VDD2.n34 VDD2.n27 104.615
R3615 VDD2.n41 VDD2.n27 104.615
R3616 VDD2.n42 VDD2.n41 104.615
R3617 VDD2.n42 VDD2.n23 104.615
R3618 VDD2.n49 VDD2.n23 104.615
R3619 VDD2.n50 VDD2.n49 104.615
R3620 VDD2.n50 VDD2.n19 104.615
R3621 VDD2.n57 VDD2.n19 104.615
R3622 VDD2.n58 VDD2.n57 104.615
R3623 VDD2.n58 VDD2.n15 104.615
R3624 VDD2.n65 VDD2.n15 104.615
R3625 VDD2.n66 VDD2.n65 104.615
R3626 VDD2.n66 VDD2.n11 104.615
R3627 VDD2.n74 VDD2.n11 104.615
R3628 VDD2.n75 VDD2.n74 104.615
R3629 VDD2.n76 VDD2.n75 104.615
R3630 VDD2.n76 VDD2.n7 104.615
R3631 VDD2.n83 VDD2.n7 104.615
R3632 VDD2.n84 VDD2.n83 104.615
R3633 VDD2.n84 VDD2.n3 104.615
R3634 VDD2.n91 VDD2.n3 104.615
R3635 VDD2.n92 VDD2.n91 104.615
R3636 VDD2.n100 VDD2.n99 64.0209
R3637 VDD2 VDD2.n201 64.018
R3638 VDD2.n200 VDD2.n199 61.8458
R3639 VDD2.n98 VDD2.n97 61.8456
R3640 VDD2.n98 VDD2.n96 53.0019
R3641 VDD2.n198 VDD2.n100 52.9976
R3642 VDD2.n136 VDD2.t7 52.3082
R3643 VDD2.n33 VDD2.t6 52.3082
R3644 VDD2.n198 VDD2.n197 50.0278
R3645 VDD2.n135 VDD2.n134 15.6677
R3646 VDD2.n32 VDD2.n31 15.6677
R3647 VDD2.n111 VDD2.n109 13.1884
R3648 VDD2.n77 VDD2.n8 13.1884
R3649 VDD2.n183 VDD2.n182 12.8005
R3650 VDD2.n179 VDD2.n178 12.8005
R3651 VDD2.n138 VDD2.n133 12.8005
R3652 VDD2.n35 VDD2.n30 12.8005
R3653 VDD2.n78 VDD2.n10 12.8005
R3654 VDD2.n82 VDD2.n81 12.8005
R3655 VDD2.n186 VDD2.n107 12.0247
R3656 VDD2.n175 VDD2.n112 12.0247
R3657 VDD2.n139 VDD2.n131 12.0247
R3658 VDD2.n36 VDD2.n28 12.0247
R3659 VDD2.n73 VDD2.n72 12.0247
R3660 VDD2.n85 VDD2.n6 12.0247
R3661 VDD2.n187 VDD2.n105 11.249
R3662 VDD2.n174 VDD2.n115 11.249
R3663 VDD2.n143 VDD2.n142 11.249
R3664 VDD2.n40 VDD2.n39 11.249
R3665 VDD2.n71 VDD2.n12 11.249
R3666 VDD2.n86 VDD2.n4 11.249
R3667 VDD2.n191 VDD2.n190 10.4732
R3668 VDD2.n171 VDD2.n170 10.4732
R3669 VDD2.n146 VDD2.n129 10.4732
R3670 VDD2.n43 VDD2.n26 10.4732
R3671 VDD2.n68 VDD2.n67 10.4732
R3672 VDD2.n90 VDD2.n89 10.4732
R3673 VDD2.n194 VDD2.n103 9.69747
R3674 VDD2.n167 VDD2.n117 9.69747
R3675 VDD2.n147 VDD2.n127 9.69747
R3676 VDD2.n44 VDD2.n24 9.69747
R3677 VDD2.n64 VDD2.n14 9.69747
R3678 VDD2.n93 VDD2.n2 9.69747
R3679 VDD2.n197 VDD2.n196 9.45567
R3680 VDD2.n96 VDD2.n95 9.45567
R3681 VDD2.n121 VDD2.n120 9.3005
R3682 VDD2.n164 VDD2.n163 9.3005
R3683 VDD2.n166 VDD2.n165 9.3005
R3684 VDD2.n117 VDD2.n116 9.3005
R3685 VDD2.n172 VDD2.n171 9.3005
R3686 VDD2.n174 VDD2.n173 9.3005
R3687 VDD2.n112 VDD2.n110 9.3005
R3688 VDD2.n180 VDD2.n179 9.3005
R3689 VDD2.n196 VDD2.n195 9.3005
R3690 VDD2.n103 VDD2.n102 9.3005
R3691 VDD2.n190 VDD2.n189 9.3005
R3692 VDD2.n188 VDD2.n187 9.3005
R3693 VDD2.n107 VDD2.n106 9.3005
R3694 VDD2.n182 VDD2.n181 9.3005
R3695 VDD2.n158 VDD2.n157 9.3005
R3696 VDD2.n156 VDD2.n155 9.3005
R3697 VDD2.n125 VDD2.n124 9.3005
R3698 VDD2.n150 VDD2.n149 9.3005
R3699 VDD2.n148 VDD2.n147 9.3005
R3700 VDD2.n129 VDD2.n128 9.3005
R3701 VDD2.n142 VDD2.n141 9.3005
R3702 VDD2.n140 VDD2.n139 9.3005
R3703 VDD2.n133 VDD2.n132 9.3005
R3704 VDD2.n95 VDD2.n94 9.3005
R3705 VDD2.n2 VDD2.n1 9.3005
R3706 VDD2.n89 VDD2.n88 9.3005
R3707 VDD2.n87 VDD2.n86 9.3005
R3708 VDD2.n6 VDD2.n5 9.3005
R3709 VDD2.n81 VDD2.n80 9.3005
R3710 VDD2.n53 VDD2.n52 9.3005
R3711 VDD2.n22 VDD2.n21 9.3005
R3712 VDD2.n47 VDD2.n46 9.3005
R3713 VDD2.n45 VDD2.n44 9.3005
R3714 VDD2.n26 VDD2.n25 9.3005
R3715 VDD2.n39 VDD2.n38 9.3005
R3716 VDD2.n37 VDD2.n36 9.3005
R3717 VDD2.n30 VDD2.n29 9.3005
R3718 VDD2.n55 VDD2.n54 9.3005
R3719 VDD2.n18 VDD2.n17 9.3005
R3720 VDD2.n61 VDD2.n60 9.3005
R3721 VDD2.n63 VDD2.n62 9.3005
R3722 VDD2.n14 VDD2.n13 9.3005
R3723 VDD2.n69 VDD2.n68 9.3005
R3724 VDD2.n71 VDD2.n70 9.3005
R3725 VDD2.n72 VDD2.n9 9.3005
R3726 VDD2.n79 VDD2.n78 9.3005
R3727 VDD2.n195 VDD2.n101 8.92171
R3728 VDD2.n166 VDD2.n119 8.92171
R3729 VDD2.n151 VDD2.n150 8.92171
R3730 VDD2.n48 VDD2.n47 8.92171
R3731 VDD2.n63 VDD2.n16 8.92171
R3732 VDD2.n94 VDD2.n0 8.92171
R3733 VDD2.n163 VDD2.n162 8.14595
R3734 VDD2.n154 VDD2.n125 8.14595
R3735 VDD2.n51 VDD2.n22 8.14595
R3736 VDD2.n60 VDD2.n59 8.14595
R3737 VDD2.n159 VDD2.n121 7.3702
R3738 VDD2.n155 VDD2.n123 7.3702
R3739 VDD2.n52 VDD2.n20 7.3702
R3740 VDD2.n56 VDD2.n18 7.3702
R3741 VDD2.n159 VDD2.n158 6.59444
R3742 VDD2.n158 VDD2.n123 6.59444
R3743 VDD2.n55 VDD2.n20 6.59444
R3744 VDD2.n56 VDD2.n55 6.59444
R3745 VDD2.n162 VDD2.n121 5.81868
R3746 VDD2.n155 VDD2.n154 5.81868
R3747 VDD2.n52 VDD2.n51 5.81868
R3748 VDD2.n59 VDD2.n18 5.81868
R3749 VDD2.n197 VDD2.n101 5.04292
R3750 VDD2.n163 VDD2.n119 5.04292
R3751 VDD2.n151 VDD2.n125 5.04292
R3752 VDD2.n48 VDD2.n22 5.04292
R3753 VDD2.n60 VDD2.n16 5.04292
R3754 VDD2.n96 VDD2.n0 5.04292
R3755 VDD2.n134 VDD2.n132 4.38563
R3756 VDD2.n31 VDD2.n29 4.38563
R3757 VDD2.n195 VDD2.n194 4.26717
R3758 VDD2.n167 VDD2.n166 4.26717
R3759 VDD2.n150 VDD2.n127 4.26717
R3760 VDD2.n47 VDD2.n24 4.26717
R3761 VDD2.n64 VDD2.n63 4.26717
R3762 VDD2.n94 VDD2.n93 4.26717
R3763 VDD2.n191 VDD2.n103 3.49141
R3764 VDD2.n170 VDD2.n117 3.49141
R3765 VDD2.n147 VDD2.n146 3.49141
R3766 VDD2.n44 VDD2.n43 3.49141
R3767 VDD2.n67 VDD2.n14 3.49141
R3768 VDD2.n90 VDD2.n2 3.49141
R3769 VDD2.n200 VDD2.n198 2.97464
R3770 VDD2.n190 VDD2.n105 2.71565
R3771 VDD2.n171 VDD2.n115 2.71565
R3772 VDD2.n143 VDD2.n129 2.71565
R3773 VDD2.n40 VDD2.n26 2.71565
R3774 VDD2.n68 VDD2.n12 2.71565
R3775 VDD2.n89 VDD2.n4 2.71565
R3776 VDD2.n187 VDD2.n186 1.93989
R3777 VDD2.n175 VDD2.n174 1.93989
R3778 VDD2.n142 VDD2.n131 1.93989
R3779 VDD2.n39 VDD2.n28 1.93989
R3780 VDD2.n73 VDD2.n71 1.93989
R3781 VDD2.n86 VDD2.n85 1.93989
R3782 VDD2.n183 VDD2.n107 1.16414
R3783 VDD2.n178 VDD2.n112 1.16414
R3784 VDD2.n139 VDD2.n138 1.16414
R3785 VDD2.n36 VDD2.n35 1.16414
R3786 VDD2.n72 VDD2.n10 1.16414
R3787 VDD2.n82 VDD2.n6 1.16414
R3788 VDD2.n201 VDD2.t2 1.12678
R3789 VDD2.n201 VDD2.t3 1.12678
R3790 VDD2.n199 VDD2.t1 1.12678
R3791 VDD2.n199 VDD2.t9 1.12678
R3792 VDD2.n99 VDD2.t8 1.12678
R3793 VDD2.n99 VDD2.t4 1.12678
R3794 VDD2.n97 VDD2.t0 1.12678
R3795 VDD2.n97 VDD2.t5 1.12678
R3796 VDD2 VDD2.n200 0.802224
R3797 VDD2.n100 VDD2.n98 0.688688
R3798 VDD2.n182 VDD2.n109 0.388379
R3799 VDD2.n179 VDD2.n111 0.388379
R3800 VDD2.n135 VDD2.n133 0.388379
R3801 VDD2.n32 VDD2.n30 0.388379
R3802 VDD2.n78 VDD2.n77 0.388379
R3803 VDD2.n81 VDD2.n8 0.388379
R3804 VDD2.n196 VDD2.n102 0.155672
R3805 VDD2.n189 VDD2.n102 0.155672
R3806 VDD2.n189 VDD2.n188 0.155672
R3807 VDD2.n188 VDD2.n106 0.155672
R3808 VDD2.n181 VDD2.n106 0.155672
R3809 VDD2.n181 VDD2.n180 0.155672
R3810 VDD2.n180 VDD2.n110 0.155672
R3811 VDD2.n173 VDD2.n110 0.155672
R3812 VDD2.n173 VDD2.n172 0.155672
R3813 VDD2.n172 VDD2.n116 0.155672
R3814 VDD2.n165 VDD2.n116 0.155672
R3815 VDD2.n165 VDD2.n164 0.155672
R3816 VDD2.n164 VDD2.n120 0.155672
R3817 VDD2.n157 VDD2.n120 0.155672
R3818 VDD2.n157 VDD2.n156 0.155672
R3819 VDD2.n156 VDD2.n124 0.155672
R3820 VDD2.n149 VDD2.n124 0.155672
R3821 VDD2.n149 VDD2.n148 0.155672
R3822 VDD2.n148 VDD2.n128 0.155672
R3823 VDD2.n141 VDD2.n128 0.155672
R3824 VDD2.n141 VDD2.n140 0.155672
R3825 VDD2.n140 VDD2.n132 0.155672
R3826 VDD2.n37 VDD2.n29 0.155672
R3827 VDD2.n38 VDD2.n37 0.155672
R3828 VDD2.n38 VDD2.n25 0.155672
R3829 VDD2.n45 VDD2.n25 0.155672
R3830 VDD2.n46 VDD2.n45 0.155672
R3831 VDD2.n46 VDD2.n21 0.155672
R3832 VDD2.n53 VDD2.n21 0.155672
R3833 VDD2.n54 VDD2.n53 0.155672
R3834 VDD2.n54 VDD2.n17 0.155672
R3835 VDD2.n61 VDD2.n17 0.155672
R3836 VDD2.n62 VDD2.n61 0.155672
R3837 VDD2.n62 VDD2.n13 0.155672
R3838 VDD2.n69 VDD2.n13 0.155672
R3839 VDD2.n70 VDD2.n69 0.155672
R3840 VDD2.n70 VDD2.n9 0.155672
R3841 VDD2.n79 VDD2.n9 0.155672
R3842 VDD2.n80 VDD2.n79 0.155672
R3843 VDD2.n80 VDD2.n5 0.155672
R3844 VDD2.n87 VDD2.n5 0.155672
R3845 VDD2.n88 VDD2.n87 0.155672
R3846 VDD2.n88 VDD2.n1 0.155672
R3847 VDD2.n95 VDD2.n1 0.155672
C0 VDD1 VN 0.155049f
C1 VDD2 VN 15.9115f
C2 VDD1 VTAIL 12.9393f
C3 VDD2 VTAIL 12.9931f
C4 VP VN 10.1912f
C5 VDD1 VDD2 2.51479f
C6 VP VTAIL 16.536098f
C7 VP VDD1 16.4026f
C8 VP VDD2 0.650805f
C9 VN VTAIL 16.521801f
C10 VDD2 B 8.786064f
C11 VDD1 B 8.77225f
C12 VTAIL B 10.866854f
C13 VN B 21.052319f
C14 VP B 19.550865f
C15 VDD2.n0 B 0.033535f
C16 VDD2.n1 B 0.023632f
C17 VDD2.n2 B 0.012699f
C18 VDD2.n3 B 0.030015f
C19 VDD2.n4 B 0.013446f
C20 VDD2.n5 B 0.023632f
C21 VDD2.n6 B 0.012699f
C22 VDD2.n7 B 0.030015f
C23 VDD2.n8 B 0.013072f
C24 VDD2.n9 B 0.023632f
C25 VDD2.n10 B 0.013446f
C26 VDD2.n11 B 0.030015f
C27 VDD2.n12 B 0.013446f
C28 VDD2.n13 B 0.023632f
C29 VDD2.n14 B 0.012699f
C30 VDD2.n15 B 0.030015f
C31 VDD2.n16 B 0.013446f
C32 VDD2.n17 B 0.023632f
C33 VDD2.n18 B 0.012699f
C34 VDD2.n19 B 0.030015f
C35 VDD2.n20 B 0.013446f
C36 VDD2.n21 B 0.023632f
C37 VDD2.n22 B 0.012699f
C38 VDD2.n23 B 0.030015f
C39 VDD2.n24 B 0.013446f
C40 VDD2.n25 B 0.023632f
C41 VDD2.n26 B 0.012699f
C42 VDD2.n27 B 0.030015f
C43 VDD2.n28 B 0.013446f
C44 VDD2.n29 B 1.81694f
C45 VDD2.n30 B 0.012699f
C46 VDD2.t6 B 0.0497f
C47 VDD2.n31 B 0.169418f
C48 VDD2.n32 B 0.017731f
C49 VDD2.n33 B 0.022511f
C50 VDD2.n34 B 0.030015f
C51 VDD2.n35 B 0.013446f
C52 VDD2.n36 B 0.012699f
C53 VDD2.n37 B 0.023632f
C54 VDD2.n38 B 0.023632f
C55 VDD2.n39 B 0.012699f
C56 VDD2.n40 B 0.013446f
C57 VDD2.n41 B 0.030015f
C58 VDD2.n42 B 0.030015f
C59 VDD2.n43 B 0.013446f
C60 VDD2.n44 B 0.012699f
C61 VDD2.n45 B 0.023632f
C62 VDD2.n46 B 0.023632f
C63 VDD2.n47 B 0.012699f
C64 VDD2.n48 B 0.013446f
C65 VDD2.n49 B 0.030015f
C66 VDD2.n50 B 0.030015f
C67 VDD2.n51 B 0.013446f
C68 VDD2.n52 B 0.012699f
C69 VDD2.n53 B 0.023632f
C70 VDD2.n54 B 0.023632f
C71 VDD2.n55 B 0.012699f
C72 VDD2.n56 B 0.013446f
C73 VDD2.n57 B 0.030015f
C74 VDD2.n58 B 0.030015f
C75 VDD2.n59 B 0.013446f
C76 VDD2.n60 B 0.012699f
C77 VDD2.n61 B 0.023632f
C78 VDD2.n62 B 0.023632f
C79 VDD2.n63 B 0.012699f
C80 VDD2.n64 B 0.013446f
C81 VDD2.n65 B 0.030015f
C82 VDD2.n66 B 0.030015f
C83 VDD2.n67 B 0.013446f
C84 VDD2.n68 B 0.012699f
C85 VDD2.n69 B 0.023632f
C86 VDD2.n70 B 0.023632f
C87 VDD2.n71 B 0.012699f
C88 VDD2.n72 B 0.012699f
C89 VDD2.n73 B 0.013446f
C90 VDD2.n74 B 0.030015f
C91 VDD2.n75 B 0.030015f
C92 VDD2.n76 B 0.030015f
C93 VDD2.n77 B 0.013072f
C94 VDD2.n78 B 0.012699f
C95 VDD2.n79 B 0.023632f
C96 VDD2.n80 B 0.023632f
C97 VDD2.n81 B 0.012699f
C98 VDD2.n82 B 0.013446f
C99 VDD2.n83 B 0.030015f
C100 VDD2.n84 B 0.030015f
C101 VDD2.n85 B 0.013446f
C102 VDD2.n86 B 0.012699f
C103 VDD2.n87 B 0.023632f
C104 VDD2.n88 B 0.023632f
C105 VDD2.n89 B 0.012699f
C106 VDD2.n90 B 0.013446f
C107 VDD2.n91 B 0.030015f
C108 VDD2.n92 B 0.065541f
C109 VDD2.n93 B 0.013446f
C110 VDD2.n94 B 0.012699f
C111 VDD2.n95 B 0.056561f
C112 VDD2.n96 B 0.068416f
C113 VDD2.t0 B 0.328298f
C114 VDD2.t5 B 0.328298f
C115 VDD2.n97 B 2.98908f
C116 VDD2.n98 B 0.732287f
C117 VDD2.t8 B 0.328298f
C118 VDD2.t4 B 0.328298f
C119 VDD2.n99 B 3.00935f
C120 VDD2.n100 B 3.33378f
C121 VDD2.n101 B 0.033535f
C122 VDD2.n102 B 0.023632f
C123 VDD2.n103 B 0.012699f
C124 VDD2.n104 B 0.030015f
C125 VDD2.n105 B 0.013446f
C126 VDD2.n106 B 0.023632f
C127 VDD2.n107 B 0.012699f
C128 VDD2.n108 B 0.030015f
C129 VDD2.n109 B 0.013072f
C130 VDD2.n110 B 0.023632f
C131 VDD2.n111 B 0.013072f
C132 VDD2.n112 B 0.012699f
C133 VDD2.n113 B 0.030015f
C134 VDD2.n114 B 0.030015f
C135 VDD2.n115 B 0.013446f
C136 VDD2.n116 B 0.023632f
C137 VDD2.n117 B 0.012699f
C138 VDD2.n118 B 0.030015f
C139 VDD2.n119 B 0.013446f
C140 VDD2.n120 B 0.023632f
C141 VDD2.n121 B 0.012699f
C142 VDD2.n122 B 0.030015f
C143 VDD2.n123 B 0.013446f
C144 VDD2.n124 B 0.023632f
C145 VDD2.n125 B 0.012699f
C146 VDD2.n126 B 0.030015f
C147 VDD2.n127 B 0.013446f
C148 VDD2.n128 B 0.023632f
C149 VDD2.n129 B 0.012699f
C150 VDD2.n130 B 0.030015f
C151 VDD2.n131 B 0.013446f
C152 VDD2.n132 B 1.81694f
C153 VDD2.n133 B 0.012699f
C154 VDD2.t7 B 0.0497f
C155 VDD2.n134 B 0.169418f
C156 VDD2.n135 B 0.017731f
C157 VDD2.n136 B 0.022511f
C158 VDD2.n137 B 0.030015f
C159 VDD2.n138 B 0.013446f
C160 VDD2.n139 B 0.012699f
C161 VDD2.n140 B 0.023632f
C162 VDD2.n141 B 0.023632f
C163 VDD2.n142 B 0.012699f
C164 VDD2.n143 B 0.013446f
C165 VDD2.n144 B 0.030015f
C166 VDD2.n145 B 0.030015f
C167 VDD2.n146 B 0.013446f
C168 VDD2.n147 B 0.012699f
C169 VDD2.n148 B 0.023632f
C170 VDD2.n149 B 0.023632f
C171 VDD2.n150 B 0.012699f
C172 VDD2.n151 B 0.013446f
C173 VDD2.n152 B 0.030015f
C174 VDD2.n153 B 0.030015f
C175 VDD2.n154 B 0.013446f
C176 VDD2.n155 B 0.012699f
C177 VDD2.n156 B 0.023632f
C178 VDD2.n157 B 0.023632f
C179 VDD2.n158 B 0.012699f
C180 VDD2.n159 B 0.013446f
C181 VDD2.n160 B 0.030015f
C182 VDD2.n161 B 0.030015f
C183 VDD2.n162 B 0.013446f
C184 VDD2.n163 B 0.012699f
C185 VDD2.n164 B 0.023632f
C186 VDD2.n165 B 0.023632f
C187 VDD2.n166 B 0.012699f
C188 VDD2.n167 B 0.013446f
C189 VDD2.n168 B 0.030015f
C190 VDD2.n169 B 0.030015f
C191 VDD2.n170 B 0.013446f
C192 VDD2.n171 B 0.012699f
C193 VDD2.n172 B 0.023632f
C194 VDD2.n173 B 0.023632f
C195 VDD2.n174 B 0.012699f
C196 VDD2.n175 B 0.013446f
C197 VDD2.n176 B 0.030015f
C198 VDD2.n177 B 0.030015f
C199 VDD2.n178 B 0.013446f
C200 VDD2.n179 B 0.012699f
C201 VDD2.n180 B 0.023632f
C202 VDD2.n181 B 0.023632f
C203 VDD2.n182 B 0.012699f
C204 VDD2.n183 B 0.013446f
C205 VDD2.n184 B 0.030015f
C206 VDD2.n185 B 0.030015f
C207 VDD2.n186 B 0.013446f
C208 VDD2.n187 B 0.012699f
C209 VDD2.n188 B 0.023632f
C210 VDD2.n189 B 0.023632f
C211 VDD2.n190 B 0.012699f
C212 VDD2.n191 B 0.013446f
C213 VDD2.n192 B 0.030015f
C214 VDD2.n193 B 0.065541f
C215 VDD2.n194 B 0.013446f
C216 VDD2.n195 B 0.012699f
C217 VDD2.n196 B 0.056561f
C218 VDD2.n197 B 0.053092f
C219 VDD2.n198 B 3.32615f
C220 VDD2.t1 B 0.328298f
C221 VDD2.t9 B 0.328298f
C222 VDD2.n199 B 2.98908f
C223 VDD2.n200 B 0.482367f
C224 VDD2.t2 B 0.328298f
C225 VDD2.t3 B 0.328298f
C226 VDD2.n201 B 3.00931f
C227 VN.t5 B 2.73716f
C228 VN.n0 B 1.01987f
C229 VN.n1 B 0.018151f
C230 VN.n2 B 0.022619f
C231 VN.n3 B 0.018151f
C232 VN.t1 B 2.73716f
C233 VN.n4 B 0.946638f
C234 VN.n5 B 0.018151f
C235 VN.n6 B 0.02513f
C236 VN.n7 B 0.018151f
C237 VN.t4 B 2.73716f
C238 VN.n8 B 0.033659f
C239 VN.n9 B 0.018151f
C240 VN.n10 B 0.033659f
C241 VN.t3 B 2.94976f
C242 VN.n11 B 0.969659f
C243 VN.t9 B 2.73716f
C244 VN.n12 B 1.01234f
C245 VN.n13 B 0.031998f
C246 VN.n14 B 0.207471f
C247 VN.n15 B 0.018151f
C248 VN.n16 B 0.018151f
C249 VN.n17 B 0.027641f
C250 VN.n18 B 0.02513f
C251 VN.n19 B 0.033659f
C252 VN.n20 B 0.018151f
C253 VN.n21 B 0.018151f
C254 VN.n22 B 0.018151f
C255 VN.n23 B 0.96368f
C256 VN.n24 B 0.033659f
C257 VN.n25 B 0.033659f
C258 VN.n26 B 0.018151f
C259 VN.n27 B 0.018151f
C260 VN.n28 B 0.018151f
C261 VN.n29 B 0.027641f
C262 VN.n30 B 0.033659f
C263 VN.n31 B 0.031998f
C264 VN.n32 B 0.018151f
C265 VN.n33 B 0.018151f
C266 VN.n34 B 0.018704f
C267 VN.n35 B 0.033659f
C268 VN.n36 B 0.033659f
C269 VN.n37 B 0.018151f
C270 VN.n38 B 0.018151f
C271 VN.n39 B 0.018151f
C272 VN.n40 B 0.030152f
C273 VN.n41 B 0.033659f
C274 VN.n42 B 0.030336f
C275 VN.n43 B 0.029291f
C276 VN.n44 B 0.038824f
C277 VN.t2 B 2.73716f
C278 VN.n45 B 1.01987f
C279 VN.n46 B 0.018151f
C280 VN.n47 B 0.022619f
C281 VN.n48 B 0.018151f
C282 VN.t8 B 2.73716f
C283 VN.n49 B 0.946638f
C284 VN.n50 B 0.018151f
C285 VN.n51 B 0.02513f
C286 VN.n52 B 0.018151f
C287 VN.t0 B 2.73716f
C288 VN.n53 B 0.033659f
C289 VN.n54 B 0.018151f
C290 VN.n55 B 0.033659f
C291 VN.t6 B 2.94976f
C292 VN.n56 B 0.969659f
C293 VN.t7 B 2.73716f
C294 VN.n57 B 1.01234f
C295 VN.n58 B 0.031998f
C296 VN.n59 B 0.207471f
C297 VN.n60 B 0.018151f
C298 VN.n61 B 0.018151f
C299 VN.n62 B 0.027641f
C300 VN.n63 B 0.02513f
C301 VN.n64 B 0.033659f
C302 VN.n65 B 0.018151f
C303 VN.n66 B 0.018151f
C304 VN.n67 B 0.018151f
C305 VN.n68 B 0.96368f
C306 VN.n69 B 0.033659f
C307 VN.n70 B 0.033659f
C308 VN.n71 B 0.018151f
C309 VN.n72 B 0.018151f
C310 VN.n73 B 0.018151f
C311 VN.n74 B 0.027641f
C312 VN.n75 B 0.033659f
C313 VN.n76 B 0.031998f
C314 VN.n77 B 0.018151f
C315 VN.n78 B 0.018151f
C316 VN.n79 B 0.018704f
C317 VN.n80 B 0.033659f
C318 VN.n81 B 0.033659f
C319 VN.n82 B 0.018151f
C320 VN.n83 B 0.018151f
C321 VN.n84 B 0.018151f
C322 VN.n85 B 0.030152f
C323 VN.n86 B 0.033659f
C324 VN.n87 B 0.030336f
C325 VN.n88 B 0.029291f
C326 VN.n89 B 1.34045f
C327 VTAIL.t5 B 0.332621f
C328 VTAIL.t6 B 0.332621f
C329 VTAIL.n0 B 2.95722f
C330 VTAIL.n1 B 0.563652f
C331 VTAIL.n2 B 0.033977f
C332 VTAIL.n3 B 0.023943f
C333 VTAIL.n4 B 0.012866f
C334 VTAIL.n5 B 0.03041f
C335 VTAIL.n6 B 0.013623f
C336 VTAIL.n7 B 0.023943f
C337 VTAIL.n8 B 0.012866f
C338 VTAIL.n9 B 0.03041f
C339 VTAIL.n10 B 0.013244f
C340 VTAIL.n11 B 0.023943f
C341 VTAIL.n12 B 0.013623f
C342 VTAIL.n13 B 0.03041f
C343 VTAIL.n14 B 0.013623f
C344 VTAIL.n15 B 0.023943f
C345 VTAIL.n16 B 0.012866f
C346 VTAIL.n17 B 0.03041f
C347 VTAIL.n18 B 0.013623f
C348 VTAIL.n19 B 0.023943f
C349 VTAIL.n20 B 0.012866f
C350 VTAIL.n21 B 0.03041f
C351 VTAIL.n22 B 0.013623f
C352 VTAIL.n23 B 0.023943f
C353 VTAIL.n24 B 0.012866f
C354 VTAIL.n25 B 0.03041f
C355 VTAIL.n26 B 0.013623f
C356 VTAIL.n27 B 0.023943f
C357 VTAIL.n28 B 0.012866f
C358 VTAIL.n29 B 0.03041f
C359 VTAIL.n30 B 0.013623f
C360 VTAIL.n31 B 1.84086f
C361 VTAIL.n32 B 0.012866f
C362 VTAIL.t17 B 0.050355f
C363 VTAIL.n33 B 0.171649f
C364 VTAIL.n34 B 0.017964f
C365 VTAIL.n35 B 0.022808f
C366 VTAIL.n36 B 0.03041f
C367 VTAIL.n37 B 0.013623f
C368 VTAIL.n38 B 0.012866f
C369 VTAIL.n39 B 0.023943f
C370 VTAIL.n40 B 0.023943f
C371 VTAIL.n41 B 0.012866f
C372 VTAIL.n42 B 0.013623f
C373 VTAIL.n43 B 0.03041f
C374 VTAIL.n44 B 0.03041f
C375 VTAIL.n45 B 0.013623f
C376 VTAIL.n46 B 0.012866f
C377 VTAIL.n47 B 0.023943f
C378 VTAIL.n48 B 0.023943f
C379 VTAIL.n49 B 0.012866f
C380 VTAIL.n50 B 0.013623f
C381 VTAIL.n51 B 0.03041f
C382 VTAIL.n52 B 0.03041f
C383 VTAIL.n53 B 0.013623f
C384 VTAIL.n54 B 0.012866f
C385 VTAIL.n55 B 0.023943f
C386 VTAIL.n56 B 0.023943f
C387 VTAIL.n57 B 0.012866f
C388 VTAIL.n58 B 0.013623f
C389 VTAIL.n59 B 0.03041f
C390 VTAIL.n60 B 0.03041f
C391 VTAIL.n61 B 0.013623f
C392 VTAIL.n62 B 0.012866f
C393 VTAIL.n63 B 0.023943f
C394 VTAIL.n64 B 0.023943f
C395 VTAIL.n65 B 0.012866f
C396 VTAIL.n66 B 0.013623f
C397 VTAIL.n67 B 0.03041f
C398 VTAIL.n68 B 0.03041f
C399 VTAIL.n69 B 0.013623f
C400 VTAIL.n70 B 0.012866f
C401 VTAIL.n71 B 0.023943f
C402 VTAIL.n72 B 0.023943f
C403 VTAIL.n73 B 0.012866f
C404 VTAIL.n74 B 0.012866f
C405 VTAIL.n75 B 0.013623f
C406 VTAIL.n76 B 0.03041f
C407 VTAIL.n77 B 0.03041f
C408 VTAIL.n78 B 0.03041f
C409 VTAIL.n79 B 0.013244f
C410 VTAIL.n80 B 0.012866f
C411 VTAIL.n81 B 0.023943f
C412 VTAIL.n82 B 0.023943f
C413 VTAIL.n83 B 0.012866f
C414 VTAIL.n84 B 0.013623f
C415 VTAIL.n85 B 0.03041f
C416 VTAIL.n86 B 0.03041f
C417 VTAIL.n87 B 0.013623f
C418 VTAIL.n88 B 0.012866f
C419 VTAIL.n89 B 0.023943f
C420 VTAIL.n90 B 0.023943f
C421 VTAIL.n91 B 0.012866f
C422 VTAIL.n92 B 0.013623f
C423 VTAIL.n93 B 0.03041f
C424 VTAIL.n94 B 0.066404f
C425 VTAIL.n95 B 0.013623f
C426 VTAIL.n96 B 0.012866f
C427 VTAIL.n97 B 0.057305f
C428 VTAIL.n98 B 0.037274f
C429 VTAIL.n99 B 0.401984f
C430 VTAIL.t16 B 0.332621f
C431 VTAIL.t11 B 0.332621f
C432 VTAIL.n100 B 2.95722f
C433 VTAIL.n101 B 0.695006f
C434 VTAIL.t15 B 0.332621f
C435 VTAIL.t14 B 0.332621f
C436 VTAIL.n102 B 2.95722f
C437 VTAIL.n103 B 2.41891f
C438 VTAIL.t8 B 0.332621f
C439 VTAIL.t7 B 0.332621f
C440 VTAIL.n104 B 2.95723f
C441 VTAIL.n105 B 2.41889f
C442 VTAIL.t0 B 0.332621f
C443 VTAIL.t9 B 0.332621f
C444 VTAIL.n106 B 2.95723f
C445 VTAIL.n107 B 0.694993f
C446 VTAIL.n108 B 0.033977f
C447 VTAIL.n109 B 0.023943f
C448 VTAIL.n110 B 0.012866f
C449 VTAIL.n111 B 0.03041f
C450 VTAIL.n112 B 0.013623f
C451 VTAIL.n113 B 0.023943f
C452 VTAIL.n114 B 0.012866f
C453 VTAIL.n115 B 0.03041f
C454 VTAIL.n116 B 0.013244f
C455 VTAIL.n117 B 0.023943f
C456 VTAIL.n118 B 0.013244f
C457 VTAIL.n119 B 0.012866f
C458 VTAIL.n120 B 0.03041f
C459 VTAIL.n121 B 0.03041f
C460 VTAIL.n122 B 0.013623f
C461 VTAIL.n123 B 0.023943f
C462 VTAIL.n124 B 0.012866f
C463 VTAIL.n125 B 0.03041f
C464 VTAIL.n126 B 0.013623f
C465 VTAIL.n127 B 0.023943f
C466 VTAIL.n128 B 0.012866f
C467 VTAIL.n129 B 0.03041f
C468 VTAIL.n130 B 0.013623f
C469 VTAIL.n131 B 0.023943f
C470 VTAIL.n132 B 0.012866f
C471 VTAIL.n133 B 0.03041f
C472 VTAIL.n134 B 0.013623f
C473 VTAIL.n135 B 0.023943f
C474 VTAIL.n136 B 0.012866f
C475 VTAIL.n137 B 0.03041f
C476 VTAIL.n138 B 0.013623f
C477 VTAIL.n139 B 1.84087f
C478 VTAIL.n140 B 0.012866f
C479 VTAIL.t1 B 0.050355f
C480 VTAIL.n141 B 0.171649f
C481 VTAIL.n142 B 0.017964f
C482 VTAIL.n143 B 0.022808f
C483 VTAIL.n144 B 0.03041f
C484 VTAIL.n145 B 0.013623f
C485 VTAIL.n146 B 0.012866f
C486 VTAIL.n147 B 0.023943f
C487 VTAIL.n148 B 0.023943f
C488 VTAIL.n149 B 0.012866f
C489 VTAIL.n150 B 0.013623f
C490 VTAIL.n151 B 0.03041f
C491 VTAIL.n152 B 0.03041f
C492 VTAIL.n153 B 0.013623f
C493 VTAIL.n154 B 0.012866f
C494 VTAIL.n155 B 0.023943f
C495 VTAIL.n156 B 0.023943f
C496 VTAIL.n157 B 0.012866f
C497 VTAIL.n158 B 0.013623f
C498 VTAIL.n159 B 0.03041f
C499 VTAIL.n160 B 0.03041f
C500 VTAIL.n161 B 0.013623f
C501 VTAIL.n162 B 0.012866f
C502 VTAIL.n163 B 0.023943f
C503 VTAIL.n164 B 0.023943f
C504 VTAIL.n165 B 0.012866f
C505 VTAIL.n166 B 0.013623f
C506 VTAIL.n167 B 0.03041f
C507 VTAIL.n168 B 0.03041f
C508 VTAIL.n169 B 0.013623f
C509 VTAIL.n170 B 0.012866f
C510 VTAIL.n171 B 0.023943f
C511 VTAIL.n172 B 0.023943f
C512 VTAIL.n173 B 0.012866f
C513 VTAIL.n174 B 0.013623f
C514 VTAIL.n175 B 0.03041f
C515 VTAIL.n176 B 0.03041f
C516 VTAIL.n177 B 0.013623f
C517 VTAIL.n178 B 0.012866f
C518 VTAIL.n179 B 0.023943f
C519 VTAIL.n180 B 0.023943f
C520 VTAIL.n181 B 0.012866f
C521 VTAIL.n182 B 0.013623f
C522 VTAIL.n183 B 0.03041f
C523 VTAIL.n184 B 0.03041f
C524 VTAIL.n185 B 0.013623f
C525 VTAIL.n186 B 0.012866f
C526 VTAIL.n187 B 0.023943f
C527 VTAIL.n188 B 0.023943f
C528 VTAIL.n189 B 0.012866f
C529 VTAIL.n190 B 0.013623f
C530 VTAIL.n191 B 0.03041f
C531 VTAIL.n192 B 0.03041f
C532 VTAIL.n193 B 0.013623f
C533 VTAIL.n194 B 0.012866f
C534 VTAIL.n195 B 0.023943f
C535 VTAIL.n196 B 0.023943f
C536 VTAIL.n197 B 0.012866f
C537 VTAIL.n198 B 0.013623f
C538 VTAIL.n199 B 0.03041f
C539 VTAIL.n200 B 0.066404f
C540 VTAIL.n201 B 0.013623f
C541 VTAIL.n202 B 0.012866f
C542 VTAIL.n203 B 0.057305f
C543 VTAIL.n204 B 0.037274f
C544 VTAIL.n205 B 0.401984f
C545 VTAIL.t12 B 0.332621f
C546 VTAIL.t19 B 0.332621f
C547 VTAIL.n206 B 2.95723f
C548 VTAIL.n207 B 0.616513f
C549 VTAIL.t13 B 0.332621f
C550 VTAIL.t18 B 0.332621f
C551 VTAIL.n208 B 2.95723f
C552 VTAIL.n209 B 0.694993f
C553 VTAIL.n210 B 0.033977f
C554 VTAIL.n211 B 0.023943f
C555 VTAIL.n212 B 0.012866f
C556 VTAIL.n213 B 0.03041f
C557 VTAIL.n214 B 0.013623f
C558 VTAIL.n215 B 0.023943f
C559 VTAIL.n216 B 0.012866f
C560 VTAIL.n217 B 0.03041f
C561 VTAIL.n218 B 0.013244f
C562 VTAIL.n219 B 0.023943f
C563 VTAIL.n220 B 0.013244f
C564 VTAIL.n221 B 0.012866f
C565 VTAIL.n222 B 0.03041f
C566 VTAIL.n223 B 0.03041f
C567 VTAIL.n224 B 0.013623f
C568 VTAIL.n225 B 0.023943f
C569 VTAIL.n226 B 0.012866f
C570 VTAIL.n227 B 0.03041f
C571 VTAIL.n228 B 0.013623f
C572 VTAIL.n229 B 0.023943f
C573 VTAIL.n230 B 0.012866f
C574 VTAIL.n231 B 0.03041f
C575 VTAIL.n232 B 0.013623f
C576 VTAIL.n233 B 0.023943f
C577 VTAIL.n234 B 0.012866f
C578 VTAIL.n235 B 0.03041f
C579 VTAIL.n236 B 0.013623f
C580 VTAIL.n237 B 0.023943f
C581 VTAIL.n238 B 0.012866f
C582 VTAIL.n239 B 0.03041f
C583 VTAIL.n240 B 0.013623f
C584 VTAIL.n241 B 1.84087f
C585 VTAIL.n242 B 0.012866f
C586 VTAIL.t10 B 0.050355f
C587 VTAIL.n243 B 0.171649f
C588 VTAIL.n244 B 0.017964f
C589 VTAIL.n245 B 0.022808f
C590 VTAIL.n246 B 0.03041f
C591 VTAIL.n247 B 0.013623f
C592 VTAIL.n248 B 0.012866f
C593 VTAIL.n249 B 0.023943f
C594 VTAIL.n250 B 0.023943f
C595 VTAIL.n251 B 0.012866f
C596 VTAIL.n252 B 0.013623f
C597 VTAIL.n253 B 0.03041f
C598 VTAIL.n254 B 0.03041f
C599 VTAIL.n255 B 0.013623f
C600 VTAIL.n256 B 0.012866f
C601 VTAIL.n257 B 0.023943f
C602 VTAIL.n258 B 0.023943f
C603 VTAIL.n259 B 0.012866f
C604 VTAIL.n260 B 0.013623f
C605 VTAIL.n261 B 0.03041f
C606 VTAIL.n262 B 0.03041f
C607 VTAIL.n263 B 0.013623f
C608 VTAIL.n264 B 0.012866f
C609 VTAIL.n265 B 0.023943f
C610 VTAIL.n266 B 0.023943f
C611 VTAIL.n267 B 0.012866f
C612 VTAIL.n268 B 0.013623f
C613 VTAIL.n269 B 0.03041f
C614 VTAIL.n270 B 0.03041f
C615 VTAIL.n271 B 0.013623f
C616 VTAIL.n272 B 0.012866f
C617 VTAIL.n273 B 0.023943f
C618 VTAIL.n274 B 0.023943f
C619 VTAIL.n275 B 0.012866f
C620 VTAIL.n276 B 0.013623f
C621 VTAIL.n277 B 0.03041f
C622 VTAIL.n278 B 0.03041f
C623 VTAIL.n279 B 0.013623f
C624 VTAIL.n280 B 0.012866f
C625 VTAIL.n281 B 0.023943f
C626 VTAIL.n282 B 0.023943f
C627 VTAIL.n283 B 0.012866f
C628 VTAIL.n284 B 0.013623f
C629 VTAIL.n285 B 0.03041f
C630 VTAIL.n286 B 0.03041f
C631 VTAIL.n287 B 0.013623f
C632 VTAIL.n288 B 0.012866f
C633 VTAIL.n289 B 0.023943f
C634 VTAIL.n290 B 0.023943f
C635 VTAIL.n291 B 0.012866f
C636 VTAIL.n292 B 0.013623f
C637 VTAIL.n293 B 0.03041f
C638 VTAIL.n294 B 0.03041f
C639 VTAIL.n295 B 0.013623f
C640 VTAIL.n296 B 0.012866f
C641 VTAIL.n297 B 0.023943f
C642 VTAIL.n298 B 0.023943f
C643 VTAIL.n299 B 0.012866f
C644 VTAIL.n300 B 0.013623f
C645 VTAIL.n301 B 0.03041f
C646 VTAIL.n302 B 0.066404f
C647 VTAIL.n303 B 0.013623f
C648 VTAIL.n304 B 0.012866f
C649 VTAIL.n305 B 0.057305f
C650 VTAIL.n306 B 0.037274f
C651 VTAIL.n307 B 1.97491f
C652 VTAIL.n308 B 0.033977f
C653 VTAIL.n309 B 0.023943f
C654 VTAIL.n310 B 0.012866f
C655 VTAIL.n311 B 0.03041f
C656 VTAIL.n312 B 0.013623f
C657 VTAIL.n313 B 0.023943f
C658 VTAIL.n314 B 0.012866f
C659 VTAIL.n315 B 0.03041f
C660 VTAIL.n316 B 0.013244f
C661 VTAIL.n317 B 0.023943f
C662 VTAIL.n318 B 0.013623f
C663 VTAIL.n319 B 0.03041f
C664 VTAIL.n320 B 0.013623f
C665 VTAIL.n321 B 0.023943f
C666 VTAIL.n322 B 0.012866f
C667 VTAIL.n323 B 0.03041f
C668 VTAIL.n324 B 0.013623f
C669 VTAIL.n325 B 0.023943f
C670 VTAIL.n326 B 0.012866f
C671 VTAIL.n327 B 0.03041f
C672 VTAIL.n328 B 0.013623f
C673 VTAIL.n329 B 0.023943f
C674 VTAIL.n330 B 0.012866f
C675 VTAIL.n331 B 0.03041f
C676 VTAIL.n332 B 0.013623f
C677 VTAIL.n333 B 0.023943f
C678 VTAIL.n334 B 0.012866f
C679 VTAIL.n335 B 0.03041f
C680 VTAIL.n336 B 0.013623f
C681 VTAIL.n337 B 1.84086f
C682 VTAIL.n338 B 0.012866f
C683 VTAIL.t2 B 0.050355f
C684 VTAIL.n339 B 0.171649f
C685 VTAIL.n340 B 0.017964f
C686 VTAIL.n341 B 0.022808f
C687 VTAIL.n342 B 0.03041f
C688 VTAIL.n343 B 0.013623f
C689 VTAIL.n344 B 0.012866f
C690 VTAIL.n345 B 0.023943f
C691 VTAIL.n346 B 0.023943f
C692 VTAIL.n347 B 0.012866f
C693 VTAIL.n348 B 0.013623f
C694 VTAIL.n349 B 0.03041f
C695 VTAIL.n350 B 0.03041f
C696 VTAIL.n351 B 0.013623f
C697 VTAIL.n352 B 0.012866f
C698 VTAIL.n353 B 0.023943f
C699 VTAIL.n354 B 0.023943f
C700 VTAIL.n355 B 0.012866f
C701 VTAIL.n356 B 0.013623f
C702 VTAIL.n357 B 0.03041f
C703 VTAIL.n358 B 0.03041f
C704 VTAIL.n359 B 0.013623f
C705 VTAIL.n360 B 0.012866f
C706 VTAIL.n361 B 0.023943f
C707 VTAIL.n362 B 0.023943f
C708 VTAIL.n363 B 0.012866f
C709 VTAIL.n364 B 0.013623f
C710 VTAIL.n365 B 0.03041f
C711 VTAIL.n366 B 0.03041f
C712 VTAIL.n367 B 0.013623f
C713 VTAIL.n368 B 0.012866f
C714 VTAIL.n369 B 0.023943f
C715 VTAIL.n370 B 0.023943f
C716 VTAIL.n371 B 0.012866f
C717 VTAIL.n372 B 0.013623f
C718 VTAIL.n373 B 0.03041f
C719 VTAIL.n374 B 0.03041f
C720 VTAIL.n375 B 0.013623f
C721 VTAIL.n376 B 0.012866f
C722 VTAIL.n377 B 0.023943f
C723 VTAIL.n378 B 0.023943f
C724 VTAIL.n379 B 0.012866f
C725 VTAIL.n380 B 0.012866f
C726 VTAIL.n381 B 0.013623f
C727 VTAIL.n382 B 0.03041f
C728 VTAIL.n383 B 0.03041f
C729 VTAIL.n384 B 0.03041f
C730 VTAIL.n385 B 0.013244f
C731 VTAIL.n386 B 0.012866f
C732 VTAIL.n387 B 0.023943f
C733 VTAIL.n388 B 0.023943f
C734 VTAIL.n389 B 0.012866f
C735 VTAIL.n390 B 0.013623f
C736 VTAIL.n391 B 0.03041f
C737 VTAIL.n392 B 0.03041f
C738 VTAIL.n393 B 0.013623f
C739 VTAIL.n394 B 0.012866f
C740 VTAIL.n395 B 0.023943f
C741 VTAIL.n396 B 0.023943f
C742 VTAIL.n397 B 0.012866f
C743 VTAIL.n398 B 0.013623f
C744 VTAIL.n399 B 0.03041f
C745 VTAIL.n400 B 0.066404f
C746 VTAIL.n401 B 0.013623f
C747 VTAIL.n402 B 0.012866f
C748 VTAIL.n403 B 0.057305f
C749 VTAIL.n404 B 0.037274f
C750 VTAIL.n405 B 1.97491f
C751 VTAIL.t3 B 0.332621f
C752 VTAIL.t4 B 0.332621f
C753 VTAIL.n406 B 2.95722f
C754 VTAIL.n407 B 0.518427f
C755 VDD1.n0 B 0.033868f
C756 VDD1.n1 B 0.023866f
C757 VDD1.n2 B 0.012825f
C758 VDD1.n3 B 0.030313f
C759 VDD1.n4 B 0.013579f
C760 VDD1.n5 B 0.023866f
C761 VDD1.n6 B 0.012825f
C762 VDD1.n7 B 0.030313f
C763 VDD1.n8 B 0.013202f
C764 VDD1.n9 B 0.023866f
C765 VDD1.n10 B 0.013202f
C766 VDD1.n11 B 0.012825f
C767 VDD1.n12 B 0.030313f
C768 VDD1.n13 B 0.030313f
C769 VDD1.n14 B 0.013579f
C770 VDD1.n15 B 0.023866f
C771 VDD1.n16 B 0.012825f
C772 VDD1.n17 B 0.030313f
C773 VDD1.n18 B 0.013579f
C774 VDD1.n19 B 0.023866f
C775 VDD1.n20 B 0.012825f
C776 VDD1.n21 B 0.030313f
C777 VDD1.n22 B 0.013579f
C778 VDD1.n23 B 0.023866f
C779 VDD1.n24 B 0.012825f
C780 VDD1.n25 B 0.030313f
C781 VDD1.n26 B 0.013579f
C782 VDD1.n27 B 0.023866f
C783 VDD1.n28 B 0.012825f
C784 VDD1.n29 B 0.030313f
C785 VDD1.n30 B 0.013579f
C786 VDD1.n31 B 1.83498f
C787 VDD1.n32 B 0.012825f
C788 VDD1.t6 B 0.050194f
C789 VDD1.n33 B 0.1711f
C790 VDD1.n34 B 0.017907f
C791 VDD1.n35 B 0.022735f
C792 VDD1.n36 B 0.030313f
C793 VDD1.n37 B 0.013579f
C794 VDD1.n38 B 0.012825f
C795 VDD1.n39 B 0.023866f
C796 VDD1.n40 B 0.023866f
C797 VDD1.n41 B 0.012825f
C798 VDD1.n42 B 0.013579f
C799 VDD1.n43 B 0.030313f
C800 VDD1.n44 B 0.030313f
C801 VDD1.n45 B 0.013579f
C802 VDD1.n46 B 0.012825f
C803 VDD1.n47 B 0.023866f
C804 VDD1.n48 B 0.023866f
C805 VDD1.n49 B 0.012825f
C806 VDD1.n50 B 0.013579f
C807 VDD1.n51 B 0.030313f
C808 VDD1.n52 B 0.030313f
C809 VDD1.n53 B 0.013579f
C810 VDD1.n54 B 0.012825f
C811 VDD1.n55 B 0.023866f
C812 VDD1.n56 B 0.023866f
C813 VDD1.n57 B 0.012825f
C814 VDD1.n58 B 0.013579f
C815 VDD1.n59 B 0.030313f
C816 VDD1.n60 B 0.030313f
C817 VDD1.n61 B 0.013579f
C818 VDD1.n62 B 0.012825f
C819 VDD1.n63 B 0.023866f
C820 VDD1.n64 B 0.023866f
C821 VDD1.n65 B 0.012825f
C822 VDD1.n66 B 0.013579f
C823 VDD1.n67 B 0.030313f
C824 VDD1.n68 B 0.030313f
C825 VDD1.n69 B 0.013579f
C826 VDD1.n70 B 0.012825f
C827 VDD1.n71 B 0.023866f
C828 VDD1.n72 B 0.023866f
C829 VDD1.n73 B 0.012825f
C830 VDD1.n74 B 0.013579f
C831 VDD1.n75 B 0.030313f
C832 VDD1.n76 B 0.030313f
C833 VDD1.n77 B 0.013579f
C834 VDD1.n78 B 0.012825f
C835 VDD1.n79 B 0.023866f
C836 VDD1.n80 B 0.023866f
C837 VDD1.n81 B 0.012825f
C838 VDD1.n82 B 0.013579f
C839 VDD1.n83 B 0.030313f
C840 VDD1.n84 B 0.030313f
C841 VDD1.n85 B 0.013579f
C842 VDD1.n86 B 0.012825f
C843 VDD1.n87 B 0.023866f
C844 VDD1.n88 B 0.023866f
C845 VDD1.n89 B 0.012825f
C846 VDD1.n90 B 0.013579f
C847 VDD1.n91 B 0.030313f
C848 VDD1.n92 B 0.066192f
C849 VDD1.n93 B 0.013579f
C850 VDD1.n94 B 0.012825f
C851 VDD1.n95 B 0.057122f
C852 VDD1.n96 B 0.069095f
C853 VDD1.t1 B 0.331558f
C854 VDD1.t7 B 0.331558f
C855 VDD1.n97 B 3.01877f
C856 VDD1.n98 B 0.747478f
C857 VDD1.n99 B 0.033868f
C858 VDD1.n100 B 0.023866f
C859 VDD1.n101 B 0.012825f
C860 VDD1.n102 B 0.030313f
C861 VDD1.n103 B 0.013579f
C862 VDD1.n104 B 0.023866f
C863 VDD1.n105 B 0.012825f
C864 VDD1.n106 B 0.030313f
C865 VDD1.n107 B 0.013202f
C866 VDD1.n108 B 0.023866f
C867 VDD1.n109 B 0.013579f
C868 VDD1.n110 B 0.030313f
C869 VDD1.n111 B 0.013579f
C870 VDD1.n112 B 0.023866f
C871 VDD1.n113 B 0.012825f
C872 VDD1.n114 B 0.030313f
C873 VDD1.n115 B 0.013579f
C874 VDD1.n116 B 0.023866f
C875 VDD1.n117 B 0.012825f
C876 VDD1.n118 B 0.030313f
C877 VDD1.n119 B 0.013579f
C878 VDD1.n120 B 0.023866f
C879 VDD1.n121 B 0.012825f
C880 VDD1.n122 B 0.030313f
C881 VDD1.n123 B 0.013579f
C882 VDD1.n124 B 0.023866f
C883 VDD1.n125 B 0.012825f
C884 VDD1.n126 B 0.030313f
C885 VDD1.n127 B 0.013579f
C886 VDD1.n128 B 1.83498f
C887 VDD1.n129 B 0.012825f
C888 VDD1.t9 B 0.050194f
C889 VDD1.n130 B 0.1711f
C890 VDD1.n131 B 0.017907f
C891 VDD1.n132 B 0.022735f
C892 VDD1.n133 B 0.030313f
C893 VDD1.n134 B 0.013579f
C894 VDD1.n135 B 0.012825f
C895 VDD1.n136 B 0.023866f
C896 VDD1.n137 B 0.023866f
C897 VDD1.n138 B 0.012825f
C898 VDD1.n139 B 0.013579f
C899 VDD1.n140 B 0.030313f
C900 VDD1.n141 B 0.030313f
C901 VDD1.n142 B 0.013579f
C902 VDD1.n143 B 0.012825f
C903 VDD1.n144 B 0.023866f
C904 VDD1.n145 B 0.023866f
C905 VDD1.n146 B 0.012825f
C906 VDD1.n147 B 0.013579f
C907 VDD1.n148 B 0.030313f
C908 VDD1.n149 B 0.030313f
C909 VDD1.n150 B 0.013579f
C910 VDD1.n151 B 0.012825f
C911 VDD1.n152 B 0.023866f
C912 VDD1.n153 B 0.023866f
C913 VDD1.n154 B 0.012825f
C914 VDD1.n155 B 0.013579f
C915 VDD1.n156 B 0.030313f
C916 VDD1.n157 B 0.030313f
C917 VDD1.n158 B 0.013579f
C918 VDD1.n159 B 0.012825f
C919 VDD1.n160 B 0.023866f
C920 VDD1.n161 B 0.023866f
C921 VDD1.n162 B 0.012825f
C922 VDD1.n163 B 0.013579f
C923 VDD1.n164 B 0.030313f
C924 VDD1.n165 B 0.030313f
C925 VDD1.n166 B 0.013579f
C926 VDD1.n167 B 0.012825f
C927 VDD1.n168 B 0.023866f
C928 VDD1.n169 B 0.023866f
C929 VDD1.n170 B 0.012825f
C930 VDD1.n171 B 0.012825f
C931 VDD1.n172 B 0.013579f
C932 VDD1.n173 B 0.030313f
C933 VDD1.n174 B 0.030313f
C934 VDD1.n175 B 0.030313f
C935 VDD1.n176 B 0.013202f
C936 VDD1.n177 B 0.012825f
C937 VDD1.n178 B 0.023866f
C938 VDD1.n179 B 0.023866f
C939 VDD1.n180 B 0.012825f
C940 VDD1.n181 B 0.013579f
C941 VDD1.n182 B 0.030313f
C942 VDD1.n183 B 0.030313f
C943 VDD1.n184 B 0.013579f
C944 VDD1.n185 B 0.012825f
C945 VDD1.n186 B 0.023866f
C946 VDD1.n187 B 0.023866f
C947 VDD1.n188 B 0.012825f
C948 VDD1.n189 B 0.013579f
C949 VDD1.n190 B 0.030313f
C950 VDD1.n191 B 0.066192f
C951 VDD1.n192 B 0.013579f
C952 VDD1.n193 B 0.012825f
C953 VDD1.n194 B 0.057122f
C954 VDD1.n195 B 0.069095f
C955 VDD1.t8 B 0.331558f
C956 VDD1.t2 B 0.331558f
C957 VDD1.n196 B 3.01876f
C958 VDD1.n197 B 0.73956f
C959 VDD1.t5 B 0.331558f
C960 VDD1.t3 B 0.331558f
C961 VDD1.n198 B 3.03924f
C962 VDD1.n199 B 3.50329f
C963 VDD1.t0 B 0.331558f
C964 VDD1.t4 B 0.331558f
C965 VDD1.n200 B 3.01876f
C966 VDD1.n201 B 3.63732f
C967 VP.t2 B 2.77095f
C968 VP.n0 B 1.03246f
C969 VP.n1 B 0.018375f
C970 VP.n2 B 0.022898f
C971 VP.n3 B 0.018375f
C972 VP.t8 B 2.77095f
C973 VP.n4 B 0.958322f
C974 VP.n5 B 0.018375f
C975 VP.n6 B 0.02544f
C976 VP.n7 B 0.018375f
C977 VP.t3 B 2.77095f
C978 VP.n8 B 0.034075f
C979 VP.n9 B 0.018375f
C980 VP.n10 B 0.034075f
C981 VP.n11 B 0.018375f
C982 VP.t5 B 2.77095f
C983 VP.n12 B 0.034075f
C984 VP.n13 B 0.018375f
C985 VP.n14 B 0.03071f
C986 VP.t9 B 2.77095f
C987 VP.n15 B 1.03246f
C988 VP.n16 B 0.018375f
C989 VP.n17 B 0.022898f
C990 VP.n18 B 0.018375f
C991 VP.t1 B 2.77095f
C992 VP.n19 B 0.958322f
C993 VP.n20 B 0.018375f
C994 VP.n21 B 0.02544f
C995 VP.n22 B 0.018375f
C996 VP.t6 B 2.77095f
C997 VP.n23 B 0.034075f
C998 VP.n24 B 0.018375f
C999 VP.n25 B 0.034075f
C1000 VP.t7 B 2.98617f
C1001 VP.n26 B 0.981629f
C1002 VP.t0 B 2.77095f
C1003 VP.n27 B 1.02484f
C1004 VP.n28 B 0.032393f
C1005 VP.n29 B 0.210032f
C1006 VP.n30 B 0.018375f
C1007 VP.n31 B 0.018375f
C1008 VP.n32 B 0.027982f
C1009 VP.n33 B 0.02544f
C1010 VP.n34 B 0.034075f
C1011 VP.n35 B 0.018375f
C1012 VP.n36 B 0.018375f
C1013 VP.n37 B 0.018375f
C1014 VP.n38 B 0.975575f
C1015 VP.n39 B 0.034075f
C1016 VP.n40 B 0.034075f
C1017 VP.n41 B 0.018375f
C1018 VP.n42 B 0.018375f
C1019 VP.n43 B 0.018375f
C1020 VP.n44 B 0.027982f
C1021 VP.n45 B 0.034075f
C1022 VP.n46 B 0.032393f
C1023 VP.n47 B 0.018375f
C1024 VP.n48 B 0.018375f
C1025 VP.n49 B 0.018935f
C1026 VP.n50 B 0.034075f
C1027 VP.n51 B 0.034075f
C1028 VP.n52 B 0.018375f
C1029 VP.n53 B 0.018375f
C1030 VP.n54 B 0.018375f
C1031 VP.n55 B 0.030524f
C1032 VP.n56 B 0.034075f
C1033 VP.n57 B 0.03071f
C1034 VP.n58 B 0.029652f
C1035 VP.n59 B 1.34993f
C1036 VP.t4 B 2.77095f
C1037 VP.n60 B 1.03246f
C1038 VP.n61 B 1.36091f
C1039 VP.n62 B 0.029652f
C1040 VP.n63 B 0.018375f
C1041 VP.n64 B 0.034075f
C1042 VP.n65 B 0.030524f
C1043 VP.n66 B 0.022898f
C1044 VP.n67 B 0.018375f
C1045 VP.n68 B 0.018375f
C1046 VP.n69 B 0.018375f
C1047 VP.n70 B 0.034075f
C1048 VP.n71 B 0.018935f
C1049 VP.n72 B 0.958322f
C1050 VP.n73 B 0.032393f
C1051 VP.n74 B 0.018375f
C1052 VP.n75 B 0.018375f
C1053 VP.n76 B 0.018375f
C1054 VP.n77 B 0.027982f
C1055 VP.n78 B 0.02544f
C1056 VP.n79 B 0.034075f
C1057 VP.n80 B 0.018375f
C1058 VP.n81 B 0.018375f
C1059 VP.n82 B 0.018375f
C1060 VP.n83 B 0.975575f
C1061 VP.n84 B 0.034075f
C1062 VP.n85 B 0.034075f
C1063 VP.n86 B 0.018375f
C1064 VP.n87 B 0.018375f
C1065 VP.n88 B 0.018375f
C1066 VP.n89 B 0.027982f
C1067 VP.n90 B 0.034075f
C1068 VP.n91 B 0.032393f
C1069 VP.n92 B 0.018375f
C1070 VP.n93 B 0.018375f
C1071 VP.n94 B 0.018935f
C1072 VP.n95 B 0.034075f
C1073 VP.n96 B 0.034075f
C1074 VP.n97 B 0.018375f
C1075 VP.n98 B 0.018375f
C1076 VP.n99 B 0.018375f
C1077 VP.n100 B 0.030524f
C1078 VP.n101 B 0.034075f
C1079 VP.n102 B 0.03071f
C1080 VP.n103 B 0.029652f
C1081 VP.n104 B 0.039303f
.ends

