* NGSPICE file created from diff_pair_sample_1653.ext - technology: sky130A

.subckt diff_pair_sample_1653 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t7 VN.t0 VTAIL.t12 B.t3 sky130_fd_pr__nfet_01v8 ad=0.77715 pd=5.04 as=1.8369 ps=10.2 w=4.71 l=3.19
X1 B.t21 B.t19 B.t20 B.t13 sky130_fd_pr__nfet_01v8 ad=1.8369 pd=10.2 as=0 ps=0 w=4.71 l=3.19
X2 VDD2.t6 VN.t1 VTAIL.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=0.77715 pd=5.04 as=0.77715 ps=5.04 w=4.71 l=3.19
X3 VTAIL.t15 VN.t2 VDD2.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=0.77715 pd=5.04 as=0.77715 ps=5.04 w=4.71 l=3.19
X4 VTAIL.t10 VN.t3 VDD2.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=0.77715 pd=5.04 as=0.77715 ps=5.04 w=4.71 l=3.19
X5 VTAIL.t4 VP.t0 VDD1.t7 B.t4 sky130_fd_pr__nfet_01v8 ad=0.77715 pd=5.04 as=0.77715 ps=5.04 w=4.71 l=3.19
X6 VTAIL.t11 VN.t4 VDD2.t3 B.t6 sky130_fd_pr__nfet_01v8 ad=1.8369 pd=10.2 as=0.77715 ps=5.04 w=4.71 l=3.19
X7 VTAIL.t9 VN.t5 VDD2.t2 B.t1 sky130_fd_pr__nfet_01v8 ad=1.8369 pd=10.2 as=0.77715 ps=5.04 w=4.71 l=3.19
X8 VTAIL.t6 VP.t1 VDD1.t6 B.t6 sky130_fd_pr__nfet_01v8 ad=1.8369 pd=10.2 as=0.77715 ps=5.04 w=4.71 l=3.19
X9 B.t18 B.t16 B.t17 B.t9 sky130_fd_pr__nfet_01v8 ad=1.8369 pd=10.2 as=0 ps=0 w=4.71 l=3.19
X10 VDD1.t5 VP.t2 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=0.77715 pd=5.04 as=0.77715 ps=5.04 w=4.71 l=3.19
X11 B.t15 B.t12 B.t14 B.t13 sky130_fd_pr__nfet_01v8 ad=1.8369 pd=10.2 as=0 ps=0 w=4.71 l=3.19
X12 VTAIL.t1 VP.t3 VDD1.t4 B.t1 sky130_fd_pr__nfet_01v8 ad=1.8369 pd=10.2 as=0.77715 ps=5.04 w=4.71 l=3.19
X13 VDD2.t1 VN.t6 VTAIL.t13 B.t2 sky130_fd_pr__nfet_01v8 ad=0.77715 pd=5.04 as=1.8369 ps=10.2 w=4.71 l=3.19
X14 VDD1.t3 VP.t4 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=0.77715 pd=5.04 as=1.8369 ps=10.2 w=4.71 l=3.19
X15 VDD1.t2 VP.t5 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=0.77715 pd=5.04 as=1.8369 ps=10.2 w=4.71 l=3.19
X16 VTAIL.t5 VP.t6 VDD1.t1 B.t5 sky130_fd_pr__nfet_01v8 ad=0.77715 pd=5.04 as=0.77715 ps=5.04 w=4.71 l=3.19
X17 VDD1.t0 VP.t7 VTAIL.t7 B.t7 sky130_fd_pr__nfet_01v8 ad=0.77715 pd=5.04 as=0.77715 ps=5.04 w=4.71 l=3.19
X18 VDD2.t0 VN.t7 VTAIL.t14 B.t0 sky130_fd_pr__nfet_01v8 ad=0.77715 pd=5.04 as=0.77715 ps=5.04 w=4.71 l=3.19
X19 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=1.8369 pd=10.2 as=0 ps=0 w=4.71 l=3.19
R0 VN.n64 VN.n63 161.3
R1 VN.n62 VN.n34 161.3
R2 VN.n61 VN.n60 161.3
R3 VN.n59 VN.n35 161.3
R4 VN.n58 VN.n57 161.3
R5 VN.n56 VN.n36 161.3
R6 VN.n55 VN.n54 161.3
R7 VN.n53 VN.n52 161.3
R8 VN.n51 VN.n38 161.3
R9 VN.n50 VN.n49 161.3
R10 VN.n48 VN.n39 161.3
R11 VN.n47 VN.n46 161.3
R12 VN.n45 VN.n40 161.3
R13 VN.n44 VN.n43 161.3
R14 VN.n31 VN.n30 161.3
R15 VN.n29 VN.n1 161.3
R16 VN.n28 VN.n27 161.3
R17 VN.n26 VN.n2 161.3
R18 VN.n25 VN.n24 161.3
R19 VN.n23 VN.n3 161.3
R20 VN.n22 VN.n21 161.3
R21 VN.n20 VN.n19 161.3
R22 VN.n18 VN.n5 161.3
R23 VN.n17 VN.n16 161.3
R24 VN.n15 VN.n6 161.3
R25 VN.n14 VN.n13 161.3
R26 VN.n12 VN.n7 161.3
R27 VN.n11 VN.n10 161.3
R28 VN.n32 VN.n0 76.3659
R29 VN.n65 VN.n33 76.3659
R30 VN.n42 VN.t6 68.4265
R31 VN.n9 VN.t4 68.4265
R32 VN.n9 VN.n8 61.53
R33 VN.n42 VN.n41 61.53
R34 VN VN.n65 48.3692
R35 VN.n28 VN.n2 42.4359
R36 VN.n61 VN.n35 42.4359
R37 VN.n13 VN.n6 40.4934
R38 VN.n17 VN.n6 40.4934
R39 VN.n46 VN.n39 40.4934
R40 VN.n50 VN.n39 40.4934
R41 VN.n24 VN.n2 38.5509
R42 VN.n57 VN.n35 38.5509
R43 VN.n8 VN.t1 35.5839
R44 VN.n4 VN.t3 35.5839
R45 VN.n0 VN.t0 35.5839
R46 VN.n41 VN.t2 35.5839
R47 VN.n37 VN.t7 35.5839
R48 VN.n33 VN.t5 35.5839
R49 VN.n12 VN.n11 24.4675
R50 VN.n13 VN.n12 24.4675
R51 VN.n18 VN.n17 24.4675
R52 VN.n19 VN.n18 24.4675
R53 VN.n23 VN.n22 24.4675
R54 VN.n24 VN.n23 24.4675
R55 VN.n29 VN.n28 24.4675
R56 VN.n30 VN.n29 24.4675
R57 VN.n46 VN.n45 24.4675
R58 VN.n45 VN.n44 24.4675
R59 VN.n57 VN.n56 24.4675
R60 VN.n56 VN.n55 24.4675
R61 VN.n52 VN.n51 24.4675
R62 VN.n51 VN.n50 24.4675
R63 VN.n63 VN.n62 24.4675
R64 VN.n62 VN.n61 24.4675
R65 VN.n30 VN.n0 13.702
R66 VN.n63 VN.n33 13.702
R67 VN.n11 VN.n8 12.7233
R68 VN.n19 VN.n4 12.7233
R69 VN.n44 VN.n41 12.7233
R70 VN.n52 VN.n37 12.7233
R71 VN.n22 VN.n4 11.7447
R72 VN.n55 VN.n37 11.7447
R73 VN.n43 VN.n42 4.20582
R74 VN.n10 VN.n9 4.20582
R75 VN.n65 VN.n64 0.354971
R76 VN.n32 VN.n31 0.354971
R77 VN VN.n32 0.26696
R78 VN.n64 VN.n34 0.189894
R79 VN.n60 VN.n34 0.189894
R80 VN.n60 VN.n59 0.189894
R81 VN.n59 VN.n58 0.189894
R82 VN.n58 VN.n36 0.189894
R83 VN.n54 VN.n36 0.189894
R84 VN.n54 VN.n53 0.189894
R85 VN.n53 VN.n38 0.189894
R86 VN.n49 VN.n38 0.189894
R87 VN.n49 VN.n48 0.189894
R88 VN.n48 VN.n47 0.189894
R89 VN.n47 VN.n40 0.189894
R90 VN.n43 VN.n40 0.189894
R91 VN.n10 VN.n7 0.189894
R92 VN.n14 VN.n7 0.189894
R93 VN.n15 VN.n14 0.189894
R94 VN.n16 VN.n15 0.189894
R95 VN.n16 VN.n5 0.189894
R96 VN.n20 VN.n5 0.189894
R97 VN.n21 VN.n20 0.189894
R98 VN.n21 VN.n3 0.189894
R99 VN.n25 VN.n3 0.189894
R100 VN.n26 VN.n25 0.189894
R101 VN.n27 VN.n26 0.189894
R102 VN.n27 VN.n1 0.189894
R103 VN.n31 VN.n1 0.189894
R104 VTAIL.n194 VTAIL.n176 289.615
R105 VTAIL.n20 VTAIL.n2 289.615
R106 VTAIL.n44 VTAIL.n26 289.615
R107 VTAIL.n70 VTAIL.n52 289.615
R108 VTAIL.n170 VTAIL.n152 289.615
R109 VTAIL.n144 VTAIL.n126 289.615
R110 VTAIL.n120 VTAIL.n102 289.615
R111 VTAIL.n94 VTAIL.n76 289.615
R112 VTAIL.n185 VTAIL.n184 185
R113 VTAIL.n187 VTAIL.n186 185
R114 VTAIL.n180 VTAIL.n179 185
R115 VTAIL.n193 VTAIL.n192 185
R116 VTAIL.n195 VTAIL.n194 185
R117 VTAIL.n11 VTAIL.n10 185
R118 VTAIL.n13 VTAIL.n12 185
R119 VTAIL.n6 VTAIL.n5 185
R120 VTAIL.n19 VTAIL.n18 185
R121 VTAIL.n21 VTAIL.n20 185
R122 VTAIL.n35 VTAIL.n34 185
R123 VTAIL.n37 VTAIL.n36 185
R124 VTAIL.n30 VTAIL.n29 185
R125 VTAIL.n43 VTAIL.n42 185
R126 VTAIL.n45 VTAIL.n44 185
R127 VTAIL.n61 VTAIL.n60 185
R128 VTAIL.n63 VTAIL.n62 185
R129 VTAIL.n56 VTAIL.n55 185
R130 VTAIL.n69 VTAIL.n68 185
R131 VTAIL.n71 VTAIL.n70 185
R132 VTAIL.n171 VTAIL.n170 185
R133 VTAIL.n169 VTAIL.n168 185
R134 VTAIL.n156 VTAIL.n155 185
R135 VTAIL.n163 VTAIL.n162 185
R136 VTAIL.n161 VTAIL.n160 185
R137 VTAIL.n145 VTAIL.n144 185
R138 VTAIL.n143 VTAIL.n142 185
R139 VTAIL.n130 VTAIL.n129 185
R140 VTAIL.n137 VTAIL.n136 185
R141 VTAIL.n135 VTAIL.n134 185
R142 VTAIL.n121 VTAIL.n120 185
R143 VTAIL.n119 VTAIL.n118 185
R144 VTAIL.n106 VTAIL.n105 185
R145 VTAIL.n113 VTAIL.n112 185
R146 VTAIL.n111 VTAIL.n110 185
R147 VTAIL.n95 VTAIL.n94 185
R148 VTAIL.n93 VTAIL.n92 185
R149 VTAIL.n80 VTAIL.n79 185
R150 VTAIL.n87 VTAIL.n86 185
R151 VTAIL.n85 VTAIL.n84 185
R152 VTAIL.n183 VTAIL.t12 147.714
R153 VTAIL.n9 VTAIL.t11 147.714
R154 VTAIL.n33 VTAIL.t2 147.714
R155 VTAIL.n59 VTAIL.t1 147.714
R156 VTAIL.n159 VTAIL.t3 147.714
R157 VTAIL.n133 VTAIL.t6 147.714
R158 VTAIL.n109 VTAIL.t13 147.714
R159 VTAIL.n83 VTAIL.t9 147.714
R160 VTAIL.n186 VTAIL.n185 104.615
R161 VTAIL.n186 VTAIL.n179 104.615
R162 VTAIL.n193 VTAIL.n179 104.615
R163 VTAIL.n194 VTAIL.n193 104.615
R164 VTAIL.n12 VTAIL.n11 104.615
R165 VTAIL.n12 VTAIL.n5 104.615
R166 VTAIL.n19 VTAIL.n5 104.615
R167 VTAIL.n20 VTAIL.n19 104.615
R168 VTAIL.n36 VTAIL.n35 104.615
R169 VTAIL.n36 VTAIL.n29 104.615
R170 VTAIL.n43 VTAIL.n29 104.615
R171 VTAIL.n44 VTAIL.n43 104.615
R172 VTAIL.n62 VTAIL.n61 104.615
R173 VTAIL.n62 VTAIL.n55 104.615
R174 VTAIL.n69 VTAIL.n55 104.615
R175 VTAIL.n70 VTAIL.n69 104.615
R176 VTAIL.n170 VTAIL.n169 104.615
R177 VTAIL.n169 VTAIL.n155 104.615
R178 VTAIL.n162 VTAIL.n155 104.615
R179 VTAIL.n162 VTAIL.n161 104.615
R180 VTAIL.n144 VTAIL.n143 104.615
R181 VTAIL.n143 VTAIL.n129 104.615
R182 VTAIL.n136 VTAIL.n129 104.615
R183 VTAIL.n136 VTAIL.n135 104.615
R184 VTAIL.n120 VTAIL.n119 104.615
R185 VTAIL.n119 VTAIL.n105 104.615
R186 VTAIL.n112 VTAIL.n105 104.615
R187 VTAIL.n112 VTAIL.n111 104.615
R188 VTAIL.n94 VTAIL.n93 104.615
R189 VTAIL.n93 VTAIL.n79 104.615
R190 VTAIL.n86 VTAIL.n79 104.615
R191 VTAIL.n86 VTAIL.n85 104.615
R192 VTAIL.n151 VTAIL.n150 56.8721
R193 VTAIL.n101 VTAIL.n100 56.8721
R194 VTAIL.n1 VTAIL.n0 56.8719
R195 VTAIL.n51 VTAIL.n50 56.8719
R196 VTAIL.n185 VTAIL.t12 52.3082
R197 VTAIL.n11 VTAIL.t11 52.3082
R198 VTAIL.n35 VTAIL.t2 52.3082
R199 VTAIL.n61 VTAIL.t1 52.3082
R200 VTAIL.n161 VTAIL.t3 52.3082
R201 VTAIL.n135 VTAIL.t6 52.3082
R202 VTAIL.n111 VTAIL.t13 52.3082
R203 VTAIL.n85 VTAIL.t9 52.3082
R204 VTAIL.n199 VTAIL.n198 35.0944
R205 VTAIL.n25 VTAIL.n24 35.0944
R206 VTAIL.n49 VTAIL.n48 35.0944
R207 VTAIL.n75 VTAIL.n74 35.0944
R208 VTAIL.n175 VTAIL.n174 35.0944
R209 VTAIL.n149 VTAIL.n148 35.0944
R210 VTAIL.n125 VTAIL.n124 35.0944
R211 VTAIL.n99 VTAIL.n98 35.0944
R212 VTAIL.n199 VTAIL.n175 19.4617
R213 VTAIL.n99 VTAIL.n75 19.4617
R214 VTAIL.n184 VTAIL.n183 15.6631
R215 VTAIL.n10 VTAIL.n9 15.6631
R216 VTAIL.n34 VTAIL.n33 15.6631
R217 VTAIL.n60 VTAIL.n59 15.6631
R218 VTAIL.n160 VTAIL.n159 15.6631
R219 VTAIL.n134 VTAIL.n133 15.6631
R220 VTAIL.n110 VTAIL.n109 15.6631
R221 VTAIL.n84 VTAIL.n83 15.6631
R222 VTAIL.n187 VTAIL.n182 12.8005
R223 VTAIL.n13 VTAIL.n8 12.8005
R224 VTAIL.n37 VTAIL.n32 12.8005
R225 VTAIL.n63 VTAIL.n58 12.8005
R226 VTAIL.n163 VTAIL.n158 12.8005
R227 VTAIL.n137 VTAIL.n132 12.8005
R228 VTAIL.n113 VTAIL.n108 12.8005
R229 VTAIL.n87 VTAIL.n82 12.8005
R230 VTAIL.n188 VTAIL.n180 12.0247
R231 VTAIL.n14 VTAIL.n6 12.0247
R232 VTAIL.n38 VTAIL.n30 12.0247
R233 VTAIL.n64 VTAIL.n56 12.0247
R234 VTAIL.n164 VTAIL.n156 12.0247
R235 VTAIL.n138 VTAIL.n130 12.0247
R236 VTAIL.n114 VTAIL.n106 12.0247
R237 VTAIL.n88 VTAIL.n80 12.0247
R238 VTAIL.n192 VTAIL.n191 11.249
R239 VTAIL.n18 VTAIL.n17 11.249
R240 VTAIL.n42 VTAIL.n41 11.249
R241 VTAIL.n68 VTAIL.n67 11.249
R242 VTAIL.n168 VTAIL.n167 11.249
R243 VTAIL.n142 VTAIL.n141 11.249
R244 VTAIL.n118 VTAIL.n117 11.249
R245 VTAIL.n92 VTAIL.n91 11.249
R246 VTAIL.n195 VTAIL.n178 10.4732
R247 VTAIL.n21 VTAIL.n4 10.4732
R248 VTAIL.n45 VTAIL.n28 10.4732
R249 VTAIL.n71 VTAIL.n54 10.4732
R250 VTAIL.n171 VTAIL.n154 10.4732
R251 VTAIL.n145 VTAIL.n128 10.4732
R252 VTAIL.n121 VTAIL.n104 10.4732
R253 VTAIL.n95 VTAIL.n78 10.4732
R254 VTAIL.n196 VTAIL.n176 9.69747
R255 VTAIL.n22 VTAIL.n2 9.69747
R256 VTAIL.n46 VTAIL.n26 9.69747
R257 VTAIL.n72 VTAIL.n52 9.69747
R258 VTAIL.n172 VTAIL.n152 9.69747
R259 VTAIL.n146 VTAIL.n126 9.69747
R260 VTAIL.n122 VTAIL.n102 9.69747
R261 VTAIL.n96 VTAIL.n76 9.69747
R262 VTAIL.n198 VTAIL.n197 9.45567
R263 VTAIL.n24 VTAIL.n23 9.45567
R264 VTAIL.n48 VTAIL.n47 9.45567
R265 VTAIL.n74 VTAIL.n73 9.45567
R266 VTAIL.n174 VTAIL.n173 9.45567
R267 VTAIL.n148 VTAIL.n147 9.45567
R268 VTAIL.n124 VTAIL.n123 9.45567
R269 VTAIL.n98 VTAIL.n97 9.45567
R270 VTAIL.n197 VTAIL.n196 9.3005
R271 VTAIL.n178 VTAIL.n177 9.3005
R272 VTAIL.n191 VTAIL.n190 9.3005
R273 VTAIL.n189 VTAIL.n188 9.3005
R274 VTAIL.n182 VTAIL.n181 9.3005
R275 VTAIL.n23 VTAIL.n22 9.3005
R276 VTAIL.n4 VTAIL.n3 9.3005
R277 VTAIL.n17 VTAIL.n16 9.3005
R278 VTAIL.n15 VTAIL.n14 9.3005
R279 VTAIL.n8 VTAIL.n7 9.3005
R280 VTAIL.n47 VTAIL.n46 9.3005
R281 VTAIL.n28 VTAIL.n27 9.3005
R282 VTAIL.n41 VTAIL.n40 9.3005
R283 VTAIL.n39 VTAIL.n38 9.3005
R284 VTAIL.n32 VTAIL.n31 9.3005
R285 VTAIL.n73 VTAIL.n72 9.3005
R286 VTAIL.n54 VTAIL.n53 9.3005
R287 VTAIL.n67 VTAIL.n66 9.3005
R288 VTAIL.n65 VTAIL.n64 9.3005
R289 VTAIL.n58 VTAIL.n57 9.3005
R290 VTAIL.n173 VTAIL.n172 9.3005
R291 VTAIL.n154 VTAIL.n153 9.3005
R292 VTAIL.n167 VTAIL.n166 9.3005
R293 VTAIL.n165 VTAIL.n164 9.3005
R294 VTAIL.n158 VTAIL.n157 9.3005
R295 VTAIL.n147 VTAIL.n146 9.3005
R296 VTAIL.n128 VTAIL.n127 9.3005
R297 VTAIL.n141 VTAIL.n140 9.3005
R298 VTAIL.n139 VTAIL.n138 9.3005
R299 VTAIL.n132 VTAIL.n131 9.3005
R300 VTAIL.n123 VTAIL.n122 9.3005
R301 VTAIL.n104 VTAIL.n103 9.3005
R302 VTAIL.n117 VTAIL.n116 9.3005
R303 VTAIL.n115 VTAIL.n114 9.3005
R304 VTAIL.n108 VTAIL.n107 9.3005
R305 VTAIL.n97 VTAIL.n96 9.3005
R306 VTAIL.n78 VTAIL.n77 9.3005
R307 VTAIL.n91 VTAIL.n90 9.3005
R308 VTAIL.n89 VTAIL.n88 9.3005
R309 VTAIL.n82 VTAIL.n81 9.3005
R310 VTAIL.n183 VTAIL.n181 4.39059
R311 VTAIL.n9 VTAIL.n7 4.39059
R312 VTAIL.n33 VTAIL.n31 4.39059
R313 VTAIL.n59 VTAIL.n57 4.39059
R314 VTAIL.n159 VTAIL.n157 4.39059
R315 VTAIL.n133 VTAIL.n131 4.39059
R316 VTAIL.n109 VTAIL.n107 4.39059
R317 VTAIL.n83 VTAIL.n81 4.39059
R318 VTAIL.n198 VTAIL.n176 4.26717
R319 VTAIL.n24 VTAIL.n2 4.26717
R320 VTAIL.n48 VTAIL.n26 4.26717
R321 VTAIL.n74 VTAIL.n52 4.26717
R322 VTAIL.n174 VTAIL.n152 4.26717
R323 VTAIL.n148 VTAIL.n126 4.26717
R324 VTAIL.n124 VTAIL.n102 4.26717
R325 VTAIL.n98 VTAIL.n76 4.26717
R326 VTAIL.n0 VTAIL.t8 4.20432
R327 VTAIL.n0 VTAIL.t10 4.20432
R328 VTAIL.n50 VTAIL.t0 4.20432
R329 VTAIL.n50 VTAIL.t5 4.20432
R330 VTAIL.n150 VTAIL.t7 4.20432
R331 VTAIL.n150 VTAIL.t4 4.20432
R332 VTAIL.n100 VTAIL.t14 4.20432
R333 VTAIL.n100 VTAIL.t15 4.20432
R334 VTAIL.n196 VTAIL.n195 3.49141
R335 VTAIL.n22 VTAIL.n21 3.49141
R336 VTAIL.n46 VTAIL.n45 3.49141
R337 VTAIL.n72 VTAIL.n71 3.49141
R338 VTAIL.n172 VTAIL.n171 3.49141
R339 VTAIL.n146 VTAIL.n145 3.49141
R340 VTAIL.n122 VTAIL.n121 3.49141
R341 VTAIL.n96 VTAIL.n95 3.49141
R342 VTAIL.n101 VTAIL.n99 3.03498
R343 VTAIL.n125 VTAIL.n101 3.03498
R344 VTAIL.n151 VTAIL.n149 3.03498
R345 VTAIL.n175 VTAIL.n151 3.03498
R346 VTAIL.n75 VTAIL.n51 3.03498
R347 VTAIL.n51 VTAIL.n49 3.03498
R348 VTAIL.n25 VTAIL.n1 3.03498
R349 VTAIL VTAIL.n199 2.97679
R350 VTAIL.n192 VTAIL.n178 2.71565
R351 VTAIL.n18 VTAIL.n4 2.71565
R352 VTAIL.n42 VTAIL.n28 2.71565
R353 VTAIL.n68 VTAIL.n54 2.71565
R354 VTAIL.n168 VTAIL.n154 2.71565
R355 VTAIL.n142 VTAIL.n128 2.71565
R356 VTAIL.n118 VTAIL.n104 2.71565
R357 VTAIL.n92 VTAIL.n78 2.71565
R358 VTAIL.n191 VTAIL.n180 1.93989
R359 VTAIL.n17 VTAIL.n6 1.93989
R360 VTAIL.n41 VTAIL.n30 1.93989
R361 VTAIL.n67 VTAIL.n56 1.93989
R362 VTAIL.n167 VTAIL.n156 1.93989
R363 VTAIL.n141 VTAIL.n130 1.93989
R364 VTAIL.n117 VTAIL.n106 1.93989
R365 VTAIL.n91 VTAIL.n80 1.93989
R366 VTAIL.n188 VTAIL.n187 1.16414
R367 VTAIL.n14 VTAIL.n13 1.16414
R368 VTAIL.n38 VTAIL.n37 1.16414
R369 VTAIL.n64 VTAIL.n63 1.16414
R370 VTAIL.n164 VTAIL.n163 1.16414
R371 VTAIL.n138 VTAIL.n137 1.16414
R372 VTAIL.n114 VTAIL.n113 1.16414
R373 VTAIL.n88 VTAIL.n87 1.16414
R374 VTAIL.n149 VTAIL.n125 0.470328
R375 VTAIL.n49 VTAIL.n25 0.470328
R376 VTAIL.n184 VTAIL.n182 0.388379
R377 VTAIL.n10 VTAIL.n8 0.388379
R378 VTAIL.n34 VTAIL.n32 0.388379
R379 VTAIL.n60 VTAIL.n58 0.388379
R380 VTAIL.n160 VTAIL.n158 0.388379
R381 VTAIL.n134 VTAIL.n132 0.388379
R382 VTAIL.n110 VTAIL.n108 0.388379
R383 VTAIL.n84 VTAIL.n82 0.388379
R384 VTAIL.n189 VTAIL.n181 0.155672
R385 VTAIL.n190 VTAIL.n189 0.155672
R386 VTAIL.n190 VTAIL.n177 0.155672
R387 VTAIL.n197 VTAIL.n177 0.155672
R388 VTAIL.n15 VTAIL.n7 0.155672
R389 VTAIL.n16 VTAIL.n15 0.155672
R390 VTAIL.n16 VTAIL.n3 0.155672
R391 VTAIL.n23 VTAIL.n3 0.155672
R392 VTAIL.n39 VTAIL.n31 0.155672
R393 VTAIL.n40 VTAIL.n39 0.155672
R394 VTAIL.n40 VTAIL.n27 0.155672
R395 VTAIL.n47 VTAIL.n27 0.155672
R396 VTAIL.n65 VTAIL.n57 0.155672
R397 VTAIL.n66 VTAIL.n65 0.155672
R398 VTAIL.n66 VTAIL.n53 0.155672
R399 VTAIL.n73 VTAIL.n53 0.155672
R400 VTAIL.n173 VTAIL.n153 0.155672
R401 VTAIL.n166 VTAIL.n153 0.155672
R402 VTAIL.n166 VTAIL.n165 0.155672
R403 VTAIL.n165 VTAIL.n157 0.155672
R404 VTAIL.n147 VTAIL.n127 0.155672
R405 VTAIL.n140 VTAIL.n127 0.155672
R406 VTAIL.n140 VTAIL.n139 0.155672
R407 VTAIL.n139 VTAIL.n131 0.155672
R408 VTAIL.n123 VTAIL.n103 0.155672
R409 VTAIL.n116 VTAIL.n103 0.155672
R410 VTAIL.n116 VTAIL.n115 0.155672
R411 VTAIL.n115 VTAIL.n107 0.155672
R412 VTAIL.n97 VTAIL.n77 0.155672
R413 VTAIL.n90 VTAIL.n77 0.155672
R414 VTAIL.n90 VTAIL.n89 0.155672
R415 VTAIL.n89 VTAIL.n81 0.155672
R416 VTAIL VTAIL.n1 0.0586897
R417 VDD2.n2 VDD2.n1 75.0126
R418 VDD2.n2 VDD2.n0 75.0126
R419 VDD2 VDD2.n5 75.0098
R420 VDD2.n4 VDD2.n3 73.5509
R421 VDD2.n4 VDD2.n2 41.4308
R422 VDD2.n5 VDD2.t5 4.20432
R423 VDD2.n5 VDD2.t1 4.20432
R424 VDD2.n3 VDD2.t2 4.20432
R425 VDD2.n3 VDD2.t0 4.20432
R426 VDD2.n1 VDD2.t4 4.20432
R427 VDD2.n1 VDD2.t7 4.20432
R428 VDD2.n0 VDD2.t3 4.20432
R429 VDD2.n0 VDD2.t6 4.20432
R430 VDD2 VDD2.n4 1.57593
R431 B.n742 B.n741 585
R432 B.n236 B.n135 585
R433 B.n235 B.n234 585
R434 B.n233 B.n232 585
R435 B.n231 B.n230 585
R436 B.n229 B.n228 585
R437 B.n227 B.n226 585
R438 B.n225 B.n224 585
R439 B.n223 B.n222 585
R440 B.n221 B.n220 585
R441 B.n219 B.n218 585
R442 B.n217 B.n216 585
R443 B.n215 B.n214 585
R444 B.n213 B.n212 585
R445 B.n211 B.n210 585
R446 B.n209 B.n208 585
R447 B.n207 B.n206 585
R448 B.n205 B.n204 585
R449 B.n203 B.n202 585
R450 B.n201 B.n200 585
R451 B.n199 B.n198 585
R452 B.n197 B.n196 585
R453 B.n195 B.n194 585
R454 B.n193 B.n192 585
R455 B.n191 B.n190 585
R456 B.n189 B.n188 585
R457 B.n187 B.n186 585
R458 B.n185 B.n184 585
R459 B.n183 B.n182 585
R460 B.n181 B.n180 585
R461 B.n179 B.n178 585
R462 B.n177 B.n176 585
R463 B.n175 B.n174 585
R464 B.n173 B.n172 585
R465 B.n171 B.n170 585
R466 B.n169 B.n168 585
R467 B.n167 B.n166 585
R468 B.n165 B.n164 585
R469 B.n163 B.n162 585
R470 B.n161 B.n160 585
R471 B.n159 B.n158 585
R472 B.n157 B.n156 585
R473 B.n155 B.n154 585
R474 B.n153 B.n152 585
R475 B.n151 B.n150 585
R476 B.n149 B.n148 585
R477 B.n147 B.n146 585
R478 B.n145 B.n144 585
R479 B.n143 B.n142 585
R480 B.n109 B.n108 585
R481 B.n740 B.n110 585
R482 B.n745 B.n110 585
R483 B.n739 B.n738 585
R484 B.n738 B.n106 585
R485 B.n737 B.n105 585
R486 B.n751 B.n105 585
R487 B.n736 B.n104 585
R488 B.n752 B.n104 585
R489 B.n735 B.n103 585
R490 B.n753 B.n103 585
R491 B.n734 B.n733 585
R492 B.n733 B.n99 585
R493 B.n732 B.n98 585
R494 B.n759 B.n98 585
R495 B.n731 B.n97 585
R496 B.n760 B.n97 585
R497 B.n730 B.n96 585
R498 B.n761 B.n96 585
R499 B.n729 B.n728 585
R500 B.n728 B.n92 585
R501 B.n727 B.n91 585
R502 B.n767 B.n91 585
R503 B.n726 B.n90 585
R504 B.n768 B.n90 585
R505 B.n725 B.n89 585
R506 B.n769 B.n89 585
R507 B.n724 B.n723 585
R508 B.n723 B.n85 585
R509 B.n722 B.n84 585
R510 B.n775 B.n84 585
R511 B.n721 B.n83 585
R512 B.n776 B.n83 585
R513 B.n720 B.n82 585
R514 B.n777 B.n82 585
R515 B.n719 B.n718 585
R516 B.n718 B.n78 585
R517 B.n717 B.n77 585
R518 B.n783 B.n77 585
R519 B.n716 B.n76 585
R520 B.n784 B.n76 585
R521 B.n715 B.n75 585
R522 B.n785 B.n75 585
R523 B.n714 B.n713 585
R524 B.n713 B.n71 585
R525 B.n712 B.n70 585
R526 B.n791 B.n70 585
R527 B.n711 B.n69 585
R528 B.n792 B.n69 585
R529 B.n710 B.n68 585
R530 B.n793 B.n68 585
R531 B.n709 B.n708 585
R532 B.n708 B.n64 585
R533 B.n707 B.n63 585
R534 B.n799 B.n63 585
R535 B.n706 B.n62 585
R536 B.n800 B.n62 585
R537 B.n705 B.n61 585
R538 B.n801 B.n61 585
R539 B.n704 B.n703 585
R540 B.n703 B.n57 585
R541 B.n702 B.n56 585
R542 B.n807 B.n56 585
R543 B.n701 B.n55 585
R544 B.n808 B.n55 585
R545 B.n700 B.n54 585
R546 B.n809 B.n54 585
R547 B.n699 B.n698 585
R548 B.n698 B.n50 585
R549 B.n697 B.n49 585
R550 B.n815 B.n49 585
R551 B.n696 B.n48 585
R552 B.n816 B.n48 585
R553 B.n695 B.n47 585
R554 B.n817 B.n47 585
R555 B.n694 B.n693 585
R556 B.n693 B.n43 585
R557 B.n692 B.n42 585
R558 B.n823 B.n42 585
R559 B.n691 B.n41 585
R560 B.n824 B.n41 585
R561 B.n690 B.n40 585
R562 B.n825 B.n40 585
R563 B.n689 B.n688 585
R564 B.n688 B.n36 585
R565 B.n687 B.n35 585
R566 B.n831 B.n35 585
R567 B.n686 B.n34 585
R568 B.n832 B.n34 585
R569 B.n685 B.n33 585
R570 B.n833 B.n33 585
R571 B.n684 B.n683 585
R572 B.n683 B.n29 585
R573 B.n682 B.n28 585
R574 B.n839 B.n28 585
R575 B.n681 B.n27 585
R576 B.n840 B.n27 585
R577 B.n680 B.n26 585
R578 B.n841 B.n26 585
R579 B.n679 B.n678 585
R580 B.n678 B.n22 585
R581 B.n677 B.n21 585
R582 B.n847 B.n21 585
R583 B.n676 B.n20 585
R584 B.n848 B.n20 585
R585 B.n675 B.n19 585
R586 B.n849 B.n19 585
R587 B.n674 B.n673 585
R588 B.n673 B.n18 585
R589 B.n672 B.n14 585
R590 B.n855 B.n14 585
R591 B.n671 B.n13 585
R592 B.n856 B.n13 585
R593 B.n670 B.n12 585
R594 B.n857 B.n12 585
R595 B.n669 B.n668 585
R596 B.n668 B.n8 585
R597 B.n667 B.n7 585
R598 B.n863 B.n7 585
R599 B.n666 B.n6 585
R600 B.n864 B.n6 585
R601 B.n665 B.n5 585
R602 B.n865 B.n5 585
R603 B.n664 B.n663 585
R604 B.n663 B.n4 585
R605 B.n662 B.n237 585
R606 B.n662 B.n661 585
R607 B.n652 B.n238 585
R608 B.n239 B.n238 585
R609 B.n654 B.n653 585
R610 B.n655 B.n654 585
R611 B.n651 B.n244 585
R612 B.n244 B.n243 585
R613 B.n650 B.n649 585
R614 B.n649 B.n648 585
R615 B.n246 B.n245 585
R616 B.n641 B.n246 585
R617 B.n640 B.n639 585
R618 B.n642 B.n640 585
R619 B.n638 B.n251 585
R620 B.n251 B.n250 585
R621 B.n637 B.n636 585
R622 B.n636 B.n635 585
R623 B.n253 B.n252 585
R624 B.n254 B.n253 585
R625 B.n628 B.n627 585
R626 B.n629 B.n628 585
R627 B.n626 B.n259 585
R628 B.n259 B.n258 585
R629 B.n625 B.n624 585
R630 B.n624 B.n623 585
R631 B.n261 B.n260 585
R632 B.n262 B.n261 585
R633 B.n616 B.n615 585
R634 B.n617 B.n616 585
R635 B.n614 B.n267 585
R636 B.n267 B.n266 585
R637 B.n613 B.n612 585
R638 B.n612 B.n611 585
R639 B.n269 B.n268 585
R640 B.n270 B.n269 585
R641 B.n604 B.n603 585
R642 B.n605 B.n604 585
R643 B.n602 B.n275 585
R644 B.n275 B.n274 585
R645 B.n601 B.n600 585
R646 B.n600 B.n599 585
R647 B.n277 B.n276 585
R648 B.n278 B.n277 585
R649 B.n592 B.n591 585
R650 B.n593 B.n592 585
R651 B.n590 B.n283 585
R652 B.n283 B.n282 585
R653 B.n589 B.n588 585
R654 B.n588 B.n587 585
R655 B.n285 B.n284 585
R656 B.n286 B.n285 585
R657 B.n580 B.n579 585
R658 B.n581 B.n580 585
R659 B.n578 B.n291 585
R660 B.n291 B.n290 585
R661 B.n577 B.n576 585
R662 B.n576 B.n575 585
R663 B.n293 B.n292 585
R664 B.n294 B.n293 585
R665 B.n568 B.n567 585
R666 B.n569 B.n568 585
R667 B.n566 B.n299 585
R668 B.n299 B.n298 585
R669 B.n565 B.n564 585
R670 B.n564 B.n563 585
R671 B.n301 B.n300 585
R672 B.n302 B.n301 585
R673 B.n556 B.n555 585
R674 B.n557 B.n556 585
R675 B.n554 B.n307 585
R676 B.n307 B.n306 585
R677 B.n553 B.n552 585
R678 B.n552 B.n551 585
R679 B.n309 B.n308 585
R680 B.n310 B.n309 585
R681 B.n544 B.n543 585
R682 B.n545 B.n544 585
R683 B.n542 B.n315 585
R684 B.n315 B.n314 585
R685 B.n541 B.n540 585
R686 B.n540 B.n539 585
R687 B.n317 B.n316 585
R688 B.n318 B.n317 585
R689 B.n532 B.n531 585
R690 B.n533 B.n532 585
R691 B.n530 B.n323 585
R692 B.n323 B.n322 585
R693 B.n529 B.n528 585
R694 B.n528 B.n527 585
R695 B.n325 B.n324 585
R696 B.n326 B.n325 585
R697 B.n520 B.n519 585
R698 B.n521 B.n520 585
R699 B.n518 B.n331 585
R700 B.n331 B.n330 585
R701 B.n517 B.n516 585
R702 B.n516 B.n515 585
R703 B.n333 B.n332 585
R704 B.n334 B.n333 585
R705 B.n508 B.n507 585
R706 B.n509 B.n508 585
R707 B.n506 B.n339 585
R708 B.n339 B.n338 585
R709 B.n505 B.n504 585
R710 B.n504 B.n503 585
R711 B.n341 B.n340 585
R712 B.n342 B.n341 585
R713 B.n496 B.n495 585
R714 B.n497 B.n496 585
R715 B.n494 B.n347 585
R716 B.n347 B.n346 585
R717 B.n493 B.n492 585
R718 B.n492 B.n491 585
R719 B.n349 B.n348 585
R720 B.n350 B.n349 585
R721 B.n484 B.n483 585
R722 B.n485 B.n484 585
R723 B.n353 B.n352 585
R724 B.n384 B.n382 585
R725 B.n385 B.n381 585
R726 B.n385 B.n354 585
R727 B.n388 B.n387 585
R728 B.n389 B.n380 585
R729 B.n391 B.n390 585
R730 B.n393 B.n379 585
R731 B.n396 B.n395 585
R732 B.n397 B.n378 585
R733 B.n399 B.n398 585
R734 B.n401 B.n377 585
R735 B.n404 B.n403 585
R736 B.n405 B.n376 585
R737 B.n407 B.n406 585
R738 B.n409 B.n375 585
R739 B.n412 B.n411 585
R740 B.n413 B.n374 585
R741 B.n415 B.n414 585
R742 B.n417 B.n373 585
R743 B.n420 B.n419 585
R744 B.n422 B.n370 585
R745 B.n424 B.n423 585
R746 B.n426 B.n369 585
R747 B.n429 B.n428 585
R748 B.n430 B.n368 585
R749 B.n432 B.n431 585
R750 B.n434 B.n367 585
R751 B.n437 B.n436 585
R752 B.n438 B.n366 585
R753 B.n443 B.n442 585
R754 B.n445 B.n365 585
R755 B.n448 B.n447 585
R756 B.n449 B.n364 585
R757 B.n451 B.n450 585
R758 B.n453 B.n363 585
R759 B.n456 B.n455 585
R760 B.n457 B.n362 585
R761 B.n459 B.n458 585
R762 B.n461 B.n361 585
R763 B.n464 B.n463 585
R764 B.n465 B.n360 585
R765 B.n467 B.n466 585
R766 B.n469 B.n359 585
R767 B.n472 B.n471 585
R768 B.n473 B.n358 585
R769 B.n475 B.n474 585
R770 B.n477 B.n357 585
R771 B.n478 B.n356 585
R772 B.n481 B.n480 585
R773 B.n482 B.n355 585
R774 B.n355 B.n354 585
R775 B.n487 B.n486 585
R776 B.n486 B.n485 585
R777 B.n488 B.n351 585
R778 B.n351 B.n350 585
R779 B.n490 B.n489 585
R780 B.n491 B.n490 585
R781 B.n345 B.n344 585
R782 B.n346 B.n345 585
R783 B.n499 B.n498 585
R784 B.n498 B.n497 585
R785 B.n500 B.n343 585
R786 B.n343 B.n342 585
R787 B.n502 B.n501 585
R788 B.n503 B.n502 585
R789 B.n337 B.n336 585
R790 B.n338 B.n337 585
R791 B.n511 B.n510 585
R792 B.n510 B.n509 585
R793 B.n512 B.n335 585
R794 B.n335 B.n334 585
R795 B.n514 B.n513 585
R796 B.n515 B.n514 585
R797 B.n329 B.n328 585
R798 B.n330 B.n329 585
R799 B.n523 B.n522 585
R800 B.n522 B.n521 585
R801 B.n524 B.n327 585
R802 B.n327 B.n326 585
R803 B.n526 B.n525 585
R804 B.n527 B.n526 585
R805 B.n321 B.n320 585
R806 B.n322 B.n321 585
R807 B.n535 B.n534 585
R808 B.n534 B.n533 585
R809 B.n536 B.n319 585
R810 B.n319 B.n318 585
R811 B.n538 B.n537 585
R812 B.n539 B.n538 585
R813 B.n313 B.n312 585
R814 B.n314 B.n313 585
R815 B.n547 B.n546 585
R816 B.n546 B.n545 585
R817 B.n548 B.n311 585
R818 B.n311 B.n310 585
R819 B.n550 B.n549 585
R820 B.n551 B.n550 585
R821 B.n305 B.n304 585
R822 B.n306 B.n305 585
R823 B.n559 B.n558 585
R824 B.n558 B.n557 585
R825 B.n560 B.n303 585
R826 B.n303 B.n302 585
R827 B.n562 B.n561 585
R828 B.n563 B.n562 585
R829 B.n297 B.n296 585
R830 B.n298 B.n297 585
R831 B.n571 B.n570 585
R832 B.n570 B.n569 585
R833 B.n572 B.n295 585
R834 B.n295 B.n294 585
R835 B.n574 B.n573 585
R836 B.n575 B.n574 585
R837 B.n289 B.n288 585
R838 B.n290 B.n289 585
R839 B.n583 B.n582 585
R840 B.n582 B.n581 585
R841 B.n584 B.n287 585
R842 B.n287 B.n286 585
R843 B.n586 B.n585 585
R844 B.n587 B.n586 585
R845 B.n281 B.n280 585
R846 B.n282 B.n281 585
R847 B.n595 B.n594 585
R848 B.n594 B.n593 585
R849 B.n596 B.n279 585
R850 B.n279 B.n278 585
R851 B.n598 B.n597 585
R852 B.n599 B.n598 585
R853 B.n273 B.n272 585
R854 B.n274 B.n273 585
R855 B.n607 B.n606 585
R856 B.n606 B.n605 585
R857 B.n608 B.n271 585
R858 B.n271 B.n270 585
R859 B.n610 B.n609 585
R860 B.n611 B.n610 585
R861 B.n265 B.n264 585
R862 B.n266 B.n265 585
R863 B.n619 B.n618 585
R864 B.n618 B.n617 585
R865 B.n620 B.n263 585
R866 B.n263 B.n262 585
R867 B.n622 B.n621 585
R868 B.n623 B.n622 585
R869 B.n257 B.n256 585
R870 B.n258 B.n257 585
R871 B.n631 B.n630 585
R872 B.n630 B.n629 585
R873 B.n632 B.n255 585
R874 B.n255 B.n254 585
R875 B.n634 B.n633 585
R876 B.n635 B.n634 585
R877 B.n249 B.n248 585
R878 B.n250 B.n249 585
R879 B.n644 B.n643 585
R880 B.n643 B.n642 585
R881 B.n645 B.n247 585
R882 B.n641 B.n247 585
R883 B.n647 B.n646 585
R884 B.n648 B.n647 585
R885 B.n242 B.n241 585
R886 B.n243 B.n242 585
R887 B.n657 B.n656 585
R888 B.n656 B.n655 585
R889 B.n658 B.n240 585
R890 B.n240 B.n239 585
R891 B.n660 B.n659 585
R892 B.n661 B.n660 585
R893 B.n2 B.n0 585
R894 B.n4 B.n2 585
R895 B.n3 B.n1 585
R896 B.n864 B.n3 585
R897 B.n862 B.n861 585
R898 B.n863 B.n862 585
R899 B.n860 B.n9 585
R900 B.n9 B.n8 585
R901 B.n859 B.n858 585
R902 B.n858 B.n857 585
R903 B.n11 B.n10 585
R904 B.n856 B.n11 585
R905 B.n854 B.n853 585
R906 B.n855 B.n854 585
R907 B.n852 B.n15 585
R908 B.n18 B.n15 585
R909 B.n851 B.n850 585
R910 B.n850 B.n849 585
R911 B.n17 B.n16 585
R912 B.n848 B.n17 585
R913 B.n846 B.n845 585
R914 B.n847 B.n846 585
R915 B.n844 B.n23 585
R916 B.n23 B.n22 585
R917 B.n843 B.n842 585
R918 B.n842 B.n841 585
R919 B.n25 B.n24 585
R920 B.n840 B.n25 585
R921 B.n838 B.n837 585
R922 B.n839 B.n838 585
R923 B.n836 B.n30 585
R924 B.n30 B.n29 585
R925 B.n835 B.n834 585
R926 B.n834 B.n833 585
R927 B.n32 B.n31 585
R928 B.n832 B.n32 585
R929 B.n830 B.n829 585
R930 B.n831 B.n830 585
R931 B.n828 B.n37 585
R932 B.n37 B.n36 585
R933 B.n827 B.n826 585
R934 B.n826 B.n825 585
R935 B.n39 B.n38 585
R936 B.n824 B.n39 585
R937 B.n822 B.n821 585
R938 B.n823 B.n822 585
R939 B.n820 B.n44 585
R940 B.n44 B.n43 585
R941 B.n819 B.n818 585
R942 B.n818 B.n817 585
R943 B.n46 B.n45 585
R944 B.n816 B.n46 585
R945 B.n814 B.n813 585
R946 B.n815 B.n814 585
R947 B.n812 B.n51 585
R948 B.n51 B.n50 585
R949 B.n811 B.n810 585
R950 B.n810 B.n809 585
R951 B.n53 B.n52 585
R952 B.n808 B.n53 585
R953 B.n806 B.n805 585
R954 B.n807 B.n806 585
R955 B.n804 B.n58 585
R956 B.n58 B.n57 585
R957 B.n803 B.n802 585
R958 B.n802 B.n801 585
R959 B.n60 B.n59 585
R960 B.n800 B.n60 585
R961 B.n798 B.n797 585
R962 B.n799 B.n798 585
R963 B.n796 B.n65 585
R964 B.n65 B.n64 585
R965 B.n795 B.n794 585
R966 B.n794 B.n793 585
R967 B.n67 B.n66 585
R968 B.n792 B.n67 585
R969 B.n790 B.n789 585
R970 B.n791 B.n790 585
R971 B.n788 B.n72 585
R972 B.n72 B.n71 585
R973 B.n787 B.n786 585
R974 B.n786 B.n785 585
R975 B.n74 B.n73 585
R976 B.n784 B.n74 585
R977 B.n782 B.n781 585
R978 B.n783 B.n782 585
R979 B.n780 B.n79 585
R980 B.n79 B.n78 585
R981 B.n779 B.n778 585
R982 B.n778 B.n777 585
R983 B.n81 B.n80 585
R984 B.n776 B.n81 585
R985 B.n774 B.n773 585
R986 B.n775 B.n774 585
R987 B.n772 B.n86 585
R988 B.n86 B.n85 585
R989 B.n771 B.n770 585
R990 B.n770 B.n769 585
R991 B.n88 B.n87 585
R992 B.n768 B.n88 585
R993 B.n766 B.n765 585
R994 B.n767 B.n766 585
R995 B.n764 B.n93 585
R996 B.n93 B.n92 585
R997 B.n763 B.n762 585
R998 B.n762 B.n761 585
R999 B.n95 B.n94 585
R1000 B.n760 B.n95 585
R1001 B.n758 B.n757 585
R1002 B.n759 B.n758 585
R1003 B.n756 B.n100 585
R1004 B.n100 B.n99 585
R1005 B.n755 B.n754 585
R1006 B.n754 B.n753 585
R1007 B.n102 B.n101 585
R1008 B.n752 B.n102 585
R1009 B.n750 B.n749 585
R1010 B.n751 B.n750 585
R1011 B.n748 B.n107 585
R1012 B.n107 B.n106 585
R1013 B.n747 B.n746 585
R1014 B.n746 B.n745 585
R1015 B.n867 B.n866 585
R1016 B.n866 B.n865 585
R1017 B.n486 B.n353 473.281
R1018 B.n746 B.n109 473.281
R1019 B.n484 B.n355 473.281
R1020 B.n742 B.n110 473.281
R1021 B.n744 B.n743 256.663
R1022 B.n744 B.n134 256.663
R1023 B.n744 B.n133 256.663
R1024 B.n744 B.n132 256.663
R1025 B.n744 B.n131 256.663
R1026 B.n744 B.n130 256.663
R1027 B.n744 B.n129 256.663
R1028 B.n744 B.n128 256.663
R1029 B.n744 B.n127 256.663
R1030 B.n744 B.n126 256.663
R1031 B.n744 B.n125 256.663
R1032 B.n744 B.n124 256.663
R1033 B.n744 B.n123 256.663
R1034 B.n744 B.n122 256.663
R1035 B.n744 B.n121 256.663
R1036 B.n744 B.n120 256.663
R1037 B.n744 B.n119 256.663
R1038 B.n744 B.n118 256.663
R1039 B.n744 B.n117 256.663
R1040 B.n744 B.n116 256.663
R1041 B.n744 B.n115 256.663
R1042 B.n744 B.n114 256.663
R1043 B.n744 B.n113 256.663
R1044 B.n744 B.n112 256.663
R1045 B.n744 B.n111 256.663
R1046 B.n383 B.n354 256.663
R1047 B.n386 B.n354 256.663
R1048 B.n392 B.n354 256.663
R1049 B.n394 B.n354 256.663
R1050 B.n400 B.n354 256.663
R1051 B.n402 B.n354 256.663
R1052 B.n408 B.n354 256.663
R1053 B.n410 B.n354 256.663
R1054 B.n416 B.n354 256.663
R1055 B.n418 B.n354 256.663
R1056 B.n425 B.n354 256.663
R1057 B.n427 B.n354 256.663
R1058 B.n433 B.n354 256.663
R1059 B.n435 B.n354 256.663
R1060 B.n444 B.n354 256.663
R1061 B.n446 B.n354 256.663
R1062 B.n452 B.n354 256.663
R1063 B.n454 B.n354 256.663
R1064 B.n460 B.n354 256.663
R1065 B.n462 B.n354 256.663
R1066 B.n468 B.n354 256.663
R1067 B.n470 B.n354 256.663
R1068 B.n476 B.n354 256.663
R1069 B.n479 B.n354 256.663
R1070 B.n439 B.t12 244.375
R1071 B.n371 B.t19 244.375
R1072 B.n139 B.t8 244.375
R1073 B.n136 B.t16 244.375
R1074 B.n439 B.t15 225.43
R1075 B.n136 B.t17 225.43
R1076 B.n371 B.t21 225.43
R1077 B.n139 B.t10 225.43
R1078 B.n486 B.n351 163.367
R1079 B.n490 B.n351 163.367
R1080 B.n490 B.n345 163.367
R1081 B.n498 B.n345 163.367
R1082 B.n498 B.n343 163.367
R1083 B.n502 B.n343 163.367
R1084 B.n502 B.n337 163.367
R1085 B.n510 B.n337 163.367
R1086 B.n510 B.n335 163.367
R1087 B.n514 B.n335 163.367
R1088 B.n514 B.n329 163.367
R1089 B.n522 B.n329 163.367
R1090 B.n522 B.n327 163.367
R1091 B.n526 B.n327 163.367
R1092 B.n526 B.n321 163.367
R1093 B.n534 B.n321 163.367
R1094 B.n534 B.n319 163.367
R1095 B.n538 B.n319 163.367
R1096 B.n538 B.n313 163.367
R1097 B.n546 B.n313 163.367
R1098 B.n546 B.n311 163.367
R1099 B.n550 B.n311 163.367
R1100 B.n550 B.n305 163.367
R1101 B.n558 B.n305 163.367
R1102 B.n558 B.n303 163.367
R1103 B.n562 B.n303 163.367
R1104 B.n562 B.n297 163.367
R1105 B.n570 B.n297 163.367
R1106 B.n570 B.n295 163.367
R1107 B.n574 B.n295 163.367
R1108 B.n574 B.n289 163.367
R1109 B.n582 B.n289 163.367
R1110 B.n582 B.n287 163.367
R1111 B.n586 B.n287 163.367
R1112 B.n586 B.n281 163.367
R1113 B.n594 B.n281 163.367
R1114 B.n594 B.n279 163.367
R1115 B.n598 B.n279 163.367
R1116 B.n598 B.n273 163.367
R1117 B.n606 B.n273 163.367
R1118 B.n606 B.n271 163.367
R1119 B.n610 B.n271 163.367
R1120 B.n610 B.n265 163.367
R1121 B.n618 B.n265 163.367
R1122 B.n618 B.n263 163.367
R1123 B.n622 B.n263 163.367
R1124 B.n622 B.n257 163.367
R1125 B.n630 B.n257 163.367
R1126 B.n630 B.n255 163.367
R1127 B.n634 B.n255 163.367
R1128 B.n634 B.n249 163.367
R1129 B.n643 B.n249 163.367
R1130 B.n643 B.n247 163.367
R1131 B.n647 B.n247 163.367
R1132 B.n647 B.n242 163.367
R1133 B.n656 B.n242 163.367
R1134 B.n656 B.n240 163.367
R1135 B.n660 B.n240 163.367
R1136 B.n660 B.n2 163.367
R1137 B.n866 B.n2 163.367
R1138 B.n866 B.n3 163.367
R1139 B.n862 B.n3 163.367
R1140 B.n862 B.n9 163.367
R1141 B.n858 B.n9 163.367
R1142 B.n858 B.n11 163.367
R1143 B.n854 B.n11 163.367
R1144 B.n854 B.n15 163.367
R1145 B.n850 B.n15 163.367
R1146 B.n850 B.n17 163.367
R1147 B.n846 B.n17 163.367
R1148 B.n846 B.n23 163.367
R1149 B.n842 B.n23 163.367
R1150 B.n842 B.n25 163.367
R1151 B.n838 B.n25 163.367
R1152 B.n838 B.n30 163.367
R1153 B.n834 B.n30 163.367
R1154 B.n834 B.n32 163.367
R1155 B.n830 B.n32 163.367
R1156 B.n830 B.n37 163.367
R1157 B.n826 B.n37 163.367
R1158 B.n826 B.n39 163.367
R1159 B.n822 B.n39 163.367
R1160 B.n822 B.n44 163.367
R1161 B.n818 B.n44 163.367
R1162 B.n818 B.n46 163.367
R1163 B.n814 B.n46 163.367
R1164 B.n814 B.n51 163.367
R1165 B.n810 B.n51 163.367
R1166 B.n810 B.n53 163.367
R1167 B.n806 B.n53 163.367
R1168 B.n806 B.n58 163.367
R1169 B.n802 B.n58 163.367
R1170 B.n802 B.n60 163.367
R1171 B.n798 B.n60 163.367
R1172 B.n798 B.n65 163.367
R1173 B.n794 B.n65 163.367
R1174 B.n794 B.n67 163.367
R1175 B.n790 B.n67 163.367
R1176 B.n790 B.n72 163.367
R1177 B.n786 B.n72 163.367
R1178 B.n786 B.n74 163.367
R1179 B.n782 B.n74 163.367
R1180 B.n782 B.n79 163.367
R1181 B.n778 B.n79 163.367
R1182 B.n778 B.n81 163.367
R1183 B.n774 B.n81 163.367
R1184 B.n774 B.n86 163.367
R1185 B.n770 B.n86 163.367
R1186 B.n770 B.n88 163.367
R1187 B.n766 B.n88 163.367
R1188 B.n766 B.n93 163.367
R1189 B.n762 B.n93 163.367
R1190 B.n762 B.n95 163.367
R1191 B.n758 B.n95 163.367
R1192 B.n758 B.n100 163.367
R1193 B.n754 B.n100 163.367
R1194 B.n754 B.n102 163.367
R1195 B.n750 B.n102 163.367
R1196 B.n750 B.n107 163.367
R1197 B.n746 B.n107 163.367
R1198 B.n385 B.n384 163.367
R1199 B.n387 B.n385 163.367
R1200 B.n391 B.n380 163.367
R1201 B.n395 B.n393 163.367
R1202 B.n399 B.n378 163.367
R1203 B.n403 B.n401 163.367
R1204 B.n407 B.n376 163.367
R1205 B.n411 B.n409 163.367
R1206 B.n415 B.n374 163.367
R1207 B.n419 B.n417 163.367
R1208 B.n424 B.n370 163.367
R1209 B.n428 B.n426 163.367
R1210 B.n432 B.n368 163.367
R1211 B.n436 B.n434 163.367
R1212 B.n443 B.n366 163.367
R1213 B.n447 B.n445 163.367
R1214 B.n451 B.n364 163.367
R1215 B.n455 B.n453 163.367
R1216 B.n459 B.n362 163.367
R1217 B.n463 B.n461 163.367
R1218 B.n467 B.n360 163.367
R1219 B.n471 B.n469 163.367
R1220 B.n475 B.n358 163.367
R1221 B.n478 B.n477 163.367
R1222 B.n480 B.n355 163.367
R1223 B.n484 B.n349 163.367
R1224 B.n492 B.n349 163.367
R1225 B.n492 B.n347 163.367
R1226 B.n496 B.n347 163.367
R1227 B.n496 B.n341 163.367
R1228 B.n504 B.n341 163.367
R1229 B.n504 B.n339 163.367
R1230 B.n508 B.n339 163.367
R1231 B.n508 B.n333 163.367
R1232 B.n516 B.n333 163.367
R1233 B.n516 B.n331 163.367
R1234 B.n520 B.n331 163.367
R1235 B.n520 B.n325 163.367
R1236 B.n528 B.n325 163.367
R1237 B.n528 B.n323 163.367
R1238 B.n532 B.n323 163.367
R1239 B.n532 B.n317 163.367
R1240 B.n540 B.n317 163.367
R1241 B.n540 B.n315 163.367
R1242 B.n544 B.n315 163.367
R1243 B.n544 B.n309 163.367
R1244 B.n552 B.n309 163.367
R1245 B.n552 B.n307 163.367
R1246 B.n556 B.n307 163.367
R1247 B.n556 B.n301 163.367
R1248 B.n564 B.n301 163.367
R1249 B.n564 B.n299 163.367
R1250 B.n568 B.n299 163.367
R1251 B.n568 B.n293 163.367
R1252 B.n576 B.n293 163.367
R1253 B.n576 B.n291 163.367
R1254 B.n580 B.n291 163.367
R1255 B.n580 B.n285 163.367
R1256 B.n588 B.n285 163.367
R1257 B.n588 B.n283 163.367
R1258 B.n592 B.n283 163.367
R1259 B.n592 B.n277 163.367
R1260 B.n600 B.n277 163.367
R1261 B.n600 B.n275 163.367
R1262 B.n604 B.n275 163.367
R1263 B.n604 B.n269 163.367
R1264 B.n612 B.n269 163.367
R1265 B.n612 B.n267 163.367
R1266 B.n616 B.n267 163.367
R1267 B.n616 B.n261 163.367
R1268 B.n624 B.n261 163.367
R1269 B.n624 B.n259 163.367
R1270 B.n628 B.n259 163.367
R1271 B.n628 B.n253 163.367
R1272 B.n636 B.n253 163.367
R1273 B.n636 B.n251 163.367
R1274 B.n640 B.n251 163.367
R1275 B.n640 B.n246 163.367
R1276 B.n649 B.n246 163.367
R1277 B.n649 B.n244 163.367
R1278 B.n654 B.n244 163.367
R1279 B.n654 B.n238 163.367
R1280 B.n662 B.n238 163.367
R1281 B.n663 B.n662 163.367
R1282 B.n663 B.n5 163.367
R1283 B.n6 B.n5 163.367
R1284 B.n7 B.n6 163.367
R1285 B.n668 B.n7 163.367
R1286 B.n668 B.n12 163.367
R1287 B.n13 B.n12 163.367
R1288 B.n14 B.n13 163.367
R1289 B.n673 B.n14 163.367
R1290 B.n673 B.n19 163.367
R1291 B.n20 B.n19 163.367
R1292 B.n21 B.n20 163.367
R1293 B.n678 B.n21 163.367
R1294 B.n678 B.n26 163.367
R1295 B.n27 B.n26 163.367
R1296 B.n28 B.n27 163.367
R1297 B.n683 B.n28 163.367
R1298 B.n683 B.n33 163.367
R1299 B.n34 B.n33 163.367
R1300 B.n35 B.n34 163.367
R1301 B.n688 B.n35 163.367
R1302 B.n688 B.n40 163.367
R1303 B.n41 B.n40 163.367
R1304 B.n42 B.n41 163.367
R1305 B.n693 B.n42 163.367
R1306 B.n693 B.n47 163.367
R1307 B.n48 B.n47 163.367
R1308 B.n49 B.n48 163.367
R1309 B.n698 B.n49 163.367
R1310 B.n698 B.n54 163.367
R1311 B.n55 B.n54 163.367
R1312 B.n56 B.n55 163.367
R1313 B.n703 B.n56 163.367
R1314 B.n703 B.n61 163.367
R1315 B.n62 B.n61 163.367
R1316 B.n63 B.n62 163.367
R1317 B.n708 B.n63 163.367
R1318 B.n708 B.n68 163.367
R1319 B.n69 B.n68 163.367
R1320 B.n70 B.n69 163.367
R1321 B.n713 B.n70 163.367
R1322 B.n713 B.n75 163.367
R1323 B.n76 B.n75 163.367
R1324 B.n77 B.n76 163.367
R1325 B.n718 B.n77 163.367
R1326 B.n718 B.n82 163.367
R1327 B.n83 B.n82 163.367
R1328 B.n84 B.n83 163.367
R1329 B.n723 B.n84 163.367
R1330 B.n723 B.n89 163.367
R1331 B.n90 B.n89 163.367
R1332 B.n91 B.n90 163.367
R1333 B.n728 B.n91 163.367
R1334 B.n728 B.n96 163.367
R1335 B.n97 B.n96 163.367
R1336 B.n98 B.n97 163.367
R1337 B.n733 B.n98 163.367
R1338 B.n733 B.n103 163.367
R1339 B.n104 B.n103 163.367
R1340 B.n105 B.n104 163.367
R1341 B.n738 B.n105 163.367
R1342 B.n738 B.n110 163.367
R1343 B.n144 B.n143 163.367
R1344 B.n148 B.n147 163.367
R1345 B.n152 B.n151 163.367
R1346 B.n156 B.n155 163.367
R1347 B.n160 B.n159 163.367
R1348 B.n164 B.n163 163.367
R1349 B.n168 B.n167 163.367
R1350 B.n172 B.n171 163.367
R1351 B.n176 B.n175 163.367
R1352 B.n180 B.n179 163.367
R1353 B.n184 B.n183 163.367
R1354 B.n188 B.n187 163.367
R1355 B.n192 B.n191 163.367
R1356 B.n196 B.n195 163.367
R1357 B.n200 B.n199 163.367
R1358 B.n204 B.n203 163.367
R1359 B.n208 B.n207 163.367
R1360 B.n212 B.n211 163.367
R1361 B.n216 B.n215 163.367
R1362 B.n220 B.n219 163.367
R1363 B.n224 B.n223 163.367
R1364 B.n228 B.n227 163.367
R1365 B.n232 B.n231 163.367
R1366 B.n234 B.n135 163.367
R1367 B.n440 B.t14 157.163
R1368 B.n137 B.t18 157.163
R1369 B.n372 B.t20 157.163
R1370 B.n140 B.t11 157.163
R1371 B.n485 B.n354 126.691
R1372 B.n745 B.n744 126.691
R1373 B.n485 B.n350 74.9129
R1374 B.n491 B.n350 74.9129
R1375 B.n491 B.n346 74.9129
R1376 B.n497 B.n346 74.9129
R1377 B.n497 B.n342 74.9129
R1378 B.n503 B.n342 74.9129
R1379 B.n503 B.n338 74.9129
R1380 B.n509 B.n338 74.9129
R1381 B.n515 B.n334 74.9129
R1382 B.n515 B.n330 74.9129
R1383 B.n521 B.n330 74.9129
R1384 B.n521 B.n326 74.9129
R1385 B.n527 B.n326 74.9129
R1386 B.n527 B.n322 74.9129
R1387 B.n533 B.n322 74.9129
R1388 B.n533 B.n318 74.9129
R1389 B.n539 B.n318 74.9129
R1390 B.n539 B.n314 74.9129
R1391 B.n545 B.n314 74.9129
R1392 B.n545 B.n310 74.9129
R1393 B.n551 B.n310 74.9129
R1394 B.n557 B.n306 74.9129
R1395 B.n557 B.n302 74.9129
R1396 B.n563 B.n302 74.9129
R1397 B.n563 B.n298 74.9129
R1398 B.n569 B.n298 74.9129
R1399 B.n569 B.n294 74.9129
R1400 B.n575 B.n294 74.9129
R1401 B.n575 B.n290 74.9129
R1402 B.n581 B.n290 74.9129
R1403 B.n587 B.n286 74.9129
R1404 B.n587 B.n282 74.9129
R1405 B.n593 B.n282 74.9129
R1406 B.n593 B.n278 74.9129
R1407 B.n599 B.n278 74.9129
R1408 B.n599 B.n274 74.9129
R1409 B.n605 B.n274 74.9129
R1410 B.n605 B.n270 74.9129
R1411 B.n611 B.n270 74.9129
R1412 B.n617 B.n266 74.9129
R1413 B.n617 B.n262 74.9129
R1414 B.n623 B.n262 74.9129
R1415 B.n623 B.n258 74.9129
R1416 B.n629 B.n258 74.9129
R1417 B.n629 B.n254 74.9129
R1418 B.n635 B.n254 74.9129
R1419 B.n635 B.n250 74.9129
R1420 B.n642 B.n250 74.9129
R1421 B.n642 B.n641 74.9129
R1422 B.n648 B.n243 74.9129
R1423 B.n655 B.n243 74.9129
R1424 B.n655 B.n239 74.9129
R1425 B.n661 B.n239 74.9129
R1426 B.n661 B.n4 74.9129
R1427 B.n865 B.n4 74.9129
R1428 B.n865 B.n864 74.9129
R1429 B.n864 B.n863 74.9129
R1430 B.n863 B.n8 74.9129
R1431 B.n857 B.n8 74.9129
R1432 B.n857 B.n856 74.9129
R1433 B.n856 B.n855 74.9129
R1434 B.n849 B.n18 74.9129
R1435 B.n849 B.n848 74.9129
R1436 B.n848 B.n847 74.9129
R1437 B.n847 B.n22 74.9129
R1438 B.n841 B.n22 74.9129
R1439 B.n841 B.n840 74.9129
R1440 B.n840 B.n839 74.9129
R1441 B.n839 B.n29 74.9129
R1442 B.n833 B.n29 74.9129
R1443 B.n833 B.n832 74.9129
R1444 B.n831 B.n36 74.9129
R1445 B.n825 B.n36 74.9129
R1446 B.n825 B.n824 74.9129
R1447 B.n824 B.n823 74.9129
R1448 B.n823 B.n43 74.9129
R1449 B.n817 B.n43 74.9129
R1450 B.n817 B.n816 74.9129
R1451 B.n816 B.n815 74.9129
R1452 B.n815 B.n50 74.9129
R1453 B.n809 B.n808 74.9129
R1454 B.n808 B.n807 74.9129
R1455 B.n807 B.n57 74.9129
R1456 B.n801 B.n57 74.9129
R1457 B.n801 B.n800 74.9129
R1458 B.n800 B.n799 74.9129
R1459 B.n799 B.n64 74.9129
R1460 B.n793 B.n64 74.9129
R1461 B.n793 B.n792 74.9129
R1462 B.n791 B.n71 74.9129
R1463 B.n785 B.n71 74.9129
R1464 B.n785 B.n784 74.9129
R1465 B.n784 B.n783 74.9129
R1466 B.n783 B.n78 74.9129
R1467 B.n777 B.n78 74.9129
R1468 B.n777 B.n776 74.9129
R1469 B.n776 B.n775 74.9129
R1470 B.n775 B.n85 74.9129
R1471 B.n769 B.n85 74.9129
R1472 B.n769 B.n768 74.9129
R1473 B.n768 B.n767 74.9129
R1474 B.n767 B.n92 74.9129
R1475 B.n761 B.n760 74.9129
R1476 B.n760 B.n759 74.9129
R1477 B.n759 B.n99 74.9129
R1478 B.n753 B.n99 74.9129
R1479 B.n753 B.n752 74.9129
R1480 B.n752 B.n751 74.9129
R1481 B.n751 B.n106 74.9129
R1482 B.n745 B.n106 74.9129
R1483 B.n383 B.n353 71.676
R1484 B.n387 B.n386 71.676
R1485 B.n392 B.n391 71.676
R1486 B.n395 B.n394 71.676
R1487 B.n400 B.n399 71.676
R1488 B.n403 B.n402 71.676
R1489 B.n408 B.n407 71.676
R1490 B.n411 B.n410 71.676
R1491 B.n416 B.n415 71.676
R1492 B.n419 B.n418 71.676
R1493 B.n425 B.n424 71.676
R1494 B.n428 B.n427 71.676
R1495 B.n433 B.n432 71.676
R1496 B.n436 B.n435 71.676
R1497 B.n444 B.n443 71.676
R1498 B.n447 B.n446 71.676
R1499 B.n452 B.n451 71.676
R1500 B.n455 B.n454 71.676
R1501 B.n460 B.n459 71.676
R1502 B.n463 B.n462 71.676
R1503 B.n468 B.n467 71.676
R1504 B.n471 B.n470 71.676
R1505 B.n476 B.n475 71.676
R1506 B.n479 B.n478 71.676
R1507 B.n111 B.n109 71.676
R1508 B.n144 B.n112 71.676
R1509 B.n148 B.n113 71.676
R1510 B.n152 B.n114 71.676
R1511 B.n156 B.n115 71.676
R1512 B.n160 B.n116 71.676
R1513 B.n164 B.n117 71.676
R1514 B.n168 B.n118 71.676
R1515 B.n172 B.n119 71.676
R1516 B.n176 B.n120 71.676
R1517 B.n180 B.n121 71.676
R1518 B.n184 B.n122 71.676
R1519 B.n188 B.n123 71.676
R1520 B.n192 B.n124 71.676
R1521 B.n196 B.n125 71.676
R1522 B.n200 B.n126 71.676
R1523 B.n204 B.n127 71.676
R1524 B.n208 B.n128 71.676
R1525 B.n212 B.n129 71.676
R1526 B.n216 B.n130 71.676
R1527 B.n220 B.n131 71.676
R1528 B.n224 B.n132 71.676
R1529 B.n228 B.n133 71.676
R1530 B.n232 B.n134 71.676
R1531 B.n743 B.n135 71.676
R1532 B.n743 B.n742 71.676
R1533 B.n234 B.n134 71.676
R1534 B.n231 B.n133 71.676
R1535 B.n227 B.n132 71.676
R1536 B.n223 B.n131 71.676
R1537 B.n219 B.n130 71.676
R1538 B.n215 B.n129 71.676
R1539 B.n211 B.n128 71.676
R1540 B.n207 B.n127 71.676
R1541 B.n203 B.n126 71.676
R1542 B.n199 B.n125 71.676
R1543 B.n195 B.n124 71.676
R1544 B.n191 B.n123 71.676
R1545 B.n187 B.n122 71.676
R1546 B.n183 B.n121 71.676
R1547 B.n179 B.n120 71.676
R1548 B.n175 B.n119 71.676
R1549 B.n171 B.n118 71.676
R1550 B.n167 B.n117 71.676
R1551 B.n163 B.n116 71.676
R1552 B.n159 B.n115 71.676
R1553 B.n155 B.n114 71.676
R1554 B.n151 B.n113 71.676
R1555 B.n147 B.n112 71.676
R1556 B.n143 B.n111 71.676
R1557 B.n384 B.n383 71.676
R1558 B.n386 B.n380 71.676
R1559 B.n393 B.n392 71.676
R1560 B.n394 B.n378 71.676
R1561 B.n401 B.n400 71.676
R1562 B.n402 B.n376 71.676
R1563 B.n409 B.n408 71.676
R1564 B.n410 B.n374 71.676
R1565 B.n417 B.n416 71.676
R1566 B.n418 B.n370 71.676
R1567 B.n426 B.n425 71.676
R1568 B.n427 B.n368 71.676
R1569 B.n434 B.n433 71.676
R1570 B.n435 B.n366 71.676
R1571 B.n445 B.n444 71.676
R1572 B.n446 B.n364 71.676
R1573 B.n453 B.n452 71.676
R1574 B.n454 B.n362 71.676
R1575 B.n461 B.n460 71.676
R1576 B.n462 B.n360 71.676
R1577 B.n469 B.n468 71.676
R1578 B.n470 B.n358 71.676
R1579 B.n477 B.n476 71.676
R1580 B.n480 B.n479 71.676
R1581 B.n440 B.n439 68.2672
R1582 B.n372 B.n371 68.2672
R1583 B.n140 B.n139 68.2672
R1584 B.n137 B.n136 68.2672
R1585 B.n611 B.t5 64.998
R1586 B.t7 B.n831 64.998
R1587 B.t1 B.n306 62.7947
R1588 B.n792 B.t3 62.7947
R1589 B.n441 B.n440 59.5399
R1590 B.n421 B.n372 59.5399
R1591 B.n141 B.n140 59.5399
R1592 B.n138 B.n137 59.5399
R1593 B.n648 B.t2 58.3881
R1594 B.n855 B.t6 58.3881
R1595 B.n509 B.t13 45.1683
R1596 B.n761 B.t9 45.1683
R1597 B.n581 B.t0 38.5583
R1598 B.n809 B.t4 38.5583
R1599 B.t0 B.n286 36.355
R1600 B.t4 B.n50 36.355
R1601 B.n747 B.n108 30.7517
R1602 B.n741 B.n740 30.7517
R1603 B.n483 B.n482 30.7517
R1604 B.n487 B.n352 30.7517
R1605 B.t13 B.n334 29.7451
R1606 B.t9 B.n92 29.7451
R1607 B B.n867 18.0485
R1608 B.n641 B.t2 16.5253
R1609 B.n18 B.t6 16.5253
R1610 B.n551 B.t1 12.1187
R1611 B.t3 B.n791 12.1187
R1612 B.n142 B.n108 10.6151
R1613 B.n145 B.n142 10.6151
R1614 B.n146 B.n145 10.6151
R1615 B.n149 B.n146 10.6151
R1616 B.n150 B.n149 10.6151
R1617 B.n153 B.n150 10.6151
R1618 B.n154 B.n153 10.6151
R1619 B.n157 B.n154 10.6151
R1620 B.n158 B.n157 10.6151
R1621 B.n161 B.n158 10.6151
R1622 B.n162 B.n161 10.6151
R1623 B.n165 B.n162 10.6151
R1624 B.n166 B.n165 10.6151
R1625 B.n169 B.n166 10.6151
R1626 B.n170 B.n169 10.6151
R1627 B.n173 B.n170 10.6151
R1628 B.n174 B.n173 10.6151
R1629 B.n177 B.n174 10.6151
R1630 B.n178 B.n177 10.6151
R1631 B.n182 B.n181 10.6151
R1632 B.n185 B.n182 10.6151
R1633 B.n186 B.n185 10.6151
R1634 B.n189 B.n186 10.6151
R1635 B.n190 B.n189 10.6151
R1636 B.n193 B.n190 10.6151
R1637 B.n194 B.n193 10.6151
R1638 B.n197 B.n194 10.6151
R1639 B.n198 B.n197 10.6151
R1640 B.n202 B.n201 10.6151
R1641 B.n205 B.n202 10.6151
R1642 B.n206 B.n205 10.6151
R1643 B.n209 B.n206 10.6151
R1644 B.n210 B.n209 10.6151
R1645 B.n213 B.n210 10.6151
R1646 B.n214 B.n213 10.6151
R1647 B.n217 B.n214 10.6151
R1648 B.n218 B.n217 10.6151
R1649 B.n221 B.n218 10.6151
R1650 B.n222 B.n221 10.6151
R1651 B.n225 B.n222 10.6151
R1652 B.n226 B.n225 10.6151
R1653 B.n229 B.n226 10.6151
R1654 B.n230 B.n229 10.6151
R1655 B.n233 B.n230 10.6151
R1656 B.n235 B.n233 10.6151
R1657 B.n236 B.n235 10.6151
R1658 B.n741 B.n236 10.6151
R1659 B.n483 B.n348 10.6151
R1660 B.n493 B.n348 10.6151
R1661 B.n494 B.n493 10.6151
R1662 B.n495 B.n494 10.6151
R1663 B.n495 B.n340 10.6151
R1664 B.n505 B.n340 10.6151
R1665 B.n506 B.n505 10.6151
R1666 B.n507 B.n506 10.6151
R1667 B.n507 B.n332 10.6151
R1668 B.n517 B.n332 10.6151
R1669 B.n518 B.n517 10.6151
R1670 B.n519 B.n518 10.6151
R1671 B.n519 B.n324 10.6151
R1672 B.n529 B.n324 10.6151
R1673 B.n530 B.n529 10.6151
R1674 B.n531 B.n530 10.6151
R1675 B.n531 B.n316 10.6151
R1676 B.n541 B.n316 10.6151
R1677 B.n542 B.n541 10.6151
R1678 B.n543 B.n542 10.6151
R1679 B.n543 B.n308 10.6151
R1680 B.n553 B.n308 10.6151
R1681 B.n554 B.n553 10.6151
R1682 B.n555 B.n554 10.6151
R1683 B.n555 B.n300 10.6151
R1684 B.n565 B.n300 10.6151
R1685 B.n566 B.n565 10.6151
R1686 B.n567 B.n566 10.6151
R1687 B.n567 B.n292 10.6151
R1688 B.n577 B.n292 10.6151
R1689 B.n578 B.n577 10.6151
R1690 B.n579 B.n578 10.6151
R1691 B.n579 B.n284 10.6151
R1692 B.n589 B.n284 10.6151
R1693 B.n590 B.n589 10.6151
R1694 B.n591 B.n590 10.6151
R1695 B.n591 B.n276 10.6151
R1696 B.n601 B.n276 10.6151
R1697 B.n602 B.n601 10.6151
R1698 B.n603 B.n602 10.6151
R1699 B.n603 B.n268 10.6151
R1700 B.n613 B.n268 10.6151
R1701 B.n614 B.n613 10.6151
R1702 B.n615 B.n614 10.6151
R1703 B.n615 B.n260 10.6151
R1704 B.n625 B.n260 10.6151
R1705 B.n626 B.n625 10.6151
R1706 B.n627 B.n626 10.6151
R1707 B.n627 B.n252 10.6151
R1708 B.n637 B.n252 10.6151
R1709 B.n638 B.n637 10.6151
R1710 B.n639 B.n638 10.6151
R1711 B.n639 B.n245 10.6151
R1712 B.n650 B.n245 10.6151
R1713 B.n651 B.n650 10.6151
R1714 B.n653 B.n651 10.6151
R1715 B.n653 B.n652 10.6151
R1716 B.n652 B.n237 10.6151
R1717 B.n664 B.n237 10.6151
R1718 B.n665 B.n664 10.6151
R1719 B.n666 B.n665 10.6151
R1720 B.n667 B.n666 10.6151
R1721 B.n669 B.n667 10.6151
R1722 B.n670 B.n669 10.6151
R1723 B.n671 B.n670 10.6151
R1724 B.n672 B.n671 10.6151
R1725 B.n674 B.n672 10.6151
R1726 B.n675 B.n674 10.6151
R1727 B.n676 B.n675 10.6151
R1728 B.n677 B.n676 10.6151
R1729 B.n679 B.n677 10.6151
R1730 B.n680 B.n679 10.6151
R1731 B.n681 B.n680 10.6151
R1732 B.n682 B.n681 10.6151
R1733 B.n684 B.n682 10.6151
R1734 B.n685 B.n684 10.6151
R1735 B.n686 B.n685 10.6151
R1736 B.n687 B.n686 10.6151
R1737 B.n689 B.n687 10.6151
R1738 B.n690 B.n689 10.6151
R1739 B.n691 B.n690 10.6151
R1740 B.n692 B.n691 10.6151
R1741 B.n694 B.n692 10.6151
R1742 B.n695 B.n694 10.6151
R1743 B.n696 B.n695 10.6151
R1744 B.n697 B.n696 10.6151
R1745 B.n699 B.n697 10.6151
R1746 B.n700 B.n699 10.6151
R1747 B.n701 B.n700 10.6151
R1748 B.n702 B.n701 10.6151
R1749 B.n704 B.n702 10.6151
R1750 B.n705 B.n704 10.6151
R1751 B.n706 B.n705 10.6151
R1752 B.n707 B.n706 10.6151
R1753 B.n709 B.n707 10.6151
R1754 B.n710 B.n709 10.6151
R1755 B.n711 B.n710 10.6151
R1756 B.n712 B.n711 10.6151
R1757 B.n714 B.n712 10.6151
R1758 B.n715 B.n714 10.6151
R1759 B.n716 B.n715 10.6151
R1760 B.n717 B.n716 10.6151
R1761 B.n719 B.n717 10.6151
R1762 B.n720 B.n719 10.6151
R1763 B.n721 B.n720 10.6151
R1764 B.n722 B.n721 10.6151
R1765 B.n724 B.n722 10.6151
R1766 B.n725 B.n724 10.6151
R1767 B.n726 B.n725 10.6151
R1768 B.n727 B.n726 10.6151
R1769 B.n729 B.n727 10.6151
R1770 B.n730 B.n729 10.6151
R1771 B.n731 B.n730 10.6151
R1772 B.n732 B.n731 10.6151
R1773 B.n734 B.n732 10.6151
R1774 B.n735 B.n734 10.6151
R1775 B.n736 B.n735 10.6151
R1776 B.n737 B.n736 10.6151
R1777 B.n739 B.n737 10.6151
R1778 B.n740 B.n739 10.6151
R1779 B.n382 B.n352 10.6151
R1780 B.n382 B.n381 10.6151
R1781 B.n388 B.n381 10.6151
R1782 B.n389 B.n388 10.6151
R1783 B.n390 B.n389 10.6151
R1784 B.n390 B.n379 10.6151
R1785 B.n396 B.n379 10.6151
R1786 B.n397 B.n396 10.6151
R1787 B.n398 B.n397 10.6151
R1788 B.n398 B.n377 10.6151
R1789 B.n404 B.n377 10.6151
R1790 B.n405 B.n404 10.6151
R1791 B.n406 B.n405 10.6151
R1792 B.n406 B.n375 10.6151
R1793 B.n412 B.n375 10.6151
R1794 B.n413 B.n412 10.6151
R1795 B.n414 B.n413 10.6151
R1796 B.n414 B.n373 10.6151
R1797 B.n420 B.n373 10.6151
R1798 B.n423 B.n422 10.6151
R1799 B.n423 B.n369 10.6151
R1800 B.n429 B.n369 10.6151
R1801 B.n430 B.n429 10.6151
R1802 B.n431 B.n430 10.6151
R1803 B.n431 B.n367 10.6151
R1804 B.n437 B.n367 10.6151
R1805 B.n438 B.n437 10.6151
R1806 B.n442 B.n438 10.6151
R1807 B.n448 B.n365 10.6151
R1808 B.n449 B.n448 10.6151
R1809 B.n450 B.n449 10.6151
R1810 B.n450 B.n363 10.6151
R1811 B.n456 B.n363 10.6151
R1812 B.n457 B.n456 10.6151
R1813 B.n458 B.n457 10.6151
R1814 B.n458 B.n361 10.6151
R1815 B.n464 B.n361 10.6151
R1816 B.n465 B.n464 10.6151
R1817 B.n466 B.n465 10.6151
R1818 B.n466 B.n359 10.6151
R1819 B.n472 B.n359 10.6151
R1820 B.n473 B.n472 10.6151
R1821 B.n474 B.n473 10.6151
R1822 B.n474 B.n357 10.6151
R1823 B.n357 B.n356 10.6151
R1824 B.n481 B.n356 10.6151
R1825 B.n482 B.n481 10.6151
R1826 B.n488 B.n487 10.6151
R1827 B.n489 B.n488 10.6151
R1828 B.n489 B.n344 10.6151
R1829 B.n499 B.n344 10.6151
R1830 B.n500 B.n499 10.6151
R1831 B.n501 B.n500 10.6151
R1832 B.n501 B.n336 10.6151
R1833 B.n511 B.n336 10.6151
R1834 B.n512 B.n511 10.6151
R1835 B.n513 B.n512 10.6151
R1836 B.n513 B.n328 10.6151
R1837 B.n523 B.n328 10.6151
R1838 B.n524 B.n523 10.6151
R1839 B.n525 B.n524 10.6151
R1840 B.n525 B.n320 10.6151
R1841 B.n535 B.n320 10.6151
R1842 B.n536 B.n535 10.6151
R1843 B.n537 B.n536 10.6151
R1844 B.n537 B.n312 10.6151
R1845 B.n547 B.n312 10.6151
R1846 B.n548 B.n547 10.6151
R1847 B.n549 B.n548 10.6151
R1848 B.n549 B.n304 10.6151
R1849 B.n559 B.n304 10.6151
R1850 B.n560 B.n559 10.6151
R1851 B.n561 B.n560 10.6151
R1852 B.n561 B.n296 10.6151
R1853 B.n571 B.n296 10.6151
R1854 B.n572 B.n571 10.6151
R1855 B.n573 B.n572 10.6151
R1856 B.n573 B.n288 10.6151
R1857 B.n583 B.n288 10.6151
R1858 B.n584 B.n583 10.6151
R1859 B.n585 B.n584 10.6151
R1860 B.n585 B.n280 10.6151
R1861 B.n595 B.n280 10.6151
R1862 B.n596 B.n595 10.6151
R1863 B.n597 B.n596 10.6151
R1864 B.n597 B.n272 10.6151
R1865 B.n607 B.n272 10.6151
R1866 B.n608 B.n607 10.6151
R1867 B.n609 B.n608 10.6151
R1868 B.n609 B.n264 10.6151
R1869 B.n619 B.n264 10.6151
R1870 B.n620 B.n619 10.6151
R1871 B.n621 B.n620 10.6151
R1872 B.n621 B.n256 10.6151
R1873 B.n631 B.n256 10.6151
R1874 B.n632 B.n631 10.6151
R1875 B.n633 B.n632 10.6151
R1876 B.n633 B.n248 10.6151
R1877 B.n644 B.n248 10.6151
R1878 B.n645 B.n644 10.6151
R1879 B.n646 B.n645 10.6151
R1880 B.n646 B.n241 10.6151
R1881 B.n657 B.n241 10.6151
R1882 B.n658 B.n657 10.6151
R1883 B.n659 B.n658 10.6151
R1884 B.n659 B.n0 10.6151
R1885 B.n861 B.n1 10.6151
R1886 B.n861 B.n860 10.6151
R1887 B.n860 B.n859 10.6151
R1888 B.n859 B.n10 10.6151
R1889 B.n853 B.n10 10.6151
R1890 B.n853 B.n852 10.6151
R1891 B.n852 B.n851 10.6151
R1892 B.n851 B.n16 10.6151
R1893 B.n845 B.n16 10.6151
R1894 B.n845 B.n844 10.6151
R1895 B.n844 B.n843 10.6151
R1896 B.n843 B.n24 10.6151
R1897 B.n837 B.n24 10.6151
R1898 B.n837 B.n836 10.6151
R1899 B.n836 B.n835 10.6151
R1900 B.n835 B.n31 10.6151
R1901 B.n829 B.n31 10.6151
R1902 B.n829 B.n828 10.6151
R1903 B.n828 B.n827 10.6151
R1904 B.n827 B.n38 10.6151
R1905 B.n821 B.n38 10.6151
R1906 B.n821 B.n820 10.6151
R1907 B.n820 B.n819 10.6151
R1908 B.n819 B.n45 10.6151
R1909 B.n813 B.n45 10.6151
R1910 B.n813 B.n812 10.6151
R1911 B.n812 B.n811 10.6151
R1912 B.n811 B.n52 10.6151
R1913 B.n805 B.n52 10.6151
R1914 B.n805 B.n804 10.6151
R1915 B.n804 B.n803 10.6151
R1916 B.n803 B.n59 10.6151
R1917 B.n797 B.n59 10.6151
R1918 B.n797 B.n796 10.6151
R1919 B.n796 B.n795 10.6151
R1920 B.n795 B.n66 10.6151
R1921 B.n789 B.n66 10.6151
R1922 B.n789 B.n788 10.6151
R1923 B.n788 B.n787 10.6151
R1924 B.n787 B.n73 10.6151
R1925 B.n781 B.n73 10.6151
R1926 B.n781 B.n780 10.6151
R1927 B.n780 B.n779 10.6151
R1928 B.n779 B.n80 10.6151
R1929 B.n773 B.n80 10.6151
R1930 B.n773 B.n772 10.6151
R1931 B.n772 B.n771 10.6151
R1932 B.n771 B.n87 10.6151
R1933 B.n765 B.n87 10.6151
R1934 B.n765 B.n764 10.6151
R1935 B.n764 B.n763 10.6151
R1936 B.n763 B.n94 10.6151
R1937 B.n757 B.n94 10.6151
R1938 B.n757 B.n756 10.6151
R1939 B.n756 B.n755 10.6151
R1940 B.n755 B.n101 10.6151
R1941 B.n749 B.n101 10.6151
R1942 B.n749 B.n748 10.6151
R1943 B.n748 B.n747 10.6151
R1944 B.t5 B.n266 9.91537
R1945 B.n832 B.t7 9.91537
R1946 B.n178 B.n141 9.36635
R1947 B.n201 B.n138 9.36635
R1948 B.n421 B.n420 9.36635
R1949 B.n441 B.n365 9.36635
R1950 B.n867 B.n0 2.81026
R1951 B.n867 B.n1 2.81026
R1952 B.n181 B.n141 1.24928
R1953 B.n198 B.n138 1.24928
R1954 B.n422 B.n421 1.24928
R1955 B.n442 B.n441 1.24928
R1956 VP.n24 VP.n23 161.3
R1957 VP.n25 VP.n20 161.3
R1958 VP.n27 VP.n26 161.3
R1959 VP.n28 VP.n19 161.3
R1960 VP.n30 VP.n29 161.3
R1961 VP.n31 VP.n18 161.3
R1962 VP.n33 VP.n32 161.3
R1963 VP.n35 VP.n34 161.3
R1964 VP.n36 VP.n16 161.3
R1965 VP.n38 VP.n37 161.3
R1966 VP.n39 VP.n15 161.3
R1967 VP.n41 VP.n40 161.3
R1968 VP.n42 VP.n14 161.3
R1969 VP.n44 VP.n43 161.3
R1970 VP.n79 VP.n78 161.3
R1971 VP.n77 VP.n1 161.3
R1972 VP.n76 VP.n75 161.3
R1973 VP.n74 VP.n2 161.3
R1974 VP.n73 VP.n72 161.3
R1975 VP.n71 VP.n3 161.3
R1976 VP.n70 VP.n69 161.3
R1977 VP.n68 VP.n67 161.3
R1978 VP.n66 VP.n5 161.3
R1979 VP.n65 VP.n64 161.3
R1980 VP.n63 VP.n6 161.3
R1981 VP.n62 VP.n61 161.3
R1982 VP.n60 VP.n7 161.3
R1983 VP.n59 VP.n58 161.3
R1984 VP.n57 VP.n56 161.3
R1985 VP.n55 VP.n9 161.3
R1986 VP.n54 VP.n53 161.3
R1987 VP.n52 VP.n10 161.3
R1988 VP.n51 VP.n50 161.3
R1989 VP.n49 VP.n11 161.3
R1990 VP.n48 VP.n47 161.3
R1991 VP.n46 VP.n12 76.3659
R1992 VP.n80 VP.n0 76.3659
R1993 VP.n45 VP.n13 76.3659
R1994 VP.n22 VP.t1 68.4263
R1995 VP.n22 VP.n21 61.5301
R1996 VP.n46 VP.n45 48.2039
R1997 VP.n50 VP.n10 42.4359
R1998 VP.n76 VP.n2 42.4359
R1999 VP.n41 VP.n15 42.4359
R2000 VP.n61 VP.n6 40.4934
R2001 VP.n65 VP.n6 40.4934
R2002 VP.n30 VP.n19 40.4934
R2003 VP.n26 VP.n19 40.4934
R2004 VP.n54 VP.n10 38.5509
R2005 VP.n72 VP.n2 38.5509
R2006 VP.n37 VP.n15 38.5509
R2007 VP.n12 VP.t3 35.5839
R2008 VP.n8 VP.t2 35.5839
R2009 VP.n4 VP.t6 35.5839
R2010 VP.n0 VP.t4 35.5839
R2011 VP.n13 VP.t5 35.5839
R2012 VP.n17 VP.t0 35.5839
R2013 VP.n21 VP.t7 35.5839
R2014 VP.n49 VP.n48 24.4675
R2015 VP.n50 VP.n49 24.4675
R2016 VP.n55 VP.n54 24.4675
R2017 VP.n56 VP.n55 24.4675
R2018 VP.n60 VP.n59 24.4675
R2019 VP.n61 VP.n60 24.4675
R2020 VP.n66 VP.n65 24.4675
R2021 VP.n67 VP.n66 24.4675
R2022 VP.n71 VP.n70 24.4675
R2023 VP.n72 VP.n71 24.4675
R2024 VP.n77 VP.n76 24.4675
R2025 VP.n78 VP.n77 24.4675
R2026 VP.n42 VP.n41 24.4675
R2027 VP.n43 VP.n42 24.4675
R2028 VP.n31 VP.n30 24.4675
R2029 VP.n32 VP.n31 24.4675
R2030 VP.n36 VP.n35 24.4675
R2031 VP.n37 VP.n36 24.4675
R2032 VP.n25 VP.n24 24.4675
R2033 VP.n26 VP.n25 24.4675
R2034 VP.n48 VP.n12 13.702
R2035 VP.n78 VP.n0 13.702
R2036 VP.n43 VP.n13 13.702
R2037 VP.n59 VP.n8 12.7233
R2038 VP.n67 VP.n4 12.7233
R2039 VP.n32 VP.n17 12.7233
R2040 VP.n24 VP.n21 12.7233
R2041 VP.n56 VP.n8 11.7447
R2042 VP.n70 VP.n4 11.7447
R2043 VP.n35 VP.n17 11.7447
R2044 VP.n23 VP.n22 4.2058
R2045 VP.n45 VP.n44 0.354971
R2046 VP.n47 VP.n46 0.354971
R2047 VP.n80 VP.n79 0.354971
R2048 VP VP.n80 0.26696
R2049 VP.n23 VP.n20 0.189894
R2050 VP.n27 VP.n20 0.189894
R2051 VP.n28 VP.n27 0.189894
R2052 VP.n29 VP.n28 0.189894
R2053 VP.n29 VP.n18 0.189894
R2054 VP.n33 VP.n18 0.189894
R2055 VP.n34 VP.n33 0.189894
R2056 VP.n34 VP.n16 0.189894
R2057 VP.n38 VP.n16 0.189894
R2058 VP.n39 VP.n38 0.189894
R2059 VP.n40 VP.n39 0.189894
R2060 VP.n40 VP.n14 0.189894
R2061 VP.n44 VP.n14 0.189894
R2062 VP.n47 VP.n11 0.189894
R2063 VP.n51 VP.n11 0.189894
R2064 VP.n52 VP.n51 0.189894
R2065 VP.n53 VP.n52 0.189894
R2066 VP.n53 VP.n9 0.189894
R2067 VP.n57 VP.n9 0.189894
R2068 VP.n58 VP.n57 0.189894
R2069 VP.n58 VP.n7 0.189894
R2070 VP.n62 VP.n7 0.189894
R2071 VP.n63 VP.n62 0.189894
R2072 VP.n64 VP.n63 0.189894
R2073 VP.n64 VP.n5 0.189894
R2074 VP.n68 VP.n5 0.189894
R2075 VP.n69 VP.n68 0.189894
R2076 VP.n69 VP.n3 0.189894
R2077 VP.n73 VP.n3 0.189894
R2078 VP.n74 VP.n73 0.189894
R2079 VP.n75 VP.n74 0.189894
R2080 VP.n75 VP.n1 0.189894
R2081 VP.n79 VP.n1 0.189894
R2082 VDD1 VDD1.n0 75.1263
R2083 VDD1.n3 VDD1.n2 75.0126
R2084 VDD1.n3 VDD1.n1 75.0126
R2085 VDD1.n5 VDD1.n4 73.5507
R2086 VDD1.n5 VDD1.n3 42.0138
R2087 VDD1.n4 VDD1.t7 4.20432
R2088 VDD1.n4 VDD1.t2 4.20432
R2089 VDD1.n0 VDD1.t6 4.20432
R2090 VDD1.n0 VDD1.t0 4.20432
R2091 VDD1.n2 VDD1.t1 4.20432
R2092 VDD1.n2 VDD1.t3 4.20432
R2093 VDD1.n1 VDD1.t4 4.20432
R2094 VDD1.n1 VDD1.t5 4.20432
R2095 VDD1 VDD1.n5 1.45955
C0 VDD1 VP 4.26037f
C1 VDD2 VDD1 2.08194f
C2 VN VP 7.03765f
C3 VDD2 VN 3.83254f
C4 VDD2 VP 0.586513f
C5 VTAIL VDD1 6.07094f
C6 VTAIL VN 4.98653f
C7 VTAIL VP 5.00064f
C8 VDD2 VTAIL 6.12931f
C9 VN VDD1 0.156305f
C10 VDD2 B 5.481031f
C11 VDD1 B 6.002371f
C12 VTAIL B 6.031063f
C13 VN B 17.076471f
C14 VP B 15.687818f
C15 VDD1.t6 B 0.111624f
C16 VDD1.t0 B 0.111624f
C17 VDD1.n0 B 0.915394f
C18 VDD1.t4 B 0.111624f
C19 VDD1.t5 B 0.111624f
C20 VDD1.n1 B 0.914155f
C21 VDD1.t1 B 0.111624f
C22 VDD1.t3 B 0.111624f
C23 VDD1.n2 B 0.914155f
C24 VDD1.n3 B 3.84971f
C25 VDD1.t7 B 0.111624f
C26 VDD1.t2 B 0.111624f
C27 VDD1.n4 B 0.900811f
C28 VDD1.n5 B 3.13894f
C29 VP.t4 B 0.941428f
C30 VP.n0 B 0.450224f
C31 VP.n1 B 0.024061f
C32 VP.n2 B 0.019575f
C33 VP.n3 B 0.024061f
C34 VP.t6 B 0.941428f
C35 VP.n4 B 0.359849f
C36 VP.n5 B 0.024061f
C37 VP.n6 B 0.019451f
C38 VP.n7 B 0.024061f
C39 VP.t2 B 0.941428f
C40 VP.n8 B 0.359849f
C41 VP.n9 B 0.024061f
C42 VP.n10 B 0.019575f
C43 VP.n11 B 0.024061f
C44 VP.t3 B 0.941428f
C45 VP.n12 B 0.450224f
C46 VP.t5 B 0.941428f
C47 VP.n13 B 0.450224f
C48 VP.n14 B 0.024061f
C49 VP.n15 B 0.019575f
C50 VP.n16 B 0.024061f
C51 VP.t0 B 0.941428f
C52 VP.n17 B 0.359849f
C53 VP.n18 B 0.024061f
C54 VP.n19 B 0.019451f
C55 VP.n20 B 0.024061f
C56 VP.t7 B 0.941428f
C57 VP.n21 B 0.439327f
C58 VP.t1 B 1.19472f
C59 VP.n22 B 0.421995f
C60 VP.n23 B 0.279873f
C61 VP.n24 B 0.034217f
C62 VP.n25 B 0.044843f
C63 VP.n26 B 0.047821f
C64 VP.n27 B 0.024061f
C65 VP.n28 B 0.024061f
C66 VP.n29 B 0.024061f
C67 VP.n30 B 0.047821f
C68 VP.n31 B 0.044843f
C69 VP.n32 B 0.034217f
C70 VP.n33 B 0.024061f
C71 VP.n34 B 0.024061f
C72 VP.n35 B 0.033331f
C73 VP.n36 B 0.044843f
C74 VP.n37 B 0.048239f
C75 VP.n38 B 0.024061f
C76 VP.n39 B 0.024061f
C77 VP.n40 B 0.024061f
C78 VP.n41 B 0.047279f
C79 VP.n42 B 0.044843f
C80 VP.n43 B 0.035102f
C81 VP.n44 B 0.038834f
C82 VP.n45 B 1.29676f
C83 VP.n46 B 1.3147f
C84 VP.n47 B 0.038834f
C85 VP.n48 B 0.035102f
C86 VP.n49 B 0.044843f
C87 VP.n50 B 0.047279f
C88 VP.n51 B 0.024061f
C89 VP.n52 B 0.024061f
C90 VP.n53 B 0.024061f
C91 VP.n54 B 0.048239f
C92 VP.n55 B 0.044843f
C93 VP.n56 B 0.033331f
C94 VP.n57 B 0.024061f
C95 VP.n58 B 0.024061f
C96 VP.n59 B 0.034217f
C97 VP.n60 B 0.044843f
C98 VP.n61 B 0.047821f
C99 VP.n62 B 0.024061f
C100 VP.n63 B 0.024061f
C101 VP.n64 B 0.024061f
C102 VP.n65 B 0.047821f
C103 VP.n66 B 0.044843f
C104 VP.n67 B 0.034217f
C105 VP.n68 B 0.024061f
C106 VP.n69 B 0.024061f
C107 VP.n70 B 0.033331f
C108 VP.n71 B 0.044843f
C109 VP.n72 B 0.048239f
C110 VP.n73 B 0.024061f
C111 VP.n74 B 0.024061f
C112 VP.n75 B 0.024061f
C113 VP.n76 B 0.047279f
C114 VP.n77 B 0.044843f
C115 VP.n78 B 0.035102f
C116 VP.n79 B 0.038834f
C117 VP.n80 B 0.058029f
C118 VDD2.t3 B 0.108117f
C119 VDD2.t6 B 0.108117f
C120 VDD2.n0 B 0.885435f
C121 VDD2.t4 B 0.108117f
C122 VDD2.t7 B 0.108117f
C123 VDD2.n1 B 0.885435f
C124 VDD2.n2 B 3.66841f
C125 VDD2.t2 B 0.108117f
C126 VDD2.t0 B 0.108117f
C127 VDD2.n3 B 0.872515f
C128 VDD2.n4 B 3.00428f
C129 VDD2.t5 B 0.108117f
C130 VDD2.t1 B 0.108117f
C131 VDD2.n5 B 0.885396f
C132 VTAIL.t8 B 0.09625f
C133 VTAIL.t10 B 0.09625f
C134 VTAIL.n0 B 0.718099f
C135 VTAIL.n1 B 0.486093f
C136 VTAIL.n2 B 0.03757f
C137 VTAIL.n3 B 0.02586f
C138 VTAIL.n4 B 0.013896f
C139 VTAIL.n5 B 0.032845f
C140 VTAIL.n6 B 0.014713f
C141 VTAIL.n7 B 0.460643f
C142 VTAIL.n8 B 0.013896f
C143 VTAIL.t11 B 0.054042f
C144 VTAIL.n9 B 0.103477f
C145 VTAIL.n10 B 0.019383f
C146 VTAIL.n11 B 0.024634f
C147 VTAIL.n12 B 0.032845f
C148 VTAIL.n13 B 0.014713f
C149 VTAIL.n14 B 0.013896f
C150 VTAIL.n15 B 0.02586f
C151 VTAIL.n16 B 0.02586f
C152 VTAIL.n17 B 0.013896f
C153 VTAIL.n18 B 0.014713f
C154 VTAIL.n19 B 0.032845f
C155 VTAIL.n20 B 0.073264f
C156 VTAIL.n21 B 0.014713f
C157 VTAIL.n22 B 0.013896f
C158 VTAIL.n23 B 0.065073f
C159 VTAIL.n24 B 0.041373f
C160 VTAIL.n25 B 0.317086f
C161 VTAIL.n26 B 0.03757f
C162 VTAIL.n27 B 0.02586f
C163 VTAIL.n28 B 0.013896f
C164 VTAIL.n29 B 0.032845f
C165 VTAIL.n30 B 0.014713f
C166 VTAIL.n31 B 0.460643f
C167 VTAIL.n32 B 0.013896f
C168 VTAIL.t2 B 0.054042f
C169 VTAIL.n33 B 0.103477f
C170 VTAIL.n34 B 0.019383f
C171 VTAIL.n35 B 0.024634f
C172 VTAIL.n36 B 0.032845f
C173 VTAIL.n37 B 0.014713f
C174 VTAIL.n38 B 0.013896f
C175 VTAIL.n39 B 0.02586f
C176 VTAIL.n40 B 0.02586f
C177 VTAIL.n41 B 0.013896f
C178 VTAIL.n42 B 0.014713f
C179 VTAIL.n43 B 0.032845f
C180 VTAIL.n44 B 0.073264f
C181 VTAIL.n45 B 0.014713f
C182 VTAIL.n46 B 0.013896f
C183 VTAIL.n47 B 0.065073f
C184 VTAIL.n48 B 0.041373f
C185 VTAIL.n49 B 0.317086f
C186 VTAIL.t0 B 0.09625f
C187 VTAIL.t5 B 0.09625f
C188 VTAIL.n50 B 0.718099f
C189 VTAIL.n51 B 0.734097f
C190 VTAIL.n52 B 0.03757f
C191 VTAIL.n53 B 0.02586f
C192 VTAIL.n54 B 0.013896f
C193 VTAIL.n55 B 0.032845f
C194 VTAIL.n56 B 0.014713f
C195 VTAIL.n57 B 0.460643f
C196 VTAIL.n58 B 0.013896f
C197 VTAIL.t1 B 0.054042f
C198 VTAIL.n59 B 0.103477f
C199 VTAIL.n60 B 0.019383f
C200 VTAIL.n61 B 0.024634f
C201 VTAIL.n62 B 0.032845f
C202 VTAIL.n63 B 0.014713f
C203 VTAIL.n64 B 0.013896f
C204 VTAIL.n65 B 0.02586f
C205 VTAIL.n66 B 0.02586f
C206 VTAIL.n67 B 0.013896f
C207 VTAIL.n68 B 0.014713f
C208 VTAIL.n69 B 0.032845f
C209 VTAIL.n70 B 0.073264f
C210 VTAIL.n71 B 0.014713f
C211 VTAIL.n72 B 0.013896f
C212 VTAIL.n73 B 0.065073f
C213 VTAIL.n74 B 0.041373f
C214 VTAIL.n75 B 1.2204f
C215 VTAIL.n76 B 0.03757f
C216 VTAIL.n77 B 0.02586f
C217 VTAIL.n78 B 0.013896f
C218 VTAIL.n79 B 0.032845f
C219 VTAIL.n80 B 0.014713f
C220 VTAIL.n81 B 0.460643f
C221 VTAIL.n82 B 0.013896f
C222 VTAIL.t9 B 0.054042f
C223 VTAIL.n83 B 0.103477f
C224 VTAIL.n84 B 0.019383f
C225 VTAIL.n85 B 0.024634f
C226 VTAIL.n86 B 0.032845f
C227 VTAIL.n87 B 0.014713f
C228 VTAIL.n88 B 0.013896f
C229 VTAIL.n89 B 0.02586f
C230 VTAIL.n90 B 0.02586f
C231 VTAIL.n91 B 0.013896f
C232 VTAIL.n92 B 0.014713f
C233 VTAIL.n93 B 0.032845f
C234 VTAIL.n94 B 0.073264f
C235 VTAIL.n95 B 0.014713f
C236 VTAIL.n96 B 0.013896f
C237 VTAIL.n97 B 0.065073f
C238 VTAIL.n98 B 0.041373f
C239 VTAIL.n99 B 1.2204f
C240 VTAIL.t14 B 0.09625f
C241 VTAIL.t15 B 0.09625f
C242 VTAIL.n100 B 0.718104f
C243 VTAIL.n101 B 0.734092f
C244 VTAIL.n102 B 0.03757f
C245 VTAIL.n103 B 0.02586f
C246 VTAIL.n104 B 0.013896f
C247 VTAIL.n105 B 0.032845f
C248 VTAIL.n106 B 0.014713f
C249 VTAIL.n107 B 0.460643f
C250 VTAIL.n108 B 0.013896f
C251 VTAIL.t13 B 0.054042f
C252 VTAIL.n109 B 0.103477f
C253 VTAIL.n110 B 0.019383f
C254 VTAIL.n111 B 0.024634f
C255 VTAIL.n112 B 0.032845f
C256 VTAIL.n113 B 0.014713f
C257 VTAIL.n114 B 0.013896f
C258 VTAIL.n115 B 0.02586f
C259 VTAIL.n116 B 0.02586f
C260 VTAIL.n117 B 0.013896f
C261 VTAIL.n118 B 0.014713f
C262 VTAIL.n119 B 0.032845f
C263 VTAIL.n120 B 0.073264f
C264 VTAIL.n121 B 0.014713f
C265 VTAIL.n122 B 0.013896f
C266 VTAIL.n123 B 0.065073f
C267 VTAIL.n124 B 0.041373f
C268 VTAIL.n125 B 0.317086f
C269 VTAIL.n126 B 0.03757f
C270 VTAIL.n127 B 0.02586f
C271 VTAIL.n128 B 0.013896f
C272 VTAIL.n129 B 0.032845f
C273 VTAIL.n130 B 0.014713f
C274 VTAIL.n131 B 0.460643f
C275 VTAIL.n132 B 0.013896f
C276 VTAIL.t6 B 0.054042f
C277 VTAIL.n133 B 0.103477f
C278 VTAIL.n134 B 0.019383f
C279 VTAIL.n135 B 0.024634f
C280 VTAIL.n136 B 0.032845f
C281 VTAIL.n137 B 0.014713f
C282 VTAIL.n138 B 0.013896f
C283 VTAIL.n139 B 0.02586f
C284 VTAIL.n140 B 0.02586f
C285 VTAIL.n141 B 0.013896f
C286 VTAIL.n142 B 0.014713f
C287 VTAIL.n143 B 0.032845f
C288 VTAIL.n144 B 0.073264f
C289 VTAIL.n145 B 0.014713f
C290 VTAIL.n146 B 0.013896f
C291 VTAIL.n147 B 0.065073f
C292 VTAIL.n148 B 0.041373f
C293 VTAIL.n149 B 0.317086f
C294 VTAIL.t7 B 0.09625f
C295 VTAIL.t4 B 0.09625f
C296 VTAIL.n150 B 0.718104f
C297 VTAIL.n151 B 0.734092f
C298 VTAIL.n152 B 0.03757f
C299 VTAIL.n153 B 0.02586f
C300 VTAIL.n154 B 0.013896f
C301 VTAIL.n155 B 0.032845f
C302 VTAIL.n156 B 0.014713f
C303 VTAIL.n157 B 0.460643f
C304 VTAIL.n158 B 0.013896f
C305 VTAIL.t3 B 0.054042f
C306 VTAIL.n159 B 0.103477f
C307 VTAIL.n160 B 0.019383f
C308 VTAIL.n161 B 0.024634f
C309 VTAIL.n162 B 0.032845f
C310 VTAIL.n163 B 0.014713f
C311 VTAIL.n164 B 0.013896f
C312 VTAIL.n165 B 0.02586f
C313 VTAIL.n166 B 0.02586f
C314 VTAIL.n167 B 0.013896f
C315 VTAIL.n168 B 0.014713f
C316 VTAIL.n169 B 0.032845f
C317 VTAIL.n170 B 0.073264f
C318 VTAIL.n171 B 0.014713f
C319 VTAIL.n172 B 0.013896f
C320 VTAIL.n173 B 0.065073f
C321 VTAIL.n174 B 0.041373f
C322 VTAIL.n175 B 1.2204f
C323 VTAIL.n176 B 0.03757f
C324 VTAIL.n177 B 0.02586f
C325 VTAIL.n178 B 0.013896f
C326 VTAIL.n179 B 0.032845f
C327 VTAIL.n180 B 0.014713f
C328 VTAIL.n181 B 0.460643f
C329 VTAIL.n182 B 0.013896f
C330 VTAIL.t12 B 0.054042f
C331 VTAIL.n183 B 0.103477f
C332 VTAIL.n184 B 0.019383f
C333 VTAIL.n185 B 0.024634f
C334 VTAIL.n186 B 0.032845f
C335 VTAIL.n187 B 0.014713f
C336 VTAIL.n188 B 0.013896f
C337 VTAIL.n189 B 0.02586f
C338 VTAIL.n190 B 0.02586f
C339 VTAIL.n191 B 0.013896f
C340 VTAIL.n192 B 0.014713f
C341 VTAIL.n193 B 0.032845f
C342 VTAIL.n194 B 0.073264f
C343 VTAIL.n195 B 0.014713f
C344 VTAIL.n196 B 0.013896f
C345 VTAIL.n197 B 0.065073f
C346 VTAIL.n198 B 0.041373f
C347 VTAIL.n199 B 1.21555f
C348 VN.t0 B 0.910661f
C349 VN.n0 B 0.43551f
C350 VN.n1 B 0.023275f
C351 VN.n2 B 0.018935f
C352 VN.n3 B 0.023275f
C353 VN.t3 B 0.910661f
C354 VN.n4 B 0.348089f
C355 VN.n5 B 0.023275f
C356 VN.n6 B 0.018815f
C357 VN.n7 B 0.023275f
C358 VN.t1 B 0.910661f
C359 VN.n8 B 0.424969f
C360 VN.t4 B 1.15568f
C361 VN.n9 B 0.408203f
C362 VN.n10 B 0.270726f
C363 VN.n11 B 0.033098f
C364 VN.n12 B 0.043378f
C365 VN.n13 B 0.046258f
C366 VN.n14 B 0.023275f
C367 VN.n15 B 0.023275f
C368 VN.n16 B 0.023275f
C369 VN.n17 B 0.046258f
C370 VN.n18 B 0.043378f
C371 VN.n19 B 0.033098f
C372 VN.n20 B 0.023275f
C373 VN.n21 B 0.023275f
C374 VN.n22 B 0.032242f
C375 VN.n23 B 0.043378f
C376 VN.n24 B 0.046662f
C377 VN.n25 B 0.023275f
C378 VN.n26 B 0.023275f
C379 VN.n27 B 0.023275f
C380 VN.n28 B 0.045734f
C381 VN.n29 B 0.043378f
C382 VN.n30 B 0.033955f
C383 VN.n31 B 0.037565f
C384 VN.n32 B 0.056132f
C385 VN.t5 B 0.910661f
C386 VN.n33 B 0.43551f
C387 VN.n34 B 0.023275f
C388 VN.n35 B 0.018935f
C389 VN.n36 B 0.023275f
C390 VN.t7 B 0.910661f
C391 VN.n37 B 0.348089f
C392 VN.n38 B 0.023275f
C393 VN.n39 B 0.018815f
C394 VN.n40 B 0.023275f
C395 VN.t2 B 0.910661f
C396 VN.n41 B 0.424969f
C397 VN.t6 B 1.15568f
C398 VN.n42 B 0.408203f
C399 VN.n43 B 0.270726f
C400 VN.n44 B 0.033098f
C401 VN.n45 B 0.043378f
C402 VN.n46 B 0.046258f
C403 VN.n47 B 0.023275f
C404 VN.n48 B 0.023275f
C405 VN.n49 B 0.023275f
C406 VN.n50 B 0.046258f
C407 VN.n51 B 0.043378f
C408 VN.n52 B 0.033098f
C409 VN.n53 B 0.023275f
C410 VN.n54 B 0.023275f
C411 VN.n55 B 0.032242f
C412 VN.n56 B 0.043378f
C413 VN.n57 B 0.046662f
C414 VN.n58 B 0.023275f
C415 VN.n59 B 0.023275f
C416 VN.n60 B 0.023275f
C417 VN.n61 B 0.045734f
C418 VN.n62 B 0.043378f
C419 VN.n63 B 0.033955f
C420 VN.n64 B 0.037565f
C421 VN.n65 B 1.26403f
.ends

