* NGSPICE file created from diff_pair_sample_0454.ext - technology: sky130A

.subckt diff_pair_sample_0454 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t5 VN.t0 VDD2.t3 B.t0 sky130_fd_pr__nfet_01v8 ad=5.2026 pd=27.46 as=2.2011 ps=13.67 w=13.34 l=2.82
X1 VDD1.t3 VP.t0 VTAIL.t7 B.t3 sky130_fd_pr__nfet_01v8 ad=2.2011 pd=13.67 as=5.2026 ps=27.46 w=13.34 l=2.82
X2 B.t17 B.t15 B.t16 B.t9 sky130_fd_pr__nfet_01v8 ad=5.2026 pd=27.46 as=0 ps=0 w=13.34 l=2.82
X3 VTAIL.t6 VP.t1 VDD1.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=5.2026 pd=27.46 as=2.2011 ps=13.67 w=13.34 l=2.82
X4 VDD2.t0 VN.t1 VTAIL.t4 B.t1 sky130_fd_pr__nfet_01v8 ad=2.2011 pd=13.67 as=5.2026 ps=27.46 w=13.34 l=2.82
X5 B.t14 B.t12 B.t13 B.t5 sky130_fd_pr__nfet_01v8 ad=5.2026 pd=27.46 as=0 ps=0 w=13.34 l=2.82
X6 VDD2.t2 VN.t2 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=2.2011 pd=13.67 as=5.2026 ps=27.46 w=13.34 l=2.82
X7 VTAIL.t2 VN.t3 VDD2.t1 B.t2 sky130_fd_pr__nfet_01v8 ad=5.2026 pd=27.46 as=2.2011 ps=13.67 w=13.34 l=2.82
X8 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=5.2026 pd=27.46 as=0 ps=0 w=13.34 l=2.82
X9 VDD1.t1 VP.t2 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=2.2011 pd=13.67 as=5.2026 ps=27.46 w=13.34 l=2.82
X10 VTAIL.t0 VP.t3 VDD1.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=5.2026 pd=27.46 as=2.2011 ps=13.67 w=13.34 l=2.82
X11 B.t7 B.t4 B.t6 B.t5 sky130_fd_pr__nfet_01v8 ad=5.2026 pd=27.46 as=0 ps=0 w=13.34 l=2.82
R0 VN.n0 VN.t3 149.218
R1 VN.n1 VN.t2 149.218
R2 VN.n0 VN.t1 148.325
R3 VN.n1 VN.t0 148.325
R4 VN VN.n1 51.7366
R5 VN VN.n0 3.46761
R6 VDD2.n2 VDD2.n0 107.195
R7 VDD2.n2 VDD2.n1 63.8346
R8 VDD2.n1 VDD2.t3 1.48476
R9 VDD2.n1 VDD2.t2 1.48476
R10 VDD2.n0 VDD2.t1 1.48476
R11 VDD2.n0 VDD2.t0 1.48476
R12 VDD2 VDD2.n2 0.0586897
R13 VTAIL.n570 VTAIL.n504 214.453
R14 VTAIL.n66 VTAIL.n0 214.453
R15 VTAIL.n138 VTAIL.n72 214.453
R16 VTAIL.n210 VTAIL.n144 214.453
R17 VTAIL.n498 VTAIL.n432 214.453
R18 VTAIL.n426 VTAIL.n360 214.453
R19 VTAIL.n354 VTAIL.n288 214.453
R20 VTAIL.n282 VTAIL.n216 214.453
R21 VTAIL.n529 VTAIL.n528 185
R22 VTAIL.n531 VTAIL.n530 185
R23 VTAIL.n524 VTAIL.n523 185
R24 VTAIL.n537 VTAIL.n536 185
R25 VTAIL.n539 VTAIL.n538 185
R26 VTAIL.n520 VTAIL.n519 185
R27 VTAIL.n545 VTAIL.n544 185
R28 VTAIL.n547 VTAIL.n546 185
R29 VTAIL.n516 VTAIL.n515 185
R30 VTAIL.n553 VTAIL.n552 185
R31 VTAIL.n555 VTAIL.n554 185
R32 VTAIL.n512 VTAIL.n511 185
R33 VTAIL.n561 VTAIL.n560 185
R34 VTAIL.n563 VTAIL.n562 185
R35 VTAIL.n508 VTAIL.n507 185
R36 VTAIL.n569 VTAIL.n568 185
R37 VTAIL.n571 VTAIL.n570 185
R38 VTAIL.n25 VTAIL.n24 185
R39 VTAIL.n27 VTAIL.n26 185
R40 VTAIL.n20 VTAIL.n19 185
R41 VTAIL.n33 VTAIL.n32 185
R42 VTAIL.n35 VTAIL.n34 185
R43 VTAIL.n16 VTAIL.n15 185
R44 VTAIL.n41 VTAIL.n40 185
R45 VTAIL.n43 VTAIL.n42 185
R46 VTAIL.n12 VTAIL.n11 185
R47 VTAIL.n49 VTAIL.n48 185
R48 VTAIL.n51 VTAIL.n50 185
R49 VTAIL.n8 VTAIL.n7 185
R50 VTAIL.n57 VTAIL.n56 185
R51 VTAIL.n59 VTAIL.n58 185
R52 VTAIL.n4 VTAIL.n3 185
R53 VTAIL.n65 VTAIL.n64 185
R54 VTAIL.n67 VTAIL.n66 185
R55 VTAIL.n97 VTAIL.n96 185
R56 VTAIL.n99 VTAIL.n98 185
R57 VTAIL.n92 VTAIL.n91 185
R58 VTAIL.n105 VTAIL.n104 185
R59 VTAIL.n107 VTAIL.n106 185
R60 VTAIL.n88 VTAIL.n87 185
R61 VTAIL.n113 VTAIL.n112 185
R62 VTAIL.n115 VTAIL.n114 185
R63 VTAIL.n84 VTAIL.n83 185
R64 VTAIL.n121 VTAIL.n120 185
R65 VTAIL.n123 VTAIL.n122 185
R66 VTAIL.n80 VTAIL.n79 185
R67 VTAIL.n129 VTAIL.n128 185
R68 VTAIL.n131 VTAIL.n130 185
R69 VTAIL.n76 VTAIL.n75 185
R70 VTAIL.n137 VTAIL.n136 185
R71 VTAIL.n139 VTAIL.n138 185
R72 VTAIL.n169 VTAIL.n168 185
R73 VTAIL.n171 VTAIL.n170 185
R74 VTAIL.n164 VTAIL.n163 185
R75 VTAIL.n177 VTAIL.n176 185
R76 VTAIL.n179 VTAIL.n178 185
R77 VTAIL.n160 VTAIL.n159 185
R78 VTAIL.n185 VTAIL.n184 185
R79 VTAIL.n187 VTAIL.n186 185
R80 VTAIL.n156 VTAIL.n155 185
R81 VTAIL.n193 VTAIL.n192 185
R82 VTAIL.n195 VTAIL.n194 185
R83 VTAIL.n152 VTAIL.n151 185
R84 VTAIL.n201 VTAIL.n200 185
R85 VTAIL.n203 VTAIL.n202 185
R86 VTAIL.n148 VTAIL.n147 185
R87 VTAIL.n209 VTAIL.n208 185
R88 VTAIL.n211 VTAIL.n210 185
R89 VTAIL.n499 VTAIL.n498 185
R90 VTAIL.n497 VTAIL.n496 185
R91 VTAIL.n436 VTAIL.n435 185
R92 VTAIL.n491 VTAIL.n490 185
R93 VTAIL.n489 VTAIL.n488 185
R94 VTAIL.n440 VTAIL.n439 185
R95 VTAIL.n483 VTAIL.n482 185
R96 VTAIL.n481 VTAIL.n480 185
R97 VTAIL.n444 VTAIL.n443 185
R98 VTAIL.n475 VTAIL.n474 185
R99 VTAIL.n473 VTAIL.n472 185
R100 VTAIL.n448 VTAIL.n447 185
R101 VTAIL.n467 VTAIL.n466 185
R102 VTAIL.n465 VTAIL.n464 185
R103 VTAIL.n452 VTAIL.n451 185
R104 VTAIL.n459 VTAIL.n458 185
R105 VTAIL.n457 VTAIL.n456 185
R106 VTAIL.n427 VTAIL.n426 185
R107 VTAIL.n425 VTAIL.n424 185
R108 VTAIL.n364 VTAIL.n363 185
R109 VTAIL.n419 VTAIL.n418 185
R110 VTAIL.n417 VTAIL.n416 185
R111 VTAIL.n368 VTAIL.n367 185
R112 VTAIL.n411 VTAIL.n410 185
R113 VTAIL.n409 VTAIL.n408 185
R114 VTAIL.n372 VTAIL.n371 185
R115 VTAIL.n403 VTAIL.n402 185
R116 VTAIL.n401 VTAIL.n400 185
R117 VTAIL.n376 VTAIL.n375 185
R118 VTAIL.n395 VTAIL.n394 185
R119 VTAIL.n393 VTAIL.n392 185
R120 VTAIL.n380 VTAIL.n379 185
R121 VTAIL.n387 VTAIL.n386 185
R122 VTAIL.n385 VTAIL.n384 185
R123 VTAIL.n355 VTAIL.n354 185
R124 VTAIL.n353 VTAIL.n352 185
R125 VTAIL.n292 VTAIL.n291 185
R126 VTAIL.n347 VTAIL.n346 185
R127 VTAIL.n345 VTAIL.n344 185
R128 VTAIL.n296 VTAIL.n295 185
R129 VTAIL.n339 VTAIL.n338 185
R130 VTAIL.n337 VTAIL.n336 185
R131 VTAIL.n300 VTAIL.n299 185
R132 VTAIL.n331 VTAIL.n330 185
R133 VTAIL.n329 VTAIL.n328 185
R134 VTAIL.n304 VTAIL.n303 185
R135 VTAIL.n323 VTAIL.n322 185
R136 VTAIL.n321 VTAIL.n320 185
R137 VTAIL.n308 VTAIL.n307 185
R138 VTAIL.n315 VTAIL.n314 185
R139 VTAIL.n313 VTAIL.n312 185
R140 VTAIL.n283 VTAIL.n282 185
R141 VTAIL.n281 VTAIL.n280 185
R142 VTAIL.n220 VTAIL.n219 185
R143 VTAIL.n275 VTAIL.n274 185
R144 VTAIL.n273 VTAIL.n272 185
R145 VTAIL.n224 VTAIL.n223 185
R146 VTAIL.n267 VTAIL.n266 185
R147 VTAIL.n265 VTAIL.n264 185
R148 VTAIL.n228 VTAIL.n227 185
R149 VTAIL.n259 VTAIL.n258 185
R150 VTAIL.n257 VTAIL.n256 185
R151 VTAIL.n232 VTAIL.n231 185
R152 VTAIL.n251 VTAIL.n250 185
R153 VTAIL.n249 VTAIL.n248 185
R154 VTAIL.n236 VTAIL.n235 185
R155 VTAIL.n243 VTAIL.n242 185
R156 VTAIL.n241 VTAIL.n240 185
R157 VTAIL.n527 VTAIL.t4 147.659
R158 VTAIL.n23 VTAIL.t2 147.659
R159 VTAIL.n95 VTAIL.t7 147.659
R160 VTAIL.n167 VTAIL.t0 147.659
R161 VTAIL.n455 VTAIL.t1 147.659
R162 VTAIL.n383 VTAIL.t6 147.659
R163 VTAIL.n311 VTAIL.t3 147.659
R164 VTAIL.n239 VTAIL.t5 147.659
R165 VTAIL.n530 VTAIL.n529 104.615
R166 VTAIL.n530 VTAIL.n523 104.615
R167 VTAIL.n537 VTAIL.n523 104.615
R168 VTAIL.n538 VTAIL.n537 104.615
R169 VTAIL.n538 VTAIL.n519 104.615
R170 VTAIL.n545 VTAIL.n519 104.615
R171 VTAIL.n546 VTAIL.n545 104.615
R172 VTAIL.n546 VTAIL.n515 104.615
R173 VTAIL.n553 VTAIL.n515 104.615
R174 VTAIL.n554 VTAIL.n553 104.615
R175 VTAIL.n554 VTAIL.n511 104.615
R176 VTAIL.n561 VTAIL.n511 104.615
R177 VTAIL.n562 VTAIL.n561 104.615
R178 VTAIL.n562 VTAIL.n507 104.615
R179 VTAIL.n569 VTAIL.n507 104.615
R180 VTAIL.n570 VTAIL.n569 104.615
R181 VTAIL.n26 VTAIL.n25 104.615
R182 VTAIL.n26 VTAIL.n19 104.615
R183 VTAIL.n33 VTAIL.n19 104.615
R184 VTAIL.n34 VTAIL.n33 104.615
R185 VTAIL.n34 VTAIL.n15 104.615
R186 VTAIL.n41 VTAIL.n15 104.615
R187 VTAIL.n42 VTAIL.n41 104.615
R188 VTAIL.n42 VTAIL.n11 104.615
R189 VTAIL.n49 VTAIL.n11 104.615
R190 VTAIL.n50 VTAIL.n49 104.615
R191 VTAIL.n50 VTAIL.n7 104.615
R192 VTAIL.n57 VTAIL.n7 104.615
R193 VTAIL.n58 VTAIL.n57 104.615
R194 VTAIL.n58 VTAIL.n3 104.615
R195 VTAIL.n65 VTAIL.n3 104.615
R196 VTAIL.n66 VTAIL.n65 104.615
R197 VTAIL.n98 VTAIL.n97 104.615
R198 VTAIL.n98 VTAIL.n91 104.615
R199 VTAIL.n105 VTAIL.n91 104.615
R200 VTAIL.n106 VTAIL.n105 104.615
R201 VTAIL.n106 VTAIL.n87 104.615
R202 VTAIL.n113 VTAIL.n87 104.615
R203 VTAIL.n114 VTAIL.n113 104.615
R204 VTAIL.n114 VTAIL.n83 104.615
R205 VTAIL.n121 VTAIL.n83 104.615
R206 VTAIL.n122 VTAIL.n121 104.615
R207 VTAIL.n122 VTAIL.n79 104.615
R208 VTAIL.n129 VTAIL.n79 104.615
R209 VTAIL.n130 VTAIL.n129 104.615
R210 VTAIL.n130 VTAIL.n75 104.615
R211 VTAIL.n137 VTAIL.n75 104.615
R212 VTAIL.n138 VTAIL.n137 104.615
R213 VTAIL.n170 VTAIL.n169 104.615
R214 VTAIL.n170 VTAIL.n163 104.615
R215 VTAIL.n177 VTAIL.n163 104.615
R216 VTAIL.n178 VTAIL.n177 104.615
R217 VTAIL.n178 VTAIL.n159 104.615
R218 VTAIL.n185 VTAIL.n159 104.615
R219 VTAIL.n186 VTAIL.n185 104.615
R220 VTAIL.n186 VTAIL.n155 104.615
R221 VTAIL.n193 VTAIL.n155 104.615
R222 VTAIL.n194 VTAIL.n193 104.615
R223 VTAIL.n194 VTAIL.n151 104.615
R224 VTAIL.n201 VTAIL.n151 104.615
R225 VTAIL.n202 VTAIL.n201 104.615
R226 VTAIL.n202 VTAIL.n147 104.615
R227 VTAIL.n209 VTAIL.n147 104.615
R228 VTAIL.n210 VTAIL.n209 104.615
R229 VTAIL.n498 VTAIL.n497 104.615
R230 VTAIL.n497 VTAIL.n435 104.615
R231 VTAIL.n490 VTAIL.n435 104.615
R232 VTAIL.n490 VTAIL.n489 104.615
R233 VTAIL.n489 VTAIL.n439 104.615
R234 VTAIL.n482 VTAIL.n439 104.615
R235 VTAIL.n482 VTAIL.n481 104.615
R236 VTAIL.n481 VTAIL.n443 104.615
R237 VTAIL.n474 VTAIL.n443 104.615
R238 VTAIL.n474 VTAIL.n473 104.615
R239 VTAIL.n473 VTAIL.n447 104.615
R240 VTAIL.n466 VTAIL.n447 104.615
R241 VTAIL.n466 VTAIL.n465 104.615
R242 VTAIL.n465 VTAIL.n451 104.615
R243 VTAIL.n458 VTAIL.n451 104.615
R244 VTAIL.n458 VTAIL.n457 104.615
R245 VTAIL.n426 VTAIL.n425 104.615
R246 VTAIL.n425 VTAIL.n363 104.615
R247 VTAIL.n418 VTAIL.n363 104.615
R248 VTAIL.n418 VTAIL.n417 104.615
R249 VTAIL.n417 VTAIL.n367 104.615
R250 VTAIL.n410 VTAIL.n367 104.615
R251 VTAIL.n410 VTAIL.n409 104.615
R252 VTAIL.n409 VTAIL.n371 104.615
R253 VTAIL.n402 VTAIL.n371 104.615
R254 VTAIL.n402 VTAIL.n401 104.615
R255 VTAIL.n401 VTAIL.n375 104.615
R256 VTAIL.n394 VTAIL.n375 104.615
R257 VTAIL.n394 VTAIL.n393 104.615
R258 VTAIL.n393 VTAIL.n379 104.615
R259 VTAIL.n386 VTAIL.n379 104.615
R260 VTAIL.n386 VTAIL.n385 104.615
R261 VTAIL.n354 VTAIL.n353 104.615
R262 VTAIL.n353 VTAIL.n291 104.615
R263 VTAIL.n346 VTAIL.n291 104.615
R264 VTAIL.n346 VTAIL.n345 104.615
R265 VTAIL.n345 VTAIL.n295 104.615
R266 VTAIL.n338 VTAIL.n295 104.615
R267 VTAIL.n338 VTAIL.n337 104.615
R268 VTAIL.n337 VTAIL.n299 104.615
R269 VTAIL.n330 VTAIL.n299 104.615
R270 VTAIL.n330 VTAIL.n329 104.615
R271 VTAIL.n329 VTAIL.n303 104.615
R272 VTAIL.n322 VTAIL.n303 104.615
R273 VTAIL.n322 VTAIL.n321 104.615
R274 VTAIL.n321 VTAIL.n307 104.615
R275 VTAIL.n314 VTAIL.n307 104.615
R276 VTAIL.n314 VTAIL.n313 104.615
R277 VTAIL.n282 VTAIL.n281 104.615
R278 VTAIL.n281 VTAIL.n219 104.615
R279 VTAIL.n274 VTAIL.n219 104.615
R280 VTAIL.n274 VTAIL.n273 104.615
R281 VTAIL.n273 VTAIL.n223 104.615
R282 VTAIL.n266 VTAIL.n223 104.615
R283 VTAIL.n266 VTAIL.n265 104.615
R284 VTAIL.n265 VTAIL.n227 104.615
R285 VTAIL.n258 VTAIL.n227 104.615
R286 VTAIL.n258 VTAIL.n257 104.615
R287 VTAIL.n257 VTAIL.n231 104.615
R288 VTAIL.n250 VTAIL.n231 104.615
R289 VTAIL.n250 VTAIL.n249 104.615
R290 VTAIL.n249 VTAIL.n235 104.615
R291 VTAIL.n242 VTAIL.n235 104.615
R292 VTAIL.n242 VTAIL.n241 104.615
R293 VTAIL.n529 VTAIL.t4 52.3082
R294 VTAIL.n25 VTAIL.t2 52.3082
R295 VTAIL.n97 VTAIL.t7 52.3082
R296 VTAIL.n169 VTAIL.t0 52.3082
R297 VTAIL.n457 VTAIL.t1 52.3082
R298 VTAIL.n385 VTAIL.t6 52.3082
R299 VTAIL.n313 VTAIL.t3 52.3082
R300 VTAIL.n241 VTAIL.t5 52.3082
R301 VTAIL.n575 VTAIL.n574 34.9005
R302 VTAIL.n71 VTAIL.n70 34.9005
R303 VTAIL.n143 VTAIL.n142 34.9005
R304 VTAIL.n215 VTAIL.n214 34.9005
R305 VTAIL.n503 VTAIL.n502 34.9005
R306 VTAIL.n431 VTAIL.n430 34.9005
R307 VTAIL.n359 VTAIL.n358 34.9005
R308 VTAIL.n287 VTAIL.n286 34.9005
R309 VTAIL.n575 VTAIL.n503 26.5824
R310 VTAIL.n287 VTAIL.n215 26.5824
R311 VTAIL.n528 VTAIL.n527 15.6677
R312 VTAIL.n24 VTAIL.n23 15.6677
R313 VTAIL.n96 VTAIL.n95 15.6677
R314 VTAIL.n168 VTAIL.n167 15.6677
R315 VTAIL.n456 VTAIL.n455 15.6677
R316 VTAIL.n384 VTAIL.n383 15.6677
R317 VTAIL.n312 VTAIL.n311 15.6677
R318 VTAIL.n240 VTAIL.n239 15.6677
R319 VTAIL.n531 VTAIL.n526 12.8005
R320 VTAIL.n572 VTAIL.n571 12.8005
R321 VTAIL.n27 VTAIL.n22 12.8005
R322 VTAIL.n68 VTAIL.n67 12.8005
R323 VTAIL.n99 VTAIL.n94 12.8005
R324 VTAIL.n140 VTAIL.n139 12.8005
R325 VTAIL.n171 VTAIL.n166 12.8005
R326 VTAIL.n212 VTAIL.n211 12.8005
R327 VTAIL.n500 VTAIL.n499 12.8005
R328 VTAIL.n459 VTAIL.n454 12.8005
R329 VTAIL.n428 VTAIL.n427 12.8005
R330 VTAIL.n387 VTAIL.n382 12.8005
R331 VTAIL.n356 VTAIL.n355 12.8005
R332 VTAIL.n315 VTAIL.n310 12.8005
R333 VTAIL.n284 VTAIL.n283 12.8005
R334 VTAIL.n243 VTAIL.n238 12.8005
R335 VTAIL.n532 VTAIL.n524 12.0247
R336 VTAIL.n568 VTAIL.n506 12.0247
R337 VTAIL.n28 VTAIL.n20 12.0247
R338 VTAIL.n64 VTAIL.n2 12.0247
R339 VTAIL.n100 VTAIL.n92 12.0247
R340 VTAIL.n136 VTAIL.n74 12.0247
R341 VTAIL.n172 VTAIL.n164 12.0247
R342 VTAIL.n208 VTAIL.n146 12.0247
R343 VTAIL.n496 VTAIL.n434 12.0247
R344 VTAIL.n460 VTAIL.n452 12.0247
R345 VTAIL.n424 VTAIL.n362 12.0247
R346 VTAIL.n388 VTAIL.n380 12.0247
R347 VTAIL.n352 VTAIL.n290 12.0247
R348 VTAIL.n316 VTAIL.n308 12.0247
R349 VTAIL.n280 VTAIL.n218 12.0247
R350 VTAIL.n244 VTAIL.n236 12.0247
R351 VTAIL.n536 VTAIL.n535 11.249
R352 VTAIL.n567 VTAIL.n508 11.249
R353 VTAIL.n32 VTAIL.n31 11.249
R354 VTAIL.n63 VTAIL.n4 11.249
R355 VTAIL.n104 VTAIL.n103 11.249
R356 VTAIL.n135 VTAIL.n76 11.249
R357 VTAIL.n176 VTAIL.n175 11.249
R358 VTAIL.n207 VTAIL.n148 11.249
R359 VTAIL.n495 VTAIL.n436 11.249
R360 VTAIL.n464 VTAIL.n463 11.249
R361 VTAIL.n423 VTAIL.n364 11.249
R362 VTAIL.n392 VTAIL.n391 11.249
R363 VTAIL.n351 VTAIL.n292 11.249
R364 VTAIL.n320 VTAIL.n319 11.249
R365 VTAIL.n279 VTAIL.n220 11.249
R366 VTAIL.n248 VTAIL.n247 11.249
R367 VTAIL.n539 VTAIL.n522 10.4732
R368 VTAIL.n564 VTAIL.n563 10.4732
R369 VTAIL.n35 VTAIL.n18 10.4732
R370 VTAIL.n60 VTAIL.n59 10.4732
R371 VTAIL.n107 VTAIL.n90 10.4732
R372 VTAIL.n132 VTAIL.n131 10.4732
R373 VTAIL.n179 VTAIL.n162 10.4732
R374 VTAIL.n204 VTAIL.n203 10.4732
R375 VTAIL.n492 VTAIL.n491 10.4732
R376 VTAIL.n467 VTAIL.n450 10.4732
R377 VTAIL.n420 VTAIL.n419 10.4732
R378 VTAIL.n395 VTAIL.n378 10.4732
R379 VTAIL.n348 VTAIL.n347 10.4732
R380 VTAIL.n323 VTAIL.n306 10.4732
R381 VTAIL.n276 VTAIL.n275 10.4732
R382 VTAIL.n251 VTAIL.n234 10.4732
R383 VTAIL.n540 VTAIL.n520 9.69747
R384 VTAIL.n560 VTAIL.n510 9.69747
R385 VTAIL.n36 VTAIL.n16 9.69747
R386 VTAIL.n56 VTAIL.n6 9.69747
R387 VTAIL.n108 VTAIL.n88 9.69747
R388 VTAIL.n128 VTAIL.n78 9.69747
R389 VTAIL.n180 VTAIL.n160 9.69747
R390 VTAIL.n200 VTAIL.n150 9.69747
R391 VTAIL.n488 VTAIL.n438 9.69747
R392 VTAIL.n468 VTAIL.n448 9.69747
R393 VTAIL.n416 VTAIL.n366 9.69747
R394 VTAIL.n396 VTAIL.n376 9.69747
R395 VTAIL.n344 VTAIL.n294 9.69747
R396 VTAIL.n324 VTAIL.n304 9.69747
R397 VTAIL.n272 VTAIL.n222 9.69747
R398 VTAIL.n252 VTAIL.n232 9.69747
R399 VTAIL.n574 VTAIL.n573 9.45567
R400 VTAIL.n70 VTAIL.n69 9.45567
R401 VTAIL.n142 VTAIL.n141 9.45567
R402 VTAIL.n214 VTAIL.n213 9.45567
R403 VTAIL.n502 VTAIL.n501 9.45567
R404 VTAIL.n430 VTAIL.n429 9.45567
R405 VTAIL.n358 VTAIL.n357 9.45567
R406 VTAIL.n286 VTAIL.n285 9.45567
R407 VTAIL.n549 VTAIL.n548 9.3005
R408 VTAIL.n518 VTAIL.n517 9.3005
R409 VTAIL.n543 VTAIL.n542 9.3005
R410 VTAIL.n541 VTAIL.n540 9.3005
R411 VTAIL.n522 VTAIL.n521 9.3005
R412 VTAIL.n535 VTAIL.n534 9.3005
R413 VTAIL.n533 VTAIL.n532 9.3005
R414 VTAIL.n526 VTAIL.n525 9.3005
R415 VTAIL.n551 VTAIL.n550 9.3005
R416 VTAIL.n514 VTAIL.n513 9.3005
R417 VTAIL.n557 VTAIL.n556 9.3005
R418 VTAIL.n559 VTAIL.n558 9.3005
R419 VTAIL.n510 VTAIL.n509 9.3005
R420 VTAIL.n565 VTAIL.n564 9.3005
R421 VTAIL.n567 VTAIL.n566 9.3005
R422 VTAIL.n506 VTAIL.n505 9.3005
R423 VTAIL.n573 VTAIL.n572 9.3005
R424 VTAIL.n45 VTAIL.n44 9.3005
R425 VTAIL.n14 VTAIL.n13 9.3005
R426 VTAIL.n39 VTAIL.n38 9.3005
R427 VTAIL.n37 VTAIL.n36 9.3005
R428 VTAIL.n18 VTAIL.n17 9.3005
R429 VTAIL.n31 VTAIL.n30 9.3005
R430 VTAIL.n29 VTAIL.n28 9.3005
R431 VTAIL.n22 VTAIL.n21 9.3005
R432 VTAIL.n47 VTAIL.n46 9.3005
R433 VTAIL.n10 VTAIL.n9 9.3005
R434 VTAIL.n53 VTAIL.n52 9.3005
R435 VTAIL.n55 VTAIL.n54 9.3005
R436 VTAIL.n6 VTAIL.n5 9.3005
R437 VTAIL.n61 VTAIL.n60 9.3005
R438 VTAIL.n63 VTAIL.n62 9.3005
R439 VTAIL.n2 VTAIL.n1 9.3005
R440 VTAIL.n69 VTAIL.n68 9.3005
R441 VTAIL.n117 VTAIL.n116 9.3005
R442 VTAIL.n86 VTAIL.n85 9.3005
R443 VTAIL.n111 VTAIL.n110 9.3005
R444 VTAIL.n109 VTAIL.n108 9.3005
R445 VTAIL.n90 VTAIL.n89 9.3005
R446 VTAIL.n103 VTAIL.n102 9.3005
R447 VTAIL.n101 VTAIL.n100 9.3005
R448 VTAIL.n94 VTAIL.n93 9.3005
R449 VTAIL.n119 VTAIL.n118 9.3005
R450 VTAIL.n82 VTAIL.n81 9.3005
R451 VTAIL.n125 VTAIL.n124 9.3005
R452 VTAIL.n127 VTAIL.n126 9.3005
R453 VTAIL.n78 VTAIL.n77 9.3005
R454 VTAIL.n133 VTAIL.n132 9.3005
R455 VTAIL.n135 VTAIL.n134 9.3005
R456 VTAIL.n74 VTAIL.n73 9.3005
R457 VTAIL.n141 VTAIL.n140 9.3005
R458 VTAIL.n189 VTAIL.n188 9.3005
R459 VTAIL.n158 VTAIL.n157 9.3005
R460 VTAIL.n183 VTAIL.n182 9.3005
R461 VTAIL.n181 VTAIL.n180 9.3005
R462 VTAIL.n162 VTAIL.n161 9.3005
R463 VTAIL.n175 VTAIL.n174 9.3005
R464 VTAIL.n173 VTAIL.n172 9.3005
R465 VTAIL.n166 VTAIL.n165 9.3005
R466 VTAIL.n191 VTAIL.n190 9.3005
R467 VTAIL.n154 VTAIL.n153 9.3005
R468 VTAIL.n197 VTAIL.n196 9.3005
R469 VTAIL.n199 VTAIL.n198 9.3005
R470 VTAIL.n150 VTAIL.n149 9.3005
R471 VTAIL.n205 VTAIL.n204 9.3005
R472 VTAIL.n207 VTAIL.n206 9.3005
R473 VTAIL.n146 VTAIL.n145 9.3005
R474 VTAIL.n213 VTAIL.n212 9.3005
R475 VTAIL.n442 VTAIL.n441 9.3005
R476 VTAIL.n485 VTAIL.n484 9.3005
R477 VTAIL.n487 VTAIL.n486 9.3005
R478 VTAIL.n438 VTAIL.n437 9.3005
R479 VTAIL.n493 VTAIL.n492 9.3005
R480 VTAIL.n495 VTAIL.n494 9.3005
R481 VTAIL.n434 VTAIL.n433 9.3005
R482 VTAIL.n501 VTAIL.n500 9.3005
R483 VTAIL.n479 VTAIL.n478 9.3005
R484 VTAIL.n477 VTAIL.n476 9.3005
R485 VTAIL.n446 VTAIL.n445 9.3005
R486 VTAIL.n471 VTAIL.n470 9.3005
R487 VTAIL.n469 VTAIL.n468 9.3005
R488 VTAIL.n450 VTAIL.n449 9.3005
R489 VTAIL.n463 VTAIL.n462 9.3005
R490 VTAIL.n461 VTAIL.n460 9.3005
R491 VTAIL.n454 VTAIL.n453 9.3005
R492 VTAIL.n370 VTAIL.n369 9.3005
R493 VTAIL.n413 VTAIL.n412 9.3005
R494 VTAIL.n415 VTAIL.n414 9.3005
R495 VTAIL.n366 VTAIL.n365 9.3005
R496 VTAIL.n421 VTAIL.n420 9.3005
R497 VTAIL.n423 VTAIL.n422 9.3005
R498 VTAIL.n362 VTAIL.n361 9.3005
R499 VTAIL.n429 VTAIL.n428 9.3005
R500 VTAIL.n407 VTAIL.n406 9.3005
R501 VTAIL.n405 VTAIL.n404 9.3005
R502 VTAIL.n374 VTAIL.n373 9.3005
R503 VTAIL.n399 VTAIL.n398 9.3005
R504 VTAIL.n397 VTAIL.n396 9.3005
R505 VTAIL.n378 VTAIL.n377 9.3005
R506 VTAIL.n391 VTAIL.n390 9.3005
R507 VTAIL.n389 VTAIL.n388 9.3005
R508 VTAIL.n382 VTAIL.n381 9.3005
R509 VTAIL.n298 VTAIL.n297 9.3005
R510 VTAIL.n341 VTAIL.n340 9.3005
R511 VTAIL.n343 VTAIL.n342 9.3005
R512 VTAIL.n294 VTAIL.n293 9.3005
R513 VTAIL.n349 VTAIL.n348 9.3005
R514 VTAIL.n351 VTAIL.n350 9.3005
R515 VTAIL.n290 VTAIL.n289 9.3005
R516 VTAIL.n357 VTAIL.n356 9.3005
R517 VTAIL.n335 VTAIL.n334 9.3005
R518 VTAIL.n333 VTAIL.n332 9.3005
R519 VTAIL.n302 VTAIL.n301 9.3005
R520 VTAIL.n327 VTAIL.n326 9.3005
R521 VTAIL.n325 VTAIL.n324 9.3005
R522 VTAIL.n306 VTAIL.n305 9.3005
R523 VTAIL.n319 VTAIL.n318 9.3005
R524 VTAIL.n317 VTAIL.n316 9.3005
R525 VTAIL.n310 VTAIL.n309 9.3005
R526 VTAIL.n226 VTAIL.n225 9.3005
R527 VTAIL.n269 VTAIL.n268 9.3005
R528 VTAIL.n271 VTAIL.n270 9.3005
R529 VTAIL.n222 VTAIL.n221 9.3005
R530 VTAIL.n277 VTAIL.n276 9.3005
R531 VTAIL.n279 VTAIL.n278 9.3005
R532 VTAIL.n218 VTAIL.n217 9.3005
R533 VTAIL.n285 VTAIL.n284 9.3005
R534 VTAIL.n263 VTAIL.n262 9.3005
R535 VTAIL.n261 VTAIL.n260 9.3005
R536 VTAIL.n230 VTAIL.n229 9.3005
R537 VTAIL.n255 VTAIL.n254 9.3005
R538 VTAIL.n253 VTAIL.n252 9.3005
R539 VTAIL.n234 VTAIL.n233 9.3005
R540 VTAIL.n247 VTAIL.n246 9.3005
R541 VTAIL.n245 VTAIL.n244 9.3005
R542 VTAIL.n238 VTAIL.n237 9.3005
R543 VTAIL.n544 VTAIL.n543 8.92171
R544 VTAIL.n559 VTAIL.n512 8.92171
R545 VTAIL.n40 VTAIL.n39 8.92171
R546 VTAIL.n55 VTAIL.n8 8.92171
R547 VTAIL.n112 VTAIL.n111 8.92171
R548 VTAIL.n127 VTAIL.n80 8.92171
R549 VTAIL.n184 VTAIL.n183 8.92171
R550 VTAIL.n199 VTAIL.n152 8.92171
R551 VTAIL.n487 VTAIL.n440 8.92171
R552 VTAIL.n472 VTAIL.n471 8.92171
R553 VTAIL.n415 VTAIL.n368 8.92171
R554 VTAIL.n400 VTAIL.n399 8.92171
R555 VTAIL.n343 VTAIL.n296 8.92171
R556 VTAIL.n328 VTAIL.n327 8.92171
R557 VTAIL.n271 VTAIL.n224 8.92171
R558 VTAIL.n256 VTAIL.n255 8.92171
R559 VTAIL.n574 VTAIL.n504 8.2187
R560 VTAIL.n70 VTAIL.n0 8.2187
R561 VTAIL.n142 VTAIL.n72 8.2187
R562 VTAIL.n214 VTAIL.n144 8.2187
R563 VTAIL.n502 VTAIL.n432 8.2187
R564 VTAIL.n430 VTAIL.n360 8.2187
R565 VTAIL.n358 VTAIL.n288 8.2187
R566 VTAIL.n286 VTAIL.n216 8.2187
R567 VTAIL.n547 VTAIL.n518 8.14595
R568 VTAIL.n556 VTAIL.n555 8.14595
R569 VTAIL.n43 VTAIL.n14 8.14595
R570 VTAIL.n52 VTAIL.n51 8.14595
R571 VTAIL.n115 VTAIL.n86 8.14595
R572 VTAIL.n124 VTAIL.n123 8.14595
R573 VTAIL.n187 VTAIL.n158 8.14595
R574 VTAIL.n196 VTAIL.n195 8.14595
R575 VTAIL.n484 VTAIL.n483 8.14595
R576 VTAIL.n475 VTAIL.n446 8.14595
R577 VTAIL.n412 VTAIL.n411 8.14595
R578 VTAIL.n403 VTAIL.n374 8.14595
R579 VTAIL.n340 VTAIL.n339 8.14595
R580 VTAIL.n331 VTAIL.n302 8.14595
R581 VTAIL.n268 VTAIL.n267 8.14595
R582 VTAIL.n259 VTAIL.n230 8.14595
R583 VTAIL.n548 VTAIL.n516 7.3702
R584 VTAIL.n552 VTAIL.n514 7.3702
R585 VTAIL.n44 VTAIL.n12 7.3702
R586 VTAIL.n48 VTAIL.n10 7.3702
R587 VTAIL.n116 VTAIL.n84 7.3702
R588 VTAIL.n120 VTAIL.n82 7.3702
R589 VTAIL.n188 VTAIL.n156 7.3702
R590 VTAIL.n192 VTAIL.n154 7.3702
R591 VTAIL.n480 VTAIL.n442 7.3702
R592 VTAIL.n476 VTAIL.n444 7.3702
R593 VTAIL.n408 VTAIL.n370 7.3702
R594 VTAIL.n404 VTAIL.n372 7.3702
R595 VTAIL.n336 VTAIL.n298 7.3702
R596 VTAIL.n332 VTAIL.n300 7.3702
R597 VTAIL.n264 VTAIL.n226 7.3702
R598 VTAIL.n260 VTAIL.n228 7.3702
R599 VTAIL.n551 VTAIL.n516 6.59444
R600 VTAIL.n552 VTAIL.n551 6.59444
R601 VTAIL.n47 VTAIL.n12 6.59444
R602 VTAIL.n48 VTAIL.n47 6.59444
R603 VTAIL.n119 VTAIL.n84 6.59444
R604 VTAIL.n120 VTAIL.n119 6.59444
R605 VTAIL.n191 VTAIL.n156 6.59444
R606 VTAIL.n192 VTAIL.n191 6.59444
R607 VTAIL.n480 VTAIL.n479 6.59444
R608 VTAIL.n479 VTAIL.n444 6.59444
R609 VTAIL.n408 VTAIL.n407 6.59444
R610 VTAIL.n407 VTAIL.n372 6.59444
R611 VTAIL.n336 VTAIL.n335 6.59444
R612 VTAIL.n335 VTAIL.n300 6.59444
R613 VTAIL.n264 VTAIL.n263 6.59444
R614 VTAIL.n263 VTAIL.n228 6.59444
R615 VTAIL.n548 VTAIL.n547 5.81868
R616 VTAIL.n555 VTAIL.n514 5.81868
R617 VTAIL.n44 VTAIL.n43 5.81868
R618 VTAIL.n51 VTAIL.n10 5.81868
R619 VTAIL.n116 VTAIL.n115 5.81868
R620 VTAIL.n123 VTAIL.n82 5.81868
R621 VTAIL.n188 VTAIL.n187 5.81868
R622 VTAIL.n195 VTAIL.n154 5.81868
R623 VTAIL.n483 VTAIL.n442 5.81868
R624 VTAIL.n476 VTAIL.n475 5.81868
R625 VTAIL.n411 VTAIL.n370 5.81868
R626 VTAIL.n404 VTAIL.n403 5.81868
R627 VTAIL.n339 VTAIL.n298 5.81868
R628 VTAIL.n332 VTAIL.n331 5.81868
R629 VTAIL.n267 VTAIL.n226 5.81868
R630 VTAIL.n260 VTAIL.n259 5.81868
R631 VTAIL.n572 VTAIL.n504 5.3904
R632 VTAIL.n68 VTAIL.n0 5.3904
R633 VTAIL.n140 VTAIL.n72 5.3904
R634 VTAIL.n212 VTAIL.n144 5.3904
R635 VTAIL.n500 VTAIL.n432 5.3904
R636 VTAIL.n428 VTAIL.n360 5.3904
R637 VTAIL.n356 VTAIL.n288 5.3904
R638 VTAIL.n284 VTAIL.n216 5.3904
R639 VTAIL.n544 VTAIL.n518 5.04292
R640 VTAIL.n556 VTAIL.n512 5.04292
R641 VTAIL.n40 VTAIL.n14 5.04292
R642 VTAIL.n52 VTAIL.n8 5.04292
R643 VTAIL.n112 VTAIL.n86 5.04292
R644 VTAIL.n124 VTAIL.n80 5.04292
R645 VTAIL.n184 VTAIL.n158 5.04292
R646 VTAIL.n196 VTAIL.n152 5.04292
R647 VTAIL.n484 VTAIL.n440 5.04292
R648 VTAIL.n472 VTAIL.n446 5.04292
R649 VTAIL.n412 VTAIL.n368 5.04292
R650 VTAIL.n400 VTAIL.n374 5.04292
R651 VTAIL.n340 VTAIL.n296 5.04292
R652 VTAIL.n328 VTAIL.n302 5.04292
R653 VTAIL.n268 VTAIL.n224 5.04292
R654 VTAIL.n256 VTAIL.n230 5.04292
R655 VTAIL.n527 VTAIL.n525 4.38563
R656 VTAIL.n23 VTAIL.n21 4.38563
R657 VTAIL.n95 VTAIL.n93 4.38563
R658 VTAIL.n167 VTAIL.n165 4.38563
R659 VTAIL.n455 VTAIL.n453 4.38563
R660 VTAIL.n383 VTAIL.n381 4.38563
R661 VTAIL.n311 VTAIL.n309 4.38563
R662 VTAIL.n239 VTAIL.n237 4.38563
R663 VTAIL.n543 VTAIL.n520 4.26717
R664 VTAIL.n560 VTAIL.n559 4.26717
R665 VTAIL.n39 VTAIL.n16 4.26717
R666 VTAIL.n56 VTAIL.n55 4.26717
R667 VTAIL.n111 VTAIL.n88 4.26717
R668 VTAIL.n128 VTAIL.n127 4.26717
R669 VTAIL.n183 VTAIL.n160 4.26717
R670 VTAIL.n200 VTAIL.n199 4.26717
R671 VTAIL.n488 VTAIL.n487 4.26717
R672 VTAIL.n471 VTAIL.n448 4.26717
R673 VTAIL.n416 VTAIL.n415 4.26717
R674 VTAIL.n399 VTAIL.n376 4.26717
R675 VTAIL.n344 VTAIL.n343 4.26717
R676 VTAIL.n327 VTAIL.n304 4.26717
R677 VTAIL.n272 VTAIL.n271 4.26717
R678 VTAIL.n255 VTAIL.n232 4.26717
R679 VTAIL.n540 VTAIL.n539 3.49141
R680 VTAIL.n563 VTAIL.n510 3.49141
R681 VTAIL.n36 VTAIL.n35 3.49141
R682 VTAIL.n59 VTAIL.n6 3.49141
R683 VTAIL.n108 VTAIL.n107 3.49141
R684 VTAIL.n131 VTAIL.n78 3.49141
R685 VTAIL.n180 VTAIL.n179 3.49141
R686 VTAIL.n203 VTAIL.n150 3.49141
R687 VTAIL.n491 VTAIL.n438 3.49141
R688 VTAIL.n468 VTAIL.n467 3.49141
R689 VTAIL.n419 VTAIL.n366 3.49141
R690 VTAIL.n396 VTAIL.n395 3.49141
R691 VTAIL.n347 VTAIL.n294 3.49141
R692 VTAIL.n324 VTAIL.n323 3.49141
R693 VTAIL.n275 VTAIL.n222 3.49141
R694 VTAIL.n252 VTAIL.n251 3.49141
R695 VTAIL.n359 VTAIL.n287 2.71602
R696 VTAIL.n503 VTAIL.n431 2.71602
R697 VTAIL.n215 VTAIL.n143 2.71602
R698 VTAIL.n536 VTAIL.n522 2.71565
R699 VTAIL.n564 VTAIL.n508 2.71565
R700 VTAIL.n32 VTAIL.n18 2.71565
R701 VTAIL.n60 VTAIL.n4 2.71565
R702 VTAIL.n104 VTAIL.n90 2.71565
R703 VTAIL.n132 VTAIL.n76 2.71565
R704 VTAIL.n176 VTAIL.n162 2.71565
R705 VTAIL.n204 VTAIL.n148 2.71565
R706 VTAIL.n492 VTAIL.n436 2.71565
R707 VTAIL.n464 VTAIL.n450 2.71565
R708 VTAIL.n420 VTAIL.n364 2.71565
R709 VTAIL.n392 VTAIL.n378 2.71565
R710 VTAIL.n348 VTAIL.n292 2.71565
R711 VTAIL.n320 VTAIL.n306 2.71565
R712 VTAIL.n276 VTAIL.n220 2.71565
R713 VTAIL.n248 VTAIL.n234 2.71565
R714 VTAIL.n535 VTAIL.n524 1.93989
R715 VTAIL.n568 VTAIL.n567 1.93989
R716 VTAIL.n31 VTAIL.n20 1.93989
R717 VTAIL.n64 VTAIL.n63 1.93989
R718 VTAIL.n103 VTAIL.n92 1.93989
R719 VTAIL.n136 VTAIL.n135 1.93989
R720 VTAIL.n175 VTAIL.n164 1.93989
R721 VTAIL.n208 VTAIL.n207 1.93989
R722 VTAIL.n496 VTAIL.n495 1.93989
R723 VTAIL.n463 VTAIL.n452 1.93989
R724 VTAIL.n424 VTAIL.n423 1.93989
R725 VTAIL.n391 VTAIL.n380 1.93989
R726 VTAIL.n352 VTAIL.n351 1.93989
R727 VTAIL.n319 VTAIL.n308 1.93989
R728 VTAIL.n280 VTAIL.n279 1.93989
R729 VTAIL.n247 VTAIL.n236 1.93989
R730 VTAIL VTAIL.n71 1.41645
R731 VTAIL VTAIL.n575 1.30007
R732 VTAIL.n532 VTAIL.n531 1.16414
R733 VTAIL.n571 VTAIL.n506 1.16414
R734 VTAIL.n28 VTAIL.n27 1.16414
R735 VTAIL.n67 VTAIL.n2 1.16414
R736 VTAIL.n100 VTAIL.n99 1.16414
R737 VTAIL.n139 VTAIL.n74 1.16414
R738 VTAIL.n172 VTAIL.n171 1.16414
R739 VTAIL.n211 VTAIL.n146 1.16414
R740 VTAIL.n499 VTAIL.n434 1.16414
R741 VTAIL.n460 VTAIL.n459 1.16414
R742 VTAIL.n427 VTAIL.n362 1.16414
R743 VTAIL.n388 VTAIL.n387 1.16414
R744 VTAIL.n355 VTAIL.n290 1.16414
R745 VTAIL.n316 VTAIL.n315 1.16414
R746 VTAIL.n283 VTAIL.n218 1.16414
R747 VTAIL.n244 VTAIL.n243 1.16414
R748 VTAIL.n431 VTAIL.n359 0.470328
R749 VTAIL.n143 VTAIL.n71 0.470328
R750 VTAIL.n528 VTAIL.n526 0.388379
R751 VTAIL.n24 VTAIL.n22 0.388379
R752 VTAIL.n96 VTAIL.n94 0.388379
R753 VTAIL.n168 VTAIL.n166 0.388379
R754 VTAIL.n456 VTAIL.n454 0.388379
R755 VTAIL.n384 VTAIL.n382 0.388379
R756 VTAIL.n312 VTAIL.n310 0.388379
R757 VTAIL.n240 VTAIL.n238 0.388379
R758 VTAIL.n533 VTAIL.n525 0.155672
R759 VTAIL.n534 VTAIL.n533 0.155672
R760 VTAIL.n534 VTAIL.n521 0.155672
R761 VTAIL.n541 VTAIL.n521 0.155672
R762 VTAIL.n542 VTAIL.n541 0.155672
R763 VTAIL.n542 VTAIL.n517 0.155672
R764 VTAIL.n549 VTAIL.n517 0.155672
R765 VTAIL.n550 VTAIL.n549 0.155672
R766 VTAIL.n550 VTAIL.n513 0.155672
R767 VTAIL.n557 VTAIL.n513 0.155672
R768 VTAIL.n558 VTAIL.n557 0.155672
R769 VTAIL.n558 VTAIL.n509 0.155672
R770 VTAIL.n565 VTAIL.n509 0.155672
R771 VTAIL.n566 VTAIL.n565 0.155672
R772 VTAIL.n566 VTAIL.n505 0.155672
R773 VTAIL.n573 VTAIL.n505 0.155672
R774 VTAIL.n29 VTAIL.n21 0.155672
R775 VTAIL.n30 VTAIL.n29 0.155672
R776 VTAIL.n30 VTAIL.n17 0.155672
R777 VTAIL.n37 VTAIL.n17 0.155672
R778 VTAIL.n38 VTAIL.n37 0.155672
R779 VTAIL.n38 VTAIL.n13 0.155672
R780 VTAIL.n45 VTAIL.n13 0.155672
R781 VTAIL.n46 VTAIL.n45 0.155672
R782 VTAIL.n46 VTAIL.n9 0.155672
R783 VTAIL.n53 VTAIL.n9 0.155672
R784 VTAIL.n54 VTAIL.n53 0.155672
R785 VTAIL.n54 VTAIL.n5 0.155672
R786 VTAIL.n61 VTAIL.n5 0.155672
R787 VTAIL.n62 VTAIL.n61 0.155672
R788 VTAIL.n62 VTAIL.n1 0.155672
R789 VTAIL.n69 VTAIL.n1 0.155672
R790 VTAIL.n101 VTAIL.n93 0.155672
R791 VTAIL.n102 VTAIL.n101 0.155672
R792 VTAIL.n102 VTAIL.n89 0.155672
R793 VTAIL.n109 VTAIL.n89 0.155672
R794 VTAIL.n110 VTAIL.n109 0.155672
R795 VTAIL.n110 VTAIL.n85 0.155672
R796 VTAIL.n117 VTAIL.n85 0.155672
R797 VTAIL.n118 VTAIL.n117 0.155672
R798 VTAIL.n118 VTAIL.n81 0.155672
R799 VTAIL.n125 VTAIL.n81 0.155672
R800 VTAIL.n126 VTAIL.n125 0.155672
R801 VTAIL.n126 VTAIL.n77 0.155672
R802 VTAIL.n133 VTAIL.n77 0.155672
R803 VTAIL.n134 VTAIL.n133 0.155672
R804 VTAIL.n134 VTAIL.n73 0.155672
R805 VTAIL.n141 VTAIL.n73 0.155672
R806 VTAIL.n173 VTAIL.n165 0.155672
R807 VTAIL.n174 VTAIL.n173 0.155672
R808 VTAIL.n174 VTAIL.n161 0.155672
R809 VTAIL.n181 VTAIL.n161 0.155672
R810 VTAIL.n182 VTAIL.n181 0.155672
R811 VTAIL.n182 VTAIL.n157 0.155672
R812 VTAIL.n189 VTAIL.n157 0.155672
R813 VTAIL.n190 VTAIL.n189 0.155672
R814 VTAIL.n190 VTAIL.n153 0.155672
R815 VTAIL.n197 VTAIL.n153 0.155672
R816 VTAIL.n198 VTAIL.n197 0.155672
R817 VTAIL.n198 VTAIL.n149 0.155672
R818 VTAIL.n205 VTAIL.n149 0.155672
R819 VTAIL.n206 VTAIL.n205 0.155672
R820 VTAIL.n206 VTAIL.n145 0.155672
R821 VTAIL.n213 VTAIL.n145 0.155672
R822 VTAIL.n501 VTAIL.n433 0.155672
R823 VTAIL.n494 VTAIL.n433 0.155672
R824 VTAIL.n494 VTAIL.n493 0.155672
R825 VTAIL.n493 VTAIL.n437 0.155672
R826 VTAIL.n486 VTAIL.n437 0.155672
R827 VTAIL.n486 VTAIL.n485 0.155672
R828 VTAIL.n485 VTAIL.n441 0.155672
R829 VTAIL.n478 VTAIL.n441 0.155672
R830 VTAIL.n478 VTAIL.n477 0.155672
R831 VTAIL.n477 VTAIL.n445 0.155672
R832 VTAIL.n470 VTAIL.n445 0.155672
R833 VTAIL.n470 VTAIL.n469 0.155672
R834 VTAIL.n469 VTAIL.n449 0.155672
R835 VTAIL.n462 VTAIL.n449 0.155672
R836 VTAIL.n462 VTAIL.n461 0.155672
R837 VTAIL.n461 VTAIL.n453 0.155672
R838 VTAIL.n429 VTAIL.n361 0.155672
R839 VTAIL.n422 VTAIL.n361 0.155672
R840 VTAIL.n422 VTAIL.n421 0.155672
R841 VTAIL.n421 VTAIL.n365 0.155672
R842 VTAIL.n414 VTAIL.n365 0.155672
R843 VTAIL.n414 VTAIL.n413 0.155672
R844 VTAIL.n413 VTAIL.n369 0.155672
R845 VTAIL.n406 VTAIL.n369 0.155672
R846 VTAIL.n406 VTAIL.n405 0.155672
R847 VTAIL.n405 VTAIL.n373 0.155672
R848 VTAIL.n398 VTAIL.n373 0.155672
R849 VTAIL.n398 VTAIL.n397 0.155672
R850 VTAIL.n397 VTAIL.n377 0.155672
R851 VTAIL.n390 VTAIL.n377 0.155672
R852 VTAIL.n390 VTAIL.n389 0.155672
R853 VTAIL.n389 VTAIL.n381 0.155672
R854 VTAIL.n357 VTAIL.n289 0.155672
R855 VTAIL.n350 VTAIL.n289 0.155672
R856 VTAIL.n350 VTAIL.n349 0.155672
R857 VTAIL.n349 VTAIL.n293 0.155672
R858 VTAIL.n342 VTAIL.n293 0.155672
R859 VTAIL.n342 VTAIL.n341 0.155672
R860 VTAIL.n341 VTAIL.n297 0.155672
R861 VTAIL.n334 VTAIL.n297 0.155672
R862 VTAIL.n334 VTAIL.n333 0.155672
R863 VTAIL.n333 VTAIL.n301 0.155672
R864 VTAIL.n326 VTAIL.n301 0.155672
R865 VTAIL.n326 VTAIL.n325 0.155672
R866 VTAIL.n325 VTAIL.n305 0.155672
R867 VTAIL.n318 VTAIL.n305 0.155672
R868 VTAIL.n318 VTAIL.n317 0.155672
R869 VTAIL.n317 VTAIL.n309 0.155672
R870 VTAIL.n285 VTAIL.n217 0.155672
R871 VTAIL.n278 VTAIL.n217 0.155672
R872 VTAIL.n278 VTAIL.n277 0.155672
R873 VTAIL.n277 VTAIL.n221 0.155672
R874 VTAIL.n270 VTAIL.n221 0.155672
R875 VTAIL.n270 VTAIL.n269 0.155672
R876 VTAIL.n269 VTAIL.n225 0.155672
R877 VTAIL.n262 VTAIL.n225 0.155672
R878 VTAIL.n262 VTAIL.n261 0.155672
R879 VTAIL.n261 VTAIL.n229 0.155672
R880 VTAIL.n254 VTAIL.n229 0.155672
R881 VTAIL.n254 VTAIL.n253 0.155672
R882 VTAIL.n253 VTAIL.n233 0.155672
R883 VTAIL.n246 VTAIL.n233 0.155672
R884 VTAIL.n246 VTAIL.n245 0.155672
R885 VTAIL.n245 VTAIL.n237 0.155672
R886 B.n806 B.n805 585
R887 B.n807 B.n806 585
R888 B.n322 B.n119 585
R889 B.n321 B.n320 585
R890 B.n319 B.n318 585
R891 B.n317 B.n316 585
R892 B.n315 B.n314 585
R893 B.n313 B.n312 585
R894 B.n311 B.n310 585
R895 B.n309 B.n308 585
R896 B.n307 B.n306 585
R897 B.n305 B.n304 585
R898 B.n303 B.n302 585
R899 B.n301 B.n300 585
R900 B.n299 B.n298 585
R901 B.n297 B.n296 585
R902 B.n295 B.n294 585
R903 B.n293 B.n292 585
R904 B.n291 B.n290 585
R905 B.n289 B.n288 585
R906 B.n287 B.n286 585
R907 B.n285 B.n284 585
R908 B.n283 B.n282 585
R909 B.n281 B.n280 585
R910 B.n279 B.n278 585
R911 B.n277 B.n276 585
R912 B.n275 B.n274 585
R913 B.n273 B.n272 585
R914 B.n271 B.n270 585
R915 B.n269 B.n268 585
R916 B.n267 B.n266 585
R917 B.n265 B.n264 585
R918 B.n263 B.n262 585
R919 B.n261 B.n260 585
R920 B.n259 B.n258 585
R921 B.n257 B.n256 585
R922 B.n255 B.n254 585
R923 B.n253 B.n252 585
R924 B.n251 B.n250 585
R925 B.n249 B.n248 585
R926 B.n247 B.n246 585
R927 B.n245 B.n244 585
R928 B.n243 B.n242 585
R929 B.n241 B.n240 585
R930 B.n239 B.n238 585
R931 B.n237 B.n236 585
R932 B.n235 B.n234 585
R933 B.n232 B.n231 585
R934 B.n230 B.n229 585
R935 B.n228 B.n227 585
R936 B.n226 B.n225 585
R937 B.n224 B.n223 585
R938 B.n222 B.n221 585
R939 B.n220 B.n219 585
R940 B.n218 B.n217 585
R941 B.n216 B.n215 585
R942 B.n214 B.n213 585
R943 B.n212 B.n211 585
R944 B.n210 B.n209 585
R945 B.n208 B.n207 585
R946 B.n206 B.n205 585
R947 B.n204 B.n203 585
R948 B.n202 B.n201 585
R949 B.n200 B.n199 585
R950 B.n198 B.n197 585
R951 B.n196 B.n195 585
R952 B.n194 B.n193 585
R953 B.n192 B.n191 585
R954 B.n190 B.n189 585
R955 B.n188 B.n187 585
R956 B.n186 B.n185 585
R957 B.n184 B.n183 585
R958 B.n182 B.n181 585
R959 B.n180 B.n179 585
R960 B.n178 B.n177 585
R961 B.n176 B.n175 585
R962 B.n174 B.n173 585
R963 B.n172 B.n171 585
R964 B.n170 B.n169 585
R965 B.n168 B.n167 585
R966 B.n166 B.n165 585
R967 B.n164 B.n163 585
R968 B.n162 B.n161 585
R969 B.n160 B.n159 585
R970 B.n158 B.n157 585
R971 B.n156 B.n155 585
R972 B.n154 B.n153 585
R973 B.n152 B.n151 585
R974 B.n150 B.n149 585
R975 B.n148 B.n147 585
R976 B.n146 B.n145 585
R977 B.n144 B.n143 585
R978 B.n142 B.n141 585
R979 B.n140 B.n139 585
R980 B.n138 B.n137 585
R981 B.n136 B.n135 585
R982 B.n134 B.n133 585
R983 B.n132 B.n131 585
R984 B.n130 B.n129 585
R985 B.n128 B.n127 585
R986 B.n126 B.n125 585
R987 B.n67 B.n66 585
R988 B.n804 B.n68 585
R989 B.n808 B.n68 585
R990 B.n803 B.n802 585
R991 B.n802 B.n64 585
R992 B.n801 B.n63 585
R993 B.n814 B.n63 585
R994 B.n800 B.n62 585
R995 B.n815 B.n62 585
R996 B.n799 B.n61 585
R997 B.n816 B.n61 585
R998 B.n798 B.n797 585
R999 B.n797 B.n57 585
R1000 B.n796 B.n56 585
R1001 B.n822 B.n56 585
R1002 B.n795 B.n55 585
R1003 B.n823 B.n55 585
R1004 B.n794 B.n54 585
R1005 B.n824 B.n54 585
R1006 B.n793 B.n792 585
R1007 B.n792 B.n50 585
R1008 B.n791 B.n49 585
R1009 B.n830 B.n49 585
R1010 B.n790 B.n48 585
R1011 B.n831 B.n48 585
R1012 B.n789 B.n47 585
R1013 B.n832 B.n47 585
R1014 B.n788 B.n787 585
R1015 B.n787 B.n43 585
R1016 B.n786 B.n42 585
R1017 B.n838 B.n42 585
R1018 B.n785 B.n41 585
R1019 B.n839 B.n41 585
R1020 B.n784 B.n40 585
R1021 B.n840 B.n40 585
R1022 B.n783 B.n782 585
R1023 B.n782 B.n36 585
R1024 B.n781 B.n35 585
R1025 B.n846 B.n35 585
R1026 B.n780 B.n34 585
R1027 B.n847 B.n34 585
R1028 B.n779 B.n33 585
R1029 B.n848 B.n33 585
R1030 B.n778 B.n777 585
R1031 B.n777 B.n29 585
R1032 B.n776 B.n28 585
R1033 B.n854 B.n28 585
R1034 B.n775 B.n27 585
R1035 B.n855 B.n27 585
R1036 B.n774 B.n26 585
R1037 B.n856 B.n26 585
R1038 B.n773 B.n772 585
R1039 B.n772 B.n22 585
R1040 B.n771 B.n21 585
R1041 B.n862 B.n21 585
R1042 B.n770 B.n20 585
R1043 B.n863 B.n20 585
R1044 B.n769 B.n19 585
R1045 B.n864 B.n19 585
R1046 B.n768 B.n767 585
R1047 B.n767 B.n18 585
R1048 B.n766 B.n14 585
R1049 B.n870 B.n14 585
R1050 B.n765 B.n13 585
R1051 B.n871 B.n13 585
R1052 B.n764 B.n12 585
R1053 B.n872 B.n12 585
R1054 B.n763 B.n762 585
R1055 B.n762 B.n8 585
R1056 B.n761 B.n7 585
R1057 B.n878 B.n7 585
R1058 B.n760 B.n6 585
R1059 B.n879 B.n6 585
R1060 B.n759 B.n5 585
R1061 B.n880 B.n5 585
R1062 B.n758 B.n757 585
R1063 B.n757 B.n4 585
R1064 B.n756 B.n323 585
R1065 B.n756 B.n755 585
R1066 B.n746 B.n324 585
R1067 B.n325 B.n324 585
R1068 B.n748 B.n747 585
R1069 B.n749 B.n748 585
R1070 B.n745 B.n330 585
R1071 B.n330 B.n329 585
R1072 B.n744 B.n743 585
R1073 B.n743 B.n742 585
R1074 B.n332 B.n331 585
R1075 B.n735 B.n332 585
R1076 B.n734 B.n733 585
R1077 B.n736 B.n734 585
R1078 B.n732 B.n337 585
R1079 B.n337 B.n336 585
R1080 B.n731 B.n730 585
R1081 B.n730 B.n729 585
R1082 B.n339 B.n338 585
R1083 B.n340 B.n339 585
R1084 B.n722 B.n721 585
R1085 B.n723 B.n722 585
R1086 B.n720 B.n345 585
R1087 B.n345 B.n344 585
R1088 B.n719 B.n718 585
R1089 B.n718 B.n717 585
R1090 B.n347 B.n346 585
R1091 B.n348 B.n347 585
R1092 B.n710 B.n709 585
R1093 B.n711 B.n710 585
R1094 B.n708 B.n353 585
R1095 B.n353 B.n352 585
R1096 B.n707 B.n706 585
R1097 B.n706 B.n705 585
R1098 B.n355 B.n354 585
R1099 B.n356 B.n355 585
R1100 B.n698 B.n697 585
R1101 B.n699 B.n698 585
R1102 B.n696 B.n361 585
R1103 B.n361 B.n360 585
R1104 B.n695 B.n694 585
R1105 B.n694 B.n693 585
R1106 B.n363 B.n362 585
R1107 B.n364 B.n363 585
R1108 B.n686 B.n685 585
R1109 B.n687 B.n686 585
R1110 B.n684 B.n369 585
R1111 B.n369 B.n368 585
R1112 B.n683 B.n682 585
R1113 B.n682 B.n681 585
R1114 B.n371 B.n370 585
R1115 B.n372 B.n371 585
R1116 B.n674 B.n673 585
R1117 B.n675 B.n674 585
R1118 B.n672 B.n377 585
R1119 B.n377 B.n376 585
R1120 B.n671 B.n670 585
R1121 B.n670 B.n669 585
R1122 B.n379 B.n378 585
R1123 B.n380 B.n379 585
R1124 B.n662 B.n661 585
R1125 B.n663 B.n662 585
R1126 B.n660 B.n385 585
R1127 B.n385 B.n384 585
R1128 B.n659 B.n658 585
R1129 B.n658 B.n657 585
R1130 B.n387 B.n386 585
R1131 B.n388 B.n387 585
R1132 B.n650 B.n649 585
R1133 B.n651 B.n650 585
R1134 B.n391 B.n390 585
R1135 B.n448 B.n446 585
R1136 B.n449 B.n445 585
R1137 B.n449 B.n392 585
R1138 B.n452 B.n451 585
R1139 B.n453 B.n444 585
R1140 B.n455 B.n454 585
R1141 B.n457 B.n443 585
R1142 B.n460 B.n459 585
R1143 B.n461 B.n442 585
R1144 B.n463 B.n462 585
R1145 B.n465 B.n441 585
R1146 B.n468 B.n467 585
R1147 B.n469 B.n440 585
R1148 B.n471 B.n470 585
R1149 B.n473 B.n439 585
R1150 B.n476 B.n475 585
R1151 B.n477 B.n438 585
R1152 B.n479 B.n478 585
R1153 B.n481 B.n437 585
R1154 B.n484 B.n483 585
R1155 B.n485 B.n436 585
R1156 B.n487 B.n486 585
R1157 B.n489 B.n435 585
R1158 B.n492 B.n491 585
R1159 B.n493 B.n434 585
R1160 B.n495 B.n494 585
R1161 B.n497 B.n433 585
R1162 B.n500 B.n499 585
R1163 B.n501 B.n432 585
R1164 B.n503 B.n502 585
R1165 B.n505 B.n431 585
R1166 B.n508 B.n507 585
R1167 B.n509 B.n430 585
R1168 B.n511 B.n510 585
R1169 B.n513 B.n429 585
R1170 B.n516 B.n515 585
R1171 B.n517 B.n428 585
R1172 B.n519 B.n518 585
R1173 B.n521 B.n427 585
R1174 B.n524 B.n523 585
R1175 B.n525 B.n426 585
R1176 B.n527 B.n526 585
R1177 B.n529 B.n425 585
R1178 B.n532 B.n531 585
R1179 B.n533 B.n424 585
R1180 B.n538 B.n537 585
R1181 B.n540 B.n423 585
R1182 B.n543 B.n542 585
R1183 B.n544 B.n422 585
R1184 B.n546 B.n545 585
R1185 B.n548 B.n421 585
R1186 B.n551 B.n550 585
R1187 B.n552 B.n420 585
R1188 B.n554 B.n553 585
R1189 B.n556 B.n419 585
R1190 B.n559 B.n558 585
R1191 B.n560 B.n415 585
R1192 B.n562 B.n561 585
R1193 B.n564 B.n414 585
R1194 B.n567 B.n566 585
R1195 B.n568 B.n413 585
R1196 B.n570 B.n569 585
R1197 B.n572 B.n412 585
R1198 B.n575 B.n574 585
R1199 B.n576 B.n411 585
R1200 B.n578 B.n577 585
R1201 B.n580 B.n410 585
R1202 B.n583 B.n582 585
R1203 B.n584 B.n409 585
R1204 B.n586 B.n585 585
R1205 B.n588 B.n408 585
R1206 B.n591 B.n590 585
R1207 B.n592 B.n407 585
R1208 B.n594 B.n593 585
R1209 B.n596 B.n406 585
R1210 B.n599 B.n598 585
R1211 B.n600 B.n405 585
R1212 B.n602 B.n601 585
R1213 B.n604 B.n404 585
R1214 B.n607 B.n606 585
R1215 B.n608 B.n403 585
R1216 B.n610 B.n609 585
R1217 B.n612 B.n402 585
R1218 B.n615 B.n614 585
R1219 B.n616 B.n401 585
R1220 B.n618 B.n617 585
R1221 B.n620 B.n400 585
R1222 B.n623 B.n622 585
R1223 B.n624 B.n399 585
R1224 B.n626 B.n625 585
R1225 B.n628 B.n398 585
R1226 B.n631 B.n630 585
R1227 B.n632 B.n397 585
R1228 B.n634 B.n633 585
R1229 B.n636 B.n396 585
R1230 B.n639 B.n638 585
R1231 B.n640 B.n395 585
R1232 B.n642 B.n641 585
R1233 B.n644 B.n394 585
R1234 B.n647 B.n646 585
R1235 B.n648 B.n393 585
R1236 B.n653 B.n652 585
R1237 B.n652 B.n651 585
R1238 B.n654 B.n389 585
R1239 B.n389 B.n388 585
R1240 B.n656 B.n655 585
R1241 B.n657 B.n656 585
R1242 B.n383 B.n382 585
R1243 B.n384 B.n383 585
R1244 B.n665 B.n664 585
R1245 B.n664 B.n663 585
R1246 B.n666 B.n381 585
R1247 B.n381 B.n380 585
R1248 B.n668 B.n667 585
R1249 B.n669 B.n668 585
R1250 B.n375 B.n374 585
R1251 B.n376 B.n375 585
R1252 B.n677 B.n676 585
R1253 B.n676 B.n675 585
R1254 B.n678 B.n373 585
R1255 B.n373 B.n372 585
R1256 B.n680 B.n679 585
R1257 B.n681 B.n680 585
R1258 B.n367 B.n366 585
R1259 B.n368 B.n367 585
R1260 B.n689 B.n688 585
R1261 B.n688 B.n687 585
R1262 B.n690 B.n365 585
R1263 B.n365 B.n364 585
R1264 B.n692 B.n691 585
R1265 B.n693 B.n692 585
R1266 B.n359 B.n358 585
R1267 B.n360 B.n359 585
R1268 B.n701 B.n700 585
R1269 B.n700 B.n699 585
R1270 B.n702 B.n357 585
R1271 B.n357 B.n356 585
R1272 B.n704 B.n703 585
R1273 B.n705 B.n704 585
R1274 B.n351 B.n350 585
R1275 B.n352 B.n351 585
R1276 B.n713 B.n712 585
R1277 B.n712 B.n711 585
R1278 B.n714 B.n349 585
R1279 B.n349 B.n348 585
R1280 B.n716 B.n715 585
R1281 B.n717 B.n716 585
R1282 B.n343 B.n342 585
R1283 B.n344 B.n343 585
R1284 B.n725 B.n724 585
R1285 B.n724 B.n723 585
R1286 B.n726 B.n341 585
R1287 B.n341 B.n340 585
R1288 B.n728 B.n727 585
R1289 B.n729 B.n728 585
R1290 B.n335 B.n334 585
R1291 B.n336 B.n335 585
R1292 B.n738 B.n737 585
R1293 B.n737 B.n736 585
R1294 B.n739 B.n333 585
R1295 B.n735 B.n333 585
R1296 B.n741 B.n740 585
R1297 B.n742 B.n741 585
R1298 B.n328 B.n327 585
R1299 B.n329 B.n328 585
R1300 B.n751 B.n750 585
R1301 B.n750 B.n749 585
R1302 B.n752 B.n326 585
R1303 B.n326 B.n325 585
R1304 B.n754 B.n753 585
R1305 B.n755 B.n754 585
R1306 B.n2 B.n0 585
R1307 B.n4 B.n2 585
R1308 B.n3 B.n1 585
R1309 B.n879 B.n3 585
R1310 B.n877 B.n876 585
R1311 B.n878 B.n877 585
R1312 B.n875 B.n9 585
R1313 B.n9 B.n8 585
R1314 B.n874 B.n873 585
R1315 B.n873 B.n872 585
R1316 B.n11 B.n10 585
R1317 B.n871 B.n11 585
R1318 B.n869 B.n868 585
R1319 B.n870 B.n869 585
R1320 B.n867 B.n15 585
R1321 B.n18 B.n15 585
R1322 B.n866 B.n865 585
R1323 B.n865 B.n864 585
R1324 B.n17 B.n16 585
R1325 B.n863 B.n17 585
R1326 B.n861 B.n860 585
R1327 B.n862 B.n861 585
R1328 B.n859 B.n23 585
R1329 B.n23 B.n22 585
R1330 B.n858 B.n857 585
R1331 B.n857 B.n856 585
R1332 B.n25 B.n24 585
R1333 B.n855 B.n25 585
R1334 B.n853 B.n852 585
R1335 B.n854 B.n853 585
R1336 B.n851 B.n30 585
R1337 B.n30 B.n29 585
R1338 B.n850 B.n849 585
R1339 B.n849 B.n848 585
R1340 B.n32 B.n31 585
R1341 B.n847 B.n32 585
R1342 B.n845 B.n844 585
R1343 B.n846 B.n845 585
R1344 B.n843 B.n37 585
R1345 B.n37 B.n36 585
R1346 B.n842 B.n841 585
R1347 B.n841 B.n840 585
R1348 B.n39 B.n38 585
R1349 B.n839 B.n39 585
R1350 B.n837 B.n836 585
R1351 B.n838 B.n837 585
R1352 B.n835 B.n44 585
R1353 B.n44 B.n43 585
R1354 B.n834 B.n833 585
R1355 B.n833 B.n832 585
R1356 B.n46 B.n45 585
R1357 B.n831 B.n46 585
R1358 B.n829 B.n828 585
R1359 B.n830 B.n829 585
R1360 B.n827 B.n51 585
R1361 B.n51 B.n50 585
R1362 B.n826 B.n825 585
R1363 B.n825 B.n824 585
R1364 B.n53 B.n52 585
R1365 B.n823 B.n53 585
R1366 B.n821 B.n820 585
R1367 B.n822 B.n821 585
R1368 B.n819 B.n58 585
R1369 B.n58 B.n57 585
R1370 B.n818 B.n817 585
R1371 B.n817 B.n816 585
R1372 B.n60 B.n59 585
R1373 B.n815 B.n60 585
R1374 B.n813 B.n812 585
R1375 B.n814 B.n813 585
R1376 B.n811 B.n65 585
R1377 B.n65 B.n64 585
R1378 B.n810 B.n809 585
R1379 B.n809 B.n808 585
R1380 B.n882 B.n881 585
R1381 B.n881 B.n880 585
R1382 B.n652 B.n391 458.866
R1383 B.n809 B.n67 458.866
R1384 B.n650 B.n393 458.866
R1385 B.n806 B.n68 458.866
R1386 B.n416 B.t11 366.135
R1387 B.n120 B.t6 366.135
R1388 B.n534 B.t17 366.135
R1389 B.n122 B.t13 366.135
R1390 B.n416 B.t8 322.361
R1391 B.n534 B.t15 322.361
R1392 B.n122 B.t12 322.361
R1393 B.n120 B.t4 322.361
R1394 B.n417 B.t10 305.046
R1395 B.n121 B.t7 305.046
R1396 B.n535 B.t16 305.045
R1397 B.n123 B.t14 305.045
R1398 B.n807 B.n118 256.663
R1399 B.n807 B.n117 256.663
R1400 B.n807 B.n116 256.663
R1401 B.n807 B.n115 256.663
R1402 B.n807 B.n114 256.663
R1403 B.n807 B.n113 256.663
R1404 B.n807 B.n112 256.663
R1405 B.n807 B.n111 256.663
R1406 B.n807 B.n110 256.663
R1407 B.n807 B.n109 256.663
R1408 B.n807 B.n108 256.663
R1409 B.n807 B.n107 256.663
R1410 B.n807 B.n106 256.663
R1411 B.n807 B.n105 256.663
R1412 B.n807 B.n104 256.663
R1413 B.n807 B.n103 256.663
R1414 B.n807 B.n102 256.663
R1415 B.n807 B.n101 256.663
R1416 B.n807 B.n100 256.663
R1417 B.n807 B.n99 256.663
R1418 B.n807 B.n98 256.663
R1419 B.n807 B.n97 256.663
R1420 B.n807 B.n96 256.663
R1421 B.n807 B.n95 256.663
R1422 B.n807 B.n94 256.663
R1423 B.n807 B.n93 256.663
R1424 B.n807 B.n92 256.663
R1425 B.n807 B.n91 256.663
R1426 B.n807 B.n90 256.663
R1427 B.n807 B.n89 256.663
R1428 B.n807 B.n88 256.663
R1429 B.n807 B.n87 256.663
R1430 B.n807 B.n86 256.663
R1431 B.n807 B.n85 256.663
R1432 B.n807 B.n84 256.663
R1433 B.n807 B.n83 256.663
R1434 B.n807 B.n82 256.663
R1435 B.n807 B.n81 256.663
R1436 B.n807 B.n80 256.663
R1437 B.n807 B.n79 256.663
R1438 B.n807 B.n78 256.663
R1439 B.n807 B.n77 256.663
R1440 B.n807 B.n76 256.663
R1441 B.n807 B.n75 256.663
R1442 B.n807 B.n74 256.663
R1443 B.n807 B.n73 256.663
R1444 B.n807 B.n72 256.663
R1445 B.n807 B.n71 256.663
R1446 B.n807 B.n70 256.663
R1447 B.n807 B.n69 256.663
R1448 B.n447 B.n392 256.663
R1449 B.n450 B.n392 256.663
R1450 B.n456 B.n392 256.663
R1451 B.n458 B.n392 256.663
R1452 B.n464 B.n392 256.663
R1453 B.n466 B.n392 256.663
R1454 B.n472 B.n392 256.663
R1455 B.n474 B.n392 256.663
R1456 B.n480 B.n392 256.663
R1457 B.n482 B.n392 256.663
R1458 B.n488 B.n392 256.663
R1459 B.n490 B.n392 256.663
R1460 B.n496 B.n392 256.663
R1461 B.n498 B.n392 256.663
R1462 B.n504 B.n392 256.663
R1463 B.n506 B.n392 256.663
R1464 B.n512 B.n392 256.663
R1465 B.n514 B.n392 256.663
R1466 B.n520 B.n392 256.663
R1467 B.n522 B.n392 256.663
R1468 B.n528 B.n392 256.663
R1469 B.n530 B.n392 256.663
R1470 B.n539 B.n392 256.663
R1471 B.n541 B.n392 256.663
R1472 B.n547 B.n392 256.663
R1473 B.n549 B.n392 256.663
R1474 B.n555 B.n392 256.663
R1475 B.n557 B.n392 256.663
R1476 B.n563 B.n392 256.663
R1477 B.n565 B.n392 256.663
R1478 B.n571 B.n392 256.663
R1479 B.n573 B.n392 256.663
R1480 B.n579 B.n392 256.663
R1481 B.n581 B.n392 256.663
R1482 B.n587 B.n392 256.663
R1483 B.n589 B.n392 256.663
R1484 B.n595 B.n392 256.663
R1485 B.n597 B.n392 256.663
R1486 B.n603 B.n392 256.663
R1487 B.n605 B.n392 256.663
R1488 B.n611 B.n392 256.663
R1489 B.n613 B.n392 256.663
R1490 B.n619 B.n392 256.663
R1491 B.n621 B.n392 256.663
R1492 B.n627 B.n392 256.663
R1493 B.n629 B.n392 256.663
R1494 B.n635 B.n392 256.663
R1495 B.n637 B.n392 256.663
R1496 B.n643 B.n392 256.663
R1497 B.n645 B.n392 256.663
R1498 B.n652 B.n389 163.367
R1499 B.n656 B.n389 163.367
R1500 B.n656 B.n383 163.367
R1501 B.n664 B.n383 163.367
R1502 B.n664 B.n381 163.367
R1503 B.n668 B.n381 163.367
R1504 B.n668 B.n375 163.367
R1505 B.n676 B.n375 163.367
R1506 B.n676 B.n373 163.367
R1507 B.n680 B.n373 163.367
R1508 B.n680 B.n367 163.367
R1509 B.n688 B.n367 163.367
R1510 B.n688 B.n365 163.367
R1511 B.n692 B.n365 163.367
R1512 B.n692 B.n359 163.367
R1513 B.n700 B.n359 163.367
R1514 B.n700 B.n357 163.367
R1515 B.n704 B.n357 163.367
R1516 B.n704 B.n351 163.367
R1517 B.n712 B.n351 163.367
R1518 B.n712 B.n349 163.367
R1519 B.n716 B.n349 163.367
R1520 B.n716 B.n343 163.367
R1521 B.n724 B.n343 163.367
R1522 B.n724 B.n341 163.367
R1523 B.n728 B.n341 163.367
R1524 B.n728 B.n335 163.367
R1525 B.n737 B.n335 163.367
R1526 B.n737 B.n333 163.367
R1527 B.n741 B.n333 163.367
R1528 B.n741 B.n328 163.367
R1529 B.n750 B.n328 163.367
R1530 B.n750 B.n326 163.367
R1531 B.n754 B.n326 163.367
R1532 B.n754 B.n2 163.367
R1533 B.n881 B.n2 163.367
R1534 B.n881 B.n3 163.367
R1535 B.n877 B.n3 163.367
R1536 B.n877 B.n9 163.367
R1537 B.n873 B.n9 163.367
R1538 B.n873 B.n11 163.367
R1539 B.n869 B.n11 163.367
R1540 B.n869 B.n15 163.367
R1541 B.n865 B.n15 163.367
R1542 B.n865 B.n17 163.367
R1543 B.n861 B.n17 163.367
R1544 B.n861 B.n23 163.367
R1545 B.n857 B.n23 163.367
R1546 B.n857 B.n25 163.367
R1547 B.n853 B.n25 163.367
R1548 B.n853 B.n30 163.367
R1549 B.n849 B.n30 163.367
R1550 B.n849 B.n32 163.367
R1551 B.n845 B.n32 163.367
R1552 B.n845 B.n37 163.367
R1553 B.n841 B.n37 163.367
R1554 B.n841 B.n39 163.367
R1555 B.n837 B.n39 163.367
R1556 B.n837 B.n44 163.367
R1557 B.n833 B.n44 163.367
R1558 B.n833 B.n46 163.367
R1559 B.n829 B.n46 163.367
R1560 B.n829 B.n51 163.367
R1561 B.n825 B.n51 163.367
R1562 B.n825 B.n53 163.367
R1563 B.n821 B.n53 163.367
R1564 B.n821 B.n58 163.367
R1565 B.n817 B.n58 163.367
R1566 B.n817 B.n60 163.367
R1567 B.n813 B.n60 163.367
R1568 B.n813 B.n65 163.367
R1569 B.n809 B.n65 163.367
R1570 B.n449 B.n448 163.367
R1571 B.n451 B.n449 163.367
R1572 B.n455 B.n444 163.367
R1573 B.n459 B.n457 163.367
R1574 B.n463 B.n442 163.367
R1575 B.n467 B.n465 163.367
R1576 B.n471 B.n440 163.367
R1577 B.n475 B.n473 163.367
R1578 B.n479 B.n438 163.367
R1579 B.n483 B.n481 163.367
R1580 B.n487 B.n436 163.367
R1581 B.n491 B.n489 163.367
R1582 B.n495 B.n434 163.367
R1583 B.n499 B.n497 163.367
R1584 B.n503 B.n432 163.367
R1585 B.n507 B.n505 163.367
R1586 B.n511 B.n430 163.367
R1587 B.n515 B.n513 163.367
R1588 B.n519 B.n428 163.367
R1589 B.n523 B.n521 163.367
R1590 B.n527 B.n426 163.367
R1591 B.n531 B.n529 163.367
R1592 B.n538 B.n424 163.367
R1593 B.n542 B.n540 163.367
R1594 B.n546 B.n422 163.367
R1595 B.n550 B.n548 163.367
R1596 B.n554 B.n420 163.367
R1597 B.n558 B.n556 163.367
R1598 B.n562 B.n415 163.367
R1599 B.n566 B.n564 163.367
R1600 B.n570 B.n413 163.367
R1601 B.n574 B.n572 163.367
R1602 B.n578 B.n411 163.367
R1603 B.n582 B.n580 163.367
R1604 B.n586 B.n409 163.367
R1605 B.n590 B.n588 163.367
R1606 B.n594 B.n407 163.367
R1607 B.n598 B.n596 163.367
R1608 B.n602 B.n405 163.367
R1609 B.n606 B.n604 163.367
R1610 B.n610 B.n403 163.367
R1611 B.n614 B.n612 163.367
R1612 B.n618 B.n401 163.367
R1613 B.n622 B.n620 163.367
R1614 B.n626 B.n399 163.367
R1615 B.n630 B.n628 163.367
R1616 B.n634 B.n397 163.367
R1617 B.n638 B.n636 163.367
R1618 B.n642 B.n395 163.367
R1619 B.n646 B.n644 163.367
R1620 B.n650 B.n387 163.367
R1621 B.n658 B.n387 163.367
R1622 B.n658 B.n385 163.367
R1623 B.n662 B.n385 163.367
R1624 B.n662 B.n379 163.367
R1625 B.n670 B.n379 163.367
R1626 B.n670 B.n377 163.367
R1627 B.n674 B.n377 163.367
R1628 B.n674 B.n371 163.367
R1629 B.n682 B.n371 163.367
R1630 B.n682 B.n369 163.367
R1631 B.n686 B.n369 163.367
R1632 B.n686 B.n363 163.367
R1633 B.n694 B.n363 163.367
R1634 B.n694 B.n361 163.367
R1635 B.n698 B.n361 163.367
R1636 B.n698 B.n355 163.367
R1637 B.n706 B.n355 163.367
R1638 B.n706 B.n353 163.367
R1639 B.n710 B.n353 163.367
R1640 B.n710 B.n347 163.367
R1641 B.n718 B.n347 163.367
R1642 B.n718 B.n345 163.367
R1643 B.n722 B.n345 163.367
R1644 B.n722 B.n339 163.367
R1645 B.n730 B.n339 163.367
R1646 B.n730 B.n337 163.367
R1647 B.n734 B.n337 163.367
R1648 B.n734 B.n332 163.367
R1649 B.n743 B.n332 163.367
R1650 B.n743 B.n330 163.367
R1651 B.n748 B.n330 163.367
R1652 B.n748 B.n324 163.367
R1653 B.n756 B.n324 163.367
R1654 B.n757 B.n756 163.367
R1655 B.n757 B.n5 163.367
R1656 B.n6 B.n5 163.367
R1657 B.n7 B.n6 163.367
R1658 B.n762 B.n7 163.367
R1659 B.n762 B.n12 163.367
R1660 B.n13 B.n12 163.367
R1661 B.n14 B.n13 163.367
R1662 B.n767 B.n14 163.367
R1663 B.n767 B.n19 163.367
R1664 B.n20 B.n19 163.367
R1665 B.n21 B.n20 163.367
R1666 B.n772 B.n21 163.367
R1667 B.n772 B.n26 163.367
R1668 B.n27 B.n26 163.367
R1669 B.n28 B.n27 163.367
R1670 B.n777 B.n28 163.367
R1671 B.n777 B.n33 163.367
R1672 B.n34 B.n33 163.367
R1673 B.n35 B.n34 163.367
R1674 B.n782 B.n35 163.367
R1675 B.n782 B.n40 163.367
R1676 B.n41 B.n40 163.367
R1677 B.n42 B.n41 163.367
R1678 B.n787 B.n42 163.367
R1679 B.n787 B.n47 163.367
R1680 B.n48 B.n47 163.367
R1681 B.n49 B.n48 163.367
R1682 B.n792 B.n49 163.367
R1683 B.n792 B.n54 163.367
R1684 B.n55 B.n54 163.367
R1685 B.n56 B.n55 163.367
R1686 B.n797 B.n56 163.367
R1687 B.n797 B.n61 163.367
R1688 B.n62 B.n61 163.367
R1689 B.n63 B.n62 163.367
R1690 B.n802 B.n63 163.367
R1691 B.n802 B.n68 163.367
R1692 B.n127 B.n126 163.367
R1693 B.n131 B.n130 163.367
R1694 B.n135 B.n134 163.367
R1695 B.n139 B.n138 163.367
R1696 B.n143 B.n142 163.367
R1697 B.n147 B.n146 163.367
R1698 B.n151 B.n150 163.367
R1699 B.n155 B.n154 163.367
R1700 B.n159 B.n158 163.367
R1701 B.n163 B.n162 163.367
R1702 B.n167 B.n166 163.367
R1703 B.n171 B.n170 163.367
R1704 B.n175 B.n174 163.367
R1705 B.n179 B.n178 163.367
R1706 B.n183 B.n182 163.367
R1707 B.n187 B.n186 163.367
R1708 B.n191 B.n190 163.367
R1709 B.n195 B.n194 163.367
R1710 B.n199 B.n198 163.367
R1711 B.n203 B.n202 163.367
R1712 B.n207 B.n206 163.367
R1713 B.n211 B.n210 163.367
R1714 B.n215 B.n214 163.367
R1715 B.n219 B.n218 163.367
R1716 B.n223 B.n222 163.367
R1717 B.n227 B.n226 163.367
R1718 B.n231 B.n230 163.367
R1719 B.n236 B.n235 163.367
R1720 B.n240 B.n239 163.367
R1721 B.n244 B.n243 163.367
R1722 B.n248 B.n247 163.367
R1723 B.n252 B.n251 163.367
R1724 B.n256 B.n255 163.367
R1725 B.n260 B.n259 163.367
R1726 B.n264 B.n263 163.367
R1727 B.n268 B.n267 163.367
R1728 B.n272 B.n271 163.367
R1729 B.n276 B.n275 163.367
R1730 B.n280 B.n279 163.367
R1731 B.n284 B.n283 163.367
R1732 B.n288 B.n287 163.367
R1733 B.n292 B.n291 163.367
R1734 B.n296 B.n295 163.367
R1735 B.n300 B.n299 163.367
R1736 B.n304 B.n303 163.367
R1737 B.n308 B.n307 163.367
R1738 B.n312 B.n311 163.367
R1739 B.n316 B.n315 163.367
R1740 B.n320 B.n319 163.367
R1741 B.n806 B.n119 163.367
R1742 B.n447 B.n391 71.676
R1743 B.n451 B.n450 71.676
R1744 B.n456 B.n455 71.676
R1745 B.n459 B.n458 71.676
R1746 B.n464 B.n463 71.676
R1747 B.n467 B.n466 71.676
R1748 B.n472 B.n471 71.676
R1749 B.n475 B.n474 71.676
R1750 B.n480 B.n479 71.676
R1751 B.n483 B.n482 71.676
R1752 B.n488 B.n487 71.676
R1753 B.n491 B.n490 71.676
R1754 B.n496 B.n495 71.676
R1755 B.n499 B.n498 71.676
R1756 B.n504 B.n503 71.676
R1757 B.n507 B.n506 71.676
R1758 B.n512 B.n511 71.676
R1759 B.n515 B.n514 71.676
R1760 B.n520 B.n519 71.676
R1761 B.n523 B.n522 71.676
R1762 B.n528 B.n527 71.676
R1763 B.n531 B.n530 71.676
R1764 B.n539 B.n538 71.676
R1765 B.n542 B.n541 71.676
R1766 B.n547 B.n546 71.676
R1767 B.n550 B.n549 71.676
R1768 B.n555 B.n554 71.676
R1769 B.n558 B.n557 71.676
R1770 B.n563 B.n562 71.676
R1771 B.n566 B.n565 71.676
R1772 B.n571 B.n570 71.676
R1773 B.n574 B.n573 71.676
R1774 B.n579 B.n578 71.676
R1775 B.n582 B.n581 71.676
R1776 B.n587 B.n586 71.676
R1777 B.n590 B.n589 71.676
R1778 B.n595 B.n594 71.676
R1779 B.n598 B.n597 71.676
R1780 B.n603 B.n602 71.676
R1781 B.n606 B.n605 71.676
R1782 B.n611 B.n610 71.676
R1783 B.n614 B.n613 71.676
R1784 B.n619 B.n618 71.676
R1785 B.n622 B.n621 71.676
R1786 B.n627 B.n626 71.676
R1787 B.n630 B.n629 71.676
R1788 B.n635 B.n634 71.676
R1789 B.n638 B.n637 71.676
R1790 B.n643 B.n642 71.676
R1791 B.n646 B.n645 71.676
R1792 B.n69 B.n67 71.676
R1793 B.n127 B.n70 71.676
R1794 B.n131 B.n71 71.676
R1795 B.n135 B.n72 71.676
R1796 B.n139 B.n73 71.676
R1797 B.n143 B.n74 71.676
R1798 B.n147 B.n75 71.676
R1799 B.n151 B.n76 71.676
R1800 B.n155 B.n77 71.676
R1801 B.n159 B.n78 71.676
R1802 B.n163 B.n79 71.676
R1803 B.n167 B.n80 71.676
R1804 B.n171 B.n81 71.676
R1805 B.n175 B.n82 71.676
R1806 B.n179 B.n83 71.676
R1807 B.n183 B.n84 71.676
R1808 B.n187 B.n85 71.676
R1809 B.n191 B.n86 71.676
R1810 B.n195 B.n87 71.676
R1811 B.n199 B.n88 71.676
R1812 B.n203 B.n89 71.676
R1813 B.n207 B.n90 71.676
R1814 B.n211 B.n91 71.676
R1815 B.n215 B.n92 71.676
R1816 B.n219 B.n93 71.676
R1817 B.n223 B.n94 71.676
R1818 B.n227 B.n95 71.676
R1819 B.n231 B.n96 71.676
R1820 B.n236 B.n97 71.676
R1821 B.n240 B.n98 71.676
R1822 B.n244 B.n99 71.676
R1823 B.n248 B.n100 71.676
R1824 B.n252 B.n101 71.676
R1825 B.n256 B.n102 71.676
R1826 B.n260 B.n103 71.676
R1827 B.n264 B.n104 71.676
R1828 B.n268 B.n105 71.676
R1829 B.n272 B.n106 71.676
R1830 B.n276 B.n107 71.676
R1831 B.n280 B.n108 71.676
R1832 B.n284 B.n109 71.676
R1833 B.n288 B.n110 71.676
R1834 B.n292 B.n111 71.676
R1835 B.n296 B.n112 71.676
R1836 B.n300 B.n113 71.676
R1837 B.n304 B.n114 71.676
R1838 B.n308 B.n115 71.676
R1839 B.n312 B.n116 71.676
R1840 B.n316 B.n117 71.676
R1841 B.n320 B.n118 71.676
R1842 B.n119 B.n118 71.676
R1843 B.n319 B.n117 71.676
R1844 B.n315 B.n116 71.676
R1845 B.n311 B.n115 71.676
R1846 B.n307 B.n114 71.676
R1847 B.n303 B.n113 71.676
R1848 B.n299 B.n112 71.676
R1849 B.n295 B.n111 71.676
R1850 B.n291 B.n110 71.676
R1851 B.n287 B.n109 71.676
R1852 B.n283 B.n108 71.676
R1853 B.n279 B.n107 71.676
R1854 B.n275 B.n106 71.676
R1855 B.n271 B.n105 71.676
R1856 B.n267 B.n104 71.676
R1857 B.n263 B.n103 71.676
R1858 B.n259 B.n102 71.676
R1859 B.n255 B.n101 71.676
R1860 B.n251 B.n100 71.676
R1861 B.n247 B.n99 71.676
R1862 B.n243 B.n98 71.676
R1863 B.n239 B.n97 71.676
R1864 B.n235 B.n96 71.676
R1865 B.n230 B.n95 71.676
R1866 B.n226 B.n94 71.676
R1867 B.n222 B.n93 71.676
R1868 B.n218 B.n92 71.676
R1869 B.n214 B.n91 71.676
R1870 B.n210 B.n90 71.676
R1871 B.n206 B.n89 71.676
R1872 B.n202 B.n88 71.676
R1873 B.n198 B.n87 71.676
R1874 B.n194 B.n86 71.676
R1875 B.n190 B.n85 71.676
R1876 B.n186 B.n84 71.676
R1877 B.n182 B.n83 71.676
R1878 B.n178 B.n82 71.676
R1879 B.n174 B.n81 71.676
R1880 B.n170 B.n80 71.676
R1881 B.n166 B.n79 71.676
R1882 B.n162 B.n78 71.676
R1883 B.n158 B.n77 71.676
R1884 B.n154 B.n76 71.676
R1885 B.n150 B.n75 71.676
R1886 B.n146 B.n74 71.676
R1887 B.n142 B.n73 71.676
R1888 B.n138 B.n72 71.676
R1889 B.n134 B.n71 71.676
R1890 B.n130 B.n70 71.676
R1891 B.n126 B.n69 71.676
R1892 B.n448 B.n447 71.676
R1893 B.n450 B.n444 71.676
R1894 B.n457 B.n456 71.676
R1895 B.n458 B.n442 71.676
R1896 B.n465 B.n464 71.676
R1897 B.n466 B.n440 71.676
R1898 B.n473 B.n472 71.676
R1899 B.n474 B.n438 71.676
R1900 B.n481 B.n480 71.676
R1901 B.n482 B.n436 71.676
R1902 B.n489 B.n488 71.676
R1903 B.n490 B.n434 71.676
R1904 B.n497 B.n496 71.676
R1905 B.n498 B.n432 71.676
R1906 B.n505 B.n504 71.676
R1907 B.n506 B.n430 71.676
R1908 B.n513 B.n512 71.676
R1909 B.n514 B.n428 71.676
R1910 B.n521 B.n520 71.676
R1911 B.n522 B.n426 71.676
R1912 B.n529 B.n528 71.676
R1913 B.n530 B.n424 71.676
R1914 B.n540 B.n539 71.676
R1915 B.n541 B.n422 71.676
R1916 B.n548 B.n547 71.676
R1917 B.n549 B.n420 71.676
R1918 B.n556 B.n555 71.676
R1919 B.n557 B.n415 71.676
R1920 B.n564 B.n563 71.676
R1921 B.n565 B.n413 71.676
R1922 B.n572 B.n571 71.676
R1923 B.n573 B.n411 71.676
R1924 B.n580 B.n579 71.676
R1925 B.n581 B.n409 71.676
R1926 B.n588 B.n587 71.676
R1927 B.n589 B.n407 71.676
R1928 B.n596 B.n595 71.676
R1929 B.n597 B.n405 71.676
R1930 B.n604 B.n603 71.676
R1931 B.n605 B.n403 71.676
R1932 B.n612 B.n611 71.676
R1933 B.n613 B.n401 71.676
R1934 B.n620 B.n619 71.676
R1935 B.n621 B.n399 71.676
R1936 B.n628 B.n627 71.676
R1937 B.n629 B.n397 71.676
R1938 B.n636 B.n635 71.676
R1939 B.n637 B.n395 71.676
R1940 B.n644 B.n643 71.676
R1941 B.n645 B.n393 71.676
R1942 B.n651 B.n392 69.1383
R1943 B.n808 B.n807 69.1383
R1944 B.n417 B.n416 61.0914
R1945 B.n535 B.n534 61.0914
R1946 B.n123 B.n122 61.0914
R1947 B.n121 B.n120 61.0914
R1948 B.n418 B.n417 59.5399
R1949 B.n536 B.n535 59.5399
R1950 B.n124 B.n123 59.5399
R1951 B.n233 B.n121 59.5399
R1952 B.n651 B.n388 40.1831
R1953 B.n657 B.n388 40.1831
R1954 B.n657 B.n384 40.1831
R1955 B.n663 B.n384 40.1831
R1956 B.n663 B.n380 40.1831
R1957 B.n669 B.n380 40.1831
R1958 B.n669 B.n376 40.1831
R1959 B.n675 B.n376 40.1831
R1960 B.n681 B.n372 40.1831
R1961 B.n681 B.n368 40.1831
R1962 B.n687 B.n368 40.1831
R1963 B.n687 B.n364 40.1831
R1964 B.n693 B.n364 40.1831
R1965 B.n693 B.n360 40.1831
R1966 B.n699 B.n360 40.1831
R1967 B.n699 B.n356 40.1831
R1968 B.n705 B.n356 40.1831
R1969 B.n705 B.n352 40.1831
R1970 B.n711 B.n352 40.1831
R1971 B.n717 B.n348 40.1831
R1972 B.n717 B.n344 40.1831
R1973 B.n723 B.n344 40.1831
R1974 B.n723 B.n340 40.1831
R1975 B.n729 B.n340 40.1831
R1976 B.n729 B.n336 40.1831
R1977 B.n736 B.n336 40.1831
R1978 B.n736 B.n735 40.1831
R1979 B.n742 B.n329 40.1831
R1980 B.n749 B.n329 40.1831
R1981 B.n749 B.n325 40.1831
R1982 B.n755 B.n325 40.1831
R1983 B.n755 B.n4 40.1831
R1984 B.n880 B.n4 40.1831
R1985 B.n880 B.n879 40.1831
R1986 B.n879 B.n878 40.1831
R1987 B.n878 B.n8 40.1831
R1988 B.n872 B.n8 40.1831
R1989 B.n872 B.n871 40.1831
R1990 B.n871 B.n870 40.1831
R1991 B.n864 B.n18 40.1831
R1992 B.n864 B.n863 40.1831
R1993 B.n863 B.n862 40.1831
R1994 B.n862 B.n22 40.1831
R1995 B.n856 B.n22 40.1831
R1996 B.n856 B.n855 40.1831
R1997 B.n855 B.n854 40.1831
R1998 B.n854 B.n29 40.1831
R1999 B.n848 B.n847 40.1831
R2000 B.n847 B.n846 40.1831
R2001 B.n846 B.n36 40.1831
R2002 B.n840 B.n36 40.1831
R2003 B.n840 B.n839 40.1831
R2004 B.n839 B.n838 40.1831
R2005 B.n838 B.n43 40.1831
R2006 B.n832 B.n43 40.1831
R2007 B.n832 B.n831 40.1831
R2008 B.n831 B.n830 40.1831
R2009 B.n830 B.n50 40.1831
R2010 B.n824 B.n823 40.1831
R2011 B.n823 B.n822 40.1831
R2012 B.n822 B.n57 40.1831
R2013 B.n816 B.n57 40.1831
R2014 B.n816 B.n815 40.1831
R2015 B.n815 B.n814 40.1831
R2016 B.n814 B.n64 40.1831
R2017 B.n808 B.n64 40.1831
R2018 B.t9 B.n372 39.0013
R2019 B.t5 B.n50 39.0013
R2020 B.n735 B.t3 30.7284
R2021 B.n18 B.t2 30.7284
R2022 B.n810 B.n66 29.8151
R2023 B.n805 B.n804 29.8151
R2024 B.n649 B.n648 29.8151
R2025 B.n653 B.n390 29.8151
R2026 B.n711 B.t0 20.0918
R2027 B.t0 B.n348 20.0918
R2028 B.t1 B.n29 20.0918
R2029 B.n848 B.t1 20.0918
R2030 B B.n882 18.0485
R2031 B.n125 B.n66 10.6151
R2032 B.n128 B.n125 10.6151
R2033 B.n129 B.n128 10.6151
R2034 B.n132 B.n129 10.6151
R2035 B.n133 B.n132 10.6151
R2036 B.n136 B.n133 10.6151
R2037 B.n137 B.n136 10.6151
R2038 B.n140 B.n137 10.6151
R2039 B.n141 B.n140 10.6151
R2040 B.n144 B.n141 10.6151
R2041 B.n145 B.n144 10.6151
R2042 B.n148 B.n145 10.6151
R2043 B.n149 B.n148 10.6151
R2044 B.n152 B.n149 10.6151
R2045 B.n153 B.n152 10.6151
R2046 B.n156 B.n153 10.6151
R2047 B.n157 B.n156 10.6151
R2048 B.n160 B.n157 10.6151
R2049 B.n161 B.n160 10.6151
R2050 B.n164 B.n161 10.6151
R2051 B.n165 B.n164 10.6151
R2052 B.n168 B.n165 10.6151
R2053 B.n169 B.n168 10.6151
R2054 B.n172 B.n169 10.6151
R2055 B.n173 B.n172 10.6151
R2056 B.n176 B.n173 10.6151
R2057 B.n177 B.n176 10.6151
R2058 B.n180 B.n177 10.6151
R2059 B.n181 B.n180 10.6151
R2060 B.n184 B.n181 10.6151
R2061 B.n185 B.n184 10.6151
R2062 B.n188 B.n185 10.6151
R2063 B.n189 B.n188 10.6151
R2064 B.n192 B.n189 10.6151
R2065 B.n193 B.n192 10.6151
R2066 B.n196 B.n193 10.6151
R2067 B.n197 B.n196 10.6151
R2068 B.n200 B.n197 10.6151
R2069 B.n201 B.n200 10.6151
R2070 B.n204 B.n201 10.6151
R2071 B.n205 B.n204 10.6151
R2072 B.n208 B.n205 10.6151
R2073 B.n209 B.n208 10.6151
R2074 B.n212 B.n209 10.6151
R2075 B.n213 B.n212 10.6151
R2076 B.n217 B.n216 10.6151
R2077 B.n220 B.n217 10.6151
R2078 B.n221 B.n220 10.6151
R2079 B.n224 B.n221 10.6151
R2080 B.n225 B.n224 10.6151
R2081 B.n228 B.n225 10.6151
R2082 B.n229 B.n228 10.6151
R2083 B.n232 B.n229 10.6151
R2084 B.n237 B.n234 10.6151
R2085 B.n238 B.n237 10.6151
R2086 B.n241 B.n238 10.6151
R2087 B.n242 B.n241 10.6151
R2088 B.n245 B.n242 10.6151
R2089 B.n246 B.n245 10.6151
R2090 B.n249 B.n246 10.6151
R2091 B.n250 B.n249 10.6151
R2092 B.n253 B.n250 10.6151
R2093 B.n254 B.n253 10.6151
R2094 B.n257 B.n254 10.6151
R2095 B.n258 B.n257 10.6151
R2096 B.n261 B.n258 10.6151
R2097 B.n262 B.n261 10.6151
R2098 B.n265 B.n262 10.6151
R2099 B.n266 B.n265 10.6151
R2100 B.n269 B.n266 10.6151
R2101 B.n270 B.n269 10.6151
R2102 B.n273 B.n270 10.6151
R2103 B.n274 B.n273 10.6151
R2104 B.n277 B.n274 10.6151
R2105 B.n278 B.n277 10.6151
R2106 B.n281 B.n278 10.6151
R2107 B.n282 B.n281 10.6151
R2108 B.n285 B.n282 10.6151
R2109 B.n286 B.n285 10.6151
R2110 B.n289 B.n286 10.6151
R2111 B.n290 B.n289 10.6151
R2112 B.n293 B.n290 10.6151
R2113 B.n294 B.n293 10.6151
R2114 B.n297 B.n294 10.6151
R2115 B.n298 B.n297 10.6151
R2116 B.n301 B.n298 10.6151
R2117 B.n302 B.n301 10.6151
R2118 B.n305 B.n302 10.6151
R2119 B.n306 B.n305 10.6151
R2120 B.n309 B.n306 10.6151
R2121 B.n310 B.n309 10.6151
R2122 B.n313 B.n310 10.6151
R2123 B.n314 B.n313 10.6151
R2124 B.n317 B.n314 10.6151
R2125 B.n318 B.n317 10.6151
R2126 B.n321 B.n318 10.6151
R2127 B.n322 B.n321 10.6151
R2128 B.n805 B.n322 10.6151
R2129 B.n649 B.n386 10.6151
R2130 B.n659 B.n386 10.6151
R2131 B.n660 B.n659 10.6151
R2132 B.n661 B.n660 10.6151
R2133 B.n661 B.n378 10.6151
R2134 B.n671 B.n378 10.6151
R2135 B.n672 B.n671 10.6151
R2136 B.n673 B.n672 10.6151
R2137 B.n673 B.n370 10.6151
R2138 B.n683 B.n370 10.6151
R2139 B.n684 B.n683 10.6151
R2140 B.n685 B.n684 10.6151
R2141 B.n685 B.n362 10.6151
R2142 B.n695 B.n362 10.6151
R2143 B.n696 B.n695 10.6151
R2144 B.n697 B.n696 10.6151
R2145 B.n697 B.n354 10.6151
R2146 B.n707 B.n354 10.6151
R2147 B.n708 B.n707 10.6151
R2148 B.n709 B.n708 10.6151
R2149 B.n709 B.n346 10.6151
R2150 B.n719 B.n346 10.6151
R2151 B.n720 B.n719 10.6151
R2152 B.n721 B.n720 10.6151
R2153 B.n721 B.n338 10.6151
R2154 B.n731 B.n338 10.6151
R2155 B.n732 B.n731 10.6151
R2156 B.n733 B.n732 10.6151
R2157 B.n733 B.n331 10.6151
R2158 B.n744 B.n331 10.6151
R2159 B.n745 B.n744 10.6151
R2160 B.n747 B.n745 10.6151
R2161 B.n747 B.n746 10.6151
R2162 B.n746 B.n323 10.6151
R2163 B.n758 B.n323 10.6151
R2164 B.n759 B.n758 10.6151
R2165 B.n760 B.n759 10.6151
R2166 B.n761 B.n760 10.6151
R2167 B.n763 B.n761 10.6151
R2168 B.n764 B.n763 10.6151
R2169 B.n765 B.n764 10.6151
R2170 B.n766 B.n765 10.6151
R2171 B.n768 B.n766 10.6151
R2172 B.n769 B.n768 10.6151
R2173 B.n770 B.n769 10.6151
R2174 B.n771 B.n770 10.6151
R2175 B.n773 B.n771 10.6151
R2176 B.n774 B.n773 10.6151
R2177 B.n775 B.n774 10.6151
R2178 B.n776 B.n775 10.6151
R2179 B.n778 B.n776 10.6151
R2180 B.n779 B.n778 10.6151
R2181 B.n780 B.n779 10.6151
R2182 B.n781 B.n780 10.6151
R2183 B.n783 B.n781 10.6151
R2184 B.n784 B.n783 10.6151
R2185 B.n785 B.n784 10.6151
R2186 B.n786 B.n785 10.6151
R2187 B.n788 B.n786 10.6151
R2188 B.n789 B.n788 10.6151
R2189 B.n790 B.n789 10.6151
R2190 B.n791 B.n790 10.6151
R2191 B.n793 B.n791 10.6151
R2192 B.n794 B.n793 10.6151
R2193 B.n795 B.n794 10.6151
R2194 B.n796 B.n795 10.6151
R2195 B.n798 B.n796 10.6151
R2196 B.n799 B.n798 10.6151
R2197 B.n800 B.n799 10.6151
R2198 B.n801 B.n800 10.6151
R2199 B.n803 B.n801 10.6151
R2200 B.n804 B.n803 10.6151
R2201 B.n446 B.n390 10.6151
R2202 B.n446 B.n445 10.6151
R2203 B.n452 B.n445 10.6151
R2204 B.n453 B.n452 10.6151
R2205 B.n454 B.n453 10.6151
R2206 B.n454 B.n443 10.6151
R2207 B.n460 B.n443 10.6151
R2208 B.n461 B.n460 10.6151
R2209 B.n462 B.n461 10.6151
R2210 B.n462 B.n441 10.6151
R2211 B.n468 B.n441 10.6151
R2212 B.n469 B.n468 10.6151
R2213 B.n470 B.n469 10.6151
R2214 B.n470 B.n439 10.6151
R2215 B.n476 B.n439 10.6151
R2216 B.n477 B.n476 10.6151
R2217 B.n478 B.n477 10.6151
R2218 B.n478 B.n437 10.6151
R2219 B.n484 B.n437 10.6151
R2220 B.n485 B.n484 10.6151
R2221 B.n486 B.n485 10.6151
R2222 B.n486 B.n435 10.6151
R2223 B.n492 B.n435 10.6151
R2224 B.n493 B.n492 10.6151
R2225 B.n494 B.n493 10.6151
R2226 B.n494 B.n433 10.6151
R2227 B.n500 B.n433 10.6151
R2228 B.n501 B.n500 10.6151
R2229 B.n502 B.n501 10.6151
R2230 B.n502 B.n431 10.6151
R2231 B.n508 B.n431 10.6151
R2232 B.n509 B.n508 10.6151
R2233 B.n510 B.n509 10.6151
R2234 B.n510 B.n429 10.6151
R2235 B.n516 B.n429 10.6151
R2236 B.n517 B.n516 10.6151
R2237 B.n518 B.n517 10.6151
R2238 B.n518 B.n427 10.6151
R2239 B.n524 B.n427 10.6151
R2240 B.n525 B.n524 10.6151
R2241 B.n526 B.n525 10.6151
R2242 B.n526 B.n425 10.6151
R2243 B.n532 B.n425 10.6151
R2244 B.n533 B.n532 10.6151
R2245 B.n537 B.n533 10.6151
R2246 B.n543 B.n423 10.6151
R2247 B.n544 B.n543 10.6151
R2248 B.n545 B.n544 10.6151
R2249 B.n545 B.n421 10.6151
R2250 B.n551 B.n421 10.6151
R2251 B.n552 B.n551 10.6151
R2252 B.n553 B.n552 10.6151
R2253 B.n553 B.n419 10.6151
R2254 B.n560 B.n559 10.6151
R2255 B.n561 B.n560 10.6151
R2256 B.n561 B.n414 10.6151
R2257 B.n567 B.n414 10.6151
R2258 B.n568 B.n567 10.6151
R2259 B.n569 B.n568 10.6151
R2260 B.n569 B.n412 10.6151
R2261 B.n575 B.n412 10.6151
R2262 B.n576 B.n575 10.6151
R2263 B.n577 B.n576 10.6151
R2264 B.n577 B.n410 10.6151
R2265 B.n583 B.n410 10.6151
R2266 B.n584 B.n583 10.6151
R2267 B.n585 B.n584 10.6151
R2268 B.n585 B.n408 10.6151
R2269 B.n591 B.n408 10.6151
R2270 B.n592 B.n591 10.6151
R2271 B.n593 B.n592 10.6151
R2272 B.n593 B.n406 10.6151
R2273 B.n599 B.n406 10.6151
R2274 B.n600 B.n599 10.6151
R2275 B.n601 B.n600 10.6151
R2276 B.n601 B.n404 10.6151
R2277 B.n607 B.n404 10.6151
R2278 B.n608 B.n607 10.6151
R2279 B.n609 B.n608 10.6151
R2280 B.n609 B.n402 10.6151
R2281 B.n615 B.n402 10.6151
R2282 B.n616 B.n615 10.6151
R2283 B.n617 B.n616 10.6151
R2284 B.n617 B.n400 10.6151
R2285 B.n623 B.n400 10.6151
R2286 B.n624 B.n623 10.6151
R2287 B.n625 B.n624 10.6151
R2288 B.n625 B.n398 10.6151
R2289 B.n631 B.n398 10.6151
R2290 B.n632 B.n631 10.6151
R2291 B.n633 B.n632 10.6151
R2292 B.n633 B.n396 10.6151
R2293 B.n639 B.n396 10.6151
R2294 B.n640 B.n639 10.6151
R2295 B.n641 B.n640 10.6151
R2296 B.n641 B.n394 10.6151
R2297 B.n647 B.n394 10.6151
R2298 B.n648 B.n647 10.6151
R2299 B.n654 B.n653 10.6151
R2300 B.n655 B.n654 10.6151
R2301 B.n655 B.n382 10.6151
R2302 B.n665 B.n382 10.6151
R2303 B.n666 B.n665 10.6151
R2304 B.n667 B.n666 10.6151
R2305 B.n667 B.n374 10.6151
R2306 B.n677 B.n374 10.6151
R2307 B.n678 B.n677 10.6151
R2308 B.n679 B.n678 10.6151
R2309 B.n679 B.n366 10.6151
R2310 B.n689 B.n366 10.6151
R2311 B.n690 B.n689 10.6151
R2312 B.n691 B.n690 10.6151
R2313 B.n691 B.n358 10.6151
R2314 B.n701 B.n358 10.6151
R2315 B.n702 B.n701 10.6151
R2316 B.n703 B.n702 10.6151
R2317 B.n703 B.n350 10.6151
R2318 B.n713 B.n350 10.6151
R2319 B.n714 B.n713 10.6151
R2320 B.n715 B.n714 10.6151
R2321 B.n715 B.n342 10.6151
R2322 B.n725 B.n342 10.6151
R2323 B.n726 B.n725 10.6151
R2324 B.n727 B.n726 10.6151
R2325 B.n727 B.n334 10.6151
R2326 B.n738 B.n334 10.6151
R2327 B.n739 B.n738 10.6151
R2328 B.n740 B.n739 10.6151
R2329 B.n740 B.n327 10.6151
R2330 B.n751 B.n327 10.6151
R2331 B.n752 B.n751 10.6151
R2332 B.n753 B.n752 10.6151
R2333 B.n753 B.n0 10.6151
R2334 B.n876 B.n1 10.6151
R2335 B.n876 B.n875 10.6151
R2336 B.n875 B.n874 10.6151
R2337 B.n874 B.n10 10.6151
R2338 B.n868 B.n10 10.6151
R2339 B.n868 B.n867 10.6151
R2340 B.n867 B.n866 10.6151
R2341 B.n866 B.n16 10.6151
R2342 B.n860 B.n16 10.6151
R2343 B.n860 B.n859 10.6151
R2344 B.n859 B.n858 10.6151
R2345 B.n858 B.n24 10.6151
R2346 B.n852 B.n24 10.6151
R2347 B.n852 B.n851 10.6151
R2348 B.n851 B.n850 10.6151
R2349 B.n850 B.n31 10.6151
R2350 B.n844 B.n31 10.6151
R2351 B.n844 B.n843 10.6151
R2352 B.n843 B.n842 10.6151
R2353 B.n842 B.n38 10.6151
R2354 B.n836 B.n38 10.6151
R2355 B.n836 B.n835 10.6151
R2356 B.n835 B.n834 10.6151
R2357 B.n834 B.n45 10.6151
R2358 B.n828 B.n45 10.6151
R2359 B.n828 B.n827 10.6151
R2360 B.n827 B.n826 10.6151
R2361 B.n826 B.n52 10.6151
R2362 B.n820 B.n52 10.6151
R2363 B.n820 B.n819 10.6151
R2364 B.n819 B.n818 10.6151
R2365 B.n818 B.n59 10.6151
R2366 B.n812 B.n59 10.6151
R2367 B.n812 B.n811 10.6151
R2368 B.n811 B.n810 10.6151
R2369 B.n742 B.t3 9.45524
R2370 B.n870 B.t2 9.45524
R2371 B.n216 B.n124 6.5566
R2372 B.n233 B.n232 6.5566
R2373 B.n536 B.n423 6.5566
R2374 B.n419 B.n418 6.5566
R2375 B.n213 B.n124 4.05904
R2376 B.n234 B.n233 4.05904
R2377 B.n537 B.n536 4.05904
R2378 B.n559 B.n418 4.05904
R2379 B.n882 B.n0 2.81026
R2380 B.n882 B.n1 2.81026
R2381 B.n675 B.t9 1.18234
R2382 B.n824 B.t5 1.18234
R2383 VP.n16 VP.n0 161.3
R2384 VP.n15 VP.n14 161.3
R2385 VP.n13 VP.n1 161.3
R2386 VP.n12 VP.n11 161.3
R2387 VP.n10 VP.n2 161.3
R2388 VP.n9 VP.n8 161.3
R2389 VP.n7 VP.n3 161.3
R2390 VP.n4 VP.t1 149.218
R2391 VP.n4 VP.t2 148.325
R2392 VP.n5 VP.t3 114.005
R2393 VP.n17 VP.t0 114.005
R2394 VP.n6 VP.n5 107.219
R2395 VP.n18 VP.n17 107.219
R2396 VP.n6 VP.n4 51.4577
R2397 VP.n11 VP.n10 40.577
R2398 VP.n11 VP.n1 40.577
R2399 VP.n9 VP.n3 24.5923
R2400 VP.n10 VP.n9 24.5923
R2401 VP.n15 VP.n1 24.5923
R2402 VP.n16 VP.n15 24.5923
R2403 VP.n5 VP.n3 3.68928
R2404 VP.n17 VP.n16 3.68928
R2405 VP.n7 VP.n6 0.278335
R2406 VP.n18 VP.n0 0.278335
R2407 VP.n8 VP.n7 0.189894
R2408 VP.n8 VP.n2 0.189894
R2409 VP.n12 VP.n2 0.189894
R2410 VP.n13 VP.n12 0.189894
R2411 VP.n14 VP.n13 0.189894
R2412 VP.n14 VP.n0 0.189894
R2413 VP VP.n18 0.153485
R2414 VDD1 VDD1.n1 107.721
R2415 VDD1 VDD1.n0 63.8928
R2416 VDD1.n0 VDD1.t2 1.48476
R2417 VDD1.n0 VDD1.t1 1.48476
R2418 VDD1.n1 VDD1.t0 1.48476
R2419 VDD1.n1 VDD1.t3 1.48476
C0 VDD1 VN 0.149371f
C1 VDD2 VP 0.408477f
C2 VDD1 VTAIL 5.75679f
C3 VDD1 VP 5.58279f
C4 VN VTAIL 5.20279f
C5 VP VN 6.59288f
C6 VP VTAIL 5.2169f
C7 VDD1 VDD2 1.07487f
C8 VDD2 VN 5.324471f
C9 VDD2 VTAIL 5.81247f
C10 VDD2 B 3.997682f
C11 VDD1 B 8.38278f
C12 VTAIL B 11.007309f
C13 VN B 11.20776f
C14 VP B 9.486737f
C15 VDD1.t2 B 0.28676f
C16 VDD1.t1 B 0.28676f
C17 VDD1.n0 B 2.58075f
C18 VDD1.t0 B 0.28676f
C19 VDD1.t3 B 0.28676f
C20 VDD1.n1 B 3.33388f
C21 VP.n0 B 0.031962f
C22 VP.t0 B 2.4921f
C23 VP.n1 B 0.047932f
C24 VP.n2 B 0.024244f
C25 VP.n3 B 0.026093f
C26 VP.t2 B 2.73183f
C27 VP.t1 B 2.73787f
C28 VP.n4 B 3.12365f
C29 VP.t3 B 2.4921f
C30 VP.n5 B 0.953678f
C31 VP.n6 B 1.39664f
C32 VP.n7 B 0.031962f
C33 VP.n8 B 0.024244f
C34 VP.n9 B 0.044959f
C35 VP.n10 B 0.047932f
C36 VP.n11 B 0.019581f
C37 VP.n12 B 0.024244f
C38 VP.n13 B 0.024244f
C39 VP.n14 B 0.024244f
C40 VP.n15 B 0.044959f
C41 VP.n16 B 0.026093f
C42 VP.n17 B 0.953678f
C43 VP.n18 B 0.044968f
C44 VTAIL.n0 B 0.022085f
C45 VTAIL.n1 B 0.01623f
C46 VTAIL.n2 B 0.008721f
C47 VTAIL.n3 B 0.020614f
C48 VTAIL.n4 B 0.009234f
C49 VTAIL.n5 B 0.01623f
C50 VTAIL.n6 B 0.008721f
C51 VTAIL.n7 B 0.020614f
C52 VTAIL.n8 B 0.009234f
C53 VTAIL.n9 B 0.01623f
C54 VTAIL.n10 B 0.008721f
C55 VTAIL.n11 B 0.020614f
C56 VTAIL.n12 B 0.009234f
C57 VTAIL.n13 B 0.01623f
C58 VTAIL.n14 B 0.008721f
C59 VTAIL.n15 B 0.020614f
C60 VTAIL.n16 B 0.009234f
C61 VTAIL.n17 B 0.01623f
C62 VTAIL.n18 B 0.008721f
C63 VTAIL.n19 B 0.020614f
C64 VTAIL.n20 B 0.009234f
C65 VTAIL.n21 B 0.932454f
C66 VTAIL.n22 B 0.008721f
C67 VTAIL.t2 B 0.033897f
C68 VTAIL.n23 B 0.099099f
C69 VTAIL.n24 B 0.012177f
C70 VTAIL.n25 B 0.01546f
C71 VTAIL.n26 B 0.020614f
C72 VTAIL.n27 B 0.009234f
C73 VTAIL.n28 B 0.008721f
C74 VTAIL.n29 B 0.01623f
C75 VTAIL.n30 B 0.01623f
C76 VTAIL.n31 B 0.008721f
C77 VTAIL.n32 B 0.009234f
C78 VTAIL.n33 B 0.020614f
C79 VTAIL.n34 B 0.020614f
C80 VTAIL.n35 B 0.009234f
C81 VTAIL.n36 B 0.008721f
C82 VTAIL.n37 B 0.01623f
C83 VTAIL.n38 B 0.01623f
C84 VTAIL.n39 B 0.008721f
C85 VTAIL.n40 B 0.009234f
C86 VTAIL.n41 B 0.020614f
C87 VTAIL.n42 B 0.020614f
C88 VTAIL.n43 B 0.009234f
C89 VTAIL.n44 B 0.008721f
C90 VTAIL.n45 B 0.01623f
C91 VTAIL.n46 B 0.01623f
C92 VTAIL.n47 B 0.008721f
C93 VTAIL.n48 B 0.009234f
C94 VTAIL.n49 B 0.020614f
C95 VTAIL.n50 B 0.020614f
C96 VTAIL.n51 B 0.009234f
C97 VTAIL.n52 B 0.008721f
C98 VTAIL.n53 B 0.01623f
C99 VTAIL.n54 B 0.01623f
C100 VTAIL.n55 B 0.008721f
C101 VTAIL.n56 B 0.009234f
C102 VTAIL.n57 B 0.020614f
C103 VTAIL.n58 B 0.020614f
C104 VTAIL.n59 B 0.009234f
C105 VTAIL.n60 B 0.008721f
C106 VTAIL.n61 B 0.01623f
C107 VTAIL.n62 B 0.01623f
C108 VTAIL.n63 B 0.008721f
C109 VTAIL.n64 B 0.009234f
C110 VTAIL.n65 B 0.020614f
C111 VTAIL.n66 B 0.042081f
C112 VTAIL.n67 B 0.009234f
C113 VTAIL.n68 B 0.017053f
C114 VTAIL.n69 B 0.040618f
C115 VTAIL.n70 B 0.043296f
C116 VTAIL.n71 B 0.114235f
C117 VTAIL.n72 B 0.022085f
C118 VTAIL.n73 B 0.01623f
C119 VTAIL.n74 B 0.008721f
C120 VTAIL.n75 B 0.020614f
C121 VTAIL.n76 B 0.009234f
C122 VTAIL.n77 B 0.01623f
C123 VTAIL.n78 B 0.008721f
C124 VTAIL.n79 B 0.020614f
C125 VTAIL.n80 B 0.009234f
C126 VTAIL.n81 B 0.01623f
C127 VTAIL.n82 B 0.008721f
C128 VTAIL.n83 B 0.020614f
C129 VTAIL.n84 B 0.009234f
C130 VTAIL.n85 B 0.01623f
C131 VTAIL.n86 B 0.008721f
C132 VTAIL.n87 B 0.020614f
C133 VTAIL.n88 B 0.009234f
C134 VTAIL.n89 B 0.01623f
C135 VTAIL.n90 B 0.008721f
C136 VTAIL.n91 B 0.020614f
C137 VTAIL.n92 B 0.009234f
C138 VTAIL.n93 B 0.932454f
C139 VTAIL.n94 B 0.008721f
C140 VTAIL.t7 B 0.033897f
C141 VTAIL.n95 B 0.099099f
C142 VTAIL.n96 B 0.012177f
C143 VTAIL.n97 B 0.01546f
C144 VTAIL.n98 B 0.020614f
C145 VTAIL.n99 B 0.009234f
C146 VTAIL.n100 B 0.008721f
C147 VTAIL.n101 B 0.01623f
C148 VTAIL.n102 B 0.01623f
C149 VTAIL.n103 B 0.008721f
C150 VTAIL.n104 B 0.009234f
C151 VTAIL.n105 B 0.020614f
C152 VTAIL.n106 B 0.020614f
C153 VTAIL.n107 B 0.009234f
C154 VTAIL.n108 B 0.008721f
C155 VTAIL.n109 B 0.01623f
C156 VTAIL.n110 B 0.01623f
C157 VTAIL.n111 B 0.008721f
C158 VTAIL.n112 B 0.009234f
C159 VTAIL.n113 B 0.020614f
C160 VTAIL.n114 B 0.020614f
C161 VTAIL.n115 B 0.009234f
C162 VTAIL.n116 B 0.008721f
C163 VTAIL.n117 B 0.01623f
C164 VTAIL.n118 B 0.01623f
C165 VTAIL.n119 B 0.008721f
C166 VTAIL.n120 B 0.009234f
C167 VTAIL.n121 B 0.020614f
C168 VTAIL.n122 B 0.020614f
C169 VTAIL.n123 B 0.009234f
C170 VTAIL.n124 B 0.008721f
C171 VTAIL.n125 B 0.01623f
C172 VTAIL.n126 B 0.01623f
C173 VTAIL.n127 B 0.008721f
C174 VTAIL.n128 B 0.009234f
C175 VTAIL.n129 B 0.020614f
C176 VTAIL.n130 B 0.020614f
C177 VTAIL.n131 B 0.009234f
C178 VTAIL.n132 B 0.008721f
C179 VTAIL.n133 B 0.01623f
C180 VTAIL.n134 B 0.01623f
C181 VTAIL.n135 B 0.008721f
C182 VTAIL.n136 B 0.009234f
C183 VTAIL.n137 B 0.020614f
C184 VTAIL.n138 B 0.042081f
C185 VTAIL.n139 B 0.009234f
C186 VTAIL.n140 B 0.017053f
C187 VTAIL.n141 B 0.040618f
C188 VTAIL.n142 B 0.043296f
C189 VTAIL.n143 B 0.182196f
C190 VTAIL.n144 B 0.022085f
C191 VTAIL.n145 B 0.01623f
C192 VTAIL.n146 B 0.008721f
C193 VTAIL.n147 B 0.020614f
C194 VTAIL.n148 B 0.009234f
C195 VTAIL.n149 B 0.01623f
C196 VTAIL.n150 B 0.008721f
C197 VTAIL.n151 B 0.020614f
C198 VTAIL.n152 B 0.009234f
C199 VTAIL.n153 B 0.01623f
C200 VTAIL.n154 B 0.008721f
C201 VTAIL.n155 B 0.020614f
C202 VTAIL.n156 B 0.009234f
C203 VTAIL.n157 B 0.01623f
C204 VTAIL.n158 B 0.008721f
C205 VTAIL.n159 B 0.020614f
C206 VTAIL.n160 B 0.009234f
C207 VTAIL.n161 B 0.01623f
C208 VTAIL.n162 B 0.008721f
C209 VTAIL.n163 B 0.020614f
C210 VTAIL.n164 B 0.009234f
C211 VTAIL.n165 B 0.932454f
C212 VTAIL.n166 B 0.008721f
C213 VTAIL.t0 B 0.033897f
C214 VTAIL.n167 B 0.099099f
C215 VTAIL.n168 B 0.012177f
C216 VTAIL.n169 B 0.01546f
C217 VTAIL.n170 B 0.020614f
C218 VTAIL.n171 B 0.009234f
C219 VTAIL.n172 B 0.008721f
C220 VTAIL.n173 B 0.01623f
C221 VTAIL.n174 B 0.01623f
C222 VTAIL.n175 B 0.008721f
C223 VTAIL.n176 B 0.009234f
C224 VTAIL.n177 B 0.020614f
C225 VTAIL.n178 B 0.020614f
C226 VTAIL.n179 B 0.009234f
C227 VTAIL.n180 B 0.008721f
C228 VTAIL.n181 B 0.01623f
C229 VTAIL.n182 B 0.01623f
C230 VTAIL.n183 B 0.008721f
C231 VTAIL.n184 B 0.009234f
C232 VTAIL.n185 B 0.020614f
C233 VTAIL.n186 B 0.020614f
C234 VTAIL.n187 B 0.009234f
C235 VTAIL.n188 B 0.008721f
C236 VTAIL.n189 B 0.01623f
C237 VTAIL.n190 B 0.01623f
C238 VTAIL.n191 B 0.008721f
C239 VTAIL.n192 B 0.009234f
C240 VTAIL.n193 B 0.020614f
C241 VTAIL.n194 B 0.020614f
C242 VTAIL.n195 B 0.009234f
C243 VTAIL.n196 B 0.008721f
C244 VTAIL.n197 B 0.01623f
C245 VTAIL.n198 B 0.01623f
C246 VTAIL.n199 B 0.008721f
C247 VTAIL.n200 B 0.009234f
C248 VTAIL.n201 B 0.020614f
C249 VTAIL.n202 B 0.020614f
C250 VTAIL.n203 B 0.009234f
C251 VTAIL.n204 B 0.008721f
C252 VTAIL.n205 B 0.01623f
C253 VTAIL.n206 B 0.01623f
C254 VTAIL.n207 B 0.008721f
C255 VTAIL.n208 B 0.009234f
C256 VTAIL.n209 B 0.020614f
C257 VTAIL.n210 B 0.042081f
C258 VTAIL.n211 B 0.009234f
C259 VTAIL.n212 B 0.017053f
C260 VTAIL.n213 B 0.040618f
C261 VTAIL.n214 B 0.043296f
C262 VTAIL.n215 B 1.1215f
C263 VTAIL.n216 B 0.022085f
C264 VTAIL.n217 B 0.01623f
C265 VTAIL.n218 B 0.008721f
C266 VTAIL.n219 B 0.020614f
C267 VTAIL.n220 B 0.009234f
C268 VTAIL.n221 B 0.01623f
C269 VTAIL.n222 B 0.008721f
C270 VTAIL.n223 B 0.020614f
C271 VTAIL.n224 B 0.009234f
C272 VTAIL.n225 B 0.01623f
C273 VTAIL.n226 B 0.008721f
C274 VTAIL.n227 B 0.020614f
C275 VTAIL.n228 B 0.009234f
C276 VTAIL.n229 B 0.01623f
C277 VTAIL.n230 B 0.008721f
C278 VTAIL.n231 B 0.020614f
C279 VTAIL.n232 B 0.009234f
C280 VTAIL.n233 B 0.01623f
C281 VTAIL.n234 B 0.008721f
C282 VTAIL.n235 B 0.020614f
C283 VTAIL.n236 B 0.009234f
C284 VTAIL.n237 B 0.932454f
C285 VTAIL.n238 B 0.008721f
C286 VTAIL.t5 B 0.033897f
C287 VTAIL.n239 B 0.099099f
C288 VTAIL.n240 B 0.012177f
C289 VTAIL.n241 B 0.01546f
C290 VTAIL.n242 B 0.020614f
C291 VTAIL.n243 B 0.009234f
C292 VTAIL.n244 B 0.008721f
C293 VTAIL.n245 B 0.01623f
C294 VTAIL.n246 B 0.01623f
C295 VTAIL.n247 B 0.008721f
C296 VTAIL.n248 B 0.009234f
C297 VTAIL.n249 B 0.020614f
C298 VTAIL.n250 B 0.020614f
C299 VTAIL.n251 B 0.009234f
C300 VTAIL.n252 B 0.008721f
C301 VTAIL.n253 B 0.01623f
C302 VTAIL.n254 B 0.01623f
C303 VTAIL.n255 B 0.008721f
C304 VTAIL.n256 B 0.009234f
C305 VTAIL.n257 B 0.020614f
C306 VTAIL.n258 B 0.020614f
C307 VTAIL.n259 B 0.009234f
C308 VTAIL.n260 B 0.008721f
C309 VTAIL.n261 B 0.01623f
C310 VTAIL.n262 B 0.01623f
C311 VTAIL.n263 B 0.008721f
C312 VTAIL.n264 B 0.009234f
C313 VTAIL.n265 B 0.020614f
C314 VTAIL.n266 B 0.020614f
C315 VTAIL.n267 B 0.009234f
C316 VTAIL.n268 B 0.008721f
C317 VTAIL.n269 B 0.01623f
C318 VTAIL.n270 B 0.01623f
C319 VTAIL.n271 B 0.008721f
C320 VTAIL.n272 B 0.009234f
C321 VTAIL.n273 B 0.020614f
C322 VTAIL.n274 B 0.020614f
C323 VTAIL.n275 B 0.009234f
C324 VTAIL.n276 B 0.008721f
C325 VTAIL.n277 B 0.01623f
C326 VTAIL.n278 B 0.01623f
C327 VTAIL.n279 B 0.008721f
C328 VTAIL.n280 B 0.009234f
C329 VTAIL.n281 B 0.020614f
C330 VTAIL.n282 B 0.042081f
C331 VTAIL.n283 B 0.009234f
C332 VTAIL.n284 B 0.017053f
C333 VTAIL.n285 B 0.040618f
C334 VTAIL.n286 B 0.043296f
C335 VTAIL.n287 B 1.1215f
C336 VTAIL.n288 B 0.022085f
C337 VTAIL.n289 B 0.01623f
C338 VTAIL.n290 B 0.008721f
C339 VTAIL.n291 B 0.020614f
C340 VTAIL.n292 B 0.009234f
C341 VTAIL.n293 B 0.01623f
C342 VTAIL.n294 B 0.008721f
C343 VTAIL.n295 B 0.020614f
C344 VTAIL.n296 B 0.009234f
C345 VTAIL.n297 B 0.01623f
C346 VTAIL.n298 B 0.008721f
C347 VTAIL.n299 B 0.020614f
C348 VTAIL.n300 B 0.009234f
C349 VTAIL.n301 B 0.01623f
C350 VTAIL.n302 B 0.008721f
C351 VTAIL.n303 B 0.020614f
C352 VTAIL.n304 B 0.009234f
C353 VTAIL.n305 B 0.01623f
C354 VTAIL.n306 B 0.008721f
C355 VTAIL.n307 B 0.020614f
C356 VTAIL.n308 B 0.009234f
C357 VTAIL.n309 B 0.932454f
C358 VTAIL.n310 B 0.008721f
C359 VTAIL.t3 B 0.033897f
C360 VTAIL.n311 B 0.099099f
C361 VTAIL.n312 B 0.012177f
C362 VTAIL.n313 B 0.01546f
C363 VTAIL.n314 B 0.020614f
C364 VTAIL.n315 B 0.009234f
C365 VTAIL.n316 B 0.008721f
C366 VTAIL.n317 B 0.01623f
C367 VTAIL.n318 B 0.01623f
C368 VTAIL.n319 B 0.008721f
C369 VTAIL.n320 B 0.009234f
C370 VTAIL.n321 B 0.020614f
C371 VTAIL.n322 B 0.020614f
C372 VTAIL.n323 B 0.009234f
C373 VTAIL.n324 B 0.008721f
C374 VTAIL.n325 B 0.01623f
C375 VTAIL.n326 B 0.01623f
C376 VTAIL.n327 B 0.008721f
C377 VTAIL.n328 B 0.009234f
C378 VTAIL.n329 B 0.020614f
C379 VTAIL.n330 B 0.020614f
C380 VTAIL.n331 B 0.009234f
C381 VTAIL.n332 B 0.008721f
C382 VTAIL.n333 B 0.01623f
C383 VTAIL.n334 B 0.01623f
C384 VTAIL.n335 B 0.008721f
C385 VTAIL.n336 B 0.009234f
C386 VTAIL.n337 B 0.020614f
C387 VTAIL.n338 B 0.020614f
C388 VTAIL.n339 B 0.009234f
C389 VTAIL.n340 B 0.008721f
C390 VTAIL.n341 B 0.01623f
C391 VTAIL.n342 B 0.01623f
C392 VTAIL.n343 B 0.008721f
C393 VTAIL.n344 B 0.009234f
C394 VTAIL.n345 B 0.020614f
C395 VTAIL.n346 B 0.020614f
C396 VTAIL.n347 B 0.009234f
C397 VTAIL.n348 B 0.008721f
C398 VTAIL.n349 B 0.01623f
C399 VTAIL.n350 B 0.01623f
C400 VTAIL.n351 B 0.008721f
C401 VTAIL.n352 B 0.009234f
C402 VTAIL.n353 B 0.020614f
C403 VTAIL.n354 B 0.042081f
C404 VTAIL.n355 B 0.009234f
C405 VTAIL.n356 B 0.017053f
C406 VTAIL.n357 B 0.040618f
C407 VTAIL.n358 B 0.043296f
C408 VTAIL.n359 B 0.182196f
C409 VTAIL.n360 B 0.022085f
C410 VTAIL.n361 B 0.01623f
C411 VTAIL.n362 B 0.008721f
C412 VTAIL.n363 B 0.020614f
C413 VTAIL.n364 B 0.009234f
C414 VTAIL.n365 B 0.01623f
C415 VTAIL.n366 B 0.008721f
C416 VTAIL.n367 B 0.020614f
C417 VTAIL.n368 B 0.009234f
C418 VTAIL.n369 B 0.01623f
C419 VTAIL.n370 B 0.008721f
C420 VTAIL.n371 B 0.020614f
C421 VTAIL.n372 B 0.009234f
C422 VTAIL.n373 B 0.01623f
C423 VTAIL.n374 B 0.008721f
C424 VTAIL.n375 B 0.020614f
C425 VTAIL.n376 B 0.009234f
C426 VTAIL.n377 B 0.01623f
C427 VTAIL.n378 B 0.008721f
C428 VTAIL.n379 B 0.020614f
C429 VTAIL.n380 B 0.009234f
C430 VTAIL.n381 B 0.932454f
C431 VTAIL.n382 B 0.008721f
C432 VTAIL.t6 B 0.033897f
C433 VTAIL.n383 B 0.099099f
C434 VTAIL.n384 B 0.012177f
C435 VTAIL.n385 B 0.01546f
C436 VTAIL.n386 B 0.020614f
C437 VTAIL.n387 B 0.009234f
C438 VTAIL.n388 B 0.008721f
C439 VTAIL.n389 B 0.01623f
C440 VTAIL.n390 B 0.01623f
C441 VTAIL.n391 B 0.008721f
C442 VTAIL.n392 B 0.009234f
C443 VTAIL.n393 B 0.020614f
C444 VTAIL.n394 B 0.020614f
C445 VTAIL.n395 B 0.009234f
C446 VTAIL.n396 B 0.008721f
C447 VTAIL.n397 B 0.01623f
C448 VTAIL.n398 B 0.01623f
C449 VTAIL.n399 B 0.008721f
C450 VTAIL.n400 B 0.009234f
C451 VTAIL.n401 B 0.020614f
C452 VTAIL.n402 B 0.020614f
C453 VTAIL.n403 B 0.009234f
C454 VTAIL.n404 B 0.008721f
C455 VTAIL.n405 B 0.01623f
C456 VTAIL.n406 B 0.01623f
C457 VTAIL.n407 B 0.008721f
C458 VTAIL.n408 B 0.009234f
C459 VTAIL.n409 B 0.020614f
C460 VTAIL.n410 B 0.020614f
C461 VTAIL.n411 B 0.009234f
C462 VTAIL.n412 B 0.008721f
C463 VTAIL.n413 B 0.01623f
C464 VTAIL.n414 B 0.01623f
C465 VTAIL.n415 B 0.008721f
C466 VTAIL.n416 B 0.009234f
C467 VTAIL.n417 B 0.020614f
C468 VTAIL.n418 B 0.020614f
C469 VTAIL.n419 B 0.009234f
C470 VTAIL.n420 B 0.008721f
C471 VTAIL.n421 B 0.01623f
C472 VTAIL.n422 B 0.01623f
C473 VTAIL.n423 B 0.008721f
C474 VTAIL.n424 B 0.009234f
C475 VTAIL.n425 B 0.020614f
C476 VTAIL.n426 B 0.042081f
C477 VTAIL.n427 B 0.009234f
C478 VTAIL.n428 B 0.017053f
C479 VTAIL.n429 B 0.040618f
C480 VTAIL.n430 B 0.043296f
C481 VTAIL.n431 B 0.182196f
C482 VTAIL.n432 B 0.022085f
C483 VTAIL.n433 B 0.01623f
C484 VTAIL.n434 B 0.008721f
C485 VTAIL.n435 B 0.020614f
C486 VTAIL.n436 B 0.009234f
C487 VTAIL.n437 B 0.01623f
C488 VTAIL.n438 B 0.008721f
C489 VTAIL.n439 B 0.020614f
C490 VTAIL.n440 B 0.009234f
C491 VTAIL.n441 B 0.01623f
C492 VTAIL.n442 B 0.008721f
C493 VTAIL.n443 B 0.020614f
C494 VTAIL.n444 B 0.009234f
C495 VTAIL.n445 B 0.01623f
C496 VTAIL.n446 B 0.008721f
C497 VTAIL.n447 B 0.020614f
C498 VTAIL.n448 B 0.009234f
C499 VTAIL.n449 B 0.01623f
C500 VTAIL.n450 B 0.008721f
C501 VTAIL.n451 B 0.020614f
C502 VTAIL.n452 B 0.009234f
C503 VTAIL.n453 B 0.932454f
C504 VTAIL.n454 B 0.008721f
C505 VTAIL.t1 B 0.033897f
C506 VTAIL.n455 B 0.099099f
C507 VTAIL.n456 B 0.012177f
C508 VTAIL.n457 B 0.01546f
C509 VTAIL.n458 B 0.020614f
C510 VTAIL.n459 B 0.009234f
C511 VTAIL.n460 B 0.008721f
C512 VTAIL.n461 B 0.01623f
C513 VTAIL.n462 B 0.01623f
C514 VTAIL.n463 B 0.008721f
C515 VTAIL.n464 B 0.009234f
C516 VTAIL.n465 B 0.020614f
C517 VTAIL.n466 B 0.020614f
C518 VTAIL.n467 B 0.009234f
C519 VTAIL.n468 B 0.008721f
C520 VTAIL.n469 B 0.01623f
C521 VTAIL.n470 B 0.01623f
C522 VTAIL.n471 B 0.008721f
C523 VTAIL.n472 B 0.009234f
C524 VTAIL.n473 B 0.020614f
C525 VTAIL.n474 B 0.020614f
C526 VTAIL.n475 B 0.009234f
C527 VTAIL.n476 B 0.008721f
C528 VTAIL.n477 B 0.01623f
C529 VTAIL.n478 B 0.01623f
C530 VTAIL.n479 B 0.008721f
C531 VTAIL.n480 B 0.009234f
C532 VTAIL.n481 B 0.020614f
C533 VTAIL.n482 B 0.020614f
C534 VTAIL.n483 B 0.009234f
C535 VTAIL.n484 B 0.008721f
C536 VTAIL.n485 B 0.01623f
C537 VTAIL.n486 B 0.01623f
C538 VTAIL.n487 B 0.008721f
C539 VTAIL.n488 B 0.009234f
C540 VTAIL.n489 B 0.020614f
C541 VTAIL.n490 B 0.020614f
C542 VTAIL.n491 B 0.009234f
C543 VTAIL.n492 B 0.008721f
C544 VTAIL.n493 B 0.01623f
C545 VTAIL.n494 B 0.01623f
C546 VTAIL.n495 B 0.008721f
C547 VTAIL.n496 B 0.009234f
C548 VTAIL.n497 B 0.020614f
C549 VTAIL.n498 B 0.042081f
C550 VTAIL.n499 B 0.009234f
C551 VTAIL.n500 B 0.017053f
C552 VTAIL.n501 B 0.040618f
C553 VTAIL.n502 B 0.043296f
C554 VTAIL.n503 B 1.1215f
C555 VTAIL.n504 B 0.022085f
C556 VTAIL.n505 B 0.01623f
C557 VTAIL.n506 B 0.008721f
C558 VTAIL.n507 B 0.020614f
C559 VTAIL.n508 B 0.009234f
C560 VTAIL.n509 B 0.01623f
C561 VTAIL.n510 B 0.008721f
C562 VTAIL.n511 B 0.020614f
C563 VTAIL.n512 B 0.009234f
C564 VTAIL.n513 B 0.01623f
C565 VTAIL.n514 B 0.008721f
C566 VTAIL.n515 B 0.020614f
C567 VTAIL.n516 B 0.009234f
C568 VTAIL.n517 B 0.01623f
C569 VTAIL.n518 B 0.008721f
C570 VTAIL.n519 B 0.020614f
C571 VTAIL.n520 B 0.009234f
C572 VTAIL.n521 B 0.01623f
C573 VTAIL.n522 B 0.008721f
C574 VTAIL.n523 B 0.020614f
C575 VTAIL.n524 B 0.009234f
C576 VTAIL.n525 B 0.932454f
C577 VTAIL.n526 B 0.008721f
C578 VTAIL.t4 B 0.033897f
C579 VTAIL.n527 B 0.099099f
C580 VTAIL.n528 B 0.012177f
C581 VTAIL.n529 B 0.01546f
C582 VTAIL.n530 B 0.020614f
C583 VTAIL.n531 B 0.009234f
C584 VTAIL.n532 B 0.008721f
C585 VTAIL.n533 B 0.01623f
C586 VTAIL.n534 B 0.01623f
C587 VTAIL.n535 B 0.008721f
C588 VTAIL.n536 B 0.009234f
C589 VTAIL.n537 B 0.020614f
C590 VTAIL.n538 B 0.020614f
C591 VTAIL.n539 B 0.009234f
C592 VTAIL.n540 B 0.008721f
C593 VTAIL.n541 B 0.01623f
C594 VTAIL.n542 B 0.01623f
C595 VTAIL.n543 B 0.008721f
C596 VTAIL.n544 B 0.009234f
C597 VTAIL.n545 B 0.020614f
C598 VTAIL.n546 B 0.020614f
C599 VTAIL.n547 B 0.009234f
C600 VTAIL.n548 B 0.008721f
C601 VTAIL.n549 B 0.01623f
C602 VTAIL.n550 B 0.01623f
C603 VTAIL.n551 B 0.008721f
C604 VTAIL.n552 B 0.009234f
C605 VTAIL.n553 B 0.020614f
C606 VTAIL.n554 B 0.020614f
C607 VTAIL.n555 B 0.009234f
C608 VTAIL.n556 B 0.008721f
C609 VTAIL.n557 B 0.01623f
C610 VTAIL.n558 B 0.01623f
C611 VTAIL.n559 B 0.008721f
C612 VTAIL.n560 B 0.009234f
C613 VTAIL.n561 B 0.020614f
C614 VTAIL.n562 B 0.020614f
C615 VTAIL.n563 B 0.009234f
C616 VTAIL.n564 B 0.008721f
C617 VTAIL.n565 B 0.01623f
C618 VTAIL.n566 B 0.01623f
C619 VTAIL.n567 B 0.008721f
C620 VTAIL.n568 B 0.009234f
C621 VTAIL.n569 B 0.020614f
C622 VTAIL.n570 B 0.042081f
C623 VTAIL.n571 B 0.009234f
C624 VTAIL.n572 B 0.017053f
C625 VTAIL.n573 B 0.040618f
C626 VTAIL.n574 B 0.043296f
C627 VTAIL.n575 B 1.04745f
C628 VDD2.t1 B 0.281696f
C629 VDD2.t0 B 0.281696f
C630 VDD2.n0 B 3.24833f
C631 VDD2.t3 B 0.281696f
C632 VDD2.t2 B 0.281696f
C633 VDD2.n1 B 2.53476f
C634 VDD2.n2 B 3.95055f
C635 VN.t3 B 2.68541f
C636 VN.t1 B 2.67948f
C637 VN.n0 B 1.68566f
C638 VN.t2 B 2.68541f
C639 VN.t0 B 2.67948f
C640 VN.n1 B 3.07634f
.ends

