* NGSPICE file created from diff_pair_sample_0375.ext - technology: sky130A

.subckt diff_pair_sample_0375 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t9 VP.t0 VTAIL.t12 B.t5 sky130_fd_pr__nfet_01v8 ad=1.9371 pd=12.07 as=1.9371 ps=12.07 w=11.74 l=2.12
X1 VTAIL.t14 VP.t1 VDD1.t8 B.t9 sky130_fd_pr__nfet_01v8 ad=1.9371 pd=12.07 as=1.9371 ps=12.07 w=11.74 l=2.12
X2 VTAIL.t1 VN.t0 VDD2.t9 B.t1 sky130_fd_pr__nfet_01v8 ad=1.9371 pd=12.07 as=1.9371 ps=12.07 w=11.74 l=2.12
X3 VDD1.t7 VP.t2 VTAIL.t10 B.t7 sky130_fd_pr__nfet_01v8 ad=1.9371 pd=12.07 as=4.5786 ps=24.26 w=11.74 l=2.12
X4 VDD2.t8 VN.t1 VTAIL.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=1.9371 pd=12.07 as=1.9371 ps=12.07 w=11.74 l=2.12
X5 B.t23 B.t21 B.t22 B.t15 sky130_fd_pr__nfet_01v8 ad=4.5786 pd=24.26 as=0 ps=0 w=11.74 l=2.12
X6 B.t20 B.t18 B.t19 B.t11 sky130_fd_pr__nfet_01v8 ad=4.5786 pd=24.26 as=0 ps=0 w=11.74 l=2.12
X7 VTAIL.t0 VN.t2 VDD2.t7 B.t0 sky130_fd_pr__nfet_01v8 ad=1.9371 pd=12.07 as=1.9371 ps=12.07 w=11.74 l=2.12
X8 VTAIL.t9 VP.t3 VDD1.t6 B.t1 sky130_fd_pr__nfet_01v8 ad=1.9371 pd=12.07 as=1.9371 ps=12.07 w=11.74 l=2.12
X9 VDD1.t5 VP.t4 VTAIL.t11 B.t2 sky130_fd_pr__nfet_01v8 ad=4.5786 pd=24.26 as=1.9371 ps=12.07 w=11.74 l=2.12
X10 VDD2.t6 VN.t3 VTAIL.t6 B.t6 sky130_fd_pr__nfet_01v8 ad=4.5786 pd=24.26 as=1.9371 ps=12.07 w=11.74 l=2.12
X11 VDD2.t5 VN.t4 VTAIL.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=1.9371 pd=12.07 as=1.9371 ps=12.07 w=11.74 l=2.12
X12 VTAIL.t15 VP.t5 VDD1.t4 B.t0 sky130_fd_pr__nfet_01v8 ad=1.9371 pd=12.07 as=1.9371 ps=12.07 w=11.74 l=2.12
X13 B.t17 B.t14 B.t16 B.t15 sky130_fd_pr__nfet_01v8 ad=4.5786 pd=24.26 as=0 ps=0 w=11.74 l=2.12
X14 VDD1.t3 VP.t6 VTAIL.t18 B.t6 sky130_fd_pr__nfet_01v8 ad=4.5786 pd=24.26 as=1.9371 ps=12.07 w=11.74 l=2.12
X15 VDD2.t4 VN.t5 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=1.9371 pd=12.07 as=4.5786 ps=24.26 w=11.74 l=2.12
X16 VTAIL.t19 VN.t6 VDD2.t3 B.t9 sky130_fd_pr__nfet_01v8 ad=1.9371 pd=12.07 as=1.9371 ps=12.07 w=11.74 l=2.12
X17 VDD1.t2 VP.t7 VTAIL.t13 B.t3 sky130_fd_pr__nfet_01v8 ad=1.9371 pd=12.07 as=4.5786 ps=24.26 w=11.74 l=2.12
X18 B.t13 B.t10 B.t12 B.t11 sky130_fd_pr__nfet_01v8 ad=4.5786 pd=24.26 as=0 ps=0 w=11.74 l=2.12
X19 VTAIL.t16 VP.t8 VDD1.t1 B.t8 sky130_fd_pr__nfet_01v8 ad=1.9371 pd=12.07 as=1.9371 ps=12.07 w=11.74 l=2.12
X20 VDD1.t0 VP.t9 VTAIL.t17 B.t4 sky130_fd_pr__nfet_01v8 ad=1.9371 pd=12.07 as=1.9371 ps=12.07 w=11.74 l=2.12
X21 VDD2.t2 VN.t7 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=4.5786 pd=24.26 as=1.9371 ps=12.07 w=11.74 l=2.12
X22 VTAIL.t8 VN.t8 VDD2.t1 B.t8 sky130_fd_pr__nfet_01v8 ad=1.9371 pd=12.07 as=1.9371 ps=12.07 w=11.74 l=2.12
X23 VDD2.t0 VN.t9 VTAIL.t7 B.t7 sky130_fd_pr__nfet_01v8 ad=1.9371 pd=12.07 as=4.5786 ps=24.26 w=11.74 l=2.12
R0 VP.n18 VP.t4 167.464
R1 VP.n20 VP.n19 161.3
R2 VP.n21 VP.n16 161.3
R3 VP.n23 VP.n22 161.3
R4 VP.n24 VP.n15 161.3
R5 VP.n26 VP.n25 161.3
R6 VP.n27 VP.n14 161.3
R7 VP.n29 VP.n28 161.3
R8 VP.n30 VP.n13 161.3
R9 VP.n32 VP.n31 161.3
R10 VP.n34 VP.n12 161.3
R11 VP.n36 VP.n35 161.3
R12 VP.n37 VP.n11 161.3
R13 VP.n39 VP.n38 161.3
R14 VP.n40 VP.n10 161.3
R15 VP.n74 VP.n0 161.3
R16 VP.n73 VP.n72 161.3
R17 VP.n71 VP.n1 161.3
R18 VP.n70 VP.n69 161.3
R19 VP.n68 VP.n2 161.3
R20 VP.n66 VP.n65 161.3
R21 VP.n64 VP.n3 161.3
R22 VP.n63 VP.n62 161.3
R23 VP.n61 VP.n4 161.3
R24 VP.n60 VP.n59 161.3
R25 VP.n58 VP.n5 161.3
R26 VP.n57 VP.n56 161.3
R27 VP.n55 VP.n6 161.3
R28 VP.n54 VP.n53 161.3
R29 VP.n52 VP.n51 161.3
R30 VP.n50 VP.n8 161.3
R31 VP.n49 VP.n48 161.3
R32 VP.n47 VP.n9 161.3
R33 VP.n46 VP.n45 161.3
R34 VP.n60 VP.t0 133.459
R35 VP.n44 VP.t6 133.459
R36 VP.n7 VP.t8 133.459
R37 VP.n67 VP.t5 133.459
R38 VP.n75 VP.t7 133.459
R39 VP.n26 VP.t9 133.459
R40 VP.n41 VP.t2 133.459
R41 VP.n33 VP.t3 133.459
R42 VP.n17 VP.t1 133.459
R43 VP.n44 VP.n43 91.1314
R44 VP.n76 VP.n75 91.1314
R45 VP.n42 VP.n41 91.1314
R46 VP.n49 VP.n9 56.4773
R47 VP.n56 VP.n55 56.4773
R48 VP.n62 VP.n3 56.4773
R49 VP.n73 VP.n1 56.4773
R50 VP.n39 VP.n11 56.4773
R51 VP.n28 VP.n13 56.4773
R52 VP.n22 VP.n21 56.4773
R53 VP.n43 VP.n42 50.3594
R54 VP.n18 VP.n17 48.3597
R55 VP.n45 VP.n9 24.3439
R56 VP.n50 VP.n49 24.3439
R57 VP.n51 VP.n50 24.3439
R58 VP.n55 VP.n54 24.3439
R59 VP.n56 VP.n5 24.3439
R60 VP.n60 VP.n5 24.3439
R61 VP.n61 VP.n60 24.3439
R62 VP.n62 VP.n61 24.3439
R63 VP.n66 VP.n3 24.3439
R64 VP.n69 VP.n68 24.3439
R65 VP.n69 VP.n1 24.3439
R66 VP.n74 VP.n73 24.3439
R67 VP.n40 VP.n39 24.3439
R68 VP.n32 VP.n13 24.3439
R69 VP.n35 VP.n34 24.3439
R70 VP.n35 VP.n11 24.3439
R71 VP.n22 VP.n15 24.3439
R72 VP.n26 VP.n15 24.3439
R73 VP.n27 VP.n26 24.3439
R74 VP.n28 VP.n27 24.3439
R75 VP.n21 VP.n20 24.3439
R76 VP.n54 VP.n7 21.9096
R77 VP.n67 VP.n66 21.9096
R78 VP.n33 VP.n32 21.9096
R79 VP.n20 VP.n17 21.9096
R80 VP.n45 VP.n44 19.4752
R81 VP.n75 VP.n74 19.4752
R82 VP.n41 VP.n40 19.4752
R83 VP.n19 VP.n18 9.03227
R84 VP.n51 VP.n7 2.43484
R85 VP.n68 VP.n67 2.43484
R86 VP.n34 VP.n33 2.43484
R87 VP.n42 VP.n10 0.278398
R88 VP.n46 VP.n43 0.278398
R89 VP.n76 VP.n0 0.278398
R90 VP.n19 VP.n16 0.189894
R91 VP.n23 VP.n16 0.189894
R92 VP.n24 VP.n23 0.189894
R93 VP.n25 VP.n24 0.189894
R94 VP.n25 VP.n14 0.189894
R95 VP.n29 VP.n14 0.189894
R96 VP.n30 VP.n29 0.189894
R97 VP.n31 VP.n30 0.189894
R98 VP.n31 VP.n12 0.189894
R99 VP.n36 VP.n12 0.189894
R100 VP.n37 VP.n36 0.189894
R101 VP.n38 VP.n37 0.189894
R102 VP.n38 VP.n10 0.189894
R103 VP.n47 VP.n46 0.189894
R104 VP.n48 VP.n47 0.189894
R105 VP.n48 VP.n8 0.189894
R106 VP.n52 VP.n8 0.189894
R107 VP.n53 VP.n52 0.189894
R108 VP.n53 VP.n6 0.189894
R109 VP.n57 VP.n6 0.189894
R110 VP.n58 VP.n57 0.189894
R111 VP.n59 VP.n58 0.189894
R112 VP.n59 VP.n4 0.189894
R113 VP.n63 VP.n4 0.189894
R114 VP.n64 VP.n63 0.189894
R115 VP.n65 VP.n64 0.189894
R116 VP.n65 VP.n2 0.189894
R117 VP.n70 VP.n2 0.189894
R118 VP.n71 VP.n70 0.189894
R119 VP.n72 VP.n71 0.189894
R120 VP.n72 VP.n0 0.189894
R121 VP VP.n76 0.153422
R122 VTAIL.n11 VTAIL.t3 46.5999
R123 VTAIL.n17 VTAIL.t7 46.5997
R124 VTAIL.n2 VTAIL.t13 46.5997
R125 VTAIL.n16 VTAIL.t10 46.5997
R126 VTAIL.n15 VTAIL.n14 44.9134
R127 VTAIL.n13 VTAIL.n12 44.9134
R128 VTAIL.n10 VTAIL.n9 44.9134
R129 VTAIL.n8 VTAIL.n7 44.9134
R130 VTAIL.n19 VTAIL.n18 44.9131
R131 VTAIL.n1 VTAIL.n0 44.9131
R132 VTAIL.n4 VTAIL.n3 44.9131
R133 VTAIL.n6 VTAIL.n5 44.9131
R134 VTAIL.n8 VTAIL.n6 26.7117
R135 VTAIL.n17 VTAIL.n16 24.5996
R136 VTAIL.n10 VTAIL.n8 2.11257
R137 VTAIL.n11 VTAIL.n10 2.11257
R138 VTAIL.n15 VTAIL.n13 2.11257
R139 VTAIL.n16 VTAIL.n15 2.11257
R140 VTAIL.n6 VTAIL.n4 2.11257
R141 VTAIL.n4 VTAIL.n2 2.11257
R142 VTAIL.n19 VTAIL.n17 2.11257
R143 VTAIL.n18 VTAIL.t4 1.68704
R144 VTAIL.n18 VTAIL.t1 1.68704
R145 VTAIL.n0 VTAIL.t2 1.68704
R146 VTAIL.n0 VTAIL.t19 1.68704
R147 VTAIL.n3 VTAIL.t12 1.68704
R148 VTAIL.n3 VTAIL.t15 1.68704
R149 VTAIL.n5 VTAIL.t18 1.68704
R150 VTAIL.n5 VTAIL.t16 1.68704
R151 VTAIL.n14 VTAIL.t17 1.68704
R152 VTAIL.n14 VTAIL.t9 1.68704
R153 VTAIL.n12 VTAIL.t11 1.68704
R154 VTAIL.n12 VTAIL.t14 1.68704
R155 VTAIL.n9 VTAIL.t5 1.68704
R156 VTAIL.n9 VTAIL.t0 1.68704
R157 VTAIL.n7 VTAIL.t6 1.68704
R158 VTAIL.n7 VTAIL.t8 1.68704
R159 VTAIL VTAIL.n1 1.64274
R160 VTAIL.n13 VTAIL.n11 1.52636
R161 VTAIL.n2 VTAIL.n1 1.52636
R162 VTAIL VTAIL.n19 0.470328
R163 VDD1.n1 VDD1.t5 65.3908
R164 VDD1.n3 VDD1.t3 65.3905
R165 VDD1.n5 VDD1.n4 63.1206
R166 VDD1.n1 VDD1.n0 61.5921
R167 VDD1.n7 VDD1.n6 61.592
R168 VDD1.n3 VDD1.n2 61.5919
R169 VDD1.n7 VDD1.n5 45.5074
R170 VDD1.n6 VDD1.t6 1.68704
R171 VDD1.n6 VDD1.t7 1.68704
R172 VDD1.n0 VDD1.t8 1.68704
R173 VDD1.n0 VDD1.t0 1.68704
R174 VDD1.n4 VDD1.t4 1.68704
R175 VDD1.n4 VDD1.t2 1.68704
R176 VDD1.n2 VDD1.t1 1.68704
R177 VDD1.n2 VDD1.t9 1.68704
R178 VDD1 VDD1.n7 1.52636
R179 VDD1 VDD1.n1 0.586707
R180 VDD1.n5 VDD1.n3 0.473171
R181 B.n877 B.n876 585
R182 B.n878 B.n877 585
R183 B.n323 B.n141 585
R184 B.n322 B.n321 585
R185 B.n320 B.n319 585
R186 B.n318 B.n317 585
R187 B.n316 B.n315 585
R188 B.n314 B.n313 585
R189 B.n312 B.n311 585
R190 B.n310 B.n309 585
R191 B.n308 B.n307 585
R192 B.n306 B.n305 585
R193 B.n304 B.n303 585
R194 B.n302 B.n301 585
R195 B.n300 B.n299 585
R196 B.n298 B.n297 585
R197 B.n296 B.n295 585
R198 B.n294 B.n293 585
R199 B.n292 B.n291 585
R200 B.n290 B.n289 585
R201 B.n288 B.n287 585
R202 B.n286 B.n285 585
R203 B.n284 B.n283 585
R204 B.n282 B.n281 585
R205 B.n280 B.n279 585
R206 B.n278 B.n277 585
R207 B.n276 B.n275 585
R208 B.n274 B.n273 585
R209 B.n272 B.n271 585
R210 B.n270 B.n269 585
R211 B.n268 B.n267 585
R212 B.n266 B.n265 585
R213 B.n264 B.n263 585
R214 B.n262 B.n261 585
R215 B.n260 B.n259 585
R216 B.n258 B.n257 585
R217 B.n256 B.n255 585
R218 B.n254 B.n253 585
R219 B.n252 B.n251 585
R220 B.n250 B.n249 585
R221 B.n248 B.n247 585
R222 B.n246 B.n245 585
R223 B.n244 B.n243 585
R224 B.n242 B.n241 585
R225 B.n240 B.n239 585
R226 B.n238 B.n237 585
R227 B.n236 B.n235 585
R228 B.n234 B.n233 585
R229 B.n232 B.n231 585
R230 B.n230 B.n229 585
R231 B.n228 B.n227 585
R232 B.n225 B.n224 585
R233 B.n223 B.n222 585
R234 B.n221 B.n220 585
R235 B.n219 B.n218 585
R236 B.n217 B.n216 585
R237 B.n215 B.n214 585
R238 B.n213 B.n212 585
R239 B.n211 B.n210 585
R240 B.n209 B.n208 585
R241 B.n207 B.n206 585
R242 B.n205 B.n204 585
R243 B.n203 B.n202 585
R244 B.n201 B.n200 585
R245 B.n199 B.n198 585
R246 B.n197 B.n196 585
R247 B.n195 B.n194 585
R248 B.n193 B.n192 585
R249 B.n191 B.n190 585
R250 B.n189 B.n188 585
R251 B.n187 B.n186 585
R252 B.n185 B.n184 585
R253 B.n183 B.n182 585
R254 B.n181 B.n180 585
R255 B.n179 B.n178 585
R256 B.n177 B.n176 585
R257 B.n175 B.n174 585
R258 B.n173 B.n172 585
R259 B.n171 B.n170 585
R260 B.n169 B.n168 585
R261 B.n167 B.n166 585
R262 B.n165 B.n164 585
R263 B.n163 B.n162 585
R264 B.n161 B.n160 585
R265 B.n159 B.n158 585
R266 B.n157 B.n156 585
R267 B.n155 B.n154 585
R268 B.n153 B.n152 585
R269 B.n151 B.n150 585
R270 B.n149 B.n148 585
R271 B.n96 B.n95 585
R272 B.n881 B.n880 585
R273 B.n875 B.n142 585
R274 B.n142 B.n93 585
R275 B.n874 B.n92 585
R276 B.n885 B.n92 585
R277 B.n873 B.n91 585
R278 B.n886 B.n91 585
R279 B.n872 B.n90 585
R280 B.n887 B.n90 585
R281 B.n871 B.n870 585
R282 B.n870 B.n86 585
R283 B.n869 B.n85 585
R284 B.n893 B.n85 585
R285 B.n868 B.n84 585
R286 B.n894 B.n84 585
R287 B.n867 B.n83 585
R288 B.n895 B.n83 585
R289 B.n866 B.n865 585
R290 B.n865 B.n79 585
R291 B.n864 B.n78 585
R292 B.n901 B.n78 585
R293 B.n863 B.n77 585
R294 B.n902 B.n77 585
R295 B.n862 B.n76 585
R296 B.n903 B.n76 585
R297 B.n861 B.n860 585
R298 B.n860 B.n72 585
R299 B.n859 B.n71 585
R300 B.n909 B.n71 585
R301 B.n858 B.n70 585
R302 B.n910 B.n70 585
R303 B.n857 B.n69 585
R304 B.n911 B.n69 585
R305 B.n856 B.n855 585
R306 B.n855 B.n65 585
R307 B.n854 B.n64 585
R308 B.n917 B.n64 585
R309 B.n853 B.n63 585
R310 B.n918 B.n63 585
R311 B.n852 B.n62 585
R312 B.n919 B.n62 585
R313 B.n851 B.n850 585
R314 B.n850 B.n58 585
R315 B.n849 B.n57 585
R316 B.n925 B.n57 585
R317 B.n848 B.n56 585
R318 B.n926 B.n56 585
R319 B.n847 B.n55 585
R320 B.n927 B.n55 585
R321 B.n846 B.n845 585
R322 B.n845 B.n54 585
R323 B.n844 B.n50 585
R324 B.n933 B.n50 585
R325 B.n843 B.n49 585
R326 B.n934 B.n49 585
R327 B.n842 B.n48 585
R328 B.n935 B.n48 585
R329 B.n841 B.n840 585
R330 B.n840 B.n44 585
R331 B.n839 B.n43 585
R332 B.n941 B.n43 585
R333 B.n838 B.n42 585
R334 B.n942 B.n42 585
R335 B.n837 B.n41 585
R336 B.n943 B.n41 585
R337 B.n836 B.n835 585
R338 B.n835 B.n37 585
R339 B.n834 B.n36 585
R340 B.n949 B.n36 585
R341 B.n833 B.n35 585
R342 B.n950 B.n35 585
R343 B.n832 B.n34 585
R344 B.n951 B.n34 585
R345 B.n831 B.n830 585
R346 B.n830 B.n30 585
R347 B.n829 B.n29 585
R348 B.n957 B.n29 585
R349 B.n828 B.n28 585
R350 B.n958 B.n28 585
R351 B.n827 B.n27 585
R352 B.n959 B.n27 585
R353 B.n826 B.n825 585
R354 B.n825 B.n23 585
R355 B.n824 B.n22 585
R356 B.n965 B.n22 585
R357 B.n823 B.n21 585
R358 B.n966 B.n21 585
R359 B.n822 B.n20 585
R360 B.n967 B.n20 585
R361 B.n821 B.n820 585
R362 B.n820 B.n16 585
R363 B.n819 B.n15 585
R364 B.n973 B.n15 585
R365 B.n818 B.n14 585
R366 B.n974 B.n14 585
R367 B.n817 B.n13 585
R368 B.n975 B.n13 585
R369 B.n816 B.n815 585
R370 B.n815 B.n12 585
R371 B.n814 B.n813 585
R372 B.n814 B.n8 585
R373 B.n812 B.n7 585
R374 B.n982 B.n7 585
R375 B.n811 B.n6 585
R376 B.n983 B.n6 585
R377 B.n810 B.n5 585
R378 B.n984 B.n5 585
R379 B.n809 B.n808 585
R380 B.n808 B.n4 585
R381 B.n807 B.n324 585
R382 B.n807 B.n806 585
R383 B.n797 B.n325 585
R384 B.n326 B.n325 585
R385 B.n799 B.n798 585
R386 B.n800 B.n799 585
R387 B.n796 B.n330 585
R388 B.n334 B.n330 585
R389 B.n795 B.n794 585
R390 B.n794 B.n793 585
R391 B.n332 B.n331 585
R392 B.n333 B.n332 585
R393 B.n786 B.n785 585
R394 B.n787 B.n786 585
R395 B.n784 B.n339 585
R396 B.n339 B.n338 585
R397 B.n783 B.n782 585
R398 B.n782 B.n781 585
R399 B.n341 B.n340 585
R400 B.n342 B.n341 585
R401 B.n774 B.n773 585
R402 B.n775 B.n774 585
R403 B.n772 B.n347 585
R404 B.n347 B.n346 585
R405 B.n771 B.n770 585
R406 B.n770 B.n769 585
R407 B.n349 B.n348 585
R408 B.n350 B.n349 585
R409 B.n762 B.n761 585
R410 B.n763 B.n762 585
R411 B.n760 B.n355 585
R412 B.n355 B.n354 585
R413 B.n759 B.n758 585
R414 B.n758 B.n757 585
R415 B.n357 B.n356 585
R416 B.n358 B.n357 585
R417 B.n750 B.n749 585
R418 B.n751 B.n750 585
R419 B.n748 B.n363 585
R420 B.n363 B.n362 585
R421 B.n747 B.n746 585
R422 B.n746 B.n745 585
R423 B.n365 B.n364 585
R424 B.n366 B.n365 585
R425 B.n738 B.n737 585
R426 B.n739 B.n738 585
R427 B.n736 B.n371 585
R428 B.n371 B.n370 585
R429 B.n735 B.n734 585
R430 B.n734 B.n733 585
R431 B.n373 B.n372 585
R432 B.n726 B.n373 585
R433 B.n725 B.n724 585
R434 B.n727 B.n725 585
R435 B.n723 B.n378 585
R436 B.n378 B.n377 585
R437 B.n722 B.n721 585
R438 B.n721 B.n720 585
R439 B.n380 B.n379 585
R440 B.n381 B.n380 585
R441 B.n713 B.n712 585
R442 B.n714 B.n713 585
R443 B.n711 B.n386 585
R444 B.n386 B.n385 585
R445 B.n710 B.n709 585
R446 B.n709 B.n708 585
R447 B.n388 B.n387 585
R448 B.n389 B.n388 585
R449 B.n701 B.n700 585
R450 B.n702 B.n701 585
R451 B.n699 B.n394 585
R452 B.n394 B.n393 585
R453 B.n698 B.n697 585
R454 B.n697 B.n696 585
R455 B.n396 B.n395 585
R456 B.n397 B.n396 585
R457 B.n689 B.n688 585
R458 B.n690 B.n689 585
R459 B.n687 B.n402 585
R460 B.n402 B.n401 585
R461 B.n686 B.n685 585
R462 B.n685 B.n684 585
R463 B.n404 B.n403 585
R464 B.n405 B.n404 585
R465 B.n677 B.n676 585
R466 B.n678 B.n677 585
R467 B.n675 B.n410 585
R468 B.n410 B.n409 585
R469 B.n674 B.n673 585
R470 B.n673 B.n672 585
R471 B.n412 B.n411 585
R472 B.n413 B.n412 585
R473 B.n665 B.n664 585
R474 B.n666 B.n665 585
R475 B.n663 B.n418 585
R476 B.n418 B.n417 585
R477 B.n662 B.n661 585
R478 B.n661 B.n660 585
R479 B.n420 B.n419 585
R480 B.n421 B.n420 585
R481 B.n656 B.n655 585
R482 B.n424 B.n423 585
R483 B.n652 B.n651 585
R484 B.n653 B.n652 585
R485 B.n650 B.n469 585
R486 B.n649 B.n648 585
R487 B.n647 B.n646 585
R488 B.n645 B.n644 585
R489 B.n643 B.n642 585
R490 B.n641 B.n640 585
R491 B.n639 B.n638 585
R492 B.n637 B.n636 585
R493 B.n635 B.n634 585
R494 B.n633 B.n632 585
R495 B.n631 B.n630 585
R496 B.n629 B.n628 585
R497 B.n627 B.n626 585
R498 B.n625 B.n624 585
R499 B.n623 B.n622 585
R500 B.n621 B.n620 585
R501 B.n619 B.n618 585
R502 B.n617 B.n616 585
R503 B.n615 B.n614 585
R504 B.n613 B.n612 585
R505 B.n611 B.n610 585
R506 B.n609 B.n608 585
R507 B.n607 B.n606 585
R508 B.n605 B.n604 585
R509 B.n603 B.n602 585
R510 B.n601 B.n600 585
R511 B.n599 B.n598 585
R512 B.n597 B.n596 585
R513 B.n595 B.n594 585
R514 B.n593 B.n592 585
R515 B.n591 B.n590 585
R516 B.n589 B.n588 585
R517 B.n587 B.n586 585
R518 B.n585 B.n584 585
R519 B.n583 B.n582 585
R520 B.n581 B.n580 585
R521 B.n579 B.n578 585
R522 B.n577 B.n576 585
R523 B.n575 B.n574 585
R524 B.n573 B.n572 585
R525 B.n571 B.n570 585
R526 B.n569 B.n568 585
R527 B.n567 B.n566 585
R528 B.n565 B.n564 585
R529 B.n563 B.n562 585
R530 B.n561 B.n560 585
R531 B.n559 B.n558 585
R532 B.n556 B.n555 585
R533 B.n554 B.n553 585
R534 B.n552 B.n551 585
R535 B.n550 B.n549 585
R536 B.n548 B.n547 585
R537 B.n546 B.n545 585
R538 B.n544 B.n543 585
R539 B.n542 B.n541 585
R540 B.n540 B.n539 585
R541 B.n538 B.n537 585
R542 B.n536 B.n535 585
R543 B.n534 B.n533 585
R544 B.n532 B.n531 585
R545 B.n530 B.n529 585
R546 B.n528 B.n527 585
R547 B.n526 B.n525 585
R548 B.n524 B.n523 585
R549 B.n522 B.n521 585
R550 B.n520 B.n519 585
R551 B.n518 B.n517 585
R552 B.n516 B.n515 585
R553 B.n514 B.n513 585
R554 B.n512 B.n511 585
R555 B.n510 B.n509 585
R556 B.n508 B.n507 585
R557 B.n506 B.n505 585
R558 B.n504 B.n503 585
R559 B.n502 B.n501 585
R560 B.n500 B.n499 585
R561 B.n498 B.n497 585
R562 B.n496 B.n495 585
R563 B.n494 B.n493 585
R564 B.n492 B.n491 585
R565 B.n490 B.n489 585
R566 B.n488 B.n487 585
R567 B.n486 B.n485 585
R568 B.n484 B.n483 585
R569 B.n482 B.n481 585
R570 B.n480 B.n479 585
R571 B.n478 B.n477 585
R572 B.n476 B.n475 585
R573 B.n657 B.n422 585
R574 B.n422 B.n421 585
R575 B.n659 B.n658 585
R576 B.n660 B.n659 585
R577 B.n416 B.n415 585
R578 B.n417 B.n416 585
R579 B.n668 B.n667 585
R580 B.n667 B.n666 585
R581 B.n669 B.n414 585
R582 B.n414 B.n413 585
R583 B.n671 B.n670 585
R584 B.n672 B.n671 585
R585 B.n408 B.n407 585
R586 B.n409 B.n408 585
R587 B.n680 B.n679 585
R588 B.n679 B.n678 585
R589 B.n681 B.n406 585
R590 B.n406 B.n405 585
R591 B.n683 B.n682 585
R592 B.n684 B.n683 585
R593 B.n400 B.n399 585
R594 B.n401 B.n400 585
R595 B.n692 B.n691 585
R596 B.n691 B.n690 585
R597 B.n693 B.n398 585
R598 B.n398 B.n397 585
R599 B.n695 B.n694 585
R600 B.n696 B.n695 585
R601 B.n392 B.n391 585
R602 B.n393 B.n392 585
R603 B.n704 B.n703 585
R604 B.n703 B.n702 585
R605 B.n705 B.n390 585
R606 B.n390 B.n389 585
R607 B.n707 B.n706 585
R608 B.n708 B.n707 585
R609 B.n384 B.n383 585
R610 B.n385 B.n384 585
R611 B.n716 B.n715 585
R612 B.n715 B.n714 585
R613 B.n717 B.n382 585
R614 B.n382 B.n381 585
R615 B.n719 B.n718 585
R616 B.n720 B.n719 585
R617 B.n376 B.n375 585
R618 B.n377 B.n376 585
R619 B.n729 B.n728 585
R620 B.n728 B.n727 585
R621 B.n730 B.n374 585
R622 B.n726 B.n374 585
R623 B.n732 B.n731 585
R624 B.n733 B.n732 585
R625 B.n369 B.n368 585
R626 B.n370 B.n369 585
R627 B.n741 B.n740 585
R628 B.n740 B.n739 585
R629 B.n742 B.n367 585
R630 B.n367 B.n366 585
R631 B.n744 B.n743 585
R632 B.n745 B.n744 585
R633 B.n361 B.n360 585
R634 B.n362 B.n361 585
R635 B.n753 B.n752 585
R636 B.n752 B.n751 585
R637 B.n754 B.n359 585
R638 B.n359 B.n358 585
R639 B.n756 B.n755 585
R640 B.n757 B.n756 585
R641 B.n353 B.n352 585
R642 B.n354 B.n353 585
R643 B.n765 B.n764 585
R644 B.n764 B.n763 585
R645 B.n766 B.n351 585
R646 B.n351 B.n350 585
R647 B.n768 B.n767 585
R648 B.n769 B.n768 585
R649 B.n345 B.n344 585
R650 B.n346 B.n345 585
R651 B.n777 B.n776 585
R652 B.n776 B.n775 585
R653 B.n778 B.n343 585
R654 B.n343 B.n342 585
R655 B.n780 B.n779 585
R656 B.n781 B.n780 585
R657 B.n337 B.n336 585
R658 B.n338 B.n337 585
R659 B.n789 B.n788 585
R660 B.n788 B.n787 585
R661 B.n790 B.n335 585
R662 B.n335 B.n333 585
R663 B.n792 B.n791 585
R664 B.n793 B.n792 585
R665 B.n329 B.n328 585
R666 B.n334 B.n329 585
R667 B.n802 B.n801 585
R668 B.n801 B.n800 585
R669 B.n803 B.n327 585
R670 B.n327 B.n326 585
R671 B.n805 B.n804 585
R672 B.n806 B.n805 585
R673 B.n3 B.n0 585
R674 B.n4 B.n3 585
R675 B.n981 B.n1 585
R676 B.n982 B.n981 585
R677 B.n980 B.n979 585
R678 B.n980 B.n8 585
R679 B.n978 B.n9 585
R680 B.n12 B.n9 585
R681 B.n977 B.n976 585
R682 B.n976 B.n975 585
R683 B.n11 B.n10 585
R684 B.n974 B.n11 585
R685 B.n972 B.n971 585
R686 B.n973 B.n972 585
R687 B.n970 B.n17 585
R688 B.n17 B.n16 585
R689 B.n969 B.n968 585
R690 B.n968 B.n967 585
R691 B.n19 B.n18 585
R692 B.n966 B.n19 585
R693 B.n964 B.n963 585
R694 B.n965 B.n964 585
R695 B.n962 B.n24 585
R696 B.n24 B.n23 585
R697 B.n961 B.n960 585
R698 B.n960 B.n959 585
R699 B.n26 B.n25 585
R700 B.n958 B.n26 585
R701 B.n956 B.n955 585
R702 B.n957 B.n956 585
R703 B.n954 B.n31 585
R704 B.n31 B.n30 585
R705 B.n953 B.n952 585
R706 B.n952 B.n951 585
R707 B.n33 B.n32 585
R708 B.n950 B.n33 585
R709 B.n948 B.n947 585
R710 B.n949 B.n948 585
R711 B.n946 B.n38 585
R712 B.n38 B.n37 585
R713 B.n945 B.n944 585
R714 B.n944 B.n943 585
R715 B.n40 B.n39 585
R716 B.n942 B.n40 585
R717 B.n940 B.n939 585
R718 B.n941 B.n940 585
R719 B.n938 B.n45 585
R720 B.n45 B.n44 585
R721 B.n937 B.n936 585
R722 B.n936 B.n935 585
R723 B.n47 B.n46 585
R724 B.n934 B.n47 585
R725 B.n932 B.n931 585
R726 B.n933 B.n932 585
R727 B.n930 B.n51 585
R728 B.n54 B.n51 585
R729 B.n929 B.n928 585
R730 B.n928 B.n927 585
R731 B.n53 B.n52 585
R732 B.n926 B.n53 585
R733 B.n924 B.n923 585
R734 B.n925 B.n924 585
R735 B.n922 B.n59 585
R736 B.n59 B.n58 585
R737 B.n921 B.n920 585
R738 B.n920 B.n919 585
R739 B.n61 B.n60 585
R740 B.n918 B.n61 585
R741 B.n916 B.n915 585
R742 B.n917 B.n916 585
R743 B.n914 B.n66 585
R744 B.n66 B.n65 585
R745 B.n913 B.n912 585
R746 B.n912 B.n911 585
R747 B.n68 B.n67 585
R748 B.n910 B.n68 585
R749 B.n908 B.n907 585
R750 B.n909 B.n908 585
R751 B.n906 B.n73 585
R752 B.n73 B.n72 585
R753 B.n905 B.n904 585
R754 B.n904 B.n903 585
R755 B.n75 B.n74 585
R756 B.n902 B.n75 585
R757 B.n900 B.n899 585
R758 B.n901 B.n900 585
R759 B.n898 B.n80 585
R760 B.n80 B.n79 585
R761 B.n897 B.n896 585
R762 B.n896 B.n895 585
R763 B.n82 B.n81 585
R764 B.n894 B.n82 585
R765 B.n892 B.n891 585
R766 B.n893 B.n892 585
R767 B.n890 B.n87 585
R768 B.n87 B.n86 585
R769 B.n889 B.n888 585
R770 B.n888 B.n887 585
R771 B.n89 B.n88 585
R772 B.n886 B.n89 585
R773 B.n884 B.n883 585
R774 B.n885 B.n884 585
R775 B.n882 B.n94 585
R776 B.n94 B.n93 585
R777 B.n985 B.n984 585
R778 B.n983 B.n2 585
R779 B.n880 B.n94 497.305
R780 B.n877 B.n142 497.305
R781 B.n475 B.n420 497.305
R782 B.n655 B.n422 497.305
R783 B.n146 B.t21 340.646
R784 B.n143 B.t14 340.646
R785 B.n473 B.t18 340.646
R786 B.n470 B.t10 340.646
R787 B.n878 B.n140 256.663
R788 B.n878 B.n139 256.663
R789 B.n878 B.n138 256.663
R790 B.n878 B.n137 256.663
R791 B.n878 B.n136 256.663
R792 B.n878 B.n135 256.663
R793 B.n878 B.n134 256.663
R794 B.n878 B.n133 256.663
R795 B.n878 B.n132 256.663
R796 B.n878 B.n131 256.663
R797 B.n878 B.n130 256.663
R798 B.n878 B.n129 256.663
R799 B.n878 B.n128 256.663
R800 B.n878 B.n127 256.663
R801 B.n878 B.n126 256.663
R802 B.n878 B.n125 256.663
R803 B.n878 B.n124 256.663
R804 B.n878 B.n123 256.663
R805 B.n878 B.n122 256.663
R806 B.n878 B.n121 256.663
R807 B.n878 B.n120 256.663
R808 B.n878 B.n119 256.663
R809 B.n878 B.n118 256.663
R810 B.n878 B.n117 256.663
R811 B.n878 B.n116 256.663
R812 B.n878 B.n115 256.663
R813 B.n878 B.n114 256.663
R814 B.n878 B.n113 256.663
R815 B.n878 B.n112 256.663
R816 B.n878 B.n111 256.663
R817 B.n878 B.n110 256.663
R818 B.n878 B.n109 256.663
R819 B.n878 B.n108 256.663
R820 B.n878 B.n107 256.663
R821 B.n878 B.n106 256.663
R822 B.n878 B.n105 256.663
R823 B.n878 B.n104 256.663
R824 B.n878 B.n103 256.663
R825 B.n878 B.n102 256.663
R826 B.n878 B.n101 256.663
R827 B.n878 B.n100 256.663
R828 B.n878 B.n99 256.663
R829 B.n878 B.n98 256.663
R830 B.n878 B.n97 256.663
R831 B.n879 B.n878 256.663
R832 B.n654 B.n653 256.663
R833 B.n653 B.n425 256.663
R834 B.n653 B.n426 256.663
R835 B.n653 B.n427 256.663
R836 B.n653 B.n428 256.663
R837 B.n653 B.n429 256.663
R838 B.n653 B.n430 256.663
R839 B.n653 B.n431 256.663
R840 B.n653 B.n432 256.663
R841 B.n653 B.n433 256.663
R842 B.n653 B.n434 256.663
R843 B.n653 B.n435 256.663
R844 B.n653 B.n436 256.663
R845 B.n653 B.n437 256.663
R846 B.n653 B.n438 256.663
R847 B.n653 B.n439 256.663
R848 B.n653 B.n440 256.663
R849 B.n653 B.n441 256.663
R850 B.n653 B.n442 256.663
R851 B.n653 B.n443 256.663
R852 B.n653 B.n444 256.663
R853 B.n653 B.n445 256.663
R854 B.n653 B.n446 256.663
R855 B.n653 B.n447 256.663
R856 B.n653 B.n448 256.663
R857 B.n653 B.n449 256.663
R858 B.n653 B.n450 256.663
R859 B.n653 B.n451 256.663
R860 B.n653 B.n452 256.663
R861 B.n653 B.n453 256.663
R862 B.n653 B.n454 256.663
R863 B.n653 B.n455 256.663
R864 B.n653 B.n456 256.663
R865 B.n653 B.n457 256.663
R866 B.n653 B.n458 256.663
R867 B.n653 B.n459 256.663
R868 B.n653 B.n460 256.663
R869 B.n653 B.n461 256.663
R870 B.n653 B.n462 256.663
R871 B.n653 B.n463 256.663
R872 B.n653 B.n464 256.663
R873 B.n653 B.n465 256.663
R874 B.n653 B.n466 256.663
R875 B.n653 B.n467 256.663
R876 B.n653 B.n468 256.663
R877 B.n987 B.n986 256.663
R878 B.n148 B.n96 163.367
R879 B.n152 B.n151 163.367
R880 B.n156 B.n155 163.367
R881 B.n160 B.n159 163.367
R882 B.n164 B.n163 163.367
R883 B.n168 B.n167 163.367
R884 B.n172 B.n171 163.367
R885 B.n176 B.n175 163.367
R886 B.n180 B.n179 163.367
R887 B.n184 B.n183 163.367
R888 B.n188 B.n187 163.367
R889 B.n192 B.n191 163.367
R890 B.n196 B.n195 163.367
R891 B.n200 B.n199 163.367
R892 B.n204 B.n203 163.367
R893 B.n208 B.n207 163.367
R894 B.n212 B.n211 163.367
R895 B.n216 B.n215 163.367
R896 B.n220 B.n219 163.367
R897 B.n224 B.n223 163.367
R898 B.n229 B.n228 163.367
R899 B.n233 B.n232 163.367
R900 B.n237 B.n236 163.367
R901 B.n241 B.n240 163.367
R902 B.n245 B.n244 163.367
R903 B.n249 B.n248 163.367
R904 B.n253 B.n252 163.367
R905 B.n257 B.n256 163.367
R906 B.n261 B.n260 163.367
R907 B.n265 B.n264 163.367
R908 B.n269 B.n268 163.367
R909 B.n273 B.n272 163.367
R910 B.n277 B.n276 163.367
R911 B.n281 B.n280 163.367
R912 B.n285 B.n284 163.367
R913 B.n289 B.n288 163.367
R914 B.n293 B.n292 163.367
R915 B.n297 B.n296 163.367
R916 B.n301 B.n300 163.367
R917 B.n305 B.n304 163.367
R918 B.n309 B.n308 163.367
R919 B.n313 B.n312 163.367
R920 B.n317 B.n316 163.367
R921 B.n321 B.n320 163.367
R922 B.n877 B.n141 163.367
R923 B.n661 B.n420 163.367
R924 B.n661 B.n418 163.367
R925 B.n665 B.n418 163.367
R926 B.n665 B.n412 163.367
R927 B.n673 B.n412 163.367
R928 B.n673 B.n410 163.367
R929 B.n677 B.n410 163.367
R930 B.n677 B.n404 163.367
R931 B.n685 B.n404 163.367
R932 B.n685 B.n402 163.367
R933 B.n689 B.n402 163.367
R934 B.n689 B.n396 163.367
R935 B.n697 B.n396 163.367
R936 B.n697 B.n394 163.367
R937 B.n701 B.n394 163.367
R938 B.n701 B.n388 163.367
R939 B.n709 B.n388 163.367
R940 B.n709 B.n386 163.367
R941 B.n713 B.n386 163.367
R942 B.n713 B.n380 163.367
R943 B.n721 B.n380 163.367
R944 B.n721 B.n378 163.367
R945 B.n725 B.n378 163.367
R946 B.n725 B.n373 163.367
R947 B.n734 B.n373 163.367
R948 B.n734 B.n371 163.367
R949 B.n738 B.n371 163.367
R950 B.n738 B.n365 163.367
R951 B.n746 B.n365 163.367
R952 B.n746 B.n363 163.367
R953 B.n750 B.n363 163.367
R954 B.n750 B.n357 163.367
R955 B.n758 B.n357 163.367
R956 B.n758 B.n355 163.367
R957 B.n762 B.n355 163.367
R958 B.n762 B.n349 163.367
R959 B.n770 B.n349 163.367
R960 B.n770 B.n347 163.367
R961 B.n774 B.n347 163.367
R962 B.n774 B.n341 163.367
R963 B.n782 B.n341 163.367
R964 B.n782 B.n339 163.367
R965 B.n786 B.n339 163.367
R966 B.n786 B.n332 163.367
R967 B.n794 B.n332 163.367
R968 B.n794 B.n330 163.367
R969 B.n799 B.n330 163.367
R970 B.n799 B.n325 163.367
R971 B.n807 B.n325 163.367
R972 B.n808 B.n807 163.367
R973 B.n808 B.n5 163.367
R974 B.n6 B.n5 163.367
R975 B.n7 B.n6 163.367
R976 B.n814 B.n7 163.367
R977 B.n815 B.n814 163.367
R978 B.n815 B.n13 163.367
R979 B.n14 B.n13 163.367
R980 B.n15 B.n14 163.367
R981 B.n820 B.n15 163.367
R982 B.n820 B.n20 163.367
R983 B.n21 B.n20 163.367
R984 B.n22 B.n21 163.367
R985 B.n825 B.n22 163.367
R986 B.n825 B.n27 163.367
R987 B.n28 B.n27 163.367
R988 B.n29 B.n28 163.367
R989 B.n830 B.n29 163.367
R990 B.n830 B.n34 163.367
R991 B.n35 B.n34 163.367
R992 B.n36 B.n35 163.367
R993 B.n835 B.n36 163.367
R994 B.n835 B.n41 163.367
R995 B.n42 B.n41 163.367
R996 B.n43 B.n42 163.367
R997 B.n840 B.n43 163.367
R998 B.n840 B.n48 163.367
R999 B.n49 B.n48 163.367
R1000 B.n50 B.n49 163.367
R1001 B.n845 B.n50 163.367
R1002 B.n845 B.n55 163.367
R1003 B.n56 B.n55 163.367
R1004 B.n57 B.n56 163.367
R1005 B.n850 B.n57 163.367
R1006 B.n850 B.n62 163.367
R1007 B.n63 B.n62 163.367
R1008 B.n64 B.n63 163.367
R1009 B.n855 B.n64 163.367
R1010 B.n855 B.n69 163.367
R1011 B.n70 B.n69 163.367
R1012 B.n71 B.n70 163.367
R1013 B.n860 B.n71 163.367
R1014 B.n860 B.n76 163.367
R1015 B.n77 B.n76 163.367
R1016 B.n78 B.n77 163.367
R1017 B.n865 B.n78 163.367
R1018 B.n865 B.n83 163.367
R1019 B.n84 B.n83 163.367
R1020 B.n85 B.n84 163.367
R1021 B.n870 B.n85 163.367
R1022 B.n870 B.n90 163.367
R1023 B.n91 B.n90 163.367
R1024 B.n92 B.n91 163.367
R1025 B.n142 B.n92 163.367
R1026 B.n652 B.n424 163.367
R1027 B.n652 B.n469 163.367
R1028 B.n648 B.n647 163.367
R1029 B.n644 B.n643 163.367
R1030 B.n640 B.n639 163.367
R1031 B.n636 B.n635 163.367
R1032 B.n632 B.n631 163.367
R1033 B.n628 B.n627 163.367
R1034 B.n624 B.n623 163.367
R1035 B.n620 B.n619 163.367
R1036 B.n616 B.n615 163.367
R1037 B.n612 B.n611 163.367
R1038 B.n608 B.n607 163.367
R1039 B.n604 B.n603 163.367
R1040 B.n600 B.n599 163.367
R1041 B.n596 B.n595 163.367
R1042 B.n592 B.n591 163.367
R1043 B.n588 B.n587 163.367
R1044 B.n584 B.n583 163.367
R1045 B.n580 B.n579 163.367
R1046 B.n576 B.n575 163.367
R1047 B.n572 B.n571 163.367
R1048 B.n568 B.n567 163.367
R1049 B.n564 B.n563 163.367
R1050 B.n560 B.n559 163.367
R1051 B.n555 B.n554 163.367
R1052 B.n551 B.n550 163.367
R1053 B.n547 B.n546 163.367
R1054 B.n543 B.n542 163.367
R1055 B.n539 B.n538 163.367
R1056 B.n535 B.n534 163.367
R1057 B.n531 B.n530 163.367
R1058 B.n527 B.n526 163.367
R1059 B.n523 B.n522 163.367
R1060 B.n519 B.n518 163.367
R1061 B.n515 B.n514 163.367
R1062 B.n511 B.n510 163.367
R1063 B.n507 B.n506 163.367
R1064 B.n503 B.n502 163.367
R1065 B.n499 B.n498 163.367
R1066 B.n495 B.n494 163.367
R1067 B.n491 B.n490 163.367
R1068 B.n487 B.n486 163.367
R1069 B.n483 B.n482 163.367
R1070 B.n479 B.n478 163.367
R1071 B.n659 B.n422 163.367
R1072 B.n659 B.n416 163.367
R1073 B.n667 B.n416 163.367
R1074 B.n667 B.n414 163.367
R1075 B.n671 B.n414 163.367
R1076 B.n671 B.n408 163.367
R1077 B.n679 B.n408 163.367
R1078 B.n679 B.n406 163.367
R1079 B.n683 B.n406 163.367
R1080 B.n683 B.n400 163.367
R1081 B.n691 B.n400 163.367
R1082 B.n691 B.n398 163.367
R1083 B.n695 B.n398 163.367
R1084 B.n695 B.n392 163.367
R1085 B.n703 B.n392 163.367
R1086 B.n703 B.n390 163.367
R1087 B.n707 B.n390 163.367
R1088 B.n707 B.n384 163.367
R1089 B.n715 B.n384 163.367
R1090 B.n715 B.n382 163.367
R1091 B.n719 B.n382 163.367
R1092 B.n719 B.n376 163.367
R1093 B.n728 B.n376 163.367
R1094 B.n728 B.n374 163.367
R1095 B.n732 B.n374 163.367
R1096 B.n732 B.n369 163.367
R1097 B.n740 B.n369 163.367
R1098 B.n740 B.n367 163.367
R1099 B.n744 B.n367 163.367
R1100 B.n744 B.n361 163.367
R1101 B.n752 B.n361 163.367
R1102 B.n752 B.n359 163.367
R1103 B.n756 B.n359 163.367
R1104 B.n756 B.n353 163.367
R1105 B.n764 B.n353 163.367
R1106 B.n764 B.n351 163.367
R1107 B.n768 B.n351 163.367
R1108 B.n768 B.n345 163.367
R1109 B.n776 B.n345 163.367
R1110 B.n776 B.n343 163.367
R1111 B.n780 B.n343 163.367
R1112 B.n780 B.n337 163.367
R1113 B.n788 B.n337 163.367
R1114 B.n788 B.n335 163.367
R1115 B.n792 B.n335 163.367
R1116 B.n792 B.n329 163.367
R1117 B.n801 B.n329 163.367
R1118 B.n801 B.n327 163.367
R1119 B.n805 B.n327 163.367
R1120 B.n805 B.n3 163.367
R1121 B.n985 B.n3 163.367
R1122 B.n981 B.n2 163.367
R1123 B.n981 B.n980 163.367
R1124 B.n980 B.n9 163.367
R1125 B.n976 B.n9 163.367
R1126 B.n976 B.n11 163.367
R1127 B.n972 B.n11 163.367
R1128 B.n972 B.n17 163.367
R1129 B.n968 B.n17 163.367
R1130 B.n968 B.n19 163.367
R1131 B.n964 B.n19 163.367
R1132 B.n964 B.n24 163.367
R1133 B.n960 B.n24 163.367
R1134 B.n960 B.n26 163.367
R1135 B.n956 B.n26 163.367
R1136 B.n956 B.n31 163.367
R1137 B.n952 B.n31 163.367
R1138 B.n952 B.n33 163.367
R1139 B.n948 B.n33 163.367
R1140 B.n948 B.n38 163.367
R1141 B.n944 B.n38 163.367
R1142 B.n944 B.n40 163.367
R1143 B.n940 B.n40 163.367
R1144 B.n940 B.n45 163.367
R1145 B.n936 B.n45 163.367
R1146 B.n936 B.n47 163.367
R1147 B.n932 B.n47 163.367
R1148 B.n932 B.n51 163.367
R1149 B.n928 B.n51 163.367
R1150 B.n928 B.n53 163.367
R1151 B.n924 B.n53 163.367
R1152 B.n924 B.n59 163.367
R1153 B.n920 B.n59 163.367
R1154 B.n920 B.n61 163.367
R1155 B.n916 B.n61 163.367
R1156 B.n916 B.n66 163.367
R1157 B.n912 B.n66 163.367
R1158 B.n912 B.n68 163.367
R1159 B.n908 B.n68 163.367
R1160 B.n908 B.n73 163.367
R1161 B.n904 B.n73 163.367
R1162 B.n904 B.n75 163.367
R1163 B.n900 B.n75 163.367
R1164 B.n900 B.n80 163.367
R1165 B.n896 B.n80 163.367
R1166 B.n896 B.n82 163.367
R1167 B.n892 B.n82 163.367
R1168 B.n892 B.n87 163.367
R1169 B.n888 B.n87 163.367
R1170 B.n888 B.n89 163.367
R1171 B.n884 B.n89 163.367
R1172 B.n884 B.n94 163.367
R1173 B.n143 B.t16 118.832
R1174 B.n473 B.t20 118.832
R1175 B.n146 B.t22 118.817
R1176 B.n470 B.t13 118.817
R1177 B.n653 B.n421 73.0537
R1178 B.n878 B.n93 73.0537
R1179 B.n880 B.n879 71.676
R1180 B.n148 B.n97 71.676
R1181 B.n152 B.n98 71.676
R1182 B.n156 B.n99 71.676
R1183 B.n160 B.n100 71.676
R1184 B.n164 B.n101 71.676
R1185 B.n168 B.n102 71.676
R1186 B.n172 B.n103 71.676
R1187 B.n176 B.n104 71.676
R1188 B.n180 B.n105 71.676
R1189 B.n184 B.n106 71.676
R1190 B.n188 B.n107 71.676
R1191 B.n192 B.n108 71.676
R1192 B.n196 B.n109 71.676
R1193 B.n200 B.n110 71.676
R1194 B.n204 B.n111 71.676
R1195 B.n208 B.n112 71.676
R1196 B.n212 B.n113 71.676
R1197 B.n216 B.n114 71.676
R1198 B.n220 B.n115 71.676
R1199 B.n224 B.n116 71.676
R1200 B.n229 B.n117 71.676
R1201 B.n233 B.n118 71.676
R1202 B.n237 B.n119 71.676
R1203 B.n241 B.n120 71.676
R1204 B.n245 B.n121 71.676
R1205 B.n249 B.n122 71.676
R1206 B.n253 B.n123 71.676
R1207 B.n257 B.n124 71.676
R1208 B.n261 B.n125 71.676
R1209 B.n265 B.n126 71.676
R1210 B.n269 B.n127 71.676
R1211 B.n273 B.n128 71.676
R1212 B.n277 B.n129 71.676
R1213 B.n281 B.n130 71.676
R1214 B.n285 B.n131 71.676
R1215 B.n289 B.n132 71.676
R1216 B.n293 B.n133 71.676
R1217 B.n297 B.n134 71.676
R1218 B.n301 B.n135 71.676
R1219 B.n305 B.n136 71.676
R1220 B.n309 B.n137 71.676
R1221 B.n313 B.n138 71.676
R1222 B.n317 B.n139 71.676
R1223 B.n321 B.n140 71.676
R1224 B.n141 B.n140 71.676
R1225 B.n320 B.n139 71.676
R1226 B.n316 B.n138 71.676
R1227 B.n312 B.n137 71.676
R1228 B.n308 B.n136 71.676
R1229 B.n304 B.n135 71.676
R1230 B.n300 B.n134 71.676
R1231 B.n296 B.n133 71.676
R1232 B.n292 B.n132 71.676
R1233 B.n288 B.n131 71.676
R1234 B.n284 B.n130 71.676
R1235 B.n280 B.n129 71.676
R1236 B.n276 B.n128 71.676
R1237 B.n272 B.n127 71.676
R1238 B.n268 B.n126 71.676
R1239 B.n264 B.n125 71.676
R1240 B.n260 B.n124 71.676
R1241 B.n256 B.n123 71.676
R1242 B.n252 B.n122 71.676
R1243 B.n248 B.n121 71.676
R1244 B.n244 B.n120 71.676
R1245 B.n240 B.n119 71.676
R1246 B.n236 B.n118 71.676
R1247 B.n232 B.n117 71.676
R1248 B.n228 B.n116 71.676
R1249 B.n223 B.n115 71.676
R1250 B.n219 B.n114 71.676
R1251 B.n215 B.n113 71.676
R1252 B.n211 B.n112 71.676
R1253 B.n207 B.n111 71.676
R1254 B.n203 B.n110 71.676
R1255 B.n199 B.n109 71.676
R1256 B.n195 B.n108 71.676
R1257 B.n191 B.n107 71.676
R1258 B.n187 B.n106 71.676
R1259 B.n183 B.n105 71.676
R1260 B.n179 B.n104 71.676
R1261 B.n175 B.n103 71.676
R1262 B.n171 B.n102 71.676
R1263 B.n167 B.n101 71.676
R1264 B.n163 B.n100 71.676
R1265 B.n159 B.n99 71.676
R1266 B.n155 B.n98 71.676
R1267 B.n151 B.n97 71.676
R1268 B.n879 B.n96 71.676
R1269 B.n655 B.n654 71.676
R1270 B.n469 B.n425 71.676
R1271 B.n647 B.n426 71.676
R1272 B.n643 B.n427 71.676
R1273 B.n639 B.n428 71.676
R1274 B.n635 B.n429 71.676
R1275 B.n631 B.n430 71.676
R1276 B.n627 B.n431 71.676
R1277 B.n623 B.n432 71.676
R1278 B.n619 B.n433 71.676
R1279 B.n615 B.n434 71.676
R1280 B.n611 B.n435 71.676
R1281 B.n607 B.n436 71.676
R1282 B.n603 B.n437 71.676
R1283 B.n599 B.n438 71.676
R1284 B.n595 B.n439 71.676
R1285 B.n591 B.n440 71.676
R1286 B.n587 B.n441 71.676
R1287 B.n583 B.n442 71.676
R1288 B.n579 B.n443 71.676
R1289 B.n575 B.n444 71.676
R1290 B.n571 B.n445 71.676
R1291 B.n567 B.n446 71.676
R1292 B.n563 B.n447 71.676
R1293 B.n559 B.n448 71.676
R1294 B.n554 B.n449 71.676
R1295 B.n550 B.n450 71.676
R1296 B.n546 B.n451 71.676
R1297 B.n542 B.n452 71.676
R1298 B.n538 B.n453 71.676
R1299 B.n534 B.n454 71.676
R1300 B.n530 B.n455 71.676
R1301 B.n526 B.n456 71.676
R1302 B.n522 B.n457 71.676
R1303 B.n518 B.n458 71.676
R1304 B.n514 B.n459 71.676
R1305 B.n510 B.n460 71.676
R1306 B.n506 B.n461 71.676
R1307 B.n502 B.n462 71.676
R1308 B.n498 B.n463 71.676
R1309 B.n494 B.n464 71.676
R1310 B.n490 B.n465 71.676
R1311 B.n486 B.n466 71.676
R1312 B.n482 B.n467 71.676
R1313 B.n478 B.n468 71.676
R1314 B.n654 B.n424 71.676
R1315 B.n648 B.n425 71.676
R1316 B.n644 B.n426 71.676
R1317 B.n640 B.n427 71.676
R1318 B.n636 B.n428 71.676
R1319 B.n632 B.n429 71.676
R1320 B.n628 B.n430 71.676
R1321 B.n624 B.n431 71.676
R1322 B.n620 B.n432 71.676
R1323 B.n616 B.n433 71.676
R1324 B.n612 B.n434 71.676
R1325 B.n608 B.n435 71.676
R1326 B.n604 B.n436 71.676
R1327 B.n600 B.n437 71.676
R1328 B.n596 B.n438 71.676
R1329 B.n592 B.n439 71.676
R1330 B.n588 B.n440 71.676
R1331 B.n584 B.n441 71.676
R1332 B.n580 B.n442 71.676
R1333 B.n576 B.n443 71.676
R1334 B.n572 B.n444 71.676
R1335 B.n568 B.n445 71.676
R1336 B.n564 B.n446 71.676
R1337 B.n560 B.n447 71.676
R1338 B.n555 B.n448 71.676
R1339 B.n551 B.n449 71.676
R1340 B.n547 B.n450 71.676
R1341 B.n543 B.n451 71.676
R1342 B.n539 B.n452 71.676
R1343 B.n535 B.n453 71.676
R1344 B.n531 B.n454 71.676
R1345 B.n527 B.n455 71.676
R1346 B.n523 B.n456 71.676
R1347 B.n519 B.n457 71.676
R1348 B.n515 B.n458 71.676
R1349 B.n511 B.n459 71.676
R1350 B.n507 B.n460 71.676
R1351 B.n503 B.n461 71.676
R1352 B.n499 B.n462 71.676
R1353 B.n495 B.n463 71.676
R1354 B.n491 B.n464 71.676
R1355 B.n487 B.n465 71.676
R1356 B.n483 B.n466 71.676
R1357 B.n479 B.n467 71.676
R1358 B.n475 B.n468 71.676
R1359 B.n986 B.n985 71.676
R1360 B.n986 B.n2 71.676
R1361 B.n144 B.t17 71.3168
R1362 B.n474 B.t19 71.3168
R1363 B.n147 B.t23 71.3021
R1364 B.n471 B.t12 71.3021
R1365 B.n226 B.n147 59.5399
R1366 B.n145 B.n144 59.5399
R1367 B.n557 B.n474 59.5399
R1368 B.n472 B.n471 59.5399
R1369 B.n147 B.n146 47.5157
R1370 B.n144 B.n143 47.5157
R1371 B.n474 B.n473 47.5157
R1372 B.n471 B.n470 47.5157
R1373 B.n660 B.n421 43.9617
R1374 B.n660 B.n417 43.9617
R1375 B.n666 B.n417 43.9617
R1376 B.n666 B.n413 43.9617
R1377 B.n672 B.n413 43.9617
R1378 B.n672 B.n409 43.9617
R1379 B.n678 B.n409 43.9617
R1380 B.n684 B.n405 43.9617
R1381 B.n684 B.n401 43.9617
R1382 B.n690 B.n401 43.9617
R1383 B.n690 B.n397 43.9617
R1384 B.n696 B.n397 43.9617
R1385 B.n696 B.n393 43.9617
R1386 B.n702 B.n393 43.9617
R1387 B.n702 B.n389 43.9617
R1388 B.n708 B.n389 43.9617
R1389 B.n714 B.n385 43.9617
R1390 B.n714 B.n381 43.9617
R1391 B.n720 B.n381 43.9617
R1392 B.n720 B.n377 43.9617
R1393 B.n727 B.n377 43.9617
R1394 B.n727 B.n726 43.9617
R1395 B.n733 B.n370 43.9617
R1396 B.n739 B.n370 43.9617
R1397 B.n739 B.n366 43.9617
R1398 B.n745 B.n366 43.9617
R1399 B.n745 B.n362 43.9617
R1400 B.n751 B.n362 43.9617
R1401 B.n757 B.n358 43.9617
R1402 B.n757 B.n354 43.9617
R1403 B.n763 B.n354 43.9617
R1404 B.n763 B.n350 43.9617
R1405 B.n769 B.n350 43.9617
R1406 B.n769 B.n346 43.9617
R1407 B.n775 B.n346 43.9617
R1408 B.n781 B.n342 43.9617
R1409 B.n781 B.n338 43.9617
R1410 B.n787 B.n338 43.9617
R1411 B.n787 B.n333 43.9617
R1412 B.n793 B.n333 43.9617
R1413 B.n793 B.n334 43.9617
R1414 B.n800 B.n326 43.9617
R1415 B.n806 B.n326 43.9617
R1416 B.n806 B.n4 43.9617
R1417 B.n984 B.n4 43.9617
R1418 B.n984 B.n983 43.9617
R1419 B.n983 B.n982 43.9617
R1420 B.n982 B.n8 43.9617
R1421 B.n12 B.n8 43.9617
R1422 B.n975 B.n12 43.9617
R1423 B.n974 B.n973 43.9617
R1424 B.n973 B.n16 43.9617
R1425 B.n967 B.n16 43.9617
R1426 B.n967 B.n966 43.9617
R1427 B.n966 B.n965 43.9617
R1428 B.n965 B.n23 43.9617
R1429 B.n959 B.n958 43.9617
R1430 B.n958 B.n957 43.9617
R1431 B.n957 B.n30 43.9617
R1432 B.n951 B.n30 43.9617
R1433 B.n951 B.n950 43.9617
R1434 B.n950 B.n949 43.9617
R1435 B.n949 B.n37 43.9617
R1436 B.n943 B.n942 43.9617
R1437 B.n942 B.n941 43.9617
R1438 B.n941 B.n44 43.9617
R1439 B.n935 B.n44 43.9617
R1440 B.n935 B.n934 43.9617
R1441 B.n934 B.n933 43.9617
R1442 B.n927 B.n54 43.9617
R1443 B.n927 B.n926 43.9617
R1444 B.n926 B.n925 43.9617
R1445 B.n925 B.n58 43.9617
R1446 B.n919 B.n58 43.9617
R1447 B.n919 B.n918 43.9617
R1448 B.n917 B.n65 43.9617
R1449 B.n911 B.n65 43.9617
R1450 B.n911 B.n910 43.9617
R1451 B.n910 B.n909 43.9617
R1452 B.n909 B.n72 43.9617
R1453 B.n903 B.n72 43.9617
R1454 B.n903 B.n902 43.9617
R1455 B.n902 B.n901 43.9617
R1456 B.n901 B.n79 43.9617
R1457 B.n895 B.n894 43.9617
R1458 B.n894 B.n893 43.9617
R1459 B.n893 B.n86 43.9617
R1460 B.n887 B.n86 43.9617
R1461 B.n887 B.n886 43.9617
R1462 B.n886 B.n885 43.9617
R1463 B.n885 B.n93 43.9617
R1464 B.t11 B.n405 41.3758
R1465 B.t15 B.n79 41.3758
R1466 B.t0 B.n342 40.0828
R1467 B.t9 B.n23 40.0828
R1468 B.n751 B.t5 38.7898
R1469 B.n943 B.t4 38.7898
R1470 B.n657 B.n656 32.3127
R1471 B.n476 B.n419 32.3127
R1472 B.n876 B.n875 32.3127
R1473 B.n882 B.n881 32.3127
R1474 B.n800 B.t3 31.0319
R1475 B.n975 B.t2 31.0319
R1476 B.n726 B.t8 29.739
R1477 B.n54 B.t1 29.739
R1478 B.t6 B.n385 23.2741
R1479 B.n918 B.t7 23.2741
R1480 B.n708 B.t6 20.6881
R1481 B.t7 B.n917 20.6881
R1482 B B.n987 18.0485
R1483 B.n733 B.t8 14.2232
R1484 B.n933 B.t1 14.2232
R1485 B.n334 B.t3 12.9303
R1486 B.t2 B.n974 12.9303
R1487 B.n658 B.n657 10.6151
R1488 B.n658 B.n415 10.6151
R1489 B.n668 B.n415 10.6151
R1490 B.n669 B.n668 10.6151
R1491 B.n670 B.n669 10.6151
R1492 B.n670 B.n407 10.6151
R1493 B.n680 B.n407 10.6151
R1494 B.n681 B.n680 10.6151
R1495 B.n682 B.n681 10.6151
R1496 B.n682 B.n399 10.6151
R1497 B.n692 B.n399 10.6151
R1498 B.n693 B.n692 10.6151
R1499 B.n694 B.n693 10.6151
R1500 B.n694 B.n391 10.6151
R1501 B.n704 B.n391 10.6151
R1502 B.n705 B.n704 10.6151
R1503 B.n706 B.n705 10.6151
R1504 B.n706 B.n383 10.6151
R1505 B.n716 B.n383 10.6151
R1506 B.n717 B.n716 10.6151
R1507 B.n718 B.n717 10.6151
R1508 B.n718 B.n375 10.6151
R1509 B.n729 B.n375 10.6151
R1510 B.n730 B.n729 10.6151
R1511 B.n731 B.n730 10.6151
R1512 B.n731 B.n368 10.6151
R1513 B.n741 B.n368 10.6151
R1514 B.n742 B.n741 10.6151
R1515 B.n743 B.n742 10.6151
R1516 B.n743 B.n360 10.6151
R1517 B.n753 B.n360 10.6151
R1518 B.n754 B.n753 10.6151
R1519 B.n755 B.n754 10.6151
R1520 B.n755 B.n352 10.6151
R1521 B.n765 B.n352 10.6151
R1522 B.n766 B.n765 10.6151
R1523 B.n767 B.n766 10.6151
R1524 B.n767 B.n344 10.6151
R1525 B.n777 B.n344 10.6151
R1526 B.n778 B.n777 10.6151
R1527 B.n779 B.n778 10.6151
R1528 B.n779 B.n336 10.6151
R1529 B.n789 B.n336 10.6151
R1530 B.n790 B.n789 10.6151
R1531 B.n791 B.n790 10.6151
R1532 B.n791 B.n328 10.6151
R1533 B.n802 B.n328 10.6151
R1534 B.n803 B.n802 10.6151
R1535 B.n804 B.n803 10.6151
R1536 B.n804 B.n0 10.6151
R1537 B.n656 B.n423 10.6151
R1538 B.n651 B.n423 10.6151
R1539 B.n651 B.n650 10.6151
R1540 B.n650 B.n649 10.6151
R1541 B.n649 B.n646 10.6151
R1542 B.n646 B.n645 10.6151
R1543 B.n645 B.n642 10.6151
R1544 B.n642 B.n641 10.6151
R1545 B.n641 B.n638 10.6151
R1546 B.n638 B.n637 10.6151
R1547 B.n637 B.n634 10.6151
R1548 B.n634 B.n633 10.6151
R1549 B.n633 B.n630 10.6151
R1550 B.n630 B.n629 10.6151
R1551 B.n629 B.n626 10.6151
R1552 B.n626 B.n625 10.6151
R1553 B.n625 B.n622 10.6151
R1554 B.n622 B.n621 10.6151
R1555 B.n621 B.n618 10.6151
R1556 B.n618 B.n617 10.6151
R1557 B.n617 B.n614 10.6151
R1558 B.n614 B.n613 10.6151
R1559 B.n613 B.n610 10.6151
R1560 B.n610 B.n609 10.6151
R1561 B.n609 B.n606 10.6151
R1562 B.n606 B.n605 10.6151
R1563 B.n605 B.n602 10.6151
R1564 B.n602 B.n601 10.6151
R1565 B.n601 B.n598 10.6151
R1566 B.n598 B.n597 10.6151
R1567 B.n597 B.n594 10.6151
R1568 B.n594 B.n593 10.6151
R1569 B.n593 B.n590 10.6151
R1570 B.n590 B.n589 10.6151
R1571 B.n589 B.n586 10.6151
R1572 B.n586 B.n585 10.6151
R1573 B.n585 B.n582 10.6151
R1574 B.n582 B.n581 10.6151
R1575 B.n581 B.n578 10.6151
R1576 B.n578 B.n577 10.6151
R1577 B.n574 B.n573 10.6151
R1578 B.n573 B.n570 10.6151
R1579 B.n570 B.n569 10.6151
R1580 B.n569 B.n566 10.6151
R1581 B.n566 B.n565 10.6151
R1582 B.n565 B.n562 10.6151
R1583 B.n562 B.n561 10.6151
R1584 B.n561 B.n558 10.6151
R1585 B.n556 B.n553 10.6151
R1586 B.n553 B.n552 10.6151
R1587 B.n552 B.n549 10.6151
R1588 B.n549 B.n548 10.6151
R1589 B.n548 B.n545 10.6151
R1590 B.n545 B.n544 10.6151
R1591 B.n544 B.n541 10.6151
R1592 B.n541 B.n540 10.6151
R1593 B.n540 B.n537 10.6151
R1594 B.n537 B.n536 10.6151
R1595 B.n536 B.n533 10.6151
R1596 B.n533 B.n532 10.6151
R1597 B.n532 B.n529 10.6151
R1598 B.n529 B.n528 10.6151
R1599 B.n528 B.n525 10.6151
R1600 B.n525 B.n524 10.6151
R1601 B.n524 B.n521 10.6151
R1602 B.n521 B.n520 10.6151
R1603 B.n520 B.n517 10.6151
R1604 B.n517 B.n516 10.6151
R1605 B.n516 B.n513 10.6151
R1606 B.n513 B.n512 10.6151
R1607 B.n512 B.n509 10.6151
R1608 B.n509 B.n508 10.6151
R1609 B.n508 B.n505 10.6151
R1610 B.n505 B.n504 10.6151
R1611 B.n504 B.n501 10.6151
R1612 B.n501 B.n500 10.6151
R1613 B.n500 B.n497 10.6151
R1614 B.n497 B.n496 10.6151
R1615 B.n496 B.n493 10.6151
R1616 B.n493 B.n492 10.6151
R1617 B.n492 B.n489 10.6151
R1618 B.n489 B.n488 10.6151
R1619 B.n488 B.n485 10.6151
R1620 B.n485 B.n484 10.6151
R1621 B.n484 B.n481 10.6151
R1622 B.n481 B.n480 10.6151
R1623 B.n480 B.n477 10.6151
R1624 B.n477 B.n476 10.6151
R1625 B.n662 B.n419 10.6151
R1626 B.n663 B.n662 10.6151
R1627 B.n664 B.n663 10.6151
R1628 B.n664 B.n411 10.6151
R1629 B.n674 B.n411 10.6151
R1630 B.n675 B.n674 10.6151
R1631 B.n676 B.n675 10.6151
R1632 B.n676 B.n403 10.6151
R1633 B.n686 B.n403 10.6151
R1634 B.n687 B.n686 10.6151
R1635 B.n688 B.n687 10.6151
R1636 B.n688 B.n395 10.6151
R1637 B.n698 B.n395 10.6151
R1638 B.n699 B.n698 10.6151
R1639 B.n700 B.n699 10.6151
R1640 B.n700 B.n387 10.6151
R1641 B.n710 B.n387 10.6151
R1642 B.n711 B.n710 10.6151
R1643 B.n712 B.n711 10.6151
R1644 B.n712 B.n379 10.6151
R1645 B.n722 B.n379 10.6151
R1646 B.n723 B.n722 10.6151
R1647 B.n724 B.n723 10.6151
R1648 B.n724 B.n372 10.6151
R1649 B.n735 B.n372 10.6151
R1650 B.n736 B.n735 10.6151
R1651 B.n737 B.n736 10.6151
R1652 B.n737 B.n364 10.6151
R1653 B.n747 B.n364 10.6151
R1654 B.n748 B.n747 10.6151
R1655 B.n749 B.n748 10.6151
R1656 B.n749 B.n356 10.6151
R1657 B.n759 B.n356 10.6151
R1658 B.n760 B.n759 10.6151
R1659 B.n761 B.n760 10.6151
R1660 B.n761 B.n348 10.6151
R1661 B.n771 B.n348 10.6151
R1662 B.n772 B.n771 10.6151
R1663 B.n773 B.n772 10.6151
R1664 B.n773 B.n340 10.6151
R1665 B.n783 B.n340 10.6151
R1666 B.n784 B.n783 10.6151
R1667 B.n785 B.n784 10.6151
R1668 B.n785 B.n331 10.6151
R1669 B.n795 B.n331 10.6151
R1670 B.n796 B.n795 10.6151
R1671 B.n798 B.n796 10.6151
R1672 B.n798 B.n797 10.6151
R1673 B.n797 B.n324 10.6151
R1674 B.n809 B.n324 10.6151
R1675 B.n810 B.n809 10.6151
R1676 B.n811 B.n810 10.6151
R1677 B.n812 B.n811 10.6151
R1678 B.n813 B.n812 10.6151
R1679 B.n816 B.n813 10.6151
R1680 B.n817 B.n816 10.6151
R1681 B.n818 B.n817 10.6151
R1682 B.n819 B.n818 10.6151
R1683 B.n821 B.n819 10.6151
R1684 B.n822 B.n821 10.6151
R1685 B.n823 B.n822 10.6151
R1686 B.n824 B.n823 10.6151
R1687 B.n826 B.n824 10.6151
R1688 B.n827 B.n826 10.6151
R1689 B.n828 B.n827 10.6151
R1690 B.n829 B.n828 10.6151
R1691 B.n831 B.n829 10.6151
R1692 B.n832 B.n831 10.6151
R1693 B.n833 B.n832 10.6151
R1694 B.n834 B.n833 10.6151
R1695 B.n836 B.n834 10.6151
R1696 B.n837 B.n836 10.6151
R1697 B.n838 B.n837 10.6151
R1698 B.n839 B.n838 10.6151
R1699 B.n841 B.n839 10.6151
R1700 B.n842 B.n841 10.6151
R1701 B.n843 B.n842 10.6151
R1702 B.n844 B.n843 10.6151
R1703 B.n846 B.n844 10.6151
R1704 B.n847 B.n846 10.6151
R1705 B.n848 B.n847 10.6151
R1706 B.n849 B.n848 10.6151
R1707 B.n851 B.n849 10.6151
R1708 B.n852 B.n851 10.6151
R1709 B.n853 B.n852 10.6151
R1710 B.n854 B.n853 10.6151
R1711 B.n856 B.n854 10.6151
R1712 B.n857 B.n856 10.6151
R1713 B.n858 B.n857 10.6151
R1714 B.n859 B.n858 10.6151
R1715 B.n861 B.n859 10.6151
R1716 B.n862 B.n861 10.6151
R1717 B.n863 B.n862 10.6151
R1718 B.n864 B.n863 10.6151
R1719 B.n866 B.n864 10.6151
R1720 B.n867 B.n866 10.6151
R1721 B.n868 B.n867 10.6151
R1722 B.n869 B.n868 10.6151
R1723 B.n871 B.n869 10.6151
R1724 B.n872 B.n871 10.6151
R1725 B.n873 B.n872 10.6151
R1726 B.n874 B.n873 10.6151
R1727 B.n875 B.n874 10.6151
R1728 B.n979 B.n1 10.6151
R1729 B.n979 B.n978 10.6151
R1730 B.n978 B.n977 10.6151
R1731 B.n977 B.n10 10.6151
R1732 B.n971 B.n10 10.6151
R1733 B.n971 B.n970 10.6151
R1734 B.n970 B.n969 10.6151
R1735 B.n969 B.n18 10.6151
R1736 B.n963 B.n18 10.6151
R1737 B.n963 B.n962 10.6151
R1738 B.n962 B.n961 10.6151
R1739 B.n961 B.n25 10.6151
R1740 B.n955 B.n25 10.6151
R1741 B.n955 B.n954 10.6151
R1742 B.n954 B.n953 10.6151
R1743 B.n953 B.n32 10.6151
R1744 B.n947 B.n32 10.6151
R1745 B.n947 B.n946 10.6151
R1746 B.n946 B.n945 10.6151
R1747 B.n945 B.n39 10.6151
R1748 B.n939 B.n39 10.6151
R1749 B.n939 B.n938 10.6151
R1750 B.n938 B.n937 10.6151
R1751 B.n937 B.n46 10.6151
R1752 B.n931 B.n46 10.6151
R1753 B.n931 B.n930 10.6151
R1754 B.n930 B.n929 10.6151
R1755 B.n929 B.n52 10.6151
R1756 B.n923 B.n52 10.6151
R1757 B.n923 B.n922 10.6151
R1758 B.n922 B.n921 10.6151
R1759 B.n921 B.n60 10.6151
R1760 B.n915 B.n60 10.6151
R1761 B.n915 B.n914 10.6151
R1762 B.n914 B.n913 10.6151
R1763 B.n913 B.n67 10.6151
R1764 B.n907 B.n67 10.6151
R1765 B.n907 B.n906 10.6151
R1766 B.n906 B.n905 10.6151
R1767 B.n905 B.n74 10.6151
R1768 B.n899 B.n74 10.6151
R1769 B.n899 B.n898 10.6151
R1770 B.n898 B.n897 10.6151
R1771 B.n897 B.n81 10.6151
R1772 B.n891 B.n81 10.6151
R1773 B.n891 B.n890 10.6151
R1774 B.n890 B.n889 10.6151
R1775 B.n889 B.n88 10.6151
R1776 B.n883 B.n88 10.6151
R1777 B.n883 B.n882 10.6151
R1778 B.n881 B.n95 10.6151
R1779 B.n149 B.n95 10.6151
R1780 B.n150 B.n149 10.6151
R1781 B.n153 B.n150 10.6151
R1782 B.n154 B.n153 10.6151
R1783 B.n157 B.n154 10.6151
R1784 B.n158 B.n157 10.6151
R1785 B.n161 B.n158 10.6151
R1786 B.n162 B.n161 10.6151
R1787 B.n165 B.n162 10.6151
R1788 B.n166 B.n165 10.6151
R1789 B.n169 B.n166 10.6151
R1790 B.n170 B.n169 10.6151
R1791 B.n173 B.n170 10.6151
R1792 B.n174 B.n173 10.6151
R1793 B.n177 B.n174 10.6151
R1794 B.n178 B.n177 10.6151
R1795 B.n181 B.n178 10.6151
R1796 B.n182 B.n181 10.6151
R1797 B.n185 B.n182 10.6151
R1798 B.n186 B.n185 10.6151
R1799 B.n189 B.n186 10.6151
R1800 B.n190 B.n189 10.6151
R1801 B.n193 B.n190 10.6151
R1802 B.n194 B.n193 10.6151
R1803 B.n197 B.n194 10.6151
R1804 B.n198 B.n197 10.6151
R1805 B.n201 B.n198 10.6151
R1806 B.n202 B.n201 10.6151
R1807 B.n205 B.n202 10.6151
R1808 B.n206 B.n205 10.6151
R1809 B.n209 B.n206 10.6151
R1810 B.n210 B.n209 10.6151
R1811 B.n213 B.n210 10.6151
R1812 B.n214 B.n213 10.6151
R1813 B.n217 B.n214 10.6151
R1814 B.n218 B.n217 10.6151
R1815 B.n221 B.n218 10.6151
R1816 B.n222 B.n221 10.6151
R1817 B.n225 B.n222 10.6151
R1818 B.n230 B.n227 10.6151
R1819 B.n231 B.n230 10.6151
R1820 B.n234 B.n231 10.6151
R1821 B.n235 B.n234 10.6151
R1822 B.n238 B.n235 10.6151
R1823 B.n239 B.n238 10.6151
R1824 B.n242 B.n239 10.6151
R1825 B.n243 B.n242 10.6151
R1826 B.n247 B.n246 10.6151
R1827 B.n250 B.n247 10.6151
R1828 B.n251 B.n250 10.6151
R1829 B.n254 B.n251 10.6151
R1830 B.n255 B.n254 10.6151
R1831 B.n258 B.n255 10.6151
R1832 B.n259 B.n258 10.6151
R1833 B.n262 B.n259 10.6151
R1834 B.n263 B.n262 10.6151
R1835 B.n266 B.n263 10.6151
R1836 B.n267 B.n266 10.6151
R1837 B.n270 B.n267 10.6151
R1838 B.n271 B.n270 10.6151
R1839 B.n274 B.n271 10.6151
R1840 B.n275 B.n274 10.6151
R1841 B.n278 B.n275 10.6151
R1842 B.n279 B.n278 10.6151
R1843 B.n282 B.n279 10.6151
R1844 B.n283 B.n282 10.6151
R1845 B.n286 B.n283 10.6151
R1846 B.n287 B.n286 10.6151
R1847 B.n290 B.n287 10.6151
R1848 B.n291 B.n290 10.6151
R1849 B.n294 B.n291 10.6151
R1850 B.n295 B.n294 10.6151
R1851 B.n298 B.n295 10.6151
R1852 B.n299 B.n298 10.6151
R1853 B.n302 B.n299 10.6151
R1854 B.n303 B.n302 10.6151
R1855 B.n306 B.n303 10.6151
R1856 B.n307 B.n306 10.6151
R1857 B.n310 B.n307 10.6151
R1858 B.n311 B.n310 10.6151
R1859 B.n314 B.n311 10.6151
R1860 B.n315 B.n314 10.6151
R1861 B.n318 B.n315 10.6151
R1862 B.n319 B.n318 10.6151
R1863 B.n322 B.n319 10.6151
R1864 B.n323 B.n322 10.6151
R1865 B.n876 B.n323 10.6151
R1866 B.n987 B.n0 8.11757
R1867 B.n987 B.n1 8.11757
R1868 B.n574 B.n472 6.5566
R1869 B.n558 B.n557 6.5566
R1870 B.n227 B.n226 6.5566
R1871 B.n243 B.n145 6.5566
R1872 B.t5 B.n358 5.17241
R1873 B.t4 B.n37 5.17241
R1874 B.n577 B.n472 4.05904
R1875 B.n557 B.n556 4.05904
R1876 B.n226 B.n225 4.05904
R1877 B.n246 B.n145 4.05904
R1878 B.n775 B.t0 3.87943
R1879 B.n959 B.t9 3.87943
R1880 B.n678 B.t11 2.58645
R1881 B.n895 B.t15 2.58645
R1882 VN.n8 VN.t7 167.464
R1883 VN.n41 VN.t5 167.464
R1884 VN.n63 VN.n33 161.3
R1885 VN.n62 VN.n61 161.3
R1886 VN.n60 VN.n34 161.3
R1887 VN.n59 VN.n58 161.3
R1888 VN.n57 VN.n35 161.3
R1889 VN.n55 VN.n54 161.3
R1890 VN.n53 VN.n36 161.3
R1891 VN.n52 VN.n51 161.3
R1892 VN.n50 VN.n37 161.3
R1893 VN.n49 VN.n48 161.3
R1894 VN.n47 VN.n38 161.3
R1895 VN.n46 VN.n45 161.3
R1896 VN.n44 VN.n39 161.3
R1897 VN.n43 VN.n42 161.3
R1898 VN.n30 VN.n0 161.3
R1899 VN.n29 VN.n28 161.3
R1900 VN.n27 VN.n1 161.3
R1901 VN.n26 VN.n25 161.3
R1902 VN.n24 VN.n2 161.3
R1903 VN.n22 VN.n21 161.3
R1904 VN.n20 VN.n3 161.3
R1905 VN.n19 VN.n18 161.3
R1906 VN.n17 VN.n4 161.3
R1907 VN.n16 VN.n15 161.3
R1908 VN.n14 VN.n5 161.3
R1909 VN.n13 VN.n12 161.3
R1910 VN.n11 VN.n6 161.3
R1911 VN.n10 VN.n9 161.3
R1912 VN.n16 VN.t4 133.459
R1913 VN.n7 VN.t6 133.459
R1914 VN.n23 VN.t0 133.459
R1915 VN.n31 VN.t9 133.459
R1916 VN.n49 VN.t1 133.459
R1917 VN.n40 VN.t2 133.459
R1918 VN.n56 VN.t8 133.459
R1919 VN.n64 VN.t3 133.459
R1920 VN.n32 VN.n31 91.1314
R1921 VN.n65 VN.n64 91.1314
R1922 VN.n12 VN.n11 56.4773
R1923 VN.n18 VN.n3 56.4773
R1924 VN.n29 VN.n1 56.4773
R1925 VN.n45 VN.n44 56.4773
R1926 VN.n51 VN.n36 56.4773
R1927 VN.n62 VN.n34 56.4773
R1928 VN VN.n65 50.6383
R1929 VN.n8 VN.n7 48.3597
R1930 VN.n41 VN.n40 48.3597
R1931 VN.n11 VN.n10 24.3439
R1932 VN.n12 VN.n5 24.3439
R1933 VN.n16 VN.n5 24.3439
R1934 VN.n17 VN.n16 24.3439
R1935 VN.n18 VN.n17 24.3439
R1936 VN.n22 VN.n3 24.3439
R1937 VN.n25 VN.n24 24.3439
R1938 VN.n25 VN.n1 24.3439
R1939 VN.n30 VN.n29 24.3439
R1940 VN.n44 VN.n43 24.3439
R1941 VN.n51 VN.n50 24.3439
R1942 VN.n50 VN.n49 24.3439
R1943 VN.n49 VN.n38 24.3439
R1944 VN.n45 VN.n38 24.3439
R1945 VN.n58 VN.n34 24.3439
R1946 VN.n58 VN.n57 24.3439
R1947 VN.n55 VN.n36 24.3439
R1948 VN.n63 VN.n62 24.3439
R1949 VN.n10 VN.n7 21.9096
R1950 VN.n23 VN.n22 21.9096
R1951 VN.n43 VN.n40 21.9096
R1952 VN.n56 VN.n55 21.9096
R1953 VN.n31 VN.n30 19.4752
R1954 VN.n64 VN.n63 19.4752
R1955 VN.n42 VN.n41 9.03227
R1956 VN.n9 VN.n8 9.03227
R1957 VN.n24 VN.n23 2.43484
R1958 VN.n57 VN.n56 2.43484
R1959 VN.n65 VN.n33 0.278398
R1960 VN.n32 VN.n0 0.278398
R1961 VN.n61 VN.n33 0.189894
R1962 VN.n61 VN.n60 0.189894
R1963 VN.n60 VN.n59 0.189894
R1964 VN.n59 VN.n35 0.189894
R1965 VN.n54 VN.n35 0.189894
R1966 VN.n54 VN.n53 0.189894
R1967 VN.n53 VN.n52 0.189894
R1968 VN.n52 VN.n37 0.189894
R1969 VN.n48 VN.n37 0.189894
R1970 VN.n48 VN.n47 0.189894
R1971 VN.n47 VN.n46 0.189894
R1972 VN.n46 VN.n39 0.189894
R1973 VN.n42 VN.n39 0.189894
R1974 VN.n9 VN.n6 0.189894
R1975 VN.n13 VN.n6 0.189894
R1976 VN.n14 VN.n13 0.189894
R1977 VN.n15 VN.n14 0.189894
R1978 VN.n15 VN.n4 0.189894
R1979 VN.n19 VN.n4 0.189894
R1980 VN.n20 VN.n19 0.189894
R1981 VN.n21 VN.n20 0.189894
R1982 VN.n21 VN.n2 0.189894
R1983 VN.n26 VN.n2 0.189894
R1984 VN.n27 VN.n26 0.189894
R1985 VN.n28 VN.n27 0.189894
R1986 VN.n28 VN.n0 0.189894
R1987 VN VN.n32 0.153422
R1988 VDD2.n1 VDD2.t2 65.3905
R1989 VDD2.n4 VDD2.t6 63.2787
R1990 VDD2.n3 VDD2.n2 63.1206
R1991 VDD2 VDD2.n7 63.1178
R1992 VDD2.n6 VDD2.n5 61.5921
R1993 VDD2.n1 VDD2.n0 61.5919
R1994 VDD2.n4 VDD2.n3 43.8683
R1995 VDD2.n6 VDD2.n4 2.11257
R1996 VDD2.n7 VDD2.t7 1.68704
R1997 VDD2.n7 VDD2.t4 1.68704
R1998 VDD2.n5 VDD2.t1 1.68704
R1999 VDD2.n5 VDD2.t8 1.68704
R2000 VDD2.n2 VDD2.t9 1.68704
R2001 VDD2.n2 VDD2.t0 1.68704
R2002 VDD2.n0 VDD2.t3 1.68704
R2003 VDD2.n0 VDD2.t5 1.68704
R2004 VDD2 VDD2.n6 0.586707
R2005 VDD2.n3 VDD2.n1 0.473171
C0 VDD2 VTAIL 10.316299f
C1 VDD1 VN 0.152082f
C2 VN VP 7.6487f
C3 VN VTAIL 10.437201f
C4 VDD2 VN 9.98429f
C5 VDD1 VP 10.3505f
C6 VDD1 VTAIL 10.269099f
C7 VDD2 VDD1 1.86312f
C8 VTAIL VP 10.4516f
C9 VDD2 VP 0.522166f
C10 VDD2 B 6.576189f
C11 VDD1 B 6.569395f
C12 VTAIL B 7.73404f
C13 VN B 15.859269f
C14 VP B 14.343278f
C15 VDD2.t2 B 2.34316f
C16 VDD2.t3 B 0.205477f
C17 VDD2.t5 B 0.205477f
C18 VDD2.n0 B 1.82798f
C19 VDD2.n1 B 0.757449f
C20 VDD2.t9 B 0.205477f
C21 VDD2.t0 B 0.205477f
C22 VDD2.n2 B 1.83894f
C23 VDD2.n3 B 2.33824f
C24 VDD2.t6 B 2.3302f
C25 VDD2.n4 B 2.58538f
C26 VDD2.t1 B 0.205477f
C27 VDD2.t8 B 0.205477f
C28 VDD2.n5 B 1.82799f
C29 VDD2.n6 B 0.376078f
C30 VDD2.t7 B 0.205477f
C31 VDD2.t4 B 0.205477f
C32 VDD2.n7 B 1.83891f
C33 VN.n0 B 0.032134f
C34 VN.t9 B 1.65171f
C35 VN.n1 B 0.030604f
C36 VN.n2 B 0.024372f
C37 VN.t0 B 1.65171f
C38 VN.n3 B 0.037444f
C39 VN.n4 B 0.024372f
C40 VN.t4 B 1.65171f
C41 VN.n5 B 0.045652f
C42 VN.n6 B 0.024372f
C43 VN.t6 B 1.65171f
C44 VN.n7 B 0.660204f
C45 VN.t7 B 1.79835f
C46 VN.n8 B 0.643049f
C47 VN.n9 B 0.20563f
C48 VN.n10 B 0.043398f
C49 VN.n11 B 0.037444f
C50 VN.n12 B 0.034024f
C51 VN.n13 B 0.024372f
C52 VN.n14 B 0.024372f
C53 VN.n15 B 0.024372f
C54 VN.n16 B 0.612311f
C55 VN.n17 B 0.045652f
C56 VN.n18 B 0.034024f
C57 VN.n19 B 0.024372f
C58 VN.n20 B 0.024372f
C59 VN.n21 B 0.024372f
C60 VN.n22 B 0.043398f
C61 VN.n23 B 0.5892f
C62 VN.n24 B 0.025366f
C63 VN.n25 B 0.045652f
C64 VN.n26 B 0.024372f
C65 VN.n27 B 0.024372f
C66 VN.n28 B 0.024372f
C67 VN.n29 B 0.040864f
C68 VN.n30 B 0.041144f
C69 VN.n31 B 0.668462f
C70 VN.n32 B 0.030232f
C71 VN.n33 B 0.032134f
C72 VN.t3 B 1.65171f
C73 VN.n34 B 0.030604f
C74 VN.n35 B 0.024372f
C75 VN.t8 B 1.65171f
C76 VN.n36 B 0.037444f
C77 VN.n37 B 0.024372f
C78 VN.t1 B 1.65171f
C79 VN.n38 B 0.045652f
C80 VN.n39 B 0.024372f
C81 VN.t2 B 1.65171f
C82 VN.n40 B 0.660204f
C83 VN.t5 B 1.79835f
C84 VN.n41 B 0.643049f
C85 VN.n42 B 0.20563f
C86 VN.n43 B 0.043398f
C87 VN.n44 B 0.037444f
C88 VN.n45 B 0.034024f
C89 VN.n46 B 0.024372f
C90 VN.n47 B 0.024372f
C91 VN.n48 B 0.024372f
C92 VN.n49 B 0.612311f
C93 VN.n50 B 0.045652f
C94 VN.n51 B 0.034024f
C95 VN.n52 B 0.024372f
C96 VN.n53 B 0.024372f
C97 VN.n54 B 0.024372f
C98 VN.n55 B 0.043398f
C99 VN.n56 B 0.5892f
C100 VN.n57 B 0.025366f
C101 VN.n58 B 0.045652f
C102 VN.n59 B 0.024372f
C103 VN.n60 B 0.024372f
C104 VN.n61 B 0.024372f
C105 VN.n62 B 0.040864f
C106 VN.n63 B 0.041144f
C107 VN.n64 B 0.668462f
C108 VN.n65 B 1.37395f
C109 VDD1.t5 B 2.37974f
C110 VDD1.t8 B 0.208684f
C111 VDD1.t0 B 0.208684f
C112 VDD1.n0 B 1.85653f
C113 VDD1.n1 B 0.776392f
C114 VDD1.t3 B 2.37974f
C115 VDD1.t1 B 0.208684f
C116 VDD1.t9 B 0.208684f
C117 VDD1.n2 B 1.85652f
C118 VDD1.n3 B 0.769274f
C119 VDD1.t4 B 0.208684f
C120 VDD1.t2 B 0.208684f
C121 VDD1.n4 B 1.86765f
C122 VDD1.n5 B 2.47567f
C123 VDD1.t6 B 0.208684f
C124 VDD1.t7 B 0.208684f
C125 VDD1.n6 B 1.85652f
C126 VDD1.n7 B 2.6594f
C127 VTAIL.t2 B 0.229535f
C128 VTAIL.t19 B 0.229535f
C129 VTAIL.n0 B 1.96764f
C130 VTAIL.n1 B 0.498324f
C131 VTAIL.t13 B 2.50808f
C132 VTAIL.n2 B 0.621343f
C133 VTAIL.t12 B 0.229535f
C134 VTAIL.t15 B 0.229535f
C135 VTAIL.n3 B 1.96764f
C136 VTAIL.n4 B 0.582514f
C137 VTAIL.t18 B 0.229535f
C138 VTAIL.t16 B 0.229535f
C139 VTAIL.n5 B 1.96764f
C140 VTAIL.n6 B 1.89383f
C141 VTAIL.t6 B 0.229535f
C142 VTAIL.t8 B 0.229535f
C143 VTAIL.n7 B 1.96765f
C144 VTAIL.n8 B 1.89383f
C145 VTAIL.t5 B 0.229535f
C146 VTAIL.t0 B 0.229535f
C147 VTAIL.n9 B 1.96765f
C148 VTAIL.n10 B 0.582508f
C149 VTAIL.t3 B 2.50809f
C150 VTAIL.n11 B 0.621336f
C151 VTAIL.t11 B 0.229535f
C152 VTAIL.t14 B 0.229535f
C153 VTAIL.n12 B 1.96765f
C154 VTAIL.n13 B 0.535774f
C155 VTAIL.t17 B 0.229535f
C156 VTAIL.t9 B 0.229535f
C157 VTAIL.n14 B 1.96765f
C158 VTAIL.n15 B 0.582508f
C159 VTAIL.t10 B 2.50808f
C160 VTAIL.n16 B 1.81101f
C161 VTAIL.t7 B 2.50808f
C162 VTAIL.n17 B 1.81101f
C163 VTAIL.t4 B 0.229535f
C164 VTAIL.t1 B 0.229535f
C165 VTAIL.n18 B 1.96764f
C166 VTAIL.n19 B 0.45159f
C167 VP.n0 B 0.032748f
C168 VP.t7 B 1.68327f
C169 VP.n1 B 0.031189f
C170 VP.n2 B 0.024838f
C171 VP.t5 B 1.68327f
C172 VP.n3 B 0.03816f
C173 VP.n4 B 0.024838f
C174 VP.t0 B 1.68327f
C175 VP.n5 B 0.046524f
C176 VP.n6 B 0.024838f
C177 VP.t8 B 1.68327f
C178 VP.n7 B 0.600456f
C179 VP.n8 B 0.024838f
C180 VP.n9 B 0.041645f
C181 VP.n10 B 0.032748f
C182 VP.t2 B 1.68327f
C183 VP.n11 B 0.031189f
C184 VP.n12 B 0.024838f
C185 VP.t3 B 1.68327f
C186 VP.n13 B 0.038159f
C187 VP.n14 B 0.024838f
C188 VP.t9 B 1.68327f
C189 VP.n15 B 0.046524f
C190 VP.n16 B 0.024838f
C191 VP.t1 B 1.68327f
C192 VP.n17 B 0.672817f
C193 VP.t4 B 1.83271f
C194 VP.n18 B 0.655334f
C195 VP.n19 B 0.209558f
C196 VP.n20 B 0.044227f
C197 VP.n21 B 0.03816f
C198 VP.n22 B 0.034674f
C199 VP.n23 B 0.024838f
C200 VP.n24 B 0.024838f
C201 VP.n25 B 0.024838f
C202 VP.n26 B 0.624009f
C203 VP.n27 B 0.046524f
C204 VP.n28 B 0.034674f
C205 VP.n29 B 0.024838f
C206 VP.n30 B 0.024838f
C207 VP.n31 B 0.024838f
C208 VP.n32 B 0.044227f
C209 VP.n33 B 0.600456f
C210 VP.n34 B 0.02585f
C211 VP.n35 B 0.046524f
C212 VP.n36 B 0.024838f
C213 VP.n37 B 0.024838f
C214 VP.n38 B 0.024838f
C215 VP.n39 B 0.041645f
C216 VP.n40 B 0.04193f
C217 VP.n41 B 0.681232f
C218 VP.n42 B 1.38687f
C219 VP.n43 B 1.40455f
C220 VP.t6 B 1.68327f
C221 VP.n44 B 0.681232f
C222 VP.n45 B 0.04193f
C223 VP.n46 B 0.032748f
C224 VP.n47 B 0.024838f
C225 VP.n48 B 0.024838f
C226 VP.n49 B 0.031189f
C227 VP.n50 B 0.046524f
C228 VP.n51 B 0.02585f
C229 VP.n52 B 0.024838f
C230 VP.n53 B 0.024838f
C231 VP.n54 B 0.044227f
C232 VP.n55 B 0.038159f
C233 VP.n56 B 0.034674f
C234 VP.n57 B 0.024838f
C235 VP.n58 B 0.024838f
C236 VP.n59 B 0.024838f
C237 VP.n60 B 0.624009f
C238 VP.n61 B 0.046524f
C239 VP.n62 B 0.034674f
C240 VP.n63 B 0.024838f
C241 VP.n64 B 0.024838f
C242 VP.n65 B 0.024838f
C243 VP.n66 B 0.044227f
C244 VP.n67 B 0.600456f
C245 VP.n68 B 0.02585f
C246 VP.n69 B 0.046524f
C247 VP.n70 B 0.024838f
C248 VP.n71 B 0.024838f
C249 VP.n72 B 0.024838f
C250 VP.n73 B 0.041645f
C251 VP.n74 B 0.04193f
C252 VP.n75 B 0.681232f
C253 VP.n76 B 0.030809f
.ends

