* NGSPICE file created from diff_pair_sample_1501.ext - technology: sky130A

.subckt diff_pair_sample_1501 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t9 VN.t0 VTAIL.t17 w_n5830_n1814# sky130_fd_pr__pfet_01v8 ad=0.69795 pd=4.56 as=1.6497 ps=9.24 w=4.23 l=3.72
X1 VTAIL.t11 VN.t1 VDD2.t8 w_n5830_n1814# sky130_fd_pr__pfet_01v8 ad=0.69795 pd=4.56 as=0.69795 ps=4.56 w=4.23 l=3.72
X2 VDD1.t9 VP.t0 VTAIL.t5 w_n5830_n1814# sky130_fd_pr__pfet_01v8 ad=1.6497 pd=9.24 as=0.69795 ps=4.56 w=4.23 l=3.72
X3 VDD2.t7 VN.t2 VTAIL.t15 w_n5830_n1814# sky130_fd_pr__pfet_01v8 ad=0.69795 pd=4.56 as=0.69795 ps=4.56 w=4.23 l=3.72
X4 VTAIL.t18 VP.t1 VDD1.t8 w_n5830_n1814# sky130_fd_pr__pfet_01v8 ad=0.69795 pd=4.56 as=0.69795 ps=4.56 w=4.23 l=3.72
X5 VTAIL.t7 VP.t2 VDD1.t7 w_n5830_n1814# sky130_fd_pr__pfet_01v8 ad=0.69795 pd=4.56 as=0.69795 ps=4.56 w=4.23 l=3.72
X6 VDD2.t6 VN.t3 VTAIL.t16 w_n5830_n1814# sky130_fd_pr__pfet_01v8 ad=0.69795 pd=4.56 as=0.69795 ps=4.56 w=4.23 l=3.72
X7 VDD1.t6 VP.t3 VTAIL.t1 w_n5830_n1814# sky130_fd_pr__pfet_01v8 ad=0.69795 pd=4.56 as=0.69795 ps=4.56 w=4.23 l=3.72
X8 VTAIL.t9 VN.t4 VDD2.t5 w_n5830_n1814# sky130_fd_pr__pfet_01v8 ad=0.69795 pd=4.56 as=0.69795 ps=4.56 w=4.23 l=3.72
X9 B.t11 B.t9 B.t10 w_n5830_n1814# sky130_fd_pr__pfet_01v8 ad=1.6497 pd=9.24 as=0 ps=0 w=4.23 l=3.72
X10 B.t8 B.t6 B.t7 w_n5830_n1814# sky130_fd_pr__pfet_01v8 ad=1.6497 pd=9.24 as=0 ps=0 w=4.23 l=3.72
X11 B.t5 B.t3 B.t4 w_n5830_n1814# sky130_fd_pr__pfet_01v8 ad=1.6497 pd=9.24 as=0 ps=0 w=4.23 l=3.72
X12 VDD2.t4 VN.t5 VTAIL.t12 w_n5830_n1814# sky130_fd_pr__pfet_01v8 ad=0.69795 pd=4.56 as=1.6497 ps=9.24 w=4.23 l=3.72
X13 VDD2.t3 VN.t6 VTAIL.t10 w_n5830_n1814# sky130_fd_pr__pfet_01v8 ad=1.6497 pd=9.24 as=0.69795 ps=4.56 w=4.23 l=3.72
X14 VDD1.t5 VP.t4 VTAIL.t19 w_n5830_n1814# sky130_fd_pr__pfet_01v8 ad=0.69795 pd=4.56 as=1.6497 ps=9.24 w=4.23 l=3.72
X15 VTAIL.t4 VP.t5 VDD1.t4 w_n5830_n1814# sky130_fd_pr__pfet_01v8 ad=0.69795 pd=4.56 as=0.69795 ps=4.56 w=4.23 l=3.72
X16 VDD1.t3 VP.t6 VTAIL.t6 w_n5830_n1814# sky130_fd_pr__pfet_01v8 ad=0.69795 pd=4.56 as=0.69795 ps=4.56 w=4.23 l=3.72
X17 VTAIL.t3 VP.t7 VDD1.t2 w_n5830_n1814# sky130_fd_pr__pfet_01v8 ad=0.69795 pd=4.56 as=0.69795 ps=4.56 w=4.23 l=3.72
X18 VDD1.t1 VP.t8 VTAIL.t2 w_n5830_n1814# sky130_fd_pr__pfet_01v8 ad=0.69795 pd=4.56 as=1.6497 ps=9.24 w=4.23 l=3.72
X19 VTAIL.t13 VN.t7 VDD2.t2 w_n5830_n1814# sky130_fd_pr__pfet_01v8 ad=0.69795 pd=4.56 as=0.69795 ps=4.56 w=4.23 l=3.72
X20 B.t2 B.t0 B.t1 w_n5830_n1814# sky130_fd_pr__pfet_01v8 ad=1.6497 pd=9.24 as=0 ps=0 w=4.23 l=3.72
X21 VDD1.t0 VP.t9 VTAIL.t0 w_n5830_n1814# sky130_fd_pr__pfet_01v8 ad=1.6497 pd=9.24 as=0.69795 ps=4.56 w=4.23 l=3.72
X22 VTAIL.t14 VN.t8 VDD2.t1 w_n5830_n1814# sky130_fd_pr__pfet_01v8 ad=0.69795 pd=4.56 as=0.69795 ps=4.56 w=4.23 l=3.72
X23 VDD2.t0 VN.t9 VTAIL.t8 w_n5830_n1814# sky130_fd_pr__pfet_01v8 ad=1.6497 pd=9.24 as=0.69795 ps=4.56 w=4.23 l=3.72
R0 VN.n108 VN.n107 161.3
R1 VN.n106 VN.n56 161.3
R2 VN.n105 VN.n104 161.3
R3 VN.n103 VN.n57 161.3
R4 VN.n102 VN.n101 161.3
R5 VN.n100 VN.n58 161.3
R6 VN.n99 VN.n98 161.3
R7 VN.n97 VN.n59 161.3
R8 VN.n96 VN.n95 161.3
R9 VN.n94 VN.n60 161.3
R10 VN.n93 VN.n92 161.3
R11 VN.n91 VN.n62 161.3
R12 VN.n90 VN.n89 161.3
R13 VN.n88 VN.n63 161.3
R14 VN.n87 VN.n86 161.3
R15 VN.n85 VN.n64 161.3
R16 VN.n84 VN.n83 161.3
R17 VN.n82 VN.n65 161.3
R18 VN.n81 VN.n80 161.3
R19 VN.n79 VN.n66 161.3
R20 VN.n78 VN.n77 161.3
R21 VN.n76 VN.n67 161.3
R22 VN.n75 VN.n74 161.3
R23 VN.n73 VN.n68 161.3
R24 VN.n72 VN.n71 161.3
R25 VN.n53 VN.n52 161.3
R26 VN.n51 VN.n1 161.3
R27 VN.n50 VN.n49 161.3
R28 VN.n48 VN.n2 161.3
R29 VN.n47 VN.n46 161.3
R30 VN.n45 VN.n3 161.3
R31 VN.n44 VN.n43 161.3
R32 VN.n42 VN.n4 161.3
R33 VN.n41 VN.n40 161.3
R34 VN.n38 VN.n5 161.3
R35 VN.n37 VN.n36 161.3
R36 VN.n35 VN.n6 161.3
R37 VN.n34 VN.n33 161.3
R38 VN.n32 VN.n7 161.3
R39 VN.n31 VN.n30 161.3
R40 VN.n29 VN.n8 161.3
R41 VN.n28 VN.n27 161.3
R42 VN.n26 VN.n9 161.3
R43 VN.n25 VN.n24 161.3
R44 VN.n23 VN.n10 161.3
R45 VN.n22 VN.n21 161.3
R46 VN.n20 VN.n11 161.3
R47 VN.n19 VN.n18 161.3
R48 VN.n17 VN.n12 161.3
R49 VN.n16 VN.n15 161.3
R50 VN.n54 VN.n0 85.174
R51 VN.n109 VN.n55 85.174
R52 VN.n14 VN.n13 72.4354
R53 VN.n70 VN.n69 72.4354
R54 VN.n69 VN.t5 59.772
R55 VN.n13 VN.t9 59.772
R56 VN VN.n109 53.5473
R57 VN.n46 VN.n2 47.7779
R58 VN.n101 VN.n57 47.7779
R59 VN.n21 VN.n20 42.9216
R60 VN.n33 VN.n6 42.9216
R61 VN.n77 VN.n76 42.9216
R62 VN.n89 VN.n62 42.9216
R63 VN.n21 VN.n10 38.0652
R64 VN.n33 VN.n32 38.0652
R65 VN.n77 VN.n66 38.0652
R66 VN.n89 VN.n88 38.0652
R67 VN.n46 VN.n45 33.2089
R68 VN.n101 VN.n100 33.2089
R69 VN.n27 VN.t2 27.4045
R70 VN.n14 VN.t8 27.4045
R71 VN.n39 VN.t1 27.4045
R72 VN.n0 VN.t0 27.4045
R73 VN.n83 VN.t3 27.4045
R74 VN.n70 VN.t7 27.4045
R75 VN.n61 VN.t4 27.4045
R76 VN.n55 VN.t6 27.4045
R77 VN.n15 VN.n12 24.4675
R78 VN.n19 VN.n12 24.4675
R79 VN.n20 VN.n19 24.4675
R80 VN.n25 VN.n10 24.4675
R81 VN.n26 VN.n25 24.4675
R82 VN.n27 VN.n26 24.4675
R83 VN.n27 VN.n8 24.4675
R84 VN.n31 VN.n8 24.4675
R85 VN.n32 VN.n31 24.4675
R86 VN.n37 VN.n6 24.4675
R87 VN.n38 VN.n37 24.4675
R88 VN.n40 VN.n38 24.4675
R89 VN.n44 VN.n4 24.4675
R90 VN.n45 VN.n44 24.4675
R91 VN.n50 VN.n2 24.4675
R92 VN.n51 VN.n50 24.4675
R93 VN.n52 VN.n51 24.4675
R94 VN.n76 VN.n75 24.4675
R95 VN.n75 VN.n68 24.4675
R96 VN.n71 VN.n68 24.4675
R97 VN.n88 VN.n87 24.4675
R98 VN.n87 VN.n64 24.4675
R99 VN.n83 VN.n64 24.4675
R100 VN.n83 VN.n82 24.4675
R101 VN.n82 VN.n81 24.4675
R102 VN.n81 VN.n66 24.4675
R103 VN.n100 VN.n99 24.4675
R104 VN.n99 VN.n59 24.4675
R105 VN.n95 VN.n94 24.4675
R106 VN.n94 VN.n93 24.4675
R107 VN.n93 VN.n62 24.4675
R108 VN.n107 VN.n106 24.4675
R109 VN.n106 VN.n105 24.4675
R110 VN.n105 VN.n57 24.4675
R111 VN.n39 VN.n4 22.0208
R112 VN.n61 VN.n59 22.0208
R113 VN.n52 VN.n0 4.8939
R114 VN.n107 VN.n55 4.8939
R115 VN.n72 VN.n69 3.31409
R116 VN.n16 VN.n13 3.31409
R117 VN.n15 VN.n14 2.4472
R118 VN.n40 VN.n39 2.4472
R119 VN.n71 VN.n70 2.4472
R120 VN.n95 VN.n61 2.4472
R121 VN.n109 VN.n108 0.354971
R122 VN.n54 VN.n53 0.354971
R123 VN VN.n54 0.26696
R124 VN.n108 VN.n56 0.189894
R125 VN.n104 VN.n56 0.189894
R126 VN.n104 VN.n103 0.189894
R127 VN.n103 VN.n102 0.189894
R128 VN.n102 VN.n58 0.189894
R129 VN.n98 VN.n58 0.189894
R130 VN.n98 VN.n97 0.189894
R131 VN.n97 VN.n96 0.189894
R132 VN.n96 VN.n60 0.189894
R133 VN.n92 VN.n60 0.189894
R134 VN.n92 VN.n91 0.189894
R135 VN.n91 VN.n90 0.189894
R136 VN.n90 VN.n63 0.189894
R137 VN.n86 VN.n63 0.189894
R138 VN.n86 VN.n85 0.189894
R139 VN.n85 VN.n84 0.189894
R140 VN.n84 VN.n65 0.189894
R141 VN.n80 VN.n65 0.189894
R142 VN.n80 VN.n79 0.189894
R143 VN.n79 VN.n78 0.189894
R144 VN.n78 VN.n67 0.189894
R145 VN.n74 VN.n67 0.189894
R146 VN.n74 VN.n73 0.189894
R147 VN.n73 VN.n72 0.189894
R148 VN.n17 VN.n16 0.189894
R149 VN.n18 VN.n17 0.189894
R150 VN.n18 VN.n11 0.189894
R151 VN.n22 VN.n11 0.189894
R152 VN.n23 VN.n22 0.189894
R153 VN.n24 VN.n23 0.189894
R154 VN.n24 VN.n9 0.189894
R155 VN.n28 VN.n9 0.189894
R156 VN.n29 VN.n28 0.189894
R157 VN.n30 VN.n29 0.189894
R158 VN.n30 VN.n7 0.189894
R159 VN.n34 VN.n7 0.189894
R160 VN.n35 VN.n34 0.189894
R161 VN.n36 VN.n35 0.189894
R162 VN.n36 VN.n5 0.189894
R163 VN.n41 VN.n5 0.189894
R164 VN.n42 VN.n41 0.189894
R165 VN.n43 VN.n42 0.189894
R166 VN.n43 VN.n3 0.189894
R167 VN.n47 VN.n3 0.189894
R168 VN.n48 VN.n47 0.189894
R169 VN.n49 VN.n48 0.189894
R170 VN.n49 VN.n1 0.189894
R171 VN.n53 VN.n1 0.189894
R172 VTAIL.n11 VTAIL.t12 99.9741
R173 VTAIL.n17 VTAIL.t17 99.9738
R174 VTAIL.n2 VTAIL.t19 99.9738
R175 VTAIL.n16 VTAIL.t2 99.9738
R176 VTAIL.n15 VTAIL.n14 92.2897
R177 VTAIL.n13 VTAIL.n12 92.2897
R178 VTAIL.n10 VTAIL.n9 92.2897
R179 VTAIL.n8 VTAIL.n7 92.2897
R180 VTAIL.n19 VTAIL.n18 92.2894
R181 VTAIL.n1 VTAIL.n0 92.2894
R182 VTAIL.n4 VTAIL.n3 92.2894
R183 VTAIL.n6 VTAIL.n5 92.2894
R184 VTAIL.n8 VTAIL.n6 22.9962
R185 VTAIL.n17 VTAIL.n16 19.5048
R186 VTAIL.n18 VTAIL.t15 7.6849
R187 VTAIL.n18 VTAIL.t11 7.6849
R188 VTAIL.n0 VTAIL.t8 7.6849
R189 VTAIL.n0 VTAIL.t14 7.6849
R190 VTAIL.n3 VTAIL.t1 7.6849
R191 VTAIL.n3 VTAIL.t4 7.6849
R192 VTAIL.n5 VTAIL.t5 7.6849
R193 VTAIL.n5 VTAIL.t7 7.6849
R194 VTAIL.n14 VTAIL.t6 7.6849
R195 VTAIL.n14 VTAIL.t3 7.6849
R196 VTAIL.n12 VTAIL.t0 7.6849
R197 VTAIL.n12 VTAIL.t18 7.6849
R198 VTAIL.n9 VTAIL.t16 7.6849
R199 VTAIL.n9 VTAIL.t13 7.6849
R200 VTAIL.n7 VTAIL.t10 7.6849
R201 VTAIL.n7 VTAIL.t9 7.6849
R202 VTAIL.n10 VTAIL.n8 3.49188
R203 VTAIL.n11 VTAIL.n10 3.49188
R204 VTAIL.n15 VTAIL.n13 3.49188
R205 VTAIL.n16 VTAIL.n15 3.49188
R206 VTAIL.n6 VTAIL.n4 3.49188
R207 VTAIL.n4 VTAIL.n2 3.49188
R208 VTAIL.n19 VTAIL.n17 3.49188
R209 VTAIL VTAIL.n1 2.67722
R210 VTAIL.n13 VTAIL.n11 2.21602
R211 VTAIL.n2 VTAIL.n1 2.21602
R212 VTAIL VTAIL.n19 0.815155
R213 VDD2.n1 VDD2.t0 120.144
R214 VDD2.n4 VDD2.t3 116.653
R215 VDD2.n3 VDD2.n2 111.531
R216 VDD2 VDD2.n7 111.528
R217 VDD2.n6 VDD2.n5 108.969
R218 VDD2.n1 VDD2.n0 108.969
R219 VDD2.n4 VDD2.n3 43.9459
R220 VDD2.n7 VDD2.t2 7.6849
R221 VDD2.n7 VDD2.t4 7.6849
R222 VDD2.n5 VDD2.t5 7.6849
R223 VDD2.n5 VDD2.t6 7.6849
R224 VDD2.n2 VDD2.t8 7.6849
R225 VDD2.n2 VDD2.t9 7.6849
R226 VDD2.n0 VDD2.t1 7.6849
R227 VDD2.n0 VDD2.t7 7.6849
R228 VDD2.n6 VDD2.n4 3.49188
R229 VDD2 VDD2.n6 0.931535
R230 VDD2.n3 VDD2.n1 0.817999
R231 VP.n33 VP.n32 161.3
R232 VP.n34 VP.n29 161.3
R233 VP.n36 VP.n35 161.3
R234 VP.n37 VP.n28 161.3
R235 VP.n39 VP.n38 161.3
R236 VP.n40 VP.n27 161.3
R237 VP.n42 VP.n41 161.3
R238 VP.n43 VP.n26 161.3
R239 VP.n45 VP.n44 161.3
R240 VP.n46 VP.n25 161.3
R241 VP.n48 VP.n47 161.3
R242 VP.n49 VP.n24 161.3
R243 VP.n51 VP.n50 161.3
R244 VP.n52 VP.n23 161.3
R245 VP.n54 VP.n53 161.3
R246 VP.n55 VP.n22 161.3
R247 VP.n58 VP.n57 161.3
R248 VP.n59 VP.n21 161.3
R249 VP.n61 VP.n60 161.3
R250 VP.n62 VP.n20 161.3
R251 VP.n64 VP.n63 161.3
R252 VP.n65 VP.n19 161.3
R253 VP.n67 VP.n66 161.3
R254 VP.n68 VP.n18 161.3
R255 VP.n70 VP.n69 161.3
R256 VP.n125 VP.n124 161.3
R257 VP.n123 VP.n1 161.3
R258 VP.n122 VP.n121 161.3
R259 VP.n120 VP.n2 161.3
R260 VP.n119 VP.n118 161.3
R261 VP.n117 VP.n3 161.3
R262 VP.n116 VP.n115 161.3
R263 VP.n114 VP.n4 161.3
R264 VP.n113 VP.n112 161.3
R265 VP.n110 VP.n5 161.3
R266 VP.n109 VP.n108 161.3
R267 VP.n107 VP.n6 161.3
R268 VP.n106 VP.n105 161.3
R269 VP.n104 VP.n7 161.3
R270 VP.n103 VP.n102 161.3
R271 VP.n101 VP.n8 161.3
R272 VP.n100 VP.n99 161.3
R273 VP.n98 VP.n9 161.3
R274 VP.n97 VP.n96 161.3
R275 VP.n95 VP.n10 161.3
R276 VP.n94 VP.n93 161.3
R277 VP.n92 VP.n11 161.3
R278 VP.n91 VP.n90 161.3
R279 VP.n89 VP.n12 161.3
R280 VP.n88 VP.n87 161.3
R281 VP.n85 VP.n13 161.3
R282 VP.n84 VP.n83 161.3
R283 VP.n82 VP.n14 161.3
R284 VP.n81 VP.n80 161.3
R285 VP.n79 VP.n15 161.3
R286 VP.n78 VP.n77 161.3
R287 VP.n76 VP.n16 161.3
R288 VP.n75 VP.n74 161.3
R289 VP.n73 VP.n72 85.174
R290 VP.n126 VP.n0 85.174
R291 VP.n71 VP.n17 85.174
R292 VP.n31 VP.n30 72.4355
R293 VP.n30 VP.t9 59.7719
R294 VP.n72 VP.n71 53.3819
R295 VP.n80 VP.n79 47.7779
R296 VP.n118 VP.n2 47.7779
R297 VP.n63 VP.n19 47.7779
R298 VP.n93 VP.n92 42.9216
R299 VP.n105 VP.n6 42.9216
R300 VP.n50 VP.n23 42.9216
R301 VP.n38 VP.n37 42.9216
R302 VP.n93 VP.n10 38.0652
R303 VP.n105 VP.n104 38.0652
R304 VP.n50 VP.n49 38.0652
R305 VP.n38 VP.n27 38.0652
R306 VP.n80 VP.n14 33.2089
R307 VP.n118 VP.n117 33.2089
R308 VP.n63 VP.n62 33.2089
R309 VP.n99 VP.t3 27.4045
R310 VP.n73 VP.t0 27.4045
R311 VP.n86 VP.t2 27.4045
R312 VP.n111 VP.t5 27.4045
R313 VP.n0 VP.t4 27.4045
R314 VP.n44 VP.t6 27.4045
R315 VP.n17 VP.t8 27.4045
R316 VP.n56 VP.t7 27.4045
R317 VP.n31 VP.t1 27.4045
R318 VP.n74 VP.n16 24.4675
R319 VP.n78 VP.n16 24.4675
R320 VP.n79 VP.n78 24.4675
R321 VP.n84 VP.n14 24.4675
R322 VP.n85 VP.n84 24.4675
R323 VP.n87 VP.n12 24.4675
R324 VP.n91 VP.n12 24.4675
R325 VP.n92 VP.n91 24.4675
R326 VP.n97 VP.n10 24.4675
R327 VP.n98 VP.n97 24.4675
R328 VP.n99 VP.n98 24.4675
R329 VP.n99 VP.n8 24.4675
R330 VP.n103 VP.n8 24.4675
R331 VP.n104 VP.n103 24.4675
R332 VP.n109 VP.n6 24.4675
R333 VP.n110 VP.n109 24.4675
R334 VP.n112 VP.n110 24.4675
R335 VP.n116 VP.n4 24.4675
R336 VP.n117 VP.n116 24.4675
R337 VP.n122 VP.n2 24.4675
R338 VP.n123 VP.n122 24.4675
R339 VP.n124 VP.n123 24.4675
R340 VP.n67 VP.n19 24.4675
R341 VP.n68 VP.n67 24.4675
R342 VP.n69 VP.n68 24.4675
R343 VP.n54 VP.n23 24.4675
R344 VP.n55 VP.n54 24.4675
R345 VP.n57 VP.n55 24.4675
R346 VP.n61 VP.n21 24.4675
R347 VP.n62 VP.n61 24.4675
R348 VP.n42 VP.n27 24.4675
R349 VP.n43 VP.n42 24.4675
R350 VP.n44 VP.n43 24.4675
R351 VP.n44 VP.n25 24.4675
R352 VP.n48 VP.n25 24.4675
R353 VP.n49 VP.n48 24.4675
R354 VP.n32 VP.n29 24.4675
R355 VP.n36 VP.n29 24.4675
R356 VP.n37 VP.n36 24.4675
R357 VP.n86 VP.n85 22.0208
R358 VP.n111 VP.n4 22.0208
R359 VP.n56 VP.n21 22.0208
R360 VP.n74 VP.n73 4.8939
R361 VP.n124 VP.n0 4.8939
R362 VP.n69 VP.n17 4.8939
R363 VP.n33 VP.n30 3.31408
R364 VP.n87 VP.n86 2.4472
R365 VP.n112 VP.n111 2.4472
R366 VP.n57 VP.n56 2.4472
R367 VP.n32 VP.n31 2.4472
R368 VP.n71 VP.n70 0.354971
R369 VP.n75 VP.n72 0.354971
R370 VP.n126 VP.n125 0.354971
R371 VP VP.n126 0.26696
R372 VP.n34 VP.n33 0.189894
R373 VP.n35 VP.n34 0.189894
R374 VP.n35 VP.n28 0.189894
R375 VP.n39 VP.n28 0.189894
R376 VP.n40 VP.n39 0.189894
R377 VP.n41 VP.n40 0.189894
R378 VP.n41 VP.n26 0.189894
R379 VP.n45 VP.n26 0.189894
R380 VP.n46 VP.n45 0.189894
R381 VP.n47 VP.n46 0.189894
R382 VP.n47 VP.n24 0.189894
R383 VP.n51 VP.n24 0.189894
R384 VP.n52 VP.n51 0.189894
R385 VP.n53 VP.n52 0.189894
R386 VP.n53 VP.n22 0.189894
R387 VP.n58 VP.n22 0.189894
R388 VP.n59 VP.n58 0.189894
R389 VP.n60 VP.n59 0.189894
R390 VP.n60 VP.n20 0.189894
R391 VP.n64 VP.n20 0.189894
R392 VP.n65 VP.n64 0.189894
R393 VP.n66 VP.n65 0.189894
R394 VP.n66 VP.n18 0.189894
R395 VP.n70 VP.n18 0.189894
R396 VP.n76 VP.n75 0.189894
R397 VP.n77 VP.n76 0.189894
R398 VP.n77 VP.n15 0.189894
R399 VP.n81 VP.n15 0.189894
R400 VP.n82 VP.n81 0.189894
R401 VP.n83 VP.n82 0.189894
R402 VP.n83 VP.n13 0.189894
R403 VP.n88 VP.n13 0.189894
R404 VP.n89 VP.n88 0.189894
R405 VP.n90 VP.n89 0.189894
R406 VP.n90 VP.n11 0.189894
R407 VP.n94 VP.n11 0.189894
R408 VP.n95 VP.n94 0.189894
R409 VP.n96 VP.n95 0.189894
R410 VP.n96 VP.n9 0.189894
R411 VP.n100 VP.n9 0.189894
R412 VP.n101 VP.n100 0.189894
R413 VP.n102 VP.n101 0.189894
R414 VP.n102 VP.n7 0.189894
R415 VP.n106 VP.n7 0.189894
R416 VP.n107 VP.n106 0.189894
R417 VP.n108 VP.n107 0.189894
R418 VP.n108 VP.n5 0.189894
R419 VP.n113 VP.n5 0.189894
R420 VP.n114 VP.n113 0.189894
R421 VP.n115 VP.n114 0.189894
R422 VP.n115 VP.n3 0.189894
R423 VP.n119 VP.n3 0.189894
R424 VP.n120 VP.n119 0.189894
R425 VP.n121 VP.n120 0.189894
R426 VP.n121 VP.n1 0.189894
R427 VP.n125 VP.n1 0.189894
R428 VDD1.n1 VDD1.t0 120.144
R429 VDD1.n3 VDD1.t9 120.144
R430 VDD1.n5 VDD1.n4 111.531
R431 VDD1.n1 VDD1.n0 108.969
R432 VDD1.n7 VDD1.n6 108.969
R433 VDD1.n3 VDD1.n2 108.969
R434 VDD1.n7 VDD1.n5 46.2746
R435 VDD1.n6 VDD1.t2 7.6849
R436 VDD1.n6 VDD1.t1 7.6849
R437 VDD1.n0 VDD1.t8 7.6849
R438 VDD1.n0 VDD1.t3 7.6849
R439 VDD1.n4 VDD1.t4 7.6849
R440 VDD1.n4 VDD1.t5 7.6849
R441 VDD1.n2 VDD1.t7 7.6849
R442 VDD1.n2 VDD1.t6 7.6849
R443 VDD1 VDD1.n7 2.56084
R444 VDD1 VDD1.n1 0.931535
R445 VDD1.n5 VDD1.n3 0.817999
R446 B.n404 B.n149 585
R447 B.n403 B.n402 585
R448 B.n401 B.n150 585
R449 B.n400 B.n399 585
R450 B.n398 B.n151 585
R451 B.n397 B.n396 585
R452 B.n395 B.n152 585
R453 B.n394 B.n393 585
R454 B.n392 B.n153 585
R455 B.n391 B.n390 585
R456 B.n389 B.n154 585
R457 B.n388 B.n387 585
R458 B.n386 B.n155 585
R459 B.n385 B.n384 585
R460 B.n383 B.n156 585
R461 B.n382 B.n381 585
R462 B.n380 B.n157 585
R463 B.n379 B.n378 585
R464 B.n377 B.n158 585
R465 B.n376 B.n375 585
R466 B.n371 B.n159 585
R467 B.n370 B.n369 585
R468 B.n368 B.n160 585
R469 B.n367 B.n366 585
R470 B.n365 B.n161 585
R471 B.n364 B.n363 585
R472 B.n362 B.n162 585
R473 B.n361 B.n360 585
R474 B.n358 B.n163 585
R475 B.n357 B.n356 585
R476 B.n355 B.n166 585
R477 B.n354 B.n353 585
R478 B.n352 B.n167 585
R479 B.n351 B.n350 585
R480 B.n349 B.n168 585
R481 B.n348 B.n347 585
R482 B.n346 B.n169 585
R483 B.n345 B.n344 585
R484 B.n343 B.n170 585
R485 B.n342 B.n341 585
R486 B.n340 B.n171 585
R487 B.n339 B.n338 585
R488 B.n337 B.n172 585
R489 B.n336 B.n335 585
R490 B.n334 B.n173 585
R491 B.n333 B.n332 585
R492 B.n331 B.n174 585
R493 B.n406 B.n405 585
R494 B.n407 B.n148 585
R495 B.n409 B.n408 585
R496 B.n410 B.n147 585
R497 B.n412 B.n411 585
R498 B.n413 B.n146 585
R499 B.n415 B.n414 585
R500 B.n416 B.n145 585
R501 B.n418 B.n417 585
R502 B.n419 B.n144 585
R503 B.n421 B.n420 585
R504 B.n422 B.n143 585
R505 B.n424 B.n423 585
R506 B.n425 B.n142 585
R507 B.n427 B.n426 585
R508 B.n428 B.n141 585
R509 B.n430 B.n429 585
R510 B.n431 B.n140 585
R511 B.n433 B.n432 585
R512 B.n434 B.n139 585
R513 B.n436 B.n435 585
R514 B.n437 B.n138 585
R515 B.n439 B.n438 585
R516 B.n440 B.n137 585
R517 B.n442 B.n441 585
R518 B.n443 B.n136 585
R519 B.n445 B.n444 585
R520 B.n446 B.n135 585
R521 B.n448 B.n447 585
R522 B.n449 B.n134 585
R523 B.n451 B.n450 585
R524 B.n452 B.n133 585
R525 B.n454 B.n453 585
R526 B.n455 B.n132 585
R527 B.n457 B.n456 585
R528 B.n458 B.n131 585
R529 B.n460 B.n459 585
R530 B.n461 B.n130 585
R531 B.n463 B.n462 585
R532 B.n464 B.n129 585
R533 B.n466 B.n465 585
R534 B.n467 B.n128 585
R535 B.n469 B.n468 585
R536 B.n470 B.n127 585
R537 B.n472 B.n471 585
R538 B.n473 B.n126 585
R539 B.n475 B.n474 585
R540 B.n476 B.n125 585
R541 B.n478 B.n477 585
R542 B.n479 B.n124 585
R543 B.n481 B.n480 585
R544 B.n482 B.n123 585
R545 B.n484 B.n483 585
R546 B.n485 B.n122 585
R547 B.n487 B.n486 585
R548 B.n488 B.n121 585
R549 B.n490 B.n489 585
R550 B.n491 B.n120 585
R551 B.n493 B.n492 585
R552 B.n494 B.n119 585
R553 B.n496 B.n495 585
R554 B.n497 B.n118 585
R555 B.n499 B.n498 585
R556 B.n500 B.n117 585
R557 B.n502 B.n501 585
R558 B.n503 B.n116 585
R559 B.n505 B.n504 585
R560 B.n506 B.n115 585
R561 B.n508 B.n507 585
R562 B.n509 B.n114 585
R563 B.n511 B.n510 585
R564 B.n512 B.n113 585
R565 B.n514 B.n513 585
R566 B.n515 B.n112 585
R567 B.n517 B.n516 585
R568 B.n518 B.n111 585
R569 B.n520 B.n519 585
R570 B.n521 B.n110 585
R571 B.n523 B.n522 585
R572 B.n524 B.n109 585
R573 B.n526 B.n525 585
R574 B.n527 B.n108 585
R575 B.n529 B.n528 585
R576 B.n530 B.n107 585
R577 B.n532 B.n531 585
R578 B.n533 B.n106 585
R579 B.n535 B.n534 585
R580 B.n536 B.n105 585
R581 B.n538 B.n537 585
R582 B.n539 B.n104 585
R583 B.n541 B.n540 585
R584 B.n542 B.n103 585
R585 B.n544 B.n543 585
R586 B.n545 B.n102 585
R587 B.n547 B.n546 585
R588 B.n548 B.n101 585
R589 B.n550 B.n549 585
R590 B.n551 B.n100 585
R591 B.n553 B.n552 585
R592 B.n554 B.n99 585
R593 B.n556 B.n555 585
R594 B.n557 B.n98 585
R595 B.n559 B.n558 585
R596 B.n560 B.n97 585
R597 B.n562 B.n561 585
R598 B.n563 B.n96 585
R599 B.n565 B.n564 585
R600 B.n566 B.n95 585
R601 B.n568 B.n567 585
R602 B.n569 B.n94 585
R603 B.n571 B.n570 585
R604 B.n572 B.n93 585
R605 B.n574 B.n573 585
R606 B.n575 B.n92 585
R607 B.n577 B.n576 585
R608 B.n578 B.n91 585
R609 B.n580 B.n579 585
R610 B.n581 B.n90 585
R611 B.n583 B.n582 585
R612 B.n584 B.n89 585
R613 B.n586 B.n585 585
R614 B.n587 B.n88 585
R615 B.n589 B.n588 585
R616 B.n590 B.n87 585
R617 B.n592 B.n591 585
R618 B.n593 B.n86 585
R619 B.n595 B.n594 585
R620 B.n596 B.n85 585
R621 B.n598 B.n597 585
R622 B.n599 B.n84 585
R623 B.n601 B.n600 585
R624 B.n602 B.n83 585
R625 B.n604 B.n603 585
R626 B.n605 B.n82 585
R627 B.n607 B.n606 585
R628 B.n608 B.n81 585
R629 B.n610 B.n609 585
R630 B.n611 B.n80 585
R631 B.n613 B.n612 585
R632 B.n614 B.n79 585
R633 B.n616 B.n615 585
R634 B.n617 B.n78 585
R635 B.n619 B.n618 585
R636 B.n620 B.n77 585
R637 B.n622 B.n621 585
R638 B.n623 B.n76 585
R639 B.n625 B.n624 585
R640 B.n626 B.n75 585
R641 B.n628 B.n627 585
R642 B.n629 B.n74 585
R643 B.n631 B.n630 585
R644 B.n632 B.n73 585
R645 B.n634 B.n633 585
R646 B.n635 B.n72 585
R647 B.n637 B.n636 585
R648 B.n638 B.n71 585
R649 B.n640 B.n639 585
R650 B.n641 B.n70 585
R651 B.n643 B.n642 585
R652 B.n644 B.n69 585
R653 B.n717 B.n716 585
R654 B.n715 B.n42 585
R655 B.n714 B.n713 585
R656 B.n712 B.n43 585
R657 B.n711 B.n710 585
R658 B.n709 B.n44 585
R659 B.n708 B.n707 585
R660 B.n706 B.n45 585
R661 B.n705 B.n704 585
R662 B.n703 B.n46 585
R663 B.n702 B.n701 585
R664 B.n700 B.n47 585
R665 B.n699 B.n698 585
R666 B.n697 B.n48 585
R667 B.n696 B.n695 585
R668 B.n694 B.n49 585
R669 B.n693 B.n692 585
R670 B.n691 B.n50 585
R671 B.n690 B.n689 585
R672 B.n687 B.n51 585
R673 B.n686 B.n685 585
R674 B.n684 B.n54 585
R675 B.n683 B.n682 585
R676 B.n681 B.n55 585
R677 B.n680 B.n679 585
R678 B.n678 B.n56 585
R679 B.n677 B.n676 585
R680 B.n675 B.n57 585
R681 B.n673 B.n672 585
R682 B.n671 B.n60 585
R683 B.n670 B.n669 585
R684 B.n668 B.n61 585
R685 B.n667 B.n666 585
R686 B.n665 B.n62 585
R687 B.n664 B.n663 585
R688 B.n662 B.n63 585
R689 B.n661 B.n660 585
R690 B.n659 B.n64 585
R691 B.n658 B.n657 585
R692 B.n656 B.n65 585
R693 B.n655 B.n654 585
R694 B.n653 B.n66 585
R695 B.n652 B.n651 585
R696 B.n650 B.n67 585
R697 B.n649 B.n648 585
R698 B.n647 B.n68 585
R699 B.n646 B.n645 585
R700 B.n718 B.n41 585
R701 B.n720 B.n719 585
R702 B.n721 B.n40 585
R703 B.n723 B.n722 585
R704 B.n724 B.n39 585
R705 B.n726 B.n725 585
R706 B.n727 B.n38 585
R707 B.n729 B.n728 585
R708 B.n730 B.n37 585
R709 B.n732 B.n731 585
R710 B.n733 B.n36 585
R711 B.n735 B.n734 585
R712 B.n736 B.n35 585
R713 B.n738 B.n737 585
R714 B.n739 B.n34 585
R715 B.n741 B.n740 585
R716 B.n742 B.n33 585
R717 B.n744 B.n743 585
R718 B.n745 B.n32 585
R719 B.n747 B.n746 585
R720 B.n748 B.n31 585
R721 B.n750 B.n749 585
R722 B.n751 B.n30 585
R723 B.n753 B.n752 585
R724 B.n754 B.n29 585
R725 B.n756 B.n755 585
R726 B.n757 B.n28 585
R727 B.n759 B.n758 585
R728 B.n760 B.n27 585
R729 B.n762 B.n761 585
R730 B.n763 B.n26 585
R731 B.n765 B.n764 585
R732 B.n766 B.n25 585
R733 B.n768 B.n767 585
R734 B.n769 B.n24 585
R735 B.n771 B.n770 585
R736 B.n772 B.n23 585
R737 B.n774 B.n773 585
R738 B.n775 B.n22 585
R739 B.n777 B.n776 585
R740 B.n778 B.n21 585
R741 B.n780 B.n779 585
R742 B.n781 B.n20 585
R743 B.n783 B.n782 585
R744 B.n784 B.n19 585
R745 B.n786 B.n785 585
R746 B.n787 B.n18 585
R747 B.n789 B.n788 585
R748 B.n790 B.n17 585
R749 B.n792 B.n791 585
R750 B.n793 B.n16 585
R751 B.n795 B.n794 585
R752 B.n796 B.n15 585
R753 B.n798 B.n797 585
R754 B.n799 B.n14 585
R755 B.n801 B.n800 585
R756 B.n802 B.n13 585
R757 B.n804 B.n803 585
R758 B.n805 B.n12 585
R759 B.n807 B.n806 585
R760 B.n808 B.n11 585
R761 B.n810 B.n809 585
R762 B.n811 B.n10 585
R763 B.n813 B.n812 585
R764 B.n814 B.n9 585
R765 B.n816 B.n815 585
R766 B.n817 B.n8 585
R767 B.n819 B.n818 585
R768 B.n820 B.n7 585
R769 B.n822 B.n821 585
R770 B.n823 B.n6 585
R771 B.n825 B.n824 585
R772 B.n826 B.n5 585
R773 B.n828 B.n827 585
R774 B.n829 B.n4 585
R775 B.n831 B.n830 585
R776 B.n832 B.n3 585
R777 B.n834 B.n833 585
R778 B.n835 B.n0 585
R779 B.n2 B.n1 585
R780 B.n214 B.n213 585
R781 B.n216 B.n215 585
R782 B.n217 B.n212 585
R783 B.n219 B.n218 585
R784 B.n220 B.n211 585
R785 B.n222 B.n221 585
R786 B.n223 B.n210 585
R787 B.n225 B.n224 585
R788 B.n226 B.n209 585
R789 B.n228 B.n227 585
R790 B.n229 B.n208 585
R791 B.n231 B.n230 585
R792 B.n232 B.n207 585
R793 B.n234 B.n233 585
R794 B.n235 B.n206 585
R795 B.n237 B.n236 585
R796 B.n238 B.n205 585
R797 B.n240 B.n239 585
R798 B.n241 B.n204 585
R799 B.n243 B.n242 585
R800 B.n244 B.n203 585
R801 B.n246 B.n245 585
R802 B.n247 B.n202 585
R803 B.n249 B.n248 585
R804 B.n250 B.n201 585
R805 B.n252 B.n251 585
R806 B.n253 B.n200 585
R807 B.n255 B.n254 585
R808 B.n256 B.n199 585
R809 B.n258 B.n257 585
R810 B.n259 B.n198 585
R811 B.n261 B.n260 585
R812 B.n262 B.n197 585
R813 B.n264 B.n263 585
R814 B.n265 B.n196 585
R815 B.n267 B.n266 585
R816 B.n268 B.n195 585
R817 B.n270 B.n269 585
R818 B.n271 B.n194 585
R819 B.n273 B.n272 585
R820 B.n274 B.n193 585
R821 B.n276 B.n275 585
R822 B.n277 B.n192 585
R823 B.n279 B.n278 585
R824 B.n280 B.n191 585
R825 B.n282 B.n281 585
R826 B.n283 B.n190 585
R827 B.n285 B.n284 585
R828 B.n286 B.n189 585
R829 B.n288 B.n287 585
R830 B.n289 B.n188 585
R831 B.n291 B.n290 585
R832 B.n292 B.n187 585
R833 B.n294 B.n293 585
R834 B.n295 B.n186 585
R835 B.n297 B.n296 585
R836 B.n298 B.n185 585
R837 B.n300 B.n299 585
R838 B.n301 B.n184 585
R839 B.n303 B.n302 585
R840 B.n304 B.n183 585
R841 B.n306 B.n305 585
R842 B.n307 B.n182 585
R843 B.n309 B.n308 585
R844 B.n310 B.n181 585
R845 B.n312 B.n311 585
R846 B.n313 B.n180 585
R847 B.n315 B.n314 585
R848 B.n316 B.n179 585
R849 B.n318 B.n317 585
R850 B.n319 B.n178 585
R851 B.n321 B.n320 585
R852 B.n322 B.n177 585
R853 B.n324 B.n323 585
R854 B.n325 B.n176 585
R855 B.n327 B.n326 585
R856 B.n328 B.n175 585
R857 B.n330 B.n329 585
R858 B.n331 B.n330 521.33
R859 B.n406 B.n149 521.33
R860 B.n646 B.n69 521.33
R861 B.n716 B.n41 521.33
R862 B.n837 B.n836 256.663
R863 B.n164 B.t3 236.685
R864 B.n372 B.t0 236.685
R865 B.n58 B.t6 236.685
R866 B.n52 B.t9 236.685
R867 B.n836 B.n835 235.042
R868 B.n836 B.n2 235.042
R869 B.n372 B.t1 200.263
R870 B.n58 B.t8 200.263
R871 B.n164 B.t4 200.26
R872 B.n52 B.t11 200.26
R873 B.n332 B.n331 163.367
R874 B.n332 B.n173 163.367
R875 B.n336 B.n173 163.367
R876 B.n337 B.n336 163.367
R877 B.n338 B.n337 163.367
R878 B.n338 B.n171 163.367
R879 B.n342 B.n171 163.367
R880 B.n343 B.n342 163.367
R881 B.n344 B.n343 163.367
R882 B.n344 B.n169 163.367
R883 B.n348 B.n169 163.367
R884 B.n349 B.n348 163.367
R885 B.n350 B.n349 163.367
R886 B.n350 B.n167 163.367
R887 B.n354 B.n167 163.367
R888 B.n355 B.n354 163.367
R889 B.n356 B.n355 163.367
R890 B.n356 B.n163 163.367
R891 B.n361 B.n163 163.367
R892 B.n362 B.n361 163.367
R893 B.n363 B.n362 163.367
R894 B.n363 B.n161 163.367
R895 B.n367 B.n161 163.367
R896 B.n368 B.n367 163.367
R897 B.n369 B.n368 163.367
R898 B.n369 B.n159 163.367
R899 B.n376 B.n159 163.367
R900 B.n377 B.n376 163.367
R901 B.n378 B.n377 163.367
R902 B.n378 B.n157 163.367
R903 B.n382 B.n157 163.367
R904 B.n383 B.n382 163.367
R905 B.n384 B.n383 163.367
R906 B.n384 B.n155 163.367
R907 B.n388 B.n155 163.367
R908 B.n389 B.n388 163.367
R909 B.n390 B.n389 163.367
R910 B.n390 B.n153 163.367
R911 B.n394 B.n153 163.367
R912 B.n395 B.n394 163.367
R913 B.n396 B.n395 163.367
R914 B.n396 B.n151 163.367
R915 B.n400 B.n151 163.367
R916 B.n401 B.n400 163.367
R917 B.n402 B.n401 163.367
R918 B.n402 B.n149 163.367
R919 B.n642 B.n69 163.367
R920 B.n642 B.n641 163.367
R921 B.n641 B.n640 163.367
R922 B.n640 B.n71 163.367
R923 B.n636 B.n71 163.367
R924 B.n636 B.n635 163.367
R925 B.n635 B.n634 163.367
R926 B.n634 B.n73 163.367
R927 B.n630 B.n73 163.367
R928 B.n630 B.n629 163.367
R929 B.n629 B.n628 163.367
R930 B.n628 B.n75 163.367
R931 B.n624 B.n75 163.367
R932 B.n624 B.n623 163.367
R933 B.n623 B.n622 163.367
R934 B.n622 B.n77 163.367
R935 B.n618 B.n77 163.367
R936 B.n618 B.n617 163.367
R937 B.n617 B.n616 163.367
R938 B.n616 B.n79 163.367
R939 B.n612 B.n79 163.367
R940 B.n612 B.n611 163.367
R941 B.n611 B.n610 163.367
R942 B.n610 B.n81 163.367
R943 B.n606 B.n81 163.367
R944 B.n606 B.n605 163.367
R945 B.n605 B.n604 163.367
R946 B.n604 B.n83 163.367
R947 B.n600 B.n83 163.367
R948 B.n600 B.n599 163.367
R949 B.n599 B.n598 163.367
R950 B.n598 B.n85 163.367
R951 B.n594 B.n85 163.367
R952 B.n594 B.n593 163.367
R953 B.n593 B.n592 163.367
R954 B.n592 B.n87 163.367
R955 B.n588 B.n87 163.367
R956 B.n588 B.n587 163.367
R957 B.n587 B.n586 163.367
R958 B.n586 B.n89 163.367
R959 B.n582 B.n89 163.367
R960 B.n582 B.n581 163.367
R961 B.n581 B.n580 163.367
R962 B.n580 B.n91 163.367
R963 B.n576 B.n91 163.367
R964 B.n576 B.n575 163.367
R965 B.n575 B.n574 163.367
R966 B.n574 B.n93 163.367
R967 B.n570 B.n93 163.367
R968 B.n570 B.n569 163.367
R969 B.n569 B.n568 163.367
R970 B.n568 B.n95 163.367
R971 B.n564 B.n95 163.367
R972 B.n564 B.n563 163.367
R973 B.n563 B.n562 163.367
R974 B.n562 B.n97 163.367
R975 B.n558 B.n97 163.367
R976 B.n558 B.n557 163.367
R977 B.n557 B.n556 163.367
R978 B.n556 B.n99 163.367
R979 B.n552 B.n99 163.367
R980 B.n552 B.n551 163.367
R981 B.n551 B.n550 163.367
R982 B.n550 B.n101 163.367
R983 B.n546 B.n101 163.367
R984 B.n546 B.n545 163.367
R985 B.n545 B.n544 163.367
R986 B.n544 B.n103 163.367
R987 B.n540 B.n103 163.367
R988 B.n540 B.n539 163.367
R989 B.n539 B.n538 163.367
R990 B.n538 B.n105 163.367
R991 B.n534 B.n105 163.367
R992 B.n534 B.n533 163.367
R993 B.n533 B.n532 163.367
R994 B.n532 B.n107 163.367
R995 B.n528 B.n107 163.367
R996 B.n528 B.n527 163.367
R997 B.n527 B.n526 163.367
R998 B.n526 B.n109 163.367
R999 B.n522 B.n109 163.367
R1000 B.n522 B.n521 163.367
R1001 B.n521 B.n520 163.367
R1002 B.n520 B.n111 163.367
R1003 B.n516 B.n111 163.367
R1004 B.n516 B.n515 163.367
R1005 B.n515 B.n514 163.367
R1006 B.n514 B.n113 163.367
R1007 B.n510 B.n113 163.367
R1008 B.n510 B.n509 163.367
R1009 B.n509 B.n508 163.367
R1010 B.n508 B.n115 163.367
R1011 B.n504 B.n115 163.367
R1012 B.n504 B.n503 163.367
R1013 B.n503 B.n502 163.367
R1014 B.n502 B.n117 163.367
R1015 B.n498 B.n117 163.367
R1016 B.n498 B.n497 163.367
R1017 B.n497 B.n496 163.367
R1018 B.n496 B.n119 163.367
R1019 B.n492 B.n119 163.367
R1020 B.n492 B.n491 163.367
R1021 B.n491 B.n490 163.367
R1022 B.n490 B.n121 163.367
R1023 B.n486 B.n121 163.367
R1024 B.n486 B.n485 163.367
R1025 B.n485 B.n484 163.367
R1026 B.n484 B.n123 163.367
R1027 B.n480 B.n123 163.367
R1028 B.n480 B.n479 163.367
R1029 B.n479 B.n478 163.367
R1030 B.n478 B.n125 163.367
R1031 B.n474 B.n125 163.367
R1032 B.n474 B.n473 163.367
R1033 B.n473 B.n472 163.367
R1034 B.n472 B.n127 163.367
R1035 B.n468 B.n127 163.367
R1036 B.n468 B.n467 163.367
R1037 B.n467 B.n466 163.367
R1038 B.n466 B.n129 163.367
R1039 B.n462 B.n129 163.367
R1040 B.n462 B.n461 163.367
R1041 B.n461 B.n460 163.367
R1042 B.n460 B.n131 163.367
R1043 B.n456 B.n131 163.367
R1044 B.n456 B.n455 163.367
R1045 B.n455 B.n454 163.367
R1046 B.n454 B.n133 163.367
R1047 B.n450 B.n133 163.367
R1048 B.n450 B.n449 163.367
R1049 B.n449 B.n448 163.367
R1050 B.n448 B.n135 163.367
R1051 B.n444 B.n135 163.367
R1052 B.n444 B.n443 163.367
R1053 B.n443 B.n442 163.367
R1054 B.n442 B.n137 163.367
R1055 B.n438 B.n137 163.367
R1056 B.n438 B.n437 163.367
R1057 B.n437 B.n436 163.367
R1058 B.n436 B.n139 163.367
R1059 B.n432 B.n139 163.367
R1060 B.n432 B.n431 163.367
R1061 B.n431 B.n430 163.367
R1062 B.n430 B.n141 163.367
R1063 B.n426 B.n141 163.367
R1064 B.n426 B.n425 163.367
R1065 B.n425 B.n424 163.367
R1066 B.n424 B.n143 163.367
R1067 B.n420 B.n143 163.367
R1068 B.n420 B.n419 163.367
R1069 B.n419 B.n418 163.367
R1070 B.n418 B.n145 163.367
R1071 B.n414 B.n145 163.367
R1072 B.n414 B.n413 163.367
R1073 B.n413 B.n412 163.367
R1074 B.n412 B.n147 163.367
R1075 B.n408 B.n147 163.367
R1076 B.n408 B.n407 163.367
R1077 B.n407 B.n406 163.367
R1078 B.n716 B.n715 163.367
R1079 B.n715 B.n714 163.367
R1080 B.n714 B.n43 163.367
R1081 B.n710 B.n43 163.367
R1082 B.n710 B.n709 163.367
R1083 B.n709 B.n708 163.367
R1084 B.n708 B.n45 163.367
R1085 B.n704 B.n45 163.367
R1086 B.n704 B.n703 163.367
R1087 B.n703 B.n702 163.367
R1088 B.n702 B.n47 163.367
R1089 B.n698 B.n47 163.367
R1090 B.n698 B.n697 163.367
R1091 B.n697 B.n696 163.367
R1092 B.n696 B.n49 163.367
R1093 B.n692 B.n49 163.367
R1094 B.n692 B.n691 163.367
R1095 B.n691 B.n690 163.367
R1096 B.n690 B.n51 163.367
R1097 B.n685 B.n51 163.367
R1098 B.n685 B.n684 163.367
R1099 B.n684 B.n683 163.367
R1100 B.n683 B.n55 163.367
R1101 B.n679 B.n55 163.367
R1102 B.n679 B.n678 163.367
R1103 B.n678 B.n677 163.367
R1104 B.n677 B.n57 163.367
R1105 B.n672 B.n57 163.367
R1106 B.n672 B.n671 163.367
R1107 B.n671 B.n670 163.367
R1108 B.n670 B.n61 163.367
R1109 B.n666 B.n61 163.367
R1110 B.n666 B.n665 163.367
R1111 B.n665 B.n664 163.367
R1112 B.n664 B.n63 163.367
R1113 B.n660 B.n63 163.367
R1114 B.n660 B.n659 163.367
R1115 B.n659 B.n658 163.367
R1116 B.n658 B.n65 163.367
R1117 B.n654 B.n65 163.367
R1118 B.n654 B.n653 163.367
R1119 B.n653 B.n652 163.367
R1120 B.n652 B.n67 163.367
R1121 B.n648 B.n67 163.367
R1122 B.n648 B.n647 163.367
R1123 B.n647 B.n646 163.367
R1124 B.n720 B.n41 163.367
R1125 B.n721 B.n720 163.367
R1126 B.n722 B.n721 163.367
R1127 B.n722 B.n39 163.367
R1128 B.n726 B.n39 163.367
R1129 B.n727 B.n726 163.367
R1130 B.n728 B.n727 163.367
R1131 B.n728 B.n37 163.367
R1132 B.n732 B.n37 163.367
R1133 B.n733 B.n732 163.367
R1134 B.n734 B.n733 163.367
R1135 B.n734 B.n35 163.367
R1136 B.n738 B.n35 163.367
R1137 B.n739 B.n738 163.367
R1138 B.n740 B.n739 163.367
R1139 B.n740 B.n33 163.367
R1140 B.n744 B.n33 163.367
R1141 B.n745 B.n744 163.367
R1142 B.n746 B.n745 163.367
R1143 B.n746 B.n31 163.367
R1144 B.n750 B.n31 163.367
R1145 B.n751 B.n750 163.367
R1146 B.n752 B.n751 163.367
R1147 B.n752 B.n29 163.367
R1148 B.n756 B.n29 163.367
R1149 B.n757 B.n756 163.367
R1150 B.n758 B.n757 163.367
R1151 B.n758 B.n27 163.367
R1152 B.n762 B.n27 163.367
R1153 B.n763 B.n762 163.367
R1154 B.n764 B.n763 163.367
R1155 B.n764 B.n25 163.367
R1156 B.n768 B.n25 163.367
R1157 B.n769 B.n768 163.367
R1158 B.n770 B.n769 163.367
R1159 B.n770 B.n23 163.367
R1160 B.n774 B.n23 163.367
R1161 B.n775 B.n774 163.367
R1162 B.n776 B.n775 163.367
R1163 B.n776 B.n21 163.367
R1164 B.n780 B.n21 163.367
R1165 B.n781 B.n780 163.367
R1166 B.n782 B.n781 163.367
R1167 B.n782 B.n19 163.367
R1168 B.n786 B.n19 163.367
R1169 B.n787 B.n786 163.367
R1170 B.n788 B.n787 163.367
R1171 B.n788 B.n17 163.367
R1172 B.n792 B.n17 163.367
R1173 B.n793 B.n792 163.367
R1174 B.n794 B.n793 163.367
R1175 B.n794 B.n15 163.367
R1176 B.n798 B.n15 163.367
R1177 B.n799 B.n798 163.367
R1178 B.n800 B.n799 163.367
R1179 B.n800 B.n13 163.367
R1180 B.n804 B.n13 163.367
R1181 B.n805 B.n804 163.367
R1182 B.n806 B.n805 163.367
R1183 B.n806 B.n11 163.367
R1184 B.n810 B.n11 163.367
R1185 B.n811 B.n810 163.367
R1186 B.n812 B.n811 163.367
R1187 B.n812 B.n9 163.367
R1188 B.n816 B.n9 163.367
R1189 B.n817 B.n816 163.367
R1190 B.n818 B.n817 163.367
R1191 B.n818 B.n7 163.367
R1192 B.n822 B.n7 163.367
R1193 B.n823 B.n822 163.367
R1194 B.n824 B.n823 163.367
R1195 B.n824 B.n5 163.367
R1196 B.n828 B.n5 163.367
R1197 B.n829 B.n828 163.367
R1198 B.n830 B.n829 163.367
R1199 B.n830 B.n3 163.367
R1200 B.n834 B.n3 163.367
R1201 B.n835 B.n834 163.367
R1202 B.n213 B.n2 163.367
R1203 B.n216 B.n213 163.367
R1204 B.n217 B.n216 163.367
R1205 B.n218 B.n217 163.367
R1206 B.n218 B.n211 163.367
R1207 B.n222 B.n211 163.367
R1208 B.n223 B.n222 163.367
R1209 B.n224 B.n223 163.367
R1210 B.n224 B.n209 163.367
R1211 B.n228 B.n209 163.367
R1212 B.n229 B.n228 163.367
R1213 B.n230 B.n229 163.367
R1214 B.n230 B.n207 163.367
R1215 B.n234 B.n207 163.367
R1216 B.n235 B.n234 163.367
R1217 B.n236 B.n235 163.367
R1218 B.n236 B.n205 163.367
R1219 B.n240 B.n205 163.367
R1220 B.n241 B.n240 163.367
R1221 B.n242 B.n241 163.367
R1222 B.n242 B.n203 163.367
R1223 B.n246 B.n203 163.367
R1224 B.n247 B.n246 163.367
R1225 B.n248 B.n247 163.367
R1226 B.n248 B.n201 163.367
R1227 B.n252 B.n201 163.367
R1228 B.n253 B.n252 163.367
R1229 B.n254 B.n253 163.367
R1230 B.n254 B.n199 163.367
R1231 B.n258 B.n199 163.367
R1232 B.n259 B.n258 163.367
R1233 B.n260 B.n259 163.367
R1234 B.n260 B.n197 163.367
R1235 B.n264 B.n197 163.367
R1236 B.n265 B.n264 163.367
R1237 B.n266 B.n265 163.367
R1238 B.n266 B.n195 163.367
R1239 B.n270 B.n195 163.367
R1240 B.n271 B.n270 163.367
R1241 B.n272 B.n271 163.367
R1242 B.n272 B.n193 163.367
R1243 B.n276 B.n193 163.367
R1244 B.n277 B.n276 163.367
R1245 B.n278 B.n277 163.367
R1246 B.n278 B.n191 163.367
R1247 B.n282 B.n191 163.367
R1248 B.n283 B.n282 163.367
R1249 B.n284 B.n283 163.367
R1250 B.n284 B.n189 163.367
R1251 B.n288 B.n189 163.367
R1252 B.n289 B.n288 163.367
R1253 B.n290 B.n289 163.367
R1254 B.n290 B.n187 163.367
R1255 B.n294 B.n187 163.367
R1256 B.n295 B.n294 163.367
R1257 B.n296 B.n295 163.367
R1258 B.n296 B.n185 163.367
R1259 B.n300 B.n185 163.367
R1260 B.n301 B.n300 163.367
R1261 B.n302 B.n301 163.367
R1262 B.n302 B.n183 163.367
R1263 B.n306 B.n183 163.367
R1264 B.n307 B.n306 163.367
R1265 B.n308 B.n307 163.367
R1266 B.n308 B.n181 163.367
R1267 B.n312 B.n181 163.367
R1268 B.n313 B.n312 163.367
R1269 B.n314 B.n313 163.367
R1270 B.n314 B.n179 163.367
R1271 B.n318 B.n179 163.367
R1272 B.n319 B.n318 163.367
R1273 B.n320 B.n319 163.367
R1274 B.n320 B.n177 163.367
R1275 B.n324 B.n177 163.367
R1276 B.n325 B.n324 163.367
R1277 B.n326 B.n325 163.367
R1278 B.n326 B.n175 163.367
R1279 B.n330 B.n175 163.367
R1280 B.n373 B.t2 121.718
R1281 B.n59 B.t7 121.718
R1282 B.n165 B.t5 121.713
R1283 B.n53 B.t10 121.713
R1284 B.n165 B.n164 78.546
R1285 B.n373 B.n372 78.546
R1286 B.n59 B.n58 78.546
R1287 B.n53 B.n52 78.546
R1288 B.n359 B.n165 59.5399
R1289 B.n374 B.n373 59.5399
R1290 B.n674 B.n59 59.5399
R1291 B.n688 B.n53 59.5399
R1292 B.n718 B.n717 33.8737
R1293 B.n645 B.n644 33.8737
R1294 B.n405 B.n404 33.8737
R1295 B.n329 B.n174 33.8737
R1296 B B.n837 18.0485
R1297 B.n719 B.n718 10.6151
R1298 B.n719 B.n40 10.6151
R1299 B.n723 B.n40 10.6151
R1300 B.n724 B.n723 10.6151
R1301 B.n725 B.n724 10.6151
R1302 B.n725 B.n38 10.6151
R1303 B.n729 B.n38 10.6151
R1304 B.n730 B.n729 10.6151
R1305 B.n731 B.n730 10.6151
R1306 B.n731 B.n36 10.6151
R1307 B.n735 B.n36 10.6151
R1308 B.n736 B.n735 10.6151
R1309 B.n737 B.n736 10.6151
R1310 B.n737 B.n34 10.6151
R1311 B.n741 B.n34 10.6151
R1312 B.n742 B.n741 10.6151
R1313 B.n743 B.n742 10.6151
R1314 B.n743 B.n32 10.6151
R1315 B.n747 B.n32 10.6151
R1316 B.n748 B.n747 10.6151
R1317 B.n749 B.n748 10.6151
R1318 B.n749 B.n30 10.6151
R1319 B.n753 B.n30 10.6151
R1320 B.n754 B.n753 10.6151
R1321 B.n755 B.n754 10.6151
R1322 B.n755 B.n28 10.6151
R1323 B.n759 B.n28 10.6151
R1324 B.n760 B.n759 10.6151
R1325 B.n761 B.n760 10.6151
R1326 B.n761 B.n26 10.6151
R1327 B.n765 B.n26 10.6151
R1328 B.n766 B.n765 10.6151
R1329 B.n767 B.n766 10.6151
R1330 B.n767 B.n24 10.6151
R1331 B.n771 B.n24 10.6151
R1332 B.n772 B.n771 10.6151
R1333 B.n773 B.n772 10.6151
R1334 B.n773 B.n22 10.6151
R1335 B.n777 B.n22 10.6151
R1336 B.n778 B.n777 10.6151
R1337 B.n779 B.n778 10.6151
R1338 B.n779 B.n20 10.6151
R1339 B.n783 B.n20 10.6151
R1340 B.n784 B.n783 10.6151
R1341 B.n785 B.n784 10.6151
R1342 B.n785 B.n18 10.6151
R1343 B.n789 B.n18 10.6151
R1344 B.n790 B.n789 10.6151
R1345 B.n791 B.n790 10.6151
R1346 B.n791 B.n16 10.6151
R1347 B.n795 B.n16 10.6151
R1348 B.n796 B.n795 10.6151
R1349 B.n797 B.n796 10.6151
R1350 B.n797 B.n14 10.6151
R1351 B.n801 B.n14 10.6151
R1352 B.n802 B.n801 10.6151
R1353 B.n803 B.n802 10.6151
R1354 B.n803 B.n12 10.6151
R1355 B.n807 B.n12 10.6151
R1356 B.n808 B.n807 10.6151
R1357 B.n809 B.n808 10.6151
R1358 B.n809 B.n10 10.6151
R1359 B.n813 B.n10 10.6151
R1360 B.n814 B.n813 10.6151
R1361 B.n815 B.n814 10.6151
R1362 B.n815 B.n8 10.6151
R1363 B.n819 B.n8 10.6151
R1364 B.n820 B.n819 10.6151
R1365 B.n821 B.n820 10.6151
R1366 B.n821 B.n6 10.6151
R1367 B.n825 B.n6 10.6151
R1368 B.n826 B.n825 10.6151
R1369 B.n827 B.n826 10.6151
R1370 B.n827 B.n4 10.6151
R1371 B.n831 B.n4 10.6151
R1372 B.n832 B.n831 10.6151
R1373 B.n833 B.n832 10.6151
R1374 B.n833 B.n0 10.6151
R1375 B.n717 B.n42 10.6151
R1376 B.n713 B.n42 10.6151
R1377 B.n713 B.n712 10.6151
R1378 B.n712 B.n711 10.6151
R1379 B.n711 B.n44 10.6151
R1380 B.n707 B.n44 10.6151
R1381 B.n707 B.n706 10.6151
R1382 B.n706 B.n705 10.6151
R1383 B.n705 B.n46 10.6151
R1384 B.n701 B.n46 10.6151
R1385 B.n701 B.n700 10.6151
R1386 B.n700 B.n699 10.6151
R1387 B.n699 B.n48 10.6151
R1388 B.n695 B.n48 10.6151
R1389 B.n695 B.n694 10.6151
R1390 B.n694 B.n693 10.6151
R1391 B.n693 B.n50 10.6151
R1392 B.n689 B.n50 10.6151
R1393 B.n687 B.n686 10.6151
R1394 B.n686 B.n54 10.6151
R1395 B.n682 B.n54 10.6151
R1396 B.n682 B.n681 10.6151
R1397 B.n681 B.n680 10.6151
R1398 B.n680 B.n56 10.6151
R1399 B.n676 B.n56 10.6151
R1400 B.n676 B.n675 10.6151
R1401 B.n673 B.n60 10.6151
R1402 B.n669 B.n60 10.6151
R1403 B.n669 B.n668 10.6151
R1404 B.n668 B.n667 10.6151
R1405 B.n667 B.n62 10.6151
R1406 B.n663 B.n62 10.6151
R1407 B.n663 B.n662 10.6151
R1408 B.n662 B.n661 10.6151
R1409 B.n661 B.n64 10.6151
R1410 B.n657 B.n64 10.6151
R1411 B.n657 B.n656 10.6151
R1412 B.n656 B.n655 10.6151
R1413 B.n655 B.n66 10.6151
R1414 B.n651 B.n66 10.6151
R1415 B.n651 B.n650 10.6151
R1416 B.n650 B.n649 10.6151
R1417 B.n649 B.n68 10.6151
R1418 B.n645 B.n68 10.6151
R1419 B.n644 B.n643 10.6151
R1420 B.n643 B.n70 10.6151
R1421 B.n639 B.n70 10.6151
R1422 B.n639 B.n638 10.6151
R1423 B.n638 B.n637 10.6151
R1424 B.n637 B.n72 10.6151
R1425 B.n633 B.n72 10.6151
R1426 B.n633 B.n632 10.6151
R1427 B.n632 B.n631 10.6151
R1428 B.n631 B.n74 10.6151
R1429 B.n627 B.n74 10.6151
R1430 B.n627 B.n626 10.6151
R1431 B.n626 B.n625 10.6151
R1432 B.n625 B.n76 10.6151
R1433 B.n621 B.n76 10.6151
R1434 B.n621 B.n620 10.6151
R1435 B.n620 B.n619 10.6151
R1436 B.n619 B.n78 10.6151
R1437 B.n615 B.n78 10.6151
R1438 B.n615 B.n614 10.6151
R1439 B.n614 B.n613 10.6151
R1440 B.n613 B.n80 10.6151
R1441 B.n609 B.n80 10.6151
R1442 B.n609 B.n608 10.6151
R1443 B.n608 B.n607 10.6151
R1444 B.n607 B.n82 10.6151
R1445 B.n603 B.n82 10.6151
R1446 B.n603 B.n602 10.6151
R1447 B.n602 B.n601 10.6151
R1448 B.n601 B.n84 10.6151
R1449 B.n597 B.n84 10.6151
R1450 B.n597 B.n596 10.6151
R1451 B.n596 B.n595 10.6151
R1452 B.n595 B.n86 10.6151
R1453 B.n591 B.n86 10.6151
R1454 B.n591 B.n590 10.6151
R1455 B.n590 B.n589 10.6151
R1456 B.n589 B.n88 10.6151
R1457 B.n585 B.n88 10.6151
R1458 B.n585 B.n584 10.6151
R1459 B.n584 B.n583 10.6151
R1460 B.n583 B.n90 10.6151
R1461 B.n579 B.n90 10.6151
R1462 B.n579 B.n578 10.6151
R1463 B.n578 B.n577 10.6151
R1464 B.n577 B.n92 10.6151
R1465 B.n573 B.n92 10.6151
R1466 B.n573 B.n572 10.6151
R1467 B.n572 B.n571 10.6151
R1468 B.n571 B.n94 10.6151
R1469 B.n567 B.n94 10.6151
R1470 B.n567 B.n566 10.6151
R1471 B.n566 B.n565 10.6151
R1472 B.n565 B.n96 10.6151
R1473 B.n561 B.n96 10.6151
R1474 B.n561 B.n560 10.6151
R1475 B.n560 B.n559 10.6151
R1476 B.n559 B.n98 10.6151
R1477 B.n555 B.n98 10.6151
R1478 B.n555 B.n554 10.6151
R1479 B.n554 B.n553 10.6151
R1480 B.n553 B.n100 10.6151
R1481 B.n549 B.n100 10.6151
R1482 B.n549 B.n548 10.6151
R1483 B.n548 B.n547 10.6151
R1484 B.n547 B.n102 10.6151
R1485 B.n543 B.n102 10.6151
R1486 B.n543 B.n542 10.6151
R1487 B.n542 B.n541 10.6151
R1488 B.n541 B.n104 10.6151
R1489 B.n537 B.n104 10.6151
R1490 B.n537 B.n536 10.6151
R1491 B.n536 B.n535 10.6151
R1492 B.n535 B.n106 10.6151
R1493 B.n531 B.n106 10.6151
R1494 B.n531 B.n530 10.6151
R1495 B.n530 B.n529 10.6151
R1496 B.n529 B.n108 10.6151
R1497 B.n525 B.n108 10.6151
R1498 B.n525 B.n524 10.6151
R1499 B.n524 B.n523 10.6151
R1500 B.n523 B.n110 10.6151
R1501 B.n519 B.n110 10.6151
R1502 B.n519 B.n518 10.6151
R1503 B.n518 B.n517 10.6151
R1504 B.n517 B.n112 10.6151
R1505 B.n513 B.n112 10.6151
R1506 B.n513 B.n512 10.6151
R1507 B.n512 B.n511 10.6151
R1508 B.n511 B.n114 10.6151
R1509 B.n507 B.n114 10.6151
R1510 B.n507 B.n506 10.6151
R1511 B.n506 B.n505 10.6151
R1512 B.n505 B.n116 10.6151
R1513 B.n501 B.n116 10.6151
R1514 B.n501 B.n500 10.6151
R1515 B.n500 B.n499 10.6151
R1516 B.n499 B.n118 10.6151
R1517 B.n495 B.n118 10.6151
R1518 B.n495 B.n494 10.6151
R1519 B.n494 B.n493 10.6151
R1520 B.n493 B.n120 10.6151
R1521 B.n489 B.n120 10.6151
R1522 B.n489 B.n488 10.6151
R1523 B.n488 B.n487 10.6151
R1524 B.n487 B.n122 10.6151
R1525 B.n483 B.n122 10.6151
R1526 B.n483 B.n482 10.6151
R1527 B.n482 B.n481 10.6151
R1528 B.n481 B.n124 10.6151
R1529 B.n477 B.n124 10.6151
R1530 B.n477 B.n476 10.6151
R1531 B.n476 B.n475 10.6151
R1532 B.n475 B.n126 10.6151
R1533 B.n471 B.n126 10.6151
R1534 B.n471 B.n470 10.6151
R1535 B.n470 B.n469 10.6151
R1536 B.n469 B.n128 10.6151
R1537 B.n465 B.n128 10.6151
R1538 B.n465 B.n464 10.6151
R1539 B.n464 B.n463 10.6151
R1540 B.n463 B.n130 10.6151
R1541 B.n459 B.n130 10.6151
R1542 B.n459 B.n458 10.6151
R1543 B.n458 B.n457 10.6151
R1544 B.n457 B.n132 10.6151
R1545 B.n453 B.n132 10.6151
R1546 B.n453 B.n452 10.6151
R1547 B.n452 B.n451 10.6151
R1548 B.n451 B.n134 10.6151
R1549 B.n447 B.n134 10.6151
R1550 B.n447 B.n446 10.6151
R1551 B.n446 B.n445 10.6151
R1552 B.n445 B.n136 10.6151
R1553 B.n441 B.n136 10.6151
R1554 B.n441 B.n440 10.6151
R1555 B.n440 B.n439 10.6151
R1556 B.n439 B.n138 10.6151
R1557 B.n435 B.n138 10.6151
R1558 B.n435 B.n434 10.6151
R1559 B.n434 B.n433 10.6151
R1560 B.n433 B.n140 10.6151
R1561 B.n429 B.n140 10.6151
R1562 B.n429 B.n428 10.6151
R1563 B.n428 B.n427 10.6151
R1564 B.n427 B.n142 10.6151
R1565 B.n423 B.n142 10.6151
R1566 B.n423 B.n422 10.6151
R1567 B.n422 B.n421 10.6151
R1568 B.n421 B.n144 10.6151
R1569 B.n417 B.n144 10.6151
R1570 B.n417 B.n416 10.6151
R1571 B.n416 B.n415 10.6151
R1572 B.n415 B.n146 10.6151
R1573 B.n411 B.n146 10.6151
R1574 B.n411 B.n410 10.6151
R1575 B.n410 B.n409 10.6151
R1576 B.n409 B.n148 10.6151
R1577 B.n405 B.n148 10.6151
R1578 B.n214 B.n1 10.6151
R1579 B.n215 B.n214 10.6151
R1580 B.n215 B.n212 10.6151
R1581 B.n219 B.n212 10.6151
R1582 B.n220 B.n219 10.6151
R1583 B.n221 B.n220 10.6151
R1584 B.n221 B.n210 10.6151
R1585 B.n225 B.n210 10.6151
R1586 B.n226 B.n225 10.6151
R1587 B.n227 B.n226 10.6151
R1588 B.n227 B.n208 10.6151
R1589 B.n231 B.n208 10.6151
R1590 B.n232 B.n231 10.6151
R1591 B.n233 B.n232 10.6151
R1592 B.n233 B.n206 10.6151
R1593 B.n237 B.n206 10.6151
R1594 B.n238 B.n237 10.6151
R1595 B.n239 B.n238 10.6151
R1596 B.n239 B.n204 10.6151
R1597 B.n243 B.n204 10.6151
R1598 B.n244 B.n243 10.6151
R1599 B.n245 B.n244 10.6151
R1600 B.n245 B.n202 10.6151
R1601 B.n249 B.n202 10.6151
R1602 B.n250 B.n249 10.6151
R1603 B.n251 B.n250 10.6151
R1604 B.n251 B.n200 10.6151
R1605 B.n255 B.n200 10.6151
R1606 B.n256 B.n255 10.6151
R1607 B.n257 B.n256 10.6151
R1608 B.n257 B.n198 10.6151
R1609 B.n261 B.n198 10.6151
R1610 B.n262 B.n261 10.6151
R1611 B.n263 B.n262 10.6151
R1612 B.n263 B.n196 10.6151
R1613 B.n267 B.n196 10.6151
R1614 B.n268 B.n267 10.6151
R1615 B.n269 B.n268 10.6151
R1616 B.n269 B.n194 10.6151
R1617 B.n273 B.n194 10.6151
R1618 B.n274 B.n273 10.6151
R1619 B.n275 B.n274 10.6151
R1620 B.n275 B.n192 10.6151
R1621 B.n279 B.n192 10.6151
R1622 B.n280 B.n279 10.6151
R1623 B.n281 B.n280 10.6151
R1624 B.n281 B.n190 10.6151
R1625 B.n285 B.n190 10.6151
R1626 B.n286 B.n285 10.6151
R1627 B.n287 B.n286 10.6151
R1628 B.n287 B.n188 10.6151
R1629 B.n291 B.n188 10.6151
R1630 B.n292 B.n291 10.6151
R1631 B.n293 B.n292 10.6151
R1632 B.n293 B.n186 10.6151
R1633 B.n297 B.n186 10.6151
R1634 B.n298 B.n297 10.6151
R1635 B.n299 B.n298 10.6151
R1636 B.n299 B.n184 10.6151
R1637 B.n303 B.n184 10.6151
R1638 B.n304 B.n303 10.6151
R1639 B.n305 B.n304 10.6151
R1640 B.n305 B.n182 10.6151
R1641 B.n309 B.n182 10.6151
R1642 B.n310 B.n309 10.6151
R1643 B.n311 B.n310 10.6151
R1644 B.n311 B.n180 10.6151
R1645 B.n315 B.n180 10.6151
R1646 B.n316 B.n315 10.6151
R1647 B.n317 B.n316 10.6151
R1648 B.n317 B.n178 10.6151
R1649 B.n321 B.n178 10.6151
R1650 B.n322 B.n321 10.6151
R1651 B.n323 B.n322 10.6151
R1652 B.n323 B.n176 10.6151
R1653 B.n327 B.n176 10.6151
R1654 B.n328 B.n327 10.6151
R1655 B.n329 B.n328 10.6151
R1656 B.n333 B.n174 10.6151
R1657 B.n334 B.n333 10.6151
R1658 B.n335 B.n334 10.6151
R1659 B.n335 B.n172 10.6151
R1660 B.n339 B.n172 10.6151
R1661 B.n340 B.n339 10.6151
R1662 B.n341 B.n340 10.6151
R1663 B.n341 B.n170 10.6151
R1664 B.n345 B.n170 10.6151
R1665 B.n346 B.n345 10.6151
R1666 B.n347 B.n346 10.6151
R1667 B.n347 B.n168 10.6151
R1668 B.n351 B.n168 10.6151
R1669 B.n352 B.n351 10.6151
R1670 B.n353 B.n352 10.6151
R1671 B.n353 B.n166 10.6151
R1672 B.n357 B.n166 10.6151
R1673 B.n358 B.n357 10.6151
R1674 B.n360 B.n162 10.6151
R1675 B.n364 B.n162 10.6151
R1676 B.n365 B.n364 10.6151
R1677 B.n366 B.n365 10.6151
R1678 B.n366 B.n160 10.6151
R1679 B.n370 B.n160 10.6151
R1680 B.n371 B.n370 10.6151
R1681 B.n375 B.n371 10.6151
R1682 B.n379 B.n158 10.6151
R1683 B.n380 B.n379 10.6151
R1684 B.n381 B.n380 10.6151
R1685 B.n381 B.n156 10.6151
R1686 B.n385 B.n156 10.6151
R1687 B.n386 B.n385 10.6151
R1688 B.n387 B.n386 10.6151
R1689 B.n387 B.n154 10.6151
R1690 B.n391 B.n154 10.6151
R1691 B.n392 B.n391 10.6151
R1692 B.n393 B.n392 10.6151
R1693 B.n393 B.n152 10.6151
R1694 B.n397 B.n152 10.6151
R1695 B.n398 B.n397 10.6151
R1696 B.n399 B.n398 10.6151
R1697 B.n399 B.n150 10.6151
R1698 B.n403 B.n150 10.6151
R1699 B.n404 B.n403 10.6151
R1700 B.n837 B.n0 8.11757
R1701 B.n837 B.n1 8.11757
R1702 B.n688 B.n687 6.5566
R1703 B.n675 B.n674 6.5566
R1704 B.n360 B.n359 6.5566
R1705 B.n375 B.n374 6.5566
R1706 B.n689 B.n688 4.05904
R1707 B.n674 B.n673 4.05904
R1708 B.n359 B.n358 4.05904
R1709 B.n374 B.n158 4.05904
C0 VP B 2.81987f
C1 VN w_n5830_n1814# 12.699401f
C2 VDD2 VP 0.73061f
C3 VN B 1.53167f
C4 VDD2 VN 4.36179f
C5 VDD1 w_n5830_n1814# 2.6768f
C6 VTAIL w_n5830_n1814# 2.30067f
C7 VN VP 8.617241f
C8 VDD1 B 2.28805f
C9 VDD2 VDD1 2.90175f
C10 VTAIL B 2.25954f
C11 VDD2 VTAIL 7.97671f
C12 VDD1 VP 4.92869f
C13 VTAIL VP 6.1881f
C14 VDD1 VN 0.15986f
C15 VTAIL VN 6.17383f
C16 VDD1 VTAIL 7.9161f
C17 B w_n5830_n1814# 10.283099f
C18 VDD2 w_n5830_n1814# 2.87821f
C19 VP w_n5830_n1814# 13.4613f
C20 VDD2 B 2.44978f
C21 VDD2 VSUBS 2.545888f
C22 VDD1 VSUBS 2.271761f
C23 VTAIL VSUBS 0.771119f
C24 VN VSUBS 9.39312f
C25 VP VSUBS 4.968506f
C26 B VSUBS 5.721764f
C27 w_n5830_n1814# VSUBS 0.132994p
C28 B.n0 VSUBS 0.011511f
C29 B.n1 VSUBS 0.011511f
C30 B.n2 VSUBS 0.017024f
C31 B.n3 VSUBS 0.013046f
C32 B.n4 VSUBS 0.013046f
C33 B.n5 VSUBS 0.013046f
C34 B.n6 VSUBS 0.013046f
C35 B.n7 VSUBS 0.013046f
C36 B.n8 VSUBS 0.013046f
C37 B.n9 VSUBS 0.013046f
C38 B.n10 VSUBS 0.013046f
C39 B.n11 VSUBS 0.013046f
C40 B.n12 VSUBS 0.013046f
C41 B.n13 VSUBS 0.013046f
C42 B.n14 VSUBS 0.013046f
C43 B.n15 VSUBS 0.013046f
C44 B.n16 VSUBS 0.013046f
C45 B.n17 VSUBS 0.013046f
C46 B.n18 VSUBS 0.013046f
C47 B.n19 VSUBS 0.013046f
C48 B.n20 VSUBS 0.013046f
C49 B.n21 VSUBS 0.013046f
C50 B.n22 VSUBS 0.013046f
C51 B.n23 VSUBS 0.013046f
C52 B.n24 VSUBS 0.013046f
C53 B.n25 VSUBS 0.013046f
C54 B.n26 VSUBS 0.013046f
C55 B.n27 VSUBS 0.013046f
C56 B.n28 VSUBS 0.013046f
C57 B.n29 VSUBS 0.013046f
C58 B.n30 VSUBS 0.013046f
C59 B.n31 VSUBS 0.013046f
C60 B.n32 VSUBS 0.013046f
C61 B.n33 VSUBS 0.013046f
C62 B.n34 VSUBS 0.013046f
C63 B.n35 VSUBS 0.013046f
C64 B.n36 VSUBS 0.013046f
C65 B.n37 VSUBS 0.013046f
C66 B.n38 VSUBS 0.013046f
C67 B.n39 VSUBS 0.013046f
C68 B.n40 VSUBS 0.013046f
C69 B.n41 VSUBS 0.030528f
C70 B.n42 VSUBS 0.013046f
C71 B.n43 VSUBS 0.013046f
C72 B.n44 VSUBS 0.013046f
C73 B.n45 VSUBS 0.013046f
C74 B.n46 VSUBS 0.013046f
C75 B.n47 VSUBS 0.013046f
C76 B.n48 VSUBS 0.013046f
C77 B.n49 VSUBS 0.013046f
C78 B.n50 VSUBS 0.013046f
C79 B.n51 VSUBS 0.013046f
C80 B.t10 VSUBS 0.210409f
C81 B.t11 VSUBS 0.256962f
C82 B.t9 VSUBS 1.42493f
C83 B.n52 VSUBS 0.19253f
C84 B.n53 VSUBS 0.1373f
C85 B.n54 VSUBS 0.013046f
C86 B.n55 VSUBS 0.013046f
C87 B.n56 VSUBS 0.013046f
C88 B.n57 VSUBS 0.013046f
C89 B.t7 VSUBS 0.210409f
C90 B.t8 VSUBS 0.256962f
C91 B.t6 VSUBS 1.42493f
C92 B.n58 VSUBS 0.19253f
C93 B.n59 VSUBS 0.1373f
C94 B.n60 VSUBS 0.013046f
C95 B.n61 VSUBS 0.013046f
C96 B.n62 VSUBS 0.013046f
C97 B.n63 VSUBS 0.013046f
C98 B.n64 VSUBS 0.013046f
C99 B.n65 VSUBS 0.013046f
C100 B.n66 VSUBS 0.013046f
C101 B.n67 VSUBS 0.013046f
C102 B.n68 VSUBS 0.013046f
C103 B.n69 VSUBS 0.030528f
C104 B.n70 VSUBS 0.013046f
C105 B.n71 VSUBS 0.013046f
C106 B.n72 VSUBS 0.013046f
C107 B.n73 VSUBS 0.013046f
C108 B.n74 VSUBS 0.013046f
C109 B.n75 VSUBS 0.013046f
C110 B.n76 VSUBS 0.013046f
C111 B.n77 VSUBS 0.013046f
C112 B.n78 VSUBS 0.013046f
C113 B.n79 VSUBS 0.013046f
C114 B.n80 VSUBS 0.013046f
C115 B.n81 VSUBS 0.013046f
C116 B.n82 VSUBS 0.013046f
C117 B.n83 VSUBS 0.013046f
C118 B.n84 VSUBS 0.013046f
C119 B.n85 VSUBS 0.013046f
C120 B.n86 VSUBS 0.013046f
C121 B.n87 VSUBS 0.013046f
C122 B.n88 VSUBS 0.013046f
C123 B.n89 VSUBS 0.013046f
C124 B.n90 VSUBS 0.013046f
C125 B.n91 VSUBS 0.013046f
C126 B.n92 VSUBS 0.013046f
C127 B.n93 VSUBS 0.013046f
C128 B.n94 VSUBS 0.013046f
C129 B.n95 VSUBS 0.013046f
C130 B.n96 VSUBS 0.013046f
C131 B.n97 VSUBS 0.013046f
C132 B.n98 VSUBS 0.013046f
C133 B.n99 VSUBS 0.013046f
C134 B.n100 VSUBS 0.013046f
C135 B.n101 VSUBS 0.013046f
C136 B.n102 VSUBS 0.013046f
C137 B.n103 VSUBS 0.013046f
C138 B.n104 VSUBS 0.013046f
C139 B.n105 VSUBS 0.013046f
C140 B.n106 VSUBS 0.013046f
C141 B.n107 VSUBS 0.013046f
C142 B.n108 VSUBS 0.013046f
C143 B.n109 VSUBS 0.013046f
C144 B.n110 VSUBS 0.013046f
C145 B.n111 VSUBS 0.013046f
C146 B.n112 VSUBS 0.013046f
C147 B.n113 VSUBS 0.013046f
C148 B.n114 VSUBS 0.013046f
C149 B.n115 VSUBS 0.013046f
C150 B.n116 VSUBS 0.013046f
C151 B.n117 VSUBS 0.013046f
C152 B.n118 VSUBS 0.013046f
C153 B.n119 VSUBS 0.013046f
C154 B.n120 VSUBS 0.013046f
C155 B.n121 VSUBS 0.013046f
C156 B.n122 VSUBS 0.013046f
C157 B.n123 VSUBS 0.013046f
C158 B.n124 VSUBS 0.013046f
C159 B.n125 VSUBS 0.013046f
C160 B.n126 VSUBS 0.013046f
C161 B.n127 VSUBS 0.013046f
C162 B.n128 VSUBS 0.013046f
C163 B.n129 VSUBS 0.013046f
C164 B.n130 VSUBS 0.013046f
C165 B.n131 VSUBS 0.013046f
C166 B.n132 VSUBS 0.013046f
C167 B.n133 VSUBS 0.013046f
C168 B.n134 VSUBS 0.013046f
C169 B.n135 VSUBS 0.013046f
C170 B.n136 VSUBS 0.013046f
C171 B.n137 VSUBS 0.013046f
C172 B.n138 VSUBS 0.013046f
C173 B.n139 VSUBS 0.013046f
C174 B.n140 VSUBS 0.013046f
C175 B.n141 VSUBS 0.013046f
C176 B.n142 VSUBS 0.013046f
C177 B.n143 VSUBS 0.013046f
C178 B.n144 VSUBS 0.013046f
C179 B.n145 VSUBS 0.013046f
C180 B.n146 VSUBS 0.013046f
C181 B.n147 VSUBS 0.013046f
C182 B.n148 VSUBS 0.013046f
C183 B.n149 VSUBS 0.032014f
C184 B.n150 VSUBS 0.013046f
C185 B.n151 VSUBS 0.013046f
C186 B.n152 VSUBS 0.013046f
C187 B.n153 VSUBS 0.013046f
C188 B.n154 VSUBS 0.013046f
C189 B.n155 VSUBS 0.013046f
C190 B.n156 VSUBS 0.013046f
C191 B.n157 VSUBS 0.013046f
C192 B.n158 VSUBS 0.009017f
C193 B.n159 VSUBS 0.013046f
C194 B.n160 VSUBS 0.013046f
C195 B.n161 VSUBS 0.013046f
C196 B.n162 VSUBS 0.013046f
C197 B.n163 VSUBS 0.013046f
C198 B.t5 VSUBS 0.210409f
C199 B.t4 VSUBS 0.256962f
C200 B.t3 VSUBS 1.42493f
C201 B.n164 VSUBS 0.19253f
C202 B.n165 VSUBS 0.1373f
C203 B.n166 VSUBS 0.013046f
C204 B.n167 VSUBS 0.013046f
C205 B.n168 VSUBS 0.013046f
C206 B.n169 VSUBS 0.013046f
C207 B.n170 VSUBS 0.013046f
C208 B.n171 VSUBS 0.013046f
C209 B.n172 VSUBS 0.013046f
C210 B.n173 VSUBS 0.013046f
C211 B.n174 VSUBS 0.032014f
C212 B.n175 VSUBS 0.013046f
C213 B.n176 VSUBS 0.013046f
C214 B.n177 VSUBS 0.013046f
C215 B.n178 VSUBS 0.013046f
C216 B.n179 VSUBS 0.013046f
C217 B.n180 VSUBS 0.013046f
C218 B.n181 VSUBS 0.013046f
C219 B.n182 VSUBS 0.013046f
C220 B.n183 VSUBS 0.013046f
C221 B.n184 VSUBS 0.013046f
C222 B.n185 VSUBS 0.013046f
C223 B.n186 VSUBS 0.013046f
C224 B.n187 VSUBS 0.013046f
C225 B.n188 VSUBS 0.013046f
C226 B.n189 VSUBS 0.013046f
C227 B.n190 VSUBS 0.013046f
C228 B.n191 VSUBS 0.013046f
C229 B.n192 VSUBS 0.013046f
C230 B.n193 VSUBS 0.013046f
C231 B.n194 VSUBS 0.013046f
C232 B.n195 VSUBS 0.013046f
C233 B.n196 VSUBS 0.013046f
C234 B.n197 VSUBS 0.013046f
C235 B.n198 VSUBS 0.013046f
C236 B.n199 VSUBS 0.013046f
C237 B.n200 VSUBS 0.013046f
C238 B.n201 VSUBS 0.013046f
C239 B.n202 VSUBS 0.013046f
C240 B.n203 VSUBS 0.013046f
C241 B.n204 VSUBS 0.013046f
C242 B.n205 VSUBS 0.013046f
C243 B.n206 VSUBS 0.013046f
C244 B.n207 VSUBS 0.013046f
C245 B.n208 VSUBS 0.013046f
C246 B.n209 VSUBS 0.013046f
C247 B.n210 VSUBS 0.013046f
C248 B.n211 VSUBS 0.013046f
C249 B.n212 VSUBS 0.013046f
C250 B.n213 VSUBS 0.013046f
C251 B.n214 VSUBS 0.013046f
C252 B.n215 VSUBS 0.013046f
C253 B.n216 VSUBS 0.013046f
C254 B.n217 VSUBS 0.013046f
C255 B.n218 VSUBS 0.013046f
C256 B.n219 VSUBS 0.013046f
C257 B.n220 VSUBS 0.013046f
C258 B.n221 VSUBS 0.013046f
C259 B.n222 VSUBS 0.013046f
C260 B.n223 VSUBS 0.013046f
C261 B.n224 VSUBS 0.013046f
C262 B.n225 VSUBS 0.013046f
C263 B.n226 VSUBS 0.013046f
C264 B.n227 VSUBS 0.013046f
C265 B.n228 VSUBS 0.013046f
C266 B.n229 VSUBS 0.013046f
C267 B.n230 VSUBS 0.013046f
C268 B.n231 VSUBS 0.013046f
C269 B.n232 VSUBS 0.013046f
C270 B.n233 VSUBS 0.013046f
C271 B.n234 VSUBS 0.013046f
C272 B.n235 VSUBS 0.013046f
C273 B.n236 VSUBS 0.013046f
C274 B.n237 VSUBS 0.013046f
C275 B.n238 VSUBS 0.013046f
C276 B.n239 VSUBS 0.013046f
C277 B.n240 VSUBS 0.013046f
C278 B.n241 VSUBS 0.013046f
C279 B.n242 VSUBS 0.013046f
C280 B.n243 VSUBS 0.013046f
C281 B.n244 VSUBS 0.013046f
C282 B.n245 VSUBS 0.013046f
C283 B.n246 VSUBS 0.013046f
C284 B.n247 VSUBS 0.013046f
C285 B.n248 VSUBS 0.013046f
C286 B.n249 VSUBS 0.013046f
C287 B.n250 VSUBS 0.013046f
C288 B.n251 VSUBS 0.013046f
C289 B.n252 VSUBS 0.013046f
C290 B.n253 VSUBS 0.013046f
C291 B.n254 VSUBS 0.013046f
C292 B.n255 VSUBS 0.013046f
C293 B.n256 VSUBS 0.013046f
C294 B.n257 VSUBS 0.013046f
C295 B.n258 VSUBS 0.013046f
C296 B.n259 VSUBS 0.013046f
C297 B.n260 VSUBS 0.013046f
C298 B.n261 VSUBS 0.013046f
C299 B.n262 VSUBS 0.013046f
C300 B.n263 VSUBS 0.013046f
C301 B.n264 VSUBS 0.013046f
C302 B.n265 VSUBS 0.013046f
C303 B.n266 VSUBS 0.013046f
C304 B.n267 VSUBS 0.013046f
C305 B.n268 VSUBS 0.013046f
C306 B.n269 VSUBS 0.013046f
C307 B.n270 VSUBS 0.013046f
C308 B.n271 VSUBS 0.013046f
C309 B.n272 VSUBS 0.013046f
C310 B.n273 VSUBS 0.013046f
C311 B.n274 VSUBS 0.013046f
C312 B.n275 VSUBS 0.013046f
C313 B.n276 VSUBS 0.013046f
C314 B.n277 VSUBS 0.013046f
C315 B.n278 VSUBS 0.013046f
C316 B.n279 VSUBS 0.013046f
C317 B.n280 VSUBS 0.013046f
C318 B.n281 VSUBS 0.013046f
C319 B.n282 VSUBS 0.013046f
C320 B.n283 VSUBS 0.013046f
C321 B.n284 VSUBS 0.013046f
C322 B.n285 VSUBS 0.013046f
C323 B.n286 VSUBS 0.013046f
C324 B.n287 VSUBS 0.013046f
C325 B.n288 VSUBS 0.013046f
C326 B.n289 VSUBS 0.013046f
C327 B.n290 VSUBS 0.013046f
C328 B.n291 VSUBS 0.013046f
C329 B.n292 VSUBS 0.013046f
C330 B.n293 VSUBS 0.013046f
C331 B.n294 VSUBS 0.013046f
C332 B.n295 VSUBS 0.013046f
C333 B.n296 VSUBS 0.013046f
C334 B.n297 VSUBS 0.013046f
C335 B.n298 VSUBS 0.013046f
C336 B.n299 VSUBS 0.013046f
C337 B.n300 VSUBS 0.013046f
C338 B.n301 VSUBS 0.013046f
C339 B.n302 VSUBS 0.013046f
C340 B.n303 VSUBS 0.013046f
C341 B.n304 VSUBS 0.013046f
C342 B.n305 VSUBS 0.013046f
C343 B.n306 VSUBS 0.013046f
C344 B.n307 VSUBS 0.013046f
C345 B.n308 VSUBS 0.013046f
C346 B.n309 VSUBS 0.013046f
C347 B.n310 VSUBS 0.013046f
C348 B.n311 VSUBS 0.013046f
C349 B.n312 VSUBS 0.013046f
C350 B.n313 VSUBS 0.013046f
C351 B.n314 VSUBS 0.013046f
C352 B.n315 VSUBS 0.013046f
C353 B.n316 VSUBS 0.013046f
C354 B.n317 VSUBS 0.013046f
C355 B.n318 VSUBS 0.013046f
C356 B.n319 VSUBS 0.013046f
C357 B.n320 VSUBS 0.013046f
C358 B.n321 VSUBS 0.013046f
C359 B.n322 VSUBS 0.013046f
C360 B.n323 VSUBS 0.013046f
C361 B.n324 VSUBS 0.013046f
C362 B.n325 VSUBS 0.013046f
C363 B.n326 VSUBS 0.013046f
C364 B.n327 VSUBS 0.013046f
C365 B.n328 VSUBS 0.013046f
C366 B.n329 VSUBS 0.030528f
C367 B.n330 VSUBS 0.030528f
C368 B.n331 VSUBS 0.032014f
C369 B.n332 VSUBS 0.013046f
C370 B.n333 VSUBS 0.013046f
C371 B.n334 VSUBS 0.013046f
C372 B.n335 VSUBS 0.013046f
C373 B.n336 VSUBS 0.013046f
C374 B.n337 VSUBS 0.013046f
C375 B.n338 VSUBS 0.013046f
C376 B.n339 VSUBS 0.013046f
C377 B.n340 VSUBS 0.013046f
C378 B.n341 VSUBS 0.013046f
C379 B.n342 VSUBS 0.013046f
C380 B.n343 VSUBS 0.013046f
C381 B.n344 VSUBS 0.013046f
C382 B.n345 VSUBS 0.013046f
C383 B.n346 VSUBS 0.013046f
C384 B.n347 VSUBS 0.013046f
C385 B.n348 VSUBS 0.013046f
C386 B.n349 VSUBS 0.013046f
C387 B.n350 VSUBS 0.013046f
C388 B.n351 VSUBS 0.013046f
C389 B.n352 VSUBS 0.013046f
C390 B.n353 VSUBS 0.013046f
C391 B.n354 VSUBS 0.013046f
C392 B.n355 VSUBS 0.013046f
C393 B.n356 VSUBS 0.013046f
C394 B.n357 VSUBS 0.013046f
C395 B.n358 VSUBS 0.009017f
C396 B.n359 VSUBS 0.030225f
C397 B.n360 VSUBS 0.010552f
C398 B.n361 VSUBS 0.013046f
C399 B.n362 VSUBS 0.013046f
C400 B.n363 VSUBS 0.013046f
C401 B.n364 VSUBS 0.013046f
C402 B.n365 VSUBS 0.013046f
C403 B.n366 VSUBS 0.013046f
C404 B.n367 VSUBS 0.013046f
C405 B.n368 VSUBS 0.013046f
C406 B.n369 VSUBS 0.013046f
C407 B.n370 VSUBS 0.013046f
C408 B.n371 VSUBS 0.013046f
C409 B.t2 VSUBS 0.210409f
C410 B.t1 VSUBS 0.256962f
C411 B.t0 VSUBS 1.42493f
C412 B.n372 VSUBS 0.19253f
C413 B.n373 VSUBS 0.1373f
C414 B.n374 VSUBS 0.030225f
C415 B.n375 VSUBS 0.010552f
C416 B.n376 VSUBS 0.013046f
C417 B.n377 VSUBS 0.013046f
C418 B.n378 VSUBS 0.013046f
C419 B.n379 VSUBS 0.013046f
C420 B.n380 VSUBS 0.013046f
C421 B.n381 VSUBS 0.013046f
C422 B.n382 VSUBS 0.013046f
C423 B.n383 VSUBS 0.013046f
C424 B.n384 VSUBS 0.013046f
C425 B.n385 VSUBS 0.013046f
C426 B.n386 VSUBS 0.013046f
C427 B.n387 VSUBS 0.013046f
C428 B.n388 VSUBS 0.013046f
C429 B.n389 VSUBS 0.013046f
C430 B.n390 VSUBS 0.013046f
C431 B.n391 VSUBS 0.013046f
C432 B.n392 VSUBS 0.013046f
C433 B.n393 VSUBS 0.013046f
C434 B.n394 VSUBS 0.013046f
C435 B.n395 VSUBS 0.013046f
C436 B.n396 VSUBS 0.013046f
C437 B.n397 VSUBS 0.013046f
C438 B.n398 VSUBS 0.013046f
C439 B.n399 VSUBS 0.013046f
C440 B.n400 VSUBS 0.013046f
C441 B.n401 VSUBS 0.013046f
C442 B.n402 VSUBS 0.013046f
C443 B.n403 VSUBS 0.013046f
C444 B.n404 VSUBS 0.030528f
C445 B.n405 VSUBS 0.032014f
C446 B.n406 VSUBS 0.030528f
C447 B.n407 VSUBS 0.013046f
C448 B.n408 VSUBS 0.013046f
C449 B.n409 VSUBS 0.013046f
C450 B.n410 VSUBS 0.013046f
C451 B.n411 VSUBS 0.013046f
C452 B.n412 VSUBS 0.013046f
C453 B.n413 VSUBS 0.013046f
C454 B.n414 VSUBS 0.013046f
C455 B.n415 VSUBS 0.013046f
C456 B.n416 VSUBS 0.013046f
C457 B.n417 VSUBS 0.013046f
C458 B.n418 VSUBS 0.013046f
C459 B.n419 VSUBS 0.013046f
C460 B.n420 VSUBS 0.013046f
C461 B.n421 VSUBS 0.013046f
C462 B.n422 VSUBS 0.013046f
C463 B.n423 VSUBS 0.013046f
C464 B.n424 VSUBS 0.013046f
C465 B.n425 VSUBS 0.013046f
C466 B.n426 VSUBS 0.013046f
C467 B.n427 VSUBS 0.013046f
C468 B.n428 VSUBS 0.013046f
C469 B.n429 VSUBS 0.013046f
C470 B.n430 VSUBS 0.013046f
C471 B.n431 VSUBS 0.013046f
C472 B.n432 VSUBS 0.013046f
C473 B.n433 VSUBS 0.013046f
C474 B.n434 VSUBS 0.013046f
C475 B.n435 VSUBS 0.013046f
C476 B.n436 VSUBS 0.013046f
C477 B.n437 VSUBS 0.013046f
C478 B.n438 VSUBS 0.013046f
C479 B.n439 VSUBS 0.013046f
C480 B.n440 VSUBS 0.013046f
C481 B.n441 VSUBS 0.013046f
C482 B.n442 VSUBS 0.013046f
C483 B.n443 VSUBS 0.013046f
C484 B.n444 VSUBS 0.013046f
C485 B.n445 VSUBS 0.013046f
C486 B.n446 VSUBS 0.013046f
C487 B.n447 VSUBS 0.013046f
C488 B.n448 VSUBS 0.013046f
C489 B.n449 VSUBS 0.013046f
C490 B.n450 VSUBS 0.013046f
C491 B.n451 VSUBS 0.013046f
C492 B.n452 VSUBS 0.013046f
C493 B.n453 VSUBS 0.013046f
C494 B.n454 VSUBS 0.013046f
C495 B.n455 VSUBS 0.013046f
C496 B.n456 VSUBS 0.013046f
C497 B.n457 VSUBS 0.013046f
C498 B.n458 VSUBS 0.013046f
C499 B.n459 VSUBS 0.013046f
C500 B.n460 VSUBS 0.013046f
C501 B.n461 VSUBS 0.013046f
C502 B.n462 VSUBS 0.013046f
C503 B.n463 VSUBS 0.013046f
C504 B.n464 VSUBS 0.013046f
C505 B.n465 VSUBS 0.013046f
C506 B.n466 VSUBS 0.013046f
C507 B.n467 VSUBS 0.013046f
C508 B.n468 VSUBS 0.013046f
C509 B.n469 VSUBS 0.013046f
C510 B.n470 VSUBS 0.013046f
C511 B.n471 VSUBS 0.013046f
C512 B.n472 VSUBS 0.013046f
C513 B.n473 VSUBS 0.013046f
C514 B.n474 VSUBS 0.013046f
C515 B.n475 VSUBS 0.013046f
C516 B.n476 VSUBS 0.013046f
C517 B.n477 VSUBS 0.013046f
C518 B.n478 VSUBS 0.013046f
C519 B.n479 VSUBS 0.013046f
C520 B.n480 VSUBS 0.013046f
C521 B.n481 VSUBS 0.013046f
C522 B.n482 VSUBS 0.013046f
C523 B.n483 VSUBS 0.013046f
C524 B.n484 VSUBS 0.013046f
C525 B.n485 VSUBS 0.013046f
C526 B.n486 VSUBS 0.013046f
C527 B.n487 VSUBS 0.013046f
C528 B.n488 VSUBS 0.013046f
C529 B.n489 VSUBS 0.013046f
C530 B.n490 VSUBS 0.013046f
C531 B.n491 VSUBS 0.013046f
C532 B.n492 VSUBS 0.013046f
C533 B.n493 VSUBS 0.013046f
C534 B.n494 VSUBS 0.013046f
C535 B.n495 VSUBS 0.013046f
C536 B.n496 VSUBS 0.013046f
C537 B.n497 VSUBS 0.013046f
C538 B.n498 VSUBS 0.013046f
C539 B.n499 VSUBS 0.013046f
C540 B.n500 VSUBS 0.013046f
C541 B.n501 VSUBS 0.013046f
C542 B.n502 VSUBS 0.013046f
C543 B.n503 VSUBS 0.013046f
C544 B.n504 VSUBS 0.013046f
C545 B.n505 VSUBS 0.013046f
C546 B.n506 VSUBS 0.013046f
C547 B.n507 VSUBS 0.013046f
C548 B.n508 VSUBS 0.013046f
C549 B.n509 VSUBS 0.013046f
C550 B.n510 VSUBS 0.013046f
C551 B.n511 VSUBS 0.013046f
C552 B.n512 VSUBS 0.013046f
C553 B.n513 VSUBS 0.013046f
C554 B.n514 VSUBS 0.013046f
C555 B.n515 VSUBS 0.013046f
C556 B.n516 VSUBS 0.013046f
C557 B.n517 VSUBS 0.013046f
C558 B.n518 VSUBS 0.013046f
C559 B.n519 VSUBS 0.013046f
C560 B.n520 VSUBS 0.013046f
C561 B.n521 VSUBS 0.013046f
C562 B.n522 VSUBS 0.013046f
C563 B.n523 VSUBS 0.013046f
C564 B.n524 VSUBS 0.013046f
C565 B.n525 VSUBS 0.013046f
C566 B.n526 VSUBS 0.013046f
C567 B.n527 VSUBS 0.013046f
C568 B.n528 VSUBS 0.013046f
C569 B.n529 VSUBS 0.013046f
C570 B.n530 VSUBS 0.013046f
C571 B.n531 VSUBS 0.013046f
C572 B.n532 VSUBS 0.013046f
C573 B.n533 VSUBS 0.013046f
C574 B.n534 VSUBS 0.013046f
C575 B.n535 VSUBS 0.013046f
C576 B.n536 VSUBS 0.013046f
C577 B.n537 VSUBS 0.013046f
C578 B.n538 VSUBS 0.013046f
C579 B.n539 VSUBS 0.013046f
C580 B.n540 VSUBS 0.013046f
C581 B.n541 VSUBS 0.013046f
C582 B.n542 VSUBS 0.013046f
C583 B.n543 VSUBS 0.013046f
C584 B.n544 VSUBS 0.013046f
C585 B.n545 VSUBS 0.013046f
C586 B.n546 VSUBS 0.013046f
C587 B.n547 VSUBS 0.013046f
C588 B.n548 VSUBS 0.013046f
C589 B.n549 VSUBS 0.013046f
C590 B.n550 VSUBS 0.013046f
C591 B.n551 VSUBS 0.013046f
C592 B.n552 VSUBS 0.013046f
C593 B.n553 VSUBS 0.013046f
C594 B.n554 VSUBS 0.013046f
C595 B.n555 VSUBS 0.013046f
C596 B.n556 VSUBS 0.013046f
C597 B.n557 VSUBS 0.013046f
C598 B.n558 VSUBS 0.013046f
C599 B.n559 VSUBS 0.013046f
C600 B.n560 VSUBS 0.013046f
C601 B.n561 VSUBS 0.013046f
C602 B.n562 VSUBS 0.013046f
C603 B.n563 VSUBS 0.013046f
C604 B.n564 VSUBS 0.013046f
C605 B.n565 VSUBS 0.013046f
C606 B.n566 VSUBS 0.013046f
C607 B.n567 VSUBS 0.013046f
C608 B.n568 VSUBS 0.013046f
C609 B.n569 VSUBS 0.013046f
C610 B.n570 VSUBS 0.013046f
C611 B.n571 VSUBS 0.013046f
C612 B.n572 VSUBS 0.013046f
C613 B.n573 VSUBS 0.013046f
C614 B.n574 VSUBS 0.013046f
C615 B.n575 VSUBS 0.013046f
C616 B.n576 VSUBS 0.013046f
C617 B.n577 VSUBS 0.013046f
C618 B.n578 VSUBS 0.013046f
C619 B.n579 VSUBS 0.013046f
C620 B.n580 VSUBS 0.013046f
C621 B.n581 VSUBS 0.013046f
C622 B.n582 VSUBS 0.013046f
C623 B.n583 VSUBS 0.013046f
C624 B.n584 VSUBS 0.013046f
C625 B.n585 VSUBS 0.013046f
C626 B.n586 VSUBS 0.013046f
C627 B.n587 VSUBS 0.013046f
C628 B.n588 VSUBS 0.013046f
C629 B.n589 VSUBS 0.013046f
C630 B.n590 VSUBS 0.013046f
C631 B.n591 VSUBS 0.013046f
C632 B.n592 VSUBS 0.013046f
C633 B.n593 VSUBS 0.013046f
C634 B.n594 VSUBS 0.013046f
C635 B.n595 VSUBS 0.013046f
C636 B.n596 VSUBS 0.013046f
C637 B.n597 VSUBS 0.013046f
C638 B.n598 VSUBS 0.013046f
C639 B.n599 VSUBS 0.013046f
C640 B.n600 VSUBS 0.013046f
C641 B.n601 VSUBS 0.013046f
C642 B.n602 VSUBS 0.013046f
C643 B.n603 VSUBS 0.013046f
C644 B.n604 VSUBS 0.013046f
C645 B.n605 VSUBS 0.013046f
C646 B.n606 VSUBS 0.013046f
C647 B.n607 VSUBS 0.013046f
C648 B.n608 VSUBS 0.013046f
C649 B.n609 VSUBS 0.013046f
C650 B.n610 VSUBS 0.013046f
C651 B.n611 VSUBS 0.013046f
C652 B.n612 VSUBS 0.013046f
C653 B.n613 VSUBS 0.013046f
C654 B.n614 VSUBS 0.013046f
C655 B.n615 VSUBS 0.013046f
C656 B.n616 VSUBS 0.013046f
C657 B.n617 VSUBS 0.013046f
C658 B.n618 VSUBS 0.013046f
C659 B.n619 VSUBS 0.013046f
C660 B.n620 VSUBS 0.013046f
C661 B.n621 VSUBS 0.013046f
C662 B.n622 VSUBS 0.013046f
C663 B.n623 VSUBS 0.013046f
C664 B.n624 VSUBS 0.013046f
C665 B.n625 VSUBS 0.013046f
C666 B.n626 VSUBS 0.013046f
C667 B.n627 VSUBS 0.013046f
C668 B.n628 VSUBS 0.013046f
C669 B.n629 VSUBS 0.013046f
C670 B.n630 VSUBS 0.013046f
C671 B.n631 VSUBS 0.013046f
C672 B.n632 VSUBS 0.013046f
C673 B.n633 VSUBS 0.013046f
C674 B.n634 VSUBS 0.013046f
C675 B.n635 VSUBS 0.013046f
C676 B.n636 VSUBS 0.013046f
C677 B.n637 VSUBS 0.013046f
C678 B.n638 VSUBS 0.013046f
C679 B.n639 VSUBS 0.013046f
C680 B.n640 VSUBS 0.013046f
C681 B.n641 VSUBS 0.013046f
C682 B.n642 VSUBS 0.013046f
C683 B.n643 VSUBS 0.013046f
C684 B.n644 VSUBS 0.030528f
C685 B.n645 VSUBS 0.032014f
C686 B.n646 VSUBS 0.032014f
C687 B.n647 VSUBS 0.013046f
C688 B.n648 VSUBS 0.013046f
C689 B.n649 VSUBS 0.013046f
C690 B.n650 VSUBS 0.013046f
C691 B.n651 VSUBS 0.013046f
C692 B.n652 VSUBS 0.013046f
C693 B.n653 VSUBS 0.013046f
C694 B.n654 VSUBS 0.013046f
C695 B.n655 VSUBS 0.013046f
C696 B.n656 VSUBS 0.013046f
C697 B.n657 VSUBS 0.013046f
C698 B.n658 VSUBS 0.013046f
C699 B.n659 VSUBS 0.013046f
C700 B.n660 VSUBS 0.013046f
C701 B.n661 VSUBS 0.013046f
C702 B.n662 VSUBS 0.013046f
C703 B.n663 VSUBS 0.013046f
C704 B.n664 VSUBS 0.013046f
C705 B.n665 VSUBS 0.013046f
C706 B.n666 VSUBS 0.013046f
C707 B.n667 VSUBS 0.013046f
C708 B.n668 VSUBS 0.013046f
C709 B.n669 VSUBS 0.013046f
C710 B.n670 VSUBS 0.013046f
C711 B.n671 VSUBS 0.013046f
C712 B.n672 VSUBS 0.013046f
C713 B.n673 VSUBS 0.009017f
C714 B.n674 VSUBS 0.030225f
C715 B.n675 VSUBS 0.010552f
C716 B.n676 VSUBS 0.013046f
C717 B.n677 VSUBS 0.013046f
C718 B.n678 VSUBS 0.013046f
C719 B.n679 VSUBS 0.013046f
C720 B.n680 VSUBS 0.013046f
C721 B.n681 VSUBS 0.013046f
C722 B.n682 VSUBS 0.013046f
C723 B.n683 VSUBS 0.013046f
C724 B.n684 VSUBS 0.013046f
C725 B.n685 VSUBS 0.013046f
C726 B.n686 VSUBS 0.013046f
C727 B.n687 VSUBS 0.010552f
C728 B.n688 VSUBS 0.030225f
C729 B.n689 VSUBS 0.009017f
C730 B.n690 VSUBS 0.013046f
C731 B.n691 VSUBS 0.013046f
C732 B.n692 VSUBS 0.013046f
C733 B.n693 VSUBS 0.013046f
C734 B.n694 VSUBS 0.013046f
C735 B.n695 VSUBS 0.013046f
C736 B.n696 VSUBS 0.013046f
C737 B.n697 VSUBS 0.013046f
C738 B.n698 VSUBS 0.013046f
C739 B.n699 VSUBS 0.013046f
C740 B.n700 VSUBS 0.013046f
C741 B.n701 VSUBS 0.013046f
C742 B.n702 VSUBS 0.013046f
C743 B.n703 VSUBS 0.013046f
C744 B.n704 VSUBS 0.013046f
C745 B.n705 VSUBS 0.013046f
C746 B.n706 VSUBS 0.013046f
C747 B.n707 VSUBS 0.013046f
C748 B.n708 VSUBS 0.013046f
C749 B.n709 VSUBS 0.013046f
C750 B.n710 VSUBS 0.013046f
C751 B.n711 VSUBS 0.013046f
C752 B.n712 VSUBS 0.013046f
C753 B.n713 VSUBS 0.013046f
C754 B.n714 VSUBS 0.013046f
C755 B.n715 VSUBS 0.013046f
C756 B.n716 VSUBS 0.032014f
C757 B.n717 VSUBS 0.032014f
C758 B.n718 VSUBS 0.030528f
C759 B.n719 VSUBS 0.013046f
C760 B.n720 VSUBS 0.013046f
C761 B.n721 VSUBS 0.013046f
C762 B.n722 VSUBS 0.013046f
C763 B.n723 VSUBS 0.013046f
C764 B.n724 VSUBS 0.013046f
C765 B.n725 VSUBS 0.013046f
C766 B.n726 VSUBS 0.013046f
C767 B.n727 VSUBS 0.013046f
C768 B.n728 VSUBS 0.013046f
C769 B.n729 VSUBS 0.013046f
C770 B.n730 VSUBS 0.013046f
C771 B.n731 VSUBS 0.013046f
C772 B.n732 VSUBS 0.013046f
C773 B.n733 VSUBS 0.013046f
C774 B.n734 VSUBS 0.013046f
C775 B.n735 VSUBS 0.013046f
C776 B.n736 VSUBS 0.013046f
C777 B.n737 VSUBS 0.013046f
C778 B.n738 VSUBS 0.013046f
C779 B.n739 VSUBS 0.013046f
C780 B.n740 VSUBS 0.013046f
C781 B.n741 VSUBS 0.013046f
C782 B.n742 VSUBS 0.013046f
C783 B.n743 VSUBS 0.013046f
C784 B.n744 VSUBS 0.013046f
C785 B.n745 VSUBS 0.013046f
C786 B.n746 VSUBS 0.013046f
C787 B.n747 VSUBS 0.013046f
C788 B.n748 VSUBS 0.013046f
C789 B.n749 VSUBS 0.013046f
C790 B.n750 VSUBS 0.013046f
C791 B.n751 VSUBS 0.013046f
C792 B.n752 VSUBS 0.013046f
C793 B.n753 VSUBS 0.013046f
C794 B.n754 VSUBS 0.013046f
C795 B.n755 VSUBS 0.013046f
C796 B.n756 VSUBS 0.013046f
C797 B.n757 VSUBS 0.013046f
C798 B.n758 VSUBS 0.013046f
C799 B.n759 VSUBS 0.013046f
C800 B.n760 VSUBS 0.013046f
C801 B.n761 VSUBS 0.013046f
C802 B.n762 VSUBS 0.013046f
C803 B.n763 VSUBS 0.013046f
C804 B.n764 VSUBS 0.013046f
C805 B.n765 VSUBS 0.013046f
C806 B.n766 VSUBS 0.013046f
C807 B.n767 VSUBS 0.013046f
C808 B.n768 VSUBS 0.013046f
C809 B.n769 VSUBS 0.013046f
C810 B.n770 VSUBS 0.013046f
C811 B.n771 VSUBS 0.013046f
C812 B.n772 VSUBS 0.013046f
C813 B.n773 VSUBS 0.013046f
C814 B.n774 VSUBS 0.013046f
C815 B.n775 VSUBS 0.013046f
C816 B.n776 VSUBS 0.013046f
C817 B.n777 VSUBS 0.013046f
C818 B.n778 VSUBS 0.013046f
C819 B.n779 VSUBS 0.013046f
C820 B.n780 VSUBS 0.013046f
C821 B.n781 VSUBS 0.013046f
C822 B.n782 VSUBS 0.013046f
C823 B.n783 VSUBS 0.013046f
C824 B.n784 VSUBS 0.013046f
C825 B.n785 VSUBS 0.013046f
C826 B.n786 VSUBS 0.013046f
C827 B.n787 VSUBS 0.013046f
C828 B.n788 VSUBS 0.013046f
C829 B.n789 VSUBS 0.013046f
C830 B.n790 VSUBS 0.013046f
C831 B.n791 VSUBS 0.013046f
C832 B.n792 VSUBS 0.013046f
C833 B.n793 VSUBS 0.013046f
C834 B.n794 VSUBS 0.013046f
C835 B.n795 VSUBS 0.013046f
C836 B.n796 VSUBS 0.013046f
C837 B.n797 VSUBS 0.013046f
C838 B.n798 VSUBS 0.013046f
C839 B.n799 VSUBS 0.013046f
C840 B.n800 VSUBS 0.013046f
C841 B.n801 VSUBS 0.013046f
C842 B.n802 VSUBS 0.013046f
C843 B.n803 VSUBS 0.013046f
C844 B.n804 VSUBS 0.013046f
C845 B.n805 VSUBS 0.013046f
C846 B.n806 VSUBS 0.013046f
C847 B.n807 VSUBS 0.013046f
C848 B.n808 VSUBS 0.013046f
C849 B.n809 VSUBS 0.013046f
C850 B.n810 VSUBS 0.013046f
C851 B.n811 VSUBS 0.013046f
C852 B.n812 VSUBS 0.013046f
C853 B.n813 VSUBS 0.013046f
C854 B.n814 VSUBS 0.013046f
C855 B.n815 VSUBS 0.013046f
C856 B.n816 VSUBS 0.013046f
C857 B.n817 VSUBS 0.013046f
C858 B.n818 VSUBS 0.013046f
C859 B.n819 VSUBS 0.013046f
C860 B.n820 VSUBS 0.013046f
C861 B.n821 VSUBS 0.013046f
C862 B.n822 VSUBS 0.013046f
C863 B.n823 VSUBS 0.013046f
C864 B.n824 VSUBS 0.013046f
C865 B.n825 VSUBS 0.013046f
C866 B.n826 VSUBS 0.013046f
C867 B.n827 VSUBS 0.013046f
C868 B.n828 VSUBS 0.013046f
C869 B.n829 VSUBS 0.013046f
C870 B.n830 VSUBS 0.013046f
C871 B.n831 VSUBS 0.013046f
C872 B.n832 VSUBS 0.013046f
C873 B.n833 VSUBS 0.013046f
C874 B.n834 VSUBS 0.013046f
C875 B.n835 VSUBS 0.017024f
C876 B.n836 VSUBS 0.018135f
C877 B.n837 VSUBS 0.036062f
C878 VDD1.t0 VSUBS 1.06602f
C879 VDD1.t8 VSUBS 0.126606f
C880 VDD1.t3 VSUBS 0.126606f
C881 VDD1.n0 VSUBS 0.754248f
C882 VDD1.n1 VSUBS 2.1082f
C883 VDD1.t9 VSUBS 1.06602f
C884 VDD1.t7 VSUBS 0.126606f
C885 VDD1.t6 VSUBS 0.126606f
C886 VDD1.n2 VSUBS 0.754245f
C887 VDD1.n3 VSUBS 2.09542f
C888 VDD1.t4 VSUBS 0.126606f
C889 VDD1.t5 VSUBS 0.126606f
C890 VDD1.n4 VSUBS 0.784152f
C891 VDD1.n5 VSUBS 5.03444f
C892 VDD1.t2 VSUBS 0.126606f
C893 VDD1.t1 VSUBS 0.126606f
C894 VDD1.n6 VSUBS 0.754244f
C895 VDD1.n7 VSUBS 4.84405f
C896 VP.t4 VSUBS 1.6417f
C897 VP.n0 VSUBS 0.784225f
C898 VP.n1 VSUBS 0.040413f
C899 VP.n2 VSUBS 0.076045f
C900 VP.n3 VSUBS 0.040413f
C901 VP.n4 VSUBS 0.071601f
C902 VP.n5 VSUBS 0.040413f
C903 VP.n6 VSUBS 0.079156f
C904 VP.n7 VSUBS 0.040413f
C905 VP.n8 VSUBS 0.075319f
C906 VP.n9 VSUBS 0.040413f
C907 VP.t3 VSUBS 1.6417f
C908 VP.n10 VSUBS 0.081164f
C909 VP.n11 VSUBS 0.040413f
C910 VP.n12 VSUBS 0.075319f
C911 VP.n13 VSUBS 0.040413f
C912 VP.t2 VSUBS 1.6417f
C913 VP.n14 VSUBS 0.081584f
C914 VP.n15 VSUBS 0.040413f
C915 VP.n16 VSUBS 0.075319f
C916 VP.t8 VSUBS 1.6417f
C917 VP.n17 VSUBS 0.784225f
C918 VP.n18 VSUBS 0.040413f
C919 VP.n19 VSUBS 0.076045f
C920 VP.n20 VSUBS 0.040413f
C921 VP.n21 VSUBS 0.071601f
C922 VP.n22 VSUBS 0.040413f
C923 VP.n23 VSUBS 0.079156f
C924 VP.n24 VSUBS 0.040413f
C925 VP.n25 VSUBS 0.075319f
C926 VP.n26 VSUBS 0.040413f
C927 VP.t6 VSUBS 1.6417f
C928 VP.n27 VSUBS 0.081164f
C929 VP.n28 VSUBS 0.040413f
C930 VP.n29 VSUBS 0.075319f
C931 VP.t9 VSUBS 2.15116f
C932 VP.n30 VSUBS 0.759891f
C933 VP.t1 VSUBS 1.6417f
C934 VP.n31 VSUBS 0.761132f
C935 VP.n32 VSUBS 0.041852f
C936 VP.n33 VSUBS 0.513604f
C937 VP.n34 VSUBS 0.040413f
C938 VP.n35 VSUBS 0.040413f
C939 VP.n36 VSUBS 0.075319f
C940 VP.n37 VSUBS 0.079156f
C941 VP.n38 VSUBS 0.032997f
C942 VP.n39 VSUBS 0.040413f
C943 VP.n40 VSUBS 0.040413f
C944 VP.n41 VSUBS 0.040413f
C945 VP.n42 VSUBS 0.075319f
C946 VP.n43 VSUBS 0.075319f
C947 VP.n44 VSUBS 0.669365f
C948 VP.n45 VSUBS 0.040413f
C949 VP.n46 VSUBS 0.040413f
C950 VP.n47 VSUBS 0.040413f
C951 VP.n48 VSUBS 0.075319f
C952 VP.n49 VSUBS 0.081164f
C953 VP.n50 VSUBS 0.032997f
C954 VP.n51 VSUBS 0.040413f
C955 VP.n52 VSUBS 0.040413f
C956 VP.n53 VSUBS 0.040413f
C957 VP.n54 VSUBS 0.075319f
C958 VP.n55 VSUBS 0.075319f
C959 VP.t7 VSUBS 1.6417f
C960 VP.n56 VSUBS 0.631231f
C961 VP.n57 VSUBS 0.041852f
C962 VP.n58 VSUBS 0.040413f
C963 VP.n59 VSUBS 0.040413f
C964 VP.n60 VSUBS 0.040413f
C965 VP.n61 VSUBS 0.075319f
C966 VP.n62 VSUBS 0.081584f
C967 VP.n63 VSUBS 0.035689f
C968 VP.n64 VSUBS 0.040413f
C969 VP.n65 VSUBS 0.040413f
C970 VP.n66 VSUBS 0.040413f
C971 VP.n67 VSUBS 0.075319f
C972 VP.n68 VSUBS 0.075319f
C973 VP.n69 VSUBS 0.045571f
C974 VP.n70 VSUBS 0.065225f
C975 VP.n71 VSUBS 2.54493f
C976 VP.n72 VSUBS 2.57214f
C977 VP.t0 VSUBS 1.6417f
C978 VP.n73 VSUBS 0.784225f
C979 VP.n74 VSUBS 0.045571f
C980 VP.n75 VSUBS 0.065225f
C981 VP.n76 VSUBS 0.040413f
C982 VP.n77 VSUBS 0.040413f
C983 VP.n78 VSUBS 0.075319f
C984 VP.n79 VSUBS 0.076045f
C985 VP.n80 VSUBS 0.035689f
C986 VP.n81 VSUBS 0.040413f
C987 VP.n82 VSUBS 0.040413f
C988 VP.n83 VSUBS 0.040413f
C989 VP.n84 VSUBS 0.075319f
C990 VP.n85 VSUBS 0.071601f
C991 VP.n86 VSUBS 0.631231f
C992 VP.n87 VSUBS 0.041852f
C993 VP.n88 VSUBS 0.040413f
C994 VP.n89 VSUBS 0.040413f
C995 VP.n90 VSUBS 0.040413f
C996 VP.n91 VSUBS 0.075319f
C997 VP.n92 VSUBS 0.079156f
C998 VP.n93 VSUBS 0.032997f
C999 VP.n94 VSUBS 0.040413f
C1000 VP.n95 VSUBS 0.040413f
C1001 VP.n96 VSUBS 0.040413f
C1002 VP.n97 VSUBS 0.075319f
C1003 VP.n98 VSUBS 0.075319f
C1004 VP.n99 VSUBS 0.669365f
C1005 VP.n100 VSUBS 0.040413f
C1006 VP.n101 VSUBS 0.040413f
C1007 VP.n102 VSUBS 0.040413f
C1008 VP.n103 VSUBS 0.075319f
C1009 VP.n104 VSUBS 0.081164f
C1010 VP.n105 VSUBS 0.032997f
C1011 VP.n106 VSUBS 0.040413f
C1012 VP.n107 VSUBS 0.040413f
C1013 VP.n108 VSUBS 0.040413f
C1014 VP.n109 VSUBS 0.075319f
C1015 VP.n110 VSUBS 0.075319f
C1016 VP.t5 VSUBS 1.6417f
C1017 VP.n111 VSUBS 0.631231f
C1018 VP.n112 VSUBS 0.041852f
C1019 VP.n113 VSUBS 0.040413f
C1020 VP.n114 VSUBS 0.040413f
C1021 VP.n115 VSUBS 0.040413f
C1022 VP.n116 VSUBS 0.075319f
C1023 VP.n117 VSUBS 0.081584f
C1024 VP.n118 VSUBS 0.035689f
C1025 VP.n119 VSUBS 0.040413f
C1026 VP.n120 VSUBS 0.040413f
C1027 VP.n121 VSUBS 0.040413f
C1028 VP.n122 VSUBS 0.075319f
C1029 VP.n123 VSUBS 0.075319f
C1030 VP.n124 VSUBS 0.045571f
C1031 VP.n125 VSUBS 0.065225f
C1032 VP.n126 VSUBS 0.119916f
C1033 VDD2.t0 VSUBS 1.06809f
C1034 VDD2.t1 VSUBS 0.126852f
C1035 VDD2.t7 VSUBS 0.126852f
C1036 VDD2.n0 VSUBS 0.755709f
C1037 VDD2.n1 VSUBS 2.09949f
C1038 VDD2.t8 VSUBS 0.126852f
C1039 VDD2.t9 VSUBS 0.126852f
C1040 VDD2.n2 VSUBS 0.785674f
C1041 VDD2.n3 VSUBS 4.81893f
C1042 VDD2.t3 VSUBS 1.03745f
C1043 VDD2.n4 VSUBS 4.68969f
C1044 VDD2.t5 VSUBS 0.126852f
C1045 VDD2.t6 VSUBS 0.126852f
C1046 VDD2.n5 VSUBS 0.755712f
C1047 VDD2.n6 VSUBS 1.08864f
C1048 VDD2.t2 VSUBS 0.126852f
C1049 VDD2.t4 VSUBS 0.126852f
C1050 VDD2.n7 VSUBS 0.785625f
C1051 VTAIL.t8 VSUBS 0.127397f
C1052 VTAIL.t14 VSUBS 0.127397f
C1053 VTAIL.n0 VSUBS 0.660833f
C1054 VTAIL.n1 VSUBS 1.19735f
C1055 VTAIL.t19 VSUBS 0.940572f
C1056 VTAIL.n2 VSUBS 1.3651f
C1057 VTAIL.t1 VSUBS 0.127397f
C1058 VTAIL.t4 VSUBS 0.127397f
C1059 VTAIL.n3 VSUBS 0.660833f
C1060 VTAIL.n4 VSUBS 1.45408f
C1061 VTAIL.t5 VSUBS 0.127397f
C1062 VTAIL.t7 VSUBS 0.127397f
C1063 VTAIL.n5 VSUBS 0.660833f
C1064 VTAIL.n6 VSUBS 2.84837f
C1065 VTAIL.t10 VSUBS 0.127397f
C1066 VTAIL.t9 VSUBS 0.127397f
C1067 VTAIL.n7 VSUBS 0.660837f
C1068 VTAIL.n8 VSUBS 2.84837f
C1069 VTAIL.t16 VSUBS 0.127397f
C1070 VTAIL.t13 VSUBS 0.127397f
C1071 VTAIL.n9 VSUBS 0.660837f
C1072 VTAIL.n10 VSUBS 1.45407f
C1073 VTAIL.t12 VSUBS 0.940576f
C1074 VTAIL.n11 VSUBS 1.3651f
C1075 VTAIL.t0 VSUBS 0.127397f
C1076 VTAIL.t18 VSUBS 0.127397f
C1077 VTAIL.n12 VSUBS 0.660837f
C1078 VTAIL.n13 VSUBS 1.29739f
C1079 VTAIL.t6 VSUBS 0.127397f
C1080 VTAIL.t3 VSUBS 0.127397f
C1081 VTAIL.n14 VSUBS 0.660837f
C1082 VTAIL.n15 VSUBS 1.45407f
C1083 VTAIL.t2 VSUBS 0.940572f
C1084 VTAIL.n16 VSUBS 2.48732f
C1085 VTAIL.t17 VSUBS 0.940572f
C1086 VTAIL.n17 VSUBS 2.48732f
C1087 VTAIL.t15 VSUBS 0.127397f
C1088 VTAIL.t11 VSUBS 0.127397f
C1089 VTAIL.n18 VSUBS 0.660833f
C1090 VTAIL.n19 VSUBS 1.12536f
C1091 VN.t0 VSUBS 1.45244f
C1092 VN.n0 VSUBS 0.693816f
C1093 VN.n1 VSUBS 0.035754f
C1094 VN.n2 VSUBS 0.067278f
C1095 VN.n3 VSUBS 0.035754f
C1096 VN.n4 VSUBS 0.063346f
C1097 VN.n5 VSUBS 0.035754f
C1098 VN.n6 VSUBS 0.070031f
C1099 VN.n7 VSUBS 0.035754f
C1100 VN.n8 VSUBS 0.066636f
C1101 VN.n9 VSUBS 0.035754f
C1102 VN.t2 VSUBS 1.45244f
C1103 VN.n10 VSUBS 0.071807f
C1104 VN.n11 VSUBS 0.035754f
C1105 VN.n12 VSUBS 0.066636f
C1106 VN.t9 VSUBS 1.90316f
C1107 VN.n13 VSUBS 0.672286f
C1108 VN.t8 VSUBS 1.45244f
C1109 VN.n14 VSUBS 0.673385f
C1110 VN.n15 VSUBS 0.037027f
C1111 VN.n16 VSUBS 0.454393f
C1112 VN.n17 VSUBS 0.035754f
C1113 VN.n18 VSUBS 0.035754f
C1114 VN.n19 VSUBS 0.066636f
C1115 VN.n20 VSUBS 0.070031f
C1116 VN.n21 VSUBS 0.029193f
C1117 VN.n22 VSUBS 0.035754f
C1118 VN.n23 VSUBS 0.035754f
C1119 VN.n24 VSUBS 0.035754f
C1120 VN.n25 VSUBS 0.066636f
C1121 VN.n26 VSUBS 0.066636f
C1122 VN.n27 VSUBS 0.592197f
C1123 VN.n28 VSUBS 0.035754f
C1124 VN.n29 VSUBS 0.035754f
C1125 VN.n30 VSUBS 0.035754f
C1126 VN.n31 VSUBS 0.066636f
C1127 VN.n32 VSUBS 0.071807f
C1128 VN.n33 VSUBS 0.029193f
C1129 VN.n34 VSUBS 0.035754f
C1130 VN.n35 VSUBS 0.035754f
C1131 VN.n36 VSUBS 0.035754f
C1132 VN.n37 VSUBS 0.066636f
C1133 VN.n38 VSUBS 0.066636f
C1134 VN.t1 VSUBS 1.45244f
C1135 VN.n39 VSUBS 0.55846f
C1136 VN.n40 VSUBS 0.037027f
C1137 VN.n41 VSUBS 0.035754f
C1138 VN.n42 VSUBS 0.035754f
C1139 VN.n43 VSUBS 0.035754f
C1140 VN.n44 VSUBS 0.066636f
C1141 VN.n45 VSUBS 0.072178f
C1142 VN.n46 VSUBS 0.031574f
C1143 VN.n47 VSUBS 0.035754f
C1144 VN.n48 VSUBS 0.035754f
C1145 VN.n49 VSUBS 0.035754f
C1146 VN.n50 VSUBS 0.066636f
C1147 VN.n51 VSUBS 0.066636f
C1148 VN.n52 VSUBS 0.040317f
C1149 VN.n53 VSUBS 0.057706f
C1150 VN.n54 VSUBS 0.106091f
C1151 VN.t6 VSUBS 1.45244f
C1152 VN.n55 VSUBS 0.693816f
C1153 VN.n56 VSUBS 0.035754f
C1154 VN.n57 VSUBS 0.067278f
C1155 VN.n58 VSUBS 0.035754f
C1156 VN.n59 VSUBS 0.063346f
C1157 VN.n60 VSUBS 0.035754f
C1158 VN.t4 VSUBS 1.45244f
C1159 VN.n61 VSUBS 0.55846f
C1160 VN.n62 VSUBS 0.070031f
C1161 VN.n63 VSUBS 0.035754f
C1162 VN.n64 VSUBS 0.066636f
C1163 VN.n65 VSUBS 0.035754f
C1164 VN.t3 VSUBS 1.45244f
C1165 VN.n66 VSUBS 0.071807f
C1166 VN.n67 VSUBS 0.035754f
C1167 VN.n68 VSUBS 0.066636f
C1168 VN.t5 VSUBS 1.90316f
C1169 VN.n69 VSUBS 0.672286f
C1170 VN.t7 VSUBS 1.45244f
C1171 VN.n70 VSUBS 0.673385f
C1172 VN.n71 VSUBS 0.037027f
C1173 VN.n72 VSUBS 0.454392f
C1174 VN.n73 VSUBS 0.035754f
C1175 VN.n74 VSUBS 0.035754f
C1176 VN.n75 VSUBS 0.066636f
C1177 VN.n76 VSUBS 0.070031f
C1178 VN.n77 VSUBS 0.029193f
C1179 VN.n78 VSUBS 0.035754f
C1180 VN.n79 VSUBS 0.035754f
C1181 VN.n80 VSUBS 0.035754f
C1182 VN.n81 VSUBS 0.066636f
C1183 VN.n82 VSUBS 0.066636f
C1184 VN.n83 VSUBS 0.592197f
C1185 VN.n84 VSUBS 0.035754f
C1186 VN.n85 VSUBS 0.035754f
C1187 VN.n86 VSUBS 0.035754f
C1188 VN.n87 VSUBS 0.066636f
C1189 VN.n88 VSUBS 0.071807f
C1190 VN.n89 VSUBS 0.029193f
C1191 VN.n90 VSUBS 0.035754f
C1192 VN.n91 VSUBS 0.035754f
C1193 VN.n92 VSUBS 0.035754f
C1194 VN.n93 VSUBS 0.066636f
C1195 VN.n94 VSUBS 0.066636f
C1196 VN.n95 VSUBS 0.037027f
C1197 VN.n96 VSUBS 0.035754f
C1198 VN.n97 VSUBS 0.035754f
C1199 VN.n98 VSUBS 0.035754f
C1200 VN.n99 VSUBS 0.066636f
C1201 VN.n100 VSUBS 0.072178f
C1202 VN.n101 VSUBS 0.031574f
C1203 VN.n102 VSUBS 0.035754f
C1204 VN.n103 VSUBS 0.035754f
C1205 VN.n104 VSUBS 0.035754f
C1206 VN.n105 VSUBS 0.066636f
C1207 VN.n106 VSUBS 0.066636f
C1208 VN.n107 VSUBS 0.040317f
C1209 VN.n108 VSUBS 0.057706f
C1210 VN.n109 VSUBS 2.26584f
.ends

