* NGSPICE file created from diff_pair_sample_0571.ext - technology: sky130A

.subckt diff_pair_sample_0571 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t3 VP.t0 VTAIL.t4 B.t1 sky130_fd_pr__nfet_01v8 ad=0.3861 pd=2.67 as=0.9126 ps=5.46 w=2.34 l=1.98
X1 VTAIL.t5 VP.t1 VDD1.t2 B.t0 sky130_fd_pr__nfet_01v8 ad=0.9126 pd=5.46 as=0.3861 ps=2.67 w=2.34 l=1.98
X2 B.t17 B.t15 B.t16 B.t5 sky130_fd_pr__nfet_01v8 ad=0.9126 pd=5.46 as=0 ps=0 w=2.34 l=1.98
X3 B.t14 B.t12 B.t13 B.t9 sky130_fd_pr__nfet_01v8 ad=0.9126 pd=5.46 as=0 ps=0 w=2.34 l=1.98
X4 VTAIL.t0 VN.t0 VDD2.t3 B.t0 sky130_fd_pr__nfet_01v8 ad=0.9126 pd=5.46 as=0.3861 ps=2.67 w=2.34 l=1.98
X5 VDD2.t2 VN.t1 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=0.3861 pd=2.67 as=0.9126 ps=5.46 w=2.34 l=1.98
X6 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=0.9126 pd=5.46 as=0 ps=0 w=2.34 l=1.98
X7 VTAIL.t7 VP.t2 VDD1.t1 B.t3 sky130_fd_pr__nfet_01v8 ad=0.9126 pd=5.46 as=0.3861 ps=2.67 w=2.34 l=1.98
X8 VDD2.t1 VN.t2 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=0.3861 pd=2.67 as=0.9126 ps=5.46 w=2.34 l=1.98
X9 B.t7 B.t4 B.t6 B.t5 sky130_fd_pr__nfet_01v8 ad=0.9126 pd=5.46 as=0 ps=0 w=2.34 l=1.98
X10 VTAIL.t3 VN.t3 VDD2.t0 B.t3 sky130_fd_pr__nfet_01v8 ad=0.9126 pd=5.46 as=0.3861 ps=2.67 w=2.34 l=1.98
X11 VDD1.t0 VP.t3 VTAIL.t6 B.t2 sky130_fd_pr__nfet_01v8 ad=0.3861 pd=2.67 as=0.9126 ps=5.46 w=2.34 l=1.98
R0 VP.n10 VP.n0 161.3
R1 VP.n9 VP.n8 161.3
R2 VP.n7 VP.n1 161.3
R3 VP.n6 VP.n5 161.3
R4 VP.n4 VP.n3 90.9889
R5 VP.n12 VP.n11 90.9889
R6 VP.n2 VP.t2 64.0351
R7 VP.n2 VP.t0 63.5056
R8 VP.n9 VP.n1 56.5617
R9 VP.n3 VP.n2 44.3789
R10 VP.n4 VP.t1 28.4823
R11 VP.n11 VP.t3 28.4823
R12 VP.n5 VP.n1 24.5923
R13 VP.n10 VP.n9 24.5923
R14 VP.n5 VP.n4 19.9199
R15 VP.n11 VP.n10 19.9199
R16 VP.n6 VP.n3 0.278335
R17 VP.n12 VP.n0 0.278335
R18 VP.n7 VP.n6 0.189894
R19 VP.n8 VP.n7 0.189894
R20 VP.n8 VP.n0 0.189894
R21 VP VP.n12 0.153485
R22 VTAIL.n5 VTAIL.t7 83.0938
R23 VTAIL.n4 VTAIL.t2 83.0938
R24 VTAIL.n3 VTAIL.t0 83.0938
R25 VTAIL.n6 VTAIL.t4 83.0938
R26 VTAIL.n7 VTAIL.t1 83.0937
R27 VTAIL.n0 VTAIL.t3 83.0937
R28 VTAIL.n1 VTAIL.t6 83.0937
R29 VTAIL.n2 VTAIL.t5 83.0937
R30 VTAIL.n7 VTAIL.n6 16.3755
R31 VTAIL.n3 VTAIL.n2 16.3755
R32 VTAIL.n4 VTAIL.n3 1.99188
R33 VTAIL.n6 VTAIL.n5 1.99188
R34 VTAIL.n2 VTAIL.n1 1.99188
R35 VTAIL VTAIL.n0 1.05438
R36 VTAIL VTAIL.n7 0.938
R37 VTAIL.n5 VTAIL.n4 0.470328
R38 VTAIL.n1 VTAIL.n0 0.470328
R39 VDD1 VDD1.n1 123.541
R40 VDD1 VDD1.n0 91.3692
R41 VDD1.n0 VDD1.t1 8.46204
R42 VDD1.n0 VDD1.t3 8.46204
R43 VDD1.n1 VDD1.t2 8.46204
R44 VDD1.n1 VDD1.t0 8.46204
R45 B.n419 B.n418 585
R46 B.n146 B.n73 585
R47 B.n145 B.n144 585
R48 B.n143 B.n142 585
R49 B.n141 B.n140 585
R50 B.n139 B.n138 585
R51 B.n137 B.n136 585
R52 B.n135 B.n134 585
R53 B.n133 B.n132 585
R54 B.n131 B.n130 585
R55 B.n129 B.n128 585
R56 B.n127 B.n126 585
R57 B.n125 B.n124 585
R58 B.n122 B.n121 585
R59 B.n120 B.n119 585
R60 B.n118 B.n117 585
R61 B.n116 B.n115 585
R62 B.n114 B.n113 585
R63 B.n112 B.n111 585
R64 B.n110 B.n109 585
R65 B.n108 B.n107 585
R66 B.n106 B.n105 585
R67 B.n104 B.n103 585
R68 B.n101 B.n100 585
R69 B.n99 B.n98 585
R70 B.n97 B.n96 585
R71 B.n95 B.n94 585
R72 B.n93 B.n92 585
R73 B.n91 B.n90 585
R74 B.n89 B.n88 585
R75 B.n87 B.n86 585
R76 B.n85 B.n84 585
R77 B.n83 B.n82 585
R78 B.n81 B.n80 585
R79 B.n79 B.n78 585
R80 B.n54 B.n53 585
R81 B.n417 B.n55 585
R82 B.n422 B.n55 585
R83 B.n416 B.n415 585
R84 B.n415 B.n51 585
R85 B.n414 B.n50 585
R86 B.n428 B.n50 585
R87 B.n413 B.n49 585
R88 B.n429 B.n49 585
R89 B.n412 B.n48 585
R90 B.n430 B.n48 585
R91 B.n411 B.n410 585
R92 B.n410 B.n44 585
R93 B.n409 B.n43 585
R94 B.n436 B.n43 585
R95 B.n408 B.n42 585
R96 B.n437 B.n42 585
R97 B.n407 B.n41 585
R98 B.n438 B.n41 585
R99 B.n406 B.n405 585
R100 B.n405 B.n37 585
R101 B.n404 B.n36 585
R102 B.n444 B.n36 585
R103 B.n403 B.n35 585
R104 B.n445 B.n35 585
R105 B.n402 B.n34 585
R106 B.n446 B.n34 585
R107 B.n401 B.n400 585
R108 B.n400 B.n30 585
R109 B.n399 B.n29 585
R110 B.n452 B.n29 585
R111 B.n398 B.n28 585
R112 B.n453 B.n28 585
R113 B.n397 B.n27 585
R114 B.n454 B.n27 585
R115 B.n396 B.n395 585
R116 B.n395 B.n23 585
R117 B.n394 B.n22 585
R118 B.n460 B.n22 585
R119 B.n393 B.n21 585
R120 B.n461 B.n21 585
R121 B.n392 B.n20 585
R122 B.n462 B.n20 585
R123 B.n391 B.n390 585
R124 B.n390 B.n16 585
R125 B.n389 B.n15 585
R126 B.n468 B.n15 585
R127 B.n388 B.n14 585
R128 B.n469 B.n14 585
R129 B.n387 B.n13 585
R130 B.n470 B.n13 585
R131 B.n386 B.n385 585
R132 B.n385 B.n12 585
R133 B.n384 B.n383 585
R134 B.n384 B.n8 585
R135 B.n382 B.n7 585
R136 B.n477 B.n7 585
R137 B.n381 B.n6 585
R138 B.n478 B.n6 585
R139 B.n380 B.n5 585
R140 B.n479 B.n5 585
R141 B.n379 B.n378 585
R142 B.n378 B.n4 585
R143 B.n377 B.n147 585
R144 B.n377 B.n376 585
R145 B.n367 B.n148 585
R146 B.n149 B.n148 585
R147 B.n369 B.n368 585
R148 B.n370 B.n369 585
R149 B.n366 B.n153 585
R150 B.n157 B.n153 585
R151 B.n365 B.n364 585
R152 B.n364 B.n363 585
R153 B.n155 B.n154 585
R154 B.n156 B.n155 585
R155 B.n356 B.n355 585
R156 B.n357 B.n356 585
R157 B.n354 B.n162 585
R158 B.n162 B.n161 585
R159 B.n353 B.n352 585
R160 B.n352 B.n351 585
R161 B.n164 B.n163 585
R162 B.n165 B.n164 585
R163 B.n344 B.n343 585
R164 B.n345 B.n344 585
R165 B.n342 B.n170 585
R166 B.n170 B.n169 585
R167 B.n341 B.n340 585
R168 B.n340 B.n339 585
R169 B.n172 B.n171 585
R170 B.n173 B.n172 585
R171 B.n332 B.n331 585
R172 B.n333 B.n332 585
R173 B.n330 B.n178 585
R174 B.n178 B.n177 585
R175 B.n329 B.n328 585
R176 B.n328 B.n327 585
R177 B.n180 B.n179 585
R178 B.n181 B.n180 585
R179 B.n320 B.n319 585
R180 B.n321 B.n320 585
R181 B.n318 B.n186 585
R182 B.n186 B.n185 585
R183 B.n317 B.n316 585
R184 B.n316 B.n315 585
R185 B.n188 B.n187 585
R186 B.n189 B.n188 585
R187 B.n308 B.n307 585
R188 B.n309 B.n308 585
R189 B.n306 B.n194 585
R190 B.n194 B.n193 585
R191 B.n305 B.n304 585
R192 B.n304 B.n303 585
R193 B.n196 B.n195 585
R194 B.n197 B.n196 585
R195 B.n296 B.n295 585
R196 B.n297 B.n296 585
R197 B.n200 B.n199 585
R198 B.n227 B.n226 585
R199 B.n228 B.n224 585
R200 B.n224 B.n201 585
R201 B.n230 B.n229 585
R202 B.n232 B.n223 585
R203 B.n235 B.n234 585
R204 B.n236 B.n222 585
R205 B.n238 B.n237 585
R206 B.n240 B.n221 585
R207 B.n243 B.n242 585
R208 B.n244 B.n220 585
R209 B.n246 B.n245 585
R210 B.n248 B.n219 585
R211 B.n251 B.n250 585
R212 B.n252 B.n215 585
R213 B.n254 B.n253 585
R214 B.n256 B.n214 585
R215 B.n259 B.n258 585
R216 B.n260 B.n213 585
R217 B.n262 B.n261 585
R218 B.n264 B.n212 585
R219 B.n267 B.n266 585
R220 B.n268 B.n209 585
R221 B.n271 B.n270 585
R222 B.n273 B.n208 585
R223 B.n276 B.n275 585
R224 B.n277 B.n207 585
R225 B.n279 B.n278 585
R226 B.n281 B.n206 585
R227 B.n284 B.n283 585
R228 B.n285 B.n205 585
R229 B.n287 B.n286 585
R230 B.n289 B.n204 585
R231 B.n290 B.n203 585
R232 B.n293 B.n292 585
R233 B.n294 B.n202 585
R234 B.n202 B.n201 585
R235 B.n299 B.n298 585
R236 B.n298 B.n297 585
R237 B.n300 B.n198 585
R238 B.n198 B.n197 585
R239 B.n302 B.n301 585
R240 B.n303 B.n302 585
R241 B.n192 B.n191 585
R242 B.n193 B.n192 585
R243 B.n311 B.n310 585
R244 B.n310 B.n309 585
R245 B.n312 B.n190 585
R246 B.n190 B.n189 585
R247 B.n314 B.n313 585
R248 B.n315 B.n314 585
R249 B.n184 B.n183 585
R250 B.n185 B.n184 585
R251 B.n323 B.n322 585
R252 B.n322 B.n321 585
R253 B.n324 B.n182 585
R254 B.n182 B.n181 585
R255 B.n326 B.n325 585
R256 B.n327 B.n326 585
R257 B.n176 B.n175 585
R258 B.n177 B.n176 585
R259 B.n335 B.n334 585
R260 B.n334 B.n333 585
R261 B.n336 B.n174 585
R262 B.n174 B.n173 585
R263 B.n338 B.n337 585
R264 B.n339 B.n338 585
R265 B.n168 B.n167 585
R266 B.n169 B.n168 585
R267 B.n347 B.n346 585
R268 B.n346 B.n345 585
R269 B.n348 B.n166 585
R270 B.n166 B.n165 585
R271 B.n350 B.n349 585
R272 B.n351 B.n350 585
R273 B.n160 B.n159 585
R274 B.n161 B.n160 585
R275 B.n359 B.n358 585
R276 B.n358 B.n357 585
R277 B.n360 B.n158 585
R278 B.n158 B.n156 585
R279 B.n362 B.n361 585
R280 B.n363 B.n362 585
R281 B.n152 B.n151 585
R282 B.n157 B.n152 585
R283 B.n372 B.n371 585
R284 B.n371 B.n370 585
R285 B.n373 B.n150 585
R286 B.n150 B.n149 585
R287 B.n375 B.n374 585
R288 B.n376 B.n375 585
R289 B.n3 B.n0 585
R290 B.n4 B.n3 585
R291 B.n476 B.n1 585
R292 B.n477 B.n476 585
R293 B.n475 B.n474 585
R294 B.n475 B.n8 585
R295 B.n473 B.n9 585
R296 B.n12 B.n9 585
R297 B.n472 B.n471 585
R298 B.n471 B.n470 585
R299 B.n11 B.n10 585
R300 B.n469 B.n11 585
R301 B.n467 B.n466 585
R302 B.n468 B.n467 585
R303 B.n465 B.n17 585
R304 B.n17 B.n16 585
R305 B.n464 B.n463 585
R306 B.n463 B.n462 585
R307 B.n19 B.n18 585
R308 B.n461 B.n19 585
R309 B.n459 B.n458 585
R310 B.n460 B.n459 585
R311 B.n457 B.n24 585
R312 B.n24 B.n23 585
R313 B.n456 B.n455 585
R314 B.n455 B.n454 585
R315 B.n26 B.n25 585
R316 B.n453 B.n26 585
R317 B.n451 B.n450 585
R318 B.n452 B.n451 585
R319 B.n449 B.n31 585
R320 B.n31 B.n30 585
R321 B.n448 B.n447 585
R322 B.n447 B.n446 585
R323 B.n33 B.n32 585
R324 B.n445 B.n33 585
R325 B.n443 B.n442 585
R326 B.n444 B.n443 585
R327 B.n441 B.n38 585
R328 B.n38 B.n37 585
R329 B.n440 B.n439 585
R330 B.n439 B.n438 585
R331 B.n40 B.n39 585
R332 B.n437 B.n40 585
R333 B.n435 B.n434 585
R334 B.n436 B.n435 585
R335 B.n433 B.n45 585
R336 B.n45 B.n44 585
R337 B.n432 B.n431 585
R338 B.n431 B.n430 585
R339 B.n47 B.n46 585
R340 B.n429 B.n47 585
R341 B.n427 B.n426 585
R342 B.n428 B.n427 585
R343 B.n425 B.n52 585
R344 B.n52 B.n51 585
R345 B.n424 B.n423 585
R346 B.n423 B.n422 585
R347 B.n480 B.n479 585
R348 B.n478 B.n2 585
R349 B.n423 B.n54 497.305
R350 B.n419 B.n55 497.305
R351 B.n296 B.n202 497.305
R352 B.n298 B.n200 497.305
R353 B.n421 B.n420 256.663
R354 B.n421 B.n72 256.663
R355 B.n421 B.n71 256.663
R356 B.n421 B.n70 256.663
R357 B.n421 B.n69 256.663
R358 B.n421 B.n68 256.663
R359 B.n421 B.n67 256.663
R360 B.n421 B.n66 256.663
R361 B.n421 B.n65 256.663
R362 B.n421 B.n64 256.663
R363 B.n421 B.n63 256.663
R364 B.n421 B.n62 256.663
R365 B.n421 B.n61 256.663
R366 B.n421 B.n60 256.663
R367 B.n421 B.n59 256.663
R368 B.n421 B.n58 256.663
R369 B.n421 B.n57 256.663
R370 B.n421 B.n56 256.663
R371 B.n225 B.n201 256.663
R372 B.n231 B.n201 256.663
R373 B.n233 B.n201 256.663
R374 B.n239 B.n201 256.663
R375 B.n241 B.n201 256.663
R376 B.n247 B.n201 256.663
R377 B.n249 B.n201 256.663
R378 B.n255 B.n201 256.663
R379 B.n257 B.n201 256.663
R380 B.n263 B.n201 256.663
R381 B.n265 B.n201 256.663
R382 B.n272 B.n201 256.663
R383 B.n274 B.n201 256.663
R384 B.n280 B.n201 256.663
R385 B.n282 B.n201 256.663
R386 B.n288 B.n201 256.663
R387 B.n291 B.n201 256.663
R388 B.n482 B.n481 256.663
R389 B.n76 B.t8 235.352
R390 B.n74 B.t12 235.352
R391 B.n210 B.t15 235.352
R392 B.n216 B.t4 235.352
R393 B.n297 B.n201 177.677
R394 B.n422 B.n421 177.677
R395 B.n80 B.n79 163.367
R396 B.n84 B.n83 163.367
R397 B.n88 B.n87 163.367
R398 B.n92 B.n91 163.367
R399 B.n96 B.n95 163.367
R400 B.n100 B.n99 163.367
R401 B.n105 B.n104 163.367
R402 B.n109 B.n108 163.367
R403 B.n113 B.n112 163.367
R404 B.n117 B.n116 163.367
R405 B.n121 B.n120 163.367
R406 B.n126 B.n125 163.367
R407 B.n130 B.n129 163.367
R408 B.n134 B.n133 163.367
R409 B.n138 B.n137 163.367
R410 B.n142 B.n141 163.367
R411 B.n144 B.n73 163.367
R412 B.n296 B.n196 163.367
R413 B.n304 B.n196 163.367
R414 B.n304 B.n194 163.367
R415 B.n308 B.n194 163.367
R416 B.n308 B.n188 163.367
R417 B.n316 B.n188 163.367
R418 B.n316 B.n186 163.367
R419 B.n320 B.n186 163.367
R420 B.n320 B.n180 163.367
R421 B.n328 B.n180 163.367
R422 B.n328 B.n178 163.367
R423 B.n332 B.n178 163.367
R424 B.n332 B.n172 163.367
R425 B.n340 B.n172 163.367
R426 B.n340 B.n170 163.367
R427 B.n344 B.n170 163.367
R428 B.n344 B.n164 163.367
R429 B.n352 B.n164 163.367
R430 B.n352 B.n162 163.367
R431 B.n356 B.n162 163.367
R432 B.n356 B.n155 163.367
R433 B.n364 B.n155 163.367
R434 B.n364 B.n153 163.367
R435 B.n369 B.n153 163.367
R436 B.n369 B.n148 163.367
R437 B.n377 B.n148 163.367
R438 B.n378 B.n377 163.367
R439 B.n378 B.n5 163.367
R440 B.n6 B.n5 163.367
R441 B.n7 B.n6 163.367
R442 B.n384 B.n7 163.367
R443 B.n385 B.n384 163.367
R444 B.n385 B.n13 163.367
R445 B.n14 B.n13 163.367
R446 B.n15 B.n14 163.367
R447 B.n390 B.n15 163.367
R448 B.n390 B.n20 163.367
R449 B.n21 B.n20 163.367
R450 B.n22 B.n21 163.367
R451 B.n395 B.n22 163.367
R452 B.n395 B.n27 163.367
R453 B.n28 B.n27 163.367
R454 B.n29 B.n28 163.367
R455 B.n400 B.n29 163.367
R456 B.n400 B.n34 163.367
R457 B.n35 B.n34 163.367
R458 B.n36 B.n35 163.367
R459 B.n405 B.n36 163.367
R460 B.n405 B.n41 163.367
R461 B.n42 B.n41 163.367
R462 B.n43 B.n42 163.367
R463 B.n410 B.n43 163.367
R464 B.n410 B.n48 163.367
R465 B.n49 B.n48 163.367
R466 B.n50 B.n49 163.367
R467 B.n415 B.n50 163.367
R468 B.n415 B.n55 163.367
R469 B.n226 B.n224 163.367
R470 B.n230 B.n224 163.367
R471 B.n234 B.n232 163.367
R472 B.n238 B.n222 163.367
R473 B.n242 B.n240 163.367
R474 B.n246 B.n220 163.367
R475 B.n250 B.n248 163.367
R476 B.n254 B.n215 163.367
R477 B.n258 B.n256 163.367
R478 B.n262 B.n213 163.367
R479 B.n266 B.n264 163.367
R480 B.n271 B.n209 163.367
R481 B.n275 B.n273 163.367
R482 B.n279 B.n207 163.367
R483 B.n283 B.n281 163.367
R484 B.n287 B.n205 163.367
R485 B.n290 B.n289 163.367
R486 B.n292 B.n202 163.367
R487 B.n298 B.n198 163.367
R488 B.n302 B.n198 163.367
R489 B.n302 B.n192 163.367
R490 B.n310 B.n192 163.367
R491 B.n310 B.n190 163.367
R492 B.n314 B.n190 163.367
R493 B.n314 B.n184 163.367
R494 B.n322 B.n184 163.367
R495 B.n322 B.n182 163.367
R496 B.n326 B.n182 163.367
R497 B.n326 B.n176 163.367
R498 B.n334 B.n176 163.367
R499 B.n334 B.n174 163.367
R500 B.n338 B.n174 163.367
R501 B.n338 B.n168 163.367
R502 B.n346 B.n168 163.367
R503 B.n346 B.n166 163.367
R504 B.n350 B.n166 163.367
R505 B.n350 B.n160 163.367
R506 B.n358 B.n160 163.367
R507 B.n358 B.n158 163.367
R508 B.n362 B.n158 163.367
R509 B.n362 B.n152 163.367
R510 B.n371 B.n152 163.367
R511 B.n371 B.n150 163.367
R512 B.n375 B.n150 163.367
R513 B.n375 B.n3 163.367
R514 B.n480 B.n3 163.367
R515 B.n476 B.n2 163.367
R516 B.n476 B.n475 163.367
R517 B.n475 B.n9 163.367
R518 B.n471 B.n9 163.367
R519 B.n471 B.n11 163.367
R520 B.n467 B.n11 163.367
R521 B.n467 B.n17 163.367
R522 B.n463 B.n17 163.367
R523 B.n463 B.n19 163.367
R524 B.n459 B.n19 163.367
R525 B.n459 B.n24 163.367
R526 B.n455 B.n24 163.367
R527 B.n455 B.n26 163.367
R528 B.n451 B.n26 163.367
R529 B.n451 B.n31 163.367
R530 B.n447 B.n31 163.367
R531 B.n447 B.n33 163.367
R532 B.n443 B.n33 163.367
R533 B.n443 B.n38 163.367
R534 B.n439 B.n38 163.367
R535 B.n439 B.n40 163.367
R536 B.n435 B.n40 163.367
R537 B.n435 B.n45 163.367
R538 B.n431 B.n45 163.367
R539 B.n431 B.n47 163.367
R540 B.n427 B.n47 163.367
R541 B.n427 B.n52 163.367
R542 B.n423 B.n52 163.367
R543 B.n74 B.t13 132.685
R544 B.n210 B.t17 132.685
R545 B.n76 B.t10 132.685
R546 B.n216 B.t7 132.685
R547 B.n297 B.n197 98.2277
R548 B.n303 B.n197 98.2277
R549 B.n303 B.n193 98.2277
R550 B.n309 B.n193 98.2277
R551 B.n309 B.n189 98.2277
R552 B.n315 B.n189 98.2277
R553 B.n321 B.n185 98.2277
R554 B.n321 B.n181 98.2277
R555 B.n327 B.n181 98.2277
R556 B.n327 B.n177 98.2277
R557 B.n333 B.n177 98.2277
R558 B.n333 B.n173 98.2277
R559 B.n339 B.n173 98.2277
R560 B.n339 B.n169 98.2277
R561 B.n345 B.n169 98.2277
R562 B.n351 B.n165 98.2277
R563 B.n351 B.n161 98.2277
R564 B.n357 B.n161 98.2277
R565 B.n357 B.n156 98.2277
R566 B.n363 B.n156 98.2277
R567 B.n363 B.n157 98.2277
R568 B.n370 B.n149 98.2277
R569 B.n376 B.n149 98.2277
R570 B.n376 B.n4 98.2277
R571 B.n479 B.n4 98.2277
R572 B.n479 B.n478 98.2277
R573 B.n478 B.n477 98.2277
R574 B.n477 B.n8 98.2277
R575 B.n12 B.n8 98.2277
R576 B.n470 B.n12 98.2277
R577 B.n469 B.n468 98.2277
R578 B.n468 B.n16 98.2277
R579 B.n462 B.n16 98.2277
R580 B.n462 B.n461 98.2277
R581 B.n461 B.n460 98.2277
R582 B.n460 B.n23 98.2277
R583 B.n454 B.n453 98.2277
R584 B.n453 B.n452 98.2277
R585 B.n452 B.n30 98.2277
R586 B.n446 B.n30 98.2277
R587 B.n446 B.n445 98.2277
R588 B.n445 B.n444 98.2277
R589 B.n444 B.n37 98.2277
R590 B.n438 B.n37 98.2277
R591 B.n438 B.n437 98.2277
R592 B.n436 B.n44 98.2277
R593 B.n430 B.n44 98.2277
R594 B.n430 B.n429 98.2277
R595 B.n429 B.n428 98.2277
R596 B.n428 B.n51 98.2277
R597 B.n422 B.n51 98.2277
R598 B.n75 B.t14 87.8845
R599 B.n211 B.t16 87.8845
R600 B.n77 B.t11 87.8842
R601 B.n217 B.t6 87.8842
R602 B.n56 B.n54 71.676
R603 B.n80 B.n57 71.676
R604 B.n84 B.n58 71.676
R605 B.n88 B.n59 71.676
R606 B.n92 B.n60 71.676
R607 B.n96 B.n61 71.676
R608 B.n100 B.n62 71.676
R609 B.n105 B.n63 71.676
R610 B.n109 B.n64 71.676
R611 B.n113 B.n65 71.676
R612 B.n117 B.n66 71.676
R613 B.n121 B.n67 71.676
R614 B.n126 B.n68 71.676
R615 B.n130 B.n69 71.676
R616 B.n134 B.n70 71.676
R617 B.n138 B.n71 71.676
R618 B.n142 B.n72 71.676
R619 B.n420 B.n73 71.676
R620 B.n420 B.n419 71.676
R621 B.n144 B.n72 71.676
R622 B.n141 B.n71 71.676
R623 B.n137 B.n70 71.676
R624 B.n133 B.n69 71.676
R625 B.n129 B.n68 71.676
R626 B.n125 B.n67 71.676
R627 B.n120 B.n66 71.676
R628 B.n116 B.n65 71.676
R629 B.n112 B.n64 71.676
R630 B.n108 B.n63 71.676
R631 B.n104 B.n62 71.676
R632 B.n99 B.n61 71.676
R633 B.n95 B.n60 71.676
R634 B.n91 B.n59 71.676
R635 B.n87 B.n58 71.676
R636 B.n83 B.n57 71.676
R637 B.n79 B.n56 71.676
R638 B.n225 B.n200 71.676
R639 B.n231 B.n230 71.676
R640 B.n234 B.n233 71.676
R641 B.n239 B.n238 71.676
R642 B.n242 B.n241 71.676
R643 B.n247 B.n246 71.676
R644 B.n250 B.n249 71.676
R645 B.n255 B.n254 71.676
R646 B.n258 B.n257 71.676
R647 B.n263 B.n262 71.676
R648 B.n266 B.n265 71.676
R649 B.n272 B.n271 71.676
R650 B.n275 B.n274 71.676
R651 B.n280 B.n279 71.676
R652 B.n283 B.n282 71.676
R653 B.n288 B.n287 71.676
R654 B.n291 B.n290 71.676
R655 B.n226 B.n225 71.676
R656 B.n232 B.n231 71.676
R657 B.n233 B.n222 71.676
R658 B.n240 B.n239 71.676
R659 B.n241 B.n220 71.676
R660 B.n248 B.n247 71.676
R661 B.n249 B.n215 71.676
R662 B.n256 B.n255 71.676
R663 B.n257 B.n213 71.676
R664 B.n264 B.n263 71.676
R665 B.n265 B.n209 71.676
R666 B.n273 B.n272 71.676
R667 B.n274 B.n207 71.676
R668 B.n281 B.n280 71.676
R669 B.n282 B.n205 71.676
R670 B.n289 B.n288 71.676
R671 B.n292 B.n291 71.676
R672 B.n481 B.n480 71.676
R673 B.n481 B.n2 71.676
R674 B.n315 B.t5 69.3373
R675 B.n345 B.t0 69.3373
R676 B.n454 B.t1 69.3373
R677 B.t9 B.n436 69.3373
R678 B.n102 B.n77 59.5399
R679 B.n123 B.n75 59.5399
R680 B.n269 B.n211 59.5399
R681 B.n218 B.n217 59.5399
R682 B.n157 B.t2 49.1141
R683 B.n370 B.t2 49.1141
R684 B.n470 B.t3 49.1141
R685 B.t3 B.n469 49.1141
R686 B.n77 B.n76 44.8005
R687 B.n75 B.n74 44.8005
R688 B.n211 B.n210 44.8005
R689 B.n217 B.n216 44.8005
R690 B.n299 B.n199 32.3127
R691 B.n295 B.n294 32.3127
R692 B.n418 B.n417 32.3127
R693 B.n424 B.n53 32.3127
R694 B.t5 B.n185 28.8908
R695 B.t0 B.n165 28.8908
R696 B.t1 B.n23 28.8908
R697 B.n437 B.t9 28.8908
R698 B B.n482 18.0485
R699 B.n300 B.n299 10.6151
R700 B.n301 B.n300 10.6151
R701 B.n301 B.n191 10.6151
R702 B.n311 B.n191 10.6151
R703 B.n312 B.n311 10.6151
R704 B.n313 B.n312 10.6151
R705 B.n313 B.n183 10.6151
R706 B.n323 B.n183 10.6151
R707 B.n324 B.n323 10.6151
R708 B.n325 B.n324 10.6151
R709 B.n325 B.n175 10.6151
R710 B.n335 B.n175 10.6151
R711 B.n336 B.n335 10.6151
R712 B.n337 B.n336 10.6151
R713 B.n337 B.n167 10.6151
R714 B.n347 B.n167 10.6151
R715 B.n348 B.n347 10.6151
R716 B.n349 B.n348 10.6151
R717 B.n349 B.n159 10.6151
R718 B.n359 B.n159 10.6151
R719 B.n360 B.n359 10.6151
R720 B.n361 B.n360 10.6151
R721 B.n361 B.n151 10.6151
R722 B.n372 B.n151 10.6151
R723 B.n373 B.n372 10.6151
R724 B.n374 B.n373 10.6151
R725 B.n374 B.n0 10.6151
R726 B.n227 B.n199 10.6151
R727 B.n228 B.n227 10.6151
R728 B.n229 B.n228 10.6151
R729 B.n229 B.n223 10.6151
R730 B.n235 B.n223 10.6151
R731 B.n236 B.n235 10.6151
R732 B.n237 B.n236 10.6151
R733 B.n237 B.n221 10.6151
R734 B.n243 B.n221 10.6151
R735 B.n244 B.n243 10.6151
R736 B.n245 B.n244 10.6151
R737 B.n245 B.n219 10.6151
R738 B.n252 B.n251 10.6151
R739 B.n253 B.n252 10.6151
R740 B.n253 B.n214 10.6151
R741 B.n259 B.n214 10.6151
R742 B.n260 B.n259 10.6151
R743 B.n261 B.n260 10.6151
R744 B.n261 B.n212 10.6151
R745 B.n267 B.n212 10.6151
R746 B.n268 B.n267 10.6151
R747 B.n270 B.n208 10.6151
R748 B.n276 B.n208 10.6151
R749 B.n277 B.n276 10.6151
R750 B.n278 B.n277 10.6151
R751 B.n278 B.n206 10.6151
R752 B.n284 B.n206 10.6151
R753 B.n285 B.n284 10.6151
R754 B.n286 B.n285 10.6151
R755 B.n286 B.n204 10.6151
R756 B.n204 B.n203 10.6151
R757 B.n293 B.n203 10.6151
R758 B.n294 B.n293 10.6151
R759 B.n295 B.n195 10.6151
R760 B.n305 B.n195 10.6151
R761 B.n306 B.n305 10.6151
R762 B.n307 B.n306 10.6151
R763 B.n307 B.n187 10.6151
R764 B.n317 B.n187 10.6151
R765 B.n318 B.n317 10.6151
R766 B.n319 B.n318 10.6151
R767 B.n319 B.n179 10.6151
R768 B.n329 B.n179 10.6151
R769 B.n330 B.n329 10.6151
R770 B.n331 B.n330 10.6151
R771 B.n331 B.n171 10.6151
R772 B.n341 B.n171 10.6151
R773 B.n342 B.n341 10.6151
R774 B.n343 B.n342 10.6151
R775 B.n343 B.n163 10.6151
R776 B.n353 B.n163 10.6151
R777 B.n354 B.n353 10.6151
R778 B.n355 B.n354 10.6151
R779 B.n355 B.n154 10.6151
R780 B.n365 B.n154 10.6151
R781 B.n366 B.n365 10.6151
R782 B.n368 B.n366 10.6151
R783 B.n368 B.n367 10.6151
R784 B.n367 B.n147 10.6151
R785 B.n379 B.n147 10.6151
R786 B.n380 B.n379 10.6151
R787 B.n381 B.n380 10.6151
R788 B.n382 B.n381 10.6151
R789 B.n383 B.n382 10.6151
R790 B.n386 B.n383 10.6151
R791 B.n387 B.n386 10.6151
R792 B.n388 B.n387 10.6151
R793 B.n389 B.n388 10.6151
R794 B.n391 B.n389 10.6151
R795 B.n392 B.n391 10.6151
R796 B.n393 B.n392 10.6151
R797 B.n394 B.n393 10.6151
R798 B.n396 B.n394 10.6151
R799 B.n397 B.n396 10.6151
R800 B.n398 B.n397 10.6151
R801 B.n399 B.n398 10.6151
R802 B.n401 B.n399 10.6151
R803 B.n402 B.n401 10.6151
R804 B.n403 B.n402 10.6151
R805 B.n404 B.n403 10.6151
R806 B.n406 B.n404 10.6151
R807 B.n407 B.n406 10.6151
R808 B.n408 B.n407 10.6151
R809 B.n409 B.n408 10.6151
R810 B.n411 B.n409 10.6151
R811 B.n412 B.n411 10.6151
R812 B.n413 B.n412 10.6151
R813 B.n414 B.n413 10.6151
R814 B.n416 B.n414 10.6151
R815 B.n417 B.n416 10.6151
R816 B.n474 B.n1 10.6151
R817 B.n474 B.n473 10.6151
R818 B.n473 B.n472 10.6151
R819 B.n472 B.n10 10.6151
R820 B.n466 B.n10 10.6151
R821 B.n466 B.n465 10.6151
R822 B.n465 B.n464 10.6151
R823 B.n464 B.n18 10.6151
R824 B.n458 B.n18 10.6151
R825 B.n458 B.n457 10.6151
R826 B.n457 B.n456 10.6151
R827 B.n456 B.n25 10.6151
R828 B.n450 B.n25 10.6151
R829 B.n450 B.n449 10.6151
R830 B.n449 B.n448 10.6151
R831 B.n448 B.n32 10.6151
R832 B.n442 B.n32 10.6151
R833 B.n442 B.n441 10.6151
R834 B.n441 B.n440 10.6151
R835 B.n440 B.n39 10.6151
R836 B.n434 B.n39 10.6151
R837 B.n434 B.n433 10.6151
R838 B.n433 B.n432 10.6151
R839 B.n432 B.n46 10.6151
R840 B.n426 B.n46 10.6151
R841 B.n426 B.n425 10.6151
R842 B.n425 B.n424 10.6151
R843 B.n78 B.n53 10.6151
R844 B.n81 B.n78 10.6151
R845 B.n82 B.n81 10.6151
R846 B.n85 B.n82 10.6151
R847 B.n86 B.n85 10.6151
R848 B.n89 B.n86 10.6151
R849 B.n90 B.n89 10.6151
R850 B.n93 B.n90 10.6151
R851 B.n94 B.n93 10.6151
R852 B.n97 B.n94 10.6151
R853 B.n98 B.n97 10.6151
R854 B.n101 B.n98 10.6151
R855 B.n106 B.n103 10.6151
R856 B.n107 B.n106 10.6151
R857 B.n110 B.n107 10.6151
R858 B.n111 B.n110 10.6151
R859 B.n114 B.n111 10.6151
R860 B.n115 B.n114 10.6151
R861 B.n118 B.n115 10.6151
R862 B.n119 B.n118 10.6151
R863 B.n122 B.n119 10.6151
R864 B.n127 B.n124 10.6151
R865 B.n128 B.n127 10.6151
R866 B.n131 B.n128 10.6151
R867 B.n132 B.n131 10.6151
R868 B.n135 B.n132 10.6151
R869 B.n136 B.n135 10.6151
R870 B.n139 B.n136 10.6151
R871 B.n140 B.n139 10.6151
R872 B.n143 B.n140 10.6151
R873 B.n145 B.n143 10.6151
R874 B.n146 B.n145 10.6151
R875 B.n418 B.n146 10.6151
R876 B.n219 B.n218 9.36635
R877 B.n270 B.n269 9.36635
R878 B.n102 B.n101 9.36635
R879 B.n124 B.n123 9.36635
R880 B.n482 B.n0 8.11757
R881 B.n482 B.n1 8.11757
R882 B.n251 B.n218 1.24928
R883 B.n269 B.n268 1.24928
R884 B.n103 B.n102 1.24928
R885 B.n123 B.n122 1.24928
R886 VN.n0 VN.t3 64.0351
R887 VN.n1 VN.t2 64.0351
R888 VN.n0 VN.t1 63.5056
R889 VN.n1 VN.t0 63.5056
R890 VN VN.n1 44.6578
R891 VN VN.n0 7.3358
R892 VDD2.n2 VDD2.n0 123.017
R893 VDD2.n2 VDD2.n1 91.311
R894 VDD2.n1 VDD2.t3 8.46204
R895 VDD2.n1 VDD2.t1 8.46204
R896 VDD2.n0 VDD2.t0 8.46204
R897 VDD2.n0 VDD2.t2 8.46204
R898 VDD2 VDD2.n2 0.0586897
C0 VDD1 VN 0.154332f
C1 VDD2 VDD1 0.878951f
C2 VP VTAIL 1.53327f
C3 VP VN 3.96076f
C4 VTAIL VN 1.51916f
C5 VP VDD2 0.36148f
C6 VDD2 VTAIL 2.86601f
C7 VP VDD1 1.33295f
C8 VTAIL VDD1 2.81596f
C9 VDD2 VN 1.12721f
C10 VDD2 B 2.611456f
C11 VDD1 B 4.70772f
C12 VTAIL B 3.648216f
C13 VN B 8.02538f
C14 VP B 6.780477f
C15 VDD2.t0 B 0.037654f
C16 VDD2.t2 B 0.037654f
C17 VDD2.n0 B 0.446269f
C18 VDD2.t3 B 0.037654f
C19 VDD2.t1 B 0.037654f
C20 VDD2.n1 B 0.251295f
C21 VDD2.n2 B 1.91677f
C22 VN.t3 B 0.387213f
C23 VN.t1 B 0.385263f
C24 VN.n0 B 0.267304f
C25 VN.t2 B 0.387213f
C26 VN.t0 B 0.385263f
C27 VN.n1 B 1.06057f
C28 VDD1.t1 B 0.035436f
C29 VDD1.t3 B 0.035436f
C30 VDD1.n0 B 0.236677f
C31 VDD1.t2 B 0.035436f
C32 VDD1.t0 B 0.035436f
C33 VDD1.n1 B 0.432428f
C34 VTAIL.t3 B 0.229863f
C35 VTAIL.n0 B 0.232817f
C36 VTAIL.t6 B 0.229863f
C37 VTAIL.n1 B 0.28146f
C38 VTAIL.t5 B 0.229863f
C39 VTAIL.n2 B 0.683813f
C40 VTAIL.t0 B 0.229864f
C41 VTAIL.n3 B 0.683812f
C42 VTAIL.t2 B 0.229864f
C43 VTAIL.n4 B 0.281459f
C44 VTAIL.t7 B 0.229864f
C45 VTAIL.n5 B 0.281459f
C46 VTAIL.t4 B 0.229864f
C47 VTAIL.n6 B 0.683812f
C48 VTAIL.t1 B 0.229863f
C49 VTAIL.n7 B 0.629131f
C50 VP.n0 B 0.030392f
C51 VP.t3 B 0.256694f
C52 VP.n1 B 0.033512f
C53 VP.t0 B 0.388384f
C54 VP.t2 B 0.39035f
C55 VP.n2 B 1.05724f
C56 VP.n3 B 0.964335f
C57 VP.t1 B 0.256694f
C58 VP.n4 B 0.190487f
C59 VP.n5 B 0.03874f
C60 VP.n6 B 0.030392f
C61 VP.n7 B 0.023053f
C62 VP.n8 B 0.023053f
C63 VP.n9 B 0.033512f
C64 VP.n10 B 0.03874f
C65 VP.n11 B 0.190487f
C66 VP.n12 B 0.027886f
.ends

