* NGSPICE file created from diff_pair_sample_1756.ext - technology: sky130A

.subckt diff_pair_sample_1756 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t7 VP.t0 VDD1.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=6.8679 pd=36 as=2.90565 ps=17.94 w=17.61 l=2.84
X1 VDD1.t1 VP.t1 VTAIL.t6 B.t1 sky130_fd_pr__nfet_01v8 ad=2.90565 pd=17.94 as=6.8679 ps=36 w=17.61 l=2.84
X2 B.t17 B.t15 B.t16 B.t9 sky130_fd_pr__nfet_01v8 ad=6.8679 pd=36 as=0 ps=0 w=17.61 l=2.84
X3 VDD1.t3 VP.t2 VTAIL.t5 B.t3 sky130_fd_pr__nfet_01v8 ad=2.90565 pd=17.94 as=6.8679 ps=36 w=17.61 l=2.84
X4 B.t14 B.t12 B.t13 B.t5 sky130_fd_pr__nfet_01v8 ad=6.8679 pd=36 as=0 ps=0 w=17.61 l=2.84
X5 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=6.8679 pd=36 as=0 ps=0 w=17.61 l=2.84
X6 VDD2.t3 VN.t0 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=2.90565 pd=17.94 as=6.8679 ps=36 w=17.61 l=2.84
X7 VTAIL.t2 VN.t1 VDD2.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=6.8679 pd=36 as=2.90565 ps=17.94 w=17.61 l=2.84
X8 VTAIL.t0 VN.t2 VDD2.t1 B.t0 sky130_fd_pr__nfet_01v8 ad=6.8679 pd=36 as=2.90565 ps=17.94 w=17.61 l=2.84
X9 B.t7 B.t4 B.t6 B.t5 sky130_fd_pr__nfet_01v8 ad=6.8679 pd=36 as=0 ps=0 w=17.61 l=2.84
X10 VTAIL.t4 VP.t3 VDD1.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=6.8679 pd=36 as=2.90565 ps=17.94 w=17.61 l=2.84
X11 VDD2.t0 VN.t3 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=2.90565 pd=17.94 as=6.8679 ps=36 w=17.61 l=2.84
R0 VP.n4 VP.t0 184.751
R1 VP.n4 VP.t1 183.856
R2 VP.n16 VP.n0 161.3
R3 VP.n15 VP.n14 161.3
R4 VP.n13 VP.n1 161.3
R5 VP.n12 VP.n11 161.3
R6 VP.n10 VP.n2 161.3
R7 VP.n9 VP.n8 161.3
R8 VP.n7 VP.n3 161.3
R9 VP.n5 VP.t3 149.438
R10 VP.n17 VP.t2 149.438
R11 VP.n6 VP.n5 106.597
R12 VP.n18 VP.n17 106.597
R13 VP.n6 VP.n4 54.7515
R14 VP.n11 VP.n10 40.4934
R15 VP.n11 VP.n1 40.4934
R16 VP.n9 VP.n3 24.4675
R17 VP.n10 VP.n9 24.4675
R18 VP.n15 VP.n1 24.4675
R19 VP.n16 VP.n15 24.4675
R20 VP.n5 VP.n3 4.15989
R21 VP.n17 VP.n16 4.15989
R22 VP.n7 VP.n6 0.278367
R23 VP.n18 VP.n0 0.278367
R24 VP.n8 VP.n7 0.189894
R25 VP.n8 VP.n2 0.189894
R26 VP.n12 VP.n2 0.189894
R27 VP.n13 VP.n12 0.189894
R28 VP.n14 VP.n13 0.189894
R29 VP.n14 VP.n0 0.189894
R30 VP VP.n18 0.153454
R31 VDD1 VDD1.n1 110.046
R32 VDD1 VDD1.n0 62.4856
R33 VDD1.n0 VDD1.t2 1.12486
R34 VDD1.n0 VDD1.t1 1.12486
R35 VDD1.n1 VDD1.t0 1.12486
R36 VDD1.n1 VDD1.t3 1.12486
R37 VTAIL.n778 VTAIL.n686 289.615
R38 VTAIL.n92 VTAIL.n0 289.615
R39 VTAIL.n190 VTAIL.n98 289.615
R40 VTAIL.n288 VTAIL.n196 289.615
R41 VTAIL.n680 VTAIL.n588 289.615
R42 VTAIL.n582 VTAIL.n490 289.615
R43 VTAIL.n484 VTAIL.n392 289.615
R44 VTAIL.n386 VTAIL.n294 289.615
R45 VTAIL.n719 VTAIL.n718 185
R46 VTAIL.n721 VTAIL.n720 185
R47 VTAIL.n714 VTAIL.n713 185
R48 VTAIL.n727 VTAIL.n726 185
R49 VTAIL.n729 VTAIL.n728 185
R50 VTAIL.n710 VTAIL.n709 185
R51 VTAIL.n735 VTAIL.n734 185
R52 VTAIL.n737 VTAIL.n736 185
R53 VTAIL.n706 VTAIL.n705 185
R54 VTAIL.n743 VTAIL.n742 185
R55 VTAIL.n745 VTAIL.n744 185
R56 VTAIL.n702 VTAIL.n701 185
R57 VTAIL.n751 VTAIL.n750 185
R58 VTAIL.n753 VTAIL.n752 185
R59 VTAIL.n698 VTAIL.n697 185
R60 VTAIL.n760 VTAIL.n759 185
R61 VTAIL.n761 VTAIL.n696 185
R62 VTAIL.n763 VTAIL.n762 185
R63 VTAIL.n694 VTAIL.n693 185
R64 VTAIL.n769 VTAIL.n768 185
R65 VTAIL.n771 VTAIL.n770 185
R66 VTAIL.n690 VTAIL.n689 185
R67 VTAIL.n777 VTAIL.n776 185
R68 VTAIL.n779 VTAIL.n778 185
R69 VTAIL.n33 VTAIL.n32 185
R70 VTAIL.n35 VTAIL.n34 185
R71 VTAIL.n28 VTAIL.n27 185
R72 VTAIL.n41 VTAIL.n40 185
R73 VTAIL.n43 VTAIL.n42 185
R74 VTAIL.n24 VTAIL.n23 185
R75 VTAIL.n49 VTAIL.n48 185
R76 VTAIL.n51 VTAIL.n50 185
R77 VTAIL.n20 VTAIL.n19 185
R78 VTAIL.n57 VTAIL.n56 185
R79 VTAIL.n59 VTAIL.n58 185
R80 VTAIL.n16 VTAIL.n15 185
R81 VTAIL.n65 VTAIL.n64 185
R82 VTAIL.n67 VTAIL.n66 185
R83 VTAIL.n12 VTAIL.n11 185
R84 VTAIL.n74 VTAIL.n73 185
R85 VTAIL.n75 VTAIL.n10 185
R86 VTAIL.n77 VTAIL.n76 185
R87 VTAIL.n8 VTAIL.n7 185
R88 VTAIL.n83 VTAIL.n82 185
R89 VTAIL.n85 VTAIL.n84 185
R90 VTAIL.n4 VTAIL.n3 185
R91 VTAIL.n91 VTAIL.n90 185
R92 VTAIL.n93 VTAIL.n92 185
R93 VTAIL.n131 VTAIL.n130 185
R94 VTAIL.n133 VTAIL.n132 185
R95 VTAIL.n126 VTAIL.n125 185
R96 VTAIL.n139 VTAIL.n138 185
R97 VTAIL.n141 VTAIL.n140 185
R98 VTAIL.n122 VTAIL.n121 185
R99 VTAIL.n147 VTAIL.n146 185
R100 VTAIL.n149 VTAIL.n148 185
R101 VTAIL.n118 VTAIL.n117 185
R102 VTAIL.n155 VTAIL.n154 185
R103 VTAIL.n157 VTAIL.n156 185
R104 VTAIL.n114 VTAIL.n113 185
R105 VTAIL.n163 VTAIL.n162 185
R106 VTAIL.n165 VTAIL.n164 185
R107 VTAIL.n110 VTAIL.n109 185
R108 VTAIL.n172 VTAIL.n171 185
R109 VTAIL.n173 VTAIL.n108 185
R110 VTAIL.n175 VTAIL.n174 185
R111 VTAIL.n106 VTAIL.n105 185
R112 VTAIL.n181 VTAIL.n180 185
R113 VTAIL.n183 VTAIL.n182 185
R114 VTAIL.n102 VTAIL.n101 185
R115 VTAIL.n189 VTAIL.n188 185
R116 VTAIL.n191 VTAIL.n190 185
R117 VTAIL.n229 VTAIL.n228 185
R118 VTAIL.n231 VTAIL.n230 185
R119 VTAIL.n224 VTAIL.n223 185
R120 VTAIL.n237 VTAIL.n236 185
R121 VTAIL.n239 VTAIL.n238 185
R122 VTAIL.n220 VTAIL.n219 185
R123 VTAIL.n245 VTAIL.n244 185
R124 VTAIL.n247 VTAIL.n246 185
R125 VTAIL.n216 VTAIL.n215 185
R126 VTAIL.n253 VTAIL.n252 185
R127 VTAIL.n255 VTAIL.n254 185
R128 VTAIL.n212 VTAIL.n211 185
R129 VTAIL.n261 VTAIL.n260 185
R130 VTAIL.n263 VTAIL.n262 185
R131 VTAIL.n208 VTAIL.n207 185
R132 VTAIL.n270 VTAIL.n269 185
R133 VTAIL.n271 VTAIL.n206 185
R134 VTAIL.n273 VTAIL.n272 185
R135 VTAIL.n204 VTAIL.n203 185
R136 VTAIL.n279 VTAIL.n278 185
R137 VTAIL.n281 VTAIL.n280 185
R138 VTAIL.n200 VTAIL.n199 185
R139 VTAIL.n287 VTAIL.n286 185
R140 VTAIL.n289 VTAIL.n288 185
R141 VTAIL.n681 VTAIL.n680 185
R142 VTAIL.n679 VTAIL.n678 185
R143 VTAIL.n592 VTAIL.n591 185
R144 VTAIL.n673 VTAIL.n672 185
R145 VTAIL.n671 VTAIL.n670 185
R146 VTAIL.n596 VTAIL.n595 185
R147 VTAIL.n600 VTAIL.n598 185
R148 VTAIL.n665 VTAIL.n664 185
R149 VTAIL.n663 VTAIL.n662 185
R150 VTAIL.n602 VTAIL.n601 185
R151 VTAIL.n657 VTAIL.n656 185
R152 VTAIL.n655 VTAIL.n654 185
R153 VTAIL.n606 VTAIL.n605 185
R154 VTAIL.n649 VTAIL.n648 185
R155 VTAIL.n647 VTAIL.n646 185
R156 VTAIL.n610 VTAIL.n609 185
R157 VTAIL.n641 VTAIL.n640 185
R158 VTAIL.n639 VTAIL.n638 185
R159 VTAIL.n614 VTAIL.n613 185
R160 VTAIL.n633 VTAIL.n632 185
R161 VTAIL.n631 VTAIL.n630 185
R162 VTAIL.n618 VTAIL.n617 185
R163 VTAIL.n625 VTAIL.n624 185
R164 VTAIL.n623 VTAIL.n622 185
R165 VTAIL.n583 VTAIL.n582 185
R166 VTAIL.n581 VTAIL.n580 185
R167 VTAIL.n494 VTAIL.n493 185
R168 VTAIL.n575 VTAIL.n574 185
R169 VTAIL.n573 VTAIL.n572 185
R170 VTAIL.n498 VTAIL.n497 185
R171 VTAIL.n502 VTAIL.n500 185
R172 VTAIL.n567 VTAIL.n566 185
R173 VTAIL.n565 VTAIL.n564 185
R174 VTAIL.n504 VTAIL.n503 185
R175 VTAIL.n559 VTAIL.n558 185
R176 VTAIL.n557 VTAIL.n556 185
R177 VTAIL.n508 VTAIL.n507 185
R178 VTAIL.n551 VTAIL.n550 185
R179 VTAIL.n549 VTAIL.n548 185
R180 VTAIL.n512 VTAIL.n511 185
R181 VTAIL.n543 VTAIL.n542 185
R182 VTAIL.n541 VTAIL.n540 185
R183 VTAIL.n516 VTAIL.n515 185
R184 VTAIL.n535 VTAIL.n534 185
R185 VTAIL.n533 VTAIL.n532 185
R186 VTAIL.n520 VTAIL.n519 185
R187 VTAIL.n527 VTAIL.n526 185
R188 VTAIL.n525 VTAIL.n524 185
R189 VTAIL.n485 VTAIL.n484 185
R190 VTAIL.n483 VTAIL.n482 185
R191 VTAIL.n396 VTAIL.n395 185
R192 VTAIL.n477 VTAIL.n476 185
R193 VTAIL.n475 VTAIL.n474 185
R194 VTAIL.n400 VTAIL.n399 185
R195 VTAIL.n404 VTAIL.n402 185
R196 VTAIL.n469 VTAIL.n468 185
R197 VTAIL.n467 VTAIL.n466 185
R198 VTAIL.n406 VTAIL.n405 185
R199 VTAIL.n461 VTAIL.n460 185
R200 VTAIL.n459 VTAIL.n458 185
R201 VTAIL.n410 VTAIL.n409 185
R202 VTAIL.n453 VTAIL.n452 185
R203 VTAIL.n451 VTAIL.n450 185
R204 VTAIL.n414 VTAIL.n413 185
R205 VTAIL.n445 VTAIL.n444 185
R206 VTAIL.n443 VTAIL.n442 185
R207 VTAIL.n418 VTAIL.n417 185
R208 VTAIL.n437 VTAIL.n436 185
R209 VTAIL.n435 VTAIL.n434 185
R210 VTAIL.n422 VTAIL.n421 185
R211 VTAIL.n429 VTAIL.n428 185
R212 VTAIL.n427 VTAIL.n426 185
R213 VTAIL.n387 VTAIL.n386 185
R214 VTAIL.n385 VTAIL.n384 185
R215 VTAIL.n298 VTAIL.n297 185
R216 VTAIL.n379 VTAIL.n378 185
R217 VTAIL.n377 VTAIL.n376 185
R218 VTAIL.n302 VTAIL.n301 185
R219 VTAIL.n306 VTAIL.n304 185
R220 VTAIL.n371 VTAIL.n370 185
R221 VTAIL.n369 VTAIL.n368 185
R222 VTAIL.n308 VTAIL.n307 185
R223 VTAIL.n363 VTAIL.n362 185
R224 VTAIL.n361 VTAIL.n360 185
R225 VTAIL.n312 VTAIL.n311 185
R226 VTAIL.n355 VTAIL.n354 185
R227 VTAIL.n353 VTAIL.n352 185
R228 VTAIL.n316 VTAIL.n315 185
R229 VTAIL.n347 VTAIL.n346 185
R230 VTAIL.n345 VTAIL.n344 185
R231 VTAIL.n320 VTAIL.n319 185
R232 VTAIL.n339 VTAIL.n338 185
R233 VTAIL.n337 VTAIL.n336 185
R234 VTAIL.n324 VTAIL.n323 185
R235 VTAIL.n331 VTAIL.n330 185
R236 VTAIL.n329 VTAIL.n328 185
R237 VTAIL.n717 VTAIL.t1 147.659
R238 VTAIL.n31 VTAIL.t2 147.659
R239 VTAIL.n129 VTAIL.t5 147.659
R240 VTAIL.n227 VTAIL.t4 147.659
R241 VTAIL.n621 VTAIL.t6 147.659
R242 VTAIL.n523 VTAIL.t7 147.659
R243 VTAIL.n425 VTAIL.t3 147.659
R244 VTAIL.n327 VTAIL.t0 147.659
R245 VTAIL.n720 VTAIL.n719 104.615
R246 VTAIL.n720 VTAIL.n713 104.615
R247 VTAIL.n727 VTAIL.n713 104.615
R248 VTAIL.n728 VTAIL.n727 104.615
R249 VTAIL.n728 VTAIL.n709 104.615
R250 VTAIL.n735 VTAIL.n709 104.615
R251 VTAIL.n736 VTAIL.n735 104.615
R252 VTAIL.n736 VTAIL.n705 104.615
R253 VTAIL.n743 VTAIL.n705 104.615
R254 VTAIL.n744 VTAIL.n743 104.615
R255 VTAIL.n744 VTAIL.n701 104.615
R256 VTAIL.n751 VTAIL.n701 104.615
R257 VTAIL.n752 VTAIL.n751 104.615
R258 VTAIL.n752 VTAIL.n697 104.615
R259 VTAIL.n760 VTAIL.n697 104.615
R260 VTAIL.n761 VTAIL.n760 104.615
R261 VTAIL.n762 VTAIL.n761 104.615
R262 VTAIL.n762 VTAIL.n693 104.615
R263 VTAIL.n769 VTAIL.n693 104.615
R264 VTAIL.n770 VTAIL.n769 104.615
R265 VTAIL.n770 VTAIL.n689 104.615
R266 VTAIL.n777 VTAIL.n689 104.615
R267 VTAIL.n778 VTAIL.n777 104.615
R268 VTAIL.n34 VTAIL.n33 104.615
R269 VTAIL.n34 VTAIL.n27 104.615
R270 VTAIL.n41 VTAIL.n27 104.615
R271 VTAIL.n42 VTAIL.n41 104.615
R272 VTAIL.n42 VTAIL.n23 104.615
R273 VTAIL.n49 VTAIL.n23 104.615
R274 VTAIL.n50 VTAIL.n49 104.615
R275 VTAIL.n50 VTAIL.n19 104.615
R276 VTAIL.n57 VTAIL.n19 104.615
R277 VTAIL.n58 VTAIL.n57 104.615
R278 VTAIL.n58 VTAIL.n15 104.615
R279 VTAIL.n65 VTAIL.n15 104.615
R280 VTAIL.n66 VTAIL.n65 104.615
R281 VTAIL.n66 VTAIL.n11 104.615
R282 VTAIL.n74 VTAIL.n11 104.615
R283 VTAIL.n75 VTAIL.n74 104.615
R284 VTAIL.n76 VTAIL.n75 104.615
R285 VTAIL.n76 VTAIL.n7 104.615
R286 VTAIL.n83 VTAIL.n7 104.615
R287 VTAIL.n84 VTAIL.n83 104.615
R288 VTAIL.n84 VTAIL.n3 104.615
R289 VTAIL.n91 VTAIL.n3 104.615
R290 VTAIL.n92 VTAIL.n91 104.615
R291 VTAIL.n132 VTAIL.n131 104.615
R292 VTAIL.n132 VTAIL.n125 104.615
R293 VTAIL.n139 VTAIL.n125 104.615
R294 VTAIL.n140 VTAIL.n139 104.615
R295 VTAIL.n140 VTAIL.n121 104.615
R296 VTAIL.n147 VTAIL.n121 104.615
R297 VTAIL.n148 VTAIL.n147 104.615
R298 VTAIL.n148 VTAIL.n117 104.615
R299 VTAIL.n155 VTAIL.n117 104.615
R300 VTAIL.n156 VTAIL.n155 104.615
R301 VTAIL.n156 VTAIL.n113 104.615
R302 VTAIL.n163 VTAIL.n113 104.615
R303 VTAIL.n164 VTAIL.n163 104.615
R304 VTAIL.n164 VTAIL.n109 104.615
R305 VTAIL.n172 VTAIL.n109 104.615
R306 VTAIL.n173 VTAIL.n172 104.615
R307 VTAIL.n174 VTAIL.n173 104.615
R308 VTAIL.n174 VTAIL.n105 104.615
R309 VTAIL.n181 VTAIL.n105 104.615
R310 VTAIL.n182 VTAIL.n181 104.615
R311 VTAIL.n182 VTAIL.n101 104.615
R312 VTAIL.n189 VTAIL.n101 104.615
R313 VTAIL.n190 VTAIL.n189 104.615
R314 VTAIL.n230 VTAIL.n229 104.615
R315 VTAIL.n230 VTAIL.n223 104.615
R316 VTAIL.n237 VTAIL.n223 104.615
R317 VTAIL.n238 VTAIL.n237 104.615
R318 VTAIL.n238 VTAIL.n219 104.615
R319 VTAIL.n245 VTAIL.n219 104.615
R320 VTAIL.n246 VTAIL.n245 104.615
R321 VTAIL.n246 VTAIL.n215 104.615
R322 VTAIL.n253 VTAIL.n215 104.615
R323 VTAIL.n254 VTAIL.n253 104.615
R324 VTAIL.n254 VTAIL.n211 104.615
R325 VTAIL.n261 VTAIL.n211 104.615
R326 VTAIL.n262 VTAIL.n261 104.615
R327 VTAIL.n262 VTAIL.n207 104.615
R328 VTAIL.n270 VTAIL.n207 104.615
R329 VTAIL.n271 VTAIL.n270 104.615
R330 VTAIL.n272 VTAIL.n271 104.615
R331 VTAIL.n272 VTAIL.n203 104.615
R332 VTAIL.n279 VTAIL.n203 104.615
R333 VTAIL.n280 VTAIL.n279 104.615
R334 VTAIL.n280 VTAIL.n199 104.615
R335 VTAIL.n287 VTAIL.n199 104.615
R336 VTAIL.n288 VTAIL.n287 104.615
R337 VTAIL.n680 VTAIL.n679 104.615
R338 VTAIL.n679 VTAIL.n591 104.615
R339 VTAIL.n672 VTAIL.n591 104.615
R340 VTAIL.n672 VTAIL.n671 104.615
R341 VTAIL.n671 VTAIL.n595 104.615
R342 VTAIL.n600 VTAIL.n595 104.615
R343 VTAIL.n664 VTAIL.n600 104.615
R344 VTAIL.n664 VTAIL.n663 104.615
R345 VTAIL.n663 VTAIL.n601 104.615
R346 VTAIL.n656 VTAIL.n601 104.615
R347 VTAIL.n656 VTAIL.n655 104.615
R348 VTAIL.n655 VTAIL.n605 104.615
R349 VTAIL.n648 VTAIL.n605 104.615
R350 VTAIL.n648 VTAIL.n647 104.615
R351 VTAIL.n647 VTAIL.n609 104.615
R352 VTAIL.n640 VTAIL.n609 104.615
R353 VTAIL.n640 VTAIL.n639 104.615
R354 VTAIL.n639 VTAIL.n613 104.615
R355 VTAIL.n632 VTAIL.n613 104.615
R356 VTAIL.n632 VTAIL.n631 104.615
R357 VTAIL.n631 VTAIL.n617 104.615
R358 VTAIL.n624 VTAIL.n617 104.615
R359 VTAIL.n624 VTAIL.n623 104.615
R360 VTAIL.n582 VTAIL.n581 104.615
R361 VTAIL.n581 VTAIL.n493 104.615
R362 VTAIL.n574 VTAIL.n493 104.615
R363 VTAIL.n574 VTAIL.n573 104.615
R364 VTAIL.n573 VTAIL.n497 104.615
R365 VTAIL.n502 VTAIL.n497 104.615
R366 VTAIL.n566 VTAIL.n502 104.615
R367 VTAIL.n566 VTAIL.n565 104.615
R368 VTAIL.n565 VTAIL.n503 104.615
R369 VTAIL.n558 VTAIL.n503 104.615
R370 VTAIL.n558 VTAIL.n557 104.615
R371 VTAIL.n557 VTAIL.n507 104.615
R372 VTAIL.n550 VTAIL.n507 104.615
R373 VTAIL.n550 VTAIL.n549 104.615
R374 VTAIL.n549 VTAIL.n511 104.615
R375 VTAIL.n542 VTAIL.n511 104.615
R376 VTAIL.n542 VTAIL.n541 104.615
R377 VTAIL.n541 VTAIL.n515 104.615
R378 VTAIL.n534 VTAIL.n515 104.615
R379 VTAIL.n534 VTAIL.n533 104.615
R380 VTAIL.n533 VTAIL.n519 104.615
R381 VTAIL.n526 VTAIL.n519 104.615
R382 VTAIL.n526 VTAIL.n525 104.615
R383 VTAIL.n484 VTAIL.n483 104.615
R384 VTAIL.n483 VTAIL.n395 104.615
R385 VTAIL.n476 VTAIL.n395 104.615
R386 VTAIL.n476 VTAIL.n475 104.615
R387 VTAIL.n475 VTAIL.n399 104.615
R388 VTAIL.n404 VTAIL.n399 104.615
R389 VTAIL.n468 VTAIL.n404 104.615
R390 VTAIL.n468 VTAIL.n467 104.615
R391 VTAIL.n467 VTAIL.n405 104.615
R392 VTAIL.n460 VTAIL.n405 104.615
R393 VTAIL.n460 VTAIL.n459 104.615
R394 VTAIL.n459 VTAIL.n409 104.615
R395 VTAIL.n452 VTAIL.n409 104.615
R396 VTAIL.n452 VTAIL.n451 104.615
R397 VTAIL.n451 VTAIL.n413 104.615
R398 VTAIL.n444 VTAIL.n413 104.615
R399 VTAIL.n444 VTAIL.n443 104.615
R400 VTAIL.n443 VTAIL.n417 104.615
R401 VTAIL.n436 VTAIL.n417 104.615
R402 VTAIL.n436 VTAIL.n435 104.615
R403 VTAIL.n435 VTAIL.n421 104.615
R404 VTAIL.n428 VTAIL.n421 104.615
R405 VTAIL.n428 VTAIL.n427 104.615
R406 VTAIL.n386 VTAIL.n385 104.615
R407 VTAIL.n385 VTAIL.n297 104.615
R408 VTAIL.n378 VTAIL.n297 104.615
R409 VTAIL.n378 VTAIL.n377 104.615
R410 VTAIL.n377 VTAIL.n301 104.615
R411 VTAIL.n306 VTAIL.n301 104.615
R412 VTAIL.n370 VTAIL.n306 104.615
R413 VTAIL.n370 VTAIL.n369 104.615
R414 VTAIL.n369 VTAIL.n307 104.615
R415 VTAIL.n362 VTAIL.n307 104.615
R416 VTAIL.n362 VTAIL.n361 104.615
R417 VTAIL.n361 VTAIL.n311 104.615
R418 VTAIL.n354 VTAIL.n311 104.615
R419 VTAIL.n354 VTAIL.n353 104.615
R420 VTAIL.n353 VTAIL.n315 104.615
R421 VTAIL.n346 VTAIL.n315 104.615
R422 VTAIL.n346 VTAIL.n345 104.615
R423 VTAIL.n345 VTAIL.n319 104.615
R424 VTAIL.n338 VTAIL.n319 104.615
R425 VTAIL.n338 VTAIL.n337 104.615
R426 VTAIL.n337 VTAIL.n323 104.615
R427 VTAIL.n330 VTAIL.n323 104.615
R428 VTAIL.n330 VTAIL.n329 104.615
R429 VTAIL.n719 VTAIL.t1 52.3082
R430 VTAIL.n33 VTAIL.t2 52.3082
R431 VTAIL.n131 VTAIL.t5 52.3082
R432 VTAIL.n229 VTAIL.t4 52.3082
R433 VTAIL.n623 VTAIL.t6 52.3082
R434 VTAIL.n525 VTAIL.t7 52.3082
R435 VTAIL.n427 VTAIL.t3 52.3082
R436 VTAIL.n329 VTAIL.t0 52.3082
R437 VTAIL.n783 VTAIL.n782 33.9308
R438 VTAIL.n97 VTAIL.n96 33.9308
R439 VTAIL.n195 VTAIL.n194 33.9308
R440 VTAIL.n293 VTAIL.n292 33.9308
R441 VTAIL.n685 VTAIL.n684 33.9308
R442 VTAIL.n587 VTAIL.n586 33.9308
R443 VTAIL.n489 VTAIL.n488 33.9308
R444 VTAIL.n391 VTAIL.n390 33.9308
R445 VTAIL.n783 VTAIL.n685 30.2807
R446 VTAIL.n391 VTAIL.n293 30.2807
R447 VTAIL.n718 VTAIL.n717 15.6677
R448 VTAIL.n32 VTAIL.n31 15.6677
R449 VTAIL.n130 VTAIL.n129 15.6677
R450 VTAIL.n228 VTAIL.n227 15.6677
R451 VTAIL.n622 VTAIL.n621 15.6677
R452 VTAIL.n524 VTAIL.n523 15.6677
R453 VTAIL.n426 VTAIL.n425 15.6677
R454 VTAIL.n328 VTAIL.n327 15.6677
R455 VTAIL.n763 VTAIL.n694 13.1884
R456 VTAIL.n77 VTAIL.n8 13.1884
R457 VTAIL.n175 VTAIL.n106 13.1884
R458 VTAIL.n273 VTAIL.n204 13.1884
R459 VTAIL.n598 VTAIL.n596 13.1884
R460 VTAIL.n500 VTAIL.n498 13.1884
R461 VTAIL.n402 VTAIL.n400 13.1884
R462 VTAIL.n304 VTAIL.n302 13.1884
R463 VTAIL.n721 VTAIL.n716 12.8005
R464 VTAIL.n764 VTAIL.n696 12.8005
R465 VTAIL.n768 VTAIL.n767 12.8005
R466 VTAIL.n35 VTAIL.n30 12.8005
R467 VTAIL.n78 VTAIL.n10 12.8005
R468 VTAIL.n82 VTAIL.n81 12.8005
R469 VTAIL.n133 VTAIL.n128 12.8005
R470 VTAIL.n176 VTAIL.n108 12.8005
R471 VTAIL.n180 VTAIL.n179 12.8005
R472 VTAIL.n231 VTAIL.n226 12.8005
R473 VTAIL.n274 VTAIL.n206 12.8005
R474 VTAIL.n278 VTAIL.n277 12.8005
R475 VTAIL.n670 VTAIL.n669 12.8005
R476 VTAIL.n666 VTAIL.n665 12.8005
R477 VTAIL.n625 VTAIL.n620 12.8005
R478 VTAIL.n572 VTAIL.n571 12.8005
R479 VTAIL.n568 VTAIL.n567 12.8005
R480 VTAIL.n527 VTAIL.n522 12.8005
R481 VTAIL.n474 VTAIL.n473 12.8005
R482 VTAIL.n470 VTAIL.n469 12.8005
R483 VTAIL.n429 VTAIL.n424 12.8005
R484 VTAIL.n376 VTAIL.n375 12.8005
R485 VTAIL.n372 VTAIL.n371 12.8005
R486 VTAIL.n331 VTAIL.n326 12.8005
R487 VTAIL.n722 VTAIL.n714 12.0247
R488 VTAIL.n759 VTAIL.n758 12.0247
R489 VTAIL.n771 VTAIL.n692 12.0247
R490 VTAIL.n36 VTAIL.n28 12.0247
R491 VTAIL.n73 VTAIL.n72 12.0247
R492 VTAIL.n85 VTAIL.n6 12.0247
R493 VTAIL.n134 VTAIL.n126 12.0247
R494 VTAIL.n171 VTAIL.n170 12.0247
R495 VTAIL.n183 VTAIL.n104 12.0247
R496 VTAIL.n232 VTAIL.n224 12.0247
R497 VTAIL.n269 VTAIL.n268 12.0247
R498 VTAIL.n281 VTAIL.n202 12.0247
R499 VTAIL.n673 VTAIL.n594 12.0247
R500 VTAIL.n662 VTAIL.n599 12.0247
R501 VTAIL.n626 VTAIL.n618 12.0247
R502 VTAIL.n575 VTAIL.n496 12.0247
R503 VTAIL.n564 VTAIL.n501 12.0247
R504 VTAIL.n528 VTAIL.n520 12.0247
R505 VTAIL.n477 VTAIL.n398 12.0247
R506 VTAIL.n466 VTAIL.n403 12.0247
R507 VTAIL.n430 VTAIL.n422 12.0247
R508 VTAIL.n379 VTAIL.n300 12.0247
R509 VTAIL.n368 VTAIL.n305 12.0247
R510 VTAIL.n332 VTAIL.n324 12.0247
R511 VTAIL.n726 VTAIL.n725 11.249
R512 VTAIL.n757 VTAIL.n698 11.249
R513 VTAIL.n772 VTAIL.n690 11.249
R514 VTAIL.n40 VTAIL.n39 11.249
R515 VTAIL.n71 VTAIL.n12 11.249
R516 VTAIL.n86 VTAIL.n4 11.249
R517 VTAIL.n138 VTAIL.n137 11.249
R518 VTAIL.n169 VTAIL.n110 11.249
R519 VTAIL.n184 VTAIL.n102 11.249
R520 VTAIL.n236 VTAIL.n235 11.249
R521 VTAIL.n267 VTAIL.n208 11.249
R522 VTAIL.n282 VTAIL.n200 11.249
R523 VTAIL.n674 VTAIL.n592 11.249
R524 VTAIL.n661 VTAIL.n602 11.249
R525 VTAIL.n630 VTAIL.n629 11.249
R526 VTAIL.n576 VTAIL.n494 11.249
R527 VTAIL.n563 VTAIL.n504 11.249
R528 VTAIL.n532 VTAIL.n531 11.249
R529 VTAIL.n478 VTAIL.n396 11.249
R530 VTAIL.n465 VTAIL.n406 11.249
R531 VTAIL.n434 VTAIL.n433 11.249
R532 VTAIL.n380 VTAIL.n298 11.249
R533 VTAIL.n367 VTAIL.n308 11.249
R534 VTAIL.n336 VTAIL.n335 11.249
R535 VTAIL.n729 VTAIL.n712 10.4732
R536 VTAIL.n754 VTAIL.n753 10.4732
R537 VTAIL.n776 VTAIL.n775 10.4732
R538 VTAIL.n43 VTAIL.n26 10.4732
R539 VTAIL.n68 VTAIL.n67 10.4732
R540 VTAIL.n90 VTAIL.n89 10.4732
R541 VTAIL.n141 VTAIL.n124 10.4732
R542 VTAIL.n166 VTAIL.n165 10.4732
R543 VTAIL.n188 VTAIL.n187 10.4732
R544 VTAIL.n239 VTAIL.n222 10.4732
R545 VTAIL.n264 VTAIL.n263 10.4732
R546 VTAIL.n286 VTAIL.n285 10.4732
R547 VTAIL.n678 VTAIL.n677 10.4732
R548 VTAIL.n658 VTAIL.n657 10.4732
R549 VTAIL.n633 VTAIL.n616 10.4732
R550 VTAIL.n580 VTAIL.n579 10.4732
R551 VTAIL.n560 VTAIL.n559 10.4732
R552 VTAIL.n535 VTAIL.n518 10.4732
R553 VTAIL.n482 VTAIL.n481 10.4732
R554 VTAIL.n462 VTAIL.n461 10.4732
R555 VTAIL.n437 VTAIL.n420 10.4732
R556 VTAIL.n384 VTAIL.n383 10.4732
R557 VTAIL.n364 VTAIL.n363 10.4732
R558 VTAIL.n339 VTAIL.n322 10.4732
R559 VTAIL.n730 VTAIL.n710 9.69747
R560 VTAIL.n750 VTAIL.n700 9.69747
R561 VTAIL.n779 VTAIL.n688 9.69747
R562 VTAIL.n44 VTAIL.n24 9.69747
R563 VTAIL.n64 VTAIL.n14 9.69747
R564 VTAIL.n93 VTAIL.n2 9.69747
R565 VTAIL.n142 VTAIL.n122 9.69747
R566 VTAIL.n162 VTAIL.n112 9.69747
R567 VTAIL.n191 VTAIL.n100 9.69747
R568 VTAIL.n240 VTAIL.n220 9.69747
R569 VTAIL.n260 VTAIL.n210 9.69747
R570 VTAIL.n289 VTAIL.n198 9.69747
R571 VTAIL.n681 VTAIL.n590 9.69747
R572 VTAIL.n654 VTAIL.n604 9.69747
R573 VTAIL.n634 VTAIL.n614 9.69747
R574 VTAIL.n583 VTAIL.n492 9.69747
R575 VTAIL.n556 VTAIL.n506 9.69747
R576 VTAIL.n536 VTAIL.n516 9.69747
R577 VTAIL.n485 VTAIL.n394 9.69747
R578 VTAIL.n458 VTAIL.n408 9.69747
R579 VTAIL.n438 VTAIL.n418 9.69747
R580 VTAIL.n387 VTAIL.n296 9.69747
R581 VTAIL.n360 VTAIL.n310 9.69747
R582 VTAIL.n340 VTAIL.n320 9.69747
R583 VTAIL.n782 VTAIL.n781 9.45567
R584 VTAIL.n96 VTAIL.n95 9.45567
R585 VTAIL.n194 VTAIL.n193 9.45567
R586 VTAIL.n292 VTAIL.n291 9.45567
R587 VTAIL.n684 VTAIL.n683 9.45567
R588 VTAIL.n586 VTAIL.n585 9.45567
R589 VTAIL.n488 VTAIL.n487 9.45567
R590 VTAIL.n390 VTAIL.n389 9.45567
R591 VTAIL.n781 VTAIL.n780 9.3005
R592 VTAIL.n688 VTAIL.n687 9.3005
R593 VTAIL.n775 VTAIL.n774 9.3005
R594 VTAIL.n773 VTAIL.n772 9.3005
R595 VTAIL.n692 VTAIL.n691 9.3005
R596 VTAIL.n767 VTAIL.n766 9.3005
R597 VTAIL.n739 VTAIL.n738 9.3005
R598 VTAIL.n708 VTAIL.n707 9.3005
R599 VTAIL.n733 VTAIL.n732 9.3005
R600 VTAIL.n731 VTAIL.n730 9.3005
R601 VTAIL.n712 VTAIL.n711 9.3005
R602 VTAIL.n725 VTAIL.n724 9.3005
R603 VTAIL.n723 VTAIL.n722 9.3005
R604 VTAIL.n716 VTAIL.n715 9.3005
R605 VTAIL.n741 VTAIL.n740 9.3005
R606 VTAIL.n704 VTAIL.n703 9.3005
R607 VTAIL.n747 VTAIL.n746 9.3005
R608 VTAIL.n749 VTAIL.n748 9.3005
R609 VTAIL.n700 VTAIL.n699 9.3005
R610 VTAIL.n755 VTAIL.n754 9.3005
R611 VTAIL.n757 VTAIL.n756 9.3005
R612 VTAIL.n758 VTAIL.n695 9.3005
R613 VTAIL.n765 VTAIL.n764 9.3005
R614 VTAIL.n95 VTAIL.n94 9.3005
R615 VTAIL.n2 VTAIL.n1 9.3005
R616 VTAIL.n89 VTAIL.n88 9.3005
R617 VTAIL.n87 VTAIL.n86 9.3005
R618 VTAIL.n6 VTAIL.n5 9.3005
R619 VTAIL.n81 VTAIL.n80 9.3005
R620 VTAIL.n53 VTAIL.n52 9.3005
R621 VTAIL.n22 VTAIL.n21 9.3005
R622 VTAIL.n47 VTAIL.n46 9.3005
R623 VTAIL.n45 VTAIL.n44 9.3005
R624 VTAIL.n26 VTAIL.n25 9.3005
R625 VTAIL.n39 VTAIL.n38 9.3005
R626 VTAIL.n37 VTAIL.n36 9.3005
R627 VTAIL.n30 VTAIL.n29 9.3005
R628 VTAIL.n55 VTAIL.n54 9.3005
R629 VTAIL.n18 VTAIL.n17 9.3005
R630 VTAIL.n61 VTAIL.n60 9.3005
R631 VTAIL.n63 VTAIL.n62 9.3005
R632 VTAIL.n14 VTAIL.n13 9.3005
R633 VTAIL.n69 VTAIL.n68 9.3005
R634 VTAIL.n71 VTAIL.n70 9.3005
R635 VTAIL.n72 VTAIL.n9 9.3005
R636 VTAIL.n79 VTAIL.n78 9.3005
R637 VTAIL.n193 VTAIL.n192 9.3005
R638 VTAIL.n100 VTAIL.n99 9.3005
R639 VTAIL.n187 VTAIL.n186 9.3005
R640 VTAIL.n185 VTAIL.n184 9.3005
R641 VTAIL.n104 VTAIL.n103 9.3005
R642 VTAIL.n179 VTAIL.n178 9.3005
R643 VTAIL.n151 VTAIL.n150 9.3005
R644 VTAIL.n120 VTAIL.n119 9.3005
R645 VTAIL.n145 VTAIL.n144 9.3005
R646 VTAIL.n143 VTAIL.n142 9.3005
R647 VTAIL.n124 VTAIL.n123 9.3005
R648 VTAIL.n137 VTAIL.n136 9.3005
R649 VTAIL.n135 VTAIL.n134 9.3005
R650 VTAIL.n128 VTAIL.n127 9.3005
R651 VTAIL.n153 VTAIL.n152 9.3005
R652 VTAIL.n116 VTAIL.n115 9.3005
R653 VTAIL.n159 VTAIL.n158 9.3005
R654 VTAIL.n161 VTAIL.n160 9.3005
R655 VTAIL.n112 VTAIL.n111 9.3005
R656 VTAIL.n167 VTAIL.n166 9.3005
R657 VTAIL.n169 VTAIL.n168 9.3005
R658 VTAIL.n170 VTAIL.n107 9.3005
R659 VTAIL.n177 VTAIL.n176 9.3005
R660 VTAIL.n291 VTAIL.n290 9.3005
R661 VTAIL.n198 VTAIL.n197 9.3005
R662 VTAIL.n285 VTAIL.n284 9.3005
R663 VTAIL.n283 VTAIL.n282 9.3005
R664 VTAIL.n202 VTAIL.n201 9.3005
R665 VTAIL.n277 VTAIL.n276 9.3005
R666 VTAIL.n249 VTAIL.n248 9.3005
R667 VTAIL.n218 VTAIL.n217 9.3005
R668 VTAIL.n243 VTAIL.n242 9.3005
R669 VTAIL.n241 VTAIL.n240 9.3005
R670 VTAIL.n222 VTAIL.n221 9.3005
R671 VTAIL.n235 VTAIL.n234 9.3005
R672 VTAIL.n233 VTAIL.n232 9.3005
R673 VTAIL.n226 VTAIL.n225 9.3005
R674 VTAIL.n251 VTAIL.n250 9.3005
R675 VTAIL.n214 VTAIL.n213 9.3005
R676 VTAIL.n257 VTAIL.n256 9.3005
R677 VTAIL.n259 VTAIL.n258 9.3005
R678 VTAIL.n210 VTAIL.n209 9.3005
R679 VTAIL.n265 VTAIL.n264 9.3005
R680 VTAIL.n267 VTAIL.n266 9.3005
R681 VTAIL.n268 VTAIL.n205 9.3005
R682 VTAIL.n275 VTAIL.n274 9.3005
R683 VTAIL.n608 VTAIL.n607 9.3005
R684 VTAIL.n651 VTAIL.n650 9.3005
R685 VTAIL.n653 VTAIL.n652 9.3005
R686 VTAIL.n604 VTAIL.n603 9.3005
R687 VTAIL.n659 VTAIL.n658 9.3005
R688 VTAIL.n661 VTAIL.n660 9.3005
R689 VTAIL.n599 VTAIL.n597 9.3005
R690 VTAIL.n667 VTAIL.n666 9.3005
R691 VTAIL.n683 VTAIL.n682 9.3005
R692 VTAIL.n590 VTAIL.n589 9.3005
R693 VTAIL.n677 VTAIL.n676 9.3005
R694 VTAIL.n675 VTAIL.n674 9.3005
R695 VTAIL.n594 VTAIL.n593 9.3005
R696 VTAIL.n669 VTAIL.n668 9.3005
R697 VTAIL.n645 VTAIL.n644 9.3005
R698 VTAIL.n643 VTAIL.n642 9.3005
R699 VTAIL.n612 VTAIL.n611 9.3005
R700 VTAIL.n637 VTAIL.n636 9.3005
R701 VTAIL.n635 VTAIL.n634 9.3005
R702 VTAIL.n616 VTAIL.n615 9.3005
R703 VTAIL.n629 VTAIL.n628 9.3005
R704 VTAIL.n627 VTAIL.n626 9.3005
R705 VTAIL.n620 VTAIL.n619 9.3005
R706 VTAIL.n510 VTAIL.n509 9.3005
R707 VTAIL.n553 VTAIL.n552 9.3005
R708 VTAIL.n555 VTAIL.n554 9.3005
R709 VTAIL.n506 VTAIL.n505 9.3005
R710 VTAIL.n561 VTAIL.n560 9.3005
R711 VTAIL.n563 VTAIL.n562 9.3005
R712 VTAIL.n501 VTAIL.n499 9.3005
R713 VTAIL.n569 VTAIL.n568 9.3005
R714 VTAIL.n585 VTAIL.n584 9.3005
R715 VTAIL.n492 VTAIL.n491 9.3005
R716 VTAIL.n579 VTAIL.n578 9.3005
R717 VTAIL.n577 VTAIL.n576 9.3005
R718 VTAIL.n496 VTAIL.n495 9.3005
R719 VTAIL.n571 VTAIL.n570 9.3005
R720 VTAIL.n547 VTAIL.n546 9.3005
R721 VTAIL.n545 VTAIL.n544 9.3005
R722 VTAIL.n514 VTAIL.n513 9.3005
R723 VTAIL.n539 VTAIL.n538 9.3005
R724 VTAIL.n537 VTAIL.n536 9.3005
R725 VTAIL.n518 VTAIL.n517 9.3005
R726 VTAIL.n531 VTAIL.n530 9.3005
R727 VTAIL.n529 VTAIL.n528 9.3005
R728 VTAIL.n522 VTAIL.n521 9.3005
R729 VTAIL.n412 VTAIL.n411 9.3005
R730 VTAIL.n455 VTAIL.n454 9.3005
R731 VTAIL.n457 VTAIL.n456 9.3005
R732 VTAIL.n408 VTAIL.n407 9.3005
R733 VTAIL.n463 VTAIL.n462 9.3005
R734 VTAIL.n465 VTAIL.n464 9.3005
R735 VTAIL.n403 VTAIL.n401 9.3005
R736 VTAIL.n471 VTAIL.n470 9.3005
R737 VTAIL.n487 VTAIL.n486 9.3005
R738 VTAIL.n394 VTAIL.n393 9.3005
R739 VTAIL.n481 VTAIL.n480 9.3005
R740 VTAIL.n479 VTAIL.n478 9.3005
R741 VTAIL.n398 VTAIL.n397 9.3005
R742 VTAIL.n473 VTAIL.n472 9.3005
R743 VTAIL.n449 VTAIL.n448 9.3005
R744 VTAIL.n447 VTAIL.n446 9.3005
R745 VTAIL.n416 VTAIL.n415 9.3005
R746 VTAIL.n441 VTAIL.n440 9.3005
R747 VTAIL.n439 VTAIL.n438 9.3005
R748 VTAIL.n420 VTAIL.n419 9.3005
R749 VTAIL.n433 VTAIL.n432 9.3005
R750 VTAIL.n431 VTAIL.n430 9.3005
R751 VTAIL.n424 VTAIL.n423 9.3005
R752 VTAIL.n314 VTAIL.n313 9.3005
R753 VTAIL.n357 VTAIL.n356 9.3005
R754 VTAIL.n359 VTAIL.n358 9.3005
R755 VTAIL.n310 VTAIL.n309 9.3005
R756 VTAIL.n365 VTAIL.n364 9.3005
R757 VTAIL.n367 VTAIL.n366 9.3005
R758 VTAIL.n305 VTAIL.n303 9.3005
R759 VTAIL.n373 VTAIL.n372 9.3005
R760 VTAIL.n389 VTAIL.n388 9.3005
R761 VTAIL.n296 VTAIL.n295 9.3005
R762 VTAIL.n383 VTAIL.n382 9.3005
R763 VTAIL.n381 VTAIL.n380 9.3005
R764 VTAIL.n300 VTAIL.n299 9.3005
R765 VTAIL.n375 VTAIL.n374 9.3005
R766 VTAIL.n351 VTAIL.n350 9.3005
R767 VTAIL.n349 VTAIL.n348 9.3005
R768 VTAIL.n318 VTAIL.n317 9.3005
R769 VTAIL.n343 VTAIL.n342 9.3005
R770 VTAIL.n341 VTAIL.n340 9.3005
R771 VTAIL.n322 VTAIL.n321 9.3005
R772 VTAIL.n335 VTAIL.n334 9.3005
R773 VTAIL.n333 VTAIL.n332 9.3005
R774 VTAIL.n326 VTAIL.n325 9.3005
R775 VTAIL.n734 VTAIL.n733 8.92171
R776 VTAIL.n749 VTAIL.n702 8.92171
R777 VTAIL.n780 VTAIL.n686 8.92171
R778 VTAIL.n48 VTAIL.n47 8.92171
R779 VTAIL.n63 VTAIL.n16 8.92171
R780 VTAIL.n94 VTAIL.n0 8.92171
R781 VTAIL.n146 VTAIL.n145 8.92171
R782 VTAIL.n161 VTAIL.n114 8.92171
R783 VTAIL.n192 VTAIL.n98 8.92171
R784 VTAIL.n244 VTAIL.n243 8.92171
R785 VTAIL.n259 VTAIL.n212 8.92171
R786 VTAIL.n290 VTAIL.n196 8.92171
R787 VTAIL.n682 VTAIL.n588 8.92171
R788 VTAIL.n653 VTAIL.n606 8.92171
R789 VTAIL.n638 VTAIL.n637 8.92171
R790 VTAIL.n584 VTAIL.n490 8.92171
R791 VTAIL.n555 VTAIL.n508 8.92171
R792 VTAIL.n540 VTAIL.n539 8.92171
R793 VTAIL.n486 VTAIL.n392 8.92171
R794 VTAIL.n457 VTAIL.n410 8.92171
R795 VTAIL.n442 VTAIL.n441 8.92171
R796 VTAIL.n388 VTAIL.n294 8.92171
R797 VTAIL.n359 VTAIL.n312 8.92171
R798 VTAIL.n344 VTAIL.n343 8.92171
R799 VTAIL.n737 VTAIL.n708 8.14595
R800 VTAIL.n746 VTAIL.n745 8.14595
R801 VTAIL.n51 VTAIL.n22 8.14595
R802 VTAIL.n60 VTAIL.n59 8.14595
R803 VTAIL.n149 VTAIL.n120 8.14595
R804 VTAIL.n158 VTAIL.n157 8.14595
R805 VTAIL.n247 VTAIL.n218 8.14595
R806 VTAIL.n256 VTAIL.n255 8.14595
R807 VTAIL.n650 VTAIL.n649 8.14595
R808 VTAIL.n641 VTAIL.n612 8.14595
R809 VTAIL.n552 VTAIL.n551 8.14595
R810 VTAIL.n543 VTAIL.n514 8.14595
R811 VTAIL.n454 VTAIL.n453 8.14595
R812 VTAIL.n445 VTAIL.n416 8.14595
R813 VTAIL.n356 VTAIL.n355 8.14595
R814 VTAIL.n347 VTAIL.n318 8.14595
R815 VTAIL.n738 VTAIL.n706 7.3702
R816 VTAIL.n742 VTAIL.n704 7.3702
R817 VTAIL.n52 VTAIL.n20 7.3702
R818 VTAIL.n56 VTAIL.n18 7.3702
R819 VTAIL.n150 VTAIL.n118 7.3702
R820 VTAIL.n154 VTAIL.n116 7.3702
R821 VTAIL.n248 VTAIL.n216 7.3702
R822 VTAIL.n252 VTAIL.n214 7.3702
R823 VTAIL.n646 VTAIL.n608 7.3702
R824 VTAIL.n642 VTAIL.n610 7.3702
R825 VTAIL.n548 VTAIL.n510 7.3702
R826 VTAIL.n544 VTAIL.n512 7.3702
R827 VTAIL.n450 VTAIL.n412 7.3702
R828 VTAIL.n446 VTAIL.n414 7.3702
R829 VTAIL.n352 VTAIL.n314 7.3702
R830 VTAIL.n348 VTAIL.n316 7.3702
R831 VTAIL.n741 VTAIL.n706 6.59444
R832 VTAIL.n742 VTAIL.n741 6.59444
R833 VTAIL.n55 VTAIL.n20 6.59444
R834 VTAIL.n56 VTAIL.n55 6.59444
R835 VTAIL.n153 VTAIL.n118 6.59444
R836 VTAIL.n154 VTAIL.n153 6.59444
R837 VTAIL.n251 VTAIL.n216 6.59444
R838 VTAIL.n252 VTAIL.n251 6.59444
R839 VTAIL.n646 VTAIL.n645 6.59444
R840 VTAIL.n645 VTAIL.n610 6.59444
R841 VTAIL.n548 VTAIL.n547 6.59444
R842 VTAIL.n547 VTAIL.n512 6.59444
R843 VTAIL.n450 VTAIL.n449 6.59444
R844 VTAIL.n449 VTAIL.n414 6.59444
R845 VTAIL.n352 VTAIL.n351 6.59444
R846 VTAIL.n351 VTAIL.n316 6.59444
R847 VTAIL.n738 VTAIL.n737 5.81868
R848 VTAIL.n745 VTAIL.n704 5.81868
R849 VTAIL.n52 VTAIL.n51 5.81868
R850 VTAIL.n59 VTAIL.n18 5.81868
R851 VTAIL.n150 VTAIL.n149 5.81868
R852 VTAIL.n157 VTAIL.n116 5.81868
R853 VTAIL.n248 VTAIL.n247 5.81868
R854 VTAIL.n255 VTAIL.n214 5.81868
R855 VTAIL.n649 VTAIL.n608 5.81868
R856 VTAIL.n642 VTAIL.n641 5.81868
R857 VTAIL.n551 VTAIL.n510 5.81868
R858 VTAIL.n544 VTAIL.n543 5.81868
R859 VTAIL.n453 VTAIL.n412 5.81868
R860 VTAIL.n446 VTAIL.n445 5.81868
R861 VTAIL.n355 VTAIL.n314 5.81868
R862 VTAIL.n348 VTAIL.n347 5.81868
R863 VTAIL.n734 VTAIL.n708 5.04292
R864 VTAIL.n746 VTAIL.n702 5.04292
R865 VTAIL.n782 VTAIL.n686 5.04292
R866 VTAIL.n48 VTAIL.n22 5.04292
R867 VTAIL.n60 VTAIL.n16 5.04292
R868 VTAIL.n96 VTAIL.n0 5.04292
R869 VTAIL.n146 VTAIL.n120 5.04292
R870 VTAIL.n158 VTAIL.n114 5.04292
R871 VTAIL.n194 VTAIL.n98 5.04292
R872 VTAIL.n244 VTAIL.n218 5.04292
R873 VTAIL.n256 VTAIL.n212 5.04292
R874 VTAIL.n292 VTAIL.n196 5.04292
R875 VTAIL.n684 VTAIL.n588 5.04292
R876 VTAIL.n650 VTAIL.n606 5.04292
R877 VTAIL.n638 VTAIL.n612 5.04292
R878 VTAIL.n586 VTAIL.n490 5.04292
R879 VTAIL.n552 VTAIL.n508 5.04292
R880 VTAIL.n540 VTAIL.n514 5.04292
R881 VTAIL.n488 VTAIL.n392 5.04292
R882 VTAIL.n454 VTAIL.n410 5.04292
R883 VTAIL.n442 VTAIL.n416 5.04292
R884 VTAIL.n390 VTAIL.n294 5.04292
R885 VTAIL.n356 VTAIL.n312 5.04292
R886 VTAIL.n344 VTAIL.n318 5.04292
R887 VTAIL.n717 VTAIL.n715 4.38563
R888 VTAIL.n31 VTAIL.n29 4.38563
R889 VTAIL.n129 VTAIL.n127 4.38563
R890 VTAIL.n227 VTAIL.n225 4.38563
R891 VTAIL.n621 VTAIL.n619 4.38563
R892 VTAIL.n523 VTAIL.n521 4.38563
R893 VTAIL.n425 VTAIL.n423 4.38563
R894 VTAIL.n327 VTAIL.n325 4.38563
R895 VTAIL.n733 VTAIL.n710 4.26717
R896 VTAIL.n750 VTAIL.n749 4.26717
R897 VTAIL.n780 VTAIL.n779 4.26717
R898 VTAIL.n47 VTAIL.n24 4.26717
R899 VTAIL.n64 VTAIL.n63 4.26717
R900 VTAIL.n94 VTAIL.n93 4.26717
R901 VTAIL.n145 VTAIL.n122 4.26717
R902 VTAIL.n162 VTAIL.n161 4.26717
R903 VTAIL.n192 VTAIL.n191 4.26717
R904 VTAIL.n243 VTAIL.n220 4.26717
R905 VTAIL.n260 VTAIL.n259 4.26717
R906 VTAIL.n290 VTAIL.n289 4.26717
R907 VTAIL.n682 VTAIL.n681 4.26717
R908 VTAIL.n654 VTAIL.n653 4.26717
R909 VTAIL.n637 VTAIL.n614 4.26717
R910 VTAIL.n584 VTAIL.n583 4.26717
R911 VTAIL.n556 VTAIL.n555 4.26717
R912 VTAIL.n539 VTAIL.n516 4.26717
R913 VTAIL.n486 VTAIL.n485 4.26717
R914 VTAIL.n458 VTAIL.n457 4.26717
R915 VTAIL.n441 VTAIL.n418 4.26717
R916 VTAIL.n388 VTAIL.n387 4.26717
R917 VTAIL.n360 VTAIL.n359 4.26717
R918 VTAIL.n343 VTAIL.n320 4.26717
R919 VTAIL.n730 VTAIL.n729 3.49141
R920 VTAIL.n753 VTAIL.n700 3.49141
R921 VTAIL.n776 VTAIL.n688 3.49141
R922 VTAIL.n44 VTAIL.n43 3.49141
R923 VTAIL.n67 VTAIL.n14 3.49141
R924 VTAIL.n90 VTAIL.n2 3.49141
R925 VTAIL.n142 VTAIL.n141 3.49141
R926 VTAIL.n165 VTAIL.n112 3.49141
R927 VTAIL.n188 VTAIL.n100 3.49141
R928 VTAIL.n240 VTAIL.n239 3.49141
R929 VTAIL.n263 VTAIL.n210 3.49141
R930 VTAIL.n286 VTAIL.n198 3.49141
R931 VTAIL.n678 VTAIL.n590 3.49141
R932 VTAIL.n657 VTAIL.n604 3.49141
R933 VTAIL.n634 VTAIL.n633 3.49141
R934 VTAIL.n580 VTAIL.n492 3.49141
R935 VTAIL.n559 VTAIL.n506 3.49141
R936 VTAIL.n536 VTAIL.n535 3.49141
R937 VTAIL.n482 VTAIL.n394 3.49141
R938 VTAIL.n461 VTAIL.n408 3.49141
R939 VTAIL.n438 VTAIL.n437 3.49141
R940 VTAIL.n384 VTAIL.n296 3.49141
R941 VTAIL.n363 VTAIL.n310 3.49141
R942 VTAIL.n340 VTAIL.n339 3.49141
R943 VTAIL.n489 VTAIL.n391 2.73326
R944 VTAIL.n685 VTAIL.n587 2.73326
R945 VTAIL.n293 VTAIL.n195 2.73326
R946 VTAIL.n726 VTAIL.n712 2.71565
R947 VTAIL.n754 VTAIL.n698 2.71565
R948 VTAIL.n775 VTAIL.n690 2.71565
R949 VTAIL.n40 VTAIL.n26 2.71565
R950 VTAIL.n68 VTAIL.n12 2.71565
R951 VTAIL.n89 VTAIL.n4 2.71565
R952 VTAIL.n138 VTAIL.n124 2.71565
R953 VTAIL.n166 VTAIL.n110 2.71565
R954 VTAIL.n187 VTAIL.n102 2.71565
R955 VTAIL.n236 VTAIL.n222 2.71565
R956 VTAIL.n264 VTAIL.n208 2.71565
R957 VTAIL.n285 VTAIL.n200 2.71565
R958 VTAIL.n677 VTAIL.n592 2.71565
R959 VTAIL.n658 VTAIL.n602 2.71565
R960 VTAIL.n630 VTAIL.n616 2.71565
R961 VTAIL.n579 VTAIL.n494 2.71565
R962 VTAIL.n560 VTAIL.n504 2.71565
R963 VTAIL.n532 VTAIL.n518 2.71565
R964 VTAIL.n481 VTAIL.n396 2.71565
R965 VTAIL.n462 VTAIL.n406 2.71565
R966 VTAIL.n434 VTAIL.n420 2.71565
R967 VTAIL.n383 VTAIL.n298 2.71565
R968 VTAIL.n364 VTAIL.n308 2.71565
R969 VTAIL.n336 VTAIL.n322 2.71565
R970 VTAIL.n725 VTAIL.n714 1.93989
R971 VTAIL.n759 VTAIL.n757 1.93989
R972 VTAIL.n772 VTAIL.n771 1.93989
R973 VTAIL.n39 VTAIL.n28 1.93989
R974 VTAIL.n73 VTAIL.n71 1.93989
R975 VTAIL.n86 VTAIL.n85 1.93989
R976 VTAIL.n137 VTAIL.n126 1.93989
R977 VTAIL.n171 VTAIL.n169 1.93989
R978 VTAIL.n184 VTAIL.n183 1.93989
R979 VTAIL.n235 VTAIL.n224 1.93989
R980 VTAIL.n269 VTAIL.n267 1.93989
R981 VTAIL.n282 VTAIL.n281 1.93989
R982 VTAIL.n674 VTAIL.n673 1.93989
R983 VTAIL.n662 VTAIL.n661 1.93989
R984 VTAIL.n629 VTAIL.n618 1.93989
R985 VTAIL.n576 VTAIL.n575 1.93989
R986 VTAIL.n564 VTAIL.n563 1.93989
R987 VTAIL.n531 VTAIL.n520 1.93989
R988 VTAIL.n478 VTAIL.n477 1.93989
R989 VTAIL.n466 VTAIL.n465 1.93989
R990 VTAIL.n433 VTAIL.n422 1.93989
R991 VTAIL.n380 VTAIL.n379 1.93989
R992 VTAIL.n368 VTAIL.n367 1.93989
R993 VTAIL.n335 VTAIL.n324 1.93989
R994 VTAIL VTAIL.n97 1.42507
R995 VTAIL VTAIL.n783 1.30869
R996 VTAIL.n722 VTAIL.n721 1.16414
R997 VTAIL.n758 VTAIL.n696 1.16414
R998 VTAIL.n768 VTAIL.n692 1.16414
R999 VTAIL.n36 VTAIL.n35 1.16414
R1000 VTAIL.n72 VTAIL.n10 1.16414
R1001 VTAIL.n82 VTAIL.n6 1.16414
R1002 VTAIL.n134 VTAIL.n133 1.16414
R1003 VTAIL.n170 VTAIL.n108 1.16414
R1004 VTAIL.n180 VTAIL.n104 1.16414
R1005 VTAIL.n232 VTAIL.n231 1.16414
R1006 VTAIL.n268 VTAIL.n206 1.16414
R1007 VTAIL.n278 VTAIL.n202 1.16414
R1008 VTAIL.n670 VTAIL.n594 1.16414
R1009 VTAIL.n665 VTAIL.n599 1.16414
R1010 VTAIL.n626 VTAIL.n625 1.16414
R1011 VTAIL.n572 VTAIL.n496 1.16414
R1012 VTAIL.n567 VTAIL.n501 1.16414
R1013 VTAIL.n528 VTAIL.n527 1.16414
R1014 VTAIL.n474 VTAIL.n398 1.16414
R1015 VTAIL.n469 VTAIL.n403 1.16414
R1016 VTAIL.n430 VTAIL.n429 1.16414
R1017 VTAIL.n376 VTAIL.n300 1.16414
R1018 VTAIL.n371 VTAIL.n305 1.16414
R1019 VTAIL.n332 VTAIL.n331 1.16414
R1020 VTAIL.n587 VTAIL.n489 0.470328
R1021 VTAIL.n195 VTAIL.n97 0.470328
R1022 VTAIL.n718 VTAIL.n716 0.388379
R1023 VTAIL.n764 VTAIL.n763 0.388379
R1024 VTAIL.n767 VTAIL.n694 0.388379
R1025 VTAIL.n32 VTAIL.n30 0.388379
R1026 VTAIL.n78 VTAIL.n77 0.388379
R1027 VTAIL.n81 VTAIL.n8 0.388379
R1028 VTAIL.n130 VTAIL.n128 0.388379
R1029 VTAIL.n176 VTAIL.n175 0.388379
R1030 VTAIL.n179 VTAIL.n106 0.388379
R1031 VTAIL.n228 VTAIL.n226 0.388379
R1032 VTAIL.n274 VTAIL.n273 0.388379
R1033 VTAIL.n277 VTAIL.n204 0.388379
R1034 VTAIL.n669 VTAIL.n596 0.388379
R1035 VTAIL.n666 VTAIL.n598 0.388379
R1036 VTAIL.n622 VTAIL.n620 0.388379
R1037 VTAIL.n571 VTAIL.n498 0.388379
R1038 VTAIL.n568 VTAIL.n500 0.388379
R1039 VTAIL.n524 VTAIL.n522 0.388379
R1040 VTAIL.n473 VTAIL.n400 0.388379
R1041 VTAIL.n470 VTAIL.n402 0.388379
R1042 VTAIL.n426 VTAIL.n424 0.388379
R1043 VTAIL.n375 VTAIL.n302 0.388379
R1044 VTAIL.n372 VTAIL.n304 0.388379
R1045 VTAIL.n328 VTAIL.n326 0.388379
R1046 VTAIL.n723 VTAIL.n715 0.155672
R1047 VTAIL.n724 VTAIL.n723 0.155672
R1048 VTAIL.n724 VTAIL.n711 0.155672
R1049 VTAIL.n731 VTAIL.n711 0.155672
R1050 VTAIL.n732 VTAIL.n731 0.155672
R1051 VTAIL.n732 VTAIL.n707 0.155672
R1052 VTAIL.n739 VTAIL.n707 0.155672
R1053 VTAIL.n740 VTAIL.n739 0.155672
R1054 VTAIL.n740 VTAIL.n703 0.155672
R1055 VTAIL.n747 VTAIL.n703 0.155672
R1056 VTAIL.n748 VTAIL.n747 0.155672
R1057 VTAIL.n748 VTAIL.n699 0.155672
R1058 VTAIL.n755 VTAIL.n699 0.155672
R1059 VTAIL.n756 VTAIL.n755 0.155672
R1060 VTAIL.n756 VTAIL.n695 0.155672
R1061 VTAIL.n765 VTAIL.n695 0.155672
R1062 VTAIL.n766 VTAIL.n765 0.155672
R1063 VTAIL.n766 VTAIL.n691 0.155672
R1064 VTAIL.n773 VTAIL.n691 0.155672
R1065 VTAIL.n774 VTAIL.n773 0.155672
R1066 VTAIL.n774 VTAIL.n687 0.155672
R1067 VTAIL.n781 VTAIL.n687 0.155672
R1068 VTAIL.n37 VTAIL.n29 0.155672
R1069 VTAIL.n38 VTAIL.n37 0.155672
R1070 VTAIL.n38 VTAIL.n25 0.155672
R1071 VTAIL.n45 VTAIL.n25 0.155672
R1072 VTAIL.n46 VTAIL.n45 0.155672
R1073 VTAIL.n46 VTAIL.n21 0.155672
R1074 VTAIL.n53 VTAIL.n21 0.155672
R1075 VTAIL.n54 VTAIL.n53 0.155672
R1076 VTAIL.n54 VTAIL.n17 0.155672
R1077 VTAIL.n61 VTAIL.n17 0.155672
R1078 VTAIL.n62 VTAIL.n61 0.155672
R1079 VTAIL.n62 VTAIL.n13 0.155672
R1080 VTAIL.n69 VTAIL.n13 0.155672
R1081 VTAIL.n70 VTAIL.n69 0.155672
R1082 VTAIL.n70 VTAIL.n9 0.155672
R1083 VTAIL.n79 VTAIL.n9 0.155672
R1084 VTAIL.n80 VTAIL.n79 0.155672
R1085 VTAIL.n80 VTAIL.n5 0.155672
R1086 VTAIL.n87 VTAIL.n5 0.155672
R1087 VTAIL.n88 VTAIL.n87 0.155672
R1088 VTAIL.n88 VTAIL.n1 0.155672
R1089 VTAIL.n95 VTAIL.n1 0.155672
R1090 VTAIL.n135 VTAIL.n127 0.155672
R1091 VTAIL.n136 VTAIL.n135 0.155672
R1092 VTAIL.n136 VTAIL.n123 0.155672
R1093 VTAIL.n143 VTAIL.n123 0.155672
R1094 VTAIL.n144 VTAIL.n143 0.155672
R1095 VTAIL.n144 VTAIL.n119 0.155672
R1096 VTAIL.n151 VTAIL.n119 0.155672
R1097 VTAIL.n152 VTAIL.n151 0.155672
R1098 VTAIL.n152 VTAIL.n115 0.155672
R1099 VTAIL.n159 VTAIL.n115 0.155672
R1100 VTAIL.n160 VTAIL.n159 0.155672
R1101 VTAIL.n160 VTAIL.n111 0.155672
R1102 VTAIL.n167 VTAIL.n111 0.155672
R1103 VTAIL.n168 VTAIL.n167 0.155672
R1104 VTAIL.n168 VTAIL.n107 0.155672
R1105 VTAIL.n177 VTAIL.n107 0.155672
R1106 VTAIL.n178 VTAIL.n177 0.155672
R1107 VTAIL.n178 VTAIL.n103 0.155672
R1108 VTAIL.n185 VTAIL.n103 0.155672
R1109 VTAIL.n186 VTAIL.n185 0.155672
R1110 VTAIL.n186 VTAIL.n99 0.155672
R1111 VTAIL.n193 VTAIL.n99 0.155672
R1112 VTAIL.n233 VTAIL.n225 0.155672
R1113 VTAIL.n234 VTAIL.n233 0.155672
R1114 VTAIL.n234 VTAIL.n221 0.155672
R1115 VTAIL.n241 VTAIL.n221 0.155672
R1116 VTAIL.n242 VTAIL.n241 0.155672
R1117 VTAIL.n242 VTAIL.n217 0.155672
R1118 VTAIL.n249 VTAIL.n217 0.155672
R1119 VTAIL.n250 VTAIL.n249 0.155672
R1120 VTAIL.n250 VTAIL.n213 0.155672
R1121 VTAIL.n257 VTAIL.n213 0.155672
R1122 VTAIL.n258 VTAIL.n257 0.155672
R1123 VTAIL.n258 VTAIL.n209 0.155672
R1124 VTAIL.n265 VTAIL.n209 0.155672
R1125 VTAIL.n266 VTAIL.n265 0.155672
R1126 VTAIL.n266 VTAIL.n205 0.155672
R1127 VTAIL.n275 VTAIL.n205 0.155672
R1128 VTAIL.n276 VTAIL.n275 0.155672
R1129 VTAIL.n276 VTAIL.n201 0.155672
R1130 VTAIL.n283 VTAIL.n201 0.155672
R1131 VTAIL.n284 VTAIL.n283 0.155672
R1132 VTAIL.n284 VTAIL.n197 0.155672
R1133 VTAIL.n291 VTAIL.n197 0.155672
R1134 VTAIL.n683 VTAIL.n589 0.155672
R1135 VTAIL.n676 VTAIL.n589 0.155672
R1136 VTAIL.n676 VTAIL.n675 0.155672
R1137 VTAIL.n675 VTAIL.n593 0.155672
R1138 VTAIL.n668 VTAIL.n593 0.155672
R1139 VTAIL.n668 VTAIL.n667 0.155672
R1140 VTAIL.n667 VTAIL.n597 0.155672
R1141 VTAIL.n660 VTAIL.n597 0.155672
R1142 VTAIL.n660 VTAIL.n659 0.155672
R1143 VTAIL.n659 VTAIL.n603 0.155672
R1144 VTAIL.n652 VTAIL.n603 0.155672
R1145 VTAIL.n652 VTAIL.n651 0.155672
R1146 VTAIL.n651 VTAIL.n607 0.155672
R1147 VTAIL.n644 VTAIL.n607 0.155672
R1148 VTAIL.n644 VTAIL.n643 0.155672
R1149 VTAIL.n643 VTAIL.n611 0.155672
R1150 VTAIL.n636 VTAIL.n611 0.155672
R1151 VTAIL.n636 VTAIL.n635 0.155672
R1152 VTAIL.n635 VTAIL.n615 0.155672
R1153 VTAIL.n628 VTAIL.n615 0.155672
R1154 VTAIL.n628 VTAIL.n627 0.155672
R1155 VTAIL.n627 VTAIL.n619 0.155672
R1156 VTAIL.n585 VTAIL.n491 0.155672
R1157 VTAIL.n578 VTAIL.n491 0.155672
R1158 VTAIL.n578 VTAIL.n577 0.155672
R1159 VTAIL.n577 VTAIL.n495 0.155672
R1160 VTAIL.n570 VTAIL.n495 0.155672
R1161 VTAIL.n570 VTAIL.n569 0.155672
R1162 VTAIL.n569 VTAIL.n499 0.155672
R1163 VTAIL.n562 VTAIL.n499 0.155672
R1164 VTAIL.n562 VTAIL.n561 0.155672
R1165 VTAIL.n561 VTAIL.n505 0.155672
R1166 VTAIL.n554 VTAIL.n505 0.155672
R1167 VTAIL.n554 VTAIL.n553 0.155672
R1168 VTAIL.n553 VTAIL.n509 0.155672
R1169 VTAIL.n546 VTAIL.n509 0.155672
R1170 VTAIL.n546 VTAIL.n545 0.155672
R1171 VTAIL.n545 VTAIL.n513 0.155672
R1172 VTAIL.n538 VTAIL.n513 0.155672
R1173 VTAIL.n538 VTAIL.n537 0.155672
R1174 VTAIL.n537 VTAIL.n517 0.155672
R1175 VTAIL.n530 VTAIL.n517 0.155672
R1176 VTAIL.n530 VTAIL.n529 0.155672
R1177 VTAIL.n529 VTAIL.n521 0.155672
R1178 VTAIL.n487 VTAIL.n393 0.155672
R1179 VTAIL.n480 VTAIL.n393 0.155672
R1180 VTAIL.n480 VTAIL.n479 0.155672
R1181 VTAIL.n479 VTAIL.n397 0.155672
R1182 VTAIL.n472 VTAIL.n397 0.155672
R1183 VTAIL.n472 VTAIL.n471 0.155672
R1184 VTAIL.n471 VTAIL.n401 0.155672
R1185 VTAIL.n464 VTAIL.n401 0.155672
R1186 VTAIL.n464 VTAIL.n463 0.155672
R1187 VTAIL.n463 VTAIL.n407 0.155672
R1188 VTAIL.n456 VTAIL.n407 0.155672
R1189 VTAIL.n456 VTAIL.n455 0.155672
R1190 VTAIL.n455 VTAIL.n411 0.155672
R1191 VTAIL.n448 VTAIL.n411 0.155672
R1192 VTAIL.n448 VTAIL.n447 0.155672
R1193 VTAIL.n447 VTAIL.n415 0.155672
R1194 VTAIL.n440 VTAIL.n415 0.155672
R1195 VTAIL.n440 VTAIL.n439 0.155672
R1196 VTAIL.n439 VTAIL.n419 0.155672
R1197 VTAIL.n432 VTAIL.n419 0.155672
R1198 VTAIL.n432 VTAIL.n431 0.155672
R1199 VTAIL.n431 VTAIL.n423 0.155672
R1200 VTAIL.n389 VTAIL.n295 0.155672
R1201 VTAIL.n382 VTAIL.n295 0.155672
R1202 VTAIL.n382 VTAIL.n381 0.155672
R1203 VTAIL.n381 VTAIL.n299 0.155672
R1204 VTAIL.n374 VTAIL.n299 0.155672
R1205 VTAIL.n374 VTAIL.n373 0.155672
R1206 VTAIL.n373 VTAIL.n303 0.155672
R1207 VTAIL.n366 VTAIL.n303 0.155672
R1208 VTAIL.n366 VTAIL.n365 0.155672
R1209 VTAIL.n365 VTAIL.n309 0.155672
R1210 VTAIL.n358 VTAIL.n309 0.155672
R1211 VTAIL.n358 VTAIL.n357 0.155672
R1212 VTAIL.n357 VTAIL.n313 0.155672
R1213 VTAIL.n350 VTAIL.n313 0.155672
R1214 VTAIL.n350 VTAIL.n349 0.155672
R1215 VTAIL.n349 VTAIL.n317 0.155672
R1216 VTAIL.n342 VTAIL.n317 0.155672
R1217 VTAIL.n342 VTAIL.n341 0.155672
R1218 VTAIL.n341 VTAIL.n321 0.155672
R1219 VTAIL.n334 VTAIL.n321 0.155672
R1220 VTAIL.n334 VTAIL.n333 0.155672
R1221 VTAIL.n333 VTAIL.n325 0.155672
R1222 B.n930 B.n929 585
R1223 B.n384 B.n131 585
R1224 B.n383 B.n382 585
R1225 B.n381 B.n380 585
R1226 B.n379 B.n378 585
R1227 B.n377 B.n376 585
R1228 B.n375 B.n374 585
R1229 B.n373 B.n372 585
R1230 B.n371 B.n370 585
R1231 B.n369 B.n368 585
R1232 B.n367 B.n366 585
R1233 B.n365 B.n364 585
R1234 B.n363 B.n362 585
R1235 B.n361 B.n360 585
R1236 B.n359 B.n358 585
R1237 B.n357 B.n356 585
R1238 B.n355 B.n354 585
R1239 B.n353 B.n352 585
R1240 B.n351 B.n350 585
R1241 B.n349 B.n348 585
R1242 B.n347 B.n346 585
R1243 B.n345 B.n344 585
R1244 B.n343 B.n342 585
R1245 B.n341 B.n340 585
R1246 B.n339 B.n338 585
R1247 B.n337 B.n336 585
R1248 B.n335 B.n334 585
R1249 B.n333 B.n332 585
R1250 B.n331 B.n330 585
R1251 B.n329 B.n328 585
R1252 B.n327 B.n326 585
R1253 B.n325 B.n324 585
R1254 B.n323 B.n322 585
R1255 B.n321 B.n320 585
R1256 B.n319 B.n318 585
R1257 B.n317 B.n316 585
R1258 B.n315 B.n314 585
R1259 B.n313 B.n312 585
R1260 B.n311 B.n310 585
R1261 B.n309 B.n308 585
R1262 B.n307 B.n306 585
R1263 B.n305 B.n304 585
R1264 B.n303 B.n302 585
R1265 B.n301 B.n300 585
R1266 B.n299 B.n298 585
R1267 B.n297 B.n296 585
R1268 B.n295 B.n294 585
R1269 B.n293 B.n292 585
R1270 B.n291 B.n290 585
R1271 B.n289 B.n288 585
R1272 B.n287 B.n286 585
R1273 B.n285 B.n284 585
R1274 B.n283 B.n282 585
R1275 B.n281 B.n280 585
R1276 B.n279 B.n278 585
R1277 B.n277 B.n276 585
R1278 B.n275 B.n274 585
R1279 B.n273 B.n272 585
R1280 B.n271 B.n270 585
R1281 B.n269 B.n268 585
R1282 B.n267 B.n266 585
R1283 B.n265 B.n264 585
R1284 B.n263 B.n262 585
R1285 B.n261 B.n260 585
R1286 B.n259 B.n258 585
R1287 B.n257 B.n256 585
R1288 B.n255 B.n254 585
R1289 B.n253 B.n252 585
R1290 B.n251 B.n250 585
R1291 B.n249 B.n248 585
R1292 B.n247 B.n246 585
R1293 B.n245 B.n244 585
R1294 B.n243 B.n242 585
R1295 B.n241 B.n240 585
R1296 B.n239 B.n238 585
R1297 B.n237 B.n236 585
R1298 B.n235 B.n234 585
R1299 B.n233 B.n232 585
R1300 B.n231 B.n230 585
R1301 B.n229 B.n228 585
R1302 B.n227 B.n226 585
R1303 B.n225 B.n224 585
R1304 B.n223 B.n222 585
R1305 B.n221 B.n220 585
R1306 B.n219 B.n218 585
R1307 B.n217 B.n216 585
R1308 B.n215 B.n214 585
R1309 B.n213 B.n212 585
R1310 B.n211 B.n210 585
R1311 B.n209 B.n208 585
R1312 B.n207 B.n206 585
R1313 B.n205 B.n204 585
R1314 B.n203 B.n202 585
R1315 B.n201 B.n200 585
R1316 B.n199 B.n198 585
R1317 B.n197 B.n196 585
R1318 B.n195 B.n194 585
R1319 B.n193 B.n192 585
R1320 B.n191 B.n190 585
R1321 B.n189 B.n188 585
R1322 B.n187 B.n186 585
R1323 B.n185 B.n184 585
R1324 B.n183 B.n182 585
R1325 B.n181 B.n180 585
R1326 B.n179 B.n178 585
R1327 B.n177 B.n176 585
R1328 B.n175 B.n174 585
R1329 B.n173 B.n172 585
R1330 B.n171 B.n170 585
R1331 B.n169 B.n168 585
R1332 B.n167 B.n166 585
R1333 B.n165 B.n164 585
R1334 B.n163 B.n162 585
R1335 B.n161 B.n160 585
R1336 B.n159 B.n158 585
R1337 B.n157 B.n156 585
R1338 B.n155 B.n154 585
R1339 B.n153 B.n152 585
R1340 B.n151 B.n150 585
R1341 B.n149 B.n148 585
R1342 B.n147 B.n146 585
R1343 B.n145 B.n144 585
R1344 B.n143 B.n142 585
R1345 B.n141 B.n140 585
R1346 B.n139 B.n138 585
R1347 B.n67 B.n66 585
R1348 B.n928 B.n68 585
R1349 B.n933 B.n68 585
R1350 B.n927 B.n926 585
R1351 B.n926 B.n64 585
R1352 B.n925 B.n63 585
R1353 B.n939 B.n63 585
R1354 B.n924 B.n62 585
R1355 B.n940 B.n62 585
R1356 B.n923 B.n61 585
R1357 B.n941 B.n61 585
R1358 B.n922 B.n921 585
R1359 B.n921 B.n57 585
R1360 B.n920 B.n56 585
R1361 B.n947 B.n56 585
R1362 B.n919 B.n55 585
R1363 B.n948 B.n55 585
R1364 B.n918 B.n54 585
R1365 B.n949 B.n54 585
R1366 B.n917 B.n916 585
R1367 B.n916 B.n50 585
R1368 B.n915 B.n49 585
R1369 B.n955 B.n49 585
R1370 B.n914 B.n48 585
R1371 B.n956 B.n48 585
R1372 B.n913 B.n47 585
R1373 B.n957 B.n47 585
R1374 B.n912 B.n911 585
R1375 B.n911 B.n43 585
R1376 B.n910 B.n42 585
R1377 B.n963 B.n42 585
R1378 B.n909 B.n41 585
R1379 B.n964 B.n41 585
R1380 B.n908 B.n40 585
R1381 B.n965 B.n40 585
R1382 B.n907 B.n906 585
R1383 B.n906 B.n36 585
R1384 B.n905 B.n35 585
R1385 B.n971 B.n35 585
R1386 B.n904 B.n34 585
R1387 B.n972 B.n34 585
R1388 B.n903 B.n33 585
R1389 B.n973 B.n33 585
R1390 B.n902 B.n901 585
R1391 B.n901 B.n29 585
R1392 B.n900 B.n28 585
R1393 B.n979 B.n28 585
R1394 B.n899 B.n27 585
R1395 B.n980 B.n27 585
R1396 B.n898 B.n26 585
R1397 B.n981 B.n26 585
R1398 B.n897 B.n896 585
R1399 B.n896 B.n22 585
R1400 B.n895 B.n21 585
R1401 B.n987 B.n21 585
R1402 B.n894 B.n20 585
R1403 B.n988 B.n20 585
R1404 B.n893 B.n19 585
R1405 B.n989 B.n19 585
R1406 B.n892 B.n891 585
R1407 B.n891 B.n18 585
R1408 B.n890 B.n14 585
R1409 B.n995 B.n14 585
R1410 B.n889 B.n13 585
R1411 B.n996 B.n13 585
R1412 B.n888 B.n12 585
R1413 B.n997 B.n12 585
R1414 B.n887 B.n886 585
R1415 B.n886 B.n8 585
R1416 B.n885 B.n7 585
R1417 B.n1003 B.n7 585
R1418 B.n884 B.n6 585
R1419 B.n1004 B.n6 585
R1420 B.n883 B.n5 585
R1421 B.n1005 B.n5 585
R1422 B.n882 B.n881 585
R1423 B.n881 B.n4 585
R1424 B.n880 B.n385 585
R1425 B.n880 B.n879 585
R1426 B.n870 B.n386 585
R1427 B.n387 B.n386 585
R1428 B.n872 B.n871 585
R1429 B.n873 B.n872 585
R1430 B.n869 B.n392 585
R1431 B.n392 B.n391 585
R1432 B.n868 B.n867 585
R1433 B.n867 B.n866 585
R1434 B.n394 B.n393 585
R1435 B.n859 B.n394 585
R1436 B.n858 B.n857 585
R1437 B.n860 B.n858 585
R1438 B.n856 B.n399 585
R1439 B.n399 B.n398 585
R1440 B.n855 B.n854 585
R1441 B.n854 B.n853 585
R1442 B.n401 B.n400 585
R1443 B.n402 B.n401 585
R1444 B.n846 B.n845 585
R1445 B.n847 B.n846 585
R1446 B.n844 B.n407 585
R1447 B.n407 B.n406 585
R1448 B.n843 B.n842 585
R1449 B.n842 B.n841 585
R1450 B.n409 B.n408 585
R1451 B.n410 B.n409 585
R1452 B.n834 B.n833 585
R1453 B.n835 B.n834 585
R1454 B.n832 B.n415 585
R1455 B.n415 B.n414 585
R1456 B.n831 B.n830 585
R1457 B.n830 B.n829 585
R1458 B.n417 B.n416 585
R1459 B.n418 B.n417 585
R1460 B.n822 B.n821 585
R1461 B.n823 B.n822 585
R1462 B.n820 B.n423 585
R1463 B.n423 B.n422 585
R1464 B.n819 B.n818 585
R1465 B.n818 B.n817 585
R1466 B.n425 B.n424 585
R1467 B.n426 B.n425 585
R1468 B.n810 B.n809 585
R1469 B.n811 B.n810 585
R1470 B.n808 B.n431 585
R1471 B.n431 B.n430 585
R1472 B.n807 B.n806 585
R1473 B.n806 B.n805 585
R1474 B.n433 B.n432 585
R1475 B.n434 B.n433 585
R1476 B.n798 B.n797 585
R1477 B.n799 B.n798 585
R1478 B.n796 B.n438 585
R1479 B.n442 B.n438 585
R1480 B.n795 B.n794 585
R1481 B.n794 B.n793 585
R1482 B.n440 B.n439 585
R1483 B.n441 B.n440 585
R1484 B.n786 B.n785 585
R1485 B.n787 B.n786 585
R1486 B.n784 B.n447 585
R1487 B.n447 B.n446 585
R1488 B.n783 B.n782 585
R1489 B.n782 B.n781 585
R1490 B.n449 B.n448 585
R1491 B.n450 B.n449 585
R1492 B.n774 B.n773 585
R1493 B.n775 B.n774 585
R1494 B.n453 B.n452 585
R1495 B.n522 B.n520 585
R1496 B.n523 B.n519 585
R1497 B.n523 B.n454 585
R1498 B.n526 B.n525 585
R1499 B.n527 B.n518 585
R1500 B.n529 B.n528 585
R1501 B.n531 B.n517 585
R1502 B.n534 B.n533 585
R1503 B.n535 B.n516 585
R1504 B.n537 B.n536 585
R1505 B.n539 B.n515 585
R1506 B.n542 B.n541 585
R1507 B.n543 B.n514 585
R1508 B.n545 B.n544 585
R1509 B.n547 B.n513 585
R1510 B.n550 B.n549 585
R1511 B.n551 B.n512 585
R1512 B.n553 B.n552 585
R1513 B.n555 B.n511 585
R1514 B.n558 B.n557 585
R1515 B.n559 B.n510 585
R1516 B.n561 B.n560 585
R1517 B.n563 B.n509 585
R1518 B.n566 B.n565 585
R1519 B.n567 B.n508 585
R1520 B.n569 B.n568 585
R1521 B.n571 B.n507 585
R1522 B.n574 B.n573 585
R1523 B.n575 B.n506 585
R1524 B.n577 B.n576 585
R1525 B.n579 B.n505 585
R1526 B.n582 B.n581 585
R1527 B.n583 B.n504 585
R1528 B.n585 B.n584 585
R1529 B.n587 B.n503 585
R1530 B.n590 B.n589 585
R1531 B.n591 B.n502 585
R1532 B.n593 B.n592 585
R1533 B.n595 B.n501 585
R1534 B.n598 B.n597 585
R1535 B.n599 B.n500 585
R1536 B.n601 B.n600 585
R1537 B.n603 B.n499 585
R1538 B.n606 B.n605 585
R1539 B.n607 B.n498 585
R1540 B.n609 B.n608 585
R1541 B.n611 B.n497 585
R1542 B.n614 B.n613 585
R1543 B.n615 B.n496 585
R1544 B.n617 B.n616 585
R1545 B.n619 B.n495 585
R1546 B.n622 B.n621 585
R1547 B.n623 B.n494 585
R1548 B.n625 B.n624 585
R1549 B.n627 B.n493 585
R1550 B.n630 B.n629 585
R1551 B.n631 B.n492 585
R1552 B.n636 B.n635 585
R1553 B.n638 B.n491 585
R1554 B.n641 B.n640 585
R1555 B.n642 B.n490 585
R1556 B.n644 B.n643 585
R1557 B.n646 B.n489 585
R1558 B.n649 B.n648 585
R1559 B.n650 B.n488 585
R1560 B.n652 B.n651 585
R1561 B.n654 B.n487 585
R1562 B.n657 B.n656 585
R1563 B.n659 B.n484 585
R1564 B.n661 B.n660 585
R1565 B.n663 B.n483 585
R1566 B.n666 B.n665 585
R1567 B.n667 B.n482 585
R1568 B.n669 B.n668 585
R1569 B.n671 B.n481 585
R1570 B.n674 B.n673 585
R1571 B.n675 B.n480 585
R1572 B.n677 B.n676 585
R1573 B.n679 B.n479 585
R1574 B.n682 B.n681 585
R1575 B.n683 B.n478 585
R1576 B.n685 B.n684 585
R1577 B.n687 B.n477 585
R1578 B.n690 B.n689 585
R1579 B.n691 B.n476 585
R1580 B.n693 B.n692 585
R1581 B.n695 B.n475 585
R1582 B.n698 B.n697 585
R1583 B.n699 B.n474 585
R1584 B.n701 B.n700 585
R1585 B.n703 B.n473 585
R1586 B.n706 B.n705 585
R1587 B.n707 B.n472 585
R1588 B.n709 B.n708 585
R1589 B.n711 B.n471 585
R1590 B.n714 B.n713 585
R1591 B.n715 B.n470 585
R1592 B.n717 B.n716 585
R1593 B.n719 B.n469 585
R1594 B.n722 B.n721 585
R1595 B.n723 B.n468 585
R1596 B.n725 B.n724 585
R1597 B.n727 B.n467 585
R1598 B.n730 B.n729 585
R1599 B.n731 B.n466 585
R1600 B.n733 B.n732 585
R1601 B.n735 B.n465 585
R1602 B.n738 B.n737 585
R1603 B.n739 B.n464 585
R1604 B.n741 B.n740 585
R1605 B.n743 B.n463 585
R1606 B.n746 B.n745 585
R1607 B.n747 B.n462 585
R1608 B.n749 B.n748 585
R1609 B.n751 B.n461 585
R1610 B.n754 B.n753 585
R1611 B.n755 B.n460 585
R1612 B.n757 B.n756 585
R1613 B.n759 B.n459 585
R1614 B.n762 B.n761 585
R1615 B.n763 B.n458 585
R1616 B.n765 B.n764 585
R1617 B.n767 B.n457 585
R1618 B.n768 B.n456 585
R1619 B.n771 B.n770 585
R1620 B.n772 B.n455 585
R1621 B.n455 B.n454 585
R1622 B.n777 B.n776 585
R1623 B.n776 B.n775 585
R1624 B.n778 B.n451 585
R1625 B.n451 B.n450 585
R1626 B.n780 B.n779 585
R1627 B.n781 B.n780 585
R1628 B.n445 B.n444 585
R1629 B.n446 B.n445 585
R1630 B.n789 B.n788 585
R1631 B.n788 B.n787 585
R1632 B.n790 B.n443 585
R1633 B.n443 B.n441 585
R1634 B.n792 B.n791 585
R1635 B.n793 B.n792 585
R1636 B.n437 B.n436 585
R1637 B.n442 B.n437 585
R1638 B.n801 B.n800 585
R1639 B.n800 B.n799 585
R1640 B.n802 B.n435 585
R1641 B.n435 B.n434 585
R1642 B.n804 B.n803 585
R1643 B.n805 B.n804 585
R1644 B.n429 B.n428 585
R1645 B.n430 B.n429 585
R1646 B.n813 B.n812 585
R1647 B.n812 B.n811 585
R1648 B.n814 B.n427 585
R1649 B.n427 B.n426 585
R1650 B.n816 B.n815 585
R1651 B.n817 B.n816 585
R1652 B.n421 B.n420 585
R1653 B.n422 B.n421 585
R1654 B.n825 B.n824 585
R1655 B.n824 B.n823 585
R1656 B.n826 B.n419 585
R1657 B.n419 B.n418 585
R1658 B.n828 B.n827 585
R1659 B.n829 B.n828 585
R1660 B.n413 B.n412 585
R1661 B.n414 B.n413 585
R1662 B.n837 B.n836 585
R1663 B.n836 B.n835 585
R1664 B.n838 B.n411 585
R1665 B.n411 B.n410 585
R1666 B.n840 B.n839 585
R1667 B.n841 B.n840 585
R1668 B.n405 B.n404 585
R1669 B.n406 B.n405 585
R1670 B.n849 B.n848 585
R1671 B.n848 B.n847 585
R1672 B.n850 B.n403 585
R1673 B.n403 B.n402 585
R1674 B.n852 B.n851 585
R1675 B.n853 B.n852 585
R1676 B.n397 B.n396 585
R1677 B.n398 B.n397 585
R1678 B.n862 B.n861 585
R1679 B.n861 B.n860 585
R1680 B.n863 B.n395 585
R1681 B.n859 B.n395 585
R1682 B.n865 B.n864 585
R1683 B.n866 B.n865 585
R1684 B.n390 B.n389 585
R1685 B.n391 B.n390 585
R1686 B.n875 B.n874 585
R1687 B.n874 B.n873 585
R1688 B.n876 B.n388 585
R1689 B.n388 B.n387 585
R1690 B.n878 B.n877 585
R1691 B.n879 B.n878 585
R1692 B.n2 B.n0 585
R1693 B.n4 B.n2 585
R1694 B.n3 B.n1 585
R1695 B.n1004 B.n3 585
R1696 B.n1002 B.n1001 585
R1697 B.n1003 B.n1002 585
R1698 B.n1000 B.n9 585
R1699 B.n9 B.n8 585
R1700 B.n999 B.n998 585
R1701 B.n998 B.n997 585
R1702 B.n11 B.n10 585
R1703 B.n996 B.n11 585
R1704 B.n994 B.n993 585
R1705 B.n995 B.n994 585
R1706 B.n992 B.n15 585
R1707 B.n18 B.n15 585
R1708 B.n991 B.n990 585
R1709 B.n990 B.n989 585
R1710 B.n17 B.n16 585
R1711 B.n988 B.n17 585
R1712 B.n986 B.n985 585
R1713 B.n987 B.n986 585
R1714 B.n984 B.n23 585
R1715 B.n23 B.n22 585
R1716 B.n983 B.n982 585
R1717 B.n982 B.n981 585
R1718 B.n25 B.n24 585
R1719 B.n980 B.n25 585
R1720 B.n978 B.n977 585
R1721 B.n979 B.n978 585
R1722 B.n976 B.n30 585
R1723 B.n30 B.n29 585
R1724 B.n975 B.n974 585
R1725 B.n974 B.n973 585
R1726 B.n32 B.n31 585
R1727 B.n972 B.n32 585
R1728 B.n970 B.n969 585
R1729 B.n971 B.n970 585
R1730 B.n968 B.n37 585
R1731 B.n37 B.n36 585
R1732 B.n967 B.n966 585
R1733 B.n966 B.n965 585
R1734 B.n39 B.n38 585
R1735 B.n964 B.n39 585
R1736 B.n962 B.n961 585
R1737 B.n963 B.n962 585
R1738 B.n960 B.n44 585
R1739 B.n44 B.n43 585
R1740 B.n959 B.n958 585
R1741 B.n958 B.n957 585
R1742 B.n46 B.n45 585
R1743 B.n956 B.n46 585
R1744 B.n954 B.n953 585
R1745 B.n955 B.n954 585
R1746 B.n952 B.n51 585
R1747 B.n51 B.n50 585
R1748 B.n951 B.n950 585
R1749 B.n950 B.n949 585
R1750 B.n53 B.n52 585
R1751 B.n948 B.n53 585
R1752 B.n946 B.n945 585
R1753 B.n947 B.n946 585
R1754 B.n944 B.n58 585
R1755 B.n58 B.n57 585
R1756 B.n943 B.n942 585
R1757 B.n942 B.n941 585
R1758 B.n60 B.n59 585
R1759 B.n940 B.n60 585
R1760 B.n938 B.n937 585
R1761 B.n939 B.n938 585
R1762 B.n936 B.n65 585
R1763 B.n65 B.n64 585
R1764 B.n935 B.n934 585
R1765 B.n934 B.n933 585
R1766 B.n1007 B.n1006 585
R1767 B.n1006 B.n1005 585
R1768 B.n776 B.n453 497.305
R1769 B.n934 B.n67 497.305
R1770 B.n774 B.n455 497.305
R1771 B.n930 B.n68 497.305
R1772 B.n485 B.t14 440.483
R1773 B.n132 B.t16 440.483
R1774 B.n632 B.t7 440.483
R1775 B.n135 B.t10 440.483
R1776 B.n486 B.t13 379.005
R1777 B.n133 B.t17 379.005
R1778 B.n633 B.t6 379.005
R1779 B.n136 B.t11 379.005
R1780 B.n485 B.t12 357.82
R1781 B.n632 B.t4 357.82
R1782 B.n135 B.t8 357.82
R1783 B.n132 B.t15 357.82
R1784 B.n932 B.n931 256.663
R1785 B.n932 B.n130 256.663
R1786 B.n932 B.n129 256.663
R1787 B.n932 B.n128 256.663
R1788 B.n932 B.n127 256.663
R1789 B.n932 B.n126 256.663
R1790 B.n932 B.n125 256.663
R1791 B.n932 B.n124 256.663
R1792 B.n932 B.n123 256.663
R1793 B.n932 B.n122 256.663
R1794 B.n932 B.n121 256.663
R1795 B.n932 B.n120 256.663
R1796 B.n932 B.n119 256.663
R1797 B.n932 B.n118 256.663
R1798 B.n932 B.n117 256.663
R1799 B.n932 B.n116 256.663
R1800 B.n932 B.n115 256.663
R1801 B.n932 B.n114 256.663
R1802 B.n932 B.n113 256.663
R1803 B.n932 B.n112 256.663
R1804 B.n932 B.n111 256.663
R1805 B.n932 B.n110 256.663
R1806 B.n932 B.n109 256.663
R1807 B.n932 B.n108 256.663
R1808 B.n932 B.n107 256.663
R1809 B.n932 B.n106 256.663
R1810 B.n932 B.n105 256.663
R1811 B.n932 B.n104 256.663
R1812 B.n932 B.n103 256.663
R1813 B.n932 B.n102 256.663
R1814 B.n932 B.n101 256.663
R1815 B.n932 B.n100 256.663
R1816 B.n932 B.n99 256.663
R1817 B.n932 B.n98 256.663
R1818 B.n932 B.n97 256.663
R1819 B.n932 B.n96 256.663
R1820 B.n932 B.n95 256.663
R1821 B.n932 B.n94 256.663
R1822 B.n932 B.n93 256.663
R1823 B.n932 B.n92 256.663
R1824 B.n932 B.n91 256.663
R1825 B.n932 B.n90 256.663
R1826 B.n932 B.n89 256.663
R1827 B.n932 B.n88 256.663
R1828 B.n932 B.n87 256.663
R1829 B.n932 B.n86 256.663
R1830 B.n932 B.n85 256.663
R1831 B.n932 B.n84 256.663
R1832 B.n932 B.n83 256.663
R1833 B.n932 B.n82 256.663
R1834 B.n932 B.n81 256.663
R1835 B.n932 B.n80 256.663
R1836 B.n932 B.n79 256.663
R1837 B.n932 B.n78 256.663
R1838 B.n932 B.n77 256.663
R1839 B.n932 B.n76 256.663
R1840 B.n932 B.n75 256.663
R1841 B.n932 B.n74 256.663
R1842 B.n932 B.n73 256.663
R1843 B.n932 B.n72 256.663
R1844 B.n932 B.n71 256.663
R1845 B.n932 B.n70 256.663
R1846 B.n932 B.n69 256.663
R1847 B.n521 B.n454 256.663
R1848 B.n524 B.n454 256.663
R1849 B.n530 B.n454 256.663
R1850 B.n532 B.n454 256.663
R1851 B.n538 B.n454 256.663
R1852 B.n540 B.n454 256.663
R1853 B.n546 B.n454 256.663
R1854 B.n548 B.n454 256.663
R1855 B.n554 B.n454 256.663
R1856 B.n556 B.n454 256.663
R1857 B.n562 B.n454 256.663
R1858 B.n564 B.n454 256.663
R1859 B.n570 B.n454 256.663
R1860 B.n572 B.n454 256.663
R1861 B.n578 B.n454 256.663
R1862 B.n580 B.n454 256.663
R1863 B.n586 B.n454 256.663
R1864 B.n588 B.n454 256.663
R1865 B.n594 B.n454 256.663
R1866 B.n596 B.n454 256.663
R1867 B.n602 B.n454 256.663
R1868 B.n604 B.n454 256.663
R1869 B.n610 B.n454 256.663
R1870 B.n612 B.n454 256.663
R1871 B.n618 B.n454 256.663
R1872 B.n620 B.n454 256.663
R1873 B.n626 B.n454 256.663
R1874 B.n628 B.n454 256.663
R1875 B.n637 B.n454 256.663
R1876 B.n639 B.n454 256.663
R1877 B.n645 B.n454 256.663
R1878 B.n647 B.n454 256.663
R1879 B.n653 B.n454 256.663
R1880 B.n655 B.n454 256.663
R1881 B.n662 B.n454 256.663
R1882 B.n664 B.n454 256.663
R1883 B.n670 B.n454 256.663
R1884 B.n672 B.n454 256.663
R1885 B.n678 B.n454 256.663
R1886 B.n680 B.n454 256.663
R1887 B.n686 B.n454 256.663
R1888 B.n688 B.n454 256.663
R1889 B.n694 B.n454 256.663
R1890 B.n696 B.n454 256.663
R1891 B.n702 B.n454 256.663
R1892 B.n704 B.n454 256.663
R1893 B.n710 B.n454 256.663
R1894 B.n712 B.n454 256.663
R1895 B.n718 B.n454 256.663
R1896 B.n720 B.n454 256.663
R1897 B.n726 B.n454 256.663
R1898 B.n728 B.n454 256.663
R1899 B.n734 B.n454 256.663
R1900 B.n736 B.n454 256.663
R1901 B.n742 B.n454 256.663
R1902 B.n744 B.n454 256.663
R1903 B.n750 B.n454 256.663
R1904 B.n752 B.n454 256.663
R1905 B.n758 B.n454 256.663
R1906 B.n760 B.n454 256.663
R1907 B.n766 B.n454 256.663
R1908 B.n769 B.n454 256.663
R1909 B.n776 B.n451 163.367
R1910 B.n780 B.n451 163.367
R1911 B.n780 B.n445 163.367
R1912 B.n788 B.n445 163.367
R1913 B.n788 B.n443 163.367
R1914 B.n792 B.n443 163.367
R1915 B.n792 B.n437 163.367
R1916 B.n800 B.n437 163.367
R1917 B.n800 B.n435 163.367
R1918 B.n804 B.n435 163.367
R1919 B.n804 B.n429 163.367
R1920 B.n812 B.n429 163.367
R1921 B.n812 B.n427 163.367
R1922 B.n816 B.n427 163.367
R1923 B.n816 B.n421 163.367
R1924 B.n824 B.n421 163.367
R1925 B.n824 B.n419 163.367
R1926 B.n828 B.n419 163.367
R1927 B.n828 B.n413 163.367
R1928 B.n836 B.n413 163.367
R1929 B.n836 B.n411 163.367
R1930 B.n840 B.n411 163.367
R1931 B.n840 B.n405 163.367
R1932 B.n848 B.n405 163.367
R1933 B.n848 B.n403 163.367
R1934 B.n852 B.n403 163.367
R1935 B.n852 B.n397 163.367
R1936 B.n861 B.n397 163.367
R1937 B.n861 B.n395 163.367
R1938 B.n865 B.n395 163.367
R1939 B.n865 B.n390 163.367
R1940 B.n874 B.n390 163.367
R1941 B.n874 B.n388 163.367
R1942 B.n878 B.n388 163.367
R1943 B.n878 B.n2 163.367
R1944 B.n1006 B.n2 163.367
R1945 B.n1006 B.n3 163.367
R1946 B.n1002 B.n3 163.367
R1947 B.n1002 B.n9 163.367
R1948 B.n998 B.n9 163.367
R1949 B.n998 B.n11 163.367
R1950 B.n994 B.n11 163.367
R1951 B.n994 B.n15 163.367
R1952 B.n990 B.n15 163.367
R1953 B.n990 B.n17 163.367
R1954 B.n986 B.n17 163.367
R1955 B.n986 B.n23 163.367
R1956 B.n982 B.n23 163.367
R1957 B.n982 B.n25 163.367
R1958 B.n978 B.n25 163.367
R1959 B.n978 B.n30 163.367
R1960 B.n974 B.n30 163.367
R1961 B.n974 B.n32 163.367
R1962 B.n970 B.n32 163.367
R1963 B.n970 B.n37 163.367
R1964 B.n966 B.n37 163.367
R1965 B.n966 B.n39 163.367
R1966 B.n962 B.n39 163.367
R1967 B.n962 B.n44 163.367
R1968 B.n958 B.n44 163.367
R1969 B.n958 B.n46 163.367
R1970 B.n954 B.n46 163.367
R1971 B.n954 B.n51 163.367
R1972 B.n950 B.n51 163.367
R1973 B.n950 B.n53 163.367
R1974 B.n946 B.n53 163.367
R1975 B.n946 B.n58 163.367
R1976 B.n942 B.n58 163.367
R1977 B.n942 B.n60 163.367
R1978 B.n938 B.n60 163.367
R1979 B.n938 B.n65 163.367
R1980 B.n934 B.n65 163.367
R1981 B.n523 B.n522 163.367
R1982 B.n525 B.n523 163.367
R1983 B.n529 B.n518 163.367
R1984 B.n533 B.n531 163.367
R1985 B.n537 B.n516 163.367
R1986 B.n541 B.n539 163.367
R1987 B.n545 B.n514 163.367
R1988 B.n549 B.n547 163.367
R1989 B.n553 B.n512 163.367
R1990 B.n557 B.n555 163.367
R1991 B.n561 B.n510 163.367
R1992 B.n565 B.n563 163.367
R1993 B.n569 B.n508 163.367
R1994 B.n573 B.n571 163.367
R1995 B.n577 B.n506 163.367
R1996 B.n581 B.n579 163.367
R1997 B.n585 B.n504 163.367
R1998 B.n589 B.n587 163.367
R1999 B.n593 B.n502 163.367
R2000 B.n597 B.n595 163.367
R2001 B.n601 B.n500 163.367
R2002 B.n605 B.n603 163.367
R2003 B.n609 B.n498 163.367
R2004 B.n613 B.n611 163.367
R2005 B.n617 B.n496 163.367
R2006 B.n621 B.n619 163.367
R2007 B.n625 B.n494 163.367
R2008 B.n629 B.n627 163.367
R2009 B.n636 B.n492 163.367
R2010 B.n640 B.n638 163.367
R2011 B.n644 B.n490 163.367
R2012 B.n648 B.n646 163.367
R2013 B.n652 B.n488 163.367
R2014 B.n656 B.n654 163.367
R2015 B.n661 B.n484 163.367
R2016 B.n665 B.n663 163.367
R2017 B.n669 B.n482 163.367
R2018 B.n673 B.n671 163.367
R2019 B.n677 B.n480 163.367
R2020 B.n681 B.n679 163.367
R2021 B.n685 B.n478 163.367
R2022 B.n689 B.n687 163.367
R2023 B.n693 B.n476 163.367
R2024 B.n697 B.n695 163.367
R2025 B.n701 B.n474 163.367
R2026 B.n705 B.n703 163.367
R2027 B.n709 B.n472 163.367
R2028 B.n713 B.n711 163.367
R2029 B.n717 B.n470 163.367
R2030 B.n721 B.n719 163.367
R2031 B.n725 B.n468 163.367
R2032 B.n729 B.n727 163.367
R2033 B.n733 B.n466 163.367
R2034 B.n737 B.n735 163.367
R2035 B.n741 B.n464 163.367
R2036 B.n745 B.n743 163.367
R2037 B.n749 B.n462 163.367
R2038 B.n753 B.n751 163.367
R2039 B.n757 B.n460 163.367
R2040 B.n761 B.n759 163.367
R2041 B.n765 B.n458 163.367
R2042 B.n768 B.n767 163.367
R2043 B.n770 B.n455 163.367
R2044 B.n774 B.n449 163.367
R2045 B.n782 B.n449 163.367
R2046 B.n782 B.n447 163.367
R2047 B.n786 B.n447 163.367
R2048 B.n786 B.n440 163.367
R2049 B.n794 B.n440 163.367
R2050 B.n794 B.n438 163.367
R2051 B.n798 B.n438 163.367
R2052 B.n798 B.n433 163.367
R2053 B.n806 B.n433 163.367
R2054 B.n806 B.n431 163.367
R2055 B.n810 B.n431 163.367
R2056 B.n810 B.n425 163.367
R2057 B.n818 B.n425 163.367
R2058 B.n818 B.n423 163.367
R2059 B.n822 B.n423 163.367
R2060 B.n822 B.n417 163.367
R2061 B.n830 B.n417 163.367
R2062 B.n830 B.n415 163.367
R2063 B.n834 B.n415 163.367
R2064 B.n834 B.n409 163.367
R2065 B.n842 B.n409 163.367
R2066 B.n842 B.n407 163.367
R2067 B.n846 B.n407 163.367
R2068 B.n846 B.n401 163.367
R2069 B.n854 B.n401 163.367
R2070 B.n854 B.n399 163.367
R2071 B.n858 B.n399 163.367
R2072 B.n858 B.n394 163.367
R2073 B.n867 B.n394 163.367
R2074 B.n867 B.n392 163.367
R2075 B.n872 B.n392 163.367
R2076 B.n872 B.n386 163.367
R2077 B.n880 B.n386 163.367
R2078 B.n881 B.n880 163.367
R2079 B.n881 B.n5 163.367
R2080 B.n6 B.n5 163.367
R2081 B.n7 B.n6 163.367
R2082 B.n886 B.n7 163.367
R2083 B.n886 B.n12 163.367
R2084 B.n13 B.n12 163.367
R2085 B.n14 B.n13 163.367
R2086 B.n891 B.n14 163.367
R2087 B.n891 B.n19 163.367
R2088 B.n20 B.n19 163.367
R2089 B.n21 B.n20 163.367
R2090 B.n896 B.n21 163.367
R2091 B.n896 B.n26 163.367
R2092 B.n27 B.n26 163.367
R2093 B.n28 B.n27 163.367
R2094 B.n901 B.n28 163.367
R2095 B.n901 B.n33 163.367
R2096 B.n34 B.n33 163.367
R2097 B.n35 B.n34 163.367
R2098 B.n906 B.n35 163.367
R2099 B.n906 B.n40 163.367
R2100 B.n41 B.n40 163.367
R2101 B.n42 B.n41 163.367
R2102 B.n911 B.n42 163.367
R2103 B.n911 B.n47 163.367
R2104 B.n48 B.n47 163.367
R2105 B.n49 B.n48 163.367
R2106 B.n916 B.n49 163.367
R2107 B.n916 B.n54 163.367
R2108 B.n55 B.n54 163.367
R2109 B.n56 B.n55 163.367
R2110 B.n921 B.n56 163.367
R2111 B.n921 B.n61 163.367
R2112 B.n62 B.n61 163.367
R2113 B.n63 B.n62 163.367
R2114 B.n926 B.n63 163.367
R2115 B.n926 B.n68 163.367
R2116 B.n140 B.n139 163.367
R2117 B.n144 B.n143 163.367
R2118 B.n148 B.n147 163.367
R2119 B.n152 B.n151 163.367
R2120 B.n156 B.n155 163.367
R2121 B.n160 B.n159 163.367
R2122 B.n164 B.n163 163.367
R2123 B.n168 B.n167 163.367
R2124 B.n172 B.n171 163.367
R2125 B.n176 B.n175 163.367
R2126 B.n180 B.n179 163.367
R2127 B.n184 B.n183 163.367
R2128 B.n188 B.n187 163.367
R2129 B.n192 B.n191 163.367
R2130 B.n196 B.n195 163.367
R2131 B.n200 B.n199 163.367
R2132 B.n204 B.n203 163.367
R2133 B.n208 B.n207 163.367
R2134 B.n212 B.n211 163.367
R2135 B.n216 B.n215 163.367
R2136 B.n220 B.n219 163.367
R2137 B.n224 B.n223 163.367
R2138 B.n228 B.n227 163.367
R2139 B.n232 B.n231 163.367
R2140 B.n236 B.n235 163.367
R2141 B.n240 B.n239 163.367
R2142 B.n244 B.n243 163.367
R2143 B.n248 B.n247 163.367
R2144 B.n252 B.n251 163.367
R2145 B.n256 B.n255 163.367
R2146 B.n260 B.n259 163.367
R2147 B.n264 B.n263 163.367
R2148 B.n268 B.n267 163.367
R2149 B.n272 B.n271 163.367
R2150 B.n276 B.n275 163.367
R2151 B.n280 B.n279 163.367
R2152 B.n284 B.n283 163.367
R2153 B.n288 B.n287 163.367
R2154 B.n292 B.n291 163.367
R2155 B.n296 B.n295 163.367
R2156 B.n300 B.n299 163.367
R2157 B.n304 B.n303 163.367
R2158 B.n308 B.n307 163.367
R2159 B.n312 B.n311 163.367
R2160 B.n316 B.n315 163.367
R2161 B.n320 B.n319 163.367
R2162 B.n324 B.n323 163.367
R2163 B.n328 B.n327 163.367
R2164 B.n332 B.n331 163.367
R2165 B.n336 B.n335 163.367
R2166 B.n340 B.n339 163.367
R2167 B.n344 B.n343 163.367
R2168 B.n348 B.n347 163.367
R2169 B.n352 B.n351 163.367
R2170 B.n356 B.n355 163.367
R2171 B.n360 B.n359 163.367
R2172 B.n364 B.n363 163.367
R2173 B.n368 B.n367 163.367
R2174 B.n372 B.n371 163.367
R2175 B.n376 B.n375 163.367
R2176 B.n380 B.n379 163.367
R2177 B.n382 B.n131 163.367
R2178 B.n521 B.n453 71.676
R2179 B.n525 B.n524 71.676
R2180 B.n530 B.n529 71.676
R2181 B.n533 B.n532 71.676
R2182 B.n538 B.n537 71.676
R2183 B.n541 B.n540 71.676
R2184 B.n546 B.n545 71.676
R2185 B.n549 B.n548 71.676
R2186 B.n554 B.n553 71.676
R2187 B.n557 B.n556 71.676
R2188 B.n562 B.n561 71.676
R2189 B.n565 B.n564 71.676
R2190 B.n570 B.n569 71.676
R2191 B.n573 B.n572 71.676
R2192 B.n578 B.n577 71.676
R2193 B.n581 B.n580 71.676
R2194 B.n586 B.n585 71.676
R2195 B.n589 B.n588 71.676
R2196 B.n594 B.n593 71.676
R2197 B.n597 B.n596 71.676
R2198 B.n602 B.n601 71.676
R2199 B.n605 B.n604 71.676
R2200 B.n610 B.n609 71.676
R2201 B.n613 B.n612 71.676
R2202 B.n618 B.n617 71.676
R2203 B.n621 B.n620 71.676
R2204 B.n626 B.n625 71.676
R2205 B.n629 B.n628 71.676
R2206 B.n637 B.n636 71.676
R2207 B.n640 B.n639 71.676
R2208 B.n645 B.n644 71.676
R2209 B.n648 B.n647 71.676
R2210 B.n653 B.n652 71.676
R2211 B.n656 B.n655 71.676
R2212 B.n662 B.n661 71.676
R2213 B.n665 B.n664 71.676
R2214 B.n670 B.n669 71.676
R2215 B.n673 B.n672 71.676
R2216 B.n678 B.n677 71.676
R2217 B.n681 B.n680 71.676
R2218 B.n686 B.n685 71.676
R2219 B.n689 B.n688 71.676
R2220 B.n694 B.n693 71.676
R2221 B.n697 B.n696 71.676
R2222 B.n702 B.n701 71.676
R2223 B.n705 B.n704 71.676
R2224 B.n710 B.n709 71.676
R2225 B.n713 B.n712 71.676
R2226 B.n718 B.n717 71.676
R2227 B.n721 B.n720 71.676
R2228 B.n726 B.n725 71.676
R2229 B.n729 B.n728 71.676
R2230 B.n734 B.n733 71.676
R2231 B.n737 B.n736 71.676
R2232 B.n742 B.n741 71.676
R2233 B.n745 B.n744 71.676
R2234 B.n750 B.n749 71.676
R2235 B.n753 B.n752 71.676
R2236 B.n758 B.n757 71.676
R2237 B.n761 B.n760 71.676
R2238 B.n766 B.n765 71.676
R2239 B.n769 B.n768 71.676
R2240 B.n69 B.n67 71.676
R2241 B.n140 B.n70 71.676
R2242 B.n144 B.n71 71.676
R2243 B.n148 B.n72 71.676
R2244 B.n152 B.n73 71.676
R2245 B.n156 B.n74 71.676
R2246 B.n160 B.n75 71.676
R2247 B.n164 B.n76 71.676
R2248 B.n168 B.n77 71.676
R2249 B.n172 B.n78 71.676
R2250 B.n176 B.n79 71.676
R2251 B.n180 B.n80 71.676
R2252 B.n184 B.n81 71.676
R2253 B.n188 B.n82 71.676
R2254 B.n192 B.n83 71.676
R2255 B.n196 B.n84 71.676
R2256 B.n200 B.n85 71.676
R2257 B.n204 B.n86 71.676
R2258 B.n208 B.n87 71.676
R2259 B.n212 B.n88 71.676
R2260 B.n216 B.n89 71.676
R2261 B.n220 B.n90 71.676
R2262 B.n224 B.n91 71.676
R2263 B.n228 B.n92 71.676
R2264 B.n232 B.n93 71.676
R2265 B.n236 B.n94 71.676
R2266 B.n240 B.n95 71.676
R2267 B.n244 B.n96 71.676
R2268 B.n248 B.n97 71.676
R2269 B.n252 B.n98 71.676
R2270 B.n256 B.n99 71.676
R2271 B.n260 B.n100 71.676
R2272 B.n264 B.n101 71.676
R2273 B.n268 B.n102 71.676
R2274 B.n272 B.n103 71.676
R2275 B.n276 B.n104 71.676
R2276 B.n280 B.n105 71.676
R2277 B.n284 B.n106 71.676
R2278 B.n288 B.n107 71.676
R2279 B.n292 B.n108 71.676
R2280 B.n296 B.n109 71.676
R2281 B.n300 B.n110 71.676
R2282 B.n304 B.n111 71.676
R2283 B.n308 B.n112 71.676
R2284 B.n312 B.n113 71.676
R2285 B.n316 B.n114 71.676
R2286 B.n320 B.n115 71.676
R2287 B.n324 B.n116 71.676
R2288 B.n328 B.n117 71.676
R2289 B.n332 B.n118 71.676
R2290 B.n336 B.n119 71.676
R2291 B.n340 B.n120 71.676
R2292 B.n344 B.n121 71.676
R2293 B.n348 B.n122 71.676
R2294 B.n352 B.n123 71.676
R2295 B.n356 B.n124 71.676
R2296 B.n360 B.n125 71.676
R2297 B.n364 B.n126 71.676
R2298 B.n368 B.n127 71.676
R2299 B.n372 B.n128 71.676
R2300 B.n376 B.n129 71.676
R2301 B.n380 B.n130 71.676
R2302 B.n931 B.n131 71.676
R2303 B.n931 B.n930 71.676
R2304 B.n382 B.n130 71.676
R2305 B.n379 B.n129 71.676
R2306 B.n375 B.n128 71.676
R2307 B.n371 B.n127 71.676
R2308 B.n367 B.n126 71.676
R2309 B.n363 B.n125 71.676
R2310 B.n359 B.n124 71.676
R2311 B.n355 B.n123 71.676
R2312 B.n351 B.n122 71.676
R2313 B.n347 B.n121 71.676
R2314 B.n343 B.n120 71.676
R2315 B.n339 B.n119 71.676
R2316 B.n335 B.n118 71.676
R2317 B.n331 B.n117 71.676
R2318 B.n327 B.n116 71.676
R2319 B.n323 B.n115 71.676
R2320 B.n319 B.n114 71.676
R2321 B.n315 B.n113 71.676
R2322 B.n311 B.n112 71.676
R2323 B.n307 B.n111 71.676
R2324 B.n303 B.n110 71.676
R2325 B.n299 B.n109 71.676
R2326 B.n295 B.n108 71.676
R2327 B.n291 B.n107 71.676
R2328 B.n287 B.n106 71.676
R2329 B.n283 B.n105 71.676
R2330 B.n279 B.n104 71.676
R2331 B.n275 B.n103 71.676
R2332 B.n271 B.n102 71.676
R2333 B.n267 B.n101 71.676
R2334 B.n263 B.n100 71.676
R2335 B.n259 B.n99 71.676
R2336 B.n255 B.n98 71.676
R2337 B.n251 B.n97 71.676
R2338 B.n247 B.n96 71.676
R2339 B.n243 B.n95 71.676
R2340 B.n239 B.n94 71.676
R2341 B.n235 B.n93 71.676
R2342 B.n231 B.n92 71.676
R2343 B.n227 B.n91 71.676
R2344 B.n223 B.n90 71.676
R2345 B.n219 B.n89 71.676
R2346 B.n215 B.n88 71.676
R2347 B.n211 B.n87 71.676
R2348 B.n207 B.n86 71.676
R2349 B.n203 B.n85 71.676
R2350 B.n199 B.n84 71.676
R2351 B.n195 B.n83 71.676
R2352 B.n191 B.n82 71.676
R2353 B.n187 B.n81 71.676
R2354 B.n183 B.n80 71.676
R2355 B.n179 B.n79 71.676
R2356 B.n175 B.n78 71.676
R2357 B.n171 B.n77 71.676
R2358 B.n167 B.n76 71.676
R2359 B.n163 B.n75 71.676
R2360 B.n159 B.n74 71.676
R2361 B.n155 B.n73 71.676
R2362 B.n151 B.n72 71.676
R2363 B.n147 B.n71 71.676
R2364 B.n143 B.n70 71.676
R2365 B.n139 B.n69 71.676
R2366 B.n522 B.n521 71.676
R2367 B.n524 B.n518 71.676
R2368 B.n531 B.n530 71.676
R2369 B.n532 B.n516 71.676
R2370 B.n539 B.n538 71.676
R2371 B.n540 B.n514 71.676
R2372 B.n547 B.n546 71.676
R2373 B.n548 B.n512 71.676
R2374 B.n555 B.n554 71.676
R2375 B.n556 B.n510 71.676
R2376 B.n563 B.n562 71.676
R2377 B.n564 B.n508 71.676
R2378 B.n571 B.n570 71.676
R2379 B.n572 B.n506 71.676
R2380 B.n579 B.n578 71.676
R2381 B.n580 B.n504 71.676
R2382 B.n587 B.n586 71.676
R2383 B.n588 B.n502 71.676
R2384 B.n595 B.n594 71.676
R2385 B.n596 B.n500 71.676
R2386 B.n603 B.n602 71.676
R2387 B.n604 B.n498 71.676
R2388 B.n611 B.n610 71.676
R2389 B.n612 B.n496 71.676
R2390 B.n619 B.n618 71.676
R2391 B.n620 B.n494 71.676
R2392 B.n627 B.n626 71.676
R2393 B.n628 B.n492 71.676
R2394 B.n638 B.n637 71.676
R2395 B.n639 B.n490 71.676
R2396 B.n646 B.n645 71.676
R2397 B.n647 B.n488 71.676
R2398 B.n654 B.n653 71.676
R2399 B.n655 B.n484 71.676
R2400 B.n663 B.n662 71.676
R2401 B.n664 B.n482 71.676
R2402 B.n671 B.n670 71.676
R2403 B.n672 B.n480 71.676
R2404 B.n679 B.n678 71.676
R2405 B.n680 B.n478 71.676
R2406 B.n687 B.n686 71.676
R2407 B.n688 B.n476 71.676
R2408 B.n695 B.n694 71.676
R2409 B.n696 B.n474 71.676
R2410 B.n703 B.n702 71.676
R2411 B.n704 B.n472 71.676
R2412 B.n711 B.n710 71.676
R2413 B.n712 B.n470 71.676
R2414 B.n719 B.n718 71.676
R2415 B.n720 B.n468 71.676
R2416 B.n727 B.n726 71.676
R2417 B.n728 B.n466 71.676
R2418 B.n735 B.n734 71.676
R2419 B.n736 B.n464 71.676
R2420 B.n743 B.n742 71.676
R2421 B.n744 B.n462 71.676
R2422 B.n751 B.n750 71.676
R2423 B.n752 B.n460 71.676
R2424 B.n759 B.n758 71.676
R2425 B.n760 B.n458 71.676
R2426 B.n767 B.n766 71.676
R2427 B.n770 B.n769 71.676
R2428 B.n775 B.n454 62.0062
R2429 B.n933 B.n932 62.0062
R2430 B.n486 B.n485 61.4793
R2431 B.n633 B.n632 61.4793
R2432 B.n136 B.n135 61.4793
R2433 B.n133 B.n132 61.4793
R2434 B.n658 B.n486 59.5399
R2435 B.n634 B.n633 59.5399
R2436 B.n137 B.n136 59.5399
R2437 B.n134 B.n133 59.5399
R2438 B.n775 B.n450 32.6857
R2439 B.n781 B.n450 32.6857
R2440 B.n781 B.n446 32.6857
R2441 B.n787 B.n446 32.6857
R2442 B.n787 B.n441 32.6857
R2443 B.n793 B.n441 32.6857
R2444 B.n793 B.n442 32.6857
R2445 B.n799 B.n434 32.6857
R2446 B.n805 B.n434 32.6857
R2447 B.n805 B.n430 32.6857
R2448 B.n811 B.n430 32.6857
R2449 B.n811 B.n426 32.6857
R2450 B.n817 B.n426 32.6857
R2451 B.n817 B.n422 32.6857
R2452 B.n823 B.n422 32.6857
R2453 B.n823 B.n418 32.6857
R2454 B.n829 B.n418 32.6857
R2455 B.n829 B.n414 32.6857
R2456 B.n835 B.n414 32.6857
R2457 B.n841 B.n410 32.6857
R2458 B.n841 B.n406 32.6857
R2459 B.n847 B.n406 32.6857
R2460 B.n847 B.n402 32.6857
R2461 B.n853 B.n402 32.6857
R2462 B.n853 B.n398 32.6857
R2463 B.n860 B.n398 32.6857
R2464 B.n860 B.n859 32.6857
R2465 B.n866 B.n391 32.6857
R2466 B.n873 B.n391 32.6857
R2467 B.n873 B.n387 32.6857
R2468 B.n879 B.n387 32.6857
R2469 B.n879 B.n4 32.6857
R2470 B.n1005 B.n4 32.6857
R2471 B.n1005 B.n1004 32.6857
R2472 B.n1004 B.n1003 32.6857
R2473 B.n1003 B.n8 32.6857
R2474 B.n997 B.n8 32.6857
R2475 B.n997 B.n996 32.6857
R2476 B.n996 B.n995 32.6857
R2477 B.n989 B.n18 32.6857
R2478 B.n989 B.n988 32.6857
R2479 B.n988 B.n987 32.6857
R2480 B.n987 B.n22 32.6857
R2481 B.n981 B.n22 32.6857
R2482 B.n981 B.n980 32.6857
R2483 B.n980 B.n979 32.6857
R2484 B.n979 B.n29 32.6857
R2485 B.n973 B.n972 32.6857
R2486 B.n972 B.n971 32.6857
R2487 B.n971 B.n36 32.6857
R2488 B.n965 B.n36 32.6857
R2489 B.n965 B.n964 32.6857
R2490 B.n964 B.n963 32.6857
R2491 B.n963 B.n43 32.6857
R2492 B.n957 B.n43 32.6857
R2493 B.n957 B.n956 32.6857
R2494 B.n956 B.n955 32.6857
R2495 B.n955 B.n50 32.6857
R2496 B.n949 B.n50 32.6857
R2497 B.n948 B.n947 32.6857
R2498 B.n947 B.n57 32.6857
R2499 B.n941 B.n57 32.6857
R2500 B.n941 B.n940 32.6857
R2501 B.n940 B.n939 32.6857
R2502 B.n939 B.n64 32.6857
R2503 B.n933 B.n64 32.6857
R2504 B.n935 B.n66 32.3127
R2505 B.n929 B.n928 32.3127
R2506 B.n773 B.n772 32.3127
R2507 B.n777 B.n452 32.3127
R2508 B.n442 B.t5 28.8404
R2509 B.t9 B.n948 28.8404
R2510 B.n859 B.t3 24.0337
R2511 B.n18 B.t2 24.0337
R2512 B.t0 B.n410 19.2271
R2513 B.t1 B.n29 19.2271
R2514 B B.n1007 18.0485
R2515 B.n835 B.t0 13.4591
R2516 B.n973 B.t1 13.4591
R2517 B.n138 B.n66 10.6151
R2518 B.n141 B.n138 10.6151
R2519 B.n142 B.n141 10.6151
R2520 B.n145 B.n142 10.6151
R2521 B.n146 B.n145 10.6151
R2522 B.n149 B.n146 10.6151
R2523 B.n150 B.n149 10.6151
R2524 B.n153 B.n150 10.6151
R2525 B.n154 B.n153 10.6151
R2526 B.n157 B.n154 10.6151
R2527 B.n158 B.n157 10.6151
R2528 B.n161 B.n158 10.6151
R2529 B.n162 B.n161 10.6151
R2530 B.n165 B.n162 10.6151
R2531 B.n166 B.n165 10.6151
R2532 B.n169 B.n166 10.6151
R2533 B.n170 B.n169 10.6151
R2534 B.n173 B.n170 10.6151
R2535 B.n174 B.n173 10.6151
R2536 B.n177 B.n174 10.6151
R2537 B.n178 B.n177 10.6151
R2538 B.n181 B.n178 10.6151
R2539 B.n182 B.n181 10.6151
R2540 B.n185 B.n182 10.6151
R2541 B.n186 B.n185 10.6151
R2542 B.n189 B.n186 10.6151
R2543 B.n190 B.n189 10.6151
R2544 B.n193 B.n190 10.6151
R2545 B.n194 B.n193 10.6151
R2546 B.n197 B.n194 10.6151
R2547 B.n198 B.n197 10.6151
R2548 B.n201 B.n198 10.6151
R2549 B.n202 B.n201 10.6151
R2550 B.n205 B.n202 10.6151
R2551 B.n206 B.n205 10.6151
R2552 B.n209 B.n206 10.6151
R2553 B.n210 B.n209 10.6151
R2554 B.n213 B.n210 10.6151
R2555 B.n214 B.n213 10.6151
R2556 B.n217 B.n214 10.6151
R2557 B.n218 B.n217 10.6151
R2558 B.n221 B.n218 10.6151
R2559 B.n222 B.n221 10.6151
R2560 B.n225 B.n222 10.6151
R2561 B.n226 B.n225 10.6151
R2562 B.n229 B.n226 10.6151
R2563 B.n230 B.n229 10.6151
R2564 B.n233 B.n230 10.6151
R2565 B.n234 B.n233 10.6151
R2566 B.n237 B.n234 10.6151
R2567 B.n238 B.n237 10.6151
R2568 B.n241 B.n238 10.6151
R2569 B.n242 B.n241 10.6151
R2570 B.n245 B.n242 10.6151
R2571 B.n246 B.n245 10.6151
R2572 B.n249 B.n246 10.6151
R2573 B.n250 B.n249 10.6151
R2574 B.n254 B.n253 10.6151
R2575 B.n257 B.n254 10.6151
R2576 B.n258 B.n257 10.6151
R2577 B.n261 B.n258 10.6151
R2578 B.n262 B.n261 10.6151
R2579 B.n265 B.n262 10.6151
R2580 B.n266 B.n265 10.6151
R2581 B.n269 B.n266 10.6151
R2582 B.n270 B.n269 10.6151
R2583 B.n274 B.n273 10.6151
R2584 B.n277 B.n274 10.6151
R2585 B.n278 B.n277 10.6151
R2586 B.n281 B.n278 10.6151
R2587 B.n282 B.n281 10.6151
R2588 B.n285 B.n282 10.6151
R2589 B.n286 B.n285 10.6151
R2590 B.n289 B.n286 10.6151
R2591 B.n290 B.n289 10.6151
R2592 B.n293 B.n290 10.6151
R2593 B.n294 B.n293 10.6151
R2594 B.n297 B.n294 10.6151
R2595 B.n298 B.n297 10.6151
R2596 B.n301 B.n298 10.6151
R2597 B.n302 B.n301 10.6151
R2598 B.n305 B.n302 10.6151
R2599 B.n306 B.n305 10.6151
R2600 B.n309 B.n306 10.6151
R2601 B.n310 B.n309 10.6151
R2602 B.n313 B.n310 10.6151
R2603 B.n314 B.n313 10.6151
R2604 B.n317 B.n314 10.6151
R2605 B.n318 B.n317 10.6151
R2606 B.n321 B.n318 10.6151
R2607 B.n322 B.n321 10.6151
R2608 B.n325 B.n322 10.6151
R2609 B.n326 B.n325 10.6151
R2610 B.n329 B.n326 10.6151
R2611 B.n330 B.n329 10.6151
R2612 B.n333 B.n330 10.6151
R2613 B.n334 B.n333 10.6151
R2614 B.n337 B.n334 10.6151
R2615 B.n338 B.n337 10.6151
R2616 B.n341 B.n338 10.6151
R2617 B.n342 B.n341 10.6151
R2618 B.n345 B.n342 10.6151
R2619 B.n346 B.n345 10.6151
R2620 B.n349 B.n346 10.6151
R2621 B.n350 B.n349 10.6151
R2622 B.n353 B.n350 10.6151
R2623 B.n354 B.n353 10.6151
R2624 B.n357 B.n354 10.6151
R2625 B.n358 B.n357 10.6151
R2626 B.n361 B.n358 10.6151
R2627 B.n362 B.n361 10.6151
R2628 B.n365 B.n362 10.6151
R2629 B.n366 B.n365 10.6151
R2630 B.n369 B.n366 10.6151
R2631 B.n370 B.n369 10.6151
R2632 B.n373 B.n370 10.6151
R2633 B.n374 B.n373 10.6151
R2634 B.n377 B.n374 10.6151
R2635 B.n378 B.n377 10.6151
R2636 B.n381 B.n378 10.6151
R2637 B.n383 B.n381 10.6151
R2638 B.n384 B.n383 10.6151
R2639 B.n929 B.n384 10.6151
R2640 B.n773 B.n448 10.6151
R2641 B.n783 B.n448 10.6151
R2642 B.n784 B.n783 10.6151
R2643 B.n785 B.n784 10.6151
R2644 B.n785 B.n439 10.6151
R2645 B.n795 B.n439 10.6151
R2646 B.n796 B.n795 10.6151
R2647 B.n797 B.n796 10.6151
R2648 B.n797 B.n432 10.6151
R2649 B.n807 B.n432 10.6151
R2650 B.n808 B.n807 10.6151
R2651 B.n809 B.n808 10.6151
R2652 B.n809 B.n424 10.6151
R2653 B.n819 B.n424 10.6151
R2654 B.n820 B.n819 10.6151
R2655 B.n821 B.n820 10.6151
R2656 B.n821 B.n416 10.6151
R2657 B.n831 B.n416 10.6151
R2658 B.n832 B.n831 10.6151
R2659 B.n833 B.n832 10.6151
R2660 B.n833 B.n408 10.6151
R2661 B.n843 B.n408 10.6151
R2662 B.n844 B.n843 10.6151
R2663 B.n845 B.n844 10.6151
R2664 B.n845 B.n400 10.6151
R2665 B.n855 B.n400 10.6151
R2666 B.n856 B.n855 10.6151
R2667 B.n857 B.n856 10.6151
R2668 B.n857 B.n393 10.6151
R2669 B.n868 B.n393 10.6151
R2670 B.n869 B.n868 10.6151
R2671 B.n871 B.n869 10.6151
R2672 B.n871 B.n870 10.6151
R2673 B.n870 B.n385 10.6151
R2674 B.n882 B.n385 10.6151
R2675 B.n883 B.n882 10.6151
R2676 B.n884 B.n883 10.6151
R2677 B.n885 B.n884 10.6151
R2678 B.n887 B.n885 10.6151
R2679 B.n888 B.n887 10.6151
R2680 B.n889 B.n888 10.6151
R2681 B.n890 B.n889 10.6151
R2682 B.n892 B.n890 10.6151
R2683 B.n893 B.n892 10.6151
R2684 B.n894 B.n893 10.6151
R2685 B.n895 B.n894 10.6151
R2686 B.n897 B.n895 10.6151
R2687 B.n898 B.n897 10.6151
R2688 B.n899 B.n898 10.6151
R2689 B.n900 B.n899 10.6151
R2690 B.n902 B.n900 10.6151
R2691 B.n903 B.n902 10.6151
R2692 B.n904 B.n903 10.6151
R2693 B.n905 B.n904 10.6151
R2694 B.n907 B.n905 10.6151
R2695 B.n908 B.n907 10.6151
R2696 B.n909 B.n908 10.6151
R2697 B.n910 B.n909 10.6151
R2698 B.n912 B.n910 10.6151
R2699 B.n913 B.n912 10.6151
R2700 B.n914 B.n913 10.6151
R2701 B.n915 B.n914 10.6151
R2702 B.n917 B.n915 10.6151
R2703 B.n918 B.n917 10.6151
R2704 B.n919 B.n918 10.6151
R2705 B.n920 B.n919 10.6151
R2706 B.n922 B.n920 10.6151
R2707 B.n923 B.n922 10.6151
R2708 B.n924 B.n923 10.6151
R2709 B.n925 B.n924 10.6151
R2710 B.n927 B.n925 10.6151
R2711 B.n928 B.n927 10.6151
R2712 B.n520 B.n452 10.6151
R2713 B.n520 B.n519 10.6151
R2714 B.n526 B.n519 10.6151
R2715 B.n527 B.n526 10.6151
R2716 B.n528 B.n527 10.6151
R2717 B.n528 B.n517 10.6151
R2718 B.n534 B.n517 10.6151
R2719 B.n535 B.n534 10.6151
R2720 B.n536 B.n535 10.6151
R2721 B.n536 B.n515 10.6151
R2722 B.n542 B.n515 10.6151
R2723 B.n543 B.n542 10.6151
R2724 B.n544 B.n543 10.6151
R2725 B.n544 B.n513 10.6151
R2726 B.n550 B.n513 10.6151
R2727 B.n551 B.n550 10.6151
R2728 B.n552 B.n551 10.6151
R2729 B.n552 B.n511 10.6151
R2730 B.n558 B.n511 10.6151
R2731 B.n559 B.n558 10.6151
R2732 B.n560 B.n559 10.6151
R2733 B.n560 B.n509 10.6151
R2734 B.n566 B.n509 10.6151
R2735 B.n567 B.n566 10.6151
R2736 B.n568 B.n567 10.6151
R2737 B.n568 B.n507 10.6151
R2738 B.n574 B.n507 10.6151
R2739 B.n575 B.n574 10.6151
R2740 B.n576 B.n575 10.6151
R2741 B.n576 B.n505 10.6151
R2742 B.n582 B.n505 10.6151
R2743 B.n583 B.n582 10.6151
R2744 B.n584 B.n583 10.6151
R2745 B.n584 B.n503 10.6151
R2746 B.n590 B.n503 10.6151
R2747 B.n591 B.n590 10.6151
R2748 B.n592 B.n591 10.6151
R2749 B.n592 B.n501 10.6151
R2750 B.n598 B.n501 10.6151
R2751 B.n599 B.n598 10.6151
R2752 B.n600 B.n599 10.6151
R2753 B.n600 B.n499 10.6151
R2754 B.n606 B.n499 10.6151
R2755 B.n607 B.n606 10.6151
R2756 B.n608 B.n607 10.6151
R2757 B.n608 B.n497 10.6151
R2758 B.n614 B.n497 10.6151
R2759 B.n615 B.n614 10.6151
R2760 B.n616 B.n615 10.6151
R2761 B.n616 B.n495 10.6151
R2762 B.n622 B.n495 10.6151
R2763 B.n623 B.n622 10.6151
R2764 B.n624 B.n623 10.6151
R2765 B.n624 B.n493 10.6151
R2766 B.n630 B.n493 10.6151
R2767 B.n631 B.n630 10.6151
R2768 B.n635 B.n631 10.6151
R2769 B.n641 B.n491 10.6151
R2770 B.n642 B.n641 10.6151
R2771 B.n643 B.n642 10.6151
R2772 B.n643 B.n489 10.6151
R2773 B.n649 B.n489 10.6151
R2774 B.n650 B.n649 10.6151
R2775 B.n651 B.n650 10.6151
R2776 B.n651 B.n487 10.6151
R2777 B.n657 B.n487 10.6151
R2778 B.n660 B.n659 10.6151
R2779 B.n660 B.n483 10.6151
R2780 B.n666 B.n483 10.6151
R2781 B.n667 B.n666 10.6151
R2782 B.n668 B.n667 10.6151
R2783 B.n668 B.n481 10.6151
R2784 B.n674 B.n481 10.6151
R2785 B.n675 B.n674 10.6151
R2786 B.n676 B.n675 10.6151
R2787 B.n676 B.n479 10.6151
R2788 B.n682 B.n479 10.6151
R2789 B.n683 B.n682 10.6151
R2790 B.n684 B.n683 10.6151
R2791 B.n684 B.n477 10.6151
R2792 B.n690 B.n477 10.6151
R2793 B.n691 B.n690 10.6151
R2794 B.n692 B.n691 10.6151
R2795 B.n692 B.n475 10.6151
R2796 B.n698 B.n475 10.6151
R2797 B.n699 B.n698 10.6151
R2798 B.n700 B.n699 10.6151
R2799 B.n700 B.n473 10.6151
R2800 B.n706 B.n473 10.6151
R2801 B.n707 B.n706 10.6151
R2802 B.n708 B.n707 10.6151
R2803 B.n708 B.n471 10.6151
R2804 B.n714 B.n471 10.6151
R2805 B.n715 B.n714 10.6151
R2806 B.n716 B.n715 10.6151
R2807 B.n716 B.n469 10.6151
R2808 B.n722 B.n469 10.6151
R2809 B.n723 B.n722 10.6151
R2810 B.n724 B.n723 10.6151
R2811 B.n724 B.n467 10.6151
R2812 B.n730 B.n467 10.6151
R2813 B.n731 B.n730 10.6151
R2814 B.n732 B.n731 10.6151
R2815 B.n732 B.n465 10.6151
R2816 B.n738 B.n465 10.6151
R2817 B.n739 B.n738 10.6151
R2818 B.n740 B.n739 10.6151
R2819 B.n740 B.n463 10.6151
R2820 B.n746 B.n463 10.6151
R2821 B.n747 B.n746 10.6151
R2822 B.n748 B.n747 10.6151
R2823 B.n748 B.n461 10.6151
R2824 B.n754 B.n461 10.6151
R2825 B.n755 B.n754 10.6151
R2826 B.n756 B.n755 10.6151
R2827 B.n756 B.n459 10.6151
R2828 B.n762 B.n459 10.6151
R2829 B.n763 B.n762 10.6151
R2830 B.n764 B.n763 10.6151
R2831 B.n764 B.n457 10.6151
R2832 B.n457 B.n456 10.6151
R2833 B.n771 B.n456 10.6151
R2834 B.n772 B.n771 10.6151
R2835 B.n778 B.n777 10.6151
R2836 B.n779 B.n778 10.6151
R2837 B.n779 B.n444 10.6151
R2838 B.n789 B.n444 10.6151
R2839 B.n790 B.n789 10.6151
R2840 B.n791 B.n790 10.6151
R2841 B.n791 B.n436 10.6151
R2842 B.n801 B.n436 10.6151
R2843 B.n802 B.n801 10.6151
R2844 B.n803 B.n802 10.6151
R2845 B.n803 B.n428 10.6151
R2846 B.n813 B.n428 10.6151
R2847 B.n814 B.n813 10.6151
R2848 B.n815 B.n814 10.6151
R2849 B.n815 B.n420 10.6151
R2850 B.n825 B.n420 10.6151
R2851 B.n826 B.n825 10.6151
R2852 B.n827 B.n826 10.6151
R2853 B.n827 B.n412 10.6151
R2854 B.n837 B.n412 10.6151
R2855 B.n838 B.n837 10.6151
R2856 B.n839 B.n838 10.6151
R2857 B.n839 B.n404 10.6151
R2858 B.n849 B.n404 10.6151
R2859 B.n850 B.n849 10.6151
R2860 B.n851 B.n850 10.6151
R2861 B.n851 B.n396 10.6151
R2862 B.n862 B.n396 10.6151
R2863 B.n863 B.n862 10.6151
R2864 B.n864 B.n863 10.6151
R2865 B.n864 B.n389 10.6151
R2866 B.n875 B.n389 10.6151
R2867 B.n876 B.n875 10.6151
R2868 B.n877 B.n876 10.6151
R2869 B.n877 B.n0 10.6151
R2870 B.n1001 B.n1 10.6151
R2871 B.n1001 B.n1000 10.6151
R2872 B.n1000 B.n999 10.6151
R2873 B.n999 B.n10 10.6151
R2874 B.n993 B.n10 10.6151
R2875 B.n993 B.n992 10.6151
R2876 B.n992 B.n991 10.6151
R2877 B.n991 B.n16 10.6151
R2878 B.n985 B.n16 10.6151
R2879 B.n985 B.n984 10.6151
R2880 B.n984 B.n983 10.6151
R2881 B.n983 B.n24 10.6151
R2882 B.n977 B.n24 10.6151
R2883 B.n977 B.n976 10.6151
R2884 B.n976 B.n975 10.6151
R2885 B.n975 B.n31 10.6151
R2886 B.n969 B.n31 10.6151
R2887 B.n969 B.n968 10.6151
R2888 B.n968 B.n967 10.6151
R2889 B.n967 B.n38 10.6151
R2890 B.n961 B.n38 10.6151
R2891 B.n961 B.n960 10.6151
R2892 B.n960 B.n959 10.6151
R2893 B.n959 B.n45 10.6151
R2894 B.n953 B.n45 10.6151
R2895 B.n953 B.n952 10.6151
R2896 B.n952 B.n951 10.6151
R2897 B.n951 B.n52 10.6151
R2898 B.n945 B.n52 10.6151
R2899 B.n945 B.n944 10.6151
R2900 B.n944 B.n943 10.6151
R2901 B.n943 B.n59 10.6151
R2902 B.n937 B.n59 10.6151
R2903 B.n937 B.n936 10.6151
R2904 B.n936 B.n935 10.6151
R2905 B.n250 B.n137 9.36635
R2906 B.n273 B.n134 9.36635
R2907 B.n635 B.n634 9.36635
R2908 B.n659 B.n658 9.36635
R2909 B.n866 B.t3 8.65245
R2910 B.n995 B.t2 8.65245
R2911 B.n799 B.t5 3.84581
R2912 B.n949 B.t9 3.84581
R2913 B.n1007 B.n0 2.81026
R2914 B.n1007 B.n1 2.81026
R2915 B.n253 B.n137 1.24928
R2916 B.n270 B.n134 1.24928
R2917 B.n634 B.n491 1.24928
R2918 B.n658 B.n657 1.24928
R2919 VN.n0 VN.t1 184.751
R2920 VN.n1 VN.t0 184.751
R2921 VN.n0 VN.t3 183.856
R2922 VN.n1 VN.t2 183.856
R2923 VN VN.n1 55.0304
R2924 VN VN.n0 3.45085
R2925 VDD2.n2 VDD2.n0 109.522
R2926 VDD2.n2 VDD2.n1 62.4274
R2927 VDD2.n1 VDD2.t1 1.12486
R2928 VDD2.n1 VDD2.t3 1.12486
R2929 VDD2.n0 VDD2.t2 1.12486
R2930 VDD2.n0 VDD2.t0 1.12486
R2931 VDD2 VDD2.n2 0.0586897
C0 VN VTAIL 6.62394f
C1 VN VDD2 6.93431f
C2 VP VDD1 7.19387f
C3 VTAIL VP 6.63805f
C4 VP VDD2 0.409415f
C5 VN VP 7.40156f
C6 VTAIL VDD1 6.74203f
C7 VDD1 VDD2 1.08002f
C8 VTAIL VDD2 6.79785f
C9 VN VDD1 0.149055f
C10 VDD2 B 4.340229f
C11 VDD1 B 9.12374f
C12 VTAIL B 13.593377f
C13 VN B 11.59952f
C14 VP B 9.817331f
C15 VDD2.t2 B 0.368691f
C16 VDD2.t0 B 0.368691f
C17 VDD2.n0 B 4.23647f
C18 VDD2.t1 B 0.368691f
C19 VDD2.t3 B 0.368691f
C20 VDD2.n1 B 3.3578f
C21 VDD2.n2 B 4.39197f
C22 VN.t1 B 3.37712f
C23 VN.t3 B 3.37124f
C24 VN.n0 B 2.1387f
C25 VN.t0 B 3.37712f
C26 VN.t2 B 3.37124f
C27 VN.n1 B 3.59619f
C28 VTAIL.n0 B 0.022161f
C29 VTAIL.n1 B 0.015397f
C30 VTAIL.n2 B 0.008274f
C31 VTAIL.n3 B 0.019556f
C32 VTAIL.n4 B 0.00876f
C33 VTAIL.n5 B 0.015397f
C34 VTAIL.n6 B 0.008274f
C35 VTAIL.n7 B 0.019556f
C36 VTAIL.n8 B 0.008517f
C37 VTAIL.n9 B 0.015397f
C38 VTAIL.n10 B 0.00876f
C39 VTAIL.n11 B 0.019556f
C40 VTAIL.n12 B 0.00876f
C41 VTAIL.n13 B 0.015397f
C42 VTAIL.n14 B 0.008274f
C43 VTAIL.n15 B 0.019556f
C44 VTAIL.n16 B 0.00876f
C45 VTAIL.n17 B 0.015397f
C46 VTAIL.n18 B 0.008274f
C47 VTAIL.n19 B 0.019556f
C48 VTAIL.n20 B 0.00876f
C49 VTAIL.n21 B 0.015397f
C50 VTAIL.n22 B 0.008274f
C51 VTAIL.n23 B 0.019556f
C52 VTAIL.n24 B 0.00876f
C53 VTAIL.n25 B 0.015397f
C54 VTAIL.n26 B 0.008274f
C55 VTAIL.n27 B 0.019556f
C56 VTAIL.n28 B 0.00876f
C57 VTAIL.n29 B 1.18591f
C58 VTAIL.n30 B 0.008274f
C59 VTAIL.t2 B 0.032383f
C60 VTAIL.n31 B 0.110497f
C61 VTAIL.n32 B 0.011552f
C62 VTAIL.n33 B 0.014667f
C63 VTAIL.n34 B 0.019556f
C64 VTAIL.n35 B 0.00876f
C65 VTAIL.n36 B 0.008274f
C66 VTAIL.n37 B 0.015397f
C67 VTAIL.n38 B 0.015397f
C68 VTAIL.n39 B 0.008274f
C69 VTAIL.n40 B 0.00876f
C70 VTAIL.n41 B 0.019556f
C71 VTAIL.n42 B 0.019556f
C72 VTAIL.n43 B 0.00876f
C73 VTAIL.n44 B 0.008274f
C74 VTAIL.n45 B 0.015397f
C75 VTAIL.n46 B 0.015397f
C76 VTAIL.n47 B 0.008274f
C77 VTAIL.n48 B 0.00876f
C78 VTAIL.n49 B 0.019556f
C79 VTAIL.n50 B 0.019556f
C80 VTAIL.n51 B 0.00876f
C81 VTAIL.n52 B 0.008274f
C82 VTAIL.n53 B 0.015397f
C83 VTAIL.n54 B 0.015397f
C84 VTAIL.n55 B 0.008274f
C85 VTAIL.n56 B 0.00876f
C86 VTAIL.n57 B 0.019556f
C87 VTAIL.n58 B 0.019556f
C88 VTAIL.n59 B 0.00876f
C89 VTAIL.n60 B 0.008274f
C90 VTAIL.n61 B 0.015397f
C91 VTAIL.n62 B 0.015397f
C92 VTAIL.n63 B 0.008274f
C93 VTAIL.n64 B 0.00876f
C94 VTAIL.n65 B 0.019556f
C95 VTAIL.n66 B 0.019556f
C96 VTAIL.n67 B 0.00876f
C97 VTAIL.n68 B 0.008274f
C98 VTAIL.n69 B 0.015397f
C99 VTAIL.n70 B 0.015397f
C100 VTAIL.n71 B 0.008274f
C101 VTAIL.n72 B 0.008274f
C102 VTAIL.n73 B 0.00876f
C103 VTAIL.n74 B 0.019556f
C104 VTAIL.n75 B 0.019556f
C105 VTAIL.n76 B 0.019556f
C106 VTAIL.n77 B 0.008517f
C107 VTAIL.n78 B 0.008274f
C108 VTAIL.n79 B 0.015397f
C109 VTAIL.n80 B 0.015397f
C110 VTAIL.n81 B 0.008274f
C111 VTAIL.n82 B 0.00876f
C112 VTAIL.n83 B 0.019556f
C113 VTAIL.n84 B 0.019556f
C114 VTAIL.n85 B 0.00876f
C115 VTAIL.n86 B 0.008274f
C116 VTAIL.n87 B 0.015397f
C117 VTAIL.n88 B 0.015397f
C118 VTAIL.n89 B 0.008274f
C119 VTAIL.n90 B 0.00876f
C120 VTAIL.n91 B 0.019556f
C121 VTAIL.n92 B 0.043253f
C122 VTAIL.n93 B 0.00876f
C123 VTAIL.n94 B 0.008274f
C124 VTAIL.n95 B 0.037482f
C125 VTAIL.n96 B 0.024353f
C126 VTAIL.n97 B 0.108204f
C127 VTAIL.n98 B 0.022161f
C128 VTAIL.n99 B 0.015397f
C129 VTAIL.n100 B 0.008274f
C130 VTAIL.n101 B 0.019556f
C131 VTAIL.n102 B 0.00876f
C132 VTAIL.n103 B 0.015397f
C133 VTAIL.n104 B 0.008274f
C134 VTAIL.n105 B 0.019556f
C135 VTAIL.n106 B 0.008517f
C136 VTAIL.n107 B 0.015397f
C137 VTAIL.n108 B 0.00876f
C138 VTAIL.n109 B 0.019556f
C139 VTAIL.n110 B 0.00876f
C140 VTAIL.n111 B 0.015397f
C141 VTAIL.n112 B 0.008274f
C142 VTAIL.n113 B 0.019556f
C143 VTAIL.n114 B 0.00876f
C144 VTAIL.n115 B 0.015397f
C145 VTAIL.n116 B 0.008274f
C146 VTAIL.n117 B 0.019556f
C147 VTAIL.n118 B 0.00876f
C148 VTAIL.n119 B 0.015397f
C149 VTAIL.n120 B 0.008274f
C150 VTAIL.n121 B 0.019556f
C151 VTAIL.n122 B 0.00876f
C152 VTAIL.n123 B 0.015397f
C153 VTAIL.n124 B 0.008274f
C154 VTAIL.n125 B 0.019556f
C155 VTAIL.n126 B 0.00876f
C156 VTAIL.n127 B 1.18591f
C157 VTAIL.n128 B 0.008274f
C158 VTAIL.t5 B 0.032383f
C159 VTAIL.n129 B 0.110497f
C160 VTAIL.n130 B 0.011552f
C161 VTAIL.n131 B 0.014667f
C162 VTAIL.n132 B 0.019556f
C163 VTAIL.n133 B 0.00876f
C164 VTAIL.n134 B 0.008274f
C165 VTAIL.n135 B 0.015397f
C166 VTAIL.n136 B 0.015397f
C167 VTAIL.n137 B 0.008274f
C168 VTAIL.n138 B 0.00876f
C169 VTAIL.n139 B 0.019556f
C170 VTAIL.n140 B 0.019556f
C171 VTAIL.n141 B 0.00876f
C172 VTAIL.n142 B 0.008274f
C173 VTAIL.n143 B 0.015397f
C174 VTAIL.n144 B 0.015397f
C175 VTAIL.n145 B 0.008274f
C176 VTAIL.n146 B 0.00876f
C177 VTAIL.n147 B 0.019556f
C178 VTAIL.n148 B 0.019556f
C179 VTAIL.n149 B 0.00876f
C180 VTAIL.n150 B 0.008274f
C181 VTAIL.n151 B 0.015397f
C182 VTAIL.n152 B 0.015397f
C183 VTAIL.n153 B 0.008274f
C184 VTAIL.n154 B 0.00876f
C185 VTAIL.n155 B 0.019556f
C186 VTAIL.n156 B 0.019556f
C187 VTAIL.n157 B 0.00876f
C188 VTAIL.n158 B 0.008274f
C189 VTAIL.n159 B 0.015397f
C190 VTAIL.n160 B 0.015397f
C191 VTAIL.n161 B 0.008274f
C192 VTAIL.n162 B 0.00876f
C193 VTAIL.n163 B 0.019556f
C194 VTAIL.n164 B 0.019556f
C195 VTAIL.n165 B 0.00876f
C196 VTAIL.n166 B 0.008274f
C197 VTAIL.n167 B 0.015397f
C198 VTAIL.n168 B 0.015397f
C199 VTAIL.n169 B 0.008274f
C200 VTAIL.n170 B 0.008274f
C201 VTAIL.n171 B 0.00876f
C202 VTAIL.n172 B 0.019556f
C203 VTAIL.n173 B 0.019556f
C204 VTAIL.n174 B 0.019556f
C205 VTAIL.n175 B 0.008517f
C206 VTAIL.n176 B 0.008274f
C207 VTAIL.n177 B 0.015397f
C208 VTAIL.n178 B 0.015397f
C209 VTAIL.n179 B 0.008274f
C210 VTAIL.n180 B 0.00876f
C211 VTAIL.n181 B 0.019556f
C212 VTAIL.n182 B 0.019556f
C213 VTAIL.n183 B 0.00876f
C214 VTAIL.n184 B 0.008274f
C215 VTAIL.n185 B 0.015397f
C216 VTAIL.n186 B 0.015397f
C217 VTAIL.n187 B 0.008274f
C218 VTAIL.n188 B 0.00876f
C219 VTAIL.n189 B 0.019556f
C220 VTAIL.n190 B 0.043253f
C221 VTAIL.n191 B 0.00876f
C222 VTAIL.n192 B 0.008274f
C223 VTAIL.n193 B 0.037482f
C224 VTAIL.n194 B 0.024353f
C225 VTAIL.n195 B 0.173106f
C226 VTAIL.n196 B 0.022161f
C227 VTAIL.n197 B 0.015397f
C228 VTAIL.n198 B 0.008274f
C229 VTAIL.n199 B 0.019556f
C230 VTAIL.n200 B 0.00876f
C231 VTAIL.n201 B 0.015397f
C232 VTAIL.n202 B 0.008274f
C233 VTAIL.n203 B 0.019556f
C234 VTAIL.n204 B 0.008517f
C235 VTAIL.n205 B 0.015397f
C236 VTAIL.n206 B 0.00876f
C237 VTAIL.n207 B 0.019556f
C238 VTAIL.n208 B 0.00876f
C239 VTAIL.n209 B 0.015397f
C240 VTAIL.n210 B 0.008274f
C241 VTAIL.n211 B 0.019556f
C242 VTAIL.n212 B 0.00876f
C243 VTAIL.n213 B 0.015397f
C244 VTAIL.n214 B 0.008274f
C245 VTAIL.n215 B 0.019556f
C246 VTAIL.n216 B 0.00876f
C247 VTAIL.n217 B 0.015397f
C248 VTAIL.n218 B 0.008274f
C249 VTAIL.n219 B 0.019556f
C250 VTAIL.n220 B 0.00876f
C251 VTAIL.n221 B 0.015397f
C252 VTAIL.n222 B 0.008274f
C253 VTAIL.n223 B 0.019556f
C254 VTAIL.n224 B 0.00876f
C255 VTAIL.n225 B 1.18591f
C256 VTAIL.n226 B 0.008274f
C257 VTAIL.t4 B 0.032383f
C258 VTAIL.n227 B 0.110497f
C259 VTAIL.n228 B 0.011552f
C260 VTAIL.n229 B 0.014667f
C261 VTAIL.n230 B 0.019556f
C262 VTAIL.n231 B 0.00876f
C263 VTAIL.n232 B 0.008274f
C264 VTAIL.n233 B 0.015397f
C265 VTAIL.n234 B 0.015397f
C266 VTAIL.n235 B 0.008274f
C267 VTAIL.n236 B 0.00876f
C268 VTAIL.n237 B 0.019556f
C269 VTAIL.n238 B 0.019556f
C270 VTAIL.n239 B 0.00876f
C271 VTAIL.n240 B 0.008274f
C272 VTAIL.n241 B 0.015397f
C273 VTAIL.n242 B 0.015397f
C274 VTAIL.n243 B 0.008274f
C275 VTAIL.n244 B 0.00876f
C276 VTAIL.n245 B 0.019556f
C277 VTAIL.n246 B 0.019556f
C278 VTAIL.n247 B 0.00876f
C279 VTAIL.n248 B 0.008274f
C280 VTAIL.n249 B 0.015397f
C281 VTAIL.n250 B 0.015397f
C282 VTAIL.n251 B 0.008274f
C283 VTAIL.n252 B 0.00876f
C284 VTAIL.n253 B 0.019556f
C285 VTAIL.n254 B 0.019556f
C286 VTAIL.n255 B 0.00876f
C287 VTAIL.n256 B 0.008274f
C288 VTAIL.n257 B 0.015397f
C289 VTAIL.n258 B 0.015397f
C290 VTAIL.n259 B 0.008274f
C291 VTAIL.n260 B 0.00876f
C292 VTAIL.n261 B 0.019556f
C293 VTAIL.n262 B 0.019556f
C294 VTAIL.n263 B 0.00876f
C295 VTAIL.n264 B 0.008274f
C296 VTAIL.n265 B 0.015397f
C297 VTAIL.n266 B 0.015397f
C298 VTAIL.n267 B 0.008274f
C299 VTAIL.n268 B 0.008274f
C300 VTAIL.n269 B 0.00876f
C301 VTAIL.n270 B 0.019556f
C302 VTAIL.n271 B 0.019556f
C303 VTAIL.n272 B 0.019556f
C304 VTAIL.n273 B 0.008517f
C305 VTAIL.n274 B 0.008274f
C306 VTAIL.n275 B 0.015397f
C307 VTAIL.n276 B 0.015397f
C308 VTAIL.n277 B 0.008274f
C309 VTAIL.n278 B 0.00876f
C310 VTAIL.n279 B 0.019556f
C311 VTAIL.n280 B 0.019556f
C312 VTAIL.n281 B 0.00876f
C313 VTAIL.n282 B 0.008274f
C314 VTAIL.n283 B 0.015397f
C315 VTAIL.n284 B 0.015397f
C316 VTAIL.n285 B 0.008274f
C317 VTAIL.n286 B 0.00876f
C318 VTAIL.n287 B 0.019556f
C319 VTAIL.n288 B 0.043253f
C320 VTAIL.n289 B 0.00876f
C321 VTAIL.n290 B 0.008274f
C322 VTAIL.n291 B 0.037482f
C323 VTAIL.n292 B 0.024353f
C324 VTAIL.n293 B 1.24768f
C325 VTAIL.n294 B 0.022161f
C326 VTAIL.n295 B 0.015397f
C327 VTAIL.n296 B 0.008274f
C328 VTAIL.n297 B 0.019556f
C329 VTAIL.n298 B 0.00876f
C330 VTAIL.n299 B 0.015397f
C331 VTAIL.n300 B 0.008274f
C332 VTAIL.n301 B 0.019556f
C333 VTAIL.n302 B 0.008517f
C334 VTAIL.n303 B 0.015397f
C335 VTAIL.n304 B 0.008517f
C336 VTAIL.n305 B 0.008274f
C337 VTAIL.n306 B 0.019556f
C338 VTAIL.n307 B 0.019556f
C339 VTAIL.n308 B 0.00876f
C340 VTAIL.n309 B 0.015397f
C341 VTAIL.n310 B 0.008274f
C342 VTAIL.n311 B 0.019556f
C343 VTAIL.n312 B 0.00876f
C344 VTAIL.n313 B 0.015397f
C345 VTAIL.n314 B 0.008274f
C346 VTAIL.n315 B 0.019556f
C347 VTAIL.n316 B 0.00876f
C348 VTAIL.n317 B 0.015397f
C349 VTAIL.n318 B 0.008274f
C350 VTAIL.n319 B 0.019556f
C351 VTAIL.n320 B 0.00876f
C352 VTAIL.n321 B 0.015397f
C353 VTAIL.n322 B 0.008274f
C354 VTAIL.n323 B 0.019556f
C355 VTAIL.n324 B 0.00876f
C356 VTAIL.n325 B 1.18591f
C357 VTAIL.n326 B 0.008274f
C358 VTAIL.t0 B 0.032383f
C359 VTAIL.n327 B 0.110497f
C360 VTAIL.n328 B 0.011552f
C361 VTAIL.n329 B 0.014667f
C362 VTAIL.n330 B 0.019556f
C363 VTAIL.n331 B 0.00876f
C364 VTAIL.n332 B 0.008274f
C365 VTAIL.n333 B 0.015397f
C366 VTAIL.n334 B 0.015397f
C367 VTAIL.n335 B 0.008274f
C368 VTAIL.n336 B 0.00876f
C369 VTAIL.n337 B 0.019556f
C370 VTAIL.n338 B 0.019556f
C371 VTAIL.n339 B 0.00876f
C372 VTAIL.n340 B 0.008274f
C373 VTAIL.n341 B 0.015397f
C374 VTAIL.n342 B 0.015397f
C375 VTAIL.n343 B 0.008274f
C376 VTAIL.n344 B 0.00876f
C377 VTAIL.n345 B 0.019556f
C378 VTAIL.n346 B 0.019556f
C379 VTAIL.n347 B 0.00876f
C380 VTAIL.n348 B 0.008274f
C381 VTAIL.n349 B 0.015397f
C382 VTAIL.n350 B 0.015397f
C383 VTAIL.n351 B 0.008274f
C384 VTAIL.n352 B 0.00876f
C385 VTAIL.n353 B 0.019556f
C386 VTAIL.n354 B 0.019556f
C387 VTAIL.n355 B 0.00876f
C388 VTAIL.n356 B 0.008274f
C389 VTAIL.n357 B 0.015397f
C390 VTAIL.n358 B 0.015397f
C391 VTAIL.n359 B 0.008274f
C392 VTAIL.n360 B 0.00876f
C393 VTAIL.n361 B 0.019556f
C394 VTAIL.n362 B 0.019556f
C395 VTAIL.n363 B 0.00876f
C396 VTAIL.n364 B 0.008274f
C397 VTAIL.n365 B 0.015397f
C398 VTAIL.n366 B 0.015397f
C399 VTAIL.n367 B 0.008274f
C400 VTAIL.n368 B 0.00876f
C401 VTAIL.n369 B 0.019556f
C402 VTAIL.n370 B 0.019556f
C403 VTAIL.n371 B 0.00876f
C404 VTAIL.n372 B 0.008274f
C405 VTAIL.n373 B 0.015397f
C406 VTAIL.n374 B 0.015397f
C407 VTAIL.n375 B 0.008274f
C408 VTAIL.n376 B 0.00876f
C409 VTAIL.n377 B 0.019556f
C410 VTAIL.n378 B 0.019556f
C411 VTAIL.n379 B 0.00876f
C412 VTAIL.n380 B 0.008274f
C413 VTAIL.n381 B 0.015397f
C414 VTAIL.n382 B 0.015397f
C415 VTAIL.n383 B 0.008274f
C416 VTAIL.n384 B 0.00876f
C417 VTAIL.n385 B 0.019556f
C418 VTAIL.n386 B 0.043253f
C419 VTAIL.n387 B 0.00876f
C420 VTAIL.n388 B 0.008274f
C421 VTAIL.n389 B 0.037482f
C422 VTAIL.n390 B 0.024353f
C423 VTAIL.n391 B 1.24768f
C424 VTAIL.n392 B 0.022161f
C425 VTAIL.n393 B 0.015397f
C426 VTAIL.n394 B 0.008274f
C427 VTAIL.n395 B 0.019556f
C428 VTAIL.n396 B 0.00876f
C429 VTAIL.n397 B 0.015397f
C430 VTAIL.n398 B 0.008274f
C431 VTAIL.n399 B 0.019556f
C432 VTAIL.n400 B 0.008517f
C433 VTAIL.n401 B 0.015397f
C434 VTAIL.n402 B 0.008517f
C435 VTAIL.n403 B 0.008274f
C436 VTAIL.n404 B 0.019556f
C437 VTAIL.n405 B 0.019556f
C438 VTAIL.n406 B 0.00876f
C439 VTAIL.n407 B 0.015397f
C440 VTAIL.n408 B 0.008274f
C441 VTAIL.n409 B 0.019556f
C442 VTAIL.n410 B 0.00876f
C443 VTAIL.n411 B 0.015397f
C444 VTAIL.n412 B 0.008274f
C445 VTAIL.n413 B 0.019556f
C446 VTAIL.n414 B 0.00876f
C447 VTAIL.n415 B 0.015397f
C448 VTAIL.n416 B 0.008274f
C449 VTAIL.n417 B 0.019556f
C450 VTAIL.n418 B 0.00876f
C451 VTAIL.n419 B 0.015397f
C452 VTAIL.n420 B 0.008274f
C453 VTAIL.n421 B 0.019556f
C454 VTAIL.n422 B 0.00876f
C455 VTAIL.n423 B 1.18591f
C456 VTAIL.n424 B 0.008274f
C457 VTAIL.t3 B 0.032383f
C458 VTAIL.n425 B 0.110497f
C459 VTAIL.n426 B 0.011552f
C460 VTAIL.n427 B 0.014667f
C461 VTAIL.n428 B 0.019556f
C462 VTAIL.n429 B 0.00876f
C463 VTAIL.n430 B 0.008274f
C464 VTAIL.n431 B 0.015397f
C465 VTAIL.n432 B 0.015397f
C466 VTAIL.n433 B 0.008274f
C467 VTAIL.n434 B 0.00876f
C468 VTAIL.n435 B 0.019556f
C469 VTAIL.n436 B 0.019556f
C470 VTAIL.n437 B 0.00876f
C471 VTAIL.n438 B 0.008274f
C472 VTAIL.n439 B 0.015397f
C473 VTAIL.n440 B 0.015397f
C474 VTAIL.n441 B 0.008274f
C475 VTAIL.n442 B 0.00876f
C476 VTAIL.n443 B 0.019556f
C477 VTAIL.n444 B 0.019556f
C478 VTAIL.n445 B 0.00876f
C479 VTAIL.n446 B 0.008274f
C480 VTAIL.n447 B 0.015397f
C481 VTAIL.n448 B 0.015397f
C482 VTAIL.n449 B 0.008274f
C483 VTAIL.n450 B 0.00876f
C484 VTAIL.n451 B 0.019556f
C485 VTAIL.n452 B 0.019556f
C486 VTAIL.n453 B 0.00876f
C487 VTAIL.n454 B 0.008274f
C488 VTAIL.n455 B 0.015397f
C489 VTAIL.n456 B 0.015397f
C490 VTAIL.n457 B 0.008274f
C491 VTAIL.n458 B 0.00876f
C492 VTAIL.n459 B 0.019556f
C493 VTAIL.n460 B 0.019556f
C494 VTAIL.n461 B 0.00876f
C495 VTAIL.n462 B 0.008274f
C496 VTAIL.n463 B 0.015397f
C497 VTAIL.n464 B 0.015397f
C498 VTAIL.n465 B 0.008274f
C499 VTAIL.n466 B 0.00876f
C500 VTAIL.n467 B 0.019556f
C501 VTAIL.n468 B 0.019556f
C502 VTAIL.n469 B 0.00876f
C503 VTAIL.n470 B 0.008274f
C504 VTAIL.n471 B 0.015397f
C505 VTAIL.n472 B 0.015397f
C506 VTAIL.n473 B 0.008274f
C507 VTAIL.n474 B 0.00876f
C508 VTAIL.n475 B 0.019556f
C509 VTAIL.n476 B 0.019556f
C510 VTAIL.n477 B 0.00876f
C511 VTAIL.n478 B 0.008274f
C512 VTAIL.n479 B 0.015397f
C513 VTAIL.n480 B 0.015397f
C514 VTAIL.n481 B 0.008274f
C515 VTAIL.n482 B 0.00876f
C516 VTAIL.n483 B 0.019556f
C517 VTAIL.n484 B 0.043253f
C518 VTAIL.n485 B 0.00876f
C519 VTAIL.n486 B 0.008274f
C520 VTAIL.n487 B 0.037482f
C521 VTAIL.n488 B 0.024353f
C522 VTAIL.n489 B 0.173106f
C523 VTAIL.n490 B 0.022161f
C524 VTAIL.n491 B 0.015397f
C525 VTAIL.n492 B 0.008274f
C526 VTAIL.n493 B 0.019556f
C527 VTAIL.n494 B 0.00876f
C528 VTAIL.n495 B 0.015397f
C529 VTAIL.n496 B 0.008274f
C530 VTAIL.n497 B 0.019556f
C531 VTAIL.n498 B 0.008517f
C532 VTAIL.n499 B 0.015397f
C533 VTAIL.n500 B 0.008517f
C534 VTAIL.n501 B 0.008274f
C535 VTAIL.n502 B 0.019556f
C536 VTAIL.n503 B 0.019556f
C537 VTAIL.n504 B 0.00876f
C538 VTAIL.n505 B 0.015397f
C539 VTAIL.n506 B 0.008274f
C540 VTAIL.n507 B 0.019556f
C541 VTAIL.n508 B 0.00876f
C542 VTAIL.n509 B 0.015397f
C543 VTAIL.n510 B 0.008274f
C544 VTAIL.n511 B 0.019556f
C545 VTAIL.n512 B 0.00876f
C546 VTAIL.n513 B 0.015397f
C547 VTAIL.n514 B 0.008274f
C548 VTAIL.n515 B 0.019556f
C549 VTAIL.n516 B 0.00876f
C550 VTAIL.n517 B 0.015397f
C551 VTAIL.n518 B 0.008274f
C552 VTAIL.n519 B 0.019556f
C553 VTAIL.n520 B 0.00876f
C554 VTAIL.n521 B 1.18591f
C555 VTAIL.n522 B 0.008274f
C556 VTAIL.t7 B 0.032383f
C557 VTAIL.n523 B 0.110497f
C558 VTAIL.n524 B 0.011552f
C559 VTAIL.n525 B 0.014667f
C560 VTAIL.n526 B 0.019556f
C561 VTAIL.n527 B 0.00876f
C562 VTAIL.n528 B 0.008274f
C563 VTAIL.n529 B 0.015397f
C564 VTAIL.n530 B 0.015397f
C565 VTAIL.n531 B 0.008274f
C566 VTAIL.n532 B 0.00876f
C567 VTAIL.n533 B 0.019556f
C568 VTAIL.n534 B 0.019556f
C569 VTAIL.n535 B 0.00876f
C570 VTAIL.n536 B 0.008274f
C571 VTAIL.n537 B 0.015397f
C572 VTAIL.n538 B 0.015397f
C573 VTAIL.n539 B 0.008274f
C574 VTAIL.n540 B 0.00876f
C575 VTAIL.n541 B 0.019556f
C576 VTAIL.n542 B 0.019556f
C577 VTAIL.n543 B 0.00876f
C578 VTAIL.n544 B 0.008274f
C579 VTAIL.n545 B 0.015397f
C580 VTAIL.n546 B 0.015397f
C581 VTAIL.n547 B 0.008274f
C582 VTAIL.n548 B 0.00876f
C583 VTAIL.n549 B 0.019556f
C584 VTAIL.n550 B 0.019556f
C585 VTAIL.n551 B 0.00876f
C586 VTAIL.n552 B 0.008274f
C587 VTAIL.n553 B 0.015397f
C588 VTAIL.n554 B 0.015397f
C589 VTAIL.n555 B 0.008274f
C590 VTAIL.n556 B 0.00876f
C591 VTAIL.n557 B 0.019556f
C592 VTAIL.n558 B 0.019556f
C593 VTAIL.n559 B 0.00876f
C594 VTAIL.n560 B 0.008274f
C595 VTAIL.n561 B 0.015397f
C596 VTAIL.n562 B 0.015397f
C597 VTAIL.n563 B 0.008274f
C598 VTAIL.n564 B 0.00876f
C599 VTAIL.n565 B 0.019556f
C600 VTAIL.n566 B 0.019556f
C601 VTAIL.n567 B 0.00876f
C602 VTAIL.n568 B 0.008274f
C603 VTAIL.n569 B 0.015397f
C604 VTAIL.n570 B 0.015397f
C605 VTAIL.n571 B 0.008274f
C606 VTAIL.n572 B 0.00876f
C607 VTAIL.n573 B 0.019556f
C608 VTAIL.n574 B 0.019556f
C609 VTAIL.n575 B 0.00876f
C610 VTAIL.n576 B 0.008274f
C611 VTAIL.n577 B 0.015397f
C612 VTAIL.n578 B 0.015397f
C613 VTAIL.n579 B 0.008274f
C614 VTAIL.n580 B 0.00876f
C615 VTAIL.n581 B 0.019556f
C616 VTAIL.n582 B 0.043253f
C617 VTAIL.n583 B 0.00876f
C618 VTAIL.n584 B 0.008274f
C619 VTAIL.n585 B 0.037482f
C620 VTAIL.n586 B 0.024353f
C621 VTAIL.n587 B 0.173106f
C622 VTAIL.n588 B 0.022161f
C623 VTAIL.n589 B 0.015397f
C624 VTAIL.n590 B 0.008274f
C625 VTAIL.n591 B 0.019556f
C626 VTAIL.n592 B 0.00876f
C627 VTAIL.n593 B 0.015397f
C628 VTAIL.n594 B 0.008274f
C629 VTAIL.n595 B 0.019556f
C630 VTAIL.n596 B 0.008517f
C631 VTAIL.n597 B 0.015397f
C632 VTAIL.n598 B 0.008517f
C633 VTAIL.n599 B 0.008274f
C634 VTAIL.n600 B 0.019556f
C635 VTAIL.n601 B 0.019556f
C636 VTAIL.n602 B 0.00876f
C637 VTAIL.n603 B 0.015397f
C638 VTAIL.n604 B 0.008274f
C639 VTAIL.n605 B 0.019556f
C640 VTAIL.n606 B 0.00876f
C641 VTAIL.n607 B 0.015397f
C642 VTAIL.n608 B 0.008274f
C643 VTAIL.n609 B 0.019556f
C644 VTAIL.n610 B 0.00876f
C645 VTAIL.n611 B 0.015397f
C646 VTAIL.n612 B 0.008274f
C647 VTAIL.n613 B 0.019556f
C648 VTAIL.n614 B 0.00876f
C649 VTAIL.n615 B 0.015397f
C650 VTAIL.n616 B 0.008274f
C651 VTAIL.n617 B 0.019556f
C652 VTAIL.n618 B 0.00876f
C653 VTAIL.n619 B 1.18591f
C654 VTAIL.n620 B 0.008274f
C655 VTAIL.t6 B 0.032383f
C656 VTAIL.n621 B 0.110497f
C657 VTAIL.n622 B 0.011552f
C658 VTAIL.n623 B 0.014667f
C659 VTAIL.n624 B 0.019556f
C660 VTAIL.n625 B 0.00876f
C661 VTAIL.n626 B 0.008274f
C662 VTAIL.n627 B 0.015397f
C663 VTAIL.n628 B 0.015397f
C664 VTAIL.n629 B 0.008274f
C665 VTAIL.n630 B 0.00876f
C666 VTAIL.n631 B 0.019556f
C667 VTAIL.n632 B 0.019556f
C668 VTAIL.n633 B 0.00876f
C669 VTAIL.n634 B 0.008274f
C670 VTAIL.n635 B 0.015397f
C671 VTAIL.n636 B 0.015397f
C672 VTAIL.n637 B 0.008274f
C673 VTAIL.n638 B 0.00876f
C674 VTAIL.n639 B 0.019556f
C675 VTAIL.n640 B 0.019556f
C676 VTAIL.n641 B 0.00876f
C677 VTAIL.n642 B 0.008274f
C678 VTAIL.n643 B 0.015397f
C679 VTAIL.n644 B 0.015397f
C680 VTAIL.n645 B 0.008274f
C681 VTAIL.n646 B 0.00876f
C682 VTAIL.n647 B 0.019556f
C683 VTAIL.n648 B 0.019556f
C684 VTAIL.n649 B 0.00876f
C685 VTAIL.n650 B 0.008274f
C686 VTAIL.n651 B 0.015397f
C687 VTAIL.n652 B 0.015397f
C688 VTAIL.n653 B 0.008274f
C689 VTAIL.n654 B 0.00876f
C690 VTAIL.n655 B 0.019556f
C691 VTAIL.n656 B 0.019556f
C692 VTAIL.n657 B 0.00876f
C693 VTAIL.n658 B 0.008274f
C694 VTAIL.n659 B 0.015397f
C695 VTAIL.n660 B 0.015397f
C696 VTAIL.n661 B 0.008274f
C697 VTAIL.n662 B 0.00876f
C698 VTAIL.n663 B 0.019556f
C699 VTAIL.n664 B 0.019556f
C700 VTAIL.n665 B 0.00876f
C701 VTAIL.n666 B 0.008274f
C702 VTAIL.n667 B 0.015397f
C703 VTAIL.n668 B 0.015397f
C704 VTAIL.n669 B 0.008274f
C705 VTAIL.n670 B 0.00876f
C706 VTAIL.n671 B 0.019556f
C707 VTAIL.n672 B 0.019556f
C708 VTAIL.n673 B 0.00876f
C709 VTAIL.n674 B 0.008274f
C710 VTAIL.n675 B 0.015397f
C711 VTAIL.n676 B 0.015397f
C712 VTAIL.n677 B 0.008274f
C713 VTAIL.n678 B 0.00876f
C714 VTAIL.n679 B 0.019556f
C715 VTAIL.n680 B 0.043253f
C716 VTAIL.n681 B 0.00876f
C717 VTAIL.n682 B 0.008274f
C718 VTAIL.n683 B 0.037482f
C719 VTAIL.n684 B 0.024353f
C720 VTAIL.n685 B 1.24768f
C721 VTAIL.n686 B 0.022161f
C722 VTAIL.n687 B 0.015397f
C723 VTAIL.n688 B 0.008274f
C724 VTAIL.n689 B 0.019556f
C725 VTAIL.n690 B 0.00876f
C726 VTAIL.n691 B 0.015397f
C727 VTAIL.n692 B 0.008274f
C728 VTAIL.n693 B 0.019556f
C729 VTAIL.n694 B 0.008517f
C730 VTAIL.n695 B 0.015397f
C731 VTAIL.n696 B 0.00876f
C732 VTAIL.n697 B 0.019556f
C733 VTAIL.n698 B 0.00876f
C734 VTAIL.n699 B 0.015397f
C735 VTAIL.n700 B 0.008274f
C736 VTAIL.n701 B 0.019556f
C737 VTAIL.n702 B 0.00876f
C738 VTAIL.n703 B 0.015397f
C739 VTAIL.n704 B 0.008274f
C740 VTAIL.n705 B 0.019556f
C741 VTAIL.n706 B 0.00876f
C742 VTAIL.n707 B 0.015397f
C743 VTAIL.n708 B 0.008274f
C744 VTAIL.n709 B 0.019556f
C745 VTAIL.n710 B 0.00876f
C746 VTAIL.n711 B 0.015397f
C747 VTAIL.n712 B 0.008274f
C748 VTAIL.n713 B 0.019556f
C749 VTAIL.n714 B 0.00876f
C750 VTAIL.n715 B 1.18591f
C751 VTAIL.n716 B 0.008274f
C752 VTAIL.t1 B 0.032383f
C753 VTAIL.n717 B 0.110497f
C754 VTAIL.n718 B 0.011552f
C755 VTAIL.n719 B 0.014667f
C756 VTAIL.n720 B 0.019556f
C757 VTAIL.n721 B 0.00876f
C758 VTAIL.n722 B 0.008274f
C759 VTAIL.n723 B 0.015397f
C760 VTAIL.n724 B 0.015397f
C761 VTAIL.n725 B 0.008274f
C762 VTAIL.n726 B 0.00876f
C763 VTAIL.n727 B 0.019556f
C764 VTAIL.n728 B 0.019556f
C765 VTAIL.n729 B 0.00876f
C766 VTAIL.n730 B 0.008274f
C767 VTAIL.n731 B 0.015397f
C768 VTAIL.n732 B 0.015397f
C769 VTAIL.n733 B 0.008274f
C770 VTAIL.n734 B 0.00876f
C771 VTAIL.n735 B 0.019556f
C772 VTAIL.n736 B 0.019556f
C773 VTAIL.n737 B 0.00876f
C774 VTAIL.n738 B 0.008274f
C775 VTAIL.n739 B 0.015397f
C776 VTAIL.n740 B 0.015397f
C777 VTAIL.n741 B 0.008274f
C778 VTAIL.n742 B 0.00876f
C779 VTAIL.n743 B 0.019556f
C780 VTAIL.n744 B 0.019556f
C781 VTAIL.n745 B 0.00876f
C782 VTAIL.n746 B 0.008274f
C783 VTAIL.n747 B 0.015397f
C784 VTAIL.n748 B 0.015397f
C785 VTAIL.n749 B 0.008274f
C786 VTAIL.n750 B 0.00876f
C787 VTAIL.n751 B 0.019556f
C788 VTAIL.n752 B 0.019556f
C789 VTAIL.n753 B 0.00876f
C790 VTAIL.n754 B 0.008274f
C791 VTAIL.n755 B 0.015397f
C792 VTAIL.n756 B 0.015397f
C793 VTAIL.n757 B 0.008274f
C794 VTAIL.n758 B 0.008274f
C795 VTAIL.n759 B 0.00876f
C796 VTAIL.n760 B 0.019556f
C797 VTAIL.n761 B 0.019556f
C798 VTAIL.n762 B 0.019556f
C799 VTAIL.n763 B 0.008517f
C800 VTAIL.n764 B 0.008274f
C801 VTAIL.n765 B 0.015397f
C802 VTAIL.n766 B 0.015397f
C803 VTAIL.n767 B 0.008274f
C804 VTAIL.n768 B 0.00876f
C805 VTAIL.n769 B 0.019556f
C806 VTAIL.n770 B 0.019556f
C807 VTAIL.n771 B 0.00876f
C808 VTAIL.n772 B 0.008274f
C809 VTAIL.n773 B 0.015397f
C810 VTAIL.n774 B 0.015397f
C811 VTAIL.n775 B 0.008274f
C812 VTAIL.n776 B 0.00876f
C813 VTAIL.n777 B 0.019556f
C814 VTAIL.n778 B 0.043253f
C815 VTAIL.n779 B 0.00876f
C816 VTAIL.n780 B 0.008274f
C817 VTAIL.n781 B 0.037482f
C818 VTAIL.n782 B 0.024353f
C819 VTAIL.n783 B 1.17701f
C820 VDD1.t2 B 0.37142f
C821 VDD1.t1 B 0.37142f
C822 VDD1.n0 B 3.3831f
C823 VDD1.t0 B 0.37142f
C824 VDD1.t3 B 0.37142f
C825 VDD1.n1 B 4.29611f
C826 VP.n0 B 0.030574f
C827 VP.t2 B 3.18873f
C828 VP.n1 B 0.04609f
C829 VP.n2 B 0.02319f
C830 VP.n3 B 0.025509f
C831 VP.t1 B 3.42489f
C832 VP.t0 B 3.43086f
C833 VP.n4 B 3.64127f
C834 VP.t3 B 3.18873f
C835 VP.n5 B 1.18248f
C836 VP.n6 B 1.46193f
C837 VP.n7 B 0.030574f
C838 VP.n8 B 0.02319f
C839 VP.n9 B 0.04322f
C840 VP.n10 B 0.04609f
C841 VP.n11 B 0.018747f
C842 VP.n12 B 0.02319f
C843 VP.n13 B 0.02319f
C844 VP.n14 B 0.02319f
C845 VP.n15 B 0.04322f
C846 VP.n16 B 0.025509f
C847 VP.n17 B 1.18248f
C848 VP.n18 B 0.042968f
.ends

