* NGSPICE file created from diff_pair_sample_0561.ext - technology: sky130A

.subckt diff_pair_sample_0561 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t9 VP.t0 VTAIL.t6 B.t9 sky130_fd_pr__nfet_01v8 ad=2.409 pd=14.93 as=2.409 ps=14.93 w=14.6 l=2.45
X1 VTAIL.t8 VP.t1 VDD1.t8 B.t2 sky130_fd_pr__nfet_01v8 ad=2.409 pd=14.93 as=2.409 ps=14.93 w=14.6 l=2.45
X2 VTAIL.t19 VN.t0 VDD2.t9 B.t8 sky130_fd_pr__nfet_01v8 ad=2.409 pd=14.93 as=2.409 ps=14.93 w=14.6 l=2.45
X3 VTAIL.t5 VP.t2 VDD1.t7 B.t0 sky130_fd_pr__nfet_01v8 ad=2.409 pd=14.93 as=2.409 ps=14.93 w=14.6 l=2.45
X4 VDD2.t8 VN.t1 VTAIL.t17 B.t4 sky130_fd_pr__nfet_01v8 ad=5.694 pd=29.98 as=2.409 ps=14.93 w=14.6 l=2.45
X5 VTAIL.t3 VN.t2 VDD2.t7 B.t3 sky130_fd_pr__nfet_01v8 ad=2.409 pd=14.93 as=2.409 ps=14.93 w=14.6 l=2.45
X6 VTAIL.t11 VP.t3 VDD1.t6 B.t8 sky130_fd_pr__nfet_01v8 ad=2.409 pd=14.93 as=2.409 ps=14.93 w=14.6 l=2.45
X7 VTAIL.t2 VN.t3 VDD2.t6 B.t2 sky130_fd_pr__nfet_01v8 ad=2.409 pd=14.93 as=2.409 ps=14.93 w=14.6 l=2.45
X8 VDD1.t5 VP.t4 VTAIL.t10 B.t7 sky130_fd_pr__nfet_01v8 ad=5.694 pd=29.98 as=2.409 ps=14.93 w=14.6 l=2.45
X9 B.t23 B.t21 B.t22 B.t18 sky130_fd_pr__nfet_01v8 ad=5.694 pd=29.98 as=0 ps=0 w=14.6 l=2.45
X10 VTAIL.t13 VP.t5 VDD1.t4 B.t3 sky130_fd_pr__nfet_01v8 ad=2.409 pd=14.93 as=2.409 ps=14.93 w=14.6 l=2.45
X11 B.t20 B.t17 B.t19 B.t18 sky130_fd_pr__nfet_01v8 ad=5.694 pd=29.98 as=0 ps=0 w=14.6 l=2.45
X12 VDD1.t3 VP.t6 VTAIL.t12 B.t6 sky130_fd_pr__nfet_01v8 ad=2.409 pd=14.93 as=2.409 ps=14.93 w=14.6 l=2.45
X13 VDD2.t5 VN.t4 VTAIL.t14 B.t6 sky130_fd_pr__nfet_01v8 ad=2.409 pd=14.93 as=2.409 ps=14.93 w=14.6 l=2.45
X14 VDD1.t2 VP.t7 VTAIL.t7 B.t5 sky130_fd_pr__nfet_01v8 ad=2.409 pd=14.93 as=5.694 ps=29.98 w=14.6 l=2.45
X15 VDD1.t1 VP.t8 VTAIL.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=5.694 pd=29.98 as=2.409 ps=14.93 w=14.6 l=2.45
X16 VDD1.t0 VP.t9 VTAIL.t9 B.t1 sky130_fd_pr__nfet_01v8 ad=2.409 pd=14.93 as=5.694 ps=29.98 w=14.6 l=2.45
X17 VDD2.t4 VN.t5 VTAIL.t15 B.t7 sky130_fd_pr__nfet_01v8 ad=5.694 pd=29.98 as=2.409 ps=14.93 w=14.6 l=2.45
X18 VDD2.t3 VN.t6 VTAIL.t16 B.t5 sky130_fd_pr__nfet_01v8 ad=2.409 pd=14.93 as=5.694 ps=29.98 w=14.6 l=2.45
X19 VDD2.t2 VN.t7 VTAIL.t18 B.t9 sky130_fd_pr__nfet_01v8 ad=2.409 pd=14.93 as=2.409 ps=14.93 w=14.6 l=2.45
X20 VDD2.t1 VN.t8 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=2.409 pd=14.93 as=5.694 ps=29.98 w=14.6 l=2.45
X21 B.t16 B.t14 B.t15 B.t11 sky130_fd_pr__nfet_01v8 ad=5.694 pd=29.98 as=0 ps=0 w=14.6 l=2.45
X22 VTAIL.t0 VN.t9 VDD2.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=2.409 pd=14.93 as=2.409 ps=14.93 w=14.6 l=2.45
X23 B.t13 B.t10 B.t12 B.t11 sky130_fd_pr__nfet_01v8 ad=5.694 pd=29.98 as=0 ps=0 w=14.6 l=2.45
R0 VP.n21 VP.t4 176.114
R1 VP.n23 VP.n20 161.3
R2 VP.n25 VP.n24 161.3
R3 VP.n26 VP.n19 161.3
R4 VP.n28 VP.n27 161.3
R5 VP.n29 VP.n18 161.3
R6 VP.n32 VP.n31 161.3
R7 VP.n33 VP.n17 161.3
R8 VP.n35 VP.n34 161.3
R9 VP.n36 VP.n16 161.3
R10 VP.n38 VP.n37 161.3
R11 VP.n39 VP.n15 161.3
R12 VP.n41 VP.n40 161.3
R13 VP.n43 VP.n14 161.3
R14 VP.n45 VP.n44 161.3
R15 VP.n46 VP.n13 161.3
R16 VP.n48 VP.n47 161.3
R17 VP.n49 VP.n12 161.3
R18 VP.n88 VP.n0 161.3
R19 VP.n87 VP.n86 161.3
R20 VP.n85 VP.n1 161.3
R21 VP.n84 VP.n83 161.3
R22 VP.n82 VP.n2 161.3
R23 VP.n80 VP.n79 161.3
R24 VP.n78 VP.n3 161.3
R25 VP.n77 VP.n76 161.3
R26 VP.n75 VP.n4 161.3
R27 VP.n74 VP.n73 161.3
R28 VP.n72 VP.n5 161.3
R29 VP.n71 VP.n70 161.3
R30 VP.n68 VP.n6 161.3
R31 VP.n67 VP.n66 161.3
R32 VP.n65 VP.n7 161.3
R33 VP.n64 VP.n63 161.3
R34 VP.n62 VP.n8 161.3
R35 VP.n60 VP.n59 161.3
R36 VP.n58 VP.n9 161.3
R37 VP.n57 VP.n56 161.3
R38 VP.n55 VP.n10 161.3
R39 VP.n54 VP.n53 161.3
R40 VP.n11 VP.t8 143.617
R41 VP.n61 VP.t3 143.617
R42 VP.n69 VP.t6 143.617
R43 VP.n81 VP.t2 143.617
R44 VP.n89 VP.t7 143.617
R45 VP.n50 VP.t9 143.617
R46 VP.n42 VP.t1 143.617
R47 VP.n30 VP.t0 143.617
R48 VP.n22 VP.t5 143.617
R49 VP.n52 VP.n11 95.6613
R50 VP.n90 VP.n89 95.6613
R51 VP.n51 VP.n50 95.6613
R52 VP.n22 VP.n21 71.1838
R53 VP.n52 VP.n51 54.333
R54 VP.n67 VP.n7 54.1398
R55 VP.n76 VP.n75 54.1398
R56 VP.n37 VP.n36 54.1398
R57 VP.n28 VP.n19 54.1398
R58 VP.n56 VP.n9 48.3272
R59 VP.n83 VP.n1 48.3272
R60 VP.n44 VP.n13 48.3272
R61 VP.n56 VP.n55 32.8269
R62 VP.n87 VP.n1 32.8269
R63 VP.n48 VP.n13 32.8269
R64 VP.n68 VP.n67 27.0143
R65 VP.n75 VP.n74 27.0143
R66 VP.n36 VP.n35 27.0143
R67 VP.n29 VP.n28 27.0143
R68 VP.n55 VP.n54 24.5923
R69 VP.n60 VP.n9 24.5923
R70 VP.n63 VP.n62 24.5923
R71 VP.n63 VP.n7 24.5923
R72 VP.n70 VP.n68 24.5923
R73 VP.n74 VP.n5 24.5923
R74 VP.n76 VP.n3 24.5923
R75 VP.n80 VP.n3 24.5923
R76 VP.n83 VP.n82 24.5923
R77 VP.n88 VP.n87 24.5923
R78 VP.n49 VP.n48 24.5923
R79 VP.n37 VP.n15 24.5923
R80 VP.n41 VP.n15 24.5923
R81 VP.n44 VP.n43 24.5923
R82 VP.n31 VP.n29 24.5923
R83 VP.n35 VP.n17 24.5923
R84 VP.n24 VP.n23 24.5923
R85 VP.n24 VP.n19 24.5923
R86 VP.n61 VP.n60 23.1168
R87 VP.n82 VP.n81 23.1168
R88 VP.n43 VP.n42 23.1168
R89 VP.n54 VP.n11 15.2474
R90 VP.n89 VP.n88 15.2474
R91 VP.n50 VP.n49 15.2474
R92 VP.n70 VP.n69 12.2964
R93 VP.n69 VP.n5 12.2964
R94 VP.n31 VP.n30 12.2964
R95 VP.n30 VP.n17 12.2964
R96 VP.n21 VP.n20 9.47955
R97 VP.n62 VP.n61 1.47601
R98 VP.n81 VP.n80 1.47601
R99 VP.n42 VP.n41 1.47601
R100 VP.n23 VP.n22 1.47601
R101 VP.n51 VP.n12 0.278335
R102 VP.n53 VP.n52 0.278335
R103 VP.n90 VP.n0 0.278335
R104 VP.n25 VP.n20 0.189894
R105 VP.n26 VP.n25 0.189894
R106 VP.n27 VP.n26 0.189894
R107 VP.n27 VP.n18 0.189894
R108 VP.n32 VP.n18 0.189894
R109 VP.n33 VP.n32 0.189894
R110 VP.n34 VP.n33 0.189894
R111 VP.n34 VP.n16 0.189894
R112 VP.n38 VP.n16 0.189894
R113 VP.n39 VP.n38 0.189894
R114 VP.n40 VP.n39 0.189894
R115 VP.n40 VP.n14 0.189894
R116 VP.n45 VP.n14 0.189894
R117 VP.n46 VP.n45 0.189894
R118 VP.n47 VP.n46 0.189894
R119 VP.n47 VP.n12 0.189894
R120 VP.n53 VP.n10 0.189894
R121 VP.n57 VP.n10 0.189894
R122 VP.n58 VP.n57 0.189894
R123 VP.n59 VP.n58 0.189894
R124 VP.n59 VP.n8 0.189894
R125 VP.n64 VP.n8 0.189894
R126 VP.n65 VP.n64 0.189894
R127 VP.n66 VP.n65 0.189894
R128 VP.n66 VP.n6 0.189894
R129 VP.n71 VP.n6 0.189894
R130 VP.n72 VP.n71 0.189894
R131 VP.n73 VP.n72 0.189894
R132 VP.n73 VP.n4 0.189894
R133 VP.n77 VP.n4 0.189894
R134 VP.n78 VP.n77 0.189894
R135 VP.n79 VP.n78 0.189894
R136 VP.n79 VP.n2 0.189894
R137 VP.n84 VP.n2 0.189894
R138 VP.n85 VP.n84 0.189894
R139 VP.n86 VP.n85 0.189894
R140 VP.n86 VP.n0 0.189894
R141 VP VP.n90 0.153485
R142 VTAIL.n11 VTAIL.t16 45.2741
R143 VTAIL.n16 VTAIL.t9 45.2741
R144 VTAIL.n17 VTAIL.t1 45.2739
R145 VTAIL.n2 VTAIL.t7 45.2739
R146 VTAIL.n15 VTAIL.n14 43.9179
R147 VTAIL.n13 VTAIL.n12 43.9179
R148 VTAIL.n10 VTAIL.n9 43.9179
R149 VTAIL.n8 VTAIL.n7 43.9179
R150 VTAIL.n19 VTAIL.n18 43.9179
R151 VTAIL.n1 VTAIL.n0 43.9179
R152 VTAIL.n4 VTAIL.n3 43.9179
R153 VTAIL.n6 VTAIL.n5 43.9179
R154 VTAIL.n8 VTAIL.n6 29.7462
R155 VTAIL.n17 VTAIL.n16 27.3496
R156 VTAIL.n10 VTAIL.n8 2.39705
R157 VTAIL.n11 VTAIL.n10 2.39705
R158 VTAIL.n15 VTAIL.n13 2.39705
R159 VTAIL.n16 VTAIL.n15 2.39705
R160 VTAIL.n6 VTAIL.n4 2.39705
R161 VTAIL.n4 VTAIL.n2 2.39705
R162 VTAIL.n19 VTAIL.n17 2.39705
R163 VTAIL VTAIL.n1 1.8561
R164 VTAIL.n13 VTAIL.n11 1.6686
R165 VTAIL.n2 VTAIL.n1 1.6686
R166 VTAIL.n18 VTAIL.t18 1.35666
R167 VTAIL.n18 VTAIL.t2 1.35666
R168 VTAIL.n0 VTAIL.t15 1.35666
R169 VTAIL.n0 VTAIL.t3 1.35666
R170 VTAIL.n3 VTAIL.t12 1.35666
R171 VTAIL.n3 VTAIL.t5 1.35666
R172 VTAIL.n5 VTAIL.t4 1.35666
R173 VTAIL.n5 VTAIL.t11 1.35666
R174 VTAIL.n14 VTAIL.t6 1.35666
R175 VTAIL.n14 VTAIL.t8 1.35666
R176 VTAIL.n12 VTAIL.t10 1.35666
R177 VTAIL.n12 VTAIL.t13 1.35666
R178 VTAIL.n9 VTAIL.t14 1.35666
R179 VTAIL.n9 VTAIL.t0 1.35666
R180 VTAIL.n7 VTAIL.t17 1.35666
R181 VTAIL.n7 VTAIL.t19 1.35666
R182 VTAIL VTAIL.n19 0.541448
R183 VDD1.n1 VDD1.t5 64.3494
R184 VDD1.n3 VDD1.t1 64.3492
R185 VDD1.n5 VDD1.n4 62.3387
R186 VDD1.n7 VDD1.n6 60.5967
R187 VDD1.n1 VDD1.n0 60.5967
R188 VDD1.n3 VDD1.n2 60.5967
R189 VDD1.n7 VDD1.n5 49.4664
R190 VDD1 VDD1.n7 1.73972
R191 VDD1.n6 VDD1.t8 1.35666
R192 VDD1.n6 VDD1.t0 1.35666
R193 VDD1.n0 VDD1.t4 1.35666
R194 VDD1.n0 VDD1.t9 1.35666
R195 VDD1.n4 VDD1.t7 1.35666
R196 VDD1.n4 VDD1.t2 1.35666
R197 VDD1.n2 VDD1.t6 1.35666
R198 VDD1.n2 VDD1.t3 1.35666
R199 VDD1 VDD1.n1 0.657828
R200 VDD1.n5 VDD1.n3 0.544292
R201 B.n1009 B.n1008 585
R202 B.n377 B.n158 585
R203 B.n376 B.n375 585
R204 B.n374 B.n373 585
R205 B.n372 B.n371 585
R206 B.n370 B.n369 585
R207 B.n368 B.n367 585
R208 B.n366 B.n365 585
R209 B.n364 B.n363 585
R210 B.n362 B.n361 585
R211 B.n360 B.n359 585
R212 B.n358 B.n357 585
R213 B.n356 B.n355 585
R214 B.n354 B.n353 585
R215 B.n352 B.n351 585
R216 B.n350 B.n349 585
R217 B.n348 B.n347 585
R218 B.n346 B.n345 585
R219 B.n344 B.n343 585
R220 B.n342 B.n341 585
R221 B.n340 B.n339 585
R222 B.n338 B.n337 585
R223 B.n336 B.n335 585
R224 B.n334 B.n333 585
R225 B.n332 B.n331 585
R226 B.n330 B.n329 585
R227 B.n328 B.n327 585
R228 B.n326 B.n325 585
R229 B.n324 B.n323 585
R230 B.n322 B.n321 585
R231 B.n320 B.n319 585
R232 B.n318 B.n317 585
R233 B.n316 B.n315 585
R234 B.n314 B.n313 585
R235 B.n312 B.n311 585
R236 B.n310 B.n309 585
R237 B.n308 B.n307 585
R238 B.n306 B.n305 585
R239 B.n304 B.n303 585
R240 B.n302 B.n301 585
R241 B.n300 B.n299 585
R242 B.n298 B.n297 585
R243 B.n296 B.n295 585
R244 B.n294 B.n293 585
R245 B.n292 B.n291 585
R246 B.n290 B.n289 585
R247 B.n288 B.n287 585
R248 B.n286 B.n285 585
R249 B.n284 B.n283 585
R250 B.n281 B.n280 585
R251 B.n279 B.n278 585
R252 B.n277 B.n276 585
R253 B.n275 B.n274 585
R254 B.n273 B.n272 585
R255 B.n271 B.n270 585
R256 B.n269 B.n268 585
R257 B.n267 B.n266 585
R258 B.n265 B.n264 585
R259 B.n263 B.n262 585
R260 B.n260 B.n259 585
R261 B.n258 B.n257 585
R262 B.n256 B.n255 585
R263 B.n254 B.n253 585
R264 B.n252 B.n251 585
R265 B.n250 B.n249 585
R266 B.n248 B.n247 585
R267 B.n246 B.n245 585
R268 B.n244 B.n243 585
R269 B.n242 B.n241 585
R270 B.n240 B.n239 585
R271 B.n238 B.n237 585
R272 B.n236 B.n235 585
R273 B.n234 B.n233 585
R274 B.n232 B.n231 585
R275 B.n230 B.n229 585
R276 B.n228 B.n227 585
R277 B.n226 B.n225 585
R278 B.n224 B.n223 585
R279 B.n222 B.n221 585
R280 B.n220 B.n219 585
R281 B.n218 B.n217 585
R282 B.n216 B.n215 585
R283 B.n214 B.n213 585
R284 B.n212 B.n211 585
R285 B.n210 B.n209 585
R286 B.n208 B.n207 585
R287 B.n206 B.n205 585
R288 B.n204 B.n203 585
R289 B.n202 B.n201 585
R290 B.n200 B.n199 585
R291 B.n198 B.n197 585
R292 B.n196 B.n195 585
R293 B.n194 B.n193 585
R294 B.n192 B.n191 585
R295 B.n190 B.n189 585
R296 B.n188 B.n187 585
R297 B.n186 B.n185 585
R298 B.n184 B.n183 585
R299 B.n182 B.n181 585
R300 B.n180 B.n179 585
R301 B.n178 B.n177 585
R302 B.n176 B.n175 585
R303 B.n174 B.n173 585
R304 B.n172 B.n171 585
R305 B.n170 B.n169 585
R306 B.n168 B.n167 585
R307 B.n166 B.n165 585
R308 B.n164 B.n163 585
R309 B.n1007 B.n104 585
R310 B.n1012 B.n104 585
R311 B.n1006 B.n103 585
R312 B.n1013 B.n103 585
R313 B.n1005 B.n1004 585
R314 B.n1004 B.n99 585
R315 B.n1003 B.n98 585
R316 B.n1019 B.n98 585
R317 B.n1002 B.n97 585
R318 B.n1020 B.n97 585
R319 B.n1001 B.n96 585
R320 B.n1021 B.n96 585
R321 B.n1000 B.n999 585
R322 B.n999 B.n92 585
R323 B.n998 B.n91 585
R324 B.n1027 B.n91 585
R325 B.n997 B.n90 585
R326 B.n1028 B.n90 585
R327 B.n996 B.n89 585
R328 B.n1029 B.n89 585
R329 B.n995 B.n994 585
R330 B.n994 B.n85 585
R331 B.n993 B.n84 585
R332 B.n1035 B.n84 585
R333 B.n992 B.n83 585
R334 B.n1036 B.n83 585
R335 B.n991 B.n82 585
R336 B.n1037 B.n82 585
R337 B.n990 B.n989 585
R338 B.n989 B.n78 585
R339 B.n988 B.n77 585
R340 B.n1043 B.n77 585
R341 B.n987 B.n76 585
R342 B.n1044 B.n76 585
R343 B.n986 B.n75 585
R344 B.n1045 B.n75 585
R345 B.n985 B.n984 585
R346 B.n984 B.n74 585
R347 B.n983 B.n70 585
R348 B.n1051 B.n70 585
R349 B.n982 B.n69 585
R350 B.n1052 B.n69 585
R351 B.n981 B.n68 585
R352 B.n1053 B.n68 585
R353 B.n980 B.n979 585
R354 B.n979 B.n64 585
R355 B.n978 B.n63 585
R356 B.n1059 B.n63 585
R357 B.n977 B.n62 585
R358 B.n1060 B.n62 585
R359 B.n976 B.n61 585
R360 B.n1061 B.n61 585
R361 B.n975 B.n974 585
R362 B.n974 B.n60 585
R363 B.n973 B.n56 585
R364 B.n1067 B.n56 585
R365 B.n972 B.n55 585
R366 B.n1068 B.n55 585
R367 B.n971 B.n54 585
R368 B.n1069 B.n54 585
R369 B.n970 B.n969 585
R370 B.n969 B.n50 585
R371 B.n968 B.n49 585
R372 B.n1075 B.n49 585
R373 B.n967 B.n48 585
R374 B.n1076 B.n48 585
R375 B.n966 B.n47 585
R376 B.n1077 B.n47 585
R377 B.n965 B.n964 585
R378 B.n964 B.n46 585
R379 B.n963 B.n42 585
R380 B.n1083 B.n42 585
R381 B.n962 B.n41 585
R382 B.n1084 B.n41 585
R383 B.n961 B.n40 585
R384 B.n1085 B.n40 585
R385 B.n960 B.n959 585
R386 B.n959 B.n36 585
R387 B.n958 B.n35 585
R388 B.n1091 B.n35 585
R389 B.n957 B.n34 585
R390 B.n1092 B.n34 585
R391 B.n956 B.n33 585
R392 B.n1093 B.n33 585
R393 B.n955 B.n954 585
R394 B.n954 B.n29 585
R395 B.n953 B.n28 585
R396 B.n1099 B.n28 585
R397 B.n952 B.n27 585
R398 B.n1100 B.n27 585
R399 B.n951 B.n26 585
R400 B.n1101 B.n26 585
R401 B.n950 B.n949 585
R402 B.n949 B.n22 585
R403 B.n948 B.n21 585
R404 B.n1107 B.n21 585
R405 B.n947 B.n20 585
R406 B.n1108 B.n20 585
R407 B.n946 B.n19 585
R408 B.n1109 B.n19 585
R409 B.n945 B.n944 585
R410 B.n944 B.n15 585
R411 B.n943 B.n14 585
R412 B.n1115 B.n14 585
R413 B.n942 B.n13 585
R414 B.n1116 B.n13 585
R415 B.n941 B.n12 585
R416 B.n1117 B.n12 585
R417 B.n940 B.n939 585
R418 B.n939 B.n8 585
R419 B.n938 B.n7 585
R420 B.n1123 B.n7 585
R421 B.n937 B.n6 585
R422 B.n1124 B.n6 585
R423 B.n936 B.n5 585
R424 B.n1125 B.n5 585
R425 B.n935 B.n934 585
R426 B.n934 B.n4 585
R427 B.n933 B.n378 585
R428 B.n933 B.n932 585
R429 B.n923 B.n379 585
R430 B.n380 B.n379 585
R431 B.n925 B.n924 585
R432 B.n926 B.n925 585
R433 B.n922 B.n385 585
R434 B.n385 B.n384 585
R435 B.n921 B.n920 585
R436 B.n920 B.n919 585
R437 B.n387 B.n386 585
R438 B.n388 B.n387 585
R439 B.n912 B.n911 585
R440 B.n913 B.n912 585
R441 B.n910 B.n393 585
R442 B.n393 B.n392 585
R443 B.n909 B.n908 585
R444 B.n908 B.n907 585
R445 B.n395 B.n394 585
R446 B.n396 B.n395 585
R447 B.n900 B.n899 585
R448 B.n901 B.n900 585
R449 B.n898 B.n401 585
R450 B.n401 B.n400 585
R451 B.n897 B.n896 585
R452 B.n896 B.n895 585
R453 B.n403 B.n402 585
R454 B.n404 B.n403 585
R455 B.n888 B.n887 585
R456 B.n889 B.n888 585
R457 B.n886 B.n409 585
R458 B.n409 B.n408 585
R459 B.n885 B.n884 585
R460 B.n884 B.n883 585
R461 B.n411 B.n410 585
R462 B.n412 B.n411 585
R463 B.n876 B.n875 585
R464 B.n877 B.n876 585
R465 B.n874 B.n417 585
R466 B.n417 B.n416 585
R467 B.n873 B.n872 585
R468 B.n872 B.n871 585
R469 B.n419 B.n418 585
R470 B.n864 B.n419 585
R471 B.n863 B.n862 585
R472 B.n865 B.n863 585
R473 B.n861 B.n424 585
R474 B.n424 B.n423 585
R475 B.n860 B.n859 585
R476 B.n859 B.n858 585
R477 B.n426 B.n425 585
R478 B.n427 B.n426 585
R479 B.n851 B.n850 585
R480 B.n852 B.n851 585
R481 B.n849 B.n432 585
R482 B.n432 B.n431 585
R483 B.n848 B.n847 585
R484 B.n847 B.n846 585
R485 B.n434 B.n433 585
R486 B.n839 B.n434 585
R487 B.n838 B.n837 585
R488 B.n840 B.n838 585
R489 B.n836 B.n439 585
R490 B.n439 B.n438 585
R491 B.n835 B.n834 585
R492 B.n834 B.n833 585
R493 B.n441 B.n440 585
R494 B.n442 B.n441 585
R495 B.n826 B.n825 585
R496 B.n827 B.n826 585
R497 B.n824 B.n447 585
R498 B.n447 B.n446 585
R499 B.n823 B.n822 585
R500 B.n822 B.n821 585
R501 B.n449 B.n448 585
R502 B.n814 B.n449 585
R503 B.n813 B.n812 585
R504 B.n815 B.n813 585
R505 B.n811 B.n454 585
R506 B.n454 B.n453 585
R507 B.n810 B.n809 585
R508 B.n809 B.n808 585
R509 B.n456 B.n455 585
R510 B.n457 B.n456 585
R511 B.n801 B.n800 585
R512 B.n802 B.n801 585
R513 B.n799 B.n462 585
R514 B.n462 B.n461 585
R515 B.n798 B.n797 585
R516 B.n797 B.n796 585
R517 B.n464 B.n463 585
R518 B.n465 B.n464 585
R519 B.n789 B.n788 585
R520 B.n790 B.n789 585
R521 B.n787 B.n470 585
R522 B.n470 B.n469 585
R523 B.n786 B.n785 585
R524 B.n785 B.n784 585
R525 B.n472 B.n471 585
R526 B.n473 B.n472 585
R527 B.n777 B.n776 585
R528 B.n778 B.n777 585
R529 B.n775 B.n478 585
R530 B.n478 B.n477 585
R531 B.n774 B.n773 585
R532 B.n773 B.n772 585
R533 B.n480 B.n479 585
R534 B.n481 B.n480 585
R535 B.n765 B.n764 585
R536 B.n766 B.n765 585
R537 B.n763 B.n486 585
R538 B.n486 B.n485 585
R539 B.n758 B.n757 585
R540 B.n756 B.n542 585
R541 B.n755 B.n541 585
R542 B.n760 B.n541 585
R543 B.n754 B.n753 585
R544 B.n752 B.n751 585
R545 B.n750 B.n749 585
R546 B.n748 B.n747 585
R547 B.n746 B.n745 585
R548 B.n744 B.n743 585
R549 B.n742 B.n741 585
R550 B.n740 B.n739 585
R551 B.n738 B.n737 585
R552 B.n736 B.n735 585
R553 B.n734 B.n733 585
R554 B.n732 B.n731 585
R555 B.n730 B.n729 585
R556 B.n728 B.n727 585
R557 B.n726 B.n725 585
R558 B.n724 B.n723 585
R559 B.n722 B.n721 585
R560 B.n720 B.n719 585
R561 B.n718 B.n717 585
R562 B.n716 B.n715 585
R563 B.n714 B.n713 585
R564 B.n712 B.n711 585
R565 B.n710 B.n709 585
R566 B.n708 B.n707 585
R567 B.n706 B.n705 585
R568 B.n704 B.n703 585
R569 B.n702 B.n701 585
R570 B.n700 B.n699 585
R571 B.n698 B.n697 585
R572 B.n696 B.n695 585
R573 B.n694 B.n693 585
R574 B.n692 B.n691 585
R575 B.n690 B.n689 585
R576 B.n688 B.n687 585
R577 B.n686 B.n685 585
R578 B.n684 B.n683 585
R579 B.n682 B.n681 585
R580 B.n680 B.n679 585
R581 B.n678 B.n677 585
R582 B.n676 B.n675 585
R583 B.n674 B.n673 585
R584 B.n672 B.n671 585
R585 B.n670 B.n669 585
R586 B.n668 B.n667 585
R587 B.n666 B.n665 585
R588 B.n664 B.n663 585
R589 B.n662 B.n661 585
R590 B.n660 B.n659 585
R591 B.n658 B.n657 585
R592 B.n656 B.n655 585
R593 B.n654 B.n653 585
R594 B.n652 B.n651 585
R595 B.n650 B.n649 585
R596 B.n648 B.n647 585
R597 B.n646 B.n645 585
R598 B.n644 B.n643 585
R599 B.n642 B.n641 585
R600 B.n640 B.n639 585
R601 B.n638 B.n637 585
R602 B.n636 B.n635 585
R603 B.n634 B.n633 585
R604 B.n632 B.n631 585
R605 B.n630 B.n629 585
R606 B.n628 B.n627 585
R607 B.n626 B.n625 585
R608 B.n624 B.n623 585
R609 B.n622 B.n621 585
R610 B.n620 B.n619 585
R611 B.n618 B.n617 585
R612 B.n616 B.n615 585
R613 B.n614 B.n613 585
R614 B.n612 B.n611 585
R615 B.n610 B.n609 585
R616 B.n608 B.n607 585
R617 B.n606 B.n605 585
R618 B.n604 B.n603 585
R619 B.n602 B.n601 585
R620 B.n600 B.n599 585
R621 B.n598 B.n597 585
R622 B.n596 B.n595 585
R623 B.n594 B.n593 585
R624 B.n592 B.n591 585
R625 B.n590 B.n589 585
R626 B.n588 B.n587 585
R627 B.n586 B.n585 585
R628 B.n584 B.n583 585
R629 B.n582 B.n581 585
R630 B.n580 B.n579 585
R631 B.n578 B.n577 585
R632 B.n576 B.n575 585
R633 B.n574 B.n573 585
R634 B.n572 B.n571 585
R635 B.n570 B.n569 585
R636 B.n568 B.n567 585
R637 B.n566 B.n565 585
R638 B.n564 B.n563 585
R639 B.n562 B.n561 585
R640 B.n560 B.n559 585
R641 B.n558 B.n557 585
R642 B.n556 B.n555 585
R643 B.n554 B.n553 585
R644 B.n552 B.n551 585
R645 B.n550 B.n549 585
R646 B.n488 B.n487 585
R647 B.n762 B.n761 585
R648 B.n761 B.n760 585
R649 B.n484 B.n483 585
R650 B.n485 B.n484 585
R651 B.n768 B.n767 585
R652 B.n767 B.n766 585
R653 B.n769 B.n482 585
R654 B.n482 B.n481 585
R655 B.n771 B.n770 585
R656 B.n772 B.n771 585
R657 B.n476 B.n475 585
R658 B.n477 B.n476 585
R659 B.n780 B.n779 585
R660 B.n779 B.n778 585
R661 B.n781 B.n474 585
R662 B.n474 B.n473 585
R663 B.n783 B.n782 585
R664 B.n784 B.n783 585
R665 B.n468 B.n467 585
R666 B.n469 B.n468 585
R667 B.n792 B.n791 585
R668 B.n791 B.n790 585
R669 B.n793 B.n466 585
R670 B.n466 B.n465 585
R671 B.n795 B.n794 585
R672 B.n796 B.n795 585
R673 B.n460 B.n459 585
R674 B.n461 B.n460 585
R675 B.n804 B.n803 585
R676 B.n803 B.n802 585
R677 B.n805 B.n458 585
R678 B.n458 B.n457 585
R679 B.n807 B.n806 585
R680 B.n808 B.n807 585
R681 B.n452 B.n451 585
R682 B.n453 B.n452 585
R683 B.n817 B.n816 585
R684 B.n816 B.n815 585
R685 B.n818 B.n450 585
R686 B.n814 B.n450 585
R687 B.n820 B.n819 585
R688 B.n821 B.n820 585
R689 B.n445 B.n444 585
R690 B.n446 B.n445 585
R691 B.n829 B.n828 585
R692 B.n828 B.n827 585
R693 B.n830 B.n443 585
R694 B.n443 B.n442 585
R695 B.n832 B.n831 585
R696 B.n833 B.n832 585
R697 B.n437 B.n436 585
R698 B.n438 B.n437 585
R699 B.n842 B.n841 585
R700 B.n841 B.n840 585
R701 B.n843 B.n435 585
R702 B.n839 B.n435 585
R703 B.n845 B.n844 585
R704 B.n846 B.n845 585
R705 B.n430 B.n429 585
R706 B.n431 B.n430 585
R707 B.n854 B.n853 585
R708 B.n853 B.n852 585
R709 B.n855 B.n428 585
R710 B.n428 B.n427 585
R711 B.n857 B.n856 585
R712 B.n858 B.n857 585
R713 B.n422 B.n421 585
R714 B.n423 B.n422 585
R715 B.n867 B.n866 585
R716 B.n866 B.n865 585
R717 B.n868 B.n420 585
R718 B.n864 B.n420 585
R719 B.n870 B.n869 585
R720 B.n871 B.n870 585
R721 B.n415 B.n414 585
R722 B.n416 B.n415 585
R723 B.n879 B.n878 585
R724 B.n878 B.n877 585
R725 B.n880 B.n413 585
R726 B.n413 B.n412 585
R727 B.n882 B.n881 585
R728 B.n883 B.n882 585
R729 B.n407 B.n406 585
R730 B.n408 B.n407 585
R731 B.n891 B.n890 585
R732 B.n890 B.n889 585
R733 B.n892 B.n405 585
R734 B.n405 B.n404 585
R735 B.n894 B.n893 585
R736 B.n895 B.n894 585
R737 B.n399 B.n398 585
R738 B.n400 B.n399 585
R739 B.n903 B.n902 585
R740 B.n902 B.n901 585
R741 B.n904 B.n397 585
R742 B.n397 B.n396 585
R743 B.n906 B.n905 585
R744 B.n907 B.n906 585
R745 B.n391 B.n390 585
R746 B.n392 B.n391 585
R747 B.n915 B.n914 585
R748 B.n914 B.n913 585
R749 B.n916 B.n389 585
R750 B.n389 B.n388 585
R751 B.n918 B.n917 585
R752 B.n919 B.n918 585
R753 B.n383 B.n382 585
R754 B.n384 B.n383 585
R755 B.n928 B.n927 585
R756 B.n927 B.n926 585
R757 B.n929 B.n381 585
R758 B.n381 B.n380 585
R759 B.n931 B.n930 585
R760 B.n932 B.n931 585
R761 B.n2 B.n0 585
R762 B.n4 B.n2 585
R763 B.n3 B.n1 585
R764 B.n1124 B.n3 585
R765 B.n1122 B.n1121 585
R766 B.n1123 B.n1122 585
R767 B.n1120 B.n9 585
R768 B.n9 B.n8 585
R769 B.n1119 B.n1118 585
R770 B.n1118 B.n1117 585
R771 B.n11 B.n10 585
R772 B.n1116 B.n11 585
R773 B.n1114 B.n1113 585
R774 B.n1115 B.n1114 585
R775 B.n1112 B.n16 585
R776 B.n16 B.n15 585
R777 B.n1111 B.n1110 585
R778 B.n1110 B.n1109 585
R779 B.n18 B.n17 585
R780 B.n1108 B.n18 585
R781 B.n1106 B.n1105 585
R782 B.n1107 B.n1106 585
R783 B.n1104 B.n23 585
R784 B.n23 B.n22 585
R785 B.n1103 B.n1102 585
R786 B.n1102 B.n1101 585
R787 B.n25 B.n24 585
R788 B.n1100 B.n25 585
R789 B.n1098 B.n1097 585
R790 B.n1099 B.n1098 585
R791 B.n1096 B.n30 585
R792 B.n30 B.n29 585
R793 B.n1095 B.n1094 585
R794 B.n1094 B.n1093 585
R795 B.n32 B.n31 585
R796 B.n1092 B.n32 585
R797 B.n1090 B.n1089 585
R798 B.n1091 B.n1090 585
R799 B.n1088 B.n37 585
R800 B.n37 B.n36 585
R801 B.n1087 B.n1086 585
R802 B.n1086 B.n1085 585
R803 B.n39 B.n38 585
R804 B.n1084 B.n39 585
R805 B.n1082 B.n1081 585
R806 B.n1083 B.n1082 585
R807 B.n1080 B.n43 585
R808 B.n46 B.n43 585
R809 B.n1079 B.n1078 585
R810 B.n1078 B.n1077 585
R811 B.n45 B.n44 585
R812 B.n1076 B.n45 585
R813 B.n1074 B.n1073 585
R814 B.n1075 B.n1074 585
R815 B.n1072 B.n51 585
R816 B.n51 B.n50 585
R817 B.n1071 B.n1070 585
R818 B.n1070 B.n1069 585
R819 B.n53 B.n52 585
R820 B.n1068 B.n53 585
R821 B.n1066 B.n1065 585
R822 B.n1067 B.n1066 585
R823 B.n1064 B.n57 585
R824 B.n60 B.n57 585
R825 B.n1063 B.n1062 585
R826 B.n1062 B.n1061 585
R827 B.n59 B.n58 585
R828 B.n1060 B.n59 585
R829 B.n1058 B.n1057 585
R830 B.n1059 B.n1058 585
R831 B.n1056 B.n65 585
R832 B.n65 B.n64 585
R833 B.n1055 B.n1054 585
R834 B.n1054 B.n1053 585
R835 B.n67 B.n66 585
R836 B.n1052 B.n67 585
R837 B.n1050 B.n1049 585
R838 B.n1051 B.n1050 585
R839 B.n1048 B.n71 585
R840 B.n74 B.n71 585
R841 B.n1047 B.n1046 585
R842 B.n1046 B.n1045 585
R843 B.n73 B.n72 585
R844 B.n1044 B.n73 585
R845 B.n1042 B.n1041 585
R846 B.n1043 B.n1042 585
R847 B.n1040 B.n79 585
R848 B.n79 B.n78 585
R849 B.n1039 B.n1038 585
R850 B.n1038 B.n1037 585
R851 B.n81 B.n80 585
R852 B.n1036 B.n81 585
R853 B.n1034 B.n1033 585
R854 B.n1035 B.n1034 585
R855 B.n1032 B.n86 585
R856 B.n86 B.n85 585
R857 B.n1031 B.n1030 585
R858 B.n1030 B.n1029 585
R859 B.n88 B.n87 585
R860 B.n1028 B.n88 585
R861 B.n1026 B.n1025 585
R862 B.n1027 B.n1026 585
R863 B.n1024 B.n93 585
R864 B.n93 B.n92 585
R865 B.n1023 B.n1022 585
R866 B.n1022 B.n1021 585
R867 B.n95 B.n94 585
R868 B.n1020 B.n95 585
R869 B.n1018 B.n1017 585
R870 B.n1019 B.n1018 585
R871 B.n1016 B.n100 585
R872 B.n100 B.n99 585
R873 B.n1015 B.n1014 585
R874 B.n1014 B.n1013 585
R875 B.n102 B.n101 585
R876 B.n1012 B.n102 585
R877 B.n1127 B.n1126 585
R878 B.n1126 B.n1125 585
R879 B.n758 B.n484 535.745
R880 B.n163 B.n102 535.745
R881 B.n761 B.n486 535.745
R882 B.n1009 B.n104 535.745
R883 B.n546 B.t10 351.425
R884 B.n543 B.t14 351.425
R885 B.n161 B.t21 351.425
R886 B.n159 B.t17 351.425
R887 B.n1011 B.n1010 256.663
R888 B.n1011 B.n157 256.663
R889 B.n1011 B.n156 256.663
R890 B.n1011 B.n155 256.663
R891 B.n1011 B.n154 256.663
R892 B.n1011 B.n153 256.663
R893 B.n1011 B.n152 256.663
R894 B.n1011 B.n151 256.663
R895 B.n1011 B.n150 256.663
R896 B.n1011 B.n149 256.663
R897 B.n1011 B.n148 256.663
R898 B.n1011 B.n147 256.663
R899 B.n1011 B.n146 256.663
R900 B.n1011 B.n145 256.663
R901 B.n1011 B.n144 256.663
R902 B.n1011 B.n143 256.663
R903 B.n1011 B.n142 256.663
R904 B.n1011 B.n141 256.663
R905 B.n1011 B.n140 256.663
R906 B.n1011 B.n139 256.663
R907 B.n1011 B.n138 256.663
R908 B.n1011 B.n137 256.663
R909 B.n1011 B.n136 256.663
R910 B.n1011 B.n135 256.663
R911 B.n1011 B.n134 256.663
R912 B.n1011 B.n133 256.663
R913 B.n1011 B.n132 256.663
R914 B.n1011 B.n131 256.663
R915 B.n1011 B.n130 256.663
R916 B.n1011 B.n129 256.663
R917 B.n1011 B.n128 256.663
R918 B.n1011 B.n127 256.663
R919 B.n1011 B.n126 256.663
R920 B.n1011 B.n125 256.663
R921 B.n1011 B.n124 256.663
R922 B.n1011 B.n123 256.663
R923 B.n1011 B.n122 256.663
R924 B.n1011 B.n121 256.663
R925 B.n1011 B.n120 256.663
R926 B.n1011 B.n119 256.663
R927 B.n1011 B.n118 256.663
R928 B.n1011 B.n117 256.663
R929 B.n1011 B.n116 256.663
R930 B.n1011 B.n115 256.663
R931 B.n1011 B.n114 256.663
R932 B.n1011 B.n113 256.663
R933 B.n1011 B.n112 256.663
R934 B.n1011 B.n111 256.663
R935 B.n1011 B.n110 256.663
R936 B.n1011 B.n109 256.663
R937 B.n1011 B.n108 256.663
R938 B.n1011 B.n107 256.663
R939 B.n1011 B.n106 256.663
R940 B.n1011 B.n105 256.663
R941 B.n760 B.n759 256.663
R942 B.n760 B.n489 256.663
R943 B.n760 B.n490 256.663
R944 B.n760 B.n491 256.663
R945 B.n760 B.n492 256.663
R946 B.n760 B.n493 256.663
R947 B.n760 B.n494 256.663
R948 B.n760 B.n495 256.663
R949 B.n760 B.n496 256.663
R950 B.n760 B.n497 256.663
R951 B.n760 B.n498 256.663
R952 B.n760 B.n499 256.663
R953 B.n760 B.n500 256.663
R954 B.n760 B.n501 256.663
R955 B.n760 B.n502 256.663
R956 B.n760 B.n503 256.663
R957 B.n760 B.n504 256.663
R958 B.n760 B.n505 256.663
R959 B.n760 B.n506 256.663
R960 B.n760 B.n507 256.663
R961 B.n760 B.n508 256.663
R962 B.n760 B.n509 256.663
R963 B.n760 B.n510 256.663
R964 B.n760 B.n511 256.663
R965 B.n760 B.n512 256.663
R966 B.n760 B.n513 256.663
R967 B.n760 B.n514 256.663
R968 B.n760 B.n515 256.663
R969 B.n760 B.n516 256.663
R970 B.n760 B.n517 256.663
R971 B.n760 B.n518 256.663
R972 B.n760 B.n519 256.663
R973 B.n760 B.n520 256.663
R974 B.n760 B.n521 256.663
R975 B.n760 B.n522 256.663
R976 B.n760 B.n523 256.663
R977 B.n760 B.n524 256.663
R978 B.n760 B.n525 256.663
R979 B.n760 B.n526 256.663
R980 B.n760 B.n527 256.663
R981 B.n760 B.n528 256.663
R982 B.n760 B.n529 256.663
R983 B.n760 B.n530 256.663
R984 B.n760 B.n531 256.663
R985 B.n760 B.n532 256.663
R986 B.n760 B.n533 256.663
R987 B.n760 B.n534 256.663
R988 B.n760 B.n535 256.663
R989 B.n760 B.n536 256.663
R990 B.n760 B.n537 256.663
R991 B.n760 B.n538 256.663
R992 B.n760 B.n539 256.663
R993 B.n760 B.n540 256.663
R994 B.n767 B.n484 163.367
R995 B.n767 B.n482 163.367
R996 B.n771 B.n482 163.367
R997 B.n771 B.n476 163.367
R998 B.n779 B.n476 163.367
R999 B.n779 B.n474 163.367
R1000 B.n783 B.n474 163.367
R1001 B.n783 B.n468 163.367
R1002 B.n791 B.n468 163.367
R1003 B.n791 B.n466 163.367
R1004 B.n795 B.n466 163.367
R1005 B.n795 B.n460 163.367
R1006 B.n803 B.n460 163.367
R1007 B.n803 B.n458 163.367
R1008 B.n807 B.n458 163.367
R1009 B.n807 B.n452 163.367
R1010 B.n816 B.n452 163.367
R1011 B.n816 B.n450 163.367
R1012 B.n820 B.n450 163.367
R1013 B.n820 B.n445 163.367
R1014 B.n828 B.n445 163.367
R1015 B.n828 B.n443 163.367
R1016 B.n832 B.n443 163.367
R1017 B.n832 B.n437 163.367
R1018 B.n841 B.n437 163.367
R1019 B.n841 B.n435 163.367
R1020 B.n845 B.n435 163.367
R1021 B.n845 B.n430 163.367
R1022 B.n853 B.n430 163.367
R1023 B.n853 B.n428 163.367
R1024 B.n857 B.n428 163.367
R1025 B.n857 B.n422 163.367
R1026 B.n866 B.n422 163.367
R1027 B.n866 B.n420 163.367
R1028 B.n870 B.n420 163.367
R1029 B.n870 B.n415 163.367
R1030 B.n878 B.n415 163.367
R1031 B.n878 B.n413 163.367
R1032 B.n882 B.n413 163.367
R1033 B.n882 B.n407 163.367
R1034 B.n890 B.n407 163.367
R1035 B.n890 B.n405 163.367
R1036 B.n894 B.n405 163.367
R1037 B.n894 B.n399 163.367
R1038 B.n902 B.n399 163.367
R1039 B.n902 B.n397 163.367
R1040 B.n906 B.n397 163.367
R1041 B.n906 B.n391 163.367
R1042 B.n914 B.n391 163.367
R1043 B.n914 B.n389 163.367
R1044 B.n918 B.n389 163.367
R1045 B.n918 B.n383 163.367
R1046 B.n927 B.n383 163.367
R1047 B.n927 B.n381 163.367
R1048 B.n931 B.n381 163.367
R1049 B.n931 B.n2 163.367
R1050 B.n1126 B.n2 163.367
R1051 B.n1126 B.n3 163.367
R1052 B.n1122 B.n3 163.367
R1053 B.n1122 B.n9 163.367
R1054 B.n1118 B.n9 163.367
R1055 B.n1118 B.n11 163.367
R1056 B.n1114 B.n11 163.367
R1057 B.n1114 B.n16 163.367
R1058 B.n1110 B.n16 163.367
R1059 B.n1110 B.n18 163.367
R1060 B.n1106 B.n18 163.367
R1061 B.n1106 B.n23 163.367
R1062 B.n1102 B.n23 163.367
R1063 B.n1102 B.n25 163.367
R1064 B.n1098 B.n25 163.367
R1065 B.n1098 B.n30 163.367
R1066 B.n1094 B.n30 163.367
R1067 B.n1094 B.n32 163.367
R1068 B.n1090 B.n32 163.367
R1069 B.n1090 B.n37 163.367
R1070 B.n1086 B.n37 163.367
R1071 B.n1086 B.n39 163.367
R1072 B.n1082 B.n39 163.367
R1073 B.n1082 B.n43 163.367
R1074 B.n1078 B.n43 163.367
R1075 B.n1078 B.n45 163.367
R1076 B.n1074 B.n45 163.367
R1077 B.n1074 B.n51 163.367
R1078 B.n1070 B.n51 163.367
R1079 B.n1070 B.n53 163.367
R1080 B.n1066 B.n53 163.367
R1081 B.n1066 B.n57 163.367
R1082 B.n1062 B.n57 163.367
R1083 B.n1062 B.n59 163.367
R1084 B.n1058 B.n59 163.367
R1085 B.n1058 B.n65 163.367
R1086 B.n1054 B.n65 163.367
R1087 B.n1054 B.n67 163.367
R1088 B.n1050 B.n67 163.367
R1089 B.n1050 B.n71 163.367
R1090 B.n1046 B.n71 163.367
R1091 B.n1046 B.n73 163.367
R1092 B.n1042 B.n73 163.367
R1093 B.n1042 B.n79 163.367
R1094 B.n1038 B.n79 163.367
R1095 B.n1038 B.n81 163.367
R1096 B.n1034 B.n81 163.367
R1097 B.n1034 B.n86 163.367
R1098 B.n1030 B.n86 163.367
R1099 B.n1030 B.n88 163.367
R1100 B.n1026 B.n88 163.367
R1101 B.n1026 B.n93 163.367
R1102 B.n1022 B.n93 163.367
R1103 B.n1022 B.n95 163.367
R1104 B.n1018 B.n95 163.367
R1105 B.n1018 B.n100 163.367
R1106 B.n1014 B.n100 163.367
R1107 B.n1014 B.n102 163.367
R1108 B.n542 B.n541 163.367
R1109 B.n753 B.n541 163.367
R1110 B.n751 B.n750 163.367
R1111 B.n747 B.n746 163.367
R1112 B.n743 B.n742 163.367
R1113 B.n739 B.n738 163.367
R1114 B.n735 B.n734 163.367
R1115 B.n731 B.n730 163.367
R1116 B.n727 B.n726 163.367
R1117 B.n723 B.n722 163.367
R1118 B.n719 B.n718 163.367
R1119 B.n715 B.n714 163.367
R1120 B.n711 B.n710 163.367
R1121 B.n707 B.n706 163.367
R1122 B.n703 B.n702 163.367
R1123 B.n699 B.n698 163.367
R1124 B.n695 B.n694 163.367
R1125 B.n691 B.n690 163.367
R1126 B.n687 B.n686 163.367
R1127 B.n683 B.n682 163.367
R1128 B.n679 B.n678 163.367
R1129 B.n675 B.n674 163.367
R1130 B.n671 B.n670 163.367
R1131 B.n667 B.n666 163.367
R1132 B.n663 B.n662 163.367
R1133 B.n659 B.n658 163.367
R1134 B.n655 B.n654 163.367
R1135 B.n651 B.n650 163.367
R1136 B.n647 B.n646 163.367
R1137 B.n643 B.n642 163.367
R1138 B.n639 B.n638 163.367
R1139 B.n635 B.n634 163.367
R1140 B.n631 B.n630 163.367
R1141 B.n627 B.n626 163.367
R1142 B.n623 B.n622 163.367
R1143 B.n619 B.n618 163.367
R1144 B.n615 B.n614 163.367
R1145 B.n611 B.n610 163.367
R1146 B.n607 B.n606 163.367
R1147 B.n603 B.n602 163.367
R1148 B.n599 B.n598 163.367
R1149 B.n595 B.n594 163.367
R1150 B.n591 B.n590 163.367
R1151 B.n587 B.n586 163.367
R1152 B.n583 B.n582 163.367
R1153 B.n579 B.n578 163.367
R1154 B.n575 B.n574 163.367
R1155 B.n571 B.n570 163.367
R1156 B.n567 B.n566 163.367
R1157 B.n563 B.n562 163.367
R1158 B.n559 B.n558 163.367
R1159 B.n555 B.n554 163.367
R1160 B.n551 B.n550 163.367
R1161 B.n761 B.n488 163.367
R1162 B.n765 B.n486 163.367
R1163 B.n765 B.n480 163.367
R1164 B.n773 B.n480 163.367
R1165 B.n773 B.n478 163.367
R1166 B.n777 B.n478 163.367
R1167 B.n777 B.n472 163.367
R1168 B.n785 B.n472 163.367
R1169 B.n785 B.n470 163.367
R1170 B.n789 B.n470 163.367
R1171 B.n789 B.n464 163.367
R1172 B.n797 B.n464 163.367
R1173 B.n797 B.n462 163.367
R1174 B.n801 B.n462 163.367
R1175 B.n801 B.n456 163.367
R1176 B.n809 B.n456 163.367
R1177 B.n809 B.n454 163.367
R1178 B.n813 B.n454 163.367
R1179 B.n813 B.n449 163.367
R1180 B.n822 B.n449 163.367
R1181 B.n822 B.n447 163.367
R1182 B.n826 B.n447 163.367
R1183 B.n826 B.n441 163.367
R1184 B.n834 B.n441 163.367
R1185 B.n834 B.n439 163.367
R1186 B.n838 B.n439 163.367
R1187 B.n838 B.n434 163.367
R1188 B.n847 B.n434 163.367
R1189 B.n847 B.n432 163.367
R1190 B.n851 B.n432 163.367
R1191 B.n851 B.n426 163.367
R1192 B.n859 B.n426 163.367
R1193 B.n859 B.n424 163.367
R1194 B.n863 B.n424 163.367
R1195 B.n863 B.n419 163.367
R1196 B.n872 B.n419 163.367
R1197 B.n872 B.n417 163.367
R1198 B.n876 B.n417 163.367
R1199 B.n876 B.n411 163.367
R1200 B.n884 B.n411 163.367
R1201 B.n884 B.n409 163.367
R1202 B.n888 B.n409 163.367
R1203 B.n888 B.n403 163.367
R1204 B.n896 B.n403 163.367
R1205 B.n896 B.n401 163.367
R1206 B.n900 B.n401 163.367
R1207 B.n900 B.n395 163.367
R1208 B.n908 B.n395 163.367
R1209 B.n908 B.n393 163.367
R1210 B.n912 B.n393 163.367
R1211 B.n912 B.n387 163.367
R1212 B.n920 B.n387 163.367
R1213 B.n920 B.n385 163.367
R1214 B.n925 B.n385 163.367
R1215 B.n925 B.n379 163.367
R1216 B.n933 B.n379 163.367
R1217 B.n934 B.n933 163.367
R1218 B.n934 B.n5 163.367
R1219 B.n6 B.n5 163.367
R1220 B.n7 B.n6 163.367
R1221 B.n939 B.n7 163.367
R1222 B.n939 B.n12 163.367
R1223 B.n13 B.n12 163.367
R1224 B.n14 B.n13 163.367
R1225 B.n944 B.n14 163.367
R1226 B.n944 B.n19 163.367
R1227 B.n20 B.n19 163.367
R1228 B.n21 B.n20 163.367
R1229 B.n949 B.n21 163.367
R1230 B.n949 B.n26 163.367
R1231 B.n27 B.n26 163.367
R1232 B.n28 B.n27 163.367
R1233 B.n954 B.n28 163.367
R1234 B.n954 B.n33 163.367
R1235 B.n34 B.n33 163.367
R1236 B.n35 B.n34 163.367
R1237 B.n959 B.n35 163.367
R1238 B.n959 B.n40 163.367
R1239 B.n41 B.n40 163.367
R1240 B.n42 B.n41 163.367
R1241 B.n964 B.n42 163.367
R1242 B.n964 B.n47 163.367
R1243 B.n48 B.n47 163.367
R1244 B.n49 B.n48 163.367
R1245 B.n969 B.n49 163.367
R1246 B.n969 B.n54 163.367
R1247 B.n55 B.n54 163.367
R1248 B.n56 B.n55 163.367
R1249 B.n974 B.n56 163.367
R1250 B.n974 B.n61 163.367
R1251 B.n62 B.n61 163.367
R1252 B.n63 B.n62 163.367
R1253 B.n979 B.n63 163.367
R1254 B.n979 B.n68 163.367
R1255 B.n69 B.n68 163.367
R1256 B.n70 B.n69 163.367
R1257 B.n984 B.n70 163.367
R1258 B.n984 B.n75 163.367
R1259 B.n76 B.n75 163.367
R1260 B.n77 B.n76 163.367
R1261 B.n989 B.n77 163.367
R1262 B.n989 B.n82 163.367
R1263 B.n83 B.n82 163.367
R1264 B.n84 B.n83 163.367
R1265 B.n994 B.n84 163.367
R1266 B.n994 B.n89 163.367
R1267 B.n90 B.n89 163.367
R1268 B.n91 B.n90 163.367
R1269 B.n999 B.n91 163.367
R1270 B.n999 B.n96 163.367
R1271 B.n97 B.n96 163.367
R1272 B.n98 B.n97 163.367
R1273 B.n1004 B.n98 163.367
R1274 B.n1004 B.n103 163.367
R1275 B.n104 B.n103 163.367
R1276 B.n167 B.n166 163.367
R1277 B.n171 B.n170 163.367
R1278 B.n175 B.n174 163.367
R1279 B.n179 B.n178 163.367
R1280 B.n183 B.n182 163.367
R1281 B.n187 B.n186 163.367
R1282 B.n191 B.n190 163.367
R1283 B.n195 B.n194 163.367
R1284 B.n199 B.n198 163.367
R1285 B.n203 B.n202 163.367
R1286 B.n207 B.n206 163.367
R1287 B.n211 B.n210 163.367
R1288 B.n215 B.n214 163.367
R1289 B.n219 B.n218 163.367
R1290 B.n223 B.n222 163.367
R1291 B.n227 B.n226 163.367
R1292 B.n231 B.n230 163.367
R1293 B.n235 B.n234 163.367
R1294 B.n239 B.n238 163.367
R1295 B.n243 B.n242 163.367
R1296 B.n247 B.n246 163.367
R1297 B.n251 B.n250 163.367
R1298 B.n255 B.n254 163.367
R1299 B.n259 B.n258 163.367
R1300 B.n264 B.n263 163.367
R1301 B.n268 B.n267 163.367
R1302 B.n272 B.n271 163.367
R1303 B.n276 B.n275 163.367
R1304 B.n280 B.n279 163.367
R1305 B.n285 B.n284 163.367
R1306 B.n289 B.n288 163.367
R1307 B.n293 B.n292 163.367
R1308 B.n297 B.n296 163.367
R1309 B.n301 B.n300 163.367
R1310 B.n305 B.n304 163.367
R1311 B.n309 B.n308 163.367
R1312 B.n313 B.n312 163.367
R1313 B.n317 B.n316 163.367
R1314 B.n321 B.n320 163.367
R1315 B.n325 B.n324 163.367
R1316 B.n329 B.n328 163.367
R1317 B.n333 B.n332 163.367
R1318 B.n337 B.n336 163.367
R1319 B.n341 B.n340 163.367
R1320 B.n345 B.n344 163.367
R1321 B.n349 B.n348 163.367
R1322 B.n353 B.n352 163.367
R1323 B.n357 B.n356 163.367
R1324 B.n361 B.n360 163.367
R1325 B.n365 B.n364 163.367
R1326 B.n369 B.n368 163.367
R1327 B.n373 B.n372 163.367
R1328 B.n375 B.n158 163.367
R1329 B.n546 B.t13 127.621
R1330 B.n159 B.t19 127.621
R1331 B.n543 B.t16 127.603
R1332 B.n161 B.t22 127.603
R1333 B.n760 B.n485 74.7175
R1334 B.n1012 B.n1011 74.7175
R1335 B.n547 B.t12 73.7056
R1336 B.n160 B.t20 73.7056
R1337 B.n544 B.t15 73.6869
R1338 B.n162 B.t23 73.6869
R1339 B.n759 B.n758 71.676
R1340 B.n753 B.n489 71.676
R1341 B.n750 B.n490 71.676
R1342 B.n746 B.n491 71.676
R1343 B.n742 B.n492 71.676
R1344 B.n738 B.n493 71.676
R1345 B.n734 B.n494 71.676
R1346 B.n730 B.n495 71.676
R1347 B.n726 B.n496 71.676
R1348 B.n722 B.n497 71.676
R1349 B.n718 B.n498 71.676
R1350 B.n714 B.n499 71.676
R1351 B.n710 B.n500 71.676
R1352 B.n706 B.n501 71.676
R1353 B.n702 B.n502 71.676
R1354 B.n698 B.n503 71.676
R1355 B.n694 B.n504 71.676
R1356 B.n690 B.n505 71.676
R1357 B.n686 B.n506 71.676
R1358 B.n682 B.n507 71.676
R1359 B.n678 B.n508 71.676
R1360 B.n674 B.n509 71.676
R1361 B.n670 B.n510 71.676
R1362 B.n666 B.n511 71.676
R1363 B.n662 B.n512 71.676
R1364 B.n658 B.n513 71.676
R1365 B.n654 B.n514 71.676
R1366 B.n650 B.n515 71.676
R1367 B.n646 B.n516 71.676
R1368 B.n642 B.n517 71.676
R1369 B.n638 B.n518 71.676
R1370 B.n634 B.n519 71.676
R1371 B.n630 B.n520 71.676
R1372 B.n626 B.n521 71.676
R1373 B.n622 B.n522 71.676
R1374 B.n618 B.n523 71.676
R1375 B.n614 B.n524 71.676
R1376 B.n610 B.n525 71.676
R1377 B.n606 B.n526 71.676
R1378 B.n602 B.n527 71.676
R1379 B.n598 B.n528 71.676
R1380 B.n594 B.n529 71.676
R1381 B.n590 B.n530 71.676
R1382 B.n586 B.n531 71.676
R1383 B.n582 B.n532 71.676
R1384 B.n578 B.n533 71.676
R1385 B.n574 B.n534 71.676
R1386 B.n570 B.n535 71.676
R1387 B.n566 B.n536 71.676
R1388 B.n562 B.n537 71.676
R1389 B.n558 B.n538 71.676
R1390 B.n554 B.n539 71.676
R1391 B.n550 B.n540 71.676
R1392 B.n163 B.n105 71.676
R1393 B.n167 B.n106 71.676
R1394 B.n171 B.n107 71.676
R1395 B.n175 B.n108 71.676
R1396 B.n179 B.n109 71.676
R1397 B.n183 B.n110 71.676
R1398 B.n187 B.n111 71.676
R1399 B.n191 B.n112 71.676
R1400 B.n195 B.n113 71.676
R1401 B.n199 B.n114 71.676
R1402 B.n203 B.n115 71.676
R1403 B.n207 B.n116 71.676
R1404 B.n211 B.n117 71.676
R1405 B.n215 B.n118 71.676
R1406 B.n219 B.n119 71.676
R1407 B.n223 B.n120 71.676
R1408 B.n227 B.n121 71.676
R1409 B.n231 B.n122 71.676
R1410 B.n235 B.n123 71.676
R1411 B.n239 B.n124 71.676
R1412 B.n243 B.n125 71.676
R1413 B.n247 B.n126 71.676
R1414 B.n251 B.n127 71.676
R1415 B.n255 B.n128 71.676
R1416 B.n259 B.n129 71.676
R1417 B.n264 B.n130 71.676
R1418 B.n268 B.n131 71.676
R1419 B.n272 B.n132 71.676
R1420 B.n276 B.n133 71.676
R1421 B.n280 B.n134 71.676
R1422 B.n285 B.n135 71.676
R1423 B.n289 B.n136 71.676
R1424 B.n293 B.n137 71.676
R1425 B.n297 B.n138 71.676
R1426 B.n301 B.n139 71.676
R1427 B.n305 B.n140 71.676
R1428 B.n309 B.n141 71.676
R1429 B.n313 B.n142 71.676
R1430 B.n317 B.n143 71.676
R1431 B.n321 B.n144 71.676
R1432 B.n325 B.n145 71.676
R1433 B.n329 B.n146 71.676
R1434 B.n333 B.n147 71.676
R1435 B.n337 B.n148 71.676
R1436 B.n341 B.n149 71.676
R1437 B.n345 B.n150 71.676
R1438 B.n349 B.n151 71.676
R1439 B.n353 B.n152 71.676
R1440 B.n357 B.n153 71.676
R1441 B.n361 B.n154 71.676
R1442 B.n365 B.n155 71.676
R1443 B.n369 B.n156 71.676
R1444 B.n373 B.n157 71.676
R1445 B.n1010 B.n158 71.676
R1446 B.n1010 B.n1009 71.676
R1447 B.n375 B.n157 71.676
R1448 B.n372 B.n156 71.676
R1449 B.n368 B.n155 71.676
R1450 B.n364 B.n154 71.676
R1451 B.n360 B.n153 71.676
R1452 B.n356 B.n152 71.676
R1453 B.n352 B.n151 71.676
R1454 B.n348 B.n150 71.676
R1455 B.n344 B.n149 71.676
R1456 B.n340 B.n148 71.676
R1457 B.n336 B.n147 71.676
R1458 B.n332 B.n146 71.676
R1459 B.n328 B.n145 71.676
R1460 B.n324 B.n144 71.676
R1461 B.n320 B.n143 71.676
R1462 B.n316 B.n142 71.676
R1463 B.n312 B.n141 71.676
R1464 B.n308 B.n140 71.676
R1465 B.n304 B.n139 71.676
R1466 B.n300 B.n138 71.676
R1467 B.n296 B.n137 71.676
R1468 B.n292 B.n136 71.676
R1469 B.n288 B.n135 71.676
R1470 B.n284 B.n134 71.676
R1471 B.n279 B.n133 71.676
R1472 B.n275 B.n132 71.676
R1473 B.n271 B.n131 71.676
R1474 B.n267 B.n130 71.676
R1475 B.n263 B.n129 71.676
R1476 B.n258 B.n128 71.676
R1477 B.n254 B.n127 71.676
R1478 B.n250 B.n126 71.676
R1479 B.n246 B.n125 71.676
R1480 B.n242 B.n124 71.676
R1481 B.n238 B.n123 71.676
R1482 B.n234 B.n122 71.676
R1483 B.n230 B.n121 71.676
R1484 B.n226 B.n120 71.676
R1485 B.n222 B.n119 71.676
R1486 B.n218 B.n118 71.676
R1487 B.n214 B.n117 71.676
R1488 B.n210 B.n116 71.676
R1489 B.n206 B.n115 71.676
R1490 B.n202 B.n114 71.676
R1491 B.n198 B.n113 71.676
R1492 B.n194 B.n112 71.676
R1493 B.n190 B.n111 71.676
R1494 B.n186 B.n110 71.676
R1495 B.n182 B.n109 71.676
R1496 B.n178 B.n108 71.676
R1497 B.n174 B.n107 71.676
R1498 B.n170 B.n106 71.676
R1499 B.n166 B.n105 71.676
R1500 B.n759 B.n542 71.676
R1501 B.n751 B.n489 71.676
R1502 B.n747 B.n490 71.676
R1503 B.n743 B.n491 71.676
R1504 B.n739 B.n492 71.676
R1505 B.n735 B.n493 71.676
R1506 B.n731 B.n494 71.676
R1507 B.n727 B.n495 71.676
R1508 B.n723 B.n496 71.676
R1509 B.n719 B.n497 71.676
R1510 B.n715 B.n498 71.676
R1511 B.n711 B.n499 71.676
R1512 B.n707 B.n500 71.676
R1513 B.n703 B.n501 71.676
R1514 B.n699 B.n502 71.676
R1515 B.n695 B.n503 71.676
R1516 B.n691 B.n504 71.676
R1517 B.n687 B.n505 71.676
R1518 B.n683 B.n506 71.676
R1519 B.n679 B.n507 71.676
R1520 B.n675 B.n508 71.676
R1521 B.n671 B.n509 71.676
R1522 B.n667 B.n510 71.676
R1523 B.n663 B.n511 71.676
R1524 B.n659 B.n512 71.676
R1525 B.n655 B.n513 71.676
R1526 B.n651 B.n514 71.676
R1527 B.n647 B.n515 71.676
R1528 B.n643 B.n516 71.676
R1529 B.n639 B.n517 71.676
R1530 B.n635 B.n518 71.676
R1531 B.n631 B.n519 71.676
R1532 B.n627 B.n520 71.676
R1533 B.n623 B.n521 71.676
R1534 B.n619 B.n522 71.676
R1535 B.n615 B.n523 71.676
R1536 B.n611 B.n524 71.676
R1537 B.n607 B.n525 71.676
R1538 B.n603 B.n526 71.676
R1539 B.n599 B.n527 71.676
R1540 B.n595 B.n528 71.676
R1541 B.n591 B.n529 71.676
R1542 B.n587 B.n530 71.676
R1543 B.n583 B.n531 71.676
R1544 B.n579 B.n532 71.676
R1545 B.n575 B.n533 71.676
R1546 B.n571 B.n534 71.676
R1547 B.n567 B.n535 71.676
R1548 B.n563 B.n536 71.676
R1549 B.n559 B.n537 71.676
R1550 B.n555 B.n538 71.676
R1551 B.n551 B.n539 71.676
R1552 B.n540 B.n488 71.676
R1553 B.n548 B.n547 59.5399
R1554 B.n545 B.n544 59.5399
R1555 B.n261 B.n162 59.5399
R1556 B.n282 B.n160 59.5399
R1557 B.n547 B.n546 53.9157
R1558 B.n544 B.n543 53.9157
R1559 B.n162 B.n161 53.9157
R1560 B.n160 B.n159 53.9157
R1561 B.n766 B.n485 37.6357
R1562 B.n766 B.n481 37.6357
R1563 B.n772 B.n481 37.6357
R1564 B.n772 B.n477 37.6357
R1565 B.n778 B.n477 37.6357
R1566 B.n778 B.n473 37.6357
R1567 B.n784 B.n473 37.6357
R1568 B.n790 B.n469 37.6357
R1569 B.n790 B.n465 37.6357
R1570 B.n796 B.n465 37.6357
R1571 B.n796 B.n461 37.6357
R1572 B.n802 B.n461 37.6357
R1573 B.n802 B.n457 37.6357
R1574 B.n808 B.n457 37.6357
R1575 B.n808 B.n453 37.6357
R1576 B.n815 B.n453 37.6357
R1577 B.n815 B.n814 37.6357
R1578 B.n821 B.n446 37.6357
R1579 B.n827 B.n446 37.6357
R1580 B.n827 B.n442 37.6357
R1581 B.n833 B.n442 37.6357
R1582 B.n833 B.n438 37.6357
R1583 B.n840 B.n438 37.6357
R1584 B.n840 B.n839 37.6357
R1585 B.n846 B.n431 37.6357
R1586 B.n852 B.n431 37.6357
R1587 B.n852 B.n427 37.6357
R1588 B.n858 B.n427 37.6357
R1589 B.n858 B.n423 37.6357
R1590 B.n865 B.n423 37.6357
R1591 B.n865 B.n864 37.6357
R1592 B.n871 B.n416 37.6357
R1593 B.n877 B.n416 37.6357
R1594 B.n877 B.n412 37.6357
R1595 B.n883 B.n412 37.6357
R1596 B.n883 B.n408 37.6357
R1597 B.n889 B.n408 37.6357
R1598 B.n889 B.n404 37.6357
R1599 B.n895 B.n404 37.6357
R1600 B.n901 B.n400 37.6357
R1601 B.n901 B.n396 37.6357
R1602 B.n907 B.n396 37.6357
R1603 B.n907 B.n392 37.6357
R1604 B.n913 B.n392 37.6357
R1605 B.n913 B.n388 37.6357
R1606 B.n919 B.n388 37.6357
R1607 B.n926 B.n384 37.6357
R1608 B.n926 B.n380 37.6357
R1609 B.n932 B.n380 37.6357
R1610 B.n932 B.n4 37.6357
R1611 B.n1125 B.n4 37.6357
R1612 B.n1125 B.n1124 37.6357
R1613 B.n1124 B.n1123 37.6357
R1614 B.n1123 B.n8 37.6357
R1615 B.n1117 B.n8 37.6357
R1616 B.n1117 B.n1116 37.6357
R1617 B.n1115 B.n15 37.6357
R1618 B.n1109 B.n15 37.6357
R1619 B.n1109 B.n1108 37.6357
R1620 B.n1108 B.n1107 37.6357
R1621 B.n1107 B.n22 37.6357
R1622 B.n1101 B.n22 37.6357
R1623 B.n1101 B.n1100 37.6357
R1624 B.n1099 B.n29 37.6357
R1625 B.n1093 B.n29 37.6357
R1626 B.n1093 B.n1092 37.6357
R1627 B.n1092 B.n1091 37.6357
R1628 B.n1091 B.n36 37.6357
R1629 B.n1085 B.n36 37.6357
R1630 B.n1085 B.n1084 37.6357
R1631 B.n1084 B.n1083 37.6357
R1632 B.n1077 B.n46 37.6357
R1633 B.n1077 B.n1076 37.6357
R1634 B.n1076 B.n1075 37.6357
R1635 B.n1075 B.n50 37.6357
R1636 B.n1069 B.n50 37.6357
R1637 B.n1069 B.n1068 37.6357
R1638 B.n1068 B.n1067 37.6357
R1639 B.n1061 B.n60 37.6357
R1640 B.n1061 B.n1060 37.6357
R1641 B.n1060 B.n1059 37.6357
R1642 B.n1059 B.n64 37.6357
R1643 B.n1053 B.n64 37.6357
R1644 B.n1053 B.n1052 37.6357
R1645 B.n1052 B.n1051 37.6357
R1646 B.n1045 B.n74 37.6357
R1647 B.n1045 B.n1044 37.6357
R1648 B.n1044 B.n1043 37.6357
R1649 B.n1043 B.n78 37.6357
R1650 B.n1037 B.n78 37.6357
R1651 B.n1037 B.n1036 37.6357
R1652 B.n1036 B.n1035 37.6357
R1653 B.n1035 B.n85 37.6357
R1654 B.n1029 B.n85 37.6357
R1655 B.n1029 B.n1028 37.6357
R1656 B.n1027 B.n92 37.6357
R1657 B.n1021 B.n92 37.6357
R1658 B.n1021 B.n1020 37.6357
R1659 B.n1020 B.n1019 37.6357
R1660 B.n1019 B.n99 37.6357
R1661 B.n1013 B.n99 37.6357
R1662 B.n1013 B.n1012 37.6357
R1663 B.n864 B.t6 35.9753
R1664 B.n46 B.t9 35.9753
R1665 B.n1008 B.n1007 34.8103
R1666 B.n164 B.n101 34.8103
R1667 B.n763 B.n762 34.8103
R1668 B.n757 B.n483 34.8103
R1669 B.t0 B.n400 32.6546
R1670 B.n1100 B.t3 32.6546
R1671 B.t11 B.n469 29.3338
R1672 B.n839 B.t8 29.3338
R1673 B.n60 B.t2 29.3338
R1674 B.n1028 B.t18 29.3338
R1675 B.t5 B.n384 26.0131
R1676 B.n1116 B.t7 26.0131
R1677 B.n814 B.t4 22.6923
R1678 B.n74 B.t1 22.6923
R1679 B B.n1127 18.0485
R1680 B.n821 B.t4 14.9439
R1681 B.n1051 B.t1 14.9439
R1682 B.n919 B.t5 11.6231
R1683 B.t7 B.n1115 11.6231
R1684 B.n165 B.n164 10.6151
R1685 B.n168 B.n165 10.6151
R1686 B.n169 B.n168 10.6151
R1687 B.n172 B.n169 10.6151
R1688 B.n173 B.n172 10.6151
R1689 B.n176 B.n173 10.6151
R1690 B.n177 B.n176 10.6151
R1691 B.n180 B.n177 10.6151
R1692 B.n181 B.n180 10.6151
R1693 B.n184 B.n181 10.6151
R1694 B.n185 B.n184 10.6151
R1695 B.n188 B.n185 10.6151
R1696 B.n189 B.n188 10.6151
R1697 B.n192 B.n189 10.6151
R1698 B.n193 B.n192 10.6151
R1699 B.n196 B.n193 10.6151
R1700 B.n197 B.n196 10.6151
R1701 B.n200 B.n197 10.6151
R1702 B.n201 B.n200 10.6151
R1703 B.n204 B.n201 10.6151
R1704 B.n205 B.n204 10.6151
R1705 B.n208 B.n205 10.6151
R1706 B.n209 B.n208 10.6151
R1707 B.n212 B.n209 10.6151
R1708 B.n213 B.n212 10.6151
R1709 B.n216 B.n213 10.6151
R1710 B.n217 B.n216 10.6151
R1711 B.n220 B.n217 10.6151
R1712 B.n221 B.n220 10.6151
R1713 B.n224 B.n221 10.6151
R1714 B.n225 B.n224 10.6151
R1715 B.n228 B.n225 10.6151
R1716 B.n229 B.n228 10.6151
R1717 B.n232 B.n229 10.6151
R1718 B.n233 B.n232 10.6151
R1719 B.n236 B.n233 10.6151
R1720 B.n237 B.n236 10.6151
R1721 B.n240 B.n237 10.6151
R1722 B.n241 B.n240 10.6151
R1723 B.n244 B.n241 10.6151
R1724 B.n245 B.n244 10.6151
R1725 B.n248 B.n245 10.6151
R1726 B.n249 B.n248 10.6151
R1727 B.n252 B.n249 10.6151
R1728 B.n253 B.n252 10.6151
R1729 B.n256 B.n253 10.6151
R1730 B.n257 B.n256 10.6151
R1731 B.n260 B.n257 10.6151
R1732 B.n265 B.n262 10.6151
R1733 B.n266 B.n265 10.6151
R1734 B.n269 B.n266 10.6151
R1735 B.n270 B.n269 10.6151
R1736 B.n273 B.n270 10.6151
R1737 B.n274 B.n273 10.6151
R1738 B.n277 B.n274 10.6151
R1739 B.n278 B.n277 10.6151
R1740 B.n281 B.n278 10.6151
R1741 B.n286 B.n283 10.6151
R1742 B.n287 B.n286 10.6151
R1743 B.n290 B.n287 10.6151
R1744 B.n291 B.n290 10.6151
R1745 B.n294 B.n291 10.6151
R1746 B.n295 B.n294 10.6151
R1747 B.n298 B.n295 10.6151
R1748 B.n299 B.n298 10.6151
R1749 B.n302 B.n299 10.6151
R1750 B.n303 B.n302 10.6151
R1751 B.n306 B.n303 10.6151
R1752 B.n307 B.n306 10.6151
R1753 B.n310 B.n307 10.6151
R1754 B.n311 B.n310 10.6151
R1755 B.n314 B.n311 10.6151
R1756 B.n315 B.n314 10.6151
R1757 B.n318 B.n315 10.6151
R1758 B.n319 B.n318 10.6151
R1759 B.n322 B.n319 10.6151
R1760 B.n323 B.n322 10.6151
R1761 B.n326 B.n323 10.6151
R1762 B.n327 B.n326 10.6151
R1763 B.n330 B.n327 10.6151
R1764 B.n331 B.n330 10.6151
R1765 B.n334 B.n331 10.6151
R1766 B.n335 B.n334 10.6151
R1767 B.n338 B.n335 10.6151
R1768 B.n339 B.n338 10.6151
R1769 B.n342 B.n339 10.6151
R1770 B.n343 B.n342 10.6151
R1771 B.n346 B.n343 10.6151
R1772 B.n347 B.n346 10.6151
R1773 B.n350 B.n347 10.6151
R1774 B.n351 B.n350 10.6151
R1775 B.n354 B.n351 10.6151
R1776 B.n355 B.n354 10.6151
R1777 B.n358 B.n355 10.6151
R1778 B.n359 B.n358 10.6151
R1779 B.n362 B.n359 10.6151
R1780 B.n363 B.n362 10.6151
R1781 B.n366 B.n363 10.6151
R1782 B.n367 B.n366 10.6151
R1783 B.n370 B.n367 10.6151
R1784 B.n371 B.n370 10.6151
R1785 B.n374 B.n371 10.6151
R1786 B.n376 B.n374 10.6151
R1787 B.n377 B.n376 10.6151
R1788 B.n1008 B.n377 10.6151
R1789 B.n764 B.n763 10.6151
R1790 B.n764 B.n479 10.6151
R1791 B.n774 B.n479 10.6151
R1792 B.n775 B.n774 10.6151
R1793 B.n776 B.n775 10.6151
R1794 B.n776 B.n471 10.6151
R1795 B.n786 B.n471 10.6151
R1796 B.n787 B.n786 10.6151
R1797 B.n788 B.n787 10.6151
R1798 B.n788 B.n463 10.6151
R1799 B.n798 B.n463 10.6151
R1800 B.n799 B.n798 10.6151
R1801 B.n800 B.n799 10.6151
R1802 B.n800 B.n455 10.6151
R1803 B.n810 B.n455 10.6151
R1804 B.n811 B.n810 10.6151
R1805 B.n812 B.n811 10.6151
R1806 B.n812 B.n448 10.6151
R1807 B.n823 B.n448 10.6151
R1808 B.n824 B.n823 10.6151
R1809 B.n825 B.n824 10.6151
R1810 B.n825 B.n440 10.6151
R1811 B.n835 B.n440 10.6151
R1812 B.n836 B.n835 10.6151
R1813 B.n837 B.n836 10.6151
R1814 B.n837 B.n433 10.6151
R1815 B.n848 B.n433 10.6151
R1816 B.n849 B.n848 10.6151
R1817 B.n850 B.n849 10.6151
R1818 B.n850 B.n425 10.6151
R1819 B.n860 B.n425 10.6151
R1820 B.n861 B.n860 10.6151
R1821 B.n862 B.n861 10.6151
R1822 B.n862 B.n418 10.6151
R1823 B.n873 B.n418 10.6151
R1824 B.n874 B.n873 10.6151
R1825 B.n875 B.n874 10.6151
R1826 B.n875 B.n410 10.6151
R1827 B.n885 B.n410 10.6151
R1828 B.n886 B.n885 10.6151
R1829 B.n887 B.n886 10.6151
R1830 B.n887 B.n402 10.6151
R1831 B.n897 B.n402 10.6151
R1832 B.n898 B.n897 10.6151
R1833 B.n899 B.n898 10.6151
R1834 B.n899 B.n394 10.6151
R1835 B.n909 B.n394 10.6151
R1836 B.n910 B.n909 10.6151
R1837 B.n911 B.n910 10.6151
R1838 B.n911 B.n386 10.6151
R1839 B.n921 B.n386 10.6151
R1840 B.n922 B.n921 10.6151
R1841 B.n924 B.n922 10.6151
R1842 B.n924 B.n923 10.6151
R1843 B.n923 B.n378 10.6151
R1844 B.n935 B.n378 10.6151
R1845 B.n936 B.n935 10.6151
R1846 B.n937 B.n936 10.6151
R1847 B.n938 B.n937 10.6151
R1848 B.n940 B.n938 10.6151
R1849 B.n941 B.n940 10.6151
R1850 B.n942 B.n941 10.6151
R1851 B.n943 B.n942 10.6151
R1852 B.n945 B.n943 10.6151
R1853 B.n946 B.n945 10.6151
R1854 B.n947 B.n946 10.6151
R1855 B.n948 B.n947 10.6151
R1856 B.n950 B.n948 10.6151
R1857 B.n951 B.n950 10.6151
R1858 B.n952 B.n951 10.6151
R1859 B.n953 B.n952 10.6151
R1860 B.n955 B.n953 10.6151
R1861 B.n956 B.n955 10.6151
R1862 B.n957 B.n956 10.6151
R1863 B.n958 B.n957 10.6151
R1864 B.n960 B.n958 10.6151
R1865 B.n961 B.n960 10.6151
R1866 B.n962 B.n961 10.6151
R1867 B.n963 B.n962 10.6151
R1868 B.n965 B.n963 10.6151
R1869 B.n966 B.n965 10.6151
R1870 B.n967 B.n966 10.6151
R1871 B.n968 B.n967 10.6151
R1872 B.n970 B.n968 10.6151
R1873 B.n971 B.n970 10.6151
R1874 B.n972 B.n971 10.6151
R1875 B.n973 B.n972 10.6151
R1876 B.n975 B.n973 10.6151
R1877 B.n976 B.n975 10.6151
R1878 B.n977 B.n976 10.6151
R1879 B.n978 B.n977 10.6151
R1880 B.n980 B.n978 10.6151
R1881 B.n981 B.n980 10.6151
R1882 B.n982 B.n981 10.6151
R1883 B.n983 B.n982 10.6151
R1884 B.n985 B.n983 10.6151
R1885 B.n986 B.n985 10.6151
R1886 B.n987 B.n986 10.6151
R1887 B.n988 B.n987 10.6151
R1888 B.n990 B.n988 10.6151
R1889 B.n991 B.n990 10.6151
R1890 B.n992 B.n991 10.6151
R1891 B.n993 B.n992 10.6151
R1892 B.n995 B.n993 10.6151
R1893 B.n996 B.n995 10.6151
R1894 B.n997 B.n996 10.6151
R1895 B.n998 B.n997 10.6151
R1896 B.n1000 B.n998 10.6151
R1897 B.n1001 B.n1000 10.6151
R1898 B.n1002 B.n1001 10.6151
R1899 B.n1003 B.n1002 10.6151
R1900 B.n1005 B.n1003 10.6151
R1901 B.n1006 B.n1005 10.6151
R1902 B.n1007 B.n1006 10.6151
R1903 B.n757 B.n756 10.6151
R1904 B.n756 B.n755 10.6151
R1905 B.n755 B.n754 10.6151
R1906 B.n754 B.n752 10.6151
R1907 B.n752 B.n749 10.6151
R1908 B.n749 B.n748 10.6151
R1909 B.n748 B.n745 10.6151
R1910 B.n745 B.n744 10.6151
R1911 B.n744 B.n741 10.6151
R1912 B.n741 B.n740 10.6151
R1913 B.n740 B.n737 10.6151
R1914 B.n737 B.n736 10.6151
R1915 B.n736 B.n733 10.6151
R1916 B.n733 B.n732 10.6151
R1917 B.n732 B.n729 10.6151
R1918 B.n729 B.n728 10.6151
R1919 B.n728 B.n725 10.6151
R1920 B.n725 B.n724 10.6151
R1921 B.n724 B.n721 10.6151
R1922 B.n721 B.n720 10.6151
R1923 B.n720 B.n717 10.6151
R1924 B.n717 B.n716 10.6151
R1925 B.n716 B.n713 10.6151
R1926 B.n713 B.n712 10.6151
R1927 B.n712 B.n709 10.6151
R1928 B.n709 B.n708 10.6151
R1929 B.n708 B.n705 10.6151
R1930 B.n705 B.n704 10.6151
R1931 B.n704 B.n701 10.6151
R1932 B.n701 B.n700 10.6151
R1933 B.n700 B.n697 10.6151
R1934 B.n697 B.n696 10.6151
R1935 B.n696 B.n693 10.6151
R1936 B.n693 B.n692 10.6151
R1937 B.n692 B.n689 10.6151
R1938 B.n689 B.n688 10.6151
R1939 B.n688 B.n685 10.6151
R1940 B.n685 B.n684 10.6151
R1941 B.n684 B.n681 10.6151
R1942 B.n681 B.n680 10.6151
R1943 B.n680 B.n677 10.6151
R1944 B.n677 B.n676 10.6151
R1945 B.n676 B.n673 10.6151
R1946 B.n673 B.n672 10.6151
R1947 B.n672 B.n669 10.6151
R1948 B.n669 B.n668 10.6151
R1949 B.n668 B.n665 10.6151
R1950 B.n665 B.n664 10.6151
R1951 B.n661 B.n660 10.6151
R1952 B.n660 B.n657 10.6151
R1953 B.n657 B.n656 10.6151
R1954 B.n656 B.n653 10.6151
R1955 B.n653 B.n652 10.6151
R1956 B.n652 B.n649 10.6151
R1957 B.n649 B.n648 10.6151
R1958 B.n648 B.n645 10.6151
R1959 B.n645 B.n644 10.6151
R1960 B.n641 B.n640 10.6151
R1961 B.n640 B.n637 10.6151
R1962 B.n637 B.n636 10.6151
R1963 B.n636 B.n633 10.6151
R1964 B.n633 B.n632 10.6151
R1965 B.n632 B.n629 10.6151
R1966 B.n629 B.n628 10.6151
R1967 B.n628 B.n625 10.6151
R1968 B.n625 B.n624 10.6151
R1969 B.n624 B.n621 10.6151
R1970 B.n621 B.n620 10.6151
R1971 B.n620 B.n617 10.6151
R1972 B.n617 B.n616 10.6151
R1973 B.n616 B.n613 10.6151
R1974 B.n613 B.n612 10.6151
R1975 B.n612 B.n609 10.6151
R1976 B.n609 B.n608 10.6151
R1977 B.n608 B.n605 10.6151
R1978 B.n605 B.n604 10.6151
R1979 B.n604 B.n601 10.6151
R1980 B.n601 B.n600 10.6151
R1981 B.n600 B.n597 10.6151
R1982 B.n597 B.n596 10.6151
R1983 B.n596 B.n593 10.6151
R1984 B.n593 B.n592 10.6151
R1985 B.n592 B.n589 10.6151
R1986 B.n589 B.n588 10.6151
R1987 B.n588 B.n585 10.6151
R1988 B.n585 B.n584 10.6151
R1989 B.n584 B.n581 10.6151
R1990 B.n581 B.n580 10.6151
R1991 B.n580 B.n577 10.6151
R1992 B.n577 B.n576 10.6151
R1993 B.n576 B.n573 10.6151
R1994 B.n573 B.n572 10.6151
R1995 B.n572 B.n569 10.6151
R1996 B.n569 B.n568 10.6151
R1997 B.n568 B.n565 10.6151
R1998 B.n565 B.n564 10.6151
R1999 B.n564 B.n561 10.6151
R2000 B.n561 B.n560 10.6151
R2001 B.n560 B.n557 10.6151
R2002 B.n557 B.n556 10.6151
R2003 B.n556 B.n553 10.6151
R2004 B.n553 B.n552 10.6151
R2005 B.n552 B.n549 10.6151
R2006 B.n549 B.n487 10.6151
R2007 B.n762 B.n487 10.6151
R2008 B.n768 B.n483 10.6151
R2009 B.n769 B.n768 10.6151
R2010 B.n770 B.n769 10.6151
R2011 B.n770 B.n475 10.6151
R2012 B.n780 B.n475 10.6151
R2013 B.n781 B.n780 10.6151
R2014 B.n782 B.n781 10.6151
R2015 B.n782 B.n467 10.6151
R2016 B.n792 B.n467 10.6151
R2017 B.n793 B.n792 10.6151
R2018 B.n794 B.n793 10.6151
R2019 B.n794 B.n459 10.6151
R2020 B.n804 B.n459 10.6151
R2021 B.n805 B.n804 10.6151
R2022 B.n806 B.n805 10.6151
R2023 B.n806 B.n451 10.6151
R2024 B.n817 B.n451 10.6151
R2025 B.n818 B.n817 10.6151
R2026 B.n819 B.n818 10.6151
R2027 B.n819 B.n444 10.6151
R2028 B.n829 B.n444 10.6151
R2029 B.n830 B.n829 10.6151
R2030 B.n831 B.n830 10.6151
R2031 B.n831 B.n436 10.6151
R2032 B.n842 B.n436 10.6151
R2033 B.n843 B.n842 10.6151
R2034 B.n844 B.n843 10.6151
R2035 B.n844 B.n429 10.6151
R2036 B.n854 B.n429 10.6151
R2037 B.n855 B.n854 10.6151
R2038 B.n856 B.n855 10.6151
R2039 B.n856 B.n421 10.6151
R2040 B.n867 B.n421 10.6151
R2041 B.n868 B.n867 10.6151
R2042 B.n869 B.n868 10.6151
R2043 B.n869 B.n414 10.6151
R2044 B.n879 B.n414 10.6151
R2045 B.n880 B.n879 10.6151
R2046 B.n881 B.n880 10.6151
R2047 B.n881 B.n406 10.6151
R2048 B.n891 B.n406 10.6151
R2049 B.n892 B.n891 10.6151
R2050 B.n893 B.n892 10.6151
R2051 B.n893 B.n398 10.6151
R2052 B.n903 B.n398 10.6151
R2053 B.n904 B.n903 10.6151
R2054 B.n905 B.n904 10.6151
R2055 B.n905 B.n390 10.6151
R2056 B.n915 B.n390 10.6151
R2057 B.n916 B.n915 10.6151
R2058 B.n917 B.n916 10.6151
R2059 B.n917 B.n382 10.6151
R2060 B.n928 B.n382 10.6151
R2061 B.n929 B.n928 10.6151
R2062 B.n930 B.n929 10.6151
R2063 B.n930 B.n0 10.6151
R2064 B.n1121 B.n1 10.6151
R2065 B.n1121 B.n1120 10.6151
R2066 B.n1120 B.n1119 10.6151
R2067 B.n1119 B.n10 10.6151
R2068 B.n1113 B.n10 10.6151
R2069 B.n1113 B.n1112 10.6151
R2070 B.n1112 B.n1111 10.6151
R2071 B.n1111 B.n17 10.6151
R2072 B.n1105 B.n17 10.6151
R2073 B.n1105 B.n1104 10.6151
R2074 B.n1104 B.n1103 10.6151
R2075 B.n1103 B.n24 10.6151
R2076 B.n1097 B.n24 10.6151
R2077 B.n1097 B.n1096 10.6151
R2078 B.n1096 B.n1095 10.6151
R2079 B.n1095 B.n31 10.6151
R2080 B.n1089 B.n31 10.6151
R2081 B.n1089 B.n1088 10.6151
R2082 B.n1088 B.n1087 10.6151
R2083 B.n1087 B.n38 10.6151
R2084 B.n1081 B.n38 10.6151
R2085 B.n1081 B.n1080 10.6151
R2086 B.n1080 B.n1079 10.6151
R2087 B.n1079 B.n44 10.6151
R2088 B.n1073 B.n44 10.6151
R2089 B.n1073 B.n1072 10.6151
R2090 B.n1072 B.n1071 10.6151
R2091 B.n1071 B.n52 10.6151
R2092 B.n1065 B.n52 10.6151
R2093 B.n1065 B.n1064 10.6151
R2094 B.n1064 B.n1063 10.6151
R2095 B.n1063 B.n58 10.6151
R2096 B.n1057 B.n58 10.6151
R2097 B.n1057 B.n1056 10.6151
R2098 B.n1056 B.n1055 10.6151
R2099 B.n1055 B.n66 10.6151
R2100 B.n1049 B.n66 10.6151
R2101 B.n1049 B.n1048 10.6151
R2102 B.n1048 B.n1047 10.6151
R2103 B.n1047 B.n72 10.6151
R2104 B.n1041 B.n72 10.6151
R2105 B.n1041 B.n1040 10.6151
R2106 B.n1040 B.n1039 10.6151
R2107 B.n1039 B.n80 10.6151
R2108 B.n1033 B.n80 10.6151
R2109 B.n1033 B.n1032 10.6151
R2110 B.n1032 B.n1031 10.6151
R2111 B.n1031 B.n87 10.6151
R2112 B.n1025 B.n87 10.6151
R2113 B.n1025 B.n1024 10.6151
R2114 B.n1024 B.n1023 10.6151
R2115 B.n1023 B.n94 10.6151
R2116 B.n1017 B.n94 10.6151
R2117 B.n1017 B.n1016 10.6151
R2118 B.n1016 B.n1015 10.6151
R2119 B.n1015 B.n101 10.6151
R2120 B.n261 B.n260 9.36635
R2121 B.n283 B.n282 9.36635
R2122 B.n664 B.n545 9.36635
R2123 B.n641 B.n548 9.36635
R2124 B.n784 B.t11 8.30239
R2125 B.n846 B.t8 8.30239
R2126 B.n1067 B.t2 8.30239
R2127 B.t18 B.n1027 8.30239
R2128 B.n895 B.t0 4.98163
R2129 B.t3 B.n1099 4.98163
R2130 B.n1127 B.n0 2.81026
R2131 B.n1127 B.n1 2.81026
R2132 B.n871 B.t6 1.66088
R2133 B.n1083 B.t9 1.66088
R2134 B.n262 B.n261 1.24928
R2135 B.n282 B.n281 1.24928
R2136 B.n661 B.n545 1.24928
R2137 B.n644 B.n548 1.24928
R2138 VN.n9 VN.t5 176.114
R2139 VN.n50 VN.t6 176.114
R2140 VN.n77 VN.n40 161.3
R2141 VN.n76 VN.n75 161.3
R2142 VN.n74 VN.n41 161.3
R2143 VN.n73 VN.n72 161.3
R2144 VN.n71 VN.n42 161.3
R2145 VN.n69 VN.n68 161.3
R2146 VN.n67 VN.n43 161.3
R2147 VN.n66 VN.n65 161.3
R2148 VN.n64 VN.n44 161.3
R2149 VN.n63 VN.n62 161.3
R2150 VN.n61 VN.n45 161.3
R2151 VN.n60 VN.n59 161.3
R2152 VN.n58 VN.n46 161.3
R2153 VN.n57 VN.n56 161.3
R2154 VN.n55 VN.n48 161.3
R2155 VN.n54 VN.n53 161.3
R2156 VN.n52 VN.n49 161.3
R2157 VN.n37 VN.n0 161.3
R2158 VN.n36 VN.n35 161.3
R2159 VN.n34 VN.n1 161.3
R2160 VN.n33 VN.n32 161.3
R2161 VN.n31 VN.n2 161.3
R2162 VN.n29 VN.n28 161.3
R2163 VN.n27 VN.n3 161.3
R2164 VN.n26 VN.n25 161.3
R2165 VN.n24 VN.n4 161.3
R2166 VN.n23 VN.n22 161.3
R2167 VN.n21 VN.n5 161.3
R2168 VN.n20 VN.n19 161.3
R2169 VN.n17 VN.n6 161.3
R2170 VN.n16 VN.n15 161.3
R2171 VN.n14 VN.n7 161.3
R2172 VN.n13 VN.n12 161.3
R2173 VN.n11 VN.n8 161.3
R2174 VN.n10 VN.t2 143.617
R2175 VN.n18 VN.t7 143.617
R2176 VN.n30 VN.t3 143.617
R2177 VN.n38 VN.t8 143.617
R2178 VN.n51 VN.t9 143.617
R2179 VN.n47 VN.t4 143.617
R2180 VN.n70 VN.t0 143.617
R2181 VN.n78 VN.t1 143.617
R2182 VN.n39 VN.n38 95.6613
R2183 VN.n79 VN.n78 95.6613
R2184 VN.n10 VN.n9 71.1838
R2185 VN.n51 VN.n50 71.1838
R2186 VN VN.n79 54.6118
R2187 VN.n16 VN.n7 54.1398
R2188 VN.n25 VN.n24 54.1398
R2189 VN.n57 VN.n48 54.1398
R2190 VN.n65 VN.n64 54.1398
R2191 VN.n32 VN.n1 48.3272
R2192 VN.n72 VN.n41 48.3272
R2193 VN.n36 VN.n1 32.8269
R2194 VN.n76 VN.n41 32.8269
R2195 VN.n17 VN.n16 27.0143
R2196 VN.n24 VN.n23 27.0143
R2197 VN.n58 VN.n57 27.0143
R2198 VN.n64 VN.n63 27.0143
R2199 VN.n12 VN.n11 24.5923
R2200 VN.n12 VN.n7 24.5923
R2201 VN.n19 VN.n17 24.5923
R2202 VN.n23 VN.n5 24.5923
R2203 VN.n25 VN.n3 24.5923
R2204 VN.n29 VN.n3 24.5923
R2205 VN.n32 VN.n31 24.5923
R2206 VN.n37 VN.n36 24.5923
R2207 VN.n53 VN.n48 24.5923
R2208 VN.n53 VN.n52 24.5923
R2209 VN.n63 VN.n45 24.5923
R2210 VN.n59 VN.n58 24.5923
R2211 VN.n72 VN.n71 24.5923
R2212 VN.n69 VN.n43 24.5923
R2213 VN.n65 VN.n43 24.5923
R2214 VN.n77 VN.n76 24.5923
R2215 VN.n31 VN.n30 23.1168
R2216 VN.n71 VN.n70 23.1168
R2217 VN.n38 VN.n37 15.2474
R2218 VN.n78 VN.n77 15.2474
R2219 VN.n19 VN.n18 12.2964
R2220 VN.n18 VN.n5 12.2964
R2221 VN.n47 VN.n45 12.2964
R2222 VN.n59 VN.n47 12.2964
R2223 VN.n50 VN.n49 9.47955
R2224 VN.n9 VN.n8 9.47955
R2225 VN.n11 VN.n10 1.47601
R2226 VN.n30 VN.n29 1.47601
R2227 VN.n52 VN.n51 1.47601
R2228 VN.n70 VN.n69 1.47601
R2229 VN.n79 VN.n40 0.278335
R2230 VN.n39 VN.n0 0.278335
R2231 VN.n75 VN.n40 0.189894
R2232 VN.n75 VN.n74 0.189894
R2233 VN.n74 VN.n73 0.189894
R2234 VN.n73 VN.n42 0.189894
R2235 VN.n68 VN.n42 0.189894
R2236 VN.n68 VN.n67 0.189894
R2237 VN.n67 VN.n66 0.189894
R2238 VN.n66 VN.n44 0.189894
R2239 VN.n62 VN.n44 0.189894
R2240 VN.n62 VN.n61 0.189894
R2241 VN.n61 VN.n60 0.189894
R2242 VN.n60 VN.n46 0.189894
R2243 VN.n56 VN.n46 0.189894
R2244 VN.n56 VN.n55 0.189894
R2245 VN.n55 VN.n54 0.189894
R2246 VN.n54 VN.n49 0.189894
R2247 VN.n13 VN.n8 0.189894
R2248 VN.n14 VN.n13 0.189894
R2249 VN.n15 VN.n14 0.189894
R2250 VN.n15 VN.n6 0.189894
R2251 VN.n20 VN.n6 0.189894
R2252 VN.n21 VN.n20 0.189894
R2253 VN.n22 VN.n21 0.189894
R2254 VN.n22 VN.n4 0.189894
R2255 VN.n26 VN.n4 0.189894
R2256 VN.n27 VN.n26 0.189894
R2257 VN.n28 VN.n27 0.189894
R2258 VN.n28 VN.n2 0.189894
R2259 VN.n33 VN.n2 0.189894
R2260 VN.n34 VN.n33 0.189894
R2261 VN.n35 VN.n34 0.189894
R2262 VN.n35 VN.n0 0.189894
R2263 VN VN.n39 0.153485
R2264 VDD2.n1 VDD2.t4 64.3492
R2265 VDD2.n3 VDD2.n2 62.3387
R2266 VDD2 VDD2.n7 62.3359
R2267 VDD2.n4 VDD2.t8 61.9529
R2268 VDD2.n6 VDD2.n5 60.5967
R2269 VDD2.n1 VDD2.n0 60.5967
R2270 VDD2.n4 VDD2.n3 47.6851
R2271 VDD2.n6 VDD2.n4 2.39705
R2272 VDD2.n7 VDD2.t0 1.35666
R2273 VDD2.n7 VDD2.t3 1.35666
R2274 VDD2.n5 VDD2.t9 1.35666
R2275 VDD2.n5 VDD2.t5 1.35666
R2276 VDD2.n2 VDD2.t6 1.35666
R2277 VDD2.n2 VDD2.t1 1.35666
R2278 VDD2.n0 VDD2.t7 1.35666
R2279 VDD2.n0 VDD2.t2 1.35666
R2280 VDD2 VDD2.n6 0.657828
R2281 VDD2.n3 VDD2.n1 0.544292
C0 VDD1 VN 0.153294f
C1 VDD2 VDD1 2.07672f
C2 VN VTAIL 13.1763f
C3 VDD2 VTAIL 11.656401f
C4 VDD1 VTAIL 11.6073f
C5 VN VP 8.6499f
C6 VDD2 VP 0.564943f
C7 VDD1 VP 13.1197f
C8 VP VTAIL 13.190599f
C9 VDD2 VN 12.7124f
C10 VDD2 B 7.50705f
C11 VDD1 B 7.46786f
C12 VTAIL B 9.119318f
C13 VN B 17.634401f
C14 VP B 16.108639f
C15 VDD2.t4 B 3.18419f
C16 VDD2.t7 B 0.275504f
C17 VDD2.t2 B 0.275504f
C18 VDD2.n0 B 2.48039f
C19 VDD2.n1 B 0.872514f
C20 VDD2.t6 B 0.275504f
C21 VDD2.t1 B 0.275504f
C22 VDD2.n2 B 2.4952f
C23 VDD2.n3 B 2.85929f
C24 VDD2.t8 B 3.16705f
C25 VDD2.n4 B 3.12567f
C26 VDD2.t9 B 0.275504f
C27 VDD2.t5 B 0.275504f
C28 VDD2.n5 B 2.48039f
C29 VDD2.n6 B 0.436813f
C30 VDD2.t0 B 0.275504f
C31 VDD2.t3 B 0.275504f
C32 VDD2.n7 B 2.49516f
C33 VN.n0 B 0.028733f
C34 VN.t8 B 2.13499f
C35 VN.n1 B 0.019449f
C36 VN.n2 B 0.021796f
C37 VN.t3 B 2.13499f
C38 VN.n3 B 0.040418f
C39 VN.n4 B 0.021796f
C40 VN.n5 B 0.030441f
C41 VN.n6 B 0.021796f
C42 VN.n7 B 0.038022f
C43 VN.n8 B 0.190915f
C44 VN.t2 B 2.13499f
C45 VN.t5 B 2.29634f
C46 VN.n9 B 0.792564f
C47 VN.n10 B 0.800731f
C48 VN.n11 B 0.021662f
C49 VN.n12 B 0.040418f
C50 VN.n13 B 0.021796f
C51 VN.n14 B 0.021796f
C52 VN.n15 B 0.021796f
C53 VN.n16 B 0.023734f
C54 VN.n17 B 0.042028f
C55 VN.t7 B 2.13499f
C56 VN.n18 B 0.748243f
C57 VN.n19 B 0.030441f
C58 VN.n20 B 0.021796f
C59 VN.n21 B 0.021796f
C60 VN.n22 B 0.021796f
C61 VN.n23 B 0.042028f
C62 VN.n24 B 0.023734f
C63 VN.n25 B 0.038022f
C64 VN.n26 B 0.021796f
C65 VN.n27 B 0.021796f
C66 VN.n28 B 0.021796f
C67 VN.n29 B 0.021662f
C68 VN.n30 B 0.748243f
C69 VN.n31 B 0.039221f
C70 VN.n32 B 0.040614f
C71 VN.n33 B 0.021796f
C72 VN.n34 B 0.021796f
C73 VN.n35 B 0.021796f
C74 VN.n36 B 0.043721f
C75 VN.n37 B 0.032835f
C76 VN.n38 B 0.823004f
C77 VN.n39 B 0.03139f
C78 VN.n40 B 0.028733f
C79 VN.t1 B 2.13499f
C80 VN.n41 B 0.019449f
C81 VN.n42 B 0.021796f
C82 VN.t0 B 2.13499f
C83 VN.n43 B 0.040418f
C84 VN.n44 B 0.021796f
C85 VN.n45 B 0.030441f
C86 VN.n46 B 0.021796f
C87 VN.t4 B 2.13499f
C88 VN.n47 B 0.748243f
C89 VN.n48 B 0.038022f
C90 VN.n49 B 0.190915f
C91 VN.t9 B 2.13499f
C92 VN.t6 B 2.29634f
C93 VN.n50 B 0.792564f
C94 VN.n51 B 0.800731f
C95 VN.n52 B 0.021662f
C96 VN.n53 B 0.040418f
C97 VN.n54 B 0.021796f
C98 VN.n55 B 0.021796f
C99 VN.n56 B 0.021796f
C100 VN.n57 B 0.023734f
C101 VN.n58 B 0.042028f
C102 VN.n59 B 0.030441f
C103 VN.n60 B 0.021796f
C104 VN.n61 B 0.021796f
C105 VN.n62 B 0.021796f
C106 VN.n63 B 0.042028f
C107 VN.n64 B 0.023734f
C108 VN.n65 B 0.038022f
C109 VN.n66 B 0.021796f
C110 VN.n67 B 0.021796f
C111 VN.n68 B 0.021796f
C112 VN.n69 B 0.021662f
C113 VN.n70 B 0.748243f
C114 VN.n71 B 0.039221f
C115 VN.n72 B 0.040614f
C116 VN.n73 B 0.021796f
C117 VN.n74 B 0.021796f
C118 VN.n75 B 0.021796f
C119 VN.n76 B 0.043721f
C120 VN.n77 B 0.032835f
C121 VN.n78 B 0.823004f
C122 VN.n79 B 1.37491f
C123 VDD1.t5 B 3.20956f
C124 VDD1.t4 B 0.277698f
C125 VDD1.t9 B 0.277698f
C126 VDD1.n0 B 2.50015f
C127 VDD1.n1 B 0.88724f
C128 VDD1.t1 B 3.20956f
C129 VDD1.t6 B 0.277698f
C130 VDD1.t3 B 0.277698f
C131 VDD1.n2 B 2.50015f
C132 VDD1.n3 B 0.879464f
C133 VDD1.t7 B 0.277698f
C134 VDD1.t2 B 0.277698f
C135 VDD1.n4 B 2.51508f
C136 VDD1.n5 B 3.00018f
C137 VDD1.t8 B 0.277698f
C138 VDD1.t0 B 0.277698f
C139 VDD1.n6 B 2.50015f
C140 VDD1.n7 B 3.19101f
C141 VTAIL.t15 B 0.279712f
C142 VTAIL.t3 B 0.279712f
C143 VTAIL.n0 B 2.44221f
C144 VTAIL.n1 B 0.523305f
C145 VTAIL.t7 B 3.11742f
C146 VTAIL.n2 B 0.653201f
C147 VTAIL.t12 B 0.279712f
C148 VTAIL.t5 B 0.279712f
C149 VTAIL.n3 B 2.44221f
C150 VTAIL.n4 B 0.62247f
C151 VTAIL.t4 B 0.279712f
C152 VTAIL.t11 B 0.279712f
C153 VTAIL.n5 B 2.44221f
C154 VTAIL.n6 B 2.12225f
C155 VTAIL.t17 B 0.279712f
C156 VTAIL.t19 B 0.279712f
C157 VTAIL.n7 B 2.44221f
C158 VTAIL.n8 B 2.12225f
C159 VTAIL.t14 B 0.279712f
C160 VTAIL.t0 B 0.279712f
C161 VTAIL.n9 B 2.44221f
C162 VTAIL.n10 B 0.622471f
C163 VTAIL.t16 B 3.11743f
C164 VTAIL.n11 B 0.653194f
C165 VTAIL.t10 B 0.279712f
C166 VTAIL.t13 B 0.279712f
C167 VTAIL.n12 B 2.44221f
C168 VTAIL.n13 B 0.565565f
C169 VTAIL.t6 B 0.279712f
C170 VTAIL.t8 B 0.279712f
C171 VTAIL.n14 B 2.44221f
C172 VTAIL.n15 B 0.622471f
C173 VTAIL.t9 B 3.11744f
C174 VTAIL.n16 B 2.02265f
C175 VTAIL.t1 B 3.11742f
C176 VTAIL.n17 B 2.02267f
C177 VTAIL.t18 B 0.279712f
C178 VTAIL.t2 B 0.279712f
C179 VTAIL.n18 B 2.44221f
C180 VTAIL.n19 B 0.477511f
C181 VP.n0 B 0.029092f
C182 VP.t7 B 2.16166f
C183 VP.n1 B 0.019692f
C184 VP.n2 B 0.022068f
C185 VP.t2 B 2.16166f
C186 VP.n3 B 0.040923f
C187 VP.n4 B 0.022068f
C188 VP.n5 B 0.030821f
C189 VP.n6 B 0.022068f
C190 VP.n7 B 0.038497f
C191 VP.n8 B 0.022068f
C192 VP.t3 B 2.16166f
C193 VP.n9 B 0.041121f
C194 VP.n10 B 0.022068f
C195 VP.t8 B 2.16166f
C196 VP.n11 B 0.833286f
C197 VP.n12 B 0.029092f
C198 VP.t9 B 2.16166f
C199 VP.n13 B 0.019692f
C200 VP.n14 B 0.022068f
C201 VP.t1 B 2.16166f
C202 VP.n15 B 0.040923f
C203 VP.n16 B 0.022068f
C204 VP.n17 B 0.030821f
C205 VP.n18 B 0.022068f
C206 VP.n19 B 0.038497f
C207 VP.n20 B 0.1933f
C208 VP.t5 B 2.16166f
C209 VP.t4 B 2.32503f
C210 VP.n21 B 0.802465f
C211 VP.n22 B 0.810735f
C212 VP.n23 B 0.021932f
C213 VP.n24 B 0.040923f
C214 VP.n25 B 0.022068f
C215 VP.n26 B 0.022068f
C216 VP.n27 B 0.022068f
C217 VP.n28 B 0.024031f
C218 VP.n29 B 0.042553f
C219 VP.t0 B 2.16166f
C220 VP.n30 B 0.757591f
C221 VP.n31 B 0.030821f
C222 VP.n32 B 0.022068f
C223 VP.n33 B 0.022068f
C224 VP.n34 B 0.022068f
C225 VP.n35 B 0.042553f
C226 VP.n36 B 0.024031f
C227 VP.n37 B 0.038497f
C228 VP.n38 B 0.022068f
C229 VP.n39 B 0.022068f
C230 VP.n40 B 0.022068f
C231 VP.n41 B 0.021932f
C232 VP.n42 B 0.757591f
C233 VP.n43 B 0.03971f
C234 VP.n44 B 0.041121f
C235 VP.n45 B 0.022068f
C236 VP.n46 B 0.022068f
C237 VP.n47 B 0.022068f
C238 VP.n48 B 0.044267f
C239 VP.n49 B 0.033246f
C240 VP.n50 B 0.833286f
C241 VP.n51 B 1.38038f
C242 VP.n52 B 1.39503f
C243 VP.n53 B 0.029092f
C244 VP.n54 B 0.033246f
C245 VP.n55 B 0.044267f
C246 VP.n56 B 0.019692f
C247 VP.n57 B 0.022068f
C248 VP.n58 B 0.022068f
C249 VP.n59 B 0.022068f
C250 VP.n60 B 0.03971f
C251 VP.n61 B 0.757591f
C252 VP.n62 B 0.021932f
C253 VP.n63 B 0.040923f
C254 VP.n64 B 0.022068f
C255 VP.n65 B 0.022068f
C256 VP.n66 B 0.022068f
C257 VP.n67 B 0.024031f
C258 VP.n68 B 0.042553f
C259 VP.t6 B 2.16166f
C260 VP.n69 B 0.757591f
C261 VP.n70 B 0.030821f
C262 VP.n71 B 0.022068f
C263 VP.n72 B 0.022068f
C264 VP.n73 B 0.022068f
C265 VP.n74 B 0.042553f
C266 VP.n75 B 0.024031f
C267 VP.n76 B 0.038497f
C268 VP.n77 B 0.022068f
C269 VP.n78 B 0.022068f
C270 VP.n79 B 0.022068f
C271 VP.n80 B 0.021932f
C272 VP.n81 B 0.757591f
C273 VP.n82 B 0.03971f
C274 VP.n83 B 0.041121f
C275 VP.n84 B 0.022068f
C276 VP.n85 B 0.022068f
C277 VP.n86 B 0.022068f
C278 VP.n87 B 0.044267f
C279 VP.n88 B 0.033246f
C280 VP.n89 B 0.833286f
C281 VP.n90 B 0.031782f
.ends

