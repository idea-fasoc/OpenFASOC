* NGSPICE file created from diff_pair_sample_0163.ext - technology: sky130A

.subckt diff_pair_sample_0163 VTAIL VN VP B VDD2 VDD1
X0 B.t21 B.t19 B.t20 B.t9 sky130_fd_pr__nfet_01v8 ad=0.8151 pd=4.96 as=0 ps=0 w=2.09 l=3.35
X1 VDD2.t7 VN.t0 VTAIL.t13 B.t4 sky130_fd_pr__nfet_01v8 ad=0.34485 pd=2.42 as=0.8151 ps=4.96 w=2.09 l=3.35
X2 VDD1.t7 VP.t0 VTAIL.t6 B.t5 sky130_fd_pr__nfet_01v8 ad=0.34485 pd=2.42 as=0.34485 ps=2.42 w=2.09 l=3.35
X3 VTAIL.t11 VN.t1 VDD2.t6 B.t7 sky130_fd_pr__nfet_01v8 ad=0.34485 pd=2.42 as=0.34485 ps=2.42 w=2.09 l=3.35
X4 B.t18 B.t16 B.t17 B.t13 sky130_fd_pr__nfet_01v8 ad=0.8151 pd=4.96 as=0 ps=0 w=2.09 l=3.35
X5 VTAIL.t4 VP.t1 VDD1.t6 B.t1 sky130_fd_pr__nfet_01v8 ad=0.8151 pd=4.96 as=0.34485 ps=2.42 w=2.09 l=3.35
X6 VTAIL.t3 VP.t2 VDD1.t5 B.t7 sky130_fd_pr__nfet_01v8 ad=0.34485 pd=2.42 as=0.34485 ps=2.42 w=2.09 l=3.35
X7 VTAIL.t12 VN.t2 VDD2.t5 B.t6 sky130_fd_pr__nfet_01v8 ad=0.8151 pd=4.96 as=0.34485 ps=2.42 w=2.09 l=3.35
X8 VTAIL.t5 VP.t3 VDD1.t4 B.t3 sky130_fd_pr__nfet_01v8 ad=0.34485 pd=2.42 as=0.34485 ps=2.42 w=2.09 l=3.35
X9 VDD1.t3 VP.t4 VTAIL.t2 B.t0 sky130_fd_pr__nfet_01v8 ad=0.34485 pd=2.42 as=0.34485 ps=2.42 w=2.09 l=3.35
X10 VDD2.t4 VN.t3 VTAIL.t14 B.t5 sky130_fd_pr__nfet_01v8 ad=0.34485 pd=2.42 as=0.34485 ps=2.42 w=2.09 l=3.35
X11 VDD1.t2 VP.t5 VTAIL.t1 B.t2 sky130_fd_pr__nfet_01v8 ad=0.34485 pd=2.42 as=0.8151 ps=4.96 w=2.09 l=3.35
X12 VDD1.t1 VP.t6 VTAIL.t0 B.t4 sky130_fd_pr__nfet_01v8 ad=0.34485 pd=2.42 as=0.8151 ps=4.96 w=2.09 l=3.35
X13 VTAIL.t7 VP.t7 VDD1.t0 B.t6 sky130_fd_pr__nfet_01v8 ad=0.8151 pd=4.96 as=0.34485 ps=2.42 w=2.09 l=3.35
X14 VDD2.t3 VN.t4 VTAIL.t9 B.t2 sky130_fd_pr__nfet_01v8 ad=0.34485 pd=2.42 as=0.8151 ps=4.96 w=2.09 l=3.35
X15 B.t15 B.t12 B.t14 B.t13 sky130_fd_pr__nfet_01v8 ad=0.8151 pd=4.96 as=0 ps=0 w=2.09 l=3.35
X16 VDD2.t2 VN.t5 VTAIL.t8 B.t0 sky130_fd_pr__nfet_01v8 ad=0.34485 pd=2.42 as=0.34485 ps=2.42 w=2.09 l=3.35
X17 VTAIL.t10 VN.t6 VDD2.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=0.8151 pd=4.96 as=0.34485 ps=2.42 w=2.09 l=3.35
X18 VTAIL.t15 VN.t7 VDD2.t0 B.t3 sky130_fd_pr__nfet_01v8 ad=0.34485 pd=2.42 as=0.34485 ps=2.42 w=2.09 l=3.35
X19 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=0.8151 pd=4.96 as=0 ps=0 w=2.09 l=3.35
R0 B.n616 B.n136 585
R1 B.n136 B.n113 585
R2 B.n618 B.n617 585
R3 B.n620 B.n135 585
R4 B.n623 B.n622 585
R5 B.n624 B.n134 585
R6 B.n626 B.n625 585
R7 B.n628 B.n133 585
R8 B.n631 B.n630 585
R9 B.n632 B.n132 585
R10 B.n634 B.n633 585
R11 B.n636 B.n131 585
R12 B.n638 B.n637 585
R13 B.n640 B.n639 585
R14 B.n643 B.n642 585
R15 B.n644 B.n126 585
R16 B.n646 B.n645 585
R17 B.n648 B.n125 585
R18 B.n651 B.n650 585
R19 B.n652 B.n124 585
R20 B.n654 B.n653 585
R21 B.n656 B.n123 585
R22 B.n659 B.n658 585
R23 B.n661 B.n120 585
R24 B.n663 B.n662 585
R25 B.n665 B.n119 585
R26 B.n668 B.n667 585
R27 B.n669 B.n118 585
R28 B.n671 B.n670 585
R29 B.n673 B.n117 585
R30 B.n676 B.n675 585
R31 B.n677 B.n116 585
R32 B.n679 B.n678 585
R33 B.n681 B.n115 585
R34 B.n684 B.n683 585
R35 B.n685 B.n114 585
R36 B.n615 B.n112 585
R37 B.n688 B.n112 585
R38 B.n614 B.n111 585
R39 B.n689 B.n111 585
R40 B.n613 B.n110 585
R41 B.n690 B.n110 585
R42 B.n612 B.n611 585
R43 B.n611 B.n106 585
R44 B.n610 B.n105 585
R45 B.n696 B.n105 585
R46 B.n609 B.n104 585
R47 B.n697 B.n104 585
R48 B.n608 B.n103 585
R49 B.n698 B.n103 585
R50 B.n607 B.n606 585
R51 B.n606 B.n99 585
R52 B.n605 B.n98 585
R53 B.n704 B.n98 585
R54 B.n604 B.n97 585
R55 B.n705 B.n97 585
R56 B.n603 B.n96 585
R57 B.n706 B.n96 585
R58 B.n602 B.n601 585
R59 B.n601 B.n92 585
R60 B.n600 B.n91 585
R61 B.n712 B.n91 585
R62 B.n599 B.n90 585
R63 B.n713 B.n90 585
R64 B.n598 B.n89 585
R65 B.n714 B.n89 585
R66 B.n597 B.n596 585
R67 B.n596 B.n85 585
R68 B.n595 B.n84 585
R69 B.n720 B.n84 585
R70 B.n594 B.n83 585
R71 B.n721 B.n83 585
R72 B.n593 B.n82 585
R73 B.n722 B.n82 585
R74 B.n592 B.n591 585
R75 B.n591 B.n78 585
R76 B.n590 B.n77 585
R77 B.n728 B.n77 585
R78 B.n589 B.n76 585
R79 B.n729 B.n76 585
R80 B.n588 B.n75 585
R81 B.n730 B.n75 585
R82 B.n587 B.n586 585
R83 B.n586 B.n71 585
R84 B.n585 B.n70 585
R85 B.n736 B.n70 585
R86 B.n584 B.n69 585
R87 B.n737 B.n69 585
R88 B.n583 B.n68 585
R89 B.n738 B.n68 585
R90 B.n582 B.n581 585
R91 B.n581 B.n64 585
R92 B.n580 B.n63 585
R93 B.n744 B.n63 585
R94 B.n579 B.n62 585
R95 B.n745 B.n62 585
R96 B.n578 B.n61 585
R97 B.n746 B.n61 585
R98 B.n577 B.n576 585
R99 B.n576 B.n57 585
R100 B.n575 B.n56 585
R101 B.n752 B.n56 585
R102 B.n574 B.n55 585
R103 B.n753 B.n55 585
R104 B.n573 B.n54 585
R105 B.n754 B.n54 585
R106 B.n572 B.n571 585
R107 B.n571 B.n50 585
R108 B.n570 B.n49 585
R109 B.n760 B.n49 585
R110 B.n569 B.n48 585
R111 B.n761 B.n48 585
R112 B.n568 B.n47 585
R113 B.n762 B.n47 585
R114 B.n567 B.n566 585
R115 B.n566 B.n43 585
R116 B.n565 B.n42 585
R117 B.n768 B.n42 585
R118 B.n564 B.n41 585
R119 B.n769 B.n41 585
R120 B.n563 B.n40 585
R121 B.n770 B.n40 585
R122 B.n562 B.n561 585
R123 B.n561 B.n36 585
R124 B.n560 B.n35 585
R125 B.n776 B.n35 585
R126 B.n559 B.n34 585
R127 B.n777 B.n34 585
R128 B.n558 B.n33 585
R129 B.n778 B.n33 585
R130 B.n557 B.n556 585
R131 B.n556 B.n29 585
R132 B.n555 B.n28 585
R133 B.n784 B.n28 585
R134 B.n554 B.n27 585
R135 B.n785 B.n27 585
R136 B.n553 B.n26 585
R137 B.n786 B.n26 585
R138 B.n552 B.n551 585
R139 B.n551 B.n22 585
R140 B.n550 B.n21 585
R141 B.n792 B.n21 585
R142 B.n549 B.n20 585
R143 B.n793 B.n20 585
R144 B.n548 B.n19 585
R145 B.n794 B.n19 585
R146 B.n547 B.n546 585
R147 B.n546 B.n15 585
R148 B.n545 B.n14 585
R149 B.n800 B.n14 585
R150 B.n544 B.n13 585
R151 B.n801 B.n13 585
R152 B.n543 B.n12 585
R153 B.n802 B.n12 585
R154 B.n542 B.n541 585
R155 B.n541 B.n8 585
R156 B.n540 B.n7 585
R157 B.n808 B.n7 585
R158 B.n539 B.n6 585
R159 B.n809 B.n6 585
R160 B.n538 B.n5 585
R161 B.n810 B.n5 585
R162 B.n537 B.n536 585
R163 B.n536 B.n4 585
R164 B.n535 B.n137 585
R165 B.n535 B.n534 585
R166 B.n525 B.n138 585
R167 B.n139 B.n138 585
R168 B.n527 B.n526 585
R169 B.n528 B.n527 585
R170 B.n524 B.n144 585
R171 B.n144 B.n143 585
R172 B.n523 B.n522 585
R173 B.n522 B.n521 585
R174 B.n146 B.n145 585
R175 B.n147 B.n146 585
R176 B.n514 B.n513 585
R177 B.n515 B.n514 585
R178 B.n512 B.n152 585
R179 B.n152 B.n151 585
R180 B.n511 B.n510 585
R181 B.n510 B.n509 585
R182 B.n154 B.n153 585
R183 B.n155 B.n154 585
R184 B.n502 B.n501 585
R185 B.n503 B.n502 585
R186 B.n500 B.n160 585
R187 B.n160 B.n159 585
R188 B.n499 B.n498 585
R189 B.n498 B.n497 585
R190 B.n162 B.n161 585
R191 B.n163 B.n162 585
R192 B.n490 B.n489 585
R193 B.n491 B.n490 585
R194 B.n488 B.n168 585
R195 B.n168 B.n167 585
R196 B.n487 B.n486 585
R197 B.n486 B.n485 585
R198 B.n170 B.n169 585
R199 B.n171 B.n170 585
R200 B.n478 B.n477 585
R201 B.n479 B.n478 585
R202 B.n476 B.n176 585
R203 B.n176 B.n175 585
R204 B.n475 B.n474 585
R205 B.n474 B.n473 585
R206 B.n178 B.n177 585
R207 B.n179 B.n178 585
R208 B.n466 B.n465 585
R209 B.n467 B.n466 585
R210 B.n464 B.n184 585
R211 B.n184 B.n183 585
R212 B.n463 B.n462 585
R213 B.n462 B.n461 585
R214 B.n186 B.n185 585
R215 B.n187 B.n186 585
R216 B.n454 B.n453 585
R217 B.n455 B.n454 585
R218 B.n452 B.n191 585
R219 B.n195 B.n191 585
R220 B.n451 B.n450 585
R221 B.n450 B.n449 585
R222 B.n193 B.n192 585
R223 B.n194 B.n193 585
R224 B.n442 B.n441 585
R225 B.n443 B.n442 585
R226 B.n440 B.n200 585
R227 B.n200 B.n199 585
R228 B.n439 B.n438 585
R229 B.n438 B.n437 585
R230 B.n202 B.n201 585
R231 B.n203 B.n202 585
R232 B.n430 B.n429 585
R233 B.n431 B.n430 585
R234 B.n428 B.n208 585
R235 B.n208 B.n207 585
R236 B.n427 B.n426 585
R237 B.n426 B.n425 585
R238 B.n210 B.n209 585
R239 B.n211 B.n210 585
R240 B.n418 B.n417 585
R241 B.n419 B.n418 585
R242 B.n416 B.n216 585
R243 B.n216 B.n215 585
R244 B.n415 B.n414 585
R245 B.n414 B.n413 585
R246 B.n218 B.n217 585
R247 B.n219 B.n218 585
R248 B.n406 B.n405 585
R249 B.n407 B.n406 585
R250 B.n404 B.n224 585
R251 B.n224 B.n223 585
R252 B.n403 B.n402 585
R253 B.n402 B.n401 585
R254 B.n226 B.n225 585
R255 B.n227 B.n226 585
R256 B.n394 B.n393 585
R257 B.n395 B.n394 585
R258 B.n392 B.n232 585
R259 B.n232 B.n231 585
R260 B.n391 B.n390 585
R261 B.n390 B.n389 585
R262 B.n234 B.n233 585
R263 B.n235 B.n234 585
R264 B.n382 B.n381 585
R265 B.n383 B.n382 585
R266 B.n380 B.n240 585
R267 B.n240 B.n239 585
R268 B.n379 B.n378 585
R269 B.n378 B.n377 585
R270 B.n242 B.n241 585
R271 B.n243 B.n242 585
R272 B.n370 B.n369 585
R273 B.n371 B.n370 585
R274 B.n368 B.n248 585
R275 B.n248 B.n247 585
R276 B.n367 B.n366 585
R277 B.n366 B.n365 585
R278 B.n250 B.n249 585
R279 B.n251 B.n250 585
R280 B.n358 B.n357 585
R281 B.n359 B.n358 585
R282 B.n356 B.n256 585
R283 B.n256 B.n255 585
R284 B.n355 B.n354 585
R285 B.n354 B.n353 585
R286 B.n350 B.n260 585
R287 B.n349 B.n348 585
R288 B.n346 B.n261 585
R289 B.n346 B.n259 585
R290 B.n345 B.n344 585
R291 B.n343 B.n342 585
R292 B.n341 B.n263 585
R293 B.n339 B.n338 585
R294 B.n337 B.n264 585
R295 B.n336 B.n335 585
R296 B.n333 B.n265 585
R297 B.n331 B.n330 585
R298 B.n329 B.n266 585
R299 B.n328 B.n327 585
R300 B.n325 B.n324 585
R301 B.n323 B.n322 585
R302 B.n321 B.n271 585
R303 B.n319 B.n318 585
R304 B.n317 B.n272 585
R305 B.n316 B.n315 585
R306 B.n313 B.n273 585
R307 B.n311 B.n310 585
R308 B.n309 B.n274 585
R309 B.n307 B.n306 585
R310 B.n304 B.n277 585
R311 B.n302 B.n301 585
R312 B.n300 B.n278 585
R313 B.n299 B.n298 585
R314 B.n296 B.n279 585
R315 B.n294 B.n293 585
R316 B.n292 B.n280 585
R317 B.n291 B.n290 585
R318 B.n288 B.n281 585
R319 B.n286 B.n285 585
R320 B.n284 B.n283 585
R321 B.n258 B.n257 585
R322 B.n352 B.n351 585
R323 B.n353 B.n352 585
R324 B.n254 B.n253 585
R325 B.n255 B.n254 585
R326 B.n361 B.n360 585
R327 B.n360 B.n359 585
R328 B.n362 B.n252 585
R329 B.n252 B.n251 585
R330 B.n364 B.n363 585
R331 B.n365 B.n364 585
R332 B.n246 B.n245 585
R333 B.n247 B.n246 585
R334 B.n373 B.n372 585
R335 B.n372 B.n371 585
R336 B.n374 B.n244 585
R337 B.n244 B.n243 585
R338 B.n376 B.n375 585
R339 B.n377 B.n376 585
R340 B.n238 B.n237 585
R341 B.n239 B.n238 585
R342 B.n385 B.n384 585
R343 B.n384 B.n383 585
R344 B.n386 B.n236 585
R345 B.n236 B.n235 585
R346 B.n388 B.n387 585
R347 B.n389 B.n388 585
R348 B.n230 B.n229 585
R349 B.n231 B.n230 585
R350 B.n397 B.n396 585
R351 B.n396 B.n395 585
R352 B.n398 B.n228 585
R353 B.n228 B.n227 585
R354 B.n400 B.n399 585
R355 B.n401 B.n400 585
R356 B.n222 B.n221 585
R357 B.n223 B.n222 585
R358 B.n409 B.n408 585
R359 B.n408 B.n407 585
R360 B.n410 B.n220 585
R361 B.n220 B.n219 585
R362 B.n412 B.n411 585
R363 B.n413 B.n412 585
R364 B.n214 B.n213 585
R365 B.n215 B.n214 585
R366 B.n421 B.n420 585
R367 B.n420 B.n419 585
R368 B.n422 B.n212 585
R369 B.n212 B.n211 585
R370 B.n424 B.n423 585
R371 B.n425 B.n424 585
R372 B.n206 B.n205 585
R373 B.n207 B.n206 585
R374 B.n433 B.n432 585
R375 B.n432 B.n431 585
R376 B.n434 B.n204 585
R377 B.n204 B.n203 585
R378 B.n436 B.n435 585
R379 B.n437 B.n436 585
R380 B.n198 B.n197 585
R381 B.n199 B.n198 585
R382 B.n445 B.n444 585
R383 B.n444 B.n443 585
R384 B.n446 B.n196 585
R385 B.n196 B.n194 585
R386 B.n448 B.n447 585
R387 B.n449 B.n448 585
R388 B.n190 B.n189 585
R389 B.n195 B.n190 585
R390 B.n457 B.n456 585
R391 B.n456 B.n455 585
R392 B.n458 B.n188 585
R393 B.n188 B.n187 585
R394 B.n460 B.n459 585
R395 B.n461 B.n460 585
R396 B.n182 B.n181 585
R397 B.n183 B.n182 585
R398 B.n469 B.n468 585
R399 B.n468 B.n467 585
R400 B.n470 B.n180 585
R401 B.n180 B.n179 585
R402 B.n472 B.n471 585
R403 B.n473 B.n472 585
R404 B.n174 B.n173 585
R405 B.n175 B.n174 585
R406 B.n481 B.n480 585
R407 B.n480 B.n479 585
R408 B.n482 B.n172 585
R409 B.n172 B.n171 585
R410 B.n484 B.n483 585
R411 B.n485 B.n484 585
R412 B.n166 B.n165 585
R413 B.n167 B.n166 585
R414 B.n493 B.n492 585
R415 B.n492 B.n491 585
R416 B.n494 B.n164 585
R417 B.n164 B.n163 585
R418 B.n496 B.n495 585
R419 B.n497 B.n496 585
R420 B.n158 B.n157 585
R421 B.n159 B.n158 585
R422 B.n505 B.n504 585
R423 B.n504 B.n503 585
R424 B.n506 B.n156 585
R425 B.n156 B.n155 585
R426 B.n508 B.n507 585
R427 B.n509 B.n508 585
R428 B.n150 B.n149 585
R429 B.n151 B.n150 585
R430 B.n517 B.n516 585
R431 B.n516 B.n515 585
R432 B.n518 B.n148 585
R433 B.n148 B.n147 585
R434 B.n520 B.n519 585
R435 B.n521 B.n520 585
R436 B.n142 B.n141 585
R437 B.n143 B.n142 585
R438 B.n530 B.n529 585
R439 B.n529 B.n528 585
R440 B.n531 B.n140 585
R441 B.n140 B.n139 585
R442 B.n533 B.n532 585
R443 B.n534 B.n533 585
R444 B.n2 B.n0 585
R445 B.n4 B.n2 585
R446 B.n3 B.n1 585
R447 B.n809 B.n3 585
R448 B.n807 B.n806 585
R449 B.n808 B.n807 585
R450 B.n805 B.n9 585
R451 B.n9 B.n8 585
R452 B.n804 B.n803 585
R453 B.n803 B.n802 585
R454 B.n11 B.n10 585
R455 B.n801 B.n11 585
R456 B.n799 B.n798 585
R457 B.n800 B.n799 585
R458 B.n797 B.n16 585
R459 B.n16 B.n15 585
R460 B.n796 B.n795 585
R461 B.n795 B.n794 585
R462 B.n18 B.n17 585
R463 B.n793 B.n18 585
R464 B.n791 B.n790 585
R465 B.n792 B.n791 585
R466 B.n789 B.n23 585
R467 B.n23 B.n22 585
R468 B.n788 B.n787 585
R469 B.n787 B.n786 585
R470 B.n25 B.n24 585
R471 B.n785 B.n25 585
R472 B.n783 B.n782 585
R473 B.n784 B.n783 585
R474 B.n781 B.n30 585
R475 B.n30 B.n29 585
R476 B.n780 B.n779 585
R477 B.n779 B.n778 585
R478 B.n32 B.n31 585
R479 B.n777 B.n32 585
R480 B.n775 B.n774 585
R481 B.n776 B.n775 585
R482 B.n773 B.n37 585
R483 B.n37 B.n36 585
R484 B.n772 B.n771 585
R485 B.n771 B.n770 585
R486 B.n39 B.n38 585
R487 B.n769 B.n39 585
R488 B.n767 B.n766 585
R489 B.n768 B.n767 585
R490 B.n765 B.n44 585
R491 B.n44 B.n43 585
R492 B.n764 B.n763 585
R493 B.n763 B.n762 585
R494 B.n46 B.n45 585
R495 B.n761 B.n46 585
R496 B.n759 B.n758 585
R497 B.n760 B.n759 585
R498 B.n757 B.n51 585
R499 B.n51 B.n50 585
R500 B.n756 B.n755 585
R501 B.n755 B.n754 585
R502 B.n53 B.n52 585
R503 B.n753 B.n53 585
R504 B.n751 B.n750 585
R505 B.n752 B.n751 585
R506 B.n749 B.n58 585
R507 B.n58 B.n57 585
R508 B.n748 B.n747 585
R509 B.n747 B.n746 585
R510 B.n60 B.n59 585
R511 B.n745 B.n60 585
R512 B.n743 B.n742 585
R513 B.n744 B.n743 585
R514 B.n741 B.n65 585
R515 B.n65 B.n64 585
R516 B.n740 B.n739 585
R517 B.n739 B.n738 585
R518 B.n67 B.n66 585
R519 B.n737 B.n67 585
R520 B.n735 B.n734 585
R521 B.n736 B.n735 585
R522 B.n733 B.n72 585
R523 B.n72 B.n71 585
R524 B.n732 B.n731 585
R525 B.n731 B.n730 585
R526 B.n74 B.n73 585
R527 B.n729 B.n74 585
R528 B.n727 B.n726 585
R529 B.n728 B.n727 585
R530 B.n725 B.n79 585
R531 B.n79 B.n78 585
R532 B.n724 B.n723 585
R533 B.n723 B.n722 585
R534 B.n81 B.n80 585
R535 B.n721 B.n81 585
R536 B.n719 B.n718 585
R537 B.n720 B.n719 585
R538 B.n717 B.n86 585
R539 B.n86 B.n85 585
R540 B.n716 B.n715 585
R541 B.n715 B.n714 585
R542 B.n88 B.n87 585
R543 B.n713 B.n88 585
R544 B.n711 B.n710 585
R545 B.n712 B.n711 585
R546 B.n709 B.n93 585
R547 B.n93 B.n92 585
R548 B.n708 B.n707 585
R549 B.n707 B.n706 585
R550 B.n95 B.n94 585
R551 B.n705 B.n95 585
R552 B.n703 B.n702 585
R553 B.n704 B.n703 585
R554 B.n701 B.n100 585
R555 B.n100 B.n99 585
R556 B.n700 B.n699 585
R557 B.n699 B.n698 585
R558 B.n102 B.n101 585
R559 B.n697 B.n102 585
R560 B.n695 B.n694 585
R561 B.n696 B.n695 585
R562 B.n693 B.n107 585
R563 B.n107 B.n106 585
R564 B.n692 B.n691 585
R565 B.n691 B.n690 585
R566 B.n109 B.n108 585
R567 B.n689 B.n109 585
R568 B.n687 B.n686 585
R569 B.n688 B.n687 585
R570 B.n812 B.n811 585
R571 B.n811 B.n810 585
R572 B.n352 B.n260 497.305
R573 B.n687 B.n114 497.305
R574 B.n354 B.n258 497.305
R575 B.n136 B.n112 497.305
R576 B.n619 B.n113 256.663
R577 B.n621 B.n113 256.663
R578 B.n627 B.n113 256.663
R579 B.n629 B.n113 256.663
R580 B.n635 B.n113 256.663
R581 B.n130 B.n113 256.663
R582 B.n641 B.n113 256.663
R583 B.n647 B.n113 256.663
R584 B.n649 B.n113 256.663
R585 B.n655 B.n113 256.663
R586 B.n657 B.n113 256.663
R587 B.n664 B.n113 256.663
R588 B.n666 B.n113 256.663
R589 B.n672 B.n113 256.663
R590 B.n674 B.n113 256.663
R591 B.n680 B.n113 256.663
R592 B.n682 B.n113 256.663
R593 B.n347 B.n259 256.663
R594 B.n262 B.n259 256.663
R595 B.n340 B.n259 256.663
R596 B.n334 B.n259 256.663
R597 B.n332 B.n259 256.663
R598 B.n326 B.n259 256.663
R599 B.n270 B.n259 256.663
R600 B.n320 B.n259 256.663
R601 B.n314 B.n259 256.663
R602 B.n312 B.n259 256.663
R603 B.n305 B.n259 256.663
R604 B.n303 B.n259 256.663
R605 B.n297 B.n259 256.663
R606 B.n295 B.n259 256.663
R607 B.n289 B.n259 256.663
R608 B.n287 B.n259 256.663
R609 B.n282 B.n259 256.663
R610 B.n275 B.t8 223.989
R611 B.n267 B.t19 223.989
R612 B.n121 B.t16 223.989
R613 B.n127 B.t12 223.989
R614 B.n353 B.n259 207.605
R615 B.n688 B.n113 207.605
R616 B.n352 B.n254 163.367
R617 B.n360 B.n254 163.367
R618 B.n360 B.n252 163.367
R619 B.n364 B.n252 163.367
R620 B.n364 B.n246 163.367
R621 B.n372 B.n246 163.367
R622 B.n372 B.n244 163.367
R623 B.n376 B.n244 163.367
R624 B.n376 B.n238 163.367
R625 B.n384 B.n238 163.367
R626 B.n384 B.n236 163.367
R627 B.n388 B.n236 163.367
R628 B.n388 B.n230 163.367
R629 B.n396 B.n230 163.367
R630 B.n396 B.n228 163.367
R631 B.n400 B.n228 163.367
R632 B.n400 B.n222 163.367
R633 B.n408 B.n222 163.367
R634 B.n408 B.n220 163.367
R635 B.n412 B.n220 163.367
R636 B.n412 B.n214 163.367
R637 B.n420 B.n214 163.367
R638 B.n420 B.n212 163.367
R639 B.n424 B.n212 163.367
R640 B.n424 B.n206 163.367
R641 B.n432 B.n206 163.367
R642 B.n432 B.n204 163.367
R643 B.n436 B.n204 163.367
R644 B.n436 B.n198 163.367
R645 B.n444 B.n198 163.367
R646 B.n444 B.n196 163.367
R647 B.n448 B.n196 163.367
R648 B.n448 B.n190 163.367
R649 B.n456 B.n190 163.367
R650 B.n456 B.n188 163.367
R651 B.n460 B.n188 163.367
R652 B.n460 B.n182 163.367
R653 B.n468 B.n182 163.367
R654 B.n468 B.n180 163.367
R655 B.n472 B.n180 163.367
R656 B.n472 B.n174 163.367
R657 B.n480 B.n174 163.367
R658 B.n480 B.n172 163.367
R659 B.n484 B.n172 163.367
R660 B.n484 B.n166 163.367
R661 B.n492 B.n166 163.367
R662 B.n492 B.n164 163.367
R663 B.n496 B.n164 163.367
R664 B.n496 B.n158 163.367
R665 B.n504 B.n158 163.367
R666 B.n504 B.n156 163.367
R667 B.n508 B.n156 163.367
R668 B.n508 B.n150 163.367
R669 B.n516 B.n150 163.367
R670 B.n516 B.n148 163.367
R671 B.n520 B.n148 163.367
R672 B.n520 B.n142 163.367
R673 B.n529 B.n142 163.367
R674 B.n529 B.n140 163.367
R675 B.n533 B.n140 163.367
R676 B.n533 B.n2 163.367
R677 B.n811 B.n2 163.367
R678 B.n811 B.n3 163.367
R679 B.n807 B.n3 163.367
R680 B.n807 B.n9 163.367
R681 B.n803 B.n9 163.367
R682 B.n803 B.n11 163.367
R683 B.n799 B.n11 163.367
R684 B.n799 B.n16 163.367
R685 B.n795 B.n16 163.367
R686 B.n795 B.n18 163.367
R687 B.n791 B.n18 163.367
R688 B.n791 B.n23 163.367
R689 B.n787 B.n23 163.367
R690 B.n787 B.n25 163.367
R691 B.n783 B.n25 163.367
R692 B.n783 B.n30 163.367
R693 B.n779 B.n30 163.367
R694 B.n779 B.n32 163.367
R695 B.n775 B.n32 163.367
R696 B.n775 B.n37 163.367
R697 B.n771 B.n37 163.367
R698 B.n771 B.n39 163.367
R699 B.n767 B.n39 163.367
R700 B.n767 B.n44 163.367
R701 B.n763 B.n44 163.367
R702 B.n763 B.n46 163.367
R703 B.n759 B.n46 163.367
R704 B.n759 B.n51 163.367
R705 B.n755 B.n51 163.367
R706 B.n755 B.n53 163.367
R707 B.n751 B.n53 163.367
R708 B.n751 B.n58 163.367
R709 B.n747 B.n58 163.367
R710 B.n747 B.n60 163.367
R711 B.n743 B.n60 163.367
R712 B.n743 B.n65 163.367
R713 B.n739 B.n65 163.367
R714 B.n739 B.n67 163.367
R715 B.n735 B.n67 163.367
R716 B.n735 B.n72 163.367
R717 B.n731 B.n72 163.367
R718 B.n731 B.n74 163.367
R719 B.n727 B.n74 163.367
R720 B.n727 B.n79 163.367
R721 B.n723 B.n79 163.367
R722 B.n723 B.n81 163.367
R723 B.n719 B.n81 163.367
R724 B.n719 B.n86 163.367
R725 B.n715 B.n86 163.367
R726 B.n715 B.n88 163.367
R727 B.n711 B.n88 163.367
R728 B.n711 B.n93 163.367
R729 B.n707 B.n93 163.367
R730 B.n707 B.n95 163.367
R731 B.n703 B.n95 163.367
R732 B.n703 B.n100 163.367
R733 B.n699 B.n100 163.367
R734 B.n699 B.n102 163.367
R735 B.n695 B.n102 163.367
R736 B.n695 B.n107 163.367
R737 B.n691 B.n107 163.367
R738 B.n691 B.n109 163.367
R739 B.n687 B.n109 163.367
R740 B.n348 B.n346 163.367
R741 B.n346 B.n345 163.367
R742 B.n342 B.n341 163.367
R743 B.n339 B.n264 163.367
R744 B.n335 B.n333 163.367
R745 B.n331 B.n266 163.367
R746 B.n327 B.n325 163.367
R747 B.n322 B.n321 163.367
R748 B.n319 B.n272 163.367
R749 B.n315 B.n313 163.367
R750 B.n311 B.n274 163.367
R751 B.n306 B.n304 163.367
R752 B.n302 B.n278 163.367
R753 B.n298 B.n296 163.367
R754 B.n294 B.n280 163.367
R755 B.n290 B.n288 163.367
R756 B.n286 B.n283 163.367
R757 B.n354 B.n256 163.367
R758 B.n358 B.n256 163.367
R759 B.n358 B.n250 163.367
R760 B.n366 B.n250 163.367
R761 B.n366 B.n248 163.367
R762 B.n370 B.n248 163.367
R763 B.n370 B.n242 163.367
R764 B.n378 B.n242 163.367
R765 B.n378 B.n240 163.367
R766 B.n382 B.n240 163.367
R767 B.n382 B.n234 163.367
R768 B.n390 B.n234 163.367
R769 B.n390 B.n232 163.367
R770 B.n394 B.n232 163.367
R771 B.n394 B.n226 163.367
R772 B.n402 B.n226 163.367
R773 B.n402 B.n224 163.367
R774 B.n406 B.n224 163.367
R775 B.n406 B.n218 163.367
R776 B.n414 B.n218 163.367
R777 B.n414 B.n216 163.367
R778 B.n418 B.n216 163.367
R779 B.n418 B.n210 163.367
R780 B.n426 B.n210 163.367
R781 B.n426 B.n208 163.367
R782 B.n430 B.n208 163.367
R783 B.n430 B.n202 163.367
R784 B.n438 B.n202 163.367
R785 B.n438 B.n200 163.367
R786 B.n442 B.n200 163.367
R787 B.n442 B.n193 163.367
R788 B.n450 B.n193 163.367
R789 B.n450 B.n191 163.367
R790 B.n454 B.n191 163.367
R791 B.n454 B.n186 163.367
R792 B.n462 B.n186 163.367
R793 B.n462 B.n184 163.367
R794 B.n466 B.n184 163.367
R795 B.n466 B.n178 163.367
R796 B.n474 B.n178 163.367
R797 B.n474 B.n176 163.367
R798 B.n478 B.n176 163.367
R799 B.n478 B.n170 163.367
R800 B.n486 B.n170 163.367
R801 B.n486 B.n168 163.367
R802 B.n490 B.n168 163.367
R803 B.n490 B.n162 163.367
R804 B.n498 B.n162 163.367
R805 B.n498 B.n160 163.367
R806 B.n502 B.n160 163.367
R807 B.n502 B.n154 163.367
R808 B.n510 B.n154 163.367
R809 B.n510 B.n152 163.367
R810 B.n514 B.n152 163.367
R811 B.n514 B.n146 163.367
R812 B.n522 B.n146 163.367
R813 B.n522 B.n144 163.367
R814 B.n527 B.n144 163.367
R815 B.n527 B.n138 163.367
R816 B.n535 B.n138 163.367
R817 B.n536 B.n535 163.367
R818 B.n536 B.n5 163.367
R819 B.n6 B.n5 163.367
R820 B.n7 B.n6 163.367
R821 B.n541 B.n7 163.367
R822 B.n541 B.n12 163.367
R823 B.n13 B.n12 163.367
R824 B.n14 B.n13 163.367
R825 B.n546 B.n14 163.367
R826 B.n546 B.n19 163.367
R827 B.n20 B.n19 163.367
R828 B.n21 B.n20 163.367
R829 B.n551 B.n21 163.367
R830 B.n551 B.n26 163.367
R831 B.n27 B.n26 163.367
R832 B.n28 B.n27 163.367
R833 B.n556 B.n28 163.367
R834 B.n556 B.n33 163.367
R835 B.n34 B.n33 163.367
R836 B.n35 B.n34 163.367
R837 B.n561 B.n35 163.367
R838 B.n561 B.n40 163.367
R839 B.n41 B.n40 163.367
R840 B.n42 B.n41 163.367
R841 B.n566 B.n42 163.367
R842 B.n566 B.n47 163.367
R843 B.n48 B.n47 163.367
R844 B.n49 B.n48 163.367
R845 B.n571 B.n49 163.367
R846 B.n571 B.n54 163.367
R847 B.n55 B.n54 163.367
R848 B.n56 B.n55 163.367
R849 B.n576 B.n56 163.367
R850 B.n576 B.n61 163.367
R851 B.n62 B.n61 163.367
R852 B.n63 B.n62 163.367
R853 B.n581 B.n63 163.367
R854 B.n581 B.n68 163.367
R855 B.n69 B.n68 163.367
R856 B.n70 B.n69 163.367
R857 B.n586 B.n70 163.367
R858 B.n586 B.n75 163.367
R859 B.n76 B.n75 163.367
R860 B.n77 B.n76 163.367
R861 B.n591 B.n77 163.367
R862 B.n591 B.n82 163.367
R863 B.n83 B.n82 163.367
R864 B.n84 B.n83 163.367
R865 B.n596 B.n84 163.367
R866 B.n596 B.n89 163.367
R867 B.n90 B.n89 163.367
R868 B.n91 B.n90 163.367
R869 B.n601 B.n91 163.367
R870 B.n601 B.n96 163.367
R871 B.n97 B.n96 163.367
R872 B.n98 B.n97 163.367
R873 B.n606 B.n98 163.367
R874 B.n606 B.n103 163.367
R875 B.n104 B.n103 163.367
R876 B.n105 B.n104 163.367
R877 B.n611 B.n105 163.367
R878 B.n611 B.n110 163.367
R879 B.n111 B.n110 163.367
R880 B.n112 B.n111 163.367
R881 B.n683 B.n681 163.367
R882 B.n679 B.n116 163.367
R883 B.n675 B.n673 163.367
R884 B.n671 B.n118 163.367
R885 B.n667 B.n665 163.367
R886 B.n663 B.n120 163.367
R887 B.n658 B.n656 163.367
R888 B.n654 B.n124 163.367
R889 B.n650 B.n648 163.367
R890 B.n646 B.n126 163.367
R891 B.n642 B.n640 163.367
R892 B.n637 B.n636 163.367
R893 B.n634 B.n132 163.367
R894 B.n630 B.n628 163.367
R895 B.n626 B.n134 163.367
R896 B.n622 B.n620 163.367
R897 B.n618 B.n136 163.367
R898 B.n275 B.t11 155.417
R899 B.n127 B.t14 155.417
R900 B.n267 B.t21 155.417
R901 B.n121 B.t17 155.417
R902 B.n353 B.n255 101.561
R903 B.n359 B.n255 101.561
R904 B.n359 B.n251 101.561
R905 B.n365 B.n251 101.561
R906 B.n365 B.n247 101.561
R907 B.n371 B.n247 101.561
R908 B.n371 B.n243 101.561
R909 B.n377 B.n243 101.561
R910 B.n383 B.n239 101.561
R911 B.n383 B.n235 101.561
R912 B.n389 B.n235 101.561
R913 B.n389 B.n231 101.561
R914 B.n395 B.n231 101.561
R915 B.n395 B.n227 101.561
R916 B.n401 B.n227 101.561
R917 B.n401 B.n223 101.561
R918 B.n407 B.n223 101.561
R919 B.n407 B.n219 101.561
R920 B.n413 B.n219 101.561
R921 B.n413 B.n215 101.561
R922 B.n419 B.n215 101.561
R923 B.n425 B.n211 101.561
R924 B.n425 B.n207 101.561
R925 B.n431 B.n207 101.561
R926 B.n431 B.n203 101.561
R927 B.n437 B.n203 101.561
R928 B.n437 B.n199 101.561
R929 B.n443 B.n199 101.561
R930 B.n443 B.n194 101.561
R931 B.n449 B.n194 101.561
R932 B.n449 B.n195 101.561
R933 B.n455 B.n187 101.561
R934 B.n461 B.n187 101.561
R935 B.n461 B.n183 101.561
R936 B.n467 B.n183 101.561
R937 B.n467 B.n179 101.561
R938 B.n473 B.n179 101.561
R939 B.n473 B.n175 101.561
R940 B.n479 B.n175 101.561
R941 B.n479 B.n171 101.561
R942 B.n485 B.n171 101.561
R943 B.n491 B.n167 101.561
R944 B.n491 B.n163 101.561
R945 B.n497 B.n163 101.561
R946 B.n497 B.n159 101.561
R947 B.n503 B.n159 101.561
R948 B.n503 B.n155 101.561
R949 B.n509 B.n155 101.561
R950 B.n509 B.n151 101.561
R951 B.n515 B.n151 101.561
R952 B.n521 B.n147 101.561
R953 B.n521 B.n143 101.561
R954 B.n528 B.n143 101.561
R955 B.n528 B.n139 101.561
R956 B.n534 B.n139 101.561
R957 B.n534 B.n4 101.561
R958 B.n810 B.n4 101.561
R959 B.n810 B.n809 101.561
R960 B.n809 B.n808 101.561
R961 B.n808 B.n8 101.561
R962 B.n802 B.n8 101.561
R963 B.n802 B.n801 101.561
R964 B.n801 B.n800 101.561
R965 B.n800 B.n15 101.561
R966 B.n794 B.n793 101.561
R967 B.n793 B.n792 101.561
R968 B.n792 B.n22 101.561
R969 B.n786 B.n22 101.561
R970 B.n786 B.n785 101.561
R971 B.n785 B.n784 101.561
R972 B.n784 B.n29 101.561
R973 B.n778 B.n29 101.561
R974 B.n778 B.n777 101.561
R975 B.n776 B.n36 101.561
R976 B.n770 B.n36 101.561
R977 B.n770 B.n769 101.561
R978 B.n769 B.n768 101.561
R979 B.n768 B.n43 101.561
R980 B.n762 B.n43 101.561
R981 B.n762 B.n761 101.561
R982 B.n761 B.n760 101.561
R983 B.n760 B.n50 101.561
R984 B.n754 B.n50 101.561
R985 B.n753 B.n752 101.561
R986 B.n752 B.n57 101.561
R987 B.n746 B.n57 101.561
R988 B.n746 B.n745 101.561
R989 B.n745 B.n744 101.561
R990 B.n744 B.n64 101.561
R991 B.n738 B.n64 101.561
R992 B.n738 B.n737 101.561
R993 B.n737 B.n736 101.561
R994 B.n736 B.n71 101.561
R995 B.n730 B.n729 101.561
R996 B.n729 B.n728 101.561
R997 B.n728 B.n78 101.561
R998 B.n722 B.n78 101.561
R999 B.n722 B.n721 101.561
R1000 B.n721 B.n720 101.561
R1001 B.n720 B.n85 101.561
R1002 B.n714 B.n85 101.561
R1003 B.n714 B.n713 101.561
R1004 B.n713 B.n712 101.561
R1005 B.n712 B.n92 101.561
R1006 B.n706 B.n92 101.561
R1007 B.n706 B.n705 101.561
R1008 B.n704 B.n99 101.561
R1009 B.n698 B.n99 101.561
R1010 B.n698 B.n697 101.561
R1011 B.n697 B.n696 101.561
R1012 B.n696 B.n106 101.561
R1013 B.n690 B.n106 101.561
R1014 B.n690 B.n689 101.561
R1015 B.n689 B.n688 101.561
R1016 B.n515 B.t2 100.069
R1017 B.n794 B.t1 100.069
R1018 B.t3 B.n167 85.1329
R1019 B.n777 B.t0 85.1329
R1020 B.n276 B.t10 84.0481
R1021 B.n128 B.t15 84.0481
R1022 B.n268 B.t20 84.0478
R1023 B.n122 B.t18 84.0478
R1024 B.n347 B.n260 71.676
R1025 B.n345 B.n262 71.676
R1026 B.n341 B.n340 71.676
R1027 B.n334 B.n264 71.676
R1028 B.n333 B.n332 71.676
R1029 B.n326 B.n266 71.676
R1030 B.n325 B.n270 71.676
R1031 B.n321 B.n320 71.676
R1032 B.n314 B.n272 71.676
R1033 B.n313 B.n312 71.676
R1034 B.n305 B.n274 71.676
R1035 B.n304 B.n303 71.676
R1036 B.n297 B.n278 71.676
R1037 B.n296 B.n295 71.676
R1038 B.n289 B.n280 71.676
R1039 B.n288 B.n287 71.676
R1040 B.n283 B.n282 71.676
R1041 B.n682 B.n114 71.676
R1042 B.n681 B.n680 71.676
R1043 B.n674 B.n116 71.676
R1044 B.n673 B.n672 71.676
R1045 B.n666 B.n118 71.676
R1046 B.n665 B.n664 71.676
R1047 B.n657 B.n120 71.676
R1048 B.n656 B.n655 71.676
R1049 B.n649 B.n124 71.676
R1050 B.n648 B.n647 71.676
R1051 B.n641 B.n126 71.676
R1052 B.n640 B.n130 71.676
R1053 B.n636 B.n635 71.676
R1054 B.n629 B.n132 71.676
R1055 B.n628 B.n627 71.676
R1056 B.n621 B.n134 71.676
R1057 B.n620 B.n619 71.676
R1058 B.n619 B.n618 71.676
R1059 B.n622 B.n621 71.676
R1060 B.n627 B.n626 71.676
R1061 B.n630 B.n629 71.676
R1062 B.n635 B.n634 71.676
R1063 B.n637 B.n130 71.676
R1064 B.n642 B.n641 71.676
R1065 B.n647 B.n646 71.676
R1066 B.n650 B.n649 71.676
R1067 B.n655 B.n654 71.676
R1068 B.n658 B.n657 71.676
R1069 B.n664 B.n663 71.676
R1070 B.n667 B.n666 71.676
R1071 B.n672 B.n671 71.676
R1072 B.n675 B.n674 71.676
R1073 B.n680 B.n679 71.676
R1074 B.n683 B.n682 71.676
R1075 B.n348 B.n347 71.676
R1076 B.n342 B.n262 71.676
R1077 B.n340 B.n339 71.676
R1078 B.n335 B.n334 71.676
R1079 B.n332 B.n331 71.676
R1080 B.n327 B.n326 71.676
R1081 B.n322 B.n270 71.676
R1082 B.n320 B.n319 71.676
R1083 B.n315 B.n314 71.676
R1084 B.n312 B.n311 71.676
R1085 B.n306 B.n305 71.676
R1086 B.n303 B.n302 71.676
R1087 B.n298 B.n297 71.676
R1088 B.n295 B.n294 71.676
R1089 B.n290 B.n289 71.676
R1090 B.n287 B.n286 71.676
R1091 B.n282 B.n258 71.676
R1092 B.n276 B.n275 71.3702
R1093 B.n268 B.n267 71.3702
R1094 B.n122 B.n121 71.3702
R1095 B.n128 B.n127 71.3702
R1096 B.n455 B.t5 67.2103
R1097 B.n754 B.t7 67.2103
R1098 B.n308 B.n276 59.5399
R1099 B.n269 B.n268 59.5399
R1100 B.n660 B.n122 59.5399
R1101 B.n129 B.n128 59.5399
R1102 B.t9 B.n239 52.2748
R1103 B.n419 B.t6 52.2748
R1104 B.n730 B.t4 52.2748
R1105 B.n705 B.t13 52.2748
R1106 B.n377 B.t9 49.2877
R1107 B.t6 B.n211 49.2877
R1108 B.t4 B.n71 49.2877
R1109 B.t13 B.n704 49.2877
R1110 B.n195 B.t5 34.3522
R1111 B.t7 B.n753 34.3522
R1112 B.n686 B.n685 32.3127
R1113 B.n616 B.n615 32.3127
R1114 B.n355 B.n257 32.3127
R1115 B.n351 B.n350 32.3127
R1116 B B.n812 18.0485
R1117 B.n485 B.t3 16.4296
R1118 B.t0 B.n776 16.4296
R1119 B.n685 B.n684 10.6151
R1120 B.n684 B.n115 10.6151
R1121 B.n678 B.n115 10.6151
R1122 B.n678 B.n677 10.6151
R1123 B.n677 B.n676 10.6151
R1124 B.n676 B.n117 10.6151
R1125 B.n670 B.n117 10.6151
R1126 B.n670 B.n669 10.6151
R1127 B.n669 B.n668 10.6151
R1128 B.n668 B.n119 10.6151
R1129 B.n662 B.n119 10.6151
R1130 B.n662 B.n661 10.6151
R1131 B.n659 B.n123 10.6151
R1132 B.n653 B.n123 10.6151
R1133 B.n653 B.n652 10.6151
R1134 B.n652 B.n651 10.6151
R1135 B.n651 B.n125 10.6151
R1136 B.n645 B.n125 10.6151
R1137 B.n645 B.n644 10.6151
R1138 B.n644 B.n643 10.6151
R1139 B.n639 B.n638 10.6151
R1140 B.n638 B.n131 10.6151
R1141 B.n633 B.n131 10.6151
R1142 B.n633 B.n632 10.6151
R1143 B.n632 B.n631 10.6151
R1144 B.n631 B.n133 10.6151
R1145 B.n625 B.n133 10.6151
R1146 B.n625 B.n624 10.6151
R1147 B.n624 B.n623 10.6151
R1148 B.n623 B.n135 10.6151
R1149 B.n617 B.n135 10.6151
R1150 B.n617 B.n616 10.6151
R1151 B.n356 B.n355 10.6151
R1152 B.n357 B.n356 10.6151
R1153 B.n357 B.n249 10.6151
R1154 B.n367 B.n249 10.6151
R1155 B.n368 B.n367 10.6151
R1156 B.n369 B.n368 10.6151
R1157 B.n369 B.n241 10.6151
R1158 B.n379 B.n241 10.6151
R1159 B.n380 B.n379 10.6151
R1160 B.n381 B.n380 10.6151
R1161 B.n381 B.n233 10.6151
R1162 B.n391 B.n233 10.6151
R1163 B.n392 B.n391 10.6151
R1164 B.n393 B.n392 10.6151
R1165 B.n393 B.n225 10.6151
R1166 B.n403 B.n225 10.6151
R1167 B.n404 B.n403 10.6151
R1168 B.n405 B.n404 10.6151
R1169 B.n405 B.n217 10.6151
R1170 B.n415 B.n217 10.6151
R1171 B.n416 B.n415 10.6151
R1172 B.n417 B.n416 10.6151
R1173 B.n417 B.n209 10.6151
R1174 B.n427 B.n209 10.6151
R1175 B.n428 B.n427 10.6151
R1176 B.n429 B.n428 10.6151
R1177 B.n429 B.n201 10.6151
R1178 B.n439 B.n201 10.6151
R1179 B.n440 B.n439 10.6151
R1180 B.n441 B.n440 10.6151
R1181 B.n441 B.n192 10.6151
R1182 B.n451 B.n192 10.6151
R1183 B.n452 B.n451 10.6151
R1184 B.n453 B.n452 10.6151
R1185 B.n453 B.n185 10.6151
R1186 B.n463 B.n185 10.6151
R1187 B.n464 B.n463 10.6151
R1188 B.n465 B.n464 10.6151
R1189 B.n465 B.n177 10.6151
R1190 B.n475 B.n177 10.6151
R1191 B.n476 B.n475 10.6151
R1192 B.n477 B.n476 10.6151
R1193 B.n477 B.n169 10.6151
R1194 B.n487 B.n169 10.6151
R1195 B.n488 B.n487 10.6151
R1196 B.n489 B.n488 10.6151
R1197 B.n489 B.n161 10.6151
R1198 B.n499 B.n161 10.6151
R1199 B.n500 B.n499 10.6151
R1200 B.n501 B.n500 10.6151
R1201 B.n501 B.n153 10.6151
R1202 B.n511 B.n153 10.6151
R1203 B.n512 B.n511 10.6151
R1204 B.n513 B.n512 10.6151
R1205 B.n513 B.n145 10.6151
R1206 B.n523 B.n145 10.6151
R1207 B.n524 B.n523 10.6151
R1208 B.n526 B.n524 10.6151
R1209 B.n526 B.n525 10.6151
R1210 B.n525 B.n137 10.6151
R1211 B.n537 B.n137 10.6151
R1212 B.n538 B.n537 10.6151
R1213 B.n539 B.n538 10.6151
R1214 B.n540 B.n539 10.6151
R1215 B.n542 B.n540 10.6151
R1216 B.n543 B.n542 10.6151
R1217 B.n544 B.n543 10.6151
R1218 B.n545 B.n544 10.6151
R1219 B.n547 B.n545 10.6151
R1220 B.n548 B.n547 10.6151
R1221 B.n549 B.n548 10.6151
R1222 B.n550 B.n549 10.6151
R1223 B.n552 B.n550 10.6151
R1224 B.n553 B.n552 10.6151
R1225 B.n554 B.n553 10.6151
R1226 B.n555 B.n554 10.6151
R1227 B.n557 B.n555 10.6151
R1228 B.n558 B.n557 10.6151
R1229 B.n559 B.n558 10.6151
R1230 B.n560 B.n559 10.6151
R1231 B.n562 B.n560 10.6151
R1232 B.n563 B.n562 10.6151
R1233 B.n564 B.n563 10.6151
R1234 B.n565 B.n564 10.6151
R1235 B.n567 B.n565 10.6151
R1236 B.n568 B.n567 10.6151
R1237 B.n569 B.n568 10.6151
R1238 B.n570 B.n569 10.6151
R1239 B.n572 B.n570 10.6151
R1240 B.n573 B.n572 10.6151
R1241 B.n574 B.n573 10.6151
R1242 B.n575 B.n574 10.6151
R1243 B.n577 B.n575 10.6151
R1244 B.n578 B.n577 10.6151
R1245 B.n579 B.n578 10.6151
R1246 B.n580 B.n579 10.6151
R1247 B.n582 B.n580 10.6151
R1248 B.n583 B.n582 10.6151
R1249 B.n584 B.n583 10.6151
R1250 B.n585 B.n584 10.6151
R1251 B.n587 B.n585 10.6151
R1252 B.n588 B.n587 10.6151
R1253 B.n589 B.n588 10.6151
R1254 B.n590 B.n589 10.6151
R1255 B.n592 B.n590 10.6151
R1256 B.n593 B.n592 10.6151
R1257 B.n594 B.n593 10.6151
R1258 B.n595 B.n594 10.6151
R1259 B.n597 B.n595 10.6151
R1260 B.n598 B.n597 10.6151
R1261 B.n599 B.n598 10.6151
R1262 B.n600 B.n599 10.6151
R1263 B.n602 B.n600 10.6151
R1264 B.n603 B.n602 10.6151
R1265 B.n604 B.n603 10.6151
R1266 B.n605 B.n604 10.6151
R1267 B.n607 B.n605 10.6151
R1268 B.n608 B.n607 10.6151
R1269 B.n609 B.n608 10.6151
R1270 B.n610 B.n609 10.6151
R1271 B.n612 B.n610 10.6151
R1272 B.n613 B.n612 10.6151
R1273 B.n614 B.n613 10.6151
R1274 B.n615 B.n614 10.6151
R1275 B.n350 B.n349 10.6151
R1276 B.n349 B.n261 10.6151
R1277 B.n344 B.n261 10.6151
R1278 B.n344 B.n343 10.6151
R1279 B.n343 B.n263 10.6151
R1280 B.n338 B.n263 10.6151
R1281 B.n338 B.n337 10.6151
R1282 B.n337 B.n336 10.6151
R1283 B.n336 B.n265 10.6151
R1284 B.n330 B.n265 10.6151
R1285 B.n330 B.n329 10.6151
R1286 B.n329 B.n328 10.6151
R1287 B.n324 B.n323 10.6151
R1288 B.n323 B.n271 10.6151
R1289 B.n318 B.n271 10.6151
R1290 B.n318 B.n317 10.6151
R1291 B.n317 B.n316 10.6151
R1292 B.n316 B.n273 10.6151
R1293 B.n310 B.n273 10.6151
R1294 B.n310 B.n309 10.6151
R1295 B.n307 B.n277 10.6151
R1296 B.n301 B.n277 10.6151
R1297 B.n301 B.n300 10.6151
R1298 B.n300 B.n299 10.6151
R1299 B.n299 B.n279 10.6151
R1300 B.n293 B.n279 10.6151
R1301 B.n293 B.n292 10.6151
R1302 B.n292 B.n291 10.6151
R1303 B.n291 B.n281 10.6151
R1304 B.n285 B.n281 10.6151
R1305 B.n285 B.n284 10.6151
R1306 B.n284 B.n257 10.6151
R1307 B.n351 B.n253 10.6151
R1308 B.n361 B.n253 10.6151
R1309 B.n362 B.n361 10.6151
R1310 B.n363 B.n362 10.6151
R1311 B.n363 B.n245 10.6151
R1312 B.n373 B.n245 10.6151
R1313 B.n374 B.n373 10.6151
R1314 B.n375 B.n374 10.6151
R1315 B.n375 B.n237 10.6151
R1316 B.n385 B.n237 10.6151
R1317 B.n386 B.n385 10.6151
R1318 B.n387 B.n386 10.6151
R1319 B.n387 B.n229 10.6151
R1320 B.n397 B.n229 10.6151
R1321 B.n398 B.n397 10.6151
R1322 B.n399 B.n398 10.6151
R1323 B.n399 B.n221 10.6151
R1324 B.n409 B.n221 10.6151
R1325 B.n410 B.n409 10.6151
R1326 B.n411 B.n410 10.6151
R1327 B.n411 B.n213 10.6151
R1328 B.n421 B.n213 10.6151
R1329 B.n422 B.n421 10.6151
R1330 B.n423 B.n422 10.6151
R1331 B.n423 B.n205 10.6151
R1332 B.n433 B.n205 10.6151
R1333 B.n434 B.n433 10.6151
R1334 B.n435 B.n434 10.6151
R1335 B.n435 B.n197 10.6151
R1336 B.n445 B.n197 10.6151
R1337 B.n446 B.n445 10.6151
R1338 B.n447 B.n446 10.6151
R1339 B.n447 B.n189 10.6151
R1340 B.n457 B.n189 10.6151
R1341 B.n458 B.n457 10.6151
R1342 B.n459 B.n458 10.6151
R1343 B.n459 B.n181 10.6151
R1344 B.n469 B.n181 10.6151
R1345 B.n470 B.n469 10.6151
R1346 B.n471 B.n470 10.6151
R1347 B.n471 B.n173 10.6151
R1348 B.n481 B.n173 10.6151
R1349 B.n482 B.n481 10.6151
R1350 B.n483 B.n482 10.6151
R1351 B.n483 B.n165 10.6151
R1352 B.n493 B.n165 10.6151
R1353 B.n494 B.n493 10.6151
R1354 B.n495 B.n494 10.6151
R1355 B.n495 B.n157 10.6151
R1356 B.n505 B.n157 10.6151
R1357 B.n506 B.n505 10.6151
R1358 B.n507 B.n506 10.6151
R1359 B.n507 B.n149 10.6151
R1360 B.n517 B.n149 10.6151
R1361 B.n518 B.n517 10.6151
R1362 B.n519 B.n518 10.6151
R1363 B.n519 B.n141 10.6151
R1364 B.n530 B.n141 10.6151
R1365 B.n531 B.n530 10.6151
R1366 B.n532 B.n531 10.6151
R1367 B.n532 B.n0 10.6151
R1368 B.n806 B.n1 10.6151
R1369 B.n806 B.n805 10.6151
R1370 B.n805 B.n804 10.6151
R1371 B.n804 B.n10 10.6151
R1372 B.n798 B.n10 10.6151
R1373 B.n798 B.n797 10.6151
R1374 B.n797 B.n796 10.6151
R1375 B.n796 B.n17 10.6151
R1376 B.n790 B.n17 10.6151
R1377 B.n790 B.n789 10.6151
R1378 B.n789 B.n788 10.6151
R1379 B.n788 B.n24 10.6151
R1380 B.n782 B.n24 10.6151
R1381 B.n782 B.n781 10.6151
R1382 B.n781 B.n780 10.6151
R1383 B.n780 B.n31 10.6151
R1384 B.n774 B.n31 10.6151
R1385 B.n774 B.n773 10.6151
R1386 B.n773 B.n772 10.6151
R1387 B.n772 B.n38 10.6151
R1388 B.n766 B.n38 10.6151
R1389 B.n766 B.n765 10.6151
R1390 B.n765 B.n764 10.6151
R1391 B.n764 B.n45 10.6151
R1392 B.n758 B.n45 10.6151
R1393 B.n758 B.n757 10.6151
R1394 B.n757 B.n756 10.6151
R1395 B.n756 B.n52 10.6151
R1396 B.n750 B.n52 10.6151
R1397 B.n750 B.n749 10.6151
R1398 B.n749 B.n748 10.6151
R1399 B.n748 B.n59 10.6151
R1400 B.n742 B.n59 10.6151
R1401 B.n742 B.n741 10.6151
R1402 B.n741 B.n740 10.6151
R1403 B.n740 B.n66 10.6151
R1404 B.n734 B.n66 10.6151
R1405 B.n734 B.n733 10.6151
R1406 B.n733 B.n732 10.6151
R1407 B.n732 B.n73 10.6151
R1408 B.n726 B.n73 10.6151
R1409 B.n726 B.n725 10.6151
R1410 B.n725 B.n724 10.6151
R1411 B.n724 B.n80 10.6151
R1412 B.n718 B.n80 10.6151
R1413 B.n718 B.n717 10.6151
R1414 B.n717 B.n716 10.6151
R1415 B.n716 B.n87 10.6151
R1416 B.n710 B.n87 10.6151
R1417 B.n710 B.n709 10.6151
R1418 B.n709 B.n708 10.6151
R1419 B.n708 B.n94 10.6151
R1420 B.n702 B.n94 10.6151
R1421 B.n702 B.n701 10.6151
R1422 B.n701 B.n700 10.6151
R1423 B.n700 B.n101 10.6151
R1424 B.n694 B.n101 10.6151
R1425 B.n694 B.n693 10.6151
R1426 B.n693 B.n692 10.6151
R1427 B.n692 B.n108 10.6151
R1428 B.n686 B.n108 10.6151
R1429 B.n660 B.n659 6.5566
R1430 B.n643 B.n129 6.5566
R1431 B.n324 B.n269 6.5566
R1432 B.n309 B.n308 6.5566
R1433 B.n661 B.n660 4.05904
R1434 B.n639 B.n129 4.05904
R1435 B.n328 B.n269 4.05904
R1436 B.n308 B.n307 4.05904
R1437 B.n812 B.n0 2.81026
R1438 B.n812 B.n1 2.81026
R1439 B.t2 B.n147 1.49405
R1440 B.t1 B.n15 1.49405
R1441 VN.n68 VN.n67 161.3
R1442 VN.n66 VN.n36 161.3
R1443 VN.n65 VN.n64 161.3
R1444 VN.n63 VN.n37 161.3
R1445 VN.n62 VN.n61 161.3
R1446 VN.n60 VN.n38 161.3
R1447 VN.n59 VN.n58 161.3
R1448 VN.n57 VN.n56 161.3
R1449 VN.n55 VN.n40 161.3
R1450 VN.n54 VN.n53 161.3
R1451 VN.n52 VN.n41 161.3
R1452 VN.n51 VN.n50 161.3
R1453 VN.n49 VN.n42 161.3
R1454 VN.n48 VN.n47 161.3
R1455 VN.n46 VN.n43 161.3
R1456 VN.n33 VN.n32 161.3
R1457 VN.n31 VN.n1 161.3
R1458 VN.n30 VN.n29 161.3
R1459 VN.n28 VN.n2 161.3
R1460 VN.n27 VN.n26 161.3
R1461 VN.n25 VN.n3 161.3
R1462 VN.n24 VN.n23 161.3
R1463 VN.n22 VN.n21 161.3
R1464 VN.n20 VN.n5 161.3
R1465 VN.n19 VN.n18 161.3
R1466 VN.n17 VN.n6 161.3
R1467 VN.n16 VN.n15 161.3
R1468 VN.n14 VN.n7 161.3
R1469 VN.n13 VN.n12 161.3
R1470 VN.n11 VN.n8 161.3
R1471 VN.n34 VN.n0 76.8552
R1472 VN.n69 VN.n35 76.8552
R1473 VN.n10 VN.n9 70.1795
R1474 VN.n45 VN.n44 70.1795
R1475 VN.n15 VN.n6 56.5193
R1476 VN.n50 VN.n41 56.5193
R1477 VN.n45 VN.t4 47.6961
R1478 VN.n10 VN.t6 47.6961
R1479 VN.n26 VN.n2 47.2923
R1480 VN.n61 VN.n37 47.2923
R1481 VN VN.n69 47.1647
R1482 VN.n30 VN.n2 33.6945
R1483 VN.n65 VN.n37 33.6945
R1484 VN.n13 VN.n8 24.4675
R1485 VN.n14 VN.n13 24.4675
R1486 VN.n15 VN.n14 24.4675
R1487 VN.n19 VN.n6 24.4675
R1488 VN.n20 VN.n19 24.4675
R1489 VN.n21 VN.n20 24.4675
R1490 VN.n25 VN.n24 24.4675
R1491 VN.n26 VN.n25 24.4675
R1492 VN.n31 VN.n30 24.4675
R1493 VN.n32 VN.n31 24.4675
R1494 VN.n50 VN.n49 24.4675
R1495 VN.n49 VN.n48 24.4675
R1496 VN.n48 VN.n43 24.4675
R1497 VN.n61 VN.n60 24.4675
R1498 VN.n60 VN.n59 24.4675
R1499 VN.n56 VN.n55 24.4675
R1500 VN.n55 VN.n54 24.4675
R1501 VN.n54 VN.n41 24.4675
R1502 VN.n67 VN.n66 24.4675
R1503 VN.n66 VN.n65 24.4675
R1504 VN.n24 VN.n4 20.0634
R1505 VN.n59 VN.n39 20.0634
R1506 VN.n9 VN.t5 15.036
R1507 VN.n4 VN.t1 15.036
R1508 VN.n0 VN.t0 15.036
R1509 VN.n44 VN.t7 15.036
R1510 VN.n39 VN.t3 15.036
R1511 VN.n35 VN.t2 15.036
R1512 VN.n32 VN.n0 13.2127
R1513 VN.n67 VN.n35 13.2127
R1514 VN.n9 VN.n8 4.40456
R1515 VN.n21 VN.n4 4.40456
R1516 VN.n44 VN.n43 4.40456
R1517 VN.n56 VN.n39 4.40456
R1518 VN.n46 VN.n45 4.24011
R1519 VN.n11 VN.n10 4.24011
R1520 VN.n69 VN.n68 0.354971
R1521 VN.n34 VN.n33 0.354971
R1522 VN VN.n34 0.26696
R1523 VN.n68 VN.n36 0.189894
R1524 VN.n64 VN.n36 0.189894
R1525 VN.n64 VN.n63 0.189894
R1526 VN.n63 VN.n62 0.189894
R1527 VN.n62 VN.n38 0.189894
R1528 VN.n58 VN.n38 0.189894
R1529 VN.n58 VN.n57 0.189894
R1530 VN.n57 VN.n40 0.189894
R1531 VN.n53 VN.n40 0.189894
R1532 VN.n53 VN.n52 0.189894
R1533 VN.n52 VN.n51 0.189894
R1534 VN.n51 VN.n42 0.189894
R1535 VN.n47 VN.n42 0.189894
R1536 VN.n47 VN.n46 0.189894
R1537 VN.n12 VN.n11 0.189894
R1538 VN.n12 VN.n7 0.189894
R1539 VN.n16 VN.n7 0.189894
R1540 VN.n17 VN.n16 0.189894
R1541 VN.n18 VN.n17 0.189894
R1542 VN.n18 VN.n5 0.189894
R1543 VN.n22 VN.n5 0.189894
R1544 VN.n23 VN.n22 0.189894
R1545 VN.n23 VN.n3 0.189894
R1546 VN.n27 VN.n3 0.189894
R1547 VN.n28 VN.n27 0.189894
R1548 VN.n29 VN.n28 0.189894
R1549 VN.n29 VN.n1 0.189894
R1550 VN.n33 VN.n1 0.189894
R1551 VTAIL.n15 VTAIL.t13 84.517
R1552 VTAIL.n2 VTAIL.t10 84.517
R1553 VTAIL.n3 VTAIL.t1 84.517
R1554 VTAIL.n6 VTAIL.t7 84.517
R1555 VTAIL.n14 VTAIL.t0 84.517
R1556 VTAIL.n11 VTAIL.t4 84.5169
R1557 VTAIL.n10 VTAIL.t9 84.5169
R1558 VTAIL.n7 VTAIL.t12 84.5169
R1559 VTAIL.n13 VTAIL.n12 75.0434
R1560 VTAIL.n9 VTAIL.n8 75.0434
R1561 VTAIL.n1 VTAIL.n0 75.0432
R1562 VTAIL.n5 VTAIL.n4 75.0432
R1563 VTAIL.n15 VTAIL.n14 17.341
R1564 VTAIL.n7 VTAIL.n6 17.341
R1565 VTAIL.n0 VTAIL.t8 9.47418
R1566 VTAIL.n0 VTAIL.t11 9.47418
R1567 VTAIL.n4 VTAIL.t6 9.47418
R1568 VTAIL.n4 VTAIL.t5 9.47418
R1569 VTAIL.n12 VTAIL.t2 9.47418
R1570 VTAIL.n12 VTAIL.t3 9.47418
R1571 VTAIL.n8 VTAIL.t14 9.47418
R1572 VTAIL.n8 VTAIL.t15 9.47418
R1573 VTAIL.n9 VTAIL.n7 3.17291
R1574 VTAIL.n10 VTAIL.n9 3.17291
R1575 VTAIL.n13 VTAIL.n11 3.17291
R1576 VTAIL.n14 VTAIL.n13 3.17291
R1577 VTAIL.n6 VTAIL.n5 3.17291
R1578 VTAIL.n5 VTAIL.n3 3.17291
R1579 VTAIL.n2 VTAIL.n1 3.17291
R1580 VTAIL VTAIL.n15 3.11472
R1581 VTAIL.n11 VTAIL.n10 0.470328
R1582 VTAIL.n3 VTAIL.n2 0.470328
R1583 VTAIL VTAIL.n1 0.0586897
R1584 VDD2.n2 VDD2.n1 93.2528
R1585 VDD2.n2 VDD2.n0 93.2528
R1586 VDD2 VDD2.n5 93.2502
R1587 VDD2.n4 VDD2.n3 91.7222
R1588 VDD2.n4 VDD2.n2 39.7929
R1589 VDD2.n5 VDD2.t0 9.47418
R1590 VDD2.n5 VDD2.t3 9.47418
R1591 VDD2.n3 VDD2.t5 9.47418
R1592 VDD2.n3 VDD2.t4 9.47418
R1593 VDD2.n1 VDD2.t6 9.47418
R1594 VDD2.n1 VDD2.t7 9.47418
R1595 VDD2.n0 VDD2.t1 9.47418
R1596 VDD2.n0 VDD2.t2 9.47418
R1597 VDD2 VDD2.n4 1.6449
R1598 VP.n24 VP.n21 161.3
R1599 VP.n26 VP.n25 161.3
R1600 VP.n27 VP.n20 161.3
R1601 VP.n29 VP.n28 161.3
R1602 VP.n30 VP.n19 161.3
R1603 VP.n32 VP.n31 161.3
R1604 VP.n33 VP.n18 161.3
R1605 VP.n35 VP.n34 161.3
R1606 VP.n37 VP.n36 161.3
R1607 VP.n38 VP.n16 161.3
R1608 VP.n40 VP.n39 161.3
R1609 VP.n41 VP.n15 161.3
R1610 VP.n43 VP.n42 161.3
R1611 VP.n44 VP.n14 161.3
R1612 VP.n46 VP.n45 161.3
R1613 VP.n83 VP.n82 161.3
R1614 VP.n81 VP.n1 161.3
R1615 VP.n80 VP.n79 161.3
R1616 VP.n78 VP.n2 161.3
R1617 VP.n77 VP.n76 161.3
R1618 VP.n75 VP.n3 161.3
R1619 VP.n74 VP.n73 161.3
R1620 VP.n72 VP.n71 161.3
R1621 VP.n70 VP.n5 161.3
R1622 VP.n69 VP.n68 161.3
R1623 VP.n67 VP.n6 161.3
R1624 VP.n66 VP.n65 161.3
R1625 VP.n64 VP.n7 161.3
R1626 VP.n63 VP.n62 161.3
R1627 VP.n61 VP.n8 161.3
R1628 VP.n60 VP.n59 161.3
R1629 VP.n57 VP.n9 161.3
R1630 VP.n56 VP.n55 161.3
R1631 VP.n54 VP.n10 161.3
R1632 VP.n53 VP.n52 161.3
R1633 VP.n51 VP.n11 161.3
R1634 VP.n50 VP.n49 161.3
R1635 VP.n48 VP.n12 76.8552
R1636 VP.n84 VP.n0 76.8552
R1637 VP.n47 VP.n13 76.8552
R1638 VP.n23 VP.n22 70.1795
R1639 VP.n65 VP.n6 56.5193
R1640 VP.n28 VP.n19 56.5193
R1641 VP.n23 VP.t1 47.6959
R1642 VP.n56 VP.n10 47.2923
R1643 VP.n76 VP.n2 47.2923
R1644 VP.n39 VP.n15 47.2923
R1645 VP.n48 VP.n47 46.9993
R1646 VP.n52 VP.n10 33.6945
R1647 VP.n80 VP.n2 33.6945
R1648 VP.n43 VP.n15 33.6945
R1649 VP.n51 VP.n50 24.4675
R1650 VP.n52 VP.n51 24.4675
R1651 VP.n57 VP.n56 24.4675
R1652 VP.n59 VP.n57 24.4675
R1653 VP.n63 VP.n8 24.4675
R1654 VP.n64 VP.n63 24.4675
R1655 VP.n65 VP.n64 24.4675
R1656 VP.n69 VP.n6 24.4675
R1657 VP.n70 VP.n69 24.4675
R1658 VP.n71 VP.n70 24.4675
R1659 VP.n75 VP.n74 24.4675
R1660 VP.n76 VP.n75 24.4675
R1661 VP.n81 VP.n80 24.4675
R1662 VP.n82 VP.n81 24.4675
R1663 VP.n44 VP.n43 24.4675
R1664 VP.n45 VP.n44 24.4675
R1665 VP.n32 VP.n19 24.4675
R1666 VP.n33 VP.n32 24.4675
R1667 VP.n34 VP.n33 24.4675
R1668 VP.n38 VP.n37 24.4675
R1669 VP.n39 VP.n38 24.4675
R1670 VP.n26 VP.n21 24.4675
R1671 VP.n27 VP.n26 24.4675
R1672 VP.n28 VP.n27 24.4675
R1673 VP.n59 VP.n58 20.0634
R1674 VP.n74 VP.n4 20.0634
R1675 VP.n37 VP.n17 20.0634
R1676 VP.n12 VP.t7 15.036
R1677 VP.n58 VP.t0 15.036
R1678 VP.n4 VP.t3 15.036
R1679 VP.n0 VP.t5 15.036
R1680 VP.n13 VP.t6 15.036
R1681 VP.n17 VP.t2 15.036
R1682 VP.n22 VP.t4 15.036
R1683 VP.n50 VP.n12 13.2127
R1684 VP.n82 VP.n0 13.2127
R1685 VP.n45 VP.n13 13.2127
R1686 VP.n58 VP.n8 4.40456
R1687 VP.n71 VP.n4 4.40456
R1688 VP.n34 VP.n17 4.40456
R1689 VP.n22 VP.n21 4.40456
R1690 VP.n24 VP.n23 4.24008
R1691 VP.n47 VP.n46 0.354971
R1692 VP.n49 VP.n48 0.354971
R1693 VP.n84 VP.n83 0.354971
R1694 VP VP.n84 0.26696
R1695 VP.n25 VP.n24 0.189894
R1696 VP.n25 VP.n20 0.189894
R1697 VP.n29 VP.n20 0.189894
R1698 VP.n30 VP.n29 0.189894
R1699 VP.n31 VP.n30 0.189894
R1700 VP.n31 VP.n18 0.189894
R1701 VP.n35 VP.n18 0.189894
R1702 VP.n36 VP.n35 0.189894
R1703 VP.n36 VP.n16 0.189894
R1704 VP.n40 VP.n16 0.189894
R1705 VP.n41 VP.n40 0.189894
R1706 VP.n42 VP.n41 0.189894
R1707 VP.n42 VP.n14 0.189894
R1708 VP.n46 VP.n14 0.189894
R1709 VP.n49 VP.n11 0.189894
R1710 VP.n53 VP.n11 0.189894
R1711 VP.n54 VP.n53 0.189894
R1712 VP.n55 VP.n54 0.189894
R1713 VP.n55 VP.n9 0.189894
R1714 VP.n60 VP.n9 0.189894
R1715 VP.n61 VP.n60 0.189894
R1716 VP.n62 VP.n61 0.189894
R1717 VP.n62 VP.n7 0.189894
R1718 VP.n66 VP.n7 0.189894
R1719 VP.n67 VP.n66 0.189894
R1720 VP.n68 VP.n67 0.189894
R1721 VP.n68 VP.n5 0.189894
R1722 VP.n72 VP.n5 0.189894
R1723 VP.n73 VP.n72 0.189894
R1724 VP.n73 VP.n3 0.189894
R1725 VP.n77 VP.n3 0.189894
R1726 VP.n78 VP.n77 0.189894
R1727 VP.n79 VP.n78 0.189894
R1728 VP.n79 VP.n1 0.189894
R1729 VP.n83 VP.n1 0.189894
R1730 VDD1 VDD1.n0 93.3666
R1731 VDD1.n3 VDD1.n2 93.2528
R1732 VDD1.n3 VDD1.n1 93.2528
R1733 VDD1.n5 VDD1.n4 91.7222
R1734 VDD1.n5 VDD1.n3 40.3759
R1735 VDD1.n4 VDD1.t5 9.47418
R1736 VDD1.n4 VDD1.t1 9.47418
R1737 VDD1.n0 VDD1.t6 9.47418
R1738 VDD1.n0 VDD1.t3 9.47418
R1739 VDD1.n2 VDD1.t4 9.47418
R1740 VDD1.n2 VDD1.t2 9.47418
R1741 VDD1.n1 VDD1.t0 9.47418
R1742 VDD1.n1 VDD1.t7 9.47418
R1743 VDD1 VDD1.n5 1.52852
C0 VN VP 6.7534f
C1 VTAIL VP 3.43929f
C2 VDD1 VP 2.4241f
C3 VDD2 VP 0.606296f
C4 VTAIL VN 3.42518f
C5 VDD1 VN 0.158595f
C6 VDD2 VN 1.97983f
C7 VDD1 VTAIL 5.42783f
C8 VDD2 VTAIL 5.48728f
C9 VDD2 VDD1 2.16395f
C10 VDD2 B 5.28014f
C11 VDD1 B 6.01702f
C12 VTAIL B 4.486934f
C13 VN B 17.430628f
C14 VP B 16.075586f
C15 VDD1.t6 B 0.0526f
C16 VDD1.t3 B 0.0526f
C17 VDD1.n0 B 0.369402f
C18 VDD1.t0 B 0.0526f
C19 VDD1.t7 B 0.0526f
C20 VDD1.n1 B 0.368342f
C21 VDD1.t4 B 0.0526f
C22 VDD1.t2 B 0.0526f
C23 VDD1.n2 B 0.368342f
C24 VDD1.n3 B 3.95594f
C25 VDD1.t5 B 0.0526f
C26 VDD1.t1 B 0.0526f
C27 VDD1.n4 B 0.356505f
C28 VDD1.n5 B 3.11585f
C29 VP.t5 B 0.472899f
C30 VP.n0 B 0.325663f
C31 VP.n1 B 0.028674f
C32 VP.n2 B 0.025037f
C33 VP.n3 B 0.028674f
C34 VP.t3 B 0.472899f
C35 VP.n4 B 0.213929f
C36 VP.n5 B 0.028674f
C37 VP.n6 B 0.041859f
C38 VP.n7 B 0.028674f
C39 VP.n8 B 0.031807f
C40 VP.n9 B 0.028674f
C41 VP.n10 B 0.025037f
C42 VP.n11 B 0.028674f
C43 VP.t7 B 0.472899f
C44 VP.n12 B 0.325663f
C45 VP.t6 B 0.472899f
C46 VP.n13 B 0.325663f
C47 VP.n14 B 0.028674f
C48 VP.n15 B 0.025037f
C49 VP.n16 B 0.028674f
C50 VP.t2 B 0.472899f
C51 VP.n17 B 0.213929f
C52 VP.n18 B 0.028674f
C53 VP.n19 B 0.041859f
C54 VP.n20 B 0.028674f
C55 VP.n21 B 0.031807f
C56 VP.t1 B 0.759842f
C57 VP.t4 B 0.472899f
C58 VP.n22 B 0.303048f
C59 VP.n23 B 0.321303f
C60 VP.n24 B 0.339575f
C61 VP.n25 B 0.028674f
C62 VP.n26 B 0.053442f
C63 VP.n27 B 0.053442f
C64 VP.n28 B 0.041859f
C65 VP.n29 B 0.028674f
C66 VP.n30 B 0.028674f
C67 VP.n31 B 0.028674f
C68 VP.n32 B 0.053442f
C69 VP.n33 B 0.053442f
C70 VP.n34 B 0.031807f
C71 VP.n35 B 0.028674f
C72 VP.n36 B 0.028674f
C73 VP.n37 B 0.048693f
C74 VP.n38 B 0.053442f
C75 VP.n39 B 0.054203f
C76 VP.n40 B 0.028674f
C77 VP.n41 B 0.028674f
C78 VP.n42 B 0.028674f
C79 VP.n43 B 0.05792f
C80 VP.n44 B 0.053442f
C81 VP.n45 B 0.041305f
C82 VP.n46 B 0.04628f
C83 VP.n47 B 1.49279f
C84 VP.n48 B 1.51472f
C85 VP.n49 B 0.04628f
C86 VP.n50 B 0.041305f
C87 VP.n51 B 0.053442f
C88 VP.n52 B 0.05792f
C89 VP.n53 B 0.028674f
C90 VP.n54 B 0.028674f
C91 VP.n55 B 0.028674f
C92 VP.n56 B 0.054203f
C93 VP.n57 B 0.053442f
C94 VP.t0 B 0.472899f
C95 VP.n58 B 0.213929f
C96 VP.n59 B 0.048693f
C97 VP.n60 B 0.028674f
C98 VP.n61 B 0.028674f
C99 VP.n62 B 0.028674f
C100 VP.n63 B 0.053442f
C101 VP.n64 B 0.053442f
C102 VP.n65 B 0.041859f
C103 VP.n66 B 0.028674f
C104 VP.n67 B 0.028674f
C105 VP.n68 B 0.028674f
C106 VP.n69 B 0.053442f
C107 VP.n70 B 0.053442f
C108 VP.n71 B 0.031807f
C109 VP.n72 B 0.028674f
C110 VP.n73 B 0.028674f
C111 VP.n74 B 0.048693f
C112 VP.n75 B 0.053442f
C113 VP.n76 B 0.054203f
C114 VP.n77 B 0.028674f
C115 VP.n78 B 0.028674f
C116 VP.n79 B 0.028674f
C117 VP.n80 B 0.05792f
C118 VP.n81 B 0.053442f
C119 VP.n82 B 0.041305f
C120 VP.n83 B 0.04628f
C121 VP.n84 B 0.07165f
C122 VDD2.t1 B 0.040984f
C123 VDD2.t2 B 0.040984f
C124 VDD2.n0 B 0.286999f
C125 VDD2.t6 B 0.040984f
C126 VDD2.t7 B 0.040984f
C127 VDD2.n1 B 0.286999f
C128 VDD2.n2 B 3.03084f
C129 VDD2.t5 B 0.040984f
C130 VDD2.t4 B 0.040984f
C131 VDD2.n3 B 0.277778f
C132 VDD2.n4 B 2.3969f
C133 VDD2.t0 B 0.040984f
C134 VDD2.t3 B 0.040984f
C135 VDD2.n5 B 0.286972f
C136 VTAIL.t8 B 0.054124f
C137 VTAIL.t11 B 0.054124f
C138 VTAIL.n0 B 0.316762f
C139 VTAIL.n1 B 0.578222f
C140 VTAIL.t10 B 0.418387f
C141 VTAIL.n2 B 0.667676f
C142 VTAIL.t1 B 0.418387f
C143 VTAIL.n3 B 0.667676f
C144 VTAIL.t6 B 0.054124f
C145 VTAIL.t5 B 0.054124f
C146 VTAIL.n4 B 0.316762f
C147 VTAIL.n5 B 0.907071f
C148 VTAIL.t7 B 0.418387f
C149 VTAIL.n6 B 1.58847f
C150 VTAIL.t12 B 0.418389f
C151 VTAIL.n7 B 1.58847f
C152 VTAIL.t14 B 0.054124f
C153 VTAIL.t15 B 0.054124f
C154 VTAIL.n8 B 0.316763f
C155 VTAIL.n9 B 0.90707f
C156 VTAIL.t9 B 0.418389f
C157 VTAIL.n10 B 0.667673f
C158 VTAIL.t4 B 0.418389f
C159 VTAIL.n11 B 0.667673f
C160 VTAIL.t2 B 0.054124f
C161 VTAIL.t3 B 0.054124f
C162 VTAIL.n12 B 0.316763f
C163 VTAIL.n13 B 0.90707f
C164 VTAIL.t0 B 0.418387f
C165 VTAIL.n14 B 1.58847f
C166 VTAIL.t13 B 0.418387f
C167 VTAIL.n15 B 1.58233f
C168 VN.t0 B 0.381602f
C169 VN.n0 B 0.262791f
C170 VN.n1 B 0.023139f
C171 VN.n2 B 0.020204f
C172 VN.n3 B 0.023139f
C173 VN.t1 B 0.381602f
C174 VN.n4 B 0.172628f
C175 VN.n5 B 0.023139f
C176 VN.n6 B 0.033778f
C177 VN.n7 B 0.023139f
C178 VN.n8 B 0.025666f
C179 VN.t5 B 0.381602f
C180 VN.n9 B 0.244542f
C181 VN.t6 B 0.61315f
C182 VN.n10 B 0.259273f
C183 VN.n11 B 0.274017f
C184 VN.n12 B 0.023139f
C185 VN.n13 B 0.043124f
C186 VN.n14 B 0.043124f
C187 VN.n15 B 0.033778f
C188 VN.n16 B 0.023139f
C189 VN.n17 B 0.023139f
C190 VN.n18 B 0.023139f
C191 VN.n19 B 0.043124f
C192 VN.n20 B 0.043124f
C193 VN.n21 B 0.025666f
C194 VN.n22 B 0.023139f
C195 VN.n23 B 0.023139f
C196 VN.n24 B 0.039292f
C197 VN.n25 B 0.043124f
C198 VN.n26 B 0.043739f
C199 VN.n27 B 0.023139f
C200 VN.n28 B 0.023139f
C201 VN.n29 B 0.023139f
C202 VN.n30 B 0.046738f
C203 VN.n31 B 0.043124f
C204 VN.n32 B 0.033331f
C205 VN.n33 B 0.037345f
C206 VN.n34 B 0.057818f
C207 VN.t2 B 0.381602f
C208 VN.n35 B 0.262791f
C209 VN.n36 B 0.023139f
C210 VN.n37 B 0.020204f
C211 VN.n38 B 0.023139f
C212 VN.t3 B 0.381602f
C213 VN.n39 B 0.172628f
C214 VN.n40 B 0.023139f
C215 VN.n41 B 0.033778f
C216 VN.n42 B 0.023139f
C217 VN.n43 B 0.025666f
C218 VN.t4 B 0.61315f
C219 VN.t7 B 0.381602f
C220 VN.n44 B 0.244542f
C221 VN.n45 B 0.259273f
C222 VN.n46 B 0.274017f
C223 VN.n47 B 0.023139f
C224 VN.n48 B 0.043124f
C225 VN.n49 B 0.043124f
C226 VN.n50 B 0.033778f
C227 VN.n51 B 0.023139f
C228 VN.n52 B 0.023139f
C229 VN.n53 B 0.023139f
C230 VN.n54 B 0.043124f
C231 VN.n55 B 0.043124f
C232 VN.n56 B 0.025666f
C233 VN.n57 B 0.023139f
C234 VN.n58 B 0.023139f
C235 VN.n59 B 0.039292f
C236 VN.n60 B 0.043124f
C237 VN.n61 B 0.043739f
C238 VN.n62 B 0.023139f
C239 VN.n63 B 0.023139f
C240 VN.n64 B 0.023139f
C241 VN.n65 B 0.046738f
C242 VN.n66 B 0.043124f
C243 VN.n67 B 0.033331f
C244 VN.n68 B 0.037345f
C245 VN.n69 B 1.21427f
.ends

