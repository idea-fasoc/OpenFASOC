* NGSPICE file created from diff_pair_sample_1486.ext - technology: sky130A

.subckt diff_pair_sample_1486 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t15 VP.t0 VDD1.t7 B.t3 sky130_fd_pr__nfet_01v8 ad=2.7423 pd=16.95 as=2.7423 ps=16.95 w=16.62 l=1.97
X1 VTAIL.t2 VN.t0 VDD2.t7 B.t2 sky130_fd_pr__nfet_01v8 ad=6.4818 pd=34.02 as=2.7423 ps=16.95 w=16.62 l=1.97
X2 B.t21 B.t19 B.t20 B.t16 sky130_fd_pr__nfet_01v8 ad=6.4818 pd=34.02 as=0 ps=0 w=16.62 l=1.97
X3 VDD2.t6 VN.t1 VTAIL.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=2.7423 pd=16.95 as=2.7423 ps=16.95 w=16.62 l=1.97
X4 B.t18 B.t15 B.t17 B.t16 sky130_fd_pr__nfet_01v8 ad=6.4818 pd=34.02 as=0 ps=0 w=16.62 l=1.97
X5 VDD2.t5 VN.t2 VTAIL.t7 B.t7 sky130_fd_pr__nfet_01v8 ad=2.7423 pd=16.95 as=6.4818 ps=34.02 w=16.62 l=1.97
X6 VTAIL.t5 VN.t3 VDD2.t4 B.t5 sky130_fd_pr__nfet_01v8 ad=2.7423 pd=16.95 as=2.7423 ps=16.95 w=16.62 l=1.97
X7 VTAIL.t14 VP.t1 VDD1.t6 B.t1 sky130_fd_pr__nfet_01v8 ad=6.4818 pd=34.02 as=2.7423 ps=16.95 w=16.62 l=1.97
X8 B.t14 B.t12 B.t13 B.t9 sky130_fd_pr__nfet_01v8 ad=6.4818 pd=34.02 as=0 ps=0 w=16.62 l=1.97
X9 VTAIL.t13 VP.t2 VDD1.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=2.7423 pd=16.95 as=2.7423 ps=16.95 w=16.62 l=1.97
X10 VDD1.t4 VP.t3 VTAIL.t12 B.t6 sky130_fd_pr__nfet_01v8 ad=2.7423 pd=16.95 as=2.7423 ps=16.95 w=16.62 l=1.97
X11 VDD2.t3 VN.t4 VTAIL.t6 B.t6 sky130_fd_pr__nfet_01v8 ad=2.7423 pd=16.95 as=2.7423 ps=16.95 w=16.62 l=1.97
X12 VDD1.t1 VP.t4 VTAIL.t11 B.t7 sky130_fd_pr__nfet_01v8 ad=2.7423 pd=16.95 as=6.4818 ps=34.02 w=16.62 l=1.97
X13 VDD1.t0 VP.t5 VTAIL.t10 B.t4 sky130_fd_pr__nfet_01v8 ad=2.7423 pd=16.95 as=2.7423 ps=16.95 w=16.62 l=1.97
X14 VTAIL.t3 VN.t5 VDD2.t2 B.t3 sky130_fd_pr__nfet_01v8 ad=2.7423 pd=16.95 as=2.7423 ps=16.95 w=16.62 l=1.97
X15 VDD2.t1 VN.t6 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=2.7423 pd=16.95 as=6.4818 ps=34.02 w=16.62 l=1.97
X16 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=6.4818 pd=34.02 as=0 ps=0 w=16.62 l=1.97
X17 VTAIL.t1 VN.t7 VDD2.t0 B.t1 sky130_fd_pr__nfet_01v8 ad=6.4818 pd=34.02 as=2.7423 ps=16.95 w=16.62 l=1.97
X18 VDD1.t3 VP.t6 VTAIL.t9 B.t0 sky130_fd_pr__nfet_01v8 ad=2.7423 pd=16.95 as=6.4818 ps=34.02 w=16.62 l=1.97
X19 VTAIL.t8 VP.t7 VDD1.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=6.4818 pd=34.02 as=2.7423 ps=16.95 w=16.62 l=1.97
R0 VP.n12 VP.t1 234.126
R1 VP.n31 VP.t7 203.321
R2 VP.n38 VP.t3 203.321
R3 VP.n46 VP.t2 203.321
R4 VP.n53 VP.t6 203.321
R5 VP.n28 VP.t4 203.321
R6 VP.n21 VP.t0 203.321
R7 VP.n13 VP.t5 203.321
R8 VP.n14 VP.n11 161.3
R9 VP.n16 VP.n15 161.3
R10 VP.n17 VP.n10 161.3
R11 VP.n19 VP.n18 161.3
R12 VP.n20 VP.n9 161.3
R13 VP.n23 VP.n22 161.3
R14 VP.n24 VP.n8 161.3
R15 VP.n26 VP.n25 161.3
R16 VP.n27 VP.n7 161.3
R17 VP.n52 VP.n0 161.3
R18 VP.n51 VP.n50 161.3
R19 VP.n49 VP.n1 161.3
R20 VP.n48 VP.n47 161.3
R21 VP.n45 VP.n2 161.3
R22 VP.n44 VP.n43 161.3
R23 VP.n42 VP.n3 161.3
R24 VP.n41 VP.n40 161.3
R25 VP.n39 VP.n4 161.3
R26 VP.n37 VP.n36 161.3
R27 VP.n35 VP.n5 161.3
R28 VP.n34 VP.n33 161.3
R29 VP.n32 VP.n6 161.3
R30 VP.n31 VP.n30 88.7756
R31 VP.n54 VP.n53 88.7756
R32 VP.n29 VP.n28 88.7756
R33 VP.n13 VP.n12 62.9301
R34 VP.n33 VP.n5 56.5617
R35 VP.n51 VP.n1 56.5617
R36 VP.n26 VP.n8 56.5617
R37 VP.n30 VP.n29 51.4997
R38 VP.n40 VP.n3 40.577
R39 VP.n44 VP.n3 40.577
R40 VP.n19 VP.n10 40.577
R41 VP.n15 VP.n10 40.577
R42 VP.n33 VP.n32 24.5923
R43 VP.n37 VP.n5 24.5923
R44 VP.n40 VP.n39 24.5923
R45 VP.n45 VP.n44 24.5923
R46 VP.n47 VP.n1 24.5923
R47 VP.n52 VP.n51 24.5923
R48 VP.n27 VP.n26 24.5923
R49 VP.n20 VP.n19 24.5923
R50 VP.n22 VP.n8 24.5923
R51 VP.n15 VP.n14 24.5923
R52 VP.n32 VP.n31 22.1332
R53 VP.n53 VP.n52 22.1332
R54 VP.n28 VP.n27 22.1332
R55 VP.n38 VP.n37 17.2148
R56 VP.n47 VP.n46 17.2148
R57 VP.n22 VP.n21 17.2148
R58 VP.n12 VP.n11 12.9948
R59 VP.n39 VP.n38 7.37805
R60 VP.n46 VP.n45 7.37805
R61 VP.n21 VP.n20 7.37805
R62 VP.n14 VP.n13 7.37805
R63 VP.n29 VP.n7 0.278335
R64 VP.n30 VP.n6 0.278335
R65 VP.n54 VP.n0 0.278335
R66 VP.n16 VP.n11 0.189894
R67 VP.n17 VP.n16 0.189894
R68 VP.n18 VP.n17 0.189894
R69 VP.n18 VP.n9 0.189894
R70 VP.n23 VP.n9 0.189894
R71 VP.n24 VP.n23 0.189894
R72 VP.n25 VP.n24 0.189894
R73 VP.n25 VP.n7 0.189894
R74 VP.n34 VP.n6 0.189894
R75 VP.n35 VP.n34 0.189894
R76 VP.n36 VP.n35 0.189894
R77 VP.n36 VP.n4 0.189894
R78 VP.n41 VP.n4 0.189894
R79 VP.n42 VP.n41 0.189894
R80 VP.n43 VP.n42 0.189894
R81 VP.n43 VP.n2 0.189894
R82 VP.n48 VP.n2 0.189894
R83 VP.n49 VP.n48 0.189894
R84 VP.n50 VP.n49 0.189894
R85 VP.n50 VP.n0 0.189894
R86 VP VP.n54 0.153485
R87 VDD1 VDD1.n0 65.2901
R88 VDD1.n3 VDD1.n2 65.1763
R89 VDD1.n3 VDD1.n1 65.1763
R90 VDD1.n5 VDD1.n4 64.2404
R91 VDD1.n5 VDD1.n3 47.5483
R92 VDD1.n4 VDD1.t7 1.19184
R93 VDD1.n4 VDD1.t1 1.19184
R94 VDD1.n0 VDD1.t6 1.19184
R95 VDD1.n0 VDD1.t0 1.19184
R96 VDD1.n2 VDD1.t5 1.19184
R97 VDD1.n2 VDD1.t3 1.19184
R98 VDD1.n1 VDD1.t2 1.19184
R99 VDD1.n1 VDD1.t4 1.19184
R100 VDD1 VDD1.n5 0.93369
R101 VTAIL.n11 VTAIL.t14 48.7531
R102 VTAIL.n10 VTAIL.t0 48.7531
R103 VTAIL.n7 VTAIL.t2 48.7531
R104 VTAIL.n14 VTAIL.t11 48.7529
R105 VTAIL.n15 VTAIL.t7 48.7529
R106 VTAIL.n2 VTAIL.t1 48.7529
R107 VTAIL.n3 VTAIL.t9 48.7529
R108 VTAIL.n6 VTAIL.t8 48.7529
R109 VTAIL.n13 VTAIL.n12 47.5618
R110 VTAIL.n9 VTAIL.n8 47.5618
R111 VTAIL.n1 VTAIL.n0 47.5615
R112 VTAIL.n5 VTAIL.n4 47.5615
R113 VTAIL.n15 VTAIL.n14 28.6772
R114 VTAIL.n7 VTAIL.n6 28.6772
R115 VTAIL.n9 VTAIL.n7 1.98326
R116 VTAIL.n10 VTAIL.n9 1.98326
R117 VTAIL.n13 VTAIL.n11 1.98326
R118 VTAIL.n14 VTAIL.n13 1.98326
R119 VTAIL.n6 VTAIL.n5 1.98326
R120 VTAIL.n5 VTAIL.n3 1.98326
R121 VTAIL.n2 VTAIL.n1 1.98326
R122 VTAIL VTAIL.n15 1.92507
R123 VTAIL.n0 VTAIL.t4 1.19184
R124 VTAIL.n0 VTAIL.t3 1.19184
R125 VTAIL.n4 VTAIL.t12 1.19184
R126 VTAIL.n4 VTAIL.t13 1.19184
R127 VTAIL.n12 VTAIL.t10 1.19184
R128 VTAIL.n12 VTAIL.t15 1.19184
R129 VTAIL.n8 VTAIL.t6 1.19184
R130 VTAIL.n8 VTAIL.t5 1.19184
R131 VTAIL.n11 VTAIL.n10 0.470328
R132 VTAIL.n3 VTAIL.n2 0.470328
R133 VTAIL VTAIL.n1 0.0586897
R134 B.n711 B.n710 585
R135 B.n713 B.n143 585
R136 B.n716 B.n715 585
R137 B.n717 B.n142 585
R138 B.n719 B.n718 585
R139 B.n721 B.n141 585
R140 B.n724 B.n723 585
R141 B.n725 B.n140 585
R142 B.n727 B.n726 585
R143 B.n729 B.n139 585
R144 B.n732 B.n731 585
R145 B.n733 B.n138 585
R146 B.n735 B.n734 585
R147 B.n737 B.n137 585
R148 B.n740 B.n739 585
R149 B.n741 B.n136 585
R150 B.n743 B.n742 585
R151 B.n745 B.n135 585
R152 B.n748 B.n747 585
R153 B.n749 B.n134 585
R154 B.n751 B.n750 585
R155 B.n753 B.n133 585
R156 B.n756 B.n755 585
R157 B.n757 B.n132 585
R158 B.n759 B.n758 585
R159 B.n761 B.n131 585
R160 B.n764 B.n763 585
R161 B.n765 B.n130 585
R162 B.n767 B.n766 585
R163 B.n769 B.n129 585
R164 B.n772 B.n771 585
R165 B.n773 B.n128 585
R166 B.n775 B.n774 585
R167 B.n777 B.n127 585
R168 B.n780 B.n779 585
R169 B.n781 B.n126 585
R170 B.n783 B.n782 585
R171 B.n785 B.n125 585
R172 B.n788 B.n787 585
R173 B.n789 B.n124 585
R174 B.n791 B.n790 585
R175 B.n793 B.n123 585
R176 B.n796 B.n795 585
R177 B.n797 B.n122 585
R178 B.n799 B.n798 585
R179 B.n801 B.n121 585
R180 B.n804 B.n803 585
R181 B.n805 B.n120 585
R182 B.n807 B.n806 585
R183 B.n809 B.n119 585
R184 B.n812 B.n811 585
R185 B.n813 B.n118 585
R186 B.n815 B.n814 585
R187 B.n817 B.n117 585
R188 B.n820 B.n819 585
R189 B.n822 B.n114 585
R190 B.n824 B.n823 585
R191 B.n826 B.n113 585
R192 B.n829 B.n828 585
R193 B.n830 B.n112 585
R194 B.n832 B.n831 585
R195 B.n834 B.n111 585
R196 B.n837 B.n836 585
R197 B.n838 B.n107 585
R198 B.n840 B.n839 585
R199 B.n842 B.n106 585
R200 B.n845 B.n844 585
R201 B.n846 B.n105 585
R202 B.n848 B.n847 585
R203 B.n850 B.n104 585
R204 B.n853 B.n852 585
R205 B.n854 B.n103 585
R206 B.n856 B.n855 585
R207 B.n858 B.n102 585
R208 B.n861 B.n860 585
R209 B.n862 B.n101 585
R210 B.n864 B.n863 585
R211 B.n866 B.n100 585
R212 B.n869 B.n868 585
R213 B.n870 B.n99 585
R214 B.n872 B.n871 585
R215 B.n874 B.n98 585
R216 B.n877 B.n876 585
R217 B.n878 B.n97 585
R218 B.n880 B.n879 585
R219 B.n882 B.n96 585
R220 B.n885 B.n884 585
R221 B.n886 B.n95 585
R222 B.n888 B.n887 585
R223 B.n890 B.n94 585
R224 B.n893 B.n892 585
R225 B.n894 B.n93 585
R226 B.n896 B.n895 585
R227 B.n898 B.n92 585
R228 B.n901 B.n900 585
R229 B.n902 B.n91 585
R230 B.n904 B.n903 585
R231 B.n906 B.n90 585
R232 B.n909 B.n908 585
R233 B.n910 B.n89 585
R234 B.n912 B.n911 585
R235 B.n914 B.n88 585
R236 B.n917 B.n916 585
R237 B.n918 B.n87 585
R238 B.n920 B.n919 585
R239 B.n922 B.n86 585
R240 B.n925 B.n924 585
R241 B.n926 B.n85 585
R242 B.n928 B.n927 585
R243 B.n930 B.n84 585
R244 B.n933 B.n932 585
R245 B.n934 B.n83 585
R246 B.n936 B.n935 585
R247 B.n938 B.n82 585
R248 B.n941 B.n940 585
R249 B.n942 B.n81 585
R250 B.n944 B.n943 585
R251 B.n946 B.n80 585
R252 B.n949 B.n948 585
R253 B.n950 B.n79 585
R254 B.n709 B.n77 585
R255 B.n953 B.n77 585
R256 B.n708 B.n76 585
R257 B.n954 B.n76 585
R258 B.n707 B.n75 585
R259 B.n955 B.n75 585
R260 B.n706 B.n705 585
R261 B.n705 B.n71 585
R262 B.n704 B.n70 585
R263 B.n961 B.n70 585
R264 B.n703 B.n69 585
R265 B.n962 B.n69 585
R266 B.n702 B.n68 585
R267 B.n963 B.n68 585
R268 B.n701 B.n700 585
R269 B.n700 B.n64 585
R270 B.n699 B.n63 585
R271 B.n969 B.n63 585
R272 B.n698 B.n62 585
R273 B.n970 B.n62 585
R274 B.n697 B.n61 585
R275 B.n971 B.n61 585
R276 B.n696 B.n695 585
R277 B.n695 B.n57 585
R278 B.n694 B.n56 585
R279 B.n977 B.n56 585
R280 B.n693 B.n55 585
R281 B.n978 B.n55 585
R282 B.n692 B.n54 585
R283 B.n979 B.n54 585
R284 B.n691 B.n690 585
R285 B.n690 B.n50 585
R286 B.n689 B.n49 585
R287 B.n985 B.n49 585
R288 B.n688 B.n48 585
R289 B.n986 B.n48 585
R290 B.n687 B.n47 585
R291 B.n987 B.n47 585
R292 B.n686 B.n685 585
R293 B.n685 B.n43 585
R294 B.n684 B.n42 585
R295 B.n993 B.n42 585
R296 B.n683 B.n41 585
R297 B.n994 B.n41 585
R298 B.n682 B.n40 585
R299 B.n995 B.n40 585
R300 B.n681 B.n680 585
R301 B.n680 B.n39 585
R302 B.n679 B.n35 585
R303 B.n1001 B.n35 585
R304 B.n678 B.n34 585
R305 B.n1002 B.n34 585
R306 B.n677 B.n33 585
R307 B.n1003 B.n33 585
R308 B.n676 B.n675 585
R309 B.n675 B.n29 585
R310 B.n674 B.n28 585
R311 B.n1009 B.n28 585
R312 B.n673 B.n27 585
R313 B.n1010 B.n27 585
R314 B.n672 B.n26 585
R315 B.n1011 B.n26 585
R316 B.n671 B.n670 585
R317 B.n670 B.n22 585
R318 B.n669 B.n21 585
R319 B.n1017 B.n21 585
R320 B.n668 B.n20 585
R321 B.n1018 B.n20 585
R322 B.n667 B.n19 585
R323 B.n1019 B.n19 585
R324 B.n666 B.n665 585
R325 B.n665 B.n15 585
R326 B.n664 B.n14 585
R327 B.n1025 B.n14 585
R328 B.n663 B.n13 585
R329 B.n1026 B.n13 585
R330 B.n662 B.n12 585
R331 B.n1027 B.n12 585
R332 B.n661 B.n660 585
R333 B.n660 B.n8 585
R334 B.n659 B.n7 585
R335 B.n1033 B.n7 585
R336 B.n658 B.n6 585
R337 B.n1034 B.n6 585
R338 B.n657 B.n5 585
R339 B.n1035 B.n5 585
R340 B.n656 B.n655 585
R341 B.n655 B.n4 585
R342 B.n654 B.n144 585
R343 B.n654 B.n653 585
R344 B.n644 B.n145 585
R345 B.n146 B.n145 585
R346 B.n646 B.n645 585
R347 B.n647 B.n646 585
R348 B.n643 B.n150 585
R349 B.n154 B.n150 585
R350 B.n642 B.n641 585
R351 B.n641 B.n640 585
R352 B.n152 B.n151 585
R353 B.n153 B.n152 585
R354 B.n633 B.n632 585
R355 B.n634 B.n633 585
R356 B.n631 B.n159 585
R357 B.n159 B.n158 585
R358 B.n630 B.n629 585
R359 B.n629 B.n628 585
R360 B.n161 B.n160 585
R361 B.n162 B.n161 585
R362 B.n621 B.n620 585
R363 B.n622 B.n621 585
R364 B.n619 B.n167 585
R365 B.n167 B.n166 585
R366 B.n618 B.n617 585
R367 B.n617 B.n616 585
R368 B.n169 B.n168 585
R369 B.n170 B.n169 585
R370 B.n609 B.n608 585
R371 B.n610 B.n609 585
R372 B.n607 B.n175 585
R373 B.n175 B.n174 585
R374 B.n606 B.n605 585
R375 B.n605 B.n604 585
R376 B.n177 B.n176 585
R377 B.n597 B.n177 585
R378 B.n596 B.n595 585
R379 B.n598 B.n596 585
R380 B.n594 B.n182 585
R381 B.n182 B.n181 585
R382 B.n593 B.n592 585
R383 B.n592 B.n591 585
R384 B.n184 B.n183 585
R385 B.n185 B.n184 585
R386 B.n584 B.n583 585
R387 B.n585 B.n584 585
R388 B.n582 B.n190 585
R389 B.n190 B.n189 585
R390 B.n581 B.n580 585
R391 B.n580 B.n579 585
R392 B.n192 B.n191 585
R393 B.n193 B.n192 585
R394 B.n572 B.n571 585
R395 B.n573 B.n572 585
R396 B.n570 B.n198 585
R397 B.n198 B.n197 585
R398 B.n569 B.n568 585
R399 B.n568 B.n567 585
R400 B.n200 B.n199 585
R401 B.n201 B.n200 585
R402 B.n560 B.n559 585
R403 B.n561 B.n560 585
R404 B.n558 B.n206 585
R405 B.n206 B.n205 585
R406 B.n557 B.n556 585
R407 B.n556 B.n555 585
R408 B.n208 B.n207 585
R409 B.n209 B.n208 585
R410 B.n548 B.n547 585
R411 B.n549 B.n548 585
R412 B.n546 B.n214 585
R413 B.n214 B.n213 585
R414 B.n545 B.n544 585
R415 B.n544 B.n543 585
R416 B.n216 B.n215 585
R417 B.n217 B.n216 585
R418 B.n536 B.n535 585
R419 B.n537 B.n536 585
R420 B.n534 B.n222 585
R421 B.n222 B.n221 585
R422 B.n533 B.n532 585
R423 B.n532 B.n531 585
R424 B.n528 B.n226 585
R425 B.n527 B.n526 585
R426 B.n524 B.n227 585
R427 B.n524 B.n225 585
R428 B.n523 B.n522 585
R429 B.n521 B.n520 585
R430 B.n519 B.n229 585
R431 B.n517 B.n516 585
R432 B.n515 B.n230 585
R433 B.n514 B.n513 585
R434 B.n511 B.n231 585
R435 B.n509 B.n508 585
R436 B.n507 B.n232 585
R437 B.n506 B.n505 585
R438 B.n503 B.n233 585
R439 B.n501 B.n500 585
R440 B.n499 B.n234 585
R441 B.n498 B.n497 585
R442 B.n495 B.n235 585
R443 B.n493 B.n492 585
R444 B.n491 B.n236 585
R445 B.n490 B.n489 585
R446 B.n487 B.n237 585
R447 B.n485 B.n484 585
R448 B.n483 B.n238 585
R449 B.n482 B.n481 585
R450 B.n479 B.n239 585
R451 B.n477 B.n476 585
R452 B.n475 B.n240 585
R453 B.n474 B.n473 585
R454 B.n471 B.n241 585
R455 B.n469 B.n468 585
R456 B.n467 B.n242 585
R457 B.n466 B.n465 585
R458 B.n463 B.n243 585
R459 B.n461 B.n460 585
R460 B.n459 B.n244 585
R461 B.n458 B.n457 585
R462 B.n455 B.n245 585
R463 B.n453 B.n452 585
R464 B.n451 B.n246 585
R465 B.n450 B.n449 585
R466 B.n447 B.n247 585
R467 B.n445 B.n444 585
R468 B.n443 B.n248 585
R469 B.n442 B.n441 585
R470 B.n439 B.n249 585
R471 B.n437 B.n436 585
R472 B.n435 B.n250 585
R473 B.n434 B.n433 585
R474 B.n431 B.n251 585
R475 B.n429 B.n428 585
R476 B.n427 B.n252 585
R477 B.n426 B.n425 585
R478 B.n423 B.n253 585
R479 B.n421 B.n420 585
R480 B.n418 B.n254 585
R481 B.n417 B.n416 585
R482 B.n414 B.n257 585
R483 B.n412 B.n411 585
R484 B.n410 B.n258 585
R485 B.n409 B.n408 585
R486 B.n406 B.n259 585
R487 B.n404 B.n403 585
R488 B.n402 B.n260 585
R489 B.n401 B.n400 585
R490 B.n398 B.n397 585
R491 B.n396 B.n395 585
R492 B.n394 B.n265 585
R493 B.n392 B.n391 585
R494 B.n390 B.n266 585
R495 B.n389 B.n388 585
R496 B.n386 B.n267 585
R497 B.n384 B.n383 585
R498 B.n382 B.n268 585
R499 B.n381 B.n380 585
R500 B.n378 B.n269 585
R501 B.n376 B.n375 585
R502 B.n374 B.n270 585
R503 B.n373 B.n372 585
R504 B.n370 B.n271 585
R505 B.n368 B.n367 585
R506 B.n366 B.n272 585
R507 B.n365 B.n364 585
R508 B.n362 B.n273 585
R509 B.n360 B.n359 585
R510 B.n358 B.n274 585
R511 B.n357 B.n356 585
R512 B.n354 B.n275 585
R513 B.n352 B.n351 585
R514 B.n350 B.n276 585
R515 B.n349 B.n348 585
R516 B.n346 B.n277 585
R517 B.n344 B.n343 585
R518 B.n342 B.n278 585
R519 B.n341 B.n340 585
R520 B.n338 B.n279 585
R521 B.n336 B.n335 585
R522 B.n334 B.n280 585
R523 B.n333 B.n332 585
R524 B.n330 B.n281 585
R525 B.n328 B.n327 585
R526 B.n326 B.n282 585
R527 B.n325 B.n324 585
R528 B.n322 B.n283 585
R529 B.n320 B.n319 585
R530 B.n318 B.n284 585
R531 B.n317 B.n316 585
R532 B.n314 B.n285 585
R533 B.n312 B.n311 585
R534 B.n310 B.n286 585
R535 B.n309 B.n308 585
R536 B.n306 B.n287 585
R537 B.n304 B.n303 585
R538 B.n302 B.n288 585
R539 B.n301 B.n300 585
R540 B.n298 B.n289 585
R541 B.n296 B.n295 585
R542 B.n294 B.n290 585
R543 B.n293 B.n292 585
R544 B.n224 B.n223 585
R545 B.n225 B.n224 585
R546 B.n530 B.n529 585
R547 B.n531 B.n530 585
R548 B.n220 B.n219 585
R549 B.n221 B.n220 585
R550 B.n539 B.n538 585
R551 B.n538 B.n537 585
R552 B.n540 B.n218 585
R553 B.n218 B.n217 585
R554 B.n542 B.n541 585
R555 B.n543 B.n542 585
R556 B.n212 B.n211 585
R557 B.n213 B.n212 585
R558 B.n551 B.n550 585
R559 B.n550 B.n549 585
R560 B.n552 B.n210 585
R561 B.n210 B.n209 585
R562 B.n554 B.n553 585
R563 B.n555 B.n554 585
R564 B.n204 B.n203 585
R565 B.n205 B.n204 585
R566 B.n563 B.n562 585
R567 B.n562 B.n561 585
R568 B.n564 B.n202 585
R569 B.n202 B.n201 585
R570 B.n566 B.n565 585
R571 B.n567 B.n566 585
R572 B.n196 B.n195 585
R573 B.n197 B.n196 585
R574 B.n575 B.n574 585
R575 B.n574 B.n573 585
R576 B.n576 B.n194 585
R577 B.n194 B.n193 585
R578 B.n578 B.n577 585
R579 B.n579 B.n578 585
R580 B.n188 B.n187 585
R581 B.n189 B.n188 585
R582 B.n587 B.n586 585
R583 B.n586 B.n585 585
R584 B.n588 B.n186 585
R585 B.n186 B.n185 585
R586 B.n590 B.n589 585
R587 B.n591 B.n590 585
R588 B.n180 B.n179 585
R589 B.n181 B.n180 585
R590 B.n600 B.n599 585
R591 B.n599 B.n598 585
R592 B.n601 B.n178 585
R593 B.n597 B.n178 585
R594 B.n603 B.n602 585
R595 B.n604 B.n603 585
R596 B.n173 B.n172 585
R597 B.n174 B.n173 585
R598 B.n612 B.n611 585
R599 B.n611 B.n610 585
R600 B.n613 B.n171 585
R601 B.n171 B.n170 585
R602 B.n615 B.n614 585
R603 B.n616 B.n615 585
R604 B.n165 B.n164 585
R605 B.n166 B.n165 585
R606 B.n624 B.n623 585
R607 B.n623 B.n622 585
R608 B.n625 B.n163 585
R609 B.n163 B.n162 585
R610 B.n627 B.n626 585
R611 B.n628 B.n627 585
R612 B.n157 B.n156 585
R613 B.n158 B.n157 585
R614 B.n636 B.n635 585
R615 B.n635 B.n634 585
R616 B.n637 B.n155 585
R617 B.n155 B.n153 585
R618 B.n639 B.n638 585
R619 B.n640 B.n639 585
R620 B.n149 B.n148 585
R621 B.n154 B.n149 585
R622 B.n649 B.n648 585
R623 B.n648 B.n647 585
R624 B.n650 B.n147 585
R625 B.n147 B.n146 585
R626 B.n652 B.n651 585
R627 B.n653 B.n652 585
R628 B.n2 B.n0 585
R629 B.n4 B.n2 585
R630 B.n3 B.n1 585
R631 B.n1034 B.n3 585
R632 B.n1032 B.n1031 585
R633 B.n1033 B.n1032 585
R634 B.n1030 B.n9 585
R635 B.n9 B.n8 585
R636 B.n1029 B.n1028 585
R637 B.n1028 B.n1027 585
R638 B.n11 B.n10 585
R639 B.n1026 B.n11 585
R640 B.n1024 B.n1023 585
R641 B.n1025 B.n1024 585
R642 B.n1022 B.n16 585
R643 B.n16 B.n15 585
R644 B.n1021 B.n1020 585
R645 B.n1020 B.n1019 585
R646 B.n18 B.n17 585
R647 B.n1018 B.n18 585
R648 B.n1016 B.n1015 585
R649 B.n1017 B.n1016 585
R650 B.n1014 B.n23 585
R651 B.n23 B.n22 585
R652 B.n1013 B.n1012 585
R653 B.n1012 B.n1011 585
R654 B.n25 B.n24 585
R655 B.n1010 B.n25 585
R656 B.n1008 B.n1007 585
R657 B.n1009 B.n1008 585
R658 B.n1006 B.n30 585
R659 B.n30 B.n29 585
R660 B.n1005 B.n1004 585
R661 B.n1004 B.n1003 585
R662 B.n32 B.n31 585
R663 B.n1002 B.n32 585
R664 B.n1000 B.n999 585
R665 B.n1001 B.n1000 585
R666 B.n998 B.n36 585
R667 B.n39 B.n36 585
R668 B.n997 B.n996 585
R669 B.n996 B.n995 585
R670 B.n38 B.n37 585
R671 B.n994 B.n38 585
R672 B.n992 B.n991 585
R673 B.n993 B.n992 585
R674 B.n990 B.n44 585
R675 B.n44 B.n43 585
R676 B.n989 B.n988 585
R677 B.n988 B.n987 585
R678 B.n46 B.n45 585
R679 B.n986 B.n46 585
R680 B.n984 B.n983 585
R681 B.n985 B.n984 585
R682 B.n982 B.n51 585
R683 B.n51 B.n50 585
R684 B.n981 B.n980 585
R685 B.n980 B.n979 585
R686 B.n53 B.n52 585
R687 B.n978 B.n53 585
R688 B.n976 B.n975 585
R689 B.n977 B.n976 585
R690 B.n974 B.n58 585
R691 B.n58 B.n57 585
R692 B.n973 B.n972 585
R693 B.n972 B.n971 585
R694 B.n60 B.n59 585
R695 B.n970 B.n60 585
R696 B.n968 B.n967 585
R697 B.n969 B.n968 585
R698 B.n966 B.n65 585
R699 B.n65 B.n64 585
R700 B.n965 B.n964 585
R701 B.n964 B.n963 585
R702 B.n67 B.n66 585
R703 B.n962 B.n67 585
R704 B.n960 B.n959 585
R705 B.n961 B.n960 585
R706 B.n958 B.n72 585
R707 B.n72 B.n71 585
R708 B.n957 B.n956 585
R709 B.n956 B.n955 585
R710 B.n74 B.n73 585
R711 B.n954 B.n74 585
R712 B.n952 B.n951 585
R713 B.n953 B.n952 585
R714 B.n1037 B.n1036 585
R715 B.n1036 B.n1035 585
R716 B.n530 B.n226 487.695
R717 B.n952 B.n79 487.695
R718 B.n532 B.n224 487.695
R719 B.n711 B.n77 487.695
R720 B.n261 B.t12 410.168
R721 B.n255 B.t8 410.168
R722 B.n108 B.t19 410.168
R723 B.n115 B.t15 410.168
R724 B.n712 B.n78 256.663
R725 B.n714 B.n78 256.663
R726 B.n720 B.n78 256.663
R727 B.n722 B.n78 256.663
R728 B.n728 B.n78 256.663
R729 B.n730 B.n78 256.663
R730 B.n736 B.n78 256.663
R731 B.n738 B.n78 256.663
R732 B.n744 B.n78 256.663
R733 B.n746 B.n78 256.663
R734 B.n752 B.n78 256.663
R735 B.n754 B.n78 256.663
R736 B.n760 B.n78 256.663
R737 B.n762 B.n78 256.663
R738 B.n768 B.n78 256.663
R739 B.n770 B.n78 256.663
R740 B.n776 B.n78 256.663
R741 B.n778 B.n78 256.663
R742 B.n784 B.n78 256.663
R743 B.n786 B.n78 256.663
R744 B.n792 B.n78 256.663
R745 B.n794 B.n78 256.663
R746 B.n800 B.n78 256.663
R747 B.n802 B.n78 256.663
R748 B.n808 B.n78 256.663
R749 B.n810 B.n78 256.663
R750 B.n816 B.n78 256.663
R751 B.n818 B.n78 256.663
R752 B.n825 B.n78 256.663
R753 B.n827 B.n78 256.663
R754 B.n833 B.n78 256.663
R755 B.n835 B.n78 256.663
R756 B.n841 B.n78 256.663
R757 B.n843 B.n78 256.663
R758 B.n849 B.n78 256.663
R759 B.n851 B.n78 256.663
R760 B.n857 B.n78 256.663
R761 B.n859 B.n78 256.663
R762 B.n865 B.n78 256.663
R763 B.n867 B.n78 256.663
R764 B.n873 B.n78 256.663
R765 B.n875 B.n78 256.663
R766 B.n881 B.n78 256.663
R767 B.n883 B.n78 256.663
R768 B.n889 B.n78 256.663
R769 B.n891 B.n78 256.663
R770 B.n897 B.n78 256.663
R771 B.n899 B.n78 256.663
R772 B.n905 B.n78 256.663
R773 B.n907 B.n78 256.663
R774 B.n913 B.n78 256.663
R775 B.n915 B.n78 256.663
R776 B.n921 B.n78 256.663
R777 B.n923 B.n78 256.663
R778 B.n929 B.n78 256.663
R779 B.n931 B.n78 256.663
R780 B.n937 B.n78 256.663
R781 B.n939 B.n78 256.663
R782 B.n945 B.n78 256.663
R783 B.n947 B.n78 256.663
R784 B.n525 B.n225 256.663
R785 B.n228 B.n225 256.663
R786 B.n518 B.n225 256.663
R787 B.n512 B.n225 256.663
R788 B.n510 B.n225 256.663
R789 B.n504 B.n225 256.663
R790 B.n502 B.n225 256.663
R791 B.n496 B.n225 256.663
R792 B.n494 B.n225 256.663
R793 B.n488 B.n225 256.663
R794 B.n486 B.n225 256.663
R795 B.n480 B.n225 256.663
R796 B.n478 B.n225 256.663
R797 B.n472 B.n225 256.663
R798 B.n470 B.n225 256.663
R799 B.n464 B.n225 256.663
R800 B.n462 B.n225 256.663
R801 B.n456 B.n225 256.663
R802 B.n454 B.n225 256.663
R803 B.n448 B.n225 256.663
R804 B.n446 B.n225 256.663
R805 B.n440 B.n225 256.663
R806 B.n438 B.n225 256.663
R807 B.n432 B.n225 256.663
R808 B.n430 B.n225 256.663
R809 B.n424 B.n225 256.663
R810 B.n422 B.n225 256.663
R811 B.n415 B.n225 256.663
R812 B.n413 B.n225 256.663
R813 B.n407 B.n225 256.663
R814 B.n405 B.n225 256.663
R815 B.n399 B.n225 256.663
R816 B.n264 B.n225 256.663
R817 B.n393 B.n225 256.663
R818 B.n387 B.n225 256.663
R819 B.n385 B.n225 256.663
R820 B.n379 B.n225 256.663
R821 B.n377 B.n225 256.663
R822 B.n371 B.n225 256.663
R823 B.n369 B.n225 256.663
R824 B.n363 B.n225 256.663
R825 B.n361 B.n225 256.663
R826 B.n355 B.n225 256.663
R827 B.n353 B.n225 256.663
R828 B.n347 B.n225 256.663
R829 B.n345 B.n225 256.663
R830 B.n339 B.n225 256.663
R831 B.n337 B.n225 256.663
R832 B.n331 B.n225 256.663
R833 B.n329 B.n225 256.663
R834 B.n323 B.n225 256.663
R835 B.n321 B.n225 256.663
R836 B.n315 B.n225 256.663
R837 B.n313 B.n225 256.663
R838 B.n307 B.n225 256.663
R839 B.n305 B.n225 256.663
R840 B.n299 B.n225 256.663
R841 B.n297 B.n225 256.663
R842 B.n291 B.n225 256.663
R843 B.n530 B.n220 163.367
R844 B.n538 B.n220 163.367
R845 B.n538 B.n218 163.367
R846 B.n542 B.n218 163.367
R847 B.n542 B.n212 163.367
R848 B.n550 B.n212 163.367
R849 B.n550 B.n210 163.367
R850 B.n554 B.n210 163.367
R851 B.n554 B.n204 163.367
R852 B.n562 B.n204 163.367
R853 B.n562 B.n202 163.367
R854 B.n566 B.n202 163.367
R855 B.n566 B.n196 163.367
R856 B.n574 B.n196 163.367
R857 B.n574 B.n194 163.367
R858 B.n578 B.n194 163.367
R859 B.n578 B.n188 163.367
R860 B.n586 B.n188 163.367
R861 B.n586 B.n186 163.367
R862 B.n590 B.n186 163.367
R863 B.n590 B.n180 163.367
R864 B.n599 B.n180 163.367
R865 B.n599 B.n178 163.367
R866 B.n603 B.n178 163.367
R867 B.n603 B.n173 163.367
R868 B.n611 B.n173 163.367
R869 B.n611 B.n171 163.367
R870 B.n615 B.n171 163.367
R871 B.n615 B.n165 163.367
R872 B.n623 B.n165 163.367
R873 B.n623 B.n163 163.367
R874 B.n627 B.n163 163.367
R875 B.n627 B.n157 163.367
R876 B.n635 B.n157 163.367
R877 B.n635 B.n155 163.367
R878 B.n639 B.n155 163.367
R879 B.n639 B.n149 163.367
R880 B.n648 B.n149 163.367
R881 B.n648 B.n147 163.367
R882 B.n652 B.n147 163.367
R883 B.n652 B.n2 163.367
R884 B.n1036 B.n2 163.367
R885 B.n1036 B.n3 163.367
R886 B.n1032 B.n3 163.367
R887 B.n1032 B.n9 163.367
R888 B.n1028 B.n9 163.367
R889 B.n1028 B.n11 163.367
R890 B.n1024 B.n11 163.367
R891 B.n1024 B.n16 163.367
R892 B.n1020 B.n16 163.367
R893 B.n1020 B.n18 163.367
R894 B.n1016 B.n18 163.367
R895 B.n1016 B.n23 163.367
R896 B.n1012 B.n23 163.367
R897 B.n1012 B.n25 163.367
R898 B.n1008 B.n25 163.367
R899 B.n1008 B.n30 163.367
R900 B.n1004 B.n30 163.367
R901 B.n1004 B.n32 163.367
R902 B.n1000 B.n32 163.367
R903 B.n1000 B.n36 163.367
R904 B.n996 B.n36 163.367
R905 B.n996 B.n38 163.367
R906 B.n992 B.n38 163.367
R907 B.n992 B.n44 163.367
R908 B.n988 B.n44 163.367
R909 B.n988 B.n46 163.367
R910 B.n984 B.n46 163.367
R911 B.n984 B.n51 163.367
R912 B.n980 B.n51 163.367
R913 B.n980 B.n53 163.367
R914 B.n976 B.n53 163.367
R915 B.n976 B.n58 163.367
R916 B.n972 B.n58 163.367
R917 B.n972 B.n60 163.367
R918 B.n968 B.n60 163.367
R919 B.n968 B.n65 163.367
R920 B.n964 B.n65 163.367
R921 B.n964 B.n67 163.367
R922 B.n960 B.n67 163.367
R923 B.n960 B.n72 163.367
R924 B.n956 B.n72 163.367
R925 B.n956 B.n74 163.367
R926 B.n952 B.n74 163.367
R927 B.n526 B.n524 163.367
R928 B.n524 B.n523 163.367
R929 B.n520 B.n519 163.367
R930 B.n517 B.n230 163.367
R931 B.n513 B.n511 163.367
R932 B.n509 B.n232 163.367
R933 B.n505 B.n503 163.367
R934 B.n501 B.n234 163.367
R935 B.n497 B.n495 163.367
R936 B.n493 B.n236 163.367
R937 B.n489 B.n487 163.367
R938 B.n485 B.n238 163.367
R939 B.n481 B.n479 163.367
R940 B.n477 B.n240 163.367
R941 B.n473 B.n471 163.367
R942 B.n469 B.n242 163.367
R943 B.n465 B.n463 163.367
R944 B.n461 B.n244 163.367
R945 B.n457 B.n455 163.367
R946 B.n453 B.n246 163.367
R947 B.n449 B.n447 163.367
R948 B.n445 B.n248 163.367
R949 B.n441 B.n439 163.367
R950 B.n437 B.n250 163.367
R951 B.n433 B.n431 163.367
R952 B.n429 B.n252 163.367
R953 B.n425 B.n423 163.367
R954 B.n421 B.n254 163.367
R955 B.n416 B.n414 163.367
R956 B.n412 B.n258 163.367
R957 B.n408 B.n406 163.367
R958 B.n404 B.n260 163.367
R959 B.n400 B.n398 163.367
R960 B.n395 B.n394 163.367
R961 B.n392 B.n266 163.367
R962 B.n388 B.n386 163.367
R963 B.n384 B.n268 163.367
R964 B.n380 B.n378 163.367
R965 B.n376 B.n270 163.367
R966 B.n372 B.n370 163.367
R967 B.n368 B.n272 163.367
R968 B.n364 B.n362 163.367
R969 B.n360 B.n274 163.367
R970 B.n356 B.n354 163.367
R971 B.n352 B.n276 163.367
R972 B.n348 B.n346 163.367
R973 B.n344 B.n278 163.367
R974 B.n340 B.n338 163.367
R975 B.n336 B.n280 163.367
R976 B.n332 B.n330 163.367
R977 B.n328 B.n282 163.367
R978 B.n324 B.n322 163.367
R979 B.n320 B.n284 163.367
R980 B.n316 B.n314 163.367
R981 B.n312 B.n286 163.367
R982 B.n308 B.n306 163.367
R983 B.n304 B.n288 163.367
R984 B.n300 B.n298 163.367
R985 B.n296 B.n290 163.367
R986 B.n292 B.n224 163.367
R987 B.n532 B.n222 163.367
R988 B.n536 B.n222 163.367
R989 B.n536 B.n216 163.367
R990 B.n544 B.n216 163.367
R991 B.n544 B.n214 163.367
R992 B.n548 B.n214 163.367
R993 B.n548 B.n208 163.367
R994 B.n556 B.n208 163.367
R995 B.n556 B.n206 163.367
R996 B.n560 B.n206 163.367
R997 B.n560 B.n200 163.367
R998 B.n568 B.n200 163.367
R999 B.n568 B.n198 163.367
R1000 B.n572 B.n198 163.367
R1001 B.n572 B.n192 163.367
R1002 B.n580 B.n192 163.367
R1003 B.n580 B.n190 163.367
R1004 B.n584 B.n190 163.367
R1005 B.n584 B.n184 163.367
R1006 B.n592 B.n184 163.367
R1007 B.n592 B.n182 163.367
R1008 B.n596 B.n182 163.367
R1009 B.n596 B.n177 163.367
R1010 B.n605 B.n177 163.367
R1011 B.n605 B.n175 163.367
R1012 B.n609 B.n175 163.367
R1013 B.n609 B.n169 163.367
R1014 B.n617 B.n169 163.367
R1015 B.n617 B.n167 163.367
R1016 B.n621 B.n167 163.367
R1017 B.n621 B.n161 163.367
R1018 B.n629 B.n161 163.367
R1019 B.n629 B.n159 163.367
R1020 B.n633 B.n159 163.367
R1021 B.n633 B.n152 163.367
R1022 B.n641 B.n152 163.367
R1023 B.n641 B.n150 163.367
R1024 B.n646 B.n150 163.367
R1025 B.n646 B.n145 163.367
R1026 B.n654 B.n145 163.367
R1027 B.n655 B.n654 163.367
R1028 B.n655 B.n5 163.367
R1029 B.n6 B.n5 163.367
R1030 B.n7 B.n6 163.367
R1031 B.n660 B.n7 163.367
R1032 B.n660 B.n12 163.367
R1033 B.n13 B.n12 163.367
R1034 B.n14 B.n13 163.367
R1035 B.n665 B.n14 163.367
R1036 B.n665 B.n19 163.367
R1037 B.n20 B.n19 163.367
R1038 B.n21 B.n20 163.367
R1039 B.n670 B.n21 163.367
R1040 B.n670 B.n26 163.367
R1041 B.n27 B.n26 163.367
R1042 B.n28 B.n27 163.367
R1043 B.n675 B.n28 163.367
R1044 B.n675 B.n33 163.367
R1045 B.n34 B.n33 163.367
R1046 B.n35 B.n34 163.367
R1047 B.n680 B.n35 163.367
R1048 B.n680 B.n40 163.367
R1049 B.n41 B.n40 163.367
R1050 B.n42 B.n41 163.367
R1051 B.n685 B.n42 163.367
R1052 B.n685 B.n47 163.367
R1053 B.n48 B.n47 163.367
R1054 B.n49 B.n48 163.367
R1055 B.n690 B.n49 163.367
R1056 B.n690 B.n54 163.367
R1057 B.n55 B.n54 163.367
R1058 B.n56 B.n55 163.367
R1059 B.n695 B.n56 163.367
R1060 B.n695 B.n61 163.367
R1061 B.n62 B.n61 163.367
R1062 B.n63 B.n62 163.367
R1063 B.n700 B.n63 163.367
R1064 B.n700 B.n68 163.367
R1065 B.n69 B.n68 163.367
R1066 B.n70 B.n69 163.367
R1067 B.n705 B.n70 163.367
R1068 B.n705 B.n75 163.367
R1069 B.n76 B.n75 163.367
R1070 B.n77 B.n76 163.367
R1071 B.n948 B.n946 163.367
R1072 B.n944 B.n81 163.367
R1073 B.n940 B.n938 163.367
R1074 B.n936 B.n83 163.367
R1075 B.n932 B.n930 163.367
R1076 B.n928 B.n85 163.367
R1077 B.n924 B.n922 163.367
R1078 B.n920 B.n87 163.367
R1079 B.n916 B.n914 163.367
R1080 B.n912 B.n89 163.367
R1081 B.n908 B.n906 163.367
R1082 B.n904 B.n91 163.367
R1083 B.n900 B.n898 163.367
R1084 B.n896 B.n93 163.367
R1085 B.n892 B.n890 163.367
R1086 B.n888 B.n95 163.367
R1087 B.n884 B.n882 163.367
R1088 B.n880 B.n97 163.367
R1089 B.n876 B.n874 163.367
R1090 B.n872 B.n99 163.367
R1091 B.n868 B.n866 163.367
R1092 B.n864 B.n101 163.367
R1093 B.n860 B.n858 163.367
R1094 B.n856 B.n103 163.367
R1095 B.n852 B.n850 163.367
R1096 B.n848 B.n105 163.367
R1097 B.n844 B.n842 163.367
R1098 B.n840 B.n107 163.367
R1099 B.n836 B.n834 163.367
R1100 B.n832 B.n112 163.367
R1101 B.n828 B.n826 163.367
R1102 B.n824 B.n114 163.367
R1103 B.n819 B.n817 163.367
R1104 B.n815 B.n118 163.367
R1105 B.n811 B.n809 163.367
R1106 B.n807 B.n120 163.367
R1107 B.n803 B.n801 163.367
R1108 B.n799 B.n122 163.367
R1109 B.n795 B.n793 163.367
R1110 B.n791 B.n124 163.367
R1111 B.n787 B.n785 163.367
R1112 B.n783 B.n126 163.367
R1113 B.n779 B.n777 163.367
R1114 B.n775 B.n128 163.367
R1115 B.n771 B.n769 163.367
R1116 B.n767 B.n130 163.367
R1117 B.n763 B.n761 163.367
R1118 B.n759 B.n132 163.367
R1119 B.n755 B.n753 163.367
R1120 B.n751 B.n134 163.367
R1121 B.n747 B.n745 163.367
R1122 B.n743 B.n136 163.367
R1123 B.n739 B.n737 163.367
R1124 B.n735 B.n138 163.367
R1125 B.n731 B.n729 163.367
R1126 B.n727 B.n140 163.367
R1127 B.n723 B.n721 163.367
R1128 B.n719 B.n142 163.367
R1129 B.n715 B.n713 163.367
R1130 B.n261 B.t14 117.761
R1131 B.n115 B.t17 117.761
R1132 B.n255 B.t11 117.74
R1133 B.n108 B.t20 117.74
R1134 B.n262 B.t13 73.1559
R1135 B.n116 B.t18 73.1559
R1136 B.n256 B.t10 73.1342
R1137 B.n109 B.t21 73.1342
R1138 B.n525 B.n226 71.676
R1139 B.n523 B.n228 71.676
R1140 B.n519 B.n518 71.676
R1141 B.n512 B.n230 71.676
R1142 B.n511 B.n510 71.676
R1143 B.n504 B.n232 71.676
R1144 B.n503 B.n502 71.676
R1145 B.n496 B.n234 71.676
R1146 B.n495 B.n494 71.676
R1147 B.n488 B.n236 71.676
R1148 B.n487 B.n486 71.676
R1149 B.n480 B.n238 71.676
R1150 B.n479 B.n478 71.676
R1151 B.n472 B.n240 71.676
R1152 B.n471 B.n470 71.676
R1153 B.n464 B.n242 71.676
R1154 B.n463 B.n462 71.676
R1155 B.n456 B.n244 71.676
R1156 B.n455 B.n454 71.676
R1157 B.n448 B.n246 71.676
R1158 B.n447 B.n446 71.676
R1159 B.n440 B.n248 71.676
R1160 B.n439 B.n438 71.676
R1161 B.n432 B.n250 71.676
R1162 B.n431 B.n430 71.676
R1163 B.n424 B.n252 71.676
R1164 B.n423 B.n422 71.676
R1165 B.n415 B.n254 71.676
R1166 B.n414 B.n413 71.676
R1167 B.n407 B.n258 71.676
R1168 B.n406 B.n405 71.676
R1169 B.n399 B.n260 71.676
R1170 B.n398 B.n264 71.676
R1171 B.n394 B.n393 71.676
R1172 B.n387 B.n266 71.676
R1173 B.n386 B.n385 71.676
R1174 B.n379 B.n268 71.676
R1175 B.n378 B.n377 71.676
R1176 B.n371 B.n270 71.676
R1177 B.n370 B.n369 71.676
R1178 B.n363 B.n272 71.676
R1179 B.n362 B.n361 71.676
R1180 B.n355 B.n274 71.676
R1181 B.n354 B.n353 71.676
R1182 B.n347 B.n276 71.676
R1183 B.n346 B.n345 71.676
R1184 B.n339 B.n278 71.676
R1185 B.n338 B.n337 71.676
R1186 B.n331 B.n280 71.676
R1187 B.n330 B.n329 71.676
R1188 B.n323 B.n282 71.676
R1189 B.n322 B.n321 71.676
R1190 B.n315 B.n284 71.676
R1191 B.n314 B.n313 71.676
R1192 B.n307 B.n286 71.676
R1193 B.n306 B.n305 71.676
R1194 B.n299 B.n288 71.676
R1195 B.n298 B.n297 71.676
R1196 B.n291 B.n290 71.676
R1197 B.n947 B.n79 71.676
R1198 B.n946 B.n945 71.676
R1199 B.n939 B.n81 71.676
R1200 B.n938 B.n937 71.676
R1201 B.n931 B.n83 71.676
R1202 B.n930 B.n929 71.676
R1203 B.n923 B.n85 71.676
R1204 B.n922 B.n921 71.676
R1205 B.n915 B.n87 71.676
R1206 B.n914 B.n913 71.676
R1207 B.n907 B.n89 71.676
R1208 B.n906 B.n905 71.676
R1209 B.n899 B.n91 71.676
R1210 B.n898 B.n897 71.676
R1211 B.n891 B.n93 71.676
R1212 B.n890 B.n889 71.676
R1213 B.n883 B.n95 71.676
R1214 B.n882 B.n881 71.676
R1215 B.n875 B.n97 71.676
R1216 B.n874 B.n873 71.676
R1217 B.n867 B.n99 71.676
R1218 B.n866 B.n865 71.676
R1219 B.n859 B.n101 71.676
R1220 B.n858 B.n857 71.676
R1221 B.n851 B.n103 71.676
R1222 B.n850 B.n849 71.676
R1223 B.n843 B.n105 71.676
R1224 B.n842 B.n841 71.676
R1225 B.n835 B.n107 71.676
R1226 B.n834 B.n833 71.676
R1227 B.n827 B.n112 71.676
R1228 B.n826 B.n825 71.676
R1229 B.n818 B.n114 71.676
R1230 B.n817 B.n816 71.676
R1231 B.n810 B.n118 71.676
R1232 B.n809 B.n808 71.676
R1233 B.n802 B.n120 71.676
R1234 B.n801 B.n800 71.676
R1235 B.n794 B.n122 71.676
R1236 B.n793 B.n792 71.676
R1237 B.n786 B.n124 71.676
R1238 B.n785 B.n784 71.676
R1239 B.n778 B.n126 71.676
R1240 B.n777 B.n776 71.676
R1241 B.n770 B.n128 71.676
R1242 B.n769 B.n768 71.676
R1243 B.n762 B.n130 71.676
R1244 B.n761 B.n760 71.676
R1245 B.n754 B.n132 71.676
R1246 B.n753 B.n752 71.676
R1247 B.n746 B.n134 71.676
R1248 B.n745 B.n744 71.676
R1249 B.n738 B.n136 71.676
R1250 B.n737 B.n736 71.676
R1251 B.n730 B.n138 71.676
R1252 B.n729 B.n728 71.676
R1253 B.n722 B.n140 71.676
R1254 B.n721 B.n720 71.676
R1255 B.n714 B.n142 71.676
R1256 B.n713 B.n712 71.676
R1257 B.n712 B.n711 71.676
R1258 B.n715 B.n714 71.676
R1259 B.n720 B.n719 71.676
R1260 B.n723 B.n722 71.676
R1261 B.n728 B.n727 71.676
R1262 B.n731 B.n730 71.676
R1263 B.n736 B.n735 71.676
R1264 B.n739 B.n738 71.676
R1265 B.n744 B.n743 71.676
R1266 B.n747 B.n746 71.676
R1267 B.n752 B.n751 71.676
R1268 B.n755 B.n754 71.676
R1269 B.n760 B.n759 71.676
R1270 B.n763 B.n762 71.676
R1271 B.n768 B.n767 71.676
R1272 B.n771 B.n770 71.676
R1273 B.n776 B.n775 71.676
R1274 B.n779 B.n778 71.676
R1275 B.n784 B.n783 71.676
R1276 B.n787 B.n786 71.676
R1277 B.n792 B.n791 71.676
R1278 B.n795 B.n794 71.676
R1279 B.n800 B.n799 71.676
R1280 B.n803 B.n802 71.676
R1281 B.n808 B.n807 71.676
R1282 B.n811 B.n810 71.676
R1283 B.n816 B.n815 71.676
R1284 B.n819 B.n818 71.676
R1285 B.n825 B.n824 71.676
R1286 B.n828 B.n827 71.676
R1287 B.n833 B.n832 71.676
R1288 B.n836 B.n835 71.676
R1289 B.n841 B.n840 71.676
R1290 B.n844 B.n843 71.676
R1291 B.n849 B.n848 71.676
R1292 B.n852 B.n851 71.676
R1293 B.n857 B.n856 71.676
R1294 B.n860 B.n859 71.676
R1295 B.n865 B.n864 71.676
R1296 B.n868 B.n867 71.676
R1297 B.n873 B.n872 71.676
R1298 B.n876 B.n875 71.676
R1299 B.n881 B.n880 71.676
R1300 B.n884 B.n883 71.676
R1301 B.n889 B.n888 71.676
R1302 B.n892 B.n891 71.676
R1303 B.n897 B.n896 71.676
R1304 B.n900 B.n899 71.676
R1305 B.n905 B.n904 71.676
R1306 B.n908 B.n907 71.676
R1307 B.n913 B.n912 71.676
R1308 B.n916 B.n915 71.676
R1309 B.n921 B.n920 71.676
R1310 B.n924 B.n923 71.676
R1311 B.n929 B.n928 71.676
R1312 B.n932 B.n931 71.676
R1313 B.n937 B.n936 71.676
R1314 B.n940 B.n939 71.676
R1315 B.n945 B.n944 71.676
R1316 B.n948 B.n947 71.676
R1317 B.n526 B.n525 71.676
R1318 B.n520 B.n228 71.676
R1319 B.n518 B.n517 71.676
R1320 B.n513 B.n512 71.676
R1321 B.n510 B.n509 71.676
R1322 B.n505 B.n504 71.676
R1323 B.n502 B.n501 71.676
R1324 B.n497 B.n496 71.676
R1325 B.n494 B.n493 71.676
R1326 B.n489 B.n488 71.676
R1327 B.n486 B.n485 71.676
R1328 B.n481 B.n480 71.676
R1329 B.n478 B.n477 71.676
R1330 B.n473 B.n472 71.676
R1331 B.n470 B.n469 71.676
R1332 B.n465 B.n464 71.676
R1333 B.n462 B.n461 71.676
R1334 B.n457 B.n456 71.676
R1335 B.n454 B.n453 71.676
R1336 B.n449 B.n448 71.676
R1337 B.n446 B.n445 71.676
R1338 B.n441 B.n440 71.676
R1339 B.n438 B.n437 71.676
R1340 B.n433 B.n432 71.676
R1341 B.n430 B.n429 71.676
R1342 B.n425 B.n424 71.676
R1343 B.n422 B.n421 71.676
R1344 B.n416 B.n415 71.676
R1345 B.n413 B.n412 71.676
R1346 B.n408 B.n407 71.676
R1347 B.n405 B.n404 71.676
R1348 B.n400 B.n399 71.676
R1349 B.n395 B.n264 71.676
R1350 B.n393 B.n392 71.676
R1351 B.n388 B.n387 71.676
R1352 B.n385 B.n384 71.676
R1353 B.n380 B.n379 71.676
R1354 B.n377 B.n376 71.676
R1355 B.n372 B.n371 71.676
R1356 B.n369 B.n368 71.676
R1357 B.n364 B.n363 71.676
R1358 B.n361 B.n360 71.676
R1359 B.n356 B.n355 71.676
R1360 B.n353 B.n352 71.676
R1361 B.n348 B.n347 71.676
R1362 B.n345 B.n344 71.676
R1363 B.n340 B.n339 71.676
R1364 B.n337 B.n336 71.676
R1365 B.n332 B.n331 71.676
R1366 B.n329 B.n328 71.676
R1367 B.n324 B.n323 71.676
R1368 B.n321 B.n320 71.676
R1369 B.n316 B.n315 71.676
R1370 B.n313 B.n312 71.676
R1371 B.n308 B.n307 71.676
R1372 B.n305 B.n304 71.676
R1373 B.n300 B.n299 71.676
R1374 B.n297 B.n296 71.676
R1375 B.n292 B.n291 71.676
R1376 B.n531 B.n225 59.7858
R1377 B.n953 B.n78 59.7858
R1378 B.n263 B.n262 59.5399
R1379 B.n419 B.n256 59.5399
R1380 B.n110 B.n109 59.5399
R1381 B.n821 B.n116 59.5399
R1382 B.n262 B.n261 44.6066
R1383 B.n256 B.n255 44.6066
R1384 B.n109 B.n108 44.6066
R1385 B.n116 B.n115 44.6066
R1386 B.n531 B.n221 34.1636
R1387 B.n537 B.n221 34.1636
R1388 B.n537 B.n217 34.1636
R1389 B.n543 B.n217 34.1636
R1390 B.n543 B.n213 34.1636
R1391 B.n549 B.n213 34.1636
R1392 B.n555 B.n209 34.1636
R1393 B.n555 B.n205 34.1636
R1394 B.n561 B.n205 34.1636
R1395 B.n561 B.n201 34.1636
R1396 B.n567 B.n201 34.1636
R1397 B.n567 B.n197 34.1636
R1398 B.n573 B.n197 34.1636
R1399 B.n573 B.n193 34.1636
R1400 B.n579 B.n193 34.1636
R1401 B.n585 B.n189 34.1636
R1402 B.n585 B.n185 34.1636
R1403 B.n591 B.n185 34.1636
R1404 B.n591 B.n181 34.1636
R1405 B.n598 B.n181 34.1636
R1406 B.n598 B.n597 34.1636
R1407 B.n604 B.n174 34.1636
R1408 B.n610 B.n174 34.1636
R1409 B.n610 B.n170 34.1636
R1410 B.n616 B.n170 34.1636
R1411 B.n616 B.n166 34.1636
R1412 B.n622 B.n166 34.1636
R1413 B.n628 B.n162 34.1636
R1414 B.n628 B.n158 34.1636
R1415 B.n634 B.n158 34.1636
R1416 B.n634 B.n153 34.1636
R1417 B.n640 B.n153 34.1636
R1418 B.n640 B.n154 34.1636
R1419 B.n647 B.n146 34.1636
R1420 B.n653 B.n146 34.1636
R1421 B.n653 B.n4 34.1636
R1422 B.n1035 B.n4 34.1636
R1423 B.n1035 B.n1034 34.1636
R1424 B.n1034 B.n1033 34.1636
R1425 B.n1033 B.n8 34.1636
R1426 B.n1027 B.n8 34.1636
R1427 B.n1026 B.n1025 34.1636
R1428 B.n1025 B.n15 34.1636
R1429 B.n1019 B.n15 34.1636
R1430 B.n1019 B.n1018 34.1636
R1431 B.n1018 B.n1017 34.1636
R1432 B.n1017 B.n22 34.1636
R1433 B.n1011 B.n1010 34.1636
R1434 B.n1010 B.n1009 34.1636
R1435 B.n1009 B.n29 34.1636
R1436 B.n1003 B.n29 34.1636
R1437 B.n1003 B.n1002 34.1636
R1438 B.n1002 B.n1001 34.1636
R1439 B.n995 B.n39 34.1636
R1440 B.n995 B.n994 34.1636
R1441 B.n994 B.n993 34.1636
R1442 B.n993 B.n43 34.1636
R1443 B.n987 B.n43 34.1636
R1444 B.n987 B.n986 34.1636
R1445 B.n985 B.n50 34.1636
R1446 B.n979 B.n50 34.1636
R1447 B.n979 B.n978 34.1636
R1448 B.n978 B.n977 34.1636
R1449 B.n977 B.n57 34.1636
R1450 B.n971 B.n57 34.1636
R1451 B.n971 B.n970 34.1636
R1452 B.n970 B.n969 34.1636
R1453 B.n969 B.n64 34.1636
R1454 B.n963 B.n962 34.1636
R1455 B.n962 B.n961 34.1636
R1456 B.n961 B.n71 34.1636
R1457 B.n955 B.n71 34.1636
R1458 B.n955 B.n954 34.1636
R1459 B.n954 B.n953 34.1636
R1460 B.n647 B.t0 33.6612
R1461 B.n1027 B.t1 33.6612
R1462 B.n951 B.n950 31.6883
R1463 B.n710 B.n709 31.6883
R1464 B.n533 B.n223 31.6883
R1465 B.n529 B.n528 31.6883
R1466 B.n549 B.t9 25.6228
R1467 B.t5 B.n162 25.6228
R1468 B.t4 B.n22 25.6228
R1469 B.n963 B.t16 25.6228
R1470 B.n579 B.t2 24.618
R1471 B.t7 B.n985 24.618
R1472 B B.n1037 18.0485
R1473 B.n604 B.t6 17.5844
R1474 B.n1001 B.t3 17.5844
R1475 B.n597 B.t6 16.5796
R1476 B.n39 B.t3 16.5796
R1477 B.n950 B.n949 10.6151
R1478 B.n949 B.n80 10.6151
R1479 B.n943 B.n80 10.6151
R1480 B.n943 B.n942 10.6151
R1481 B.n942 B.n941 10.6151
R1482 B.n941 B.n82 10.6151
R1483 B.n935 B.n82 10.6151
R1484 B.n935 B.n934 10.6151
R1485 B.n934 B.n933 10.6151
R1486 B.n933 B.n84 10.6151
R1487 B.n927 B.n84 10.6151
R1488 B.n927 B.n926 10.6151
R1489 B.n926 B.n925 10.6151
R1490 B.n925 B.n86 10.6151
R1491 B.n919 B.n86 10.6151
R1492 B.n919 B.n918 10.6151
R1493 B.n918 B.n917 10.6151
R1494 B.n917 B.n88 10.6151
R1495 B.n911 B.n88 10.6151
R1496 B.n911 B.n910 10.6151
R1497 B.n910 B.n909 10.6151
R1498 B.n909 B.n90 10.6151
R1499 B.n903 B.n90 10.6151
R1500 B.n903 B.n902 10.6151
R1501 B.n902 B.n901 10.6151
R1502 B.n901 B.n92 10.6151
R1503 B.n895 B.n92 10.6151
R1504 B.n895 B.n894 10.6151
R1505 B.n894 B.n893 10.6151
R1506 B.n893 B.n94 10.6151
R1507 B.n887 B.n94 10.6151
R1508 B.n887 B.n886 10.6151
R1509 B.n886 B.n885 10.6151
R1510 B.n885 B.n96 10.6151
R1511 B.n879 B.n96 10.6151
R1512 B.n879 B.n878 10.6151
R1513 B.n878 B.n877 10.6151
R1514 B.n877 B.n98 10.6151
R1515 B.n871 B.n98 10.6151
R1516 B.n871 B.n870 10.6151
R1517 B.n870 B.n869 10.6151
R1518 B.n869 B.n100 10.6151
R1519 B.n863 B.n100 10.6151
R1520 B.n863 B.n862 10.6151
R1521 B.n862 B.n861 10.6151
R1522 B.n861 B.n102 10.6151
R1523 B.n855 B.n102 10.6151
R1524 B.n855 B.n854 10.6151
R1525 B.n854 B.n853 10.6151
R1526 B.n853 B.n104 10.6151
R1527 B.n847 B.n104 10.6151
R1528 B.n847 B.n846 10.6151
R1529 B.n846 B.n845 10.6151
R1530 B.n845 B.n106 10.6151
R1531 B.n839 B.n838 10.6151
R1532 B.n838 B.n837 10.6151
R1533 B.n837 B.n111 10.6151
R1534 B.n831 B.n111 10.6151
R1535 B.n831 B.n830 10.6151
R1536 B.n830 B.n829 10.6151
R1537 B.n829 B.n113 10.6151
R1538 B.n823 B.n113 10.6151
R1539 B.n823 B.n822 10.6151
R1540 B.n820 B.n117 10.6151
R1541 B.n814 B.n117 10.6151
R1542 B.n814 B.n813 10.6151
R1543 B.n813 B.n812 10.6151
R1544 B.n812 B.n119 10.6151
R1545 B.n806 B.n119 10.6151
R1546 B.n806 B.n805 10.6151
R1547 B.n805 B.n804 10.6151
R1548 B.n804 B.n121 10.6151
R1549 B.n798 B.n121 10.6151
R1550 B.n798 B.n797 10.6151
R1551 B.n797 B.n796 10.6151
R1552 B.n796 B.n123 10.6151
R1553 B.n790 B.n123 10.6151
R1554 B.n790 B.n789 10.6151
R1555 B.n789 B.n788 10.6151
R1556 B.n788 B.n125 10.6151
R1557 B.n782 B.n125 10.6151
R1558 B.n782 B.n781 10.6151
R1559 B.n781 B.n780 10.6151
R1560 B.n780 B.n127 10.6151
R1561 B.n774 B.n127 10.6151
R1562 B.n774 B.n773 10.6151
R1563 B.n773 B.n772 10.6151
R1564 B.n772 B.n129 10.6151
R1565 B.n766 B.n129 10.6151
R1566 B.n766 B.n765 10.6151
R1567 B.n765 B.n764 10.6151
R1568 B.n764 B.n131 10.6151
R1569 B.n758 B.n131 10.6151
R1570 B.n758 B.n757 10.6151
R1571 B.n757 B.n756 10.6151
R1572 B.n756 B.n133 10.6151
R1573 B.n750 B.n133 10.6151
R1574 B.n750 B.n749 10.6151
R1575 B.n749 B.n748 10.6151
R1576 B.n748 B.n135 10.6151
R1577 B.n742 B.n135 10.6151
R1578 B.n742 B.n741 10.6151
R1579 B.n741 B.n740 10.6151
R1580 B.n740 B.n137 10.6151
R1581 B.n734 B.n137 10.6151
R1582 B.n734 B.n733 10.6151
R1583 B.n733 B.n732 10.6151
R1584 B.n732 B.n139 10.6151
R1585 B.n726 B.n139 10.6151
R1586 B.n726 B.n725 10.6151
R1587 B.n725 B.n724 10.6151
R1588 B.n724 B.n141 10.6151
R1589 B.n718 B.n141 10.6151
R1590 B.n718 B.n717 10.6151
R1591 B.n717 B.n716 10.6151
R1592 B.n716 B.n143 10.6151
R1593 B.n710 B.n143 10.6151
R1594 B.n534 B.n533 10.6151
R1595 B.n535 B.n534 10.6151
R1596 B.n535 B.n215 10.6151
R1597 B.n545 B.n215 10.6151
R1598 B.n546 B.n545 10.6151
R1599 B.n547 B.n546 10.6151
R1600 B.n547 B.n207 10.6151
R1601 B.n557 B.n207 10.6151
R1602 B.n558 B.n557 10.6151
R1603 B.n559 B.n558 10.6151
R1604 B.n559 B.n199 10.6151
R1605 B.n569 B.n199 10.6151
R1606 B.n570 B.n569 10.6151
R1607 B.n571 B.n570 10.6151
R1608 B.n571 B.n191 10.6151
R1609 B.n581 B.n191 10.6151
R1610 B.n582 B.n581 10.6151
R1611 B.n583 B.n582 10.6151
R1612 B.n583 B.n183 10.6151
R1613 B.n593 B.n183 10.6151
R1614 B.n594 B.n593 10.6151
R1615 B.n595 B.n594 10.6151
R1616 B.n595 B.n176 10.6151
R1617 B.n606 B.n176 10.6151
R1618 B.n607 B.n606 10.6151
R1619 B.n608 B.n607 10.6151
R1620 B.n608 B.n168 10.6151
R1621 B.n618 B.n168 10.6151
R1622 B.n619 B.n618 10.6151
R1623 B.n620 B.n619 10.6151
R1624 B.n620 B.n160 10.6151
R1625 B.n630 B.n160 10.6151
R1626 B.n631 B.n630 10.6151
R1627 B.n632 B.n631 10.6151
R1628 B.n632 B.n151 10.6151
R1629 B.n642 B.n151 10.6151
R1630 B.n643 B.n642 10.6151
R1631 B.n645 B.n643 10.6151
R1632 B.n645 B.n644 10.6151
R1633 B.n644 B.n144 10.6151
R1634 B.n656 B.n144 10.6151
R1635 B.n657 B.n656 10.6151
R1636 B.n658 B.n657 10.6151
R1637 B.n659 B.n658 10.6151
R1638 B.n661 B.n659 10.6151
R1639 B.n662 B.n661 10.6151
R1640 B.n663 B.n662 10.6151
R1641 B.n664 B.n663 10.6151
R1642 B.n666 B.n664 10.6151
R1643 B.n667 B.n666 10.6151
R1644 B.n668 B.n667 10.6151
R1645 B.n669 B.n668 10.6151
R1646 B.n671 B.n669 10.6151
R1647 B.n672 B.n671 10.6151
R1648 B.n673 B.n672 10.6151
R1649 B.n674 B.n673 10.6151
R1650 B.n676 B.n674 10.6151
R1651 B.n677 B.n676 10.6151
R1652 B.n678 B.n677 10.6151
R1653 B.n679 B.n678 10.6151
R1654 B.n681 B.n679 10.6151
R1655 B.n682 B.n681 10.6151
R1656 B.n683 B.n682 10.6151
R1657 B.n684 B.n683 10.6151
R1658 B.n686 B.n684 10.6151
R1659 B.n687 B.n686 10.6151
R1660 B.n688 B.n687 10.6151
R1661 B.n689 B.n688 10.6151
R1662 B.n691 B.n689 10.6151
R1663 B.n692 B.n691 10.6151
R1664 B.n693 B.n692 10.6151
R1665 B.n694 B.n693 10.6151
R1666 B.n696 B.n694 10.6151
R1667 B.n697 B.n696 10.6151
R1668 B.n698 B.n697 10.6151
R1669 B.n699 B.n698 10.6151
R1670 B.n701 B.n699 10.6151
R1671 B.n702 B.n701 10.6151
R1672 B.n703 B.n702 10.6151
R1673 B.n704 B.n703 10.6151
R1674 B.n706 B.n704 10.6151
R1675 B.n707 B.n706 10.6151
R1676 B.n708 B.n707 10.6151
R1677 B.n709 B.n708 10.6151
R1678 B.n528 B.n527 10.6151
R1679 B.n527 B.n227 10.6151
R1680 B.n522 B.n227 10.6151
R1681 B.n522 B.n521 10.6151
R1682 B.n521 B.n229 10.6151
R1683 B.n516 B.n229 10.6151
R1684 B.n516 B.n515 10.6151
R1685 B.n515 B.n514 10.6151
R1686 B.n514 B.n231 10.6151
R1687 B.n508 B.n231 10.6151
R1688 B.n508 B.n507 10.6151
R1689 B.n507 B.n506 10.6151
R1690 B.n506 B.n233 10.6151
R1691 B.n500 B.n233 10.6151
R1692 B.n500 B.n499 10.6151
R1693 B.n499 B.n498 10.6151
R1694 B.n498 B.n235 10.6151
R1695 B.n492 B.n235 10.6151
R1696 B.n492 B.n491 10.6151
R1697 B.n491 B.n490 10.6151
R1698 B.n490 B.n237 10.6151
R1699 B.n484 B.n237 10.6151
R1700 B.n484 B.n483 10.6151
R1701 B.n483 B.n482 10.6151
R1702 B.n482 B.n239 10.6151
R1703 B.n476 B.n239 10.6151
R1704 B.n476 B.n475 10.6151
R1705 B.n475 B.n474 10.6151
R1706 B.n474 B.n241 10.6151
R1707 B.n468 B.n241 10.6151
R1708 B.n468 B.n467 10.6151
R1709 B.n467 B.n466 10.6151
R1710 B.n466 B.n243 10.6151
R1711 B.n460 B.n243 10.6151
R1712 B.n460 B.n459 10.6151
R1713 B.n459 B.n458 10.6151
R1714 B.n458 B.n245 10.6151
R1715 B.n452 B.n245 10.6151
R1716 B.n452 B.n451 10.6151
R1717 B.n451 B.n450 10.6151
R1718 B.n450 B.n247 10.6151
R1719 B.n444 B.n247 10.6151
R1720 B.n444 B.n443 10.6151
R1721 B.n443 B.n442 10.6151
R1722 B.n442 B.n249 10.6151
R1723 B.n436 B.n249 10.6151
R1724 B.n436 B.n435 10.6151
R1725 B.n435 B.n434 10.6151
R1726 B.n434 B.n251 10.6151
R1727 B.n428 B.n251 10.6151
R1728 B.n428 B.n427 10.6151
R1729 B.n427 B.n426 10.6151
R1730 B.n426 B.n253 10.6151
R1731 B.n420 B.n253 10.6151
R1732 B.n418 B.n417 10.6151
R1733 B.n417 B.n257 10.6151
R1734 B.n411 B.n257 10.6151
R1735 B.n411 B.n410 10.6151
R1736 B.n410 B.n409 10.6151
R1737 B.n409 B.n259 10.6151
R1738 B.n403 B.n259 10.6151
R1739 B.n403 B.n402 10.6151
R1740 B.n402 B.n401 10.6151
R1741 B.n397 B.n396 10.6151
R1742 B.n396 B.n265 10.6151
R1743 B.n391 B.n265 10.6151
R1744 B.n391 B.n390 10.6151
R1745 B.n390 B.n389 10.6151
R1746 B.n389 B.n267 10.6151
R1747 B.n383 B.n267 10.6151
R1748 B.n383 B.n382 10.6151
R1749 B.n382 B.n381 10.6151
R1750 B.n381 B.n269 10.6151
R1751 B.n375 B.n269 10.6151
R1752 B.n375 B.n374 10.6151
R1753 B.n374 B.n373 10.6151
R1754 B.n373 B.n271 10.6151
R1755 B.n367 B.n271 10.6151
R1756 B.n367 B.n366 10.6151
R1757 B.n366 B.n365 10.6151
R1758 B.n365 B.n273 10.6151
R1759 B.n359 B.n273 10.6151
R1760 B.n359 B.n358 10.6151
R1761 B.n358 B.n357 10.6151
R1762 B.n357 B.n275 10.6151
R1763 B.n351 B.n275 10.6151
R1764 B.n351 B.n350 10.6151
R1765 B.n350 B.n349 10.6151
R1766 B.n349 B.n277 10.6151
R1767 B.n343 B.n277 10.6151
R1768 B.n343 B.n342 10.6151
R1769 B.n342 B.n341 10.6151
R1770 B.n341 B.n279 10.6151
R1771 B.n335 B.n279 10.6151
R1772 B.n335 B.n334 10.6151
R1773 B.n334 B.n333 10.6151
R1774 B.n333 B.n281 10.6151
R1775 B.n327 B.n281 10.6151
R1776 B.n327 B.n326 10.6151
R1777 B.n326 B.n325 10.6151
R1778 B.n325 B.n283 10.6151
R1779 B.n319 B.n283 10.6151
R1780 B.n319 B.n318 10.6151
R1781 B.n318 B.n317 10.6151
R1782 B.n317 B.n285 10.6151
R1783 B.n311 B.n285 10.6151
R1784 B.n311 B.n310 10.6151
R1785 B.n310 B.n309 10.6151
R1786 B.n309 B.n287 10.6151
R1787 B.n303 B.n287 10.6151
R1788 B.n303 B.n302 10.6151
R1789 B.n302 B.n301 10.6151
R1790 B.n301 B.n289 10.6151
R1791 B.n295 B.n289 10.6151
R1792 B.n295 B.n294 10.6151
R1793 B.n294 B.n293 10.6151
R1794 B.n293 B.n223 10.6151
R1795 B.n529 B.n219 10.6151
R1796 B.n539 B.n219 10.6151
R1797 B.n540 B.n539 10.6151
R1798 B.n541 B.n540 10.6151
R1799 B.n541 B.n211 10.6151
R1800 B.n551 B.n211 10.6151
R1801 B.n552 B.n551 10.6151
R1802 B.n553 B.n552 10.6151
R1803 B.n553 B.n203 10.6151
R1804 B.n563 B.n203 10.6151
R1805 B.n564 B.n563 10.6151
R1806 B.n565 B.n564 10.6151
R1807 B.n565 B.n195 10.6151
R1808 B.n575 B.n195 10.6151
R1809 B.n576 B.n575 10.6151
R1810 B.n577 B.n576 10.6151
R1811 B.n577 B.n187 10.6151
R1812 B.n587 B.n187 10.6151
R1813 B.n588 B.n587 10.6151
R1814 B.n589 B.n588 10.6151
R1815 B.n589 B.n179 10.6151
R1816 B.n600 B.n179 10.6151
R1817 B.n601 B.n600 10.6151
R1818 B.n602 B.n601 10.6151
R1819 B.n602 B.n172 10.6151
R1820 B.n612 B.n172 10.6151
R1821 B.n613 B.n612 10.6151
R1822 B.n614 B.n613 10.6151
R1823 B.n614 B.n164 10.6151
R1824 B.n624 B.n164 10.6151
R1825 B.n625 B.n624 10.6151
R1826 B.n626 B.n625 10.6151
R1827 B.n626 B.n156 10.6151
R1828 B.n636 B.n156 10.6151
R1829 B.n637 B.n636 10.6151
R1830 B.n638 B.n637 10.6151
R1831 B.n638 B.n148 10.6151
R1832 B.n649 B.n148 10.6151
R1833 B.n650 B.n649 10.6151
R1834 B.n651 B.n650 10.6151
R1835 B.n651 B.n0 10.6151
R1836 B.n1031 B.n1 10.6151
R1837 B.n1031 B.n1030 10.6151
R1838 B.n1030 B.n1029 10.6151
R1839 B.n1029 B.n10 10.6151
R1840 B.n1023 B.n10 10.6151
R1841 B.n1023 B.n1022 10.6151
R1842 B.n1022 B.n1021 10.6151
R1843 B.n1021 B.n17 10.6151
R1844 B.n1015 B.n17 10.6151
R1845 B.n1015 B.n1014 10.6151
R1846 B.n1014 B.n1013 10.6151
R1847 B.n1013 B.n24 10.6151
R1848 B.n1007 B.n24 10.6151
R1849 B.n1007 B.n1006 10.6151
R1850 B.n1006 B.n1005 10.6151
R1851 B.n1005 B.n31 10.6151
R1852 B.n999 B.n31 10.6151
R1853 B.n999 B.n998 10.6151
R1854 B.n998 B.n997 10.6151
R1855 B.n997 B.n37 10.6151
R1856 B.n991 B.n37 10.6151
R1857 B.n991 B.n990 10.6151
R1858 B.n990 B.n989 10.6151
R1859 B.n989 B.n45 10.6151
R1860 B.n983 B.n45 10.6151
R1861 B.n983 B.n982 10.6151
R1862 B.n982 B.n981 10.6151
R1863 B.n981 B.n52 10.6151
R1864 B.n975 B.n52 10.6151
R1865 B.n975 B.n974 10.6151
R1866 B.n974 B.n973 10.6151
R1867 B.n973 B.n59 10.6151
R1868 B.n967 B.n59 10.6151
R1869 B.n967 B.n966 10.6151
R1870 B.n966 B.n965 10.6151
R1871 B.n965 B.n66 10.6151
R1872 B.n959 B.n66 10.6151
R1873 B.n959 B.n958 10.6151
R1874 B.n958 B.n957 10.6151
R1875 B.n957 B.n73 10.6151
R1876 B.n951 B.n73 10.6151
R1877 B.t2 B.n189 9.54606
R1878 B.n986 B.t7 9.54606
R1879 B.n110 B.n106 9.36635
R1880 B.n821 B.n820 9.36635
R1881 B.n420 B.n419 9.36635
R1882 B.n397 B.n263 9.36635
R1883 B.t9 B.n209 8.54126
R1884 B.n622 B.t5 8.54126
R1885 B.n1011 B.t4 8.54126
R1886 B.t16 B.n64 8.54126
R1887 B.n1037 B.n0 2.81026
R1888 B.n1037 B.n1 2.81026
R1889 B.n839 B.n110 1.24928
R1890 B.n822 B.n821 1.24928
R1891 B.n419 B.n418 1.24928
R1892 B.n401 B.n263 1.24928
R1893 B.n154 B.t0 0.502898
R1894 B.t1 B.n1026 0.502898
R1895 VN.n5 VN.t7 234.126
R1896 VN.n28 VN.t6 234.126
R1897 VN.n6 VN.t1 203.321
R1898 VN.n14 VN.t5 203.321
R1899 VN.n21 VN.t2 203.321
R1900 VN.n29 VN.t3 203.321
R1901 VN.n37 VN.t4 203.321
R1902 VN.n44 VN.t0 203.321
R1903 VN.n43 VN.n23 161.3
R1904 VN.n42 VN.n41 161.3
R1905 VN.n40 VN.n24 161.3
R1906 VN.n39 VN.n38 161.3
R1907 VN.n36 VN.n25 161.3
R1908 VN.n35 VN.n34 161.3
R1909 VN.n33 VN.n26 161.3
R1910 VN.n32 VN.n31 161.3
R1911 VN.n30 VN.n27 161.3
R1912 VN.n20 VN.n0 161.3
R1913 VN.n19 VN.n18 161.3
R1914 VN.n17 VN.n1 161.3
R1915 VN.n16 VN.n15 161.3
R1916 VN.n13 VN.n2 161.3
R1917 VN.n12 VN.n11 161.3
R1918 VN.n10 VN.n3 161.3
R1919 VN.n9 VN.n8 161.3
R1920 VN.n7 VN.n4 161.3
R1921 VN.n22 VN.n21 88.7756
R1922 VN.n45 VN.n44 88.7756
R1923 VN.n6 VN.n5 62.9301
R1924 VN.n29 VN.n28 62.9301
R1925 VN.n19 VN.n1 56.5617
R1926 VN.n42 VN.n24 56.5617
R1927 VN VN.n45 51.7785
R1928 VN.n8 VN.n3 40.577
R1929 VN.n12 VN.n3 40.577
R1930 VN.n31 VN.n26 40.577
R1931 VN.n35 VN.n26 40.577
R1932 VN.n8 VN.n7 24.5923
R1933 VN.n13 VN.n12 24.5923
R1934 VN.n15 VN.n1 24.5923
R1935 VN.n20 VN.n19 24.5923
R1936 VN.n31 VN.n30 24.5923
R1937 VN.n38 VN.n24 24.5923
R1938 VN.n36 VN.n35 24.5923
R1939 VN.n43 VN.n42 24.5923
R1940 VN.n21 VN.n20 22.1332
R1941 VN.n44 VN.n43 22.1332
R1942 VN.n15 VN.n14 17.2148
R1943 VN.n38 VN.n37 17.2148
R1944 VN.n28 VN.n27 12.9948
R1945 VN.n5 VN.n4 12.9948
R1946 VN.n7 VN.n6 7.37805
R1947 VN.n14 VN.n13 7.37805
R1948 VN.n30 VN.n29 7.37805
R1949 VN.n37 VN.n36 7.37805
R1950 VN.n45 VN.n23 0.278335
R1951 VN.n22 VN.n0 0.278335
R1952 VN.n41 VN.n23 0.189894
R1953 VN.n41 VN.n40 0.189894
R1954 VN.n40 VN.n39 0.189894
R1955 VN.n39 VN.n25 0.189894
R1956 VN.n34 VN.n25 0.189894
R1957 VN.n34 VN.n33 0.189894
R1958 VN.n33 VN.n32 0.189894
R1959 VN.n32 VN.n27 0.189894
R1960 VN.n9 VN.n4 0.189894
R1961 VN.n10 VN.n9 0.189894
R1962 VN.n11 VN.n10 0.189894
R1963 VN.n11 VN.n2 0.189894
R1964 VN.n16 VN.n2 0.189894
R1965 VN.n17 VN.n16 0.189894
R1966 VN.n18 VN.n17 0.189894
R1967 VN.n18 VN.n0 0.189894
R1968 VN VN.n22 0.153485
R1969 VDD2.n2 VDD2.n1 65.1763
R1970 VDD2.n2 VDD2.n0 65.1763
R1971 VDD2 VDD2.n5 65.1736
R1972 VDD2.n4 VDD2.n3 64.2406
R1973 VDD2.n4 VDD2.n2 46.9653
R1974 VDD2.n5 VDD2.t4 1.19184
R1975 VDD2.n5 VDD2.t1 1.19184
R1976 VDD2.n3 VDD2.t7 1.19184
R1977 VDD2.n3 VDD2.t3 1.19184
R1978 VDD2.n1 VDD2.t2 1.19184
R1979 VDD2.n1 VDD2.t5 1.19184
R1980 VDD2.n0 VDD2.t0 1.19184
R1981 VDD2.n0 VDD2.t6 1.19184
R1982 VDD2 VDD2.n4 1.05007
C0 VDD1 VTAIL 9.93112f
C1 VN VP 7.74335f
C2 VDD2 VP 0.453049f
C3 VTAIL VP 11.171401f
C4 VDD1 VP 11.4486f
C5 VN VDD2 11.147699f
C6 VN VTAIL 11.1573f
C7 VTAIL VDD2 9.981309f
C8 VN VDD1 0.151006f
C9 VDD1 VDD2 1.45017f
C10 VDD2 B 5.098616f
C11 VDD1 B 5.465209f
C12 VTAIL B 12.76652f
C13 VN B 13.54313f
C14 VP B 11.932442f
C15 VDD2.t0 B 0.322774f
C16 VDD2.t6 B 0.322774f
C17 VDD2.n0 B 2.94091f
C18 VDD2.t2 B 0.322774f
C19 VDD2.t5 B 0.322774f
C20 VDD2.n1 B 2.94091f
C21 VDD2.n2 B 3.14212f
C22 VDD2.t7 B 0.322774f
C23 VDD2.t3 B 0.322774f
C24 VDD2.n3 B 2.93458f
C25 VDD2.n4 B 3.02769f
C26 VDD2.t4 B 0.322774f
C27 VDD2.t1 B 0.322774f
C28 VDD2.n5 B 2.94087f
C29 VN.n0 B 0.033731f
C30 VN.t2 B 2.30063f
C31 VN.n1 B 0.040733f
C32 VN.n2 B 0.025586f
C33 VN.t5 B 2.30063f
C34 VN.n3 B 0.020665f
C35 VN.n4 B 0.190824f
C36 VN.t1 B 2.30063f
C37 VN.t7 B 2.42312f
C38 VN.n5 B 0.872832f
C39 VN.n6 B 0.861853f
C40 VN.n7 B 0.031051f
C41 VN.n8 B 0.050585f
C42 VN.n9 B 0.025586f
C43 VN.n10 B 0.025586f
C44 VN.n11 B 0.025586f
C45 VN.n12 B 0.050585f
C46 VN.n13 B 0.031051f
C47 VN.n14 B 0.805997f
C48 VN.n15 B 0.04042f
C49 VN.n16 B 0.025586f
C50 VN.n17 B 0.025586f
C51 VN.n18 B 0.025586f
C52 VN.n19 B 0.033654f
C53 VN.n20 B 0.045105f
C54 VN.n21 B 0.886287f
C55 VN.n22 B 0.029222f
C56 VN.n23 B 0.033731f
C57 VN.t0 B 2.30063f
C58 VN.n24 B 0.040733f
C59 VN.n25 B 0.025586f
C60 VN.t4 B 2.30063f
C61 VN.n26 B 0.020665f
C62 VN.n27 B 0.190824f
C63 VN.t3 B 2.30063f
C64 VN.t6 B 2.42312f
C65 VN.n28 B 0.872832f
C66 VN.n29 B 0.861853f
C67 VN.n30 B 0.031051f
C68 VN.n31 B 0.050585f
C69 VN.n32 B 0.025586f
C70 VN.n33 B 0.025586f
C71 VN.n34 B 0.025586f
C72 VN.n35 B 0.050585f
C73 VN.n36 B 0.031051f
C74 VN.n37 B 0.805997f
C75 VN.n38 B 0.04042f
C76 VN.n39 B 0.025586f
C77 VN.n40 B 0.025586f
C78 VN.n41 B 0.025586f
C79 VN.n42 B 0.033654f
C80 VN.n43 B 0.045105f
C81 VN.n44 B 0.886287f
C82 VN.n45 B 1.48724f
C83 VTAIL.t4 B 0.243845f
C84 VTAIL.t3 B 0.243845f
C85 VTAIL.n0 B 2.16544f
C86 VTAIL.n1 B 0.298891f
C87 VTAIL.t1 B 2.76726f
C88 VTAIL.n2 B 0.386725f
C89 VTAIL.t9 B 2.76726f
C90 VTAIL.n3 B 0.386725f
C91 VTAIL.t12 B 0.243845f
C92 VTAIL.t13 B 0.243845f
C93 VTAIL.n4 B 2.16544f
C94 VTAIL.n5 B 0.414029f
C95 VTAIL.t8 B 2.76726f
C96 VTAIL.n6 B 1.58659f
C97 VTAIL.t2 B 2.76727f
C98 VTAIL.n7 B 1.58659f
C99 VTAIL.t6 B 0.243845f
C100 VTAIL.t5 B 0.243845f
C101 VTAIL.n8 B 2.16544f
C102 VTAIL.n9 B 0.414026f
C103 VTAIL.t0 B 2.76727f
C104 VTAIL.n10 B 0.386722f
C105 VTAIL.t14 B 2.76727f
C106 VTAIL.n11 B 0.386722f
C107 VTAIL.t10 B 0.243845f
C108 VTAIL.t15 B 0.243845f
C109 VTAIL.n12 B 2.16544f
C110 VTAIL.n13 B 0.414026f
C111 VTAIL.t11 B 2.76726f
C112 VTAIL.n14 B 1.58659f
C113 VTAIL.t7 B 2.76726f
C114 VTAIL.n15 B 1.58311f
C115 VDD1.t6 B 0.324438f
C116 VDD1.t0 B 0.324438f
C117 VDD1.n0 B 2.95696f
C118 VDD1.t2 B 0.324438f
C119 VDD1.t4 B 0.324438f
C120 VDD1.n1 B 2.95607f
C121 VDD1.t5 B 0.324438f
C122 VDD1.t3 B 0.324438f
C123 VDD1.n2 B 2.95607f
C124 VDD1.n3 B 3.20993f
C125 VDD1.t7 B 0.324438f
C126 VDD1.t1 B 0.324438f
C127 VDD1.n4 B 2.94969f
C128 VDD1.n5 B 3.07367f
C129 VP.n0 B 0.034109f
C130 VP.t6 B 2.32643f
C131 VP.n1 B 0.04119f
C132 VP.n2 B 0.025873f
C133 VP.t2 B 2.32643f
C134 VP.n3 B 0.020897f
C135 VP.n4 B 0.025873f
C136 VP.t3 B 2.32643f
C137 VP.n5 B 0.04119f
C138 VP.n6 B 0.034109f
C139 VP.t7 B 2.32643f
C140 VP.n7 B 0.034109f
C141 VP.t4 B 2.32643f
C142 VP.n8 B 0.04119f
C143 VP.n9 B 0.025873f
C144 VP.t0 B 2.32643f
C145 VP.n10 B 0.020897f
C146 VP.n11 B 0.192963f
C147 VP.t5 B 2.32643f
C148 VP.t1 B 2.45029f
C149 VP.n12 B 0.882618f
C150 VP.n13 B 0.871516f
C151 VP.n14 B 0.031399f
C152 VP.n15 B 0.051152f
C153 VP.n16 B 0.025873f
C154 VP.n17 B 0.025873f
C155 VP.n18 B 0.025873f
C156 VP.n19 B 0.051152f
C157 VP.n20 B 0.031399f
C158 VP.n21 B 0.815034f
C159 VP.n22 B 0.040874f
C160 VP.n23 B 0.025873f
C161 VP.n24 B 0.025873f
C162 VP.n25 B 0.025873f
C163 VP.n26 B 0.034031f
C164 VP.n27 B 0.045611f
C165 VP.n28 B 0.896224f
C166 VP.n29 B 1.49008f
C167 VP.n30 B 1.50819f
C168 VP.n31 B 0.896224f
C169 VP.n32 B 0.045611f
C170 VP.n33 B 0.034031f
C171 VP.n34 B 0.025873f
C172 VP.n35 B 0.025873f
C173 VP.n36 B 0.025873f
C174 VP.n37 B 0.040874f
C175 VP.n38 B 0.815034f
C176 VP.n39 B 0.031399f
C177 VP.n40 B 0.051152f
C178 VP.n41 B 0.025873f
C179 VP.n42 B 0.025873f
C180 VP.n43 B 0.025873f
C181 VP.n44 B 0.051152f
C182 VP.n45 B 0.031399f
C183 VP.n46 B 0.815034f
C184 VP.n47 B 0.040874f
C185 VP.n48 B 0.025873f
C186 VP.n49 B 0.025873f
C187 VP.n50 B 0.025873f
C188 VP.n51 B 0.034031f
C189 VP.n52 B 0.045611f
C190 VP.n53 B 0.896224f
C191 VP.n54 B 0.029549f
.ends

