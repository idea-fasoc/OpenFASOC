* NGSPICE file created from diff_pair_sample_1125.ext - technology: sky130A

.subckt diff_pair_sample_1125 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t15 VP.t0 VDD1.t3 w_n4880_n3920# sky130_fd_pr__pfet_01v8 ad=5.7564 pd=30.3 as=2.4354 ps=15.09 w=14.76 l=3.58
X1 VDD1.t2 VP.t1 VTAIL.t14 w_n4880_n3920# sky130_fd_pr__pfet_01v8 ad=2.4354 pd=15.09 as=5.7564 ps=30.3 w=14.76 l=3.58
X2 B.t11 B.t9 B.t10 w_n4880_n3920# sky130_fd_pr__pfet_01v8 ad=5.7564 pd=30.3 as=0 ps=0 w=14.76 l=3.58
X3 VDD1.t5 VP.t2 VTAIL.t13 w_n4880_n3920# sky130_fd_pr__pfet_01v8 ad=2.4354 pd=15.09 as=2.4354 ps=15.09 w=14.76 l=3.58
X4 VTAIL.t12 VP.t3 VDD1.t4 w_n4880_n3920# sky130_fd_pr__pfet_01v8 ad=2.4354 pd=15.09 as=2.4354 ps=15.09 w=14.76 l=3.58
X5 VDD2.t7 VN.t0 VTAIL.t7 w_n4880_n3920# sky130_fd_pr__pfet_01v8 ad=2.4354 pd=15.09 as=5.7564 ps=30.3 w=14.76 l=3.58
X6 VTAIL.t4 VN.t1 VDD2.t6 w_n4880_n3920# sky130_fd_pr__pfet_01v8 ad=5.7564 pd=30.3 as=2.4354 ps=15.09 w=14.76 l=3.58
X7 VDD1.t1 VP.t4 VTAIL.t11 w_n4880_n3920# sky130_fd_pr__pfet_01v8 ad=2.4354 pd=15.09 as=2.4354 ps=15.09 w=14.76 l=3.58
X8 VDD2.t5 VN.t2 VTAIL.t3 w_n4880_n3920# sky130_fd_pr__pfet_01v8 ad=2.4354 pd=15.09 as=2.4354 ps=15.09 w=14.76 l=3.58
X9 B.t8 B.t6 B.t7 w_n4880_n3920# sky130_fd_pr__pfet_01v8 ad=5.7564 pd=30.3 as=0 ps=0 w=14.76 l=3.58
X10 VTAIL.t10 VP.t5 VDD1.t0 w_n4880_n3920# sky130_fd_pr__pfet_01v8 ad=2.4354 pd=15.09 as=2.4354 ps=15.09 w=14.76 l=3.58
X11 VTAIL.t2 VN.t3 VDD2.t4 w_n4880_n3920# sky130_fd_pr__pfet_01v8 ad=2.4354 pd=15.09 as=2.4354 ps=15.09 w=14.76 l=3.58
X12 B.t5 B.t3 B.t4 w_n4880_n3920# sky130_fd_pr__pfet_01v8 ad=5.7564 pd=30.3 as=0 ps=0 w=14.76 l=3.58
X13 VDD2.t3 VN.t4 VTAIL.t5 w_n4880_n3920# sky130_fd_pr__pfet_01v8 ad=2.4354 pd=15.09 as=5.7564 ps=30.3 w=14.76 l=3.58
X14 VTAIL.t1 VN.t5 VDD2.t2 w_n4880_n3920# sky130_fd_pr__pfet_01v8 ad=5.7564 pd=30.3 as=2.4354 ps=15.09 w=14.76 l=3.58
X15 VDD2.t1 VN.t6 VTAIL.t6 w_n4880_n3920# sky130_fd_pr__pfet_01v8 ad=2.4354 pd=15.09 as=2.4354 ps=15.09 w=14.76 l=3.58
X16 VDD1.t7 VP.t6 VTAIL.t9 w_n4880_n3920# sky130_fd_pr__pfet_01v8 ad=2.4354 pd=15.09 as=5.7564 ps=30.3 w=14.76 l=3.58
X17 B.t2 B.t0 B.t1 w_n4880_n3920# sky130_fd_pr__pfet_01v8 ad=5.7564 pd=30.3 as=0 ps=0 w=14.76 l=3.58
X18 VTAIL.t0 VN.t7 VDD2.t0 w_n4880_n3920# sky130_fd_pr__pfet_01v8 ad=2.4354 pd=15.09 as=2.4354 ps=15.09 w=14.76 l=3.58
X19 VTAIL.t8 VP.t7 VDD1.t6 w_n4880_n3920# sky130_fd_pr__pfet_01v8 ad=5.7564 pd=30.3 as=2.4354 ps=15.09 w=14.76 l=3.58
R0 VP.n24 VP.n21 161.3
R1 VP.n26 VP.n25 161.3
R2 VP.n27 VP.n20 161.3
R3 VP.n29 VP.n28 161.3
R4 VP.n30 VP.n19 161.3
R5 VP.n32 VP.n31 161.3
R6 VP.n33 VP.n18 161.3
R7 VP.n36 VP.n35 161.3
R8 VP.n37 VP.n17 161.3
R9 VP.n39 VP.n38 161.3
R10 VP.n40 VP.n16 161.3
R11 VP.n42 VP.n41 161.3
R12 VP.n43 VP.n15 161.3
R13 VP.n45 VP.n44 161.3
R14 VP.n46 VP.n14 161.3
R15 VP.n48 VP.n47 161.3
R16 VP.n89 VP.n88 161.3
R17 VP.n87 VP.n1 161.3
R18 VP.n86 VP.n85 161.3
R19 VP.n84 VP.n2 161.3
R20 VP.n83 VP.n82 161.3
R21 VP.n81 VP.n3 161.3
R22 VP.n80 VP.n79 161.3
R23 VP.n78 VP.n4 161.3
R24 VP.n77 VP.n76 161.3
R25 VP.n74 VP.n5 161.3
R26 VP.n73 VP.n72 161.3
R27 VP.n71 VP.n6 161.3
R28 VP.n70 VP.n69 161.3
R29 VP.n68 VP.n7 161.3
R30 VP.n67 VP.n66 161.3
R31 VP.n65 VP.n8 161.3
R32 VP.n64 VP.n63 161.3
R33 VP.n61 VP.n9 161.3
R34 VP.n60 VP.n59 161.3
R35 VP.n58 VP.n10 161.3
R36 VP.n57 VP.n56 161.3
R37 VP.n55 VP.n11 161.3
R38 VP.n54 VP.n53 161.3
R39 VP.n52 VP.n12 161.3
R40 VP.n23 VP.t0 132.018
R41 VP.n50 VP.t7 99.3625
R42 VP.n62 VP.t2 99.3625
R43 VP.n75 VP.t3 99.3625
R44 VP.n0 VP.t1 99.3625
R45 VP.n13 VP.t6 99.3625
R46 VP.n34 VP.t5 99.3625
R47 VP.n22 VP.t4 99.3625
R48 VP.n51 VP.n50 84.5894
R49 VP.n90 VP.n0 84.5894
R50 VP.n49 VP.n13 84.5894
R51 VP.n23 VP.n22 64.6381
R52 VP.n51 VP.n49 57.6132
R53 VP.n69 VP.n6 56.5617
R54 VP.n28 VP.n19 56.5617
R55 VP.n56 VP.n10 56.0773
R56 VP.n82 VP.n2 56.0773
R57 VP.n41 VP.n15 56.0773
R58 VP.n60 VP.n10 25.0767
R59 VP.n82 VP.n81 25.0767
R60 VP.n41 VP.n40 25.0767
R61 VP.n54 VP.n12 24.5923
R62 VP.n55 VP.n54 24.5923
R63 VP.n56 VP.n55 24.5923
R64 VP.n61 VP.n60 24.5923
R65 VP.n63 VP.n61 24.5923
R66 VP.n67 VP.n8 24.5923
R67 VP.n68 VP.n67 24.5923
R68 VP.n69 VP.n68 24.5923
R69 VP.n73 VP.n6 24.5923
R70 VP.n74 VP.n73 24.5923
R71 VP.n76 VP.n74 24.5923
R72 VP.n80 VP.n4 24.5923
R73 VP.n81 VP.n80 24.5923
R74 VP.n86 VP.n2 24.5923
R75 VP.n87 VP.n86 24.5923
R76 VP.n88 VP.n87 24.5923
R77 VP.n45 VP.n15 24.5923
R78 VP.n46 VP.n45 24.5923
R79 VP.n47 VP.n46 24.5923
R80 VP.n32 VP.n19 24.5923
R81 VP.n33 VP.n32 24.5923
R82 VP.n35 VP.n33 24.5923
R83 VP.n39 VP.n17 24.5923
R84 VP.n40 VP.n39 24.5923
R85 VP.n26 VP.n21 24.5923
R86 VP.n27 VP.n26 24.5923
R87 VP.n28 VP.n27 24.5923
R88 VP.n63 VP.n62 14.5097
R89 VP.n75 VP.n4 14.5097
R90 VP.n34 VP.n17 14.5097
R91 VP.n62 VP.n8 10.0832
R92 VP.n76 VP.n75 10.0832
R93 VP.n35 VP.n34 10.0832
R94 VP.n22 VP.n21 10.0832
R95 VP.n50 VP.n12 5.65662
R96 VP.n88 VP.n0 5.65662
R97 VP.n47 VP.n13 5.65662
R98 VP.n24 VP.n23 3.28578
R99 VP.n49 VP.n48 0.354861
R100 VP.n52 VP.n51 0.354861
R101 VP.n90 VP.n89 0.354861
R102 VP VP.n90 0.267071
R103 VP.n25 VP.n24 0.189894
R104 VP.n25 VP.n20 0.189894
R105 VP.n29 VP.n20 0.189894
R106 VP.n30 VP.n29 0.189894
R107 VP.n31 VP.n30 0.189894
R108 VP.n31 VP.n18 0.189894
R109 VP.n36 VP.n18 0.189894
R110 VP.n37 VP.n36 0.189894
R111 VP.n38 VP.n37 0.189894
R112 VP.n38 VP.n16 0.189894
R113 VP.n42 VP.n16 0.189894
R114 VP.n43 VP.n42 0.189894
R115 VP.n44 VP.n43 0.189894
R116 VP.n44 VP.n14 0.189894
R117 VP.n48 VP.n14 0.189894
R118 VP.n53 VP.n52 0.189894
R119 VP.n53 VP.n11 0.189894
R120 VP.n57 VP.n11 0.189894
R121 VP.n58 VP.n57 0.189894
R122 VP.n59 VP.n58 0.189894
R123 VP.n59 VP.n9 0.189894
R124 VP.n64 VP.n9 0.189894
R125 VP.n65 VP.n64 0.189894
R126 VP.n66 VP.n65 0.189894
R127 VP.n66 VP.n7 0.189894
R128 VP.n70 VP.n7 0.189894
R129 VP.n71 VP.n70 0.189894
R130 VP.n72 VP.n71 0.189894
R131 VP.n72 VP.n5 0.189894
R132 VP.n77 VP.n5 0.189894
R133 VP.n78 VP.n77 0.189894
R134 VP.n79 VP.n78 0.189894
R135 VP.n79 VP.n3 0.189894
R136 VP.n83 VP.n3 0.189894
R137 VP.n84 VP.n83 0.189894
R138 VP.n85 VP.n84 0.189894
R139 VP.n85 VP.n1 0.189894
R140 VP.n89 VP.n1 0.189894
R141 VDD1 VDD1.n0 74.8374
R142 VDD1.n3 VDD1.n2 74.7237
R143 VDD1.n3 VDD1.n1 74.7237
R144 VDD1.n5 VDD1.n4 73.0936
R145 VDD1.n5 VDD1.n3 52.1906
R146 VDD1.n4 VDD1.t0 2.20274
R147 VDD1.n4 VDD1.t7 2.20274
R148 VDD1.n0 VDD1.t3 2.20274
R149 VDD1.n0 VDD1.t1 2.20274
R150 VDD1.n2 VDD1.t4 2.20274
R151 VDD1.n2 VDD1.t2 2.20274
R152 VDD1.n1 VDD1.t6 2.20274
R153 VDD1.n1 VDD1.t5 2.20274
R154 VDD1 VDD1.n5 1.62766
R155 VTAIL.n658 VTAIL.n582 756.745
R156 VTAIL.n78 VTAIL.n2 756.745
R157 VTAIL.n160 VTAIL.n84 756.745
R158 VTAIL.n244 VTAIL.n168 756.745
R159 VTAIL.n576 VTAIL.n500 756.745
R160 VTAIL.n492 VTAIL.n416 756.745
R161 VTAIL.n410 VTAIL.n334 756.745
R162 VTAIL.n326 VTAIL.n250 756.745
R163 VTAIL.n609 VTAIL.n608 585
R164 VTAIL.n606 VTAIL.n605 585
R165 VTAIL.n615 VTAIL.n614 585
R166 VTAIL.n617 VTAIL.n616 585
R167 VTAIL.n602 VTAIL.n601 585
R168 VTAIL.n623 VTAIL.n622 585
R169 VTAIL.n625 VTAIL.n624 585
R170 VTAIL.n598 VTAIL.n597 585
R171 VTAIL.n631 VTAIL.n630 585
R172 VTAIL.n633 VTAIL.n632 585
R173 VTAIL.n594 VTAIL.n593 585
R174 VTAIL.n639 VTAIL.n638 585
R175 VTAIL.n641 VTAIL.n640 585
R176 VTAIL.n590 VTAIL.n589 585
R177 VTAIL.n647 VTAIL.n646 585
R178 VTAIL.n650 VTAIL.n649 585
R179 VTAIL.n648 VTAIL.n586 585
R180 VTAIL.n655 VTAIL.n585 585
R181 VTAIL.n657 VTAIL.n656 585
R182 VTAIL.n659 VTAIL.n658 585
R183 VTAIL.n29 VTAIL.n28 585
R184 VTAIL.n26 VTAIL.n25 585
R185 VTAIL.n35 VTAIL.n34 585
R186 VTAIL.n37 VTAIL.n36 585
R187 VTAIL.n22 VTAIL.n21 585
R188 VTAIL.n43 VTAIL.n42 585
R189 VTAIL.n45 VTAIL.n44 585
R190 VTAIL.n18 VTAIL.n17 585
R191 VTAIL.n51 VTAIL.n50 585
R192 VTAIL.n53 VTAIL.n52 585
R193 VTAIL.n14 VTAIL.n13 585
R194 VTAIL.n59 VTAIL.n58 585
R195 VTAIL.n61 VTAIL.n60 585
R196 VTAIL.n10 VTAIL.n9 585
R197 VTAIL.n67 VTAIL.n66 585
R198 VTAIL.n70 VTAIL.n69 585
R199 VTAIL.n68 VTAIL.n6 585
R200 VTAIL.n75 VTAIL.n5 585
R201 VTAIL.n77 VTAIL.n76 585
R202 VTAIL.n79 VTAIL.n78 585
R203 VTAIL.n111 VTAIL.n110 585
R204 VTAIL.n108 VTAIL.n107 585
R205 VTAIL.n117 VTAIL.n116 585
R206 VTAIL.n119 VTAIL.n118 585
R207 VTAIL.n104 VTAIL.n103 585
R208 VTAIL.n125 VTAIL.n124 585
R209 VTAIL.n127 VTAIL.n126 585
R210 VTAIL.n100 VTAIL.n99 585
R211 VTAIL.n133 VTAIL.n132 585
R212 VTAIL.n135 VTAIL.n134 585
R213 VTAIL.n96 VTAIL.n95 585
R214 VTAIL.n141 VTAIL.n140 585
R215 VTAIL.n143 VTAIL.n142 585
R216 VTAIL.n92 VTAIL.n91 585
R217 VTAIL.n149 VTAIL.n148 585
R218 VTAIL.n152 VTAIL.n151 585
R219 VTAIL.n150 VTAIL.n88 585
R220 VTAIL.n157 VTAIL.n87 585
R221 VTAIL.n159 VTAIL.n158 585
R222 VTAIL.n161 VTAIL.n160 585
R223 VTAIL.n195 VTAIL.n194 585
R224 VTAIL.n192 VTAIL.n191 585
R225 VTAIL.n201 VTAIL.n200 585
R226 VTAIL.n203 VTAIL.n202 585
R227 VTAIL.n188 VTAIL.n187 585
R228 VTAIL.n209 VTAIL.n208 585
R229 VTAIL.n211 VTAIL.n210 585
R230 VTAIL.n184 VTAIL.n183 585
R231 VTAIL.n217 VTAIL.n216 585
R232 VTAIL.n219 VTAIL.n218 585
R233 VTAIL.n180 VTAIL.n179 585
R234 VTAIL.n225 VTAIL.n224 585
R235 VTAIL.n227 VTAIL.n226 585
R236 VTAIL.n176 VTAIL.n175 585
R237 VTAIL.n233 VTAIL.n232 585
R238 VTAIL.n236 VTAIL.n235 585
R239 VTAIL.n234 VTAIL.n172 585
R240 VTAIL.n241 VTAIL.n171 585
R241 VTAIL.n243 VTAIL.n242 585
R242 VTAIL.n245 VTAIL.n244 585
R243 VTAIL.n577 VTAIL.n576 585
R244 VTAIL.n575 VTAIL.n574 585
R245 VTAIL.n573 VTAIL.n503 585
R246 VTAIL.n507 VTAIL.n504 585
R247 VTAIL.n568 VTAIL.n567 585
R248 VTAIL.n566 VTAIL.n565 585
R249 VTAIL.n509 VTAIL.n508 585
R250 VTAIL.n560 VTAIL.n559 585
R251 VTAIL.n558 VTAIL.n557 585
R252 VTAIL.n513 VTAIL.n512 585
R253 VTAIL.n552 VTAIL.n551 585
R254 VTAIL.n550 VTAIL.n549 585
R255 VTAIL.n517 VTAIL.n516 585
R256 VTAIL.n544 VTAIL.n543 585
R257 VTAIL.n542 VTAIL.n541 585
R258 VTAIL.n521 VTAIL.n520 585
R259 VTAIL.n536 VTAIL.n535 585
R260 VTAIL.n534 VTAIL.n533 585
R261 VTAIL.n525 VTAIL.n524 585
R262 VTAIL.n528 VTAIL.n527 585
R263 VTAIL.n493 VTAIL.n492 585
R264 VTAIL.n491 VTAIL.n490 585
R265 VTAIL.n489 VTAIL.n419 585
R266 VTAIL.n423 VTAIL.n420 585
R267 VTAIL.n484 VTAIL.n483 585
R268 VTAIL.n482 VTAIL.n481 585
R269 VTAIL.n425 VTAIL.n424 585
R270 VTAIL.n476 VTAIL.n475 585
R271 VTAIL.n474 VTAIL.n473 585
R272 VTAIL.n429 VTAIL.n428 585
R273 VTAIL.n468 VTAIL.n467 585
R274 VTAIL.n466 VTAIL.n465 585
R275 VTAIL.n433 VTAIL.n432 585
R276 VTAIL.n460 VTAIL.n459 585
R277 VTAIL.n458 VTAIL.n457 585
R278 VTAIL.n437 VTAIL.n436 585
R279 VTAIL.n452 VTAIL.n451 585
R280 VTAIL.n450 VTAIL.n449 585
R281 VTAIL.n441 VTAIL.n440 585
R282 VTAIL.n444 VTAIL.n443 585
R283 VTAIL.n411 VTAIL.n410 585
R284 VTAIL.n409 VTAIL.n408 585
R285 VTAIL.n407 VTAIL.n337 585
R286 VTAIL.n341 VTAIL.n338 585
R287 VTAIL.n402 VTAIL.n401 585
R288 VTAIL.n400 VTAIL.n399 585
R289 VTAIL.n343 VTAIL.n342 585
R290 VTAIL.n394 VTAIL.n393 585
R291 VTAIL.n392 VTAIL.n391 585
R292 VTAIL.n347 VTAIL.n346 585
R293 VTAIL.n386 VTAIL.n385 585
R294 VTAIL.n384 VTAIL.n383 585
R295 VTAIL.n351 VTAIL.n350 585
R296 VTAIL.n378 VTAIL.n377 585
R297 VTAIL.n376 VTAIL.n375 585
R298 VTAIL.n355 VTAIL.n354 585
R299 VTAIL.n370 VTAIL.n369 585
R300 VTAIL.n368 VTAIL.n367 585
R301 VTAIL.n359 VTAIL.n358 585
R302 VTAIL.n362 VTAIL.n361 585
R303 VTAIL.n327 VTAIL.n326 585
R304 VTAIL.n325 VTAIL.n324 585
R305 VTAIL.n323 VTAIL.n253 585
R306 VTAIL.n257 VTAIL.n254 585
R307 VTAIL.n318 VTAIL.n317 585
R308 VTAIL.n316 VTAIL.n315 585
R309 VTAIL.n259 VTAIL.n258 585
R310 VTAIL.n310 VTAIL.n309 585
R311 VTAIL.n308 VTAIL.n307 585
R312 VTAIL.n263 VTAIL.n262 585
R313 VTAIL.n302 VTAIL.n301 585
R314 VTAIL.n300 VTAIL.n299 585
R315 VTAIL.n267 VTAIL.n266 585
R316 VTAIL.n294 VTAIL.n293 585
R317 VTAIL.n292 VTAIL.n291 585
R318 VTAIL.n271 VTAIL.n270 585
R319 VTAIL.n286 VTAIL.n285 585
R320 VTAIL.n284 VTAIL.n283 585
R321 VTAIL.n275 VTAIL.n274 585
R322 VTAIL.n278 VTAIL.n277 585
R323 VTAIL.t9 VTAIL.n526 327.466
R324 VTAIL.t15 VTAIL.n442 327.466
R325 VTAIL.t7 VTAIL.n360 327.466
R326 VTAIL.t4 VTAIL.n276 327.466
R327 VTAIL.t5 VTAIL.n607 327.466
R328 VTAIL.t1 VTAIL.n27 327.466
R329 VTAIL.t14 VTAIL.n109 327.466
R330 VTAIL.t8 VTAIL.n193 327.466
R331 VTAIL.n608 VTAIL.n605 171.744
R332 VTAIL.n615 VTAIL.n605 171.744
R333 VTAIL.n616 VTAIL.n615 171.744
R334 VTAIL.n616 VTAIL.n601 171.744
R335 VTAIL.n623 VTAIL.n601 171.744
R336 VTAIL.n624 VTAIL.n623 171.744
R337 VTAIL.n624 VTAIL.n597 171.744
R338 VTAIL.n631 VTAIL.n597 171.744
R339 VTAIL.n632 VTAIL.n631 171.744
R340 VTAIL.n632 VTAIL.n593 171.744
R341 VTAIL.n639 VTAIL.n593 171.744
R342 VTAIL.n640 VTAIL.n639 171.744
R343 VTAIL.n640 VTAIL.n589 171.744
R344 VTAIL.n647 VTAIL.n589 171.744
R345 VTAIL.n649 VTAIL.n647 171.744
R346 VTAIL.n649 VTAIL.n648 171.744
R347 VTAIL.n648 VTAIL.n585 171.744
R348 VTAIL.n657 VTAIL.n585 171.744
R349 VTAIL.n658 VTAIL.n657 171.744
R350 VTAIL.n28 VTAIL.n25 171.744
R351 VTAIL.n35 VTAIL.n25 171.744
R352 VTAIL.n36 VTAIL.n35 171.744
R353 VTAIL.n36 VTAIL.n21 171.744
R354 VTAIL.n43 VTAIL.n21 171.744
R355 VTAIL.n44 VTAIL.n43 171.744
R356 VTAIL.n44 VTAIL.n17 171.744
R357 VTAIL.n51 VTAIL.n17 171.744
R358 VTAIL.n52 VTAIL.n51 171.744
R359 VTAIL.n52 VTAIL.n13 171.744
R360 VTAIL.n59 VTAIL.n13 171.744
R361 VTAIL.n60 VTAIL.n59 171.744
R362 VTAIL.n60 VTAIL.n9 171.744
R363 VTAIL.n67 VTAIL.n9 171.744
R364 VTAIL.n69 VTAIL.n67 171.744
R365 VTAIL.n69 VTAIL.n68 171.744
R366 VTAIL.n68 VTAIL.n5 171.744
R367 VTAIL.n77 VTAIL.n5 171.744
R368 VTAIL.n78 VTAIL.n77 171.744
R369 VTAIL.n110 VTAIL.n107 171.744
R370 VTAIL.n117 VTAIL.n107 171.744
R371 VTAIL.n118 VTAIL.n117 171.744
R372 VTAIL.n118 VTAIL.n103 171.744
R373 VTAIL.n125 VTAIL.n103 171.744
R374 VTAIL.n126 VTAIL.n125 171.744
R375 VTAIL.n126 VTAIL.n99 171.744
R376 VTAIL.n133 VTAIL.n99 171.744
R377 VTAIL.n134 VTAIL.n133 171.744
R378 VTAIL.n134 VTAIL.n95 171.744
R379 VTAIL.n141 VTAIL.n95 171.744
R380 VTAIL.n142 VTAIL.n141 171.744
R381 VTAIL.n142 VTAIL.n91 171.744
R382 VTAIL.n149 VTAIL.n91 171.744
R383 VTAIL.n151 VTAIL.n149 171.744
R384 VTAIL.n151 VTAIL.n150 171.744
R385 VTAIL.n150 VTAIL.n87 171.744
R386 VTAIL.n159 VTAIL.n87 171.744
R387 VTAIL.n160 VTAIL.n159 171.744
R388 VTAIL.n194 VTAIL.n191 171.744
R389 VTAIL.n201 VTAIL.n191 171.744
R390 VTAIL.n202 VTAIL.n201 171.744
R391 VTAIL.n202 VTAIL.n187 171.744
R392 VTAIL.n209 VTAIL.n187 171.744
R393 VTAIL.n210 VTAIL.n209 171.744
R394 VTAIL.n210 VTAIL.n183 171.744
R395 VTAIL.n217 VTAIL.n183 171.744
R396 VTAIL.n218 VTAIL.n217 171.744
R397 VTAIL.n218 VTAIL.n179 171.744
R398 VTAIL.n225 VTAIL.n179 171.744
R399 VTAIL.n226 VTAIL.n225 171.744
R400 VTAIL.n226 VTAIL.n175 171.744
R401 VTAIL.n233 VTAIL.n175 171.744
R402 VTAIL.n235 VTAIL.n233 171.744
R403 VTAIL.n235 VTAIL.n234 171.744
R404 VTAIL.n234 VTAIL.n171 171.744
R405 VTAIL.n243 VTAIL.n171 171.744
R406 VTAIL.n244 VTAIL.n243 171.744
R407 VTAIL.n576 VTAIL.n575 171.744
R408 VTAIL.n575 VTAIL.n503 171.744
R409 VTAIL.n507 VTAIL.n503 171.744
R410 VTAIL.n567 VTAIL.n507 171.744
R411 VTAIL.n567 VTAIL.n566 171.744
R412 VTAIL.n566 VTAIL.n508 171.744
R413 VTAIL.n559 VTAIL.n508 171.744
R414 VTAIL.n559 VTAIL.n558 171.744
R415 VTAIL.n558 VTAIL.n512 171.744
R416 VTAIL.n551 VTAIL.n512 171.744
R417 VTAIL.n551 VTAIL.n550 171.744
R418 VTAIL.n550 VTAIL.n516 171.744
R419 VTAIL.n543 VTAIL.n516 171.744
R420 VTAIL.n543 VTAIL.n542 171.744
R421 VTAIL.n542 VTAIL.n520 171.744
R422 VTAIL.n535 VTAIL.n520 171.744
R423 VTAIL.n535 VTAIL.n534 171.744
R424 VTAIL.n534 VTAIL.n524 171.744
R425 VTAIL.n527 VTAIL.n524 171.744
R426 VTAIL.n492 VTAIL.n491 171.744
R427 VTAIL.n491 VTAIL.n419 171.744
R428 VTAIL.n423 VTAIL.n419 171.744
R429 VTAIL.n483 VTAIL.n423 171.744
R430 VTAIL.n483 VTAIL.n482 171.744
R431 VTAIL.n482 VTAIL.n424 171.744
R432 VTAIL.n475 VTAIL.n424 171.744
R433 VTAIL.n475 VTAIL.n474 171.744
R434 VTAIL.n474 VTAIL.n428 171.744
R435 VTAIL.n467 VTAIL.n428 171.744
R436 VTAIL.n467 VTAIL.n466 171.744
R437 VTAIL.n466 VTAIL.n432 171.744
R438 VTAIL.n459 VTAIL.n432 171.744
R439 VTAIL.n459 VTAIL.n458 171.744
R440 VTAIL.n458 VTAIL.n436 171.744
R441 VTAIL.n451 VTAIL.n436 171.744
R442 VTAIL.n451 VTAIL.n450 171.744
R443 VTAIL.n450 VTAIL.n440 171.744
R444 VTAIL.n443 VTAIL.n440 171.744
R445 VTAIL.n410 VTAIL.n409 171.744
R446 VTAIL.n409 VTAIL.n337 171.744
R447 VTAIL.n341 VTAIL.n337 171.744
R448 VTAIL.n401 VTAIL.n341 171.744
R449 VTAIL.n401 VTAIL.n400 171.744
R450 VTAIL.n400 VTAIL.n342 171.744
R451 VTAIL.n393 VTAIL.n342 171.744
R452 VTAIL.n393 VTAIL.n392 171.744
R453 VTAIL.n392 VTAIL.n346 171.744
R454 VTAIL.n385 VTAIL.n346 171.744
R455 VTAIL.n385 VTAIL.n384 171.744
R456 VTAIL.n384 VTAIL.n350 171.744
R457 VTAIL.n377 VTAIL.n350 171.744
R458 VTAIL.n377 VTAIL.n376 171.744
R459 VTAIL.n376 VTAIL.n354 171.744
R460 VTAIL.n369 VTAIL.n354 171.744
R461 VTAIL.n369 VTAIL.n368 171.744
R462 VTAIL.n368 VTAIL.n358 171.744
R463 VTAIL.n361 VTAIL.n358 171.744
R464 VTAIL.n326 VTAIL.n325 171.744
R465 VTAIL.n325 VTAIL.n253 171.744
R466 VTAIL.n257 VTAIL.n253 171.744
R467 VTAIL.n317 VTAIL.n257 171.744
R468 VTAIL.n317 VTAIL.n316 171.744
R469 VTAIL.n316 VTAIL.n258 171.744
R470 VTAIL.n309 VTAIL.n258 171.744
R471 VTAIL.n309 VTAIL.n308 171.744
R472 VTAIL.n308 VTAIL.n262 171.744
R473 VTAIL.n301 VTAIL.n262 171.744
R474 VTAIL.n301 VTAIL.n300 171.744
R475 VTAIL.n300 VTAIL.n266 171.744
R476 VTAIL.n293 VTAIL.n266 171.744
R477 VTAIL.n293 VTAIL.n292 171.744
R478 VTAIL.n292 VTAIL.n270 171.744
R479 VTAIL.n285 VTAIL.n270 171.744
R480 VTAIL.n285 VTAIL.n284 171.744
R481 VTAIL.n284 VTAIL.n274 171.744
R482 VTAIL.n277 VTAIL.n274 171.744
R483 VTAIL.n608 VTAIL.t5 85.8723
R484 VTAIL.n28 VTAIL.t1 85.8723
R485 VTAIL.n110 VTAIL.t14 85.8723
R486 VTAIL.n194 VTAIL.t8 85.8723
R487 VTAIL.n527 VTAIL.t9 85.8723
R488 VTAIL.n443 VTAIL.t15 85.8723
R489 VTAIL.n361 VTAIL.t7 85.8723
R490 VTAIL.n277 VTAIL.t4 85.8723
R491 VTAIL.n499 VTAIL.n498 56.4151
R492 VTAIL.n333 VTAIL.n332 56.4151
R493 VTAIL.n1 VTAIL.n0 56.4149
R494 VTAIL.n167 VTAIL.n166 56.4149
R495 VTAIL.n663 VTAIL.n662 34.5126
R496 VTAIL.n83 VTAIL.n82 34.5126
R497 VTAIL.n165 VTAIL.n164 34.5126
R498 VTAIL.n249 VTAIL.n248 34.5126
R499 VTAIL.n581 VTAIL.n580 34.5126
R500 VTAIL.n497 VTAIL.n496 34.5126
R501 VTAIL.n415 VTAIL.n414 34.5126
R502 VTAIL.n331 VTAIL.n330 34.5126
R503 VTAIL.n663 VTAIL.n581 28.4617
R504 VTAIL.n331 VTAIL.n249 28.4617
R505 VTAIL.n609 VTAIL.n607 16.3895
R506 VTAIL.n29 VTAIL.n27 16.3895
R507 VTAIL.n111 VTAIL.n109 16.3895
R508 VTAIL.n195 VTAIL.n193 16.3895
R509 VTAIL.n528 VTAIL.n526 16.3895
R510 VTAIL.n444 VTAIL.n442 16.3895
R511 VTAIL.n362 VTAIL.n360 16.3895
R512 VTAIL.n278 VTAIL.n276 16.3895
R513 VTAIL.n656 VTAIL.n655 13.1884
R514 VTAIL.n76 VTAIL.n75 13.1884
R515 VTAIL.n158 VTAIL.n157 13.1884
R516 VTAIL.n242 VTAIL.n241 13.1884
R517 VTAIL.n574 VTAIL.n573 13.1884
R518 VTAIL.n490 VTAIL.n489 13.1884
R519 VTAIL.n408 VTAIL.n407 13.1884
R520 VTAIL.n324 VTAIL.n323 13.1884
R521 VTAIL.n610 VTAIL.n606 12.8005
R522 VTAIL.n654 VTAIL.n586 12.8005
R523 VTAIL.n659 VTAIL.n584 12.8005
R524 VTAIL.n30 VTAIL.n26 12.8005
R525 VTAIL.n74 VTAIL.n6 12.8005
R526 VTAIL.n79 VTAIL.n4 12.8005
R527 VTAIL.n112 VTAIL.n108 12.8005
R528 VTAIL.n156 VTAIL.n88 12.8005
R529 VTAIL.n161 VTAIL.n86 12.8005
R530 VTAIL.n196 VTAIL.n192 12.8005
R531 VTAIL.n240 VTAIL.n172 12.8005
R532 VTAIL.n245 VTAIL.n170 12.8005
R533 VTAIL.n577 VTAIL.n502 12.8005
R534 VTAIL.n572 VTAIL.n504 12.8005
R535 VTAIL.n529 VTAIL.n525 12.8005
R536 VTAIL.n493 VTAIL.n418 12.8005
R537 VTAIL.n488 VTAIL.n420 12.8005
R538 VTAIL.n445 VTAIL.n441 12.8005
R539 VTAIL.n411 VTAIL.n336 12.8005
R540 VTAIL.n406 VTAIL.n338 12.8005
R541 VTAIL.n363 VTAIL.n359 12.8005
R542 VTAIL.n327 VTAIL.n252 12.8005
R543 VTAIL.n322 VTAIL.n254 12.8005
R544 VTAIL.n279 VTAIL.n275 12.8005
R545 VTAIL.n614 VTAIL.n613 12.0247
R546 VTAIL.n651 VTAIL.n650 12.0247
R547 VTAIL.n660 VTAIL.n582 12.0247
R548 VTAIL.n34 VTAIL.n33 12.0247
R549 VTAIL.n71 VTAIL.n70 12.0247
R550 VTAIL.n80 VTAIL.n2 12.0247
R551 VTAIL.n116 VTAIL.n115 12.0247
R552 VTAIL.n153 VTAIL.n152 12.0247
R553 VTAIL.n162 VTAIL.n84 12.0247
R554 VTAIL.n200 VTAIL.n199 12.0247
R555 VTAIL.n237 VTAIL.n236 12.0247
R556 VTAIL.n246 VTAIL.n168 12.0247
R557 VTAIL.n578 VTAIL.n500 12.0247
R558 VTAIL.n569 VTAIL.n568 12.0247
R559 VTAIL.n533 VTAIL.n532 12.0247
R560 VTAIL.n494 VTAIL.n416 12.0247
R561 VTAIL.n485 VTAIL.n484 12.0247
R562 VTAIL.n449 VTAIL.n448 12.0247
R563 VTAIL.n412 VTAIL.n334 12.0247
R564 VTAIL.n403 VTAIL.n402 12.0247
R565 VTAIL.n367 VTAIL.n366 12.0247
R566 VTAIL.n328 VTAIL.n250 12.0247
R567 VTAIL.n319 VTAIL.n318 12.0247
R568 VTAIL.n283 VTAIL.n282 12.0247
R569 VTAIL.n617 VTAIL.n604 11.249
R570 VTAIL.n646 VTAIL.n588 11.249
R571 VTAIL.n37 VTAIL.n24 11.249
R572 VTAIL.n66 VTAIL.n8 11.249
R573 VTAIL.n119 VTAIL.n106 11.249
R574 VTAIL.n148 VTAIL.n90 11.249
R575 VTAIL.n203 VTAIL.n190 11.249
R576 VTAIL.n232 VTAIL.n174 11.249
R577 VTAIL.n565 VTAIL.n506 11.249
R578 VTAIL.n536 VTAIL.n523 11.249
R579 VTAIL.n481 VTAIL.n422 11.249
R580 VTAIL.n452 VTAIL.n439 11.249
R581 VTAIL.n399 VTAIL.n340 11.249
R582 VTAIL.n370 VTAIL.n357 11.249
R583 VTAIL.n315 VTAIL.n256 11.249
R584 VTAIL.n286 VTAIL.n273 11.249
R585 VTAIL.n618 VTAIL.n602 10.4732
R586 VTAIL.n645 VTAIL.n590 10.4732
R587 VTAIL.n38 VTAIL.n22 10.4732
R588 VTAIL.n65 VTAIL.n10 10.4732
R589 VTAIL.n120 VTAIL.n104 10.4732
R590 VTAIL.n147 VTAIL.n92 10.4732
R591 VTAIL.n204 VTAIL.n188 10.4732
R592 VTAIL.n231 VTAIL.n176 10.4732
R593 VTAIL.n564 VTAIL.n509 10.4732
R594 VTAIL.n537 VTAIL.n521 10.4732
R595 VTAIL.n480 VTAIL.n425 10.4732
R596 VTAIL.n453 VTAIL.n437 10.4732
R597 VTAIL.n398 VTAIL.n343 10.4732
R598 VTAIL.n371 VTAIL.n355 10.4732
R599 VTAIL.n314 VTAIL.n259 10.4732
R600 VTAIL.n287 VTAIL.n271 10.4732
R601 VTAIL.n622 VTAIL.n621 9.69747
R602 VTAIL.n642 VTAIL.n641 9.69747
R603 VTAIL.n42 VTAIL.n41 9.69747
R604 VTAIL.n62 VTAIL.n61 9.69747
R605 VTAIL.n124 VTAIL.n123 9.69747
R606 VTAIL.n144 VTAIL.n143 9.69747
R607 VTAIL.n208 VTAIL.n207 9.69747
R608 VTAIL.n228 VTAIL.n227 9.69747
R609 VTAIL.n561 VTAIL.n560 9.69747
R610 VTAIL.n541 VTAIL.n540 9.69747
R611 VTAIL.n477 VTAIL.n476 9.69747
R612 VTAIL.n457 VTAIL.n456 9.69747
R613 VTAIL.n395 VTAIL.n394 9.69747
R614 VTAIL.n375 VTAIL.n374 9.69747
R615 VTAIL.n311 VTAIL.n310 9.69747
R616 VTAIL.n291 VTAIL.n290 9.69747
R617 VTAIL.n662 VTAIL.n661 9.45567
R618 VTAIL.n82 VTAIL.n81 9.45567
R619 VTAIL.n164 VTAIL.n163 9.45567
R620 VTAIL.n248 VTAIL.n247 9.45567
R621 VTAIL.n580 VTAIL.n579 9.45567
R622 VTAIL.n496 VTAIL.n495 9.45567
R623 VTAIL.n414 VTAIL.n413 9.45567
R624 VTAIL.n330 VTAIL.n329 9.45567
R625 VTAIL.n661 VTAIL.n660 9.3005
R626 VTAIL.n584 VTAIL.n583 9.3005
R627 VTAIL.n629 VTAIL.n628 9.3005
R628 VTAIL.n627 VTAIL.n626 9.3005
R629 VTAIL.n600 VTAIL.n599 9.3005
R630 VTAIL.n621 VTAIL.n620 9.3005
R631 VTAIL.n619 VTAIL.n618 9.3005
R632 VTAIL.n604 VTAIL.n603 9.3005
R633 VTAIL.n613 VTAIL.n612 9.3005
R634 VTAIL.n611 VTAIL.n610 9.3005
R635 VTAIL.n596 VTAIL.n595 9.3005
R636 VTAIL.n635 VTAIL.n634 9.3005
R637 VTAIL.n637 VTAIL.n636 9.3005
R638 VTAIL.n592 VTAIL.n591 9.3005
R639 VTAIL.n643 VTAIL.n642 9.3005
R640 VTAIL.n645 VTAIL.n644 9.3005
R641 VTAIL.n588 VTAIL.n587 9.3005
R642 VTAIL.n652 VTAIL.n651 9.3005
R643 VTAIL.n654 VTAIL.n653 9.3005
R644 VTAIL.n81 VTAIL.n80 9.3005
R645 VTAIL.n4 VTAIL.n3 9.3005
R646 VTAIL.n49 VTAIL.n48 9.3005
R647 VTAIL.n47 VTAIL.n46 9.3005
R648 VTAIL.n20 VTAIL.n19 9.3005
R649 VTAIL.n41 VTAIL.n40 9.3005
R650 VTAIL.n39 VTAIL.n38 9.3005
R651 VTAIL.n24 VTAIL.n23 9.3005
R652 VTAIL.n33 VTAIL.n32 9.3005
R653 VTAIL.n31 VTAIL.n30 9.3005
R654 VTAIL.n16 VTAIL.n15 9.3005
R655 VTAIL.n55 VTAIL.n54 9.3005
R656 VTAIL.n57 VTAIL.n56 9.3005
R657 VTAIL.n12 VTAIL.n11 9.3005
R658 VTAIL.n63 VTAIL.n62 9.3005
R659 VTAIL.n65 VTAIL.n64 9.3005
R660 VTAIL.n8 VTAIL.n7 9.3005
R661 VTAIL.n72 VTAIL.n71 9.3005
R662 VTAIL.n74 VTAIL.n73 9.3005
R663 VTAIL.n163 VTAIL.n162 9.3005
R664 VTAIL.n86 VTAIL.n85 9.3005
R665 VTAIL.n131 VTAIL.n130 9.3005
R666 VTAIL.n129 VTAIL.n128 9.3005
R667 VTAIL.n102 VTAIL.n101 9.3005
R668 VTAIL.n123 VTAIL.n122 9.3005
R669 VTAIL.n121 VTAIL.n120 9.3005
R670 VTAIL.n106 VTAIL.n105 9.3005
R671 VTAIL.n115 VTAIL.n114 9.3005
R672 VTAIL.n113 VTAIL.n112 9.3005
R673 VTAIL.n98 VTAIL.n97 9.3005
R674 VTAIL.n137 VTAIL.n136 9.3005
R675 VTAIL.n139 VTAIL.n138 9.3005
R676 VTAIL.n94 VTAIL.n93 9.3005
R677 VTAIL.n145 VTAIL.n144 9.3005
R678 VTAIL.n147 VTAIL.n146 9.3005
R679 VTAIL.n90 VTAIL.n89 9.3005
R680 VTAIL.n154 VTAIL.n153 9.3005
R681 VTAIL.n156 VTAIL.n155 9.3005
R682 VTAIL.n247 VTAIL.n246 9.3005
R683 VTAIL.n170 VTAIL.n169 9.3005
R684 VTAIL.n215 VTAIL.n214 9.3005
R685 VTAIL.n213 VTAIL.n212 9.3005
R686 VTAIL.n186 VTAIL.n185 9.3005
R687 VTAIL.n207 VTAIL.n206 9.3005
R688 VTAIL.n205 VTAIL.n204 9.3005
R689 VTAIL.n190 VTAIL.n189 9.3005
R690 VTAIL.n199 VTAIL.n198 9.3005
R691 VTAIL.n197 VTAIL.n196 9.3005
R692 VTAIL.n182 VTAIL.n181 9.3005
R693 VTAIL.n221 VTAIL.n220 9.3005
R694 VTAIL.n223 VTAIL.n222 9.3005
R695 VTAIL.n178 VTAIL.n177 9.3005
R696 VTAIL.n229 VTAIL.n228 9.3005
R697 VTAIL.n231 VTAIL.n230 9.3005
R698 VTAIL.n174 VTAIL.n173 9.3005
R699 VTAIL.n238 VTAIL.n237 9.3005
R700 VTAIL.n240 VTAIL.n239 9.3005
R701 VTAIL.n554 VTAIL.n553 9.3005
R702 VTAIL.n556 VTAIL.n555 9.3005
R703 VTAIL.n511 VTAIL.n510 9.3005
R704 VTAIL.n562 VTAIL.n561 9.3005
R705 VTAIL.n564 VTAIL.n563 9.3005
R706 VTAIL.n506 VTAIL.n505 9.3005
R707 VTAIL.n570 VTAIL.n569 9.3005
R708 VTAIL.n572 VTAIL.n571 9.3005
R709 VTAIL.n579 VTAIL.n578 9.3005
R710 VTAIL.n502 VTAIL.n501 9.3005
R711 VTAIL.n515 VTAIL.n514 9.3005
R712 VTAIL.n548 VTAIL.n547 9.3005
R713 VTAIL.n546 VTAIL.n545 9.3005
R714 VTAIL.n519 VTAIL.n518 9.3005
R715 VTAIL.n540 VTAIL.n539 9.3005
R716 VTAIL.n538 VTAIL.n537 9.3005
R717 VTAIL.n523 VTAIL.n522 9.3005
R718 VTAIL.n532 VTAIL.n531 9.3005
R719 VTAIL.n530 VTAIL.n529 9.3005
R720 VTAIL.n470 VTAIL.n469 9.3005
R721 VTAIL.n472 VTAIL.n471 9.3005
R722 VTAIL.n427 VTAIL.n426 9.3005
R723 VTAIL.n478 VTAIL.n477 9.3005
R724 VTAIL.n480 VTAIL.n479 9.3005
R725 VTAIL.n422 VTAIL.n421 9.3005
R726 VTAIL.n486 VTAIL.n485 9.3005
R727 VTAIL.n488 VTAIL.n487 9.3005
R728 VTAIL.n495 VTAIL.n494 9.3005
R729 VTAIL.n418 VTAIL.n417 9.3005
R730 VTAIL.n431 VTAIL.n430 9.3005
R731 VTAIL.n464 VTAIL.n463 9.3005
R732 VTAIL.n462 VTAIL.n461 9.3005
R733 VTAIL.n435 VTAIL.n434 9.3005
R734 VTAIL.n456 VTAIL.n455 9.3005
R735 VTAIL.n454 VTAIL.n453 9.3005
R736 VTAIL.n439 VTAIL.n438 9.3005
R737 VTAIL.n448 VTAIL.n447 9.3005
R738 VTAIL.n446 VTAIL.n445 9.3005
R739 VTAIL.n388 VTAIL.n387 9.3005
R740 VTAIL.n390 VTAIL.n389 9.3005
R741 VTAIL.n345 VTAIL.n344 9.3005
R742 VTAIL.n396 VTAIL.n395 9.3005
R743 VTAIL.n398 VTAIL.n397 9.3005
R744 VTAIL.n340 VTAIL.n339 9.3005
R745 VTAIL.n404 VTAIL.n403 9.3005
R746 VTAIL.n406 VTAIL.n405 9.3005
R747 VTAIL.n413 VTAIL.n412 9.3005
R748 VTAIL.n336 VTAIL.n335 9.3005
R749 VTAIL.n349 VTAIL.n348 9.3005
R750 VTAIL.n382 VTAIL.n381 9.3005
R751 VTAIL.n380 VTAIL.n379 9.3005
R752 VTAIL.n353 VTAIL.n352 9.3005
R753 VTAIL.n374 VTAIL.n373 9.3005
R754 VTAIL.n372 VTAIL.n371 9.3005
R755 VTAIL.n357 VTAIL.n356 9.3005
R756 VTAIL.n366 VTAIL.n365 9.3005
R757 VTAIL.n364 VTAIL.n363 9.3005
R758 VTAIL.n304 VTAIL.n303 9.3005
R759 VTAIL.n306 VTAIL.n305 9.3005
R760 VTAIL.n261 VTAIL.n260 9.3005
R761 VTAIL.n312 VTAIL.n311 9.3005
R762 VTAIL.n314 VTAIL.n313 9.3005
R763 VTAIL.n256 VTAIL.n255 9.3005
R764 VTAIL.n320 VTAIL.n319 9.3005
R765 VTAIL.n322 VTAIL.n321 9.3005
R766 VTAIL.n329 VTAIL.n328 9.3005
R767 VTAIL.n252 VTAIL.n251 9.3005
R768 VTAIL.n265 VTAIL.n264 9.3005
R769 VTAIL.n298 VTAIL.n297 9.3005
R770 VTAIL.n296 VTAIL.n295 9.3005
R771 VTAIL.n269 VTAIL.n268 9.3005
R772 VTAIL.n290 VTAIL.n289 9.3005
R773 VTAIL.n288 VTAIL.n287 9.3005
R774 VTAIL.n273 VTAIL.n272 9.3005
R775 VTAIL.n282 VTAIL.n281 9.3005
R776 VTAIL.n280 VTAIL.n279 9.3005
R777 VTAIL.n625 VTAIL.n600 8.92171
R778 VTAIL.n638 VTAIL.n592 8.92171
R779 VTAIL.n45 VTAIL.n20 8.92171
R780 VTAIL.n58 VTAIL.n12 8.92171
R781 VTAIL.n127 VTAIL.n102 8.92171
R782 VTAIL.n140 VTAIL.n94 8.92171
R783 VTAIL.n211 VTAIL.n186 8.92171
R784 VTAIL.n224 VTAIL.n178 8.92171
R785 VTAIL.n557 VTAIL.n511 8.92171
R786 VTAIL.n544 VTAIL.n519 8.92171
R787 VTAIL.n473 VTAIL.n427 8.92171
R788 VTAIL.n460 VTAIL.n435 8.92171
R789 VTAIL.n391 VTAIL.n345 8.92171
R790 VTAIL.n378 VTAIL.n353 8.92171
R791 VTAIL.n307 VTAIL.n261 8.92171
R792 VTAIL.n294 VTAIL.n269 8.92171
R793 VTAIL.n626 VTAIL.n598 8.14595
R794 VTAIL.n637 VTAIL.n594 8.14595
R795 VTAIL.n46 VTAIL.n18 8.14595
R796 VTAIL.n57 VTAIL.n14 8.14595
R797 VTAIL.n128 VTAIL.n100 8.14595
R798 VTAIL.n139 VTAIL.n96 8.14595
R799 VTAIL.n212 VTAIL.n184 8.14595
R800 VTAIL.n223 VTAIL.n180 8.14595
R801 VTAIL.n556 VTAIL.n513 8.14595
R802 VTAIL.n545 VTAIL.n517 8.14595
R803 VTAIL.n472 VTAIL.n429 8.14595
R804 VTAIL.n461 VTAIL.n433 8.14595
R805 VTAIL.n390 VTAIL.n347 8.14595
R806 VTAIL.n379 VTAIL.n351 8.14595
R807 VTAIL.n306 VTAIL.n263 8.14595
R808 VTAIL.n295 VTAIL.n267 8.14595
R809 VTAIL.n630 VTAIL.n629 7.3702
R810 VTAIL.n634 VTAIL.n633 7.3702
R811 VTAIL.n50 VTAIL.n49 7.3702
R812 VTAIL.n54 VTAIL.n53 7.3702
R813 VTAIL.n132 VTAIL.n131 7.3702
R814 VTAIL.n136 VTAIL.n135 7.3702
R815 VTAIL.n216 VTAIL.n215 7.3702
R816 VTAIL.n220 VTAIL.n219 7.3702
R817 VTAIL.n553 VTAIL.n552 7.3702
R818 VTAIL.n549 VTAIL.n548 7.3702
R819 VTAIL.n469 VTAIL.n468 7.3702
R820 VTAIL.n465 VTAIL.n464 7.3702
R821 VTAIL.n387 VTAIL.n386 7.3702
R822 VTAIL.n383 VTAIL.n382 7.3702
R823 VTAIL.n303 VTAIL.n302 7.3702
R824 VTAIL.n299 VTAIL.n298 7.3702
R825 VTAIL.n630 VTAIL.n596 6.59444
R826 VTAIL.n633 VTAIL.n596 6.59444
R827 VTAIL.n50 VTAIL.n16 6.59444
R828 VTAIL.n53 VTAIL.n16 6.59444
R829 VTAIL.n132 VTAIL.n98 6.59444
R830 VTAIL.n135 VTAIL.n98 6.59444
R831 VTAIL.n216 VTAIL.n182 6.59444
R832 VTAIL.n219 VTAIL.n182 6.59444
R833 VTAIL.n552 VTAIL.n515 6.59444
R834 VTAIL.n549 VTAIL.n515 6.59444
R835 VTAIL.n468 VTAIL.n431 6.59444
R836 VTAIL.n465 VTAIL.n431 6.59444
R837 VTAIL.n386 VTAIL.n349 6.59444
R838 VTAIL.n383 VTAIL.n349 6.59444
R839 VTAIL.n302 VTAIL.n265 6.59444
R840 VTAIL.n299 VTAIL.n265 6.59444
R841 VTAIL.n629 VTAIL.n598 5.81868
R842 VTAIL.n634 VTAIL.n594 5.81868
R843 VTAIL.n49 VTAIL.n18 5.81868
R844 VTAIL.n54 VTAIL.n14 5.81868
R845 VTAIL.n131 VTAIL.n100 5.81868
R846 VTAIL.n136 VTAIL.n96 5.81868
R847 VTAIL.n215 VTAIL.n184 5.81868
R848 VTAIL.n220 VTAIL.n180 5.81868
R849 VTAIL.n553 VTAIL.n513 5.81868
R850 VTAIL.n548 VTAIL.n517 5.81868
R851 VTAIL.n469 VTAIL.n429 5.81868
R852 VTAIL.n464 VTAIL.n433 5.81868
R853 VTAIL.n387 VTAIL.n347 5.81868
R854 VTAIL.n382 VTAIL.n351 5.81868
R855 VTAIL.n303 VTAIL.n263 5.81868
R856 VTAIL.n298 VTAIL.n267 5.81868
R857 VTAIL.n626 VTAIL.n625 5.04292
R858 VTAIL.n638 VTAIL.n637 5.04292
R859 VTAIL.n46 VTAIL.n45 5.04292
R860 VTAIL.n58 VTAIL.n57 5.04292
R861 VTAIL.n128 VTAIL.n127 5.04292
R862 VTAIL.n140 VTAIL.n139 5.04292
R863 VTAIL.n212 VTAIL.n211 5.04292
R864 VTAIL.n224 VTAIL.n223 5.04292
R865 VTAIL.n557 VTAIL.n556 5.04292
R866 VTAIL.n545 VTAIL.n544 5.04292
R867 VTAIL.n473 VTAIL.n472 5.04292
R868 VTAIL.n461 VTAIL.n460 5.04292
R869 VTAIL.n391 VTAIL.n390 5.04292
R870 VTAIL.n379 VTAIL.n378 5.04292
R871 VTAIL.n307 VTAIL.n306 5.04292
R872 VTAIL.n295 VTAIL.n294 5.04292
R873 VTAIL.n622 VTAIL.n600 4.26717
R874 VTAIL.n641 VTAIL.n592 4.26717
R875 VTAIL.n42 VTAIL.n20 4.26717
R876 VTAIL.n61 VTAIL.n12 4.26717
R877 VTAIL.n124 VTAIL.n102 4.26717
R878 VTAIL.n143 VTAIL.n94 4.26717
R879 VTAIL.n208 VTAIL.n186 4.26717
R880 VTAIL.n227 VTAIL.n178 4.26717
R881 VTAIL.n560 VTAIL.n511 4.26717
R882 VTAIL.n541 VTAIL.n519 4.26717
R883 VTAIL.n476 VTAIL.n427 4.26717
R884 VTAIL.n457 VTAIL.n435 4.26717
R885 VTAIL.n394 VTAIL.n345 4.26717
R886 VTAIL.n375 VTAIL.n353 4.26717
R887 VTAIL.n310 VTAIL.n261 4.26717
R888 VTAIL.n291 VTAIL.n269 4.26717
R889 VTAIL.n611 VTAIL.n607 3.70982
R890 VTAIL.n31 VTAIL.n27 3.70982
R891 VTAIL.n113 VTAIL.n109 3.70982
R892 VTAIL.n197 VTAIL.n193 3.70982
R893 VTAIL.n530 VTAIL.n526 3.70982
R894 VTAIL.n446 VTAIL.n442 3.70982
R895 VTAIL.n364 VTAIL.n360 3.70982
R896 VTAIL.n280 VTAIL.n276 3.70982
R897 VTAIL.n621 VTAIL.n602 3.49141
R898 VTAIL.n642 VTAIL.n590 3.49141
R899 VTAIL.n41 VTAIL.n22 3.49141
R900 VTAIL.n62 VTAIL.n10 3.49141
R901 VTAIL.n123 VTAIL.n104 3.49141
R902 VTAIL.n144 VTAIL.n92 3.49141
R903 VTAIL.n207 VTAIL.n188 3.49141
R904 VTAIL.n228 VTAIL.n176 3.49141
R905 VTAIL.n561 VTAIL.n509 3.49141
R906 VTAIL.n540 VTAIL.n521 3.49141
R907 VTAIL.n477 VTAIL.n425 3.49141
R908 VTAIL.n456 VTAIL.n437 3.49141
R909 VTAIL.n395 VTAIL.n343 3.49141
R910 VTAIL.n374 VTAIL.n355 3.49141
R911 VTAIL.n311 VTAIL.n259 3.49141
R912 VTAIL.n290 VTAIL.n271 3.49141
R913 VTAIL.n333 VTAIL.n331 3.37119
R914 VTAIL.n415 VTAIL.n333 3.37119
R915 VTAIL.n499 VTAIL.n497 3.37119
R916 VTAIL.n581 VTAIL.n499 3.37119
R917 VTAIL.n249 VTAIL.n167 3.37119
R918 VTAIL.n167 VTAIL.n165 3.37119
R919 VTAIL.n83 VTAIL.n1 3.37119
R920 VTAIL VTAIL.n663 3.313
R921 VTAIL.n618 VTAIL.n617 2.71565
R922 VTAIL.n646 VTAIL.n645 2.71565
R923 VTAIL.n38 VTAIL.n37 2.71565
R924 VTAIL.n66 VTAIL.n65 2.71565
R925 VTAIL.n120 VTAIL.n119 2.71565
R926 VTAIL.n148 VTAIL.n147 2.71565
R927 VTAIL.n204 VTAIL.n203 2.71565
R928 VTAIL.n232 VTAIL.n231 2.71565
R929 VTAIL.n565 VTAIL.n564 2.71565
R930 VTAIL.n537 VTAIL.n536 2.71565
R931 VTAIL.n481 VTAIL.n480 2.71565
R932 VTAIL.n453 VTAIL.n452 2.71565
R933 VTAIL.n399 VTAIL.n398 2.71565
R934 VTAIL.n371 VTAIL.n370 2.71565
R935 VTAIL.n315 VTAIL.n314 2.71565
R936 VTAIL.n287 VTAIL.n286 2.71565
R937 VTAIL.n0 VTAIL.t6 2.20274
R938 VTAIL.n0 VTAIL.t2 2.20274
R939 VTAIL.n166 VTAIL.t13 2.20274
R940 VTAIL.n166 VTAIL.t12 2.20274
R941 VTAIL.n498 VTAIL.t11 2.20274
R942 VTAIL.n498 VTAIL.t10 2.20274
R943 VTAIL.n332 VTAIL.t3 2.20274
R944 VTAIL.n332 VTAIL.t0 2.20274
R945 VTAIL.n614 VTAIL.n604 1.93989
R946 VTAIL.n650 VTAIL.n588 1.93989
R947 VTAIL.n662 VTAIL.n582 1.93989
R948 VTAIL.n34 VTAIL.n24 1.93989
R949 VTAIL.n70 VTAIL.n8 1.93989
R950 VTAIL.n82 VTAIL.n2 1.93989
R951 VTAIL.n116 VTAIL.n106 1.93989
R952 VTAIL.n152 VTAIL.n90 1.93989
R953 VTAIL.n164 VTAIL.n84 1.93989
R954 VTAIL.n200 VTAIL.n190 1.93989
R955 VTAIL.n236 VTAIL.n174 1.93989
R956 VTAIL.n248 VTAIL.n168 1.93989
R957 VTAIL.n580 VTAIL.n500 1.93989
R958 VTAIL.n568 VTAIL.n506 1.93989
R959 VTAIL.n533 VTAIL.n523 1.93989
R960 VTAIL.n496 VTAIL.n416 1.93989
R961 VTAIL.n484 VTAIL.n422 1.93989
R962 VTAIL.n449 VTAIL.n439 1.93989
R963 VTAIL.n414 VTAIL.n334 1.93989
R964 VTAIL.n402 VTAIL.n340 1.93989
R965 VTAIL.n367 VTAIL.n357 1.93989
R966 VTAIL.n330 VTAIL.n250 1.93989
R967 VTAIL.n318 VTAIL.n256 1.93989
R968 VTAIL.n283 VTAIL.n273 1.93989
R969 VTAIL.n613 VTAIL.n606 1.16414
R970 VTAIL.n651 VTAIL.n586 1.16414
R971 VTAIL.n660 VTAIL.n659 1.16414
R972 VTAIL.n33 VTAIL.n26 1.16414
R973 VTAIL.n71 VTAIL.n6 1.16414
R974 VTAIL.n80 VTAIL.n79 1.16414
R975 VTAIL.n115 VTAIL.n108 1.16414
R976 VTAIL.n153 VTAIL.n88 1.16414
R977 VTAIL.n162 VTAIL.n161 1.16414
R978 VTAIL.n199 VTAIL.n192 1.16414
R979 VTAIL.n237 VTAIL.n172 1.16414
R980 VTAIL.n246 VTAIL.n245 1.16414
R981 VTAIL.n578 VTAIL.n577 1.16414
R982 VTAIL.n569 VTAIL.n504 1.16414
R983 VTAIL.n532 VTAIL.n525 1.16414
R984 VTAIL.n494 VTAIL.n493 1.16414
R985 VTAIL.n485 VTAIL.n420 1.16414
R986 VTAIL.n448 VTAIL.n441 1.16414
R987 VTAIL.n412 VTAIL.n411 1.16414
R988 VTAIL.n403 VTAIL.n338 1.16414
R989 VTAIL.n366 VTAIL.n359 1.16414
R990 VTAIL.n328 VTAIL.n327 1.16414
R991 VTAIL.n319 VTAIL.n254 1.16414
R992 VTAIL.n282 VTAIL.n275 1.16414
R993 VTAIL.n497 VTAIL.n415 0.470328
R994 VTAIL.n165 VTAIL.n83 0.470328
R995 VTAIL.n610 VTAIL.n609 0.388379
R996 VTAIL.n655 VTAIL.n654 0.388379
R997 VTAIL.n656 VTAIL.n584 0.388379
R998 VTAIL.n30 VTAIL.n29 0.388379
R999 VTAIL.n75 VTAIL.n74 0.388379
R1000 VTAIL.n76 VTAIL.n4 0.388379
R1001 VTAIL.n112 VTAIL.n111 0.388379
R1002 VTAIL.n157 VTAIL.n156 0.388379
R1003 VTAIL.n158 VTAIL.n86 0.388379
R1004 VTAIL.n196 VTAIL.n195 0.388379
R1005 VTAIL.n241 VTAIL.n240 0.388379
R1006 VTAIL.n242 VTAIL.n170 0.388379
R1007 VTAIL.n574 VTAIL.n502 0.388379
R1008 VTAIL.n573 VTAIL.n572 0.388379
R1009 VTAIL.n529 VTAIL.n528 0.388379
R1010 VTAIL.n490 VTAIL.n418 0.388379
R1011 VTAIL.n489 VTAIL.n488 0.388379
R1012 VTAIL.n445 VTAIL.n444 0.388379
R1013 VTAIL.n408 VTAIL.n336 0.388379
R1014 VTAIL.n407 VTAIL.n406 0.388379
R1015 VTAIL.n363 VTAIL.n362 0.388379
R1016 VTAIL.n324 VTAIL.n252 0.388379
R1017 VTAIL.n323 VTAIL.n322 0.388379
R1018 VTAIL.n279 VTAIL.n278 0.388379
R1019 VTAIL.n612 VTAIL.n611 0.155672
R1020 VTAIL.n612 VTAIL.n603 0.155672
R1021 VTAIL.n619 VTAIL.n603 0.155672
R1022 VTAIL.n620 VTAIL.n619 0.155672
R1023 VTAIL.n620 VTAIL.n599 0.155672
R1024 VTAIL.n627 VTAIL.n599 0.155672
R1025 VTAIL.n628 VTAIL.n627 0.155672
R1026 VTAIL.n628 VTAIL.n595 0.155672
R1027 VTAIL.n635 VTAIL.n595 0.155672
R1028 VTAIL.n636 VTAIL.n635 0.155672
R1029 VTAIL.n636 VTAIL.n591 0.155672
R1030 VTAIL.n643 VTAIL.n591 0.155672
R1031 VTAIL.n644 VTAIL.n643 0.155672
R1032 VTAIL.n644 VTAIL.n587 0.155672
R1033 VTAIL.n652 VTAIL.n587 0.155672
R1034 VTAIL.n653 VTAIL.n652 0.155672
R1035 VTAIL.n653 VTAIL.n583 0.155672
R1036 VTAIL.n661 VTAIL.n583 0.155672
R1037 VTAIL.n32 VTAIL.n31 0.155672
R1038 VTAIL.n32 VTAIL.n23 0.155672
R1039 VTAIL.n39 VTAIL.n23 0.155672
R1040 VTAIL.n40 VTAIL.n39 0.155672
R1041 VTAIL.n40 VTAIL.n19 0.155672
R1042 VTAIL.n47 VTAIL.n19 0.155672
R1043 VTAIL.n48 VTAIL.n47 0.155672
R1044 VTAIL.n48 VTAIL.n15 0.155672
R1045 VTAIL.n55 VTAIL.n15 0.155672
R1046 VTAIL.n56 VTAIL.n55 0.155672
R1047 VTAIL.n56 VTAIL.n11 0.155672
R1048 VTAIL.n63 VTAIL.n11 0.155672
R1049 VTAIL.n64 VTAIL.n63 0.155672
R1050 VTAIL.n64 VTAIL.n7 0.155672
R1051 VTAIL.n72 VTAIL.n7 0.155672
R1052 VTAIL.n73 VTAIL.n72 0.155672
R1053 VTAIL.n73 VTAIL.n3 0.155672
R1054 VTAIL.n81 VTAIL.n3 0.155672
R1055 VTAIL.n114 VTAIL.n113 0.155672
R1056 VTAIL.n114 VTAIL.n105 0.155672
R1057 VTAIL.n121 VTAIL.n105 0.155672
R1058 VTAIL.n122 VTAIL.n121 0.155672
R1059 VTAIL.n122 VTAIL.n101 0.155672
R1060 VTAIL.n129 VTAIL.n101 0.155672
R1061 VTAIL.n130 VTAIL.n129 0.155672
R1062 VTAIL.n130 VTAIL.n97 0.155672
R1063 VTAIL.n137 VTAIL.n97 0.155672
R1064 VTAIL.n138 VTAIL.n137 0.155672
R1065 VTAIL.n138 VTAIL.n93 0.155672
R1066 VTAIL.n145 VTAIL.n93 0.155672
R1067 VTAIL.n146 VTAIL.n145 0.155672
R1068 VTAIL.n146 VTAIL.n89 0.155672
R1069 VTAIL.n154 VTAIL.n89 0.155672
R1070 VTAIL.n155 VTAIL.n154 0.155672
R1071 VTAIL.n155 VTAIL.n85 0.155672
R1072 VTAIL.n163 VTAIL.n85 0.155672
R1073 VTAIL.n198 VTAIL.n197 0.155672
R1074 VTAIL.n198 VTAIL.n189 0.155672
R1075 VTAIL.n205 VTAIL.n189 0.155672
R1076 VTAIL.n206 VTAIL.n205 0.155672
R1077 VTAIL.n206 VTAIL.n185 0.155672
R1078 VTAIL.n213 VTAIL.n185 0.155672
R1079 VTAIL.n214 VTAIL.n213 0.155672
R1080 VTAIL.n214 VTAIL.n181 0.155672
R1081 VTAIL.n221 VTAIL.n181 0.155672
R1082 VTAIL.n222 VTAIL.n221 0.155672
R1083 VTAIL.n222 VTAIL.n177 0.155672
R1084 VTAIL.n229 VTAIL.n177 0.155672
R1085 VTAIL.n230 VTAIL.n229 0.155672
R1086 VTAIL.n230 VTAIL.n173 0.155672
R1087 VTAIL.n238 VTAIL.n173 0.155672
R1088 VTAIL.n239 VTAIL.n238 0.155672
R1089 VTAIL.n239 VTAIL.n169 0.155672
R1090 VTAIL.n247 VTAIL.n169 0.155672
R1091 VTAIL.n579 VTAIL.n501 0.155672
R1092 VTAIL.n571 VTAIL.n501 0.155672
R1093 VTAIL.n571 VTAIL.n570 0.155672
R1094 VTAIL.n570 VTAIL.n505 0.155672
R1095 VTAIL.n563 VTAIL.n505 0.155672
R1096 VTAIL.n563 VTAIL.n562 0.155672
R1097 VTAIL.n562 VTAIL.n510 0.155672
R1098 VTAIL.n555 VTAIL.n510 0.155672
R1099 VTAIL.n555 VTAIL.n554 0.155672
R1100 VTAIL.n554 VTAIL.n514 0.155672
R1101 VTAIL.n547 VTAIL.n514 0.155672
R1102 VTAIL.n547 VTAIL.n546 0.155672
R1103 VTAIL.n546 VTAIL.n518 0.155672
R1104 VTAIL.n539 VTAIL.n518 0.155672
R1105 VTAIL.n539 VTAIL.n538 0.155672
R1106 VTAIL.n538 VTAIL.n522 0.155672
R1107 VTAIL.n531 VTAIL.n522 0.155672
R1108 VTAIL.n531 VTAIL.n530 0.155672
R1109 VTAIL.n495 VTAIL.n417 0.155672
R1110 VTAIL.n487 VTAIL.n417 0.155672
R1111 VTAIL.n487 VTAIL.n486 0.155672
R1112 VTAIL.n486 VTAIL.n421 0.155672
R1113 VTAIL.n479 VTAIL.n421 0.155672
R1114 VTAIL.n479 VTAIL.n478 0.155672
R1115 VTAIL.n478 VTAIL.n426 0.155672
R1116 VTAIL.n471 VTAIL.n426 0.155672
R1117 VTAIL.n471 VTAIL.n470 0.155672
R1118 VTAIL.n470 VTAIL.n430 0.155672
R1119 VTAIL.n463 VTAIL.n430 0.155672
R1120 VTAIL.n463 VTAIL.n462 0.155672
R1121 VTAIL.n462 VTAIL.n434 0.155672
R1122 VTAIL.n455 VTAIL.n434 0.155672
R1123 VTAIL.n455 VTAIL.n454 0.155672
R1124 VTAIL.n454 VTAIL.n438 0.155672
R1125 VTAIL.n447 VTAIL.n438 0.155672
R1126 VTAIL.n447 VTAIL.n446 0.155672
R1127 VTAIL.n413 VTAIL.n335 0.155672
R1128 VTAIL.n405 VTAIL.n335 0.155672
R1129 VTAIL.n405 VTAIL.n404 0.155672
R1130 VTAIL.n404 VTAIL.n339 0.155672
R1131 VTAIL.n397 VTAIL.n339 0.155672
R1132 VTAIL.n397 VTAIL.n396 0.155672
R1133 VTAIL.n396 VTAIL.n344 0.155672
R1134 VTAIL.n389 VTAIL.n344 0.155672
R1135 VTAIL.n389 VTAIL.n388 0.155672
R1136 VTAIL.n388 VTAIL.n348 0.155672
R1137 VTAIL.n381 VTAIL.n348 0.155672
R1138 VTAIL.n381 VTAIL.n380 0.155672
R1139 VTAIL.n380 VTAIL.n352 0.155672
R1140 VTAIL.n373 VTAIL.n352 0.155672
R1141 VTAIL.n373 VTAIL.n372 0.155672
R1142 VTAIL.n372 VTAIL.n356 0.155672
R1143 VTAIL.n365 VTAIL.n356 0.155672
R1144 VTAIL.n365 VTAIL.n364 0.155672
R1145 VTAIL.n329 VTAIL.n251 0.155672
R1146 VTAIL.n321 VTAIL.n251 0.155672
R1147 VTAIL.n321 VTAIL.n320 0.155672
R1148 VTAIL.n320 VTAIL.n255 0.155672
R1149 VTAIL.n313 VTAIL.n255 0.155672
R1150 VTAIL.n313 VTAIL.n312 0.155672
R1151 VTAIL.n312 VTAIL.n260 0.155672
R1152 VTAIL.n305 VTAIL.n260 0.155672
R1153 VTAIL.n305 VTAIL.n304 0.155672
R1154 VTAIL.n304 VTAIL.n264 0.155672
R1155 VTAIL.n297 VTAIL.n264 0.155672
R1156 VTAIL.n297 VTAIL.n296 0.155672
R1157 VTAIL.n296 VTAIL.n268 0.155672
R1158 VTAIL.n289 VTAIL.n268 0.155672
R1159 VTAIL.n289 VTAIL.n288 0.155672
R1160 VTAIL.n288 VTAIL.n272 0.155672
R1161 VTAIL.n281 VTAIL.n272 0.155672
R1162 VTAIL.n281 VTAIL.n280 0.155672
R1163 VTAIL VTAIL.n1 0.0586897
R1164 B.n511 B.n510 585
R1165 B.n509 B.n160 585
R1166 B.n508 B.n507 585
R1167 B.n506 B.n161 585
R1168 B.n505 B.n504 585
R1169 B.n503 B.n162 585
R1170 B.n502 B.n501 585
R1171 B.n500 B.n163 585
R1172 B.n499 B.n498 585
R1173 B.n497 B.n164 585
R1174 B.n496 B.n495 585
R1175 B.n494 B.n165 585
R1176 B.n493 B.n492 585
R1177 B.n491 B.n166 585
R1178 B.n490 B.n489 585
R1179 B.n488 B.n167 585
R1180 B.n487 B.n486 585
R1181 B.n485 B.n168 585
R1182 B.n484 B.n483 585
R1183 B.n482 B.n169 585
R1184 B.n481 B.n480 585
R1185 B.n479 B.n170 585
R1186 B.n478 B.n477 585
R1187 B.n476 B.n171 585
R1188 B.n475 B.n474 585
R1189 B.n473 B.n172 585
R1190 B.n472 B.n471 585
R1191 B.n470 B.n173 585
R1192 B.n469 B.n468 585
R1193 B.n467 B.n174 585
R1194 B.n466 B.n465 585
R1195 B.n464 B.n175 585
R1196 B.n463 B.n462 585
R1197 B.n461 B.n176 585
R1198 B.n460 B.n459 585
R1199 B.n458 B.n177 585
R1200 B.n457 B.n456 585
R1201 B.n455 B.n178 585
R1202 B.n454 B.n453 585
R1203 B.n452 B.n179 585
R1204 B.n451 B.n450 585
R1205 B.n449 B.n180 585
R1206 B.n448 B.n447 585
R1207 B.n446 B.n181 585
R1208 B.n445 B.n444 585
R1209 B.n443 B.n182 585
R1210 B.n442 B.n441 585
R1211 B.n440 B.n183 585
R1212 B.n439 B.n438 585
R1213 B.n437 B.n184 585
R1214 B.n436 B.n435 585
R1215 B.n431 B.n185 585
R1216 B.n430 B.n429 585
R1217 B.n428 B.n186 585
R1218 B.n427 B.n426 585
R1219 B.n425 B.n187 585
R1220 B.n424 B.n423 585
R1221 B.n422 B.n188 585
R1222 B.n421 B.n420 585
R1223 B.n418 B.n189 585
R1224 B.n417 B.n416 585
R1225 B.n415 B.n192 585
R1226 B.n414 B.n413 585
R1227 B.n412 B.n193 585
R1228 B.n411 B.n410 585
R1229 B.n409 B.n194 585
R1230 B.n408 B.n407 585
R1231 B.n406 B.n195 585
R1232 B.n405 B.n404 585
R1233 B.n403 B.n196 585
R1234 B.n402 B.n401 585
R1235 B.n400 B.n197 585
R1236 B.n399 B.n398 585
R1237 B.n397 B.n198 585
R1238 B.n396 B.n395 585
R1239 B.n394 B.n199 585
R1240 B.n393 B.n392 585
R1241 B.n391 B.n200 585
R1242 B.n390 B.n389 585
R1243 B.n388 B.n201 585
R1244 B.n387 B.n386 585
R1245 B.n385 B.n202 585
R1246 B.n384 B.n383 585
R1247 B.n382 B.n203 585
R1248 B.n381 B.n380 585
R1249 B.n379 B.n204 585
R1250 B.n378 B.n377 585
R1251 B.n376 B.n205 585
R1252 B.n375 B.n374 585
R1253 B.n373 B.n206 585
R1254 B.n372 B.n371 585
R1255 B.n370 B.n207 585
R1256 B.n369 B.n368 585
R1257 B.n367 B.n208 585
R1258 B.n366 B.n365 585
R1259 B.n364 B.n209 585
R1260 B.n363 B.n362 585
R1261 B.n361 B.n210 585
R1262 B.n360 B.n359 585
R1263 B.n358 B.n211 585
R1264 B.n357 B.n356 585
R1265 B.n355 B.n212 585
R1266 B.n354 B.n353 585
R1267 B.n352 B.n213 585
R1268 B.n351 B.n350 585
R1269 B.n349 B.n214 585
R1270 B.n348 B.n347 585
R1271 B.n346 B.n215 585
R1272 B.n345 B.n344 585
R1273 B.n512 B.n159 585
R1274 B.n514 B.n513 585
R1275 B.n515 B.n158 585
R1276 B.n517 B.n516 585
R1277 B.n518 B.n157 585
R1278 B.n520 B.n519 585
R1279 B.n521 B.n156 585
R1280 B.n523 B.n522 585
R1281 B.n524 B.n155 585
R1282 B.n526 B.n525 585
R1283 B.n527 B.n154 585
R1284 B.n529 B.n528 585
R1285 B.n530 B.n153 585
R1286 B.n532 B.n531 585
R1287 B.n533 B.n152 585
R1288 B.n535 B.n534 585
R1289 B.n536 B.n151 585
R1290 B.n538 B.n537 585
R1291 B.n539 B.n150 585
R1292 B.n541 B.n540 585
R1293 B.n542 B.n149 585
R1294 B.n544 B.n543 585
R1295 B.n545 B.n148 585
R1296 B.n547 B.n546 585
R1297 B.n548 B.n147 585
R1298 B.n550 B.n549 585
R1299 B.n551 B.n146 585
R1300 B.n553 B.n552 585
R1301 B.n554 B.n145 585
R1302 B.n556 B.n555 585
R1303 B.n557 B.n144 585
R1304 B.n559 B.n558 585
R1305 B.n560 B.n143 585
R1306 B.n562 B.n561 585
R1307 B.n563 B.n142 585
R1308 B.n565 B.n564 585
R1309 B.n566 B.n141 585
R1310 B.n568 B.n567 585
R1311 B.n569 B.n140 585
R1312 B.n571 B.n570 585
R1313 B.n572 B.n139 585
R1314 B.n574 B.n573 585
R1315 B.n575 B.n138 585
R1316 B.n577 B.n576 585
R1317 B.n578 B.n137 585
R1318 B.n580 B.n579 585
R1319 B.n581 B.n136 585
R1320 B.n583 B.n582 585
R1321 B.n584 B.n135 585
R1322 B.n586 B.n585 585
R1323 B.n587 B.n134 585
R1324 B.n589 B.n588 585
R1325 B.n590 B.n133 585
R1326 B.n592 B.n591 585
R1327 B.n593 B.n132 585
R1328 B.n595 B.n594 585
R1329 B.n596 B.n131 585
R1330 B.n598 B.n597 585
R1331 B.n599 B.n130 585
R1332 B.n601 B.n600 585
R1333 B.n602 B.n129 585
R1334 B.n604 B.n603 585
R1335 B.n605 B.n128 585
R1336 B.n607 B.n606 585
R1337 B.n608 B.n127 585
R1338 B.n610 B.n609 585
R1339 B.n611 B.n126 585
R1340 B.n613 B.n612 585
R1341 B.n614 B.n125 585
R1342 B.n616 B.n615 585
R1343 B.n617 B.n124 585
R1344 B.n619 B.n618 585
R1345 B.n620 B.n123 585
R1346 B.n622 B.n621 585
R1347 B.n623 B.n122 585
R1348 B.n625 B.n624 585
R1349 B.n626 B.n121 585
R1350 B.n628 B.n627 585
R1351 B.n629 B.n120 585
R1352 B.n631 B.n630 585
R1353 B.n632 B.n119 585
R1354 B.n634 B.n633 585
R1355 B.n635 B.n118 585
R1356 B.n637 B.n636 585
R1357 B.n638 B.n117 585
R1358 B.n640 B.n639 585
R1359 B.n641 B.n116 585
R1360 B.n643 B.n642 585
R1361 B.n644 B.n115 585
R1362 B.n646 B.n645 585
R1363 B.n647 B.n114 585
R1364 B.n649 B.n648 585
R1365 B.n650 B.n113 585
R1366 B.n652 B.n651 585
R1367 B.n653 B.n112 585
R1368 B.n655 B.n654 585
R1369 B.n656 B.n111 585
R1370 B.n658 B.n657 585
R1371 B.n659 B.n110 585
R1372 B.n661 B.n660 585
R1373 B.n662 B.n109 585
R1374 B.n664 B.n663 585
R1375 B.n665 B.n108 585
R1376 B.n667 B.n666 585
R1377 B.n668 B.n107 585
R1378 B.n670 B.n669 585
R1379 B.n671 B.n106 585
R1380 B.n673 B.n672 585
R1381 B.n674 B.n105 585
R1382 B.n676 B.n675 585
R1383 B.n677 B.n104 585
R1384 B.n679 B.n678 585
R1385 B.n680 B.n103 585
R1386 B.n682 B.n681 585
R1387 B.n683 B.n102 585
R1388 B.n685 B.n684 585
R1389 B.n686 B.n101 585
R1390 B.n688 B.n687 585
R1391 B.n689 B.n100 585
R1392 B.n691 B.n690 585
R1393 B.n692 B.n99 585
R1394 B.n694 B.n693 585
R1395 B.n695 B.n98 585
R1396 B.n697 B.n696 585
R1397 B.n698 B.n97 585
R1398 B.n700 B.n699 585
R1399 B.n701 B.n96 585
R1400 B.n703 B.n702 585
R1401 B.n704 B.n95 585
R1402 B.n706 B.n705 585
R1403 B.n707 B.n94 585
R1404 B.n709 B.n708 585
R1405 B.n874 B.n873 585
R1406 B.n872 B.n35 585
R1407 B.n871 B.n870 585
R1408 B.n869 B.n36 585
R1409 B.n868 B.n867 585
R1410 B.n866 B.n37 585
R1411 B.n865 B.n864 585
R1412 B.n863 B.n38 585
R1413 B.n862 B.n861 585
R1414 B.n860 B.n39 585
R1415 B.n859 B.n858 585
R1416 B.n857 B.n40 585
R1417 B.n856 B.n855 585
R1418 B.n854 B.n41 585
R1419 B.n853 B.n852 585
R1420 B.n851 B.n42 585
R1421 B.n850 B.n849 585
R1422 B.n848 B.n43 585
R1423 B.n847 B.n846 585
R1424 B.n845 B.n44 585
R1425 B.n844 B.n843 585
R1426 B.n842 B.n45 585
R1427 B.n841 B.n840 585
R1428 B.n839 B.n46 585
R1429 B.n838 B.n837 585
R1430 B.n836 B.n47 585
R1431 B.n835 B.n834 585
R1432 B.n833 B.n48 585
R1433 B.n832 B.n831 585
R1434 B.n830 B.n49 585
R1435 B.n829 B.n828 585
R1436 B.n827 B.n50 585
R1437 B.n826 B.n825 585
R1438 B.n824 B.n51 585
R1439 B.n823 B.n822 585
R1440 B.n821 B.n52 585
R1441 B.n820 B.n819 585
R1442 B.n818 B.n53 585
R1443 B.n817 B.n816 585
R1444 B.n815 B.n54 585
R1445 B.n814 B.n813 585
R1446 B.n812 B.n55 585
R1447 B.n811 B.n810 585
R1448 B.n809 B.n56 585
R1449 B.n808 B.n807 585
R1450 B.n806 B.n57 585
R1451 B.n805 B.n804 585
R1452 B.n803 B.n58 585
R1453 B.n802 B.n801 585
R1454 B.n800 B.n59 585
R1455 B.n798 B.n797 585
R1456 B.n796 B.n62 585
R1457 B.n795 B.n794 585
R1458 B.n793 B.n63 585
R1459 B.n792 B.n791 585
R1460 B.n790 B.n64 585
R1461 B.n789 B.n788 585
R1462 B.n787 B.n65 585
R1463 B.n786 B.n785 585
R1464 B.n784 B.n783 585
R1465 B.n782 B.n69 585
R1466 B.n781 B.n780 585
R1467 B.n779 B.n70 585
R1468 B.n778 B.n777 585
R1469 B.n776 B.n71 585
R1470 B.n775 B.n774 585
R1471 B.n773 B.n72 585
R1472 B.n772 B.n771 585
R1473 B.n770 B.n73 585
R1474 B.n769 B.n768 585
R1475 B.n767 B.n74 585
R1476 B.n766 B.n765 585
R1477 B.n764 B.n75 585
R1478 B.n763 B.n762 585
R1479 B.n761 B.n76 585
R1480 B.n760 B.n759 585
R1481 B.n758 B.n77 585
R1482 B.n757 B.n756 585
R1483 B.n755 B.n78 585
R1484 B.n754 B.n753 585
R1485 B.n752 B.n79 585
R1486 B.n751 B.n750 585
R1487 B.n749 B.n80 585
R1488 B.n748 B.n747 585
R1489 B.n746 B.n81 585
R1490 B.n745 B.n744 585
R1491 B.n743 B.n82 585
R1492 B.n742 B.n741 585
R1493 B.n740 B.n83 585
R1494 B.n739 B.n738 585
R1495 B.n737 B.n84 585
R1496 B.n736 B.n735 585
R1497 B.n734 B.n85 585
R1498 B.n733 B.n732 585
R1499 B.n731 B.n86 585
R1500 B.n730 B.n729 585
R1501 B.n728 B.n87 585
R1502 B.n727 B.n726 585
R1503 B.n725 B.n88 585
R1504 B.n724 B.n723 585
R1505 B.n722 B.n89 585
R1506 B.n721 B.n720 585
R1507 B.n719 B.n90 585
R1508 B.n718 B.n717 585
R1509 B.n716 B.n91 585
R1510 B.n715 B.n714 585
R1511 B.n713 B.n92 585
R1512 B.n712 B.n711 585
R1513 B.n710 B.n93 585
R1514 B.n875 B.n34 585
R1515 B.n877 B.n876 585
R1516 B.n878 B.n33 585
R1517 B.n880 B.n879 585
R1518 B.n881 B.n32 585
R1519 B.n883 B.n882 585
R1520 B.n884 B.n31 585
R1521 B.n886 B.n885 585
R1522 B.n887 B.n30 585
R1523 B.n889 B.n888 585
R1524 B.n890 B.n29 585
R1525 B.n892 B.n891 585
R1526 B.n893 B.n28 585
R1527 B.n895 B.n894 585
R1528 B.n896 B.n27 585
R1529 B.n898 B.n897 585
R1530 B.n899 B.n26 585
R1531 B.n901 B.n900 585
R1532 B.n902 B.n25 585
R1533 B.n904 B.n903 585
R1534 B.n905 B.n24 585
R1535 B.n907 B.n906 585
R1536 B.n908 B.n23 585
R1537 B.n910 B.n909 585
R1538 B.n911 B.n22 585
R1539 B.n913 B.n912 585
R1540 B.n914 B.n21 585
R1541 B.n916 B.n915 585
R1542 B.n917 B.n20 585
R1543 B.n919 B.n918 585
R1544 B.n920 B.n19 585
R1545 B.n922 B.n921 585
R1546 B.n923 B.n18 585
R1547 B.n925 B.n924 585
R1548 B.n926 B.n17 585
R1549 B.n928 B.n927 585
R1550 B.n929 B.n16 585
R1551 B.n931 B.n930 585
R1552 B.n932 B.n15 585
R1553 B.n934 B.n933 585
R1554 B.n935 B.n14 585
R1555 B.n937 B.n936 585
R1556 B.n938 B.n13 585
R1557 B.n940 B.n939 585
R1558 B.n941 B.n12 585
R1559 B.n943 B.n942 585
R1560 B.n944 B.n11 585
R1561 B.n946 B.n945 585
R1562 B.n947 B.n10 585
R1563 B.n949 B.n948 585
R1564 B.n950 B.n9 585
R1565 B.n952 B.n951 585
R1566 B.n953 B.n8 585
R1567 B.n955 B.n954 585
R1568 B.n956 B.n7 585
R1569 B.n958 B.n957 585
R1570 B.n959 B.n6 585
R1571 B.n961 B.n960 585
R1572 B.n962 B.n5 585
R1573 B.n964 B.n963 585
R1574 B.n965 B.n4 585
R1575 B.n967 B.n966 585
R1576 B.n968 B.n3 585
R1577 B.n970 B.n969 585
R1578 B.n971 B.n0 585
R1579 B.n2 B.n1 585
R1580 B.n249 B.n248 585
R1581 B.n250 B.n247 585
R1582 B.n252 B.n251 585
R1583 B.n253 B.n246 585
R1584 B.n255 B.n254 585
R1585 B.n256 B.n245 585
R1586 B.n258 B.n257 585
R1587 B.n259 B.n244 585
R1588 B.n261 B.n260 585
R1589 B.n262 B.n243 585
R1590 B.n264 B.n263 585
R1591 B.n265 B.n242 585
R1592 B.n267 B.n266 585
R1593 B.n268 B.n241 585
R1594 B.n270 B.n269 585
R1595 B.n271 B.n240 585
R1596 B.n273 B.n272 585
R1597 B.n274 B.n239 585
R1598 B.n276 B.n275 585
R1599 B.n277 B.n238 585
R1600 B.n279 B.n278 585
R1601 B.n280 B.n237 585
R1602 B.n282 B.n281 585
R1603 B.n283 B.n236 585
R1604 B.n285 B.n284 585
R1605 B.n286 B.n235 585
R1606 B.n288 B.n287 585
R1607 B.n289 B.n234 585
R1608 B.n291 B.n290 585
R1609 B.n292 B.n233 585
R1610 B.n294 B.n293 585
R1611 B.n295 B.n232 585
R1612 B.n297 B.n296 585
R1613 B.n298 B.n231 585
R1614 B.n300 B.n299 585
R1615 B.n301 B.n230 585
R1616 B.n303 B.n302 585
R1617 B.n304 B.n229 585
R1618 B.n306 B.n305 585
R1619 B.n307 B.n228 585
R1620 B.n309 B.n308 585
R1621 B.n310 B.n227 585
R1622 B.n312 B.n311 585
R1623 B.n313 B.n226 585
R1624 B.n315 B.n314 585
R1625 B.n316 B.n225 585
R1626 B.n318 B.n317 585
R1627 B.n319 B.n224 585
R1628 B.n321 B.n320 585
R1629 B.n322 B.n223 585
R1630 B.n324 B.n323 585
R1631 B.n325 B.n222 585
R1632 B.n327 B.n326 585
R1633 B.n328 B.n221 585
R1634 B.n330 B.n329 585
R1635 B.n331 B.n220 585
R1636 B.n333 B.n332 585
R1637 B.n334 B.n219 585
R1638 B.n336 B.n335 585
R1639 B.n337 B.n218 585
R1640 B.n339 B.n338 585
R1641 B.n340 B.n217 585
R1642 B.n342 B.n341 585
R1643 B.n343 B.n216 585
R1644 B.n344 B.n343 521.33
R1645 B.n510 B.n159 521.33
R1646 B.n708 B.n93 521.33
R1647 B.n875 B.n874 521.33
R1648 B.n432 B.t4 501.127
R1649 B.n66 B.t2 501.127
R1650 B.n190 B.t7 501.127
R1651 B.n60 B.t11 501.127
R1652 B.n433 B.t5 425.296
R1653 B.n67 B.t1 425.296
R1654 B.n191 B.t8 425.296
R1655 B.n61 B.t10 425.296
R1656 B.n190 B.t6 308.526
R1657 B.n432 B.t3 308.526
R1658 B.n66 B.t0 308.526
R1659 B.n60 B.t9 308.526
R1660 B.n973 B.n972 256.663
R1661 B.n972 B.n971 235.042
R1662 B.n972 B.n2 235.042
R1663 B.n344 B.n215 163.367
R1664 B.n348 B.n215 163.367
R1665 B.n349 B.n348 163.367
R1666 B.n350 B.n349 163.367
R1667 B.n350 B.n213 163.367
R1668 B.n354 B.n213 163.367
R1669 B.n355 B.n354 163.367
R1670 B.n356 B.n355 163.367
R1671 B.n356 B.n211 163.367
R1672 B.n360 B.n211 163.367
R1673 B.n361 B.n360 163.367
R1674 B.n362 B.n361 163.367
R1675 B.n362 B.n209 163.367
R1676 B.n366 B.n209 163.367
R1677 B.n367 B.n366 163.367
R1678 B.n368 B.n367 163.367
R1679 B.n368 B.n207 163.367
R1680 B.n372 B.n207 163.367
R1681 B.n373 B.n372 163.367
R1682 B.n374 B.n373 163.367
R1683 B.n374 B.n205 163.367
R1684 B.n378 B.n205 163.367
R1685 B.n379 B.n378 163.367
R1686 B.n380 B.n379 163.367
R1687 B.n380 B.n203 163.367
R1688 B.n384 B.n203 163.367
R1689 B.n385 B.n384 163.367
R1690 B.n386 B.n385 163.367
R1691 B.n386 B.n201 163.367
R1692 B.n390 B.n201 163.367
R1693 B.n391 B.n390 163.367
R1694 B.n392 B.n391 163.367
R1695 B.n392 B.n199 163.367
R1696 B.n396 B.n199 163.367
R1697 B.n397 B.n396 163.367
R1698 B.n398 B.n397 163.367
R1699 B.n398 B.n197 163.367
R1700 B.n402 B.n197 163.367
R1701 B.n403 B.n402 163.367
R1702 B.n404 B.n403 163.367
R1703 B.n404 B.n195 163.367
R1704 B.n408 B.n195 163.367
R1705 B.n409 B.n408 163.367
R1706 B.n410 B.n409 163.367
R1707 B.n410 B.n193 163.367
R1708 B.n414 B.n193 163.367
R1709 B.n415 B.n414 163.367
R1710 B.n416 B.n415 163.367
R1711 B.n416 B.n189 163.367
R1712 B.n421 B.n189 163.367
R1713 B.n422 B.n421 163.367
R1714 B.n423 B.n422 163.367
R1715 B.n423 B.n187 163.367
R1716 B.n427 B.n187 163.367
R1717 B.n428 B.n427 163.367
R1718 B.n429 B.n428 163.367
R1719 B.n429 B.n185 163.367
R1720 B.n436 B.n185 163.367
R1721 B.n437 B.n436 163.367
R1722 B.n438 B.n437 163.367
R1723 B.n438 B.n183 163.367
R1724 B.n442 B.n183 163.367
R1725 B.n443 B.n442 163.367
R1726 B.n444 B.n443 163.367
R1727 B.n444 B.n181 163.367
R1728 B.n448 B.n181 163.367
R1729 B.n449 B.n448 163.367
R1730 B.n450 B.n449 163.367
R1731 B.n450 B.n179 163.367
R1732 B.n454 B.n179 163.367
R1733 B.n455 B.n454 163.367
R1734 B.n456 B.n455 163.367
R1735 B.n456 B.n177 163.367
R1736 B.n460 B.n177 163.367
R1737 B.n461 B.n460 163.367
R1738 B.n462 B.n461 163.367
R1739 B.n462 B.n175 163.367
R1740 B.n466 B.n175 163.367
R1741 B.n467 B.n466 163.367
R1742 B.n468 B.n467 163.367
R1743 B.n468 B.n173 163.367
R1744 B.n472 B.n173 163.367
R1745 B.n473 B.n472 163.367
R1746 B.n474 B.n473 163.367
R1747 B.n474 B.n171 163.367
R1748 B.n478 B.n171 163.367
R1749 B.n479 B.n478 163.367
R1750 B.n480 B.n479 163.367
R1751 B.n480 B.n169 163.367
R1752 B.n484 B.n169 163.367
R1753 B.n485 B.n484 163.367
R1754 B.n486 B.n485 163.367
R1755 B.n486 B.n167 163.367
R1756 B.n490 B.n167 163.367
R1757 B.n491 B.n490 163.367
R1758 B.n492 B.n491 163.367
R1759 B.n492 B.n165 163.367
R1760 B.n496 B.n165 163.367
R1761 B.n497 B.n496 163.367
R1762 B.n498 B.n497 163.367
R1763 B.n498 B.n163 163.367
R1764 B.n502 B.n163 163.367
R1765 B.n503 B.n502 163.367
R1766 B.n504 B.n503 163.367
R1767 B.n504 B.n161 163.367
R1768 B.n508 B.n161 163.367
R1769 B.n509 B.n508 163.367
R1770 B.n510 B.n509 163.367
R1771 B.n708 B.n707 163.367
R1772 B.n707 B.n706 163.367
R1773 B.n706 B.n95 163.367
R1774 B.n702 B.n95 163.367
R1775 B.n702 B.n701 163.367
R1776 B.n701 B.n700 163.367
R1777 B.n700 B.n97 163.367
R1778 B.n696 B.n97 163.367
R1779 B.n696 B.n695 163.367
R1780 B.n695 B.n694 163.367
R1781 B.n694 B.n99 163.367
R1782 B.n690 B.n99 163.367
R1783 B.n690 B.n689 163.367
R1784 B.n689 B.n688 163.367
R1785 B.n688 B.n101 163.367
R1786 B.n684 B.n101 163.367
R1787 B.n684 B.n683 163.367
R1788 B.n683 B.n682 163.367
R1789 B.n682 B.n103 163.367
R1790 B.n678 B.n103 163.367
R1791 B.n678 B.n677 163.367
R1792 B.n677 B.n676 163.367
R1793 B.n676 B.n105 163.367
R1794 B.n672 B.n105 163.367
R1795 B.n672 B.n671 163.367
R1796 B.n671 B.n670 163.367
R1797 B.n670 B.n107 163.367
R1798 B.n666 B.n107 163.367
R1799 B.n666 B.n665 163.367
R1800 B.n665 B.n664 163.367
R1801 B.n664 B.n109 163.367
R1802 B.n660 B.n109 163.367
R1803 B.n660 B.n659 163.367
R1804 B.n659 B.n658 163.367
R1805 B.n658 B.n111 163.367
R1806 B.n654 B.n111 163.367
R1807 B.n654 B.n653 163.367
R1808 B.n653 B.n652 163.367
R1809 B.n652 B.n113 163.367
R1810 B.n648 B.n113 163.367
R1811 B.n648 B.n647 163.367
R1812 B.n647 B.n646 163.367
R1813 B.n646 B.n115 163.367
R1814 B.n642 B.n115 163.367
R1815 B.n642 B.n641 163.367
R1816 B.n641 B.n640 163.367
R1817 B.n640 B.n117 163.367
R1818 B.n636 B.n117 163.367
R1819 B.n636 B.n635 163.367
R1820 B.n635 B.n634 163.367
R1821 B.n634 B.n119 163.367
R1822 B.n630 B.n119 163.367
R1823 B.n630 B.n629 163.367
R1824 B.n629 B.n628 163.367
R1825 B.n628 B.n121 163.367
R1826 B.n624 B.n121 163.367
R1827 B.n624 B.n623 163.367
R1828 B.n623 B.n622 163.367
R1829 B.n622 B.n123 163.367
R1830 B.n618 B.n123 163.367
R1831 B.n618 B.n617 163.367
R1832 B.n617 B.n616 163.367
R1833 B.n616 B.n125 163.367
R1834 B.n612 B.n125 163.367
R1835 B.n612 B.n611 163.367
R1836 B.n611 B.n610 163.367
R1837 B.n610 B.n127 163.367
R1838 B.n606 B.n127 163.367
R1839 B.n606 B.n605 163.367
R1840 B.n605 B.n604 163.367
R1841 B.n604 B.n129 163.367
R1842 B.n600 B.n129 163.367
R1843 B.n600 B.n599 163.367
R1844 B.n599 B.n598 163.367
R1845 B.n598 B.n131 163.367
R1846 B.n594 B.n131 163.367
R1847 B.n594 B.n593 163.367
R1848 B.n593 B.n592 163.367
R1849 B.n592 B.n133 163.367
R1850 B.n588 B.n133 163.367
R1851 B.n588 B.n587 163.367
R1852 B.n587 B.n586 163.367
R1853 B.n586 B.n135 163.367
R1854 B.n582 B.n135 163.367
R1855 B.n582 B.n581 163.367
R1856 B.n581 B.n580 163.367
R1857 B.n580 B.n137 163.367
R1858 B.n576 B.n137 163.367
R1859 B.n576 B.n575 163.367
R1860 B.n575 B.n574 163.367
R1861 B.n574 B.n139 163.367
R1862 B.n570 B.n139 163.367
R1863 B.n570 B.n569 163.367
R1864 B.n569 B.n568 163.367
R1865 B.n568 B.n141 163.367
R1866 B.n564 B.n141 163.367
R1867 B.n564 B.n563 163.367
R1868 B.n563 B.n562 163.367
R1869 B.n562 B.n143 163.367
R1870 B.n558 B.n143 163.367
R1871 B.n558 B.n557 163.367
R1872 B.n557 B.n556 163.367
R1873 B.n556 B.n145 163.367
R1874 B.n552 B.n145 163.367
R1875 B.n552 B.n551 163.367
R1876 B.n551 B.n550 163.367
R1877 B.n550 B.n147 163.367
R1878 B.n546 B.n147 163.367
R1879 B.n546 B.n545 163.367
R1880 B.n545 B.n544 163.367
R1881 B.n544 B.n149 163.367
R1882 B.n540 B.n149 163.367
R1883 B.n540 B.n539 163.367
R1884 B.n539 B.n538 163.367
R1885 B.n538 B.n151 163.367
R1886 B.n534 B.n151 163.367
R1887 B.n534 B.n533 163.367
R1888 B.n533 B.n532 163.367
R1889 B.n532 B.n153 163.367
R1890 B.n528 B.n153 163.367
R1891 B.n528 B.n527 163.367
R1892 B.n527 B.n526 163.367
R1893 B.n526 B.n155 163.367
R1894 B.n522 B.n155 163.367
R1895 B.n522 B.n521 163.367
R1896 B.n521 B.n520 163.367
R1897 B.n520 B.n157 163.367
R1898 B.n516 B.n157 163.367
R1899 B.n516 B.n515 163.367
R1900 B.n515 B.n514 163.367
R1901 B.n514 B.n159 163.367
R1902 B.n874 B.n35 163.367
R1903 B.n870 B.n35 163.367
R1904 B.n870 B.n869 163.367
R1905 B.n869 B.n868 163.367
R1906 B.n868 B.n37 163.367
R1907 B.n864 B.n37 163.367
R1908 B.n864 B.n863 163.367
R1909 B.n863 B.n862 163.367
R1910 B.n862 B.n39 163.367
R1911 B.n858 B.n39 163.367
R1912 B.n858 B.n857 163.367
R1913 B.n857 B.n856 163.367
R1914 B.n856 B.n41 163.367
R1915 B.n852 B.n41 163.367
R1916 B.n852 B.n851 163.367
R1917 B.n851 B.n850 163.367
R1918 B.n850 B.n43 163.367
R1919 B.n846 B.n43 163.367
R1920 B.n846 B.n845 163.367
R1921 B.n845 B.n844 163.367
R1922 B.n844 B.n45 163.367
R1923 B.n840 B.n45 163.367
R1924 B.n840 B.n839 163.367
R1925 B.n839 B.n838 163.367
R1926 B.n838 B.n47 163.367
R1927 B.n834 B.n47 163.367
R1928 B.n834 B.n833 163.367
R1929 B.n833 B.n832 163.367
R1930 B.n832 B.n49 163.367
R1931 B.n828 B.n49 163.367
R1932 B.n828 B.n827 163.367
R1933 B.n827 B.n826 163.367
R1934 B.n826 B.n51 163.367
R1935 B.n822 B.n51 163.367
R1936 B.n822 B.n821 163.367
R1937 B.n821 B.n820 163.367
R1938 B.n820 B.n53 163.367
R1939 B.n816 B.n53 163.367
R1940 B.n816 B.n815 163.367
R1941 B.n815 B.n814 163.367
R1942 B.n814 B.n55 163.367
R1943 B.n810 B.n55 163.367
R1944 B.n810 B.n809 163.367
R1945 B.n809 B.n808 163.367
R1946 B.n808 B.n57 163.367
R1947 B.n804 B.n57 163.367
R1948 B.n804 B.n803 163.367
R1949 B.n803 B.n802 163.367
R1950 B.n802 B.n59 163.367
R1951 B.n797 B.n59 163.367
R1952 B.n797 B.n796 163.367
R1953 B.n796 B.n795 163.367
R1954 B.n795 B.n63 163.367
R1955 B.n791 B.n63 163.367
R1956 B.n791 B.n790 163.367
R1957 B.n790 B.n789 163.367
R1958 B.n789 B.n65 163.367
R1959 B.n785 B.n65 163.367
R1960 B.n785 B.n784 163.367
R1961 B.n784 B.n69 163.367
R1962 B.n780 B.n69 163.367
R1963 B.n780 B.n779 163.367
R1964 B.n779 B.n778 163.367
R1965 B.n778 B.n71 163.367
R1966 B.n774 B.n71 163.367
R1967 B.n774 B.n773 163.367
R1968 B.n773 B.n772 163.367
R1969 B.n772 B.n73 163.367
R1970 B.n768 B.n73 163.367
R1971 B.n768 B.n767 163.367
R1972 B.n767 B.n766 163.367
R1973 B.n766 B.n75 163.367
R1974 B.n762 B.n75 163.367
R1975 B.n762 B.n761 163.367
R1976 B.n761 B.n760 163.367
R1977 B.n760 B.n77 163.367
R1978 B.n756 B.n77 163.367
R1979 B.n756 B.n755 163.367
R1980 B.n755 B.n754 163.367
R1981 B.n754 B.n79 163.367
R1982 B.n750 B.n79 163.367
R1983 B.n750 B.n749 163.367
R1984 B.n749 B.n748 163.367
R1985 B.n748 B.n81 163.367
R1986 B.n744 B.n81 163.367
R1987 B.n744 B.n743 163.367
R1988 B.n743 B.n742 163.367
R1989 B.n742 B.n83 163.367
R1990 B.n738 B.n83 163.367
R1991 B.n738 B.n737 163.367
R1992 B.n737 B.n736 163.367
R1993 B.n736 B.n85 163.367
R1994 B.n732 B.n85 163.367
R1995 B.n732 B.n731 163.367
R1996 B.n731 B.n730 163.367
R1997 B.n730 B.n87 163.367
R1998 B.n726 B.n87 163.367
R1999 B.n726 B.n725 163.367
R2000 B.n725 B.n724 163.367
R2001 B.n724 B.n89 163.367
R2002 B.n720 B.n89 163.367
R2003 B.n720 B.n719 163.367
R2004 B.n719 B.n718 163.367
R2005 B.n718 B.n91 163.367
R2006 B.n714 B.n91 163.367
R2007 B.n714 B.n713 163.367
R2008 B.n713 B.n712 163.367
R2009 B.n712 B.n93 163.367
R2010 B.n876 B.n875 163.367
R2011 B.n876 B.n33 163.367
R2012 B.n880 B.n33 163.367
R2013 B.n881 B.n880 163.367
R2014 B.n882 B.n881 163.367
R2015 B.n882 B.n31 163.367
R2016 B.n886 B.n31 163.367
R2017 B.n887 B.n886 163.367
R2018 B.n888 B.n887 163.367
R2019 B.n888 B.n29 163.367
R2020 B.n892 B.n29 163.367
R2021 B.n893 B.n892 163.367
R2022 B.n894 B.n893 163.367
R2023 B.n894 B.n27 163.367
R2024 B.n898 B.n27 163.367
R2025 B.n899 B.n898 163.367
R2026 B.n900 B.n899 163.367
R2027 B.n900 B.n25 163.367
R2028 B.n904 B.n25 163.367
R2029 B.n905 B.n904 163.367
R2030 B.n906 B.n905 163.367
R2031 B.n906 B.n23 163.367
R2032 B.n910 B.n23 163.367
R2033 B.n911 B.n910 163.367
R2034 B.n912 B.n911 163.367
R2035 B.n912 B.n21 163.367
R2036 B.n916 B.n21 163.367
R2037 B.n917 B.n916 163.367
R2038 B.n918 B.n917 163.367
R2039 B.n918 B.n19 163.367
R2040 B.n922 B.n19 163.367
R2041 B.n923 B.n922 163.367
R2042 B.n924 B.n923 163.367
R2043 B.n924 B.n17 163.367
R2044 B.n928 B.n17 163.367
R2045 B.n929 B.n928 163.367
R2046 B.n930 B.n929 163.367
R2047 B.n930 B.n15 163.367
R2048 B.n934 B.n15 163.367
R2049 B.n935 B.n934 163.367
R2050 B.n936 B.n935 163.367
R2051 B.n936 B.n13 163.367
R2052 B.n940 B.n13 163.367
R2053 B.n941 B.n940 163.367
R2054 B.n942 B.n941 163.367
R2055 B.n942 B.n11 163.367
R2056 B.n946 B.n11 163.367
R2057 B.n947 B.n946 163.367
R2058 B.n948 B.n947 163.367
R2059 B.n948 B.n9 163.367
R2060 B.n952 B.n9 163.367
R2061 B.n953 B.n952 163.367
R2062 B.n954 B.n953 163.367
R2063 B.n954 B.n7 163.367
R2064 B.n958 B.n7 163.367
R2065 B.n959 B.n958 163.367
R2066 B.n960 B.n959 163.367
R2067 B.n960 B.n5 163.367
R2068 B.n964 B.n5 163.367
R2069 B.n965 B.n964 163.367
R2070 B.n966 B.n965 163.367
R2071 B.n966 B.n3 163.367
R2072 B.n970 B.n3 163.367
R2073 B.n971 B.n970 163.367
R2074 B.n248 B.n2 163.367
R2075 B.n248 B.n247 163.367
R2076 B.n252 B.n247 163.367
R2077 B.n253 B.n252 163.367
R2078 B.n254 B.n253 163.367
R2079 B.n254 B.n245 163.367
R2080 B.n258 B.n245 163.367
R2081 B.n259 B.n258 163.367
R2082 B.n260 B.n259 163.367
R2083 B.n260 B.n243 163.367
R2084 B.n264 B.n243 163.367
R2085 B.n265 B.n264 163.367
R2086 B.n266 B.n265 163.367
R2087 B.n266 B.n241 163.367
R2088 B.n270 B.n241 163.367
R2089 B.n271 B.n270 163.367
R2090 B.n272 B.n271 163.367
R2091 B.n272 B.n239 163.367
R2092 B.n276 B.n239 163.367
R2093 B.n277 B.n276 163.367
R2094 B.n278 B.n277 163.367
R2095 B.n278 B.n237 163.367
R2096 B.n282 B.n237 163.367
R2097 B.n283 B.n282 163.367
R2098 B.n284 B.n283 163.367
R2099 B.n284 B.n235 163.367
R2100 B.n288 B.n235 163.367
R2101 B.n289 B.n288 163.367
R2102 B.n290 B.n289 163.367
R2103 B.n290 B.n233 163.367
R2104 B.n294 B.n233 163.367
R2105 B.n295 B.n294 163.367
R2106 B.n296 B.n295 163.367
R2107 B.n296 B.n231 163.367
R2108 B.n300 B.n231 163.367
R2109 B.n301 B.n300 163.367
R2110 B.n302 B.n301 163.367
R2111 B.n302 B.n229 163.367
R2112 B.n306 B.n229 163.367
R2113 B.n307 B.n306 163.367
R2114 B.n308 B.n307 163.367
R2115 B.n308 B.n227 163.367
R2116 B.n312 B.n227 163.367
R2117 B.n313 B.n312 163.367
R2118 B.n314 B.n313 163.367
R2119 B.n314 B.n225 163.367
R2120 B.n318 B.n225 163.367
R2121 B.n319 B.n318 163.367
R2122 B.n320 B.n319 163.367
R2123 B.n320 B.n223 163.367
R2124 B.n324 B.n223 163.367
R2125 B.n325 B.n324 163.367
R2126 B.n326 B.n325 163.367
R2127 B.n326 B.n221 163.367
R2128 B.n330 B.n221 163.367
R2129 B.n331 B.n330 163.367
R2130 B.n332 B.n331 163.367
R2131 B.n332 B.n219 163.367
R2132 B.n336 B.n219 163.367
R2133 B.n337 B.n336 163.367
R2134 B.n338 B.n337 163.367
R2135 B.n338 B.n217 163.367
R2136 B.n342 B.n217 163.367
R2137 B.n343 B.n342 163.367
R2138 B.n191 B.n190 75.8308
R2139 B.n433 B.n432 75.8308
R2140 B.n67 B.n66 75.8308
R2141 B.n61 B.n60 75.8308
R2142 B.n419 B.n191 59.5399
R2143 B.n434 B.n433 59.5399
R2144 B.n68 B.n67 59.5399
R2145 B.n799 B.n61 59.5399
R2146 B.n873 B.n34 33.8737
R2147 B.n710 B.n709 33.8737
R2148 B.n512 B.n511 33.8737
R2149 B.n345 B.n216 33.8737
R2150 B B.n973 18.0485
R2151 B.n877 B.n34 10.6151
R2152 B.n878 B.n877 10.6151
R2153 B.n879 B.n878 10.6151
R2154 B.n879 B.n32 10.6151
R2155 B.n883 B.n32 10.6151
R2156 B.n884 B.n883 10.6151
R2157 B.n885 B.n884 10.6151
R2158 B.n885 B.n30 10.6151
R2159 B.n889 B.n30 10.6151
R2160 B.n890 B.n889 10.6151
R2161 B.n891 B.n890 10.6151
R2162 B.n891 B.n28 10.6151
R2163 B.n895 B.n28 10.6151
R2164 B.n896 B.n895 10.6151
R2165 B.n897 B.n896 10.6151
R2166 B.n897 B.n26 10.6151
R2167 B.n901 B.n26 10.6151
R2168 B.n902 B.n901 10.6151
R2169 B.n903 B.n902 10.6151
R2170 B.n903 B.n24 10.6151
R2171 B.n907 B.n24 10.6151
R2172 B.n908 B.n907 10.6151
R2173 B.n909 B.n908 10.6151
R2174 B.n909 B.n22 10.6151
R2175 B.n913 B.n22 10.6151
R2176 B.n914 B.n913 10.6151
R2177 B.n915 B.n914 10.6151
R2178 B.n915 B.n20 10.6151
R2179 B.n919 B.n20 10.6151
R2180 B.n920 B.n919 10.6151
R2181 B.n921 B.n920 10.6151
R2182 B.n921 B.n18 10.6151
R2183 B.n925 B.n18 10.6151
R2184 B.n926 B.n925 10.6151
R2185 B.n927 B.n926 10.6151
R2186 B.n927 B.n16 10.6151
R2187 B.n931 B.n16 10.6151
R2188 B.n932 B.n931 10.6151
R2189 B.n933 B.n932 10.6151
R2190 B.n933 B.n14 10.6151
R2191 B.n937 B.n14 10.6151
R2192 B.n938 B.n937 10.6151
R2193 B.n939 B.n938 10.6151
R2194 B.n939 B.n12 10.6151
R2195 B.n943 B.n12 10.6151
R2196 B.n944 B.n943 10.6151
R2197 B.n945 B.n944 10.6151
R2198 B.n945 B.n10 10.6151
R2199 B.n949 B.n10 10.6151
R2200 B.n950 B.n949 10.6151
R2201 B.n951 B.n950 10.6151
R2202 B.n951 B.n8 10.6151
R2203 B.n955 B.n8 10.6151
R2204 B.n956 B.n955 10.6151
R2205 B.n957 B.n956 10.6151
R2206 B.n957 B.n6 10.6151
R2207 B.n961 B.n6 10.6151
R2208 B.n962 B.n961 10.6151
R2209 B.n963 B.n962 10.6151
R2210 B.n963 B.n4 10.6151
R2211 B.n967 B.n4 10.6151
R2212 B.n968 B.n967 10.6151
R2213 B.n969 B.n968 10.6151
R2214 B.n969 B.n0 10.6151
R2215 B.n873 B.n872 10.6151
R2216 B.n872 B.n871 10.6151
R2217 B.n871 B.n36 10.6151
R2218 B.n867 B.n36 10.6151
R2219 B.n867 B.n866 10.6151
R2220 B.n866 B.n865 10.6151
R2221 B.n865 B.n38 10.6151
R2222 B.n861 B.n38 10.6151
R2223 B.n861 B.n860 10.6151
R2224 B.n860 B.n859 10.6151
R2225 B.n859 B.n40 10.6151
R2226 B.n855 B.n40 10.6151
R2227 B.n855 B.n854 10.6151
R2228 B.n854 B.n853 10.6151
R2229 B.n853 B.n42 10.6151
R2230 B.n849 B.n42 10.6151
R2231 B.n849 B.n848 10.6151
R2232 B.n848 B.n847 10.6151
R2233 B.n847 B.n44 10.6151
R2234 B.n843 B.n44 10.6151
R2235 B.n843 B.n842 10.6151
R2236 B.n842 B.n841 10.6151
R2237 B.n841 B.n46 10.6151
R2238 B.n837 B.n46 10.6151
R2239 B.n837 B.n836 10.6151
R2240 B.n836 B.n835 10.6151
R2241 B.n835 B.n48 10.6151
R2242 B.n831 B.n48 10.6151
R2243 B.n831 B.n830 10.6151
R2244 B.n830 B.n829 10.6151
R2245 B.n829 B.n50 10.6151
R2246 B.n825 B.n50 10.6151
R2247 B.n825 B.n824 10.6151
R2248 B.n824 B.n823 10.6151
R2249 B.n823 B.n52 10.6151
R2250 B.n819 B.n52 10.6151
R2251 B.n819 B.n818 10.6151
R2252 B.n818 B.n817 10.6151
R2253 B.n817 B.n54 10.6151
R2254 B.n813 B.n54 10.6151
R2255 B.n813 B.n812 10.6151
R2256 B.n812 B.n811 10.6151
R2257 B.n811 B.n56 10.6151
R2258 B.n807 B.n56 10.6151
R2259 B.n807 B.n806 10.6151
R2260 B.n806 B.n805 10.6151
R2261 B.n805 B.n58 10.6151
R2262 B.n801 B.n58 10.6151
R2263 B.n801 B.n800 10.6151
R2264 B.n798 B.n62 10.6151
R2265 B.n794 B.n62 10.6151
R2266 B.n794 B.n793 10.6151
R2267 B.n793 B.n792 10.6151
R2268 B.n792 B.n64 10.6151
R2269 B.n788 B.n64 10.6151
R2270 B.n788 B.n787 10.6151
R2271 B.n787 B.n786 10.6151
R2272 B.n783 B.n782 10.6151
R2273 B.n782 B.n781 10.6151
R2274 B.n781 B.n70 10.6151
R2275 B.n777 B.n70 10.6151
R2276 B.n777 B.n776 10.6151
R2277 B.n776 B.n775 10.6151
R2278 B.n775 B.n72 10.6151
R2279 B.n771 B.n72 10.6151
R2280 B.n771 B.n770 10.6151
R2281 B.n770 B.n769 10.6151
R2282 B.n769 B.n74 10.6151
R2283 B.n765 B.n74 10.6151
R2284 B.n765 B.n764 10.6151
R2285 B.n764 B.n763 10.6151
R2286 B.n763 B.n76 10.6151
R2287 B.n759 B.n76 10.6151
R2288 B.n759 B.n758 10.6151
R2289 B.n758 B.n757 10.6151
R2290 B.n757 B.n78 10.6151
R2291 B.n753 B.n78 10.6151
R2292 B.n753 B.n752 10.6151
R2293 B.n752 B.n751 10.6151
R2294 B.n751 B.n80 10.6151
R2295 B.n747 B.n80 10.6151
R2296 B.n747 B.n746 10.6151
R2297 B.n746 B.n745 10.6151
R2298 B.n745 B.n82 10.6151
R2299 B.n741 B.n82 10.6151
R2300 B.n741 B.n740 10.6151
R2301 B.n740 B.n739 10.6151
R2302 B.n739 B.n84 10.6151
R2303 B.n735 B.n84 10.6151
R2304 B.n735 B.n734 10.6151
R2305 B.n734 B.n733 10.6151
R2306 B.n733 B.n86 10.6151
R2307 B.n729 B.n86 10.6151
R2308 B.n729 B.n728 10.6151
R2309 B.n728 B.n727 10.6151
R2310 B.n727 B.n88 10.6151
R2311 B.n723 B.n88 10.6151
R2312 B.n723 B.n722 10.6151
R2313 B.n722 B.n721 10.6151
R2314 B.n721 B.n90 10.6151
R2315 B.n717 B.n90 10.6151
R2316 B.n717 B.n716 10.6151
R2317 B.n716 B.n715 10.6151
R2318 B.n715 B.n92 10.6151
R2319 B.n711 B.n92 10.6151
R2320 B.n711 B.n710 10.6151
R2321 B.n709 B.n94 10.6151
R2322 B.n705 B.n94 10.6151
R2323 B.n705 B.n704 10.6151
R2324 B.n704 B.n703 10.6151
R2325 B.n703 B.n96 10.6151
R2326 B.n699 B.n96 10.6151
R2327 B.n699 B.n698 10.6151
R2328 B.n698 B.n697 10.6151
R2329 B.n697 B.n98 10.6151
R2330 B.n693 B.n98 10.6151
R2331 B.n693 B.n692 10.6151
R2332 B.n692 B.n691 10.6151
R2333 B.n691 B.n100 10.6151
R2334 B.n687 B.n100 10.6151
R2335 B.n687 B.n686 10.6151
R2336 B.n686 B.n685 10.6151
R2337 B.n685 B.n102 10.6151
R2338 B.n681 B.n102 10.6151
R2339 B.n681 B.n680 10.6151
R2340 B.n680 B.n679 10.6151
R2341 B.n679 B.n104 10.6151
R2342 B.n675 B.n104 10.6151
R2343 B.n675 B.n674 10.6151
R2344 B.n674 B.n673 10.6151
R2345 B.n673 B.n106 10.6151
R2346 B.n669 B.n106 10.6151
R2347 B.n669 B.n668 10.6151
R2348 B.n668 B.n667 10.6151
R2349 B.n667 B.n108 10.6151
R2350 B.n663 B.n108 10.6151
R2351 B.n663 B.n662 10.6151
R2352 B.n662 B.n661 10.6151
R2353 B.n661 B.n110 10.6151
R2354 B.n657 B.n110 10.6151
R2355 B.n657 B.n656 10.6151
R2356 B.n656 B.n655 10.6151
R2357 B.n655 B.n112 10.6151
R2358 B.n651 B.n112 10.6151
R2359 B.n651 B.n650 10.6151
R2360 B.n650 B.n649 10.6151
R2361 B.n649 B.n114 10.6151
R2362 B.n645 B.n114 10.6151
R2363 B.n645 B.n644 10.6151
R2364 B.n644 B.n643 10.6151
R2365 B.n643 B.n116 10.6151
R2366 B.n639 B.n116 10.6151
R2367 B.n639 B.n638 10.6151
R2368 B.n638 B.n637 10.6151
R2369 B.n637 B.n118 10.6151
R2370 B.n633 B.n118 10.6151
R2371 B.n633 B.n632 10.6151
R2372 B.n632 B.n631 10.6151
R2373 B.n631 B.n120 10.6151
R2374 B.n627 B.n120 10.6151
R2375 B.n627 B.n626 10.6151
R2376 B.n626 B.n625 10.6151
R2377 B.n625 B.n122 10.6151
R2378 B.n621 B.n122 10.6151
R2379 B.n621 B.n620 10.6151
R2380 B.n620 B.n619 10.6151
R2381 B.n619 B.n124 10.6151
R2382 B.n615 B.n124 10.6151
R2383 B.n615 B.n614 10.6151
R2384 B.n614 B.n613 10.6151
R2385 B.n613 B.n126 10.6151
R2386 B.n609 B.n126 10.6151
R2387 B.n609 B.n608 10.6151
R2388 B.n608 B.n607 10.6151
R2389 B.n607 B.n128 10.6151
R2390 B.n603 B.n128 10.6151
R2391 B.n603 B.n602 10.6151
R2392 B.n602 B.n601 10.6151
R2393 B.n601 B.n130 10.6151
R2394 B.n597 B.n130 10.6151
R2395 B.n597 B.n596 10.6151
R2396 B.n596 B.n595 10.6151
R2397 B.n595 B.n132 10.6151
R2398 B.n591 B.n132 10.6151
R2399 B.n591 B.n590 10.6151
R2400 B.n590 B.n589 10.6151
R2401 B.n589 B.n134 10.6151
R2402 B.n585 B.n134 10.6151
R2403 B.n585 B.n584 10.6151
R2404 B.n584 B.n583 10.6151
R2405 B.n583 B.n136 10.6151
R2406 B.n579 B.n136 10.6151
R2407 B.n579 B.n578 10.6151
R2408 B.n578 B.n577 10.6151
R2409 B.n577 B.n138 10.6151
R2410 B.n573 B.n138 10.6151
R2411 B.n573 B.n572 10.6151
R2412 B.n572 B.n571 10.6151
R2413 B.n571 B.n140 10.6151
R2414 B.n567 B.n140 10.6151
R2415 B.n567 B.n566 10.6151
R2416 B.n566 B.n565 10.6151
R2417 B.n565 B.n142 10.6151
R2418 B.n561 B.n142 10.6151
R2419 B.n561 B.n560 10.6151
R2420 B.n560 B.n559 10.6151
R2421 B.n559 B.n144 10.6151
R2422 B.n555 B.n144 10.6151
R2423 B.n555 B.n554 10.6151
R2424 B.n554 B.n553 10.6151
R2425 B.n553 B.n146 10.6151
R2426 B.n549 B.n146 10.6151
R2427 B.n549 B.n548 10.6151
R2428 B.n548 B.n547 10.6151
R2429 B.n547 B.n148 10.6151
R2430 B.n543 B.n148 10.6151
R2431 B.n543 B.n542 10.6151
R2432 B.n542 B.n541 10.6151
R2433 B.n541 B.n150 10.6151
R2434 B.n537 B.n150 10.6151
R2435 B.n537 B.n536 10.6151
R2436 B.n536 B.n535 10.6151
R2437 B.n535 B.n152 10.6151
R2438 B.n531 B.n152 10.6151
R2439 B.n531 B.n530 10.6151
R2440 B.n530 B.n529 10.6151
R2441 B.n529 B.n154 10.6151
R2442 B.n525 B.n154 10.6151
R2443 B.n525 B.n524 10.6151
R2444 B.n524 B.n523 10.6151
R2445 B.n523 B.n156 10.6151
R2446 B.n519 B.n156 10.6151
R2447 B.n519 B.n518 10.6151
R2448 B.n518 B.n517 10.6151
R2449 B.n517 B.n158 10.6151
R2450 B.n513 B.n158 10.6151
R2451 B.n513 B.n512 10.6151
R2452 B.n249 B.n1 10.6151
R2453 B.n250 B.n249 10.6151
R2454 B.n251 B.n250 10.6151
R2455 B.n251 B.n246 10.6151
R2456 B.n255 B.n246 10.6151
R2457 B.n256 B.n255 10.6151
R2458 B.n257 B.n256 10.6151
R2459 B.n257 B.n244 10.6151
R2460 B.n261 B.n244 10.6151
R2461 B.n262 B.n261 10.6151
R2462 B.n263 B.n262 10.6151
R2463 B.n263 B.n242 10.6151
R2464 B.n267 B.n242 10.6151
R2465 B.n268 B.n267 10.6151
R2466 B.n269 B.n268 10.6151
R2467 B.n269 B.n240 10.6151
R2468 B.n273 B.n240 10.6151
R2469 B.n274 B.n273 10.6151
R2470 B.n275 B.n274 10.6151
R2471 B.n275 B.n238 10.6151
R2472 B.n279 B.n238 10.6151
R2473 B.n280 B.n279 10.6151
R2474 B.n281 B.n280 10.6151
R2475 B.n281 B.n236 10.6151
R2476 B.n285 B.n236 10.6151
R2477 B.n286 B.n285 10.6151
R2478 B.n287 B.n286 10.6151
R2479 B.n287 B.n234 10.6151
R2480 B.n291 B.n234 10.6151
R2481 B.n292 B.n291 10.6151
R2482 B.n293 B.n292 10.6151
R2483 B.n293 B.n232 10.6151
R2484 B.n297 B.n232 10.6151
R2485 B.n298 B.n297 10.6151
R2486 B.n299 B.n298 10.6151
R2487 B.n299 B.n230 10.6151
R2488 B.n303 B.n230 10.6151
R2489 B.n304 B.n303 10.6151
R2490 B.n305 B.n304 10.6151
R2491 B.n305 B.n228 10.6151
R2492 B.n309 B.n228 10.6151
R2493 B.n310 B.n309 10.6151
R2494 B.n311 B.n310 10.6151
R2495 B.n311 B.n226 10.6151
R2496 B.n315 B.n226 10.6151
R2497 B.n316 B.n315 10.6151
R2498 B.n317 B.n316 10.6151
R2499 B.n317 B.n224 10.6151
R2500 B.n321 B.n224 10.6151
R2501 B.n322 B.n321 10.6151
R2502 B.n323 B.n322 10.6151
R2503 B.n323 B.n222 10.6151
R2504 B.n327 B.n222 10.6151
R2505 B.n328 B.n327 10.6151
R2506 B.n329 B.n328 10.6151
R2507 B.n329 B.n220 10.6151
R2508 B.n333 B.n220 10.6151
R2509 B.n334 B.n333 10.6151
R2510 B.n335 B.n334 10.6151
R2511 B.n335 B.n218 10.6151
R2512 B.n339 B.n218 10.6151
R2513 B.n340 B.n339 10.6151
R2514 B.n341 B.n340 10.6151
R2515 B.n341 B.n216 10.6151
R2516 B.n346 B.n345 10.6151
R2517 B.n347 B.n346 10.6151
R2518 B.n347 B.n214 10.6151
R2519 B.n351 B.n214 10.6151
R2520 B.n352 B.n351 10.6151
R2521 B.n353 B.n352 10.6151
R2522 B.n353 B.n212 10.6151
R2523 B.n357 B.n212 10.6151
R2524 B.n358 B.n357 10.6151
R2525 B.n359 B.n358 10.6151
R2526 B.n359 B.n210 10.6151
R2527 B.n363 B.n210 10.6151
R2528 B.n364 B.n363 10.6151
R2529 B.n365 B.n364 10.6151
R2530 B.n365 B.n208 10.6151
R2531 B.n369 B.n208 10.6151
R2532 B.n370 B.n369 10.6151
R2533 B.n371 B.n370 10.6151
R2534 B.n371 B.n206 10.6151
R2535 B.n375 B.n206 10.6151
R2536 B.n376 B.n375 10.6151
R2537 B.n377 B.n376 10.6151
R2538 B.n377 B.n204 10.6151
R2539 B.n381 B.n204 10.6151
R2540 B.n382 B.n381 10.6151
R2541 B.n383 B.n382 10.6151
R2542 B.n383 B.n202 10.6151
R2543 B.n387 B.n202 10.6151
R2544 B.n388 B.n387 10.6151
R2545 B.n389 B.n388 10.6151
R2546 B.n389 B.n200 10.6151
R2547 B.n393 B.n200 10.6151
R2548 B.n394 B.n393 10.6151
R2549 B.n395 B.n394 10.6151
R2550 B.n395 B.n198 10.6151
R2551 B.n399 B.n198 10.6151
R2552 B.n400 B.n399 10.6151
R2553 B.n401 B.n400 10.6151
R2554 B.n401 B.n196 10.6151
R2555 B.n405 B.n196 10.6151
R2556 B.n406 B.n405 10.6151
R2557 B.n407 B.n406 10.6151
R2558 B.n407 B.n194 10.6151
R2559 B.n411 B.n194 10.6151
R2560 B.n412 B.n411 10.6151
R2561 B.n413 B.n412 10.6151
R2562 B.n413 B.n192 10.6151
R2563 B.n417 B.n192 10.6151
R2564 B.n418 B.n417 10.6151
R2565 B.n420 B.n188 10.6151
R2566 B.n424 B.n188 10.6151
R2567 B.n425 B.n424 10.6151
R2568 B.n426 B.n425 10.6151
R2569 B.n426 B.n186 10.6151
R2570 B.n430 B.n186 10.6151
R2571 B.n431 B.n430 10.6151
R2572 B.n435 B.n431 10.6151
R2573 B.n439 B.n184 10.6151
R2574 B.n440 B.n439 10.6151
R2575 B.n441 B.n440 10.6151
R2576 B.n441 B.n182 10.6151
R2577 B.n445 B.n182 10.6151
R2578 B.n446 B.n445 10.6151
R2579 B.n447 B.n446 10.6151
R2580 B.n447 B.n180 10.6151
R2581 B.n451 B.n180 10.6151
R2582 B.n452 B.n451 10.6151
R2583 B.n453 B.n452 10.6151
R2584 B.n453 B.n178 10.6151
R2585 B.n457 B.n178 10.6151
R2586 B.n458 B.n457 10.6151
R2587 B.n459 B.n458 10.6151
R2588 B.n459 B.n176 10.6151
R2589 B.n463 B.n176 10.6151
R2590 B.n464 B.n463 10.6151
R2591 B.n465 B.n464 10.6151
R2592 B.n465 B.n174 10.6151
R2593 B.n469 B.n174 10.6151
R2594 B.n470 B.n469 10.6151
R2595 B.n471 B.n470 10.6151
R2596 B.n471 B.n172 10.6151
R2597 B.n475 B.n172 10.6151
R2598 B.n476 B.n475 10.6151
R2599 B.n477 B.n476 10.6151
R2600 B.n477 B.n170 10.6151
R2601 B.n481 B.n170 10.6151
R2602 B.n482 B.n481 10.6151
R2603 B.n483 B.n482 10.6151
R2604 B.n483 B.n168 10.6151
R2605 B.n487 B.n168 10.6151
R2606 B.n488 B.n487 10.6151
R2607 B.n489 B.n488 10.6151
R2608 B.n489 B.n166 10.6151
R2609 B.n493 B.n166 10.6151
R2610 B.n494 B.n493 10.6151
R2611 B.n495 B.n494 10.6151
R2612 B.n495 B.n164 10.6151
R2613 B.n499 B.n164 10.6151
R2614 B.n500 B.n499 10.6151
R2615 B.n501 B.n500 10.6151
R2616 B.n501 B.n162 10.6151
R2617 B.n505 B.n162 10.6151
R2618 B.n506 B.n505 10.6151
R2619 B.n507 B.n506 10.6151
R2620 B.n507 B.n160 10.6151
R2621 B.n511 B.n160 10.6151
R2622 B.n973 B.n0 8.11757
R2623 B.n973 B.n1 8.11757
R2624 B.n799 B.n798 6.5566
R2625 B.n786 B.n68 6.5566
R2626 B.n420 B.n419 6.5566
R2627 B.n435 B.n434 6.5566
R2628 B.n800 B.n799 4.05904
R2629 B.n783 B.n68 4.05904
R2630 B.n419 B.n418 4.05904
R2631 B.n434 B.n184 4.05904
R2632 VN.n72 VN.n71 161.3
R2633 VN.n70 VN.n38 161.3
R2634 VN.n69 VN.n68 161.3
R2635 VN.n67 VN.n39 161.3
R2636 VN.n66 VN.n65 161.3
R2637 VN.n64 VN.n40 161.3
R2638 VN.n63 VN.n62 161.3
R2639 VN.n61 VN.n41 161.3
R2640 VN.n60 VN.n59 161.3
R2641 VN.n58 VN.n42 161.3
R2642 VN.n57 VN.n56 161.3
R2643 VN.n55 VN.n44 161.3
R2644 VN.n54 VN.n53 161.3
R2645 VN.n52 VN.n45 161.3
R2646 VN.n51 VN.n50 161.3
R2647 VN.n49 VN.n46 161.3
R2648 VN.n35 VN.n34 161.3
R2649 VN.n33 VN.n1 161.3
R2650 VN.n32 VN.n31 161.3
R2651 VN.n30 VN.n2 161.3
R2652 VN.n29 VN.n28 161.3
R2653 VN.n27 VN.n3 161.3
R2654 VN.n26 VN.n25 161.3
R2655 VN.n24 VN.n4 161.3
R2656 VN.n23 VN.n22 161.3
R2657 VN.n20 VN.n5 161.3
R2658 VN.n19 VN.n18 161.3
R2659 VN.n17 VN.n6 161.3
R2660 VN.n16 VN.n15 161.3
R2661 VN.n14 VN.n7 161.3
R2662 VN.n13 VN.n12 161.3
R2663 VN.n11 VN.n8 161.3
R2664 VN.n48 VN.t0 132.018
R2665 VN.n10 VN.t5 132.018
R2666 VN.n9 VN.t6 99.3625
R2667 VN.n21 VN.t3 99.3625
R2668 VN.n0 VN.t4 99.3625
R2669 VN.n47 VN.t7 99.3625
R2670 VN.n43 VN.t2 99.3625
R2671 VN.n37 VN.t1 99.3625
R2672 VN.n36 VN.n0 84.5894
R2673 VN.n73 VN.n37 84.5894
R2674 VN.n10 VN.n9 64.6381
R2675 VN.n48 VN.n47 64.6381
R2676 VN VN.n73 57.7784
R2677 VN.n15 VN.n6 56.5617
R2678 VN.n53 VN.n44 56.5617
R2679 VN.n28 VN.n2 56.0773
R2680 VN.n65 VN.n39 56.0773
R2681 VN.n28 VN.n27 25.0767
R2682 VN.n65 VN.n64 25.0767
R2683 VN.n13 VN.n8 24.5923
R2684 VN.n14 VN.n13 24.5923
R2685 VN.n15 VN.n14 24.5923
R2686 VN.n19 VN.n6 24.5923
R2687 VN.n20 VN.n19 24.5923
R2688 VN.n22 VN.n20 24.5923
R2689 VN.n26 VN.n4 24.5923
R2690 VN.n27 VN.n26 24.5923
R2691 VN.n32 VN.n2 24.5923
R2692 VN.n33 VN.n32 24.5923
R2693 VN.n34 VN.n33 24.5923
R2694 VN.n53 VN.n52 24.5923
R2695 VN.n52 VN.n51 24.5923
R2696 VN.n51 VN.n46 24.5923
R2697 VN.n64 VN.n63 24.5923
R2698 VN.n63 VN.n41 24.5923
R2699 VN.n59 VN.n58 24.5923
R2700 VN.n58 VN.n57 24.5923
R2701 VN.n57 VN.n44 24.5923
R2702 VN.n71 VN.n70 24.5923
R2703 VN.n70 VN.n69 24.5923
R2704 VN.n69 VN.n39 24.5923
R2705 VN.n21 VN.n4 14.5097
R2706 VN.n43 VN.n41 14.5097
R2707 VN.n9 VN.n8 10.0832
R2708 VN.n22 VN.n21 10.0832
R2709 VN.n47 VN.n46 10.0832
R2710 VN.n59 VN.n43 10.0832
R2711 VN.n34 VN.n0 5.65662
R2712 VN.n71 VN.n37 5.65662
R2713 VN.n49 VN.n48 3.2858
R2714 VN.n11 VN.n10 3.2858
R2715 VN.n73 VN.n72 0.354861
R2716 VN.n36 VN.n35 0.354861
R2717 VN VN.n36 0.267071
R2718 VN.n72 VN.n38 0.189894
R2719 VN.n68 VN.n38 0.189894
R2720 VN.n68 VN.n67 0.189894
R2721 VN.n67 VN.n66 0.189894
R2722 VN.n66 VN.n40 0.189894
R2723 VN.n62 VN.n40 0.189894
R2724 VN.n62 VN.n61 0.189894
R2725 VN.n61 VN.n60 0.189894
R2726 VN.n60 VN.n42 0.189894
R2727 VN.n56 VN.n42 0.189894
R2728 VN.n56 VN.n55 0.189894
R2729 VN.n55 VN.n54 0.189894
R2730 VN.n54 VN.n45 0.189894
R2731 VN.n50 VN.n45 0.189894
R2732 VN.n50 VN.n49 0.189894
R2733 VN.n12 VN.n11 0.189894
R2734 VN.n12 VN.n7 0.189894
R2735 VN.n16 VN.n7 0.189894
R2736 VN.n17 VN.n16 0.189894
R2737 VN.n18 VN.n17 0.189894
R2738 VN.n18 VN.n5 0.189894
R2739 VN.n23 VN.n5 0.189894
R2740 VN.n24 VN.n23 0.189894
R2741 VN.n25 VN.n24 0.189894
R2742 VN.n25 VN.n3 0.189894
R2743 VN.n29 VN.n3 0.189894
R2744 VN.n30 VN.n29 0.189894
R2745 VN.n31 VN.n30 0.189894
R2746 VN.n31 VN.n1 0.189894
R2747 VN.n35 VN.n1 0.189894
R2748 VDD2.n2 VDD2.n1 74.7237
R2749 VDD2.n2 VDD2.n0 74.7237
R2750 VDD2 VDD2.n5 74.7208
R2751 VDD2.n4 VDD2.n3 73.0938
R2752 VDD2.n4 VDD2.n2 51.6075
R2753 VDD2.n5 VDD2.t0 2.20274
R2754 VDD2.n5 VDD2.t7 2.20274
R2755 VDD2.n3 VDD2.t6 2.20274
R2756 VDD2.n3 VDD2.t5 2.20274
R2757 VDD2.n1 VDD2.t4 2.20274
R2758 VDD2.n1 VDD2.t3 2.20274
R2759 VDD2.n0 VDD2.t2 2.20274
R2760 VDD2.n0 VDD2.t1 2.20274
R2761 VDD2 VDD2.n4 1.74403
C0 VDD1 VP 11.648f
C1 B VDD1 2.02293f
C2 VDD1 VDD2 2.28623f
C3 B VP 2.56242f
C4 VP VDD2 0.624391f
C5 B VDD2 2.14979f
C6 w_n4880_n3920# VTAIL 4.90464f
C7 w_n4880_n3920# VN 10.2447f
C8 VTAIL VN 11.7745f
C9 w_n4880_n3920# VDD1 2.34572f
C10 VTAIL VDD1 9.26129f
C11 VDD1 VN 0.153937f
C12 w_n4880_n3920# VP 10.8811f
C13 VTAIL VP 11.7886f
C14 VP VN 9.36758f
C15 w_n4880_n3920# B 12.3892f
C16 w_n4880_n3920# VDD2 2.50154f
C17 B VTAIL 6.33929f
C18 B VN 1.49034f
C19 VTAIL VDD2 9.322269f
C20 VN VDD2 11.1794f
C21 VDD2 VSUBS 2.46042f
C22 VDD1 VSUBS 3.27324f
C23 VTAIL VSUBS 1.632401f
C24 VN VSUBS 8.132481f
C25 VP VSUBS 4.690831f
C26 B VSUBS 6.329934f
C27 w_n4880_n3920# VSUBS 0.23465p
C28 VDD2.t2 VSUBS 0.375069f
C29 VDD2.t1 VSUBS 0.375069f
C30 VDD2.n0 VSUBS 3.07212f
C31 VDD2.t4 VSUBS 0.375069f
C32 VDD2.t3 VSUBS 0.375069f
C33 VDD2.n1 VSUBS 3.07212f
C34 VDD2.n2 VSUBS 5.83808f
C35 VDD2.t6 VSUBS 0.375069f
C36 VDD2.t5 VSUBS 0.375069f
C37 VDD2.n3 VSUBS 3.04738f
C38 VDD2.n4 VSUBS 4.83901f
C39 VDD2.t0 VSUBS 0.375069f
C40 VDD2.t7 VSUBS 0.375069f
C41 VDD2.n5 VSUBS 3.07206f
C42 VN.t4 VSUBS 3.32546f
C43 VN.n0 VSUBS 1.23935f
C44 VN.n1 VSUBS 0.022975f
C45 VN.n2 VSUBS 0.039063f
C46 VN.n3 VSUBS 0.022975f
C47 VN.n4 VSUBS 0.033982f
C48 VN.n5 VSUBS 0.022975f
C49 VN.n6 VSUBS 0.033398f
C50 VN.n7 VSUBS 0.022975f
C51 VN.n8 VSUBS 0.030196f
C52 VN.t6 VSUBS 3.32546f
C53 VN.n9 VSUBS 1.23232f
C54 VN.t5 VSUBS 3.65361f
C55 VN.n10 VSUBS 1.17611f
C56 VN.n11 VSUBS 0.287416f
C57 VN.n12 VSUBS 0.022975f
C58 VN.n13 VSUBS 0.042606f
C59 VN.n14 VSUBS 0.042606f
C60 VN.n15 VSUBS 0.033398f
C61 VN.n16 VSUBS 0.022975f
C62 VN.n17 VSUBS 0.022975f
C63 VN.n18 VSUBS 0.022975f
C64 VN.n19 VSUBS 0.042606f
C65 VN.n20 VSUBS 0.042606f
C66 VN.t3 VSUBS 3.32546f
C67 VN.n21 VSUBS 1.15513f
C68 VN.n22 VSUBS 0.030196f
C69 VN.n23 VSUBS 0.022975f
C70 VN.n24 VSUBS 0.022975f
C71 VN.n25 VSUBS 0.022975f
C72 VN.n26 VSUBS 0.042606f
C73 VN.n27 VSUBS 0.043004f
C74 VN.n28 VSUBS 0.027335f
C75 VN.n29 VSUBS 0.022975f
C76 VN.n30 VSUBS 0.022975f
C77 VN.n31 VSUBS 0.022975f
C78 VN.n32 VSUBS 0.042606f
C79 VN.n33 VSUBS 0.042606f
C80 VN.n34 VSUBS 0.02641f
C81 VN.n35 VSUBS 0.037076f
C82 VN.n36 VSUBS 0.06586f
C83 VN.t1 VSUBS 3.32546f
C84 VN.n37 VSUBS 1.23935f
C85 VN.n38 VSUBS 0.022975f
C86 VN.n39 VSUBS 0.039063f
C87 VN.n40 VSUBS 0.022975f
C88 VN.n41 VSUBS 0.033982f
C89 VN.n42 VSUBS 0.022975f
C90 VN.t2 VSUBS 3.32546f
C91 VN.n43 VSUBS 1.15513f
C92 VN.n44 VSUBS 0.033398f
C93 VN.n45 VSUBS 0.022975f
C94 VN.n46 VSUBS 0.030196f
C95 VN.t0 VSUBS 3.65361f
C96 VN.t7 VSUBS 3.32546f
C97 VN.n47 VSUBS 1.23232f
C98 VN.n48 VSUBS 1.17611f
C99 VN.n49 VSUBS 0.287416f
C100 VN.n50 VSUBS 0.022975f
C101 VN.n51 VSUBS 0.042606f
C102 VN.n52 VSUBS 0.042606f
C103 VN.n53 VSUBS 0.033398f
C104 VN.n54 VSUBS 0.022975f
C105 VN.n55 VSUBS 0.022975f
C106 VN.n56 VSUBS 0.022975f
C107 VN.n57 VSUBS 0.042606f
C108 VN.n58 VSUBS 0.042606f
C109 VN.n59 VSUBS 0.030196f
C110 VN.n60 VSUBS 0.022975f
C111 VN.n61 VSUBS 0.022975f
C112 VN.n62 VSUBS 0.022975f
C113 VN.n63 VSUBS 0.042606f
C114 VN.n64 VSUBS 0.043004f
C115 VN.n65 VSUBS 0.027335f
C116 VN.n66 VSUBS 0.022975f
C117 VN.n67 VSUBS 0.022975f
C118 VN.n68 VSUBS 0.022975f
C119 VN.n69 VSUBS 0.042606f
C120 VN.n70 VSUBS 0.042606f
C121 VN.n71 VSUBS 0.02641f
C122 VN.n72 VSUBS 0.037076f
C123 VN.n73 VSUBS 1.61138f
C124 B.n0 VSUBS 0.007058f
C125 B.n1 VSUBS 0.007058f
C126 B.n2 VSUBS 0.010439f
C127 B.n3 VSUBS 0.007999f
C128 B.n4 VSUBS 0.007999f
C129 B.n5 VSUBS 0.007999f
C130 B.n6 VSUBS 0.007999f
C131 B.n7 VSUBS 0.007999f
C132 B.n8 VSUBS 0.007999f
C133 B.n9 VSUBS 0.007999f
C134 B.n10 VSUBS 0.007999f
C135 B.n11 VSUBS 0.007999f
C136 B.n12 VSUBS 0.007999f
C137 B.n13 VSUBS 0.007999f
C138 B.n14 VSUBS 0.007999f
C139 B.n15 VSUBS 0.007999f
C140 B.n16 VSUBS 0.007999f
C141 B.n17 VSUBS 0.007999f
C142 B.n18 VSUBS 0.007999f
C143 B.n19 VSUBS 0.007999f
C144 B.n20 VSUBS 0.007999f
C145 B.n21 VSUBS 0.007999f
C146 B.n22 VSUBS 0.007999f
C147 B.n23 VSUBS 0.007999f
C148 B.n24 VSUBS 0.007999f
C149 B.n25 VSUBS 0.007999f
C150 B.n26 VSUBS 0.007999f
C151 B.n27 VSUBS 0.007999f
C152 B.n28 VSUBS 0.007999f
C153 B.n29 VSUBS 0.007999f
C154 B.n30 VSUBS 0.007999f
C155 B.n31 VSUBS 0.007999f
C156 B.n32 VSUBS 0.007999f
C157 B.n33 VSUBS 0.007999f
C158 B.n34 VSUBS 0.018675f
C159 B.n35 VSUBS 0.007999f
C160 B.n36 VSUBS 0.007999f
C161 B.n37 VSUBS 0.007999f
C162 B.n38 VSUBS 0.007999f
C163 B.n39 VSUBS 0.007999f
C164 B.n40 VSUBS 0.007999f
C165 B.n41 VSUBS 0.007999f
C166 B.n42 VSUBS 0.007999f
C167 B.n43 VSUBS 0.007999f
C168 B.n44 VSUBS 0.007999f
C169 B.n45 VSUBS 0.007999f
C170 B.n46 VSUBS 0.007999f
C171 B.n47 VSUBS 0.007999f
C172 B.n48 VSUBS 0.007999f
C173 B.n49 VSUBS 0.007999f
C174 B.n50 VSUBS 0.007999f
C175 B.n51 VSUBS 0.007999f
C176 B.n52 VSUBS 0.007999f
C177 B.n53 VSUBS 0.007999f
C178 B.n54 VSUBS 0.007999f
C179 B.n55 VSUBS 0.007999f
C180 B.n56 VSUBS 0.007999f
C181 B.n57 VSUBS 0.007999f
C182 B.n58 VSUBS 0.007999f
C183 B.n59 VSUBS 0.007999f
C184 B.t10 VSUBS 0.313079f
C185 B.t11 VSUBS 0.361975f
C186 B.t9 VSUBS 2.77396f
C187 B.n60 VSUBS 0.575776f
C188 B.n61 VSUBS 0.334535f
C189 B.n62 VSUBS 0.007999f
C190 B.n63 VSUBS 0.007999f
C191 B.n64 VSUBS 0.007999f
C192 B.n65 VSUBS 0.007999f
C193 B.t1 VSUBS 0.313083f
C194 B.t2 VSUBS 0.361978f
C195 B.t0 VSUBS 2.77396f
C196 B.n66 VSUBS 0.575773f
C197 B.n67 VSUBS 0.334531f
C198 B.n68 VSUBS 0.018534f
C199 B.n69 VSUBS 0.007999f
C200 B.n70 VSUBS 0.007999f
C201 B.n71 VSUBS 0.007999f
C202 B.n72 VSUBS 0.007999f
C203 B.n73 VSUBS 0.007999f
C204 B.n74 VSUBS 0.007999f
C205 B.n75 VSUBS 0.007999f
C206 B.n76 VSUBS 0.007999f
C207 B.n77 VSUBS 0.007999f
C208 B.n78 VSUBS 0.007999f
C209 B.n79 VSUBS 0.007999f
C210 B.n80 VSUBS 0.007999f
C211 B.n81 VSUBS 0.007999f
C212 B.n82 VSUBS 0.007999f
C213 B.n83 VSUBS 0.007999f
C214 B.n84 VSUBS 0.007999f
C215 B.n85 VSUBS 0.007999f
C216 B.n86 VSUBS 0.007999f
C217 B.n87 VSUBS 0.007999f
C218 B.n88 VSUBS 0.007999f
C219 B.n89 VSUBS 0.007999f
C220 B.n90 VSUBS 0.007999f
C221 B.n91 VSUBS 0.007999f
C222 B.n92 VSUBS 0.007999f
C223 B.n93 VSUBS 0.019675f
C224 B.n94 VSUBS 0.007999f
C225 B.n95 VSUBS 0.007999f
C226 B.n96 VSUBS 0.007999f
C227 B.n97 VSUBS 0.007999f
C228 B.n98 VSUBS 0.007999f
C229 B.n99 VSUBS 0.007999f
C230 B.n100 VSUBS 0.007999f
C231 B.n101 VSUBS 0.007999f
C232 B.n102 VSUBS 0.007999f
C233 B.n103 VSUBS 0.007999f
C234 B.n104 VSUBS 0.007999f
C235 B.n105 VSUBS 0.007999f
C236 B.n106 VSUBS 0.007999f
C237 B.n107 VSUBS 0.007999f
C238 B.n108 VSUBS 0.007999f
C239 B.n109 VSUBS 0.007999f
C240 B.n110 VSUBS 0.007999f
C241 B.n111 VSUBS 0.007999f
C242 B.n112 VSUBS 0.007999f
C243 B.n113 VSUBS 0.007999f
C244 B.n114 VSUBS 0.007999f
C245 B.n115 VSUBS 0.007999f
C246 B.n116 VSUBS 0.007999f
C247 B.n117 VSUBS 0.007999f
C248 B.n118 VSUBS 0.007999f
C249 B.n119 VSUBS 0.007999f
C250 B.n120 VSUBS 0.007999f
C251 B.n121 VSUBS 0.007999f
C252 B.n122 VSUBS 0.007999f
C253 B.n123 VSUBS 0.007999f
C254 B.n124 VSUBS 0.007999f
C255 B.n125 VSUBS 0.007999f
C256 B.n126 VSUBS 0.007999f
C257 B.n127 VSUBS 0.007999f
C258 B.n128 VSUBS 0.007999f
C259 B.n129 VSUBS 0.007999f
C260 B.n130 VSUBS 0.007999f
C261 B.n131 VSUBS 0.007999f
C262 B.n132 VSUBS 0.007999f
C263 B.n133 VSUBS 0.007999f
C264 B.n134 VSUBS 0.007999f
C265 B.n135 VSUBS 0.007999f
C266 B.n136 VSUBS 0.007999f
C267 B.n137 VSUBS 0.007999f
C268 B.n138 VSUBS 0.007999f
C269 B.n139 VSUBS 0.007999f
C270 B.n140 VSUBS 0.007999f
C271 B.n141 VSUBS 0.007999f
C272 B.n142 VSUBS 0.007999f
C273 B.n143 VSUBS 0.007999f
C274 B.n144 VSUBS 0.007999f
C275 B.n145 VSUBS 0.007999f
C276 B.n146 VSUBS 0.007999f
C277 B.n147 VSUBS 0.007999f
C278 B.n148 VSUBS 0.007999f
C279 B.n149 VSUBS 0.007999f
C280 B.n150 VSUBS 0.007999f
C281 B.n151 VSUBS 0.007999f
C282 B.n152 VSUBS 0.007999f
C283 B.n153 VSUBS 0.007999f
C284 B.n154 VSUBS 0.007999f
C285 B.n155 VSUBS 0.007999f
C286 B.n156 VSUBS 0.007999f
C287 B.n157 VSUBS 0.007999f
C288 B.n158 VSUBS 0.007999f
C289 B.n159 VSUBS 0.018675f
C290 B.n160 VSUBS 0.007999f
C291 B.n161 VSUBS 0.007999f
C292 B.n162 VSUBS 0.007999f
C293 B.n163 VSUBS 0.007999f
C294 B.n164 VSUBS 0.007999f
C295 B.n165 VSUBS 0.007999f
C296 B.n166 VSUBS 0.007999f
C297 B.n167 VSUBS 0.007999f
C298 B.n168 VSUBS 0.007999f
C299 B.n169 VSUBS 0.007999f
C300 B.n170 VSUBS 0.007999f
C301 B.n171 VSUBS 0.007999f
C302 B.n172 VSUBS 0.007999f
C303 B.n173 VSUBS 0.007999f
C304 B.n174 VSUBS 0.007999f
C305 B.n175 VSUBS 0.007999f
C306 B.n176 VSUBS 0.007999f
C307 B.n177 VSUBS 0.007999f
C308 B.n178 VSUBS 0.007999f
C309 B.n179 VSUBS 0.007999f
C310 B.n180 VSUBS 0.007999f
C311 B.n181 VSUBS 0.007999f
C312 B.n182 VSUBS 0.007999f
C313 B.n183 VSUBS 0.007999f
C314 B.n184 VSUBS 0.005529f
C315 B.n185 VSUBS 0.007999f
C316 B.n186 VSUBS 0.007999f
C317 B.n187 VSUBS 0.007999f
C318 B.n188 VSUBS 0.007999f
C319 B.n189 VSUBS 0.007999f
C320 B.t8 VSUBS 0.313079f
C321 B.t7 VSUBS 0.361975f
C322 B.t6 VSUBS 2.77396f
C323 B.n190 VSUBS 0.575776f
C324 B.n191 VSUBS 0.334535f
C325 B.n192 VSUBS 0.007999f
C326 B.n193 VSUBS 0.007999f
C327 B.n194 VSUBS 0.007999f
C328 B.n195 VSUBS 0.007999f
C329 B.n196 VSUBS 0.007999f
C330 B.n197 VSUBS 0.007999f
C331 B.n198 VSUBS 0.007999f
C332 B.n199 VSUBS 0.007999f
C333 B.n200 VSUBS 0.007999f
C334 B.n201 VSUBS 0.007999f
C335 B.n202 VSUBS 0.007999f
C336 B.n203 VSUBS 0.007999f
C337 B.n204 VSUBS 0.007999f
C338 B.n205 VSUBS 0.007999f
C339 B.n206 VSUBS 0.007999f
C340 B.n207 VSUBS 0.007999f
C341 B.n208 VSUBS 0.007999f
C342 B.n209 VSUBS 0.007999f
C343 B.n210 VSUBS 0.007999f
C344 B.n211 VSUBS 0.007999f
C345 B.n212 VSUBS 0.007999f
C346 B.n213 VSUBS 0.007999f
C347 B.n214 VSUBS 0.007999f
C348 B.n215 VSUBS 0.007999f
C349 B.n216 VSUBS 0.018675f
C350 B.n217 VSUBS 0.007999f
C351 B.n218 VSUBS 0.007999f
C352 B.n219 VSUBS 0.007999f
C353 B.n220 VSUBS 0.007999f
C354 B.n221 VSUBS 0.007999f
C355 B.n222 VSUBS 0.007999f
C356 B.n223 VSUBS 0.007999f
C357 B.n224 VSUBS 0.007999f
C358 B.n225 VSUBS 0.007999f
C359 B.n226 VSUBS 0.007999f
C360 B.n227 VSUBS 0.007999f
C361 B.n228 VSUBS 0.007999f
C362 B.n229 VSUBS 0.007999f
C363 B.n230 VSUBS 0.007999f
C364 B.n231 VSUBS 0.007999f
C365 B.n232 VSUBS 0.007999f
C366 B.n233 VSUBS 0.007999f
C367 B.n234 VSUBS 0.007999f
C368 B.n235 VSUBS 0.007999f
C369 B.n236 VSUBS 0.007999f
C370 B.n237 VSUBS 0.007999f
C371 B.n238 VSUBS 0.007999f
C372 B.n239 VSUBS 0.007999f
C373 B.n240 VSUBS 0.007999f
C374 B.n241 VSUBS 0.007999f
C375 B.n242 VSUBS 0.007999f
C376 B.n243 VSUBS 0.007999f
C377 B.n244 VSUBS 0.007999f
C378 B.n245 VSUBS 0.007999f
C379 B.n246 VSUBS 0.007999f
C380 B.n247 VSUBS 0.007999f
C381 B.n248 VSUBS 0.007999f
C382 B.n249 VSUBS 0.007999f
C383 B.n250 VSUBS 0.007999f
C384 B.n251 VSUBS 0.007999f
C385 B.n252 VSUBS 0.007999f
C386 B.n253 VSUBS 0.007999f
C387 B.n254 VSUBS 0.007999f
C388 B.n255 VSUBS 0.007999f
C389 B.n256 VSUBS 0.007999f
C390 B.n257 VSUBS 0.007999f
C391 B.n258 VSUBS 0.007999f
C392 B.n259 VSUBS 0.007999f
C393 B.n260 VSUBS 0.007999f
C394 B.n261 VSUBS 0.007999f
C395 B.n262 VSUBS 0.007999f
C396 B.n263 VSUBS 0.007999f
C397 B.n264 VSUBS 0.007999f
C398 B.n265 VSUBS 0.007999f
C399 B.n266 VSUBS 0.007999f
C400 B.n267 VSUBS 0.007999f
C401 B.n268 VSUBS 0.007999f
C402 B.n269 VSUBS 0.007999f
C403 B.n270 VSUBS 0.007999f
C404 B.n271 VSUBS 0.007999f
C405 B.n272 VSUBS 0.007999f
C406 B.n273 VSUBS 0.007999f
C407 B.n274 VSUBS 0.007999f
C408 B.n275 VSUBS 0.007999f
C409 B.n276 VSUBS 0.007999f
C410 B.n277 VSUBS 0.007999f
C411 B.n278 VSUBS 0.007999f
C412 B.n279 VSUBS 0.007999f
C413 B.n280 VSUBS 0.007999f
C414 B.n281 VSUBS 0.007999f
C415 B.n282 VSUBS 0.007999f
C416 B.n283 VSUBS 0.007999f
C417 B.n284 VSUBS 0.007999f
C418 B.n285 VSUBS 0.007999f
C419 B.n286 VSUBS 0.007999f
C420 B.n287 VSUBS 0.007999f
C421 B.n288 VSUBS 0.007999f
C422 B.n289 VSUBS 0.007999f
C423 B.n290 VSUBS 0.007999f
C424 B.n291 VSUBS 0.007999f
C425 B.n292 VSUBS 0.007999f
C426 B.n293 VSUBS 0.007999f
C427 B.n294 VSUBS 0.007999f
C428 B.n295 VSUBS 0.007999f
C429 B.n296 VSUBS 0.007999f
C430 B.n297 VSUBS 0.007999f
C431 B.n298 VSUBS 0.007999f
C432 B.n299 VSUBS 0.007999f
C433 B.n300 VSUBS 0.007999f
C434 B.n301 VSUBS 0.007999f
C435 B.n302 VSUBS 0.007999f
C436 B.n303 VSUBS 0.007999f
C437 B.n304 VSUBS 0.007999f
C438 B.n305 VSUBS 0.007999f
C439 B.n306 VSUBS 0.007999f
C440 B.n307 VSUBS 0.007999f
C441 B.n308 VSUBS 0.007999f
C442 B.n309 VSUBS 0.007999f
C443 B.n310 VSUBS 0.007999f
C444 B.n311 VSUBS 0.007999f
C445 B.n312 VSUBS 0.007999f
C446 B.n313 VSUBS 0.007999f
C447 B.n314 VSUBS 0.007999f
C448 B.n315 VSUBS 0.007999f
C449 B.n316 VSUBS 0.007999f
C450 B.n317 VSUBS 0.007999f
C451 B.n318 VSUBS 0.007999f
C452 B.n319 VSUBS 0.007999f
C453 B.n320 VSUBS 0.007999f
C454 B.n321 VSUBS 0.007999f
C455 B.n322 VSUBS 0.007999f
C456 B.n323 VSUBS 0.007999f
C457 B.n324 VSUBS 0.007999f
C458 B.n325 VSUBS 0.007999f
C459 B.n326 VSUBS 0.007999f
C460 B.n327 VSUBS 0.007999f
C461 B.n328 VSUBS 0.007999f
C462 B.n329 VSUBS 0.007999f
C463 B.n330 VSUBS 0.007999f
C464 B.n331 VSUBS 0.007999f
C465 B.n332 VSUBS 0.007999f
C466 B.n333 VSUBS 0.007999f
C467 B.n334 VSUBS 0.007999f
C468 B.n335 VSUBS 0.007999f
C469 B.n336 VSUBS 0.007999f
C470 B.n337 VSUBS 0.007999f
C471 B.n338 VSUBS 0.007999f
C472 B.n339 VSUBS 0.007999f
C473 B.n340 VSUBS 0.007999f
C474 B.n341 VSUBS 0.007999f
C475 B.n342 VSUBS 0.007999f
C476 B.n343 VSUBS 0.018675f
C477 B.n344 VSUBS 0.019675f
C478 B.n345 VSUBS 0.019675f
C479 B.n346 VSUBS 0.007999f
C480 B.n347 VSUBS 0.007999f
C481 B.n348 VSUBS 0.007999f
C482 B.n349 VSUBS 0.007999f
C483 B.n350 VSUBS 0.007999f
C484 B.n351 VSUBS 0.007999f
C485 B.n352 VSUBS 0.007999f
C486 B.n353 VSUBS 0.007999f
C487 B.n354 VSUBS 0.007999f
C488 B.n355 VSUBS 0.007999f
C489 B.n356 VSUBS 0.007999f
C490 B.n357 VSUBS 0.007999f
C491 B.n358 VSUBS 0.007999f
C492 B.n359 VSUBS 0.007999f
C493 B.n360 VSUBS 0.007999f
C494 B.n361 VSUBS 0.007999f
C495 B.n362 VSUBS 0.007999f
C496 B.n363 VSUBS 0.007999f
C497 B.n364 VSUBS 0.007999f
C498 B.n365 VSUBS 0.007999f
C499 B.n366 VSUBS 0.007999f
C500 B.n367 VSUBS 0.007999f
C501 B.n368 VSUBS 0.007999f
C502 B.n369 VSUBS 0.007999f
C503 B.n370 VSUBS 0.007999f
C504 B.n371 VSUBS 0.007999f
C505 B.n372 VSUBS 0.007999f
C506 B.n373 VSUBS 0.007999f
C507 B.n374 VSUBS 0.007999f
C508 B.n375 VSUBS 0.007999f
C509 B.n376 VSUBS 0.007999f
C510 B.n377 VSUBS 0.007999f
C511 B.n378 VSUBS 0.007999f
C512 B.n379 VSUBS 0.007999f
C513 B.n380 VSUBS 0.007999f
C514 B.n381 VSUBS 0.007999f
C515 B.n382 VSUBS 0.007999f
C516 B.n383 VSUBS 0.007999f
C517 B.n384 VSUBS 0.007999f
C518 B.n385 VSUBS 0.007999f
C519 B.n386 VSUBS 0.007999f
C520 B.n387 VSUBS 0.007999f
C521 B.n388 VSUBS 0.007999f
C522 B.n389 VSUBS 0.007999f
C523 B.n390 VSUBS 0.007999f
C524 B.n391 VSUBS 0.007999f
C525 B.n392 VSUBS 0.007999f
C526 B.n393 VSUBS 0.007999f
C527 B.n394 VSUBS 0.007999f
C528 B.n395 VSUBS 0.007999f
C529 B.n396 VSUBS 0.007999f
C530 B.n397 VSUBS 0.007999f
C531 B.n398 VSUBS 0.007999f
C532 B.n399 VSUBS 0.007999f
C533 B.n400 VSUBS 0.007999f
C534 B.n401 VSUBS 0.007999f
C535 B.n402 VSUBS 0.007999f
C536 B.n403 VSUBS 0.007999f
C537 B.n404 VSUBS 0.007999f
C538 B.n405 VSUBS 0.007999f
C539 B.n406 VSUBS 0.007999f
C540 B.n407 VSUBS 0.007999f
C541 B.n408 VSUBS 0.007999f
C542 B.n409 VSUBS 0.007999f
C543 B.n410 VSUBS 0.007999f
C544 B.n411 VSUBS 0.007999f
C545 B.n412 VSUBS 0.007999f
C546 B.n413 VSUBS 0.007999f
C547 B.n414 VSUBS 0.007999f
C548 B.n415 VSUBS 0.007999f
C549 B.n416 VSUBS 0.007999f
C550 B.n417 VSUBS 0.007999f
C551 B.n418 VSUBS 0.005529f
C552 B.n419 VSUBS 0.018534f
C553 B.n420 VSUBS 0.00647f
C554 B.n421 VSUBS 0.007999f
C555 B.n422 VSUBS 0.007999f
C556 B.n423 VSUBS 0.007999f
C557 B.n424 VSUBS 0.007999f
C558 B.n425 VSUBS 0.007999f
C559 B.n426 VSUBS 0.007999f
C560 B.n427 VSUBS 0.007999f
C561 B.n428 VSUBS 0.007999f
C562 B.n429 VSUBS 0.007999f
C563 B.n430 VSUBS 0.007999f
C564 B.n431 VSUBS 0.007999f
C565 B.t5 VSUBS 0.313083f
C566 B.t4 VSUBS 0.361978f
C567 B.t3 VSUBS 2.77396f
C568 B.n432 VSUBS 0.575773f
C569 B.n433 VSUBS 0.334531f
C570 B.n434 VSUBS 0.018534f
C571 B.n435 VSUBS 0.00647f
C572 B.n436 VSUBS 0.007999f
C573 B.n437 VSUBS 0.007999f
C574 B.n438 VSUBS 0.007999f
C575 B.n439 VSUBS 0.007999f
C576 B.n440 VSUBS 0.007999f
C577 B.n441 VSUBS 0.007999f
C578 B.n442 VSUBS 0.007999f
C579 B.n443 VSUBS 0.007999f
C580 B.n444 VSUBS 0.007999f
C581 B.n445 VSUBS 0.007999f
C582 B.n446 VSUBS 0.007999f
C583 B.n447 VSUBS 0.007999f
C584 B.n448 VSUBS 0.007999f
C585 B.n449 VSUBS 0.007999f
C586 B.n450 VSUBS 0.007999f
C587 B.n451 VSUBS 0.007999f
C588 B.n452 VSUBS 0.007999f
C589 B.n453 VSUBS 0.007999f
C590 B.n454 VSUBS 0.007999f
C591 B.n455 VSUBS 0.007999f
C592 B.n456 VSUBS 0.007999f
C593 B.n457 VSUBS 0.007999f
C594 B.n458 VSUBS 0.007999f
C595 B.n459 VSUBS 0.007999f
C596 B.n460 VSUBS 0.007999f
C597 B.n461 VSUBS 0.007999f
C598 B.n462 VSUBS 0.007999f
C599 B.n463 VSUBS 0.007999f
C600 B.n464 VSUBS 0.007999f
C601 B.n465 VSUBS 0.007999f
C602 B.n466 VSUBS 0.007999f
C603 B.n467 VSUBS 0.007999f
C604 B.n468 VSUBS 0.007999f
C605 B.n469 VSUBS 0.007999f
C606 B.n470 VSUBS 0.007999f
C607 B.n471 VSUBS 0.007999f
C608 B.n472 VSUBS 0.007999f
C609 B.n473 VSUBS 0.007999f
C610 B.n474 VSUBS 0.007999f
C611 B.n475 VSUBS 0.007999f
C612 B.n476 VSUBS 0.007999f
C613 B.n477 VSUBS 0.007999f
C614 B.n478 VSUBS 0.007999f
C615 B.n479 VSUBS 0.007999f
C616 B.n480 VSUBS 0.007999f
C617 B.n481 VSUBS 0.007999f
C618 B.n482 VSUBS 0.007999f
C619 B.n483 VSUBS 0.007999f
C620 B.n484 VSUBS 0.007999f
C621 B.n485 VSUBS 0.007999f
C622 B.n486 VSUBS 0.007999f
C623 B.n487 VSUBS 0.007999f
C624 B.n488 VSUBS 0.007999f
C625 B.n489 VSUBS 0.007999f
C626 B.n490 VSUBS 0.007999f
C627 B.n491 VSUBS 0.007999f
C628 B.n492 VSUBS 0.007999f
C629 B.n493 VSUBS 0.007999f
C630 B.n494 VSUBS 0.007999f
C631 B.n495 VSUBS 0.007999f
C632 B.n496 VSUBS 0.007999f
C633 B.n497 VSUBS 0.007999f
C634 B.n498 VSUBS 0.007999f
C635 B.n499 VSUBS 0.007999f
C636 B.n500 VSUBS 0.007999f
C637 B.n501 VSUBS 0.007999f
C638 B.n502 VSUBS 0.007999f
C639 B.n503 VSUBS 0.007999f
C640 B.n504 VSUBS 0.007999f
C641 B.n505 VSUBS 0.007999f
C642 B.n506 VSUBS 0.007999f
C643 B.n507 VSUBS 0.007999f
C644 B.n508 VSUBS 0.007999f
C645 B.n509 VSUBS 0.007999f
C646 B.n510 VSUBS 0.019675f
C647 B.n511 VSUBS 0.018764f
C648 B.n512 VSUBS 0.019586f
C649 B.n513 VSUBS 0.007999f
C650 B.n514 VSUBS 0.007999f
C651 B.n515 VSUBS 0.007999f
C652 B.n516 VSUBS 0.007999f
C653 B.n517 VSUBS 0.007999f
C654 B.n518 VSUBS 0.007999f
C655 B.n519 VSUBS 0.007999f
C656 B.n520 VSUBS 0.007999f
C657 B.n521 VSUBS 0.007999f
C658 B.n522 VSUBS 0.007999f
C659 B.n523 VSUBS 0.007999f
C660 B.n524 VSUBS 0.007999f
C661 B.n525 VSUBS 0.007999f
C662 B.n526 VSUBS 0.007999f
C663 B.n527 VSUBS 0.007999f
C664 B.n528 VSUBS 0.007999f
C665 B.n529 VSUBS 0.007999f
C666 B.n530 VSUBS 0.007999f
C667 B.n531 VSUBS 0.007999f
C668 B.n532 VSUBS 0.007999f
C669 B.n533 VSUBS 0.007999f
C670 B.n534 VSUBS 0.007999f
C671 B.n535 VSUBS 0.007999f
C672 B.n536 VSUBS 0.007999f
C673 B.n537 VSUBS 0.007999f
C674 B.n538 VSUBS 0.007999f
C675 B.n539 VSUBS 0.007999f
C676 B.n540 VSUBS 0.007999f
C677 B.n541 VSUBS 0.007999f
C678 B.n542 VSUBS 0.007999f
C679 B.n543 VSUBS 0.007999f
C680 B.n544 VSUBS 0.007999f
C681 B.n545 VSUBS 0.007999f
C682 B.n546 VSUBS 0.007999f
C683 B.n547 VSUBS 0.007999f
C684 B.n548 VSUBS 0.007999f
C685 B.n549 VSUBS 0.007999f
C686 B.n550 VSUBS 0.007999f
C687 B.n551 VSUBS 0.007999f
C688 B.n552 VSUBS 0.007999f
C689 B.n553 VSUBS 0.007999f
C690 B.n554 VSUBS 0.007999f
C691 B.n555 VSUBS 0.007999f
C692 B.n556 VSUBS 0.007999f
C693 B.n557 VSUBS 0.007999f
C694 B.n558 VSUBS 0.007999f
C695 B.n559 VSUBS 0.007999f
C696 B.n560 VSUBS 0.007999f
C697 B.n561 VSUBS 0.007999f
C698 B.n562 VSUBS 0.007999f
C699 B.n563 VSUBS 0.007999f
C700 B.n564 VSUBS 0.007999f
C701 B.n565 VSUBS 0.007999f
C702 B.n566 VSUBS 0.007999f
C703 B.n567 VSUBS 0.007999f
C704 B.n568 VSUBS 0.007999f
C705 B.n569 VSUBS 0.007999f
C706 B.n570 VSUBS 0.007999f
C707 B.n571 VSUBS 0.007999f
C708 B.n572 VSUBS 0.007999f
C709 B.n573 VSUBS 0.007999f
C710 B.n574 VSUBS 0.007999f
C711 B.n575 VSUBS 0.007999f
C712 B.n576 VSUBS 0.007999f
C713 B.n577 VSUBS 0.007999f
C714 B.n578 VSUBS 0.007999f
C715 B.n579 VSUBS 0.007999f
C716 B.n580 VSUBS 0.007999f
C717 B.n581 VSUBS 0.007999f
C718 B.n582 VSUBS 0.007999f
C719 B.n583 VSUBS 0.007999f
C720 B.n584 VSUBS 0.007999f
C721 B.n585 VSUBS 0.007999f
C722 B.n586 VSUBS 0.007999f
C723 B.n587 VSUBS 0.007999f
C724 B.n588 VSUBS 0.007999f
C725 B.n589 VSUBS 0.007999f
C726 B.n590 VSUBS 0.007999f
C727 B.n591 VSUBS 0.007999f
C728 B.n592 VSUBS 0.007999f
C729 B.n593 VSUBS 0.007999f
C730 B.n594 VSUBS 0.007999f
C731 B.n595 VSUBS 0.007999f
C732 B.n596 VSUBS 0.007999f
C733 B.n597 VSUBS 0.007999f
C734 B.n598 VSUBS 0.007999f
C735 B.n599 VSUBS 0.007999f
C736 B.n600 VSUBS 0.007999f
C737 B.n601 VSUBS 0.007999f
C738 B.n602 VSUBS 0.007999f
C739 B.n603 VSUBS 0.007999f
C740 B.n604 VSUBS 0.007999f
C741 B.n605 VSUBS 0.007999f
C742 B.n606 VSUBS 0.007999f
C743 B.n607 VSUBS 0.007999f
C744 B.n608 VSUBS 0.007999f
C745 B.n609 VSUBS 0.007999f
C746 B.n610 VSUBS 0.007999f
C747 B.n611 VSUBS 0.007999f
C748 B.n612 VSUBS 0.007999f
C749 B.n613 VSUBS 0.007999f
C750 B.n614 VSUBS 0.007999f
C751 B.n615 VSUBS 0.007999f
C752 B.n616 VSUBS 0.007999f
C753 B.n617 VSUBS 0.007999f
C754 B.n618 VSUBS 0.007999f
C755 B.n619 VSUBS 0.007999f
C756 B.n620 VSUBS 0.007999f
C757 B.n621 VSUBS 0.007999f
C758 B.n622 VSUBS 0.007999f
C759 B.n623 VSUBS 0.007999f
C760 B.n624 VSUBS 0.007999f
C761 B.n625 VSUBS 0.007999f
C762 B.n626 VSUBS 0.007999f
C763 B.n627 VSUBS 0.007999f
C764 B.n628 VSUBS 0.007999f
C765 B.n629 VSUBS 0.007999f
C766 B.n630 VSUBS 0.007999f
C767 B.n631 VSUBS 0.007999f
C768 B.n632 VSUBS 0.007999f
C769 B.n633 VSUBS 0.007999f
C770 B.n634 VSUBS 0.007999f
C771 B.n635 VSUBS 0.007999f
C772 B.n636 VSUBS 0.007999f
C773 B.n637 VSUBS 0.007999f
C774 B.n638 VSUBS 0.007999f
C775 B.n639 VSUBS 0.007999f
C776 B.n640 VSUBS 0.007999f
C777 B.n641 VSUBS 0.007999f
C778 B.n642 VSUBS 0.007999f
C779 B.n643 VSUBS 0.007999f
C780 B.n644 VSUBS 0.007999f
C781 B.n645 VSUBS 0.007999f
C782 B.n646 VSUBS 0.007999f
C783 B.n647 VSUBS 0.007999f
C784 B.n648 VSUBS 0.007999f
C785 B.n649 VSUBS 0.007999f
C786 B.n650 VSUBS 0.007999f
C787 B.n651 VSUBS 0.007999f
C788 B.n652 VSUBS 0.007999f
C789 B.n653 VSUBS 0.007999f
C790 B.n654 VSUBS 0.007999f
C791 B.n655 VSUBS 0.007999f
C792 B.n656 VSUBS 0.007999f
C793 B.n657 VSUBS 0.007999f
C794 B.n658 VSUBS 0.007999f
C795 B.n659 VSUBS 0.007999f
C796 B.n660 VSUBS 0.007999f
C797 B.n661 VSUBS 0.007999f
C798 B.n662 VSUBS 0.007999f
C799 B.n663 VSUBS 0.007999f
C800 B.n664 VSUBS 0.007999f
C801 B.n665 VSUBS 0.007999f
C802 B.n666 VSUBS 0.007999f
C803 B.n667 VSUBS 0.007999f
C804 B.n668 VSUBS 0.007999f
C805 B.n669 VSUBS 0.007999f
C806 B.n670 VSUBS 0.007999f
C807 B.n671 VSUBS 0.007999f
C808 B.n672 VSUBS 0.007999f
C809 B.n673 VSUBS 0.007999f
C810 B.n674 VSUBS 0.007999f
C811 B.n675 VSUBS 0.007999f
C812 B.n676 VSUBS 0.007999f
C813 B.n677 VSUBS 0.007999f
C814 B.n678 VSUBS 0.007999f
C815 B.n679 VSUBS 0.007999f
C816 B.n680 VSUBS 0.007999f
C817 B.n681 VSUBS 0.007999f
C818 B.n682 VSUBS 0.007999f
C819 B.n683 VSUBS 0.007999f
C820 B.n684 VSUBS 0.007999f
C821 B.n685 VSUBS 0.007999f
C822 B.n686 VSUBS 0.007999f
C823 B.n687 VSUBS 0.007999f
C824 B.n688 VSUBS 0.007999f
C825 B.n689 VSUBS 0.007999f
C826 B.n690 VSUBS 0.007999f
C827 B.n691 VSUBS 0.007999f
C828 B.n692 VSUBS 0.007999f
C829 B.n693 VSUBS 0.007999f
C830 B.n694 VSUBS 0.007999f
C831 B.n695 VSUBS 0.007999f
C832 B.n696 VSUBS 0.007999f
C833 B.n697 VSUBS 0.007999f
C834 B.n698 VSUBS 0.007999f
C835 B.n699 VSUBS 0.007999f
C836 B.n700 VSUBS 0.007999f
C837 B.n701 VSUBS 0.007999f
C838 B.n702 VSUBS 0.007999f
C839 B.n703 VSUBS 0.007999f
C840 B.n704 VSUBS 0.007999f
C841 B.n705 VSUBS 0.007999f
C842 B.n706 VSUBS 0.007999f
C843 B.n707 VSUBS 0.007999f
C844 B.n708 VSUBS 0.018675f
C845 B.n709 VSUBS 0.018675f
C846 B.n710 VSUBS 0.019675f
C847 B.n711 VSUBS 0.007999f
C848 B.n712 VSUBS 0.007999f
C849 B.n713 VSUBS 0.007999f
C850 B.n714 VSUBS 0.007999f
C851 B.n715 VSUBS 0.007999f
C852 B.n716 VSUBS 0.007999f
C853 B.n717 VSUBS 0.007999f
C854 B.n718 VSUBS 0.007999f
C855 B.n719 VSUBS 0.007999f
C856 B.n720 VSUBS 0.007999f
C857 B.n721 VSUBS 0.007999f
C858 B.n722 VSUBS 0.007999f
C859 B.n723 VSUBS 0.007999f
C860 B.n724 VSUBS 0.007999f
C861 B.n725 VSUBS 0.007999f
C862 B.n726 VSUBS 0.007999f
C863 B.n727 VSUBS 0.007999f
C864 B.n728 VSUBS 0.007999f
C865 B.n729 VSUBS 0.007999f
C866 B.n730 VSUBS 0.007999f
C867 B.n731 VSUBS 0.007999f
C868 B.n732 VSUBS 0.007999f
C869 B.n733 VSUBS 0.007999f
C870 B.n734 VSUBS 0.007999f
C871 B.n735 VSUBS 0.007999f
C872 B.n736 VSUBS 0.007999f
C873 B.n737 VSUBS 0.007999f
C874 B.n738 VSUBS 0.007999f
C875 B.n739 VSUBS 0.007999f
C876 B.n740 VSUBS 0.007999f
C877 B.n741 VSUBS 0.007999f
C878 B.n742 VSUBS 0.007999f
C879 B.n743 VSUBS 0.007999f
C880 B.n744 VSUBS 0.007999f
C881 B.n745 VSUBS 0.007999f
C882 B.n746 VSUBS 0.007999f
C883 B.n747 VSUBS 0.007999f
C884 B.n748 VSUBS 0.007999f
C885 B.n749 VSUBS 0.007999f
C886 B.n750 VSUBS 0.007999f
C887 B.n751 VSUBS 0.007999f
C888 B.n752 VSUBS 0.007999f
C889 B.n753 VSUBS 0.007999f
C890 B.n754 VSUBS 0.007999f
C891 B.n755 VSUBS 0.007999f
C892 B.n756 VSUBS 0.007999f
C893 B.n757 VSUBS 0.007999f
C894 B.n758 VSUBS 0.007999f
C895 B.n759 VSUBS 0.007999f
C896 B.n760 VSUBS 0.007999f
C897 B.n761 VSUBS 0.007999f
C898 B.n762 VSUBS 0.007999f
C899 B.n763 VSUBS 0.007999f
C900 B.n764 VSUBS 0.007999f
C901 B.n765 VSUBS 0.007999f
C902 B.n766 VSUBS 0.007999f
C903 B.n767 VSUBS 0.007999f
C904 B.n768 VSUBS 0.007999f
C905 B.n769 VSUBS 0.007999f
C906 B.n770 VSUBS 0.007999f
C907 B.n771 VSUBS 0.007999f
C908 B.n772 VSUBS 0.007999f
C909 B.n773 VSUBS 0.007999f
C910 B.n774 VSUBS 0.007999f
C911 B.n775 VSUBS 0.007999f
C912 B.n776 VSUBS 0.007999f
C913 B.n777 VSUBS 0.007999f
C914 B.n778 VSUBS 0.007999f
C915 B.n779 VSUBS 0.007999f
C916 B.n780 VSUBS 0.007999f
C917 B.n781 VSUBS 0.007999f
C918 B.n782 VSUBS 0.007999f
C919 B.n783 VSUBS 0.005529f
C920 B.n784 VSUBS 0.007999f
C921 B.n785 VSUBS 0.007999f
C922 B.n786 VSUBS 0.00647f
C923 B.n787 VSUBS 0.007999f
C924 B.n788 VSUBS 0.007999f
C925 B.n789 VSUBS 0.007999f
C926 B.n790 VSUBS 0.007999f
C927 B.n791 VSUBS 0.007999f
C928 B.n792 VSUBS 0.007999f
C929 B.n793 VSUBS 0.007999f
C930 B.n794 VSUBS 0.007999f
C931 B.n795 VSUBS 0.007999f
C932 B.n796 VSUBS 0.007999f
C933 B.n797 VSUBS 0.007999f
C934 B.n798 VSUBS 0.00647f
C935 B.n799 VSUBS 0.018534f
C936 B.n800 VSUBS 0.005529f
C937 B.n801 VSUBS 0.007999f
C938 B.n802 VSUBS 0.007999f
C939 B.n803 VSUBS 0.007999f
C940 B.n804 VSUBS 0.007999f
C941 B.n805 VSUBS 0.007999f
C942 B.n806 VSUBS 0.007999f
C943 B.n807 VSUBS 0.007999f
C944 B.n808 VSUBS 0.007999f
C945 B.n809 VSUBS 0.007999f
C946 B.n810 VSUBS 0.007999f
C947 B.n811 VSUBS 0.007999f
C948 B.n812 VSUBS 0.007999f
C949 B.n813 VSUBS 0.007999f
C950 B.n814 VSUBS 0.007999f
C951 B.n815 VSUBS 0.007999f
C952 B.n816 VSUBS 0.007999f
C953 B.n817 VSUBS 0.007999f
C954 B.n818 VSUBS 0.007999f
C955 B.n819 VSUBS 0.007999f
C956 B.n820 VSUBS 0.007999f
C957 B.n821 VSUBS 0.007999f
C958 B.n822 VSUBS 0.007999f
C959 B.n823 VSUBS 0.007999f
C960 B.n824 VSUBS 0.007999f
C961 B.n825 VSUBS 0.007999f
C962 B.n826 VSUBS 0.007999f
C963 B.n827 VSUBS 0.007999f
C964 B.n828 VSUBS 0.007999f
C965 B.n829 VSUBS 0.007999f
C966 B.n830 VSUBS 0.007999f
C967 B.n831 VSUBS 0.007999f
C968 B.n832 VSUBS 0.007999f
C969 B.n833 VSUBS 0.007999f
C970 B.n834 VSUBS 0.007999f
C971 B.n835 VSUBS 0.007999f
C972 B.n836 VSUBS 0.007999f
C973 B.n837 VSUBS 0.007999f
C974 B.n838 VSUBS 0.007999f
C975 B.n839 VSUBS 0.007999f
C976 B.n840 VSUBS 0.007999f
C977 B.n841 VSUBS 0.007999f
C978 B.n842 VSUBS 0.007999f
C979 B.n843 VSUBS 0.007999f
C980 B.n844 VSUBS 0.007999f
C981 B.n845 VSUBS 0.007999f
C982 B.n846 VSUBS 0.007999f
C983 B.n847 VSUBS 0.007999f
C984 B.n848 VSUBS 0.007999f
C985 B.n849 VSUBS 0.007999f
C986 B.n850 VSUBS 0.007999f
C987 B.n851 VSUBS 0.007999f
C988 B.n852 VSUBS 0.007999f
C989 B.n853 VSUBS 0.007999f
C990 B.n854 VSUBS 0.007999f
C991 B.n855 VSUBS 0.007999f
C992 B.n856 VSUBS 0.007999f
C993 B.n857 VSUBS 0.007999f
C994 B.n858 VSUBS 0.007999f
C995 B.n859 VSUBS 0.007999f
C996 B.n860 VSUBS 0.007999f
C997 B.n861 VSUBS 0.007999f
C998 B.n862 VSUBS 0.007999f
C999 B.n863 VSUBS 0.007999f
C1000 B.n864 VSUBS 0.007999f
C1001 B.n865 VSUBS 0.007999f
C1002 B.n866 VSUBS 0.007999f
C1003 B.n867 VSUBS 0.007999f
C1004 B.n868 VSUBS 0.007999f
C1005 B.n869 VSUBS 0.007999f
C1006 B.n870 VSUBS 0.007999f
C1007 B.n871 VSUBS 0.007999f
C1008 B.n872 VSUBS 0.007999f
C1009 B.n873 VSUBS 0.019675f
C1010 B.n874 VSUBS 0.019675f
C1011 B.n875 VSUBS 0.018675f
C1012 B.n876 VSUBS 0.007999f
C1013 B.n877 VSUBS 0.007999f
C1014 B.n878 VSUBS 0.007999f
C1015 B.n879 VSUBS 0.007999f
C1016 B.n880 VSUBS 0.007999f
C1017 B.n881 VSUBS 0.007999f
C1018 B.n882 VSUBS 0.007999f
C1019 B.n883 VSUBS 0.007999f
C1020 B.n884 VSUBS 0.007999f
C1021 B.n885 VSUBS 0.007999f
C1022 B.n886 VSUBS 0.007999f
C1023 B.n887 VSUBS 0.007999f
C1024 B.n888 VSUBS 0.007999f
C1025 B.n889 VSUBS 0.007999f
C1026 B.n890 VSUBS 0.007999f
C1027 B.n891 VSUBS 0.007999f
C1028 B.n892 VSUBS 0.007999f
C1029 B.n893 VSUBS 0.007999f
C1030 B.n894 VSUBS 0.007999f
C1031 B.n895 VSUBS 0.007999f
C1032 B.n896 VSUBS 0.007999f
C1033 B.n897 VSUBS 0.007999f
C1034 B.n898 VSUBS 0.007999f
C1035 B.n899 VSUBS 0.007999f
C1036 B.n900 VSUBS 0.007999f
C1037 B.n901 VSUBS 0.007999f
C1038 B.n902 VSUBS 0.007999f
C1039 B.n903 VSUBS 0.007999f
C1040 B.n904 VSUBS 0.007999f
C1041 B.n905 VSUBS 0.007999f
C1042 B.n906 VSUBS 0.007999f
C1043 B.n907 VSUBS 0.007999f
C1044 B.n908 VSUBS 0.007999f
C1045 B.n909 VSUBS 0.007999f
C1046 B.n910 VSUBS 0.007999f
C1047 B.n911 VSUBS 0.007999f
C1048 B.n912 VSUBS 0.007999f
C1049 B.n913 VSUBS 0.007999f
C1050 B.n914 VSUBS 0.007999f
C1051 B.n915 VSUBS 0.007999f
C1052 B.n916 VSUBS 0.007999f
C1053 B.n917 VSUBS 0.007999f
C1054 B.n918 VSUBS 0.007999f
C1055 B.n919 VSUBS 0.007999f
C1056 B.n920 VSUBS 0.007999f
C1057 B.n921 VSUBS 0.007999f
C1058 B.n922 VSUBS 0.007999f
C1059 B.n923 VSUBS 0.007999f
C1060 B.n924 VSUBS 0.007999f
C1061 B.n925 VSUBS 0.007999f
C1062 B.n926 VSUBS 0.007999f
C1063 B.n927 VSUBS 0.007999f
C1064 B.n928 VSUBS 0.007999f
C1065 B.n929 VSUBS 0.007999f
C1066 B.n930 VSUBS 0.007999f
C1067 B.n931 VSUBS 0.007999f
C1068 B.n932 VSUBS 0.007999f
C1069 B.n933 VSUBS 0.007999f
C1070 B.n934 VSUBS 0.007999f
C1071 B.n935 VSUBS 0.007999f
C1072 B.n936 VSUBS 0.007999f
C1073 B.n937 VSUBS 0.007999f
C1074 B.n938 VSUBS 0.007999f
C1075 B.n939 VSUBS 0.007999f
C1076 B.n940 VSUBS 0.007999f
C1077 B.n941 VSUBS 0.007999f
C1078 B.n942 VSUBS 0.007999f
C1079 B.n943 VSUBS 0.007999f
C1080 B.n944 VSUBS 0.007999f
C1081 B.n945 VSUBS 0.007999f
C1082 B.n946 VSUBS 0.007999f
C1083 B.n947 VSUBS 0.007999f
C1084 B.n948 VSUBS 0.007999f
C1085 B.n949 VSUBS 0.007999f
C1086 B.n950 VSUBS 0.007999f
C1087 B.n951 VSUBS 0.007999f
C1088 B.n952 VSUBS 0.007999f
C1089 B.n953 VSUBS 0.007999f
C1090 B.n954 VSUBS 0.007999f
C1091 B.n955 VSUBS 0.007999f
C1092 B.n956 VSUBS 0.007999f
C1093 B.n957 VSUBS 0.007999f
C1094 B.n958 VSUBS 0.007999f
C1095 B.n959 VSUBS 0.007999f
C1096 B.n960 VSUBS 0.007999f
C1097 B.n961 VSUBS 0.007999f
C1098 B.n962 VSUBS 0.007999f
C1099 B.n963 VSUBS 0.007999f
C1100 B.n964 VSUBS 0.007999f
C1101 B.n965 VSUBS 0.007999f
C1102 B.n966 VSUBS 0.007999f
C1103 B.n967 VSUBS 0.007999f
C1104 B.n968 VSUBS 0.007999f
C1105 B.n969 VSUBS 0.007999f
C1106 B.n970 VSUBS 0.007999f
C1107 B.n971 VSUBS 0.010439f
C1108 B.n972 VSUBS 0.01112f
C1109 B.n973 VSUBS 0.022113f
C1110 VTAIL.t6 VSUBS 0.291674f
C1111 VTAIL.t2 VSUBS 0.291674f
C1112 VTAIL.n0 VSUBS 2.23249f
C1113 VTAIL.n1 VSUBS 0.848758f
C1114 VTAIL.n2 VSUBS 0.026524f
C1115 VTAIL.n3 VSUBS 0.025007f
C1116 VTAIL.n4 VSUBS 0.013438f
C1117 VTAIL.n5 VSUBS 0.031761f
C1118 VTAIL.n6 VSUBS 0.014228f
C1119 VTAIL.n7 VSUBS 0.025007f
C1120 VTAIL.n8 VSUBS 0.013438f
C1121 VTAIL.n9 VSUBS 0.031761f
C1122 VTAIL.n10 VSUBS 0.014228f
C1123 VTAIL.n11 VSUBS 0.025007f
C1124 VTAIL.n12 VSUBS 0.013438f
C1125 VTAIL.n13 VSUBS 0.031761f
C1126 VTAIL.n14 VSUBS 0.014228f
C1127 VTAIL.n15 VSUBS 0.025007f
C1128 VTAIL.n16 VSUBS 0.013438f
C1129 VTAIL.n17 VSUBS 0.031761f
C1130 VTAIL.n18 VSUBS 0.014228f
C1131 VTAIL.n19 VSUBS 0.025007f
C1132 VTAIL.n20 VSUBS 0.013438f
C1133 VTAIL.n21 VSUBS 0.031761f
C1134 VTAIL.n22 VSUBS 0.014228f
C1135 VTAIL.n23 VSUBS 0.025007f
C1136 VTAIL.n24 VSUBS 0.013438f
C1137 VTAIL.n25 VSUBS 0.031761f
C1138 VTAIL.n26 VSUBS 0.014228f
C1139 VTAIL.n27 VSUBS 0.174506f
C1140 VTAIL.t1 VSUBS 0.06798f
C1141 VTAIL.n28 VSUBS 0.023821f
C1142 VTAIL.n29 VSUBS 0.020205f
C1143 VTAIL.n30 VSUBS 0.013438f
C1144 VTAIL.n31 VSUBS 1.56949f
C1145 VTAIL.n32 VSUBS 0.025007f
C1146 VTAIL.n33 VSUBS 0.013438f
C1147 VTAIL.n34 VSUBS 0.014228f
C1148 VTAIL.n35 VSUBS 0.031761f
C1149 VTAIL.n36 VSUBS 0.031761f
C1150 VTAIL.n37 VSUBS 0.014228f
C1151 VTAIL.n38 VSUBS 0.013438f
C1152 VTAIL.n39 VSUBS 0.025007f
C1153 VTAIL.n40 VSUBS 0.025007f
C1154 VTAIL.n41 VSUBS 0.013438f
C1155 VTAIL.n42 VSUBS 0.014228f
C1156 VTAIL.n43 VSUBS 0.031761f
C1157 VTAIL.n44 VSUBS 0.031761f
C1158 VTAIL.n45 VSUBS 0.014228f
C1159 VTAIL.n46 VSUBS 0.013438f
C1160 VTAIL.n47 VSUBS 0.025007f
C1161 VTAIL.n48 VSUBS 0.025007f
C1162 VTAIL.n49 VSUBS 0.013438f
C1163 VTAIL.n50 VSUBS 0.014228f
C1164 VTAIL.n51 VSUBS 0.031761f
C1165 VTAIL.n52 VSUBS 0.031761f
C1166 VTAIL.n53 VSUBS 0.014228f
C1167 VTAIL.n54 VSUBS 0.013438f
C1168 VTAIL.n55 VSUBS 0.025007f
C1169 VTAIL.n56 VSUBS 0.025007f
C1170 VTAIL.n57 VSUBS 0.013438f
C1171 VTAIL.n58 VSUBS 0.014228f
C1172 VTAIL.n59 VSUBS 0.031761f
C1173 VTAIL.n60 VSUBS 0.031761f
C1174 VTAIL.n61 VSUBS 0.014228f
C1175 VTAIL.n62 VSUBS 0.013438f
C1176 VTAIL.n63 VSUBS 0.025007f
C1177 VTAIL.n64 VSUBS 0.025007f
C1178 VTAIL.n65 VSUBS 0.013438f
C1179 VTAIL.n66 VSUBS 0.014228f
C1180 VTAIL.n67 VSUBS 0.031761f
C1181 VTAIL.n68 VSUBS 0.031761f
C1182 VTAIL.n69 VSUBS 0.031761f
C1183 VTAIL.n70 VSUBS 0.014228f
C1184 VTAIL.n71 VSUBS 0.013438f
C1185 VTAIL.n72 VSUBS 0.025007f
C1186 VTAIL.n73 VSUBS 0.025007f
C1187 VTAIL.n74 VSUBS 0.013438f
C1188 VTAIL.n75 VSUBS 0.013833f
C1189 VTAIL.n76 VSUBS 0.013833f
C1190 VTAIL.n77 VSUBS 0.031761f
C1191 VTAIL.n78 VSUBS 0.073646f
C1192 VTAIL.n79 VSUBS 0.014228f
C1193 VTAIL.n80 VSUBS 0.013438f
C1194 VTAIL.n81 VSUBS 0.061901f
C1195 VTAIL.n82 VSUBS 0.037014f
C1196 VTAIL.n83 VSUBS 0.333134f
C1197 VTAIL.n84 VSUBS 0.026524f
C1198 VTAIL.n85 VSUBS 0.025007f
C1199 VTAIL.n86 VSUBS 0.013438f
C1200 VTAIL.n87 VSUBS 0.031761f
C1201 VTAIL.n88 VSUBS 0.014228f
C1202 VTAIL.n89 VSUBS 0.025007f
C1203 VTAIL.n90 VSUBS 0.013438f
C1204 VTAIL.n91 VSUBS 0.031761f
C1205 VTAIL.n92 VSUBS 0.014228f
C1206 VTAIL.n93 VSUBS 0.025007f
C1207 VTAIL.n94 VSUBS 0.013438f
C1208 VTAIL.n95 VSUBS 0.031761f
C1209 VTAIL.n96 VSUBS 0.014228f
C1210 VTAIL.n97 VSUBS 0.025007f
C1211 VTAIL.n98 VSUBS 0.013438f
C1212 VTAIL.n99 VSUBS 0.031761f
C1213 VTAIL.n100 VSUBS 0.014228f
C1214 VTAIL.n101 VSUBS 0.025007f
C1215 VTAIL.n102 VSUBS 0.013438f
C1216 VTAIL.n103 VSUBS 0.031761f
C1217 VTAIL.n104 VSUBS 0.014228f
C1218 VTAIL.n105 VSUBS 0.025007f
C1219 VTAIL.n106 VSUBS 0.013438f
C1220 VTAIL.n107 VSUBS 0.031761f
C1221 VTAIL.n108 VSUBS 0.014228f
C1222 VTAIL.n109 VSUBS 0.174506f
C1223 VTAIL.t14 VSUBS 0.06798f
C1224 VTAIL.n110 VSUBS 0.023821f
C1225 VTAIL.n111 VSUBS 0.020205f
C1226 VTAIL.n112 VSUBS 0.013438f
C1227 VTAIL.n113 VSUBS 1.56949f
C1228 VTAIL.n114 VSUBS 0.025007f
C1229 VTAIL.n115 VSUBS 0.013438f
C1230 VTAIL.n116 VSUBS 0.014228f
C1231 VTAIL.n117 VSUBS 0.031761f
C1232 VTAIL.n118 VSUBS 0.031761f
C1233 VTAIL.n119 VSUBS 0.014228f
C1234 VTAIL.n120 VSUBS 0.013438f
C1235 VTAIL.n121 VSUBS 0.025007f
C1236 VTAIL.n122 VSUBS 0.025007f
C1237 VTAIL.n123 VSUBS 0.013438f
C1238 VTAIL.n124 VSUBS 0.014228f
C1239 VTAIL.n125 VSUBS 0.031761f
C1240 VTAIL.n126 VSUBS 0.031761f
C1241 VTAIL.n127 VSUBS 0.014228f
C1242 VTAIL.n128 VSUBS 0.013438f
C1243 VTAIL.n129 VSUBS 0.025007f
C1244 VTAIL.n130 VSUBS 0.025007f
C1245 VTAIL.n131 VSUBS 0.013438f
C1246 VTAIL.n132 VSUBS 0.014228f
C1247 VTAIL.n133 VSUBS 0.031761f
C1248 VTAIL.n134 VSUBS 0.031761f
C1249 VTAIL.n135 VSUBS 0.014228f
C1250 VTAIL.n136 VSUBS 0.013438f
C1251 VTAIL.n137 VSUBS 0.025007f
C1252 VTAIL.n138 VSUBS 0.025007f
C1253 VTAIL.n139 VSUBS 0.013438f
C1254 VTAIL.n140 VSUBS 0.014228f
C1255 VTAIL.n141 VSUBS 0.031761f
C1256 VTAIL.n142 VSUBS 0.031761f
C1257 VTAIL.n143 VSUBS 0.014228f
C1258 VTAIL.n144 VSUBS 0.013438f
C1259 VTAIL.n145 VSUBS 0.025007f
C1260 VTAIL.n146 VSUBS 0.025007f
C1261 VTAIL.n147 VSUBS 0.013438f
C1262 VTAIL.n148 VSUBS 0.014228f
C1263 VTAIL.n149 VSUBS 0.031761f
C1264 VTAIL.n150 VSUBS 0.031761f
C1265 VTAIL.n151 VSUBS 0.031761f
C1266 VTAIL.n152 VSUBS 0.014228f
C1267 VTAIL.n153 VSUBS 0.013438f
C1268 VTAIL.n154 VSUBS 0.025007f
C1269 VTAIL.n155 VSUBS 0.025007f
C1270 VTAIL.n156 VSUBS 0.013438f
C1271 VTAIL.n157 VSUBS 0.013833f
C1272 VTAIL.n158 VSUBS 0.013833f
C1273 VTAIL.n159 VSUBS 0.031761f
C1274 VTAIL.n160 VSUBS 0.073646f
C1275 VTAIL.n161 VSUBS 0.014228f
C1276 VTAIL.n162 VSUBS 0.013438f
C1277 VTAIL.n163 VSUBS 0.061901f
C1278 VTAIL.n164 VSUBS 0.037014f
C1279 VTAIL.n165 VSUBS 0.333134f
C1280 VTAIL.t13 VSUBS 0.291674f
C1281 VTAIL.t12 VSUBS 0.291674f
C1282 VTAIL.n166 VSUBS 2.23249f
C1283 VTAIL.n167 VSUBS 1.11567f
C1284 VTAIL.n168 VSUBS 0.026524f
C1285 VTAIL.n169 VSUBS 0.025007f
C1286 VTAIL.n170 VSUBS 0.013438f
C1287 VTAIL.n171 VSUBS 0.031761f
C1288 VTAIL.n172 VSUBS 0.014228f
C1289 VTAIL.n173 VSUBS 0.025007f
C1290 VTAIL.n174 VSUBS 0.013438f
C1291 VTAIL.n175 VSUBS 0.031761f
C1292 VTAIL.n176 VSUBS 0.014228f
C1293 VTAIL.n177 VSUBS 0.025007f
C1294 VTAIL.n178 VSUBS 0.013438f
C1295 VTAIL.n179 VSUBS 0.031761f
C1296 VTAIL.n180 VSUBS 0.014228f
C1297 VTAIL.n181 VSUBS 0.025007f
C1298 VTAIL.n182 VSUBS 0.013438f
C1299 VTAIL.n183 VSUBS 0.031761f
C1300 VTAIL.n184 VSUBS 0.014228f
C1301 VTAIL.n185 VSUBS 0.025007f
C1302 VTAIL.n186 VSUBS 0.013438f
C1303 VTAIL.n187 VSUBS 0.031761f
C1304 VTAIL.n188 VSUBS 0.014228f
C1305 VTAIL.n189 VSUBS 0.025007f
C1306 VTAIL.n190 VSUBS 0.013438f
C1307 VTAIL.n191 VSUBS 0.031761f
C1308 VTAIL.n192 VSUBS 0.014228f
C1309 VTAIL.n193 VSUBS 0.174506f
C1310 VTAIL.t8 VSUBS 0.06798f
C1311 VTAIL.n194 VSUBS 0.023821f
C1312 VTAIL.n195 VSUBS 0.020205f
C1313 VTAIL.n196 VSUBS 0.013438f
C1314 VTAIL.n197 VSUBS 1.56949f
C1315 VTAIL.n198 VSUBS 0.025007f
C1316 VTAIL.n199 VSUBS 0.013438f
C1317 VTAIL.n200 VSUBS 0.014228f
C1318 VTAIL.n201 VSUBS 0.031761f
C1319 VTAIL.n202 VSUBS 0.031761f
C1320 VTAIL.n203 VSUBS 0.014228f
C1321 VTAIL.n204 VSUBS 0.013438f
C1322 VTAIL.n205 VSUBS 0.025007f
C1323 VTAIL.n206 VSUBS 0.025007f
C1324 VTAIL.n207 VSUBS 0.013438f
C1325 VTAIL.n208 VSUBS 0.014228f
C1326 VTAIL.n209 VSUBS 0.031761f
C1327 VTAIL.n210 VSUBS 0.031761f
C1328 VTAIL.n211 VSUBS 0.014228f
C1329 VTAIL.n212 VSUBS 0.013438f
C1330 VTAIL.n213 VSUBS 0.025007f
C1331 VTAIL.n214 VSUBS 0.025007f
C1332 VTAIL.n215 VSUBS 0.013438f
C1333 VTAIL.n216 VSUBS 0.014228f
C1334 VTAIL.n217 VSUBS 0.031761f
C1335 VTAIL.n218 VSUBS 0.031761f
C1336 VTAIL.n219 VSUBS 0.014228f
C1337 VTAIL.n220 VSUBS 0.013438f
C1338 VTAIL.n221 VSUBS 0.025007f
C1339 VTAIL.n222 VSUBS 0.025007f
C1340 VTAIL.n223 VSUBS 0.013438f
C1341 VTAIL.n224 VSUBS 0.014228f
C1342 VTAIL.n225 VSUBS 0.031761f
C1343 VTAIL.n226 VSUBS 0.031761f
C1344 VTAIL.n227 VSUBS 0.014228f
C1345 VTAIL.n228 VSUBS 0.013438f
C1346 VTAIL.n229 VSUBS 0.025007f
C1347 VTAIL.n230 VSUBS 0.025007f
C1348 VTAIL.n231 VSUBS 0.013438f
C1349 VTAIL.n232 VSUBS 0.014228f
C1350 VTAIL.n233 VSUBS 0.031761f
C1351 VTAIL.n234 VSUBS 0.031761f
C1352 VTAIL.n235 VSUBS 0.031761f
C1353 VTAIL.n236 VSUBS 0.014228f
C1354 VTAIL.n237 VSUBS 0.013438f
C1355 VTAIL.n238 VSUBS 0.025007f
C1356 VTAIL.n239 VSUBS 0.025007f
C1357 VTAIL.n240 VSUBS 0.013438f
C1358 VTAIL.n241 VSUBS 0.013833f
C1359 VTAIL.n242 VSUBS 0.013833f
C1360 VTAIL.n243 VSUBS 0.031761f
C1361 VTAIL.n244 VSUBS 0.073646f
C1362 VTAIL.n245 VSUBS 0.014228f
C1363 VTAIL.n246 VSUBS 0.013438f
C1364 VTAIL.n247 VSUBS 0.061901f
C1365 VTAIL.n248 VSUBS 0.037014f
C1366 VTAIL.n249 VSUBS 1.93184f
C1367 VTAIL.n250 VSUBS 0.026524f
C1368 VTAIL.n251 VSUBS 0.025007f
C1369 VTAIL.n252 VSUBS 0.013438f
C1370 VTAIL.n253 VSUBS 0.031761f
C1371 VTAIL.n254 VSUBS 0.014228f
C1372 VTAIL.n255 VSUBS 0.025007f
C1373 VTAIL.n256 VSUBS 0.013438f
C1374 VTAIL.n257 VSUBS 0.031761f
C1375 VTAIL.n258 VSUBS 0.031761f
C1376 VTAIL.n259 VSUBS 0.014228f
C1377 VTAIL.n260 VSUBS 0.025007f
C1378 VTAIL.n261 VSUBS 0.013438f
C1379 VTAIL.n262 VSUBS 0.031761f
C1380 VTAIL.n263 VSUBS 0.014228f
C1381 VTAIL.n264 VSUBS 0.025007f
C1382 VTAIL.n265 VSUBS 0.013438f
C1383 VTAIL.n266 VSUBS 0.031761f
C1384 VTAIL.n267 VSUBS 0.014228f
C1385 VTAIL.n268 VSUBS 0.025007f
C1386 VTAIL.n269 VSUBS 0.013438f
C1387 VTAIL.n270 VSUBS 0.031761f
C1388 VTAIL.n271 VSUBS 0.014228f
C1389 VTAIL.n272 VSUBS 0.025007f
C1390 VTAIL.n273 VSUBS 0.013438f
C1391 VTAIL.n274 VSUBS 0.031761f
C1392 VTAIL.n275 VSUBS 0.014228f
C1393 VTAIL.n276 VSUBS 0.174506f
C1394 VTAIL.t4 VSUBS 0.06798f
C1395 VTAIL.n277 VSUBS 0.023821f
C1396 VTAIL.n278 VSUBS 0.020205f
C1397 VTAIL.n279 VSUBS 0.013438f
C1398 VTAIL.n280 VSUBS 1.56949f
C1399 VTAIL.n281 VSUBS 0.025007f
C1400 VTAIL.n282 VSUBS 0.013438f
C1401 VTAIL.n283 VSUBS 0.014228f
C1402 VTAIL.n284 VSUBS 0.031761f
C1403 VTAIL.n285 VSUBS 0.031761f
C1404 VTAIL.n286 VSUBS 0.014228f
C1405 VTAIL.n287 VSUBS 0.013438f
C1406 VTAIL.n288 VSUBS 0.025007f
C1407 VTAIL.n289 VSUBS 0.025007f
C1408 VTAIL.n290 VSUBS 0.013438f
C1409 VTAIL.n291 VSUBS 0.014228f
C1410 VTAIL.n292 VSUBS 0.031761f
C1411 VTAIL.n293 VSUBS 0.031761f
C1412 VTAIL.n294 VSUBS 0.014228f
C1413 VTAIL.n295 VSUBS 0.013438f
C1414 VTAIL.n296 VSUBS 0.025007f
C1415 VTAIL.n297 VSUBS 0.025007f
C1416 VTAIL.n298 VSUBS 0.013438f
C1417 VTAIL.n299 VSUBS 0.014228f
C1418 VTAIL.n300 VSUBS 0.031761f
C1419 VTAIL.n301 VSUBS 0.031761f
C1420 VTAIL.n302 VSUBS 0.014228f
C1421 VTAIL.n303 VSUBS 0.013438f
C1422 VTAIL.n304 VSUBS 0.025007f
C1423 VTAIL.n305 VSUBS 0.025007f
C1424 VTAIL.n306 VSUBS 0.013438f
C1425 VTAIL.n307 VSUBS 0.014228f
C1426 VTAIL.n308 VSUBS 0.031761f
C1427 VTAIL.n309 VSUBS 0.031761f
C1428 VTAIL.n310 VSUBS 0.014228f
C1429 VTAIL.n311 VSUBS 0.013438f
C1430 VTAIL.n312 VSUBS 0.025007f
C1431 VTAIL.n313 VSUBS 0.025007f
C1432 VTAIL.n314 VSUBS 0.013438f
C1433 VTAIL.n315 VSUBS 0.014228f
C1434 VTAIL.n316 VSUBS 0.031761f
C1435 VTAIL.n317 VSUBS 0.031761f
C1436 VTAIL.n318 VSUBS 0.014228f
C1437 VTAIL.n319 VSUBS 0.013438f
C1438 VTAIL.n320 VSUBS 0.025007f
C1439 VTAIL.n321 VSUBS 0.025007f
C1440 VTAIL.n322 VSUBS 0.013438f
C1441 VTAIL.n323 VSUBS 0.013833f
C1442 VTAIL.n324 VSUBS 0.013833f
C1443 VTAIL.n325 VSUBS 0.031761f
C1444 VTAIL.n326 VSUBS 0.073646f
C1445 VTAIL.n327 VSUBS 0.014228f
C1446 VTAIL.n328 VSUBS 0.013438f
C1447 VTAIL.n329 VSUBS 0.061901f
C1448 VTAIL.n330 VSUBS 0.037014f
C1449 VTAIL.n331 VSUBS 1.93184f
C1450 VTAIL.t3 VSUBS 0.291674f
C1451 VTAIL.t0 VSUBS 0.291674f
C1452 VTAIL.n332 VSUBS 2.23251f
C1453 VTAIL.n333 VSUBS 1.11566f
C1454 VTAIL.n334 VSUBS 0.026524f
C1455 VTAIL.n335 VSUBS 0.025007f
C1456 VTAIL.n336 VSUBS 0.013438f
C1457 VTAIL.n337 VSUBS 0.031761f
C1458 VTAIL.n338 VSUBS 0.014228f
C1459 VTAIL.n339 VSUBS 0.025007f
C1460 VTAIL.n340 VSUBS 0.013438f
C1461 VTAIL.n341 VSUBS 0.031761f
C1462 VTAIL.n342 VSUBS 0.031761f
C1463 VTAIL.n343 VSUBS 0.014228f
C1464 VTAIL.n344 VSUBS 0.025007f
C1465 VTAIL.n345 VSUBS 0.013438f
C1466 VTAIL.n346 VSUBS 0.031761f
C1467 VTAIL.n347 VSUBS 0.014228f
C1468 VTAIL.n348 VSUBS 0.025007f
C1469 VTAIL.n349 VSUBS 0.013438f
C1470 VTAIL.n350 VSUBS 0.031761f
C1471 VTAIL.n351 VSUBS 0.014228f
C1472 VTAIL.n352 VSUBS 0.025007f
C1473 VTAIL.n353 VSUBS 0.013438f
C1474 VTAIL.n354 VSUBS 0.031761f
C1475 VTAIL.n355 VSUBS 0.014228f
C1476 VTAIL.n356 VSUBS 0.025007f
C1477 VTAIL.n357 VSUBS 0.013438f
C1478 VTAIL.n358 VSUBS 0.031761f
C1479 VTAIL.n359 VSUBS 0.014228f
C1480 VTAIL.n360 VSUBS 0.174506f
C1481 VTAIL.t7 VSUBS 0.06798f
C1482 VTAIL.n361 VSUBS 0.023821f
C1483 VTAIL.n362 VSUBS 0.020205f
C1484 VTAIL.n363 VSUBS 0.013438f
C1485 VTAIL.n364 VSUBS 1.56949f
C1486 VTAIL.n365 VSUBS 0.025007f
C1487 VTAIL.n366 VSUBS 0.013438f
C1488 VTAIL.n367 VSUBS 0.014228f
C1489 VTAIL.n368 VSUBS 0.031761f
C1490 VTAIL.n369 VSUBS 0.031761f
C1491 VTAIL.n370 VSUBS 0.014228f
C1492 VTAIL.n371 VSUBS 0.013438f
C1493 VTAIL.n372 VSUBS 0.025007f
C1494 VTAIL.n373 VSUBS 0.025007f
C1495 VTAIL.n374 VSUBS 0.013438f
C1496 VTAIL.n375 VSUBS 0.014228f
C1497 VTAIL.n376 VSUBS 0.031761f
C1498 VTAIL.n377 VSUBS 0.031761f
C1499 VTAIL.n378 VSUBS 0.014228f
C1500 VTAIL.n379 VSUBS 0.013438f
C1501 VTAIL.n380 VSUBS 0.025007f
C1502 VTAIL.n381 VSUBS 0.025007f
C1503 VTAIL.n382 VSUBS 0.013438f
C1504 VTAIL.n383 VSUBS 0.014228f
C1505 VTAIL.n384 VSUBS 0.031761f
C1506 VTAIL.n385 VSUBS 0.031761f
C1507 VTAIL.n386 VSUBS 0.014228f
C1508 VTAIL.n387 VSUBS 0.013438f
C1509 VTAIL.n388 VSUBS 0.025007f
C1510 VTAIL.n389 VSUBS 0.025007f
C1511 VTAIL.n390 VSUBS 0.013438f
C1512 VTAIL.n391 VSUBS 0.014228f
C1513 VTAIL.n392 VSUBS 0.031761f
C1514 VTAIL.n393 VSUBS 0.031761f
C1515 VTAIL.n394 VSUBS 0.014228f
C1516 VTAIL.n395 VSUBS 0.013438f
C1517 VTAIL.n396 VSUBS 0.025007f
C1518 VTAIL.n397 VSUBS 0.025007f
C1519 VTAIL.n398 VSUBS 0.013438f
C1520 VTAIL.n399 VSUBS 0.014228f
C1521 VTAIL.n400 VSUBS 0.031761f
C1522 VTAIL.n401 VSUBS 0.031761f
C1523 VTAIL.n402 VSUBS 0.014228f
C1524 VTAIL.n403 VSUBS 0.013438f
C1525 VTAIL.n404 VSUBS 0.025007f
C1526 VTAIL.n405 VSUBS 0.025007f
C1527 VTAIL.n406 VSUBS 0.013438f
C1528 VTAIL.n407 VSUBS 0.013833f
C1529 VTAIL.n408 VSUBS 0.013833f
C1530 VTAIL.n409 VSUBS 0.031761f
C1531 VTAIL.n410 VSUBS 0.073646f
C1532 VTAIL.n411 VSUBS 0.014228f
C1533 VTAIL.n412 VSUBS 0.013438f
C1534 VTAIL.n413 VSUBS 0.061901f
C1535 VTAIL.n414 VSUBS 0.037014f
C1536 VTAIL.n415 VSUBS 0.333134f
C1537 VTAIL.n416 VSUBS 0.026524f
C1538 VTAIL.n417 VSUBS 0.025007f
C1539 VTAIL.n418 VSUBS 0.013438f
C1540 VTAIL.n419 VSUBS 0.031761f
C1541 VTAIL.n420 VSUBS 0.014228f
C1542 VTAIL.n421 VSUBS 0.025007f
C1543 VTAIL.n422 VSUBS 0.013438f
C1544 VTAIL.n423 VSUBS 0.031761f
C1545 VTAIL.n424 VSUBS 0.031761f
C1546 VTAIL.n425 VSUBS 0.014228f
C1547 VTAIL.n426 VSUBS 0.025007f
C1548 VTAIL.n427 VSUBS 0.013438f
C1549 VTAIL.n428 VSUBS 0.031761f
C1550 VTAIL.n429 VSUBS 0.014228f
C1551 VTAIL.n430 VSUBS 0.025007f
C1552 VTAIL.n431 VSUBS 0.013438f
C1553 VTAIL.n432 VSUBS 0.031761f
C1554 VTAIL.n433 VSUBS 0.014228f
C1555 VTAIL.n434 VSUBS 0.025007f
C1556 VTAIL.n435 VSUBS 0.013438f
C1557 VTAIL.n436 VSUBS 0.031761f
C1558 VTAIL.n437 VSUBS 0.014228f
C1559 VTAIL.n438 VSUBS 0.025007f
C1560 VTAIL.n439 VSUBS 0.013438f
C1561 VTAIL.n440 VSUBS 0.031761f
C1562 VTAIL.n441 VSUBS 0.014228f
C1563 VTAIL.n442 VSUBS 0.174506f
C1564 VTAIL.t15 VSUBS 0.06798f
C1565 VTAIL.n443 VSUBS 0.023821f
C1566 VTAIL.n444 VSUBS 0.020205f
C1567 VTAIL.n445 VSUBS 0.013438f
C1568 VTAIL.n446 VSUBS 1.56949f
C1569 VTAIL.n447 VSUBS 0.025007f
C1570 VTAIL.n448 VSUBS 0.013438f
C1571 VTAIL.n449 VSUBS 0.014228f
C1572 VTAIL.n450 VSUBS 0.031761f
C1573 VTAIL.n451 VSUBS 0.031761f
C1574 VTAIL.n452 VSUBS 0.014228f
C1575 VTAIL.n453 VSUBS 0.013438f
C1576 VTAIL.n454 VSUBS 0.025007f
C1577 VTAIL.n455 VSUBS 0.025007f
C1578 VTAIL.n456 VSUBS 0.013438f
C1579 VTAIL.n457 VSUBS 0.014228f
C1580 VTAIL.n458 VSUBS 0.031761f
C1581 VTAIL.n459 VSUBS 0.031761f
C1582 VTAIL.n460 VSUBS 0.014228f
C1583 VTAIL.n461 VSUBS 0.013438f
C1584 VTAIL.n462 VSUBS 0.025007f
C1585 VTAIL.n463 VSUBS 0.025007f
C1586 VTAIL.n464 VSUBS 0.013438f
C1587 VTAIL.n465 VSUBS 0.014228f
C1588 VTAIL.n466 VSUBS 0.031761f
C1589 VTAIL.n467 VSUBS 0.031761f
C1590 VTAIL.n468 VSUBS 0.014228f
C1591 VTAIL.n469 VSUBS 0.013438f
C1592 VTAIL.n470 VSUBS 0.025007f
C1593 VTAIL.n471 VSUBS 0.025007f
C1594 VTAIL.n472 VSUBS 0.013438f
C1595 VTAIL.n473 VSUBS 0.014228f
C1596 VTAIL.n474 VSUBS 0.031761f
C1597 VTAIL.n475 VSUBS 0.031761f
C1598 VTAIL.n476 VSUBS 0.014228f
C1599 VTAIL.n477 VSUBS 0.013438f
C1600 VTAIL.n478 VSUBS 0.025007f
C1601 VTAIL.n479 VSUBS 0.025007f
C1602 VTAIL.n480 VSUBS 0.013438f
C1603 VTAIL.n481 VSUBS 0.014228f
C1604 VTAIL.n482 VSUBS 0.031761f
C1605 VTAIL.n483 VSUBS 0.031761f
C1606 VTAIL.n484 VSUBS 0.014228f
C1607 VTAIL.n485 VSUBS 0.013438f
C1608 VTAIL.n486 VSUBS 0.025007f
C1609 VTAIL.n487 VSUBS 0.025007f
C1610 VTAIL.n488 VSUBS 0.013438f
C1611 VTAIL.n489 VSUBS 0.013833f
C1612 VTAIL.n490 VSUBS 0.013833f
C1613 VTAIL.n491 VSUBS 0.031761f
C1614 VTAIL.n492 VSUBS 0.073646f
C1615 VTAIL.n493 VSUBS 0.014228f
C1616 VTAIL.n494 VSUBS 0.013438f
C1617 VTAIL.n495 VSUBS 0.061901f
C1618 VTAIL.n496 VSUBS 0.037014f
C1619 VTAIL.n497 VSUBS 0.333134f
C1620 VTAIL.t11 VSUBS 0.291674f
C1621 VTAIL.t10 VSUBS 0.291674f
C1622 VTAIL.n498 VSUBS 2.23251f
C1623 VTAIL.n499 VSUBS 1.11566f
C1624 VTAIL.n500 VSUBS 0.026524f
C1625 VTAIL.n501 VSUBS 0.025007f
C1626 VTAIL.n502 VSUBS 0.013438f
C1627 VTAIL.n503 VSUBS 0.031761f
C1628 VTAIL.n504 VSUBS 0.014228f
C1629 VTAIL.n505 VSUBS 0.025007f
C1630 VTAIL.n506 VSUBS 0.013438f
C1631 VTAIL.n507 VSUBS 0.031761f
C1632 VTAIL.n508 VSUBS 0.031761f
C1633 VTAIL.n509 VSUBS 0.014228f
C1634 VTAIL.n510 VSUBS 0.025007f
C1635 VTAIL.n511 VSUBS 0.013438f
C1636 VTAIL.n512 VSUBS 0.031761f
C1637 VTAIL.n513 VSUBS 0.014228f
C1638 VTAIL.n514 VSUBS 0.025007f
C1639 VTAIL.n515 VSUBS 0.013438f
C1640 VTAIL.n516 VSUBS 0.031761f
C1641 VTAIL.n517 VSUBS 0.014228f
C1642 VTAIL.n518 VSUBS 0.025007f
C1643 VTAIL.n519 VSUBS 0.013438f
C1644 VTAIL.n520 VSUBS 0.031761f
C1645 VTAIL.n521 VSUBS 0.014228f
C1646 VTAIL.n522 VSUBS 0.025007f
C1647 VTAIL.n523 VSUBS 0.013438f
C1648 VTAIL.n524 VSUBS 0.031761f
C1649 VTAIL.n525 VSUBS 0.014228f
C1650 VTAIL.n526 VSUBS 0.174506f
C1651 VTAIL.t9 VSUBS 0.06798f
C1652 VTAIL.n527 VSUBS 0.023821f
C1653 VTAIL.n528 VSUBS 0.020205f
C1654 VTAIL.n529 VSUBS 0.013438f
C1655 VTAIL.n530 VSUBS 1.56949f
C1656 VTAIL.n531 VSUBS 0.025007f
C1657 VTAIL.n532 VSUBS 0.013438f
C1658 VTAIL.n533 VSUBS 0.014228f
C1659 VTAIL.n534 VSUBS 0.031761f
C1660 VTAIL.n535 VSUBS 0.031761f
C1661 VTAIL.n536 VSUBS 0.014228f
C1662 VTAIL.n537 VSUBS 0.013438f
C1663 VTAIL.n538 VSUBS 0.025007f
C1664 VTAIL.n539 VSUBS 0.025007f
C1665 VTAIL.n540 VSUBS 0.013438f
C1666 VTAIL.n541 VSUBS 0.014228f
C1667 VTAIL.n542 VSUBS 0.031761f
C1668 VTAIL.n543 VSUBS 0.031761f
C1669 VTAIL.n544 VSUBS 0.014228f
C1670 VTAIL.n545 VSUBS 0.013438f
C1671 VTAIL.n546 VSUBS 0.025007f
C1672 VTAIL.n547 VSUBS 0.025007f
C1673 VTAIL.n548 VSUBS 0.013438f
C1674 VTAIL.n549 VSUBS 0.014228f
C1675 VTAIL.n550 VSUBS 0.031761f
C1676 VTAIL.n551 VSUBS 0.031761f
C1677 VTAIL.n552 VSUBS 0.014228f
C1678 VTAIL.n553 VSUBS 0.013438f
C1679 VTAIL.n554 VSUBS 0.025007f
C1680 VTAIL.n555 VSUBS 0.025007f
C1681 VTAIL.n556 VSUBS 0.013438f
C1682 VTAIL.n557 VSUBS 0.014228f
C1683 VTAIL.n558 VSUBS 0.031761f
C1684 VTAIL.n559 VSUBS 0.031761f
C1685 VTAIL.n560 VSUBS 0.014228f
C1686 VTAIL.n561 VSUBS 0.013438f
C1687 VTAIL.n562 VSUBS 0.025007f
C1688 VTAIL.n563 VSUBS 0.025007f
C1689 VTAIL.n564 VSUBS 0.013438f
C1690 VTAIL.n565 VSUBS 0.014228f
C1691 VTAIL.n566 VSUBS 0.031761f
C1692 VTAIL.n567 VSUBS 0.031761f
C1693 VTAIL.n568 VSUBS 0.014228f
C1694 VTAIL.n569 VSUBS 0.013438f
C1695 VTAIL.n570 VSUBS 0.025007f
C1696 VTAIL.n571 VSUBS 0.025007f
C1697 VTAIL.n572 VSUBS 0.013438f
C1698 VTAIL.n573 VSUBS 0.013833f
C1699 VTAIL.n574 VSUBS 0.013833f
C1700 VTAIL.n575 VSUBS 0.031761f
C1701 VTAIL.n576 VSUBS 0.073646f
C1702 VTAIL.n577 VSUBS 0.014228f
C1703 VTAIL.n578 VSUBS 0.013438f
C1704 VTAIL.n579 VSUBS 0.061901f
C1705 VTAIL.n580 VSUBS 0.037014f
C1706 VTAIL.n581 VSUBS 1.93184f
C1707 VTAIL.n582 VSUBS 0.026524f
C1708 VTAIL.n583 VSUBS 0.025007f
C1709 VTAIL.n584 VSUBS 0.013438f
C1710 VTAIL.n585 VSUBS 0.031761f
C1711 VTAIL.n586 VSUBS 0.014228f
C1712 VTAIL.n587 VSUBS 0.025007f
C1713 VTAIL.n588 VSUBS 0.013438f
C1714 VTAIL.n589 VSUBS 0.031761f
C1715 VTAIL.n590 VSUBS 0.014228f
C1716 VTAIL.n591 VSUBS 0.025007f
C1717 VTAIL.n592 VSUBS 0.013438f
C1718 VTAIL.n593 VSUBS 0.031761f
C1719 VTAIL.n594 VSUBS 0.014228f
C1720 VTAIL.n595 VSUBS 0.025007f
C1721 VTAIL.n596 VSUBS 0.013438f
C1722 VTAIL.n597 VSUBS 0.031761f
C1723 VTAIL.n598 VSUBS 0.014228f
C1724 VTAIL.n599 VSUBS 0.025007f
C1725 VTAIL.n600 VSUBS 0.013438f
C1726 VTAIL.n601 VSUBS 0.031761f
C1727 VTAIL.n602 VSUBS 0.014228f
C1728 VTAIL.n603 VSUBS 0.025007f
C1729 VTAIL.n604 VSUBS 0.013438f
C1730 VTAIL.n605 VSUBS 0.031761f
C1731 VTAIL.n606 VSUBS 0.014228f
C1732 VTAIL.n607 VSUBS 0.174506f
C1733 VTAIL.t5 VSUBS 0.06798f
C1734 VTAIL.n608 VSUBS 0.023821f
C1735 VTAIL.n609 VSUBS 0.020205f
C1736 VTAIL.n610 VSUBS 0.013438f
C1737 VTAIL.n611 VSUBS 1.56949f
C1738 VTAIL.n612 VSUBS 0.025007f
C1739 VTAIL.n613 VSUBS 0.013438f
C1740 VTAIL.n614 VSUBS 0.014228f
C1741 VTAIL.n615 VSUBS 0.031761f
C1742 VTAIL.n616 VSUBS 0.031761f
C1743 VTAIL.n617 VSUBS 0.014228f
C1744 VTAIL.n618 VSUBS 0.013438f
C1745 VTAIL.n619 VSUBS 0.025007f
C1746 VTAIL.n620 VSUBS 0.025007f
C1747 VTAIL.n621 VSUBS 0.013438f
C1748 VTAIL.n622 VSUBS 0.014228f
C1749 VTAIL.n623 VSUBS 0.031761f
C1750 VTAIL.n624 VSUBS 0.031761f
C1751 VTAIL.n625 VSUBS 0.014228f
C1752 VTAIL.n626 VSUBS 0.013438f
C1753 VTAIL.n627 VSUBS 0.025007f
C1754 VTAIL.n628 VSUBS 0.025007f
C1755 VTAIL.n629 VSUBS 0.013438f
C1756 VTAIL.n630 VSUBS 0.014228f
C1757 VTAIL.n631 VSUBS 0.031761f
C1758 VTAIL.n632 VSUBS 0.031761f
C1759 VTAIL.n633 VSUBS 0.014228f
C1760 VTAIL.n634 VSUBS 0.013438f
C1761 VTAIL.n635 VSUBS 0.025007f
C1762 VTAIL.n636 VSUBS 0.025007f
C1763 VTAIL.n637 VSUBS 0.013438f
C1764 VTAIL.n638 VSUBS 0.014228f
C1765 VTAIL.n639 VSUBS 0.031761f
C1766 VTAIL.n640 VSUBS 0.031761f
C1767 VTAIL.n641 VSUBS 0.014228f
C1768 VTAIL.n642 VSUBS 0.013438f
C1769 VTAIL.n643 VSUBS 0.025007f
C1770 VTAIL.n644 VSUBS 0.025007f
C1771 VTAIL.n645 VSUBS 0.013438f
C1772 VTAIL.n646 VSUBS 0.014228f
C1773 VTAIL.n647 VSUBS 0.031761f
C1774 VTAIL.n648 VSUBS 0.031761f
C1775 VTAIL.n649 VSUBS 0.031761f
C1776 VTAIL.n650 VSUBS 0.014228f
C1777 VTAIL.n651 VSUBS 0.013438f
C1778 VTAIL.n652 VSUBS 0.025007f
C1779 VTAIL.n653 VSUBS 0.025007f
C1780 VTAIL.n654 VSUBS 0.013438f
C1781 VTAIL.n655 VSUBS 0.013833f
C1782 VTAIL.n656 VSUBS 0.013833f
C1783 VTAIL.n657 VSUBS 0.031761f
C1784 VTAIL.n658 VSUBS 0.073646f
C1785 VTAIL.n659 VSUBS 0.014228f
C1786 VTAIL.n660 VSUBS 0.013438f
C1787 VTAIL.n661 VSUBS 0.061901f
C1788 VTAIL.n662 VSUBS 0.037014f
C1789 VTAIL.n663 VSUBS 1.92715f
C1790 VDD1.t3 VSUBS 0.374814f
C1791 VDD1.t1 VSUBS 0.374814f
C1792 VDD1.n0 VSUBS 3.07199f
C1793 VDD1.t6 VSUBS 0.374814f
C1794 VDD1.t5 VSUBS 0.374814f
C1795 VDD1.n1 VSUBS 3.07003f
C1796 VDD1.t4 VSUBS 0.374814f
C1797 VDD1.t2 VSUBS 0.374814f
C1798 VDD1.n2 VSUBS 3.07003f
C1799 VDD1.n3 VSUBS 5.900259f
C1800 VDD1.t0 VSUBS 0.374814f
C1801 VDD1.t7 VSUBS 0.374814f
C1802 VDD1.n4 VSUBS 3.04529f
C1803 VDD1.n5 VSUBS 4.8762f
C1804 VP.t1 VSUBS 3.61703f
C1805 VP.n0 VSUBS 1.34801f
C1806 VP.n1 VSUBS 0.02499f
C1807 VP.n2 VSUBS 0.042488f
C1808 VP.n3 VSUBS 0.02499f
C1809 VP.n4 VSUBS 0.036961f
C1810 VP.n5 VSUBS 0.02499f
C1811 VP.n6 VSUBS 0.036327f
C1812 VP.n7 VSUBS 0.02499f
C1813 VP.n8 VSUBS 0.032843f
C1814 VP.n9 VSUBS 0.02499f
C1815 VP.n10 VSUBS 0.029732f
C1816 VP.n11 VSUBS 0.02499f
C1817 VP.n12 VSUBS 0.028726f
C1818 VP.t6 VSUBS 3.61703f
C1819 VP.n13 VSUBS 1.34801f
C1820 VP.n14 VSUBS 0.02499f
C1821 VP.n15 VSUBS 0.042488f
C1822 VP.n16 VSUBS 0.02499f
C1823 VP.n17 VSUBS 0.036961f
C1824 VP.n18 VSUBS 0.02499f
C1825 VP.n19 VSUBS 0.036327f
C1826 VP.n20 VSUBS 0.02499f
C1827 VP.n21 VSUBS 0.032843f
C1828 VP.t0 VSUBS 3.97395f
C1829 VP.t4 VSUBS 3.61703f
C1830 VP.n22 VSUBS 1.34036f
C1831 VP.n23 VSUBS 1.27923f
C1832 VP.n24 VSUBS 0.312617f
C1833 VP.n25 VSUBS 0.02499f
C1834 VP.n26 VSUBS 0.046341f
C1835 VP.n27 VSUBS 0.046341f
C1836 VP.n28 VSUBS 0.036327f
C1837 VP.n29 VSUBS 0.02499f
C1838 VP.n30 VSUBS 0.02499f
C1839 VP.n31 VSUBS 0.02499f
C1840 VP.n32 VSUBS 0.046341f
C1841 VP.n33 VSUBS 0.046341f
C1842 VP.t5 VSUBS 3.61703f
C1843 VP.n34 VSUBS 1.25641f
C1844 VP.n35 VSUBS 0.032843f
C1845 VP.n36 VSUBS 0.02499f
C1846 VP.n37 VSUBS 0.02499f
C1847 VP.n38 VSUBS 0.02499f
C1848 VP.n39 VSUBS 0.046341f
C1849 VP.n40 VSUBS 0.046774f
C1850 VP.n41 VSUBS 0.029732f
C1851 VP.n42 VSUBS 0.02499f
C1852 VP.n43 VSUBS 0.02499f
C1853 VP.n44 VSUBS 0.02499f
C1854 VP.n45 VSUBS 0.046341f
C1855 VP.n46 VSUBS 0.046341f
C1856 VP.n47 VSUBS 0.028726f
C1857 VP.n48 VSUBS 0.040327f
C1858 VP.n49 VSUBS 1.74291f
C1859 VP.t7 VSUBS 3.61703f
C1860 VP.n50 VSUBS 1.34801f
C1861 VP.n51 VSUBS 1.75855f
C1862 VP.n52 VSUBS 0.040327f
C1863 VP.n53 VSUBS 0.02499f
C1864 VP.n54 VSUBS 0.046341f
C1865 VP.n55 VSUBS 0.046341f
C1866 VP.n56 VSUBS 0.042488f
C1867 VP.n57 VSUBS 0.02499f
C1868 VP.n58 VSUBS 0.02499f
C1869 VP.n59 VSUBS 0.02499f
C1870 VP.n60 VSUBS 0.046774f
C1871 VP.n61 VSUBS 0.046341f
C1872 VP.t2 VSUBS 3.61703f
C1873 VP.n62 VSUBS 1.25641f
C1874 VP.n63 VSUBS 0.036961f
C1875 VP.n64 VSUBS 0.02499f
C1876 VP.n65 VSUBS 0.02499f
C1877 VP.n66 VSUBS 0.02499f
C1878 VP.n67 VSUBS 0.046341f
C1879 VP.n68 VSUBS 0.046341f
C1880 VP.n69 VSUBS 0.036327f
C1881 VP.n70 VSUBS 0.02499f
C1882 VP.n71 VSUBS 0.02499f
C1883 VP.n72 VSUBS 0.02499f
C1884 VP.n73 VSUBS 0.046341f
C1885 VP.n74 VSUBS 0.046341f
C1886 VP.t3 VSUBS 3.61703f
C1887 VP.n75 VSUBS 1.25641f
C1888 VP.n76 VSUBS 0.032843f
C1889 VP.n77 VSUBS 0.02499f
C1890 VP.n78 VSUBS 0.02499f
C1891 VP.n79 VSUBS 0.02499f
C1892 VP.n80 VSUBS 0.046341f
C1893 VP.n81 VSUBS 0.046774f
C1894 VP.n82 VSUBS 0.029732f
C1895 VP.n83 VSUBS 0.02499f
C1896 VP.n84 VSUBS 0.02499f
C1897 VP.n85 VSUBS 0.02499f
C1898 VP.n86 VSUBS 0.046341f
C1899 VP.n87 VSUBS 0.046341f
C1900 VP.n88 VSUBS 0.028726f
C1901 VP.n89 VSUBS 0.040327f
C1902 VP.n90 VSUBS 0.071634f
.ends

