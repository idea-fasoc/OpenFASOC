* NGSPICE file created from diff_pair_sample_0536.ext - technology: sky130A

.subckt diff_pair_sample_0536 VTAIL VN VP B VDD2 VDD1
X0 B.t11 B.t9 B.t10 w_n3274_n4326# sky130_fd_pr__pfet_01v8 ad=6.5481 pd=34.36 as=0 ps=0 w=16.79 l=3.51
X1 B.t8 B.t6 B.t7 w_n3274_n4326# sky130_fd_pr__pfet_01v8 ad=6.5481 pd=34.36 as=0 ps=0 w=16.79 l=3.51
X2 VDD1.t3 VP.t0 VTAIL.t5 w_n3274_n4326# sky130_fd_pr__pfet_01v8 ad=2.77035 pd=17.12 as=6.5481 ps=34.36 w=16.79 l=3.51
X3 VTAIL.t2 VN.t0 VDD2.t3 w_n3274_n4326# sky130_fd_pr__pfet_01v8 ad=6.5481 pd=34.36 as=2.77035 ps=17.12 w=16.79 l=3.51
X4 VDD2.t2 VN.t1 VTAIL.t3 w_n3274_n4326# sky130_fd_pr__pfet_01v8 ad=2.77035 pd=17.12 as=6.5481 ps=34.36 w=16.79 l=3.51
X5 VTAIL.t1 VN.t2 VDD2.t1 w_n3274_n4326# sky130_fd_pr__pfet_01v8 ad=6.5481 pd=34.36 as=2.77035 ps=17.12 w=16.79 l=3.51
X6 VDD1.t2 VP.t1 VTAIL.t7 w_n3274_n4326# sky130_fd_pr__pfet_01v8 ad=2.77035 pd=17.12 as=6.5481 ps=34.36 w=16.79 l=3.51
X7 VTAIL.t6 VP.t2 VDD1.t1 w_n3274_n4326# sky130_fd_pr__pfet_01v8 ad=6.5481 pd=34.36 as=2.77035 ps=17.12 w=16.79 l=3.51
X8 B.t5 B.t3 B.t4 w_n3274_n4326# sky130_fd_pr__pfet_01v8 ad=6.5481 pd=34.36 as=0 ps=0 w=16.79 l=3.51
X9 VTAIL.t4 VP.t3 VDD1.t0 w_n3274_n4326# sky130_fd_pr__pfet_01v8 ad=6.5481 pd=34.36 as=2.77035 ps=17.12 w=16.79 l=3.51
X10 VDD2.t0 VN.t3 VTAIL.t0 w_n3274_n4326# sky130_fd_pr__pfet_01v8 ad=2.77035 pd=17.12 as=6.5481 ps=34.36 w=16.79 l=3.51
X11 B.t2 B.t0 B.t1 w_n3274_n4326# sky130_fd_pr__pfet_01v8 ad=6.5481 pd=34.36 as=0 ps=0 w=16.79 l=3.51
R0 B.n588 B.n87 585
R1 B.n590 B.n589 585
R2 B.n591 B.n86 585
R3 B.n593 B.n592 585
R4 B.n594 B.n85 585
R5 B.n596 B.n595 585
R6 B.n597 B.n84 585
R7 B.n599 B.n598 585
R8 B.n600 B.n83 585
R9 B.n602 B.n601 585
R10 B.n603 B.n82 585
R11 B.n605 B.n604 585
R12 B.n606 B.n81 585
R13 B.n608 B.n607 585
R14 B.n609 B.n80 585
R15 B.n611 B.n610 585
R16 B.n612 B.n79 585
R17 B.n614 B.n613 585
R18 B.n615 B.n78 585
R19 B.n617 B.n616 585
R20 B.n618 B.n77 585
R21 B.n620 B.n619 585
R22 B.n621 B.n76 585
R23 B.n623 B.n622 585
R24 B.n624 B.n75 585
R25 B.n626 B.n625 585
R26 B.n627 B.n74 585
R27 B.n629 B.n628 585
R28 B.n630 B.n73 585
R29 B.n632 B.n631 585
R30 B.n633 B.n72 585
R31 B.n635 B.n634 585
R32 B.n636 B.n71 585
R33 B.n638 B.n637 585
R34 B.n639 B.n70 585
R35 B.n641 B.n640 585
R36 B.n642 B.n69 585
R37 B.n644 B.n643 585
R38 B.n645 B.n68 585
R39 B.n647 B.n646 585
R40 B.n648 B.n67 585
R41 B.n650 B.n649 585
R42 B.n651 B.n66 585
R43 B.n653 B.n652 585
R44 B.n654 B.n65 585
R45 B.n656 B.n655 585
R46 B.n657 B.n64 585
R47 B.n659 B.n658 585
R48 B.n660 B.n63 585
R49 B.n662 B.n661 585
R50 B.n663 B.n62 585
R51 B.n665 B.n664 585
R52 B.n666 B.n61 585
R53 B.n668 B.n667 585
R54 B.n669 B.n60 585
R55 B.n671 B.n670 585
R56 B.n673 B.n57 585
R57 B.n675 B.n674 585
R58 B.n676 B.n56 585
R59 B.n678 B.n677 585
R60 B.n679 B.n55 585
R61 B.n681 B.n680 585
R62 B.n682 B.n54 585
R63 B.n684 B.n683 585
R64 B.n685 B.n51 585
R65 B.n688 B.n687 585
R66 B.n689 B.n50 585
R67 B.n691 B.n690 585
R68 B.n692 B.n49 585
R69 B.n694 B.n693 585
R70 B.n695 B.n48 585
R71 B.n697 B.n696 585
R72 B.n698 B.n47 585
R73 B.n700 B.n699 585
R74 B.n701 B.n46 585
R75 B.n703 B.n702 585
R76 B.n704 B.n45 585
R77 B.n706 B.n705 585
R78 B.n707 B.n44 585
R79 B.n709 B.n708 585
R80 B.n710 B.n43 585
R81 B.n712 B.n711 585
R82 B.n713 B.n42 585
R83 B.n715 B.n714 585
R84 B.n716 B.n41 585
R85 B.n718 B.n717 585
R86 B.n719 B.n40 585
R87 B.n721 B.n720 585
R88 B.n722 B.n39 585
R89 B.n724 B.n723 585
R90 B.n725 B.n38 585
R91 B.n727 B.n726 585
R92 B.n728 B.n37 585
R93 B.n730 B.n729 585
R94 B.n731 B.n36 585
R95 B.n733 B.n732 585
R96 B.n734 B.n35 585
R97 B.n736 B.n735 585
R98 B.n737 B.n34 585
R99 B.n739 B.n738 585
R100 B.n740 B.n33 585
R101 B.n742 B.n741 585
R102 B.n743 B.n32 585
R103 B.n745 B.n744 585
R104 B.n746 B.n31 585
R105 B.n748 B.n747 585
R106 B.n749 B.n30 585
R107 B.n751 B.n750 585
R108 B.n752 B.n29 585
R109 B.n754 B.n753 585
R110 B.n755 B.n28 585
R111 B.n757 B.n756 585
R112 B.n758 B.n27 585
R113 B.n760 B.n759 585
R114 B.n761 B.n26 585
R115 B.n763 B.n762 585
R116 B.n764 B.n25 585
R117 B.n766 B.n765 585
R118 B.n767 B.n24 585
R119 B.n769 B.n768 585
R120 B.n770 B.n23 585
R121 B.n587 B.n586 585
R122 B.n585 B.n88 585
R123 B.n584 B.n583 585
R124 B.n582 B.n89 585
R125 B.n581 B.n580 585
R126 B.n579 B.n90 585
R127 B.n578 B.n577 585
R128 B.n576 B.n91 585
R129 B.n575 B.n574 585
R130 B.n573 B.n92 585
R131 B.n572 B.n571 585
R132 B.n570 B.n93 585
R133 B.n569 B.n568 585
R134 B.n567 B.n94 585
R135 B.n566 B.n565 585
R136 B.n564 B.n95 585
R137 B.n563 B.n562 585
R138 B.n561 B.n96 585
R139 B.n560 B.n559 585
R140 B.n558 B.n97 585
R141 B.n557 B.n556 585
R142 B.n555 B.n98 585
R143 B.n554 B.n553 585
R144 B.n552 B.n99 585
R145 B.n551 B.n550 585
R146 B.n549 B.n100 585
R147 B.n548 B.n547 585
R148 B.n546 B.n101 585
R149 B.n545 B.n544 585
R150 B.n543 B.n102 585
R151 B.n542 B.n541 585
R152 B.n540 B.n103 585
R153 B.n539 B.n538 585
R154 B.n537 B.n104 585
R155 B.n536 B.n535 585
R156 B.n534 B.n105 585
R157 B.n533 B.n532 585
R158 B.n531 B.n106 585
R159 B.n530 B.n529 585
R160 B.n528 B.n107 585
R161 B.n527 B.n526 585
R162 B.n525 B.n108 585
R163 B.n524 B.n523 585
R164 B.n522 B.n109 585
R165 B.n521 B.n520 585
R166 B.n519 B.n110 585
R167 B.n518 B.n517 585
R168 B.n516 B.n111 585
R169 B.n515 B.n514 585
R170 B.n513 B.n112 585
R171 B.n512 B.n511 585
R172 B.n510 B.n113 585
R173 B.n509 B.n508 585
R174 B.n507 B.n114 585
R175 B.n506 B.n505 585
R176 B.n504 B.n115 585
R177 B.n503 B.n502 585
R178 B.n501 B.n116 585
R179 B.n500 B.n499 585
R180 B.n498 B.n117 585
R181 B.n497 B.n496 585
R182 B.n495 B.n118 585
R183 B.n494 B.n493 585
R184 B.n492 B.n119 585
R185 B.n491 B.n490 585
R186 B.n489 B.n120 585
R187 B.n488 B.n487 585
R188 B.n486 B.n121 585
R189 B.n485 B.n484 585
R190 B.n483 B.n122 585
R191 B.n482 B.n481 585
R192 B.n480 B.n123 585
R193 B.n479 B.n478 585
R194 B.n477 B.n124 585
R195 B.n476 B.n475 585
R196 B.n474 B.n125 585
R197 B.n473 B.n472 585
R198 B.n471 B.n126 585
R199 B.n470 B.n469 585
R200 B.n468 B.n127 585
R201 B.n467 B.n466 585
R202 B.n465 B.n128 585
R203 B.n464 B.n463 585
R204 B.n462 B.n129 585
R205 B.n461 B.n460 585
R206 B.n278 B.n277 585
R207 B.n279 B.n194 585
R208 B.n281 B.n280 585
R209 B.n282 B.n193 585
R210 B.n284 B.n283 585
R211 B.n285 B.n192 585
R212 B.n287 B.n286 585
R213 B.n288 B.n191 585
R214 B.n290 B.n289 585
R215 B.n291 B.n190 585
R216 B.n293 B.n292 585
R217 B.n294 B.n189 585
R218 B.n296 B.n295 585
R219 B.n297 B.n188 585
R220 B.n299 B.n298 585
R221 B.n300 B.n187 585
R222 B.n302 B.n301 585
R223 B.n303 B.n186 585
R224 B.n305 B.n304 585
R225 B.n306 B.n185 585
R226 B.n308 B.n307 585
R227 B.n309 B.n184 585
R228 B.n311 B.n310 585
R229 B.n312 B.n183 585
R230 B.n314 B.n313 585
R231 B.n315 B.n182 585
R232 B.n317 B.n316 585
R233 B.n318 B.n181 585
R234 B.n320 B.n319 585
R235 B.n321 B.n180 585
R236 B.n323 B.n322 585
R237 B.n324 B.n179 585
R238 B.n326 B.n325 585
R239 B.n327 B.n178 585
R240 B.n329 B.n328 585
R241 B.n330 B.n177 585
R242 B.n332 B.n331 585
R243 B.n333 B.n176 585
R244 B.n335 B.n334 585
R245 B.n336 B.n175 585
R246 B.n338 B.n337 585
R247 B.n339 B.n174 585
R248 B.n341 B.n340 585
R249 B.n342 B.n173 585
R250 B.n344 B.n343 585
R251 B.n345 B.n172 585
R252 B.n347 B.n346 585
R253 B.n348 B.n171 585
R254 B.n350 B.n349 585
R255 B.n351 B.n170 585
R256 B.n353 B.n352 585
R257 B.n354 B.n169 585
R258 B.n356 B.n355 585
R259 B.n357 B.n168 585
R260 B.n359 B.n358 585
R261 B.n360 B.n165 585
R262 B.n363 B.n362 585
R263 B.n364 B.n164 585
R264 B.n366 B.n365 585
R265 B.n367 B.n163 585
R266 B.n369 B.n368 585
R267 B.n370 B.n162 585
R268 B.n372 B.n371 585
R269 B.n373 B.n161 585
R270 B.n375 B.n374 585
R271 B.n377 B.n376 585
R272 B.n378 B.n157 585
R273 B.n380 B.n379 585
R274 B.n381 B.n156 585
R275 B.n383 B.n382 585
R276 B.n384 B.n155 585
R277 B.n386 B.n385 585
R278 B.n387 B.n154 585
R279 B.n389 B.n388 585
R280 B.n390 B.n153 585
R281 B.n392 B.n391 585
R282 B.n393 B.n152 585
R283 B.n395 B.n394 585
R284 B.n396 B.n151 585
R285 B.n398 B.n397 585
R286 B.n399 B.n150 585
R287 B.n401 B.n400 585
R288 B.n402 B.n149 585
R289 B.n404 B.n403 585
R290 B.n405 B.n148 585
R291 B.n407 B.n406 585
R292 B.n408 B.n147 585
R293 B.n410 B.n409 585
R294 B.n411 B.n146 585
R295 B.n413 B.n412 585
R296 B.n414 B.n145 585
R297 B.n416 B.n415 585
R298 B.n417 B.n144 585
R299 B.n419 B.n418 585
R300 B.n420 B.n143 585
R301 B.n422 B.n421 585
R302 B.n423 B.n142 585
R303 B.n425 B.n424 585
R304 B.n426 B.n141 585
R305 B.n428 B.n427 585
R306 B.n429 B.n140 585
R307 B.n431 B.n430 585
R308 B.n432 B.n139 585
R309 B.n434 B.n433 585
R310 B.n435 B.n138 585
R311 B.n437 B.n436 585
R312 B.n438 B.n137 585
R313 B.n440 B.n439 585
R314 B.n441 B.n136 585
R315 B.n443 B.n442 585
R316 B.n444 B.n135 585
R317 B.n446 B.n445 585
R318 B.n447 B.n134 585
R319 B.n449 B.n448 585
R320 B.n450 B.n133 585
R321 B.n452 B.n451 585
R322 B.n453 B.n132 585
R323 B.n455 B.n454 585
R324 B.n456 B.n131 585
R325 B.n458 B.n457 585
R326 B.n459 B.n130 585
R327 B.n276 B.n195 585
R328 B.n275 B.n274 585
R329 B.n273 B.n196 585
R330 B.n272 B.n271 585
R331 B.n270 B.n197 585
R332 B.n269 B.n268 585
R333 B.n267 B.n198 585
R334 B.n266 B.n265 585
R335 B.n264 B.n199 585
R336 B.n263 B.n262 585
R337 B.n261 B.n200 585
R338 B.n260 B.n259 585
R339 B.n258 B.n201 585
R340 B.n257 B.n256 585
R341 B.n255 B.n202 585
R342 B.n254 B.n253 585
R343 B.n252 B.n203 585
R344 B.n251 B.n250 585
R345 B.n249 B.n204 585
R346 B.n248 B.n247 585
R347 B.n246 B.n205 585
R348 B.n245 B.n244 585
R349 B.n243 B.n206 585
R350 B.n242 B.n241 585
R351 B.n240 B.n207 585
R352 B.n239 B.n238 585
R353 B.n237 B.n208 585
R354 B.n236 B.n235 585
R355 B.n234 B.n209 585
R356 B.n233 B.n232 585
R357 B.n231 B.n210 585
R358 B.n230 B.n229 585
R359 B.n228 B.n211 585
R360 B.n227 B.n226 585
R361 B.n225 B.n212 585
R362 B.n224 B.n223 585
R363 B.n222 B.n213 585
R364 B.n221 B.n220 585
R365 B.n219 B.n214 585
R366 B.n218 B.n217 585
R367 B.n216 B.n215 585
R368 B.n2 B.n0 585
R369 B.n833 B.n1 585
R370 B.n832 B.n831 585
R371 B.n830 B.n3 585
R372 B.n829 B.n828 585
R373 B.n827 B.n4 585
R374 B.n826 B.n825 585
R375 B.n824 B.n5 585
R376 B.n823 B.n822 585
R377 B.n821 B.n6 585
R378 B.n820 B.n819 585
R379 B.n818 B.n7 585
R380 B.n817 B.n816 585
R381 B.n815 B.n8 585
R382 B.n814 B.n813 585
R383 B.n812 B.n9 585
R384 B.n811 B.n810 585
R385 B.n809 B.n10 585
R386 B.n808 B.n807 585
R387 B.n806 B.n11 585
R388 B.n805 B.n804 585
R389 B.n803 B.n12 585
R390 B.n802 B.n801 585
R391 B.n800 B.n13 585
R392 B.n799 B.n798 585
R393 B.n797 B.n14 585
R394 B.n796 B.n795 585
R395 B.n794 B.n15 585
R396 B.n793 B.n792 585
R397 B.n791 B.n16 585
R398 B.n790 B.n789 585
R399 B.n788 B.n17 585
R400 B.n787 B.n786 585
R401 B.n785 B.n18 585
R402 B.n784 B.n783 585
R403 B.n782 B.n19 585
R404 B.n781 B.n780 585
R405 B.n779 B.n20 585
R406 B.n778 B.n777 585
R407 B.n776 B.n21 585
R408 B.n775 B.n774 585
R409 B.n773 B.n22 585
R410 B.n772 B.n771 585
R411 B.n835 B.n834 585
R412 B.n158 B.t11 536.319
R413 B.n58 B.t7 536.319
R414 B.n166 B.t2 536.319
R415 B.n52 B.t4 536.319
R416 B.n278 B.n195 497.305
R417 B.n772 B.n23 497.305
R418 B.n460 B.n459 497.305
R419 B.n586 B.n87 497.305
R420 B.n159 B.t10 461.846
R421 B.n59 B.t8 461.846
R422 B.n167 B.t1 461.846
R423 B.n53 B.t5 461.846
R424 B.n158 B.t9 324.385
R425 B.n166 B.t0 324.385
R426 B.n52 B.t3 324.385
R427 B.n58 B.t6 324.385
R428 B.n274 B.n195 163.367
R429 B.n274 B.n273 163.367
R430 B.n273 B.n272 163.367
R431 B.n272 B.n197 163.367
R432 B.n268 B.n197 163.367
R433 B.n268 B.n267 163.367
R434 B.n267 B.n266 163.367
R435 B.n266 B.n199 163.367
R436 B.n262 B.n199 163.367
R437 B.n262 B.n261 163.367
R438 B.n261 B.n260 163.367
R439 B.n260 B.n201 163.367
R440 B.n256 B.n201 163.367
R441 B.n256 B.n255 163.367
R442 B.n255 B.n254 163.367
R443 B.n254 B.n203 163.367
R444 B.n250 B.n203 163.367
R445 B.n250 B.n249 163.367
R446 B.n249 B.n248 163.367
R447 B.n248 B.n205 163.367
R448 B.n244 B.n205 163.367
R449 B.n244 B.n243 163.367
R450 B.n243 B.n242 163.367
R451 B.n242 B.n207 163.367
R452 B.n238 B.n207 163.367
R453 B.n238 B.n237 163.367
R454 B.n237 B.n236 163.367
R455 B.n236 B.n209 163.367
R456 B.n232 B.n209 163.367
R457 B.n232 B.n231 163.367
R458 B.n231 B.n230 163.367
R459 B.n230 B.n211 163.367
R460 B.n226 B.n211 163.367
R461 B.n226 B.n225 163.367
R462 B.n225 B.n224 163.367
R463 B.n224 B.n213 163.367
R464 B.n220 B.n213 163.367
R465 B.n220 B.n219 163.367
R466 B.n219 B.n218 163.367
R467 B.n218 B.n215 163.367
R468 B.n215 B.n2 163.367
R469 B.n834 B.n2 163.367
R470 B.n834 B.n833 163.367
R471 B.n833 B.n832 163.367
R472 B.n832 B.n3 163.367
R473 B.n828 B.n3 163.367
R474 B.n828 B.n827 163.367
R475 B.n827 B.n826 163.367
R476 B.n826 B.n5 163.367
R477 B.n822 B.n5 163.367
R478 B.n822 B.n821 163.367
R479 B.n821 B.n820 163.367
R480 B.n820 B.n7 163.367
R481 B.n816 B.n7 163.367
R482 B.n816 B.n815 163.367
R483 B.n815 B.n814 163.367
R484 B.n814 B.n9 163.367
R485 B.n810 B.n9 163.367
R486 B.n810 B.n809 163.367
R487 B.n809 B.n808 163.367
R488 B.n808 B.n11 163.367
R489 B.n804 B.n11 163.367
R490 B.n804 B.n803 163.367
R491 B.n803 B.n802 163.367
R492 B.n802 B.n13 163.367
R493 B.n798 B.n13 163.367
R494 B.n798 B.n797 163.367
R495 B.n797 B.n796 163.367
R496 B.n796 B.n15 163.367
R497 B.n792 B.n15 163.367
R498 B.n792 B.n791 163.367
R499 B.n791 B.n790 163.367
R500 B.n790 B.n17 163.367
R501 B.n786 B.n17 163.367
R502 B.n786 B.n785 163.367
R503 B.n785 B.n784 163.367
R504 B.n784 B.n19 163.367
R505 B.n780 B.n19 163.367
R506 B.n780 B.n779 163.367
R507 B.n779 B.n778 163.367
R508 B.n778 B.n21 163.367
R509 B.n774 B.n21 163.367
R510 B.n774 B.n773 163.367
R511 B.n773 B.n772 163.367
R512 B.n279 B.n278 163.367
R513 B.n280 B.n279 163.367
R514 B.n280 B.n193 163.367
R515 B.n284 B.n193 163.367
R516 B.n285 B.n284 163.367
R517 B.n286 B.n285 163.367
R518 B.n286 B.n191 163.367
R519 B.n290 B.n191 163.367
R520 B.n291 B.n290 163.367
R521 B.n292 B.n291 163.367
R522 B.n292 B.n189 163.367
R523 B.n296 B.n189 163.367
R524 B.n297 B.n296 163.367
R525 B.n298 B.n297 163.367
R526 B.n298 B.n187 163.367
R527 B.n302 B.n187 163.367
R528 B.n303 B.n302 163.367
R529 B.n304 B.n303 163.367
R530 B.n304 B.n185 163.367
R531 B.n308 B.n185 163.367
R532 B.n309 B.n308 163.367
R533 B.n310 B.n309 163.367
R534 B.n310 B.n183 163.367
R535 B.n314 B.n183 163.367
R536 B.n315 B.n314 163.367
R537 B.n316 B.n315 163.367
R538 B.n316 B.n181 163.367
R539 B.n320 B.n181 163.367
R540 B.n321 B.n320 163.367
R541 B.n322 B.n321 163.367
R542 B.n322 B.n179 163.367
R543 B.n326 B.n179 163.367
R544 B.n327 B.n326 163.367
R545 B.n328 B.n327 163.367
R546 B.n328 B.n177 163.367
R547 B.n332 B.n177 163.367
R548 B.n333 B.n332 163.367
R549 B.n334 B.n333 163.367
R550 B.n334 B.n175 163.367
R551 B.n338 B.n175 163.367
R552 B.n339 B.n338 163.367
R553 B.n340 B.n339 163.367
R554 B.n340 B.n173 163.367
R555 B.n344 B.n173 163.367
R556 B.n345 B.n344 163.367
R557 B.n346 B.n345 163.367
R558 B.n346 B.n171 163.367
R559 B.n350 B.n171 163.367
R560 B.n351 B.n350 163.367
R561 B.n352 B.n351 163.367
R562 B.n352 B.n169 163.367
R563 B.n356 B.n169 163.367
R564 B.n357 B.n356 163.367
R565 B.n358 B.n357 163.367
R566 B.n358 B.n165 163.367
R567 B.n363 B.n165 163.367
R568 B.n364 B.n363 163.367
R569 B.n365 B.n364 163.367
R570 B.n365 B.n163 163.367
R571 B.n369 B.n163 163.367
R572 B.n370 B.n369 163.367
R573 B.n371 B.n370 163.367
R574 B.n371 B.n161 163.367
R575 B.n375 B.n161 163.367
R576 B.n376 B.n375 163.367
R577 B.n376 B.n157 163.367
R578 B.n380 B.n157 163.367
R579 B.n381 B.n380 163.367
R580 B.n382 B.n381 163.367
R581 B.n382 B.n155 163.367
R582 B.n386 B.n155 163.367
R583 B.n387 B.n386 163.367
R584 B.n388 B.n387 163.367
R585 B.n388 B.n153 163.367
R586 B.n392 B.n153 163.367
R587 B.n393 B.n392 163.367
R588 B.n394 B.n393 163.367
R589 B.n394 B.n151 163.367
R590 B.n398 B.n151 163.367
R591 B.n399 B.n398 163.367
R592 B.n400 B.n399 163.367
R593 B.n400 B.n149 163.367
R594 B.n404 B.n149 163.367
R595 B.n405 B.n404 163.367
R596 B.n406 B.n405 163.367
R597 B.n406 B.n147 163.367
R598 B.n410 B.n147 163.367
R599 B.n411 B.n410 163.367
R600 B.n412 B.n411 163.367
R601 B.n412 B.n145 163.367
R602 B.n416 B.n145 163.367
R603 B.n417 B.n416 163.367
R604 B.n418 B.n417 163.367
R605 B.n418 B.n143 163.367
R606 B.n422 B.n143 163.367
R607 B.n423 B.n422 163.367
R608 B.n424 B.n423 163.367
R609 B.n424 B.n141 163.367
R610 B.n428 B.n141 163.367
R611 B.n429 B.n428 163.367
R612 B.n430 B.n429 163.367
R613 B.n430 B.n139 163.367
R614 B.n434 B.n139 163.367
R615 B.n435 B.n434 163.367
R616 B.n436 B.n435 163.367
R617 B.n436 B.n137 163.367
R618 B.n440 B.n137 163.367
R619 B.n441 B.n440 163.367
R620 B.n442 B.n441 163.367
R621 B.n442 B.n135 163.367
R622 B.n446 B.n135 163.367
R623 B.n447 B.n446 163.367
R624 B.n448 B.n447 163.367
R625 B.n448 B.n133 163.367
R626 B.n452 B.n133 163.367
R627 B.n453 B.n452 163.367
R628 B.n454 B.n453 163.367
R629 B.n454 B.n131 163.367
R630 B.n458 B.n131 163.367
R631 B.n459 B.n458 163.367
R632 B.n460 B.n129 163.367
R633 B.n464 B.n129 163.367
R634 B.n465 B.n464 163.367
R635 B.n466 B.n465 163.367
R636 B.n466 B.n127 163.367
R637 B.n470 B.n127 163.367
R638 B.n471 B.n470 163.367
R639 B.n472 B.n471 163.367
R640 B.n472 B.n125 163.367
R641 B.n476 B.n125 163.367
R642 B.n477 B.n476 163.367
R643 B.n478 B.n477 163.367
R644 B.n478 B.n123 163.367
R645 B.n482 B.n123 163.367
R646 B.n483 B.n482 163.367
R647 B.n484 B.n483 163.367
R648 B.n484 B.n121 163.367
R649 B.n488 B.n121 163.367
R650 B.n489 B.n488 163.367
R651 B.n490 B.n489 163.367
R652 B.n490 B.n119 163.367
R653 B.n494 B.n119 163.367
R654 B.n495 B.n494 163.367
R655 B.n496 B.n495 163.367
R656 B.n496 B.n117 163.367
R657 B.n500 B.n117 163.367
R658 B.n501 B.n500 163.367
R659 B.n502 B.n501 163.367
R660 B.n502 B.n115 163.367
R661 B.n506 B.n115 163.367
R662 B.n507 B.n506 163.367
R663 B.n508 B.n507 163.367
R664 B.n508 B.n113 163.367
R665 B.n512 B.n113 163.367
R666 B.n513 B.n512 163.367
R667 B.n514 B.n513 163.367
R668 B.n514 B.n111 163.367
R669 B.n518 B.n111 163.367
R670 B.n519 B.n518 163.367
R671 B.n520 B.n519 163.367
R672 B.n520 B.n109 163.367
R673 B.n524 B.n109 163.367
R674 B.n525 B.n524 163.367
R675 B.n526 B.n525 163.367
R676 B.n526 B.n107 163.367
R677 B.n530 B.n107 163.367
R678 B.n531 B.n530 163.367
R679 B.n532 B.n531 163.367
R680 B.n532 B.n105 163.367
R681 B.n536 B.n105 163.367
R682 B.n537 B.n536 163.367
R683 B.n538 B.n537 163.367
R684 B.n538 B.n103 163.367
R685 B.n542 B.n103 163.367
R686 B.n543 B.n542 163.367
R687 B.n544 B.n543 163.367
R688 B.n544 B.n101 163.367
R689 B.n548 B.n101 163.367
R690 B.n549 B.n548 163.367
R691 B.n550 B.n549 163.367
R692 B.n550 B.n99 163.367
R693 B.n554 B.n99 163.367
R694 B.n555 B.n554 163.367
R695 B.n556 B.n555 163.367
R696 B.n556 B.n97 163.367
R697 B.n560 B.n97 163.367
R698 B.n561 B.n560 163.367
R699 B.n562 B.n561 163.367
R700 B.n562 B.n95 163.367
R701 B.n566 B.n95 163.367
R702 B.n567 B.n566 163.367
R703 B.n568 B.n567 163.367
R704 B.n568 B.n93 163.367
R705 B.n572 B.n93 163.367
R706 B.n573 B.n572 163.367
R707 B.n574 B.n573 163.367
R708 B.n574 B.n91 163.367
R709 B.n578 B.n91 163.367
R710 B.n579 B.n578 163.367
R711 B.n580 B.n579 163.367
R712 B.n580 B.n89 163.367
R713 B.n584 B.n89 163.367
R714 B.n585 B.n584 163.367
R715 B.n586 B.n585 163.367
R716 B.n768 B.n23 163.367
R717 B.n768 B.n767 163.367
R718 B.n767 B.n766 163.367
R719 B.n766 B.n25 163.367
R720 B.n762 B.n25 163.367
R721 B.n762 B.n761 163.367
R722 B.n761 B.n760 163.367
R723 B.n760 B.n27 163.367
R724 B.n756 B.n27 163.367
R725 B.n756 B.n755 163.367
R726 B.n755 B.n754 163.367
R727 B.n754 B.n29 163.367
R728 B.n750 B.n29 163.367
R729 B.n750 B.n749 163.367
R730 B.n749 B.n748 163.367
R731 B.n748 B.n31 163.367
R732 B.n744 B.n31 163.367
R733 B.n744 B.n743 163.367
R734 B.n743 B.n742 163.367
R735 B.n742 B.n33 163.367
R736 B.n738 B.n33 163.367
R737 B.n738 B.n737 163.367
R738 B.n737 B.n736 163.367
R739 B.n736 B.n35 163.367
R740 B.n732 B.n35 163.367
R741 B.n732 B.n731 163.367
R742 B.n731 B.n730 163.367
R743 B.n730 B.n37 163.367
R744 B.n726 B.n37 163.367
R745 B.n726 B.n725 163.367
R746 B.n725 B.n724 163.367
R747 B.n724 B.n39 163.367
R748 B.n720 B.n39 163.367
R749 B.n720 B.n719 163.367
R750 B.n719 B.n718 163.367
R751 B.n718 B.n41 163.367
R752 B.n714 B.n41 163.367
R753 B.n714 B.n713 163.367
R754 B.n713 B.n712 163.367
R755 B.n712 B.n43 163.367
R756 B.n708 B.n43 163.367
R757 B.n708 B.n707 163.367
R758 B.n707 B.n706 163.367
R759 B.n706 B.n45 163.367
R760 B.n702 B.n45 163.367
R761 B.n702 B.n701 163.367
R762 B.n701 B.n700 163.367
R763 B.n700 B.n47 163.367
R764 B.n696 B.n47 163.367
R765 B.n696 B.n695 163.367
R766 B.n695 B.n694 163.367
R767 B.n694 B.n49 163.367
R768 B.n690 B.n49 163.367
R769 B.n690 B.n689 163.367
R770 B.n689 B.n688 163.367
R771 B.n688 B.n51 163.367
R772 B.n683 B.n51 163.367
R773 B.n683 B.n682 163.367
R774 B.n682 B.n681 163.367
R775 B.n681 B.n55 163.367
R776 B.n677 B.n55 163.367
R777 B.n677 B.n676 163.367
R778 B.n676 B.n675 163.367
R779 B.n675 B.n57 163.367
R780 B.n670 B.n57 163.367
R781 B.n670 B.n669 163.367
R782 B.n669 B.n668 163.367
R783 B.n668 B.n61 163.367
R784 B.n664 B.n61 163.367
R785 B.n664 B.n663 163.367
R786 B.n663 B.n662 163.367
R787 B.n662 B.n63 163.367
R788 B.n658 B.n63 163.367
R789 B.n658 B.n657 163.367
R790 B.n657 B.n656 163.367
R791 B.n656 B.n65 163.367
R792 B.n652 B.n65 163.367
R793 B.n652 B.n651 163.367
R794 B.n651 B.n650 163.367
R795 B.n650 B.n67 163.367
R796 B.n646 B.n67 163.367
R797 B.n646 B.n645 163.367
R798 B.n645 B.n644 163.367
R799 B.n644 B.n69 163.367
R800 B.n640 B.n69 163.367
R801 B.n640 B.n639 163.367
R802 B.n639 B.n638 163.367
R803 B.n638 B.n71 163.367
R804 B.n634 B.n71 163.367
R805 B.n634 B.n633 163.367
R806 B.n633 B.n632 163.367
R807 B.n632 B.n73 163.367
R808 B.n628 B.n73 163.367
R809 B.n628 B.n627 163.367
R810 B.n627 B.n626 163.367
R811 B.n626 B.n75 163.367
R812 B.n622 B.n75 163.367
R813 B.n622 B.n621 163.367
R814 B.n621 B.n620 163.367
R815 B.n620 B.n77 163.367
R816 B.n616 B.n77 163.367
R817 B.n616 B.n615 163.367
R818 B.n615 B.n614 163.367
R819 B.n614 B.n79 163.367
R820 B.n610 B.n79 163.367
R821 B.n610 B.n609 163.367
R822 B.n609 B.n608 163.367
R823 B.n608 B.n81 163.367
R824 B.n604 B.n81 163.367
R825 B.n604 B.n603 163.367
R826 B.n603 B.n602 163.367
R827 B.n602 B.n83 163.367
R828 B.n598 B.n83 163.367
R829 B.n598 B.n597 163.367
R830 B.n597 B.n596 163.367
R831 B.n596 B.n85 163.367
R832 B.n592 B.n85 163.367
R833 B.n592 B.n591 163.367
R834 B.n591 B.n590 163.367
R835 B.n590 B.n87 163.367
R836 B.n159 B.n158 74.4732
R837 B.n167 B.n166 74.4732
R838 B.n53 B.n52 74.4732
R839 B.n59 B.n58 74.4732
R840 B.n160 B.n159 59.5399
R841 B.n361 B.n167 59.5399
R842 B.n686 B.n53 59.5399
R843 B.n672 B.n59 59.5399
R844 B.n771 B.n770 32.3127
R845 B.n588 B.n587 32.3127
R846 B.n461 B.n130 32.3127
R847 B.n277 B.n276 32.3127
R848 B B.n835 18.0485
R849 B.n770 B.n769 10.6151
R850 B.n769 B.n24 10.6151
R851 B.n765 B.n24 10.6151
R852 B.n765 B.n764 10.6151
R853 B.n764 B.n763 10.6151
R854 B.n763 B.n26 10.6151
R855 B.n759 B.n26 10.6151
R856 B.n759 B.n758 10.6151
R857 B.n758 B.n757 10.6151
R858 B.n757 B.n28 10.6151
R859 B.n753 B.n28 10.6151
R860 B.n753 B.n752 10.6151
R861 B.n752 B.n751 10.6151
R862 B.n751 B.n30 10.6151
R863 B.n747 B.n30 10.6151
R864 B.n747 B.n746 10.6151
R865 B.n746 B.n745 10.6151
R866 B.n745 B.n32 10.6151
R867 B.n741 B.n32 10.6151
R868 B.n741 B.n740 10.6151
R869 B.n740 B.n739 10.6151
R870 B.n739 B.n34 10.6151
R871 B.n735 B.n34 10.6151
R872 B.n735 B.n734 10.6151
R873 B.n734 B.n733 10.6151
R874 B.n733 B.n36 10.6151
R875 B.n729 B.n36 10.6151
R876 B.n729 B.n728 10.6151
R877 B.n728 B.n727 10.6151
R878 B.n727 B.n38 10.6151
R879 B.n723 B.n38 10.6151
R880 B.n723 B.n722 10.6151
R881 B.n722 B.n721 10.6151
R882 B.n721 B.n40 10.6151
R883 B.n717 B.n40 10.6151
R884 B.n717 B.n716 10.6151
R885 B.n716 B.n715 10.6151
R886 B.n715 B.n42 10.6151
R887 B.n711 B.n42 10.6151
R888 B.n711 B.n710 10.6151
R889 B.n710 B.n709 10.6151
R890 B.n709 B.n44 10.6151
R891 B.n705 B.n44 10.6151
R892 B.n705 B.n704 10.6151
R893 B.n704 B.n703 10.6151
R894 B.n703 B.n46 10.6151
R895 B.n699 B.n46 10.6151
R896 B.n699 B.n698 10.6151
R897 B.n698 B.n697 10.6151
R898 B.n697 B.n48 10.6151
R899 B.n693 B.n48 10.6151
R900 B.n693 B.n692 10.6151
R901 B.n692 B.n691 10.6151
R902 B.n691 B.n50 10.6151
R903 B.n687 B.n50 10.6151
R904 B.n685 B.n684 10.6151
R905 B.n684 B.n54 10.6151
R906 B.n680 B.n54 10.6151
R907 B.n680 B.n679 10.6151
R908 B.n679 B.n678 10.6151
R909 B.n678 B.n56 10.6151
R910 B.n674 B.n56 10.6151
R911 B.n674 B.n673 10.6151
R912 B.n671 B.n60 10.6151
R913 B.n667 B.n60 10.6151
R914 B.n667 B.n666 10.6151
R915 B.n666 B.n665 10.6151
R916 B.n665 B.n62 10.6151
R917 B.n661 B.n62 10.6151
R918 B.n661 B.n660 10.6151
R919 B.n660 B.n659 10.6151
R920 B.n659 B.n64 10.6151
R921 B.n655 B.n64 10.6151
R922 B.n655 B.n654 10.6151
R923 B.n654 B.n653 10.6151
R924 B.n653 B.n66 10.6151
R925 B.n649 B.n66 10.6151
R926 B.n649 B.n648 10.6151
R927 B.n648 B.n647 10.6151
R928 B.n647 B.n68 10.6151
R929 B.n643 B.n68 10.6151
R930 B.n643 B.n642 10.6151
R931 B.n642 B.n641 10.6151
R932 B.n641 B.n70 10.6151
R933 B.n637 B.n70 10.6151
R934 B.n637 B.n636 10.6151
R935 B.n636 B.n635 10.6151
R936 B.n635 B.n72 10.6151
R937 B.n631 B.n72 10.6151
R938 B.n631 B.n630 10.6151
R939 B.n630 B.n629 10.6151
R940 B.n629 B.n74 10.6151
R941 B.n625 B.n74 10.6151
R942 B.n625 B.n624 10.6151
R943 B.n624 B.n623 10.6151
R944 B.n623 B.n76 10.6151
R945 B.n619 B.n76 10.6151
R946 B.n619 B.n618 10.6151
R947 B.n618 B.n617 10.6151
R948 B.n617 B.n78 10.6151
R949 B.n613 B.n78 10.6151
R950 B.n613 B.n612 10.6151
R951 B.n612 B.n611 10.6151
R952 B.n611 B.n80 10.6151
R953 B.n607 B.n80 10.6151
R954 B.n607 B.n606 10.6151
R955 B.n606 B.n605 10.6151
R956 B.n605 B.n82 10.6151
R957 B.n601 B.n82 10.6151
R958 B.n601 B.n600 10.6151
R959 B.n600 B.n599 10.6151
R960 B.n599 B.n84 10.6151
R961 B.n595 B.n84 10.6151
R962 B.n595 B.n594 10.6151
R963 B.n594 B.n593 10.6151
R964 B.n593 B.n86 10.6151
R965 B.n589 B.n86 10.6151
R966 B.n589 B.n588 10.6151
R967 B.n462 B.n461 10.6151
R968 B.n463 B.n462 10.6151
R969 B.n463 B.n128 10.6151
R970 B.n467 B.n128 10.6151
R971 B.n468 B.n467 10.6151
R972 B.n469 B.n468 10.6151
R973 B.n469 B.n126 10.6151
R974 B.n473 B.n126 10.6151
R975 B.n474 B.n473 10.6151
R976 B.n475 B.n474 10.6151
R977 B.n475 B.n124 10.6151
R978 B.n479 B.n124 10.6151
R979 B.n480 B.n479 10.6151
R980 B.n481 B.n480 10.6151
R981 B.n481 B.n122 10.6151
R982 B.n485 B.n122 10.6151
R983 B.n486 B.n485 10.6151
R984 B.n487 B.n486 10.6151
R985 B.n487 B.n120 10.6151
R986 B.n491 B.n120 10.6151
R987 B.n492 B.n491 10.6151
R988 B.n493 B.n492 10.6151
R989 B.n493 B.n118 10.6151
R990 B.n497 B.n118 10.6151
R991 B.n498 B.n497 10.6151
R992 B.n499 B.n498 10.6151
R993 B.n499 B.n116 10.6151
R994 B.n503 B.n116 10.6151
R995 B.n504 B.n503 10.6151
R996 B.n505 B.n504 10.6151
R997 B.n505 B.n114 10.6151
R998 B.n509 B.n114 10.6151
R999 B.n510 B.n509 10.6151
R1000 B.n511 B.n510 10.6151
R1001 B.n511 B.n112 10.6151
R1002 B.n515 B.n112 10.6151
R1003 B.n516 B.n515 10.6151
R1004 B.n517 B.n516 10.6151
R1005 B.n517 B.n110 10.6151
R1006 B.n521 B.n110 10.6151
R1007 B.n522 B.n521 10.6151
R1008 B.n523 B.n522 10.6151
R1009 B.n523 B.n108 10.6151
R1010 B.n527 B.n108 10.6151
R1011 B.n528 B.n527 10.6151
R1012 B.n529 B.n528 10.6151
R1013 B.n529 B.n106 10.6151
R1014 B.n533 B.n106 10.6151
R1015 B.n534 B.n533 10.6151
R1016 B.n535 B.n534 10.6151
R1017 B.n535 B.n104 10.6151
R1018 B.n539 B.n104 10.6151
R1019 B.n540 B.n539 10.6151
R1020 B.n541 B.n540 10.6151
R1021 B.n541 B.n102 10.6151
R1022 B.n545 B.n102 10.6151
R1023 B.n546 B.n545 10.6151
R1024 B.n547 B.n546 10.6151
R1025 B.n547 B.n100 10.6151
R1026 B.n551 B.n100 10.6151
R1027 B.n552 B.n551 10.6151
R1028 B.n553 B.n552 10.6151
R1029 B.n553 B.n98 10.6151
R1030 B.n557 B.n98 10.6151
R1031 B.n558 B.n557 10.6151
R1032 B.n559 B.n558 10.6151
R1033 B.n559 B.n96 10.6151
R1034 B.n563 B.n96 10.6151
R1035 B.n564 B.n563 10.6151
R1036 B.n565 B.n564 10.6151
R1037 B.n565 B.n94 10.6151
R1038 B.n569 B.n94 10.6151
R1039 B.n570 B.n569 10.6151
R1040 B.n571 B.n570 10.6151
R1041 B.n571 B.n92 10.6151
R1042 B.n575 B.n92 10.6151
R1043 B.n576 B.n575 10.6151
R1044 B.n577 B.n576 10.6151
R1045 B.n577 B.n90 10.6151
R1046 B.n581 B.n90 10.6151
R1047 B.n582 B.n581 10.6151
R1048 B.n583 B.n582 10.6151
R1049 B.n583 B.n88 10.6151
R1050 B.n587 B.n88 10.6151
R1051 B.n277 B.n194 10.6151
R1052 B.n281 B.n194 10.6151
R1053 B.n282 B.n281 10.6151
R1054 B.n283 B.n282 10.6151
R1055 B.n283 B.n192 10.6151
R1056 B.n287 B.n192 10.6151
R1057 B.n288 B.n287 10.6151
R1058 B.n289 B.n288 10.6151
R1059 B.n289 B.n190 10.6151
R1060 B.n293 B.n190 10.6151
R1061 B.n294 B.n293 10.6151
R1062 B.n295 B.n294 10.6151
R1063 B.n295 B.n188 10.6151
R1064 B.n299 B.n188 10.6151
R1065 B.n300 B.n299 10.6151
R1066 B.n301 B.n300 10.6151
R1067 B.n301 B.n186 10.6151
R1068 B.n305 B.n186 10.6151
R1069 B.n306 B.n305 10.6151
R1070 B.n307 B.n306 10.6151
R1071 B.n307 B.n184 10.6151
R1072 B.n311 B.n184 10.6151
R1073 B.n312 B.n311 10.6151
R1074 B.n313 B.n312 10.6151
R1075 B.n313 B.n182 10.6151
R1076 B.n317 B.n182 10.6151
R1077 B.n318 B.n317 10.6151
R1078 B.n319 B.n318 10.6151
R1079 B.n319 B.n180 10.6151
R1080 B.n323 B.n180 10.6151
R1081 B.n324 B.n323 10.6151
R1082 B.n325 B.n324 10.6151
R1083 B.n325 B.n178 10.6151
R1084 B.n329 B.n178 10.6151
R1085 B.n330 B.n329 10.6151
R1086 B.n331 B.n330 10.6151
R1087 B.n331 B.n176 10.6151
R1088 B.n335 B.n176 10.6151
R1089 B.n336 B.n335 10.6151
R1090 B.n337 B.n336 10.6151
R1091 B.n337 B.n174 10.6151
R1092 B.n341 B.n174 10.6151
R1093 B.n342 B.n341 10.6151
R1094 B.n343 B.n342 10.6151
R1095 B.n343 B.n172 10.6151
R1096 B.n347 B.n172 10.6151
R1097 B.n348 B.n347 10.6151
R1098 B.n349 B.n348 10.6151
R1099 B.n349 B.n170 10.6151
R1100 B.n353 B.n170 10.6151
R1101 B.n354 B.n353 10.6151
R1102 B.n355 B.n354 10.6151
R1103 B.n355 B.n168 10.6151
R1104 B.n359 B.n168 10.6151
R1105 B.n360 B.n359 10.6151
R1106 B.n362 B.n164 10.6151
R1107 B.n366 B.n164 10.6151
R1108 B.n367 B.n366 10.6151
R1109 B.n368 B.n367 10.6151
R1110 B.n368 B.n162 10.6151
R1111 B.n372 B.n162 10.6151
R1112 B.n373 B.n372 10.6151
R1113 B.n374 B.n373 10.6151
R1114 B.n378 B.n377 10.6151
R1115 B.n379 B.n378 10.6151
R1116 B.n379 B.n156 10.6151
R1117 B.n383 B.n156 10.6151
R1118 B.n384 B.n383 10.6151
R1119 B.n385 B.n384 10.6151
R1120 B.n385 B.n154 10.6151
R1121 B.n389 B.n154 10.6151
R1122 B.n390 B.n389 10.6151
R1123 B.n391 B.n390 10.6151
R1124 B.n391 B.n152 10.6151
R1125 B.n395 B.n152 10.6151
R1126 B.n396 B.n395 10.6151
R1127 B.n397 B.n396 10.6151
R1128 B.n397 B.n150 10.6151
R1129 B.n401 B.n150 10.6151
R1130 B.n402 B.n401 10.6151
R1131 B.n403 B.n402 10.6151
R1132 B.n403 B.n148 10.6151
R1133 B.n407 B.n148 10.6151
R1134 B.n408 B.n407 10.6151
R1135 B.n409 B.n408 10.6151
R1136 B.n409 B.n146 10.6151
R1137 B.n413 B.n146 10.6151
R1138 B.n414 B.n413 10.6151
R1139 B.n415 B.n414 10.6151
R1140 B.n415 B.n144 10.6151
R1141 B.n419 B.n144 10.6151
R1142 B.n420 B.n419 10.6151
R1143 B.n421 B.n420 10.6151
R1144 B.n421 B.n142 10.6151
R1145 B.n425 B.n142 10.6151
R1146 B.n426 B.n425 10.6151
R1147 B.n427 B.n426 10.6151
R1148 B.n427 B.n140 10.6151
R1149 B.n431 B.n140 10.6151
R1150 B.n432 B.n431 10.6151
R1151 B.n433 B.n432 10.6151
R1152 B.n433 B.n138 10.6151
R1153 B.n437 B.n138 10.6151
R1154 B.n438 B.n437 10.6151
R1155 B.n439 B.n438 10.6151
R1156 B.n439 B.n136 10.6151
R1157 B.n443 B.n136 10.6151
R1158 B.n444 B.n443 10.6151
R1159 B.n445 B.n444 10.6151
R1160 B.n445 B.n134 10.6151
R1161 B.n449 B.n134 10.6151
R1162 B.n450 B.n449 10.6151
R1163 B.n451 B.n450 10.6151
R1164 B.n451 B.n132 10.6151
R1165 B.n455 B.n132 10.6151
R1166 B.n456 B.n455 10.6151
R1167 B.n457 B.n456 10.6151
R1168 B.n457 B.n130 10.6151
R1169 B.n276 B.n275 10.6151
R1170 B.n275 B.n196 10.6151
R1171 B.n271 B.n196 10.6151
R1172 B.n271 B.n270 10.6151
R1173 B.n270 B.n269 10.6151
R1174 B.n269 B.n198 10.6151
R1175 B.n265 B.n198 10.6151
R1176 B.n265 B.n264 10.6151
R1177 B.n264 B.n263 10.6151
R1178 B.n263 B.n200 10.6151
R1179 B.n259 B.n200 10.6151
R1180 B.n259 B.n258 10.6151
R1181 B.n258 B.n257 10.6151
R1182 B.n257 B.n202 10.6151
R1183 B.n253 B.n202 10.6151
R1184 B.n253 B.n252 10.6151
R1185 B.n252 B.n251 10.6151
R1186 B.n251 B.n204 10.6151
R1187 B.n247 B.n204 10.6151
R1188 B.n247 B.n246 10.6151
R1189 B.n246 B.n245 10.6151
R1190 B.n245 B.n206 10.6151
R1191 B.n241 B.n206 10.6151
R1192 B.n241 B.n240 10.6151
R1193 B.n240 B.n239 10.6151
R1194 B.n239 B.n208 10.6151
R1195 B.n235 B.n208 10.6151
R1196 B.n235 B.n234 10.6151
R1197 B.n234 B.n233 10.6151
R1198 B.n233 B.n210 10.6151
R1199 B.n229 B.n210 10.6151
R1200 B.n229 B.n228 10.6151
R1201 B.n228 B.n227 10.6151
R1202 B.n227 B.n212 10.6151
R1203 B.n223 B.n212 10.6151
R1204 B.n223 B.n222 10.6151
R1205 B.n222 B.n221 10.6151
R1206 B.n221 B.n214 10.6151
R1207 B.n217 B.n214 10.6151
R1208 B.n217 B.n216 10.6151
R1209 B.n216 B.n0 10.6151
R1210 B.n831 B.n1 10.6151
R1211 B.n831 B.n830 10.6151
R1212 B.n830 B.n829 10.6151
R1213 B.n829 B.n4 10.6151
R1214 B.n825 B.n4 10.6151
R1215 B.n825 B.n824 10.6151
R1216 B.n824 B.n823 10.6151
R1217 B.n823 B.n6 10.6151
R1218 B.n819 B.n6 10.6151
R1219 B.n819 B.n818 10.6151
R1220 B.n818 B.n817 10.6151
R1221 B.n817 B.n8 10.6151
R1222 B.n813 B.n8 10.6151
R1223 B.n813 B.n812 10.6151
R1224 B.n812 B.n811 10.6151
R1225 B.n811 B.n10 10.6151
R1226 B.n807 B.n10 10.6151
R1227 B.n807 B.n806 10.6151
R1228 B.n806 B.n805 10.6151
R1229 B.n805 B.n12 10.6151
R1230 B.n801 B.n12 10.6151
R1231 B.n801 B.n800 10.6151
R1232 B.n800 B.n799 10.6151
R1233 B.n799 B.n14 10.6151
R1234 B.n795 B.n14 10.6151
R1235 B.n795 B.n794 10.6151
R1236 B.n794 B.n793 10.6151
R1237 B.n793 B.n16 10.6151
R1238 B.n789 B.n16 10.6151
R1239 B.n789 B.n788 10.6151
R1240 B.n788 B.n787 10.6151
R1241 B.n787 B.n18 10.6151
R1242 B.n783 B.n18 10.6151
R1243 B.n783 B.n782 10.6151
R1244 B.n782 B.n781 10.6151
R1245 B.n781 B.n20 10.6151
R1246 B.n777 B.n20 10.6151
R1247 B.n777 B.n776 10.6151
R1248 B.n776 B.n775 10.6151
R1249 B.n775 B.n22 10.6151
R1250 B.n771 B.n22 10.6151
R1251 B.n686 B.n685 6.5566
R1252 B.n673 B.n672 6.5566
R1253 B.n362 B.n361 6.5566
R1254 B.n374 B.n160 6.5566
R1255 B.n687 B.n686 4.05904
R1256 B.n672 B.n671 4.05904
R1257 B.n361 B.n360 4.05904
R1258 B.n377 B.n160 4.05904
R1259 B.n835 B.n0 2.81026
R1260 B.n835 B.n1 2.81026
R1261 VP.n19 VP.n18 161.3
R1262 VP.n17 VP.n1 161.3
R1263 VP.n16 VP.n15 161.3
R1264 VP.n14 VP.n2 161.3
R1265 VP.n13 VP.n12 161.3
R1266 VP.n11 VP.n3 161.3
R1267 VP.n10 VP.n9 161.3
R1268 VP.n8 VP.n4 161.3
R1269 VP.n5 VP.t2 149.768
R1270 VP.n5 VP.t1 148.547
R1271 VP.n6 VP.t3 115.282
R1272 VP.n0 VP.t0 115.282
R1273 VP.n7 VP.n6 81.7486
R1274 VP.n20 VP.n0 81.7486
R1275 VP.n12 VP.n2 56.5193
R1276 VP.n7 VP.n5 54.9532
R1277 VP.n10 VP.n4 24.4675
R1278 VP.n11 VP.n10 24.4675
R1279 VP.n12 VP.n11 24.4675
R1280 VP.n16 VP.n2 24.4675
R1281 VP.n17 VP.n16 24.4675
R1282 VP.n18 VP.n17 24.4675
R1283 VP.n6 VP.n4 8.31928
R1284 VP.n18 VP.n0 8.31928
R1285 VP.n8 VP.n7 0.354971
R1286 VP.n20 VP.n19 0.354971
R1287 VP VP.n20 0.26696
R1288 VP.n9 VP.n8 0.189894
R1289 VP.n9 VP.n3 0.189894
R1290 VP.n13 VP.n3 0.189894
R1291 VP.n14 VP.n13 0.189894
R1292 VP.n15 VP.n14 0.189894
R1293 VP.n15 VP.n1 0.189894
R1294 VP.n19 VP.n1 0.189894
R1295 VTAIL.n746 VTAIL.n658 756.745
R1296 VTAIL.n88 VTAIL.n0 756.745
R1297 VTAIL.n182 VTAIL.n94 756.745
R1298 VTAIL.n276 VTAIL.n188 756.745
R1299 VTAIL.n652 VTAIL.n564 756.745
R1300 VTAIL.n558 VTAIL.n470 756.745
R1301 VTAIL.n464 VTAIL.n376 756.745
R1302 VTAIL.n370 VTAIL.n282 756.745
R1303 VTAIL.n689 VTAIL.n688 585
R1304 VTAIL.n686 VTAIL.n685 585
R1305 VTAIL.n695 VTAIL.n694 585
R1306 VTAIL.n697 VTAIL.n696 585
R1307 VTAIL.n682 VTAIL.n681 585
R1308 VTAIL.n703 VTAIL.n702 585
R1309 VTAIL.n705 VTAIL.n704 585
R1310 VTAIL.n678 VTAIL.n677 585
R1311 VTAIL.n711 VTAIL.n710 585
R1312 VTAIL.n713 VTAIL.n712 585
R1313 VTAIL.n674 VTAIL.n673 585
R1314 VTAIL.n719 VTAIL.n718 585
R1315 VTAIL.n721 VTAIL.n720 585
R1316 VTAIL.n670 VTAIL.n669 585
R1317 VTAIL.n727 VTAIL.n726 585
R1318 VTAIL.n730 VTAIL.n729 585
R1319 VTAIL.n728 VTAIL.n666 585
R1320 VTAIL.n735 VTAIL.n665 585
R1321 VTAIL.n737 VTAIL.n736 585
R1322 VTAIL.n739 VTAIL.n738 585
R1323 VTAIL.n662 VTAIL.n661 585
R1324 VTAIL.n745 VTAIL.n744 585
R1325 VTAIL.n747 VTAIL.n746 585
R1326 VTAIL.n31 VTAIL.n30 585
R1327 VTAIL.n28 VTAIL.n27 585
R1328 VTAIL.n37 VTAIL.n36 585
R1329 VTAIL.n39 VTAIL.n38 585
R1330 VTAIL.n24 VTAIL.n23 585
R1331 VTAIL.n45 VTAIL.n44 585
R1332 VTAIL.n47 VTAIL.n46 585
R1333 VTAIL.n20 VTAIL.n19 585
R1334 VTAIL.n53 VTAIL.n52 585
R1335 VTAIL.n55 VTAIL.n54 585
R1336 VTAIL.n16 VTAIL.n15 585
R1337 VTAIL.n61 VTAIL.n60 585
R1338 VTAIL.n63 VTAIL.n62 585
R1339 VTAIL.n12 VTAIL.n11 585
R1340 VTAIL.n69 VTAIL.n68 585
R1341 VTAIL.n72 VTAIL.n71 585
R1342 VTAIL.n70 VTAIL.n8 585
R1343 VTAIL.n77 VTAIL.n7 585
R1344 VTAIL.n79 VTAIL.n78 585
R1345 VTAIL.n81 VTAIL.n80 585
R1346 VTAIL.n4 VTAIL.n3 585
R1347 VTAIL.n87 VTAIL.n86 585
R1348 VTAIL.n89 VTAIL.n88 585
R1349 VTAIL.n125 VTAIL.n124 585
R1350 VTAIL.n122 VTAIL.n121 585
R1351 VTAIL.n131 VTAIL.n130 585
R1352 VTAIL.n133 VTAIL.n132 585
R1353 VTAIL.n118 VTAIL.n117 585
R1354 VTAIL.n139 VTAIL.n138 585
R1355 VTAIL.n141 VTAIL.n140 585
R1356 VTAIL.n114 VTAIL.n113 585
R1357 VTAIL.n147 VTAIL.n146 585
R1358 VTAIL.n149 VTAIL.n148 585
R1359 VTAIL.n110 VTAIL.n109 585
R1360 VTAIL.n155 VTAIL.n154 585
R1361 VTAIL.n157 VTAIL.n156 585
R1362 VTAIL.n106 VTAIL.n105 585
R1363 VTAIL.n163 VTAIL.n162 585
R1364 VTAIL.n166 VTAIL.n165 585
R1365 VTAIL.n164 VTAIL.n102 585
R1366 VTAIL.n171 VTAIL.n101 585
R1367 VTAIL.n173 VTAIL.n172 585
R1368 VTAIL.n175 VTAIL.n174 585
R1369 VTAIL.n98 VTAIL.n97 585
R1370 VTAIL.n181 VTAIL.n180 585
R1371 VTAIL.n183 VTAIL.n182 585
R1372 VTAIL.n219 VTAIL.n218 585
R1373 VTAIL.n216 VTAIL.n215 585
R1374 VTAIL.n225 VTAIL.n224 585
R1375 VTAIL.n227 VTAIL.n226 585
R1376 VTAIL.n212 VTAIL.n211 585
R1377 VTAIL.n233 VTAIL.n232 585
R1378 VTAIL.n235 VTAIL.n234 585
R1379 VTAIL.n208 VTAIL.n207 585
R1380 VTAIL.n241 VTAIL.n240 585
R1381 VTAIL.n243 VTAIL.n242 585
R1382 VTAIL.n204 VTAIL.n203 585
R1383 VTAIL.n249 VTAIL.n248 585
R1384 VTAIL.n251 VTAIL.n250 585
R1385 VTAIL.n200 VTAIL.n199 585
R1386 VTAIL.n257 VTAIL.n256 585
R1387 VTAIL.n260 VTAIL.n259 585
R1388 VTAIL.n258 VTAIL.n196 585
R1389 VTAIL.n265 VTAIL.n195 585
R1390 VTAIL.n267 VTAIL.n266 585
R1391 VTAIL.n269 VTAIL.n268 585
R1392 VTAIL.n192 VTAIL.n191 585
R1393 VTAIL.n275 VTAIL.n274 585
R1394 VTAIL.n277 VTAIL.n276 585
R1395 VTAIL.n653 VTAIL.n652 585
R1396 VTAIL.n651 VTAIL.n650 585
R1397 VTAIL.n568 VTAIL.n567 585
R1398 VTAIL.n645 VTAIL.n644 585
R1399 VTAIL.n643 VTAIL.n642 585
R1400 VTAIL.n641 VTAIL.n571 585
R1401 VTAIL.n575 VTAIL.n572 585
R1402 VTAIL.n636 VTAIL.n635 585
R1403 VTAIL.n634 VTAIL.n633 585
R1404 VTAIL.n577 VTAIL.n576 585
R1405 VTAIL.n628 VTAIL.n627 585
R1406 VTAIL.n626 VTAIL.n625 585
R1407 VTAIL.n581 VTAIL.n580 585
R1408 VTAIL.n620 VTAIL.n619 585
R1409 VTAIL.n618 VTAIL.n617 585
R1410 VTAIL.n585 VTAIL.n584 585
R1411 VTAIL.n612 VTAIL.n611 585
R1412 VTAIL.n610 VTAIL.n609 585
R1413 VTAIL.n589 VTAIL.n588 585
R1414 VTAIL.n604 VTAIL.n603 585
R1415 VTAIL.n602 VTAIL.n601 585
R1416 VTAIL.n593 VTAIL.n592 585
R1417 VTAIL.n596 VTAIL.n595 585
R1418 VTAIL.n559 VTAIL.n558 585
R1419 VTAIL.n557 VTAIL.n556 585
R1420 VTAIL.n474 VTAIL.n473 585
R1421 VTAIL.n551 VTAIL.n550 585
R1422 VTAIL.n549 VTAIL.n548 585
R1423 VTAIL.n547 VTAIL.n477 585
R1424 VTAIL.n481 VTAIL.n478 585
R1425 VTAIL.n542 VTAIL.n541 585
R1426 VTAIL.n540 VTAIL.n539 585
R1427 VTAIL.n483 VTAIL.n482 585
R1428 VTAIL.n534 VTAIL.n533 585
R1429 VTAIL.n532 VTAIL.n531 585
R1430 VTAIL.n487 VTAIL.n486 585
R1431 VTAIL.n526 VTAIL.n525 585
R1432 VTAIL.n524 VTAIL.n523 585
R1433 VTAIL.n491 VTAIL.n490 585
R1434 VTAIL.n518 VTAIL.n517 585
R1435 VTAIL.n516 VTAIL.n515 585
R1436 VTAIL.n495 VTAIL.n494 585
R1437 VTAIL.n510 VTAIL.n509 585
R1438 VTAIL.n508 VTAIL.n507 585
R1439 VTAIL.n499 VTAIL.n498 585
R1440 VTAIL.n502 VTAIL.n501 585
R1441 VTAIL.n465 VTAIL.n464 585
R1442 VTAIL.n463 VTAIL.n462 585
R1443 VTAIL.n380 VTAIL.n379 585
R1444 VTAIL.n457 VTAIL.n456 585
R1445 VTAIL.n455 VTAIL.n454 585
R1446 VTAIL.n453 VTAIL.n383 585
R1447 VTAIL.n387 VTAIL.n384 585
R1448 VTAIL.n448 VTAIL.n447 585
R1449 VTAIL.n446 VTAIL.n445 585
R1450 VTAIL.n389 VTAIL.n388 585
R1451 VTAIL.n440 VTAIL.n439 585
R1452 VTAIL.n438 VTAIL.n437 585
R1453 VTAIL.n393 VTAIL.n392 585
R1454 VTAIL.n432 VTAIL.n431 585
R1455 VTAIL.n430 VTAIL.n429 585
R1456 VTAIL.n397 VTAIL.n396 585
R1457 VTAIL.n424 VTAIL.n423 585
R1458 VTAIL.n422 VTAIL.n421 585
R1459 VTAIL.n401 VTAIL.n400 585
R1460 VTAIL.n416 VTAIL.n415 585
R1461 VTAIL.n414 VTAIL.n413 585
R1462 VTAIL.n405 VTAIL.n404 585
R1463 VTAIL.n408 VTAIL.n407 585
R1464 VTAIL.n371 VTAIL.n370 585
R1465 VTAIL.n369 VTAIL.n368 585
R1466 VTAIL.n286 VTAIL.n285 585
R1467 VTAIL.n363 VTAIL.n362 585
R1468 VTAIL.n361 VTAIL.n360 585
R1469 VTAIL.n359 VTAIL.n289 585
R1470 VTAIL.n293 VTAIL.n290 585
R1471 VTAIL.n354 VTAIL.n353 585
R1472 VTAIL.n352 VTAIL.n351 585
R1473 VTAIL.n295 VTAIL.n294 585
R1474 VTAIL.n346 VTAIL.n345 585
R1475 VTAIL.n344 VTAIL.n343 585
R1476 VTAIL.n299 VTAIL.n298 585
R1477 VTAIL.n338 VTAIL.n337 585
R1478 VTAIL.n336 VTAIL.n335 585
R1479 VTAIL.n303 VTAIL.n302 585
R1480 VTAIL.n330 VTAIL.n329 585
R1481 VTAIL.n328 VTAIL.n327 585
R1482 VTAIL.n307 VTAIL.n306 585
R1483 VTAIL.n322 VTAIL.n321 585
R1484 VTAIL.n320 VTAIL.n319 585
R1485 VTAIL.n311 VTAIL.n310 585
R1486 VTAIL.n314 VTAIL.n313 585
R1487 VTAIL.t7 VTAIL.n594 327.466
R1488 VTAIL.t6 VTAIL.n500 327.466
R1489 VTAIL.t3 VTAIL.n406 327.466
R1490 VTAIL.t1 VTAIL.n312 327.466
R1491 VTAIL.t0 VTAIL.n687 327.466
R1492 VTAIL.t2 VTAIL.n29 327.466
R1493 VTAIL.t5 VTAIL.n123 327.466
R1494 VTAIL.t4 VTAIL.n217 327.466
R1495 VTAIL.n688 VTAIL.n685 171.744
R1496 VTAIL.n695 VTAIL.n685 171.744
R1497 VTAIL.n696 VTAIL.n695 171.744
R1498 VTAIL.n696 VTAIL.n681 171.744
R1499 VTAIL.n703 VTAIL.n681 171.744
R1500 VTAIL.n704 VTAIL.n703 171.744
R1501 VTAIL.n704 VTAIL.n677 171.744
R1502 VTAIL.n711 VTAIL.n677 171.744
R1503 VTAIL.n712 VTAIL.n711 171.744
R1504 VTAIL.n712 VTAIL.n673 171.744
R1505 VTAIL.n719 VTAIL.n673 171.744
R1506 VTAIL.n720 VTAIL.n719 171.744
R1507 VTAIL.n720 VTAIL.n669 171.744
R1508 VTAIL.n727 VTAIL.n669 171.744
R1509 VTAIL.n729 VTAIL.n727 171.744
R1510 VTAIL.n729 VTAIL.n728 171.744
R1511 VTAIL.n728 VTAIL.n665 171.744
R1512 VTAIL.n737 VTAIL.n665 171.744
R1513 VTAIL.n738 VTAIL.n737 171.744
R1514 VTAIL.n738 VTAIL.n661 171.744
R1515 VTAIL.n745 VTAIL.n661 171.744
R1516 VTAIL.n746 VTAIL.n745 171.744
R1517 VTAIL.n30 VTAIL.n27 171.744
R1518 VTAIL.n37 VTAIL.n27 171.744
R1519 VTAIL.n38 VTAIL.n37 171.744
R1520 VTAIL.n38 VTAIL.n23 171.744
R1521 VTAIL.n45 VTAIL.n23 171.744
R1522 VTAIL.n46 VTAIL.n45 171.744
R1523 VTAIL.n46 VTAIL.n19 171.744
R1524 VTAIL.n53 VTAIL.n19 171.744
R1525 VTAIL.n54 VTAIL.n53 171.744
R1526 VTAIL.n54 VTAIL.n15 171.744
R1527 VTAIL.n61 VTAIL.n15 171.744
R1528 VTAIL.n62 VTAIL.n61 171.744
R1529 VTAIL.n62 VTAIL.n11 171.744
R1530 VTAIL.n69 VTAIL.n11 171.744
R1531 VTAIL.n71 VTAIL.n69 171.744
R1532 VTAIL.n71 VTAIL.n70 171.744
R1533 VTAIL.n70 VTAIL.n7 171.744
R1534 VTAIL.n79 VTAIL.n7 171.744
R1535 VTAIL.n80 VTAIL.n79 171.744
R1536 VTAIL.n80 VTAIL.n3 171.744
R1537 VTAIL.n87 VTAIL.n3 171.744
R1538 VTAIL.n88 VTAIL.n87 171.744
R1539 VTAIL.n124 VTAIL.n121 171.744
R1540 VTAIL.n131 VTAIL.n121 171.744
R1541 VTAIL.n132 VTAIL.n131 171.744
R1542 VTAIL.n132 VTAIL.n117 171.744
R1543 VTAIL.n139 VTAIL.n117 171.744
R1544 VTAIL.n140 VTAIL.n139 171.744
R1545 VTAIL.n140 VTAIL.n113 171.744
R1546 VTAIL.n147 VTAIL.n113 171.744
R1547 VTAIL.n148 VTAIL.n147 171.744
R1548 VTAIL.n148 VTAIL.n109 171.744
R1549 VTAIL.n155 VTAIL.n109 171.744
R1550 VTAIL.n156 VTAIL.n155 171.744
R1551 VTAIL.n156 VTAIL.n105 171.744
R1552 VTAIL.n163 VTAIL.n105 171.744
R1553 VTAIL.n165 VTAIL.n163 171.744
R1554 VTAIL.n165 VTAIL.n164 171.744
R1555 VTAIL.n164 VTAIL.n101 171.744
R1556 VTAIL.n173 VTAIL.n101 171.744
R1557 VTAIL.n174 VTAIL.n173 171.744
R1558 VTAIL.n174 VTAIL.n97 171.744
R1559 VTAIL.n181 VTAIL.n97 171.744
R1560 VTAIL.n182 VTAIL.n181 171.744
R1561 VTAIL.n218 VTAIL.n215 171.744
R1562 VTAIL.n225 VTAIL.n215 171.744
R1563 VTAIL.n226 VTAIL.n225 171.744
R1564 VTAIL.n226 VTAIL.n211 171.744
R1565 VTAIL.n233 VTAIL.n211 171.744
R1566 VTAIL.n234 VTAIL.n233 171.744
R1567 VTAIL.n234 VTAIL.n207 171.744
R1568 VTAIL.n241 VTAIL.n207 171.744
R1569 VTAIL.n242 VTAIL.n241 171.744
R1570 VTAIL.n242 VTAIL.n203 171.744
R1571 VTAIL.n249 VTAIL.n203 171.744
R1572 VTAIL.n250 VTAIL.n249 171.744
R1573 VTAIL.n250 VTAIL.n199 171.744
R1574 VTAIL.n257 VTAIL.n199 171.744
R1575 VTAIL.n259 VTAIL.n257 171.744
R1576 VTAIL.n259 VTAIL.n258 171.744
R1577 VTAIL.n258 VTAIL.n195 171.744
R1578 VTAIL.n267 VTAIL.n195 171.744
R1579 VTAIL.n268 VTAIL.n267 171.744
R1580 VTAIL.n268 VTAIL.n191 171.744
R1581 VTAIL.n275 VTAIL.n191 171.744
R1582 VTAIL.n276 VTAIL.n275 171.744
R1583 VTAIL.n652 VTAIL.n651 171.744
R1584 VTAIL.n651 VTAIL.n567 171.744
R1585 VTAIL.n644 VTAIL.n567 171.744
R1586 VTAIL.n644 VTAIL.n643 171.744
R1587 VTAIL.n643 VTAIL.n571 171.744
R1588 VTAIL.n575 VTAIL.n571 171.744
R1589 VTAIL.n635 VTAIL.n575 171.744
R1590 VTAIL.n635 VTAIL.n634 171.744
R1591 VTAIL.n634 VTAIL.n576 171.744
R1592 VTAIL.n627 VTAIL.n576 171.744
R1593 VTAIL.n627 VTAIL.n626 171.744
R1594 VTAIL.n626 VTAIL.n580 171.744
R1595 VTAIL.n619 VTAIL.n580 171.744
R1596 VTAIL.n619 VTAIL.n618 171.744
R1597 VTAIL.n618 VTAIL.n584 171.744
R1598 VTAIL.n611 VTAIL.n584 171.744
R1599 VTAIL.n611 VTAIL.n610 171.744
R1600 VTAIL.n610 VTAIL.n588 171.744
R1601 VTAIL.n603 VTAIL.n588 171.744
R1602 VTAIL.n603 VTAIL.n602 171.744
R1603 VTAIL.n602 VTAIL.n592 171.744
R1604 VTAIL.n595 VTAIL.n592 171.744
R1605 VTAIL.n558 VTAIL.n557 171.744
R1606 VTAIL.n557 VTAIL.n473 171.744
R1607 VTAIL.n550 VTAIL.n473 171.744
R1608 VTAIL.n550 VTAIL.n549 171.744
R1609 VTAIL.n549 VTAIL.n477 171.744
R1610 VTAIL.n481 VTAIL.n477 171.744
R1611 VTAIL.n541 VTAIL.n481 171.744
R1612 VTAIL.n541 VTAIL.n540 171.744
R1613 VTAIL.n540 VTAIL.n482 171.744
R1614 VTAIL.n533 VTAIL.n482 171.744
R1615 VTAIL.n533 VTAIL.n532 171.744
R1616 VTAIL.n532 VTAIL.n486 171.744
R1617 VTAIL.n525 VTAIL.n486 171.744
R1618 VTAIL.n525 VTAIL.n524 171.744
R1619 VTAIL.n524 VTAIL.n490 171.744
R1620 VTAIL.n517 VTAIL.n490 171.744
R1621 VTAIL.n517 VTAIL.n516 171.744
R1622 VTAIL.n516 VTAIL.n494 171.744
R1623 VTAIL.n509 VTAIL.n494 171.744
R1624 VTAIL.n509 VTAIL.n508 171.744
R1625 VTAIL.n508 VTAIL.n498 171.744
R1626 VTAIL.n501 VTAIL.n498 171.744
R1627 VTAIL.n464 VTAIL.n463 171.744
R1628 VTAIL.n463 VTAIL.n379 171.744
R1629 VTAIL.n456 VTAIL.n379 171.744
R1630 VTAIL.n456 VTAIL.n455 171.744
R1631 VTAIL.n455 VTAIL.n383 171.744
R1632 VTAIL.n387 VTAIL.n383 171.744
R1633 VTAIL.n447 VTAIL.n387 171.744
R1634 VTAIL.n447 VTAIL.n446 171.744
R1635 VTAIL.n446 VTAIL.n388 171.744
R1636 VTAIL.n439 VTAIL.n388 171.744
R1637 VTAIL.n439 VTAIL.n438 171.744
R1638 VTAIL.n438 VTAIL.n392 171.744
R1639 VTAIL.n431 VTAIL.n392 171.744
R1640 VTAIL.n431 VTAIL.n430 171.744
R1641 VTAIL.n430 VTAIL.n396 171.744
R1642 VTAIL.n423 VTAIL.n396 171.744
R1643 VTAIL.n423 VTAIL.n422 171.744
R1644 VTAIL.n422 VTAIL.n400 171.744
R1645 VTAIL.n415 VTAIL.n400 171.744
R1646 VTAIL.n415 VTAIL.n414 171.744
R1647 VTAIL.n414 VTAIL.n404 171.744
R1648 VTAIL.n407 VTAIL.n404 171.744
R1649 VTAIL.n370 VTAIL.n369 171.744
R1650 VTAIL.n369 VTAIL.n285 171.744
R1651 VTAIL.n362 VTAIL.n285 171.744
R1652 VTAIL.n362 VTAIL.n361 171.744
R1653 VTAIL.n361 VTAIL.n289 171.744
R1654 VTAIL.n293 VTAIL.n289 171.744
R1655 VTAIL.n353 VTAIL.n293 171.744
R1656 VTAIL.n353 VTAIL.n352 171.744
R1657 VTAIL.n352 VTAIL.n294 171.744
R1658 VTAIL.n345 VTAIL.n294 171.744
R1659 VTAIL.n345 VTAIL.n344 171.744
R1660 VTAIL.n344 VTAIL.n298 171.744
R1661 VTAIL.n337 VTAIL.n298 171.744
R1662 VTAIL.n337 VTAIL.n336 171.744
R1663 VTAIL.n336 VTAIL.n302 171.744
R1664 VTAIL.n329 VTAIL.n302 171.744
R1665 VTAIL.n329 VTAIL.n328 171.744
R1666 VTAIL.n328 VTAIL.n306 171.744
R1667 VTAIL.n321 VTAIL.n306 171.744
R1668 VTAIL.n321 VTAIL.n320 171.744
R1669 VTAIL.n320 VTAIL.n310 171.744
R1670 VTAIL.n313 VTAIL.n310 171.744
R1671 VTAIL.n688 VTAIL.t0 85.8723
R1672 VTAIL.n30 VTAIL.t2 85.8723
R1673 VTAIL.n124 VTAIL.t5 85.8723
R1674 VTAIL.n218 VTAIL.t4 85.8723
R1675 VTAIL.n595 VTAIL.t7 85.8723
R1676 VTAIL.n501 VTAIL.t6 85.8723
R1677 VTAIL.n407 VTAIL.t3 85.8723
R1678 VTAIL.n313 VTAIL.t1 85.8723
R1679 VTAIL.n751 VTAIL.n750 31.9914
R1680 VTAIL.n93 VTAIL.n92 31.9914
R1681 VTAIL.n187 VTAIL.n186 31.9914
R1682 VTAIL.n281 VTAIL.n280 31.9914
R1683 VTAIL.n657 VTAIL.n656 31.9914
R1684 VTAIL.n563 VTAIL.n562 31.9914
R1685 VTAIL.n469 VTAIL.n468 31.9914
R1686 VTAIL.n375 VTAIL.n374 31.9914
R1687 VTAIL.n751 VTAIL.n657 30.1514
R1688 VTAIL.n375 VTAIL.n281 30.1514
R1689 VTAIL.n689 VTAIL.n687 16.3895
R1690 VTAIL.n31 VTAIL.n29 16.3895
R1691 VTAIL.n125 VTAIL.n123 16.3895
R1692 VTAIL.n219 VTAIL.n217 16.3895
R1693 VTAIL.n596 VTAIL.n594 16.3895
R1694 VTAIL.n502 VTAIL.n500 16.3895
R1695 VTAIL.n408 VTAIL.n406 16.3895
R1696 VTAIL.n314 VTAIL.n312 16.3895
R1697 VTAIL.n736 VTAIL.n735 13.1884
R1698 VTAIL.n78 VTAIL.n77 13.1884
R1699 VTAIL.n172 VTAIL.n171 13.1884
R1700 VTAIL.n266 VTAIL.n265 13.1884
R1701 VTAIL.n642 VTAIL.n641 13.1884
R1702 VTAIL.n548 VTAIL.n547 13.1884
R1703 VTAIL.n454 VTAIL.n453 13.1884
R1704 VTAIL.n360 VTAIL.n359 13.1884
R1705 VTAIL.n690 VTAIL.n686 12.8005
R1706 VTAIL.n734 VTAIL.n666 12.8005
R1707 VTAIL.n739 VTAIL.n664 12.8005
R1708 VTAIL.n32 VTAIL.n28 12.8005
R1709 VTAIL.n76 VTAIL.n8 12.8005
R1710 VTAIL.n81 VTAIL.n6 12.8005
R1711 VTAIL.n126 VTAIL.n122 12.8005
R1712 VTAIL.n170 VTAIL.n102 12.8005
R1713 VTAIL.n175 VTAIL.n100 12.8005
R1714 VTAIL.n220 VTAIL.n216 12.8005
R1715 VTAIL.n264 VTAIL.n196 12.8005
R1716 VTAIL.n269 VTAIL.n194 12.8005
R1717 VTAIL.n645 VTAIL.n570 12.8005
R1718 VTAIL.n640 VTAIL.n572 12.8005
R1719 VTAIL.n597 VTAIL.n593 12.8005
R1720 VTAIL.n551 VTAIL.n476 12.8005
R1721 VTAIL.n546 VTAIL.n478 12.8005
R1722 VTAIL.n503 VTAIL.n499 12.8005
R1723 VTAIL.n457 VTAIL.n382 12.8005
R1724 VTAIL.n452 VTAIL.n384 12.8005
R1725 VTAIL.n409 VTAIL.n405 12.8005
R1726 VTAIL.n363 VTAIL.n288 12.8005
R1727 VTAIL.n358 VTAIL.n290 12.8005
R1728 VTAIL.n315 VTAIL.n311 12.8005
R1729 VTAIL.n694 VTAIL.n693 12.0247
R1730 VTAIL.n731 VTAIL.n730 12.0247
R1731 VTAIL.n740 VTAIL.n662 12.0247
R1732 VTAIL.n36 VTAIL.n35 12.0247
R1733 VTAIL.n73 VTAIL.n72 12.0247
R1734 VTAIL.n82 VTAIL.n4 12.0247
R1735 VTAIL.n130 VTAIL.n129 12.0247
R1736 VTAIL.n167 VTAIL.n166 12.0247
R1737 VTAIL.n176 VTAIL.n98 12.0247
R1738 VTAIL.n224 VTAIL.n223 12.0247
R1739 VTAIL.n261 VTAIL.n260 12.0247
R1740 VTAIL.n270 VTAIL.n192 12.0247
R1741 VTAIL.n646 VTAIL.n568 12.0247
R1742 VTAIL.n637 VTAIL.n636 12.0247
R1743 VTAIL.n601 VTAIL.n600 12.0247
R1744 VTAIL.n552 VTAIL.n474 12.0247
R1745 VTAIL.n543 VTAIL.n542 12.0247
R1746 VTAIL.n507 VTAIL.n506 12.0247
R1747 VTAIL.n458 VTAIL.n380 12.0247
R1748 VTAIL.n449 VTAIL.n448 12.0247
R1749 VTAIL.n413 VTAIL.n412 12.0247
R1750 VTAIL.n364 VTAIL.n286 12.0247
R1751 VTAIL.n355 VTAIL.n354 12.0247
R1752 VTAIL.n319 VTAIL.n318 12.0247
R1753 VTAIL.n697 VTAIL.n684 11.249
R1754 VTAIL.n726 VTAIL.n668 11.249
R1755 VTAIL.n744 VTAIL.n743 11.249
R1756 VTAIL.n39 VTAIL.n26 11.249
R1757 VTAIL.n68 VTAIL.n10 11.249
R1758 VTAIL.n86 VTAIL.n85 11.249
R1759 VTAIL.n133 VTAIL.n120 11.249
R1760 VTAIL.n162 VTAIL.n104 11.249
R1761 VTAIL.n180 VTAIL.n179 11.249
R1762 VTAIL.n227 VTAIL.n214 11.249
R1763 VTAIL.n256 VTAIL.n198 11.249
R1764 VTAIL.n274 VTAIL.n273 11.249
R1765 VTAIL.n650 VTAIL.n649 11.249
R1766 VTAIL.n633 VTAIL.n574 11.249
R1767 VTAIL.n604 VTAIL.n591 11.249
R1768 VTAIL.n556 VTAIL.n555 11.249
R1769 VTAIL.n539 VTAIL.n480 11.249
R1770 VTAIL.n510 VTAIL.n497 11.249
R1771 VTAIL.n462 VTAIL.n461 11.249
R1772 VTAIL.n445 VTAIL.n386 11.249
R1773 VTAIL.n416 VTAIL.n403 11.249
R1774 VTAIL.n368 VTAIL.n367 11.249
R1775 VTAIL.n351 VTAIL.n292 11.249
R1776 VTAIL.n322 VTAIL.n309 11.249
R1777 VTAIL.n698 VTAIL.n682 10.4732
R1778 VTAIL.n725 VTAIL.n670 10.4732
R1779 VTAIL.n747 VTAIL.n660 10.4732
R1780 VTAIL.n40 VTAIL.n24 10.4732
R1781 VTAIL.n67 VTAIL.n12 10.4732
R1782 VTAIL.n89 VTAIL.n2 10.4732
R1783 VTAIL.n134 VTAIL.n118 10.4732
R1784 VTAIL.n161 VTAIL.n106 10.4732
R1785 VTAIL.n183 VTAIL.n96 10.4732
R1786 VTAIL.n228 VTAIL.n212 10.4732
R1787 VTAIL.n255 VTAIL.n200 10.4732
R1788 VTAIL.n277 VTAIL.n190 10.4732
R1789 VTAIL.n653 VTAIL.n566 10.4732
R1790 VTAIL.n632 VTAIL.n577 10.4732
R1791 VTAIL.n605 VTAIL.n589 10.4732
R1792 VTAIL.n559 VTAIL.n472 10.4732
R1793 VTAIL.n538 VTAIL.n483 10.4732
R1794 VTAIL.n511 VTAIL.n495 10.4732
R1795 VTAIL.n465 VTAIL.n378 10.4732
R1796 VTAIL.n444 VTAIL.n389 10.4732
R1797 VTAIL.n417 VTAIL.n401 10.4732
R1798 VTAIL.n371 VTAIL.n284 10.4732
R1799 VTAIL.n350 VTAIL.n295 10.4732
R1800 VTAIL.n323 VTAIL.n307 10.4732
R1801 VTAIL.n702 VTAIL.n701 9.69747
R1802 VTAIL.n722 VTAIL.n721 9.69747
R1803 VTAIL.n748 VTAIL.n658 9.69747
R1804 VTAIL.n44 VTAIL.n43 9.69747
R1805 VTAIL.n64 VTAIL.n63 9.69747
R1806 VTAIL.n90 VTAIL.n0 9.69747
R1807 VTAIL.n138 VTAIL.n137 9.69747
R1808 VTAIL.n158 VTAIL.n157 9.69747
R1809 VTAIL.n184 VTAIL.n94 9.69747
R1810 VTAIL.n232 VTAIL.n231 9.69747
R1811 VTAIL.n252 VTAIL.n251 9.69747
R1812 VTAIL.n278 VTAIL.n188 9.69747
R1813 VTAIL.n654 VTAIL.n564 9.69747
R1814 VTAIL.n629 VTAIL.n628 9.69747
R1815 VTAIL.n609 VTAIL.n608 9.69747
R1816 VTAIL.n560 VTAIL.n470 9.69747
R1817 VTAIL.n535 VTAIL.n534 9.69747
R1818 VTAIL.n515 VTAIL.n514 9.69747
R1819 VTAIL.n466 VTAIL.n376 9.69747
R1820 VTAIL.n441 VTAIL.n440 9.69747
R1821 VTAIL.n421 VTAIL.n420 9.69747
R1822 VTAIL.n372 VTAIL.n282 9.69747
R1823 VTAIL.n347 VTAIL.n346 9.69747
R1824 VTAIL.n327 VTAIL.n326 9.69747
R1825 VTAIL.n750 VTAIL.n749 9.45567
R1826 VTAIL.n92 VTAIL.n91 9.45567
R1827 VTAIL.n186 VTAIL.n185 9.45567
R1828 VTAIL.n280 VTAIL.n279 9.45567
R1829 VTAIL.n656 VTAIL.n655 9.45567
R1830 VTAIL.n562 VTAIL.n561 9.45567
R1831 VTAIL.n468 VTAIL.n467 9.45567
R1832 VTAIL.n374 VTAIL.n373 9.45567
R1833 VTAIL.n749 VTAIL.n748 9.3005
R1834 VTAIL.n660 VTAIL.n659 9.3005
R1835 VTAIL.n743 VTAIL.n742 9.3005
R1836 VTAIL.n741 VTAIL.n740 9.3005
R1837 VTAIL.n664 VTAIL.n663 9.3005
R1838 VTAIL.n709 VTAIL.n708 9.3005
R1839 VTAIL.n707 VTAIL.n706 9.3005
R1840 VTAIL.n680 VTAIL.n679 9.3005
R1841 VTAIL.n701 VTAIL.n700 9.3005
R1842 VTAIL.n699 VTAIL.n698 9.3005
R1843 VTAIL.n684 VTAIL.n683 9.3005
R1844 VTAIL.n693 VTAIL.n692 9.3005
R1845 VTAIL.n691 VTAIL.n690 9.3005
R1846 VTAIL.n676 VTAIL.n675 9.3005
R1847 VTAIL.n715 VTAIL.n714 9.3005
R1848 VTAIL.n717 VTAIL.n716 9.3005
R1849 VTAIL.n672 VTAIL.n671 9.3005
R1850 VTAIL.n723 VTAIL.n722 9.3005
R1851 VTAIL.n725 VTAIL.n724 9.3005
R1852 VTAIL.n668 VTAIL.n667 9.3005
R1853 VTAIL.n732 VTAIL.n731 9.3005
R1854 VTAIL.n734 VTAIL.n733 9.3005
R1855 VTAIL.n91 VTAIL.n90 9.3005
R1856 VTAIL.n2 VTAIL.n1 9.3005
R1857 VTAIL.n85 VTAIL.n84 9.3005
R1858 VTAIL.n83 VTAIL.n82 9.3005
R1859 VTAIL.n6 VTAIL.n5 9.3005
R1860 VTAIL.n51 VTAIL.n50 9.3005
R1861 VTAIL.n49 VTAIL.n48 9.3005
R1862 VTAIL.n22 VTAIL.n21 9.3005
R1863 VTAIL.n43 VTAIL.n42 9.3005
R1864 VTAIL.n41 VTAIL.n40 9.3005
R1865 VTAIL.n26 VTAIL.n25 9.3005
R1866 VTAIL.n35 VTAIL.n34 9.3005
R1867 VTAIL.n33 VTAIL.n32 9.3005
R1868 VTAIL.n18 VTAIL.n17 9.3005
R1869 VTAIL.n57 VTAIL.n56 9.3005
R1870 VTAIL.n59 VTAIL.n58 9.3005
R1871 VTAIL.n14 VTAIL.n13 9.3005
R1872 VTAIL.n65 VTAIL.n64 9.3005
R1873 VTAIL.n67 VTAIL.n66 9.3005
R1874 VTAIL.n10 VTAIL.n9 9.3005
R1875 VTAIL.n74 VTAIL.n73 9.3005
R1876 VTAIL.n76 VTAIL.n75 9.3005
R1877 VTAIL.n185 VTAIL.n184 9.3005
R1878 VTAIL.n96 VTAIL.n95 9.3005
R1879 VTAIL.n179 VTAIL.n178 9.3005
R1880 VTAIL.n177 VTAIL.n176 9.3005
R1881 VTAIL.n100 VTAIL.n99 9.3005
R1882 VTAIL.n145 VTAIL.n144 9.3005
R1883 VTAIL.n143 VTAIL.n142 9.3005
R1884 VTAIL.n116 VTAIL.n115 9.3005
R1885 VTAIL.n137 VTAIL.n136 9.3005
R1886 VTAIL.n135 VTAIL.n134 9.3005
R1887 VTAIL.n120 VTAIL.n119 9.3005
R1888 VTAIL.n129 VTAIL.n128 9.3005
R1889 VTAIL.n127 VTAIL.n126 9.3005
R1890 VTAIL.n112 VTAIL.n111 9.3005
R1891 VTAIL.n151 VTAIL.n150 9.3005
R1892 VTAIL.n153 VTAIL.n152 9.3005
R1893 VTAIL.n108 VTAIL.n107 9.3005
R1894 VTAIL.n159 VTAIL.n158 9.3005
R1895 VTAIL.n161 VTAIL.n160 9.3005
R1896 VTAIL.n104 VTAIL.n103 9.3005
R1897 VTAIL.n168 VTAIL.n167 9.3005
R1898 VTAIL.n170 VTAIL.n169 9.3005
R1899 VTAIL.n279 VTAIL.n278 9.3005
R1900 VTAIL.n190 VTAIL.n189 9.3005
R1901 VTAIL.n273 VTAIL.n272 9.3005
R1902 VTAIL.n271 VTAIL.n270 9.3005
R1903 VTAIL.n194 VTAIL.n193 9.3005
R1904 VTAIL.n239 VTAIL.n238 9.3005
R1905 VTAIL.n237 VTAIL.n236 9.3005
R1906 VTAIL.n210 VTAIL.n209 9.3005
R1907 VTAIL.n231 VTAIL.n230 9.3005
R1908 VTAIL.n229 VTAIL.n228 9.3005
R1909 VTAIL.n214 VTAIL.n213 9.3005
R1910 VTAIL.n223 VTAIL.n222 9.3005
R1911 VTAIL.n221 VTAIL.n220 9.3005
R1912 VTAIL.n206 VTAIL.n205 9.3005
R1913 VTAIL.n245 VTAIL.n244 9.3005
R1914 VTAIL.n247 VTAIL.n246 9.3005
R1915 VTAIL.n202 VTAIL.n201 9.3005
R1916 VTAIL.n253 VTAIL.n252 9.3005
R1917 VTAIL.n255 VTAIL.n254 9.3005
R1918 VTAIL.n198 VTAIL.n197 9.3005
R1919 VTAIL.n262 VTAIL.n261 9.3005
R1920 VTAIL.n264 VTAIL.n263 9.3005
R1921 VTAIL.n622 VTAIL.n621 9.3005
R1922 VTAIL.n624 VTAIL.n623 9.3005
R1923 VTAIL.n579 VTAIL.n578 9.3005
R1924 VTAIL.n630 VTAIL.n629 9.3005
R1925 VTAIL.n632 VTAIL.n631 9.3005
R1926 VTAIL.n574 VTAIL.n573 9.3005
R1927 VTAIL.n638 VTAIL.n637 9.3005
R1928 VTAIL.n640 VTAIL.n639 9.3005
R1929 VTAIL.n655 VTAIL.n654 9.3005
R1930 VTAIL.n566 VTAIL.n565 9.3005
R1931 VTAIL.n649 VTAIL.n648 9.3005
R1932 VTAIL.n647 VTAIL.n646 9.3005
R1933 VTAIL.n570 VTAIL.n569 9.3005
R1934 VTAIL.n583 VTAIL.n582 9.3005
R1935 VTAIL.n616 VTAIL.n615 9.3005
R1936 VTAIL.n614 VTAIL.n613 9.3005
R1937 VTAIL.n587 VTAIL.n586 9.3005
R1938 VTAIL.n608 VTAIL.n607 9.3005
R1939 VTAIL.n606 VTAIL.n605 9.3005
R1940 VTAIL.n591 VTAIL.n590 9.3005
R1941 VTAIL.n600 VTAIL.n599 9.3005
R1942 VTAIL.n598 VTAIL.n597 9.3005
R1943 VTAIL.n528 VTAIL.n527 9.3005
R1944 VTAIL.n530 VTAIL.n529 9.3005
R1945 VTAIL.n485 VTAIL.n484 9.3005
R1946 VTAIL.n536 VTAIL.n535 9.3005
R1947 VTAIL.n538 VTAIL.n537 9.3005
R1948 VTAIL.n480 VTAIL.n479 9.3005
R1949 VTAIL.n544 VTAIL.n543 9.3005
R1950 VTAIL.n546 VTAIL.n545 9.3005
R1951 VTAIL.n561 VTAIL.n560 9.3005
R1952 VTAIL.n472 VTAIL.n471 9.3005
R1953 VTAIL.n555 VTAIL.n554 9.3005
R1954 VTAIL.n553 VTAIL.n552 9.3005
R1955 VTAIL.n476 VTAIL.n475 9.3005
R1956 VTAIL.n489 VTAIL.n488 9.3005
R1957 VTAIL.n522 VTAIL.n521 9.3005
R1958 VTAIL.n520 VTAIL.n519 9.3005
R1959 VTAIL.n493 VTAIL.n492 9.3005
R1960 VTAIL.n514 VTAIL.n513 9.3005
R1961 VTAIL.n512 VTAIL.n511 9.3005
R1962 VTAIL.n497 VTAIL.n496 9.3005
R1963 VTAIL.n506 VTAIL.n505 9.3005
R1964 VTAIL.n504 VTAIL.n503 9.3005
R1965 VTAIL.n434 VTAIL.n433 9.3005
R1966 VTAIL.n436 VTAIL.n435 9.3005
R1967 VTAIL.n391 VTAIL.n390 9.3005
R1968 VTAIL.n442 VTAIL.n441 9.3005
R1969 VTAIL.n444 VTAIL.n443 9.3005
R1970 VTAIL.n386 VTAIL.n385 9.3005
R1971 VTAIL.n450 VTAIL.n449 9.3005
R1972 VTAIL.n452 VTAIL.n451 9.3005
R1973 VTAIL.n467 VTAIL.n466 9.3005
R1974 VTAIL.n378 VTAIL.n377 9.3005
R1975 VTAIL.n461 VTAIL.n460 9.3005
R1976 VTAIL.n459 VTAIL.n458 9.3005
R1977 VTAIL.n382 VTAIL.n381 9.3005
R1978 VTAIL.n395 VTAIL.n394 9.3005
R1979 VTAIL.n428 VTAIL.n427 9.3005
R1980 VTAIL.n426 VTAIL.n425 9.3005
R1981 VTAIL.n399 VTAIL.n398 9.3005
R1982 VTAIL.n420 VTAIL.n419 9.3005
R1983 VTAIL.n418 VTAIL.n417 9.3005
R1984 VTAIL.n403 VTAIL.n402 9.3005
R1985 VTAIL.n412 VTAIL.n411 9.3005
R1986 VTAIL.n410 VTAIL.n409 9.3005
R1987 VTAIL.n340 VTAIL.n339 9.3005
R1988 VTAIL.n342 VTAIL.n341 9.3005
R1989 VTAIL.n297 VTAIL.n296 9.3005
R1990 VTAIL.n348 VTAIL.n347 9.3005
R1991 VTAIL.n350 VTAIL.n349 9.3005
R1992 VTAIL.n292 VTAIL.n291 9.3005
R1993 VTAIL.n356 VTAIL.n355 9.3005
R1994 VTAIL.n358 VTAIL.n357 9.3005
R1995 VTAIL.n373 VTAIL.n372 9.3005
R1996 VTAIL.n284 VTAIL.n283 9.3005
R1997 VTAIL.n367 VTAIL.n366 9.3005
R1998 VTAIL.n365 VTAIL.n364 9.3005
R1999 VTAIL.n288 VTAIL.n287 9.3005
R2000 VTAIL.n301 VTAIL.n300 9.3005
R2001 VTAIL.n334 VTAIL.n333 9.3005
R2002 VTAIL.n332 VTAIL.n331 9.3005
R2003 VTAIL.n305 VTAIL.n304 9.3005
R2004 VTAIL.n326 VTAIL.n325 9.3005
R2005 VTAIL.n324 VTAIL.n323 9.3005
R2006 VTAIL.n309 VTAIL.n308 9.3005
R2007 VTAIL.n318 VTAIL.n317 9.3005
R2008 VTAIL.n316 VTAIL.n315 9.3005
R2009 VTAIL.n705 VTAIL.n680 8.92171
R2010 VTAIL.n718 VTAIL.n672 8.92171
R2011 VTAIL.n47 VTAIL.n22 8.92171
R2012 VTAIL.n60 VTAIL.n14 8.92171
R2013 VTAIL.n141 VTAIL.n116 8.92171
R2014 VTAIL.n154 VTAIL.n108 8.92171
R2015 VTAIL.n235 VTAIL.n210 8.92171
R2016 VTAIL.n248 VTAIL.n202 8.92171
R2017 VTAIL.n625 VTAIL.n579 8.92171
R2018 VTAIL.n612 VTAIL.n587 8.92171
R2019 VTAIL.n531 VTAIL.n485 8.92171
R2020 VTAIL.n518 VTAIL.n493 8.92171
R2021 VTAIL.n437 VTAIL.n391 8.92171
R2022 VTAIL.n424 VTAIL.n399 8.92171
R2023 VTAIL.n343 VTAIL.n297 8.92171
R2024 VTAIL.n330 VTAIL.n305 8.92171
R2025 VTAIL.n706 VTAIL.n678 8.14595
R2026 VTAIL.n717 VTAIL.n674 8.14595
R2027 VTAIL.n48 VTAIL.n20 8.14595
R2028 VTAIL.n59 VTAIL.n16 8.14595
R2029 VTAIL.n142 VTAIL.n114 8.14595
R2030 VTAIL.n153 VTAIL.n110 8.14595
R2031 VTAIL.n236 VTAIL.n208 8.14595
R2032 VTAIL.n247 VTAIL.n204 8.14595
R2033 VTAIL.n624 VTAIL.n581 8.14595
R2034 VTAIL.n613 VTAIL.n585 8.14595
R2035 VTAIL.n530 VTAIL.n487 8.14595
R2036 VTAIL.n519 VTAIL.n491 8.14595
R2037 VTAIL.n436 VTAIL.n393 8.14595
R2038 VTAIL.n425 VTAIL.n397 8.14595
R2039 VTAIL.n342 VTAIL.n299 8.14595
R2040 VTAIL.n331 VTAIL.n303 8.14595
R2041 VTAIL.n710 VTAIL.n709 7.3702
R2042 VTAIL.n714 VTAIL.n713 7.3702
R2043 VTAIL.n52 VTAIL.n51 7.3702
R2044 VTAIL.n56 VTAIL.n55 7.3702
R2045 VTAIL.n146 VTAIL.n145 7.3702
R2046 VTAIL.n150 VTAIL.n149 7.3702
R2047 VTAIL.n240 VTAIL.n239 7.3702
R2048 VTAIL.n244 VTAIL.n243 7.3702
R2049 VTAIL.n621 VTAIL.n620 7.3702
R2050 VTAIL.n617 VTAIL.n616 7.3702
R2051 VTAIL.n527 VTAIL.n526 7.3702
R2052 VTAIL.n523 VTAIL.n522 7.3702
R2053 VTAIL.n433 VTAIL.n432 7.3702
R2054 VTAIL.n429 VTAIL.n428 7.3702
R2055 VTAIL.n339 VTAIL.n338 7.3702
R2056 VTAIL.n335 VTAIL.n334 7.3702
R2057 VTAIL.n710 VTAIL.n676 6.59444
R2058 VTAIL.n713 VTAIL.n676 6.59444
R2059 VTAIL.n52 VTAIL.n18 6.59444
R2060 VTAIL.n55 VTAIL.n18 6.59444
R2061 VTAIL.n146 VTAIL.n112 6.59444
R2062 VTAIL.n149 VTAIL.n112 6.59444
R2063 VTAIL.n240 VTAIL.n206 6.59444
R2064 VTAIL.n243 VTAIL.n206 6.59444
R2065 VTAIL.n620 VTAIL.n583 6.59444
R2066 VTAIL.n617 VTAIL.n583 6.59444
R2067 VTAIL.n526 VTAIL.n489 6.59444
R2068 VTAIL.n523 VTAIL.n489 6.59444
R2069 VTAIL.n432 VTAIL.n395 6.59444
R2070 VTAIL.n429 VTAIL.n395 6.59444
R2071 VTAIL.n338 VTAIL.n301 6.59444
R2072 VTAIL.n335 VTAIL.n301 6.59444
R2073 VTAIL.n709 VTAIL.n678 5.81868
R2074 VTAIL.n714 VTAIL.n674 5.81868
R2075 VTAIL.n51 VTAIL.n20 5.81868
R2076 VTAIL.n56 VTAIL.n16 5.81868
R2077 VTAIL.n145 VTAIL.n114 5.81868
R2078 VTAIL.n150 VTAIL.n110 5.81868
R2079 VTAIL.n239 VTAIL.n208 5.81868
R2080 VTAIL.n244 VTAIL.n204 5.81868
R2081 VTAIL.n621 VTAIL.n581 5.81868
R2082 VTAIL.n616 VTAIL.n585 5.81868
R2083 VTAIL.n527 VTAIL.n487 5.81868
R2084 VTAIL.n522 VTAIL.n491 5.81868
R2085 VTAIL.n433 VTAIL.n393 5.81868
R2086 VTAIL.n428 VTAIL.n397 5.81868
R2087 VTAIL.n339 VTAIL.n299 5.81868
R2088 VTAIL.n334 VTAIL.n303 5.81868
R2089 VTAIL.n706 VTAIL.n705 5.04292
R2090 VTAIL.n718 VTAIL.n717 5.04292
R2091 VTAIL.n48 VTAIL.n47 5.04292
R2092 VTAIL.n60 VTAIL.n59 5.04292
R2093 VTAIL.n142 VTAIL.n141 5.04292
R2094 VTAIL.n154 VTAIL.n153 5.04292
R2095 VTAIL.n236 VTAIL.n235 5.04292
R2096 VTAIL.n248 VTAIL.n247 5.04292
R2097 VTAIL.n625 VTAIL.n624 5.04292
R2098 VTAIL.n613 VTAIL.n612 5.04292
R2099 VTAIL.n531 VTAIL.n530 5.04292
R2100 VTAIL.n519 VTAIL.n518 5.04292
R2101 VTAIL.n437 VTAIL.n436 5.04292
R2102 VTAIL.n425 VTAIL.n424 5.04292
R2103 VTAIL.n343 VTAIL.n342 5.04292
R2104 VTAIL.n331 VTAIL.n330 5.04292
R2105 VTAIL.n702 VTAIL.n680 4.26717
R2106 VTAIL.n721 VTAIL.n672 4.26717
R2107 VTAIL.n750 VTAIL.n658 4.26717
R2108 VTAIL.n44 VTAIL.n22 4.26717
R2109 VTAIL.n63 VTAIL.n14 4.26717
R2110 VTAIL.n92 VTAIL.n0 4.26717
R2111 VTAIL.n138 VTAIL.n116 4.26717
R2112 VTAIL.n157 VTAIL.n108 4.26717
R2113 VTAIL.n186 VTAIL.n94 4.26717
R2114 VTAIL.n232 VTAIL.n210 4.26717
R2115 VTAIL.n251 VTAIL.n202 4.26717
R2116 VTAIL.n280 VTAIL.n188 4.26717
R2117 VTAIL.n656 VTAIL.n564 4.26717
R2118 VTAIL.n628 VTAIL.n579 4.26717
R2119 VTAIL.n609 VTAIL.n587 4.26717
R2120 VTAIL.n562 VTAIL.n470 4.26717
R2121 VTAIL.n534 VTAIL.n485 4.26717
R2122 VTAIL.n515 VTAIL.n493 4.26717
R2123 VTAIL.n468 VTAIL.n376 4.26717
R2124 VTAIL.n440 VTAIL.n391 4.26717
R2125 VTAIL.n421 VTAIL.n399 4.26717
R2126 VTAIL.n374 VTAIL.n282 4.26717
R2127 VTAIL.n346 VTAIL.n297 4.26717
R2128 VTAIL.n327 VTAIL.n305 4.26717
R2129 VTAIL.n691 VTAIL.n687 3.70982
R2130 VTAIL.n33 VTAIL.n29 3.70982
R2131 VTAIL.n127 VTAIL.n123 3.70982
R2132 VTAIL.n221 VTAIL.n217 3.70982
R2133 VTAIL.n598 VTAIL.n594 3.70982
R2134 VTAIL.n504 VTAIL.n500 3.70982
R2135 VTAIL.n410 VTAIL.n406 3.70982
R2136 VTAIL.n316 VTAIL.n312 3.70982
R2137 VTAIL.n701 VTAIL.n682 3.49141
R2138 VTAIL.n722 VTAIL.n670 3.49141
R2139 VTAIL.n748 VTAIL.n747 3.49141
R2140 VTAIL.n43 VTAIL.n24 3.49141
R2141 VTAIL.n64 VTAIL.n12 3.49141
R2142 VTAIL.n90 VTAIL.n89 3.49141
R2143 VTAIL.n137 VTAIL.n118 3.49141
R2144 VTAIL.n158 VTAIL.n106 3.49141
R2145 VTAIL.n184 VTAIL.n183 3.49141
R2146 VTAIL.n231 VTAIL.n212 3.49141
R2147 VTAIL.n252 VTAIL.n200 3.49141
R2148 VTAIL.n278 VTAIL.n277 3.49141
R2149 VTAIL.n654 VTAIL.n653 3.49141
R2150 VTAIL.n629 VTAIL.n577 3.49141
R2151 VTAIL.n608 VTAIL.n589 3.49141
R2152 VTAIL.n560 VTAIL.n559 3.49141
R2153 VTAIL.n535 VTAIL.n483 3.49141
R2154 VTAIL.n514 VTAIL.n495 3.49141
R2155 VTAIL.n466 VTAIL.n465 3.49141
R2156 VTAIL.n441 VTAIL.n389 3.49141
R2157 VTAIL.n420 VTAIL.n401 3.49141
R2158 VTAIL.n372 VTAIL.n371 3.49141
R2159 VTAIL.n347 VTAIL.n295 3.49141
R2160 VTAIL.n326 VTAIL.n307 3.49141
R2161 VTAIL.n469 VTAIL.n375 3.31084
R2162 VTAIL.n657 VTAIL.n563 3.31084
R2163 VTAIL.n281 VTAIL.n187 3.31084
R2164 VTAIL.n698 VTAIL.n697 2.71565
R2165 VTAIL.n726 VTAIL.n725 2.71565
R2166 VTAIL.n744 VTAIL.n660 2.71565
R2167 VTAIL.n40 VTAIL.n39 2.71565
R2168 VTAIL.n68 VTAIL.n67 2.71565
R2169 VTAIL.n86 VTAIL.n2 2.71565
R2170 VTAIL.n134 VTAIL.n133 2.71565
R2171 VTAIL.n162 VTAIL.n161 2.71565
R2172 VTAIL.n180 VTAIL.n96 2.71565
R2173 VTAIL.n228 VTAIL.n227 2.71565
R2174 VTAIL.n256 VTAIL.n255 2.71565
R2175 VTAIL.n274 VTAIL.n190 2.71565
R2176 VTAIL.n650 VTAIL.n566 2.71565
R2177 VTAIL.n633 VTAIL.n632 2.71565
R2178 VTAIL.n605 VTAIL.n604 2.71565
R2179 VTAIL.n556 VTAIL.n472 2.71565
R2180 VTAIL.n539 VTAIL.n538 2.71565
R2181 VTAIL.n511 VTAIL.n510 2.71565
R2182 VTAIL.n462 VTAIL.n378 2.71565
R2183 VTAIL.n445 VTAIL.n444 2.71565
R2184 VTAIL.n417 VTAIL.n416 2.71565
R2185 VTAIL.n368 VTAIL.n284 2.71565
R2186 VTAIL.n351 VTAIL.n350 2.71565
R2187 VTAIL.n323 VTAIL.n322 2.71565
R2188 VTAIL.n694 VTAIL.n684 1.93989
R2189 VTAIL.n730 VTAIL.n668 1.93989
R2190 VTAIL.n743 VTAIL.n662 1.93989
R2191 VTAIL.n36 VTAIL.n26 1.93989
R2192 VTAIL.n72 VTAIL.n10 1.93989
R2193 VTAIL.n85 VTAIL.n4 1.93989
R2194 VTAIL.n130 VTAIL.n120 1.93989
R2195 VTAIL.n166 VTAIL.n104 1.93989
R2196 VTAIL.n179 VTAIL.n98 1.93989
R2197 VTAIL.n224 VTAIL.n214 1.93989
R2198 VTAIL.n260 VTAIL.n198 1.93989
R2199 VTAIL.n273 VTAIL.n192 1.93989
R2200 VTAIL.n649 VTAIL.n568 1.93989
R2201 VTAIL.n636 VTAIL.n574 1.93989
R2202 VTAIL.n601 VTAIL.n591 1.93989
R2203 VTAIL.n555 VTAIL.n474 1.93989
R2204 VTAIL.n542 VTAIL.n480 1.93989
R2205 VTAIL.n507 VTAIL.n497 1.93989
R2206 VTAIL.n461 VTAIL.n380 1.93989
R2207 VTAIL.n448 VTAIL.n386 1.93989
R2208 VTAIL.n413 VTAIL.n403 1.93989
R2209 VTAIL.n367 VTAIL.n286 1.93989
R2210 VTAIL.n354 VTAIL.n292 1.93989
R2211 VTAIL.n319 VTAIL.n309 1.93989
R2212 VTAIL VTAIL.n93 1.71386
R2213 VTAIL VTAIL.n751 1.59748
R2214 VTAIL.n693 VTAIL.n686 1.16414
R2215 VTAIL.n731 VTAIL.n666 1.16414
R2216 VTAIL.n740 VTAIL.n739 1.16414
R2217 VTAIL.n35 VTAIL.n28 1.16414
R2218 VTAIL.n73 VTAIL.n8 1.16414
R2219 VTAIL.n82 VTAIL.n81 1.16414
R2220 VTAIL.n129 VTAIL.n122 1.16414
R2221 VTAIL.n167 VTAIL.n102 1.16414
R2222 VTAIL.n176 VTAIL.n175 1.16414
R2223 VTAIL.n223 VTAIL.n216 1.16414
R2224 VTAIL.n261 VTAIL.n196 1.16414
R2225 VTAIL.n270 VTAIL.n269 1.16414
R2226 VTAIL.n646 VTAIL.n645 1.16414
R2227 VTAIL.n637 VTAIL.n572 1.16414
R2228 VTAIL.n600 VTAIL.n593 1.16414
R2229 VTAIL.n552 VTAIL.n551 1.16414
R2230 VTAIL.n543 VTAIL.n478 1.16414
R2231 VTAIL.n506 VTAIL.n499 1.16414
R2232 VTAIL.n458 VTAIL.n457 1.16414
R2233 VTAIL.n449 VTAIL.n384 1.16414
R2234 VTAIL.n412 VTAIL.n405 1.16414
R2235 VTAIL.n364 VTAIL.n363 1.16414
R2236 VTAIL.n355 VTAIL.n290 1.16414
R2237 VTAIL.n318 VTAIL.n311 1.16414
R2238 VTAIL.n563 VTAIL.n469 0.470328
R2239 VTAIL.n187 VTAIL.n93 0.470328
R2240 VTAIL.n690 VTAIL.n689 0.388379
R2241 VTAIL.n735 VTAIL.n734 0.388379
R2242 VTAIL.n736 VTAIL.n664 0.388379
R2243 VTAIL.n32 VTAIL.n31 0.388379
R2244 VTAIL.n77 VTAIL.n76 0.388379
R2245 VTAIL.n78 VTAIL.n6 0.388379
R2246 VTAIL.n126 VTAIL.n125 0.388379
R2247 VTAIL.n171 VTAIL.n170 0.388379
R2248 VTAIL.n172 VTAIL.n100 0.388379
R2249 VTAIL.n220 VTAIL.n219 0.388379
R2250 VTAIL.n265 VTAIL.n264 0.388379
R2251 VTAIL.n266 VTAIL.n194 0.388379
R2252 VTAIL.n642 VTAIL.n570 0.388379
R2253 VTAIL.n641 VTAIL.n640 0.388379
R2254 VTAIL.n597 VTAIL.n596 0.388379
R2255 VTAIL.n548 VTAIL.n476 0.388379
R2256 VTAIL.n547 VTAIL.n546 0.388379
R2257 VTAIL.n503 VTAIL.n502 0.388379
R2258 VTAIL.n454 VTAIL.n382 0.388379
R2259 VTAIL.n453 VTAIL.n452 0.388379
R2260 VTAIL.n409 VTAIL.n408 0.388379
R2261 VTAIL.n360 VTAIL.n288 0.388379
R2262 VTAIL.n359 VTAIL.n358 0.388379
R2263 VTAIL.n315 VTAIL.n314 0.388379
R2264 VTAIL.n692 VTAIL.n691 0.155672
R2265 VTAIL.n692 VTAIL.n683 0.155672
R2266 VTAIL.n699 VTAIL.n683 0.155672
R2267 VTAIL.n700 VTAIL.n699 0.155672
R2268 VTAIL.n700 VTAIL.n679 0.155672
R2269 VTAIL.n707 VTAIL.n679 0.155672
R2270 VTAIL.n708 VTAIL.n707 0.155672
R2271 VTAIL.n708 VTAIL.n675 0.155672
R2272 VTAIL.n715 VTAIL.n675 0.155672
R2273 VTAIL.n716 VTAIL.n715 0.155672
R2274 VTAIL.n716 VTAIL.n671 0.155672
R2275 VTAIL.n723 VTAIL.n671 0.155672
R2276 VTAIL.n724 VTAIL.n723 0.155672
R2277 VTAIL.n724 VTAIL.n667 0.155672
R2278 VTAIL.n732 VTAIL.n667 0.155672
R2279 VTAIL.n733 VTAIL.n732 0.155672
R2280 VTAIL.n733 VTAIL.n663 0.155672
R2281 VTAIL.n741 VTAIL.n663 0.155672
R2282 VTAIL.n742 VTAIL.n741 0.155672
R2283 VTAIL.n742 VTAIL.n659 0.155672
R2284 VTAIL.n749 VTAIL.n659 0.155672
R2285 VTAIL.n34 VTAIL.n33 0.155672
R2286 VTAIL.n34 VTAIL.n25 0.155672
R2287 VTAIL.n41 VTAIL.n25 0.155672
R2288 VTAIL.n42 VTAIL.n41 0.155672
R2289 VTAIL.n42 VTAIL.n21 0.155672
R2290 VTAIL.n49 VTAIL.n21 0.155672
R2291 VTAIL.n50 VTAIL.n49 0.155672
R2292 VTAIL.n50 VTAIL.n17 0.155672
R2293 VTAIL.n57 VTAIL.n17 0.155672
R2294 VTAIL.n58 VTAIL.n57 0.155672
R2295 VTAIL.n58 VTAIL.n13 0.155672
R2296 VTAIL.n65 VTAIL.n13 0.155672
R2297 VTAIL.n66 VTAIL.n65 0.155672
R2298 VTAIL.n66 VTAIL.n9 0.155672
R2299 VTAIL.n74 VTAIL.n9 0.155672
R2300 VTAIL.n75 VTAIL.n74 0.155672
R2301 VTAIL.n75 VTAIL.n5 0.155672
R2302 VTAIL.n83 VTAIL.n5 0.155672
R2303 VTAIL.n84 VTAIL.n83 0.155672
R2304 VTAIL.n84 VTAIL.n1 0.155672
R2305 VTAIL.n91 VTAIL.n1 0.155672
R2306 VTAIL.n128 VTAIL.n127 0.155672
R2307 VTAIL.n128 VTAIL.n119 0.155672
R2308 VTAIL.n135 VTAIL.n119 0.155672
R2309 VTAIL.n136 VTAIL.n135 0.155672
R2310 VTAIL.n136 VTAIL.n115 0.155672
R2311 VTAIL.n143 VTAIL.n115 0.155672
R2312 VTAIL.n144 VTAIL.n143 0.155672
R2313 VTAIL.n144 VTAIL.n111 0.155672
R2314 VTAIL.n151 VTAIL.n111 0.155672
R2315 VTAIL.n152 VTAIL.n151 0.155672
R2316 VTAIL.n152 VTAIL.n107 0.155672
R2317 VTAIL.n159 VTAIL.n107 0.155672
R2318 VTAIL.n160 VTAIL.n159 0.155672
R2319 VTAIL.n160 VTAIL.n103 0.155672
R2320 VTAIL.n168 VTAIL.n103 0.155672
R2321 VTAIL.n169 VTAIL.n168 0.155672
R2322 VTAIL.n169 VTAIL.n99 0.155672
R2323 VTAIL.n177 VTAIL.n99 0.155672
R2324 VTAIL.n178 VTAIL.n177 0.155672
R2325 VTAIL.n178 VTAIL.n95 0.155672
R2326 VTAIL.n185 VTAIL.n95 0.155672
R2327 VTAIL.n222 VTAIL.n221 0.155672
R2328 VTAIL.n222 VTAIL.n213 0.155672
R2329 VTAIL.n229 VTAIL.n213 0.155672
R2330 VTAIL.n230 VTAIL.n229 0.155672
R2331 VTAIL.n230 VTAIL.n209 0.155672
R2332 VTAIL.n237 VTAIL.n209 0.155672
R2333 VTAIL.n238 VTAIL.n237 0.155672
R2334 VTAIL.n238 VTAIL.n205 0.155672
R2335 VTAIL.n245 VTAIL.n205 0.155672
R2336 VTAIL.n246 VTAIL.n245 0.155672
R2337 VTAIL.n246 VTAIL.n201 0.155672
R2338 VTAIL.n253 VTAIL.n201 0.155672
R2339 VTAIL.n254 VTAIL.n253 0.155672
R2340 VTAIL.n254 VTAIL.n197 0.155672
R2341 VTAIL.n262 VTAIL.n197 0.155672
R2342 VTAIL.n263 VTAIL.n262 0.155672
R2343 VTAIL.n263 VTAIL.n193 0.155672
R2344 VTAIL.n271 VTAIL.n193 0.155672
R2345 VTAIL.n272 VTAIL.n271 0.155672
R2346 VTAIL.n272 VTAIL.n189 0.155672
R2347 VTAIL.n279 VTAIL.n189 0.155672
R2348 VTAIL.n655 VTAIL.n565 0.155672
R2349 VTAIL.n648 VTAIL.n565 0.155672
R2350 VTAIL.n648 VTAIL.n647 0.155672
R2351 VTAIL.n647 VTAIL.n569 0.155672
R2352 VTAIL.n639 VTAIL.n569 0.155672
R2353 VTAIL.n639 VTAIL.n638 0.155672
R2354 VTAIL.n638 VTAIL.n573 0.155672
R2355 VTAIL.n631 VTAIL.n573 0.155672
R2356 VTAIL.n631 VTAIL.n630 0.155672
R2357 VTAIL.n630 VTAIL.n578 0.155672
R2358 VTAIL.n623 VTAIL.n578 0.155672
R2359 VTAIL.n623 VTAIL.n622 0.155672
R2360 VTAIL.n622 VTAIL.n582 0.155672
R2361 VTAIL.n615 VTAIL.n582 0.155672
R2362 VTAIL.n615 VTAIL.n614 0.155672
R2363 VTAIL.n614 VTAIL.n586 0.155672
R2364 VTAIL.n607 VTAIL.n586 0.155672
R2365 VTAIL.n607 VTAIL.n606 0.155672
R2366 VTAIL.n606 VTAIL.n590 0.155672
R2367 VTAIL.n599 VTAIL.n590 0.155672
R2368 VTAIL.n599 VTAIL.n598 0.155672
R2369 VTAIL.n561 VTAIL.n471 0.155672
R2370 VTAIL.n554 VTAIL.n471 0.155672
R2371 VTAIL.n554 VTAIL.n553 0.155672
R2372 VTAIL.n553 VTAIL.n475 0.155672
R2373 VTAIL.n545 VTAIL.n475 0.155672
R2374 VTAIL.n545 VTAIL.n544 0.155672
R2375 VTAIL.n544 VTAIL.n479 0.155672
R2376 VTAIL.n537 VTAIL.n479 0.155672
R2377 VTAIL.n537 VTAIL.n536 0.155672
R2378 VTAIL.n536 VTAIL.n484 0.155672
R2379 VTAIL.n529 VTAIL.n484 0.155672
R2380 VTAIL.n529 VTAIL.n528 0.155672
R2381 VTAIL.n528 VTAIL.n488 0.155672
R2382 VTAIL.n521 VTAIL.n488 0.155672
R2383 VTAIL.n521 VTAIL.n520 0.155672
R2384 VTAIL.n520 VTAIL.n492 0.155672
R2385 VTAIL.n513 VTAIL.n492 0.155672
R2386 VTAIL.n513 VTAIL.n512 0.155672
R2387 VTAIL.n512 VTAIL.n496 0.155672
R2388 VTAIL.n505 VTAIL.n496 0.155672
R2389 VTAIL.n505 VTAIL.n504 0.155672
R2390 VTAIL.n467 VTAIL.n377 0.155672
R2391 VTAIL.n460 VTAIL.n377 0.155672
R2392 VTAIL.n460 VTAIL.n459 0.155672
R2393 VTAIL.n459 VTAIL.n381 0.155672
R2394 VTAIL.n451 VTAIL.n381 0.155672
R2395 VTAIL.n451 VTAIL.n450 0.155672
R2396 VTAIL.n450 VTAIL.n385 0.155672
R2397 VTAIL.n443 VTAIL.n385 0.155672
R2398 VTAIL.n443 VTAIL.n442 0.155672
R2399 VTAIL.n442 VTAIL.n390 0.155672
R2400 VTAIL.n435 VTAIL.n390 0.155672
R2401 VTAIL.n435 VTAIL.n434 0.155672
R2402 VTAIL.n434 VTAIL.n394 0.155672
R2403 VTAIL.n427 VTAIL.n394 0.155672
R2404 VTAIL.n427 VTAIL.n426 0.155672
R2405 VTAIL.n426 VTAIL.n398 0.155672
R2406 VTAIL.n419 VTAIL.n398 0.155672
R2407 VTAIL.n419 VTAIL.n418 0.155672
R2408 VTAIL.n418 VTAIL.n402 0.155672
R2409 VTAIL.n411 VTAIL.n402 0.155672
R2410 VTAIL.n411 VTAIL.n410 0.155672
R2411 VTAIL.n373 VTAIL.n283 0.155672
R2412 VTAIL.n366 VTAIL.n283 0.155672
R2413 VTAIL.n366 VTAIL.n365 0.155672
R2414 VTAIL.n365 VTAIL.n287 0.155672
R2415 VTAIL.n357 VTAIL.n287 0.155672
R2416 VTAIL.n357 VTAIL.n356 0.155672
R2417 VTAIL.n356 VTAIL.n291 0.155672
R2418 VTAIL.n349 VTAIL.n291 0.155672
R2419 VTAIL.n349 VTAIL.n348 0.155672
R2420 VTAIL.n348 VTAIL.n296 0.155672
R2421 VTAIL.n341 VTAIL.n296 0.155672
R2422 VTAIL.n341 VTAIL.n340 0.155672
R2423 VTAIL.n340 VTAIL.n300 0.155672
R2424 VTAIL.n333 VTAIL.n300 0.155672
R2425 VTAIL.n333 VTAIL.n332 0.155672
R2426 VTAIL.n332 VTAIL.n304 0.155672
R2427 VTAIL.n325 VTAIL.n304 0.155672
R2428 VTAIL.n325 VTAIL.n324 0.155672
R2429 VTAIL.n324 VTAIL.n308 0.155672
R2430 VTAIL.n317 VTAIL.n308 0.155672
R2431 VTAIL.n317 VTAIL.n316 0.155672
R2432 VDD1 VDD1.n1 117.843
R2433 VDD1 VDD1.n0 69.2561
R2434 VDD1.n0 VDD1.t1 1.93647
R2435 VDD1.n0 VDD1.t2 1.93647
R2436 VDD1.n1 VDD1.t0 1.93647
R2437 VDD1.n1 VDD1.t3 1.93647
R2438 VN.n1 VN.t1 149.768
R2439 VN.n0 VN.t0 149.768
R2440 VN.n0 VN.t3 148.547
R2441 VN.n1 VN.t2 148.547
R2442 VN VN.n1 55.1186
R2443 VN VN.n0 2.19057
R2444 VDD2.n2 VDD2.n0 117.317
R2445 VDD2.n2 VDD2.n1 69.1979
R2446 VDD2.n1 VDD2.t1 1.93647
R2447 VDD2.n1 VDD2.t2 1.93647
R2448 VDD2.n0 VDD2.t3 1.93647
R2449 VDD2.n0 VDD2.t0 1.93647
R2450 VDD2 VDD2.n2 0.0586897
C0 VDD2 VN 6.835f
C1 VP VN 7.73552f
C2 VN VTAIL 6.65846f
C3 VDD1 VDD2 1.24418f
C4 VDD1 VP 7.13642f
C5 VDD1 VTAIL 6.66696f
C6 VDD2 VP 0.452361f
C7 VDD2 VTAIL 6.72726f
C8 VP VTAIL 6.67257f
C9 B VN 1.33765f
C10 w_n3274_n4326# VN 5.80409f
C11 VDD1 B 1.55186f
C12 VDD1 w_n3274_n4326# 1.75483f
C13 VDD2 B 1.61908f
C14 B VP 2.04415f
C15 VDD2 w_n3274_n4326# 1.83102f
C16 B VTAIL 6.96299f
C17 w_n3274_n4326# VP 6.22728f
C18 w_n3274_n4326# VTAIL 5.05564f
C19 w_n3274_n4326# B 11.7075f
C20 VDD1 VN 0.149973f
C21 VDD2 VSUBS 1.209129f
C22 VDD1 VSUBS 6.842639f
C23 VTAIL VSUBS 1.544344f
C24 VN VSUBS 6.0981f
C25 VP VSUBS 2.941612f
C26 B VSUBS 5.46428f
C27 w_n3274_n4326# VSUBS 0.173378p
C28 VDD2.t3 VSUBS 0.353343f
C29 VDD2.t0 VSUBS 0.353343f
C30 VDD2.n0 VSUBS 3.8711f
C31 VDD2.t1 VSUBS 0.353343f
C32 VDD2.t2 VSUBS 0.353343f
C33 VDD2.n1 VSUBS 2.90844f
C34 VDD2.n2 VSUBS 5.01729f
C35 VN.t3 VSUBS 4.456759f
C36 VN.t0 VSUBS 4.46942f
C37 VN.n0 VSUBS 2.72933f
C38 VN.t1 VSUBS 4.46942f
C39 VN.t2 VSUBS 4.456759f
C40 VN.n1 VSUBS 4.49228f
C41 VDD1.t1 VSUBS 0.358582f
C42 VDD1.t2 VSUBS 0.358582f
C43 VDD1.n0 VSUBS 2.95227f
C44 VDD1.t0 VSUBS 0.358582f
C45 VDD1.t3 VSUBS 0.358582f
C46 VDD1.n1 VSUBS 3.95658f
C47 VTAIL.n0 VSUBS 0.024405f
C48 VTAIL.n1 VSUBS 0.023101f
C49 VTAIL.n2 VSUBS 0.012414f
C50 VTAIL.n3 VSUBS 0.029341f
C51 VTAIL.n4 VSUBS 0.013144f
C52 VTAIL.n5 VSUBS 0.023101f
C53 VTAIL.n6 VSUBS 0.012414f
C54 VTAIL.n7 VSUBS 0.029341f
C55 VTAIL.n8 VSUBS 0.013144f
C56 VTAIL.n9 VSUBS 0.023101f
C57 VTAIL.n10 VSUBS 0.012414f
C58 VTAIL.n11 VSUBS 0.029341f
C59 VTAIL.n12 VSUBS 0.013144f
C60 VTAIL.n13 VSUBS 0.023101f
C61 VTAIL.n14 VSUBS 0.012414f
C62 VTAIL.n15 VSUBS 0.029341f
C63 VTAIL.n16 VSUBS 0.013144f
C64 VTAIL.n17 VSUBS 0.023101f
C65 VTAIL.n18 VSUBS 0.012414f
C66 VTAIL.n19 VSUBS 0.029341f
C67 VTAIL.n20 VSUBS 0.013144f
C68 VTAIL.n21 VSUBS 0.023101f
C69 VTAIL.n22 VSUBS 0.012414f
C70 VTAIL.n23 VSUBS 0.029341f
C71 VTAIL.n24 VSUBS 0.013144f
C72 VTAIL.n25 VSUBS 0.023101f
C73 VTAIL.n26 VSUBS 0.012414f
C74 VTAIL.n27 VSUBS 0.029341f
C75 VTAIL.n28 VSUBS 0.013144f
C76 VTAIL.n29 VSUBS 0.175041f
C77 VTAIL.t2 VSUBS 0.062917f
C78 VTAIL.n30 VSUBS 0.022006f
C79 VTAIL.n31 VSUBS 0.018666f
C80 VTAIL.n32 VSUBS 0.012414f
C81 VTAIL.n33 VSUBS 1.66279f
C82 VTAIL.n34 VSUBS 0.023101f
C83 VTAIL.n35 VSUBS 0.012414f
C84 VTAIL.n36 VSUBS 0.013144f
C85 VTAIL.n37 VSUBS 0.029341f
C86 VTAIL.n38 VSUBS 0.029341f
C87 VTAIL.n39 VSUBS 0.013144f
C88 VTAIL.n40 VSUBS 0.012414f
C89 VTAIL.n41 VSUBS 0.023101f
C90 VTAIL.n42 VSUBS 0.023101f
C91 VTAIL.n43 VSUBS 0.012414f
C92 VTAIL.n44 VSUBS 0.013144f
C93 VTAIL.n45 VSUBS 0.029341f
C94 VTAIL.n46 VSUBS 0.029341f
C95 VTAIL.n47 VSUBS 0.013144f
C96 VTAIL.n48 VSUBS 0.012414f
C97 VTAIL.n49 VSUBS 0.023101f
C98 VTAIL.n50 VSUBS 0.023101f
C99 VTAIL.n51 VSUBS 0.012414f
C100 VTAIL.n52 VSUBS 0.013144f
C101 VTAIL.n53 VSUBS 0.029341f
C102 VTAIL.n54 VSUBS 0.029341f
C103 VTAIL.n55 VSUBS 0.013144f
C104 VTAIL.n56 VSUBS 0.012414f
C105 VTAIL.n57 VSUBS 0.023101f
C106 VTAIL.n58 VSUBS 0.023101f
C107 VTAIL.n59 VSUBS 0.012414f
C108 VTAIL.n60 VSUBS 0.013144f
C109 VTAIL.n61 VSUBS 0.029341f
C110 VTAIL.n62 VSUBS 0.029341f
C111 VTAIL.n63 VSUBS 0.013144f
C112 VTAIL.n64 VSUBS 0.012414f
C113 VTAIL.n65 VSUBS 0.023101f
C114 VTAIL.n66 VSUBS 0.023101f
C115 VTAIL.n67 VSUBS 0.012414f
C116 VTAIL.n68 VSUBS 0.013144f
C117 VTAIL.n69 VSUBS 0.029341f
C118 VTAIL.n70 VSUBS 0.029341f
C119 VTAIL.n71 VSUBS 0.029341f
C120 VTAIL.n72 VSUBS 0.013144f
C121 VTAIL.n73 VSUBS 0.012414f
C122 VTAIL.n74 VSUBS 0.023101f
C123 VTAIL.n75 VSUBS 0.023101f
C124 VTAIL.n76 VSUBS 0.012414f
C125 VTAIL.n77 VSUBS 0.012779f
C126 VTAIL.n78 VSUBS 0.012779f
C127 VTAIL.n79 VSUBS 0.029341f
C128 VTAIL.n80 VSUBS 0.029341f
C129 VTAIL.n81 VSUBS 0.013144f
C130 VTAIL.n82 VSUBS 0.012414f
C131 VTAIL.n83 VSUBS 0.023101f
C132 VTAIL.n84 VSUBS 0.023101f
C133 VTAIL.n85 VSUBS 0.012414f
C134 VTAIL.n86 VSUBS 0.013144f
C135 VTAIL.n87 VSUBS 0.029341f
C136 VTAIL.n88 VSUBS 0.067701f
C137 VTAIL.n89 VSUBS 0.013144f
C138 VTAIL.n90 VSUBS 0.012414f
C139 VTAIL.n91 VSUBS 0.053082f
C140 VTAIL.n92 VSUBS 0.033889f
C141 VTAIL.n93 VSUBS 0.182064f
C142 VTAIL.n94 VSUBS 0.024405f
C143 VTAIL.n95 VSUBS 0.023101f
C144 VTAIL.n96 VSUBS 0.012414f
C145 VTAIL.n97 VSUBS 0.029341f
C146 VTAIL.n98 VSUBS 0.013144f
C147 VTAIL.n99 VSUBS 0.023101f
C148 VTAIL.n100 VSUBS 0.012414f
C149 VTAIL.n101 VSUBS 0.029341f
C150 VTAIL.n102 VSUBS 0.013144f
C151 VTAIL.n103 VSUBS 0.023101f
C152 VTAIL.n104 VSUBS 0.012414f
C153 VTAIL.n105 VSUBS 0.029341f
C154 VTAIL.n106 VSUBS 0.013144f
C155 VTAIL.n107 VSUBS 0.023101f
C156 VTAIL.n108 VSUBS 0.012414f
C157 VTAIL.n109 VSUBS 0.029341f
C158 VTAIL.n110 VSUBS 0.013144f
C159 VTAIL.n111 VSUBS 0.023101f
C160 VTAIL.n112 VSUBS 0.012414f
C161 VTAIL.n113 VSUBS 0.029341f
C162 VTAIL.n114 VSUBS 0.013144f
C163 VTAIL.n115 VSUBS 0.023101f
C164 VTAIL.n116 VSUBS 0.012414f
C165 VTAIL.n117 VSUBS 0.029341f
C166 VTAIL.n118 VSUBS 0.013144f
C167 VTAIL.n119 VSUBS 0.023101f
C168 VTAIL.n120 VSUBS 0.012414f
C169 VTAIL.n121 VSUBS 0.029341f
C170 VTAIL.n122 VSUBS 0.013144f
C171 VTAIL.n123 VSUBS 0.175041f
C172 VTAIL.t5 VSUBS 0.062917f
C173 VTAIL.n124 VSUBS 0.022006f
C174 VTAIL.n125 VSUBS 0.018666f
C175 VTAIL.n126 VSUBS 0.012414f
C176 VTAIL.n127 VSUBS 1.66279f
C177 VTAIL.n128 VSUBS 0.023101f
C178 VTAIL.n129 VSUBS 0.012414f
C179 VTAIL.n130 VSUBS 0.013144f
C180 VTAIL.n131 VSUBS 0.029341f
C181 VTAIL.n132 VSUBS 0.029341f
C182 VTAIL.n133 VSUBS 0.013144f
C183 VTAIL.n134 VSUBS 0.012414f
C184 VTAIL.n135 VSUBS 0.023101f
C185 VTAIL.n136 VSUBS 0.023101f
C186 VTAIL.n137 VSUBS 0.012414f
C187 VTAIL.n138 VSUBS 0.013144f
C188 VTAIL.n139 VSUBS 0.029341f
C189 VTAIL.n140 VSUBS 0.029341f
C190 VTAIL.n141 VSUBS 0.013144f
C191 VTAIL.n142 VSUBS 0.012414f
C192 VTAIL.n143 VSUBS 0.023101f
C193 VTAIL.n144 VSUBS 0.023101f
C194 VTAIL.n145 VSUBS 0.012414f
C195 VTAIL.n146 VSUBS 0.013144f
C196 VTAIL.n147 VSUBS 0.029341f
C197 VTAIL.n148 VSUBS 0.029341f
C198 VTAIL.n149 VSUBS 0.013144f
C199 VTAIL.n150 VSUBS 0.012414f
C200 VTAIL.n151 VSUBS 0.023101f
C201 VTAIL.n152 VSUBS 0.023101f
C202 VTAIL.n153 VSUBS 0.012414f
C203 VTAIL.n154 VSUBS 0.013144f
C204 VTAIL.n155 VSUBS 0.029341f
C205 VTAIL.n156 VSUBS 0.029341f
C206 VTAIL.n157 VSUBS 0.013144f
C207 VTAIL.n158 VSUBS 0.012414f
C208 VTAIL.n159 VSUBS 0.023101f
C209 VTAIL.n160 VSUBS 0.023101f
C210 VTAIL.n161 VSUBS 0.012414f
C211 VTAIL.n162 VSUBS 0.013144f
C212 VTAIL.n163 VSUBS 0.029341f
C213 VTAIL.n164 VSUBS 0.029341f
C214 VTAIL.n165 VSUBS 0.029341f
C215 VTAIL.n166 VSUBS 0.013144f
C216 VTAIL.n167 VSUBS 0.012414f
C217 VTAIL.n168 VSUBS 0.023101f
C218 VTAIL.n169 VSUBS 0.023101f
C219 VTAIL.n170 VSUBS 0.012414f
C220 VTAIL.n171 VSUBS 0.012779f
C221 VTAIL.n172 VSUBS 0.012779f
C222 VTAIL.n173 VSUBS 0.029341f
C223 VTAIL.n174 VSUBS 0.029341f
C224 VTAIL.n175 VSUBS 0.013144f
C225 VTAIL.n176 VSUBS 0.012414f
C226 VTAIL.n177 VSUBS 0.023101f
C227 VTAIL.n178 VSUBS 0.023101f
C228 VTAIL.n179 VSUBS 0.012414f
C229 VTAIL.n180 VSUBS 0.013144f
C230 VTAIL.n181 VSUBS 0.029341f
C231 VTAIL.n182 VSUBS 0.067701f
C232 VTAIL.n183 VSUBS 0.013144f
C233 VTAIL.n184 VSUBS 0.012414f
C234 VTAIL.n185 VSUBS 0.053082f
C235 VTAIL.n186 VSUBS 0.033889f
C236 VTAIL.n187 VSUBS 0.300939f
C237 VTAIL.n188 VSUBS 0.024405f
C238 VTAIL.n189 VSUBS 0.023101f
C239 VTAIL.n190 VSUBS 0.012414f
C240 VTAIL.n191 VSUBS 0.029341f
C241 VTAIL.n192 VSUBS 0.013144f
C242 VTAIL.n193 VSUBS 0.023101f
C243 VTAIL.n194 VSUBS 0.012414f
C244 VTAIL.n195 VSUBS 0.029341f
C245 VTAIL.n196 VSUBS 0.013144f
C246 VTAIL.n197 VSUBS 0.023101f
C247 VTAIL.n198 VSUBS 0.012414f
C248 VTAIL.n199 VSUBS 0.029341f
C249 VTAIL.n200 VSUBS 0.013144f
C250 VTAIL.n201 VSUBS 0.023101f
C251 VTAIL.n202 VSUBS 0.012414f
C252 VTAIL.n203 VSUBS 0.029341f
C253 VTAIL.n204 VSUBS 0.013144f
C254 VTAIL.n205 VSUBS 0.023101f
C255 VTAIL.n206 VSUBS 0.012414f
C256 VTAIL.n207 VSUBS 0.029341f
C257 VTAIL.n208 VSUBS 0.013144f
C258 VTAIL.n209 VSUBS 0.023101f
C259 VTAIL.n210 VSUBS 0.012414f
C260 VTAIL.n211 VSUBS 0.029341f
C261 VTAIL.n212 VSUBS 0.013144f
C262 VTAIL.n213 VSUBS 0.023101f
C263 VTAIL.n214 VSUBS 0.012414f
C264 VTAIL.n215 VSUBS 0.029341f
C265 VTAIL.n216 VSUBS 0.013144f
C266 VTAIL.n217 VSUBS 0.175041f
C267 VTAIL.t4 VSUBS 0.062917f
C268 VTAIL.n218 VSUBS 0.022006f
C269 VTAIL.n219 VSUBS 0.018666f
C270 VTAIL.n220 VSUBS 0.012414f
C271 VTAIL.n221 VSUBS 1.66279f
C272 VTAIL.n222 VSUBS 0.023101f
C273 VTAIL.n223 VSUBS 0.012414f
C274 VTAIL.n224 VSUBS 0.013144f
C275 VTAIL.n225 VSUBS 0.029341f
C276 VTAIL.n226 VSUBS 0.029341f
C277 VTAIL.n227 VSUBS 0.013144f
C278 VTAIL.n228 VSUBS 0.012414f
C279 VTAIL.n229 VSUBS 0.023101f
C280 VTAIL.n230 VSUBS 0.023101f
C281 VTAIL.n231 VSUBS 0.012414f
C282 VTAIL.n232 VSUBS 0.013144f
C283 VTAIL.n233 VSUBS 0.029341f
C284 VTAIL.n234 VSUBS 0.029341f
C285 VTAIL.n235 VSUBS 0.013144f
C286 VTAIL.n236 VSUBS 0.012414f
C287 VTAIL.n237 VSUBS 0.023101f
C288 VTAIL.n238 VSUBS 0.023101f
C289 VTAIL.n239 VSUBS 0.012414f
C290 VTAIL.n240 VSUBS 0.013144f
C291 VTAIL.n241 VSUBS 0.029341f
C292 VTAIL.n242 VSUBS 0.029341f
C293 VTAIL.n243 VSUBS 0.013144f
C294 VTAIL.n244 VSUBS 0.012414f
C295 VTAIL.n245 VSUBS 0.023101f
C296 VTAIL.n246 VSUBS 0.023101f
C297 VTAIL.n247 VSUBS 0.012414f
C298 VTAIL.n248 VSUBS 0.013144f
C299 VTAIL.n249 VSUBS 0.029341f
C300 VTAIL.n250 VSUBS 0.029341f
C301 VTAIL.n251 VSUBS 0.013144f
C302 VTAIL.n252 VSUBS 0.012414f
C303 VTAIL.n253 VSUBS 0.023101f
C304 VTAIL.n254 VSUBS 0.023101f
C305 VTAIL.n255 VSUBS 0.012414f
C306 VTAIL.n256 VSUBS 0.013144f
C307 VTAIL.n257 VSUBS 0.029341f
C308 VTAIL.n258 VSUBS 0.029341f
C309 VTAIL.n259 VSUBS 0.029341f
C310 VTAIL.n260 VSUBS 0.013144f
C311 VTAIL.n261 VSUBS 0.012414f
C312 VTAIL.n262 VSUBS 0.023101f
C313 VTAIL.n263 VSUBS 0.023101f
C314 VTAIL.n264 VSUBS 0.012414f
C315 VTAIL.n265 VSUBS 0.012779f
C316 VTAIL.n266 VSUBS 0.012779f
C317 VTAIL.n267 VSUBS 0.029341f
C318 VTAIL.n268 VSUBS 0.029341f
C319 VTAIL.n269 VSUBS 0.013144f
C320 VTAIL.n270 VSUBS 0.012414f
C321 VTAIL.n271 VSUBS 0.023101f
C322 VTAIL.n272 VSUBS 0.023101f
C323 VTAIL.n273 VSUBS 0.012414f
C324 VTAIL.n274 VSUBS 0.013144f
C325 VTAIL.n275 VSUBS 0.029341f
C326 VTAIL.n276 VSUBS 0.067701f
C327 VTAIL.n277 VSUBS 0.013144f
C328 VTAIL.n278 VSUBS 0.012414f
C329 VTAIL.n279 VSUBS 0.053082f
C330 VTAIL.n280 VSUBS 0.033889f
C331 VTAIL.n281 VSUBS 1.90361f
C332 VTAIL.n282 VSUBS 0.024405f
C333 VTAIL.n283 VSUBS 0.023101f
C334 VTAIL.n284 VSUBS 0.012414f
C335 VTAIL.n285 VSUBS 0.029341f
C336 VTAIL.n286 VSUBS 0.013144f
C337 VTAIL.n287 VSUBS 0.023101f
C338 VTAIL.n288 VSUBS 0.012414f
C339 VTAIL.n289 VSUBS 0.029341f
C340 VTAIL.n290 VSUBS 0.013144f
C341 VTAIL.n291 VSUBS 0.023101f
C342 VTAIL.n292 VSUBS 0.012414f
C343 VTAIL.n293 VSUBS 0.029341f
C344 VTAIL.n294 VSUBS 0.029341f
C345 VTAIL.n295 VSUBS 0.013144f
C346 VTAIL.n296 VSUBS 0.023101f
C347 VTAIL.n297 VSUBS 0.012414f
C348 VTAIL.n298 VSUBS 0.029341f
C349 VTAIL.n299 VSUBS 0.013144f
C350 VTAIL.n300 VSUBS 0.023101f
C351 VTAIL.n301 VSUBS 0.012414f
C352 VTAIL.n302 VSUBS 0.029341f
C353 VTAIL.n303 VSUBS 0.013144f
C354 VTAIL.n304 VSUBS 0.023101f
C355 VTAIL.n305 VSUBS 0.012414f
C356 VTAIL.n306 VSUBS 0.029341f
C357 VTAIL.n307 VSUBS 0.013144f
C358 VTAIL.n308 VSUBS 0.023101f
C359 VTAIL.n309 VSUBS 0.012414f
C360 VTAIL.n310 VSUBS 0.029341f
C361 VTAIL.n311 VSUBS 0.013144f
C362 VTAIL.n312 VSUBS 0.175041f
C363 VTAIL.t1 VSUBS 0.062917f
C364 VTAIL.n313 VSUBS 0.022006f
C365 VTAIL.n314 VSUBS 0.018666f
C366 VTAIL.n315 VSUBS 0.012414f
C367 VTAIL.n316 VSUBS 1.66279f
C368 VTAIL.n317 VSUBS 0.023101f
C369 VTAIL.n318 VSUBS 0.012414f
C370 VTAIL.n319 VSUBS 0.013144f
C371 VTAIL.n320 VSUBS 0.029341f
C372 VTAIL.n321 VSUBS 0.029341f
C373 VTAIL.n322 VSUBS 0.013144f
C374 VTAIL.n323 VSUBS 0.012414f
C375 VTAIL.n324 VSUBS 0.023101f
C376 VTAIL.n325 VSUBS 0.023101f
C377 VTAIL.n326 VSUBS 0.012414f
C378 VTAIL.n327 VSUBS 0.013144f
C379 VTAIL.n328 VSUBS 0.029341f
C380 VTAIL.n329 VSUBS 0.029341f
C381 VTAIL.n330 VSUBS 0.013144f
C382 VTAIL.n331 VSUBS 0.012414f
C383 VTAIL.n332 VSUBS 0.023101f
C384 VTAIL.n333 VSUBS 0.023101f
C385 VTAIL.n334 VSUBS 0.012414f
C386 VTAIL.n335 VSUBS 0.013144f
C387 VTAIL.n336 VSUBS 0.029341f
C388 VTAIL.n337 VSUBS 0.029341f
C389 VTAIL.n338 VSUBS 0.013144f
C390 VTAIL.n339 VSUBS 0.012414f
C391 VTAIL.n340 VSUBS 0.023101f
C392 VTAIL.n341 VSUBS 0.023101f
C393 VTAIL.n342 VSUBS 0.012414f
C394 VTAIL.n343 VSUBS 0.013144f
C395 VTAIL.n344 VSUBS 0.029341f
C396 VTAIL.n345 VSUBS 0.029341f
C397 VTAIL.n346 VSUBS 0.013144f
C398 VTAIL.n347 VSUBS 0.012414f
C399 VTAIL.n348 VSUBS 0.023101f
C400 VTAIL.n349 VSUBS 0.023101f
C401 VTAIL.n350 VSUBS 0.012414f
C402 VTAIL.n351 VSUBS 0.013144f
C403 VTAIL.n352 VSUBS 0.029341f
C404 VTAIL.n353 VSUBS 0.029341f
C405 VTAIL.n354 VSUBS 0.013144f
C406 VTAIL.n355 VSUBS 0.012414f
C407 VTAIL.n356 VSUBS 0.023101f
C408 VTAIL.n357 VSUBS 0.023101f
C409 VTAIL.n358 VSUBS 0.012414f
C410 VTAIL.n359 VSUBS 0.012779f
C411 VTAIL.n360 VSUBS 0.012779f
C412 VTAIL.n361 VSUBS 0.029341f
C413 VTAIL.n362 VSUBS 0.029341f
C414 VTAIL.n363 VSUBS 0.013144f
C415 VTAIL.n364 VSUBS 0.012414f
C416 VTAIL.n365 VSUBS 0.023101f
C417 VTAIL.n366 VSUBS 0.023101f
C418 VTAIL.n367 VSUBS 0.012414f
C419 VTAIL.n368 VSUBS 0.013144f
C420 VTAIL.n369 VSUBS 0.029341f
C421 VTAIL.n370 VSUBS 0.067701f
C422 VTAIL.n371 VSUBS 0.013144f
C423 VTAIL.n372 VSUBS 0.012414f
C424 VTAIL.n373 VSUBS 0.053082f
C425 VTAIL.n374 VSUBS 0.033889f
C426 VTAIL.n375 VSUBS 1.90361f
C427 VTAIL.n376 VSUBS 0.024405f
C428 VTAIL.n377 VSUBS 0.023101f
C429 VTAIL.n378 VSUBS 0.012414f
C430 VTAIL.n379 VSUBS 0.029341f
C431 VTAIL.n380 VSUBS 0.013144f
C432 VTAIL.n381 VSUBS 0.023101f
C433 VTAIL.n382 VSUBS 0.012414f
C434 VTAIL.n383 VSUBS 0.029341f
C435 VTAIL.n384 VSUBS 0.013144f
C436 VTAIL.n385 VSUBS 0.023101f
C437 VTAIL.n386 VSUBS 0.012414f
C438 VTAIL.n387 VSUBS 0.029341f
C439 VTAIL.n388 VSUBS 0.029341f
C440 VTAIL.n389 VSUBS 0.013144f
C441 VTAIL.n390 VSUBS 0.023101f
C442 VTAIL.n391 VSUBS 0.012414f
C443 VTAIL.n392 VSUBS 0.029341f
C444 VTAIL.n393 VSUBS 0.013144f
C445 VTAIL.n394 VSUBS 0.023101f
C446 VTAIL.n395 VSUBS 0.012414f
C447 VTAIL.n396 VSUBS 0.029341f
C448 VTAIL.n397 VSUBS 0.013144f
C449 VTAIL.n398 VSUBS 0.023101f
C450 VTAIL.n399 VSUBS 0.012414f
C451 VTAIL.n400 VSUBS 0.029341f
C452 VTAIL.n401 VSUBS 0.013144f
C453 VTAIL.n402 VSUBS 0.023101f
C454 VTAIL.n403 VSUBS 0.012414f
C455 VTAIL.n404 VSUBS 0.029341f
C456 VTAIL.n405 VSUBS 0.013144f
C457 VTAIL.n406 VSUBS 0.175041f
C458 VTAIL.t3 VSUBS 0.062917f
C459 VTAIL.n407 VSUBS 0.022006f
C460 VTAIL.n408 VSUBS 0.018666f
C461 VTAIL.n409 VSUBS 0.012414f
C462 VTAIL.n410 VSUBS 1.66279f
C463 VTAIL.n411 VSUBS 0.023101f
C464 VTAIL.n412 VSUBS 0.012414f
C465 VTAIL.n413 VSUBS 0.013144f
C466 VTAIL.n414 VSUBS 0.029341f
C467 VTAIL.n415 VSUBS 0.029341f
C468 VTAIL.n416 VSUBS 0.013144f
C469 VTAIL.n417 VSUBS 0.012414f
C470 VTAIL.n418 VSUBS 0.023101f
C471 VTAIL.n419 VSUBS 0.023101f
C472 VTAIL.n420 VSUBS 0.012414f
C473 VTAIL.n421 VSUBS 0.013144f
C474 VTAIL.n422 VSUBS 0.029341f
C475 VTAIL.n423 VSUBS 0.029341f
C476 VTAIL.n424 VSUBS 0.013144f
C477 VTAIL.n425 VSUBS 0.012414f
C478 VTAIL.n426 VSUBS 0.023101f
C479 VTAIL.n427 VSUBS 0.023101f
C480 VTAIL.n428 VSUBS 0.012414f
C481 VTAIL.n429 VSUBS 0.013144f
C482 VTAIL.n430 VSUBS 0.029341f
C483 VTAIL.n431 VSUBS 0.029341f
C484 VTAIL.n432 VSUBS 0.013144f
C485 VTAIL.n433 VSUBS 0.012414f
C486 VTAIL.n434 VSUBS 0.023101f
C487 VTAIL.n435 VSUBS 0.023101f
C488 VTAIL.n436 VSUBS 0.012414f
C489 VTAIL.n437 VSUBS 0.013144f
C490 VTAIL.n438 VSUBS 0.029341f
C491 VTAIL.n439 VSUBS 0.029341f
C492 VTAIL.n440 VSUBS 0.013144f
C493 VTAIL.n441 VSUBS 0.012414f
C494 VTAIL.n442 VSUBS 0.023101f
C495 VTAIL.n443 VSUBS 0.023101f
C496 VTAIL.n444 VSUBS 0.012414f
C497 VTAIL.n445 VSUBS 0.013144f
C498 VTAIL.n446 VSUBS 0.029341f
C499 VTAIL.n447 VSUBS 0.029341f
C500 VTAIL.n448 VSUBS 0.013144f
C501 VTAIL.n449 VSUBS 0.012414f
C502 VTAIL.n450 VSUBS 0.023101f
C503 VTAIL.n451 VSUBS 0.023101f
C504 VTAIL.n452 VSUBS 0.012414f
C505 VTAIL.n453 VSUBS 0.012779f
C506 VTAIL.n454 VSUBS 0.012779f
C507 VTAIL.n455 VSUBS 0.029341f
C508 VTAIL.n456 VSUBS 0.029341f
C509 VTAIL.n457 VSUBS 0.013144f
C510 VTAIL.n458 VSUBS 0.012414f
C511 VTAIL.n459 VSUBS 0.023101f
C512 VTAIL.n460 VSUBS 0.023101f
C513 VTAIL.n461 VSUBS 0.012414f
C514 VTAIL.n462 VSUBS 0.013144f
C515 VTAIL.n463 VSUBS 0.029341f
C516 VTAIL.n464 VSUBS 0.067701f
C517 VTAIL.n465 VSUBS 0.013144f
C518 VTAIL.n466 VSUBS 0.012414f
C519 VTAIL.n467 VSUBS 0.053082f
C520 VTAIL.n468 VSUBS 0.033889f
C521 VTAIL.n469 VSUBS 0.300939f
C522 VTAIL.n470 VSUBS 0.024405f
C523 VTAIL.n471 VSUBS 0.023101f
C524 VTAIL.n472 VSUBS 0.012414f
C525 VTAIL.n473 VSUBS 0.029341f
C526 VTAIL.n474 VSUBS 0.013144f
C527 VTAIL.n475 VSUBS 0.023101f
C528 VTAIL.n476 VSUBS 0.012414f
C529 VTAIL.n477 VSUBS 0.029341f
C530 VTAIL.n478 VSUBS 0.013144f
C531 VTAIL.n479 VSUBS 0.023101f
C532 VTAIL.n480 VSUBS 0.012414f
C533 VTAIL.n481 VSUBS 0.029341f
C534 VTAIL.n482 VSUBS 0.029341f
C535 VTAIL.n483 VSUBS 0.013144f
C536 VTAIL.n484 VSUBS 0.023101f
C537 VTAIL.n485 VSUBS 0.012414f
C538 VTAIL.n486 VSUBS 0.029341f
C539 VTAIL.n487 VSUBS 0.013144f
C540 VTAIL.n488 VSUBS 0.023101f
C541 VTAIL.n489 VSUBS 0.012414f
C542 VTAIL.n490 VSUBS 0.029341f
C543 VTAIL.n491 VSUBS 0.013144f
C544 VTAIL.n492 VSUBS 0.023101f
C545 VTAIL.n493 VSUBS 0.012414f
C546 VTAIL.n494 VSUBS 0.029341f
C547 VTAIL.n495 VSUBS 0.013144f
C548 VTAIL.n496 VSUBS 0.023101f
C549 VTAIL.n497 VSUBS 0.012414f
C550 VTAIL.n498 VSUBS 0.029341f
C551 VTAIL.n499 VSUBS 0.013144f
C552 VTAIL.n500 VSUBS 0.175041f
C553 VTAIL.t6 VSUBS 0.062917f
C554 VTAIL.n501 VSUBS 0.022006f
C555 VTAIL.n502 VSUBS 0.018666f
C556 VTAIL.n503 VSUBS 0.012414f
C557 VTAIL.n504 VSUBS 1.66279f
C558 VTAIL.n505 VSUBS 0.023101f
C559 VTAIL.n506 VSUBS 0.012414f
C560 VTAIL.n507 VSUBS 0.013144f
C561 VTAIL.n508 VSUBS 0.029341f
C562 VTAIL.n509 VSUBS 0.029341f
C563 VTAIL.n510 VSUBS 0.013144f
C564 VTAIL.n511 VSUBS 0.012414f
C565 VTAIL.n512 VSUBS 0.023101f
C566 VTAIL.n513 VSUBS 0.023101f
C567 VTAIL.n514 VSUBS 0.012414f
C568 VTAIL.n515 VSUBS 0.013144f
C569 VTAIL.n516 VSUBS 0.029341f
C570 VTAIL.n517 VSUBS 0.029341f
C571 VTAIL.n518 VSUBS 0.013144f
C572 VTAIL.n519 VSUBS 0.012414f
C573 VTAIL.n520 VSUBS 0.023101f
C574 VTAIL.n521 VSUBS 0.023101f
C575 VTAIL.n522 VSUBS 0.012414f
C576 VTAIL.n523 VSUBS 0.013144f
C577 VTAIL.n524 VSUBS 0.029341f
C578 VTAIL.n525 VSUBS 0.029341f
C579 VTAIL.n526 VSUBS 0.013144f
C580 VTAIL.n527 VSUBS 0.012414f
C581 VTAIL.n528 VSUBS 0.023101f
C582 VTAIL.n529 VSUBS 0.023101f
C583 VTAIL.n530 VSUBS 0.012414f
C584 VTAIL.n531 VSUBS 0.013144f
C585 VTAIL.n532 VSUBS 0.029341f
C586 VTAIL.n533 VSUBS 0.029341f
C587 VTAIL.n534 VSUBS 0.013144f
C588 VTAIL.n535 VSUBS 0.012414f
C589 VTAIL.n536 VSUBS 0.023101f
C590 VTAIL.n537 VSUBS 0.023101f
C591 VTAIL.n538 VSUBS 0.012414f
C592 VTAIL.n539 VSUBS 0.013144f
C593 VTAIL.n540 VSUBS 0.029341f
C594 VTAIL.n541 VSUBS 0.029341f
C595 VTAIL.n542 VSUBS 0.013144f
C596 VTAIL.n543 VSUBS 0.012414f
C597 VTAIL.n544 VSUBS 0.023101f
C598 VTAIL.n545 VSUBS 0.023101f
C599 VTAIL.n546 VSUBS 0.012414f
C600 VTAIL.n547 VSUBS 0.012779f
C601 VTAIL.n548 VSUBS 0.012779f
C602 VTAIL.n549 VSUBS 0.029341f
C603 VTAIL.n550 VSUBS 0.029341f
C604 VTAIL.n551 VSUBS 0.013144f
C605 VTAIL.n552 VSUBS 0.012414f
C606 VTAIL.n553 VSUBS 0.023101f
C607 VTAIL.n554 VSUBS 0.023101f
C608 VTAIL.n555 VSUBS 0.012414f
C609 VTAIL.n556 VSUBS 0.013144f
C610 VTAIL.n557 VSUBS 0.029341f
C611 VTAIL.n558 VSUBS 0.067701f
C612 VTAIL.n559 VSUBS 0.013144f
C613 VTAIL.n560 VSUBS 0.012414f
C614 VTAIL.n561 VSUBS 0.053082f
C615 VTAIL.n562 VSUBS 0.033889f
C616 VTAIL.n563 VSUBS 0.300939f
C617 VTAIL.n564 VSUBS 0.024405f
C618 VTAIL.n565 VSUBS 0.023101f
C619 VTAIL.n566 VSUBS 0.012414f
C620 VTAIL.n567 VSUBS 0.029341f
C621 VTAIL.n568 VSUBS 0.013144f
C622 VTAIL.n569 VSUBS 0.023101f
C623 VTAIL.n570 VSUBS 0.012414f
C624 VTAIL.n571 VSUBS 0.029341f
C625 VTAIL.n572 VSUBS 0.013144f
C626 VTAIL.n573 VSUBS 0.023101f
C627 VTAIL.n574 VSUBS 0.012414f
C628 VTAIL.n575 VSUBS 0.029341f
C629 VTAIL.n576 VSUBS 0.029341f
C630 VTAIL.n577 VSUBS 0.013144f
C631 VTAIL.n578 VSUBS 0.023101f
C632 VTAIL.n579 VSUBS 0.012414f
C633 VTAIL.n580 VSUBS 0.029341f
C634 VTAIL.n581 VSUBS 0.013144f
C635 VTAIL.n582 VSUBS 0.023101f
C636 VTAIL.n583 VSUBS 0.012414f
C637 VTAIL.n584 VSUBS 0.029341f
C638 VTAIL.n585 VSUBS 0.013144f
C639 VTAIL.n586 VSUBS 0.023101f
C640 VTAIL.n587 VSUBS 0.012414f
C641 VTAIL.n588 VSUBS 0.029341f
C642 VTAIL.n589 VSUBS 0.013144f
C643 VTAIL.n590 VSUBS 0.023101f
C644 VTAIL.n591 VSUBS 0.012414f
C645 VTAIL.n592 VSUBS 0.029341f
C646 VTAIL.n593 VSUBS 0.013144f
C647 VTAIL.n594 VSUBS 0.175041f
C648 VTAIL.t7 VSUBS 0.062917f
C649 VTAIL.n595 VSUBS 0.022006f
C650 VTAIL.n596 VSUBS 0.018666f
C651 VTAIL.n597 VSUBS 0.012414f
C652 VTAIL.n598 VSUBS 1.66279f
C653 VTAIL.n599 VSUBS 0.023101f
C654 VTAIL.n600 VSUBS 0.012414f
C655 VTAIL.n601 VSUBS 0.013144f
C656 VTAIL.n602 VSUBS 0.029341f
C657 VTAIL.n603 VSUBS 0.029341f
C658 VTAIL.n604 VSUBS 0.013144f
C659 VTAIL.n605 VSUBS 0.012414f
C660 VTAIL.n606 VSUBS 0.023101f
C661 VTAIL.n607 VSUBS 0.023101f
C662 VTAIL.n608 VSUBS 0.012414f
C663 VTAIL.n609 VSUBS 0.013144f
C664 VTAIL.n610 VSUBS 0.029341f
C665 VTAIL.n611 VSUBS 0.029341f
C666 VTAIL.n612 VSUBS 0.013144f
C667 VTAIL.n613 VSUBS 0.012414f
C668 VTAIL.n614 VSUBS 0.023101f
C669 VTAIL.n615 VSUBS 0.023101f
C670 VTAIL.n616 VSUBS 0.012414f
C671 VTAIL.n617 VSUBS 0.013144f
C672 VTAIL.n618 VSUBS 0.029341f
C673 VTAIL.n619 VSUBS 0.029341f
C674 VTAIL.n620 VSUBS 0.013144f
C675 VTAIL.n621 VSUBS 0.012414f
C676 VTAIL.n622 VSUBS 0.023101f
C677 VTAIL.n623 VSUBS 0.023101f
C678 VTAIL.n624 VSUBS 0.012414f
C679 VTAIL.n625 VSUBS 0.013144f
C680 VTAIL.n626 VSUBS 0.029341f
C681 VTAIL.n627 VSUBS 0.029341f
C682 VTAIL.n628 VSUBS 0.013144f
C683 VTAIL.n629 VSUBS 0.012414f
C684 VTAIL.n630 VSUBS 0.023101f
C685 VTAIL.n631 VSUBS 0.023101f
C686 VTAIL.n632 VSUBS 0.012414f
C687 VTAIL.n633 VSUBS 0.013144f
C688 VTAIL.n634 VSUBS 0.029341f
C689 VTAIL.n635 VSUBS 0.029341f
C690 VTAIL.n636 VSUBS 0.013144f
C691 VTAIL.n637 VSUBS 0.012414f
C692 VTAIL.n638 VSUBS 0.023101f
C693 VTAIL.n639 VSUBS 0.023101f
C694 VTAIL.n640 VSUBS 0.012414f
C695 VTAIL.n641 VSUBS 0.012779f
C696 VTAIL.n642 VSUBS 0.012779f
C697 VTAIL.n643 VSUBS 0.029341f
C698 VTAIL.n644 VSUBS 0.029341f
C699 VTAIL.n645 VSUBS 0.013144f
C700 VTAIL.n646 VSUBS 0.012414f
C701 VTAIL.n647 VSUBS 0.023101f
C702 VTAIL.n648 VSUBS 0.023101f
C703 VTAIL.n649 VSUBS 0.012414f
C704 VTAIL.n650 VSUBS 0.013144f
C705 VTAIL.n651 VSUBS 0.029341f
C706 VTAIL.n652 VSUBS 0.067701f
C707 VTAIL.n653 VSUBS 0.013144f
C708 VTAIL.n654 VSUBS 0.012414f
C709 VTAIL.n655 VSUBS 0.053082f
C710 VTAIL.n656 VSUBS 0.033889f
C711 VTAIL.n657 VSUBS 1.90361f
C712 VTAIL.n658 VSUBS 0.024405f
C713 VTAIL.n659 VSUBS 0.023101f
C714 VTAIL.n660 VSUBS 0.012414f
C715 VTAIL.n661 VSUBS 0.029341f
C716 VTAIL.n662 VSUBS 0.013144f
C717 VTAIL.n663 VSUBS 0.023101f
C718 VTAIL.n664 VSUBS 0.012414f
C719 VTAIL.n665 VSUBS 0.029341f
C720 VTAIL.n666 VSUBS 0.013144f
C721 VTAIL.n667 VSUBS 0.023101f
C722 VTAIL.n668 VSUBS 0.012414f
C723 VTAIL.n669 VSUBS 0.029341f
C724 VTAIL.n670 VSUBS 0.013144f
C725 VTAIL.n671 VSUBS 0.023101f
C726 VTAIL.n672 VSUBS 0.012414f
C727 VTAIL.n673 VSUBS 0.029341f
C728 VTAIL.n674 VSUBS 0.013144f
C729 VTAIL.n675 VSUBS 0.023101f
C730 VTAIL.n676 VSUBS 0.012414f
C731 VTAIL.n677 VSUBS 0.029341f
C732 VTAIL.n678 VSUBS 0.013144f
C733 VTAIL.n679 VSUBS 0.023101f
C734 VTAIL.n680 VSUBS 0.012414f
C735 VTAIL.n681 VSUBS 0.029341f
C736 VTAIL.n682 VSUBS 0.013144f
C737 VTAIL.n683 VSUBS 0.023101f
C738 VTAIL.n684 VSUBS 0.012414f
C739 VTAIL.n685 VSUBS 0.029341f
C740 VTAIL.n686 VSUBS 0.013144f
C741 VTAIL.n687 VSUBS 0.175041f
C742 VTAIL.t0 VSUBS 0.062917f
C743 VTAIL.n688 VSUBS 0.022006f
C744 VTAIL.n689 VSUBS 0.018666f
C745 VTAIL.n690 VSUBS 0.012414f
C746 VTAIL.n691 VSUBS 1.66279f
C747 VTAIL.n692 VSUBS 0.023101f
C748 VTAIL.n693 VSUBS 0.012414f
C749 VTAIL.n694 VSUBS 0.013144f
C750 VTAIL.n695 VSUBS 0.029341f
C751 VTAIL.n696 VSUBS 0.029341f
C752 VTAIL.n697 VSUBS 0.013144f
C753 VTAIL.n698 VSUBS 0.012414f
C754 VTAIL.n699 VSUBS 0.023101f
C755 VTAIL.n700 VSUBS 0.023101f
C756 VTAIL.n701 VSUBS 0.012414f
C757 VTAIL.n702 VSUBS 0.013144f
C758 VTAIL.n703 VSUBS 0.029341f
C759 VTAIL.n704 VSUBS 0.029341f
C760 VTAIL.n705 VSUBS 0.013144f
C761 VTAIL.n706 VSUBS 0.012414f
C762 VTAIL.n707 VSUBS 0.023101f
C763 VTAIL.n708 VSUBS 0.023101f
C764 VTAIL.n709 VSUBS 0.012414f
C765 VTAIL.n710 VSUBS 0.013144f
C766 VTAIL.n711 VSUBS 0.029341f
C767 VTAIL.n712 VSUBS 0.029341f
C768 VTAIL.n713 VSUBS 0.013144f
C769 VTAIL.n714 VSUBS 0.012414f
C770 VTAIL.n715 VSUBS 0.023101f
C771 VTAIL.n716 VSUBS 0.023101f
C772 VTAIL.n717 VSUBS 0.012414f
C773 VTAIL.n718 VSUBS 0.013144f
C774 VTAIL.n719 VSUBS 0.029341f
C775 VTAIL.n720 VSUBS 0.029341f
C776 VTAIL.n721 VSUBS 0.013144f
C777 VTAIL.n722 VSUBS 0.012414f
C778 VTAIL.n723 VSUBS 0.023101f
C779 VTAIL.n724 VSUBS 0.023101f
C780 VTAIL.n725 VSUBS 0.012414f
C781 VTAIL.n726 VSUBS 0.013144f
C782 VTAIL.n727 VSUBS 0.029341f
C783 VTAIL.n728 VSUBS 0.029341f
C784 VTAIL.n729 VSUBS 0.029341f
C785 VTAIL.n730 VSUBS 0.013144f
C786 VTAIL.n731 VSUBS 0.012414f
C787 VTAIL.n732 VSUBS 0.023101f
C788 VTAIL.n733 VSUBS 0.023101f
C789 VTAIL.n734 VSUBS 0.012414f
C790 VTAIL.n735 VSUBS 0.012779f
C791 VTAIL.n736 VSUBS 0.012779f
C792 VTAIL.n737 VSUBS 0.029341f
C793 VTAIL.n738 VSUBS 0.029341f
C794 VTAIL.n739 VSUBS 0.013144f
C795 VTAIL.n740 VSUBS 0.012414f
C796 VTAIL.n741 VSUBS 0.023101f
C797 VTAIL.n742 VSUBS 0.023101f
C798 VTAIL.n743 VSUBS 0.012414f
C799 VTAIL.n744 VSUBS 0.013144f
C800 VTAIL.n745 VSUBS 0.029341f
C801 VTAIL.n746 VSUBS 0.067701f
C802 VTAIL.n747 VSUBS 0.013144f
C803 VTAIL.n748 VSUBS 0.012414f
C804 VTAIL.n749 VSUBS 0.053082f
C805 VTAIL.n750 VSUBS 0.033889f
C806 VTAIL.n751 VSUBS 1.77607f
C807 VP.t0 VSUBS 4.51345f
C808 VP.n0 VSUBS 1.66576f
C809 VP.n1 VSUBS 0.027882f
C810 VP.n2 VSUBS 0.040702f
C811 VP.n3 VSUBS 0.027882f
C812 VP.n4 VSUBS 0.035032f
C813 VP.t2 VSUBS 4.92285f
C814 VP.t1 VSUBS 4.9089f
C815 VP.n5 VSUBS 4.93702f
C816 VP.t3 VSUBS 4.51345f
C817 VP.n6 VSUBS 1.66576f
C818 VP.n7 VSUBS 1.82366f
C819 VP.n8 VSUBS 0.045001f
C820 VP.n9 VSUBS 0.027882f
C821 VP.n10 VSUBS 0.051965f
C822 VP.n11 VSUBS 0.051965f
C823 VP.n12 VSUBS 0.040702f
C824 VP.n13 VSUBS 0.027882f
C825 VP.n14 VSUBS 0.027882f
C826 VP.n15 VSUBS 0.027882f
C827 VP.n16 VSUBS 0.051965f
C828 VP.n17 VSUBS 0.051965f
C829 VP.n18 VSUBS 0.035032f
C830 VP.n19 VSUBS 0.045001f
C831 VP.n20 VSUBS 0.076634f
C832 B.n0 VSUBS 0.003976f
C833 B.n1 VSUBS 0.003976f
C834 B.n2 VSUBS 0.006288f
C835 B.n3 VSUBS 0.006288f
C836 B.n4 VSUBS 0.006288f
C837 B.n5 VSUBS 0.006288f
C838 B.n6 VSUBS 0.006288f
C839 B.n7 VSUBS 0.006288f
C840 B.n8 VSUBS 0.006288f
C841 B.n9 VSUBS 0.006288f
C842 B.n10 VSUBS 0.006288f
C843 B.n11 VSUBS 0.006288f
C844 B.n12 VSUBS 0.006288f
C845 B.n13 VSUBS 0.006288f
C846 B.n14 VSUBS 0.006288f
C847 B.n15 VSUBS 0.006288f
C848 B.n16 VSUBS 0.006288f
C849 B.n17 VSUBS 0.006288f
C850 B.n18 VSUBS 0.006288f
C851 B.n19 VSUBS 0.006288f
C852 B.n20 VSUBS 0.006288f
C853 B.n21 VSUBS 0.006288f
C854 B.n22 VSUBS 0.006288f
C855 B.n23 VSUBS 0.014967f
C856 B.n24 VSUBS 0.006288f
C857 B.n25 VSUBS 0.006288f
C858 B.n26 VSUBS 0.006288f
C859 B.n27 VSUBS 0.006288f
C860 B.n28 VSUBS 0.006288f
C861 B.n29 VSUBS 0.006288f
C862 B.n30 VSUBS 0.006288f
C863 B.n31 VSUBS 0.006288f
C864 B.n32 VSUBS 0.006288f
C865 B.n33 VSUBS 0.006288f
C866 B.n34 VSUBS 0.006288f
C867 B.n35 VSUBS 0.006288f
C868 B.n36 VSUBS 0.006288f
C869 B.n37 VSUBS 0.006288f
C870 B.n38 VSUBS 0.006288f
C871 B.n39 VSUBS 0.006288f
C872 B.n40 VSUBS 0.006288f
C873 B.n41 VSUBS 0.006288f
C874 B.n42 VSUBS 0.006288f
C875 B.n43 VSUBS 0.006288f
C876 B.n44 VSUBS 0.006288f
C877 B.n45 VSUBS 0.006288f
C878 B.n46 VSUBS 0.006288f
C879 B.n47 VSUBS 0.006288f
C880 B.n48 VSUBS 0.006288f
C881 B.n49 VSUBS 0.006288f
C882 B.n50 VSUBS 0.006288f
C883 B.n51 VSUBS 0.006288f
C884 B.t5 VSUBS 0.289161f
C885 B.t4 VSUBS 0.327567f
C886 B.t3 VSUBS 2.4098f
C887 B.n52 VSUBS 0.520105f
C888 B.n53 VSUBS 0.285553f
C889 B.n54 VSUBS 0.006288f
C890 B.n55 VSUBS 0.006288f
C891 B.n56 VSUBS 0.006288f
C892 B.n57 VSUBS 0.006288f
C893 B.t8 VSUBS 0.289164f
C894 B.t7 VSUBS 0.32757f
C895 B.t6 VSUBS 2.4098f
C896 B.n58 VSUBS 0.520102f
C897 B.n59 VSUBS 0.28555f
C898 B.n60 VSUBS 0.006288f
C899 B.n61 VSUBS 0.006288f
C900 B.n62 VSUBS 0.006288f
C901 B.n63 VSUBS 0.006288f
C902 B.n64 VSUBS 0.006288f
C903 B.n65 VSUBS 0.006288f
C904 B.n66 VSUBS 0.006288f
C905 B.n67 VSUBS 0.006288f
C906 B.n68 VSUBS 0.006288f
C907 B.n69 VSUBS 0.006288f
C908 B.n70 VSUBS 0.006288f
C909 B.n71 VSUBS 0.006288f
C910 B.n72 VSUBS 0.006288f
C911 B.n73 VSUBS 0.006288f
C912 B.n74 VSUBS 0.006288f
C913 B.n75 VSUBS 0.006288f
C914 B.n76 VSUBS 0.006288f
C915 B.n77 VSUBS 0.006288f
C916 B.n78 VSUBS 0.006288f
C917 B.n79 VSUBS 0.006288f
C918 B.n80 VSUBS 0.006288f
C919 B.n81 VSUBS 0.006288f
C920 B.n82 VSUBS 0.006288f
C921 B.n83 VSUBS 0.006288f
C922 B.n84 VSUBS 0.006288f
C923 B.n85 VSUBS 0.006288f
C924 B.n86 VSUBS 0.006288f
C925 B.n87 VSUBS 0.014967f
C926 B.n88 VSUBS 0.006288f
C927 B.n89 VSUBS 0.006288f
C928 B.n90 VSUBS 0.006288f
C929 B.n91 VSUBS 0.006288f
C930 B.n92 VSUBS 0.006288f
C931 B.n93 VSUBS 0.006288f
C932 B.n94 VSUBS 0.006288f
C933 B.n95 VSUBS 0.006288f
C934 B.n96 VSUBS 0.006288f
C935 B.n97 VSUBS 0.006288f
C936 B.n98 VSUBS 0.006288f
C937 B.n99 VSUBS 0.006288f
C938 B.n100 VSUBS 0.006288f
C939 B.n101 VSUBS 0.006288f
C940 B.n102 VSUBS 0.006288f
C941 B.n103 VSUBS 0.006288f
C942 B.n104 VSUBS 0.006288f
C943 B.n105 VSUBS 0.006288f
C944 B.n106 VSUBS 0.006288f
C945 B.n107 VSUBS 0.006288f
C946 B.n108 VSUBS 0.006288f
C947 B.n109 VSUBS 0.006288f
C948 B.n110 VSUBS 0.006288f
C949 B.n111 VSUBS 0.006288f
C950 B.n112 VSUBS 0.006288f
C951 B.n113 VSUBS 0.006288f
C952 B.n114 VSUBS 0.006288f
C953 B.n115 VSUBS 0.006288f
C954 B.n116 VSUBS 0.006288f
C955 B.n117 VSUBS 0.006288f
C956 B.n118 VSUBS 0.006288f
C957 B.n119 VSUBS 0.006288f
C958 B.n120 VSUBS 0.006288f
C959 B.n121 VSUBS 0.006288f
C960 B.n122 VSUBS 0.006288f
C961 B.n123 VSUBS 0.006288f
C962 B.n124 VSUBS 0.006288f
C963 B.n125 VSUBS 0.006288f
C964 B.n126 VSUBS 0.006288f
C965 B.n127 VSUBS 0.006288f
C966 B.n128 VSUBS 0.006288f
C967 B.n129 VSUBS 0.006288f
C968 B.n130 VSUBS 0.014967f
C969 B.n131 VSUBS 0.006288f
C970 B.n132 VSUBS 0.006288f
C971 B.n133 VSUBS 0.006288f
C972 B.n134 VSUBS 0.006288f
C973 B.n135 VSUBS 0.006288f
C974 B.n136 VSUBS 0.006288f
C975 B.n137 VSUBS 0.006288f
C976 B.n138 VSUBS 0.006288f
C977 B.n139 VSUBS 0.006288f
C978 B.n140 VSUBS 0.006288f
C979 B.n141 VSUBS 0.006288f
C980 B.n142 VSUBS 0.006288f
C981 B.n143 VSUBS 0.006288f
C982 B.n144 VSUBS 0.006288f
C983 B.n145 VSUBS 0.006288f
C984 B.n146 VSUBS 0.006288f
C985 B.n147 VSUBS 0.006288f
C986 B.n148 VSUBS 0.006288f
C987 B.n149 VSUBS 0.006288f
C988 B.n150 VSUBS 0.006288f
C989 B.n151 VSUBS 0.006288f
C990 B.n152 VSUBS 0.006288f
C991 B.n153 VSUBS 0.006288f
C992 B.n154 VSUBS 0.006288f
C993 B.n155 VSUBS 0.006288f
C994 B.n156 VSUBS 0.006288f
C995 B.n157 VSUBS 0.006288f
C996 B.t10 VSUBS 0.289164f
C997 B.t11 VSUBS 0.32757f
C998 B.t9 VSUBS 2.4098f
C999 B.n158 VSUBS 0.520102f
C1000 B.n159 VSUBS 0.28555f
C1001 B.n160 VSUBS 0.014568f
C1002 B.n161 VSUBS 0.006288f
C1003 B.n162 VSUBS 0.006288f
C1004 B.n163 VSUBS 0.006288f
C1005 B.n164 VSUBS 0.006288f
C1006 B.n165 VSUBS 0.006288f
C1007 B.t1 VSUBS 0.289161f
C1008 B.t2 VSUBS 0.327567f
C1009 B.t0 VSUBS 2.4098f
C1010 B.n166 VSUBS 0.520105f
C1011 B.n167 VSUBS 0.285553f
C1012 B.n168 VSUBS 0.006288f
C1013 B.n169 VSUBS 0.006288f
C1014 B.n170 VSUBS 0.006288f
C1015 B.n171 VSUBS 0.006288f
C1016 B.n172 VSUBS 0.006288f
C1017 B.n173 VSUBS 0.006288f
C1018 B.n174 VSUBS 0.006288f
C1019 B.n175 VSUBS 0.006288f
C1020 B.n176 VSUBS 0.006288f
C1021 B.n177 VSUBS 0.006288f
C1022 B.n178 VSUBS 0.006288f
C1023 B.n179 VSUBS 0.006288f
C1024 B.n180 VSUBS 0.006288f
C1025 B.n181 VSUBS 0.006288f
C1026 B.n182 VSUBS 0.006288f
C1027 B.n183 VSUBS 0.006288f
C1028 B.n184 VSUBS 0.006288f
C1029 B.n185 VSUBS 0.006288f
C1030 B.n186 VSUBS 0.006288f
C1031 B.n187 VSUBS 0.006288f
C1032 B.n188 VSUBS 0.006288f
C1033 B.n189 VSUBS 0.006288f
C1034 B.n190 VSUBS 0.006288f
C1035 B.n191 VSUBS 0.006288f
C1036 B.n192 VSUBS 0.006288f
C1037 B.n193 VSUBS 0.006288f
C1038 B.n194 VSUBS 0.006288f
C1039 B.n195 VSUBS 0.014253f
C1040 B.n196 VSUBS 0.006288f
C1041 B.n197 VSUBS 0.006288f
C1042 B.n198 VSUBS 0.006288f
C1043 B.n199 VSUBS 0.006288f
C1044 B.n200 VSUBS 0.006288f
C1045 B.n201 VSUBS 0.006288f
C1046 B.n202 VSUBS 0.006288f
C1047 B.n203 VSUBS 0.006288f
C1048 B.n204 VSUBS 0.006288f
C1049 B.n205 VSUBS 0.006288f
C1050 B.n206 VSUBS 0.006288f
C1051 B.n207 VSUBS 0.006288f
C1052 B.n208 VSUBS 0.006288f
C1053 B.n209 VSUBS 0.006288f
C1054 B.n210 VSUBS 0.006288f
C1055 B.n211 VSUBS 0.006288f
C1056 B.n212 VSUBS 0.006288f
C1057 B.n213 VSUBS 0.006288f
C1058 B.n214 VSUBS 0.006288f
C1059 B.n215 VSUBS 0.006288f
C1060 B.n216 VSUBS 0.006288f
C1061 B.n217 VSUBS 0.006288f
C1062 B.n218 VSUBS 0.006288f
C1063 B.n219 VSUBS 0.006288f
C1064 B.n220 VSUBS 0.006288f
C1065 B.n221 VSUBS 0.006288f
C1066 B.n222 VSUBS 0.006288f
C1067 B.n223 VSUBS 0.006288f
C1068 B.n224 VSUBS 0.006288f
C1069 B.n225 VSUBS 0.006288f
C1070 B.n226 VSUBS 0.006288f
C1071 B.n227 VSUBS 0.006288f
C1072 B.n228 VSUBS 0.006288f
C1073 B.n229 VSUBS 0.006288f
C1074 B.n230 VSUBS 0.006288f
C1075 B.n231 VSUBS 0.006288f
C1076 B.n232 VSUBS 0.006288f
C1077 B.n233 VSUBS 0.006288f
C1078 B.n234 VSUBS 0.006288f
C1079 B.n235 VSUBS 0.006288f
C1080 B.n236 VSUBS 0.006288f
C1081 B.n237 VSUBS 0.006288f
C1082 B.n238 VSUBS 0.006288f
C1083 B.n239 VSUBS 0.006288f
C1084 B.n240 VSUBS 0.006288f
C1085 B.n241 VSUBS 0.006288f
C1086 B.n242 VSUBS 0.006288f
C1087 B.n243 VSUBS 0.006288f
C1088 B.n244 VSUBS 0.006288f
C1089 B.n245 VSUBS 0.006288f
C1090 B.n246 VSUBS 0.006288f
C1091 B.n247 VSUBS 0.006288f
C1092 B.n248 VSUBS 0.006288f
C1093 B.n249 VSUBS 0.006288f
C1094 B.n250 VSUBS 0.006288f
C1095 B.n251 VSUBS 0.006288f
C1096 B.n252 VSUBS 0.006288f
C1097 B.n253 VSUBS 0.006288f
C1098 B.n254 VSUBS 0.006288f
C1099 B.n255 VSUBS 0.006288f
C1100 B.n256 VSUBS 0.006288f
C1101 B.n257 VSUBS 0.006288f
C1102 B.n258 VSUBS 0.006288f
C1103 B.n259 VSUBS 0.006288f
C1104 B.n260 VSUBS 0.006288f
C1105 B.n261 VSUBS 0.006288f
C1106 B.n262 VSUBS 0.006288f
C1107 B.n263 VSUBS 0.006288f
C1108 B.n264 VSUBS 0.006288f
C1109 B.n265 VSUBS 0.006288f
C1110 B.n266 VSUBS 0.006288f
C1111 B.n267 VSUBS 0.006288f
C1112 B.n268 VSUBS 0.006288f
C1113 B.n269 VSUBS 0.006288f
C1114 B.n270 VSUBS 0.006288f
C1115 B.n271 VSUBS 0.006288f
C1116 B.n272 VSUBS 0.006288f
C1117 B.n273 VSUBS 0.006288f
C1118 B.n274 VSUBS 0.006288f
C1119 B.n275 VSUBS 0.006288f
C1120 B.n276 VSUBS 0.014253f
C1121 B.n277 VSUBS 0.014967f
C1122 B.n278 VSUBS 0.014967f
C1123 B.n279 VSUBS 0.006288f
C1124 B.n280 VSUBS 0.006288f
C1125 B.n281 VSUBS 0.006288f
C1126 B.n282 VSUBS 0.006288f
C1127 B.n283 VSUBS 0.006288f
C1128 B.n284 VSUBS 0.006288f
C1129 B.n285 VSUBS 0.006288f
C1130 B.n286 VSUBS 0.006288f
C1131 B.n287 VSUBS 0.006288f
C1132 B.n288 VSUBS 0.006288f
C1133 B.n289 VSUBS 0.006288f
C1134 B.n290 VSUBS 0.006288f
C1135 B.n291 VSUBS 0.006288f
C1136 B.n292 VSUBS 0.006288f
C1137 B.n293 VSUBS 0.006288f
C1138 B.n294 VSUBS 0.006288f
C1139 B.n295 VSUBS 0.006288f
C1140 B.n296 VSUBS 0.006288f
C1141 B.n297 VSUBS 0.006288f
C1142 B.n298 VSUBS 0.006288f
C1143 B.n299 VSUBS 0.006288f
C1144 B.n300 VSUBS 0.006288f
C1145 B.n301 VSUBS 0.006288f
C1146 B.n302 VSUBS 0.006288f
C1147 B.n303 VSUBS 0.006288f
C1148 B.n304 VSUBS 0.006288f
C1149 B.n305 VSUBS 0.006288f
C1150 B.n306 VSUBS 0.006288f
C1151 B.n307 VSUBS 0.006288f
C1152 B.n308 VSUBS 0.006288f
C1153 B.n309 VSUBS 0.006288f
C1154 B.n310 VSUBS 0.006288f
C1155 B.n311 VSUBS 0.006288f
C1156 B.n312 VSUBS 0.006288f
C1157 B.n313 VSUBS 0.006288f
C1158 B.n314 VSUBS 0.006288f
C1159 B.n315 VSUBS 0.006288f
C1160 B.n316 VSUBS 0.006288f
C1161 B.n317 VSUBS 0.006288f
C1162 B.n318 VSUBS 0.006288f
C1163 B.n319 VSUBS 0.006288f
C1164 B.n320 VSUBS 0.006288f
C1165 B.n321 VSUBS 0.006288f
C1166 B.n322 VSUBS 0.006288f
C1167 B.n323 VSUBS 0.006288f
C1168 B.n324 VSUBS 0.006288f
C1169 B.n325 VSUBS 0.006288f
C1170 B.n326 VSUBS 0.006288f
C1171 B.n327 VSUBS 0.006288f
C1172 B.n328 VSUBS 0.006288f
C1173 B.n329 VSUBS 0.006288f
C1174 B.n330 VSUBS 0.006288f
C1175 B.n331 VSUBS 0.006288f
C1176 B.n332 VSUBS 0.006288f
C1177 B.n333 VSUBS 0.006288f
C1178 B.n334 VSUBS 0.006288f
C1179 B.n335 VSUBS 0.006288f
C1180 B.n336 VSUBS 0.006288f
C1181 B.n337 VSUBS 0.006288f
C1182 B.n338 VSUBS 0.006288f
C1183 B.n339 VSUBS 0.006288f
C1184 B.n340 VSUBS 0.006288f
C1185 B.n341 VSUBS 0.006288f
C1186 B.n342 VSUBS 0.006288f
C1187 B.n343 VSUBS 0.006288f
C1188 B.n344 VSUBS 0.006288f
C1189 B.n345 VSUBS 0.006288f
C1190 B.n346 VSUBS 0.006288f
C1191 B.n347 VSUBS 0.006288f
C1192 B.n348 VSUBS 0.006288f
C1193 B.n349 VSUBS 0.006288f
C1194 B.n350 VSUBS 0.006288f
C1195 B.n351 VSUBS 0.006288f
C1196 B.n352 VSUBS 0.006288f
C1197 B.n353 VSUBS 0.006288f
C1198 B.n354 VSUBS 0.006288f
C1199 B.n355 VSUBS 0.006288f
C1200 B.n356 VSUBS 0.006288f
C1201 B.n357 VSUBS 0.006288f
C1202 B.n358 VSUBS 0.006288f
C1203 B.n359 VSUBS 0.006288f
C1204 B.n360 VSUBS 0.004346f
C1205 B.n361 VSUBS 0.014568f
C1206 B.n362 VSUBS 0.005086f
C1207 B.n363 VSUBS 0.006288f
C1208 B.n364 VSUBS 0.006288f
C1209 B.n365 VSUBS 0.006288f
C1210 B.n366 VSUBS 0.006288f
C1211 B.n367 VSUBS 0.006288f
C1212 B.n368 VSUBS 0.006288f
C1213 B.n369 VSUBS 0.006288f
C1214 B.n370 VSUBS 0.006288f
C1215 B.n371 VSUBS 0.006288f
C1216 B.n372 VSUBS 0.006288f
C1217 B.n373 VSUBS 0.006288f
C1218 B.n374 VSUBS 0.005086f
C1219 B.n375 VSUBS 0.006288f
C1220 B.n376 VSUBS 0.006288f
C1221 B.n377 VSUBS 0.004346f
C1222 B.n378 VSUBS 0.006288f
C1223 B.n379 VSUBS 0.006288f
C1224 B.n380 VSUBS 0.006288f
C1225 B.n381 VSUBS 0.006288f
C1226 B.n382 VSUBS 0.006288f
C1227 B.n383 VSUBS 0.006288f
C1228 B.n384 VSUBS 0.006288f
C1229 B.n385 VSUBS 0.006288f
C1230 B.n386 VSUBS 0.006288f
C1231 B.n387 VSUBS 0.006288f
C1232 B.n388 VSUBS 0.006288f
C1233 B.n389 VSUBS 0.006288f
C1234 B.n390 VSUBS 0.006288f
C1235 B.n391 VSUBS 0.006288f
C1236 B.n392 VSUBS 0.006288f
C1237 B.n393 VSUBS 0.006288f
C1238 B.n394 VSUBS 0.006288f
C1239 B.n395 VSUBS 0.006288f
C1240 B.n396 VSUBS 0.006288f
C1241 B.n397 VSUBS 0.006288f
C1242 B.n398 VSUBS 0.006288f
C1243 B.n399 VSUBS 0.006288f
C1244 B.n400 VSUBS 0.006288f
C1245 B.n401 VSUBS 0.006288f
C1246 B.n402 VSUBS 0.006288f
C1247 B.n403 VSUBS 0.006288f
C1248 B.n404 VSUBS 0.006288f
C1249 B.n405 VSUBS 0.006288f
C1250 B.n406 VSUBS 0.006288f
C1251 B.n407 VSUBS 0.006288f
C1252 B.n408 VSUBS 0.006288f
C1253 B.n409 VSUBS 0.006288f
C1254 B.n410 VSUBS 0.006288f
C1255 B.n411 VSUBS 0.006288f
C1256 B.n412 VSUBS 0.006288f
C1257 B.n413 VSUBS 0.006288f
C1258 B.n414 VSUBS 0.006288f
C1259 B.n415 VSUBS 0.006288f
C1260 B.n416 VSUBS 0.006288f
C1261 B.n417 VSUBS 0.006288f
C1262 B.n418 VSUBS 0.006288f
C1263 B.n419 VSUBS 0.006288f
C1264 B.n420 VSUBS 0.006288f
C1265 B.n421 VSUBS 0.006288f
C1266 B.n422 VSUBS 0.006288f
C1267 B.n423 VSUBS 0.006288f
C1268 B.n424 VSUBS 0.006288f
C1269 B.n425 VSUBS 0.006288f
C1270 B.n426 VSUBS 0.006288f
C1271 B.n427 VSUBS 0.006288f
C1272 B.n428 VSUBS 0.006288f
C1273 B.n429 VSUBS 0.006288f
C1274 B.n430 VSUBS 0.006288f
C1275 B.n431 VSUBS 0.006288f
C1276 B.n432 VSUBS 0.006288f
C1277 B.n433 VSUBS 0.006288f
C1278 B.n434 VSUBS 0.006288f
C1279 B.n435 VSUBS 0.006288f
C1280 B.n436 VSUBS 0.006288f
C1281 B.n437 VSUBS 0.006288f
C1282 B.n438 VSUBS 0.006288f
C1283 B.n439 VSUBS 0.006288f
C1284 B.n440 VSUBS 0.006288f
C1285 B.n441 VSUBS 0.006288f
C1286 B.n442 VSUBS 0.006288f
C1287 B.n443 VSUBS 0.006288f
C1288 B.n444 VSUBS 0.006288f
C1289 B.n445 VSUBS 0.006288f
C1290 B.n446 VSUBS 0.006288f
C1291 B.n447 VSUBS 0.006288f
C1292 B.n448 VSUBS 0.006288f
C1293 B.n449 VSUBS 0.006288f
C1294 B.n450 VSUBS 0.006288f
C1295 B.n451 VSUBS 0.006288f
C1296 B.n452 VSUBS 0.006288f
C1297 B.n453 VSUBS 0.006288f
C1298 B.n454 VSUBS 0.006288f
C1299 B.n455 VSUBS 0.006288f
C1300 B.n456 VSUBS 0.006288f
C1301 B.n457 VSUBS 0.006288f
C1302 B.n458 VSUBS 0.006288f
C1303 B.n459 VSUBS 0.014967f
C1304 B.n460 VSUBS 0.014253f
C1305 B.n461 VSUBS 0.014253f
C1306 B.n462 VSUBS 0.006288f
C1307 B.n463 VSUBS 0.006288f
C1308 B.n464 VSUBS 0.006288f
C1309 B.n465 VSUBS 0.006288f
C1310 B.n466 VSUBS 0.006288f
C1311 B.n467 VSUBS 0.006288f
C1312 B.n468 VSUBS 0.006288f
C1313 B.n469 VSUBS 0.006288f
C1314 B.n470 VSUBS 0.006288f
C1315 B.n471 VSUBS 0.006288f
C1316 B.n472 VSUBS 0.006288f
C1317 B.n473 VSUBS 0.006288f
C1318 B.n474 VSUBS 0.006288f
C1319 B.n475 VSUBS 0.006288f
C1320 B.n476 VSUBS 0.006288f
C1321 B.n477 VSUBS 0.006288f
C1322 B.n478 VSUBS 0.006288f
C1323 B.n479 VSUBS 0.006288f
C1324 B.n480 VSUBS 0.006288f
C1325 B.n481 VSUBS 0.006288f
C1326 B.n482 VSUBS 0.006288f
C1327 B.n483 VSUBS 0.006288f
C1328 B.n484 VSUBS 0.006288f
C1329 B.n485 VSUBS 0.006288f
C1330 B.n486 VSUBS 0.006288f
C1331 B.n487 VSUBS 0.006288f
C1332 B.n488 VSUBS 0.006288f
C1333 B.n489 VSUBS 0.006288f
C1334 B.n490 VSUBS 0.006288f
C1335 B.n491 VSUBS 0.006288f
C1336 B.n492 VSUBS 0.006288f
C1337 B.n493 VSUBS 0.006288f
C1338 B.n494 VSUBS 0.006288f
C1339 B.n495 VSUBS 0.006288f
C1340 B.n496 VSUBS 0.006288f
C1341 B.n497 VSUBS 0.006288f
C1342 B.n498 VSUBS 0.006288f
C1343 B.n499 VSUBS 0.006288f
C1344 B.n500 VSUBS 0.006288f
C1345 B.n501 VSUBS 0.006288f
C1346 B.n502 VSUBS 0.006288f
C1347 B.n503 VSUBS 0.006288f
C1348 B.n504 VSUBS 0.006288f
C1349 B.n505 VSUBS 0.006288f
C1350 B.n506 VSUBS 0.006288f
C1351 B.n507 VSUBS 0.006288f
C1352 B.n508 VSUBS 0.006288f
C1353 B.n509 VSUBS 0.006288f
C1354 B.n510 VSUBS 0.006288f
C1355 B.n511 VSUBS 0.006288f
C1356 B.n512 VSUBS 0.006288f
C1357 B.n513 VSUBS 0.006288f
C1358 B.n514 VSUBS 0.006288f
C1359 B.n515 VSUBS 0.006288f
C1360 B.n516 VSUBS 0.006288f
C1361 B.n517 VSUBS 0.006288f
C1362 B.n518 VSUBS 0.006288f
C1363 B.n519 VSUBS 0.006288f
C1364 B.n520 VSUBS 0.006288f
C1365 B.n521 VSUBS 0.006288f
C1366 B.n522 VSUBS 0.006288f
C1367 B.n523 VSUBS 0.006288f
C1368 B.n524 VSUBS 0.006288f
C1369 B.n525 VSUBS 0.006288f
C1370 B.n526 VSUBS 0.006288f
C1371 B.n527 VSUBS 0.006288f
C1372 B.n528 VSUBS 0.006288f
C1373 B.n529 VSUBS 0.006288f
C1374 B.n530 VSUBS 0.006288f
C1375 B.n531 VSUBS 0.006288f
C1376 B.n532 VSUBS 0.006288f
C1377 B.n533 VSUBS 0.006288f
C1378 B.n534 VSUBS 0.006288f
C1379 B.n535 VSUBS 0.006288f
C1380 B.n536 VSUBS 0.006288f
C1381 B.n537 VSUBS 0.006288f
C1382 B.n538 VSUBS 0.006288f
C1383 B.n539 VSUBS 0.006288f
C1384 B.n540 VSUBS 0.006288f
C1385 B.n541 VSUBS 0.006288f
C1386 B.n542 VSUBS 0.006288f
C1387 B.n543 VSUBS 0.006288f
C1388 B.n544 VSUBS 0.006288f
C1389 B.n545 VSUBS 0.006288f
C1390 B.n546 VSUBS 0.006288f
C1391 B.n547 VSUBS 0.006288f
C1392 B.n548 VSUBS 0.006288f
C1393 B.n549 VSUBS 0.006288f
C1394 B.n550 VSUBS 0.006288f
C1395 B.n551 VSUBS 0.006288f
C1396 B.n552 VSUBS 0.006288f
C1397 B.n553 VSUBS 0.006288f
C1398 B.n554 VSUBS 0.006288f
C1399 B.n555 VSUBS 0.006288f
C1400 B.n556 VSUBS 0.006288f
C1401 B.n557 VSUBS 0.006288f
C1402 B.n558 VSUBS 0.006288f
C1403 B.n559 VSUBS 0.006288f
C1404 B.n560 VSUBS 0.006288f
C1405 B.n561 VSUBS 0.006288f
C1406 B.n562 VSUBS 0.006288f
C1407 B.n563 VSUBS 0.006288f
C1408 B.n564 VSUBS 0.006288f
C1409 B.n565 VSUBS 0.006288f
C1410 B.n566 VSUBS 0.006288f
C1411 B.n567 VSUBS 0.006288f
C1412 B.n568 VSUBS 0.006288f
C1413 B.n569 VSUBS 0.006288f
C1414 B.n570 VSUBS 0.006288f
C1415 B.n571 VSUBS 0.006288f
C1416 B.n572 VSUBS 0.006288f
C1417 B.n573 VSUBS 0.006288f
C1418 B.n574 VSUBS 0.006288f
C1419 B.n575 VSUBS 0.006288f
C1420 B.n576 VSUBS 0.006288f
C1421 B.n577 VSUBS 0.006288f
C1422 B.n578 VSUBS 0.006288f
C1423 B.n579 VSUBS 0.006288f
C1424 B.n580 VSUBS 0.006288f
C1425 B.n581 VSUBS 0.006288f
C1426 B.n582 VSUBS 0.006288f
C1427 B.n583 VSUBS 0.006288f
C1428 B.n584 VSUBS 0.006288f
C1429 B.n585 VSUBS 0.006288f
C1430 B.n586 VSUBS 0.014253f
C1431 B.n587 VSUBS 0.015004f
C1432 B.n588 VSUBS 0.014216f
C1433 B.n589 VSUBS 0.006288f
C1434 B.n590 VSUBS 0.006288f
C1435 B.n591 VSUBS 0.006288f
C1436 B.n592 VSUBS 0.006288f
C1437 B.n593 VSUBS 0.006288f
C1438 B.n594 VSUBS 0.006288f
C1439 B.n595 VSUBS 0.006288f
C1440 B.n596 VSUBS 0.006288f
C1441 B.n597 VSUBS 0.006288f
C1442 B.n598 VSUBS 0.006288f
C1443 B.n599 VSUBS 0.006288f
C1444 B.n600 VSUBS 0.006288f
C1445 B.n601 VSUBS 0.006288f
C1446 B.n602 VSUBS 0.006288f
C1447 B.n603 VSUBS 0.006288f
C1448 B.n604 VSUBS 0.006288f
C1449 B.n605 VSUBS 0.006288f
C1450 B.n606 VSUBS 0.006288f
C1451 B.n607 VSUBS 0.006288f
C1452 B.n608 VSUBS 0.006288f
C1453 B.n609 VSUBS 0.006288f
C1454 B.n610 VSUBS 0.006288f
C1455 B.n611 VSUBS 0.006288f
C1456 B.n612 VSUBS 0.006288f
C1457 B.n613 VSUBS 0.006288f
C1458 B.n614 VSUBS 0.006288f
C1459 B.n615 VSUBS 0.006288f
C1460 B.n616 VSUBS 0.006288f
C1461 B.n617 VSUBS 0.006288f
C1462 B.n618 VSUBS 0.006288f
C1463 B.n619 VSUBS 0.006288f
C1464 B.n620 VSUBS 0.006288f
C1465 B.n621 VSUBS 0.006288f
C1466 B.n622 VSUBS 0.006288f
C1467 B.n623 VSUBS 0.006288f
C1468 B.n624 VSUBS 0.006288f
C1469 B.n625 VSUBS 0.006288f
C1470 B.n626 VSUBS 0.006288f
C1471 B.n627 VSUBS 0.006288f
C1472 B.n628 VSUBS 0.006288f
C1473 B.n629 VSUBS 0.006288f
C1474 B.n630 VSUBS 0.006288f
C1475 B.n631 VSUBS 0.006288f
C1476 B.n632 VSUBS 0.006288f
C1477 B.n633 VSUBS 0.006288f
C1478 B.n634 VSUBS 0.006288f
C1479 B.n635 VSUBS 0.006288f
C1480 B.n636 VSUBS 0.006288f
C1481 B.n637 VSUBS 0.006288f
C1482 B.n638 VSUBS 0.006288f
C1483 B.n639 VSUBS 0.006288f
C1484 B.n640 VSUBS 0.006288f
C1485 B.n641 VSUBS 0.006288f
C1486 B.n642 VSUBS 0.006288f
C1487 B.n643 VSUBS 0.006288f
C1488 B.n644 VSUBS 0.006288f
C1489 B.n645 VSUBS 0.006288f
C1490 B.n646 VSUBS 0.006288f
C1491 B.n647 VSUBS 0.006288f
C1492 B.n648 VSUBS 0.006288f
C1493 B.n649 VSUBS 0.006288f
C1494 B.n650 VSUBS 0.006288f
C1495 B.n651 VSUBS 0.006288f
C1496 B.n652 VSUBS 0.006288f
C1497 B.n653 VSUBS 0.006288f
C1498 B.n654 VSUBS 0.006288f
C1499 B.n655 VSUBS 0.006288f
C1500 B.n656 VSUBS 0.006288f
C1501 B.n657 VSUBS 0.006288f
C1502 B.n658 VSUBS 0.006288f
C1503 B.n659 VSUBS 0.006288f
C1504 B.n660 VSUBS 0.006288f
C1505 B.n661 VSUBS 0.006288f
C1506 B.n662 VSUBS 0.006288f
C1507 B.n663 VSUBS 0.006288f
C1508 B.n664 VSUBS 0.006288f
C1509 B.n665 VSUBS 0.006288f
C1510 B.n666 VSUBS 0.006288f
C1511 B.n667 VSUBS 0.006288f
C1512 B.n668 VSUBS 0.006288f
C1513 B.n669 VSUBS 0.006288f
C1514 B.n670 VSUBS 0.006288f
C1515 B.n671 VSUBS 0.004346f
C1516 B.n672 VSUBS 0.014568f
C1517 B.n673 VSUBS 0.005086f
C1518 B.n674 VSUBS 0.006288f
C1519 B.n675 VSUBS 0.006288f
C1520 B.n676 VSUBS 0.006288f
C1521 B.n677 VSUBS 0.006288f
C1522 B.n678 VSUBS 0.006288f
C1523 B.n679 VSUBS 0.006288f
C1524 B.n680 VSUBS 0.006288f
C1525 B.n681 VSUBS 0.006288f
C1526 B.n682 VSUBS 0.006288f
C1527 B.n683 VSUBS 0.006288f
C1528 B.n684 VSUBS 0.006288f
C1529 B.n685 VSUBS 0.005086f
C1530 B.n686 VSUBS 0.014568f
C1531 B.n687 VSUBS 0.004346f
C1532 B.n688 VSUBS 0.006288f
C1533 B.n689 VSUBS 0.006288f
C1534 B.n690 VSUBS 0.006288f
C1535 B.n691 VSUBS 0.006288f
C1536 B.n692 VSUBS 0.006288f
C1537 B.n693 VSUBS 0.006288f
C1538 B.n694 VSUBS 0.006288f
C1539 B.n695 VSUBS 0.006288f
C1540 B.n696 VSUBS 0.006288f
C1541 B.n697 VSUBS 0.006288f
C1542 B.n698 VSUBS 0.006288f
C1543 B.n699 VSUBS 0.006288f
C1544 B.n700 VSUBS 0.006288f
C1545 B.n701 VSUBS 0.006288f
C1546 B.n702 VSUBS 0.006288f
C1547 B.n703 VSUBS 0.006288f
C1548 B.n704 VSUBS 0.006288f
C1549 B.n705 VSUBS 0.006288f
C1550 B.n706 VSUBS 0.006288f
C1551 B.n707 VSUBS 0.006288f
C1552 B.n708 VSUBS 0.006288f
C1553 B.n709 VSUBS 0.006288f
C1554 B.n710 VSUBS 0.006288f
C1555 B.n711 VSUBS 0.006288f
C1556 B.n712 VSUBS 0.006288f
C1557 B.n713 VSUBS 0.006288f
C1558 B.n714 VSUBS 0.006288f
C1559 B.n715 VSUBS 0.006288f
C1560 B.n716 VSUBS 0.006288f
C1561 B.n717 VSUBS 0.006288f
C1562 B.n718 VSUBS 0.006288f
C1563 B.n719 VSUBS 0.006288f
C1564 B.n720 VSUBS 0.006288f
C1565 B.n721 VSUBS 0.006288f
C1566 B.n722 VSUBS 0.006288f
C1567 B.n723 VSUBS 0.006288f
C1568 B.n724 VSUBS 0.006288f
C1569 B.n725 VSUBS 0.006288f
C1570 B.n726 VSUBS 0.006288f
C1571 B.n727 VSUBS 0.006288f
C1572 B.n728 VSUBS 0.006288f
C1573 B.n729 VSUBS 0.006288f
C1574 B.n730 VSUBS 0.006288f
C1575 B.n731 VSUBS 0.006288f
C1576 B.n732 VSUBS 0.006288f
C1577 B.n733 VSUBS 0.006288f
C1578 B.n734 VSUBS 0.006288f
C1579 B.n735 VSUBS 0.006288f
C1580 B.n736 VSUBS 0.006288f
C1581 B.n737 VSUBS 0.006288f
C1582 B.n738 VSUBS 0.006288f
C1583 B.n739 VSUBS 0.006288f
C1584 B.n740 VSUBS 0.006288f
C1585 B.n741 VSUBS 0.006288f
C1586 B.n742 VSUBS 0.006288f
C1587 B.n743 VSUBS 0.006288f
C1588 B.n744 VSUBS 0.006288f
C1589 B.n745 VSUBS 0.006288f
C1590 B.n746 VSUBS 0.006288f
C1591 B.n747 VSUBS 0.006288f
C1592 B.n748 VSUBS 0.006288f
C1593 B.n749 VSUBS 0.006288f
C1594 B.n750 VSUBS 0.006288f
C1595 B.n751 VSUBS 0.006288f
C1596 B.n752 VSUBS 0.006288f
C1597 B.n753 VSUBS 0.006288f
C1598 B.n754 VSUBS 0.006288f
C1599 B.n755 VSUBS 0.006288f
C1600 B.n756 VSUBS 0.006288f
C1601 B.n757 VSUBS 0.006288f
C1602 B.n758 VSUBS 0.006288f
C1603 B.n759 VSUBS 0.006288f
C1604 B.n760 VSUBS 0.006288f
C1605 B.n761 VSUBS 0.006288f
C1606 B.n762 VSUBS 0.006288f
C1607 B.n763 VSUBS 0.006288f
C1608 B.n764 VSUBS 0.006288f
C1609 B.n765 VSUBS 0.006288f
C1610 B.n766 VSUBS 0.006288f
C1611 B.n767 VSUBS 0.006288f
C1612 B.n768 VSUBS 0.006288f
C1613 B.n769 VSUBS 0.006288f
C1614 B.n770 VSUBS 0.014967f
C1615 B.n771 VSUBS 0.014253f
C1616 B.n772 VSUBS 0.014253f
C1617 B.n773 VSUBS 0.006288f
C1618 B.n774 VSUBS 0.006288f
C1619 B.n775 VSUBS 0.006288f
C1620 B.n776 VSUBS 0.006288f
C1621 B.n777 VSUBS 0.006288f
C1622 B.n778 VSUBS 0.006288f
C1623 B.n779 VSUBS 0.006288f
C1624 B.n780 VSUBS 0.006288f
C1625 B.n781 VSUBS 0.006288f
C1626 B.n782 VSUBS 0.006288f
C1627 B.n783 VSUBS 0.006288f
C1628 B.n784 VSUBS 0.006288f
C1629 B.n785 VSUBS 0.006288f
C1630 B.n786 VSUBS 0.006288f
C1631 B.n787 VSUBS 0.006288f
C1632 B.n788 VSUBS 0.006288f
C1633 B.n789 VSUBS 0.006288f
C1634 B.n790 VSUBS 0.006288f
C1635 B.n791 VSUBS 0.006288f
C1636 B.n792 VSUBS 0.006288f
C1637 B.n793 VSUBS 0.006288f
C1638 B.n794 VSUBS 0.006288f
C1639 B.n795 VSUBS 0.006288f
C1640 B.n796 VSUBS 0.006288f
C1641 B.n797 VSUBS 0.006288f
C1642 B.n798 VSUBS 0.006288f
C1643 B.n799 VSUBS 0.006288f
C1644 B.n800 VSUBS 0.006288f
C1645 B.n801 VSUBS 0.006288f
C1646 B.n802 VSUBS 0.006288f
C1647 B.n803 VSUBS 0.006288f
C1648 B.n804 VSUBS 0.006288f
C1649 B.n805 VSUBS 0.006288f
C1650 B.n806 VSUBS 0.006288f
C1651 B.n807 VSUBS 0.006288f
C1652 B.n808 VSUBS 0.006288f
C1653 B.n809 VSUBS 0.006288f
C1654 B.n810 VSUBS 0.006288f
C1655 B.n811 VSUBS 0.006288f
C1656 B.n812 VSUBS 0.006288f
C1657 B.n813 VSUBS 0.006288f
C1658 B.n814 VSUBS 0.006288f
C1659 B.n815 VSUBS 0.006288f
C1660 B.n816 VSUBS 0.006288f
C1661 B.n817 VSUBS 0.006288f
C1662 B.n818 VSUBS 0.006288f
C1663 B.n819 VSUBS 0.006288f
C1664 B.n820 VSUBS 0.006288f
C1665 B.n821 VSUBS 0.006288f
C1666 B.n822 VSUBS 0.006288f
C1667 B.n823 VSUBS 0.006288f
C1668 B.n824 VSUBS 0.006288f
C1669 B.n825 VSUBS 0.006288f
C1670 B.n826 VSUBS 0.006288f
C1671 B.n827 VSUBS 0.006288f
C1672 B.n828 VSUBS 0.006288f
C1673 B.n829 VSUBS 0.006288f
C1674 B.n830 VSUBS 0.006288f
C1675 B.n831 VSUBS 0.006288f
C1676 B.n832 VSUBS 0.006288f
C1677 B.n833 VSUBS 0.006288f
C1678 B.n834 VSUBS 0.006288f
C1679 B.n835 VSUBS 0.014238f
.ends

