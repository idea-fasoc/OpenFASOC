* NGSPICE file created from diff_pair_sample_0226.ext - technology: sky130A

.subckt diff_pair_sample_0226 VTAIL VN VP B VDD2 VDD1
X0 B.t15 B.t13 B.t14 B.t7 sky130_fd_pr__nfet_01v8 ad=1.2714 pd=7.3 as=0 ps=0 w=3.26 l=3.41
X1 VDD1.t1 VP.t0 VTAIL.t2 B.t0 sky130_fd_pr__nfet_01v8 ad=1.2714 pd=7.3 as=1.2714 ps=7.3 w=3.26 l=3.41
X2 VDD1.t0 VP.t1 VTAIL.t3 B.t1 sky130_fd_pr__nfet_01v8 ad=1.2714 pd=7.3 as=1.2714 ps=7.3 w=3.26 l=3.41
X3 B.t12 B.t10 B.t11 B.t3 sky130_fd_pr__nfet_01v8 ad=1.2714 pd=7.3 as=0 ps=0 w=3.26 l=3.41
X4 VDD2.t1 VN.t0 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=1.2714 pd=7.3 as=1.2714 ps=7.3 w=3.26 l=3.41
X5 B.t9 B.t6 B.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=1.2714 pd=7.3 as=0 ps=0 w=3.26 l=3.41
X6 B.t5 B.t2 B.t4 B.t3 sky130_fd_pr__nfet_01v8 ad=1.2714 pd=7.3 as=0 ps=0 w=3.26 l=3.41
X7 VDD2.t0 VN.t1 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=1.2714 pd=7.3 as=1.2714 ps=7.3 w=3.26 l=3.41
R0 B.n377 B.n82 585
R1 B.n82 B.n57 585
R2 B.n379 B.n378 585
R3 B.n381 B.n81 585
R4 B.n384 B.n383 585
R5 B.n385 B.n80 585
R6 B.n387 B.n386 585
R7 B.n389 B.n79 585
R8 B.n392 B.n391 585
R9 B.n393 B.n78 585
R10 B.n395 B.n394 585
R11 B.n397 B.n77 585
R12 B.n400 B.n399 585
R13 B.n401 B.n76 585
R14 B.n403 B.n402 585
R15 B.n405 B.n75 585
R16 B.n408 B.n407 585
R17 B.n410 B.n72 585
R18 B.n412 B.n411 585
R19 B.n414 B.n71 585
R20 B.n417 B.n416 585
R21 B.n418 B.n70 585
R22 B.n420 B.n419 585
R23 B.n422 B.n69 585
R24 B.n425 B.n424 585
R25 B.n426 B.n66 585
R26 B.n429 B.n428 585
R27 B.n431 B.n65 585
R28 B.n434 B.n433 585
R29 B.n435 B.n64 585
R30 B.n437 B.n436 585
R31 B.n439 B.n63 585
R32 B.n442 B.n441 585
R33 B.n443 B.n62 585
R34 B.n445 B.n444 585
R35 B.n447 B.n61 585
R36 B.n450 B.n449 585
R37 B.n451 B.n60 585
R38 B.n453 B.n452 585
R39 B.n455 B.n59 585
R40 B.n458 B.n457 585
R41 B.n459 B.n58 585
R42 B.n376 B.n56 585
R43 B.n462 B.n56 585
R44 B.n375 B.n55 585
R45 B.n463 B.n55 585
R46 B.n374 B.n54 585
R47 B.n464 B.n54 585
R48 B.n373 B.n372 585
R49 B.n372 B.n50 585
R50 B.n371 B.n49 585
R51 B.n470 B.n49 585
R52 B.n370 B.n48 585
R53 B.n471 B.n48 585
R54 B.n369 B.n47 585
R55 B.n472 B.n47 585
R56 B.n368 B.n367 585
R57 B.n367 B.n43 585
R58 B.n366 B.n42 585
R59 B.n478 B.n42 585
R60 B.n365 B.n41 585
R61 B.n479 B.n41 585
R62 B.n364 B.n40 585
R63 B.n480 B.n40 585
R64 B.n363 B.n362 585
R65 B.n362 B.n36 585
R66 B.n361 B.n35 585
R67 B.n486 B.n35 585
R68 B.n360 B.n34 585
R69 B.n487 B.n34 585
R70 B.n359 B.n33 585
R71 B.n488 B.n33 585
R72 B.n358 B.n357 585
R73 B.n357 B.n29 585
R74 B.n356 B.n28 585
R75 B.n494 B.n28 585
R76 B.n355 B.n27 585
R77 B.n495 B.n27 585
R78 B.n354 B.n26 585
R79 B.n496 B.n26 585
R80 B.n353 B.n352 585
R81 B.n352 B.n22 585
R82 B.n351 B.n21 585
R83 B.n502 B.n21 585
R84 B.n350 B.n20 585
R85 B.n503 B.n20 585
R86 B.n349 B.n19 585
R87 B.n504 B.n19 585
R88 B.n348 B.n347 585
R89 B.n347 B.n15 585
R90 B.n346 B.n14 585
R91 B.n510 B.n14 585
R92 B.n345 B.n13 585
R93 B.n511 B.n13 585
R94 B.n344 B.n12 585
R95 B.n512 B.n12 585
R96 B.n343 B.n342 585
R97 B.n342 B.n8 585
R98 B.n341 B.n7 585
R99 B.n518 B.n7 585
R100 B.n340 B.n6 585
R101 B.n519 B.n6 585
R102 B.n339 B.n5 585
R103 B.n520 B.n5 585
R104 B.n338 B.n337 585
R105 B.n337 B.n4 585
R106 B.n336 B.n83 585
R107 B.n336 B.n335 585
R108 B.n326 B.n84 585
R109 B.n85 B.n84 585
R110 B.n328 B.n327 585
R111 B.n329 B.n328 585
R112 B.n325 B.n90 585
R113 B.n90 B.n89 585
R114 B.n324 B.n323 585
R115 B.n323 B.n322 585
R116 B.n92 B.n91 585
R117 B.n93 B.n92 585
R118 B.n315 B.n314 585
R119 B.n316 B.n315 585
R120 B.n313 B.n98 585
R121 B.n98 B.n97 585
R122 B.n312 B.n311 585
R123 B.n311 B.n310 585
R124 B.n100 B.n99 585
R125 B.n101 B.n100 585
R126 B.n303 B.n302 585
R127 B.n304 B.n303 585
R128 B.n301 B.n106 585
R129 B.n106 B.n105 585
R130 B.n300 B.n299 585
R131 B.n299 B.n298 585
R132 B.n108 B.n107 585
R133 B.n109 B.n108 585
R134 B.n291 B.n290 585
R135 B.n292 B.n291 585
R136 B.n289 B.n114 585
R137 B.n114 B.n113 585
R138 B.n288 B.n287 585
R139 B.n287 B.n286 585
R140 B.n116 B.n115 585
R141 B.n117 B.n116 585
R142 B.n279 B.n278 585
R143 B.n280 B.n279 585
R144 B.n277 B.n122 585
R145 B.n122 B.n121 585
R146 B.n276 B.n275 585
R147 B.n275 B.n274 585
R148 B.n124 B.n123 585
R149 B.n125 B.n124 585
R150 B.n267 B.n266 585
R151 B.n268 B.n267 585
R152 B.n265 B.n130 585
R153 B.n130 B.n129 585
R154 B.n264 B.n263 585
R155 B.n263 B.n262 585
R156 B.n132 B.n131 585
R157 B.n133 B.n132 585
R158 B.n255 B.n254 585
R159 B.n256 B.n255 585
R160 B.n253 B.n138 585
R161 B.n138 B.n137 585
R162 B.n252 B.n251 585
R163 B.n251 B.n250 585
R164 B.n247 B.n142 585
R165 B.n246 B.n245 585
R166 B.n243 B.n143 585
R167 B.n243 B.n141 585
R168 B.n242 B.n241 585
R169 B.n240 B.n239 585
R170 B.n238 B.n145 585
R171 B.n236 B.n235 585
R172 B.n234 B.n146 585
R173 B.n233 B.n232 585
R174 B.n230 B.n147 585
R175 B.n228 B.n227 585
R176 B.n226 B.n148 585
R177 B.n225 B.n224 585
R178 B.n222 B.n149 585
R179 B.n220 B.n219 585
R180 B.n218 B.n150 585
R181 B.n216 B.n215 585
R182 B.n213 B.n153 585
R183 B.n211 B.n210 585
R184 B.n209 B.n154 585
R185 B.n208 B.n207 585
R186 B.n205 B.n155 585
R187 B.n203 B.n202 585
R188 B.n201 B.n156 585
R189 B.n200 B.n199 585
R190 B.n197 B.n196 585
R191 B.n195 B.n194 585
R192 B.n193 B.n161 585
R193 B.n191 B.n190 585
R194 B.n189 B.n162 585
R195 B.n188 B.n187 585
R196 B.n185 B.n163 585
R197 B.n183 B.n182 585
R198 B.n181 B.n164 585
R199 B.n180 B.n179 585
R200 B.n177 B.n165 585
R201 B.n175 B.n174 585
R202 B.n173 B.n166 585
R203 B.n172 B.n171 585
R204 B.n169 B.n167 585
R205 B.n140 B.n139 585
R206 B.n249 B.n248 585
R207 B.n250 B.n249 585
R208 B.n136 B.n135 585
R209 B.n137 B.n136 585
R210 B.n258 B.n257 585
R211 B.n257 B.n256 585
R212 B.n259 B.n134 585
R213 B.n134 B.n133 585
R214 B.n261 B.n260 585
R215 B.n262 B.n261 585
R216 B.n128 B.n127 585
R217 B.n129 B.n128 585
R218 B.n270 B.n269 585
R219 B.n269 B.n268 585
R220 B.n271 B.n126 585
R221 B.n126 B.n125 585
R222 B.n273 B.n272 585
R223 B.n274 B.n273 585
R224 B.n120 B.n119 585
R225 B.n121 B.n120 585
R226 B.n282 B.n281 585
R227 B.n281 B.n280 585
R228 B.n283 B.n118 585
R229 B.n118 B.n117 585
R230 B.n285 B.n284 585
R231 B.n286 B.n285 585
R232 B.n112 B.n111 585
R233 B.n113 B.n112 585
R234 B.n294 B.n293 585
R235 B.n293 B.n292 585
R236 B.n295 B.n110 585
R237 B.n110 B.n109 585
R238 B.n297 B.n296 585
R239 B.n298 B.n297 585
R240 B.n104 B.n103 585
R241 B.n105 B.n104 585
R242 B.n306 B.n305 585
R243 B.n305 B.n304 585
R244 B.n307 B.n102 585
R245 B.n102 B.n101 585
R246 B.n309 B.n308 585
R247 B.n310 B.n309 585
R248 B.n96 B.n95 585
R249 B.n97 B.n96 585
R250 B.n318 B.n317 585
R251 B.n317 B.n316 585
R252 B.n319 B.n94 585
R253 B.n94 B.n93 585
R254 B.n321 B.n320 585
R255 B.n322 B.n321 585
R256 B.n88 B.n87 585
R257 B.n89 B.n88 585
R258 B.n331 B.n330 585
R259 B.n330 B.n329 585
R260 B.n332 B.n86 585
R261 B.n86 B.n85 585
R262 B.n334 B.n333 585
R263 B.n335 B.n334 585
R264 B.n2 B.n0 585
R265 B.n4 B.n2 585
R266 B.n3 B.n1 585
R267 B.n519 B.n3 585
R268 B.n517 B.n516 585
R269 B.n518 B.n517 585
R270 B.n515 B.n9 585
R271 B.n9 B.n8 585
R272 B.n514 B.n513 585
R273 B.n513 B.n512 585
R274 B.n11 B.n10 585
R275 B.n511 B.n11 585
R276 B.n509 B.n508 585
R277 B.n510 B.n509 585
R278 B.n507 B.n16 585
R279 B.n16 B.n15 585
R280 B.n506 B.n505 585
R281 B.n505 B.n504 585
R282 B.n18 B.n17 585
R283 B.n503 B.n18 585
R284 B.n501 B.n500 585
R285 B.n502 B.n501 585
R286 B.n499 B.n23 585
R287 B.n23 B.n22 585
R288 B.n498 B.n497 585
R289 B.n497 B.n496 585
R290 B.n25 B.n24 585
R291 B.n495 B.n25 585
R292 B.n493 B.n492 585
R293 B.n494 B.n493 585
R294 B.n491 B.n30 585
R295 B.n30 B.n29 585
R296 B.n490 B.n489 585
R297 B.n489 B.n488 585
R298 B.n32 B.n31 585
R299 B.n487 B.n32 585
R300 B.n485 B.n484 585
R301 B.n486 B.n485 585
R302 B.n483 B.n37 585
R303 B.n37 B.n36 585
R304 B.n482 B.n481 585
R305 B.n481 B.n480 585
R306 B.n39 B.n38 585
R307 B.n479 B.n39 585
R308 B.n477 B.n476 585
R309 B.n478 B.n477 585
R310 B.n475 B.n44 585
R311 B.n44 B.n43 585
R312 B.n474 B.n473 585
R313 B.n473 B.n472 585
R314 B.n46 B.n45 585
R315 B.n471 B.n46 585
R316 B.n469 B.n468 585
R317 B.n470 B.n469 585
R318 B.n467 B.n51 585
R319 B.n51 B.n50 585
R320 B.n466 B.n465 585
R321 B.n465 B.n464 585
R322 B.n53 B.n52 585
R323 B.n463 B.n53 585
R324 B.n461 B.n460 585
R325 B.n462 B.n461 585
R326 B.n522 B.n521 585
R327 B.n521 B.n520 585
R328 B.n249 B.n142 550.159
R329 B.n461 B.n58 550.159
R330 B.n251 B.n140 550.159
R331 B.n82 B.n56 550.159
R332 B.n380 B.n57 256.663
R333 B.n382 B.n57 256.663
R334 B.n388 B.n57 256.663
R335 B.n390 B.n57 256.663
R336 B.n396 B.n57 256.663
R337 B.n398 B.n57 256.663
R338 B.n404 B.n57 256.663
R339 B.n406 B.n57 256.663
R340 B.n413 B.n57 256.663
R341 B.n415 B.n57 256.663
R342 B.n421 B.n57 256.663
R343 B.n423 B.n57 256.663
R344 B.n430 B.n57 256.663
R345 B.n432 B.n57 256.663
R346 B.n438 B.n57 256.663
R347 B.n440 B.n57 256.663
R348 B.n446 B.n57 256.663
R349 B.n448 B.n57 256.663
R350 B.n454 B.n57 256.663
R351 B.n456 B.n57 256.663
R352 B.n244 B.n141 256.663
R353 B.n144 B.n141 256.663
R354 B.n237 B.n141 256.663
R355 B.n231 B.n141 256.663
R356 B.n229 B.n141 256.663
R357 B.n223 B.n141 256.663
R358 B.n221 B.n141 256.663
R359 B.n214 B.n141 256.663
R360 B.n212 B.n141 256.663
R361 B.n206 B.n141 256.663
R362 B.n204 B.n141 256.663
R363 B.n198 B.n141 256.663
R364 B.n160 B.n141 256.663
R365 B.n192 B.n141 256.663
R366 B.n186 B.n141 256.663
R367 B.n184 B.n141 256.663
R368 B.n178 B.n141 256.663
R369 B.n176 B.n141 256.663
R370 B.n170 B.n141 256.663
R371 B.n168 B.n141 256.663
R372 B.n157 B.t10 232.052
R373 B.n151 B.t2 232.052
R374 B.n67 B.t13 232.052
R375 B.n73 B.t6 232.052
R376 B.n157 B.t12 205.876
R377 B.n73 B.t8 205.876
R378 B.n151 B.t5 205.876
R379 B.n67 B.t14 205.876
R380 B.n250 B.n141 168.834
R381 B.n462 B.n57 168.834
R382 B.n249 B.n136 163.367
R383 B.n257 B.n136 163.367
R384 B.n257 B.n134 163.367
R385 B.n261 B.n134 163.367
R386 B.n261 B.n128 163.367
R387 B.n269 B.n128 163.367
R388 B.n269 B.n126 163.367
R389 B.n273 B.n126 163.367
R390 B.n273 B.n120 163.367
R391 B.n281 B.n120 163.367
R392 B.n281 B.n118 163.367
R393 B.n285 B.n118 163.367
R394 B.n285 B.n112 163.367
R395 B.n293 B.n112 163.367
R396 B.n293 B.n110 163.367
R397 B.n297 B.n110 163.367
R398 B.n297 B.n104 163.367
R399 B.n305 B.n104 163.367
R400 B.n305 B.n102 163.367
R401 B.n309 B.n102 163.367
R402 B.n309 B.n96 163.367
R403 B.n317 B.n96 163.367
R404 B.n317 B.n94 163.367
R405 B.n321 B.n94 163.367
R406 B.n321 B.n88 163.367
R407 B.n330 B.n88 163.367
R408 B.n330 B.n86 163.367
R409 B.n334 B.n86 163.367
R410 B.n334 B.n2 163.367
R411 B.n521 B.n2 163.367
R412 B.n521 B.n3 163.367
R413 B.n517 B.n3 163.367
R414 B.n517 B.n9 163.367
R415 B.n513 B.n9 163.367
R416 B.n513 B.n11 163.367
R417 B.n509 B.n11 163.367
R418 B.n509 B.n16 163.367
R419 B.n505 B.n16 163.367
R420 B.n505 B.n18 163.367
R421 B.n501 B.n18 163.367
R422 B.n501 B.n23 163.367
R423 B.n497 B.n23 163.367
R424 B.n497 B.n25 163.367
R425 B.n493 B.n25 163.367
R426 B.n493 B.n30 163.367
R427 B.n489 B.n30 163.367
R428 B.n489 B.n32 163.367
R429 B.n485 B.n32 163.367
R430 B.n485 B.n37 163.367
R431 B.n481 B.n37 163.367
R432 B.n481 B.n39 163.367
R433 B.n477 B.n39 163.367
R434 B.n477 B.n44 163.367
R435 B.n473 B.n44 163.367
R436 B.n473 B.n46 163.367
R437 B.n469 B.n46 163.367
R438 B.n469 B.n51 163.367
R439 B.n465 B.n51 163.367
R440 B.n465 B.n53 163.367
R441 B.n461 B.n53 163.367
R442 B.n245 B.n243 163.367
R443 B.n243 B.n242 163.367
R444 B.n239 B.n238 163.367
R445 B.n236 B.n146 163.367
R446 B.n232 B.n230 163.367
R447 B.n228 B.n148 163.367
R448 B.n224 B.n222 163.367
R449 B.n220 B.n150 163.367
R450 B.n215 B.n213 163.367
R451 B.n211 B.n154 163.367
R452 B.n207 B.n205 163.367
R453 B.n203 B.n156 163.367
R454 B.n199 B.n197 163.367
R455 B.n194 B.n193 163.367
R456 B.n191 B.n162 163.367
R457 B.n187 B.n185 163.367
R458 B.n183 B.n164 163.367
R459 B.n179 B.n177 163.367
R460 B.n175 B.n166 163.367
R461 B.n171 B.n169 163.367
R462 B.n251 B.n138 163.367
R463 B.n255 B.n138 163.367
R464 B.n255 B.n132 163.367
R465 B.n263 B.n132 163.367
R466 B.n263 B.n130 163.367
R467 B.n267 B.n130 163.367
R468 B.n267 B.n124 163.367
R469 B.n275 B.n124 163.367
R470 B.n275 B.n122 163.367
R471 B.n279 B.n122 163.367
R472 B.n279 B.n116 163.367
R473 B.n287 B.n116 163.367
R474 B.n287 B.n114 163.367
R475 B.n291 B.n114 163.367
R476 B.n291 B.n108 163.367
R477 B.n299 B.n108 163.367
R478 B.n299 B.n106 163.367
R479 B.n303 B.n106 163.367
R480 B.n303 B.n100 163.367
R481 B.n311 B.n100 163.367
R482 B.n311 B.n98 163.367
R483 B.n315 B.n98 163.367
R484 B.n315 B.n92 163.367
R485 B.n323 B.n92 163.367
R486 B.n323 B.n90 163.367
R487 B.n328 B.n90 163.367
R488 B.n328 B.n84 163.367
R489 B.n336 B.n84 163.367
R490 B.n337 B.n336 163.367
R491 B.n337 B.n5 163.367
R492 B.n6 B.n5 163.367
R493 B.n7 B.n6 163.367
R494 B.n342 B.n7 163.367
R495 B.n342 B.n12 163.367
R496 B.n13 B.n12 163.367
R497 B.n14 B.n13 163.367
R498 B.n347 B.n14 163.367
R499 B.n347 B.n19 163.367
R500 B.n20 B.n19 163.367
R501 B.n21 B.n20 163.367
R502 B.n352 B.n21 163.367
R503 B.n352 B.n26 163.367
R504 B.n27 B.n26 163.367
R505 B.n28 B.n27 163.367
R506 B.n357 B.n28 163.367
R507 B.n357 B.n33 163.367
R508 B.n34 B.n33 163.367
R509 B.n35 B.n34 163.367
R510 B.n362 B.n35 163.367
R511 B.n362 B.n40 163.367
R512 B.n41 B.n40 163.367
R513 B.n42 B.n41 163.367
R514 B.n367 B.n42 163.367
R515 B.n367 B.n47 163.367
R516 B.n48 B.n47 163.367
R517 B.n49 B.n48 163.367
R518 B.n372 B.n49 163.367
R519 B.n372 B.n54 163.367
R520 B.n55 B.n54 163.367
R521 B.n56 B.n55 163.367
R522 B.n457 B.n455 163.367
R523 B.n453 B.n60 163.367
R524 B.n449 B.n447 163.367
R525 B.n445 B.n62 163.367
R526 B.n441 B.n439 163.367
R527 B.n437 B.n64 163.367
R528 B.n433 B.n431 163.367
R529 B.n429 B.n66 163.367
R530 B.n424 B.n422 163.367
R531 B.n420 B.n70 163.367
R532 B.n416 B.n414 163.367
R533 B.n412 B.n72 163.367
R534 B.n407 B.n405 163.367
R535 B.n403 B.n76 163.367
R536 B.n399 B.n397 163.367
R537 B.n395 B.n78 163.367
R538 B.n391 B.n389 163.367
R539 B.n387 B.n80 163.367
R540 B.n383 B.n381 163.367
R541 B.n379 B.n82 163.367
R542 B.n158 B.t11 133.343
R543 B.n74 B.t9 133.343
R544 B.n152 B.t4 133.343
R545 B.n68 B.t15 133.343
R546 B.n250 B.n137 87.6396
R547 B.n256 B.n137 87.6396
R548 B.n256 B.n133 87.6396
R549 B.n262 B.n133 87.6396
R550 B.n262 B.n129 87.6396
R551 B.n268 B.n129 87.6396
R552 B.n268 B.n125 87.6396
R553 B.n274 B.n125 87.6396
R554 B.n280 B.n121 87.6396
R555 B.n280 B.n117 87.6396
R556 B.n286 B.n117 87.6396
R557 B.n286 B.n113 87.6396
R558 B.n292 B.n113 87.6396
R559 B.n292 B.n109 87.6396
R560 B.n298 B.n109 87.6396
R561 B.n298 B.n105 87.6396
R562 B.n304 B.n105 87.6396
R563 B.n304 B.n101 87.6396
R564 B.n310 B.n101 87.6396
R565 B.n310 B.n97 87.6396
R566 B.n316 B.n97 87.6396
R567 B.n322 B.n93 87.6396
R568 B.n322 B.n89 87.6396
R569 B.n329 B.n89 87.6396
R570 B.n329 B.n85 87.6396
R571 B.n335 B.n85 87.6396
R572 B.n335 B.n4 87.6396
R573 B.n520 B.n4 87.6396
R574 B.n520 B.n519 87.6396
R575 B.n519 B.n518 87.6396
R576 B.n518 B.n8 87.6396
R577 B.n512 B.n8 87.6396
R578 B.n512 B.n511 87.6396
R579 B.n511 B.n510 87.6396
R580 B.n510 B.n15 87.6396
R581 B.n504 B.n503 87.6396
R582 B.n503 B.n502 87.6396
R583 B.n502 B.n22 87.6396
R584 B.n496 B.n22 87.6396
R585 B.n496 B.n495 87.6396
R586 B.n495 B.n494 87.6396
R587 B.n494 B.n29 87.6396
R588 B.n488 B.n29 87.6396
R589 B.n488 B.n487 87.6396
R590 B.n487 B.n486 87.6396
R591 B.n486 B.n36 87.6396
R592 B.n480 B.n36 87.6396
R593 B.n480 B.n479 87.6396
R594 B.n478 B.n43 87.6396
R595 B.n472 B.n43 87.6396
R596 B.n472 B.n471 87.6396
R597 B.n471 B.n470 87.6396
R598 B.n470 B.n50 87.6396
R599 B.n464 B.n50 87.6396
R600 B.n464 B.n463 87.6396
R601 B.n463 B.n462 87.6396
R602 B.n316 B.t0 78.618
R603 B.n504 B.t1 78.618
R604 B.n158 B.n157 72.5338
R605 B.n152 B.n151 72.5338
R606 B.n68 B.n67 72.5338
R607 B.n74 B.n73 72.5338
R608 B.n244 B.n142 71.676
R609 B.n242 B.n144 71.676
R610 B.n238 B.n237 71.676
R611 B.n231 B.n146 71.676
R612 B.n230 B.n229 71.676
R613 B.n223 B.n148 71.676
R614 B.n222 B.n221 71.676
R615 B.n214 B.n150 71.676
R616 B.n213 B.n212 71.676
R617 B.n206 B.n154 71.676
R618 B.n205 B.n204 71.676
R619 B.n198 B.n156 71.676
R620 B.n197 B.n160 71.676
R621 B.n193 B.n192 71.676
R622 B.n186 B.n162 71.676
R623 B.n185 B.n184 71.676
R624 B.n178 B.n164 71.676
R625 B.n177 B.n176 71.676
R626 B.n170 B.n166 71.676
R627 B.n169 B.n168 71.676
R628 B.n456 B.n58 71.676
R629 B.n455 B.n454 71.676
R630 B.n448 B.n60 71.676
R631 B.n447 B.n446 71.676
R632 B.n440 B.n62 71.676
R633 B.n439 B.n438 71.676
R634 B.n432 B.n64 71.676
R635 B.n431 B.n430 71.676
R636 B.n423 B.n66 71.676
R637 B.n422 B.n421 71.676
R638 B.n415 B.n70 71.676
R639 B.n414 B.n413 71.676
R640 B.n406 B.n72 71.676
R641 B.n405 B.n404 71.676
R642 B.n398 B.n76 71.676
R643 B.n397 B.n396 71.676
R644 B.n390 B.n78 71.676
R645 B.n389 B.n388 71.676
R646 B.n382 B.n80 71.676
R647 B.n381 B.n380 71.676
R648 B.n380 B.n379 71.676
R649 B.n383 B.n382 71.676
R650 B.n388 B.n387 71.676
R651 B.n391 B.n390 71.676
R652 B.n396 B.n395 71.676
R653 B.n399 B.n398 71.676
R654 B.n404 B.n403 71.676
R655 B.n407 B.n406 71.676
R656 B.n413 B.n412 71.676
R657 B.n416 B.n415 71.676
R658 B.n421 B.n420 71.676
R659 B.n424 B.n423 71.676
R660 B.n430 B.n429 71.676
R661 B.n433 B.n432 71.676
R662 B.n438 B.n437 71.676
R663 B.n441 B.n440 71.676
R664 B.n446 B.n445 71.676
R665 B.n449 B.n448 71.676
R666 B.n454 B.n453 71.676
R667 B.n457 B.n456 71.676
R668 B.n245 B.n244 71.676
R669 B.n239 B.n144 71.676
R670 B.n237 B.n236 71.676
R671 B.n232 B.n231 71.676
R672 B.n229 B.n228 71.676
R673 B.n224 B.n223 71.676
R674 B.n221 B.n220 71.676
R675 B.n215 B.n214 71.676
R676 B.n212 B.n211 71.676
R677 B.n207 B.n206 71.676
R678 B.n204 B.n203 71.676
R679 B.n199 B.n198 71.676
R680 B.n194 B.n160 71.676
R681 B.n192 B.n191 71.676
R682 B.n187 B.n186 71.676
R683 B.n184 B.n183 71.676
R684 B.n179 B.n178 71.676
R685 B.n176 B.n175 71.676
R686 B.n171 B.n170 71.676
R687 B.n168 B.n140 71.676
R688 B.n274 B.t3 60.5746
R689 B.t7 B.n478 60.5746
R690 B.n159 B.n158 59.5399
R691 B.n217 B.n152 59.5399
R692 B.n427 B.n68 59.5399
R693 B.n409 B.n74 59.5399
R694 B.n460 B.n459 35.7468
R695 B.n252 B.n139 35.7468
R696 B.n248 B.n247 35.7468
R697 B.n377 B.n376 35.7468
R698 B.t3 B.n121 27.0655
R699 B.n479 B.t7 27.0655
R700 B B.n522 18.0485
R701 B.n459 B.n458 10.6151
R702 B.n458 B.n59 10.6151
R703 B.n452 B.n59 10.6151
R704 B.n452 B.n451 10.6151
R705 B.n451 B.n450 10.6151
R706 B.n450 B.n61 10.6151
R707 B.n444 B.n61 10.6151
R708 B.n444 B.n443 10.6151
R709 B.n443 B.n442 10.6151
R710 B.n442 B.n63 10.6151
R711 B.n436 B.n63 10.6151
R712 B.n436 B.n435 10.6151
R713 B.n435 B.n434 10.6151
R714 B.n434 B.n65 10.6151
R715 B.n428 B.n65 10.6151
R716 B.n426 B.n425 10.6151
R717 B.n425 B.n69 10.6151
R718 B.n419 B.n69 10.6151
R719 B.n419 B.n418 10.6151
R720 B.n418 B.n417 10.6151
R721 B.n417 B.n71 10.6151
R722 B.n411 B.n71 10.6151
R723 B.n411 B.n410 10.6151
R724 B.n408 B.n75 10.6151
R725 B.n402 B.n75 10.6151
R726 B.n402 B.n401 10.6151
R727 B.n401 B.n400 10.6151
R728 B.n400 B.n77 10.6151
R729 B.n394 B.n77 10.6151
R730 B.n394 B.n393 10.6151
R731 B.n393 B.n392 10.6151
R732 B.n392 B.n79 10.6151
R733 B.n386 B.n79 10.6151
R734 B.n386 B.n385 10.6151
R735 B.n385 B.n384 10.6151
R736 B.n384 B.n81 10.6151
R737 B.n378 B.n81 10.6151
R738 B.n378 B.n377 10.6151
R739 B.n253 B.n252 10.6151
R740 B.n254 B.n253 10.6151
R741 B.n254 B.n131 10.6151
R742 B.n264 B.n131 10.6151
R743 B.n265 B.n264 10.6151
R744 B.n266 B.n265 10.6151
R745 B.n266 B.n123 10.6151
R746 B.n276 B.n123 10.6151
R747 B.n277 B.n276 10.6151
R748 B.n278 B.n277 10.6151
R749 B.n278 B.n115 10.6151
R750 B.n288 B.n115 10.6151
R751 B.n289 B.n288 10.6151
R752 B.n290 B.n289 10.6151
R753 B.n290 B.n107 10.6151
R754 B.n300 B.n107 10.6151
R755 B.n301 B.n300 10.6151
R756 B.n302 B.n301 10.6151
R757 B.n302 B.n99 10.6151
R758 B.n312 B.n99 10.6151
R759 B.n313 B.n312 10.6151
R760 B.n314 B.n313 10.6151
R761 B.n314 B.n91 10.6151
R762 B.n324 B.n91 10.6151
R763 B.n325 B.n324 10.6151
R764 B.n327 B.n325 10.6151
R765 B.n327 B.n326 10.6151
R766 B.n326 B.n83 10.6151
R767 B.n338 B.n83 10.6151
R768 B.n339 B.n338 10.6151
R769 B.n340 B.n339 10.6151
R770 B.n341 B.n340 10.6151
R771 B.n343 B.n341 10.6151
R772 B.n344 B.n343 10.6151
R773 B.n345 B.n344 10.6151
R774 B.n346 B.n345 10.6151
R775 B.n348 B.n346 10.6151
R776 B.n349 B.n348 10.6151
R777 B.n350 B.n349 10.6151
R778 B.n351 B.n350 10.6151
R779 B.n353 B.n351 10.6151
R780 B.n354 B.n353 10.6151
R781 B.n355 B.n354 10.6151
R782 B.n356 B.n355 10.6151
R783 B.n358 B.n356 10.6151
R784 B.n359 B.n358 10.6151
R785 B.n360 B.n359 10.6151
R786 B.n361 B.n360 10.6151
R787 B.n363 B.n361 10.6151
R788 B.n364 B.n363 10.6151
R789 B.n365 B.n364 10.6151
R790 B.n366 B.n365 10.6151
R791 B.n368 B.n366 10.6151
R792 B.n369 B.n368 10.6151
R793 B.n370 B.n369 10.6151
R794 B.n371 B.n370 10.6151
R795 B.n373 B.n371 10.6151
R796 B.n374 B.n373 10.6151
R797 B.n375 B.n374 10.6151
R798 B.n376 B.n375 10.6151
R799 B.n247 B.n246 10.6151
R800 B.n246 B.n143 10.6151
R801 B.n241 B.n143 10.6151
R802 B.n241 B.n240 10.6151
R803 B.n240 B.n145 10.6151
R804 B.n235 B.n145 10.6151
R805 B.n235 B.n234 10.6151
R806 B.n234 B.n233 10.6151
R807 B.n233 B.n147 10.6151
R808 B.n227 B.n147 10.6151
R809 B.n227 B.n226 10.6151
R810 B.n226 B.n225 10.6151
R811 B.n225 B.n149 10.6151
R812 B.n219 B.n149 10.6151
R813 B.n219 B.n218 10.6151
R814 B.n216 B.n153 10.6151
R815 B.n210 B.n153 10.6151
R816 B.n210 B.n209 10.6151
R817 B.n209 B.n208 10.6151
R818 B.n208 B.n155 10.6151
R819 B.n202 B.n155 10.6151
R820 B.n202 B.n201 10.6151
R821 B.n201 B.n200 10.6151
R822 B.n196 B.n195 10.6151
R823 B.n195 B.n161 10.6151
R824 B.n190 B.n161 10.6151
R825 B.n190 B.n189 10.6151
R826 B.n189 B.n188 10.6151
R827 B.n188 B.n163 10.6151
R828 B.n182 B.n163 10.6151
R829 B.n182 B.n181 10.6151
R830 B.n181 B.n180 10.6151
R831 B.n180 B.n165 10.6151
R832 B.n174 B.n165 10.6151
R833 B.n174 B.n173 10.6151
R834 B.n173 B.n172 10.6151
R835 B.n172 B.n167 10.6151
R836 B.n167 B.n139 10.6151
R837 B.n248 B.n135 10.6151
R838 B.n258 B.n135 10.6151
R839 B.n259 B.n258 10.6151
R840 B.n260 B.n259 10.6151
R841 B.n260 B.n127 10.6151
R842 B.n270 B.n127 10.6151
R843 B.n271 B.n270 10.6151
R844 B.n272 B.n271 10.6151
R845 B.n272 B.n119 10.6151
R846 B.n282 B.n119 10.6151
R847 B.n283 B.n282 10.6151
R848 B.n284 B.n283 10.6151
R849 B.n284 B.n111 10.6151
R850 B.n294 B.n111 10.6151
R851 B.n295 B.n294 10.6151
R852 B.n296 B.n295 10.6151
R853 B.n296 B.n103 10.6151
R854 B.n306 B.n103 10.6151
R855 B.n307 B.n306 10.6151
R856 B.n308 B.n307 10.6151
R857 B.n308 B.n95 10.6151
R858 B.n318 B.n95 10.6151
R859 B.n319 B.n318 10.6151
R860 B.n320 B.n319 10.6151
R861 B.n320 B.n87 10.6151
R862 B.n331 B.n87 10.6151
R863 B.n332 B.n331 10.6151
R864 B.n333 B.n332 10.6151
R865 B.n333 B.n0 10.6151
R866 B.n516 B.n1 10.6151
R867 B.n516 B.n515 10.6151
R868 B.n515 B.n514 10.6151
R869 B.n514 B.n10 10.6151
R870 B.n508 B.n10 10.6151
R871 B.n508 B.n507 10.6151
R872 B.n507 B.n506 10.6151
R873 B.n506 B.n17 10.6151
R874 B.n500 B.n17 10.6151
R875 B.n500 B.n499 10.6151
R876 B.n499 B.n498 10.6151
R877 B.n498 B.n24 10.6151
R878 B.n492 B.n24 10.6151
R879 B.n492 B.n491 10.6151
R880 B.n491 B.n490 10.6151
R881 B.n490 B.n31 10.6151
R882 B.n484 B.n31 10.6151
R883 B.n484 B.n483 10.6151
R884 B.n483 B.n482 10.6151
R885 B.n482 B.n38 10.6151
R886 B.n476 B.n38 10.6151
R887 B.n476 B.n475 10.6151
R888 B.n475 B.n474 10.6151
R889 B.n474 B.n45 10.6151
R890 B.n468 B.n45 10.6151
R891 B.n468 B.n467 10.6151
R892 B.n467 B.n466 10.6151
R893 B.n466 B.n52 10.6151
R894 B.n460 B.n52 10.6151
R895 B.t0 B.n93 9.02218
R896 B.t1 B.n15 9.02218
R897 B.n427 B.n426 6.5566
R898 B.n410 B.n409 6.5566
R899 B.n217 B.n216 6.5566
R900 B.n200 B.n159 6.5566
R901 B.n428 B.n427 4.05904
R902 B.n409 B.n408 4.05904
R903 B.n218 B.n217 4.05904
R904 B.n196 B.n159 4.05904
R905 B.n522 B.n0 2.81026
R906 B.n522 B.n1 2.81026
R907 VP.n0 VP.t1 102.07
R908 VP.n0 VP.t0 61.8861
R909 VP VP.n0 0.526373
R910 VTAIL.n58 VTAIL.n48 289.615
R911 VTAIL.n10 VTAIL.n0 289.615
R912 VTAIL.n42 VTAIL.n32 289.615
R913 VTAIL.n26 VTAIL.n16 289.615
R914 VTAIL.n52 VTAIL.n51 185
R915 VTAIL.n57 VTAIL.n56 185
R916 VTAIL.n59 VTAIL.n58 185
R917 VTAIL.n4 VTAIL.n3 185
R918 VTAIL.n9 VTAIL.n8 185
R919 VTAIL.n11 VTAIL.n10 185
R920 VTAIL.n43 VTAIL.n42 185
R921 VTAIL.n41 VTAIL.n40 185
R922 VTAIL.n36 VTAIL.n35 185
R923 VTAIL.n27 VTAIL.n26 185
R924 VTAIL.n25 VTAIL.n24 185
R925 VTAIL.n20 VTAIL.n19 185
R926 VTAIL.n53 VTAIL.t1 148.606
R927 VTAIL.n5 VTAIL.t2 148.606
R928 VTAIL.n37 VTAIL.t3 148.606
R929 VTAIL.n21 VTAIL.t0 148.606
R930 VTAIL.n57 VTAIL.n51 104.615
R931 VTAIL.n58 VTAIL.n57 104.615
R932 VTAIL.n9 VTAIL.n3 104.615
R933 VTAIL.n10 VTAIL.n9 104.615
R934 VTAIL.n42 VTAIL.n41 104.615
R935 VTAIL.n41 VTAIL.n35 104.615
R936 VTAIL.n26 VTAIL.n25 104.615
R937 VTAIL.n25 VTAIL.n19 104.615
R938 VTAIL.t1 VTAIL.n51 52.3082
R939 VTAIL.t2 VTAIL.n3 52.3082
R940 VTAIL.t3 VTAIL.n35 52.3082
R941 VTAIL.t0 VTAIL.n19 52.3082
R942 VTAIL.n63 VTAIL.n62 34.9005
R943 VTAIL.n15 VTAIL.n14 34.9005
R944 VTAIL.n47 VTAIL.n46 34.9005
R945 VTAIL.n31 VTAIL.n30 34.9005
R946 VTAIL.n31 VTAIL.n15 21.6255
R947 VTAIL.n63 VTAIL.n47 18.4014
R948 VTAIL.n53 VTAIL.n52 15.5966
R949 VTAIL.n5 VTAIL.n4 15.5966
R950 VTAIL.n37 VTAIL.n36 15.5966
R951 VTAIL.n21 VTAIL.n20 15.5966
R952 VTAIL.n56 VTAIL.n55 12.8005
R953 VTAIL.n8 VTAIL.n7 12.8005
R954 VTAIL.n40 VTAIL.n39 12.8005
R955 VTAIL.n24 VTAIL.n23 12.8005
R956 VTAIL.n59 VTAIL.n50 12.0247
R957 VTAIL.n11 VTAIL.n2 12.0247
R958 VTAIL.n43 VTAIL.n34 12.0247
R959 VTAIL.n27 VTAIL.n18 12.0247
R960 VTAIL.n60 VTAIL.n48 11.249
R961 VTAIL.n12 VTAIL.n0 11.249
R962 VTAIL.n44 VTAIL.n32 11.249
R963 VTAIL.n28 VTAIL.n16 11.249
R964 VTAIL.n62 VTAIL.n61 9.45567
R965 VTAIL.n14 VTAIL.n13 9.45567
R966 VTAIL.n46 VTAIL.n45 9.45567
R967 VTAIL.n30 VTAIL.n29 9.45567
R968 VTAIL.n61 VTAIL.n60 9.3005
R969 VTAIL.n50 VTAIL.n49 9.3005
R970 VTAIL.n55 VTAIL.n54 9.3005
R971 VTAIL.n13 VTAIL.n12 9.3005
R972 VTAIL.n2 VTAIL.n1 9.3005
R973 VTAIL.n7 VTAIL.n6 9.3005
R974 VTAIL.n45 VTAIL.n44 9.3005
R975 VTAIL.n34 VTAIL.n33 9.3005
R976 VTAIL.n39 VTAIL.n38 9.3005
R977 VTAIL.n29 VTAIL.n28 9.3005
R978 VTAIL.n18 VTAIL.n17 9.3005
R979 VTAIL.n23 VTAIL.n22 9.3005
R980 VTAIL.n54 VTAIL.n53 4.46457
R981 VTAIL.n6 VTAIL.n5 4.46457
R982 VTAIL.n38 VTAIL.n37 4.46457
R983 VTAIL.n22 VTAIL.n21 4.46457
R984 VTAIL.n62 VTAIL.n48 2.71565
R985 VTAIL.n14 VTAIL.n0 2.71565
R986 VTAIL.n46 VTAIL.n32 2.71565
R987 VTAIL.n30 VTAIL.n16 2.71565
R988 VTAIL.n47 VTAIL.n31 2.0824
R989 VTAIL.n60 VTAIL.n59 1.93989
R990 VTAIL.n12 VTAIL.n11 1.93989
R991 VTAIL.n44 VTAIL.n43 1.93989
R992 VTAIL.n28 VTAIL.n27 1.93989
R993 VTAIL VTAIL.n15 1.33455
R994 VTAIL.n56 VTAIL.n50 1.16414
R995 VTAIL.n8 VTAIL.n2 1.16414
R996 VTAIL.n40 VTAIL.n34 1.16414
R997 VTAIL.n24 VTAIL.n18 1.16414
R998 VTAIL VTAIL.n63 0.748345
R999 VTAIL.n55 VTAIL.n52 0.388379
R1000 VTAIL.n7 VTAIL.n4 0.388379
R1001 VTAIL.n39 VTAIL.n36 0.388379
R1002 VTAIL.n23 VTAIL.n20 0.388379
R1003 VTAIL.n54 VTAIL.n49 0.155672
R1004 VTAIL.n61 VTAIL.n49 0.155672
R1005 VTAIL.n6 VTAIL.n1 0.155672
R1006 VTAIL.n13 VTAIL.n1 0.155672
R1007 VTAIL.n45 VTAIL.n33 0.155672
R1008 VTAIL.n38 VTAIL.n33 0.155672
R1009 VTAIL.n29 VTAIL.n17 0.155672
R1010 VTAIL.n22 VTAIL.n17 0.155672
R1011 VDD1.n10 VDD1.n0 289.615
R1012 VDD1.n25 VDD1.n15 289.615
R1013 VDD1.n11 VDD1.n10 185
R1014 VDD1.n9 VDD1.n8 185
R1015 VDD1.n4 VDD1.n3 185
R1016 VDD1.n19 VDD1.n18 185
R1017 VDD1.n24 VDD1.n23 185
R1018 VDD1.n26 VDD1.n25 185
R1019 VDD1.n5 VDD1.t0 148.606
R1020 VDD1.n20 VDD1.t1 148.606
R1021 VDD1.n10 VDD1.n9 104.615
R1022 VDD1.n9 VDD1.n3 104.615
R1023 VDD1.n24 VDD1.n18 104.615
R1024 VDD1.n25 VDD1.n24 104.615
R1025 VDD1 VDD1.n29 85.8282
R1026 VDD1 VDD1.n14 52.4435
R1027 VDD1.t0 VDD1.n3 52.3082
R1028 VDD1.t1 VDD1.n18 52.3082
R1029 VDD1.n5 VDD1.n4 15.5966
R1030 VDD1.n20 VDD1.n19 15.5966
R1031 VDD1.n8 VDD1.n7 12.8005
R1032 VDD1.n23 VDD1.n22 12.8005
R1033 VDD1.n11 VDD1.n2 12.0247
R1034 VDD1.n26 VDD1.n17 12.0247
R1035 VDD1.n12 VDD1.n0 11.249
R1036 VDD1.n27 VDD1.n15 11.249
R1037 VDD1.n14 VDD1.n13 9.45567
R1038 VDD1.n29 VDD1.n28 9.45567
R1039 VDD1.n13 VDD1.n12 9.3005
R1040 VDD1.n2 VDD1.n1 9.3005
R1041 VDD1.n7 VDD1.n6 9.3005
R1042 VDD1.n28 VDD1.n27 9.3005
R1043 VDD1.n17 VDD1.n16 9.3005
R1044 VDD1.n22 VDD1.n21 9.3005
R1045 VDD1.n6 VDD1.n5 4.46457
R1046 VDD1.n21 VDD1.n20 4.46457
R1047 VDD1.n14 VDD1.n0 2.71565
R1048 VDD1.n29 VDD1.n15 2.71565
R1049 VDD1.n12 VDD1.n11 1.93989
R1050 VDD1.n27 VDD1.n26 1.93989
R1051 VDD1.n8 VDD1.n2 1.16414
R1052 VDD1.n23 VDD1.n17 1.16414
R1053 VDD1.n7 VDD1.n4 0.388379
R1054 VDD1.n22 VDD1.n19 0.388379
R1055 VDD1.n13 VDD1.n1 0.155672
R1056 VDD1.n6 VDD1.n1 0.155672
R1057 VDD1.n21 VDD1.n16 0.155672
R1058 VDD1.n28 VDD1.n16 0.155672
R1059 VN VN.t0 101.977
R1060 VN VN.t1 62.4119
R1061 VDD2.n25 VDD2.n15 289.615
R1062 VDD2.n10 VDD2.n0 289.615
R1063 VDD2.n26 VDD2.n25 185
R1064 VDD2.n24 VDD2.n23 185
R1065 VDD2.n19 VDD2.n18 185
R1066 VDD2.n4 VDD2.n3 185
R1067 VDD2.n9 VDD2.n8 185
R1068 VDD2.n11 VDD2.n10 185
R1069 VDD2.n20 VDD2.t1 148.606
R1070 VDD2.n5 VDD2.t0 148.606
R1071 VDD2.n25 VDD2.n24 104.615
R1072 VDD2.n24 VDD2.n18 104.615
R1073 VDD2.n9 VDD2.n3 104.615
R1074 VDD2.n10 VDD2.n9 104.615
R1075 VDD2.n30 VDD2.n14 84.4973
R1076 VDD2.t1 VDD2.n18 52.3082
R1077 VDD2.t0 VDD2.n3 52.3082
R1078 VDD2.n30 VDD2.n29 51.5793
R1079 VDD2.n20 VDD2.n19 15.5966
R1080 VDD2.n5 VDD2.n4 15.5966
R1081 VDD2.n23 VDD2.n22 12.8005
R1082 VDD2.n8 VDD2.n7 12.8005
R1083 VDD2.n26 VDD2.n17 12.0247
R1084 VDD2.n11 VDD2.n2 12.0247
R1085 VDD2.n27 VDD2.n15 11.249
R1086 VDD2.n12 VDD2.n0 11.249
R1087 VDD2.n29 VDD2.n28 9.45567
R1088 VDD2.n14 VDD2.n13 9.45567
R1089 VDD2.n28 VDD2.n27 9.3005
R1090 VDD2.n17 VDD2.n16 9.3005
R1091 VDD2.n22 VDD2.n21 9.3005
R1092 VDD2.n13 VDD2.n12 9.3005
R1093 VDD2.n2 VDD2.n1 9.3005
R1094 VDD2.n7 VDD2.n6 9.3005
R1095 VDD2.n21 VDD2.n20 4.46457
R1096 VDD2.n6 VDD2.n5 4.46457
R1097 VDD2.n29 VDD2.n15 2.71565
R1098 VDD2.n14 VDD2.n0 2.71565
R1099 VDD2.n27 VDD2.n26 1.93989
R1100 VDD2.n12 VDD2.n11 1.93989
R1101 VDD2.n23 VDD2.n17 1.16414
R1102 VDD2.n8 VDD2.n2 1.16414
R1103 VDD2 VDD2.n30 0.864724
R1104 VDD2.n22 VDD2.n19 0.388379
R1105 VDD2.n7 VDD2.n4 0.388379
R1106 VDD2.n28 VDD2.n16 0.155672
R1107 VDD2.n21 VDD2.n16 0.155672
R1108 VDD2.n6 VDD2.n1 0.155672
R1109 VDD2.n13 VDD2.n1 0.155672
C0 VN VP 4.22013f
C1 VP VDD2 0.372219f
C2 VTAIL VP 1.26919f
C3 VP VDD1 1.18993f
C4 VN VDD2 0.972931f
C5 VTAIL VN 1.25505f
C6 VN VDD1 0.153667f
C7 VTAIL VDD2 3.06708f
C8 VDD1 VDD2 0.772713f
C9 VTAIL VDD1 3.0088f
C10 VDD2 B 3.104391f
C11 VDD1 B 4.83978f
C12 VTAIL B 3.82454f
C13 VN B 8.62443f
C14 VP B 6.611557f
C15 VDD2.n0 B 0.023673f
C16 VDD2.n1 B 0.017005f
C17 VDD2.n2 B 0.009138f
C18 VDD2.n3 B 0.016199f
C19 VDD2.n4 B 0.012594f
C20 VDD2.t0 B 0.036618f
C21 VDD2.n5 B 0.063532f
C22 VDD2.n6 B 0.187229f
C23 VDD2.n7 B 0.009138f
C24 VDD2.n8 B 0.009675f
C25 VDD2.n9 B 0.021599f
C26 VDD2.n10 B 0.046352f
C27 VDD2.n11 B 0.009675f
C28 VDD2.n12 B 0.009138f
C29 VDD2.n13 B 0.04256f
C30 VDD2.n14 B 0.329801f
C31 VDD2.n15 B 0.023673f
C32 VDD2.n16 B 0.017005f
C33 VDD2.n17 B 0.009138f
C34 VDD2.n18 B 0.016199f
C35 VDD2.n19 B 0.012594f
C36 VDD2.t1 B 0.036618f
C37 VDD2.n20 B 0.063532f
C38 VDD2.n21 B 0.187229f
C39 VDD2.n22 B 0.009138f
C40 VDD2.n23 B 0.009675f
C41 VDD2.n24 B 0.021599f
C42 VDD2.n25 B 0.046352f
C43 VDD2.n26 B 0.009675f
C44 VDD2.n27 B 0.009138f
C45 VDD2.n28 B 0.04256f
C46 VDD2.n29 B 0.037709f
C47 VDD2.n30 B 1.56808f
C48 VN.t1 B 0.893211f
C49 VN.t0 B 1.35748f
C50 VDD1.n0 B 0.022455f
C51 VDD1.n1 B 0.01613f
C52 VDD1.n2 B 0.008668f
C53 VDD1.n3 B 0.015365f
C54 VDD1.n4 B 0.011946f
C55 VDD1.t0 B 0.034733f
C56 VDD1.n5 B 0.060261f
C57 VDD1.n6 B 0.177591f
C58 VDD1.n7 B 0.008668f
C59 VDD1.n8 B 0.009177f
C60 VDD1.n9 B 0.020487f
C61 VDD1.n10 B 0.043966f
C62 VDD1.n11 B 0.009177f
C63 VDD1.n12 B 0.008668f
C64 VDD1.n13 B 0.040369f
C65 VDD1.n14 B 0.037049f
C66 VDD1.n15 B 0.022455f
C67 VDD1.n16 B 0.01613f
C68 VDD1.n17 B 0.008668f
C69 VDD1.n18 B 0.015365f
C70 VDD1.n19 B 0.011946f
C71 VDD1.t1 B 0.034733f
C72 VDD1.n20 B 0.060261f
C73 VDD1.n21 B 0.177591f
C74 VDD1.n22 B 0.008668f
C75 VDD1.n23 B 0.009177f
C76 VDD1.n24 B 0.020487f
C77 VDD1.n25 B 0.043966f
C78 VDD1.n26 B 0.009177f
C79 VDD1.n27 B 0.008668f
C80 VDD1.n28 B 0.040369f
C81 VDD1.n29 B 0.342248f
C82 VTAIL.n0 B 0.027338f
C83 VTAIL.n1 B 0.019638f
C84 VTAIL.n2 B 0.010553f
C85 VTAIL.n3 B 0.018707f
C86 VTAIL.n4 B 0.014544f
C87 VTAIL.t2 B 0.042287f
C88 VTAIL.n5 B 0.073368f
C89 VTAIL.n6 B 0.216216f
C90 VTAIL.n7 B 0.010553f
C91 VTAIL.n8 B 0.011174f
C92 VTAIL.n9 B 0.024943f
C93 VTAIL.n10 B 0.053528f
C94 VTAIL.n11 B 0.011174f
C95 VTAIL.n12 B 0.010553f
C96 VTAIL.n13 B 0.049149f
C97 VTAIL.n14 B 0.030014f
C98 VTAIL.n15 B 0.955949f
C99 VTAIL.n16 B 0.027338f
C100 VTAIL.n17 B 0.019638f
C101 VTAIL.n18 B 0.010553f
C102 VTAIL.n19 B 0.018707f
C103 VTAIL.n20 B 0.014544f
C104 VTAIL.t0 B 0.042287f
C105 VTAIL.n21 B 0.073368f
C106 VTAIL.n22 B 0.216216f
C107 VTAIL.n23 B 0.010553f
C108 VTAIL.n24 B 0.011174f
C109 VTAIL.n25 B 0.024943f
C110 VTAIL.n26 B 0.053528f
C111 VTAIL.n27 B 0.011174f
C112 VTAIL.n28 B 0.010553f
C113 VTAIL.n29 B 0.049149f
C114 VTAIL.n30 B 0.030014f
C115 VTAIL.n31 B 1.00327f
C116 VTAIL.n32 B 0.027338f
C117 VTAIL.n33 B 0.019638f
C118 VTAIL.n34 B 0.010553f
C119 VTAIL.n35 B 0.018707f
C120 VTAIL.n36 B 0.014544f
C121 VTAIL.t3 B 0.042287f
C122 VTAIL.n37 B 0.073368f
C123 VTAIL.n38 B 0.216216f
C124 VTAIL.n39 B 0.010553f
C125 VTAIL.n40 B 0.011174f
C126 VTAIL.n41 B 0.024943f
C127 VTAIL.n42 B 0.053528f
C128 VTAIL.n43 B 0.011174f
C129 VTAIL.n44 B 0.010553f
C130 VTAIL.n45 B 0.049149f
C131 VTAIL.n46 B 0.030014f
C132 VTAIL.n47 B 0.799252f
C133 VTAIL.n48 B 0.027338f
C134 VTAIL.n49 B 0.019638f
C135 VTAIL.n50 B 0.010553f
C136 VTAIL.n51 B 0.018707f
C137 VTAIL.n52 B 0.014544f
C138 VTAIL.t1 B 0.042287f
C139 VTAIL.n53 B 0.073368f
C140 VTAIL.n54 B 0.216216f
C141 VTAIL.n55 B 0.010553f
C142 VTAIL.n56 B 0.011174f
C143 VTAIL.n57 B 0.024943f
C144 VTAIL.n58 B 0.053528f
C145 VTAIL.n59 B 0.011174f
C146 VTAIL.n60 B 0.010553f
C147 VTAIL.n61 B 0.049149f
C148 VTAIL.n62 B 0.030014f
C149 VTAIL.n63 B 0.714835f
C150 VP.t1 B 1.36682f
C151 VP.t0 B 0.897291f
C152 VP.n0 B 1.85438f
.ends

