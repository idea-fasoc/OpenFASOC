* NGSPICE file created from diff_pair_sample_1150.ext - technology: sky130A

.subckt diff_pair_sample_1150 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t15 VP.t0 VDD1.t3 w_n2290_n1844# sky130_fd_pr__pfet_01v8 ad=0.7227 pd=4.71 as=0.7227 ps=4.71 w=4.38 l=0.99
X1 B.t11 B.t9 B.t10 w_n2290_n1844# sky130_fd_pr__pfet_01v8 ad=1.7082 pd=9.54 as=0 ps=0 w=4.38 l=0.99
X2 VDD2.t7 VN.t0 VTAIL.t7 w_n2290_n1844# sky130_fd_pr__pfet_01v8 ad=0.7227 pd=4.71 as=1.7082 ps=9.54 w=4.38 l=0.99
X3 VDD1.t2 VP.t1 VTAIL.t14 w_n2290_n1844# sky130_fd_pr__pfet_01v8 ad=0.7227 pd=4.71 as=0.7227 ps=4.71 w=4.38 l=0.99
X4 VTAIL.t2 VN.t1 VDD2.t6 w_n2290_n1844# sky130_fd_pr__pfet_01v8 ad=0.7227 pd=4.71 as=0.7227 ps=4.71 w=4.38 l=0.99
X5 VTAIL.t13 VP.t2 VDD1.t4 w_n2290_n1844# sky130_fd_pr__pfet_01v8 ad=1.7082 pd=9.54 as=0.7227 ps=4.71 w=4.38 l=0.99
X6 VDD2.t5 VN.t2 VTAIL.t6 w_n2290_n1844# sky130_fd_pr__pfet_01v8 ad=0.7227 pd=4.71 as=1.7082 ps=9.54 w=4.38 l=0.99
X7 VTAIL.t12 VP.t3 VDD1.t5 w_n2290_n1844# sky130_fd_pr__pfet_01v8 ad=1.7082 pd=9.54 as=0.7227 ps=4.71 w=4.38 l=0.99
X8 VTAIL.t0 VN.t3 VDD2.t4 w_n2290_n1844# sky130_fd_pr__pfet_01v8 ad=1.7082 pd=9.54 as=0.7227 ps=4.71 w=4.38 l=0.99
X9 VDD1.t6 VP.t4 VTAIL.t11 w_n2290_n1844# sky130_fd_pr__pfet_01v8 ad=0.7227 pd=4.71 as=1.7082 ps=9.54 w=4.38 l=0.99
X10 VDD1.t0 VP.t5 VTAIL.t10 w_n2290_n1844# sky130_fd_pr__pfet_01v8 ad=0.7227 pd=4.71 as=1.7082 ps=9.54 w=4.38 l=0.99
X11 B.t8 B.t6 B.t7 w_n2290_n1844# sky130_fd_pr__pfet_01v8 ad=1.7082 pd=9.54 as=0 ps=0 w=4.38 l=0.99
X12 VTAIL.t1 VN.t4 VDD2.t3 w_n2290_n1844# sky130_fd_pr__pfet_01v8 ad=1.7082 pd=9.54 as=0.7227 ps=4.71 w=4.38 l=0.99
X13 B.t5 B.t3 B.t4 w_n2290_n1844# sky130_fd_pr__pfet_01v8 ad=1.7082 pd=9.54 as=0 ps=0 w=4.38 l=0.99
X14 VDD2.t2 VN.t5 VTAIL.t3 w_n2290_n1844# sky130_fd_pr__pfet_01v8 ad=0.7227 pd=4.71 as=0.7227 ps=4.71 w=4.38 l=0.99
X15 VTAIL.t9 VP.t6 VDD1.t7 w_n2290_n1844# sky130_fd_pr__pfet_01v8 ad=0.7227 pd=4.71 as=0.7227 ps=4.71 w=4.38 l=0.99
X16 VDD2.t1 VN.t6 VTAIL.t4 w_n2290_n1844# sky130_fd_pr__pfet_01v8 ad=0.7227 pd=4.71 as=0.7227 ps=4.71 w=4.38 l=0.99
X17 B.t2 B.t0 B.t1 w_n2290_n1844# sky130_fd_pr__pfet_01v8 ad=1.7082 pd=9.54 as=0 ps=0 w=4.38 l=0.99
X18 VTAIL.t5 VN.t7 VDD2.t0 w_n2290_n1844# sky130_fd_pr__pfet_01v8 ad=0.7227 pd=4.71 as=0.7227 ps=4.71 w=4.38 l=0.99
X19 VDD1.t1 VP.t7 VTAIL.t8 w_n2290_n1844# sky130_fd_pr__pfet_01v8 ad=0.7227 pd=4.71 as=0.7227 ps=4.71 w=4.38 l=0.99
R0 VP.n5 VP.t2 161.457
R1 VP.n8 VP.n7 161.3
R2 VP.n9 VP.n4 161.3
R3 VP.n11 VP.n10 161.3
R4 VP.n13 VP.n3 161.3
R5 VP.n26 VP.n0 161.3
R6 VP.n24 VP.n23 161.3
R7 VP.n22 VP.n1 161.3
R8 VP.n21 VP.n20 161.3
R9 VP.n18 VP.n2 161.3
R10 VP.n17 VP.t3 146.304
R11 VP.n27 VP.t5 146.304
R12 VP.n14 VP.t4 146.304
R13 VP.n19 VP.t7 106.624
R14 VP.n25 VP.t0 106.624
R15 VP.n12 VP.t6 106.624
R16 VP.n6 VP.t1 106.624
R17 VP.n15 VP.n14 80.6037
R18 VP.n28 VP.n27 80.6037
R19 VP.n17 VP.n16 80.6037
R20 VP.n18 VP.n17 55.824
R21 VP.n27 VP.n26 55.824
R22 VP.n14 VP.n13 55.824
R23 VP.n6 VP.n5 46.9382
R24 VP.n8 VP.n5 43.9713
R25 VP.n20 VP.n1 40.577
R26 VP.n24 VP.n1 40.577
R27 VP.n11 VP.n4 40.577
R28 VP.n7 VP.n4 40.577
R29 VP.n16 VP.n15 37.7893
R30 VP.n19 VP.n18 16.7229
R31 VP.n26 VP.n25 16.7229
R32 VP.n13 VP.n12 16.7229
R33 VP.n20 VP.n19 7.86989
R34 VP.n25 VP.n24 7.86989
R35 VP.n12 VP.n11 7.86989
R36 VP.n7 VP.n6 7.86989
R37 VP.n15 VP.n3 0.285035
R38 VP.n16 VP.n2 0.285035
R39 VP.n28 VP.n0 0.285035
R40 VP.n9 VP.n8 0.189894
R41 VP.n10 VP.n9 0.189894
R42 VP.n10 VP.n3 0.189894
R43 VP.n21 VP.n2 0.189894
R44 VP.n22 VP.n21 0.189894
R45 VP.n23 VP.n22 0.189894
R46 VP.n23 VP.n0 0.189894
R47 VP VP.n28 0.146778
R48 VDD1 VDD1.n0 112.504
R49 VDD1.n3 VDD1.n2 112.391
R50 VDD1.n3 VDD1.n1 112.391
R51 VDD1.n5 VDD1.n4 111.877
R52 VDD1.n5 VDD1.n3 33.1949
R53 VDD1.n4 VDD1.t7 7.42173
R54 VDD1.n4 VDD1.t6 7.42173
R55 VDD1.n0 VDD1.t4 7.42173
R56 VDD1.n0 VDD1.t2 7.42173
R57 VDD1.n2 VDD1.t3 7.42173
R58 VDD1.n2 VDD1.t0 7.42173
R59 VDD1.n1 VDD1.t5 7.42173
R60 VDD1.n1 VDD1.t1 7.42173
R61 VDD1 VDD1.n5 0.511276
R62 VTAIL.n11 VTAIL.t13 102.62
R63 VTAIL.n10 VTAIL.t6 102.62
R64 VTAIL.n7 VTAIL.t1 102.62
R65 VTAIL.n15 VTAIL.t7 102.62
R66 VTAIL.n2 VTAIL.t0 102.62
R67 VTAIL.n3 VTAIL.t10 102.62
R68 VTAIL.n6 VTAIL.t12 102.62
R69 VTAIL.n14 VTAIL.t11 102.62
R70 VTAIL.n13 VTAIL.n12 95.1987
R71 VTAIL.n9 VTAIL.n8 95.1987
R72 VTAIL.n1 VTAIL.n0 95.1985
R73 VTAIL.n5 VTAIL.n4 95.1985
R74 VTAIL.n15 VTAIL.n14 17.2807
R75 VTAIL.n7 VTAIL.n6 17.2807
R76 VTAIL.n0 VTAIL.t3 7.42173
R77 VTAIL.n0 VTAIL.t5 7.42173
R78 VTAIL.n4 VTAIL.t8 7.42173
R79 VTAIL.n4 VTAIL.t15 7.42173
R80 VTAIL.n12 VTAIL.t14 7.42173
R81 VTAIL.n12 VTAIL.t9 7.42173
R82 VTAIL.n8 VTAIL.t4 7.42173
R83 VTAIL.n8 VTAIL.t2 7.42173
R84 VTAIL.n9 VTAIL.n7 1.13843
R85 VTAIL.n10 VTAIL.n9 1.13843
R86 VTAIL.n13 VTAIL.n11 1.13843
R87 VTAIL.n14 VTAIL.n13 1.13843
R88 VTAIL.n6 VTAIL.n5 1.13843
R89 VTAIL.n5 VTAIL.n3 1.13843
R90 VTAIL.n2 VTAIL.n1 1.13843
R91 VTAIL VTAIL.n15 1.08024
R92 VTAIL.n11 VTAIL.n10 0.470328
R93 VTAIL.n3 VTAIL.n2 0.470328
R94 VTAIL VTAIL.n1 0.0586897
R95 B.n225 B.n72 585
R96 B.n224 B.n223 585
R97 B.n222 B.n73 585
R98 B.n221 B.n220 585
R99 B.n219 B.n74 585
R100 B.n218 B.n217 585
R101 B.n216 B.n75 585
R102 B.n215 B.n214 585
R103 B.n213 B.n76 585
R104 B.n212 B.n211 585
R105 B.n210 B.n77 585
R106 B.n209 B.n208 585
R107 B.n207 B.n78 585
R108 B.n206 B.n205 585
R109 B.n204 B.n79 585
R110 B.n203 B.n202 585
R111 B.n201 B.n80 585
R112 B.n200 B.n199 585
R113 B.n198 B.n81 585
R114 B.n196 B.n195 585
R115 B.n194 B.n84 585
R116 B.n193 B.n192 585
R117 B.n191 B.n85 585
R118 B.n190 B.n189 585
R119 B.n188 B.n86 585
R120 B.n187 B.n186 585
R121 B.n185 B.n87 585
R122 B.n184 B.n183 585
R123 B.n182 B.n88 585
R124 B.n181 B.n180 585
R125 B.n176 B.n89 585
R126 B.n175 B.n174 585
R127 B.n173 B.n90 585
R128 B.n172 B.n171 585
R129 B.n170 B.n91 585
R130 B.n169 B.n168 585
R131 B.n167 B.n92 585
R132 B.n166 B.n165 585
R133 B.n164 B.n93 585
R134 B.n163 B.n162 585
R135 B.n161 B.n94 585
R136 B.n160 B.n159 585
R137 B.n158 B.n95 585
R138 B.n157 B.n156 585
R139 B.n155 B.n96 585
R140 B.n154 B.n153 585
R141 B.n152 B.n97 585
R142 B.n151 B.n150 585
R143 B.n227 B.n226 585
R144 B.n228 B.n71 585
R145 B.n230 B.n229 585
R146 B.n231 B.n70 585
R147 B.n233 B.n232 585
R148 B.n234 B.n69 585
R149 B.n236 B.n235 585
R150 B.n237 B.n68 585
R151 B.n239 B.n238 585
R152 B.n240 B.n67 585
R153 B.n242 B.n241 585
R154 B.n243 B.n66 585
R155 B.n245 B.n244 585
R156 B.n246 B.n65 585
R157 B.n248 B.n247 585
R158 B.n249 B.n64 585
R159 B.n251 B.n250 585
R160 B.n252 B.n63 585
R161 B.n254 B.n253 585
R162 B.n255 B.n62 585
R163 B.n257 B.n256 585
R164 B.n258 B.n61 585
R165 B.n260 B.n259 585
R166 B.n261 B.n60 585
R167 B.n263 B.n262 585
R168 B.n264 B.n59 585
R169 B.n266 B.n265 585
R170 B.n267 B.n58 585
R171 B.n269 B.n268 585
R172 B.n270 B.n57 585
R173 B.n272 B.n271 585
R174 B.n273 B.n56 585
R175 B.n275 B.n274 585
R176 B.n276 B.n55 585
R177 B.n278 B.n277 585
R178 B.n279 B.n54 585
R179 B.n281 B.n280 585
R180 B.n282 B.n53 585
R181 B.n284 B.n283 585
R182 B.n285 B.n52 585
R183 B.n287 B.n286 585
R184 B.n288 B.n51 585
R185 B.n290 B.n289 585
R186 B.n291 B.n50 585
R187 B.n293 B.n292 585
R188 B.n294 B.n49 585
R189 B.n296 B.n295 585
R190 B.n297 B.n48 585
R191 B.n299 B.n298 585
R192 B.n300 B.n47 585
R193 B.n302 B.n301 585
R194 B.n303 B.n46 585
R195 B.n305 B.n304 585
R196 B.n306 B.n45 585
R197 B.n308 B.n307 585
R198 B.n309 B.n44 585
R199 B.n383 B.n382 585
R200 B.n381 B.n16 585
R201 B.n380 B.n379 585
R202 B.n378 B.n17 585
R203 B.n377 B.n376 585
R204 B.n375 B.n18 585
R205 B.n374 B.n373 585
R206 B.n372 B.n19 585
R207 B.n371 B.n370 585
R208 B.n369 B.n20 585
R209 B.n368 B.n367 585
R210 B.n366 B.n21 585
R211 B.n365 B.n364 585
R212 B.n363 B.n22 585
R213 B.n362 B.n361 585
R214 B.n360 B.n23 585
R215 B.n359 B.n358 585
R216 B.n357 B.n24 585
R217 B.n356 B.n355 585
R218 B.n353 B.n25 585
R219 B.n352 B.n351 585
R220 B.n350 B.n28 585
R221 B.n349 B.n348 585
R222 B.n347 B.n29 585
R223 B.n346 B.n345 585
R224 B.n344 B.n30 585
R225 B.n343 B.n342 585
R226 B.n341 B.n31 585
R227 B.n340 B.n339 585
R228 B.n338 B.n337 585
R229 B.n336 B.n35 585
R230 B.n335 B.n334 585
R231 B.n333 B.n36 585
R232 B.n332 B.n331 585
R233 B.n330 B.n37 585
R234 B.n329 B.n328 585
R235 B.n327 B.n38 585
R236 B.n326 B.n325 585
R237 B.n324 B.n39 585
R238 B.n323 B.n322 585
R239 B.n321 B.n40 585
R240 B.n320 B.n319 585
R241 B.n318 B.n41 585
R242 B.n317 B.n316 585
R243 B.n315 B.n42 585
R244 B.n314 B.n313 585
R245 B.n312 B.n43 585
R246 B.n311 B.n310 585
R247 B.n384 B.n15 585
R248 B.n386 B.n385 585
R249 B.n387 B.n14 585
R250 B.n389 B.n388 585
R251 B.n390 B.n13 585
R252 B.n392 B.n391 585
R253 B.n393 B.n12 585
R254 B.n395 B.n394 585
R255 B.n396 B.n11 585
R256 B.n398 B.n397 585
R257 B.n399 B.n10 585
R258 B.n401 B.n400 585
R259 B.n402 B.n9 585
R260 B.n404 B.n403 585
R261 B.n405 B.n8 585
R262 B.n407 B.n406 585
R263 B.n408 B.n7 585
R264 B.n410 B.n409 585
R265 B.n411 B.n6 585
R266 B.n413 B.n412 585
R267 B.n414 B.n5 585
R268 B.n416 B.n415 585
R269 B.n417 B.n4 585
R270 B.n419 B.n418 585
R271 B.n420 B.n3 585
R272 B.n422 B.n421 585
R273 B.n423 B.n0 585
R274 B.n2 B.n1 585
R275 B.n112 B.n111 585
R276 B.n113 B.n110 585
R277 B.n115 B.n114 585
R278 B.n116 B.n109 585
R279 B.n118 B.n117 585
R280 B.n119 B.n108 585
R281 B.n121 B.n120 585
R282 B.n122 B.n107 585
R283 B.n124 B.n123 585
R284 B.n125 B.n106 585
R285 B.n127 B.n126 585
R286 B.n128 B.n105 585
R287 B.n130 B.n129 585
R288 B.n131 B.n104 585
R289 B.n133 B.n132 585
R290 B.n134 B.n103 585
R291 B.n136 B.n135 585
R292 B.n137 B.n102 585
R293 B.n139 B.n138 585
R294 B.n140 B.n101 585
R295 B.n142 B.n141 585
R296 B.n143 B.n100 585
R297 B.n145 B.n144 585
R298 B.n146 B.n99 585
R299 B.n148 B.n147 585
R300 B.n149 B.n98 585
R301 B.n150 B.n149 502.111
R302 B.n226 B.n225 502.111
R303 B.n310 B.n309 502.111
R304 B.n382 B.n15 502.111
R305 B.n177 B.t0 309.483
R306 B.n82 B.t6 309.483
R307 B.n32 B.t3 309.483
R308 B.n26 B.t9 309.483
R309 B.n425 B.n424 256.663
R310 B.n424 B.n423 235.042
R311 B.n424 B.n2 235.042
R312 B.n150 B.n97 163.367
R313 B.n154 B.n97 163.367
R314 B.n155 B.n154 163.367
R315 B.n156 B.n155 163.367
R316 B.n156 B.n95 163.367
R317 B.n160 B.n95 163.367
R318 B.n161 B.n160 163.367
R319 B.n162 B.n161 163.367
R320 B.n162 B.n93 163.367
R321 B.n166 B.n93 163.367
R322 B.n167 B.n166 163.367
R323 B.n168 B.n167 163.367
R324 B.n168 B.n91 163.367
R325 B.n172 B.n91 163.367
R326 B.n173 B.n172 163.367
R327 B.n174 B.n173 163.367
R328 B.n174 B.n89 163.367
R329 B.n181 B.n89 163.367
R330 B.n182 B.n181 163.367
R331 B.n183 B.n182 163.367
R332 B.n183 B.n87 163.367
R333 B.n187 B.n87 163.367
R334 B.n188 B.n187 163.367
R335 B.n189 B.n188 163.367
R336 B.n189 B.n85 163.367
R337 B.n193 B.n85 163.367
R338 B.n194 B.n193 163.367
R339 B.n195 B.n194 163.367
R340 B.n195 B.n81 163.367
R341 B.n200 B.n81 163.367
R342 B.n201 B.n200 163.367
R343 B.n202 B.n201 163.367
R344 B.n202 B.n79 163.367
R345 B.n206 B.n79 163.367
R346 B.n207 B.n206 163.367
R347 B.n208 B.n207 163.367
R348 B.n208 B.n77 163.367
R349 B.n212 B.n77 163.367
R350 B.n213 B.n212 163.367
R351 B.n214 B.n213 163.367
R352 B.n214 B.n75 163.367
R353 B.n218 B.n75 163.367
R354 B.n219 B.n218 163.367
R355 B.n220 B.n219 163.367
R356 B.n220 B.n73 163.367
R357 B.n224 B.n73 163.367
R358 B.n225 B.n224 163.367
R359 B.n309 B.n308 163.367
R360 B.n308 B.n45 163.367
R361 B.n304 B.n45 163.367
R362 B.n304 B.n303 163.367
R363 B.n303 B.n302 163.367
R364 B.n302 B.n47 163.367
R365 B.n298 B.n47 163.367
R366 B.n298 B.n297 163.367
R367 B.n297 B.n296 163.367
R368 B.n296 B.n49 163.367
R369 B.n292 B.n49 163.367
R370 B.n292 B.n291 163.367
R371 B.n291 B.n290 163.367
R372 B.n290 B.n51 163.367
R373 B.n286 B.n51 163.367
R374 B.n286 B.n285 163.367
R375 B.n285 B.n284 163.367
R376 B.n284 B.n53 163.367
R377 B.n280 B.n53 163.367
R378 B.n280 B.n279 163.367
R379 B.n279 B.n278 163.367
R380 B.n278 B.n55 163.367
R381 B.n274 B.n55 163.367
R382 B.n274 B.n273 163.367
R383 B.n273 B.n272 163.367
R384 B.n272 B.n57 163.367
R385 B.n268 B.n57 163.367
R386 B.n268 B.n267 163.367
R387 B.n267 B.n266 163.367
R388 B.n266 B.n59 163.367
R389 B.n262 B.n59 163.367
R390 B.n262 B.n261 163.367
R391 B.n261 B.n260 163.367
R392 B.n260 B.n61 163.367
R393 B.n256 B.n61 163.367
R394 B.n256 B.n255 163.367
R395 B.n255 B.n254 163.367
R396 B.n254 B.n63 163.367
R397 B.n250 B.n63 163.367
R398 B.n250 B.n249 163.367
R399 B.n249 B.n248 163.367
R400 B.n248 B.n65 163.367
R401 B.n244 B.n65 163.367
R402 B.n244 B.n243 163.367
R403 B.n243 B.n242 163.367
R404 B.n242 B.n67 163.367
R405 B.n238 B.n67 163.367
R406 B.n238 B.n237 163.367
R407 B.n237 B.n236 163.367
R408 B.n236 B.n69 163.367
R409 B.n232 B.n69 163.367
R410 B.n232 B.n231 163.367
R411 B.n231 B.n230 163.367
R412 B.n230 B.n71 163.367
R413 B.n226 B.n71 163.367
R414 B.n382 B.n381 163.367
R415 B.n381 B.n380 163.367
R416 B.n380 B.n17 163.367
R417 B.n376 B.n17 163.367
R418 B.n376 B.n375 163.367
R419 B.n375 B.n374 163.367
R420 B.n374 B.n19 163.367
R421 B.n370 B.n19 163.367
R422 B.n370 B.n369 163.367
R423 B.n369 B.n368 163.367
R424 B.n368 B.n21 163.367
R425 B.n364 B.n21 163.367
R426 B.n364 B.n363 163.367
R427 B.n363 B.n362 163.367
R428 B.n362 B.n23 163.367
R429 B.n358 B.n23 163.367
R430 B.n358 B.n357 163.367
R431 B.n357 B.n356 163.367
R432 B.n356 B.n25 163.367
R433 B.n351 B.n25 163.367
R434 B.n351 B.n350 163.367
R435 B.n350 B.n349 163.367
R436 B.n349 B.n29 163.367
R437 B.n345 B.n29 163.367
R438 B.n345 B.n344 163.367
R439 B.n344 B.n343 163.367
R440 B.n343 B.n31 163.367
R441 B.n339 B.n31 163.367
R442 B.n339 B.n338 163.367
R443 B.n338 B.n35 163.367
R444 B.n334 B.n35 163.367
R445 B.n334 B.n333 163.367
R446 B.n333 B.n332 163.367
R447 B.n332 B.n37 163.367
R448 B.n328 B.n37 163.367
R449 B.n328 B.n327 163.367
R450 B.n327 B.n326 163.367
R451 B.n326 B.n39 163.367
R452 B.n322 B.n39 163.367
R453 B.n322 B.n321 163.367
R454 B.n321 B.n320 163.367
R455 B.n320 B.n41 163.367
R456 B.n316 B.n41 163.367
R457 B.n316 B.n315 163.367
R458 B.n315 B.n314 163.367
R459 B.n314 B.n43 163.367
R460 B.n310 B.n43 163.367
R461 B.n386 B.n15 163.367
R462 B.n387 B.n386 163.367
R463 B.n388 B.n387 163.367
R464 B.n388 B.n13 163.367
R465 B.n392 B.n13 163.367
R466 B.n393 B.n392 163.367
R467 B.n394 B.n393 163.367
R468 B.n394 B.n11 163.367
R469 B.n398 B.n11 163.367
R470 B.n399 B.n398 163.367
R471 B.n400 B.n399 163.367
R472 B.n400 B.n9 163.367
R473 B.n404 B.n9 163.367
R474 B.n405 B.n404 163.367
R475 B.n406 B.n405 163.367
R476 B.n406 B.n7 163.367
R477 B.n410 B.n7 163.367
R478 B.n411 B.n410 163.367
R479 B.n412 B.n411 163.367
R480 B.n412 B.n5 163.367
R481 B.n416 B.n5 163.367
R482 B.n417 B.n416 163.367
R483 B.n418 B.n417 163.367
R484 B.n418 B.n3 163.367
R485 B.n422 B.n3 163.367
R486 B.n423 B.n422 163.367
R487 B.n112 B.n2 163.367
R488 B.n113 B.n112 163.367
R489 B.n114 B.n113 163.367
R490 B.n114 B.n109 163.367
R491 B.n118 B.n109 163.367
R492 B.n119 B.n118 163.367
R493 B.n120 B.n119 163.367
R494 B.n120 B.n107 163.367
R495 B.n124 B.n107 163.367
R496 B.n125 B.n124 163.367
R497 B.n126 B.n125 163.367
R498 B.n126 B.n105 163.367
R499 B.n130 B.n105 163.367
R500 B.n131 B.n130 163.367
R501 B.n132 B.n131 163.367
R502 B.n132 B.n103 163.367
R503 B.n136 B.n103 163.367
R504 B.n137 B.n136 163.367
R505 B.n138 B.n137 163.367
R506 B.n138 B.n101 163.367
R507 B.n142 B.n101 163.367
R508 B.n143 B.n142 163.367
R509 B.n144 B.n143 163.367
R510 B.n144 B.n99 163.367
R511 B.n148 B.n99 163.367
R512 B.n149 B.n148 163.367
R513 B.n82 B.t7 149.964
R514 B.n32 B.t5 149.964
R515 B.n177 B.t1 149.959
R516 B.n26 B.t11 149.959
R517 B.n83 B.t8 124.364
R518 B.n33 B.t4 124.364
R519 B.n178 B.t2 124.359
R520 B.n27 B.t10 124.359
R521 B.n179 B.n178 59.5399
R522 B.n197 B.n83 59.5399
R523 B.n34 B.n33 59.5399
R524 B.n354 B.n27 59.5399
R525 B.n384 B.n383 32.6249
R526 B.n311 B.n44 32.6249
R527 B.n227 B.n72 32.6249
R528 B.n151 B.n98 32.6249
R529 B.n178 B.n177 25.6005
R530 B.n83 B.n82 25.6005
R531 B.n33 B.n32 25.6005
R532 B.n27 B.n26 25.6005
R533 B B.n425 18.0485
R534 B.n385 B.n384 10.6151
R535 B.n385 B.n14 10.6151
R536 B.n389 B.n14 10.6151
R537 B.n390 B.n389 10.6151
R538 B.n391 B.n390 10.6151
R539 B.n391 B.n12 10.6151
R540 B.n395 B.n12 10.6151
R541 B.n396 B.n395 10.6151
R542 B.n397 B.n396 10.6151
R543 B.n397 B.n10 10.6151
R544 B.n401 B.n10 10.6151
R545 B.n402 B.n401 10.6151
R546 B.n403 B.n402 10.6151
R547 B.n403 B.n8 10.6151
R548 B.n407 B.n8 10.6151
R549 B.n408 B.n407 10.6151
R550 B.n409 B.n408 10.6151
R551 B.n409 B.n6 10.6151
R552 B.n413 B.n6 10.6151
R553 B.n414 B.n413 10.6151
R554 B.n415 B.n414 10.6151
R555 B.n415 B.n4 10.6151
R556 B.n419 B.n4 10.6151
R557 B.n420 B.n419 10.6151
R558 B.n421 B.n420 10.6151
R559 B.n421 B.n0 10.6151
R560 B.n383 B.n16 10.6151
R561 B.n379 B.n16 10.6151
R562 B.n379 B.n378 10.6151
R563 B.n378 B.n377 10.6151
R564 B.n377 B.n18 10.6151
R565 B.n373 B.n18 10.6151
R566 B.n373 B.n372 10.6151
R567 B.n372 B.n371 10.6151
R568 B.n371 B.n20 10.6151
R569 B.n367 B.n20 10.6151
R570 B.n367 B.n366 10.6151
R571 B.n366 B.n365 10.6151
R572 B.n365 B.n22 10.6151
R573 B.n361 B.n22 10.6151
R574 B.n361 B.n360 10.6151
R575 B.n360 B.n359 10.6151
R576 B.n359 B.n24 10.6151
R577 B.n355 B.n24 10.6151
R578 B.n353 B.n352 10.6151
R579 B.n352 B.n28 10.6151
R580 B.n348 B.n28 10.6151
R581 B.n348 B.n347 10.6151
R582 B.n347 B.n346 10.6151
R583 B.n346 B.n30 10.6151
R584 B.n342 B.n30 10.6151
R585 B.n342 B.n341 10.6151
R586 B.n341 B.n340 10.6151
R587 B.n337 B.n336 10.6151
R588 B.n336 B.n335 10.6151
R589 B.n335 B.n36 10.6151
R590 B.n331 B.n36 10.6151
R591 B.n331 B.n330 10.6151
R592 B.n330 B.n329 10.6151
R593 B.n329 B.n38 10.6151
R594 B.n325 B.n38 10.6151
R595 B.n325 B.n324 10.6151
R596 B.n324 B.n323 10.6151
R597 B.n323 B.n40 10.6151
R598 B.n319 B.n40 10.6151
R599 B.n319 B.n318 10.6151
R600 B.n318 B.n317 10.6151
R601 B.n317 B.n42 10.6151
R602 B.n313 B.n42 10.6151
R603 B.n313 B.n312 10.6151
R604 B.n312 B.n311 10.6151
R605 B.n307 B.n44 10.6151
R606 B.n307 B.n306 10.6151
R607 B.n306 B.n305 10.6151
R608 B.n305 B.n46 10.6151
R609 B.n301 B.n46 10.6151
R610 B.n301 B.n300 10.6151
R611 B.n300 B.n299 10.6151
R612 B.n299 B.n48 10.6151
R613 B.n295 B.n48 10.6151
R614 B.n295 B.n294 10.6151
R615 B.n294 B.n293 10.6151
R616 B.n293 B.n50 10.6151
R617 B.n289 B.n50 10.6151
R618 B.n289 B.n288 10.6151
R619 B.n288 B.n287 10.6151
R620 B.n287 B.n52 10.6151
R621 B.n283 B.n52 10.6151
R622 B.n283 B.n282 10.6151
R623 B.n282 B.n281 10.6151
R624 B.n281 B.n54 10.6151
R625 B.n277 B.n54 10.6151
R626 B.n277 B.n276 10.6151
R627 B.n276 B.n275 10.6151
R628 B.n275 B.n56 10.6151
R629 B.n271 B.n56 10.6151
R630 B.n271 B.n270 10.6151
R631 B.n270 B.n269 10.6151
R632 B.n269 B.n58 10.6151
R633 B.n265 B.n58 10.6151
R634 B.n265 B.n264 10.6151
R635 B.n264 B.n263 10.6151
R636 B.n263 B.n60 10.6151
R637 B.n259 B.n60 10.6151
R638 B.n259 B.n258 10.6151
R639 B.n258 B.n257 10.6151
R640 B.n257 B.n62 10.6151
R641 B.n253 B.n62 10.6151
R642 B.n253 B.n252 10.6151
R643 B.n252 B.n251 10.6151
R644 B.n251 B.n64 10.6151
R645 B.n247 B.n64 10.6151
R646 B.n247 B.n246 10.6151
R647 B.n246 B.n245 10.6151
R648 B.n245 B.n66 10.6151
R649 B.n241 B.n66 10.6151
R650 B.n241 B.n240 10.6151
R651 B.n240 B.n239 10.6151
R652 B.n239 B.n68 10.6151
R653 B.n235 B.n68 10.6151
R654 B.n235 B.n234 10.6151
R655 B.n234 B.n233 10.6151
R656 B.n233 B.n70 10.6151
R657 B.n229 B.n70 10.6151
R658 B.n229 B.n228 10.6151
R659 B.n228 B.n227 10.6151
R660 B.n111 B.n1 10.6151
R661 B.n111 B.n110 10.6151
R662 B.n115 B.n110 10.6151
R663 B.n116 B.n115 10.6151
R664 B.n117 B.n116 10.6151
R665 B.n117 B.n108 10.6151
R666 B.n121 B.n108 10.6151
R667 B.n122 B.n121 10.6151
R668 B.n123 B.n122 10.6151
R669 B.n123 B.n106 10.6151
R670 B.n127 B.n106 10.6151
R671 B.n128 B.n127 10.6151
R672 B.n129 B.n128 10.6151
R673 B.n129 B.n104 10.6151
R674 B.n133 B.n104 10.6151
R675 B.n134 B.n133 10.6151
R676 B.n135 B.n134 10.6151
R677 B.n135 B.n102 10.6151
R678 B.n139 B.n102 10.6151
R679 B.n140 B.n139 10.6151
R680 B.n141 B.n140 10.6151
R681 B.n141 B.n100 10.6151
R682 B.n145 B.n100 10.6151
R683 B.n146 B.n145 10.6151
R684 B.n147 B.n146 10.6151
R685 B.n147 B.n98 10.6151
R686 B.n152 B.n151 10.6151
R687 B.n153 B.n152 10.6151
R688 B.n153 B.n96 10.6151
R689 B.n157 B.n96 10.6151
R690 B.n158 B.n157 10.6151
R691 B.n159 B.n158 10.6151
R692 B.n159 B.n94 10.6151
R693 B.n163 B.n94 10.6151
R694 B.n164 B.n163 10.6151
R695 B.n165 B.n164 10.6151
R696 B.n165 B.n92 10.6151
R697 B.n169 B.n92 10.6151
R698 B.n170 B.n169 10.6151
R699 B.n171 B.n170 10.6151
R700 B.n171 B.n90 10.6151
R701 B.n175 B.n90 10.6151
R702 B.n176 B.n175 10.6151
R703 B.n180 B.n176 10.6151
R704 B.n184 B.n88 10.6151
R705 B.n185 B.n184 10.6151
R706 B.n186 B.n185 10.6151
R707 B.n186 B.n86 10.6151
R708 B.n190 B.n86 10.6151
R709 B.n191 B.n190 10.6151
R710 B.n192 B.n191 10.6151
R711 B.n192 B.n84 10.6151
R712 B.n196 B.n84 10.6151
R713 B.n199 B.n198 10.6151
R714 B.n199 B.n80 10.6151
R715 B.n203 B.n80 10.6151
R716 B.n204 B.n203 10.6151
R717 B.n205 B.n204 10.6151
R718 B.n205 B.n78 10.6151
R719 B.n209 B.n78 10.6151
R720 B.n210 B.n209 10.6151
R721 B.n211 B.n210 10.6151
R722 B.n211 B.n76 10.6151
R723 B.n215 B.n76 10.6151
R724 B.n216 B.n215 10.6151
R725 B.n217 B.n216 10.6151
R726 B.n217 B.n74 10.6151
R727 B.n221 B.n74 10.6151
R728 B.n222 B.n221 10.6151
R729 B.n223 B.n222 10.6151
R730 B.n223 B.n72 10.6151
R731 B.n355 B.n354 9.36635
R732 B.n337 B.n34 9.36635
R733 B.n180 B.n179 9.36635
R734 B.n198 B.n197 9.36635
R735 B.n425 B.n0 8.11757
R736 B.n425 B.n1 8.11757
R737 B.n354 B.n353 1.24928
R738 B.n340 B.n34 1.24928
R739 B.n179 B.n88 1.24928
R740 B.n197 B.n196 1.24928
R741 VN.n2 VN.t3 161.457
R742 VN.n15 VN.t2 161.457
R743 VN.n23 VN.n13 161.3
R744 VN.n21 VN.n20 161.3
R745 VN.n19 VN.n14 161.3
R746 VN.n18 VN.n17 161.3
R747 VN.n10 VN.n0 161.3
R748 VN.n8 VN.n7 161.3
R749 VN.n6 VN.n1 161.3
R750 VN.n5 VN.n4 161.3
R751 VN.n11 VN.t0 146.304
R752 VN.n24 VN.t4 146.304
R753 VN.n3 VN.t5 106.624
R754 VN.n9 VN.t7 106.624
R755 VN.n16 VN.t1 106.624
R756 VN.n22 VN.t6 106.624
R757 VN.n25 VN.n24 80.6037
R758 VN.n12 VN.n11 80.6037
R759 VN.n11 VN.n10 55.824
R760 VN.n24 VN.n23 55.824
R761 VN.n3 VN.n2 46.9382
R762 VN.n16 VN.n15 46.9382
R763 VN.n18 VN.n15 43.9713
R764 VN.n5 VN.n2 43.9713
R765 VN.n4 VN.n1 40.577
R766 VN.n8 VN.n1 40.577
R767 VN.n17 VN.n14 40.577
R768 VN.n21 VN.n14 40.577
R769 VN VN.n25 38.0748
R770 VN.n10 VN.n9 16.7229
R771 VN.n23 VN.n22 16.7229
R772 VN.n4 VN.n3 7.86989
R773 VN.n9 VN.n8 7.86989
R774 VN.n17 VN.n16 7.86989
R775 VN.n22 VN.n21 7.86989
R776 VN.n25 VN.n13 0.285035
R777 VN.n12 VN.n0 0.285035
R778 VN.n20 VN.n13 0.189894
R779 VN.n20 VN.n19 0.189894
R780 VN.n19 VN.n18 0.189894
R781 VN.n6 VN.n5 0.189894
R782 VN.n7 VN.n6 0.189894
R783 VN.n7 VN.n0 0.189894
R784 VN VN.n12 0.146778
R785 VDD2.n2 VDD2.n1 112.391
R786 VDD2.n2 VDD2.n0 112.391
R787 VDD2 VDD2.n5 112.388
R788 VDD2.n4 VDD2.n3 111.877
R789 VDD2.n4 VDD2.n2 32.6118
R790 VDD2.n5 VDD2.t6 7.42173
R791 VDD2.n5 VDD2.t5 7.42173
R792 VDD2.n3 VDD2.t3 7.42173
R793 VDD2.n3 VDD2.t1 7.42173
R794 VDD2.n1 VDD2.t0 7.42173
R795 VDD2.n1 VDD2.t7 7.42173
R796 VDD2.n0 VDD2.t4 7.42173
R797 VDD2.n0 VDD2.t2 7.42173
R798 VDD2 VDD2.n4 0.627655
C0 B VN 0.770708f
C1 VTAIL VN 2.8901f
C2 B VP 1.2524f
C3 B VDD2 0.998748f
C4 VTAIL VP 2.9042f
C5 w_n2290_n1844# VN 4.05705f
C6 VTAIL VDD2 5.07633f
C7 B VDD1 0.953047f
C8 VDD1 VTAIL 5.03271f
C9 w_n2290_n1844# VDD2 1.25246f
C10 VP w_n2290_n1844# 4.34921f
C11 VDD1 w_n2290_n1844# 1.20589f
C12 VP VN 4.28298f
C13 VDD2 VN 2.61797f
C14 VDD1 VN 0.153292f
C15 VP VDD2 0.353194f
C16 VDD1 VP 2.81689f
C17 VDD1 VDD2 0.971179f
C18 B VTAIL 1.89432f
C19 B w_n2290_n1844# 5.51679f
C20 VTAIL w_n2290_n1844# 2.28352f
C21 VDD2 VSUBS 1.078389f
C22 VDD1 VSUBS 1.43462f
C23 VTAIL VSUBS 0.485555f
C24 VN VSUBS 4.45611f
C25 VP VSUBS 1.551301f
C26 B VSUBS 2.441043f
C27 w_n2290_n1844# VSUBS 53.063896f
C28 VDD2.t4 VSUBS 0.088401f
C29 VDD2.t2 VSUBS 0.088401f
C30 VDD2.n0 VSUBS 0.535783f
C31 VDD2.t0 VSUBS 0.088401f
C32 VDD2.t7 VSUBS 0.088401f
C33 VDD2.n1 VSUBS 0.535783f
C34 VDD2.n2 VSUBS 2.25261f
C35 VDD2.t3 VSUBS 0.088401f
C36 VDD2.t1 VSUBS 0.088401f
C37 VDD2.n3 VSUBS 0.533409f
C38 VDD2.n4 VSUBS 1.98946f
C39 VDD2.t6 VSUBS 0.088401f
C40 VDD2.t5 VSUBS 0.088401f
C41 VDD2.n5 VSUBS 0.535763f
C42 VN.n0 VSUBS 0.076919f
C43 VN.t7 VSUBS 0.64719f
C44 VN.n1 VSUBS 0.046558f
C45 VN.t3 VSUBS 0.769208f
C46 VN.n2 VSUBS 0.367669f
C47 VN.t5 VSUBS 0.64719f
C48 VN.n3 VSUBS 0.336386f
C49 VN.n4 VSUBS 0.07808f
C50 VN.n5 VSUBS 0.245365f
C51 VN.n6 VSUBS 0.057645f
C52 VN.n7 VSUBS 0.057645f
C53 VN.n8 VSUBS 0.07808f
C54 VN.n9 VSUBS 0.286272f
C55 VN.n10 VSUBS 0.077849f
C56 VN.t0 VSUBS 0.734086f
C57 VN.n11 VSUBS 0.37385f
C58 VN.n12 VSUBS 0.053986f
C59 VN.n13 VSUBS 0.076919f
C60 VN.t6 VSUBS 0.64719f
C61 VN.n14 VSUBS 0.046558f
C62 VN.t2 VSUBS 0.769208f
C63 VN.n15 VSUBS 0.367669f
C64 VN.t1 VSUBS 0.64719f
C65 VN.n16 VSUBS 0.336386f
C66 VN.n17 VSUBS 0.07808f
C67 VN.n18 VSUBS 0.245365f
C68 VN.n19 VSUBS 0.057645f
C69 VN.n20 VSUBS 0.057645f
C70 VN.n21 VSUBS 0.07808f
C71 VN.n22 VSUBS 0.286272f
C72 VN.n23 VSUBS 0.077849f
C73 VN.t4 VSUBS 0.734086f
C74 VN.n24 VSUBS 0.37385f
C75 VN.n25 VSUBS 2.03498f
C76 B.n0 VSUBS 0.006213f
C77 B.n1 VSUBS 0.006213f
C78 B.n2 VSUBS 0.009189f
C79 B.n3 VSUBS 0.007042f
C80 B.n4 VSUBS 0.007042f
C81 B.n5 VSUBS 0.007042f
C82 B.n6 VSUBS 0.007042f
C83 B.n7 VSUBS 0.007042f
C84 B.n8 VSUBS 0.007042f
C85 B.n9 VSUBS 0.007042f
C86 B.n10 VSUBS 0.007042f
C87 B.n11 VSUBS 0.007042f
C88 B.n12 VSUBS 0.007042f
C89 B.n13 VSUBS 0.007042f
C90 B.n14 VSUBS 0.007042f
C91 B.n15 VSUBS 0.016049f
C92 B.n16 VSUBS 0.007042f
C93 B.n17 VSUBS 0.007042f
C94 B.n18 VSUBS 0.007042f
C95 B.n19 VSUBS 0.007042f
C96 B.n20 VSUBS 0.007042f
C97 B.n21 VSUBS 0.007042f
C98 B.n22 VSUBS 0.007042f
C99 B.n23 VSUBS 0.007042f
C100 B.n24 VSUBS 0.007042f
C101 B.n25 VSUBS 0.007042f
C102 B.t10 VSUBS 0.118469f
C103 B.t11 VSUBS 0.12756f
C104 B.t9 VSUBS 0.19847f
C105 B.n26 VSUBS 0.081232f
C106 B.n27 VSUBS 0.063294f
C107 B.n28 VSUBS 0.007042f
C108 B.n29 VSUBS 0.007042f
C109 B.n30 VSUBS 0.007042f
C110 B.n31 VSUBS 0.007042f
C111 B.t4 VSUBS 0.118469f
C112 B.t5 VSUBS 0.127559f
C113 B.t3 VSUBS 0.19847f
C114 B.n32 VSUBS 0.081232f
C115 B.n33 VSUBS 0.063294f
C116 B.n34 VSUBS 0.016315f
C117 B.n35 VSUBS 0.007042f
C118 B.n36 VSUBS 0.007042f
C119 B.n37 VSUBS 0.007042f
C120 B.n38 VSUBS 0.007042f
C121 B.n39 VSUBS 0.007042f
C122 B.n40 VSUBS 0.007042f
C123 B.n41 VSUBS 0.007042f
C124 B.n42 VSUBS 0.007042f
C125 B.n43 VSUBS 0.007042f
C126 B.n44 VSUBS 0.016049f
C127 B.n45 VSUBS 0.007042f
C128 B.n46 VSUBS 0.007042f
C129 B.n47 VSUBS 0.007042f
C130 B.n48 VSUBS 0.007042f
C131 B.n49 VSUBS 0.007042f
C132 B.n50 VSUBS 0.007042f
C133 B.n51 VSUBS 0.007042f
C134 B.n52 VSUBS 0.007042f
C135 B.n53 VSUBS 0.007042f
C136 B.n54 VSUBS 0.007042f
C137 B.n55 VSUBS 0.007042f
C138 B.n56 VSUBS 0.007042f
C139 B.n57 VSUBS 0.007042f
C140 B.n58 VSUBS 0.007042f
C141 B.n59 VSUBS 0.007042f
C142 B.n60 VSUBS 0.007042f
C143 B.n61 VSUBS 0.007042f
C144 B.n62 VSUBS 0.007042f
C145 B.n63 VSUBS 0.007042f
C146 B.n64 VSUBS 0.007042f
C147 B.n65 VSUBS 0.007042f
C148 B.n66 VSUBS 0.007042f
C149 B.n67 VSUBS 0.007042f
C150 B.n68 VSUBS 0.007042f
C151 B.n69 VSUBS 0.007042f
C152 B.n70 VSUBS 0.007042f
C153 B.n71 VSUBS 0.007042f
C154 B.n72 VSUBS 0.016049f
C155 B.n73 VSUBS 0.007042f
C156 B.n74 VSUBS 0.007042f
C157 B.n75 VSUBS 0.007042f
C158 B.n76 VSUBS 0.007042f
C159 B.n77 VSUBS 0.007042f
C160 B.n78 VSUBS 0.007042f
C161 B.n79 VSUBS 0.007042f
C162 B.n80 VSUBS 0.007042f
C163 B.n81 VSUBS 0.007042f
C164 B.t8 VSUBS 0.118469f
C165 B.t7 VSUBS 0.127559f
C166 B.t6 VSUBS 0.19847f
C167 B.n82 VSUBS 0.081232f
C168 B.n83 VSUBS 0.063294f
C169 B.n84 VSUBS 0.007042f
C170 B.n85 VSUBS 0.007042f
C171 B.n86 VSUBS 0.007042f
C172 B.n87 VSUBS 0.007042f
C173 B.n88 VSUBS 0.003935f
C174 B.n89 VSUBS 0.007042f
C175 B.n90 VSUBS 0.007042f
C176 B.n91 VSUBS 0.007042f
C177 B.n92 VSUBS 0.007042f
C178 B.n93 VSUBS 0.007042f
C179 B.n94 VSUBS 0.007042f
C180 B.n95 VSUBS 0.007042f
C181 B.n96 VSUBS 0.007042f
C182 B.n97 VSUBS 0.007042f
C183 B.n98 VSUBS 0.016049f
C184 B.n99 VSUBS 0.007042f
C185 B.n100 VSUBS 0.007042f
C186 B.n101 VSUBS 0.007042f
C187 B.n102 VSUBS 0.007042f
C188 B.n103 VSUBS 0.007042f
C189 B.n104 VSUBS 0.007042f
C190 B.n105 VSUBS 0.007042f
C191 B.n106 VSUBS 0.007042f
C192 B.n107 VSUBS 0.007042f
C193 B.n108 VSUBS 0.007042f
C194 B.n109 VSUBS 0.007042f
C195 B.n110 VSUBS 0.007042f
C196 B.n111 VSUBS 0.007042f
C197 B.n112 VSUBS 0.007042f
C198 B.n113 VSUBS 0.007042f
C199 B.n114 VSUBS 0.007042f
C200 B.n115 VSUBS 0.007042f
C201 B.n116 VSUBS 0.007042f
C202 B.n117 VSUBS 0.007042f
C203 B.n118 VSUBS 0.007042f
C204 B.n119 VSUBS 0.007042f
C205 B.n120 VSUBS 0.007042f
C206 B.n121 VSUBS 0.007042f
C207 B.n122 VSUBS 0.007042f
C208 B.n123 VSUBS 0.007042f
C209 B.n124 VSUBS 0.007042f
C210 B.n125 VSUBS 0.007042f
C211 B.n126 VSUBS 0.007042f
C212 B.n127 VSUBS 0.007042f
C213 B.n128 VSUBS 0.007042f
C214 B.n129 VSUBS 0.007042f
C215 B.n130 VSUBS 0.007042f
C216 B.n131 VSUBS 0.007042f
C217 B.n132 VSUBS 0.007042f
C218 B.n133 VSUBS 0.007042f
C219 B.n134 VSUBS 0.007042f
C220 B.n135 VSUBS 0.007042f
C221 B.n136 VSUBS 0.007042f
C222 B.n137 VSUBS 0.007042f
C223 B.n138 VSUBS 0.007042f
C224 B.n139 VSUBS 0.007042f
C225 B.n140 VSUBS 0.007042f
C226 B.n141 VSUBS 0.007042f
C227 B.n142 VSUBS 0.007042f
C228 B.n143 VSUBS 0.007042f
C229 B.n144 VSUBS 0.007042f
C230 B.n145 VSUBS 0.007042f
C231 B.n146 VSUBS 0.007042f
C232 B.n147 VSUBS 0.007042f
C233 B.n148 VSUBS 0.007042f
C234 B.n149 VSUBS 0.016049f
C235 B.n150 VSUBS 0.016882f
C236 B.n151 VSUBS 0.016882f
C237 B.n152 VSUBS 0.007042f
C238 B.n153 VSUBS 0.007042f
C239 B.n154 VSUBS 0.007042f
C240 B.n155 VSUBS 0.007042f
C241 B.n156 VSUBS 0.007042f
C242 B.n157 VSUBS 0.007042f
C243 B.n158 VSUBS 0.007042f
C244 B.n159 VSUBS 0.007042f
C245 B.n160 VSUBS 0.007042f
C246 B.n161 VSUBS 0.007042f
C247 B.n162 VSUBS 0.007042f
C248 B.n163 VSUBS 0.007042f
C249 B.n164 VSUBS 0.007042f
C250 B.n165 VSUBS 0.007042f
C251 B.n166 VSUBS 0.007042f
C252 B.n167 VSUBS 0.007042f
C253 B.n168 VSUBS 0.007042f
C254 B.n169 VSUBS 0.007042f
C255 B.n170 VSUBS 0.007042f
C256 B.n171 VSUBS 0.007042f
C257 B.n172 VSUBS 0.007042f
C258 B.n173 VSUBS 0.007042f
C259 B.n174 VSUBS 0.007042f
C260 B.n175 VSUBS 0.007042f
C261 B.n176 VSUBS 0.007042f
C262 B.t2 VSUBS 0.118469f
C263 B.t1 VSUBS 0.12756f
C264 B.t0 VSUBS 0.19847f
C265 B.n177 VSUBS 0.081232f
C266 B.n178 VSUBS 0.063294f
C267 B.n179 VSUBS 0.016315f
C268 B.n180 VSUBS 0.006627f
C269 B.n181 VSUBS 0.007042f
C270 B.n182 VSUBS 0.007042f
C271 B.n183 VSUBS 0.007042f
C272 B.n184 VSUBS 0.007042f
C273 B.n185 VSUBS 0.007042f
C274 B.n186 VSUBS 0.007042f
C275 B.n187 VSUBS 0.007042f
C276 B.n188 VSUBS 0.007042f
C277 B.n189 VSUBS 0.007042f
C278 B.n190 VSUBS 0.007042f
C279 B.n191 VSUBS 0.007042f
C280 B.n192 VSUBS 0.007042f
C281 B.n193 VSUBS 0.007042f
C282 B.n194 VSUBS 0.007042f
C283 B.n195 VSUBS 0.007042f
C284 B.n196 VSUBS 0.003935f
C285 B.n197 VSUBS 0.016315f
C286 B.n198 VSUBS 0.006627f
C287 B.n199 VSUBS 0.007042f
C288 B.n200 VSUBS 0.007042f
C289 B.n201 VSUBS 0.007042f
C290 B.n202 VSUBS 0.007042f
C291 B.n203 VSUBS 0.007042f
C292 B.n204 VSUBS 0.007042f
C293 B.n205 VSUBS 0.007042f
C294 B.n206 VSUBS 0.007042f
C295 B.n207 VSUBS 0.007042f
C296 B.n208 VSUBS 0.007042f
C297 B.n209 VSUBS 0.007042f
C298 B.n210 VSUBS 0.007042f
C299 B.n211 VSUBS 0.007042f
C300 B.n212 VSUBS 0.007042f
C301 B.n213 VSUBS 0.007042f
C302 B.n214 VSUBS 0.007042f
C303 B.n215 VSUBS 0.007042f
C304 B.n216 VSUBS 0.007042f
C305 B.n217 VSUBS 0.007042f
C306 B.n218 VSUBS 0.007042f
C307 B.n219 VSUBS 0.007042f
C308 B.n220 VSUBS 0.007042f
C309 B.n221 VSUBS 0.007042f
C310 B.n222 VSUBS 0.007042f
C311 B.n223 VSUBS 0.007042f
C312 B.n224 VSUBS 0.007042f
C313 B.n225 VSUBS 0.016882f
C314 B.n226 VSUBS 0.016049f
C315 B.n227 VSUBS 0.016882f
C316 B.n228 VSUBS 0.007042f
C317 B.n229 VSUBS 0.007042f
C318 B.n230 VSUBS 0.007042f
C319 B.n231 VSUBS 0.007042f
C320 B.n232 VSUBS 0.007042f
C321 B.n233 VSUBS 0.007042f
C322 B.n234 VSUBS 0.007042f
C323 B.n235 VSUBS 0.007042f
C324 B.n236 VSUBS 0.007042f
C325 B.n237 VSUBS 0.007042f
C326 B.n238 VSUBS 0.007042f
C327 B.n239 VSUBS 0.007042f
C328 B.n240 VSUBS 0.007042f
C329 B.n241 VSUBS 0.007042f
C330 B.n242 VSUBS 0.007042f
C331 B.n243 VSUBS 0.007042f
C332 B.n244 VSUBS 0.007042f
C333 B.n245 VSUBS 0.007042f
C334 B.n246 VSUBS 0.007042f
C335 B.n247 VSUBS 0.007042f
C336 B.n248 VSUBS 0.007042f
C337 B.n249 VSUBS 0.007042f
C338 B.n250 VSUBS 0.007042f
C339 B.n251 VSUBS 0.007042f
C340 B.n252 VSUBS 0.007042f
C341 B.n253 VSUBS 0.007042f
C342 B.n254 VSUBS 0.007042f
C343 B.n255 VSUBS 0.007042f
C344 B.n256 VSUBS 0.007042f
C345 B.n257 VSUBS 0.007042f
C346 B.n258 VSUBS 0.007042f
C347 B.n259 VSUBS 0.007042f
C348 B.n260 VSUBS 0.007042f
C349 B.n261 VSUBS 0.007042f
C350 B.n262 VSUBS 0.007042f
C351 B.n263 VSUBS 0.007042f
C352 B.n264 VSUBS 0.007042f
C353 B.n265 VSUBS 0.007042f
C354 B.n266 VSUBS 0.007042f
C355 B.n267 VSUBS 0.007042f
C356 B.n268 VSUBS 0.007042f
C357 B.n269 VSUBS 0.007042f
C358 B.n270 VSUBS 0.007042f
C359 B.n271 VSUBS 0.007042f
C360 B.n272 VSUBS 0.007042f
C361 B.n273 VSUBS 0.007042f
C362 B.n274 VSUBS 0.007042f
C363 B.n275 VSUBS 0.007042f
C364 B.n276 VSUBS 0.007042f
C365 B.n277 VSUBS 0.007042f
C366 B.n278 VSUBS 0.007042f
C367 B.n279 VSUBS 0.007042f
C368 B.n280 VSUBS 0.007042f
C369 B.n281 VSUBS 0.007042f
C370 B.n282 VSUBS 0.007042f
C371 B.n283 VSUBS 0.007042f
C372 B.n284 VSUBS 0.007042f
C373 B.n285 VSUBS 0.007042f
C374 B.n286 VSUBS 0.007042f
C375 B.n287 VSUBS 0.007042f
C376 B.n288 VSUBS 0.007042f
C377 B.n289 VSUBS 0.007042f
C378 B.n290 VSUBS 0.007042f
C379 B.n291 VSUBS 0.007042f
C380 B.n292 VSUBS 0.007042f
C381 B.n293 VSUBS 0.007042f
C382 B.n294 VSUBS 0.007042f
C383 B.n295 VSUBS 0.007042f
C384 B.n296 VSUBS 0.007042f
C385 B.n297 VSUBS 0.007042f
C386 B.n298 VSUBS 0.007042f
C387 B.n299 VSUBS 0.007042f
C388 B.n300 VSUBS 0.007042f
C389 B.n301 VSUBS 0.007042f
C390 B.n302 VSUBS 0.007042f
C391 B.n303 VSUBS 0.007042f
C392 B.n304 VSUBS 0.007042f
C393 B.n305 VSUBS 0.007042f
C394 B.n306 VSUBS 0.007042f
C395 B.n307 VSUBS 0.007042f
C396 B.n308 VSUBS 0.007042f
C397 B.n309 VSUBS 0.016049f
C398 B.n310 VSUBS 0.016882f
C399 B.n311 VSUBS 0.016882f
C400 B.n312 VSUBS 0.007042f
C401 B.n313 VSUBS 0.007042f
C402 B.n314 VSUBS 0.007042f
C403 B.n315 VSUBS 0.007042f
C404 B.n316 VSUBS 0.007042f
C405 B.n317 VSUBS 0.007042f
C406 B.n318 VSUBS 0.007042f
C407 B.n319 VSUBS 0.007042f
C408 B.n320 VSUBS 0.007042f
C409 B.n321 VSUBS 0.007042f
C410 B.n322 VSUBS 0.007042f
C411 B.n323 VSUBS 0.007042f
C412 B.n324 VSUBS 0.007042f
C413 B.n325 VSUBS 0.007042f
C414 B.n326 VSUBS 0.007042f
C415 B.n327 VSUBS 0.007042f
C416 B.n328 VSUBS 0.007042f
C417 B.n329 VSUBS 0.007042f
C418 B.n330 VSUBS 0.007042f
C419 B.n331 VSUBS 0.007042f
C420 B.n332 VSUBS 0.007042f
C421 B.n333 VSUBS 0.007042f
C422 B.n334 VSUBS 0.007042f
C423 B.n335 VSUBS 0.007042f
C424 B.n336 VSUBS 0.007042f
C425 B.n337 VSUBS 0.006627f
C426 B.n338 VSUBS 0.007042f
C427 B.n339 VSUBS 0.007042f
C428 B.n340 VSUBS 0.003935f
C429 B.n341 VSUBS 0.007042f
C430 B.n342 VSUBS 0.007042f
C431 B.n343 VSUBS 0.007042f
C432 B.n344 VSUBS 0.007042f
C433 B.n345 VSUBS 0.007042f
C434 B.n346 VSUBS 0.007042f
C435 B.n347 VSUBS 0.007042f
C436 B.n348 VSUBS 0.007042f
C437 B.n349 VSUBS 0.007042f
C438 B.n350 VSUBS 0.007042f
C439 B.n351 VSUBS 0.007042f
C440 B.n352 VSUBS 0.007042f
C441 B.n353 VSUBS 0.003935f
C442 B.n354 VSUBS 0.016315f
C443 B.n355 VSUBS 0.006627f
C444 B.n356 VSUBS 0.007042f
C445 B.n357 VSUBS 0.007042f
C446 B.n358 VSUBS 0.007042f
C447 B.n359 VSUBS 0.007042f
C448 B.n360 VSUBS 0.007042f
C449 B.n361 VSUBS 0.007042f
C450 B.n362 VSUBS 0.007042f
C451 B.n363 VSUBS 0.007042f
C452 B.n364 VSUBS 0.007042f
C453 B.n365 VSUBS 0.007042f
C454 B.n366 VSUBS 0.007042f
C455 B.n367 VSUBS 0.007042f
C456 B.n368 VSUBS 0.007042f
C457 B.n369 VSUBS 0.007042f
C458 B.n370 VSUBS 0.007042f
C459 B.n371 VSUBS 0.007042f
C460 B.n372 VSUBS 0.007042f
C461 B.n373 VSUBS 0.007042f
C462 B.n374 VSUBS 0.007042f
C463 B.n375 VSUBS 0.007042f
C464 B.n376 VSUBS 0.007042f
C465 B.n377 VSUBS 0.007042f
C466 B.n378 VSUBS 0.007042f
C467 B.n379 VSUBS 0.007042f
C468 B.n380 VSUBS 0.007042f
C469 B.n381 VSUBS 0.007042f
C470 B.n382 VSUBS 0.016882f
C471 B.n383 VSUBS 0.016882f
C472 B.n384 VSUBS 0.016049f
C473 B.n385 VSUBS 0.007042f
C474 B.n386 VSUBS 0.007042f
C475 B.n387 VSUBS 0.007042f
C476 B.n388 VSUBS 0.007042f
C477 B.n389 VSUBS 0.007042f
C478 B.n390 VSUBS 0.007042f
C479 B.n391 VSUBS 0.007042f
C480 B.n392 VSUBS 0.007042f
C481 B.n393 VSUBS 0.007042f
C482 B.n394 VSUBS 0.007042f
C483 B.n395 VSUBS 0.007042f
C484 B.n396 VSUBS 0.007042f
C485 B.n397 VSUBS 0.007042f
C486 B.n398 VSUBS 0.007042f
C487 B.n399 VSUBS 0.007042f
C488 B.n400 VSUBS 0.007042f
C489 B.n401 VSUBS 0.007042f
C490 B.n402 VSUBS 0.007042f
C491 B.n403 VSUBS 0.007042f
C492 B.n404 VSUBS 0.007042f
C493 B.n405 VSUBS 0.007042f
C494 B.n406 VSUBS 0.007042f
C495 B.n407 VSUBS 0.007042f
C496 B.n408 VSUBS 0.007042f
C497 B.n409 VSUBS 0.007042f
C498 B.n410 VSUBS 0.007042f
C499 B.n411 VSUBS 0.007042f
C500 B.n412 VSUBS 0.007042f
C501 B.n413 VSUBS 0.007042f
C502 B.n414 VSUBS 0.007042f
C503 B.n415 VSUBS 0.007042f
C504 B.n416 VSUBS 0.007042f
C505 B.n417 VSUBS 0.007042f
C506 B.n418 VSUBS 0.007042f
C507 B.n419 VSUBS 0.007042f
C508 B.n420 VSUBS 0.007042f
C509 B.n421 VSUBS 0.007042f
C510 B.n422 VSUBS 0.007042f
C511 B.n423 VSUBS 0.009189f
C512 B.n424 VSUBS 0.009789f
C513 B.n425 VSUBS 0.019466f
C514 VTAIL.t3 VSUBS 0.090635f
C515 VTAIL.t5 VSUBS 0.090635f
C516 VTAIL.n0 VSUBS 0.480809f
C517 VTAIL.n1 VSUBS 0.513562f
C518 VTAIL.t0 VSUBS 0.681903f
C519 VTAIL.n2 VSUBS 0.594387f
C520 VTAIL.t10 VSUBS 0.681903f
C521 VTAIL.n3 VSUBS 0.594387f
C522 VTAIL.t8 VSUBS 0.090635f
C523 VTAIL.t15 VSUBS 0.090635f
C524 VTAIL.n4 VSUBS 0.480809f
C525 VTAIL.n5 VSUBS 0.604667f
C526 VTAIL.t12 VSUBS 0.681903f
C527 VTAIL.n6 VSUBS 1.32506f
C528 VTAIL.t1 VSUBS 0.681905f
C529 VTAIL.n7 VSUBS 1.32506f
C530 VTAIL.t4 VSUBS 0.090635f
C531 VTAIL.t2 VSUBS 0.090635f
C532 VTAIL.n8 VSUBS 0.480812f
C533 VTAIL.n9 VSUBS 0.604665f
C534 VTAIL.t6 VSUBS 0.681905f
C535 VTAIL.n10 VSUBS 0.594385f
C536 VTAIL.t13 VSUBS 0.681905f
C537 VTAIL.n11 VSUBS 0.594385f
C538 VTAIL.t14 VSUBS 0.090635f
C539 VTAIL.t9 VSUBS 0.090635f
C540 VTAIL.n12 VSUBS 0.480812f
C541 VTAIL.n13 VSUBS 0.604665f
C542 VTAIL.t11 VSUBS 0.681903f
C543 VTAIL.n14 VSUBS 1.32506f
C544 VTAIL.t7 VSUBS 0.681903f
C545 VTAIL.n15 VSUBS 1.32015f
C546 VDD1.t4 VSUBS 0.088465f
C547 VDD1.t2 VSUBS 0.088465f
C548 VDD1.n0 VSUBS 0.536743f
C549 VDD1.t5 VSUBS 0.088465f
C550 VDD1.t1 VSUBS 0.088465f
C551 VDD1.n1 VSUBS 0.536173f
C552 VDD1.t3 VSUBS 0.088465f
C553 VDD1.t0 VSUBS 0.088465f
C554 VDD1.n2 VSUBS 0.536173f
C555 VDD1.n3 VSUBS 2.3088f
C556 VDD1.t7 VSUBS 0.088465f
C557 VDD1.t6 VSUBS 0.088465f
C558 VDD1.n4 VSUBS 0.533794f
C559 VDD1.n5 VSUBS 2.02116f
C560 VP.n0 VSUBS 0.079597f
C561 VP.t0 VSUBS 0.669718f
C562 VP.n1 VSUBS 0.048178f
C563 VP.n2 VSUBS 0.079597f
C564 VP.t7 VSUBS 0.669718f
C565 VP.n3 VSUBS 0.079597f
C566 VP.t4 VSUBS 0.759639f
C567 VP.t6 VSUBS 0.669718f
C568 VP.n4 VSUBS 0.048178f
C569 VP.t2 VSUBS 0.795984f
C570 VP.n5 VSUBS 0.380467f
C571 VP.t1 VSUBS 0.669718f
C572 VP.n6 VSUBS 0.348095f
C573 VP.n7 VSUBS 0.080798f
C574 VP.n8 VSUBS 0.253907f
C575 VP.n9 VSUBS 0.059651f
C576 VP.n10 VSUBS 0.059651f
C577 VP.n11 VSUBS 0.080798f
C578 VP.n12 VSUBS 0.296237f
C579 VP.n13 VSUBS 0.080559f
C580 VP.n14 VSUBS 0.386864f
C581 VP.n15 VSUBS 2.07169f
C582 VP.n16 VSUBS 2.12859f
C583 VP.t3 VSUBS 0.759639f
C584 VP.n17 VSUBS 0.386864f
C585 VP.n18 VSUBS 0.080559f
C586 VP.n19 VSUBS 0.296237f
C587 VP.n20 VSUBS 0.080798f
C588 VP.n21 VSUBS 0.059651f
C589 VP.n22 VSUBS 0.059651f
C590 VP.n23 VSUBS 0.059651f
C591 VP.n24 VSUBS 0.080798f
C592 VP.n25 VSUBS 0.296237f
C593 VP.n26 VSUBS 0.080559f
C594 VP.t5 VSUBS 0.759639f
C595 VP.n27 VSUBS 0.386864f
C596 VP.n28 VSUBS 0.055866f
.ends

