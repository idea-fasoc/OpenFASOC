* NGSPICE file created from diff_pair_sample_0666.ext - technology: sky130A

.subckt diff_pair_sample_0666 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t18 VP.t0 VDD1.t0 B.t2 sky130_fd_pr__nfet_01v8 ad=0.28545 pd=2.06 as=0.28545 ps=2.06 w=1.73 l=0.83
X1 VDD1.t2 VP.t1 VTAIL.t17 B.t23 sky130_fd_pr__nfet_01v8 ad=0.6747 pd=4.24 as=0.28545 ps=2.06 w=1.73 l=0.83
X2 VDD1.t9 VP.t2 VTAIL.t16 B.t4 sky130_fd_pr__nfet_01v8 ad=0.28545 pd=2.06 as=0.28545 ps=2.06 w=1.73 l=0.83
X3 VDD1.t8 VP.t3 VTAIL.t15 B.t3 sky130_fd_pr__nfet_01v8 ad=0.28545 pd=2.06 as=0.6747 ps=4.24 w=1.73 l=0.83
X4 VDD1.t7 VP.t4 VTAIL.t14 B.t8 sky130_fd_pr__nfet_01v8 ad=0.28545 pd=2.06 as=0.6747 ps=4.24 w=1.73 l=0.83
X5 VTAIL.t13 VP.t5 VDD1.t4 B.t7 sky130_fd_pr__nfet_01v8 ad=0.28545 pd=2.06 as=0.28545 ps=2.06 w=1.73 l=0.83
X6 VTAIL.t12 VP.t6 VDD1.t3 B.t0 sky130_fd_pr__nfet_01v8 ad=0.28545 pd=2.06 as=0.28545 ps=2.06 w=1.73 l=0.83
X7 VTAIL.t11 VP.t7 VDD1.t1 B.t6 sky130_fd_pr__nfet_01v8 ad=0.28545 pd=2.06 as=0.28545 ps=2.06 w=1.73 l=0.83
X8 VDD2.t9 VN.t0 VTAIL.t19 B.t23 sky130_fd_pr__nfet_01v8 ad=0.6747 pd=4.24 as=0.28545 ps=2.06 w=1.73 l=0.83
X9 B.t22 B.t20 B.t21 B.t17 sky130_fd_pr__nfet_01v8 ad=0.6747 pd=4.24 as=0 ps=0 w=1.73 l=0.83
X10 VDD1.t6 VP.t8 VTAIL.t10 B.t5 sky130_fd_pr__nfet_01v8 ad=0.6747 pd=4.24 as=0.28545 ps=2.06 w=1.73 l=0.83
X11 VTAIL.t2 VN.t1 VDD2.t8 B.t2 sky130_fd_pr__nfet_01v8 ad=0.28545 pd=2.06 as=0.28545 ps=2.06 w=1.73 l=0.83
X12 VTAIL.t6 VN.t2 VDD2.t7 B.t6 sky130_fd_pr__nfet_01v8 ad=0.28545 pd=2.06 as=0.28545 ps=2.06 w=1.73 l=0.83
X13 B.t19 B.t16 B.t18 B.t17 sky130_fd_pr__nfet_01v8 ad=0.6747 pd=4.24 as=0 ps=0 w=1.73 l=0.83
X14 VDD2.t6 VN.t3 VTAIL.t8 B.t8 sky130_fd_pr__nfet_01v8 ad=0.28545 pd=2.06 as=0.6747 ps=4.24 w=1.73 l=0.83
X15 B.t15 B.t13 B.t14 B.t10 sky130_fd_pr__nfet_01v8 ad=0.6747 pd=4.24 as=0 ps=0 w=1.73 l=0.83
X16 B.t12 B.t9 B.t11 B.t10 sky130_fd_pr__nfet_01v8 ad=0.6747 pd=4.24 as=0 ps=0 w=1.73 l=0.83
X17 VTAIL.t7 VN.t4 VDD2.t5 B.t7 sky130_fd_pr__nfet_01v8 ad=0.28545 pd=2.06 as=0.28545 ps=2.06 w=1.73 l=0.83
X18 VDD2.t4 VN.t5 VTAIL.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=0.28545 pd=2.06 as=0.28545 ps=2.06 w=1.73 l=0.83
X19 VTAIL.t0 VN.t6 VDD2.t3 B.t0 sky130_fd_pr__nfet_01v8 ad=0.28545 pd=2.06 as=0.28545 ps=2.06 w=1.73 l=0.83
X20 VDD2.t2 VN.t7 VTAIL.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=0.6747 pd=4.24 as=0.28545 ps=2.06 w=1.73 l=0.83
X21 VDD2.t1 VN.t8 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=0.28545 pd=2.06 as=0.28545 ps=2.06 w=1.73 l=0.83
X22 VDD2.t0 VN.t9 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=0.28545 pd=2.06 as=0.6747 ps=4.24 w=1.73 l=0.83
X23 VDD1.t5 VP.t9 VTAIL.t9 B.t1 sky130_fd_pr__nfet_01v8 ad=0.28545 pd=2.06 as=0.28545 ps=2.06 w=1.73 l=0.83
R0 VP.n40 VP.n39 161.3
R1 VP.n11 VP.n8 161.3
R2 VP.n13 VP.n12 161.3
R3 VP.n15 VP.n7 161.3
R4 VP.n17 VP.n16 161.3
R5 VP.n19 VP.n18 161.3
R6 VP.n20 VP.n5 161.3
R7 VP.n22 VP.n21 161.3
R8 VP.n38 VP.n0 161.3
R9 VP.n37 VP.n36 161.3
R10 VP.n35 VP.n34 161.3
R11 VP.n33 VP.n2 161.3
R12 VP.n31 VP.n30 161.3
R13 VP.n29 VP.n3 161.3
R14 VP.n28 VP.n27 161.3
R15 VP.n25 VP.n4 161.3
R16 VP.n24 VP.n23 161.3
R17 VP.n10 VP.t1 122.052
R18 VP.n24 VP.t8 97.8523
R19 VP.n39 VP.t4 97.8523
R20 VP.n21 VP.t3 97.8523
R21 VP.n31 VP.n3 56.5193
R22 VP.n34 VP.n33 56.5193
R23 VP.n16 VP.n15 56.5193
R24 VP.n13 VP.n8 56.5193
R25 VP.n26 VP.t6 50.233
R26 VP.n32 VP.t2 50.233
R27 VP.n1 VP.t7 50.233
R28 VP.n6 VP.t5 50.233
R29 VP.n14 VP.t9 50.233
R30 VP.n9 VP.t0 50.233
R31 VP.n11 VP.n10 42.3937
R32 VP.n27 VP.n25 41.4647
R33 VP.n38 VP.n37 41.4647
R34 VP.n20 VP.n19 41.4647
R35 VP.n23 VP.n22 35.7505
R36 VP.n10 VP.n9 33.4547
R37 VP.n25 VP.n24 22.6399
R38 VP.n39 VP.n38 22.6399
R39 VP.n21 VP.n20 22.6399
R40 VP.n26 VP.n3 20.0634
R41 VP.n34 VP.n1 20.0634
R42 VP.n16 VP.n6 20.0634
R43 VP.n9 VP.n8 20.0634
R44 VP.n32 VP.n31 12.234
R45 VP.n33 VP.n32 12.234
R46 VP.n14 VP.n13 12.234
R47 VP.n15 VP.n14 12.234
R48 VP.n27 VP.n26 4.40456
R49 VP.n37 VP.n1 4.40456
R50 VP.n19 VP.n6 4.40456
R51 VP.n12 VP.n11 0.189894
R52 VP.n12 VP.n7 0.189894
R53 VP.n17 VP.n7 0.189894
R54 VP.n18 VP.n17 0.189894
R55 VP.n18 VP.n5 0.189894
R56 VP.n22 VP.n5 0.189894
R57 VP.n23 VP.n4 0.189894
R58 VP.n28 VP.n4 0.189894
R59 VP.n29 VP.n28 0.189894
R60 VP.n30 VP.n29 0.189894
R61 VP.n30 VP.n2 0.189894
R62 VP.n35 VP.n2 0.189894
R63 VP.n36 VP.n35 0.189894
R64 VP.n36 VP.n0 0.189894
R65 VP.n40 VP.n0 0.189894
R66 VP VP.n40 0.0516364
R67 VDD1.n2 VDD1.n0 289.615
R68 VDD1.n11 VDD1.n9 289.615
R69 VDD1.n3 VDD1.n2 185
R70 VDD1.n12 VDD1.n11 185
R71 VDD1.t2 VDD1.n1 164.876
R72 VDD1.t6 VDD1.n10 164.876
R73 VDD1.n19 VDD1.n18 101.147
R74 VDD1.n21 VDD1.n20 100.454
R75 VDD1.n8 VDD1.n7 100.454
R76 VDD1.n17 VDD1.n16 100.454
R77 VDD1.n2 VDD1.t2 52.3082
R78 VDD1.n11 VDD1.t6 52.3082
R79 VDD1.n8 VDD1.n6 50.8338
R80 VDD1.n17 VDD1.n15 50.8338
R81 VDD1.n21 VDD1.n19 31.0397
R82 VDD1.n3 VDD1.n1 14.7318
R83 VDD1.n12 VDD1.n10 14.7318
R84 VDD1.n4 VDD1.n0 12.8005
R85 VDD1.n13 VDD1.n9 12.8005
R86 VDD1.n20 VDD1.t4 11.4456
R87 VDD1.n20 VDD1.t8 11.4456
R88 VDD1.n7 VDD1.t0 11.4456
R89 VDD1.n7 VDD1.t5 11.4456
R90 VDD1.n18 VDD1.t1 11.4456
R91 VDD1.n18 VDD1.t7 11.4456
R92 VDD1.n16 VDD1.t3 11.4456
R93 VDD1.n16 VDD1.t9 11.4456
R94 VDD1.n6 VDD1.n5 9.45567
R95 VDD1.n15 VDD1.n14 9.45567
R96 VDD1.n5 VDD1.n4 9.3005
R97 VDD1.n14 VDD1.n13 9.3005
R98 VDD1.n5 VDD1.n1 5.62509
R99 VDD1.n14 VDD1.n10 5.62509
R100 VDD1.n6 VDD1.n0 1.16414
R101 VDD1.n15 VDD1.n9 1.16414
R102 VDD1 VDD1.n21 0.69231
R103 VDD1.n4 VDD1.n3 0.388379
R104 VDD1.n13 VDD1.n12 0.388379
R105 VDD1 VDD1.n8 0.30869
R106 VDD1.n19 VDD1.n17 0.195154
R107 VTAIL.n40 VTAIL.n38 289.615
R108 VTAIL.n4 VTAIL.n2 289.615
R109 VTAIL.n32 VTAIL.n30 289.615
R110 VTAIL.n20 VTAIL.n18 289.615
R111 VTAIL.n41 VTAIL.n40 185
R112 VTAIL.n5 VTAIL.n4 185
R113 VTAIL.n33 VTAIL.n32 185
R114 VTAIL.n21 VTAIL.n20 185
R115 VTAIL.t3 VTAIL.n39 164.876
R116 VTAIL.t14 VTAIL.n3 164.876
R117 VTAIL.t15 VTAIL.n31 164.876
R118 VTAIL.t8 VTAIL.n19 164.876
R119 VTAIL.n29 VTAIL.n28 83.7746
R120 VTAIL.n27 VTAIL.n26 83.7746
R121 VTAIL.n17 VTAIL.n16 83.7746
R122 VTAIL.n15 VTAIL.n14 83.7746
R123 VTAIL.n47 VTAIL.n46 83.7746
R124 VTAIL.n1 VTAIL.n0 83.7746
R125 VTAIL.n11 VTAIL.n10 83.7746
R126 VTAIL.n13 VTAIL.n12 83.7746
R127 VTAIL.n40 VTAIL.t3 52.3082
R128 VTAIL.n4 VTAIL.t14 52.3082
R129 VTAIL.n32 VTAIL.t15 52.3082
R130 VTAIL.n20 VTAIL.t8 52.3082
R131 VTAIL.n45 VTAIL.n44 33.155
R132 VTAIL.n9 VTAIL.n8 33.155
R133 VTAIL.n37 VTAIL.n36 33.155
R134 VTAIL.n25 VTAIL.n24 33.155
R135 VTAIL.n15 VTAIL.n13 15.8583
R136 VTAIL.n45 VTAIL.n37 14.8583
R137 VTAIL.n41 VTAIL.n39 14.7318
R138 VTAIL.n5 VTAIL.n3 14.7318
R139 VTAIL.n33 VTAIL.n31 14.7318
R140 VTAIL.n21 VTAIL.n19 14.7318
R141 VTAIL.n42 VTAIL.n38 12.8005
R142 VTAIL.n6 VTAIL.n2 12.8005
R143 VTAIL.n34 VTAIL.n30 12.8005
R144 VTAIL.n22 VTAIL.n18 12.8005
R145 VTAIL.n46 VTAIL.t1 11.4456
R146 VTAIL.n46 VTAIL.t7 11.4456
R147 VTAIL.n0 VTAIL.t19 11.4456
R148 VTAIL.n0 VTAIL.t2 11.4456
R149 VTAIL.n10 VTAIL.t16 11.4456
R150 VTAIL.n10 VTAIL.t11 11.4456
R151 VTAIL.n12 VTAIL.t10 11.4456
R152 VTAIL.n12 VTAIL.t12 11.4456
R153 VTAIL.n28 VTAIL.t9 11.4456
R154 VTAIL.n28 VTAIL.t13 11.4456
R155 VTAIL.n26 VTAIL.t17 11.4456
R156 VTAIL.n26 VTAIL.t18 11.4456
R157 VTAIL.n16 VTAIL.t4 11.4456
R158 VTAIL.n16 VTAIL.t6 11.4456
R159 VTAIL.n14 VTAIL.t5 11.4456
R160 VTAIL.n14 VTAIL.t0 11.4456
R161 VTAIL.n44 VTAIL.n43 9.45567
R162 VTAIL.n8 VTAIL.n7 9.45567
R163 VTAIL.n36 VTAIL.n35 9.45567
R164 VTAIL.n24 VTAIL.n23 9.45567
R165 VTAIL.n43 VTAIL.n42 9.3005
R166 VTAIL.n7 VTAIL.n6 9.3005
R167 VTAIL.n35 VTAIL.n34 9.3005
R168 VTAIL.n23 VTAIL.n22 9.3005
R169 VTAIL.n43 VTAIL.n39 5.62509
R170 VTAIL.n7 VTAIL.n3 5.62509
R171 VTAIL.n35 VTAIL.n31 5.62509
R172 VTAIL.n23 VTAIL.n19 5.62509
R173 VTAIL.n44 VTAIL.n38 1.16414
R174 VTAIL.n8 VTAIL.n2 1.16414
R175 VTAIL.n36 VTAIL.n30 1.16414
R176 VTAIL.n24 VTAIL.n18 1.16414
R177 VTAIL.n17 VTAIL.n15 1.0005
R178 VTAIL.n25 VTAIL.n17 1.0005
R179 VTAIL.n29 VTAIL.n27 1.0005
R180 VTAIL.n37 VTAIL.n29 1.0005
R181 VTAIL.n13 VTAIL.n11 1.0005
R182 VTAIL.n11 VTAIL.n9 1.0005
R183 VTAIL.n47 VTAIL.n45 1.0005
R184 VTAIL.n27 VTAIL.n25 0.970328
R185 VTAIL.n9 VTAIL.n1 0.970328
R186 VTAIL VTAIL.n1 0.80869
R187 VTAIL.n42 VTAIL.n41 0.388379
R188 VTAIL.n6 VTAIL.n5 0.388379
R189 VTAIL.n34 VTAIL.n33 0.388379
R190 VTAIL.n22 VTAIL.n21 0.388379
R191 VTAIL VTAIL.n47 0.19231
R192 B.n399 B.n398 585
R193 B.n136 B.n71 585
R194 B.n135 B.n134 585
R195 B.n133 B.n132 585
R196 B.n131 B.n130 585
R197 B.n129 B.n128 585
R198 B.n127 B.n126 585
R199 B.n125 B.n124 585
R200 B.n123 B.n122 585
R201 B.n121 B.n120 585
R202 B.n119 B.n118 585
R203 B.n116 B.n115 585
R204 B.n114 B.n113 585
R205 B.n112 B.n111 585
R206 B.n110 B.n109 585
R207 B.n108 B.n107 585
R208 B.n106 B.n105 585
R209 B.n104 B.n103 585
R210 B.n102 B.n101 585
R211 B.n100 B.n99 585
R212 B.n98 B.n97 585
R213 B.n95 B.n94 585
R214 B.n93 B.n92 585
R215 B.n91 B.n90 585
R216 B.n89 B.n88 585
R217 B.n87 B.n86 585
R218 B.n85 B.n84 585
R219 B.n83 B.n82 585
R220 B.n81 B.n80 585
R221 B.n79 B.n78 585
R222 B.n77 B.n76 585
R223 B.n54 B.n53 585
R224 B.n397 B.n55 585
R225 B.n402 B.n55 585
R226 B.n396 B.n395 585
R227 B.n395 B.n51 585
R228 B.n394 B.n50 585
R229 B.n408 B.n50 585
R230 B.n393 B.n49 585
R231 B.n409 B.n49 585
R232 B.n392 B.n48 585
R233 B.n410 B.n48 585
R234 B.n391 B.n390 585
R235 B.n390 B.n44 585
R236 B.n389 B.n43 585
R237 B.n416 B.n43 585
R238 B.n388 B.n42 585
R239 B.n417 B.n42 585
R240 B.n387 B.n41 585
R241 B.n418 B.n41 585
R242 B.n386 B.n385 585
R243 B.n385 B.n37 585
R244 B.n384 B.n36 585
R245 B.n424 B.n36 585
R246 B.n383 B.n35 585
R247 B.n425 B.n35 585
R248 B.n382 B.n34 585
R249 B.n426 B.n34 585
R250 B.n381 B.n380 585
R251 B.n380 B.n30 585
R252 B.n379 B.n29 585
R253 B.n432 B.n29 585
R254 B.n378 B.n28 585
R255 B.n433 B.n28 585
R256 B.n377 B.n27 585
R257 B.n434 B.n27 585
R258 B.n376 B.n375 585
R259 B.n375 B.n23 585
R260 B.n374 B.n22 585
R261 B.n440 B.n22 585
R262 B.n373 B.n21 585
R263 B.n441 B.n21 585
R264 B.n372 B.n20 585
R265 B.n442 B.n20 585
R266 B.n371 B.n370 585
R267 B.n370 B.n19 585
R268 B.n369 B.n15 585
R269 B.n448 B.n15 585
R270 B.n368 B.n14 585
R271 B.n449 B.n14 585
R272 B.n367 B.n13 585
R273 B.n450 B.n13 585
R274 B.n366 B.n365 585
R275 B.n365 B.n12 585
R276 B.n364 B.n363 585
R277 B.n364 B.n8 585
R278 B.n362 B.n7 585
R279 B.n457 B.n7 585
R280 B.n361 B.n6 585
R281 B.n458 B.n6 585
R282 B.n360 B.n5 585
R283 B.n459 B.n5 585
R284 B.n359 B.n358 585
R285 B.n358 B.n4 585
R286 B.n357 B.n137 585
R287 B.n357 B.n356 585
R288 B.n346 B.n138 585
R289 B.n349 B.n138 585
R290 B.n348 B.n347 585
R291 B.n350 B.n348 585
R292 B.n345 B.n143 585
R293 B.n143 B.n142 585
R294 B.n344 B.n343 585
R295 B.n343 B.n342 585
R296 B.n145 B.n144 585
R297 B.n335 B.n145 585
R298 B.n334 B.n333 585
R299 B.n336 B.n334 585
R300 B.n332 B.n150 585
R301 B.n150 B.n149 585
R302 B.n331 B.n330 585
R303 B.n330 B.n329 585
R304 B.n152 B.n151 585
R305 B.n153 B.n152 585
R306 B.n322 B.n321 585
R307 B.n323 B.n322 585
R308 B.n320 B.n158 585
R309 B.n158 B.n157 585
R310 B.n319 B.n318 585
R311 B.n318 B.n317 585
R312 B.n160 B.n159 585
R313 B.n161 B.n160 585
R314 B.n310 B.n309 585
R315 B.n311 B.n310 585
R316 B.n308 B.n165 585
R317 B.n169 B.n165 585
R318 B.n307 B.n306 585
R319 B.n306 B.n305 585
R320 B.n167 B.n166 585
R321 B.n168 B.n167 585
R322 B.n298 B.n297 585
R323 B.n299 B.n298 585
R324 B.n296 B.n174 585
R325 B.n174 B.n173 585
R326 B.n295 B.n294 585
R327 B.n294 B.n293 585
R328 B.n176 B.n175 585
R329 B.n177 B.n176 585
R330 B.n286 B.n285 585
R331 B.n287 B.n286 585
R332 B.n284 B.n182 585
R333 B.n182 B.n181 585
R334 B.n283 B.n282 585
R335 B.n282 B.n281 585
R336 B.n184 B.n183 585
R337 B.n185 B.n184 585
R338 B.n274 B.n273 585
R339 B.n275 B.n274 585
R340 B.n188 B.n187 585
R341 B.n213 B.n212 585
R342 B.n214 B.n210 585
R343 B.n210 B.n189 585
R344 B.n216 B.n215 585
R345 B.n218 B.n209 585
R346 B.n221 B.n220 585
R347 B.n222 B.n208 585
R348 B.n224 B.n223 585
R349 B.n226 B.n207 585
R350 B.n229 B.n228 585
R351 B.n230 B.n204 585
R352 B.n233 B.n232 585
R353 B.n235 B.n203 585
R354 B.n238 B.n237 585
R355 B.n239 B.n202 585
R356 B.n241 B.n240 585
R357 B.n243 B.n201 585
R358 B.n246 B.n245 585
R359 B.n247 B.n200 585
R360 B.n249 B.n248 585
R361 B.n251 B.n199 585
R362 B.n254 B.n253 585
R363 B.n255 B.n195 585
R364 B.n257 B.n256 585
R365 B.n259 B.n194 585
R366 B.n262 B.n261 585
R367 B.n263 B.n193 585
R368 B.n265 B.n264 585
R369 B.n267 B.n192 585
R370 B.n268 B.n191 585
R371 B.n271 B.n270 585
R372 B.n272 B.n190 585
R373 B.n190 B.n189 585
R374 B.n277 B.n276 585
R375 B.n276 B.n275 585
R376 B.n278 B.n186 585
R377 B.n186 B.n185 585
R378 B.n280 B.n279 585
R379 B.n281 B.n280 585
R380 B.n180 B.n179 585
R381 B.n181 B.n180 585
R382 B.n289 B.n288 585
R383 B.n288 B.n287 585
R384 B.n290 B.n178 585
R385 B.n178 B.n177 585
R386 B.n292 B.n291 585
R387 B.n293 B.n292 585
R388 B.n172 B.n171 585
R389 B.n173 B.n172 585
R390 B.n301 B.n300 585
R391 B.n300 B.n299 585
R392 B.n302 B.n170 585
R393 B.n170 B.n168 585
R394 B.n304 B.n303 585
R395 B.n305 B.n304 585
R396 B.n164 B.n163 585
R397 B.n169 B.n164 585
R398 B.n313 B.n312 585
R399 B.n312 B.n311 585
R400 B.n314 B.n162 585
R401 B.n162 B.n161 585
R402 B.n316 B.n315 585
R403 B.n317 B.n316 585
R404 B.n156 B.n155 585
R405 B.n157 B.n156 585
R406 B.n325 B.n324 585
R407 B.n324 B.n323 585
R408 B.n326 B.n154 585
R409 B.n154 B.n153 585
R410 B.n328 B.n327 585
R411 B.n329 B.n328 585
R412 B.n148 B.n147 585
R413 B.n149 B.n148 585
R414 B.n338 B.n337 585
R415 B.n337 B.n336 585
R416 B.n339 B.n146 585
R417 B.n335 B.n146 585
R418 B.n341 B.n340 585
R419 B.n342 B.n341 585
R420 B.n141 B.n140 585
R421 B.n142 B.n141 585
R422 B.n352 B.n351 585
R423 B.n351 B.n350 585
R424 B.n353 B.n139 585
R425 B.n349 B.n139 585
R426 B.n355 B.n354 585
R427 B.n356 B.n355 585
R428 B.n3 B.n0 585
R429 B.n4 B.n3 585
R430 B.n456 B.n1 585
R431 B.n457 B.n456 585
R432 B.n455 B.n454 585
R433 B.n455 B.n8 585
R434 B.n453 B.n9 585
R435 B.n12 B.n9 585
R436 B.n452 B.n451 585
R437 B.n451 B.n450 585
R438 B.n11 B.n10 585
R439 B.n449 B.n11 585
R440 B.n447 B.n446 585
R441 B.n448 B.n447 585
R442 B.n445 B.n16 585
R443 B.n19 B.n16 585
R444 B.n444 B.n443 585
R445 B.n443 B.n442 585
R446 B.n18 B.n17 585
R447 B.n441 B.n18 585
R448 B.n439 B.n438 585
R449 B.n440 B.n439 585
R450 B.n437 B.n24 585
R451 B.n24 B.n23 585
R452 B.n436 B.n435 585
R453 B.n435 B.n434 585
R454 B.n26 B.n25 585
R455 B.n433 B.n26 585
R456 B.n431 B.n430 585
R457 B.n432 B.n431 585
R458 B.n429 B.n31 585
R459 B.n31 B.n30 585
R460 B.n428 B.n427 585
R461 B.n427 B.n426 585
R462 B.n33 B.n32 585
R463 B.n425 B.n33 585
R464 B.n423 B.n422 585
R465 B.n424 B.n423 585
R466 B.n421 B.n38 585
R467 B.n38 B.n37 585
R468 B.n420 B.n419 585
R469 B.n419 B.n418 585
R470 B.n40 B.n39 585
R471 B.n417 B.n40 585
R472 B.n415 B.n414 585
R473 B.n416 B.n415 585
R474 B.n413 B.n45 585
R475 B.n45 B.n44 585
R476 B.n412 B.n411 585
R477 B.n411 B.n410 585
R478 B.n47 B.n46 585
R479 B.n409 B.n47 585
R480 B.n407 B.n406 585
R481 B.n408 B.n407 585
R482 B.n405 B.n52 585
R483 B.n52 B.n51 585
R484 B.n404 B.n403 585
R485 B.n403 B.n402 585
R486 B.n460 B.n459 585
R487 B.n458 B.n2 585
R488 B.n403 B.n54 545.355
R489 B.n399 B.n55 545.355
R490 B.n274 B.n190 545.355
R491 B.n276 B.n188 545.355
R492 B.n401 B.n400 256.663
R493 B.n401 B.n70 256.663
R494 B.n401 B.n69 256.663
R495 B.n401 B.n68 256.663
R496 B.n401 B.n67 256.663
R497 B.n401 B.n66 256.663
R498 B.n401 B.n65 256.663
R499 B.n401 B.n64 256.663
R500 B.n401 B.n63 256.663
R501 B.n401 B.n62 256.663
R502 B.n401 B.n61 256.663
R503 B.n401 B.n60 256.663
R504 B.n401 B.n59 256.663
R505 B.n401 B.n58 256.663
R506 B.n401 B.n57 256.663
R507 B.n401 B.n56 256.663
R508 B.n211 B.n189 256.663
R509 B.n217 B.n189 256.663
R510 B.n219 B.n189 256.663
R511 B.n225 B.n189 256.663
R512 B.n227 B.n189 256.663
R513 B.n234 B.n189 256.663
R514 B.n236 B.n189 256.663
R515 B.n242 B.n189 256.663
R516 B.n244 B.n189 256.663
R517 B.n250 B.n189 256.663
R518 B.n252 B.n189 256.663
R519 B.n258 B.n189 256.663
R520 B.n260 B.n189 256.663
R521 B.n266 B.n189 256.663
R522 B.n269 B.n189 256.663
R523 B.n462 B.n461 256.663
R524 B.n74 B.t16 251.85
R525 B.n72 B.t20 251.85
R526 B.n196 B.t9 251.85
R527 B.n205 B.t13 251.85
R528 B.n275 B.n189 202.571
R529 B.n402 B.n401 202.571
R530 B.n78 B.n77 163.367
R531 B.n82 B.n81 163.367
R532 B.n86 B.n85 163.367
R533 B.n90 B.n89 163.367
R534 B.n94 B.n93 163.367
R535 B.n99 B.n98 163.367
R536 B.n103 B.n102 163.367
R537 B.n107 B.n106 163.367
R538 B.n111 B.n110 163.367
R539 B.n115 B.n114 163.367
R540 B.n120 B.n119 163.367
R541 B.n124 B.n123 163.367
R542 B.n128 B.n127 163.367
R543 B.n132 B.n131 163.367
R544 B.n134 B.n71 163.367
R545 B.n274 B.n184 163.367
R546 B.n282 B.n184 163.367
R547 B.n282 B.n182 163.367
R548 B.n286 B.n182 163.367
R549 B.n286 B.n176 163.367
R550 B.n294 B.n176 163.367
R551 B.n294 B.n174 163.367
R552 B.n298 B.n174 163.367
R553 B.n298 B.n167 163.367
R554 B.n306 B.n167 163.367
R555 B.n306 B.n165 163.367
R556 B.n310 B.n165 163.367
R557 B.n310 B.n160 163.367
R558 B.n318 B.n160 163.367
R559 B.n318 B.n158 163.367
R560 B.n322 B.n158 163.367
R561 B.n322 B.n152 163.367
R562 B.n330 B.n152 163.367
R563 B.n330 B.n150 163.367
R564 B.n334 B.n150 163.367
R565 B.n334 B.n145 163.367
R566 B.n343 B.n145 163.367
R567 B.n343 B.n143 163.367
R568 B.n348 B.n143 163.367
R569 B.n348 B.n138 163.367
R570 B.n357 B.n138 163.367
R571 B.n358 B.n357 163.367
R572 B.n358 B.n5 163.367
R573 B.n6 B.n5 163.367
R574 B.n7 B.n6 163.367
R575 B.n364 B.n7 163.367
R576 B.n365 B.n364 163.367
R577 B.n365 B.n13 163.367
R578 B.n14 B.n13 163.367
R579 B.n15 B.n14 163.367
R580 B.n370 B.n15 163.367
R581 B.n370 B.n20 163.367
R582 B.n21 B.n20 163.367
R583 B.n22 B.n21 163.367
R584 B.n375 B.n22 163.367
R585 B.n375 B.n27 163.367
R586 B.n28 B.n27 163.367
R587 B.n29 B.n28 163.367
R588 B.n380 B.n29 163.367
R589 B.n380 B.n34 163.367
R590 B.n35 B.n34 163.367
R591 B.n36 B.n35 163.367
R592 B.n385 B.n36 163.367
R593 B.n385 B.n41 163.367
R594 B.n42 B.n41 163.367
R595 B.n43 B.n42 163.367
R596 B.n390 B.n43 163.367
R597 B.n390 B.n48 163.367
R598 B.n49 B.n48 163.367
R599 B.n50 B.n49 163.367
R600 B.n395 B.n50 163.367
R601 B.n395 B.n55 163.367
R602 B.n212 B.n210 163.367
R603 B.n216 B.n210 163.367
R604 B.n220 B.n218 163.367
R605 B.n224 B.n208 163.367
R606 B.n228 B.n226 163.367
R607 B.n233 B.n204 163.367
R608 B.n237 B.n235 163.367
R609 B.n241 B.n202 163.367
R610 B.n245 B.n243 163.367
R611 B.n249 B.n200 163.367
R612 B.n253 B.n251 163.367
R613 B.n257 B.n195 163.367
R614 B.n261 B.n259 163.367
R615 B.n265 B.n193 163.367
R616 B.n268 B.n267 163.367
R617 B.n270 B.n190 163.367
R618 B.n276 B.n186 163.367
R619 B.n280 B.n186 163.367
R620 B.n280 B.n180 163.367
R621 B.n288 B.n180 163.367
R622 B.n288 B.n178 163.367
R623 B.n292 B.n178 163.367
R624 B.n292 B.n172 163.367
R625 B.n300 B.n172 163.367
R626 B.n300 B.n170 163.367
R627 B.n304 B.n170 163.367
R628 B.n304 B.n164 163.367
R629 B.n312 B.n164 163.367
R630 B.n312 B.n162 163.367
R631 B.n316 B.n162 163.367
R632 B.n316 B.n156 163.367
R633 B.n324 B.n156 163.367
R634 B.n324 B.n154 163.367
R635 B.n328 B.n154 163.367
R636 B.n328 B.n148 163.367
R637 B.n337 B.n148 163.367
R638 B.n337 B.n146 163.367
R639 B.n341 B.n146 163.367
R640 B.n341 B.n141 163.367
R641 B.n351 B.n141 163.367
R642 B.n351 B.n139 163.367
R643 B.n355 B.n139 163.367
R644 B.n355 B.n3 163.367
R645 B.n460 B.n3 163.367
R646 B.n456 B.n2 163.367
R647 B.n456 B.n455 163.367
R648 B.n455 B.n9 163.367
R649 B.n451 B.n9 163.367
R650 B.n451 B.n11 163.367
R651 B.n447 B.n11 163.367
R652 B.n447 B.n16 163.367
R653 B.n443 B.n16 163.367
R654 B.n443 B.n18 163.367
R655 B.n439 B.n18 163.367
R656 B.n439 B.n24 163.367
R657 B.n435 B.n24 163.367
R658 B.n435 B.n26 163.367
R659 B.n431 B.n26 163.367
R660 B.n431 B.n31 163.367
R661 B.n427 B.n31 163.367
R662 B.n427 B.n33 163.367
R663 B.n423 B.n33 163.367
R664 B.n423 B.n38 163.367
R665 B.n419 B.n38 163.367
R666 B.n419 B.n40 163.367
R667 B.n415 B.n40 163.367
R668 B.n415 B.n45 163.367
R669 B.n411 B.n45 163.367
R670 B.n411 B.n47 163.367
R671 B.n407 B.n47 163.367
R672 B.n407 B.n52 163.367
R673 B.n403 B.n52 163.367
R674 B.n72 B.t21 140.28
R675 B.n196 B.t12 140.28
R676 B.n74 B.t18 140.279
R677 B.n205 B.t15 140.279
R678 B.n73 B.t22 117.782
R679 B.n197 B.t11 117.782
R680 B.n75 B.t19 117.781
R681 B.n206 B.t14 117.781
R682 B.n275 B.n185 106.781
R683 B.n281 B.n185 106.781
R684 B.n281 B.n181 106.781
R685 B.n287 B.n181 106.781
R686 B.n293 B.n177 106.781
R687 B.n293 B.n173 106.781
R688 B.n299 B.n173 106.781
R689 B.n299 B.n168 106.781
R690 B.n305 B.n168 106.781
R691 B.n305 B.n169 106.781
R692 B.n311 B.n161 106.781
R693 B.n317 B.n161 106.781
R694 B.n323 B.n157 106.781
R695 B.n323 B.n153 106.781
R696 B.n329 B.n153 106.781
R697 B.n336 B.n149 106.781
R698 B.n336 B.n335 106.781
R699 B.n342 B.n142 106.781
R700 B.n350 B.n142 106.781
R701 B.n350 B.n349 106.781
R702 B.n356 B.n4 106.781
R703 B.n459 B.n4 106.781
R704 B.n459 B.n458 106.781
R705 B.n458 B.n457 106.781
R706 B.n457 B.n8 106.781
R707 B.n450 B.n12 106.781
R708 B.n450 B.n449 106.781
R709 B.n449 B.n448 106.781
R710 B.n442 B.n19 106.781
R711 B.n442 B.n441 106.781
R712 B.n440 B.n23 106.781
R713 B.n434 B.n23 106.781
R714 B.n434 B.n433 106.781
R715 B.n432 B.n30 106.781
R716 B.n426 B.n30 106.781
R717 B.n425 B.n424 106.781
R718 B.n424 B.n37 106.781
R719 B.n418 B.n37 106.781
R720 B.n418 B.n417 106.781
R721 B.n417 B.n416 106.781
R722 B.n416 B.n44 106.781
R723 B.n410 B.n409 106.781
R724 B.n409 B.n408 106.781
R725 B.n408 B.n51 106.781
R726 B.n402 B.n51 106.781
R727 B.n317 B.t0 102.07
R728 B.t7 B.n432 102.07
R729 B.n287 B.t10 98.9298
R730 B.n410 B.t17 98.9298
R731 B.n356 B.t8 86.3674
R732 B.t23 B.n8 86.3674
R733 B.n335 B.t6 83.2268
R734 B.n19 B.t2 83.2268
R735 B.n56 B.n54 71.676
R736 B.n78 B.n57 71.676
R737 B.n82 B.n58 71.676
R738 B.n86 B.n59 71.676
R739 B.n90 B.n60 71.676
R740 B.n94 B.n61 71.676
R741 B.n99 B.n62 71.676
R742 B.n103 B.n63 71.676
R743 B.n107 B.n64 71.676
R744 B.n111 B.n65 71.676
R745 B.n115 B.n66 71.676
R746 B.n120 B.n67 71.676
R747 B.n124 B.n68 71.676
R748 B.n128 B.n69 71.676
R749 B.n132 B.n70 71.676
R750 B.n400 B.n71 71.676
R751 B.n400 B.n399 71.676
R752 B.n134 B.n70 71.676
R753 B.n131 B.n69 71.676
R754 B.n127 B.n68 71.676
R755 B.n123 B.n67 71.676
R756 B.n119 B.n66 71.676
R757 B.n114 B.n65 71.676
R758 B.n110 B.n64 71.676
R759 B.n106 B.n63 71.676
R760 B.n102 B.n62 71.676
R761 B.n98 B.n61 71.676
R762 B.n93 B.n60 71.676
R763 B.n89 B.n59 71.676
R764 B.n85 B.n58 71.676
R765 B.n81 B.n57 71.676
R766 B.n77 B.n56 71.676
R767 B.n211 B.n188 71.676
R768 B.n217 B.n216 71.676
R769 B.n220 B.n219 71.676
R770 B.n225 B.n224 71.676
R771 B.n228 B.n227 71.676
R772 B.n234 B.n233 71.676
R773 B.n237 B.n236 71.676
R774 B.n242 B.n241 71.676
R775 B.n245 B.n244 71.676
R776 B.n250 B.n249 71.676
R777 B.n253 B.n252 71.676
R778 B.n258 B.n257 71.676
R779 B.n261 B.n260 71.676
R780 B.n266 B.n265 71.676
R781 B.n269 B.n268 71.676
R782 B.n212 B.n211 71.676
R783 B.n218 B.n217 71.676
R784 B.n219 B.n208 71.676
R785 B.n226 B.n225 71.676
R786 B.n227 B.n204 71.676
R787 B.n235 B.n234 71.676
R788 B.n236 B.n202 71.676
R789 B.n243 B.n242 71.676
R790 B.n244 B.n200 71.676
R791 B.n251 B.n250 71.676
R792 B.n252 B.n195 71.676
R793 B.n259 B.n258 71.676
R794 B.n260 B.n193 71.676
R795 B.n267 B.n266 71.676
R796 B.n270 B.n269 71.676
R797 B.n461 B.n460 71.676
R798 B.n461 B.n2 71.676
R799 B.t4 B.n149 67.5237
R800 B.n441 B.t1 67.5237
R801 B.n96 B.n75 59.5399
R802 B.n117 B.n73 59.5399
R803 B.n198 B.n197 59.5399
R804 B.n231 B.n206 59.5399
R805 B.n169 B.t5 58.1019
R806 B.t3 B.n425 58.1019
R807 B.n311 B.t5 48.68
R808 B.n426 B.t3 48.68
R809 B.n329 B.t4 39.2582
R810 B.t1 B.n440 39.2582
R811 B.n277 B.n187 35.4346
R812 B.n273 B.n272 35.4346
R813 B.n404 B.n53 35.4346
R814 B.n398 B.n397 35.4346
R815 B.n342 B.t6 23.5551
R816 B.n448 B.t2 23.5551
R817 B.n75 B.n74 22.4975
R818 B.n73 B.n72 22.4975
R819 B.n197 B.n196 22.4975
R820 B.n206 B.n205 22.4975
R821 B.n349 B.t8 20.4145
R822 B.n12 B.t23 20.4145
R823 B B.n462 18.0485
R824 B.n278 B.n277 10.6151
R825 B.n279 B.n278 10.6151
R826 B.n279 B.n179 10.6151
R827 B.n289 B.n179 10.6151
R828 B.n290 B.n289 10.6151
R829 B.n291 B.n290 10.6151
R830 B.n291 B.n171 10.6151
R831 B.n301 B.n171 10.6151
R832 B.n302 B.n301 10.6151
R833 B.n303 B.n302 10.6151
R834 B.n303 B.n163 10.6151
R835 B.n313 B.n163 10.6151
R836 B.n314 B.n313 10.6151
R837 B.n315 B.n314 10.6151
R838 B.n315 B.n155 10.6151
R839 B.n325 B.n155 10.6151
R840 B.n326 B.n325 10.6151
R841 B.n327 B.n326 10.6151
R842 B.n327 B.n147 10.6151
R843 B.n338 B.n147 10.6151
R844 B.n339 B.n338 10.6151
R845 B.n340 B.n339 10.6151
R846 B.n340 B.n140 10.6151
R847 B.n352 B.n140 10.6151
R848 B.n353 B.n352 10.6151
R849 B.n354 B.n353 10.6151
R850 B.n354 B.n0 10.6151
R851 B.n213 B.n187 10.6151
R852 B.n214 B.n213 10.6151
R853 B.n215 B.n214 10.6151
R854 B.n215 B.n209 10.6151
R855 B.n221 B.n209 10.6151
R856 B.n222 B.n221 10.6151
R857 B.n223 B.n222 10.6151
R858 B.n223 B.n207 10.6151
R859 B.n229 B.n207 10.6151
R860 B.n230 B.n229 10.6151
R861 B.n232 B.n203 10.6151
R862 B.n238 B.n203 10.6151
R863 B.n239 B.n238 10.6151
R864 B.n240 B.n239 10.6151
R865 B.n240 B.n201 10.6151
R866 B.n246 B.n201 10.6151
R867 B.n247 B.n246 10.6151
R868 B.n248 B.n247 10.6151
R869 B.n248 B.n199 10.6151
R870 B.n255 B.n254 10.6151
R871 B.n256 B.n255 10.6151
R872 B.n256 B.n194 10.6151
R873 B.n262 B.n194 10.6151
R874 B.n263 B.n262 10.6151
R875 B.n264 B.n263 10.6151
R876 B.n264 B.n192 10.6151
R877 B.n192 B.n191 10.6151
R878 B.n271 B.n191 10.6151
R879 B.n272 B.n271 10.6151
R880 B.n273 B.n183 10.6151
R881 B.n283 B.n183 10.6151
R882 B.n284 B.n283 10.6151
R883 B.n285 B.n284 10.6151
R884 B.n285 B.n175 10.6151
R885 B.n295 B.n175 10.6151
R886 B.n296 B.n295 10.6151
R887 B.n297 B.n296 10.6151
R888 B.n297 B.n166 10.6151
R889 B.n307 B.n166 10.6151
R890 B.n308 B.n307 10.6151
R891 B.n309 B.n308 10.6151
R892 B.n309 B.n159 10.6151
R893 B.n319 B.n159 10.6151
R894 B.n320 B.n319 10.6151
R895 B.n321 B.n320 10.6151
R896 B.n321 B.n151 10.6151
R897 B.n331 B.n151 10.6151
R898 B.n332 B.n331 10.6151
R899 B.n333 B.n332 10.6151
R900 B.n333 B.n144 10.6151
R901 B.n344 B.n144 10.6151
R902 B.n345 B.n344 10.6151
R903 B.n347 B.n345 10.6151
R904 B.n347 B.n346 10.6151
R905 B.n346 B.n137 10.6151
R906 B.n359 B.n137 10.6151
R907 B.n360 B.n359 10.6151
R908 B.n361 B.n360 10.6151
R909 B.n362 B.n361 10.6151
R910 B.n363 B.n362 10.6151
R911 B.n366 B.n363 10.6151
R912 B.n367 B.n366 10.6151
R913 B.n368 B.n367 10.6151
R914 B.n369 B.n368 10.6151
R915 B.n371 B.n369 10.6151
R916 B.n372 B.n371 10.6151
R917 B.n373 B.n372 10.6151
R918 B.n374 B.n373 10.6151
R919 B.n376 B.n374 10.6151
R920 B.n377 B.n376 10.6151
R921 B.n378 B.n377 10.6151
R922 B.n379 B.n378 10.6151
R923 B.n381 B.n379 10.6151
R924 B.n382 B.n381 10.6151
R925 B.n383 B.n382 10.6151
R926 B.n384 B.n383 10.6151
R927 B.n386 B.n384 10.6151
R928 B.n387 B.n386 10.6151
R929 B.n388 B.n387 10.6151
R930 B.n389 B.n388 10.6151
R931 B.n391 B.n389 10.6151
R932 B.n392 B.n391 10.6151
R933 B.n393 B.n392 10.6151
R934 B.n394 B.n393 10.6151
R935 B.n396 B.n394 10.6151
R936 B.n397 B.n396 10.6151
R937 B.n454 B.n1 10.6151
R938 B.n454 B.n453 10.6151
R939 B.n453 B.n452 10.6151
R940 B.n452 B.n10 10.6151
R941 B.n446 B.n10 10.6151
R942 B.n446 B.n445 10.6151
R943 B.n445 B.n444 10.6151
R944 B.n444 B.n17 10.6151
R945 B.n438 B.n17 10.6151
R946 B.n438 B.n437 10.6151
R947 B.n437 B.n436 10.6151
R948 B.n436 B.n25 10.6151
R949 B.n430 B.n25 10.6151
R950 B.n430 B.n429 10.6151
R951 B.n429 B.n428 10.6151
R952 B.n428 B.n32 10.6151
R953 B.n422 B.n32 10.6151
R954 B.n422 B.n421 10.6151
R955 B.n421 B.n420 10.6151
R956 B.n420 B.n39 10.6151
R957 B.n414 B.n39 10.6151
R958 B.n414 B.n413 10.6151
R959 B.n413 B.n412 10.6151
R960 B.n412 B.n46 10.6151
R961 B.n406 B.n46 10.6151
R962 B.n406 B.n405 10.6151
R963 B.n405 B.n404 10.6151
R964 B.n76 B.n53 10.6151
R965 B.n79 B.n76 10.6151
R966 B.n80 B.n79 10.6151
R967 B.n83 B.n80 10.6151
R968 B.n84 B.n83 10.6151
R969 B.n87 B.n84 10.6151
R970 B.n88 B.n87 10.6151
R971 B.n91 B.n88 10.6151
R972 B.n92 B.n91 10.6151
R973 B.n95 B.n92 10.6151
R974 B.n100 B.n97 10.6151
R975 B.n101 B.n100 10.6151
R976 B.n104 B.n101 10.6151
R977 B.n105 B.n104 10.6151
R978 B.n108 B.n105 10.6151
R979 B.n109 B.n108 10.6151
R980 B.n112 B.n109 10.6151
R981 B.n113 B.n112 10.6151
R982 B.n116 B.n113 10.6151
R983 B.n121 B.n118 10.6151
R984 B.n122 B.n121 10.6151
R985 B.n125 B.n122 10.6151
R986 B.n126 B.n125 10.6151
R987 B.n129 B.n126 10.6151
R988 B.n130 B.n129 10.6151
R989 B.n133 B.n130 10.6151
R990 B.n135 B.n133 10.6151
R991 B.n136 B.n135 10.6151
R992 B.n398 B.n136 10.6151
R993 B.n231 B.n230 9.36635
R994 B.n254 B.n198 9.36635
R995 B.n96 B.n95 9.36635
R996 B.n118 B.n117 9.36635
R997 B.n462 B.n0 8.11757
R998 B.n462 B.n1 8.11757
R999 B.t10 B.n177 7.85203
R1000 B.t17 B.n44 7.85203
R1001 B.t0 B.n157 4.71142
R1002 B.n433 B.t7 4.71142
R1003 B.n232 B.n231 1.24928
R1004 B.n199 B.n198 1.24928
R1005 B.n97 B.n96 1.24928
R1006 B.n117 B.n116 1.24928
R1007 VN.n17 VN.n16 161.3
R1008 VN.n35 VN.n34 161.3
R1009 VN.n33 VN.n18 161.3
R1010 VN.n32 VN.n31 161.3
R1011 VN.n30 VN.n29 161.3
R1012 VN.n28 VN.n20 161.3
R1013 VN.n26 VN.n25 161.3
R1014 VN.n24 VN.n21 161.3
R1015 VN.n15 VN.n0 161.3
R1016 VN.n14 VN.n13 161.3
R1017 VN.n12 VN.n11 161.3
R1018 VN.n10 VN.n2 161.3
R1019 VN.n8 VN.n7 161.3
R1020 VN.n6 VN.n3 161.3
R1021 VN.n5 VN.t0 122.052
R1022 VN.n23 VN.t3 122.052
R1023 VN.n16 VN.t9 97.8523
R1024 VN.n34 VN.t7 97.8523
R1025 VN.n8 VN.n3 56.5193
R1026 VN.n11 VN.n10 56.5193
R1027 VN.n26 VN.n21 56.5193
R1028 VN.n29 VN.n28 56.5193
R1029 VN.n4 VN.t1 50.233
R1030 VN.n9 VN.t8 50.233
R1031 VN.n1 VN.t4 50.233
R1032 VN.n22 VN.t2 50.233
R1033 VN.n27 VN.t5 50.233
R1034 VN.n19 VN.t6 50.233
R1035 VN.n24 VN.n23 42.3937
R1036 VN.n6 VN.n5 42.3937
R1037 VN.n15 VN.n14 41.4647
R1038 VN.n33 VN.n32 41.4647
R1039 VN VN.n35 36.1312
R1040 VN.n5 VN.n4 33.4547
R1041 VN.n23 VN.n22 33.4547
R1042 VN.n16 VN.n15 22.6399
R1043 VN.n34 VN.n33 22.6399
R1044 VN.n4 VN.n3 20.0634
R1045 VN.n11 VN.n1 20.0634
R1046 VN.n22 VN.n21 20.0634
R1047 VN.n29 VN.n19 20.0634
R1048 VN.n9 VN.n8 12.234
R1049 VN.n10 VN.n9 12.234
R1050 VN.n28 VN.n27 12.234
R1051 VN.n27 VN.n26 12.234
R1052 VN.n14 VN.n1 4.40456
R1053 VN.n32 VN.n19 4.40456
R1054 VN.n35 VN.n18 0.189894
R1055 VN.n31 VN.n18 0.189894
R1056 VN.n31 VN.n30 0.189894
R1057 VN.n30 VN.n20 0.189894
R1058 VN.n25 VN.n20 0.189894
R1059 VN.n25 VN.n24 0.189894
R1060 VN.n7 VN.n6 0.189894
R1061 VN.n7 VN.n2 0.189894
R1062 VN.n12 VN.n2 0.189894
R1063 VN.n13 VN.n12 0.189894
R1064 VN.n13 VN.n0 0.189894
R1065 VN.n17 VN.n0 0.189894
R1066 VN VN.n17 0.0516364
R1067 VDD2.n13 VDD2.n11 289.615
R1068 VDD2.n2 VDD2.n0 289.615
R1069 VDD2.n14 VDD2.n13 185
R1070 VDD2.n3 VDD2.n2 185
R1071 VDD2.t2 VDD2.n12 164.876
R1072 VDD2.t9 VDD2.n1 164.876
R1073 VDD2.n10 VDD2.n9 101.147
R1074 VDD2 VDD2.n21 101.145
R1075 VDD2.n20 VDD2.n19 100.454
R1076 VDD2.n8 VDD2.n7 100.454
R1077 VDD2.n13 VDD2.t2 52.3082
R1078 VDD2.n2 VDD2.t9 52.3082
R1079 VDD2.n8 VDD2.n6 50.8338
R1080 VDD2.n18 VDD2.n17 49.8338
R1081 VDD2.n18 VDD2.n10 29.9567
R1082 VDD2.n14 VDD2.n12 14.7318
R1083 VDD2.n3 VDD2.n1 14.7318
R1084 VDD2.n15 VDD2.n11 12.8005
R1085 VDD2.n4 VDD2.n0 12.8005
R1086 VDD2.n21 VDD2.t7 11.4456
R1087 VDD2.n21 VDD2.t6 11.4456
R1088 VDD2.n19 VDD2.t3 11.4456
R1089 VDD2.n19 VDD2.t4 11.4456
R1090 VDD2.n9 VDD2.t5 11.4456
R1091 VDD2.n9 VDD2.t0 11.4456
R1092 VDD2.n7 VDD2.t8 11.4456
R1093 VDD2.n7 VDD2.t1 11.4456
R1094 VDD2.n17 VDD2.n16 9.45567
R1095 VDD2.n6 VDD2.n5 9.45567
R1096 VDD2.n16 VDD2.n15 9.3005
R1097 VDD2.n5 VDD2.n4 9.3005
R1098 VDD2.n16 VDD2.n12 5.62509
R1099 VDD2.n5 VDD2.n1 5.62509
R1100 VDD2.n17 VDD2.n11 1.16414
R1101 VDD2.n6 VDD2.n0 1.16414
R1102 VDD2.n20 VDD2.n18 1.0005
R1103 VDD2.n15 VDD2.n14 0.388379
R1104 VDD2.n4 VDD2.n3 0.388379
R1105 VDD2 VDD2.n20 0.30869
R1106 VDD2.n10 VDD2.n8 0.195154
C0 VN VTAIL 1.88316f
C1 VDD1 VN 0.156017f
C2 VP VTAIL 1.89733f
C3 VN VDD2 1.43389f
C4 VP VDD1 1.63987f
C5 VP VDD2 0.364241f
C6 VP VN 3.8935f
C7 VDD1 VTAIL 4.1927f
C8 VTAIL VDD2 4.23356f
C9 VDD1 VDD2 1.05027f
C10 VDD2 B 3.15236f
C11 VDD1 B 3.192209f
C12 VTAIL B 2.578878f
C13 VN B 8.148117f
C14 VP B 7.240658f
C15 VDD2.n0 B 0.023023f
C16 VDD2.n1 B 0.053931f
C17 VDD2.t9 B 0.038976f
C18 VDD2.n2 B 0.039748f
C19 VDD2.n3 B 0.011931f
C20 VDD2.n4 B 0.009685f
C21 VDD2.n5 B 0.104569f
C22 VDD2.n6 B 0.039334f
C23 VDD2.t8 B 0.024639f
C24 VDD2.t1 B 0.024639f
C25 VDD2.n7 B 0.157371f
C26 VDD2.n8 B 0.286108f
C27 VDD2.t5 B 0.024639f
C28 VDD2.t0 B 0.024639f
C29 VDD2.n9 B 0.158945f
C30 VDD2.n10 B 0.965566f
C31 VDD2.n11 B 0.023023f
C32 VDD2.n12 B 0.053931f
C33 VDD2.t2 B 0.038976f
C34 VDD2.n13 B 0.039748f
C35 VDD2.n14 B 0.011931f
C36 VDD2.n15 B 0.009685f
C37 VDD2.n16 B 0.104569f
C38 VDD2.n17 B 0.037495f
C39 VDD2.n18 B 0.994167f
C40 VDD2.t3 B 0.024639f
C41 VDD2.t4 B 0.024639f
C42 VDD2.n19 B 0.157371f
C43 VDD2.n20 B 0.19891f
C44 VDD2.t7 B 0.024639f
C45 VDD2.t6 B 0.024639f
C46 VDD2.n21 B 0.158934f
C47 VN.n0 B 0.023894f
C48 VN.t4 B 0.077623f
C49 VN.n1 B 0.054035f
C50 VN.n2 B 0.023894f
C51 VN.t8 B 0.077623f
C52 VN.n3 B 0.025596f
C53 VN.t0 B 0.124453f
C54 VN.t1 B 0.077623f
C55 VN.n4 B 0.081494f
C56 VN.n5 B 0.075218f
C57 VN.n6 B 0.101975f
C58 VN.n7 B 0.023894f
C59 VN.n8 B 0.029214f
C60 VN.n9 B 0.054035f
C61 VN.n10 B 0.029214f
C62 VN.n11 B 0.025596f
C63 VN.n12 B 0.023894f
C64 VN.n13 B 0.023894f
C65 VN.n14 B 0.029205f
C66 VN.n15 B 0.011892f
C67 VN.t9 B 0.108006f
C68 VN.n16 B 0.077503f
C69 VN.n17 B 0.018517f
C70 VN.n18 B 0.023894f
C71 VN.t6 B 0.077623f
C72 VN.n19 B 0.054035f
C73 VN.n20 B 0.023894f
C74 VN.t5 B 0.077623f
C75 VN.n21 B 0.025596f
C76 VN.t3 B 0.124453f
C77 VN.t2 B 0.077623f
C78 VN.n22 B 0.081494f
C79 VN.n23 B 0.075218f
C80 VN.n24 B 0.101975f
C81 VN.n25 B 0.023894f
C82 VN.n26 B 0.029214f
C83 VN.n27 B 0.054035f
C84 VN.n28 B 0.029214f
C85 VN.n29 B 0.025596f
C86 VN.n30 B 0.023894f
C87 VN.n31 B 0.023894f
C88 VN.n32 B 0.029205f
C89 VN.n33 B 0.011892f
C90 VN.t7 B 0.108006f
C91 VN.n34 B 0.077503f
C92 VN.n35 B 0.757274f
C93 VTAIL.t19 B 0.031544f
C94 VTAIL.t2 B 0.031544f
C95 VTAIL.n0 B 0.171008f
C96 VTAIL.n1 B 0.288676f
C97 VTAIL.n2 B 0.029474f
C98 VTAIL.n3 B 0.069042f
C99 VTAIL.t14 B 0.049897f
C100 VTAIL.n4 B 0.050885f
C101 VTAIL.n5 B 0.015275f
C102 VTAIL.n6 B 0.012399f
C103 VTAIL.n7 B 0.13387f
C104 VTAIL.n8 B 0.032082f
C105 VTAIL.n9 B 0.167048f
C106 VTAIL.t16 B 0.031544f
C107 VTAIL.t11 B 0.031544f
C108 VTAIL.n10 B 0.171008f
C109 VTAIL.n11 B 0.30518f
C110 VTAIL.t10 B 0.031544f
C111 VTAIL.t12 B 0.031544f
C112 VTAIL.n12 B 0.171008f
C113 VTAIL.n13 B 0.803832f
C114 VTAIL.t5 B 0.031544f
C115 VTAIL.t0 B 0.031544f
C116 VTAIL.n14 B 0.171009f
C117 VTAIL.n15 B 0.803831f
C118 VTAIL.t4 B 0.031544f
C119 VTAIL.t6 B 0.031544f
C120 VTAIL.n16 B 0.171009f
C121 VTAIL.n17 B 0.305178f
C122 VTAIL.n18 B 0.029474f
C123 VTAIL.n19 B 0.069042f
C124 VTAIL.t8 B 0.049897f
C125 VTAIL.n20 B 0.050885f
C126 VTAIL.n21 B 0.015275f
C127 VTAIL.n22 B 0.012399f
C128 VTAIL.n23 B 0.13387f
C129 VTAIL.n24 B 0.032082f
C130 VTAIL.n25 B 0.167048f
C131 VTAIL.t17 B 0.031544f
C132 VTAIL.t18 B 0.031544f
C133 VTAIL.n26 B 0.171009f
C134 VTAIL.n27 B 0.302935f
C135 VTAIL.t9 B 0.031544f
C136 VTAIL.t13 B 0.031544f
C137 VTAIL.n28 B 0.171009f
C138 VTAIL.n29 B 0.305178f
C139 VTAIL.n30 B 0.029474f
C140 VTAIL.n31 B 0.069042f
C141 VTAIL.t15 B 0.049897f
C142 VTAIL.n32 B 0.050885f
C143 VTAIL.n33 B 0.015275f
C144 VTAIL.n34 B 0.012399f
C145 VTAIL.n35 B 0.13387f
C146 VTAIL.n36 B 0.032082f
C147 VTAIL.n37 B 0.593597f
C148 VTAIL.n38 B 0.029474f
C149 VTAIL.n39 B 0.069042f
C150 VTAIL.t3 B 0.049897f
C151 VTAIL.n40 B 0.050885f
C152 VTAIL.n41 B 0.015275f
C153 VTAIL.n42 B 0.012399f
C154 VTAIL.n43 B 0.13387f
C155 VTAIL.n44 B 0.032082f
C156 VTAIL.n45 B 0.593597f
C157 VTAIL.t1 B 0.031544f
C158 VTAIL.t7 B 0.031544f
C159 VTAIL.n46 B 0.171008f
C160 VTAIL.n47 B 0.245093f
C161 VDD1.n0 B 0.022664f
C162 VDD1.n1 B 0.053089f
C163 VDD1.t2 B 0.038367f
C164 VDD1.n2 B 0.039127f
C165 VDD1.n3 B 0.011745f
C166 VDD1.n4 B 0.009534f
C167 VDD1.n5 B 0.102937f
C168 VDD1.n6 B 0.03872f
C169 VDD1.t0 B 0.024255f
C170 VDD1.t5 B 0.024255f
C171 VDD1.n7 B 0.154916f
C172 VDD1.n8 B 0.286021f
C173 VDD1.n9 B 0.022664f
C174 VDD1.n10 B 0.053089f
C175 VDD1.t6 B 0.038367f
C176 VDD1.n11 B 0.039127f
C177 VDD1.n12 B 0.011745f
C178 VDD1.n13 B 0.009534f
C179 VDD1.n14 B 0.102937f
C180 VDD1.n15 B 0.03872f
C181 VDD1.t3 B 0.024255f
C182 VDD1.t9 B 0.024255f
C183 VDD1.n16 B 0.154915f
C184 VDD1.n17 B 0.281645f
C185 VDD1.t1 B 0.024255f
C186 VDD1.t7 B 0.024255f
C187 VDD1.n18 B 0.156465f
C188 VDD1.n19 B 1.00338f
C189 VDD1.t4 B 0.024255f
C190 VDD1.t8 B 0.024255f
C191 VDD1.n20 B 0.154916f
C192 VDD1.n21 B 1.12416f
C193 VP.n0 B 0.024101f
C194 VP.t7 B 0.078298f
C195 VP.n1 B 0.054505f
C196 VP.n2 B 0.024101f
C197 VP.t2 B 0.078298f
C198 VP.n3 B 0.025819f
C199 VP.n4 B 0.024101f
C200 VP.n5 B 0.024101f
C201 VP.t3 B 0.108944f
C202 VP.t5 B 0.078298f
C203 VP.n6 B 0.054505f
C204 VP.n7 B 0.024101f
C205 VP.t9 B 0.078298f
C206 VP.n8 B 0.025819f
C207 VP.t0 B 0.078298f
C208 VP.n9 B 0.082202f
C209 VP.t1 B 0.125534f
C210 VP.n10 B 0.075872f
C211 VP.n11 B 0.102861f
C212 VP.n12 B 0.024101f
C213 VP.n13 B 0.029468f
C214 VP.n14 B 0.054505f
C215 VP.n15 B 0.029468f
C216 VP.n16 B 0.025819f
C217 VP.n17 B 0.024101f
C218 VP.n18 B 0.024101f
C219 VP.n19 B 0.029459f
C220 VP.n20 B 0.011995f
C221 VP.n21 B 0.078177f
C222 VP.n22 B 0.747858f
C223 VP.n23 B 0.772092f
C224 VP.t8 B 0.108944f
C225 VP.n24 B 0.078177f
C226 VP.n25 B 0.011995f
C227 VP.t6 B 0.078298f
C228 VP.n26 B 0.054505f
C229 VP.n27 B 0.029459f
C230 VP.n28 B 0.024101f
C231 VP.n29 B 0.024101f
C232 VP.n30 B 0.024101f
C233 VP.n31 B 0.029468f
C234 VP.n32 B 0.054505f
C235 VP.n33 B 0.029468f
C236 VP.n34 B 0.025819f
C237 VP.n35 B 0.024101f
C238 VP.n36 B 0.024101f
C239 VP.n37 B 0.029459f
C240 VP.n38 B 0.011995f
C241 VP.t4 B 0.108944f
C242 VP.n39 B 0.078177f
C243 VP.n40 B 0.018677f
.ends

