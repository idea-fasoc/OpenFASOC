* NGSPICE file created from diff_pair_sample_0357.ext - technology: sky130A

.subckt diff_pair_sample_0357 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t9 VN.t0 VTAIL.t12 B.t3 sky130_fd_pr__nfet_01v8 ad=2.2737 pd=14.11 as=2.2737 ps=14.11 w=13.78 l=2.37
X1 VTAIL.t8 VN.t1 VDD2.t8 B.t9 sky130_fd_pr__nfet_01v8 ad=2.2737 pd=14.11 as=2.2737 ps=14.11 w=13.78 l=2.37
X2 VTAIL.t14 VP.t0 VDD1.t9 B.t9 sky130_fd_pr__nfet_01v8 ad=2.2737 pd=14.11 as=2.2737 ps=14.11 w=13.78 l=2.37
X3 B.t23 B.t21 B.t22 B.t18 sky130_fd_pr__nfet_01v8 ad=5.3742 pd=28.34 as=0 ps=0 w=13.78 l=2.37
X4 VDD1.t8 VP.t1 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=5.3742 pd=28.34 as=2.2737 ps=14.11 w=13.78 l=2.37
X5 VDD1.t7 VP.t2 VTAIL.t19 B.t8 sky130_fd_pr__nfet_01v8 ad=2.2737 pd=14.11 as=5.3742 ps=28.34 w=13.78 l=2.37
X6 B.t20 B.t17 B.t19 B.t18 sky130_fd_pr__nfet_01v8 ad=5.3742 pd=28.34 as=0 ps=0 w=13.78 l=2.37
X7 VDD1.t6 VP.t3 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=2.2737 pd=14.11 as=2.2737 ps=14.11 w=13.78 l=2.37
X8 VTAIL.t11 VN.t2 VDD2.t7 B.t2 sky130_fd_pr__nfet_01v8 ad=2.2737 pd=14.11 as=2.2737 ps=14.11 w=13.78 l=2.37
X9 VDD2.t6 VN.t3 VTAIL.t9 B.t8 sky130_fd_pr__nfet_01v8 ad=2.2737 pd=14.11 as=5.3742 ps=28.34 w=13.78 l=2.37
X10 VTAIL.t2 VP.t4 VDD1.t5 B.t2 sky130_fd_pr__nfet_01v8 ad=2.2737 pd=14.11 as=2.2737 ps=14.11 w=13.78 l=2.37
X11 VTAIL.t4 VN.t4 VDD2.t5 B.t1 sky130_fd_pr__nfet_01v8 ad=2.2737 pd=14.11 as=2.2737 ps=14.11 w=13.78 l=2.37
X12 VDD1.t4 VP.t5 VTAIL.t15 B.t4 sky130_fd_pr__nfet_01v8 ad=5.3742 pd=28.34 as=2.2737 ps=14.11 w=13.78 l=2.37
X13 VDD1.t3 VP.t6 VTAIL.t16 B.t7 sky130_fd_pr__nfet_01v8 ad=2.2737 pd=14.11 as=5.3742 ps=28.34 w=13.78 l=2.37
X14 B.t16 B.t14 B.t15 B.t11 sky130_fd_pr__nfet_01v8 ad=5.3742 pd=28.34 as=0 ps=0 w=13.78 l=2.37
X15 VDD2.t4 VN.t5 VTAIL.t7 B.t7 sky130_fd_pr__nfet_01v8 ad=2.2737 pd=14.11 as=5.3742 ps=28.34 w=13.78 l=2.37
X16 B.t13 B.t10 B.t12 B.t11 sky130_fd_pr__nfet_01v8 ad=5.3742 pd=28.34 as=0 ps=0 w=13.78 l=2.37
X17 VTAIL.t13 VN.t6 VDD2.t3 B.t6 sky130_fd_pr__nfet_01v8 ad=2.2737 pd=14.11 as=2.2737 ps=14.11 w=13.78 l=2.37
X18 VDD1.t2 VP.t7 VTAIL.t17 B.t5 sky130_fd_pr__nfet_01v8 ad=2.2737 pd=14.11 as=2.2737 ps=14.11 w=13.78 l=2.37
X19 VTAIL.t18 VP.t8 VDD1.t1 B.t6 sky130_fd_pr__nfet_01v8 ad=2.2737 pd=14.11 as=2.2737 ps=14.11 w=13.78 l=2.37
X20 VDD2.t2 VN.t7 VTAIL.t10 B.t0 sky130_fd_pr__nfet_01v8 ad=5.3742 pd=28.34 as=2.2737 ps=14.11 w=13.78 l=2.37
X21 VTAIL.t1 VP.t9 VDD1.t0 B.t1 sky130_fd_pr__nfet_01v8 ad=2.2737 pd=14.11 as=2.2737 ps=14.11 w=13.78 l=2.37
X22 VDD2.t1 VN.t8 VTAIL.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=2.2737 pd=14.11 as=2.2737 ps=14.11 w=13.78 l=2.37
X23 VDD2.t0 VN.t9 VTAIL.t6 B.t4 sky130_fd_pr__nfet_01v8 ad=5.3742 pd=28.34 as=2.2737 ps=14.11 w=13.78 l=2.37
R0 VN.n9 VN.t9 173.024
R1 VN.n47 VN.t5 173.024
R2 VN.n73 VN.n38 161.3
R3 VN.n72 VN.n71 161.3
R4 VN.n70 VN.n39 161.3
R5 VN.n69 VN.n68 161.3
R6 VN.n67 VN.n40 161.3
R7 VN.n66 VN.n65 161.3
R8 VN.n64 VN.n63 161.3
R9 VN.n62 VN.n42 161.3
R10 VN.n61 VN.n60 161.3
R11 VN.n59 VN.n43 161.3
R12 VN.n58 VN.n57 161.3
R13 VN.n55 VN.n44 161.3
R14 VN.n54 VN.n53 161.3
R15 VN.n52 VN.n45 161.3
R16 VN.n51 VN.n50 161.3
R17 VN.n49 VN.n46 161.3
R18 VN.n35 VN.n0 161.3
R19 VN.n34 VN.n33 161.3
R20 VN.n32 VN.n1 161.3
R21 VN.n31 VN.n30 161.3
R22 VN.n29 VN.n2 161.3
R23 VN.n28 VN.n27 161.3
R24 VN.n26 VN.n25 161.3
R25 VN.n24 VN.n4 161.3
R26 VN.n23 VN.n22 161.3
R27 VN.n21 VN.n5 161.3
R28 VN.n20 VN.n19 161.3
R29 VN.n17 VN.n6 161.3
R30 VN.n16 VN.n15 161.3
R31 VN.n14 VN.n7 161.3
R32 VN.n13 VN.n12 161.3
R33 VN.n11 VN.n8 161.3
R34 VN.n10 VN.t4 140.126
R35 VN.n18 VN.t0 140.126
R36 VN.n3 VN.t6 140.126
R37 VN.n36 VN.t3 140.126
R38 VN.n48 VN.t1 140.126
R39 VN.n56 VN.t8 140.126
R40 VN.n41 VN.t2 140.126
R41 VN.n74 VN.t7 140.126
R42 VN.n37 VN.n36 103.531
R43 VN.n75 VN.n74 103.531
R44 VN.n30 VN.n1 56.5617
R45 VN.n68 VN.n39 56.5617
R46 VN VN.n75 53.4149
R47 VN.n10 VN.n9 50.3824
R48 VN.n48 VN.n47 50.3824
R49 VN.n12 VN.n7 50.2647
R50 VN.n24 VN.n23 50.2647
R51 VN.n50 VN.n45 50.2647
R52 VN.n62 VN.n61 50.2647
R53 VN.n16 VN.n7 30.8893
R54 VN.n23 VN.n5 30.8893
R55 VN.n54 VN.n45 30.8893
R56 VN.n61 VN.n43 30.8893
R57 VN.n12 VN.n11 24.5923
R58 VN.n17 VN.n16 24.5923
R59 VN.n19 VN.n5 24.5923
R60 VN.n25 VN.n24 24.5923
R61 VN.n29 VN.n28 24.5923
R62 VN.n30 VN.n29 24.5923
R63 VN.n34 VN.n1 24.5923
R64 VN.n35 VN.n34 24.5923
R65 VN.n50 VN.n49 24.5923
R66 VN.n57 VN.n43 24.5923
R67 VN.n55 VN.n54 24.5923
R68 VN.n68 VN.n67 24.5923
R69 VN.n67 VN.n66 24.5923
R70 VN.n63 VN.n62 24.5923
R71 VN.n73 VN.n72 24.5923
R72 VN.n72 VN.n39 24.5923
R73 VN.n11 VN.n10 22.1332
R74 VN.n25 VN.n3 22.1332
R75 VN.n49 VN.n48 22.1332
R76 VN.n63 VN.n41 22.1332
R77 VN.n18 VN.n17 12.2964
R78 VN.n19 VN.n18 12.2964
R79 VN.n57 VN.n56 12.2964
R80 VN.n56 VN.n55 12.2964
R81 VN.n36 VN.n35 7.37805
R82 VN.n74 VN.n73 7.37805
R83 VN.n47 VN.n46 6.9978
R84 VN.n9 VN.n8 6.9978
R85 VN.n28 VN.n3 2.45968
R86 VN.n66 VN.n41 2.45968
R87 VN.n75 VN.n38 0.278335
R88 VN.n37 VN.n0 0.278335
R89 VN.n71 VN.n38 0.189894
R90 VN.n71 VN.n70 0.189894
R91 VN.n70 VN.n69 0.189894
R92 VN.n69 VN.n40 0.189894
R93 VN.n65 VN.n40 0.189894
R94 VN.n65 VN.n64 0.189894
R95 VN.n64 VN.n42 0.189894
R96 VN.n60 VN.n42 0.189894
R97 VN.n60 VN.n59 0.189894
R98 VN.n59 VN.n58 0.189894
R99 VN.n58 VN.n44 0.189894
R100 VN.n53 VN.n44 0.189894
R101 VN.n53 VN.n52 0.189894
R102 VN.n52 VN.n51 0.189894
R103 VN.n51 VN.n46 0.189894
R104 VN.n13 VN.n8 0.189894
R105 VN.n14 VN.n13 0.189894
R106 VN.n15 VN.n14 0.189894
R107 VN.n15 VN.n6 0.189894
R108 VN.n20 VN.n6 0.189894
R109 VN.n21 VN.n20 0.189894
R110 VN.n22 VN.n21 0.189894
R111 VN.n22 VN.n4 0.189894
R112 VN.n26 VN.n4 0.189894
R113 VN.n27 VN.n26 0.189894
R114 VN.n27 VN.n2 0.189894
R115 VN.n31 VN.n2 0.189894
R116 VN.n32 VN.n31 0.189894
R117 VN.n33 VN.n32 0.189894
R118 VN.n33 VN.n0 0.189894
R119 VN VN.n37 0.153485
R120 VTAIL.n11 VTAIL.t7 50.0919
R121 VTAIL.n17 VTAIL.t9 50.0917
R122 VTAIL.n2 VTAIL.t16 50.0917
R123 VTAIL.n16 VTAIL.t19 50.0917
R124 VTAIL.n15 VTAIL.n14 48.655
R125 VTAIL.n13 VTAIL.n12 48.655
R126 VTAIL.n10 VTAIL.n9 48.655
R127 VTAIL.n8 VTAIL.n7 48.655
R128 VTAIL.n19 VTAIL.n18 48.6548
R129 VTAIL.n1 VTAIL.n0 48.6548
R130 VTAIL.n4 VTAIL.n3 48.6548
R131 VTAIL.n6 VTAIL.n5 48.6548
R132 VTAIL.n8 VTAIL.n6 28.9014
R133 VTAIL.n17 VTAIL.n16 26.5738
R134 VTAIL.n10 VTAIL.n8 2.32809
R135 VTAIL.n11 VTAIL.n10 2.32809
R136 VTAIL.n15 VTAIL.n13 2.32809
R137 VTAIL.n16 VTAIL.n15 2.32809
R138 VTAIL.n6 VTAIL.n4 2.32809
R139 VTAIL.n4 VTAIL.n2 2.32809
R140 VTAIL.n19 VTAIL.n17 2.32809
R141 VTAIL VTAIL.n1 1.80438
R142 VTAIL.n13 VTAIL.n11 1.63412
R143 VTAIL.n2 VTAIL.n1 1.63412
R144 VTAIL.n18 VTAIL.t12 1.43736
R145 VTAIL.n18 VTAIL.t13 1.43736
R146 VTAIL.n0 VTAIL.t6 1.43736
R147 VTAIL.n0 VTAIL.t4 1.43736
R148 VTAIL.n3 VTAIL.t17 1.43736
R149 VTAIL.n3 VTAIL.t14 1.43736
R150 VTAIL.n5 VTAIL.t0 1.43736
R151 VTAIL.n5 VTAIL.t2 1.43736
R152 VTAIL.n14 VTAIL.t3 1.43736
R153 VTAIL.n14 VTAIL.t18 1.43736
R154 VTAIL.n12 VTAIL.t15 1.43736
R155 VTAIL.n12 VTAIL.t1 1.43736
R156 VTAIL.n9 VTAIL.t5 1.43736
R157 VTAIL.n9 VTAIL.t8 1.43736
R158 VTAIL.n7 VTAIL.t10 1.43736
R159 VTAIL.n7 VTAIL.t11 1.43736
R160 VTAIL VTAIL.n19 0.524207
R161 VDD2.n1 VDD2.t0 69.098
R162 VDD2.n3 VDD2.n2 67.0239
R163 VDD2 VDD2.n7 67.0211
R164 VDD2.n4 VDD2.t2 66.7707
R165 VDD2.n6 VDD2.n5 65.3338
R166 VDD2.n1 VDD2.n0 65.3336
R167 VDD2.n4 VDD2.n3 46.6506
R168 VDD2.n6 VDD2.n4 2.32809
R169 VDD2.n7 VDD2.t8 1.43736
R170 VDD2.n7 VDD2.t4 1.43736
R171 VDD2.n5 VDD2.t7 1.43736
R172 VDD2.n5 VDD2.t1 1.43736
R173 VDD2.n2 VDD2.t3 1.43736
R174 VDD2.n2 VDD2.t6 1.43736
R175 VDD2.n0 VDD2.t5 1.43736
R176 VDD2.n0 VDD2.t9 1.43736
R177 VDD2 VDD2.n6 0.640586
R178 VDD2.n3 VDD2.n1 0.527051
R179 B.n969 B.n968 585
R180 B.n970 B.n969 585
R181 B.n360 B.n154 585
R182 B.n359 B.n358 585
R183 B.n357 B.n356 585
R184 B.n355 B.n354 585
R185 B.n353 B.n352 585
R186 B.n351 B.n350 585
R187 B.n349 B.n348 585
R188 B.n347 B.n346 585
R189 B.n345 B.n344 585
R190 B.n343 B.n342 585
R191 B.n341 B.n340 585
R192 B.n339 B.n338 585
R193 B.n337 B.n336 585
R194 B.n335 B.n334 585
R195 B.n333 B.n332 585
R196 B.n331 B.n330 585
R197 B.n329 B.n328 585
R198 B.n327 B.n326 585
R199 B.n325 B.n324 585
R200 B.n323 B.n322 585
R201 B.n321 B.n320 585
R202 B.n319 B.n318 585
R203 B.n317 B.n316 585
R204 B.n315 B.n314 585
R205 B.n313 B.n312 585
R206 B.n311 B.n310 585
R207 B.n309 B.n308 585
R208 B.n307 B.n306 585
R209 B.n305 B.n304 585
R210 B.n303 B.n302 585
R211 B.n301 B.n300 585
R212 B.n299 B.n298 585
R213 B.n297 B.n296 585
R214 B.n295 B.n294 585
R215 B.n293 B.n292 585
R216 B.n291 B.n290 585
R217 B.n289 B.n288 585
R218 B.n287 B.n286 585
R219 B.n285 B.n284 585
R220 B.n283 B.n282 585
R221 B.n281 B.n280 585
R222 B.n279 B.n278 585
R223 B.n277 B.n276 585
R224 B.n275 B.n274 585
R225 B.n273 B.n272 585
R226 B.n271 B.n270 585
R227 B.n269 B.n268 585
R228 B.n267 B.n266 585
R229 B.n265 B.n264 585
R230 B.n263 B.n262 585
R231 B.n261 B.n260 585
R232 B.n259 B.n258 585
R233 B.n257 B.n256 585
R234 B.n255 B.n254 585
R235 B.n253 B.n252 585
R236 B.n250 B.n249 585
R237 B.n248 B.n247 585
R238 B.n246 B.n245 585
R239 B.n244 B.n243 585
R240 B.n242 B.n241 585
R241 B.n240 B.n239 585
R242 B.n238 B.n237 585
R243 B.n236 B.n235 585
R244 B.n234 B.n233 585
R245 B.n232 B.n231 585
R246 B.n230 B.n229 585
R247 B.n228 B.n227 585
R248 B.n226 B.n225 585
R249 B.n224 B.n223 585
R250 B.n222 B.n221 585
R251 B.n220 B.n219 585
R252 B.n218 B.n217 585
R253 B.n216 B.n215 585
R254 B.n214 B.n213 585
R255 B.n212 B.n211 585
R256 B.n210 B.n209 585
R257 B.n208 B.n207 585
R258 B.n206 B.n205 585
R259 B.n204 B.n203 585
R260 B.n202 B.n201 585
R261 B.n200 B.n199 585
R262 B.n198 B.n197 585
R263 B.n196 B.n195 585
R264 B.n194 B.n193 585
R265 B.n192 B.n191 585
R266 B.n190 B.n189 585
R267 B.n188 B.n187 585
R268 B.n186 B.n185 585
R269 B.n184 B.n183 585
R270 B.n182 B.n181 585
R271 B.n180 B.n179 585
R272 B.n178 B.n177 585
R273 B.n176 B.n175 585
R274 B.n174 B.n173 585
R275 B.n172 B.n171 585
R276 B.n170 B.n169 585
R277 B.n168 B.n167 585
R278 B.n166 B.n165 585
R279 B.n164 B.n163 585
R280 B.n162 B.n161 585
R281 B.n103 B.n102 585
R282 B.n973 B.n972 585
R283 B.n967 B.n155 585
R284 B.n155 B.n100 585
R285 B.n966 B.n99 585
R286 B.n977 B.n99 585
R287 B.n965 B.n98 585
R288 B.n978 B.n98 585
R289 B.n964 B.n97 585
R290 B.n979 B.n97 585
R291 B.n963 B.n962 585
R292 B.n962 B.n93 585
R293 B.n961 B.n92 585
R294 B.n985 B.n92 585
R295 B.n960 B.n91 585
R296 B.n986 B.n91 585
R297 B.n959 B.n90 585
R298 B.n987 B.n90 585
R299 B.n958 B.n957 585
R300 B.n957 B.n86 585
R301 B.n956 B.n85 585
R302 B.n993 B.n85 585
R303 B.n955 B.n84 585
R304 B.n994 B.n84 585
R305 B.n954 B.n83 585
R306 B.n995 B.n83 585
R307 B.n953 B.n952 585
R308 B.n952 B.n79 585
R309 B.n951 B.n78 585
R310 B.n1001 B.n78 585
R311 B.n950 B.n77 585
R312 B.n1002 B.n77 585
R313 B.n949 B.n76 585
R314 B.n1003 B.n76 585
R315 B.n948 B.n947 585
R316 B.n947 B.n72 585
R317 B.n946 B.n71 585
R318 B.n1009 B.n71 585
R319 B.n945 B.n70 585
R320 B.n1010 B.n70 585
R321 B.n944 B.n69 585
R322 B.n1011 B.n69 585
R323 B.n943 B.n942 585
R324 B.n942 B.n65 585
R325 B.n941 B.n64 585
R326 B.n1017 B.n64 585
R327 B.n940 B.n63 585
R328 B.n1018 B.n63 585
R329 B.n939 B.n62 585
R330 B.n1019 B.n62 585
R331 B.n938 B.n937 585
R332 B.n937 B.n58 585
R333 B.n936 B.n57 585
R334 B.n1025 B.n57 585
R335 B.n935 B.n56 585
R336 B.n1026 B.n56 585
R337 B.n934 B.n55 585
R338 B.n1027 B.n55 585
R339 B.n933 B.n932 585
R340 B.n932 B.n51 585
R341 B.n931 B.n50 585
R342 B.n1033 B.n50 585
R343 B.n930 B.n49 585
R344 B.n1034 B.n49 585
R345 B.n929 B.n48 585
R346 B.n1035 B.n48 585
R347 B.n928 B.n927 585
R348 B.n927 B.n44 585
R349 B.n926 B.n43 585
R350 B.n1041 B.n43 585
R351 B.n925 B.n42 585
R352 B.n1042 B.n42 585
R353 B.n924 B.n41 585
R354 B.n1043 B.n41 585
R355 B.n923 B.n922 585
R356 B.n922 B.n37 585
R357 B.n921 B.n36 585
R358 B.n1049 B.n36 585
R359 B.n920 B.n35 585
R360 B.n1050 B.n35 585
R361 B.n919 B.n34 585
R362 B.n1051 B.n34 585
R363 B.n918 B.n917 585
R364 B.n917 B.n30 585
R365 B.n916 B.n29 585
R366 B.n1057 B.n29 585
R367 B.n915 B.n28 585
R368 B.n1058 B.n28 585
R369 B.n914 B.n27 585
R370 B.n1059 B.n27 585
R371 B.n913 B.n912 585
R372 B.n912 B.n23 585
R373 B.n911 B.n22 585
R374 B.n1065 B.n22 585
R375 B.n910 B.n21 585
R376 B.n1066 B.n21 585
R377 B.n909 B.n20 585
R378 B.n1067 B.n20 585
R379 B.n908 B.n907 585
R380 B.n907 B.n16 585
R381 B.n906 B.n15 585
R382 B.n1073 B.n15 585
R383 B.n905 B.n14 585
R384 B.n1074 B.n14 585
R385 B.n904 B.n13 585
R386 B.n1075 B.n13 585
R387 B.n903 B.n902 585
R388 B.n902 B.n12 585
R389 B.n901 B.n900 585
R390 B.n901 B.n8 585
R391 B.n899 B.n7 585
R392 B.n1082 B.n7 585
R393 B.n898 B.n6 585
R394 B.n1083 B.n6 585
R395 B.n897 B.n5 585
R396 B.n1084 B.n5 585
R397 B.n896 B.n895 585
R398 B.n895 B.n4 585
R399 B.n894 B.n361 585
R400 B.n894 B.n893 585
R401 B.n884 B.n362 585
R402 B.n363 B.n362 585
R403 B.n886 B.n885 585
R404 B.n887 B.n886 585
R405 B.n883 B.n368 585
R406 B.n368 B.n367 585
R407 B.n882 B.n881 585
R408 B.n881 B.n880 585
R409 B.n370 B.n369 585
R410 B.n371 B.n370 585
R411 B.n873 B.n872 585
R412 B.n874 B.n873 585
R413 B.n871 B.n376 585
R414 B.n376 B.n375 585
R415 B.n870 B.n869 585
R416 B.n869 B.n868 585
R417 B.n378 B.n377 585
R418 B.n379 B.n378 585
R419 B.n861 B.n860 585
R420 B.n862 B.n861 585
R421 B.n859 B.n384 585
R422 B.n384 B.n383 585
R423 B.n858 B.n857 585
R424 B.n857 B.n856 585
R425 B.n386 B.n385 585
R426 B.n387 B.n386 585
R427 B.n849 B.n848 585
R428 B.n850 B.n849 585
R429 B.n847 B.n392 585
R430 B.n392 B.n391 585
R431 B.n846 B.n845 585
R432 B.n845 B.n844 585
R433 B.n394 B.n393 585
R434 B.n395 B.n394 585
R435 B.n837 B.n836 585
R436 B.n838 B.n837 585
R437 B.n835 B.n399 585
R438 B.n403 B.n399 585
R439 B.n834 B.n833 585
R440 B.n833 B.n832 585
R441 B.n401 B.n400 585
R442 B.n402 B.n401 585
R443 B.n825 B.n824 585
R444 B.n826 B.n825 585
R445 B.n823 B.n408 585
R446 B.n408 B.n407 585
R447 B.n822 B.n821 585
R448 B.n821 B.n820 585
R449 B.n410 B.n409 585
R450 B.n411 B.n410 585
R451 B.n813 B.n812 585
R452 B.n814 B.n813 585
R453 B.n811 B.n415 585
R454 B.n419 B.n415 585
R455 B.n810 B.n809 585
R456 B.n809 B.n808 585
R457 B.n417 B.n416 585
R458 B.n418 B.n417 585
R459 B.n801 B.n800 585
R460 B.n802 B.n801 585
R461 B.n799 B.n424 585
R462 B.n424 B.n423 585
R463 B.n798 B.n797 585
R464 B.n797 B.n796 585
R465 B.n426 B.n425 585
R466 B.n427 B.n426 585
R467 B.n789 B.n788 585
R468 B.n790 B.n789 585
R469 B.n787 B.n431 585
R470 B.n435 B.n431 585
R471 B.n786 B.n785 585
R472 B.n785 B.n784 585
R473 B.n433 B.n432 585
R474 B.n434 B.n433 585
R475 B.n777 B.n776 585
R476 B.n778 B.n777 585
R477 B.n775 B.n440 585
R478 B.n440 B.n439 585
R479 B.n774 B.n773 585
R480 B.n773 B.n772 585
R481 B.n442 B.n441 585
R482 B.n443 B.n442 585
R483 B.n765 B.n764 585
R484 B.n766 B.n765 585
R485 B.n763 B.n448 585
R486 B.n448 B.n447 585
R487 B.n762 B.n761 585
R488 B.n761 B.n760 585
R489 B.n450 B.n449 585
R490 B.n451 B.n450 585
R491 B.n753 B.n752 585
R492 B.n754 B.n753 585
R493 B.n751 B.n456 585
R494 B.n456 B.n455 585
R495 B.n750 B.n749 585
R496 B.n749 B.n748 585
R497 B.n458 B.n457 585
R498 B.n459 B.n458 585
R499 B.n741 B.n740 585
R500 B.n742 B.n741 585
R501 B.n739 B.n464 585
R502 B.n464 B.n463 585
R503 B.n738 B.n737 585
R504 B.n737 B.n736 585
R505 B.n466 B.n465 585
R506 B.n467 B.n466 585
R507 B.n732 B.n731 585
R508 B.n470 B.n469 585
R509 B.n728 B.n727 585
R510 B.n729 B.n728 585
R511 B.n726 B.n521 585
R512 B.n725 B.n724 585
R513 B.n723 B.n722 585
R514 B.n721 B.n720 585
R515 B.n719 B.n718 585
R516 B.n717 B.n716 585
R517 B.n715 B.n714 585
R518 B.n713 B.n712 585
R519 B.n711 B.n710 585
R520 B.n709 B.n708 585
R521 B.n707 B.n706 585
R522 B.n705 B.n704 585
R523 B.n703 B.n702 585
R524 B.n701 B.n700 585
R525 B.n699 B.n698 585
R526 B.n697 B.n696 585
R527 B.n695 B.n694 585
R528 B.n693 B.n692 585
R529 B.n691 B.n690 585
R530 B.n689 B.n688 585
R531 B.n687 B.n686 585
R532 B.n685 B.n684 585
R533 B.n683 B.n682 585
R534 B.n681 B.n680 585
R535 B.n679 B.n678 585
R536 B.n677 B.n676 585
R537 B.n675 B.n674 585
R538 B.n673 B.n672 585
R539 B.n671 B.n670 585
R540 B.n669 B.n668 585
R541 B.n667 B.n666 585
R542 B.n665 B.n664 585
R543 B.n663 B.n662 585
R544 B.n661 B.n660 585
R545 B.n659 B.n658 585
R546 B.n657 B.n656 585
R547 B.n655 B.n654 585
R548 B.n653 B.n652 585
R549 B.n651 B.n650 585
R550 B.n649 B.n648 585
R551 B.n647 B.n646 585
R552 B.n645 B.n644 585
R553 B.n643 B.n642 585
R554 B.n641 B.n640 585
R555 B.n639 B.n638 585
R556 B.n637 B.n636 585
R557 B.n635 B.n634 585
R558 B.n633 B.n632 585
R559 B.n631 B.n630 585
R560 B.n629 B.n628 585
R561 B.n627 B.n626 585
R562 B.n625 B.n624 585
R563 B.n623 B.n622 585
R564 B.n620 B.n619 585
R565 B.n618 B.n617 585
R566 B.n616 B.n615 585
R567 B.n614 B.n613 585
R568 B.n612 B.n611 585
R569 B.n610 B.n609 585
R570 B.n608 B.n607 585
R571 B.n606 B.n605 585
R572 B.n604 B.n603 585
R573 B.n602 B.n601 585
R574 B.n600 B.n599 585
R575 B.n598 B.n597 585
R576 B.n596 B.n595 585
R577 B.n594 B.n593 585
R578 B.n592 B.n591 585
R579 B.n590 B.n589 585
R580 B.n588 B.n587 585
R581 B.n586 B.n585 585
R582 B.n584 B.n583 585
R583 B.n582 B.n581 585
R584 B.n580 B.n579 585
R585 B.n578 B.n577 585
R586 B.n576 B.n575 585
R587 B.n574 B.n573 585
R588 B.n572 B.n571 585
R589 B.n570 B.n569 585
R590 B.n568 B.n567 585
R591 B.n566 B.n565 585
R592 B.n564 B.n563 585
R593 B.n562 B.n561 585
R594 B.n560 B.n559 585
R595 B.n558 B.n557 585
R596 B.n556 B.n555 585
R597 B.n554 B.n553 585
R598 B.n552 B.n551 585
R599 B.n550 B.n549 585
R600 B.n548 B.n547 585
R601 B.n546 B.n545 585
R602 B.n544 B.n543 585
R603 B.n542 B.n541 585
R604 B.n540 B.n539 585
R605 B.n538 B.n537 585
R606 B.n536 B.n535 585
R607 B.n534 B.n533 585
R608 B.n532 B.n531 585
R609 B.n530 B.n529 585
R610 B.n528 B.n527 585
R611 B.n733 B.n468 585
R612 B.n468 B.n467 585
R613 B.n735 B.n734 585
R614 B.n736 B.n735 585
R615 B.n462 B.n461 585
R616 B.n463 B.n462 585
R617 B.n744 B.n743 585
R618 B.n743 B.n742 585
R619 B.n745 B.n460 585
R620 B.n460 B.n459 585
R621 B.n747 B.n746 585
R622 B.n748 B.n747 585
R623 B.n454 B.n453 585
R624 B.n455 B.n454 585
R625 B.n756 B.n755 585
R626 B.n755 B.n754 585
R627 B.n757 B.n452 585
R628 B.n452 B.n451 585
R629 B.n759 B.n758 585
R630 B.n760 B.n759 585
R631 B.n446 B.n445 585
R632 B.n447 B.n446 585
R633 B.n768 B.n767 585
R634 B.n767 B.n766 585
R635 B.n769 B.n444 585
R636 B.n444 B.n443 585
R637 B.n771 B.n770 585
R638 B.n772 B.n771 585
R639 B.n438 B.n437 585
R640 B.n439 B.n438 585
R641 B.n780 B.n779 585
R642 B.n779 B.n778 585
R643 B.n781 B.n436 585
R644 B.n436 B.n434 585
R645 B.n783 B.n782 585
R646 B.n784 B.n783 585
R647 B.n430 B.n429 585
R648 B.n435 B.n430 585
R649 B.n792 B.n791 585
R650 B.n791 B.n790 585
R651 B.n793 B.n428 585
R652 B.n428 B.n427 585
R653 B.n795 B.n794 585
R654 B.n796 B.n795 585
R655 B.n422 B.n421 585
R656 B.n423 B.n422 585
R657 B.n804 B.n803 585
R658 B.n803 B.n802 585
R659 B.n805 B.n420 585
R660 B.n420 B.n418 585
R661 B.n807 B.n806 585
R662 B.n808 B.n807 585
R663 B.n414 B.n413 585
R664 B.n419 B.n414 585
R665 B.n816 B.n815 585
R666 B.n815 B.n814 585
R667 B.n817 B.n412 585
R668 B.n412 B.n411 585
R669 B.n819 B.n818 585
R670 B.n820 B.n819 585
R671 B.n406 B.n405 585
R672 B.n407 B.n406 585
R673 B.n828 B.n827 585
R674 B.n827 B.n826 585
R675 B.n829 B.n404 585
R676 B.n404 B.n402 585
R677 B.n831 B.n830 585
R678 B.n832 B.n831 585
R679 B.n398 B.n397 585
R680 B.n403 B.n398 585
R681 B.n840 B.n839 585
R682 B.n839 B.n838 585
R683 B.n841 B.n396 585
R684 B.n396 B.n395 585
R685 B.n843 B.n842 585
R686 B.n844 B.n843 585
R687 B.n390 B.n389 585
R688 B.n391 B.n390 585
R689 B.n852 B.n851 585
R690 B.n851 B.n850 585
R691 B.n853 B.n388 585
R692 B.n388 B.n387 585
R693 B.n855 B.n854 585
R694 B.n856 B.n855 585
R695 B.n382 B.n381 585
R696 B.n383 B.n382 585
R697 B.n864 B.n863 585
R698 B.n863 B.n862 585
R699 B.n865 B.n380 585
R700 B.n380 B.n379 585
R701 B.n867 B.n866 585
R702 B.n868 B.n867 585
R703 B.n374 B.n373 585
R704 B.n375 B.n374 585
R705 B.n876 B.n875 585
R706 B.n875 B.n874 585
R707 B.n877 B.n372 585
R708 B.n372 B.n371 585
R709 B.n879 B.n878 585
R710 B.n880 B.n879 585
R711 B.n366 B.n365 585
R712 B.n367 B.n366 585
R713 B.n889 B.n888 585
R714 B.n888 B.n887 585
R715 B.n890 B.n364 585
R716 B.n364 B.n363 585
R717 B.n892 B.n891 585
R718 B.n893 B.n892 585
R719 B.n3 B.n0 585
R720 B.n4 B.n3 585
R721 B.n1081 B.n1 585
R722 B.n1082 B.n1081 585
R723 B.n1080 B.n1079 585
R724 B.n1080 B.n8 585
R725 B.n1078 B.n9 585
R726 B.n12 B.n9 585
R727 B.n1077 B.n1076 585
R728 B.n1076 B.n1075 585
R729 B.n11 B.n10 585
R730 B.n1074 B.n11 585
R731 B.n1072 B.n1071 585
R732 B.n1073 B.n1072 585
R733 B.n1070 B.n17 585
R734 B.n17 B.n16 585
R735 B.n1069 B.n1068 585
R736 B.n1068 B.n1067 585
R737 B.n19 B.n18 585
R738 B.n1066 B.n19 585
R739 B.n1064 B.n1063 585
R740 B.n1065 B.n1064 585
R741 B.n1062 B.n24 585
R742 B.n24 B.n23 585
R743 B.n1061 B.n1060 585
R744 B.n1060 B.n1059 585
R745 B.n26 B.n25 585
R746 B.n1058 B.n26 585
R747 B.n1056 B.n1055 585
R748 B.n1057 B.n1056 585
R749 B.n1054 B.n31 585
R750 B.n31 B.n30 585
R751 B.n1053 B.n1052 585
R752 B.n1052 B.n1051 585
R753 B.n33 B.n32 585
R754 B.n1050 B.n33 585
R755 B.n1048 B.n1047 585
R756 B.n1049 B.n1048 585
R757 B.n1046 B.n38 585
R758 B.n38 B.n37 585
R759 B.n1045 B.n1044 585
R760 B.n1044 B.n1043 585
R761 B.n40 B.n39 585
R762 B.n1042 B.n40 585
R763 B.n1040 B.n1039 585
R764 B.n1041 B.n1040 585
R765 B.n1038 B.n45 585
R766 B.n45 B.n44 585
R767 B.n1037 B.n1036 585
R768 B.n1036 B.n1035 585
R769 B.n47 B.n46 585
R770 B.n1034 B.n47 585
R771 B.n1032 B.n1031 585
R772 B.n1033 B.n1032 585
R773 B.n1030 B.n52 585
R774 B.n52 B.n51 585
R775 B.n1029 B.n1028 585
R776 B.n1028 B.n1027 585
R777 B.n54 B.n53 585
R778 B.n1026 B.n54 585
R779 B.n1024 B.n1023 585
R780 B.n1025 B.n1024 585
R781 B.n1022 B.n59 585
R782 B.n59 B.n58 585
R783 B.n1021 B.n1020 585
R784 B.n1020 B.n1019 585
R785 B.n61 B.n60 585
R786 B.n1018 B.n61 585
R787 B.n1016 B.n1015 585
R788 B.n1017 B.n1016 585
R789 B.n1014 B.n66 585
R790 B.n66 B.n65 585
R791 B.n1013 B.n1012 585
R792 B.n1012 B.n1011 585
R793 B.n68 B.n67 585
R794 B.n1010 B.n68 585
R795 B.n1008 B.n1007 585
R796 B.n1009 B.n1008 585
R797 B.n1006 B.n73 585
R798 B.n73 B.n72 585
R799 B.n1005 B.n1004 585
R800 B.n1004 B.n1003 585
R801 B.n75 B.n74 585
R802 B.n1002 B.n75 585
R803 B.n1000 B.n999 585
R804 B.n1001 B.n1000 585
R805 B.n998 B.n80 585
R806 B.n80 B.n79 585
R807 B.n997 B.n996 585
R808 B.n996 B.n995 585
R809 B.n82 B.n81 585
R810 B.n994 B.n82 585
R811 B.n992 B.n991 585
R812 B.n993 B.n992 585
R813 B.n990 B.n87 585
R814 B.n87 B.n86 585
R815 B.n989 B.n988 585
R816 B.n988 B.n987 585
R817 B.n89 B.n88 585
R818 B.n986 B.n89 585
R819 B.n984 B.n983 585
R820 B.n985 B.n984 585
R821 B.n982 B.n94 585
R822 B.n94 B.n93 585
R823 B.n981 B.n980 585
R824 B.n980 B.n979 585
R825 B.n96 B.n95 585
R826 B.n978 B.n96 585
R827 B.n976 B.n975 585
R828 B.n977 B.n976 585
R829 B.n974 B.n101 585
R830 B.n101 B.n100 585
R831 B.n1085 B.n1084 585
R832 B.n1083 B.n2 585
R833 B.n972 B.n101 564.573
R834 B.n969 B.n155 564.573
R835 B.n527 B.n466 564.573
R836 B.n731 B.n468 564.573
R837 B.n159 B.t17 347.798
R838 B.n156 B.t21 347.798
R839 B.n525 B.t14 347.798
R840 B.n522 B.t10 347.798
R841 B.n970 B.n153 256.663
R842 B.n970 B.n152 256.663
R843 B.n970 B.n151 256.663
R844 B.n970 B.n150 256.663
R845 B.n970 B.n149 256.663
R846 B.n970 B.n148 256.663
R847 B.n970 B.n147 256.663
R848 B.n970 B.n146 256.663
R849 B.n970 B.n145 256.663
R850 B.n970 B.n144 256.663
R851 B.n970 B.n143 256.663
R852 B.n970 B.n142 256.663
R853 B.n970 B.n141 256.663
R854 B.n970 B.n140 256.663
R855 B.n970 B.n139 256.663
R856 B.n970 B.n138 256.663
R857 B.n970 B.n137 256.663
R858 B.n970 B.n136 256.663
R859 B.n970 B.n135 256.663
R860 B.n970 B.n134 256.663
R861 B.n970 B.n133 256.663
R862 B.n970 B.n132 256.663
R863 B.n970 B.n131 256.663
R864 B.n970 B.n130 256.663
R865 B.n970 B.n129 256.663
R866 B.n970 B.n128 256.663
R867 B.n970 B.n127 256.663
R868 B.n970 B.n126 256.663
R869 B.n970 B.n125 256.663
R870 B.n970 B.n124 256.663
R871 B.n970 B.n123 256.663
R872 B.n970 B.n122 256.663
R873 B.n970 B.n121 256.663
R874 B.n970 B.n120 256.663
R875 B.n970 B.n119 256.663
R876 B.n970 B.n118 256.663
R877 B.n970 B.n117 256.663
R878 B.n970 B.n116 256.663
R879 B.n970 B.n115 256.663
R880 B.n970 B.n114 256.663
R881 B.n970 B.n113 256.663
R882 B.n970 B.n112 256.663
R883 B.n970 B.n111 256.663
R884 B.n970 B.n110 256.663
R885 B.n970 B.n109 256.663
R886 B.n970 B.n108 256.663
R887 B.n970 B.n107 256.663
R888 B.n970 B.n106 256.663
R889 B.n970 B.n105 256.663
R890 B.n970 B.n104 256.663
R891 B.n971 B.n970 256.663
R892 B.n730 B.n729 256.663
R893 B.n729 B.n471 256.663
R894 B.n729 B.n472 256.663
R895 B.n729 B.n473 256.663
R896 B.n729 B.n474 256.663
R897 B.n729 B.n475 256.663
R898 B.n729 B.n476 256.663
R899 B.n729 B.n477 256.663
R900 B.n729 B.n478 256.663
R901 B.n729 B.n479 256.663
R902 B.n729 B.n480 256.663
R903 B.n729 B.n481 256.663
R904 B.n729 B.n482 256.663
R905 B.n729 B.n483 256.663
R906 B.n729 B.n484 256.663
R907 B.n729 B.n485 256.663
R908 B.n729 B.n486 256.663
R909 B.n729 B.n487 256.663
R910 B.n729 B.n488 256.663
R911 B.n729 B.n489 256.663
R912 B.n729 B.n490 256.663
R913 B.n729 B.n491 256.663
R914 B.n729 B.n492 256.663
R915 B.n729 B.n493 256.663
R916 B.n729 B.n494 256.663
R917 B.n729 B.n495 256.663
R918 B.n729 B.n496 256.663
R919 B.n729 B.n497 256.663
R920 B.n729 B.n498 256.663
R921 B.n729 B.n499 256.663
R922 B.n729 B.n500 256.663
R923 B.n729 B.n501 256.663
R924 B.n729 B.n502 256.663
R925 B.n729 B.n503 256.663
R926 B.n729 B.n504 256.663
R927 B.n729 B.n505 256.663
R928 B.n729 B.n506 256.663
R929 B.n729 B.n507 256.663
R930 B.n729 B.n508 256.663
R931 B.n729 B.n509 256.663
R932 B.n729 B.n510 256.663
R933 B.n729 B.n511 256.663
R934 B.n729 B.n512 256.663
R935 B.n729 B.n513 256.663
R936 B.n729 B.n514 256.663
R937 B.n729 B.n515 256.663
R938 B.n729 B.n516 256.663
R939 B.n729 B.n517 256.663
R940 B.n729 B.n518 256.663
R941 B.n729 B.n519 256.663
R942 B.n729 B.n520 256.663
R943 B.n1087 B.n1086 256.663
R944 B.n161 B.n103 163.367
R945 B.n165 B.n164 163.367
R946 B.n169 B.n168 163.367
R947 B.n173 B.n172 163.367
R948 B.n177 B.n176 163.367
R949 B.n181 B.n180 163.367
R950 B.n185 B.n184 163.367
R951 B.n189 B.n188 163.367
R952 B.n193 B.n192 163.367
R953 B.n197 B.n196 163.367
R954 B.n201 B.n200 163.367
R955 B.n205 B.n204 163.367
R956 B.n209 B.n208 163.367
R957 B.n213 B.n212 163.367
R958 B.n217 B.n216 163.367
R959 B.n221 B.n220 163.367
R960 B.n225 B.n224 163.367
R961 B.n229 B.n228 163.367
R962 B.n233 B.n232 163.367
R963 B.n237 B.n236 163.367
R964 B.n241 B.n240 163.367
R965 B.n245 B.n244 163.367
R966 B.n249 B.n248 163.367
R967 B.n254 B.n253 163.367
R968 B.n258 B.n257 163.367
R969 B.n262 B.n261 163.367
R970 B.n266 B.n265 163.367
R971 B.n270 B.n269 163.367
R972 B.n274 B.n273 163.367
R973 B.n278 B.n277 163.367
R974 B.n282 B.n281 163.367
R975 B.n286 B.n285 163.367
R976 B.n290 B.n289 163.367
R977 B.n294 B.n293 163.367
R978 B.n298 B.n297 163.367
R979 B.n302 B.n301 163.367
R980 B.n306 B.n305 163.367
R981 B.n310 B.n309 163.367
R982 B.n314 B.n313 163.367
R983 B.n318 B.n317 163.367
R984 B.n322 B.n321 163.367
R985 B.n326 B.n325 163.367
R986 B.n330 B.n329 163.367
R987 B.n334 B.n333 163.367
R988 B.n338 B.n337 163.367
R989 B.n342 B.n341 163.367
R990 B.n346 B.n345 163.367
R991 B.n350 B.n349 163.367
R992 B.n354 B.n353 163.367
R993 B.n358 B.n357 163.367
R994 B.n969 B.n154 163.367
R995 B.n737 B.n466 163.367
R996 B.n737 B.n464 163.367
R997 B.n741 B.n464 163.367
R998 B.n741 B.n458 163.367
R999 B.n749 B.n458 163.367
R1000 B.n749 B.n456 163.367
R1001 B.n753 B.n456 163.367
R1002 B.n753 B.n450 163.367
R1003 B.n761 B.n450 163.367
R1004 B.n761 B.n448 163.367
R1005 B.n765 B.n448 163.367
R1006 B.n765 B.n442 163.367
R1007 B.n773 B.n442 163.367
R1008 B.n773 B.n440 163.367
R1009 B.n777 B.n440 163.367
R1010 B.n777 B.n433 163.367
R1011 B.n785 B.n433 163.367
R1012 B.n785 B.n431 163.367
R1013 B.n789 B.n431 163.367
R1014 B.n789 B.n426 163.367
R1015 B.n797 B.n426 163.367
R1016 B.n797 B.n424 163.367
R1017 B.n801 B.n424 163.367
R1018 B.n801 B.n417 163.367
R1019 B.n809 B.n417 163.367
R1020 B.n809 B.n415 163.367
R1021 B.n813 B.n415 163.367
R1022 B.n813 B.n410 163.367
R1023 B.n821 B.n410 163.367
R1024 B.n821 B.n408 163.367
R1025 B.n825 B.n408 163.367
R1026 B.n825 B.n401 163.367
R1027 B.n833 B.n401 163.367
R1028 B.n833 B.n399 163.367
R1029 B.n837 B.n399 163.367
R1030 B.n837 B.n394 163.367
R1031 B.n845 B.n394 163.367
R1032 B.n845 B.n392 163.367
R1033 B.n849 B.n392 163.367
R1034 B.n849 B.n386 163.367
R1035 B.n857 B.n386 163.367
R1036 B.n857 B.n384 163.367
R1037 B.n861 B.n384 163.367
R1038 B.n861 B.n378 163.367
R1039 B.n869 B.n378 163.367
R1040 B.n869 B.n376 163.367
R1041 B.n873 B.n376 163.367
R1042 B.n873 B.n370 163.367
R1043 B.n881 B.n370 163.367
R1044 B.n881 B.n368 163.367
R1045 B.n886 B.n368 163.367
R1046 B.n886 B.n362 163.367
R1047 B.n894 B.n362 163.367
R1048 B.n895 B.n894 163.367
R1049 B.n895 B.n5 163.367
R1050 B.n6 B.n5 163.367
R1051 B.n7 B.n6 163.367
R1052 B.n901 B.n7 163.367
R1053 B.n902 B.n901 163.367
R1054 B.n902 B.n13 163.367
R1055 B.n14 B.n13 163.367
R1056 B.n15 B.n14 163.367
R1057 B.n907 B.n15 163.367
R1058 B.n907 B.n20 163.367
R1059 B.n21 B.n20 163.367
R1060 B.n22 B.n21 163.367
R1061 B.n912 B.n22 163.367
R1062 B.n912 B.n27 163.367
R1063 B.n28 B.n27 163.367
R1064 B.n29 B.n28 163.367
R1065 B.n917 B.n29 163.367
R1066 B.n917 B.n34 163.367
R1067 B.n35 B.n34 163.367
R1068 B.n36 B.n35 163.367
R1069 B.n922 B.n36 163.367
R1070 B.n922 B.n41 163.367
R1071 B.n42 B.n41 163.367
R1072 B.n43 B.n42 163.367
R1073 B.n927 B.n43 163.367
R1074 B.n927 B.n48 163.367
R1075 B.n49 B.n48 163.367
R1076 B.n50 B.n49 163.367
R1077 B.n932 B.n50 163.367
R1078 B.n932 B.n55 163.367
R1079 B.n56 B.n55 163.367
R1080 B.n57 B.n56 163.367
R1081 B.n937 B.n57 163.367
R1082 B.n937 B.n62 163.367
R1083 B.n63 B.n62 163.367
R1084 B.n64 B.n63 163.367
R1085 B.n942 B.n64 163.367
R1086 B.n942 B.n69 163.367
R1087 B.n70 B.n69 163.367
R1088 B.n71 B.n70 163.367
R1089 B.n947 B.n71 163.367
R1090 B.n947 B.n76 163.367
R1091 B.n77 B.n76 163.367
R1092 B.n78 B.n77 163.367
R1093 B.n952 B.n78 163.367
R1094 B.n952 B.n83 163.367
R1095 B.n84 B.n83 163.367
R1096 B.n85 B.n84 163.367
R1097 B.n957 B.n85 163.367
R1098 B.n957 B.n90 163.367
R1099 B.n91 B.n90 163.367
R1100 B.n92 B.n91 163.367
R1101 B.n962 B.n92 163.367
R1102 B.n962 B.n97 163.367
R1103 B.n98 B.n97 163.367
R1104 B.n99 B.n98 163.367
R1105 B.n155 B.n99 163.367
R1106 B.n728 B.n470 163.367
R1107 B.n728 B.n521 163.367
R1108 B.n724 B.n723 163.367
R1109 B.n720 B.n719 163.367
R1110 B.n716 B.n715 163.367
R1111 B.n712 B.n711 163.367
R1112 B.n708 B.n707 163.367
R1113 B.n704 B.n703 163.367
R1114 B.n700 B.n699 163.367
R1115 B.n696 B.n695 163.367
R1116 B.n692 B.n691 163.367
R1117 B.n688 B.n687 163.367
R1118 B.n684 B.n683 163.367
R1119 B.n680 B.n679 163.367
R1120 B.n676 B.n675 163.367
R1121 B.n672 B.n671 163.367
R1122 B.n668 B.n667 163.367
R1123 B.n664 B.n663 163.367
R1124 B.n660 B.n659 163.367
R1125 B.n656 B.n655 163.367
R1126 B.n652 B.n651 163.367
R1127 B.n648 B.n647 163.367
R1128 B.n644 B.n643 163.367
R1129 B.n640 B.n639 163.367
R1130 B.n636 B.n635 163.367
R1131 B.n632 B.n631 163.367
R1132 B.n628 B.n627 163.367
R1133 B.n624 B.n623 163.367
R1134 B.n619 B.n618 163.367
R1135 B.n615 B.n614 163.367
R1136 B.n611 B.n610 163.367
R1137 B.n607 B.n606 163.367
R1138 B.n603 B.n602 163.367
R1139 B.n599 B.n598 163.367
R1140 B.n595 B.n594 163.367
R1141 B.n591 B.n590 163.367
R1142 B.n587 B.n586 163.367
R1143 B.n583 B.n582 163.367
R1144 B.n579 B.n578 163.367
R1145 B.n575 B.n574 163.367
R1146 B.n571 B.n570 163.367
R1147 B.n567 B.n566 163.367
R1148 B.n563 B.n562 163.367
R1149 B.n559 B.n558 163.367
R1150 B.n555 B.n554 163.367
R1151 B.n551 B.n550 163.367
R1152 B.n547 B.n546 163.367
R1153 B.n543 B.n542 163.367
R1154 B.n539 B.n538 163.367
R1155 B.n535 B.n534 163.367
R1156 B.n531 B.n530 163.367
R1157 B.n735 B.n468 163.367
R1158 B.n735 B.n462 163.367
R1159 B.n743 B.n462 163.367
R1160 B.n743 B.n460 163.367
R1161 B.n747 B.n460 163.367
R1162 B.n747 B.n454 163.367
R1163 B.n755 B.n454 163.367
R1164 B.n755 B.n452 163.367
R1165 B.n759 B.n452 163.367
R1166 B.n759 B.n446 163.367
R1167 B.n767 B.n446 163.367
R1168 B.n767 B.n444 163.367
R1169 B.n771 B.n444 163.367
R1170 B.n771 B.n438 163.367
R1171 B.n779 B.n438 163.367
R1172 B.n779 B.n436 163.367
R1173 B.n783 B.n436 163.367
R1174 B.n783 B.n430 163.367
R1175 B.n791 B.n430 163.367
R1176 B.n791 B.n428 163.367
R1177 B.n795 B.n428 163.367
R1178 B.n795 B.n422 163.367
R1179 B.n803 B.n422 163.367
R1180 B.n803 B.n420 163.367
R1181 B.n807 B.n420 163.367
R1182 B.n807 B.n414 163.367
R1183 B.n815 B.n414 163.367
R1184 B.n815 B.n412 163.367
R1185 B.n819 B.n412 163.367
R1186 B.n819 B.n406 163.367
R1187 B.n827 B.n406 163.367
R1188 B.n827 B.n404 163.367
R1189 B.n831 B.n404 163.367
R1190 B.n831 B.n398 163.367
R1191 B.n839 B.n398 163.367
R1192 B.n839 B.n396 163.367
R1193 B.n843 B.n396 163.367
R1194 B.n843 B.n390 163.367
R1195 B.n851 B.n390 163.367
R1196 B.n851 B.n388 163.367
R1197 B.n855 B.n388 163.367
R1198 B.n855 B.n382 163.367
R1199 B.n863 B.n382 163.367
R1200 B.n863 B.n380 163.367
R1201 B.n867 B.n380 163.367
R1202 B.n867 B.n374 163.367
R1203 B.n875 B.n374 163.367
R1204 B.n875 B.n372 163.367
R1205 B.n879 B.n372 163.367
R1206 B.n879 B.n366 163.367
R1207 B.n888 B.n366 163.367
R1208 B.n888 B.n364 163.367
R1209 B.n892 B.n364 163.367
R1210 B.n892 B.n3 163.367
R1211 B.n1085 B.n3 163.367
R1212 B.n1081 B.n2 163.367
R1213 B.n1081 B.n1080 163.367
R1214 B.n1080 B.n9 163.367
R1215 B.n1076 B.n9 163.367
R1216 B.n1076 B.n11 163.367
R1217 B.n1072 B.n11 163.367
R1218 B.n1072 B.n17 163.367
R1219 B.n1068 B.n17 163.367
R1220 B.n1068 B.n19 163.367
R1221 B.n1064 B.n19 163.367
R1222 B.n1064 B.n24 163.367
R1223 B.n1060 B.n24 163.367
R1224 B.n1060 B.n26 163.367
R1225 B.n1056 B.n26 163.367
R1226 B.n1056 B.n31 163.367
R1227 B.n1052 B.n31 163.367
R1228 B.n1052 B.n33 163.367
R1229 B.n1048 B.n33 163.367
R1230 B.n1048 B.n38 163.367
R1231 B.n1044 B.n38 163.367
R1232 B.n1044 B.n40 163.367
R1233 B.n1040 B.n40 163.367
R1234 B.n1040 B.n45 163.367
R1235 B.n1036 B.n45 163.367
R1236 B.n1036 B.n47 163.367
R1237 B.n1032 B.n47 163.367
R1238 B.n1032 B.n52 163.367
R1239 B.n1028 B.n52 163.367
R1240 B.n1028 B.n54 163.367
R1241 B.n1024 B.n54 163.367
R1242 B.n1024 B.n59 163.367
R1243 B.n1020 B.n59 163.367
R1244 B.n1020 B.n61 163.367
R1245 B.n1016 B.n61 163.367
R1246 B.n1016 B.n66 163.367
R1247 B.n1012 B.n66 163.367
R1248 B.n1012 B.n68 163.367
R1249 B.n1008 B.n68 163.367
R1250 B.n1008 B.n73 163.367
R1251 B.n1004 B.n73 163.367
R1252 B.n1004 B.n75 163.367
R1253 B.n1000 B.n75 163.367
R1254 B.n1000 B.n80 163.367
R1255 B.n996 B.n80 163.367
R1256 B.n996 B.n82 163.367
R1257 B.n992 B.n82 163.367
R1258 B.n992 B.n87 163.367
R1259 B.n988 B.n87 163.367
R1260 B.n988 B.n89 163.367
R1261 B.n984 B.n89 163.367
R1262 B.n984 B.n94 163.367
R1263 B.n980 B.n94 163.367
R1264 B.n980 B.n96 163.367
R1265 B.n976 B.n96 163.367
R1266 B.n976 B.n101 163.367
R1267 B.n156 B.t22 123.433
R1268 B.n525 B.t16 123.433
R1269 B.n159 B.t19 123.416
R1270 B.n522 B.t13 123.416
R1271 B.n729 B.n467 81.3965
R1272 B.n970 B.n100 81.3965
R1273 B.n972 B.n971 71.676
R1274 B.n161 B.n104 71.676
R1275 B.n165 B.n105 71.676
R1276 B.n169 B.n106 71.676
R1277 B.n173 B.n107 71.676
R1278 B.n177 B.n108 71.676
R1279 B.n181 B.n109 71.676
R1280 B.n185 B.n110 71.676
R1281 B.n189 B.n111 71.676
R1282 B.n193 B.n112 71.676
R1283 B.n197 B.n113 71.676
R1284 B.n201 B.n114 71.676
R1285 B.n205 B.n115 71.676
R1286 B.n209 B.n116 71.676
R1287 B.n213 B.n117 71.676
R1288 B.n217 B.n118 71.676
R1289 B.n221 B.n119 71.676
R1290 B.n225 B.n120 71.676
R1291 B.n229 B.n121 71.676
R1292 B.n233 B.n122 71.676
R1293 B.n237 B.n123 71.676
R1294 B.n241 B.n124 71.676
R1295 B.n245 B.n125 71.676
R1296 B.n249 B.n126 71.676
R1297 B.n254 B.n127 71.676
R1298 B.n258 B.n128 71.676
R1299 B.n262 B.n129 71.676
R1300 B.n266 B.n130 71.676
R1301 B.n270 B.n131 71.676
R1302 B.n274 B.n132 71.676
R1303 B.n278 B.n133 71.676
R1304 B.n282 B.n134 71.676
R1305 B.n286 B.n135 71.676
R1306 B.n290 B.n136 71.676
R1307 B.n294 B.n137 71.676
R1308 B.n298 B.n138 71.676
R1309 B.n302 B.n139 71.676
R1310 B.n306 B.n140 71.676
R1311 B.n310 B.n141 71.676
R1312 B.n314 B.n142 71.676
R1313 B.n318 B.n143 71.676
R1314 B.n322 B.n144 71.676
R1315 B.n326 B.n145 71.676
R1316 B.n330 B.n146 71.676
R1317 B.n334 B.n147 71.676
R1318 B.n338 B.n148 71.676
R1319 B.n342 B.n149 71.676
R1320 B.n346 B.n150 71.676
R1321 B.n350 B.n151 71.676
R1322 B.n354 B.n152 71.676
R1323 B.n358 B.n153 71.676
R1324 B.n154 B.n153 71.676
R1325 B.n357 B.n152 71.676
R1326 B.n353 B.n151 71.676
R1327 B.n349 B.n150 71.676
R1328 B.n345 B.n149 71.676
R1329 B.n341 B.n148 71.676
R1330 B.n337 B.n147 71.676
R1331 B.n333 B.n146 71.676
R1332 B.n329 B.n145 71.676
R1333 B.n325 B.n144 71.676
R1334 B.n321 B.n143 71.676
R1335 B.n317 B.n142 71.676
R1336 B.n313 B.n141 71.676
R1337 B.n309 B.n140 71.676
R1338 B.n305 B.n139 71.676
R1339 B.n301 B.n138 71.676
R1340 B.n297 B.n137 71.676
R1341 B.n293 B.n136 71.676
R1342 B.n289 B.n135 71.676
R1343 B.n285 B.n134 71.676
R1344 B.n281 B.n133 71.676
R1345 B.n277 B.n132 71.676
R1346 B.n273 B.n131 71.676
R1347 B.n269 B.n130 71.676
R1348 B.n265 B.n129 71.676
R1349 B.n261 B.n128 71.676
R1350 B.n257 B.n127 71.676
R1351 B.n253 B.n126 71.676
R1352 B.n248 B.n125 71.676
R1353 B.n244 B.n124 71.676
R1354 B.n240 B.n123 71.676
R1355 B.n236 B.n122 71.676
R1356 B.n232 B.n121 71.676
R1357 B.n228 B.n120 71.676
R1358 B.n224 B.n119 71.676
R1359 B.n220 B.n118 71.676
R1360 B.n216 B.n117 71.676
R1361 B.n212 B.n116 71.676
R1362 B.n208 B.n115 71.676
R1363 B.n204 B.n114 71.676
R1364 B.n200 B.n113 71.676
R1365 B.n196 B.n112 71.676
R1366 B.n192 B.n111 71.676
R1367 B.n188 B.n110 71.676
R1368 B.n184 B.n109 71.676
R1369 B.n180 B.n108 71.676
R1370 B.n176 B.n107 71.676
R1371 B.n172 B.n106 71.676
R1372 B.n168 B.n105 71.676
R1373 B.n164 B.n104 71.676
R1374 B.n971 B.n103 71.676
R1375 B.n731 B.n730 71.676
R1376 B.n521 B.n471 71.676
R1377 B.n723 B.n472 71.676
R1378 B.n719 B.n473 71.676
R1379 B.n715 B.n474 71.676
R1380 B.n711 B.n475 71.676
R1381 B.n707 B.n476 71.676
R1382 B.n703 B.n477 71.676
R1383 B.n699 B.n478 71.676
R1384 B.n695 B.n479 71.676
R1385 B.n691 B.n480 71.676
R1386 B.n687 B.n481 71.676
R1387 B.n683 B.n482 71.676
R1388 B.n679 B.n483 71.676
R1389 B.n675 B.n484 71.676
R1390 B.n671 B.n485 71.676
R1391 B.n667 B.n486 71.676
R1392 B.n663 B.n487 71.676
R1393 B.n659 B.n488 71.676
R1394 B.n655 B.n489 71.676
R1395 B.n651 B.n490 71.676
R1396 B.n647 B.n491 71.676
R1397 B.n643 B.n492 71.676
R1398 B.n639 B.n493 71.676
R1399 B.n635 B.n494 71.676
R1400 B.n631 B.n495 71.676
R1401 B.n627 B.n496 71.676
R1402 B.n623 B.n497 71.676
R1403 B.n618 B.n498 71.676
R1404 B.n614 B.n499 71.676
R1405 B.n610 B.n500 71.676
R1406 B.n606 B.n501 71.676
R1407 B.n602 B.n502 71.676
R1408 B.n598 B.n503 71.676
R1409 B.n594 B.n504 71.676
R1410 B.n590 B.n505 71.676
R1411 B.n586 B.n506 71.676
R1412 B.n582 B.n507 71.676
R1413 B.n578 B.n508 71.676
R1414 B.n574 B.n509 71.676
R1415 B.n570 B.n510 71.676
R1416 B.n566 B.n511 71.676
R1417 B.n562 B.n512 71.676
R1418 B.n558 B.n513 71.676
R1419 B.n554 B.n514 71.676
R1420 B.n550 B.n515 71.676
R1421 B.n546 B.n516 71.676
R1422 B.n542 B.n517 71.676
R1423 B.n538 B.n518 71.676
R1424 B.n534 B.n519 71.676
R1425 B.n530 B.n520 71.676
R1426 B.n730 B.n470 71.676
R1427 B.n724 B.n471 71.676
R1428 B.n720 B.n472 71.676
R1429 B.n716 B.n473 71.676
R1430 B.n712 B.n474 71.676
R1431 B.n708 B.n475 71.676
R1432 B.n704 B.n476 71.676
R1433 B.n700 B.n477 71.676
R1434 B.n696 B.n478 71.676
R1435 B.n692 B.n479 71.676
R1436 B.n688 B.n480 71.676
R1437 B.n684 B.n481 71.676
R1438 B.n680 B.n482 71.676
R1439 B.n676 B.n483 71.676
R1440 B.n672 B.n484 71.676
R1441 B.n668 B.n485 71.676
R1442 B.n664 B.n486 71.676
R1443 B.n660 B.n487 71.676
R1444 B.n656 B.n488 71.676
R1445 B.n652 B.n489 71.676
R1446 B.n648 B.n490 71.676
R1447 B.n644 B.n491 71.676
R1448 B.n640 B.n492 71.676
R1449 B.n636 B.n493 71.676
R1450 B.n632 B.n494 71.676
R1451 B.n628 B.n495 71.676
R1452 B.n624 B.n496 71.676
R1453 B.n619 B.n497 71.676
R1454 B.n615 B.n498 71.676
R1455 B.n611 B.n499 71.676
R1456 B.n607 B.n500 71.676
R1457 B.n603 B.n501 71.676
R1458 B.n599 B.n502 71.676
R1459 B.n595 B.n503 71.676
R1460 B.n591 B.n504 71.676
R1461 B.n587 B.n505 71.676
R1462 B.n583 B.n506 71.676
R1463 B.n579 B.n507 71.676
R1464 B.n575 B.n508 71.676
R1465 B.n571 B.n509 71.676
R1466 B.n567 B.n510 71.676
R1467 B.n563 B.n511 71.676
R1468 B.n559 B.n512 71.676
R1469 B.n555 B.n513 71.676
R1470 B.n551 B.n514 71.676
R1471 B.n547 B.n515 71.676
R1472 B.n543 B.n516 71.676
R1473 B.n539 B.n517 71.676
R1474 B.n535 B.n518 71.676
R1475 B.n531 B.n519 71.676
R1476 B.n527 B.n520 71.676
R1477 B.n1086 B.n1085 71.676
R1478 B.n1086 B.n2 71.676
R1479 B.n157 B.t23 71.0702
R1480 B.n526 B.t15 71.0702
R1481 B.n160 B.t20 71.0524
R1482 B.n523 B.t12 71.0524
R1483 B.n251 B.n160 59.5399
R1484 B.n158 B.n157 59.5399
R1485 B.n621 B.n526 59.5399
R1486 B.n524 B.n523 59.5399
R1487 B.n160 B.n159 52.3641
R1488 B.n157 B.n156 52.3641
R1489 B.n526 B.n525 52.3641
R1490 B.n523 B.n522 52.3641
R1491 B.n736 B.n467 39.2553
R1492 B.n736 B.n463 39.2553
R1493 B.n742 B.n463 39.2553
R1494 B.n742 B.n459 39.2553
R1495 B.n748 B.n459 39.2553
R1496 B.n748 B.n455 39.2553
R1497 B.n754 B.n455 39.2553
R1498 B.n760 B.n451 39.2553
R1499 B.n760 B.n447 39.2553
R1500 B.n766 B.n447 39.2553
R1501 B.n766 B.n443 39.2553
R1502 B.n772 B.n443 39.2553
R1503 B.n772 B.n439 39.2553
R1504 B.n778 B.n439 39.2553
R1505 B.n778 B.n434 39.2553
R1506 B.n784 B.n434 39.2553
R1507 B.n784 B.n435 39.2553
R1508 B.n790 B.n427 39.2553
R1509 B.n796 B.n427 39.2553
R1510 B.n796 B.n423 39.2553
R1511 B.n802 B.n423 39.2553
R1512 B.n802 B.n418 39.2553
R1513 B.n808 B.n418 39.2553
R1514 B.n808 B.n419 39.2553
R1515 B.n814 B.n411 39.2553
R1516 B.n820 B.n411 39.2553
R1517 B.n820 B.n407 39.2553
R1518 B.n826 B.n407 39.2553
R1519 B.n826 B.n402 39.2553
R1520 B.n832 B.n402 39.2553
R1521 B.n832 B.n403 39.2553
R1522 B.n838 B.n395 39.2553
R1523 B.n844 B.n395 39.2553
R1524 B.n844 B.n391 39.2553
R1525 B.n850 B.n391 39.2553
R1526 B.n850 B.n387 39.2553
R1527 B.n856 B.n387 39.2553
R1528 B.n862 B.n383 39.2553
R1529 B.n862 B.n379 39.2553
R1530 B.n868 B.n379 39.2553
R1531 B.n868 B.n375 39.2553
R1532 B.n874 B.n375 39.2553
R1533 B.n874 B.n371 39.2553
R1534 B.n880 B.n371 39.2553
R1535 B.n887 B.n367 39.2553
R1536 B.n887 B.n363 39.2553
R1537 B.n893 B.n363 39.2553
R1538 B.n893 B.n4 39.2553
R1539 B.n1084 B.n4 39.2553
R1540 B.n1084 B.n1083 39.2553
R1541 B.n1083 B.n1082 39.2553
R1542 B.n1082 B.n8 39.2553
R1543 B.n12 B.n8 39.2553
R1544 B.n1075 B.n12 39.2553
R1545 B.n1075 B.n1074 39.2553
R1546 B.n1073 B.n16 39.2553
R1547 B.n1067 B.n16 39.2553
R1548 B.n1067 B.n1066 39.2553
R1549 B.n1066 B.n1065 39.2553
R1550 B.n1065 B.n23 39.2553
R1551 B.n1059 B.n23 39.2553
R1552 B.n1059 B.n1058 39.2553
R1553 B.n1057 B.n30 39.2553
R1554 B.n1051 B.n30 39.2553
R1555 B.n1051 B.n1050 39.2553
R1556 B.n1050 B.n1049 39.2553
R1557 B.n1049 B.n37 39.2553
R1558 B.n1043 B.n37 39.2553
R1559 B.n1042 B.n1041 39.2553
R1560 B.n1041 B.n44 39.2553
R1561 B.n1035 B.n44 39.2553
R1562 B.n1035 B.n1034 39.2553
R1563 B.n1034 B.n1033 39.2553
R1564 B.n1033 B.n51 39.2553
R1565 B.n1027 B.n51 39.2553
R1566 B.n1026 B.n1025 39.2553
R1567 B.n1025 B.n58 39.2553
R1568 B.n1019 B.n58 39.2553
R1569 B.n1019 B.n1018 39.2553
R1570 B.n1018 B.n1017 39.2553
R1571 B.n1017 B.n65 39.2553
R1572 B.n1011 B.n65 39.2553
R1573 B.n1010 B.n1009 39.2553
R1574 B.n1009 B.n72 39.2553
R1575 B.n1003 B.n72 39.2553
R1576 B.n1003 B.n1002 39.2553
R1577 B.n1002 B.n1001 39.2553
R1578 B.n1001 B.n79 39.2553
R1579 B.n995 B.n79 39.2553
R1580 B.n995 B.n994 39.2553
R1581 B.n994 B.n993 39.2553
R1582 B.n993 B.n86 39.2553
R1583 B.n987 B.n986 39.2553
R1584 B.n986 B.n985 39.2553
R1585 B.n985 B.n93 39.2553
R1586 B.n979 B.n93 39.2553
R1587 B.n979 B.n978 39.2553
R1588 B.n978 B.n977 39.2553
R1589 B.n977 B.n100 39.2553
R1590 B.t11 B.n451 38.678
R1591 B.n856 B.t9 38.678
R1592 B.t1 B.n1057 38.678
R1593 B.t18 B.n86 38.678
R1594 B.n838 B.t5 37.5235
R1595 B.n1043 B.t3 37.5235
R1596 B.n733 B.n732 36.6834
R1597 B.n528 B.n465 36.6834
R1598 B.n968 B.n967 36.6834
R1599 B.n974 B.n973 36.6834
R1600 B.n880 B.t7 36.3689
R1601 B.t4 B.n1073 36.3689
R1602 B.n814 B.t2 35.2144
R1603 B.n1027 B.t6 35.2144
R1604 B.n790 B.t0 32.9053
R1605 B.n1011 B.t8 32.9053
R1606 B B.n1087 18.0485
R1607 B.n734 B.n733 10.6151
R1608 B.n734 B.n461 10.6151
R1609 B.n744 B.n461 10.6151
R1610 B.n745 B.n744 10.6151
R1611 B.n746 B.n745 10.6151
R1612 B.n746 B.n453 10.6151
R1613 B.n756 B.n453 10.6151
R1614 B.n757 B.n756 10.6151
R1615 B.n758 B.n757 10.6151
R1616 B.n758 B.n445 10.6151
R1617 B.n768 B.n445 10.6151
R1618 B.n769 B.n768 10.6151
R1619 B.n770 B.n769 10.6151
R1620 B.n770 B.n437 10.6151
R1621 B.n780 B.n437 10.6151
R1622 B.n781 B.n780 10.6151
R1623 B.n782 B.n781 10.6151
R1624 B.n782 B.n429 10.6151
R1625 B.n792 B.n429 10.6151
R1626 B.n793 B.n792 10.6151
R1627 B.n794 B.n793 10.6151
R1628 B.n794 B.n421 10.6151
R1629 B.n804 B.n421 10.6151
R1630 B.n805 B.n804 10.6151
R1631 B.n806 B.n805 10.6151
R1632 B.n806 B.n413 10.6151
R1633 B.n816 B.n413 10.6151
R1634 B.n817 B.n816 10.6151
R1635 B.n818 B.n817 10.6151
R1636 B.n818 B.n405 10.6151
R1637 B.n828 B.n405 10.6151
R1638 B.n829 B.n828 10.6151
R1639 B.n830 B.n829 10.6151
R1640 B.n830 B.n397 10.6151
R1641 B.n840 B.n397 10.6151
R1642 B.n841 B.n840 10.6151
R1643 B.n842 B.n841 10.6151
R1644 B.n842 B.n389 10.6151
R1645 B.n852 B.n389 10.6151
R1646 B.n853 B.n852 10.6151
R1647 B.n854 B.n853 10.6151
R1648 B.n854 B.n381 10.6151
R1649 B.n864 B.n381 10.6151
R1650 B.n865 B.n864 10.6151
R1651 B.n866 B.n865 10.6151
R1652 B.n866 B.n373 10.6151
R1653 B.n876 B.n373 10.6151
R1654 B.n877 B.n876 10.6151
R1655 B.n878 B.n877 10.6151
R1656 B.n878 B.n365 10.6151
R1657 B.n889 B.n365 10.6151
R1658 B.n890 B.n889 10.6151
R1659 B.n891 B.n890 10.6151
R1660 B.n891 B.n0 10.6151
R1661 B.n732 B.n469 10.6151
R1662 B.n727 B.n469 10.6151
R1663 B.n727 B.n726 10.6151
R1664 B.n726 B.n725 10.6151
R1665 B.n725 B.n722 10.6151
R1666 B.n722 B.n721 10.6151
R1667 B.n721 B.n718 10.6151
R1668 B.n718 B.n717 10.6151
R1669 B.n717 B.n714 10.6151
R1670 B.n714 B.n713 10.6151
R1671 B.n713 B.n710 10.6151
R1672 B.n710 B.n709 10.6151
R1673 B.n709 B.n706 10.6151
R1674 B.n706 B.n705 10.6151
R1675 B.n705 B.n702 10.6151
R1676 B.n702 B.n701 10.6151
R1677 B.n701 B.n698 10.6151
R1678 B.n698 B.n697 10.6151
R1679 B.n697 B.n694 10.6151
R1680 B.n694 B.n693 10.6151
R1681 B.n693 B.n690 10.6151
R1682 B.n690 B.n689 10.6151
R1683 B.n689 B.n686 10.6151
R1684 B.n686 B.n685 10.6151
R1685 B.n685 B.n682 10.6151
R1686 B.n682 B.n681 10.6151
R1687 B.n681 B.n678 10.6151
R1688 B.n678 B.n677 10.6151
R1689 B.n677 B.n674 10.6151
R1690 B.n674 B.n673 10.6151
R1691 B.n673 B.n670 10.6151
R1692 B.n670 B.n669 10.6151
R1693 B.n669 B.n666 10.6151
R1694 B.n666 B.n665 10.6151
R1695 B.n665 B.n662 10.6151
R1696 B.n662 B.n661 10.6151
R1697 B.n661 B.n658 10.6151
R1698 B.n658 B.n657 10.6151
R1699 B.n657 B.n654 10.6151
R1700 B.n654 B.n653 10.6151
R1701 B.n653 B.n650 10.6151
R1702 B.n650 B.n649 10.6151
R1703 B.n649 B.n646 10.6151
R1704 B.n646 B.n645 10.6151
R1705 B.n645 B.n642 10.6151
R1706 B.n642 B.n641 10.6151
R1707 B.n638 B.n637 10.6151
R1708 B.n637 B.n634 10.6151
R1709 B.n634 B.n633 10.6151
R1710 B.n633 B.n630 10.6151
R1711 B.n630 B.n629 10.6151
R1712 B.n629 B.n626 10.6151
R1713 B.n626 B.n625 10.6151
R1714 B.n625 B.n622 10.6151
R1715 B.n620 B.n617 10.6151
R1716 B.n617 B.n616 10.6151
R1717 B.n616 B.n613 10.6151
R1718 B.n613 B.n612 10.6151
R1719 B.n612 B.n609 10.6151
R1720 B.n609 B.n608 10.6151
R1721 B.n608 B.n605 10.6151
R1722 B.n605 B.n604 10.6151
R1723 B.n604 B.n601 10.6151
R1724 B.n601 B.n600 10.6151
R1725 B.n600 B.n597 10.6151
R1726 B.n597 B.n596 10.6151
R1727 B.n596 B.n593 10.6151
R1728 B.n593 B.n592 10.6151
R1729 B.n592 B.n589 10.6151
R1730 B.n589 B.n588 10.6151
R1731 B.n588 B.n585 10.6151
R1732 B.n585 B.n584 10.6151
R1733 B.n584 B.n581 10.6151
R1734 B.n581 B.n580 10.6151
R1735 B.n580 B.n577 10.6151
R1736 B.n577 B.n576 10.6151
R1737 B.n576 B.n573 10.6151
R1738 B.n573 B.n572 10.6151
R1739 B.n572 B.n569 10.6151
R1740 B.n569 B.n568 10.6151
R1741 B.n568 B.n565 10.6151
R1742 B.n565 B.n564 10.6151
R1743 B.n564 B.n561 10.6151
R1744 B.n561 B.n560 10.6151
R1745 B.n560 B.n557 10.6151
R1746 B.n557 B.n556 10.6151
R1747 B.n556 B.n553 10.6151
R1748 B.n553 B.n552 10.6151
R1749 B.n552 B.n549 10.6151
R1750 B.n549 B.n548 10.6151
R1751 B.n548 B.n545 10.6151
R1752 B.n545 B.n544 10.6151
R1753 B.n544 B.n541 10.6151
R1754 B.n541 B.n540 10.6151
R1755 B.n540 B.n537 10.6151
R1756 B.n537 B.n536 10.6151
R1757 B.n536 B.n533 10.6151
R1758 B.n533 B.n532 10.6151
R1759 B.n532 B.n529 10.6151
R1760 B.n529 B.n528 10.6151
R1761 B.n738 B.n465 10.6151
R1762 B.n739 B.n738 10.6151
R1763 B.n740 B.n739 10.6151
R1764 B.n740 B.n457 10.6151
R1765 B.n750 B.n457 10.6151
R1766 B.n751 B.n750 10.6151
R1767 B.n752 B.n751 10.6151
R1768 B.n752 B.n449 10.6151
R1769 B.n762 B.n449 10.6151
R1770 B.n763 B.n762 10.6151
R1771 B.n764 B.n763 10.6151
R1772 B.n764 B.n441 10.6151
R1773 B.n774 B.n441 10.6151
R1774 B.n775 B.n774 10.6151
R1775 B.n776 B.n775 10.6151
R1776 B.n776 B.n432 10.6151
R1777 B.n786 B.n432 10.6151
R1778 B.n787 B.n786 10.6151
R1779 B.n788 B.n787 10.6151
R1780 B.n788 B.n425 10.6151
R1781 B.n798 B.n425 10.6151
R1782 B.n799 B.n798 10.6151
R1783 B.n800 B.n799 10.6151
R1784 B.n800 B.n416 10.6151
R1785 B.n810 B.n416 10.6151
R1786 B.n811 B.n810 10.6151
R1787 B.n812 B.n811 10.6151
R1788 B.n812 B.n409 10.6151
R1789 B.n822 B.n409 10.6151
R1790 B.n823 B.n822 10.6151
R1791 B.n824 B.n823 10.6151
R1792 B.n824 B.n400 10.6151
R1793 B.n834 B.n400 10.6151
R1794 B.n835 B.n834 10.6151
R1795 B.n836 B.n835 10.6151
R1796 B.n836 B.n393 10.6151
R1797 B.n846 B.n393 10.6151
R1798 B.n847 B.n846 10.6151
R1799 B.n848 B.n847 10.6151
R1800 B.n848 B.n385 10.6151
R1801 B.n858 B.n385 10.6151
R1802 B.n859 B.n858 10.6151
R1803 B.n860 B.n859 10.6151
R1804 B.n860 B.n377 10.6151
R1805 B.n870 B.n377 10.6151
R1806 B.n871 B.n870 10.6151
R1807 B.n872 B.n871 10.6151
R1808 B.n872 B.n369 10.6151
R1809 B.n882 B.n369 10.6151
R1810 B.n883 B.n882 10.6151
R1811 B.n885 B.n883 10.6151
R1812 B.n885 B.n884 10.6151
R1813 B.n884 B.n361 10.6151
R1814 B.n896 B.n361 10.6151
R1815 B.n897 B.n896 10.6151
R1816 B.n898 B.n897 10.6151
R1817 B.n899 B.n898 10.6151
R1818 B.n900 B.n899 10.6151
R1819 B.n903 B.n900 10.6151
R1820 B.n904 B.n903 10.6151
R1821 B.n905 B.n904 10.6151
R1822 B.n906 B.n905 10.6151
R1823 B.n908 B.n906 10.6151
R1824 B.n909 B.n908 10.6151
R1825 B.n910 B.n909 10.6151
R1826 B.n911 B.n910 10.6151
R1827 B.n913 B.n911 10.6151
R1828 B.n914 B.n913 10.6151
R1829 B.n915 B.n914 10.6151
R1830 B.n916 B.n915 10.6151
R1831 B.n918 B.n916 10.6151
R1832 B.n919 B.n918 10.6151
R1833 B.n920 B.n919 10.6151
R1834 B.n921 B.n920 10.6151
R1835 B.n923 B.n921 10.6151
R1836 B.n924 B.n923 10.6151
R1837 B.n925 B.n924 10.6151
R1838 B.n926 B.n925 10.6151
R1839 B.n928 B.n926 10.6151
R1840 B.n929 B.n928 10.6151
R1841 B.n930 B.n929 10.6151
R1842 B.n931 B.n930 10.6151
R1843 B.n933 B.n931 10.6151
R1844 B.n934 B.n933 10.6151
R1845 B.n935 B.n934 10.6151
R1846 B.n936 B.n935 10.6151
R1847 B.n938 B.n936 10.6151
R1848 B.n939 B.n938 10.6151
R1849 B.n940 B.n939 10.6151
R1850 B.n941 B.n940 10.6151
R1851 B.n943 B.n941 10.6151
R1852 B.n944 B.n943 10.6151
R1853 B.n945 B.n944 10.6151
R1854 B.n946 B.n945 10.6151
R1855 B.n948 B.n946 10.6151
R1856 B.n949 B.n948 10.6151
R1857 B.n950 B.n949 10.6151
R1858 B.n951 B.n950 10.6151
R1859 B.n953 B.n951 10.6151
R1860 B.n954 B.n953 10.6151
R1861 B.n955 B.n954 10.6151
R1862 B.n956 B.n955 10.6151
R1863 B.n958 B.n956 10.6151
R1864 B.n959 B.n958 10.6151
R1865 B.n960 B.n959 10.6151
R1866 B.n961 B.n960 10.6151
R1867 B.n963 B.n961 10.6151
R1868 B.n964 B.n963 10.6151
R1869 B.n965 B.n964 10.6151
R1870 B.n966 B.n965 10.6151
R1871 B.n967 B.n966 10.6151
R1872 B.n1079 B.n1 10.6151
R1873 B.n1079 B.n1078 10.6151
R1874 B.n1078 B.n1077 10.6151
R1875 B.n1077 B.n10 10.6151
R1876 B.n1071 B.n10 10.6151
R1877 B.n1071 B.n1070 10.6151
R1878 B.n1070 B.n1069 10.6151
R1879 B.n1069 B.n18 10.6151
R1880 B.n1063 B.n18 10.6151
R1881 B.n1063 B.n1062 10.6151
R1882 B.n1062 B.n1061 10.6151
R1883 B.n1061 B.n25 10.6151
R1884 B.n1055 B.n25 10.6151
R1885 B.n1055 B.n1054 10.6151
R1886 B.n1054 B.n1053 10.6151
R1887 B.n1053 B.n32 10.6151
R1888 B.n1047 B.n32 10.6151
R1889 B.n1047 B.n1046 10.6151
R1890 B.n1046 B.n1045 10.6151
R1891 B.n1045 B.n39 10.6151
R1892 B.n1039 B.n39 10.6151
R1893 B.n1039 B.n1038 10.6151
R1894 B.n1038 B.n1037 10.6151
R1895 B.n1037 B.n46 10.6151
R1896 B.n1031 B.n46 10.6151
R1897 B.n1031 B.n1030 10.6151
R1898 B.n1030 B.n1029 10.6151
R1899 B.n1029 B.n53 10.6151
R1900 B.n1023 B.n53 10.6151
R1901 B.n1023 B.n1022 10.6151
R1902 B.n1022 B.n1021 10.6151
R1903 B.n1021 B.n60 10.6151
R1904 B.n1015 B.n60 10.6151
R1905 B.n1015 B.n1014 10.6151
R1906 B.n1014 B.n1013 10.6151
R1907 B.n1013 B.n67 10.6151
R1908 B.n1007 B.n67 10.6151
R1909 B.n1007 B.n1006 10.6151
R1910 B.n1006 B.n1005 10.6151
R1911 B.n1005 B.n74 10.6151
R1912 B.n999 B.n74 10.6151
R1913 B.n999 B.n998 10.6151
R1914 B.n998 B.n997 10.6151
R1915 B.n997 B.n81 10.6151
R1916 B.n991 B.n81 10.6151
R1917 B.n991 B.n990 10.6151
R1918 B.n990 B.n989 10.6151
R1919 B.n989 B.n88 10.6151
R1920 B.n983 B.n88 10.6151
R1921 B.n983 B.n982 10.6151
R1922 B.n982 B.n981 10.6151
R1923 B.n981 B.n95 10.6151
R1924 B.n975 B.n95 10.6151
R1925 B.n975 B.n974 10.6151
R1926 B.n973 B.n102 10.6151
R1927 B.n162 B.n102 10.6151
R1928 B.n163 B.n162 10.6151
R1929 B.n166 B.n163 10.6151
R1930 B.n167 B.n166 10.6151
R1931 B.n170 B.n167 10.6151
R1932 B.n171 B.n170 10.6151
R1933 B.n174 B.n171 10.6151
R1934 B.n175 B.n174 10.6151
R1935 B.n178 B.n175 10.6151
R1936 B.n179 B.n178 10.6151
R1937 B.n182 B.n179 10.6151
R1938 B.n183 B.n182 10.6151
R1939 B.n186 B.n183 10.6151
R1940 B.n187 B.n186 10.6151
R1941 B.n190 B.n187 10.6151
R1942 B.n191 B.n190 10.6151
R1943 B.n194 B.n191 10.6151
R1944 B.n195 B.n194 10.6151
R1945 B.n198 B.n195 10.6151
R1946 B.n199 B.n198 10.6151
R1947 B.n202 B.n199 10.6151
R1948 B.n203 B.n202 10.6151
R1949 B.n206 B.n203 10.6151
R1950 B.n207 B.n206 10.6151
R1951 B.n210 B.n207 10.6151
R1952 B.n211 B.n210 10.6151
R1953 B.n214 B.n211 10.6151
R1954 B.n215 B.n214 10.6151
R1955 B.n218 B.n215 10.6151
R1956 B.n219 B.n218 10.6151
R1957 B.n222 B.n219 10.6151
R1958 B.n223 B.n222 10.6151
R1959 B.n226 B.n223 10.6151
R1960 B.n227 B.n226 10.6151
R1961 B.n230 B.n227 10.6151
R1962 B.n231 B.n230 10.6151
R1963 B.n234 B.n231 10.6151
R1964 B.n235 B.n234 10.6151
R1965 B.n238 B.n235 10.6151
R1966 B.n239 B.n238 10.6151
R1967 B.n242 B.n239 10.6151
R1968 B.n243 B.n242 10.6151
R1969 B.n246 B.n243 10.6151
R1970 B.n247 B.n246 10.6151
R1971 B.n250 B.n247 10.6151
R1972 B.n255 B.n252 10.6151
R1973 B.n256 B.n255 10.6151
R1974 B.n259 B.n256 10.6151
R1975 B.n260 B.n259 10.6151
R1976 B.n263 B.n260 10.6151
R1977 B.n264 B.n263 10.6151
R1978 B.n267 B.n264 10.6151
R1979 B.n268 B.n267 10.6151
R1980 B.n272 B.n271 10.6151
R1981 B.n275 B.n272 10.6151
R1982 B.n276 B.n275 10.6151
R1983 B.n279 B.n276 10.6151
R1984 B.n280 B.n279 10.6151
R1985 B.n283 B.n280 10.6151
R1986 B.n284 B.n283 10.6151
R1987 B.n287 B.n284 10.6151
R1988 B.n288 B.n287 10.6151
R1989 B.n291 B.n288 10.6151
R1990 B.n292 B.n291 10.6151
R1991 B.n295 B.n292 10.6151
R1992 B.n296 B.n295 10.6151
R1993 B.n299 B.n296 10.6151
R1994 B.n300 B.n299 10.6151
R1995 B.n303 B.n300 10.6151
R1996 B.n304 B.n303 10.6151
R1997 B.n307 B.n304 10.6151
R1998 B.n308 B.n307 10.6151
R1999 B.n311 B.n308 10.6151
R2000 B.n312 B.n311 10.6151
R2001 B.n315 B.n312 10.6151
R2002 B.n316 B.n315 10.6151
R2003 B.n319 B.n316 10.6151
R2004 B.n320 B.n319 10.6151
R2005 B.n323 B.n320 10.6151
R2006 B.n324 B.n323 10.6151
R2007 B.n327 B.n324 10.6151
R2008 B.n328 B.n327 10.6151
R2009 B.n331 B.n328 10.6151
R2010 B.n332 B.n331 10.6151
R2011 B.n335 B.n332 10.6151
R2012 B.n336 B.n335 10.6151
R2013 B.n339 B.n336 10.6151
R2014 B.n340 B.n339 10.6151
R2015 B.n343 B.n340 10.6151
R2016 B.n344 B.n343 10.6151
R2017 B.n347 B.n344 10.6151
R2018 B.n348 B.n347 10.6151
R2019 B.n351 B.n348 10.6151
R2020 B.n352 B.n351 10.6151
R2021 B.n355 B.n352 10.6151
R2022 B.n356 B.n355 10.6151
R2023 B.n359 B.n356 10.6151
R2024 B.n360 B.n359 10.6151
R2025 B.n968 B.n360 10.6151
R2026 B.n1087 B.n0 8.11757
R2027 B.n1087 B.n1 8.11757
R2028 B.n638 B.n524 6.5566
R2029 B.n622 B.n621 6.5566
R2030 B.n252 B.n251 6.5566
R2031 B.n268 B.n158 6.5566
R2032 B.n435 B.t0 6.35054
R2033 B.t8 B.n1010 6.35054
R2034 B.n641 B.n524 4.05904
R2035 B.n621 B.n620 4.05904
R2036 B.n251 B.n250 4.05904
R2037 B.n271 B.n158 4.05904
R2038 B.n419 B.t2 4.04143
R2039 B.t6 B.n1026 4.04143
R2040 B.t7 B.n367 2.88688
R2041 B.n1074 B.t4 2.88688
R2042 B.n403 B.t5 1.73233
R2043 B.t3 B.n1042 1.73233
R2044 B.n754 B.t11 0.577776
R2045 B.t9 B.n383 0.577776
R2046 B.n1058 B.t1 0.577776
R2047 B.n987 B.t18 0.577776
R2048 VP.n21 VP.t5 173.024
R2049 VP.n23 VP.n20 161.3
R2050 VP.n25 VP.n24 161.3
R2051 VP.n26 VP.n19 161.3
R2052 VP.n28 VP.n27 161.3
R2053 VP.n29 VP.n18 161.3
R2054 VP.n32 VP.n31 161.3
R2055 VP.n33 VP.n17 161.3
R2056 VP.n35 VP.n34 161.3
R2057 VP.n36 VP.n16 161.3
R2058 VP.n38 VP.n37 161.3
R2059 VP.n40 VP.n39 161.3
R2060 VP.n41 VP.n14 161.3
R2061 VP.n43 VP.n42 161.3
R2062 VP.n44 VP.n13 161.3
R2063 VP.n46 VP.n45 161.3
R2064 VP.n47 VP.n12 161.3
R2065 VP.n86 VP.n0 161.3
R2066 VP.n85 VP.n84 161.3
R2067 VP.n83 VP.n1 161.3
R2068 VP.n82 VP.n81 161.3
R2069 VP.n80 VP.n2 161.3
R2070 VP.n79 VP.n78 161.3
R2071 VP.n77 VP.n76 161.3
R2072 VP.n75 VP.n4 161.3
R2073 VP.n74 VP.n73 161.3
R2074 VP.n72 VP.n5 161.3
R2075 VP.n71 VP.n70 161.3
R2076 VP.n68 VP.n6 161.3
R2077 VP.n67 VP.n66 161.3
R2078 VP.n65 VP.n7 161.3
R2079 VP.n64 VP.n63 161.3
R2080 VP.n62 VP.n8 161.3
R2081 VP.n60 VP.n59 161.3
R2082 VP.n58 VP.n9 161.3
R2083 VP.n57 VP.n56 161.3
R2084 VP.n55 VP.n10 161.3
R2085 VP.n54 VP.n53 161.3
R2086 VP.n52 VP.n11 161.3
R2087 VP.n50 VP.t1 140.126
R2088 VP.n61 VP.t4 140.126
R2089 VP.n69 VP.t7 140.126
R2090 VP.n3 VP.t0 140.126
R2091 VP.n87 VP.t6 140.126
R2092 VP.n48 VP.t2 140.126
R2093 VP.n15 VP.t8 140.126
R2094 VP.n30 VP.t3 140.126
R2095 VP.n22 VP.t9 140.126
R2096 VP.n51 VP.n50 103.531
R2097 VP.n88 VP.n87 103.531
R2098 VP.n49 VP.n48 103.531
R2099 VP.n56 VP.n55 56.5617
R2100 VP.n81 VP.n1 56.5617
R2101 VP.n42 VP.n13 56.5617
R2102 VP.n51 VP.n49 53.136
R2103 VP.n22 VP.n21 50.3824
R2104 VP.n63 VP.n7 50.2647
R2105 VP.n75 VP.n74 50.2647
R2106 VP.n36 VP.n35 50.2647
R2107 VP.n24 VP.n19 50.2647
R2108 VP.n67 VP.n7 30.8893
R2109 VP.n74 VP.n5 30.8893
R2110 VP.n35 VP.n17 30.8893
R2111 VP.n28 VP.n19 30.8893
R2112 VP.n54 VP.n11 24.5923
R2113 VP.n55 VP.n54 24.5923
R2114 VP.n56 VP.n9 24.5923
R2115 VP.n60 VP.n9 24.5923
R2116 VP.n63 VP.n62 24.5923
R2117 VP.n68 VP.n67 24.5923
R2118 VP.n70 VP.n5 24.5923
R2119 VP.n76 VP.n75 24.5923
R2120 VP.n80 VP.n79 24.5923
R2121 VP.n81 VP.n80 24.5923
R2122 VP.n85 VP.n1 24.5923
R2123 VP.n86 VP.n85 24.5923
R2124 VP.n46 VP.n13 24.5923
R2125 VP.n47 VP.n46 24.5923
R2126 VP.n37 VP.n36 24.5923
R2127 VP.n41 VP.n40 24.5923
R2128 VP.n42 VP.n41 24.5923
R2129 VP.n29 VP.n28 24.5923
R2130 VP.n31 VP.n17 24.5923
R2131 VP.n24 VP.n23 24.5923
R2132 VP.n62 VP.n61 22.1332
R2133 VP.n76 VP.n3 22.1332
R2134 VP.n37 VP.n15 22.1332
R2135 VP.n23 VP.n22 22.1332
R2136 VP.n69 VP.n68 12.2964
R2137 VP.n70 VP.n69 12.2964
R2138 VP.n30 VP.n29 12.2964
R2139 VP.n31 VP.n30 12.2964
R2140 VP.n50 VP.n11 7.37805
R2141 VP.n87 VP.n86 7.37805
R2142 VP.n48 VP.n47 7.37805
R2143 VP.n21 VP.n20 6.9978
R2144 VP.n61 VP.n60 2.45968
R2145 VP.n79 VP.n3 2.45968
R2146 VP.n40 VP.n15 2.45968
R2147 VP.n49 VP.n12 0.278335
R2148 VP.n52 VP.n51 0.278335
R2149 VP.n88 VP.n0 0.278335
R2150 VP.n25 VP.n20 0.189894
R2151 VP.n26 VP.n25 0.189894
R2152 VP.n27 VP.n26 0.189894
R2153 VP.n27 VP.n18 0.189894
R2154 VP.n32 VP.n18 0.189894
R2155 VP.n33 VP.n32 0.189894
R2156 VP.n34 VP.n33 0.189894
R2157 VP.n34 VP.n16 0.189894
R2158 VP.n38 VP.n16 0.189894
R2159 VP.n39 VP.n38 0.189894
R2160 VP.n39 VP.n14 0.189894
R2161 VP.n43 VP.n14 0.189894
R2162 VP.n44 VP.n43 0.189894
R2163 VP.n45 VP.n44 0.189894
R2164 VP.n45 VP.n12 0.189894
R2165 VP.n53 VP.n52 0.189894
R2166 VP.n53 VP.n10 0.189894
R2167 VP.n57 VP.n10 0.189894
R2168 VP.n58 VP.n57 0.189894
R2169 VP.n59 VP.n58 0.189894
R2170 VP.n59 VP.n8 0.189894
R2171 VP.n64 VP.n8 0.189894
R2172 VP.n65 VP.n64 0.189894
R2173 VP.n66 VP.n65 0.189894
R2174 VP.n66 VP.n6 0.189894
R2175 VP.n71 VP.n6 0.189894
R2176 VP.n72 VP.n71 0.189894
R2177 VP.n73 VP.n72 0.189894
R2178 VP.n73 VP.n4 0.189894
R2179 VP.n77 VP.n4 0.189894
R2180 VP.n78 VP.n77 0.189894
R2181 VP.n78 VP.n2 0.189894
R2182 VP.n82 VP.n2 0.189894
R2183 VP.n83 VP.n82 0.189894
R2184 VP.n84 VP.n83 0.189894
R2185 VP.n84 VP.n0 0.189894
R2186 VP VP.n88 0.153485
R2187 VDD1.n1 VDD1.t4 69.0982
R2188 VDD1.n3 VDD1.t8 69.098
R2189 VDD1.n5 VDD1.n4 67.0239
R2190 VDD1.n1 VDD1.n0 65.3338
R2191 VDD1.n7 VDD1.n6 65.3336
R2192 VDD1.n3 VDD1.n2 65.3336
R2193 VDD1.n7 VDD1.n5 48.3974
R2194 VDD1 VDD1.n7 1.688
R2195 VDD1.n6 VDD1.t1 1.43736
R2196 VDD1.n6 VDD1.t7 1.43736
R2197 VDD1.n0 VDD1.t0 1.43736
R2198 VDD1.n0 VDD1.t6 1.43736
R2199 VDD1.n4 VDD1.t9 1.43736
R2200 VDD1.n4 VDD1.t3 1.43736
R2201 VDD1.n2 VDD1.t5 1.43736
R2202 VDD1.n2 VDD1.t2 1.43736
R2203 VDD1 VDD1.n1 0.640586
R2204 VDD1.n5 VDD1.n3 0.527051
C0 VDD2 VP 0.554763f
C1 VDD2 VTAIL 11.2776f
C2 VN VDD2 11.939401f
C3 VTAIL VP 12.4211f
C4 VN VP 8.386781f
C5 VDD2 VDD1 2.02519f
C6 VN VTAIL 12.4067f
C7 VDD1 VP 12.3367f
C8 VDD1 VTAIL 11.228901f
C9 VN VDD1 0.153198f
C10 VDD2 B 7.260975f
C11 VDD1 B 7.230502f
C12 VTAIL B 8.732973f
C13 VN B 17.200882f
C14 VP B 15.67932f
C15 VDD1.t4 B 3.03438f
C16 VDD1.t0 B 0.262248f
C17 VDD1.t6 B 0.262248f
C18 VDD1.n0 B 2.36488f
C19 VDD1.n1 B 0.849796f
C20 VDD1.t8 B 3.03437f
C21 VDD1.t5 B 0.262248f
C22 VDD1.t2 B 0.262248f
C23 VDD1.n2 B 2.36488f
C24 VDD1.n3 B 0.842049f
C25 VDD1.t9 B 0.262248f
C26 VDD1.t3 B 0.262248f
C27 VDD1.n4 B 2.37783f
C28 VDD1.n5 B 2.89916f
C29 VDD1.t1 B 0.262248f
C30 VDD1.t7 B 0.262248f
C31 VDD1.n6 B 2.36488f
C32 VDD1.n7 B 3.08916f
C33 VP.n0 B 0.029916f
C34 VP.t6 B 2.02664f
C35 VP.n1 B 0.029847f
C36 VP.n2 B 0.022692f
C37 VP.t0 B 2.02664f
C38 VP.n3 B 0.713069f
C39 VP.n4 B 0.022692f
C40 VP.n5 B 0.045214f
C41 VP.n6 B 0.022692f
C42 VP.t7 B 2.02664f
C43 VP.n7 B 0.021395f
C44 VP.n8 B 0.022692f
C45 VP.t4 B 2.02664f
C46 VP.n9 B 0.04208f
C47 VP.n10 B 0.022692f
C48 VP.n11 B 0.027539f
C49 VP.n12 B 0.029916f
C50 VP.t2 B 2.02664f
C51 VP.n13 B 0.029847f
C52 VP.n14 B 0.022692f
C53 VP.t8 B 2.02664f
C54 VP.n15 B 0.713069f
C55 VP.n16 B 0.022692f
C56 VP.n17 B 0.045214f
C57 VP.n18 B 0.022692f
C58 VP.t3 B 2.02664f
C59 VP.n19 B 0.021395f
C60 VP.n20 B 0.213781f
C61 VP.t9 B 2.02664f
C62 VP.t5 B 2.18692f
C63 VP.n21 B 0.760682f
C64 VP.n22 B 0.784057f
C65 VP.n23 B 0.040003f
C66 VP.n24 B 0.041444f
C67 VP.n25 B 0.022692f
C68 VP.n26 B 0.022692f
C69 VP.n27 B 0.022692f
C70 VP.n28 B 0.045214f
C71 VP.n29 B 0.031693f
C72 VP.n30 B 0.713069f
C73 VP.n31 B 0.031693f
C74 VP.n32 B 0.022692f
C75 VP.n33 B 0.022692f
C76 VP.n34 B 0.022692f
C77 VP.n35 B 0.021395f
C78 VP.n36 B 0.041444f
C79 VP.n37 B 0.040003f
C80 VP.n38 B 0.022692f
C81 VP.n39 B 0.022692f
C82 VP.n40 B 0.023384f
C83 VP.n41 B 0.04208f
C84 VP.n42 B 0.036126f
C85 VP.n43 B 0.022692f
C86 VP.n44 B 0.022692f
C87 VP.n45 B 0.022692f
C88 VP.n46 B 0.04208f
C89 VP.n47 B 0.027539f
C90 VP.n48 B 0.778508f
C91 VP.n49 B 1.37748f
C92 VP.t1 B 2.02664f
C93 VP.n50 B 0.778508f
C94 VP.n51 B 1.39288f
C95 VP.n52 B 0.029916f
C96 VP.n53 B 0.022692f
C97 VP.n54 B 0.04208f
C98 VP.n55 B 0.029847f
C99 VP.n56 B 0.036126f
C100 VP.n57 B 0.022692f
C101 VP.n58 B 0.022692f
C102 VP.n59 B 0.022692f
C103 VP.n60 B 0.023384f
C104 VP.n61 B 0.713069f
C105 VP.n62 B 0.040003f
C106 VP.n63 B 0.041444f
C107 VP.n64 B 0.022692f
C108 VP.n65 B 0.022692f
C109 VP.n66 B 0.022692f
C110 VP.n67 B 0.045214f
C111 VP.n68 B 0.031693f
C112 VP.n69 B 0.713069f
C113 VP.n70 B 0.031693f
C114 VP.n71 B 0.022692f
C115 VP.n72 B 0.022692f
C116 VP.n73 B 0.022692f
C117 VP.n74 B 0.021395f
C118 VP.n75 B 0.041444f
C119 VP.n76 B 0.040003f
C120 VP.n77 B 0.022692f
C121 VP.n78 B 0.022692f
C122 VP.n79 B 0.023384f
C123 VP.n80 B 0.04208f
C124 VP.n81 B 0.036126f
C125 VP.n82 B 0.022692f
C126 VP.n83 B 0.022692f
C127 VP.n84 B 0.022692f
C128 VP.n85 B 0.04208f
C129 VP.n86 B 0.027539f
C130 VP.n87 B 0.778508f
C131 VP.n88 B 0.036571f
C132 VDD2.t0 B 3.00917f
C133 VDD2.t5 B 0.26007f
C134 VDD2.t9 B 0.26007f
C135 VDD2.n0 B 2.34524f
C136 VDD2.n1 B 0.835055f
C137 VDD2.t3 B 0.26007f
C138 VDD2.t6 B 0.26007f
C139 VDD2.n2 B 2.35808f
C140 VDD2.n3 B 2.7604f
C141 VDD2.t2 B 2.99439f
C142 VDD2.n4 B 3.02025f
C143 VDD2.t7 B 0.26007f
C144 VDD2.t1 B 0.26007f
C145 VDD2.n5 B 2.34524f
C146 VDD2.n6 B 0.418515f
C147 VDD2.t8 B 0.26007f
C148 VDD2.t4 B 0.26007f
C149 VDD2.n7 B 2.35805f
C150 VTAIL.t6 B 0.264936f
C151 VTAIL.t4 B 0.264936f
C152 VTAIL.n0 B 2.32431f
C153 VTAIL.n1 B 0.494922f
C154 VTAIL.t16 B 2.96707f
C155 VTAIL.n2 B 0.615778f
C156 VTAIL.t17 B 0.264936f
C157 VTAIL.t14 B 0.264936f
C158 VTAIL.n3 B 2.32431f
C159 VTAIL.n4 B 0.590383f
C160 VTAIL.t0 B 0.264936f
C161 VTAIL.t2 B 0.264936f
C162 VTAIL.n5 B 2.32431f
C163 VTAIL.n6 B 2.03464f
C164 VTAIL.t10 B 0.264936f
C165 VTAIL.t11 B 0.264936f
C166 VTAIL.n7 B 2.32432f
C167 VTAIL.n8 B 2.03464f
C168 VTAIL.t5 B 0.264936f
C169 VTAIL.t8 B 0.264936f
C170 VTAIL.n9 B 2.32432f
C171 VTAIL.n10 B 0.59038f
C172 VTAIL.t7 B 2.96707f
C173 VTAIL.n11 B 0.615776f
C174 VTAIL.t15 B 0.264936f
C175 VTAIL.t1 B 0.264936f
C176 VTAIL.n12 B 2.32432f
C177 VTAIL.n13 B 0.535976f
C178 VTAIL.t3 B 0.264936f
C179 VTAIL.t18 B 0.264936f
C180 VTAIL.n14 B 2.32432f
C181 VTAIL.n15 B 0.59038f
C182 VTAIL.t19 B 2.96707f
C183 VTAIL.n16 B 1.93197f
C184 VTAIL.t9 B 2.96707f
C185 VTAIL.n17 B 1.93197f
C186 VTAIL.t12 B 0.264936f
C187 VTAIL.t13 B 0.264936f
C188 VTAIL.n18 B 2.32431f
C189 VTAIL.n19 B 0.448966f
C190 VN.n0 B 0.029525f
C191 VN.t3 B 2.00023f
C192 VN.n1 B 0.029458f
C193 VN.n2 B 0.022396f
C194 VN.t6 B 2.00023f
C195 VN.n3 B 0.703773f
C196 VN.n4 B 0.022396f
C197 VN.n5 B 0.044625f
C198 VN.n6 B 0.022396f
C199 VN.t0 B 2.00023f
C200 VN.n7 B 0.021116f
C201 VN.n8 B 0.210994f
C202 VN.t4 B 2.00023f
C203 VN.t9 B 2.15841f
C204 VN.n9 B 0.750766f
C205 VN.n10 B 0.773836f
C206 VN.n11 B 0.039481f
C207 VN.n12 B 0.040903f
C208 VN.n13 B 0.022396f
C209 VN.n14 B 0.022396f
C210 VN.n15 B 0.022396f
C211 VN.n16 B 0.044625f
C212 VN.n17 B 0.03128f
C213 VN.n18 B 0.703773f
C214 VN.n19 B 0.03128f
C215 VN.n20 B 0.022396f
C216 VN.n21 B 0.022396f
C217 VN.n22 B 0.022396f
C218 VN.n23 B 0.021116f
C219 VN.n24 B 0.040903f
C220 VN.n25 B 0.039481f
C221 VN.n26 B 0.022396f
C222 VN.n27 B 0.022396f
C223 VN.n28 B 0.023079f
C224 VN.n29 B 0.041532f
C225 VN.n30 B 0.035655f
C226 VN.n31 B 0.022396f
C227 VN.n32 B 0.022396f
C228 VN.n33 B 0.022396f
C229 VN.n34 B 0.041532f
C230 VN.n35 B 0.02718f
C231 VN.n36 B 0.76836f
C232 VN.n37 B 0.036094f
C233 VN.n38 B 0.029525f
C234 VN.t7 B 2.00023f
C235 VN.n39 B 0.029458f
C236 VN.n40 B 0.022396f
C237 VN.t2 B 2.00023f
C238 VN.n41 B 0.703773f
C239 VN.n42 B 0.022396f
C240 VN.n43 B 0.044625f
C241 VN.n44 B 0.022396f
C242 VN.t8 B 2.00023f
C243 VN.n45 B 0.021116f
C244 VN.n46 B 0.210994f
C245 VN.t1 B 2.00023f
C246 VN.t5 B 2.15841f
C247 VN.n47 B 0.750766f
C248 VN.n48 B 0.773836f
C249 VN.n49 B 0.039481f
C250 VN.n50 B 0.040903f
C251 VN.n51 B 0.022396f
C252 VN.n52 B 0.022396f
C253 VN.n53 B 0.022396f
C254 VN.n54 B 0.044625f
C255 VN.n55 B 0.03128f
C256 VN.n56 B 0.703773f
C257 VN.n57 B 0.03128f
C258 VN.n58 B 0.022396f
C259 VN.n59 B 0.022396f
C260 VN.n60 B 0.022396f
C261 VN.n61 B 0.021116f
C262 VN.n62 B 0.040903f
C263 VN.n63 B 0.039481f
C264 VN.n64 B 0.022396f
C265 VN.n65 B 0.022396f
C266 VN.n66 B 0.023079f
C267 VN.n67 B 0.041532f
C268 VN.n68 B 0.035655f
C269 VN.n69 B 0.022396f
C270 VN.n70 B 0.022396f
C271 VN.n71 B 0.022396f
C272 VN.n72 B 0.041532f
C273 VN.n73 B 0.02718f
C274 VN.n74 B 0.76836f
C275 VN.n75 B 1.37145f
.ends

