* NGSPICE file created from diff_pair_sample_0554.ext - technology: sky130A

.subckt diff_pair_sample_0554 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t14 VN.t0 VDD2.t2 w_n2550_n2858# sky130_fd_pr__pfet_01v8 ad=3.6855 pd=19.68 as=1.55925 ps=9.78 w=9.45 l=1.25
X1 VTAIL.t5 VP.t0 VDD1.t7 w_n2550_n2858# sky130_fd_pr__pfet_01v8 ad=1.55925 pd=9.78 as=1.55925 ps=9.78 w=9.45 l=1.25
X2 VDD2.t1 VN.t1 VTAIL.t13 w_n2550_n2858# sky130_fd_pr__pfet_01v8 ad=1.55925 pd=9.78 as=1.55925 ps=9.78 w=9.45 l=1.25
X3 VDD1.t6 VP.t1 VTAIL.t15 w_n2550_n2858# sky130_fd_pr__pfet_01v8 ad=1.55925 pd=9.78 as=3.6855 ps=19.68 w=9.45 l=1.25
X4 VTAIL.t12 VN.t2 VDD2.t7 w_n2550_n2858# sky130_fd_pr__pfet_01v8 ad=1.55925 pd=9.78 as=1.55925 ps=9.78 w=9.45 l=1.25
X5 VTAIL.t6 VP.t2 VDD1.t5 w_n2550_n2858# sky130_fd_pr__pfet_01v8 ad=1.55925 pd=9.78 as=1.55925 ps=9.78 w=9.45 l=1.25
X6 VDD2.t5 VN.t3 VTAIL.t11 w_n2550_n2858# sky130_fd_pr__pfet_01v8 ad=1.55925 pd=9.78 as=3.6855 ps=19.68 w=9.45 l=1.25
X7 VTAIL.t10 VN.t4 VDD2.t0 w_n2550_n2858# sky130_fd_pr__pfet_01v8 ad=3.6855 pd=19.68 as=1.55925 ps=9.78 w=9.45 l=1.25
X8 VTAIL.t3 VP.t3 VDD1.t4 w_n2550_n2858# sky130_fd_pr__pfet_01v8 ad=3.6855 pd=19.68 as=1.55925 ps=9.78 w=9.45 l=1.25
X9 VDD2.t3 VN.t5 VTAIL.t9 w_n2550_n2858# sky130_fd_pr__pfet_01v8 ad=1.55925 pd=9.78 as=1.55925 ps=9.78 w=9.45 l=1.25
X10 VDD1.t3 VP.t4 VTAIL.t1 w_n2550_n2858# sky130_fd_pr__pfet_01v8 ad=1.55925 pd=9.78 as=3.6855 ps=19.68 w=9.45 l=1.25
X11 VDD2.t6 VN.t6 VTAIL.t8 w_n2550_n2858# sky130_fd_pr__pfet_01v8 ad=1.55925 pd=9.78 as=3.6855 ps=19.68 w=9.45 l=1.25
X12 VDD1.t2 VP.t5 VTAIL.t2 w_n2550_n2858# sky130_fd_pr__pfet_01v8 ad=1.55925 pd=9.78 as=1.55925 ps=9.78 w=9.45 l=1.25
X13 VDD1.t1 VP.t6 VTAIL.t4 w_n2550_n2858# sky130_fd_pr__pfet_01v8 ad=1.55925 pd=9.78 as=1.55925 ps=9.78 w=9.45 l=1.25
X14 B.t11 B.t9 B.t10 w_n2550_n2858# sky130_fd_pr__pfet_01v8 ad=3.6855 pd=19.68 as=0 ps=0 w=9.45 l=1.25
X15 VTAIL.t7 VN.t7 VDD2.t4 w_n2550_n2858# sky130_fd_pr__pfet_01v8 ad=1.55925 pd=9.78 as=1.55925 ps=9.78 w=9.45 l=1.25
X16 B.t8 B.t6 B.t7 w_n2550_n2858# sky130_fd_pr__pfet_01v8 ad=3.6855 pd=19.68 as=0 ps=0 w=9.45 l=1.25
X17 B.t5 B.t3 B.t4 w_n2550_n2858# sky130_fd_pr__pfet_01v8 ad=3.6855 pd=19.68 as=0 ps=0 w=9.45 l=1.25
X18 VTAIL.t0 VP.t7 VDD1.t0 w_n2550_n2858# sky130_fd_pr__pfet_01v8 ad=3.6855 pd=19.68 as=1.55925 ps=9.78 w=9.45 l=1.25
X19 B.t2 B.t0 B.t1 w_n2550_n2858# sky130_fd_pr__pfet_01v8 ad=3.6855 pd=19.68 as=0 ps=0 w=9.45 l=1.25
R0 VN.n4 VN.t4 233.855
R1 VN.n19 VN.t3 233.855
R2 VN.n13 VN.t6 213.815
R3 VN.n28 VN.t0 213.815
R4 VN.n3 VN.t5 182.196
R5 VN.n1 VN.t7 182.196
R6 VN.n18 VN.t2 182.196
R7 VN.n16 VN.t1 182.196
R8 VN.n27 VN.n15 161.3
R9 VN.n26 VN.n25 161.3
R10 VN.n24 VN.n23 161.3
R11 VN.n22 VN.n17 161.3
R12 VN.n21 VN.n20 161.3
R13 VN.n12 VN.n0 161.3
R14 VN.n11 VN.n10 161.3
R15 VN.n9 VN.n8 161.3
R16 VN.n7 VN.n2 161.3
R17 VN.n6 VN.n5 161.3
R18 VN.n29 VN.n28 80.6037
R19 VN.n14 VN.n13 80.6037
R20 VN.n4 VN.n3 43.2178
R21 VN.n19 VN.n18 43.2178
R22 VN VN.n29 43.1127
R23 VN.n7 VN.n6 40.4934
R24 VN.n8 VN.n7 40.4934
R25 VN.n22 VN.n21 40.4934
R26 VN.n23 VN.n22 40.4934
R27 VN.n13 VN.n12 35.7853
R28 VN.n28 VN.n27 35.7853
R29 VN.n12 VN.n11 32.7233
R30 VN.n27 VN.n26 32.7233
R31 VN.n20 VN.n19 29.2134
R32 VN.n5 VN.n4 29.2134
R33 VN.n6 VN.n3 14.1914
R34 VN.n8 VN.n1 14.1914
R35 VN.n21 VN.n18 14.1914
R36 VN.n23 VN.n16 14.1914
R37 VN.n11 VN.n1 10.2766
R38 VN.n26 VN.n16 10.2766
R39 VN.n29 VN.n15 0.285035
R40 VN.n14 VN.n0 0.285035
R41 VN.n25 VN.n15 0.189894
R42 VN.n25 VN.n24 0.189894
R43 VN.n24 VN.n17 0.189894
R44 VN.n20 VN.n17 0.189894
R45 VN.n5 VN.n2 0.189894
R46 VN.n9 VN.n2 0.189894
R47 VN.n10 VN.n9 0.189894
R48 VN.n10 VN.n0 0.189894
R49 VN VN.n14 0.146778
R50 VDD2.n2 VDD2.n1 83.2791
R51 VDD2.n2 VDD2.n0 83.2791
R52 VDD2 VDD2.n5 83.2763
R53 VDD2.n4 VDD2.n3 82.6536
R54 VDD2.n4 VDD2.n2 37.9912
R55 VDD2.n5 VDD2.t7 3.44018
R56 VDD2.n5 VDD2.t5 3.44018
R57 VDD2.n3 VDD2.t2 3.44018
R58 VDD2.n3 VDD2.t1 3.44018
R59 VDD2.n1 VDD2.t4 3.44018
R60 VDD2.n1 VDD2.t6 3.44018
R61 VDD2.n0 VDD2.t0 3.44018
R62 VDD2.n0 VDD2.t3 3.44018
R63 VDD2 VDD2.n4 0.739724
R64 VTAIL.n402 VTAIL.n358 756.745
R65 VTAIL.n46 VTAIL.n2 756.745
R66 VTAIL.n96 VTAIL.n52 756.745
R67 VTAIL.n148 VTAIL.n104 756.745
R68 VTAIL.n352 VTAIL.n308 756.745
R69 VTAIL.n300 VTAIL.n256 756.745
R70 VTAIL.n250 VTAIL.n206 756.745
R71 VTAIL.n198 VTAIL.n154 756.745
R72 VTAIL.n375 VTAIL.n374 585
R73 VTAIL.n377 VTAIL.n376 585
R74 VTAIL.n370 VTAIL.n369 585
R75 VTAIL.n383 VTAIL.n382 585
R76 VTAIL.n385 VTAIL.n384 585
R77 VTAIL.n366 VTAIL.n365 585
R78 VTAIL.n392 VTAIL.n391 585
R79 VTAIL.n393 VTAIL.n364 585
R80 VTAIL.n395 VTAIL.n394 585
R81 VTAIL.n362 VTAIL.n361 585
R82 VTAIL.n401 VTAIL.n400 585
R83 VTAIL.n403 VTAIL.n402 585
R84 VTAIL.n19 VTAIL.n18 585
R85 VTAIL.n21 VTAIL.n20 585
R86 VTAIL.n14 VTAIL.n13 585
R87 VTAIL.n27 VTAIL.n26 585
R88 VTAIL.n29 VTAIL.n28 585
R89 VTAIL.n10 VTAIL.n9 585
R90 VTAIL.n36 VTAIL.n35 585
R91 VTAIL.n37 VTAIL.n8 585
R92 VTAIL.n39 VTAIL.n38 585
R93 VTAIL.n6 VTAIL.n5 585
R94 VTAIL.n45 VTAIL.n44 585
R95 VTAIL.n47 VTAIL.n46 585
R96 VTAIL.n69 VTAIL.n68 585
R97 VTAIL.n71 VTAIL.n70 585
R98 VTAIL.n64 VTAIL.n63 585
R99 VTAIL.n77 VTAIL.n76 585
R100 VTAIL.n79 VTAIL.n78 585
R101 VTAIL.n60 VTAIL.n59 585
R102 VTAIL.n86 VTAIL.n85 585
R103 VTAIL.n87 VTAIL.n58 585
R104 VTAIL.n89 VTAIL.n88 585
R105 VTAIL.n56 VTAIL.n55 585
R106 VTAIL.n95 VTAIL.n94 585
R107 VTAIL.n97 VTAIL.n96 585
R108 VTAIL.n121 VTAIL.n120 585
R109 VTAIL.n123 VTAIL.n122 585
R110 VTAIL.n116 VTAIL.n115 585
R111 VTAIL.n129 VTAIL.n128 585
R112 VTAIL.n131 VTAIL.n130 585
R113 VTAIL.n112 VTAIL.n111 585
R114 VTAIL.n138 VTAIL.n137 585
R115 VTAIL.n139 VTAIL.n110 585
R116 VTAIL.n141 VTAIL.n140 585
R117 VTAIL.n108 VTAIL.n107 585
R118 VTAIL.n147 VTAIL.n146 585
R119 VTAIL.n149 VTAIL.n148 585
R120 VTAIL.n353 VTAIL.n352 585
R121 VTAIL.n351 VTAIL.n350 585
R122 VTAIL.n312 VTAIL.n311 585
R123 VTAIL.n316 VTAIL.n314 585
R124 VTAIL.n345 VTAIL.n344 585
R125 VTAIL.n343 VTAIL.n342 585
R126 VTAIL.n318 VTAIL.n317 585
R127 VTAIL.n337 VTAIL.n336 585
R128 VTAIL.n335 VTAIL.n334 585
R129 VTAIL.n322 VTAIL.n321 585
R130 VTAIL.n329 VTAIL.n328 585
R131 VTAIL.n327 VTAIL.n326 585
R132 VTAIL.n301 VTAIL.n300 585
R133 VTAIL.n299 VTAIL.n298 585
R134 VTAIL.n260 VTAIL.n259 585
R135 VTAIL.n264 VTAIL.n262 585
R136 VTAIL.n293 VTAIL.n292 585
R137 VTAIL.n291 VTAIL.n290 585
R138 VTAIL.n266 VTAIL.n265 585
R139 VTAIL.n285 VTAIL.n284 585
R140 VTAIL.n283 VTAIL.n282 585
R141 VTAIL.n270 VTAIL.n269 585
R142 VTAIL.n277 VTAIL.n276 585
R143 VTAIL.n275 VTAIL.n274 585
R144 VTAIL.n251 VTAIL.n250 585
R145 VTAIL.n249 VTAIL.n248 585
R146 VTAIL.n210 VTAIL.n209 585
R147 VTAIL.n214 VTAIL.n212 585
R148 VTAIL.n243 VTAIL.n242 585
R149 VTAIL.n241 VTAIL.n240 585
R150 VTAIL.n216 VTAIL.n215 585
R151 VTAIL.n235 VTAIL.n234 585
R152 VTAIL.n233 VTAIL.n232 585
R153 VTAIL.n220 VTAIL.n219 585
R154 VTAIL.n227 VTAIL.n226 585
R155 VTAIL.n225 VTAIL.n224 585
R156 VTAIL.n199 VTAIL.n198 585
R157 VTAIL.n197 VTAIL.n196 585
R158 VTAIL.n158 VTAIL.n157 585
R159 VTAIL.n162 VTAIL.n160 585
R160 VTAIL.n191 VTAIL.n190 585
R161 VTAIL.n189 VTAIL.n188 585
R162 VTAIL.n164 VTAIL.n163 585
R163 VTAIL.n183 VTAIL.n182 585
R164 VTAIL.n181 VTAIL.n180 585
R165 VTAIL.n168 VTAIL.n167 585
R166 VTAIL.n175 VTAIL.n174 585
R167 VTAIL.n173 VTAIL.n172 585
R168 VTAIL.n373 VTAIL.t8 329.038
R169 VTAIL.n17 VTAIL.t10 329.038
R170 VTAIL.n67 VTAIL.t1 329.038
R171 VTAIL.n119 VTAIL.t0 329.038
R172 VTAIL.n325 VTAIL.t15 329.038
R173 VTAIL.n273 VTAIL.t3 329.038
R174 VTAIL.n223 VTAIL.t11 329.038
R175 VTAIL.n171 VTAIL.t14 329.038
R176 VTAIL.n376 VTAIL.n375 171.744
R177 VTAIL.n376 VTAIL.n369 171.744
R178 VTAIL.n383 VTAIL.n369 171.744
R179 VTAIL.n384 VTAIL.n383 171.744
R180 VTAIL.n384 VTAIL.n365 171.744
R181 VTAIL.n392 VTAIL.n365 171.744
R182 VTAIL.n393 VTAIL.n392 171.744
R183 VTAIL.n394 VTAIL.n393 171.744
R184 VTAIL.n394 VTAIL.n361 171.744
R185 VTAIL.n401 VTAIL.n361 171.744
R186 VTAIL.n402 VTAIL.n401 171.744
R187 VTAIL.n20 VTAIL.n19 171.744
R188 VTAIL.n20 VTAIL.n13 171.744
R189 VTAIL.n27 VTAIL.n13 171.744
R190 VTAIL.n28 VTAIL.n27 171.744
R191 VTAIL.n28 VTAIL.n9 171.744
R192 VTAIL.n36 VTAIL.n9 171.744
R193 VTAIL.n37 VTAIL.n36 171.744
R194 VTAIL.n38 VTAIL.n37 171.744
R195 VTAIL.n38 VTAIL.n5 171.744
R196 VTAIL.n45 VTAIL.n5 171.744
R197 VTAIL.n46 VTAIL.n45 171.744
R198 VTAIL.n70 VTAIL.n69 171.744
R199 VTAIL.n70 VTAIL.n63 171.744
R200 VTAIL.n77 VTAIL.n63 171.744
R201 VTAIL.n78 VTAIL.n77 171.744
R202 VTAIL.n78 VTAIL.n59 171.744
R203 VTAIL.n86 VTAIL.n59 171.744
R204 VTAIL.n87 VTAIL.n86 171.744
R205 VTAIL.n88 VTAIL.n87 171.744
R206 VTAIL.n88 VTAIL.n55 171.744
R207 VTAIL.n95 VTAIL.n55 171.744
R208 VTAIL.n96 VTAIL.n95 171.744
R209 VTAIL.n122 VTAIL.n121 171.744
R210 VTAIL.n122 VTAIL.n115 171.744
R211 VTAIL.n129 VTAIL.n115 171.744
R212 VTAIL.n130 VTAIL.n129 171.744
R213 VTAIL.n130 VTAIL.n111 171.744
R214 VTAIL.n138 VTAIL.n111 171.744
R215 VTAIL.n139 VTAIL.n138 171.744
R216 VTAIL.n140 VTAIL.n139 171.744
R217 VTAIL.n140 VTAIL.n107 171.744
R218 VTAIL.n147 VTAIL.n107 171.744
R219 VTAIL.n148 VTAIL.n147 171.744
R220 VTAIL.n352 VTAIL.n351 171.744
R221 VTAIL.n351 VTAIL.n311 171.744
R222 VTAIL.n316 VTAIL.n311 171.744
R223 VTAIL.n344 VTAIL.n316 171.744
R224 VTAIL.n344 VTAIL.n343 171.744
R225 VTAIL.n343 VTAIL.n317 171.744
R226 VTAIL.n336 VTAIL.n317 171.744
R227 VTAIL.n336 VTAIL.n335 171.744
R228 VTAIL.n335 VTAIL.n321 171.744
R229 VTAIL.n328 VTAIL.n321 171.744
R230 VTAIL.n328 VTAIL.n327 171.744
R231 VTAIL.n300 VTAIL.n299 171.744
R232 VTAIL.n299 VTAIL.n259 171.744
R233 VTAIL.n264 VTAIL.n259 171.744
R234 VTAIL.n292 VTAIL.n264 171.744
R235 VTAIL.n292 VTAIL.n291 171.744
R236 VTAIL.n291 VTAIL.n265 171.744
R237 VTAIL.n284 VTAIL.n265 171.744
R238 VTAIL.n284 VTAIL.n283 171.744
R239 VTAIL.n283 VTAIL.n269 171.744
R240 VTAIL.n276 VTAIL.n269 171.744
R241 VTAIL.n276 VTAIL.n275 171.744
R242 VTAIL.n250 VTAIL.n249 171.744
R243 VTAIL.n249 VTAIL.n209 171.744
R244 VTAIL.n214 VTAIL.n209 171.744
R245 VTAIL.n242 VTAIL.n214 171.744
R246 VTAIL.n242 VTAIL.n241 171.744
R247 VTAIL.n241 VTAIL.n215 171.744
R248 VTAIL.n234 VTAIL.n215 171.744
R249 VTAIL.n234 VTAIL.n233 171.744
R250 VTAIL.n233 VTAIL.n219 171.744
R251 VTAIL.n226 VTAIL.n219 171.744
R252 VTAIL.n226 VTAIL.n225 171.744
R253 VTAIL.n198 VTAIL.n197 171.744
R254 VTAIL.n197 VTAIL.n157 171.744
R255 VTAIL.n162 VTAIL.n157 171.744
R256 VTAIL.n190 VTAIL.n162 171.744
R257 VTAIL.n190 VTAIL.n189 171.744
R258 VTAIL.n189 VTAIL.n163 171.744
R259 VTAIL.n182 VTAIL.n163 171.744
R260 VTAIL.n182 VTAIL.n181 171.744
R261 VTAIL.n181 VTAIL.n167 171.744
R262 VTAIL.n174 VTAIL.n167 171.744
R263 VTAIL.n174 VTAIL.n173 171.744
R264 VTAIL.n375 VTAIL.t8 85.8723
R265 VTAIL.n19 VTAIL.t10 85.8723
R266 VTAIL.n69 VTAIL.t1 85.8723
R267 VTAIL.n121 VTAIL.t0 85.8723
R268 VTAIL.n327 VTAIL.t15 85.8723
R269 VTAIL.n275 VTAIL.t3 85.8723
R270 VTAIL.n225 VTAIL.t11 85.8723
R271 VTAIL.n173 VTAIL.t14 85.8723
R272 VTAIL.n307 VTAIL.n306 65.9748
R273 VTAIL.n205 VTAIL.n204 65.9748
R274 VTAIL.n1 VTAIL.n0 65.9747
R275 VTAIL.n103 VTAIL.n102 65.9747
R276 VTAIL.n407 VTAIL.n406 36.2581
R277 VTAIL.n51 VTAIL.n50 36.2581
R278 VTAIL.n101 VTAIL.n100 36.2581
R279 VTAIL.n153 VTAIL.n152 36.2581
R280 VTAIL.n357 VTAIL.n356 36.2581
R281 VTAIL.n305 VTAIL.n304 36.2581
R282 VTAIL.n255 VTAIL.n254 36.2581
R283 VTAIL.n203 VTAIL.n202 36.2581
R284 VTAIL.n407 VTAIL.n357 21.8755
R285 VTAIL.n203 VTAIL.n153 21.8755
R286 VTAIL.n395 VTAIL.n362 13.1884
R287 VTAIL.n39 VTAIL.n6 13.1884
R288 VTAIL.n89 VTAIL.n56 13.1884
R289 VTAIL.n141 VTAIL.n108 13.1884
R290 VTAIL.n314 VTAIL.n312 13.1884
R291 VTAIL.n262 VTAIL.n260 13.1884
R292 VTAIL.n212 VTAIL.n210 13.1884
R293 VTAIL.n160 VTAIL.n158 13.1884
R294 VTAIL.n396 VTAIL.n364 12.8005
R295 VTAIL.n400 VTAIL.n399 12.8005
R296 VTAIL.n40 VTAIL.n8 12.8005
R297 VTAIL.n44 VTAIL.n43 12.8005
R298 VTAIL.n90 VTAIL.n58 12.8005
R299 VTAIL.n94 VTAIL.n93 12.8005
R300 VTAIL.n142 VTAIL.n110 12.8005
R301 VTAIL.n146 VTAIL.n145 12.8005
R302 VTAIL.n350 VTAIL.n349 12.8005
R303 VTAIL.n346 VTAIL.n345 12.8005
R304 VTAIL.n298 VTAIL.n297 12.8005
R305 VTAIL.n294 VTAIL.n293 12.8005
R306 VTAIL.n248 VTAIL.n247 12.8005
R307 VTAIL.n244 VTAIL.n243 12.8005
R308 VTAIL.n196 VTAIL.n195 12.8005
R309 VTAIL.n192 VTAIL.n191 12.8005
R310 VTAIL.n391 VTAIL.n390 12.0247
R311 VTAIL.n403 VTAIL.n360 12.0247
R312 VTAIL.n35 VTAIL.n34 12.0247
R313 VTAIL.n47 VTAIL.n4 12.0247
R314 VTAIL.n85 VTAIL.n84 12.0247
R315 VTAIL.n97 VTAIL.n54 12.0247
R316 VTAIL.n137 VTAIL.n136 12.0247
R317 VTAIL.n149 VTAIL.n106 12.0247
R318 VTAIL.n353 VTAIL.n310 12.0247
R319 VTAIL.n342 VTAIL.n315 12.0247
R320 VTAIL.n301 VTAIL.n258 12.0247
R321 VTAIL.n290 VTAIL.n263 12.0247
R322 VTAIL.n251 VTAIL.n208 12.0247
R323 VTAIL.n240 VTAIL.n213 12.0247
R324 VTAIL.n199 VTAIL.n156 12.0247
R325 VTAIL.n188 VTAIL.n161 12.0247
R326 VTAIL.n389 VTAIL.n366 11.249
R327 VTAIL.n404 VTAIL.n358 11.249
R328 VTAIL.n33 VTAIL.n10 11.249
R329 VTAIL.n48 VTAIL.n2 11.249
R330 VTAIL.n83 VTAIL.n60 11.249
R331 VTAIL.n98 VTAIL.n52 11.249
R332 VTAIL.n135 VTAIL.n112 11.249
R333 VTAIL.n150 VTAIL.n104 11.249
R334 VTAIL.n354 VTAIL.n308 11.249
R335 VTAIL.n341 VTAIL.n318 11.249
R336 VTAIL.n302 VTAIL.n256 11.249
R337 VTAIL.n289 VTAIL.n266 11.249
R338 VTAIL.n252 VTAIL.n206 11.249
R339 VTAIL.n239 VTAIL.n216 11.249
R340 VTAIL.n200 VTAIL.n154 11.249
R341 VTAIL.n187 VTAIL.n164 11.249
R342 VTAIL.n374 VTAIL.n373 10.7239
R343 VTAIL.n18 VTAIL.n17 10.7239
R344 VTAIL.n68 VTAIL.n67 10.7239
R345 VTAIL.n120 VTAIL.n119 10.7239
R346 VTAIL.n326 VTAIL.n325 10.7239
R347 VTAIL.n274 VTAIL.n273 10.7239
R348 VTAIL.n224 VTAIL.n223 10.7239
R349 VTAIL.n172 VTAIL.n171 10.7239
R350 VTAIL.n386 VTAIL.n385 10.4732
R351 VTAIL.n30 VTAIL.n29 10.4732
R352 VTAIL.n80 VTAIL.n79 10.4732
R353 VTAIL.n132 VTAIL.n131 10.4732
R354 VTAIL.n338 VTAIL.n337 10.4732
R355 VTAIL.n286 VTAIL.n285 10.4732
R356 VTAIL.n236 VTAIL.n235 10.4732
R357 VTAIL.n184 VTAIL.n183 10.4732
R358 VTAIL.n382 VTAIL.n368 9.69747
R359 VTAIL.n26 VTAIL.n12 9.69747
R360 VTAIL.n76 VTAIL.n62 9.69747
R361 VTAIL.n128 VTAIL.n114 9.69747
R362 VTAIL.n334 VTAIL.n320 9.69747
R363 VTAIL.n282 VTAIL.n268 9.69747
R364 VTAIL.n232 VTAIL.n218 9.69747
R365 VTAIL.n180 VTAIL.n166 9.69747
R366 VTAIL.n406 VTAIL.n405 9.45567
R367 VTAIL.n50 VTAIL.n49 9.45567
R368 VTAIL.n100 VTAIL.n99 9.45567
R369 VTAIL.n152 VTAIL.n151 9.45567
R370 VTAIL.n356 VTAIL.n355 9.45567
R371 VTAIL.n304 VTAIL.n303 9.45567
R372 VTAIL.n254 VTAIL.n253 9.45567
R373 VTAIL.n202 VTAIL.n201 9.45567
R374 VTAIL.n405 VTAIL.n404 9.3005
R375 VTAIL.n360 VTAIL.n359 9.3005
R376 VTAIL.n399 VTAIL.n398 9.3005
R377 VTAIL.n372 VTAIL.n371 9.3005
R378 VTAIL.n379 VTAIL.n378 9.3005
R379 VTAIL.n381 VTAIL.n380 9.3005
R380 VTAIL.n368 VTAIL.n367 9.3005
R381 VTAIL.n387 VTAIL.n386 9.3005
R382 VTAIL.n389 VTAIL.n388 9.3005
R383 VTAIL.n390 VTAIL.n363 9.3005
R384 VTAIL.n397 VTAIL.n396 9.3005
R385 VTAIL.n49 VTAIL.n48 9.3005
R386 VTAIL.n4 VTAIL.n3 9.3005
R387 VTAIL.n43 VTAIL.n42 9.3005
R388 VTAIL.n16 VTAIL.n15 9.3005
R389 VTAIL.n23 VTAIL.n22 9.3005
R390 VTAIL.n25 VTAIL.n24 9.3005
R391 VTAIL.n12 VTAIL.n11 9.3005
R392 VTAIL.n31 VTAIL.n30 9.3005
R393 VTAIL.n33 VTAIL.n32 9.3005
R394 VTAIL.n34 VTAIL.n7 9.3005
R395 VTAIL.n41 VTAIL.n40 9.3005
R396 VTAIL.n99 VTAIL.n98 9.3005
R397 VTAIL.n54 VTAIL.n53 9.3005
R398 VTAIL.n93 VTAIL.n92 9.3005
R399 VTAIL.n66 VTAIL.n65 9.3005
R400 VTAIL.n73 VTAIL.n72 9.3005
R401 VTAIL.n75 VTAIL.n74 9.3005
R402 VTAIL.n62 VTAIL.n61 9.3005
R403 VTAIL.n81 VTAIL.n80 9.3005
R404 VTAIL.n83 VTAIL.n82 9.3005
R405 VTAIL.n84 VTAIL.n57 9.3005
R406 VTAIL.n91 VTAIL.n90 9.3005
R407 VTAIL.n151 VTAIL.n150 9.3005
R408 VTAIL.n106 VTAIL.n105 9.3005
R409 VTAIL.n145 VTAIL.n144 9.3005
R410 VTAIL.n118 VTAIL.n117 9.3005
R411 VTAIL.n125 VTAIL.n124 9.3005
R412 VTAIL.n127 VTAIL.n126 9.3005
R413 VTAIL.n114 VTAIL.n113 9.3005
R414 VTAIL.n133 VTAIL.n132 9.3005
R415 VTAIL.n135 VTAIL.n134 9.3005
R416 VTAIL.n136 VTAIL.n109 9.3005
R417 VTAIL.n143 VTAIL.n142 9.3005
R418 VTAIL.n324 VTAIL.n323 9.3005
R419 VTAIL.n331 VTAIL.n330 9.3005
R420 VTAIL.n333 VTAIL.n332 9.3005
R421 VTAIL.n320 VTAIL.n319 9.3005
R422 VTAIL.n339 VTAIL.n338 9.3005
R423 VTAIL.n341 VTAIL.n340 9.3005
R424 VTAIL.n315 VTAIL.n313 9.3005
R425 VTAIL.n347 VTAIL.n346 9.3005
R426 VTAIL.n355 VTAIL.n354 9.3005
R427 VTAIL.n310 VTAIL.n309 9.3005
R428 VTAIL.n349 VTAIL.n348 9.3005
R429 VTAIL.n272 VTAIL.n271 9.3005
R430 VTAIL.n279 VTAIL.n278 9.3005
R431 VTAIL.n281 VTAIL.n280 9.3005
R432 VTAIL.n268 VTAIL.n267 9.3005
R433 VTAIL.n287 VTAIL.n286 9.3005
R434 VTAIL.n289 VTAIL.n288 9.3005
R435 VTAIL.n263 VTAIL.n261 9.3005
R436 VTAIL.n295 VTAIL.n294 9.3005
R437 VTAIL.n303 VTAIL.n302 9.3005
R438 VTAIL.n258 VTAIL.n257 9.3005
R439 VTAIL.n297 VTAIL.n296 9.3005
R440 VTAIL.n222 VTAIL.n221 9.3005
R441 VTAIL.n229 VTAIL.n228 9.3005
R442 VTAIL.n231 VTAIL.n230 9.3005
R443 VTAIL.n218 VTAIL.n217 9.3005
R444 VTAIL.n237 VTAIL.n236 9.3005
R445 VTAIL.n239 VTAIL.n238 9.3005
R446 VTAIL.n213 VTAIL.n211 9.3005
R447 VTAIL.n245 VTAIL.n244 9.3005
R448 VTAIL.n253 VTAIL.n252 9.3005
R449 VTAIL.n208 VTAIL.n207 9.3005
R450 VTAIL.n247 VTAIL.n246 9.3005
R451 VTAIL.n170 VTAIL.n169 9.3005
R452 VTAIL.n177 VTAIL.n176 9.3005
R453 VTAIL.n179 VTAIL.n178 9.3005
R454 VTAIL.n166 VTAIL.n165 9.3005
R455 VTAIL.n185 VTAIL.n184 9.3005
R456 VTAIL.n187 VTAIL.n186 9.3005
R457 VTAIL.n161 VTAIL.n159 9.3005
R458 VTAIL.n193 VTAIL.n192 9.3005
R459 VTAIL.n201 VTAIL.n200 9.3005
R460 VTAIL.n156 VTAIL.n155 9.3005
R461 VTAIL.n195 VTAIL.n194 9.3005
R462 VTAIL.n381 VTAIL.n370 8.92171
R463 VTAIL.n25 VTAIL.n14 8.92171
R464 VTAIL.n75 VTAIL.n64 8.92171
R465 VTAIL.n127 VTAIL.n116 8.92171
R466 VTAIL.n333 VTAIL.n322 8.92171
R467 VTAIL.n281 VTAIL.n270 8.92171
R468 VTAIL.n231 VTAIL.n220 8.92171
R469 VTAIL.n179 VTAIL.n168 8.92171
R470 VTAIL.n378 VTAIL.n377 8.14595
R471 VTAIL.n22 VTAIL.n21 8.14595
R472 VTAIL.n72 VTAIL.n71 8.14595
R473 VTAIL.n124 VTAIL.n123 8.14595
R474 VTAIL.n330 VTAIL.n329 8.14595
R475 VTAIL.n278 VTAIL.n277 8.14595
R476 VTAIL.n228 VTAIL.n227 8.14595
R477 VTAIL.n176 VTAIL.n175 8.14595
R478 VTAIL.n374 VTAIL.n372 7.3702
R479 VTAIL.n18 VTAIL.n16 7.3702
R480 VTAIL.n68 VTAIL.n66 7.3702
R481 VTAIL.n120 VTAIL.n118 7.3702
R482 VTAIL.n326 VTAIL.n324 7.3702
R483 VTAIL.n274 VTAIL.n272 7.3702
R484 VTAIL.n224 VTAIL.n222 7.3702
R485 VTAIL.n172 VTAIL.n170 7.3702
R486 VTAIL.n377 VTAIL.n372 5.81868
R487 VTAIL.n21 VTAIL.n16 5.81868
R488 VTAIL.n71 VTAIL.n66 5.81868
R489 VTAIL.n123 VTAIL.n118 5.81868
R490 VTAIL.n329 VTAIL.n324 5.81868
R491 VTAIL.n277 VTAIL.n272 5.81868
R492 VTAIL.n227 VTAIL.n222 5.81868
R493 VTAIL.n175 VTAIL.n170 5.81868
R494 VTAIL.n378 VTAIL.n370 5.04292
R495 VTAIL.n22 VTAIL.n14 5.04292
R496 VTAIL.n72 VTAIL.n64 5.04292
R497 VTAIL.n124 VTAIL.n116 5.04292
R498 VTAIL.n330 VTAIL.n322 5.04292
R499 VTAIL.n278 VTAIL.n270 5.04292
R500 VTAIL.n228 VTAIL.n220 5.04292
R501 VTAIL.n176 VTAIL.n168 5.04292
R502 VTAIL.n382 VTAIL.n381 4.26717
R503 VTAIL.n26 VTAIL.n25 4.26717
R504 VTAIL.n76 VTAIL.n75 4.26717
R505 VTAIL.n128 VTAIL.n127 4.26717
R506 VTAIL.n334 VTAIL.n333 4.26717
R507 VTAIL.n282 VTAIL.n281 4.26717
R508 VTAIL.n232 VTAIL.n231 4.26717
R509 VTAIL.n180 VTAIL.n179 4.26717
R510 VTAIL.n385 VTAIL.n368 3.49141
R511 VTAIL.n29 VTAIL.n12 3.49141
R512 VTAIL.n79 VTAIL.n62 3.49141
R513 VTAIL.n131 VTAIL.n114 3.49141
R514 VTAIL.n337 VTAIL.n320 3.49141
R515 VTAIL.n285 VTAIL.n268 3.49141
R516 VTAIL.n235 VTAIL.n218 3.49141
R517 VTAIL.n183 VTAIL.n166 3.49141
R518 VTAIL.n0 VTAIL.t9 3.44018
R519 VTAIL.n0 VTAIL.t7 3.44018
R520 VTAIL.n102 VTAIL.t4 3.44018
R521 VTAIL.n102 VTAIL.t5 3.44018
R522 VTAIL.n306 VTAIL.t2 3.44018
R523 VTAIL.n306 VTAIL.t6 3.44018
R524 VTAIL.n204 VTAIL.t13 3.44018
R525 VTAIL.n204 VTAIL.t12 3.44018
R526 VTAIL.n386 VTAIL.n366 2.71565
R527 VTAIL.n406 VTAIL.n358 2.71565
R528 VTAIL.n30 VTAIL.n10 2.71565
R529 VTAIL.n50 VTAIL.n2 2.71565
R530 VTAIL.n80 VTAIL.n60 2.71565
R531 VTAIL.n100 VTAIL.n52 2.71565
R532 VTAIL.n132 VTAIL.n112 2.71565
R533 VTAIL.n152 VTAIL.n104 2.71565
R534 VTAIL.n356 VTAIL.n308 2.71565
R535 VTAIL.n338 VTAIL.n318 2.71565
R536 VTAIL.n304 VTAIL.n256 2.71565
R537 VTAIL.n286 VTAIL.n266 2.71565
R538 VTAIL.n254 VTAIL.n206 2.71565
R539 VTAIL.n236 VTAIL.n216 2.71565
R540 VTAIL.n202 VTAIL.n154 2.71565
R541 VTAIL.n184 VTAIL.n164 2.71565
R542 VTAIL.n373 VTAIL.n371 2.41283
R543 VTAIL.n17 VTAIL.n15 2.41283
R544 VTAIL.n67 VTAIL.n65 2.41283
R545 VTAIL.n119 VTAIL.n117 2.41283
R546 VTAIL.n325 VTAIL.n323 2.41283
R547 VTAIL.n273 VTAIL.n271 2.41283
R548 VTAIL.n223 VTAIL.n221 2.41283
R549 VTAIL.n171 VTAIL.n169 2.41283
R550 VTAIL.n391 VTAIL.n389 1.93989
R551 VTAIL.n404 VTAIL.n403 1.93989
R552 VTAIL.n35 VTAIL.n33 1.93989
R553 VTAIL.n48 VTAIL.n47 1.93989
R554 VTAIL.n85 VTAIL.n83 1.93989
R555 VTAIL.n98 VTAIL.n97 1.93989
R556 VTAIL.n137 VTAIL.n135 1.93989
R557 VTAIL.n150 VTAIL.n149 1.93989
R558 VTAIL.n354 VTAIL.n353 1.93989
R559 VTAIL.n342 VTAIL.n341 1.93989
R560 VTAIL.n302 VTAIL.n301 1.93989
R561 VTAIL.n290 VTAIL.n289 1.93989
R562 VTAIL.n252 VTAIL.n251 1.93989
R563 VTAIL.n240 VTAIL.n239 1.93989
R564 VTAIL.n200 VTAIL.n199 1.93989
R565 VTAIL.n188 VTAIL.n187 1.93989
R566 VTAIL.n205 VTAIL.n203 1.36257
R567 VTAIL.n255 VTAIL.n205 1.36257
R568 VTAIL.n307 VTAIL.n305 1.36257
R569 VTAIL.n357 VTAIL.n307 1.36257
R570 VTAIL.n153 VTAIL.n103 1.36257
R571 VTAIL.n103 VTAIL.n101 1.36257
R572 VTAIL.n51 VTAIL.n1 1.36257
R573 VTAIL VTAIL.n407 1.30438
R574 VTAIL.n390 VTAIL.n364 1.16414
R575 VTAIL.n400 VTAIL.n360 1.16414
R576 VTAIL.n34 VTAIL.n8 1.16414
R577 VTAIL.n44 VTAIL.n4 1.16414
R578 VTAIL.n84 VTAIL.n58 1.16414
R579 VTAIL.n94 VTAIL.n54 1.16414
R580 VTAIL.n136 VTAIL.n110 1.16414
R581 VTAIL.n146 VTAIL.n106 1.16414
R582 VTAIL.n350 VTAIL.n310 1.16414
R583 VTAIL.n345 VTAIL.n315 1.16414
R584 VTAIL.n298 VTAIL.n258 1.16414
R585 VTAIL.n293 VTAIL.n263 1.16414
R586 VTAIL.n248 VTAIL.n208 1.16414
R587 VTAIL.n243 VTAIL.n213 1.16414
R588 VTAIL.n196 VTAIL.n156 1.16414
R589 VTAIL.n191 VTAIL.n161 1.16414
R590 VTAIL.n305 VTAIL.n255 0.470328
R591 VTAIL.n101 VTAIL.n51 0.470328
R592 VTAIL.n396 VTAIL.n395 0.388379
R593 VTAIL.n399 VTAIL.n362 0.388379
R594 VTAIL.n40 VTAIL.n39 0.388379
R595 VTAIL.n43 VTAIL.n6 0.388379
R596 VTAIL.n90 VTAIL.n89 0.388379
R597 VTAIL.n93 VTAIL.n56 0.388379
R598 VTAIL.n142 VTAIL.n141 0.388379
R599 VTAIL.n145 VTAIL.n108 0.388379
R600 VTAIL.n349 VTAIL.n312 0.388379
R601 VTAIL.n346 VTAIL.n314 0.388379
R602 VTAIL.n297 VTAIL.n260 0.388379
R603 VTAIL.n294 VTAIL.n262 0.388379
R604 VTAIL.n247 VTAIL.n210 0.388379
R605 VTAIL.n244 VTAIL.n212 0.388379
R606 VTAIL.n195 VTAIL.n158 0.388379
R607 VTAIL.n192 VTAIL.n160 0.388379
R608 VTAIL.n379 VTAIL.n371 0.155672
R609 VTAIL.n380 VTAIL.n379 0.155672
R610 VTAIL.n380 VTAIL.n367 0.155672
R611 VTAIL.n387 VTAIL.n367 0.155672
R612 VTAIL.n388 VTAIL.n387 0.155672
R613 VTAIL.n388 VTAIL.n363 0.155672
R614 VTAIL.n397 VTAIL.n363 0.155672
R615 VTAIL.n398 VTAIL.n397 0.155672
R616 VTAIL.n398 VTAIL.n359 0.155672
R617 VTAIL.n405 VTAIL.n359 0.155672
R618 VTAIL.n23 VTAIL.n15 0.155672
R619 VTAIL.n24 VTAIL.n23 0.155672
R620 VTAIL.n24 VTAIL.n11 0.155672
R621 VTAIL.n31 VTAIL.n11 0.155672
R622 VTAIL.n32 VTAIL.n31 0.155672
R623 VTAIL.n32 VTAIL.n7 0.155672
R624 VTAIL.n41 VTAIL.n7 0.155672
R625 VTAIL.n42 VTAIL.n41 0.155672
R626 VTAIL.n42 VTAIL.n3 0.155672
R627 VTAIL.n49 VTAIL.n3 0.155672
R628 VTAIL.n73 VTAIL.n65 0.155672
R629 VTAIL.n74 VTAIL.n73 0.155672
R630 VTAIL.n74 VTAIL.n61 0.155672
R631 VTAIL.n81 VTAIL.n61 0.155672
R632 VTAIL.n82 VTAIL.n81 0.155672
R633 VTAIL.n82 VTAIL.n57 0.155672
R634 VTAIL.n91 VTAIL.n57 0.155672
R635 VTAIL.n92 VTAIL.n91 0.155672
R636 VTAIL.n92 VTAIL.n53 0.155672
R637 VTAIL.n99 VTAIL.n53 0.155672
R638 VTAIL.n125 VTAIL.n117 0.155672
R639 VTAIL.n126 VTAIL.n125 0.155672
R640 VTAIL.n126 VTAIL.n113 0.155672
R641 VTAIL.n133 VTAIL.n113 0.155672
R642 VTAIL.n134 VTAIL.n133 0.155672
R643 VTAIL.n134 VTAIL.n109 0.155672
R644 VTAIL.n143 VTAIL.n109 0.155672
R645 VTAIL.n144 VTAIL.n143 0.155672
R646 VTAIL.n144 VTAIL.n105 0.155672
R647 VTAIL.n151 VTAIL.n105 0.155672
R648 VTAIL.n355 VTAIL.n309 0.155672
R649 VTAIL.n348 VTAIL.n309 0.155672
R650 VTAIL.n348 VTAIL.n347 0.155672
R651 VTAIL.n347 VTAIL.n313 0.155672
R652 VTAIL.n340 VTAIL.n313 0.155672
R653 VTAIL.n340 VTAIL.n339 0.155672
R654 VTAIL.n339 VTAIL.n319 0.155672
R655 VTAIL.n332 VTAIL.n319 0.155672
R656 VTAIL.n332 VTAIL.n331 0.155672
R657 VTAIL.n331 VTAIL.n323 0.155672
R658 VTAIL.n303 VTAIL.n257 0.155672
R659 VTAIL.n296 VTAIL.n257 0.155672
R660 VTAIL.n296 VTAIL.n295 0.155672
R661 VTAIL.n295 VTAIL.n261 0.155672
R662 VTAIL.n288 VTAIL.n261 0.155672
R663 VTAIL.n288 VTAIL.n287 0.155672
R664 VTAIL.n287 VTAIL.n267 0.155672
R665 VTAIL.n280 VTAIL.n267 0.155672
R666 VTAIL.n280 VTAIL.n279 0.155672
R667 VTAIL.n279 VTAIL.n271 0.155672
R668 VTAIL.n253 VTAIL.n207 0.155672
R669 VTAIL.n246 VTAIL.n207 0.155672
R670 VTAIL.n246 VTAIL.n245 0.155672
R671 VTAIL.n245 VTAIL.n211 0.155672
R672 VTAIL.n238 VTAIL.n211 0.155672
R673 VTAIL.n238 VTAIL.n237 0.155672
R674 VTAIL.n237 VTAIL.n217 0.155672
R675 VTAIL.n230 VTAIL.n217 0.155672
R676 VTAIL.n230 VTAIL.n229 0.155672
R677 VTAIL.n229 VTAIL.n221 0.155672
R678 VTAIL.n201 VTAIL.n155 0.155672
R679 VTAIL.n194 VTAIL.n155 0.155672
R680 VTAIL.n194 VTAIL.n193 0.155672
R681 VTAIL.n193 VTAIL.n159 0.155672
R682 VTAIL.n186 VTAIL.n159 0.155672
R683 VTAIL.n186 VTAIL.n185 0.155672
R684 VTAIL.n185 VTAIL.n165 0.155672
R685 VTAIL.n178 VTAIL.n165 0.155672
R686 VTAIL.n178 VTAIL.n177 0.155672
R687 VTAIL.n177 VTAIL.n169 0.155672
R688 VTAIL VTAIL.n1 0.0586897
R689 VP.n9 VP.t3 233.855
R690 VP.n21 VP.t7 213.815
R691 VP.n33 VP.t4 213.815
R692 VP.n18 VP.t1 213.815
R693 VP.n3 VP.t6 182.196
R694 VP.n1 VP.t0 182.196
R695 VP.n6 VP.t2 182.196
R696 VP.n8 VP.t5 182.196
R697 VP.n11 VP.n10 161.3
R698 VP.n12 VP.n7 161.3
R699 VP.n14 VP.n13 161.3
R700 VP.n16 VP.n15 161.3
R701 VP.n17 VP.n5 161.3
R702 VP.n32 VP.n0 161.3
R703 VP.n31 VP.n30 161.3
R704 VP.n29 VP.n28 161.3
R705 VP.n27 VP.n2 161.3
R706 VP.n26 VP.n25 161.3
R707 VP.n24 VP.n23 161.3
R708 VP.n22 VP.n4 161.3
R709 VP.n19 VP.n18 80.6037
R710 VP.n34 VP.n33 80.6037
R711 VP.n21 VP.n20 80.6037
R712 VP.n9 VP.n8 43.2178
R713 VP.n20 VP.n19 42.8271
R714 VP.n27 VP.n26 40.4934
R715 VP.n28 VP.n27 40.4934
R716 VP.n13 VP.n12 40.4934
R717 VP.n12 VP.n11 40.4934
R718 VP.n22 VP.n21 35.7853
R719 VP.n33 VP.n32 35.7853
R720 VP.n18 VP.n17 35.7853
R721 VP.n23 VP.n22 32.7233
R722 VP.n32 VP.n31 32.7233
R723 VP.n17 VP.n16 32.7233
R724 VP.n10 VP.n9 29.2134
R725 VP.n26 VP.n3 14.1914
R726 VP.n28 VP.n1 14.1914
R727 VP.n13 VP.n6 14.1914
R728 VP.n11 VP.n8 14.1914
R729 VP.n23 VP.n3 10.2766
R730 VP.n31 VP.n1 10.2766
R731 VP.n16 VP.n6 10.2766
R732 VP.n19 VP.n5 0.285035
R733 VP.n20 VP.n4 0.285035
R734 VP.n34 VP.n0 0.285035
R735 VP.n10 VP.n7 0.189894
R736 VP.n14 VP.n7 0.189894
R737 VP.n15 VP.n14 0.189894
R738 VP.n15 VP.n5 0.189894
R739 VP.n24 VP.n4 0.189894
R740 VP.n25 VP.n24 0.189894
R741 VP.n25 VP.n2 0.189894
R742 VP.n29 VP.n2 0.189894
R743 VP.n30 VP.n29 0.189894
R744 VP.n30 VP.n0 0.189894
R745 VP VP.n34 0.146778
R746 VDD1 VDD1.n0 83.3928
R747 VDD1.n3 VDD1.n2 83.2791
R748 VDD1.n3 VDD1.n1 83.2791
R749 VDD1.n5 VDD1.n4 82.6534
R750 VDD1.n5 VDD1.n3 38.5742
R751 VDD1.n4 VDD1.t5 3.44018
R752 VDD1.n4 VDD1.t6 3.44018
R753 VDD1.n0 VDD1.t4 3.44018
R754 VDD1.n0 VDD1.t2 3.44018
R755 VDD1.n2 VDD1.t7 3.44018
R756 VDD1.n2 VDD1.t3 3.44018
R757 VDD1.n1 VDD1.t0 3.44018
R758 VDD1.n1 VDD1.t1 3.44018
R759 VDD1 VDD1.n5 0.623345
R760 B.n315 B.n314 585
R761 B.n313 B.n94 585
R762 B.n312 B.n311 585
R763 B.n310 B.n95 585
R764 B.n309 B.n308 585
R765 B.n307 B.n96 585
R766 B.n306 B.n305 585
R767 B.n304 B.n97 585
R768 B.n303 B.n302 585
R769 B.n301 B.n98 585
R770 B.n300 B.n299 585
R771 B.n298 B.n99 585
R772 B.n297 B.n296 585
R773 B.n295 B.n100 585
R774 B.n294 B.n293 585
R775 B.n292 B.n101 585
R776 B.n291 B.n290 585
R777 B.n289 B.n102 585
R778 B.n288 B.n287 585
R779 B.n286 B.n103 585
R780 B.n285 B.n284 585
R781 B.n283 B.n104 585
R782 B.n282 B.n281 585
R783 B.n280 B.n105 585
R784 B.n279 B.n278 585
R785 B.n277 B.n106 585
R786 B.n276 B.n275 585
R787 B.n274 B.n107 585
R788 B.n273 B.n272 585
R789 B.n271 B.n108 585
R790 B.n270 B.n269 585
R791 B.n268 B.n109 585
R792 B.n267 B.n266 585
R793 B.n265 B.n110 585
R794 B.n263 B.n262 585
R795 B.n261 B.n113 585
R796 B.n260 B.n259 585
R797 B.n258 B.n114 585
R798 B.n257 B.n256 585
R799 B.n255 B.n115 585
R800 B.n254 B.n253 585
R801 B.n252 B.n116 585
R802 B.n251 B.n250 585
R803 B.n249 B.n117 585
R804 B.n248 B.n247 585
R805 B.n243 B.n118 585
R806 B.n242 B.n241 585
R807 B.n240 B.n119 585
R808 B.n239 B.n238 585
R809 B.n237 B.n120 585
R810 B.n236 B.n235 585
R811 B.n234 B.n121 585
R812 B.n233 B.n232 585
R813 B.n231 B.n122 585
R814 B.n230 B.n229 585
R815 B.n228 B.n123 585
R816 B.n227 B.n226 585
R817 B.n225 B.n124 585
R818 B.n224 B.n223 585
R819 B.n222 B.n125 585
R820 B.n221 B.n220 585
R821 B.n219 B.n126 585
R822 B.n218 B.n217 585
R823 B.n216 B.n127 585
R824 B.n215 B.n214 585
R825 B.n213 B.n128 585
R826 B.n212 B.n211 585
R827 B.n210 B.n129 585
R828 B.n209 B.n208 585
R829 B.n207 B.n130 585
R830 B.n206 B.n205 585
R831 B.n204 B.n131 585
R832 B.n203 B.n202 585
R833 B.n201 B.n132 585
R834 B.n200 B.n199 585
R835 B.n198 B.n133 585
R836 B.n197 B.n196 585
R837 B.n195 B.n134 585
R838 B.n316 B.n93 585
R839 B.n318 B.n317 585
R840 B.n319 B.n92 585
R841 B.n321 B.n320 585
R842 B.n322 B.n91 585
R843 B.n324 B.n323 585
R844 B.n325 B.n90 585
R845 B.n327 B.n326 585
R846 B.n328 B.n89 585
R847 B.n330 B.n329 585
R848 B.n331 B.n88 585
R849 B.n333 B.n332 585
R850 B.n334 B.n87 585
R851 B.n336 B.n335 585
R852 B.n337 B.n86 585
R853 B.n339 B.n338 585
R854 B.n340 B.n85 585
R855 B.n342 B.n341 585
R856 B.n343 B.n84 585
R857 B.n345 B.n344 585
R858 B.n346 B.n83 585
R859 B.n348 B.n347 585
R860 B.n349 B.n82 585
R861 B.n351 B.n350 585
R862 B.n352 B.n81 585
R863 B.n354 B.n353 585
R864 B.n355 B.n80 585
R865 B.n357 B.n356 585
R866 B.n358 B.n79 585
R867 B.n360 B.n359 585
R868 B.n361 B.n78 585
R869 B.n363 B.n362 585
R870 B.n364 B.n77 585
R871 B.n366 B.n365 585
R872 B.n367 B.n76 585
R873 B.n369 B.n368 585
R874 B.n370 B.n75 585
R875 B.n372 B.n371 585
R876 B.n373 B.n74 585
R877 B.n375 B.n374 585
R878 B.n376 B.n73 585
R879 B.n378 B.n377 585
R880 B.n379 B.n72 585
R881 B.n381 B.n380 585
R882 B.n382 B.n71 585
R883 B.n384 B.n383 585
R884 B.n385 B.n70 585
R885 B.n387 B.n386 585
R886 B.n388 B.n69 585
R887 B.n390 B.n389 585
R888 B.n391 B.n68 585
R889 B.n393 B.n392 585
R890 B.n394 B.n67 585
R891 B.n396 B.n395 585
R892 B.n397 B.n66 585
R893 B.n399 B.n398 585
R894 B.n400 B.n65 585
R895 B.n402 B.n401 585
R896 B.n403 B.n64 585
R897 B.n405 B.n404 585
R898 B.n406 B.n63 585
R899 B.n408 B.n407 585
R900 B.n409 B.n62 585
R901 B.n411 B.n410 585
R902 B.n529 B.n528 585
R903 B.n527 B.n18 585
R904 B.n526 B.n525 585
R905 B.n524 B.n19 585
R906 B.n523 B.n522 585
R907 B.n521 B.n20 585
R908 B.n520 B.n519 585
R909 B.n518 B.n21 585
R910 B.n517 B.n516 585
R911 B.n515 B.n22 585
R912 B.n514 B.n513 585
R913 B.n512 B.n23 585
R914 B.n511 B.n510 585
R915 B.n509 B.n24 585
R916 B.n508 B.n507 585
R917 B.n506 B.n25 585
R918 B.n505 B.n504 585
R919 B.n503 B.n26 585
R920 B.n502 B.n501 585
R921 B.n500 B.n27 585
R922 B.n499 B.n498 585
R923 B.n497 B.n28 585
R924 B.n496 B.n495 585
R925 B.n494 B.n29 585
R926 B.n493 B.n492 585
R927 B.n491 B.n30 585
R928 B.n490 B.n489 585
R929 B.n488 B.n31 585
R930 B.n487 B.n486 585
R931 B.n485 B.n32 585
R932 B.n484 B.n483 585
R933 B.n482 B.n33 585
R934 B.n481 B.n480 585
R935 B.n479 B.n34 585
R936 B.n478 B.n477 585
R937 B.n476 B.n35 585
R938 B.n475 B.n474 585
R939 B.n473 B.n39 585
R940 B.n472 B.n471 585
R941 B.n470 B.n40 585
R942 B.n469 B.n468 585
R943 B.n467 B.n41 585
R944 B.n466 B.n465 585
R945 B.n464 B.n42 585
R946 B.n462 B.n461 585
R947 B.n460 B.n45 585
R948 B.n459 B.n458 585
R949 B.n457 B.n46 585
R950 B.n456 B.n455 585
R951 B.n454 B.n47 585
R952 B.n453 B.n452 585
R953 B.n451 B.n48 585
R954 B.n450 B.n449 585
R955 B.n448 B.n49 585
R956 B.n447 B.n446 585
R957 B.n445 B.n50 585
R958 B.n444 B.n443 585
R959 B.n442 B.n51 585
R960 B.n441 B.n440 585
R961 B.n439 B.n52 585
R962 B.n438 B.n437 585
R963 B.n436 B.n53 585
R964 B.n435 B.n434 585
R965 B.n433 B.n54 585
R966 B.n432 B.n431 585
R967 B.n430 B.n55 585
R968 B.n429 B.n428 585
R969 B.n427 B.n56 585
R970 B.n426 B.n425 585
R971 B.n424 B.n57 585
R972 B.n423 B.n422 585
R973 B.n421 B.n58 585
R974 B.n420 B.n419 585
R975 B.n418 B.n59 585
R976 B.n417 B.n416 585
R977 B.n415 B.n60 585
R978 B.n414 B.n413 585
R979 B.n412 B.n61 585
R980 B.n530 B.n17 585
R981 B.n532 B.n531 585
R982 B.n533 B.n16 585
R983 B.n535 B.n534 585
R984 B.n536 B.n15 585
R985 B.n538 B.n537 585
R986 B.n539 B.n14 585
R987 B.n541 B.n540 585
R988 B.n542 B.n13 585
R989 B.n544 B.n543 585
R990 B.n545 B.n12 585
R991 B.n547 B.n546 585
R992 B.n548 B.n11 585
R993 B.n550 B.n549 585
R994 B.n551 B.n10 585
R995 B.n553 B.n552 585
R996 B.n554 B.n9 585
R997 B.n556 B.n555 585
R998 B.n557 B.n8 585
R999 B.n559 B.n558 585
R1000 B.n560 B.n7 585
R1001 B.n562 B.n561 585
R1002 B.n563 B.n6 585
R1003 B.n565 B.n564 585
R1004 B.n566 B.n5 585
R1005 B.n568 B.n567 585
R1006 B.n569 B.n4 585
R1007 B.n571 B.n570 585
R1008 B.n572 B.n3 585
R1009 B.n574 B.n573 585
R1010 B.n575 B.n0 585
R1011 B.n2 B.n1 585
R1012 B.n150 B.n149 585
R1013 B.n152 B.n151 585
R1014 B.n153 B.n148 585
R1015 B.n155 B.n154 585
R1016 B.n156 B.n147 585
R1017 B.n158 B.n157 585
R1018 B.n159 B.n146 585
R1019 B.n161 B.n160 585
R1020 B.n162 B.n145 585
R1021 B.n164 B.n163 585
R1022 B.n165 B.n144 585
R1023 B.n167 B.n166 585
R1024 B.n168 B.n143 585
R1025 B.n170 B.n169 585
R1026 B.n171 B.n142 585
R1027 B.n173 B.n172 585
R1028 B.n174 B.n141 585
R1029 B.n176 B.n175 585
R1030 B.n177 B.n140 585
R1031 B.n179 B.n178 585
R1032 B.n180 B.n139 585
R1033 B.n182 B.n181 585
R1034 B.n183 B.n138 585
R1035 B.n185 B.n184 585
R1036 B.n186 B.n137 585
R1037 B.n188 B.n187 585
R1038 B.n189 B.n136 585
R1039 B.n191 B.n190 585
R1040 B.n192 B.n135 585
R1041 B.n194 B.n193 585
R1042 B.n193 B.n134 458.866
R1043 B.n316 B.n315 458.866
R1044 B.n412 B.n411 458.866
R1045 B.n528 B.n17 458.866
R1046 B.n244 B.t9 386.567
R1047 B.n111 B.t0 386.567
R1048 B.n43 B.t6 386.567
R1049 B.n36 B.t3 386.567
R1050 B.n111 B.t1 360.505
R1051 B.n43 B.t8 360.505
R1052 B.n244 B.t10 360.505
R1053 B.n36 B.t5 360.505
R1054 B.n112 B.t2 329.863
R1055 B.n44 B.t7 329.863
R1056 B.n245 B.t11 329.863
R1057 B.n37 B.t4 329.863
R1058 B.n577 B.n576 256.663
R1059 B.n576 B.n575 235.042
R1060 B.n576 B.n2 235.042
R1061 B.n197 B.n134 163.367
R1062 B.n198 B.n197 163.367
R1063 B.n199 B.n198 163.367
R1064 B.n199 B.n132 163.367
R1065 B.n203 B.n132 163.367
R1066 B.n204 B.n203 163.367
R1067 B.n205 B.n204 163.367
R1068 B.n205 B.n130 163.367
R1069 B.n209 B.n130 163.367
R1070 B.n210 B.n209 163.367
R1071 B.n211 B.n210 163.367
R1072 B.n211 B.n128 163.367
R1073 B.n215 B.n128 163.367
R1074 B.n216 B.n215 163.367
R1075 B.n217 B.n216 163.367
R1076 B.n217 B.n126 163.367
R1077 B.n221 B.n126 163.367
R1078 B.n222 B.n221 163.367
R1079 B.n223 B.n222 163.367
R1080 B.n223 B.n124 163.367
R1081 B.n227 B.n124 163.367
R1082 B.n228 B.n227 163.367
R1083 B.n229 B.n228 163.367
R1084 B.n229 B.n122 163.367
R1085 B.n233 B.n122 163.367
R1086 B.n234 B.n233 163.367
R1087 B.n235 B.n234 163.367
R1088 B.n235 B.n120 163.367
R1089 B.n239 B.n120 163.367
R1090 B.n240 B.n239 163.367
R1091 B.n241 B.n240 163.367
R1092 B.n241 B.n118 163.367
R1093 B.n248 B.n118 163.367
R1094 B.n249 B.n248 163.367
R1095 B.n250 B.n249 163.367
R1096 B.n250 B.n116 163.367
R1097 B.n254 B.n116 163.367
R1098 B.n255 B.n254 163.367
R1099 B.n256 B.n255 163.367
R1100 B.n256 B.n114 163.367
R1101 B.n260 B.n114 163.367
R1102 B.n261 B.n260 163.367
R1103 B.n262 B.n261 163.367
R1104 B.n262 B.n110 163.367
R1105 B.n267 B.n110 163.367
R1106 B.n268 B.n267 163.367
R1107 B.n269 B.n268 163.367
R1108 B.n269 B.n108 163.367
R1109 B.n273 B.n108 163.367
R1110 B.n274 B.n273 163.367
R1111 B.n275 B.n274 163.367
R1112 B.n275 B.n106 163.367
R1113 B.n279 B.n106 163.367
R1114 B.n280 B.n279 163.367
R1115 B.n281 B.n280 163.367
R1116 B.n281 B.n104 163.367
R1117 B.n285 B.n104 163.367
R1118 B.n286 B.n285 163.367
R1119 B.n287 B.n286 163.367
R1120 B.n287 B.n102 163.367
R1121 B.n291 B.n102 163.367
R1122 B.n292 B.n291 163.367
R1123 B.n293 B.n292 163.367
R1124 B.n293 B.n100 163.367
R1125 B.n297 B.n100 163.367
R1126 B.n298 B.n297 163.367
R1127 B.n299 B.n298 163.367
R1128 B.n299 B.n98 163.367
R1129 B.n303 B.n98 163.367
R1130 B.n304 B.n303 163.367
R1131 B.n305 B.n304 163.367
R1132 B.n305 B.n96 163.367
R1133 B.n309 B.n96 163.367
R1134 B.n310 B.n309 163.367
R1135 B.n311 B.n310 163.367
R1136 B.n311 B.n94 163.367
R1137 B.n315 B.n94 163.367
R1138 B.n411 B.n62 163.367
R1139 B.n407 B.n62 163.367
R1140 B.n407 B.n406 163.367
R1141 B.n406 B.n405 163.367
R1142 B.n405 B.n64 163.367
R1143 B.n401 B.n64 163.367
R1144 B.n401 B.n400 163.367
R1145 B.n400 B.n399 163.367
R1146 B.n399 B.n66 163.367
R1147 B.n395 B.n66 163.367
R1148 B.n395 B.n394 163.367
R1149 B.n394 B.n393 163.367
R1150 B.n393 B.n68 163.367
R1151 B.n389 B.n68 163.367
R1152 B.n389 B.n388 163.367
R1153 B.n388 B.n387 163.367
R1154 B.n387 B.n70 163.367
R1155 B.n383 B.n70 163.367
R1156 B.n383 B.n382 163.367
R1157 B.n382 B.n381 163.367
R1158 B.n381 B.n72 163.367
R1159 B.n377 B.n72 163.367
R1160 B.n377 B.n376 163.367
R1161 B.n376 B.n375 163.367
R1162 B.n375 B.n74 163.367
R1163 B.n371 B.n74 163.367
R1164 B.n371 B.n370 163.367
R1165 B.n370 B.n369 163.367
R1166 B.n369 B.n76 163.367
R1167 B.n365 B.n76 163.367
R1168 B.n365 B.n364 163.367
R1169 B.n364 B.n363 163.367
R1170 B.n363 B.n78 163.367
R1171 B.n359 B.n78 163.367
R1172 B.n359 B.n358 163.367
R1173 B.n358 B.n357 163.367
R1174 B.n357 B.n80 163.367
R1175 B.n353 B.n80 163.367
R1176 B.n353 B.n352 163.367
R1177 B.n352 B.n351 163.367
R1178 B.n351 B.n82 163.367
R1179 B.n347 B.n82 163.367
R1180 B.n347 B.n346 163.367
R1181 B.n346 B.n345 163.367
R1182 B.n345 B.n84 163.367
R1183 B.n341 B.n84 163.367
R1184 B.n341 B.n340 163.367
R1185 B.n340 B.n339 163.367
R1186 B.n339 B.n86 163.367
R1187 B.n335 B.n86 163.367
R1188 B.n335 B.n334 163.367
R1189 B.n334 B.n333 163.367
R1190 B.n333 B.n88 163.367
R1191 B.n329 B.n88 163.367
R1192 B.n329 B.n328 163.367
R1193 B.n328 B.n327 163.367
R1194 B.n327 B.n90 163.367
R1195 B.n323 B.n90 163.367
R1196 B.n323 B.n322 163.367
R1197 B.n322 B.n321 163.367
R1198 B.n321 B.n92 163.367
R1199 B.n317 B.n92 163.367
R1200 B.n317 B.n316 163.367
R1201 B.n528 B.n527 163.367
R1202 B.n527 B.n526 163.367
R1203 B.n526 B.n19 163.367
R1204 B.n522 B.n19 163.367
R1205 B.n522 B.n521 163.367
R1206 B.n521 B.n520 163.367
R1207 B.n520 B.n21 163.367
R1208 B.n516 B.n21 163.367
R1209 B.n516 B.n515 163.367
R1210 B.n515 B.n514 163.367
R1211 B.n514 B.n23 163.367
R1212 B.n510 B.n23 163.367
R1213 B.n510 B.n509 163.367
R1214 B.n509 B.n508 163.367
R1215 B.n508 B.n25 163.367
R1216 B.n504 B.n25 163.367
R1217 B.n504 B.n503 163.367
R1218 B.n503 B.n502 163.367
R1219 B.n502 B.n27 163.367
R1220 B.n498 B.n27 163.367
R1221 B.n498 B.n497 163.367
R1222 B.n497 B.n496 163.367
R1223 B.n496 B.n29 163.367
R1224 B.n492 B.n29 163.367
R1225 B.n492 B.n491 163.367
R1226 B.n491 B.n490 163.367
R1227 B.n490 B.n31 163.367
R1228 B.n486 B.n31 163.367
R1229 B.n486 B.n485 163.367
R1230 B.n485 B.n484 163.367
R1231 B.n484 B.n33 163.367
R1232 B.n480 B.n33 163.367
R1233 B.n480 B.n479 163.367
R1234 B.n479 B.n478 163.367
R1235 B.n478 B.n35 163.367
R1236 B.n474 B.n35 163.367
R1237 B.n474 B.n473 163.367
R1238 B.n473 B.n472 163.367
R1239 B.n472 B.n40 163.367
R1240 B.n468 B.n40 163.367
R1241 B.n468 B.n467 163.367
R1242 B.n467 B.n466 163.367
R1243 B.n466 B.n42 163.367
R1244 B.n461 B.n42 163.367
R1245 B.n461 B.n460 163.367
R1246 B.n460 B.n459 163.367
R1247 B.n459 B.n46 163.367
R1248 B.n455 B.n46 163.367
R1249 B.n455 B.n454 163.367
R1250 B.n454 B.n453 163.367
R1251 B.n453 B.n48 163.367
R1252 B.n449 B.n48 163.367
R1253 B.n449 B.n448 163.367
R1254 B.n448 B.n447 163.367
R1255 B.n447 B.n50 163.367
R1256 B.n443 B.n50 163.367
R1257 B.n443 B.n442 163.367
R1258 B.n442 B.n441 163.367
R1259 B.n441 B.n52 163.367
R1260 B.n437 B.n52 163.367
R1261 B.n437 B.n436 163.367
R1262 B.n436 B.n435 163.367
R1263 B.n435 B.n54 163.367
R1264 B.n431 B.n54 163.367
R1265 B.n431 B.n430 163.367
R1266 B.n430 B.n429 163.367
R1267 B.n429 B.n56 163.367
R1268 B.n425 B.n56 163.367
R1269 B.n425 B.n424 163.367
R1270 B.n424 B.n423 163.367
R1271 B.n423 B.n58 163.367
R1272 B.n419 B.n58 163.367
R1273 B.n419 B.n418 163.367
R1274 B.n418 B.n417 163.367
R1275 B.n417 B.n60 163.367
R1276 B.n413 B.n60 163.367
R1277 B.n413 B.n412 163.367
R1278 B.n532 B.n17 163.367
R1279 B.n533 B.n532 163.367
R1280 B.n534 B.n533 163.367
R1281 B.n534 B.n15 163.367
R1282 B.n538 B.n15 163.367
R1283 B.n539 B.n538 163.367
R1284 B.n540 B.n539 163.367
R1285 B.n540 B.n13 163.367
R1286 B.n544 B.n13 163.367
R1287 B.n545 B.n544 163.367
R1288 B.n546 B.n545 163.367
R1289 B.n546 B.n11 163.367
R1290 B.n550 B.n11 163.367
R1291 B.n551 B.n550 163.367
R1292 B.n552 B.n551 163.367
R1293 B.n552 B.n9 163.367
R1294 B.n556 B.n9 163.367
R1295 B.n557 B.n556 163.367
R1296 B.n558 B.n557 163.367
R1297 B.n558 B.n7 163.367
R1298 B.n562 B.n7 163.367
R1299 B.n563 B.n562 163.367
R1300 B.n564 B.n563 163.367
R1301 B.n564 B.n5 163.367
R1302 B.n568 B.n5 163.367
R1303 B.n569 B.n568 163.367
R1304 B.n570 B.n569 163.367
R1305 B.n570 B.n3 163.367
R1306 B.n574 B.n3 163.367
R1307 B.n575 B.n574 163.367
R1308 B.n150 B.n2 163.367
R1309 B.n151 B.n150 163.367
R1310 B.n151 B.n148 163.367
R1311 B.n155 B.n148 163.367
R1312 B.n156 B.n155 163.367
R1313 B.n157 B.n156 163.367
R1314 B.n157 B.n146 163.367
R1315 B.n161 B.n146 163.367
R1316 B.n162 B.n161 163.367
R1317 B.n163 B.n162 163.367
R1318 B.n163 B.n144 163.367
R1319 B.n167 B.n144 163.367
R1320 B.n168 B.n167 163.367
R1321 B.n169 B.n168 163.367
R1322 B.n169 B.n142 163.367
R1323 B.n173 B.n142 163.367
R1324 B.n174 B.n173 163.367
R1325 B.n175 B.n174 163.367
R1326 B.n175 B.n140 163.367
R1327 B.n179 B.n140 163.367
R1328 B.n180 B.n179 163.367
R1329 B.n181 B.n180 163.367
R1330 B.n181 B.n138 163.367
R1331 B.n185 B.n138 163.367
R1332 B.n186 B.n185 163.367
R1333 B.n187 B.n186 163.367
R1334 B.n187 B.n136 163.367
R1335 B.n191 B.n136 163.367
R1336 B.n192 B.n191 163.367
R1337 B.n193 B.n192 163.367
R1338 B.n246 B.n245 59.5399
R1339 B.n264 B.n112 59.5399
R1340 B.n463 B.n44 59.5399
R1341 B.n38 B.n37 59.5399
R1342 B.n245 B.n244 30.6429
R1343 B.n112 B.n111 30.6429
R1344 B.n44 B.n43 30.6429
R1345 B.n37 B.n36 30.6429
R1346 B.n530 B.n529 29.8151
R1347 B.n410 B.n61 29.8151
R1348 B.n314 B.n93 29.8151
R1349 B.n195 B.n194 29.8151
R1350 B B.n577 18.0485
R1351 B.n531 B.n530 10.6151
R1352 B.n531 B.n16 10.6151
R1353 B.n535 B.n16 10.6151
R1354 B.n536 B.n535 10.6151
R1355 B.n537 B.n536 10.6151
R1356 B.n537 B.n14 10.6151
R1357 B.n541 B.n14 10.6151
R1358 B.n542 B.n541 10.6151
R1359 B.n543 B.n542 10.6151
R1360 B.n543 B.n12 10.6151
R1361 B.n547 B.n12 10.6151
R1362 B.n548 B.n547 10.6151
R1363 B.n549 B.n548 10.6151
R1364 B.n549 B.n10 10.6151
R1365 B.n553 B.n10 10.6151
R1366 B.n554 B.n553 10.6151
R1367 B.n555 B.n554 10.6151
R1368 B.n555 B.n8 10.6151
R1369 B.n559 B.n8 10.6151
R1370 B.n560 B.n559 10.6151
R1371 B.n561 B.n560 10.6151
R1372 B.n561 B.n6 10.6151
R1373 B.n565 B.n6 10.6151
R1374 B.n566 B.n565 10.6151
R1375 B.n567 B.n566 10.6151
R1376 B.n567 B.n4 10.6151
R1377 B.n571 B.n4 10.6151
R1378 B.n572 B.n571 10.6151
R1379 B.n573 B.n572 10.6151
R1380 B.n573 B.n0 10.6151
R1381 B.n529 B.n18 10.6151
R1382 B.n525 B.n18 10.6151
R1383 B.n525 B.n524 10.6151
R1384 B.n524 B.n523 10.6151
R1385 B.n523 B.n20 10.6151
R1386 B.n519 B.n20 10.6151
R1387 B.n519 B.n518 10.6151
R1388 B.n518 B.n517 10.6151
R1389 B.n517 B.n22 10.6151
R1390 B.n513 B.n22 10.6151
R1391 B.n513 B.n512 10.6151
R1392 B.n512 B.n511 10.6151
R1393 B.n511 B.n24 10.6151
R1394 B.n507 B.n24 10.6151
R1395 B.n507 B.n506 10.6151
R1396 B.n506 B.n505 10.6151
R1397 B.n505 B.n26 10.6151
R1398 B.n501 B.n26 10.6151
R1399 B.n501 B.n500 10.6151
R1400 B.n500 B.n499 10.6151
R1401 B.n499 B.n28 10.6151
R1402 B.n495 B.n28 10.6151
R1403 B.n495 B.n494 10.6151
R1404 B.n494 B.n493 10.6151
R1405 B.n493 B.n30 10.6151
R1406 B.n489 B.n30 10.6151
R1407 B.n489 B.n488 10.6151
R1408 B.n488 B.n487 10.6151
R1409 B.n487 B.n32 10.6151
R1410 B.n483 B.n32 10.6151
R1411 B.n483 B.n482 10.6151
R1412 B.n482 B.n481 10.6151
R1413 B.n481 B.n34 10.6151
R1414 B.n477 B.n476 10.6151
R1415 B.n476 B.n475 10.6151
R1416 B.n475 B.n39 10.6151
R1417 B.n471 B.n39 10.6151
R1418 B.n471 B.n470 10.6151
R1419 B.n470 B.n469 10.6151
R1420 B.n469 B.n41 10.6151
R1421 B.n465 B.n41 10.6151
R1422 B.n465 B.n464 10.6151
R1423 B.n462 B.n45 10.6151
R1424 B.n458 B.n45 10.6151
R1425 B.n458 B.n457 10.6151
R1426 B.n457 B.n456 10.6151
R1427 B.n456 B.n47 10.6151
R1428 B.n452 B.n47 10.6151
R1429 B.n452 B.n451 10.6151
R1430 B.n451 B.n450 10.6151
R1431 B.n450 B.n49 10.6151
R1432 B.n446 B.n49 10.6151
R1433 B.n446 B.n445 10.6151
R1434 B.n445 B.n444 10.6151
R1435 B.n444 B.n51 10.6151
R1436 B.n440 B.n51 10.6151
R1437 B.n440 B.n439 10.6151
R1438 B.n439 B.n438 10.6151
R1439 B.n438 B.n53 10.6151
R1440 B.n434 B.n53 10.6151
R1441 B.n434 B.n433 10.6151
R1442 B.n433 B.n432 10.6151
R1443 B.n432 B.n55 10.6151
R1444 B.n428 B.n55 10.6151
R1445 B.n428 B.n427 10.6151
R1446 B.n427 B.n426 10.6151
R1447 B.n426 B.n57 10.6151
R1448 B.n422 B.n57 10.6151
R1449 B.n422 B.n421 10.6151
R1450 B.n421 B.n420 10.6151
R1451 B.n420 B.n59 10.6151
R1452 B.n416 B.n59 10.6151
R1453 B.n416 B.n415 10.6151
R1454 B.n415 B.n414 10.6151
R1455 B.n414 B.n61 10.6151
R1456 B.n410 B.n409 10.6151
R1457 B.n409 B.n408 10.6151
R1458 B.n408 B.n63 10.6151
R1459 B.n404 B.n63 10.6151
R1460 B.n404 B.n403 10.6151
R1461 B.n403 B.n402 10.6151
R1462 B.n402 B.n65 10.6151
R1463 B.n398 B.n65 10.6151
R1464 B.n398 B.n397 10.6151
R1465 B.n397 B.n396 10.6151
R1466 B.n396 B.n67 10.6151
R1467 B.n392 B.n67 10.6151
R1468 B.n392 B.n391 10.6151
R1469 B.n391 B.n390 10.6151
R1470 B.n390 B.n69 10.6151
R1471 B.n386 B.n69 10.6151
R1472 B.n386 B.n385 10.6151
R1473 B.n385 B.n384 10.6151
R1474 B.n384 B.n71 10.6151
R1475 B.n380 B.n71 10.6151
R1476 B.n380 B.n379 10.6151
R1477 B.n379 B.n378 10.6151
R1478 B.n378 B.n73 10.6151
R1479 B.n374 B.n73 10.6151
R1480 B.n374 B.n373 10.6151
R1481 B.n373 B.n372 10.6151
R1482 B.n372 B.n75 10.6151
R1483 B.n368 B.n75 10.6151
R1484 B.n368 B.n367 10.6151
R1485 B.n367 B.n366 10.6151
R1486 B.n366 B.n77 10.6151
R1487 B.n362 B.n77 10.6151
R1488 B.n362 B.n361 10.6151
R1489 B.n361 B.n360 10.6151
R1490 B.n360 B.n79 10.6151
R1491 B.n356 B.n79 10.6151
R1492 B.n356 B.n355 10.6151
R1493 B.n355 B.n354 10.6151
R1494 B.n354 B.n81 10.6151
R1495 B.n350 B.n81 10.6151
R1496 B.n350 B.n349 10.6151
R1497 B.n349 B.n348 10.6151
R1498 B.n348 B.n83 10.6151
R1499 B.n344 B.n83 10.6151
R1500 B.n344 B.n343 10.6151
R1501 B.n343 B.n342 10.6151
R1502 B.n342 B.n85 10.6151
R1503 B.n338 B.n85 10.6151
R1504 B.n338 B.n337 10.6151
R1505 B.n337 B.n336 10.6151
R1506 B.n336 B.n87 10.6151
R1507 B.n332 B.n87 10.6151
R1508 B.n332 B.n331 10.6151
R1509 B.n331 B.n330 10.6151
R1510 B.n330 B.n89 10.6151
R1511 B.n326 B.n89 10.6151
R1512 B.n326 B.n325 10.6151
R1513 B.n325 B.n324 10.6151
R1514 B.n324 B.n91 10.6151
R1515 B.n320 B.n91 10.6151
R1516 B.n320 B.n319 10.6151
R1517 B.n319 B.n318 10.6151
R1518 B.n318 B.n93 10.6151
R1519 B.n149 B.n1 10.6151
R1520 B.n152 B.n149 10.6151
R1521 B.n153 B.n152 10.6151
R1522 B.n154 B.n153 10.6151
R1523 B.n154 B.n147 10.6151
R1524 B.n158 B.n147 10.6151
R1525 B.n159 B.n158 10.6151
R1526 B.n160 B.n159 10.6151
R1527 B.n160 B.n145 10.6151
R1528 B.n164 B.n145 10.6151
R1529 B.n165 B.n164 10.6151
R1530 B.n166 B.n165 10.6151
R1531 B.n166 B.n143 10.6151
R1532 B.n170 B.n143 10.6151
R1533 B.n171 B.n170 10.6151
R1534 B.n172 B.n171 10.6151
R1535 B.n172 B.n141 10.6151
R1536 B.n176 B.n141 10.6151
R1537 B.n177 B.n176 10.6151
R1538 B.n178 B.n177 10.6151
R1539 B.n178 B.n139 10.6151
R1540 B.n182 B.n139 10.6151
R1541 B.n183 B.n182 10.6151
R1542 B.n184 B.n183 10.6151
R1543 B.n184 B.n137 10.6151
R1544 B.n188 B.n137 10.6151
R1545 B.n189 B.n188 10.6151
R1546 B.n190 B.n189 10.6151
R1547 B.n190 B.n135 10.6151
R1548 B.n194 B.n135 10.6151
R1549 B.n196 B.n195 10.6151
R1550 B.n196 B.n133 10.6151
R1551 B.n200 B.n133 10.6151
R1552 B.n201 B.n200 10.6151
R1553 B.n202 B.n201 10.6151
R1554 B.n202 B.n131 10.6151
R1555 B.n206 B.n131 10.6151
R1556 B.n207 B.n206 10.6151
R1557 B.n208 B.n207 10.6151
R1558 B.n208 B.n129 10.6151
R1559 B.n212 B.n129 10.6151
R1560 B.n213 B.n212 10.6151
R1561 B.n214 B.n213 10.6151
R1562 B.n214 B.n127 10.6151
R1563 B.n218 B.n127 10.6151
R1564 B.n219 B.n218 10.6151
R1565 B.n220 B.n219 10.6151
R1566 B.n220 B.n125 10.6151
R1567 B.n224 B.n125 10.6151
R1568 B.n225 B.n224 10.6151
R1569 B.n226 B.n225 10.6151
R1570 B.n226 B.n123 10.6151
R1571 B.n230 B.n123 10.6151
R1572 B.n231 B.n230 10.6151
R1573 B.n232 B.n231 10.6151
R1574 B.n232 B.n121 10.6151
R1575 B.n236 B.n121 10.6151
R1576 B.n237 B.n236 10.6151
R1577 B.n238 B.n237 10.6151
R1578 B.n238 B.n119 10.6151
R1579 B.n242 B.n119 10.6151
R1580 B.n243 B.n242 10.6151
R1581 B.n247 B.n243 10.6151
R1582 B.n251 B.n117 10.6151
R1583 B.n252 B.n251 10.6151
R1584 B.n253 B.n252 10.6151
R1585 B.n253 B.n115 10.6151
R1586 B.n257 B.n115 10.6151
R1587 B.n258 B.n257 10.6151
R1588 B.n259 B.n258 10.6151
R1589 B.n259 B.n113 10.6151
R1590 B.n263 B.n113 10.6151
R1591 B.n266 B.n265 10.6151
R1592 B.n266 B.n109 10.6151
R1593 B.n270 B.n109 10.6151
R1594 B.n271 B.n270 10.6151
R1595 B.n272 B.n271 10.6151
R1596 B.n272 B.n107 10.6151
R1597 B.n276 B.n107 10.6151
R1598 B.n277 B.n276 10.6151
R1599 B.n278 B.n277 10.6151
R1600 B.n278 B.n105 10.6151
R1601 B.n282 B.n105 10.6151
R1602 B.n283 B.n282 10.6151
R1603 B.n284 B.n283 10.6151
R1604 B.n284 B.n103 10.6151
R1605 B.n288 B.n103 10.6151
R1606 B.n289 B.n288 10.6151
R1607 B.n290 B.n289 10.6151
R1608 B.n290 B.n101 10.6151
R1609 B.n294 B.n101 10.6151
R1610 B.n295 B.n294 10.6151
R1611 B.n296 B.n295 10.6151
R1612 B.n296 B.n99 10.6151
R1613 B.n300 B.n99 10.6151
R1614 B.n301 B.n300 10.6151
R1615 B.n302 B.n301 10.6151
R1616 B.n302 B.n97 10.6151
R1617 B.n306 B.n97 10.6151
R1618 B.n307 B.n306 10.6151
R1619 B.n308 B.n307 10.6151
R1620 B.n308 B.n95 10.6151
R1621 B.n312 B.n95 10.6151
R1622 B.n313 B.n312 10.6151
R1623 B.n314 B.n313 10.6151
R1624 B.n38 B.n34 9.36635
R1625 B.n463 B.n462 9.36635
R1626 B.n247 B.n246 9.36635
R1627 B.n265 B.n264 9.36635
R1628 B.n577 B.n0 8.11757
R1629 B.n577 B.n1 8.11757
R1630 B.n477 B.n38 1.24928
R1631 B.n464 B.n463 1.24928
R1632 B.n246 B.n117 1.24928
R1633 B.n264 B.n263 1.24928
C0 VN VDD1 0.149029f
C1 VN VDD2 5.68833f
C2 VTAIL VDD1 7.56118f
C3 VN w_n2550_n2858# 4.76453f
C4 VDD2 VTAIL 7.60655f
C5 VN VP 5.53752f
C6 w_n2550_n2858# VTAIL 3.53977f
C7 VN B 0.880654f
C8 VTAIL VP 5.76417f
C9 VDD2 VDD1 1.10013f
C10 VTAIL B 3.49786f
C11 w_n2550_n2858# VDD1 1.43191f
C12 VDD1 VP 5.91435f
C13 w_n2550_n2858# VDD2 1.48987f
C14 VDD2 VP 0.375759f
C15 VDD1 B 1.16943f
C16 w_n2550_n2858# VP 5.09159f
C17 VDD2 B 1.22313f
C18 VN VTAIL 5.75006f
C19 w_n2550_n2858# B 7.3336f
C20 VP B 1.42173f
C21 VDD2 VSUBS 1.338985f
C22 VDD1 VSUBS 1.745991f
C23 VTAIL VSUBS 0.948785f
C24 VN VSUBS 5.02405f
C25 VP VSUBS 2.126996f
C26 B VSUBS 3.282469f
C27 w_n2550_n2858# VSUBS 90.117004f
C28 B.n0 VSUBS 0.00702f
C29 B.n1 VSUBS 0.00702f
C30 B.n2 VSUBS 0.010382f
C31 B.n3 VSUBS 0.007956f
C32 B.n4 VSUBS 0.007956f
C33 B.n5 VSUBS 0.007956f
C34 B.n6 VSUBS 0.007956f
C35 B.n7 VSUBS 0.007956f
C36 B.n8 VSUBS 0.007956f
C37 B.n9 VSUBS 0.007956f
C38 B.n10 VSUBS 0.007956f
C39 B.n11 VSUBS 0.007956f
C40 B.n12 VSUBS 0.007956f
C41 B.n13 VSUBS 0.007956f
C42 B.n14 VSUBS 0.007956f
C43 B.n15 VSUBS 0.007956f
C44 B.n16 VSUBS 0.007956f
C45 B.n17 VSUBS 0.017111f
C46 B.n18 VSUBS 0.007956f
C47 B.n19 VSUBS 0.007956f
C48 B.n20 VSUBS 0.007956f
C49 B.n21 VSUBS 0.007956f
C50 B.n22 VSUBS 0.007956f
C51 B.n23 VSUBS 0.007956f
C52 B.n24 VSUBS 0.007956f
C53 B.n25 VSUBS 0.007956f
C54 B.n26 VSUBS 0.007956f
C55 B.n27 VSUBS 0.007956f
C56 B.n28 VSUBS 0.007956f
C57 B.n29 VSUBS 0.007956f
C58 B.n30 VSUBS 0.007956f
C59 B.n31 VSUBS 0.007956f
C60 B.n32 VSUBS 0.007956f
C61 B.n33 VSUBS 0.007956f
C62 B.n34 VSUBS 0.007488f
C63 B.n35 VSUBS 0.007956f
C64 B.t4 VSUBS 0.177496f
C65 B.t5 VSUBS 0.196714f
C66 B.t3 VSUBS 0.588656f
C67 B.n36 VSUBS 0.31351f
C68 B.n37 VSUBS 0.237444f
C69 B.n38 VSUBS 0.018434f
C70 B.n39 VSUBS 0.007956f
C71 B.n40 VSUBS 0.007956f
C72 B.n41 VSUBS 0.007956f
C73 B.n42 VSUBS 0.007956f
C74 B.t7 VSUBS 0.177499f
C75 B.t8 VSUBS 0.196717f
C76 B.t6 VSUBS 0.588656f
C77 B.n43 VSUBS 0.313508f
C78 B.n44 VSUBS 0.237441f
C79 B.n45 VSUBS 0.007956f
C80 B.n46 VSUBS 0.007956f
C81 B.n47 VSUBS 0.007956f
C82 B.n48 VSUBS 0.007956f
C83 B.n49 VSUBS 0.007956f
C84 B.n50 VSUBS 0.007956f
C85 B.n51 VSUBS 0.007956f
C86 B.n52 VSUBS 0.007956f
C87 B.n53 VSUBS 0.007956f
C88 B.n54 VSUBS 0.007956f
C89 B.n55 VSUBS 0.007956f
C90 B.n56 VSUBS 0.007956f
C91 B.n57 VSUBS 0.007956f
C92 B.n58 VSUBS 0.007956f
C93 B.n59 VSUBS 0.007956f
C94 B.n60 VSUBS 0.007956f
C95 B.n61 VSUBS 0.01799f
C96 B.n62 VSUBS 0.007956f
C97 B.n63 VSUBS 0.007956f
C98 B.n64 VSUBS 0.007956f
C99 B.n65 VSUBS 0.007956f
C100 B.n66 VSUBS 0.007956f
C101 B.n67 VSUBS 0.007956f
C102 B.n68 VSUBS 0.007956f
C103 B.n69 VSUBS 0.007956f
C104 B.n70 VSUBS 0.007956f
C105 B.n71 VSUBS 0.007956f
C106 B.n72 VSUBS 0.007956f
C107 B.n73 VSUBS 0.007956f
C108 B.n74 VSUBS 0.007956f
C109 B.n75 VSUBS 0.007956f
C110 B.n76 VSUBS 0.007956f
C111 B.n77 VSUBS 0.007956f
C112 B.n78 VSUBS 0.007956f
C113 B.n79 VSUBS 0.007956f
C114 B.n80 VSUBS 0.007956f
C115 B.n81 VSUBS 0.007956f
C116 B.n82 VSUBS 0.007956f
C117 B.n83 VSUBS 0.007956f
C118 B.n84 VSUBS 0.007956f
C119 B.n85 VSUBS 0.007956f
C120 B.n86 VSUBS 0.007956f
C121 B.n87 VSUBS 0.007956f
C122 B.n88 VSUBS 0.007956f
C123 B.n89 VSUBS 0.007956f
C124 B.n90 VSUBS 0.007956f
C125 B.n91 VSUBS 0.007956f
C126 B.n92 VSUBS 0.007956f
C127 B.n93 VSUBS 0.018141f
C128 B.n94 VSUBS 0.007956f
C129 B.n95 VSUBS 0.007956f
C130 B.n96 VSUBS 0.007956f
C131 B.n97 VSUBS 0.007956f
C132 B.n98 VSUBS 0.007956f
C133 B.n99 VSUBS 0.007956f
C134 B.n100 VSUBS 0.007956f
C135 B.n101 VSUBS 0.007956f
C136 B.n102 VSUBS 0.007956f
C137 B.n103 VSUBS 0.007956f
C138 B.n104 VSUBS 0.007956f
C139 B.n105 VSUBS 0.007956f
C140 B.n106 VSUBS 0.007956f
C141 B.n107 VSUBS 0.007956f
C142 B.n108 VSUBS 0.007956f
C143 B.n109 VSUBS 0.007956f
C144 B.n110 VSUBS 0.007956f
C145 B.t2 VSUBS 0.177499f
C146 B.t1 VSUBS 0.196717f
C147 B.t0 VSUBS 0.588656f
C148 B.n111 VSUBS 0.313508f
C149 B.n112 VSUBS 0.237441f
C150 B.n113 VSUBS 0.007956f
C151 B.n114 VSUBS 0.007956f
C152 B.n115 VSUBS 0.007956f
C153 B.n116 VSUBS 0.007956f
C154 B.n117 VSUBS 0.004446f
C155 B.n118 VSUBS 0.007956f
C156 B.n119 VSUBS 0.007956f
C157 B.n120 VSUBS 0.007956f
C158 B.n121 VSUBS 0.007956f
C159 B.n122 VSUBS 0.007956f
C160 B.n123 VSUBS 0.007956f
C161 B.n124 VSUBS 0.007956f
C162 B.n125 VSUBS 0.007956f
C163 B.n126 VSUBS 0.007956f
C164 B.n127 VSUBS 0.007956f
C165 B.n128 VSUBS 0.007956f
C166 B.n129 VSUBS 0.007956f
C167 B.n130 VSUBS 0.007956f
C168 B.n131 VSUBS 0.007956f
C169 B.n132 VSUBS 0.007956f
C170 B.n133 VSUBS 0.007956f
C171 B.n134 VSUBS 0.01799f
C172 B.n135 VSUBS 0.007956f
C173 B.n136 VSUBS 0.007956f
C174 B.n137 VSUBS 0.007956f
C175 B.n138 VSUBS 0.007956f
C176 B.n139 VSUBS 0.007956f
C177 B.n140 VSUBS 0.007956f
C178 B.n141 VSUBS 0.007956f
C179 B.n142 VSUBS 0.007956f
C180 B.n143 VSUBS 0.007956f
C181 B.n144 VSUBS 0.007956f
C182 B.n145 VSUBS 0.007956f
C183 B.n146 VSUBS 0.007956f
C184 B.n147 VSUBS 0.007956f
C185 B.n148 VSUBS 0.007956f
C186 B.n149 VSUBS 0.007956f
C187 B.n150 VSUBS 0.007956f
C188 B.n151 VSUBS 0.007956f
C189 B.n152 VSUBS 0.007956f
C190 B.n153 VSUBS 0.007956f
C191 B.n154 VSUBS 0.007956f
C192 B.n155 VSUBS 0.007956f
C193 B.n156 VSUBS 0.007956f
C194 B.n157 VSUBS 0.007956f
C195 B.n158 VSUBS 0.007956f
C196 B.n159 VSUBS 0.007956f
C197 B.n160 VSUBS 0.007956f
C198 B.n161 VSUBS 0.007956f
C199 B.n162 VSUBS 0.007956f
C200 B.n163 VSUBS 0.007956f
C201 B.n164 VSUBS 0.007956f
C202 B.n165 VSUBS 0.007956f
C203 B.n166 VSUBS 0.007956f
C204 B.n167 VSUBS 0.007956f
C205 B.n168 VSUBS 0.007956f
C206 B.n169 VSUBS 0.007956f
C207 B.n170 VSUBS 0.007956f
C208 B.n171 VSUBS 0.007956f
C209 B.n172 VSUBS 0.007956f
C210 B.n173 VSUBS 0.007956f
C211 B.n174 VSUBS 0.007956f
C212 B.n175 VSUBS 0.007956f
C213 B.n176 VSUBS 0.007956f
C214 B.n177 VSUBS 0.007956f
C215 B.n178 VSUBS 0.007956f
C216 B.n179 VSUBS 0.007956f
C217 B.n180 VSUBS 0.007956f
C218 B.n181 VSUBS 0.007956f
C219 B.n182 VSUBS 0.007956f
C220 B.n183 VSUBS 0.007956f
C221 B.n184 VSUBS 0.007956f
C222 B.n185 VSUBS 0.007956f
C223 B.n186 VSUBS 0.007956f
C224 B.n187 VSUBS 0.007956f
C225 B.n188 VSUBS 0.007956f
C226 B.n189 VSUBS 0.007956f
C227 B.n190 VSUBS 0.007956f
C228 B.n191 VSUBS 0.007956f
C229 B.n192 VSUBS 0.007956f
C230 B.n193 VSUBS 0.017111f
C231 B.n194 VSUBS 0.017111f
C232 B.n195 VSUBS 0.01799f
C233 B.n196 VSUBS 0.007956f
C234 B.n197 VSUBS 0.007956f
C235 B.n198 VSUBS 0.007956f
C236 B.n199 VSUBS 0.007956f
C237 B.n200 VSUBS 0.007956f
C238 B.n201 VSUBS 0.007956f
C239 B.n202 VSUBS 0.007956f
C240 B.n203 VSUBS 0.007956f
C241 B.n204 VSUBS 0.007956f
C242 B.n205 VSUBS 0.007956f
C243 B.n206 VSUBS 0.007956f
C244 B.n207 VSUBS 0.007956f
C245 B.n208 VSUBS 0.007956f
C246 B.n209 VSUBS 0.007956f
C247 B.n210 VSUBS 0.007956f
C248 B.n211 VSUBS 0.007956f
C249 B.n212 VSUBS 0.007956f
C250 B.n213 VSUBS 0.007956f
C251 B.n214 VSUBS 0.007956f
C252 B.n215 VSUBS 0.007956f
C253 B.n216 VSUBS 0.007956f
C254 B.n217 VSUBS 0.007956f
C255 B.n218 VSUBS 0.007956f
C256 B.n219 VSUBS 0.007956f
C257 B.n220 VSUBS 0.007956f
C258 B.n221 VSUBS 0.007956f
C259 B.n222 VSUBS 0.007956f
C260 B.n223 VSUBS 0.007956f
C261 B.n224 VSUBS 0.007956f
C262 B.n225 VSUBS 0.007956f
C263 B.n226 VSUBS 0.007956f
C264 B.n227 VSUBS 0.007956f
C265 B.n228 VSUBS 0.007956f
C266 B.n229 VSUBS 0.007956f
C267 B.n230 VSUBS 0.007956f
C268 B.n231 VSUBS 0.007956f
C269 B.n232 VSUBS 0.007956f
C270 B.n233 VSUBS 0.007956f
C271 B.n234 VSUBS 0.007956f
C272 B.n235 VSUBS 0.007956f
C273 B.n236 VSUBS 0.007956f
C274 B.n237 VSUBS 0.007956f
C275 B.n238 VSUBS 0.007956f
C276 B.n239 VSUBS 0.007956f
C277 B.n240 VSUBS 0.007956f
C278 B.n241 VSUBS 0.007956f
C279 B.n242 VSUBS 0.007956f
C280 B.n243 VSUBS 0.007956f
C281 B.t11 VSUBS 0.177496f
C282 B.t10 VSUBS 0.196714f
C283 B.t9 VSUBS 0.588656f
C284 B.n244 VSUBS 0.31351f
C285 B.n245 VSUBS 0.237444f
C286 B.n246 VSUBS 0.018434f
C287 B.n247 VSUBS 0.007488f
C288 B.n248 VSUBS 0.007956f
C289 B.n249 VSUBS 0.007956f
C290 B.n250 VSUBS 0.007956f
C291 B.n251 VSUBS 0.007956f
C292 B.n252 VSUBS 0.007956f
C293 B.n253 VSUBS 0.007956f
C294 B.n254 VSUBS 0.007956f
C295 B.n255 VSUBS 0.007956f
C296 B.n256 VSUBS 0.007956f
C297 B.n257 VSUBS 0.007956f
C298 B.n258 VSUBS 0.007956f
C299 B.n259 VSUBS 0.007956f
C300 B.n260 VSUBS 0.007956f
C301 B.n261 VSUBS 0.007956f
C302 B.n262 VSUBS 0.007956f
C303 B.n263 VSUBS 0.004446f
C304 B.n264 VSUBS 0.018434f
C305 B.n265 VSUBS 0.007488f
C306 B.n266 VSUBS 0.007956f
C307 B.n267 VSUBS 0.007956f
C308 B.n268 VSUBS 0.007956f
C309 B.n269 VSUBS 0.007956f
C310 B.n270 VSUBS 0.007956f
C311 B.n271 VSUBS 0.007956f
C312 B.n272 VSUBS 0.007956f
C313 B.n273 VSUBS 0.007956f
C314 B.n274 VSUBS 0.007956f
C315 B.n275 VSUBS 0.007956f
C316 B.n276 VSUBS 0.007956f
C317 B.n277 VSUBS 0.007956f
C318 B.n278 VSUBS 0.007956f
C319 B.n279 VSUBS 0.007956f
C320 B.n280 VSUBS 0.007956f
C321 B.n281 VSUBS 0.007956f
C322 B.n282 VSUBS 0.007956f
C323 B.n283 VSUBS 0.007956f
C324 B.n284 VSUBS 0.007956f
C325 B.n285 VSUBS 0.007956f
C326 B.n286 VSUBS 0.007956f
C327 B.n287 VSUBS 0.007956f
C328 B.n288 VSUBS 0.007956f
C329 B.n289 VSUBS 0.007956f
C330 B.n290 VSUBS 0.007956f
C331 B.n291 VSUBS 0.007956f
C332 B.n292 VSUBS 0.007956f
C333 B.n293 VSUBS 0.007956f
C334 B.n294 VSUBS 0.007956f
C335 B.n295 VSUBS 0.007956f
C336 B.n296 VSUBS 0.007956f
C337 B.n297 VSUBS 0.007956f
C338 B.n298 VSUBS 0.007956f
C339 B.n299 VSUBS 0.007956f
C340 B.n300 VSUBS 0.007956f
C341 B.n301 VSUBS 0.007956f
C342 B.n302 VSUBS 0.007956f
C343 B.n303 VSUBS 0.007956f
C344 B.n304 VSUBS 0.007956f
C345 B.n305 VSUBS 0.007956f
C346 B.n306 VSUBS 0.007956f
C347 B.n307 VSUBS 0.007956f
C348 B.n308 VSUBS 0.007956f
C349 B.n309 VSUBS 0.007956f
C350 B.n310 VSUBS 0.007956f
C351 B.n311 VSUBS 0.007956f
C352 B.n312 VSUBS 0.007956f
C353 B.n313 VSUBS 0.007956f
C354 B.n314 VSUBS 0.01696f
C355 B.n315 VSUBS 0.01799f
C356 B.n316 VSUBS 0.017111f
C357 B.n317 VSUBS 0.007956f
C358 B.n318 VSUBS 0.007956f
C359 B.n319 VSUBS 0.007956f
C360 B.n320 VSUBS 0.007956f
C361 B.n321 VSUBS 0.007956f
C362 B.n322 VSUBS 0.007956f
C363 B.n323 VSUBS 0.007956f
C364 B.n324 VSUBS 0.007956f
C365 B.n325 VSUBS 0.007956f
C366 B.n326 VSUBS 0.007956f
C367 B.n327 VSUBS 0.007956f
C368 B.n328 VSUBS 0.007956f
C369 B.n329 VSUBS 0.007956f
C370 B.n330 VSUBS 0.007956f
C371 B.n331 VSUBS 0.007956f
C372 B.n332 VSUBS 0.007956f
C373 B.n333 VSUBS 0.007956f
C374 B.n334 VSUBS 0.007956f
C375 B.n335 VSUBS 0.007956f
C376 B.n336 VSUBS 0.007956f
C377 B.n337 VSUBS 0.007956f
C378 B.n338 VSUBS 0.007956f
C379 B.n339 VSUBS 0.007956f
C380 B.n340 VSUBS 0.007956f
C381 B.n341 VSUBS 0.007956f
C382 B.n342 VSUBS 0.007956f
C383 B.n343 VSUBS 0.007956f
C384 B.n344 VSUBS 0.007956f
C385 B.n345 VSUBS 0.007956f
C386 B.n346 VSUBS 0.007956f
C387 B.n347 VSUBS 0.007956f
C388 B.n348 VSUBS 0.007956f
C389 B.n349 VSUBS 0.007956f
C390 B.n350 VSUBS 0.007956f
C391 B.n351 VSUBS 0.007956f
C392 B.n352 VSUBS 0.007956f
C393 B.n353 VSUBS 0.007956f
C394 B.n354 VSUBS 0.007956f
C395 B.n355 VSUBS 0.007956f
C396 B.n356 VSUBS 0.007956f
C397 B.n357 VSUBS 0.007956f
C398 B.n358 VSUBS 0.007956f
C399 B.n359 VSUBS 0.007956f
C400 B.n360 VSUBS 0.007956f
C401 B.n361 VSUBS 0.007956f
C402 B.n362 VSUBS 0.007956f
C403 B.n363 VSUBS 0.007956f
C404 B.n364 VSUBS 0.007956f
C405 B.n365 VSUBS 0.007956f
C406 B.n366 VSUBS 0.007956f
C407 B.n367 VSUBS 0.007956f
C408 B.n368 VSUBS 0.007956f
C409 B.n369 VSUBS 0.007956f
C410 B.n370 VSUBS 0.007956f
C411 B.n371 VSUBS 0.007956f
C412 B.n372 VSUBS 0.007956f
C413 B.n373 VSUBS 0.007956f
C414 B.n374 VSUBS 0.007956f
C415 B.n375 VSUBS 0.007956f
C416 B.n376 VSUBS 0.007956f
C417 B.n377 VSUBS 0.007956f
C418 B.n378 VSUBS 0.007956f
C419 B.n379 VSUBS 0.007956f
C420 B.n380 VSUBS 0.007956f
C421 B.n381 VSUBS 0.007956f
C422 B.n382 VSUBS 0.007956f
C423 B.n383 VSUBS 0.007956f
C424 B.n384 VSUBS 0.007956f
C425 B.n385 VSUBS 0.007956f
C426 B.n386 VSUBS 0.007956f
C427 B.n387 VSUBS 0.007956f
C428 B.n388 VSUBS 0.007956f
C429 B.n389 VSUBS 0.007956f
C430 B.n390 VSUBS 0.007956f
C431 B.n391 VSUBS 0.007956f
C432 B.n392 VSUBS 0.007956f
C433 B.n393 VSUBS 0.007956f
C434 B.n394 VSUBS 0.007956f
C435 B.n395 VSUBS 0.007956f
C436 B.n396 VSUBS 0.007956f
C437 B.n397 VSUBS 0.007956f
C438 B.n398 VSUBS 0.007956f
C439 B.n399 VSUBS 0.007956f
C440 B.n400 VSUBS 0.007956f
C441 B.n401 VSUBS 0.007956f
C442 B.n402 VSUBS 0.007956f
C443 B.n403 VSUBS 0.007956f
C444 B.n404 VSUBS 0.007956f
C445 B.n405 VSUBS 0.007956f
C446 B.n406 VSUBS 0.007956f
C447 B.n407 VSUBS 0.007956f
C448 B.n408 VSUBS 0.007956f
C449 B.n409 VSUBS 0.007956f
C450 B.n410 VSUBS 0.017111f
C451 B.n411 VSUBS 0.017111f
C452 B.n412 VSUBS 0.01799f
C453 B.n413 VSUBS 0.007956f
C454 B.n414 VSUBS 0.007956f
C455 B.n415 VSUBS 0.007956f
C456 B.n416 VSUBS 0.007956f
C457 B.n417 VSUBS 0.007956f
C458 B.n418 VSUBS 0.007956f
C459 B.n419 VSUBS 0.007956f
C460 B.n420 VSUBS 0.007956f
C461 B.n421 VSUBS 0.007956f
C462 B.n422 VSUBS 0.007956f
C463 B.n423 VSUBS 0.007956f
C464 B.n424 VSUBS 0.007956f
C465 B.n425 VSUBS 0.007956f
C466 B.n426 VSUBS 0.007956f
C467 B.n427 VSUBS 0.007956f
C468 B.n428 VSUBS 0.007956f
C469 B.n429 VSUBS 0.007956f
C470 B.n430 VSUBS 0.007956f
C471 B.n431 VSUBS 0.007956f
C472 B.n432 VSUBS 0.007956f
C473 B.n433 VSUBS 0.007956f
C474 B.n434 VSUBS 0.007956f
C475 B.n435 VSUBS 0.007956f
C476 B.n436 VSUBS 0.007956f
C477 B.n437 VSUBS 0.007956f
C478 B.n438 VSUBS 0.007956f
C479 B.n439 VSUBS 0.007956f
C480 B.n440 VSUBS 0.007956f
C481 B.n441 VSUBS 0.007956f
C482 B.n442 VSUBS 0.007956f
C483 B.n443 VSUBS 0.007956f
C484 B.n444 VSUBS 0.007956f
C485 B.n445 VSUBS 0.007956f
C486 B.n446 VSUBS 0.007956f
C487 B.n447 VSUBS 0.007956f
C488 B.n448 VSUBS 0.007956f
C489 B.n449 VSUBS 0.007956f
C490 B.n450 VSUBS 0.007956f
C491 B.n451 VSUBS 0.007956f
C492 B.n452 VSUBS 0.007956f
C493 B.n453 VSUBS 0.007956f
C494 B.n454 VSUBS 0.007956f
C495 B.n455 VSUBS 0.007956f
C496 B.n456 VSUBS 0.007956f
C497 B.n457 VSUBS 0.007956f
C498 B.n458 VSUBS 0.007956f
C499 B.n459 VSUBS 0.007956f
C500 B.n460 VSUBS 0.007956f
C501 B.n461 VSUBS 0.007956f
C502 B.n462 VSUBS 0.007488f
C503 B.n463 VSUBS 0.018434f
C504 B.n464 VSUBS 0.004446f
C505 B.n465 VSUBS 0.007956f
C506 B.n466 VSUBS 0.007956f
C507 B.n467 VSUBS 0.007956f
C508 B.n468 VSUBS 0.007956f
C509 B.n469 VSUBS 0.007956f
C510 B.n470 VSUBS 0.007956f
C511 B.n471 VSUBS 0.007956f
C512 B.n472 VSUBS 0.007956f
C513 B.n473 VSUBS 0.007956f
C514 B.n474 VSUBS 0.007956f
C515 B.n475 VSUBS 0.007956f
C516 B.n476 VSUBS 0.007956f
C517 B.n477 VSUBS 0.004446f
C518 B.n478 VSUBS 0.007956f
C519 B.n479 VSUBS 0.007956f
C520 B.n480 VSUBS 0.007956f
C521 B.n481 VSUBS 0.007956f
C522 B.n482 VSUBS 0.007956f
C523 B.n483 VSUBS 0.007956f
C524 B.n484 VSUBS 0.007956f
C525 B.n485 VSUBS 0.007956f
C526 B.n486 VSUBS 0.007956f
C527 B.n487 VSUBS 0.007956f
C528 B.n488 VSUBS 0.007956f
C529 B.n489 VSUBS 0.007956f
C530 B.n490 VSUBS 0.007956f
C531 B.n491 VSUBS 0.007956f
C532 B.n492 VSUBS 0.007956f
C533 B.n493 VSUBS 0.007956f
C534 B.n494 VSUBS 0.007956f
C535 B.n495 VSUBS 0.007956f
C536 B.n496 VSUBS 0.007956f
C537 B.n497 VSUBS 0.007956f
C538 B.n498 VSUBS 0.007956f
C539 B.n499 VSUBS 0.007956f
C540 B.n500 VSUBS 0.007956f
C541 B.n501 VSUBS 0.007956f
C542 B.n502 VSUBS 0.007956f
C543 B.n503 VSUBS 0.007956f
C544 B.n504 VSUBS 0.007956f
C545 B.n505 VSUBS 0.007956f
C546 B.n506 VSUBS 0.007956f
C547 B.n507 VSUBS 0.007956f
C548 B.n508 VSUBS 0.007956f
C549 B.n509 VSUBS 0.007956f
C550 B.n510 VSUBS 0.007956f
C551 B.n511 VSUBS 0.007956f
C552 B.n512 VSUBS 0.007956f
C553 B.n513 VSUBS 0.007956f
C554 B.n514 VSUBS 0.007956f
C555 B.n515 VSUBS 0.007956f
C556 B.n516 VSUBS 0.007956f
C557 B.n517 VSUBS 0.007956f
C558 B.n518 VSUBS 0.007956f
C559 B.n519 VSUBS 0.007956f
C560 B.n520 VSUBS 0.007956f
C561 B.n521 VSUBS 0.007956f
C562 B.n522 VSUBS 0.007956f
C563 B.n523 VSUBS 0.007956f
C564 B.n524 VSUBS 0.007956f
C565 B.n525 VSUBS 0.007956f
C566 B.n526 VSUBS 0.007956f
C567 B.n527 VSUBS 0.007956f
C568 B.n528 VSUBS 0.01799f
C569 B.n529 VSUBS 0.01799f
C570 B.n530 VSUBS 0.017111f
C571 B.n531 VSUBS 0.007956f
C572 B.n532 VSUBS 0.007956f
C573 B.n533 VSUBS 0.007956f
C574 B.n534 VSUBS 0.007956f
C575 B.n535 VSUBS 0.007956f
C576 B.n536 VSUBS 0.007956f
C577 B.n537 VSUBS 0.007956f
C578 B.n538 VSUBS 0.007956f
C579 B.n539 VSUBS 0.007956f
C580 B.n540 VSUBS 0.007956f
C581 B.n541 VSUBS 0.007956f
C582 B.n542 VSUBS 0.007956f
C583 B.n543 VSUBS 0.007956f
C584 B.n544 VSUBS 0.007956f
C585 B.n545 VSUBS 0.007956f
C586 B.n546 VSUBS 0.007956f
C587 B.n547 VSUBS 0.007956f
C588 B.n548 VSUBS 0.007956f
C589 B.n549 VSUBS 0.007956f
C590 B.n550 VSUBS 0.007956f
C591 B.n551 VSUBS 0.007956f
C592 B.n552 VSUBS 0.007956f
C593 B.n553 VSUBS 0.007956f
C594 B.n554 VSUBS 0.007956f
C595 B.n555 VSUBS 0.007956f
C596 B.n556 VSUBS 0.007956f
C597 B.n557 VSUBS 0.007956f
C598 B.n558 VSUBS 0.007956f
C599 B.n559 VSUBS 0.007956f
C600 B.n560 VSUBS 0.007956f
C601 B.n561 VSUBS 0.007956f
C602 B.n562 VSUBS 0.007956f
C603 B.n563 VSUBS 0.007956f
C604 B.n564 VSUBS 0.007956f
C605 B.n565 VSUBS 0.007956f
C606 B.n566 VSUBS 0.007956f
C607 B.n567 VSUBS 0.007956f
C608 B.n568 VSUBS 0.007956f
C609 B.n569 VSUBS 0.007956f
C610 B.n570 VSUBS 0.007956f
C611 B.n571 VSUBS 0.007956f
C612 B.n572 VSUBS 0.007956f
C613 B.n573 VSUBS 0.007956f
C614 B.n574 VSUBS 0.007956f
C615 B.n575 VSUBS 0.010382f
C616 B.n576 VSUBS 0.01106f
C617 B.n577 VSUBS 0.021994f
C618 VDD1.t4 VSUBS 0.190416f
C619 VDD1.t2 VSUBS 0.190416f
C620 VDD1.n0 VSUBS 1.43815f
C621 VDD1.t0 VSUBS 0.190416f
C622 VDD1.t1 VSUBS 0.190416f
C623 VDD1.n1 VSUBS 1.43723f
C624 VDD1.t7 VSUBS 0.190416f
C625 VDD1.t3 VSUBS 0.190416f
C626 VDD1.n2 VSUBS 1.43723f
C627 VDD1.n3 VSUBS 2.90471f
C628 VDD1.t5 VSUBS 0.190416f
C629 VDD1.t6 VSUBS 0.190416f
C630 VDD1.n4 VSUBS 1.43258f
C631 VDD1.n5 VSUBS 2.59337f
C632 VP.n0 VSUBS 0.060775f
C633 VP.t0 VSUBS 1.45457f
C634 VP.n1 VSUBS 0.544491f
C635 VP.n2 VSUBS 0.045546f
C636 VP.t6 VSUBS 1.45457f
C637 VP.n3 VSUBS 0.544491f
C638 VP.n4 VSUBS 0.060775f
C639 VP.n5 VSUBS 0.060775f
C640 VP.t1 VSUBS 1.54179f
C641 VP.t2 VSUBS 1.45457f
C642 VP.n6 VSUBS 0.544491f
C643 VP.n7 VSUBS 0.045546f
C644 VP.t5 VSUBS 1.45457f
C645 VP.n8 VSUBS 0.605867f
C646 VP.t3 VSUBS 1.597f
C647 VP.n9 VSUBS 0.620473f
C648 VP.n10 VSUBS 0.239305f
C649 VP.n11 VSUBS 0.07292f
C650 VP.n12 VSUBS 0.036819f
C651 VP.n13 VSUBS 0.07292f
C652 VP.n14 VSUBS 0.045546f
C653 VP.n15 VSUBS 0.045546f
C654 VP.n16 VSUBS 0.067554f
C655 VP.n17 VSUBS 0.033402f
C656 VP.n18 VSUBS 0.633922f
C657 VP.n19 VSUBS 1.95789f
C658 VP.n20 VSUBS 1.99612f
C659 VP.t7 VSUBS 1.54179f
C660 VP.n21 VSUBS 0.633922f
C661 VP.n22 VSUBS 0.033402f
C662 VP.n23 VSUBS 0.067554f
C663 VP.n24 VSUBS 0.045546f
C664 VP.n25 VSUBS 0.045546f
C665 VP.n26 VSUBS 0.07292f
C666 VP.n27 VSUBS 0.036819f
C667 VP.n28 VSUBS 0.07292f
C668 VP.n29 VSUBS 0.045546f
C669 VP.n30 VSUBS 0.045546f
C670 VP.n31 VSUBS 0.067554f
C671 VP.n32 VSUBS 0.033402f
C672 VP.t4 VSUBS 1.54179f
C673 VP.n33 VSUBS 0.633922f
C674 VP.n34 VSUBS 0.042655f
C675 VTAIL.t9 VSUBS 0.18798f
C676 VTAIL.t7 VSUBS 0.18798f
C677 VTAIL.n0 VSUBS 1.30462f
C678 VTAIL.n1 VSUBS 0.629073f
C679 VTAIL.n2 VSUBS 0.028087f
C680 VTAIL.n3 VSUBS 0.025172f
C681 VTAIL.n4 VSUBS 0.013527f
C682 VTAIL.n5 VSUBS 0.031972f
C683 VTAIL.n6 VSUBS 0.013924f
C684 VTAIL.n7 VSUBS 0.025172f
C685 VTAIL.n8 VSUBS 0.014322f
C686 VTAIL.n9 VSUBS 0.031972f
C687 VTAIL.n10 VSUBS 0.014322f
C688 VTAIL.n11 VSUBS 0.025172f
C689 VTAIL.n12 VSUBS 0.013527f
C690 VTAIL.n13 VSUBS 0.031972f
C691 VTAIL.n14 VSUBS 0.014322f
C692 VTAIL.n15 VSUBS 0.955455f
C693 VTAIL.n16 VSUBS 0.013527f
C694 VTAIL.t10 VSUBS 0.068729f
C695 VTAIL.n17 VSUBS 0.169266f
C696 VTAIL.n18 VSUBS 0.024051f
C697 VTAIL.n19 VSUBS 0.023979f
C698 VTAIL.n20 VSUBS 0.031972f
C699 VTAIL.n21 VSUBS 0.014322f
C700 VTAIL.n22 VSUBS 0.013527f
C701 VTAIL.n23 VSUBS 0.025172f
C702 VTAIL.n24 VSUBS 0.025172f
C703 VTAIL.n25 VSUBS 0.013527f
C704 VTAIL.n26 VSUBS 0.014322f
C705 VTAIL.n27 VSUBS 0.031972f
C706 VTAIL.n28 VSUBS 0.031972f
C707 VTAIL.n29 VSUBS 0.014322f
C708 VTAIL.n30 VSUBS 0.013527f
C709 VTAIL.n31 VSUBS 0.025172f
C710 VTAIL.n32 VSUBS 0.025172f
C711 VTAIL.n33 VSUBS 0.013527f
C712 VTAIL.n34 VSUBS 0.013527f
C713 VTAIL.n35 VSUBS 0.014322f
C714 VTAIL.n36 VSUBS 0.031972f
C715 VTAIL.n37 VSUBS 0.031972f
C716 VTAIL.n38 VSUBS 0.031972f
C717 VTAIL.n39 VSUBS 0.013924f
C718 VTAIL.n40 VSUBS 0.013527f
C719 VTAIL.n41 VSUBS 0.025172f
C720 VTAIL.n42 VSUBS 0.025172f
C721 VTAIL.n43 VSUBS 0.013527f
C722 VTAIL.n44 VSUBS 0.014322f
C723 VTAIL.n45 VSUBS 0.031972f
C724 VTAIL.n46 VSUBS 0.078859f
C725 VTAIL.n47 VSUBS 0.014322f
C726 VTAIL.n48 VSUBS 0.013527f
C727 VTAIL.n49 VSUBS 0.065406f
C728 VTAIL.n50 VSUBS 0.039933f
C729 VTAIL.n51 VSUBS 0.174174f
C730 VTAIL.n52 VSUBS 0.028087f
C731 VTAIL.n53 VSUBS 0.025172f
C732 VTAIL.n54 VSUBS 0.013527f
C733 VTAIL.n55 VSUBS 0.031972f
C734 VTAIL.n56 VSUBS 0.013924f
C735 VTAIL.n57 VSUBS 0.025172f
C736 VTAIL.n58 VSUBS 0.014322f
C737 VTAIL.n59 VSUBS 0.031972f
C738 VTAIL.n60 VSUBS 0.014322f
C739 VTAIL.n61 VSUBS 0.025172f
C740 VTAIL.n62 VSUBS 0.013527f
C741 VTAIL.n63 VSUBS 0.031972f
C742 VTAIL.n64 VSUBS 0.014322f
C743 VTAIL.n65 VSUBS 0.955455f
C744 VTAIL.n66 VSUBS 0.013527f
C745 VTAIL.t1 VSUBS 0.068729f
C746 VTAIL.n67 VSUBS 0.169266f
C747 VTAIL.n68 VSUBS 0.024051f
C748 VTAIL.n69 VSUBS 0.023979f
C749 VTAIL.n70 VSUBS 0.031972f
C750 VTAIL.n71 VSUBS 0.014322f
C751 VTAIL.n72 VSUBS 0.013527f
C752 VTAIL.n73 VSUBS 0.025172f
C753 VTAIL.n74 VSUBS 0.025172f
C754 VTAIL.n75 VSUBS 0.013527f
C755 VTAIL.n76 VSUBS 0.014322f
C756 VTAIL.n77 VSUBS 0.031972f
C757 VTAIL.n78 VSUBS 0.031972f
C758 VTAIL.n79 VSUBS 0.014322f
C759 VTAIL.n80 VSUBS 0.013527f
C760 VTAIL.n81 VSUBS 0.025172f
C761 VTAIL.n82 VSUBS 0.025172f
C762 VTAIL.n83 VSUBS 0.013527f
C763 VTAIL.n84 VSUBS 0.013527f
C764 VTAIL.n85 VSUBS 0.014322f
C765 VTAIL.n86 VSUBS 0.031972f
C766 VTAIL.n87 VSUBS 0.031972f
C767 VTAIL.n88 VSUBS 0.031972f
C768 VTAIL.n89 VSUBS 0.013924f
C769 VTAIL.n90 VSUBS 0.013527f
C770 VTAIL.n91 VSUBS 0.025172f
C771 VTAIL.n92 VSUBS 0.025172f
C772 VTAIL.n93 VSUBS 0.013527f
C773 VTAIL.n94 VSUBS 0.014322f
C774 VTAIL.n95 VSUBS 0.031972f
C775 VTAIL.n96 VSUBS 0.078859f
C776 VTAIL.n97 VSUBS 0.014322f
C777 VTAIL.n98 VSUBS 0.013527f
C778 VTAIL.n99 VSUBS 0.065406f
C779 VTAIL.n100 VSUBS 0.039933f
C780 VTAIL.n101 VSUBS 0.174174f
C781 VTAIL.t4 VSUBS 0.18798f
C782 VTAIL.t5 VSUBS 0.18798f
C783 VTAIL.n102 VSUBS 1.30462f
C784 VTAIL.n103 VSUBS 0.734832f
C785 VTAIL.n104 VSUBS 0.028087f
C786 VTAIL.n105 VSUBS 0.025172f
C787 VTAIL.n106 VSUBS 0.013527f
C788 VTAIL.n107 VSUBS 0.031972f
C789 VTAIL.n108 VSUBS 0.013924f
C790 VTAIL.n109 VSUBS 0.025172f
C791 VTAIL.n110 VSUBS 0.014322f
C792 VTAIL.n111 VSUBS 0.031972f
C793 VTAIL.n112 VSUBS 0.014322f
C794 VTAIL.n113 VSUBS 0.025172f
C795 VTAIL.n114 VSUBS 0.013527f
C796 VTAIL.n115 VSUBS 0.031972f
C797 VTAIL.n116 VSUBS 0.014322f
C798 VTAIL.n117 VSUBS 0.955455f
C799 VTAIL.n118 VSUBS 0.013527f
C800 VTAIL.t0 VSUBS 0.068729f
C801 VTAIL.n119 VSUBS 0.169266f
C802 VTAIL.n120 VSUBS 0.024051f
C803 VTAIL.n121 VSUBS 0.023979f
C804 VTAIL.n122 VSUBS 0.031972f
C805 VTAIL.n123 VSUBS 0.014322f
C806 VTAIL.n124 VSUBS 0.013527f
C807 VTAIL.n125 VSUBS 0.025172f
C808 VTAIL.n126 VSUBS 0.025172f
C809 VTAIL.n127 VSUBS 0.013527f
C810 VTAIL.n128 VSUBS 0.014322f
C811 VTAIL.n129 VSUBS 0.031972f
C812 VTAIL.n130 VSUBS 0.031972f
C813 VTAIL.n131 VSUBS 0.014322f
C814 VTAIL.n132 VSUBS 0.013527f
C815 VTAIL.n133 VSUBS 0.025172f
C816 VTAIL.n134 VSUBS 0.025172f
C817 VTAIL.n135 VSUBS 0.013527f
C818 VTAIL.n136 VSUBS 0.013527f
C819 VTAIL.n137 VSUBS 0.014322f
C820 VTAIL.n138 VSUBS 0.031972f
C821 VTAIL.n139 VSUBS 0.031972f
C822 VTAIL.n140 VSUBS 0.031972f
C823 VTAIL.n141 VSUBS 0.013924f
C824 VTAIL.n142 VSUBS 0.013527f
C825 VTAIL.n143 VSUBS 0.025172f
C826 VTAIL.n144 VSUBS 0.025172f
C827 VTAIL.n145 VSUBS 0.013527f
C828 VTAIL.n146 VSUBS 0.014322f
C829 VTAIL.n147 VSUBS 0.031972f
C830 VTAIL.n148 VSUBS 0.078859f
C831 VTAIL.n149 VSUBS 0.014322f
C832 VTAIL.n150 VSUBS 0.013527f
C833 VTAIL.n151 VSUBS 0.065406f
C834 VTAIL.n152 VSUBS 0.039933f
C835 VTAIL.n153 VSUBS 1.24926f
C836 VTAIL.n154 VSUBS 0.028087f
C837 VTAIL.n155 VSUBS 0.025172f
C838 VTAIL.n156 VSUBS 0.013527f
C839 VTAIL.n157 VSUBS 0.031972f
C840 VTAIL.n158 VSUBS 0.013924f
C841 VTAIL.n159 VSUBS 0.025172f
C842 VTAIL.n160 VSUBS 0.013924f
C843 VTAIL.n161 VSUBS 0.013527f
C844 VTAIL.n162 VSUBS 0.031972f
C845 VTAIL.n163 VSUBS 0.031972f
C846 VTAIL.n164 VSUBS 0.014322f
C847 VTAIL.n165 VSUBS 0.025172f
C848 VTAIL.n166 VSUBS 0.013527f
C849 VTAIL.n167 VSUBS 0.031972f
C850 VTAIL.n168 VSUBS 0.014322f
C851 VTAIL.n169 VSUBS 0.955455f
C852 VTAIL.n170 VSUBS 0.013527f
C853 VTAIL.t14 VSUBS 0.068729f
C854 VTAIL.n171 VSUBS 0.169266f
C855 VTAIL.n172 VSUBS 0.024051f
C856 VTAIL.n173 VSUBS 0.023979f
C857 VTAIL.n174 VSUBS 0.031972f
C858 VTAIL.n175 VSUBS 0.014322f
C859 VTAIL.n176 VSUBS 0.013527f
C860 VTAIL.n177 VSUBS 0.025172f
C861 VTAIL.n178 VSUBS 0.025172f
C862 VTAIL.n179 VSUBS 0.013527f
C863 VTAIL.n180 VSUBS 0.014322f
C864 VTAIL.n181 VSUBS 0.031972f
C865 VTAIL.n182 VSUBS 0.031972f
C866 VTAIL.n183 VSUBS 0.014322f
C867 VTAIL.n184 VSUBS 0.013527f
C868 VTAIL.n185 VSUBS 0.025172f
C869 VTAIL.n186 VSUBS 0.025172f
C870 VTAIL.n187 VSUBS 0.013527f
C871 VTAIL.n188 VSUBS 0.014322f
C872 VTAIL.n189 VSUBS 0.031972f
C873 VTAIL.n190 VSUBS 0.031972f
C874 VTAIL.n191 VSUBS 0.014322f
C875 VTAIL.n192 VSUBS 0.013527f
C876 VTAIL.n193 VSUBS 0.025172f
C877 VTAIL.n194 VSUBS 0.025172f
C878 VTAIL.n195 VSUBS 0.013527f
C879 VTAIL.n196 VSUBS 0.014322f
C880 VTAIL.n197 VSUBS 0.031972f
C881 VTAIL.n198 VSUBS 0.078859f
C882 VTAIL.n199 VSUBS 0.014322f
C883 VTAIL.n200 VSUBS 0.013527f
C884 VTAIL.n201 VSUBS 0.065406f
C885 VTAIL.n202 VSUBS 0.039933f
C886 VTAIL.n203 VSUBS 1.24926f
C887 VTAIL.t13 VSUBS 0.18798f
C888 VTAIL.t12 VSUBS 0.18798f
C889 VTAIL.n204 VSUBS 1.30463f
C890 VTAIL.n205 VSUBS 0.734823f
C891 VTAIL.n206 VSUBS 0.028087f
C892 VTAIL.n207 VSUBS 0.025172f
C893 VTAIL.n208 VSUBS 0.013527f
C894 VTAIL.n209 VSUBS 0.031972f
C895 VTAIL.n210 VSUBS 0.013924f
C896 VTAIL.n211 VSUBS 0.025172f
C897 VTAIL.n212 VSUBS 0.013924f
C898 VTAIL.n213 VSUBS 0.013527f
C899 VTAIL.n214 VSUBS 0.031972f
C900 VTAIL.n215 VSUBS 0.031972f
C901 VTAIL.n216 VSUBS 0.014322f
C902 VTAIL.n217 VSUBS 0.025172f
C903 VTAIL.n218 VSUBS 0.013527f
C904 VTAIL.n219 VSUBS 0.031972f
C905 VTAIL.n220 VSUBS 0.014322f
C906 VTAIL.n221 VSUBS 0.955455f
C907 VTAIL.n222 VSUBS 0.013527f
C908 VTAIL.t11 VSUBS 0.068729f
C909 VTAIL.n223 VSUBS 0.169266f
C910 VTAIL.n224 VSUBS 0.024051f
C911 VTAIL.n225 VSUBS 0.023979f
C912 VTAIL.n226 VSUBS 0.031972f
C913 VTAIL.n227 VSUBS 0.014322f
C914 VTAIL.n228 VSUBS 0.013527f
C915 VTAIL.n229 VSUBS 0.025172f
C916 VTAIL.n230 VSUBS 0.025172f
C917 VTAIL.n231 VSUBS 0.013527f
C918 VTAIL.n232 VSUBS 0.014322f
C919 VTAIL.n233 VSUBS 0.031972f
C920 VTAIL.n234 VSUBS 0.031972f
C921 VTAIL.n235 VSUBS 0.014322f
C922 VTAIL.n236 VSUBS 0.013527f
C923 VTAIL.n237 VSUBS 0.025172f
C924 VTAIL.n238 VSUBS 0.025172f
C925 VTAIL.n239 VSUBS 0.013527f
C926 VTAIL.n240 VSUBS 0.014322f
C927 VTAIL.n241 VSUBS 0.031972f
C928 VTAIL.n242 VSUBS 0.031972f
C929 VTAIL.n243 VSUBS 0.014322f
C930 VTAIL.n244 VSUBS 0.013527f
C931 VTAIL.n245 VSUBS 0.025172f
C932 VTAIL.n246 VSUBS 0.025172f
C933 VTAIL.n247 VSUBS 0.013527f
C934 VTAIL.n248 VSUBS 0.014322f
C935 VTAIL.n249 VSUBS 0.031972f
C936 VTAIL.n250 VSUBS 0.078859f
C937 VTAIL.n251 VSUBS 0.014322f
C938 VTAIL.n252 VSUBS 0.013527f
C939 VTAIL.n253 VSUBS 0.065406f
C940 VTAIL.n254 VSUBS 0.039933f
C941 VTAIL.n255 VSUBS 0.174174f
C942 VTAIL.n256 VSUBS 0.028087f
C943 VTAIL.n257 VSUBS 0.025172f
C944 VTAIL.n258 VSUBS 0.013527f
C945 VTAIL.n259 VSUBS 0.031972f
C946 VTAIL.n260 VSUBS 0.013924f
C947 VTAIL.n261 VSUBS 0.025172f
C948 VTAIL.n262 VSUBS 0.013924f
C949 VTAIL.n263 VSUBS 0.013527f
C950 VTAIL.n264 VSUBS 0.031972f
C951 VTAIL.n265 VSUBS 0.031972f
C952 VTAIL.n266 VSUBS 0.014322f
C953 VTAIL.n267 VSUBS 0.025172f
C954 VTAIL.n268 VSUBS 0.013527f
C955 VTAIL.n269 VSUBS 0.031972f
C956 VTAIL.n270 VSUBS 0.014322f
C957 VTAIL.n271 VSUBS 0.955455f
C958 VTAIL.n272 VSUBS 0.013527f
C959 VTAIL.t3 VSUBS 0.068729f
C960 VTAIL.n273 VSUBS 0.169266f
C961 VTAIL.n274 VSUBS 0.024051f
C962 VTAIL.n275 VSUBS 0.023979f
C963 VTAIL.n276 VSUBS 0.031972f
C964 VTAIL.n277 VSUBS 0.014322f
C965 VTAIL.n278 VSUBS 0.013527f
C966 VTAIL.n279 VSUBS 0.025172f
C967 VTAIL.n280 VSUBS 0.025172f
C968 VTAIL.n281 VSUBS 0.013527f
C969 VTAIL.n282 VSUBS 0.014322f
C970 VTAIL.n283 VSUBS 0.031972f
C971 VTAIL.n284 VSUBS 0.031972f
C972 VTAIL.n285 VSUBS 0.014322f
C973 VTAIL.n286 VSUBS 0.013527f
C974 VTAIL.n287 VSUBS 0.025172f
C975 VTAIL.n288 VSUBS 0.025172f
C976 VTAIL.n289 VSUBS 0.013527f
C977 VTAIL.n290 VSUBS 0.014322f
C978 VTAIL.n291 VSUBS 0.031972f
C979 VTAIL.n292 VSUBS 0.031972f
C980 VTAIL.n293 VSUBS 0.014322f
C981 VTAIL.n294 VSUBS 0.013527f
C982 VTAIL.n295 VSUBS 0.025172f
C983 VTAIL.n296 VSUBS 0.025172f
C984 VTAIL.n297 VSUBS 0.013527f
C985 VTAIL.n298 VSUBS 0.014322f
C986 VTAIL.n299 VSUBS 0.031972f
C987 VTAIL.n300 VSUBS 0.078859f
C988 VTAIL.n301 VSUBS 0.014322f
C989 VTAIL.n302 VSUBS 0.013527f
C990 VTAIL.n303 VSUBS 0.065406f
C991 VTAIL.n304 VSUBS 0.039933f
C992 VTAIL.n305 VSUBS 0.174174f
C993 VTAIL.t2 VSUBS 0.18798f
C994 VTAIL.t6 VSUBS 0.18798f
C995 VTAIL.n306 VSUBS 1.30463f
C996 VTAIL.n307 VSUBS 0.734823f
C997 VTAIL.n308 VSUBS 0.028087f
C998 VTAIL.n309 VSUBS 0.025172f
C999 VTAIL.n310 VSUBS 0.013527f
C1000 VTAIL.n311 VSUBS 0.031972f
C1001 VTAIL.n312 VSUBS 0.013924f
C1002 VTAIL.n313 VSUBS 0.025172f
C1003 VTAIL.n314 VSUBS 0.013924f
C1004 VTAIL.n315 VSUBS 0.013527f
C1005 VTAIL.n316 VSUBS 0.031972f
C1006 VTAIL.n317 VSUBS 0.031972f
C1007 VTAIL.n318 VSUBS 0.014322f
C1008 VTAIL.n319 VSUBS 0.025172f
C1009 VTAIL.n320 VSUBS 0.013527f
C1010 VTAIL.n321 VSUBS 0.031972f
C1011 VTAIL.n322 VSUBS 0.014322f
C1012 VTAIL.n323 VSUBS 0.955455f
C1013 VTAIL.n324 VSUBS 0.013527f
C1014 VTAIL.t15 VSUBS 0.068729f
C1015 VTAIL.n325 VSUBS 0.169266f
C1016 VTAIL.n326 VSUBS 0.024051f
C1017 VTAIL.n327 VSUBS 0.023979f
C1018 VTAIL.n328 VSUBS 0.031972f
C1019 VTAIL.n329 VSUBS 0.014322f
C1020 VTAIL.n330 VSUBS 0.013527f
C1021 VTAIL.n331 VSUBS 0.025172f
C1022 VTAIL.n332 VSUBS 0.025172f
C1023 VTAIL.n333 VSUBS 0.013527f
C1024 VTAIL.n334 VSUBS 0.014322f
C1025 VTAIL.n335 VSUBS 0.031972f
C1026 VTAIL.n336 VSUBS 0.031972f
C1027 VTAIL.n337 VSUBS 0.014322f
C1028 VTAIL.n338 VSUBS 0.013527f
C1029 VTAIL.n339 VSUBS 0.025172f
C1030 VTAIL.n340 VSUBS 0.025172f
C1031 VTAIL.n341 VSUBS 0.013527f
C1032 VTAIL.n342 VSUBS 0.014322f
C1033 VTAIL.n343 VSUBS 0.031972f
C1034 VTAIL.n344 VSUBS 0.031972f
C1035 VTAIL.n345 VSUBS 0.014322f
C1036 VTAIL.n346 VSUBS 0.013527f
C1037 VTAIL.n347 VSUBS 0.025172f
C1038 VTAIL.n348 VSUBS 0.025172f
C1039 VTAIL.n349 VSUBS 0.013527f
C1040 VTAIL.n350 VSUBS 0.014322f
C1041 VTAIL.n351 VSUBS 0.031972f
C1042 VTAIL.n352 VSUBS 0.078859f
C1043 VTAIL.n353 VSUBS 0.014322f
C1044 VTAIL.n354 VSUBS 0.013527f
C1045 VTAIL.n355 VSUBS 0.065406f
C1046 VTAIL.n356 VSUBS 0.039933f
C1047 VTAIL.n357 VSUBS 1.24926f
C1048 VTAIL.n358 VSUBS 0.028087f
C1049 VTAIL.n359 VSUBS 0.025172f
C1050 VTAIL.n360 VSUBS 0.013527f
C1051 VTAIL.n361 VSUBS 0.031972f
C1052 VTAIL.n362 VSUBS 0.013924f
C1053 VTAIL.n363 VSUBS 0.025172f
C1054 VTAIL.n364 VSUBS 0.014322f
C1055 VTAIL.n365 VSUBS 0.031972f
C1056 VTAIL.n366 VSUBS 0.014322f
C1057 VTAIL.n367 VSUBS 0.025172f
C1058 VTAIL.n368 VSUBS 0.013527f
C1059 VTAIL.n369 VSUBS 0.031972f
C1060 VTAIL.n370 VSUBS 0.014322f
C1061 VTAIL.n371 VSUBS 0.955455f
C1062 VTAIL.n372 VSUBS 0.013527f
C1063 VTAIL.t8 VSUBS 0.068729f
C1064 VTAIL.n373 VSUBS 0.169266f
C1065 VTAIL.n374 VSUBS 0.024051f
C1066 VTAIL.n375 VSUBS 0.023979f
C1067 VTAIL.n376 VSUBS 0.031972f
C1068 VTAIL.n377 VSUBS 0.014322f
C1069 VTAIL.n378 VSUBS 0.013527f
C1070 VTAIL.n379 VSUBS 0.025172f
C1071 VTAIL.n380 VSUBS 0.025172f
C1072 VTAIL.n381 VSUBS 0.013527f
C1073 VTAIL.n382 VSUBS 0.014322f
C1074 VTAIL.n383 VSUBS 0.031972f
C1075 VTAIL.n384 VSUBS 0.031972f
C1076 VTAIL.n385 VSUBS 0.014322f
C1077 VTAIL.n386 VSUBS 0.013527f
C1078 VTAIL.n387 VSUBS 0.025172f
C1079 VTAIL.n388 VSUBS 0.025172f
C1080 VTAIL.n389 VSUBS 0.013527f
C1081 VTAIL.n390 VSUBS 0.013527f
C1082 VTAIL.n391 VSUBS 0.014322f
C1083 VTAIL.n392 VSUBS 0.031972f
C1084 VTAIL.n393 VSUBS 0.031972f
C1085 VTAIL.n394 VSUBS 0.031972f
C1086 VTAIL.n395 VSUBS 0.013924f
C1087 VTAIL.n396 VSUBS 0.013527f
C1088 VTAIL.n397 VSUBS 0.025172f
C1089 VTAIL.n398 VSUBS 0.025172f
C1090 VTAIL.n399 VSUBS 0.013527f
C1091 VTAIL.n400 VSUBS 0.014322f
C1092 VTAIL.n401 VSUBS 0.031972f
C1093 VTAIL.n402 VSUBS 0.078859f
C1094 VTAIL.n403 VSUBS 0.014322f
C1095 VTAIL.n404 VSUBS 0.013527f
C1096 VTAIL.n405 VSUBS 0.065406f
C1097 VTAIL.n406 VSUBS 0.039933f
C1098 VTAIL.n407 VSUBS 1.24454f
C1099 VDD2.t0 VSUBS 0.188913f
C1100 VDD2.t3 VSUBS 0.188913f
C1101 VDD2.n0 VSUBS 1.42589f
C1102 VDD2.t4 VSUBS 0.188913f
C1103 VDD2.t6 VSUBS 0.188913f
C1104 VDD2.n1 VSUBS 1.42589f
C1105 VDD2.n2 VSUBS 2.82811f
C1106 VDD2.t2 VSUBS 0.188913f
C1107 VDD2.t1 VSUBS 0.188913f
C1108 VDD2.n3 VSUBS 1.42128f
C1109 VDD2.n4 VSUBS 2.54262f
C1110 VDD2.t7 VSUBS 0.188913f
C1111 VDD2.t5 VSUBS 0.188913f
C1112 VDD2.n5 VSUBS 1.42586f
C1113 VN.n0 VSUBS 0.059242f
C1114 VN.t7 VSUBS 1.41788f
C1115 VN.n1 VSUBS 0.530759f
C1116 VN.n2 VSUBS 0.044397f
C1117 VN.t5 VSUBS 1.41788f
C1118 VN.n3 VSUBS 0.590587f
C1119 VN.t4 VSUBS 1.55672f
C1120 VN.n4 VSUBS 0.604825f
C1121 VN.n5 VSUBS 0.233269f
C1122 VN.n6 VSUBS 0.071081f
C1123 VN.n7 VSUBS 0.035891f
C1124 VN.n8 VSUBS 0.071081f
C1125 VN.n9 VSUBS 0.044397f
C1126 VN.n10 VSUBS 0.044397f
C1127 VN.n11 VSUBS 0.06585f
C1128 VN.n12 VSUBS 0.03256f
C1129 VN.t6 VSUBS 1.5029f
C1130 VN.n13 VSUBS 0.617934f
C1131 VN.n14 VSUBS 0.041579f
C1132 VN.n15 VSUBS 0.059242f
C1133 VN.t1 VSUBS 1.41788f
C1134 VN.n16 VSUBS 0.530759f
C1135 VN.n17 VSUBS 0.044397f
C1136 VN.t2 VSUBS 1.41788f
C1137 VN.n18 VSUBS 0.590587f
C1138 VN.t3 VSUBS 1.55672f
C1139 VN.n19 VSUBS 0.604825f
C1140 VN.n20 VSUBS 0.233269f
C1141 VN.n21 VSUBS 0.071081f
C1142 VN.n22 VSUBS 0.035891f
C1143 VN.n23 VSUBS 0.071081f
C1144 VN.n24 VSUBS 0.044397f
C1145 VN.n25 VSUBS 0.044397f
C1146 VN.n26 VSUBS 0.06585f
C1147 VN.n27 VSUBS 0.03256f
C1148 VN.t0 VSUBS 1.5029f
C1149 VN.n28 VSUBS 0.617934f
C1150 VN.n29 VSUBS 1.93333f
.ends

