* NGSPICE file created from diff_pair_sample_1448.ext - technology: sky130A

.subckt diff_pair_sample_1448 VTAIL VN VP B VDD2 VDD1
X0 B.t11 B.t9 B.t10 w_n1878_n2178# sky130_fd_pr__pfet_01v8 ad=2.3595 pd=12.88 as=0 ps=0 w=6.05 l=1.94
X1 VDD1.t1 VP.t0 VTAIL.t3 w_n1878_n2178# sky130_fd_pr__pfet_01v8 ad=2.3595 pd=12.88 as=2.3595 ps=12.88 w=6.05 l=1.94
X2 B.t8 B.t6 B.t7 w_n1878_n2178# sky130_fd_pr__pfet_01v8 ad=2.3595 pd=12.88 as=0 ps=0 w=6.05 l=1.94
X3 VDD2.t1 VN.t0 VTAIL.t1 w_n1878_n2178# sky130_fd_pr__pfet_01v8 ad=2.3595 pd=12.88 as=2.3595 ps=12.88 w=6.05 l=1.94
X4 B.t5 B.t3 B.t4 w_n1878_n2178# sky130_fd_pr__pfet_01v8 ad=2.3595 pd=12.88 as=0 ps=0 w=6.05 l=1.94
X5 VDD1.t0 VP.t1 VTAIL.t2 w_n1878_n2178# sky130_fd_pr__pfet_01v8 ad=2.3595 pd=12.88 as=2.3595 ps=12.88 w=6.05 l=1.94
X6 VDD2.t0 VN.t1 VTAIL.t0 w_n1878_n2178# sky130_fd_pr__pfet_01v8 ad=2.3595 pd=12.88 as=2.3595 ps=12.88 w=6.05 l=1.94
X7 B.t2 B.t0 B.t1 w_n1878_n2178# sky130_fd_pr__pfet_01v8 ad=2.3595 pd=12.88 as=0 ps=0 w=6.05 l=1.94
R0 B.n230 B.n229 585
R1 B.n228 B.n69 585
R2 B.n227 B.n226 585
R3 B.n225 B.n70 585
R4 B.n224 B.n223 585
R5 B.n222 B.n71 585
R6 B.n221 B.n220 585
R7 B.n219 B.n72 585
R8 B.n218 B.n217 585
R9 B.n216 B.n73 585
R10 B.n215 B.n214 585
R11 B.n213 B.n74 585
R12 B.n212 B.n211 585
R13 B.n210 B.n75 585
R14 B.n209 B.n208 585
R15 B.n207 B.n76 585
R16 B.n206 B.n205 585
R17 B.n204 B.n77 585
R18 B.n203 B.n202 585
R19 B.n201 B.n78 585
R20 B.n200 B.n199 585
R21 B.n198 B.n79 585
R22 B.n197 B.n196 585
R23 B.n195 B.n80 585
R24 B.n193 B.n192 585
R25 B.n191 B.n83 585
R26 B.n190 B.n189 585
R27 B.n188 B.n84 585
R28 B.n187 B.n186 585
R29 B.n185 B.n85 585
R30 B.n184 B.n183 585
R31 B.n182 B.n86 585
R32 B.n181 B.n180 585
R33 B.n179 B.n87 585
R34 B.n178 B.n177 585
R35 B.n173 B.n88 585
R36 B.n172 B.n171 585
R37 B.n170 B.n89 585
R38 B.n169 B.n168 585
R39 B.n167 B.n90 585
R40 B.n166 B.n165 585
R41 B.n164 B.n91 585
R42 B.n163 B.n162 585
R43 B.n161 B.n92 585
R44 B.n160 B.n159 585
R45 B.n158 B.n93 585
R46 B.n157 B.n156 585
R47 B.n155 B.n94 585
R48 B.n154 B.n153 585
R49 B.n152 B.n95 585
R50 B.n151 B.n150 585
R51 B.n149 B.n96 585
R52 B.n148 B.n147 585
R53 B.n146 B.n97 585
R54 B.n145 B.n144 585
R55 B.n143 B.n98 585
R56 B.n142 B.n141 585
R57 B.n140 B.n99 585
R58 B.n231 B.n68 585
R59 B.n233 B.n232 585
R60 B.n234 B.n67 585
R61 B.n236 B.n235 585
R62 B.n237 B.n66 585
R63 B.n239 B.n238 585
R64 B.n240 B.n65 585
R65 B.n242 B.n241 585
R66 B.n243 B.n64 585
R67 B.n245 B.n244 585
R68 B.n246 B.n63 585
R69 B.n248 B.n247 585
R70 B.n249 B.n62 585
R71 B.n251 B.n250 585
R72 B.n252 B.n61 585
R73 B.n254 B.n253 585
R74 B.n255 B.n60 585
R75 B.n257 B.n256 585
R76 B.n258 B.n59 585
R77 B.n260 B.n259 585
R78 B.n261 B.n58 585
R79 B.n263 B.n262 585
R80 B.n264 B.n57 585
R81 B.n266 B.n265 585
R82 B.n267 B.n56 585
R83 B.n269 B.n268 585
R84 B.n270 B.n55 585
R85 B.n272 B.n271 585
R86 B.n273 B.n54 585
R87 B.n275 B.n274 585
R88 B.n276 B.n53 585
R89 B.n278 B.n277 585
R90 B.n279 B.n52 585
R91 B.n281 B.n280 585
R92 B.n282 B.n51 585
R93 B.n284 B.n283 585
R94 B.n285 B.n50 585
R95 B.n287 B.n286 585
R96 B.n288 B.n49 585
R97 B.n290 B.n289 585
R98 B.n291 B.n48 585
R99 B.n293 B.n292 585
R100 B.n294 B.n47 585
R101 B.n296 B.n295 585
R102 B.n384 B.n383 585
R103 B.n382 B.n13 585
R104 B.n381 B.n380 585
R105 B.n379 B.n14 585
R106 B.n378 B.n377 585
R107 B.n376 B.n15 585
R108 B.n375 B.n374 585
R109 B.n373 B.n16 585
R110 B.n372 B.n371 585
R111 B.n370 B.n17 585
R112 B.n369 B.n368 585
R113 B.n367 B.n18 585
R114 B.n366 B.n365 585
R115 B.n364 B.n19 585
R116 B.n363 B.n362 585
R117 B.n361 B.n20 585
R118 B.n360 B.n359 585
R119 B.n358 B.n21 585
R120 B.n357 B.n356 585
R121 B.n355 B.n22 585
R122 B.n354 B.n353 585
R123 B.n352 B.n23 585
R124 B.n351 B.n350 585
R125 B.n349 B.n24 585
R126 B.n348 B.n347 585
R127 B.n346 B.n25 585
R128 B.n345 B.n344 585
R129 B.n343 B.n29 585
R130 B.n342 B.n341 585
R131 B.n340 B.n30 585
R132 B.n339 B.n338 585
R133 B.n337 B.n31 585
R134 B.n336 B.n335 585
R135 B.n334 B.n32 585
R136 B.n332 B.n331 585
R137 B.n330 B.n35 585
R138 B.n329 B.n328 585
R139 B.n327 B.n36 585
R140 B.n326 B.n325 585
R141 B.n324 B.n37 585
R142 B.n323 B.n322 585
R143 B.n321 B.n38 585
R144 B.n320 B.n319 585
R145 B.n318 B.n39 585
R146 B.n317 B.n316 585
R147 B.n315 B.n40 585
R148 B.n314 B.n313 585
R149 B.n312 B.n41 585
R150 B.n311 B.n310 585
R151 B.n309 B.n42 585
R152 B.n308 B.n307 585
R153 B.n306 B.n43 585
R154 B.n305 B.n304 585
R155 B.n303 B.n44 585
R156 B.n302 B.n301 585
R157 B.n300 B.n45 585
R158 B.n299 B.n298 585
R159 B.n297 B.n46 585
R160 B.n385 B.n12 585
R161 B.n387 B.n386 585
R162 B.n388 B.n11 585
R163 B.n390 B.n389 585
R164 B.n391 B.n10 585
R165 B.n393 B.n392 585
R166 B.n394 B.n9 585
R167 B.n396 B.n395 585
R168 B.n397 B.n8 585
R169 B.n399 B.n398 585
R170 B.n400 B.n7 585
R171 B.n402 B.n401 585
R172 B.n403 B.n6 585
R173 B.n405 B.n404 585
R174 B.n406 B.n5 585
R175 B.n408 B.n407 585
R176 B.n409 B.n4 585
R177 B.n411 B.n410 585
R178 B.n412 B.n3 585
R179 B.n414 B.n413 585
R180 B.n415 B.n0 585
R181 B.n2 B.n1 585
R182 B.n110 B.n109 585
R183 B.n112 B.n111 585
R184 B.n113 B.n108 585
R185 B.n115 B.n114 585
R186 B.n116 B.n107 585
R187 B.n118 B.n117 585
R188 B.n119 B.n106 585
R189 B.n121 B.n120 585
R190 B.n122 B.n105 585
R191 B.n124 B.n123 585
R192 B.n125 B.n104 585
R193 B.n127 B.n126 585
R194 B.n128 B.n103 585
R195 B.n130 B.n129 585
R196 B.n131 B.n102 585
R197 B.n133 B.n132 585
R198 B.n134 B.n101 585
R199 B.n136 B.n135 585
R200 B.n137 B.n100 585
R201 B.n139 B.n138 585
R202 B.n140 B.n139 478.086
R203 B.n229 B.n68 478.086
R204 B.n295 B.n46 478.086
R205 B.n385 B.n384 478.086
R206 B.n81 B.t10 313.187
R207 B.n33 B.t8 313.187
R208 B.n174 B.t1 313.187
R209 B.n26 B.t5 313.187
R210 B.n174 B.t0 281.93
R211 B.n81 B.t9 281.93
R212 B.n33 B.t6 281.93
R213 B.n26 B.t3 281.93
R214 B.n82 B.t11 269.163
R215 B.n34 B.t7 269.163
R216 B.n175 B.t2 269.163
R217 B.n27 B.t4 269.163
R218 B.n417 B.n416 256.663
R219 B.n416 B.n415 235.042
R220 B.n416 B.n2 235.042
R221 B.n141 B.n140 163.367
R222 B.n141 B.n98 163.367
R223 B.n145 B.n98 163.367
R224 B.n146 B.n145 163.367
R225 B.n147 B.n146 163.367
R226 B.n147 B.n96 163.367
R227 B.n151 B.n96 163.367
R228 B.n152 B.n151 163.367
R229 B.n153 B.n152 163.367
R230 B.n153 B.n94 163.367
R231 B.n157 B.n94 163.367
R232 B.n158 B.n157 163.367
R233 B.n159 B.n158 163.367
R234 B.n159 B.n92 163.367
R235 B.n163 B.n92 163.367
R236 B.n164 B.n163 163.367
R237 B.n165 B.n164 163.367
R238 B.n165 B.n90 163.367
R239 B.n169 B.n90 163.367
R240 B.n170 B.n169 163.367
R241 B.n171 B.n170 163.367
R242 B.n171 B.n88 163.367
R243 B.n178 B.n88 163.367
R244 B.n179 B.n178 163.367
R245 B.n180 B.n179 163.367
R246 B.n180 B.n86 163.367
R247 B.n184 B.n86 163.367
R248 B.n185 B.n184 163.367
R249 B.n186 B.n185 163.367
R250 B.n186 B.n84 163.367
R251 B.n190 B.n84 163.367
R252 B.n191 B.n190 163.367
R253 B.n192 B.n191 163.367
R254 B.n192 B.n80 163.367
R255 B.n197 B.n80 163.367
R256 B.n198 B.n197 163.367
R257 B.n199 B.n198 163.367
R258 B.n199 B.n78 163.367
R259 B.n203 B.n78 163.367
R260 B.n204 B.n203 163.367
R261 B.n205 B.n204 163.367
R262 B.n205 B.n76 163.367
R263 B.n209 B.n76 163.367
R264 B.n210 B.n209 163.367
R265 B.n211 B.n210 163.367
R266 B.n211 B.n74 163.367
R267 B.n215 B.n74 163.367
R268 B.n216 B.n215 163.367
R269 B.n217 B.n216 163.367
R270 B.n217 B.n72 163.367
R271 B.n221 B.n72 163.367
R272 B.n222 B.n221 163.367
R273 B.n223 B.n222 163.367
R274 B.n223 B.n70 163.367
R275 B.n227 B.n70 163.367
R276 B.n228 B.n227 163.367
R277 B.n229 B.n228 163.367
R278 B.n295 B.n294 163.367
R279 B.n294 B.n293 163.367
R280 B.n293 B.n48 163.367
R281 B.n289 B.n48 163.367
R282 B.n289 B.n288 163.367
R283 B.n288 B.n287 163.367
R284 B.n287 B.n50 163.367
R285 B.n283 B.n50 163.367
R286 B.n283 B.n282 163.367
R287 B.n282 B.n281 163.367
R288 B.n281 B.n52 163.367
R289 B.n277 B.n52 163.367
R290 B.n277 B.n276 163.367
R291 B.n276 B.n275 163.367
R292 B.n275 B.n54 163.367
R293 B.n271 B.n54 163.367
R294 B.n271 B.n270 163.367
R295 B.n270 B.n269 163.367
R296 B.n269 B.n56 163.367
R297 B.n265 B.n56 163.367
R298 B.n265 B.n264 163.367
R299 B.n264 B.n263 163.367
R300 B.n263 B.n58 163.367
R301 B.n259 B.n58 163.367
R302 B.n259 B.n258 163.367
R303 B.n258 B.n257 163.367
R304 B.n257 B.n60 163.367
R305 B.n253 B.n60 163.367
R306 B.n253 B.n252 163.367
R307 B.n252 B.n251 163.367
R308 B.n251 B.n62 163.367
R309 B.n247 B.n62 163.367
R310 B.n247 B.n246 163.367
R311 B.n246 B.n245 163.367
R312 B.n245 B.n64 163.367
R313 B.n241 B.n64 163.367
R314 B.n241 B.n240 163.367
R315 B.n240 B.n239 163.367
R316 B.n239 B.n66 163.367
R317 B.n235 B.n66 163.367
R318 B.n235 B.n234 163.367
R319 B.n234 B.n233 163.367
R320 B.n233 B.n68 163.367
R321 B.n384 B.n13 163.367
R322 B.n380 B.n13 163.367
R323 B.n380 B.n379 163.367
R324 B.n379 B.n378 163.367
R325 B.n378 B.n15 163.367
R326 B.n374 B.n15 163.367
R327 B.n374 B.n373 163.367
R328 B.n373 B.n372 163.367
R329 B.n372 B.n17 163.367
R330 B.n368 B.n17 163.367
R331 B.n368 B.n367 163.367
R332 B.n367 B.n366 163.367
R333 B.n366 B.n19 163.367
R334 B.n362 B.n19 163.367
R335 B.n362 B.n361 163.367
R336 B.n361 B.n360 163.367
R337 B.n360 B.n21 163.367
R338 B.n356 B.n21 163.367
R339 B.n356 B.n355 163.367
R340 B.n355 B.n354 163.367
R341 B.n354 B.n23 163.367
R342 B.n350 B.n23 163.367
R343 B.n350 B.n349 163.367
R344 B.n349 B.n348 163.367
R345 B.n348 B.n25 163.367
R346 B.n344 B.n25 163.367
R347 B.n344 B.n343 163.367
R348 B.n343 B.n342 163.367
R349 B.n342 B.n30 163.367
R350 B.n338 B.n30 163.367
R351 B.n338 B.n337 163.367
R352 B.n337 B.n336 163.367
R353 B.n336 B.n32 163.367
R354 B.n331 B.n32 163.367
R355 B.n331 B.n330 163.367
R356 B.n330 B.n329 163.367
R357 B.n329 B.n36 163.367
R358 B.n325 B.n36 163.367
R359 B.n325 B.n324 163.367
R360 B.n324 B.n323 163.367
R361 B.n323 B.n38 163.367
R362 B.n319 B.n38 163.367
R363 B.n319 B.n318 163.367
R364 B.n318 B.n317 163.367
R365 B.n317 B.n40 163.367
R366 B.n313 B.n40 163.367
R367 B.n313 B.n312 163.367
R368 B.n312 B.n311 163.367
R369 B.n311 B.n42 163.367
R370 B.n307 B.n42 163.367
R371 B.n307 B.n306 163.367
R372 B.n306 B.n305 163.367
R373 B.n305 B.n44 163.367
R374 B.n301 B.n44 163.367
R375 B.n301 B.n300 163.367
R376 B.n300 B.n299 163.367
R377 B.n299 B.n46 163.367
R378 B.n386 B.n385 163.367
R379 B.n386 B.n11 163.367
R380 B.n390 B.n11 163.367
R381 B.n391 B.n390 163.367
R382 B.n392 B.n391 163.367
R383 B.n392 B.n9 163.367
R384 B.n396 B.n9 163.367
R385 B.n397 B.n396 163.367
R386 B.n398 B.n397 163.367
R387 B.n398 B.n7 163.367
R388 B.n402 B.n7 163.367
R389 B.n403 B.n402 163.367
R390 B.n404 B.n403 163.367
R391 B.n404 B.n5 163.367
R392 B.n408 B.n5 163.367
R393 B.n409 B.n408 163.367
R394 B.n410 B.n409 163.367
R395 B.n410 B.n3 163.367
R396 B.n414 B.n3 163.367
R397 B.n415 B.n414 163.367
R398 B.n110 B.n2 163.367
R399 B.n111 B.n110 163.367
R400 B.n111 B.n108 163.367
R401 B.n115 B.n108 163.367
R402 B.n116 B.n115 163.367
R403 B.n117 B.n116 163.367
R404 B.n117 B.n106 163.367
R405 B.n121 B.n106 163.367
R406 B.n122 B.n121 163.367
R407 B.n123 B.n122 163.367
R408 B.n123 B.n104 163.367
R409 B.n127 B.n104 163.367
R410 B.n128 B.n127 163.367
R411 B.n129 B.n128 163.367
R412 B.n129 B.n102 163.367
R413 B.n133 B.n102 163.367
R414 B.n134 B.n133 163.367
R415 B.n135 B.n134 163.367
R416 B.n135 B.n100 163.367
R417 B.n139 B.n100 163.367
R418 B.n176 B.n175 59.5399
R419 B.n194 B.n82 59.5399
R420 B.n333 B.n34 59.5399
R421 B.n28 B.n27 59.5399
R422 B.n175 B.n174 44.0247
R423 B.n82 B.n81 44.0247
R424 B.n34 B.n33 44.0247
R425 B.n27 B.n26 44.0247
R426 B.n383 B.n12 31.0639
R427 B.n297 B.n296 31.0639
R428 B.n231 B.n230 31.0639
R429 B.n138 B.n99 31.0639
R430 B B.n417 18.0485
R431 B.n387 B.n12 10.6151
R432 B.n388 B.n387 10.6151
R433 B.n389 B.n388 10.6151
R434 B.n389 B.n10 10.6151
R435 B.n393 B.n10 10.6151
R436 B.n394 B.n393 10.6151
R437 B.n395 B.n394 10.6151
R438 B.n395 B.n8 10.6151
R439 B.n399 B.n8 10.6151
R440 B.n400 B.n399 10.6151
R441 B.n401 B.n400 10.6151
R442 B.n401 B.n6 10.6151
R443 B.n405 B.n6 10.6151
R444 B.n406 B.n405 10.6151
R445 B.n407 B.n406 10.6151
R446 B.n407 B.n4 10.6151
R447 B.n411 B.n4 10.6151
R448 B.n412 B.n411 10.6151
R449 B.n413 B.n412 10.6151
R450 B.n413 B.n0 10.6151
R451 B.n383 B.n382 10.6151
R452 B.n382 B.n381 10.6151
R453 B.n381 B.n14 10.6151
R454 B.n377 B.n14 10.6151
R455 B.n377 B.n376 10.6151
R456 B.n376 B.n375 10.6151
R457 B.n375 B.n16 10.6151
R458 B.n371 B.n16 10.6151
R459 B.n371 B.n370 10.6151
R460 B.n370 B.n369 10.6151
R461 B.n369 B.n18 10.6151
R462 B.n365 B.n18 10.6151
R463 B.n365 B.n364 10.6151
R464 B.n364 B.n363 10.6151
R465 B.n363 B.n20 10.6151
R466 B.n359 B.n20 10.6151
R467 B.n359 B.n358 10.6151
R468 B.n358 B.n357 10.6151
R469 B.n357 B.n22 10.6151
R470 B.n353 B.n22 10.6151
R471 B.n353 B.n352 10.6151
R472 B.n352 B.n351 10.6151
R473 B.n351 B.n24 10.6151
R474 B.n347 B.n346 10.6151
R475 B.n346 B.n345 10.6151
R476 B.n345 B.n29 10.6151
R477 B.n341 B.n29 10.6151
R478 B.n341 B.n340 10.6151
R479 B.n340 B.n339 10.6151
R480 B.n339 B.n31 10.6151
R481 B.n335 B.n31 10.6151
R482 B.n335 B.n334 10.6151
R483 B.n332 B.n35 10.6151
R484 B.n328 B.n35 10.6151
R485 B.n328 B.n327 10.6151
R486 B.n327 B.n326 10.6151
R487 B.n326 B.n37 10.6151
R488 B.n322 B.n37 10.6151
R489 B.n322 B.n321 10.6151
R490 B.n321 B.n320 10.6151
R491 B.n320 B.n39 10.6151
R492 B.n316 B.n39 10.6151
R493 B.n316 B.n315 10.6151
R494 B.n315 B.n314 10.6151
R495 B.n314 B.n41 10.6151
R496 B.n310 B.n41 10.6151
R497 B.n310 B.n309 10.6151
R498 B.n309 B.n308 10.6151
R499 B.n308 B.n43 10.6151
R500 B.n304 B.n43 10.6151
R501 B.n304 B.n303 10.6151
R502 B.n303 B.n302 10.6151
R503 B.n302 B.n45 10.6151
R504 B.n298 B.n45 10.6151
R505 B.n298 B.n297 10.6151
R506 B.n296 B.n47 10.6151
R507 B.n292 B.n47 10.6151
R508 B.n292 B.n291 10.6151
R509 B.n291 B.n290 10.6151
R510 B.n290 B.n49 10.6151
R511 B.n286 B.n49 10.6151
R512 B.n286 B.n285 10.6151
R513 B.n285 B.n284 10.6151
R514 B.n284 B.n51 10.6151
R515 B.n280 B.n51 10.6151
R516 B.n280 B.n279 10.6151
R517 B.n279 B.n278 10.6151
R518 B.n278 B.n53 10.6151
R519 B.n274 B.n53 10.6151
R520 B.n274 B.n273 10.6151
R521 B.n273 B.n272 10.6151
R522 B.n272 B.n55 10.6151
R523 B.n268 B.n55 10.6151
R524 B.n268 B.n267 10.6151
R525 B.n267 B.n266 10.6151
R526 B.n266 B.n57 10.6151
R527 B.n262 B.n57 10.6151
R528 B.n262 B.n261 10.6151
R529 B.n261 B.n260 10.6151
R530 B.n260 B.n59 10.6151
R531 B.n256 B.n59 10.6151
R532 B.n256 B.n255 10.6151
R533 B.n255 B.n254 10.6151
R534 B.n254 B.n61 10.6151
R535 B.n250 B.n61 10.6151
R536 B.n250 B.n249 10.6151
R537 B.n249 B.n248 10.6151
R538 B.n248 B.n63 10.6151
R539 B.n244 B.n63 10.6151
R540 B.n244 B.n243 10.6151
R541 B.n243 B.n242 10.6151
R542 B.n242 B.n65 10.6151
R543 B.n238 B.n65 10.6151
R544 B.n238 B.n237 10.6151
R545 B.n237 B.n236 10.6151
R546 B.n236 B.n67 10.6151
R547 B.n232 B.n67 10.6151
R548 B.n232 B.n231 10.6151
R549 B.n109 B.n1 10.6151
R550 B.n112 B.n109 10.6151
R551 B.n113 B.n112 10.6151
R552 B.n114 B.n113 10.6151
R553 B.n114 B.n107 10.6151
R554 B.n118 B.n107 10.6151
R555 B.n119 B.n118 10.6151
R556 B.n120 B.n119 10.6151
R557 B.n120 B.n105 10.6151
R558 B.n124 B.n105 10.6151
R559 B.n125 B.n124 10.6151
R560 B.n126 B.n125 10.6151
R561 B.n126 B.n103 10.6151
R562 B.n130 B.n103 10.6151
R563 B.n131 B.n130 10.6151
R564 B.n132 B.n131 10.6151
R565 B.n132 B.n101 10.6151
R566 B.n136 B.n101 10.6151
R567 B.n137 B.n136 10.6151
R568 B.n138 B.n137 10.6151
R569 B.n142 B.n99 10.6151
R570 B.n143 B.n142 10.6151
R571 B.n144 B.n143 10.6151
R572 B.n144 B.n97 10.6151
R573 B.n148 B.n97 10.6151
R574 B.n149 B.n148 10.6151
R575 B.n150 B.n149 10.6151
R576 B.n150 B.n95 10.6151
R577 B.n154 B.n95 10.6151
R578 B.n155 B.n154 10.6151
R579 B.n156 B.n155 10.6151
R580 B.n156 B.n93 10.6151
R581 B.n160 B.n93 10.6151
R582 B.n161 B.n160 10.6151
R583 B.n162 B.n161 10.6151
R584 B.n162 B.n91 10.6151
R585 B.n166 B.n91 10.6151
R586 B.n167 B.n166 10.6151
R587 B.n168 B.n167 10.6151
R588 B.n168 B.n89 10.6151
R589 B.n172 B.n89 10.6151
R590 B.n173 B.n172 10.6151
R591 B.n177 B.n173 10.6151
R592 B.n181 B.n87 10.6151
R593 B.n182 B.n181 10.6151
R594 B.n183 B.n182 10.6151
R595 B.n183 B.n85 10.6151
R596 B.n187 B.n85 10.6151
R597 B.n188 B.n187 10.6151
R598 B.n189 B.n188 10.6151
R599 B.n189 B.n83 10.6151
R600 B.n193 B.n83 10.6151
R601 B.n196 B.n195 10.6151
R602 B.n196 B.n79 10.6151
R603 B.n200 B.n79 10.6151
R604 B.n201 B.n200 10.6151
R605 B.n202 B.n201 10.6151
R606 B.n202 B.n77 10.6151
R607 B.n206 B.n77 10.6151
R608 B.n207 B.n206 10.6151
R609 B.n208 B.n207 10.6151
R610 B.n208 B.n75 10.6151
R611 B.n212 B.n75 10.6151
R612 B.n213 B.n212 10.6151
R613 B.n214 B.n213 10.6151
R614 B.n214 B.n73 10.6151
R615 B.n218 B.n73 10.6151
R616 B.n219 B.n218 10.6151
R617 B.n220 B.n219 10.6151
R618 B.n220 B.n71 10.6151
R619 B.n224 B.n71 10.6151
R620 B.n225 B.n224 10.6151
R621 B.n226 B.n225 10.6151
R622 B.n226 B.n69 10.6151
R623 B.n230 B.n69 10.6151
R624 B.n28 B.n24 9.36635
R625 B.n333 B.n332 9.36635
R626 B.n177 B.n176 9.36635
R627 B.n195 B.n194 9.36635
R628 B.n417 B.n0 8.11757
R629 B.n417 B.n1 8.11757
R630 B.n347 B.n28 1.24928
R631 B.n334 B.n333 1.24928
R632 B.n176 B.n87 1.24928
R633 B.n194 B.n193 1.24928
R634 VP.n0 VP.t0 172.417
R635 VP.n0 VP.t1 134.018
R636 VP VP.n0 0.241678
R637 VTAIL.n122 VTAIL.n96 756.745
R638 VTAIL.n26 VTAIL.n0 756.745
R639 VTAIL.n90 VTAIL.n64 756.745
R640 VTAIL.n58 VTAIL.n32 756.745
R641 VTAIL.n107 VTAIL.n106 585
R642 VTAIL.n104 VTAIL.n103 585
R643 VTAIL.n113 VTAIL.n112 585
R644 VTAIL.n115 VTAIL.n114 585
R645 VTAIL.n100 VTAIL.n99 585
R646 VTAIL.n121 VTAIL.n120 585
R647 VTAIL.n123 VTAIL.n122 585
R648 VTAIL.n11 VTAIL.n10 585
R649 VTAIL.n8 VTAIL.n7 585
R650 VTAIL.n17 VTAIL.n16 585
R651 VTAIL.n19 VTAIL.n18 585
R652 VTAIL.n4 VTAIL.n3 585
R653 VTAIL.n25 VTAIL.n24 585
R654 VTAIL.n27 VTAIL.n26 585
R655 VTAIL.n91 VTAIL.n90 585
R656 VTAIL.n89 VTAIL.n88 585
R657 VTAIL.n68 VTAIL.n67 585
R658 VTAIL.n83 VTAIL.n82 585
R659 VTAIL.n81 VTAIL.n80 585
R660 VTAIL.n72 VTAIL.n71 585
R661 VTAIL.n75 VTAIL.n74 585
R662 VTAIL.n59 VTAIL.n58 585
R663 VTAIL.n57 VTAIL.n56 585
R664 VTAIL.n36 VTAIL.n35 585
R665 VTAIL.n51 VTAIL.n50 585
R666 VTAIL.n49 VTAIL.n48 585
R667 VTAIL.n40 VTAIL.n39 585
R668 VTAIL.n43 VTAIL.n42 585
R669 VTAIL.t0 VTAIL.n105 327.601
R670 VTAIL.t2 VTAIL.n9 327.601
R671 VTAIL.t3 VTAIL.n73 327.601
R672 VTAIL.t1 VTAIL.n41 327.601
R673 VTAIL.n106 VTAIL.n103 171.744
R674 VTAIL.n113 VTAIL.n103 171.744
R675 VTAIL.n114 VTAIL.n113 171.744
R676 VTAIL.n114 VTAIL.n99 171.744
R677 VTAIL.n121 VTAIL.n99 171.744
R678 VTAIL.n122 VTAIL.n121 171.744
R679 VTAIL.n10 VTAIL.n7 171.744
R680 VTAIL.n17 VTAIL.n7 171.744
R681 VTAIL.n18 VTAIL.n17 171.744
R682 VTAIL.n18 VTAIL.n3 171.744
R683 VTAIL.n25 VTAIL.n3 171.744
R684 VTAIL.n26 VTAIL.n25 171.744
R685 VTAIL.n90 VTAIL.n89 171.744
R686 VTAIL.n89 VTAIL.n67 171.744
R687 VTAIL.n82 VTAIL.n67 171.744
R688 VTAIL.n82 VTAIL.n81 171.744
R689 VTAIL.n81 VTAIL.n71 171.744
R690 VTAIL.n74 VTAIL.n71 171.744
R691 VTAIL.n58 VTAIL.n57 171.744
R692 VTAIL.n57 VTAIL.n35 171.744
R693 VTAIL.n50 VTAIL.n35 171.744
R694 VTAIL.n50 VTAIL.n49 171.744
R695 VTAIL.n49 VTAIL.n39 171.744
R696 VTAIL.n42 VTAIL.n39 171.744
R697 VTAIL.n106 VTAIL.t0 85.8723
R698 VTAIL.n10 VTAIL.t2 85.8723
R699 VTAIL.n74 VTAIL.t3 85.8723
R700 VTAIL.n42 VTAIL.t1 85.8723
R701 VTAIL.n127 VTAIL.n126 33.155
R702 VTAIL.n31 VTAIL.n30 33.155
R703 VTAIL.n95 VTAIL.n94 33.155
R704 VTAIL.n63 VTAIL.n62 33.155
R705 VTAIL.n63 VTAIL.n31 21.4962
R706 VTAIL.n127 VTAIL.n95 19.5393
R707 VTAIL.n107 VTAIL.n105 16.3865
R708 VTAIL.n11 VTAIL.n9 16.3865
R709 VTAIL.n75 VTAIL.n73 16.3865
R710 VTAIL.n43 VTAIL.n41 16.3865
R711 VTAIL.n108 VTAIL.n104 12.8005
R712 VTAIL.n12 VTAIL.n8 12.8005
R713 VTAIL.n76 VTAIL.n72 12.8005
R714 VTAIL.n44 VTAIL.n40 12.8005
R715 VTAIL.n112 VTAIL.n111 12.0247
R716 VTAIL.n16 VTAIL.n15 12.0247
R717 VTAIL.n80 VTAIL.n79 12.0247
R718 VTAIL.n48 VTAIL.n47 12.0247
R719 VTAIL.n115 VTAIL.n102 11.249
R720 VTAIL.n19 VTAIL.n6 11.249
R721 VTAIL.n83 VTAIL.n70 11.249
R722 VTAIL.n51 VTAIL.n38 11.249
R723 VTAIL.n116 VTAIL.n100 10.4732
R724 VTAIL.n20 VTAIL.n4 10.4732
R725 VTAIL.n84 VTAIL.n68 10.4732
R726 VTAIL.n52 VTAIL.n36 10.4732
R727 VTAIL.n120 VTAIL.n119 9.69747
R728 VTAIL.n24 VTAIL.n23 9.69747
R729 VTAIL.n88 VTAIL.n87 9.69747
R730 VTAIL.n56 VTAIL.n55 9.69747
R731 VTAIL.n126 VTAIL.n125 9.45567
R732 VTAIL.n30 VTAIL.n29 9.45567
R733 VTAIL.n94 VTAIL.n93 9.45567
R734 VTAIL.n62 VTAIL.n61 9.45567
R735 VTAIL.n125 VTAIL.n124 9.3005
R736 VTAIL.n98 VTAIL.n97 9.3005
R737 VTAIL.n119 VTAIL.n118 9.3005
R738 VTAIL.n117 VTAIL.n116 9.3005
R739 VTAIL.n102 VTAIL.n101 9.3005
R740 VTAIL.n111 VTAIL.n110 9.3005
R741 VTAIL.n109 VTAIL.n108 9.3005
R742 VTAIL.n29 VTAIL.n28 9.3005
R743 VTAIL.n2 VTAIL.n1 9.3005
R744 VTAIL.n23 VTAIL.n22 9.3005
R745 VTAIL.n21 VTAIL.n20 9.3005
R746 VTAIL.n6 VTAIL.n5 9.3005
R747 VTAIL.n15 VTAIL.n14 9.3005
R748 VTAIL.n13 VTAIL.n12 9.3005
R749 VTAIL.n93 VTAIL.n92 9.3005
R750 VTAIL.n66 VTAIL.n65 9.3005
R751 VTAIL.n87 VTAIL.n86 9.3005
R752 VTAIL.n85 VTAIL.n84 9.3005
R753 VTAIL.n70 VTAIL.n69 9.3005
R754 VTAIL.n79 VTAIL.n78 9.3005
R755 VTAIL.n77 VTAIL.n76 9.3005
R756 VTAIL.n61 VTAIL.n60 9.3005
R757 VTAIL.n34 VTAIL.n33 9.3005
R758 VTAIL.n55 VTAIL.n54 9.3005
R759 VTAIL.n53 VTAIL.n52 9.3005
R760 VTAIL.n38 VTAIL.n37 9.3005
R761 VTAIL.n47 VTAIL.n46 9.3005
R762 VTAIL.n45 VTAIL.n44 9.3005
R763 VTAIL.n123 VTAIL.n98 8.92171
R764 VTAIL.n27 VTAIL.n2 8.92171
R765 VTAIL.n91 VTAIL.n66 8.92171
R766 VTAIL.n59 VTAIL.n34 8.92171
R767 VTAIL.n124 VTAIL.n96 8.14595
R768 VTAIL.n28 VTAIL.n0 8.14595
R769 VTAIL.n92 VTAIL.n64 8.14595
R770 VTAIL.n60 VTAIL.n32 8.14595
R771 VTAIL.n126 VTAIL.n96 5.81868
R772 VTAIL.n30 VTAIL.n0 5.81868
R773 VTAIL.n94 VTAIL.n64 5.81868
R774 VTAIL.n62 VTAIL.n32 5.81868
R775 VTAIL.n124 VTAIL.n123 5.04292
R776 VTAIL.n28 VTAIL.n27 5.04292
R777 VTAIL.n92 VTAIL.n91 5.04292
R778 VTAIL.n60 VTAIL.n59 5.04292
R779 VTAIL.n120 VTAIL.n98 4.26717
R780 VTAIL.n24 VTAIL.n2 4.26717
R781 VTAIL.n88 VTAIL.n66 4.26717
R782 VTAIL.n56 VTAIL.n34 4.26717
R783 VTAIL.n77 VTAIL.n73 3.71286
R784 VTAIL.n45 VTAIL.n41 3.71286
R785 VTAIL.n109 VTAIL.n105 3.71286
R786 VTAIL.n13 VTAIL.n9 3.71286
R787 VTAIL.n119 VTAIL.n100 3.49141
R788 VTAIL.n23 VTAIL.n4 3.49141
R789 VTAIL.n87 VTAIL.n68 3.49141
R790 VTAIL.n55 VTAIL.n36 3.49141
R791 VTAIL.n116 VTAIL.n115 2.71565
R792 VTAIL.n20 VTAIL.n19 2.71565
R793 VTAIL.n84 VTAIL.n83 2.71565
R794 VTAIL.n52 VTAIL.n51 2.71565
R795 VTAIL.n112 VTAIL.n102 1.93989
R796 VTAIL.n16 VTAIL.n6 1.93989
R797 VTAIL.n80 VTAIL.n70 1.93989
R798 VTAIL.n48 VTAIL.n38 1.93989
R799 VTAIL.n95 VTAIL.n63 1.44878
R800 VTAIL.n111 VTAIL.n104 1.16414
R801 VTAIL.n15 VTAIL.n8 1.16414
R802 VTAIL.n79 VTAIL.n72 1.16414
R803 VTAIL.n47 VTAIL.n40 1.16414
R804 VTAIL VTAIL.n31 1.01774
R805 VTAIL VTAIL.n127 0.431534
R806 VTAIL.n108 VTAIL.n107 0.388379
R807 VTAIL.n12 VTAIL.n11 0.388379
R808 VTAIL.n76 VTAIL.n75 0.388379
R809 VTAIL.n44 VTAIL.n43 0.388379
R810 VTAIL.n110 VTAIL.n109 0.155672
R811 VTAIL.n110 VTAIL.n101 0.155672
R812 VTAIL.n117 VTAIL.n101 0.155672
R813 VTAIL.n118 VTAIL.n117 0.155672
R814 VTAIL.n118 VTAIL.n97 0.155672
R815 VTAIL.n125 VTAIL.n97 0.155672
R816 VTAIL.n14 VTAIL.n13 0.155672
R817 VTAIL.n14 VTAIL.n5 0.155672
R818 VTAIL.n21 VTAIL.n5 0.155672
R819 VTAIL.n22 VTAIL.n21 0.155672
R820 VTAIL.n22 VTAIL.n1 0.155672
R821 VTAIL.n29 VTAIL.n1 0.155672
R822 VTAIL.n93 VTAIL.n65 0.155672
R823 VTAIL.n86 VTAIL.n65 0.155672
R824 VTAIL.n86 VTAIL.n85 0.155672
R825 VTAIL.n85 VTAIL.n69 0.155672
R826 VTAIL.n78 VTAIL.n69 0.155672
R827 VTAIL.n78 VTAIL.n77 0.155672
R828 VTAIL.n61 VTAIL.n33 0.155672
R829 VTAIL.n54 VTAIL.n33 0.155672
R830 VTAIL.n54 VTAIL.n53 0.155672
R831 VTAIL.n53 VTAIL.n37 0.155672
R832 VTAIL.n46 VTAIL.n37 0.155672
R833 VTAIL.n46 VTAIL.n45 0.155672
R834 VDD1.n26 VDD1.n0 756.745
R835 VDD1.n57 VDD1.n31 756.745
R836 VDD1.n27 VDD1.n26 585
R837 VDD1.n25 VDD1.n24 585
R838 VDD1.n4 VDD1.n3 585
R839 VDD1.n19 VDD1.n18 585
R840 VDD1.n17 VDD1.n16 585
R841 VDD1.n8 VDD1.n7 585
R842 VDD1.n11 VDD1.n10 585
R843 VDD1.n42 VDD1.n41 585
R844 VDD1.n39 VDD1.n38 585
R845 VDD1.n48 VDD1.n47 585
R846 VDD1.n50 VDD1.n49 585
R847 VDD1.n35 VDD1.n34 585
R848 VDD1.n56 VDD1.n55 585
R849 VDD1.n58 VDD1.n57 585
R850 VDD1.t1 VDD1.n9 327.601
R851 VDD1.t0 VDD1.n40 327.601
R852 VDD1.n26 VDD1.n25 171.744
R853 VDD1.n25 VDD1.n3 171.744
R854 VDD1.n18 VDD1.n3 171.744
R855 VDD1.n18 VDD1.n17 171.744
R856 VDD1.n17 VDD1.n7 171.744
R857 VDD1.n10 VDD1.n7 171.744
R858 VDD1.n41 VDD1.n38 171.744
R859 VDD1.n48 VDD1.n38 171.744
R860 VDD1.n49 VDD1.n48 171.744
R861 VDD1.n49 VDD1.n34 171.744
R862 VDD1.n56 VDD1.n34 171.744
R863 VDD1.n57 VDD1.n56 171.744
R864 VDD1.n10 VDD1.t1 85.8723
R865 VDD1.n41 VDD1.t0 85.8723
R866 VDD1 VDD1.n61 83.6366
R867 VDD1 VDD1.n30 50.3812
R868 VDD1.n11 VDD1.n9 16.3865
R869 VDD1.n42 VDD1.n40 16.3865
R870 VDD1.n12 VDD1.n8 12.8005
R871 VDD1.n43 VDD1.n39 12.8005
R872 VDD1.n16 VDD1.n15 12.0247
R873 VDD1.n47 VDD1.n46 12.0247
R874 VDD1.n19 VDD1.n6 11.249
R875 VDD1.n50 VDD1.n37 11.249
R876 VDD1.n20 VDD1.n4 10.4732
R877 VDD1.n51 VDD1.n35 10.4732
R878 VDD1.n24 VDD1.n23 9.69747
R879 VDD1.n55 VDD1.n54 9.69747
R880 VDD1.n30 VDD1.n29 9.45567
R881 VDD1.n61 VDD1.n60 9.45567
R882 VDD1.n29 VDD1.n28 9.3005
R883 VDD1.n2 VDD1.n1 9.3005
R884 VDD1.n23 VDD1.n22 9.3005
R885 VDD1.n21 VDD1.n20 9.3005
R886 VDD1.n6 VDD1.n5 9.3005
R887 VDD1.n15 VDD1.n14 9.3005
R888 VDD1.n13 VDD1.n12 9.3005
R889 VDD1.n60 VDD1.n59 9.3005
R890 VDD1.n33 VDD1.n32 9.3005
R891 VDD1.n54 VDD1.n53 9.3005
R892 VDD1.n52 VDD1.n51 9.3005
R893 VDD1.n37 VDD1.n36 9.3005
R894 VDD1.n46 VDD1.n45 9.3005
R895 VDD1.n44 VDD1.n43 9.3005
R896 VDD1.n27 VDD1.n2 8.92171
R897 VDD1.n58 VDD1.n33 8.92171
R898 VDD1.n28 VDD1.n0 8.14595
R899 VDD1.n59 VDD1.n31 8.14595
R900 VDD1.n30 VDD1.n0 5.81868
R901 VDD1.n61 VDD1.n31 5.81868
R902 VDD1.n28 VDD1.n27 5.04292
R903 VDD1.n59 VDD1.n58 5.04292
R904 VDD1.n24 VDD1.n2 4.26717
R905 VDD1.n55 VDD1.n33 4.26717
R906 VDD1.n13 VDD1.n9 3.71286
R907 VDD1.n44 VDD1.n40 3.71286
R908 VDD1.n23 VDD1.n4 3.49141
R909 VDD1.n54 VDD1.n35 3.49141
R910 VDD1.n20 VDD1.n19 2.71565
R911 VDD1.n51 VDD1.n50 2.71565
R912 VDD1.n16 VDD1.n6 1.93989
R913 VDD1.n47 VDD1.n37 1.93989
R914 VDD1.n15 VDD1.n8 1.16414
R915 VDD1.n46 VDD1.n39 1.16414
R916 VDD1.n12 VDD1.n11 0.388379
R917 VDD1.n43 VDD1.n42 0.388379
R918 VDD1.n29 VDD1.n1 0.155672
R919 VDD1.n22 VDD1.n1 0.155672
R920 VDD1.n22 VDD1.n21 0.155672
R921 VDD1.n21 VDD1.n5 0.155672
R922 VDD1.n14 VDD1.n5 0.155672
R923 VDD1.n14 VDD1.n13 0.155672
R924 VDD1.n45 VDD1.n44 0.155672
R925 VDD1.n45 VDD1.n36 0.155672
R926 VDD1.n52 VDD1.n36 0.155672
R927 VDD1.n53 VDD1.n52 0.155672
R928 VDD1.n53 VDD1.n32 0.155672
R929 VDD1.n60 VDD1.n32 0.155672
R930 VN VN.t0 172.608
R931 VN VN.t1 134.26
R932 VDD2.n57 VDD2.n31 756.745
R933 VDD2.n26 VDD2.n0 756.745
R934 VDD2.n58 VDD2.n57 585
R935 VDD2.n56 VDD2.n55 585
R936 VDD2.n35 VDD2.n34 585
R937 VDD2.n50 VDD2.n49 585
R938 VDD2.n48 VDD2.n47 585
R939 VDD2.n39 VDD2.n38 585
R940 VDD2.n42 VDD2.n41 585
R941 VDD2.n11 VDD2.n10 585
R942 VDD2.n8 VDD2.n7 585
R943 VDD2.n17 VDD2.n16 585
R944 VDD2.n19 VDD2.n18 585
R945 VDD2.n4 VDD2.n3 585
R946 VDD2.n25 VDD2.n24 585
R947 VDD2.n27 VDD2.n26 585
R948 VDD2.t1 VDD2.n40 327.601
R949 VDD2.t0 VDD2.n9 327.601
R950 VDD2.n57 VDD2.n56 171.744
R951 VDD2.n56 VDD2.n34 171.744
R952 VDD2.n49 VDD2.n34 171.744
R953 VDD2.n49 VDD2.n48 171.744
R954 VDD2.n48 VDD2.n38 171.744
R955 VDD2.n41 VDD2.n38 171.744
R956 VDD2.n10 VDD2.n7 171.744
R957 VDD2.n17 VDD2.n7 171.744
R958 VDD2.n18 VDD2.n17 171.744
R959 VDD2.n18 VDD2.n3 171.744
R960 VDD2.n25 VDD2.n3 171.744
R961 VDD2.n26 VDD2.n25 171.744
R962 VDD2.n41 VDD2.t1 85.8723
R963 VDD2.n10 VDD2.t0 85.8723
R964 VDD2.n62 VDD2.n30 82.6226
R965 VDD2.n62 VDD2.n61 49.8338
R966 VDD2.n42 VDD2.n40 16.3865
R967 VDD2.n11 VDD2.n9 16.3865
R968 VDD2.n43 VDD2.n39 12.8005
R969 VDD2.n12 VDD2.n8 12.8005
R970 VDD2.n47 VDD2.n46 12.0247
R971 VDD2.n16 VDD2.n15 12.0247
R972 VDD2.n50 VDD2.n37 11.249
R973 VDD2.n19 VDD2.n6 11.249
R974 VDD2.n51 VDD2.n35 10.4732
R975 VDD2.n20 VDD2.n4 10.4732
R976 VDD2.n55 VDD2.n54 9.69747
R977 VDD2.n24 VDD2.n23 9.69747
R978 VDD2.n61 VDD2.n60 9.45567
R979 VDD2.n30 VDD2.n29 9.45567
R980 VDD2.n60 VDD2.n59 9.3005
R981 VDD2.n33 VDD2.n32 9.3005
R982 VDD2.n54 VDD2.n53 9.3005
R983 VDD2.n52 VDD2.n51 9.3005
R984 VDD2.n37 VDD2.n36 9.3005
R985 VDD2.n46 VDD2.n45 9.3005
R986 VDD2.n44 VDD2.n43 9.3005
R987 VDD2.n29 VDD2.n28 9.3005
R988 VDD2.n2 VDD2.n1 9.3005
R989 VDD2.n23 VDD2.n22 9.3005
R990 VDD2.n21 VDD2.n20 9.3005
R991 VDD2.n6 VDD2.n5 9.3005
R992 VDD2.n15 VDD2.n14 9.3005
R993 VDD2.n13 VDD2.n12 9.3005
R994 VDD2.n58 VDD2.n33 8.92171
R995 VDD2.n27 VDD2.n2 8.92171
R996 VDD2.n59 VDD2.n31 8.14595
R997 VDD2.n28 VDD2.n0 8.14595
R998 VDD2.n61 VDD2.n31 5.81868
R999 VDD2.n30 VDD2.n0 5.81868
R1000 VDD2.n59 VDD2.n58 5.04292
R1001 VDD2.n28 VDD2.n27 5.04292
R1002 VDD2.n55 VDD2.n33 4.26717
R1003 VDD2.n24 VDD2.n2 4.26717
R1004 VDD2.n44 VDD2.n40 3.71286
R1005 VDD2.n13 VDD2.n9 3.71286
R1006 VDD2.n54 VDD2.n35 3.49141
R1007 VDD2.n23 VDD2.n4 3.49141
R1008 VDD2.n51 VDD2.n50 2.71565
R1009 VDD2.n20 VDD2.n19 2.71565
R1010 VDD2.n47 VDD2.n37 1.93989
R1011 VDD2.n16 VDD2.n6 1.93989
R1012 VDD2.n46 VDD2.n39 1.16414
R1013 VDD2.n15 VDD2.n8 1.16414
R1014 VDD2 VDD2.n62 0.547914
R1015 VDD2.n43 VDD2.n42 0.388379
R1016 VDD2.n12 VDD2.n11 0.388379
R1017 VDD2.n60 VDD2.n32 0.155672
R1018 VDD2.n53 VDD2.n32 0.155672
R1019 VDD2.n53 VDD2.n52 0.155672
R1020 VDD2.n52 VDD2.n36 0.155672
R1021 VDD2.n45 VDD2.n36 0.155672
R1022 VDD2.n45 VDD2.n44 0.155672
R1023 VDD2.n14 VDD2.n13 0.155672
R1024 VDD2.n14 VDD2.n5 0.155672
R1025 VDD2.n21 VDD2.n5 0.155672
R1026 VDD2.n22 VDD2.n21 0.155672
R1027 VDD2.n22 VDD2.n1 0.155672
R1028 VDD2.n29 VDD2.n1 0.155672
C0 VN VTAIL 1.40499f
C1 B VTAIL 2.10219f
C2 VP w_n1878_n2178# 2.6598f
C3 VDD2 VTAIL 3.40136f
C4 VP VTAIL 1.41922f
C5 VDD1 VN 0.147819f
C6 VDD1 B 1.15288f
C7 VTAIL w_n1878_n2178# 1.89991f
C8 VDD1 VDD2 0.595475f
C9 B VN 0.865085f
C10 VN VDD2 1.45677f
C11 B VDD2 1.17713f
C12 VDD1 VP 1.61211f
C13 VP VN 4.042861f
C14 VP B 1.25339f
C15 VP VDD2 0.304815f
C16 VDD1 w_n1878_n2178# 1.28759f
C17 VN w_n1878_n2178# 2.42201f
C18 B w_n1878_n2178# 6.43561f
C19 VDD2 w_n1878_n2178# 1.30555f
C20 VDD1 VTAIL 3.35424f
C21 VDD2 VSUBS 0.613595f
C22 VDD1 VSUBS 2.187787f
C23 VTAIL VSUBS 0.506332f
C24 VN VSUBS 5.02136f
C25 VP VSUBS 1.175499f
C26 B VSUBS 2.901157f
C27 w_n1878_n2178# VSUBS 51.044003f
C28 VDD2.n0 VSUBS 0.016254f
C29 VDD2.n1 VSUBS 0.014567f
C30 VDD2.n2 VSUBS 0.007828f
C31 VDD2.n3 VSUBS 0.018502f
C32 VDD2.n4 VSUBS 0.008288f
C33 VDD2.n5 VSUBS 0.014567f
C34 VDD2.n6 VSUBS 0.007828f
C35 VDD2.n7 VSUBS 0.018502f
C36 VDD2.n8 VSUBS 0.008288f
C37 VDD2.n9 VSUBS 0.064662f
C38 VDD2.t0 VSUBS 0.039741f
C39 VDD2.n10 VSUBS 0.013876f
C40 VDD2.n11 VSUBS 0.011764f
C41 VDD2.n12 VSUBS 0.007828f
C42 VDD2.n13 VSUBS 0.337387f
C43 VDD2.n14 VSUBS 0.014567f
C44 VDD2.n15 VSUBS 0.007828f
C45 VDD2.n16 VSUBS 0.008288f
C46 VDD2.n17 VSUBS 0.018502f
C47 VDD2.n18 VSUBS 0.018502f
C48 VDD2.n19 VSUBS 0.008288f
C49 VDD2.n20 VSUBS 0.007828f
C50 VDD2.n21 VSUBS 0.014567f
C51 VDD2.n22 VSUBS 0.014567f
C52 VDD2.n23 VSUBS 0.007828f
C53 VDD2.n24 VSUBS 0.008288f
C54 VDD2.n25 VSUBS 0.018502f
C55 VDD2.n26 VSUBS 0.045635f
C56 VDD2.n27 VSUBS 0.008288f
C57 VDD2.n28 VSUBS 0.007828f
C58 VDD2.n29 VSUBS 0.034666f
C59 VDD2.n30 VSUBS 0.288179f
C60 VDD2.n31 VSUBS 0.016254f
C61 VDD2.n32 VSUBS 0.014567f
C62 VDD2.n33 VSUBS 0.007828f
C63 VDD2.n34 VSUBS 0.018502f
C64 VDD2.n35 VSUBS 0.008288f
C65 VDD2.n36 VSUBS 0.014567f
C66 VDD2.n37 VSUBS 0.007828f
C67 VDD2.n38 VSUBS 0.018502f
C68 VDD2.n39 VSUBS 0.008288f
C69 VDD2.n40 VSUBS 0.064662f
C70 VDD2.t1 VSUBS 0.039741f
C71 VDD2.n41 VSUBS 0.013876f
C72 VDD2.n42 VSUBS 0.011764f
C73 VDD2.n43 VSUBS 0.007828f
C74 VDD2.n44 VSUBS 0.337387f
C75 VDD2.n45 VSUBS 0.014567f
C76 VDD2.n46 VSUBS 0.007828f
C77 VDD2.n47 VSUBS 0.008288f
C78 VDD2.n48 VSUBS 0.018502f
C79 VDD2.n49 VSUBS 0.018502f
C80 VDD2.n50 VSUBS 0.008288f
C81 VDD2.n51 VSUBS 0.007828f
C82 VDD2.n52 VSUBS 0.014567f
C83 VDD2.n53 VSUBS 0.014567f
C84 VDD2.n54 VSUBS 0.007828f
C85 VDD2.n55 VSUBS 0.008288f
C86 VDD2.n56 VSUBS 0.018502f
C87 VDD2.n57 VSUBS 0.045635f
C88 VDD2.n58 VSUBS 0.008288f
C89 VDD2.n59 VSUBS 0.007828f
C90 VDD2.n60 VSUBS 0.034666f
C91 VDD2.n61 VSUBS 0.033068f
C92 VDD2.n62 VSUBS 1.33902f
C93 VN.t1 VSUBS 1.41881f
C94 VN.t0 VSUBS 1.81073f
C95 VDD1.n0 VSUBS 0.016001f
C96 VDD1.n1 VSUBS 0.01434f
C97 VDD1.n2 VSUBS 0.007706f
C98 VDD1.n3 VSUBS 0.018214f
C99 VDD1.n4 VSUBS 0.008159f
C100 VDD1.n5 VSUBS 0.01434f
C101 VDD1.n6 VSUBS 0.007706f
C102 VDD1.n7 VSUBS 0.018214f
C103 VDD1.n8 VSUBS 0.008159f
C104 VDD1.n9 VSUBS 0.063655f
C105 VDD1.t1 VSUBS 0.039122f
C106 VDD1.n10 VSUBS 0.01366f
C107 VDD1.n11 VSUBS 0.01158f
C108 VDD1.n12 VSUBS 0.007706f
C109 VDD1.n13 VSUBS 0.332131f
C110 VDD1.n14 VSUBS 0.01434f
C111 VDD1.n15 VSUBS 0.007706f
C112 VDD1.n16 VSUBS 0.008159f
C113 VDD1.n17 VSUBS 0.018214f
C114 VDD1.n18 VSUBS 0.018214f
C115 VDD1.n19 VSUBS 0.008159f
C116 VDD1.n20 VSUBS 0.007706f
C117 VDD1.n21 VSUBS 0.01434f
C118 VDD1.n22 VSUBS 0.01434f
C119 VDD1.n23 VSUBS 0.007706f
C120 VDD1.n24 VSUBS 0.008159f
C121 VDD1.n25 VSUBS 0.018214f
C122 VDD1.n26 VSUBS 0.044924f
C123 VDD1.n27 VSUBS 0.008159f
C124 VDD1.n28 VSUBS 0.007706f
C125 VDD1.n29 VSUBS 0.034126f
C126 VDD1.n30 VSUBS 0.033134f
C127 VDD1.n31 VSUBS 0.016001f
C128 VDD1.n32 VSUBS 0.01434f
C129 VDD1.n33 VSUBS 0.007706f
C130 VDD1.n34 VSUBS 0.018214f
C131 VDD1.n35 VSUBS 0.008159f
C132 VDD1.n36 VSUBS 0.01434f
C133 VDD1.n37 VSUBS 0.007706f
C134 VDD1.n38 VSUBS 0.018214f
C135 VDD1.n39 VSUBS 0.008159f
C136 VDD1.n40 VSUBS 0.063655f
C137 VDD1.t0 VSUBS 0.039122f
C138 VDD1.n41 VSUBS 0.01366f
C139 VDD1.n42 VSUBS 0.01158f
C140 VDD1.n43 VSUBS 0.007706f
C141 VDD1.n44 VSUBS 0.332131f
C142 VDD1.n45 VSUBS 0.01434f
C143 VDD1.n46 VSUBS 0.007706f
C144 VDD1.n47 VSUBS 0.008159f
C145 VDD1.n48 VSUBS 0.018214f
C146 VDD1.n49 VSUBS 0.018214f
C147 VDD1.n50 VSUBS 0.008159f
C148 VDD1.n51 VSUBS 0.007706f
C149 VDD1.n52 VSUBS 0.01434f
C150 VDD1.n53 VSUBS 0.01434f
C151 VDD1.n54 VSUBS 0.007706f
C152 VDD1.n55 VSUBS 0.008159f
C153 VDD1.n56 VSUBS 0.018214f
C154 VDD1.n57 VSUBS 0.044924f
C155 VDD1.n58 VSUBS 0.008159f
C156 VDD1.n59 VSUBS 0.007706f
C157 VDD1.n60 VSUBS 0.034126f
C158 VDD1.n61 VSUBS 0.305496f
C159 VTAIL.n0 VSUBS 0.023819f
C160 VTAIL.n1 VSUBS 0.021347f
C161 VTAIL.n2 VSUBS 0.011471f
C162 VTAIL.n3 VSUBS 0.027113f
C163 VTAIL.n4 VSUBS 0.012146f
C164 VTAIL.n5 VSUBS 0.021347f
C165 VTAIL.n6 VSUBS 0.011471f
C166 VTAIL.n7 VSUBS 0.027113f
C167 VTAIL.n8 VSUBS 0.012146f
C168 VTAIL.n9 VSUBS 0.094759f
C169 VTAIL.t2 VSUBS 0.058238f
C170 VTAIL.n10 VSUBS 0.020335f
C171 VTAIL.n11 VSUBS 0.017239f
C172 VTAIL.n12 VSUBS 0.011471f
C173 VTAIL.n13 VSUBS 0.494419f
C174 VTAIL.n14 VSUBS 0.021347f
C175 VTAIL.n15 VSUBS 0.011471f
C176 VTAIL.n16 VSUBS 0.012146f
C177 VTAIL.n17 VSUBS 0.027113f
C178 VTAIL.n18 VSUBS 0.027113f
C179 VTAIL.n19 VSUBS 0.012146f
C180 VTAIL.n20 VSUBS 0.011471f
C181 VTAIL.n21 VSUBS 0.021347f
C182 VTAIL.n22 VSUBS 0.021347f
C183 VTAIL.n23 VSUBS 0.011471f
C184 VTAIL.n24 VSUBS 0.012146f
C185 VTAIL.n25 VSUBS 0.027113f
C186 VTAIL.n26 VSUBS 0.066876f
C187 VTAIL.n27 VSUBS 0.012146f
C188 VTAIL.n28 VSUBS 0.011471f
C189 VTAIL.n29 VSUBS 0.050801f
C190 VTAIL.n30 VSUBS 0.03373f
C191 VTAIL.n31 VSUBS 1.00696f
C192 VTAIL.n32 VSUBS 0.023819f
C193 VTAIL.n33 VSUBS 0.021347f
C194 VTAIL.n34 VSUBS 0.011471f
C195 VTAIL.n35 VSUBS 0.027113f
C196 VTAIL.n36 VSUBS 0.012146f
C197 VTAIL.n37 VSUBS 0.021347f
C198 VTAIL.n38 VSUBS 0.011471f
C199 VTAIL.n39 VSUBS 0.027113f
C200 VTAIL.n40 VSUBS 0.012146f
C201 VTAIL.n41 VSUBS 0.094759f
C202 VTAIL.t1 VSUBS 0.058238f
C203 VTAIL.n42 VSUBS 0.020335f
C204 VTAIL.n43 VSUBS 0.017239f
C205 VTAIL.n44 VSUBS 0.011471f
C206 VTAIL.n45 VSUBS 0.494419f
C207 VTAIL.n46 VSUBS 0.021347f
C208 VTAIL.n47 VSUBS 0.011471f
C209 VTAIL.n48 VSUBS 0.012146f
C210 VTAIL.n49 VSUBS 0.027113f
C211 VTAIL.n50 VSUBS 0.027113f
C212 VTAIL.n51 VSUBS 0.012146f
C213 VTAIL.n52 VSUBS 0.011471f
C214 VTAIL.n53 VSUBS 0.021347f
C215 VTAIL.n54 VSUBS 0.021347f
C216 VTAIL.n55 VSUBS 0.011471f
C217 VTAIL.n56 VSUBS 0.012146f
C218 VTAIL.n57 VSUBS 0.027113f
C219 VTAIL.n58 VSUBS 0.066876f
C220 VTAIL.n59 VSUBS 0.012146f
C221 VTAIL.n60 VSUBS 0.011471f
C222 VTAIL.n61 VSUBS 0.050801f
C223 VTAIL.n62 VSUBS 0.03373f
C224 VTAIL.n63 VSUBS 1.03661f
C225 VTAIL.n64 VSUBS 0.023819f
C226 VTAIL.n65 VSUBS 0.021347f
C227 VTAIL.n66 VSUBS 0.011471f
C228 VTAIL.n67 VSUBS 0.027113f
C229 VTAIL.n68 VSUBS 0.012146f
C230 VTAIL.n69 VSUBS 0.021347f
C231 VTAIL.n70 VSUBS 0.011471f
C232 VTAIL.n71 VSUBS 0.027113f
C233 VTAIL.n72 VSUBS 0.012146f
C234 VTAIL.n73 VSUBS 0.094759f
C235 VTAIL.t3 VSUBS 0.058238f
C236 VTAIL.n74 VSUBS 0.020335f
C237 VTAIL.n75 VSUBS 0.017239f
C238 VTAIL.n76 VSUBS 0.011471f
C239 VTAIL.n77 VSUBS 0.494419f
C240 VTAIL.n78 VSUBS 0.021347f
C241 VTAIL.n79 VSUBS 0.011471f
C242 VTAIL.n80 VSUBS 0.012146f
C243 VTAIL.n81 VSUBS 0.027113f
C244 VTAIL.n82 VSUBS 0.027113f
C245 VTAIL.n83 VSUBS 0.012146f
C246 VTAIL.n84 VSUBS 0.011471f
C247 VTAIL.n85 VSUBS 0.021347f
C248 VTAIL.n86 VSUBS 0.021347f
C249 VTAIL.n87 VSUBS 0.011471f
C250 VTAIL.n88 VSUBS 0.012146f
C251 VTAIL.n89 VSUBS 0.027113f
C252 VTAIL.n90 VSUBS 0.066876f
C253 VTAIL.n91 VSUBS 0.012146f
C254 VTAIL.n92 VSUBS 0.011471f
C255 VTAIL.n93 VSUBS 0.050801f
C256 VTAIL.n94 VSUBS 0.03373f
C257 VTAIL.n95 VSUBS 0.902007f
C258 VTAIL.n96 VSUBS 0.023819f
C259 VTAIL.n97 VSUBS 0.021347f
C260 VTAIL.n98 VSUBS 0.011471f
C261 VTAIL.n99 VSUBS 0.027113f
C262 VTAIL.n100 VSUBS 0.012146f
C263 VTAIL.n101 VSUBS 0.021347f
C264 VTAIL.n102 VSUBS 0.011471f
C265 VTAIL.n103 VSUBS 0.027113f
C266 VTAIL.n104 VSUBS 0.012146f
C267 VTAIL.n105 VSUBS 0.094759f
C268 VTAIL.t0 VSUBS 0.058238f
C269 VTAIL.n106 VSUBS 0.020335f
C270 VTAIL.n107 VSUBS 0.017239f
C271 VTAIL.n108 VSUBS 0.011471f
C272 VTAIL.n109 VSUBS 0.494419f
C273 VTAIL.n110 VSUBS 0.021347f
C274 VTAIL.n111 VSUBS 0.011471f
C275 VTAIL.n112 VSUBS 0.012146f
C276 VTAIL.n113 VSUBS 0.027113f
C277 VTAIL.n114 VSUBS 0.027113f
C278 VTAIL.n115 VSUBS 0.012146f
C279 VTAIL.n116 VSUBS 0.011471f
C280 VTAIL.n117 VSUBS 0.021347f
C281 VTAIL.n118 VSUBS 0.021347f
C282 VTAIL.n119 VSUBS 0.011471f
C283 VTAIL.n120 VSUBS 0.012146f
C284 VTAIL.n121 VSUBS 0.027113f
C285 VTAIL.n122 VSUBS 0.066876f
C286 VTAIL.n123 VSUBS 0.012146f
C287 VTAIL.n124 VSUBS 0.011471f
C288 VTAIL.n125 VSUBS 0.050801f
C289 VTAIL.n126 VSUBS 0.03373f
C290 VTAIL.n127 VSUBS 0.832036f
C291 VP.t0 VSUBS 1.90527f
C292 VP.t1 VSUBS 1.49649f
C293 VP.n0 VSUBS 3.23509f
C294 B.n0 VSUBS 0.00706f
C295 B.n1 VSUBS 0.00706f
C296 B.n2 VSUBS 0.010442f
C297 B.n3 VSUBS 0.008002f
C298 B.n4 VSUBS 0.008002f
C299 B.n5 VSUBS 0.008002f
C300 B.n6 VSUBS 0.008002f
C301 B.n7 VSUBS 0.008002f
C302 B.n8 VSUBS 0.008002f
C303 B.n9 VSUBS 0.008002f
C304 B.n10 VSUBS 0.008002f
C305 B.n11 VSUBS 0.008002f
C306 B.n12 VSUBS 0.017601f
C307 B.n13 VSUBS 0.008002f
C308 B.n14 VSUBS 0.008002f
C309 B.n15 VSUBS 0.008002f
C310 B.n16 VSUBS 0.008002f
C311 B.n17 VSUBS 0.008002f
C312 B.n18 VSUBS 0.008002f
C313 B.n19 VSUBS 0.008002f
C314 B.n20 VSUBS 0.008002f
C315 B.n21 VSUBS 0.008002f
C316 B.n22 VSUBS 0.008002f
C317 B.n23 VSUBS 0.008002f
C318 B.n24 VSUBS 0.007531f
C319 B.n25 VSUBS 0.008002f
C320 B.t4 VSUBS 0.103426f
C321 B.t5 VSUBS 0.126652f
C322 B.t3 VSUBS 0.624423f
C323 B.n26 VSUBS 0.21906f
C324 B.n27 VSUBS 0.176642f
C325 B.n28 VSUBS 0.018539f
C326 B.n29 VSUBS 0.008002f
C327 B.n30 VSUBS 0.008002f
C328 B.n31 VSUBS 0.008002f
C329 B.n32 VSUBS 0.008002f
C330 B.t7 VSUBS 0.103428f
C331 B.t8 VSUBS 0.126654f
C332 B.t6 VSUBS 0.624423f
C333 B.n33 VSUBS 0.219058f
C334 B.n34 VSUBS 0.17664f
C335 B.n35 VSUBS 0.008002f
C336 B.n36 VSUBS 0.008002f
C337 B.n37 VSUBS 0.008002f
C338 B.n38 VSUBS 0.008002f
C339 B.n39 VSUBS 0.008002f
C340 B.n40 VSUBS 0.008002f
C341 B.n41 VSUBS 0.008002f
C342 B.n42 VSUBS 0.008002f
C343 B.n43 VSUBS 0.008002f
C344 B.n44 VSUBS 0.008002f
C345 B.n45 VSUBS 0.008002f
C346 B.n46 VSUBS 0.018643f
C347 B.n47 VSUBS 0.008002f
C348 B.n48 VSUBS 0.008002f
C349 B.n49 VSUBS 0.008002f
C350 B.n50 VSUBS 0.008002f
C351 B.n51 VSUBS 0.008002f
C352 B.n52 VSUBS 0.008002f
C353 B.n53 VSUBS 0.008002f
C354 B.n54 VSUBS 0.008002f
C355 B.n55 VSUBS 0.008002f
C356 B.n56 VSUBS 0.008002f
C357 B.n57 VSUBS 0.008002f
C358 B.n58 VSUBS 0.008002f
C359 B.n59 VSUBS 0.008002f
C360 B.n60 VSUBS 0.008002f
C361 B.n61 VSUBS 0.008002f
C362 B.n62 VSUBS 0.008002f
C363 B.n63 VSUBS 0.008002f
C364 B.n64 VSUBS 0.008002f
C365 B.n65 VSUBS 0.008002f
C366 B.n66 VSUBS 0.008002f
C367 B.n67 VSUBS 0.008002f
C368 B.n68 VSUBS 0.017601f
C369 B.n69 VSUBS 0.008002f
C370 B.n70 VSUBS 0.008002f
C371 B.n71 VSUBS 0.008002f
C372 B.n72 VSUBS 0.008002f
C373 B.n73 VSUBS 0.008002f
C374 B.n74 VSUBS 0.008002f
C375 B.n75 VSUBS 0.008002f
C376 B.n76 VSUBS 0.008002f
C377 B.n77 VSUBS 0.008002f
C378 B.n78 VSUBS 0.008002f
C379 B.n79 VSUBS 0.008002f
C380 B.n80 VSUBS 0.008002f
C381 B.t11 VSUBS 0.103428f
C382 B.t10 VSUBS 0.126654f
C383 B.t9 VSUBS 0.624423f
C384 B.n81 VSUBS 0.219058f
C385 B.n82 VSUBS 0.17664f
C386 B.n83 VSUBS 0.008002f
C387 B.n84 VSUBS 0.008002f
C388 B.n85 VSUBS 0.008002f
C389 B.n86 VSUBS 0.008002f
C390 B.n87 VSUBS 0.004472f
C391 B.n88 VSUBS 0.008002f
C392 B.n89 VSUBS 0.008002f
C393 B.n90 VSUBS 0.008002f
C394 B.n91 VSUBS 0.008002f
C395 B.n92 VSUBS 0.008002f
C396 B.n93 VSUBS 0.008002f
C397 B.n94 VSUBS 0.008002f
C398 B.n95 VSUBS 0.008002f
C399 B.n96 VSUBS 0.008002f
C400 B.n97 VSUBS 0.008002f
C401 B.n98 VSUBS 0.008002f
C402 B.n99 VSUBS 0.018643f
C403 B.n100 VSUBS 0.008002f
C404 B.n101 VSUBS 0.008002f
C405 B.n102 VSUBS 0.008002f
C406 B.n103 VSUBS 0.008002f
C407 B.n104 VSUBS 0.008002f
C408 B.n105 VSUBS 0.008002f
C409 B.n106 VSUBS 0.008002f
C410 B.n107 VSUBS 0.008002f
C411 B.n108 VSUBS 0.008002f
C412 B.n109 VSUBS 0.008002f
C413 B.n110 VSUBS 0.008002f
C414 B.n111 VSUBS 0.008002f
C415 B.n112 VSUBS 0.008002f
C416 B.n113 VSUBS 0.008002f
C417 B.n114 VSUBS 0.008002f
C418 B.n115 VSUBS 0.008002f
C419 B.n116 VSUBS 0.008002f
C420 B.n117 VSUBS 0.008002f
C421 B.n118 VSUBS 0.008002f
C422 B.n119 VSUBS 0.008002f
C423 B.n120 VSUBS 0.008002f
C424 B.n121 VSUBS 0.008002f
C425 B.n122 VSUBS 0.008002f
C426 B.n123 VSUBS 0.008002f
C427 B.n124 VSUBS 0.008002f
C428 B.n125 VSUBS 0.008002f
C429 B.n126 VSUBS 0.008002f
C430 B.n127 VSUBS 0.008002f
C431 B.n128 VSUBS 0.008002f
C432 B.n129 VSUBS 0.008002f
C433 B.n130 VSUBS 0.008002f
C434 B.n131 VSUBS 0.008002f
C435 B.n132 VSUBS 0.008002f
C436 B.n133 VSUBS 0.008002f
C437 B.n134 VSUBS 0.008002f
C438 B.n135 VSUBS 0.008002f
C439 B.n136 VSUBS 0.008002f
C440 B.n137 VSUBS 0.008002f
C441 B.n138 VSUBS 0.017601f
C442 B.n139 VSUBS 0.017601f
C443 B.n140 VSUBS 0.018643f
C444 B.n141 VSUBS 0.008002f
C445 B.n142 VSUBS 0.008002f
C446 B.n143 VSUBS 0.008002f
C447 B.n144 VSUBS 0.008002f
C448 B.n145 VSUBS 0.008002f
C449 B.n146 VSUBS 0.008002f
C450 B.n147 VSUBS 0.008002f
C451 B.n148 VSUBS 0.008002f
C452 B.n149 VSUBS 0.008002f
C453 B.n150 VSUBS 0.008002f
C454 B.n151 VSUBS 0.008002f
C455 B.n152 VSUBS 0.008002f
C456 B.n153 VSUBS 0.008002f
C457 B.n154 VSUBS 0.008002f
C458 B.n155 VSUBS 0.008002f
C459 B.n156 VSUBS 0.008002f
C460 B.n157 VSUBS 0.008002f
C461 B.n158 VSUBS 0.008002f
C462 B.n159 VSUBS 0.008002f
C463 B.n160 VSUBS 0.008002f
C464 B.n161 VSUBS 0.008002f
C465 B.n162 VSUBS 0.008002f
C466 B.n163 VSUBS 0.008002f
C467 B.n164 VSUBS 0.008002f
C468 B.n165 VSUBS 0.008002f
C469 B.n166 VSUBS 0.008002f
C470 B.n167 VSUBS 0.008002f
C471 B.n168 VSUBS 0.008002f
C472 B.n169 VSUBS 0.008002f
C473 B.n170 VSUBS 0.008002f
C474 B.n171 VSUBS 0.008002f
C475 B.n172 VSUBS 0.008002f
C476 B.n173 VSUBS 0.008002f
C477 B.t2 VSUBS 0.103426f
C478 B.t1 VSUBS 0.126652f
C479 B.t0 VSUBS 0.624423f
C480 B.n174 VSUBS 0.21906f
C481 B.n175 VSUBS 0.176642f
C482 B.n176 VSUBS 0.018539f
C483 B.n177 VSUBS 0.007531f
C484 B.n178 VSUBS 0.008002f
C485 B.n179 VSUBS 0.008002f
C486 B.n180 VSUBS 0.008002f
C487 B.n181 VSUBS 0.008002f
C488 B.n182 VSUBS 0.008002f
C489 B.n183 VSUBS 0.008002f
C490 B.n184 VSUBS 0.008002f
C491 B.n185 VSUBS 0.008002f
C492 B.n186 VSUBS 0.008002f
C493 B.n187 VSUBS 0.008002f
C494 B.n188 VSUBS 0.008002f
C495 B.n189 VSUBS 0.008002f
C496 B.n190 VSUBS 0.008002f
C497 B.n191 VSUBS 0.008002f
C498 B.n192 VSUBS 0.008002f
C499 B.n193 VSUBS 0.004472f
C500 B.n194 VSUBS 0.018539f
C501 B.n195 VSUBS 0.007531f
C502 B.n196 VSUBS 0.008002f
C503 B.n197 VSUBS 0.008002f
C504 B.n198 VSUBS 0.008002f
C505 B.n199 VSUBS 0.008002f
C506 B.n200 VSUBS 0.008002f
C507 B.n201 VSUBS 0.008002f
C508 B.n202 VSUBS 0.008002f
C509 B.n203 VSUBS 0.008002f
C510 B.n204 VSUBS 0.008002f
C511 B.n205 VSUBS 0.008002f
C512 B.n206 VSUBS 0.008002f
C513 B.n207 VSUBS 0.008002f
C514 B.n208 VSUBS 0.008002f
C515 B.n209 VSUBS 0.008002f
C516 B.n210 VSUBS 0.008002f
C517 B.n211 VSUBS 0.008002f
C518 B.n212 VSUBS 0.008002f
C519 B.n213 VSUBS 0.008002f
C520 B.n214 VSUBS 0.008002f
C521 B.n215 VSUBS 0.008002f
C522 B.n216 VSUBS 0.008002f
C523 B.n217 VSUBS 0.008002f
C524 B.n218 VSUBS 0.008002f
C525 B.n219 VSUBS 0.008002f
C526 B.n220 VSUBS 0.008002f
C527 B.n221 VSUBS 0.008002f
C528 B.n222 VSUBS 0.008002f
C529 B.n223 VSUBS 0.008002f
C530 B.n224 VSUBS 0.008002f
C531 B.n225 VSUBS 0.008002f
C532 B.n226 VSUBS 0.008002f
C533 B.n227 VSUBS 0.008002f
C534 B.n228 VSUBS 0.008002f
C535 B.n229 VSUBS 0.018643f
C536 B.n230 VSUBS 0.017649f
C537 B.n231 VSUBS 0.018595f
C538 B.n232 VSUBS 0.008002f
C539 B.n233 VSUBS 0.008002f
C540 B.n234 VSUBS 0.008002f
C541 B.n235 VSUBS 0.008002f
C542 B.n236 VSUBS 0.008002f
C543 B.n237 VSUBS 0.008002f
C544 B.n238 VSUBS 0.008002f
C545 B.n239 VSUBS 0.008002f
C546 B.n240 VSUBS 0.008002f
C547 B.n241 VSUBS 0.008002f
C548 B.n242 VSUBS 0.008002f
C549 B.n243 VSUBS 0.008002f
C550 B.n244 VSUBS 0.008002f
C551 B.n245 VSUBS 0.008002f
C552 B.n246 VSUBS 0.008002f
C553 B.n247 VSUBS 0.008002f
C554 B.n248 VSUBS 0.008002f
C555 B.n249 VSUBS 0.008002f
C556 B.n250 VSUBS 0.008002f
C557 B.n251 VSUBS 0.008002f
C558 B.n252 VSUBS 0.008002f
C559 B.n253 VSUBS 0.008002f
C560 B.n254 VSUBS 0.008002f
C561 B.n255 VSUBS 0.008002f
C562 B.n256 VSUBS 0.008002f
C563 B.n257 VSUBS 0.008002f
C564 B.n258 VSUBS 0.008002f
C565 B.n259 VSUBS 0.008002f
C566 B.n260 VSUBS 0.008002f
C567 B.n261 VSUBS 0.008002f
C568 B.n262 VSUBS 0.008002f
C569 B.n263 VSUBS 0.008002f
C570 B.n264 VSUBS 0.008002f
C571 B.n265 VSUBS 0.008002f
C572 B.n266 VSUBS 0.008002f
C573 B.n267 VSUBS 0.008002f
C574 B.n268 VSUBS 0.008002f
C575 B.n269 VSUBS 0.008002f
C576 B.n270 VSUBS 0.008002f
C577 B.n271 VSUBS 0.008002f
C578 B.n272 VSUBS 0.008002f
C579 B.n273 VSUBS 0.008002f
C580 B.n274 VSUBS 0.008002f
C581 B.n275 VSUBS 0.008002f
C582 B.n276 VSUBS 0.008002f
C583 B.n277 VSUBS 0.008002f
C584 B.n278 VSUBS 0.008002f
C585 B.n279 VSUBS 0.008002f
C586 B.n280 VSUBS 0.008002f
C587 B.n281 VSUBS 0.008002f
C588 B.n282 VSUBS 0.008002f
C589 B.n283 VSUBS 0.008002f
C590 B.n284 VSUBS 0.008002f
C591 B.n285 VSUBS 0.008002f
C592 B.n286 VSUBS 0.008002f
C593 B.n287 VSUBS 0.008002f
C594 B.n288 VSUBS 0.008002f
C595 B.n289 VSUBS 0.008002f
C596 B.n290 VSUBS 0.008002f
C597 B.n291 VSUBS 0.008002f
C598 B.n292 VSUBS 0.008002f
C599 B.n293 VSUBS 0.008002f
C600 B.n294 VSUBS 0.008002f
C601 B.n295 VSUBS 0.017601f
C602 B.n296 VSUBS 0.017601f
C603 B.n297 VSUBS 0.018643f
C604 B.n298 VSUBS 0.008002f
C605 B.n299 VSUBS 0.008002f
C606 B.n300 VSUBS 0.008002f
C607 B.n301 VSUBS 0.008002f
C608 B.n302 VSUBS 0.008002f
C609 B.n303 VSUBS 0.008002f
C610 B.n304 VSUBS 0.008002f
C611 B.n305 VSUBS 0.008002f
C612 B.n306 VSUBS 0.008002f
C613 B.n307 VSUBS 0.008002f
C614 B.n308 VSUBS 0.008002f
C615 B.n309 VSUBS 0.008002f
C616 B.n310 VSUBS 0.008002f
C617 B.n311 VSUBS 0.008002f
C618 B.n312 VSUBS 0.008002f
C619 B.n313 VSUBS 0.008002f
C620 B.n314 VSUBS 0.008002f
C621 B.n315 VSUBS 0.008002f
C622 B.n316 VSUBS 0.008002f
C623 B.n317 VSUBS 0.008002f
C624 B.n318 VSUBS 0.008002f
C625 B.n319 VSUBS 0.008002f
C626 B.n320 VSUBS 0.008002f
C627 B.n321 VSUBS 0.008002f
C628 B.n322 VSUBS 0.008002f
C629 B.n323 VSUBS 0.008002f
C630 B.n324 VSUBS 0.008002f
C631 B.n325 VSUBS 0.008002f
C632 B.n326 VSUBS 0.008002f
C633 B.n327 VSUBS 0.008002f
C634 B.n328 VSUBS 0.008002f
C635 B.n329 VSUBS 0.008002f
C636 B.n330 VSUBS 0.008002f
C637 B.n331 VSUBS 0.008002f
C638 B.n332 VSUBS 0.007531f
C639 B.n333 VSUBS 0.018539f
C640 B.n334 VSUBS 0.004472f
C641 B.n335 VSUBS 0.008002f
C642 B.n336 VSUBS 0.008002f
C643 B.n337 VSUBS 0.008002f
C644 B.n338 VSUBS 0.008002f
C645 B.n339 VSUBS 0.008002f
C646 B.n340 VSUBS 0.008002f
C647 B.n341 VSUBS 0.008002f
C648 B.n342 VSUBS 0.008002f
C649 B.n343 VSUBS 0.008002f
C650 B.n344 VSUBS 0.008002f
C651 B.n345 VSUBS 0.008002f
C652 B.n346 VSUBS 0.008002f
C653 B.n347 VSUBS 0.004472f
C654 B.n348 VSUBS 0.008002f
C655 B.n349 VSUBS 0.008002f
C656 B.n350 VSUBS 0.008002f
C657 B.n351 VSUBS 0.008002f
C658 B.n352 VSUBS 0.008002f
C659 B.n353 VSUBS 0.008002f
C660 B.n354 VSUBS 0.008002f
C661 B.n355 VSUBS 0.008002f
C662 B.n356 VSUBS 0.008002f
C663 B.n357 VSUBS 0.008002f
C664 B.n358 VSUBS 0.008002f
C665 B.n359 VSUBS 0.008002f
C666 B.n360 VSUBS 0.008002f
C667 B.n361 VSUBS 0.008002f
C668 B.n362 VSUBS 0.008002f
C669 B.n363 VSUBS 0.008002f
C670 B.n364 VSUBS 0.008002f
C671 B.n365 VSUBS 0.008002f
C672 B.n366 VSUBS 0.008002f
C673 B.n367 VSUBS 0.008002f
C674 B.n368 VSUBS 0.008002f
C675 B.n369 VSUBS 0.008002f
C676 B.n370 VSUBS 0.008002f
C677 B.n371 VSUBS 0.008002f
C678 B.n372 VSUBS 0.008002f
C679 B.n373 VSUBS 0.008002f
C680 B.n374 VSUBS 0.008002f
C681 B.n375 VSUBS 0.008002f
C682 B.n376 VSUBS 0.008002f
C683 B.n377 VSUBS 0.008002f
C684 B.n378 VSUBS 0.008002f
C685 B.n379 VSUBS 0.008002f
C686 B.n380 VSUBS 0.008002f
C687 B.n381 VSUBS 0.008002f
C688 B.n382 VSUBS 0.008002f
C689 B.n383 VSUBS 0.018643f
C690 B.n384 VSUBS 0.018643f
C691 B.n385 VSUBS 0.017601f
C692 B.n386 VSUBS 0.008002f
C693 B.n387 VSUBS 0.008002f
C694 B.n388 VSUBS 0.008002f
C695 B.n389 VSUBS 0.008002f
C696 B.n390 VSUBS 0.008002f
C697 B.n391 VSUBS 0.008002f
C698 B.n392 VSUBS 0.008002f
C699 B.n393 VSUBS 0.008002f
C700 B.n394 VSUBS 0.008002f
C701 B.n395 VSUBS 0.008002f
C702 B.n396 VSUBS 0.008002f
C703 B.n397 VSUBS 0.008002f
C704 B.n398 VSUBS 0.008002f
C705 B.n399 VSUBS 0.008002f
C706 B.n400 VSUBS 0.008002f
C707 B.n401 VSUBS 0.008002f
C708 B.n402 VSUBS 0.008002f
C709 B.n403 VSUBS 0.008002f
C710 B.n404 VSUBS 0.008002f
C711 B.n405 VSUBS 0.008002f
C712 B.n406 VSUBS 0.008002f
C713 B.n407 VSUBS 0.008002f
C714 B.n408 VSUBS 0.008002f
C715 B.n409 VSUBS 0.008002f
C716 B.n410 VSUBS 0.008002f
C717 B.n411 VSUBS 0.008002f
C718 B.n412 VSUBS 0.008002f
C719 B.n413 VSUBS 0.008002f
C720 B.n414 VSUBS 0.008002f
C721 B.n415 VSUBS 0.010442f
C722 B.n416 VSUBS 0.011123f
C723 B.n417 VSUBS 0.02212f
.ends

