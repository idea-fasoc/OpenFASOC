* NGSPICE file created from diff_pair_sample_0614.ext - technology: sky130A

.subckt diff_pair_sample_0614 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t5 VN.t0 VTAIL.t7 w_n2650_n2218# sky130_fd_pr__pfet_01v8 ad=2.4375 pd=13.28 as=1.03125 ps=6.58 w=6.25 l=1.77
X1 B.t11 B.t9 B.t10 w_n2650_n2218# sky130_fd_pr__pfet_01v8 ad=2.4375 pd=13.28 as=0 ps=0 w=6.25 l=1.77
X2 VDD2.t4 VN.t1 VTAIL.t5 w_n2650_n2218# sky130_fd_pr__pfet_01v8 ad=2.4375 pd=13.28 as=1.03125 ps=6.58 w=6.25 l=1.77
X3 B.t8 B.t6 B.t7 w_n2650_n2218# sky130_fd_pr__pfet_01v8 ad=2.4375 pd=13.28 as=0 ps=0 w=6.25 l=1.77
X4 VTAIL.t11 VP.t0 VDD1.t5 w_n2650_n2218# sky130_fd_pr__pfet_01v8 ad=1.03125 pd=6.58 as=1.03125 ps=6.58 w=6.25 l=1.77
X5 VDD2.t3 VN.t2 VTAIL.t6 w_n2650_n2218# sky130_fd_pr__pfet_01v8 ad=1.03125 pd=6.58 as=2.4375 ps=13.28 w=6.25 l=1.77
X6 B.t5 B.t3 B.t4 w_n2650_n2218# sky130_fd_pr__pfet_01v8 ad=2.4375 pd=13.28 as=0 ps=0 w=6.25 l=1.77
X7 VDD1.t4 VP.t1 VTAIL.t10 w_n2650_n2218# sky130_fd_pr__pfet_01v8 ad=1.03125 pd=6.58 as=2.4375 ps=13.28 w=6.25 l=1.77
X8 VDD1.t3 VP.t2 VTAIL.t3 w_n2650_n2218# sky130_fd_pr__pfet_01v8 ad=1.03125 pd=6.58 as=2.4375 ps=13.28 w=6.25 l=1.77
X9 VTAIL.t8 VN.t3 VDD2.t2 w_n2650_n2218# sky130_fd_pr__pfet_01v8 ad=1.03125 pd=6.58 as=1.03125 ps=6.58 w=6.25 l=1.77
X10 VTAIL.t1 VP.t3 VDD1.t2 w_n2650_n2218# sky130_fd_pr__pfet_01v8 ad=1.03125 pd=6.58 as=1.03125 ps=6.58 w=6.25 l=1.77
X11 VTAIL.t4 VN.t4 VDD2.t1 w_n2650_n2218# sky130_fd_pr__pfet_01v8 ad=1.03125 pd=6.58 as=1.03125 ps=6.58 w=6.25 l=1.77
X12 VDD2.t0 VN.t5 VTAIL.t9 w_n2650_n2218# sky130_fd_pr__pfet_01v8 ad=1.03125 pd=6.58 as=2.4375 ps=13.28 w=6.25 l=1.77
X13 VDD1.t1 VP.t4 VTAIL.t0 w_n2650_n2218# sky130_fd_pr__pfet_01v8 ad=2.4375 pd=13.28 as=1.03125 ps=6.58 w=6.25 l=1.77
X14 B.t2 B.t0 B.t1 w_n2650_n2218# sky130_fd_pr__pfet_01v8 ad=2.4375 pd=13.28 as=0 ps=0 w=6.25 l=1.77
X15 VDD1.t0 VP.t5 VTAIL.t2 w_n2650_n2218# sky130_fd_pr__pfet_01v8 ad=2.4375 pd=13.28 as=1.03125 ps=6.58 w=6.25 l=1.77
R0 VN.n11 VN.n10 180.875
R1 VN.n23 VN.n22 180.875
R2 VN.n21 VN.n12 161.3
R3 VN.n20 VN.n19 161.3
R4 VN.n18 VN.n13 161.3
R5 VN.n17 VN.n16 161.3
R6 VN.n9 VN.n0 161.3
R7 VN.n8 VN.n7 161.3
R8 VN.n6 VN.n1 161.3
R9 VN.n5 VN.n4 161.3
R10 VN.n2 VN.t1 120.436
R11 VN.n14 VN.t2 120.436
R12 VN.n3 VN.t3 85.0994
R13 VN.n10 VN.t5 85.0994
R14 VN.n15 VN.t4 85.0994
R15 VN.n22 VN.t0 85.0994
R16 VN.n8 VN.n1 45.3497
R17 VN.n20 VN.n13 45.3497
R18 VN.n15 VN.n14 44.5155
R19 VN.n3 VN.n2 44.5155
R20 VN VN.n23 41.3585
R21 VN.n4 VN.n1 35.6371
R22 VN.n16 VN.n13 35.6371
R23 VN.n4 VN.n3 24.4675
R24 VN.n9 VN.n8 24.4675
R25 VN.n16 VN.n15 24.4675
R26 VN.n21 VN.n20 24.4675
R27 VN.n17 VN.n14 12.2033
R28 VN.n5 VN.n2 12.2033
R29 VN.n10 VN.n9 4.8939
R30 VN.n22 VN.n21 4.8939
R31 VN.n23 VN.n12 0.189894
R32 VN.n19 VN.n12 0.189894
R33 VN.n19 VN.n18 0.189894
R34 VN.n18 VN.n17 0.189894
R35 VN.n6 VN.n5 0.189894
R36 VN.n7 VN.n6 0.189894
R37 VN.n7 VN.n0 0.189894
R38 VN.n11 VN.n0 0.189894
R39 VN VN.n11 0.0516364
R40 VTAIL.n7 VTAIL.t6 76.6171
R41 VTAIL.n11 VTAIL.t9 76.617
R42 VTAIL.n2 VTAIL.t10 76.617
R43 VTAIL.n10 VTAIL.t3 76.617
R44 VTAIL.n9 VTAIL.n8 71.4163
R45 VTAIL.n6 VTAIL.n5 71.4163
R46 VTAIL.n1 VTAIL.n0 71.4161
R47 VTAIL.n4 VTAIL.n3 71.4161
R48 VTAIL.n6 VTAIL.n4 21.3755
R49 VTAIL.n11 VTAIL.n10 19.5652
R50 VTAIL.n0 VTAIL.t5 5.2013
R51 VTAIL.n0 VTAIL.t8 5.2013
R52 VTAIL.n3 VTAIL.t2 5.2013
R53 VTAIL.n3 VTAIL.t1 5.2013
R54 VTAIL.n8 VTAIL.t0 5.2013
R55 VTAIL.n8 VTAIL.t11 5.2013
R56 VTAIL.n5 VTAIL.t7 5.2013
R57 VTAIL.n5 VTAIL.t4 5.2013
R58 VTAIL.n7 VTAIL.n6 1.81084
R59 VTAIL.n10 VTAIL.n9 1.81084
R60 VTAIL.n4 VTAIL.n2 1.81084
R61 VTAIL.n9 VTAIL.n7 1.3755
R62 VTAIL.n2 VTAIL.n1 1.3755
R63 VTAIL VTAIL.n11 1.30007
R64 VTAIL VTAIL.n1 0.511276
R65 VDD2.n1 VDD2.t4 94.5982
R66 VDD2.n2 VDD2.t5 93.2959
R67 VDD2.n1 VDD2.n0 88.4921
R68 VDD2 VDD2.n3 88.4893
R69 VDD2.n2 VDD2.n1 34.9868
R70 VDD2.n3 VDD2.t1 5.2013
R71 VDD2.n3 VDD2.t3 5.2013
R72 VDD2.n0 VDD2.t2 5.2013
R73 VDD2.n0 VDD2.t0 5.2013
R74 VDD2 VDD2.n2 1.41645
R75 B.n375 B.n374 585
R76 B.n376 B.n51 585
R77 B.n378 B.n377 585
R78 B.n379 B.n50 585
R79 B.n381 B.n380 585
R80 B.n382 B.n49 585
R81 B.n384 B.n383 585
R82 B.n385 B.n48 585
R83 B.n387 B.n386 585
R84 B.n388 B.n47 585
R85 B.n390 B.n389 585
R86 B.n391 B.n46 585
R87 B.n393 B.n392 585
R88 B.n394 B.n45 585
R89 B.n396 B.n395 585
R90 B.n397 B.n44 585
R91 B.n399 B.n398 585
R92 B.n400 B.n43 585
R93 B.n402 B.n401 585
R94 B.n403 B.n42 585
R95 B.n405 B.n404 585
R96 B.n406 B.n41 585
R97 B.n408 B.n407 585
R98 B.n409 B.n40 585
R99 B.n411 B.n410 585
R100 B.n413 B.n37 585
R101 B.n415 B.n414 585
R102 B.n416 B.n36 585
R103 B.n418 B.n417 585
R104 B.n419 B.n35 585
R105 B.n421 B.n420 585
R106 B.n422 B.n34 585
R107 B.n424 B.n423 585
R108 B.n425 B.n31 585
R109 B.n428 B.n427 585
R110 B.n429 B.n30 585
R111 B.n431 B.n430 585
R112 B.n432 B.n29 585
R113 B.n434 B.n433 585
R114 B.n435 B.n28 585
R115 B.n437 B.n436 585
R116 B.n438 B.n27 585
R117 B.n440 B.n439 585
R118 B.n441 B.n26 585
R119 B.n443 B.n442 585
R120 B.n444 B.n25 585
R121 B.n446 B.n445 585
R122 B.n447 B.n24 585
R123 B.n449 B.n448 585
R124 B.n450 B.n23 585
R125 B.n452 B.n451 585
R126 B.n453 B.n22 585
R127 B.n455 B.n454 585
R128 B.n456 B.n21 585
R129 B.n458 B.n457 585
R130 B.n459 B.n20 585
R131 B.n461 B.n460 585
R132 B.n462 B.n19 585
R133 B.n464 B.n463 585
R134 B.n373 B.n52 585
R135 B.n372 B.n371 585
R136 B.n370 B.n53 585
R137 B.n369 B.n368 585
R138 B.n367 B.n54 585
R139 B.n366 B.n365 585
R140 B.n364 B.n55 585
R141 B.n363 B.n362 585
R142 B.n361 B.n56 585
R143 B.n360 B.n359 585
R144 B.n358 B.n57 585
R145 B.n357 B.n356 585
R146 B.n355 B.n58 585
R147 B.n354 B.n353 585
R148 B.n352 B.n59 585
R149 B.n351 B.n350 585
R150 B.n349 B.n60 585
R151 B.n348 B.n347 585
R152 B.n346 B.n61 585
R153 B.n345 B.n344 585
R154 B.n343 B.n62 585
R155 B.n342 B.n341 585
R156 B.n340 B.n63 585
R157 B.n339 B.n338 585
R158 B.n337 B.n64 585
R159 B.n336 B.n335 585
R160 B.n334 B.n65 585
R161 B.n333 B.n332 585
R162 B.n331 B.n66 585
R163 B.n330 B.n329 585
R164 B.n328 B.n67 585
R165 B.n327 B.n326 585
R166 B.n325 B.n68 585
R167 B.n324 B.n323 585
R168 B.n322 B.n69 585
R169 B.n321 B.n320 585
R170 B.n319 B.n70 585
R171 B.n318 B.n317 585
R172 B.n316 B.n71 585
R173 B.n315 B.n314 585
R174 B.n313 B.n72 585
R175 B.n312 B.n311 585
R176 B.n310 B.n73 585
R177 B.n309 B.n308 585
R178 B.n307 B.n74 585
R179 B.n306 B.n305 585
R180 B.n304 B.n75 585
R181 B.n303 B.n302 585
R182 B.n301 B.n76 585
R183 B.n300 B.n299 585
R184 B.n298 B.n77 585
R185 B.n297 B.n296 585
R186 B.n295 B.n78 585
R187 B.n294 B.n293 585
R188 B.n292 B.n79 585
R189 B.n291 B.n290 585
R190 B.n289 B.n80 585
R191 B.n288 B.n287 585
R192 B.n286 B.n81 585
R193 B.n285 B.n284 585
R194 B.n283 B.n82 585
R195 B.n282 B.n281 585
R196 B.n280 B.n83 585
R197 B.n279 B.n278 585
R198 B.n277 B.n84 585
R199 B.n276 B.n275 585
R200 B.n274 B.n85 585
R201 B.n184 B.n119 585
R202 B.n186 B.n185 585
R203 B.n187 B.n118 585
R204 B.n189 B.n188 585
R205 B.n190 B.n117 585
R206 B.n192 B.n191 585
R207 B.n193 B.n116 585
R208 B.n195 B.n194 585
R209 B.n196 B.n115 585
R210 B.n198 B.n197 585
R211 B.n199 B.n114 585
R212 B.n201 B.n200 585
R213 B.n202 B.n113 585
R214 B.n204 B.n203 585
R215 B.n205 B.n112 585
R216 B.n207 B.n206 585
R217 B.n208 B.n111 585
R218 B.n210 B.n209 585
R219 B.n211 B.n110 585
R220 B.n213 B.n212 585
R221 B.n214 B.n109 585
R222 B.n216 B.n215 585
R223 B.n217 B.n108 585
R224 B.n219 B.n218 585
R225 B.n220 B.n105 585
R226 B.n223 B.n222 585
R227 B.n224 B.n104 585
R228 B.n226 B.n225 585
R229 B.n227 B.n103 585
R230 B.n229 B.n228 585
R231 B.n230 B.n102 585
R232 B.n232 B.n231 585
R233 B.n233 B.n101 585
R234 B.n235 B.n234 585
R235 B.n237 B.n236 585
R236 B.n238 B.n97 585
R237 B.n240 B.n239 585
R238 B.n241 B.n96 585
R239 B.n243 B.n242 585
R240 B.n244 B.n95 585
R241 B.n246 B.n245 585
R242 B.n247 B.n94 585
R243 B.n249 B.n248 585
R244 B.n250 B.n93 585
R245 B.n252 B.n251 585
R246 B.n253 B.n92 585
R247 B.n255 B.n254 585
R248 B.n256 B.n91 585
R249 B.n258 B.n257 585
R250 B.n259 B.n90 585
R251 B.n261 B.n260 585
R252 B.n262 B.n89 585
R253 B.n264 B.n263 585
R254 B.n265 B.n88 585
R255 B.n267 B.n266 585
R256 B.n268 B.n87 585
R257 B.n270 B.n269 585
R258 B.n271 B.n86 585
R259 B.n273 B.n272 585
R260 B.n183 B.n182 585
R261 B.n181 B.n120 585
R262 B.n180 B.n179 585
R263 B.n178 B.n121 585
R264 B.n177 B.n176 585
R265 B.n175 B.n122 585
R266 B.n174 B.n173 585
R267 B.n172 B.n123 585
R268 B.n171 B.n170 585
R269 B.n169 B.n124 585
R270 B.n168 B.n167 585
R271 B.n166 B.n125 585
R272 B.n165 B.n164 585
R273 B.n163 B.n126 585
R274 B.n162 B.n161 585
R275 B.n160 B.n127 585
R276 B.n159 B.n158 585
R277 B.n157 B.n128 585
R278 B.n156 B.n155 585
R279 B.n154 B.n129 585
R280 B.n153 B.n152 585
R281 B.n151 B.n130 585
R282 B.n150 B.n149 585
R283 B.n148 B.n131 585
R284 B.n147 B.n146 585
R285 B.n145 B.n132 585
R286 B.n144 B.n143 585
R287 B.n142 B.n133 585
R288 B.n141 B.n140 585
R289 B.n139 B.n134 585
R290 B.n138 B.n137 585
R291 B.n136 B.n135 585
R292 B.n2 B.n0 585
R293 B.n513 B.n1 585
R294 B.n512 B.n511 585
R295 B.n510 B.n3 585
R296 B.n509 B.n508 585
R297 B.n507 B.n4 585
R298 B.n506 B.n505 585
R299 B.n504 B.n5 585
R300 B.n503 B.n502 585
R301 B.n501 B.n6 585
R302 B.n500 B.n499 585
R303 B.n498 B.n7 585
R304 B.n497 B.n496 585
R305 B.n495 B.n8 585
R306 B.n494 B.n493 585
R307 B.n492 B.n9 585
R308 B.n491 B.n490 585
R309 B.n489 B.n10 585
R310 B.n488 B.n487 585
R311 B.n486 B.n11 585
R312 B.n485 B.n484 585
R313 B.n483 B.n12 585
R314 B.n482 B.n481 585
R315 B.n480 B.n13 585
R316 B.n479 B.n478 585
R317 B.n477 B.n14 585
R318 B.n476 B.n475 585
R319 B.n474 B.n15 585
R320 B.n473 B.n472 585
R321 B.n471 B.n16 585
R322 B.n470 B.n469 585
R323 B.n468 B.n17 585
R324 B.n467 B.n466 585
R325 B.n465 B.n18 585
R326 B.n515 B.n514 585
R327 B.n182 B.n119 468.476
R328 B.n465 B.n464 468.476
R329 B.n272 B.n85 468.476
R330 B.n374 B.n373 468.476
R331 B.n98 B.t9 291.421
R332 B.n106 B.t6 291.421
R333 B.n32 B.t3 291.421
R334 B.n38 B.t0 291.421
R335 B.n182 B.n181 163.367
R336 B.n181 B.n180 163.367
R337 B.n180 B.n121 163.367
R338 B.n176 B.n121 163.367
R339 B.n176 B.n175 163.367
R340 B.n175 B.n174 163.367
R341 B.n174 B.n123 163.367
R342 B.n170 B.n123 163.367
R343 B.n170 B.n169 163.367
R344 B.n169 B.n168 163.367
R345 B.n168 B.n125 163.367
R346 B.n164 B.n125 163.367
R347 B.n164 B.n163 163.367
R348 B.n163 B.n162 163.367
R349 B.n162 B.n127 163.367
R350 B.n158 B.n127 163.367
R351 B.n158 B.n157 163.367
R352 B.n157 B.n156 163.367
R353 B.n156 B.n129 163.367
R354 B.n152 B.n129 163.367
R355 B.n152 B.n151 163.367
R356 B.n151 B.n150 163.367
R357 B.n150 B.n131 163.367
R358 B.n146 B.n131 163.367
R359 B.n146 B.n145 163.367
R360 B.n145 B.n144 163.367
R361 B.n144 B.n133 163.367
R362 B.n140 B.n133 163.367
R363 B.n140 B.n139 163.367
R364 B.n139 B.n138 163.367
R365 B.n138 B.n135 163.367
R366 B.n135 B.n2 163.367
R367 B.n514 B.n2 163.367
R368 B.n514 B.n513 163.367
R369 B.n513 B.n512 163.367
R370 B.n512 B.n3 163.367
R371 B.n508 B.n3 163.367
R372 B.n508 B.n507 163.367
R373 B.n507 B.n506 163.367
R374 B.n506 B.n5 163.367
R375 B.n502 B.n5 163.367
R376 B.n502 B.n501 163.367
R377 B.n501 B.n500 163.367
R378 B.n500 B.n7 163.367
R379 B.n496 B.n7 163.367
R380 B.n496 B.n495 163.367
R381 B.n495 B.n494 163.367
R382 B.n494 B.n9 163.367
R383 B.n490 B.n9 163.367
R384 B.n490 B.n489 163.367
R385 B.n489 B.n488 163.367
R386 B.n488 B.n11 163.367
R387 B.n484 B.n11 163.367
R388 B.n484 B.n483 163.367
R389 B.n483 B.n482 163.367
R390 B.n482 B.n13 163.367
R391 B.n478 B.n13 163.367
R392 B.n478 B.n477 163.367
R393 B.n477 B.n476 163.367
R394 B.n476 B.n15 163.367
R395 B.n472 B.n15 163.367
R396 B.n472 B.n471 163.367
R397 B.n471 B.n470 163.367
R398 B.n470 B.n17 163.367
R399 B.n466 B.n17 163.367
R400 B.n466 B.n465 163.367
R401 B.n186 B.n119 163.367
R402 B.n187 B.n186 163.367
R403 B.n188 B.n187 163.367
R404 B.n188 B.n117 163.367
R405 B.n192 B.n117 163.367
R406 B.n193 B.n192 163.367
R407 B.n194 B.n193 163.367
R408 B.n194 B.n115 163.367
R409 B.n198 B.n115 163.367
R410 B.n199 B.n198 163.367
R411 B.n200 B.n199 163.367
R412 B.n200 B.n113 163.367
R413 B.n204 B.n113 163.367
R414 B.n205 B.n204 163.367
R415 B.n206 B.n205 163.367
R416 B.n206 B.n111 163.367
R417 B.n210 B.n111 163.367
R418 B.n211 B.n210 163.367
R419 B.n212 B.n211 163.367
R420 B.n212 B.n109 163.367
R421 B.n216 B.n109 163.367
R422 B.n217 B.n216 163.367
R423 B.n218 B.n217 163.367
R424 B.n218 B.n105 163.367
R425 B.n223 B.n105 163.367
R426 B.n224 B.n223 163.367
R427 B.n225 B.n224 163.367
R428 B.n225 B.n103 163.367
R429 B.n229 B.n103 163.367
R430 B.n230 B.n229 163.367
R431 B.n231 B.n230 163.367
R432 B.n231 B.n101 163.367
R433 B.n235 B.n101 163.367
R434 B.n236 B.n235 163.367
R435 B.n236 B.n97 163.367
R436 B.n240 B.n97 163.367
R437 B.n241 B.n240 163.367
R438 B.n242 B.n241 163.367
R439 B.n242 B.n95 163.367
R440 B.n246 B.n95 163.367
R441 B.n247 B.n246 163.367
R442 B.n248 B.n247 163.367
R443 B.n248 B.n93 163.367
R444 B.n252 B.n93 163.367
R445 B.n253 B.n252 163.367
R446 B.n254 B.n253 163.367
R447 B.n254 B.n91 163.367
R448 B.n258 B.n91 163.367
R449 B.n259 B.n258 163.367
R450 B.n260 B.n259 163.367
R451 B.n260 B.n89 163.367
R452 B.n264 B.n89 163.367
R453 B.n265 B.n264 163.367
R454 B.n266 B.n265 163.367
R455 B.n266 B.n87 163.367
R456 B.n270 B.n87 163.367
R457 B.n271 B.n270 163.367
R458 B.n272 B.n271 163.367
R459 B.n276 B.n85 163.367
R460 B.n277 B.n276 163.367
R461 B.n278 B.n277 163.367
R462 B.n278 B.n83 163.367
R463 B.n282 B.n83 163.367
R464 B.n283 B.n282 163.367
R465 B.n284 B.n283 163.367
R466 B.n284 B.n81 163.367
R467 B.n288 B.n81 163.367
R468 B.n289 B.n288 163.367
R469 B.n290 B.n289 163.367
R470 B.n290 B.n79 163.367
R471 B.n294 B.n79 163.367
R472 B.n295 B.n294 163.367
R473 B.n296 B.n295 163.367
R474 B.n296 B.n77 163.367
R475 B.n300 B.n77 163.367
R476 B.n301 B.n300 163.367
R477 B.n302 B.n301 163.367
R478 B.n302 B.n75 163.367
R479 B.n306 B.n75 163.367
R480 B.n307 B.n306 163.367
R481 B.n308 B.n307 163.367
R482 B.n308 B.n73 163.367
R483 B.n312 B.n73 163.367
R484 B.n313 B.n312 163.367
R485 B.n314 B.n313 163.367
R486 B.n314 B.n71 163.367
R487 B.n318 B.n71 163.367
R488 B.n319 B.n318 163.367
R489 B.n320 B.n319 163.367
R490 B.n320 B.n69 163.367
R491 B.n324 B.n69 163.367
R492 B.n325 B.n324 163.367
R493 B.n326 B.n325 163.367
R494 B.n326 B.n67 163.367
R495 B.n330 B.n67 163.367
R496 B.n331 B.n330 163.367
R497 B.n332 B.n331 163.367
R498 B.n332 B.n65 163.367
R499 B.n336 B.n65 163.367
R500 B.n337 B.n336 163.367
R501 B.n338 B.n337 163.367
R502 B.n338 B.n63 163.367
R503 B.n342 B.n63 163.367
R504 B.n343 B.n342 163.367
R505 B.n344 B.n343 163.367
R506 B.n344 B.n61 163.367
R507 B.n348 B.n61 163.367
R508 B.n349 B.n348 163.367
R509 B.n350 B.n349 163.367
R510 B.n350 B.n59 163.367
R511 B.n354 B.n59 163.367
R512 B.n355 B.n354 163.367
R513 B.n356 B.n355 163.367
R514 B.n356 B.n57 163.367
R515 B.n360 B.n57 163.367
R516 B.n361 B.n360 163.367
R517 B.n362 B.n361 163.367
R518 B.n362 B.n55 163.367
R519 B.n366 B.n55 163.367
R520 B.n367 B.n366 163.367
R521 B.n368 B.n367 163.367
R522 B.n368 B.n53 163.367
R523 B.n372 B.n53 163.367
R524 B.n373 B.n372 163.367
R525 B.n464 B.n19 163.367
R526 B.n460 B.n19 163.367
R527 B.n460 B.n459 163.367
R528 B.n459 B.n458 163.367
R529 B.n458 B.n21 163.367
R530 B.n454 B.n21 163.367
R531 B.n454 B.n453 163.367
R532 B.n453 B.n452 163.367
R533 B.n452 B.n23 163.367
R534 B.n448 B.n23 163.367
R535 B.n448 B.n447 163.367
R536 B.n447 B.n446 163.367
R537 B.n446 B.n25 163.367
R538 B.n442 B.n25 163.367
R539 B.n442 B.n441 163.367
R540 B.n441 B.n440 163.367
R541 B.n440 B.n27 163.367
R542 B.n436 B.n27 163.367
R543 B.n436 B.n435 163.367
R544 B.n435 B.n434 163.367
R545 B.n434 B.n29 163.367
R546 B.n430 B.n29 163.367
R547 B.n430 B.n429 163.367
R548 B.n429 B.n428 163.367
R549 B.n428 B.n31 163.367
R550 B.n423 B.n31 163.367
R551 B.n423 B.n422 163.367
R552 B.n422 B.n421 163.367
R553 B.n421 B.n35 163.367
R554 B.n417 B.n35 163.367
R555 B.n417 B.n416 163.367
R556 B.n416 B.n415 163.367
R557 B.n415 B.n37 163.367
R558 B.n410 B.n37 163.367
R559 B.n410 B.n409 163.367
R560 B.n409 B.n408 163.367
R561 B.n408 B.n41 163.367
R562 B.n404 B.n41 163.367
R563 B.n404 B.n403 163.367
R564 B.n403 B.n402 163.367
R565 B.n402 B.n43 163.367
R566 B.n398 B.n43 163.367
R567 B.n398 B.n397 163.367
R568 B.n397 B.n396 163.367
R569 B.n396 B.n45 163.367
R570 B.n392 B.n45 163.367
R571 B.n392 B.n391 163.367
R572 B.n391 B.n390 163.367
R573 B.n390 B.n47 163.367
R574 B.n386 B.n47 163.367
R575 B.n386 B.n385 163.367
R576 B.n385 B.n384 163.367
R577 B.n384 B.n49 163.367
R578 B.n380 B.n49 163.367
R579 B.n380 B.n379 163.367
R580 B.n379 B.n378 163.367
R581 B.n378 B.n51 163.367
R582 B.n374 B.n51 163.367
R583 B.n98 B.t11 153.911
R584 B.n38 B.t1 153.911
R585 B.n106 B.t8 153.905
R586 B.n32 B.t4 153.905
R587 B.n99 B.t10 113.183
R588 B.n39 B.t2 113.183
R589 B.n107 B.t7 113.177
R590 B.n33 B.t5 113.177
R591 B.n100 B.n99 59.5399
R592 B.n221 B.n107 59.5399
R593 B.n426 B.n33 59.5399
R594 B.n412 B.n39 59.5399
R595 B.n99 B.n98 40.7278
R596 B.n107 B.n106 40.7278
R597 B.n33 B.n32 40.7278
R598 B.n39 B.n38 40.7278
R599 B.n463 B.n18 30.4395
R600 B.n274 B.n273 30.4395
R601 B.n184 B.n183 30.4395
R602 B.n375 B.n52 30.4395
R603 B B.n515 18.0485
R604 B.n463 B.n462 10.6151
R605 B.n462 B.n461 10.6151
R606 B.n461 B.n20 10.6151
R607 B.n457 B.n20 10.6151
R608 B.n457 B.n456 10.6151
R609 B.n456 B.n455 10.6151
R610 B.n455 B.n22 10.6151
R611 B.n451 B.n22 10.6151
R612 B.n451 B.n450 10.6151
R613 B.n450 B.n449 10.6151
R614 B.n449 B.n24 10.6151
R615 B.n445 B.n24 10.6151
R616 B.n445 B.n444 10.6151
R617 B.n444 B.n443 10.6151
R618 B.n443 B.n26 10.6151
R619 B.n439 B.n26 10.6151
R620 B.n439 B.n438 10.6151
R621 B.n438 B.n437 10.6151
R622 B.n437 B.n28 10.6151
R623 B.n433 B.n28 10.6151
R624 B.n433 B.n432 10.6151
R625 B.n432 B.n431 10.6151
R626 B.n431 B.n30 10.6151
R627 B.n427 B.n30 10.6151
R628 B.n425 B.n424 10.6151
R629 B.n424 B.n34 10.6151
R630 B.n420 B.n34 10.6151
R631 B.n420 B.n419 10.6151
R632 B.n419 B.n418 10.6151
R633 B.n418 B.n36 10.6151
R634 B.n414 B.n36 10.6151
R635 B.n414 B.n413 10.6151
R636 B.n411 B.n40 10.6151
R637 B.n407 B.n40 10.6151
R638 B.n407 B.n406 10.6151
R639 B.n406 B.n405 10.6151
R640 B.n405 B.n42 10.6151
R641 B.n401 B.n42 10.6151
R642 B.n401 B.n400 10.6151
R643 B.n400 B.n399 10.6151
R644 B.n399 B.n44 10.6151
R645 B.n395 B.n44 10.6151
R646 B.n395 B.n394 10.6151
R647 B.n394 B.n393 10.6151
R648 B.n393 B.n46 10.6151
R649 B.n389 B.n46 10.6151
R650 B.n389 B.n388 10.6151
R651 B.n388 B.n387 10.6151
R652 B.n387 B.n48 10.6151
R653 B.n383 B.n48 10.6151
R654 B.n383 B.n382 10.6151
R655 B.n382 B.n381 10.6151
R656 B.n381 B.n50 10.6151
R657 B.n377 B.n50 10.6151
R658 B.n377 B.n376 10.6151
R659 B.n376 B.n375 10.6151
R660 B.n275 B.n274 10.6151
R661 B.n275 B.n84 10.6151
R662 B.n279 B.n84 10.6151
R663 B.n280 B.n279 10.6151
R664 B.n281 B.n280 10.6151
R665 B.n281 B.n82 10.6151
R666 B.n285 B.n82 10.6151
R667 B.n286 B.n285 10.6151
R668 B.n287 B.n286 10.6151
R669 B.n287 B.n80 10.6151
R670 B.n291 B.n80 10.6151
R671 B.n292 B.n291 10.6151
R672 B.n293 B.n292 10.6151
R673 B.n293 B.n78 10.6151
R674 B.n297 B.n78 10.6151
R675 B.n298 B.n297 10.6151
R676 B.n299 B.n298 10.6151
R677 B.n299 B.n76 10.6151
R678 B.n303 B.n76 10.6151
R679 B.n304 B.n303 10.6151
R680 B.n305 B.n304 10.6151
R681 B.n305 B.n74 10.6151
R682 B.n309 B.n74 10.6151
R683 B.n310 B.n309 10.6151
R684 B.n311 B.n310 10.6151
R685 B.n311 B.n72 10.6151
R686 B.n315 B.n72 10.6151
R687 B.n316 B.n315 10.6151
R688 B.n317 B.n316 10.6151
R689 B.n317 B.n70 10.6151
R690 B.n321 B.n70 10.6151
R691 B.n322 B.n321 10.6151
R692 B.n323 B.n322 10.6151
R693 B.n323 B.n68 10.6151
R694 B.n327 B.n68 10.6151
R695 B.n328 B.n327 10.6151
R696 B.n329 B.n328 10.6151
R697 B.n329 B.n66 10.6151
R698 B.n333 B.n66 10.6151
R699 B.n334 B.n333 10.6151
R700 B.n335 B.n334 10.6151
R701 B.n335 B.n64 10.6151
R702 B.n339 B.n64 10.6151
R703 B.n340 B.n339 10.6151
R704 B.n341 B.n340 10.6151
R705 B.n341 B.n62 10.6151
R706 B.n345 B.n62 10.6151
R707 B.n346 B.n345 10.6151
R708 B.n347 B.n346 10.6151
R709 B.n347 B.n60 10.6151
R710 B.n351 B.n60 10.6151
R711 B.n352 B.n351 10.6151
R712 B.n353 B.n352 10.6151
R713 B.n353 B.n58 10.6151
R714 B.n357 B.n58 10.6151
R715 B.n358 B.n357 10.6151
R716 B.n359 B.n358 10.6151
R717 B.n359 B.n56 10.6151
R718 B.n363 B.n56 10.6151
R719 B.n364 B.n363 10.6151
R720 B.n365 B.n364 10.6151
R721 B.n365 B.n54 10.6151
R722 B.n369 B.n54 10.6151
R723 B.n370 B.n369 10.6151
R724 B.n371 B.n370 10.6151
R725 B.n371 B.n52 10.6151
R726 B.n185 B.n184 10.6151
R727 B.n185 B.n118 10.6151
R728 B.n189 B.n118 10.6151
R729 B.n190 B.n189 10.6151
R730 B.n191 B.n190 10.6151
R731 B.n191 B.n116 10.6151
R732 B.n195 B.n116 10.6151
R733 B.n196 B.n195 10.6151
R734 B.n197 B.n196 10.6151
R735 B.n197 B.n114 10.6151
R736 B.n201 B.n114 10.6151
R737 B.n202 B.n201 10.6151
R738 B.n203 B.n202 10.6151
R739 B.n203 B.n112 10.6151
R740 B.n207 B.n112 10.6151
R741 B.n208 B.n207 10.6151
R742 B.n209 B.n208 10.6151
R743 B.n209 B.n110 10.6151
R744 B.n213 B.n110 10.6151
R745 B.n214 B.n213 10.6151
R746 B.n215 B.n214 10.6151
R747 B.n215 B.n108 10.6151
R748 B.n219 B.n108 10.6151
R749 B.n220 B.n219 10.6151
R750 B.n222 B.n104 10.6151
R751 B.n226 B.n104 10.6151
R752 B.n227 B.n226 10.6151
R753 B.n228 B.n227 10.6151
R754 B.n228 B.n102 10.6151
R755 B.n232 B.n102 10.6151
R756 B.n233 B.n232 10.6151
R757 B.n234 B.n233 10.6151
R758 B.n238 B.n237 10.6151
R759 B.n239 B.n238 10.6151
R760 B.n239 B.n96 10.6151
R761 B.n243 B.n96 10.6151
R762 B.n244 B.n243 10.6151
R763 B.n245 B.n244 10.6151
R764 B.n245 B.n94 10.6151
R765 B.n249 B.n94 10.6151
R766 B.n250 B.n249 10.6151
R767 B.n251 B.n250 10.6151
R768 B.n251 B.n92 10.6151
R769 B.n255 B.n92 10.6151
R770 B.n256 B.n255 10.6151
R771 B.n257 B.n256 10.6151
R772 B.n257 B.n90 10.6151
R773 B.n261 B.n90 10.6151
R774 B.n262 B.n261 10.6151
R775 B.n263 B.n262 10.6151
R776 B.n263 B.n88 10.6151
R777 B.n267 B.n88 10.6151
R778 B.n268 B.n267 10.6151
R779 B.n269 B.n268 10.6151
R780 B.n269 B.n86 10.6151
R781 B.n273 B.n86 10.6151
R782 B.n183 B.n120 10.6151
R783 B.n179 B.n120 10.6151
R784 B.n179 B.n178 10.6151
R785 B.n178 B.n177 10.6151
R786 B.n177 B.n122 10.6151
R787 B.n173 B.n122 10.6151
R788 B.n173 B.n172 10.6151
R789 B.n172 B.n171 10.6151
R790 B.n171 B.n124 10.6151
R791 B.n167 B.n124 10.6151
R792 B.n167 B.n166 10.6151
R793 B.n166 B.n165 10.6151
R794 B.n165 B.n126 10.6151
R795 B.n161 B.n126 10.6151
R796 B.n161 B.n160 10.6151
R797 B.n160 B.n159 10.6151
R798 B.n159 B.n128 10.6151
R799 B.n155 B.n128 10.6151
R800 B.n155 B.n154 10.6151
R801 B.n154 B.n153 10.6151
R802 B.n153 B.n130 10.6151
R803 B.n149 B.n130 10.6151
R804 B.n149 B.n148 10.6151
R805 B.n148 B.n147 10.6151
R806 B.n147 B.n132 10.6151
R807 B.n143 B.n132 10.6151
R808 B.n143 B.n142 10.6151
R809 B.n142 B.n141 10.6151
R810 B.n141 B.n134 10.6151
R811 B.n137 B.n134 10.6151
R812 B.n137 B.n136 10.6151
R813 B.n136 B.n0 10.6151
R814 B.n511 B.n1 10.6151
R815 B.n511 B.n510 10.6151
R816 B.n510 B.n509 10.6151
R817 B.n509 B.n4 10.6151
R818 B.n505 B.n4 10.6151
R819 B.n505 B.n504 10.6151
R820 B.n504 B.n503 10.6151
R821 B.n503 B.n6 10.6151
R822 B.n499 B.n6 10.6151
R823 B.n499 B.n498 10.6151
R824 B.n498 B.n497 10.6151
R825 B.n497 B.n8 10.6151
R826 B.n493 B.n8 10.6151
R827 B.n493 B.n492 10.6151
R828 B.n492 B.n491 10.6151
R829 B.n491 B.n10 10.6151
R830 B.n487 B.n10 10.6151
R831 B.n487 B.n486 10.6151
R832 B.n486 B.n485 10.6151
R833 B.n485 B.n12 10.6151
R834 B.n481 B.n12 10.6151
R835 B.n481 B.n480 10.6151
R836 B.n480 B.n479 10.6151
R837 B.n479 B.n14 10.6151
R838 B.n475 B.n14 10.6151
R839 B.n475 B.n474 10.6151
R840 B.n474 B.n473 10.6151
R841 B.n473 B.n16 10.6151
R842 B.n469 B.n16 10.6151
R843 B.n469 B.n468 10.6151
R844 B.n468 B.n467 10.6151
R845 B.n467 B.n18 10.6151
R846 B.n426 B.n425 6.5566
R847 B.n413 B.n412 6.5566
R848 B.n222 B.n221 6.5566
R849 B.n234 B.n100 6.5566
R850 B.n427 B.n426 4.05904
R851 B.n412 B.n411 4.05904
R852 B.n221 B.n220 4.05904
R853 B.n237 B.n100 4.05904
R854 B.n515 B.n0 2.81026
R855 B.n515 B.n1 2.81026
R856 VP.n18 VP.n17 180.875
R857 VP.n33 VP.n32 180.875
R858 VP.n16 VP.n15 180.875
R859 VP.n10 VP.n9 161.3
R860 VP.n11 VP.n6 161.3
R861 VP.n13 VP.n12 161.3
R862 VP.n14 VP.n5 161.3
R863 VP.n31 VP.n0 161.3
R864 VP.n30 VP.n29 161.3
R865 VP.n28 VP.n1 161.3
R866 VP.n27 VP.n26 161.3
R867 VP.n25 VP.n2 161.3
R868 VP.n24 VP.n23 161.3
R869 VP.n22 VP.n3 161.3
R870 VP.n21 VP.n20 161.3
R871 VP.n19 VP.n4 161.3
R872 VP.n7 VP.t4 120.436
R873 VP.n25 VP.t3 85.0994
R874 VP.n18 VP.t5 85.0994
R875 VP.n32 VP.t1 85.0994
R876 VP.n8 VP.t0 85.0994
R877 VP.n15 VP.t2 85.0994
R878 VP.n20 VP.n3 45.3497
R879 VP.n30 VP.n1 45.3497
R880 VP.n13 VP.n6 45.3497
R881 VP.n8 VP.n7 44.5155
R882 VP.n17 VP.n16 40.9778
R883 VP.n24 VP.n3 35.6371
R884 VP.n26 VP.n1 35.6371
R885 VP.n9 VP.n6 35.6371
R886 VP.n20 VP.n19 24.4675
R887 VP.n25 VP.n24 24.4675
R888 VP.n26 VP.n25 24.4675
R889 VP.n31 VP.n30 24.4675
R890 VP.n14 VP.n13 24.4675
R891 VP.n9 VP.n8 24.4675
R892 VP.n10 VP.n7 12.2033
R893 VP.n19 VP.n18 4.8939
R894 VP.n32 VP.n31 4.8939
R895 VP.n15 VP.n14 4.8939
R896 VP.n11 VP.n10 0.189894
R897 VP.n12 VP.n11 0.189894
R898 VP.n12 VP.n5 0.189894
R899 VP.n16 VP.n5 0.189894
R900 VP.n17 VP.n4 0.189894
R901 VP.n21 VP.n4 0.189894
R902 VP.n22 VP.n21 0.189894
R903 VP.n23 VP.n22 0.189894
R904 VP.n23 VP.n2 0.189894
R905 VP.n27 VP.n2 0.189894
R906 VP.n28 VP.n27 0.189894
R907 VP.n29 VP.n28 0.189894
R908 VP.n29 VP.n0 0.189894
R909 VP.n33 VP.n0 0.189894
R910 VP VP.n33 0.0516364
R911 VDD1 VDD1.t1 94.7118
R912 VDD1.n1 VDD1.t0 94.5982
R913 VDD1.n1 VDD1.n0 88.4921
R914 VDD1.n3 VDD1.n2 88.0949
R915 VDD1.n3 VDD1.n1 36.475
R916 VDD1.n2 VDD1.t5 5.2013
R917 VDD1.n2 VDD1.t3 5.2013
R918 VDD1.n0 VDD1.t2 5.2013
R919 VDD1.n0 VDD1.t4 5.2013
R920 VDD1 VDD1.n3 0.394897
C0 w_n2650_n2218# VP 5.05322f
C1 B VN 0.921599f
C2 VDD2 VTAIL 5.41339f
C3 B VTAIL 2.11755f
C4 VN VDD1 0.149462f
C5 VDD2 VP 0.387289f
C6 B VP 1.48558f
C7 VTAIL VDD1 5.3674f
C8 VTAIL VN 3.69838f
C9 VDD2 w_n2650_n2218# 1.73701f
C10 VDD1 VP 3.62625f
C11 B w_n2650_n2218# 6.92342f
C12 VN VP 5.05422f
C13 w_n2650_n2218# VDD1 1.67852f
C14 VTAIL VP 3.71263f
C15 w_n2650_n2218# VN 4.71292f
C16 VDD2 B 1.48141f
C17 w_n2650_n2218# VTAIL 2.08059f
C18 VDD2 VDD1 1.10737f
C19 VDD2 VN 3.39063f
C20 B VDD1 1.42718f
C21 VDD2 VSUBS 1.259185f
C22 VDD1 VSUBS 1.652959f
C23 VTAIL VSUBS 0.599727f
C24 VN VSUBS 4.75688f
C25 VP VSUBS 1.946599f
C26 B VSUBS 3.330397f
C27 w_n2650_n2218# VSUBS 73.298996f
C28 VDD1.t1 VSUBS 0.987952f
C29 VDD1.t0 VSUBS 0.987215f
C30 VDD1.t2 VSUBS 0.109737f
C31 VDD1.t4 VSUBS 0.109737f
C32 VDD1.n0 VSUBS 0.734528f
C33 VDD1.n1 VSUBS 2.40892f
C34 VDD1.t5 VSUBS 0.109737f
C35 VDD1.t3 VSUBS 0.109737f
C36 VDD1.n2 VSUBS 0.732117f
C37 VDD1.n3 VSUBS 2.05836f
C38 VP.n0 VSUBS 0.046054f
C39 VP.t1 VSUBS 1.35163f
C40 VP.n1 VSUBS 0.03873f
C41 VP.n2 VSUBS 0.046054f
C42 VP.t3 VSUBS 1.35163f
C43 VP.n3 VSUBS 0.03873f
C44 VP.n4 VSUBS 0.046054f
C45 VP.t5 VSUBS 1.35163f
C46 VP.n5 VSUBS 0.046054f
C47 VP.t2 VSUBS 1.35163f
C48 VP.n6 VSUBS 0.03873f
C49 VP.t4 VSUBS 1.56711f
C50 VP.n7 VSUBS 0.608911f
C51 VP.t0 VSUBS 1.35163f
C52 VP.n8 VSUBS 0.641905f
C53 VP.n9 VSUBS 0.093002f
C54 VP.n10 VSUBS 0.338898f
C55 VP.n11 VSUBS 0.046054f
C56 VP.n12 VSUBS 0.046054f
C57 VP.n13 VSUBS 0.088561f
C58 VP.n14 VSUBS 0.051932f
C59 VP.n15 VSUBS 0.62281f
C60 VP.n16 VSUBS 1.83652f
C61 VP.n17 VSUBS 1.87692f
C62 VP.n18 VSUBS 0.62281f
C63 VP.n19 VSUBS 0.051932f
C64 VP.n20 VSUBS 0.088561f
C65 VP.n21 VSUBS 0.046054f
C66 VP.n22 VSUBS 0.046054f
C67 VP.n23 VSUBS 0.046054f
C68 VP.n24 VSUBS 0.093002f
C69 VP.n25 VSUBS 0.561758f
C70 VP.n26 VSUBS 0.093002f
C71 VP.n27 VSUBS 0.046054f
C72 VP.n28 VSUBS 0.046054f
C73 VP.n29 VSUBS 0.046054f
C74 VP.n30 VSUBS 0.088561f
C75 VP.n31 VSUBS 0.051932f
C76 VP.n32 VSUBS 0.62281f
C77 VP.n33 VSUBS 0.048372f
C78 B.n0 VSUBS 0.00497f
C79 B.n1 VSUBS 0.00497f
C80 B.n2 VSUBS 0.00786f
C81 B.n3 VSUBS 0.00786f
C82 B.n4 VSUBS 0.00786f
C83 B.n5 VSUBS 0.00786f
C84 B.n6 VSUBS 0.00786f
C85 B.n7 VSUBS 0.00786f
C86 B.n8 VSUBS 0.00786f
C87 B.n9 VSUBS 0.00786f
C88 B.n10 VSUBS 0.00786f
C89 B.n11 VSUBS 0.00786f
C90 B.n12 VSUBS 0.00786f
C91 B.n13 VSUBS 0.00786f
C92 B.n14 VSUBS 0.00786f
C93 B.n15 VSUBS 0.00786f
C94 B.n16 VSUBS 0.00786f
C95 B.n17 VSUBS 0.00786f
C96 B.n18 VSUBS 0.017241f
C97 B.n19 VSUBS 0.00786f
C98 B.n20 VSUBS 0.00786f
C99 B.n21 VSUBS 0.00786f
C100 B.n22 VSUBS 0.00786f
C101 B.n23 VSUBS 0.00786f
C102 B.n24 VSUBS 0.00786f
C103 B.n25 VSUBS 0.00786f
C104 B.n26 VSUBS 0.00786f
C105 B.n27 VSUBS 0.00786f
C106 B.n28 VSUBS 0.00786f
C107 B.n29 VSUBS 0.00786f
C108 B.n30 VSUBS 0.00786f
C109 B.n31 VSUBS 0.00786f
C110 B.t5 VSUBS 0.20665f
C111 B.t4 VSUBS 0.223734f
C112 B.t3 VSUBS 0.573815f
C113 B.n32 VSUBS 0.123067f
C114 B.n33 VSUBS 0.075771f
C115 B.n34 VSUBS 0.00786f
C116 B.n35 VSUBS 0.00786f
C117 B.n36 VSUBS 0.00786f
C118 B.n37 VSUBS 0.00786f
C119 B.t2 VSUBS 0.206649f
C120 B.t1 VSUBS 0.223733f
C121 B.t0 VSUBS 0.573815f
C122 B.n38 VSUBS 0.123069f
C123 B.n39 VSUBS 0.075771f
C124 B.n40 VSUBS 0.00786f
C125 B.n41 VSUBS 0.00786f
C126 B.n42 VSUBS 0.00786f
C127 B.n43 VSUBS 0.00786f
C128 B.n44 VSUBS 0.00786f
C129 B.n45 VSUBS 0.00786f
C130 B.n46 VSUBS 0.00786f
C131 B.n47 VSUBS 0.00786f
C132 B.n48 VSUBS 0.00786f
C133 B.n49 VSUBS 0.00786f
C134 B.n50 VSUBS 0.00786f
C135 B.n51 VSUBS 0.00786f
C136 B.n52 VSUBS 0.018237f
C137 B.n53 VSUBS 0.00786f
C138 B.n54 VSUBS 0.00786f
C139 B.n55 VSUBS 0.00786f
C140 B.n56 VSUBS 0.00786f
C141 B.n57 VSUBS 0.00786f
C142 B.n58 VSUBS 0.00786f
C143 B.n59 VSUBS 0.00786f
C144 B.n60 VSUBS 0.00786f
C145 B.n61 VSUBS 0.00786f
C146 B.n62 VSUBS 0.00786f
C147 B.n63 VSUBS 0.00786f
C148 B.n64 VSUBS 0.00786f
C149 B.n65 VSUBS 0.00786f
C150 B.n66 VSUBS 0.00786f
C151 B.n67 VSUBS 0.00786f
C152 B.n68 VSUBS 0.00786f
C153 B.n69 VSUBS 0.00786f
C154 B.n70 VSUBS 0.00786f
C155 B.n71 VSUBS 0.00786f
C156 B.n72 VSUBS 0.00786f
C157 B.n73 VSUBS 0.00786f
C158 B.n74 VSUBS 0.00786f
C159 B.n75 VSUBS 0.00786f
C160 B.n76 VSUBS 0.00786f
C161 B.n77 VSUBS 0.00786f
C162 B.n78 VSUBS 0.00786f
C163 B.n79 VSUBS 0.00786f
C164 B.n80 VSUBS 0.00786f
C165 B.n81 VSUBS 0.00786f
C166 B.n82 VSUBS 0.00786f
C167 B.n83 VSUBS 0.00786f
C168 B.n84 VSUBS 0.00786f
C169 B.n85 VSUBS 0.017241f
C170 B.n86 VSUBS 0.00786f
C171 B.n87 VSUBS 0.00786f
C172 B.n88 VSUBS 0.00786f
C173 B.n89 VSUBS 0.00786f
C174 B.n90 VSUBS 0.00786f
C175 B.n91 VSUBS 0.00786f
C176 B.n92 VSUBS 0.00786f
C177 B.n93 VSUBS 0.00786f
C178 B.n94 VSUBS 0.00786f
C179 B.n95 VSUBS 0.00786f
C180 B.n96 VSUBS 0.00786f
C181 B.n97 VSUBS 0.00786f
C182 B.t10 VSUBS 0.206649f
C183 B.t11 VSUBS 0.223733f
C184 B.t9 VSUBS 0.573815f
C185 B.n98 VSUBS 0.123069f
C186 B.n99 VSUBS 0.075771f
C187 B.n100 VSUBS 0.01821f
C188 B.n101 VSUBS 0.00786f
C189 B.n102 VSUBS 0.00786f
C190 B.n103 VSUBS 0.00786f
C191 B.n104 VSUBS 0.00786f
C192 B.n105 VSUBS 0.00786f
C193 B.t7 VSUBS 0.20665f
C194 B.t8 VSUBS 0.223734f
C195 B.t6 VSUBS 0.573815f
C196 B.n106 VSUBS 0.123067f
C197 B.n107 VSUBS 0.075771f
C198 B.n108 VSUBS 0.00786f
C199 B.n109 VSUBS 0.00786f
C200 B.n110 VSUBS 0.00786f
C201 B.n111 VSUBS 0.00786f
C202 B.n112 VSUBS 0.00786f
C203 B.n113 VSUBS 0.00786f
C204 B.n114 VSUBS 0.00786f
C205 B.n115 VSUBS 0.00786f
C206 B.n116 VSUBS 0.00786f
C207 B.n117 VSUBS 0.00786f
C208 B.n118 VSUBS 0.00786f
C209 B.n119 VSUBS 0.017897f
C210 B.n120 VSUBS 0.00786f
C211 B.n121 VSUBS 0.00786f
C212 B.n122 VSUBS 0.00786f
C213 B.n123 VSUBS 0.00786f
C214 B.n124 VSUBS 0.00786f
C215 B.n125 VSUBS 0.00786f
C216 B.n126 VSUBS 0.00786f
C217 B.n127 VSUBS 0.00786f
C218 B.n128 VSUBS 0.00786f
C219 B.n129 VSUBS 0.00786f
C220 B.n130 VSUBS 0.00786f
C221 B.n131 VSUBS 0.00786f
C222 B.n132 VSUBS 0.00786f
C223 B.n133 VSUBS 0.00786f
C224 B.n134 VSUBS 0.00786f
C225 B.n135 VSUBS 0.00786f
C226 B.n136 VSUBS 0.00786f
C227 B.n137 VSUBS 0.00786f
C228 B.n138 VSUBS 0.00786f
C229 B.n139 VSUBS 0.00786f
C230 B.n140 VSUBS 0.00786f
C231 B.n141 VSUBS 0.00786f
C232 B.n142 VSUBS 0.00786f
C233 B.n143 VSUBS 0.00786f
C234 B.n144 VSUBS 0.00786f
C235 B.n145 VSUBS 0.00786f
C236 B.n146 VSUBS 0.00786f
C237 B.n147 VSUBS 0.00786f
C238 B.n148 VSUBS 0.00786f
C239 B.n149 VSUBS 0.00786f
C240 B.n150 VSUBS 0.00786f
C241 B.n151 VSUBS 0.00786f
C242 B.n152 VSUBS 0.00786f
C243 B.n153 VSUBS 0.00786f
C244 B.n154 VSUBS 0.00786f
C245 B.n155 VSUBS 0.00786f
C246 B.n156 VSUBS 0.00786f
C247 B.n157 VSUBS 0.00786f
C248 B.n158 VSUBS 0.00786f
C249 B.n159 VSUBS 0.00786f
C250 B.n160 VSUBS 0.00786f
C251 B.n161 VSUBS 0.00786f
C252 B.n162 VSUBS 0.00786f
C253 B.n163 VSUBS 0.00786f
C254 B.n164 VSUBS 0.00786f
C255 B.n165 VSUBS 0.00786f
C256 B.n166 VSUBS 0.00786f
C257 B.n167 VSUBS 0.00786f
C258 B.n168 VSUBS 0.00786f
C259 B.n169 VSUBS 0.00786f
C260 B.n170 VSUBS 0.00786f
C261 B.n171 VSUBS 0.00786f
C262 B.n172 VSUBS 0.00786f
C263 B.n173 VSUBS 0.00786f
C264 B.n174 VSUBS 0.00786f
C265 B.n175 VSUBS 0.00786f
C266 B.n176 VSUBS 0.00786f
C267 B.n177 VSUBS 0.00786f
C268 B.n178 VSUBS 0.00786f
C269 B.n179 VSUBS 0.00786f
C270 B.n180 VSUBS 0.00786f
C271 B.n181 VSUBS 0.00786f
C272 B.n182 VSUBS 0.017241f
C273 B.n183 VSUBS 0.017241f
C274 B.n184 VSUBS 0.017897f
C275 B.n185 VSUBS 0.00786f
C276 B.n186 VSUBS 0.00786f
C277 B.n187 VSUBS 0.00786f
C278 B.n188 VSUBS 0.00786f
C279 B.n189 VSUBS 0.00786f
C280 B.n190 VSUBS 0.00786f
C281 B.n191 VSUBS 0.00786f
C282 B.n192 VSUBS 0.00786f
C283 B.n193 VSUBS 0.00786f
C284 B.n194 VSUBS 0.00786f
C285 B.n195 VSUBS 0.00786f
C286 B.n196 VSUBS 0.00786f
C287 B.n197 VSUBS 0.00786f
C288 B.n198 VSUBS 0.00786f
C289 B.n199 VSUBS 0.00786f
C290 B.n200 VSUBS 0.00786f
C291 B.n201 VSUBS 0.00786f
C292 B.n202 VSUBS 0.00786f
C293 B.n203 VSUBS 0.00786f
C294 B.n204 VSUBS 0.00786f
C295 B.n205 VSUBS 0.00786f
C296 B.n206 VSUBS 0.00786f
C297 B.n207 VSUBS 0.00786f
C298 B.n208 VSUBS 0.00786f
C299 B.n209 VSUBS 0.00786f
C300 B.n210 VSUBS 0.00786f
C301 B.n211 VSUBS 0.00786f
C302 B.n212 VSUBS 0.00786f
C303 B.n213 VSUBS 0.00786f
C304 B.n214 VSUBS 0.00786f
C305 B.n215 VSUBS 0.00786f
C306 B.n216 VSUBS 0.00786f
C307 B.n217 VSUBS 0.00786f
C308 B.n218 VSUBS 0.00786f
C309 B.n219 VSUBS 0.00786f
C310 B.n220 VSUBS 0.005432f
C311 B.n221 VSUBS 0.01821f
C312 B.n222 VSUBS 0.006357f
C313 B.n223 VSUBS 0.00786f
C314 B.n224 VSUBS 0.00786f
C315 B.n225 VSUBS 0.00786f
C316 B.n226 VSUBS 0.00786f
C317 B.n227 VSUBS 0.00786f
C318 B.n228 VSUBS 0.00786f
C319 B.n229 VSUBS 0.00786f
C320 B.n230 VSUBS 0.00786f
C321 B.n231 VSUBS 0.00786f
C322 B.n232 VSUBS 0.00786f
C323 B.n233 VSUBS 0.00786f
C324 B.n234 VSUBS 0.006357f
C325 B.n235 VSUBS 0.00786f
C326 B.n236 VSUBS 0.00786f
C327 B.n237 VSUBS 0.005432f
C328 B.n238 VSUBS 0.00786f
C329 B.n239 VSUBS 0.00786f
C330 B.n240 VSUBS 0.00786f
C331 B.n241 VSUBS 0.00786f
C332 B.n242 VSUBS 0.00786f
C333 B.n243 VSUBS 0.00786f
C334 B.n244 VSUBS 0.00786f
C335 B.n245 VSUBS 0.00786f
C336 B.n246 VSUBS 0.00786f
C337 B.n247 VSUBS 0.00786f
C338 B.n248 VSUBS 0.00786f
C339 B.n249 VSUBS 0.00786f
C340 B.n250 VSUBS 0.00786f
C341 B.n251 VSUBS 0.00786f
C342 B.n252 VSUBS 0.00786f
C343 B.n253 VSUBS 0.00786f
C344 B.n254 VSUBS 0.00786f
C345 B.n255 VSUBS 0.00786f
C346 B.n256 VSUBS 0.00786f
C347 B.n257 VSUBS 0.00786f
C348 B.n258 VSUBS 0.00786f
C349 B.n259 VSUBS 0.00786f
C350 B.n260 VSUBS 0.00786f
C351 B.n261 VSUBS 0.00786f
C352 B.n262 VSUBS 0.00786f
C353 B.n263 VSUBS 0.00786f
C354 B.n264 VSUBS 0.00786f
C355 B.n265 VSUBS 0.00786f
C356 B.n266 VSUBS 0.00786f
C357 B.n267 VSUBS 0.00786f
C358 B.n268 VSUBS 0.00786f
C359 B.n269 VSUBS 0.00786f
C360 B.n270 VSUBS 0.00786f
C361 B.n271 VSUBS 0.00786f
C362 B.n272 VSUBS 0.017897f
C363 B.n273 VSUBS 0.017897f
C364 B.n274 VSUBS 0.017241f
C365 B.n275 VSUBS 0.00786f
C366 B.n276 VSUBS 0.00786f
C367 B.n277 VSUBS 0.00786f
C368 B.n278 VSUBS 0.00786f
C369 B.n279 VSUBS 0.00786f
C370 B.n280 VSUBS 0.00786f
C371 B.n281 VSUBS 0.00786f
C372 B.n282 VSUBS 0.00786f
C373 B.n283 VSUBS 0.00786f
C374 B.n284 VSUBS 0.00786f
C375 B.n285 VSUBS 0.00786f
C376 B.n286 VSUBS 0.00786f
C377 B.n287 VSUBS 0.00786f
C378 B.n288 VSUBS 0.00786f
C379 B.n289 VSUBS 0.00786f
C380 B.n290 VSUBS 0.00786f
C381 B.n291 VSUBS 0.00786f
C382 B.n292 VSUBS 0.00786f
C383 B.n293 VSUBS 0.00786f
C384 B.n294 VSUBS 0.00786f
C385 B.n295 VSUBS 0.00786f
C386 B.n296 VSUBS 0.00786f
C387 B.n297 VSUBS 0.00786f
C388 B.n298 VSUBS 0.00786f
C389 B.n299 VSUBS 0.00786f
C390 B.n300 VSUBS 0.00786f
C391 B.n301 VSUBS 0.00786f
C392 B.n302 VSUBS 0.00786f
C393 B.n303 VSUBS 0.00786f
C394 B.n304 VSUBS 0.00786f
C395 B.n305 VSUBS 0.00786f
C396 B.n306 VSUBS 0.00786f
C397 B.n307 VSUBS 0.00786f
C398 B.n308 VSUBS 0.00786f
C399 B.n309 VSUBS 0.00786f
C400 B.n310 VSUBS 0.00786f
C401 B.n311 VSUBS 0.00786f
C402 B.n312 VSUBS 0.00786f
C403 B.n313 VSUBS 0.00786f
C404 B.n314 VSUBS 0.00786f
C405 B.n315 VSUBS 0.00786f
C406 B.n316 VSUBS 0.00786f
C407 B.n317 VSUBS 0.00786f
C408 B.n318 VSUBS 0.00786f
C409 B.n319 VSUBS 0.00786f
C410 B.n320 VSUBS 0.00786f
C411 B.n321 VSUBS 0.00786f
C412 B.n322 VSUBS 0.00786f
C413 B.n323 VSUBS 0.00786f
C414 B.n324 VSUBS 0.00786f
C415 B.n325 VSUBS 0.00786f
C416 B.n326 VSUBS 0.00786f
C417 B.n327 VSUBS 0.00786f
C418 B.n328 VSUBS 0.00786f
C419 B.n329 VSUBS 0.00786f
C420 B.n330 VSUBS 0.00786f
C421 B.n331 VSUBS 0.00786f
C422 B.n332 VSUBS 0.00786f
C423 B.n333 VSUBS 0.00786f
C424 B.n334 VSUBS 0.00786f
C425 B.n335 VSUBS 0.00786f
C426 B.n336 VSUBS 0.00786f
C427 B.n337 VSUBS 0.00786f
C428 B.n338 VSUBS 0.00786f
C429 B.n339 VSUBS 0.00786f
C430 B.n340 VSUBS 0.00786f
C431 B.n341 VSUBS 0.00786f
C432 B.n342 VSUBS 0.00786f
C433 B.n343 VSUBS 0.00786f
C434 B.n344 VSUBS 0.00786f
C435 B.n345 VSUBS 0.00786f
C436 B.n346 VSUBS 0.00786f
C437 B.n347 VSUBS 0.00786f
C438 B.n348 VSUBS 0.00786f
C439 B.n349 VSUBS 0.00786f
C440 B.n350 VSUBS 0.00786f
C441 B.n351 VSUBS 0.00786f
C442 B.n352 VSUBS 0.00786f
C443 B.n353 VSUBS 0.00786f
C444 B.n354 VSUBS 0.00786f
C445 B.n355 VSUBS 0.00786f
C446 B.n356 VSUBS 0.00786f
C447 B.n357 VSUBS 0.00786f
C448 B.n358 VSUBS 0.00786f
C449 B.n359 VSUBS 0.00786f
C450 B.n360 VSUBS 0.00786f
C451 B.n361 VSUBS 0.00786f
C452 B.n362 VSUBS 0.00786f
C453 B.n363 VSUBS 0.00786f
C454 B.n364 VSUBS 0.00786f
C455 B.n365 VSUBS 0.00786f
C456 B.n366 VSUBS 0.00786f
C457 B.n367 VSUBS 0.00786f
C458 B.n368 VSUBS 0.00786f
C459 B.n369 VSUBS 0.00786f
C460 B.n370 VSUBS 0.00786f
C461 B.n371 VSUBS 0.00786f
C462 B.n372 VSUBS 0.00786f
C463 B.n373 VSUBS 0.017241f
C464 B.n374 VSUBS 0.017897f
C465 B.n375 VSUBS 0.0169f
C466 B.n376 VSUBS 0.00786f
C467 B.n377 VSUBS 0.00786f
C468 B.n378 VSUBS 0.00786f
C469 B.n379 VSUBS 0.00786f
C470 B.n380 VSUBS 0.00786f
C471 B.n381 VSUBS 0.00786f
C472 B.n382 VSUBS 0.00786f
C473 B.n383 VSUBS 0.00786f
C474 B.n384 VSUBS 0.00786f
C475 B.n385 VSUBS 0.00786f
C476 B.n386 VSUBS 0.00786f
C477 B.n387 VSUBS 0.00786f
C478 B.n388 VSUBS 0.00786f
C479 B.n389 VSUBS 0.00786f
C480 B.n390 VSUBS 0.00786f
C481 B.n391 VSUBS 0.00786f
C482 B.n392 VSUBS 0.00786f
C483 B.n393 VSUBS 0.00786f
C484 B.n394 VSUBS 0.00786f
C485 B.n395 VSUBS 0.00786f
C486 B.n396 VSUBS 0.00786f
C487 B.n397 VSUBS 0.00786f
C488 B.n398 VSUBS 0.00786f
C489 B.n399 VSUBS 0.00786f
C490 B.n400 VSUBS 0.00786f
C491 B.n401 VSUBS 0.00786f
C492 B.n402 VSUBS 0.00786f
C493 B.n403 VSUBS 0.00786f
C494 B.n404 VSUBS 0.00786f
C495 B.n405 VSUBS 0.00786f
C496 B.n406 VSUBS 0.00786f
C497 B.n407 VSUBS 0.00786f
C498 B.n408 VSUBS 0.00786f
C499 B.n409 VSUBS 0.00786f
C500 B.n410 VSUBS 0.00786f
C501 B.n411 VSUBS 0.005432f
C502 B.n412 VSUBS 0.01821f
C503 B.n413 VSUBS 0.006357f
C504 B.n414 VSUBS 0.00786f
C505 B.n415 VSUBS 0.00786f
C506 B.n416 VSUBS 0.00786f
C507 B.n417 VSUBS 0.00786f
C508 B.n418 VSUBS 0.00786f
C509 B.n419 VSUBS 0.00786f
C510 B.n420 VSUBS 0.00786f
C511 B.n421 VSUBS 0.00786f
C512 B.n422 VSUBS 0.00786f
C513 B.n423 VSUBS 0.00786f
C514 B.n424 VSUBS 0.00786f
C515 B.n425 VSUBS 0.006357f
C516 B.n426 VSUBS 0.01821f
C517 B.n427 VSUBS 0.005432f
C518 B.n428 VSUBS 0.00786f
C519 B.n429 VSUBS 0.00786f
C520 B.n430 VSUBS 0.00786f
C521 B.n431 VSUBS 0.00786f
C522 B.n432 VSUBS 0.00786f
C523 B.n433 VSUBS 0.00786f
C524 B.n434 VSUBS 0.00786f
C525 B.n435 VSUBS 0.00786f
C526 B.n436 VSUBS 0.00786f
C527 B.n437 VSUBS 0.00786f
C528 B.n438 VSUBS 0.00786f
C529 B.n439 VSUBS 0.00786f
C530 B.n440 VSUBS 0.00786f
C531 B.n441 VSUBS 0.00786f
C532 B.n442 VSUBS 0.00786f
C533 B.n443 VSUBS 0.00786f
C534 B.n444 VSUBS 0.00786f
C535 B.n445 VSUBS 0.00786f
C536 B.n446 VSUBS 0.00786f
C537 B.n447 VSUBS 0.00786f
C538 B.n448 VSUBS 0.00786f
C539 B.n449 VSUBS 0.00786f
C540 B.n450 VSUBS 0.00786f
C541 B.n451 VSUBS 0.00786f
C542 B.n452 VSUBS 0.00786f
C543 B.n453 VSUBS 0.00786f
C544 B.n454 VSUBS 0.00786f
C545 B.n455 VSUBS 0.00786f
C546 B.n456 VSUBS 0.00786f
C547 B.n457 VSUBS 0.00786f
C548 B.n458 VSUBS 0.00786f
C549 B.n459 VSUBS 0.00786f
C550 B.n460 VSUBS 0.00786f
C551 B.n461 VSUBS 0.00786f
C552 B.n462 VSUBS 0.00786f
C553 B.n463 VSUBS 0.017897f
C554 B.n464 VSUBS 0.017897f
C555 B.n465 VSUBS 0.017241f
C556 B.n466 VSUBS 0.00786f
C557 B.n467 VSUBS 0.00786f
C558 B.n468 VSUBS 0.00786f
C559 B.n469 VSUBS 0.00786f
C560 B.n470 VSUBS 0.00786f
C561 B.n471 VSUBS 0.00786f
C562 B.n472 VSUBS 0.00786f
C563 B.n473 VSUBS 0.00786f
C564 B.n474 VSUBS 0.00786f
C565 B.n475 VSUBS 0.00786f
C566 B.n476 VSUBS 0.00786f
C567 B.n477 VSUBS 0.00786f
C568 B.n478 VSUBS 0.00786f
C569 B.n479 VSUBS 0.00786f
C570 B.n480 VSUBS 0.00786f
C571 B.n481 VSUBS 0.00786f
C572 B.n482 VSUBS 0.00786f
C573 B.n483 VSUBS 0.00786f
C574 B.n484 VSUBS 0.00786f
C575 B.n485 VSUBS 0.00786f
C576 B.n486 VSUBS 0.00786f
C577 B.n487 VSUBS 0.00786f
C578 B.n488 VSUBS 0.00786f
C579 B.n489 VSUBS 0.00786f
C580 B.n490 VSUBS 0.00786f
C581 B.n491 VSUBS 0.00786f
C582 B.n492 VSUBS 0.00786f
C583 B.n493 VSUBS 0.00786f
C584 B.n494 VSUBS 0.00786f
C585 B.n495 VSUBS 0.00786f
C586 B.n496 VSUBS 0.00786f
C587 B.n497 VSUBS 0.00786f
C588 B.n498 VSUBS 0.00786f
C589 B.n499 VSUBS 0.00786f
C590 B.n500 VSUBS 0.00786f
C591 B.n501 VSUBS 0.00786f
C592 B.n502 VSUBS 0.00786f
C593 B.n503 VSUBS 0.00786f
C594 B.n504 VSUBS 0.00786f
C595 B.n505 VSUBS 0.00786f
C596 B.n506 VSUBS 0.00786f
C597 B.n507 VSUBS 0.00786f
C598 B.n508 VSUBS 0.00786f
C599 B.n509 VSUBS 0.00786f
C600 B.n510 VSUBS 0.00786f
C601 B.n511 VSUBS 0.00786f
C602 B.n512 VSUBS 0.00786f
C603 B.n513 VSUBS 0.00786f
C604 B.n514 VSUBS 0.00786f
C605 B.n515 VSUBS 0.017797f
C606 VDD2.t4 VSUBS 0.974159f
C607 VDD2.t2 VSUBS 0.108286f
C608 VDD2.t0 VSUBS 0.108286f
C609 VDD2.n0 VSUBS 0.724814f
C610 VDD2.n1 VSUBS 2.29053f
C611 VDD2.t5 VSUBS 0.967064f
C612 VDD2.n2 VSUBS 2.03166f
C613 VDD2.t1 VSUBS 0.108286f
C614 VDD2.t3 VSUBS 0.108286f
C615 VDD2.n3 VSUBS 0.72479f
C616 VTAIL.t5 VSUBS 0.157596f
C617 VTAIL.t8 VSUBS 0.157596f
C618 VTAIL.n0 VSUBS 0.929209f
C619 VTAIL.n1 VSUBS 0.802052f
C620 VTAIL.t10 VSUBS 1.27746f
C621 VTAIL.n2 VSUBS 1.01722f
C622 VTAIL.t2 VSUBS 0.157596f
C623 VTAIL.t1 VSUBS 0.157596f
C624 VTAIL.n3 VSUBS 0.929209f
C625 VTAIL.n4 VSUBS 2.15398f
C626 VTAIL.t7 VSUBS 0.157596f
C627 VTAIL.t4 VSUBS 0.157596f
C628 VTAIL.n5 VSUBS 0.929215f
C629 VTAIL.n6 VSUBS 2.15398f
C630 VTAIL.t6 VSUBS 1.27747f
C631 VTAIL.n7 VSUBS 1.01722f
C632 VTAIL.t0 VSUBS 0.157596f
C633 VTAIL.t11 VSUBS 0.157596f
C634 VTAIL.n8 VSUBS 0.929215f
C635 VTAIL.n9 VSUBS 0.935664f
C636 VTAIL.t3 VSUBS 1.27746f
C637 VTAIL.n10 VSUBS 2.0494f
C638 VTAIL.t9 VSUBS 1.27746f
C639 VTAIL.n11 VSUBS 1.99689f
C640 VN.n0 VSUBS 0.044311f
C641 VN.t5 VSUBS 1.30047f
C642 VN.n1 VSUBS 0.037265f
C643 VN.t1 VSUBS 1.5078f
C644 VN.n2 VSUBS 0.585867f
C645 VN.t3 VSUBS 1.30047f
C646 VN.n3 VSUBS 0.617612f
C647 VN.n4 VSUBS 0.089482f
C648 VN.n5 VSUBS 0.326073f
C649 VN.n6 VSUBS 0.044311f
C650 VN.n7 VSUBS 0.044311f
C651 VN.n8 VSUBS 0.085209f
C652 VN.n9 VSUBS 0.049966f
C653 VN.n10 VSUBS 0.59924f
C654 VN.n11 VSUBS 0.046541f
C655 VN.n12 VSUBS 0.044311f
C656 VN.t0 VSUBS 1.30047f
C657 VN.n13 VSUBS 0.037265f
C658 VN.t2 VSUBS 1.5078f
C659 VN.n14 VSUBS 0.585867f
C660 VN.t4 VSUBS 1.30047f
C661 VN.n15 VSUBS 0.617612f
C662 VN.n16 VSUBS 0.089482f
C663 VN.n17 VSUBS 0.326073f
C664 VN.n18 VSUBS 0.044311f
C665 VN.n19 VSUBS 0.044311f
C666 VN.n20 VSUBS 0.085209f
C667 VN.n21 VSUBS 0.049966f
C668 VN.n22 VSUBS 0.59924f
C669 VN.n23 VSUBS 1.79615f
.ends

