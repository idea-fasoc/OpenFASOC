* NGSPICE file created from diff_pair_sample_1753.ext - technology: sky130A

.subckt diff_pair_sample_1753 VTAIL VN VP B VDD2 VDD1
X0 B.t19 B.t17 B.t18 B.t11 sky130_fd_pr__nfet_01v8 ad=6.3531 pd=33.36 as=0 ps=0 w=16.29 l=0.24
X1 B.t16 B.t14 B.t15 B.t7 sky130_fd_pr__nfet_01v8 ad=6.3531 pd=33.36 as=0 ps=0 w=16.29 l=0.24
X2 B.t13 B.t10 B.t12 B.t11 sky130_fd_pr__nfet_01v8 ad=6.3531 pd=33.36 as=0 ps=0 w=16.29 l=0.24
X3 VTAIL.t9 VN.t0 VDD2.t4 B.t1 sky130_fd_pr__nfet_01v8 ad=2.68785 pd=16.62 as=2.68785 ps=16.62 w=16.29 l=0.24
X4 VTAIL.t10 VP.t0 VDD1.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=2.68785 pd=16.62 as=2.68785 ps=16.62 w=16.29 l=0.24
X5 VTAIL.t11 VP.t1 VDD1.t4 B.t1 sky130_fd_pr__nfet_01v8 ad=2.68785 pd=16.62 as=2.68785 ps=16.62 w=16.29 l=0.24
X6 VDD1.t3 VP.t2 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=6.3531 pd=33.36 as=2.68785 ps=16.62 w=16.29 l=0.24
X7 VDD1.t2 VP.t3 VTAIL.t3 B.t2 sky130_fd_pr__nfet_01v8 ad=2.68785 pd=16.62 as=6.3531 ps=33.36 w=16.29 l=0.24
X8 VDD2.t3 VN.t1 VTAIL.t8 B.t4 sky130_fd_pr__nfet_01v8 ad=6.3531 pd=33.36 as=2.68785 ps=16.62 w=16.29 l=0.24
X9 VDD2.t5 VN.t2 VTAIL.t7 B.t3 sky130_fd_pr__nfet_01v8 ad=2.68785 pd=16.62 as=6.3531 ps=33.36 w=16.29 l=0.24
X10 VDD2.t1 VN.t3 VTAIL.t6 B.t2 sky130_fd_pr__nfet_01v8 ad=2.68785 pd=16.62 as=6.3531 ps=33.36 w=16.29 l=0.24
X11 VDD1.t1 VP.t4 VTAIL.t1 B.t3 sky130_fd_pr__nfet_01v8 ad=2.68785 pd=16.62 as=6.3531 ps=33.36 w=16.29 l=0.24
X12 VTAIL.t5 VN.t4 VDD2.t2 B.t5 sky130_fd_pr__nfet_01v8 ad=2.68785 pd=16.62 as=2.68785 ps=16.62 w=16.29 l=0.24
X13 B.t9 B.t6 B.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=6.3531 pd=33.36 as=0 ps=0 w=16.29 l=0.24
X14 VDD1.t0 VP.t5 VTAIL.t2 B.t4 sky130_fd_pr__nfet_01v8 ad=6.3531 pd=33.36 as=2.68785 ps=16.62 w=16.29 l=0.24
X15 VDD2.t0 VN.t5 VTAIL.t4 B.t0 sky130_fd_pr__nfet_01v8 ad=6.3531 pd=33.36 as=2.68785 ps=16.62 w=16.29 l=0.24
R0 B.n416 B.t14 1862.1
R1 B.n414 B.t6 1862.1
R2 B.n95 B.t10 1862.1
R3 B.n92 B.t17 1862.1
R4 B.n720 B.n719 585
R5 B.n326 B.n90 585
R6 B.n325 B.n324 585
R7 B.n323 B.n322 585
R8 B.n321 B.n320 585
R9 B.n319 B.n318 585
R10 B.n317 B.n316 585
R11 B.n315 B.n314 585
R12 B.n313 B.n312 585
R13 B.n311 B.n310 585
R14 B.n309 B.n308 585
R15 B.n307 B.n306 585
R16 B.n305 B.n304 585
R17 B.n303 B.n302 585
R18 B.n301 B.n300 585
R19 B.n299 B.n298 585
R20 B.n297 B.n296 585
R21 B.n295 B.n294 585
R22 B.n293 B.n292 585
R23 B.n291 B.n290 585
R24 B.n289 B.n288 585
R25 B.n287 B.n286 585
R26 B.n285 B.n284 585
R27 B.n283 B.n282 585
R28 B.n281 B.n280 585
R29 B.n279 B.n278 585
R30 B.n277 B.n276 585
R31 B.n275 B.n274 585
R32 B.n273 B.n272 585
R33 B.n271 B.n270 585
R34 B.n269 B.n268 585
R35 B.n267 B.n266 585
R36 B.n265 B.n264 585
R37 B.n263 B.n262 585
R38 B.n261 B.n260 585
R39 B.n259 B.n258 585
R40 B.n257 B.n256 585
R41 B.n255 B.n254 585
R42 B.n253 B.n252 585
R43 B.n251 B.n250 585
R44 B.n249 B.n248 585
R45 B.n247 B.n246 585
R46 B.n245 B.n244 585
R47 B.n243 B.n242 585
R48 B.n241 B.n240 585
R49 B.n239 B.n238 585
R50 B.n237 B.n236 585
R51 B.n235 B.n234 585
R52 B.n233 B.n232 585
R53 B.n231 B.n230 585
R54 B.n229 B.n228 585
R55 B.n227 B.n226 585
R56 B.n225 B.n224 585
R57 B.n223 B.n222 585
R58 B.n221 B.n220 585
R59 B.n219 B.n218 585
R60 B.n217 B.n216 585
R61 B.n215 B.n214 585
R62 B.n213 B.n212 585
R63 B.n211 B.n210 585
R64 B.n209 B.n208 585
R65 B.n207 B.n206 585
R66 B.n205 B.n204 585
R67 B.n203 B.n202 585
R68 B.n201 B.n200 585
R69 B.n199 B.n198 585
R70 B.n197 B.n196 585
R71 B.n195 B.n194 585
R72 B.n193 B.n192 585
R73 B.n191 B.n190 585
R74 B.n189 B.n188 585
R75 B.n187 B.n186 585
R76 B.n185 B.n184 585
R77 B.n183 B.n182 585
R78 B.n181 B.n180 585
R79 B.n179 B.n178 585
R80 B.n177 B.n176 585
R81 B.n175 B.n174 585
R82 B.n173 B.n172 585
R83 B.n171 B.n170 585
R84 B.n169 B.n168 585
R85 B.n167 B.n166 585
R86 B.n165 B.n164 585
R87 B.n163 B.n162 585
R88 B.n161 B.n160 585
R89 B.n159 B.n158 585
R90 B.n157 B.n156 585
R91 B.n155 B.n154 585
R92 B.n153 B.n152 585
R93 B.n151 B.n150 585
R94 B.n149 B.n148 585
R95 B.n147 B.n146 585
R96 B.n145 B.n144 585
R97 B.n143 B.n142 585
R98 B.n141 B.n140 585
R99 B.n139 B.n138 585
R100 B.n137 B.n136 585
R101 B.n135 B.n134 585
R102 B.n133 B.n132 585
R103 B.n131 B.n130 585
R104 B.n129 B.n128 585
R105 B.n127 B.n126 585
R106 B.n125 B.n124 585
R107 B.n123 B.n122 585
R108 B.n121 B.n120 585
R109 B.n119 B.n118 585
R110 B.n117 B.n116 585
R111 B.n115 B.n114 585
R112 B.n113 B.n112 585
R113 B.n111 B.n110 585
R114 B.n109 B.n108 585
R115 B.n107 B.n106 585
R116 B.n105 B.n104 585
R117 B.n103 B.n102 585
R118 B.n101 B.n100 585
R119 B.n99 B.n98 585
R120 B.n32 B.n31 585
R121 B.n725 B.n724 585
R122 B.n718 B.n91 585
R123 B.n91 B.n29 585
R124 B.n717 B.n28 585
R125 B.n729 B.n28 585
R126 B.n716 B.n27 585
R127 B.n730 B.n27 585
R128 B.n715 B.n26 585
R129 B.n731 B.n26 585
R130 B.n714 B.n713 585
R131 B.n713 B.n25 585
R132 B.n712 B.n21 585
R133 B.n737 B.n21 585
R134 B.n711 B.n20 585
R135 B.n738 B.n20 585
R136 B.n710 B.n19 585
R137 B.n739 B.n19 585
R138 B.n709 B.n708 585
R139 B.n708 B.n15 585
R140 B.n707 B.n14 585
R141 B.n745 B.n14 585
R142 B.n706 B.n13 585
R143 B.n746 B.n13 585
R144 B.n705 B.n12 585
R145 B.n747 B.n12 585
R146 B.n704 B.n703 585
R147 B.n703 B.n11 585
R148 B.n702 B.n7 585
R149 B.n753 B.n7 585
R150 B.n701 B.n6 585
R151 B.n754 B.n6 585
R152 B.n700 B.n5 585
R153 B.n755 B.n5 585
R154 B.n699 B.n698 585
R155 B.n698 B.n4 585
R156 B.n697 B.n327 585
R157 B.n697 B.n696 585
R158 B.n686 B.n328 585
R159 B.n689 B.n328 585
R160 B.n688 B.n687 585
R161 B.n690 B.n688 585
R162 B.n685 B.n332 585
R163 B.n336 B.n332 585
R164 B.n684 B.n683 585
R165 B.n683 B.n682 585
R166 B.n334 B.n333 585
R167 B.n335 B.n334 585
R168 B.n675 B.n674 585
R169 B.n676 B.n675 585
R170 B.n673 B.n341 585
R171 B.n341 B.n340 585
R172 B.n672 B.n671 585
R173 B.n671 B.n670 585
R174 B.n343 B.n342 585
R175 B.n663 B.n343 585
R176 B.n662 B.n661 585
R177 B.n664 B.n662 585
R178 B.n660 B.n348 585
R179 B.n348 B.n347 585
R180 B.n659 B.n658 585
R181 B.n658 B.n657 585
R182 B.n350 B.n349 585
R183 B.n351 B.n350 585
R184 B.n653 B.n652 585
R185 B.n354 B.n353 585
R186 B.n649 B.n648 585
R187 B.n650 B.n649 585
R188 B.n647 B.n413 585
R189 B.n646 B.n645 585
R190 B.n644 B.n643 585
R191 B.n642 B.n641 585
R192 B.n640 B.n639 585
R193 B.n638 B.n637 585
R194 B.n636 B.n635 585
R195 B.n634 B.n633 585
R196 B.n632 B.n631 585
R197 B.n630 B.n629 585
R198 B.n628 B.n627 585
R199 B.n626 B.n625 585
R200 B.n624 B.n623 585
R201 B.n622 B.n621 585
R202 B.n620 B.n619 585
R203 B.n618 B.n617 585
R204 B.n616 B.n615 585
R205 B.n614 B.n613 585
R206 B.n612 B.n611 585
R207 B.n610 B.n609 585
R208 B.n608 B.n607 585
R209 B.n606 B.n605 585
R210 B.n604 B.n603 585
R211 B.n602 B.n601 585
R212 B.n600 B.n599 585
R213 B.n598 B.n597 585
R214 B.n596 B.n595 585
R215 B.n594 B.n593 585
R216 B.n592 B.n591 585
R217 B.n590 B.n589 585
R218 B.n588 B.n587 585
R219 B.n586 B.n585 585
R220 B.n584 B.n583 585
R221 B.n582 B.n581 585
R222 B.n580 B.n579 585
R223 B.n578 B.n577 585
R224 B.n576 B.n575 585
R225 B.n574 B.n573 585
R226 B.n572 B.n571 585
R227 B.n570 B.n569 585
R228 B.n568 B.n567 585
R229 B.n566 B.n565 585
R230 B.n564 B.n563 585
R231 B.n562 B.n561 585
R232 B.n560 B.n559 585
R233 B.n558 B.n557 585
R234 B.n556 B.n555 585
R235 B.n554 B.n553 585
R236 B.n552 B.n551 585
R237 B.n550 B.n549 585
R238 B.n548 B.n547 585
R239 B.n545 B.n544 585
R240 B.n543 B.n542 585
R241 B.n541 B.n540 585
R242 B.n539 B.n538 585
R243 B.n537 B.n536 585
R244 B.n535 B.n534 585
R245 B.n533 B.n532 585
R246 B.n531 B.n530 585
R247 B.n529 B.n528 585
R248 B.n527 B.n526 585
R249 B.n524 B.n523 585
R250 B.n522 B.n521 585
R251 B.n520 B.n519 585
R252 B.n518 B.n517 585
R253 B.n516 B.n515 585
R254 B.n514 B.n513 585
R255 B.n512 B.n511 585
R256 B.n510 B.n509 585
R257 B.n508 B.n507 585
R258 B.n506 B.n505 585
R259 B.n504 B.n503 585
R260 B.n502 B.n501 585
R261 B.n500 B.n499 585
R262 B.n498 B.n497 585
R263 B.n496 B.n495 585
R264 B.n494 B.n493 585
R265 B.n492 B.n491 585
R266 B.n490 B.n489 585
R267 B.n488 B.n487 585
R268 B.n486 B.n485 585
R269 B.n484 B.n483 585
R270 B.n482 B.n481 585
R271 B.n480 B.n479 585
R272 B.n478 B.n477 585
R273 B.n476 B.n475 585
R274 B.n474 B.n473 585
R275 B.n472 B.n471 585
R276 B.n470 B.n469 585
R277 B.n468 B.n467 585
R278 B.n466 B.n465 585
R279 B.n464 B.n463 585
R280 B.n462 B.n461 585
R281 B.n460 B.n459 585
R282 B.n458 B.n457 585
R283 B.n456 B.n455 585
R284 B.n454 B.n453 585
R285 B.n452 B.n451 585
R286 B.n450 B.n449 585
R287 B.n448 B.n447 585
R288 B.n446 B.n445 585
R289 B.n444 B.n443 585
R290 B.n442 B.n441 585
R291 B.n440 B.n439 585
R292 B.n438 B.n437 585
R293 B.n436 B.n435 585
R294 B.n434 B.n433 585
R295 B.n432 B.n431 585
R296 B.n430 B.n429 585
R297 B.n428 B.n427 585
R298 B.n426 B.n425 585
R299 B.n424 B.n423 585
R300 B.n422 B.n421 585
R301 B.n420 B.n419 585
R302 B.n418 B.n412 585
R303 B.n650 B.n412 585
R304 B.n654 B.n352 585
R305 B.n352 B.n351 585
R306 B.n656 B.n655 585
R307 B.n657 B.n656 585
R308 B.n346 B.n345 585
R309 B.n347 B.n346 585
R310 B.n666 B.n665 585
R311 B.n665 B.n664 585
R312 B.n667 B.n344 585
R313 B.n663 B.n344 585
R314 B.n669 B.n668 585
R315 B.n670 B.n669 585
R316 B.n339 B.n338 585
R317 B.n340 B.n339 585
R318 B.n678 B.n677 585
R319 B.n677 B.n676 585
R320 B.n679 B.n337 585
R321 B.n337 B.n335 585
R322 B.n681 B.n680 585
R323 B.n682 B.n681 585
R324 B.n331 B.n330 585
R325 B.n336 B.n331 585
R326 B.n692 B.n691 585
R327 B.n691 B.n690 585
R328 B.n693 B.n329 585
R329 B.n689 B.n329 585
R330 B.n695 B.n694 585
R331 B.n696 B.n695 585
R332 B.n2 B.n0 585
R333 B.n4 B.n2 585
R334 B.n3 B.n1 585
R335 B.n754 B.n3 585
R336 B.n752 B.n751 585
R337 B.n753 B.n752 585
R338 B.n750 B.n8 585
R339 B.n11 B.n8 585
R340 B.n749 B.n748 585
R341 B.n748 B.n747 585
R342 B.n10 B.n9 585
R343 B.n746 B.n10 585
R344 B.n744 B.n743 585
R345 B.n745 B.n744 585
R346 B.n742 B.n16 585
R347 B.n16 B.n15 585
R348 B.n741 B.n740 585
R349 B.n740 B.n739 585
R350 B.n18 B.n17 585
R351 B.n738 B.n18 585
R352 B.n736 B.n735 585
R353 B.n737 B.n736 585
R354 B.n734 B.n22 585
R355 B.n25 B.n22 585
R356 B.n733 B.n732 585
R357 B.n732 B.n731 585
R358 B.n24 B.n23 585
R359 B.n730 B.n24 585
R360 B.n728 B.n727 585
R361 B.n729 B.n728 585
R362 B.n726 B.n30 585
R363 B.n30 B.n29 585
R364 B.n757 B.n756 585
R365 B.n756 B.n755 585
R366 B.n652 B.n352 473.281
R367 B.n724 B.n30 473.281
R368 B.n412 B.n350 473.281
R369 B.n720 B.n91 473.281
R370 B.n416 B.t16 367.409
R371 B.n92 B.t18 367.409
R372 B.n414 B.t9 367.409
R373 B.n95 B.t12 367.409
R374 B.n417 B.t15 356.356
R375 B.n93 B.t19 356.356
R376 B.n415 B.t8 356.356
R377 B.n96 B.t13 356.356
R378 B.n722 B.n721 256.663
R379 B.n722 B.n89 256.663
R380 B.n722 B.n88 256.663
R381 B.n722 B.n87 256.663
R382 B.n722 B.n86 256.663
R383 B.n722 B.n85 256.663
R384 B.n722 B.n84 256.663
R385 B.n722 B.n83 256.663
R386 B.n722 B.n82 256.663
R387 B.n722 B.n81 256.663
R388 B.n722 B.n80 256.663
R389 B.n722 B.n79 256.663
R390 B.n722 B.n78 256.663
R391 B.n722 B.n77 256.663
R392 B.n722 B.n76 256.663
R393 B.n722 B.n75 256.663
R394 B.n722 B.n74 256.663
R395 B.n722 B.n73 256.663
R396 B.n722 B.n72 256.663
R397 B.n722 B.n71 256.663
R398 B.n722 B.n70 256.663
R399 B.n722 B.n69 256.663
R400 B.n722 B.n68 256.663
R401 B.n722 B.n67 256.663
R402 B.n722 B.n66 256.663
R403 B.n722 B.n65 256.663
R404 B.n722 B.n64 256.663
R405 B.n722 B.n63 256.663
R406 B.n722 B.n62 256.663
R407 B.n722 B.n61 256.663
R408 B.n722 B.n60 256.663
R409 B.n722 B.n59 256.663
R410 B.n722 B.n58 256.663
R411 B.n722 B.n57 256.663
R412 B.n722 B.n56 256.663
R413 B.n722 B.n55 256.663
R414 B.n722 B.n54 256.663
R415 B.n722 B.n53 256.663
R416 B.n722 B.n52 256.663
R417 B.n722 B.n51 256.663
R418 B.n722 B.n50 256.663
R419 B.n722 B.n49 256.663
R420 B.n722 B.n48 256.663
R421 B.n722 B.n47 256.663
R422 B.n722 B.n46 256.663
R423 B.n722 B.n45 256.663
R424 B.n722 B.n44 256.663
R425 B.n722 B.n43 256.663
R426 B.n722 B.n42 256.663
R427 B.n722 B.n41 256.663
R428 B.n722 B.n40 256.663
R429 B.n722 B.n39 256.663
R430 B.n722 B.n38 256.663
R431 B.n722 B.n37 256.663
R432 B.n722 B.n36 256.663
R433 B.n722 B.n35 256.663
R434 B.n722 B.n34 256.663
R435 B.n722 B.n33 256.663
R436 B.n723 B.n722 256.663
R437 B.n651 B.n650 256.663
R438 B.n650 B.n355 256.663
R439 B.n650 B.n356 256.663
R440 B.n650 B.n357 256.663
R441 B.n650 B.n358 256.663
R442 B.n650 B.n359 256.663
R443 B.n650 B.n360 256.663
R444 B.n650 B.n361 256.663
R445 B.n650 B.n362 256.663
R446 B.n650 B.n363 256.663
R447 B.n650 B.n364 256.663
R448 B.n650 B.n365 256.663
R449 B.n650 B.n366 256.663
R450 B.n650 B.n367 256.663
R451 B.n650 B.n368 256.663
R452 B.n650 B.n369 256.663
R453 B.n650 B.n370 256.663
R454 B.n650 B.n371 256.663
R455 B.n650 B.n372 256.663
R456 B.n650 B.n373 256.663
R457 B.n650 B.n374 256.663
R458 B.n650 B.n375 256.663
R459 B.n650 B.n376 256.663
R460 B.n650 B.n377 256.663
R461 B.n650 B.n378 256.663
R462 B.n650 B.n379 256.663
R463 B.n650 B.n380 256.663
R464 B.n650 B.n381 256.663
R465 B.n650 B.n382 256.663
R466 B.n650 B.n383 256.663
R467 B.n650 B.n384 256.663
R468 B.n650 B.n385 256.663
R469 B.n650 B.n386 256.663
R470 B.n650 B.n387 256.663
R471 B.n650 B.n388 256.663
R472 B.n650 B.n389 256.663
R473 B.n650 B.n390 256.663
R474 B.n650 B.n391 256.663
R475 B.n650 B.n392 256.663
R476 B.n650 B.n393 256.663
R477 B.n650 B.n394 256.663
R478 B.n650 B.n395 256.663
R479 B.n650 B.n396 256.663
R480 B.n650 B.n397 256.663
R481 B.n650 B.n398 256.663
R482 B.n650 B.n399 256.663
R483 B.n650 B.n400 256.663
R484 B.n650 B.n401 256.663
R485 B.n650 B.n402 256.663
R486 B.n650 B.n403 256.663
R487 B.n650 B.n404 256.663
R488 B.n650 B.n405 256.663
R489 B.n650 B.n406 256.663
R490 B.n650 B.n407 256.663
R491 B.n650 B.n408 256.663
R492 B.n650 B.n409 256.663
R493 B.n650 B.n410 256.663
R494 B.n650 B.n411 256.663
R495 B.n656 B.n352 163.367
R496 B.n656 B.n346 163.367
R497 B.n665 B.n346 163.367
R498 B.n665 B.n344 163.367
R499 B.n669 B.n344 163.367
R500 B.n669 B.n339 163.367
R501 B.n677 B.n339 163.367
R502 B.n677 B.n337 163.367
R503 B.n681 B.n337 163.367
R504 B.n681 B.n331 163.367
R505 B.n691 B.n331 163.367
R506 B.n691 B.n329 163.367
R507 B.n695 B.n329 163.367
R508 B.n695 B.n2 163.367
R509 B.n756 B.n2 163.367
R510 B.n756 B.n3 163.367
R511 B.n752 B.n3 163.367
R512 B.n752 B.n8 163.367
R513 B.n748 B.n8 163.367
R514 B.n748 B.n10 163.367
R515 B.n744 B.n10 163.367
R516 B.n744 B.n16 163.367
R517 B.n740 B.n16 163.367
R518 B.n740 B.n18 163.367
R519 B.n736 B.n18 163.367
R520 B.n736 B.n22 163.367
R521 B.n732 B.n22 163.367
R522 B.n732 B.n24 163.367
R523 B.n728 B.n24 163.367
R524 B.n728 B.n30 163.367
R525 B.n649 B.n354 163.367
R526 B.n649 B.n413 163.367
R527 B.n645 B.n644 163.367
R528 B.n641 B.n640 163.367
R529 B.n637 B.n636 163.367
R530 B.n633 B.n632 163.367
R531 B.n629 B.n628 163.367
R532 B.n625 B.n624 163.367
R533 B.n621 B.n620 163.367
R534 B.n617 B.n616 163.367
R535 B.n613 B.n612 163.367
R536 B.n609 B.n608 163.367
R537 B.n605 B.n604 163.367
R538 B.n601 B.n600 163.367
R539 B.n597 B.n596 163.367
R540 B.n593 B.n592 163.367
R541 B.n589 B.n588 163.367
R542 B.n585 B.n584 163.367
R543 B.n581 B.n580 163.367
R544 B.n577 B.n576 163.367
R545 B.n573 B.n572 163.367
R546 B.n569 B.n568 163.367
R547 B.n565 B.n564 163.367
R548 B.n561 B.n560 163.367
R549 B.n557 B.n556 163.367
R550 B.n553 B.n552 163.367
R551 B.n549 B.n548 163.367
R552 B.n544 B.n543 163.367
R553 B.n540 B.n539 163.367
R554 B.n536 B.n535 163.367
R555 B.n532 B.n531 163.367
R556 B.n528 B.n527 163.367
R557 B.n523 B.n522 163.367
R558 B.n519 B.n518 163.367
R559 B.n515 B.n514 163.367
R560 B.n511 B.n510 163.367
R561 B.n507 B.n506 163.367
R562 B.n503 B.n502 163.367
R563 B.n499 B.n498 163.367
R564 B.n495 B.n494 163.367
R565 B.n491 B.n490 163.367
R566 B.n487 B.n486 163.367
R567 B.n483 B.n482 163.367
R568 B.n479 B.n478 163.367
R569 B.n475 B.n474 163.367
R570 B.n471 B.n470 163.367
R571 B.n467 B.n466 163.367
R572 B.n463 B.n462 163.367
R573 B.n459 B.n458 163.367
R574 B.n455 B.n454 163.367
R575 B.n451 B.n450 163.367
R576 B.n447 B.n446 163.367
R577 B.n443 B.n442 163.367
R578 B.n439 B.n438 163.367
R579 B.n435 B.n434 163.367
R580 B.n431 B.n430 163.367
R581 B.n427 B.n426 163.367
R582 B.n423 B.n422 163.367
R583 B.n419 B.n412 163.367
R584 B.n658 B.n350 163.367
R585 B.n658 B.n348 163.367
R586 B.n662 B.n348 163.367
R587 B.n662 B.n343 163.367
R588 B.n671 B.n343 163.367
R589 B.n671 B.n341 163.367
R590 B.n675 B.n341 163.367
R591 B.n675 B.n334 163.367
R592 B.n683 B.n334 163.367
R593 B.n683 B.n332 163.367
R594 B.n688 B.n332 163.367
R595 B.n688 B.n328 163.367
R596 B.n697 B.n328 163.367
R597 B.n698 B.n697 163.367
R598 B.n698 B.n5 163.367
R599 B.n6 B.n5 163.367
R600 B.n7 B.n6 163.367
R601 B.n703 B.n7 163.367
R602 B.n703 B.n12 163.367
R603 B.n13 B.n12 163.367
R604 B.n14 B.n13 163.367
R605 B.n708 B.n14 163.367
R606 B.n708 B.n19 163.367
R607 B.n20 B.n19 163.367
R608 B.n21 B.n20 163.367
R609 B.n713 B.n21 163.367
R610 B.n713 B.n26 163.367
R611 B.n27 B.n26 163.367
R612 B.n28 B.n27 163.367
R613 B.n91 B.n28 163.367
R614 B.n98 B.n32 163.367
R615 B.n102 B.n101 163.367
R616 B.n106 B.n105 163.367
R617 B.n110 B.n109 163.367
R618 B.n114 B.n113 163.367
R619 B.n118 B.n117 163.367
R620 B.n122 B.n121 163.367
R621 B.n126 B.n125 163.367
R622 B.n130 B.n129 163.367
R623 B.n134 B.n133 163.367
R624 B.n138 B.n137 163.367
R625 B.n142 B.n141 163.367
R626 B.n146 B.n145 163.367
R627 B.n150 B.n149 163.367
R628 B.n154 B.n153 163.367
R629 B.n158 B.n157 163.367
R630 B.n162 B.n161 163.367
R631 B.n166 B.n165 163.367
R632 B.n170 B.n169 163.367
R633 B.n174 B.n173 163.367
R634 B.n178 B.n177 163.367
R635 B.n182 B.n181 163.367
R636 B.n186 B.n185 163.367
R637 B.n190 B.n189 163.367
R638 B.n194 B.n193 163.367
R639 B.n198 B.n197 163.367
R640 B.n202 B.n201 163.367
R641 B.n206 B.n205 163.367
R642 B.n210 B.n209 163.367
R643 B.n214 B.n213 163.367
R644 B.n218 B.n217 163.367
R645 B.n222 B.n221 163.367
R646 B.n226 B.n225 163.367
R647 B.n230 B.n229 163.367
R648 B.n234 B.n233 163.367
R649 B.n238 B.n237 163.367
R650 B.n242 B.n241 163.367
R651 B.n246 B.n245 163.367
R652 B.n250 B.n249 163.367
R653 B.n254 B.n253 163.367
R654 B.n258 B.n257 163.367
R655 B.n262 B.n261 163.367
R656 B.n266 B.n265 163.367
R657 B.n270 B.n269 163.367
R658 B.n274 B.n273 163.367
R659 B.n278 B.n277 163.367
R660 B.n282 B.n281 163.367
R661 B.n286 B.n285 163.367
R662 B.n290 B.n289 163.367
R663 B.n294 B.n293 163.367
R664 B.n298 B.n297 163.367
R665 B.n302 B.n301 163.367
R666 B.n306 B.n305 163.367
R667 B.n310 B.n309 163.367
R668 B.n314 B.n313 163.367
R669 B.n318 B.n317 163.367
R670 B.n322 B.n321 163.367
R671 B.n324 B.n90 163.367
R672 B.n652 B.n651 71.676
R673 B.n413 B.n355 71.676
R674 B.n644 B.n356 71.676
R675 B.n640 B.n357 71.676
R676 B.n636 B.n358 71.676
R677 B.n632 B.n359 71.676
R678 B.n628 B.n360 71.676
R679 B.n624 B.n361 71.676
R680 B.n620 B.n362 71.676
R681 B.n616 B.n363 71.676
R682 B.n612 B.n364 71.676
R683 B.n608 B.n365 71.676
R684 B.n604 B.n366 71.676
R685 B.n600 B.n367 71.676
R686 B.n596 B.n368 71.676
R687 B.n592 B.n369 71.676
R688 B.n588 B.n370 71.676
R689 B.n584 B.n371 71.676
R690 B.n580 B.n372 71.676
R691 B.n576 B.n373 71.676
R692 B.n572 B.n374 71.676
R693 B.n568 B.n375 71.676
R694 B.n564 B.n376 71.676
R695 B.n560 B.n377 71.676
R696 B.n556 B.n378 71.676
R697 B.n552 B.n379 71.676
R698 B.n548 B.n380 71.676
R699 B.n543 B.n381 71.676
R700 B.n539 B.n382 71.676
R701 B.n535 B.n383 71.676
R702 B.n531 B.n384 71.676
R703 B.n527 B.n385 71.676
R704 B.n522 B.n386 71.676
R705 B.n518 B.n387 71.676
R706 B.n514 B.n388 71.676
R707 B.n510 B.n389 71.676
R708 B.n506 B.n390 71.676
R709 B.n502 B.n391 71.676
R710 B.n498 B.n392 71.676
R711 B.n494 B.n393 71.676
R712 B.n490 B.n394 71.676
R713 B.n486 B.n395 71.676
R714 B.n482 B.n396 71.676
R715 B.n478 B.n397 71.676
R716 B.n474 B.n398 71.676
R717 B.n470 B.n399 71.676
R718 B.n466 B.n400 71.676
R719 B.n462 B.n401 71.676
R720 B.n458 B.n402 71.676
R721 B.n454 B.n403 71.676
R722 B.n450 B.n404 71.676
R723 B.n446 B.n405 71.676
R724 B.n442 B.n406 71.676
R725 B.n438 B.n407 71.676
R726 B.n434 B.n408 71.676
R727 B.n430 B.n409 71.676
R728 B.n426 B.n410 71.676
R729 B.n422 B.n411 71.676
R730 B.n724 B.n723 71.676
R731 B.n98 B.n33 71.676
R732 B.n102 B.n34 71.676
R733 B.n106 B.n35 71.676
R734 B.n110 B.n36 71.676
R735 B.n114 B.n37 71.676
R736 B.n118 B.n38 71.676
R737 B.n122 B.n39 71.676
R738 B.n126 B.n40 71.676
R739 B.n130 B.n41 71.676
R740 B.n134 B.n42 71.676
R741 B.n138 B.n43 71.676
R742 B.n142 B.n44 71.676
R743 B.n146 B.n45 71.676
R744 B.n150 B.n46 71.676
R745 B.n154 B.n47 71.676
R746 B.n158 B.n48 71.676
R747 B.n162 B.n49 71.676
R748 B.n166 B.n50 71.676
R749 B.n170 B.n51 71.676
R750 B.n174 B.n52 71.676
R751 B.n178 B.n53 71.676
R752 B.n182 B.n54 71.676
R753 B.n186 B.n55 71.676
R754 B.n190 B.n56 71.676
R755 B.n194 B.n57 71.676
R756 B.n198 B.n58 71.676
R757 B.n202 B.n59 71.676
R758 B.n206 B.n60 71.676
R759 B.n210 B.n61 71.676
R760 B.n214 B.n62 71.676
R761 B.n218 B.n63 71.676
R762 B.n222 B.n64 71.676
R763 B.n226 B.n65 71.676
R764 B.n230 B.n66 71.676
R765 B.n234 B.n67 71.676
R766 B.n238 B.n68 71.676
R767 B.n242 B.n69 71.676
R768 B.n246 B.n70 71.676
R769 B.n250 B.n71 71.676
R770 B.n254 B.n72 71.676
R771 B.n258 B.n73 71.676
R772 B.n262 B.n74 71.676
R773 B.n266 B.n75 71.676
R774 B.n270 B.n76 71.676
R775 B.n274 B.n77 71.676
R776 B.n278 B.n78 71.676
R777 B.n282 B.n79 71.676
R778 B.n286 B.n80 71.676
R779 B.n290 B.n81 71.676
R780 B.n294 B.n82 71.676
R781 B.n298 B.n83 71.676
R782 B.n302 B.n84 71.676
R783 B.n306 B.n85 71.676
R784 B.n310 B.n86 71.676
R785 B.n314 B.n87 71.676
R786 B.n318 B.n88 71.676
R787 B.n322 B.n89 71.676
R788 B.n721 B.n90 71.676
R789 B.n721 B.n720 71.676
R790 B.n324 B.n89 71.676
R791 B.n321 B.n88 71.676
R792 B.n317 B.n87 71.676
R793 B.n313 B.n86 71.676
R794 B.n309 B.n85 71.676
R795 B.n305 B.n84 71.676
R796 B.n301 B.n83 71.676
R797 B.n297 B.n82 71.676
R798 B.n293 B.n81 71.676
R799 B.n289 B.n80 71.676
R800 B.n285 B.n79 71.676
R801 B.n281 B.n78 71.676
R802 B.n277 B.n77 71.676
R803 B.n273 B.n76 71.676
R804 B.n269 B.n75 71.676
R805 B.n265 B.n74 71.676
R806 B.n261 B.n73 71.676
R807 B.n257 B.n72 71.676
R808 B.n253 B.n71 71.676
R809 B.n249 B.n70 71.676
R810 B.n245 B.n69 71.676
R811 B.n241 B.n68 71.676
R812 B.n237 B.n67 71.676
R813 B.n233 B.n66 71.676
R814 B.n229 B.n65 71.676
R815 B.n225 B.n64 71.676
R816 B.n221 B.n63 71.676
R817 B.n217 B.n62 71.676
R818 B.n213 B.n61 71.676
R819 B.n209 B.n60 71.676
R820 B.n205 B.n59 71.676
R821 B.n201 B.n58 71.676
R822 B.n197 B.n57 71.676
R823 B.n193 B.n56 71.676
R824 B.n189 B.n55 71.676
R825 B.n185 B.n54 71.676
R826 B.n181 B.n53 71.676
R827 B.n177 B.n52 71.676
R828 B.n173 B.n51 71.676
R829 B.n169 B.n50 71.676
R830 B.n165 B.n49 71.676
R831 B.n161 B.n48 71.676
R832 B.n157 B.n47 71.676
R833 B.n153 B.n46 71.676
R834 B.n149 B.n45 71.676
R835 B.n145 B.n44 71.676
R836 B.n141 B.n43 71.676
R837 B.n137 B.n42 71.676
R838 B.n133 B.n41 71.676
R839 B.n129 B.n40 71.676
R840 B.n125 B.n39 71.676
R841 B.n121 B.n38 71.676
R842 B.n117 B.n37 71.676
R843 B.n113 B.n36 71.676
R844 B.n109 B.n35 71.676
R845 B.n105 B.n34 71.676
R846 B.n101 B.n33 71.676
R847 B.n723 B.n32 71.676
R848 B.n651 B.n354 71.676
R849 B.n645 B.n355 71.676
R850 B.n641 B.n356 71.676
R851 B.n637 B.n357 71.676
R852 B.n633 B.n358 71.676
R853 B.n629 B.n359 71.676
R854 B.n625 B.n360 71.676
R855 B.n621 B.n361 71.676
R856 B.n617 B.n362 71.676
R857 B.n613 B.n363 71.676
R858 B.n609 B.n364 71.676
R859 B.n605 B.n365 71.676
R860 B.n601 B.n366 71.676
R861 B.n597 B.n367 71.676
R862 B.n593 B.n368 71.676
R863 B.n589 B.n369 71.676
R864 B.n585 B.n370 71.676
R865 B.n581 B.n371 71.676
R866 B.n577 B.n372 71.676
R867 B.n573 B.n373 71.676
R868 B.n569 B.n374 71.676
R869 B.n565 B.n375 71.676
R870 B.n561 B.n376 71.676
R871 B.n557 B.n377 71.676
R872 B.n553 B.n378 71.676
R873 B.n549 B.n379 71.676
R874 B.n544 B.n380 71.676
R875 B.n540 B.n381 71.676
R876 B.n536 B.n382 71.676
R877 B.n532 B.n383 71.676
R878 B.n528 B.n384 71.676
R879 B.n523 B.n385 71.676
R880 B.n519 B.n386 71.676
R881 B.n515 B.n387 71.676
R882 B.n511 B.n388 71.676
R883 B.n507 B.n389 71.676
R884 B.n503 B.n390 71.676
R885 B.n499 B.n391 71.676
R886 B.n495 B.n392 71.676
R887 B.n491 B.n393 71.676
R888 B.n487 B.n394 71.676
R889 B.n483 B.n395 71.676
R890 B.n479 B.n396 71.676
R891 B.n475 B.n397 71.676
R892 B.n471 B.n398 71.676
R893 B.n467 B.n399 71.676
R894 B.n463 B.n400 71.676
R895 B.n459 B.n401 71.676
R896 B.n455 B.n402 71.676
R897 B.n451 B.n403 71.676
R898 B.n447 B.n404 71.676
R899 B.n443 B.n405 71.676
R900 B.n439 B.n406 71.676
R901 B.n435 B.n407 71.676
R902 B.n431 B.n408 71.676
R903 B.n427 B.n409 71.676
R904 B.n423 B.n410 71.676
R905 B.n419 B.n411 71.676
R906 B.n525 B.n417 59.5399
R907 B.n546 B.n415 59.5399
R908 B.n97 B.n96 59.5399
R909 B.n94 B.n93 59.5399
R910 B.n650 B.n351 56.62
R911 B.n722 B.n29 56.62
R912 B.n657 B.n351 34.6863
R913 B.n657 B.n347 34.6863
R914 B.n664 B.n347 34.6863
R915 B.n664 B.n663 34.6863
R916 B.n670 B.n340 34.6863
R917 B.n676 B.n340 34.6863
R918 B.n676 B.n335 34.6863
R919 B.n682 B.n335 34.6863
R920 B.n690 B.n689 34.6863
R921 B.n696 B.n4 34.6863
R922 B.n755 B.n4 34.6863
R923 B.n755 B.n754 34.6863
R924 B.n754 B.n753 34.6863
R925 B.n747 B.n11 34.6863
R926 B.n745 B.n15 34.6863
R927 B.n739 B.n15 34.6863
R928 B.n739 B.n738 34.6863
R929 B.n738 B.n737 34.6863
R930 B.n731 B.n25 34.6863
R931 B.n731 B.n730 34.6863
R932 B.n730 B.n729 34.6863
R933 B.n729 B.n29 34.6863
R934 B.n726 B.n725 30.7517
R935 B.n418 B.n349 30.7517
R936 B.n654 B.n653 30.7517
R937 B.n719 B.n718 30.7517
R938 B.n336 B.t5 30.6056
R939 B.t1 B.n746 30.6056
R940 B.t0 B.n336 27.5451
R941 B.n746 B.t2 27.5451
R942 B.n670 B.t7 23.4644
R943 B.n737 B.t11 23.4644
R944 B.n689 B.t3 19.3838
R945 B.n11 B.t4 19.3838
R946 B B.n757 18.0485
R947 B.n696 B.t3 15.3031
R948 B.n753 B.t4 15.3031
R949 B.n663 B.t7 11.2224
R950 B.n25 B.t11 11.2224
R951 B.n417 B.n416 11.055
R952 B.n415 B.n414 11.055
R953 B.n96 B.n95 11.055
R954 B.n93 B.n92 11.055
R955 B.n725 B.n31 10.6151
R956 B.n99 B.n31 10.6151
R957 B.n100 B.n99 10.6151
R958 B.n103 B.n100 10.6151
R959 B.n104 B.n103 10.6151
R960 B.n107 B.n104 10.6151
R961 B.n108 B.n107 10.6151
R962 B.n111 B.n108 10.6151
R963 B.n112 B.n111 10.6151
R964 B.n115 B.n112 10.6151
R965 B.n116 B.n115 10.6151
R966 B.n119 B.n116 10.6151
R967 B.n120 B.n119 10.6151
R968 B.n123 B.n120 10.6151
R969 B.n124 B.n123 10.6151
R970 B.n127 B.n124 10.6151
R971 B.n128 B.n127 10.6151
R972 B.n131 B.n128 10.6151
R973 B.n132 B.n131 10.6151
R974 B.n135 B.n132 10.6151
R975 B.n136 B.n135 10.6151
R976 B.n139 B.n136 10.6151
R977 B.n140 B.n139 10.6151
R978 B.n143 B.n140 10.6151
R979 B.n144 B.n143 10.6151
R980 B.n147 B.n144 10.6151
R981 B.n148 B.n147 10.6151
R982 B.n151 B.n148 10.6151
R983 B.n152 B.n151 10.6151
R984 B.n155 B.n152 10.6151
R985 B.n156 B.n155 10.6151
R986 B.n159 B.n156 10.6151
R987 B.n160 B.n159 10.6151
R988 B.n163 B.n160 10.6151
R989 B.n164 B.n163 10.6151
R990 B.n167 B.n164 10.6151
R991 B.n168 B.n167 10.6151
R992 B.n171 B.n168 10.6151
R993 B.n172 B.n171 10.6151
R994 B.n175 B.n172 10.6151
R995 B.n176 B.n175 10.6151
R996 B.n179 B.n176 10.6151
R997 B.n180 B.n179 10.6151
R998 B.n183 B.n180 10.6151
R999 B.n184 B.n183 10.6151
R1000 B.n187 B.n184 10.6151
R1001 B.n188 B.n187 10.6151
R1002 B.n191 B.n188 10.6151
R1003 B.n192 B.n191 10.6151
R1004 B.n195 B.n192 10.6151
R1005 B.n196 B.n195 10.6151
R1006 B.n199 B.n196 10.6151
R1007 B.n200 B.n199 10.6151
R1008 B.n204 B.n203 10.6151
R1009 B.n207 B.n204 10.6151
R1010 B.n208 B.n207 10.6151
R1011 B.n211 B.n208 10.6151
R1012 B.n212 B.n211 10.6151
R1013 B.n215 B.n212 10.6151
R1014 B.n216 B.n215 10.6151
R1015 B.n219 B.n216 10.6151
R1016 B.n220 B.n219 10.6151
R1017 B.n224 B.n223 10.6151
R1018 B.n227 B.n224 10.6151
R1019 B.n228 B.n227 10.6151
R1020 B.n231 B.n228 10.6151
R1021 B.n232 B.n231 10.6151
R1022 B.n235 B.n232 10.6151
R1023 B.n236 B.n235 10.6151
R1024 B.n239 B.n236 10.6151
R1025 B.n240 B.n239 10.6151
R1026 B.n243 B.n240 10.6151
R1027 B.n244 B.n243 10.6151
R1028 B.n247 B.n244 10.6151
R1029 B.n248 B.n247 10.6151
R1030 B.n251 B.n248 10.6151
R1031 B.n252 B.n251 10.6151
R1032 B.n255 B.n252 10.6151
R1033 B.n256 B.n255 10.6151
R1034 B.n259 B.n256 10.6151
R1035 B.n260 B.n259 10.6151
R1036 B.n263 B.n260 10.6151
R1037 B.n264 B.n263 10.6151
R1038 B.n267 B.n264 10.6151
R1039 B.n268 B.n267 10.6151
R1040 B.n271 B.n268 10.6151
R1041 B.n272 B.n271 10.6151
R1042 B.n275 B.n272 10.6151
R1043 B.n276 B.n275 10.6151
R1044 B.n279 B.n276 10.6151
R1045 B.n280 B.n279 10.6151
R1046 B.n283 B.n280 10.6151
R1047 B.n284 B.n283 10.6151
R1048 B.n287 B.n284 10.6151
R1049 B.n288 B.n287 10.6151
R1050 B.n291 B.n288 10.6151
R1051 B.n292 B.n291 10.6151
R1052 B.n295 B.n292 10.6151
R1053 B.n296 B.n295 10.6151
R1054 B.n299 B.n296 10.6151
R1055 B.n300 B.n299 10.6151
R1056 B.n303 B.n300 10.6151
R1057 B.n304 B.n303 10.6151
R1058 B.n307 B.n304 10.6151
R1059 B.n308 B.n307 10.6151
R1060 B.n311 B.n308 10.6151
R1061 B.n312 B.n311 10.6151
R1062 B.n315 B.n312 10.6151
R1063 B.n316 B.n315 10.6151
R1064 B.n319 B.n316 10.6151
R1065 B.n320 B.n319 10.6151
R1066 B.n323 B.n320 10.6151
R1067 B.n325 B.n323 10.6151
R1068 B.n326 B.n325 10.6151
R1069 B.n719 B.n326 10.6151
R1070 B.n659 B.n349 10.6151
R1071 B.n660 B.n659 10.6151
R1072 B.n661 B.n660 10.6151
R1073 B.n661 B.n342 10.6151
R1074 B.n672 B.n342 10.6151
R1075 B.n673 B.n672 10.6151
R1076 B.n674 B.n673 10.6151
R1077 B.n674 B.n333 10.6151
R1078 B.n684 B.n333 10.6151
R1079 B.n685 B.n684 10.6151
R1080 B.n687 B.n685 10.6151
R1081 B.n687 B.n686 10.6151
R1082 B.n686 B.n327 10.6151
R1083 B.n699 B.n327 10.6151
R1084 B.n700 B.n699 10.6151
R1085 B.n701 B.n700 10.6151
R1086 B.n702 B.n701 10.6151
R1087 B.n704 B.n702 10.6151
R1088 B.n705 B.n704 10.6151
R1089 B.n706 B.n705 10.6151
R1090 B.n707 B.n706 10.6151
R1091 B.n709 B.n707 10.6151
R1092 B.n710 B.n709 10.6151
R1093 B.n711 B.n710 10.6151
R1094 B.n712 B.n711 10.6151
R1095 B.n714 B.n712 10.6151
R1096 B.n715 B.n714 10.6151
R1097 B.n716 B.n715 10.6151
R1098 B.n717 B.n716 10.6151
R1099 B.n718 B.n717 10.6151
R1100 B.n653 B.n353 10.6151
R1101 B.n648 B.n353 10.6151
R1102 B.n648 B.n647 10.6151
R1103 B.n647 B.n646 10.6151
R1104 B.n646 B.n643 10.6151
R1105 B.n643 B.n642 10.6151
R1106 B.n642 B.n639 10.6151
R1107 B.n639 B.n638 10.6151
R1108 B.n638 B.n635 10.6151
R1109 B.n635 B.n634 10.6151
R1110 B.n634 B.n631 10.6151
R1111 B.n631 B.n630 10.6151
R1112 B.n630 B.n627 10.6151
R1113 B.n627 B.n626 10.6151
R1114 B.n626 B.n623 10.6151
R1115 B.n623 B.n622 10.6151
R1116 B.n622 B.n619 10.6151
R1117 B.n619 B.n618 10.6151
R1118 B.n618 B.n615 10.6151
R1119 B.n615 B.n614 10.6151
R1120 B.n614 B.n611 10.6151
R1121 B.n611 B.n610 10.6151
R1122 B.n610 B.n607 10.6151
R1123 B.n607 B.n606 10.6151
R1124 B.n606 B.n603 10.6151
R1125 B.n603 B.n602 10.6151
R1126 B.n602 B.n599 10.6151
R1127 B.n599 B.n598 10.6151
R1128 B.n598 B.n595 10.6151
R1129 B.n595 B.n594 10.6151
R1130 B.n594 B.n591 10.6151
R1131 B.n591 B.n590 10.6151
R1132 B.n590 B.n587 10.6151
R1133 B.n587 B.n586 10.6151
R1134 B.n586 B.n583 10.6151
R1135 B.n583 B.n582 10.6151
R1136 B.n582 B.n579 10.6151
R1137 B.n579 B.n578 10.6151
R1138 B.n578 B.n575 10.6151
R1139 B.n575 B.n574 10.6151
R1140 B.n574 B.n571 10.6151
R1141 B.n571 B.n570 10.6151
R1142 B.n570 B.n567 10.6151
R1143 B.n567 B.n566 10.6151
R1144 B.n566 B.n563 10.6151
R1145 B.n563 B.n562 10.6151
R1146 B.n562 B.n559 10.6151
R1147 B.n559 B.n558 10.6151
R1148 B.n558 B.n555 10.6151
R1149 B.n555 B.n554 10.6151
R1150 B.n554 B.n551 10.6151
R1151 B.n551 B.n550 10.6151
R1152 B.n550 B.n547 10.6151
R1153 B.n545 B.n542 10.6151
R1154 B.n542 B.n541 10.6151
R1155 B.n541 B.n538 10.6151
R1156 B.n538 B.n537 10.6151
R1157 B.n537 B.n534 10.6151
R1158 B.n534 B.n533 10.6151
R1159 B.n533 B.n530 10.6151
R1160 B.n530 B.n529 10.6151
R1161 B.n529 B.n526 10.6151
R1162 B.n524 B.n521 10.6151
R1163 B.n521 B.n520 10.6151
R1164 B.n520 B.n517 10.6151
R1165 B.n517 B.n516 10.6151
R1166 B.n516 B.n513 10.6151
R1167 B.n513 B.n512 10.6151
R1168 B.n512 B.n509 10.6151
R1169 B.n509 B.n508 10.6151
R1170 B.n508 B.n505 10.6151
R1171 B.n505 B.n504 10.6151
R1172 B.n504 B.n501 10.6151
R1173 B.n501 B.n500 10.6151
R1174 B.n500 B.n497 10.6151
R1175 B.n497 B.n496 10.6151
R1176 B.n496 B.n493 10.6151
R1177 B.n493 B.n492 10.6151
R1178 B.n492 B.n489 10.6151
R1179 B.n489 B.n488 10.6151
R1180 B.n488 B.n485 10.6151
R1181 B.n485 B.n484 10.6151
R1182 B.n484 B.n481 10.6151
R1183 B.n481 B.n480 10.6151
R1184 B.n480 B.n477 10.6151
R1185 B.n477 B.n476 10.6151
R1186 B.n476 B.n473 10.6151
R1187 B.n473 B.n472 10.6151
R1188 B.n472 B.n469 10.6151
R1189 B.n469 B.n468 10.6151
R1190 B.n468 B.n465 10.6151
R1191 B.n465 B.n464 10.6151
R1192 B.n464 B.n461 10.6151
R1193 B.n461 B.n460 10.6151
R1194 B.n460 B.n457 10.6151
R1195 B.n457 B.n456 10.6151
R1196 B.n456 B.n453 10.6151
R1197 B.n453 B.n452 10.6151
R1198 B.n452 B.n449 10.6151
R1199 B.n449 B.n448 10.6151
R1200 B.n448 B.n445 10.6151
R1201 B.n445 B.n444 10.6151
R1202 B.n444 B.n441 10.6151
R1203 B.n441 B.n440 10.6151
R1204 B.n440 B.n437 10.6151
R1205 B.n437 B.n436 10.6151
R1206 B.n436 B.n433 10.6151
R1207 B.n433 B.n432 10.6151
R1208 B.n432 B.n429 10.6151
R1209 B.n429 B.n428 10.6151
R1210 B.n428 B.n425 10.6151
R1211 B.n425 B.n424 10.6151
R1212 B.n424 B.n421 10.6151
R1213 B.n421 B.n420 10.6151
R1214 B.n420 B.n418 10.6151
R1215 B.n655 B.n654 10.6151
R1216 B.n655 B.n345 10.6151
R1217 B.n666 B.n345 10.6151
R1218 B.n667 B.n666 10.6151
R1219 B.n668 B.n667 10.6151
R1220 B.n668 B.n338 10.6151
R1221 B.n678 B.n338 10.6151
R1222 B.n679 B.n678 10.6151
R1223 B.n680 B.n679 10.6151
R1224 B.n680 B.n330 10.6151
R1225 B.n692 B.n330 10.6151
R1226 B.n693 B.n692 10.6151
R1227 B.n694 B.n693 10.6151
R1228 B.n694 B.n0 10.6151
R1229 B.n751 B.n1 10.6151
R1230 B.n751 B.n750 10.6151
R1231 B.n750 B.n749 10.6151
R1232 B.n749 B.n9 10.6151
R1233 B.n743 B.n9 10.6151
R1234 B.n743 B.n742 10.6151
R1235 B.n742 B.n741 10.6151
R1236 B.n741 B.n17 10.6151
R1237 B.n735 B.n17 10.6151
R1238 B.n735 B.n734 10.6151
R1239 B.n734 B.n733 10.6151
R1240 B.n733 B.n23 10.6151
R1241 B.n727 B.n23 10.6151
R1242 B.n727 B.n726 10.6151
R1243 B.n200 B.n97 9.36635
R1244 B.n223 B.n94 9.36635
R1245 B.n547 B.n546 9.36635
R1246 B.n525 B.n524 9.36635
R1247 B.n682 B.t0 7.1417
R1248 B.t2 B.n745 7.1417
R1249 B.n690 B.t5 4.08119
R1250 B.n747 B.t1 4.08119
R1251 B.n757 B.n0 2.81026
R1252 B.n757 B.n1 2.81026
R1253 B.n203 B.n97 1.24928
R1254 B.n220 B.n94 1.24928
R1255 B.n546 B.n545 1.24928
R1256 B.n526 B.n525 1.24928
R1257 VN.n2 VN.t3 1814.07
R1258 VN.n0 VN.t1 1814.07
R1259 VN.n6 VN.t5 1814.07
R1260 VN.n4 VN.t2 1814.07
R1261 VN.n1 VN.t0 1767.33
R1262 VN.n5 VN.t4 1767.33
R1263 VN.n7 VN.n4 161.489
R1264 VN.n3 VN.n0 161.489
R1265 VN.n3 VN.n2 161.3
R1266 VN.n7 VN.n6 161.3
R1267 VN VN.n7 43.135
R1268 VN.n1 VN.n0 36.5157
R1269 VN.n2 VN.n1 36.5157
R1270 VN.n6 VN.n5 36.5157
R1271 VN.n5 VN.n4 36.5157
R1272 VN VN.n3 0.0516364
R1273 VDD2.n175 VDD2.n91 289.615
R1274 VDD2.n84 VDD2.n0 289.615
R1275 VDD2.n176 VDD2.n175 185
R1276 VDD2.n174 VDD2.n173 185
R1277 VDD2.n95 VDD2.n94 185
R1278 VDD2.n168 VDD2.n167 185
R1279 VDD2.n166 VDD2.n97 185
R1280 VDD2.n165 VDD2.n164 185
R1281 VDD2.n100 VDD2.n98 185
R1282 VDD2.n159 VDD2.n158 185
R1283 VDD2.n157 VDD2.n156 185
R1284 VDD2.n104 VDD2.n103 185
R1285 VDD2.n151 VDD2.n150 185
R1286 VDD2.n149 VDD2.n148 185
R1287 VDD2.n108 VDD2.n107 185
R1288 VDD2.n143 VDD2.n142 185
R1289 VDD2.n141 VDD2.n140 185
R1290 VDD2.n112 VDD2.n111 185
R1291 VDD2.n135 VDD2.n134 185
R1292 VDD2.n133 VDD2.n132 185
R1293 VDD2.n116 VDD2.n115 185
R1294 VDD2.n127 VDD2.n126 185
R1295 VDD2.n125 VDD2.n124 185
R1296 VDD2.n120 VDD2.n119 185
R1297 VDD2.n28 VDD2.n27 185
R1298 VDD2.n33 VDD2.n32 185
R1299 VDD2.n35 VDD2.n34 185
R1300 VDD2.n24 VDD2.n23 185
R1301 VDD2.n41 VDD2.n40 185
R1302 VDD2.n43 VDD2.n42 185
R1303 VDD2.n20 VDD2.n19 185
R1304 VDD2.n49 VDD2.n48 185
R1305 VDD2.n51 VDD2.n50 185
R1306 VDD2.n16 VDD2.n15 185
R1307 VDD2.n57 VDD2.n56 185
R1308 VDD2.n59 VDD2.n58 185
R1309 VDD2.n12 VDD2.n11 185
R1310 VDD2.n65 VDD2.n64 185
R1311 VDD2.n67 VDD2.n66 185
R1312 VDD2.n8 VDD2.n7 185
R1313 VDD2.n74 VDD2.n73 185
R1314 VDD2.n75 VDD2.n6 185
R1315 VDD2.n77 VDD2.n76 185
R1316 VDD2.n4 VDD2.n3 185
R1317 VDD2.n83 VDD2.n82 185
R1318 VDD2.n85 VDD2.n84 185
R1319 VDD2.n121 VDD2.t0 147.659
R1320 VDD2.n29 VDD2.t3 147.659
R1321 VDD2.n175 VDD2.n174 104.615
R1322 VDD2.n174 VDD2.n94 104.615
R1323 VDD2.n167 VDD2.n94 104.615
R1324 VDD2.n167 VDD2.n166 104.615
R1325 VDD2.n166 VDD2.n165 104.615
R1326 VDD2.n165 VDD2.n98 104.615
R1327 VDD2.n158 VDD2.n98 104.615
R1328 VDD2.n158 VDD2.n157 104.615
R1329 VDD2.n157 VDD2.n103 104.615
R1330 VDD2.n150 VDD2.n103 104.615
R1331 VDD2.n150 VDD2.n149 104.615
R1332 VDD2.n149 VDD2.n107 104.615
R1333 VDD2.n142 VDD2.n107 104.615
R1334 VDD2.n142 VDD2.n141 104.615
R1335 VDD2.n141 VDD2.n111 104.615
R1336 VDD2.n134 VDD2.n111 104.615
R1337 VDD2.n134 VDD2.n133 104.615
R1338 VDD2.n133 VDD2.n115 104.615
R1339 VDD2.n126 VDD2.n115 104.615
R1340 VDD2.n126 VDD2.n125 104.615
R1341 VDD2.n125 VDD2.n119 104.615
R1342 VDD2.n33 VDD2.n27 104.615
R1343 VDD2.n34 VDD2.n33 104.615
R1344 VDD2.n34 VDD2.n23 104.615
R1345 VDD2.n41 VDD2.n23 104.615
R1346 VDD2.n42 VDD2.n41 104.615
R1347 VDD2.n42 VDD2.n19 104.615
R1348 VDD2.n49 VDD2.n19 104.615
R1349 VDD2.n50 VDD2.n49 104.615
R1350 VDD2.n50 VDD2.n15 104.615
R1351 VDD2.n57 VDD2.n15 104.615
R1352 VDD2.n58 VDD2.n57 104.615
R1353 VDD2.n58 VDD2.n11 104.615
R1354 VDD2.n65 VDD2.n11 104.615
R1355 VDD2.n66 VDD2.n65 104.615
R1356 VDD2.n66 VDD2.n7 104.615
R1357 VDD2.n74 VDD2.n7 104.615
R1358 VDD2.n75 VDD2.n74 104.615
R1359 VDD2.n76 VDD2.n75 104.615
R1360 VDD2.n76 VDD2.n3 104.615
R1361 VDD2.n83 VDD2.n3 104.615
R1362 VDD2.n84 VDD2.n83 104.615
R1363 VDD2.n90 VDD2.n89 64.9178
R1364 VDD2 VDD2.n181 64.9149
R1365 VDD2.n90 VDD2.n88 53.25
R1366 VDD2.n180 VDD2.n179 52.9369
R1367 VDD2.t0 VDD2.n119 52.3082
R1368 VDD2.t3 VDD2.n27 52.3082
R1369 VDD2.n180 VDD2.n90 39.3554
R1370 VDD2.n121 VDD2.n120 15.6677
R1371 VDD2.n29 VDD2.n28 15.6677
R1372 VDD2.n168 VDD2.n97 13.1884
R1373 VDD2.n77 VDD2.n6 13.1884
R1374 VDD2.n169 VDD2.n95 12.8005
R1375 VDD2.n164 VDD2.n99 12.8005
R1376 VDD2.n124 VDD2.n123 12.8005
R1377 VDD2.n32 VDD2.n31 12.8005
R1378 VDD2.n73 VDD2.n72 12.8005
R1379 VDD2.n78 VDD2.n4 12.8005
R1380 VDD2.n173 VDD2.n172 12.0247
R1381 VDD2.n163 VDD2.n100 12.0247
R1382 VDD2.n127 VDD2.n118 12.0247
R1383 VDD2.n35 VDD2.n26 12.0247
R1384 VDD2.n71 VDD2.n8 12.0247
R1385 VDD2.n82 VDD2.n81 12.0247
R1386 VDD2.n176 VDD2.n93 11.249
R1387 VDD2.n160 VDD2.n159 11.249
R1388 VDD2.n128 VDD2.n116 11.249
R1389 VDD2.n36 VDD2.n24 11.249
R1390 VDD2.n68 VDD2.n67 11.249
R1391 VDD2.n85 VDD2.n2 11.249
R1392 VDD2.n177 VDD2.n91 10.4732
R1393 VDD2.n156 VDD2.n102 10.4732
R1394 VDD2.n132 VDD2.n131 10.4732
R1395 VDD2.n40 VDD2.n39 10.4732
R1396 VDD2.n64 VDD2.n10 10.4732
R1397 VDD2.n86 VDD2.n0 10.4732
R1398 VDD2.n155 VDD2.n104 9.69747
R1399 VDD2.n135 VDD2.n114 9.69747
R1400 VDD2.n43 VDD2.n22 9.69747
R1401 VDD2.n63 VDD2.n12 9.69747
R1402 VDD2.n179 VDD2.n178 9.45567
R1403 VDD2.n88 VDD2.n87 9.45567
R1404 VDD2.n147 VDD2.n146 9.3005
R1405 VDD2.n106 VDD2.n105 9.3005
R1406 VDD2.n153 VDD2.n152 9.3005
R1407 VDD2.n155 VDD2.n154 9.3005
R1408 VDD2.n102 VDD2.n101 9.3005
R1409 VDD2.n161 VDD2.n160 9.3005
R1410 VDD2.n163 VDD2.n162 9.3005
R1411 VDD2.n99 VDD2.n96 9.3005
R1412 VDD2.n178 VDD2.n177 9.3005
R1413 VDD2.n93 VDD2.n92 9.3005
R1414 VDD2.n172 VDD2.n171 9.3005
R1415 VDD2.n170 VDD2.n169 9.3005
R1416 VDD2.n145 VDD2.n144 9.3005
R1417 VDD2.n110 VDD2.n109 9.3005
R1418 VDD2.n139 VDD2.n138 9.3005
R1419 VDD2.n137 VDD2.n136 9.3005
R1420 VDD2.n114 VDD2.n113 9.3005
R1421 VDD2.n131 VDD2.n130 9.3005
R1422 VDD2.n129 VDD2.n128 9.3005
R1423 VDD2.n118 VDD2.n117 9.3005
R1424 VDD2.n123 VDD2.n122 9.3005
R1425 VDD2.n87 VDD2.n86 9.3005
R1426 VDD2.n2 VDD2.n1 9.3005
R1427 VDD2.n81 VDD2.n80 9.3005
R1428 VDD2.n79 VDD2.n78 9.3005
R1429 VDD2.n18 VDD2.n17 9.3005
R1430 VDD2.n47 VDD2.n46 9.3005
R1431 VDD2.n45 VDD2.n44 9.3005
R1432 VDD2.n22 VDD2.n21 9.3005
R1433 VDD2.n39 VDD2.n38 9.3005
R1434 VDD2.n37 VDD2.n36 9.3005
R1435 VDD2.n26 VDD2.n25 9.3005
R1436 VDD2.n31 VDD2.n30 9.3005
R1437 VDD2.n53 VDD2.n52 9.3005
R1438 VDD2.n55 VDD2.n54 9.3005
R1439 VDD2.n14 VDD2.n13 9.3005
R1440 VDD2.n61 VDD2.n60 9.3005
R1441 VDD2.n63 VDD2.n62 9.3005
R1442 VDD2.n10 VDD2.n9 9.3005
R1443 VDD2.n69 VDD2.n68 9.3005
R1444 VDD2.n71 VDD2.n70 9.3005
R1445 VDD2.n72 VDD2.n5 9.3005
R1446 VDD2.n152 VDD2.n151 8.92171
R1447 VDD2.n136 VDD2.n112 8.92171
R1448 VDD2.n44 VDD2.n20 8.92171
R1449 VDD2.n60 VDD2.n59 8.92171
R1450 VDD2.n148 VDD2.n106 8.14595
R1451 VDD2.n140 VDD2.n139 8.14595
R1452 VDD2.n48 VDD2.n47 8.14595
R1453 VDD2.n56 VDD2.n14 8.14595
R1454 VDD2.n147 VDD2.n108 7.3702
R1455 VDD2.n143 VDD2.n110 7.3702
R1456 VDD2.n51 VDD2.n18 7.3702
R1457 VDD2.n55 VDD2.n16 7.3702
R1458 VDD2.n144 VDD2.n108 6.59444
R1459 VDD2.n144 VDD2.n143 6.59444
R1460 VDD2.n52 VDD2.n51 6.59444
R1461 VDD2.n52 VDD2.n16 6.59444
R1462 VDD2.n148 VDD2.n147 5.81868
R1463 VDD2.n140 VDD2.n110 5.81868
R1464 VDD2.n48 VDD2.n18 5.81868
R1465 VDD2.n56 VDD2.n55 5.81868
R1466 VDD2.n151 VDD2.n106 5.04292
R1467 VDD2.n139 VDD2.n112 5.04292
R1468 VDD2.n47 VDD2.n20 5.04292
R1469 VDD2.n59 VDD2.n14 5.04292
R1470 VDD2.n122 VDD2.n121 4.38563
R1471 VDD2.n30 VDD2.n29 4.38563
R1472 VDD2.n152 VDD2.n104 4.26717
R1473 VDD2.n136 VDD2.n135 4.26717
R1474 VDD2.n44 VDD2.n43 4.26717
R1475 VDD2.n60 VDD2.n12 4.26717
R1476 VDD2.n179 VDD2.n91 3.49141
R1477 VDD2.n156 VDD2.n155 3.49141
R1478 VDD2.n132 VDD2.n114 3.49141
R1479 VDD2.n40 VDD2.n22 3.49141
R1480 VDD2.n64 VDD2.n63 3.49141
R1481 VDD2.n88 VDD2.n0 3.49141
R1482 VDD2.n177 VDD2.n176 2.71565
R1483 VDD2.n159 VDD2.n102 2.71565
R1484 VDD2.n131 VDD2.n116 2.71565
R1485 VDD2.n39 VDD2.n24 2.71565
R1486 VDD2.n67 VDD2.n10 2.71565
R1487 VDD2.n86 VDD2.n85 2.71565
R1488 VDD2.n173 VDD2.n93 1.93989
R1489 VDD2.n160 VDD2.n100 1.93989
R1490 VDD2.n128 VDD2.n127 1.93989
R1491 VDD2.n36 VDD2.n35 1.93989
R1492 VDD2.n68 VDD2.n8 1.93989
R1493 VDD2.n82 VDD2.n2 1.93989
R1494 VDD2.n181 VDD2.t2 1.21597
R1495 VDD2.n181 VDD2.t5 1.21597
R1496 VDD2.n89 VDD2.t4 1.21597
R1497 VDD2.n89 VDD2.t1 1.21597
R1498 VDD2.n172 VDD2.n95 1.16414
R1499 VDD2.n164 VDD2.n163 1.16414
R1500 VDD2.n124 VDD2.n118 1.16414
R1501 VDD2.n32 VDD2.n26 1.16414
R1502 VDD2.n73 VDD2.n71 1.16414
R1503 VDD2.n81 VDD2.n4 1.16414
R1504 VDD2 VDD2.n180 0.427224
R1505 VDD2.n169 VDD2.n168 0.388379
R1506 VDD2.n99 VDD2.n97 0.388379
R1507 VDD2.n123 VDD2.n120 0.388379
R1508 VDD2.n31 VDD2.n28 0.388379
R1509 VDD2.n72 VDD2.n6 0.388379
R1510 VDD2.n78 VDD2.n77 0.388379
R1511 VDD2.n178 VDD2.n92 0.155672
R1512 VDD2.n171 VDD2.n92 0.155672
R1513 VDD2.n171 VDD2.n170 0.155672
R1514 VDD2.n170 VDD2.n96 0.155672
R1515 VDD2.n162 VDD2.n96 0.155672
R1516 VDD2.n162 VDD2.n161 0.155672
R1517 VDD2.n161 VDD2.n101 0.155672
R1518 VDD2.n154 VDD2.n101 0.155672
R1519 VDD2.n154 VDD2.n153 0.155672
R1520 VDD2.n153 VDD2.n105 0.155672
R1521 VDD2.n146 VDD2.n105 0.155672
R1522 VDD2.n146 VDD2.n145 0.155672
R1523 VDD2.n145 VDD2.n109 0.155672
R1524 VDD2.n138 VDD2.n109 0.155672
R1525 VDD2.n138 VDD2.n137 0.155672
R1526 VDD2.n137 VDD2.n113 0.155672
R1527 VDD2.n130 VDD2.n113 0.155672
R1528 VDD2.n130 VDD2.n129 0.155672
R1529 VDD2.n129 VDD2.n117 0.155672
R1530 VDD2.n122 VDD2.n117 0.155672
R1531 VDD2.n30 VDD2.n25 0.155672
R1532 VDD2.n37 VDD2.n25 0.155672
R1533 VDD2.n38 VDD2.n37 0.155672
R1534 VDD2.n38 VDD2.n21 0.155672
R1535 VDD2.n45 VDD2.n21 0.155672
R1536 VDD2.n46 VDD2.n45 0.155672
R1537 VDD2.n46 VDD2.n17 0.155672
R1538 VDD2.n53 VDD2.n17 0.155672
R1539 VDD2.n54 VDD2.n53 0.155672
R1540 VDD2.n54 VDD2.n13 0.155672
R1541 VDD2.n61 VDD2.n13 0.155672
R1542 VDD2.n62 VDD2.n61 0.155672
R1543 VDD2.n62 VDD2.n9 0.155672
R1544 VDD2.n69 VDD2.n9 0.155672
R1545 VDD2.n70 VDD2.n69 0.155672
R1546 VDD2.n70 VDD2.n5 0.155672
R1547 VDD2.n79 VDD2.n5 0.155672
R1548 VDD2.n80 VDD2.n79 0.155672
R1549 VDD2.n80 VDD2.n1 0.155672
R1550 VDD2.n87 VDD2.n1 0.155672
R1551 VTAIL.n362 VTAIL.n278 289.615
R1552 VTAIL.n86 VTAIL.n2 289.615
R1553 VTAIL.n272 VTAIL.n188 289.615
R1554 VTAIL.n180 VTAIL.n96 289.615
R1555 VTAIL.n306 VTAIL.n305 185
R1556 VTAIL.n311 VTAIL.n310 185
R1557 VTAIL.n313 VTAIL.n312 185
R1558 VTAIL.n302 VTAIL.n301 185
R1559 VTAIL.n319 VTAIL.n318 185
R1560 VTAIL.n321 VTAIL.n320 185
R1561 VTAIL.n298 VTAIL.n297 185
R1562 VTAIL.n327 VTAIL.n326 185
R1563 VTAIL.n329 VTAIL.n328 185
R1564 VTAIL.n294 VTAIL.n293 185
R1565 VTAIL.n335 VTAIL.n334 185
R1566 VTAIL.n337 VTAIL.n336 185
R1567 VTAIL.n290 VTAIL.n289 185
R1568 VTAIL.n343 VTAIL.n342 185
R1569 VTAIL.n345 VTAIL.n344 185
R1570 VTAIL.n286 VTAIL.n285 185
R1571 VTAIL.n352 VTAIL.n351 185
R1572 VTAIL.n353 VTAIL.n284 185
R1573 VTAIL.n355 VTAIL.n354 185
R1574 VTAIL.n282 VTAIL.n281 185
R1575 VTAIL.n361 VTAIL.n360 185
R1576 VTAIL.n363 VTAIL.n362 185
R1577 VTAIL.n30 VTAIL.n29 185
R1578 VTAIL.n35 VTAIL.n34 185
R1579 VTAIL.n37 VTAIL.n36 185
R1580 VTAIL.n26 VTAIL.n25 185
R1581 VTAIL.n43 VTAIL.n42 185
R1582 VTAIL.n45 VTAIL.n44 185
R1583 VTAIL.n22 VTAIL.n21 185
R1584 VTAIL.n51 VTAIL.n50 185
R1585 VTAIL.n53 VTAIL.n52 185
R1586 VTAIL.n18 VTAIL.n17 185
R1587 VTAIL.n59 VTAIL.n58 185
R1588 VTAIL.n61 VTAIL.n60 185
R1589 VTAIL.n14 VTAIL.n13 185
R1590 VTAIL.n67 VTAIL.n66 185
R1591 VTAIL.n69 VTAIL.n68 185
R1592 VTAIL.n10 VTAIL.n9 185
R1593 VTAIL.n76 VTAIL.n75 185
R1594 VTAIL.n77 VTAIL.n8 185
R1595 VTAIL.n79 VTAIL.n78 185
R1596 VTAIL.n6 VTAIL.n5 185
R1597 VTAIL.n85 VTAIL.n84 185
R1598 VTAIL.n87 VTAIL.n86 185
R1599 VTAIL.n273 VTAIL.n272 185
R1600 VTAIL.n271 VTAIL.n270 185
R1601 VTAIL.n192 VTAIL.n191 185
R1602 VTAIL.n265 VTAIL.n264 185
R1603 VTAIL.n263 VTAIL.n194 185
R1604 VTAIL.n262 VTAIL.n261 185
R1605 VTAIL.n197 VTAIL.n195 185
R1606 VTAIL.n256 VTAIL.n255 185
R1607 VTAIL.n254 VTAIL.n253 185
R1608 VTAIL.n201 VTAIL.n200 185
R1609 VTAIL.n248 VTAIL.n247 185
R1610 VTAIL.n246 VTAIL.n245 185
R1611 VTAIL.n205 VTAIL.n204 185
R1612 VTAIL.n240 VTAIL.n239 185
R1613 VTAIL.n238 VTAIL.n237 185
R1614 VTAIL.n209 VTAIL.n208 185
R1615 VTAIL.n232 VTAIL.n231 185
R1616 VTAIL.n230 VTAIL.n229 185
R1617 VTAIL.n213 VTAIL.n212 185
R1618 VTAIL.n224 VTAIL.n223 185
R1619 VTAIL.n222 VTAIL.n221 185
R1620 VTAIL.n217 VTAIL.n216 185
R1621 VTAIL.n181 VTAIL.n180 185
R1622 VTAIL.n179 VTAIL.n178 185
R1623 VTAIL.n100 VTAIL.n99 185
R1624 VTAIL.n173 VTAIL.n172 185
R1625 VTAIL.n171 VTAIL.n102 185
R1626 VTAIL.n170 VTAIL.n169 185
R1627 VTAIL.n105 VTAIL.n103 185
R1628 VTAIL.n164 VTAIL.n163 185
R1629 VTAIL.n162 VTAIL.n161 185
R1630 VTAIL.n109 VTAIL.n108 185
R1631 VTAIL.n156 VTAIL.n155 185
R1632 VTAIL.n154 VTAIL.n153 185
R1633 VTAIL.n113 VTAIL.n112 185
R1634 VTAIL.n148 VTAIL.n147 185
R1635 VTAIL.n146 VTAIL.n145 185
R1636 VTAIL.n117 VTAIL.n116 185
R1637 VTAIL.n140 VTAIL.n139 185
R1638 VTAIL.n138 VTAIL.n137 185
R1639 VTAIL.n121 VTAIL.n120 185
R1640 VTAIL.n132 VTAIL.n131 185
R1641 VTAIL.n130 VTAIL.n129 185
R1642 VTAIL.n125 VTAIL.n124 185
R1643 VTAIL.n307 VTAIL.t6 147.659
R1644 VTAIL.n31 VTAIL.t1 147.659
R1645 VTAIL.n218 VTAIL.t3 147.659
R1646 VTAIL.n126 VTAIL.t7 147.659
R1647 VTAIL.n311 VTAIL.n305 104.615
R1648 VTAIL.n312 VTAIL.n311 104.615
R1649 VTAIL.n312 VTAIL.n301 104.615
R1650 VTAIL.n319 VTAIL.n301 104.615
R1651 VTAIL.n320 VTAIL.n319 104.615
R1652 VTAIL.n320 VTAIL.n297 104.615
R1653 VTAIL.n327 VTAIL.n297 104.615
R1654 VTAIL.n328 VTAIL.n327 104.615
R1655 VTAIL.n328 VTAIL.n293 104.615
R1656 VTAIL.n335 VTAIL.n293 104.615
R1657 VTAIL.n336 VTAIL.n335 104.615
R1658 VTAIL.n336 VTAIL.n289 104.615
R1659 VTAIL.n343 VTAIL.n289 104.615
R1660 VTAIL.n344 VTAIL.n343 104.615
R1661 VTAIL.n344 VTAIL.n285 104.615
R1662 VTAIL.n352 VTAIL.n285 104.615
R1663 VTAIL.n353 VTAIL.n352 104.615
R1664 VTAIL.n354 VTAIL.n353 104.615
R1665 VTAIL.n354 VTAIL.n281 104.615
R1666 VTAIL.n361 VTAIL.n281 104.615
R1667 VTAIL.n362 VTAIL.n361 104.615
R1668 VTAIL.n35 VTAIL.n29 104.615
R1669 VTAIL.n36 VTAIL.n35 104.615
R1670 VTAIL.n36 VTAIL.n25 104.615
R1671 VTAIL.n43 VTAIL.n25 104.615
R1672 VTAIL.n44 VTAIL.n43 104.615
R1673 VTAIL.n44 VTAIL.n21 104.615
R1674 VTAIL.n51 VTAIL.n21 104.615
R1675 VTAIL.n52 VTAIL.n51 104.615
R1676 VTAIL.n52 VTAIL.n17 104.615
R1677 VTAIL.n59 VTAIL.n17 104.615
R1678 VTAIL.n60 VTAIL.n59 104.615
R1679 VTAIL.n60 VTAIL.n13 104.615
R1680 VTAIL.n67 VTAIL.n13 104.615
R1681 VTAIL.n68 VTAIL.n67 104.615
R1682 VTAIL.n68 VTAIL.n9 104.615
R1683 VTAIL.n76 VTAIL.n9 104.615
R1684 VTAIL.n77 VTAIL.n76 104.615
R1685 VTAIL.n78 VTAIL.n77 104.615
R1686 VTAIL.n78 VTAIL.n5 104.615
R1687 VTAIL.n85 VTAIL.n5 104.615
R1688 VTAIL.n86 VTAIL.n85 104.615
R1689 VTAIL.n272 VTAIL.n271 104.615
R1690 VTAIL.n271 VTAIL.n191 104.615
R1691 VTAIL.n264 VTAIL.n191 104.615
R1692 VTAIL.n264 VTAIL.n263 104.615
R1693 VTAIL.n263 VTAIL.n262 104.615
R1694 VTAIL.n262 VTAIL.n195 104.615
R1695 VTAIL.n255 VTAIL.n195 104.615
R1696 VTAIL.n255 VTAIL.n254 104.615
R1697 VTAIL.n254 VTAIL.n200 104.615
R1698 VTAIL.n247 VTAIL.n200 104.615
R1699 VTAIL.n247 VTAIL.n246 104.615
R1700 VTAIL.n246 VTAIL.n204 104.615
R1701 VTAIL.n239 VTAIL.n204 104.615
R1702 VTAIL.n239 VTAIL.n238 104.615
R1703 VTAIL.n238 VTAIL.n208 104.615
R1704 VTAIL.n231 VTAIL.n208 104.615
R1705 VTAIL.n231 VTAIL.n230 104.615
R1706 VTAIL.n230 VTAIL.n212 104.615
R1707 VTAIL.n223 VTAIL.n212 104.615
R1708 VTAIL.n223 VTAIL.n222 104.615
R1709 VTAIL.n222 VTAIL.n216 104.615
R1710 VTAIL.n180 VTAIL.n179 104.615
R1711 VTAIL.n179 VTAIL.n99 104.615
R1712 VTAIL.n172 VTAIL.n99 104.615
R1713 VTAIL.n172 VTAIL.n171 104.615
R1714 VTAIL.n171 VTAIL.n170 104.615
R1715 VTAIL.n170 VTAIL.n103 104.615
R1716 VTAIL.n163 VTAIL.n103 104.615
R1717 VTAIL.n163 VTAIL.n162 104.615
R1718 VTAIL.n162 VTAIL.n108 104.615
R1719 VTAIL.n155 VTAIL.n108 104.615
R1720 VTAIL.n155 VTAIL.n154 104.615
R1721 VTAIL.n154 VTAIL.n112 104.615
R1722 VTAIL.n147 VTAIL.n112 104.615
R1723 VTAIL.n147 VTAIL.n146 104.615
R1724 VTAIL.n146 VTAIL.n116 104.615
R1725 VTAIL.n139 VTAIL.n116 104.615
R1726 VTAIL.n139 VTAIL.n138 104.615
R1727 VTAIL.n138 VTAIL.n120 104.615
R1728 VTAIL.n131 VTAIL.n120 104.615
R1729 VTAIL.n131 VTAIL.n130 104.615
R1730 VTAIL.n130 VTAIL.n124 104.615
R1731 VTAIL.t6 VTAIL.n305 52.3082
R1732 VTAIL.t1 VTAIL.n29 52.3082
R1733 VTAIL.t3 VTAIL.n216 52.3082
R1734 VTAIL.t7 VTAIL.n124 52.3082
R1735 VTAIL.n187 VTAIL.n186 48.1717
R1736 VTAIL.n95 VTAIL.n94 48.1717
R1737 VTAIL.n1 VTAIL.n0 48.1715
R1738 VTAIL.n93 VTAIL.n92 48.1715
R1739 VTAIL.n367 VTAIL.n366 36.2581
R1740 VTAIL.n91 VTAIL.n90 36.2581
R1741 VTAIL.n277 VTAIL.n276 36.2581
R1742 VTAIL.n185 VTAIL.n184 36.2581
R1743 VTAIL.n95 VTAIL.n93 27.3927
R1744 VTAIL.n367 VTAIL.n277 26.9014
R1745 VTAIL.n307 VTAIL.n306 15.6677
R1746 VTAIL.n31 VTAIL.n30 15.6677
R1747 VTAIL.n218 VTAIL.n217 15.6677
R1748 VTAIL.n126 VTAIL.n125 15.6677
R1749 VTAIL.n355 VTAIL.n284 13.1884
R1750 VTAIL.n79 VTAIL.n8 13.1884
R1751 VTAIL.n265 VTAIL.n194 13.1884
R1752 VTAIL.n173 VTAIL.n102 13.1884
R1753 VTAIL.n310 VTAIL.n309 12.8005
R1754 VTAIL.n351 VTAIL.n350 12.8005
R1755 VTAIL.n356 VTAIL.n282 12.8005
R1756 VTAIL.n34 VTAIL.n33 12.8005
R1757 VTAIL.n75 VTAIL.n74 12.8005
R1758 VTAIL.n80 VTAIL.n6 12.8005
R1759 VTAIL.n266 VTAIL.n192 12.8005
R1760 VTAIL.n261 VTAIL.n196 12.8005
R1761 VTAIL.n221 VTAIL.n220 12.8005
R1762 VTAIL.n174 VTAIL.n100 12.8005
R1763 VTAIL.n169 VTAIL.n104 12.8005
R1764 VTAIL.n129 VTAIL.n128 12.8005
R1765 VTAIL.n313 VTAIL.n304 12.0247
R1766 VTAIL.n349 VTAIL.n286 12.0247
R1767 VTAIL.n360 VTAIL.n359 12.0247
R1768 VTAIL.n37 VTAIL.n28 12.0247
R1769 VTAIL.n73 VTAIL.n10 12.0247
R1770 VTAIL.n84 VTAIL.n83 12.0247
R1771 VTAIL.n270 VTAIL.n269 12.0247
R1772 VTAIL.n260 VTAIL.n197 12.0247
R1773 VTAIL.n224 VTAIL.n215 12.0247
R1774 VTAIL.n178 VTAIL.n177 12.0247
R1775 VTAIL.n168 VTAIL.n105 12.0247
R1776 VTAIL.n132 VTAIL.n123 12.0247
R1777 VTAIL.n314 VTAIL.n302 11.249
R1778 VTAIL.n346 VTAIL.n345 11.249
R1779 VTAIL.n363 VTAIL.n280 11.249
R1780 VTAIL.n38 VTAIL.n26 11.249
R1781 VTAIL.n70 VTAIL.n69 11.249
R1782 VTAIL.n87 VTAIL.n4 11.249
R1783 VTAIL.n273 VTAIL.n190 11.249
R1784 VTAIL.n257 VTAIL.n256 11.249
R1785 VTAIL.n225 VTAIL.n213 11.249
R1786 VTAIL.n181 VTAIL.n98 11.249
R1787 VTAIL.n165 VTAIL.n164 11.249
R1788 VTAIL.n133 VTAIL.n121 11.249
R1789 VTAIL.n318 VTAIL.n317 10.4732
R1790 VTAIL.n342 VTAIL.n288 10.4732
R1791 VTAIL.n364 VTAIL.n278 10.4732
R1792 VTAIL.n42 VTAIL.n41 10.4732
R1793 VTAIL.n66 VTAIL.n12 10.4732
R1794 VTAIL.n88 VTAIL.n2 10.4732
R1795 VTAIL.n274 VTAIL.n188 10.4732
R1796 VTAIL.n253 VTAIL.n199 10.4732
R1797 VTAIL.n229 VTAIL.n228 10.4732
R1798 VTAIL.n182 VTAIL.n96 10.4732
R1799 VTAIL.n161 VTAIL.n107 10.4732
R1800 VTAIL.n137 VTAIL.n136 10.4732
R1801 VTAIL.n321 VTAIL.n300 9.69747
R1802 VTAIL.n341 VTAIL.n290 9.69747
R1803 VTAIL.n45 VTAIL.n24 9.69747
R1804 VTAIL.n65 VTAIL.n14 9.69747
R1805 VTAIL.n252 VTAIL.n201 9.69747
R1806 VTAIL.n232 VTAIL.n211 9.69747
R1807 VTAIL.n160 VTAIL.n109 9.69747
R1808 VTAIL.n140 VTAIL.n119 9.69747
R1809 VTAIL.n366 VTAIL.n365 9.45567
R1810 VTAIL.n90 VTAIL.n89 9.45567
R1811 VTAIL.n276 VTAIL.n275 9.45567
R1812 VTAIL.n184 VTAIL.n183 9.45567
R1813 VTAIL.n365 VTAIL.n364 9.3005
R1814 VTAIL.n280 VTAIL.n279 9.3005
R1815 VTAIL.n359 VTAIL.n358 9.3005
R1816 VTAIL.n357 VTAIL.n356 9.3005
R1817 VTAIL.n296 VTAIL.n295 9.3005
R1818 VTAIL.n325 VTAIL.n324 9.3005
R1819 VTAIL.n323 VTAIL.n322 9.3005
R1820 VTAIL.n300 VTAIL.n299 9.3005
R1821 VTAIL.n317 VTAIL.n316 9.3005
R1822 VTAIL.n315 VTAIL.n314 9.3005
R1823 VTAIL.n304 VTAIL.n303 9.3005
R1824 VTAIL.n309 VTAIL.n308 9.3005
R1825 VTAIL.n331 VTAIL.n330 9.3005
R1826 VTAIL.n333 VTAIL.n332 9.3005
R1827 VTAIL.n292 VTAIL.n291 9.3005
R1828 VTAIL.n339 VTAIL.n338 9.3005
R1829 VTAIL.n341 VTAIL.n340 9.3005
R1830 VTAIL.n288 VTAIL.n287 9.3005
R1831 VTAIL.n347 VTAIL.n346 9.3005
R1832 VTAIL.n349 VTAIL.n348 9.3005
R1833 VTAIL.n350 VTAIL.n283 9.3005
R1834 VTAIL.n89 VTAIL.n88 9.3005
R1835 VTAIL.n4 VTAIL.n3 9.3005
R1836 VTAIL.n83 VTAIL.n82 9.3005
R1837 VTAIL.n81 VTAIL.n80 9.3005
R1838 VTAIL.n20 VTAIL.n19 9.3005
R1839 VTAIL.n49 VTAIL.n48 9.3005
R1840 VTAIL.n47 VTAIL.n46 9.3005
R1841 VTAIL.n24 VTAIL.n23 9.3005
R1842 VTAIL.n41 VTAIL.n40 9.3005
R1843 VTAIL.n39 VTAIL.n38 9.3005
R1844 VTAIL.n28 VTAIL.n27 9.3005
R1845 VTAIL.n33 VTAIL.n32 9.3005
R1846 VTAIL.n55 VTAIL.n54 9.3005
R1847 VTAIL.n57 VTAIL.n56 9.3005
R1848 VTAIL.n16 VTAIL.n15 9.3005
R1849 VTAIL.n63 VTAIL.n62 9.3005
R1850 VTAIL.n65 VTAIL.n64 9.3005
R1851 VTAIL.n12 VTAIL.n11 9.3005
R1852 VTAIL.n71 VTAIL.n70 9.3005
R1853 VTAIL.n73 VTAIL.n72 9.3005
R1854 VTAIL.n74 VTAIL.n7 9.3005
R1855 VTAIL.n244 VTAIL.n243 9.3005
R1856 VTAIL.n203 VTAIL.n202 9.3005
R1857 VTAIL.n250 VTAIL.n249 9.3005
R1858 VTAIL.n252 VTAIL.n251 9.3005
R1859 VTAIL.n199 VTAIL.n198 9.3005
R1860 VTAIL.n258 VTAIL.n257 9.3005
R1861 VTAIL.n260 VTAIL.n259 9.3005
R1862 VTAIL.n196 VTAIL.n193 9.3005
R1863 VTAIL.n275 VTAIL.n274 9.3005
R1864 VTAIL.n190 VTAIL.n189 9.3005
R1865 VTAIL.n269 VTAIL.n268 9.3005
R1866 VTAIL.n267 VTAIL.n266 9.3005
R1867 VTAIL.n242 VTAIL.n241 9.3005
R1868 VTAIL.n207 VTAIL.n206 9.3005
R1869 VTAIL.n236 VTAIL.n235 9.3005
R1870 VTAIL.n234 VTAIL.n233 9.3005
R1871 VTAIL.n211 VTAIL.n210 9.3005
R1872 VTAIL.n228 VTAIL.n227 9.3005
R1873 VTAIL.n226 VTAIL.n225 9.3005
R1874 VTAIL.n215 VTAIL.n214 9.3005
R1875 VTAIL.n220 VTAIL.n219 9.3005
R1876 VTAIL.n152 VTAIL.n151 9.3005
R1877 VTAIL.n111 VTAIL.n110 9.3005
R1878 VTAIL.n158 VTAIL.n157 9.3005
R1879 VTAIL.n160 VTAIL.n159 9.3005
R1880 VTAIL.n107 VTAIL.n106 9.3005
R1881 VTAIL.n166 VTAIL.n165 9.3005
R1882 VTAIL.n168 VTAIL.n167 9.3005
R1883 VTAIL.n104 VTAIL.n101 9.3005
R1884 VTAIL.n183 VTAIL.n182 9.3005
R1885 VTAIL.n98 VTAIL.n97 9.3005
R1886 VTAIL.n177 VTAIL.n176 9.3005
R1887 VTAIL.n175 VTAIL.n174 9.3005
R1888 VTAIL.n150 VTAIL.n149 9.3005
R1889 VTAIL.n115 VTAIL.n114 9.3005
R1890 VTAIL.n144 VTAIL.n143 9.3005
R1891 VTAIL.n142 VTAIL.n141 9.3005
R1892 VTAIL.n119 VTAIL.n118 9.3005
R1893 VTAIL.n136 VTAIL.n135 9.3005
R1894 VTAIL.n134 VTAIL.n133 9.3005
R1895 VTAIL.n123 VTAIL.n122 9.3005
R1896 VTAIL.n128 VTAIL.n127 9.3005
R1897 VTAIL.n322 VTAIL.n298 8.92171
R1898 VTAIL.n338 VTAIL.n337 8.92171
R1899 VTAIL.n46 VTAIL.n22 8.92171
R1900 VTAIL.n62 VTAIL.n61 8.92171
R1901 VTAIL.n249 VTAIL.n248 8.92171
R1902 VTAIL.n233 VTAIL.n209 8.92171
R1903 VTAIL.n157 VTAIL.n156 8.92171
R1904 VTAIL.n141 VTAIL.n117 8.92171
R1905 VTAIL.n326 VTAIL.n325 8.14595
R1906 VTAIL.n334 VTAIL.n292 8.14595
R1907 VTAIL.n50 VTAIL.n49 8.14595
R1908 VTAIL.n58 VTAIL.n16 8.14595
R1909 VTAIL.n245 VTAIL.n203 8.14595
R1910 VTAIL.n237 VTAIL.n236 8.14595
R1911 VTAIL.n153 VTAIL.n111 8.14595
R1912 VTAIL.n145 VTAIL.n144 8.14595
R1913 VTAIL.n329 VTAIL.n296 7.3702
R1914 VTAIL.n333 VTAIL.n294 7.3702
R1915 VTAIL.n53 VTAIL.n20 7.3702
R1916 VTAIL.n57 VTAIL.n18 7.3702
R1917 VTAIL.n244 VTAIL.n205 7.3702
R1918 VTAIL.n240 VTAIL.n207 7.3702
R1919 VTAIL.n152 VTAIL.n113 7.3702
R1920 VTAIL.n148 VTAIL.n115 7.3702
R1921 VTAIL.n330 VTAIL.n329 6.59444
R1922 VTAIL.n330 VTAIL.n294 6.59444
R1923 VTAIL.n54 VTAIL.n53 6.59444
R1924 VTAIL.n54 VTAIL.n18 6.59444
R1925 VTAIL.n241 VTAIL.n205 6.59444
R1926 VTAIL.n241 VTAIL.n240 6.59444
R1927 VTAIL.n149 VTAIL.n113 6.59444
R1928 VTAIL.n149 VTAIL.n148 6.59444
R1929 VTAIL.n326 VTAIL.n296 5.81868
R1930 VTAIL.n334 VTAIL.n333 5.81868
R1931 VTAIL.n50 VTAIL.n20 5.81868
R1932 VTAIL.n58 VTAIL.n57 5.81868
R1933 VTAIL.n245 VTAIL.n244 5.81868
R1934 VTAIL.n237 VTAIL.n207 5.81868
R1935 VTAIL.n153 VTAIL.n152 5.81868
R1936 VTAIL.n145 VTAIL.n115 5.81868
R1937 VTAIL.n325 VTAIL.n298 5.04292
R1938 VTAIL.n337 VTAIL.n292 5.04292
R1939 VTAIL.n49 VTAIL.n22 5.04292
R1940 VTAIL.n61 VTAIL.n16 5.04292
R1941 VTAIL.n248 VTAIL.n203 5.04292
R1942 VTAIL.n236 VTAIL.n209 5.04292
R1943 VTAIL.n156 VTAIL.n111 5.04292
R1944 VTAIL.n144 VTAIL.n117 5.04292
R1945 VTAIL.n308 VTAIL.n307 4.38563
R1946 VTAIL.n32 VTAIL.n31 4.38563
R1947 VTAIL.n219 VTAIL.n218 4.38563
R1948 VTAIL.n127 VTAIL.n126 4.38563
R1949 VTAIL.n322 VTAIL.n321 4.26717
R1950 VTAIL.n338 VTAIL.n290 4.26717
R1951 VTAIL.n46 VTAIL.n45 4.26717
R1952 VTAIL.n62 VTAIL.n14 4.26717
R1953 VTAIL.n249 VTAIL.n201 4.26717
R1954 VTAIL.n233 VTAIL.n232 4.26717
R1955 VTAIL.n157 VTAIL.n109 4.26717
R1956 VTAIL.n141 VTAIL.n140 4.26717
R1957 VTAIL.n318 VTAIL.n300 3.49141
R1958 VTAIL.n342 VTAIL.n341 3.49141
R1959 VTAIL.n366 VTAIL.n278 3.49141
R1960 VTAIL.n42 VTAIL.n24 3.49141
R1961 VTAIL.n66 VTAIL.n65 3.49141
R1962 VTAIL.n90 VTAIL.n2 3.49141
R1963 VTAIL.n276 VTAIL.n188 3.49141
R1964 VTAIL.n253 VTAIL.n252 3.49141
R1965 VTAIL.n229 VTAIL.n211 3.49141
R1966 VTAIL.n184 VTAIL.n96 3.49141
R1967 VTAIL.n161 VTAIL.n160 3.49141
R1968 VTAIL.n137 VTAIL.n119 3.49141
R1969 VTAIL.n317 VTAIL.n302 2.71565
R1970 VTAIL.n345 VTAIL.n288 2.71565
R1971 VTAIL.n364 VTAIL.n363 2.71565
R1972 VTAIL.n41 VTAIL.n26 2.71565
R1973 VTAIL.n69 VTAIL.n12 2.71565
R1974 VTAIL.n88 VTAIL.n87 2.71565
R1975 VTAIL.n274 VTAIL.n273 2.71565
R1976 VTAIL.n256 VTAIL.n199 2.71565
R1977 VTAIL.n228 VTAIL.n213 2.71565
R1978 VTAIL.n182 VTAIL.n181 2.71565
R1979 VTAIL.n164 VTAIL.n107 2.71565
R1980 VTAIL.n136 VTAIL.n121 2.71565
R1981 VTAIL.n314 VTAIL.n313 1.93989
R1982 VTAIL.n346 VTAIL.n286 1.93989
R1983 VTAIL.n360 VTAIL.n280 1.93989
R1984 VTAIL.n38 VTAIL.n37 1.93989
R1985 VTAIL.n70 VTAIL.n10 1.93989
R1986 VTAIL.n84 VTAIL.n4 1.93989
R1987 VTAIL.n270 VTAIL.n190 1.93989
R1988 VTAIL.n257 VTAIL.n197 1.93989
R1989 VTAIL.n225 VTAIL.n224 1.93989
R1990 VTAIL.n178 VTAIL.n98 1.93989
R1991 VTAIL.n165 VTAIL.n105 1.93989
R1992 VTAIL.n133 VTAIL.n132 1.93989
R1993 VTAIL.n0 VTAIL.t8 1.21597
R1994 VTAIL.n0 VTAIL.t9 1.21597
R1995 VTAIL.n92 VTAIL.t0 1.21597
R1996 VTAIL.n92 VTAIL.t10 1.21597
R1997 VTAIL.n186 VTAIL.t2 1.21597
R1998 VTAIL.n186 VTAIL.t11 1.21597
R1999 VTAIL.n94 VTAIL.t4 1.21597
R2000 VTAIL.n94 VTAIL.t5 1.21597
R2001 VTAIL.n310 VTAIL.n304 1.16414
R2002 VTAIL.n351 VTAIL.n349 1.16414
R2003 VTAIL.n359 VTAIL.n282 1.16414
R2004 VTAIL.n34 VTAIL.n28 1.16414
R2005 VTAIL.n75 VTAIL.n73 1.16414
R2006 VTAIL.n83 VTAIL.n6 1.16414
R2007 VTAIL.n269 VTAIL.n192 1.16414
R2008 VTAIL.n261 VTAIL.n260 1.16414
R2009 VTAIL.n221 VTAIL.n215 1.16414
R2010 VTAIL.n177 VTAIL.n100 1.16414
R2011 VTAIL.n169 VTAIL.n168 1.16414
R2012 VTAIL.n129 VTAIL.n123 1.16414
R2013 VTAIL.n187 VTAIL.n185 0.716017
R2014 VTAIL.n91 VTAIL.n1 0.716017
R2015 VTAIL.n185 VTAIL.n95 0.491879
R2016 VTAIL.n277 VTAIL.n187 0.491879
R2017 VTAIL.n93 VTAIL.n91 0.491879
R2018 VTAIL.n309 VTAIL.n306 0.388379
R2019 VTAIL.n350 VTAIL.n284 0.388379
R2020 VTAIL.n356 VTAIL.n355 0.388379
R2021 VTAIL.n33 VTAIL.n30 0.388379
R2022 VTAIL.n74 VTAIL.n8 0.388379
R2023 VTAIL.n80 VTAIL.n79 0.388379
R2024 VTAIL.n266 VTAIL.n265 0.388379
R2025 VTAIL.n196 VTAIL.n194 0.388379
R2026 VTAIL.n220 VTAIL.n217 0.388379
R2027 VTAIL.n174 VTAIL.n173 0.388379
R2028 VTAIL.n104 VTAIL.n102 0.388379
R2029 VTAIL.n128 VTAIL.n125 0.388379
R2030 VTAIL VTAIL.n367 0.310845
R2031 VTAIL VTAIL.n1 0.181534
R2032 VTAIL.n308 VTAIL.n303 0.155672
R2033 VTAIL.n315 VTAIL.n303 0.155672
R2034 VTAIL.n316 VTAIL.n315 0.155672
R2035 VTAIL.n316 VTAIL.n299 0.155672
R2036 VTAIL.n323 VTAIL.n299 0.155672
R2037 VTAIL.n324 VTAIL.n323 0.155672
R2038 VTAIL.n324 VTAIL.n295 0.155672
R2039 VTAIL.n331 VTAIL.n295 0.155672
R2040 VTAIL.n332 VTAIL.n331 0.155672
R2041 VTAIL.n332 VTAIL.n291 0.155672
R2042 VTAIL.n339 VTAIL.n291 0.155672
R2043 VTAIL.n340 VTAIL.n339 0.155672
R2044 VTAIL.n340 VTAIL.n287 0.155672
R2045 VTAIL.n347 VTAIL.n287 0.155672
R2046 VTAIL.n348 VTAIL.n347 0.155672
R2047 VTAIL.n348 VTAIL.n283 0.155672
R2048 VTAIL.n357 VTAIL.n283 0.155672
R2049 VTAIL.n358 VTAIL.n357 0.155672
R2050 VTAIL.n358 VTAIL.n279 0.155672
R2051 VTAIL.n365 VTAIL.n279 0.155672
R2052 VTAIL.n32 VTAIL.n27 0.155672
R2053 VTAIL.n39 VTAIL.n27 0.155672
R2054 VTAIL.n40 VTAIL.n39 0.155672
R2055 VTAIL.n40 VTAIL.n23 0.155672
R2056 VTAIL.n47 VTAIL.n23 0.155672
R2057 VTAIL.n48 VTAIL.n47 0.155672
R2058 VTAIL.n48 VTAIL.n19 0.155672
R2059 VTAIL.n55 VTAIL.n19 0.155672
R2060 VTAIL.n56 VTAIL.n55 0.155672
R2061 VTAIL.n56 VTAIL.n15 0.155672
R2062 VTAIL.n63 VTAIL.n15 0.155672
R2063 VTAIL.n64 VTAIL.n63 0.155672
R2064 VTAIL.n64 VTAIL.n11 0.155672
R2065 VTAIL.n71 VTAIL.n11 0.155672
R2066 VTAIL.n72 VTAIL.n71 0.155672
R2067 VTAIL.n72 VTAIL.n7 0.155672
R2068 VTAIL.n81 VTAIL.n7 0.155672
R2069 VTAIL.n82 VTAIL.n81 0.155672
R2070 VTAIL.n82 VTAIL.n3 0.155672
R2071 VTAIL.n89 VTAIL.n3 0.155672
R2072 VTAIL.n275 VTAIL.n189 0.155672
R2073 VTAIL.n268 VTAIL.n189 0.155672
R2074 VTAIL.n268 VTAIL.n267 0.155672
R2075 VTAIL.n267 VTAIL.n193 0.155672
R2076 VTAIL.n259 VTAIL.n193 0.155672
R2077 VTAIL.n259 VTAIL.n258 0.155672
R2078 VTAIL.n258 VTAIL.n198 0.155672
R2079 VTAIL.n251 VTAIL.n198 0.155672
R2080 VTAIL.n251 VTAIL.n250 0.155672
R2081 VTAIL.n250 VTAIL.n202 0.155672
R2082 VTAIL.n243 VTAIL.n202 0.155672
R2083 VTAIL.n243 VTAIL.n242 0.155672
R2084 VTAIL.n242 VTAIL.n206 0.155672
R2085 VTAIL.n235 VTAIL.n206 0.155672
R2086 VTAIL.n235 VTAIL.n234 0.155672
R2087 VTAIL.n234 VTAIL.n210 0.155672
R2088 VTAIL.n227 VTAIL.n210 0.155672
R2089 VTAIL.n227 VTAIL.n226 0.155672
R2090 VTAIL.n226 VTAIL.n214 0.155672
R2091 VTAIL.n219 VTAIL.n214 0.155672
R2092 VTAIL.n183 VTAIL.n97 0.155672
R2093 VTAIL.n176 VTAIL.n97 0.155672
R2094 VTAIL.n176 VTAIL.n175 0.155672
R2095 VTAIL.n175 VTAIL.n101 0.155672
R2096 VTAIL.n167 VTAIL.n101 0.155672
R2097 VTAIL.n167 VTAIL.n166 0.155672
R2098 VTAIL.n166 VTAIL.n106 0.155672
R2099 VTAIL.n159 VTAIL.n106 0.155672
R2100 VTAIL.n159 VTAIL.n158 0.155672
R2101 VTAIL.n158 VTAIL.n110 0.155672
R2102 VTAIL.n151 VTAIL.n110 0.155672
R2103 VTAIL.n151 VTAIL.n150 0.155672
R2104 VTAIL.n150 VTAIL.n114 0.155672
R2105 VTAIL.n143 VTAIL.n114 0.155672
R2106 VTAIL.n143 VTAIL.n142 0.155672
R2107 VTAIL.n142 VTAIL.n118 0.155672
R2108 VTAIL.n135 VTAIL.n118 0.155672
R2109 VTAIL.n135 VTAIL.n134 0.155672
R2110 VTAIL.n134 VTAIL.n122 0.155672
R2111 VTAIL.n127 VTAIL.n122 0.155672
R2112 VP.n7 VP.t4 1814.07
R2113 VP.n5 VP.t2 1814.07
R2114 VP.n0 VP.t5 1814.07
R2115 VP.n2 VP.t3 1814.07
R2116 VP.n6 VP.t0 1767.33
R2117 VP.n1 VP.t1 1767.33
R2118 VP.n3 VP.n0 161.489
R2119 VP.n8 VP.n7 161.3
R2120 VP.n3 VP.n2 161.3
R2121 VP.n5 VP.n4 161.3
R2122 VP.n4 VP.n3 42.7543
R2123 VP.n6 VP.n5 36.5157
R2124 VP.n7 VP.n6 36.5157
R2125 VP.n1 VP.n0 36.5157
R2126 VP.n2 VP.n1 36.5157
R2127 VP.n8 VP.n4 0.189894
R2128 VP VP.n8 0.0516364
R2129 VDD1.n84 VDD1.n0 289.615
R2130 VDD1.n173 VDD1.n89 289.615
R2131 VDD1.n85 VDD1.n84 185
R2132 VDD1.n83 VDD1.n82 185
R2133 VDD1.n4 VDD1.n3 185
R2134 VDD1.n77 VDD1.n76 185
R2135 VDD1.n75 VDD1.n6 185
R2136 VDD1.n74 VDD1.n73 185
R2137 VDD1.n9 VDD1.n7 185
R2138 VDD1.n68 VDD1.n67 185
R2139 VDD1.n66 VDD1.n65 185
R2140 VDD1.n13 VDD1.n12 185
R2141 VDD1.n60 VDD1.n59 185
R2142 VDD1.n58 VDD1.n57 185
R2143 VDD1.n17 VDD1.n16 185
R2144 VDD1.n52 VDD1.n51 185
R2145 VDD1.n50 VDD1.n49 185
R2146 VDD1.n21 VDD1.n20 185
R2147 VDD1.n44 VDD1.n43 185
R2148 VDD1.n42 VDD1.n41 185
R2149 VDD1.n25 VDD1.n24 185
R2150 VDD1.n36 VDD1.n35 185
R2151 VDD1.n34 VDD1.n33 185
R2152 VDD1.n29 VDD1.n28 185
R2153 VDD1.n117 VDD1.n116 185
R2154 VDD1.n122 VDD1.n121 185
R2155 VDD1.n124 VDD1.n123 185
R2156 VDD1.n113 VDD1.n112 185
R2157 VDD1.n130 VDD1.n129 185
R2158 VDD1.n132 VDD1.n131 185
R2159 VDD1.n109 VDD1.n108 185
R2160 VDD1.n138 VDD1.n137 185
R2161 VDD1.n140 VDD1.n139 185
R2162 VDD1.n105 VDD1.n104 185
R2163 VDD1.n146 VDD1.n145 185
R2164 VDD1.n148 VDD1.n147 185
R2165 VDD1.n101 VDD1.n100 185
R2166 VDD1.n154 VDD1.n153 185
R2167 VDD1.n156 VDD1.n155 185
R2168 VDD1.n97 VDD1.n96 185
R2169 VDD1.n163 VDD1.n162 185
R2170 VDD1.n164 VDD1.n95 185
R2171 VDD1.n166 VDD1.n165 185
R2172 VDD1.n93 VDD1.n92 185
R2173 VDD1.n172 VDD1.n171 185
R2174 VDD1.n174 VDD1.n173 185
R2175 VDD1.n30 VDD1.t0 147.659
R2176 VDD1.n118 VDD1.t3 147.659
R2177 VDD1.n84 VDD1.n83 104.615
R2178 VDD1.n83 VDD1.n3 104.615
R2179 VDD1.n76 VDD1.n3 104.615
R2180 VDD1.n76 VDD1.n75 104.615
R2181 VDD1.n75 VDD1.n74 104.615
R2182 VDD1.n74 VDD1.n7 104.615
R2183 VDD1.n67 VDD1.n7 104.615
R2184 VDD1.n67 VDD1.n66 104.615
R2185 VDD1.n66 VDD1.n12 104.615
R2186 VDD1.n59 VDD1.n12 104.615
R2187 VDD1.n59 VDD1.n58 104.615
R2188 VDD1.n58 VDD1.n16 104.615
R2189 VDD1.n51 VDD1.n16 104.615
R2190 VDD1.n51 VDD1.n50 104.615
R2191 VDD1.n50 VDD1.n20 104.615
R2192 VDD1.n43 VDD1.n20 104.615
R2193 VDD1.n43 VDD1.n42 104.615
R2194 VDD1.n42 VDD1.n24 104.615
R2195 VDD1.n35 VDD1.n24 104.615
R2196 VDD1.n35 VDD1.n34 104.615
R2197 VDD1.n34 VDD1.n28 104.615
R2198 VDD1.n122 VDD1.n116 104.615
R2199 VDD1.n123 VDD1.n122 104.615
R2200 VDD1.n123 VDD1.n112 104.615
R2201 VDD1.n130 VDD1.n112 104.615
R2202 VDD1.n131 VDD1.n130 104.615
R2203 VDD1.n131 VDD1.n108 104.615
R2204 VDD1.n138 VDD1.n108 104.615
R2205 VDD1.n139 VDD1.n138 104.615
R2206 VDD1.n139 VDD1.n104 104.615
R2207 VDD1.n146 VDD1.n104 104.615
R2208 VDD1.n147 VDD1.n146 104.615
R2209 VDD1.n147 VDD1.n100 104.615
R2210 VDD1.n154 VDD1.n100 104.615
R2211 VDD1.n155 VDD1.n154 104.615
R2212 VDD1.n155 VDD1.n96 104.615
R2213 VDD1.n163 VDD1.n96 104.615
R2214 VDD1.n164 VDD1.n163 104.615
R2215 VDD1.n165 VDD1.n164 104.615
R2216 VDD1.n165 VDD1.n92 104.615
R2217 VDD1.n172 VDD1.n92 104.615
R2218 VDD1.n173 VDD1.n172 104.615
R2219 VDD1.n179 VDD1.n178 64.9178
R2220 VDD1.n181 VDD1.n180 64.8503
R2221 VDD1 VDD1.n88 53.3636
R2222 VDD1.n179 VDD1.n177 53.25
R2223 VDD1.t0 VDD1.n28 52.3082
R2224 VDD1.t3 VDD1.n116 52.3082
R2225 VDD1.n181 VDD1.n179 40.1841
R2226 VDD1.n30 VDD1.n29 15.6677
R2227 VDD1.n118 VDD1.n117 15.6677
R2228 VDD1.n77 VDD1.n6 13.1884
R2229 VDD1.n166 VDD1.n95 13.1884
R2230 VDD1.n78 VDD1.n4 12.8005
R2231 VDD1.n73 VDD1.n8 12.8005
R2232 VDD1.n33 VDD1.n32 12.8005
R2233 VDD1.n121 VDD1.n120 12.8005
R2234 VDD1.n162 VDD1.n161 12.8005
R2235 VDD1.n167 VDD1.n93 12.8005
R2236 VDD1.n82 VDD1.n81 12.0247
R2237 VDD1.n72 VDD1.n9 12.0247
R2238 VDD1.n36 VDD1.n27 12.0247
R2239 VDD1.n124 VDD1.n115 12.0247
R2240 VDD1.n160 VDD1.n97 12.0247
R2241 VDD1.n171 VDD1.n170 12.0247
R2242 VDD1.n85 VDD1.n2 11.249
R2243 VDD1.n69 VDD1.n68 11.249
R2244 VDD1.n37 VDD1.n25 11.249
R2245 VDD1.n125 VDD1.n113 11.249
R2246 VDD1.n157 VDD1.n156 11.249
R2247 VDD1.n174 VDD1.n91 11.249
R2248 VDD1.n86 VDD1.n0 10.4732
R2249 VDD1.n65 VDD1.n11 10.4732
R2250 VDD1.n41 VDD1.n40 10.4732
R2251 VDD1.n129 VDD1.n128 10.4732
R2252 VDD1.n153 VDD1.n99 10.4732
R2253 VDD1.n175 VDD1.n89 10.4732
R2254 VDD1.n64 VDD1.n13 9.69747
R2255 VDD1.n44 VDD1.n23 9.69747
R2256 VDD1.n132 VDD1.n111 9.69747
R2257 VDD1.n152 VDD1.n101 9.69747
R2258 VDD1.n88 VDD1.n87 9.45567
R2259 VDD1.n177 VDD1.n176 9.45567
R2260 VDD1.n56 VDD1.n55 9.3005
R2261 VDD1.n15 VDD1.n14 9.3005
R2262 VDD1.n62 VDD1.n61 9.3005
R2263 VDD1.n64 VDD1.n63 9.3005
R2264 VDD1.n11 VDD1.n10 9.3005
R2265 VDD1.n70 VDD1.n69 9.3005
R2266 VDD1.n72 VDD1.n71 9.3005
R2267 VDD1.n8 VDD1.n5 9.3005
R2268 VDD1.n87 VDD1.n86 9.3005
R2269 VDD1.n2 VDD1.n1 9.3005
R2270 VDD1.n81 VDD1.n80 9.3005
R2271 VDD1.n79 VDD1.n78 9.3005
R2272 VDD1.n54 VDD1.n53 9.3005
R2273 VDD1.n19 VDD1.n18 9.3005
R2274 VDD1.n48 VDD1.n47 9.3005
R2275 VDD1.n46 VDD1.n45 9.3005
R2276 VDD1.n23 VDD1.n22 9.3005
R2277 VDD1.n40 VDD1.n39 9.3005
R2278 VDD1.n38 VDD1.n37 9.3005
R2279 VDD1.n27 VDD1.n26 9.3005
R2280 VDD1.n32 VDD1.n31 9.3005
R2281 VDD1.n176 VDD1.n175 9.3005
R2282 VDD1.n91 VDD1.n90 9.3005
R2283 VDD1.n170 VDD1.n169 9.3005
R2284 VDD1.n168 VDD1.n167 9.3005
R2285 VDD1.n107 VDD1.n106 9.3005
R2286 VDD1.n136 VDD1.n135 9.3005
R2287 VDD1.n134 VDD1.n133 9.3005
R2288 VDD1.n111 VDD1.n110 9.3005
R2289 VDD1.n128 VDD1.n127 9.3005
R2290 VDD1.n126 VDD1.n125 9.3005
R2291 VDD1.n115 VDD1.n114 9.3005
R2292 VDD1.n120 VDD1.n119 9.3005
R2293 VDD1.n142 VDD1.n141 9.3005
R2294 VDD1.n144 VDD1.n143 9.3005
R2295 VDD1.n103 VDD1.n102 9.3005
R2296 VDD1.n150 VDD1.n149 9.3005
R2297 VDD1.n152 VDD1.n151 9.3005
R2298 VDD1.n99 VDD1.n98 9.3005
R2299 VDD1.n158 VDD1.n157 9.3005
R2300 VDD1.n160 VDD1.n159 9.3005
R2301 VDD1.n161 VDD1.n94 9.3005
R2302 VDD1.n61 VDD1.n60 8.92171
R2303 VDD1.n45 VDD1.n21 8.92171
R2304 VDD1.n133 VDD1.n109 8.92171
R2305 VDD1.n149 VDD1.n148 8.92171
R2306 VDD1.n57 VDD1.n15 8.14595
R2307 VDD1.n49 VDD1.n48 8.14595
R2308 VDD1.n137 VDD1.n136 8.14595
R2309 VDD1.n145 VDD1.n103 8.14595
R2310 VDD1.n56 VDD1.n17 7.3702
R2311 VDD1.n52 VDD1.n19 7.3702
R2312 VDD1.n140 VDD1.n107 7.3702
R2313 VDD1.n144 VDD1.n105 7.3702
R2314 VDD1.n53 VDD1.n17 6.59444
R2315 VDD1.n53 VDD1.n52 6.59444
R2316 VDD1.n141 VDD1.n140 6.59444
R2317 VDD1.n141 VDD1.n105 6.59444
R2318 VDD1.n57 VDD1.n56 5.81868
R2319 VDD1.n49 VDD1.n19 5.81868
R2320 VDD1.n137 VDD1.n107 5.81868
R2321 VDD1.n145 VDD1.n144 5.81868
R2322 VDD1.n60 VDD1.n15 5.04292
R2323 VDD1.n48 VDD1.n21 5.04292
R2324 VDD1.n136 VDD1.n109 5.04292
R2325 VDD1.n148 VDD1.n103 5.04292
R2326 VDD1.n31 VDD1.n30 4.38563
R2327 VDD1.n119 VDD1.n118 4.38563
R2328 VDD1.n61 VDD1.n13 4.26717
R2329 VDD1.n45 VDD1.n44 4.26717
R2330 VDD1.n133 VDD1.n132 4.26717
R2331 VDD1.n149 VDD1.n101 4.26717
R2332 VDD1.n88 VDD1.n0 3.49141
R2333 VDD1.n65 VDD1.n64 3.49141
R2334 VDD1.n41 VDD1.n23 3.49141
R2335 VDD1.n129 VDD1.n111 3.49141
R2336 VDD1.n153 VDD1.n152 3.49141
R2337 VDD1.n177 VDD1.n89 3.49141
R2338 VDD1.n86 VDD1.n85 2.71565
R2339 VDD1.n68 VDD1.n11 2.71565
R2340 VDD1.n40 VDD1.n25 2.71565
R2341 VDD1.n128 VDD1.n113 2.71565
R2342 VDD1.n156 VDD1.n99 2.71565
R2343 VDD1.n175 VDD1.n174 2.71565
R2344 VDD1.n82 VDD1.n2 1.93989
R2345 VDD1.n69 VDD1.n9 1.93989
R2346 VDD1.n37 VDD1.n36 1.93989
R2347 VDD1.n125 VDD1.n124 1.93989
R2348 VDD1.n157 VDD1.n97 1.93989
R2349 VDD1.n171 VDD1.n91 1.93989
R2350 VDD1.n180 VDD1.t4 1.21597
R2351 VDD1.n180 VDD1.t2 1.21597
R2352 VDD1.n178 VDD1.t5 1.21597
R2353 VDD1.n178 VDD1.t1 1.21597
R2354 VDD1.n81 VDD1.n4 1.16414
R2355 VDD1.n73 VDD1.n72 1.16414
R2356 VDD1.n33 VDD1.n27 1.16414
R2357 VDD1.n121 VDD1.n115 1.16414
R2358 VDD1.n162 VDD1.n160 1.16414
R2359 VDD1.n170 VDD1.n93 1.16414
R2360 VDD1.n78 VDD1.n77 0.388379
R2361 VDD1.n8 VDD1.n6 0.388379
R2362 VDD1.n32 VDD1.n29 0.388379
R2363 VDD1.n120 VDD1.n117 0.388379
R2364 VDD1.n161 VDD1.n95 0.388379
R2365 VDD1.n167 VDD1.n166 0.388379
R2366 VDD1.n87 VDD1.n1 0.155672
R2367 VDD1.n80 VDD1.n1 0.155672
R2368 VDD1.n80 VDD1.n79 0.155672
R2369 VDD1.n79 VDD1.n5 0.155672
R2370 VDD1.n71 VDD1.n5 0.155672
R2371 VDD1.n71 VDD1.n70 0.155672
R2372 VDD1.n70 VDD1.n10 0.155672
R2373 VDD1.n63 VDD1.n10 0.155672
R2374 VDD1.n63 VDD1.n62 0.155672
R2375 VDD1.n62 VDD1.n14 0.155672
R2376 VDD1.n55 VDD1.n14 0.155672
R2377 VDD1.n55 VDD1.n54 0.155672
R2378 VDD1.n54 VDD1.n18 0.155672
R2379 VDD1.n47 VDD1.n18 0.155672
R2380 VDD1.n47 VDD1.n46 0.155672
R2381 VDD1.n46 VDD1.n22 0.155672
R2382 VDD1.n39 VDD1.n22 0.155672
R2383 VDD1.n39 VDD1.n38 0.155672
R2384 VDD1.n38 VDD1.n26 0.155672
R2385 VDD1.n31 VDD1.n26 0.155672
R2386 VDD1.n119 VDD1.n114 0.155672
R2387 VDD1.n126 VDD1.n114 0.155672
R2388 VDD1.n127 VDD1.n126 0.155672
R2389 VDD1.n127 VDD1.n110 0.155672
R2390 VDD1.n134 VDD1.n110 0.155672
R2391 VDD1.n135 VDD1.n134 0.155672
R2392 VDD1.n135 VDD1.n106 0.155672
R2393 VDD1.n142 VDD1.n106 0.155672
R2394 VDD1.n143 VDD1.n142 0.155672
R2395 VDD1.n143 VDD1.n102 0.155672
R2396 VDD1.n150 VDD1.n102 0.155672
R2397 VDD1.n151 VDD1.n150 0.155672
R2398 VDD1.n151 VDD1.n98 0.155672
R2399 VDD1.n158 VDD1.n98 0.155672
R2400 VDD1.n159 VDD1.n158 0.155672
R2401 VDD1.n159 VDD1.n94 0.155672
R2402 VDD1.n168 VDD1.n94 0.155672
R2403 VDD1.n169 VDD1.n168 0.155672
R2404 VDD1.n169 VDD1.n90 0.155672
R2405 VDD1.n176 VDD1.n90 0.155672
R2406 VDD1 VDD1.n181 0.0651552
C0 VP VN 5.42721f
C1 VDD1 VP 3.2392f
C2 VDD1 VN 0.147327f
C3 VTAIL VP 2.46039f
C4 VDD2 VP 0.259506f
C5 VTAIL VN 2.44536f
C6 VDD2 VN 3.13406f
C7 VTAIL VDD1 20.064f
C8 VDD2 VDD1 0.550725f
C9 VDD2 VTAIL 20.0895f
C10 VDD2 B 4.930918f
C11 VDD1 B 4.874904f
C12 VTAIL B 7.474251f
C13 VN B 7.31843f
C14 VP B 4.668256f
C15 VDD1.n0 B 0.043539f
C16 VDD1.n1 B 0.029693f
C17 VDD1.n2 B 0.015956f
C18 VDD1.n3 B 0.037714f
C19 VDD1.n4 B 0.016894f
C20 VDD1.n5 B 0.029693f
C21 VDD1.n6 B 0.016425f
C22 VDD1.n7 B 0.037714f
C23 VDD1.n8 B 0.015956f
C24 VDD1.n9 B 0.016894f
C25 VDD1.n10 B 0.029693f
C26 VDD1.n11 B 0.015956f
C27 VDD1.n12 B 0.037714f
C28 VDD1.n13 B 0.016894f
C29 VDD1.n14 B 0.029693f
C30 VDD1.n15 B 0.015956f
C31 VDD1.n16 B 0.037714f
C32 VDD1.n17 B 0.016894f
C33 VDD1.n18 B 0.029693f
C34 VDD1.n19 B 0.015956f
C35 VDD1.n20 B 0.037714f
C36 VDD1.n21 B 0.016894f
C37 VDD1.n22 B 0.029693f
C38 VDD1.n23 B 0.015956f
C39 VDD1.n24 B 0.037714f
C40 VDD1.n25 B 0.016894f
C41 VDD1.n26 B 0.029693f
C42 VDD1.n27 B 0.015956f
C43 VDD1.n28 B 0.028285f
C44 VDD1.n29 B 0.022279f
C45 VDD1.t0 B 0.062316f
C46 VDD1.n30 B 0.203267f
C47 VDD1.n31 B 2.10741f
C48 VDD1.n32 B 0.015956f
C49 VDD1.n33 B 0.016894f
C50 VDD1.n34 B 0.037714f
C51 VDD1.n35 B 0.037714f
C52 VDD1.n36 B 0.016894f
C53 VDD1.n37 B 0.015956f
C54 VDD1.n38 B 0.029693f
C55 VDD1.n39 B 0.029693f
C56 VDD1.n40 B 0.015956f
C57 VDD1.n41 B 0.016894f
C58 VDD1.n42 B 0.037714f
C59 VDD1.n43 B 0.037714f
C60 VDD1.n44 B 0.016894f
C61 VDD1.n45 B 0.015956f
C62 VDD1.n46 B 0.029693f
C63 VDD1.n47 B 0.029693f
C64 VDD1.n48 B 0.015956f
C65 VDD1.n49 B 0.016894f
C66 VDD1.n50 B 0.037714f
C67 VDD1.n51 B 0.037714f
C68 VDD1.n52 B 0.016894f
C69 VDD1.n53 B 0.015956f
C70 VDD1.n54 B 0.029693f
C71 VDD1.n55 B 0.029693f
C72 VDD1.n56 B 0.015956f
C73 VDD1.n57 B 0.016894f
C74 VDD1.n58 B 0.037714f
C75 VDD1.n59 B 0.037714f
C76 VDD1.n60 B 0.016894f
C77 VDD1.n61 B 0.015956f
C78 VDD1.n62 B 0.029693f
C79 VDD1.n63 B 0.029693f
C80 VDD1.n64 B 0.015956f
C81 VDD1.n65 B 0.016894f
C82 VDD1.n66 B 0.037714f
C83 VDD1.n67 B 0.037714f
C84 VDD1.n68 B 0.016894f
C85 VDD1.n69 B 0.015956f
C86 VDD1.n70 B 0.029693f
C87 VDD1.n71 B 0.029693f
C88 VDD1.n72 B 0.015956f
C89 VDD1.n73 B 0.016894f
C90 VDD1.n74 B 0.037714f
C91 VDD1.n75 B 0.037714f
C92 VDD1.n76 B 0.037714f
C93 VDD1.n77 B 0.016425f
C94 VDD1.n78 B 0.015956f
C95 VDD1.n79 B 0.029693f
C96 VDD1.n80 B 0.029693f
C97 VDD1.n81 B 0.015956f
C98 VDD1.n82 B 0.016894f
C99 VDD1.n83 B 0.037714f
C100 VDD1.n84 B 0.084832f
C101 VDD1.n85 B 0.016894f
C102 VDD1.n86 B 0.015956f
C103 VDD1.n87 B 0.077152f
C104 VDD1.n88 B 0.069309f
C105 VDD1.n89 B 0.043539f
C106 VDD1.n90 B 0.029693f
C107 VDD1.n91 B 0.015956f
C108 VDD1.n92 B 0.037714f
C109 VDD1.n93 B 0.016894f
C110 VDD1.n94 B 0.029693f
C111 VDD1.n95 B 0.016425f
C112 VDD1.n96 B 0.037714f
C113 VDD1.n97 B 0.016894f
C114 VDD1.n98 B 0.029693f
C115 VDD1.n99 B 0.015956f
C116 VDD1.n100 B 0.037714f
C117 VDD1.n101 B 0.016894f
C118 VDD1.n102 B 0.029693f
C119 VDD1.n103 B 0.015956f
C120 VDD1.n104 B 0.037714f
C121 VDD1.n105 B 0.016894f
C122 VDD1.n106 B 0.029693f
C123 VDD1.n107 B 0.015956f
C124 VDD1.n108 B 0.037714f
C125 VDD1.n109 B 0.016894f
C126 VDD1.n110 B 0.029693f
C127 VDD1.n111 B 0.015956f
C128 VDD1.n112 B 0.037714f
C129 VDD1.n113 B 0.016894f
C130 VDD1.n114 B 0.029693f
C131 VDD1.n115 B 0.015956f
C132 VDD1.n116 B 0.028285f
C133 VDD1.n117 B 0.022279f
C134 VDD1.t3 B 0.062316f
C135 VDD1.n118 B 0.203267f
C136 VDD1.n119 B 2.10741f
C137 VDD1.n120 B 0.015956f
C138 VDD1.n121 B 0.016894f
C139 VDD1.n122 B 0.037714f
C140 VDD1.n123 B 0.037714f
C141 VDD1.n124 B 0.016894f
C142 VDD1.n125 B 0.015956f
C143 VDD1.n126 B 0.029693f
C144 VDD1.n127 B 0.029693f
C145 VDD1.n128 B 0.015956f
C146 VDD1.n129 B 0.016894f
C147 VDD1.n130 B 0.037714f
C148 VDD1.n131 B 0.037714f
C149 VDD1.n132 B 0.016894f
C150 VDD1.n133 B 0.015956f
C151 VDD1.n134 B 0.029693f
C152 VDD1.n135 B 0.029693f
C153 VDD1.n136 B 0.015956f
C154 VDD1.n137 B 0.016894f
C155 VDD1.n138 B 0.037714f
C156 VDD1.n139 B 0.037714f
C157 VDD1.n140 B 0.016894f
C158 VDD1.n141 B 0.015956f
C159 VDD1.n142 B 0.029693f
C160 VDD1.n143 B 0.029693f
C161 VDD1.n144 B 0.015956f
C162 VDD1.n145 B 0.016894f
C163 VDD1.n146 B 0.037714f
C164 VDD1.n147 B 0.037714f
C165 VDD1.n148 B 0.016894f
C166 VDD1.n149 B 0.015956f
C167 VDD1.n150 B 0.029693f
C168 VDD1.n151 B 0.029693f
C169 VDD1.n152 B 0.015956f
C170 VDD1.n153 B 0.016894f
C171 VDD1.n154 B 0.037714f
C172 VDD1.n155 B 0.037714f
C173 VDD1.n156 B 0.016894f
C174 VDD1.n157 B 0.015956f
C175 VDD1.n158 B 0.029693f
C176 VDD1.n159 B 0.029693f
C177 VDD1.n160 B 0.015956f
C178 VDD1.n161 B 0.015956f
C179 VDD1.n162 B 0.016894f
C180 VDD1.n163 B 0.037714f
C181 VDD1.n164 B 0.037714f
C182 VDD1.n165 B 0.037714f
C183 VDD1.n166 B 0.016425f
C184 VDD1.n167 B 0.015956f
C185 VDD1.n168 B 0.029693f
C186 VDD1.n169 B 0.029693f
C187 VDD1.n170 B 0.015956f
C188 VDD1.n171 B 0.016894f
C189 VDD1.n172 B 0.037714f
C190 VDD1.n173 B 0.084832f
C191 VDD1.n174 B 0.016894f
C192 VDD1.n175 B 0.015956f
C193 VDD1.n176 B 0.077152f
C194 VDD1.n177 B 0.069041f
C195 VDD1.t5 B 0.382233f
C196 VDD1.t1 B 0.382233f
C197 VDD1.n178 B 3.47324f
C198 VDD1.n179 B 2.35347f
C199 VDD1.t4 B 0.382233f
C200 VDD1.t2 B 0.382233f
C201 VDD1.n180 B 3.47292f
C202 VDD1.n181 B 2.91116f
C203 VP.t5 B 0.680472f
C204 VP.n0 B 0.278438f
C205 VP.t1 B 0.673717f
C206 VP.n1 B 0.259938f
C207 VP.t3 B 0.680472f
C208 VP.n2 B 0.27835f
C209 VP.n3 B 2.67293f
C210 VP.n4 B 2.64897f
C211 VP.t0 B 0.673717f
C212 VP.t2 B 0.680472f
C213 VP.n5 B 0.27835f
C214 VP.n6 B 0.259938f
C215 VP.t4 B 0.680472f
C216 VP.n7 B 0.27835f
C217 VP.n8 B 0.047352f
C218 VTAIL.t8 B 0.387168f
C219 VTAIL.t9 B 0.387168f
C220 VTAIL.n0 B 3.4357f
C221 VTAIL.n1 B 0.370806f
C222 VTAIL.n2 B 0.044101f
C223 VTAIL.n3 B 0.030076f
C224 VTAIL.n4 B 0.016162f
C225 VTAIL.n5 B 0.0382f
C226 VTAIL.n6 B 0.017112f
C227 VTAIL.n7 B 0.030076f
C228 VTAIL.n8 B 0.016637f
C229 VTAIL.n9 B 0.0382f
C230 VTAIL.n10 B 0.017112f
C231 VTAIL.n11 B 0.030076f
C232 VTAIL.n12 B 0.016162f
C233 VTAIL.n13 B 0.0382f
C234 VTAIL.n14 B 0.017112f
C235 VTAIL.n15 B 0.030076f
C236 VTAIL.n16 B 0.016162f
C237 VTAIL.n17 B 0.0382f
C238 VTAIL.n18 B 0.017112f
C239 VTAIL.n19 B 0.030076f
C240 VTAIL.n20 B 0.016162f
C241 VTAIL.n21 B 0.0382f
C242 VTAIL.n22 B 0.017112f
C243 VTAIL.n23 B 0.030076f
C244 VTAIL.n24 B 0.016162f
C245 VTAIL.n25 B 0.0382f
C246 VTAIL.n26 B 0.017112f
C247 VTAIL.n27 B 0.030076f
C248 VTAIL.n28 B 0.016162f
C249 VTAIL.n29 B 0.02865f
C250 VTAIL.n30 B 0.022566f
C251 VTAIL.t1 B 0.063121f
C252 VTAIL.n31 B 0.205892f
C253 VTAIL.n32 B 2.13462f
C254 VTAIL.n33 B 0.016162f
C255 VTAIL.n34 B 0.017112f
C256 VTAIL.n35 B 0.0382f
C257 VTAIL.n36 B 0.0382f
C258 VTAIL.n37 B 0.017112f
C259 VTAIL.n38 B 0.016162f
C260 VTAIL.n39 B 0.030076f
C261 VTAIL.n40 B 0.030076f
C262 VTAIL.n41 B 0.016162f
C263 VTAIL.n42 B 0.017112f
C264 VTAIL.n43 B 0.0382f
C265 VTAIL.n44 B 0.0382f
C266 VTAIL.n45 B 0.017112f
C267 VTAIL.n46 B 0.016162f
C268 VTAIL.n47 B 0.030076f
C269 VTAIL.n48 B 0.030076f
C270 VTAIL.n49 B 0.016162f
C271 VTAIL.n50 B 0.017112f
C272 VTAIL.n51 B 0.0382f
C273 VTAIL.n52 B 0.0382f
C274 VTAIL.n53 B 0.017112f
C275 VTAIL.n54 B 0.016162f
C276 VTAIL.n55 B 0.030076f
C277 VTAIL.n56 B 0.030076f
C278 VTAIL.n57 B 0.016162f
C279 VTAIL.n58 B 0.017112f
C280 VTAIL.n59 B 0.0382f
C281 VTAIL.n60 B 0.0382f
C282 VTAIL.n61 B 0.017112f
C283 VTAIL.n62 B 0.016162f
C284 VTAIL.n63 B 0.030076f
C285 VTAIL.n64 B 0.030076f
C286 VTAIL.n65 B 0.016162f
C287 VTAIL.n66 B 0.017112f
C288 VTAIL.n67 B 0.0382f
C289 VTAIL.n68 B 0.0382f
C290 VTAIL.n69 B 0.017112f
C291 VTAIL.n70 B 0.016162f
C292 VTAIL.n71 B 0.030076f
C293 VTAIL.n72 B 0.030076f
C294 VTAIL.n73 B 0.016162f
C295 VTAIL.n74 B 0.016162f
C296 VTAIL.n75 B 0.017112f
C297 VTAIL.n76 B 0.0382f
C298 VTAIL.n77 B 0.0382f
C299 VTAIL.n78 B 0.0382f
C300 VTAIL.n79 B 0.016637f
C301 VTAIL.n80 B 0.016162f
C302 VTAIL.n81 B 0.030076f
C303 VTAIL.n82 B 0.030076f
C304 VTAIL.n83 B 0.016162f
C305 VTAIL.n84 B 0.017112f
C306 VTAIL.n85 B 0.0382f
C307 VTAIL.n86 B 0.085927f
C308 VTAIL.n87 B 0.017112f
C309 VTAIL.n88 B 0.016162f
C310 VTAIL.n89 B 0.078148f
C311 VTAIL.n90 B 0.048663f
C312 VTAIL.n91 B 0.147534f
C313 VTAIL.t0 B 0.387168f
C314 VTAIL.t10 B 0.387168f
C315 VTAIL.n92 B 3.4357f
C316 VTAIL.n93 B 2.19629f
C317 VTAIL.t4 B 0.387168f
C318 VTAIL.t5 B 0.387168f
C319 VTAIL.n94 B 3.43571f
C320 VTAIL.n95 B 2.19627f
C321 VTAIL.n96 B 0.044101f
C322 VTAIL.n97 B 0.030076f
C323 VTAIL.n98 B 0.016162f
C324 VTAIL.n99 B 0.0382f
C325 VTAIL.n100 B 0.017112f
C326 VTAIL.n101 B 0.030076f
C327 VTAIL.n102 B 0.016637f
C328 VTAIL.n103 B 0.0382f
C329 VTAIL.n104 B 0.016162f
C330 VTAIL.n105 B 0.017112f
C331 VTAIL.n106 B 0.030076f
C332 VTAIL.n107 B 0.016162f
C333 VTAIL.n108 B 0.0382f
C334 VTAIL.n109 B 0.017112f
C335 VTAIL.n110 B 0.030076f
C336 VTAIL.n111 B 0.016162f
C337 VTAIL.n112 B 0.0382f
C338 VTAIL.n113 B 0.017112f
C339 VTAIL.n114 B 0.030076f
C340 VTAIL.n115 B 0.016162f
C341 VTAIL.n116 B 0.0382f
C342 VTAIL.n117 B 0.017112f
C343 VTAIL.n118 B 0.030076f
C344 VTAIL.n119 B 0.016162f
C345 VTAIL.n120 B 0.0382f
C346 VTAIL.n121 B 0.017112f
C347 VTAIL.n122 B 0.030076f
C348 VTAIL.n123 B 0.016162f
C349 VTAIL.n124 B 0.02865f
C350 VTAIL.n125 B 0.022566f
C351 VTAIL.t7 B 0.063121f
C352 VTAIL.n126 B 0.205892f
C353 VTAIL.n127 B 2.13462f
C354 VTAIL.n128 B 0.016162f
C355 VTAIL.n129 B 0.017112f
C356 VTAIL.n130 B 0.0382f
C357 VTAIL.n131 B 0.0382f
C358 VTAIL.n132 B 0.017112f
C359 VTAIL.n133 B 0.016162f
C360 VTAIL.n134 B 0.030076f
C361 VTAIL.n135 B 0.030076f
C362 VTAIL.n136 B 0.016162f
C363 VTAIL.n137 B 0.017112f
C364 VTAIL.n138 B 0.0382f
C365 VTAIL.n139 B 0.0382f
C366 VTAIL.n140 B 0.017112f
C367 VTAIL.n141 B 0.016162f
C368 VTAIL.n142 B 0.030076f
C369 VTAIL.n143 B 0.030076f
C370 VTAIL.n144 B 0.016162f
C371 VTAIL.n145 B 0.017112f
C372 VTAIL.n146 B 0.0382f
C373 VTAIL.n147 B 0.0382f
C374 VTAIL.n148 B 0.017112f
C375 VTAIL.n149 B 0.016162f
C376 VTAIL.n150 B 0.030076f
C377 VTAIL.n151 B 0.030076f
C378 VTAIL.n152 B 0.016162f
C379 VTAIL.n153 B 0.017112f
C380 VTAIL.n154 B 0.0382f
C381 VTAIL.n155 B 0.0382f
C382 VTAIL.n156 B 0.017112f
C383 VTAIL.n157 B 0.016162f
C384 VTAIL.n158 B 0.030076f
C385 VTAIL.n159 B 0.030076f
C386 VTAIL.n160 B 0.016162f
C387 VTAIL.n161 B 0.017112f
C388 VTAIL.n162 B 0.0382f
C389 VTAIL.n163 B 0.0382f
C390 VTAIL.n164 B 0.017112f
C391 VTAIL.n165 B 0.016162f
C392 VTAIL.n166 B 0.030076f
C393 VTAIL.n167 B 0.030076f
C394 VTAIL.n168 B 0.016162f
C395 VTAIL.n169 B 0.017112f
C396 VTAIL.n170 B 0.0382f
C397 VTAIL.n171 B 0.0382f
C398 VTAIL.n172 B 0.0382f
C399 VTAIL.n173 B 0.016637f
C400 VTAIL.n174 B 0.016162f
C401 VTAIL.n175 B 0.030076f
C402 VTAIL.n176 B 0.030076f
C403 VTAIL.n177 B 0.016162f
C404 VTAIL.n178 B 0.017112f
C405 VTAIL.n179 B 0.0382f
C406 VTAIL.n180 B 0.085927f
C407 VTAIL.n181 B 0.017112f
C408 VTAIL.n182 B 0.016162f
C409 VTAIL.n183 B 0.078148f
C410 VTAIL.n184 B 0.048663f
C411 VTAIL.n185 B 0.147534f
C412 VTAIL.t2 B 0.387168f
C413 VTAIL.t11 B 0.387168f
C414 VTAIL.n186 B 3.43571f
C415 VTAIL.n187 B 0.400867f
C416 VTAIL.n188 B 0.044101f
C417 VTAIL.n189 B 0.030076f
C418 VTAIL.n190 B 0.016162f
C419 VTAIL.n191 B 0.0382f
C420 VTAIL.n192 B 0.017112f
C421 VTAIL.n193 B 0.030076f
C422 VTAIL.n194 B 0.016637f
C423 VTAIL.n195 B 0.0382f
C424 VTAIL.n196 B 0.016162f
C425 VTAIL.n197 B 0.017112f
C426 VTAIL.n198 B 0.030076f
C427 VTAIL.n199 B 0.016162f
C428 VTAIL.n200 B 0.0382f
C429 VTAIL.n201 B 0.017112f
C430 VTAIL.n202 B 0.030076f
C431 VTAIL.n203 B 0.016162f
C432 VTAIL.n204 B 0.0382f
C433 VTAIL.n205 B 0.017112f
C434 VTAIL.n206 B 0.030076f
C435 VTAIL.n207 B 0.016162f
C436 VTAIL.n208 B 0.0382f
C437 VTAIL.n209 B 0.017112f
C438 VTAIL.n210 B 0.030076f
C439 VTAIL.n211 B 0.016162f
C440 VTAIL.n212 B 0.0382f
C441 VTAIL.n213 B 0.017112f
C442 VTAIL.n214 B 0.030076f
C443 VTAIL.n215 B 0.016162f
C444 VTAIL.n216 B 0.02865f
C445 VTAIL.n217 B 0.022566f
C446 VTAIL.t3 B 0.063121f
C447 VTAIL.n218 B 0.205892f
C448 VTAIL.n219 B 2.13462f
C449 VTAIL.n220 B 0.016162f
C450 VTAIL.n221 B 0.017112f
C451 VTAIL.n222 B 0.0382f
C452 VTAIL.n223 B 0.0382f
C453 VTAIL.n224 B 0.017112f
C454 VTAIL.n225 B 0.016162f
C455 VTAIL.n226 B 0.030076f
C456 VTAIL.n227 B 0.030076f
C457 VTAIL.n228 B 0.016162f
C458 VTAIL.n229 B 0.017112f
C459 VTAIL.n230 B 0.0382f
C460 VTAIL.n231 B 0.0382f
C461 VTAIL.n232 B 0.017112f
C462 VTAIL.n233 B 0.016162f
C463 VTAIL.n234 B 0.030076f
C464 VTAIL.n235 B 0.030076f
C465 VTAIL.n236 B 0.016162f
C466 VTAIL.n237 B 0.017112f
C467 VTAIL.n238 B 0.0382f
C468 VTAIL.n239 B 0.0382f
C469 VTAIL.n240 B 0.017112f
C470 VTAIL.n241 B 0.016162f
C471 VTAIL.n242 B 0.030076f
C472 VTAIL.n243 B 0.030076f
C473 VTAIL.n244 B 0.016162f
C474 VTAIL.n245 B 0.017112f
C475 VTAIL.n246 B 0.0382f
C476 VTAIL.n247 B 0.0382f
C477 VTAIL.n248 B 0.017112f
C478 VTAIL.n249 B 0.016162f
C479 VTAIL.n250 B 0.030076f
C480 VTAIL.n251 B 0.030076f
C481 VTAIL.n252 B 0.016162f
C482 VTAIL.n253 B 0.017112f
C483 VTAIL.n254 B 0.0382f
C484 VTAIL.n255 B 0.0382f
C485 VTAIL.n256 B 0.017112f
C486 VTAIL.n257 B 0.016162f
C487 VTAIL.n258 B 0.030076f
C488 VTAIL.n259 B 0.030076f
C489 VTAIL.n260 B 0.016162f
C490 VTAIL.n261 B 0.017112f
C491 VTAIL.n262 B 0.0382f
C492 VTAIL.n263 B 0.0382f
C493 VTAIL.n264 B 0.0382f
C494 VTAIL.n265 B 0.016637f
C495 VTAIL.n266 B 0.016162f
C496 VTAIL.n267 B 0.030076f
C497 VTAIL.n268 B 0.030076f
C498 VTAIL.n269 B 0.016162f
C499 VTAIL.n270 B 0.017112f
C500 VTAIL.n271 B 0.0382f
C501 VTAIL.n272 B 0.085927f
C502 VTAIL.n273 B 0.017112f
C503 VTAIL.n274 B 0.016162f
C504 VTAIL.n275 B 0.078148f
C505 VTAIL.n276 B 0.048663f
C506 VTAIL.n277 B 1.89532f
C507 VTAIL.n278 B 0.044101f
C508 VTAIL.n279 B 0.030076f
C509 VTAIL.n280 B 0.016162f
C510 VTAIL.n281 B 0.0382f
C511 VTAIL.n282 B 0.017112f
C512 VTAIL.n283 B 0.030076f
C513 VTAIL.n284 B 0.016637f
C514 VTAIL.n285 B 0.0382f
C515 VTAIL.n286 B 0.017112f
C516 VTAIL.n287 B 0.030076f
C517 VTAIL.n288 B 0.016162f
C518 VTAIL.n289 B 0.0382f
C519 VTAIL.n290 B 0.017112f
C520 VTAIL.n291 B 0.030076f
C521 VTAIL.n292 B 0.016162f
C522 VTAIL.n293 B 0.0382f
C523 VTAIL.n294 B 0.017112f
C524 VTAIL.n295 B 0.030076f
C525 VTAIL.n296 B 0.016162f
C526 VTAIL.n297 B 0.0382f
C527 VTAIL.n298 B 0.017112f
C528 VTAIL.n299 B 0.030076f
C529 VTAIL.n300 B 0.016162f
C530 VTAIL.n301 B 0.0382f
C531 VTAIL.n302 B 0.017112f
C532 VTAIL.n303 B 0.030076f
C533 VTAIL.n304 B 0.016162f
C534 VTAIL.n305 B 0.02865f
C535 VTAIL.n306 B 0.022566f
C536 VTAIL.t6 B 0.063121f
C537 VTAIL.n307 B 0.205892f
C538 VTAIL.n308 B 2.13462f
C539 VTAIL.n309 B 0.016162f
C540 VTAIL.n310 B 0.017112f
C541 VTAIL.n311 B 0.0382f
C542 VTAIL.n312 B 0.0382f
C543 VTAIL.n313 B 0.017112f
C544 VTAIL.n314 B 0.016162f
C545 VTAIL.n315 B 0.030076f
C546 VTAIL.n316 B 0.030076f
C547 VTAIL.n317 B 0.016162f
C548 VTAIL.n318 B 0.017112f
C549 VTAIL.n319 B 0.0382f
C550 VTAIL.n320 B 0.0382f
C551 VTAIL.n321 B 0.017112f
C552 VTAIL.n322 B 0.016162f
C553 VTAIL.n323 B 0.030076f
C554 VTAIL.n324 B 0.030076f
C555 VTAIL.n325 B 0.016162f
C556 VTAIL.n326 B 0.017112f
C557 VTAIL.n327 B 0.0382f
C558 VTAIL.n328 B 0.0382f
C559 VTAIL.n329 B 0.017112f
C560 VTAIL.n330 B 0.016162f
C561 VTAIL.n331 B 0.030076f
C562 VTAIL.n332 B 0.030076f
C563 VTAIL.n333 B 0.016162f
C564 VTAIL.n334 B 0.017112f
C565 VTAIL.n335 B 0.0382f
C566 VTAIL.n336 B 0.0382f
C567 VTAIL.n337 B 0.017112f
C568 VTAIL.n338 B 0.016162f
C569 VTAIL.n339 B 0.030076f
C570 VTAIL.n340 B 0.030076f
C571 VTAIL.n341 B 0.016162f
C572 VTAIL.n342 B 0.017112f
C573 VTAIL.n343 B 0.0382f
C574 VTAIL.n344 B 0.0382f
C575 VTAIL.n345 B 0.017112f
C576 VTAIL.n346 B 0.016162f
C577 VTAIL.n347 B 0.030076f
C578 VTAIL.n348 B 0.030076f
C579 VTAIL.n349 B 0.016162f
C580 VTAIL.n350 B 0.016162f
C581 VTAIL.n351 B 0.017112f
C582 VTAIL.n352 B 0.0382f
C583 VTAIL.n353 B 0.0382f
C584 VTAIL.n354 B 0.0382f
C585 VTAIL.n355 B 0.016637f
C586 VTAIL.n356 B 0.016162f
C587 VTAIL.n357 B 0.030076f
C588 VTAIL.n358 B 0.030076f
C589 VTAIL.n359 B 0.016162f
C590 VTAIL.n360 B 0.017112f
C591 VTAIL.n361 B 0.0382f
C592 VTAIL.n362 B 0.085927f
C593 VTAIL.n363 B 0.017112f
C594 VTAIL.n364 B 0.016162f
C595 VTAIL.n365 B 0.078148f
C596 VTAIL.n366 B 0.048663f
C597 VTAIL.n367 B 1.87777f
C598 VDD2.n0 B 0.043557f
C599 VDD2.n1 B 0.029705f
C600 VDD2.n2 B 0.015962f
C601 VDD2.n3 B 0.037729f
C602 VDD2.n4 B 0.016901f
C603 VDD2.n5 B 0.029705f
C604 VDD2.n6 B 0.016432f
C605 VDD2.n7 B 0.037729f
C606 VDD2.n8 B 0.016901f
C607 VDD2.n9 B 0.029705f
C608 VDD2.n10 B 0.015962f
C609 VDD2.n11 B 0.037729f
C610 VDD2.n12 B 0.016901f
C611 VDD2.n13 B 0.029705f
C612 VDD2.n14 B 0.015962f
C613 VDD2.n15 B 0.037729f
C614 VDD2.n16 B 0.016901f
C615 VDD2.n17 B 0.029705f
C616 VDD2.n18 B 0.015962f
C617 VDD2.n19 B 0.037729f
C618 VDD2.n20 B 0.016901f
C619 VDD2.n21 B 0.029705f
C620 VDD2.n22 B 0.015962f
C621 VDD2.n23 B 0.037729f
C622 VDD2.n24 B 0.016901f
C623 VDD2.n25 B 0.029705f
C624 VDD2.n26 B 0.015962f
C625 VDD2.n27 B 0.028297f
C626 VDD2.n28 B 0.022288f
C627 VDD2.t3 B 0.062342f
C628 VDD2.n29 B 0.203352f
C629 VDD2.n30 B 2.10829f
C630 VDD2.n31 B 0.015962f
C631 VDD2.n32 B 0.016901f
C632 VDD2.n33 B 0.037729f
C633 VDD2.n34 B 0.037729f
C634 VDD2.n35 B 0.016901f
C635 VDD2.n36 B 0.015962f
C636 VDD2.n37 B 0.029705f
C637 VDD2.n38 B 0.029705f
C638 VDD2.n39 B 0.015962f
C639 VDD2.n40 B 0.016901f
C640 VDD2.n41 B 0.037729f
C641 VDD2.n42 B 0.037729f
C642 VDD2.n43 B 0.016901f
C643 VDD2.n44 B 0.015962f
C644 VDD2.n45 B 0.029705f
C645 VDD2.n46 B 0.029705f
C646 VDD2.n47 B 0.015962f
C647 VDD2.n48 B 0.016901f
C648 VDD2.n49 B 0.037729f
C649 VDD2.n50 B 0.037729f
C650 VDD2.n51 B 0.016901f
C651 VDD2.n52 B 0.015962f
C652 VDD2.n53 B 0.029705f
C653 VDD2.n54 B 0.029705f
C654 VDD2.n55 B 0.015962f
C655 VDD2.n56 B 0.016901f
C656 VDD2.n57 B 0.037729f
C657 VDD2.n58 B 0.037729f
C658 VDD2.n59 B 0.016901f
C659 VDD2.n60 B 0.015962f
C660 VDD2.n61 B 0.029705f
C661 VDD2.n62 B 0.029705f
C662 VDD2.n63 B 0.015962f
C663 VDD2.n64 B 0.016901f
C664 VDD2.n65 B 0.037729f
C665 VDD2.n66 B 0.037729f
C666 VDD2.n67 B 0.016901f
C667 VDD2.n68 B 0.015962f
C668 VDD2.n69 B 0.029705f
C669 VDD2.n70 B 0.029705f
C670 VDD2.n71 B 0.015962f
C671 VDD2.n72 B 0.015962f
C672 VDD2.n73 B 0.016901f
C673 VDD2.n74 B 0.037729f
C674 VDD2.n75 B 0.037729f
C675 VDD2.n76 B 0.037729f
C676 VDD2.n77 B 0.016432f
C677 VDD2.n78 B 0.015962f
C678 VDD2.n79 B 0.029705f
C679 VDD2.n80 B 0.029705f
C680 VDD2.n81 B 0.015962f
C681 VDD2.n82 B 0.016901f
C682 VDD2.n83 B 0.037729f
C683 VDD2.n84 B 0.084867f
C684 VDD2.n85 B 0.016901f
C685 VDD2.n86 B 0.015962f
C686 VDD2.n87 B 0.077184f
C687 VDD2.n88 B 0.06907f
C688 VDD2.t4 B 0.382392f
C689 VDD2.t1 B 0.382392f
C690 VDD2.n89 B 3.47469f
C691 VDD2.n90 B 2.27458f
C692 VDD2.n91 B 0.043557f
C693 VDD2.n92 B 0.029705f
C694 VDD2.n93 B 0.015962f
C695 VDD2.n94 B 0.037729f
C696 VDD2.n95 B 0.016901f
C697 VDD2.n96 B 0.029705f
C698 VDD2.n97 B 0.016432f
C699 VDD2.n98 B 0.037729f
C700 VDD2.n99 B 0.015962f
C701 VDD2.n100 B 0.016901f
C702 VDD2.n101 B 0.029705f
C703 VDD2.n102 B 0.015962f
C704 VDD2.n103 B 0.037729f
C705 VDD2.n104 B 0.016901f
C706 VDD2.n105 B 0.029705f
C707 VDD2.n106 B 0.015962f
C708 VDD2.n107 B 0.037729f
C709 VDD2.n108 B 0.016901f
C710 VDD2.n109 B 0.029705f
C711 VDD2.n110 B 0.015962f
C712 VDD2.n111 B 0.037729f
C713 VDD2.n112 B 0.016901f
C714 VDD2.n113 B 0.029705f
C715 VDD2.n114 B 0.015962f
C716 VDD2.n115 B 0.037729f
C717 VDD2.n116 B 0.016901f
C718 VDD2.n117 B 0.029705f
C719 VDD2.n118 B 0.015962f
C720 VDD2.n119 B 0.028297f
C721 VDD2.n120 B 0.022288f
C722 VDD2.t0 B 0.062342f
C723 VDD2.n121 B 0.203352f
C724 VDD2.n122 B 2.10829f
C725 VDD2.n123 B 0.015962f
C726 VDD2.n124 B 0.016901f
C727 VDD2.n125 B 0.037729f
C728 VDD2.n126 B 0.037729f
C729 VDD2.n127 B 0.016901f
C730 VDD2.n128 B 0.015962f
C731 VDD2.n129 B 0.029705f
C732 VDD2.n130 B 0.029705f
C733 VDD2.n131 B 0.015962f
C734 VDD2.n132 B 0.016901f
C735 VDD2.n133 B 0.037729f
C736 VDD2.n134 B 0.037729f
C737 VDD2.n135 B 0.016901f
C738 VDD2.n136 B 0.015962f
C739 VDD2.n137 B 0.029705f
C740 VDD2.n138 B 0.029705f
C741 VDD2.n139 B 0.015962f
C742 VDD2.n140 B 0.016901f
C743 VDD2.n141 B 0.037729f
C744 VDD2.n142 B 0.037729f
C745 VDD2.n143 B 0.016901f
C746 VDD2.n144 B 0.015962f
C747 VDD2.n145 B 0.029705f
C748 VDD2.n146 B 0.029705f
C749 VDD2.n147 B 0.015962f
C750 VDD2.n148 B 0.016901f
C751 VDD2.n149 B 0.037729f
C752 VDD2.n150 B 0.037729f
C753 VDD2.n151 B 0.016901f
C754 VDD2.n152 B 0.015962f
C755 VDD2.n153 B 0.029705f
C756 VDD2.n154 B 0.029705f
C757 VDD2.n155 B 0.015962f
C758 VDD2.n156 B 0.016901f
C759 VDD2.n157 B 0.037729f
C760 VDD2.n158 B 0.037729f
C761 VDD2.n159 B 0.016901f
C762 VDD2.n160 B 0.015962f
C763 VDD2.n161 B 0.029705f
C764 VDD2.n162 B 0.029705f
C765 VDD2.n163 B 0.015962f
C766 VDD2.n164 B 0.016901f
C767 VDD2.n165 B 0.037729f
C768 VDD2.n166 B 0.037729f
C769 VDD2.n167 B 0.037729f
C770 VDD2.n168 B 0.016432f
C771 VDD2.n169 B 0.015962f
C772 VDD2.n170 B 0.029705f
C773 VDD2.n171 B 0.029705f
C774 VDD2.n172 B 0.015962f
C775 VDD2.n173 B 0.016901f
C776 VDD2.n174 B 0.037729f
C777 VDD2.n175 B 0.084867f
C778 VDD2.n176 B 0.016901f
C779 VDD2.n177 B 0.015962f
C780 VDD2.n178 B 0.077184f
C781 VDD2.n179 B 0.068515f
C782 VDD2.n180 B 2.68052f
C783 VDD2.t2 B 0.382392f
C784 VDD2.t5 B 0.382392f
C785 VDD2.n181 B 3.47467f
C786 VN.t1 B 0.66308f
C787 VN.n0 B 0.271322f
C788 VN.t0 B 0.656498f
C789 VN.n1 B 0.253295f
C790 VN.t3 B 0.66308f
C791 VN.n2 B 0.271236f
C792 VN.n3 B 0.119546f
C793 VN.t2 B 0.66308f
C794 VN.n4 B 0.271322f
C795 VN.t5 B 0.66308f
C796 VN.t4 B 0.656498f
C797 VN.n5 B 0.253295f
C798 VN.n6 B 0.271236f
C799 VN.n7 B 2.64365f
.ends

