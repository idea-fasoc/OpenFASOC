* NGSPICE file created from diff_pair_sample_0577.ext - technology: sky130A

.subckt diff_pair_sample_0577 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t5 VP.t0 VTAIL.t9 B.t0 sky130_fd_pr__nfet_01v8 ad=0.8877 pd=5.71 as=2.0982 ps=11.54 w=5.38 l=0.52
X1 VDD2.t5 VN.t0 VTAIL.t11 B.t5 sky130_fd_pr__nfet_01v8 ad=2.0982 pd=11.54 as=0.8877 ps=5.71 w=5.38 l=0.52
X2 VDD1.t4 VP.t1 VTAIL.t6 B.t3 sky130_fd_pr__nfet_01v8 ad=0.8877 pd=5.71 as=2.0982 ps=11.54 w=5.38 l=0.52
X3 VTAIL.t7 VP.t2 VDD1.t3 B.t4 sky130_fd_pr__nfet_01v8 ad=0.8877 pd=5.71 as=0.8877 ps=5.71 w=5.38 l=0.52
X4 B.t19 B.t17 B.t18 B.t7 sky130_fd_pr__nfet_01v8 ad=2.0982 pd=11.54 as=0 ps=0 w=5.38 l=0.52
X5 B.t16 B.t14 B.t15 B.t11 sky130_fd_pr__nfet_01v8 ad=2.0982 pd=11.54 as=0 ps=0 w=5.38 l=0.52
X6 B.t13 B.t10 B.t12 B.t11 sky130_fd_pr__nfet_01v8 ad=2.0982 pd=11.54 as=0 ps=0 w=5.38 l=0.52
X7 VDD2.t4 VN.t1 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=0.8877 pd=5.71 as=2.0982 ps=11.54 w=5.38 l=0.52
X8 VTAIL.t4 VN.t2 VDD2.t3 B.t4 sky130_fd_pr__nfet_01v8 ad=0.8877 pd=5.71 as=0.8877 ps=5.71 w=5.38 l=0.52
X9 VTAIL.t8 VP.t3 VDD1.t2 B.t1 sky130_fd_pr__nfet_01v8 ad=0.8877 pd=5.71 as=0.8877 ps=5.71 w=5.38 l=0.52
X10 B.t9 B.t6 B.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=2.0982 pd=11.54 as=0 ps=0 w=5.38 l=0.52
X11 VDD2.t2 VN.t3 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=2.0982 pd=11.54 as=0.8877 ps=5.71 w=5.38 l=0.52
X12 VTAIL.t1 VN.t4 VDD2.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=0.8877 pd=5.71 as=0.8877 ps=5.71 w=5.38 l=0.52
X13 VDD2.t0 VN.t5 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=0.8877 pd=5.71 as=2.0982 ps=11.54 w=5.38 l=0.52
X14 VDD1.t1 VP.t4 VTAIL.t10 B.t2 sky130_fd_pr__nfet_01v8 ad=2.0982 pd=11.54 as=0.8877 ps=5.71 w=5.38 l=0.52
X15 VDD1.t0 VP.t5 VTAIL.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=2.0982 pd=11.54 as=0.8877 ps=5.71 w=5.38 l=0.52
R0 VP.n1 VP.t5 351.709
R1 VP.n6 VP.t4 324.887
R2 VP.n7 VP.t3 324.887
R3 VP.n8 VP.t1 324.887
R4 VP.n3 VP.t0 324.887
R5 VP.n2 VP.t2 324.887
R6 VP.n9 VP.n8 161.3
R7 VP.n4 VP.n3 161.3
R8 VP.n6 VP.n5 161.3
R9 VP.n7 VP.n0 80.6037
R10 VP.n7 VP.n6 48.2005
R11 VP.n8 VP.n7 48.2005
R12 VP.n3 VP.n2 48.2005
R13 VP.n4 VP.n1 45.1367
R14 VP.n5 VP.n4 35.4891
R15 VP.n2 VP.n1 13.3799
R16 VP.n5 VP.n0 0.285035
R17 VP.n9 VP.n0 0.285035
R18 VP VP.n9 0.0516364
R19 VTAIL.n114 VTAIL.n92 289.615
R20 VTAIL.n24 VTAIL.n2 289.615
R21 VTAIL.n86 VTAIL.n64 289.615
R22 VTAIL.n56 VTAIL.n34 289.615
R23 VTAIL.n100 VTAIL.n99 185
R24 VTAIL.n105 VTAIL.n104 185
R25 VTAIL.n107 VTAIL.n106 185
R26 VTAIL.n96 VTAIL.n95 185
R27 VTAIL.n113 VTAIL.n112 185
R28 VTAIL.n115 VTAIL.n114 185
R29 VTAIL.n10 VTAIL.n9 185
R30 VTAIL.n15 VTAIL.n14 185
R31 VTAIL.n17 VTAIL.n16 185
R32 VTAIL.n6 VTAIL.n5 185
R33 VTAIL.n23 VTAIL.n22 185
R34 VTAIL.n25 VTAIL.n24 185
R35 VTAIL.n87 VTAIL.n86 185
R36 VTAIL.n85 VTAIL.n84 185
R37 VTAIL.n68 VTAIL.n67 185
R38 VTAIL.n79 VTAIL.n78 185
R39 VTAIL.n77 VTAIL.n76 185
R40 VTAIL.n72 VTAIL.n71 185
R41 VTAIL.n57 VTAIL.n56 185
R42 VTAIL.n55 VTAIL.n54 185
R43 VTAIL.n38 VTAIL.n37 185
R44 VTAIL.n49 VTAIL.n48 185
R45 VTAIL.n47 VTAIL.n46 185
R46 VTAIL.n42 VTAIL.n41 185
R47 VTAIL.n101 VTAIL.t0 147.672
R48 VTAIL.n11 VTAIL.t6 147.672
R49 VTAIL.n73 VTAIL.t9 147.672
R50 VTAIL.n43 VTAIL.t3 147.672
R51 VTAIL.n105 VTAIL.n99 104.615
R52 VTAIL.n106 VTAIL.n105 104.615
R53 VTAIL.n106 VTAIL.n95 104.615
R54 VTAIL.n113 VTAIL.n95 104.615
R55 VTAIL.n114 VTAIL.n113 104.615
R56 VTAIL.n15 VTAIL.n9 104.615
R57 VTAIL.n16 VTAIL.n15 104.615
R58 VTAIL.n16 VTAIL.n5 104.615
R59 VTAIL.n23 VTAIL.n5 104.615
R60 VTAIL.n24 VTAIL.n23 104.615
R61 VTAIL.n86 VTAIL.n85 104.615
R62 VTAIL.n85 VTAIL.n67 104.615
R63 VTAIL.n78 VTAIL.n67 104.615
R64 VTAIL.n78 VTAIL.n77 104.615
R65 VTAIL.n77 VTAIL.n71 104.615
R66 VTAIL.n56 VTAIL.n55 104.615
R67 VTAIL.n55 VTAIL.n37 104.615
R68 VTAIL.n48 VTAIL.n37 104.615
R69 VTAIL.n48 VTAIL.n47 104.615
R70 VTAIL.n47 VTAIL.n41 104.615
R71 VTAIL.n63 VTAIL.n62 53.9159
R72 VTAIL.n33 VTAIL.n32 53.9159
R73 VTAIL.n1 VTAIL.n0 53.9157
R74 VTAIL.n31 VTAIL.n30 53.9157
R75 VTAIL.t0 VTAIL.n99 52.3082
R76 VTAIL.t6 VTAIL.n9 52.3082
R77 VTAIL.t9 VTAIL.n71 52.3082
R78 VTAIL.t3 VTAIL.n41 52.3082
R79 VTAIL.n119 VTAIL.n118 34.1247
R80 VTAIL.n29 VTAIL.n28 34.1247
R81 VTAIL.n91 VTAIL.n90 34.1247
R82 VTAIL.n61 VTAIL.n60 34.1247
R83 VTAIL.n33 VTAIL.n31 18.4703
R84 VTAIL.n119 VTAIL.n91 17.7376
R85 VTAIL.n101 VTAIL.n100 15.6666
R86 VTAIL.n11 VTAIL.n10 15.6666
R87 VTAIL.n73 VTAIL.n72 15.6666
R88 VTAIL.n43 VTAIL.n42 15.6666
R89 VTAIL.n104 VTAIL.n103 12.8005
R90 VTAIL.n14 VTAIL.n13 12.8005
R91 VTAIL.n76 VTAIL.n75 12.8005
R92 VTAIL.n46 VTAIL.n45 12.8005
R93 VTAIL.n107 VTAIL.n98 12.0247
R94 VTAIL.n17 VTAIL.n8 12.0247
R95 VTAIL.n79 VTAIL.n70 12.0247
R96 VTAIL.n49 VTAIL.n40 12.0247
R97 VTAIL.n108 VTAIL.n96 11.249
R98 VTAIL.n18 VTAIL.n6 11.249
R99 VTAIL.n80 VTAIL.n68 11.249
R100 VTAIL.n50 VTAIL.n38 11.249
R101 VTAIL.n112 VTAIL.n111 10.4732
R102 VTAIL.n22 VTAIL.n21 10.4732
R103 VTAIL.n84 VTAIL.n83 10.4732
R104 VTAIL.n54 VTAIL.n53 10.4732
R105 VTAIL.n115 VTAIL.n94 9.69747
R106 VTAIL.n25 VTAIL.n4 9.69747
R107 VTAIL.n87 VTAIL.n66 9.69747
R108 VTAIL.n57 VTAIL.n36 9.69747
R109 VTAIL.n118 VTAIL.n117 9.45567
R110 VTAIL.n28 VTAIL.n27 9.45567
R111 VTAIL.n90 VTAIL.n89 9.45567
R112 VTAIL.n60 VTAIL.n59 9.45567
R113 VTAIL.n117 VTAIL.n116 9.3005
R114 VTAIL.n94 VTAIL.n93 9.3005
R115 VTAIL.n111 VTAIL.n110 9.3005
R116 VTAIL.n109 VTAIL.n108 9.3005
R117 VTAIL.n98 VTAIL.n97 9.3005
R118 VTAIL.n103 VTAIL.n102 9.3005
R119 VTAIL.n27 VTAIL.n26 9.3005
R120 VTAIL.n4 VTAIL.n3 9.3005
R121 VTAIL.n21 VTAIL.n20 9.3005
R122 VTAIL.n19 VTAIL.n18 9.3005
R123 VTAIL.n8 VTAIL.n7 9.3005
R124 VTAIL.n13 VTAIL.n12 9.3005
R125 VTAIL.n89 VTAIL.n88 9.3005
R126 VTAIL.n66 VTAIL.n65 9.3005
R127 VTAIL.n83 VTAIL.n82 9.3005
R128 VTAIL.n81 VTAIL.n80 9.3005
R129 VTAIL.n70 VTAIL.n69 9.3005
R130 VTAIL.n75 VTAIL.n74 9.3005
R131 VTAIL.n59 VTAIL.n58 9.3005
R132 VTAIL.n36 VTAIL.n35 9.3005
R133 VTAIL.n53 VTAIL.n52 9.3005
R134 VTAIL.n51 VTAIL.n50 9.3005
R135 VTAIL.n40 VTAIL.n39 9.3005
R136 VTAIL.n45 VTAIL.n44 9.3005
R137 VTAIL.n116 VTAIL.n92 8.92171
R138 VTAIL.n26 VTAIL.n2 8.92171
R139 VTAIL.n88 VTAIL.n64 8.92171
R140 VTAIL.n58 VTAIL.n34 8.92171
R141 VTAIL.n118 VTAIL.n92 5.04292
R142 VTAIL.n28 VTAIL.n2 5.04292
R143 VTAIL.n90 VTAIL.n64 5.04292
R144 VTAIL.n60 VTAIL.n34 5.04292
R145 VTAIL.n102 VTAIL.n101 4.38687
R146 VTAIL.n12 VTAIL.n11 4.38687
R147 VTAIL.n74 VTAIL.n73 4.38687
R148 VTAIL.n44 VTAIL.n43 4.38687
R149 VTAIL.n116 VTAIL.n115 4.26717
R150 VTAIL.n26 VTAIL.n25 4.26717
R151 VTAIL.n88 VTAIL.n87 4.26717
R152 VTAIL.n58 VTAIL.n57 4.26717
R153 VTAIL.n0 VTAIL.t11 3.6808
R154 VTAIL.n0 VTAIL.t4 3.6808
R155 VTAIL.n30 VTAIL.t10 3.6808
R156 VTAIL.n30 VTAIL.t8 3.6808
R157 VTAIL.n62 VTAIL.t5 3.6808
R158 VTAIL.n62 VTAIL.t7 3.6808
R159 VTAIL.n32 VTAIL.t2 3.6808
R160 VTAIL.n32 VTAIL.t1 3.6808
R161 VTAIL.n112 VTAIL.n94 3.49141
R162 VTAIL.n22 VTAIL.n4 3.49141
R163 VTAIL.n84 VTAIL.n66 3.49141
R164 VTAIL.n54 VTAIL.n36 3.49141
R165 VTAIL.n111 VTAIL.n96 2.71565
R166 VTAIL.n21 VTAIL.n6 2.71565
R167 VTAIL.n83 VTAIL.n68 2.71565
R168 VTAIL.n53 VTAIL.n38 2.71565
R169 VTAIL.n108 VTAIL.n107 1.93989
R170 VTAIL.n18 VTAIL.n17 1.93989
R171 VTAIL.n80 VTAIL.n79 1.93989
R172 VTAIL.n50 VTAIL.n49 1.93989
R173 VTAIL.n104 VTAIL.n98 1.16414
R174 VTAIL.n14 VTAIL.n8 1.16414
R175 VTAIL.n76 VTAIL.n70 1.16414
R176 VTAIL.n46 VTAIL.n40 1.16414
R177 VTAIL.n63 VTAIL.n61 0.836707
R178 VTAIL.n29 VTAIL.n1 0.836707
R179 VTAIL.n61 VTAIL.n33 0.733259
R180 VTAIL.n91 VTAIL.n63 0.733259
R181 VTAIL.n31 VTAIL.n29 0.733259
R182 VTAIL VTAIL.n119 0.491879
R183 VTAIL.n103 VTAIL.n100 0.388379
R184 VTAIL.n13 VTAIL.n10 0.388379
R185 VTAIL.n75 VTAIL.n72 0.388379
R186 VTAIL.n45 VTAIL.n42 0.388379
R187 VTAIL VTAIL.n1 0.241879
R188 VTAIL.n102 VTAIL.n97 0.155672
R189 VTAIL.n109 VTAIL.n97 0.155672
R190 VTAIL.n110 VTAIL.n109 0.155672
R191 VTAIL.n110 VTAIL.n93 0.155672
R192 VTAIL.n117 VTAIL.n93 0.155672
R193 VTAIL.n12 VTAIL.n7 0.155672
R194 VTAIL.n19 VTAIL.n7 0.155672
R195 VTAIL.n20 VTAIL.n19 0.155672
R196 VTAIL.n20 VTAIL.n3 0.155672
R197 VTAIL.n27 VTAIL.n3 0.155672
R198 VTAIL.n89 VTAIL.n65 0.155672
R199 VTAIL.n82 VTAIL.n65 0.155672
R200 VTAIL.n82 VTAIL.n81 0.155672
R201 VTAIL.n81 VTAIL.n69 0.155672
R202 VTAIL.n74 VTAIL.n69 0.155672
R203 VTAIL.n59 VTAIL.n35 0.155672
R204 VTAIL.n52 VTAIL.n35 0.155672
R205 VTAIL.n52 VTAIL.n51 0.155672
R206 VTAIL.n51 VTAIL.n39 0.155672
R207 VTAIL.n44 VTAIL.n39 0.155672
R208 VDD1.n22 VDD1.n0 289.615
R209 VDD1.n49 VDD1.n27 289.615
R210 VDD1.n23 VDD1.n22 185
R211 VDD1.n21 VDD1.n20 185
R212 VDD1.n4 VDD1.n3 185
R213 VDD1.n15 VDD1.n14 185
R214 VDD1.n13 VDD1.n12 185
R215 VDD1.n8 VDD1.n7 185
R216 VDD1.n35 VDD1.n34 185
R217 VDD1.n40 VDD1.n39 185
R218 VDD1.n42 VDD1.n41 185
R219 VDD1.n31 VDD1.n30 185
R220 VDD1.n48 VDD1.n47 185
R221 VDD1.n50 VDD1.n49 185
R222 VDD1.n9 VDD1.t0 147.672
R223 VDD1.n36 VDD1.t1 147.672
R224 VDD1.n22 VDD1.n21 104.615
R225 VDD1.n21 VDD1.n3 104.615
R226 VDD1.n14 VDD1.n3 104.615
R227 VDD1.n14 VDD1.n13 104.615
R228 VDD1.n13 VDD1.n7 104.615
R229 VDD1.n40 VDD1.n34 104.615
R230 VDD1.n41 VDD1.n40 104.615
R231 VDD1.n41 VDD1.n30 104.615
R232 VDD1.n48 VDD1.n30 104.615
R233 VDD1.n49 VDD1.n48 104.615
R234 VDD1.n55 VDD1.n54 70.7223
R235 VDD1.n57 VDD1.n56 70.5945
R236 VDD1.t0 VDD1.n7 52.3082
R237 VDD1.t1 VDD1.n34 52.3082
R238 VDD1 VDD1.n26 51.4113
R239 VDD1.n55 VDD1.n53 51.2978
R240 VDD1.n57 VDD1.n55 31.6841
R241 VDD1.n9 VDD1.n8 15.6666
R242 VDD1.n36 VDD1.n35 15.6666
R243 VDD1.n12 VDD1.n11 12.8005
R244 VDD1.n39 VDD1.n38 12.8005
R245 VDD1.n15 VDD1.n6 12.0247
R246 VDD1.n42 VDD1.n33 12.0247
R247 VDD1.n16 VDD1.n4 11.249
R248 VDD1.n43 VDD1.n31 11.249
R249 VDD1.n20 VDD1.n19 10.4732
R250 VDD1.n47 VDD1.n46 10.4732
R251 VDD1.n23 VDD1.n2 9.69747
R252 VDD1.n50 VDD1.n29 9.69747
R253 VDD1.n26 VDD1.n25 9.45567
R254 VDD1.n53 VDD1.n52 9.45567
R255 VDD1.n25 VDD1.n24 9.3005
R256 VDD1.n2 VDD1.n1 9.3005
R257 VDD1.n19 VDD1.n18 9.3005
R258 VDD1.n17 VDD1.n16 9.3005
R259 VDD1.n6 VDD1.n5 9.3005
R260 VDD1.n11 VDD1.n10 9.3005
R261 VDD1.n52 VDD1.n51 9.3005
R262 VDD1.n29 VDD1.n28 9.3005
R263 VDD1.n46 VDD1.n45 9.3005
R264 VDD1.n44 VDD1.n43 9.3005
R265 VDD1.n33 VDD1.n32 9.3005
R266 VDD1.n38 VDD1.n37 9.3005
R267 VDD1.n24 VDD1.n0 8.92171
R268 VDD1.n51 VDD1.n27 8.92171
R269 VDD1.n26 VDD1.n0 5.04292
R270 VDD1.n53 VDD1.n27 5.04292
R271 VDD1.n10 VDD1.n9 4.38687
R272 VDD1.n37 VDD1.n36 4.38687
R273 VDD1.n24 VDD1.n23 4.26717
R274 VDD1.n51 VDD1.n50 4.26717
R275 VDD1.n56 VDD1.t3 3.6808
R276 VDD1.n56 VDD1.t5 3.6808
R277 VDD1.n54 VDD1.t2 3.6808
R278 VDD1.n54 VDD1.t4 3.6808
R279 VDD1.n20 VDD1.n2 3.49141
R280 VDD1.n47 VDD1.n29 3.49141
R281 VDD1.n19 VDD1.n4 2.71565
R282 VDD1.n46 VDD1.n31 2.71565
R283 VDD1.n16 VDD1.n15 1.93989
R284 VDD1.n43 VDD1.n42 1.93989
R285 VDD1.n12 VDD1.n6 1.16414
R286 VDD1.n39 VDD1.n33 1.16414
R287 VDD1.n11 VDD1.n8 0.388379
R288 VDD1.n38 VDD1.n35 0.388379
R289 VDD1.n25 VDD1.n1 0.155672
R290 VDD1.n18 VDD1.n1 0.155672
R291 VDD1.n18 VDD1.n17 0.155672
R292 VDD1.n17 VDD1.n5 0.155672
R293 VDD1.n10 VDD1.n5 0.155672
R294 VDD1.n37 VDD1.n32 0.155672
R295 VDD1.n44 VDD1.n32 0.155672
R296 VDD1.n45 VDD1.n44 0.155672
R297 VDD1.n45 VDD1.n28 0.155672
R298 VDD1.n52 VDD1.n28 0.155672
R299 VDD1 VDD1.n57 0.1255
R300 B.n323 B.n322 585
R301 B.n324 B.n69 585
R302 B.n326 B.n325 585
R303 B.n328 B.n68 585
R304 B.n331 B.n330 585
R305 B.n332 B.n67 585
R306 B.n334 B.n333 585
R307 B.n336 B.n66 585
R308 B.n339 B.n338 585
R309 B.n340 B.n65 585
R310 B.n342 B.n341 585
R311 B.n344 B.n64 585
R312 B.n347 B.n346 585
R313 B.n348 B.n63 585
R314 B.n350 B.n349 585
R315 B.n352 B.n62 585
R316 B.n355 B.n354 585
R317 B.n356 B.n61 585
R318 B.n358 B.n357 585
R319 B.n360 B.n60 585
R320 B.n362 B.n361 585
R321 B.n364 B.n363 585
R322 B.n367 B.n366 585
R323 B.n368 B.n55 585
R324 B.n370 B.n369 585
R325 B.n372 B.n54 585
R326 B.n375 B.n374 585
R327 B.n376 B.n53 585
R328 B.n378 B.n377 585
R329 B.n380 B.n52 585
R330 B.n382 B.n381 585
R331 B.n384 B.n383 585
R332 B.n387 B.n386 585
R333 B.n388 B.n47 585
R334 B.n390 B.n389 585
R335 B.n392 B.n46 585
R336 B.n395 B.n394 585
R337 B.n396 B.n45 585
R338 B.n398 B.n397 585
R339 B.n400 B.n44 585
R340 B.n403 B.n402 585
R341 B.n404 B.n43 585
R342 B.n406 B.n405 585
R343 B.n408 B.n42 585
R344 B.n411 B.n410 585
R345 B.n412 B.n41 585
R346 B.n414 B.n413 585
R347 B.n416 B.n40 585
R348 B.n419 B.n418 585
R349 B.n420 B.n39 585
R350 B.n422 B.n421 585
R351 B.n424 B.n38 585
R352 B.n427 B.n426 585
R353 B.n428 B.n37 585
R354 B.n320 B.n35 585
R355 B.n431 B.n35 585
R356 B.n319 B.n34 585
R357 B.n432 B.n34 585
R358 B.n318 B.n33 585
R359 B.n433 B.n33 585
R360 B.n317 B.n316 585
R361 B.n316 B.n29 585
R362 B.n315 B.n28 585
R363 B.n439 B.n28 585
R364 B.n314 B.n27 585
R365 B.n440 B.n27 585
R366 B.n313 B.n26 585
R367 B.n441 B.n26 585
R368 B.n312 B.n311 585
R369 B.n311 B.n22 585
R370 B.n310 B.n21 585
R371 B.n447 B.n21 585
R372 B.n309 B.n20 585
R373 B.n448 B.n20 585
R374 B.n308 B.n19 585
R375 B.n449 B.n19 585
R376 B.n307 B.n306 585
R377 B.n306 B.n15 585
R378 B.n305 B.n14 585
R379 B.n455 B.n14 585
R380 B.n304 B.n13 585
R381 B.n456 B.n13 585
R382 B.n303 B.n12 585
R383 B.n457 B.n12 585
R384 B.n302 B.n301 585
R385 B.n301 B.n11 585
R386 B.n300 B.n7 585
R387 B.n463 B.n7 585
R388 B.n299 B.n6 585
R389 B.n464 B.n6 585
R390 B.n298 B.n5 585
R391 B.n465 B.n5 585
R392 B.n297 B.n296 585
R393 B.n296 B.n4 585
R394 B.n295 B.n70 585
R395 B.n295 B.n294 585
R396 B.n284 B.n71 585
R397 B.n287 B.n71 585
R398 B.n286 B.n285 585
R399 B.n288 B.n286 585
R400 B.n283 B.n76 585
R401 B.n76 B.n75 585
R402 B.n282 B.n281 585
R403 B.n281 B.n280 585
R404 B.n78 B.n77 585
R405 B.n79 B.n78 585
R406 B.n273 B.n272 585
R407 B.n274 B.n273 585
R408 B.n271 B.n84 585
R409 B.n84 B.n83 585
R410 B.n270 B.n269 585
R411 B.n269 B.n268 585
R412 B.n86 B.n85 585
R413 B.n87 B.n86 585
R414 B.n261 B.n260 585
R415 B.n262 B.n261 585
R416 B.n259 B.n92 585
R417 B.n92 B.n91 585
R418 B.n258 B.n257 585
R419 B.n257 B.n256 585
R420 B.n94 B.n93 585
R421 B.n95 B.n94 585
R422 B.n249 B.n248 585
R423 B.n250 B.n249 585
R424 B.n247 B.n100 585
R425 B.n100 B.n99 585
R426 B.n246 B.n245 585
R427 B.n245 B.n244 585
R428 B.n241 B.n104 585
R429 B.n240 B.n239 585
R430 B.n237 B.n105 585
R431 B.n237 B.n103 585
R432 B.n236 B.n235 585
R433 B.n234 B.n233 585
R434 B.n232 B.n107 585
R435 B.n230 B.n229 585
R436 B.n228 B.n108 585
R437 B.n227 B.n226 585
R438 B.n224 B.n109 585
R439 B.n222 B.n221 585
R440 B.n220 B.n110 585
R441 B.n219 B.n218 585
R442 B.n216 B.n111 585
R443 B.n214 B.n213 585
R444 B.n212 B.n112 585
R445 B.n211 B.n210 585
R446 B.n208 B.n113 585
R447 B.n206 B.n205 585
R448 B.n204 B.n114 585
R449 B.n203 B.n202 585
R450 B.n200 B.n115 585
R451 B.n198 B.n197 585
R452 B.n196 B.n116 585
R453 B.n195 B.n194 585
R454 B.n192 B.n120 585
R455 B.n190 B.n189 585
R456 B.n188 B.n121 585
R457 B.n187 B.n186 585
R458 B.n184 B.n122 585
R459 B.n182 B.n181 585
R460 B.n180 B.n123 585
R461 B.n178 B.n177 585
R462 B.n175 B.n126 585
R463 B.n173 B.n172 585
R464 B.n171 B.n127 585
R465 B.n170 B.n169 585
R466 B.n167 B.n128 585
R467 B.n165 B.n164 585
R468 B.n163 B.n129 585
R469 B.n162 B.n161 585
R470 B.n159 B.n130 585
R471 B.n157 B.n156 585
R472 B.n155 B.n131 585
R473 B.n154 B.n153 585
R474 B.n151 B.n132 585
R475 B.n149 B.n148 585
R476 B.n147 B.n133 585
R477 B.n146 B.n145 585
R478 B.n143 B.n134 585
R479 B.n141 B.n140 585
R480 B.n139 B.n135 585
R481 B.n138 B.n137 585
R482 B.n102 B.n101 585
R483 B.n103 B.n102 585
R484 B.n243 B.n242 585
R485 B.n244 B.n243 585
R486 B.n98 B.n97 585
R487 B.n99 B.n98 585
R488 B.n252 B.n251 585
R489 B.n251 B.n250 585
R490 B.n253 B.n96 585
R491 B.n96 B.n95 585
R492 B.n255 B.n254 585
R493 B.n256 B.n255 585
R494 B.n90 B.n89 585
R495 B.n91 B.n90 585
R496 B.n264 B.n263 585
R497 B.n263 B.n262 585
R498 B.n265 B.n88 585
R499 B.n88 B.n87 585
R500 B.n267 B.n266 585
R501 B.n268 B.n267 585
R502 B.n82 B.n81 585
R503 B.n83 B.n82 585
R504 B.n276 B.n275 585
R505 B.n275 B.n274 585
R506 B.n277 B.n80 585
R507 B.n80 B.n79 585
R508 B.n279 B.n278 585
R509 B.n280 B.n279 585
R510 B.n74 B.n73 585
R511 B.n75 B.n74 585
R512 B.n290 B.n289 585
R513 B.n289 B.n288 585
R514 B.n291 B.n72 585
R515 B.n287 B.n72 585
R516 B.n293 B.n292 585
R517 B.n294 B.n293 585
R518 B.n2 B.n0 585
R519 B.n4 B.n2 585
R520 B.n3 B.n1 585
R521 B.n464 B.n3 585
R522 B.n462 B.n461 585
R523 B.n463 B.n462 585
R524 B.n460 B.n8 585
R525 B.n11 B.n8 585
R526 B.n459 B.n458 585
R527 B.n458 B.n457 585
R528 B.n10 B.n9 585
R529 B.n456 B.n10 585
R530 B.n454 B.n453 585
R531 B.n455 B.n454 585
R532 B.n452 B.n16 585
R533 B.n16 B.n15 585
R534 B.n451 B.n450 585
R535 B.n450 B.n449 585
R536 B.n18 B.n17 585
R537 B.n448 B.n18 585
R538 B.n446 B.n445 585
R539 B.n447 B.n446 585
R540 B.n444 B.n23 585
R541 B.n23 B.n22 585
R542 B.n443 B.n442 585
R543 B.n442 B.n441 585
R544 B.n25 B.n24 585
R545 B.n440 B.n25 585
R546 B.n438 B.n437 585
R547 B.n439 B.n438 585
R548 B.n436 B.n30 585
R549 B.n30 B.n29 585
R550 B.n435 B.n434 585
R551 B.n434 B.n433 585
R552 B.n32 B.n31 585
R553 B.n432 B.n32 585
R554 B.n430 B.n429 585
R555 B.n431 B.n430 585
R556 B.n467 B.n466 585
R557 B.n466 B.n465 585
R558 B.n243 B.n104 506.916
R559 B.n430 B.n37 506.916
R560 B.n245 B.n102 506.916
R561 B.n322 B.n35 506.916
R562 B.n124 B.t14 455.286
R563 B.n117 B.t10 455.286
R564 B.n48 B.t6 455.286
R565 B.n56 B.t17 455.286
R566 B.n321 B.n36 256.663
R567 B.n327 B.n36 256.663
R568 B.n329 B.n36 256.663
R569 B.n335 B.n36 256.663
R570 B.n337 B.n36 256.663
R571 B.n343 B.n36 256.663
R572 B.n345 B.n36 256.663
R573 B.n351 B.n36 256.663
R574 B.n353 B.n36 256.663
R575 B.n359 B.n36 256.663
R576 B.n59 B.n36 256.663
R577 B.n365 B.n36 256.663
R578 B.n371 B.n36 256.663
R579 B.n373 B.n36 256.663
R580 B.n379 B.n36 256.663
R581 B.n51 B.n36 256.663
R582 B.n385 B.n36 256.663
R583 B.n391 B.n36 256.663
R584 B.n393 B.n36 256.663
R585 B.n399 B.n36 256.663
R586 B.n401 B.n36 256.663
R587 B.n407 B.n36 256.663
R588 B.n409 B.n36 256.663
R589 B.n415 B.n36 256.663
R590 B.n417 B.n36 256.663
R591 B.n423 B.n36 256.663
R592 B.n425 B.n36 256.663
R593 B.n238 B.n103 256.663
R594 B.n106 B.n103 256.663
R595 B.n231 B.n103 256.663
R596 B.n225 B.n103 256.663
R597 B.n223 B.n103 256.663
R598 B.n217 B.n103 256.663
R599 B.n215 B.n103 256.663
R600 B.n209 B.n103 256.663
R601 B.n207 B.n103 256.663
R602 B.n201 B.n103 256.663
R603 B.n199 B.n103 256.663
R604 B.n193 B.n103 256.663
R605 B.n191 B.n103 256.663
R606 B.n185 B.n103 256.663
R607 B.n183 B.n103 256.663
R608 B.n176 B.n103 256.663
R609 B.n174 B.n103 256.663
R610 B.n168 B.n103 256.663
R611 B.n166 B.n103 256.663
R612 B.n160 B.n103 256.663
R613 B.n158 B.n103 256.663
R614 B.n152 B.n103 256.663
R615 B.n150 B.n103 256.663
R616 B.n144 B.n103 256.663
R617 B.n142 B.n103 256.663
R618 B.n136 B.n103 256.663
R619 B.n124 B.t16 184.999
R620 B.n56 B.t18 184.999
R621 B.n117 B.t13 184.999
R622 B.n48 B.t8 184.999
R623 B.n125 B.t15 168.513
R624 B.n57 B.t19 168.513
R625 B.n118 B.t12 168.513
R626 B.n49 B.t9 168.513
R627 B.n243 B.n98 163.367
R628 B.n251 B.n98 163.367
R629 B.n251 B.n96 163.367
R630 B.n255 B.n96 163.367
R631 B.n255 B.n90 163.367
R632 B.n263 B.n90 163.367
R633 B.n263 B.n88 163.367
R634 B.n267 B.n88 163.367
R635 B.n267 B.n82 163.367
R636 B.n275 B.n82 163.367
R637 B.n275 B.n80 163.367
R638 B.n279 B.n80 163.367
R639 B.n279 B.n74 163.367
R640 B.n289 B.n74 163.367
R641 B.n289 B.n72 163.367
R642 B.n293 B.n72 163.367
R643 B.n293 B.n2 163.367
R644 B.n466 B.n2 163.367
R645 B.n466 B.n3 163.367
R646 B.n462 B.n3 163.367
R647 B.n462 B.n8 163.367
R648 B.n458 B.n8 163.367
R649 B.n458 B.n10 163.367
R650 B.n454 B.n10 163.367
R651 B.n454 B.n16 163.367
R652 B.n450 B.n16 163.367
R653 B.n450 B.n18 163.367
R654 B.n446 B.n18 163.367
R655 B.n446 B.n23 163.367
R656 B.n442 B.n23 163.367
R657 B.n442 B.n25 163.367
R658 B.n438 B.n25 163.367
R659 B.n438 B.n30 163.367
R660 B.n434 B.n30 163.367
R661 B.n434 B.n32 163.367
R662 B.n430 B.n32 163.367
R663 B.n239 B.n237 163.367
R664 B.n237 B.n236 163.367
R665 B.n233 B.n232 163.367
R666 B.n230 B.n108 163.367
R667 B.n226 B.n224 163.367
R668 B.n222 B.n110 163.367
R669 B.n218 B.n216 163.367
R670 B.n214 B.n112 163.367
R671 B.n210 B.n208 163.367
R672 B.n206 B.n114 163.367
R673 B.n202 B.n200 163.367
R674 B.n198 B.n116 163.367
R675 B.n194 B.n192 163.367
R676 B.n190 B.n121 163.367
R677 B.n186 B.n184 163.367
R678 B.n182 B.n123 163.367
R679 B.n177 B.n175 163.367
R680 B.n173 B.n127 163.367
R681 B.n169 B.n167 163.367
R682 B.n165 B.n129 163.367
R683 B.n161 B.n159 163.367
R684 B.n157 B.n131 163.367
R685 B.n153 B.n151 163.367
R686 B.n149 B.n133 163.367
R687 B.n145 B.n143 163.367
R688 B.n141 B.n135 163.367
R689 B.n137 B.n102 163.367
R690 B.n245 B.n100 163.367
R691 B.n249 B.n100 163.367
R692 B.n249 B.n94 163.367
R693 B.n257 B.n94 163.367
R694 B.n257 B.n92 163.367
R695 B.n261 B.n92 163.367
R696 B.n261 B.n86 163.367
R697 B.n269 B.n86 163.367
R698 B.n269 B.n84 163.367
R699 B.n273 B.n84 163.367
R700 B.n273 B.n78 163.367
R701 B.n281 B.n78 163.367
R702 B.n281 B.n76 163.367
R703 B.n286 B.n76 163.367
R704 B.n286 B.n71 163.367
R705 B.n295 B.n71 163.367
R706 B.n296 B.n295 163.367
R707 B.n296 B.n5 163.367
R708 B.n6 B.n5 163.367
R709 B.n7 B.n6 163.367
R710 B.n301 B.n7 163.367
R711 B.n301 B.n12 163.367
R712 B.n13 B.n12 163.367
R713 B.n14 B.n13 163.367
R714 B.n306 B.n14 163.367
R715 B.n306 B.n19 163.367
R716 B.n20 B.n19 163.367
R717 B.n21 B.n20 163.367
R718 B.n311 B.n21 163.367
R719 B.n311 B.n26 163.367
R720 B.n27 B.n26 163.367
R721 B.n28 B.n27 163.367
R722 B.n316 B.n28 163.367
R723 B.n316 B.n33 163.367
R724 B.n34 B.n33 163.367
R725 B.n35 B.n34 163.367
R726 B.n426 B.n424 163.367
R727 B.n422 B.n39 163.367
R728 B.n418 B.n416 163.367
R729 B.n414 B.n41 163.367
R730 B.n410 B.n408 163.367
R731 B.n406 B.n43 163.367
R732 B.n402 B.n400 163.367
R733 B.n398 B.n45 163.367
R734 B.n394 B.n392 163.367
R735 B.n390 B.n47 163.367
R736 B.n386 B.n384 163.367
R737 B.n381 B.n380 163.367
R738 B.n378 B.n53 163.367
R739 B.n374 B.n372 163.367
R740 B.n370 B.n55 163.367
R741 B.n366 B.n364 163.367
R742 B.n361 B.n360 163.367
R743 B.n358 B.n61 163.367
R744 B.n354 B.n352 163.367
R745 B.n350 B.n63 163.367
R746 B.n346 B.n344 163.367
R747 B.n342 B.n65 163.367
R748 B.n338 B.n336 163.367
R749 B.n334 B.n67 163.367
R750 B.n330 B.n328 163.367
R751 B.n326 B.n69 163.367
R752 B.n244 B.n103 135.243
R753 B.n431 B.n36 135.243
R754 B.n238 B.n104 71.676
R755 B.n236 B.n106 71.676
R756 B.n232 B.n231 71.676
R757 B.n225 B.n108 71.676
R758 B.n224 B.n223 71.676
R759 B.n217 B.n110 71.676
R760 B.n216 B.n215 71.676
R761 B.n209 B.n112 71.676
R762 B.n208 B.n207 71.676
R763 B.n201 B.n114 71.676
R764 B.n200 B.n199 71.676
R765 B.n193 B.n116 71.676
R766 B.n192 B.n191 71.676
R767 B.n185 B.n121 71.676
R768 B.n184 B.n183 71.676
R769 B.n176 B.n123 71.676
R770 B.n175 B.n174 71.676
R771 B.n168 B.n127 71.676
R772 B.n167 B.n166 71.676
R773 B.n160 B.n129 71.676
R774 B.n159 B.n158 71.676
R775 B.n152 B.n131 71.676
R776 B.n151 B.n150 71.676
R777 B.n144 B.n133 71.676
R778 B.n143 B.n142 71.676
R779 B.n136 B.n135 71.676
R780 B.n425 B.n37 71.676
R781 B.n424 B.n423 71.676
R782 B.n417 B.n39 71.676
R783 B.n416 B.n415 71.676
R784 B.n409 B.n41 71.676
R785 B.n408 B.n407 71.676
R786 B.n401 B.n43 71.676
R787 B.n400 B.n399 71.676
R788 B.n393 B.n45 71.676
R789 B.n392 B.n391 71.676
R790 B.n385 B.n47 71.676
R791 B.n384 B.n51 71.676
R792 B.n380 B.n379 71.676
R793 B.n373 B.n53 71.676
R794 B.n372 B.n371 71.676
R795 B.n365 B.n55 71.676
R796 B.n364 B.n59 71.676
R797 B.n360 B.n359 71.676
R798 B.n353 B.n61 71.676
R799 B.n352 B.n351 71.676
R800 B.n345 B.n63 71.676
R801 B.n344 B.n343 71.676
R802 B.n337 B.n65 71.676
R803 B.n336 B.n335 71.676
R804 B.n329 B.n67 71.676
R805 B.n328 B.n327 71.676
R806 B.n321 B.n69 71.676
R807 B.n322 B.n321 71.676
R808 B.n327 B.n326 71.676
R809 B.n330 B.n329 71.676
R810 B.n335 B.n334 71.676
R811 B.n338 B.n337 71.676
R812 B.n343 B.n342 71.676
R813 B.n346 B.n345 71.676
R814 B.n351 B.n350 71.676
R815 B.n354 B.n353 71.676
R816 B.n359 B.n358 71.676
R817 B.n361 B.n59 71.676
R818 B.n366 B.n365 71.676
R819 B.n371 B.n370 71.676
R820 B.n374 B.n373 71.676
R821 B.n379 B.n378 71.676
R822 B.n381 B.n51 71.676
R823 B.n386 B.n385 71.676
R824 B.n391 B.n390 71.676
R825 B.n394 B.n393 71.676
R826 B.n399 B.n398 71.676
R827 B.n402 B.n401 71.676
R828 B.n407 B.n406 71.676
R829 B.n410 B.n409 71.676
R830 B.n415 B.n414 71.676
R831 B.n418 B.n417 71.676
R832 B.n423 B.n422 71.676
R833 B.n426 B.n425 71.676
R834 B.n239 B.n238 71.676
R835 B.n233 B.n106 71.676
R836 B.n231 B.n230 71.676
R837 B.n226 B.n225 71.676
R838 B.n223 B.n222 71.676
R839 B.n218 B.n217 71.676
R840 B.n215 B.n214 71.676
R841 B.n210 B.n209 71.676
R842 B.n207 B.n206 71.676
R843 B.n202 B.n201 71.676
R844 B.n199 B.n198 71.676
R845 B.n194 B.n193 71.676
R846 B.n191 B.n190 71.676
R847 B.n186 B.n185 71.676
R848 B.n183 B.n182 71.676
R849 B.n177 B.n176 71.676
R850 B.n174 B.n173 71.676
R851 B.n169 B.n168 71.676
R852 B.n166 B.n165 71.676
R853 B.n161 B.n160 71.676
R854 B.n158 B.n157 71.676
R855 B.n153 B.n152 71.676
R856 B.n150 B.n149 71.676
R857 B.n145 B.n144 71.676
R858 B.n142 B.n141 71.676
R859 B.n137 B.n136 71.676
R860 B.n244 B.n99 70.2023
R861 B.n250 B.n99 70.2023
R862 B.n250 B.n95 70.2023
R863 B.n256 B.n95 70.2023
R864 B.n262 B.n91 70.2023
R865 B.n262 B.n87 70.2023
R866 B.n268 B.n87 70.2023
R867 B.n268 B.n83 70.2023
R868 B.n274 B.n83 70.2023
R869 B.n280 B.n79 70.2023
R870 B.n288 B.n75 70.2023
R871 B.n288 B.n287 70.2023
R872 B.n294 B.n4 70.2023
R873 B.n465 B.n4 70.2023
R874 B.n465 B.n464 70.2023
R875 B.n464 B.n463 70.2023
R876 B.n457 B.n11 70.2023
R877 B.n457 B.n456 70.2023
R878 B.n455 B.n15 70.2023
R879 B.n449 B.n448 70.2023
R880 B.n448 B.n447 70.2023
R881 B.n447 B.n22 70.2023
R882 B.n441 B.n22 70.2023
R883 B.n441 B.n440 70.2023
R884 B.n439 B.n29 70.2023
R885 B.n433 B.n29 70.2023
R886 B.n433 B.n432 70.2023
R887 B.n432 B.n431 70.2023
R888 B.t2 B.n79 59.8785
R889 B.n294 B.t3 59.8785
R890 B.n463 B.t5 59.8785
R891 B.t0 B.n15 59.8785
R892 B.n179 B.n125 59.5399
R893 B.n119 B.n118 59.5399
R894 B.n50 B.n49 59.5399
R895 B.n58 B.n57 59.5399
R896 B.n280 B.t1 45.4252
R897 B.t4 B.n455 45.4252
R898 B.t11 B.n91 39.2309
R899 B.n440 B.t7 39.2309
R900 B.n429 B.n428 32.9371
R901 B.n323 B.n320 32.9371
R902 B.n246 B.n101 32.9371
R903 B.n242 B.n241 32.9371
R904 B.n256 B.t11 30.9719
R905 B.t7 B.n439 30.9719
R906 B.t1 B.n75 24.7776
R907 B.n456 B.t4 24.7776
R908 B B.n467 18.0485
R909 B.n125 B.n124 16.4853
R910 B.n118 B.n117 16.4853
R911 B.n49 B.n48 16.4853
R912 B.n57 B.n56 16.4853
R913 B.n428 B.n427 10.6151
R914 B.n427 B.n38 10.6151
R915 B.n421 B.n38 10.6151
R916 B.n421 B.n420 10.6151
R917 B.n420 B.n419 10.6151
R918 B.n419 B.n40 10.6151
R919 B.n413 B.n40 10.6151
R920 B.n413 B.n412 10.6151
R921 B.n412 B.n411 10.6151
R922 B.n411 B.n42 10.6151
R923 B.n405 B.n42 10.6151
R924 B.n405 B.n404 10.6151
R925 B.n404 B.n403 10.6151
R926 B.n403 B.n44 10.6151
R927 B.n397 B.n44 10.6151
R928 B.n397 B.n396 10.6151
R929 B.n396 B.n395 10.6151
R930 B.n395 B.n46 10.6151
R931 B.n389 B.n46 10.6151
R932 B.n389 B.n388 10.6151
R933 B.n388 B.n387 10.6151
R934 B.n383 B.n382 10.6151
R935 B.n382 B.n52 10.6151
R936 B.n377 B.n52 10.6151
R937 B.n377 B.n376 10.6151
R938 B.n376 B.n375 10.6151
R939 B.n375 B.n54 10.6151
R940 B.n369 B.n54 10.6151
R941 B.n369 B.n368 10.6151
R942 B.n368 B.n367 10.6151
R943 B.n363 B.n362 10.6151
R944 B.n362 B.n60 10.6151
R945 B.n357 B.n60 10.6151
R946 B.n357 B.n356 10.6151
R947 B.n356 B.n355 10.6151
R948 B.n355 B.n62 10.6151
R949 B.n349 B.n62 10.6151
R950 B.n349 B.n348 10.6151
R951 B.n348 B.n347 10.6151
R952 B.n347 B.n64 10.6151
R953 B.n341 B.n64 10.6151
R954 B.n341 B.n340 10.6151
R955 B.n340 B.n339 10.6151
R956 B.n339 B.n66 10.6151
R957 B.n333 B.n66 10.6151
R958 B.n333 B.n332 10.6151
R959 B.n332 B.n331 10.6151
R960 B.n331 B.n68 10.6151
R961 B.n325 B.n68 10.6151
R962 B.n325 B.n324 10.6151
R963 B.n324 B.n323 10.6151
R964 B.n247 B.n246 10.6151
R965 B.n248 B.n247 10.6151
R966 B.n248 B.n93 10.6151
R967 B.n258 B.n93 10.6151
R968 B.n259 B.n258 10.6151
R969 B.n260 B.n259 10.6151
R970 B.n260 B.n85 10.6151
R971 B.n270 B.n85 10.6151
R972 B.n271 B.n270 10.6151
R973 B.n272 B.n271 10.6151
R974 B.n272 B.n77 10.6151
R975 B.n282 B.n77 10.6151
R976 B.n283 B.n282 10.6151
R977 B.n285 B.n283 10.6151
R978 B.n285 B.n284 10.6151
R979 B.n284 B.n70 10.6151
R980 B.n297 B.n70 10.6151
R981 B.n298 B.n297 10.6151
R982 B.n299 B.n298 10.6151
R983 B.n300 B.n299 10.6151
R984 B.n302 B.n300 10.6151
R985 B.n303 B.n302 10.6151
R986 B.n304 B.n303 10.6151
R987 B.n305 B.n304 10.6151
R988 B.n307 B.n305 10.6151
R989 B.n308 B.n307 10.6151
R990 B.n309 B.n308 10.6151
R991 B.n310 B.n309 10.6151
R992 B.n312 B.n310 10.6151
R993 B.n313 B.n312 10.6151
R994 B.n314 B.n313 10.6151
R995 B.n315 B.n314 10.6151
R996 B.n317 B.n315 10.6151
R997 B.n318 B.n317 10.6151
R998 B.n319 B.n318 10.6151
R999 B.n320 B.n319 10.6151
R1000 B.n241 B.n240 10.6151
R1001 B.n240 B.n105 10.6151
R1002 B.n235 B.n105 10.6151
R1003 B.n235 B.n234 10.6151
R1004 B.n234 B.n107 10.6151
R1005 B.n229 B.n107 10.6151
R1006 B.n229 B.n228 10.6151
R1007 B.n228 B.n227 10.6151
R1008 B.n227 B.n109 10.6151
R1009 B.n221 B.n109 10.6151
R1010 B.n221 B.n220 10.6151
R1011 B.n220 B.n219 10.6151
R1012 B.n219 B.n111 10.6151
R1013 B.n213 B.n111 10.6151
R1014 B.n213 B.n212 10.6151
R1015 B.n212 B.n211 10.6151
R1016 B.n211 B.n113 10.6151
R1017 B.n205 B.n113 10.6151
R1018 B.n205 B.n204 10.6151
R1019 B.n204 B.n203 10.6151
R1020 B.n203 B.n115 10.6151
R1021 B.n197 B.n196 10.6151
R1022 B.n196 B.n195 10.6151
R1023 B.n195 B.n120 10.6151
R1024 B.n189 B.n120 10.6151
R1025 B.n189 B.n188 10.6151
R1026 B.n188 B.n187 10.6151
R1027 B.n187 B.n122 10.6151
R1028 B.n181 B.n122 10.6151
R1029 B.n181 B.n180 10.6151
R1030 B.n178 B.n126 10.6151
R1031 B.n172 B.n126 10.6151
R1032 B.n172 B.n171 10.6151
R1033 B.n171 B.n170 10.6151
R1034 B.n170 B.n128 10.6151
R1035 B.n164 B.n128 10.6151
R1036 B.n164 B.n163 10.6151
R1037 B.n163 B.n162 10.6151
R1038 B.n162 B.n130 10.6151
R1039 B.n156 B.n130 10.6151
R1040 B.n156 B.n155 10.6151
R1041 B.n155 B.n154 10.6151
R1042 B.n154 B.n132 10.6151
R1043 B.n148 B.n132 10.6151
R1044 B.n148 B.n147 10.6151
R1045 B.n147 B.n146 10.6151
R1046 B.n146 B.n134 10.6151
R1047 B.n140 B.n134 10.6151
R1048 B.n140 B.n139 10.6151
R1049 B.n139 B.n138 10.6151
R1050 B.n138 B.n101 10.6151
R1051 B.n242 B.n97 10.6151
R1052 B.n252 B.n97 10.6151
R1053 B.n253 B.n252 10.6151
R1054 B.n254 B.n253 10.6151
R1055 B.n254 B.n89 10.6151
R1056 B.n264 B.n89 10.6151
R1057 B.n265 B.n264 10.6151
R1058 B.n266 B.n265 10.6151
R1059 B.n266 B.n81 10.6151
R1060 B.n276 B.n81 10.6151
R1061 B.n277 B.n276 10.6151
R1062 B.n278 B.n277 10.6151
R1063 B.n278 B.n73 10.6151
R1064 B.n290 B.n73 10.6151
R1065 B.n291 B.n290 10.6151
R1066 B.n292 B.n291 10.6151
R1067 B.n292 B.n0 10.6151
R1068 B.n461 B.n1 10.6151
R1069 B.n461 B.n460 10.6151
R1070 B.n460 B.n459 10.6151
R1071 B.n459 B.n9 10.6151
R1072 B.n453 B.n9 10.6151
R1073 B.n453 B.n452 10.6151
R1074 B.n452 B.n451 10.6151
R1075 B.n451 B.n17 10.6151
R1076 B.n445 B.n17 10.6151
R1077 B.n445 B.n444 10.6151
R1078 B.n444 B.n443 10.6151
R1079 B.n443 B.n24 10.6151
R1080 B.n437 B.n24 10.6151
R1081 B.n437 B.n436 10.6151
R1082 B.n436 B.n435 10.6151
R1083 B.n435 B.n31 10.6151
R1084 B.n429 B.n31 10.6151
R1085 B.n274 B.t2 10.3243
R1086 B.n287 B.t3 10.3243
R1087 B.n11 B.t5 10.3243
R1088 B.n449 B.t0 10.3243
R1089 B.n387 B.n50 9.36635
R1090 B.n363 B.n58 9.36635
R1091 B.n119 B.n115 9.36635
R1092 B.n179 B.n178 9.36635
R1093 B.n467 B.n0 2.81026
R1094 B.n467 B.n1 2.81026
R1095 B.n383 B.n50 1.24928
R1096 B.n367 B.n58 1.24928
R1097 B.n197 B.n119 1.24928
R1098 B.n180 B.n179 1.24928
R1099 VN.n0 VN.t0 351.709
R1100 VN.n4 VN.t1 351.709
R1101 VN.n1 VN.t2 324.887
R1102 VN.n2 VN.t5 324.887
R1103 VN.n5 VN.t4 324.887
R1104 VN.n6 VN.t3 324.887
R1105 VN.n3 VN.n2 161.3
R1106 VN.n7 VN.n6 161.3
R1107 VN.n2 VN.n1 48.2005
R1108 VN.n6 VN.n5 48.2005
R1109 VN.n7 VN.n4 45.1367
R1110 VN.n3 VN.n0 45.1367
R1111 VN VN.n7 35.8698
R1112 VN.n5 VN.n4 13.3799
R1113 VN.n1 VN.n0 13.3799
R1114 VN VN.n3 0.0516364
R1115 VDD2.n51 VDD2.n29 289.615
R1116 VDD2.n22 VDD2.n0 289.615
R1117 VDD2.n52 VDD2.n51 185
R1118 VDD2.n50 VDD2.n49 185
R1119 VDD2.n33 VDD2.n32 185
R1120 VDD2.n44 VDD2.n43 185
R1121 VDD2.n42 VDD2.n41 185
R1122 VDD2.n37 VDD2.n36 185
R1123 VDD2.n8 VDD2.n7 185
R1124 VDD2.n13 VDD2.n12 185
R1125 VDD2.n15 VDD2.n14 185
R1126 VDD2.n4 VDD2.n3 185
R1127 VDD2.n21 VDD2.n20 185
R1128 VDD2.n23 VDD2.n22 185
R1129 VDD2.n38 VDD2.t2 147.672
R1130 VDD2.n9 VDD2.t5 147.672
R1131 VDD2.n51 VDD2.n50 104.615
R1132 VDD2.n50 VDD2.n32 104.615
R1133 VDD2.n43 VDD2.n32 104.615
R1134 VDD2.n43 VDD2.n42 104.615
R1135 VDD2.n42 VDD2.n36 104.615
R1136 VDD2.n13 VDD2.n7 104.615
R1137 VDD2.n14 VDD2.n13 104.615
R1138 VDD2.n14 VDD2.n3 104.615
R1139 VDD2.n21 VDD2.n3 104.615
R1140 VDD2.n22 VDD2.n21 104.615
R1141 VDD2.n28 VDD2.n27 70.7223
R1142 VDD2 VDD2.n57 70.7195
R1143 VDD2.t2 VDD2.n36 52.3082
R1144 VDD2.t5 VDD2.n7 52.3082
R1145 VDD2.n28 VDD2.n26 51.2978
R1146 VDD2.n56 VDD2.n55 50.8035
R1147 VDD2.n56 VDD2.n28 30.7347
R1148 VDD2.n38 VDD2.n37 15.6666
R1149 VDD2.n9 VDD2.n8 15.6666
R1150 VDD2.n41 VDD2.n40 12.8005
R1151 VDD2.n12 VDD2.n11 12.8005
R1152 VDD2.n44 VDD2.n35 12.0247
R1153 VDD2.n15 VDD2.n6 12.0247
R1154 VDD2.n45 VDD2.n33 11.249
R1155 VDD2.n16 VDD2.n4 11.249
R1156 VDD2.n49 VDD2.n48 10.4732
R1157 VDD2.n20 VDD2.n19 10.4732
R1158 VDD2.n52 VDD2.n31 9.69747
R1159 VDD2.n23 VDD2.n2 9.69747
R1160 VDD2.n55 VDD2.n54 9.45567
R1161 VDD2.n26 VDD2.n25 9.45567
R1162 VDD2.n54 VDD2.n53 9.3005
R1163 VDD2.n31 VDD2.n30 9.3005
R1164 VDD2.n48 VDD2.n47 9.3005
R1165 VDD2.n46 VDD2.n45 9.3005
R1166 VDD2.n35 VDD2.n34 9.3005
R1167 VDD2.n40 VDD2.n39 9.3005
R1168 VDD2.n25 VDD2.n24 9.3005
R1169 VDD2.n2 VDD2.n1 9.3005
R1170 VDD2.n19 VDD2.n18 9.3005
R1171 VDD2.n17 VDD2.n16 9.3005
R1172 VDD2.n6 VDD2.n5 9.3005
R1173 VDD2.n11 VDD2.n10 9.3005
R1174 VDD2.n53 VDD2.n29 8.92171
R1175 VDD2.n24 VDD2.n0 8.92171
R1176 VDD2.n55 VDD2.n29 5.04292
R1177 VDD2.n26 VDD2.n0 5.04292
R1178 VDD2.n39 VDD2.n38 4.38687
R1179 VDD2.n10 VDD2.n9 4.38687
R1180 VDD2.n53 VDD2.n52 4.26717
R1181 VDD2.n24 VDD2.n23 4.26717
R1182 VDD2.n57 VDD2.t1 3.6808
R1183 VDD2.n57 VDD2.t4 3.6808
R1184 VDD2.n27 VDD2.t3 3.6808
R1185 VDD2.n27 VDD2.t0 3.6808
R1186 VDD2.n49 VDD2.n31 3.49141
R1187 VDD2.n20 VDD2.n2 3.49141
R1188 VDD2.n48 VDD2.n33 2.71565
R1189 VDD2.n19 VDD2.n4 2.71565
R1190 VDD2.n45 VDD2.n44 1.93989
R1191 VDD2.n16 VDD2.n15 1.93989
R1192 VDD2.n41 VDD2.n35 1.16414
R1193 VDD2.n12 VDD2.n6 1.16414
R1194 VDD2 VDD2.n56 0.608259
R1195 VDD2.n40 VDD2.n37 0.388379
R1196 VDD2.n11 VDD2.n8 0.388379
R1197 VDD2.n54 VDD2.n30 0.155672
R1198 VDD2.n47 VDD2.n30 0.155672
R1199 VDD2.n47 VDD2.n46 0.155672
R1200 VDD2.n46 VDD2.n34 0.155672
R1201 VDD2.n39 VDD2.n34 0.155672
R1202 VDD2.n10 VDD2.n5 0.155672
R1203 VDD2.n17 VDD2.n5 0.155672
R1204 VDD2.n18 VDD2.n17 0.155672
R1205 VDD2.n18 VDD2.n1 0.155672
R1206 VDD2.n25 VDD2.n1 0.155672
C0 VN VP 3.67912f
C1 VDD1 VDD2 0.644993f
C2 VDD1 VTAIL 5.95927f
C3 VDD1 VP 1.97543f
C4 VDD1 VN 0.148283f
C5 VTAIL VDD2 5.99546f
C6 VDD2 VP 0.285634f
C7 VTAIL VP 1.80702f
C8 VN VDD2 1.84428f
C9 VN VTAIL 1.79267f
C10 VDD2 B 3.07981f
C11 VDD1 B 3.124812f
C12 VTAIL B 3.695732f
C13 VN B 5.611774f
C14 VP B 4.693738f
C15 VDD2.n0 B 0.027074f
C16 VDD2.n1 B 0.018723f
C17 VDD2.n2 B 0.010061f
C18 VDD2.n3 B 0.02378f
C19 VDD2.n4 B 0.010653f
C20 VDD2.n5 B 0.018723f
C21 VDD2.n6 B 0.010061f
C22 VDD2.n7 B 0.017835f
C23 VDD2.n8 B 0.014044f
C24 VDD2.t5 B 0.038875f
C25 VDD2.n9 B 0.077515f
C26 VDD2.n10 B 0.391826f
C27 VDD2.n11 B 0.010061f
C28 VDD2.n12 B 0.010653f
C29 VDD2.n13 B 0.02378f
C30 VDD2.n14 B 0.02378f
C31 VDD2.n15 B 0.010653f
C32 VDD2.n16 B 0.010061f
C33 VDD2.n17 B 0.018723f
C34 VDD2.n18 B 0.018723f
C35 VDD2.n19 B 0.010061f
C36 VDD2.n20 B 0.010653f
C37 VDD2.n21 B 0.02378f
C38 VDD2.n22 B 0.05282f
C39 VDD2.n23 B 0.010653f
C40 VDD2.n24 B 0.010061f
C41 VDD2.n25 B 0.045834f
C42 VDD2.n26 B 0.043335f
C43 VDD2.t3 B 0.079598f
C44 VDD2.t0 B 0.079598f
C45 VDD2.n27 B 0.655307f
C46 VDD2.n28 B 1.03305f
C47 VDD2.n29 B 0.027074f
C48 VDD2.n30 B 0.018723f
C49 VDD2.n31 B 0.010061f
C50 VDD2.n32 B 0.02378f
C51 VDD2.n33 B 0.010653f
C52 VDD2.n34 B 0.018723f
C53 VDD2.n35 B 0.010061f
C54 VDD2.n36 B 0.017835f
C55 VDD2.n37 B 0.014044f
C56 VDD2.t2 B 0.038875f
C57 VDD2.n38 B 0.077515f
C58 VDD2.n39 B 0.391826f
C59 VDD2.n40 B 0.010061f
C60 VDD2.n41 B 0.010653f
C61 VDD2.n42 B 0.02378f
C62 VDD2.n43 B 0.02378f
C63 VDD2.n44 B 0.010653f
C64 VDD2.n45 B 0.010061f
C65 VDD2.n46 B 0.018723f
C66 VDD2.n47 B 0.018723f
C67 VDD2.n48 B 0.010061f
C68 VDD2.n49 B 0.010653f
C69 VDD2.n50 B 0.02378f
C70 VDD2.n51 B 0.05282f
C71 VDD2.n52 B 0.010653f
C72 VDD2.n53 B 0.010061f
C73 VDD2.n54 B 0.045834f
C74 VDD2.n55 B 0.042678f
C75 VDD2.n56 B 1.0998f
C76 VDD2.t1 B 0.079598f
C77 VDD2.t4 B 0.079598f
C78 VDD2.n57 B 0.655292f
C79 VN.t0 B 0.218674f
C80 VN.n0 B 0.095033f
C81 VN.t2 B 0.210866f
C82 VN.n1 B 0.10819f
C83 VN.t5 B 0.210866f
C84 VN.n2 B 0.102317f
C85 VN.n3 B 0.100703f
C86 VN.t1 B 0.218674f
C87 VN.n4 B 0.095033f
C88 VN.t4 B 0.210866f
C89 VN.n5 B 0.10819f
C90 VN.t3 B 0.210866f
C91 VN.n6 B 0.102317f
C92 VN.n7 B 0.889901f
C93 VDD1.n0 B 0.026766f
C94 VDD1.n1 B 0.018509f
C95 VDD1.n2 B 0.009946f
C96 VDD1.n3 B 0.023509f
C97 VDD1.n4 B 0.010531f
C98 VDD1.n5 B 0.018509f
C99 VDD1.n6 B 0.009946f
C100 VDD1.n7 B 0.017632f
C101 VDD1.n8 B 0.013884f
C102 VDD1.t0 B 0.038432f
C103 VDD1.n9 B 0.076632f
C104 VDD1.n10 B 0.387362f
C105 VDD1.n11 B 0.009946f
C106 VDD1.n12 B 0.010531f
C107 VDD1.n13 B 0.023509f
C108 VDD1.n14 B 0.023509f
C109 VDD1.n15 B 0.010531f
C110 VDD1.n16 B 0.009946f
C111 VDD1.n17 B 0.018509f
C112 VDD1.n18 B 0.018509f
C113 VDD1.n19 B 0.009946f
C114 VDD1.n20 B 0.010531f
C115 VDD1.n21 B 0.023509f
C116 VDD1.n22 B 0.052218f
C117 VDD1.n23 B 0.010531f
C118 VDD1.n24 B 0.009946f
C119 VDD1.n25 B 0.045312f
C120 VDD1.n26 B 0.043058f
C121 VDD1.n27 B 0.026766f
C122 VDD1.n28 B 0.018509f
C123 VDD1.n29 B 0.009946f
C124 VDD1.n30 B 0.023509f
C125 VDD1.n31 B 0.010531f
C126 VDD1.n32 B 0.018509f
C127 VDD1.n33 B 0.009946f
C128 VDD1.n34 B 0.017632f
C129 VDD1.n35 B 0.013884f
C130 VDD1.t1 B 0.038432f
C131 VDD1.n36 B 0.076632f
C132 VDD1.n37 B 0.387362f
C133 VDD1.n38 B 0.009946f
C134 VDD1.n39 B 0.010531f
C135 VDD1.n40 B 0.023509f
C136 VDD1.n41 B 0.023509f
C137 VDD1.n42 B 0.010531f
C138 VDD1.n43 B 0.009946f
C139 VDD1.n44 B 0.018509f
C140 VDD1.n45 B 0.018509f
C141 VDD1.n46 B 0.009946f
C142 VDD1.n47 B 0.010531f
C143 VDD1.n48 B 0.023509f
C144 VDD1.n49 B 0.052218f
C145 VDD1.n50 B 0.010531f
C146 VDD1.n51 B 0.009946f
C147 VDD1.n52 B 0.045312f
C148 VDD1.n53 B 0.042841f
C149 VDD1.t2 B 0.078691f
C150 VDD1.t4 B 0.078691f
C151 VDD1.n54 B 0.64784f
C152 VDD1.n55 B 1.07352f
C153 VDD1.t3 B 0.078691f
C154 VDD1.t5 B 0.078691f
C155 VDD1.n56 B 0.64746f
C156 VDD1.n57 B 1.23706f
C157 VTAIL.t11 B 0.089278f
C158 VTAIL.t4 B 0.089278f
C159 VTAIL.n0 B 0.683719f
C160 VTAIL.n1 B 0.263578f
C161 VTAIL.n2 B 0.030367f
C162 VTAIL.n3 B 0.020999f
C163 VTAIL.n4 B 0.011284f
C164 VTAIL.n5 B 0.026672f
C165 VTAIL.n6 B 0.011948f
C166 VTAIL.n7 B 0.020999f
C167 VTAIL.n8 B 0.011284f
C168 VTAIL.n9 B 0.020004f
C169 VTAIL.n10 B 0.015752f
C170 VTAIL.t6 B 0.043603f
C171 VTAIL.n11 B 0.086942f
C172 VTAIL.n12 B 0.439475f
C173 VTAIL.n13 B 0.011284f
C174 VTAIL.n14 B 0.011948f
C175 VTAIL.n15 B 0.026672f
C176 VTAIL.n16 B 0.026672f
C177 VTAIL.n17 B 0.011948f
C178 VTAIL.n18 B 0.011284f
C179 VTAIL.n19 B 0.020999f
C180 VTAIL.n20 B 0.020999f
C181 VTAIL.n21 B 0.011284f
C182 VTAIL.n22 B 0.011948f
C183 VTAIL.n23 B 0.026672f
C184 VTAIL.n24 B 0.059243f
C185 VTAIL.n25 B 0.011948f
C186 VTAIL.n26 B 0.011284f
C187 VTAIL.n27 B 0.051408f
C188 VTAIL.n28 B 0.033389f
C189 VTAIL.n29 B 0.12572f
C190 VTAIL.t10 B 0.089278f
C191 VTAIL.t8 B 0.089278f
C192 VTAIL.n30 B 0.683719f
C193 VTAIL.n31 B 0.938486f
C194 VTAIL.t2 B 0.089278f
C195 VTAIL.t1 B 0.089278f
C196 VTAIL.n32 B 0.683724f
C197 VTAIL.n33 B 0.938481f
C198 VTAIL.n34 B 0.030367f
C199 VTAIL.n35 B 0.020999f
C200 VTAIL.n36 B 0.011284f
C201 VTAIL.n37 B 0.026672f
C202 VTAIL.n38 B 0.011948f
C203 VTAIL.n39 B 0.020999f
C204 VTAIL.n40 B 0.011284f
C205 VTAIL.n41 B 0.020004f
C206 VTAIL.n42 B 0.015752f
C207 VTAIL.t3 B 0.043603f
C208 VTAIL.n43 B 0.086942f
C209 VTAIL.n44 B 0.439475f
C210 VTAIL.n45 B 0.011284f
C211 VTAIL.n46 B 0.011948f
C212 VTAIL.n47 B 0.026672f
C213 VTAIL.n48 B 0.026672f
C214 VTAIL.n49 B 0.011948f
C215 VTAIL.n50 B 0.011284f
C216 VTAIL.n51 B 0.020999f
C217 VTAIL.n52 B 0.020999f
C218 VTAIL.n53 B 0.011284f
C219 VTAIL.n54 B 0.011948f
C220 VTAIL.n55 B 0.026672f
C221 VTAIL.n56 B 0.059243f
C222 VTAIL.n57 B 0.011948f
C223 VTAIL.n58 B 0.011284f
C224 VTAIL.n59 B 0.051408f
C225 VTAIL.n60 B 0.033389f
C226 VTAIL.n61 B 0.12572f
C227 VTAIL.t5 B 0.089278f
C228 VTAIL.t7 B 0.089278f
C229 VTAIL.n62 B 0.683724f
C230 VTAIL.n63 B 0.296822f
C231 VTAIL.n64 B 0.030367f
C232 VTAIL.n65 B 0.020999f
C233 VTAIL.n66 B 0.011284f
C234 VTAIL.n67 B 0.026672f
C235 VTAIL.n68 B 0.011948f
C236 VTAIL.n69 B 0.020999f
C237 VTAIL.n70 B 0.011284f
C238 VTAIL.n71 B 0.020004f
C239 VTAIL.n72 B 0.015752f
C240 VTAIL.t9 B 0.043603f
C241 VTAIL.n73 B 0.086942f
C242 VTAIL.n74 B 0.439475f
C243 VTAIL.n75 B 0.011284f
C244 VTAIL.n76 B 0.011948f
C245 VTAIL.n77 B 0.026672f
C246 VTAIL.n78 B 0.026672f
C247 VTAIL.n79 B 0.011948f
C248 VTAIL.n80 B 0.011284f
C249 VTAIL.n81 B 0.020999f
C250 VTAIL.n82 B 0.020999f
C251 VTAIL.n83 B 0.011284f
C252 VTAIL.n84 B 0.011948f
C253 VTAIL.n85 B 0.026672f
C254 VTAIL.n86 B 0.059243f
C255 VTAIL.n87 B 0.011948f
C256 VTAIL.n88 B 0.011284f
C257 VTAIL.n89 B 0.051408f
C258 VTAIL.n90 B 0.033389f
C259 VTAIL.n91 B 0.717797f
C260 VTAIL.n92 B 0.030367f
C261 VTAIL.n93 B 0.020999f
C262 VTAIL.n94 B 0.011284f
C263 VTAIL.n95 B 0.026672f
C264 VTAIL.n96 B 0.011948f
C265 VTAIL.n97 B 0.020999f
C266 VTAIL.n98 B 0.011284f
C267 VTAIL.n99 B 0.020004f
C268 VTAIL.n100 B 0.015752f
C269 VTAIL.t0 B 0.043603f
C270 VTAIL.n101 B 0.086942f
C271 VTAIL.n102 B 0.439475f
C272 VTAIL.n103 B 0.011284f
C273 VTAIL.n104 B 0.011948f
C274 VTAIL.n105 B 0.026672f
C275 VTAIL.n106 B 0.026672f
C276 VTAIL.n107 B 0.011948f
C277 VTAIL.n108 B 0.011284f
C278 VTAIL.n109 B 0.020999f
C279 VTAIL.n110 B 0.020999f
C280 VTAIL.n111 B 0.011284f
C281 VTAIL.n112 B 0.011948f
C282 VTAIL.n113 B 0.026672f
C283 VTAIL.n114 B 0.059243f
C284 VTAIL.n115 B 0.011948f
C285 VTAIL.n116 B 0.011284f
C286 VTAIL.n117 B 0.051408f
C287 VTAIL.n118 B 0.033389f
C288 VTAIL.n119 B 0.701464f
C289 VP.n0 B 0.034802f
C290 VP.t5 B 0.220846f
C291 VP.n1 B 0.095976f
C292 VP.t0 B 0.212961f
C293 VP.t2 B 0.212961f
C294 VP.n2 B 0.109265f
C295 VP.n3 B 0.103333f
C296 VP.n4 B 0.881381f
C297 VP.n5 B 0.835234f
C298 VP.t4 B 0.212961f
C299 VP.n6 B 0.103333f
C300 VP.t3 B 0.212961f
C301 VP.n7 B 0.109265f
C302 VP.t1 B 0.212961f
C303 VP.n8 B 0.103333f
C304 VP.n9 B 0.029001f
.ends

