* NGSPICE file created from diff_pair_sample_0859.ext - technology: sky130A

.subckt diff_pair_sample_0859 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t14 VP.t0 VDD1.t6 B.t2 sky130_fd_pr__nfet_01v8 ad=0.94545 pd=6.06 as=0.94545 ps=6.06 w=5.73 l=0.37
X1 B.t20 B.t18 B.t19 B.t12 sky130_fd_pr__nfet_01v8 ad=2.2347 pd=12.24 as=0 ps=0 w=5.73 l=0.37
X2 B.t17 B.t15 B.t16 B.t8 sky130_fd_pr__nfet_01v8 ad=2.2347 pd=12.24 as=0 ps=0 w=5.73 l=0.37
X3 VDD2.t7 VN.t0 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=0.94545 pd=6.06 as=0.94545 ps=6.06 w=5.73 l=0.37
X4 VTAIL.t4 VN.t1 VDD2.t6 B.t4 sky130_fd_pr__nfet_01v8 ad=0.94545 pd=6.06 as=0.94545 ps=6.06 w=5.73 l=0.37
X5 VTAIL.t2 VN.t2 VDD2.t5 B.t2 sky130_fd_pr__nfet_01v8 ad=0.94545 pd=6.06 as=0.94545 ps=6.06 w=5.73 l=0.37
X6 VDD2.t4 VN.t3 VTAIL.t6 B.t6 sky130_fd_pr__nfet_01v8 ad=0.94545 pd=6.06 as=0.94545 ps=6.06 w=5.73 l=0.37
X7 VDD1.t0 VP.t1 VTAIL.t13 B.t6 sky130_fd_pr__nfet_01v8 ad=0.94545 pd=6.06 as=0.94545 ps=6.06 w=5.73 l=0.37
X8 B.t14 B.t11 B.t13 B.t12 sky130_fd_pr__nfet_01v8 ad=2.2347 pd=12.24 as=0 ps=0 w=5.73 l=0.37
X9 VTAIL.t3 VN.t4 VDD2.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=2.2347 pd=12.24 as=0.94545 ps=6.06 w=5.73 l=0.37
X10 B.t10 B.t7 B.t9 B.t8 sky130_fd_pr__nfet_01v8 ad=2.2347 pd=12.24 as=0 ps=0 w=5.73 l=0.37
X11 VDD2.t2 VN.t5 VTAIL.t15 B.t21 sky130_fd_pr__nfet_01v8 ad=0.94545 pd=6.06 as=2.2347 ps=12.24 w=5.73 l=0.37
X12 VDD2.t1 VN.t6 VTAIL.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=0.94545 pd=6.06 as=2.2347 ps=12.24 w=5.73 l=0.37
X13 VTAIL.t12 VP.t2 VDD1.t7 B.t4 sky130_fd_pr__nfet_01v8 ad=0.94545 pd=6.06 as=0.94545 ps=6.06 w=5.73 l=0.37
X14 VTAIL.t11 VP.t3 VDD1.t1 B.t3 sky130_fd_pr__nfet_01v8 ad=2.2347 pd=12.24 as=0.94545 ps=6.06 w=5.73 l=0.37
X15 VDD1.t4 VP.t4 VTAIL.t10 B.t5 sky130_fd_pr__nfet_01v8 ad=0.94545 pd=6.06 as=2.2347 ps=12.24 w=5.73 l=0.37
X16 VTAIL.t9 VP.t5 VDD1.t5 B.t0 sky130_fd_pr__nfet_01v8 ad=2.2347 pd=12.24 as=0.94545 ps=6.06 w=5.73 l=0.37
X17 VTAIL.t0 VN.t7 VDD2.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=2.2347 pd=12.24 as=0.94545 ps=6.06 w=5.73 l=0.37
X18 VDD1.t3 VP.t6 VTAIL.t8 B.t1 sky130_fd_pr__nfet_01v8 ad=0.94545 pd=6.06 as=0.94545 ps=6.06 w=5.73 l=0.37
X19 VDD1.t2 VP.t7 VTAIL.t7 B.t21 sky130_fd_pr__nfet_01v8 ad=0.94545 pd=6.06 as=2.2347 ps=12.24 w=5.73 l=0.37
R0 VP.n3 VP.t3 511.161
R1 VP.n12 VP.t4 496.844
R2 VP.n1 VP.t5 496.844
R3 VP.n6 VP.t7 496.844
R4 VP.n10 VP.t6 480.046
R5 VP.n11 VP.t2 480.046
R6 VP.n5 VP.t0 480.046
R7 VP.n4 VP.t1 480.046
R8 VP.n13 VP.n12 161.3
R9 VP.n5 VP.n2 161.3
R10 VP.n7 VP.n6 161.3
R11 VP.n11 VP.n0 161.3
R12 VP.n10 VP.n9 161.3
R13 VP.n8 VP.n1 161.3
R14 VP.n3 VP.n2 73.733
R15 VP.n11 VP.n10 48.2005
R16 VP.n5 VP.n4 48.2005
R17 VP.n8 VP.n7 35.8111
R18 VP.n10 VP.n1 31.4035
R19 VP.n12 VP.n11 31.4035
R20 VP.n6 VP.n5 31.4035
R21 VP.n4 VP.n3 14.302
R22 VP.n7 VP.n2 0.189894
R23 VP.n9 VP.n8 0.189894
R24 VP.n9 VP.n0 0.189894
R25 VP.n13 VP.n0 0.189894
R26 VP VP.n13 0.0516364
R27 VDD1 VDD1.n0 69.9754
R28 VDD1.n3 VDD1.n2 69.8616
R29 VDD1.n3 VDD1.n1 69.8616
R30 VDD1.n5 VDD1.n4 69.6153
R31 VDD1.n5 VDD1.n3 31.9535
R32 VDD1.n4 VDD1.t6 3.456
R33 VDD1.n4 VDD1.t2 3.456
R34 VDD1.n0 VDD1.t1 3.456
R35 VDD1.n0 VDD1.t0 3.456
R36 VDD1.n2 VDD1.t7 3.456
R37 VDD1.n2 VDD1.t4 3.456
R38 VDD1.n1 VDD1.t5 3.456
R39 VDD1.n1 VDD1.t3 3.456
R40 VDD1 VDD1.n5 0.244034
R41 VTAIL.n11 VTAIL.t11 56.3922
R42 VTAIL.n10 VTAIL.t5 56.3922
R43 VTAIL.n7 VTAIL.t0 56.3922
R44 VTAIL.n15 VTAIL.t15 56.392
R45 VTAIL.n2 VTAIL.t3 56.392
R46 VTAIL.n3 VTAIL.t10 56.392
R47 VTAIL.n6 VTAIL.t9 56.392
R48 VTAIL.n14 VTAIL.t7 56.392
R49 VTAIL.n13 VTAIL.n12 52.9367
R50 VTAIL.n9 VTAIL.n8 52.9367
R51 VTAIL.n1 VTAIL.n0 52.9365
R52 VTAIL.n5 VTAIL.n4 52.9365
R53 VTAIL.n15 VTAIL.n14 17.91
R54 VTAIL.n7 VTAIL.n6 17.91
R55 VTAIL.n0 VTAIL.t6 3.456
R56 VTAIL.n0 VTAIL.t2 3.456
R57 VTAIL.n4 VTAIL.t8 3.456
R58 VTAIL.n4 VTAIL.t12 3.456
R59 VTAIL.n12 VTAIL.t13 3.456
R60 VTAIL.n12 VTAIL.t14 3.456
R61 VTAIL.n8 VTAIL.t1 3.456
R62 VTAIL.n8 VTAIL.t4 3.456
R63 VTAIL.n9 VTAIL.n7 0.603948
R64 VTAIL.n10 VTAIL.n9 0.603948
R65 VTAIL.n13 VTAIL.n11 0.603948
R66 VTAIL.n14 VTAIL.n13 0.603948
R67 VTAIL.n6 VTAIL.n5 0.603948
R68 VTAIL.n5 VTAIL.n3 0.603948
R69 VTAIL.n2 VTAIL.n1 0.603948
R70 VTAIL VTAIL.n15 0.545759
R71 VTAIL.n11 VTAIL.n10 0.470328
R72 VTAIL.n3 VTAIL.n2 0.470328
R73 VTAIL VTAIL.n1 0.0586897
R74 B.n330 B.n329 585
R75 B.n332 B.n70 585
R76 B.n335 B.n334 585
R77 B.n336 B.n69 585
R78 B.n338 B.n337 585
R79 B.n340 B.n68 585
R80 B.n343 B.n342 585
R81 B.n344 B.n67 585
R82 B.n346 B.n345 585
R83 B.n348 B.n66 585
R84 B.n351 B.n350 585
R85 B.n352 B.n65 585
R86 B.n354 B.n353 585
R87 B.n356 B.n64 585
R88 B.n359 B.n358 585
R89 B.n360 B.n63 585
R90 B.n362 B.n361 585
R91 B.n364 B.n62 585
R92 B.n367 B.n366 585
R93 B.n368 B.n61 585
R94 B.n370 B.n369 585
R95 B.n372 B.n60 585
R96 B.n375 B.n374 585
R97 B.n377 B.n57 585
R98 B.n379 B.n378 585
R99 B.n381 B.n56 585
R100 B.n384 B.n383 585
R101 B.n385 B.n55 585
R102 B.n387 B.n386 585
R103 B.n389 B.n54 585
R104 B.n392 B.n391 585
R105 B.n393 B.n50 585
R106 B.n395 B.n394 585
R107 B.n397 B.n49 585
R108 B.n400 B.n399 585
R109 B.n401 B.n48 585
R110 B.n403 B.n402 585
R111 B.n405 B.n47 585
R112 B.n408 B.n407 585
R113 B.n409 B.n46 585
R114 B.n411 B.n410 585
R115 B.n413 B.n45 585
R116 B.n416 B.n415 585
R117 B.n417 B.n44 585
R118 B.n419 B.n418 585
R119 B.n421 B.n43 585
R120 B.n424 B.n423 585
R121 B.n425 B.n42 585
R122 B.n427 B.n426 585
R123 B.n429 B.n41 585
R124 B.n432 B.n431 585
R125 B.n433 B.n40 585
R126 B.n435 B.n434 585
R127 B.n437 B.n39 585
R128 B.n440 B.n439 585
R129 B.n441 B.n38 585
R130 B.n328 B.n36 585
R131 B.n444 B.n36 585
R132 B.n327 B.n35 585
R133 B.n445 B.n35 585
R134 B.n326 B.n34 585
R135 B.n446 B.n34 585
R136 B.n325 B.n324 585
R137 B.n324 B.n30 585
R138 B.n323 B.n29 585
R139 B.n452 B.n29 585
R140 B.n322 B.n28 585
R141 B.n453 B.n28 585
R142 B.n321 B.n27 585
R143 B.n454 B.n27 585
R144 B.n320 B.n319 585
R145 B.n319 B.n23 585
R146 B.n318 B.n22 585
R147 B.n460 B.n22 585
R148 B.n317 B.n21 585
R149 B.n461 B.n21 585
R150 B.n316 B.n20 585
R151 B.n462 B.n20 585
R152 B.n315 B.n314 585
R153 B.n314 B.n19 585
R154 B.n313 B.n15 585
R155 B.n468 B.n15 585
R156 B.n312 B.n14 585
R157 B.n469 B.n14 585
R158 B.n311 B.n13 585
R159 B.n470 B.n13 585
R160 B.n310 B.n309 585
R161 B.n309 B.n12 585
R162 B.n308 B.n307 585
R163 B.n308 B.n8 585
R164 B.n306 B.n7 585
R165 B.n477 B.n7 585
R166 B.n305 B.n6 585
R167 B.n478 B.n6 585
R168 B.n304 B.n5 585
R169 B.n479 B.n5 585
R170 B.n303 B.n302 585
R171 B.n302 B.n4 585
R172 B.n301 B.n71 585
R173 B.n301 B.n300 585
R174 B.n290 B.n72 585
R175 B.n293 B.n72 585
R176 B.n292 B.n291 585
R177 B.n294 B.n292 585
R178 B.n289 B.n76 585
R179 B.n79 B.n76 585
R180 B.n288 B.n287 585
R181 B.n287 B.n286 585
R182 B.n78 B.n77 585
R183 B.n279 B.n78 585
R184 B.n278 B.n277 585
R185 B.n280 B.n278 585
R186 B.n276 B.n83 585
R187 B.n87 B.n83 585
R188 B.n275 B.n274 585
R189 B.n274 B.n273 585
R190 B.n85 B.n84 585
R191 B.n86 B.n85 585
R192 B.n266 B.n265 585
R193 B.n267 B.n266 585
R194 B.n264 B.n92 585
R195 B.n92 B.n91 585
R196 B.n263 B.n262 585
R197 B.n262 B.n261 585
R198 B.n94 B.n93 585
R199 B.n95 B.n94 585
R200 B.n254 B.n253 585
R201 B.n255 B.n254 585
R202 B.n252 B.n100 585
R203 B.n100 B.n99 585
R204 B.n251 B.n250 585
R205 B.n250 B.n249 585
R206 B.n246 B.n104 585
R207 B.n245 B.n244 585
R208 B.n242 B.n105 585
R209 B.n242 B.n103 585
R210 B.n241 B.n240 585
R211 B.n239 B.n238 585
R212 B.n237 B.n107 585
R213 B.n235 B.n234 585
R214 B.n233 B.n108 585
R215 B.n232 B.n231 585
R216 B.n229 B.n109 585
R217 B.n227 B.n226 585
R218 B.n225 B.n110 585
R219 B.n224 B.n223 585
R220 B.n221 B.n111 585
R221 B.n219 B.n218 585
R222 B.n217 B.n112 585
R223 B.n216 B.n215 585
R224 B.n213 B.n113 585
R225 B.n211 B.n210 585
R226 B.n209 B.n114 585
R227 B.n208 B.n207 585
R228 B.n205 B.n115 585
R229 B.n203 B.n202 585
R230 B.n200 B.n116 585
R231 B.n199 B.n198 585
R232 B.n196 B.n119 585
R233 B.n194 B.n193 585
R234 B.n192 B.n120 585
R235 B.n191 B.n190 585
R236 B.n188 B.n121 585
R237 B.n186 B.n185 585
R238 B.n184 B.n122 585
R239 B.n183 B.n182 585
R240 B.n180 B.n179 585
R241 B.n178 B.n177 585
R242 B.n176 B.n127 585
R243 B.n174 B.n173 585
R244 B.n172 B.n128 585
R245 B.n171 B.n170 585
R246 B.n168 B.n129 585
R247 B.n166 B.n165 585
R248 B.n164 B.n130 585
R249 B.n163 B.n162 585
R250 B.n160 B.n131 585
R251 B.n158 B.n157 585
R252 B.n156 B.n132 585
R253 B.n155 B.n154 585
R254 B.n152 B.n133 585
R255 B.n150 B.n149 585
R256 B.n148 B.n134 585
R257 B.n147 B.n146 585
R258 B.n144 B.n135 585
R259 B.n142 B.n141 585
R260 B.n140 B.n136 585
R261 B.n139 B.n138 585
R262 B.n102 B.n101 585
R263 B.n103 B.n102 585
R264 B.n248 B.n247 585
R265 B.n249 B.n248 585
R266 B.n98 B.n97 585
R267 B.n99 B.n98 585
R268 B.n257 B.n256 585
R269 B.n256 B.n255 585
R270 B.n258 B.n96 585
R271 B.n96 B.n95 585
R272 B.n260 B.n259 585
R273 B.n261 B.n260 585
R274 B.n90 B.n89 585
R275 B.n91 B.n90 585
R276 B.n269 B.n268 585
R277 B.n268 B.n267 585
R278 B.n270 B.n88 585
R279 B.n88 B.n86 585
R280 B.n272 B.n271 585
R281 B.n273 B.n272 585
R282 B.n82 B.n81 585
R283 B.n87 B.n82 585
R284 B.n282 B.n281 585
R285 B.n281 B.n280 585
R286 B.n283 B.n80 585
R287 B.n279 B.n80 585
R288 B.n285 B.n284 585
R289 B.n286 B.n285 585
R290 B.n75 B.n74 585
R291 B.n79 B.n75 585
R292 B.n296 B.n295 585
R293 B.n295 B.n294 585
R294 B.n297 B.n73 585
R295 B.n293 B.n73 585
R296 B.n299 B.n298 585
R297 B.n300 B.n299 585
R298 B.n3 B.n0 585
R299 B.n4 B.n3 585
R300 B.n476 B.n1 585
R301 B.n477 B.n476 585
R302 B.n475 B.n474 585
R303 B.n475 B.n8 585
R304 B.n473 B.n9 585
R305 B.n12 B.n9 585
R306 B.n472 B.n471 585
R307 B.n471 B.n470 585
R308 B.n11 B.n10 585
R309 B.n469 B.n11 585
R310 B.n467 B.n466 585
R311 B.n468 B.n467 585
R312 B.n465 B.n16 585
R313 B.n19 B.n16 585
R314 B.n464 B.n463 585
R315 B.n463 B.n462 585
R316 B.n18 B.n17 585
R317 B.n461 B.n18 585
R318 B.n459 B.n458 585
R319 B.n460 B.n459 585
R320 B.n457 B.n24 585
R321 B.n24 B.n23 585
R322 B.n456 B.n455 585
R323 B.n455 B.n454 585
R324 B.n26 B.n25 585
R325 B.n453 B.n26 585
R326 B.n451 B.n450 585
R327 B.n452 B.n451 585
R328 B.n449 B.n31 585
R329 B.n31 B.n30 585
R330 B.n448 B.n447 585
R331 B.n447 B.n446 585
R332 B.n33 B.n32 585
R333 B.n445 B.n33 585
R334 B.n443 B.n442 585
R335 B.n444 B.n443 585
R336 B.n480 B.n479 585
R337 B.n478 B.n2 585
R338 B.n51 B.t15 583.866
R339 B.n58 B.t7 583.866
R340 B.n123 B.t18 583.866
R341 B.n117 B.t11 583.866
R342 B.n443 B.n38 478.086
R343 B.n330 B.n36 478.086
R344 B.n250 B.n102 478.086
R345 B.n248 B.n104 478.086
R346 B.n331 B.n37 256.663
R347 B.n333 B.n37 256.663
R348 B.n339 B.n37 256.663
R349 B.n341 B.n37 256.663
R350 B.n347 B.n37 256.663
R351 B.n349 B.n37 256.663
R352 B.n355 B.n37 256.663
R353 B.n357 B.n37 256.663
R354 B.n363 B.n37 256.663
R355 B.n365 B.n37 256.663
R356 B.n371 B.n37 256.663
R357 B.n373 B.n37 256.663
R358 B.n380 B.n37 256.663
R359 B.n382 B.n37 256.663
R360 B.n388 B.n37 256.663
R361 B.n390 B.n37 256.663
R362 B.n396 B.n37 256.663
R363 B.n398 B.n37 256.663
R364 B.n404 B.n37 256.663
R365 B.n406 B.n37 256.663
R366 B.n412 B.n37 256.663
R367 B.n414 B.n37 256.663
R368 B.n420 B.n37 256.663
R369 B.n422 B.n37 256.663
R370 B.n428 B.n37 256.663
R371 B.n430 B.n37 256.663
R372 B.n436 B.n37 256.663
R373 B.n438 B.n37 256.663
R374 B.n243 B.n103 256.663
R375 B.n106 B.n103 256.663
R376 B.n236 B.n103 256.663
R377 B.n230 B.n103 256.663
R378 B.n228 B.n103 256.663
R379 B.n222 B.n103 256.663
R380 B.n220 B.n103 256.663
R381 B.n214 B.n103 256.663
R382 B.n212 B.n103 256.663
R383 B.n206 B.n103 256.663
R384 B.n204 B.n103 256.663
R385 B.n197 B.n103 256.663
R386 B.n195 B.n103 256.663
R387 B.n189 B.n103 256.663
R388 B.n187 B.n103 256.663
R389 B.n181 B.n103 256.663
R390 B.n126 B.n103 256.663
R391 B.n175 B.n103 256.663
R392 B.n169 B.n103 256.663
R393 B.n167 B.n103 256.663
R394 B.n161 B.n103 256.663
R395 B.n159 B.n103 256.663
R396 B.n153 B.n103 256.663
R397 B.n151 B.n103 256.663
R398 B.n145 B.n103 256.663
R399 B.n143 B.n103 256.663
R400 B.n137 B.n103 256.663
R401 B.n482 B.n481 256.663
R402 B.n439 B.n437 163.367
R403 B.n435 B.n40 163.367
R404 B.n431 B.n429 163.367
R405 B.n427 B.n42 163.367
R406 B.n423 B.n421 163.367
R407 B.n419 B.n44 163.367
R408 B.n415 B.n413 163.367
R409 B.n411 B.n46 163.367
R410 B.n407 B.n405 163.367
R411 B.n403 B.n48 163.367
R412 B.n399 B.n397 163.367
R413 B.n395 B.n50 163.367
R414 B.n391 B.n389 163.367
R415 B.n387 B.n55 163.367
R416 B.n383 B.n381 163.367
R417 B.n379 B.n57 163.367
R418 B.n374 B.n372 163.367
R419 B.n370 B.n61 163.367
R420 B.n366 B.n364 163.367
R421 B.n362 B.n63 163.367
R422 B.n358 B.n356 163.367
R423 B.n354 B.n65 163.367
R424 B.n350 B.n348 163.367
R425 B.n346 B.n67 163.367
R426 B.n342 B.n340 163.367
R427 B.n338 B.n69 163.367
R428 B.n334 B.n332 163.367
R429 B.n250 B.n100 163.367
R430 B.n254 B.n100 163.367
R431 B.n254 B.n94 163.367
R432 B.n262 B.n94 163.367
R433 B.n262 B.n92 163.367
R434 B.n266 B.n92 163.367
R435 B.n266 B.n85 163.367
R436 B.n274 B.n85 163.367
R437 B.n274 B.n83 163.367
R438 B.n278 B.n83 163.367
R439 B.n278 B.n78 163.367
R440 B.n287 B.n78 163.367
R441 B.n287 B.n76 163.367
R442 B.n292 B.n76 163.367
R443 B.n292 B.n72 163.367
R444 B.n301 B.n72 163.367
R445 B.n302 B.n301 163.367
R446 B.n302 B.n5 163.367
R447 B.n6 B.n5 163.367
R448 B.n7 B.n6 163.367
R449 B.n308 B.n7 163.367
R450 B.n309 B.n308 163.367
R451 B.n309 B.n13 163.367
R452 B.n14 B.n13 163.367
R453 B.n15 B.n14 163.367
R454 B.n314 B.n15 163.367
R455 B.n314 B.n20 163.367
R456 B.n21 B.n20 163.367
R457 B.n22 B.n21 163.367
R458 B.n319 B.n22 163.367
R459 B.n319 B.n27 163.367
R460 B.n28 B.n27 163.367
R461 B.n29 B.n28 163.367
R462 B.n324 B.n29 163.367
R463 B.n324 B.n34 163.367
R464 B.n35 B.n34 163.367
R465 B.n36 B.n35 163.367
R466 B.n244 B.n242 163.367
R467 B.n242 B.n241 163.367
R468 B.n238 B.n237 163.367
R469 B.n235 B.n108 163.367
R470 B.n231 B.n229 163.367
R471 B.n227 B.n110 163.367
R472 B.n223 B.n221 163.367
R473 B.n219 B.n112 163.367
R474 B.n215 B.n213 163.367
R475 B.n211 B.n114 163.367
R476 B.n207 B.n205 163.367
R477 B.n203 B.n116 163.367
R478 B.n198 B.n196 163.367
R479 B.n194 B.n120 163.367
R480 B.n190 B.n188 163.367
R481 B.n186 B.n122 163.367
R482 B.n182 B.n180 163.367
R483 B.n177 B.n176 163.367
R484 B.n174 B.n128 163.367
R485 B.n170 B.n168 163.367
R486 B.n166 B.n130 163.367
R487 B.n162 B.n160 163.367
R488 B.n158 B.n132 163.367
R489 B.n154 B.n152 163.367
R490 B.n150 B.n134 163.367
R491 B.n146 B.n144 163.367
R492 B.n142 B.n136 163.367
R493 B.n138 B.n102 163.367
R494 B.n248 B.n98 163.367
R495 B.n256 B.n98 163.367
R496 B.n256 B.n96 163.367
R497 B.n260 B.n96 163.367
R498 B.n260 B.n90 163.367
R499 B.n268 B.n90 163.367
R500 B.n268 B.n88 163.367
R501 B.n272 B.n88 163.367
R502 B.n272 B.n82 163.367
R503 B.n281 B.n82 163.367
R504 B.n281 B.n80 163.367
R505 B.n285 B.n80 163.367
R506 B.n285 B.n75 163.367
R507 B.n295 B.n75 163.367
R508 B.n295 B.n73 163.367
R509 B.n299 B.n73 163.367
R510 B.n299 B.n3 163.367
R511 B.n480 B.n3 163.367
R512 B.n476 B.n2 163.367
R513 B.n476 B.n475 163.367
R514 B.n475 B.n9 163.367
R515 B.n471 B.n9 163.367
R516 B.n471 B.n11 163.367
R517 B.n467 B.n11 163.367
R518 B.n467 B.n16 163.367
R519 B.n463 B.n16 163.367
R520 B.n463 B.n18 163.367
R521 B.n459 B.n18 163.367
R522 B.n459 B.n24 163.367
R523 B.n455 B.n24 163.367
R524 B.n455 B.n26 163.367
R525 B.n451 B.n26 163.367
R526 B.n451 B.n31 163.367
R527 B.n447 B.n31 163.367
R528 B.n447 B.n33 163.367
R529 B.n443 B.n33 163.367
R530 B.n249 B.n103 116.948
R531 B.n444 B.n37 116.948
R532 B.n58 B.t9 88.8199
R533 B.n123 B.t20 88.8199
R534 B.n51 B.t16 88.8141
R535 B.n117 B.t14 88.8141
R536 B.n59 B.t10 75.2441
R537 B.n124 B.t19 75.2441
R538 B.n52 B.t17 75.2383
R539 B.n118 B.t13 75.2383
R540 B.n438 B.n38 71.676
R541 B.n437 B.n436 71.676
R542 B.n430 B.n40 71.676
R543 B.n429 B.n428 71.676
R544 B.n422 B.n42 71.676
R545 B.n421 B.n420 71.676
R546 B.n414 B.n44 71.676
R547 B.n413 B.n412 71.676
R548 B.n406 B.n46 71.676
R549 B.n405 B.n404 71.676
R550 B.n398 B.n48 71.676
R551 B.n397 B.n396 71.676
R552 B.n390 B.n50 71.676
R553 B.n389 B.n388 71.676
R554 B.n382 B.n55 71.676
R555 B.n381 B.n380 71.676
R556 B.n373 B.n57 71.676
R557 B.n372 B.n371 71.676
R558 B.n365 B.n61 71.676
R559 B.n364 B.n363 71.676
R560 B.n357 B.n63 71.676
R561 B.n356 B.n355 71.676
R562 B.n349 B.n65 71.676
R563 B.n348 B.n347 71.676
R564 B.n341 B.n67 71.676
R565 B.n340 B.n339 71.676
R566 B.n333 B.n69 71.676
R567 B.n332 B.n331 71.676
R568 B.n331 B.n330 71.676
R569 B.n334 B.n333 71.676
R570 B.n339 B.n338 71.676
R571 B.n342 B.n341 71.676
R572 B.n347 B.n346 71.676
R573 B.n350 B.n349 71.676
R574 B.n355 B.n354 71.676
R575 B.n358 B.n357 71.676
R576 B.n363 B.n362 71.676
R577 B.n366 B.n365 71.676
R578 B.n371 B.n370 71.676
R579 B.n374 B.n373 71.676
R580 B.n380 B.n379 71.676
R581 B.n383 B.n382 71.676
R582 B.n388 B.n387 71.676
R583 B.n391 B.n390 71.676
R584 B.n396 B.n395 71.676
R585 B.n399 B.n398 71.676
R586 B.n404 B.n403 71.676
R587 B.n407 B.n406 71.676
R588 B.n412 B.n411 71.676
R589 B.n415 B.n414 71.676
R590 B.n420 B.n419 71.676
R591 B.n423 B.n422 71.676
R592 B.n428 B.n427 71.676
R593 B.n431 B.n430 71.676
R594 B.n436 B.n435 71.676
R595 B.n439 B.n438 71.676
R596 B.n243 B.n104 71.676
R597 B.n241 B.n106 71.676
R598 B.n237 B.n236 71.676
R599 B.n230 B.n108 71.676
R600 B.n229 B.n228 71.676
R601 B.n222 B.n110 71.676
R602 B.n221 B.n220 71.676
R603 B.n214 B.n112 71.676
R604 B.n213 B.n212 71.676
R605 B.n206 B.n114 71.676
R606 B.n205 B.n204 71.676
R607 B.n197 B.n116 71.676
R608 B.n196 B.n195 71.676
R609 B.n189 B.n120 71.676
R610 B.n188 B.n187 71.676
R611 B.n181 B.n122 71.676
R612 B.n180 B.n126 71.676
R613 B.n176 B.n175 71.676
R614 B.n169 B.n128 71.676
R615 B.n168 B.n167 71.676
R616 B.n161 B.n130 71.676
R617 B.n160 B.n159 71.676
R618 B.n153 B.n132 71.676
R619 B.n152 B.n151 71.676
R620 B.n145 B.n134 71.676
R621 B.n144 B.n143 71.676
R622 B.n137 B.n136 71.676
R623 B.n244 B.n243 71.676
R624 B.n238 B.n106 71.676
R625 B.n236 B.n235 71.676
R626 B.n231 B.n230 71.676
R627 B.n228 B.n227 71.676
R628 B.n223 B.n222 71.676
R629 B.n220 B.n219 71.676
R630 B.n215 B.n214 71.676
R631 B.n212 B.n211 71.676
R632 B.n207 B.n206 71.676
R633 B.n204 B.n203 71.676
R634 B.n198 B.n197 71.676
R635 B.n195 B.n194 71.676
R636 B.n190 B.n189 71.676
R637 B.n187 B.n186 71.676
R638 B.n182 B.n181 71.676
R639 B.n177 B.n126 71.676
R640 B.n175 B.n174 71.676
R641 B.n170 B.n169 71.676
R642 B.n167 B.n166 71.676
R643 B.n162 B.n161 71.676
R644 B.n159 B.n158 71.676
R645 B.n154 B.n153 71.676
R646 B.n151 B.n150 71.676
R647 B.n146 B.n145 71.676
R648 B.n143 B.n142 71.676
R649 B.n138 B.n137 71.676
R650 B.n481 B.n480 71.676
R651 B.n481 B.n2 71.676
R652 B.n249 B.n99 67.9696
R653 B.n255 B.n99 67.9696
R654 B.n255 B.n95 67.9696
R655 B.n261 B.n95 67.9696
R656 B.n267 B.n91 67.9696
R657 B.n267 B.n86 67.9696
R658 B.n273 B.n86 67.9696
R659 B.n273 B.n87 67.9696
R660 B.n280 B.n279 67.9696
R661 B.n286 B.n79 67.9696
R662 B.n294 B.n293 67.9696
R663 B.n300 B.n4 67.9696
R664 B.n479 B.n4 67.9696
R665 B.n479 B.n478 67.9696
R666 B.n478 B.n477 67.9696
R667 B.n477 B.n8 67.9696
R668 B.n470 B.n12 67.9696
R669 B.n469 B.n468 67.9696
R670 B.n462 B.n19 67.9696
R671 B.n461 B.n460 67.9696
R672 B.n460 B.n23 67.9696
R673 B.n454 B.n23 67.9696
R674 B.n454 B.n453 67.9696
R675 B.n452 B.n30 67.9696
R676 B.n446 B.n30 67.9696
R677 B.n446 B.n445 67.9696
R678 B.n445 B.n444 67.9696
R679 B.n53 B.n52 59.5399
R680 B.n376 B.n59 59.5399
R681 B.n125 B.n124 59.5399
R682 B.n201 B.n118 59.5399
R683 B.n293 B.t5 58.9737
R684 B.n12 B.t3 58.9737
R685 B.n79 B.t4 54.9755
R686 B.t6 B.n469 54.9755
R687 B.n279 B.t1 50.9773
R688 B.n19 B.t2 50.9773
R689 B.n87 B.t0 46.9791
R690 B.t21 B.n461 46.9791
R691 B.t12 B.n91 38.9828
R692 B.n453 B.t8 38.9828
R693 B.n247 B.n246 31.0639
R694 B.n251 B.n101 31.0639
R695 B.n329 B.n328 31.0639
R696 B.n442 B.n441 31.0639
R697 B.n261 B.t12 28.9873
R698 B.t8 B.n452 28.9873
R699 B.n280 B.t0 20.991
R700 B.n462 B.t21 20.991
R701 B B.n482 18.0485
R702 B.n286 B.t1 16.9928
R703 B.n468 B.t2 16.9928
R704 B.n52 B.n51 13.5763
R705 B.n59 B.n58 13.5763
R706 B.n124 B.n123 13.5763
R707 B.n118 B.n117 13.5763
R708 B.n294 B.t4 12.9946
R709 B.n470 B.t6 12.9946
R710 B.n247 B.n97 10.6151
R711 B.n257 B.n97 10.6151
R712 B.n258 B.n257 10.6151
R713 B.n259 B.n258 10.6151
R714 B.n259 B.n89 10.6151
R715 B.n269 B.n89 10.6151
R716 B.n270 B.n269 10.6151
R717 B.n271 B.n270 10.6151
R718 B.n271 B.n81 10.6151
R719 B.n282 B.n81 10.6151
R720 B.n283 B.n282 10.6151
R721 B.n284 B.n283 10.6151
R722 B.n284 B.n74 10.6151
R723 B.n296 B.n74 10.6151
R724 B.n297 B.n296 10.6151
R725 B.n298 B.n297 10.6151
R726 B.n298 B.n0 10.6151
R727 B.n246 B.n245 10.6151
R728 B.n245 B.n105 10.6151
R729 B.n240 B.n105 10.6151
R730 B.n240 B.n239 10.6151
R731 B.n239 B.n107 10.6151
R732 B.n234 B.n107 10.6151
R733 B.n234 B.n233 10.6151
R734 B.n233 B.n232 10.6151
R735 B.n232 B.n109 10.6151
R736 B.n226 B.n109 10.6151
R737 B.n226 B.n225 10.6151
R738 B.n225 B.n224 10.6151
R739 B.n224 B.n111 10.6151
R740 B.n218 B.n111 10.6151
R741 B.n218 B.n217 10.6151
R742 B.n217 B.n216 10.6151
R743 B.n216 B.n113 10.6151
R744 B.n210 B.n113 10.6151
R745 B.n210 B.n209 10.6151
R746 B.n209 B.n208 10.6151
R747 B.n208 B.n115 10.6151
R748 B.n202 B.n115 10.6151
R749 B.n200 B.n199 10.6151
R750 B.n199 B.n119 10.6151
R751 B.n193 B.n119 10.6151
R752 B.n193 B.n192 10.6151
R753 B.n192 B.n191 10.6151
R754 B.n191 B.n121 10.6151
R755 B.n185 B.n121 10.6151
R756 B.n185 B.n184 10.6151
R757 B.n184 B.n183 10.6151
R758 B.n179 B.n178 10.6151
R759 B.n178 B.n127 10.6151
R760 B.n173 B.n127 10.6151
R761 B.n173 B.n172 10.6151
R762 B.n172 B.n171 10.6151
R763 B.n171 B.n129 10.6151
R764 B.n165 B.n129 10.6151
R765 B.n165 B.n164 10.6151
R766 B.n164 B.n163 10.6151
R767 B.n163 B.n131 10.6151
R768 B.n157 B.n131 10.6151
R769 B.n157 B.n156 10.6151
R770 B.n156 B.n155 10.6151
R771 B.n155 B.n133 10.6151
R772 B.n149 B.n133 10.6151
R773 B.n149 B.n148 10.6151
R774 B.n148 B.n147 10.6151
R775 B.n147 B.n135 10.6151
R776 B.n141 B.n135 10.6151
R777 B.n141 B.n140 10.6151
R778 B.n140 B.n139 10.6151
R779 B.n139 B.n101 10.6151
R780 B.n252 B.n251 10.6151
R781 B.n253 B.n252 10.6151
R782 B.n253 B.n93 10.6151
R783 B.n263 B.n93 10.6151
R784 B.n264 B.n263 10.6151
R785 B.n265 B.n264 10.6151
R786 B.n265 B.n84 10.6151
R787 B.n275 B.n84 10.6151
R788 B.n276 B.n275 10.6151
R789 B.n277 B.n276 10.6151
R790 B.n277 B.n77 10.6151
R791 B.n288 B.n77 10.6151
R792 B.n289 B.n288 10.6151
R793 B.n291 B.n289 10.6151
R794 B.n291 B.n290 10.6151
R795 B.n290 B.n71 10.6151
R796 B.n303 B.n71 10.6151
R797 B.n304 B.n303 10.6151
R798 B.n305 B.n304 10.6151
R799 B.n306 B.n305 10.6151
R800 B.n307 B.n306 10.6151
R801 B.n310 B.n307 10.6151
R802 B.n311 B.n310 10.6151
R803 B.n312 B.n311 10.6151
R804 B.n313 B.n312 10.6151
R805 B.n315 B.n313 10.6151
R806 B.n316 B.n315 10.6151
R807 B.n317 B.n316 10.6151
R808 B.n318 B.n317 10.6151
R809 B.n320 B.n318 10.6151
R810 B.n321 B.n320 10.6151
R811 B.n322 B.n321 10.6151
R812 B.n323 B.n322 10.6151
R813 B.n325 B.n323 10.6151
R814 B.n326 B.n325 10.6151
R815 B.n327 B.n326 10.6151
R816 B.n328 B.n327 10.6151
R817 B.n474 B.n1 10.6151
R818 B.n474 B.n473 10.6151
R819 B.n473 B.n472 10.6151
R820 B.n472 B.n10 10.6151
R821 B.n466 B.n10 10.6151
R822 B.n466 B.n465 10.6151
R823 B.n465 B.n464 10.6151
R824 B.n464 B.n17 10.6151
R825 B.n458 B.n17 10.6151
R826 B.n458 B.n457 10.6151
R827 B.n457 B.n456 10.6151
R828 B.n456 B.n25 10.6151
R829 B.n450 B.n25 10.6151
R830 B.n450 B.n449 10.6151
R831 B.n449 B.n448 10.6151
R832 B.n448 B.n32 10.6151
R833 B.n442 B.n32 10.6151
R834 B.n441 B.n440 10.6151
R835 B.n440 B.n39 10.6151
R836 B.n434 B.n39 10.6151
R837 B.n434 B.n433 10.6151
R838 B.n433 B.n432 10.6151
R839 B.n432 B.n41 10.6151
R840 B.n426 B.n41 10.6151
R841 B.n426 B.n425 10.6151
R842 B.n425 B.n424 10.6151
R843 B.n424 B.n43 10.6151
R844 B.n418 B.n43 10.6151
R845 B.n418 B.n417 10.6151
R846 B.n417 B.n416 10.6151
R847 B.n416 B.n45 10.6151
R848 B.n410 B.n45 10.6151
R849 B.n410 B.n409 10.6151
R850 B.n409 B.n408 10.6151
R851 B.n408 B.n47 10.6151
R852 B.n402 B.n47 10.6151
R853 B.n402 B.n401 10.6151
R854 B.n401 B.n400 10.6151
R855 B.n400 B.n49 10.6151
R856 B.n394 B.n393 10.6151
R857 B.n393 B.n392 10.6151
R858 B.n392 B.n54 10.6151
R859 B.n386 B.n54 10.6151
R860 B.n386 B.n385 10.6151
R861 B.n385 B.n384 10.6151
R862 B.n384 B.n56 10.6151
R863 B.n378 B.n56 10.6151
R864 B.n378 B.n377 10.6151
R865 B.n375 B.n60 10.6151
R866 B.n369 B.n60 10.6151
R867 B.n369 B.n368 10.6151
R868 B.n368 B.n367 10.6151
R869 B.n367 B.n62 10.6151
R870 B.n361 B.n62 10.6151
R871 B.n361 B.n360 10.6151
R872 B.n360 B.n359 10.6151
R873 B.n359 B.n64 10.6151
R874 B.n353 B.n64 10.6151
R875 B.n353 B.n352 10.6151
R876 B.n352 B.n351 10.6151
R877 B.n351 B.n66 10.6151
R878 B.n345 B.n66 10.6151
R879 B.n345 B.n344 10.6151
R880 B.n344 B.n343 10.6151
R881 B.n343 B.n68 10.6151
R882 B.n337 B.n68 10.6151
R883 B.n337 B.n336 10.6151
R884 B.n336 B.n335 10.6151
R885 B.n335 B.n70 10.6151
R886 B.n329 B.n70 10.6151
R887 B.n202 B.n201 9.36635
R888 B.n179 B.n125 9.36635
R889 B.n53 B.n49 9.36635
R890 B.n376 B.n375 9.36635
R891 B.n300 B.t5 8.99641
R892 B.t3 B.n8 8.99641
R893 B.n482 B.n0 8.11757
R894 B.n482 B.n1 8.11757
R895 B.n201 B.n200 1.24928
R896 B.n183 B.n125 1.24928
R897 B.n394 B.n53 1.24928
R898 B.n377 B.n376 1.24928
R899 VN.n1 VN.t4 511.161
R900 VN.n7 VN.t6 511.161
R901 VN.n4 VN.t5 496.844
R902 VN.n10 VN.t7 496.844
R903 VN.n2 VN.t3 480.046
R904 VN.n3 VN.t2 480.046
R905 VN.n8 VN.t1 480.046
R906 VN.n9 VN.t0 480.046
R907 VN.n5 VN.n4 161.3
R908 VN.n11 VN.n10 161.3
R909 VN.n9 VN.n6 161.3
R910 VN.n3 VN.n0 161.3
R911 VN.n7 VN.n6 73.733
R912 VN.n1 VN.n0 73.733
R913 VN.n3 VN.n2 48.2005
R914 VN.n9 VN.n8 48.2005
R915 VN VN.n11 36.1918
R916 VN.n4 VN.n3 31.4035
R917 VN.n10 VN.n9 31.4035
R918 VN.n8 VN.n7 14.302
R919 VN.n2 VN.n1 14.302
R920 VN.n11 VN.n6 0.189894
R921 VN.n5 VN.n0 0.189894
R922 VN VN.n5 0.0516364
R923 VDD2.n2 VDD2.n1 69.8616
R924 VDD2.n2 VDD2.n0 69.8616
R925 VDD2 VDD2.n5 69.8589
R926 VDD2.n4 VDD2.n3 69.6155
R927 VDD2.n4 VDD2.n2 31.3705
R928 VDD2.n5 VDD2.t6 3.456
R929 VDD2.n5 VDD2.t1 3.456
R930 VDD2.n3 VDD2.t0 3.456
R931 VDD2.n3 VDD2.t7 3.456
R932 VDD2.n1 VDD2.t5 3.456
R933 VDD2.n1 VDD2.t2 3.456
R934 VDD2.n0 VDD2.t3 3.456
R935 VDD2.n0 VDD2.t4 3.456
R936 VDD2 VDD2.n4 0.360414
C0 VDD1 VP 2.1482f
C1 VDD1 VN 0.147305f
C2 VN VP 3.77215f
C3 VTAIL VDD2 8.11164f
C4 VDD1 VDD2 0.662907f
C5 VDD1 VTAIL 8.07218f
C6 VDD2 VP 0.281983f
C7 VDD2 VN 2.01378f
C8 VTAIL VP 1.93345f
C9 VTAIL VN 1.91934f
C10 VDD2 B 2.687836f
C11 VDD1 B 2.888746f
C12 VTAIL B 5.009248f
C13 VN B 6.21128f
C14 VP B 4.845546f
C15 VDD2.t3 B 0.138348f
C16 VDD2.t4 B 0.138348f
C17 VDD2.n0 B 1.14901f
C18 VDD2.t5 B 0.138348f
C19 VDD2.t2 B 0.138348f
C20 VDD2.n1 B 1.14901f
C21 VDD2.n2 B 1.95328f
C22 VDD2.t0 B 0.138348f
C23 VDD2.t7 B 0.138348f
C24 VDD2.n3 B 1.1478f
C25 VDD2.n4 B 2.04488f
C26 VDD2.t6 B 0.138348f
C27 VDD2.t1 B 0.138348f
C28 VDD2.n5 B 1.14898f
C29 VN.n0 B 0.13095f
C30 VN.t4 B 0.253028f
C31 VN.n1 B 0.115735f
C32 VN.t3 B 0.24586f
C33 VN.n2 B 0.125068f
C34 VN.t2 B 0.24586f
C35 VN.n3 B 0.125068f
C36 VN.t5 B 0.249699f
C37 VN.n4 B 0.118769f
C38 VN.n5 B 0.030917f
C39 VN.n6 B 0.13095f
C40 VN.t7 B 0.249699f
C41 VN.t1 B 0.24586f
C42 VN.t6 B 0.253028f
C43 VN.n7 B 0.115735f
C44 VN.n8 B 0.125068f
C45 VN.t0 B 0.24586f
C46 VN.n9 B 0.125068f
C47 VN.n10 B 0.118769f
C48 VN.n11 B 1.26837f
C49 VTAIL.t6 B 0.088463f
C50 VTAIL.t2 B 0.088463f
C51 VTAIL.n0 B 0.685465f
C52 VTAIL.n1 B 0.221082f
C53 VTAIL.t3 B 0.875361f
C54 VTAIL.n2 B 0.298362f
C55 VTAIL.t10 B 0.875361f
C56 VTAIL.n3 B 0.298362f
C57 VTAIL.t8 B 0.088463f
C58 VTAIL.t12 B 0.088463f
C59 VTAIL.n4 B 0.685465f
C60 VTAIL.n5 B 0.255407f
C61 VTAIL.t9 B 0.875361f
C62 VTAIL.n6 B 0.883118f
C63 VTAIL.t0 B 0.875365f
C64 VTAIL.n7 B 0.883115f
C65 VTAIL.t1 B 0.088463f
C66 VTAIL.t4 B 0.088463f
C67 VTAIL.n8 B 0.685469f
C68 VTAIL.n9 B 0.255404f
C69 VTAIL.t5 B 0.875365f
C70 VTAIL.n10 B 0.298358f
C71 VTAIL.t11 B 0.875365f
C72 VTAIL.n11 B 0.298358f
C73 VTAIL.t13 B 0.088463f
C74 VTAIL.t14 B 0.088463f
C75 VTAIL.n12 B 0.685469f
C76 VTAIL.n13 B 0.255404f
C77 VTAIL.t7 B 0.875361f
C78 VTAIL.n14 B 0.883118f
C79 VTAIL.t15 B 0.875361f
C80 VTAIL.n15 B 0.879455f
C81 VDD1.t1 B 0.138174f
C82 VDD1.t0 B 0.138174f
C83 VDD1.n0 B 1.14817f
C84 VDD1.t5 B 0.138174f
C85 VDD1.t3 B 0.138174f
C86 VDD1.n1 B 1.14756f
C87 VDD1.t7 B 0.138174f
C88 VDD1.t4 B 0.138174f
C89 VDD1.n2 B 1.14756f
C90 VDD1.n3 B 2.01657f
C91 VDD1.t6 B 0.138174f
C92 VDD1.t2 B 0.138174f
C93 VDD1.n4 B 1.14635f
C94 VDD1.n5 B 2.07782f
C95 VP.n0 B 0.040979f
C96 VP.t5 B 0.256484f
C97 VP.n1 B 0.121997f
C98 VP.n2 B 0.134508f
C99 VP.t0 B 0.252541f
C100 VP.t1 B 0.252541f
C101 VP.t3 B 0.259903f
C102 VP.n3 B 0.11888f
C103 VP.n4 B 0.128466f
C104 VP.n5 B 0.128466f
C105 VP.t7 B 0.256484f
C106 VP.n6 B 0.121997f
C107 VP.n7 B 1.27565f
C108 VP.n8 B 1.31678f
C109 VP.n9 B 0.040979f
C110 VP.t6 B 0.252541f
C111 VP.n10 B 0.128466f
C112 VP.t2 B 0.252541f
C113 VP.n11 B 0.128466f
C114 VP.t4 B 0.256484f
C115 VP.n12 B 0.121997f
C116 VP.n13 B 0.031757f
.ends

