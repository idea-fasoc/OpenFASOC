* NGSPICE file created from diff_pair_sample_0394.ext - technology: sky130A

.subckt diff_pair_sample_0394 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t1 VN.t0 VTAIL.t2 w_n1382_n2314# sky130_fd_pr__pfet_01v8 ad=2.6169 pd=14.2 as=2.6169 ps=14.2 w=6.71 l=0.7
X1 B.t11 B.t9 B.t10 w_n1382_n2314# sky130_fd_pr__pfet_01v8 ad=2.6169 pd=14.2 as=0 ps=0 w=6.71 l=0.7
X2 VDD1.t1 VP.t0 VTAIL.t1 w_n1382_n2314# sky130_fd_pr__pfet_01v8 ad=2.6169 pd=14.2 as=2.6169 ps=14.2 w=6.71 l=0.7
X3 B.t8 B.t6 B.t7 w_n1382_n2314# sky130_fd_pr__pfet_01v8 ad=2.6169 pd=14.2 as=0 ps=0 w=6.71 l=0.7
X4 B.t5 B.t3 B.t4 w_n1382_n2314# sky130_fd_pr__pfet_01v8 ad=2.6169 pd=14.2 as=0 ps=0 w=6.71 l=0.7
X5 VDD2.t0 VN.t1 VTAIL.t3 w_n1382_n2314# sky130_fd_pr__pfet_01v8 ad=2.6169 pd=14.2 as=2.6169 ps=14.2 w=6.71 l=0.7
X6 B.t2 B.t0 B.t1 w_n1382_n2314# sky130_fd_pr__pfet_01v8 ad=2.6169 pd=14.2 as=0 ps=0 w=6.71 l=0.7
X7 VDD1.t0 VP.t1 VTAIL.t0 w_n1382_n2314# sky130_fd_pr__pfet_01v8 ad=2.6169 pd=14.2 as=2.6169 ps=14.2 w=6.71 l=0.7
R0 VN VN.t1 484.784
R1 VN VN.t0 448.83
R2 VTAIL.n138 VTAIL.n108 756.745
R3 VTAIL.n30 VTAIL.n0 756.745
R4 VTAIL.n102 VTAIL.n72 756.745
R5 VTAIL.n66 VTAIL.n36 756.745
R6 VTAIL.n121 VTAIL.n120 585
R7 VTAIL.n123 VTAIL.n122 585
R8 VTAIL.n116 VTAIL.n115 585
R9 VTAIL.n129 VTAIL.n128 585
R10 VTAIL.n131 VTAIL.n130 585
R11 VTAIL.n112 VTAIL.n111 585
R12 VTAIL.n137 VTAIL.n136 585
R13 VTAIL.n139 VTAIL.n138 585
R14 VTAIL.n13 VTAIL.n12 585
R15 VTAIL.n15 VTAIL.n14 585
R16 VTAIL.n8 VTAIL.n7 585
R17 VTAIL.n21 VTAIL.n20 585
R18 VTAIL.n23 VTAIL.n22 585
R19 VTAIL.n4 VTAIL.n3 585
R20 VTAIL.n29 VTAIL.n28 585
R21 VTAIL.n31 VTAIL.n30 585
R22 VTAIL.n103 VTAIL.n102 585
R23 VTAIL.n101 VTAIL.n100 585
R24 VTAIL.n76 VTAIL.n75 585
R25 VTAIL.n95 VTAIL.n94 585
R26 VTAIL.n93 VTAIL.n92 585
R27 VTAIL.n80 VTAIL.n79 585
R28 VTAIL.n87 VTAIL.n86 585
R29 VTAIL.n85 VTAIL.n84 585
R30 VTAIL.n67 VTAIL.n66 585
R31 VTAIL.n65 VTAIL.n64 585
R32 VTAIL.n40 VTAIL.n39 585
R33 VTAIL.n59 VTAIL.n58 585
R34 VTAIL.n57 VTAIL.n56 585
R35 VTAIL.n44 VTAIL.n43 585
R36 VTAIL.n51 VTAIL.n50 585
R37 VTAIL.n49 VTAIL.n48 585
R38 VTAIL.n119 VTAIL.t2 327.514
R39 VTAIL.n11 VTAIL.t0 327.514
R40 VTAIL.n83 VTAIL.t1 327.514
R41 VTAIL.n47 VTAIL.t3 327.514
R42 VTAIL.n122 VTAIL.n121 171.744
R43 VTAIL.n122 VTAIL.n115 171.744
R44 VTAIL.n129 VTAIL.n115 171.744
R45 VTAIL.n130 VTAIL.n129 171.744
R46 VTAIL.n130 VTAIL.n111 171.744
R47 VTAIL.n137 VTAIL.n111 171.744
R48 VTAIL.n138 VTAIL.n137 171.744
R49 VTAIL.n14 VTAIL.n13 171.744
R50 VTAIL.n14 VTAIL.n7 171.744
R51 VTAIL.n21 VTAIL.n7 171.744
R52 VTAIL.n22 VTAIL.n21 171.744
R53 VTAIL.n22 VTAIL.n3 171.744
R54 VTAIL.n29 VTAIL.n3 171.744
R55 VTAIL.n30 VTAIL.n29 171.744
R56 VTAIL.n102 VTAIL.n101 171.744
R57 VTAIL.n101 VTAIL.n75 171.744
R58 VTAIL.n94 VTAIL.n75 171.744
R59 VTAIL.n94 VTAIL.n93 171.744
R60 VTAIL.n93 VTAIL.n79 171.744
R61 VTAIL.n86 VTAIL.n79 171.744
R62 VTAIL.n86 VTAIL.n85 171.744
R63 VTAIL.n66 VTAIL.n65 171.744
R64 VTAIL.n65 VTAIL.n39 171.744
R65 VTAIL.n58 VTAIL.n39 171.744
R66 VTAIL.n58 VTAIL.n57 171.744
R67 VTAIL.n57 VTAIL.n43 171.744
R68 VTAIL.n50 VTAIL.n43 171.744
R69 VTAIL.n50 VTAIL.n49 171.744
R70 VTAIL.n121 VTAIL.t2 85.8723
R71 VTAIL.n13 VTAIL.t0 85.8723
R72 VTAIL.n85 VTAIL.t1 85.8723
R73 VTAIL.n49 VTAIL.t3 85.8723
R74 VTAIL.n143 VTAIL.n142 31.9914
R75 VTAIL.n35 VTAIL.n34 31.9914
R76 VTAIL.n107 VTAIL.n106 31.9914
R77 VTAIL.n71 VTAIL.n70 31.9914
R78 VTAIL.n71 VTAIL.n35 19.9445
R79 VTAIL.n143 VTAIL.n107 19.0565
R80 VTAIL.n120 VTAIL.n119 16.3884
R81 VTAIL.n12 VTAIL.n11 16.3884
R82 VTAIL.n84 VTAIL.n83 16.3884
R83 VTAIL.n48 VTAIL.n47 16.3884
R84 VTAIL.n123 VTAIL.n118 12.8005
R85 VTAIL.n15 VTAIL.n10 12.8005
R86 VTAIL.n87 VTAIL.n82 12.8005
R87 VTAIL.n51 VTAIL.n46 12.8005
R88 VTAIL.n124 VTAIL.n116 12.0247
R89 VTAIL.n16 VTAIL.n8 12.0247
R90 VTAIL.n88 VTAIL.n80 12.0247
R91 VTAIL.n52 VTAIL.n44 12.0247
R92 VTAIL.n128 VTAIL.n127 11.249
R93 VTAIL.n20 VTAIL.n19 11.249
R94 VTAIL.n92 VTAIL.n91 11.249
R95 VTAIL.n56 VTAIL.n55 11.249
R96 VTAIL.n131 VTAIL.n114 10.4732
R97 VTAIL.n23 VTAIL.n6 10.4732
R98 VTAIL.n95 VTAIL.n78 10.4732
R99 VTAIL.n59 VTAIL.n42 10.4732
R100 VTAIL.n132 VTAIL.n112 9.69747
R101 VTAIL.n24 VTAIL.n4 9.69747
R102 VTAIL.n96 VTAIL.n76 9.69747
R103 VTAIL.n60 VTAIL.n40 9.69747
R104 VTAIL.n142 VTAIL.n141 9.45567
R105 VTAIL.n34 VTAIL.n33 9.45567
R106 VTAIL.n106 VTAIL.n105 9.45567
R107 VTAIL.n70 VTAIL.n69 9.45567
R108 VTAIL.n110 VTAIL.n109 9.3005
R109 VTAIL.n135 VTAIL.n134 9.3005
R110 VTAIL.n133 VTAIL.n132 9.3005
R111 VTAIL.n114 VTAIL.n113 9.3005
R112 VTAIL.n127 VTAIL.n126 9.3005
R113 VTAIL.n125 VTAIL.n124 9.3005
R114 VTAIL.n118 VTAIL.n117 9.3005
R115 VTAIL.n141 VTAIL.n140 9.3005
R116 VTAIL.n2 VTAIL.n1 9.3005
R117 VTAIL.n27 VTAIL.n26 9.3005
R118 VTAIL.n25 VTAIL.n24 9.3005
R119 VTAIL.n6 VTAIL.n5 9.3005
R120 VTAIL.n19 VTAIL.n18 9.3005
R121 VTAIL.n17 VTAIL.n16 9.3005
R122 VTAIL.n10 VTAIL.n9 9.3005
R123 VTAIL.n33 VTAIL.n32 9.3005
R124 VTAIL.n105 VTAIL.n104 9.3005
R125 VTAIL.n74 VTAIL.n73 9.3005
R126 VTAIL.n99 VTAIL.n98 9.3005
R127 VTAIL.n97 VTAIL.n96 9.3005
R128 VTAIL.n78 VTAIL.n77 9.3005
R129 VTAIL.n91 VTAIL.n90 9.3005
R130 VTAIL.n89 VTAIL.n88 9.3005
R131 VTAIL.n82 VTAIL.n81 9.3005
R132 VTAIL.n69 VTAIL.n68 9.3005
R133 VTAIL.n38 VTAIL.n37 9.3005
R134 VTAIL.n63 VTAIL.n62 9.3005
R135 VTAIL.n61 VTAIL.n60 9.3005
R136 VTAIL.n42 VTAIL.n41 9.3005
R137 VTAIL.n55 VTAIL.n54 9.3005
R138 VTAIL.n53 VTAIL.n52 9.3005
R139 VTAIL.n46 VTAIL.n45 9.3005
R140 VTAIL.n136 VTAIL.n135 8.92171
R141 VTAIL.n28 VTAIL.n27 8.92171
R142 VTAIL.n100 VTAIL.n99 8.92171
R143 VTAIL.n64 VTAIL.n63 8.92171
R144 VTAIL.n139 VTAIL.n110 8.14595
R145 VTAIL.n31 VTAIL.n2 8.14595
R146 VTAIL.n103 VTAIL.n74 8.14595
R147 VTAIL.n67 VTAIL.n38 8.14595
R148 VTAIL.n140 VTAIL.n108 7.3702
R149 VTAIL.n32 VTAIL.n0 7.3702
R150 VTAIL.n104 VTAIL.n72 7.3702
R151 VTAIL.n68 VTAIL.n36 7.3702
R152 VTAIL.n142 VTAIL.n108 6.59444
R153 VTAIL.n34 VTAIL.n0 6.59444
R154 VTAIL.n106 VTAIL.n72 6.59444
R155 VTAIL.n70 VTAIL.n36 6.59444
R156 VTAIL.n140 VTAIL.n139 5.81868
R157 VTAIL.n32 VTAIL.n31 5.81868
R158 VTAIL.n104 VTAIL.n103 5.81868
R159 VTAIL.n68 VTAIL.n67 5.81868
R160 VTAIL.n136 VTAIL.n110 5.04292
R161 VTAIL.n28 VTAIL.n2 5.04292
R162 VTAIL.n100 VTAIL.n74 5.04292
R163 VTAIL.n64 VTAIL.n38 5.04292
R164 VTAIL.n135 VTAIL.n112 4.26717
R165 VTAIL.n27 VTAIL.n4 4.26717
R166 VTAIL.n99 VTAIL.n76 4.26717
R167 VTAIL.n63 VTAIL.n40 4.26717
R168 VTAIL.n119 VTAIL.n117 3.71088
R169 VTAIL.n11 VTAIL.n9 3.71088
R170 VTAIL.n83 VTAIL.n81 3.71088
R171 VTAIL.n47 VTAIL.n45 3.71088
R172 VTAIL.n132 VTAIL.n131 3.49141
R173 VTAIL.n24 VTAIL.n23 3.49141
R174 VTAIL.n96 VTAIL.n95 3.49141
R175 VTAIL.n60 VTAIL.n59 3.49141
R176 VTAIL.n128 VTAIL.n114 2.71565
R177 VTAIL.n20 VTAIL.n6 2.71565
R178 VTAIL.n92 VTAIL.n78 2.71565
R179 VTAIL.n56 VTAIL.n42 2.71565
R180 VTAIL.n127 VTAIL.n116 1.93989
R181 VTAIL.n19 VTAIL.n8 1.93989
R182 VTAIL.n91 VTAIL.n80 1.93989
R183 VTAIL.n55 VTAIL.n44 1.93989
R184 VTAIL.n124 VTAIL.n123 1.16414
R185 VTAIL.n16 VTAIL.n15 1.16414
R186 VTAIL.n88 VTAIL.n87 1.16414
R187 VTAIL.n52 VTAIL.n51 1.16414
R188 VTAIL.n107 VTAIL.n71 0.914293
R189 VTAIL VTAIL.n35 0.7505
R190 VTAIL.n120 VTAIL.n118 0.388379
R191 VTAIL.n12 VTAIL.n10 0.388379
R192 VTAIL.n84 VTAIL.n82 0.388379
R193 VTAIL.n48 VTAIL.n46 0.388379
R194 VTAIL VTAIL.n143 0.164293
R195 VTAIL.n125 VTAIL.n117 0.155672
R196 VTAIL.n126 VTAIL.n125 0.155672
R197 VTAIL.n126 VTAIL.n113 0.155672
R198 VTAIL.n133 VTAIL.n113 0.155672
R199 VTAIL.n134 VTAIL.n133 0.155672
R200 VTAIL.n134 VTAIL.n109 0.155672
R201 VTAIL.n141 VTAIL.n109 0.155672
R202 VTAIL.n17 VTAIL.n9 0.155672
R203 VTAIL.n18 VTAIL.n17 0.155672
R204 VTAIL.n18 VTAIL.n5 0.155672
R205 VTAIL.n25 VTAIL.n5 0.155672
R206 VTAIL.n26 VTAIL.n25 0.155672
R207 VTAIL.n26 VTAIL.n1 0.155672
R208 VTAIL.n33 VTAIL.n1 0.155672
R209 VTAIL.n105 VTAIL.n73 0.155672
R210 VTAIL.n98 VTAIL.n73 0.155672
R211 VTAIL.n98 VTAIL.n97 0.155672
R212 VTAIL.n97 VTAIL.n77 0.155672
R213 VTAIL.n90 VTAIL.n77 0.155672
R214 VTAIL.n90 VTAIL.n89 0.155672
R215 VTAIL.n89 VTAIL.n81 0.155672
R216 VTAIL.n69 VTAIL.n37 0.155672
R217 VTAIL.n62 VTAIL.n37 0.155672
R218 VTAIL.n62 VTAIL.n61 0.155672
R219 VTAIL.n61 VTAIL.n41 0.155672
R220 VTAIL.n54 VTAIL.n41 0.155672
R221 VTAIL.n54 VTAIL.n53 0.155672
R222 VTAIL.n53 VTAIL.n45 0.155672
R223 VDD2.n65 VDD2.n35 756.745
R224 VDD2.n30 VDD2.n0 756.745
R225 VDD2.n66 VDD2.n65 585
R226 VDD2.n64 VDD2.n63 585
R227 VDD2.n39 VDD2.n38 585
R228 VDD2.n58 VDD2.n57 585
R229 VDD2.n56 VDD2.n55 585
R230 VDD2.n43 VDD2.n42 585
R231 VDD2.n50 VDD2.n49 585
R232 VDD2.n48 VDD2.n47 585
R233 VDD2.n13 VDD2.n12 585
R234 VDD2.n15 VDD2.n14 585
R235 VDD2.n8 VDD2.n7 585
R236 VDD2.n21 VDD2.n20 585
R237 VDD2.n23 VDD2.n22 585
R238 VDD2.n4 VDD2.n3 585
R239 VDD2.n29 VDD2.n28 585
R240 VDD2.n31 VDD2.n30 585
R241 VDD2.n46 VDD2.t0 327.514
R242 VDD2.n11 VDD2.t1 327.514
R243 VDD2.n65 VDD2.n64 171.744
R244 VDD2.n64 VDD2.n38 171.744
R245 VDD2.n57 VDD2.n38 171.744
R246 VDD2.n57 VDD2.n56 171.744
R247 VDD2.n56 VDD2.n42 171.744
R248 VDD2.n49 VDD2.n42 171.744
R249 VDD2.n49 VDD2.n48 171.744
R250 VDD2.n14 VDD2.n13 171.744
R251 VDD2.n14 VDD2.n7 171.744
R252 VDD2.n21 VDD2.n7 171.744
R253 VDD2.n22 VDD2.n21 171.744
R254 VDD2.n22 VDD2.n3 171.744
R255 VDD2.n29 VDD2.n3 171.744
R256 VDD2.n30 VDD2.n29 171.744
R257 VDD2.n48 VDD2.t0 85.8723
R258 VDD2.n13 VDD2.t1 85.8723
R259 VDD2.n70 VDD2.n34 79.9072
R260 VDD2.n70 VDD2.n69 48.6702
R261 VDD2.n12 VDD2.n11 16.3884
R262 VDD2.n47 VDD2.n46 16.3884
R263 VDD2.n50 VDD2.n45 12.8005
R264 VDD2.n15 VDD2.n10 12.8005
R265 VDD2.n51 VDD2.n43 12.0247
R266 VDD2.n16 VDD2.n8 12.0247
R267 VDD2.n55 VDD2.n54 11.249
R268 VDD2.n20 VDD2.n19 11.249
R269 VDD2.n58 VDD2.n41 10.4732
R270 VDD2.n23 VDD2.n6 10.4732
R271 VDD2.n59 VDD2.n39 9.69747
R272 VDD2.n24 VDD2.n4 9.69747
R273 VDD2.n69 VDD2.n68 9.45567
R274 VDD2.n34 VDD2.n33 9.45567
R275 VDD2.n68 VDD2.n67 9.3005
R276 VDD2.n37 VDD2.n36 9.3005
R277 VDD2.n62 VDD2.n61 9.3005
R278 VDD2.n60 VDD2.n59 9.3005
R279 VDD2.n41 VDD2.n40 9.3005
R280 VDD2.n54 VDD2.n53 9.3005
R281 VDD2.n52 VDD2.n51 9.3005
R282 VDD2.n45 VDD2.n44 9.3005
R283 VDD2.n2 VDD2.n1 9.3005
R284 VDD2.n27 VDD2.n26 9.3005
R285 VDD2.n25 VDD2.n24 9.3005
R286 VDD2.n6 VDD2.n5 9.3005
R287 VDD2.n19 VDD2.n18 9.3005
R288 VDD2.n17 VDD2.n16 9.3005
R289 VDD2.n10 VDD2.n9 9.3005
R290 VDD2.n33 VDD2.n32 9.3005
R291 VDD2.n63 VDD2.n62 8.92171
R292 VDD2.n28 VDD2.n27 8.92171
R293 VDD2.n66 VDD2.n37 8.14595
R294 VDD2.n31 VDD2.n2 8.14595
R295 VDD2.n67 VDD2.n35 7.3702
R296 VDD2.n32 VDD2.n0 7.3702
R297 VDD2.n69 VDD2.n35 6.59444
R298 VDD2.n34 VDD2.n0 6.59444
R299 VDD2.n67 VDD2.n66 5.81868
R300 VDD2.n32 VDD2.n31 5.81868
R301 VDD2.n63 VDD2.n37 5.04292
R302 VDD2.n28 VDD2.n2 5.04292
R303 VDD2.n62 VDD2.n39 4.26717
R304 VDD2.n27 VDD2.n4 4.26717
R305 VDD2.n46 VDD2.n44 3.71088
R306 VDD2.n11 VDD2.n9 3.71088
R307 VDD2.n59 VDD2.n58 3.49141
R308 VDD2.n24 VDD2.n23 3.49141
R309 VDD2.n55 VDD2.n41 2.71565
R310 VDD2.n20 VDD2.n6 2.71565
R311 VDD2.n54 VDD2.n43 1.93989
R312 VDD2.n19 VDD2.n8 1.93989
R313 VDD2.n51 VDD2.n50 1.16414
R314 VDD2.n16 VDD2.n15 1.16414
R315 VDD2.n47 VDD2.n45 0.388379
R316 VDD2.n12 VDD2.n10 0.388379
R317 VDD2 VDD2.n70 0.280672
R318 VDD2.n68 VDD2.n36 0.155672
R319 VDD2.n61 VDD2.n36 0.155672
R320 VDD2.n61 VDD2.n60 0.155672
R321 VDD2.n60 VDD2.n40 0.155672
R322 VDD2.n53 VDD2.n40 0.155672
R323 VDD2.n53 VDD2.n52 0.155672
R324 VDD2.n52 VDD2.n44 0.155672
R325 VDD2.n17 VDD2.n9 0.155672
R326 VDD2.n18 VDD2.n17 0.155672
R327 VDD2.n18 VDD2.n5 0.155672
R328 VDD2.n25 VDD2.n5 0.155672
R329 VDD2.n26 VDD2.n25 0.155672
R330 VDD2.n26 VDD2.n1 0.155672
R331 VDD2.n33 VDD2.n1 0.155672
R332 B.n259 B.n44 585
R333 B.n261 B.n260 585
R334 B.n262 B.n43 585
R335 B.n264 B.n263 585
R336 B.n265 B.n42 585
R337 B.n267 B.n266 585
R338 B.n268 B.n41 585
R339 B.n270 B.n269 585
R340 B.n271 B.n40 585
R341 B.n273 B.n272 585
R342 B.n274 B.n39 585
R343 B.n276 B.n275 585
R344 B.n277 B.n38 585
R345 B.n279 B.n278 585
R346 B.n280 B.n37 585
R347 B.n282 B.n281 585
R348 B.n283 B.n36 585
R349 B.n285 B.n284 585
R350 B.n286 B.n35 585
R351 B.n288 B.n287 585
R352 B.n289 B.n34 585
R353 B.n291 B.n290 585
R354 B.n292 B.n33 585
R355 B.n294 B.n293 585
R356 B.n295 B.n32 585
R357 B.n297 B.n296 585
R358 B.n299 B.n29 585
R359 B.n301 B.n300 585
R360 B.n302 B.n28 585
R361 B.n304 B.n303 585
R362 B.n305 B.n27 585
R363 B.n307 B.n306 585
R364 B.n308 B.n26 585
R365 B.n310 B.n309 585
R366 B.n311 B.n25 585
R367 B.n313 B.n312 585
R368 B.n315 B.n314 585
R369 B.n316 B.n21 585
R370 B.n318 B.n317 585
R371 B.n319 B.n20 585
R372 B.n321 B.n320 585
R373 B.n322 B.n19 585
R374 B.n324 B.n323 585
R375 B.n325 B.n18 585
R376 B.n327 B.n326 585
R377 B.n328 B.n17 585
R378 B.n330 B.n329 585
R379 B.n331 B.n16 585
R380 B.n333 B.n332 585
R381 B.n334 B.n15 585
R382 B.n336 B.n335 585
R383 B.n337 B.n14 585
R384 B.n339 B.n338 585
R385 B.n340 B.n13 585
R386 B.n342 B.n341 585
R387 B.n343 B.n12 585
R388 B.n345 B.n344 585
R389 B.n346 B.n11 585
R390 B.n348 B.n347 585
R391 B.n349 B.n10 585
R392 B.n351 B.n350 585
R393 B.n352 B.n9 585
R394 B.n258 B.n257 585
R395 B.n256 B.n45 585
R396 B.n255 B.n254 585
R397 B.n253 B.n46 585
R398 B.n252 B.n251 585
R399 B.n250 B.n47 585
R400 B.n249 B.n248 585
R401 B.n247 B.n48 585
R402 B.n246 B.n245 585
R403 B.n244 B.n49 585
R404 B.n243 B.n242 585
R405 B.n241 B.n50 585
R406 B.n240 B.n239 585
R407 B.n238 B.n51 585
R408 B.n237 B.n236 585
R409 B.n235 B.n52 585
R410 B.n234 B.n233 585
R411 B.n232 B.n53 585
R412 B.n231 B.n230 585
R413 B.n229 B.n54 585
R414 B.n228 B.n227 585
R415 B.n226 B.n55 585
R416 B.n225 B.n224 585
R417 B.n223 B.n56 585
R418 B.n222 B.n221 585
R419 B.n220 B.n57 585
R420 B.n219 B.n218 585
R421 B.n217 B.n58 585
R422 B.n216 B.n215 585
R423 B.n121 B.n94 585
R424 B.n123 B.n122 585
R425 B.n124 B.n93 585
R426 B.n126 B.n125 585
R427 B.n127 B.n92 585
R428 B.n129 B.n128 585
R429 B.n130 B.n91 585
R430 B.n132 B.n131 585
R431 B.n133 B.n90 585
R432 B.n135 B.n134 585
R433 B.n136 B.n89 585
R434 B.n138 B.n137 585
R435 B.n139 B.n88 585
R436 B.n141 B.n140 585
R437 B.n142 B.n87 585
R438 B.n144 B.n143 585
R439 B.n145 B.n86 585
R440 B.n147 B.n146 585
R441 B.n148 B.n85 585
R442 B.n150 B.n149 585
R443 B.n151 B.n84 585
R444 B.n153 B.n152 585
R445 B.n154 B.n83 585
R446 B.n156 B.n155 585
R447 B.n157 B.n82 585
R448 B.n159 B.n158 585
R449 B.n161 B.n79 585
R450 B.n163 B.n162 585
R451 B.n164 B.n78 585
R452 B.n166 B.n165 585
R453 B.n167 B.n77 585
R454 B.n169 B.n168 585
R455 B.n170 B.n76 585
R456 B.n172 B.n171 585
R457 B.n173 B.n75 585
R458 B.n175 B.n174 585
R459 B.n177 B.n176 585
R460 B.n178 B.n71 585
R461 B.n180 B.n179 585
R462 B.n181 B.n70 585
R463 B.n183 B.n182 585
R464 B.n184 B.n69 585
R465 B.n186 B.n185 585
R466 B.n187 B.n68 585
R467 B.n189 B.n188 585
R468 B.n190 B.n67 585
R469 B.n192 B.n191 585
R470 B.n193 B.n66 585
R471 B.n195 B.n194 585
R472 B.n196 B.n65 585
R473 B.n198 B.n197 585
R474 B.n199 B.n64 585
R475 B.n201 B.n200 585
R476 B.n202 B.n63 585
R477 B.n204 B.n203 585
R478 B.n205 B.n62 585
R479 B.n207 B.n206 585
R480 B.n208 B.n61 585
R481 B.n210 B.n209 585
R482 B.n211 B.n60 585
R483 B.n213 B.n212 585
R484 B.n214 B.n59 585
R485 B.n120 B.n119 585
R486 B.n118 B.n95 585
R487 B.n117 B.n116 585
R488 B.n115 B.n96 585
R489 B.n114 B.n113 585
R490 B.n112 B.n97 585
R491 B.n111 B.n110 585
R492 B.n109 B.n98 585
R493 B.n108 B.n107 585
R494 B.n106 B.n99 585
R495 B.n105 B.n104 585
R496 B.n103 B.n100 585
R497 B.n102 B.n101 585
R498 B.n2 B.n0 585
R499 B.n373 B.n1 585
R500 B.n372 B.n371 585
R501 B.n370 B.n3 585
R502 B.n369 B.n368 585
R503 B.n367 B.n4 585
R504 B.n366 B.n365 585
R505 B.n364 B.n5 585
R506 B.n363 B.n362 585
R507 B.n361 B.n6 585
R508 B.n360 B.n359 585
R509 B.n358 B.n7 585
R510 B.n357 B.n356 585
R511 B.n355 B.n8 585
R512 B.n354 B.n353 585
R513 B.n375 B.n374 585
R514 B.n121 B.n120 511.721
R515 B.n354 B.n9 511.721
R516 B.n216 B.n59 511.721
R517 B.n259 B.n258 511.721
R518 B.n72 B.t3 433.981
R519 B.n80 B.t0 433.981
R520 B.n22 B.t6 433.981
R521 B.n30 B.t9 433.981
R522 B.n72 B.t5 300.745
R523 B.n30 B.t10 300.745
R524 B.n80 B.t2 300.745
R525 B.n22 B.t7 300.745
R526 B.n73 B.t4 280.769
R527 B.n31 B.t11 280.769
R528 B.n81 B.t1 280.769
R529 B.n23 B.t8 280.769
R530 B.n120 B.n95 163.367
R531 B.n116 B.n95 163.367
R532 B.n116 B.n115 163.367
R533 B.n115 B.n114 163.367
R534 B.n114 B.n97 163.367
R535 B.n110 B.n97 163.367
R536 B.n110 B.n109 163.367
R537 B.n109 B.n108 163.367
R538 B.n108 B.n99 163.367
R539 B.n104 B.n99 163.367
R540 B.n104 B.n103 163.367
R541 B.n103 B.n102 163.367
R542 B.n102 B.n2 163.367
R543 B.n374 B.n2 163.367
R544 B.n374 B.n373 163.367
R545 B.n373 B.n372 163.367
R546 B.n372 B.n3 163.367
R547 B.n368 B.n3 163.367
R548 B.n368 B.n367 163.367
R549 B.n367 B.n366 163.367
R550 B.n366 B.n5 163.367
R551 B.n362 B.n5 163.367
R552 B.n362 B.n361 163.367
R553 B.n361 B.n360 163.367
R554 B.n360 B.n7 163.367
R555 B.n356 B.n7 163.367
R556 B.n356 B.n355 163.367
R557 B.n355 B.n354 163.367
R558 B.n122 B.n121 163.367
R559 B.n122 B.n93 163.367
R560 B.n126 B.n93 163.367
R561 B.n127 B.n126 163.367
R562 B.n128 B.n127 163.367
R563 B.n128 B.n91 163.367
R564 B.n132 B.n91 163.367
R565 B.n133 B.n132 163.367
R566 B.n134 B.n133 163.367
R567 B.n134 B.n89 163.367
R568 B.n138 B.n89 163.367
R569 B.n139 B.n138 163.367
R570 B.n140 B.n139 163.367
R571 B.n140 B.n87 163.367
R572 B.n144 B.n87 163.367
R573 B.n145 B.n144 163.367
R574 B.n146 B.n145 163.367
R575 B.n146 B.n85 163.367
R576 B.n150 B.n85 163.367
R577 B.n151 B.n150 163.367
R578 B.n152 B.n151 163.367
R579 B.n152 B.n83 163.367
R580 B.n156 B.n83 163.367
R581 B.n157 B.n156 163.367
R582 B.n158 B.n157 163.367
R583 B.n158 B.n79 163.367
R584 B.n163 B.n79 163.367
R585 B.n164 B.n163 163.367
R586 B.n165 B.n164 163.367
R587 B.n165 B.n77 163.367
R588 B.n169 B.n77 163.367
R589 B.n170 B.n169 163.367
R590 B.n171 B.n170 163.367
R591 B.n171 B.n75 163.367
R592 B.n175 B.n75 163.367
R593 B.n176 B.n175 163.367
R594 B.n176 B.n71 163.367
R595 B.n180 B.n71 163.367
R596 B.n181 B.n180 163.367
R597 B.n182 B.n181 163.367
R598 B.n182 B.n69 163.367
R599 B.n186 B.n69 163.367
R600 B.n187 B.n186 163.367
R601 B.n188 B.n187 163.367
R602 B.n188 B.n67 163.367
R603 B.n192 B.n67 163.367
R604 B.n193 B.n192 163.367
R605 B.n194 B.n193 163.367
R606 B.n194 B.n65 163.367
R607 B.n198 B.n65 163.367
R608 B.n199 B.n198 163.367
R609 B.n200 B.n199 163.367
R610 B.n200 B.n63 163.367
R611 B.n204 B.n63 163.367
R612 B.n205 B.n204 163.367
R613 B.n206 B.n205 163.367
R614 B.n206 B.n61 163.367
R615 B.n210 B.n61 163.367
R616 B.n211 B.n210 163.367
R617 B.n212 B.n211 163.367
R618 B.n212 B.n59 163.367
R619 B.n217 B.n216 163.367
R620 B.n218 B.n217 163.367
R621 B.n218 B.n57 163.367
R622 B.n222 B.n57 163.367
R623 B.n223 B.n222 163.367
R624 B.n224 B.n223 163.367
R625 B.n224 B.n55 163.367
R626 B.n228 B.n55 163.367
R627 B.n229 B.n228 163.367
R628 B.n230 B.n229 163.367
R629 B.n230 B.n53 163.367
R630 B.n234 B.n53 163.367
R631 B.n235 B.n234 163.367
R632 B.n236 B.n235 163.367
R633 B.n236 B.n51 163.367
R634 B.n240 B.n51 163.367
R635 B.n241 B.n240 163.367
R636 B.n242 B.n241 163.367
R637 B.n242 B.n49 163.367
R638 B.n246 B.n49 163.367
R639 B.n247 B.n246 163.367
R640 B.n248 B.n247 163.367
R641 B.n248 B.n47 163.367
R642 B.n252 B.n47 163.367
R643 B.n253 B.n252 163.367
R644 B.n254 B.n253 163.367
R645 B.n254 B.n45 163.367
R646 B.n258 B.n45 163.367
R647 B.n350 B.n9 163.367
R648 B.n350 B.n349 163.367
R649 B.n349 B.n348 163.367
R650 B.n348 B.n11 163.367
R651 B.n344 B.n11 163.367
R652 B.n344 B.n343 163.367
R653 B.n343 B.n342 163.367
R654 B.n342 B.n13 163.367
R655 B.n338 B.n13 163.367
R656 B.n338 B.n337 163.367
R657 B.n337 B.n336 163.367
R658 B.n336 B.n15 163.367
R659 B.n332 B.n15 163.367
R660 B.n332 B.n331 163.367
R661 B.n331 B.n330 163.367
R662 B.n330 B.n17 163.367
R663 B.n326 B.n17 163.367
R664 B.n326 B.n325 163.367
R665 B.n325 B.n324 163.367
R666 B.n324 B.n19 163.367
R667 B.n320 B.n19 163.367
R668 B.n320 B.n319 163.367
R669 B.n319 B.n318 163.367
R670 B.n318 B.n21 163.367
R671 B.n314 B.n21 163.367
R672 B.n314 B.n313 163.367
R673 B.n313 B.n25 163.367
R674 B.n309 B.n25 163.367
R675 B.n309 B.n308 163.367
R676 B.n308 B.n307 163.367
R677 B.n307 B.n27 163.367
R678 B.n303 B.n27 163.367
R679 B.n303 B.n302 163.367
R680 B.n302 B.n301 163.367
R681 B.n301 B.n29 163.367
R682 B.n296 B.n29 163.367
R683 B.n296 B.n295 163.367
R684 B.n295 B.n294 163.367
R685 B.n294 B.n33 163.367
R686 B.n290 B.n33 163.367
R687 B.n290 B.n289 163.367
R688 B.n289 B.n288 163.367
R689 B.n288 B.n35 163.367
R690 B.n284 B.n35 163.367
R691 B.n284 B.n283 163.367
R692 B.n283 B.n282 163.367
R693 B.n282 B.n37 163.367
R694 B.n278 B.n37 163.367
R695 B.n278 B.n277 163.367
R696 B.n277 B.n276 163.367
R697 B.n276 B.n39 163.367
R698 B.n272 B.n39 163.367
R699 B.n272 B.n271 163.367
R700 B.n271 B.n270 163.367
R701 B.n270 B.n41 163.367
R702 B.n266 B.n41 163.367
R703 B.n266 B.n265 163.367
R704 B.n265 B.n264 163.367
R705 B.n264 B.n43 163.367
R706 B.n260 B.n43 163.367
R707 B.n260 B.n259 163.367
R708 B.n74 B.n73 59.5399
R709 B.n160 B.n81 59.5399
R710 B.n24 B.n23 59.5399
R711 B.n298 B.n31 59.5399
R712 B.n353 B.n352 33.2493
R713 B.n257 B.n44 33.2493
R714 B.n215 B.n214 33.2493
R715 B.n119 B.n94 33.2493
R716 B.n73 B.n72 19.9763
R717 B.n81 B.n80 19.9763
R718 B.n23 B.n22 19.9763
R719 B.n31 B.n30 19.9763
R720 B B.n375 18.0485
R721 B.n352 B.n351 10.6151
R722 B.n351 B.n10 10.6151
R723 B.n347 B.n10 10.6151
R724 B.n347 B.n346 10.6151
R725 B.n346 B.n345 10.6151
R726 B.n345 B.n12 10.6151
R727 B.n341 B.n12 10.6151
R728 B.n341 B.n340 10.6151
R729 B.n340 B.n339 10.6151
R730 B.n339 B.n14 10.6151
R731 B.n335 B.n14 10.6151
R732 B.n335 B.n334 10.6151
R733 B.n334 B.n333 10.6151
R734 B.n333 B.n16 10.6151
R735 B.n329 B.n16 10.6151
R736 B.n329 B.n328 10.6151
R737 B.n328 B.n327 10.6151
R738 B.n327 B.n18 10.6151
R739 B.n323 B.n18 10.6151
R740 B.n323 B.n322 10.6151
R741 B.n322 B.n321 10.6151
R742 B.n321 B.n20 10.6151
R743 B.n317 B.n20 10.6151
R744 B.n317 B.n316 10.6151
R745 B.n316 B.n315 10.6151
R746 B.n312 B.n311 10.6151
R747 B.n311 B.n310 10.6151
R748 B.n310 B.n26 10.6151
R749 B.n306 B.n26 10.6151
R750 B.n306 B.n305 10.6151
R751 B.n305 B.n304 10.6151
R752 B.n304 B.n28 10.6151
R753 B.n300 B.n28 10.6151
R754 B.n300 B.n299 10.6151
R755 B.n297 B.n32 10.6151
R756 B.n293 B.n32 10.6151
R757 B.n293 B.n292 10.6151
R758 B.n292 B.n291 10.6151
R759 B.n291 B.n34 10.6151
R760 B.n287 B.n34 10.6151
R761 B.n287 B.n286 10.6151
R762 B.n286 B.n285 10.6151
R763 B.n285 B.n36 10.6151
R764 B.n281 B.n36 10.6151
R765 B.n281 B.n280 10.6151
R766 B.n280 B.n279 10.6151
R767 B.n279 B.n38 10.6151
R768 B.n275 B.n38 10.6151
R769 B.n275 B.n274 10.6151
R770 B.n274 B.n273 10.6151
R771 B.n273 B.n40 10.6151
R772 B.n269 B.n40 10.6151
R773 B.n269 B.n268 10.6151
R774 B.n268 B.n267 10.6151
R775 B.n267 B.n42 10.6151
R776 B.n263 B.n42 10.6151
R777 B.n263 B.n262 10.6151
R778 B.n262 B.n261 10.6151
R779 B.n261 B.n44 10.6151
R780 B.n215 B.n58 10.6151
R781 B.n219 B.n58 10.6151
R782 B.n220 B.n219 10.6151
R783 B.n221 B.n220 10.6151
R784 B.n221 B.n56 10.6151
R785 B.n225 B.n56 10.6151
R786 B.n226 B.n225 10.6151
R787 B.n227 B.n226 10.6151
R788 B.n227 B.n54 10.6151
R789 B.n231 B.n54 10.6151
R790 B.n232 B.n231 10.6151
R791 B.n233 B.n232 10.6151
R792 B.n233 B.n52 10.6151
R793 B.n237 B.n52 10.6151
R794 B.n238 B.n237 10.6151
R795 B.n239 B.n238 10.6151
R796 B.n239 B.n50 10.6151
R797 B.n243 B.n50 10.6151
R798 B.n244 B.n243 10.6151
R799 B.n245 B.n244 10.6151
R800 B.n245 B.n48 10.6151
R801 B.n249 B.n48 10.6151
R802 B.n250 B.n249 10.6151
R803 B.n251 B.n250 10.6151
R804 B.n251 B.n46 10.6151
R805 B.n255 B.n46 10.6151
R806 B.n256 B.n255 10.6151
R807 B.n257 B.n256 10.6151
R808 B.n123 B.n94 10.6151
R809 B.n124 B.n123 10.6151
R810 B.n125 B.n124 10.6151
R811 B.n125 B.n92 10.6151
R812 B.n129 B.n92 10.6151
R813 B.n130 B.n129 10.6151
R814 B.n131 B.n130 10.6151
R815 B.n131 B.n90 10.6151
R816 B.n135 B.n90 10.6151
R817 B.n136 B.n135 10.6151
R818 B.n137 B.n136 10.6151
R819 B.n137 B.n88 10.6151
R820 B.n141 B.n88 10.6151
R821 B.n142 B.n141 10.6151
R822 B.n143 B.n142 10.6151
R823 B.n143 B.n86 10.6151
R824 B.n147 B.n86 10.6151
R825 B.n148 B.n147 10.6151
R826 B.n149 B.n148 10.6151
R827 B.n149 B.n84 10.6151
R828 B.n153 B.n84 10.6151
R829 B.n154 B.n153 10.6151
R830 B.n155 B.n154 10.6151
R831 B.n155 B.n82 10.6151
R832 B.n159 B.n82 10.6151
R833 B.n162 B.n161 10.6151
R834 B.n162 B.n78 10.6151
R835 B.n166 B.n78 10.6151
R836 B.n167 B.n166 10.6151
R837 B.n168 B.n167 10.6151
R838 B.n168 B.n76 10.6151
R839 B.n172 B.n76 10.6151
R840 B.n173 B.n172 10.6151
R841 B.n174 B.n173 10.6151
R842 B.n178 B.n177 10.6151
R843 B.n179 B.n178 10.6151
R844 B.n179 B.n70 10.6151
R845 B.n183 B.n70 10.6151
R846 B.n184 B.n183 10.6151
R847 B.n185 B.n184 10.6151
R848 B.n185 B.n68 10.6151
R849 B.n189 B.n68 10.6151
R850 B.n190 B.n189 10.6151
R851 B.n191 B.n190 10.6151
R852 B.n191 B.n66 10.6151
R853 B.n195 B.n66 10.6151
R854 B.n196 B.n195 10.6151
R855 B.n197 B.n196 10.6151
R856 B.n197 B.n64 10.6151
R857 B.n201 B.n64 10.6151
R858 B.n202 B.n201 10.6151
R859 B.n203 B.n202 10.6151
R860 B.n203 B.n62 10.6151
R861 B.n207 B.n62 10.6151
R862 B.n208 B.n207 10.6151
R863 B.n209 B.n208 10.6151
R864 B.n209 B.n60 10.6151
R865 B.n213 B.n60 10.6151
R866 B.n214 B.n213 10.6151
R867 B.n119 B.n118 10.6151
R868 B.n118 B.n117 10.6151
R869 B.n117 B.n96 10.6151
R870 B.n113 B.n96 10.6151
R871 B.n113 B.n112 10.6151
R872 B.n112 B.n111 10.6151
R873 B.n111 B.n98 10.6151
R874 B.n107 B.n98 10.6151
R875 B.n107 B.n106 10.6151
R876 B.n106 B.n105 10.6151
R877 B.n105 B.n100 10.6151
R878 B.n101 B.n100 10.6151
R879 B.n101 B.n0 10.6151
R880 B.n371 B.n1 10.6151
R881 B.n371 B.n370 10.6151
R882 B.n370 B.n369 10.6151
R883 B.n369 B.n4 10.6151
R884 B.n365 B.n4 10.6151
R885 B.n365 B.n364 10.6151
R886 B.n364 B.n363 10.6151
R887 B.n363 B.n6 10.6151
R888 B.n359 B.n6 10.6151
R889 B.n359 B.n358 10.6151
R890 B.n358 B.n357 10.6151
R891 B.n357 B.n8 10.6151
R892 B.n353 B.n8 10.6151
R893 B.n315 B.n24 8.74196
R894 B.n298 B.n297 8.74196
R895 B.n160 B.n159 8.74196
R896 B.n177 B.n74 8.74196
R897 B.n375 B.n0 2.81026
R898 B.n375 B.n1 2.81026
R899 B.n312 B.n24 1.87367
R900 B.n299 B.n298 1.87367
R901 B.n161 B.n160 1.87367
R902 B.n174 B.n74 1.87367
R903 VP.n0 VP.t0 484.404
R904 VP.n0 VP.t1 448.779
R905 VP VP.n0 0.0516364
R906 VDD1.n30 VDD1.n0 756.745
R907 VDD1.n65 VDD1.n35 756.745
R908 VDD1.n31 VDD1.n30 585
R909 VDD1.n29 VDD1.n28 585
R910 VDD1.n4 VDD1.n3 585
R911 VDD1.n23 VDD1.n22 585
R912 VDD1.n21 VDD1.n20 585
R913 VDD1.n8 VDD1.n7 585
R914 VDD1.n15 VDD1.n14 585
R915 VDD1.n13 VDD1.n12 585
R916 VDD1.n48 VDD1.n47 585
R917 VDD1.n50 VDD1.n49 585
R918 VDD1.n43 VDD1.n42 585
R919 VDD1.n56 VDD1.n55 585
R920 VDD1.n58 VDD1.n57 585
R921 VDD1.n39 VDD1.n38 585
R922 VDD1.n64 VDD1.n63 585
R923 VDD1.n66 VDD1.n65 585
R924 VDD1.n11 VDD1.t1 327.514
R925 VDD1.n46 VDD1.t0 327.514
R926 VDD1.n30 VDD1.n29 171.744
R927 VDD1.n29 VDD1.n3 171.744
R928 VDD1.n22 VDD1.n3 171.744
R929 VDD1.n22 VDD1.n21 171.744
R930 VDD1.n21 VDD1.n7 171.744
R931 VDD1.n14 VDD1.n7 171.744
R932 VDD1.n14 VDD1.n13 171.744
R933 VDD1.n49 VDD1.n48 171.744
R934 VDD1.n49 VDD1.n42 171.744
R935 VDD1.n56 VDD1.n42 171.744
R936 VDD1.n57 VDD1.n56 171.744
R937 VDD1.n57 VDD1.n38 171.744
R938 VDD1.n64 VDD1.n38 171.744
R939 VDD1.n65 VDD1.n64 171.744
R940 VDD1.n13 VDD1.t1 85.8723
R941 VDD1.n48 VDD1.t0 85.8723
R942 VDD1 VDD1.n69 80.654
R943 VDD1 VDD1.n34 48.9504
R944 VDD1.n47 VDD1.n46 16.3884
R945 VDD1.n12 VDD1.n11 16.3884
R946 VDD1.n15 VDD1.n10 12.8005
R947 VDD1.n50 VDD1.n45 12.8005
R948 VDD1.n16 VDD1.n8 12.0247
R949 VDD1.n51 VDD1.n43 12.0247
R950 VDD1.n20 VDD1.n19 11.249
R951 VDD1.n55 VDD1.n54 11.249
R952 VDD1.n23 VDD1.n6 10.4732
R953 VDD1.n58 VDD1.n41 10.4732
R954 VDD1.n24 VDD1.n4 9.69747
R955 VDD1.n59 VDD1.n39 9.69747
R956 VDD1.n34 VDD1.n33 9.45567
R957 VDD1.n69 VDD1.n68 9.45567
R958 VDD1.n33 VDD1.n32 9.3005
R959 VDD1.n2 VDD1.n1 9.3005
R960 VDD1.n27 VDD1.n26 9.3005
R961 VDD1.n25 VDD1.n24 9.3005
R962 VDD1.n6 VDD1.n5 9.3005
R963 VDD1.n19 VDD1.n18 9.3005
R964 VDD1.n17 VDD1.n16 9.3005
R965 VDD1.n10 VDD1.n9 9.3005
R966 VDD1.n37 VDD1.n36 9.3005
R967 VDD1.n62 VDD1.n61 9.3005
R968 VDD1.n60 VDD1.n59 9.3005
R969 VDD1.n41 VDD1.n40 9.3005
R970 VDD1.n54 VDD1.n53 9.3005
R971 VDD1.n52 VDD1.n51 9.3005
R972 VDD1.n45 VDD1.n44 9.3005
R973 VDD1.n68 VDD1.n67 9.3005
R974 VDD1.n28 VDD1.n27 8.92171
R975 VDD1.n63 VDD1.n62 8.92171
R976 VDD1.n31 VDD1.n2 8.14595
R977 VDD1.n66 VDD1.n37 8.14595
R978 VDD1.n32 VDD1.n0 7.3702
R979 VDD1.n67 VDD1.n35 7.3702
R980 VDD1.n34 VDD1.n0 6.59444
R981 VDD1.n69 VDD1.n35 6.59444
R982 VDD1.n32 VDD1.n31 5.81868
R983 VDD1.n67 VDD1.n66 5.81868
R984 VDD1.n28 VDD1.n2 5.04292
R985 VDD1.n63 VDD1.n37 5.04292
R986 VDD1.n27 VDD1.n4 4.26717
R987 VDD1.n62 VDD1.n39 4.26717
R988 VDD1.n11 VDD1.n9 3.71088
R989 VDD1.n46 VDD1.n44 3.71088
R990 VDD1.n24 VDD1.n23 3.49141
R991 VDD1.n59 VDD1.n58 3.49141
R992 VDD1.n20 VDD1.n6 2.71565
R993 VDD1.n55 VDD1.n41 2.71565
R994 VDD1.n19 VDD1.n8 1.93989
R995 VDD1.n54 VDD1.n43 1.93989
R996 VDD1.n16 VDD1.n15 1.16414
R997 VDD1.n51 VDD1.n50 1.16414
R998 VDD1.n12 VDD1.n10 0.388379
R999 VDD1.n47 VDD1.n45 0.388379
R1000 VDD1.n33 VDD1.n1 0.155672
R1001 VDD1.n26 VDD1.n1 0.155672
R1002 VDD1.n26 VDD1.n25 0.155672
R1003 VDD1.n25 VDD1.n5 0.155672
R1004 VDD1.n18 VDD1.n5 0.155672
R1005 VDD1.n18 VDD1.n17 0.155672
R1006 VDD1.n17 VDD1.n9 0.155672
R1007 VDD1.n52 VDD1.n44 0.155672
R1008 VDD1.n53 VDD1.n52 0.155672
R1009 VDD1.n53 VDD1.n40 0.155672
R1010 VDD1.n60 VDD1.n40 0.155672
R1011 VDD1.n61 VDD1.n60 0.155672
R1012 VDD1.n61 VDD1.n36 0.155672
R1013 VDD1.n68 VDD1.n36 0.155672
C0 VDD1 VN 0.148589f
C1 VTAIL VDD2 3.74157f
C2 VP VDD2 0.254194f
C3 w_n1382_n2314# VDD2 1.18627f
C4 B VDD2 1.04531f
C5 VTAIL VP 0.997339f
C6 VDD1 VDD2 0.460656f
C7 w_n1382_n2314# VTAIL 2.0376f
C8 VTAIL B 1.77161f
C9 VDD1 VTAIL 3.70478f
C10 VN VDD2 1.21566f
C11 w_n1382_n2314# VP 1.81969f
C12 B VP 0.93967f
C13 VDD1 VP 1.31875f
C14 w_n1382_n2314# B 5.27813f
C15 VTAIL VN 0.982953f
C16 w_n1382_n2314# VDD1 1.18162f
C17 VDD1 B 1.03081f
C18 VN VP 3.58214f
C19 w_n1382_n2314# VN 1.64775f
C20 VN B 0.664609f
C21 VDD2 VSUBS 0.554876f
C22 VDD1 VSUBS 2.055193f
C23 VTAIL VSUBS 0.471693f
C24 VN VSUBS 3.80289f
C25 VP VSUBS 0.857682f
C26 B VSUBS 2.047821f
C27 w_n1382_n2314# VSUBS 39.8182f
C28 VDD1.n0 VSUBS 0.017204f
C29 VDD1.n1 VSUBS 0.015537f
C30 VDD1.n2 VSUBS 0.008349f
C31 VDD1.n3 VSUBS 0.019733f
C32 VDD1.n4 VSUBS 0.00884f
C33 VDD1.n5 VSUBS 0.015537f
C34 VDD1.n6 VSUBS 0.008349f
C35 VDD1.n7 VSUBS 0.019733f
C36 VDD1.n8 VSUBS 0.00884f
C37 VDD1.n9 VSUBS 0.40679f
C38 VDD1.n10 VSUBS 0.008349f
C39 VDD1.t1 VSUBS 0.042206f
C40 VDD1.n11 VSUBS 0.071801f
C41 VDD1.n12 VSUBS 0.012551f
C42 VDD1.n13 VSUBS 0.0148f
C43 VDD1.n14 VSUBS 0.019733f
C44 VDD1.n15 VSUBS 0.00884f
C45 VDD1.n16 VSUBS 0.008349f
C46 VDD1.n17 VSUBS 0.015537f
C47 VDD1.n18 VSUBS 0.015537f
C48 VDD1.n19 VSUBS 0.008349f
C49 VDD1.n20 VSUBS 0.00884f
C50 VDD1.n21 VSUBS 0.019733f
C51 VDD1.n22 VSUBS 0.019733f
C52 VDD1.n23 VSUBS 0.00884f
C53 VDD1.n24 VSUBS 0.008349f
C54 VDD1.n25 VSUBS 0.015537f
C55 VDD1.n26 VSUBS 0.015537f
C56 VDD1.n27 VSUBS 0.008349f
C57 VDD1.n28 VSUBS 0.00884f
C58 VDD1.n29 VSUBS 0.019733f
C59 VDD1.n30 VSUBS 0.048224f
C60 VDD1.n31 VSUBS 0.00884f
C61 VDD1.n32 VSUBS 0.008349f
C62 VDD1.n33 VSUBS 0.0357f
C63 VDD1.n34 VSUBS 0.035245f
C64 VDD1.n35 VSUBS 0.017204f
C65 VDD1.n36 VSUBS 0.015537f
C66 VDD1.n37 VSUBS 0.008349f
C67 VDD1.n38 VSUBS 0.019733f
C68 VDD1.n39 VSUBS 0.00884f
C69 VDD1.n40 VSUBS 0.015537f
C70 VDD1.n41 VSUBS 0.008349f
C71 VDD1.n42 VSUBS 0.019733f
C72 VDD1.n43 VSUBS 0.00884f
C73 VDD1.n44 VSUBS 0.40679f
C74 VDD1.n45 VSUBS 0.008349f
C75 VDD1.t0 VSUBS 0.042206f
C76 VDD1.n46 VSUBS 0.071801f
C77 VDD1.n47 VSUBS 0.012551f
C78 VDD1.n48 VSUBS 0.0148f
C79 VDD1.n49 VSUBS 0.019733f
C80 VDD1.n50 VSUBS 0.00884f
C81 VDD1.n51 VSUBS 0.008349f
C82 VDD1.n52 VSUBS 0.015537f
C83 VDD1.n53 VSUBS 0.015537f
C84 VDD1.n54 VSUBS 0.008349f
C85 VDD1.n55 VSUBS 0.00884f
C86 VDD1.n56 VSUBS 0.019733f
C87 VDD1.n57 VSUBS 0.019733f
C88 VDD1.n58 VSUBS 0.00884f
C89 VDD1.n59 VSUBS 0.008349f
C90 VDD1.n60 VSUBS 0.015537f
C91 VDD1.n61 VSUBS 0.015537f
C92 VDD1.n62 VSUBS 0.008349f
C93 VDD1.n63 VSUBS 0.00884f
C94 VDD1.n64 VSUBS 0.019733f
C95 VDD1.n65 VSUBS 0.048224f
C96 VDD1.n66 VSUBS 0.00884f
C97 VDD1.n67 VSUBS 0.008349f
C98 VDD1.n68 VSUBS 0.0357f
C99 VDD1.n69 VSUBS 0.298448f
C100 VP.t0 VSUBS 0.645182f
C101 VP.t1 VSUBS 0.554941f
C102 VP.n0 VSUBS 2.38757f
C103 B.n0 VSUBS 0.004021f
C104 B.n1 VSUBS 0.004021f
C105 B.n2 VSUBS 0.006359f
C106 B.n3 VSUBS 0.006359f
C107 B.n4 VSUBS 0.006359f
C108 B.n5 VSUBS 0.006359f
C109 B.n6 VSUBS 0.006359f
C110 B.n7 VSUBS 0.006359f
C111 B.n8 VSUBS 0.006359f
C112 B.n9 VSUBS 0.01557f
C113 B.n10 VSUBS 0.006359f
C114 B.n11 VSUBS 0.006359f
C115 B.n12 VSUBS 0.006359f
C116 B.n13 VSUBS 0.006359f
C117 B.n14 VSUBS 0.006359f
C118 B.n15 VSUBS 0.006359f
C119 B.n16 VSUBS 0.006359f
C120 B.n17 VSUBS 0.006359f
C121 B.n18 VSUBS 0.006359f
C122 B.n19 VSUBS 0.006359f
C123 B.n20 VSUBS 0.006359f
C124 B.n21 VSUBS 0.006359f
C125 B.t8 VSUBS 0.09289f
C126 B.t7 VSUBS 0.102031f
C127 B.t6 VSUBS 0.183159f
C128 B.n22 VSUBS 0.172324f
C129 B.n23 VSUBS 0.146701f
C130 B.n24 VSUBS 0.014734f
C131 B.n25 VSUBS 0.006359f
C132 B.n26 VSUBS 0.006359f
C133 B.n27 VSUBS 0.006359f
C134 B.n28 VSUBS 0.006359f
C135 B.n29 VSUBS 0.006359f
C136 B.t11 VSUBS 0.092892f
C137 B.t10 VSUBS 0.102033f
C138 B.t9 VSUBS 0.183159f
C139 B.n30 VSUBS 0.172322f
C140 B.n31 VSUBS 0.146699f
C141 B.n32 VSUBS 0.006359f
C142 B.n33 VSUBS 0.006359f
C143 B.n34 VSUBS 0.006359f
C144 B.n35 VSUBS 0.006359f
C145 B.n36 VSUBS 0.006359f
C146 B.n37 VSUBS 0.006359f
C147 B.n38 VSUBS 0.006359f
C148 B.n39 VSUBS 0.006359f
C149 B.n40 VSUBS 0.006359f
C150 B.n41 VSUBS 0.006359f
C151 B.n42 VSUBS 0.006359f
C152 B.n43 VSUBS 0.006359f
C153 B.n44 VSUBS 0.014832f
C154 B.n45 VSUBS 0.006359f
C155 B.n46 VSUBS 0.006359f
C156 B.n47 VSUBS 0.006359f
C157 B.n48 VSUBS 0.006359f
C158 B.n49 VSUBS 0.006359f
C159 B.n50 VSUBS 0.006359f
C160 B.n51 VSUBS 0.006359f
C161 B.n52 VSUBS 0.006359f
C162 B.n53 VSUBS 0.006359f
C163 B.n54 VSUBS 0.006359f
C164 B.n55 VSUBS 0.006359f
C165 B.n56 VSUBS 0.006359f
C166 B.n57 VSUBS 0.006359f
C167 B.n58 VSUBS 0.006359f
C168 B.n59 VSUBS 0.01557f
C169 B.n60 VSUBS 0.006359f
C170 B.n61 VSUBS 0.006359f
C171 B.n62 VSUBS 0.006359f
C172 B.n63 VSUBS 0.006359f
C173 B.n64 VSUBS 0.006359f
C174 B.n65 VSUBS 0.006359f
C175 B.n66 VSUBS 0.006359f
C176 B.n67 VSUBS 0.006359f
C177 B.n68 VSUBS 0.006359f
C178 B.n69 VSUBS 0.006359f
C179 B.n70 VSUBS 0.006359f
C180 B.n71 VSUBS 0.006359f
C181 B.t4 VSUBS 0.092892f
C182 B.t5 VSUBS 0.102033f
C183 B.t3 VSUBS 0.183159f
C184 B.n72 VSUBS 0.172322f
C185 B.n73 VSUBS 0.146699f
C186 B.n74 VSUBS 0.014734f
C187 B.n75 VSUBS 0.006359f
C188 B.n76 VSUBS 0.006359f
C189 B.n77 VSUBS 0.006359f
C190 B.n78 VSUBS 0.006359f
C191 B.n79 VSUBS 0.006359f
C192 B.t1 VSUBS 0.09289f
C193 B.t2 VSUBS 0.102031f
C194 B.t0 VSUBS 0.183159f
C195 B.n80 VSUBS 0.172324f
C196 B.n81 VSUBS 0.146701f
C197 B.n82 VSUBS 0.006359f
C198 B.n83 VSUBS 0.006359f
C199 B.n84 VSUBS 0.006359f
C200 B.n85 VSUBS 0.006359f
C201 B.n86 VSUBS 0.006359f
C202 B.n87 VSUBS 0.006359f
C203 B.n88 VSUBS 0.006359f
C204 B.n89 VSUBS 0.006359f
C205 B.n90 VSUBS 0.006359f
C206 B.n91 VSUBS 0.006359f
C207 B.n92 VSUBS 0.006359f
C208 B.n93 VSUBS 0.006359f
C209 B.n94 VSUBS 0.01557f
C210 B.n95 VSUBS 0.006359f
C211 B.n96 VSUBS 0.006359f
C212 B.n97 VSUBS 0.006359f
C213 B.n98 VSUBS 0.006359f
C214 B.n99 VSUBS 0.006359f
C215 B.n100 VSUBS 0.006359f
C216 B.n101 VSUBS 0.006359f
C217 B.n102 VSUBS 0.006359f
C218 B.n103 VSUBS 0.006359f
C219 B.n104 VSUBS 0.006359f
C220 B.n105 VSUBS 0.006359f
C221 B.n106 VSUBS 0.006359f
C222 B.n107 VSUBS 0.006359f
C223 B.n108 VSUBS 0.006359f
C224 B.n109 VSUBS 0.006359f
C225 B.n110 VSUBS 0.006359f
C226 B.n111 VSUBS 0.006359f
C227 B.n112 VSUBS 0.006359f
C228 B.n113 VSUBS 0.006359f
C229 B.n114 VSUBS 0.006359f
C230 B.n115 VSUBS 0.006359f
C231 B.n116 VSUBS 0.006359f
C232 B.n117 VSUBS 0.006359f
C233 B.n118 VSUBS 0.006359f
C234 B.n119 VSUBS 0.014544f
C235 B.n120 VSUBS 0.014544f
C236 B.n121 VSUBS 0.01557f
C237 B.n122 VSUBS 0.006359f
C238 B.n123 VSUBS 0.006359f
C239 B.n124 VSUBS 0.006359f
C240 B.n125 VSUBS 0.006359f
C241 B.n126 VSUBS 0.006359f
C242 B.n127 VSUBS 0.006359f
C243 B.n128 VSUBS 0.006359f
C244 B.n129 VSUBS 0.006359f
C245 B.n130 VSUBS 0.006359f
C246 B.n131 VSUBS 0.006359f
C247 B.n132 VSUBS 0.006359f
C248 B.n133 VSUBS 0.006359f
C249 B.n134 VSUBS 0.006359f
C250 B.n135 VSUBS 0.006359f
C251 B.n136 VSUBS 0.006359f
C252 B.n137 VSUBS 0.006359f
C253 B.n138 VSUBS 0.006359f
C254 B.n139 VSUBS 0.006359f
C255 B.n140 VSUBS 0.006359f
C256 B.n141 VSUBS 0.006359f
C257 B.n142 VSUBS 0.006359f
C258 B.n143 VSUBS 0.006359f
C259 B.n144 VSUBS 0.006359f
C260 B.n145 VSUBS 0.006359f
C261 B.n146 VSUBS 0.006359f
C262 B.n147 VSUBS 0.006359f
C263 B.n148 VSUBS 0.006359f
C264 B.n149 VSUBS 0.006359f
C265 B.n150 VSUBS 0.006359f
C266 B.n151 VSUBS 0.006359f
C267 B.n152 VSUBS 0.006359f
C268 B.n153 VSUBS 0.006359f
C269 B.n154 VSUBS 0.006359f
C270 B.n155 VSUBS 0.006359f
C271 B.n156 VSUBS 0.006359f
C272 B.n157 VSUBS 0.006359f
C273 B.n158 VSUBS 0.006359f
C274 B.n159 VSUBS 0.005798f
C275 B.n160 VSUBS 0.014734f
C276 B.n161 VSUBS 0.003741f
C277 B.n162 VSUBS 0.006359f
C278 B.n163 VSUBS 0.006359f
C279 B.n164 VSUBS 0.006359f
C280 B.n165 VSUBS 0.006359f
C281 B.n166 VSUBS 0.006359f
C282 B.n167 VSUBS 0.006359f
C283 B.n168 VSUBS 0.006359f
C284 B.n169 VSUBS 0.006359f
C285 B.n170 VSUBS 0.006359f
C286 B.n171 VSUBS 0.006359f
C287 B.n172 VSUBS 0.006359f
C288 B.n173 VSUBS 0.006359f
C289 B.n174 VSUBS 0.003741f
C290 B.n175 VSUBS 0.006359f
C291 B.n176 VSUBS 0.006359f
C292 B.n177 VSUBS 0.005798f
C293 B.n178 VSUBS 0.006359f
C294 B.n179 VSUBS 0.006359f
C295 B.n180 VSUBS 0.006359f
C296 B.n181 VSUBS 0.006359f
C297 B.n182 VSUBS 0.006359f
C298 B.n183 VSUBS 0.006359f
C299 B.n184 VSUBS 0.006359f
C300 B.n185 VSUBS 0.006359f
C301 B.n186 VSUBS 0.006359f
C302 B.n187 VSUBS 0.006359f
C303 B.n188 VSUBS 0.006359f
C304 B.n189 VSUBS 0.006359f
C305 B.n190 VSUBS 0.006359f
C306 B.n191 VSUBS 0.006359f
C307 B.n192 VSUBS 0.006359f
C308 B.n193 VSUBS 0.006359f
C309 B.n194 VSUBS 0.006359f
C310 B.n195 VSUBS 0.006359f
C311 B.n196 VSUBS 0.006359f
C312 B.n197 VSUBS 0.006359f
C313 B.n198 VSUBS 0.006359f
C314 B.n199 VSUBS 0.006359f
C315 B.n200 VSUBS 0.006359f
C316 B.n201 VSUBS 0.006359f
C317 B.n202 VSUBS 0.006359f
C318 B.n203 VSUBS 0.006359f
C319 B.n204 VSUBS 0.006359f
C320 B.n205 VSUBS 0.006359f
C321 B.n206 VSUBS 0.006359f
C322 B.n207 VSUBS 0.006359f
C323 B.n208 VSUBS 0.006359f
C324 B.n209 VSUBS 0.006359f
C325 B.n210 VSUBS 0.006359f
C326 B.n211 VSUBS 0.006359f
C327 B.n212 VSUBS 0.006359f
C328 B.n213 VSUBS 0.006359f
C329 B.n214 VSUBS 0.01557f
C330 B.n215 VSUBS 0.014544f
C331 B.n216 VSUBS 0.014544f
C332 B.n217 VSUBS 0.006359f
C333 B.n218 VSUBS 0.006359f
C334 B.n219 VSUBS 0.006359f
C335 B.n220 VSUBS 0.006359f
C336 B.n221 VSUBS 0.006359f
C337 B.n222 VSUBS 0.006359f
C338 B.n223 VSUBS 0.006359f
C339 B.n224 VSUBS 0.006359f
C340 B.n225 VSUBS 0.006359f
C341 B.n226 VSUBS 0.006359f
C342 B.n227 VSUBS 0.006359f
C343 B.n228 VSUBS 0.006359f
C344 B.n229 VSUBS 0.006359f
C345 B.n230 VSUBS 0.006359f
C346 B.n231 VSUBS 0.006359f
C347 B.n232 VSUBS 0.006359f
C348 B.n233 VSUBS 0.006359f
C349 B.n234 VSUBS 0.006359f
C350 B.n235 VSUBS 0.006359f
C351 B.n236 VSUBS 0.006359f
C352 B.n237 VSUBS 0.006359f
C353 B.n238 VSUBS 0.006359f
C354 B.n239 VSUBS 0.006359f
C355 B.n240 VSUBS 0.006359f
C356 B.n241 VSUBS 0.006359f
C357 B.n242 VSUBS 0.006359f
C358 B.n243 VSUBS 0.006359f
C359 B.n244 VSUBS 0.006359f
C360 B.n245 VSUBS 0.006359f
C361 B.n246 VSUBS 0.006359f
C362 B.n247 VSUBS 0.006359f
C363 B.n248 VSUBS 0.006359f
C364 B.n249 VSUBS 0.006359f
C365 B.n250 VSUBS 0.006359f
C366 B.n251 VSUBS 0.006359f
C367 B.n252 VSUBS 0.006359f
C368 B.n253 VSUBS 0.006359f
C369 B.n254 VSUBS 0.006359f
C370 B.n255 VSUBS 0.006359f
C371 B.n256 VSUBS 0.006359f
C372 B.n257 VSUBS 0.015282f
C373 B.n258 VSUBS 0.014544f
C374 B.n259 VSUBS 0.01557f
C375 B.n260 VSUBS 0.006359f
C376 B.n261 VSUBS 0.006359f
C377 B.n262 VSUBS 0.006359f
C378 B.n263 VSUBS 0.006359f
C379 B.n264 VSUBS 0.006359f
C380 B.n265 VSUBS 0.006359f
C381 B.n266 VSUBS 0.006359f
C382 B.n267 VSUBS 0.006359f
C383 B.n268 VSUBS 0.006359f
C384 B.n269 VSUBS 0.006359f
C385 B.n270 VSUBS 0.006359f
C386 B.n271 VSUBS 0.006359f
C387 B.n272 VSUBS 0.006359f
C388 B.n273 VSUBS 0.006359f
C389 B.n274 VSUBS 0.006359f
C390 B.n275 VSUBS 0.006359f
C391 B.n276 VSUBS 0.006359f
C392 B.n277 VSUBS 0.006359f
C393 B.n278 VSUBS 0.006359f
C394 B.n279 VSUBS 0.006359f
C395 B.n280 VSUBS 0.006359f
C396 B.n281 VSUBS 0.006359f
C397 B.n282 VSUBS 0.006359f
C398 B.n283 VSUBS 0.006359f
C399 B.n284 VSUBS 0.006359f
C400 B.n285 VSUBS 0.006359f
C401 B.n286 VSUBS 0.006359f
C402 B.n287 VSUBS 0.006359f
C403 B.n288 VSUBS 0.006359f
C404 B.n289 VSUBS 0.006359f
C405 B.n290 VSUBS 0.006359f
C406 B.n291 VSUBS 0.006359f
C407 B.n292 VSUBS 0.006359f
C408 B.n293 VSUBS 0.006359f
C409 B.n294 VSUBS 0.006359f
C410 B.n295 VSUBS 0.006359f
C411 B.n296 VSUBS 0.006359f
C412 B.n297 VSUBS 0.005798f
C413 B.n298 VSUBS 0.014734f
C414 B.n299 VSUBS 0.003741f
C415 B.n300 VSUBS 0.006359f
C416 B.n301 VSUBS 0.006359f
C417 B.n302 VSUBS 0.006359f
C418 B.n303 VSUBS 0.006359f
C419 B.n304 VSUBS 0.006359f
C420 B.n305 VSUBS 0.006359f
C421 B.n306 VSUBS 0.006359f
C422 B.n307 VSUBS 0.006359f
C423 B.n308 VSUBS 0.006359f
C424 B.n309 VSUBS 0.006359f
C425 B.n310 VSUBS 0.006359f
C426 B.n311 VSUBS 0.006359f
C427 B.n312 VSUBS 0.003741f
C428 B.n313 VSUBS 0.006359f
C429 B.n314 VSUBS 0.006359f
C430 B.n315 VSUBS 0.005798f
C431 B.n316 VSUBS 0.006359f
C432 B.n317 VSUBS 0.006359f
C433 B.n318 VSUBS 0.006359f
C434 B.n319 VSUBS 0.006359f
C435 B.n320 VSUBS 0.006359f
C436 B.n321 VSUBS 0.006359f
C437 B.n322 VSUBS 0.006359f
C438 B.n323 VSUBS 0.006359f
C439 B.n324 VSUBS 0.006359f
C440 B.n325 VSUBS 0.006359f
C441 B.n326 VSUBS 0.006359f
C442 B.n327 VSUBS 0.006359f
C443 B.n328 VSUBS 0.006359f
C444 B.n329 VSUBS 0.006359f
C445 B.n330 VSUBS 0.006359f
C446 B.n331 VSUBS 0.006359f
C447 B.n332 VSUBS 0.006359f
C448 B.n333 VSUBS 0.006359f
C449 B.n334 VSUBS 0.006359f
C450 B.n335 VSUBS 0.006359f
C451 B.n336 VSUBS 0.006359f
C452 B.n337 VSUBS 0.006359f
C453 B.n338 VSUBS 0.006359f
C454 B.n339 VSUBS 0.006359f
C455 B.n340 VSUBS 0.006359f
C456 B.n341 VSUBS 0.006359f
C457 B.n342 VSUBS 0.006359f
C458 B.n343 VSUBS 0.006359f
C459 B.n344 VSUBS 0.006359f
C460 B.n345 VSUBS 0.006359f
C461 B.n346 VSUBS 0.006359f
C462 B.n347 VSUBS 0.006359f
C463 B.n348 VSUBS 0.006359f
C464 B.n349 VSUBS 0.006359f
C465 B.n350 VSUBS 0.006359f
C466 B.n351 VSUBS 0.006359f
C467 B.n352 VSUBS 0.01557f
C468 B.n353 VSUBS 0.014544f
C469 B.n354 VSUBS 0.014544f
C470 B.n355 VSUBS 0.006359f
C471 B.n356 VSUBS 0.006359f
C472 B.n357 VSUBS 0.006359f
C473 B.n358 VSUBS 0.006359f
C474 B.n359 VSUBS 0.006359f
C475 B.n360 VSUBS 0.006359f
C476 B.n361 VSUBS 0.006359f
C477 B.n362 VSUBS 0.006359f
C478 B.n363 VSUBS 0.006359f
C479 B.n364 VSUBS 0.006359f
C480 B.n365 VSUBS 0.006359f
C481 B.n366 VSUBS 0.006359f
C482 B.n367 VSUBS 0.006359f
C483 B.n368 VSUBS 0.006359f
C484 B.n369 VSUBS 0.006359f
C485 B.n370 VSUBS 0.006359f
C486 B.n371 VSUBS 0.006359f
C487 B.n372 VSUBS 0.006359f
C488 B.n373 VSUBS 0.006359f
C489 B.n374 VSUBS 0.006359f
C490 B.n375 VSUBS 0.0144f
C491 VDD2.n0 VSUBS 0.017475f
C492 VDD2.n1 VSUBS 0.015782f
C493 VDD2.n2 VSUBS 0.00848f
C494 VDD2.n3 VSUBS 0.020044f
C495 VDD2.n4 VSUBS 0.008979f
C496 VDD2.n5 VSUBS 0.015782f
C497 VDD2.n6 VSUBS 0.00848f
C498 VDD2.n7 VSUBS 0.020044f
C499 VDD2.n8 VSUBS 0.008979f
C500 VDD2.n9 VSUBS 0.413199f
C501 VDD2.n10 VSUBS 0.00848f
C502 VDD2.t1 VSUBS 0.042871f
C503 VDD2.n11 VSUBS 0.072933f
C504 VDD2.n12 VSUBS 0.012749f
C505 VDD2.n13 VSUBS 0.015033f
C506 VDD2.n14 VSUBS 0.020044f
C507 VDD2.n15 VSUBS 0.008979f
C508 VDD2.n16 VSUBS 0.00848f
C509 VDD2.n17 VSUBS 0.015782f
C510 VDD2.n18 VSUBS 0.015782f
C511 VDD2.n19 VSUBS 0.00848f
C512 VDD2.n20 VSUBS 0.008979f
C513 VDD2.n21 VSUBS 0.020044f
C514 VDD2.n22 VSUBS 0.020044f
C515 VDD2.n23 VSUBS 0.008979f
C516 VDD2.n24 VSUBS 0.00848f
C517 VDD2.n25 VSUBS 0.015782f
C518 VDD2.n26 VSUBS 0.015782f
C519 VDD2.n27 VSUBS 0.00848f
C520 VDD2.n28 VSUBS 0.008979f
C521 VDD2.n29 VSUBS 0.020044f
C522 VDD2.n30 VSUBS 0.048984f
C523 VDD2.n31 VSUBS 0.008979f
C524 VDD2.n32 VSUBS 0.00848f
C525 VDD2.n33 VSUBS 0.036263f
C526 VDD2.n34 VSUBS 0.284134f
C527 VDD2.n35 VSUBS 0.017475f
C528 VDD2.n36 VSUBS 0.015782f
C529 VDD2.n37 VSUBS 0.00848f
C530 VDD2.n38 VSUBS 0.020044f
C531 VDD2.n39 VSUBS 0.008979f
C532 VDD2.n40 VSUBS 0.015782f
C533 VDD2.n41 VSUBS 0.00848f
C534 VDD2.n42 VSUBS 0.020044f
C535 VDD2.n43 VSUBS 0.008979f
C536 VDD2.n44 VSUBS 0.413199f
C537 VDD2.n45 VSUBS 0.00848f
C538 VDD2.t0 VSUBS 0.042871f
C539 VDD2.n46 VSUBS 0.072933f
C540 VDD2.n47 VSUBS 0.012749f
C541 VDD2.n48 VSUBS 0.015033f
C542 VDD2.n49 VSUBS 0.020044f
C543 VDD2.n50 VSUBS 0.008979f
C544 VDD2.n51 VSUBS 0.00848f
C545 VDD2.n52 VSUBS 0.015782f
C546 VDD2.n53 VSUBS 0.015782f
C547 VDD2.n54 VSUBS 0.00848f
C548 VDD2.n55 VSUBS 0.008979f
C549 VDD2.n56 VSUBS 0.020044f
C550 VDD2.n57 VSUBS 0.020044f
C551 VDD2.n58 VSUBS 0.008979f
C552 VDD2.n59 VSUBS 0.00848f
C553 VDD2.n60 VSUBS 0.015782f
C554 VDD2.n61 VSUBS 0.015782f
C555 VDD2.n62 VSUBS 0.00848f
C556 VDD2.n63 VSUBS 0.008979f
C557 VDD2.n64 VSUBS 0.020044f
C558 VDD2.n65 VSUBS 0.048984f
C559 VDD2.n66 VSUBS 0.008979f
C560 VDD2.n67 VSUBS 0.00848f
C561 VDD2.n68 VSUBS 0.036263f
C562 VDD2.n69 VSUBS 0.035546f
C563 VDD2.n70 VSUBS 1.33274f
C564 VTAIL.n0 VSUBS 0.024639f
C565 VTAIL.n1 VSUBS 0.022251f
C566 VTAIL.n2 VSUBS 0.011957f
C567 VTAIL.n3 VSUBS 0.028261f
C568 VTAIL.n4 VSUBS 0.01266f
C569 VTAIL.n5 VSUBS 0.022251f
C570 VTAIL.n6 VSUBS 0.011957f
C571 VTAIL.n7 VSUBS 0.028261f
C572 VTAIL.n8 VSUBS 0.01266f
C573 VTAIL.n9 VSUBS 0.582577f
C574 VTAIL.n10 VSUBS 0.011957f
C575 VTAIL.t0 VSUBS 0.060444f
C576 VTAIL.n11 VSUBS 0.102829f
C577 VTAIL.n12 VSUBS 0.017975f
C578 VTAIL.n13 VSUBS 0.021196f
C579 VTAIL.n14 VSUBS 0.028261f
C580 VTAIL.n15 VSUBS 0.01266f
C581 VTAIL.n16 VSUBS 0.011957f
C582 VTAIL.n17 VSUBS 0.022251f
C583 VTAIL.n18 VSUBS 0.022251f
C584 VTAIL.n19 VSUBS 0.011957f
C585 VTAIL.n20 VSUBS 0.01266f
C586 VTAIL.n21 VSUBS 0.028261f
C587 VTAIL.n22 VSUBS 0.028261f
C588 VTAIL.n23 VSUBS 0.01266f
C589 VTAIL.n24 VSUBS 0.011957f
C590 VTAIL.n25 VSUBS 0.022251f
C591 VTAIL.n26 VSUBS 0.022251f
C592 VTAIL.n27 VSUBS 0.011957f
C593 VTAIL.n28 VSUBS 0.01266f
C594 VTAIL.n29 VSUBS 0.028261f
C595 VTAIL.n30 VSUBS 0.069064f
C596 VTAIL.n31 VSUBS 0.01266f
C597 VTAIL.n32 VSUBS 0.011957f
C598 VTAIL.n33 VSUBS 0.051127f
C599 VTAIL.n34 VSUBS 0.034751f
C600 VTAIL.n35 VSUBS 0.918143f
C601 VTAIL.n36 VSUBS 0.024639f
C602 VTAIL.n37 VSUBS 0.022251f
C603 VTAIL.n38 VSUBS 0.011957f
C604 VTAIL.n39 VSUBS 0.028261f
C605 VTAIL.n40 VSUBS 0.01266f
C606 VTAIL.n41 VSUBS 0.022251f
C607 VTAIL.n42 VSUBS 0.011957f
C608 VTAIL.n43 VSUBS 0.028261f
C609 VTAIL.n44 VSUBS 0.01266f
C610 VTAIL.n45 VSUBS 0.582577f
C611 VTAIL.n46 VSUBS 0.011957f
C612 VTAIL.t3 VSUBS 0.060444f
C613 VTAIL.n47 VSUBS 0.102829f
C614 VTAIL.n48 VSUBS 0.017975f
C615 VTAIL.n49 VSUBS 0.021196f
C616 VTAIL.n50 VSUBS 0.028261f
C617 VTAIL.n51 VSUBS 0.01266f
C618 VTAIL.n52 VSUBS 0.011957f
C619 VTAIL.n53 VSUBS 0.022251f
C620 VTAIL.n54 VSUBS 0.022251f
C621 VTAIL.n55 VSUBS 0.011957f
C622 VTAIL.n56 VSUBS 0.01266f
C623 VTAIL.n57 VSUBS 0.028261f
C624 VTAIL.n58 VSUBS 0.028261f
C625 VTAIL.n59 VSUBS 0.01266f
C626 VTAIL.n60 VSUBS 0.011957f
C627 VTAIL.n61 VSUBS 0.022251f
C628 VTAIL.n62 VSUBS 0.022251f
C629 VTAIL.n63 VSUBS 0.011957f
C630 VTAIL.n64 VSUBS 0.01266f
C631 VTAIL.n65 VSUBS 0.028261f
C632 VTAIL.n66 VSUBS 0.069064f
C633 VTAIL.n67 VSUBS 0.01266f
C634 VTAIL.n68 VSUBS 0.011957f
C635 VTAIL.n69 VSUBS 0.051127f
C636 VTAIL.n70 VSUBS 0.034751f
C637 VTAIL.n71 VSUBS 0.929887f
C638 VTAIL.n72 VSUBS 0.024639f
C639 VTAIL.n73 VSUBS 0.022251f
C640 VTAIL.n74 VSUBS 0.011957f
C641 VTAIL.n75 VSUBS 0.028261f
C642 VTAIL.n76 VSUBS 0.01266f
C643 VTAIL.n77 VSUBS 0.022251f
C644 VTAIL.n78 VSUBS 0.011957f
C645 VTAIL.n79 VSUBS 0.028261f
C646 VTAIL.n80 VSUBS 0.01266f
C647 VTAIL.n81 VSUBS 0.582577f
C648 VTAIL.n82 VSUBS 0.011957f
C649 VTAIL.t1 VSUBS 0.060444f
C650 VTAIL.n83 VSUBS 0.102829f
C651 VTAIL.n84 VSUBS 0.017975f
C652 VTAIL.n85 VSUBS 0.021196f
C653 VTAIL.n86 VSUBS 0.028261f
C654 VTAIL.n87 VSUBS 0.01266f
C655 VTAIL.n88 VSUBS 0.011957f
C656 VTAIL.n89 VSUBS 0.022251f
C657 VTAIL.n90 VSUBS 0.022251f
C658 VTAIL.n91 VSUBS 0.011957f
C659 VTAIL.n92 VSUBS 0.01266f
C660 VTAIL.n93 VSUBS 0.028261f
C661 VTAIL.n94 VSUBS 0.028261f
C662 VTAIL.n95 VSUBS 0.01266f
C663 VTAIL.n96 VSUBS 0.011957f
C664 VTAIL.n97 VSUBS 0.022251f
C665 VTAIL.n98 VSUBS 0.022251f
C666 VTAIL.n99 VSUBS 0.011957f
C667 VTAIL.n100 VSUBS 0.01266f
C668 VTAIL.n101 VSUBS 0.028261f
C669 VTAIL.n102 VSUBS 0.069064f
C670 VTAIL.n103 VSUBS 0.01266f
C671 VTAIL.n104 VSUBS 0.011957f
C672 VTAIL.n105 VSUBS 0.051127f
C673 VTAIL.n106 VSUBS 0.034751f
C674 VTAIL.n107 VSUBS 0.866225f
C675 VTAIL.n108 VSUBS 0.024639f
C676 VTAIL.n109 VSUBS 0.022251f
C677 VTAIL.n110 VSUBS 0.011957f
C678 VTAIL.n111 VSUBS 0.028261f
C679 VTAIL.n112 VSUBS 0.01266f
C680 VTAIL.n113 VSUBS 0.022251f
C681 VTAIL.n114 VSUBS 0.011957f
C682 VTAIL.n115 VSUBS 0.028261f
C683 VTAIL.n116 VSUBS 0.01266f
C684 VTAIL.n117 VSUBS 0.582577f
C685 VTAIL.n118 VSUBS 0.011957f
C686 VTAIL.t2 VSUBS 0.060444f
C687 VTAIL.n119 VSUBS 0.102829f
C688 VTAIL.n120 VSUBS 0.017975f
C689 VTAIL.n121 VSUBS 0.021196f
C690 VTAIL.n122 VSUBS 0.028261f
C691 VTAIL.n123 VSUBS 0.01266f
C692 VTAIL.n124 VSUBS 0.011957f
C693 VTAIL.n125 VSUBS 0.022251f
C694 VTAIL.n126 VSUBS 0.022251f
C695 VTAIL.n127 VSUBS 0.011957f
C696 VTAIL.n128 VSUBS 0.01266f
C697 VTAIL.n129 VSUBS 0.028261f
C698 VTAIL.n130 VSUBS 0.028261f
C699 VTAIL.n131 VSUBS 0.01266f
C700 VTAIL.n132 VSUBS 0.011957f
C701 VTAIL.n133 VSUBS 0.022251f
C702 VTAIL.n134 VSUBS 0.022251f
C703 VTAIL.n135 VSUBS 0.011957f
C704 VTAIL.n136 VSUBS 0.01266f
C705 VTAIL.n137 VSUBS 0.028261f
C706 VTAIL.n138 VSUBS 0.069064f
C707 VTAIL.n139 VSUBS 0.01266f
C708 VTAIL.n140 VSUBS 0.011957f
C709 VTAIL.n141 VSUBS 0.051127f
C710 VTAIL.n142 VSUBS 0.034751f
C711 VTAIL.n143 VSUBS 0.812452f
C712 VN.t0 VSUBS 0.547408f
C713 VN.t1 VSUBS 0.639001f
.ends

