* NGSPICE file created from diff_pair_sample_0491.ext - technology: sky130A

.subckt diff_pair_sample_0491 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t7 VN.t0 VDD2.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=5.9163 pd=31.12 as=2.50305 ps=15.5 w=15.17 l=3.16
X1 VTAIL.t1 VP.t0 VDD1.t3 B.t1 sky130_fd_pr__nfet_01v8 ad=5.9163 pd=31.12 as=2.50305 ps=15.5 w=15.17 l=3.16
X2 B.t17 B.t15 B.t16 B.t12 sky130_fd_pr__nfet_01v8 ad=5.9163 pd=31.12 as=0 ps=0 w=15.17 l=3.16
X3 B.t14 B.t11 B.t13 B.t12 sky130_fd_pr__nfet_01v8 ad=5.9163 pd=31.12 as=0 ps=0 w=15.17 l=3.16
X4 VTAIL.t2 VP.t1 VDD1.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=5.9163 pd=31.12 as=2.50305 ps=15.5 w=15.17 l=3.16
X5 VDD1.t1 VP.t2 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=2.50305 pd=15.5 as=5.9163 ps=31.12 w=15.17 l=3.16
X6 VDD2.t0 VN.t1 VTAIL.t6 B.t3 sky130_fd_pr__nfet_01v8 ad=2.50305 pd=15.5 as=5.9163 ps=31.12 w=15.17 l=3.16
X7 B.t10 B.t8 B.t9 B.t5 sky130_fd_pr__nfet_01v8 ad=5.9163 pd=31.12 as=0 ps=0 w=15.17 l=3.16
X8 VDD1.t0 VP.t3 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=2.50305 pd=15.5 as=5.9163 ps=31.12 w=15.17 l=3.16
X9 VDD2.t3 VN.t2 VTAIL.t5 B.t0 sky130_fd_pr__nfet_01v8 ad=2.50305 pd=15.5 as=5.9163 ps=31.12 w=15.17 l=3.16
X10 B.t7 B.t4 B.t6 B.t5 sky130_fd_pr__nfet_01v8 ad=5.9163 pd=31.12 as=0 ps=0 w=15.17 l=3.16
X11 VTAIL.t4 VN.t3 VDD2.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=5.9163 pd=31.12 as=2.50305 ps=15.5 w=15.17 l=3.16
R0 VN.n0 VN.t3 150.206
R1 VN.n1 VN.t1 150.206
R2 VN.n0 VN.t2 149.12
R3 VN.n1 VN.t0 149.12
R4 VN VN.n1 53.2417
R5 VN VN.n0 2.67727
R6 VDD2.n2 VDD2.n0 109.995
R7 VDD2.n2 VDD2.n1 64.1766
R8 VDD2.n1 VDD2.t2 1.30571
R9 VDD2.n1 VDD2.t0 1.30571
R10 VDD2.n0 VDD2.t1 1.30571
R11 VDD2.n0 VDD2.t3 1.30571
R12 VDD2 VDD2.n2 0.0586897
R13 VTAIL.n5 VTAIL.t1 48.8032
R14 VTAIL.n4 VTAIL.t6 48.8032
R15 VTAIL.n3 VTAIL.t7 48.8032
R16 VTAIL.n7 VTAIL.t5 48.803
R17 VTAIL.n0 VTAIL.t4 48.803
R18 VTAIL.n1 VTAIL.t3 48.803
R19 VTAIL.n2 VTAIL.t2 48.803
R20 VTAIL.n6 VTAIL.t0 48.803
R21 VTAIL.n7 VTAIL.n6 28.4531
R22 VTAIL.n3 VTAIL.n2 28.4531
R23 VTAIL.n4 VTAIL.n3 3.00912
R24 VTAIL.n6 VTAIL.n5 3.00912
R25 VTAIL.n2 VTAIL.n1 3.00912
R26 VTAIL VTAIL.n0 1.563
R27 VTAIL VTAIL.n7 1.44662
R28 VTAIL.n5 VTAIL.n4 0.470328
R29 VTAIL.n1 VTAIL.n0 0.470328
R30 B.n877 B.n876 585
R31 B.n878 B.n877 585
R32 B.n351 B.n129 585
R33 B.n350 B.n349 585
R34 B.n348 B.n347 585
R35 B.n346 B.n345 585
R36 B.n344 B.n343 585
R37 B.n342 B.n341 585
R38 B.n340 B.n339 585
R39 B.n338 B.n337 585
R40 B.n336 B.n335 585
R41 B.n334 B.n333 585
R42 B.n332 B.n331 585
R43 B.n330 B.n329 585
R44 B.n328 B.n327 585
R45 B.n326 B.n325 585
R46 B.n324 B.n323 585
R47 B.n322 B.n321 585
R48 B.n320 B.n319 585
R49 B.n318 B.n317 585
R50 B.n316 B.n315 585
R51 B.n314 B.n313 585
R52 B.n312 B.n311 585
R53 B.n310 B.n309 585
R54 B.n308 B.n307 585
R55 B.n306 B.n305 585
R56 B.n304 B.n303 585
R57 B.n302 B.n301 585
R58 B.n300 B.n299 585
R59 B.n298 B.n297 585
R60 B.n296 B.n295 585
R61 B.n294 B.n293 585
R62 B.n292 B.n291 585
R63 B.n290 B.n289 585
R64 B.n288 B.n287 585
R65 B.n286 B.n285 585
R66 B.n284 B.n283 585
R67 B.n282 B.n281 585
R68 B.n280 B.n279 585
R69 B.n278 B.n277 585
R70 B.n276 B.n275 585
R71 B.n274 B.n273 585
R72 B.n272 B.n271 585
R73 B.n270 B.n269 585
R74 B.n268 B.n267 585
R75 B.n266 B.n265 585
R76 B.n264 B.n263 585
R77 B.n262 B.n261 585
R78 B.n260 B.n259 585
R79 B.n258 B.n257 585
R80 B.n256 B.n255 585
R81 B.n254 B.n253 585
R82 B.n252 B.n251 585
R83 B.n250 B.n249 585
R84 B.n248 B.n247 585
R85 B.n246 B.n245 585
R86 B.n244 B.n243 585
R87 B.n242 B.n241 585
R88 B.n240 B.n239 585
R89 B.n238 B.n237 585
R90 B.n236 B.n235 585
R91 B.n233 B.n232 585
R92 B.n231 B.n230 585
R93 B.n229 B.n228 585
R94 B.n227 B.n226 585
R95 B.n225 B.n224 585
R96 B.n223 B.n222 585
R97 B.n221 B.n220 585
R98 B.n219 B.n218 585
R99 B.n217 B.n216 585
R100 B.n215 B.n214 585
R101 B.n213 B.n212 585
R102 B.n211 B.n210 585
R103 B.n209 B.n208 585
R104 B.n207 B.n206 585
R105 B.n205 B.n204 585
R106 B.n203 B.n202 585
R107 B.n201 B.n200 585
R108 B.n199 B.n198 585
R109 B.n197 B.n196 585
R110 B.n195 B.n194 585
R111 B.n193 B.n192 585
R112 B.n191 B.n190 585
R113 B.n189 B.n188 585
R114 B.n187 B.n186 585
R115 B.n185 B.n184 585
R116 B.n183 B.n182 585
R117 B.n181 B.n180 585
R118 B.n179 B.n178 585
R119 B.n177 B.n176 585
R120 B.n175 B.n174 585
R121 B.n173 B.n172 585
R122 B.n171 B.n170 585
R123 B.n169 B.n168 585
R124 B.n167 B.n166 585
R125 B.n165 B.n164 585
R126 B.n163 B.n162 585
R127 B.n161 B.n160 585
R128 B.n159 B.n158 585
R129 B.n157 B.n156 585
R130 B.n155 B.n154 585
R131 B.n153 B.n152 585
R132 B.n151 B.n150 585
R133 B.n149 B.n148 585
R134 B.n147 B.n146 585
R135 B.n145 B.n144 585
R136 B.n143 B.n142 585
R137 B.n141 B.n140 585
R138 B.n139 B.n138 585
R139 B.n137 B.n136 585
R140 B.n74 B.n73 585
R141 B.n881 B.n880 585
R142 B.n875 B.n130 585
R143 B.n130 B.n71 585
R144 B.n874 B.n70 585
R145 B.n885 B.n70 585
R146 B.n873 B.n69 585
R147 B.n886 B.n69 585
R148 B.n872 B.n68 585
R149 B.n887 B.n68 585
R150 B.n871 B.n870 585
R151 B.n870 B.n64 585
R152 B.n869 B.n63 585
R153 B.n893 B.n63 585
R154 B.n868 B.n62 585
R155 B.n894 B.n62 585
R156 B.n867 B.n61 585
R157 B.n895 B.n61 585
R158 B.n866 B.n865 585
R159 B.n865 B.n60 585
R160 B.n864 B.n56 585
R161 B.n901 B.n56 585
R162 B.n863 B.n55 585
R163 B.n902 B.n55 585
R164 B.n862 B.n54 585
R165 B.n903 B.n54 585
R166 B.n861 B.n860 585
R167 B.n860 B.n50 585
R168 B.n859 B.n49 585
R169 B.n909 B.n49 585
R170 B.n858 B.n48 585
R171 B.n910 B.n48 585
R172 B.n857 B.n47 585
R173 B.n911 B.n47 585
R174 B.n856 B.n855 585
R175 B.n855 B.n43 585
R176 B.n854 B.n42 585
R177 B.n917 B.n42 585
R178 B.n853 B.n41 585
R179 B.n918 B.n41 585
R180 B.n852 B.n40 585
R181 B.n919 B.n40 585
R182 B.n851 B.n850 585
R183 B.n850 B.n36 585
R184 B.n849 B.n35 585
R185 B.n925 B.n35 585
R186 B.n848 B.n34 585
R187 B.t0 B.n34 585
R188 B.n847 B.n33 585
R189 B.n926 B.n33 585
R190 B.n846 B.n845 585
R191 B.n845 B.n29 585
R192 B.n844 B.n28 585
R193 B.n932 B.n28 585
R194 B.n843 B.n27 585
R195 B.n933 B.n27 585
R196 B.n842 B.n26 585
R197 B.n934 B.n26 585
R198 B.n841 B.n840 585
R199 B.n840 B.n22 585
R200 B.n839 B.n21 585
R201 B.n940 B.n21 585
R202 B.n838 B.n20 585
R203 B.n941 B.n20 585
R204 B.n837 B.n19 585
R205 B.n942 B.n19 585
R206 B.n836 B.n835 585
R207 B.n835 B.n18 585
R208 B.n834 B.n14 585
R209 B.n948 B.n14 585
R210 B.n833 B.n13 585
R211 B.n949 B.n13 585
R212 B.n832 B.n12 585
R213 B.n950 B.n12 585
R214 B.n831 B.n830 585
R215 B.n830 B.n8 585
R216 B.n829 B.n7 585
R217 B.n956 B.n7 585
R218 B.n828 B.n6 585
R219 B.n957 B.n6 585
R220 B.n827 B.n5 585
R221 B.n958 B.n5 585
R222 B.n826 B.n825 585
R223 B.n825 B.n4 585
R224 B.n824 B.n352 585
R225 B.n824 B.n823 585
R226 B.n814 B.n353 585
R227 B.n354 B.n353 585
R228 B.n816 B.n815 585
R229 B.n817 B.n816 585
R230 B.n813 B.n359 585
R231 B.n359 B.n358 585
R232 B.n812 B.n811 585
R233 B.n811 B.n810 585
R234 B.n361 B.n360 585
R235 B.n803 B.n361 585
R236 B.n802 B.n801 585
R237 B.n804 B.n802 585
R238 B.n800 B.n366 585
R239 B.n366 B.n365 585
R240 B.n799 B.n798 585
R241 B.n798 B.n797 585
R242 B.n368 B.n367 585
R243 B.n369 B.n368 585
R244 B.n790 B.n789 585
R245 B.n791 B.n790 585
R246 B.n788 B.n374 585
R247 B.n374 B.n373 585
R248 B.n787 B.n786 585
R249 B.n786 B.n785 585
R250 B.n376 B.n375 585
R251 B.n377 B.n376 585
R252 B.n778 B.n777 585
R253 B.n779 B.n778 585
R254 B.n776 B.n381 585
R255 B.n381 B.t2 585
R256 B.n775 B.n774 585
R257 B.n774 B.n773 585
R258 B.n383 B.n382 585
R259 B.n384 B.n383 585
R260 B.n766 B.n765 585
R261 B.n767 B.n766 585
R262 B.n764 B.n389 585
R263 B.n389 B.n388 585
R264 B.n763 B.n762 585
R265 B.n762 B.n761 585
R266 B.n391 B.n390 585
R267 B.n392 B.n391 585
R268 B.n754 B.n753 585
R269 B.n755 B.n754 585
R270 B.n752 B.n397 585
R271 B.n397 B.n396 585
R272 B.n751 B.n750 585
R273 B.n750 B.n749 585
R274 B.n399 B.n398 585
R275 B.n400 B.n399 585
R276 B.n742 B.n741 585
R277 B.n743 B.n742 585
R278 B.n740 B.n405 585
R279 B.n405 B.n404 585
R280 B.n739 B.n738 585
R281 B.n738 B.n737 585
R282 B.n407 B.n406 585
R283 B.n730 B.n407 585
R284 B.n729 B.n728 585
R285 B.n731 B.n729 585
R286 B.n727 B.n412 585
R287 B.n412 B.n411 585
R288 B.n726 B.n725 585
R289 B.n725 B.n724 585
R290 B.n414 B.n413 585
R291 B.n415 B.n414 585
R292 B.n717 B.n716 585
R293 B.n718 B.n717 585
R294 B.n715 B.n420 585
R295 B.n420 B.n419 585
R296 B.n714 B.n713 585
R297 B.n713 B.n712 585
R298 B.n422 B.n421 585
R299 B.n423 B.n422 585
R300 B.n708 B.n707 585
R301 B.n426 B.n425 585
R302 B.n704 B.n703 585
R303 B.n705 B.n704 585
R304 B.n702 B.n481 585
R305 B.n701 B.n700 585
R306 B.n699 B.n698 585
R307 B.n697 B.n696 585
R308 B.n695 B.n694 585
R309 B.n693 B.n692 585
R310 B.n691 B.n690 585
R311 B.n689 B.n688 585
R312 B.n687 B.n686 585
R313 B.n685 B.n684 585
R314 B.n683 B.n682 585
R315 B.n681 B.n680 585
R316 B.n679 B.n678 585
R317 B.n677 B.n676 585
R318 B.n675 B.n674 585
R319 B.n673 B.n672 585
R320 B.n671 B.n670 585
R321 B.n669 B.n668 585
R322 B.n667 B.n666 585
R323 B.n665 B.n664 585
R324 B.n663 B.n662 585
R325 B.n661 B.n660 585
R326 B.n659 B.n658 585
R327 B.n657 B.n656 585
R328 B.n655 B.n654 585
R329 B.n653 B.n652 585
R330 B.n651 B.n650 585
R331 B.n649 B.n648 585
R332 B.n647 B.n646 585
R333 B.n645 B.n644 585
R334 B.n643 B.n642 585
R335 B.n641 B.n640 585
R336 B.n639 B.n638 585
R337 B.n637 B.n636 585
R338 B.n635 B.n634 585
R339 B.n633 B.n632 585
R340 B.n631 B.n630 585
R341 B.n629 B.n628 585
R342 B.n627 B.n626 585
R343 B.n625 B.n624 585
R344 B.n623 B.n622 585
R345 B.n621 B.n620 585
R346 B.n619 B.n618 585
R347 B.n617 B.n616 585
R348 B.n615 B.n614 585
R349 B.n613 B.n612 585
R350 B.n611 B.n610 585
R351 B.n609 B.n608 585
R352 B.n607 B.n606 585
R353 B.n605 B.n604 585
R354 B.n603 B.n602 585
R355 B.n601 B.n600 585
R356 B.n599 B.n598 585
R357 B.n597 B.n596 585
R358 B.n595 B.n594 585
R359 B.n593 B.n592 585
R360 B.n591 B.n590 585
R361 B.n588 B.n587 585
R362 B.n586 B.n585 585
R363 B.n584 B.n583 585
R364 B.n582 B.n581 585
R365 B.n580 B.n579 585
R366 B.n578 B.n577 585
R367 B.n576 B.n575 585
R368 B.n574 B.n573 585
R369 B.n572 B.n571 585
R370 B.n570 B.n569 585
R371 B.n568 B.n567 585
R372 B.n566 B.n565 585
R373 B.n564 B.n563 585
R374 B.n562 B.n561 585
R375 B.n560 B.n559 585
R376 B.n558 B.n557 585
R377 B.n556 B.n555 585
R378 B.n554 B.n553 585
R379 B.n552 B.n551 585
R380 B.n550 B.n549 585
R381 B.n548 B.n547 585
R382 B.n546 B.n545 585
R383 B.n544 B.n543 585
R384 B.n542 B.n541 585
R385 B.n540 B.n539 585
R386 B.n538 B.n537 585
R387 B.n536 B.n535 585
R388 B.n534 B.n533 585
R389 B.n532 B.n531 585
R390 B.n530 B.n529 585
R391 B.n528 B.n527 585
R392 B.n526 B.n525 585
R393 B.n524 B.n523 585
R394 B.n522 B.n521 585
R395 B.n520 B.n519 585
R396 B.n518 B.n517 585
R397 B.n516 B.n515 585
R398 B.n514 B.n513 585
R399 B.n512 B.n511 585
R400 B.n510 B.n509 585
R401 B.n508 B.n507 585
R402 B.n506 B.n505 585
R403 B.n504 B.n503 585
R404 B.n502 B.n501 585
R405 B.n500 B.n499 585
R406 B.n498 B.n497 585
R407 B.n496 B.n495 585
R408 B.n494 B.n493 585
R409 B.n492 B.n491 585
R410 B.n490 B.n489 585
R411 B.n488 B.n487 585
R412 B.n709 B.n424 585
R413 B.n424 B.n423 585
R414 B.n711 B.n710 585
R415 B.n712 B.n711 585
R416 B.n418 B.n417 585
R417 B.n419 B.n418 585
R418 B.n720 B.n719 585
R419 B.n719 B.n718 585
R420 B.n721 B.n416 585
R421 B.n416 B.n415 585
R422 B.n723 B.n722 585
R423 B.n724 B.n723 585
R424 B.n410 B.n409 585
R425 B.n411 B.n410 585
R426 B.n733 B.n732 585
R427 B.n732 B.n731 585
R428 B.n734 B.n408 585
R429 B.n730 B.n408 585
R430 B.n736 B.n735 585
R431 B.n737 B.n736 585
R432 B.n403 B.n402 585
R433 B.n404 B.n403 585
R434 B.n745 B.n744 585
R435 B.n744 B.n743 585
R436 B.n746 B.n401 585
R437 B.n401 B.n400 585
R438 B.n748 B.n747 585
R439 B.n749 B.n748 585
R440 B.n395 B.n394 585
R441 B.n396 B.n395 585
R442 B.n757 B.n756 585
R443 B.n756 B.n755 585
R444 B.n758 B.n393 585
R445 B.n393 B.n392 585
R446 B.n760 B.n759 585
R447 B.n761 B.n760 585
R448 B.n387 B.n386 585
R449 B.n388 B.n387 585
R450 B.n769 B.n768 585
R451 B.n768 B.n767 585
R452 B.n770 B.n385 585
R453 B.n385 B.n384 585
R454 B.n772 B.n771 585
R455 B.n773 B.n772 585
R456 B.n380 B.n379 585
R457 B.t2 B.n380 585
R458 B.n781 B.n780 585
R459 B.n780 B.n779 585
R460 B.n782 B.n378 585
R461 B.n378 B.n377 585
R462 B.n784 B.n783 585
R463 B.n785 B.n784 585
R464 B.n372 B.n371 585
R465 B.n373 B.n372 585
R466 B.n793 B.n792 585
R467 B.n792 B.n791 585
R468 B.n794 B.n370 585
R469 B.n370 B.n369 585
R470 B.n796 B.n795 585
R471 B.n797 B.n796 585
R472 B.n364 B.n363 585
R473 B.n365 B.n364 585
R474 B.n806 B.n805 585
R475 B.n805 B.n804 585
R476 B.n807 B.n362 585
R477 B.n803 B.n362 585
R478 B.n809 B.n808 585
R479 B.n810 B.n809 585
R480 B.n357 B.n356 585
R481 B.n358 B.n357 585
R482 B.n819 B.n818 585
R483 B.n818 B.n817 585
R484 B.n820 B.n355 585
R485 B.n355 B.n354 585
R486 B.n822 B.n821 585
R487 B.n823 B.n822 585
R488 B.n2 B.n0 585
R489 B.n4 B.n2 585
R490 B.n3 B.n1 585
R491 B.n957 B.n3 585
R492 B.n955 B.n954 585
R493 B.n956 B.n955 585
R494 B.n953 B.n9 585
R495 B.n9 B.n8 585
R496 B.n952 B.n951 585
R497 B.n951 B.n950 585
R498 B.n11 B.n10 585
R499 B.n949 B.n11 585
R500 B.n947 B.n946 585
R501 B.n948 B.n947 585
R502 B.n945 B.n15 585
R503 B.n18 B.n15 585
R504 B.n944 B.n943 585
R505 B.n943 B.n942 585
R506 B.n17 B.n16 585
R507 B.n941 B.n17 585
R508 B.n939 B.n938 585
R509 B.n940 B.n939 585
R510 B.n937 B.n23 585
R511 B.n23 B.n22 585
R512 B.n936 B.n935 585
R513 B.n935 B.n934 585
R514 B.n25 B.n24 585
R515 B.n933 B.n25 585
R516 B.n931 B.n930 585
R517 B.n932 B.n931 585
R518 B.n929 B.n30 585
R519 B.n30 B.n29 585
R520 B.n928 B.n927 585
R521 B.n927 B.n926 585
R522 B.n32 B.n31 585
R523 B.t0 B.n32 585
R524 B.n924 B.n923 585
R525 B.n925 B.n924 585
R526 B.n922 B.n37 585
R527 B.n37 B.n36 585
R528 B.n921 B.n920 585
R529 B.n920 B.n919 585
R530 B.n39 B.n38 585
R531 B.n918 B.n39 585
R532 B.n916 B.n915 585
R533 B.n917 B.n916 585
R534 B.n914 B.n44 585
R535 B.n44 B.n43 585
R536 B.n913 B.n912 585
R537 B.n912 B.n911 585
R538 B.n46 B.n45 585
R539 B.n910 B.n46 585
R540 B.n908 B.n907 585
R541 B.n909 B.n908 585
R542 B.n906 B.n51 585
R543 B.n51 B.n50 585
R544 B.n905 B.n904 585
R545 B.n904 B.n903 585
R546 B.n53 B.n52 585
R547 B.n902 B.n53 585
R548 B.n900 B.n899 585
R549 B.n901 B.n900 585
R550 B.n898 B.n57 585
R551 B.n60 B.n57 585
R552 B.n897 B.n896 585
R553 B.n896 B.n895 585
R554 B.n59 B.n58 585
R555 B.n894 B.n59 585
R556 B.n892 B.n891 585
R557 B.n893 B.n892 585
R558 B.n890 B.n65 585
R559 B.n65 B.n64 585
R560 B.n889 B.n888 585
R561 B.n888 B.n887 585
R562 B.n67 B.n66 585
R563 B.n886 B.n67 585
R564 B.n884 B.n883 585
R565 B.n885 B.n884 585
R566 B.n882 B.n72 585
R567 B.n72 B.n71 585
R568 B.n960 B.n959 585
R569 B.n959 B.n958 585
R570 B.n707 B.n424 521.33
R571 B.n880 B.n72 521.33
R572 B.n487 B.n422 521.33
R573 B.n877 B.n130 521.33
R574 B.n485 B.t11 324.455
R575 B.n482 B.t15 324.455
R576 B.n134 B.t8 324.455
R577 B.n131 B.t4 324.455
R578 B.n878 B.n128 256.663
R579 B.n878 B.n127 256.663
R580 B.n878 B.n126 256.663
R581 B.n878 B.n125 256.663
R582 B.n878 B.n124 256.663
R583 B.n878 B.n123 256.663
R584 B.n878 B.n122 256.663
R585 B.n878 B.n121 256.663
R586 B.n878 B.n120 256.663
R587 B.n878 B.n119 256.663
R588 B.n878 B.n118 256.663
R589 B.n878 B.n117 256.663
R590 B.n878 B.n116 256.663
R591 B.n878 B.n115 256.663
R592 B.n878 B.n114 256.663
R593 B.n878 B.n113 256.663
R594 B.n878 B.n112 256.663
R595 B.n878 B.n111 256.663
R596 B.n878 B.n110 256.663
R597 B.n878 B.n109 256.663
R598 B.n878 B.n108 256.663
R599 B.n878 B.n107 256.663
R600 B.n878 B.n106 256.663
R601 B.n878 B.n105 256.663
R602 B.n878 B.n104 256.663
R603 B.n878 B.n103 256.663
R604 B.n878 B.n102 256.663
R605 B.n878 B.n101 256.663
R606 B.n878 B.n100 256.663
R607 B.n878 B.n99 256.663
R608 B.n878 B.n98 256.663
R609 B.n878 B.n97 256.663
R610 B.n878 B.n96 256.663
R611 B.n878 B.n95 256.663
R612 B.n878 B.n94 256.663
R613 B.n878 B.n93 256.663
R614 B.n878 B.n92 256.663
R615 B.n878 B.n91 256.663
R616 B.n878 B.n90 256.663
R617 B.n878 B.n89 256.663
R618 B.n878 B.n88 256.663
R619 B.n878 B.n87 256.663
R620 B.n878 B.n86 256.663
R621 B.n878 B.n85 256.663
R622 B.n878 B.n84 256.663
R623 B.n878 B.n83 256.663
R624 B.n878 B.n82 256.663
R625 B.n878 B.n81 256.663
R626 B.n878 B.n80 256.663
R627 B.n878 B.n79 256.663
R628 B.n878 B.n78 256.663
R629 B.n878 B.n77 256.663
R630 B.n878 B.n76 256.663
R631 B.n878 B.n75 256.663
R632 B.n879 B.n878 256.663
R633 B.n706 B.n705 256.663
R634 B.n705 B.n427 256.663
R635 B.n705 B.n428 256.663
R636 B.n705 B.n429 256.663
R637 B.n705 B.n430 256.663
R638 B.n705 B.n431 256.663
R639 B.n705 B.n432 256.663
R640 B.n705 B.n433 256.663
R641 B.n705 B.n434 256.663
R642 B.n705 B.n435 256.663
R643 B.n705 B.n436 256.663
R644 B.n705 B.n437 256.663
R645 B.n705 B.n438 256.663
R646 B.n705 B.n439 256.663
R647 B.n705 B.n440 256.663
R648 B.n705 B.n441 256.663
R649 B.n705 B.n442 256.663
R650 B.n705 B.n443 256.663
R651 B.n705 B.n444 256.663
R652 B.n705 B.n445 256.663
R653 B.n705 B.n446 256.663
R654 B.n705 B.n447 256.663
R655 B.n705 B.n448 256.663
R656 B.n705 B.n449 256.663
R657 B.n705 B.n450 256.663
R658 B.n705 B.n451 256.663
R659 B.n705 B.n452 256.663
R660 B.n705 B.n453 256.663
R661 B.n705 B.n454 256.663
R662 B.n705 B.n455 256.663
R663 B.n705 B.n456 256.663
R664 B.n705 B.n457 256.663
R665 B.n705 B.n458 256.663
R666 B.n705 B.n459 256.663
R667 B.n705 B.n460 256.663
R668 B.n705 B.n461 256.663
R669 B.n705 B.n462 256.663
R670 B.n705 B.n463 256.663
R671 B.n705 B.n464 256.663
R672 B.n705 B.n465 256.663
R673 B.n705 B.n466 256.663
R674 B.n705 B.n467 256.663
R675 B.n705 B.n468 256.663
R676 B.n705 B.n469 256.663
R677 B.n705 B.n470 256.663
R678 B.n705 B.n471 256.663
R679 B.n705 B.n472 256.663
R680 B.n705 B.n473 256.663
R681 B.n705 B.n474 256.663
R682 B.n705 B.n475 256.663
R683 B.n705 B.n476 256.663
R684 B.n705 B.n477 256.663
R685 B.n705 B.n478 256.663
R686 B.n705 B.n479 256.663
R687 B.n705 B.n480 256.663
R688 B.n711 B.n424 163.367
R689 B.n711 B.n418 163.367
R690 B.n719 B.n418 163.367
R691 B.n719 B.n416 163.367
R692 B.n723 B.n416 163.367
R693 B.n723 B.n410 163.367
R694 B.n732 B.n410 163.367
R695 B.n732 B.n408 163.367
R696 B.n736 B.n408 163.367
R697 B.n736 B.n403 163.367
R698 B.n744 B.n403 163.367
R699 B.n744 B.n401 163.367
R700 B.n748 B.n401 163.367
R701 B.n748 B.n395 163.367
R702 B.n756 B.n395 163.367
R703 B.n756 B.n393 163.367
R704 B.n760 B.n393 163.367
R705 B.n760 B.n387 163.367
R706 B.n768 B.n387 163.367
R707 B.n768 B.n385 163.367
R708 B.n772 B.n385 163.367
R709 B.n772 B.n380 163.367
R710 B.n780 B.n380 163.367
R711 B.n780 B.n378 163.367
R712 B.n784 B.n378 163.367
R713 B.n784 B.n372 163.367
R714 B.n792 B.n372 163.367
R715 B.n792 B.n370 163.367
R716 B.n796 B.n370 163.367
R717 B.n796 B.n364 163.367
R718 B.n805 B.n364 163.367
R719 B.n805 B.n362 163.367
R720 B.n809 B.n362 163.367
R721 B.n809 B.n357 163.367
R722 B.n818 B.n357 163.367
R723 B.n818 B.n355 163.367
R724 B.n822 B.n355 163.367
R725 B.n822 B.n2 163.367
R726 B.n959 B.n2 163.367
R727 B.n959 B.n3 163.367
R728 B.n955 B.n3 163.367
R729 B.n955 B.n9 163.367
R730 B.n951 B.n9 163.367
R731 B.n951 B.n11 163.367
R732 B.n947 B.n11 163.367
R733 B.n947 B.n15 163.367
R734 B.n943 B.n15 163.367
R735 B.n943 B.n17 163.367
R736 B.n939 B.n17 163.367
R737 B.n939 B.n23 163.367
R738 B.n935 B.n23 163.367
R739 B.n935 B.n25 163.367
R740 B.n931 B.n25 163.367
R741 B.n931 B.n30 163.367
R742 B.n927 B.n30 163.367
R743 B.n927 B.n32 163.367
R744 B.n924 B.n32 163.367
R745 B.n924 B.n37 163.367
R746 B.n920 B.n37 163.367
R747 B.n920 B.n39 163.367
R748 B.n916 B.n39 163.367
R749 B.n916 B.n44 163.367
R750 B.n912 B.n44 163.367
R751 B.n912 B.n46 163.367
R752 B.n908 B.n46 163.367
R753 B.n908 B.n51 163.367
R754 B.n904 B.n51 163.367
R755 B.n904 B.n53 163.367
R756 B.n900 B.n53 163.367
R757 B.n900 B.n57 163.367
R758 B.n896 B.n57 163.367
R759 B.n896 B.n59 163.367
R760 B.n892 B.n59 163.367
R761 B.n892 B.n65 163.367
R762 B.n888 B.n65 163.367
R763 B.n888 B.n67 163.367
R764 B.n884 B.n67 163.367
R765 B.n884 B.n72 163.367
R766 B.n704 B.n426 163.367
R767 B.n704 B.n481 163.367
R768 B.n700 B.n699 163.367
R769 B.n696 B.n695 163.367
R770 B.n692 B.n691 163.367
R771 B.n688 B.n687 163.367
R772 B.n684 B.n683 163.367
R773 B.n680 B.n679 163.367
R774 B.n676 B.n675 163.367
R775 B.n672 B.n671 163.367
R776 B.n668 B.n667 163.367
R777 B.n664 B.n663 163.367
R778 B.n660 B.n659 163.367
R779 B.n656 B.n655 163.367
R780 B.n652 B.n651 163.367
R781 B.n648 B.n647 163.367
R782 B.n644 B.n643 163.367
R783 B.n640 B.n639 163.367
R784 B.n636 B.n635 163.367
R785 B.n632 B.n631 163.367
R786 B.n628 B.n627 163.367
R787 B.n624 B.n623 163.367
R788 B.n620 B.n619 163.367
R789 B.n616 B.n615 163.367
R790 B.n612 B.n611 163.367
R791 B.n608 B.n607 163.367
R792 B.n604 B.n603 163.367
R793 B.n600 B.n599 163.367
R794 B.n596 B.n595 163.367
R795 B.n592 B.n591 163.367
R796 B.n587 B.n586 163.367
R797 B.n583 B.n582 163.367
R798 B.n579 B.n578 163.367
R799 B.n575 B.n574 163.367
R800 B.n571 B.n570 163.367
R801 B.n567 B.n566 163.367
R802 B.n563 B.n562 163.367
R803 B.n559 B.n558 163.367
R804 B.n555 B.n554 163.367
R805 B.n551 B.n550 163.367
R806 B.n547 B.n546 163.367
R807 B.n543 B.n542 163.367
R808 B.n539 B.n538 163.367
R809 B.n535 B.n534 163.367
R810 B.n531 B.n530 163.367
R811 B.n527 B.n526 163.367
R812 B.n523 B.n522 163.367
R813 B.n519 B.n518 163.367
R814 B.n515 B.n514 163.367
R815 B.n511 B.n510 163.367
R816 B.n507 B.n506 163.367
R817 B.n503 B.n502 163.367
R818 B.n499 B.n498 163.367
R819 B.n495 B.n494 163.367
R820 B.n491 B.n490 163.367
R821 B.n713 B.n422 163.367
R822 B.n713 B.n420 163.367
R823 B.n717 B.n420 163.367
R824 B.n717 B.n414 163.367
R825 B.n725 B.n414 163.367
R826 B.n725 B.n412 163.367
R827 B.n729 B.n412 163.367
R828 B.n729 B.n407 163.367
R829 B.n738 B.n407 163.367
R830 B.n738 B.n405 163.367
R831 B.n742 B.n405 163.367
R832 B.n742 B.n399 163.367
R833 B.n750 B.n399 163.367
R834 B.n750 B.n397 163.367
R835 B.n754 B.n397 163.367
R836 B.n754 B.n391 163.367
R837 B.n762 B.n391 163.367
R838 B.n762 B.n389 163.367
R839 B.n766 B.n389 163.367
R840 B.n766 B.n383 163.367
R841 B.n774 B.n383 163.367
R842 B.n774 B.n381 163.367
R843 B.n778 B.n381 163.367
R844 B.n778 B.n376 163.367
R845 B.n786 B.n376 163.367
R846 B.n786 B.n374 163.367
R847 B.n790 B.n374 163.367
R848 B.n790 B.n368 163.367
R849 B.n798 B.n368 163.367
R850 B.n798 B.n366 163.367
R851 B.n802 B.n366 163.367
R852 B.n802 B.n361 163.367
R853 B.n811 B.n361 163.367
R854 B.n811 B.n359 163.367
R855 B.n816 B.n359 163.367
R856 B.n816 B.n353 163.367
R857 B.n824 B.n353 163.367
R858 B.n825 B.n824 163.367
R859 B.n825 B.n5 163.367
R860 B.n6 B.n5 163.367
R861 B.n7 B.n6 163.367
R862 B.n830 B.n7 163.367
R863 B.n830 B.n12 163.367
R864 B.n13 B.n12 163.367
R865 B.n14 B.n13 163.367
R866 B.n835 B.n14 163.367
R867 B.n835 B.n19 163.367
R868 B.n20 B.n19 163.367
R869 B.n21 B.n20 163.367
R870 B.n840 B.n21 163.367
R871 B.n840 B.n26 163.367
R872 B.n27 B.n26 163.367
R873 B.n28 B.n27 163.367
R874 B.n845 B.n28 163.367
R875 B.n845 B.n33 163.367
R876 B.n34 B.n33 163.367
R877 B.n35 B.n34 163.367
R878 B.n850 B.n35 163.367
R879 B.n850 B.n40 163.367
R880 B.n41 B.n40 163.367
R881 B.n42 B.n41 163.367
R882 B.n855 B.n42 163.367
R883 B.n855 B.n47 163.367
R884 B.n48 B.n47 163.367
R885 B.n49 B.n48 163.367
R886 B.n860 B.n49 163.367
R887 B.n860 B.n54 163.367
R888 B.n55 B.n54 163.367
R889 B.n56 B.n55 163.367
R890 B.n865 B.n56 163.367
R891 B.n865 B.n61 163.367
R892 B.n62 B.n61 163.367
R893 B.n63 B.n62 163.367
R894 B.n870 B.n63 163.367
R895 B.n870 B.n68 163.367
R896 B.n69 B.n68 163.367
R897 B.n70 B.n69 163.367
R898 B.n130 B.n70 163.367
R899 B.n136 B.n74 163.367
R900 B.n140 B.n139 163.367
R901 B.n144 B.n143 163.367
R902 B.n148 B.n147 163.367
R903 B.n152 B.n151 163.367
R904 B.n156 B.n155 163.367
R905 B.n160 B.n159 163.367
R906 B.n164 B.n163 163.367
R907 B.n168 B.n167 163.367
R908 B.n172 B.n171 163.367
R909 B.n176 B.n175 163.367
R910 B.n180 B.n179 163.367
R911 B.n184 B.n183 163.367
R912 B.n188 B.n187 163.367
R913 B.n192 B.n191 163.367
R914 B.n196 B.n195 163.367
R915 B.n200 B.n199 163.367
R916 B.n204 B.n203 163.367
R917 B.n208 B.n207 163.367
R918 B.n212 B.n211 163.367
R919 B.n216 B.n215 163.367
R920 B.n220 B.n219 163.367
R921 B.n224 B.n223 163.367
R922 B.n228 B.n227 163.367
R923 B.n232 B.n231 163.367
R924 B.n237 B.n236 163.367
R925 B.n241 B.n240 163.367
R926 B.n245 B.n244 163.367
R927 B.n249 B.n248 163.367
R928 B.n253 B.n252 163.367
R929 B.n257 B.n256 163.367
R930 B.n261 B.n260 163.367
R931 B.n265 B.n264 163.367
R932 B.n269 B.n268 163.367
R933 B.n273 B.n272 163.367
R934 B.n277 B.n276 163.367
R935 B.n281 B.n280 163.367
R936 B.n285 B.n284 163.367
R937 B.n289 B.n288 163.367
R938 B.n293 B.n292 163.367
R939 B.n297 B.n296 163.367
R940 B.n301 B.n300 163.367
R941 B.n305 B.n304 163.367
R942 B.n309 B.n308 163.367
R943 B.n313 B.n312 163.367
R944 B.n317 B.n316 163.367
R945 B.n321 B.n320 163.367
R946 B.n325 B.n324 163.367
R947 B.n329 B.n328 163.367
R948 B.n333 B.n332 163.367
R949 B.n337 B.n336 163.367
R950 B.n341 B.n340 163.367
R951 B.n345 B.n344 163.367
R952 B.n349 B.n348 163.367
R953 B.n877 B.n129 163.367
R954 B.n485 B.t14 139.208
R955 B.n131 B.t6 139.208
R956 B.n482 B.t17 139.188
R957 B.n134 B.t9 139.188
R958 B.n707 B.n706 71.676
R959 B.n481 B.n427 71.676
R960 B.n699 B.n428 71.676
R961 B.n695 B.n429 71.676
R962 B.n691 B.n430 71.676
R963 B.n687 B.n431 71.676
R964 B.n683 B.n432 71.676
R965 B.n679 B.n433 71.676
R966 B.n675 B.n434 71.676
R967 B.n671 B.n435 71.676
R968 B.n667 B.n436 71.676
R969 B.n663 B.n437 71.676
R970 B.n659 B.n438 71.676
R971 B.n655 B.n439 71.676
R972 B.n651 B.n440 71.676
R973 B.n647 B.n441 71.676
R974 B.n643 B.n442 71.676
R975 B.n639 B.n443 71.676
R976 B.n635 B.n444 71.676
R977 B.n631 B.n445 71.676
R978 B.n627 B.n446 71.676
R979 B.n623 B.n447 71.676
R980 B.n619 B.n448 71.676
R981 B.n615 B.n449 71.676
R982 B.n611 B.n450 71.676
R983 B.n607 B.n451 71.676
R984 B.n603 B.n452 71.676
R985 B.n599 B.n453 71.676
R986 B.n595 B.n454 71.676
R987 B.n591 B.n455 71.676
R988 B.n586 B.n456 71.676
R989 B.n582 B.n457 71.676
R990 B.n578 B.n458 71.676
R991 B.n574 B.n459 71.676
R992 B.n570 B.n460 71.676
R993 B.n566 B.n461 71.676
R994 B.n562 B.n462 71.676
R995 B.n558 B.n463 71.676
R996 B.n554 B.n464 71.676
R997 B.n550 B.n465 71.676
R998 B.n546 B.n466 71.676
R999 B.n542 B.n467 71.676
R1000 B.n538 B.n468 71.676
R1001 B.n534 B.n469 71.676
R1002 B.n530 B.n470 71.676
R1003 B.n526 B.n471 71.676
R1004 B.n522 B.n472 71.676
R1005 B.n518 B.n473 71.676
R1006 B.n514 B.n474 71.676
R1007 B.n510 B.n475 71.676
R1008 B.n506 B.n476 71.676
R1009 B.n502 B.n477 71.676
R1010 B.n498 B.n478 71.676
R1011 B.n494 B.n479 71.676
R1012 B.n490 B.n480 71.676
R1013 B.n880 B.n879 71.676
R1014 B.n136 B.n75 71.676
R1015 B.n140 B.n76 71.676
R1016 B.n144 B.n77 71.676
R1017 B.n148 B.n78 71.676
R1018 B.n152 B.n79 71.676
R1019 B.n156 B.n80 71.676
R1020 B.n160 B.n81 71.676
R1021 B.n164 B.n82 71.676
R1022 B.n168 B.n83 71.676
R1023 B.n172 B.n84 71.676
R1024 B.n176 B.n85 71.676
R1025 B.n180 B.n86 71.676
R1026 B.n184 B.n87 71.676
R1027 B.n188 B.n88 71.676
R1028 B.n192 B.n89 71.676
R1029 B.n196 B.n90 71.676
R1030 B.n200 B.n91 71.676
R1031 B.n204 B.n92 71.676
R1032 B.n208 B.n93 71.676
R1033 B.n212 B.n94 71.676
R1034 B.n216 B.n95 71.676
R1035 B.n220 B.n96 71.676
R1036 B.n224 B.n97 71.676
R1037 B.n228 B.n98 71.676
R1038 B.n232 B.n99 71.676
R1039 B.n237 B.n100 71.676
R1040 B.n241 B.n101 71.676
R1041 B.n245 B.n102 71.676
R1042 B.n249 B.n103 71.676
R1043 B.n253 B.n104 71.676
R1044 B.n257 B.n105 71.676
R1045 B.n261 B.n106 71.676
R1046 B.n265 B.n107 71.676
R1047 B.n269 B.n108 71.676
R1048 B.n273 B.n109 71.676
R1049 B.n277 B.n110 71.676
R1050 B.n281 B.n111 71.676
R1051 B.n285 B.n112 71.676
R1052 B.n289 B.n113 71.676
R1053 B.n293 B.n114 71.676
R1054 B.n297 B.n115 71.676
R1055 B.n301 B.n116 71.676
R1056 B.n305 B.n117 71.676
R1057 B.n309 B.n118 71.676
R1058 B.n313 B.n119 71.676
R1059 B.n317 B.n120 71.676
R1060 B.n321 B.n121 71.676
R1061 B.n325 B.n122 71.676
R1062 B.n329 B.n123 71.676
R1063 B.n333 B.n124 71.676
R1064 B.n337 B.n125 71.676
R1065 B.n341 B.n126 71.676
R1066 B.n345 B.n127 71.676
R1067 B.n349 B.n128 71.676
R1068 B.n129 B.n128 71.676
R1069 B.n348 B.n127 71.676
R1070 B.n344 B.n126 71.676
R1071 B.n340 B.n125 71.676
R1072 B.n336 B.n124 71.676
R1073 B.n332 B.n123 71.676
R1074 B.n328 B.n122 71.676
R1075 B.n324 B.n121 71.676
R1076 B.n320 B.n120 71.676
R1077 B.n316 B.n119 71.676
R1078 B.n312 B.n118 71.676
R1079 B.n308 B.n117 71.676
R1080 B.n304 B.n116 71.676
R1081 B.n300 B.n115 71.676
R1082 B.n296 B.n114 71.676
R1083 B.n292 B.n113 71.676
R1084 B.n288 B.n112 71.676
R1085 B.n284 B.n111 71.676
R1086 B.n280 B.n110 71.676
R1087 B.n276 B.n109 71.676
R1088 B.n272 B.n108 71.676
R1089 B.n268 B.n107 71.676
R1090 B.n264 B.n106 71.676
R1091 B.n260 B.n105 71.676
R1092 B.n256 B.n104 71.676
R1093 B.n252 B.n103 71.676
R1094 B.n248 B.n102 71.676
R1095 B.n244 B.n101 71.676
R1096 B.n240 B.n100 71.676
R1097 B.n236 B.n99 71.676
R1098 B.n231 B.n98 71.676
R1099 B.n227 B.n97 71.676
R1100 B.n223 B.n96 71.676
R1101 B.n219 B.n95 71.676
R1102 B.n215 B.n94 71.676
R1103 B.n211 B.n93 71.676
R1104 B.n207 B.n92 71.676
R1105 B.n203 B.n91 71.676
R1106 B.n199 B.n90 71.676
R1107 B.n195 B.n89 71.676
R1108 B.n191 B.n88 71.676
R1109 B.n187 B.n87 71.676
R1110 B.n183 B.n86 71.676
R1111 B.n179 B.n85 71.676
R1112 B.n175 B.n84 71.676
R1113 B.n171 B.n83 71.676
R1114 B.n167 B.n82 71.676
R1115 B.n163 B.n81 71.676
R1116 B.n159 B.n80 71.676
R1117 B.n155 B.n79 71.676
R1118 B.n151 B.n78 71.676
R1119 B.n147 B.n77 71.676
R1120 B.n143 B.n76 71.676
R1121 B.n139 B.n75 71.676
R1122 B.n879 B.n74 71.676
R1123 B.n706 B.n426 71.676
R1124 B.n700 B.n427 71.676
R1125 B.n696 B.n428 71.676
R1126 B.n692 B.n429 71.676
R1127 B.n688 B.n430 71.676
R1128 B.n684 B.n431 71.676
R1129 B.n680 B.n432 71.676
R1130 B.n676 B.n433 71.676
R1131 B.n672 B.n434 71.676
R1132 B.n668 B.n435 71.676
R1133 B.n664 B.n436 71.676
R1134 B.n660 B.n437 71.676
R1135 B.n656 B.n438 71.676
R1136 B.n652 B.n439 71.676
R1137 B.n648 B.n440 71.676
R1138 B.n644 B.n441 71.676
R1139 B.n640 B.n442 71.676
R1140 B.n636 B.n443 71.676
R1141 B.n632 B.n444 71.676
R1142 B.n628 B.n445 71.676
R1143 B.n624 B.n446 71.676
R1144 B.n620 B.n447 71.676
R1145 B.n616 B.n448 71.676
R1146 B.n612 B.n449 71.676
R1147 B.n608 B.n450 71.676
R1148 B.n604 B.n451 71.676
R1149 B.n600 B.n452 71.676
R1150 B.n596 B.n453 71.676
R1151 B.n592 B.n454 71.676
R1152 B.n587 B.n455 71.676
R1153 B.n583 B.n456 71.676
R1154 B.n579 B.n457 71.676
R1155 B.n575 B.n458 71.676
R1156 B.n571 B.n459 71.676
R1157 B.n567 B.n460 71.676
R1158 B.n563 B.n461 71.676
R1159 B.n559 B.n462 71.676
R1160 B.n555 B.n463 71.676
R1161 B.n551 B.n464 71.676
R1162 B.n547 B.n465 71.676
R1163 B.n543 B.n466 71.676
R1164 B.n539 B.n467 71.676
R1165 B.n535 B.n468 71.676
R1166 B.n531 B.n469 71.676
R1167 B.n527 B.n470 71.676
R1168 B.n523 B.n471 71.676
R1169 B.n519 B.n472 71.676
R1170 B.n515 B.n473 71.676
R1171 B.n511 B.n474 71.676
R1172 B.n507 B.n475 71.676
R1173 B.n503 B.n476 71.676
R1174 B.n499 B.n477 71.676
R1175 B.n495 B.n478 71.676
R1176 B.n491 B.n479 71.676
R1177 B.n487 B.n480 71.676
R1178 B.n486 B.t13 71.5223
R1179 B.n132 B.t7 71.5223
R1180 B.n483 B.t16 71.5026
R1181 B.n135 B.t10 71.5026
R1182 B.n486 B.n485 67.6854
R1183 B.n483 B.n482 67.6854
R1184 B.n135 B.n134 67.6854
R1185 B.n132 B.n131 67.6854
R1186 B.n705 B.n423 62.9499
R1187 B.n878 B.n71 62.9499
R1188 B.n589 B.n486 59.5399
R1189 B.n484 B.n483 59.5399
R1190 B.n234 B.n135 59.5399
R1191 B.n133 B.n132 59.5399
R1192 B.n712 B.n423 36.5865
R1193 B.n712 B.n419 36.5865
R1194 B.n718 B.n419 36.5865
R1195 B.n718 B.n415 36.5865
R1196 B.n724 B.n415 36.5865
R1197 B.n724 B.n411 36.5865
R1198 B.n731 B.n411 36.5865
R1199 B.n731 B.n730 36.5865
R1200 B.n737 B.n404 36.5865
R1201 B.n743 B.n404 36.5865
R1202 B.n743 B.n400 36.5865
R1203 B.n749 B.n400 36.5865
R1204 B.n749 B.n396 36.5865
R1205 B.n755 B.n396 36.5865
R1206 B.n755 B.n392 36.5865
R1207 B.n761 B.n392 36.5865
R1208 B.n761 B.n388 36.5865
R1209 B.n767 B.n388 36.5865
R1210 B.n767 B.n384 36.5865
R1211 B.n773 B.n384 36.5865
R1212 B.n773 B.t2 36.5865
R1213 B.n779 B.t2 36.5865
R1214 B.n779 B.n377 36.5865
R1215 B.n785 B.n377 36.5865
R1216 B.n785 B.n373 36.5865
R1217 B.n791 B.n373 36.5865
R1218 B.n791 B.n369 36.5865
R1219 B.n797 B.n369 36.5865
R1220 B.n797 B.n365 36.5865
R1221 B.n804 B.n365 36.5865
R1222 B.n804 B.n803 36.5865
R1223 B.n810 B.n358 36.5865
R1224 B.n817 B.n358 36.5865
R1225 B.n817 B.n354 36.5865
R1226 B.n823 B.n354 36.5865
R1227 B.n823 B.n4 36.5865
R1228 B.n958 B.n4 36.5865
R1229 B.n958 B.n957 36.5865
R1230 B.n957 B.n956 36.5865
R1231 B.n956 B.n8 36.5865
R1232 B.n950 B.n8 36.5865
R1233 B.n950 B.n949 36.5865
R1234 B.n949 B.n948 36.5865
R1235 B.n942 B.n18 36.5865
R1236 B.n942 B.n941 36.5865
R1237 B.n941 B.n940 36.5865
R1238 B.n940 B.n22 36.5865
R1239 B.n934 B.n22 36.5865
R1240 B.n934 B.n933 36.5865
R1241 B.n933 B.n932 36.5865
R1242 B.n932 B.n29 36.5865
R1243 B.n926 B.n29 36.5865
R1244 B.n926 B.t0 36.5865
R1245 B.t0 B.n925 36.5865
R1246 B.n925 B.n36 36.5865
R1247 B.n919 B.n36 36.5865
R1248 B.n919 B.n918 36.5865
R1249 B.n918 B.n917 36.5865
R1250 B.n917 B.n43 36.5865
R1251 B.n911 B.n43 36.5865
R1252 B.n911 B.n910 36.5865
R1253 B.n910 B.n909 36.5865
R1254 B.n909 B.n50 36.5865
R1255 B.n903 B.n50 36.5865
R1256 B.n903 B.n902 36.5865
R1257 B.n902 B.n901 36.5865
R1258 B.n895 B.n60 36.5865
R1259 B.n895 B.n894 36.5865
R1260 B.n894 B.n893 36.5865
R1261 B.n893 B.n64 36.5865
R1262 B.n887 B.n64 36.5865
R1263 B.n887 B.n886 36.5865
R1264 B.n886 B.n885 36.5865
R1265 B.n885 B.n71 36.5865
R1266 B.n882 B.n881 33.8737
R1267 B.n876 B.n875 33.8737
R1268 B.n488 B.n421 33.8737
R1269 B.n709 B.n708 33.8737
R1270 B.n810 B.t3 26.9019
R1271 B.n948 B.t1 26.9019
R1272 B.n730 B.t12 19.3695
R1273 B.n60 B.t5 19.3695
R1274 B B.n960 18.0485
R1275 B.n737 B.t12 17.2174
R1276 B.n901 B.t5 17.2174
R1277 B.n881 B.n73 10.6151
R1278 B.n137 B.n73 10.6151
R1279 B.n138 B.n137 10.6151
R1280 B.n141 B.n138 10.6151
R1281 B.n142 B.n141 10.6151
R1282 B.n145 B.n142 10.6151
R1283 B.n146 B.n145 10.6151
R1284 B.n149 B.n146 10.6151
R1285 B.n150 B.n149 10.6151
R1286 B.n153 B.n150 10.6151
R1287 B.n154 B.n153 10.6151
R1288 B.n157 B.n154 10.6151
R1289 B.n158 B.n157 10.6151
R1290 B.n161 B.n158 10.6151
R1291 B.n162 B.n161 10.6151
R1292 B.n165 B.n162 10.6151
R1293 B.n166 B.n165 10.6151
R1294 B.n169 B.n166 10.6151
R1295 B.n170 B.n169 10.6151
R1296 B.n173 B.n170 10.6151
R1297 B.n174 B.n173 10.6151
R1298 B.n177 B.n174 10.6151
R1299 B.n178 B.n177 10.6151
R1300 B.n181 B.n178 10.6151
R1301 B.n182 B.n181 10.6151
R1302 B.n185 B.n182 10.6151
R1303 B.n186 B.n185 10.6151
R1304 B.n189 B.n186 10.6151
R1305 B.n190 B.n189 10.6151
R1306 B.n193 B.n190 10.6151
R1307 B.n194 B.n193 10.6151
R1308 B.n197 B.n194 10.6151
R1309 B.n198 B.n197 10.6151
R1310 B.n201 B.n198 10.6151
R1311 B.n202 B.n201 10.6151
R1312 B.n205 B.n202 10.6151
R1313 B.n206 B.n205 10.6151
R1314 B.n209 B.n206 10.6151
R1315 B.n210 B.n209 10.6151
R1316 B.n213 B.n210 10.6151
R1317 B.n214 B.n213 10.6151
R1318 B.n217 B.n214 10.6151
R1319 B.n218 B.n217 10.6151
R1320 B.n221 B.n218 10.6151
R1321 B.n222 B.n221 10.6151
R1322 B.n225 B.n222 10.6151
R1323 B.n226 B.n225 10.6151
R1324 B.n229 B.n226 10.6151
R1325 B.n230 B.n229 10.6151
R1326 B.n233 B.n230 10.6151
R1327 B.n238 B.n235 10.6151
R1328 B.n239 B.n238 10.6151
R1329 B.n242 B.n239 10.6151
R1330 B.n243 B.n242 10.6151
R1331 B.n246 B.n243 10.6151
R1332 B.n247 B.n246 10.6151
R1333 B.n250 B.n247 10.6151
R1334 B.n251 B.n250 10.6151
R1335 B.n255 B.n254 10.6151
R1336 B.n258 B.n255 10.6151
R1337 B.n259 B.n258 10.6151
R1338 B.n262 B.n259 10.6151
R1339 B.n263 B.n262 10.6151
R1340 B.n266 B.n263 10.6151
R1341 B.n267 B.n266 10.6151
R1342 B.n270 B.n267 10.6151
R1343 B.n271 B.n270 10.6151
R1344 B.n274 B.n271 10.6151
R1345 B.n275 B.n274 10.6151
R1346 B.n278 B.n275 10.6151
R1347 B.n279 B.n278 10.6151
R1348 B.n282 B.n279 10.6151
R1349 B.n283 B.n282 10.6151
R1350 B.n286 B.n283 10.6151
R1351 B.n287 B.n286 10.6151
R1352 B.n290 B.n287 10.6151
R1353 B.n291 B.n290 10.6151
R1354 B.n294 B.n291 10.6151
R1355 B.n295 B.n294 10.6151
R1356 B.n298 B.n295 10.6151
R1357 B.n299 B.n298 10.6151
R1358 B.n302 B.n299 10.6151
R1359 B.n303 B.n302 10.6151
R1360 B.n306 B.n303 10.6151
R1361 B.n307 B.n306 10.6151
R1362 B.n310 B.n307 10.6151
R1363 B.n311 B.n310 10.6151
R1364 B.n314 B.n311 10.6151
R1365 B.n315 B.n314 10.6151
R1366 B.n318 B.n315 10.6151
R1367 B.n319 B.n318 10.6151
R1368 B.n322 B.n319 10.6151
R1369 B.n323 B.n322 10.6151
R1370 B.n326 B.n323 10.6151
R1371 B.n327 B.n326 10.6151
R1372 B.n330 B.n327 10.6151
R1373 B.n331 B.n330 10.6151
R1374 B.n334 B.n331 10.6151
R1375 B.n335 B.n334 10.6151
R1376 B.n338 B.n335 10.6151
R1377 B.n339 B.n338 10.6151
R1378 B.n342 B.n339 10.6151
R1379 B.n343 B.n342 10.6151
R1380 B.n346 B.n343 10.6151
R1381 B.n347 B.n346 10.6151
R1382 B.n350 B.n347 10.6151
R1383 B.n351 B.n350 10.6151
R1384 B.n876 B.n351 10.6151
R1385 B.n714 B.n421 10.6151
R1386 B.n715 B.n714 10.6151
R1387 B.n716 B.n715 10.6151
R1388 B.n716 B.n413 10.6151
R1389 B.n726 B.n413 10.6151
R1390 B.n727 B.n726 10.6151
R1391 B.n728 B.n727 10.6151
R1392 B.n728 B.n406 10.6151
R1393 B.n739 B.n406 10.6151
R1394 B.n740 B.n739 10.6151
R1395 B.n741 B.n740 10.6151
R1396 B.n741 B.n398 10.6151
R1397 B.n751 B.n398 10.6151
R1398 B.n752 B.n751 10.6151
R1399 B.n753 B.n752 10.6151
R1400 B.n753 B.n390 10.6151
R1401 B.n763 B.n390 10.6151
R1402 B.n764 B.n763 10.6151
R1403 B.n765 B.n764 10.6151
R1404 B.n765 B.n382 10.6151
R1405 B.n775 B.n382 10.6151
R1406 B.n776 B.n775 10.6151
R1407 B.n777 B.n776 10.6151
R1408 B.n777 B.n375 10.6151
R1409 B.n787 B.n375 10.6151
R1410 B.n788 B.n787 10.6151
R1411 B.n789 B.n788 10.6151
R1412 B.n789 B.n367 10.6151
R1413 B.n799 B.n367 10.6151
R1414 B.n800 B.n799 10.6151
R1415 B.n801 B.n800 10.6151
R1416 B.n801 B.n360 10.6151
R1417 B.n812 B.n360 10.6151
R1418 B.n813 B.n812 10.6151
R1419 B.n815 B.n813 10.6151
R1420 B.n815 B.n814 10.6151
R1421 B.n814 B.n352 10.6151
R1422 B.n826 B.n352 10.6151
R1423 B.n827 B.n826 10.6151
R1424 B.n828 B.n827 10.6151
R1425 B.n829 B.n828 10.6151
R1426 B.n831 B.n829 10.6151
R1427 B.n832 B.n831 10.6151
R1428 B.n833 B.n832 10.6151
R1429 B.n834 B.n833 10.6151
R1430 B.n836 B.n834 10.6151
R1431 B.n837 B.n836 10.6151
R1432 B.n838 B.n837 10.6151
R1433 B.n839 B.n838 10.6151
R1434 B.n841 B.n839 10.6151
R1435 B.n842 B.n841 10.6151
R1436 B.n843 B.n842 10.6151
R1437 B.n844 B.n843 10.6151
R1438 B.n846 B.n844 10.6151
R1439 B.n847 B.n846 10.6151
R1440 B.n848 B.n847 10.6151
R1441 B.n849 B.n848 10.6151
R1442 B.n851 B.n849 10.6151
R1443 B.n852 B.n851 10.6151
R1444 B.n853 B.n852 10.6151
R1445 B.n854 B.n853 10.6151
R1446 B.n856 B.n854 10.6151
R1447 B.n857 B.n856 10.6151
R1448 B.n858 B.n857 10.6151
R1449 B.n859 B.n858 10.6151
R1450 B.n861 B.n859 10.6151
R1451 B.n862 B.n861 10.6151
R1452 B.n863 B.n862 10.6151
R1453 B.n864 B.n863 10.6151
R1454 B.n866 B.n864 10.6151
R1455 B.n867 B.n866 10.6151
R1456 B.n868 B.n867 10.6151
R1457 B.n869 B.n868 10.6151
R1458 B.n871 B.n869 10.6151
R1459 B.n872 B.n871 10.6151
R1460 B.n873 B.n872 10.6151
R1461 B.n874 B.n873 10.6151
R1462 B.n875 B.n874 10.6151
R1463 B.n708 B.n425 10.6151
R1464 B.n703 B.n425 10.6151
R1465 B.n703 B.n702 10.6151
R1466 B.n702 B.n701 10.6151
R1467 B.n701 B.n698 10.6151
R1468 B.n698 B.n697 10.6151
R1469 B.n697 B.n694 10.6151
R1470 B.n694 B.n693 10.6151
R1471 B.n693 B.n690 10.6151
R1472 B.n690 B.n689 10.6151
R1473 B.n689 B.n686 10.6151
R1474 B.n686 B.n685 10.6151
R1475 B.n685 B.n682 10.6151
R1476 B.n682 B.n681 10.6151
R1477 B.n681 B.n678 10.6151
R1478 B.n678 B.n677 10.6151
R1479 B.n677 B.n674 10.6151
R1480 B.n674 B.n673 10.6151
R1481 B.n673 B.n670 10.6151
R1482 B.n670 B.n669 10.6151
R1483 B.n669 B.n666 10.6151
R1484 B.n666 B.n665 10.6151
R1485 B.n665 B.n662 10.6151
R1486 B.n662 B.n661 10.6151
R1487 B.n661 B.n658 10.6151
R1488 B.n658 B.n657 10.6151
R1489 B.n657 B.n654 10.6151
R1490 B.n654 B.n653 10.6151
R1491 B.n653 B.n650 10.6151
R1492 B.n650 B.n649 10.6151
R1493 B.n649 B.n646 10.6151
R1494 B.n646 B.n645 10.6151
R1495 B.n645 B.n642 10.6151
R1496 B.n642 B.n641 10.6151
R1497 B.n641 B.n638 10.6151
R1498 B.n638 B.n637 10.6151
R1499 B.n637 B.n634 10.6151
R1500 B.n634 B.n633 10.6151
R1501 B.n633 B.n630 10.6151
R1502 B.n630 B.n629 10.6151
R1503 B.n629 B.n626 10.6151
R1504 B.n626 B.n625 10.6151
R1505 B.n625 B.n622 10.6151
R1506 B.n622 B.n621 10.6151
R1507 B.n621 B.n618 10.6151
R1508 B.n618 B.n617 10.6151
R1509 B.n617 B.n614 10.6151
R1510 B.n614 B.n613 10.6151
R1511 B.n613 B.n610 10.6151
R1512 B.n610 B.n609 10.6151
R1513 B.n606 B.n605 10.6151
R1514 B.n605 B.n602 10.6151
R1515 B.n602 B.n601 10.6151
R1516 B.n601 B.n598 10.6151
R1517 B.n598 B.n597 10.6151
R1518 B.n597 B.n594 10.6151
R1519 B.n594 B.n593 10.6151
R1520 B.n593 B.n590 10.6151
R1521 B.n588 B.n585 10.6151
R1522 B.n585 B.n584 10.6151
R1523 B.n584 B.n581 10.6151
R1524 B.n581 B.n580 10.6151
R1525 B.n580 B.n577 10.6151
R1526 B.n577 B.n576 10.6151
R1527 B.n576 B.n573 10.6151
R1528 B.n573 B.n572 10.6151
R1529 B.n572 B.n569 10.6151
R1530 B.n569 B.n568 10.6151
R1531 B.n568 B.n565 10.6151
R1532 B.n565 B.n564 10.6151
R1533 B.n564 B.n561 10.6151
R1534 B.n561 B.n560 10.6151
R1535 B.n560 B.n557 10.6151
R1536 B.n557 B.n556 10.6151
R1537 B.n556 B.n553 10.6151
R1538 B.n553 B.n552 10.6151
R1539 B.n552 B.n549 10.6151
R1540 B.n549 B.n548 10.6151
R1541 B.n548 B.n545 10.6151
R1542 B.n545 B.n544 10.6151
R1543 B.n544 B.n541 10.6151
R1544 B.n541 B.n540 10.6151
R1545 B.n540 B.n537 10.6151
R1546 B.n537 B.n536 10.6151
R1547 B.n536 B.n533 10.6151
R1548 B.n533 B.n532 10.6151
R1549 B.n532 B.n529 10.6151
R1550 B.n529 B.n528 10.6151
R1551 B.n528 B.n525 10.6151
R1552 B.n525 B.n524 10.6151
R1553 B.n524 B.n521 10.6151
R1554 B.n521 B.n520 10.6151
R1555 B.n520 B.n517 10.6151
R1556 B.n517 B.n516 10.6151
R1557 B.n516 B.n513 10.6151
R1558 B.n513 B.n512 10.6151
R1559 B.n512 B.n509 10.6151
R1560 B.n509 B.n508 10.6151
R1561 B.n508 B.n505 10.6151
R1562 B.n505 B.n504 10.6151
R1563 B.n504 B.n501 10.6151
R1564 B.n501 B.n500 10.6151
R1565 B.n500 B.n497 10.6151
R1566 B.n497 B.n496 10.6151
R1567 B.n496 B.n493 10.6151
R1568 B.n493 B.n492 10.6151
R1569 B.n492 B.n489 10.6151
R1570 B.n489 B.n488 10.6151
R1571 B.n710 B.n709 10.6151
R1572 B.n710 B.n417 10.6151
R1573 B.n720 B.n417 10.6151
R1574 B.n721 B.n720 10.6151
R1575 B.n722 B.n721 10.6151
R1576 B.n722 B.n409 10.6151
R1577 B.n733 B.n409 10.6151
R1578 B.n734 B.n733 10.6151
R1579 B.n735 B.n734 10.6151
R1580 B.n735 B.n402 10.6151
R1581 B.n745 B.n402 10.6151
R1582 B.n746 B.n745 10.6151
R1583 B.n747 B.n746 10.6151
R1584 B.n747 B.n394 10.6151
R1585 B.n757 B.n394 10.6151
R1586 B.n758 B.n757 10.6151
R1587 B.n759 B.n758 10.6151
R1588 B.n759 B.n386 10.6151
R1589 B.n769 B.n386 10.6151
R1590 B.n770 B.n769 10.6151
R1591 B.n771 B.n770 10.6151
R1592 B.n771 B.n379 10.6151
R1593 B.n781 B.n379 10.6151
R1594 B.n782 B.n781 10.6151
R1595 B.n783 B.n782 10.6151
R1596 B.n783 B.n371 10.6151
R1597 B.n793 B.n371 10.6151
R1598 B.n794 B.n793 10.6151
R1599 B.n795 B.n794 10.6151
R1600 B.n795 B.n363 10.6151
R1601 B.n806 B.n363 10.6151
R1602 B.n807 B.n806 10.6151
R1603 B.n808 B.n807 10.6151
R1604 B.n808 B.n356 10.6151
R1605 B.n819 B.n356 10.6151
R1606 B.n820 B.n819 10.6151
R1607 B.n821 B.n820 10.6151
R1608 B.n821 B.n0 10.6151
R1609 B.n954 B.n1 10.6151
R1610 B.n954 B.n953 10.6151
R1611 B.n953 B.n952 10.6151
R1612 B.n952 B.n10 10.6151
R1613 B.n946 B.n10 10.6151
R1614 B.n946 B.n945 10.6151
R1615 B.n945 B.n944 10.6151
R1616 B.n944 B.n16 10.6151
R1617 B.n938 B.n16 10.6151
R1618 B.n938 B.n937 10.6151
R1619 B.n937 B.n936 10.6151
R1620 B.n936 B.n24 10.6151
R1621 B.n930 B.n24 10.6151
R1622 B.n930 B.n929 10.6151
R1623 B.n929 B.n928 10.6151
R1624 B.n928 B.n31 10.6151
R1625 B.n923 B.n31 10.6151
R1626 B.n923 B.n922 10.6151
R1627 B.n922 B.n921 10.6151
R1628 B.n921 B.n38 10.6151
R1629 B.n915 B.n38 10.6151
R1630 B.n915 B.n914 10.6151
R1631 B.n914 B.n913 10.6151
R1632 B.n913 B.n45 10.6151
R1633 B.n907 B.n45 10.6151
R1634 B.n907 B.n906 10.6151
R1635 B.n906 B.n905 10.6151
R1636 B.n905 B.n52 10.6151
R1637 B.n899 B.n52 10.6151
R1638 B.n899 B.n898 10.6151
R1639 B.n898 B.n897 10.6151
R1640 B.n897 B.n58 10.6151
R1641 B.n891 B.n58 10.6151
R1642 B.n891 B.n890 10.6151
R1643 B.n890 B.n889 10.6151
R1644 B.n889 B.n66 10.6151
R1645 B.n883 B.n66 10.6151
R1646 B.n883 B.n882 10.6151
R1647 B.n803 B.t3 9.68502
R1648 B.n18 B.t1 9.68502
R1649 B.n235 B.n234 6.5566
R1650 B.n251 B.n133 6.5566
R1651 B.n606 B.n484 6.5566
R1652 B.n590 B.n589 6.5566
R1653 B.n234 B.n233 4.05904
R1654 B.n254 B.n133 4.05904
R1655 B.n609 B.n484 4.05904
R1656 B.n589 B.n588 4.05904
R1657 B.n960 B.n0 2.81026
R1658 B.n960 B.n1 2.81026
R1659 VP.n17 VP.n16 161.3
R1660 VP.n15 VP.n1 161.3
R1661 VP.n14 VP.n13 161.3
R1662 VP.n12 VP.n2 161.3
R1663 VP.n11 VP.n10 161.3
R1664 VP.n9 VP.n3 161.3
R1665 VP.n8 VP.n7 161.3
R1666 VP.n5 VP.t0 150.206
R1667 VP.n5 VP.t3 149.12
R1668 VP.n4 VP.t1 115.695
R1669 VP.n0 VP.t2 115.695
R1670 VP.n6 VP.n4 78.0786
R1671 VP.n18 VP.n0 78.0786
R1672 VP.n6 VP.n5 53.0763
R1673 VP.n10 VP.n2 40.4934
R1674 VP.n14 VP.n2 40.4934
R1675 VP.n9 VP.n8 24.4675
R1676 VP.n10 VP.n9 24.4675
R1677 VP.n15 VP.n14 24.4675
R1678 VP.n16 VP.n15 24.4675
R1679 VP.n8 VP.n4 11.9893
R1680 VP.n16 VP.n0 11.9893
R1681 VP.n7 VP.n6 0.354971
R1682 VP.n18 VP.n17 0.354971
R1683 VP VP.n18 0.26696
R1684 VP.n7 VP.n3 0.189894
R1685 VP.n11 VP.n3 0.189894
R1686 VP.n12 VP.n11 0.189894
R1687 VP.n13 VP.n12 0.189894
R1688 VP.n13 VP.n1 0.189894
R1689 VP.n17 VP.n1 0.189894
R1690 VDD1 VDD1.n1 110.519
R1691 VDD1 VDD1.n0 64.2348
R1692 VDD1.n0 VDD1.t3 1.30571
R1693 VDD1.n0 VDD1.t0 1.30571
R1694 VDD1.n1 VDD1.t2 1.30571
R1695 VDD1.n1 VDD1.t1 1.30571
C0 VDD2 VN 6.12078f
C1 VTAIL VN 5.96526f
C2 VN VDD1 0.14935f
C3 VDD2 VP 0.429783f
C4 VTAIL VP 5.97937f
C5 VDD2 VTAIL 6.292799f
C6 VDD1 VP 6.40033f
C7 VDD2 VDD1 1.1625f
C8 VTAIL VDD1 6.23484f
C9 VN VP 7.18642f
C10 VDD2 B 4.32529f
C11 VDD1 B 8.985359f
C12 VTAIL B 12.305656f
C13 VN B 12.0371f
C14 VP B 10.35774f
C15 VDD1.t3 B 0.323251f
C16 VDD1.t0 B 0.323251f
C17 VDD1.n0 B 2.9276f
C18 VDD1.t2 B 0.323251f
C19 VDD1.t1 B 0.323251f
C20 VDD1.n1 B 3.75864f
C21 VP.t2 B 2.90322f
C22 VP.n0 B 1.08987f
C23 VP.n1 B 0.022096f
C24 VP.n2 B 0.017863f
C25 VP.n3 B 0.022096f
C26 VP.t1 B 2.90322f
C27 VP.n4 B 1.08987f
C28 VP.t0 B 3.17198f
C29 VP.t3 B 3.16376f
C30 VP.n5 B 3.38746f
C31 VP.n6 B 1.36475f
C32 VP.n7 B 0.035663f
C33 VP.n8 B 0.030811f
C34 VP.n9 B 0.041182f
C35 VP.n10 B 0.043916f
C36 VP.n11 B 0.022096f
C37 VP.n12 B 0.022096f
C38 VP.n13 B 0.022096f
C39 VP.n14 B 0.043916f
C40 VP.n15 B 0.041182f
C41 VP.n16 B 0.030811f
C42 VP.n17 B 0.035663f
C43 VP.n18 B 0.054348f
C44 VTAIL.t4 B 2.16505f
C45 VTAIL.n0 B 0.310743f
C46 VTAIL.t3 B 2.16505f
C47 VTAIL.n1 B 0.385416f
C48 VTAIL.t2 B 2.16505f
C49 VTAIL.n2 B 1.40948f
C50 VTAIL.t7 B 2.16505f
C51 VTAIL.n3 B 1.40948f
C52 VTAIL.t6 B 2.16505f
C53 VTAIL.n4 B 0.385414f
C54 VTAIL.t1 B 2.16505f
C55 VTAIL.n5 B 0.385414f
C56 VTAIL.t0 B 2.16505f
C57 VTAIL.n6 B 1.40948f
C58 VTAIL.t5 B 2.16505f
C59 VTAIL.n7 B 1.3288f
C60 VDD2.t1 B 0.320655f
C61 VDD2.t3 B 0.320655f
C62 VDD2.n0 B 3.70108f
C63 VDD2.t2 B 0.320655f
C64 VDD2.t0 B 0.320655f
C65 VDD2.n1 B 2.90364f
C66 VDD2.n2 B 4.24759f
C67 VN.t2 B 3.1104f
C68 VN.t3 B 3.11849f
C69 VN.n0 B 1.9339f
C70 VN.t0 B 3.1104f
C71 VN.t1 B 3.11849f
C72 VN.n1 B 3.339f
.ends

