* NGSPICE file created from diff_pair_sample_0913.ext - technology: sky130A

.subckt diff_pair_sample_0913 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t7 VN.t0 VTAIL.t8 w_n2420_n1178# sky130_fd_pr__pfet_01v8 ad=0.17325 pd=1.38 as=0.17325 ps=1.38 w=1.05 l=1.12
X1 VDD1.t7 VP.t0 VTAIL.t1 w_n2420_n1178# sky130_fd_pr__pfet_01v8 ad=0.17325 pd=1.38 as=0.17325 ps=1.38 w=1.05 l=1.12
X2 VTAIL.t3 VP.t1 VDD1.t6 w_n2420_n1178# sky130_fd_pr__pfet_01v8 ad=0.17325 pd=1.38 as=0.17325 ps=1.38 w=1.05 l=1.12
X3 VDD2.t6 VN.t1 VTAIL.t11 w_n2420_n1178# sky130_fd_pr__pfet_01v8 ad=0.17325 pd=1.38 as=0.4095 ps=2.88 w=1.05 l=1.12
X4 VDD2.t5 VN.t2 VTAIL.t15 w_n2420_n1178# sky130_fd_pr__pfet_01v8 ad=0.17325 pd=1.38 as=0.17325 ps=1.38 w=1.05 l=1.12
X5 B.t11 B.t9 B.t10 w_n2420_n1178# sky130_fd_pr__pfet_01v8 ad=0.4095 pd=2.88 as=0 ps=0 w=1.05 l=1.12
X6 VTAIL.t5 VP.t2 VDD1.t5 w_n2420_n1178# sky130_fd_pr__pfet_01v8 ad=0.4095 pd=2.88 as=0.17325 ps=1.38 w=1.05 l=1.12
X7 B.t8 B.t6 B.t7 w_n2420_n1178# sky130_fd_pr__pfet_01v8 ad=0.4095 pd=2.88 as=0 ps=0 w=1.05 l=1.12
X8 VTAIL.t10 VN.t3 VDD2.t4 w_n2420_n1178# sky130_fd_pr__pfet_01v8 ad=0.4095 pd=2.88 as=0.17325 ps=1.38 w=1.05 l=1.12
X9 B.t5 B.t3 B.t4 w_n2420_n1178# sky130_fd_pr__pfet_01v8 ad=0.4095 pd=2.88 as=0 ps=0 w=1.05 l=1.12
X10 VDD2.t3 VN.t4 VTAIL.t14 w_n2420_n1178# sky130_fd_pr__pfet_01v8 ad=0.17325 pd=1.38 as=0.4095 ps=2.88 w=1.05 l=1.12
X11 VTAIL.t0 VP.t3 VDD1.t4 w_n2420_n1178# sky130_fd_pr__pfet_01v8 ad=0.17325 pd=1.38 as=0.17325 ps=1.38 w=1.05 l=1.12
X12 VTAIL.t13 VN.t5 VDD2.t2 w_n2420_n1178# sky130_fd_pr__pfet_01v8 ad=0.17325 pd=1.38 as=0.17325 ps=1.38 w=1.05 l=1.12
X13 VDD1.t3 VP.t4 VTAIL.t7 w_n2420_n1178# sky130_fd_pr__pfet_01v8 ad=0.17325 pd=1.38 as=0.4095 ps=2.88 w=1.05 l=1.12
X14 B.t2 B.t0 B.t1 w_n2420_n1178# sky130_fd_pr__pfet_01v8 ad=0.4095 pd=2.88 as=0 ps=0 w=1.05 l=1.12
X15 VTAIL.t9 VN.t6 VDD2.t1 w_n2420_n1178# sky130_fd_pr__pfet_01v8 ad=0.4095 pd=2.88 as=0.17325 ps=1.38 w=1.05 l=1.12
X16 VDD1.t2 VP.t5 VTAIL.t2 w_n2420_n1178# sky130_fd_pr__pfet_01v8 ad=0.17325 pd=1.38 as=0.4095 ps=2.88 w=1.05 l=1.12
X17 VTAIL.t4 VP.t6 VDD1.t1 w_n2420_n1178# sky130_fd_pr__pfet_01v8 ad=0.4095 pd=2.88 as=0.17325 ps=1.38 w=1.05 l=1.12
X18 VDD1.t0 VP.t7 VTAIL.t6 w_n2420_n1178# sky130_fd_pr__pfet_01v8 ad=0.17325 pd=1.38 as=0.17325 ps=1.38 w=1.05 l=1.12
X19 VTAIL.t12 VN.t7 VDD2.t0 w_n2420_n1178# sky130_fd_pr__pfet_01v8 ad=0.17325 pd=1.38 as=0.17325 ps=1.38 w=1.05 l=1.12
R0 VN.n23 VN.n13 161.3
R1 VN.n22 VN.n21 161.3
R2 VN.n20 VN.n19 161.3
R3 VN.n18 VN.n15 161.3
R4 VN.n10 VN.n0 161.3
R5 VN.n9 VN.n8 161.3
R6 VN.n7 VN.n6 161.3
R7 VN.n5 VN.n2 161.3
R8 VN.n3 VN.t6 80.7457
R9 VN.n16 VN.t1 80.7457
R10 VN.n25 VN.n24 80.6037
R11 VN.n12 VN.n11 80.6037
R12 VN.n11 VN.t4 57.8835
R13 VN.n24 VN.t3 57.8835
R14 VN.n6 VN.n5 56.5193
R15 VN.n19 VN.n18 56.5193
R16 VN.n11 VN.n10 49.9132
R17 VN.n24 VN.n23 49.9132
R18 VN VN.n25 36.1506
R19 VN.n4 VN.n3 33.7295
R20 VN.n17 VN.n16 33.7295
R21 VN.n16 VN.n15 28.2143
R22 VN.n3 VN.n2 28.2143
R23 VN.n10 VN.n9 24.4675
R24 VN.n23 VN.n22 24.4675
R25 VN.n5 VN.n4 23.2442
R26 VN.n6 VN.n1 23.2442
R27 VN.n18 VN.n17 23.2442
R28 VN.n19 VN.n14 23.2442
R29 VN.n4 VN.t2 22.5943
R30 VN.n1 VN.t7 22.5943
R31 VN.n17 VN.t5 22.5943
R32 VN.n14 VN.t0 22.5943
R33 VN.n9 VN.n1 1.22385
R34 VN.n22 VN.n14 1.22385
R35 VN.n25 VN.n13 0.285035
R36 VN.n12 VN.n0 0.285035
R37 VN.n21 VN.n13 0.189894
R38 VN.n21 VN.n20 0.189894
R39 VN.n20 VN.n15 0.189894
R40 VN.n7 VN.n2 0.189894
R41 VN.n8 VN.n7 0.189894
R42 VN.n8 VN.n0 0.189894
R43 VN VN.n12 0.146778
R44 VTAIL.n15 VTAIL.t14 371.553
R45 VTAIL.n2 VTAIL.t9 371.553
R46 VTAIL.n3 VTAIL.t7 371.553
R47 VTAIL.n6 VTAIL.t5 371.553
R48 VTAIL.n14 VTAIL.t2 371.553
R49 VTAIL.n11 VTAIL.t4 371.553
R50 VTAIL.n10 VTAIL.t11 371.553
R51 VTAIL.n7 VTAIL.t10 371.553
R52 VTAIL.n1 VTAIL.n0 328.615
R53 VTAIL.n5 VTAIL.n4 328.615
R54 VTAIL.n13 VTAIL.n12 328.615
R55 VTAIL.n9 VTAIL.n8 328.615
R56 VTAIL.n0 VTAIL.t15 30.9576
R57 VTAIL.n0 VTAIL.t12 30.9576
R58 VTAIL.n4 VTAIL.t6 30.9576
R59 VTAIL.n4 VTAIL.t3 30.9576
R60 VTAIL.n12 VTAIL.t1 30.9576
R61 VTAIL.n12 VTAIL.t0 30.9576
R62 VTAIL.n8 VTAIL.t8 30.9576
R63 VTAIL.n8 VTAIL.t13 30.9576
R64 VTAIL.n15 VTAIL.n14 14.5221
R65 VTAIL.n7 VTAIL.n6 14.5221
R66 VTAIL.n9 VTAIL.n7 1.2505
R67 VTAIL.n10 VTAIL.n9 1.2505
R68 VTAIL.n13 VTAIL.n11 1.2505
R69 VTAIL.n14 VTAIL.n13 1.2505
R70 VTAIL.n6 VTAIL.n5 1.2505
R71 VTAIL.n5 VTAIL.n3 1.2505
R72 VTAIL.n2 VTAIL.n1 1.2505
R73 VTAIL VTAIL.n15 1.19231
R74 VTAIL.n11 VTAIL.n10 0.470328
R75 VTAIL.n3 VTAIL.n2 0.470328
R76 VTAIL VTAIL.n1 0.0586897
R77 VDD2.n2 VDD2.n1 345.863
R78 VDD2.n2 VDD2.n0 345.863
R79 VDD2 VDD2.n5 345.861
R80 VDD2.n4 VDD2.n3 345.293
R81 VDD2.n5 VDD2.t2 30.9576
R82 VDD2.n5 VDD2.t6 30.9576
R83 VDD2.n3 VDD2.t4 30.9576
R84 VDD2.n3 VDD2.t7 30.9576
R85 VDD2.n1 VDD2.t0 30.9576
R86 VDD2.n1 VDD2.t3 30.9576
R87 VDD2.n0 VDD2.t1 30.9576
R88 VDD2.n0 VDD2.t5 30.9576
R89 VDD2.n4 VDD2.n2 30.2455
R90 VDD2 VDD2.n4 0.68369
R91 VP.n9 VP.n6 161.3
R92 VP.n11 VP.n10 161.3
R93 VP.n13 VP.n12 161.3
R94 VP.n14 VP.n4 161.3
R95 VP.n28 VP.n0 161.3
R96 VP.n27 VP.n26 161.3
R97 VP.n25 VP.n24 161.3
R98 VP.n23 VP.n2 161.3
R99 VP.n21 VP.n20 161.3
R100 VP.n19 VP.n3 161.3
R101 VP.n7 VP.t6 80.7457
R102 VP.n16 VP.n15 80.6037
R103 VP.n30 VP.n29 80.6037
R104 VP.n18 VP.n17 80.6037
R105 VP.n17 VP.t2 57.8835
R106 VP.n29 VP.t4 57.8835
R107 VP.n15 VP.t5 57.8835
R108 VP.n24 VP.n23 56.5193
R109 VP.n10 VP.n9 56.5193
R110 VP.n17 VP.n3 49.9132
R111 VP.n29 VP.n28 49.9132
R112 VP.n15 VP.n14 49.9132
R113 VP.n18 VP.n16 35.865
R114 VP.n8 VP.n7 33.7295
R115 VP.n7 VP.n6 28.2143
R116 VP.n21 VP.n3 24.4675
R117 VP.n28 VP.n27 24.4675
R118 VP.n14 VP.n13 24.4675
R119 VP.n23 VP.n22 23.2442
R120 VP.n24 VP.n1 23.2442
R121 VP.n10 VP.n5 23.2442
R122 VP.n9 VP.n8 23.2442
R123 VP.n22 VP.t7 22.5943
R124 VP.n1 VP.t1 22.5943
R125 VP.n5 VP.t3 22.5943
R126 VP.n8 VP.t0 22.5943
R127 VP.n22 VP.n21 1.22385
R128 VP.n27 VP.n1 1.22385
R129 VP.n13 VP.n5 1.22385
R130 VP.n16 VP.n4 0.285035
R131 VP.n19 VP.n18 0.285035
R132 VP.n30 VP.n0 0.285035
R133 VP.n11 VP.n6 0.189894
R134 VP.n12 VP.n11 0.189894
R135 VP.n12 VP.n4 0.189894
R136 VP.n20 VP.n19 0.189894
R137 VP.n20 VP.n2 0.189894
R138 VP.n25 VP.n2 0.189894
R139 VP.n26 VP.n25 0.189894
R140 VP.n26 VP.n0 0.189894
R141 VP VP.n30 0.146778
R142 VDD1 VDD1.n0 345.976
R143 VDD1.n3 VDD1.n2 345.863
R144 VDD1.n3 VDD1.n1 345.863
R145 VDD1.n5 VDD1.n4 345.295
R146 VDD1.n4 VDD1.t4 30.9576
R147 VDD1.n4 VDD1.t2 30.9576
R148 VDD1.n0 VDD1.t1 30.9576
R149 VDD1.n0 VDD1.t7 30.9576
R150 VDD1.n2 VDD1.t6 30.9576
R151 VDD1.n2 VDD1.t3 30.9576
R152 VDD1.n1 VDD1.t5 30.9576
R153 VDD1.n1 VDD1.t0 30.9576
R154 VDD1.n5 VDD1.n3 30.8285
R155 VDD1 VDD1.n5 0.56731
R156 B.n182 B.n65 585
R157 B.n181 B.n180 585
R158 B.n179 B.n66 585
R159 B.n178 B.n177 585
R160 B.n176 B.n67 585
R161 B.n175 B.n174 585
R162 B.n173 B.n68 585
R163 B.n172 B.n171 585
R164 B.n170 B.n69 585
R165 B.n168 B.n167 585
R166 B.n166 B.n72 585
R167 B.n165 B.n164 585
R168 B.n163 B.n73 585
R169 B.n162 B.n161 585
R170 B.n160 B.n74 585
R171 B.n159 B.n158 585
R172 B.n157 B.n75 585
R173 B.n156 B.n155 585
R174 B.n154 B.n76 585
R175 B.n153 B.n152 585
R176 B.n148 B.n77 585
R177 B.n147 B.n146 585
R178 B.n145 B.n78 585
R179 B.n144 B.n143 585
R180 B.n142 B.n79 585
R181 B.n141 B.n140 585
R182 B.n139 B.n80 585
R183 B.n138 B.n137 585
R184 B.n184 B.n183 585
R185 B.n185 B.n64 585
R186 B.n187 B.n186 585
R187 B.n188 B.n63 585
R188 B.n190 B.n189 585
R189 B.n191 B.n62 585
R190 B.n193 B.n192 585
R191 B.n194 B.n61 585
R192 B.n196 B.n195 585
R193 B.n197 B.n60 585
R194 B.n199 B.n198 585
R195 B.n200 B.n59 585
R196 B.n202 B.n201 585
R197 B.n203 B.n58 585
R198 B.n205 B.n204 585
R199 B.n206 B.n57 585
R200 B.n208 B.n207 585
R201 B.n209 B.n56 585
R202 B.n211 B.n210 585
R203 B.n212 B.n55 585
R204 B.n214 B.n213 585
R205 B.n215 B.n54 585
R206 B.n217 B.n216 585
R207 B.n218 B.n53 585
R208 B.n220 B.n219 585
R209 B.n221 B.n52 585
R210 B.n223 B.n222 585
R211 B.n224 B.n51 585
R212 B.n226 B.n225 585
R213 B.n227 B.n50 585
R214 B.n229 B.n228 585
R215 B.n230 B.n49 585
R216 B.n232 B.n231 585
R217 B.n233 B.n48 585
R218 B.n235 B.n234 585
R219 B.n236 B.n47 585
R220 B.n238 B.n237 585
R221 B.n239 B.n46 585
R222 B.n241 B.n240 585
R223 B.n242 B.n45 585
R224 B.n244 B.n243 585
R225 B.n245 B.n44 585
R226 B.n247 B.n246 585
R227 B.n248 B.n43 585
R228 B.n250 B.n249 585
R229 B.n251 B.n42 585
R230 B.n253 B.n252 585
R231 B.n254 B.n41 585
R232 B.n256 B.n255 585
R233 B.n257 B.n40 585
R234 B.n259 B.n258 585
R235 B.n260 B.n39 585
R236 B.n262 B.n261 585
R237 B.n263 B.n38 585
R238 B.n265 B.n264 585
R239 B.n266 B.n37 585
R240 B.n268 B.n267 585
R241 B.n269 B.n36 585
R242 B.n271 B.n270 585
R243 B.n272 B.n35 585
R244 B.n316 B.n315 585
R245 B.n314 B.n17 585
R246 B.n313 B.n312 585
R247 B.n311 B.n18 585
R248 B.n310 B.n309 585
R249 B.n308 B.n19 585
R250 B.n307 B.n306 585
R251 B.n305 B.n20 585
R252 B.n304 B.n303 585
R253 B.n301 B.n21 585
R254 B.n300 B.n299 585
R255 B.n298 B.n24 585
R256 B.n297 B.n296 585
R257 B.n295 B.n25 585
R258 B.n294 B.n293 585
R259 B.n292 B.n26 585
R260 B.n291 B.n290 585
R261 B.n289 B.n27 585
R262 B.n288 B.n287 585
R263 B.n286 B.n285 585
R264 B.n284 B.n31 585
R265 B.n283 B.n282 585
R266 B.n281 B.n32 585
R267 B.n280 B.n279 585
R268 B.n278 B.n33 585
R269 B.n277 B.n276 585
R270 B.n275 B.n34 585
R271 B.n274 B.n273 585
R272 B.n317 B.n16 585
R273 B.n319 B.n318 585
R274 B.n320 B.n15 585
R275 B.n322 B.n321 585
R276 B.n323 B.n14 585
R277 B.n325 B.n324 585
R278 B.n326 B.n13 585
R279 B.n328 B.n327 585
R280 B.n329 B.n12 585
R281 B.n331 B.n330 585
R282 B.n332 B.n11 585
R283 B.n334 B.n333 585
R284 B.n335 B.n10 585
R285 B.n337 B.n336 585
R286 B.n338 B.n9 585
R287 B.n340 B.n339 585
R288 B.n341 B.n8 585
R289 B.n343 B.n342 585
R290 B.n344 B.n7 585
R291 B.n346 B.n345 585
R292 B.n347 B.n6 585
R293 B.n349 B.n348 585
R294 B.n350 B.n5 585
R295 B.n352 B.n351 585
R296 B.n353 B.n4 585
R297 B.n355 B.n354 585
R298 B.n356 B.n3 585
R299 B.n358 B.n357 585
R300 B.n359 B.n0 585
R301 B.n2 B.n1 585
R302 B.n96 B.n95 585
R303 B.n97 B.n94 585
R304 B.n99 B.n98 585
R305 B.n100 B.n93 585
R306 B.n102 B.n101 585
R307 B.n103 B.n92 585
R308 B.n105 B.n104 585
R309 B.n106 B.n91 585
R310 B.n108 B.n107 585
R311 B.n109 B.n90 585
R312 B.n111 B.n110 585
R313 B.n112 B.n89 585
R314 B.n114 B.n113 585
R315 B.n115 B.n88 585
R316 B.n117 B.n116 585
R317 B.n118 B.n87 585
R318 B.n120 B.n119 585
R319 B.n121 B.n86 585
R320 B.n123 B.n122 585
R321 B.n124 B.n85 585
R322 B.n126 B.n125 585
R323 B.n127 B.n84 585
R324 B.n129 B.n128 585
R325 B.n130 B.n83 585
R326 B.n132 B.n131 585
R327 B.n133 B.n82 585
R328 B.n135 B.n134 585
R329 B.n136 B.n81 585
R330 B.n138 B.n81 521.33
R331 B.n184 B.n65 521.33
R332 B.n274 B.n35 521.33
R333 B.n317 B.n316 521.33
R334 B.n149 B.t1 390.291
R335 B.n70 B.t4 390.291
R336 B.n28 B.t8 390.291
R337 B.n22 B.t11 390.291
R338 B.n150 B.t2 362.168
R339 B.n71 B.t5 362.168
R340 B.n29 B.t7 362.168
R341 B.n23 B.t10 362.168
R342 B.n361 B.n360 256.663
R343 B.n360 B.n359 235.042
R344 B.n360 B.n2 235.042
R345 B.n149 B.t0 226.272
R346 B.n70 B.t3 226.272
R347 B.n28 B.t6 226.272
R348 B.n22 B.t9 226.272
R349 B.n139 B.n138 163.367
R350 B.n140 B.n139 163.367
R351 B.n140 B.n79 163.367
R352 B.n144 B.n79 163.367
R353 B.n145 B.n144 163.367
R354 B.n146 B.n145 163.367
R355 B.n146 B.n77 163.367
R356 B.n153 B.n77 163.367
R357 B.n154 B.n153 163.367
R358 B.n155 B.n154 163.367
R359 B.n155 B.n75 163.367
R360 B.n159 B.n75 163.367
R361 B.n160 B.n159 163.367
R362 B.n161 B.n160 163.367
R363 B.n161 B.n73 163.367
R364 B.n165 B.n73 163.367
R365 B.n166 B.n165 163.367
R366 B.n167 B.n166 163.367
R367 B.n167 B.n69 163.367
R368 B.n172 B.n69 163.367
R369 B.n173 B.n172 163.367
R370 B.n174 B.n173 163.367
R371 B.n174 B.n67 163.367
R372 B.n178 B.n67 163.367
R373 B.n179 B.n178 163.367
R374 B.n180 B.n179 163.367
R375 B.n180 B.n65 163.367
R376 B.n270 B.n35 163.367
R377 B.n270 B.n269 163.367
R378 B.n269 B.n268 163.367
R379 B.n268 B.n37 163.367
R380 B.n264 B.n37 163.367
R381 B.n264 B.n263 163.367
R382 B.n263 B.n262 163.367
R383 B.n262 B.n39 163.367
R384 B.n258 B.n39 163.367
R385 B.n258 B.n257 163.367
R386 B.n257 B.n256 163.367
R387 B.n256 B.n41 163.367
R388 B.n252 B.n41 163.367
R389 B.n252 B.n251 163.367
R390 B.n251 B.n250 163.367
R391 B.n250 B.n43 163.367
R392 B.n246 B.n43 163.367
R393 B.n246 B.n245 163.367
R394 B.n245 B.n244 163.367
R395 B.n244 B.n45 163.367
R396 B.n240 B.n45 163.367
R397 B.n240 B.n239 163.367
R398 B.n239 B.n238 163.367
R399 B.n238 B.n47 163.367
R400 B.n234 B.n47 163.367
R401 B.n234 B.n233 163.367
R402 B.n233 B.n232 163.367
R403 B.n232 B.n49 163.367
R404 B.n228 B.n49 163.367
R405 B.n228 B.n227 163.367
R406 B.n227 B.n226 163.367
R407 B.n226 B.n51 163.367
R408 B.n222 B.n51 163.367
R409 B.n222 B.n221 163.367
R410 B.n221 B.n220 163.367
R411 B.n220 B.n53 163.367
R412 B.n216 B.n53 163.367
R413 B.n216 B.n215 163.367
R414 B.n215 B.n214 163.367
R415 B.n214 B.n55 163.367
R416 B.n210 B.n55 163.367
R417 B.n210 B.n209 163.367
R418 B.n209 B.n208 163.367
R419 B.n208 B.n57 163.367
R420 B.n204 B.n57 163.367
R421 B.n204 B.n203 163.367
R422 B.n203 B.n202 163.367
R423 B.n202 B.n59 163.367
R424 B.n198 B.n59 163.367
R425 B.n198 B.n197 163.367
R426 B.n197 B.n196 163.367
R427 B.n196 B.n61 163.367
R428 B.n192 B.n61 163.367
R429 B.n192 B.n191 163.367
R430 B.n191 B.n190 163.367
R431 B.n190 B.n63 163.367
R432 B.n186 B.n63 163.367
R433 B.n186 B.n185 163.367
R434 B.n185 B.n184 163.367
R435 B.n316 B.n17 163.367
R436 B.n312 B.n17 163.367
R437 B.n312 B.n311 163.367
R438 B.n311 B.n310 163.367
R439 B.n310 B.n19 163.367
R440 B.n306 B.n19 163.367
R441 B.n306 B.n305 163.367
R442 B.n305 B.n304 163.367
R443 B.n304 B.n21 163.367
R444 B.n299 B.n21 163.367
R445 B.n299 B.n298 163.367
R446 B.n298 B.n297 163.367
R447 B.n297 B.n25 163.367
R448 B.n293 B.n25 163.367
R449 B.n293 B.n292 163.367
R450 B.n292 B.n291 163.367
R451 B.n291 B.n27 163.367
R452 B.n287 B.n27 163.367
R453 B.n287 B.n286 163.367
R454 B.n286 B.n31 163.367
R455 B.n282 B.n31 163.367
R456 B.n282 B.n281 163.367
R457 B.n281 B.n280 163.367
R458 B.n280 B.n33 163.367
R459 B.n276 B.n33 163.367
R460 B.n276 B.n275 163.367
R461 B.n275 B.n274 163.367
R462 B.n318 B.n317 163.367
R463 B.n318 B.n15 163.367
R464 B.n322 B.n15 163.367
R465 B.n323 B.n322 163.367
R466 B.n324 B.n323 163.367
R467 B.n324 B.n13 163.367
R468 B.n328 B.n13 163.367
R469 B.n329 B.n328 163.367
R470 B.n330 B.n329 163.367
R471 B.n330 B.n11 163.367
R472 B.n334 B.n11 163.367
R473 B.n335 B.n334 163.367
R474 B.n336 B.n335 163.367
R475 B.n336 B.n9 163.367
R476 B.n340 B.n9 163.367
R477 B.n341 B.n340 163.367
R478 B.n342 B.n341 163.367
R479 B.n342 B.n7 163.367
R480 B.n346 B.n7 163.367
R481 B.n347 B.n346 163.367
R482 B.n348 B.n347 163.367
R483 B.n348 B.n5 163.367
R484 B.n352 B.n5 163.367
R485 B.n353 B.n352 163.367
R486 B.n354 B.n353 163.367
R487 B.n354 B.n3 163.367
R488 B.n358 B.n3 163.367
R489 B.n359 B.n358 163.367
R490 B.n96 B.n2 163.367
R491 B.n97 B.n96 163.367
R492 B.n98 B.n97 163.367
R493 B.n98 B.n93 163.367
R494 B.n102 B.n93 163.367
R495 B.n103 B.n102 163.367
R496 B.n104 B.n103 163.367
R497 B.n104 B.n91 163.367
R498 B.n108 B.n91 163.367
R499 B.n109 B.n108 163.367
R500 B.n110 B.n109 163.367
R501 B.n110 B.n89 163.367
R502 B.n114 B.n89 163.367
R503 B.n115 B.n114 163.367
R504 B.n116 B.n115 163.367
R505 B.n116 B.n87 163.367
R506 B.n120 B.n87 163.367
R507 B.n121 B.n120 163.367
R508 B.n122 B.n121 163.367
R509 B.n122 B.n85 163.367
R510 B.n126 B.n85 163.367
R511 B.n127 B.n126 163.367
R512 B.n128 B.n127 163.367
R513 B.n128 B.n83 163.367
R514 B.n132 B.n83 163.367
R515 B.n133 B.n132 163.367
R516 B.n134 B.n133 163.367
R517 B.n134 B.n81 163.367
R518 B.n151 B.n150 59.5399
R519 B.n169 B.n71 59.5399
R520 B.n30 B.n29 59.5399
R521 B.n302 B.n23 59.5399
R522 B.n315 B.n16 33.8737
R523 B.n273 B.n272 33.8737
R524 B.n183 B.n182 33.8737
R525 B.n137 B.n136 33.8737
R526 B.n150 B.n149 28.1217
R527 B.n71 B.n70 28.1217
R528 B.n29 B.n28 28.1217
R529 B.n23 B.n22 28.1217
R530 B B.n361 18.0485
R531 B.n319 B.n16 10.6151
R532 B.n320 B.n319 10.6151
R533 B.n321 B.n320 10.6151
R534 B.n321 B.n14 10.6151
R535 B.n325 B.n14 10.6151
R536 B.n326 B.n325 10.6151
R537 B.n327 B.n326 10.6151
R538 B.n327 B.n12 10.6151
R539 B.n331 B.n12 10.6151
R540 B.n332 B.n331 10.6151
R541 B.n333 B.n332 10.6151
R542 B.n333 B.n10 10.6151
R543 B.n337 B.n10 10.6151
R544 B.n338 B.n337 10.6151
R545 B.n339 B.n338 10.6151
R546 B.n339 B.n8 10.6151
R547 B.n343 B.n8 10.6151
R548 B.n344 B.n343 10.6151
R549 B.n345 B.n344 10.6151
R550 B.n345 B.n6 10.6151
R551 B.n349 B.n6 10.6151
R552 B.n350 B.n349 10.6151
R553 B.n351 B.n350 10.6151
R554 B.n351 B.n4 10.6151
R555 B.n355 B.n4 10.6151
R556 B.n356 B.n355 10.6151
R557 B.n357 B.n356 10.6151
R558 B.n357 B.n0 10.6151
R559 B.n315 B.n314 10.6151
R560 B.n314 B.n313 10.6151
R561 B.n313 B.n18 10.6151
R562 B.n309 B.n18 10.6151
R563 B.n309 B.n308 10.6151
R564 B.n308 B.n307 10.6151
R565 B.n307 B.n20 10.6151
R566 B.n303 B.n20 10.6151
R567 B.n301 B.n300 10.6151
R568 B.n300 B.n24 10.6151
R569 B.n296 B.n24 10.6151
R570 B.n296 B.n295 10.6151
R571 B.n295 B.n294 10.6151
R572 B.n294 B.n26 10.6151
R573 B.n290 B.n26 10.6151
R574 B.n290 B.n289 10.6151
R575 B.n289 B.n288 10.6151
R576 B.n285 B.n284 10.6151
R577 B.n284 B.n283 10.6151
R578 B.n283 B.n32 10.6151
R579 B.n279 B.n32 10.6151
R580 B.n279 B.n278 10.6151
R581 B.n278 B.n277 10.6151
R582 B.n277 B.n34 10.6151
R583 B.n273 B.n34 10.6151
R584 B.n272 B.n271 10.6151
R585 B.n271 B.n36 10.6151
R586 B.n267 B.n36 10.6151
R587 B.n267 B.n266 10.6151
R588 B.n266 B.n265 10.6151
R589 B.n265 B.n38 10.6151
R590 B.n261 B.n38 10.6151
R591 B.n261 B.n260 10.6151
R592 B.n260 B.n259 10.6151
R593 B.n259 B.n40 10.6151
R594 B.n255 B.n40 10.6151
R595 B.n255 B.n254 10.6151
R596 B.n254 B.n253 10.6151
R597 B.n253 B.n42 10.6151
R598 B.n249 B.n42 10.6151
R599 B.n249 B.n248 10.6151
R600 B.n248 B.n247 10.6151
R601 B.n247 B.n44 10.6151
R602 B.n243 B.n44 10.6151
R603 B.n243 B.n242 10.6151
R604 B.n242 B.n241 10.6151
R605 B.n241 B.n46 10.6151
R606 B.n237 B.n46 10.6151
R607 B.n237 B.n236 10.6151
R608 B.n236 B.n235 10.6151
R609 B.n235 B.n48 10.6151
R610 B.n231 B.n48 10.6151
R611 B.n231 B.n230 10.6151
R612 B.n230 B.n229 10.6151
R613 B.n229 B.n50 10.6151
R614 B.n225 B.n50 10.6151
R615 B.n225 B.n224 10.6151
R616 B.n224 B.n223 10.6151
R617 B.n223 B.n52 10.6151
R618 B.n219 B.n52 10.6151
R619 B.n219 B.n218 10.6151
R620 B.n218 B.n217 10.6151
R621 B.n217 B.n54 10.6151
R622 B.n213 B.n54 10.6151
R623 B.n213 B.n212 10.6151
R624 B.n212 B.n211 10.6151
R625 B.n211 B.n56 10.6151
R626 B.n207 B.n56 10.6151
R627 B.n207 B.n206 10.6151
R628 B.n206 B.n205 10.6151
R629 B.n205 B.n58 10.6151
R630 B.n201 B.n58 10.6151
R631 B.n201 B.n200 10.6151
R632 B.n200 B.n199 10.6151
R633 B.n199 B.n60 10.6151
R634 B.n195 B.n60 10.6151
R635 B.n195 B.n194 10.6151
R636 B.n194 B.n193 10.6151
R637 B.n193 B.n62 10.6151
R638 B.n189 B.n62 10.6151
R639 B.n189 B.n188 10.6151
R640 B.n188 B.n187 10.6151
R641 B.n187 B.n64 10.6151
R642 B.n183 B.n64 10.6151
R643 B.n95 B.n1 10.6151
R644 B.n95 B.n94 10.6151
R645 B.n99 B.n94 10.6151
R646 B.n100 B.n99 10.6151
R647 B.n101 B.n100 10.6151
R648 B.n101 B.n92 10.6151
R649 B.n105 B.n92 10.6151
R650 B.n106 B.n105 10.6151
R651 B.n107 B.n106 10.6151
R652 B.n107 B.n90 10.6151
R653 B.n111 B.n90 10.6151
R654 B.n112 B.n111 10.6151
R655 B.n113 B.n112 10.6151
R656 B.n113 B.n88 10.6151
R657 B.n117 B.n88 10.6151
R658 B.n118 B.n117 10.6151
R659 B.n119 B.n118 10.6151
R660 B.n119 B.n86 10.6151
R661 B.n123 B.n86 10.6151
R662 B.n124 B.n123 10.6151
R663 B.n125 B.n124 10.6151
R664 B.n125 B.n84 10.6151
R665 B.n129 B.n84 10.6151
R666 B.n130 B.n129 10.6151
R667 B.n131 B.n130 10.6151
R668 B.n131 B.n82 10.6151
R669 B.n135 B.n82 10.6151
R670 B.n136 B.n135 10.6151
R671 B.n137 B.n80 10.6151
R672 B.n141 B.n80 10.6151
R673 B.n142 B.n141 10.6151
R674 B.n143 B.n142 10.6151
R675 B.n143 B.n78 10.6151
R676 B.n147 B.n78 10.6151
R677 B.n148 B.n147 10.6151
R678 B.n152 B.n148 10.6151
R679 B.n156 B.n76 10.6151
R680 B.n157 B.n156 10.6151
R681 B.n158 B.n157 10.6151
R682 B.n158 B.n74 10.6151
R683 B.n162 B.n74 10.6151
R684 B.n163 B.n162 10.6151
R685 B.n164 B.n163 10.6151
R686 B.n164 B.n72 10.6151
R687 B.n168 B.n72 10.6151
R688 B.n171 B.n170 10.6151
R689 B.n171 B.n68 10.6151
R690 B.n175 B.n68 10.6151
R691 B.n176 B.n175 10.6151
R692 B.n177 B.n176 10.6151
R693 B.n177 B.n66 10.6151
R694 B.n181 B.n66 10.6151
R695 B.n182 B.n181 10.6151
R696 B.n303 B.n302 9.36635
R697 B.n285 B.n30 9.36635
R698 B.n152 B.n151 9.36635
R699 B.n170 B.n169 9.36635
R700 B.n361 B.n0 8.11757
R701 B.n361 B.n1 8.11757
R702 B.n302 B.n301 1.24928
R703 B.n288 B.n30 1.24928
R704 B.n151 B.n76 1.24928
R705 B.n169 B.n168 1.24928
C0 B VTAIL 0.919652f
C1 VP VN 3.8323f
C2 w_n2420_n1178# VDD1 1.15687f
C3 VDD2 B 0.951741f
C4 VP VTAIL 1.53861f
C5 B VDD1 0.901723f
C6 VDD2 VP 0.37061f
C7 w_n2420_n1178# B 4.78427f
C8 VTAIL VN 1.52451f
C9 VP VDD1 1.18037f
C10 w_n2420_n1178# VP 4.57371f
C11 VDD2 VN 0.968085f
C12 VDD1 VN 0.156147f
C13 VP B 1.23998f
C14 VDD2 VTAIL 3.15796f
C15 w_n2420_n1178# VN 4.27148f
C16 VDD1 VTAIL 3.11347f
C17 w_n2420_n1178# VTAIL 1.4406f
C18 B VN 0.729744f
C19 VDD2 VDD1 1.03664f
C20 w_n2420_n1178# VDD2 1.20826f
C21 VDD2 VSUBS 0.746128f
C22 VDD1 VSUBS 1.104671f
C23 VTAIL VSUBS 0.315297f
C24 VN VSUBS 4.26144f
C25 VP VSUBS 1.549925f
C26 B VSUBS 2.294001f
C27 w_n2420_n1178# VSUBS 36.735603f
C28 B.n0 VSUBS 0.008626f
C29 B.n1 VSUBS 0.008626f
C30 B.n2 VSUBS 0.012758f
C31 B.n3 VSUBS 0.009777f
C32 B.n4 VSUBS 0.009777f
C33 B.n5 VSUBS 0.009777f
C34 B.n6 VSUBS 0.009777f
C35 B.n7 VSUBS 0.009777f
C36 B.n8 VSUBS 0.009777f
C37 B.n9 VSUBS 0.009777f
C38 B.n10 VSUBS 0.009777f
C39 B.n11 VSUBS 0.009777f
C40 B.n12 VSUBS 0.009777f
C41 B.n13 VSUBS 0.009777f
C42 B.n14 VSUBS 0.009777f
C43 B.n15 VSUBS 0.009777f
C44 B.n16 VSUBS 0.02315f
C45 B.n17 VSUBS 0.009777f
C46 B.n18 VSUBS 0.009777f
C47 B.n19 VSUBS 0.009777f
C48 B.n20 VSUBS 0.009777f
C49 B.n21 VSUBS 0.009777f
C50 B.t10 VSUBS 0.027581f
C51 B.t11 VSUBS 0.030711f
C52 B.t9 VSUBS 0.083354f
C53 B.n22 VSUBS 0.063846f
C54 B.n23 VSUBS 0.057379f
C55 B.n24 VSUBS 0.009777f
C56 B.n25 VSUBS 0.009777f
C57 B.n26 VSUBS 0.009777f
C58 B.n27 VSUBS 0.009777f
C59 B.t7 VSUBS 0.027581f
C60 B.t8 VSUBS 0.030711f
C61 B.t6 VSUBS 0.083354f
C62 B.n28 VSUBS 0.063846f
C63 B.n29 VSUBS 0.057379f
C64 B.n30 VSUBS 0.022652f
C65 B.n31 VSUBS 0.009777f
C66 B.n32 VSUBS 0.009777f
C67 B.n33 VSUBS 0.009777f
C68 B.n34 VSUBS 0.009777f
C69 B.n35 VSUBS 0.02315f
C70 B.n36 VSUBS 0.009777f
C71 B.n37 VSUBS 0.009777f
C72 B.n38 VSUBS 0.009777f
C73 B.n39 VSUBS 0.009777f
C74 B.n40 VSUBS 0.009777f
C75 B.n41 VSUBS 0.009777f
C76 B.n42 VSUBS 0.009777f
C77 B.n43 VSUBS 0.009777f
C78 B.n44 VSUBS 0.009777f
C79 B.n45 VSUBS 0.009777f
C80 B.n46 VSUBS 0.009777f
C81 B.n47 VSUBS 0.009777f
C82 B.n48 VSUBS 0.009777f
C83 B.n49 VSUBS 0.009777f
C84 B.n50 VSUBS 0.009777f
C85 B.n51 VSUBS 0.009777f
C86 B.n52 VSUBS 0.009777f
C87 B.n53 VSUBS 0.009777f
C88 B.n54 VSUBS 0.009777f
C89 B.n55 VSUBS 0.009777f
C90 B.n56 VSUBS 0.009777f
C91 B.n57 VSUBS 0.009777f
C92 B.n58 VSUBS 0.009777f
C93 B.n59 VSUBS 0.009777f
C94 B.n60 VSUBS 0.009777f
C95 B.n61 VSUBS 0.009777f
C96 B.n62 VSUBS 0.009777f
C97 B.n63 VSUBS 0.009777f
C98 B.n64 VSUBS 0.009777f
C99 B.n65 VSUBS 0.023721f
C100 B.n66 VSUBS 0.009777f
C101 B.n67 VSUBS 0.009777f
C102 B.n68 VSUBS 0.009777f
C103 B.n69 VSUBS 0.009777f
C104 B.t5 VSUBS 0.027581f
C105 B.t4 VSUBS 0.030711f
C106 B.t3 VSUBS 0.083354f
C107 B.n70 VSUBS 0.063846f
C108 B.n71 VSUBS 0.057379f
C109 B.n72 VSUBS 0.009777f
C110 B.n73 VSUBS 0.009777f
C111 B.n74 VSUBS 0.009777f
C112 B.n75 VSUBS 0.009777f
C113 B.n76 VSUBS 0.005463f
C114 B.n77 VSUBS 0.009777f
C115 B.n78 VSUBS 0.009777f
C116 B.n79 VSUBS 0.009777f
C117 B.n80 VSUBS 0.009777f
C118 B.n81 VSUBS 0.02315f
C119 B.n82 VSUBS 0.009777f
C120 B.n83 VSUBS 0.009777f
C121 B.n84 VSUBS 0.009777f
C122 B.n85 VSUBS 0.009777f
C123 B.n86 VSUBS 0.009777f
C124 B.n87 VSUBS 0.009777f
C125 B.n88 VSUBS 0.009777f
C126 B.n89 VSUBS 0.009777f
C127 B.n90 VSUBS 0.009777f
C128 B.n91 VSUBS 0.009777f
C129 B.n92 VSUBS 0.009777f
C130 B.n93 VSUBS 0.009777f
C131 B.n94 VSUBS 0.009777f
C132 B.n95 VSUBS 0.009777f
C133 B.n96 VSUBS 0.009777f
C134 B.n97 VSUBS 0.009777f
C135 B.n98 VSUBS 0.009777f
C136 B.n99 VSUBS 0.009777f
C137 B.n100 VSUBS 0.009777f
C138 B.n101 VSUBS 0.009777f
C139 B.n102 VSUBS 0.009777f
C140 B.n103 VSUBS 0.009777f
C141 B.n104 VSUBS 0.009777f
C142 B.n105 VSUBS 0.009777f
C143 B.n106 VSUBS 0.009777f
C144 B.n107 VSUBS 0.009777f
C145 B.n108 VSUBS 0.009777f
C146 B.n109 VSUBS 0.009777f
C147 B.n110 VSUBS 0.009777f
C148 B.n111 VSUBS 0.009777f
C149 B.n112 VSUBS 0.009777f
C150 B.n113 VSUBS 0.009777f
C151 B.n114 VSUBS 0.009777f
C152 B.n115 VSUBS 0.009777f
C153 B.n116 VSUBS 0.009777f
C154 B.n117 VSUBS 0.009777f
C155 B.n118 VSUBS 0.009777f
C156 B.n119 VSUBS 0.009777f
C157 B.n120 VSUBS 0.009777f
C158 B.n121 VSUBS 0.009777f
C159 B.n122 VSUBS 0.009777f
C160 B.n123 VSUBS 0.009777f
C161 B.n124 VSUBS 0.009777f
C162 B.n125 VSUBS 0.009777f
C163 B.n126 VSUBS 0.009777f
C164 B.n127 VSUBS 0.009777f
C165 B.n128 VSUBS 0.009777f
C166 B.n129 VSUBS 0.009777f
C167 B.n130 VSUBS 0.009777f
C168 B.n131 VSUBS 0.009777f
C169 B.n132 VSUBS 0.009777f
C170 B.n133 VSUBS 0.009777f
C171 B.n134 VSUBS 0.009777f
C172 B.n135 VSUBS 0.009777f
C173 B.n136 VSUBS 0.02315f
C174 B.n137 VSUBS 0.023721f
C175 B.n138 VSUBS 0.023721f
C176 B.n139 VSUBS 0.009777f
C177 B.n140 VSUBS 0.009777f
C178 B.n141 VSUBS 0.009777f
C179 B.n142 VSUBS 0.009777f
C180 B.n143 VSUBS 0.009777f
C181 B.n144 VSUBS 0.009777f
C182 B.n145 VSUBS 0.009777f
C183 B.n146 VSUBS 0.009777f
C184 B.n147 VSUBS 0.009777f
C185 B.n148 VSUBS 0.009777f
C186 B.t2 VSUBS 0.027581f
C187 B.t1 VSUBS 0.030711f
C188 B.t0 VSUBS 0.083354f
C189 B.n149 VSUBS 0.063846f
C190 B.n150 VSUBS 0.057379f
C191 B.n151 VSUBS 0.022652f
C192 B.n152 VSUBS 0.009202f
C193 B.n153 VSUBS 0.009777f
C194 B.n154 VSUBS 0.009777f
C195 B.n155 VSUBS 0.009777f
C196 B.n156 VSUBS 0.009777f
C197 B.n157 VSUBS 0.009777f
C198 B.n158 VSUBS 0.009777f
C199 B.n159 VSUBS 0.009777f
C200 B.n160 VSUBS 0.009777f
C201 B.n161 VSUBS 0.009777f
C202 B.n162 VSUBS 0.009777f
C203 B.n163 VSUBS 0.009777f
C204 B.n164 VSUBS 0.009777f
C205 B.n165 VSUBS 0.009777f
C206 B.n166 VSUBS 0.009777f
C207 B.n167 VSUBS 0.009777f
C208 B.n168 VSUBS 0.005463f
C209 B.n169 VSUBS 0.022652f
C210 B.n170 VSUBS 0.009202f
C211 B.n171 VSUBS 0.009777f
C212 B.n172 VSUBS 0.009777f
C213 B.n173 VSUBS 0.009777f
C214 B.n174 VSUBS 0.009777f
C215 B.n175 VSUBS 0.009777f
C216 B.n176 VSUBS 0.009777f
C217 B.n177 VSUBS 0.009777f
C218 B.n178 VSUBS 0.009777f
C219 B.n179 VSUBS 0.009777f
C220 B.n180 VSUBS 0.009777f
C221 B.n181 VSUBS 0.009777f
C222 B.n182 VSUBS 0.022607f
C223 B.n183 VSUBS 0.024264f
C224 B.n184 VSUBS 0.02315f
C225 B.n185 VSUBS 0.009777f
C226 B.n186 VSUBS 0.009777f
C227 B.n187 VSUBS 0.009777f
C228 B.n188 VSUBS 0.009777f
C229 B.n189 VSUBS 0.009777f
C230 B.n190 VSUBS 0.009777f
C231 B.n191 VSUBS 0.009777f
C232 B.n192 VSUBS 0.009777f
C233 B.n193 VSUBS 0.009777f
C234 B.n194 VSUBS 0.009777f
C235 B.n195 VSUBS 0.009777f
C236 B.n196 VSUBS 0.009777f
C237 B.n197 VSUBS 0.009777f
C238 B.n198 VSUBS 0.009777f
C239 B.n199 VSUBS 0.009777f
C240 B.n200 VSUBS 0.009777f
C241 B.n201 VSUBS 0.009777f
C242 B.n202 VSUBS 0.009777f
C243 B.n203 VSUBS 0.009777f
C244 B.n204 VSUBS 0.009777f
C245 B.n205 VSUBS 0.009777f
C246 B.n206 VSUBS 0.009777f
C247 B.n207 VSUBS 0.009777f
C248 B.n208 VSUBS 0.009777f
C249 B.n209 VSUBS 0.009777f
C250 B.n210 VSUBS 0.009777f
C251 B.n211 VSUBS 0.009777f
C252 B.n212 VSUBS 0.009777f
C253 B.n213 VSUBS 0.009777f
C254 B.n214 VSUBS 0.009777f
C255 B.n215 VSUBS 0.009777f
C256 B.n216 VSUBS 0.009777f
C257 B.n217 VSUBS 0.009777f
C258 B.n218 VSUBS 0.009777f
C259 B.n219 VSUBS 0.009777f
C260 B.n220 VSUBS 0.009777f
C261 B.n221 VSUBS 0.009777f
C262 B.n222 VSUBS 0.009777f
C263 B.n223 VSUBS 0.009777f
C264 B.n224 VSUBS 0.009777f
C265 B.n225 VSUBS 0.009777f
C266 B.n226 VSUBS 0.009777f
C267 B.n227 VSUBS 0.009777f
C268 B.n228 VSUBS 0.009777f
C269 B.n229 VSUBS 0.009777f
C270 B.n230 VSUBS 0.009777f
C271 B.n231 VSUBS 0.009777f
C272 B.n232 VSUBS 0.009777f
C273 B.n233 VSUBS 0.009777f
C274 B.n234 VSUBS 0.009777f
C275 B.n235 VSUBS 0.009777f
C276 B.n236 VSUBS 0.009777f
C277 B.n237 VSUBS 0.009777f
C278 B.n238 VSUBS 0.009777f
C279 B.n239 VSUBS 0.009777f
C280 B.n240 VSUBS 0.009777f
C281 B.n241 VSUBS 0.009777f
C282 B.n242 VSUBS 0.009777f
C283 B.n243 VSUBS 0.009777f
C284 B.n244 VSUBS 0.009777f
C285 B.n245 VSUBS 0.009777f
C286 B.n246 VSUBS 0.009777f
C287 B.n247 VSUBS 0.009777f
C288 B.n248 VSUBS 0.009777f
C289 B.n249 VSUBS 0.009777f
C290 B.n250 VSUBS 0.009777f
C291 B.n251 VSUBS 0.009777f
C292 B.n252 VSUBS 0.009777f
C293 B.n253 VSUBS 0.009777f
C294 B.n254 VSUBS 0.009777f
C295 B.n255 VSUBS 0.009777f
C296 B.n256 VSUBS 0.009777f
C297 B.n257 VSUBS 0.009777f
C298 B.n258 VSUBS 0.009777f
C299 B.n259 VSUBS 0.009777f
C300 B.n260 VSUBS 0.009777f
C301 B.n261 VSUBS 0.009777f
C302 B.n262 VSUBS 0.009777f
C303 B.n263 VSUBS 0.009777f
C304 B.n264 VSUBS 0.009777f
C305 B.n265 VSUBS 0.009777f
C306 B.n266 VSUBS 0.009777f
C307 B.n267 VSUBS 0.009777f
C308 B.n268 VSUBS 0.009777f
C309 B.n269 VSUBS 0.009777f
C310 B.n270 VSUBS 0.009777f
C311 B.n271 VSUBS 0.009777f
C312 B.n272 VSUBS 0.02315f
C313 B.n273 VSUBS 0.023721f
C314 B.n274 VSUBS 0.023721f
C315 B.n275 VSUBS 0.009777f
C316 B.n276 VSUBS 0.009777f
C317 B.n277 VSUBS 0.009777f
C318 B.n278 VSUBS 0.009777f
C319 B.n279 VSUBS 0.009777f
C320 B.n280 VSUBS 0.009777f
C321 B.n281 VSUBS 0.009777f
C322 B.n282 VSUBS 0.009777f
C323 B.n283 VSUBS 0.009777f
C324 B.n284 VSUBS 0.009777f
C325 B.n285 VSUBS 0.009202f
C326 B.n286 VSUBS 0.009777f
C327 B.n287 VSUBS 0.009777f
C328 B.n288 VSUBS 0.005463f
C329 B.n289 VSUBS 0.009777f
C330 B.n290 VSUBS 0.009777f
C331 B.n291 VSUBS 0.009777f
C332 B.n292 VSUBS 0.009777f
C333 B.n293 VSUBS 0.009777f
C334 B.n294 VSUBS 0.009777f
C335 B.n295 VSUBS 0.009777f
C336 B.n296 VSUBS 0.009777f
C337 B.n297 VSUBS 0.009777f
C338 B.n298 VSUBS 0.009777f
C339 B.n299 VSUBS 0.009777f
C340 B.n300 VSUBS 0.009777f
C341 B.n301 VSUBS 0.005463f
C342 B.n302 VSUBS 0.022652f
C343 B.n303 VSUBS 0.009202f
C344 B.n304 VSUBS 0.009777f
C345 B.n305 VSUBS 0.009777f
C346 B.n306 VSUBS 0.009777f
C347 B.n307 VSUBS 0.009777f
C348 B.n308 VSUBS 0.009777f
C349 B.n309 VSUBS 0.009777f
C350 B.n310 VSUBS 0.009777f
C351 B.n311 VSUBS 0.009777f
C352 B.n312 VSUBS 0.009777f
C353 B.n313 VSUBS 0.009777f
C354 B.n314 VSUBS 0.009777f
C355 B.n315 VSUBS 0.023721f
C356 B.n316 VSUBS 0.023721f
C357 B.n317 VSUBS 0.02315f
C358 B.n318 VSUBS 0.009777f
C359 B.n319 VSUBS 0.009777f
C360 B.n320 VSUBS 0.009777f
C361 B.n321 VSUBS 0.009777f
C362 B.n322 VSUBS 0.009777f
C363 B.n323 VSUBS 0.009777f
C364 B.n324 VSUBS 0.009777f
C365 B.n325 VSUBS 0.009777f
C366 B.n326 VSUBS 0.009777f
C367 B.n327 VSUBS 0.009777f
C368 B.n328 VSUBS 0.009777f
C369 B.n329 VSUBS 0.009777f
C370 B.n330 VSUBS 0.009777f
C371 B.n331 VSUBS 0.009777f
C372 B.n332 VSUBS 0.009777f
C373 B.n333 VSUBS 0.009777f
C374 B.n334 VSUBS 0.009777f
C375 B.n335 VSUBS 0.009777f
C376 B.n336 VSUBS 0.009777f
C377 B.n337 VSUBS 0.009777f
C378 B.n338 VSUBS 0.009777f
C379 B.n339 VSUBS 0.009777f
C380 B.n340 VSUBS 0.009777f
C381 B.n341 VSUBS 0.009777f
C382 B.n342 VSUBS 0.009777f
C383 B.n343 VSUBS 0.009777f
C384 B.n344 VSUBS 0.009777f
C385 B.n345 VSUBS 0.009777f
C386 B.n346 VSUBS 0.009777f
C387 B.n347 VSUBS 0.009777f
C388 B.n348 VSUBS 0.009777f
C389 B.n349 VSUBS 0.009777f
C390 B.n350 VSUBS 0.009777f
C391 B.n351 VSUBS 0.009777f
C392 B.n352 VSUBS 0.009777f
C393 B.n353 VSUBS 0.009777f
C394 B.n354 VSUBS 0.009777f
C395 B.n355 VSUBS 0.009777f
C396 B.n356 VSUBS 0.009777f
C397 B.n357 VSUBS 0.009777f
C398 B.n358 VSUBS 0.009777f
C399 B.n359 VSUBS 0.012758f
C400 B.n360 VSUBS 0.013591f
C401 B.n361 VSUBS 0.027026f
C402 VDD1.t1 VSUBS 0.01502f
C403 VDD1.t7 VSUBS 0.01502f
C404 VDD1.n0 VSUBS 0.050283f
C405 VDD1.t5 VSUBS 0.01502f
C406 VDD1.t0 VSUBS 0.01502f
C407 VDD1.n1 VSUBS 0.050189f
C408 VDD1.t6 VSUBS 0.01502f
C409 VDD1.t3 VSUBS 0.01502f
C410 VDD1.n2 VSUBS 0.050189f
C411 VDD1.n3 VSUBS 1.30509f
C412 VDD1.t4 VSUBS 0.01502f
C413 VDD1.t2 VSUBS 0.01502f
C414 VDD1.n4 VSUBS 0.049771f
C415 VDD1.n5 VSUBS 1.14265f
C416 VP.n0 VSUBS 0.077801f
C417 VP.t1 VSUBS 0.131154f
C418 VP.n1 VSUBS 0.117696f
C419 VP.n2 VSUBS 0.058305f
C420 VP.t7 VSUBS 0.131154f
C421 VP.n3 VSUBS 0.073849f
C422 VP.n4 VSUBS 0.077801f
C423 VP.t5 VSUBS 0.231198f
C424 VP.t3 VSUBS 0.131154f
C425 VP.n5 VSUBS 0.117696f
C426 VP.n6 VSUBS 0.305541f
C427 VP.t0 VSUBS 0.131154f
C428 VP.t6 VSUBS 0.297436f
C429 VP.n7 VSUBS 0.194372f
C430 VP.n8 VSUBS 0.211003f
C431 VP.n9 VSUBS 0.08243f
C432 VP.n10 VSUBS 0.08243f
C433 VP.n11 VSUBS 0.058305f
C434 VP.n12 VSUBS 0.058305f
C435 VP.n13 VSUBS 0.057697f
C436 VP.n14 VSUBS 0.073849f
C437 VP.n15 VSUBS 0.219491f
C438 VP.n16 VSUBS 1.84092f
C439 VP.t2 VSUBS 0.231198f
C440 VP.n17 VSUBS 0.219491f
C441 VP.n18 VSUBS 1.89936f
C442 VP.n19 VSUBS 0.077801f
C443 VP.n20 VSUBS 0.058305f
C444 VP.n21 VSUBS 0.057697f
C445 VP.n22 VSUBS 0.117696f
C446 VP.n23 VSUBS 0.08243f
C447 VP.n24 VSUBS 0.08243f
C448 VP.n25 VSUBS 0.058305f
C449 VP.n26 VSUBS 0.058305f
C450 VP.n27 VSUBS 0.057697f
C451 VP.n28 VSUBS 0.073849f
C452 VP.t4 VSUBS 0.231198f
C453 VP.n29 VSUBS 0.219491f
C454 VP.n30 VSUBS 0.054605f
C455 VDD2.t1 VSUBS 0.015847f
C456 VDD2.t5 VSUBS 0.015847f
C457 VDD2.n0 VSUBS 0.05295f
C458 VDD2.t0 VSUBS 0.015847f
C459 VDD2.t3 VSUBS 0.015847f
C460 VDD2.n1 VSUBS 0.05295f
C461 VDD2.n2 VSUBS 1.33623f
C462 VDD2.t4 VSUBS 0.015847f
C463 VDD2.t7 VSUBS 0.015847f
C464 VDD2.n3 VSUBS 0.052509f
C465 VDD2.n4 VSUBS 1.18278f
C466 VDD2.t2 VSUBS 0.015847f
C467 VDD2.t6 VSUBS 0.015847f
C468 VDD2.n5 VSUBS 0.052946f
C469 VTAIL.t15 VSUBS 0.018257f
C470 VTAIL.t12 VSUBS 0.018257f
C471 VTAIL.n0 VSUBS 0.052121f
C472 VTAIL.n1 VSUBS 0.24043f
C473 VTAIL.t9 VSUBS 0.091751f
C474 VTAIL.n2 VSUBS 0.279777f
C475 VTAIL.t7 VSUBS 0.091751f
C476 VTAIL.n3 VSUBS 0.279777f
C477 VTAIL.t6 VSUBS 0.018257f
C478 VTAIL.t3 VSUBS 0.018257f
C479 VTAIL.n4 VSUBS 0.052121f
C480 VTAIL.n5 VSUBS 0.324929f
C481 VTAIL.t5 VSUBS 0.091751f
C482 VTAIL.n6 VSUBS 0.698157f
C483 VTAIL.t10 VSUBS 0.091751f
C484 VTAIL.n7 VSUBS 0.698157f
C485 VTAIL.t8 VSUBS 0.018257f
C486 VTAIL.t13 VSUBS 0.018257f
C487 VTAIL.n8 VSUBS 0.052121f
C488 VTAIL.n9 VSUBS 0.324929f
C489 VTAIL.t11 VSUBS 0.091751f
C490 VTAIL.n10 VSUBS 0.279777f
C491 VTAIL.t4 VSUBS 0.091751f
C492 VTAIL.n11 VSUBS 0.279777f
C493 VTAIL.t1 VSUBS 0.018257f
C494 VTAIL.t0 VSUBS 0.018257f
C495 VTAIL.n12 VSUBS 0.052121f
C496 VTAIL.n13 VSUBS 0.324929f
C497 VTAIL.t2 VSUBS 0.091751f
C498 VTAIL.n14 VSUBS 0.698157f
C499 VTAIL.t14 VSUBS 0.091751f
C500 VTAIL.n15 VSUBS 0.694031f
C501 VN.n0 VSUBS 0.074297f
C502 VN.t7 VSUBS 0.125248f
C503 VN.n1 VSUBS 0.112396f
C504 VN.n2 VSUBS 0.291782f
C505 VN.t2 VSUBS 0.125248f
C506 VN.t6 VSUBS 0.284042f
C507 VN.n3 VSUBS 0.185619f
C508 VN.n4 VSUBS 0.201501f
C509 VN.n5 VSUBS 0.078718f
C510 VN.n6 VSUBS 0.078718f
C511 VN.n7 VSUBS 0.05568f
C512 VN.n8 VSUBS 0.05568f
C513 VN.n9 VSUBS 0.055099f
C514 VN.n10 VSUBS 0.070524f
C515 VN.t4 VSUBS 0.220786f
C516 VN.n11 VSUBS 0.209607f
C517 VN.n12 VSUBS 0.052146f
C518 VN.n13 VSUBS 0.074297f
C519 VN.t0 VSUBS 0.125248f
C520 VN.n14 VSUBS 0.112396f
C521 VN.n15 VSUBS 0.291782f
C522 VN.t5 VSUBS 0.125248f
C523 VN.t1 VSUBS 0.284042f
C524 VN.n16 VSUBS 0.185619f
C525 VN.n17 VSUBS 0.201501f
C526 VN.n18 VSUBS 0.078718f
C527 VN.n19 VSUBS 0.078718f
C528 VN.n20 VSUBS 0.05568f
C529 VN.n21 VSUBS 0.05568f
C530 VN.n22 VSUBS 0.055099f
C531 VN.n23 VSUBS 0.070524f
C532 VN.t3 VSUBS 0.220786f
C533 VN.n24 VSUBS 0.209607f
C534 VN.n25 VSUBS 1.7902f
.ends

