* NGSPICE file created from diff_pair_sample_0437.ext - technology: sky130A

.subckt diff_pair_sample_0437 VTAIL VN VP B VDD2 VDD1
X0 B.t17 B.t15 B.t16 B.t9 sky130_fd_pr__nfet_01v8 ad=6.8211 pd=35.76 as=0 ps=0 w=17.49 l=1.36
X1 VTAIL.t7 VP.t0 VDD1.t0 B.t1 sky130_fd_pr__nfet_01v8 ad=6.8211 pd=35.76 as=2.88585 ps=17.82 w=17.49 l=1.36
X2 VTAIL.t3 VN.t0 VDD2.t3 B.t1 sky130_fd_pr__nfet_01v8 ad=6.8211 pd=35.76 as=2.88585 ps=17.82 w=17.49 l=1.36
X3 VDD2.t2 VN.t1 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=2.88585 pd=17.82 as=6.8211 ps=35.76 w=17.49 l=1.36
X4 VDD1.t1 VP.t1 VTAIL.t6 B.t2 sky130_fd_pr__nfet_01v8 ad=2.88585 pd=17.82 as=6.8211 ps=35.76 w=17.49 l=1.36
X5 VDD2.t1 VN.t2 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=2.88585 pd=17.82 as=6.8211 ps=35.76 w=17.49 l=1.36
X6 VTAIL.t5 VP.t2 VDD1.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=6.8211 pd=35.76 as=2.88585 ps=17.82 w=17.49 l=1.36
X7 VDD1.t2 VP.t3 VTAIL.t4 B.t0 sky130_fd_pr__nfet_01v8 ad=2.88585 pd=17.82 as=6.8211 ps=35.76 w=17.49 l=1.36
X8 B.t14 B.t12 B.t13 B.t5 sky130_fd_pr__nfet_01v8 ad=6.8211 pd=35.76 as=0 ps=0 w=17.49 l=1.36
X9 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=6.8211 pd=35.76 as=0 ps=0 w=17.49 l=1.36
X10 B.t7 B.t4 B.t6 B.t5 sky130_fd_pr__nfet_01v8 ad=6.8211 pd=35.76 as=0 ps=0 w=17.49 l=1.36
X11 VTAIL.t1 VN.t3 VDD2.t0 B.t3 sky130_fd_pr__nfet_01v8 ad=6.8211 pd=35.76 as=2.88585 ps=17.82 w=17.49 l=1.36
R0 B.n820 B.n819 585
R1 B.n821 B.n820 585
R2 B.n358 B.n108 585
R3 B.n357 B.n356 585
R4 B.n355 B.n354 585
R5 B.n353 B.n352 585
R6 B.n351 B.n350 585
R7 B.n349 B.n348 585
R8 B.n347 B.n346 585
R9 B.n345 B.n344 585
R10 B.n343 B.n342 585
R11 B.n341 B.n340 585
R12 B.n339 B.n338 585
R13 B.n337 B.n336 585
R14 B.n335 B.n334 585
R15 B.n333 B.n332 585
R16 B.n331 B.n330 585
R17 B.n329 B.n328 585
R18 B.n327 B.n326 585
R19 B.n325 B.n324 585
R20 B.n323 B.n322 585
R21 B.n321 B.n320 585
R22 B.n319 B.n318 585
R23 B.n317 B.n316 585
R24 B.n315 B.n314 585
R25 B.n313 B.n312 585
R26 B.n311 B.n310 585
R27 B.n309 B.n308 585
R28 B.n307 B.n306 585
R29 B.n305 B.n304 585
R30 B.n303 B.n302 585
R31 B.n301 B.n300 585
R32 B.n299 B.n298 585
R33 B.n297 B.n296 585
R34 B.n295 B.n294 585
R35 B.n293 B.n292 585
R36 B.n291 B.n290 585
R37 B.n289 B.n288 585
R38 B.n287 B.n286 585
R39 B.n285 B.n284 585
R40 B.n283 B.n282 585
R41 B.n281 B.n280 585
R42 B.n279 B.n278 585
R43 B.n277 B.n276 585
R44 B.n275 B.n274 585
R45 B.n273 B.n272 585
R46 B.n271 B.n270 585
R47 B.n269 B.n268 585
R48 B.n267 B.n266 585
R49 B.n265 B.n264 585
R50 B.n263 B.n262 585
R51 B.n261 B.n260 585
R52 B.n259 B.n258 585
R53 B.n257 B.n256 585
R54 B.n255 B.n254 585
R55 B.n253 B.n252 585
R56 B.n251 B.n250 585
R57 B.n249 B.n248 585
R58 B.n247 B.n246 585
R59 B.n244 B.n243 585
R60 B.n242 B.n241 585
R61 B.n240 B.n239 585
R62 B.n238 B.n237 585
R63 B.n236 B.n235 585
R64 B.n234 B.n233 585
R65 B.n232 B.n231 585
R66 B.n230 B.n229 585
R67 B.n228 B.n227 585
R68 B.n226 B.n225 585
R69 B.n224 B.n223 585
R70 B.n222 B.n221 585
R71 B.n220 B.n219 585
R72 B.n218 B.n217 585
R73 B.n216 B.n215 585
R74 B.n214 B.n213 585
R75 B.n212 B.n211 585
R76 B.n210 B.n209 585
R77 B.n208 B.n207 585
R78 B.n206 B.n205 585
R79 B.n204 B.n203 585
R80 B.n202 B.n201 585
R81 B.n200 B.n199 585
R82 B.n198 B.n197 585
R83 B.n196 B.n195 585
R84 B.n194 B.n193 585
R85 B.n192 B.n191 585
R86 B.n190 B.n189 585
R87 B.n188 B.n187 585
R88 B.n186 B.n185 585
R89 B.n184 B.n183 585
R90 B.n182 B.n181 585
R91 B.n180 B.n179 585
R92 B.n178 B.n177 585
R93 B.n176 B.n175 585
R94 B.n174 B.n173 585
R95 B.n172 B.n171 585
R96 B.n170 B.n169 585
R97 B.n168 B.n167 585
R98 B.n166 B.n165 585
R99 B.n164 B.n163 585
R100 B.n162 B.n161 585
R101 B.n160 B.n159 585
R102 B.n158 B.n157 585
R103 B.n156 B.n155 585
R104 B.n154 B.n153 585
R105 B.n152 B.n151 585
R106 B.n150 B.n149 585
R107 B.n148 B.n147 585
R108 B.n146 B.n145 585
R109 B.n144 B.n143 585
R110 B.n142 B.n141 585
R111 B.n140 B.n139 585
R112 B.n138 B.n137 585
R113 B.n136 B.n135 585
R114 B.n134 B.n133 585
R115 B.n132 B.n131 585
R116 B.n130 B.n129 585
R117 B.n128 B.n127 585
R118 B.n126 B.n125 585
R119 B.n124 B.n123 585
R120 B.n122 B.n121 585
R121 B.n120 B.n119 585
R122 B.n118 B.n117 585
R123 B.n116 B.n115 585
R124 B.n46 B.n45 585
R125 B.n824 B.n823 585
R126 B.n818 B.n109 585
R127 B.n109 B.n43 585
R128 B.n817 B.n42 585
R129 B.n828 B.n42 585
R130 B.n816 B.n41 585
R131 B.n829 B.n41 585
R132 B.n815 B.n40 585
R133 B.n830 B.n40 585
R134 B.n814 B.n813 585
R135 B.n813 B.n36 585
R136 B.n812 B.n35 585
R137 B.n836 B.n35 585
R138 B.n811 B.n34 585
R139 B.n837 B.n34 585
R140 B.n810 B.n33 585
R141 B.n838 B.n33 585
R142 B.n809 B.n808 585
R143 B.n808 B.n29 585
R144 B.n807 B.n28 585
R145 B.n844 B.n28 585
R146 B.n806 B.n27 585
R147 B.n845 B.n27 585
R148 B.n805 B.n26 585
R149 B.n846 B.n26 585
R150 B.n804 B.n803 585
R151 B.n803 B.n22 585
R152 B.n802 B.n21 585
R153 B.n852 B.n21 585
R154 B.n801 B.n20 585
R155 B.n853 B.n20 585
R156 B.n800 B.n19 585
R157 B.n854 B.n19 585
R158 B.n799 B.n798 585
R159 B.n798 B.n15 585
R160 B.n797 B.n14 585
R161 B.n860 B.n14 585
R162 B.n796 B.n13 585
R163 B.n861 B.n13 585
R164 B.n795 B.n12 585
R165 B.n862 B.n12 585
R166 B.n794 B.n793 585
R167 B.n793 B.n8 585
R168 B.n792 B.n7 585
R169 B.n868 B.n7 585
R170 B.n791 B.n6 585
R171 B.n869 B.n6 585
R172 B.n790 B.n5 585
R173 B.n870 B.n5 585
R174 B.n789 B.n788 585
R175 B.n788 B.n4 585
R176 B.n787 B.n359 585
R177 B.n787 B.n786 585
R178 B.n777 B.n360 585
R179 B.n361 B.n360 585
R180 B.n779 B.n778 585
R181 B.n780 B.n779 585
R182 B.n776 B.n365 585
R183 B.n369 B.n365 585
R184 B.n775 B.n774 585
R185 B.n774 B.n773 585
R186 B.n367 B.n366 585
R187 B.n368 B.n367 585
R188 B.n766 B.n765 585
R189 B.n767 B.n766 585
R190 B.n764 B.n374 585
R191 B.n374 B.n373 585
R192 B.n763 B.n762 585
R193 B.n762 B.n761 585
R194 B.n376 B.n375 585
R195 B.n377 B.n376 585
R196 B.n754 B.n753 585
R197 B.n755 B.n754 585
R198 B.n752 B.n382 585
R199 B.n382 B.n381 585
R200 B.n751 B.n750 585
R201 B.n750 B.n749 585
R202 B.n384 B.n383 585
R203 B.n385 B.n384 585
R204 B.n742 B.n741 585
R205 B.n743 B.n742 585
R206 B.n740 B.n390 585
R207 B.n390 B.n389 585
R208 B.n739 B.n738 585
R209 B.n738 B.n737 585
R210 B.n392 B.n391 585
R211 B.n393 B.n392 585
R212 B.n730 B.n729 585
R213 B.n731 B.n730 585
R214 B.n728 B.n398 585
R215 B.n398 B.n397 585
R216 B.n727 B.n726 585
R217 B.n726 B.n725 585
R218 B.n400 B.n399 585
R219 B.n401 B.n400 585
R220 B.n721 B.n720 585
R221 B.n404 B.n403 585
R222 B.n717 B.n716 585
R223 B.n718 B.n717 585
R224 B.n715 B.n466 585
R225 B.n714 B.n713 585
R226 B.n712 B.n711 585
R227 B.n710 B.n709 585
R228 B.n708 B.n707 585
R229 B.n706 B.n705 585
R230 B.n704 B.n703 585
R231 B.n702 B.n701 585
R232 B.n700 B.n699 585
R233 B.n698 B.n697 585
R234 B.n696 B.n695 585
R235 B.n694 B.n693 585
R236 B.n692 B.n691 585
R237 B.n690 B.n689 585
R238 B.n688 B.n687 585
R239 B.n686 B.n685 585
R240 B.n684 B.n683 585
R241 B.n682 B.n681 585
R242 B.n680 B.n679 585
R243 B.n678 B.n677 585
R244 B.n676 B.n675 585
R245 B.n674 B.n673 585
R246 B.n672 B.n671 585
R247 B.n670 B.n669 585
R248 B.n668 B.n667 585
R249 B.n666 B.n665 585
R250 B.n664 B.n663 585
R251 B.n662 B.n661 585
R252 B.n660 B.n659 585
R253 B.n658 B.n657 585
R254 B.n656 B.n655 585
R255 B.n654 B.n653 585
R256 B.n652 B.n651 585
R257 B.n650 B.n649 585
R258 B.n648 B.n647 585
R259 B.n646 B.n645 585
R260 B.n644 B.n643 585
R261 B.n642 B.n641 585
R262 B.n640 B.n639 585
R263 B.n638 B.n637 585
R264 B.n636 B.n635 585
R265 B.n634 B.n633 585
R266 B.n632 B.n631 585
R267 B.n630 B.n629 585
R268 B.n628 B.n627 585
R269 B.n626 B.n625 585
R270 B.n624 B.n623 585
R271 B.n622 B.n621 585
R272 B.n620 B.n619 585
R273 B.n618 B.n617 585
R274 B.n616 B.n615 585
R275 B.n614 B.n613 585
R276 B.n612 B.n611 585
R277 B.n610 B.n609 585
R278 B.n608 B.n607 585
R279 B.n605 B.n604 585
R280 B.n603 B.n602 585
R281 B.n601 B.n600 585
R282 B.n599 B.n598 585
R283 B.n597 B.n596 585
R284 B.n595 B.n594 585
R285 B.n593 B.n592 585
R286 B.n591 B.n590 585
R287 B.n589 B.n588 585
R288 B.n587 B.n586 585
R289 B.n585 B.n584 585
R290 B.n583 B.n582 585
R291 B.n581 B.n580 585
R292 B.n579 B.n578 585
R293 B.n577 B.n576 585
R294 B.n575 B.n574 585
R295 B.n573 B.n572 585
R296 B.n571 B.n570 585
R297 B.n569 B.n568 585
R298 B.n567 B.n566 585
R299 B.n565 B.n564 585
R300 B.n563 B.n562 585
R301 B.n561 B.n560 585
R302 B.n559 B.n558 585
R303 B.n557 B.n556 585
R304 B.n555 B.n554 585
R305 B.n553 B.n552 585
R306 B.n551 B.n550 585
R307 B.n549 B.n548 585
R308 B.n547 B.n546 585
R309 B.n545 B.n544 585
R310 B.n543 B.n542 585
R311 B.n541 B.n540 585
R312 B.n539 B.n538 585
R313 B.n537 B.n536 585
R314 B.n535 B.n534 585
R315 B.n533 B.n532 585
R316 B.n531 B.n530 585
R317 B.n529 B.n528 585
R318 B.n527 B.n526 585
R319 B.n525 B.n524 585
R320 B.n523 B.n522 585
R321 B.n521 B.n520 585
R322 B.n519 B.n518 585
R323 B.n517 B.n516 585
R324 B.n515 B.n514 585
R325 B.n513 B.n512 585
R326 B.n511 B.n510 585
R327 B.n509 B.n508 585
R328 B.n507 B.n506 585
R329 B.n505 B.n504 585
R330 B.n503 B.n502 585
R331 B.n501 B.n500 585
R332 B.n499 B.n498 585
R333 B.n497 B.n496 585
R334 B.n495 B.n494 585
R335 B.n493 B.n492 585
R336 B.n491 B.n490 585
R337 B.n489 B.n488 585
R338 B.n487 B.n486 585
R339 B.n485 B.n484 585
R340 B.n483 B.n482 585
R341 B.n481 B.n480 585
R342 B.n479 B.n478 585
R343 B.n477 B.n476 585
R344 B.n475 B.n474 585
R345 B.n473 B.n472 585
R346 B.n722 B.n402 585
R347 B.n402 B.n401 585
R348 B.n724 B.n723 585
R349 B.n725 B.n724 585
R350 B.n396 B.n395 585
R351 B.n397 B.n396 585
R352 B.n733 B.n732 585
R353 B.n732 B.n731 585
R354 B.n734 B.n394 585
R355 B.n394 B.n393 585
R356 B.n736 B.n735 585
R357 B.n737 B.n736 585
R358 B.n388 B.n387 585
R359 B.n389 B.n388 585
R360 B.n745 B.n744 585
R361 B.n744 B.n743 585
R362 B.n746 B.n386 585
R363 B.n386 B.n385 585
R364 B.n748 B.n747 585
R365 B.n749 B.n748 585
R366 B.n380 B.n379 585
R367 B.n381 B.n380 585
R368 B.n757 B.n756 585
R369 B.n756 B.n755 585
R370 B.n758 B.n378 585
R371 B.n378 B.n377 585
R372 B.n760 B.n759 585
R373 B.n761 B.n760 585
R374 B.n372 B.n371 585
R375 B.n373 B.n372 585
R376 B.n769 B.n768 585
R377 B.n768 B.n767 585
R378 B.n770 B.n370 585
R379 B.n370 B.n368 585
R380 B.n772 B.n771 585
R381 B.n773 B.n772 585
R382 B.n364 B.n363 585
R383 B.n369 B.n364 585
R384 B.n782 B.n781 585
R385 B.n781 B.n780 585
R386 B.n783 B.n362 585
R387 B.n362 B.n361 585
R388 B.n785 B.n784 585
R389 B.n786 B.n785 585
R390 B.n2 B.n0 585
R391 B.n4 B.n2 585
R392 B.n3 B.n1 585
R393 B.n869 B.n3 585
R394 B.n867 B.n866 585
R395 B.n868 B.n867 585
R396 B.n865 B.n9 585
R397 B.n9 B.n8 585
R398 B.n864 B.n863 585
R399 B.n863 B.n862 585
R400 B.n11 B.n10 585
R401 B.n861 B.n11 585
R402 B.n859 B.n858 585
R403 B.n860 B.n859 585
R404 B.n857 B.n16 585
R405 B.n16 B.n15 585
R406 B.n856 B.n855 585
R407 B.n855 B.n854 585
R408 B.n18 B.n17 585
R409 B.n853 B.n18 585
R410 B.n851 B.n850 585
R411 B.n852 B.n851 585
R412 B.n849 B.n23 585
R413 B.n23 B.n22 585
R414 B.n848 B.n847 585
R415 B.n847 B.n846 585
R416 B.n25 B.n24 585
R417 B.n845 B.n25 585
R418 B.n843 B.n842 585
R419 B.n844 B.n843 585
R420 B.n841 B.n30 585
R421 B.n30 B.n29 585
R422 B.n840 B.n839 585
R423 B.n839 B.n838 585
R424 B.n32 B.n31 585
R425 B.n837 B.n32 585
R426 B.n835 B.n834 585
R427 B.n836 B.n835 585
R428 B.n833 B.n37 585
R429 B.n37 B.n36 585
R430 B.n832 B.n831 585
R431 B.n831 B.n830 585
R432 B.n39 B.n38 585
R433 B.n829 B.n39 585
R434 B.n827 B.n826 585
R435 B.n828 B.n827 585
R436 B.n825 B.n44 585
R437 B.n44 B.n43 585
R438 B.n872 B.n871 585
R439 B.n871 B.n870 585
R440 B.n469 B.t12 514.811
R441 B.n467 B.t4 514.811
R442 B.n112 B.t8 514.811
R443 B.n110 B.t15 514.811
R444 B.n720 B.n402 511.721
R445 B.n823 B.n44 511.721
R446 B.n472 B.n400 511.721
R447 B.n820 B.n109 511.721
R448 B.n469 B.t14 409.452
R449 B.n110 B.t16 409.452
R450 B.n467 B.t7 409.452
R451 B.n112 B.t10 409.452
R452 B.n470 B.t13 376.678
R453 B.n111 B.t17 376.678
R454 B.n468 B.t6 376.678
R455 B.n113 B.t11 376.678
R456 B.n821 B.n107 256.663
R457 B.n821 B.n106 256.663
R458 B.n821 B.n105 256.663
R459 B.n821 B.n104 256.663
R460 B.n821 B.n103 256.663
R461 B.n821 B.n102 256.663
R462 B.n821 B.n101 256.663
R463 B.n821 B.n100 256.663
R464 B.n821 B.n99 256.663
R465 B.n821 B.n98 256.663
R466 B.n821 B.n97 256.663
R467 B.n821 B.n96 256.663
R468 B.n821 B.n95 256.663
R469 B.n821 B.n94 256.663
R470 B.n821 B.n93 256.663
R471 B.n821 B.n92 256.663
R472 B.n821 B.n91 256.663
R473 B.n821 B.n90 256.663
R474 B.n821 B.n89 256.663
R475 B.n821 B.n88 256.663
R476 B.n821 B.n87 256.663
R477 B.n821 B.n86 256.663
R478 B.n821 B.n85 256.663
R479 B.n821 B.n84 256.663
R480 B.n821 B.n83 256.663
R481 B.n821 B.n82 256.663
R482 B.n821 B.n81 256.663
R483 B.n821 B.n80 256.663
R484 B.n821 B.n79 256.663
R485 B.n821 B.n78 256.663
R486 B.n821 B.n77 256.663
R487 B.n821 B.n76 256.663
R488 B.n821 B.n75 256.663
R489 B.n821 B.n74 256.663
R490 B.n821 B.n73 256.663
R491 B.n821 B.n72 256.663
R492 B.n821 B.n71 256.663
R493 B.n821 B.n70 256.663
R494 B.n821 B.n69 256.663
R495 B.n821 B.n68 256.663
R496 B.n821 B.n67 256.663
R497 B.n821 B.n66 256.663
R498 B.n821 B.n65 256.663
R499 B.n821 B.n64 256.663
R500 B.n821 B.n63 256.663
R501 B.n821 B.n62 256.663
R502 B.n821 B.n61 256.663
R503 B.n821 B.n60 256.663
R504 B.n821 B.n59 256.663
R505 B.n821 B.n58 256.663
R506 B.n821 B.n57 256.663
R507 B.n821 B.n56 256.663
R508 B.n821 B.n55 256.663
R509 B.n821 B.n54 256.663
R510 B.n821 B.n53 256.663
R511 B.n821 B.n52 256.663
R512 B.n821 B.n51 256.663
R513 B.n821 B.n50 256.663
R514 B.n821 B.n49 256.663
R515 B.n821 B.n48 256.663
R516 B.n821 B.n47 256.663
R517 B.n822 B.n821 256.663
R518 B.n719 B.n718 256.663
R519 B.n718 B.n405 256.663
R520 B.n718 B.n406 256.663
R521 B.n718 B.n407 256.663
R522 B.n718 B.n408 256.663
R523 B.n718 B.n409 256.663
R524 B.n718 B.n410 256.663
R525 B.n718 B.n411 256.663
R526 B.n718 B.n412 256.663
R527 B.n718 B.n413 256.663
R528 B.n718 B.n414 256.663
R529 B.n718 B.n415 256.663
R530 B.n718 B.n416 256.663
R531 B.n718 B.n417 256.663
R532 B.n718 B.n418 256.663
R533 B.n718 B.n419 256.663
R534 B.n718 B.n420 256.663
R535 B.n718 B.n421 256.663
R536 B.n718 B.n422 256.663
R537 B.n718 B.n423 256.663
R538 B.n718 B.n424 256.663
R539 B.n718 B.n425 256.663
R540 B.n718 B.n426 256.663
R541 B.n718 B.n427 256.663
R542 B.n718 B.n428 256.663
R543 B.n718 B.n429 256.663
R544 B.n718 B.n430 256.663
R545 B.n718 B.n431 256.663
R546 B.n718 B.n432 256.663
R547 B.n718 B.n433 256.663
R548 B.n718 B.n434 256.663
R549 B.n718 B.n435 256.663
R550 B.n718 B.n436 256.663
R551 B.n718 B.n437 256.663
R552 B.n718 B.n438 256.663
R553 B.n718 B.n439 256.663
R554 B.n718 B.n440 256.663
R555 B.n718 B.n441 256.663
R556 B.n718 B.n442 256.663
R557 B.n718 B.n443 256.663
R558 B.n718 B.n444 256.663
R559 B.n718 B.n445 256.663
R560 B.n718 B.n446 256.663
R561 B.n718 B.n447 256.663
R562 B.n718 B.n448 256.663
R563 B.n718 B.n449 256.663
R564 B.n718 B.n450 256.663
R565 B.n718 B.n451 256.663
R566 B.n718 B.n452 256.663
R567 B.n718 B.n453 256.663
R568 B.n718 B.n454 256.663
R569 B.n718 B.n455 256.663
R570 B.n718 B.n456 256.663
R571 B.n718 B.n457 256.663
R572 B.n718 B.n458 256.663
R573 B.n718 B.n459 256.663
R574 B.n718 B.n460 256.663
R575 B.n718 B.n461 256.663
R576 B.n718 B.n462 256.663
R577 B.n718 B.n463 256.663
R578 B.n718 B.n464 256.663
R579 B.n718 B.n465 256.663
R580 B.n724 B.n402 163.367
R581 B.n724 B.n396 163.367
R582 B.n732 B.n396 163.367
R583 B.n732 B.n394 163.367
R584 B.n736 B.n394 163.367
R585 B.n736 B.n388 163.367
R586 B.n744 B.n388 163.367
R587 B.n744 B.n386 163.367
R588 B.n748 B.n386 163.367
R589 B.n748 B.n380 163.367
R590 B.n756 B.n380 163.367
R591 B.n756 B.n378 163.367
R592 B.n760 B.n378 163.367
R593 B.n760 B.n372 163.367
R594 B.n768 B.n372 163.367
R595 B.n768 B.n370 163.367
R596 B.n772 B.n370 163.367
R597 B.n772 B.n364 163.367
R598 B.n781 B.n364 163.367
R599 B.n781 B.n362 163.367
R600 B.n785 B.n362 163.367
R601 B.n785 B.n2 163.367
R602 B.n871 B.n2 163.367
R603 B.n871 B.n3 163.367
R604 B.n867 B.n3 163.367
R605 B.n867 B.n9 163.367
R606 B.n863 B.n9 163.367
R607 B.n863 B.n11 163.367
R608 B.n859 B.n11 163.367
R609 B.n859 B.n16 163.367
R610 B.n855 B.n16 163.367
R611 B.n855 B.n18 163.367
R612 B.n851 B.n18 163.367
R613 B.n851 B.n23 163.367
R614 B.n847 B.n23 163.367
R615 B.n847 B.n25 163.367
R616 B.n843 B.n25 163.367
R617 B.n843 B.n30 163.367
R618 B.n839 B.n30 163.367
R619 B.n839 B.n32 163.367
R620 B.n835 B.n32 163.367
R621 B.n835 B.n37 163.367
R622 B.n831 B.n37 163.367
R623 B.n831 B.n39 163.367
R624 B.n827 B.n39 163.367
R625 B.n827 B.n44 163.367
R626 B.n717 B.n404 163.367
R627 B.n717 B.n466 163.367
R628 B.n713 B.n712 163.367
R629 B.n709 B.n708 163.367
R630 B.n705 B.n704 163.367
R631 B.n701 B.n700 163.367
R632 B.n697 B.n696 163.367
R633 B.n693 B.n692 163.367
R634 B.n689 B.n688 163.367
R635 B.n685 B.n684 163.367
R636 B.n681 B.n680 163.367
R637 B.n677 B.n676 163.367
R638 B.n673 B.n672 163.367
R639 B.n669 B.n668 163.367
R640 B.n665 B.n664 163.367
R641 B.n661 B.n660 163.367
R642 B.n657 B.n656 163.367
R643 B.n653 B.n652 163.367
R644 B.n649 B.n648 163.367
R645 B.n645 B.n644 163.367
R646 B.n641 B.n640 163.367
R647 B.n637 B.n636 163.367
R648 B.n633 B.n632 163.367
R649 B.n629 B.n628 163.367
R650 B.n625 B.n624 163.367
R651 B.n621 B.n620 163.367
R652 B.n617 B.n616 163.367
R653 B.n613 B.n612 163.367
R654 B.n609 B.n608 163.367
R655 B.n604 B.n603 163.367
R656 B.n600 B.n599 163.367
R657 B.n596 B.n595 163.367
R658 B.n592 B.n591 163.367
R659 B.n588 B.n587 163.367
R660 B.n584 B.n583 163.367
R661 B.n580 B.n579 163.367
R662 B.n576 B.n575 163.367
R663 B.n572 B.n571 163.367
R664 B.n568 B.n567 163.367
R665 B.n564 B.n563 163.367
R666 B.n560 B.n559 163.367
R667 B.n556 B.n555 163.367
R668 B.n552 B.n551 163.367
R669 B.n548 B.n547 163.367
R670 B.n544 B.n543 163.367
R671 B.n540 B.n539 163.367
R672 B.n536 B.n535 163.367
R673 B.n532 B.n531 163.367
R674 B.n528 B.n527 163.367
R675 B.n524 B.n523 163.367
R676 B.n520 B.n519 163.367
R677 B.n516 B.n515 163.367
R678 B.n512 B.n511 163.367
R679 B.n508 B.n507 163.367
R680 B.n504 B.n503 163.367
R681 B.n500 B.n499 163.367
R682 B.n496 B.n495 163.367
R683 B.n492 B.n491 163.367
R684 B.n488 B.n487 163.367
R685 B.n484 B.n483 163.367
R686 B.n480 B.n479 163.367
R687 B.n476 B.n475 163.367
R688 B.n726 B.n400 163.367
R689 B.n726 B.n398 163.367
R690 B.n730 B.n398 163.367
R691 B.n730 B.n392 163.367
R692 B.n738 B.n392 163.367
R693 B.n738 B.n390 163.367
R694 B.n742 B.n390 163.367
R695 B.n742 B.n384 163.367
R696 B.n750 B.n384 163.367
R697 B.n750 B.n382 163.367
R698 B.n754 B.n382 163.367
R699 B.n754 B.n376 163.367
R700 B.n762 B.n376 163.367
R701 B.n762 B.n374 163.367
R702 B.n766 B.n374 163.367
R703 B.n766 B.n367 163.367
R704 B.n774 B.n367 163.367
R705 B.n774 B.n365 163.367
R706 B.n779 B.n365 163.367
R707 B.n779 B.n360 163.367
R708 B.n787 B.n360 163.367
R709 B.n788 B.n787 163.367
R710 B.n788 B.n5 163.367
R711 B.n6 B.n5 163.367
R712 B.n7 B.n6 163.367
R713 B.n793 B.n7 163.367
R714 B.n793 B.n12 163.367
R715 B.n13 B.n12 163.367
R716 B.n14 B.n13 163.367
R717 B.n798 B.n14 163.367
R718 B.n798 B.n19 163.367
R719 B.n20 B.n19 163.367
R720 B.n21 B.n20 163.367
R721 B.n803 B.n21 163.367
R722 B.n803 B.n26 163.367
R723 B.n27 B.n26 163.367
R724 B.n28 B.n27 163.367
R725 B.n808 B.n28 163.367
R726 B.n808 B.n33 163.367
R727 B.n34 B.n33 163.367
R728 B.n35 B.n34 163.367
R729 B.n813 B.n35 163.367
R730 B.n813 B.n40 163.367
R731 B.n41 B.n40 163.367
R732 B.n42 B.n41 163.367
R733 B.n109 B.n42 163.367
R734 B.n115 B.n46 163.367
R735 B.n119 B.n118 163.367
R736 B.n123 B.n122 163.367
R737 B.n127 B.n126 163.367
R738 B.n131 B.n130 163.367
R739 B.n135 B.n134 163.367
R740 B.n139 B.n138 163.367
R741 B.n143 B.n142 163.367
R742 B.n147 B.n146 163.367
R743 B.n151 B.n150 163.367
R744 B.n155 B.n154 163.367
R745 B.n159 B.n158 163.367
R746 B.n163 B.n162 163.367
R747 B.n167 B.n166 163.367
R748 B.n171 B.n170 163.367
R749 B.n175 B.n174 163.367
R750 B.n179 B.n178 163.367
R751 B.n183 B.n182 163.367
R752 B.n187 B.n186 163.367
R753 B.n191 B.n190 163.367
R754 B.n195 B.n194 163.367
R755 B.n199 B.n198 163.367
R756 B.n203 B.n202 163.367
R757 B.n207 B.n206 163.367
R758 B.n211 B.n210 163.367
R759 B.n215 B.n214 163.367
R760 B.n219 B.n218 163.367
R761 B.n223 B.n222 163.367
R762 B.n227 B.n226 163.367
R763 B.n231 B.n230 163.367
R764 B.n235 B.n234 163.367
R765 B.n239 B.n238 163.367
R766 B.n243 B.n242 163.367
R767 B.n248 B.n247 163.367
R768 B.n252 B.n251 163.367
R769 B.n256 B.n255 163.367
R770 B.n260 B.n259 163.367
R771 B.n264 B.n263 163.367
R772 B.n268 B.n267 163.367
R773 B.n272 B.n271 163.367
R774 B.n276 B.n275 163.367
R775 B.n280 B.n279 163.367
R776 B.n284 B.n283 163.367
R777 B.n288 B.n287 163.367
R778 B.n292 B.n291 163.367
R779 B.n296 B.n295 163.367
R780 B.n300 B.n299 163.367
R781 B.n304 B.n303 163.367
R782 B.n308 B.n307 163.367
R783 B.n312 B.n311 163.367
R784 B.n316 B.n315 163.367
R785 B.n320 B.n319 163.367
R786 B.n324 B.n323 163.367
R787 B.n328 B.n327 163.367
R788 B.n332 B.n331 163.367
R789 B.n336 B.n335 163.367
R790 B.n340 B.n339 163.367
R791 B.n344 B.n343 163.367
R792 B.n348 B.n347 163.367
R793 B.n352 B.n351 163.367
R794 B.n356 B.n355 163.367
R795 B.n820 B.n108 163.367
R796 B.n720 B.n719 71.676
R797 B.n466 B.n405 71.676
R798 B.n712 B.n406 71.676
R799 B.n708 B.n407 71.676
R800 B.n704 B.n408 71.676
R801 B.n700 B.n409 71.676
R802 B.n696 B.n410 71.676
R803 B.n692 B.n411 71.676
R804 B.n688 B.n412 71.676
R805 B.n684 B.n413 71.676
R806 B.n680 B.n414 71.676
R807 B.n676 B.n415 71.676
R808 B.n672 B.n416 71.676
R809 B.n668 B.n417 71.676
R810 B.n664 B.n418 71.676
R811 B.n660 B.n419 71.676
R812 B.n656 B.n420 71.676
R813 B.n652 B.n421 71.676
R814 B.n648 B.n422 71.676
R815 B.n644 B.n423 71.676
R816 B.n640 B.n424 71.676
R817 B.n636 B.n425 71.676
R818 B.n632 B.n426 71.676
R819 B.n628 B.n427 71.676
R820 B.n624 B.n428 71.676
R821 B.n620 B.n429 71.676
R822 B.n616 B.n430 71.676
R823 B.n612 B.n431 71.676
R824 B.n608 B.n432 71.676
R825 B.n603 B.n433 71.676
R826 B.n599 B.n434 71.676
R827 B.n595 B.n435 71.676
R828 B.n591 B.n436 71.676
R829 B.n587 B.n437 71.676
R830 B.n583 B.n438 71.676
R831 B.n579 B.n439 71.676
R832 B.n575 B.n440 71.676
R833 B.n571 B.n441 71.676
R834 B.n567 B.n442 71.676
R835 B.n563 B.n443 71.676
R836 B.n559 B.n444 71.676
R837 B.n555 B.n445 71.676
R838 B.n551 B.n446 71.676
R839 B.n547 B.n447 71.676
R840 B.n543 B.n448 71.676
R841 B.n539 B.n449 71.676
R842 B.n535 B.n450 71.676
R843 B.n531 B.n451 71.676
R844 B.n527 B.n452 71.676
R845 B.n523 B.n453 71.676
R846 B.n519 B.n454 71.676
R847 B.n515 B.n455 71.676
R848 B.n511 B.n456 71.676
R849 B.n507 B.n457 71.676
R850 B.n503 B.n458 71.676
R851 B.n499 B.n459 71.676
R852 B.n495 B.n460 71.676
R853 B.n491 B.n461 71.676
R854 B.n487 B.n462 71.676
R855 B.n483 B.n463 71.676
R856 B.n479 B.n464 71.676
R857 B.n475 B.n465 71.676
R858 B.n823 B.n822 71.676
R859 B.n115 B.n47 71.676
R860 B.n119 B.n48 71.676
R861 B.n123 B.n49 71.676
R862 B.n127 B.n50 71.676
R863 B.n131 B.n51 71.676
R864 B.n135 B.n52 71.676
R865 B.n139 B.n53 71.676
R866 B.n143 B.n54 71.676
R867 B.n147 B.n55 71.676
R868 B.n151 B.n56 71.676
R869 B.n155 B.n57 71.676
R870 B.n159 B.n58 71.676
R871 B.n163 B.n59 71.676
R872 B.n167 B.n60 71.676
R873 B.n171 B.n61 71.676
R874 B.n175 B.n62 71.676
R875 B.n179 B.n63 71.676
R876 B.n183 B.n64 71.676
R877 B.n187 B.n65 71.676
R878 B.n191 B.n66 71.676
R879 B.n195 B.n67 71.676
R880 B.n199 B.n68 71.676
R881 B.n203 B.n69 71.676
R882 B.n207 B.n70 71.676
R883 B.n211 B.n71 71.676
R884 B.n215 B.n72 71.676
R885 B.n219 B.n73 71.676
R886 B.n223 B.n74 71.676
R887 B.n227 B.n75 71.676
R888 B.n231 B.n76 71.676
R889 B.n235 B.n77 71.676
R890 B.n239 B.n78 71.676
R891 B.n243 B.n79 71.676
R892 B.n248 B.n80 71.676
R893 B.n252 B.n81 71.676
R894 B.n256 B.n82 71.676
R895 B.n260 B.n83 71.676
R896 B.n264 B.n84 71.676
R897 B.n268 B.n85 71.676
R898 B.n272 B.n86 71.676
R899 B.n276 B.n87 71.676
R900 B.n280 B.n88 71.676
R901 B.n284 B.n89 71.676
R902 B.n288 B.n90 71.676
R903 B.n292 B.n91 71.676
R904 B.n296 B.n92 71.676
R905 B.n300 B.n93 71.676
R906 B.n304 B.n94 71.676
R907 B.n308 B.n95 71.676
R908 B.n312 B.n96 71.676
R909 B.n316 B.n97 71.676
R910 B.n320 B.n98 71.676
R911 B.n324 B.n99 71.676
R912 B.n328 B.n100 71.676
R913 B.n332 B.n101 71.676
R914 B.n336 B.n102 71.676
R915 B.n340 B.n103 71.676
R916 B.n344 B.n104 71.676
R917 B.n348 B.n105 71.676
R918 B.n352 B.n106 71.676
R919 B.n356 B.n107 71.676
R920 B.n108 B.n107 71.676
R921 B.n355 B.n106 71.676
R922 B.n351 B.n105 71.676
R923 B.n347 B.n104 71.676
R924 B.n343 B.n103 71.676
R925 B.n339 B.n102 71.676
R926 B.n335 B.n101 71.676
R927 B.n331 B.n100 71.676
R928 B.n327 B.n99 71.676
R929 B.n323 B.n98 71.676
R930 B.n319 B.n97 71.676
R931 B.n315 B.n96 71.676
R932 B.n311 B.n95 71.676
R933 B.n307 B.n94 71.676
R934 B.n303 B.n93 71.676
R935 B.n299 B.n92 71.676
R936 B.n295 B.n91 71.676
R937 B.n291 B.n90 71.676
R938 B.n287 B.n89 71.676
R939 B.n283 B.n88 71.676
R940 B.n279 B.n87 71.676
R941 B.n275 B.n86 71.676
R942 B.n271 B.n85 71.676
R943 B.n267 B.n84 71.676
R944 B.n263 B.n83 71.676
R945 B.n259 B.n82 71.676
R946 B.n255 B.n81 71.676
R947 B.n251 B.n80 71.676
R948 B.n247 B.n79 71.676
R949 B.n242 B.n78 71.676
R950 B.n238 B.n77 71.676
R951 B.n234 B.n76 71.676
R952 B.n230 B.n75 71.676
R953 B.n226 B.n74 71.676
R954 B.n222 B.n73 71.676
R955 B.n218 B.n72 71.676
R956 B.n214 B.n71 71.676
R957 B.n210 B.n70 71.676
R958 B.n206 B.n69 71.676
R959 B.n202 B.n68 71.676
R960 B.n198 B.n67 71.676
R961 B.n194 B.n66 71.676
R962 B.n190 B.n65 71.676
R963 B.n186 B.n64 71.676
R964 B.n182 B.n63 71.676
R965 B.n178 B.n62 71.676
R966 B.n174 B.n61 71.676
R967 B.n170 B.n60 71.676
R968 B.n166 B.n59 71.676
R969 B.n162 B.n58 71.676
R970 B.n158 B.n57 71.676
R971 B.n154 B.n56 71.676
R972 B.n150 B.n55 71.676
R973 B.n146 B.n54 71.676
R974 B.n142 B.n53 71.676
R975 B.n138 B.n52 71.676
R976 B.n134 B.n51 71.676
R977 B.n130 B.n50 71.676
R978 B.n126 B.n49 71.676
R979 B.n122 B.n48 71.676
R980 B.n118 B.n47 71.676
R981 B.n822 B.n46 71.676
R982 B.n719 B.n404 71.676
R983 B.n713 B.n405 71.676
R984 B.n709 B.n406 71.676
R985 B.n705 B.n407 71.676
R986 B.n701 B.n408 71.676
R987 B.n697 B.n409 71.676
R988 B.n693 B.n410 71.676
R989 B.n689 B.n411 71.676
R990 B.n685 B.n412 71.676
R991 B.n681 B.n413 71.676
R992 B.n677 B.n414 71.676
R993 B.n673 B.n415 71.676
R994 B.n669 B.n416 71.676
R995 B.n665 B.n417 71.676
R996 B.n661 B.n418 71.676
R997 B.n657 B.n419 71.676
R998 B.n653 B.n420 71.676
R999 B.n649 B.n421 71.676
R1000 B.n645 B.n422 71.676
R1001 B.n641 B.n423 71.676
R1002 B.n637 B.n424 71.676
R1003 B.n633 B.n425 71.676
R1004 B.n629 B.n426 71.676
R1005 B.n625 B.n427 71.676
R1006 B.n621 B.n428 71.676
R1007 B.n617 B.n429 71.676
R1008 B.n613 B.n430 71.676
R1009 B.n609 B.n431 71.676
R1010 B.n604 B.n432 71.676
R1011 B.n600 B.n433 71.676
R1012 B.n596 B.n434 71.676
R1013 B.n592 B.n435 71.676
R1014 B.n588 B.n436 71.676
R1015 B.n584 B.n437 71.676
R1016 B.n580 B.n438 71.676
R1017 B.n576 B.n439 71.676
R1018 B.n572 B.n440 71.676
R1019 B.n568 B.n441 71.676
R1020 B.n564 B.n442 71.676
R1021 B.n560 B.n443 71.676
R1022 B.n556 B.n444 71.676
R1023 B.n552 B.n445 71.676
R1024 B.n548 B.n446 71.676
R1025 B.n544 B.n447 71.676
R1026 B.n540 B.n448 71.676
R1027 B.n536 B.n449 71.676
R1028 B.n532 B.n450 71.676
R1029 B.n528 B.n451 71.676
R1030 B.n524 B.n452 71.676
R1031 B.n520 B.n453 71.676
R1032 B.n516 B.n454 71.676
R1033 B.n512 B.n455 71.676
R1034 B.n508 B.n456 71.676
R1035 B.n504 B.n457 71.676
R1036 B.n500 B.n458 71.676
R1037 B.n496 B.n459 71.676
R1038 B.n492 B.n460 71.676
R1039 B.n488 B.n461 71.676
R1040 B.n484 B.n462 71.676
R1041 B.n480 B.n463 71.676
R1042 B.n476 B.n464 71.676
R1043 B.n472 B.n465 71.676
R1044 B.n718 B.n401 60.4002
R1045 B.n821 B.n43 60.4002
R1046 B.n471 B.n470 59.5399
R1047 B.n606 B.n468 59.5399
R1048 B.n114 B.n113 59.5399
R1049 B.n245 B.n111 59.5399
R1050 B.n825 B.n824 33.2493
R1051 B.n819 B.n818 33.2493
R1052 B.n473 B.n399 33.2493
R1053 B.n722 B.n721 33.2493
R1054 B.n725 B.n401 32.858
R1055 B.n725 B.n397 32.858
R1056 B.n731 B.n397 32.858
R1057 B.n731 B.n393 32.858
R1058 B.n737 B.n393 32.858
R1059 B.n743 B.n389 32.858
R1060 B.n743 B.n385 32.858
R1061 B.n749 B.n385 32.858
R1062 B.n749 B.n381 32.858
R1063 B.n755 B.n381 32.858
R1064 B.n755 B.n377 32.858
R1065 B.n761 B.n377 32.858
R1066 B.n767 B.n373 32.858
R1067 B.n767 B.n368 32.858
R1068 B.n773 B.n368 32.858
R1069 B.n773 B.n369 32.858
R1070 B.n780 B.n361 32.858
R1071 B.n786 B.n361 32.858
R1072 B.n786 B.n4 32.858
R1073 B.n870 B.n4 32.858
R1074 B.n870 B.n869 32.858
R1075 B.n869 B.n868 32.858
R1076 B.n868 B.n8 32.858
R1077 B.n862 B.n8 32.858
R1078 B.n861 B.n860 32.858
R1079 B.n860 B.n15 32.858
R1080 B.n854 B.n15 32.858
R1081 B.n854 B.n853 32.858
R1082 B.n852 B.n22 32.858
R1083 B.n846 B.n22 32.858
R1084 B.n846 B.n845 32.858
R1085 B.n845 B.n844 32.858
R1086 B.n844 B.n29 32.858
R1087 B.n838 B.n29 32.858
R1088 B.n838 B.n837 32.858
R1089 B.n836 B.n36 32.858
R1090 B.n830 B.n36 32.858
R1091 B.n830 B.n829 32.858
R1092 B.n829 B.n828 32.858
R1093 B.n828 B.n43 32.858
R1094 B.n470 B.n469 32.7763
R1095 B.n468 B.n467 32.7763
R1096 B.n113 B.n112 32.7763
R1097 B.n111 B.n110 32.7763
R1098 B.n761 B.t1 30.9252
R1099 B.t2 B.n852 30.9252
R1100 B.n369 B.t0 29.9588
R1101 B.t3 B.n861 29.9588
R1102 B.n737 B.t5 25.1268
R1103 B.t9 B.n836 25.1268
R1104 B B.n872 18.0485
R1105 B.n824 B.n45 10.6151
R1106 B.n116 B.n45 10.6151
R1107 B.n117 B.n116 10.6151
R1108 B.n120 B.n117 10.6151
R1109 B.n121 B.n120 10.6151
R1110 B.n124 B.n121 10.6151
R1111 B.n125 B.n124 10.6151
R1112 B.n128 B.n125 10.6151
R1113 B.n129 B.n128 10.6151
R1114 B.n132 B.n129 10.6151
R1115 B.n133 B.n132 10.6151
R1116 B.n136 B.n133 10.6151
R1117 B.n137 B.n136 10.6151
R1118 B.n140 B.n137 10.6151
R1119 B.n141 B.n140 10.6151
R1120 B.n144 B.n141 10.6151
R1121 B.n145 B.n144 10.6151
R1122 B.n148 B.n145 10.6151
R1123 B.n149 B.n148 10.6151
R1124 B.n152 B.n149 10.6151
R1125 B.n153 B.n152 10.6151
R1126 B.n156 B.n153 10.6151
R1127 B.n157 B.n156 10.6151
R1128 B.n160 B.n157 10.6151
R1129 B.n161 B.n160 10.6151
R1130 B.n164 B.n161 10.6151
R1131 B.n165 B.n164 10.6151
R1132 B.n168 B.n165 10.6151
R1133 B.n169 B.n168 10.6151
R1134 B.n172 B.n169 10.6151
R1135 B.n173 B.n172 10.6151
R1136 B.n176 B.n173 10.6151
R1137 B.n177 B.n176 10.6151
R1138 B.n180 B.n177 10.6151
R1139 B.n181 B.n180 10.6151
R1140 B.n184 B.n181 10.6151
R1141 B.n185 B.n184 10.6151
R1142 B.n188 B.n185 10.6151
R1143 B.n189 B.n188 10.6151
R1144 B.n192 B.n189 10.6151
R1145 B.n193 B.n192 10.6151
R1146 B.n196 B.n193 10.6151
R1147 B.n197 B.n196 10.6151
R1148 B.n200 B.n197 10.6151
R1149 B.n201 B.n200 10.6151
R1150 B.n204 B.n201 10.6151
R1151 B.n205 B.n204 10.6151
R1152 B.n208 B.n205 10.6151
R1153 B.n209 B.n208 10.6151
R1154 B.n212 B.n209 10.6151
R1155 B.n213 B.n212 10.6151
R1156 B.n216 B.n213 10.6151
R1157 B.n217 B.n216 10.6151
R1158 B.n220 B.n217 10.6151
R1159 B.n221 B.n220 10.6151
R1160 B.n224 B.n221 10.6151
R1161 B.n225 B.n224 10.6151
R1162 B.n229 B.n228 10.6151
R1163 B.n232 B.n229 10.6151
R1164 B.n233 B.n232 10.6151
R1165 B.n236 B.n233 10.6151
R1166 B.n237 B.n236 10.6151
R1167 B.n240 B.n237 10.6151
R1168 B.n241 B.n240 10.6151
R1169 B.n244 B.n241 10.6151
R1170 B.n249 B.n246 10.6151
R1171 B.n250 B.n249 10.6151
R1172 B.n253 B.n250 10.6151
R1173 B.n254 B.n253 10.6151
R1174 B.n257 B.n254 10.6151
R1175 B.n258 B.n257 10.6151
R1176 B.n261 B.n258 10.6151
R1177 B.n262 B.n261 10.6151
R1178 B.n265 B.n262 10.6151
R1179 B.n266 B.n265 10.6151
R1180 B.n269 B.n266 10.6151
R1181 B.n270 B.n269 10.6151
R1182 B.n273 B.n270 10.6151
R1183 B.n274 B.n273 10.6151
R1184 B.n277 B.n274 10.6151
R1185 B.n278 B.n277 10.6151
R1186 B.n281 B.n278 10.6151
R1187 B.n282 B.n281 10.6151
R1188 B.n285 B.n282 10.6151
R1189 B.n286 B.n285 10.6151
R1190 B.n289 B.n286 10.6151
R1191 B.n290 B.n289 10.6151
R1192 B.n293 B.n290 10.6151
R1193 B.n294 B.n293 10.6151
R1194 B.n297 B.n294 10.6151
R1195 B.n298 B.n297 10.6151
R1196 B.n301 B.n298 10.6151
R1197 B.n302 B.n301 10.6151
R1198 B.n305 B.n302 10.6151
R1199 B.n306 B.n305 10.6151
R1200 B.n309 B.n306 10.6151
R1201 B.n310 B.n309 10.6151
R1202 B.n313 B.n310 10.6151
R1203 B.n314 B.n313 10.6151
R1204 B.n317 B.n314 10.6151
R1205 B.n318 B.n317 10.6151
R1206 B.n321 B.n318 10.6151
R1207 B.n322 B.n321 10.6151
R1208 B.n325 B.n322 10.6151
R1209 B.n326 B.n325 10.6151
R1210 B.n329 B.n326 10.6151
R1211 B.n330 B.n329 10.6151
R1212 B.n333 B.n330 10.6151
R1213 B.n334 B.n333 10.6151
R1214 B.n337 B.n334 10.6151
R1215 B.n338 B.n337 10.6151
R1216 B.n341 B.n338 10.6151
R1217 B.n342 B.n341 10.6151
R1218 B.n345 B.n342 10.6151
R1219 B.n346 B.n345 10.6151
R1220 B.n349 B.n346 10.6151
R1221 B.n350 B.n349 10.6151
R1222 B.n353 B.n350 10.6151
R1223 B.n354 B.n353 10.6151
R1224 B.n357 B.n354 10.6151
R1225 B.n358 B.n357 10.6151
R1226 B.n819 B.n358 10.6151
R1227 B.n727 B.n399 10.6151
R1228 B.n728 B.n727 10.6151
R1229 B.n729 B.n728 10.6151
R1230 B.n729 B.n391 10.6151
R1231 B.n739 B.n391 10.6151
R1232 B.n740 B.n739 10.6151
R1233 B.n741 B.n740 10.6151
R1234 B.n741 B.n383 10.6151
R1235 B.n751 B.n383 10.6151
R1236 B.n752 B.n751 10.6151
R1237 B.n753 B.n752 10.6151
R1238 B.n753 B.n375 10.6151
R1239 B.n763 B.n375 10.6151
R1240 B.n764 B.n763 10.6151
R1241 B.n765 B.n764 10.6151
R1242 B.n765 B.n366 10.6151
R1243 B.n775 B.n366 10.6151
R1244 B.n776 B.n775 10.6151
R1245 B.n778 B.n776 10.6151
R1246 B.n778 B.n777 10.6151
R1247 B.n777 B.n359 10.6151
R1248 B.n789 B.n359 10.6151
R1249 B.n790 B.n789 10.6151
R1250 B.n791 B.n790 10.6151
R1251 B.n792 B.n791 10.6151
R1252 B.n794 B.n792 10.6151
R1253 B.n795 B.n794 10.6151
R1254 B.n796 B.n795 10.6151
R1255 B.n797 B.n796 10.6151
R1256 B.n799 B.n797 10.6151
R1257 B.n800 B.n799 10.6151
R1258 B.n801 B.n800 10.6151
R1259 B.n802 B.n801 10.6151
R1260 B.n804 B.n802 10.6151
R1261 B.n805 B.n804 10.6151
R1262 B.n806 B.n805 10.6151
R1263 B.n807 B.n806 10.6151
R1264 B.n809 B.n807 10.6151
R1265 B.n810 B.n809 10.6151
R1266 B.n811 B.n810 10.6151
R1267 B.n812 B.n811 10.6151
R1268 B.n814 B.n812 10.6151
R1269 B.n815 B.n814 10.6151
R1270 B.n816 B.n815 10.6151
R1271 B.n817 B.n816 10.6151
R1272 B.n818 B.n817 10.6151
R1273 B.n721 B.n403 10.6151
R1274 B.n716 B.n403 10.6151
R1275 B.n716 B.n715 10.6151
R1276 B.n715 B.n714 10.6151
R1277 B.n714 B.n711 10.6151
R1278 B.n711 B.n710 10.6151
R1279 B.n710 B.n707 10.6151
R1280 B.n707 B.n706 10.6151
R1281 B.n706 B.n703 10.6151
R1282 B.n703 B.n702 10.6151
R1283 B.n702 B.n699 10.6151
R1284 B.n699 B.n698 10.6151
R1285 B.n698 B.n695 10.6151
R1286 B.n695 B.n694 10.6151
R1287 B.n694 B.n691 10.6151
R1288 B.n691 B.n690 10.6151
R1289 B.n690 B.n687 10.6151
R1290 B.n687 B.n686 10.6151
R1291 B.n686 B.n683 10.6151
R1292 B.n683 B.n682 10.6151
R1293 B.n682 B.n679 10.6151
R1294 B.n679 B.n678 10.6151
R1295 B.n678 B.n675 10.6151
R1296 B.n675 B.n674 10.6151
R1297 B.n674 B.n671 10.6151
R1298 B.n671 B.n670 10.6151
R1299 B.n670 B.n667 10.6151
R1300 B.n667 B.n666 10.6151
R1301 B.n666 B.n663 10.6151
R1302 B.n663 B.n662 10.6151
R1303 B.n662 B.n659 10.6151
R1304 B.n659 B.n658 10.6151
R1305 B.n658 B.n655 10.6151
R1306 B.n655 B.n654 10.6151
R1307 B.n654 B.n651 10.6151
R1308 B.n651 B.n650 10.6151
R1309 B.n650 B.n647 10.6151
R1310 B.n647 B.n646 10.6151
R1311 B.n646 B.n643 10.6151
R1312 B.n643 B.n642 10.6151
R1313 B.n642 B.n639 10.6151
R1314 B.n639 B.n638 10.6151
R1315 B.n638 B.n635 10.6151
R1316 B.n635 B.n634 10.6151
R1317 B.n634 B.n631 10.6151
R1318 B.n631 B.n630 10.6151
R1319 B.n630 B.n627 10.6151
R1320 B.n627 B.n626 10.6151
R1321 B.n626 B.n623 10.6151
R1322 B.n623 B.n622 10.6151
R1323 B.n622 B.n619 10.6151
R1324 B.n619 B.n618 10.6151
R1325 B.n618 B.n615 10.6151
R1326 B.n615 B.n614 10.6151
R1327 B.n614 B.n611 10.6151
R1328 B.n611 B.n610 10.6151
R1329 B.n610 B.n607 10.6151
R1330 B.n605 B.n602 10.6151
R1331 B.n602 B.n601 10.6151
R1332 B.n601 B.n598 10.6151
R1333 B.n598 B.n597 10.6151
R1334 B.n597 B.n594 10.6151
R1335 B.n594 B.n593 10.6151
R1336 B.n593 B.n590 10.6151
R1337 B.n590 B.n589 10.6151
R1338 B.n586 B.n585 10.6151
R1339 B.n585 B.n582 10.6151
R1340 B.n582 B.n581 10.6151
R1341 B.n581 B.n578 10.6151
R1342 B.n578 B.n577 10.6151
R1343 B.n577 B.n574 10.6151
R1344 B.n574 B.n573 10.6151
R1345 B.n573 B.n570 10.6151
R1346 B.n570 B.n569 10.6151
R1347 B.n569 B.n566 10.6151
R1348 B.n566 B.n565 10.6151
R1349 B.n565 B.n562 10.6151
R1350 B.n562 B.n561 10.6151
R1351 B.n561 B.n558 10.6151
R1352 B.n558 B.n557 10.6151
R1353 B.n557 B.n554 10.6151
R1354 B.n554 B.n553 10.6151
R1355 B.n553 B.n550 10.6151
R1356 B.n550 B.n549 10.6151
R1357 B.n549 B.n546 10.6151
R1358 B.n546 B.n545 10.6151
R1359 B.n545 B.n542 10.6151
R1360 B.n542 B.n541 10.6151
R1361 B.n541 B.n538 10.6151
R1362 B.n538 B.n537 10.6151
R1363 B.n537 B.n534 10.6151
R1364 B.n534 B.n533 10.6151
R1365 B.n533 B.n530 10.6151
R1366 B.n530 B.n529 10.6151
R1367 B.n529 B.n526 10.6151
R1368 B.n526 B.n525 10.6151
R1369 B.n525 B.n522 10.6151
R1370 B.n522 B.n521 10.6151
R1371 B.n521 B.n518 10.6151
R1372 B.n518 B.n517 10.6151
R1373 B.n517 B.n514 10.6151
R1374 B.n514 B.n513 10.6151
R1375 B.n513 B.n510 10.6151
R1376 B.n510 B.n509 10.6151
R1377 B.n509 B.n506 10.6151
R1378 B.n506 B.n505 10.6151
R1379 B.n505 B.n502 10.6151
R1380 B.n502 B.n501 10.6151
R1381 B.n501 B.n498 10.6151
R1382 B.n498 B.n497 10.6151
R1383 B.n497 B.n494 10.6151
R1384 B.n494 B.n493 10.6151
R1385 B.n493 B.n490 10.6151
R1386 B.n490 B.n489 10.6151
R1387 B.n489 B.n486 10.6151
R1388 B.n486 B.n485 10.6151
R1389 B.n485 B.n482 10.6151
R1390 B.n482 B.n481 10.6151
R1391 B.n481 B.n478 10.6151
R1392 B.n478 B.n477 10.6151
R1393 B.n477 B.n474 10.6151
R1394 B.n474 B.n473 10.6151
R1395 B.n723 B.n722 10.6151
R1396 B.n723 B.n395 10.6151
R1397 B.n733 B.n395 10.6151
R1398 B.n734 B.n733 10.6151
R1399 B.n735 B.n734 10.6151
R1400 B.n735 B.n387 10.6151
R1401 B.n745 B.n387 10.6151
R1402 B.n746 B.n745 10.6151
R1403 B.n747 B.n746 10.6151
R1404 B.n747 B.n379 10.6151
R1405 B.n757 B.n379 10.6151
R1406 B.n758 B.n757 10.6151
R1407 B.n759 B.n758 10.6151
R1408 B.n759 B.n371 10.6151
R1409 B.n769 B.n371 10.6151
R1410 B.n770 B.n769 10.6151
R1411 B.n771 B.n770 10.6151
R1412 B.n771 B.n363 10.6151
R1413 B.n782 B.n363 10.6151
R1414 B.n783 B.n782 10.6151
R1415 B.n784 B.n783 10.6151
R1416 B.n784 B.n0 10.6151
R1417 B.n866 B.n1 10.6151
R1418 B.n866 B.n865 10.6151
R1419 B.n865 B.n864 10.6151
R1420 B.n864 B.n10 10.6151
R1421 B.n858 B.n10 10.6151
R1422 B.n858 B.n857 10.6151
R1423 B.n857 B.n856 10.6151
R1424 B.n856 B.n17 10.6151
R1425 B.n850 B.n17 10.6151
R1426 B.n850 B.n849 10.6151
R1427 B.n849 B.n848 10.6151
R1428 B.n848 B.n24 10.6151
R1429 B.n842 B.n24 10.6151
R1430 B.n842 B.n841 10.6151
R1431 B.n841 B.n840 10.6151
R1432 B.n840 B.n31 10.6151
R1433 B.n834 B.n31 10.6151
R1434 B.n834 B.n833 10.6151
R1435 B.n833 B.n832 10.6151
R1436 B.n832 B.n38 10.6151
R1437 B.n826 B.n38 10.6151
R1438 B.n826 B.n825 10.6151
R1439 B.t5 B.n389 7.73167
R1440 B.n837 B.t9 7.73167
R1441 B.n228 B.n114 6.5566
R1442 B.n245 B.n244 6.5566
R1443 B.n606 B.n605 6.5566
R1444 B.n589 B.n471 6.5566
R1445 B.n225 B.n114 4.05904
R1446 B.n246 B.n245 4.05904
R1447 B.n607 B.n606 4.05904
R1448 B.n586 B.n471 4.05904
R1449 B.n780 B.t0 2.89969
R1450 B.n862 B.t3 2.89969
R1451 B.n872 B.n0 2.81026
R1452 B.n872 B.n1 2.81026
R1453 B.t1 B.n373 1.93329
R1454 B.n853 B.t2 1.93329
R1455 VP.n2 VP.t2 348.219
R1456 VP.n2 VP.t1 347.986
R1457 VP.n3 VP.t0 309.933
R1458 VP.n9 VP.t3 309.933
R1459 VP.n4 VP.n3 168.886
R1460 VP.n10 VP.n9 168.886
R1461 VP.n8 VP.n0 161.3
R1462 VP.n7 VP.n6 161.3
R1463 VP.n5 VP.n1 161.3
R1464 VP.n4 VP.n2 64.328
R1465 VP.n7 VP.n1 40.4934
R1466 VP.n8 VP.n7 40.4934
R1467 VP.n3 VP.n1 16.8827
R1468 VP.n9 VP.n8 16.8827
R1469 VP.n5 VP.n4 0.189894
R1470 VP.n6 VP.n5 0.189894
R1471 VP.n6 VP.n0 0.189894
R1472 VP.n10 VP.n0 0.189894
R1473 VP VP.n10 0.0516364
R1474 VDD1 VDD1.n1 103.788
R1475 VDD1 VDD1.n0 60.1583
R1476 VDD1.n0 VDD1.t3 1.13258
R1477 VDD1.n0 VDD1.t1 1.13258
R1478 VDD1.n1 VDD1.t0 1.13258
R1479 VDD1.n1 VDD1.t2 1.13258
R1480 VTAIL.n778 VTAIL.n686 289.615
R1481 VTAIL.n92 VTAIL.n0 289.615
R1482 VTAIL.n190 VTAIL.n98 289.615
R1483 VTAIL.n288 VTAIL.n196 289.615
R1484 VTAIL.n680 VTAIL.n588 289.615
R1485 VTAIL.n582 VTAIL.n490 289.615
R1486 VTAIL.n484 VTAIL.n392 289.615
R1487 VTAIL.n386 VTAIL.n294 289.615
R1488 VTAIL.n719 VTAIL.n718 185
R1489 VTAIL.n721 VTAIL.n720 185
R1490 VTAIL.n714 VTAIL.n713 185
R1491 VTAIL.n727 VTAIL.n726 185
R1492 VTAIL.n729 VTAIL.n728 185
R1493 VTAIL.n710 VTAIL.n709 185
R1494 VTAIL.n735 VTAIL.n734 185
R1495 VTAIL.n737 VTAIL.n736 185
R1496 VTAIL.n706 VTAIL.n705 185
R1497 VTAIL.n743 VTAIL.n742 185
R1498 VTAIL.n745 VTAIL.n744 185
R1499 VTAIL.n702 VTAIL.n701 185
R1500 VTAIL.n751 VTAIL.n750 185
R1501 VTAIL.n753 VTAIL.n752 185
R1502 VTAIL.n698 VTAIL.n697 185
R1503 VTAIL.n760 VTAIL.n759 185
R1504 VTAIL.n761 VTAIL.n696 185
R1505 VTAIL.n763 VTAIL.n762 185
R1506 VTAIL.n694 VTAIL.n693 185
R1507 VTAIL.n769 VTAIL.n768 185
R1508 VTAIL.n771 VTAIL.n770 185
R1509 VTAIL.n690 VTAIL.n689 185
R1510 VTAIL.n777 VTAIL.n776 185
R1511 VTAIL.n779 VTAIL.n778 185
R1512 VTAIL.n33 VTAIL.n32 185
R1513 VTAIL.n35 VTAIL.n34 185
R1514 VTAIL.n28 VTAIL.n27 185
R1515 VTAIL.n41 VTAIL.n40 185
R1516 VTAIL.n43 VTAIL.n42 185
R1517 VTAIL.n24 VTAIL.n23 185
R1518 VTAIL.n49 VTAIL.n48 185
R1519 VTAIL.n51 VTAIL.n50 185
R1520 VTAIL.n20 VTAIL.n19 185
R1521 VTAIL.n57 VTAIL.n56 185
R1522 VTAIL.n59 VTAIL.n58 185
R1523 VTAIL.n16 VTAIL.n15 185
R1524 VTAIL.n65 VTAIL.n64 185
R1525 VTAIL.n67 VTAIL.n66 185
R1526 VTAIL.n12 VTAIL.n11 185
R1527 VTAIL.n74 VTAIL.n73 185
R1528 VTAIL.n75 VTAIL.n10 185
R1529 VTAIL.n77 VTAIL.n76 185
R1530 VTAIL.n8 VTAIL.n7 185
R1531 VTAIL.n83 VTAIL.n82 185
R1532 VTAIL.n85 VTAIL.n84 185
R1533 VTAIL.n4 VTAIL.n3 185
R1534 VTAIL.n91 VTAIL.n90 185
R1535 VTAIL.n93 VTAIL.n92 185
R1536 VTAIL.n131 VTAIL.n130 185
R1537 VTAIL.n133 VTAIL.n132 185
R1538 VTAIL.n126 VTAIL.n125 185
R1539 VTAIL.n139 VTAIL.n138 185
R1540 VTAIL.n141 VTAIL.n140 185
R1541 VTAIL.n122 VTAIL.n121 185
R1542 VTAIL.n147 VTAIL.n146 185
R1543 VTAIL.n149 VTAIL.n148 185
R1544 VTAIL.n118 VTAIL.n117 185
R1545 VTAIL.n155 VTAIL.n154 185
R1546 VTAIL.n157 VTAIL.n156 185
R1547 VTAIL.n114 VTAIL.n113 185
R1548 VTAIL.n163 VTAIL.n162 185
R1549 VTAIL.n165 VTAIL.n164 185
R1550 VTAIL.n110 VTAIL.n109 185
R1551 VTAIL.n172 VTAIL.n171 185
R1552 VTAIL.n173 VTAIL.n108 185
R1553 VTAIL.n175 VTAIL.n174 185
R1554 VTAIL.n106 VTAIL.n105 185
R1555 VTAIL.n181 VTAIL.n180 185
R1556 VTAIL.n183 VTAIL.n182 185
R1557 VTAIL.n102 VTAIL.n101 185
R1558 VTAIL.n189 VTAIL.n188 185
R1559 VTAIL.n191 VTAIL.n190 185
R1560 VTAIL.n229 VTAIL.n228 185
R1561 VTAIL.n231 VTAIL.n230 185
R1562 VTAIL.n224 VTAIL.n223 185
R1563 VTAIL.n237 VTAIL.n236 185
R1564 VTAIL.n239 VTAIL.n238 185
R1565 VTAIL.n220 VTAIL.n219 185
R1566 VTAIL.n245 VTAIL.n244 185
R1567 VTAIL.n247 VTAIL.n246 185
R1568 VTAIL.n216 VTAIL.n215 185
R1569 VTAIL.n253 VTAIL.n252 185
R1570 VTAIL.n255 VTAIL.n254 185
R1571 VTAIL.n212 VTAIL.n211 185
R1572 VTAIL.n261 VTAIL.n260 185
R1573 VTAIL.n263 VTAIL.n262 185
R1574 VTAIL.n208 VTAIL.n207 185
R1575 VTAIL.n270 VTAIL.n269 185
R1576 VTAIL.n271 VTAIL.n206 185
R1577 VTAIL.n273 VTAIL.n272 185
R1578 VTAIL.n204 VTAIL.n203 185
R1579 VTAIL.n279 VTAIL.n278 185
R1580 VTAIL.n281 VTAIL.n280 185
R1581 VTAIL.n200 VTAIL.n199 185
R1582 VTAIL.n287 VTAIL.n286 185
R1583 VTAIL.n289 VTAIL.n288 185
R1584 VTAIL.n681 VTAIL.n680 185
R1585 VTAIL.n679 VTAIL.n678 185
R1586 VTAIL.n592 VTAIL.n591 185
R1587 VTAIL.n673 VTAIL.n672 185
R1588 VTAIL.n671 VTAIL.n670 185
R1589 VTAIL.n596 VTAIL.n595 185
R1590 VTAIL.n600 VTAIL.n598 185
R1591 VTAIL.n665 VTAIL.n664 185
R1592 VTAIL.n663 VTAIL.n662 185
R1593 VTAIL.n602 VTAIL.n601 185
R1594 VTAIL.n657 VTAIL.n656 185
R1595 VTAIL.n655 VTAIL.n654 185
R1596 VTAIL.n606 VTAIL.n605 185
R1597 VTAIL.n649 VTAIL.n648 185
R1598 VTAIL.n647 VTAIL.n646 185
R1599 VTAIL.n610 VTAIL.n609 185
R1600 VTAIL.n641 VTAIL.n640 185
R1601 VTAIL.n639 VTAIL.n638 185
R1602 VTAIL.n614 VTAIL.n613 185
R1603 VTAIL.n633 VTAIL.n632 185
R1604 VTAIL.n631 VTAIL.n630 185
R1605 VTAIL.n618 VTAIL.n617 185
R1606 VTAIL.n625 VTAIL.n624 185
R1607 VTAIL.n623 VTAIL.n622 185
R1608 VTAIL.n583 VTAIL.n582 185
R1609 VTAIL.n581 VTAIL.n580 185
R1610 VTAIL.n494 VTAIL.n493 185
R1611 VTAIL.n575 VTAIL.n574 185
R1612 VTAIL.n573 VTAIL.n572 185
R1613 VTAIL.n498 VTAIL.n497 185
R1614 VTAIL.n502 VTAIL.n500 185
R1615 VTAIL.n567 VTAIL.n566 185
R1616 VTAIL.n565 VTAIL.n564 185
R1617 VTAIL.n504 VTAIL.n503 185
R1618 VTAIL.n559 VTAIL.n558 185
R1619 VTAIL.n557 VTAIL.n556 185
R1620 VTAIL.n508 VTAIL.n507 185
R1621 VTAIL.n551 VTAIL.n550 185
R1622 VTAIL.n549 VTAIL.n548 185
R1623 VTAIL.n512 VTAIL.n511 185
R1624 VTAIL.n543 VTAIL.n542 185
R1625 VTAIL.n541 VTAIL.n540 185
R1626 VTAIL.n516 VTAIL.n515 185
R1627 VTAIL.n535 VTAIL.n534 185
R1628 VTAIL.n533 VTAIL.n532 185
R1629 VTAIL.n520 VTAIL.n519 185
R1630 VTAIL.n527 VTAIL.n526 185
R1631 VTAIL.n525 VTAIL.n524 185
R1632 VTAIL.n485 VTAIL.n484 185
R1633 VTAIL.n483 VTAIL.n482 185
R1634 VTAIL.n396 VTAIL.n395 185
R1635 VTAIL.n477 VTAIL.n476 185
R1636 VTAIL.n475 VTAIL.n474 185
R1637 VTAIL.n400 VTAIL.n399 185
R1638 VTAIL.n404 VTAIL.n402 185
R1639 VTAIL.n469 VTAIL.n468 185
R1640 VTAIL.n467 VTAIL.n466 185
R1641 VTAIL.n406 VTAIL.n405 185
R1642 VTAIL.n461 VTAIL.n460 185
R1643 VTAIL.n459 VTAIL.n458 185
R1644 VTAIL.n410 VTAIL.n409 185
R1645 VTAIL.n453 VTAIL.n452 185
R1646 VTAIL.n451 VTAIL.n450 185
R1647 VTAIL.n414 VTAIL.n413 185
R1648 VTAIL.n445 VTAIL.n444 185
R1649 VTAIL.n443 VTAIL.n442 185
R1650 VTAIL.n418 VTAIL.n417 185
R1651 VTAIL.n437 VTAIL.n436 185
R1652 VTAIL.n435 VTAIL.n434 185
R1653 VTAIL.n422 VTAIL.n421 185
R1654 VTAIL.n429 VTAIL.n428 185
R1655 VTAIL.n427 VTAIL.n426 185
R1656 VTAIL.n387 VTAIL.n386 185
R1657 VTAIL.n385 VTAIL.n384 185
R1658 VTAIL.n298 VTAIL.n297 185
R1659 VTAIL.n379 VTAIL.n378 185
R1660 VTAIL.n377 VTAIL.n376 185
R1661 VTAIL.n302 VTAIL.n301 185
R1662 VTAIL.n306 VTAIL.n304 185
R1663 VTAIL.n371 VTAIL.n370 185
R1664 VTAIL.n369 VTAIL.n368 185
R1665 VTAIL.n308 VTAIL.n307 185
R1666 VTAIL.n363 VTAIL.n362 185
R1667 VTAIL.n361 VTAIL.n360 185
R1668 VTAIL.n312 VTAIL.n311 185
R1669 VTAIL.n355 VTAIL.n354 185
R1670 VTAIL.n353 VTAIL.n352 185
R1671 VTAIL.n316 VTAIL.n315 185
R1672 VTAIL.n347 VTAIL.n346 185
R1673 VTAIL.n345 VTAIL.n344 185
R1674 VTAIL.n320 VTAIL.n319 185
R1675 VTAIL.n339 VTAIL.n338 185
R1676 VTAIL.n337 VTAIL.n336 185
R1677 VTAIL.n324 VTAIL.n323 185
R1678 VTAIL.n331 VTAIL.n330 185
R1679 VTAIL.n329 VTAIL.n328 185
R1680 VTAIL.n717 VTAIL.t2 147.659
R1681 VTAIL.n31 VTAIL.t1 147.659
R1682 VTAIL.n129 VTAIL.t4 147.659
R1683 VTAIL.n227 VTAIL.t7 147.659
R1684 VTAIL.n621 VTAIL.t6 147.659
R1685 VTAIL.n523 VTAIL.t5 147.659
R1686 VTAIL.n425 VTAIL.t0 147.659
R1687 VTAIL.n327 VTAIL.t3 147.659
R1688 VTAIL.n720 VTAIL.n719 104.615
R1689 VTAIL.n720 VTAIL.n713 104.615
R1690 VTAIL.n727 VTAIL.n713 104.615
R1691 VTAIL.n728 VTAIL.n727 104.615
R1692 VTAIL.n728 VTAIL.n709 104.615
R1693 VTAIL.n735 VTAIL.n709 104.615
R1694 VTAIL.n736 VTAIL.n735 104.615
R1695 VTAIL.n736 VTAIL.n705 104.615
R1696 VTAIL.n743 VTAIL.n705 104.615
R1697 VTAIL.n744 VTAIL.n743 104.615
R1698 VTAIL.n744 VTAIL.n701 104.615
R1699 VTAIL.n751 VTAIL.n701 104.615
R1700 VTAIL.n752 VTAIL.n751 104.615
R1701 VTAIL.n752 VTAIL.n697 104.615
R1702 VTAIL.n760 VTAIL.n697 104.615
R1703 VTAIL.n761 VTAIL.n760 104.615
R1704 VTAIL.n762 VTAIL.n761 104.615
R1705 VTAIL.n762 VTAIL.n693 104.615
R1706 VTAIL.n769 VTAIL.n693 104.615
R1707 VTAIL.n770 VTAIL.n769 104.615
R1708 VTAIL.n770 VTAIL.n689 104.615
R1709 VTAIL.n777 VTAIL.n689 104.615
R1710 VTAIL.n778 VTAIL.n777 104.615
R1711 VTAIL.n34 VTAIL.n33 104.615
R1712 VTAIL.n34 VTAIL.n27 104.615
R1713 VTAIL.n41 VTAIL.n27 104.615
R1714 VTAIL.n42 VTAIL.n41 104.615
R1715 VTAIL.n42 VTAIL.n23 104.615
R1716 VTAIL.n49 VTAIL.n23 104.615
R1717 VTAIL.n50 VTAIL.n49 104.615
R1718 VTAIL.n50 VTAIL.n19 104.615
R1719 VTAIL.n57 VTAIL.n19 104.615
R1720 VTAIL.n58 VTAIL.n57 104.615
R1721 VTAIL.n58 VTAIL.n15 104.615
R1722 VTAIL.n65 VTAIL.n15 104.615
R1723 VTAIL.n66 VTAIL.n65 104.615
R1724 VTAIL.n66 VTAIL.n11 104.615
R1725 VTAIL.n74 VTAIL.n11 104.615
R1726 VTAIL.n75 VTAIL.n74 104.615
R1727 VTAIL.n76 VTAIL.n75 104.615
R1728 VTAIL.n76 VTAIL.n7 104.615
R1729 VTAIL.n83 VTAIL.n7 104.615
R1730 VTAIL.n84 VTAIL.n83 104.615
R1731 VTAIL.n84 VTAIL.n3 104.615
R1732 VTAIL.n91 VTAIL.n3 104.615
R1733 VTAIL.n92 VTAIL.n91 104.615
R1734 VTAIL.n132 VTAIL.n131 104.615
R1735 VTAIL.n132 VTAIL.n125 104.615
R1736 VTAIL.n139 VTAIL.n125 104.615
R1737 VTAIL.n140 VTAIL.n139 104.615
R1738 VTAIL.n140 VTAIL.n121 104.615
R1739 VTAIL.n147 VTAIL.n121 104.615
R1740 VTAIL.n148 VTAIL.n147 104.615
R1741 VTAIL.n148 VTAIL.n117 104.615
R1742 VTAIL.n155 VTAIL.n117 104.615
R1743 VTAIL.n156 VTAIL.n155 104.615
R1744 VTAIL.n156 VTAIL.n113 104.615
R1745 VTAIL.n163 VTAIL.n113 104.615
R1746 VTAIL.n164 VTAIL.n163 104.615
R1747 VTAIL.n164 VTAIL.n109 104.615
R1748 VTAIL.n172 VTAIL.n109 104.615
R1749 VTAIL.n173 VTAIL.n172 104.615
R1750 VTAIL.n174 VTAIL.n173 104.615
R1751 VTAIL.n174 VTAIL.n105 104.615
R1752 VTAIL.n181 VTAIL.n105 104.615
R1753 VTAIL.n182 VTAIL.n181 104.615
R1754 VTAIL.n182 VTAIL.n101 104.615
R1755 VTAIL.n189 VTAIL.n101 104.615
R1756 VTAIL.n190 VTAIL.n189 104.615
R1757 VTAIL.n230 VTAIL.n229 104.615
R1758 VTAIL.n230 VTAIL.n223 104.615
R1759 VTAIL.n237 VTAIL.n223 104.615
R1760 VTAIL.n238 VTAIL.n237 104.615
R1761 VTAIL.n238 VTAIL.n219 104.615
R1762 VTAIL.n245 VTAIL.n219 104.615
R1763 VTAIL.n246 VTAIL.n245 104.615
R1764 VTAIL.n246 VTAIL.n215 104.615
R1765 VTAIL.n253 VTAIL.n215 104.615
R1766 VTAIL.n254 VTAIL.n253 104.615
R1767 VTAIL.n254 VTAIL.n211 104.615
R1768 VTAIL.n261 VTAIL.n211 104.615
R1769 VTAIL.n262 VTAIL.n261 104.615
R1770 VTAIL.n262 VTAIL.n207 104.615
R1771 VTAIL.n270 VTAIL.n207 104.615
R1772 VTAIL.n271 VTAIL.n270 104.615
R1773 VTAIL.n272 VTAIL.n271 104.615
R1774 VTAIL.n272 VTAIL.n203 104.615
R1775 VTAIL.n279 VTAIL.n203 104.615
R1776 VTAIL.n280 VTAIL.n279 104.615
R1777 VTAIL.n280 VTAIL.n199 104.615
R1778 VTAIL.n287 VTAIL.n199 104.615
R1779 VTAIL.n288 VTAIL.n287 104.615
R1780 VTAIL.n680 VTAIL.n679 104.615
R1781 VTAIL.n679 VTAIL.n591 104.615
R1782 VTAIL.n672 VTAIL.n591 104.615
R1783 VTAIL.n672 VTAIL.n671 104.615
R1784 VTAIL.n671 VTAIL.n595 104.615
R1785 VTAIL.n600 VTAIL.n595 104.615
R1786 VTAIL.n664 VTAIL.n600 104.615
R1787 VTAIL.n664 VTAIL.n663 104.615
R1788 VTAIL.n663 VTAIL.n601 104.615
R1789 VTAIL.n656 VTAIL.n601 104.615
R1790 VTAIL.n656 VTAIL.n655 104.615
R1791 VTAIL.n655 VTAIL.n605 104.615
R1792 VTAIL.n648 VTAIL.n605 104.615
R1793 VTAIL.n648 VTAIL.n647 104.615
R1794 VTAIL.n647 VTAIL.n609 104.615
R1795 VTAIL.n640 VTAIL.n609 104.615
R1796 VTAIL.n640 VTAIL.n639 104.615
R1797 VTAIL.n639 VTAIL.n613 104.615
R1798 VTAIL.n632 VTAIL.n613 104.615
R1799 VTAIL.n632 VTAIL.n631 104.615
R1800 VTAIL.n631 VTAIL.n617 104.615
R1801 VTAIL.n624 VTAIL.n617 104.615
R1802 VTAIL.n624 VTAIL.n623 104.615
R1803 VTAIL.n582 VTAIL.n581 104.615
R1804 VTAIL.n581 VTAIL.n493 104.615
R1805 VTAIL.n574 VTAIL.n493 104.615
R1806 VTAIL.n574 VTAIL.n573 104.615
R1807 VTAIL.n573 VTAIL.n497 104.615
R1808 VTAIL.n502 VTAIL.n497 104.615
R1809 VTAIL.n566 VTAIL.n502 104.615
R1810 VTAIL.n566 VTAIL.n565 104.615
R1811 VTAIL.n565 VTAIL.n503 104.615
R1812 VTAIL.n558 VTAIL.n503 104.615
R1813 VTAIL.n558 VTAIL.n557 104.615
R1814 VTAIL.n557 VTAIL.n507 104.615
R1815 VTAIL.n550 VTAIL.n507 104.615
R1816 VTAIL.n550 VTAIL.n549 104.615
R1817 VTAIL.n549 VTAIL.n511 104.615
R1818 VTAIL.n542 VTAIL.n511 104.615
R1819 VTAIL.n542 VTAIL.n541 104.615
R1820 VTAIL.n541 VTAIL.n515 104.615
R1821 VTAIL.n534 VTAIL.n515 104.615
R1822 VTAIL.n534 VTAIL.n533 104.615
R1823 VTAIL.n533 VTAIL.n519 104.615
R1824 VTAIL.n526 VTAIL.n519 104.615
R1825 VTAIL.n526 VTAIL.n525 104.615
R1826 VTAIL.n484 VTAIL.n483 104.615
R1827 VTAIL.n483 VTAIL.n395 104.615
R1828 VTAIL.n476 VTAIL.n395 104.615
R1829 VTAIL.n476 VTAIL.n475 104.615
R1830 VTAIL.n475 VTAIL.n399 104.615
R1831 VTAIL.n404 VTAIL.n399 104.615
R1832 VTAIL.n468 VTAIL.n404 104.615
R1833 VTAIL.n468 VTAIL.n467 104.615
R1834 VTAIL.n467 VTAIL.n405 104.615
R1835 VTAIL.n460 VTAIL.n405 104.615
R1836 VTAIL.n460 VTAIL.n459 104.615
R1837 VTAIL.n459 VTAIL.n409 104.615
R1838 VTAIL.n452 VTAIL.n409 104.615
R1839 VTAIL.n452 VTAIL.n451 104.615
R1840 VTAIL.n451 VTAIL.n413 104.615
R1841 VTAIL.n444 VTAIL.n413 104.615
R1842 VTAIL.n444 VTAIL.n443 104.615
R1843 VTAIL.n443 VTAIL.n417 104.615
R1844 VTAIL.n436 VTAIL.n417 104.615
R1845 VTAIL.n436 VTAIL.n435 104.615
R1846 VTAIL.n435 VTAIL.n421 104.615
R1847 VTAIL.n428 VTAIL.n421 104.615
R1848 VTAIL.n428 VTAIL.n427 104.615
R1849 VTAIL.n386 VTAIL.n385 104.615
R1850 VTAIL.n385 VTAIL.n297 104.615
R1851 VTAIL.n378 VTAIL.n297 104.615
R1852 VTAIL.n378 VTAIL.n377 104.615
R1853 VTAIL.n377 VTAIL.n301 104.615
R1854 VTAIL.n306 VTAIL.n301 104.615
R1855 VTAIL.n370 VTAIL.n306 104.615
R1856 VTAIL.n370 VTAIL.n369 104.615
R1857 VTAIL.n369 VTAIL.n307 104.615
R1858 VTAIL.n362 VTAIL.n307 104.615
R1859 VTAIL.n362 VTAIL.n361 104.615
R1860 VTAIL.n361 VTAIL.n311 104.615
R1861 VTAIL.n354 VTAIL.n311 104.615
R1862 VTAIL.n354 VTAIL.n353 104.615
R1863 VTAIL.n353 VTAIL.n315 104.615
R1864 VTAIL.n346 VTAIL.n315 104.615
R1865 VTAIL.n346 VTAIL.n345 104.615
R1866 VTAIL.n345 VTAIL.n319 104.615
R1867 VTAIL.n338 VTAIL.n319 104.615
R1868 VTAIL.n338 VTAIL.n337 104.615
R1869 VTAIL.n337 VTAIL.n323 104.615
R1870 VTAIL.n330 VTAIL.n323 104.615
R1871 VTAIL.n330 VTAIL.n329 104.615
R1872 VTAIL.n719 VTAIL.t2 52.3082
R1873 VTAIL.n33 VTAIL.t1 52.3082
R1874 VTAIL.n131 VTAIL.t4 52.3082
R1875 VTAIL.n229 VTAIL.t7 52.3082
R1876 VTAIL.n623 VTAIL.t6 52.3082
R1877 VTAIL.n525 VTAIL.t5 52.3082
R1878 VTAIL.n427 VTAIL.t0 52.3082
R1879 VTAIL.n329 VTAIL.t3 52.3082
R1880 VTAIL.n783 VTAIL.n782 31.6035
R1881 VTAIL.n97 VTAIL.n96 31.6035
R1882 VTAIL.n195 VTAIL.n194 31.6035
R1883 VTAIL.n293 VTAIL.n292 31.6035
R1884 VTAIL.n685 VTAIL.n684 31.6035
R1885 VTAIL.n587 VTAIL.n586 31.6035
R1886 VTAIL.n489 VTAIL.n488 31.6035
R1887 VTAIL.n391 VTAIL.n390 31.6035
R1888 VTAIL.n783 VTAIL.n685 28.9014
R1889 VTAIL.n391 VTAIL.n293 28.9014
R1890 VTAIL.n718 VTAIL.n717 15.6677
R1891 VTAIL.n32 VTAIL.n31 15.6677
R1892 VTAIL.n130 VTAIL.n129 15.6677
R1893 VTAIL.n228 VTAIL.n227 15.6677
R1894 VTAIL.n622 VTAIL.n621 15.6677
R1895 VTAIL.n524 VTAIL.n523 15.6677
R1896 VTAIL.n426 VTAIL.n425 15.6677
R1897 VTAIL.n328 VTAIL.n327 15.6677
R1898 VTAIL.n763 VTAIL.n694 13.1884
R1899 VTAIL.n77 VTAIL.n8 13.1884
R1900 VTAIL.n175 VTAIL.n106 13.1884
R1901 VTAIL.n273 VTAIL.n204 13.1884
R1902 VTAIL.n598 VTAIL.n596 13.1884
R1903 VTAIL.n500 VTAIL.n498 13.1884
R1904 VTAIL.n402 VTAIL.n400 13.1884
R1905 VTAIL.n304 VTAIL.n302 13.1884
R1906 VTAIL.n721 VTAIL.n716 12.8005
R1907 VTAIL.n764 VTAIL.n696 12.8005
R1908 VTAIL.n768 VTAIL.n767 12.8005
R1909 VTAIL.n35 VTAIL.n30 12.8005
R1910 VTAIL.n78 VTAIL.n10 12.8005
R1911 VTAIL.n82 VTAIL.n81 12.8005
R1912 VTAIL.n133 VTAIL.n128 12.8005
R1913 VTAIL.n176 VTAIL.n108 12.8005
R1914 VTAIL.n180 VTAIL.n179 12.8005
R1915 VTAIL.n231 VTAIL.n226 12.8005
R1916 VTAIL.n274 VTAIL.n206 12.8005
R1917 VTAIL.n278 VTAIL.n277 12.8005
R1918 VTAIL.n670 VTAIL.n669 12.8005
R1919 VTAIL.n666 VTAIL.n665 12.8005
R1920 VTAIL.n625 VTAIL.n620 12.8005
R1921 VTAIL.n572 VTAIL.n571 12.8005
R1922 VTAIL.n568 VTAIL.n567 12.8005
R1923 VTAIL.n527 VTAIL.n522 12.8005
R1924 VTAIL.n474 VTAIL.n473 12.8005
R1925 VTAIL.n470 VTAIL.n469 12.8005
R1926 VTAIL.n429 VTAIL.n424 12.8005
R1927 VTAIL.n376 VTAIL.n375 12.8005
R1928 VTAIL.n372 VTAIL.n371 12.8005
R1929 VTAIL.n331 VTAIL.n326 12.8005
R1930 VTAIL.n722 VTAIL.n714 12.0247
R1931 VTAIL.n759 VTAIL.n758 12.0247
R1932 VTAIL.n771 VTAIL.n692 12.0247
R1933 VTAIL.n36 VTAIL.n28 12.0247
R1934 VTAIL.n73 VTAIL.n72 12.0247
R1935 VTAIL.n85 VTAIL.n6 12.0247
R1936 VTAIL.n134 VTAIL.n126 12.0247
R1937 VTAIL.n171 VTAIL.n170 12.0247
R1938 VTAIL.n183 VTAIL.n104 12.0247
R1939 VTAIL.n232 VTAIL.n224 12.0247
R1940 VTAIL.n269 VTAIL.n268 12.0247
R1941 VTAIL.n281 VTAIL.n202 12.0247
R1942 VTAIL.n673 VTAIL.n594 12.0247
R1943 VTAIL.n662 VTAIL.n599 12.0247
R1944 VTAIL.n626 VTAIL.n618 12.0247
R1945 VTAIL.n575 VTAIL.n496 12.0247
R1946 VTAIL.n564 VTAIL.n501 12.0247
R1947 VTAIL.n528 VTAIL.n520 12.0247
R1948 VTAIL.n477 VTAIL.n398 12.0247
R1949 VTAIL.n466 VTAIL.n403 12.0247
R1950 VTAIL.n430 VTAIL.n422 12.0247
R1951 VTAIL.n379 VTAIL.n300 12.0247
R1952 VTAIL.n368 VTAIL.n305 12.0247
R1953 VTAIL.n332 VTAIL.n324 12.0247
R1954 VTAIL.n726 VTAIL.n725 11.249
R1955 VTAIL.n757 VTAIL.n698 11.249
R1956 VTAIL.n772 VTAIL.n690 11.249
R1957 VTAIL.n40 VTAIL.n39 11.249
R1958 VTAIL.n71 VTAIL.n12 11.249
R1959 VTAIL.n86 VTAIL.n4 11.249
R1960 VTAIL.n138 VTAIL.n137 11.249
R1961 VTAIL.n169 VTAIL.n110 11.249
R1962 VTAIL.n184 VTAIL.n102 11.249
R1963 VTAIL.n236 VTAIL.n235 11.249
R1964 VTAIL.n267 VTAIL.n208 11.249
R1965 VTAIL.n282 VTAIL.n200 11.249
R1966 VTAIL.n674 VTAIL.n592 11.249
R1967 VTAIL.n661 VTAIL.n602 11.249
R1968 VTAIL.n630 VTAIL.n629 11.249
R1969 VTAIL.n576 VTAIL.n494 11.249
R1970 VTAIL.n563 VTAIL.n504 11.249
R1971 VTAIL.n532 VTAIL.n531 11.249
R1972 VTAIL.n478 VTAIL.n396 11.249
R1973 VTAIL.n465 VTAIL.n406 11.249
R1974 VTAIL.n434 VTAIL.n433 11.249
R1975 VTAIL.n380 VTAIL.n298 11.249
R1976 VTAIL.n367 VTAIL.n308 11.249
R1977 VTAIL.n336 VTAIL.n335 11.249
R1978 VTAIL.n729 VTAIL.n712 10.4732
R1979 VTAIL.n754 VTAIL.n753 10.4732
R1980 VTAIL.n776 VTAIL.n775 10.4732
R1981 VTAIL.n43 VTAIL.n26 10.4732
R1982 VTAIL.n68 VTAIL.n67 10.4732
R1983 VTAIL.n90 VTAIL.n89 10.4732
R1984 VTAIL.n141 VTAIL.n124 10.4732
R1985 VTAIL.n166 VTAIL.n165 10.4732
R1986 VTAIL.n188 VTAIL.n187 10.4732
R1987 VTAIL.n239 VTAIL.n222 10.4732
R1988 VTAIL.n264 VTAIL.n263 10.4732
R1989 VTAIL.n286 VTAIL.n285 10.4732
R1990 VTAIL.n678 VTAIL.n677 10.4732
R1991 VTAIL.n658 VTAIL.n657 10.4732
R1992 VTAIL.n633 VTAIL.n616 10.4732
R1993 VTAIL.n580 VTAIL.n579 10.4732
R1994 VTAIL.n560 VTAIL.n559 10.4732
R1995 VTAIL.n535 VTAIL.n518 10.4732
R1996 VTAIL.n482 VTAIL.n481 10.4732
R1997 VTAIL.n462 VTAIL.n461 10.4732
R1998 VTAIL.n437 VTAIL.n420 10.4732
R1999 VTAIL.n384 VTAIL.n383 10.4732
R2000 VTAIL.n364 VTAIL.n363 10.4732
R2001 VTAIL.n339 VTAIL.n322 10.4732
R2002 VTAIL.n730 VTAIL.n710 9.69747
R2003 VTAIL.n750 VTAIL.n700 9.69747
R2004 VTAIL.n779 VTAIL.n688 9.69747
R2005 VTAIL.n44 VTAIL.n24 9.69747
R2006 VTAIL.n64 VTAIL.n14 9.69747
R2007 VTAIL.n93 VTAIL.n2 9.69747
R2008 VTAIL.n142 VTAIL.n122 9.69747
R2009 VTAIL.n162 VTAIL.n112 9.69747
R2010 VTAIL.n191 VTAIL.n100 9.69747
R2011 VTAIL.n240 VTAIL.n220 9.69747
R2012 VTAIL.n260 VTAIL.n210 9.69747
R2013 VTAIL.n289 VTAIL.n198 9.69747
R2014 VTAIL.n681 VTAIL.n590 9.69747
R2015 VTAIL.n654 VTAIL.n604 9.69747
R2016 VTAIL.n634 VTAIL.n614 9.69747
R2017 VTAIL.n583 VTAIL.n492 9.69747
R2018 VTAIL.n556 VTAIL.n506 9.69747
R2019 VTAIL.n536 VTAIL.n516 9.69747
R2020 VTAIL.n485 VTAIL.n394 9.69747
R2021 VTAIL.n458 VTAIL.n408 9.69747
R2022 VTAIL.n438 VTAIL.n418 9.69747
R2023 VTAIL.n387 VTAIL.n296 9.69747
R2024 VTAIL.n360 VTAIL.n310 9.69747
R2025 VTAIL.n340 VTAIL.n320 9.69747
R2026 VTAIL.n782 VTAIL.n781 9.45567
R2027 VTAIL.n96 VTAIL.n95 9.45567
R2028 VTAIL.n194 VTAIL.n193 9.45567
R2029 VTAIL.n292 VTAIL.n291 9.45567
R2030 VTAIL.n684 VTAIL.n683 9.45567
R2031 VTAIL.n586 VTAIL.n585 9.45567
R2032 VTAIL.n488 VTAIL.n487 9.45567
R2033 VTAIL.n390 VTAIL.n389 9.45567
R2034 VTAIL.n781 VTAIL.n780 9.3005
R2035 VTAIL.n688 VTAIL.n687 9.3005
R2036 VTAIL.n775 VTAIL.n774 9.3005
R2037 VTAIL.n773 VTAIL.n772 9.3005
R2038 VTAIL.n692 VTAIL.n691 9.3005
R2039 VTAIL.n767 VTAIL.n766 9.3005
R2040 VTAIL.n739 VTAIL.n738 9.3005
R2041 VTAIL.n708 VTAIL.n707 9.3005
R2042 VTAIL.n733 VTAIL.n732 9.3005
R2043 VTAIL.n731 VTAIL.n730 9.3005
R2044 VTAIL.n712 VTAIL.n711 9.3005
R2045 VTAIL.n725 VTAIL.n724 9.3005
R2046 VTAIL.n723 VTAIL.n722 9.3005
R2047 VTAIL.n716 VTAIL.n715 9.3005
R2048 VTAIL.n741 VTAIL.n740 9.3005
R2049 VTAIL.n704 VTAIL.n703 9.3005
R2050 VTAIL.n747 VTAIL.n746 9.3005
R2051 VTAIL.n749 VTAIL.n748 9.3005
R2052 VTAIL.n700 VTAIL.n699 9.3005
R2053 VTAIL.n755 VTAIL.n754 9.3005
R2054 VTAIL.n757 VTAIL.n756 9.3005
R2055 VTAIL.n758 VTAIL.n695 9.3005
R2056 VTAIL.n765 VTAIL.n764 9.3005
R2057 VTAIL.n95 VTAIL.n94 9.3005
R2058 VTAIL.n2 VTAIL.n1 9.3005
R2059 VTAIL.n89 VTAIL.n88 9.3005
R2060 VTAIL.n87 VTAIL.n86 9.3005
R2061 VTAIL.n6 VTAIL.n5 9.3005
R2062 VTAIL.n81 VTAIL.n80 9.3005
R2063 VTAIL.n53 VTAIL.n52 9.3005
R2064 VTAIL.n22 VTAIL.n21 9.3005
R2065 VTAIL.n47 VTAIL.n46 9.3005
R2066 VTAIL.n45 VTAIL.n44 9.3005
R2067 VTAIL.n26 VTAIL.n25 9.3005
R2068 VTAIL.n39 VTAIL.n38 9.3005
R2069 VTAIL.n37 VTAIL.n36 9.3005
R2070 VTAIL.n30 VTAIL.n29 9.3005
R2071 VTAIL.n55 VTAIL.n54 9.3005
R2072 VTAIL.n18 VTAIL.n17 9.3005
R2073 VTAIL.n61 VTAIL.n60 9.3005
R2074 VTAIL.n63 VTAIL.n62 9.3005
R2075 VTAIL.n14 VTAIL.n13 9.3005
R2076 VTAIL.n69 VTAIL.n68 9.3005
R2077 VTAIL.n71 VTAIL.n70 9.3005
R2078 VTAIL.n72 VTAIL.n9 9.3005
R2079 VTAIL.n79 VTAIL.n78 9.3005
R2080 VTAIL.n193 VTAIL.n192 9.3005
R2081 VTAIL.n100 VTAIL.n99 9.3005
R2082 VTAIL.n187 VTAIL.n186 9.3005
R2083 VTAIL.n185 VTAIL.n184 9.3005
R2084 VTAIL.n104 VTAIL.n103 9.3005
R2085 VTAIL.n179 VTAIL.n178 9.3005
R2086 VTAIL.n151 VTAIL.n150 9.3005
R2087 VTAIL.n120 VTAIL.n119 9.3005
R2088 VTAIL.n145 VTAIL.n144 9.3005
R2089 VTAIL.n143 VTAIL.n142 9.3005
R2090 VTAIL.n124 VTAIL.n123 9.3005
R2091 VTAIL.n137 VTAIL.n136 9.3005
R2092 VTAIL.n135 VTAIL.n134 9.3005
R2093 VTAIL.n128 VTAIL.n127 9.3005
R2094 VTAIL.n153 VTAIL.n152 9.3005
R2095 VTAIL.n116 VTAIL.n115 9.3005
R2096 VTAIL.n159 VTAIL.n158 9.3005
R2097 VTAIL.n161 VTAIL.n160 9.3005
R2098 VTAIL.n112 VTAIL.n111 9.3005
R2099 VTAIL.n167 VTAIL.n166 9.3005
R2100 VTAIL.n169 VTAIL.n168 9.3005
R2101 VTAIL.n170 VTAIL.n107 9.3005
R2102 VTAIL.n177 VTAIL.n176 9.3005
R2103 VTAIL.n291 VTAIL.n290 9.3005
R2104 VTAIL.n198 VTAIL.n197 9.3005
R2105 VTAIL.n285 VTAIL.n284 9.3005
R2106 VTAIL.n283 VTAIL.n282 9.3005
R2107 VTAIL.n202 VTAIL.n201 9.3005
R2108 VTAIL.n277 VTAIL.n276 9.3005
R2109 VTAIL.n249 VTAIL.n248 9.3005
R2110 VTAIL.n218 VTAIL.n217 9.3005
R2111 VTAIL.n243 VTAIL.n242 9.3005
R2112 VTAIL.n241 VTAIL.n240 9.3005
R2113 VTAIL.n222 VTAIL.n221 9.3005
R2114 VTAIL.n235 VTAIL.n234 9.3005
R2115 VTAIL.n233 VTAIL.n232 9.3005
R2116 VTAIL.n226 VTAIL.n225 9.3005
R2117 VTAIL.n251 VTAIL.n250 9.3005
R2118 VTAIL.n214 VTAIL.n213 9.3005
R2119 VTAIL.n257 VTAIL.n256 9.3005
R2120 VTAIL.n259 VTAIL.n258 9.3005
R2121 VTAIL.n210 VTAIL.n209 9.3005
R2122 VTAIL.n265 VTAIL.n264 9.3005
R2123 VTAIL.n267 VTAIL.n266 9.3005
R2124 VTAIL.n268 VTAIL.n205 9.3005
R2125 VTAIL.n275 VTAIL.n274 9.3005
R2126 VTAIL.n608 VTAIL.n607 9.3005
R2127 VTAIL.n651 VTAIL.n650 9.3005
R2128 VTAIL.n653 VTAIL.n652 9.3005
R2129 VTAIL.n604 VTAIL.n603 9.3005
R2130 VTAIL.n659 VTAIL.n658 9.3005
R2131 VTAIL.n661 VTAIL.n660 9.3005
R2132 VTAIL.n599 VTAIL.n597 9.3005
R2133 VTAIL.n667 VTAIL.n666 9.3005
R2134 VTAIL.n683 VTAIL.n682 9.3005
R2135 VTAIL.n590 VTAIL.n589 9.3005
R2136 VTAIL.n677 VTAIL.n676 9.3005
R2137 VTAIL.n675 VTAIL.n674 9.3005
R2138 VTAIL.n594 VTAIL.n593 9.3005
R2139 VTAIL.n669 VTAIL.n668 9.3005
R2140 VTAIL.n645 VTAIL.n644 9.3005
R2141 VTAIL.n643 VTAIL.n642 9.3005
R2142 VTAIL.n612 VTAIL.n611 9.3005
R2143 VTAIL.n637 VTAIL.n636 9.3005
R2144 VTAIL.n635 VTAIL.n634 9.3005
R2145 VTAIL.n616 VTAIL.n615 9.3005
R2146 VTAIL.n629 VTAIL.n628 9.3005
R2147 VTAIL.n627 VTAIL.n626 9.3005
R2148 VTAIL.n620 VTAIL.n619 9.3005
R2149 VTAIL.n510 VTAIL.n509 9.3005
R2150 VTAIL.n553 VTAIL.n552 9.3005
R2151 VTAIL.n555 VTAIL.n554 9.3005
R2152 VTAIL.n506 VTAIL.n505 9.3005
R2153 VTAIL.n561 VTAIL.n560 9.3005
R2154 VTAIL.n563 VTAIL.n562 9.3005
R2155 VTAIL.n501 VTAIL.n499 9.3005
R2156 VTAIL.n569 VTAIL.n568 9.3005
R2157 VTAIL.n585 VTAIL.n584 9.3005
R2158 VTAIL.n492 VTAIL.n491 9.3005
R2159 VTAIL.n579 VTAIL.n578 9.3005
R2160 VTAIL.n577 VTAIL.n576 9.3005
R2161 VTAIL.n496 VTAIL.n495 9.3005
R2162 VTAIL.n571 VTAIL.n570 9.3005
R2163 VTAIL.n547 VTAIL.n546 9.3005
R2164 VTAIL.n545 VTAIL.n544 9.3005
R2165 VTAIL.n514 VTAIL.n513 9.3005
R2166 VTAIL.n539 VTAIL.n538 9.3005
R2167 VTAIL.n537 VTAIL.n536 9.3005
R2168 VTAIL.n518 VTAIL.n517 9.3005
R2169 VTAIL.n531 VTAIL.n530 9.3005
R2170 VTAIL.n529 VTAIL.n528 9.3005
R2171 VTAIL.n522 VTAIL.n521 9.3005
R2172 VTAIL.n412 VTAIL.n411 9.3005
R2173 VTAIL.n455 VTAIL.n454 9.3005
R2174 VTAIL.n457 VTAIL.n456 9.3005
R2175 VTAIL.n408 VTAIL.n407 9.3005
R2176 VTAIL.n463 VTAIL.n462 9.3005
R2177 VTAIL.n465 VTAIL.n464 9.3005
R2178 VTAIL.n403 VTAIL.n401 9.3005
R2179 VTAIL.n471 VTAIL.n470 9.3005
R2180 VTAIL.n487 VTAIL.n486 9.3005
R2181 VTAIL.n394 VTAIL.n393 9.3005
R2182 VTAIL.n481 VTAIL.n480 9.3005
R2183 VTAIL.n479 VTAIL.n478 9.3005
R2184 VTAIL.n398 VTAIL.n397 9.3005
R2185 VTAIL.n473 VTAIL.n472 9.3005
R2186 VTAIL.n449 VTAIL.n448 9.3005
R2187 VTAIL.n447 VTAIL.n446 9.3005
R2188 VTAIL.n416 VTAIL.n415 9.3005
R2189 VTAIL.n441 VTAIL.n440 9.3005
R2190 VTAIL.n439 VTAIL.n438 9.3005
R2191 VTAIL.n420 VTAIL.n419 9.3005
R2192 VTAIL.n433 VTAIL.n432 9.3005
R2193 VTAIL.n431 VTAIL.n430 9.3005
R2194 VTAIL.n424 VTAIL.n423 9.3005
R2195 VTAIL.n314 VTAIL.n313 9.3005
R2196 VTAIL.n357 VTAIL.n356 9.3005
R2197 VTAIL.n359 VTAIL.n358 9.3005
R2198 VTAIL.n310 VTAIL.n309 9.3005
R2199 VTAIL.n365 VTAIL.n364 9.3005
R2200 VTAIL.n367 VTAIL.n366 9.3005
R2201 VTAIL.n305 VTAIL.n303 9.3005
R2202 VTAIL.n373 VTAIL.n372 9.3005
R2203 VTAIL.n389 VTAIL.n388 9.3005
R2204 VTAIL.n296 VTAIL.n295 9.3005
R2205 VTAIL.n383 VTAIL.n382 9.3005
R2206 VTAIL.n381 VTAIL.n380 9.3005
R2207 VTAIL.n300 VTAIL.n299 9.3005
R2208 VTAIL.n375 VTAIL.n374 9.3005
R2209 VTAIL.n351 VTAIL.n350 9.3005
R2210 VTAIL.n349 VTAIL.n348 9.3005
R2211 VTAIL.n318 VTAIL.n317 9.3005
R2212 VTAIL.n343 VTAIL.n342 9.3005
R2213 VTAIL.n341 VTAIL.n340 9.3005
R2214 VTAIL.n322 VTAIL.n321 9.3005
R2215 VTAIL.n335 VTAIL.n334 9.3005
R2216 VTAIL.n333 VTAIL.n332 9.3005
R2217 VTAIL.n326 VTAIL.n325 9.3005
R2218 VTAIL.n734 VTAIL.n733 8.92171
R2219 VTAIL.n749 VTAIL.n702 8.92171
R2220 VTAIL.n780 VTAIL.n686 8.92171
R2221 VTAIL.n48 VTAIL.n47 8.92171
R2222 VTAIL.n63 VTAIL.n16 8.92171
R2223 VTAIL.n94 VTAIL.n0 8.92171
R2224 VTAIL.n146 VTAIL.n145 8.92171
R2225 VTAIL.n161 VTAIL.n114 8.92171
R2226 VTAIL.n192 VTAIL.n98 8.92171
R2227 VTAIL.n244 VTAIL.n243 8.92171
R2228 VTAIL.n259 VTAIL.n212 8.92171
R2229 VTAIL.n290 VTAIL.n196 8.92171
R2230 VTAIL.n682 VTAIL.n588 8.92171
R2231 VTAIL.n653 VTAIL.n606 8.92171
R2232 VTAIL.n638 VTAIL.n637 8.92171
R2233 VTAIL.n584 VTAIL.n490 8.92171
R2234 VTAIL.n555 VTAIL.n508 8.92171
R2235 VTAIL.n540 VTAIL.n539 8.92171
R2236 VTAIL.n486 VTAIL.n392 8.92171
R2237 VTAIL.n457 VTAIL.n410 8.92171
R2238 VTAIL.n442 VTAIL.n441 8.92171
R2239 VTAIL.n388 VTAIL.n294 8.92171
R2240 VTAIL.n359 VTAIL.n312 8.92171
R2241 VTAIL.n344 VTAIL.n343 8.92171
R2242 VTAIL.n737 VTAIL.n708 8.14595
R2243 VTAIL.n746 VTAIL.n745 8.14595
R2244 VTAIL.n51 VTAIL.n22 8.14595
R2245 VTAIL.n60 VTAIL.n59 8.14595
R2246 VTAIL.n149 VTAIL.n120 8.14595
R2247 VTAIL.n158 VTAIL.n157 8.14595
R2248 VTAIL.n247 VTAIL.n218 8.14595
R2249 VTAIL.n256 VTAIL.n255 8.14595
R2250 VTAIL.n650 VTAIL.n649 8.14595
R2251 VTAIL.n641 VTAIL.n612 8.14595
R2252 VTAIL.n552 VTAIL.n551 8.14595
R2253 VTAIL.n543 VTAIL.n514 8.14595
R2254 VTAIL.n454 VTAIL.n453 8.14595
R2255 VTAIL.n445 VTAIL.n416 8.14595
R2256 VTAIL.n356 VTAIL.n355 8.14595
R2257 VTAIL.n347 VTAIL.n318 8.14595
R2258 VTAIL.n738 VTAIL.n706 7.3702
R2259 VTAIL.n742 VTAIL.n704 7.3702
R2260 VTAIL.n52 VTAIL.n20 7.3702
R2261 VTAIL.n56 VTAIL.n18 7.3702
R2262 VTAIL.n150 VTAIL.n118 7.3702
R2263 VTAIL.n154 VTAIL.n116 7.3702
R2264 VTAIL.n248 VTAIL.n216 7.3702
R2265 VTAIL.n252 VTAIL.n214 7.3702
R2266 VTAIL.n646 VTAIL.n608 7.3702
R2267 VTAIL.n642 VTAIL.n610 7.3702
R2268 VTAIL.n548 VTAIL.n510 7.3702
R2269 VTAIL.n544 VTAIL.n512 7.3702
R2270 VTAIL.n450 VTAIL.n412 7.3702
R2271 VTAIL.n446 VTAIL.n414 7.3702
R2272 VTAIL.n352 VTAIL.n314 7.3702
R2273 VTAIL.n348 VTAIL.n316 7.3702
R2274 VTAIL.n741 VTAIL.n706 6.59444
R2275 VTAIL.n742 VTAIL.n741 6.59444
R2276 VTAIL.n55 VTAIL.n20 6.59444
R2277 VTAIL.n56 VTAIL.n55 6.59444
R2278 VTAIL.n153 VTAIL.n118 6.59444
R2279 VTAIL.n154 VTAIL.n153 6.59444
R2280 VTAIL.n251 VTAIL.n216 6.59444
R2281 VTAIL.n252 VTAIL.n251 6.59444
R2282 VTAIL.n646 VTAIL.n645 6.59444
R2283 VTAIL.n645 VTAIL.n610 6.59444
R2284 VTAIL.n548 VTAIL.n547 6.59444
R2285 VTAIL.n547 VTAIL.n512 6.59444
R2286 VTAIL.n450 VTAIL.n449 6.59444
R2287 VTAIL.n449 VTAIL.n414 6.59444
R2288 VTAIL.n352 VTAIL.n351 6.59444
R2289 VTAIL.n351 VTAIL.n316 6.59444
R2290 VTAIL.n738 VTAIL.n737 5.81868
R2291 VTAIL.n745 VTAIL.n704 5.81868
R2292 VTAIL.n52 VTAIL.n51 5.81868
R2293 VTAIL.n59 VTAIL.n18 5.81868
R2294 VTAIL.n150 VTAIL.n149 5.81868
R2295 VTAIL.n157 VTAIL.n116 5.81868
R2296 VTAIL.n248 VTAIL.n247 5.81868
R2297 VTAIL.n255 VTAIL.n214 5.81868
R2298 VTAIL.n649 VTAIL.n608 5.81868
R2299 VTAIL.n642 VTAIL.n641 5.81868
R2300 VTAIL.n551 VTAIL.n510 5.81868
R2301 VTAIL.n544 VTAIL.n543 5.81868
R2302 VTAIL.n453 VTAIL.n412 5.81868
R2303 VTAIL.n446 VTAIL.n445 5.81868
R2304 VTAIL.n355 VTAIL.n314 5.81868
R2305 VTAIL.n348 VTAIL.n347 5.81868
R2306 VTAIL.n734 VTAIL.n708 5.04292
R2307 VTAIL.n746 VTAIL.n702 5.04292
R2308 VTAIL.n782 VTAIL.n686 5.04292
R2309 VTAIL.n48 VTAIL.n22 5.04292
R2310 VTAIL.n60 VTAIL.n16 5.04292
R2311 VTAIL.n96 VTAIL.n0 5.04292
R2312 VTAIL.n146 VTAIL.n120 5.04292
R2313 VTAIL.n158 VTAIL.n114 5.04292
R2314 VTAIL.n194 VTAIL.n98 5.04292
R2315 VTAIL.n244 VTAIL.n218 5.04292
R2316 VTAIL.n256 VTAIL.n212 5.04292
R2317 VTAIL.n292 VTAIL.n196 5.04292
R2318 VTAIL.n684 VTAIL.n588 5.04292
R2319 VTAIL.n650 VTAIL.n606 5.04292
R2320 VTAIL.n638 VTAIL.n612 5.04292
R2321 VTAIL.n586 VTAIL.n490 5.04292
R2322 VTAIL.n552 VTAIL.n508 5.04292
R2323 VTAIL.n540 VTAIL.n514 5.04292
R2324 VTAIL.n488 VTAIL.n392 5.04292
R2325 VTAIL.n454 VTAIL.n410 5.04292
R2326 VTAIL.n442 VTAIL.n416 5.04292
R2327 VTAIL.n390 VTAIL.n294 5.04292
R2328 VTAIL.n356 VTAIL.n312 5.04292
R2329 VTAIL.n344 VTAIL.n318 5.04292
R2330 VTAIL.n717 VTAIL.n715 4.38563
R2331 VTAIL.n31 VTAIL.n29 4.38563
R2332 VTAIL.n129 VTAIL.n127 4.38563
R2333 VTAIL.n227 VTAIL.n225 4.38563
R2334 VTAIL.n621 VTAIL.n619 4.38563
R2335 VTAIL.n523 VTAIL.n521 4.38563
R2336 VTAIL.n425 VTAIL.n423 4.38563
R2337 VTAIL.n327 VTAIL.n325 4.38563
R2338 VTAIL.n733 VTAIL.n710 4.26717
R2339 VTAIL.n750 VTAIL.n749 4.26717
R2340 VTAIL.n780 VTAIL.n779 4.26717
R2341 VTAIL.n47 VTAIL.n24 4.26717
R2342 VTAIL.n64 VTAIL.n63 4.26717
R2343 VTAIL.n94 VTAIL.n93 4.26717
R2344 VTAIL.n145 VTAIL.n122 4.26717
R2345 VTAIL.n162 VTAIL.n161 4.26717
R2346 VTAIL.n192 VTAIL.n191 4.26717
R2347 VTAIL.n243 VTAIL.n220 4.26717
R2348 VTAIL.n260 VTAIL.n259 4.26717
R2349 VTAIL.n290 VTAIL.n289 4.26717
R2350 VTAIL.n682 VTAIL.n681 4.26717
R2351 VTAIL.n654 VTAIL.n653 4.26717
R2352 VTAIL.n637 VTAIL.n614 4.26717
R2353 VTAIL.n584 VTAIL.n583 4.26717
R2354 VTAIL.n556 VTAIL.n555 4.26717
R2355 VTAIL.n539 VTAIL.n516 4.26717
R2356 VTAIL.n486 VTAIL.n485 4.26717
R2357 VTAIL.n458 VTAIL.n457 4.26717
R2358 VTAIL.n441 VTAIL.n418 4.26717
R2359 VTAIL.n388 VTAIL.n387 4.26717
R2360 VTAIL.n360 VTAIL.n359 4.26717
R2361 VTAIL.n343 VTAIL.n320 4.26717
R2362 VTAIL.n730 VTAIL.n729 3.49141
R2363 VTAIL.n753 VTAIL.n700 3.49141
R2364 VTAIL.n776 VTAIL.n688 3.49141
R2365 VTAIL.n44 VTAIL.n43 3.49141
R2366 VTAIL.n67 VTAIL.n14 3.49141
R2367 VTAIL.n90 VTAIL.n2 3.49141
R2368 VTAIL.n142 VTAIL.n141 3.49141
R2369 VTAIL.n165 VTAIL.n112 3.49141
R2370 VTAIL.n188 VTAIL.n100 3.49141
R2371 VTAIL.n240 VTAIL.n239 3.49141
R2372 VTAIL.n263 VTAIL.n210 3.49141
R2373 VTAIL.n286 VTAIL.n198 3.49141
R2374 VTAIL.n678 VTAIL.n590 3.49141
R2375 VTAIL.n657 VTAIL.n604 3.49141
R2376 VTAIL.n634 VTAIL.n633 3.49141
R2377 VTAIL.n580 VTAIL.n492 3.49141
R2378 VTAIL.n559 VTAIL.n506 3.49141
R2379 VTAIL.n536 VTAIL.n535 3.49141
R2380 VTAIL.n482 VTAIL.n394 3.49141
R2381 VTAIL.n461 VTAIL.n408 3.49141
R2382 VTAIL.n438 VTAIL.n437 3.49141
R2383 VTAIL.n384 VTAIL.n296 3.49141
R2384 VTAIL.n363 VTAIL.n310 3.49141
R2385 VTAIL.n340 VTAIL.n339 3.49141
R2386 VTAIL.n726 VTAIL.n712 2.71565
R2387 VTAIL.n754 VTAIL.n698 2.71565
R2388 VTAIL.n775 VTAIL.n690 2.71565
R2389 VTAIL.n40 VTAIL.n26 2.71565
R2390 VTAIL.n68 VTAIL.n12 2.71565
R2391 VTAIL.n89 VTAIL.n4 2.71565
R2392 VTAIL.n138 VTAIL.n124 2.71565
R2393 VTAIL.n166 VTAIL.n110 2.71565
R2394 VTAIL.n187 VTAIL.n102 2.71565
R2395 VTAIL.n236 VTAIL.n222 2.71565
R2396 VTAIL.n264 VTAIL.n208 2.71565
R2397 VTAIL.n285 VTAIL.n200 2.71565
R2398 VTAIL.n677 VTAIL.n592 2.71565
R2399 VTAIL.n658 VTAIL.n602 2.71565
R2400 VTAIL.n630 VTAIL.n616 2.71565
R2401 VTAIL.n579 VTAIL.n494 2.71565
R2402 VTAIL.n560 VTAIL.n504 2.71565
R2403 VTAIL.n532 VTAIL.n518 2.71565
R2404 VTAIL.n481 VTAIL.n396 2.71565
R2405 VTAIL.n462 VTAIL.n406 2.71565
R2406 VTAIL.n434 VTAIL.n420 2.71565
R2407 VTAIL.n383 VTAIL.n298 2.71565
R2408 VTAIL.n364 VTAIL.n308 2.71565
R2409 VTAIL.n336 VTAIL.n322 2.71565
R2410 VTAIL.n725 VTAIL.n714 1.93989
R2411 VTAIL.n759 VTAIL.n757 1.93989
R2412 VTAIL.n772 VTAIL.n771 1.93989
R2413 VTAIL.n39 VTAIL.n28 1.93989
R2414 VTAIL.n73 VTAIL.n71 1.93989
R2415 VTAIL.n86 VTAIL.n85 1.93989
R2416 VTAIL.n137 VTAIL.n126 1.93989
R2417 VTAIL.n171 VTAIL.n169 1.93989
R2418 VTAIL.n184 VTAIL.n183 1.93989
R2419 VTAIL.n235 VTAIL.n224 1.93989
R2420 VTAIL.n269 VTAIL.n267 1.93989
R2421 VTAIL.n282 VTAIL.n281 1.93989
R2422 VTAIL.n674 VTAIL.n673 1.93989
R2423 VTAIL.n662 VTAIL.n661 1.93989
R2424 VTAIL.n629 VTAIL.n618 1.93989
R2425 VTAIL.n576 VTAIL.n575 1.93989
R2426 VTAIL.n564 VTAIL.n563 1.93989
R2427 VTAIL.n531 VTAIL.n520 1.93989
R2428 VTAIL.n478 VTAIL.n477 1.93989
R2429 VTAIL.n466 VTAIL.n465 1.93989
R2430 VTAIL.n433 VTAIL.n422 1.93989
R2431 VTAIL.n380 VTAIL.n379 1.93989
R2432 VTAIL.n368 VTAIL.n367 1.93989
R2433 VTAIL.n335 VTAIL.n324 1.93989
R2434 VTAIL.n489 VTAIL.n391 1.4574
R2435 VTAIL.n685 VTAIL.n587 1.4574
R2436 VTAIL.n293 VTAIL.n195 1.4574
R2437 VTAIL.n722 VTAIL.n721 1.16414
R2438 VTAIL.n758 VTAIL.n696 1.16414
R2439 VTAIL.n768 VTAIL.n692 1.16414
R2440 VTAIL.n36 VTAIL.n35 1.16414
R2441 VTAIL.n72 VTAIL.n10 1.16414
R2442 VTAIL.n82 VTAIL.n6 1.16414
R2443 VTAIL.n134 VTAIL.n133 1.16414
R2444 VTAIL.n170 VTAIL.n108 1.16414
R2445 VTAIL.n180 VTAIL.n104 1.16414
R2446 VTAIL.n232 VTAIL.n231 1.16414
R2447 VTAIL.n268 VTAIL.n206 1.16414
R2448 VTAIL.n278 VTAIL.n202 1.16414
R2449 VTAIL.n670 VTAIL.n594 1.16414
R2450 VTAIL.n665 VTAIL.n599 1.16414
R2451 VTAIL.n626 VTAIL.n625 1.16414
R2452 VTAIL.n572 VTAIL.n496 1.16414
R2453 VTAIL.n567 VTAIL.n501 1.16414
R2454 VTAIL.n528 VTAIL.n527 1.16414
R2455 VTAIL.n474 VTAIL.n398 1.16414
R2456 VTAIL.n469 VTAIL.n403 1.16414
R2457 VTAIL.n430 VTAIL.n429 1.16414
R2458 VTAIL.n376 VTAIL.n300 1.16414
R2459 VTAIL.n371 VTAIL.n305 1.16414
R2460 VTAIL.n332 VTAIL.n331 1.16414
R2461 VTAIL VTAIL.n97 0.787138
R2462 VTAIL VTAIL.n783 0.670759
R2463 VTAIL.n587 VTAIL.n489 0.470328
R2464 VTAIL.n195 VTAIL.n97 0.470328
R2465 VTAIL.n718 VTAIL.n716 0.388379
R2466 VTAIL.n764 VTAIL.n763 0.388379
R2467 VTAIL.n767 VTAIL.n694 0.388379
R2468 VTAIL.n32 VTAIL.n30 0.388379
R2469 VTAIL.n78 VTAIL.n77 0.388379
R2470 VTAIL.n81 VTAIL.n8 0.388379
R2471 VTAIL.n130 VTAIL.n128 0.388379
R2472 VTAIL.n176 VTAIL.n175 0.388379
R2473 VTAIL.n179 VTAIL.n106 0.388379
R2474 VTAIL.n228 VTAIL.n226 0.388379
R2475 VTAIL.n274 VTAIL.n273 0.388379
R2476 VTAIL.n277 VTAIL.n204 0.388379
R2477 VTAIL.n669 VTAIL.n596 0.388379
R2478 VTAIL.n666 VTAIL.n598 0.388379
R2479 VTAIL.n622 VTAIL.n620 0.388379
R2480 VTAIL.n571 VTAIL.n498 0.388379
R2481 VTAIL.n568 VTAIL.n500 0.388379
R2482 VTAIL.n524 VTAIL.n522 0.388379
R2483 VTAIL.n473 VTAIL.n400 0.388379
R2484 VTAIL.n470 VTAIL.n402 0.388379
R2485 VTAIL.n426 VTAIL.n424 0.388379
R2486 VTAIL.n375 VTAIL.n302 0.388379
R2487 VTAIL.n372 VTAIL.n304 0.388379
R2488 VTAIL.n328 VTAIL.n326 0.388379
R2489 VTAIL.n723 VTAIL.n715 0.155672
R2490 VTAIL.n724 VTAIL.n723 0.155672
R2491 VTAIL.n724 VTAIL.n711 0.155672
R2492 VTAIL.n731 VTAIL.n711 0.155672
R2493 VTAIL.n732 VTAIL.n731 0.155672
R2494 VTAIL.n732 VTAIL.n707 0.155672
R2495 VTAIL.n739 VTAIL.n707 0.155672
R2496 VTAIL.n740 VTAIL.n739 0.155672
R2497 VTAIL.n740 VTAIL.n703 0.155672
R2498 VTAIL.n747 VTAIL.n703 0.155672
R2499 VTAIL.n748 VTAIL.n747 0.155672
R2500 VTAIL.n748 VTAIL.n699 0.155672
R2501 VTAIL.n755 VTAIL.n699 0.155672
R2502 VTAIL.n756 VTAIL.n755 0.155672
R2503 VTAIL.n756 VTAIL.n695 0.155672
R2504 VTAIL.n765 VTAIL.n695 0.155672
R2505 VTAIL.n766 VTAIL.n765 0.155672
R2506 VTAIL.n766 VTAIL.n691 0.155672
R2507 VTAIL.n773 VTAIL.n691 0.155672
R2508 VTAIL.n774 VTAIL.n773 0.155672
R2509 VTAIL.n774 VTAIL.n687 0.155672
R2510 VTAIL.n781 VTAIL.n687 0.155672
R2511 VTAIL.n37 VTAIL.n29 0.155672
R2512 VTAIL.n38 VTAIL.n37 0.155672
R2513 VTAIL.n38 VTAIL.n25 0.155672
R2514 VTAIL.n45 VTAIL.n25 0.155672
R2515 VTAIL.n46 VTAIL.n45 0.155672
R2516 VTAIL.n46 VTAIL.n21 0.155672
R2517 VTAIL.n53 VTAIL.n21 0.155672
R2518 VTAIL.n54 VTAIL.n53 0.155672
R2519 VTAIL.n54 VTAIL.n17 0.155672
R2520 VTAIL.n61 VTAIL.n17 0.155672
R2521 VTAIL.n62 VTAIL.n61 0.155672
R2522 VTAIL.n62 VTAIL.n13 0.155672
R2523 VTAIL.n69 VTAIL.n13 0.155672
R2524 VTAIL.n70 VTAIL.n69 0.155672
R2525 VTAIL.n70 VTAIL.n9 0.155672
R2526 VTAIL.n79 VTAIL.n9 0.155672
R2527 VTAIL.n80 VTAIL.n79 0.155672
R2528 VTAIL.n80 VTAIL.n5 0.155672
R2529 VTAIL.n87 VTAIL.n5 0.155672
R2530 VTAIL.n88 VTAIL.n87 0.155672
R2531 VTAIL.n88 VTAIL.n1 0.155672
R2532 VTAIL.n95 VTAIL.n1 0.155672
R2533 VTAIL.n135 VTAIL.n127 0.155672
R2534 VTAIL.n136 VTAIL.n135 0.155672
R2535 VTAIL.n136 VTAIL.n123 0.155672
R2536 VTAIL.n143 VTAIL.n123 0.155672
R2537 VTAIL.n144 VTAIL.n143 0.155672
R2538 VTAIL.n144 VTAIL.n119 0.155672
R2539 VTAIL.n151 VTAIL.n119 0.155672
R2540 VTAIL.n152 VTAIL.n151 0.155672
R2541 VTAIL.n152 VTAIL.n115 0.155672
R2542 VTAIL.n159 VTAIL.n115 0.155672
R2543 VTAIL.n160 VTAIL.n159 0.155672
R2544 VTAIL.n160 VTAIL.n111 0.155672
R2545 VTAIL.n167 VTAIL.n111 0.155672
R2546 VTAIL.n168 VTAIL.n167 0.155672
R2547 VTAIL.n168 VTAIL.n107 0.155672
R2548 VTAIL.n177 VTAIL.n107 0.155672
R2549 VTAIL.n178 VTAIL.n177 0.155672
R2550 VTAIL.n178 VTAIL.n103 0.155672
R2551 VTAIL.n185 VTAIL.n103 0.155672
R2552 VTAIL.n186 VTAIL.n185 0.155672
R2553 VTAIL.n186 VTAIL.n99 0.155672
R2554 VTAIL.n193 VTAIL.n99 0.155672
R2555 VTAIL.n233 VTAIL.n225 0.155672
R2556 VTAIL.n234 VTAIL.n233 0.155672
R2557 VTAIL.n234 VTAIL.n221 0.155672
R2558 VTAIL.n241 VTAIL.n221 0.155672
R2559 VTAIL.n242 VTAIL.n241 0.155672
R2560 VTAIL.n242 VTAIL.n217 0.155672
R2561 VTAIL.n249 VTAIL.n217 0.155672
R2562 VTAIL.n250 VTAIL.n249 0.155672
R2563 VTAIL.n250 VTAIL.n213 0.155672
R2564 VTAIL.n257 VTAIL.n213 0.155672
R2565 VTAIL.n258 VTAIL.n257 0.155672
R2566 VTAIL.n258 VTAIL.n209 0.155672
R2567 VTAIL.n265 VTAIL.n209 0.155672
R2568 VTAIL.n266 VTAIL.n265 0.155672
R2569 VTAIL.n266 VTAIL.n205 0.155672
R2570 VTAIL.n275 VTAIL.n205 0.155672
R2571 VTAIL.n276 VTAIL.n275 0.155672
R2572 VTAIL.n276 VTAIL.n201 0.155672
R2573 VTAIL.n283 VTAIL.n201 0.155672
R2574 VTAIL.n284 VTAIL.n283 0.155672
R2575 VTAIL.n284 VTAIL.n197 0.155672
R2576 VTAIL.n291 VTAIL.n197 0.155672
R2577 VTAIL.n683 VTAIL.n589 0.155672
R2578 VTAIL.n676 VTAIL.n589 0.155672
R2579 VTAIL.n676 VTAIL.n675 0.155672
R2580 VTAIL.n675 VTAIL.n593 0.155672
R2581 VTAIL.n668 VTAIL.n593 0.155672
R2582 VTAIL.n668 VTAIL.n667 0.155672
R2583 VTAIL.n667 VTAIL.n597 0.155672
R2584 VTAIL.n660 VTAIL.n597 0.155672
R2585 VTAIL.n660 VTAIL.n659 0.155672
R2586 VTAIL.n659 VTAIL.n603 0.155672
R2587 VTAIL.n652 VTAIL.n603 0.155672
R2588 VTAIL.n652 VTAIL.n651 0.155672
R2589 VTAIL.n651 VTAIL.n607 0.155672
R2590 VTAIL.n644 VTAIL.n607 0.155672
R2591 VTAIL.n644 VTAIL.n643 0.155672
R2592 VTAIL.n643 VTAIL.n611 0.155672
R2593 VTAIL.n636 VTAIL.n611 0.155672
R2594 VTAIL.n636 VTAIL.n635 0.155672
R2595 VTAIL.n635 VTAIL.n615 0.155672
R2596 VTAIL.n628 VTAIL.n615 0.155672
R2597 VTAIL.n628 VTAIL.n627 0.155672
R2598 VTAIL.n627 VTAIL.n619 0.155672
R2599 VTAIL.n585 VTAIL.n491 0.155672
R2600 VTAIL.n578 VTAIL.n491 0.155672
R2601 VTAIL.n578 VTAIL.n577 0.155672
R2602 VTAIL.n577 VTAIL.n495 0.155672
R2603 VTAIL.n570 VTAIL.n495 0.155672
R2604 VTAIL.n570 VTAIL.n569 0.155672
R2605 VTAIL.n569 VTAIL.n499 0.155672
R2606 VTAIL.n562 VTAIL.n499 0.155672
R2607 VTAIL.n562 VTAIL.n561 0.155672
R2608 VTAIL.n561 VTAIL.n505 0.155672
R2609 VTAIL.n554 VTAIL.n505 0.155672
R2610 VTAIL.n554 VTAIL.n553 0.155672
R2611 VTAIL.n553 VTAIL.n509 0.155672
R2612 VTAIL.n546 VTAIL.n509 0.155672
R2613 VTAIL.n546 VTAIL.n545 0.155672
R2614 VTAIL.n545 VTAIL.n513 0.155672
R2615 VTAIL.n538 VTAIL.n513 0.155672
R2616 VTAIL.n538 VTAIL.n537 0.155672
R2617 VTAIL.n537 VTAIL.n517 0.155672
R2618 VTAIL.n530 VTAIL.n517 0.155672
R2619 VTAIL.n530 VTAIL.n529 0.155672
R2620 VTAIL.n529 VTAIL.n521 0.155672
R2621 VTAIL.n487 VTAIL.n393 0.155672
R2622 VTAIL.n480 VTAIL.n393 0.155672
R2623 VTAIL.n480 VTAIL.n479 0.155672
R2624 VTAIL.n479 VTAIL.n397 0.155672
R2625 VTAIL.n472 VTAIL.n397 0.155672
R2626 VTAIL.n472 VTAIL.n471 0.155672
R2627 VTAIL.n471 VTAIL.n401 0.155672
R2628 VTAIL.n464 VTAIL.n401 0.155672
R2629 VTAIL.n464 VTAIL.n463 0.155672
R2630 VTAIL.n463 VTAIL.n407 0.155672
R2631 VTAIL.n456 VTAIL.n407 0.155672
R2632 VTAIL.n456 VTAIL.n455 0.155672
R2633 VTAIL.n455 VTAIL.n411 0.155672
R2634 VTAIL.n448 VTAIL.n411 0.155672
R2635 VTAIL.n448 VTAIL.n447 0.155672
R2636 VTAIL.n447 VTAIL.n415 0.155672
R2637 VTAIL.n440 VTAIL.n415 0.155672
R2638 VTAIL.n440 VTAIL.n439 0.155672
R2639 VTAIL.n439 VTAIL.n419 0.155672
R2640 VTAIL.n432 VTAIL.n419 0.155672
R2641 VTAIL.n432 VTAIL.n431 0.155672
R2642 VTAIL.n431 VTAIL.n423 0.155672
R2643 VTAIL.n389 VTAIL.n295 0.155672
R2644 VTAIL.n382 VTAIL.n295 0.155672
R2645 VTAIL.n382 VTAIL.n381 0.155672
R2646 VTAIL.n381 VTAIL.n299 0.155672
R2647 VTAIL.n374 VTAIL.n299 0.155672
R2648 VTAIL.n374 VTAIL.n373 0.155672
R2649 VTAIL.n373 VTAIL.n303 0.155672
R2650 VTAIL.n366 VTAIL.n303 0.155672
R2651 VTAIL.n366 VTAIL.n365 0.155672
R2652 VTAIL.n365 VTAIL.n309 0.155672
R2653 VTAIL.n358 VTAIL.n309 0.155672
R2654 VTAIL.n358 VTAIL.n357 0.155672
R2655 VTAIL.n357 VTAIL.n313 0.155672
R2656 VTAIL.n350 VTAIL.n313 0.155672
R2657 VTAIL.n350 VTAIL.n349 0.155672
R2658 VTAIL.n349 VTAIL.n317 0.155672
R2659 VTAIL.n342 VTAIL.n317 0.155672
R2660 VTAIL.n342 VTAIL.n341 0.155672
R2661 VTAIL.n341 VTAIL.n321 0.155672
R2662 VTAIL.n334 VTAIL.n321 0.155672
R2663 VTAIL.n334 VTAIL.n333 0.155672
R2664 VTAIL.n333 VTAIL.n325 0.155672
R2665 VN.n0 VN.t3 348.219
R2666 VN.n1 VN.t2 348.219
R2667 VN.n0 VN.t1 347.986
R2668 VN.n1 VN.t0 347.986
R2669 VN VN.n1 64.7087
R2670 VN VN.n0 17.6897
R2671 VDD2.n2 VDD2.n0 103.263
R2672 VDD2.n2 VDD2.n1 60.1001
R2673 VDD2.n1 VDD2.t3 1.13258
R2674 VDD2.n1 VDD2.t1 1.13258
R2675 VDD2.n0 VDD2.t0 1.13258
R2676 VDD2.n0 VDD2.t2 1.13258
R2677 VDD2 VDD2.n2 0.0586897
C0 VN VDD2 5.79485f
C1 VTAIL VDD2 7.40502f
C2 VN VTAIL 5.28107f
C3 VDD1 VP 5.96195f
C4 VDD2 VP 0.315217f
C5 VN VP 6.31133f
C6 VDD1 VDD2 0.723287f
C7 VTAIL VP 5.29517f
C8 VN VDD1 0.147694f
C9 VTAIL VDD1 7.35913f
C10 VDD2 B 3.497063f
C11 VDD1 B 7.85878f
C12 VTAIL B 12.488223f
C13 VN B 9.2796f
C14 VP B 6.659454f
C15 VDD2.t0 B 0.369541f
C16 VDD2.t2 B 0.369541f
C17 VDD2.n0 B 4.17871f
C18 VDD2.t3 B 0.369541f
C19 VDD2.t1 B 0.369541f
C20 VDD2.n1 B 3.36154f
C21 VDD2.n2 B 4.05031f
C22 VN.t3 B 2.47581f
C23 VN.t1 B 2.47516f
C24 VN.n0 B 1.77407f
C25 VN.t2 B 2.47581f
C26 VN.t0 B 2.47516f
C27 VN.n1 B 3.19907f
C28 VTAIL.n0 B 0.020609f
C29 VTAIL.n1 B 0.015172f
C30 VTAIL.n2 B 0.008153f
C31 VTAIL.n3 B 0.01927f
C32 VTAIL.n4 B 0.008632f
C33 VTAIL.n5 B 0.015172f
C34 VTAIL.n6 B 0.008153f
C35 VTAIL.n7 B 0.01927f
C36 VTAIL.n8 B 0.008392f
C37 VTAIL.n9 B 0.015172f
C38 VTAIL.n10 B 0.008632f
C39 VTAIL.n11 B 0.01927f
C40 VTAIL.n12 B 0.008632f
C41 VTAIL.n13 B 0.015172f
C42 VTAIL.n14 B 0.008153f
C43 VTAIL.n15 B 0.01927f
C44 VTAIL.n16 B 0.008632f
C45 VTAIL.n17 B 0.015172f
C46 VTAIL.n18 B 0.008153f
C47 VTAIL.n19 B 0.01927f
C48 VTAIL.n20 B 0.008632f
C49 VTAIL.n21 B 0.015172f
C50 VTAIL.n22 B 0.008153f
C51 VTAIL.n23 B 0.01927f
C52 VTAIL.n24 B 0.008632f
C53 VTAIL.n25 B 0.015172f
C54 VTAIL.n26 B 0.008153f
C55 VTAIL.n27 B 0.01927f
C56 VTAIL.n28 B 0.008632f
C57 VTAIL.n29 B 1.16023f
C58 VTAIL.n30 B 0.008153f
C59 VTAIL.t1 B 0.031903f
C60 VTAIL.n31 B 0.108425f
C61 VTAIL.n32 B 0.011383f
C62 VTAIL.n33 B 0.014452f
C63 VTAIL.n34 B 0.01927f
C64 VTAIL.n35 B 0.008632f
C65 VTAIL.n36 B 0.008153f
C66 VTAIL.n37 B 0.015172f
C67 VTAIL.n38 B 0.015172f
C68 VTAIL.n39 B 0.008153f
C69 VTAIL.n40 B 0.008632f
C70 VTAIL.n41 B 0.01927f
C71 VTAIL.n42 B 0.01927f
C72 VTAIL.n43 B 0.008632f
C73 VTAIL.n44 B 0.008153f
C74 VTAIL.n45 B 0.015172f
C75 VTAIL.n46 B 0.015172f
C76 VTAIL.n47 B 0.008153f
C77 VTAIL.n48 B 0.008632f
C78 VTAIL.n49 B 0.01927f
C79 VTAIL.n50 B 0.01927f
C80 VTAIL.n51 B 0.008632f
C81 VTAIL.n52 B 0.008153f
C82 VTAIL.n53 B 0.015172f
C83 VTAIL.n54 B 0.015172f
C84 VTAIL.n55 B 0.008153f
C85 VTAIL.n56 B 0.008632f
C86 VTAIL.n57 B 0.01927f
C87 VTAIL.n58 B 0.01927f
C88 VTAIL.n59 B 0.008632f
C89 VTAIL.n60 B 0.008153f
C90 VTAIL.n61 B 0.015172f
C91 VTAIL.n62 B 0.015172f
C92 VTAIL.n63 B 0.008153f
C93 VTAIL.n64 B 0.008632f
C94 VTAIL.n65 B 0.01927f
C95 VTAIL.n66 B 0.01927f
C96 VTAIL.n67 B 0.008632f
C97 VTAIL.n68 B 0.008153f
C98 VTAIL.n69 B 0.015172f
C99 VTAIL.n70 B 0.015172f
C100 VTAIL.n71 B 0.008153f
C101 VTAIL.n72 B 0.008153f
C102 VTAIL.n73 B 0.008632f
C103 VTAIL.n74 B 0.01927f
C104 VTAIL.n75 B 0.01927f
C105 VTAIL.n76 B 0.01927f
C106 VTAIL.n77 B 0.008392f
C107 VTAIL.n78 B 0.008153f
C108 VTAIL.n79 B 0.015172f
C109 VTAIL.n80 B 0.015172f
C110 VTAIL.n81 B 0.008153f
C111 VTAIL.n82 B 0.008632f
C112 VTAIL.n83 B 0.01927f
C113 VTAIL.n84 B 0.01927f
C114 VTAIL.n85 B 0.008632f
C115 VTAIL.n86 B 0.008153f
C116 VTAIL.n87 B 0.015172f
C117 VTAIL.n88 B 0.015172f
C118 VTAIL.n89 B 0.008153f
C119 VTAIL.n90 B 0.008632f
C120 VTAIL.n91 B 0.01927f
C121 VTAIL.n92 B 0.040449f
C122 VTAIL.n93 B 0.008632f
C123 VTAIL.n94 B 0.008153f
C124 VTAIL.n95 B 0.034447f
C125 VTAIL.n96 B 0.022483f
C126 VTAIL.n97 B 0.074031f
C127 VTAIL.n98 B 0.020609f
C128 VTAIL.n99 B 0.015172f
C129 VTAIL.n100 B 0.008153f
C130 VTAIL.n101 B 0.01927f
C131 VTAIL.n102 B 0.008632f
C132 VTAIL.n103 B 0.015172f
C133 VTAIL.n104 B 0.008153f
C134 VTAIL.n105 B 0.01927f
C135 VTAIL.n106 B 0.008392f
C136 VTAIL.n107 B 0.015172f
C137 VTAIL.n108 B 0.008632f
C138 VTAIL.n109 B 0.01927f
C139 VTAIL.n110 B 0.008632f
C140 VTAIL.n111 B 0.015172f
C141 VTAIL.n112 B 0.008153f
C142 VTAIL.n113 B 0.01927f
C143 VTAIL.n114 B 0.008632f
C144 VTAIL.n115 B 0.015172f
C145 VTAIL.n116 B 0.008153f
C146 VTAIL.n117 B 0.01927f
C147 VTAIL.n118 B 0.008632f
C148 VTAIL.n119 B 0.015172f
C149 VTAIL.n120 B 0.008153f
C150 VTAIL.n121 B 0.01927f
C151 VTAIL.n122 B 0.008632f
C152 VTAIL.n123 B 0.015172f
C153 VTAIL.n124 B 0.008153f
C154 VTAIL.n125 B 0.01927f
C155 VTAIL.n126 B 0.008632f
C156 VTAIL.n127 B 1.16023f
C157 VTAIL.n128 B 0.008153f
C158 VTAIL.t4 B 0.031903f
C159 VTAIL.n129 B 0.108425f
C160 VTAIL.n130 B 0.011383f
C161 VTAIL.n131 B 0.014452f
C162 VTAIL.n132 B 0.01927f
C163 VTAIL.n133 B 0.008632f
C164 VTAIL.n134 B 0.008153f
C165 VTAIL.n135 B 0.015172f
C166 VTAIL.n136 B 0.015172f
C167 VTAIL.n137 B 0.008153f
C168 VTAIL.n138 B 0.008632f
C169 VTAIL.n139 B 0.01927f
C170 VTAIL.n140 B 0.01927f
C171 VTAIL.n141 B 0.008632f
C172 VTAIL.n142 B 0.008153f
C173 VTAIL.n143 B 0.015172f
C174 VTAIL.n144 B 0.015172f
C175 VTAIL.n145 B 0.008153f
C176 VTAIL.n146 B 0.008632f
C177 VTAIL.n147 B 0.01927f
C178 VTAIL.n148 B 0.01927f
C179 VTAIL.n149 B 0.008632f
C180 VTAIL.n150 B 0.008153f
C181 VTAIL.n151 B 0.015172f
C182 VTAIL.n152 B 0.015172f
C183 VTAIL.n153 B 0.008153f
C184 VTAIL.n154 B 0.008632f
C185 VTAIL.n155 B 0.01927f
C186 VTAIL.n156 B 0.01927f
C187 VTAIL.n157 B 0.008632f
C188 VTAIL.n158 B 0.008153f
C189 VTAIL.n159 B 0.015172f
C190 VTAIL.n160 B 0.015172f
C191 VTAIL.n161 B 0.008153f
C192 VTAIL.n162 B 0.008632f
C193 VTAIL.n163 B 0.01927f
C194 VTAIL.n164 B 0.01927f
C195 VTAIL.n165 B 0.008632f
C196 VTAIL.n166 B 0.008153f
C197 VTAIL.n167 B 0.015172f
C198 VTAIL.n168 B 0.015172f
C199 VTAIL.n169 B 0.008153f
C200 VTAIL.n170 B 0.008153f
C201 VTAIL.n171 B 0.008632f
C202 VTAIL.n172 B 0.01927f
C203 VTAIL.n173 B 0.01927f
C204 VTAIL.n174 B 0.01927f
C205 VTAIL.n175 B 0.008392f
C206 VTAIL.n176 B 0.008153f
C207 VTAIL.n177 B 0.015172f
C208 VTAIL.n178 B 0.015172f
C209 VTAIL.n179 B 0.008153f
C210 VTAIL.n180 B 0.008632f
C211 VTAIL.n181 B 0.01927f
C212 VTAIL.n182 B 0.01927f
C213 VTAIL.n183 B 0.008632f
C214 VTAIL.n184 B 0.008153f
C215 VTAIL.n185 B 0.015172f
C216 VTAIL.n186 B 0.015172f
C217 VTAIL.n187 B 0.008153f
C218 VTAIL.n188 B 0.008632f
C219 VTAIL.n189 B 0.01927f
C220 VTAIL.n190 B 0.040449f
C221 VTAIL.n191 B 0.008632f
C222 VTAIL.n192 B 0.008153f
C223 VTAIL.n193 B 0.034447f
C224 VTAIL.n194 B 0.022483f
C225 VTAIL.n195 B 0.106798f
C226 VTAIL.n196 B 0.020609f
C227 VTAIL.n197 B 0.015172f
C228 VTAIL.n198 B 0.008153f
C229 VTAIL.n199 B 0.01927f
C230 VTAIL.n200 B 0.008632f
C231 VTAIL.n201 B 0.015172f
C232 VTAIL.n202 B 0.008153f
C233 VTAIL.n203 B 0.01927f
C234 VTAIL.n204 B 0.008392f
C235 VTAIL.n205 B 0.015172f
C236 VTAIL.n206 B 0.008632f
C237 VTAIL.n207 B 0.01927f
C238 VTAIL.n208 B 0.008632f
C239 VTAIL.n209 B 0.015172f
C240 VTAIL.n210 B 0.008153f
C241 VTAIL.n211 B 0.01927f
C242 VTAIL.n212 B 0.008632f
C243 VTAIL.n213 B 0.015172f
C244 VTAIL.n214 B 0.008153f
C245 VTAIL.n215 B 0.01927f
C246 VTAIL.n216 B 0.008632f
C247 VTAIL.n217 B 0.015172f
C248 VTAIL.n218 B 0.008153f
C249 VTAIL.n219 B 0.01927f
C250 VTAIL.n220 B 0.008632f
C251 VTAIL.n221 B 0.015172f
C252 VTAIL.n222 B 0.008153f
C253 VTAIL.n223 B 0.01927f
C254 VTAIL.n224 B 0.008632f
C255 VTAIL.n225 B 1.16023f
C256 VTAIL.n226 B 0.008153f
C257 VTAIL.t7 B 0.031903f
C258 VTAIL.n227 B 0.108425f
C259 VTAIL.n228 B 0.011383f
C260 VTAIL.n229 B 0.014452f
C261 VTAIL.n230 B 0.01927f
C262 VTAIL.n231 B 0.008632f
C263 VTAIL.n232 B 0.008153f
C264 VTAIL.n233 B 0.015172f
C265 VTAIL.n234 B 0.015172f
C266 VTAIL.n235 B 0.008153f
C267 VTAIL.n236 B 0.008632f
C268 VTAIL.n237 B 0.01927f
C269 VTAIL.n238 B 0.01927f
C270 VTAIL.n239 B 0.008632f
C271 VTAIL.n240 B 0.008153f
C272 VTAIL.n241 B 0.015172f
C273 VTAIL.n242 B 0.015172f
C274 VTAIL.n243 B 0.008153f
C275 VTAIL.n244 B 0.008632f
C276 VTAIL.n245 B 0.01927f
C277 VTAIL.n246 B 0.01927f
C278 VTAIL.n247 B 0.008632f
C279 VTAIL.n248 B 0.008153f
C280 VTAIL.n249 B 0.015172f
C281 VTAIL.n250 B 0.015172f
C282 VTAIL.n251 B 0.008153f
C283 VTAIL.n252 B 0.008632f
C284 VTAIL.n253 B 0.01927f
C285 VTAIL.n254 B 0.01927f
C286 VTAIL.n255 B 0.008632f
C287 VTAIL.n256 B 0.008153f
C288 VTAIL.n257 B 0.015172f
C289 VTAIL.n258 B 0.015172f
C290 VTAIL.n259 B 0.008153f
C291 VTAIL.n260 B 0.008632f
C292 VTAIL.n261 B 0.01927f
C293 VTAIL.n262 B 0.01927f
C294 VTAIL.n263 B 0.008632f
C295 VTAIL.n264 B 0.008153f
C296 VTAIL.n265 B 0.015172f
C297 VTAIL.n266 B 0.015172f
C298 VTAIL.n267 B 0.008153f
C299 VTAIL.n268 B 0.008153f
C300 VTAIL.n269 B 0.008632f
C301 VTAIL.n270 B 0.01927f
C302 VTAIL.n271 B 0.01927f
C303 VTAIL.n272 B 0.01927f
C304 VTAIL.n273 B 0.008392f
C305 VTAIL.n274 B 0.008153f
C306 VTAIL.n275 B 0.015172f
C307 VTAIL.n276 B 0.015172f
C308 VTAIL.n277 B 0.008153f
C309 VTAIL.n278 B 0.008632f
C310 VTAIL.n279 B 0.01927f
C311 VTAIL.n280 B 0.01927f
C312 VTAIL.n281 B 0.008632f
C313 VTAIL.n282 B 0.008153f
C314 VTAIL.n283 B 0.015172f
C315 VTAIL.n284 B 0.015172f
C316 VTAIL.n285 B 0.008153f
C317 VTAIL.n286 B 0.008632f
C318 VTAIL.n287 B 0.01927f
C319 VTAIL.n288 B 0.040449f
C320 VTAIL.n289 B 0.008632f
C321 VTAIL.n290 B 0.008153f
C322 VTAIL.n291 B 0.034447f
C323 VTAIL.n292 B 0.022483f
C324 VTAIL.n293 B 1.09823f
C325 VTAIL.n294 B 0.020609f
C326 VTAIL.n295 B 0.015172f
C327 VTAIL.n296 B 0.008153f
C328 VTAIL.n297 B 0.01927f
C329 VTAIL.n298 B 0.008632f
C330 VTAIL.n299 B 0.015172f
C331 VTAIL.n300 B 0.008153f
C332 VTAIL.n301 B 0.01927f
C333 VTAIL.n302 B 0.008392f
C334 VTAIL.n303 B 0.015172f
C335 VTAIL.n304 B 0.008392f
C336 VTAIL.n305 B 0.008153f
C337 VTAIL.n306 B 0.01927f
C338 VTAIL.n307 B 0.01927f
C339 VTAIL.n308 B 0.008632f
C340 VTAIL.n309 B 0.015172f
C341 VTAIL.n310 B 0.008153f
C342 VTAIL.n311 B 0.01927f
C343 VTAIL.n312 B 0.008632f
C344 VTAIL.n313 B 0.015172f
C345 VTAIL.n314 B 0.008153f
C346 VTAIL.n315 B 0.01927f
C347 VTAIL.n316 B 0.008632f
C348 VTAIL.n317 B 0.015172f
C349 VTAIL.n318 B 0.008153f
C350 VTAIL.n319 B 0.01927f
C351 VTAIL.n320 B 0.008632f
C352 VTAIL.n321 B 0.015172f
C353 VTAIL.n322 B 0.008153f
C354 VTAIL.n323 B 0.01927f
C355 VTAIL.n324 B 0.008632f
C356 VTAIL.n325 B 1.16023f
C357 VTAIL.n326 B 0.008153f
C358 VTAIL.t3 B 0.031903f
C359 VTAIL.n327 B 0.108425f
C360 VTAIL.n328 B 0.011383f
C361 VTAIL.n329 B 0.014452f
C362 VTAIL.n330 B 0.01927f
C363 VTAIL.n331 B 0.008632f
C364 VTAIL.n332 B 0.008153f
C365 VTAIL.n333 B 0.015172f
C366 VTAIL.n334 B 0.015172f
C367 VTAIL.n335 B 0.008153f
C368 VTAIL.n336 B 0.008632f
C369 VTAIL.n337 B 0.01927f
C370 VTAIL.n338 B 0.01927f
C371 VTAIL.n339 B 0.008632f
C372 VTAIL.n340 B 0.008153f
C373 VTAIL.n341 B 0.015172f
C374 VTAIL.n342 B 0.015172f
C375 VTAIL.n343 B 0.008153f
C376 VTAIL.n344 B 0.008632f
C377 VTAIL.n345 B 0.01927f
C378 VTAIL.n346 B 0.01927f
C379 VTAIL.n347 B 0.008632f
C380 VTAIL.n348 B 0.008153f
C381 VTAIL.n349 B 0.015172f
C382 VTAIL.n350 B 0.015172f
C383 VTAIL.n351 B 0.008153f
C384 VTAIL.n352 B 0.008632f
C385 VTAIL.n353 B 0.01927f
C386 VTAIL.n354 B 0.01927f
C387 VTAIL.n355 B 0.008632f
C388 VTAIL.n356 B 0.008153f
C389 VTAIL.n357 B 0.015172f
C390 VTAIL.n358 B 0.015172f
C391 VTAIL.n359 B 0.008153f
C392 VTAIL.n360 B 0.008632f
C393 VTAIL.n361 B 0.01927f
C394 VTAIL.n362 B 0.01927f
C395 VTAIL.n363 B 0.008632f
C396 VTAIL.n364 B 0.008153f
C397 VTAIL.n365 B 0.015172f
C398 VTAIL.n366 B 0.015172f
C399 VTAIL.n367 B 0.008153f
C400 VTAIL.n368 B 0.008632f
C401 VTAIL.n369 B 0.01927f
C402 VTAIL.n370 B 0.01927f
C403 VTAIL.n371 B 0.008632f
C404 VTAIL.n372 B 0.008153f
C405 VTAIL.n373 B 0.015172f
C406 VTAIL.n374 B 0.015172f
C407 VTAIL.n375 B 0.008153f
C408 VTAIL.n376 B 0.008632f
C409 VTAIL.n377 B 0.01927f
C410 VTAIL.n378 B 0.01927f
C411 VTAIL.n379 B 0.008632f
C412 VTAIL.n380 B 0.008153f
C413 VTAIL.n381 B 0.015172f
C414 VTAIL.n382 B 0.015172f
C415 VTAIL.n383 B 0.008153f
C416 VTAIL.n384 B 0.008632f
C417 VTAIL.n385 B 0.01927f
C418 VTAIL.n386 B 0.040449f
C419 VTAIL.n387 B 0.008632f
C420 VTAIL.n388 B 0.008153f
C421 VTAIL.n389 B 0.034447f
C422 VTAIL.n390 B 0.022483f
C423 VTAIL.n391 B 1.09823f
C424 VTAIL.n392 B 0.020609f
C425 VTAIL.n393 B 0.015172f
C426 VTAIL.n394 B 0.008153f
C427 VTAIL.n395 B 0.01927f
C428 VTAIL.n396 B 0.008632f
C429 VTAIL.n397 B 0.015172f
C430 VTAIL.n398 B 0.008153f
C431 VTAIL.n399 B 0.01927f
C432 VTAIL.n400 B 0.008392f
C433 VTAIL.n401 B 0.015172f
C434 VTAIL.n402 B 0.008392f
C435 VTAIL.n403 B 0.008153f
C436 VTAIL.n404 B 0.01927f
C437 VTAIL.n405 B 0.01927f
C438 VTAIL.n406 B 0.008632f
C439 VTAIL.n407 B 0.015172f
C440 VTAIL.n408 B 0.008153f
C441 VTAIL.n409 B 0.01927f
C442 VTAIL.n410 B 0.008632f
C443 VTAIL.n411 B 0.015172f
C444 VTAIL.n412 B 0.008153f
C445 VTAIL.n413 B 0.01927f
C446 VTAIL.n414 B 0.008632f
C447 VTAIL.n415 B 0.015172f
C448 VTAIL.n416 B 0.008153f
C449 VTAIL.n417 B 0.01927f
C450 VTAIL.n418 B 0.008632f
C451 VTAIL.n419 B 0.015172f
C452 VTAIL.n420 B 0.008153f
C453 VTAIL.n421 B 0.01927f
C454 VTAIL.n422 B 0.008632f
C455 VTAIL.n423 B 1.16023f
C456 VTAIL.n424 B 0.008153f
C457 VTAIL.t0 B 0.031903f
C458 VTAIL.n425 B 0.108425f
C459 VTAIL.n426 B 0.011383f
C460 VTAIL.n427 B 0.014452f
C461 VTAIL.n428 B 0.01927f
C462 VTAIL.n429 B 0.008632f
C463 VTAIL.n430 B 0.008153f
C464 VTAIL.n431 B 0.015172f
C465 VTAIL.n432 B 0.015172f
C466 VTAIL.n433 B 0.008153f
C467 VTAIL.n434 B 0.008632f
C468 VTAIL.n435 B 0.01927f
C469 VTAIL.n436 B 0.01927f
C470 VTAIL.n437 B 0.008632f
C471 VTAIL.n438 B 0.008153f
C472 VTAIL.n439 B 0.015172f
C473 VTAIL.n440 B 0.015172f
C474 VTAIL.n441 B 0.008153f
C475 VTAIL.n442 B 0.008632f
C476 VTAIL.n443 B 0.01927f
C477 VTAIL.n444 B 0.01927f
C478 VTAIL.n445 B 0.008632f
C479 VTAIL.n446 B 0.008153f
C480 VTAIL.n447 B 0.015172f
C481 VTAIL.n448 B 0.015172f
C482 VTAIL.n449 B 0.008153f
C483 VTAIL.n450 B 0.008632f
C484 VTAIL.n451 B 0.01927f
C485 VTAIL.n452 B 0.01927f
C486 VTAIL.n453 B 0.008632f
C487 VTAIL.n454 B 0.008153f
C488 VTAIL.n455 B 0.015172f
C489 VTAIL.n456 B 0.015172f
C490 VTAIL.n457 B 0.008153f
C491 VTAIL.n458 B 0.008632f
C492 VTAIL.n459 B 0.01927f
C493 VTAIL.n460 B 0.01927f
C494 VTAIL.n461 B 0.008632f
C495 VTAIL.n462 B 0.008153f
C496 VTAIL.n463 B 0.015172f
C497 VTAIL.n464 B 0.015172f
C498 VTAIL.n465 B 0.008153f
C499 VTAIL.n466 B 0.008632f
C500 VTAIL.n467 B 0.01927f
C501 VTAIL.n468 B 0.01927f
C502 VTAIL.n469 B 0.008632f
C503 VTAIL.n470 B 0.008153f
C504 VTAIL.n471 B 0.015172f
C505 VTAIL.n472 B 0.015172f
C506 VTAIL.n473 B 0.008153f
C507 VTAIL.n474 B 0.008632f
C508 VTAIL.n475 B 0.01927f
C509 VTAIL.n476 B 0.01927f
C510 VTAIL.n477 B 0.008632f
C511 VTAIL.n478 B 0.008153f
C512 VTAIL.n479 B 0.015172f
C513 VTAIL.n480 B 0.015172f
C514 VTAIL.n481 B 0.008153f
C515 VTAIL.n482 B 0.008632f
C516 VTAIL.n483 B 0.01927f
C517 VTAIL.n484 B 0.040449f
C518 VTAIL.n485 B 0.008632f
C519 VTAIL.n486 B 0.008153f
C520 VTAIL.n487 B 0.034447f
C521 VTAIL.n488 B 0.022483f
C522 VTAIL.n489 B 0.106798f
C523 VTAIL.n490 B 0.020609f
C524 VTAIL.n491 B 0.015172f
C525 VTAIL.n492 B 0.008153f
C526 VTAIL.n493 B 0.01927f
C527 VTAIL.n494 B 0.008632f
C528 VTAIL.n495 B 0.015172f
C529 VTAIL.n496 B 0.008153f
C530 VTAIL.n497 B 0.01927f
C531 VTAIL.n498 B 0.008392f
C532 VTAIL.n499 B 0.015172f
C533 VTAIL.n500 B 0.008392f
C534 VTAIL.n501 B 0.008153f
C535 VTAIL.n502 B 0.01927f
C536 VTAIL.n503 B 0.01927f
C537 VTAIL.n504 B 0.008632f
C538 VTAIL.n505 B 0.015172f
C539 VTAIL.n506 B 0.008153f
C540 VTAIL.n507 B 0.01927f
C541 VTAIL.n508 B 0.008632f
C542 VTAIL.n509 B 0.015172f
C543 VTAIL.n510 B 0.008153f
C544 VTAIL.n511 B 0.01927f
C545 VTAIL.n512 B 0.008632f
C546 VTAIL.n513 B 0.015172f
C547 VTAIL.n514 B 0.008153f
C548 VTAIL.n515 B 0.01927f
C549 VTAIL.n516 B 0.008632f
C550 VTAIL.n517 B 0.015172f
C551 VTAIL.n518 B 0.008153f
C552 VTAIL.n519 B 0.01927f
C553 VTAIL.n520 B 0.008632f
C554 VTAIL.n521 B 1.16023f
C555 VTAIL.n522 B 0.008153f
C556 VTAIL.t5 B 0.031903f
C557 VTAIL.n523 B 0.108425f
C558 VTAIL.n524 B 0.011383f
C559 VTAIL.n525 B 0.014452f
C560 VTAIL.n526 B 0.01927f
C561 VTAIL.n527 B 0.008632f
C562 VTAIL.n528 B 0.008153f
C563 VTAIL.n529 B 0.015172f
C564 VTAIL.n530 B 0.015172f
C565 VTAIL.n531 B 0.008153f
C566 VTAIL.n532 B 0.008632f
C567 VTAIL.n533 B 0.01927f
C568 VTAIL.n534 B 0.01927f
C569 VTAIL.n535 B 0.008632f
C570 VTAIL.n536 B 0.008153f
C571 VTAIL.n537 B 0.015172f
C572 VTAIL.n538 B 0.015172f
C573 VTAIL.n539 B 0.008153f
C574 VTAIL.n540 B 0.008632f
C575 VTAIL.n541 B 0.01927f
C576 VTAIL.n542 B 0.01927f
C577 VTAIL.n543 B 0.008632f
C578 VTAIL.n544 B 0.008153f
C579 VTAIL.n545 B 0.015172f
C580 VTAIL.n546 B 0.015172f
C581 VTAIL.n547 B 0.008153f
C582 VTAIL.n548 B 0.008632f
C583 VTAIL.n549 B 0.01927f
C584 VTAIL.n550 B 0.01927f
C585 VTAIL.n551 B 0.008632f
C586 VTAIL.n552 B 0.008153f
C587 VTAIL.n553 B 0.015172f
C588 VTAIL.n554 B 0.015172f
C589 VTAIL.n555 B 0.008153f
C590 VTAIL.n556 B 0.008632f
C591 VTAIL.n557 B 0.01927f
C592 VTAIL.n558 B 0.01927f
C593 VTAIL.n559 B 0.008632f
C594 VTAIL.n560 B 0.008153f
C595 VTAIL.n561 B 0.015172f
C596 VTAIL.n562 B 0.015172f
C597 VTAIL.n563 B 0.008153f
C598 VTAIL.n564 B 0.008632f
C599 VTAIL.n565 B 0.01927f
C600 VTAIL.n566 B 0.01927f
C601 VTAIL.n567 B 0.008632f
C602 VTAIL.n568 B 0.008153f
C603 VTAIL.n569 B 0.015172f
C604 VTAIL.n570 B 0.015172f
C605 VTAIL.n571 B 0.008153f
C606 VTAIL.n572 B 0.008632f
C607 VTAIL.n573 B 0.01927f
C608 VTAIL.n574 B 0.01927f
C609 VTAIL.n575 B 0.008632f
C610 VTAIL.n576 B 0.008153f
C611 VTAIL.n577 B 0.015172f
C612 VTAIL.n578 B 0.015172f
C613 VTAIL.n579 B 0.008153f
C614 VTAIL.n580 B 0.008632f
C615 VTAIL.n581 B 0.01927f
C616 VTAIL.n582 B 0.040449f
C617 VTAIL.n583 B 0.008632f
C618 VTAIL.n584 B 0.008153f
C619 VTAIL.n585 B 0.034447f
C620 VTAIL.n586 B 0.022483f
C621 VTAIL.n587 B 0.106798f
C622 VTAIL.n588 B 0.020609f
C623 VTAIL.n589 B 0.015172f
C624 VTAIL.n590 B 0.008153f
C625 VTAIL.n591 B 0.01927f
C626 VTAIL.n592 B 0.008632f
C627 VTAIL.n593 B 0.015172f
C628 VTAIL.n594 B 0.008153f
C629 VTAIL.n595 B 0.01927f
C630 VTAIL.n596 B 0.008392f
C631 VTAIL.n597 B 0.015172f
C632 VTAIL.n598 B 0.008392f
C633 VTAIL.n599 B 0.008153f
C634 VTAIL.n600 B 0.01927f
C635 VTAIL.n601 B 0.01927f
C636 VTAIL.n602 B 0.008632f
C637 VTAIL.n603 B 0.015172f
C638 VTAIL.n604 B 0.008153f
C639 VTAIL.n605 B 0.01927f
C640 VTAIL.n606 B 0.008632f
C641 VTAIL.n607 B 0.015172f
C642 VTAIL.n608 B 0.008153f
C643 VTAIL.n609 B 0.01927f
C644 VTAIL.n610 B 0.008632f
C645 VTAIL.n611 B 0.015172f
C646 VTAIL.n612 B 0.008153f
C647 VTAIL.n613 B 0.01927f
C648 VTAIL.n614 B 0.008632f
C649 VTAIL.n615 B 0.015172f
C650 VTAIL.n616 B 0.008153f
C651 VTAIL.n617 B 0.01927f
C652 VTAIL.n618 B 0.008632f
C653 VTAIL.n619 B 1.16023f
C654 VTAIL.n620 B 0.008153f
C655 VTAIL.t6 B 0.031903f
C656 VTAIL.n621 B 0.108425f
C657 VTAIL.n622 B 0.011383f
C658 VTAIL.n623 B 0.014452f
C659 VTAIL.n624 B 0.01927f
C660 VTAIL.n625 B 0.008632f
C661 VTAIL.n626 B 0.008153f
C662 VTAIL.n627 B 0.015172f
C663 VTAIL.n628 B 0.015172f
C664 VTAIL.n629 B 0.008153f
C665 VTAIL.n630 B 0.008632f
C666 VTAIL.n631 B 0.01927f
C667 VTAIL.n632 B 0.01927f
C668 VTAIL.n633 B 0.008632f
C669 VTAIL.n634 B 0.008153f
C670 VTAIL.n635 B 0.015172f
C671 VTAIL.n636 B 0.015172f
C672 VTAIL.n637 B 0.008153f
C673 VTAIL.n638 B 0.008632f
C674 VTAIL.n639 B 0.01927f
C675 VTAIL.n640 B 0.01927f
C676 VTAIL.n641 B 0.008632f
C677 VTAIL.n642 B 0.008153f
C678 VTAIL.n643 B 0.015172f
C679 VTAIL.n644 B 0.015172f
C680 VTAIL.n645 B 0.008153f
C681 VTAIL.n646 B 0.008632f
C682 VTAIL.n647 B 0.01927f
C683 VTAIL.n648 B 0.01927f
C684 VTAIL.n649 B 0.008632f
C685 VTAIL.n650 B 0.008153f
C686 VTAIL.n651 B 0.015172f
C687 VTAIL.n652 B 0.015172f
C688 VTAIL.n653 B 0.008153f
C689 VTAIL.n654 B 0.008632f
C690 VTAIL.n655 B 0.01927f
C691 VTAIL.n656 B 0.01927f
C692 VTAIL.n657 B 0.008632f
C693 VTAIL.n658 B 0.008153f
C694 VTAIL.n659 B 0.015172f
C695 VTAIL.n660 B 0.015172f
C696 VTAIL.n661 B 0.008153f
C697 VTAIL.n662 B 0.008632f
C698 VTAIL.n663 B 0.01927f
C699 VTAIL.n664 B 0.01927f
C700 VTAIL.n665 B 0.008632f
C701 VTAIL.n666 B 0.008153f
C702 VTAIL.n667 B 0.015172f
C703 VTAIL.n668 B 0.015172f
C704 VTAIL.n669 B 0.008153f
C705 VTAIL.n670 B 0.008632f
C706 VTAIL.n671 B 0.01927f
C707 VTAIL.n672 B 0.01927f
C708 VTAIL.n673 B 0.008632f
C709 VTAIL.n674 B 0.008153f
C710 VTAIL.n675 B 0.015172f
C711 VTAIL.n676 B 0.015172f
C712 VTAIL.n677 B 0.008153f
C713 VTAIL.n678 B 0.008632f
C714 VTAIL.n679 B 0.01927f
C715 VTAIL.n680 B 0.040449f
C716 VTAIL.n681 B 0.008632f
C717 VTAIL.n682 B 0.008153f
C718 VTAIL.n683 B 0.034447f
C719 VTAIL.n684 B 0.022483f
C720 VTAIL.n685 B 1.09823f
C721 VTAIL.n686 B 0.020609f
C722 VTAIL.n687 B 0.015172f
C723 VTAIL.n688 B 0.008153f
C724 VTAIL.n689 B 0.01927f
C725 VTAIL.n690 B 0.008632f
C726 VTAIL.n691 B 0.015172f
C727 VTAIL.n692 B 0.008153f
C728 VTAIL.n693 B 0.01927f
C729 VTAIL.n694 B 0.008392f
C730 VTAIL.n695 B 0.015172f
C731 VTAIL.n696 B 0.008632f
C732 VTAIL.n697 B 0.01927f
C733 VTAIL.n698 B 0.008632f
C734 VTAIL.n699 B 0.015172f
C735 VTAIL.n700 B 0.008153f
C736 VTAIL.n701 B 0.01927f
C737 VTAIL.n702 B 0.008632f
C738 VTAIL.n703 B 0.015172f
C739 VTAIL.n704 B 0.008153f
C740 VTAIL.n705 B 0.01927f
C741 VTAIL.n706 B 0.008632f
C742 VTAIL.n707 B 0.015172f
C743 VTAIL.n708 B 0.008153f
C744 VTAIL.n709 B 0.01927f
C745 VTAIL.n710 B 0.008632f
C746 VTAIL.n711 B 0.015172f
C747 VTAIL.n712 B 0.008153f
C748 VTAIL.n713 B 0.01927f
C749 VTAIL.n714 B 0.008632f
C750 VTAIL.n715 B 1.16023f
C751 VTAIL.n716 B 0.008153f
C752 VTAIL.t2 B 0.031903f
C753 VTAIL.n717 B 0.108425f
C754 VTAIL.n718 B 0.011383f
C755 VTAIL.n719 B 0.014452f
C756 VTAIL.n720 B 0.01927f
C757 VTAIL.n721 B 0.008632f
C758 VTAIL.n722 B 0.008153f
C759 VTAIL.n723 B 0.015172f
C760 VTAIL.n724 B 0.015172f
C761 VTAIL.n725 B 0.008153f
C762 VTAIL.n726 B 0.008632f
C763 VTAIL.n727 B 0.01927f
C764 VTAIL.n728 B 0.01927f
C765 VTAIL.n729 B 0.008632f
C766 VTAIL.n730 B 0.008153f
C767 VTAIL.n731 B 0.015172f
C768 VTAIL.n732 B 0.015172f
C769 VTAIL.n733 B 0.008153f
C770 VTAIL.n734 B 0.008632f
C771 VTAIL.n735 B 0.01927f
C772 VTAIL.n736 B 0.01927f
C773 VTAIL.n737 B 0.008632f
C774 VTAIL.n738 B 0.008153f
C775 VTAIL.n739 B 0.015172f
C776 VTAIL.n740 B 0.015172f
C777 VTAIL.n741 B 0.008153f
C778 VTAIL.n742 B 0.008632f
C779 VTAIL.n743 B 0.01927f
C780 VTAIL.n744 B 0.01927f
C781 VTAIL.n745 B 0.008632f
C782 VTAIL.n746 B 0.008153f
C783 VTAIL.n747 B 0.015172f
C784 VTAIL.n748 B 0.015172f
C785 VTAIL.n749 B 0.008153f
C786 VTAIL.n750 B 0.008632f
C787 VTAIL.n751 B 0.01927f
C788 VTAIL.n752 B 0.01927f
C789 VTAIL.n753 B 0.008632f
C790 VTAIL.n754 B 0.008153f
C791 VTAIL.n755 B 0.015172f
C792 VTAIL.n756 B 0.015172f
C793 VTAIL.n757 B 0.008153f
C794 VTAIL.n758 B 0.008153f
C795 VTAIL.n759 B 0.008632f
C796 VTAIL.n760 B 0.01927f
C797 VTAIL.n761 B 0.01927f
C798 VTAIL.n762 B 0.01927f
C799 VTAIL.n763 B 0.008392f
C800 VTAIL.n764 B 0.008153f
C801 VTAIL.n765 B 0.015172f
C802 VTAIL.n766 B 0.015172f
C803 VTAIL.n767 B 0.008153f
C804 VTAIL.n768 B 0.008632f
C805 VTAIL.n769 B 0.01927f
C806 VTAIL.n770 B 0.01927f
C807 VTAIL.n771 B 0.008632f
C808 VTAIL.n772 B 0.008153f
C809 VTAIL.n773 B 0.015172f
C810 VTAIL.n774 B 0.015172f
C811 VTAIL.n775 B 0.008153f
C812 VTAIL.n776 B 0.008632f
C813 VTAIL.n777 B 0.01927f
C814 VTAIL.n778 B 0.040449f
C815 VTAIL.n779 B 0.008632f
C816 VTAIL.n780 B 0.008153f
C817 VTAIL.n781 B 0.034447f
C818 VTAIL.n782 B 0.022483f
C819 VTAIL.n783 B 1.05978f
C820 VDD1.t3 B 0.372355f
C821 VDD1.t1 B 0.372355f
C822 VDD1.n0 B 3.38749f
C823 VDD1.t0 B 0.372355f
C824 VDD1.t2 B 0.372355f
C825 VDD1.n1 B 4.23889f
C826 VP.n0 B 0.036754f
C827 VP.t3 B 2.40332f
C828 VP.n1 B 0.062562f
C829 VP.t2 B 2.51162f
C830 VP.t1 B 2.51095f
C831 VP.n2 B 3.22473f
C832 VP.t0 B 2.40332f
C833 VP.n3 B 0.929149f
C834 VP.n4 B 2.36975f
C835 VP.n5 B 0.036754f
C836 VP.n6 B 0.036754f
C837 VP.n7 B 0.029712f
C838 VP.n8 B 0.062562f
C839 VP.n9 B 0.929149f
C840 VP.n10 B 0.032181f
.ends

