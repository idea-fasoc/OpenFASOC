* NGSPICE file created from diff_pair_sample_0788.ext - technology: sky130A

.subckt diff_pair_sample_0788 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t9 VP.t0 VTAIL.t12 B.t5 sky130_fd_pr__nfet_01v8 ad=2.847 pd=15.38 as=1.2045 ps=7.63 w=7.3 l=0.95
X1 VDD1.t8 VP.t1 VTAIL.t9 B.t8 sky130_fd_pr__nfet_01v8 ad=2.847 pd=15.38 as=1.2045 ps=7.63 w=7.3 l=0.95
X2 VDD2.t9 VN.t0 VTAIL.t8 B.t8 sky130_fd_pr__nfet_01v8 ad=2.847 pd=15.38 as=1.2045 ps=7.63 w=7.3 l=0.95
X3 VDD2.t8 VN.t1 VTAIL.t19 B.t9 sky130_fd_pr__nfet_01v8 ad=1.2045 pd=7.63 as=1.2045 ps=7.63 w=7.3 l=0.95
X4 B.t23 B.t21 B.t22 B.t18 sky130_fd_pr__nfet_01v8 ad=2.847 pd=15.38 as=0 ps=0 w=7.3 l=0.95
X5 VDD1.t7 VP.t2 VTAIL.t15 B.t6 sky130_fd_pr__nfet_01v8 ad=1.2045 pd=7.63 as=2.847 ps=15.38 w=7.3 l=0.95
X6 VTAIL.t14 VP.t3 VDD1.t6 B.t0 sky130_fd_pr__nfet_01v8 ad=1.2045 pd=7.63 as=1.2045 ps=7.63 w=7.3 l=0.95
X7 VTAIL.t10 VP.t4 VDD1.t5 B.t1 sky130_fd_pr__nfet_01v8 ad=1.2045 pd=7.63 as=1.2045 ps=7.63 w=7.3 l=0.95
X8 VDD1.t4 VP.t5 VTAIL.t16 B.t9 sky130_fd_pr__nfet_01v8 ad=1.2045 pd=7.63 as=1.2045 ps=7.63 w=7.3 l=0.95
X9 VDD2.t7 VN.t2 VTAIL.t6 B.t6 sky130_fd_pr__nfet_01v8 ad=1.2045 pd=7.63 as=2.847 ps=15.38 w=7.3 l=0.95
X10 VDD2.t6 VN.t3 VTAIL.t7 B.t7 sky130_fd_pr__nfet_01v8 ad=1.2045 pd=7.63 as=2.847 ps=15.38 w=7.3 l=0.95
X11 VTAIL.t1 VN.t4 VDD2.t5 B.t1 sky130_fd_pr__nfet_01v8 ad=1.2045 pd=7.63 as=1.2045 ps=7.63 w=7.3 l=0.95
X12 B.t20 B.t17 B.t19 B.t18 sky130_fd_pr__nfet_01v8 ad=2.847 pd=15.38 as=0 ps=0 w=7.3 l=0.95
X13 VTAIL.t17 VP.t6 VDD1.t3 B.t4 sky130_fd_pr__nfet_01v8 ad=1.2045 pd=7.63 as=1.2045 ps=7.63 w=7.3 l=0.95
X14 VTAIL.t2 VN.t5 VDD2.t4 B.t2 sky130_fd_pr__nfet_01v8 ad=1.2045 pd=7.63 as=1.2045 ps=7.63 w=7.3 l=0.95
X15 VDD1.t2 VP.t7 VTAIL.t18 B.t3 sky130_fd_pr__nfet_01v8 ad=1.2045 pd=7.63 as=1.2045 ps=7.63 w=7.3 l=0.95
X16 VTAIL.t4 VN.t6 VDD2.t3 B.t4 sky130_fd_pr__nfet_01v8 ad=1.2045 pd=7.63 as=1.2045 ps=7.63 w=7.3 l=0.95
X17 VDD1.t1 VP.t8 VTAIL.t11 B.t7 sky130_fd_pr__nfet_01v8 ad=1.2045 pd=7.63 as=2.847 ps=15.38 w=7.3 l=0.95
X18 B.t16 B.t14 B.t15 B.t11 sky130_fd_pr__nfet_01v8 ad=2.847 pd=15.38 as=0 ps=0 w=7.3 l=0.95
X19 B.t13 B.t10 B.t12 B.t11 sky130_fd_pr__nfet_01v8 ad=2.847 pd=15.38 as=0 ps=0 w=7.3 l=0.95
X20 VTAIL.t13 VP.t9 VDD1.t0 B.t2 sky130_fd_pr__nfet_01v8 ad=1.2045 pd=7.63 as=1.2045 ps=7.63 w=7.3 l=0.95
X21 VDD2.t2 VN.t7 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=1.2045 pd=7.63 as=1.2045 ps=7.63 w=7.3 l=0.95
X22 VDD2.t1 VN.t8 VTAIL.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=2.847 pd=15.38 as=1.2045 ps=7.63 w=7.3 l=0.95
X23 VTAIL.t0 VN.t9 VDD2.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=1.2045 pd=7.63 as=1.2045 ps=7.63 w=7.3 l=0.95
R0 VP.n10 VP.t1 246.935
R1 VP.n5 VP.t0 226.541
R2 VP.n41 VP.t8 226.541
R3 VP.n23 VP.t2 226.541
R4 VP.n34 VP.t5 185.19
R5 VP.n29 VP.t4 185.19
R6 VP.n1 VP.t6 185.19
R7 VP.n16 VP.t7 185.19
R8 VP.n7 VP.t9 185.19
R9 VP.n11 VP.t3 185.19
R10 VP.n42 VP.n41 161.3
R11 VP.n13 VP.n12 161.3
R12 VP.n14 VP.n9 161.3
R13 VP.n16 VP.n15 161.3
R14 VP.n17 VP.n8 161.3
R15 VP.n19 VP.n18 161.3
R16 VP.n21 VP.n20 161.3
R17 VP.n22 VP.n6 161.3
R18 VP.n24 VP.n23 161.3
R19 VP.n40 VP.n0 161.3
R20 VP.n39 VP.n38 161.3
R21 VP.n37 VP.n36 161.3
R22 VP.n35 VP.n2 161.3
R23 VP.n34 VP.n33 161.3
R24 VP.n32 VP.n3 161.3
R25 VP.n31 VP.n30 161.3
R26 VP.n28 VP.n4 161.3
R27 VP.n27 VP.n26 161.3
R28 VP.n25 VP.n5 161.3
R29 VP.n30 VP.n3 54.1398
R30 VP.n36 VP.n35 54.1398
R31 VP.n18 VP.n17 54.1398
R32 VP.n12 VP.n9 54.1398
R33 VP.n28 VP.n27 48.3272
R34 VP.n40 VP.n39 48.3272
R35 VP.n22 VP.n21 48.3272
R36 VP.n13 VP.n10 43.0014
R37 VP.n11 VP.n10 40.664
R38 VP.n25 VP.n24 40.6444
R39 VP.n34 VP.n3 27.0143
R40 VP.n35 VP.n34 27.0143
R41 VP.n17 VP.n16 27.0143
R42 VP.n16 VP.n9 27.0143
R43 VP.n30 VP.n29 13.7719
R44 VP.n36 VP.n1 13.7719
R45 VP.n18 VP.n7 13.7719
R46 VP.n12 VP.n11 13.7719
R47 VP.n27 VP.n5 12.4157
R48 VP.n41 VP.n40 12.4157
R49 VP.n23 VP.n22 12.4157
R50 VP.n29 VP.n28 10.8209
R51 VP.n39 VP.n1 10.8209
R52 VP.n21 VP.n7 10.8209
R53 VP.n14 VP.n13 0.189894
R54 VP.n15 VP.n14 0.189894
R55 VP.n15 VP.n8 0.189894
R56 VP.n19 VP.n8 0.189894
R57 VP.n20 VP.n19 0.189894
R58 VP.n20 VP.n6 0.189894
R59 VP.n24 VP.n6 0.189894
R60 VP.n26 VP.n25 0.189894
R61 VP.n26 VP.n4 0.189894
R62 VP.n31 VP.n4 0.189894
R63 VP.n32 VP.n31 0.189894
R64 VP.n33 VP.n32 0.189894
R65 VP.n33 VP.n2 0.189894
R66 VP.n37 VP.n2 0.189894
R67 VP.n38 VP.n37 0.189894
R68 VP.n38 VP.n0 0.189894
R69 VP.n42 VP.n0 0.189894
R70 VP VP.n42 0.0516364
R71 VTAIL.n152 VTAIL.n122 214.453
R72 VTAIL.n32 VTAIL.n2 214.453
R73 VTAIL.n116 VTAIL.n86 214.453
R74 VTAIL.n76 VTAIL.n46 214.453
R75 VTAIL.n135 VTAIL.n134 185
R76 VTAIL.n137 VTAIL.n136 185
R77 VTAIL.n130 VTAIL.n129 185
R78 VTAIL.n143 VTAIL.n142 185
R79 VTAIL.n145 VTAIL.n144 185
R80 VTAIL.n126 VTAIL.n125 185
R81 VTAIL.n151 VTAIL.n150 185
R82 VTAIL.n153 VTAIL.n152 185
R83 VTAIL.n15 VTAIL.n14 185
R84 VTAIL.n17 VTAIL.n16 185
R85 VTAIL.n10 VTAIL.n9 185
R86 VTAIL.n23 VTAIL.n22 185
R87 VTAIL.n25 VTAIL.n24 185
R88 VTAIL.n6 VTAIL.n5 185
R89 VTAIL.n31 VTAIL.n30 185
R90 VTAIL.n33 VTAIL.n32 185
R91 VTAIL.n117 VTAIL.n116 185
R92 VTAIL.n115 VTAIL.n114 185
R93 VTAIL.n90 VTAIL.n89 185
R94 VTAIL.n109 VTAIL.n108 185
R95 VTAIL.n107 VTAIL.n106 185
R96 VTAIL.n94 VTAIL.n93 185
R97 VTAIL.n101 VTAIL.n100 185
R98 VTAIL.n99 VTAIL.n98 185
R99 VTAIL.n77 VTAIL.n76 185
R100 VTAIL.n75 VTAIL.n74 185
R101 VTAIL.n50 VTAIL.n49 185
R102 VTAIL.n69 VTAIL.n68 185
R103 VTAIL.n67 VTAIL.n66 185
R104 VTAIL.n54 VTAIL.n53 185
R105 VTAIL.n61 VTAIL.n60 185
R106 VTAIL.n59 VTAIL.n58 185
R107 VTAIL.n133 VTAIL.t6 149.524
R108 VTAIL.n13 VTAIL.t11 149.524
R109 VTAIL.n97 VTAIL.t15 149.524
R110 VTAIL.n57 VTAIL.t7 149.524
R111 VTAIL.n136 VTAIL.n135 104.615
R112 VTAIL.n136 VTAIL.n129 104.615
R113 VTAIL.n143 VTAIL.n129 104.615
R114 VTAIL.n144 VTAIL.n143 104.615
R115 VTAIL.n144 VTAIL.n125 104.615
R116 VTAIL.n151 VTAIL.n125 104.615
R117 VTAIL.n152 VTAIL.n151 104.615
R118 VTAIL.n16 VTAIL.n15 104.615
R119 VTAIL.n16 VTAIL.n9 104.615
R120 VTAIL.n23 VTAIL.n9 104.615
R121 VTAIL.n24 VTAIL.n23 104.615
R122 VTAIL.n24 VTAIL.n5 104.615
R123 VTAIL.n31 VTAIL.n5 104.615
R124 VTAIL.n32 VTAIL.n31 104.615
R125 VTAIL.n116 VTAIL.n115 104.615
R126 VTAIL.n115 VTAIL.n89 104.615
R127 VTAIL.n108 VTAIL.n89 104.615
R128 VTAIL.n108 VTAIL.n107 104.615
R129 VTAIL.n107 VTAIL.n93 104.615
R130 VTAIL.n100 VTAIL.n93 104.615
R131 VTAIL.n100 VTAIL.n99 104.615
R132 VTAIL.n76 VTAIL.n75 104.615
R133 VTAIL.n75 VTAIL.n49 104.615
R134 VTAIL.n68 VTAIL.n49 104.615
R135 VTAIL.n68 VTAIL.n67 104.615
R136 VTAIL.n67 VTAIL.n53 104.615
R137 VTAIL.n60 VTAIL.n53 104.615
R138 VTAIL.n60 VTAIL.n59 104.615
R139 VTAIL.n135 VTAIL.t6 52.3082
R140 VTAIL.n15 VTAIL.t11 52.3082
R141 VTAIL.n99 VTAIL.t15 52.3082
R142 VTAIL.n59 VTAIL.t7 52.3082
R143 VTAIL.n85 VTAIL.n84 52.2228
R144 VTAIL.n83 VTAIL.n82 52.2228
R145 VTAIL.n45 VTAIL.n44 52.2228
R146 VTAIL.n43 VTAIL.n42 52.2228
R147 VTAIL.n159 VTAIL.n158 52.2227
R148 VTAIL.n1 VTAIL.n0 52.2227
R149 VTAIL.n39 VTAIL.n38 52.2227
R150 VTAIL.n41 VTAIL.n40 52.2227
R151 VTAIL.n157 VTAIL.n156 36.452
R152 VTAIL.n37 VTAIL.n36 36.452
R153 VTAIL.n121 VTAIL.n120 36.452
R154 VTAIL.n81 VTAIL.n80 36.452
R155 VTAIL.n43 VTAIL.n41 20.8669
R156 VTAIL.n157 VTAIL.n121 19.7634
R157 VTAIL.n154 VTAIL.n153 12.8005
R158 VTAIL.n34 VTAIL.n33 12.8005
R159 VTAIL.n118 VTAIL.n117 12.8005
R160 VTAIL.n78 VTAIL.n77 12.8005
R161 VTAIL.n150 VTAIL.n124 12.0247
R162 VTAIL.n30 VTAIL.n4 12.0247
R163 VTAIL.n114 VTAIL.n88 12.0247
R164 VTAIL.n74 VTAIL.n48 12.0247
R165 VTAIL.n149 VTAIL.n126 11.249
R166 VTAIL.n29 VTAIL.n6 11.249
R167 VTAIL.n113 VTAIL.n90 11.249
R168 VTAIL.n73 VTAIL.n50 11.249
R169 VTAIL.n146 VTAIL.n145 10.4732
R170 VTAIL.n26 VTAIL.n25 10.4732
R171 VTAIL.n110 VTAIL.n109 10.4732
R172 VTAIL.n70 VTAIL.n69 10.4732
R173 VTAIL.n134 VTAIL.n133 10.2747
R174 VTAIL.n14 VTAIL.n13 10.2747
R175 VTAIL.n98 VTAIL.n97 10.2747
R176 VTAIL.n58 VTAIL.n57 10.2747
R177 VTAIL.n142 VTAIL.n128 9.69747
R178 VTAIL.n22 VTAIL.n8 9.69747
R179 VTAIL.n106 VTAIL.n92 9.69747
R180 VTAIL.n66 VTAIL.n52 9.69747
R181 VTAIL.n156 VTAIL.n155 9.45567
R182 VTAIL.n36 VTAIL.n35 9.45567
R183 VTAIL.n120 VTAIL.n119 9.45567
R184 VTAIL.n80 VTAIL.n79 9.45567
R185 VTAIL.n132 VTAIL.n131 9.3005
R186 VTAIL.n139 VTAIL.n138 9.3005
R187 VTAIL.n141 VTAIL.n140 9.3005
R188 VTAIL.n128 VTAIL.n127 9.3005
R189 VTAIL.n147 VTAIL.n146 9.3005
R190 VTAIL.n149 VTAIL.n148 9.3005
R191 VTAIL.n124 VTAIL.n123 9.3005
R192 VTAIL.n155 VTAIL.n154 9.3005
R193 VTAIL.n12 VTAIL.n11 9.3005
R194 VTAIL.n19 VTAIL.n18 9.3005
R195 VTAIL.n21 VTAIL.n20 9.3005
R196 VTAIL.n8 VTAIL.n7 9.3005
R197 VTAIL.n27 VTAIL.n26 9.3005
R198 VTAIL.n29 VTAIL.n28 9.3005
R199 VTAIL.n4 VTAIL.n3 9.3005
R200 VTAIL.n35 VTAIL.n34 9.3005
R201 VTAIL.n96 VTAIL.n95 9.3005
R202 VTAIL.n103 VTAIL.n102 9.3005
R203 VTAIL.n105 VTAIL.n104 9.3005
R204 VTAIL.n92 VTAIL.n91 9.3005
R205 VTAIL.n111 VTAIL.n110 9.3005
R206 VTAIL.n113 VTAIL.n112 9.3005
R207 VTAIL.n88 VTAIL.n87 9.3005
R208 VTAIL.n119 VTAIL.n118 9.3005
R209 VTAIL.n56 VTAIL.n55 9.3005
R210 VTAIL.n63 VTAIL.n62 9.3005
R211 VTAIL.n65 VTAIL.n64 9.3005
R212 VTAIL.n52 VTAIL.n51 9.3005
R213 VTAIL.n71 VTAIL.n70 9.3005
R214 VTAIL.n73 VTAIL.n72 9.3005
R215 VTAIL.n48 VTAIL.n47 9.3005
R216 VTAIL.n79 VTAIL.n78 9.3005
R217 VTAIL.n141 VTAIL.n130 8.92171
R218 VTAIL.n21 VTAIL.n10 8.92171
R219 VTAIL.n105 VTAIL.n94 8.92171
R220 VTAIL.n65 VTAIL.n54 8.92171
R221 VTAIL.n156 VTAIL.n122 8.2187
R222 VTAIL.n36 VTAIL.n2 8.2187
R223 VTAIL.n120 VTAIL.n86 8.2187
R224 VTAIL.n80 VTAIL.n46 8.2187
R225 VTAIL.n138 VTAIL.n137 8.14595
R226 VTAIL.n18 VTAIL.n17 8.14595
R227 VTAIL.n102 VTAIL.n101 8.14595
R228 VTAIL.n62 VTAIL.n61 8.14595
R229 VTAIL.n134 VTAIL.n132 7.3702
R230 VTAIL.n14 VTAIL.n12 7.3702
R231 VTAIL.n98 VTAIL.n96 7.3702
R232 VTAIL.n58 VTAIL.n56 7.3702
R233 VTAIL.n137 VTAIL.n132 5.81868
R234 VTAIL.n17 VTAIL.n12 5.81868
R235 VTAIL.n101 VTAIL.n96 5.81868
R236 VTAIL.n61 VTAIL.n56 5.81868
R237 VTAIL.n154 VTAIL.n122 5.3904
R238 VTAIL.n34 VTAIL.n2 5.3904
R239 VTAIL.n118 VTAIL.n86 5.3904
R240 VTAIL.n78 VTAIL.n46 5.3904
R241 VTAIL.n138 VTAIL.n130 5.04292
R242 VTAIL.n18 VTAIL.n10 5.04292
R243 VTAIL.n102 VTAIL.n94 5.04292
R244 VTAIL.n62 VTAIL.n54 5.04292
R245 VTAIL.n142 VTAIL.n141 4.26717
R246 VTAIL.n22 VTAIL.n21 4.26717
R247 VTAIL.n106 VTAIL.n105 4.26717
R248 VTAIL.n66 VTAIL.n65 4.26717
R249 VTAIL.n145 VTAIL.n128 3.49141
R250 VTAIL.n25 VTAIL.n8 3.49141
R251 VTAIL.n109 VTAIL.n92 3.49141
R252 VTAIL.n69 VTAIL.n52 3.49141
R253 VTAIL.n133 VTAIL.n131 2.84305
R254 VTAIL.n13 VTAIL.n11 2.84305
R255 VTAIL.n97 VTAIL.n95 2.84305
R256 VTAIL.n57 VTAIL.n55 2.84305
R257 VTAIL.n146 VTAIL.n126 2.71565
R258 VTAIL.n26 VTAIL.n6 2.71565
R259 VTAIL.n110 VTAIL.n90 2.71565
R260 VTAIL.n70 VTAIL.n50 2.71565
R261 VTAIL.n158 VTAIL.t3 2.71283
R262 VTAIL.n158 VTAIL.t2 2.71283
R263 VTAIL.n0 VTAIL.t8 2.71283
R264 VTAIL.n0 VTAIL.t0 2.71283
R265 VTAIL.n38 VTAIL.t16 2.71283
R266 VTAIL.n38 VTAIL.t17 2.71283
R267 VTAIL.n40 VTAIL.t12 2.71283
R268 VTAIL.n40 VTAIL.t10 2.71283
R269 VTAIL.n84 VTAIL.t18 2.71283
R270 VTAIL.n84 VTAIL.t13 2.71283
R271 VTAIL.n82 VTAIL.t9 2.71283
R272 VTAIL.n82 VTAIL.t14 2.71283
R273 VTAIL.n44 VTAIL.t19 2.71283
R274 VTAIL.n44 VTAIL.t4 2.71283
R275 VTAIL.n42 VTAIL.t5 2.71283
R276 VTAIL.n42 VTAIL.t1 2.71283
R277 VTAIL.n150 VTAIL.n149 1.93989
R278 VTAIL.n30 VTAIL.n29 1.93989
R279 VTAIL.n114 VTAIL.n113 1.93989
R280 VTAIL.n74 VTAIL.n73 1.93989
R281 VTAIL.n153 VTAIL.n124 1.16414
R282 VTAIL.n33 VTAIL.n4 1.16414
R283 VTAIL.n117 VTAIL.n88 1.16414
R284 VTAIL.n77 VTAIL.n48 1.16414
R285 VTAIL.n45 VTAIL.n43 1.10395
R286 VTAIL.n81 VTAIL.n45 1.10395
R287 VTAIL.n85 VTAIL.n83 1.10395
R288 VTAIL.n121 VTAIL.n85 1.10395
R289 VTAIL.n41 VTAIL.n39 1.10395
R290 VTAIL.n39 VTAIL.n37 1.10395
R291 VTAIL.n159 VTAIL.n157 1.10395
R292 VTAIL.n83 VTAIL.n81 1.02205
R293 VTAIL.n37 VTAIL.n1 1.02205
R294 VTAIL VTAIL.n1 0.886276
R295 VTAIL VTAIL.n159 0.218172
R296 VTAIL.n139 VTAIL.n131 0.155672
R297 VTAIL.n140 VTAIL.n139 0.155672
R298 VTAIL.n140 VTAIL.n127 0.155672
R299 VTAIL.n147 VTAIL.n127 0.155672
R300 VTAIL.n148 VTAIL.n147 0.155672
R301 VTAIL.n148 VTAIL.n123 0.155672
R302 VTAIL.n155 VTAIL.n123 0.155672
R303 VTAIL.n19 VTAIL.n11 0.155672
R304 VTAIL.n20 VTAIL.n19 0.155672
R305 VTAIL.n20 VTAIL.n7 0.155672
R306 VTAIL.n27 VTAIL.n7 0.155672
R307 VTAIL.n28 VTAIL.n27 0.155672
R308 VTAIL.n28 VTAIL.n3 0.155672
R309 VTAIL.n35 VTAIL.n3 0.155672
R310 VTAIL.n119 VTAIL.n87 0.155672
R311 VTAIL.n112 VTAIL.n87 0.155672
R312 VTAIL.n112 VTAIL.n111 0.155672
R313 VTAIL.n111 VTAIL.n91 0.155672
R314 VTAIL.n104 VTAIL.n91 0.155672
R315 VTAIL.n104 VTAIL.n103 0.155672
R316 VTAIL.n103 VTAIL.n95 0.155672
R317 VTAIL.n79 VTAIL.n47 0.155672
R318 VTAIL.n72 VTAIL.n47 0.155672
R319 VTAIL.n72 VTAIL.n71 0.155672
R320 VTAIL.n71 VTAIL.n51 0.155672
R321 VTAIL.n64 VTAIL.n51 0.155672
R322 VTAIL.n64 VTAIL.n63 0.155672
R323 VTAIL.n63 VTAIL.n55 0.155672
R324 VDD1.n30 VDD1.n0 214.453
R325 VDD1.n67 VDD1.n37 214.453
R326 VDD1.n31 VDD1.n30 185
R327 VDD1.n29 VDD1.n28 185
R328 VDD1.n4 VDD1.n3 185
R329 VDD1.n23 VDD1.n22 185
R330 VDD1.n21 VDD1.n20 185
R331 VDD1.n8 VDD1.n7 185
R332 VDD1.n15 VDD1.n14 185
R333 VDD1.n13 VDD1.n12 185
R334 VDD1.n50 VDD1.n49 185
R335 VDD1.n52 VDD1.n51 185
R336 VDD1.n45 VDD1.n44 185
R337 VDD1.n58 VDD1.n57 185
R338 VDD1.n60 VDD1.n59 185
R339 VDD1.n41 VDD1.n40 185
R340 VDD1.n66 VDD1.n65 185
R341 VDD1.n68 VDD1.n67 185
R342 VDD1.n48 VDD1.t9 149.524
R343 VDD1.n11 VDD1.t8 149.524
R344 VDD1.n30 VDD1.n29 104.615
R345 VDD1.n29 VDD1.n3 104.615
R346 VDD1.n22 VDD1.n3 104.615
R347 VDD1.n22 VDD1.n21 104.615
R348 VDD1.n21 VDD1.n7 104.615
R349 VDD1.n14 VDD1.n7 104.615
R350 VDD1.n14 VDD1.n13 104.615
R351 VDD1.n51 VDD1.n50 104.615
R352 VDD1.n51 VDD1.n44 104.615
R353 VDD1.n58 VDD1.n44 104.615
R354 VDD1.n59 VDD1.n58 104.615
R355 VDD1.n59 VDD1.n40 104.615
R356 VDD1.n66 VDD1.n40 104.615
R357 VDD1.n67 VDD1.n66 104.615
R358 VDD1.n75 VDD1.n74 69.6737
R359 VDD1.n36 VDD1.n35 68.9016
R360 VDD1.n77 VDD1.n76 68.9015
R361 VDD1.n73 VDD1.n72 68.9015
R362 VDD1.n36 VDD1.n34 54.2343
R363 VDD1.n73 VDD1.n71 54.2343
R364 VDD1.n13 VDD1.t8 52.3082
R365 VDD1.n50 VDD1.t9 52.3082
R366 VDD1.n77 VDD1.n75 36.3845
R367 VDD1.n32 VDD1.n31 12.8005
R368 VDD1.n69 VDD1.n68 12.8005
R369 VDD1.n28 VDD1.n2 12.0247
R370 VDD1.n65 VDD1.n39 12.0247
R371 VDD1.n27 VDD1.n4 11.249
R372 VDD1.n64 VDD1.n41 11.249
R373 VDD1.n24 VDD1.n23 10.4732
R374 VDD1.n61 VDD1.n60 10.4732
R375 VDD1.n12 VDD1.n11 10.2747
R376 VDD1.n49 VDD1.n48 10.2747
R377 VDD1.n20 VDD1.n6 9.69747
R378 VDD1.n57 VDD1.n43 9.69747
R379 VDD1.n34 VDD1.n33 9.45567
R380 VDD1.n71 VDD1.n70 9.45567
R381 VDD1.n10 VDD1.n9 9.3005
R382 VDD1.n17 VDD1.n16 9.3005
R383 VDD1.n19 VDD1.n18 9.3005
R384 VDD1.n6 VDD1.n5 9.3005
R385 VDD1.n25 VDD1.n24 9.3005
R386 VDD1.n27 VDD1.n26 9.3005
R387 VDD1.n2 VDD1.n1 9.3005
R388 VDD1.n33 VDD1.n32 9.3005
R389 VDD1.n47 VDD1.n46 9.3005
R390 VDD1.n54 VDD1.n53 9.3005
R391 VDD1.n56 VDD1.n55 9.3005
R392 VDD1.n43 VDD1.n42 9.3005
R393 VDD1.n62 VDD1.n61 9.3005
R394 VDD1.n64 VDD1.n63 9.3005
R395 VDD1.n39 VDD1.n38 9.3005
R396 VDD1.n70 VDD1.n69 9.3005
R397 VDD1.n19 VDD1.n8 8.92171
R398 VDD1.n56 VDD1.n45 8.92171
R399 VDD1.n34 VDD1.n0 8.2187
R400 VDD1.n71 VDD1.n37 8.2187
R401 VDD1.n16 VDD1.n15 8.14595
R402 VDD1.n53 VDD1.n52 8.14595
R403 VDD1.n12 VDD1.n10 7.3702
R404 VDD1.n49 VDD1.n47 7.3702
R405 VDD1.n15 VDD1.n10 5.81868
R406 VDD1.n52 VDD1.n47 5.81868
R407 VDD1.n32 VDD1.n0 5.3904
R408 VDD1.n69 VDD1.n37 5.3904
R409 VDD1.n16 VDD1.n8 5.04292
R410 VDD1.n53 VDD1.n45 5.04292
R411 VDD1.n20 VDD1.n19 4.26717
R412 VDD1.n57 VDD1.n56 4.26717
R413 VDD1.n23 VDD1.n6 3.49141
R414 VDD1.n60 VDD1.n43 3.49141
R415 VDD1.n11 VDD1.n9 2.84305
R416 VDD1.n48 VDD1.n46 2.84305
R417 VDD1.n24 VDD1.n4 2.71565
R418 VDD1.n61 VDD1.n41 2.71565
R419 VDD1.n76 VDD1.t0 2.71283
R420 VDD1.n76 VDD1.t7 2.71283
R421 VDD1.n35 VDD1.t6 2.71283
R422 VDD1.n35 VDD1.t2 2.71283
R423 VDD1.n74 VDD1.t3 2.71283
R424 VDD1.n74 VDD1.t1 2.71283
R425 VDD1.n72 VDD1.t5 2.71283
R426 VDD1.n72 VDD1.t4 2.71283
R427 VDD1.n28 VDD1.n27 1.93989
R428 VDD1.n65 VDD1.n64 1.93989
R429 VDD1.n31 VDD1.n2 1.16414
R430 VDD1.n68 VDD1.n39 1.16414
R431 VDD1 VDD1.n77 0.769897
R432 VDD1 VDD1.n36 0.334552
R433 VDD1.n75 VDD1.n73 0.221016
R434 VDD1.n33 VDD1.n1 0.155672
R435 VDD1.n26 VDD1.n1 0.155672
R436 VDD1.n26 VDD1.n25 0.155672
R437 VDD1.n25 VDD1.n5 0.155672
R438 VDD1.n18 VDD1.n5 0.155672
R439 VDD1.n18 VDD1.n17 0.155672
R440 VDD1.n17 VDD1.n9 0.155672
R441 VDD1.n54 VDD1.n46 0.155672
R442 VDD1.n55 VDD1.n54 0.155672
R443 VDD1.n55 VDD1.n42 0.155672
R444 VDD1.n62 VDD1.n42 0.155672
R445 VDD1.n63 VDD1.n62 0.155672
R446 VDD1.n63 VDD1.n38 0.155672
R447 VDD1.n70 VDD1.n38 0.155672
R448 B.n452 B.n95 585
R449 B.n95 B.n58 585
R450 B.n454 B.n453 585
R451 B.n456 B.n94 585
R452 B.n459 B.n458 585
R453 B.n460 B.n93 585
R454 B.n462 B.n461 585
R455 B.n464 B.n92 585
R456 B.n467 B.n466 585
R457 B.n468 B.n91 585
R458 B.n470 B.n469 585
R459 B.n472 B.n90 585
R460 B.n475 B.n474 585
R461 B.n476 B.n89 585
R462 B.n478 B.n477 585
R463 B.n480 B.n88 585
R464 B.n483 B.n482 585
R465 B.n484 B.n87 585
R466 B.n486 B.n485 585
R467 B.n488 B.n86 585
R468 B.n491 B.n490 585
R469 B.n492 B.n85 585
R470 B.n494 B.n493 585
R471 B.n496 B.n84 585
R472 B.n499 B.n498 585
R473 B.n500 B.n83 585
R474 B.n502 B.n501 585
R475 B.n504 B.n82 585
R476 B.n507 B.n506 585
R477 B.n509 B.n79 585
R478 B.n511 B.n510 585
R479 B.n513 B.n78 585
R480 B.n516 B.n515 585
R481 B.n517 B.n77 585
R482 B.n519 B.n518 585
R483 B.n521 B.n76 585
R484 B.n524 B.n523 585
R485 B.n525 B.n73 585
R486 B.n528 B.n527 585
R487 B.n530 B.n72 585
R488 B.n533 B.n532 585
R489 B.n534 B.n71 585
R490 B.n536 B.n535 585
R491 B.n538 B.n70 585
R492 B.n541 B.n540 585
R493 B.n542 B.n69 585
R494 B.n544 B.n543 585
R495 B.n546 B.n68 585
R496 B.n549 B.n548 585
R497 B.n550 B.n67 585
R498 B.n552 B.n551 585
R499 B.n554 B.n66 585
R500 B.n557 B.n556 585
R501 B.n558 B.n65 585
R502 B.n560 B.n559 585
R503 B.n562 B.n64 585
R504 B.n565 B.n564 585
R505 B.n566 B.n63 585
R506 B.n568 B.n567 585
R507 B.n570 B.n62 585
R508 B.n573 B.n572 585
R509 B.n574 B.n61 585
R510 B.n576 B.n575 585
R511 B.n578 B.n60 585
R512 B.n581 B.n580 585
R513 B.n582 B.n59 585
R514 B.n451 B.n57 585
R515 B.n585 B.n57 585
R516 B.n450 B.n56 585
R517 B.n586 B.n56 585
R518 B.n449 B.n55 585
R519 B.n587 B.n55 585
R520 B.n448 B.n447 585
R521 B.n447 B.n51 585
R522 B.n446 B.n50 585
R523 B.n593 B.n50 585
R524 B.n445 B.n49 585
R525 B.n594 B.n49 585
R526 B.n444 B.n48 585
R527 B.n595 B.n48 585
R528 B.n443 B.n442 585
R529 B.n442 B.n44 585
R530 B.n441 B.n43 585
R531 B.n601 B.n43 585
R532 B.n440 B.n42 585
R533 B.n602 B.n42 585
R534 B.n439 B.n41 585
R535 B.n603 B.n41 585
R536 B.n438 B.n437 585
R537 B.n437 B.n40 585
R538 B.n436 B.n36 585
R539 B.n609 B.n36 585
R540 B.n435 B.n35 585
R541 B.n610 B.n35 585
R542 B.n434 B.n34 585
R543 B.n611 B.n34 585
R544 B.n433 B.n432 585
R545 B.n432 B.n33 585
R546 B.n431 B.n29 585
R547 B.n617 B.n29 585
R548 B.n430 B.n28 585
R549 B.n618 B.n28 585
R550 B.n429 B.n27 585
R551 B.n619 B.n27 585
R552 B.n428 B.n427 585
R553 B.n427 B.n26 585
R554 B.n426 B.n22 585
R555 B.n625 B.n22 585
R556 B.n425 B.n21 585
R557 B.n626 B.n21 585
R558 B.n424 B.n20 585
R559 B.n627 B.n20 585
R560 B.n423 B.n422 585
R561 B.n422 B.n19 585
R562 B.n421 B.n15 585
R563 B.n633 B.n15 585
R564 B.n420 B.n14 585
R565 B.n634 B.n14 585
R566 B.n419 B.n13 585
R567 B.n635 B.n13 585
R568 B.n418 B.n417 585
R569 B.n417 B.n12 585
R570 B.n416 B.n415 585
R571 B.n416 B.n8 585
R572 B.n414 B.n7 585
R573 B.n642 B.n7 585
R574 B.n413 B.n6 585
R575 B.n643 B.n6 585
R576 B.n412 B.n5 585
R577 B.n644 B.n5 585
R578 B.n411 B.n410 585
R579 B.n410 B.n4 585
R580 B.n409 B.n96 585
R581 B.n409 B.n408 585
R582 B.n398 B.n97 585
R583 B.n401 B.n97 585
R584 B.n400 B.n399 585
R585 B.n402 B.n400 585
R586 B.n397 B.n102 585
R587 B.n102 B.n101 585
R588 B.n396 B.n395 585
R589 B.n395 B.n394 585
R590 B.n104 B.n103 585
R591 B.n387 B.n104 585
R592 B.n386 B.n385 585
R593 B.n388 B.n386 585
R594 B.n384 B.n109 585
R595 B.n109 B.n108 585
R596 B.n383 B.n382 585
R597 B.n382 B.n381 585
R598 B.n111 B.n110 585
R599 B.n374 B.n111 585
R600 B.n373 B.n372 585
R601 B.n375 B.n373 585
R602 B.n371 B.n116 585
R603 B.n116 B.n115 585
R604 B.n370 B.n369 585
R605 B.n369 B.n368 585
R606 B.n118 B.n117 585
R607 B.n361 B.n118 585
R608 B.n360 B.n359 585
R609 B.n362 B.n360 585
R610 B.n358 B.n123 585
R611 B.n123 B.n122 585
R612 B.n357 B.n356 585
R613 B.n356 B.n355 585
R614 B.n125 B.n124 585
R615 B.n348 B.n125 585
R616 B.n347 B.n346 585
R617 B.n349 B.n347 585
R618 B.n345 B.n130 585
R619 B.n130 B.n129 585
R620 B.n344 B.n343 585
R621 B.n343 B.n342 585
R622 B.n132 B.n131 585
R623 B.n133 B.n132 585
R624 B.n335 B.n334 585
R625 B.n336 B.n335 585
R626 B.n333 B.n138 585
R627 B.n138 B.n137 585
R628 B.n332 B.n331 585
R629 B.n331 B.n330 585
R630 B.n140 B.n139 585
R631 B.n141 B.n140 585
R632 B.n323 B.n322 585
R633 B.n324 B.n323 585
R634 B.n321 B.n146 585
R635 B.n146 B.n145 585
R636 B.n320 B.n319 585
R637 B.n319 B.n318 585
R638 B.n315 B.n150 585
R639 B.n314 B.n313 585
R640 B.n311 B.n151 585
R641 B.n311 B.n149 585
R642 B.n310 B.n309 585
R643 B.n308 B.n307 585
R644 B.n306 B.n153 585
R645 B.n304 B.n303 585
R646 B.n302 B.n154 585
R647 B.n301 B.n300 585
R648 B.n298 B.n155 585
R649 B.n296 B.n295 585
R650 B.n294 B.n156 585
R651 B.n293 B.n292 585
R652 B.n290 B.n157 585
R653 B.n288 B.n287 585
R654 B.n286 B.n158 585
R655 B.n285 B.n284 585
R656 B.n282 B.n159 585
R657 B.n280 B.n279 585
R658 B.n278 B.n160 585
R659 B.n277 B.n276 585
R660 B.n274 B.n161 585
R661 B.n272 B.n271 585
R662 B.n270 B.n162 585
R663 B.n269 B.n268 585
R664 B.n266 B.n163 585
R665 B.n264 B.n263 585
R666 B.n262 B.n164 585
R667 B.n260 B.n259 585
R668 B.n257 B.n167 585
R669 B.n255 B.n254 585
R670 B.n253 B.n168 585
R671 B.n252 B.n251 585
R672 B.n249 B.n169 585
R673 B.n247 B.n246 585
R674 B.n245 B.n170 585
R675 B.n244 B.n243 585
R676 B.n241 B.n240 585
R677 B.n239 B.n238 585
R678 B.n237 B.n175 585
R679 B.n235 B.n234 585
R680 B.n233 B.n176 585
R681 B.n232 B.n231 585
R682 B.n229 B.n177 585
R683 B.n227 B.n226 585
R684 B.n225 B.n178 585
R685 B.n224 B.n223 585
R686 B.n221 B.n179 585
R687 B.n219 B.n218 585
R688 B.n217 B.n180 585
R689 B.n216 B.n215 585
R690 B.n213 B.n181 585
R691 B.n211 B.n210 585
R692 B.n209 B.n182 585
R693 B.n208 B.n207 585
R694 B.n205 B.n183 585
R695 B.n203 B.n202 585
R696 B.n201 B.n184 585
R697 B.n200 B.n199 585
R698 B.n197 B.n185 585
R699 B.n195 B.n194 585
R700 B.n193 B.n186 585
R701 B.n192 B.n191 585
R702 B.n189 B.n187 585
R703 B.n148 B.n147 585
R704 B.n317 B.n316 585
R705 B.n318 B.n317 585
R706 B.n144 B.n143 585
R707 B.n145 B.n144 585
R708 B.n326 B.n325 585
R709 B.n325 B.n324 585
R710 B.n327 B.n142 585
R711 B.n142 B.n141 585
R712 B.n329 B.n328 585
R713 B.n330 B.n329 585
R714 B.n136 B.n135 585
R715 B.n137 B.n136 585
R716 B.n338 B.n337 585
R717 B.n337 B.n336 585
R718 B.n339 B.n134 585
R719 B.n134 B.n133 585
R720 B.n341 B.n340 585
R721 B.n342 B.n341 585
R722 B.n128 B.n127 585
R723 B.n129 B.n128 585
R724 B.n351 B.n350 585
R725 B.n350 B.n349 585
R726 B.n352 B.n126 585
R727 B.n348 B.n126 585
R728 B.n354 B.n353 585
R729 B.n355 B.n354 585
R730 B.n121 B.n120 585
R731 B.n122 B.n121 585
R732 B.n364 B.n363 585
R733 B.n363 B.n362 585
R734 B.n365 B.n119 585
R735 B.n361 B.n119 585
R736 B.n367 B.n366 585
R737 B.n368 B.n367 585
R738 B.n114 B.n113 585
R739 B.n115 B.n114 585
R740 B.n377 B.n376 585
R741 B.n376 B.n375 585
R742 B.n378 B.n112 585
R743 B.n374 B.n112 585
R744 B.n380 B.n379 585
R745 B.n381 B.n380 585
R746 B.n107 B.n106 585
R747 B.n108 B.n107 585
R748 B.n390 B.n389 585
R749 B.n389 B.n388 585
R750 B.n391 B.n105 585
R751 B.n387 B.n105 585
R752 B.n393 B.n392 585
R753 B.n394 B.n393 585
R754 B.n100 B.n99 585
R755 B.n101 B.n100 585
R756 B.n404 B.n403 585
R757 B.n403 B.n402 585
R758 B.n405 B.n98 585
R759 B.n401 B.n98 585
R760 B.n407 B.n406 585
R761 B.n408 B.n407 585
R762 B.n3 B.n0 585
R763 B.n4 B.n3 585
R764 B.n641 B.n1 585
R765 B.n642 B.n641 585
R766 B.n640 B.n639 585
R767 B.n640 B.n8 585
R768 B.n638 B.n9 585
R769 B.n12 B.n9 585
R770 B.n637 B.n636 585
R771 B.n636 B.n635 585
R772 B.n11 B.n10 585
R773 B.n634 B.n11 585
R774 B.n632 B.n631 585
R775 B.n633 B.n632 585
R776 B.n630 B.n16 585
R777 B.n19 B.n16 585
R778 B.n629 B.n628 585
R779 B.n628 B.n627 585
R780 B.n18 B.n17 585
R781 B.n626 B.n18 585
R782 B.n624 B.n623 585
R783 B.n625 B.n624 585
R784 B.n622 B.n23 585
R785 B.n26 B.n23 585
R786 B.n621 B.n620 585
R787 B.n620 B.n619 585
R788 B.n25 B.n24 585
R789 B.n618 B.n25 585
R790 B.n616 B.n615 585
R791 B.n617 B.n616 585
R792 B.n614 B.n30 585
R793 B.n33 B.n30 585
R794 B.n613 B.n612 585
R795 B.n612 B.n611 585
R796 B.n32 B.n31 585
R797 B.n610 B.n32 585
R798 B.n608 B.n607 585
R799 B.n609 B.n608 585
R800 B.n606 B.n37 585
R801 B.n40 B.n37 585
R802 B.n605 B.n604 585
R803 B.n604 B.n603 585
R804 B.n39 B.n38 585
R805 B.n602 B.n39 585
R806 B.n600 B.n599 585
R807 B.n601 B.n600 585
R808 B.n598 B.n45 585
R809 B.n45 B.n44 585
R810 B.n597 B.n596 585
R811 B.n596 B.n595 585
R812 B.n47 B.n46 585
R813 B.n594 B.n47 585
R814 B.n592 B.n591 585
R815 B.n593 B.n592 585
R816 B.n590 B.n52 585
R817 B.n52 B.n51 585
R818 B.n589 B.n588 585
R819 B.n588 B.n587 585
R820 B.n54 B.n53 585
R821 B.n586 B.n54 585
R822 B.n584 B.n583 585
R823 B.n585 B.n584 585
R824 B.n645 B.n644 585
R825 B.n643 B.n2 585
R826 B.n584 B.n59 545.355
R827 B.n95 B.n57 545.355
R828 B.n319 B.n148 545.355
R829 B.n317 B.n150 545.355
R830 B.n74 B.t21 387.764
R831 B.n80 B.t17 387.764
R832 B.n171 B.t10 387.764
R833 B.n165 B.t14 387.764
R834 B.n455 B.n58 256.663
R835 B.n457 B.n58 256.663
R836 B.n463 B.n58 256.663
R837 B.n465 B.n58 256.663
R838 B.n471 B.n58 256.663
R839 B.n473 B.n58 256.663
R840 B.n479 B.n58 256.663
R841 B.n481 B.n58 256.663
R842 B.n487 B.n58 256.663
R843 B.n489 B.n58 256.663
R844 B.n495 B.n58 256.663
R845 B.n497 B.n58 256.663
R846 B.n503 B.n58 256.663
R847 B.n505 B.n58 256.663
R848 B.n512 B.n58 256.663
R849 B.n514 B.n58 256.663
R850 B.n520 B.n58 256.663
R851 B.n522 B.n58 256.663
R852 B.n529 B.n58 256.663
R853 B.n531 B.n58 256.663
R854 B.n537 B.n58 256.663
R855 B.n539 B.n58 256.663
R856 B.n545 B.n58 256.663
R857 B.n547 B.n58 256.663
R858 B.n553 B.n58 256.663
R859 B.n555 B.n58 256.663
R860 B.n561 B.n58 256.663
R861 B.n563 B.n58 256.663
R862 B.n569 B.n58 256.663
R863 B.n571 B.n58 256.663
R864 B.n577 B.n58 256.663
R865 B.n579 B.n58 256.663
R866 B.n312 B.n149 256.663
R867 B.n152 B.n149 256.663
R868 B.n305 B.n149 256.663
R869 B.n299 B.n149 256.663
R870 B.n297 B.n149 256.663
R871 B.n291 B.n149 256.663
R872 B.n289 B.n149 256.663
R873 B.n283 B.n149 256.663
R874 B.n281 B.n149 256.663
R875 B.n275 B.n149 256.663
R876 B.n273 B.n149 256.663
R877 B.n267 B.n149 256.663
R878 B.n265 B.n149 256.663
R879 B.n258 B.n149 256.663
R880 B.n256 B.n149 256.663
R881 B.n250 B.n149 256.663
R882 B.n248 B.n149 256.663
R883 B.n242 B.n149 256.663
R884 B.n174 B.n149 256.663
R885 B.n236 B.n149 256.663
R886 B.n230 B.n149 256.663
R887 B.n228 B.n149 256.663
R888 B.n222 B.n149 256.663
R889 B.n220 B.n149 256.663
R890 B.n214 B.n149 256.663
R891 B.n212 B.n149 256.663
R892 B.n206 B.n149 256.663
R893 B.n204 B.n149 256.663
R894 B.n198 B.n149 256.663
R895 B.n196 B.n149 256.663
R896 B.n190 B.n149 256.663
R897 B.n188 B.n149 256.663
R898 B.n647 B.n646 256.663
R899 B.n80 B.t19 226.023
R900 B.n171 B.t13 226.023
R901 B.n74 B.t22 226.023
R902 B.n165 B.t16 226.023
R903 B.n81 B.t20 201.197
R904 B.n172 B.t12 201.197
R905 B.n75 B.t23 201.197
R906 B.n166 B.t15 201.197
R907 B.n580 B.n578 163.367
R908 B.n576 B.n61 163.367
R909 B.n572 B.n570 163.367
R910 B.n568 B.n63 163.367
R911 B.n564 B.n562 163.367
R912 B.n560 B.n65 163.367
R913 B.n556 B.n554 163.367
R914 B.n552 B.n67 163.367
R915 B.n548 B.n546 163.367
R916 B.n544 B.n69 163.367
R917 B.n540 B.n538 163.367
R918 B.n536 B.n71 163.367
R919 B.n532 B.n530 163.367
R920 B.n528 B.n73 163.367
R921 B.n523 B.n521 163.367
R922 B.n519 B.n77 163.367
R923 B.n515 B.n513 163.367
R924 B.n511 B.n79 163.367
R925 B.n506 B.n504 163.367
R926 B.n502 B.n83 163.367
R927 B.n498 B.n496 163.367
R928 B.n494 B.n85 163.367
R929 B.n490 B.n488 163.367
R930 B.n486 B.n87 163.367
R931 B.n482 B.n480 163.367
R932 B.n478 B.n89 163.367
R933 B.n474 B.n472 163.367
R934 B.n470 B.n91 163.367
R935 B.n466 B.n464 163.367
R936 B.n462 B.n93 163.367
R937 B.n458 B.n456 163.367
R938 B.n454 B.n95 163.367
R939 B.n319 B.n146 163.367
R940 B.n323 B.n146 163.367
R941 B.n323 B.n140 163.367
R942 B.n331 B.n140 163.367
R943 B.n331 B.n138 163.367
R944 B.n335 B.n138 163.367
R945 B.n335 B.n132 163.367
R946 B.n343 B.n132 163.367
R947 B.n343 B.n130 163.367
R948 B.n347 B.n130 163.367
R949 B.n347 B.n125 163.367
R950 B.n356 B.n125 163.367
R951 B.n356 B.n123 163.367
R952 B.n360 B.n123 163.367
R953 B.n360 B.n118 163.367
R954 B.n369 B.n118 163.367
R955 B.n369 B.n116 163.367
R956 B.n373 B.n116 163.367
R957 B.n373 B.n111 163.367
R958 B.n382 B.n111 163.367
R959 B.n382 B.n109 163.367
R960 B.n386 B.n109 163.367
R961 B.n386 B.n104 163.367
R962 B.n395 B.n104 163.367
R963 B.n395 B.n102 163.367
R964 B.n400 B.n102 163.367
R965 B.n400 B.n97 163.367
R966 B.n409 B.n97 163.367
R967 B.n410 B.n409 163.367
R968 B.n410 B.n5 163.367
R969 B.n6 B.n5 163.367
R970 B.n7 B.n6 163.367
R971 B.n416 B.n7 163.367
R972 B.n417 B.n416 163.367
R973 B.n417 B.n13 163.367
R974 B.n14 B.n13 163.367
R975 B.n15 B.n14 163.367
R976 B.n422 B.n15 163.367
R977 B.n422 B.n20 163.367
R978 B.n21 B.n20 163.367
R979 B.n22 B.n21 163.367
R980 B.n427 B.n22 163.367
R981 B.n427 B.n27 163.367
R982 B.n28 B.n27 163.367
R983 B.n29 B.n28 163.367
R984 B.n432 B.n29 163.367
R985 B.n432 B.n34 163.367
R986 B.n35 B.n34 163.367
R987 B.n36 B.n35 163.367
R988 B.n437 B.n36 163.367
R989 B.n437 B.n41 163.367
R990 B.n42 B.n41 163.367
R991 B.n43 B.n42 163.367
R992 B.n442 B.n43 163.367
R993 B.n442 B.n48 163.367
R994 B.n49 B.n48 163.367
R995 B.n50 B.n49 163.367
R996 B.n447 B.n50 163.367
R997 B.n447 B.n55 163.367
R998 B.n56 B.n55 163.367
R999 B.n57 B.n56 163.367
R1000 B.n313 B.n311 163.367
R1001 B.n311 B.n310 163.367
R1002 B.n307 B.n306 163.367
R1003 B.n304 B.n154 163.367
R1004 B.n300 B.n298 163.367
R1005 B.n296 B.n156 163.367
R1006 B.n292 B.n290 163.367
R1007 B.n288 B.n158 163.367
R1008 B.n284 B.n282 163.367
R1009 B.n280 B.n160 163.367
R1010 B.n276 B.n274 163.367
R1011 B.n272 B.n162 163.367
R1012 B.n268 B.n266 163.367
R1013 B.n264 B.n164 163.367
R1014 B.n259 B.n257 163.367
R1015 B.n255 B.n168 163.367
R1016 B.n251 B.n249 163.367
R1017 B.n247 B.n170 163.367
R1018 B.n243 B.n241 163.367
R1019 B.n238 B.n237 163.367
R1020 B.n235 B.n176 163.367
R1021 B.n231 B.n229 163.367
R1022 B.n227 B.n178 163.367
R1023 B.n223 B.n221 163.367
R1024 B.n219 B.n180 163.367
R1025 B.n215 B.n213 163.367
R1026 B.n211 B.n182 163.367
R1027 B.n207 B.n205 163.367
R1028 B.n203 B.n184 163.367
R1029 B.n199 B.n197 163.367
R1030 B.n195 B.n186 163.367
R1031 B.n191 B.n189 163.367
R1032 B.n317 B.n144 163.367
R1033 B.n325 B.n144 163.367
R1034 B.n325 B.n142 163.367
R1035 B.n329 B.n142 163.367
R1036 B.n329 B.n136 163.367
R1037 B.n337 B.n136 163.367
R1038 B.n337 B.n134 163.367
R1039 B.n341 B.n134 163.367
R1040 B.n341 B.n128 163.367
R1041 B.n350 B.n128 163.367
R1042 B.n350 B.n126 163.367
R1043 B.n354 B.n126 163.367
R1044 B.n354 B.n121 163.367
R1045 B.n363 B.n121 163.367
R1046 B.n363 B.n119 163.367
R1047 B.n367 B.n119 163.367
R1048 B.n367 B.n114 163.367
R1049 B.n376 B.n114 163.367
R1050 B.n376 B.n112 163.367
R1051 B.n380 B.n112 163.367
R1052 B.n380 B.n107 163.367
R1053 B.n389 B.n107 163.367
R1054 B.n389 B.n105 163.367
R1055 B.n393 B.n105 163.367
R1056 B.n393 B.n100 163.367
R1057 B.n403 B.n100 163.367
R1058 B.n403 B.n98 163.367
R1059 B.n407 B.n98 163.367
R1060 B.n407 B.n3 163.367
R1061 B.n645 B.n3 163.367
R1062 B.n641 B.n2 163.367
R1063 B.n641 B.n640 163.367
R1064 B.n640 B.n9 163.367
R1065 B.n636 B.n9 163.367
R1066 B.n636 B.n11 163.367
R1067 B.n632 B.n11 163.367
R1068 B.n632 B.n16 163.367
R1069 B.n628 B.n16 163.367
R1070 B.n628 B.n18 163.367
R1071 B.n624 B.n18 163.367
R1072 B.n624 B.n23 163.367
R1073 B.n620 B.n23 163.367
R1074 B.n620 B.n25 163.367
R1075 B.n616 B.n25 163.367
R1076 B.n616 B.n30 163.367
R1077 B.n612 B.n30 163.367
R1078 B.n612 B.n32 163.367
R1079 B.n608 B.n32 163.367
R1080 B.n608 B.n37 163.367
R1081 B.n604 B.n37 163.367
R1082 B.n604 B.n39 163.367
R1083 B.n600 B.n39 163.367
R1084 B.n600 B.n45 163.367
R1085 B.n596 B.n45 163.367
R1086 B.n596 B.n47 163.367
R1087 B.n592 B.n47 163.367
R1088 B.n592 B.n52 163.367
R1089 B.n588 B.n52 163.367
R1090 B.n588 B.n54 163.367
R1091 B.n584 B.n54 163.367
R1092 B.n318 B.n149 119.841
R1093 B.n585 B.n58 119.841
R1094 B.n579 B.n59 71.676
R1095 B.n578 B.n577 71.676
R1096 B.n571 B.n61 71.676
R1097 B.n570 B.n569 71.676
R1098 B.n563 B.n63 71.676
R1099 B.n562 B.n561 71.676
R1100 B.n555 B.n65 71.676
R1101 B.n554 B.n553 71.676
R1102 B.n547 B.n67 71.676
R1103 B.n546 B.n545 71.676
R1104 B.n539 B.n69 71.676
R1105 B.n538 B.n537 71.676
R1106 B.n531 B.n71 71.676
R1107 B.n530 B.n529 71.676
R1108 B.n522 B.n73 71.676
R1109 B.n521 B.n520 71.676
R1110 B.n514 B.n77 71.676
R1111 B.n513 B.n512 71.676
R1112 B.n505 B.n79 71.676
R1113 B.n504 B.n503 71.676
R1114 B.n497 B.n83 71.676
R1115 B.n496 B.n495 71.676
R1116 B.n489 B.n85 71.676
R1117 B.n488 B.n487 71.676
R1118 B.n481 B.n87 71.676
R1119 B.n480 B.n479 71.676
R1120 B.n473 B.n89 71.676
R1121 B.n472 B.n471 71.676
R1122 B.n465 B.n91 71.676
R1123 B.n464 B.n463 71.676
R1124 B.n457 B.n93 71.676
R1125 B.n456 B.n455 71.676
R1126 B.n455 B.n454 71.676
R1127 B.n458 B.n457 71.676
R1128 B.n463 B.n462 71.676
R1129 B.n466 B.n465 71.676
R1130 B.n471 B.n470 71.676
R1131 B.n474 B.n473 71.676
R1132 B.n479 B.n478 71.676
R1133 B.n482 B.n481 71.676
R1134 B.n487 B.n486 71.676
R1135 B.n490 B.n489 71.676
R1136 B.n495 B.n494 71.676
R1137 B.n498 B.n497 71.676
R1138 B.n503 B.n502 71.676
R1139 B.n506 B.n505 71.676
R1140 B.n512 B.n511 71.676
R1141 B.n515 B.n514 71.676
R1142 B.n520 B.n519 71.676
R1143 B.n523 B.n522 71.676
R1144 B.n529 B.n528 71.676
R1145 B.n532 B.n531 71.676
R1146 B.n537 B.n536 71.676
R1147 B.n540 B.n539 71.676
R1148 B.n545 B.n544 71.676
R1149 B.n548 B.n547 71.676
R1150 B.n553 B.n552 71.676
R1151 B.n556 B.n555 71.676
R1152 B.n561 B.n560 71.676
R1153 B.n564 B.n563 71.676
R1154 B.n569 B.n568 71.676
R1155 B.n572 B.n571 71.676
R1156 B.n577 B.n576 71.676
R1157 B.n580 B.n579 71.676
R1158 B.n312 B.n150 71.676
R1159 B.n310 B.n152 71.676
R1160 B.n306 B.n305 71.676
R1161 B.n299 B.n154 71.676
R1162 B.n298 B.n297 71.676
R1163 B.n291 B.n156 71.676
R1164 B.n290 B.n289 71.676
R1165 B.n283 B.n158 71.676
R1166 B.n282 B.n281 71.676
R1167 B.n275 B.n160 71.676
R1168 B.n274 B.n273 71.676
R1169 B.n267 B.n162 71.676
R1170 B.n266 B.n265 71.676
R1171 B.n258 B.n164 71.676
R1172 B.n257 B.n256 71.676
R1173 B.n250 B.n168 71.676
R1174 B.n249 B.n248 71.676
R1175 B.n242 B.n170 71.676
R1176 B.n241 B.n174 71.676
R1177 B.n237 B.n236 71.676
R1178 B.n230 B.n176 71.676
R1179 B.n229 B.n228 71.676
R1180 B.n222 B.n178 71.676
R1181 B.n221 B.n220 71.676
R1182 B.n214 B.n180 71.676
R1183 B.n213 B.n212 71.676
R1184 B.n206 B.n182 71.676
R1185 B.n205 B.n204 71.676
R1186 B.n198 B.n184 71.676
R1187 B.n197 B.n196 71.676
R1188 B.n190 B.n186 71.676
R1189 B.n189 B.n188 71.676
R1190 B.n313 B.n312 71.676
R1191 B.n307 B.n152 71.676
R1192 B.n305 B.n304 71.676
R1193 B.n300 B.n299 71.676
R1194 B.n297 B.n296 71.676
R1195 B.n292 B.n291 71.676
R1196 B.n289 B.n288 71.676
R1197 B.n284 B.n283 71.676
R1198 B.n281 B.n280 71.676
R1199 B.n276 B.n275 71.676
R1200 B.n273 B.n272 71.676
R1201 B.n268 B.n267 71.676
R1202 B.n265 B.n264 71.676
R1203 B.n259 B.n258 71.676
R1204 B.n256 B.n255 71.676
R1205 B.n251 B.n250 71.676
R1206 B.n248 B.n247 71.676
R1207 B.n243 B.n242 71.676
R1208 B.n238 B.n174 71.676
R1209 B.n236 B.n235 71.676
R1210 B.n231 B.n230 71.676
R1211 B.n228 B.n227 71.676
R1212 B.n223 B.n222 71.676
R1213 B.n220 B.n219 71.676
R1214 B.n215 B.n214 71.676
R1215 B.n212 B.n211 71.676
R1216 B.n207 B.n206 71.676
R1217 B.n204 B.n203 71.676
R1218 B.n199 B.n198 71.676
R1219 B.n196 B.n195 71.676
R1220 B.n191 B.n190 71.676
R1221 B.n188 B.n148 71.676
R1222 B.n646 B.n645 71.676
R1223 B.n646 B.n2 71.676
R1224 B.n526 B.n75 59.5399
R1225 B.n508 B.n81 59.5399
R1226 B.n173 B.n172 59.5399
R1227 B.n261 B.n166 59.5399
R1228 B.n318 B.n145 59.4836
R1229 B.n324 B.n145 59.4836
R1230 B.n324 B.n141 59.4836
R1231 B.n330 B.n141 59.4836
R1232 B.n336 B.n137 59.4836
R1233 B.n336 B.n133 59.4836
R1234 B.n342 B.n133 59.4836
R1235 B.n342 B.n129 59.4836
R1236 B.n349 B.n129 59.4836
R1237 B.n349 B.n348 59.4836
R1238 B.n355 B.n122 59.4836
R1239 B.n362 B.n122 59.4836
R1240 B.n362 B.n361 59.4836
R1241 B.n368 B.n115 59.4836
R1242 B.n375 B.n115 59.4836
R1243 B.n375 B.n374 59.4836
R1244 B.n381 B.n108 59.4836
R1245 B.n388 B.n108 59.4836
R1246 B.n388 B.n387 59.4836
R1247 B.n394 B.n101 59.4836
R1248 B.n402 B.n101 59.4836
R1249 B.n402 B.n401 59.4836
R1250 B.n408 B.n4 59.4836
R1251 B.n644 B.n4 59.4836
R1252 B.n644 B.n643 59.4836
R1253 B.n643 B.n642 59.4836
R1254 B.n642 B.n8 59.4836
R1255 B.n635 B.n12 59.4836
R1256 B.n635 B.n634 59.4836
R1257 B.n634 B.n633 59.4836
R1258 B.n627 B.n19 59.4836
R1259 B.n627 B.n626 59.4836
R1260 B.n626 B.n625 59.4836
R1261 B.n619 B.n26 59.4836
R1262 B.n619 B.n618 59.4836
R1263 B.n618 B.n617 59.4836
R1264 B.n611 B.n33 59.4836
R1265 B.n611 B.n610 59.4836
R1266 B.n610 B.n609 59.4836
R1267 B.n603 B.n40 59.4836
R1268 B.n603 B.n602 59.4836
R1269 B.n602 B.n601 59.4836
R1270 B.n601 B.n44 59.4836
R1271 B.n595 B.n44 59.4836
R1272 B.n595 B.n594 59.4836
R1273 B.n593 B.n51 59.4836
R1274 B.n587 B.n51 59.4836
R1275 B.n587 B.n586 59.4836
R1276 B.n586 B.n585 59.4836
R1277 B.n330 B.t11 58.6089
R1278 B.n408 B.t7 58.6089
R1279 B.t8 B.n8 58.6089
R1280 B.t18 B.n593 58.6089
R1281 B.n348 B.t5 56.8593
R1282 B.n40 B.t6 56.8593
R1283 B.n394 B.t4 44.6128
R1284 B.n633 B.t0 44.6128
R1285 B.n361 B.t1 42.8633
R1286 B.n33 B.t2 42.8633
R1287 B.n452 B.n451 35.4346
R1288 B.n316 B.n315 35.4346
R1289 B.n320 B.n147 35.4346
R1290 B.n583 B.n582 35.4346
R1291 B.n381 B.t9 30.6168
R1292 B.n625 B.t3 30.6168
R1293 B.n374 B.t9 28.8673
R1294 B.n26 B.t3 28.8673
R1295 B.n75 B.n74 24.8247
R1296 B.n81 B.n80 24.8247
R1297 B.n172 B.n171 24.8247
R1298 B.n166 B.n165 24.8247
R1299 B B.n647 18.0485
R1300 B.n368 B.t1 16.6208
R1301 B.n617 B.t2 16.6208
R1302 B.n387 B.t4 14.8713
R1303 B.n19 B.t0 14.8713
R1304 B.n316 B.n143 10.6151
R1305 B.n326 B.n143 10.6151
R1306 B.n327 B.n326 10.6151
R1307 B.n328 B.n327 10.6151
R1308 B.n328 B.n135 10.6151
R1309 B.n338 B.n135 10.6151
R1310 B.n339 B.n338 10.6151
R1311 B.n340 B.n339 10.6151
R1312 B.n340 B.n127 10.6151
R1313 B.n351 B.n127 10.6151
R1314 B.n352 B.n351 10.6151
R1315 B.n353 B.n352 10.6151
R1316 B.n353 B.n120 10.6151
R1317 B.n364 B.n120 10.6151
R1318 B.n365 B.n364 10.6151
R1319 B.n366 B.n365 10.6151
R1320 B.n366 B.n113 10.6151
R1321 B.n377 B.n113 10.6151
R1322 B.n378 B.n377 10.6151
R1323 B.n379 B.n378 10.6151
R1324 B.n379 B.n106 10.6151
R1325 B.n390 B.n106 10.6151
R1326 B.n391 B.n390 10.6151
R1327 B.n392 B.n391 10.6151
R1328 B.n392 B.n99 10.6151
R1329 B.n404 B.n99 10.6151
R1330 B.n405 B.n404 10.6151
R1331 B.n406 B.n405 10.6151
R1332 B.n406 B.n0 10.6151
R1333 B.n315 B.n314 10.6151
R1334 B.n314 B.n151 10.6151
R1335 B.n309 B.n151 10.6151
R1336 B.n309 B.n308 10.6151
R1337 B.n308 B.n153 10.6151
R1338 B.n303 B.n153 10.6151
R1339 B.n303 B.n302 10.6151
R1340 B.n302 B.n301 10.6151
R1341 B.n301 B.n155 10.6151
R1342 B.n295 B.n155 10.6151
R1343 B.n295 B.n294 10.6151
R1344 B.n294 B.n293 10.6151
R1345 B.n293 B.n157 10.6151
R1346 B.n287 B.n157 10.6151
R1347 B.n287 B.n286 10.6151
R1348 B.n286 B.n285 10.6151
R1349 B.n285 B.n159 10.6151
R1350 B.n279 B.n159 10.6151
R1351 B.n279 B.n278 10.6151
R1352 B.n278 B.n277 10.6151
R1353 B.n277 B.n161 10.6151
R1354 B.n271 B.n161 10.6151
R1355 B.n271 B.n270 10.6151
R1356 B.n270 B.n269 10.6151
R1357 B.n269 B.n163 10.6151
R1358 B.n263 B.n163 10.6151
R1359 B.n263 B.n262 10.6151
R1360 B.n260 B.n167 10.6151
R1361 B.n254 B.n167 10.6151
R1362 B.n254 B.n253 10.6151
R1363 B.n253 B.n252 10.6151
R1364 B.n252 B.n169 10.6151
R1365 B.n246 B.n169 10.6151
R1366 B.n246 B.n245 10.6151
R1367 B.n245 B.n244 10.6151
R1368 B.n240 B.n239 10.6151
R1369 B.n239 B.n175 10.6151
R1370 B.n234 B.n175 10.6151
R1371 B.n234 B.n233 10.6151
R1372 B.n233 B.n232 10.6151
R1373 B.n232 B.n177 10.6151
R1374 B.n226 B.n177 10.6151
R1375 B.n226 B.n225 10.6151
R1376 B.n225 B.n224 10.6151
R1377 B.n224 B.n179 10.6151
R1378 B.n218 B.n179 10.6151
R1379 B.n218 B.n217 10.6151
R1380 B.n217 B.n216 10.6151
R1381 B.n216 B.n181 10.6151
R1382 B.n210 B.n181 10.6151
R1383 B.n210 B.n209 10.6151
R1384 B.n209 B.n208 10.6151
R1385 B.n208 B.n183 10.6151
R1386 B.n202 B.n183 10.6151
R1387 B.n202 B.n201 10.6151
R1388 B.n201 B.n200 10.6151
R1389 B.n200 B.n185 10.6151
R1390 B.n194 B.n185 10.6151
R1391 B.n194 B.n193 10.6151
R1392 B.n193 B.n192 10.6151
R1393 B.n192 B.n187 10.6151
R1394 B.n187 B.n147 10.6151
R1395 B.n321 B.n320 10.6151
R1396 B.n322 B.n321 10.6151
R1397 B.n322 B.n139 10.6151
R1398 B.n332 B.n139 10.6151
R1399 B.n333 B.n332 10.6151
R1400 B.n334 B.n333 10.6151
R1401 B.n334 B.n131 10.6151
R1402 B.n344 B.n131 10.6151
R1403 B.n345 B.n344 10.6151
R1404 B.n346 B.n345 10.6151
R1405 B.n346 B.n124 10.6151
R1406 B.n357 B.n124 10.6151
R1407 B.n358 B.n357 10.6151
R1408 B.n359 B.n358 10.6151
R1409 B.n359 B.n117 10.6151
R1410 B.n370 B.n117 10.6151
R1411 B.n371 B.n370 10.6151
R1412 B.n372 B.n371 10.6151
R1413 B.n372 B.n110 10.6151
R1414 B.n383 B.n110 10.6151
R1415 B.n384 B.n383 10.6151
R1416 B.n385 B.n384 10.6151
R1417 B.n385 B.n103 10.6151
R1418 B.n396 B.n103 10.6151
R1419 B.n397 B.n396 10.6151
R1420 B.n399 B.n397 10.6151
R1421 B.n399 B.n398 10.6151
R1422 B.n398 B.n96 10.6151
R1423 B.n411 B.n96 10.6151
R1424 B.n412 B.n411 10.6151
R1425 B.n413 B.n412 10.6151
R1426 B.n414 B.n413 10.6151
R1427 B.n415 B.n414 10.6151
R1428 B.n418 B.n415 10.6151
R1429 B.n419 B.n418 10.6151
R1430 B.n420 B.n419 10.6151
R1431 B.n421 B.n420 10.6151
R1432 B.n423 B.n421 10.6151
R1433 B.n424 B.n423 10.6151
R1434 B.n425 B.n424 10.6151
R1435 B.n426 B.n425 10.6151
R1436 B.n428 B.n426 10.6151
R1437 B.n429 B.n428 10.6151
R1438 B.n430 B.n429 10.6151
R1439 B.n431 B.n430 10.6151
R1440 B.n433 B.n431 10.6151
R1441 B.n434 B.n433 10.6151
R1442 B.n435 B.n434 10.6151
R1443 B.n436 B.n435 10.6151
R1444 B.n438 B.n436 10.6151
R1445 B.n439 B.n438 10.6151
R1446 B.n440 B.n439 10.6151
R1447 B.n441 B.n440 10.6151
R1448 B.n443 B.n441 10.6151
R1449 B.n444 B.n443 10.6151
R1450 B.n445 B.n444 10.6151
R1451 B.n446 B.n445 10.6151
R1452 B.n448 B.n446 10.6151
R1453 B.n449 B.n448 10.6151
R1454 B.n450 B.n449 10.6151
R1455 B.n451 B.n450 10.6151
R1456 B.n639 B.n1 10.6151
R1457 B.n639 B.n638 10.6151
R1458 B.n638 B.n637 10.6151
R1459 B.n637 B.n10 10.6151
R1460 B.n631 B.n10 10.6151
R1461 B.n631 B.n630 10.6151
R1462 B.n630 B.n629 10.6151
R1463 B.n629 B.n17 10.6151
R1464 B.n623 B.n17 10.6151
R1465 B.n623 B.n622 10.6151
R1466 B.n622 B.n621 10.6151
R1467 B.n621 B.n24 10.6151
R1468 B.n615 B.n24 10.6151
R1469 B.n615 B.n614 10.6151
R1470 B.n614 B.n613 10.6151
R1471 B.n613 B.n31 10.6151
R1472 B.n607 B.n31 10.6151
R1473 B.n607 B.n606 10.6151
R1474 B.n606 B.n605 10.6151
R1475 B.n605 B.n38 10.6151
R1476 B.n599 B.n38 10.6151
R1477 B.n599 B.n598 10.6151
R1478 B.n598 B.n597 10.6151
R1479 B.n597 B.n46 10.6151
R1480 B.n591 B.n46 10.6151
R1481 B.n591 B.n590 10.6151
R1482 B.n590 B.n589 10.6151
R1483 B.n589 B.n53 10.6151
R1484 B.n583 B.n53 10.6151
R1485 B.n582 B.n581 10.6151
R1486 B.n581 B.n60 10.6151
R1487 B.n575 B.n60 10.6151
R1488 B.n575 B.n574 10.6151
R1489 B.n574 B.n573 10.6151
R1490 B.n573 B.n62 10.6151
R1491 B.n567 B.n62 10.6151
R1492 B.n567 B.n566 10.6151
R1493 B.n566 B.n565 10.6151
R1494 B.n565 B.n64 10.6151
R1495 B.n559 B.n64 10.6151
R1496 B.n559 B.n558 10.6151
R1497 B.n558 B.n557 10.6151
R1498 B.n557 B.n66 10.6151
R1499 B.n551 B.n66 10.6151
R1500 B.n551 B.n550 10.6151
R1501 B.n550 B.n549 10.6151
R1502 B.n549 B.n68 10.6151
R1503 B.n543 B.n68 10.6151
R1504 B.n543 B.n542 10.6151
R1505 B.n542 B.n541 10.6151
R1506 B.n541 B.n70 10.6151
R1507 B.n535 B.n70 10.6151
R1508 B.n535 B.n534 10.6151
R1509 B.n534 B.n533 10.6151
R1510 B.n533 B.n72 10.6151
R1511 B.n527 B.n72 10.6151
R1512 B.n525 B.n524 10.6151
R1513 B.n524 B.n76 10.6151
R1514 B.n518 B.n76 10.6151
R1515 B.n518 B.n517 10.6151
R1516 B.n517 B.n516 10.6151
R1517 B.n516 B.n78 10.6151
R1518 B.n510 B.n78 10.6151
R1519 B.n510 B.n509 10.6151
R1520 B.n507 B.n82 10.6151
R1521 B.n501 B.n82 10.6151
R1522 B.n501 B.n500 10.6151
R1523 B.n500 B.n499 10.6151
R1524 B.n499 B.n84 10.6151
R1525 B.n493 B.n84 10.6151
R1526 B.n493 B.n492 10.6151
R1527 B.n492 B.n491 10.6151
R1528 B.n491 B.n86 10.6151
R1529 B.n485 B.n86 10.6151
R1530 B.n485 B.n484 10.6151
R1531 B.n484 B.n483 10.6151
R1532 B.n483 B.n88 10.6151
R1533 B.n477 B.n88 10.6151
R1534 B.n477 B.n476 10.6151
R1535 B.n476 B.n475 10.6151
R1536 B.n475 B.n90 10.6151
R1537 B.n469 B.n90 10.6151
R1538 B.n469 B.n468 10.6151
R1539 B.n468 B.n467 10.6151
R1540 B.n467 B.n92 10.6151
R1541 B.n461 B.n92 10.6151
R1542 B.n461 B.n460 10.6151
R1543 B.n460 B.n459 10.6151
R1544 B.n459 B.n94 10.6151
R1545 B.n453 B.n94 10.6151
R1546 B.n453 B.n452 10.6151
R1547 B.n647 B.n0 8.11757
R1548 B.n647 B.n1 8.11757
R1549 B.n261 B.n260 6.5566
R1550 B.n244 B.n173 6.5566
R1551 B.n526 B.n525 6.5566
R1552 B.n509 B.n508 6.5566
R1553 B.n262 B.n261 4.05904
R1554 B.n240 B.n173 4.05904
R1555 B.n527 B.n526 4.05904
R1556 B.n508 B.n507 4.05904
R1557 B.n355 B.t5 2.62475
R1558 B.n609 B.t6 2.62475
R1559 B.t11 B.n137 0.875251
R1560 B.n401 B.t7 0.875251
R1561 B.n12 B.t8 0.875251
R1562 B.n594 B.t18 0.875251
R1563 VN.n4 VN.t0 246.935
R1564 VN.n23 VN.t3 246.935
R1565 VN.n17 VN.t2 226.541
R1566 VN.n36 VN.t8 226.541
R1567 VN.n10 VN.t7 185.19
R1568 VN.n5 VN.t9 185.19
R1569 VN.n1 VN.t5 185.19
R1570 VN.n29 VN.t1 185.19
R1571 VN.n24 VN.t6 185.19
R1572 VN.n20 VN.t4 185.19
R1573 VN.n18 VN.n17 161.3
R1574 VN.n37 VN.n36 161.3
R1575 VN.n35 VN.n19 161.3
R1576 VN.n34 VN.n33 161.3
R1577 VN.n32 VN.n31 161.3
R1578 VN.n30 VN.n21 161.3
R1579 VN.n29 VN.n28 161.3
R1580 VN.n27 VN.n22 161.3
R1581 VN.n26 VN.n25 161.3
R1582 VN.n16 VN.n0 161.3
R1583 VN.n15 VN.n14 161.3
R1584 VN.n13 VN.n12 161.3
R1585 VN.n11 VN.n2 161.3
R1586 VN.n10 VN.n9 161.3
R1587 VN.n8 VN.n3 161.3
R1588 VN.n7 VN.n6 161.3
R1589 VN.n6 VN.n3 54.1398
R1590 VN.n12 VN.n11 54.1398
R1591 VN.n25 VN.n22 54.1398
R1592 VN.n31 VN.n30 54.1398
R1593 VN.n16 VN.n15 48.3272
R1594 VN.n35 VN.n34 48.3272
R1595 VN.n26 VN.n23 43.0014
R1596 VN.n7 VN.n4 43.0014
R1597 VN VN.n37 41.0251
R1598 VN.n5 VN.n4 40.664
R1599 VN.n24 VN.n23 40.664
R1600 VN.n10 VN.n3 27.0143
R1601 VN.n11 VN.n10 27.0143
R1602 VN.n29 VN.n22 27.0143
R1603 VN.n30 VN.n29 27.0143
R1604 VN.n6 VN.n5 13.7719
R1605 VN.n12 VN.n1 13.7719
R1606 VN.n25 VN.n24 13.7719
R1607 VN.n31 VN.n20 13.7719
R1608 VN.n17 VN.n16 12.4157
R1609 VN.n36 VN.n35 12.4157
R1610 VN.n15 VN.n1 10.8209
R1611 VN.n34 VN.n20 10.8209
R1612 VN.n37 VN.n19 0.189894
R1613 VN.n33 VN.n19 0.189894
R1614 VN.n33 VN.n32 0.189894
R1615 VN.n32 VN.n21 0.189894
R1616 VN.n28 VN.n21 0.189894
R1617 VN.n28 VN.n27 0.189894
R1618 VN.n27 VN.n26 0.189894
R1619 VN.n8 VN.n7 0.189894
R1620 VN.n9 VN.n8 0.189894
R1621 VN.n9 VN.n2 0.189894
R1622 VN.n13 VN.n2 0.189894
R1623 VN.n14 VN.n13 0.189894
R1624 VN.n14 VN.n0 0.189894
R1625 VN.n18 VN.n0 0.189894
R1626 VN VN.n18 0.0516364
R1627 VDD2.n69 VDD2.n39 214.453
R1628 VDD2.n30 VDD2.n0 214.453
R1629 VDD2.n70 VDD2.n69 185
R1630 VDD2.n68 VDD2.n67 185
R1631 VDD2.n43 VDD2.n42 185
R1632 VDD2.n62 VDD2.n61 185
R1633 VDD2.n60 VDD2.n59 185
R1634 VDD2.n47 VDD2.n46 185
R1635 VDD2.n54 VDD2.n53 185
R1636 VDD2.n52 VDD2.n51 185
R1637 VDD2.n13 VDD2.n12 185
R1638 VDD2.n15 VDD2.n14 185
R1639 VDD2.n8 VDD2.n7 185
R1640 VDD2.n21 VDD2.n20 185
R1641 VDD2.n23 VDD2.n22 185
R1642 VDD2.n4 VDD2.n3 185
R1643 VDD2.n29 VDD2.n28 185
R1644 VDD2.n31 VDD2.n30 185
R1645 VDD2.n11 VDD2.t9 149.524
R1646 VDD2.n50 VDD2.t1 149.524
R1647 VDD2.n69 VDD2.n68 104.615
R1648 VDD2.n68 VDD2.n42 104.615
R1649 VDD2.n61 VDD2.n42 104.615
R1650 VDD2.n61 VDD2.n60 104.615
R1651 VDD2.n60 VDD2.n46 104.615
R1652 VDD2.n53 VDD2.n46 104.615
R1653 VDD2.n53 VDD2.n52 104.615
R1654 VDD2.n14 VDD2.n13 104.615
R1655 VDD2.n14 VDD2.n7 104.615
R1656 VDD2.n21 VDD2.n7 104.615
R1657 VDD2.n22 VDD2.n21 104.615
R1658 VDD2.n22 VDD2.n3 104.615
R1659 VDD2.n29 VDD2.n3 104.615
R1660 VDD2.n30 VDD2.n29 104.615
R1661 VDD2.n38 VDD2.n37 69.6737
R1662 VDD2 VDD2.n77 69.6709
R1663 VDD2.n76 VDD2.n75 68.9016
R1664 VDD2.n36 VDD2.n35 68.9015
R1665 VDD2.n36 VDD2.n34 54.2343
R1666 VDD2.n74 VDD2.n73 53.1308
R1667 VDD2.n52 VDD2.t1 52.3082
R1668 VDD2.n13 VDD2.t9 52.3082
R1669 VDD2.n74 VDD2.n38 35.2498
R1670 VDD2.n71 VDD2.n70 12.8005
R1671 VDD2.n32 VDD2.n31 12.8005
R1672 VDD2.n67 VDD2.n41 12.0247
R1673 VDD2.n28 VDD2.n2 12.0247
R1674 VDD2.n66 VDD2.n43 11.249
R1675 VDD2.n27 VDD2.n4 11.249
R1676 VDD2.n63 VDD2.n62 10.4732
R1677 VDD2.n24 VDD2.n23 10.4732
R1678 VDD2.n51 VDD2.n50 10.2747
R1679 VDD2.n12 VDD2.n11 10.2747
R1680 VDD2.n59 VDD2.n45 9.69747
R1681 VDD2.n20 VDD2.n6 9.69747
R1682 VDD2.n73 VDD2.n72 9.45567
R1683 VDD2.n34 VDD2.n33 9.45567
R1684 VDD2.n49 VDD2.n48 9.3005
R1685 VDD2.n56 VDD2.n55 9.3005
R1686 VDD2.n58 VDD2.n57 9.3005
R1687 VDD2.n45 VDD2.n44 9.3005
R1688 VDD2.n64 VDD2.n63 9.3005
R1689 VDD2.n66 VDD2.n65 9.3005
R1690 VDD2.n41 VDD2.n40 9.3005
R1691 VDD2.n72 VDD2.n71 9.3005
R1692 VDD2.n10 VDD2.n9 9.3005
R1693 VDD2.n17 VDD2.n16 9.3005
R1694 VDD2.n19 VDD2.n18 9.3005
R1695 VDD2.n6 VDD2.n5 9.3005
R1696 VDD2.n25 VDD2.n24 9.3005
R1697 VDD2.n27 VDD2.n26 9.3005
R1698 VDD2.n2 VDD2.n1 9.3005
R1699 VDD2.n33 VDD2.n32 9.3005
R1700 VDD2.n58 VDD2.n47 8.92171
R1701 VDD2.n19 VDD2.n8 8.92171
R1702 VDD2.n73 VDD2.n39 8.2187
R1703 VDD2.n34 VDD2.n0 8.2187
R1704 VDD2.n55 VDD2.n54 8.14595
R1705 VDD2.n16 VDD2.n15 8.14595
R1706 VDD2.n51 VDD2.n49 7.3702
R1707 VDD2.n12 VDD2.n10 7.3702
R1708 VDD2.n54 VDD2.n49 5.81868
R1709 VDD2.n15 VDD2.n10 5.81868
R1710 VDD2.n71 VDD2.n39 5.3904
R1711 VDD2.n32 VDD2.n0 5.3904
R1712 VDD2.n55 VDD2.n47 5.04292
R1713 VDD2.n16 VDD2.n8 5.04292
R1714 VDD2.n59 VDD2.n58 4.26717
R1715 VDD2.n20 VDD2.n19 4.26717
R1716 VDD2.n62 VDD2.n45 3.49141
R1717 VDD2.n23 VDD2.n6 3.49141
R1718 VDD2.n50 VDD2.n48 2.84305
R1719 VDD2.n11 VDD2.n9 2.84305
R1720 VDD2.n63 VDD2.n43 2.71565
R1721 VDD2.n24 VDD2.n4 2.71565
R1722 VDD2.n77 VDD2.t3 2.71283
R1723 VDD2.n77 VDD2.t6 2.71283
R1724 VDD2.n75 VDD2.t5 2.71283
R1725 VDD2.n75 VDD2.t8 2.71283
R1726 VDD2.n37 VDD2.t4 2.71283
R1727 VDD2.n37 VDD2.t7 2.71283
R1728 VDD2.n35 VDD2.t0 2.71283
R1729 VDD2.n35 VDD2.t2 2.71283
R1730 VDD2.n67 VDD2.n66 1.93989
R1731 VDD2.n28 VDD2.n27 1.93989
R1732 VDD2.n70 VDD2.n41 1.16414
R1733 VDD2.n31 VDD2.n2 1.16414
R1734 VDD2.n76 VDD2.n74 1.10395
R1735 VDD2 VDD2.n76 0.334552
R1736 VDD2.n38 VDD2.n36 0.221016
R1737 VDD2.n72 VDD2.n40 0.155672
R1738 VDD2.n65 VDD2.n40 0.155672
R1739 VDD2.n65 VDD2.n64 0.155672
R1740 VDD2.n64 VDD2.n44 0.155672
R1741 VDD2.n57 VDD2.n44 0.155672
R1742 VDD2.n57 VDD2.n56 0.155672
R1743 VDD2.n56 VDD2.n48 0.155672
R1744 VDD2.n17 VDD2.n9 0.155672
R1745 VDD2.n18 VDD2.n17 0.155672
R1746 VDD2.n18 VDD2.n5 0.155672
R1747 VDD2.n25 VDD2.n5 0.155672
R1748 VDD2.n26 VDD2.n25 0.155672
R1749 VDD2.n26 VDD2.n1 0.155672
R1750 VDD2.n33 VDD2.n1 0.155672
C0 VP VDD1 5.12026f
C1 VDD2 VTAIL 8.776549f
C2 VP VDD2 0.372968f
C3 VN VTAIL 5.03852f
C4 VP VN 5.08837f
C5 VDD2 VDD1 1.12799f
C6 VN VDD1 0.14984f
C7 VP VTAIL 5.05289f
C8 VN VDD2 4.90011f
C9 VDD1 VTAIL 8.737519f
C10 VDD2 B 4.41893f
C11 VDD1 B 4.36859f
C12 VTAIL B 5.02956f
C13 VN B 10.017962f
C14 VP B 8.372352f
C15 VDD2.n0 B 0.033246f
C16 VDD2.n1 B 0.02358f
C17 VDD2.n2 B 0.012671f
C18 VDD2.n3 B 0.02995f
C19 VDD2.n4 B 0.013416f
C20 VDD2.n5 B 0.02358f
C21 VDD2.n6 B 0.012671f
C22 VDD2.n7 B 0.02995f
C23 VDD2.n8 B 0.013416f
C24 VDD2.n9 B 0.696542f
C25 VDD2.n10 B 0.012671f
C26 VDD2.t9 B 0.050024f
C27 VDD2.n11 B 0.127529f
C28 VDD2.n12 B 0.021172f
C29 VDD2.n13 B 0.022462f
C30 VDD2.n14 B 0.02995f
C31 VDD2.n15 B 0.013416f
C32 VDD2.n16 B 0.012671f
C33 VDD2.n17 B 0.02358f
C34 VDD2.n18 B 0.02358f
C35 VDD2.n19 B 0.012671f
C36 VDD2.n20 B 0.013416f
C37 VDD2.n21 B 0.02995f
C38 VDD2.n22 B 0.02995f
C39 VDD2.n23 B 0.013416f
C40 VDD2.n24 B 0.012671f
C41 VDD2.n25 B 0.02358f
C42 VDD2.n26 B 0.02358f
C43 VDD2.n27 B 0.012671f
C44 VDD2.n28 B 0.013416f
C45 VDD2.n29 B 0.02995f
C46 VDD2.n30 B 0.062293f
C47 VDD2.n31 B 0.013416f
C48 VDD2.n32 B 0.024776f
C49 VDD2.n33 B 0.061592f
C50 VDD2.n34 B 0.084628f
C51 VDD2.t0 B 0.136028f
C52 VDD2.t2 B 0.136028f
C53 VDD2.n35 B 1.16964f
C54 VDD2.n36 B 0.418365f
C55 VDD2.t4 B 0.136028f
C56 VDD2.t7 B 0.136028f
C57 VDD2.n37 B 1.17338f
C58 VDD2.n38 B 1.64599f
C59 VDD2.n39 B 0.033246f
C60 VDD2.n40 B 0.02358f
C61 VDD2.n41 B 0.012671f
C62 VDD2.n42 B 0.02995f
C63 VDD2.n43 B 0.013416f
C64 VDD2.n44 B 0.02358f
C65 VDD2.n45 B 0.012671f
C66 VDD2.n46 B 0.02995f
C67 VDD2.n47 B 0.013416f
C68 VDD2.n48 B 0.696542f
C69 VDD2.n49 B 0.012671f
C70 VDD2.t1 B 0.050024f
C71 VDD2.n50 B 0.127529f
C72 VDD2.n51 B 0.021172f
C73 VDD2.n52 B 0.022462f
C74 VDD2.n53 B 0.02995f
C75 VDD2.n54 B 0.013416f
C76 VDD2.n55 B 0.012671f
C77 VDD2.n56 B 0.02358f
C78 VDD2.n57 B 0.02358f
C79 VDD2.n58 B 0.012671f
C80 VDD2.n59 B 0.013416f
C81 VDD2.n60 B 0.02995f
C82 VDD2.n61 B 0.02995f
C83 VDD2.n62 B 0.013416f
C84 VDD2.n63 B 0.012671f
C85 VDD2.n64 B 0.02358f
C86 VDD2.n65 B 0.02358f
C87 VDD2.n66 B 0.012671f
C88 VDD2.n67 B 0.013416f
C89 VDD2.n68 B 0.02995f
C90 VDD2.n69 B 0.062293f
C91 VDD2.n70 B 0.013416f
C92 VDD2.n71 B 0.024776f
C93 VDD2.n72 B 0.061592f
C94 VDD2.n73 B 0.081916f
C95 VDD2.n74 B 1.77748f
C96 VDD2.t5 B 0.136028f
C97 VDD2.t8 B 0.136028f
C98 VDD2.n75 B 1.16964f
C99 VDD2.n76 B 0.293912f
C100 VDD2.t3 B 0.136028f
C101 VDD2.t6 B 0.136028f
C102 VDD2.n77 B 1.17335f
C103 VN.n0 B 0.038469f
C104 VN.t5 B 0.713509f
C105 VN.n1 B 0.284433f
C106 VN.n2 B 0.038469f
C107 VN.t7 B 0.713509f
C108 VN.n3 B 0.041891f
C109 VN.t0 B 0.797228f
C110 VN.n4 B 0.33061f
C111 VN.t9 B 0.713509f
C112 VN.n5 B 0.323771f
C113 VN.n6 B 0.051613f
C114 VN.n7 B 0.166547f
C115 VN.n8 B 0.038469f
C116 VN.n9 B 0.038469f
C117 VN.n10 B 0.326236f
C118 VN.n11 B 0.041891f
C119 VN.n12 B 0.051613f
C120 VN.n13 B 0.038469f
C121 VN.n14 B 0.038469f
C122 VN.n15 B 0.051961f
C123 VN.n16 B 0.014899f
C124 VN.t2 B 0.769155f
C125 VN.n17 B 0.330313f
C126 VN.n18 B 0.029812f
C127 VN.n19 B 0.038469f
C128 VN.t4 B 0.713509f
C129 VN.n20 B 0.284433f
C130 VN.n21 B 0.038469f
C131 VN.t1 B 0.713509f
C132 VN.n22 B 0.041891f
C133 VN.t3 B 0.797228f
C134 VN.n23 B 0.33061f
C135 VN.t6 B 0.713509f
C136 VN.n24 B 0.323771f
C137 VN.n25 B 0.051613f
C138 VN.n26 B 0.166547f
C139 VN.n27 B 0.038469f
C140 VN.n28 B 0.038469f
C141 VN.n29 B 0.326236f
C142 VN.n30 B 0.041891f
C143 VN.n31 B 0.051613f
C144 VN.n32 B 0.038469f
C145 VN.n33 B 0.038469f
C146 VN.n34 B 0.051961f
C147 VN.n35 B 0.014899f
C148 VN.t8 B 0.769155f
C149 VN.n36 B 0.330313f
C150 VN.n37 B 1.52771f
C151 VDD1.n0 B 0.033277f
C152 VDD1.n1 B 0.023603f
C153 VDD1.n2 B 0.012683f
C154 VDD1.n3 B 0.029978f
C155 VDD1.n4 B 0.013429f
C156 VDD1.n5 B 0.023603f
C157 VDD1.n6 B 0.012683f
C158 VDD1.n7 B 0.029978f
C159 VDD1.n8 B 0.013429f
C160 VDD1.n9 B 0.697194f
C161 VDD1.n10 B 0.012683f
C162 VDD1.t8 B 0.050071f
C163 VDD1.n11 B 0.127649f
C164 VDD1.n12 B 0.021192f
C165 VDD1.n13 B 0.022483f
C166 VDD1.n14 B 0.029978f
C167 VDD1.n15 B 0.013429f
C168 VDD1.n16 B 0.012683f
C169 VDD1.n17 B 0.023603f
C170 VDD1.n18 B 0.023603f
C171 VDD1.n19 B 0.012683f
C172 VDD1.n20 B 0.013429f
C173 VDD1.n21 B 0.029978f
C174 VDD1.n22 B 0.029978f
C175 VDD1.n23 B 0.013429f
C176 VDD1.n24 B 0.012683f
C177 VDD1.n25 B 0.023603f
C178 VDD1.n26 B 0.023603f
C179 VDD1.n27 B 0.012683f
C180 VDD1.n28 B 0.013429f
C181 VDD1.n29 B 0.029978f
C182 VDD1.n30 B 0.062351f
C183 VDD1.n31 B 0.013429f
C184 VDD1.n32 B 0.024799f
C185 VDD1.n33 B 0.06165f
C186 VDD1.n34 B 0.084707f
C187 VDD1.t6 B 0.136155f
C188 VDD1.t2 B 0.136155f
C189 VDD1.n35 B 1.17074f
C190 VDD1.n36 B 0.424904f
C191 VDD1.n37 B 0.033277f
C192 VDD1.n38 B 0.023603f
C193 VDD1.n39 B 0.012683f
C194 VDD1.n40 B 0.029978f
C195 VDD1.n41 B 0.013429f
C196 VDD1.n42 B 0.023603f
C197 VDD1.n43 B 0.012683f
C198 VDD1.n44 B 0.029978f
C199 VDD1.n45 B 0.013429f
C200 VDD1.n46 B 0.697194f
C201 VDD1.n47 B 0.012683f
C202 VDD1.t9 B 0.050071f
C203 VDD1.n48 B 0.127649f
C204 VDD1.n49 B 0.021192f
C205 VDD1.n50 B 0.022483f
C206 VDD1.n51 B 0.029978f
C207 VDD1.n52 B 0.013429f
C208 VDD1.n53 B 0.012683f
C209 VDD1.n54 B 0.023603f
C210 VDD1.n55 B 0.023603f
C211 VDD1.n56 B 0.012683f
C212 VDD1.n57 B 0.013429f
C213 VDD1.n58 B 0.029978f
C214 VDD1.n59 B 0.029978f
C215 VDD1.n60 B 0.013429f
C216 VDD1.n61 B 0.012683f
C217 VDD1.n62 B 0.023603f
C218 VDD1.n63 B 0.023603f
C219 VDD1.n64 B 0.012683f
C220 VDD1.n65 B 0.013429f
C221 VDD1.n66 B 0.029978f
C222 VDD1.n67 B 0.062351f
C223 VDD1.n68 B 0.013429f
C224 VDD1.n69 B 0.024799f
C225 VDD1.n70 B 0.06165f
C226 VDD1.n71 B 0.084707f
C227 VDD1.t5 B 0.136155f
C228 VDD1.t4 B 0.136155f
C229 VDD1.n72 B 1.17073f
C230 VDD1.n73 B 0.418756f
C231 VDD1.t3 B 0.136155f
C232 VDD1.t1 B 0.136155f
C233 VDD1.n74 B 1.17447f
C234 VDD1.n75 B 1.72379f
C235 VDD1.t0 B 0.136155f
C236 VDD1.t7 B 0.136155f
C237 VDD1.n76 B 1.17073f
C238 VDD1.n77 B 1.99344f
C239 VTAIL.t8 B 0.15092f
C240 VTAIL.t0 B 0.15092f
C241 VTAIL.n0 B 1.23383f
C242 VTAIL.n1 B 0.393996f
C243 VTAIL.n2 B 0.036885f
C244 VTAIL.n3 B 0.026162f
C245 VTAIL.n4 B 0.014058f
C246 VTAIL.n5 B 0.033229f
C247 VTAIL.n6 B 0.014885f
C248 VTAIL.n7 B 0.026162f
C249 VTAIL.n8 B 0.014058f
C250 VTAIL.n9 B 0.033229f
C251 VTAIL.n10 B 0.014885f
C252 VTAIL.n11 B 0.772796f
C253 VTAIL.n12 B 0.014058f
C254 VTAIL.t11 B 0.0555f
C255 VTAIL.n13 B 0.14149f
C256 VTAIL.n14 B 0.02349f
C257 VTAIL.n15 B 0.024921f
C258 VTAIL.n16 B 0.033229f
C259 VTAIL.n17 B 0.014885f
C260 VTAIL.n18 B 0.014058f
C261 VTAIL.n19 B 0.026162f
C262 VTAIL.n20 B 0.026162f
C263 VTAIL.n21 B 0.014058f
C264 VTAIL.n22 B 0.014885f
C265 VTAIL.n23 B 0.033229f
C266 VTAIL.n24 B 0.033229f
C267 VTAIL.n25 B 0.014885f
C268 VTAIL.n26 B 0.014058f
C269 VTAIL.n27 B 0.026162f
C270 VTAIL.n28 B 0.026162f
C271 VTAIL.n29 B 0.014058f
C272 VTAIL.n30 B 0.014885f
C273 VTAIL.n31 B 0.033229f
C274 VTAIL.n32 B 0.069113f
C275 VTAIL.n33 B 0.014885f
C276 VTAIL.n34 B 0.027489f
C277 VTAIL.n35 B 0.068335f
C278 VTAIL.n36 B 0.072873f
C279 VTAIL.n37 B 0.205932f
C280 VTAIL.t16 B 0.15092f
C281 VTAIL.t17 B 0.15092f
C282 VTAIL.n38 B 1.23383f
C283 VTAIL.n39 B 0.419249f
C284 VTAIL.t12 B 0.15092f
C285 VTAIL.t10 B 0.15092f
C286 VTAIL.n40 B 1.23383f
C287 VTAIL.n41 B 1.39815f
C288 VTAIL.t5 B 0.15092f
C289 VTAIL.t1 B 0.15092f
C290 VTAIL.n42 B 1.23384f
C291 VTAIL.n43 B 1.39815f
C292 VTAIL.t19 B 0.15092f
C293 VTAIL.t4 B 0.15092f
C294 VTAIL.n44 B 1.23384f
C295 VTAIL.n45 B 0.419241f
C296 VTAIL.n46 B 0.036885f
C297 VTAIL.n47 B 0.026162f
C298 VTAIL.n48 B 0.014058f
C299 VTAIL.n49 B 0.033229f
C300 VTAIL.n50 B 0.014885f
C301 VTAIL.n51 B 0.026162f
C302 VTAIL.n52 B 0.014058f
C303 VTAIL.n53 B 0.033229f
C304 VTAIL.n54 B 0.014885f
C305 VTAIL.n55 B 0.772796f
C306 VTAIL.n56 B 0.014058f
C307 VTAIL.t7 B 0.0555f
C308 VTAIL.n57 B 0.14149f
C309 VTAIL.n58 B 0.02349f
C310 VTAIL.n59 B 0.024921f
C311 VTAIL.n60 B 0.033229f
C312 VTAIL.n61 B 0.014885f
C313 VTAIL.n62 B 0.014058f
C314 VTAIL.n63 B 0.026162f
C315 VTAIL.n64 B 0.026162f
C316 VTAIL.n65 B 0.014058f
C317 VTAIL.n66 B 0.014885f
C318 VTAIL.n67 B 0.033229f
C319 VTAIL.n68 B 0.033229f
C320 VTAIL.n69 B 0.014885f
C321 VTAIL.n70 B 0.014058f
C322 VTAIL.n71 B 0.026162f
C323 VTAIL.n72 B 0.026162f
C324 VTAIL.n73 B 0.014058f
C325 VTAIL.n74 B 0.014885f
C326 VTAIL.n75 B 0.033229f
C327 VTAIL.n76 B 0.069113f
C328 VTAIL.n77 B 0.014885f
C329 VTAIL.n78 B 0.027489f
C330 VTAIL.n79 B 0.068335f
C331 VTAIL.n80 B 0.072873f
C332 VTAIL.n81 B 0.205932f
C333 VTAIL.t9 B 0.15092f
C334 VTAIL.t14 B 0.15092f
C335 VTAIL.n82 B 1.23384f
C336 VTAIL.n83 B 0.412337f
C337 VTAIL.t18 B 0.15092f
C338 VTAIL.t13 B 0.15092f
C339 VTAIL.n84 B 1.23384f
C340 VTAIL.n85 B 0.419241f
C341 VTAIL.n86 B 0.036885f
C342 VTAIL.n87 B 0.026162f
C343 VTAIL.n88 B 0.014058f
C344 VTAIL.n89 B 0.033229f
C345 VTAIL.n90 B 0.014885f
C346 VTAIL.n91 B 0.026162f
C347 VTAIL.n92 B 0.014058f
C348 VTAIL.n93 B 0.033229f
C349 VTAIL.n94 B 0.014885f
C350 VTAIL.n95 B 0.772796f
C351 VTAIL.n96 B 0.014058f
C352 VTAIL.t15 B 0.0555f
C353 VTAIL.n97 B 0.14149f
C354 VTAIL.n98 B 0.02349f
C355 VTAIL.n99 B 0.024921f
C356 VTAIL.n100 B 0.033229f
C357 VTAIL.n101 B 0.014885f
C358 VTAIL.n102 B 0.014058f
C359 VTAIL.n103 B 0.026162f
C360 VTAIL.n104 B 0.026162f
C361 VTAIL.n105 B 0.014058f
C362 VTAIL.n106 B 0.014885f
C363 VTAIL.n107 B 0.033229f
C364 VTAIL.n108 B 0.033229f
C365 VTAIL.n109 B 0.014885f
C366 VTAIL.n110 B 0.014058f
C367 VTAIL.n111 B 0.026162f
C368 VTAIL.n112 B 0.026162f
C369 VTAIL.n113 B 0.014058f
C370 VTAIL.n114 B 0.014885f
C371 VTAIL.n115 B 0.033229f
C372 VTAIL.n116 B 0.069113f
C373 VTAIL.n117 B 0.014885f
C374 VTAIL.n118 B 0.027489f
C375 VTAIL.n119 B 0.068335f
C376 VTAIL.n120 B 0.072873f
C377 VTAIL.n121 B 1.09872f
C378 VTAIL.n122 B 0.036885f
C379 VTAIL.n123 B 0.026162f
C380 VTAIL.n124 B 0.014058f
C381 VTAIL.n125 B 0.033229f
C382 VTAIL.n126 B 0.014885f
C383 VTAIL.n127 B 0.026162f
C384 VTAIL.n128 B 0.014058f
C385 VTAIL.n129 B 0.033229f
C386 VTAIL.n130 B 0.014885f
C387 VTAIL.n131 B 0.772796f
C388 VTAIL.n132 B 0.014058f
C389 VTAIL.t6 B 0.0555f
C390 VTAIL.n133 B 0.14149f
C391 VTAIL.n134 B 0.02349f
C392 VTAIL.n135 B 0.024921f
C393 VTAIL.n136 B 0.033229f
C394 VTAIL.n137 B 0.014885f
C395 VTAIL.n138 B 0.014058f
C396 VTAIL.n139 B 0.026162f
C397 VTAIL.n140 B 0.026162f
C398 VTAIL.n141 B 0.014058f
C399 VTAIL.n142 B 0.014885f
C400 VTAIL.n143 B 0.033229f
C401 VTAIL.n144 B 0.033229f
C402 VTAIL.n145 B 0.014885f
C403 VTAIL.n146 B 0.014058f
C404 VTAIL.n147 B 0.026162f
C405 VTAIL.n148 B 0.026162f
C406 VTAIL.n149 B 0.014058f
C407 VTAIL.n150 B 0.014885f
C408 VTAIL.n151 B 0.033229f
C409 VTAIL.n152 B 0.069113f
C410 VTAIL.n153 B 0.014885f
C411 VTAIL.n154 B 0.027489f
C412 VTAIL.n155 B 0.068335f
C413 VTAIL.n156 B 0.072873f
C414 VTAIL.n157 B 1.09872f
C415 VTAIL.t3 B 0.15092f
C416 VTAIL.t2 B 0.15092f
C417 VTAIL.n158 B 1.23383f
C418 VTAIL.n159 B 0.344579f
C419 VP.n0 B 0.03938f
C420 VP.t6 B 0.730412f
C421 VP.n1 B 0.291172f
C422 VP.n2 B 0.03938f
C423 VP.t5 B 0.730412f
C424 VP.n3 B 0.042883f
C425 VP.n4 B 0.03938f
C426 VP.t4 B 0.730412f
C427 VP.t0 B 0.787377f
C428 VP.n5 B 0.338138f
C429 VP.n6 B 0.03938f
C430 VP.t2 B 0.787377f
C431 VP.t9 B 0.730412f
C432 VP.n7 B 0.291172f
C433 VP.n8 B 0.03938f
C434 VP.t7 B 0.730412f
C435 VP.n9 B 0.042883f
C436 VP.t1 B 0.816115f
C437 VP.n10 B 0.338443f
C438 VP.t3 B 0.730412f
C439 VP.n11 B 0.331441f
C440 VP.n12 B 0.052836f
C441 VP.n13 B 0.170493f
C442 VP.n14 B 0.03938f
C443 VP.n15 B 0.03938f
C444 VP.n16 B 0.333965f
C445 VP.n17 B 0.042883f
C446 VP.n18 B 0.052836f
C447 VP.n19 B 0.03938f
C448 VP.n20 B 0.03938f
C449 VP.n21 B 0.053192f
C450 VP.n22 B 0.015252f
C451 VP.n23 B 0.338138f
C452 VP.n24 B 1.53799f
C453 VP.n25 B 1.57292f
C454 VP.n26 B 0.03938f
C455 VP.n27 B 0.015252f
C456 VP.n28 B 0.053192f
C457 VP.n29 B 0.291172f
C458 VP.n30 B 0.052836f
C459 VP.n31 B 0.03938f
C460 VP.n32 B 0.03938f
C461 VP.n33 B 0.03938f
C462 VP.n34 B 0.333965f
C463 VP.n35 B 0.042883f
C464 VP.n36 B 0.052836f
C465 VP.n37 B 0.03938f
C466 VP.n38 B 0.03938f
C467 VP.n39 B 0.053192f
C468 VP.n40 B 0.015252f
C469 VP.t8 B 0.787377f
C470 VP.n41 B 0.338138f
C471 VP.n42 B 0.030518f
.ends

