* NGSPICE file created from diff_pair_sample_1325.ext - technology: sky130A

.subckt diff_pair_sample_1325 VTAIL VN VP B VDD2 VDD1
X0 B.t15 B.t13 B.t14 B.t7 sky130_fd_pr__nfet_01v8 ad=1.4664 pd=8.3 as=0 ps=0 w=3.76 l=1.62
X1 B.t12 B.t10 B.t11 B.t3 sky130_fd_pr__nfet_01v8 ad=1.4664 pd=8.3 as=0 ps=0 w=3.76 l=1.62
X2 VDD2.t1 VN.t0 VTAIL.t2 B.t0 sky130_fd_pr__nfet_01v8 ad=1.4664 pd=8.3 as=1.4664 ps=8.3 w=3.76 l=1.62
X3 B.t9 B.t6 B.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=1.4664 pd=8.3 as=0 ps=0 w=3.76 l=1.62
X4 VDD2.t0 VN.t1 VTAIL.t3 B.t1 sky130_fd_pr__nfet_01v8 ad=1.4664 pd=8.3 as=1.4664 ps=8.3 w=3.76 l=1.62
X5 B.t5 B.t2 B.t4 B.t3 sky130_fd_pr__nfet_01v8 ad=1.4664 pd=8.3 as=0 ps=0 w=3.76 l=1.62
X6 VDD1.t1 VP.t0 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=1.4664 pd=8.3 as=1.4664 ps=8.3 w=3.76 l=1.62
X7 VDD1.t0 VP.t1 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=1.4664 pd=8.3 as=1.4664 ps=8.3 w=3.76 l=1.62
R0 B.n385 B.n384 585
R1 B.n148 B.n60 585
R2 B.n147 B.n146 585
R3 B.n145 B.n144 585
R4 B.n143 B.n142 585
R5 B.n141 B.n140 585
R6 B.n139 B.n138 585
R7 B.n137 B.n136 585
R8 B.n135 B.n134 585
R9 B.n133 B.n132 585
R10 B.n131 B.n130 585
R11 B.n129 B.n128 585
R12 B.n127 B.n126 585
R13 B.n125 B.n124 585
R14 B.n123 B.n122 585
R15 B.n121 B.n120 585
R16 B.n119 B.n118 585
R17 B.n116 B.n115 585
R18 B.n114 B.n113 585
R19 B.n112 B.n111 585
R20 B.n110 B.n109 585
R21 B.n108 B.n107 585
R22 B.n106 B.n105 585
R23 B.n104 B.n103 585
R24 B.n102 B.n101 585
R25 B.n100 B.n99 585
R26 B.n98 B.n97 585
R27 B.n95 B.n94 585
R28 B.n93 B.n92 585
R29 B.n91 B.n90 585
R30 B.n89 B.n88 585
R31 B.n87 B.n86 585
R32 B.n85 B.n84 585
R33 B.n83 B.n82 585
R34 B.n81 B.n80 585
R35 B.n79 B.n78 585
R36 B.n77 B.n76 585
R37 B.n75 B.n74 585
R38 B.n73 B.n72 585
R39 B.n71 B.n70 585
R40 B.n69 B.n68 585
R41 B.n67 B.n66 585
R42 B.n39 B.n38 585
R43 B.n390 B.n389 585
R44 B.n383 B.n61 585
R45 B.n61 B.n36 585
R46 B.n382 B.n35 585
R47 B.n394 B.n35 585
R48 B.n381 B.n34 585
R49 B.n395 B.n34 585
R50 B.n380 B.n33 585
R51 B.n396 B.n33 585
R52 B.n379 B.n378 585
R53 B.n378 B.n29 585
R54 B.n377 B.n28 585
R55 B.n402 B.n28 585
R56 B.n376 B.n27 585
R57 B.n403 B.n27 585
R58 B.n375 B.n26 585
R59 B.n404 B.n26 585
R60 B.n374 B.n373 585
R61 B.n373 B.n22 585
R62 B.n372 B.n21 585
R63 B.n410 B.n21 585
R64 B.n371 B.n20 585
R65 B.n411 B.n20 585
R66 B.n370 B.n19 585
R67 B.n412 B.n19 585
R68 B.n369 B.n368 585
R69 B.n368 B.n15 585
R70 B.n367 B.n14 585
R71 B.n418 B.n14 585
R72 B.n366 B.n13 585
R73 B.n419 B.n13 585
R74 B.n365 B.n12 585
R75 B.n420 B.n12 585
R76 B.n364 B.n363 585
R77 B.n363 B.n362 585
R78 B.n361 B.n360 585
R79 B.n361 B.n8 585
R80 B.n359 B.n7 585
R81 B.n427 B.n7 585
R82 B.n358 B.n6 585
R83 B.n428 B.n6 585
R84 B.n357 B.n5 585
R85 B.n429 B.n5 585
R86 B.n356 B.n355 585
R87 B.n355 B.n4 585
R88 B.n354 B.n149 585
R89 B.n354 B.n353 585
R90 B.n344 B.n150 585
R91 B.n151 B.n150 585
R92 B.n346 B.n345 585
R93 B.n347 B.n346 585
R94 B.n343 B.n156 585
R95 B.n156 B.n155 585
R96 B.n342 B.n341 585
R97 B.n341 B.n340 585
R98 B.n158 B.n157 585
R99 B.n159 B.n158 585
R100 B.n333 B.n332 585
R101 B.n334 B.n333 585
R102 B.n331 B.n164 585
R103 B.n164 B.n163 585
R104 B.n330 B.n329 585
R105 B.n329 B.n328 585
R106 B.n166 B.n165 585
R107 B.n167 B.n166 585
R108 B.n321 B.n320 585
R109 B.n322 B.n321 585
R110 B.n319 B.n171 585
R111 B.n175 B.n171 585
R112 B.n318 B.n317 585
R113 B.n317 B.n316 585
R114 B.n173 B.n172 585
R115 B.n174 B.n173 585
R116 B.n309 B.n308 585
R117 B.n310 B.n309 585
R118 B.n307 B.n180 585
R119 B.n180 B.n179 585
R120 B.n306 B.n305 585
R121 B.n305 B.n304 585
R122 B.n182 B.n181 585
R123 B.n183 B.n182 585
R124 B.n300 B.n299 585
R125 B.n186 B.n185 585
R126 B.n296 B.n295 585
R127 B.n297 B.n296 585
R128 B.n294 B.n208 585
R129 B.n293 B.n292 585
R130 B.n291 B.n290 585
R131 B.n289 B.n288 585
R132 B.n287 B.n286 585
R133 B.n285 B.n284 585
R134 B.n283 B.n282 585
R135 B.n281 B.n280 585
R136 B.n279 B.n278 585
R137 B.n277 B.n276 585
R138 B.n275 B.n274 585
R139 B.n273 B.n272 585
R140 B.n271 B.n270 585
R141 B.n269 B.n268 585
R142 B.n267 B.n266 585
R143 B.n265 B.n264 585
R144 B.n263 B.n262 585
R145 B.n261 B.n260 585
R146 B.n259 B.n258 585
R147 B.n257 B.n256 585
R148 B.n255 B.n254 585
R149 B.n253 B.n252 585
R150 B.n251 B.n250 585
R151 B.n249 B.n248 585
R152 B.n247 B.n246 585
R153 B.n245 B.n244 585
R154 B.n243 B.n242 585
R155 B.n241 B.n240 585
R156 B.n239 B.n238 585
R157 B.n237 B.n236 585
R158 B.n235 B.n234 585
R159 B.n233 B.n232 585
R160 B.n231 B.n230 585
R161 B.n229 B.n228 585
R162 B.n227 B.n226 585
R163 B.n225 B.n224 585
R164 B.n223 B.n222 585
R165 B.n221 B.n220 585
R166 B.n219 B.n218 585
R167 B.n217 B.n216 585
R168 B.n215 B.n207 585
R169 B.n297 B.n207 585
R170 B.n301 B.n184 585
R171 B.n184 B.n183 585
R172 B.n303 B.n302 585
R173 B.n304 B.n303 585
R174 B.n178 B.n177 585
R175 B.n179 B.n178 585
R176 B.n312 B.n311 585
R177 B.n311 B.n310 585
R178 B.n313 B.n176 585
R179 B.n176 B.n174 585
R180 B.n315 B.n314 585
R181 B.n316 B.n315 585
R182 B.n170 B.n169 585
R183 B.n175 B.n170 585
R184 B.n324 B.n323 585
R185 B.n323 B.n322 585
R186 B.n325 B.n168 585
R187 B.n168 B.n167 585
R188 B.n327 B.n326 585
R189 B.n328 B.n327 585
R190 B.n162 B.n161 585
R191 B.n163 B.n162 585
R192 B.n336 B.n335 585
R193 B.n335 B.n334 585
R194 B.n337 B.n160 585
R195 B.n160 B.n159 585
R196 B.n339 B.n338 585
R197 B.n340 B.n339 585
R198 B.n154 B.n153 585
R199 B.n155 B.n154 585
R200 B.n349 B.n348 585
R201 B.n348 B.n347 585
R202 B.n350 B.n152 585
R203 B.n152 B.n151 585
R204 B.n352 B.n351 585
R205 B.n353 B.n352 585
R206 B.n3 B.n0 585
R207 B.n4 B.n3 585
R208 B.n426 B.n1 585
R209 B.n427 B.n426 585
R210 B.n425 B.n424 585
R211 B.n425 B.n8 585
R212 B.n423 B.n9 585
R213 B.n362 B.n9 585
R214 B.n422 B.n421 585
R215 B.n421 B.n420 585
R216 B.n11 B.n10 585
R217 B.n419 B.n11 585
R218 B.n417 B.n416 585
R219 B.n418 B.n417 585
R220 B.n415 B.n16 585
R221 B.n16 B.n15 585
R222 B.n414 B.n413 585
R223 B.n413 B.n412 585
R224 B.n18 B.n17 585
R225 B.n411 B.n18 585
R226 B.n409 B.n408 585
R227 B.n410 B.n409 585
R228 B.n407 B.n23 585
R229 B.n23 B.n22 585
R230 B.n406 B.n405 585
R231 B.n405 B.n404 585
R232 B.n25 B.n24 585
R233 B.n403 B.n25 585
R234 B.n401 B.n400 585
R235 B.n402 B.n401 585
R236 B.n399 B.n30 585
R237 B.n30 B.n29 585
R238 B.n398 B.n397 585
R239 B.n397 B.n396 585
R240 B.n32 B.n31 585
R241 B.n395 B.n32 585
R242 B.n393 B.n392 585
R243 B.n394 B.n393 585
R244 B.n391 B.n37 585
R245 B.n37 B.n36 585
R246 B.n430 B.n429 585
R247 B.n428 B.n2 585
R248 B.n389 B.n37 540.549
R249 B.n385 B.n61 540.549
R250 B.n207 B.n182 540.549
R251 B.n299 B.n184 540.549
R252 B.n64 B.t6 261.796
R253 B.n62 B.t13 261.796
R254 B.n212 B.t2 261.796
R255 B.n209 B.t10 261.796
R256 B.n387 B.n386 256.663
R257 B.n387 B.n59 256.663
R258 B.n387 B.n58 256.663
R259 B.n387 B.n57 256.663
R260 B.n387 B.n56 256.663
R261 B.n387 B.n55 256.663
R262 B.n387 B.n54 256.663
R263 B.n387 B.n53 256.663
R264 B.n387 B.n52 256.663
R265 B.n387 B.n51 256.663
R266 B.n387 B.n50 256.663
R267 B.n387 B.n49 256.663
R268 B.n387 B.n48 256.663
R269 B.n387 B.n47 256.663
R270 B.n387 B.n46 256.663
R271 B.n387 B.n45 256.663
R272 B.n387 B.n44 256.663
R273 B.n387 B.n43 256.663
R274 B.n387 B.n42 256.663
R275 B.n387 B.n41 256.663
R276 B.n387 B.n40 256.663
R277 B.n388 B.n387 256.663
R278 B.n298 B.n297 256.663
R279 B.n297 B.n187 256.663
R280 B.n297 B.n188 256.663
R281 B.n297 B.n189 256.663
R282 B.n297 B.n190 256.663
R283 B.n297 B.n191 256.663
R284 B.n297 B.n192 256.663
R285 B.n297 B.n193 256.663
R286 B.n297 B.n194 256.663
R287 B.n297 B.n195 256.663
R288 B.n297 B.n196 256.663
R289 B.n297 B.n197 256.663
R290 B.n297 B.n198 256.663
R291 B.n297 B.n199 256.663
R292 B.n297 B.n200 256.663
R293 B.n297 B.n201 256.663
R294 B.n297 B.n202 256.663
R295 B.n297 B.n203 256.663
R296 B.n297 B.n204 256.663
R297 B.n297 B.n205 256.663
R298 B.n297 B.n206 256.663
R299 B.n432 B.n431 256.663
R300 B.n62 B.t14 178.423
R301 B.n212 B.t5 178.423
R302 B.n64 B.t8 178.423
R303 B.n209 B.t12 178.423
R304 B.n66 B.n39 163.367
R305 B.n70 B.n69 163.367
R306 B.n74 B.n73 163.367
R307 B.n78 B.n77 163.367
R308 B.n82 B.n81 163.367
R309 B.n86 B.n85 163.367
R310 B.n90 B.n89 163.367
R311 B.n94 B.n93 163.367
R312 B.n99 B.n98 163.367
R313 B.n103 B.n102 163.367
R314 B.n107 B.n106 163.367
R315 B.n111 B.n110 163.367
R316 B.n115 B.n114 163.367
R317 B.n120 B.n119 163.367
R318 B.n124 B.n123 163.367
R319 B.n128 B.n127 163.367
R320 B.n132 B.n131 163.367
R321 B.n136 B.n135 163.367
R322 B.n140 B.n139 163.367
R323 B.n144 B.n143 163.367
R324 B.n146 B.n60 163.367
R325 B.n305 B.n182 163.367
R326 B.n305 B.n180 163.367
R327 B.n309 B.n180 163.367
R328 B.n309 B.n173 163.367
R329 B.n317 B.n173 163.367
R330 B.n317 B.n171 163.367
R331 B.n321 B.n171 163.367
R332 B.n321 B.n166 163.367
R333 B.n329 B.n166 163.367
R334 B.n329 B.n164 163.367
R335 B.n333 B.n164 163.367
R336 B.n333 B.n158 163.367
R337 B.n341 B.n158 163.367
R338 B.n341 B.n156 163.367
R339 B.n346 B.n156 163.367
R340 B.n346 B.n150 163.367
R341 B.n354 B.n150 163.367
R342 B.n355 B.n354 163.367
R343 B.n355 B.n5 163.367
R344 B.n6 B.n5 163.367
R345 B.n7 B.n6 163.367
R346 B.n361 B.n7 163.367
R347 B.n363 B.n361 163.367
R348 B.n363 B.n12 163.367
R349 B.n13 B.n12 163.367
R350 B.n14 B.n13 163.367
R351 B.n368 B.n14 163.367
R352 B.n368 B.n19 163.367
R353 B.n20 B.n19 163.367
R354 B.n21 B.n20 163.367
R355 B.n373 B.n21 163.367
R356 B.n373 B.n26 163.367
R357 B.n27 B.n26 163.367
R358 B.n28 B.n27 163.367
R359 B.n378 B.n28 163.367
R360 B.n378 B.n33 163.367
R361 B.n34 B.n33 163.367
R362 B.n35 B.n34 163.367
R363 B.n61 B.n35 163.367
R364 B.n296 B.n186 163.367
R365 B.n296 B.n208 163.367
R366 B.n292 B.n291 163.367
R367 B.n288 B.n287 163.367
R368 B.n284 B.n283 163.367
R369 B.n280 B.n279 163.367
R370 B.n276 B.n275 163.367
R371 B.n272 B.n271 163.367
R372 B.n268 B.n267 163.367
R373 B.n264 B.n263 163.367
R374 B.n260 B.n259 163.367
R375 B.n256 B.n255 163.367
R376 B.n252 B.n251 163.367
R377 B.n248 B.n247 163.367
R378 B.n244 B.n243 163.367
R379 B.n240 B.n239 163.367
R380 B.n236 B.n235 163.367
R381 B.n232 B.n231 163.367
R382 B.n228 B.n227 163.367
R383 B.n224 B.n223 163.367
R384 B.n220 B.n219 163.367
R385 B.n216 B.n207 163.367
R386 B.n303 B.n184 163.367
R387 B.n303 B.n178 163.367
R388 B.n311 B.n178 163.367
R389 B.n311 B.n176 163.367
R390 B.n315 B.n176 163.367
R391 B.n315 B.n170 163.367
R392 B.n323 B.n170 163.367
R393 B.n323 B.n168 163.367
R394 B.n327 B.n168 163.367
R395 B.n327 B.n162 163.367
R396 B.n335 B.n162 163.367
R397 B.n335 B.n160 163.367
R398 B.n339 B.n160 163.367
R399 B.n339 B.n154 163.367
R400 B.n348 B.n154 163.367
R401 B.n348 B.n152 163.367
R402 B.n352 B.n152 163.367
R403 B.n352 B.n3 163.367
R404 B.n430 B.n3 163.367
R405 B.n426 B.n2 163.367
R406 B.n426 B.n425 163.367
R407 B.n425 B.n9 163.367
R408 B.n421 B.n9 163.367
R409 B.n421 B.n11 163.367
R410 B.n417 B.n11 163.367
R411 B.n417 B.n16 163.367
R412 B.n413 B.n16 163.367
R413 B.n413 B.n18 163.367
R414 B.n409 B.n18 163.367
R415 B.n409 B.n23 163.367
R416 B.n405 B.n23 163.367
R417 B.n405 B.n25 163.367
R418 B.n401 B.n25 163.367
R419 B.n401 B.n30 163.367
R420 B.n397 B.n30 163.367
R421 B.n397 B.n32 163.367
R422 B.n393 B.n32 163.367
R423 B.n393 B.n37 163.367
R424 B.n297 B.n183 157.056
R425 B.n387 B.n36 157.056
R426 B.n63 B.t15 140.606
R427 B.n213 B.t4 140.606
R428 B.n65 B.t9 140.606
R429 B.n210 B.t11 140.606
R430 B.n304 B.n183 82.7897
R431 B.n304 B.n179 82.7897
R432 B.n310 B.n179 82.7897
R433 B.n310 B.n174 82.7897
R434 B.n316 B.n174 82.7897
R435 B.n316 B.n175 82.7897
R436 B.n322 B.n167 82.7897
R437 B.n328 B.n167 82.7897
R438 B.n328 B.n163 82.7897
R439 B.n334 B.n163 82.7897
R440 B.n334 B.n159 82.7897
R441 B.n340 B.n159 82.7897
R442 B.n340 B.n155 82.7897
R443 B.n347 B.n155 82.7897
R444 B.n353 B.n151 82.7897
R445 B.n353 B.n4 82.7897
R446 B.n429 B.n4 82.7897
R447 B.n429 B.n428 82.7897
R448 B.n428 B.n427 82.7897
R449 B.n427 B.n8 82.7897
R450 B.n362 B.n8 82.7897
R451 B.n420 B.n419 82.7897
R452 B.n419 B.n418 82.7897
R453 B.n418 B.n15 82.7897
R454 B.n412 B.n15 82.7897
R455 B.n412 B.n411 82.7897
R456 B.n411 B.n410 82.7897
R457 B.n410 B.n22 82.7897
R458 B.n404 B.n22 82.7897
R459 B.n403 B.n402 82.7897
R460 B.n402 B.n29 82.7897
R461 B.n396 B.n29 82.7897
R462 B.n396 B.n395 82.7897
R463 B.n395 B.n394 82.7897
R464 B.n394 B.n36 82.7897
R465 B.t1 B.n151 80.3547
R466 B.n362 B.t0 80.3547
R467 B.n322 B.t3 75.4847
R468 B.n404 B.t7 75.4847
R469 B.n389 B.n388 71.676
R470 B.n66 B.n40 71.676
R471 B.n70 B.n41 71.676
R472 B.n74 B.n42 71.676
R473 B.n78 B.n43 71.676
R474 B.n82 B.n44 71.676
R475 B.n86 B.n45 71.676
R476 B.n90 B.n46 71.676
R477 B.n94 B.n47 71.676
R478 B.n99 B.n48 71.676
R479 B.n103 B.n49 71.676
R480 B.n107 B.n50 71.676
R481 B.n111 B.n51 71.676
R482 B.n115 B.n52 71.676
R483 B.n120 B.n53 71.676
R484 B.n124 B.n54 71.676
R485 B.n128 B.n55 71.676
R486 B.n132 B.n56 71.676
R487 B.n136 B.n57 71.676
R488 B.n140 B.n58 71.676
R489 B.n144 B.n59 71.676
R490 B.n386 B.n60 71.676
R491 B.n386 B.n385 71.676
R492 B.n146 B.n59 71.676
R493 B.n143 B.n58 71.676
R494 B.n139 B.n57 71.676
R495 B.n135 B.n56 71.676
R496 B.n131 B.n55 71.676
R497 B.n127 B.n54 71.676
R498 B.n123 B.n53 71.676
R499 B.n119 B.n52 71.676
R500 B.n114 B.n51 71.676
R501 B.n110 B.n50 71.676
R502 B.n106 B.n49 71.676
R503 B.n102 B.n48 71.676
R504 B.n98 B.n47 71.676
R505 B.n93 B.n46 71.676
R506 B.n89 B.n45 71.676
R507 B.n85 B.n44 71.676
R508 B.n81 B.n43 71.676
R509 B.n77 B.n42 71.676
R510 B.n73 B.n41 71.676
R511 B.n69 B.n40 71.676
R512 B.n388 B.n39 71.676
R513 B.n299 B.n298 71.676
R514 B.n208 B.n187 71.676
R515 B.n291 B.n188 71.676
R516 B.n287 B.n189 71.676
R517 B.n283 B.n190 71.676
R518 B.n279 B.n191 71.676
R519 B.n275 B.n192 71.676
R520 B.n271 B.n193 71.676
R521 B.n267 B.n194 71.676
R522 B.n263 B.n195 71.676
R523 B.n259 B.n196 71.676
R524 B.n255 B.n197 71.676
R525 B.n251 B.n198 71.676
R526 B.n247 B.n199 71.676
R527 B.n243 B.n200 71.676
R528 B.n239 B.n201 71.676
R529 B.n235 B.n202 71.676
R530 B.n231 B.n203 71.676
R531 B.n227 B.n204 71.676
R532 B.n223 B.n205 71.676
R533 B.n219 B.n206 71.676
R534 B.n298 B.n186 71.676
R535 B.n292 B.n187 71.676
R536 B.n288 B.n188 71.676
R537 B.n284 B.n189 71.676
R538 B.n280 B.n190 71.676
R539 B.n276 B.n191 71.676
R540 B.n272 B.n192 71.676
R541 B.n268 B.n193 71.676
R542 B.n264 B.n194 71.676
R543 B.n260 B.n195 71.676
R544 B.n256 B.n196 71.676
R545 B.n252 B.n197 71.676
R546 B.n248 B.n198 71.676
R547 B.n244 B.n199 71.676
R548 B.n240 B.n200 71.676
R549 B.n236 B.n201 71.676
R550 B.n232 B.n202 71.676
R551 B.n228 B.n203 71.676
R552 B.n224 B.n204 71.676
R553 B.n220 B.n205 71.676
R554 B.n216 B.n206 71.676
R555 B.n431 B.n430 71.676
R556 B.n431 B.n2 71.676
R557 B.n96 B.n65 59.5399
R558 B.n117 B.n63 59.5399
R559 B.n214 B.n213 59.5399
R560 B.n211 B.n210 59.5399
R561 B.n65 B.n64 37.8187
R562 B.n63 B.n62 37.8187
R563 B.n213 B.n212 37.8187
R564 B.n210 B.n209 37.8187
R565 B.n301 B.n300 35.1225
R566 B.n215 B.n181 35.1225
R567 B.n391 B.n390 35.1225
R568 B.n384 B.n383 35.1224
R569 B B.n432 18.0485
R570 B.n302 B.n301 10.6151
R571 B.n302 B.n177 10.6151
R572 B.n312 B.n177 10.6151
R573 B.n313 B.n312 10.6151
R574 B.n314 B.n313 10.6151
R575 B.n314 B.n169 10.6151
R576 B.n324 B.n169 10.6151
R577 B.n325 B.n324 10.6151
R578 B.n326 B.n325 10.6151
R579 B.n326 B.n161 10.6151
R580 B.n336 B.n161 10.6151
R581 B.n337 B.n336 10.6151
R582 B.n338 B.n337 10.6151
R583 B.n338 B.n153 10.6151
R584 B.n349 B.n153 10.6151
R585 B.n350 B.n349 10.6151
R586 B.n351 B.n350 10.6151
R587 B.n351 B.n0 10.6151
R588 B.n300 B.n185 10.6151
R589 B.n295 B.n185 10.6151
R590 B.n295 B.n294 10.6151
R591 B.n294 B.n293 10.6151
R592 B.n293 B.n290 10.6151
R593 B.n290 B.n289 10.6151
R594 B.n289 B.n286 10.6151
R595 B.n286 B.n285 10.6151
R596 B.n285 B.n282 10.6151
R597 B.n282 B.n281 10.6151
R598 B.n281 B.n278 10.6151
R599 B.n278 B.n277 10.6151
R600 B.n277 B.n274 10.6151
R601 B.n274 B.n273 10.6151
R602 B.n273 B.n270 10.6151
R603 B.n270 B.n269 10.6151
R604 B.n266 B.n265 10.6151
R605 B.n265 B.n262 10.6151
R606 B.n262 B.n261 10.6151
R607 B.n261 B.n258 10.6151
R608 B.n258 B.n257 10.6151
R609 B.n257 B.n254 10.6151
R610 B.n254 B.n253 10.6151
R611 B.n253 B.n250 10.6151
R612 B.n250 B.n249 10.6151
R613 B.n246 B.n245 10.6151
R614 B.n245 B.n242 10.6151
R615 B.n242 B.n241 10.6151
R616 B.n241 B.n238 10.6151
R617 B.n238 B.n237 10.6151
R618 B.n237 B.n234 10.6151
R619 B.n234 B.n233 10.6151
R620 B.n233 B.n230 10.6151
R621 B.n230 B.n229 10.6151
R622 B.n229 B.n226 10.6151
R623 B.n226 B.n225 10.6151
R624 B.n225 B.n222 10.6151
R625 B.n222 B.n221 10.6151
R626 B.n221 B.n218 10.6151
R627 B.n218 B.n217 10.6151
R628 B.n217 B.n215 10.6151
R629 B.n306 B.n181 10.6151
R630 B.n307 B.n306 10.6151
R631 B.n308 B.n307 10.6151
R632 B.n308 B.n172 10.6151
R633 B.n318 B.n172 10.6151
R634 B.n319 B.n318 10.6151
R635 B.n320 B.n319 10.6151
R636 B.n320 B.n165 10.6151
R637 B.n330 B.n165 10.6151
R638 B.n331 B.n330 10.6151
R639 B.n332 B.n331 10.6151
R640 B.n332 B.n157 10.6151
R641 B.n342 B.n157 10.6151
R642 B.n343 B.n342 10.6151
R643 B.n345 B.n343 10.6151
R644 B.n345 B.n344 10.6151
R645 B.n344 B.n149 10.6151
R646 B.n356 B.n149 10.6151
R647 B.n357 B.n356 10.6151
R648 B.n358 B.n357 10.6151
R649 B.n359 B.n358 10.6151
R650 B.n360 B.n359 10.6151
R651 B.n364 B.n360 10.6151
R652 B.n365 B.n364 10.6151
R653 B.n366 B.n365 10.6151
R654 B.n367 B.n366 10.6151
R655 B.n369 B.n367 10.6151
R656 B.n370 B.n369 10.6151
R657 B.n371 B.n370 10.6151
R658 B.n372 B.n371 10.6151
R659 B.n374 B.n372 10.6151
R660 B.n375 B.n374 10.6151
R661 B.n376 B.n375 10.6151
R662 B.n377 B.n376 10.6151
R663 B.n379 B.n377 10.6151
R664 B.n380 B.n379 10.6151
R665 B.n381 B.n380 10.6151
R666 B.n382 B.n381 10.6151
R667 B.n383 B.n382 10.6151
R668 B.n424 B.n1 10.6151
R669 B.n424 B.n423 10.6151
R670 B.n423 B.n422 10.6151
R671 B.n422 B.n10 10.6151
R672 B.n416 B.n10 10.6151
R673 B.n416 B.n415 10.6151
R674 B.n415 B.n414 10.6151
R675 B.n414 B.n17 10.6151
R676 B.n408 B.n17 10.6151
R677 B.n408 B.n407 10.6151
R678 B.n407 B.n406 10.6151
R679 B.n406 B.n24 10.6151
R680 B.n400 B.n24 10.6151
R681 B.n400 B.n399 10.6151
R682 B.n399 B.n398 10.6151
R683 B.n398 B.n31 10.6151
R684 B.n392 B.n31 10.6151
R685 B.n392 B.n391 10.6151
R686 B.n390 B.n38 10.6151
R687 B.n67 B.n38 10.6151
R688 B.n68 B.n67 10.6151
R689 B.n71 B.n68 10.6151
R690 B.n72 B.n71 10.6151
R691 B.n75 B.n72 10.6151
R692 B.n76 B.n75 10.6151
R693 B.n79 B.n76 10.6151
R694 B.n80 B.n79 10.6151
R695 B.n83 B.n80 10.6151
R696 B.n84 B.n83 10.6151
R697 B.n87 B.n84 10.6151
R698 B.n88 B.n87 10.6151
R699 B.n91 B.n88 10.6151
R700 B.n92 B.n91 10.6151
R701 B.n95 B.n92 10.6151
R702 B.n100 B.n97 10.6151
R703 B.n101 B.n100 10.6151
R704 B.n104 B.n101 10.6151
R705 B.n105 B.n104 10.6151
R706 B.n108 B.n105 10.6151
R707 B.n109 B.n108 10.6151
R708 B.n112 B.n109 10.6151
R709 B.n113 B.n112 10.6151
R710 B.n116 B.n113 10.6151
R711 B.n121 B.n118 10.6151
R712 B.n122 B.n121 10.6151
R713 B.n125 B.n122 10.6151
R714 B.n126 B.n125 10.6151
R715 B.n129 B.n126 10.6151
R716 B.n130 B.n129 10.6151
R717 B.n133 B.n130 10.6151
R718 B.n134 B.n133 10.6151
R719 B.n137 B.n134 10.6151
R720 B.n138 B.n137 10.6151
R721 B.n141 B.n138 10.6151
R722 B.n142 B.n141 10.6151
R723 B.n145 B.n142 10.6151
R724 B.n147 B.n145 10.6151
R725 B.n148 B.n147 10.6151
R726 B.n384 B.n148 10.6151
R727 B.n269 B.n211 9.36635
R728 B.n246 B.n214 9.36635
R729 B.n96 B.n95 9.36635
R730 B.n118 B.n117 9.36635
R731 B.n432 B.n0 8.11757
R732 B.n432 B.n1 8.11757
R733 B.n175 B.t3 7.30543
R734 B.t7 B.n403 7.30543
R735 B.n347 B.t1 2.43548
R736 B.n420 B.t0 2.43548
R737 B.n266 B.n211 1.24928
R738 B.n249 B.n214 1.24928
R739 B.n97 B.n96 1.24928
R740 B.n117 B.n116 1.24928
R741 VN VN.t1 150.828
R742 VN VN.t0 115.064
R743 VTAIL.n74 VTAIL.n60 289.615
R744 VTAIL.n14 VTAIL.n0 289.615
R745 VTAIL.n54 VTAIL.n40 289.615
R746 VTAIL.n34 VTAIL.n20 289.615
R747 VTAIL.n67 VTAIL.n66 185
R748 VTAIL.n64 VTAIL.n63 185
R749 VTAIL.n73 VTAIL.n72 185
R750 VTAIL.n75 VTAIL.n74 185
R751 VTAIL.n7 VTAIL.n6 185
R752 VTAIL.n4 VTAIL.n3 185
R753 VTAIL.n13 VTAIL.n12 185
R754 VTAIL.n15 VTAIL.n14 185
R755 VTAIL.n55 VTAIL.n54 185
R756 VTAIL.n53 VTAIL.n52 185
R757 VTAIL.n44 VTAIL.n43 185
R758 VTAIL.n47 VTAIL.n46 185
R759 VTAIL.n35 VTAIL.n34 185
R760 VTAIL.n33 VTAIL.n32 185
R761 VTAIL.n24 VTAIL.n23 185
R762 VTAIL.n27 VTAIL.n26 185
R763 VTAIL.t2 VTAIL.n65 147.888
R764 VTAIL.t1 VTAIL.n5 147.888
R765 VTAIL.t0 VTAIL.n45 147.888
R766 VTAIL.t3 VTAIL.n25 147.888
R767 VTAIL.n66 VTAIL.n63 104.615
R768 VTAIL.n73 VTAIL.n63 104.615
R769 VTAIL.n74 VTAIL.n73 104.615
R770 VTAIL.n6 VTAIL.n3 104.615
R771 VTAIL.n13 VTAIL.n3 104.615
R772 VTAIL.n14 VTAIL.n13 104.615
R773 VTAIL.n54 VTAIL.n53 104.615
R774 VTAIL.n53 VTAIL.n43 104.615
R775 VTAIL.n46 VTAIL.n43 104.615
R776 VTAIL.n34 VTAIL.n33 104.615
R777 VTAIL.n33 VTAIL.n23 104.615
R778 VTAIL.n26 VTAIL.n23 104.615
R779 VTAIL.n66 VTAIL.t2 52.3082
R780 VTAIL.n6 VTAIL.t1 52.3082
R781 VTAIL.n46 VTAIL.t0 52.3082
R782 VTAIL.n26 VTAIL.t3 52.3082
R783 VTAIL.n79 VTAIL.n78 30.6338
R784 VTAIL.n19 VTAIL.n18 30.6338
R785 VTAIL.n59 VTAIL.n58 30.6338
R786 VTAIL.n39 VTAIL.n38 30.6338
R787 VTAIL.n39 VTAIL.n19 18.9703
R788 VTAIL.n79 VTAIL.n59 17.2893
R789 VTAIL.n67 VTAIL.n65 15.6496
R790 VTAIL.n7 VTAIL.n5 15.6496
R791 VTAIL.n47 VTAIL.n45 15.6496
R792 VTAIL.n27 VTAIL.n25 15.6496
R793 VTAIL.n68 VTAIL.n64 12.8005
R794 VTAIL.n8 VTAIL.n4 12.8005
R795 VTAIL.n48 VTAIL.n44 12.8005
R796 VTAIL.n28 VTAIL.n24 12.8005
R797 VTAIL.n72 VTAIL.n71 12.0247
R798 VTAIL.n12 VTAIL.n11 12.0247
R799 VTAIL.n52 VTAIL.n51 12.0247
R800 VTAIL.n32 VTAIL.n31 12.0247
R801 VTAIL.n75 VTAIL.n62 11.249
R802 VTAIL.n15 VTAIL.n2 11.249
R803 VTAIL.n55 VTAIL.n42 11.249
R804 VTAIL.n35 VTAIL.n22 11.249
R805 VTAIL.n76 VTAIL.n60 10.4732
R806 VTAIL.n16 VTAIL.n0 10.4732
R807 VTAIL.n56 VTAIL.n40 10.4732
R808 VTAIL.n36 VTAIL.n20 10.4732
R809 VTAIL.n78 VTAIL.n77 9.45567
R810 VTAIL.n18 VTAIL.n17 9.45567
R811 VTAIL.n58 VTAIL.n57 9.45567
R812 VTAIL.n38 VTAIL.n37 9.45567
R813 VTAIL.n77 VTAIL.n76 9.3005
R814 VTAIL.n62 VTAIL.n61 9.3005
R815 VTAIL.n71 VTAIL.n70 9.3005
R816 VTAIL.n69 VTAIL.n68 9.3005
R817 VTAIL.n17 VTAIL.n16 9.3005
R818 VTAIL.n2 VTAIL.n1 9.3005
R819 VTAIL.n11 VTAIL.n10 9.3005
R820 VTAIL.n9 VTAIL.n8 9.3005
R821 VTAIL.n57 VTAIL.n56 9.3005
R822 VTAIL.n42 VTAIL.n41 9.3005
R823 VTAIL.n51 VTAIL.n50 9.3005
R824 VTAIL.n49 VTAIL.n48 9.3005
R825 VTAIL.n37 VTAIL.n36 9.3005
R826 VTAIL.n22 VTAIL.n21 9.3005
R827 VTAIL.n31 VTAIL.n30 9.3005
R828 VTAIL.n29 VTAIL.n28 9.3005
R829 VTAIL.n69 VTAIL.n65 4.40546
R830 VTAIL.n9 VTAIL.n5 4.40546
R831 VTAIL.n49 VTAIL.n45 4.40546
R832 VTAIL.n29 VTAIL.n25 4.40546
R833 VTAIL.n78 VTAIL.n60 3.49141
R834 VTAIL.n18 VTAIL.n0 3.49141
R835 VTAIL.n58 VTAIL.n40 3.49141
R836 VTAIL.n38 VTAIL.n20 3.49141
R837 VTAIL.n76 VTAIL.n75 2.71565
R838 VTAIL.n16 VTAIL.n15 2.71565
R839 VTAIL.n56 VTAIL.n55 2.71565
R840 VTAIL.n36 VTAIL.n35 2.71565
R841 VTAIL.n72 VTAIL.n62 1.93989
R842 VTAIL.n12 VTAIL.n2 1.93989
R843 VTAIL.n52 VTAIL.n42 1.93989
R844 VTAIL.n32 VTAIL.n22 1.93989
R845 VTAIL.n59 VTAIL.n39 1.31084
R846 VTAIL.n71 VTAIL.n64 1.16414
R847 VTAIL.n11 VTAIL.n4 1.16414
R848 VTAIL.n51 VTAIL.n44 1.16414
R849 VTAIL.n31 VTAIL.n24 1.16414
R850 VTAIL VTAIL.n19 0.948776
R851 VTAIL.n68 VTAIL.n67 0.388379
R852 VTAIL.n8 VTAIL.n7 0.388379
R853 VTAIL.n48 VTAIL.n47 0.388379
R854 VTAIL.n28 VTAIL.n27 0.388379
R855 VTAIL VTAIL.n79 0.362569
R856 VTAIL.n70 VTAIL.n69 0.155672
R857 VTAIL.n70 VTAIL.n61 0.155672
R858 VTAIL.n77 VTAIL.n61 0.155672
R859 VTAIL.n10 VTAIL.n9 0.155672
R860 VTAIL.n10 VTAIL.n1 0.155672
R861 VTAIL.n17 VTAIL.n1 0.155672
R862 VTAIL.n57 VTAIL.n41 0.155672
R863 VTAIL.n50 VTAIL.n41 0.155672
R864 VTAIL.n50 VTAIL.n49 0.155672
R865 VTAIL.n37 VTAIL.n21 0.155672
R866 VTAIL.n30 VTAIL.n21 0.155672
R867 VTAIL.n30 VTAIL.n29 0.155672
R868 VDD2.n33 VDD2.n19 289.615
R869 VDD2.n14 VDD2.n0 289.615
R870 VDD2.n34 VDD2.n33 185
R871 VDD2.n32 VDD2.n31 185
R872 VDD2.n23 VDD2.n22 185
R873 VDD2.n26 VDD2.n25 185
R874 VDD2.n7 VDD2.n6 185
R875 VDD2.n4 VDD2.n3 185
R876 VDD2.n13 VDD2.n12 185
R877 VDD2.n15 VDD2.n14 185
R878 VDD2.t0 VDD2.n24 147.888
R879 VDD2.t1 VDD2.n5 147.888
R880 VDD2.n33 VDD2.n32 104.615
R881 VDD2.n32 VDD2.n22 104.615
R882 VDD2.n25 VDD2.n22 104.615
R883 VDD2.n6 VDD2.n3 104.615
R884 VDD2.n13 VDD2.n3 104.615
R885 VDD2.n14 VDD2.n13 104.615
R886 VDD2.n38 VDD2.n18 77.5755
R887 VDD2.n25 VDD2.t0 52.3082
R888 VDD2.n6 VDD2.t1 52.3082
R889 VDD2.n38 VDD2.n37 47.3126
R890 VDD2.n26 VDD2.n24 15.6496
R891 VDD2.n7 VDD2.n5 15.6496
R892 VDD2.n27 VDD2.n23 12.8005
R893 VDD2.n8 VDD2.n4 12.8005
R894 VDD2.n31 VDD2.n30 12.0247
R895 VDD2.n12 VDD2.n11 12.0247
R896 VDD2.n34 VDD2.n21 11.249
R897 VDD2.n15 VDD2.n2 11.249
R898 VDD2.n35 VDD2.n19 10.4732
R899 VDD2.n16 VDD2.n0 10.4732
R900 VDD2.n37 VDD2.n36 9.45567
R901 VDD2.n18 VDD2.n17 9.45567
R902 VDD2.n36 VDD2.n35 9.3005
R903 VDD2.n21 VDD2.n20 9.3005
R904 VDD2.n30 VDD2.n29 9.3005
R905 VDD2.n28 VDD2.n27 9.3005
R906 VDD2.n17 VDD2.n16 9.3005
R907 VDD2.n2 VDD2.n1 9.3005
R908 VDD2.n11 VDD2.n10 9.3005
R909 VDD2.n9 VDD2.n8 9.3005
R910 VDD2.n28 VDD2.n24 4.40546
R911 VDD2.n9 VDD2.n5 4.40546
R912 VDD2.n37 VDD2.n19 3.49141
R913 VDD2.n18 VDD2.n0 3.49141
R914 VDD2.n35 VDD2.n34 2.71565
R915 VDD2.n16 VDD2.n15 2.71565
R916 VDD2.n31 VDD2.n21 1.93989
R917 VDD2.n12 VDD2.n2 1.93989
R918 VDD2.n30 VDD2.n23 1.16414
R919 VDD2.n11 VDD2.n4 1.16414
R920 VDD2 VDD2.n38 0.478948
R921 VDD2.n27 VDD2.n26 0.388379
R922 VDD2.n8 VDD2.n7 0.388379
R923 VDD2.n36 VDD2.n20 0.155672
R924 VDD2.n29 VDD2.n20 0.155672
R925 VDD2.n29 VDD2.n28 0.155672
R926 VDD2.n10 VDD2.n9 0.155672
R927 VDD2.n10 VDD2.n1 0.155672
R928 VDD2.n17 VDD2.n1 0.155672
R929 VP.n0 VP.t0 150.637
R930 VP.n0 VP.t1 114.823
R931 VP VP.n0 0.241678
R932 VDD1.n14 VDD1.n0 289.615
R933 VDD1.n33 VDD1.n19 289.615
R934 VDD1.n15 VDD1.n14 185
R935 VDD1.n13 VDD1.n12 185
R936 VDD1.n4 VDD1.n3 185
R937 VDD1.n7 VDD1.n6 185
R938 VDD1.n26 VDD1.n25 185
R939 VDD1.n23 VDD1.n22 185
R940 VDD1.n32 VDD1.n31 185
R941 VDD1.n34 VDD1.n33 185
R942 VDD1.t1 VDD1.n5 147.888
R943 VDD1.t0 VDD1.n24 147.888
R944 VDD1.n14 VDD1.n13 104.615
R945 VDD1.n13 VDD1.n3 104.615
R946 VDD1.n6 VDD1.n3 104.615
R947 VDD1.n25 VDD1.n22 104.615
R948 VDD1.n32 VDD1.n22 104.615
R949 VDD1.n33 VDD1.n32 104.615
R950 VDD1 VDD1.n37 78.5206
R951 VDD1.n6 VDD1.t1 52.3082
R952 VDD1.n25 VDD1.t0 52.3082
R953 VDD1 VDD1.n18 47.7911
R954 VDD1.n7 VDD1.n5 15.6496
R955 VDD1.n26 VDD1.n24 15.6496
R956 VDD1.n8 VDD1.n4 12.8005
R957 VDD1.n27 VDD1.n23 12.8005
R958 VDD1.n12 VDD1.n11 12.0247
R959 VDD1.n31 VDD1.n30 12.0247
R960 VDD1.n15 VDD1.n2 11.249
R961 VDD1.n34 VDD1.n21 11.249
R962 VDD1.n16 VDD1.n0 10.4732
R963 VDD1.n35 VDD1.n19 10.4732
R964 VDD1.n18 VDD1.n17 9.45567
R965 VDD1.n37 VDD1.n36 9.45567
R966 VDD1.n17 VDD1.n16 9.3005
R967 VDD1.n2 VDD1.n1 9.3005
R968 VDD1.n11 VDD1.n10 9.3005
R969 VDD1.n9 VDD1.n8 9.3005
R970 VDD1.n36 VDD1.n35 9.3005
R971 VDD1.n21 VDD1.n20 9.3005
R972 VDD1.n30 VDD1.n29 9.3005
R973 VDD1.n28 VDD1.n27 9.3005
R974 VDD1.n9 VDD1.n5 4.40546
R975 VDD1.n28 VDD1.n24 4.40546
R976 VDD1.n18 VDD1.n0 3.49141
R977 VDD1.n37 VDD1.n19 3.49141
R978 VDD1.n16 VDD1.n15 2.71565
R979 VDD1.n35 VDD1.n34 2.71565
R980 VDD1.n12 VDD1.n2 1.93989
R981 VDD1.n31 VDD1.n21 1.93989
R982 VDD1.n11 VDD1.n4 1.16414
R983 VDD1.n30 VDD1.n23 1.16414
R984 VDD1.n8 VDD1.n7 0.388379
R985 VDD1.n27 VDD1.n26 0.388379
R986 VDD1.n17 VDD1.n1 0.155672
R987 VDD1.n10 VDD1.n1 0.155672
R988 VDD1.n10 VDD1.n9 0.155672
R989 VDD1.n29 VDD1.n28 0.155672
R990 VDD1.n29 VDD1.n20 0.155672
R991 VDD1.n36 VDD1.n20 0.155672
C0 VTAIL VN 1.00845f
C1 VDD2 VP 0.296232f
C2 VDD2 VDD1 0.558246f
C3 VDD2 VN 0.967203f
C4 VP VDD1 1.10941f
C5 VDD2 VTAIL 2.68823f
C6 VP VN 3.47679f
C7 VP VTAIL 1.02265f
C8 VDD1 VN 0.152403f
C9 VTAIL VDD1 2.64276f
C10 VDD2 B 2.571186f
C11 VDD1 B 3.93709f
C12 VTAIL B 3.422646f
C13 VN B 6.59205f
C14 VP B 4.497505f
C15 VDD1.n0 B 0.018764f
C16 VDD1.n1 B 0.014767f
C17 VDD1.n2 B 0.007935f
C18 VDD1.n3 B 0.018756f
C19 VDD1.n4 B 0.008402f
C20 VDD1.n5 B 0.055491f
C21 VDD1.t1 B 0.030841f
C22 VDD1.n6 B 0.014067f
C23 VDD1.n7 B 0.011039f
C24 VDD1.n8 B 0.007935f
C25 VDD1.n9 B 0.198836f
C26 VDD1.n10 B 0.014767f
C27 VDD1.n11 B 0.007935f
C28 VDD1.n12 B 0.008402f
C29 VDD1.n13 B 0.018756f
C30 VDD1.n14 B 0.03708f
C31 VDD1.n15 B 0.008402f
C32 VDD1.n16 B 0.007935f
C33 VDD1.n17 B 0.03252f
C34 VDD1.n18 B 0.031048f
C35 VDD1.n19 B 0.018764f
C36 VDD1.n20 B 0.014767f
C37 VDD1.n21 B 0.007935f
C38 VDD1.n22 B 0.018756f
C39 VDD1.n23 B 0.008402f
C40 VDD1.n24 B 0.055491f
C41 VDD1.t0 B 0.030841f
C42 VDD1.n25 B 0.014067f
C43 VDD1.n26 B 0.011039f
C44 VDD1.n27 B 0.007935f
C45 VDD1.n28 B 0.198836f
C46 VDD1.n29 B 0.014767f
C47 VDD1.n30 B 0.007935f
C48 VDD1.n31 B 0.008402f
C49 VDD1.n32 B 0.018756f
C50 VDD1.n33 B 0.03708f
C51 VDD1.n34 B 0.008402f
C52 VDD1.n35 B 0.007935f
C53 VDD1.n36 B 0.03252f
C54 VDD1.n37 B 0.266504f
C55 VP.t0 B 0.882837f
C56 VP.t1 B 0.616895f
C57 VP.n0 B 1.96034f
C58 VDD2.n0 B 0.019903f
C59 VDD2.n1 B 0.015664f
C60 VDD2.n2 B 0.008417f
C61 VDD2.n3 B 0.019895f
C62 VDD2.n4 B 0.008912f
C63 VDD2.n5 B 0.05886f
C64 VDD2.t1 B 0.032713f
C65 VDD2.n6 B 0.014921f
C66 VDD2.n7 B 0.011709f
C67 VDD2.n8 B 0.008417f
C68 VDD2.n9 B 0.210908f
C69 VDD2.n10 B 0.015664f
C70 VDD2.n11 B 0.008417f
C71 VDD2.n12 B 0.008912f
C72 VDD2.n13 B 0.019895f
C73 VDD2.n14 B 0.039331f
C74 VDD2.n15 B 0.008912f
C75 VDD2.n16 B 0.008417f
C76 VDD2.n17 B 0.034494f
C77 VDD2.n18 B 0.261042f
C78 VDD2.n19 B 0.019903f
C79 VDD2.n20 B 0.015664f
C80 VDD2.n21 B 0.008417f
C81 VDD2.n22 B 0.019895f
C82 VDD2.n23 B 0.008912f
C83 VDD2.n24 B 0.05886f
C84 VDD2.t0 B 0.032713f
C85 VDD2.n25 B 0.014921f
C86 VDD2.n26 B 0.011709f
C87 VDD2.n27 B 0.008417f
C88 VDD2.n28 B 0.210908f
C89 VDD2.n29 B 0.015664f
C90 VDD2.n30 B 0.008417f
C91 VDD2.n31 B 0.008912f
C92 VDD2.n32 B 0.019895f
C93 VDD2.n33 B 0.039331f
C94 VDD2.n34 B 0.008912f
C95 VDD2.n35 B 0.008417f
C96 VDD2.n36 B 0.034494f
C97 VDD2.n37 B 0.032399f
C98 VDD2.n38 B 1.23083f
C99 VTAIL.n0 B 0.022771f
C100 VTAIL.n1 B 0.017921f
C101 VTAIL.n2 B 0.00963f
C102 VTAIL.n3 B 0.022761f
C103 VTAIL.n4 B 0.010196f
C104 VTAIL.n5 B 0.067341f
C105 VTAIL.t1 B 0.037427f
C106 VTAIL.n6 B 0.017071f
C107 VTAIL.n7 B 0.013397f
C108 VTAIL.n8 B 0.00963f
C109 VTAIL.n9 B 0.241299f
C110 VTAIL.n10 B 0.017921f
C111 VTAIL.n11 B 0.00963f
C112 VTAIL.n12 B 0.010196f
C113 VTAIL.n13 B 0.022761f
C114 VTAIL.n14 B 0.044999f
C115 VTAIL.n15 B 0.010196f
C116 VTAIL.n16 B 0.00963f
C117 VTAIL.n17 B 0.039465f
C118 VTAIL.n18 B 0.024677f
C119 VTAIL.n19 B 0.693708f
C120 VTAIL.n20 B 0.022771f
C121 VTAIL.n21 B 0.017921f
C122 VTAIL.n22 B 0.00963f
C123 VTAIL.n23 B 0.022761f
C124 VTAIL.n24 B 0.010196f
C125 VTAIL.n25 B 0.067341f
C126 VTAIL.t3 B 0.037427f
C127 VTAIL.n26 B 0.017071f
C128 VTAIL.n27 B 0.013397f
C129 VTAIL.n28 B 0.00963f
C130 VTAIL.n29 B 0.241299f
C131 VTAIL.n30 B 0.017921f
C132 VTAIL.n31 B 0.00963f
C133 VTAIL.n32 B 0.010196f
C134 VTAIL.n33 B 0.022761f
C135 VTAIL.n34 B 0.044999f
C136 VTAIL.n35 B 0.010196f
C137 VTAIL.n36 B 0.00963f
C138 VTAIL.n37 B 0.039465f
C139 VTAIL.n38 B 0.024677f
C140 VTAIL.n39 B 0.714616f
C141 VTAIL.n40 B 0.022771f
C142 VTAIL.n41 B 0.017921f
C143 VTAIL.n42 B 0.00963f
C144 VTAIL.n43 B 0.022761f
C145 VTAIL.n44 B 0.010196f
C146 VTAIL.n45 B 0.067341f
C147 VTAIL.t0 B 0.037427f
C148 VTAIL.n46 B 0.017071f
C149 VTAIL.n47 B 0.013397f
C150 VTAIL.n48 B 0.00963f
C151 VTAIL.n49 B 0.241299f
C152 VTAIL.n50 B 0.017921f
C153 VTAIL.n51 B 0.00963f
C154 VTAIL.n52 B 0.010196f
C155 VTAIL.n53 B 0.022761f
C156 VTAIL.n54 B 0.044999f
C157 VTAIL.n55 B 0.010196f
C158 VTAIL.n56 B 0.00963f
C159 VTAIL.n57 B 0.039465f
C160 VTAIL.n58 B 0.024677f
C161 VTAIL.n59 B 0.617545f
C162 VTAIL.n60 B 0.022771f
C163 VTAIL.n61 B 0.017921f
C164 VTAIL.n62 B 0.00963f
C165 VTAIL.n63 B 0.022761f
C166 VTAIL.n64 B 0.010196f
C167 VTAIL.n65 B 0.067341f
C168 VTAIL.t2 B 0.037427f
C169 VTAIL.n66 B 0.017071f
C170 VTAIL.n67 B 0.013397f
C171 VTAIL.n68 B 0.00963f
C172 VTAIL.n69 B 0.241299f
C173 VTAIL.n70 B 0.017921f
C174 VTAIL.n71 B 0.00963f
C175 VTAIL.n72 B 0.010196f
C176 VTAIL.n73 B 0.022761f
C177 VTAIL.n74 B 0.044999f
C178 VTAIL.n75 B 0.010196f
C179 VTAIL.n76 B 0.00963f
C180 VTAIL.n77 B 0.039465f
C181 VTAIL.n78 B 0.024677f
C182 VTAIL.n79 B 0.562787f
C183 VN.t0 B 0.610258f
C184 VN.t1 B 0.877094f
.ends

