* NGSPICE file created from diff_pair_sample_0929.ext - technology: sky130A

.subckt diff_pair_sample_0929 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t15 VN.t0 VDD2.t6 B.t0 sky130_fd_pr__nfet_01v8 ad=1.73085 pd=10.82 as=1.73085 ps=10.82 w=10.49 l=2.08
X1 VTAIL.t14 VN.t1 VDD2.t3 B.t2 sky130_fd_pr__nfet_01v8 ad=4.0911 pd=21.76 as=1.73085 ps=10.82 w=10.49 l=2.08
X2 VDD1.t7 VP.t0 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=1.73085 pd=10.82 as=4.0911 ps=21.76 w=10.49 l=2.08
X3 VTAIL.t2 VP.t1 VDD1.t6 B.t2 sky130_fd_pr__nfet_01v8 ad=4.0911 pd=21.76 as=1.73085 ps=10.82 w=10.49 l=2.08
X4 B.t20 B.t18 B.t19 B.t15 sky130_fd_pr__nfet_01v8 ad=4.0911 pd=21.76 as=0 ps=0 w=10.49 l=2.08
X5 B.t17 B.t14 B.t16 B.t15 sky130_fd_pr__nfet_01v8 ad=4.0911 pd=21.76 as=0 ps=0 w=10.49 l=2.08
X6 B.t13 B.t11 B.t12 B.t8 sky130_fd_pr__nfet_01v8 ad=4.0911 pd=21.76 as=0 ps=0 w=10.49 l=2.08
X7 VDD1.t5 VP.t2 VTAIL.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=1.73085 pd=10.82 as=1.73085 ps=10.82 w=10.49 l=2.08
X8 VDD2.t7 VN.t2 VTAIL.t13 B.t4 sky130_fd_pr__nfet_01v8 ad=1.73085 pd=10.82 as=1.73085 ps=10.82 w=10.49 l=2.08
X9 VDD2.t2 VN.t3 VTAIL.t12 B.t5 sky130_fd_pr__nfet_01v8 ad=1.73085 pd=10.82 as=1.73085 ps=10.82 w=10.49 l=2.08
X10 VTAIL.t0 VP.t3 VDD1.t4 B.t0 sky130_fd_pr__nfet_01v8 ad=1.73085 pd=10.82 as=1.73085 ps=10.82 w=10.49 l=2.08
X11 VTAIL.t11 VN.t4 VDD2.t4 B.t3 sky130_fd_pr__nfet_01v8 ad=4.0911 pd=21.76 as=1.73085 ps=10.82 w=10.49 l=2.08
X12 VTAIL.t10 VN.t5 VDD2.t1 B.t6 sky130_fd_pr__nfet_01v8 ad=1.73085 pd=10.82 as=1.73085 ps=10.82 w=10.49 l=2.08
X13 VDD2.t5 VN.t6 VTAIL.t9 B.t1 sky130_fd_pr__nfet_01v8 ad=1.73085 pd=10.82 as=4.0911 ps=21.76 w=10.49 l=2.08
X14 VTAIL.t6 VP.t4 VDD1.t3 B.t6 sky130_fd_pr__nfet_01v8 ad=1.73085 pd=10.82 as=1.73085 ps=10.82 w=10.49 l=2.08
X15 B.t10 B.t7 B.t9 B.t8 sky130_fd_pr__nfet_01v8 ad=4.0911 pd=21.76 as=0 ps=0 w=10.49 l=2.08
X16 VDD1.t2 VP.t5 VTAIL.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=1.73085 pd=10.82 as=1.73085 ps=10.82 w=10.49 l=2.08
X17 VDD1.t1 VP.t6 VTAIL.t7 B.t21 sky130_fd_pr__nfet_01v8 ad=1.73085 pd=10.82 as=4.0911 ps=21.76 w=10.49 l=2.08
X18 VTAIL.t3 VP.t7 VDD1.t0 B.t3 sky130_fd_pr__nfet_01v8 ad=4.0911 pd=21.76 as=1.73085 ps=10.82 w=10.49 l=2.08
X19 VDD2.t0 VN.t7 VTAIL.t8 B.t21 sky130_fd_pr__nfet_01v8 ad=1.73085 pd=10.82 as=4.0911 ps=21.76 w=10.49 l=2.08
R0 VN.n43 VN.n23 161.3
R1 VN.n42 VN.n41 161.3
R2 VN.n40 VN.n24 161.3
R3 VN.n39 VN.n38 161.3
R4 VN.n37 VN.n25 161.3
R5 VN.n35 VN.n34 161.3
R6 VN.n33 VN.n26 161.3
R7 VN.n32 VN.n31 161.3
R8 VN.n30 VN.n27 161.3
R9 VN.n20 VN.n0 161.3
R10 VN.n19 VN.n18 161.3
R11 VN.n17 VN.n1 161.3
R12 VN.n16 VN.n15 161.3
R13 VN.n14 VN.n2 161.3
R14 VN.n12 VN.n11 161.3
R15 VN.n10 VN.n3 161.3
R16 VN.n9 VN.n8 161.3
R17 VN.n7 VN.n4 161.3
R18 VN.n5 VN.t1 155.309
R19 VN.n28 VN.t6 155.309
R20 VN.n6 VN.t2 121.543
R21 VN.n13 VN.t5 121.543
R22 VN.n21 VN.t7 121.543
R23 VN.n29 VN.t0 121.543
R24 VN.n36 VN.t3 121.543
R25 VN.n44 VN.t4 121.543
R26 VN.n22 VN.n21 92.8955
R27 VN.n45 VN.n44 92.8955
R28 VN.n8 VN.n3 56.5193
R29 VN.n31 VN.n26 56.5193
R30 VN.n19 VN.n1 56.0336
R31 VN.n42 VN.n24 56.0336
R32 VN.n6 VN.n5 48.1291
R33 VN.n29 VN.n28 48.1291
R34 VN VN.n45 47.6118
R35 VN.n15 VN.n1 24.9531
R36 VN.n38 VN.n24 24.9531
R37 VN.n8 VN.n7 24.4675
R38 VN.n12 VN.n3 24.4675
R39 VN.n15 VN.n14 24.4675
R40 VN.n20 VN.n19 24.4675
R41 VN.n31 VN.n30 24.4675
R42 VN.n38 VN.n37 24.4675
R43 VN.n35 VN.n26 24.4675
R44 VN.n43 VN.n42 24.4675
R45 VN.n7 VN.n6 22.2655
R46 VN.n13 VN.n12 22.2655
R47 VN.n30 VN.n29 22.2655
R48 VN.n36 VN.n35 22.2655
R49 VN.n21 VN.n20 17.8614
R50 VN.n44 VN.n43 17.8614
R51 VN.n28 VN.n27 9.16971
R52 VN.n5 VN.n4 9.16971
R53 VN.n14 VN.n13 2.20253
R54 VN.n37 VN.n36 2.20253
R55 VN.n45 VN.n23 0.278367
R56 VN.n22 VN.n0 0.278367
R57 VN.n41 VN.n23 0.189894
R58 VN.n41 VN.n40 0.189894
R59 VN.n40 VN.n39 0.189894
R60 VN.n39 VN.n25 0.189894
R61 VN.n34 VN.n25 0.189894
R62 VN.n34 VN.n33 0.189894
R63 VN.n33 VN.n32 0.189894
R64 VN.n32 VN.n27 0.189894
R65 VN.n9 VN.n4 0.189894
R66 VN.n10 VN.n9 0.189894
R67 VN.n11 VN.n10 0.189894
R68 VN.n11 VN.n2 0.189894
R69 VN.n16 VN.n2 0.189894
R70 VN.n17 VN.n16 0.189894
R71 VN.n18 VN.n17 0.189894
R72 VN.n18 VN.n0 0.189894
R73 VN VN.n22 0.153454
R74 VDD2.n2 VDD2.n1 66.7632
R75 VDD2.n2 VDD2.n0 66.7632
R76 VDD2 VDD2.n5 66.7604
R77 VDD2.n4 VDD2.n3 65.78
R78 VDD2.n4 VDD2.n2 42.1075
R79 VDD2.n5 VDD2.t6 1.88801
R80 VDD2.n5 VDD2.t5 1.88801
R81 VDD2.n3 VDD2.t4 1.88801
R82 VDD2.n3 VDD2.t2 1.88801
R83 VDD2.n1 VDD2.t1 1.88801
R84 VDD2.n1 VDD2.t0 1.88801
R85 VDD2.n0 VDD2.t3 1.88801
R86 VDD2.n0 VDD2.t7 1.88801
R87 VDD2 VDD2.n4 1.09748
R88 VTAIL.n11 VTAIL.t2 50.9887
R89 VTAIL.n10 VTAIL.t9 50.9887
R90 VTAIL.n7 VTAIL.t11 50.9887
R91 VTAIL.n15 VTAIL.t8 50.9885
R92 VTAIL.n2 VTAIL.t14 50.9885
R93 VTAIL.n3 VTAIL.t1 50.9885
R94 VTAIL.n6 VTAIL.t3 50.9885
R95 VTAIL.n14 VTAIL.t7 50.9885
R96 VTAIL.n13 VTAIL.n12 49.1012
R97 VTAIL.n9 VTAIL.n8 49.1012
R98 VTAIL.n1 VTAIL.n0 49.1009
R99 VTAIL.n5 VTAIL.n4 49.1009
R100 VTAIL.n15 VTAIL.n14 23.4876
R101 VTAIL.n7 VTAIL.n6 23.4876
R102 VTAIL.n9 VTAIL.n7 2.07809
R103 VTAIL.n10 VTAIL.n9 2.07809
R104 VTAIL.n13 VTAIL.n11 2.07809
R105 VTAIL.n14 VTAIL.n13 2.07809
R106 VTAIL.n6 VTAIL.n5 2.07809
R107 VTAIL.n5 VTAIL.n3 2.07809
R108 VTAIL.n2 VTAIL.n1 2.07809
R109 VTAIL VTAIL.n15 2.0199
R110 VTAIL.n0 VTAIL.t13 1.88801
R111 VTAIL.n0 VTAIL.t10 1.88801
R112 VTAIL.n4 VTAIL.t5 1.88801
R113 VTAIL.n4 VTAIL.t0 1.88801
R114 VTAIL.n12 VTAIL.t4 1.88801
R115 VTAIL.n12 VTAIL.t6 1.88801
R116 VTAIL.n8 VTAIL.t12 1.88801
R117 VTAIL.n8 VTAIL.t15 1.88801
R118 VTAIL.n11 VTAIL.n10 0.470328
R119 VTAIL.n3 VTAIL.n2 0.470328
R120 VTAIL VTAIL.n1 0.0586897
R121 B.n777 B.n776 585
R122 B.n291 B.n123 585
R123 B.n290 B.n289 585
R124 B.n288 B.n287 585
R125 B.n286 B.n285 585
R126 B.n284 B.n283 585
R127 B.n282 B.n281 585
R128 B.n280 B.n279 585
R129 B.n278 B.n277 585
R130 B.n276 B.n275 585
R131 B.n274 B.n273 585
R132 B.n272 B.n271 585
R133 B.n270 B.n269 585
R134 B.n268 B.n267 585
R135 B.n266 B.n265 585
R136 B.n264 B.n263 585
R137 B.n262 B.n261 585
R138 B.n260 B.n259 585
R139 B.n258 B.n257 585
R140 B.n256 B.n255 585
R141 B.n254 B.n253 585
R142 B.n252 B.n251 585
R143 B.n250 B.n249 585
R144 B.n248 B.n247 585
R145 B.n246 B.n245 585
R146 B.n244 B.n243 585
R147 B.n242 B.n241 585
R148 B.n240 B.n239 585
R149 B.n238 B.n237 585
R150 B.n236 B.n235 585
R151 B.n234 B.n233 585
R152 B.n232 B.n231 585
R153 B.n230 B.n229 585
R154 B.n228 B.n227 585
R155 B.n226 B.n225 585
R156 B.n224 B.n223 585
R157 B.n222 B.n221 585
R158 B.n219 B.n218 585
R159 B.n217 B.n216 585
R160 B.n215 B.n214 585
R161 B.n213 B.n212 585
R162 B.n211 B.n210 585
R163 B.n209 B.n208 585
R164 B.n207 B.n206 585
R165 B.n205 B.n204 585
R166 B.n203 B.n202 585
R167 B.n201 B.n200 585
R168 B.n198 B.n197 585
R169 B.n196 B.n195 585
R170 B.n194 B.n193 585
R171 B.n192 B.n191 585
R172 B.n190 B.n189 585
R173 B.n188 B.n187 585
R174 B.n186 B.n185 585
R175 B.n184 B.n183 585
R176 B.n182 B.n181 585
R177 B.n180 B.n179 585
R178 B.n178 B.n177 585
R179 B.n176 B.n175 585
R180 B.n174 B.n173 585
R181 B.n172 B.n171 585
R182 B.n170 B.n169 585
R183 B.n168 B.n167 585
R184 B.n166 B.n165 585
R185 B.n164 B.n163 585
R186 B.n162 B.n161 585
R187 B.n160 B.n159 585
R188 B.n158 B.n157 585
R189 B.n156 B.n155 585
R190 B.n154 B.n153 585
R191 B.n152 B.n151 585
R192 B.n150 B.n149 585
R193 B.n148 B.n147 585
R194 B.n146 B.n145 585
R195 B.n144 B.n143 585
R196 B.n142 B.n141 585
R197 B.n140 B.n139 585
R198 B.n138 B.n137 585
R199 B.n136 B.n135 585
R200 B.n134 B.n133 585
R201 B.n132 B.n131 585
R202 B.n130 B.n129 585
R203 B.n82 B.n81 585
R204 B.n782 B.n781 585
R205 B.n775 B.n124 585
R206 B.n124 B.n79 585
R207 B.n774 B.n78 585
R208 B.n786 B.n78 585
R209 B.n773 B.n77 585
R210 B.n787 B.n77 585
R211 B.n772 B.n76 585
R212 B.n788 B.n76 585
R213 B.n771 B.n770 585
R214 B.n770 B.n72 585
R215 B.n769 B.n71 585
R216 B.n794 B.n71 585
R217 B.n768 B.n70 585
R218 B.n795 B.n70 585
R219 B.n767 B.n69 585
R220 B.n796 B.n69 585
R221 B.n766 B.n765 585
R222 B.n765 B.n65 585
R223 B.n764 B.n64 585
R224 B.n802 B.n64 585
R225 B.n763 B.n63 585
R226 B.n803 B.n63 585
R227 B.n762 B.n62 585
R228 B.n804 B.n62 585
R229 B.n761 B.n760 585
R230 B.n760 B.n58 585
R231 B.n759 B.n57 585
R232 B.n810 B.n57 585
R233 B.n758 B.n56 585
R234 B.n811 B.n56 585
R235 B.n757 B.n55 585
R236 B.n812 B.n55 585
R237 B.n756 B.n755 585
R238 B.n755 B.n51 585
R239 B.n754 B.n50 585
R240 B.n818 B.n50 585
R241 B.n753 B.n49 585
R242 B.n819 B.n49 585
R243 B.n752 B.n48 585
R244 B.n820 B.n48 585
R245 B.n751 B.n750 585
R246 B.n750 B.n44 585
R247 B.n749 B.n43 585
R248 B.n826 B.n43 585
R249 B.n748 B.n42 585
R250 B.n827 B.n42 585
R251 B.n747 B.n41 585
R252 B.n828 B.n41 585
R253 B.n746 B.n745 585
R254 B.n745 B.n40 585
R255 B.n744 B.n36 585
R256 B.n834 B.n36 585
R257 B.n743 B.n35 585
R258 B.n835 B.n35 585
R259 B.n742 B.n34 585
R260 B.n836 B.n34 585
R261 B.n741 B.n740 585
R262 B.n740 B.n30 585
R263 B.n739 B.n29 585
R264 B.n842 B.n29 585
R265 B.n738 B.n28 585
R266 B.n843 B.n28 585
R267 B.n737 B.n27 585
R268 B.n844 B.n27 585
R269 B.n736 B.n735 585
R270 B.n735 B.n23 585
R271 B.n734 B.n22 585
R272 B.n850 B.n22 585
R273 B.n733 B.n21 585
R274 B.n851 B.n21 585
R275 B.n732 B.n20 585
R276 B.n852 B.n20 585
R277 B.n731 B.n730 585
R278 B.n730 B.n16 585
R279 B.n729 B.n15 585
R280 B.n858 B.n15 585
R281 B.n728 B.n14 585
R282 B.n859 B.n14 585
R283 B.n727 B.n13 585
R284 B.n860 B.n13 585
R285 B.n726 B.n725 585
R286 B.n725 B.n12 585
R287 B.n724 B.n723 585
R288 B.n724 B.n8 585
R289 B.n722 B.n7 585
R290 B.n867 B.n7 585
R291 B.n721 B.n6 585
R292 B.n868 B.n6 585
R293 B.n720 B.n5 585
R294 B.n869 B.n5 585
R295 B.n719 B.n718 585
R296 B.n718 B.n4 585
R297 B.n717 B.n292 585
R298 B.n717 B.n716 585
R299 B.n707 B.n293 585
R300 B.n294 B.n293 585
R301 B.n709 B.n708 585
R302 B.n710 B.n709 585
R303 B.n706 B.n298 585
R304 B.n302 B.n298 585
R305 B.n705 B.n704 585
R306 B.n704 B.n703 585
R307 B.n300 B.n299 585
R308 B.n301 B.n300 585
R309 B.n696 B.n695 585
R310 B.n697 B.n696 585
R311 B.n694 B.n307 585
R312 B.n307 B.n306 585
R313 B.n693 B.n692 585
R314 B.n692 B.n691 585
R315 B.n309 B.n308 585
R316 B.n310 B.n309 585
R317 B.n684 B.n683 585
R318 B.n685 B.n684 585
R319 B.n682 B.n315 585
R320 B.n315 B.n314 585
R321 B.n681 B.n680 585
R322 B.n680 B.n679 585
R323 B.n317 B.n316 585
R324 B.n318 B.n317 585
R325 B.n672 B.n671 585
R326 B.n673 B.n672 585
R327 B.n670 B.n323 585
R328 B.n323 B.n322 585
R329 B.n669 B.n668 585
R330 B.n668 B.n667 585
R331 B.n325 B.n324 585
R332 B.n660 B.n325 585
R333 B.n659 B.n658 585
R334 B.n661 B.n659 585
R335 B.n657 B.n330 585
R336 B.n330 B.n329 585
R337 B.n656 B.n655 585
R338 B.n655 B.n654 585
R339 B.n332 B.n331 585
R340 B.n333 B.n332 585
R341 B.n647 B.n646 585
R342 B.n648 B.n647 585
R343 B.n645 B.n338 585
R344 B.n338 B.n337 585
R345 B.n644 B.n643 585
R346 B.n643 B.n642 585
R347 B.n340 B.n339 585
R348 B.n341 B.n340 585
R349 B.n635 B.n634 585
R350 B.n636 B.n635 585
R351 B.n633 B.n346 585
R352 B.n346 B.n345 585
R353 B.n632 B.n631 585
R354 B.n631 B.n630 585
R355 B.n348 B.n347 585
R356 B.n349 B.n348 585
R357 B.n623 B.n622 585
R358 B.n624 B.n623 585
R359 B.n621 B.n354 585
R360 B.n354 B.n353 585
R361 B.n620 B.n619 585
R362 B.n619 B.n618 585
R363 B.n356 B.n355 585
R364 B.n357 B.n356 585
R365 B.n611 B.n610 585
R366 B.n612 B.n611 585
R367 B.n609 B.n361 585
R368 B.n365 B.n361 585
R369 B.n608 B.n607 585
R370 B.n607 B.n606 585
R371 B.n363 B.n362 585
R372 B.n364 B.n363 585
R373 B.n599 B.n598 585
R374 B.n600 B.n599 585
R375 B.n597 B.n370 585
R376 B.n370 B.n369 585
R377 B.n596 B.n595 585
R378 B.n595 B.n594 585
R379 B.n372 B.n371 585
R380 B.n373 B.n372 585
R381 B.n590 B.n589 585
R382 B.n376 B.n375 585
R383 B.n586 B.n585 585
R384 B.n587 B.n586 585
R385 B.n584 B.n418 585
R386 B.n583 B.n582 585
R387 B.n581 B.n580 585
R388 B.n579 B.n578 585
R389 B.n577 B.n576 585
R390 B.n575 B.n574 585
R391 B.n573 B.n572 585
R392 B.n571 B.n570 585
R393 B.n569 B.n568 585
R394 B.n567 B.n566 585
R395 B.n565 B.n564 585
R396 B.n563 B.n562 585
R397 B.n561 B.n560 585
R398 B.n559 B.n558 585
R399 B.n557 B.n556 585
R400 B.n555 B.n554 585
R401 B.n553 B.n552 585
R402 B.n551 B.n550 585
R403 B.n549 B.n548 585
R404 B.n547 B.n546 585
R405 B.n545 B.n544 585
R406 B.n543 B.n542 585
R407 B.n541 B.n540 585
R408 B.n539 B.n538 585
R409 B.n537 B.n536 585
R410 B.n535 B.n534 585
R411 B.n533 B.n532 585
R412 B.n531 B.n530 585
R413 B.n529 B.n528 585
R414 B.n527 B.n526 585
R415 B.n525 B.n524 585
R416 B.n523 B.n522 585
R417 B.n521 B.n520 585
R418 B.n519 B.n518 585
R419 B.n517 B.n516 585
R420 B.n515 B.n514 585
R421 B.n513 B.n512 585
R422 B.n511 B.n510 585
R423 B.n509 B.n508 585
R424 B.n507 B.n506 585
R425 B.n505 B.n504 585
R426 B.n503 B.n502 585
R427 B.n501 B.n500 585
R428 B.n499 B.n498 585
R429 B.n497 B.n496 585
R430 B.n495 B.n494 585
R431 B.n493 B.n492 585
R432 B.n491 B.n490 585
R433 B.n489 B.n488 585
R434 B.n487 B.n486 585
R435 B.n485 B.n484 585
R436 B.n483 B.n482 585
R437 B.n481 B.n480 585
R438 B.n479 B.n478 585
R439 B.n477 B.n476 585
R440 B.n475 B.n474 585
R441 B.n473 B.n472 585
R442 B.n471 B.n470 585
R443 B.n469 B.n468 585
R444 B.n467 B.n466 585
R445 B.n465 B.n464 585
R446 B.n463 B.n462 585
R447 B.n461 B.n460 585
R448 B.n459 B.n458 585
R449 B.n457 B.n456 585
R450 B.n455 B.n454 585
R451 B.n453 B.n452 585
R452 B.n451 B.n450 585
R453 B.n449 B.n448 585
R454 B.n447 B.n446 585
R455 B.n445 B.n444 585
R456 B.n443 B.n442 585
R457 B.n441 B.n440 585
R458 B.n439 B.n438 585
R459 B.n437 B.n436 585
R460 B.n435 B.n434 585
R461 B.n433 B.n432 585
R462 B.n431 B.n430 585
R463 B.n429 B.n428 585
R464 B.n427 B.n426 585
R465 B.n425 B.n417 585
R466 B.n587 B.n417 585
R467 B.n591 B.n374 585
R468 B.n374 B.n373 585
R469 B.n593 B.n592 585
R470 B.n594 B.n593 585
R471 B.n368 B.n367 585
R472 B.n369 B.n368 585
R473 B.n602 B.n601 585
R474 B.n601 B.n600 585
R475 B.n603 B.n366 585
R476 B.n366 B.n364 585
R477 B.n605 B.n604 585
R478 B.n606 B.n605 585
R479 B.n360 B.n359 585
R480 B.n365 B.n360 585
R481 B.n614 B.n613 585
R482 B.n613 B.n612 585
R483 B.n615 B.n358 585
R484 B.n358 B.n357 585
R485 B.n617 B.n616 585
R486 B.n618 B.n617 585
R487 B.n352 B.n351 585
R488 B.n353 B.n352 585
R489 B.n626 B.n625 585
R490 B.n625 B.n624 585
R491 B.n627 B.n350 585
R492 B.n350 B.n349 585
R493 B.n629 B.n628 585
R494 B.n630 B.n629 585
R495 B.n344 B.n343 585
R496 B.n345 B.n344 585
R497 B.n638 B.n637 585
R498 B.n637 B.n636 585
R499 B.n639 B.n342 585
R500 B.n342 B.n341 585
R501 B.n641 B.n640 585
R502 B.n642 B.n641 585
R503 B.n336 B.n335 585
R504 B.n337 B.n336 585
R505 B.n650 B.n649 585
R506 B.n649 B.n648 585
R507 B.n651 B.n334 585
R508 B.n334 B.n333 585
R509 B.n653 B.n652 585
R510 B.n654 B.n653 585
R511 B.n328 B.n327 585
R512 B.n329 B.n328 585
R513 B.n663 B.n662 585
R514 B.n662 B.n661 585
R515 B.n664 B.n326 585
R516 B.n660 B.n326 585
R517 B.n666 B.n665 585
R518 B.n667 B.n666 585
R519 B.n321 B.n320 585
R520 B.n322 B.n321 585
R521 B.n675 B.n674 585
R522 B.n674 B.n673 585
R523 B.n676 B.n319 585
R524 B.n319 B.n318 585
R525 B.n678 B.n677 585
R526 B.n679 B.n678 585
R527 B.n313 B.n312 585
R528 B.n314 B.n313 585
R529 B.n687 B.n686 585
R530 B.n686 B.n685 585
R531 B.n688 B.n311 585
R532 B.n311 B.n310 585
R533 B.n690 B.n689 585
R534 B.n691 B.n690 585
R535 B.n305 B.n304 585
R536 B.n306 B.n305 585
R537 B.n699 B.n698 585
R538 B.n698 B.n697 585
R539 B.n700 B.n303 585
R540 B.n303 B.n301 585
R541 B.n702 B.n701 585
R542 B.n703 B.n702 585
R543 B.n297 B.n296 585
R544 B.n302 B.n297 585
R545 B.n712 B.n711 585
R546 B.n711 B.n710 585
R547 B.n713 B.n295 585
R548 B.n295 B.n294 585
R549 B.n715 B.n714 585
R550 B.n716 B.n715 585
R551 B.n3 B.n0 585
R552 B.n4 B.n3 585
R553 B.n866 B.n1 585
R554 B.n867 B.n866 585
R555 B.n865 B.n864 585
R556 B.n865 B.n8 585
R557 B.n863 B.n9 585
R558 B.n12 B.n9 585
R559 B.n862 B.n861 585
R560 B.n861 B.n860 585
R561 B.n11 B.n10 585
R562 B.n859 B.n11 585
R563 B.n857 B.n856 585
R564 B.n858 B.n857 585
R565 B.n855 B.n17 585
R566 B.n17 B.n16 585
R567 B.n854 B.n853 585
R568 B.n853 B.n852 585
R569 B.n19 B.n18 585
R570 B.n851 B.n19 585
R571 B.n849 B.n848 585
R572 B.n850 B.n849 585
R573 B.n847 B.n24 585
R574 B.n24 B.n23 585
R575 B.n846 B.n845 585
R576 B.n845 B.n844 585
R577 B.n26 B.n25 585
R578 B.n843 B.n26 585
R579 B.n841 B.n840 585
R580 B.n842 B.n841 585
R581 B.n839 B.n31 585
R582 B.n31 B.n30 585
R583 B.n838 B.n837 585
R584 B.n837 B.n836 585
R585 B.n33 B.n32 585
R586 B.n835 B.n33 585
R587 B.n833 B.n832 585
R588 B.n834 B.n833 585
R589 B.n831 B.n37 585
R590 B.n40 B.n37 585
R591 B.n830 B.n829 585
R592 B.n829 B.n828 585
R593 B.n39 B.n38 585
R594 B.n827 B.n39 585
R595 B.n825 B.n824 585
R596 B.n826 B.n825 585
R597 B.n823 B.n45 585
R598 B.n45 B.n44 585
R599 B.n822 B.n821 585
R600 B.n821 B.n820 585
R601 B.n47 B.n46 585
R602 B.n819 B.n47 585
R603 B.n817 B.n816 585
R604 B.n818 B.n817 585
R605 B.n815 B.n52 585
R606 B.n52 B.n51 585
R607 B.n814 B.n813 585
R608 B.n813 B.n812 585
R609 B.n54 B.n53 585
R610 B.n811 B.n54 585
R611 B.n809 B.n808 585
R612 B.n810 B.n809 585
R613 B.n807 B.n59 585
R614 B.n59 B.n58 585
R615 B.n806 B.n805 585
R616 B.n805 B.n804 585
R617 B.n61 B.n60 585
R618 B.n803 B.n61 585
R619 B.n801 B.n800 585
R620 B.n802 B.n801 585
R621 B.n799 B.n66 585
R622 B.n66 B.n65 585
R623 B.n798 B.n797 585
R624 B.n797 B.n796 585
R625 B.n68 B.n67 585
R626 B.n795 B.n68 585
R627 B.n793 B.n792 585
R628 B.n794 B.n793 585
R629 B.n791 B.n73 585
R630 B.n73 B.n72 585
R631 B.n790 B.n789 585
R632 B.n789 B.n788 585
R633 B.n75 B.n74 585
R634 B.n787 B.n75 585
R635 B.n785 B.n784 585
R636 B.n786 B.n785 585
R637 B.n783 B.n80 585
R638 B.n80 B.n79 585
R639 B.n870 B.n869 585
R640 B.n868 B.n2 585
R641 B.n781 B.n80 502.111
R642 B.n777 B.n124 502.111
R643 B.n417 B.n372 502.111
R644 B.n589 B.n374 502.111
R645 B.n127 B.t7 328.642
R646 B.n125 B.t11 328.642
R647 B.n422 B.t18 328.642
R648 B.n419 B.t14 328.642
R649 B.n779 B.n778 256.663
R650 B.n779 B.n122 256.663
R651 B.n779 B.n121 256.663
R652 B.n779 B.n120 256.663
R653 B.n779 B.n119 256.663
R654 B.n779 B.n118 256.663
R655 B.n779 B.n117 256.663
R656 B.n779 B.n116 256.663
R657 B.n779 B.n115 256.663
R658 B.n779 B.n114 256.663
R659 B.n779 B.n113 256.663
R660 B.n779 B.n112 256.663
R661 B.n779 B.n111 256.663
R662 B.n779 B.n110 256.663
R663 B.n779 B.n109 256.663
R664 B.n779 B.n108 256.663
R665 B.n779 B.n107 256.663
R666 B.n779 B.n106 256.663
R667 B.n779 B.n105 256.663
R668 B.n779 B.n104 256.663
R669 B.n779 B.n103 256.663
R670 B.n779 B.n102 256.663
R671 B.n779 B.n101 256.663
R672 B.n779 B.n100 256.663
R673 B.n779 B.n99 256.663
R674 B.n779 B.n98 256.663
R675 B.n779 B.n97 256.663
R676 B.n779 B.n96 256.663
R677 B.n779 B.n95 256.663
R678 B.n779 B.n94 256.663
R679 B.n779 B.n93 256.663
R680 B.n779 B.n92 256.663
R681 B.n779 B.n91 256.663
R682 B.n779 B.n90 256.663
R683 B.n779 B.n89 256.663
R684 B.n779 B.n88 256.663
R685 B.n779 B.n87 256.663
R686 B.n779 B.n86 256.663
R687 B.n779 B.n85 256.663
R688 B.n779 B.n84 256.663
R689 B.n779 B.n83 256.663
R690 B.n780 B.n779 256.663
R691 B.n588 B.n587 256.663
R692 B.n587 B.n377 256.663
R693 B.n587 B.n378 256.663
R694 B.n587 B.n379 256.663
R695 B.n587 B.n380 256.663
R696 B.n587 B.n381 256.663
R697 B.n587 B.n382 256.663
R698 B.n587 B.n383 256.663
R699 B.n587 B.n384 256.663
R700 B.n587 B.n385 256.663
R701 B.n587 B.n386 256.663
R702 B.n587 B.n387 256.663
R703 B.n587 B.n388 256.663
R704 B.n587 B.n389 256.663
R705 B.n587 B.n390 256.663
R706 B.n587 B.n391 256.663
R707 B.n587 B.n392 256.663
R708 B.n587 B.n393 256.663
R709 B.n587 B.n394 256.663
R710 B.n587 B.n395 256.663
R711 B.n587 B.n396 256.663
R712 B.n587 B.n397 256.663
R713 B.n587 B.n398 256.663
R714 B.n587 B.n399 256.663
R715 B.n587 B.n400 256.663
R716 B.n587 B.n401 256.663
R717 B.n587 B.n402 256.663
R718 B.n587 B.n403 256.663
R719 B.n587 B.n404 256.663
R720 B.n587 B.n405 256.663
R721 B.n587 B.n406 256.663
R722 B.n587 B.n407 256.663
R723 B.n587 B.n408 256.663
R724 B.n587 B.n409 256.663
R725 B.n587 B.n410 256.663
R726 B.n587 B.n411 256.663
R727 B.n587 B.n412 256.663
R728 B.n587 B.n413 256.663
R729 B.n587 B.n414 256.663
R730 B.n587 B.n415 256.663
R731 B.n587 B.n416 256.663
R732 B.n872 B.n871 256.663
R733 B.n129 B.n82 163.367
R734 B.n133 B.n132 163.367
R735 B.n137 B.n136 163.367
R736 B.n141 B.n140 163.367
R737 B.n145 B.n144 163.367
R738 B.n149 B.n148 163.367
R739 B.n153 B.n152 163.367
R740 B.n157 B.n156 163.367
R741 B.n161 B.n160 163.367
R742 B.n165 B.n164 163.367
R743 B.n169 B.n168 163.367
R744 B.n173 B.n172 163.367
R745 B.n177 B.n176 163.367
R746 B.n181 B.n180 163.367
R747 B.n185 B.n184 163.367
R748 B.n189 B.n188 163.367
R749 B.n193 B.n192 163.367
R750 B.n197 B.n196 163.367
R751 B.n202 B.n201 163.367
R752 B.n206 B.n205 163.367
R753 B.n210 B.n209 163.367
R754 B.n214 B.n213 163.367
R755 B.n218 B.n217 163.367
R756 B.n223 B.n222 163.367
R757 B.n227 B.n226 163.367
R758 B.n231 B.n230 163.367
R759 B.n235 B.n234 163.367
R760 B.n239 B.n238 163.367
R761 B.n243 B.n242 163.367
R762 B.n247 B.n246 163.367
R763 B.n251 B.n250 163.367
R764 B.n255 B.n254 163.367
R765 B.n259 B.n258 163.367
R766 B.n263 B.n262 163.367
R767 B.n267 B.n266 163.367
R768 B.n271 B.n270 163.367
R769 B.n275 B.n274 163.367
R770 B.n279 B.n278 163.367
R771 B.n283 B.n282 163.367
R772 B.n287 B.n286 163.367
R773 B.n289 B.n123 163.367
R774 B.n595 B.n372 163.367
R775 B.n595 B.n370 163.367
R776 B.n599 B.n370 163.367
R777 B.n599 B.n363 163.367
R778 B.n607 B.n363 163.367
R779 B.n607 B.n361 163.367
R780 B.n611 B.n361 163.367
R781 B.n611 B.n356 163.367
R782 B.n619 B.n356 163.367
R783 B.n619 B.n354 163.367
R784 B.n623 B.n354 163.367
R785 B.n623 B.n348 163.367
R786 B.n631 B.n348 163.367
R787 B.n631 B.n346 163.367
R788 B.n635 B.n346 163.367
R789 B.n635 B.n340 163.367
R790 B.n643 B.n340 163.367
R791 B.n643 B.n338 163.367
R792 B.n647 B.n338 163.367
R793 B.n647 B.n332 163.367
R794 B.n655 B.n332 163.367
R795 B.n655 B.n330 163.367
R796 B.n659 B.n330 163.367
R797 B.n659 B.n325 163.367
R798 B.n668 B.n325 163.367
R799 B.n668 B.n323 163.367
R800 B.n672 B.n323 163.367
R801 B.n672 B.n317 163.367
R802 B.n680 B.n317 163.367
R803 B.n680 B.n315 163.367
R804 B.n684 B.n315 163.367
R805 B.n684 B.n309 163.367
R806 B.n692 B.n309 163.367
R807 B.n692 B.n307 163.367
R808 B.n696 B.n307 163.367
R809 B.n696 B.n300 163.367
R810 B.n704 B.n300 163.367
R811 B.n704 B.n298 163.367
R812 B.n709 B.n298 163.367
R813 B.n709 B.n293 163.367
R814 B.n717 B.n293 163.367
R815 B.n718 B.n717 163.367
R816 B.n718 B.n5 163.367
R817 B.n6 B.n5 163.367
R818 B.n7 B.n6 163.367
R819 B.n724 B.n7 163.367
R820 B.n725 B.n724 163.367
R821 B.n725 B.n13 163.367
R822 B.n14 B.n13 163.367
R823 B.n15 B.n14 163.367
R824 B.n730 B.n15 163.367
R825 B.n730 B.n20 163.367
R826 B.n21 B.n20 163.367
R827 B.n22 B.n21 163.367
R828 B.n735 B.n22 163.367
R829 B.n735 B.n27 163.367
R830 B.n28 B.n27 163.367
R831 B.n29 B.n28 163.367
R832 B.n740 B.n29 163.367
R833 B.n740 B.n34 163.367
R834 B.n35 B.n34 163.367
R835 B.n36 B.n35 163.367
R836 B.n745 B.n36 163.367
R837 B.n745 B.n41 163.367
R838 B.n42 B.n41 163.367
R839 B.n43 B.n42 163.367
R840 B.n750 B.n43 163.367
R841 B.n750 B.n48 163.367
R842 B.n49 B.n48 163.367
R843 B.n50 B.n49 163.367
R844 B.n755 B.n50 163.367
R845 B.n755 B.n55 163.367
R846 B.n56 B.n55 163.367
R847 B.n57 B.n56 163.367
R848 B.n760 B.n57 163.367
R849 B.n760 B.n62 163.367
R850 B.n63 B.n62 163.367
R851 B.n64 B.n63 163.367
R852 B.n765 B.n64 163.367
R853 B.n765 B.n69 163.367
R854 B.n70 B.n69 163.367
R855 B.n71 B.n70 163.367
R856 B.n770 B.n71 163.367
R857 B.n770 B.n76 163.367
R858 B.n77 B.n76 163.367
R859 B.n78 B.n77 163.367
R860 B.n124 B.n78 163.367
R861 B.n586 B.n376 163.367
R862 B.n586 B.n418 163.367
R863 B.n582 B.n581 163.367
R864 B.n578 B.n577 163.367
R865 B.n574 B.n573 163.367
R866 B.n570 B.n569 163.367
R867 B.n566 B.n565 163.367
R868 B.n562 B.n561 163.367
R869 B.n558 B.n557 163.367
R870 B.n554 B.n553 163.367
R871 B.n550 B.n549 163.367
R872 B.n546 B.n545 163.367
R873 B.n542 B.n541 163.367
R874 B.n538 B.n537 163.367
R875 B.n534 B.n533 163.367
R876 B.n530 B.n529 163.367
R877 B.n526 B.n525 163.367
R878 B.n522 B.n521 163.367
R879 B.n518 B.n517 163.367
R880 B.n514 B.n513 163.367
R881 B.n510 B.n509 163.367
R882 B.n506 B.n505 163.367
R883 B.n502 B.n501 163.367
R884 B.n498 B.n497 163.367
R885 B.n494 B.n493 163.367
R886 B.n490 B.n489 163.367
R887 B.n486 B.n485 163.367
R888 B.n482 B.n481 163.367
R889 B.n478 B.n477 163.367
R890 B.n474 B.n473 163.367
R891 B.n470 B.n469 163.367
R892 B.n466 B.n465 163.367
R893 B.n462 B.n461 163.367
R894 B.n458 B.n457 163.367
R895 B.n454 B.n453 163.367
R896 B.n450 B.n449 163.367
R897 B.n446 B.n445 163.367
R898 B.n442 B.n441 163.367
R899 B.n438 B.n437 163.367
R900 B.n434 B.n433 163.367
R901 B.n430 B.n429 163.367
R902 B.n426 B.n417 163.367
R903 B.n593 B.n374 163.367
R904 B.n593 B.n368 163.367
R905 B.n601 B.n368 163.367
R906 B.n601 B.n366 163.367
R907 B.n605 B.n366 163.367
R908 B.n605 B.n360 163.367
R909 B.n613 B.n360 163.367
R910 B.n613 B.n358 163.367
R911 B.n617 B.n358 163.367
R912 B.n617 B.n352 163.367
R913 B.n625 B.n352 163.367
R914 B.n625 B.n350 163.367
R915 B.n629 B.n350 163.367
R916 B.n629 B.n344 163.367
R917 B.n637 B.n344 163.367
R918 B.n637 B.n342 163.367
R919 B.n641 B.n342 163.367
R920 B.n641 B.n336 163.367
R921 B.n649 B.n336 163.367
R922 B.n649 B.n334 163.367
R923 B.n653 B.n334 163.367
R924 B.n653 B.n328 163.367
R925 B.n662 B.n328 163.367
R926 B.n662 B.n326 163.367
R927 B.n666 B.n326 163.367
R928 B.n666 B.n321 163.367
R929 B.n674 B.n321 163.367
R930 B.n674 B.n319 163.367
R931 B.n678 B.n319 163.367
R932 B.n678 B.n313 163.367
R933 B.n686 B.n313 163.367
R934 B.n686 B.n311 163.367
R935 B.n690 B.n311 163.367
R936 B.n690 B.n305 163.367
R937 B.n698 B.n305 163.367
R938 B.n698 B.n303 163.367
R939 B.n702 B.n303 163.367
R940 B.n702 B.n297 163.367
R941 B.n711 B.n297 163.367
R942 B.n711 B.n295 163.367
R943 B.n715 B.n295 163.367
R944 B.n715 B.n3 163.367
R945 B.n870 B.n3 163.367
R946 B.n866 B.n2 163.367
R947 B.n866 B.n865 163.367
R948 B.n865 B.n9 163.367
R949 B.n861 B.n9 163.367
R950 B.n861 B.n11 163.367
R951 B.n857 B.n11 163.367
R952 B.n857 B.n17 163.367
R953 B.n853 B.n17 163.367
R954 B.n853 B.n19 163.367
R955 B.n849 B.n19 163.367
R956 B.n849 B.n24 163.367
R957 B.n845 B.n24 163.367
R958 B.n845 B.n26 163.367
R959 B.n841 B.n26 163.367
R960 B.n841 B.n31 163.367
R961 B.n837 B.n31 163.367
R962 B.n837 B.n33 163.367
R963 B.n833 B.n33 163.367
R964 B.n833 B.n37 163.367
R965 B.n829 B.n37 163.367
R966 B.n829 B.n39 163.367
R967 B.n825 B.n39 163.367
R968 B.n825 B.n45 163.367
R969 B.n821 B.n45 163.367
R970 B.n821 B.n47 163.367
R971 B.n817 B.n47 163.367
R972 B.n817 B.n52 163.367
R973 B.n813 B.n52 163.367
R974 B.n813 B.n54 163.367
R975 B.n809 B.n54 163.367
R976 B.n809 B.n59 163.367
R977 B.n805 B.n59 163.367
R978 B.n805 B.n61 163.367
R979 B.n801 B.n61 163.367
R980 B.n801 B.n66 163.367
R981 B.n797 B.n66 163.367
R982 B.n797 B.n68 163.367
R983 B.n793 B.n68 163.367
R984 B.n793 B.n73 163.367
R985 B.n789 B.n73 163.367
R986 B.n789 B.n75 163.367
R987 B.n785 B.n75 163.367
R988 B.n785 B.n80 163.367
R989 B.n125 B.t12 120.388
R990 B.n422 B.t20 120.388
R991 B.n127 B.t9 120.376
R992 B.n419 B.t17 120.376
R993 B.n587 B.n373 88.6145
R994 B.n779 B.n79 88.6145
R995 B.n126 B.t13 73.6492
R996 B.n423 B.t19 73.6492
R997 B.n128 B.t10 73.6364
R998 B.n420 B.t16 73.6364
R999 B.n781 B.n780 71.676
R1000 B.n129 B.n83 71.676
R1001 B.n133 B.n84 71.676
R1002 B.n137 B.n85 71.676
R1003 B.n141 B.n86 71.676
R1004 B.n145 B.n87 71.676
R1005 B.n149 B.n88 71.676
R1006 B.n153 B.n89 71.676
R1007 B.n157 B.n90 71.676
R1008 B.n161 B.n91 71.676
R1009 B.n165 B.n92 71.676
R1010 B.n169 B.n93 71.676
R1011 B.n173 B.n94 71.676
R1012 B.n177 B.n95 71.676
R1013 B.n181 B.n96 71.676
R1014 B.n185 B.n97 71.676
R1015 B.n189 B.n98 71.676
R1016 B.n193 B.n99 71.676
R1017 B.n197 B.n100 71.676
R1018 B.n202 B.n101 71.676
R1019 B.n206 B.n102 71.676
R1020 B.n210 B.n103 71.676
R1021 B.n214 B.n104 71.676
R1022 B.n218 B.n105 71.676
R1023 B.n223 B.n106 71.676
R1024 B.n227 B.n107 71.676
R1025 B.n231 B.n108 71.676
R1026 B.n235 B.n109 71.676
R1027 B.n239 B.n110 71.676
R1028 B.n243 B.n111 71.676
R1029 B.n247 B.n112 71.676
R1030 B.n251 B.n113 71.676
R1031 B.n255 B.n114 71.676
R1032 B.n259 B.n115 71.676
R1033 B.n263 B.n116 71.676
R1034 B.n267 B.n117 71.676
R1035 B.n271 B.n118 71.676
R1036 B.n275 B.n119 71.676
R1037 B.n279 B.n120 71.676
R1038 B.n283 B.n121 71.676
R1039 B.n287 B.n122 71.676
R1040 B.n778 B.n123 71.676
R1041 B.n778 B.n777 71.676
R1042 B.n289 B.n122 71.676
R1043 B.n286 B.n121 71.676
R1044 B.n282 B.n120 71.676
R1045 B.n278 B.n119 71.676
R1046 B.n274 B.n118 71.676
R1047 B.n270 B.n117 71.676
R1048 B.n266 B.n116 71.676
R1049 B.n262 B.n115 71.676
R1050 B.n258 B.n114 71.676
R1051 B.n254 B.n113 71.676
R1052 B.n250 B.n112 71.676
R1053 B.n246 B.n111 71.676
R1054 B.n242 B.n110 71.676
R1055 B.n238 B.n109 71.676
R1056 B.n234 B.n108 71.676
R1057 B.n230 B.n107 71.676
R1058 B.n226 B.n106 71.676
R1059 B.n222 B.n105 71.676
R1060 B.n217 B.n104 71.676
R1061 B.n213 B.n103 71.676
R1062 B.n209 B.n102 71.676
R1063 B.n205 B.n101 71.676
R1064 B.n201 B.n100 71.676
R1065 B.n196 B.n99 71.676
R1066 B.n192 B.n98 71.676
R1067 B.n188 B.n97 71.676
R1068 B.n184 B.n96 71.676
R1069 B.n180 B.n95 71.676
R1070 B.n176 B.n94 71.676
R1071 B.n172 B.n93 71.676
R1072 B.n168 B.n92 71.676
R1073 B.n164 B.n91 71.676
R1074 B.n160 B.n90 71.676
R1075 B.n156 B.n89 71.676
R1076 B.n152 B.n88 71.676
R1077 B.n148 B.n87 71.676
R1078 B.n144 B.n86 71.676
R1079 B.n140 B.n85 71.676
R1080 B.n136 B.n84 71.676
R1081 B.n132 B.n83 71.676
R1082 B.n780 B.n82 71.676
R1083 B.n589 B.n588 71.676
R1084 B.n418 B.n377 71.676
R1085 B.n581 B.n378 71.676
R1086 B.n577 B.n379 71.676
R1087 B.n573 B.n380 71.676
R1088 B.n569 B.n381 71.676
R1089 B.n565 B.n382 71.676
R1090 B.n561 B.n383 71.676
R1091 B.n557 B.n384 71.676
R1092 B.n553 B.n385 71.676
R1093 B.n549 B.n386 71.676
R1094 B.n545 B.n387 71.676
R1095 B.n541 B.n388 71.676
R1096 B.n537 B.n389 71.676
R1097 B.n533 B.n390 71.676
R1098 B.n529 B.n391 71.676
R1099 B.n525 B.n392 71.676
R1100 B.n521 B.n393 71.676
R1101 B.n517 B.n394 71.676
R1102 B.n513 B.n395 71.676
R1103 B.n509 B.n396 71.676
R1104 B.n505 B.n397 71.676
R1105 B.n501 B.n398 71.676
R1106 B.n497 B.n399 71.676
R1107 B.n493 B.n400 71.676
R1108 B.n489 B.n401 71.676
R1109 B.n485 B.n402 71.676
R1110 B.n481 B.n403 71.676
R1111 B.n477 B.n404 71.676
R1112 B.n473 B.n405 71.676
R1113 B.n469 B.n406 71.676
R1114 B.n465 B.n407 71.676
R1115 B.n461 B.n408 71.676
R1116 B.n457 B.n409 71.676
R1117 B.n453 B.n410 71.676
R1118 B.n449 B.n411 71.676
R1119 B.n445 B.n412 71.676
R1120 B.n441 B.n413 71.676
R1121 B.n437 B.n414 71.676
R1122 B.n433 B.n415 71.676
R1123 B.n429 B.n416 71.676
R1124 B.n588 B.n376 71.676
R1125 B.n582 B.n377 71.676
R1126 B.n578 B.n378 71.676
R1127 B.n574 B.n379 71.676
R1128 B.n570 B.n380 71.676
R1129 B.n566 B.n381 71.676
R1130 B.n562 B.n382 71.676
R1131 B.n558 B.n383 71.676
R1132 B.n554 B.n384 71.676
R1133 B.n550 B.n385 71.676
R1134 B.n546 B.n386 71.676
R1135 B.n542 B.n387 71.676
R1136 B.n538 B.n388 71.676
R1137 B.n534 B.n389 71.676
R1138 B.n530 B.n390 71.676
R1139 B.n526 B.n391 71.676
R1140 B.n522 B.n392 71.676
R1141 B.n518 B.n393 71.676
R1142 B.n514 B.n394 71.676
R1143 B.n510 B.n395 71.676
R1144 B.n506 B.n396 71.676
R1145 B.n502 B.n397 71.676
R1146 B.n498 B.n398 71.676
R1147 B.n494 B.n399 71.676
R1148 B.n490 B.n400 71.676
R1149 B.n486 B.n401 71.676
R1150 B.n482 B.n402 71.676
R1151 B.n478 B.n403 71.676
R1152 B.n474 B.n404 71.676
R1153 B.n470 B.n405 71.676
R1154 B.n466 B.n406 71.676
R1155 B.n462 B.n407 71.676
R1156 B.n458 B.n408 71.676
R1157 B.n454 B.n409 71.676
R1158 B.n450 B.n410 71.676
R1159 B.n446 B.n411 71.676
R1160 B.n442 B.n412 71.676
R1161 B.n438 B.n413 71.676
R1162 B.n434 B.n414 71.676
R1163 B.n430 B.n415 71.676
R1164 B.n426 B.n416 71.676
R1165 B.n871 B.n870 71.676
R1166 B.n871 B.n2 71.676
R1167 B.n199 B.n128 59.5399
R1168 B.n220 B.n126 59.5399
R1169 B.n424 B.n423 59.5399
R1170 B.n421 B.n420 59.5399
R1171 B.n594 B.n373 47.4474
R1172 B.n594 B.n369 47.4474
R1173 B.n600 B.n369 47.4474
R1174 B.n600 B.n364 47.4474
R1175 B.n606 B.n364 47.4474
R1176 B.n606 B.n365 47.4474
R1177 B.n612 B.n357 47.4474
R1178 B.n618 B.n357 47.4474
R1179 B.n618 B.n353 47.4474
R1180 B.n624 B.n353 47.4474
R1181 B.n624 B.n349 47.4474
R1182 B.n630 B.n349 47.4474
R1183 B.n630 B.n345 47.4474
R1184 B.n636 B.n345 47.4474
R1185 B.n636 B.n341 47.4474
R1186 B.n642 B.n341 47.4474
R1187 B.n648 B.n337 47.4474
R1188 B.n648 B.n333 47.4474
R1189 B.n654 B.n333 47.4474
R1190 B.n654 B.n329 47.4474
R1191 B.n661 B.n329 47.4474
R1192 B.n661 B.n660 47.4474
R1193 B.n667 B.n322 47.4474
R1194 B.n673 B.n322 47.4474
R1195 B.n673 B.n318 47.4474
R1196 B.n679 B.n318 47.4474
R1197 B.n679 B.n314 47.4474
R1198 B.n685 B.n314 47.4474
R1199 B.n691 B.n310 47.4474
R1200 B.n691 B.n306 47.4474
R1201 B.n697 B.n306 47.4474
R1202 B.n697 B.n301 47.4474
R1203 B.n703 B.n301 47.4474
R1204 B.n703 B.n302 47.4474
R1205 B.n710 B.n294 47.4474
R1206 B.n716 B.n294 47.4474
R1207 B.n716 B.n4 47.4474
R1208 B.n869 B.n4 47.4474
R1209 B.n869 B.n868 47.4474
R1210 B.n868 B.n867 47.4474
R1211 B.n867 B.n8 47.4474
R1212 B.n12 B.n8 47.4474
R1213 B.n860 B.n12 47.4474
R1214 B.n859 B.n858 47.4474
R1215 B.n858 B.n16 47.4474
R1216 B.n852 B.n16 47.4474
R1217 B.n852 B.n851 47.4474
R1218 B.n851 B.n850 47.4474
R1219 B.n850 B.n23 47.4474
R1220 B.n844 B.n843 47.4474
R1221 B.n843 B.n842 47.4474
R1222 B.n842 B.n30 47.4474
R1223 B.n836 B.n30 47.4474
R1224 B.n836 B.n835 47.4474
R1225 B.n835 B.n834 47.4474
R1226 B.n828 B.n40 47.4474
R1227 B.n828 B.n827 47.4474
R1228 B.n827 B.n826 47.4474
R1229 B.n826 B.n44 47.4474
R1230 B.n820 B.n44 47.4474
R1231 B.n820 B.n819 47.4474
R1232 B.n818 B.n51 47.4474
R1233 B.n812 B.n51 47.4474
R1234 B.n812 B.n811 47.4474
R1235 B.n811 B.n810 47.4474
R1236 B.n810 B.n58 47.4474
R1237 B.n804 B.n58 47.4474
R1238 B.n804 B.n803 47.4474
R1239 B.n803 B.n802 47.4474
R1240 B.n802 B.n65 47.4474
R1241 B.n796 B.n65 47.4474
R1242 B.n795 B.n794 47.4474
R1243 B.n794 B.n72 47.4474
R1244 B.n788 B.n72 47.4474
R1245 B.n788 B.n787 47.4474
R1246 B.n787 B.n786 47.4474
R1247 B.n786 B.n79 47.4474
R1248 B.n128 B.n127 46.7399
R1249 B.n126 B.n125 46.7399
R1250 B.n423 B.n422 46.7399
R1251 B.n420 B.n419 46.7399
R1252 B.t3 B.n337 43.2609
R1253 B.n819 B.t21 43.2609
R1254 B.n667 B.t5 39.0744
R1255 B.n834 B.t6 39.0744
R1256 B.n365 B.t15 37.6789
R1257 B.t8 B.n795 37.6789
R1258 B.t0 B.n310 34.8879
R1259 B.t4 B.n23 34.8879
R1260 B.n591 B.n590 32.6249
R1261 B.n425 B.n371 32.6249
R1262 B.n776 B.n775 32.6249
R1263 B.n783 B.n782 32.6249
R1264 B.n710 B.t1 30.7014
R1265 B.n860 B.t2 30.7014
R1266 B B.n872 18.0485
R1267 B.n302 B.t1 16.7465
R1268 B.t2 B.n859 16.7465
R1269 B.n685 B.t0 12.56
R1270 B.n844 B.t4 12.56
R1271 B.n592 B.n591 10.6151
R1272 B.n592 B.n367 10.6151
R1273 B.n602 B.n367 10.6151
R1274 B.n603 B.n602 10.6151
R1275 B.n604 B.n603 10.6151
R1276 B.n604 B.n359 10.6151
R1277 B.n614 B.n359 10.6151
R1278 B.n615 B.n614 10.6151
R1279 B.n616 B.n615 10.6151
R1280 B.n616 B.n351 10.6151
R1281 B.n626 B.n351 10.6151
R1282 B.n627 B.n626 10.6151
R1283 B.n628 B.n627 10.6151
R1284 B.n628 B.n343 10.6151
R1285 B.n638 B.n343 10.6151
R1286 B.n639 B.n638 10.6151
R1287 B.n640 B.n639 10.6151
R1288 B.n640 B.n335 10.6151
R1289 B.n650 B.n335 10.6151
R1290 B.n651 B.n650 10.6151
R1291 B.n652 B.n651 10.6151
R1292 B.n652 B.n327 10.6151
R1293 B.n663 B.n327 10.6151
R1294 B.n664 B.n663 10.6151
R1295 B.n665 B.n664 10.6151
R1296 B.n665 B.n320 10.6151
R1297 B.n675 B.n320 10.6151
R1298 B.n676 B.n675 10.6151
R1299 B.n677 B.n676 10.6151
R1300 B.n677 B.n312 10.6151
R1301 B.n687 B.n312 10.6151
R1302 B.n688 B.n687 10.6151
R1303 B.n689 B.n688 10.6151
R1304 B.n689 B.n304 10.6151
R1305 B.n699 B.n304 10.6151
R1306 B.n700 B.n699 10.6151
R1307 B.n701 B.n700 10.6151
R1308 B.n701 B.n296 10.6151
R1309 B.n712 B.n296 10.6151
R1310 B.n713 B.n712 10.6151
R1311 B.n714 B.n713 10.6151
R1312 B.n714 B.n0 10.6151
R1313 B.n590 B.n375 10.6151
R1314 B.n585 B.n375 10.6151
R1315 B.n585 B.n584 10.6151
R1316 B.n584 B.n583 10.6151
R1317 B.n583 B.n580 10.6151
R1318 B.n580 B.n579 10.6151
R1319 B.n579 B.n576 10.6151
R1320 B.n576 B.n575 10.6151
R1321 B.n575 B.n572 10.6151
R1322 B.n572 B.n571 10.6151
R1323 B.n571 B.n568 10.6151
R1324 B.n568 B.n567 10.6151
R1325 B.n567 B.n564 10.6151
R1326 B.n564 B.n563 10.6151
R1327 B.n563 B.n560 10.6151
R1328 B.n560 B.n559 10.6151
R1329 B.n559 B.n556 10.6151
R1330 B.n556 B.n555 10.6151
R1331 B.n555 B.n552 10.6151
R1332 B.n552 B.n551 10.6151
R1333 B.n551 B.n548 10.6151
R1334 B.n548 B.n547 10.6151
R1335 B.n547 B.n544 10.6151
R1336 B.n544 B.n543 10.6151
R1337 B.n543 B.n540 10.6151
R1338 B.n540 B.n539 10.6151
R1339 B.n539 B.n536 10.6151
R1340 B.n536 B.n535 10.6151
R1341 B.n535 B.n532 10.6151
R1342 B.n532 B.n531 10.6151
R1343 B.n531 B.n528 10.6151
R1344 B.n528 B.n527 10.6151
R1345 B.n527 B.n524 10.6151
R1346 B.n524 B.n523 10.6151
R1347 B.n523 B.n520 10.6151
R1348 B.n520 B.n519 10.6151
R1349 B.n516 B.n515 10.6151
R1350 B.n515 B.n512 10.6151
R1351 B.n512 B.n511 10.6151
R1352 B.n511 B.n508 10.6151
R1353 B.n508 B.n507 10.6151
R1354 B.n507 B.n504 10.6151
R1355 B.n504 B.n503 10.6151
R1356 B.n503 B.n500 10.6151
R1357 B.n500 B.n499 10.6151
R1358 B.n496 B.n495 10.6151
R1359 B.n495 B.n492 10.6151
R1360 B.n492 B.n491 10.6151
R1361 B.n491 B.n488 10.6151
R1362 B.n488 B.n487 10.6151
R1363 B.n487 B.n484 10.6151
R1364 B.n484 B.n483 10.6151
R1365 B.n483 B.n480 10.6151
R1366 B.n480 B.n479 10.6151
R1367 B.n479 B.n476 10.6151
R1368 B.n476 B.n475 10.6151
R1369 B.n475 B.n472 10.6151
R1370 B.n472 B.n471 10.6151
R1371 B.n471 B.n468 10.6151
R1372 B.n468 B.n467 10.6151
R1373 B.n467 B.n464 10.6151
R1374 B.n464 B.n463 10.6151
R1375 B.n463 B.n460 10.6151
R1376 B.n460 B.n459 10.6151
R1377 B.n459 B.n456 10.6151
R1378 B.n456 B.n455 10.6151
R1379 B.n455 B.n452 10.6151
R1380 B.n452 B.n451 10.6151
R1381 B.n451 B.n448 10.6151
R1382 B.n448 B.n447 10.6151
R1383 B.n447 B.n444 10.6151
R1384 B.n444 B.n443 10.6151
R1385 B.n443 B.n440 10.6151
R1386 B.n440 B.n439 10.6151
R1387 B.n439 B.n436 10.6151
R1388 B.n436 B.n435 10.6151
R1389 B.n435 B.n432 10.6151
R1390 B.n432 B.n431 10.6151
R1391 B.n431 B.n428 10.6151
R1392 B.n428 B.n427 10.6151
R1393 B.n427 B.n425 10.6151
R1394 B.n596 B.n371 10.6151
R1395 B.n597 B.n596 10.6151
R1396 B.n598 B.n597 10.6151
R1397 B.n598 B.n362 10.6151
R1398 B.n608 B.n362 10.6151
R1399 B.n609 B.n608 10.6151
R1400 B.n610 B.n609 10.6151
R1401 B.n610 B.n355 10.6151
R1402 B.n620 B.n355 10.6151
R1403 B.n621 B.n620 10.6151
R1404 B.n622 B.n621 10.6151
R1405 B.n622 B.n347 10.6151
R1406 B.n632 B.n347 10.6151
R1407 B.n633 B.n632 10.6151
R1408 B.n634 B.n633 10.6151
R1409 B.n634 B.n339 10.6151
R1410 B.n644 B.n339 10.6151
R1411 B.n645 B.n644 10.6151
R1412 B.n646 B.n645 10.6151
R1413 B.n646 B.n331 10.6151
R1414 B.n656 B.n331 10.6151
R1415 B.n657 B.n656 10.6151
R1416 B.n658 B.n657 10.6151
R1417 B.n658 B.n324 10.6151
R1418 B.n669 B.n324 10.6151
R1419 B.n670 B.n669 10.6151
R1420 B.n671 B.n670 10.6151
R1421 B.n671 B.n316 10.6151
R1422 B.n681 B.n316 10.6151
R1423 B.n682 B.n681 10.6151
R1424 B.n683 B.n682 10.6151
R1425 B.n683 B.n308 10.6151
R1426 B.n693 B.n308 10.6151
R1427 B.n694 B.n693 10.6151
R1428 B.n695 B.n694 10.6151
R1429 B.n695 B.n299 10.6151
R1430 B.n705 B.n299 10.6151
R1431 B.n706 B.n705 10.6151
R1432 B.n708 B.n706 10.6151
R1433 B.n708 B.n707 10.6151
R1434 B.n707 B.n292 10.6151
R1435 B.n719 B.n292 10.6151
R1436 B.n720 B.n719 10.6151
R1437 B.n721 B.n720 10.6151
R1438 B.n722 B.n721 10.6151
R1439 B.n723 B.n722 10.6151
R1440 B.n726 B.n723 10.6151
R1441 B.n727 B.n726 10.6151
R1442 B.n728 B.n727 10.6151
R1443 B.n729 B.n728 10.6151
R1444 B.n731 B.n729 10.6151
R1445 B.n732 B.n731 10.6151
R1446 B.n733 B.n732 10.6151
R1447 B.n734 B.n733 10.6151
R1448 B.n736 B.n734 10.6151
R1449 B.n737 B.n736 10.6151
R1450 B.n738 B.n737 10.6151
R1451 B.n739 B.n738 10.6151
R1452 B.n741 B.n739 10.6151
R1453 B.n742 B.n741 10.6151
R1454 B.n743 B.n742 10.6151
R1455 B.n744 B.n743 10.6151
R1456 B.n746 B.n744 10.6151
R1457 B.n747 B.n746 10.6151
R1458 B.n748 B.n747 10.6151
R1459 B.n749 B.n748 10.6151
R1460 B.n751 B.n749 10.6151
R1461 B.n752 B.n751 10.6151
R1462 B.n753 B.n752 10.6151
R1463 B.n754 B.n753 10.6151
R1464 B.n756 B.n754 10.6151
R1465 B.n757 B.n756 10.6151
R1466 B.n758 B.n757 10.6151
R1467 B.n759 B.n758 10.6151
R1468 B.n761 B.n759 10.6151
R1469 B.n762 B.n761 10.6151
R1470 B.n763 B.n762 10.6151
R1471 B.n764 B.n763 10.6151
R1472 B.n766 B.n764 10.6151
R1473 B.n767 B.n766 10.6151
R1474 B.n768 B.n767 10.6151
R1475 B.n769 B.n768 10.6151
R1476 B.n771 B.n769 10.6151
R1477 B.n772 B.n771 10.6151
R1478 B.n773 B.n772 10.6151
R1479 B.n774 B.n773 10.6151
R1480 B.n775 B.n774 10.6151
R1481 B.n864 B.n1 10.6151
R1482 B.n864 B.n863 10.6151
R1483 B.n863 B.n862 10.6151
R1484 B.n862 B.n10 10.6151
R1485 B.n856 B.n10 10.6151
R1486 B.n856 B.n855 10.6151
R1487 B.n855 B.n854 10.6151
R1488 B.n854 B.n18 10.6151
R1489 B.n848 B.n18 10.6151
R1490 B.n848 B.n847 10.6151
R1491 B.n847 B.n846 10.6151
R1492 B.n846 B.n25 10.6151
R1493 B.n840 B.n25 10.6151
R1494 B.n840 B.n839 10.6151
R1495 B.n839 B.n838 10.6151
R1496 B.n838 B.n32 10.6151
R1497 B.n832 B.n32 10.6151
R1498 B.n832 B.n831 10.6151
R1499 B.n831 B.n830 10.6151
R1500 B.n830 B.n38 10.6151
R1501 B.n824 B.n38 10.6151
R1502 B.n824 B.n823 10.6151
R1503 B.n823 B.n822 10.6151
R1504 B.n822 B.n46 10.6151
R1505 B.n816 B.n46 10.6151
R1506 B.n816 B.n815 10.6151
R1507 B.n815 B.n814 10.6151
R1508 B.n814 B.n53 10.6151
R1509 B.n808 B.n53 10.6151
R1510 B.n808 B.n807 10.6151
R1511 B.n807 B.n806 10.6151
R1512 B.n806 B.n60 10.6151
R1513 B.n800 B.n60 10.6151
R1514 B.n800 B.n799 10.6151
R1515 B.n799 B.n798 10.6151
R1516 B.n798 B.n67 10.6151
R1517 B.n792 B.n67 10.6151
R1518 B.n792 B.n791 10.6151
R1519 B.n791 B.n790 10.6151
R1520 B.n790 B.n74 10.6151
R1521 B.n784 B.n74 10.6151
R1522 B.n784 B.n783 10.6151
R1523 B.n782 B.n81 10.6151
R1524 B.n130 B.n81 10.6151
R1525 B.n131 B.n130 10.6151
R1526 B.n134 B.n131 10.6151
R1527 B.n135 B.n134 10.6151
R1528 B.n138 B.n135 10.6151
R1529 B.n139 B.n138 10.6151
R1530 B.n142 B.n139 10.6151
R1531 B.n143 B.n142 10.6151
R1532 B.n146 B.n143 10.6151
R1533 B.n147 B.n146 10.6151
R1534 B.n150 B.n147 10.6151
R1535 B.n151 B.n150 10.6151
R1536 B.n154 B.n151 10.6151
R1537 B.n155 B.n154 10.6151
R1538 B.n158 B.n155 10.6151
R1539 B.n159 B.n158 10.6151
R1540 B.n162 B.n159 10.6151
R1541 B.n163 B.n162 10.6151
R1542 B.n166 B.n163 10.6151
R1543 B.n167 B.n166 10.6151
R1544 B.n170 B.n167 10.6151
R1545 B.n171 B.n170 10.6151
R1546 B.n174 B.n171 10.6151
R1547 B.n175 B.n174 10.6151
R1548 B.n178 B.n175 10.6151
R1549 B.n179 B.n178 10.6151
R1550 B.n182 B.n179 10.6151
R1551 B.n183 B.n182 10.6151
R1552 B.n186 B.n183 10.6151
R1553 B.n187 B.n186 10.6151
R1554 B.n190 B.n187 10.6151
R1555 B.n191 B.n190 10.6151
R1556 B.n194 B.n191 10.6151
R1557 B.n195 B.n194 10.6151
R1558 B.n198 B.n195 10.6151
R1559 B.n203 B.n200 10.6151
R1560 B.n204 B.n203 10.6151
R1561 B.n207 B.n204 10.6151
R1562 B.n208 B.n207 10.6151
R1563 B.n211 B.n208 10.6151
R1564 B.n212 B.n211 10.6151
R1565 B.n215 B.n212 10.6151
R1566 B.n216 B.n215 10.6151
R1567 B.n219 B.n216 10.6151
R1568 B.n224 B.n221 10.6151
R1569 B.n225 B.n224 10.6151
R1570 B.n228 B.n225 10.6151
R1571 B.n229 B.n228 10.6151
R1572 B.n232 B.n229 10.6151
R1573 B.n233 B.n232 10.6151
R1574 B.n236 B.n233 10.6151
R1575 B.n237 B.n236 10.6151
R1576 B.n240 B.n237 10.6151
R1577 B.n241 B.n240 10.6151
R1578 B.n244 B.n241 10.6151
R1579 B.n245 B.n244 10.6151
R1580 B.n248 B.n245 10.6151
R1581 B.n249 B.n248 10.6151
R1582 B.n252 B.n249 10.6151
R1583 B.n253 B.n252 10.6151
R1584 B.n256 B.n253 10.6151
R1585 B.n257 B.n256 10.6151
R1586 B.n260 B.n257 10.6151
R1587 B.n261 B.n260 10.6151
R1588 B.n264 B.n261 10.6151
R1589 B.n265 B.n264 10.6151
R1590 B.n268 B.n265 10.6151
R1591 B.n269 B.n268 10.6151
R1592 B.n272 B.n269 10.6151
R1593 B.n273 B.n272 10.6151
R1594 B.n276 B.n273 10.6151
R1595 B.n277 B.n276 10.6151
R1596 B.n280 B.n277 10.6151
R1597 B.n281 B.n280 10.6151
R1598 B.n284 B.n281 10.6151
R1599 B.n285 B.n284 10.6151
R1600 B.n288 B.n285 10.6151
R1601 B.n290 B.n288 10.6151
R1602 B.n291 B.n290 10.6151
R1603 B.n776 B.n291 10.6151
R1604 B.n612 B.t15 9.76897
R1605 B.n796 B.t8 9.76897
R1606 B.n519 B.n421 9.36635
R1607 B.n496 B.n424 9.36635
R1608 B.n199 B.n198 9.36635
R1609 B.n221 B.n220 9.36635
R1610 B.n660 B.t5 8.37348
R1611 B.n40 B.t6 8.37348
R1612 B.n872 B.n0 8.11757
R1613 B.n872 B.n1 8.11757
R1614 B.n642 B.t3 4.18699
R1615 B.t21 B.n818 4.18699
R1616 B.n516 B.n421 1.24928
R1617 B.n499 B.n424 1.24928
R1618 B.n200 B.n199 1.24928
R1619 B.n220 B.n219 1.24928
R1620 VP.n15 VP.n12 161.3
R1621 VP.n17 VP.n16 161.3
R1622 VP.n18 VP.n11 161.3
R1623 VP.n20 VP.n19 161.3
R1624 VP.n22 VP.n10 161.3
R1625 VP.n24 VP.n23 161.3
R1626 VP.n25 VP.n9 161.3
R1627 VP.n27 VP.n26 161.3
R1628 VP.n28 VP.n8 161.3
R1629 VP.n54 VP.n0 161.3
R1630 VP.n53 VP.n52 161.3
R1631 VP.n51 VP.n1 161.3
R1632 VP.n50 VP.n49 161.3
R1633 VP.n48 VP.n2 161.3
R1634 VP.n46 VP.n45 161.3
R1635 VP.n44 VP.n3 161.3
R1636 VP.n43 VP.n42 161.3
R1637 VP.n41 VP.n4 161.3
R1638 VP.n39 VP.n38 161.3
R1639 VP.n37 VP.n5 161.3
R1640 VP.n36 VP.n35 161.3
R1641 VP.n34 VP.n6 161.3
R1642 VP.n33 VP.n32 161.3
R1643 VP.n13 VP.t1 155.309
R1644 VP.n7 VP.t7 121.543
R1645 VP.n40 VP.t5 121.543
R1646 VP.n47 VP.t3 121.543
R1647 VP.n55 VP.t0 121.543
R1648 VP.n29 VP.t6 121.543
R1649 VP.n21 VP.t4 121.543
R1650 VP.n14 VP.t2 121.543
R1651 VP.n31 VP.n7 92.8955
R1652 VP.n56 VP.n55 92.8955
R1653 VP.n30 VP.n29 92.8955
R1654 VP.n42 VP.n3 56.5193
R1655 VP.n16 VP.n11 56.5193
R1656 VP.n35 VP.n34 56.0336
R1657 VP.n53 VP.n1 56.0336
R1658 VP.n27 VP.n9 56.0336
R1659 VP.n14 VP.n13 48.1291
R1660 VP.n31 VP.n30 47.3329
R1661 VP.n35 VP.n5 24.9531
R1662 VP.n49 VP.n1 24.9531
R1663 VP.n23 VP.n9 24.9531
R1664 VP.n34 VP.n33 24.4675
R1665 VP.n39 VP.n5 24.4675
R1666 VP.n42 VP.n41 24.4675
R1667 VP.n46 VP.n3 24.4675
R1668 VP.n49 VP.n48 24.4675
R1669 VP.n54 VP.n53 24.4675
R1670 VP.n28 VP.n27 24.4675
R1671 VP.n20 VP.n11 24.4675
R1672 VP.n23 VP.n22 24.4675
R1673 VP.n16 VP.n15 24.4675
R1674 VP.n41 VP.n40 22.2655
R1675 VP.n47 VP.n46 22.2655
R1676 VP.n21 VP.n20 22.2655
R1677 VP.n15 VP.n14 22.2655
R1678 VP.n33 VP.n7 17.8614
R1679 VP.n55 VP.n54 17.8614
R1680 VP.n29 VP.n28 17.8614
R1681 VP.n13 VP.n12 9.16971
R1682 VP.n40 VP.n39 2.20253
R1683 VP.n48 VP.n47 2.20253
R1684 VP.n22 VP.n21 2.20253
R1685 VP.n30 VP.n8 0.278367
R1686 VP.n32 VP.n31 0.278367
R1687 VP.n56 VP.n0 0.278367
R1688 VP.n17 VP.n12 0.189894
R1689 VP.n18 VP.n17 0.189894
R1690 VP.n19 VP.n18 0.189894
R1691 VP.n19 VP.n10 0.189894
R1692 VP.n24 VP.n10 0.189894
R1693 VP.n25 VP.n24 0.189894
R1694 VP.n26 VP.n25 0.189894
R1695 VP.n26 VP.n8 0.189894
R1696 VP.n32 VP.n6 0.189894
R1697 VP.n36 VP.n6 0.189894
R1698 VP.n37 VP.n36 0.189894
R1699 VP.n38 VP.n37 0.189894
R1700 VP.n38 VP.n4 0.189894
R1701 VP.n43 VP.n4 0.189894
R1702 VP.n44 VP.n43 0.189894
R1703 VP.n45 VP.n44 0.189894
R1704 VP.n45 VP.n2 0.189894
R1705 VP.n50 VP.n2 0.189894
R1706 VP.n51 VP.n50 0.189894
R1707 VP.n52 VP.n51 0.189894
R1708 VP.n52 VP.n0 0.189894
R1709 VP VP.n56 0.153454
R1710 VDD1 VDD1.n0 66.8769
R1711 VDD1.n3 VDD1.n2 66.7632
R1712 VDD1.n3 VDD1.n1 66.7632
R1713 VDD1.n5 VDD1.n4 65.7798
R1714 VDD1.n5 VDD1.n3 42.6905
R1715 VDD1.n4 VDD1.t3 1.88801
R1716 VDD1.n4 VDD1.t1 1.88801
R1717 VDD1.n0 VDD1.t6 1.88801
R1718 VDD1.n0 VDD1.t5 1.88801
R1719 VDD1.n2 VDD1.t4 1.88801
R1720 VDD1.n2 VDD1.t7 1.88801
R1721 VDD1.n1 VDD1.t0 1.88801
R1722 VDD1.n1 VDD1.t2 1.88801
R1723 VDD1 VDD1.n5 0.981103
C0 VDD2 VP 0.46439f
C1 VDD2 VN 7.28939f
C2 VDD2 VTAIL 7.55656f
C3 VDD2 VDD1 1.50716f
C4 VN VP 6.74875f
C5 VTAIL VP 7.59676f
C6 VDD1 VP 7.601799f
C7 VTAIL VN 7.58265f
C8 VDD1 VN 0.150841f
C9 VDD1 VTAIL 7.50563f
C10 VDD2 B 4.732098f
C11 VDD1 B 5.111438f
C12 VTAIL B 9.227307f
C13 VN B 13.40582f
C14 VP B 11.953016f
C15 VDD1.t6 B 0.205213f
C16 VDD1.t5 B 0.205213f
C17 VDD1.n0 B 1.82323f
C18 VDD1.t0 B 0.205213f
C19 VDD1.t2 B 0.205213f
C20 VDD1.n1 B 1.82233f
C21 VDD1.t4 B 0.205213f
C22 VDD1.t7 B 0.205213f
C23 VDD1.n2 B 1.82233f
C24 VDD1.n3 B 2.89961f
C25 VDD1.t3 B 0.205213f
C26 VDD1.t1 B 0.205213f
C27 VDD1.n4 B 1.81563f
C28 VDD1.n5 B 2.65385f
C29 VP.n0 B 0.034549f
C30 VP.t0 B 1.55146f
C31 VP.n1 B 0.031289f
C32 VP.n2 B 0.026205f
C33 VP.t3 B 1.55146f
C34 VP.n3 B 0.038255f
C35 VP.n4 B 0.026205f
C36 VP.t5 B 1.55146f
C37 VP.n5 B 0.049298f
C38 VP.n6 B 0.026205f
C39 VP.t7 B 1.55146f
C40 VP.n7 B 0.638701f
C41 VP.n8 B 0.034549f
C42 VP.t6 B 1.55146f
C43 VP.n9 B 0.031289f
C44 VP.n10 B 0.026205f
C45 VP.t4 B 1.55146f
C46 VP.n11 B 0.038255f
C47 VP.n12 B 0.220171f
C48 VP.t2 B 1.55146f
C49 VP.t1 B 1.70295f
C50 VP.n13 B 0.615495f
C51 VP.n14 B 0.633569f
C52 VP.n15 B 0.046668f
C53 VP.n16 B 0.038255f
C54 VP.n17 B 0.026205f
C55 VP.n18 B 0.026205f
C56 VP.n19 B 0.026205f
C57 VP.n20 B 0.046668f
C58 VP.n21 B 0.558237f
C59 VP.n22 B 0.026896f
C60 VP.n23 B 0.049298f
C61 VP.n24 B 0.026205f
C62 VP.n25 B 0.026205f
C63 VP.n26 B 0.026205f
C64 VP.n27 B 0.044762f
C65 VP.n28 B 0.042328f
C66 VP.n29 B 0.638701f
C67 VP.n30 B 1.33413f
C68 VP.n31 B 1.35404f
C69 VP.n32 B 0.034549f
C70 VP.n33 B 0.042328f
C71 VP.n34 B 0.044762f
C72 VP.n35 B 0.031289f
C73 VP.n36 B 0.026205f
C74 VP.n37 B 0.026205f
C75 VP.n38 B 0.026205f
C76 VP.n39 B 0.026896f
C77 VP.n40 B 0.558237f
C78 VP.n41 B 0.046668f
C79 VP.n42 B 0.038255f
C80 VP.n43 B 0.026205f
C81 VP.n44 B 0.026205f
C82 VP.n45 B 0.026205f
C83 VP.n46 B 0.046668f
C84 VP.n47 B 0.558237f
C85 VP.n48 B 0.026896f
C86 VP.n49 B 0.049298f
C87 VP.n50 B 0.026205f
C88 VP.n51 B 0.026205f
C89 VP.n52 B 0.026205f
C90 VP.n53 B 0.044762f
C91 VP.n54 B 0.042328f
C92 VP.n55 B 0.638701f
C93 VP.n56 B 0.03362f
C94 VTAIL.t13 B 0.165381f
C95 VTAIL.t10 B 0.165381f
C96 VTAIL.n0 B 1.40976f
C97 VTAIL.n1 B 0.324814f
C98 VTAIL.t14 B 1.79804f
C99 VTAIL.n2 B 0.414038f
C100 VTAIL.t1 B 1.79804f
C101 VTAIL.n3 B 0.414038f
C102 VTAIL.t5 B 0.165381f
C103 VTAIL.t0 B 0.165381f
C104 VTAIL.n4 B 1.40976f
C105 VTAIL.n5 B 0.454631f
C106 VTAIL.t3 B 1.79804f
C107 VTAIL.n6 B 1.36974f
C108 VTAIL.t11 B 1.79804f
C109 VTAIL.n7 B 1.36973f
C110 VTAIL.t12 B 0.165381f
C111 VTAIL.t15 B 0.165381f
C112 VTAIL.n8 B 1.40976f
C113 VTAIL.n9 B 0.454627f
C114 VTAIL.t9 B 1.79804f
C115 VTAIL.n10 B 0.414034f
C116 VTAIL.t2 B 1.79804f
C117 VTAIL.n11 B 0.414034f
C118 VTAIL.t4 B 0.165381f
C119 VTAIL.t6 B 0.165381f
C120 VTAIL.n12 B 1.40976f
C121 VTAIL.n13 B 0.454627f
C122 VTAIL.t7 B 1.79804f
C123 VTAIL.n14 B 1.36974f
C124 VTAIL.t8 B 1.79804f
C125 VTAIL.n15 B 1.366f
C126 VDD2.t3 B 0.203729f
C127 VDD2.t7 B 0.203729f
C128 VDD2.n0 B 1.80915f
C129 VDD2.t1 B 0.203729f
C130 VDD2.t0 B 0.203729f
C131 VDD2.n1 B 1.80915f
C132 VDD2.n2 B 2.82708f
C133 VDD2.t4 B 0.203729f
C134 VDD2.t2 B 0.203729f
C135 VDD2.n3 B 1.8025f
C136 VDD2.n4 B 2.60464f
C137 VDD2.t6 B 0.203729f
C138 VDD2.t5 B 0.203729f
C139 VDD2.n5 B 1.80911f
C140 VN.n0 B 0.034018f
C141 VN.t7 B 1.52764f
C142 VN.n1 B 0.030808f
C143 VN.n2 B 0.025803f
C144 VN.t5 B 1.52764f
C145 VN.n3 B 0.037667f
C146 VN.n4 B 0.21679f
C147 VN.t2 B 1.52764f
C148 VN.t1 B 1.6768f
C149 VN.n5 B 0.606044f
C150 VN.n6 B 0.623841f
C151 VN.n7 B 0.045952f
C152 VN.n8 B 0.037667f
C153 VN.n9 B 0.025803f
C154 VN.n10 B 0.025803f
C155 VN.n11 B 0.025803f
C156 VN.n12 B 0.045952f
C157 VN.n13 B 0.549665f
C158 VN.n14 B 0.026483f
C159 VN.n15 B 0.048541f
C160 VN.n16 B 0.025803f
C161 VN.n17 B 0.025803f
C162 VN.n18 B 0.025803f
C163 VN.n19 B 0.044075f
C164 VN.n20 B 0.041678f
C165 VN.n21 B 0.628894f
C166 VN.n22 B 0.033104f
C167 VN.n23 B 0.034018f
C168 VN.t4 B 1.52764f
C169 VN.n24 B 0.030808f
C170 VN.n25 B 0.025803f
C171 VN.t3 B 1.52764f
C172 VN.n26 B 0.037667f
C173 VN.n27 B 0.21679f
C174 VN.t0 B 1.52764f
C175 VN.t6 B 1.6768f
C176 VN.n28 B 0.606044f
C177 VN.n29 B 0.623841f
C178 VN.n30 B 0.045952f
C179 VN.n31 B 0.037667f
C180 VN.n32 B 0.025803f
C181 VN.n33 B 0.025803f
C182 VN.n34 B 0.025803f
C183 VN.n35 B 0.045952f
C184 VN.n36 B 0.549665f
C185 VN.n37 B 0.026483f
C186 VN.n38 B 0.048541f
C187 VN.n39 B 0.025803f
C188 VN.n40 B 0.025803f
C189 VN.n41 B 0.025803f
C190 VN.n42 B 0.044075f
C191 VN.n43 B 0.041678f
C192 VN.n44 B 0.628894f
C193 VN.n45 B 1.32764f
.ends

