* NGSPICE file created from diff_pair_sample_0758.ext - technology: sky130A

.subckt diff_pair_sample_0758 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t11 VP.t0 VDD1.t4 B.t3 sky130_fd_pr__nfet_01v8 ad=1.68135 pd=10.52 as=1.68135 ps=10.52 w=10.19 l=2.52
X1 VDD1.t3 VP.t1 VTAIL.t10 B.t4 sky130_fd_pr__nfet_01v8 ad=1.68135 pd=10.52 as=3.9741 ps=21.16 w=10.19 l=2.52
X2 VDD2.t5 VN.t0 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=3.9741 pd=21.16 as=1.68135 ps=10.52 w=10.19 l=2.52
X3 VDD2.t4 VN.t1 VTAIL.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=3.9741 pd=21.16 as=1.68135 ps=10.52 w=10.19 l=2.52
X4 B.t19 B.t17 B.t18 B.t14 sky130_fd_pr__nfet_01v8 ad=3.9741 pd=21.16 as=0 ps=0 w=10.19 l=2.52
X5 VTAIL.t3 VN.t2 VDD2.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=1.68135 pd=10.52 as=1.68135 ps=10.52 w=10.19 l=2.52
X6 B.t16 B.t13 B.t15 B.t14 sky130_fd_pr__nfet_01v8 ad=3.9741 pd=21.16 as=0 ps=0 w=10.19 l=2.52
X7 VDD2.t2 VN.t3 VTAIL.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=1.68135 pd=10.52 as=3.9741 ps=21.16 w=10.19 l=2.52
X8 VTAIL.t9 VP.t2 VDD1.t5 B.t0 sky130_fd_pr__nfet_01v8 ad=1.68135 pd=10.52 as=1.68135 ps=10.52 w=10.19 l=2.52
X9 VDD2.t1 VN.t4 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=1.68135 pd=10.52 as=3.9741 ps=21.16 w=10.19 l=2.52
X10 B.t12 B.t10 B.t11 B.t7 sky130_fd_pr__nfet_01v8 ad=3.9741 pd=21.16 as=0 ps=0 w=10.19 l=2.52
X11 VDD1.t1 VP.t3 VTAIL.t8 B.t5 sky130_fd_pr__nfet_01v8 ad=3.9741 pd=21.16 as=1.68135 ps=10.52 w=10.19 l=2.52
X12 VTAIL.t0 VN.t5 VDD2.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=1.68135 pd=10.52 as=1.68135 ps=10.52 w=10.19 l=2.52
X13 VDD1.t0 VP.t4 VTAIL.t7 B.t1 sky130_fd_pr__nfet_01v8 ad=3.9741 pd=21.16 as=1.68135 ps=10.52 w=10.19 l=2.52
X14 B.t9 B.t6 B.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=3.9741 pd=21.16 as=0 ps=0 w=10.19 l=2.52
X15 VDD1.t2 VP.t5 VTAIL.t6 B.t2 sky130_fd_pr__nfet_01v8 ad=1.68135 pd=10.52 as=3.9741 ps=21.16 w=10.19 l=2.52
R0 VP.n13 VP.n12 161.3
R1 VP.n14 VP.n9 161.3
R2 VP.n16 VP.n15 161.3
R3 VP.n17 VP.n8 161.3
R4 VP.n19 VP.n18 161.3
R5 VP.n20 VP.n7 161.3
R6 VP.n42 VP.n0 161.3
R7 VP.n41 VP.n40 161.3
R8 VP.n39 VP.n1 161.3
R9 VP.n38 VP.n37 161.3
R10 VP.n36 VP.n2 161.3
R11 VP.n35 VP.n34 161.3
R12 VP.n33 VP.n32 161.3
R13 VP.n31 VP.n4 161.3
R14 VP.n30 VP.n29 161.3
R15 VP.n28 VP.n5 161.3
R16 VP.n27 VP.n26 161.3
R17 VP.n25 VP.n6 161.3
R18 VP.n11 VP.t3 129.466
R19 VP.n24 VP.n23 105.864
R20 VP.n44 VP.n43 105.864
R21 VP.n22 VP.n21 105.864
R22 VP.n24 VP.t4 97.4525
R23 VP.n3 VP.t0 97.4525
R24 VP.n43 VP.t5 97.4525
R25 VP.n21 VP.t1 97.4525
R26 VP.n10 VP.t2 97.4525
R27 VP.n11 VP.n10 59.8984
R28 VP.n30 VP.n5 56.5193
R29 VP.n37 VP.n1 56.5193
R30 VP.n15 VP.n8 56.5193
R31 VP.n23 VP.n22 46.9125
R32 VP.n26 VP.n25 24.4675
R33 VP.n26 VP.n5 24.4675
R34 VP.n31 VP.n30 24.4675
R35 VP.n32 VP.n31 24.4675
R36 VP.n36 VP.n35 24.4675
R37 VP.n37 VP.n36 24.4675
R38 VP.n41 VP.n1 24.4675
R39 VP.n42 VP.n41 24.4675
R40 VP.n19 VP.n8 24.4675
R41 VP.n20 VP.n19 24.4675
R42 VP.n14 VP.n13 24.4675
R43 VP.n15 VP.n14 24.4675
R44 VP.n32 VP.n3 12.234
R45 VP.n35 VP.n3 12.234
R46 VP.n13 VP.n10 12.234
R47 VP.n12 VP.n11 7.17115
R48 VP.n25 VP.n24 4.8939
R49 VP.n43 VP.n42 4.8939
R50 VP.n21 VP.n20 4.8939
R51 VP.n22 VP.n7 0.278367
R52 VP.n23 VP.n6 0.278367
R53 VP.n44 VP.n0 0.278367
R54 VP.n12 VP.n9 0.189894
R55 VP.n16 VP.n9 0.189894
R56 VP.n17 VP.n16 0.189894
R57 VP.n18 VP.n17 0.189894
R58 VP.n18 VP.n7 0.189894
R59 VP.n27 VP.n6 0.189894
R60 VP.n28 VP.n27 0.189894
R61 VP.n29 VP.n28 0.189894
R62 VP.n29 VP.n4 0.189894
R63 VP.n33 VP.n4 0.189894
R64 VP.n34 VP.n33 0.189894
R65 VP.n34 VP.n2 0.189894
R66 VP.n38 VP.n2 0.189894
R67 VP.n39 VP.n38 0.189894
R68 VP.n40 VP.n39 0.189894
R69 VP.n40 VP.n0 0.189894
R70 VP VP.n44 0.153454
R71 VDD1.n48 VDD1.n0 289.615
R72 VDD1.n101 VDD1.n53 289.615
R73 VDD1.n49 VDD1.n48 185
R74 VDD1.n47 VDD1.n46 185
R75 VDD1.n4 VDD1.n3 185
R76 VDD1.n41 VDD1.n40 185
R77 VDD1.n39 VDD1.n6 185
R78 VDD1.n38 VDD1.n37 185
R79 VDD1.n9 VDD1.n7 185
R80 VDD1.n32 VDD1.n31 185
R81 VDD1.n30 VDD1.n29 185
R82 VDD1.n13 VDD1.n12 185
R83 VDD1.n24 VDD1.n23 185
R84 VDD1.n22 VDD1.n21 185
R85 VDD1.n17 VDD1.n16 185
R86 VDD1.n69 VDD1.n68 185
R87 VDD1.n74 VDD1.n73 185
R88 VDD1.n76 VDD1.n75 185
R89 VDD1.n65 VDD1.n64 185
R90 VDD1.n82 VDD1.n81 185
R91 VDD1.n84 VDD1.n83 185
R92 VDD1.n61 VDD1.n60 185
R93 VDD1.n91 VDD1.n90 185
R94 VDD1.n92 VDD1.n59 185
R95 VDD1.n94 VDD1.n93 185
R96 VDD1.n57 VDD1.n56 185
R97 VDD1.n100 VDD1.n99 185
R98 VDD1.n102 VDD1.n101 185
R99 VDD1.n18 VDD1.t1 149.524
R100 VDD1.n70 VDD1.t0 149.524
R101 VDD1.n48 VDD1.n47 104.615
R102 VDD1.n47 VDD1.n3 104.615
R103 VDD1.n40 VDD1.n3 104.615
R104 VDD1.n40 VDD1.n39 104.615
R105 VDD1.n39 VDD1.n38 104.615
R106 VDD1.n38 VDD1.n7 104.615
R107 VDD1.n31 VDD1.n7 104.615
R108 VDD1.n31 VDD1.n30 104.615
R109 VDD1.n30 VDD1.n12 104.615
R110 VDD1.n23 VDD1.n12 104.615
R111 VDD1.n23 VDD1.n22 104.615
R112 VDD1.n22 VDD1.n16 104.615
R113 VDD1.n74 VDD1.n68 104.615
R114 VDD1.n75 VDD1.n74 104.615
R115 VDD1.n75 VDD1.n64 104.615
R116 VDD1.n82 VDD1.n64 104.615
R117 VDD1.n83 VDD1.n82 104.615
R118 VDD1.n83 VDD1.n60 104.615
R119 VDD1.n91 VDD1.n60 104.615
R120 VDD1.n92 VDD1.n91 104.615
R121 VDD1.n93 VDD1.n92 104.615
R122 VDD1.n93 VDD1.n56 104.615
R123 VDD1.n100 VDD1.n56 104.615
R124 VDD1.n101 VDD1.n100 104.615
R125 VDD1.n107 VDD1.n106 67.6596
R126 VDD1.n109 VDD1.n108 67.1008
R127 VDD1 VDD1.n52 55.2256
R128 VDD1.n107 VDD1.n105 55.1121
R129 VDD1.t1 VDD1.n16 52.3082
R130 VDD1.t0 VDD1.n68 52.3082
R131 VDD1.n109 VDD1.n107 42.2962
R132 VDD1.n41 VDD1.n6 13.1884
R133 VDD1.n94 VDD1.n59 13.1884
R134 VDD1.n42 VDD1.n4 12.8005
R135 VDD1.n37 VDD1.n8 12.8005
R136 VDD1.n90 VDD1.n89 12.8005
R137 VDD1.n95 VDD1.n57 12.8005
R138 VDD1.n46 VDD1.n45 12.0247
R139 VDD1.n36 VDD1.n9 12.0247
R140 VDD1.n88 VDD1.n61 12.0247
R141 VDD1.n99 VDD1.n98 12.0247
R142 VDD1.n49 VDD1.n2 11.249
R143 VDD1.n33 VDD1.n32 11.249
R144 VDD1.n85 VDD1.n84 11.249
R145 VDD1.n102 VDD1.n55 11.249
R146 VDD1.n50 VDD1.n0 10.4732
R147 VDD1.n29 VDD1.n11 10.4732
R148 VDD1.n81 VDD1.n63 10.4732
R149 VDD1.n103 VDD1.n53 10.4732
R150 VDD1.n18 VDD1.n17 10.2747
R151 VDD1.n70 VDD1.n69 10.2747
R152 VDD1.n28 VDD1.n13 9.69747
R153 VDD1.n80 VDD1.n65 9.69747
R154 VDD1.n52 VDD1.n51 9.45567
R155 VDD1.n105 VDD1.n104 9.45567
R156 VDD1.n20 VDD1.n19 9.3005
R157 VDD1.n15 VDD1.n14 9.3005
R158 VDD1.n26 VDD1.n25 9.3005
R159 VDD1.n28 VDD1.n27 9.3005
R160 VDD1.n11 VDD1.n10 9.3005
R161 VDD1.n34 VDD1.n33 9.3005
R162 VDD1.n36 VDD1.n35 9.3005
R163 VDD1.n8 VDD1.n5 9.3005
R164 VDD1.n51 VDD1.n50 9.3005
R165 VDD1.n2 VDD1.n1 9.3005
R166 VDD1.n45 VDD1.n44 9.3005
R167 VDD1.n43 VDD1.n42 9.3005
R168 VDD1.n104 VDD1.n103 9.3005
R169 VDD1.n55 VDD1.n54 9.3005
R170 VDD1.n98 VDD1.n97 9.3005
R171 VDD1.n96 VDD1.n95 9.3005
R172 VDD1.n72 VDD1.n71 9.3005
R173 VDD1.n67 VDD1.n66 9.3005
R174 VDD1.n78 VDD1.n77 9.3005
R175 VDD1.n80 VDD1.n79 9.3005
R176 VDD1.n63 VDD1.n62 9.3005
R177 VDD1.n86 VDD1.n85 9.3005
R178 VDD1.n88 VDD1.n87 9.3005
R179 VDD1.n89 VDD1.n58 9.3005
R180 VDD1.n25 VDD1.n24 8.92171
R181 VDD1.n77 VDD1.n76 8.92171
R182 VDD1.n21 VDD1.n15 8.14595
R183 VDD1.n73 VDD1.n67 8.14595
R184 VDD1.n20 VDD1.n17 7.3702
R185 VDD1.n72 VDD1.n69 7.3702
R186 VDD1.n21 VDD1.n20 5.81868
R187 VDD1.n73 VDD1.n72 5.81868
R188 VDD1.n24 VDD1.n15 5.04292
R189 VDD1.n76 VDD1.n67 5.04292
R190 VDD1.n25 VDD1.n13 4.26717
R191 VDD1.n77 VDD1.n65 4.26717
R192 VDD1.n52 VDD1.n0 3.49141
R193 VDD1.n29 VDD1.n28 3.49141
R194 VDD1.n81 VDD1.n80 3.49141
R195 VDD1.n105 VDD1.n53 3.49141
R196 VDD1.n19 VDD1.n18 2.84303
R197 VDD1.n71 VDD1.n70 2.84303
R198 VDD1.n50 VDD1.n49 2.71565
R199 VDD1.n32 VDD1.n11 2.71565
R200 VDD1.n84 VDD1.n63 2.71565
R201 VDD1.n103 VDD1.n102 2.71565
R202 VDD1.n108 VDD1.t5 1.94358
R203 VDD1.n108 VDD1.t3 1.94358
R204 VDD1.n106 VDD1.t4 1.94358
R205 VDD1.n106 VDD1.t2 1.94358
R206 VDD1.n46 VDD1.n2 1.93989
R207 VDD1.n33 VDD1.n9 1.93989
R208 VDD1.n85 VDD1.n61 1.93989
R209 VDD1.n99 VDD1.n55 1.93989
R210 VDD1.n45 VDD1.n4 1.16414
R211 VDD1.n37 VDD1.n36 1.16414
R212 VDD1.n90 VDD1.n88 1.16414
R213 VDD1.n98 VDD1.n57 1.16414
R214 VDD1 VDD1.n109 0.556535
R215 VDD1.n42 VDD1.n41 0.388379
R216 VDD1.n8 VDD1.n6 0.388379
R217 VDD1.n89 VDD1.n59 0.388379
R218 VDD1.n95 VDD1.n94 0.388379
R219 VDD1.n51 VDD1.n1 0.155672
R220 VDD1.n44 VDD1.n1 0.155672
R221 VDD1.n44 VDD1.n43 0.155672
R222 VDD1.n43 VDD1.n5 0.155672
R223 VDD1.n35 VDD1.n5 0.155672
R224 VDD1.n35 VDD1.n34 0.155672
R225 VDD1.n34 VDD1.n10 0.155672
R226 VDD1.n27 VDD1.n10 0.155672
R227 VDD1.n27 VDD1.n26 0.155672
R228 VDD1.n26 VDD1.n14 0.155672
R229 VDD1.n19 VDD1.n14 0.155672
R230 VDD1.n71 VDD1.n66 0.155672
R231 VDD1.n78 VDD1.n66 0.155672
R232 VDD1.n79 VDD1.n78 0.155672
R233 VDD1.n79 VDD1.n62 0.155672
R234 VDD1.n86 VDD1.n62 0.155672
R235 VDD1.n87 VDD1.n86 0.155672
R236 VDD1.n87 VDD1.n58 0.155672
R237 VDD1.n96 VDD1.n58 0.155672
R238 VDD1.n97 VDD1.n96 0.155672
R239 VDD1.n97 VDD1.n54 0.155672
R240 VDD1.n104 VDD1.n54 0.155672
R241 VTAIL.n218 VTAIL.n170 289.615
R242 VTAIL.n50 VTAIL.n2 289.615
R243 VTAIL.n164 VTAIL.n116 289.615
R244 VTAIL.n108 VTAIL.n60 289.615
R245 VTAIL.n186 VTAIL.n185 185
R246 VTAIL.n191 VTAIL.n190 185
R247 VTAIL.n193 VTAIL.n192 185
R248 VTAIL.n182 VTAIL.n181 185
R249 VTAIL.n199 VTAIL.n198 185
R250 VTAIL.n201 VTAIL.n200 185
R251 VTAIL.n178 VTAIL.n177 185
R252 VTAIL.n208 VTAIL.n207 185
R253 VTAIL.n209 VTAIL.n176 185
R254 VTAIL.n211 VTAIL.n210 185
R255 VTAIL.n174 VTAIL.n173 185
R256 VTAIL.n217 VTAIL.n216 185
R257 VTAIL.n219 VTAIL.n218 185
R258 VTAIL.n18 VTAIL.n17 185
R259 VTAIL.n23 VTAIL.n22 185
R260 VTAIL.n25 VTAIL.n24 185
R261 VTAIL.n14 VTAIL.n13 185
R262 VTAIL.n31 VTAIL.n30 185
R263 VTAIL.n33 VTAIL.n32 185
R264 VTAIL.n10 VTAIL.n9 185
R265 VTAIL.n40 VTAIL.n39 185
R266 VTAIL.n41 VTAIL.n8 185
R267 VTAIL.n43 VTAIL.n42 185
R268 VTAIL.n6 VTAIL.n5 185
R269 VTAIL.n49 VTAIL.n48 185
R270 VTAIL.n51 VTAIL.n50 185
R271 VTAIL.n165 VTAIL.n164 185
R272 VTAIL.n163 VTAIL.n162 185
R273 VTAIL.n120 VTAIL.n119 185
R274 VTAIL.n157 VTAIL.n156 185
R275 VTAIL.n155 VTAIL.n122 185
R276 VTAIL.n154 VTAIL.n153 185
R277 VTAIL.n125 VTAIL.n123 185
R278 VTAIL.n148 VTAIL.n147 185
R279 VTAIL.n146 VTAIL.n145 185
R280 VTAIL.n129 VTAIL.n128 185
R281 VTAIL.n140 VTAIL.n139 185
R282 VTAIL.n138 VTAIL.n137 185
R283 VTAIL.n133 VTAIL.n132 185
R284 VTAIL.n109 VTAIL.n108 185
R285 VTAIL.n107 VTAIL.n106 185
R286 VTAIL.n64 VTAIL.n63 185
R287 VTAIL.n101 VTAIL.n100 185
R288 VTAIL.n99 VTAIL.n66 185
R289 VTAIL.n98 VTAIL.n97 185
R290 VTAIL.n69 VTAIL.n67 185
R291 VTAIL.n92 VTAIL.n91 185
R292 VTAIL.n90 VTAIL.n89 185
R293 VTAIL.n73 VTAIL.n72 185
R294 VTAIL.n84 VTAIL.n83 185
R295 VTAIL.n82 VTAIL.n81 185
R296 VTAIL.n77 VTAIL.n76 185
R297 VTAIL.n187 VTAIL.t4 149.524
R298 VTAIL.n19 VTAIL.t6 149.524
R299 VTAIL.n134 VTAIL.t10 149.524
R300 VTAIL.n78 VTAIL.t2 149.524
R301 VTAIL.n191 VTAIL.n185 104.615
R302 VTAIL.n192 VTAIL.n191 104.615
R303 VTAIL.n192 VTAIL.n181 104.615
R304 VTAIL.n199 VTAIL.n181 104.615
R305 VTAIL.n200 VTAIL.n199 104.615
R306 VTAIL.n200 VTAIL.n177 104.615
R307 VTAIL.n208 VTAIL.n177 104.615
R308 VTAIL.n209 VTAIL.n208 104.615
R309 VTAIL.n210 VTAIL.n209 104.615
R310 VTAIL.n210 VTAIL.n173 104.615
R311 VTAIL.n217 VTAIL.n173 104.615
R312 VTAIL.n218 VTAIL.n217 104.615
R313 VTAIL.n23 VTAIL.n17 104.615
R314 VTAIL.n24 VTAIL.n23 104.615
R315 VTAIL.n24 VTAIL.n13 104.615
R316 VTAIL.n31 VTAIL.n13 104.615
R317 VTAIL.n32 VTAIL.n31 104.615
R318 VTAIL.n32 VTAIL.n9 104.615
R319 VTAIL.n40 VTAIL.n9 104.615
R320 VTAIL.n41 VTAIL.n40 104.615
R321 VTAIL.n42 VTAIL.n41 104.615
R322 VTAIL.n42 VTAIL.n5 104.615
R323 VTAIL.n49 VTAIL.n5 104.615
R324 VTAIL.n50 VTAIL.n49 104.615
R325 VTAIL.n164 VTAIL.n163 104.615
R326 VTAIL.n163 VTAIL.n119 104.615
R327 VTAIL.n156 VTAIL.n119 104.615
R328 VTAIL.n156 VTAIL.n155 104.615
R329 VTAIL.n155 VTAIL.n154 104.615
R330 VTAIL.n154 VTAIL.n123 104.615
R331 VTAIL.n147 VTAIL.n123 104.615
R332 VTAIL.n147 VTAIL.n146 104.615
R333 VTAIL.n146 VTAIL.n128 104.615
R334 VTAIL.n139 VTAIL.n128 104.615
R335 VTAIL.n139 VTAIL.n138 104.615
R336 VTAIL.n138 VTAIL.n132 104.615
R337 VTAIL.n108 VTAIL.n107 104.615
R338 VTAIL.n107 VTAIL.n63 104.615
R339 VTAIL.n100 VTAIL.n63 104.615
R340 VTAIL.n100 VTAIL.n99 104.615
R341 VTAIL.n99 VTAIL.n98 104.615
R342 VTAIL.n98 VTAIL.n67 104.615
R343 VTAIL.n91 VTAIL.n67 104.615
R344 VTAIL.n91 VTAIL.n90 104.615
R345 VTAIL.n90 VTAIL.n72 104.615
R346 VTAIL.n83 VTAIL.n72 104.615
R347 VTAIL.n83 VTAIL.n82 104.615
R348 VTAIL.n82 VTAIL.n76 104.615
R349 VTAIL.t4 VTAIL.n185 52.3082
R350 VTAIL.t6 VTAIL.n17 52.3082
R351 VTAIL.t10 VTAIL.n132 52.3082
R352 VTAIL.t2 VTAIL.n76 52.3082
R353 VTAIL.n115 VTAIL.n114 50.4221
R354 VTAIL.n59 VTAIL.n58 50.4221
R355 VTAIL.n1 VTAIL.n0 50.422
R356 VTAIL.n57 VTAIL.n56 50.422
R357 VTAIL.n223 VTAIL.n222 36.646
R358 VTAIL.n55 VTAIL.n54 36.646
R359 VTAIL.n169 VTAIL.n168 36.646
R360 VTAIL.n113 VTAIL.n112 36.646
R361 VTAIL.n59 VTAIL.n57 26.0652
R362 VTAIL.n223 VTAIL.n169 23.6083
R363 VTAIL.n211 VTAIL.n176 13.1884
R364 VTAIL.n43 VTAIL.n8 13.1884
R365 VTAIL.n157 VTAIL.n122 13.1884
R366 VTAIL.n101 VTAIL.n66 13.1884
R367 VTAIL.n207 VTAIL.n206 12.8005
R368 VTAIL.n212 VTAIL.n174 12.8005
R369 VTAIL.n39 VTAIL.n38 12.8005
R370 VTAIL.n44 VTAIL.n6 12.8005
R371 VTAIL.n158 VTAIL.n120 12.8005
R372 VTAIL.n153 VTAIL.n124 12.8005
R373 VTAIL.n102 VTAIL.n64 12.8005
R374 VTAIL.n97 VTAIL.n68 12.8005
R375 VTAIL.n205 VTAIL.n178 12.0247
R376 VTAIL.n216 VTAIL.n215 12.0247
R377 VTAIL.n37 VTAIL.n10 12.0247
R378 VTAIL.n48 VTAIL.n47 12.0247
R379 VTAIL.n162 VTAIL.n161 12.0247
R380 VTAIL.n152 VTAIL.n125 12.0247
R381 VTAIL.n106 VTAIL.n105 12.0247
R382 VTAIL.n96 VTAIL.n69 12.0247
R383 VTAIL.n202 VTAIL.n201 11.249
R384 VTAIL.n219 VTAIL.n172 11.249
R385 VTAIL.n34 VTAIL.n33 11.249
R386 VTAIL.n51 VTAIL.n4 11.249
R387 VTAIL.n165 VTAIL.n118 11.249
R388 VTAIL.n149 VTAIL.n148 11.249
R389 VTAIL.n109 VTAIL.n62 11.249
R390 VTAIL.n93 VTAIL.n92 11.249
R391 VTAIL.n198 VTAIL.n180 10.4732
R392 VTAIL.n220 VTAIL.n170 10.4732
R393 VTAIL.n30 VTAIL.n12 10.4732
R394 VTAIL.n52 VTAIL.n2 10.4732
R395 VTAIL.n166 VTAIL.n116 10.4732
R396 VTAIL.n145 VTAIL.n127 10.4732
R397 VTAIL.n110 VTAIL.n60 10.4732
R398 VTAIL.n89 VTAIL.n71 10.4732
R399 VTAIL.n187 VTAIL.n186 10.2747
R400 VTAIL.n19 VTAIL.n18 10.2747
R401 VTAIL.n134 VTAIL.n133 10.2747
R402 VTAIL.n78 VTAIL.n77 10.2747
R403 VTAIL.n197 VTAIL.n182 9.69747
R404 VTAIL.n29 VTAIL.n14 9.69747
R405 VTAIL.n144 VTAIL.n129 9.69747
R406 VTAIL.n88 VTAIL.n73 9.69747
R407 VTAIL.n222 VTAIL.n221 9.45567
R408 VTAIL.n54 VTAIL.n53 9.45567
R409 VTAIL.n168 VTAIL.n167 9.45567
R410 VTAIL.n112 VTAIL.n111 9.45567
R411 VTAIL.n221 VTAIL.n220 9.3005
R412 VTAIL.n172 VTAIL.n171 9.3005
R413 VTAIL.n215 VTAIL.n214 9.3005
R414 VTAIL.n213 VTAIL.n212 9.3005
R415 VTAIL.n189 VTAIL.n188 9.3005
R416 VTAIL.n184 VTAIL.n183 9.3005
R417 VTAIL.n195 VTAIL.n194 9.3005
R418 VTAIL.n197 VTAIL.n196 9.3005
R419 VTAIL.n180 VTAIL.n179 9.3005
R420 VTAIL.n203 VTAIL.n202 9.3005
R421 VTAIL.n205 VTAIL.n204 9.3005
R422 VTAIL.n206 VTAIL.n175 9.3005
R423 VTAIL.n53 VTAIL.n52 9.3005
R424 VTAIL.n4 VTAIL.n3 9.3005
R425 VTAIL.n47 VTAIL.n46 9.3005
R426 VTAIL.n45 VTAIL.n44 9.3005
R427 VTAIL.n21 VTAIL.n20 9.3005
R428 VTAIL.n16 VTAIL.n15 9.3005
R429 VTAIL.n27 VTAIL.n26 9.3005
R430 VTAIL.n29 VTAIL.n28 9.3005
R431 VTAIL.n12 VTAIL.n11 9.3005
R432 VTAIL.n35 VTAIL.n34 9.3005
R433 VTAIL.n37 VTAIL.n36 9.3005
R434 VTAIL.n38 VTAIL.n7 9.3005
R435 VTAIL.n136 VTAIL.n135 9.3005
R436 VTAIL.n131 VTAIL.n130 9.3005
R437 VTAIL.n142 VTAIL.n141 9.3005
R438 VTAIL.n144 VTAIL.n143 9.3005
R439 VTAIL.n127 VTAIL.n126 9.3005
R440 VTAIL.n150 VTAIL.n149 9.3005
R441 VTAIL.n152 VTAIL.n151 9.3005
R442 VTAIL.n124 VTAIL.n121 9.3005
R443 VTAIL.n167 VTAIL.n166 9.3005
R444 VTAIL.n118 VTAIL.n117 9.3005
R445 VTAIL.n161 VTAIL.n160 9.3005
R446 VTAIL.n159 VTAIL.n158 9.3005
R447 VTAIL.n80 VTAIL.n79 9.3005
R448 VTAIL.n75 VTAIL.n74 9.3005
R449 VTAIL.n86 VTAIL.n85 9.3005
R450 VTAIL.n88 VTAIL.n87 9.3005
R451 VTAIL.n71 VTAIL.n70 9.3005
R452 VTAIL.n94 VTAIL.n93 9.3005
R453 VTAIL.n96 VTAIL.n95 9.3005
R454 VTAIL.n68 VTAIL.n65 9.3005
R455 VTAIL.n111 VTAIL.n110 9.3005
R456 VTAIL.n62 VTAIL.n61 9.3005
R457 VTAIL.n105 VTAIL.n104 9.3005
R458 VTAIL.n103 VTAIL.n102 9.3005
R459 VTAIL.n194 VTAIL.n193 8.92171
R460 VTAIL.n26 VTAIL.n25 8.92171
R461 VTAIL.n141 VTAIL.n140 8.92171
R462 VTAIL.n85 VTAIL.n84 8.92171
R463 VTAIL.n190 VTAIL.n184 8.14595
R464 VTAIL.n22 VTAIL.n16 8.14595
R465 VTAIL.n137 VTAIL.n131 8.14595
R466 VTAIL.n81 VTAIL.n75 8.14595
R467 VTAIL.n189 VTAIL.n186 7.3702
R468 VTAIL.n21 VTAIL.n18 7.3702
R469 VTAIL.n136 VTAIL.n133 7.3702
R470 VTAIL.n80 VTAIL.n77 7.3702
R471 VTAIL.n190 VTAIL.n189 5.81868
R472 VTAIL.n22 VTAIL.n21 5.81868
R473 VTAIL.n137 VTAIL.n136 5.81868
R474 VTAIL.n81 VTAIL.n80 5.81868
R475 VTAIL.n193 VTAIL.n184 5.04292
R476 VTAIL.n25 VTAIL.n16 5.04292
R477 VTAIL.n140 VTAIL.n131 5.04292
R478 VTAIL.n84 VTAIL.n75 5.04292
R479 VTAIL.n194 VTAIL.n182 4.26717
R480 VTAIL.n26 VTAIL.n14 4.26717
R481 VTAIL.n141 VTAIL.n129 4.26717
R482 VTAIL.n85 VTAIL.n73 4.26717
R483 VTAIL.n198 VTAIL.n197 3.49141
R484 VTAIL.n222 VTAIL.n170 3.49141
R485 VTAIL.n30 VTAIL.n29 3.49141
R486 VTAIL.n54 VTAIL.n2 3.49141
R487 VTAIL.n168 VTAIL.n116 3.49141
R488 VTAIL.n145 VTAIL.n144 3.49141
R489 VTAIL.n112 VTAIL.n60 3.49141
R490 VTAIL.n89 VTAIL.n88 3.49141
R491 VTAIL.n188 VTAIL.n187 2.84303
R492 VTAIL.n20 VTAIL.n19 2.84303
R493 VTAIL.n135 VTAIL.n134 2.84303
R494 VTAIL.n79 VTAIL.n78 2.84303
R495 VTAIL.n201 VTAIL.n180 2.71565
R496 VTAIL.n220 VTAIL.n219 2.71565
R497 VTAIL.n33 VTAIL.n12 2.71565
R498 VTAIL.n52 VTAIL.n51 2.71565
R499 VTAIL.n166 VTAIL.n165 2.71565
R500 VTAIL.n148 VTAIL.n127 2.71565
R501 VTAIL.n110 VTAIL.n109 2.71565
R502 VTAIL.n92 VTAIL.n71 2.71565
R503 VTAIL.n113 VTAIL.n59 2.4574
R504 VTAIL.n169 VTAIL.n115 2.4574
R505 VTAIL.n57 VTAIL.n55 2.4574
R506 VTAIL.n0 VTAIL.t5 1.94358
R507 VTAIL.n0 VTAIL.t0 1.94358
R508 VTAIL.n56 VTAIL.t7 1.94358
R509 VTAIL.n56 VTAIL.t11 1.94358
R510 VTAIL.n114 VTAIL.t8 1.94358
R511 VTAIL.n114 VTAIL.t9 1.94358
R512 VTAIL.n58 VTAIL.t1 1.94358
R513 VTAIL.n58 VTAIL.t3 1.94358
R514 VTAIL.n202 VTAIL.n178 1.93989
R515 VTAIL.n216 VTAIL.n172 1.93989
R516 VTAIL.n34 VTAIL.n10 1.93989
R517 VTAIL.n48 VTAIL.n4 1.93989
R518 VTAIL.n162 VTAIL.n118 1.93989
R519 VTAIL.n149 VTAIL.n125 1.93989
R520 VTAIL.n106 VTAIL.n62 1.93989
R521 VTAIL.n93 VTAIL.n69 1.93989
R522 VTAIL VTAIL.n223 1.78498
R523 VTAIL.n115 VTAIL.n113 1.69878
R524 VTAIL.n55 VTAIL.n1 1.69878
R525 VTAIL.n207 VTAIL.n205 1.16414
R526 VTAIL.n215 VTAIL.n174 1.16414
R527 VTAIL.n39 VTAIL.n37 1.16414
R528 VTAIL.n47 VTAIL.n6 1.16414
R529 VTAIL.n161 VTAIL.n120 1.16414
R530 VTAIL.n153 VTAIL.n152 1.16414
R531 VTAIL.n105 VTAIL.n64 1.16414
R532 VTAIL.n97 VTAIL.n96 1.16414
R533 VTAIL VTAIL.n1 0.672914
R534 VTAIL.n206 VTAIL.n176 0.388379
R535 VTAIL.n212 VTAIL.n211 0.388379
R536 VTAIL.n38 VTAIL.n8 0.388379
R537 VTAIL.n44 VTAIL.n43 0.388379
R538 VTAIL.n158 VTAIL.n157 0.388379
R539 VTAIL.n124 VTAIL.n122 0.388379
R540 VTAIL.n102 VTAIL.n101 0.388379
R541 VTAIL.n68 VTAIL.n66 0.388379
R542 VTAIL.n188 VTAIL.n183 0.155672
R543 VTAIL.n195 VTAIL.n183 0.155672
R544 VTAIL.n196 VTAIL.n195 0.155672
R545 VTAIL.n196 VTAIL.n179 0.155672
R546 VTAIL.n203 VTAIL.n179 0.155672
R547 VTAIL.n204 VTAIL.n203 0.155672
R548 VTAIL.n204 VTAIL.n175 0.155672
R549 VTAIL.n213 VTAIL.n175 0.155672
R550 VTAIL.n214 VTAIL.n213 0.155672
R551 VTAIL.n214 VTAIL.n171 0.155672
R552 VTAIL.n221 VTAIL.n171 0.155672
R553 VTAIL.n20 VTAIL.n15 0.155672
R554 VTAIL.n27 VTAIL.n15 0.155672
R555 VTAIL.n28 VTAIL.n27 0.155672
R556 VTAIL.n28 VTAIL.n11 0.155672
R557 VTAIL.n35 VTAIL.n11 0.155672
R558 VTAIL.n36 VTAIL.n35 0.155672
R559 VTAIL.n36 VTAIL.n7 0.155672
R560 VTAIL.n45 VTAIL.n7 0.155672
R561 VTAIL.n46 VTAIL.n45 0.155672
R562 VTAIL.n46 VTAIL.n3 0.155672
R563 VTAIL.n53 VTAIL.n3 0.155672
R564 VTAIL.n167 VTAIL.n117 0.155672
R565 VTAIL.n160 VTAIL.n117 0.155672
R566 VTAIL.n160 VTAIL.n159 0.155672
R567 VTAIL.n159 VTAIL.n121 0.155672
R568 VTAIL.n151 VTAIL.n121 0.155672
R569 VTAIL.n151 VTAIL.n150 0.155672
R570 VTAIL.n150 VTAIL.n126 0.155672
R571 VTAIL.n143 VTAIL.n126 0.155672
R572 VTAIL.n143 VTAIL.n142 0.155672
R573 VTAIL.n142 VTAIL.n130 0.155672
R574 VTAIL.n135 VTAIL.n130 0.155672
R575 VTAIL.n111 VTAIL.n61 0.155672
R576 VTAIL.n104 VTAIL.n61 0.155672
R577 VTAIL.n104 VTAIL.n103 0.155672
R578 VTAIL.n103 VTAIL.n65 0.155672
R579 VTAIL.n95 VTAIL.n65 0.155672
R580 VTAIL.n95 VTAIL.n94 0.155672
R581 VTAIL.n94 VTAIL.n70 0.155672
R582 VTAIL.n87 VTAIL.n70 0.155672
R583 VTAIL.n87 VTAIL.n86 0.155672
R584 VTAIL.n86 VTAIL.n74 0.155672
R585 VTAIL.n79 VTAIL.n74 0.155672
R586 B.n754 B.n753 585
R587 B.n285 B.n118 585
R588 B.n284 B.n283 585
R589 B.n282 B.n281 585
R590 B.n280 B.n279 585
R591 B.n278 B.n277 585
R592 B.n276 B.n275 585
R593 B.n274 B.n273 585
R594 B.n272 B.n271 585
R595 B.n270 B.n269 585
R596 B.n268 B.n267 585
R597 B.n266 B.n265 585
R598 B.n264 B.n263 585
R599 B.n262 B.n261 585
R600 B.n260 B.n259 585
R601 B.n258 B.n257 585
R602 B.n256 B.n255 585
R603 B.n254 B.n253 585
R604 B.n252 B.n251 585
R605 B.n250 B.n249 585
R606 B.n248 B.n247 585
R607 B.n246 B.n245 585
R608 B.n244 B.n243 585
R609 B.n242 B.n241 585
R610 B.n240 B.n239 585
R611 B.n238 B.n237 585
R612 B.n236 B.n235 585
R613 B.n234 B.n233 585
R614 B.n232 B.n231 585
R615 B.n230 B.n229 585
R616 B.n228 B.n227 585
R617 B.n226 B.n225 585
R618 B.n224 B.n223 585
R619 B.n222 B.n221 585
R620 B.n220 B.n219 585
R621 B.n218 B.n217 585
R622 B.n216 B.n215 585
R623 B.n214 B.n213 585
R624 B.n212 B.n211 585
R625 B.n210 B.n209 585
R626 B.n208 B.n207 585
R627 B.n206 B.n205 585
R628 B.n204 B.n203 585
R629 B.n202 B.n201 585
R630 B.n200 B.n199 585
R631 B.n198 B.n197 585
R632 B.n196 B.n195 585
R633 B.n194 B.n193 585
R634 B.n192 B.n191 585
R635 B.n190 B.n189 585
R636 B.n188 B.n187 585
R637 B.n186 B.n185 585
R638 B.n184 B.n183 585
R639 B.n182 B.n181 585
R640 B.n180 B.n179 585
R641 B.n178 B.n177 585
R642 B.n176 B.n175 585
R643 B.n174 B.n173 585
R644 B.n172 B.n171 585
R645 B.n170 B.n169 585
R646 B.n168 B.n167 585
R647 B.n166 B.n165 585
R648 B.n164 B.n163 585
R649 B.n162 B.n161 585
R650 B.n160 B.n159 585
R651 B.n158 B.n157 585
R652 B.n156 B.n155 585
R653 B.n154 B.n153 585
R654 B.n152 B.n151 585
R655 B.n150 B.n149 585
R656 B.n148 B.n147 585
R657 B.n146 B.n145 585
R658 B.n144 B.n143 585
R659 B.n142 B.n141 585
R660 B.n140 B.n139 585
R661 B.n138 B.n137 585
R662 B.n136 B.n135 585
R663 B.n134 B.n133 585
R664 B.n132 B.n131 585
R665 B.n130 B.n129 585
R666 B.n128 B.n127 585
R667 B.n126 B.n125 585
R668 B.n752 B.n77 585
R669 B.n757 B.n77 585
R670 B.n751 B.n76 585
R671 B.n758 B.n76 585
R672 B.n750 B.n749 585
R673 B.n749 B.n72 585
R674 B.n748 B.n71 585
R675 B.n764 B.n71 585
R676 B.n747 B.n70 585
R677 B.n765 B.n70 585
R678 B.n746 B.n69 585
R679 B.n766 B.n69 585
R680 B.n745 B.n744 585
R681 B.n744 B.n65 585
R682 B.n743 B.n64 585
R683 B.n772 B.n64 585
R684 B.n742 B.n63 585
R685 B.n773 B.n63 585
R686 B.n741 B.n62 585
R687 B.n774 B.n62 585
R688 B.n740 B.n739 585
R689 B.n739 B.n58 585
R690 B.n738 B.n57 585
R691 B.n780 B.n57 585
R692 B.n737 B.n56 585
R693 B.n781 B.n56 585
R694 B.n736 B.n55 585
R695 B.n782 B.n55 585
R696 B.n735 B.n734 585
R697 B.n734 B.n51 585
R698 B.n733 B.n50 585
R699 B.n788 B.n50 585
R700 B.n732 B.n49 585
R701 B.n789 B.n49 585
R702 B.n731 B.n48 585
R703 B.n790 B.n48 585
R704 B.n730 B.n729 585
R705 B.n729 B.n47 585
R706 B.n728 B.n43 585
R707 B.n796 B.n43 585
R708 B.n727 B.n42 585
R709 B.n797 B.n42 585
R710 B.n726 B.n41 585
R711 B.n798 B.n41 585
R712 B.n725 B.n724 585
R713 B.n724 B.n37 585
R714 B.n723 B.n36 585
R715 B.n804 B.n36 585
R716 B.n722 B.n35 585
R717 B.n805 B.n35 585
R718 B.n721 B.n34 585
R719 B.n806 B.n34 585
R720 B.n720 B.n719 585
R721 B.n719 B.n30 585
R722 B.n718 B.n29 585
R723 B.n812 B.n29 585
R724 B.n717 B.n28 585
R725 B.n813 B.n28 585
R726 B.n716 B.n27 585
R727 B.n814 B.n27 585
R728 B.n715 B.n714 585
R729 B.n714 B.n23 585
R730 B.n713 B.n22 585
R731 B.n820 B.n22 585
R732 B.n712 B.n21 585
R733 B.n821 B.n21 585
R734 B.n711 B.n20 585
R735 B.n822 B.n20 585
R736 B.n710 B.n709 585
R737 B.n709 B.n16 585
R738 B.n708 B.n15 585
R739 B.n828 B.n15 585
R740 B.n707 B.n14 585
R741 B.n829 B.n14 585
R742 B.n706 B.n13 585
R743 B.n830 B.n13 585
R744 B.n705 B.n704 585
R745 B.n704 B.n12 585
R746 B.n703 B.n702 585
R747 B.n703 B.n8 585
R748 B.n701 B.n7 585
R749 B.n837 B.n7 585
R750 B.n700 B.n6 585
R751 B.n838 B.n6 585
R752 B.n699 B.n5 585
R753 B.n839 B.n5 585
R754 B.n698 B.n697 585
R755 B.n697 B.n4 585
R756 B.n696 B.n286 585
R757 B.n696 B.n695 585
R758 B.n686 B.n287 585
R759 B.n288 B.n287 585
R760 B.n688 B.n687 585
R761 B.n689 B.n688 585
R762 B.n685 B.n293 585
R763 B.n293 B.n292 585
R764 B.n684 B.n683 585
R765 B.n683 B.n682 585
R766 B.n295 B.n294 585
R767 B.n296 B.n295 585
R768 B.n675 B.n674 585
R769 B.n676 B.n675 585
R770 B.n673 B.n301 585
R771 B.n301 B.n300 585
R772 B.n672 B.n671 585
R773 B.n671 B.n670 585
R774 B.n303 B.n302 585
R775 B.n304 B.n303 585
R776 B.n663 B.n662 585
R777 B.n664 B.n663 585
R778 B.n661 B.n309 585
R779 B.n309 B.n308 585
R780 B.n660 B.n659 585
R781 B.n659 B.n658 585
R782 B.n311 B.n310 585
R783 B.n312 B.n311 585
R784 B.n651 B.n650 585
R785 B.n652 B.n651 585
R786 B.n649 B.n317 585
R787 B.n317 B.n316 585
R788 B.n648 B.n647 585
R789 B.n647 B.n646 585
R790 B.n319 B.n318 585
R791 B.n320 B.n319 585
R792 B.n639 B.n638 585
R793 B.n640 B.n639 585
R794 B.n637 B.n325 585
R795 B.n325 B.n324 585
R796 B.n636 B.n635 585
R797 B.n635 B.n634 585
R798 B.n327 B.n326 585
R799 B.n627 B.n327 585
R800 B.n626 B.n625 585
R801 B.n628 B.n626 585
R802 B.n624 B.n332 585
R803 B.n332 B.n331 585
R804 B.n623 B.n622 585
R805 B.n622 B.n621 585
R806 B.n334 B.n333 585
R807 B.n335 B.n334 585
R808 B.n614 B.n613 585
R809 B.n615 B.n614 585
R810 B.n612 B.n340 585
R811 B.n340 B.n339 585
R812 B.n611 B.n610 585
R813 B.n610 B.n609 585
R814 B.n342 B.n341 585
R815 B.n343 B.n342 585
R816 B.n602 B.n601 585
R817 B.n603 B.n602 585
R818 B.n600 B.n348 585
R819 B.n348 B.n347 585
R820 B.n599 B.n598 585
R821 B.n598 B.n597 585
R822 B.n350 B.n349 585
R823 B.n351 B.n350 585
R824 B.n590 B.n589 585
R825 B.n591 B.n590 585
R826 B.n588 B.n356 585
R827 B.n356 B.n355 585
R828 B.n587 B.n586 585
R829 B.n586 B.n585 585
R830 B.n358 B.n357 585
R831 B.n359 B.n358 585
R832 B.n578 B.n577 585
R833 B.n579 B.n578 585
R834 B.n576 B.n364 585
R835 B.n364 B.n363 585
R836 B.n571 B.n570 585
R837 B.n569 B.n407 585
R838 B.n568 B.n406 585
R839 B.n573 B.n406 585
R840 B.n567 B.n566 585
R841 B.n565 B.n564 585
R842 B.n563 B.n562 585
R843 B.n561 B.n560 585
R844 B.n559 B.n558 585
R845 B.n557 B.n556 585
R846 B.n555 B.n554 585
R847 B.n553 B.n552 585
R848 B.n551 B.n550 585
R849 B.n549 B.n548 585
R850 B.n547 B.n546 585
R851 B.n545 B.n544 585
R852 B.n543 B.n542 585
R853 B.n541 B.n540 585
R854 B.n539 B.n538 585
R855 B.n537 B.n536 585
R856 B.n535 B.n534 585
R857 B.n533 B.n532 585
R858 B.n531 B.n530 585
R859 B.n529 B.n528 585
R860 B.n527 B.n526 585
R861 B.n525 B.n524 585
R862 B.n523 B.n522 585
R863 B.n521 B.n520 585
R864 B.n519 B.n518 585
R865 B.n517 B.n516 585
R866 B.n515 B.n514 585
R867 B.n513 B.n512 585
R868 B.n511 B.n510 585
R869 B.n509 B.n508 585
R870 B.n507 B.n506 585
R871 B.n505 B.n504 585
R872 B.n503 B.n502 585
R873 B.n500 B.n499 585
R874 B.n498 B.n497 585
R875 B.n496 B.n495 585
R876 B.n494 B.n493 585
R877 B.n492 B.n491 585
R878 B.n490 B.n489 585
R879 B.n488 B.n487 585
R880 B.n486 B.n485 585
R881 B.n484 B.n483 585
R882 B.n482 B.n481 585
R883 B.n479 B.n478 585
R884 B.n477 B.n476 585
R885 B.n475 B.n474 585
R886 B.n473 B.n472 585
R887 B.n471 B.n470 585
R888 B.n469 B.n468 585
R889 B.n467 B.n466 585
R890 B.n465 B.n464 585
R891 B.n463 B.n462 585
R892 B.n461 B.n460 585
R893 B.n459 B.n458 585
R894 B.n457 B.n456 585
R895 B.n455 B.n454 585
R896 B.n453 B.n452 585
R897 B.n451 B.n450 585
R898 B.n449 B.n448 585
R899 B.n447 B.n446 585
R900 B.n445 B.n444 585
R901 B.n443 B.n442 585
R902 B.n441 B.n440 585
R903 B.n439 B.n438 585
R904 B.n437 B.n436 585
R905 B.n435 B.n434 585
R906 B.n433 B.n432 585
R907 B.n431 B.n430 585
R908 B.n429 B.n428 585
R909 B.n427 B.n426 585
R910 B.n425 B.n424 585
R911 B.n423 B.n422 585
R912 B.n421 B.n420 585
R913 B.n419 B.n418 585
R914 B.n417 B.n416 585
R915 B.n415 B.n414 585
R916 B.n413 B.n412 585
R917 B.n366 B.n365 585
R918 B.n575 B.n574 585
R919 B.n574 B.n573 585
R920 B.n362 B.n361 585
R921 B.n363 B.n362 585
R922 B.n581 B.n580 585
R923 B.n580 B.n579 585
R924 B.n582 B.n360 585
R925 B.n360 B.n359 585
R926 B.n584 B.n583 585
R927 B.n585 B.n584 585
R928 B.n354 B.n353 585
R929 B.n355 B.n354 585
R930 B.n593 B.n592 585
R931 B.n592 B.n591 585
R932 B.n594 B.n352 585
R933 B.n352 B.n351 585
R934 B.n596 B.n595 585
R935 B.n597 B.n596 585
R936 B.n346 B.n345 585
R937 B.n347 B.n346 585
R938 B.n605 B.n604 585
R939 B.n604 B.n603 585
R940 B.n606 B.n344 585
R941 B.n344 B.n343 585
R942 B.n608 B.n607 585
R943 B.n609 B.n608 585
R944 B.n338 B.n337 585
R945 B.n339 B.n338 585
R946 B.n617 B.n616 585
R947 B.n616 B.n615 585
R948 B.n618 B.n336 585
R949 B.n336 B.n335 585
R950 B.n620 B.n619 585
R951 B.n621 B.n620 585
R952 B.n330 B.n329 585
R953 B.n331 B.n330 585
R954 B.n630 B.n629 585
R955 B.n629 B.n628 585
R956 B.n631 B.n328 585
R957 B.n627 B.n328 585
R958 B.n633 B.n632 585
R959 B.n634 B.n633 585
R960 B.n323 B.n322 585
R961 B.n324 B.n323 585
R962 B.n642 B.n641 585
R963 B.n641 B.n640 585
R964 B.n643 B.n321 585
R965 B.n321 B.n320 585
R966 B.n645 B.n644 585
R967 B.n646 B.n645 585
R968 B.n315 B.n314 585
R969 B.n316 B.n315 585
R970 B.n654 B.n653 585
R971 B.n653 B.n652 585
R972 B.n655 B.n313 585
R973 B.n313 B.n312 585
R974 B.n657 B.n656 585
R975 B.n658 B.n657 585
R976 B.n307 B.n306 585
R977 B.n308 B.n307 585
R978 B.n666 B.n665 585
R979 B.n665 B.n664 585
R980 B.n667 B.n305 585
R981 B.n305 B.n304 585
R982 B.n669 B.n668 585
R983 B.n670 B.n669 585
R984 B.n299 B.n298 585
R985 B.n300 B.n299 585
R986 B.n678 B.n677 585
R987 B.n677 B.n676 585
R988 B.n679 B.n297 585
R989 B.n297 B.n296 585
R990 B.n681 B.n680 585
R991 B.n682 B.n681 585
R992 B.n291 B.n290 585
R993 B.n292 B.n291 585
R994 B.n691 B.n690 585
R995 B.n690 B.n689 585
R996 B.n692 B.n289 585
R997 B.n289 B.n288 585
R998 B.n694 B.n693 585
R999 B.n695 B.n694 585
R1000 B.n3 B.n0 585
R1001 B.n4 B.n3 585
R1002 B.n836 B.n1 585
R1003 B.n837 B.n836 585
R1004 B.n835 B.n834 585
R1005 B.n835 B.n8 585
R1006 B.n833 B.n9 585
R1007 B.n12 B.n9 585
R1008 B.n832 B.n831 585
R1009 B.n831 B.n830 585
R1010 B.n11 B.n10 585
R1011 B.n829 B.n11 585
R1012 B.n827 B.n826 585
R1013 B.n828 B.n827 585
R1014 B.n825 B.n17 585
R1015 B.n17 B.n16 585
R1016 B.n824 B.n823 585
R1017 B.n823 B.n822 585
R1018 B.n19 B.n18 585
R1019 B.n821 B.n19 585
R1020 B.n819 B.n818 585
R1021 B.n820 B.n819 585
R1022 B.n817 B.n24 585
R1023 B.n24 B.n23 585
R1024 B.n816 B.n815 585
R1025 B.n815 B.n814 585
R1026 B.n26 B.n25 585
R1027 B.n813 B.n26 585
R1028 B.n811 B.n810 585
R1029 B.n812 B.n811 585
R1030 B.n809 B.n31 585
R1031 B.n31 B.n30 585
R1032 B.n808 B.n807 585
R1033 B.n807 B.n806 585
R1034 B.n33 B.n32 585
R1035 B.n805 B.n33 585
R1036 B.n803 B.n802 585
R1037 B.n804 B.n803 585
R1038 B.n801 B.n38 585
R1039 B.n38 B.n37 585
R1040 B.n800 B.n799 585
R1041 B.n799 B.n798 585
R1042 B.n40 B.n39 585
R1043 B.n797 B.n40 585
R1044 B.n795 B.n794 585
R1045 B.n796 B.n795 585
R1046 B.n793 B.n44 585
R1047 B.n47 B.n44 585
R1048 B.n792 B.n791 585
R1049 B.n791 B.n790 585
R1050 B.n46 B.n45 585
R1051 B.n789 B.n46 585
R1052 B.n787 B.n786 585
R1053 B.n788 B.n787 585
R1054 B.n785 B.n52 585
R1055 B.n52 B.n51 585
R1056 B.n784 B.n783 585
R1057 B.n783 B.n782 585
R1058 B.n54 B.n53 585
R1059 B.n781 B.n54 585
R1060 B.n779 B.n778 585
R1061 B.n780 B.n779 585
R1062 B.n777 B.n59 585
R1063 B.n59 B.n58 585
R1064 B.n776 B.n775 585
R1065 B.n775 B.n774 585
R1066 B.n61 B.n60 585
R1067 B.n773 B.n61 585
R1068 B.n771 B.n770 585
R1069 B.n772 B.n771 585
R1070 B.n769 B.n66 585
R1071 B.n66 B.n65 585
R1072 B.n768 B.n767 585
R1073 B.n767 B.n766 585
R1074 B.n68 B.n67 585
R1075 B.n765 B.n68 585
R1076 B.n763 B.n762 585
R1077 B.n764 B.n763 585
R1078 B.n761 B.n73 585
R1079 B.n73 B.n72 585
R1080 B.n760 B.n759 585
R1081 B.n759 B.n758 585
R1082 B.n75 B.n74 585
R1083 B.n757 B.n75 585
R1084 B.n840 B.n839 585
R1085 B.n838 B.n2 585
R1086 B.n125 B.n75 535.745
R1087 B.n754 B.n77 535.745
R1088 B.n574 B.n364 535.745
R1089 B.n571 B.n362 535.745
R1090 B.n119 B.t15 306.604
R1091 B.n410 B.t9 306.604
R1092 B.n122 B.t18 306.604
R1093 B.n408 B.t12 306.604
R1094 B.n122 B.t17 305.375
R1095 B.n119 B.t13 305.375
R1096 B.n410 B.t6 305.375
R1097 B.n408 B.t10 305.375
R1098 B.n756 B.n755 256.663
R1099 B.n756 B.n117 256.663
R1100 B.n756 B.n116 256.663
R1101 B.n756 B.n115 256.663
R1102 B.n756 B.n114 256.663
R1103 B.n756 B.n113 256.663
R1104 B.n756 B.n112 256.663
R1105 B.n756 B.n111 256.663
R1106 B.n756 B.n110 256.663
R1107 B.n756 B.n109 256.663
R1108 B.n756 B.n108 256.663
R1109 B.n756 B.n107 256.663
R1110 B.n756 B.n106 256.663
R1111 B.n756 B.n105 256.663
R1112 B.n756 B.n104 256.663
R1113 B.n756 B.n103 256.663
R1114 B.n756 B.n102 256.663
R1115 B.n756 B.n101 256.663
R1116 B.n756 B.n100 256.663
R1117 B.n756 B.n99 256.663
R1118 B.n756 B.n98 256.663
R1119 B.n756 B.n97 256.663
R1120 B.n756 B.n96 256.663
R1121 B.n756 B.n95 256.663
R1122 B.n756 B.n94 256.663
R1123 B.n756 B.n93 256.663
R1124 B.n756 B.n92 256.663
R1125 B.n756 B.n91 256.663
R1126 B.n756 B.n90 256.663
R1127 B.n756 B.n89 256.663
R1128 B.n756 B.n88 256.663
R1129 B.n756 B.n87 256.663
R1130 B.n756 B.n86 256.663
R1131 B.n756 B.n85 256.663
R1132 B.n756 B.n84 256.663
R1133 B.n756 B.n83 256.663
R1134 B.n756 B.n82 256.663
R1135 B.n756 B.n81 256.663
R1136 B.n756 B.n80 256.663
R1137 B.n756 B.n79 256.663
R1138 B.n756 B.n78 256.663
R1139 B.n573 B.n572 256.663
R1140 B.n573 B.n367 256.663
R1141 B.n573 B.n368 256.663
R1142 B.n573 B.n369 256.663
R1143 B.n573 B.n370 256.663
R1144 B.n573 B.n371 256.663
R1145 B.n573 B.n372 256.663
R1146 B.n573 B.n373 256.663
R1147 B.n573 B.n374 256.663
R1148 B.n573 B.n375 256.663
R1149 B.n573 B.n376 256.663
R1150 B.n573 B.n377 256.663
R1151 B.n573 B.n378 256.663
R1152 B.n573 B.n379 256.663
R1153 B.n573 B.n380 256.663
R1154 B.n573 B.n381 256.663
R1155 B.n573 B.n382 256.663
R1156 B.n573 B.n383 256.663
R1157 B.n573 B.n384 256.663
R1158 B.n573 B.n385 256.663
R1159 B.n573 B.n386 256.663
R1160 B.n573 B.n387 256.663
R1161 B.n573 B.n388 256.663
R1162 B.n573 B.n389 256.663
R1163 B.n573 B.n390 256.663
R1164 B.n573 B.n391 256.663
R1165 B.n573 B.n392 256.663
R1166 B.n573 B.n393 256.663
R1167 B.n573 B.n394 256.663
R1168 B.n573 B.n395 256.663
R1169 B.n573 B.n396 256.663
R1170 B.n573 B.n397 256.663
R1171 B.n573 B.n398 256.663
R1172 B.n573 B.n399 256.663
R1173 B.n573 B.n400 256.663
R1174 B.n573 B.n401 256.663
R1175 B.n573 B.n402 256.663
R1176 B.n573 B.n403 256.663
R1177 B.n573 B.n404 256.663
R1178 B.n573 B.n405 256.663
R1179 B.n842 B.n841 256.663
R1180 B.n120 B.t16 251.333
R1181 B.n411 B.t8 251.333
R1182 B.n123 B.t19 251.332
R1183 B.n409 B.t11 251.332
R1184 B.n129 B.n128 163.367
R1185 B.n133 B.n132 163.367
R1186 B.n137 B.n136 163.367
R1187 B.n141 B.n140 163.367
R1188 B.n145 B.n144 163.367
R1189 B.n149 B.n148 163.367
R1190 B.n153 B.n152 163.367
R1191 B.n157 B.n156 163.367
R1192 B.n161 B.n160 163.367
R1193 B.n165 B.n164 163.367
R1194 B.n169 B.n168 163.367
R1195 B.n173 B.n172 163.367
R1196 B.n177 B.n176 163.367
R1197 B.n181 B.n180 163.367
R1198 B.n185 B.n184 163.367
R1199 B.n189 B.n188 163.367
R1200 B.n193 B.n192 163.367
R1201 B.n197 B.n196 163.367
R1202 B.n201 B.n200 163.367
R1203 B.n205 B.n204 163.367
R1204 B.n209 B.n208 163.367
R1205 B.n213 B.n212 163.367
R1206 B.n217 B.n216 163.367
R1207 B.n221 B.n220 163.367
R1208 B.n225 B.n224 163.367
R1209 B.n229 B.n228 163.367
R1210 B.n233 B.n232 163.367
R1211 B.n237 B.n236 163.367
R1212 B.n241 B.n240 163.367
R1213 B.n245 B.n244 163.367
R1214 B.n249 B.n248 163.367
R1215 B.n253 B.n252 163.367
R1216 B.n257 B.n256 163.367
R1217 B.n261 B.n260 163.367
R1218 B.n265 B.n264 163.367
R1219 B.n269 B.n268 163.367
R1220 B.n273 B.n272 163.367
R1221 B.n277 B.n276 163.367
R1222 B.n281 B.n280 163.367
R1223 B.n283 B.n118 163.367
R1224 B.n578 B.n364 163.367
R1225 B.n578 B.n358 163.367
R1226 B.n586 B.n358 163.367
R1227 B.n586 B.n356 163.367
R1228 B.n590 B.n356 163.367
R1229 B.n590 B.n350 163.367
R1230 B.n598 B.n350 163.367
R1231 B.n598 B.n348 163.367
R1232 B.n602 B.n348 163.367
R1233 B.n602 B.n342 163.367
R1234 B.n610 B.n342 163.367
R1235 B.n610 B.n340 163.367
R1236 B.n614 B.n340 163.367
R1237 B.n614 B.n334 163.367
R1238 B.n622 B.n334 163.367
R1239 B.n622 B.n332 163.367
R1240 B.n626 B.n332 163.367
R1241 B.n626 B.n327 163.367
R1242 B.n635 B.n327 163.367
R1243 B.n635 B.n325 163.367
R1244 B.n639 B.n325 163.367
R1245 B.n639 B.n319 163.367
R1246 B.n647 B.n319 163.367
R1247 B.n647 B.n317 163.367
R1248 B.n651 B.n317 163.367
R1249 B.n651 B.n311 163.367
R1250 B.n659 B.n311 163.367
R1251 B.n659 B.n309 163.367
R1252 B.n663 B.n309 163.367
R1253 B.n663 B.n303 163.367
R1254 B.n671 B.n303 163.367
R1255 B.n671 B.n301 163.367
R1256 B.n675 B.n301 163.367
R1257 B.n675 B.n295 163.367
R1258 B.n683 B.n295 163.367
R1259 B.n683 B.n293 163.367
R1260 B.n688 B.n293 163.367
R1261 B.n688 B.n287 163.367
R1262 B.n696 B.n287 163.367
R1263 B.n697 B.n696 163.367
R1264 B.n697 B.n5 163.367
R1265 B.n6 B.n5 163.367
R1266 B.n7 B.n6 163.367
R1267 B.n703 B.n7 163.367
R1268 B.n704 B.n703 163.367
R1269 B.n704 B.n13 163.367
R1270 B.n14 B.n13 163.367
R1271 B.n15 B.n14 163.367
R1272 B.n709 B.n15 163.367
R1273 B.n709 B.n20 163.367
R1274 B.n21 B.n20 163.367
R1275 B.n22 B.n21 163.367
R1276 B.n714 B.n22 163.367
R1277 B.n714 B.n27 163.367
R1278 B.n28 B.n27 163.367
R1279 B.n29 B.n28 163.367
R1280 B.n719 B.n29 163.367
R1281 B.n719 B.n34 163.367
R1282 B.n35 B.n34 163.367
R1283 B.n36 B.n35 163.367
R1284 B.n724 B.n36 163.367
R1285 B.n724 B.n41 163.367
R1286 B.n42 B.n41 163.367
R1287 B.n43 B.n42 163.367
R1288 B.n729 B.n43 163.367
R1289 B.n729 B.n48 163.367
R1290 B.n49 B.n48 163.367
R1291 B.n50 B.n49 163.367
R1292 B.n734 B.n50 163.367
R1293 B.n734 B.n55 163.367
R1294 B.n56 B.n55 163.367
R1295 B.n57 B.n56 163.367
R1296 B.n739 B.n57 163.367
R1297 B.n739 B.n62 163.367
R1298 B.n63 B.n62 163.367
R1299 B.n64 B.n63 163.367
R1300 B.n744 B.n64 163.367
R1301 B.n744 B.n69 163.367
R1302 B.n70 B.n69 163.367
R1303 B.n71 B.n70 163.367
R1304 B.n749 B.n71 163.367
R1305 B.n749 B.n76 163.367
R1306 B.n77 B.n76 163.367
R1307 B.n407 B.n406 163.367
R1308 B.n566 B.n406 163.367
R1309 B.n564 B.n563 163.367
R1310 B.n560 B.n559 163.367
R1311 B.n556 B.n555 163.367
R1312 B.n552 B.n551 163.367
R1313 B.n548 B.n547 163.367
R1314 B.n544 B.n543 163.367
R1315 B.n540 B.n539 163.367
R1316 B.n536 B.n535 163.367
R1317 B.n532 B.n531 163.367
R1318 B.n528 B.n527 163.367
R1319 B.n524 B.n523 163.367
R1320 B.n520 B.n519 163.367
R1321 B.n516 B.n515 163.367
R1322 B.n512 B.n511 163.367
R1323 B.n508 B.n507 163.367
R1324 B.n504 B.n503 163.367
R1325 B.n499 B.n498 163.367
R1326 B.n495 B.n494 163.367
R1327 B.n491 B.n490 163.367
R1328 B.n487 B.n486 163.367
R1329 B.n483 B.n482 163.367
R1330 B.n478 B.n477 163.367
R1331 B.n474 B.n473 163.367
R1332 B.n470 B.n469 163.367
R1333 B.n466 B.n465 163.367
R1334 B.n462 B.n461 163.367
R1335 B.n458 B.n457 163.367
R1336 B.n454 B.n453 163.367
R1337 B.n450 B.n449 163.367
R1338 B.n446 B.n445 163.367
R1339 B.n442 B.n441 163.367
R1340 B.n438 B.n437 163.367
R1341 B.n434 B.n433 163.367
R1342 B.n430 B.n429 163.367
R1343 B.n426 B.n425 163.367
R1344 B.n422 B.n421 163.367
R1345 B.n418 B.n417 163.367
R1346 B.n414 B.n413 163.367
R1347 B.n574 B.n366 163.367
R1348 B.n580 B.n362 163.367
R1349 B.n580 B.n360 163.367
R1350 B.n584 B.n360 163.367
R1351 B.n584 B.n354 163.367
R1352 B.n592 B.n354 163.367
R1353 B.n592 B.n352 163.367
R1354 B.n596 B.n352 163.367
R1355 B.n596 B.n346 163.367
R1356 B.n604 B.n346 163.367
R1357 B.n604 B.n344 163.367
R1358 B.n608 B.n344 163.367
R1359 B.n608 B.n338 163.367
R1360 B.n616 B.n338 163.367
R1361 B.n616 B.n336 163.367
R1362 B.n620 B.n336 163.367
R1363 B.n620 B.n330 163.367
R1364 B.n629 B.n330 163.367
R1365 B.n629 B.n328 163.367
R1366 B.n633 B.n328 163.367
R1367 B.n633 B.n323 163.367
R1368 B.n641 B.n323 163.367
R1369 B.n641 B.n321 163.367
R1370 B.n645 B.n321 163.367
R1371 B.n645 B.n315 163.367
R1372 B.n653 B.n315 163.367
R1373 B.n653 B.n313 163.367
R1374 B.n657 B.n313 163.367
R1375 B.n657 B.n307 163.367
R1376 B.n665 B.n307 163.367
R1377 B.n665 B.n305 163.367
R1378 B.n669 B.n305 163.367
R1379 B.n669 B.n299 163.367
R1380 B.n677 B.n299 163.367
R1381 B.n677 B.n297 163.367
R1382 B.n681 B.n297 163.367
R1383 B.n681 B.n291 163.367
R1384 B.n690 B.n291 163.367
R1385 B.n690 B.n289 163.367
R1386 B.n694 B.n289 163.367
R1387 B.n694 B.n3 163.367
R1388 B.n840 B.n3 163.367
R1389 B.n836 B.n2 163.367
R1390 B.n836 B.n835 163.367
R1391 B.n835 B.n9 163.367
R1392 B.n831 B.n9 163.367
R1393 B.n831 B.n11 163.367
R1394 B.n827 B.n11 163.367
R1395 B.n827 B.n17 163.367
R1396 B.n823 B.n17 163.367
R1397 B.n823 B.n19 163.367
R1398 B.n819 B.n19 163.367
R1399 B.n819 B.n24 163.367
R1400 B.n815 B.n24 163.367
R1401 B.n815 B.n26 163.367
R1402 B.n811 B.n26 163.367
R1403 B.n811 B.n31 163.367
R1404 B.n807 B.n31 163.367
R1405 B.n807 B.n33 163.367
R1406 B.n803 B.n33 163.367
R1407 B.n803 B.n38 163.367
R1408 B.n799 B.n38 163.367
R1409 B.n799 B.n40 163.367
R1410 B.n795 B.n40 163.367
R1411 B.n795 B.n44 163.367
R1412 B.n791 B.n44 163.367
R1413 B.n791 B.n46 163.367
R1414 B.n787 B.n46 163.367
R1415 B.n787 B.n52 163.367
R1416 B.n783 B.n52 163.367
R1417 B.n783 B.n54 163.367
R1418 B.n779 B.n54 163.367
R1419 B.n779 B.n59 163.367
R1420 B.n775 B.n59 163.367
R1421 B.n775 B.n61 163.367
R1422 B.n771 B.n61 163.367
R1423 B.n771 B.n66 163.367
R1424 B.n767 B.n66 163.367
R1425 B.n767 B.n68 163.367
R1426 B.n763 B.n68 163.367
R1427 B.n763 B.n73 163.367
R1428 B.n759 B.n73 163.367
R1429 B.n759 B.n75 163.367
R1430 B.n573 B.n363 94.6012
R1431 B.n757 B.n756 94.6012
R1432 B.n125 B.n78 71.676
R1433 B.n129 B.n79 71.676
R1434 B.n133 B.n80 71.676
R1435 B.n137 B.n81 71.676
R1436 B.n141 B.n82 71.676
R1437 B.n145 B.n83 71.676
R1438 B.n149 B.n84 71.676
R1439 B.n153 B.n85 71.676
R1440 B.n157 B.n86 71.676
R1441 B.n161 B.n87 71.676
R1442 B.n165 B.n88 71.676
R1443 B.n169 B.n89 71.676
R1444 B.n173 B.n90 71.676
R1445 B.n177 B.n91 71.676
R1446 B.n181 B.n92 71.676
R1447 B.n185 B.n93 71.676
R1448 B.n189 B.n94 71.676
R1449 B.n193 B.n95 71.676
R1450 B.n197 B.n96 71.676
R1451 B.n201 B.n97 71.676
R1452 B.n205 B.n98 71.676
R1453 B.n209 B.n99 71.676
R1454 B.n213 B.n100 71.676
R1455 B.n217 B.n101 71.676
R1456 B.n221 B.n102 71.676
R1457 B.n225 B.n103 71.676
R1458 B.n229 B.n104 71.676
R1459 B.n233 B.n105 71.676
R1460 B.n237 B.n106 71.676
R1461 B.n241 B.n107 71.676
R1462 B.n245 B.n108 71.676
R1463 B.n249 B.n109 71.676
R1464 B.n253 B.n110 71.676
R1465 B.n257 B.n111 71.676
R1466 B.n261 B.n112 71.676
R1467 B.n265 B.n113 71.676
R1468 B.n269 B.n114 71.676
R1469 B.n273 B.n115 71.676
R1470 B.n277 B.n116 71.676
R1471 B.n281 B.n117 71.676
R1472 B.n755 B.n118 71.676
R1473 B.n755 B.n754 71.676
R1474 B.n283 B.n117 71.676
R1475 B.n280 B.n116 71.676
R1476 B.n276 B.n115 71.676
R1477 B.n272 B.n114 71.676
R1478 B.n268 B.n113 71.676
R1479 B.n264 B.n112 71.676
R1480 B.n260 B.n111 71.676
R1481 B.n256 B.n110 71.676
R1482 B.n252 B.n109 71.676
R1483 B.n248 B.n108 71.676
R1484 B.n244 B.n107 71.676
R1485 B.n240 B.n106 71.676
R1486 B.n236 B.n105 71.676
R1487 B.n232 B.n104 71.676
R1488 B.n228 B.n103 71.676
R1489 B.n224 B.n102 71.676
R1490 B.n220 B.n101 71.676
R1491 B.n216 B.n100 71.676
R1492 B.n212 B.n99 71.676
R1493 B.n208 B.n98 71.676
R1494 B.n204 B.n97 71.676
R1495 B.n200 B.n96 71.676
R1496 B.n196 B.n95 71.676
R1497 B.n192 B.n94 71.676
R1498 B.n188 B.n93 71.676
R1499 B.n184 B.n92 71.676
R1500 B.n180 B.n91 71.676
R1501 B.n176 B.n90 71.676
R1502 B.n172 B.n89 71.676
R1503 B.n168 B.n88 71.676
R1504 B.n164 B.n87 71.676
R1505 B.n160 B.n86 71.676
R1506 B.n156 B.n85 71.676
R1507 B.n152 B.n84 71.676
R1508 B.n148 B.n83 71.676
R1509 B.n144 B.n82 71.676
R1510 B.n140 B.n81 71.676
R1511 B.n136 B.n80 71.676
R1512 B.n132 B.n79 71.676
R1513 B.n128 B.n78 71.676
R1514 B.n572 B.n571 71.676
R1515 B.n566 B.n367 71.676
R1516 B.n563 B.n368 71.676
R1517 B.n559 B.n369 71.676
R1518 B.n555 B.n370 71.676
R1519 B.n551 B.n371 71.676
R1520 B.n547 B.n372 71.676
R1521 B.n543 B.n373 71.676
R1522 B.n539 B.n374 71.676
R1523 B.n535 B.n375 71.676
R1524 B.n531 B.n376 71.676
R1525 B.n527 B.n377 71.676
R1526 B.n523 B.n378 71.676
R1527 B.n519 B.n379 71.676
R1528 B.n515 B.n380 71.676
R1529 B.n511 B.n381 71.676
R1530 B.n507 B.n382 71.676
R1531 B.n503 B.n383 71.676
R1532 B.n498 B.n384 71.676
R1533 B.n494 B.n385 71.676
R1534 B.n490 B.n386 71.676
R1535 B.n486 B.n387 71.676
R1536 B.n482 B.n388 71.676
R1537 B.n477 B.n389 71.676
R1538 B.n473 B.n390 71.676
R1539 B.n469 B.n391 71.676
R1540 B.n465 B.n392 71.676
R1541 B.n461 B.n393 71.676
R1542 B.n457 B.n394 71.676
R1543 B.n453 B.n395 71.676
R1544 B.n449 B.n396 71.676
R1545 B.n445 B.n397 71.676
R1546 B.n441 B.n398 71.676
R1547 B.n437 B.n399 71.676
R1548 B.n433 B.n400 71.676
R1549 B.n429 B.n401 71.676
R1550 B.n425 B.n402 71.676
R1551 B.n421 B.n403 71.676
R1552 B.n417 B.n404 71.676
R1553 B.n413 B.n405 71.676
R1554 B.n572 B.n407 71.676
R1555 B.n564 B.n367 71.676
R1556 B.n560 B.n368 71.676
R1557 B.n556 B.n369 71.676
R1558 B.n552 B.n370 71.676
R1559 B.n548 B.n371 71.676
R1560 B.n544 B.n372 71.676
R1561 B.n540 B.n373 71.676
R1562 B.n536 B.n374 71.676
R1563 B.n532 B.n375 71.676
R1564 B.n528 B.n376 71.676
R1565 B.n524 B.n377 71.676
R1566 B.n520 B.n378 71.676
R1567 B.n516 B.n379 71.676
R1568 B.n512 B.n380 71.676
R1569 B.n508 B.n381 71.676
R1570 B.n504 B.n382 71.676
R1571 B.n499 B.n383 71.676
R1572 B.n495 B.n384 71.676
R1573 B.n491 B.n385 71.676
R1574 B.n487 B.n386 71.676
R1575 B.n483 B.n387 71.676
R1576 B.n478 B.n388 71.676
R1577 B.n474 B.n389 71.676
R1578 B.n470 B.n390 71.676
R1579 B.n466 B.n391 71.676
R1580 B.n462 B.n392 71.676
R1581 B.n458 B.n393 71.676
R1582 B.n454 B.n394 71.676
R1583 B.n450 B.n395 71.676
R1584 B.n446 B.n396 71.676
R1585 B.n442 B.n397 71.676
R1586 B.n438 B.n398 71.676
R1587 B.n434 B.n399 71.676
R1588 B.n430 B.n400 71.676
R1589 B.n426 B.n401 71.676
R1590 B.n422 B.n402 71.676
R1591 B.n418 B.n403 71.676
R1592 B.n414 B.n404 71.676
R1593 B.n405 B.n366 71.676
R1594 B.n841 B.n840 71.676
R1595 B.n841 B.n2 71.676
R1596 B.n124 B.n123 59.5399
R1597 B.n121 B.n120 59.5399
R1598 B.n480 B.n411 59.5399
R1599 B.n501 B.n409 59.5399
R1600 B.n123 B.n122 55.2732
R1601 B.n120 B.n119 55.2732
R1602 B.n411 B.n410 55.2732
R1603 B.n409 B.n408 55.2732
R1604 B.n579 B.n363 48.3678
R1605 B.n579 B.n359 48.3678
R1606 B.n585 B.n359 48.3678
R1607 B.n585 B.n355 48.3678
R1608 B.n591 B.n355 48.3678
R1609 B.n591 B.n351 48.3678
R1610 B.n597 B.n351 48.3678
R1611 B.n603 B.n347 48.3678
R1612 B.n603 B.n343 48.3678
R1613 B.n609 B.n343 48.3678
R1614 B.n609 B.n339 48.3678
R1615 B.n615 B.n339 48.3678
R1616 B.n615 B.n335 48.3678
R1617 B.n621 B.n335 48.3678
R1618 B.n621 B.n331 48.3678
R1619 B.n628 B.n331 48.3678
R1620 B.n628 B.n627 48.3678
R1621 B.n634 B.n324 48.3678
R1622 B.n640 B.n324 48.3678
R1623 B.n640 B.n320 48.3678
R1624 B.n646 B.n320 48.3678
R1625 B.n646 B.n316 48.3678
R1626 B.n652 B.n316 48.3678
R1627 B.n652 B.n312 48.3678
R1628 B.n658 B.n312 48.3678
R1629 B.n664 B.n308 48.3678
R1630 B.n664 B.n304 48.3678
R1631 B.n670 B.n304 48.3678
R1632 B.n670 B.n300 48.3678
R1633 B.n676 B.n300 48.3678
R1634 B.n676 B.n296 48.3678
R1635 B.n682 B.n296 48.3678
R1636 B.n689 B.n292 48.3678
R1637 B.n689 B.n288 48.3678
R1638 B.n695 B.n288 48.3678
R1639 B.n695 B.n4 48.3678
R1640 B.n839 B.n4 48.3678
R1641 B.n839 B.n838 48.3678
R1642 B.n838 B.n837 48.3678
R1643 B.n837 B.n8 48.3678
R1644 B.n12 B.n8 48.3678
R1645 B.n830 B.n12 48.3678
R1646 B.n830 B.n829 48.3678
R1647 B.n828 B.n16 48.3678
R1648 B.n822 B.n16 48.3678
R1649 B.n822 B.n821 48.3678
R1650 B.n821 B.n820 48.3678
R1651 B.n820 B.n23 48.3678
R1652 B.n814 B.n23 48.3678
R1653 B.n814 B.n813 48.3678
R1654 B.n812 B.n30 48.3678
R1655 B.n806 B.n30 48.3678
R1656 B.n806 B.n805 48.3678
R1657 B.n805 B.n804 48.3678
R1658 B.n804 B.n37 48.3678
R1659 B.n798 B.n37 48.3678
R1660 B.n798 B.n797 48.3678
R1661 B.n797 B.n796 48.3678
R1662 B.n790 B.n47 48.3678
R1663 B.n790 B.n789 48.3678
R1664 B.n789 B.n788 48.3678
R1665 B.n788 B.n51 48.3678
R1666 B.n782 B.n51 48.3678
R1667 B.n782 B.n781 48.3678
R1668 B.n781 B.n780 48.3678
R1669 B.n780 B.n58 48.3678
R1670 B.n774 B.n58 48.3678
R1671 B.n774 B.n773 48.3678
R1672 B.n772 B.n65 48.3678
R1673 B.n766 B.n65 48.3678
R1674 B.n766 B.n765 48.3678
R1675 B.n765 B.n764 48.3678
R1676 B.n764 B.n72 48.3678
R1677 B.n758 B.n72 48.3678
R1678 B.n758 B.n757 48.3678
R1679 B.n627 B.t1 45.5226
R1680 B.n47 B.t4 45.5226
R1681 B.n570 B.n361 34.8103
R1682 B.n576 B.n575 34.8103
R1683 B.n753 B.n752 34.8103
R1684 B.n126 B.n74 34.8103
R1685 B.n682 B.t2 34.1421
R1686 B.t5 B.n828 34.1421
R1687 B.t3 B.n308 32.7195
R1688 B.n813 B.t0 32.7195
R1689 B.t7 B.n347 31.297
R1690 B.n773 B.t14 31.297
R1691 B B.n842 18.0485
R1692 B.n597 B.t7 17.0713
R1693 B.t14 B.n772 17.0713
R1694 B.n658 B.t3 15.6487
R1695 B.t0 B.n812 15.6487
R1696 B.t2 B.n292 14.2262
R1697 B.n829 B.t5 14.2262
R1698 B.n581 B.n361 10.6151
R1699 B.n582 B.n581 10.6151
R1700 B.n583 B.n582 10.6151
R1701 B.n583 B.n353 10.6151
R1702 B.n593 B.n353 10.6151
R1703 B.n594 B.n593 10.6151
R1704 B.n595 B.n594 10.6151
R1705 B.n595 B.n345 10.6151
R1706 B.n605 B.n345 10.6151
R1707 B.n606 B.n605 10.6151
R1708 B.n607 B.n606 10.6151
R1709 B.n607 B.n337 10.6151
R1710 B.n617 B.n337 10.6151
R1711 B.n618 B.n617 10.6151
R1712 B.n619 B.n618 10.6151
R1713 B.n619 B.n329 10.6151
R1714 B.n630 B.n329 10.6151
R1715 B.n631 B.n630 10.6151
R1716 B.n632 B.n631 10.6151
R1717 B.n632 B.n322 10.6151
R1718 B.n642 B.n322 10.6151
R1719 B.n643 B.n642 10.6151
R1720 B.n644 B.n643 10.6151
R1721 B.n644 B.n314 10.6151
R1722 B.n654 B.n314 10.6151
R1723 B.n655 B.n654 10.6151
R1724 B.n656 B.n655 10.6151
R1725 B.n656 B.n306 10.6151
R1726 B.n666 B.n306 10.6151
R1727 B.n667 B.n666 10.6151
R1728 B.n668 B.n667 10.6151
R1729 B.n668 B.n298 10.6151
R1730 B.n678 B.n298 10.6151
R1731 B.n679 B.n678 10.6151
R1732 B.n680 B.n679 10.6151
R1733 B.n680 B.n290 10.6151
R1734 B.n691 B.n290 10.6151
R1735 B.n692 B.n691 10.6151
R1736 B.n693 B.n692 10.6151
R1737 B.n693 B.n0 10.6151
R1738 B.n570 B.n569 10.6151
R1739 B.n569 B.n568 10.6151
R1740 B.n568 B.n567 10.6151
R1741 B.n567 B.n565 10.6151
R1742 B.n565 B.n562 10.6151
R1743 B.n562 B.n561 10.6151
R1744 B.n561 B.n558 10.6151
R1745 B.n558 B.n557 10.6151
R1746 B.n557 B.n554 10.6151
R1747 B.n554 B.n553 10.6151
R1748 B.n553 B.n550 10.6151
R1749 B.n550 B.n549 10.6151
R1750 B.n549 B.n546 10.6151
R1751 B.n546 B.n545 10.6151
R1752 B.n545 B.n542 10.6151
R1753 B.n542 B.n541 10.6151
R1754 B.n541 B.n538 10.6151
R1755 B.n538 B.n537 10.6151
R1756 B.n537 B.n534 10.6151
R1757 B.n534 B.n533 10.6151
R1758 B.n533 B.n530 10.6151
R1759 B.n530 B.n529 10.6151
R1760 B.n529 B.n526 10.6151
R1761 B.n526 B.n525 10.6151
R1762 B.n525 B.n522 10.6151
R1763 B.n522 B.n521 10.6151
R1764 B.n521 B.n518 10.6151
R1765 B.n518 B.n517 10.6151
R1766 B.n517 B.n514 10.6151
R1767 B.n514 B.n513 10.6151
R1768 B.n513 B.n510 10.6151
R1769 B.n510 B.n509 10.6151
R1770 B.n509 B.n506 10.6151
R1771 B.n506 B.n505 10.6151
R1772 B.n505 B.n502 10.6151
R1773 B.n500 B.n497 10.6151
R1774 B.n497 B.n496 10.6151
R1775 B.n496 B.n493 10.6151
R1776 B.n493 B.n492 10.6151
R1777 B.n492 B.n489 10.6151
R1778 B.n489 B.n488 10.6151
R1779 B.n488 B.n485 10.6151
R1780 B.n485 B.n484 10.6151
R1781 B.n484 B.n481 10.6151
R1782 B.n479 B.n476 10.6151
R1783 B.n476 B.n475 10.6151
R1784 B.n475 B.n472 10.6151
R1785 B.n472 B.n471 10.6151
R1786 B.n471 B.n468 10.6151
R1787 B.n468 B.n467 10.6151
R1788 B.n467 B.n464 10.6151
R1789 B.n464 B.n463 10.6151
R1790 B.n463 B.n460 10.6151
R1791 B.n460 B.n459 10.6151
R1792 B.n459 B.n456 10.6151
R1793 B.n456 B.n455 10.6151
R1794 B.n455 B.n452 10.6151
R1795 B.n452 B.n451 10.6151
R1796 B.n451 B.n448 10.6151
R1797 B.n448 B.n447 10.6151
R1798 B.n447 B.n444 10.6151
R1799 B.n444 B.n443 10.6151
R1800 B.n443 B.n440 10.6151
R1801 B.n440 B.n439 10.6151
R1802 B.n439 B.n436 10.6151
R1803 B.n436 B.n435 10.6151
R1804 B.n435 B.n432 10.6151
R1805 B.n432 B.n431 10.6151
R1806 B.n431 B.n428 10.6151
R1807 B.n428 B.n427 10.6151
R1808 B.n427 B.n424 10.6151
R1809 B.n424 B.n423 10.6151
R1810 B.n423 B.n420 10.6151
R1811 B.n420 B.n419 10.6151
R1812 B.n419 B.n416 10.6151
R1813 B.n416 B.n415 10.6151
R1814 B.n415 B.n412 10.6151
R1815 B.n412 B.n365 10.6151
R1816 B.n575 B.n365 10.6151
R1817 B.n577 B.n576 10.6151
R1818 B.n577 B.n357 10.6151
R1819 B.n587 B.n357 10.6151
R1820 B.n588 B.n587 10.6151
R1821 B.n589 B.n588 10.6151
R1822 B.n589 B.n349 10.6151
R1823 B.n599 B.n349 10.6151
R1824 B.n600 B.n599 10.6151
R1825 B.n601 B.n600 10.6151
R1826 B.n601 B.n341 10.6151
R1827 B.n611 B.n341 10.6151
R1828 B.n612 B.n611 10.6151
R1829 B.n613 B.n612 10.6151
R1830 B.n613 B.n333 10.6151
R1831 B.n623 B.n333 10.6151
R1832 B.n624 B.n623 10.6151
R1833 B.n625 B.n624 10.6151
R1834 B.n625 B.n326 10.6151
R1835 B.n636 B.n326 10.6151
R1836 B.n637 B.n636 10.6151
R1837 B.n638 B.n637 10.6151
R1838 B.n638 B.n318 10.6151
R1839 B.n648 B.n318 10.6151
R1840 B.n649 B.n648 10.6151
R1841 B.n650 B.n649 10.6151
R1842 B.n650 B.n310 10.6151
R1843 B.n660 B.n310 10.6151
R1844 B.n661 B.n660 10.6151
R1845 B.n662 B.n661 10.6151
R1846 B.n662 B.n302 10.6151
R1847 B.n672 B.n302 10.6151
R1848 B.n673 B.n672 10.6151
R1849 B.n674 B.n673 10.6151
R1850 B.n674 B.n294 10.6151
R1851 B.n684 B.n294 10.6151
R1852 B.n685 B.n684 10.6151
R1853 B.n687 B.n685 10.6151
R1854 B.n687 B.n686 10.6151
R1855 B.n686 B.n286 10.6151
R1856 B.n698 B.n286 10.6151
R1857 B.n699 B.n698 10.6151
R1858 B.n700 B.n699 10.6151
R1859 B.n701 B.n700 10.6151
R1860 B.n702 B.n701 10.6151
R1861 B.n705 B.n702 10.6151
R1862 B.n706 B.n705 10.6151
R1863 B.n707 B.n706 10.6151
R1864 B.n708 B.n707 10.6151
R1865 B.n710 B.n708 10.6151
R1866 B.n711 B.n710 10.6151
R1867 B.n712 B.n711 10.6151
R1868 B.n713 B.n712 10.6151
R1869 B.n715 B.n713 10.6151
R1870 B.n716 B.n715 10.6151
R1871 B.n717 B.n716 10.6151
R1872 B.n718 B.n717 10.6151
R1873 B.n720 B.n718 10.6151
R1874 B.n721 B.n720 10.6151
R1875 B.n722 B.n721 10.6151
R1876 B.n723 B.n722 10.6151
R1877 B.n725 B.n723 10.6151
R1878 B.n726 B.n725 10.6151
R1879 B.n727 B.n726 10.6151
R1880 B.n728 B.n727 10.6151
R1881 B.n730 B.n728 10.6151
R1882 B.n731 B.n730 10.6151
R1883 B.n732 B.n731 10.6151
R1884 B.n733 B.n732 10.6151
R1885 B.n735 B.n733 10.6151
R1886 B.n736 B.n735 10.6151
R1887 B.n737 B.n736 10.6151
R1888 B.n738 B.n737 10.6151
R1889 B.n740 B.n738 10.6151
R1890 B.n741 B.n740 10.6151
R1891 B.n742 B.n741 10.6151
R1892 B.n743 B.n742 10.6151
R1893 B.n745 B.n743 10.6151
R1894 B.n746 B.n745 10.6151
R1895 B.n747 B.n746 10.6151
R1896 B.n748 B.n747 10.6151
R1897 B.n750 B.n748 10.6151
R1898 B.n751 B.n750 10.6151
R1899 B.n752 B.n751 10.6151
R1900 B.n834 B.n1 10.6151
R1901 B.n834 B.n833 10.6151
R1902 B.n833 B.n832 10.6151
R1903 B.n832 B.n10 10.6151
R1904 B.n826 B.n10 10.6151
R1905 B.n826 B.n825 10.6151
R1906 B.n825 B.n824 10.6151
R1907 B.n824 B.n18 10.6151
R1908 B.n818 B.n18 10.6151
R1909 B.n818 B.n817 10.6151
R1910 B.n817 B.n816 10.6151
R1911 B.n816 B.n25 10.6151
R1912 B.n810 B.n25 10.6151
R1913 B.n810 B.n809 10.6151
R1914 B.n809 B.n808 10.6151
R1915 B.n808 B.n32 10.6151
R1916 B.n802 B.n32 10.6151
R1917 B.n802 B.n801 10.6151
R1918 B.n801 B.n800 10.6151
R1919 B.n800 B.n39 10.6151
R1920 B.n794 B.n39 10.6151
R1921 B.n794 B.n793 10.6151
R1922 B.n793 B.n792 10.6151
R1923 B.n792 B.n45 10.6151
R1924 B.n786 B.n45 10.6151
R1925 B.n786 B.n785 10.6151
R1926 B.n785 B.n784 10.6151
R1927 B.n784 B.n53 10.6151
R1928 B.n778 B.n53 10.6151
R1929 B.n778 B.n777 10.6151
R1930 B.n777 B.n776 10.6151
R1931 B.n776 B.n60 10.6151
R1932 B.n770 B.n60 10.6151
R1933 B.n770 B.n769 10.6151
R1934 B.n769 B.n768 10.6151
R1935 B.n768 B.n67 10.6151
R1936 B.n762 B.n67 10.6151
R1937 B.n762 B.n761 10.6151
R1938 B.n761 B.n760 10.6151
R1939 B.n760 B.n74 10.6151
R1940 B.n127 B.n126 10.6151
R1941 B.n130 B.n127 10.6151
R1942 B.n131 B.n130 10.6151
R1943 B.n134 B.n131 10.6151
R1944 B.n135 B.n134 10.6151
R1945 B.n138 B.n135 10.6151
R1946 B.n139 B.n138 10.6151
R1947 B.n142 B.n139 10.6151
R1948 B.n143 B.n142 10.6151
R1949 B.n146 B.n143 10.6151
R1950 B.n147 B.n146 10.6151
R1951 B.n150 B.n147 10.6151
R1952 B.n151 B.n150 10.6151
R1953 B.n154 B.n151 10.6151
R1954 B.n155 B.n154 10.6151
R1955 B.n158 B.n155 10.6151
R1956 B.n159 B.n158 10.6151
R1957 B.n162 B.n159 10.6151
R1958 B.n163 B.n162 10.6151
R1959 B.n166 B.n163 10.6151
R1960 B.n167 B.n166 10.6151
R1961 B.n170 B.n167 10.6151
R1962 B.n171 B.n170 10.6151
R1963 B.n174 B.n171 10.6151
R1964 B.n175 B.n174 10.6151
R1965 B.n178 B.n175 10.6151
R1966 B.n179 B.n178 10.6151
R1967 B.n182 B.n179 10.6151
R1968 B.n183 B.n182 10.6151
R1969 B.n186 B.n183 10.6151
R1970 B.n187 B.n186 10.6151
R1971 B.n190 B.n187 10.6151
R1972 B.n191 B.n190 10.6151
R1973 B.n194 B.n191 10.6151
R1974 B.n195 B.n194 10.6151
R1975 B.n199 B.n198 10.6151
R1976 B.n202 B.n199 10.6151
R1977 B.n203 B.n202 10.6151
R1978 B.n206 B.n203 10.6151
R1979 B.n207 B.n206 10.6151
R1980 B.n210 B.n207 10.6151
R1981 B.n211 B.n210 10.6151
R1982 B.n214 B.n211 10.6151
R1983 B.n215 B.n214 10.6151
R1984 B.n219 B.n218 10.6151
R1985 B.n222 B.n219 10.6151
R1986 B.n223 B.n222 10.6151
R1987 B.n226 B.n223 10.6151
R1988 B.n227 B.n226 10.6151
R1989 B.n230 B.n227 10.6151
R1990 B.n231 B.n230 10.6151
R1991 B.n234 B.n231 10.6151
R1992 B.n235 B.n234 10.6151
R1993 B.n238 B.n235 10.6151
R1994 B.n239 B.n238 10.6151
R1995 B.n242 B.n239 10.6151
R1996 B.n243 B.n242 10.6151
R1997 B.n246 B.n243 10.6151
R1998 B.n247 B.n246 10.6151
R1999 B.n250 B.n247 10.6151
R2000 B.n251 B.n250 10.6151
R2001 B.n254 B.n251 10.6151
R2002 B.n255 B.n254 10.6151
R2003 B.n258 B.n255 10.6151
R2004 B.n259 B.n258 10.6151
R2005 B.n262 B.n259 10.6151
R2006 B.n263 B.n262 10.6151
R2007 B.n266 B.n263 10.6151
R2008 B.n267 B.n266 10.6151
R2009 B.n270 B.n267 10.6151
R2010 B.n271 B.n270 10.6151
R2011 B.n274 B.n271 10.6151
R2012 B.n275 B.n274 10.6151
R2013 B.n278 B.n275 10.6151
R2014 B.n279 B.n278 10.6151
R2015 B.n282 B.n279 10.6151
R2016 B.n284 B.n282 10.6151
R2017 B.n285 B.n284 10.6151
R2018 B.n753 B.n285 10.6151
R2019 B.n502 B.n501 9.36635
R2020 B.n480 B.n479 9.36635
R2021 B.n195 B.n124 9.36635
R2022 B.n218 B.n121 9.36635
R2023 B.n842 B.n0 8.11757
R2024 B.n842 B.n1 8.11757
R2025 B.n634 B.t1 2.84563
R2026 B.n796 B.t4 2.84563
R2027 B.n501 B.n500 1.24928
R2028 B.n481 B.n480 1.24928
R2029 B.n198 B.n124 1.24928
R2030 B.n215 B.n121 1.24928
R2031 VN.n29 VN.n16 161.3
R2032 VN.n28 VN.n27 161.3
R2033 VN.n26 VN.n17 161.3
R2034 VN.n25 VN.n24 161.3
R2035 VN.n23 VN.n18 161.3
R2036 VN.n22 VN.n21 161.3
R2037 VN.n13 VN.n0 161.3
R2038 VN.n12 VN.n11 161.3
R2039 VN.n10 VN.n1 161.3
R2040 VN.n9 VN.n8 161.3
R2041 VN.n7 VN.n2 161.3
R2042 VN.n6 VN.n5 161.3
R2043 VN.n4 VN.t1 129.466
R2044 VN.n20 VN.t4 129.466
R2045 VN.n15 VN.n14 105.864
R2046 VN.n31 VN.n30 105.864
R2047 VN.n3 VN.t5 97.4525
R2048 VN.n14 VN.t3 97.4525
R2049 VN.n19 VN.t2 97.4525
R2050 VN.n30 VN.t0 97.4525
R2051 VN.n4 VN.n3 59.8984
R2052 VN.n20 VN.n19 59.8984
R2053 VN.n8 VN.n1 56.5193
R2054 VN.n24 VN.n17 56.5193
R2055 VN VN.n31 47.1913
R2056 VN.n7 VN.n6 24.4675
R2057 VN.n8 VN.n7 24.4675
R2058 VN.n12 VN.n1 24.4675
R2059 VN.n13 VN.n12 24.4675
R2060 VN.n24 VN.n23 24.4675
R2061 VN.n23 VN.n22 24.4675
R2062 VN.n29 VN.n28 24.4675
R2063 VN.n28 VN.n17 24.4675
R2064 VN.n6 VN.n3 12.234
R2065 VN.n22 VN.n19 12.234
R2066 VN.n21 VN.n20 7.17115
R2067 VN.n5 VN.n4 7.17115
R2068 VN.n14 VN.n13 4.8939
R2069 VN.n30 VN.n29 4.8939
R2070 VN.n31 VN.n16 0.278367
R2071 VN.n15 VN.n0 0.278367
R2072 VN.n27 VN.n16 0.189894
R2073 VN.n27 VN.n26 0.189894
R2074 VN.n26 VN.n25 0.189894
R2075 VN.n25 VN.n18 0.189894
R2076 VN.n21 VN.n18 0.189894
R2077 VN.n5 VN.n2 0.189894
R2078 VN.n9 VN.n2 0.189894
R2079 VN.n10 VN.n9 0.189894
R2080 VN.n11 VN.n10 0.189894
R2081 VN.n11 VN.n0 0.189894
R2082 VN VN.n15 0.153454
R2083 VDD2.n103 VDD2.n55 289.615
R2084 VDD2.n48 VDD2.n0 289.615
R2085 VDD2.n104 VDD2.n103 185
R2086 VDD2.n102 VDD2.n101 185
R2087 VDD2.n59 VDD2.n58 185
R2088 VDD2.n96 VDD2.n95 185
R2089 VDD2.n94 VDD2.n61 185
R2090 VDD2.n93 VDD2.n92 185
R2091 VDD2.n64 VDD2.n62 185
R2092 VDD2.n87 VDD2.n86 185
R2093 VDD2.n85 VDD2.n84 185
R2094 VDD2.n68 VDD2.n67 185
R2095 VDD2.n79 VDD2.n78 185
R2096 VDD2.n77 VDD2.n76 185
R2097 VDD2.n72 VDD2.n71 185
R2098 VDD2.n16 VDD2.n15 185
R2099 VDD2.n21 VDD2.n20 185
R2100 VDD2.n23 VDD2.n22 185
R2101 VDD2.n12 VDD2.n11 185
R2102 VDD2.n29 VDD2.n28 185
R2103 VDD2.n31 VDD2.n30 185
R2104 VDD2.n8 VDD2.n7 185
R2105 VDD2.n38 VDD2.n37 185
R2106 VDD2.n39 VDD2.n6 185
R2107 VDD2.n41 VDD2.n40 185
R2108 VDD2.n4 VDD2.n3 185
R2109 VDD2.n47 VDD2.n46 185
R2110 VDD2.n49 VDD2.n48 185
R2111 VDD2.n73 VDD2.t5 149.524
R2112 VDD2.n17 VDD2.t4 149.524
R2113 VDD2.n103 VDD2.n102 104.615
R2114 VDD2.n102 VDD2.n58 104.615
R2115 VDD2.n95 VDD2.n58 104.615
R2116 VDD2.n95 VDD2.n94 104.615
R2117 VDD2.n94 VDD2.n93 104.615
R2118 VDD2.n93 VDD2.n62 104.615
R2119 VDD2.n86 VDD2.n62 104.615
R2120 VDD2.n86 VDD2.n85 104.615
R2121 VDD2.n85 VDD2.n67 104.615
R2122 VDD2.n78 VDD2.n67 104.615
R2123 VDD2.n78 VDD2.n77 104.615
R2124 VDD2.n77 VDD2.n71 104.615
R2125 VDD2.n21 VDD2.n15 104.615
R2126 VDD2.n22 VDD2.n21 104.615
R2127 VDD2.n22 VDD2.n11 104.615
R2128 VDD2.n29 VDD2.n11 104.615
R2129 VDD2.n30 VDD2.n29 104.615
R2130 VDD2.n30 VDD2.n7 104.615
R2131 VDD2.n38 VDD2.n7 104.615
R2132 VDD2.n39 VDD2.n38 104.615
R2133 VDD2.n40 VDD2.n39 104.615
R2134 VDD2.n40 VDD2.n3 104.615
R2135 VDD2.n47 VDD2.n3 104.615
R2136 VDD2.n48 VDD2.n47 104.615
R2137 VDD2.n54 VDD2.n53 67.6596
R2138 VDD2 VDD2.n109 67.6568
R2139 VDD2.n54 VDD2.n52 55.1121
R2140 VDD2.n108 VDD2.n107 53.3247
R2141 VDD2.t5 VDD2.n71 52.3082
R2142 VDD2.t4 VDD2.n15 52.3082
R2143 VDD2.n108 VDD2.n54 40.4847
R2144 VDD2.n96 VDD2.n61 13.1884
R2145 VDD2.n41 VDD2.n6 13.1884
R2146 VDD2.n97 VDD2.n59 12.8005
R2147 VDD2.n92 VDD2.n63 12.8005
R2148 VDD2.n37 VDD2.n36 12.8005
R2149 VDD2.n42 VDD2.n4 12.8005
R2150 VDD2.n101 VDD2.n100 12.0247
R2151 VDD2.n91 VDD2.n64 12.0247
R2152 VDD2.n35 VDD2.n8 12.0247
R2153 VDD2.n46 VDD2.n45 12.0247
R2154 VDD2.n104 VDD2.n57 11.249
R2155 VDD2.n88 VDD2.n87 11.249
R2156 VDD2.n32 VDD2.n31 11.249
R2157 VDD2.n49 VDD2.n2 11.249
R2158 VDD2.n105 VDD2.n55 10.4732
R2159 VDD2.n84 VDD2.n66 10.4732
R2160 VDD2.n28 VDD2.n10 10.4732
R2161 VDD2.n50 VDD2.n0 10.4732
R2162 VDD2.n73 VDD2.n72 10.2747
R2163 VDD2.n17 VDD2.n16 10.2747
R2164 VDD2.n83 VDD2.n68 9.69747
R2165 VDD2.n27 VDD2.n12 9.69747
R2166 VDD2.n107 VDD2.n106 9.45567
R2167 VDD2.n52 VDD2.n51 9.45567
R2168 VDD2.n75 VDD2.n74 9.3005
R2169 VDD2.n70 VDD2.n69 9.3005
R2170 VDD2.n81 VDD2.n80 9.3005
R2171 VDD2.n83 VDD2.n82 9.3005
R2172 VDD2.n66 VDD2.n65 9.3005
R2173 VDD2.n89 VDD2.n88 9.3005
R2174 VDD2.n91 VDD2.n90 9.3005
R2175 VDD2.n63 VDD2.n60 9.3005
R2176 VDD2.n106 VDD2.n105 9.3005
R2177 VDD2.n57 VDD2.n56 9.3005
R2178 VDD2.n100 VDD2.n99 9.3005
R2179 VDD2.n98 VDD2.n97 9.3005
R2180 VDD2.n51 VDD2.n50 9.3005
R2181 VDD2.n2 VDD2.n1 9.3005
R2182 VDD2.n45 VDD2.n44 9.3005
R2183 VDD2.n43 VDD2.n42 9.3005
R2184 VDD2.n19 VDD2.n18 9.3005
R2185 VDD2.n14 VDD2.n13 9.3005
R2186 VDD2.n25 VDD2.n24 9.3005
R2187 VDD2.n27 VDD2.n26 9.3005
R2188 VDD2.n10 VDD2.n9 9.3005
R2189 VDD2.n33 VDD2.n32 9.3005
R2190 VDD2.n35 VDD2.n34 9.3005
R2191 VDD2.n36 VDD2.n5 9.3005
R2192 VDD2.n80 VDD2.n79 8.92171
R2193 VDD2.n24 VDD2.n23 8.92171
R2194 VDD2.n76 VDD2.n70 8.14595
R2195 VDD2.n20 VDD2.n14 8.14595
R2196 VDD2.n75 VDD2.n72 7.3702
R2197 VDD2.n19 VDD2.n16 7.3702
R2198 VDD2.n76 VDD2.n75 5.81868
R2199 VDD2.n20 VDD2.n19 5.81868
R2200 VDD2.n79 VDD2.n70 5.04292
R2201 VDD2.n23 VDD2.n14 5.04292
R2202 VDD2.n80 VDD2.n68 4.26717
R2203 VDD2.n24 VDD2.n12 4.26717
R2204 VDD2.n107 VDD2.n55 3.49141
R2205 VDD2.n84 VDD2.n83 3.49141
R2206 VDD2.n28 VDD2.n27 3.49141
R2207 VDD2.n52 VDD2.n0 3.49141
R2208 VDD2.n74 VDD2.n73 2.84303
R2209 VDD2.n18 VDD2.n17 2.84303
R2210 VDD2.n105 VDD2.n104 2.71565
R2211 VDD2.n87 VDD2.n66 2.71565
R2212 VDD2.n31 VDD2.n10 2.71565
R2213 VDD2.n50 VDD2.n49 2.71565
R2214 VDD2.n109 VDD2.t3 1.94358
R2215 VDD2.n109 VDD2.t1 1.94358
R2216 VDD2.n53 VDD2.t0 1.94358
R2217 VDD2.n53 VDD2.t2 1.94358
R2218 VDD2.n101 VDD2.n57 1.93989
R2219 VDD2.n88 VDD2.n64 1.93989
R2220 VDD2.n32 VDD2.n8 1.93989
R2221 VDD2.n46 VDD2.n2 1.93989
R2222 VDD2 VDD2.n108 1.90136
R2223 VDD2.n100 VDD2.n59 1.16414
R2224 VDD2.n92 VDD2.n91 1.16414
R2225 VDD2.n37 VDD2.n35 1.16414
R2226 VDD2.n45 VDD2.n4 1.16414
R2227 VDD2.n97 VDD2.n96 0.388379
R2228 VDD2.n63 VDD2.n61 0.388379
R2229 VDD2.n36 VDD2.n6 0.388379
R2230 VDD2.n42 VDD2.n41 0.388379
R2231 VDD2.n106 VDD2.n56 0.155672
R2232 VDD2.n99 VDD2.n56 0.155672
R2233 VDD2.n99 VDD2.n98 0.155672
R2234 VDD2.n98 VDD2.n60 0.155672
R2235 VDD2.n90 VDD2.n60 0.155672
R2236 VDD2.n90 VDD2.n89 0.155672
R2237 VDD2.n89 VDD2.n65 0.155672
R2238 VDD2.n82 VDD2.n65 0.155672
R2239 VDD2.n82 VDD2.n81 0.155672
R2240 VDD2.n81 VDD2.n69 0.155672
R2241 VDD2.n74 VDD2.n69 0.155672
R2242 VDD2.n18 VDD2.n13 0.155672
R2243 VDD2.n25 VDD2.n13 0.155672
R2244 VDD2.n26 VDD2.n25 0.155672
R2245 VDD2.n26 VDD2.n9 0.155672
R2246 VDD2.n33 VDD2.n9 0.155672
R2247 VDD2.n34 VDD2.n33 0.155672
R2248 VDD2.n34 VDD2.n5 0.155672
R2249 VDD2.n43 VDD2.n5 0.155672
R2250 VDD2.n44 VDD2.n43 0.155672
R2251 VDD2.n44 VDD2.n1 0.155672
R2252 VDD2.n51 VDD2.n1 0.155672
C0 VDD2 VP 0.451473f
C1 VTAIL VDD1 7.05327f
C2 VTAIL VN 5.94813f
C3 VDD1 VN 0.15071f
C4 VTAIL VP 5.9624f
C5 VDD1 VP 6.02786f
C6 VN VP 6.51729f
C7 VTAIL VDD2 7.10392f
C8 VDD1 VDD2 1.37617f
C9 VN VDD2 5.72999f
C10 VDD2 B 5.602246f
C11 VDD1 B 5.734435f
C12 VTAIL B 7.04176f
C13 VN B 12.501109f
C14 VP B 11.151477f
C15 VDD2.n0 B 0.031715f
C16 VDD2.n1 B 0.021432f
C17 VDD2.n2 B 0.011517f
C18 VDD2.n3 B 0.027221f
C19 VDD2.n4 B 0.012194f
C20 VDD2.n5 B 0.021432f
C21 VDD2.n6 B 0.011855f
C22 VDD2.n7 B 0.027221f
C23 VDD2.n8 B 0.012194f
C24 VDD2.n9 B 0.021432f
C25 VDD2.n10 B 0.011517f
C26 VDD2.n11 B 0.027221f
C27 VDD2.n12 B 0.012194f
C28 VDD2.n13 B 0.021432f
C29 VDD2.n14 B 0.011517f
C30 VDD2.n15 B 0.020416f
C31 VDD2.n16 B 0.019243f
C32 VDD2.t4 B 0.045768f
C33 VDD2.n17 B 0.139633f
C34 VDD2.n18 B 0.908656f
C35 VDD2.n19 B 0.011517f
C36 VDD2.n20 B 0.012194f
C37 VDD2.n21 B 0.027221f
C38 VDD2.n22 B 0.027221f
C39 VDD2.n23 B 0.012194f
C40 VDD2.n24 B 0.011517f
C41 VDD2.n25 B 0.021432f
C42 VDD2.n26 B 0.021432f
C43 VDD2.n27 B 0.011517f
C44 VDD2.n28 B 0.012194f
C45 VDD2.n29 B 0.027221f
C46 VDD2.n30 B 0.027221f
C47 VDD2.n31 B 0.012194f
C48 VDD2.n32 B 0.011517f
C49 VDD2.n33 B 0.021432f
C50 VDD2.n34 B 0.021432f
C51 VDD2.n35 B 0.011517f
C52 VDD2.n36 B 0.011517f
C53 VDD2.n37 B 0.012194f
C54 VDD2.n38 B 0.027221f
C55 VDD2.n39 B 0.027221f
C56 VDD2.n40 B 0.027221f
C57 VDD2.n41 B 0.011855f
C58 VDD2.n42 B 0.011517f
C59 VDD2.n43 B 0.021432f
C60 VDD2.n44 B 0.021432f
C61 VDD2.n45 B 0.011517f
C62 VDD2.n46 B 0.012194f
C63 VDD2.n47 B 0.027221f
C64 VDD2.n48 B 0.061742f
C65 VDD2.n49 B 0.012194f
C66 VDD2.n50 B 0.011517f
C67 VDD2.n51 B 0.056273f
C68 VDD2.n52 B 0.05526f
C69 VDD2.t0 B 0.172579f
C70 VDD2.t2 B 0.172579f
C71 VDD2.n53 B 1.52778f
C72 VDD2.n54 B 2.17116f
C73 VDD2.n55 B 0.031715f
C74 VDD2.n56 B 0.021432f
C75 VDD2.n57 B 0.011517f
C76 VDD2.n58 B 0.027221f
C77 VDD2.n59 B 0.012194f
C78 VDD2.n60 B 0.021432f
C79 VDD2.n61 B 0.011855f
C80 VDD2.n62 B 0.027221f
C81 VDD2.n63 B 0.011517f
C82 VDD2.n64 B 0.012194f
C83 VDD2.n65 B 0.021432f
C84 VDD2.n66 B 0.011517f
C85 VDD2.n67 B 0.027221f
C86 VDD2.n68 B 0.012194f
C87 VDD2.n69 B 0.021432f
C88 VDD2.n70 B 0.011517f
C89 VDD2.n71 B 0.020416f
C90 VDD2.n72 B 0.019243f
C91 VDD2.t5 B 0.045768f
C92 VDD2.n73 B 0.139633f
C93 VDD2.n74 B 0.908656f
C94 VDD2.n75 B 0.011517f
C95 VDD2.n76 B 0.012194f
C96 VDD2.n77 B 0.027221f
C97 VDD2.n78 B 0.027221f
C98 VDD2.n79 B 0.012194f
C99 VDD2.n80 B 0.011517f
C100 VDD2.n81 B 0.021432f
C101 VDD2.n82 B 0.021432f
C102 VDD2.n83 B 0.011517f
C103 VDD2.n84 B 0.012194f
C104 VDD2.n85 B 0.027221f
C105 VDD2.n86 B 0.027221f
C106 VDD2.n87 B 0.012194f
C107 VDD2.n88 B 0.011517f
C108 VDD2.n89 B 0.021432f
C109 VDD2.n90 B 0.021432f
C110 VDD2.n91 B 0.011517f
C111 VDD2.n92 B 0.012194f
C112 VDD2.n93 B 0.027221f
C113 VDD2.n94 B 0.027221f
C114 VDD2.n95 B 0.027221f
C115 VDD2.n96 B 0.011855f
C116 VDD2.n97 B 0.011517f
C117 VDD2.n98 B 0.021432f
C118 VDD2.n99 B 0.021432f
C119 VDD2.n100 B 0.011517f
C120 VDD2.n101 B 0.012194f
C121 VDD2.n102 B 0.027221f
C122 VDD2.n103 B 0.061742f
C123 VDD2.n104 B 0.012194f
C124 VDD2.n105 B 0.011517f
C125 VDD2.n106 B 0.056273f
C126 VDD2.n107 B 0.049784f
C127 VDD2.n108 B 2.06059f
C128 VDD2.t3 B 0.172579f
C129 VDD2.t1 B 0.172579f
C130 VDD2.n109 B 1.52776f
C131 VN.n0 B 0.031816f
C132 VN.t3 B 1.67985f
C133 VN.n1 B 0.040275f
C134 VN.n2 B 0.024132f
C135 VN.t5 B 1.67985f
C136 VN.n3 B 0.669337f
C137 VN.t1 B 1.86417f
C138 VN.n4 B 0.654914f
C139 VN.n5 B 0.230857f
C140 VN.n6 B 0.033874f
C141 VN.n7 B 0.044977f
C142 VN.n8 B 0.030188f
C143 VN.n9 B 0.024132f
C144 VN.n10 B 0.024132f
C145 VN.n11 B 0.024132f
C146 VN.n12 B 0.044977f
C147 VN.n13 B 0.027212f
C148 VN.n14 B 0.672879f
C149 VN.n15 B 0.041396f
C150 VN.n16 B 0.031816f
C151 VN.t0 B 1.67985f
C152 VN.n17 B 0.040275f
C153 VN.n18 B 0.024132f
C154 VN.t2 B 1.67985f
C155 VN.n19 B 0.669337f
C156 VN.t4 B 1.86417f
C157 VN.n20 B 0.654914f
C158 VN.n21 B 0.230857f
C159 VN.n22 B 0.033874f
C160 VN.n23 B 0.044977f
C161 VN.n24 B 0.030188f
C162 VN.n25 B 0.024132f
C163 VN.n26 B 0.024132f
C164 VN.n27 B 0.024132f
C165 VN.n28 B 0.044977f
C166 VN.n29 B 0.027212f
C167 VN.n30 B 0.672879f
C168 VN.n31 B 1.2352f
C169 VTAIL.t5 B 0.195508f
C170 VTAIL.t0 B 0.195508f
C171 VTAIL.n0 B 1.66415f
C172 VTAIL.n1 B 0.410382f
C173 VTAIL.n2 B 0.035929f
C174 VTAIL.n3 B 0.024279f
C175 VTAIL.n4 B 0.013047f
C176 VTAIL.n5 B 0.030837f
C177 VTAIL.n6 B 0.013814f
C178 VTAIL.n7 B 0.024279f
C179 VTAIL.n8 B 0.01343f
C180 VTAIL.n9 B 0.030837f
C181 VTAIL.n10 B 0.013814f
C182 VTAIL.n11 B 0.024279f
C183 VTAIL.n12 B 0.013047f
C184 VTAIL.n13 B 0.030837f
C185 VTAIL.n14 B 0.013814f
C186 VTAIL.n15 B 0.024279f
C187 VTAIL.n16 B 0.013047f
C188 VTAIL.n17 B 0.023128f
C189 VTAIL.n18 B 0.0218f
C190 VTAIL.t6 B 0.051849f
C191 VTAIL.n19 B 0.158184f
C192 VTAIL.n20 B 1.02938f
C193 VTAIL.n21 B 0.013047f
C194 VTAIL.n22 B 0.013814f
C195 VTAIL.n23 B 0.030837f
C196 VTAIL.n24 B 0.030837f
C197 VTAIL.n25 B 0.013814f
C198 VTAIL.n26 B 0.013047f
C199 VTAIL.n27 B 0.024279f
C200 VTAIL.n28 B 0.024279f
C201 VTAIL.n29 B 0.013047f
C202 VTAIL.n30 B 0.013814f
C203 VTAIL.n31 B 0.030837f
C204 VTAIL.n32 B 0.030837f
C205 VTAIL.n33 B 0.013814f
C206 VTAIL.n34 B 0.013047f
C207 VTAIL.n35 B 0.024279f
C208 VTAIL.n36 B 0.024279f
C209 VTAIL.n37 B 0.013047f
C210 VTAIL.n38 B 0.013047f
C211 VTAIL.n39 B 0.013814f
C212 VTAIL.n40 B 0.030837f
C213 VTAIL.n41 B 0.030837f
C214 VTAIL.n42 B 0.030837f
C215 VTAIL.n43 B 0.01343f
C216 VTAIL.n44 B 0.013047f
C217 VTAIL.n45 B 0.024279f
C218 VTAIL.n46 B 0.024279f
C219 VTAIL.n47 B 0.013047f
C220 VTAIL.n48 B 0.013814f
C221 VTAIL.n49 B 0.030837f
C222 VTAIL.n50 B 0.069945f
C223 VTAIL.n51 B 0.013814f
C224 VTAIL.n52 B 0.013047f
C225 VTAIL.n53 B 0.063749f
C226 VTAIL.n54 B 0.039686f
C227 VTAIL.n55 B 0.350128f
C228 VTAIL.t7 B 0.195508f
C229 VTAIL.t11 B 0.195508f
C230 VTAIL.n56 B 1.66415f
C231 VTAIL.n57 B 1.81859f
C232 VTAIL.t1 B 0.195508f
C233 VTAIL.t3 B 0.195508f
C234 VTAIL.n58 B 1.66416f
C235 VTAIL.n59 B 1.81859f
C236 VTAIL.n60 B 0.035929f
C237 VTAIL.n61 B 0.024279f
C238 VTAIL.n62 B 0.013047f
C239 VTAIL.n63 B 0.030837f
C240 VTAIL.n64 B 0.013814f
C241 VTAIL.n65 B 0.024279f
C242 VTAIL.n66 B 0.01343f
C243 VTAIL.n67 B 0.030837f
C244 VTAIL.n68 B 0.013047f
C245 VTAIL.n69 B 0.013814f
C246 VTAIL.n70 B 0.024279f
C247 VTAIL.n71 B 0.013047f
C248 VTAIL.n72 B 0.030837f
C249 VTAIL.n73 B 0.013814f
C250 VTAIL.n74 B 0.024279f
C251 VTAIL.n75 B 0.013047f
C252 VTAIL.n76 B 0.023128f
C253 VTAIL.n77 B 0.0218f
C254 VTAIL.t2 B 0.051849f
C255 VTAIL.n78 B 0.158184f
C256 VTAIL.n79 B 1.02938f
C257 VTAIL.n80 B 0.013047f
C258 VTAIL.n81 B 0.013814f
C259 VTAIL.n82 B 0.030837f
C260 VTAIL.n83 B 0.030837f
C261 VTAIL.n84 B 0.013814f
C262 VTAIL.n85 B 0.013047f
C263 VTAIL.n86 B 0.024279f
C264 VTAIL.n87 B 0.024279f
C265 VTAIL.n88 B 0.013047f
C266 VTAIL.n89 B 0.013814f
C267 VTAIL.n90 B 0.030837f
C268 VTAIL.n91 B 0.030837f
C269 VTAIL.n92 B 0.013814f
C270 VTAIL.n93 B 0.013047f
C271 VTAIL.n94 B 0.024279f
C272 VTAIL.n95 B 0.024279f
C273 VTAIL.n96 B 0.013047f
C274 VTAIL.n97 B 0.013814f
C275 VTAIL.n98 B 0.030837f
C276 VTAIL.n99 B 0.030837f
C277 VTAIL.n100 B 0.030837f
C278 VTAIL.n101 B 0.01343f
C279 VTAIL.n102 B 0.013047f
C280 VTAIL.n103 B 0.024279f
C281 VTAIL.n104 B 0.024279f
C282 VTAIL.n105 B 0.013047f
C283 VTAIL.n106 B 0.013814f
C284 VTAIL.n107 B 0.030837f
C285 VTAIL.n108 B 0.069945f
C286 VTAIL.n109 B 0.013814f
C287 VTAIL.n110 B 0.013047f
C288 VTAIL.n111 B 0.063749f
C289 VTAIL.n112 B 0.039686f
C290 VTAIL.n113 B 0.350128f
C291 VTAIL.t8 B 0.195508f
C292 VTAIL.t9 B 0.195508f
C293 VTAIL.n114 B 1.66416f
C294 VTAIL.n115 B 0.549979f
C295 VTAIL.n116 B 0.035929f
C296 VTAIL.n117 B 0.024279f
C297 VTAIL.n118 B 0.013047f
C298 VTAIL.n119 B 0.030837f
C299 VTAIL.n120 B 0.013814f
C300 VTAIL.n121 B 0.024279f
C301 VTAIL.n122 B 0.01343f
C302 VTAIL.n123 B 0.030837f
C303 VTAIL.n124 B 0.013047f
C304 VTAIL.n125 B 0.013814f
C305 VTAIL.n126 B 0.024279f
C306 VTAIL.n127 B 0.013047f
C307 VTAIL.n128 B 0.030837f
C308 VTAIL.n129 B 0.013814f
C309 VTAIL.n130 B 0.024279f
C310 VTAIL.n131 B 0.013047f
C311 VTAIL.n132 B 0.023128f
C312 VTAIL.n133 B 0.0218f
C313 VTAIL.t10 B 0.051849f
C314 VTAIL.n134 B 0.158184f
C315 VTAIL.n135 B 1.02938f
C316 VTAIL.n136 B 0.013047f
C317 VTAIL.n137 B 0.013814f
C318 VTAIL.n138 B 0.030837f
C319 VTAIL.n139 B 0.030837f
C320 VTAIL.n140 B 0.013814f
C321 VTAIL.n141 B 0.013047f
C322 VTAIL.n142 B 0.024279f
C323 VTAIL.n143 B 0.024279f
C324 VTAIL.n144 B 0.013047f
C325 VTAIL.n145 B 0.013814f
C326 VTAIL.n146 B 0.030837f
C327 VTAIL.n147 B 0.030837f
C328 VTAIL.n148 B 0.013814f
C329 VTAIL.n149 B 0.013047f
C330 VTAIL.n150 B 0.024279f
C331 VTAIL.n151 B 0.024279f
C332 VTAIL.n152 B 0.013047f
C333 VTAIL.n153 B 0.013814f
C334 VTAIL.n154 B 0.030837f
C335 VTAIL.n155 B 0.030837f
C336 VTAIL.n156 B 0.030837f
C337 VTAIL.n157 B 0.01343f
C338 VTAIL.n158 B 0.013047f
C339 VTAIL.n159 B 0.024279f
C340 VTAIL.n160 B 0.024279f
C341 VTAIL.n161 B 0.013047f
C342 VTAIL.n162 B 0.013814f
C343 VTAIL.n163 B 0.030837f
C344 VTAIL.n164 B 0.069945f
C345 VTAIL.n165 B 0.013814f
C346 VTAIL.n166 B 0.013047f
C347 VTAIL.n167 B 0.063749f
C348 VTAIL.n168 B 0.039686f
C349 VTAIL.n169 B 1.42652f
C350 VTAIL.n170 B 0.035929f
C351 VTAIL.n171 B 0.024279f
C352 VTAIL.n172 B 0.013047f
C353 VTAIL.n173 B 0.030837f
C354 VTAIL.n174 B 0.013814f
C355 VTAIL.n175 B 0.024279f
C356 VTAIL.n176 B 0.01343f
C357 VTAIL.n177 B 0.030837f
C358 VTAIL.n178 B 0.013814f
C359 VTAIL.n179 B 0.024279f
C360 VTAIL.n180 B 0.013047f
C361 VTAIL.n181 B 0.030837f
C362 VTAIL.n182 B 0.013814f
C363 VTAIL.n183 B 0.024279f
C364 VTAIL.n184 B 0.013047f
C365 VTAIL.n185 B 0.023128f
C366 VTAIL.n186 B 0.0218f
C367 VTAIL.t4 B 0.051849f
C368 VTAIL.n187 B 0.158184f
C369 VTAIL.n188 B 1.02938f
C370 VTAIL.n189 B 0.013047f
C371 VTAIL.n190 B 0.013814f
C372 VTAIL.n191 B 0.030837f
C373 VTAIL.n192 B 0.030837f
C374 VTAIL.n193 B 0.013814f
C375 VTAIL.n194 B 0.013047f
C376 VTAIL.n195 B 0.024279f
C377 VTAIL.n196 B 0.024279f
C378 VTAIL.n197 B 0.013047f
C379 VTAIL.n198 B 0.013814f
C380 VTAIL.n199 B 0.030837f
C381 VTAIL.n200 B 0.030837f
C382 VTAIL.n201 B 0.013814f
C383 VTAIL.n202 B 0.013047f
C384 VTAIL.n203 B 0.024279f
C385 VTAIL.n204 B 0.024279f
C386 VTAIL.n205 B 0.013047f
C387 VTAIL.n206 B 0.013047f
C388 VTAIL.n207 B 0.013814f
C389 VTAIL.n208 B 0.030837f
C390 VTAIL.n209 B 0.030837f
C391 VTAIL.n210 B 0.030837f
C392 VTAIL.n211 B 0.01343f
C393 VTAIL.n212 B 0.013047f
C394 VTAIL.n213 B 0.024279f
C395 VTAIL.n214 B 0.024279f
C396 VTAIL.n215 B 0.013047f
C397 VTAIL.n216 B 0.013814f
C398 VTAIL.n217 B 0.030837f
C399 VTAIL.n218 B 0.069945f
C400 VTAIL.n219 B 0.013814f
C401 VTAIL.n220 B 0.013047f
C402 VTAIL.n221 B 0.063749f
C403 VTAIL.n222 B 0.039686f
C404 VTAIL.n223 B 1.37392f
C405 VDD1.n0 B 0.032259f
C406 VDD1.n1 B 0.021799f
C407 VDD1.n2 B 0.011714f
C408 VDD1.n3 B 0.027688f
C409 VDD1.n4 B 0.012403f
C410 VDD1.n5 B 0.021799f
C411 VDD1.n6 B 0.012059f
C412 VDD1.n7 B 0.027688f
C413 VDD1.n8 B 0.011714f
C414 VDD1.n9 B 0.012403f
C415 VDD1.n10 B 0.021799f
C416 VDD1.n11 B 0.011714f
C417 VDD1.n12 B 0.027688f
C418 VDD1.n13 B 0.012403f
C419 VDD1.n14 B 0.021799f
C420 VDD1.n15 B 0.011714f
C421 VDD1.n16 B 0.020766f
C422 VDD1.n17 B 0.019573f
C423 VDD1.t1 B 0.046553f
C424 VDD1.n18 B 0.142027f
C425 VDD1.n19 B 0.924237f
C426 VDD1.n20 B 0.011714f
C427 VDD1.n21 B 0.012403f
C428 VDD1.n22 B 0.027688f
C429 VDD1.n23 B 0.027688f
C430 VDD1.n24 B 0.012403f
C431 VDD1.n25 B 0.011714f
C432 VDD1.n26 B 0.021799f
C433 VDD1.n27 B 0.021799f
C434 VDD1.n28 B 0.011714f
C435 VDD1.n29 B 0.012403f
C436 VDD1.n30 B 0.027688f
C437 VDD1.n31 B 0.027688f
C438 VDD1.n32 B 0.012403f
C439 VDD1.n33 B 0.011714f
C440 VDD1.n34 B 0.021799f
C441 VDD1.n35 B 0.021799f
C442 VDD1.n36 B 0.011714f
C443 VDD1.n37 B 0.012403f
C444 VDD1.n38 B 0.027688f
C445 VDD1.n39 B 0.027688f
C446 VDD1.n40 B 0.027688f
C447 VDD1.n41 B 0.012059f
C448 VDD1.n42 B 0.011714f
C449 VDD1.n43 B 0.021799f
C450 VDD1.n44 B 0.021799f
C451 VDD1.n45 B 0.011714f
C452 VDD1.n46 B 0.012403f
C453 VDD1.n47 B 0.027688f
C454 VDD1.n48 B 0.0628f
C455 VDD1.n49 B 0.012403f
C456 VDD1.n50 B 0.011714f
C457 VDD1.n51 B 0.057238f
C458 VDD1.n52 B 0.056813f
C459 VDD1.n53 B 0.032259f
C460 VDD1.n54 B 0.021799f
C461 VDD1.n55 B 0.011714f
C462 VDD1.n56 B 0.027688f
C463 VDD1.n57 B 0.012403f
C464 VDD1.n58 B 0.021799f
C465 VDD1.n59 B 0.012059f
C466 VDD1.n60 B 0.027688f
C467 VDD1.n61 B 0.012403f
C468 VDD1.n62 B 0.021799f
C469 VDD1.n63 B 0.011714f
C470 VDD1.n64 B 0.027688f
C471 VDD1.n65 B 0.012403f
C472 VDD1.n66 B 0.021799f
C473 VDD1.n67 B 0.011714f
C474 VDD1.n68 B 0.020766f
C475 VDD1.n69 B 0.019573f
C476 VDD1.t0 B 0.046553f
C477 VDD1.n70 B 0.142027f
C478 VDD1.n71 B 0.924237f
C479 VDD1.n72 B 0.011714f
C480 VDD1.n73 B 0.012403f
C481 VDD1.n74 B 0.027688f
C482 VDD1.n75 B 0.027688f
C483 VDD1.n76 B 0.012403f
C484 VDD1.n77 B 0.011714f
C485 VDD1.n78 B 0.021799f
C486 VDD1.n79 B 0.021799f
C487 VDD1.n80 B 0.011714f
C488 VDD1.n81 B 0.012403f
C489 VDD1.n82 B 0.027688f
C490 VDD1.n83 B 0.027688f
C491 VDD1.n84 B 0.012403f
C492 VDD1.n85 B 0.011714f
C493 VDD1.n86 B 0.021799f
C494 VDD1.n87 B 0.021799f
C495 VDD1.n88 B 0.011714f
C496 VDD1.n89 B 0.011714f
C497 VDD1.n90 B 0.012403f
C498 VDD1.n91 B 0.027688f
C499 VDD1.n92 B 0.027688f
C500 VDD1.n93 B 0.027688f
C501 VDD1.n94 B 0.012059f
C502 VDD1.n95 B 0.011714f
C503 VDD1.n96 B 0.021799f
C504 VDD1.n97 B 0.021799f
C505 VDD1.n98 B 0.011714f
C506 VDD1.n99 B 0.012403f
C507 VDD1.n100 B 0.027688f
C508 VDD1.n101 B 0.0628f
C509 VDD1.n102 B 0.012403f
C510 VDD1.n103 B 0.011714f
C511 VDD1.n104 B 0.057238f
C512 VDD1.n105 B 0.056207f
C513 VDD1.t4 B 0.175539f
C514 VDD1.t2 B 0.175539f
C515 VDD1.n106 B 1.55398f
C516 VDD1.n107 B 2.31354f
C517 VDD1.t5 B 0.175539f
C518 VDD1.t3 B 0.175539f
C519 VDD1.n108 B 1.5507f
C520 VDD1.n109 B 2.28732f
C521 VP.n0 B 0.03258f
C522 VP.t5 B 1.7202f
C523 VP.n1 B 0.041242f
C524 VP.n2 B 0.024712f
C525 VP.t0 B 1.7202f
C526 VP.n3 B 0.615529f
C527 VP.n4 B 0.024712f
C528 VP.n5 B 0.041242f
C529 VP.n6 B 0.03258f
C530 VP.t4 B 1.7202f
C531 VP.n7 B 0.03258f
C532 VP.t1 B 1.7202f
C533 VP.n8 B 0.041242f
C534 VP.n9 B 0.024712f
C535 VP.t2 B 1.7202f
C536 VP.n10 B 0.685414f
C537 VP.t3 B 1.90894f
C538 VP.n11 B 0.670644f
C539 VP.n12 B 0.236402f
C540 VP.n13 B 0.034688f
C541 VP.n14 B 0.046057f
C542 VP.n15 B 0.030913f
C543 VP.n16 B 0.024712f
C544 VP.n17 B 0.024712f
C545 VP.n18 B 0.024712f
C546 VP.n19 B 0.046057f
C547 VP.n20 B 0.027866f
C548 VP.n21 B 0.68904f
C549 VP.n22 B 1.25145f
C550 VP.n23 B 1.27038f
C551 VP.n24 B 0.68904f
C552 VP.n25 B 0.027866f
C553 VP.n26 B 0.046057f
C554 VP.n27 B 0.024712f
C555 VP.n28 B 0.024712f
C556 VP.n29 B 0.024712f
C557 VP.n30 B 0.030913f
C558 VP.n31 B 0.046057f
C559 VP.n32 B 0.034688f
C560 VP.n33 B 0.024712f
C561 VP.n34 B 0.024712f
C562 VP.n35 B 0.034688f
C563 VP.n36 B 0.046057f
C564 VP.n37 B 0.030913f
C565 VP.n38 B 0.024712f
C566 VP.n39 B 0.024712f
C567 VP.n40 B 0.024712f
C568 VP.n41 B 0.046057f
C569 VP.n42 B 0.027866f
C570 VP.n43 B 0.68904f
C571 VP.n44 B 0.04239f
.ends

