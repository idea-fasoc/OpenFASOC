* NGSPICE file created from diff_pair_sample_0700.ext - technology: sky130A

.subckt diff_pair_sample_0700 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t1 VP.t0 VTAIL.t2 B.t0 sky130_fd_pr__nfet_01v8 ad=7.7454 pd=40.5 as=7.7454 ps=40.5 w=19.86 l=3.43
X1 B.t15 B.t13 B.t14 B.t3 sky130_fd_pr__nfet_01v8 ad=7.7454 pd=40.5 as=0 ps=0 w=19.86 l=3.43
X2 B.t12 B.t10 B.t11 B.t7 sky130_fd_pr__nfet_01v8 ad=7.7454 pd=40.5 as=0 ps=0 w=19.86 l=3.43
X3 B.t9 B.t6 B.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=7.7454 pd=40.5 as=0 ps=0 w=19.86 l=3.43
X4 B.t5 B.t2 B.t4 B.t3 sky130_fd_pr__nfet_01v8 ad=7.7454 pd=40.5 as=0 ps=0 w=19.86 l=3.43
X5 VDD2.t1 VN.t0 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=7.7454 pd=40.5 as=7.7454 ps=40.5 w=19.86 l=3.43
X6 VDD1.t0 VP.t1 VTAIL.t3 B.t1 sky130_fd_pr__nfet_01v8 ad=7.7454 pd=40.5 as=7.7454 ps=40.5 w=19.86 l=3.43
X7 VDD2.t0 VN.t1 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=7.7454 pd=40.5 as=7.7454 ps=40.5 w=19.86 l=3.43
R0 VP.n0 VP.t0 231.2
R1 VP.n0 VP.t1 178.387
R2 VP VP.n0 0.526373
R3 VTAIL.n1 VTAIL.t1 48.0139
R4 VTAIL.n3 VTAIL.t0 48.0137
R5 VTAIL.n0 VTAIL.t3 48.0137
R6 VTAIL.n2 VTAIL.t2 48.0137
R7 VTAIL.n1 VTAIL.n0 35.9703
R8 VTAIL.n3 VTAIL.n2 32.729
R9 VTAIL.n2 VTAIL.n1 2.09102
R10 VTAIL VTAIL.n0 1.33886
R11 VTAIL VTAIL.n3 0.752655
R12 VDD1 VDD1.t0 113.29
R13 VDD1 VDD1.t1 65.5611
R14 B.n672 B.n132 585
R15 B.n132 B.n57 585
R16 B.n674 B.n673 585
R17 B.n676 B.n131 585
R18 B.n679 B.n678 585
R19 B.n680 B.n130 585
R20 B.n682 B.n681 585
R21 B.n684 B.n129 585
R22 B.n687 B.n686 585
R23 B.n688 B.n128 585
R24 B.n690 B.n689 585
R25 B.n692 B.n127 585
R26 B.n695 B.n694 585
R27 B.n696 B.n126 585
R28 B.n698 B.n697 585
R29 B.n700 B.n125 585
R30 B.n703 B.n702 585
R31 B.n704 B.n124 585
R32 B.n706 B.n705 585
R33 B.n708 B.n123 585
R34 B.n711 B.n710 585
R35 B.n712 B.n122 585
R36 B.n714 B.n713 585
R37 B.n716 B.n121 585
R38 B.n719 B.n718 585
R39 B.n720 B.n120 585
R40 B.n722 B.n721 585
R41 B.n724 B.n119 585
R42 B.n727 B.n726 585
R43 B.n728 B.n118 585
R44 B.n730 B.n729 585
R45 B.n732 B.n117 585
R46 B.n735 B.n734 585
R47 B.n736 B.n116 585
R48 B.n738 B.n737 585
R49 B.n740 B.n115 585
R50 B.n743 B.n742 585
R51 B.n744 B.n114 585
R52 B.n746 B.n745 585
R53 B.n748 B.n113 585
R54 B.n751 B.n750 585
R55 B.n752 B.n112 585
R56 B.n754 B.n753 585
R57 B.n756 B.n111 585
R58 B.n759 B.n758 585
R59 B.n760 B.n110 585
R60 B.n762 B.n761 585
R61 B.n764 B.n109 585
R62 B.n767 B.n766 585
R63 B.n768 B.n108 585
R64 B.n770 B.n769 585
R65 B.n772 B.n107 585
R66 B.n775 B.n774 585
R67 B.n776 B.n106 585
R68 B.n778 B.n777 585
R69 B.n780 B.n105 585
R70 B.n783 B.n782 585
R71 B.n784 B.n104 585
R72 B.n786 B.n785 585
R73 B.n788 B.n103 585
R74 B.n791 B.n790 585
R75 B.n792 B.n102 585
R76 B.n794 B.n793 585
R77 B.n796 B.n101 585
R78 B.n798 B.n797 585
R79 B.n800 B.n799 585
R80 B.n803 B.n802 585
R81 B.n804 B.n96 585
R82 B.n806 B.n805 585
R83 B.n808 B.n95 585
R84 B.n811 B.n810 585
R85 B.n812 B.n94 585
R86 B.n814 B.n813 585
R87 B.n816 B.n93 585
R88 B.n819 B.n818 585
R89 B.n821 B.n90 585
R90 B.n823 B.n822 585
R91 B.n825 B.n89 585
R92 B.n828 B.n827 585
R93 B.n829 B.n88 585
R94 B.n831 B.n830 585
R95 B.n833 B.n87 585
R96 B.n836 B.n835 585
R97 B.n837 B.n86 585
R98 B.n839 B.n838 585
R99 B.n841 B.n85 585
R100 B.n844 B.n843 585
R101 B.n845 B.n84 585
R102 B.n847 B.n846 585
R103 B.n849 B.n83 585
R104 B.n852 B.n851 585
R105 B.n853 B.n82 585
R106 B.n855 B.n854 585
R107 B.n857 B.n81 585
R108 B.n860 B.n859 585
R109 B.n861 B.n80 585
R110 B.n863 B.n862 585
R111 B.n865 B.n79 585
R112 B.n868 B.n867 585
R113 B.n869 B.n78 585
R114 B.n871 B.n870 585
R115 B.n873 B.n77 585
R116 B.n876 B.n875 585
R117 B.n877 B.n76 585
R118 B.n879 B.n878 585
R119 B.n881 B.n75 585
R120 B.n884 B.n883 585
R121 B.n885 B.n74 585
R122 B.n887 B.n886 585
R123 B.n889 B.n73 585
R124 B.n892 B.n891 585
R125 B.n893 B.n72 585
R126 B.n895 B.n894 585
R127 B.n897 B.n71 585
R128 B.n900 B.n899 585
R129 B.n901 B.n70 585
R130 B.n903 B.n902 585
R131 B.n905 B.n69 585
R132 B.n908 B.n907 585
R133 B.n909 B.n68 585
R134 B.n911 B.n910 585
R135 B.n913 B.n67 585
R136 B.n916 B.n915 585
R137 B.n917 B.n66 585
R138 B.n919 B.n918 585
R139 B.n921 B.n65 585
R140 B.n924 B.n923 585
R141 B.n925 B.n64 585
R142 B.n927 B.n926 585
R143 B.n929 B.n63 585
R144 B.n932 B.n931 585
R145 B.n933 B.n62 585
R146 B.n935 B.n934 585
R147 B.n937 B.n61 585
R148 B.n940 B.n939 585
R149 B.n941 B.n60 585
R150 B.n943 B.n942 585
R151 B.n945 B.n59 585
R152 B.n948 B.n947 585
R153 B.n949 B.n58 585
R154 B.n671 B.n56 585
R155 B.n952 B.n56 585
R156 B.n670 B.n55 585
R157 B.n953 B.n55 585
R158 B.n669 B.n54 585
R159 B.n954 B.n54 585
R160 B.n668 B.n667 585
R161 B.n667 B.n50 585
R162 B.n666 B.n49 585
R163 B.n960 B.n49 585
R164 B.n665 B.n48 585
R165 B.n961 B.n48 585
R166 B.n664 B.n47 585
R167 B.n962 B.n47 585
R168 B.n663 B.n662 585
R169 B.n662 B.n43 585
R170 B.n661 B.n42 585
R171 B.n968 B.n42 585
R172 B.n660 B.n41 585
R173 B.n969 B.n41 585
R174 B.n659 B.n40 585
R175 B.n970 B.n40 585
R176 B.n658 B.n657 585
R177 B.n657 B.n36 585
R178 B.n656 B.n35 585
R179 B.n976 B.n35 585
R180 B.n655 B.n34 585
R181 B.n977 B.n34 585
R182 B.n654 B.n33 585
R183 B.n978 B.n33 585
R184 B.n653 B.n652 585
R185 B.n652 B.n29 585
R186 B.n651 B.n28 585
R187 B.n984 B.n28 585
R188 B.n650 B.n27 585
R189 B.n985 B.n27 585
R190 B.n649 B.n26 585
R191 B.n986 B.n26 585
R192 B.n648 B.n647 585
R193 B.n647 B.n22 585
R194 B.n646 B.n21 585
R195 B.n992 B.n21 585
R196 B.n645 B.n20 585
R197 B.n993 B.n20 585
R198 B.n644 B.n19 585
R199 B.n994 B.n19 585
R200 B.n643 B.n642 585
R201 B.n642 B.n15 585
R202 B.n641 B.n14 585
R203 B.n1000 B.n14 585
R204 B.n640 B.n13 585
R205 B.n1001 B.n13 585
R206 B.n639 B.n12 585
R207 B.n1002 B.n12 585
R208 B.n638 B.n637 585
R209 B.n637 B.n8 585
R210 B.n636 B.n7 585
R211 B.n1008 B.n7 585
R212 B.n635 B.n6 585
R213 B.n1009 B.n6 585
R214 B.n634 B.n5 585
R215 B.n1010 B.n5 585
R216 B.n633 B.n632 585
R217 B.n632 B.n4 585
R218 B.n631 B.n133 585
R219 B.n631 B.n630 585
R220 B.n621 B.n134 585
R221 B.n135 B.n134 585
R222 B.n623 B.n622 585
R223 B.n624 B.n623 585
R224 B.n620 B.n140 585
R225 B.n140 B.n139 585
R226 B.n619 B.n618 585
R227 B.n618 B.n617 585
R228 B.n142 B.n141 585
R229 B.n143 B.n142 585
R230 B.n610 B.n609 585
R231 B.n611 B.n610 585
R232 B.n608 B.n148 585
R233 B.n148 B.n147 585
R234 B.n607 B.n606 585
R235 B.n606 B.n605 585
R236 B.n150 B.n149 585
R237 B.n151 B.n150 585
R238 B.n598 B.n597 585
R239 B.n599 B.n598 585
R240 B.n596 B.n156 585
R241 B.n156 B.n155 585
R242 B.n595 B.n594 585
R243 B.n594 B.n593 585
R244 B.n158 B.n157 585
R245 B.n159 B.n158 585
R246 B.n586 B.n585 585
R247 B.n587 B.n586 585
R248 B.n584 B.n164 585
R249 B.n164 B.n163 585
R250 B.n583 B.n582 585
R251 B.n582 B.n581 585
R252 B.n166 B.n165 585
R253 B.n167 B.n166 585
R254 B.n574 B.n573 585
R255 B.n575 B.n574 585
R256 B.n572 B.n172 585
R257 B.n172 B.n171 585
R258 B.n571 B.n570 585
R259 B.n570 B.n569 585
R260 B.n174 B.n173 585
R261 B.n175 B.n174 585
R262 B.n562 B.n561 585
R263 B.n563 B.n562 585
R264 B.n560 B.n180 585
R265 B.n180 B.n179 585
R266 B.n559 B.n558 585
R267 B.n558 B.n557 585
R268 B.n182 B.n181 585
R269 B.n183 B.n182 585
R270 B.n550 B.n549 585
R271 B.n551 B.n550 585
R272 B.n548 B.n188 585
R273 B.n188 B.n187 585
R274 B.n547 B.n546 585
R275 B.n546 B.n545 585
R276 B.n542 B.n192 585
R277 B.n541 B.n540 585
R278 B.n538 B.n193 585
R279 B.n538 B.n191 585
R280 B.n537 B.n536 585
R281 B.n535 B.n534 585
R282 B.n533 B.n195 585
R283 B.n531 B.n530 585
R284 B.n529 B.n196 585
R285 B.n528 B.n527 585
R286 B.n525 B.n197 585
R287 B.n523 B.n522 585
R288 B.n521 B.n198 585
R289 B.n520 B.n519 585
R290 B.n517 B.n199 585
R291 B.n515 B.n514 585
R292 B.n513 B.n200 585
R293 B.n512 B.n511 585
R294 B.n509 B.n201 585
R295 B.n507 B.n506 585
R296 B.n505 B.n202 585
R297 B.n504 B.n503 585
R298 B.n501 B.n203 585
R299 B.n499 B.n498 585
R300 B.n497 B.n204 585
R301 B.n496 B.n495 585
R302 B.n493 B.n205 585
R303 B.n491 B.n490 585
R304 B.n489 B.n206 585
R305 B.n488 B.n487 585
R306 B.n485 B.n207 585
R307 B.n483 B.n482 585
R308 B.n481 B.n208 585
R309 B.n480 B.n479 585
R310 B.n477 B.n209 585
R311 B.n475 B.n474 585
R312 B.n473 B.n210 585
R313 B.n472 B.n471 585
R314 B.n469 B.n211 585
R315 B.n467 B.n466 585
R316 B.n465 B.n212 585
R317 B.n464 B.n463 585
R318 B.n461 B.n213 585
R319 B.n459 B.n458 585
R320 B.n457 B.n214 585
R321 B.n456 B.n455 585
R322 B.n453 B.n215 585
R323 B.n451 B.n450 585
R324 B.n449 B.n216 585
R325 B.n448 B.n447 585
R326 B.n445 B.n217 585
R327 B.n443 B.n442 585
R328 B.n441 B.n218 585
R329 B.n440 B.n439 585
R330 B.n437 B.n219 585
R331 B.n435 B.n434 585
R332 B.n433 B.n220 585
R333 B.n432 B.n431 585
R334 B.n429 B.n221 585
R335 B.n427 B.n426 585
R336 B.n425 B.n222 585
R337 B.n424 B.n423 585
R338 B.n421 B.n223 585
R339 B.n419 B.n418 585
R340 B.n417 B.n224 585
R341 B.n416 B.n415 585
R342 B.n413 B.n412 585
R343 B.n411 B.n410 585
R344 B.n409 B.n229 585
R345 B.n407 B.n406 585
R346 B.n405 B.n230 585
R347 B.n404 B.n403 585
R348 B.n401 B.n231 585
R349 B.n399 B.n398 585
R350 B.n397 B.n232 585
R351 B.n395 B.n394 585
R352 B.n392 B.n235 585
R353 B.n390 B.n389 585
R354 B.n388 B.n236 585
R355 B.n387 B.n386 585
R356 B.n384 B.n237 585
R357 B.n382 B.n381 585
R358 B.n380 B.n238 585
R359 B.n379 B.n378 585
R360 B.n376 B.n239 585
R361 B.n374 B.n373 585
R362 B.n372 B.n240 585
R363 B.n371 B.n370 585
R364 B.n368 B.n241 585
R365 B.n366 B.n365 585
R366 B.n364 B.n242 585
R367 B.n363 B.n362 585
R368 B.n360 B.n243 585
R369 B.n358 B.n357 585
R370 B.n356 B.n244 585
R371 B.n355 B.n354 585
R372 B.n352 B.n245 585
R373 B.n350 B.n349 585
R374 B.n348 B.n246 585
R375 B.n347 B.n346 585
R376 B.n344 B.n247 585
R377 B.n342 B.n341 585
R378 B.n340 B.n248 585
R379 B.n339 B.n338 585
R380 B.n336 B.n249 585
R381 B.n334 B.n333 585
R382 B.n332 B.n250 585
R383 B.n331 B.n330 585
R384 B.n328 B.n251 585
R385 B.n326 B.n325 585
R386 B.n324 B.n252 585
R387 B.n323 B.n322 585
R388 B.n320 B.n253 585
R389 B.n318 B.n317 585
R390 B.n316 B.n254 585
R391 B.n315 B.n314 585
R392 B.n312 B.n255 585
R393 B.n310 B.n309 585
R394 B.n308 B.n256 585
R395 B.n307 B.n306 585
R396 B.n304 B.n257 585
R397 B.n302 B.n301 585
R398 B.n300 B.n258 585
R399 B.n299 B.n298 585
R400 B.n296 B.n259 585
R401 B.n294 B.n293 585
R402 B.n292 B.n260 585
R403 B.n291 B.n290 585
R404 B.n288 B.n261 585
R405 B.n286 B.n285 585
R406 B.n284 B.n262 585
R407 B.n283 B.n282 585
R408 B.n280 B.n263 585
R409 B.n278 B.n277 585
R410 B.n276 B.n264 585
R411 B.n275 B.n274 585
R412 B.n272 B.n265 585
R413 B.n270 B.n269 585
R414 B.n268 B.n267 585
R415 B.n190 B.n189 585
R416 B.n544 B.n543 585
R417 B.n545 B.n544 585
R418 B.n186 B.n185 585
R419 B.n187 B.n186 585
R420 B.n553 B.n552 585
R421 B.n552 B.n551 585
R422 B.n554 B.n184 585
R423 B.n184 B.n183 585
R424 B.n556 B.n555 585
R425 B.n557 B.n556 585
R426 B.n178 B.n177 585
R427 B.n179 B.n178 585
R428 B.n565 B.n564 585
R429 B.n564 B.n563 585
R430 B.n566 B.n176 585
R431 B.n176 B.n175 585
R432 B.n568 B.n567 585
R433 B.n569 B.n568 585
R434 B.n170 B.n169 585
R435 B.n171 B.n170 585
R436 B.n577 B.n576 585
R437 B.n576 B.n575 585
R438 B.n578 B.n168 585
R439 B.n168 B.n167 585
R440 B.n580 B.n579 585
R441 B.n581 B.n580 585
R442 B.n162 B.n161 585
R443 B.n163 B.n162 585
R444 B.n589 B.n588 585
R445 B.n588 B.n587 585
R446 B.n590 B.n160 585
R447 B.n160 B.n159 585
R448 B.n592 B.n591 585
R449 B.n593 B.n592 585
R450 B.n154 B.n153 585
R451 B.n155 B.n154 585
R452 B.n601 B.n600 585
R453 B.n600 B.n599 585
R454 B.n602 B.n152 585
R455 B.n152 B.n151 585
R456 B.n604 B.n603 585
R457 B.n605 B.n604 585
R458 B.n146 B.n145 585
R459 B.n147 B.n146 585
R460 B.n613 B.n612 585
R461 B.n612 B.n611 585
R462 B.n614 B.n144 585
R463 B.n144 B.n143 585
R464 B.n616 B.n615 585
R465 B.n617 B.n616 585
R466 B.n138 B.n137 585
R467 B.n139 B.n138 585
R468 B.n626 B.n625 585
R469 B.n625 B.n624 585
R470 B.n627 B.n136 585
R471 B.n136 B.n135 585
R472 B.n629 B.n628 585
R473 B.n630 B.n629 585
R474 B.n2 B.n0 585
R475 B.n4 B.n2 585
R476 B.n3 B.n1 585
R477 B.n1009 B.n3 585
R478 B.n1007 B.n1006 585
R479 B.n1008 B.n1007 585
R480 B.n1005 B.n9 585
R481 B.n9 B.n8 585
R482 B.n1004 B.n1003 585
R483 B.n1003 B.n1002 585
R484 B.n11 B.n10 585
R485 B.n1001 B.n11 585
R486 B.n999 B.n998 585
R487 B.n1000 B.n999 585
R488 B.n997 B.n16 585
R489 B.n16 B.n15 585
R490 B.n996 B.n995 585
R491 B.n995 B.n994 585
R492 B.n18 B.n17 585
R493 B.n993 B.n18 585
R494 B.n991 B.n990 585
R495 B.n992 B.n991 585
R496 B.n989 B.n23 585
R497 B.n23 B.n22 585
R498 B.n988 B.n987 585
R499 B.n987 B.n986 585
R500 B.n25 B.n24 585
R501 B.n985 B.n25 585
R502 B.n983 B.n982 585
R503 B.n984 B.n983 585
R504 B.n981 B.n30 585
R505 B.n30 B.n29 585
R506 B.n980 B.n979 585
R507 B.n979 B.n978 585
R508 B.n32 B.n31 585
R509 B.n977 B.n32 585
R510 B.n975 B.n974 585
R511 B.n976 B.n975 585
R512 B.n973 B.n37 585
R513 B.n37 B.n36 585
R514 B.n972 B.n971 585
R515 B.n971 B.n970 585
R516 B.n39 B.n38 585
R517 B.n969 B.n39 585
R518 B.n967 B.n966 585
R519 B.n968 B.n967 585
R520 B.n965 B.n44 585
R521 B.n44 B.n43 585
R522 B.n964 B.n963 585
R523 B.n963 B.n962 585
R524 B.n46 B.n45 585
R525 B.n961 B.n46 585
R526 B.n959 B.n958 585
R527 B.n960 B.n959 585
R528 B.n957 B.n51 585
R529 B.n51 B.n50 585
R530 B.n956 B.n955 585
R531 B.n955 B.n954 585
R532 B.n53 B.n52 585
R533 B.n953 B.n53 585
R534 B.n951 B.n950 585
R535 B.n952 B.n951 585
R536 B.n1012 B.n1011 585
R537 B.n1011 B.n1010 585
R538 B.n544 B.n192 540.549
R539 B.n951 B.n58 540.549
R540 B.n546 B.n190 540.549
R541 B.n132 B.n56 540.549
R542 B.n233 B.t13 348.572
R543 B.n225 B.t2 348.572
R544 B.n91 B.t6 348.572
R545 B.n97 B.t10 348.572
R546 B.n675 B.n57 256.663
R547 B.n677 B.n57 256.663
R548 B.n683 B.n57 256.663
R549 B.n685 B.n57 256.663
R550 B.n691 B.n57 256.663
R551 B.n693 B.n57 256.663
R552 B.n699 B.n57 256.663
R553 B.n701 B.n57 256.663
R554 B.n707 B.n57 256.663
R555 B.n709 B.n57 256.663
R556 B.n715 B.n57 256.663
R557 B.n717 B.n57 256.663
R558 B.n723 B.n57 256.663
R559 B.n725 B.n57 256.663
R560 B.n731 B.n57 256.663
R561 B.n733 B.n57 256.663
R562 B.n739 B.n57 256.663
R563 B.n741 B.n57 256.663
R564 B.n747 B.n57 256.663
R565 B.n749 B.n57 256.663
R566 B.n755 B.n57 256.663
R567 B.n757 B.n57 256.663
R568 B.n763 B.n57 256.663
R569 B.n765 B.n57 256.663
R570 B.n771 B.n57 256.663
R571 B.n773 B.n57 256.663
R572 B.n779 B.n57 256.663
R573 B.n781 B.n57 256.663
R574 B.n787 B.n57 256.663
R575 B.n789 B.n57 256.663
R576 B.n795 B.n57 256.663
R577 B.n100 B.n57 256.663
R578 B.n801 B.n57 256.663
R579 B.n807 B.n57 256.663
R580 B.n809 B.n57 256.663
R581 B.n815 B.n57 256.663
R582 B.n817 B.n57 256.663
R583 B.n824 B.n57 256.663
R584 B.n826 B.n57 256.663
R585 B.n832 B.n57 256.663
R586 B.n834 B.n57 256.663
R587 B.n840 B.n57 256.663
R588 B.n842 B.n57 256.663
R589 B.n848 B.n57 256.663
R590 B.n850 B.n57 256.663
R591 B.n856 B.n57 256.663
R592 B.n858 B.n57 256.663
R593 B.n864 B.n57 256.663
R594 B.n866 B.n57 256.663
R595 B.n872 B.n57 256.663
R596 B.n874 B.n57 256.663
R597 B.n880 B.n57 256.663
R598 B.n882 B.n57 256.663
R599 B.n888 B.n57 256.663
R600 B.n890 B.n57 256.663
R601 B.n896 B.n57 256.663
R602 B.n898 B.n57 256.663
R603 B.n904 B.n57 256.663
R604 B.n906 B.n57 256.663
R605 B.n912 B.n57 256.663
R606 B.n914 B.n57 256.663
R607 B.n920 B.n57 256.663
R608 B.n922 B.n57 256.663
R609 B.n928 B.n57 256.663
R610 B.n930 B.n57 256.663
R611 B.n936 B.n57 256.663
R612 B.n938 B.n57 256.663
R613 B.n944 B.n57 256.663
R614 B.n946 B.n57 256.663
R615 B.n539 B.n191 256.663
R616 B.n194 B.n191 256.663
R617 B.n532 B.n191 256.663
R618 B.n526 B.n191 256.663
R619 B.n524 B.n191 256.663
R620 B.n518 B.n191 256.663
R621 B.n516 B.n191 256.663
R622 B.n510 B.n191 256.663
R623 B.n508 B.n191 256.663
R624 B.n502 B.n191 256.663
R625 B.n500 B.n191 256.663
R626 B.n494 B.n191 256.663
R627 B.n492 B.n191 256.663
R628 B.n486 B.n191 256.663
R629 B.n484 B.n191 256.663
R630 B.n478 B.n191 256.663
R631 B.n476 B.n191 256.663
R632 B.n470 B.n191 256.663
R633 B.n468 B.n191 256.663
R634 B.n462 B.n191 256.663
R635 B.n460 B.n191 256.663
R636 B.n454 B.n191 256.663
R637 B.n452 B.n191 256.663
R638 B.n446 B.n191 256.663
R639 B.n444 B.n191 256.663
R640 B.n438 B.n191 256.663
R641 B.n436 B.n191 256.663
R642 B.n430 B.n191 256.663
R643 B.n428 B.n191 256.663
R644 B.n422 B.n191 256.663
R645 B.n420 B.n191 256.663
R646 B.n414 B.n191 256.663
R647 B.n228 B.n191 256.663
R648 B.n408 B.n191 256.663
R649 B.n402 B.n191 256.663
R650 B.n400 B.n191 256.663
R651 B.n393 B.n191 256.663
R652 B.n391 B.n191 256.663
R653 B.n385 B.n191 256.663
R654 B.n383 B.n191 256.663
R655 B.n377 B.n191 256.663
R656 B.n375 B.n191 256.663
R657 B.n369 B.n191 256.663
R658 B.n367 B.n191 256.663
R659 B.n361 B.n191 256.663
R660 B.n359 B.n191 256.663
R661 B.n353 B.n191 256.663
R662 B.n351 B.n191 256.663
R663 B.n345 B.n191 256.663
R664 B.n343 B.n191 256.663
R665 B.n337 B.n191 256.663
R666 B.n335 B.n191 256.663
R667 B.n329 B.n191 256.663
R668 B.n327 B.n191 256.663
R669 B.n321 B.n191 256.663
R670 B.n319 B.n191 256.663
R671 B.n313 B.n191 256.663
R672 B.n311 B.n191 256.663
R673 B.n305 B.n191 256.663
R674 B.n303 B.n191 256.663
R675 B.n297 B.n191 256.663
R676 B.n295 B.n191 256.663
R677 B.n289 B.n191 256.663
R678 B.n287 B.n191 256.663
R679 B.n281 B.n191 256.663
R680 B.n279 B.n191 256.663
R681 B.n273 B.n191 256.663
R682 B.n271 B.n191 256.663
R683 B.n266 B.n191 256.663
R684 B.n544 B.n186 163.367
R685 B.n552 B.n186 163.367
R686 B.n552 B.n184 163.367
R687 B.n556 B.n184 163.367
R688 B.n556 B.n178 163.367
R689 B.n564 B.n178 163.367
R690 B.n564 B.n176 163.367
R691 B.n568 B.n176 163.367
R692 B.n568 B.n170 163.367
R693 B.n576 B.n170 163.367
R694 B.n576 B.n168 163.367
R695 B.n580 B.n168 163.367
R696 B.n580 B.n162 163.367
R697 B.n588 B.n162 163.367
R698 B.n588 B.n160 163.367
R699 B.n592 B.n160 163.367
R700 B.n592 B.n154 163.367
R701 B.n600 B.n154 163.367
R702 B.n600 B.n152 163.367
R703 B.n604 B.n152 163.367
R704 B.n604 B.n146 163.367
R705 B.n612 B.n146 163.367
R706 B.n612 B.n144 163.367
R707 B.n616 B.n144 163.367
R708 B.n616 B.n138 163.367
R709 B.n625 B.n138 163.367
R710 B.n625 B.n136 163.367
R711 B.n629 B.n136 163.367
R712 B.n629 B.n2 163.367
R713 B.n1011 B.n2 163.367
R714 B.n1011 B.n3 163.367
R715 B.n1007 B.n3 163.367
R716 B.n1007 B.n9 163.367
R717 B.n1003 B.n9 163.367
R718 B.n1003 B.n11 163.367
R719 B.n999 B.n11 163.367
R720 B.n999 B.n16 163.367
R721 B.n995 B.n16 163.367
R722 B.n995 B.n18 163.367
R723 B.n991 B.n18 163.367
R724 B.n991 B.n23 163.367
R725 B.n987 B.n23 163.367
R726 B.n987 B.n25 163.367
R727 B.n983 B.n25 163.367
R728 B.n983 B.n30 163.367
R729 B.n979 B.n30 163.367
R730 B.n979 B.n32 163.367
R731 B.n975 B.n32 163.367
R732 B.n975 B.n37 163.367
R733 B.n971 B.n37 163.367
R734 B.n971 B.n39 163.367
R735 B.n967 B.n39 163.367
R736 B.n967 B.n44 163.367
R737 B.n963 B.n44 163.367
R738 B.n963 B.n46 163.367
R739 B.n959 B.n46 163.367
R740 B.n959 B.n51 163.367
R741 B.n955 B.n51 163.367
R742 B.n955 B.n53 163.367
R743 B.n951 B.n53 163.367
R744 B.n540 B.n538 163.367
R745 B.n538 B.n537 163.367
R746 B.n534 B.n533 163.367
R747 B.n531 B.n196 163.367
R748 B.n527 B.n525 163.367
R749 B.n523 B.n198 163.367
R750 B.n519 B.n517 163.367
R751 B.n515 B.n200 163.367
R752 B.n511 B.n509 163.367
R753 B.n507 B.n202 163.367
R754 B.n503 B.n501 163.367
R755 B.n499 B.n204 163.367
R756 B.n495 B.n493 163.367
R757 B.n491 B.n206 163.367
R758 B.n487 B.n485 163.367
R759 B.n483 B.n208 163.367
R760 B.n479 B.n477 163.367
R761 B.n475 B.n210 163.367
R762 B.n471 B.n469 163.367
R763 B.n467 B.n212 163.367
R764 B.n463 B.n461 163.367
R765 B.n459 B.n214 163.367
R766 B.n455 B.n453 163.367
R767 B.n451 B.n216 163.367
R768 B.n447 B.n445 163.367
R769 B.n443 B.n218 163.367
R770 B.n439 B.n437 163.367
R771 B.n435 B.n220 163.367
R772 B.n431 B.n429 163.367
R773 B.n427 B.n222 163.367
R774 B.n423 B.n421 163.367
R775 B.n419 B.n224 163.367
R776 B.n415 B.n413 163.367
R777 B.n410 B.n409 163.367
R778 B.n407 B.n230 163.367
R779 B.n403 B.n401 163.367
R780 B.n399 B.n232 163.367
R781 B.n394 B.n392 163.367
R782 B.n390 B.n236 163.367
R783 B.n386 B.n384 163.367
R784 B.n382 B.n238 163.367
R785 B.n378 B.n376 163.367
R786 B.n374 B.n240 163.367
R787 B.n370 B.n368 163.367
R788 B.n366 B.n242 163.367
R789 B.n362 B.n360 163.367
R790 B.n358 B.n244 163.367
R791 B.n354 B.n352 163.367
R792 B.n350 B.n246 163.367
R793 B.n346 B.n344 163.367
R794 B.n342 B.n248 163.367
R795 B.n338 B.n336 163.367
R796 B.n334 B.n250 163.367
R797 B.n330 B.n328 163.367
R798 B.n326 B.n252 163.367
R799 B.n322 B.n320 163.367
R800 B.n318 B.n254 163.367
R801 B.n314 B.n312 163.367
R802 B.n310 B.n256 163.367
R803 B.n306 B.n304 163.367
R804 B.n302 B.n258 163.367
R805 B.n298 B.n296 163.367
R806 B.n294 B.n260 163.367
R807 B.n290 B.n288 163.367
R808 B.n286 B.n262 163.367
R809 B.n282 B.n280 163.367
R810 B.n278 B.n264 163.367
R811 B.n274 B.n272 163.367
R812 B.n270 B.n267 163.367
R813 B.n546 B.n188 163.367
R814 B.n550 B.n188 163.367
R815 B.n550 B.n182 163.367
R816 B.n558 B.n182 163.367
R817 B.n558 B.n180 163.367
R818 B.n562 B.n180 163.367
R819 B.n562 B.n174 163.367
R820 B.n570 B.n174 163.367
R821 B.n570 B.n172 163.367
R822 B.n574 B.n172 163.367
R823 B.n574 B.n166 163.367
R824 B.n582 B.n166 163.367
R825 B.n582 B.n164 163.367
R826 B.n586 B.n164 163.367
R827 B.n586 B.n158 163.367
R828 B.n594 B.n158 163.367
R829 B.n594 B.n156 163.367
R830 B.n598 B.n156 163.367
R831 B.n598 B.n150 163.367
R832 B.n606 B.n150 163.367
R833 B.n606 B.n148 163.367
R834 B.n610 B.n148 163.367
R835 B.n610 B.n142 163.367
R836 B.n618 B.n142 163.367
R837 B.n618 B.n140 163.367
R838 B.n623 B.n140 163.367
R839 B.n623 B.n134 163.367
R840 B.n631 B.n134 163.367
R841 B.n632 B.n631 163.367
R842 B.n632 B.n5 163.367
R843 B.n6 B.n5 163.367
R844 B.n7 B.n6 163.367
R845 B.n637 B.n7 163.367
R846 B.n637 B.n12 163.367
R847 B.n13 B.n12 163.367
R848 B.n14 B.n13 163.367
R849 B.n642 B.n14 163.367
R850 B.n642 B.n19 163.367
R851 B.n20 B.n19 163.367
R852 B.n21 B.n20 163.367
R853 B.n647 B.n21 163.367
R854 B.n647 B.n26 163.367
R855 B.n27 B.n26 163.367
R856 B.n28 B.n27 163.367
R857 B.n652 B.n28 163.367
R858 B.n652 B.n33 163.367
R859 B.n34 B.n33 163.367
R860 B.n35 B.n34 163.367
R861 B.n657 B.n35 163.367
R862 B.n657 B.n40 163.367
R863 B.n41 B.n40 163.367
R864 B.n42 B.n41 163.367
R865 B.n662 B.n42 163.367
R866 B.n662 B.n47 163.367
R867 B.n48 B.n47 163.367
R868 B.n49 B.n48 163.367
R869 B.n667 B.n49 163.367
R870 B.n667 B.n54 163.367
R871 B.n55 B.n54 163.367
R872 B.n56 B.n55 163.367
R873 B.n947 B.n945 163.367
R874 B.n943 B.n60 163.367
R875 B.n939 B.n937 163.367
R876 B.n935 B.n62 163.367
R877 B.n931 B.n929 163.367
R878 B.n927 B.n64 163.367
R879 B.n923 B.n921 163.367
R880 B.n919 B.n66 163.367
R881 B.n915 B.n913 163.367
R882 B.n911 B.n68 163.367
R883 B.n907 B.n905 163.367
R884 B.n903 B.n70 163.367
R885 B.n899 B.n897 163.367
R886 B.n895 B.n72 163.367
R887 B.n891 B.n889 163.367
R888 B.n887 B.n74 163.367
R889 B.n883 B.n881 163.367
R890 B.n879 B.n76 163.367
R891 B.n875 B.n873 163.367
R892 B.n871 B.n78 163.367
R893 B.n867 B.n865 163.367
R894 B.n863 B.n80 163.367
R895 B.n859 B.n857 163.367
R896 B.n855 B.n82 163.367
R897 B.n851 B.n849 163.367
R898 B.n847 B.n84 163.367
R899 B.n843 B.n841 163.367
R900 B.n839 B.n86 163.367
R901 B.n835 B.n833 163.367
R902 B.n831 B.n88 163.367
R903 B.n827 B.n825 163.367
R904 B.n823 B.n90 163.367
R905 B.n818 B.n816 163.367
R906 B.n814 B.n94 163.367
R907 B.n810 B.n808 163.367
R908 B.n806 B.n96 163.367
R909 B.n802 B.n800 163.367
R910 B.n797 B.n796 163.367
R911 B.n794 B.n102 163.367
R912 B.n790 B.n788 163.367
R913 B.n786 B.n104 163.367
R914 B.n782 B.n780 163.367
R915 B.n778 B.n106 163.367
R916 B.n774 B.n772 163.367
R917 B.n770 B.n108 163.367
R918 B.n766 B.n764 163.367
R919 B.n762 B.n110 163.367
R920 B.n758 B.n756 163.367
R921 B.n754 B.n112 163.367
R922 B.n750 B.n748 163.367
R923 B.n746 B.n114 163.367
R924 B.n742 B.n740 163.367
R925 B.n738 B.n116 163.367
R926 B.n734 B.n732 163.367
R927 B.n730 B.n118 163.367
R928 B.n726 B.n724 163.367
R929 B.n722 B.n120 163.367
R930 B.n718 B.n716 163.367
R931 B.n714 B.n122 163.367
R932 B.n710 B.n708 163.367
R933 B.n706 B.n124 163.367
R934 B.n702 B.n700 163.367
R935 B.n698 B.n126 163.367
R936 B.n694 B.n692 163.367
R937 B.n690 B.n128 163.367
R938 B.n686 B.n684 163.367
R939 B.n682 B.n130 163.367
R940 B.n678 B.n676 163.367
R941 B.n674 B.n132 163.367
R942 B.n233 B.t15 142.785
R943 B.n97 B.t11 142.785
R944 B.n225 B.t5 142.758
R945 B.n91 B.t8 142.758
R946 B.n234 B.n233 72.9217
R947 B.n226 B.n225 72.9217
R948 B.n92 B.n91 72.9217
R949 B.n98 B.n97 72.9217
R950 B.n539 B.n192 71.676
R951 B.n537 B.n194 71.676
R952 B.n533 B.n532 71.676
R953 B.n526 B.n196 71.676
R954 B.n525 B.n524 71.676
R955 B.n518 B.n198 71.676
R956 B.n517 B.n516 71.676
R957 B.n510 B.n200 71.676
R958 B.n509 B.n508 71.676
R959 B.n502 B.n202 71.676
R960 B.n501 B.n500 71.676
R961 B.n494 B.n204 71.676
R962 B.n493 B.n492 71.676
R963 B.n486 B.n206 71.676
R964 B.n485 B.n484 71.676
R965 B.n478 B.n208 71.676
R966 B.n477 B.n476 71.676
R967 B.n470 B.n210 71.676
R968 B.n469 B.n468 71.676
R969 B.n462 B.n212 71.676
R970 B.n461 B.n460 71.676
R971 B.n454 B.n214 71.676
R972 B.n453 B.n452 71.676
R973 B.n446 B.n216 71.676
R974 B.n445 B.n444 71.676
R975 B.n438 B.n218 71.676
R976 B.n437 B.n436 71.676
R977 B.n430 B.n220 71.676
R978 B.n429 B.n428 71.676
R979 B.n422 B.n222 71.676
R980 B.n421 B.n420 71.676
R981 B.n414 B.n224 71.676
R982 B.n413 B.n228 71.676
R983 B.n409 B.n408 71.676
R984 B.n402 B.n230 71.676
R985 B.n401 B.n400 71.676
R986 B.n393 B.n232 71.676
R987 B.n392 B.n391 71.676
R988 B.n385 B.n236 71.676
R989 B.n384 B.n383 71.676
R990 B.n377 B.n238 71.676
R991 B.n376 B.n375 71.676
R992 B.n369 B.n240 71.676
R993 B.n368 B.n367 71.676
R994 B.n361 B.n242 71.676
R995 B.n360 B.n359 71.676
R996 B.n353 B.n244 71.676
R997 B.n352 B.n351 71.676
R998 B.n345 B.n246 71.676
R999 B.n344 B.n343 71.676
R1000 B.n337 B.n248 71.676
R1001 B.n336 B.n335 71.676
R1002 B.n329 B.n250 71.676
R1003 B.n328 B.n327 71.676
R1004 B.n321 B.n252 71.676
R1005 B.n320 B.n319 71.676
R1006 B.n313 B.n254 71.676
R1007 B.n312 B.n311 71.676
R1008 B.n305 B.n256 71.676
R1009 B.n304 B.n303 71.676
R1010 B.n297 B.n258 71.676
R1011 B.n296 B.n295 71.676
R1012 B.n289 B.n260 71.676
R1013 B.n288 B.n287 71.676
R1014 B.n281 B.n262 71.676
R1015 B.n280 B.n279 71.676
R1016 B.n273 B.n264 71.676
R1017 B.n272 B.n271 71.676
R1018 B.n267 B.n266 71.676
R1019 B.n946 B.n58 71.676
R1020 B.n945 B.n944 71.676
R1021 B.n938 B.n60 71.676
R1022 B.n937 B.n936 71.676
R1023 B.n930 B.n62 71.676
R1024 B.n929 B.n928 71.676
R1025 B.n922 B.n64 71.676
R1026 B.n921 B.n920 71.676
R1027 B.n914 B.n66 71.676
R1028 B.n913 B.n912 71.676
R1029 B.n906 B.n68 71.676
R1030 B.n905 B.n904 71.676
R1031 B.n898 B.n70 71.676
R1032 B.n897 B.n896 71.676
R1033 B.n890 B.n72 71.676
R1034 B.n889 B.n888 71.676
R1035 B.n882 B.n74 71.676
R1036 B.n881 B.n880 71.676
R1037 B.n874 B.n76 71.676
R1038 B.n873 B.n872 71.676
R1039 B.n866 B.n78 71.676
R1040 B.n865 B.n864 71.676
R1041 B.n858 B.n80 71.676
R1042 B.n857 B.n856 71.676
R1043 B.n850 B.n82 71.676
R1044 B.n849 B.n848 71.676
R1045 B.n842 B.n84 71.676
R1046 B.n841 B.n840 71.676
R1047 B.n834 B.n86 71.676
R1048 B.n833 B.n832 71.676
R1049 B.n826 B.n88 71.676
R1050 B.n825 B.n824 71.676
R1051 B.n817 B.n90 71.676
R1052 B.n816 B.n815 71.676
R1053 B.n809 B.n94 71.676
R1054 B.n808 B.n807 71.676
R1055 B.n801 B.n96 71.676
R1056 B.n800 B.n100 71.676
R1057 B.n796 B.n795 71.676
R1058 B.n789 B.n102 71.676
R1059 B.n788 B.n787 71.676
R1060 B.n781 B.n104 71.676
R1061 B.n780 B.n779 71.676
R1062 B.n773 B.n106 71.676
R1063 B.n772 B.n771 71.676
R1064 B.n765 B.n108 71.676
R1065 B.n764 B.n763 71.676
R1066 B.n757 B.n110 71.676
R1067 B.n756 B.n755 71.676
R1068 B.n749 B.n112 71.676
R1069 B.n748 B.n747 71.676
R1070 B.n741 B.n114 71.676
R1071 B.n740 B.n739 71.676
R1072 B.n733 B.n116 71.676
R1073 B.n732 B.n731 71.676
R1074 B.n725 B.n118 71.676
R1075 B.n724 B.n723 71.676
R1076 B.n717 B.n120 71.676
R1077 B.n716 B.n715 71.676
R1078 B.n709 B.n122 71.676
R1079 B.n708 B.n707 71.676
R1080 B.n701 B.n124 71.676
R1081 B.n700 B.n699 71.676
R1082 B.n693 B.n126 71.676
R1083 B.n692 B.n691 71.676
R1084 B.n685 B.n128 71.676
R1085 B.n684 B.n683 71.676
R1086 B.n677 B.n130 71.676
R1087 B.n676 B.n675 71.676
R1088 B.n675 B.n674 71.676
R1089 B.n678 B.n677 71.676
R1090 B.n683 B.n682 71.676
R1091 B.n686 B.n685 71.676
R1092 B.n691 B.n690 71.676
R1093 B.n694 B.n693 71.676
R1094 B.n699 B.n698 71.676
R1095 B.n702 B.n701 71.676
R1096 B.n707 B.n706 71.676
R1097 B.n710 B.n709 71.676
R1098 B.n715 B.n714 71.676
R1099 B.n718 B.n717 71.676
R1100 B.n723 B.n722 71.676
R1101 B.n726 B.n725 71.676
R1102 B.n731 B.n730 71.676
R1103 B.n734 B.n733 71.676
R1104 B.n739 B.n738 71.676
R1105 B.n742 B.n741 71.676
R1106 B.n747 B.n746 71.676
R1107 B.n750 B.n749 71.676
R1108 B.n755 B.n754 71.676
R1109 B.n758 B.n757 71.676
R1110 B.n763 B.n762 71.676
R1111 B.n766 B.n765 71.676
R1112 B.n771 B.n770 71.676
R1113 B.n774 B.n773 71.676
R1114 B.n779 B.n778 71.676
R1115 B.n782 B.n781 71.676
R1116 B.n787 B.n786 71.676
R1117 B.n790 B.n789 71.676
R1118 B.n795 B.n794 71.676
R1119 B.n797 B.n100 71.676
R1120 B.n802 B.n801 71.676
R1121 B.n807 B.n806 71.676
R1122 B.n810 B.n809 71.676
R1123 B.n815 B.n814 71.676
R1124 B.n818 B.n817 71.676
R1125 B.n824 B.n823 71.676
R1126 B.n827 B.n826 71.676
R1127 B.n832 B.n831 71.676
R1128 B.n835 B.n834 71.676
R1129 B.n840 B.n839 71.676
R1130 B.n843 B.n842 71.676
R1131 B.n848 B.n847 71.676
R1132 B.n851 B.n850 71.676
R1133 B.n856 B.n855 71.676
R1134 B.n859 B.n858 71.676
R1135 B.n864 B.n863 71.676
R1136 B.n867 B.n866 71.676
R1137 B.n872 B.n871 71.676
R1138 B.n875 B.n874 71.676
R1139 B.n880 B.n879 71.676
R1140 B.n883 B.n882 71.676
R1141 B.n888 B.n887 71.676
R1142 B.n891 B.n890 71.676
R1143 B.n896 B.n895 71.676
R1144 B.n899 B.n898 71.676
R1145 B.n904 B.n903 71.676
R1146 B.n907 B.n906 71.676
R1147 B.n912 B.n911 71.676
R1148 B.n915 B.n914 71.676
R1149 B.n920 B.n919 71.676
R1150 B.n923 B.n922 71.676
R1151 B.n928 B.n927 71.676
R1152 B.n931 B.n930 71.676
R1153 B.n936 B.n935 71.676
R1154 B.n939 B.n938 71.676
R1155 B.n944 B.n943 71.676
R1156 B.n947 B.n946 71.676
R1157 B.n540 B.n539 71.676
R1158 B.n534 B.n194 71.676
R1159 B.n532 B.n531 71.676
R1160 B.n527 B.n526 71.676
R1161 B.n524 B.n523 71.676
R1162 B.n519 B.n518 71.676
R1163 B.n516 B.n515 71.676
R1164 B.n511 B.n510 71.676
R1165 B.n508 B.n507 71.676
R1166 B.n503 B.n502 71.676
R1167 B.n500 B.n499 71.676
R1168 B.n495 B.n494 71.676
R1169 B.n492 B.n491 71.676
R1170 B.n487 B.n486 71.676
R1171 B.n484 B.n483 71.676
R1172 B.n479 B.n478 71.676
R1173 B.n476 B.n475 71.676
R1174 B.n471 B.n470 71.676
R1175 B.n468 B.n467 71.676
R1176 B.n463 B.n462 71.676
R1177 B.n460 B.n459 71.676
R1178 B.n455 B.n454 71.676
R1179 B.n452 B.n451 71.676
R1180 B.n447 B.n446 71.676
R1181 B.n444 B.n443 71.676
R1182 B.n439 B.n438 71.676
R1183 B.n436 B.n435 71.676
R1184 B.n431 B.n430 71.676
R1185 B.n428 B.n427 71.676
R1186 B.n423 B.n422 71.676
R1187 B.n420 B.n419 71.676
R1188 B.n415 B.n414 71.676
R1189 B.n410 B.n228 71.676
R1190 B.n408 B.n407 71.676
R1191 B.n403 B.n402 71.676
R1192 B.n400 B.n399 71.676
R1193 B.n394 B.n393 71.676
R1194 B.n391 B.n390 71.676
R1195 B.n386 B.n385 71.676
R1196 B.n383 B.n382 71.676
R1197 B.n378 B.n377 71.676
R1198 B.n375 B.n374 71.676
R1199 B.n370 B.n369 71.676
R1200 B.n367 B.n366 71.676
R1201 B.n362 B.n361 71.676
R1202 B.n359 B.n358 71.676
R1203 B.n354 B.n353 71.676
R1204 B.n351 B.n350 71.676
R1205 B.n346 B.n345 71.676
R1206 B.n343 B.n342 71.676
R1207 B.n338 B.n337 71.676
R1208 B.n335 B.n334 71.676
R1209 B.n330 B.n329 71.676
R1210 B.n327 B.n326 71.676
R1211 B.n322 B.n321 71.676
R1212 B.n319 B.n318 71.676
R1213 B.n314 B.n313 71.676
R1214 B.n311 B.n310 71.676
R1215 B.n306 B.n305 71.676
R1216 B.n303 B.n302 71.676
R1217 B.n298 B.n297 71.676
R1218 B.n295 B.n294 71.676
R1219 B.n290 B.n289 71.676
R1220 B.n287 B.n286 71.676
R1221 B.n282 B.n281 71.676
R1222 B.n279 B.n278 71.676
R1223 B.n274 B.n273 71.676
R1224 B.n271 B.n270 71.676
R1225 B.n266 B.n190 71.676
R1226 B.n234 B.t14 69.8635
R1227 B.n98 B.t12 69.8635
R1228 B.n226 B.t4 69.8368
R1229 B.n92 B.t9 69.8368
R1230 B.n545 B.n191 60.832
R1231 B.n952 B.n57 60.832
R1232 B.n396 B.n234 59.5399
R1233 B.n227 B.n226 59.5399
R1234 B.n820 B.n92 59.5399
R1235 B.n99 B.n98 59.5399
R1236 B.n950 B.n949 35.1225
R1237 B.n672 B.n671 35.1225
R1238 B.n547 B.n189 35.1225
R1239 B.n543 B.n542 35.1225
R1240 B.n545 B.n187 29.7598
R1241 B.n551 B.n187 29.7598
R1242 B.n551 B.n183 29.7598
R1243 B.n557 B.n183 29.7598
R1244 B.n557 B.n179 29.7598
R1245 B.n563 B.n179 29.7598
R1246 B.n563 B.n175 29.7598
R1247 B.n569 B.n175 29.7598
R1248 B.n575 B.n171 29.7598
R1249 B.n575 B.n167 29.7598
R1250 B.n581 B.n167 29.7598
R1251 B.n581 B.n163 29.7598
R1252 B.n587 B.n163 29.7598
R1253 B.n587 B.n159 29.7598
R1254 B.n593 B.n159 29.7598
R1255 B.n593 B.n155 29.7598
R1256 B.n599 B.n155 29.7598
R1257 B.n599 B.n151 29.7598
R1258 B.n605 B.n151 29.7598
R1259 B.n605 B.n147 29.7598
R1260 B.n611 B.n147 29.7598
R1261 B.n617 B.n143 29.7598
R1262 B.n617 B.n139 29.7598
R1263 B.n624 B.n139 29.7598
R1264 B.n624 B.n135 29.7598
R1265 B.n630 B.n135 29.7598
R1266 B.n630 B.n4 29.7598
R1267 B.n1010 B.n4 29.7598
R1268 B.n1010 B.n1009 29.7598
R1269 B.n1009 B.n1008 29.7598
R1270 B.n1008 B.n8 29.7598
R1271 B.n1002 B.n8 29.7598
R1272 B.n1002 B.n1001 29.7598
R1273 B.n1001 B.n1000 29.7598
R1274 B.n1000 B.n15 29.7598
R1275 B.n994 B.n993 29.7598
R1276 B.n993 B.n992 29.7598
R1277 B.n992 B.n22 29.7598
R1278 B.n986 B.n22 29.7598
R1279 B.n986 B.n985 29.7598
R1280 B.n985 B.n984 29.7598
R1281 B.n984 B.n29 29.7598
R1282 B.n978 B.n29 29.7598
R1283 B.n978 B.n977 29.7598
R1284 B.n977 B.n976 29.7598
R1285 B.n976 B.n36 29.7598
R1286 B.n970 B.n36 29.7598
R1287 B.n970 B.n969 29.7598
R1288 B.n968 B.n43 29.7598
R1289 B.n962 B.n43 29.7598
R1290 B.n962 B.n961 29.7598
R1291 B.n961 B.n960 29.7598
R1292 B.n960 B.n50 29.7598
R1293 B.n954 B.n50 29.7598
R1294 B.n954 B.n953 29.7598
R1295 B.n953 B.n952 29.7598
R1296 B.n611 B.t1 25.8211
R1297 B.n994 B.t0 25.8211
R1298 B B.n1012 18.0485
R1299 B.n569 B.t3 17.9436
R1300 B.t7 B.n968 17.9436
R1301 B.t3 B.n171 11.8167
R1302 B.n969 B.t7 11.8167
R1303 B.n949 B.n948 10.6151
R1304 B.n948 B.n59 10.6151
R1305 B.n942 B.n59 10.6151
R1306 B.n942 B.n941 10.6151
R1307 B.n941 B.n940 10.6151
R1308 B.n940 B.n61 10.6151
R1309 B.n934 B.n61 10.6151
R1310 B.n934 B.n933 10.6151
R1311 B.n933 B.n932 10.6151
R1312 B.n932 B.n63 10.6151
R1313 B.n926 B.n63 10.6151
R1314 B.n926 B.n925 10.6151
R1315 B.n925 B.n924 10.6151
R1316 B.n924 B.n65 10.6151
R1317 B.n918 B.n65 10.6151
R1318 B.n918 B.n917 10.6151
R1319 B.n917 B.n916 10.6151
R1320 B.n916 B.n67 10.6151
R1321 B.n910 B.n67 10.6151
R1322 B.n910 B.n909 10.6151
R1323 B.n909 B.n908 10.6151
R1324 B.n908 B.n69 10.6151
R1325 B.n902 B.n69 10.6151
R1326 B.n902 B.n901 10.6151
R1327 B.n901 B.n900 10.6151
R1328 B.n900 B.n71 10.6151
R1329 B.n894 B.n71 10.6151
R1330 B.n894 B.n893 10.6151
R1331 B.n893 B.n892 10.6151
R1332 B.n892 B.n73 10.6151
R1333 B.n886 B.n73 10.6151
R1334 B.n886 B.n885 10.6151
R1335 B.n885 B.n884 10.6151
R1336 B.n884 B.n75 10.6151
R1337 B.n878 B.n75 10.6151
R1338 B.n878 B.n877 10.6151
R1339 B.n877 B.n876 10.6151
R1340 B.n876 B.n77 10.6151
R1341 B.n870 B.n77 10.6151
R1342 B.n870 B.n869 10.6151
R1343 B.n869 B.n868 10.6151
R1344 B.n868 B.n79 10.6151
R1345 B.n862 B.n79 10.6151
R1346 B.n862 B.n861 10.6151
R1347 B.n861 B.n860 10.6151
R1348 B.n860 B.n81 10.6151
R1349 B.n854 B.n81 10.6151
R1350 B.n854 B.n853 10.6151
R1351 B.n853 B.n852 10.6151
R1352 B.n852 B.n83 10.6151
R1353 B.n846 B.n83 10.6151
R1354 B.n846 B.n845 10.6151
R1355 B.n845 B.n844 10.6151
R1356 B.n844 B.n85 10.6151
R1357 B.n838 B.n85 10.6151
R1358 B.n838 B.n837 10.6151
R1359 B.n837 B.n836 10.6151
R1360 B.n836 B.n87 10.6151
R1361 B.n830 B.n87 10.6151
R1362 B.n830 B.n829 10.6151
R1363 B.n829 B.n828 10.6151
R1364 B.n828 B.n89 10.6151
R1365 B.n822 B.n89 10.6151
R1366 B.n822 B.n821 10.6151
R1367 B.n819 B.n93 10.6151
R1368 B.n813 B.n93 10.6151
R1369 B.n813 B.n812 10.6151
R1370 B.n812 B.n811 10.6151
R1371 B.n811 B.n95 10.6151
R1372 B.n805 B.n95 10.6151
R1373 B.n805 B.n804 10.6151
R1374 B.n804 B.n803 10.6151
R1375 B.n799 B.n798 10.6151
R1376 B.n798 B.n101 10.6151
R1377 B.n793 B.n101 10.6151
R1378 B.n793 B.n792 10.6151
R1379 B.n792 B.n791 10.6151
R1380 B.n791 B.n103 10.6151
R1381 B.n785 B.n103 10.6151
R1382 B.n785 B.n784 10.6151
R1383 B.n784 B.n783 10.6151
R1384 B.n783 B.n105 10.6151
R1385 B.n777 B.n105 10.6151
R1386 B.n777 B.n776 10.6151
R1387 B.n776 B.n775 10.6151
R1388 B.n775 B.n107 10.6151
R1389 B.n769 B.n107 10.6151
R1390 B.n769 B.n768 10.6151
R1391 B.n768 B.n767 10.6151
R1392 B.n767 B.n109 10.6151
R1393 B.n761 B.n109 10.6151
R1394 B.n761 B.n760 10.6151
R1395 B.n760 B.n759 10.6151
R1396 B.n759 B.n111 10.6151
R1397 B.n753 B.n111 10.6151
R1398 B.n753 B.n752 10.6151
R1399 B.n752 B.n751 10.6151
R1400 B.n751 B.n113 10.6151
R1401 B.n745 B.n113 10.6151
R1402 B.n745 B.n744 10.6151
R1403 B.n744 B.n743 10.6151
R1404 B.n743 B.n115 10.6151
R1405 B.n737 B.n115 10.6151
R1406 B.n737 B.n736 10.6151
R1407 B.n736 B.n735 10.6151
R1408 B.n735 B.n117 10.6151
R1409 B.n729 B.n117 10.6151
R1410 B.n729 B.n728 10.6151
R1411 B.n728 B.n727 10.6151
R1412 B.n727 B.n119 10.6151
R1413 B.n721 B.n119 10.6151
R1414 B.n721 B.n720 10.6151
R1415 B.n720 B.n719 10.6151
R1416 B.n719 B.n121 10.6151
R1417 B.n713 B.n121 10.6151
R1418 B.n713 B.n712 10.6151
R1419 B.n712 B.n711 10.6151
R1420 B.n711 B.n123 10.6151
R1421 B.n705 B.n123 10.6151
R1422 B.n705 B.n704 10.6151
R1423 B.n704 B.n703 10.6151
R1424 B.n703 B.n125 10.6151
R1425 B.n697 B.n125 10.6151
R1426 B.n697 B.n696 10.6151
R1427 B.n696 B.n695 10.6151
R1428 B.n695 B.n127 10.6151
R1429 B.n689 B.n127 10.6151
R1430 B.n689 B.n688 10.6151
R1431 B.n688 B.n687 10.6151
R1432 B.n687 B.n129 10.6151
R1433 B.n681 B.n129 10.6151
R1434 B.n681 B.n680 10.6151
R1435 B.n680 B.n679 10.6151
R1436 B.n679 B.n131 10.6151
R1437 B.n673 B.n131 10.6151
R1438 B.n673 B.n672 10.6151
R1439 B.n548 B.n547 10.6151
R1440 B.n549 B.n548 10.6151
R1441 B.n549 B.n181 10.6151
R1442 B.n559 B.n181 10.6151
R1443 B.n560 B.n559 10.6151
R1444 B.n561 B.n560 10.6151
R1445 B.n561 B.n173 10.6151
R1446 B.n571 B.n173 10.6151
R1447 B.n572 B.n571 10.6151
R1448 B.n573 B.n572 10.6151
R1449 B.n573 B.n165 10.6151
R1450 B.n583 B.n165 10.6151
R1451 B.n584 B.n583 10.6151
R1452 B.n585 B.n584 10.6151
R1453 B.n585 B.n157 10.6151
R1454 B.n595 B.n157 10.6151
R1455 B.n596 B.n595 10.6151
R1456 B.n597 B.n596 10.6151
R1457 B.n597 B.n149 10.6151
R1458 B.n607 B.n149 10.6151
R1459 B.n608 B.n607 10.6151
R1460 B.n609 B.n608 10.6151
R1461 B.n609 B.n141 10.6151
R1462 B.n619 B.n141 10.6151
R1463 B.n620 B.n619 10.6151
R1464 B.n622 B.n620 10.6151
R1465 B.n622 B.n621 10.6151
R1466 B.n621 B.n133 10.6151
R1467 B.n633 B.n133 10.6151
R1468 B.n634 B.n633 10.6151
R1469 B.n635 B.n634 10.6151
R1470 B.n636 B.n635 10.6151
R1471 B.n638 B.n636 10.6151
R1472 B.n639 B.n638 10.6151
R1473 B.n640 B.n639 10.6151
R1474 B.n641 B.n640 10.6151
R1475 B.n643 B.n641 10.6151
R1476 B.n644 B.n643 10.6151
R1477 B.n645 B.n644 10.6151
R1478 B.n646 B.n645 10.6151
R1479 B.n648 B.n646 10.6151
R1480 B.n649 B.n648 10.6151
R1481 B.n650 B.n649 10.6151
R1482 B.n651 B.n650 10.6151
R1483 B.n653 B.n651 10.6151
R1484 B.n654 B.n653 10.6151
R1485 B.n655 B.n654 10.6151
R1486 B.n656 B.n655 10.6151
R1487 B.n658 B.n656 10.6151
R1488 B.n659 B.n658 10.6151
R1489 B.n660 B.n659 10.6151
R1490 B.n661 B.n660 10.6151
R1491 B.n663 B.n661 10.6151
R1492 B.n664 B.n663 10.6151
R1493 B.n665 B.n664 10.6151
R1494 B.n666 B.n665 10.6151
R1495 B.n668 B.n666 10.6151
R1496 B.n669 B.n668 10.6151
R1497 B.n670 B.n669 10.6151
R1498 B.n671 B.n670 10.6151
R1499 B.n542 B.n541 10.6151
R1500 B.n541 B.n193 10.6151
R1501 B.n536 B.n193 10.6151
R1502 B.n536 B.n535 10.6151
R1503 B.n535 B.n195 10.6151
R1504 B.n530 B.n195 10.6151
R1505 B.n530 B.n529 10.6151
R1506 B.n529 B.n528 10.6151
R1507 B.n528 B.n197 10.6151
R1508 B.n522 B.n197 10.6151
R1509 B.n522 B.n521 10.6151
R1510 B.n521 B.n520 10.6151
R1511 B.n520 B.n199 10.6151
R1512 B.n514 B.n199 10.6151
R1513 B.n514 B.n513 10.6151
R1514 B.n513 B.n512 10.6151
R1515 B.n512 B.n201 10.6151
R1516 B.n506 B.n201 10.6151
R1517 B.n506 B.n505 10.6151
R1518 B.n505 B.n504 10.6151
R1519 B.n504 B.n203 10.6151
R1520 B.n498 B.n203 10.6151
R1521 B.n498 B.n497 10.6151
R1522 B.n497 B.n496 10.6151
R1523 B.n496 B.n205 10.6151
R1524 B.n490 B.n205 10.6151
R1525 B.n490 B.n489 10.6151
R1526 B.n489 B.n488 10.6151
R1527 B.n488 B.n207 10.6151
R1528 B.n482 B.n207 10.6151
R1529 B.n482 B.n481 10.6151
R1530 B.n481 B.n480 10.6151
R1531 B.n480 B.n209 10.6151
R1532 B.n474 B.n209 10.6151
R1533 B.n474 B.n473 10.6151
R1534 B.n473 B.n472 10.6151
R1535 B.n472 B.n211 10.6151
R1536 B.n466 B.n211 10.6151
R1537 B.n466 B.n465 10.6151
R1538 B.n465 B.n464 10.6151
R1539 B.n464 B.n213 10.6151
R1540 B.n458 B.n213 10.6151
R1541 B.n458 B.n457 10.6151
R1542 B.n457 B.n456 10.6151
R1543 B.n456 B.n215 10.6151
R1544 B.n450 B.n215 10.6151
R1545 B.n450 B.n449 10.6151
R1546 B.n449 B.n448 10.6151
R1547 B.n448 B.n217 10.6151
R1548 B.n442 B.n217 10.6151
R1549 B.n442 B.n441 10.6151
R1550 B.n441 B.n440 10.6151
R1551 B.n440 B.n219 10.6151
R1552 B.n434 B.n219 10.6151
R1553 B.n434 B.n433 10.6151
R1554 B.n433 B.n432 10.6151
R1555 B.n432 B.n221 10.6151
R1556 B.n426 B.n221 10.6151
R1557 B.n426 B.n425 10.6151
R1558 B.n425 B.n424 10.6151
R1559 B.n424 B.n223 10.6151
R1560 B.n418 B.n223 10.6151
R1561 B.n418 B.n417 10.6151
R1562 B.n417 B.n416 10.6151
R1563 B.n412 B.n411 10.6151
R1564 B.n411 B.n229 10.6151
R1565 B.n406 B.n229 10.6151
R1566 B.n406 B.n405 10.6151
R1567 B.n405 B.n404 10.6151
R1568 B.n404 B.n231 10.6151
R1569 B.n398 B.n231 10.6151
R1570 B.n398 B.n397 10.6151
R1571 B.n395 B.n235 10.6151
R1572 B.n389 B.n235 10.6151
R1573 B.n389 B.n388 10.6151
R1574 B.n388 B.n387 10.6151
R1575 B.n387 B.n237 10.6151
R1576 B.n381 B.n237 10.6151
R1577 B.n381 B.n380 10.6151
R1578 B.n380 B.n379 10.6151
R1579 B.n379 B.n239 10.6151
R1580 B.n373 B.n239 10.6151
R1581 B.n373 B.n372 10.6151
R1582 B.n372 B.n371 10.6151
R1583 B.n371 B.n241 10.6151
R1584 B.n365 B.n241 10.6151
R1585 B.n365 B.n364 10.6151
R1586 B.n364 B.n363 10.6151
R1587 B.n363 B.n243 10.6151
R1588 B.n357 B.n243 10.6151
R1589 B.n357 B.n356 10.6151
R1590 B.n356 B.n355 10.6151
R1591 B.n355 B.n245 10.6151
R1592 B.n349 B.n245 10.6151
R1593 B.n349 B.n348 10.6151
R1594 B.n348 B.n347 10.6151
R1595 B.n347 B.n247 10.6151
R1596 B.n341 B.n247 10.6151
R1597 B.n341 B.n340 10.6151
R1598 B.n340 B.n339 10.6151
R1599 B.n339 B.n249 10.6151
R1600 B.n333 B.n249 10.6151
R1601 B.n333 B.n332 10.6151
R1602 B.n332 B.n331 10.6151
R1603 B.n331 B.n251 10.6151
R1604 B.n325 B.n251 10.6151
R1605 B.n325 B.n324 10.6151
R1606 B.n324 B.n323 10.6151
R1607 B.n323 B.n253 10.6151
R1608 B.n317 B.n253 10.6151
R1609 B.n317 B.n316 10.6151
R1610 B.n316 B.n315 10.6151
R1611 B.n315 B.n255 10.6151
R1612 B.n309 B.n255 10.6151
R1613 B.n309 B.n308 10.6151
R1614 B.n308 B.n307 10.6151
R1615 B.n307 B.n257 10.6151
R1616 B.n301 B.n257 10.6151
R1617 B.n301 B.n300 10.6151
R1618 B.n300 B.n299 10.6151
R1619 B.n299 B.n259 10.6151
R1620 B.n293 B.n259 10.6151
R1621 B.n293 B.n292 10.6151
R1622 B.n292 B.n291 10.6151
R1623 B.n291 B.n261 10.6151
R1624 B.n285 B.n261 10.6151
R1625 B.n285 B.n284 10.6151
R1626 B.n284 B.n283 10.6151
R1627 B.n283 B.n263 10.6151
R1628 B.n277 B.n263 10.6151
R1629 B.n277 B.n276 10.6151
R1630 B.n276 B.n275 10.6151
R1631 B.n275 B.n265 10.6151
R1632 B.n269 B.n265 10.6151
R1633 B.n269 B.n268 10.6151
R1634 B.n268 B.n189 10.6151
R1635 B.n543 B.n185 10.6151
R1636 B.n553 B.n185 10.6151
R1637 B.n554 B.n553 10.6151
R1638 B.n555 B.n554 10.6151
R1639 B.n555 B.n177 10.6151
R1640 B.n565 B.n177 10.6151
R1641 B.n566 B.n565 10.6151
R1642 B.n567 B.n566 10.6151
R1643 B.n567 B.n169 10.6151
R1644 B.n577 B.n169 10.6151
R1645 B.n578 B.n577 10.6151
R1646 B.n579 B.n578 10.6151
R1647 B.n579 B.n161 10.6151
R1648 B.n589 B.n161 10.6151
R1649 B.n590 B.n589 10.6151
R1650 B.n591 B.n590 10.6151
R1651 B.n591 B.n153 10.6151
R1652 B.n601 B.n153 10.6151
R1653 B.n602 B.n601 10.6151
R1654 B.n603 B.n602 10.6151
R1655 B.n603 B.n145 10.6151
R1656 B.n613 B.n145 10.6151
R1657 B.n614 B.n613 10.6151
R1658 B.n615 B.n614 10.6151
R1659 B.n615 B.n137 10.6151
R1660 B.n626 B.n137 10.6151
R1661 B.n627 B.n626 10.6151
R1662 B.n628 B.n627 10.6151
R1663 B.n628 B.n0 10.6151
R1664 B.n1006 B.n1 10.6151
R1665 B.n1006 B.n1005 10.6151
R1666 B.n1005 B.n1004 10.6151
R1667 B.n1004 B.n10 10.6151
R1668 B.n998 B.n10 10.6151
R1669 B.n998 B.n997 10.6151
R1670 B.n997 B.n996 10.6151
R1671 B.n996 B.n17 10.6151
R1672 B.n990 B.n17 10.6151
R1673 B.n990 B.n989 10.6151
R1674 B.n989 B.n988 10.6151
R1675 B.n988 B.n24 10.6151
R1676 B.n982 B.n24 10.6151
R1677 B.n982 B.n981 10.6151
R1678 B.n981 B.n980 10.6151
R1679 B.n980 B.n31 10.6151
R1680 B.n974 B.n31 10.6151
R1681 B.n974 B.n973 10.6151
R1682 B.n973 B.n972 10.6151
R1683 B.n972 B.n38 10.6151
R1684 B.n966 B.n38 10.6151
R1685 B.n966 B.n965 10.6151
R1686 B.n965 B.n964 10.6151
R1687 B.n964 B.n45 10.6151
R1688 B.n958 B.n45 10.6151
R1689 B.n958 B.n957 10.6151
R1690 B.n957 B.n956 10.6151
R1691 B.n956 B.n52 10.6151
R1692 B.n950 B.n52 10.6151
R1693 B.n820 B.n819 6.5566
R1694 B.n803 B.n99 6.5566
R1695 B.n412 B.n227 6.5566
R1696 B.n397 B.n396 6.5566
R1697 B.n821 B.n820 4.05904
R1698 B.n799 B.n99 4.05904
R1699 B.n416 B.n227 4.05904
R1700 B.n396 B.n395 4.05904
R1701 B.t1 B.n143 3.93923
R1702 B.t0 B.n15 3.93923
R1703 B.n1012 B.n0 2.81026
R1704 B.n1012 B.n1 2.81026
R1705 VN VN.t0 231.107
R1706 VN VN.t1 178.913
R1707 VDD2.n0 VDD2.t0 111.956
R1708 VDD2.n0 VDD2.t1 64.6925
R1709 VDD2 VDD2.n0 0.869035
C0 VDD1 VN 0.148837f
C1 VN VTAIL 3.96269f
C2 VN VDD2 4.61154f
C3 VDD1 VTAIL 7.20965f
C4 VP VN 7.297141f
C5 VDD1 VDD2 0.776627f
C6 VTAIL VDD2 7.26518f
C7 VDD1 VP 4.8282f
C8 VP VTAIL 3.97701f
C9 VP VDD2 0.368773f
C10 VDD2 B 6.126414f
C11 VDD1 B 9.986441f
C12 VTAIL B 10.988797f
C13 VN B 13.34007f
C14 VP B 7.955465f
C15 VDD2.t0 B 4.46342f
C16 VDD2.t1 B 3.67462f
C17 VDD2.n0 B 3.60125f
C18 VN.t1 B 4.93931f
C19 VN.t0 B 5.61736f
C20 VDD1.t1 B 3.68635f
C21 VDD1.t0 B 4.51943f
C22 VTAIL.t3 B 3.567f
C23 VTAIL.n0 B 2.11334f
C24 VTAIL.t1 B 3.567f
C25 VTAIL.n1 B 2.16126f
C26 VTAIL.t2 B 3.567f
C27 VTAIL.n2 B 1.95474f
C28 VTAIL.t0 B 3.567f
C29 VTAIL.n3 B 1.86947f
C30 VP.t0 B 5.70065f
C31 VP.t1 B 5.0076f
C32 VP.n0 B 5.3019f
.ends

