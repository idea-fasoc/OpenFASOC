* NGSPICE file created from diff_pair_sample_1498.ext - technology: sky130A

.subckt diff_pair_sample_1498 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t1 VP.t0 VTAIL.t3 B.t0 sky130_fd_pr__nfet_01v8 ad=2.5194 pd=13.7 as=2.5194 ps=13.7 w=6.46 l=1.55
X1 VDD1.t0 VP.t1 VTAIL.t2 B.t1 sky130_fd_pr__nfet_01v8 ad=2.5194 pd=13.7 as=2.5194 ps=13.7 w=6.46 l=1.55
X2 B.t15 B.t13 B.t14 B.t10 sky130_fd_pr__nfet_01v8 ad=2.5194 pd=13.7 as=0 ps=0 w=6.46 l=1.55
X3 B.t12 B.t9 B.t11 B.t10 sky130_fd_pr__nfet_01v8 ad=2.5194 pd=13.7 as=0 ps=0 w=6.46 l=1.55
X4 VDD2.t1 VN.t0 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=2.5194 pd=13.7 as=2.5194 ps=13.7 w=6.46 l=1.55
X5 B.t8 B.t6 B.t7 B.t3 sky130_fd_pr__nfet_01v8 ad=2.5194 pd=13.7 as=0 ps=0 w=6.46 l=1.55
X6 B.t5 B.t2 B.t4 B.t3 sky130_fd_pr__nfet_01v8 ad=2.5194 pd=13.7 as=0 ps=0 w=6.46 l=1.55
X7 VDD2.t0 VN.t1 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=2.5194 pd=13.7 as=2.5194 ps=13.7 w=6.46 l=1.55
R0 VP.n0 VP.t1 244.065
R1 VP.n0 VP.t0 206.391
R2 VP VP.n0 0.146778
R3 VTAIL.n134 VTAIL.n133 289.615
R4 VTAIL.n32 VTAIL.n31 289.615
R5 VTAIL.n100 VTAIL.n99 289.615
R6 VTAIL.n66 VTAIL.n65 289.615
R7 VTAIL.n112 VTAIL.n111 185
R8 VTAIL.n117 VTAIL.n116 185
R9 VTAIL.n119 VTAIL.n118 185
R10 VTAIL.n108 VTAIL.n107 185
R11 VTAIL.n125 VTAIL.n124 185
R12 VTAIL.n127 VTAIL.n126 185
R13 VTAIL.n104 VTAIL.n103 185
R14 VTAIL.n133 VTAIL.n132 185
R15 VTAIL.n10 VTAIL.n9 185
R16 VTAIL.n15 VTAIL.n14 185
R17 VTAIL.n17 VTAIL.n16 185
R18 VTAIL.n6 VTAIL.n5 185
R19 VTAIL.n23 VTAIL.n22 185
R20 VTAIL.n25 VTAIL.n24 185
R21 VTAIL.n2 VTAIL.n1 185
R22 VTAIL.n31 VTAIL.n30 185
R23 VTAIL.n99 VTAIL.n98 185
R24 VTAIL.n70 VTAIL.n69 185
R25 VTAIL.n93 VTAIL.n92 185
R26 VTAIL.n91 VTAIL.n90 185
R27 VTAIL.n74 VTAIL.n73 185
R28 VTAIL.n85 VTAIL.n84 185
R29 VTAIL.n83 VTAIL.n82 185
R30 VTAIL.n78 VTAIL.n77 185
R31 VTAIL.n65 VTAIL.n64 185
R32 VTAIL.n36 VTAIL.n35 185
R33 VTAIL.n59 VTAIL.n58 185
R34 VTAIL.n57 VTAIL.n56 185
R35 VTAIL.n40 VTAIL.n39 185
R36 VTAIL.n51 VTAIL.n50 185
R37 VTAIL.n49 VTAIL.n48 185
R38 VTAIL.n44 VTAIL.n43 185
R39 VTAIL.n45 VTAIL.t0 149.525
R40 VTAIL.n113 VTAIL.t1 149.525
R41 VTAIL.n11 VTAIL.t3 149.525
R42 VTAIL.n79 VTAIL.t2 149.525
R43 VTAIL.n117 VTAIL.n111 104.615
R44 VTAIL.n118 VTAIL.n117 104.615
R45 VTAIL.n118 VTAIL.n107 104.615
R46 VTAIL.n125 VTAIL.n107 104.615
R47 VTAIL.n126 VTAIL.n125 104.615
R48 VTAIL.n126 VTAIL.n103 104.615
R49 VTAIL.n133 VTAIL.n103 104.615
R50 VTAIL.n15 VTAIL.n9 104.615
R51 VTAIL.n16 VTAIL.n15 104.615
R52 VTAIL.n16 VTAIL.n5 104.615
R53 VTAIL.n23 VTAIL.n5 104.615
R54 VTAIL.n24 VTAIL.n23 104.615
R55 VTAIL.n24 VTAIL.n1 104.615
R56 VTAIL.n31 VTAIL.n1 104.615
R57 VTAIL.n99 VTAIL.n69 104.615
R58 VTAIL.n92 VTAIL.n69 104.615
R59 VTAIL.n92 VTAIL.n91 104.615
R60 VTAIL.n91 VTAIL.n73 104.615
R61 VTAIL.n84 VTAIL.n73 104.615
R62 VTAIL.n84 VTAIL.n83 104.615
R63 VTAIL.n83 VTAIL.n77 104.615
R64 VTAIL.n65 VTAIL.n35 104.615
R65 VTAIL.n58 VTAIL.n35 104.615
R66 VTAIL.n58 VTAIL.n57 104.615
R67 VTAIL.n57 VTAIL.n39 104.615
R68 VTAIL.n50 VTAIL.n39 104.615
R69 VTAIL.n50 VTAIL.n49 104.615
R70 VTAIL.n49 VTAIL.n43 104.615
R71 VTAIL.t1 VTAIL.n111 52.3082
R72 VTAIL.t3 VTAIL.n9 52.3082
R73 VTAIL.t2 VTAIL.n77 52.3082
R74 VTAIL.t0 VTAIL.n43 52.3082
R75 VTAIL.n135 VTAIL.n134 33.7369
R76 VTAIL.n33 VTAIL.n32 33.7369
R77 VTAIL.n101 VTAIL.n100 33.7369
R78 VTAIL.n67 VTAIL.n66 33.7369
R79 VTAIL.n67 VTAIL.n33 21.1772
R80 VTAIL.n135 VTAIL.n101 19.5565
R81 VTAIL.n132 VTAIL.n102 12.8005
R82 VTAIL.n30 VTAIL.n0 12.8005
R83 VTAIL.n98 VTAIL.n68 12.8005
R84 VTAIL.n64 VTAIL.n34 12.8005
R85 VTAIL.n131 VTAIL.n104 12.0247
R86 VTAIL.n29 VTAIL.n2 12.0247
R87 VTAIL.n97 VTAIL.n70 12.0247
R88 VTAIL.n63 VTAIL.n36 12.0247
R89 VTAIL.n128 VTAIL.n127 11.249
R90 VTAIL.n26 VTAIL.n25 11.249
R91 VTAIL.n94 VTAIL.n93 11.249
R92 VTAIL.n60 VTAIL.n59 11.249
R93 VTAIL.n124 VTAIL.n106 10.4732
R94 VTAIL.n22 VTAIL.n4 10.4732
R95 VTAIL.n90 VTAIL.n72 10.4732
R96 VTAIL.n56 VTAIL.n38 10.4732
R97 VTAIL.n113 VTAIL.n112 10.2746
R98 VTAIL.n11 VTAIL.n10 10.2746
R99 VTAIL.n79 VTAIL.n78 10.2746
R100 VTAIL.n45 VTAIL.n44 10.2746
R101 VTAIL.n123 VTAIL.n108 9.69747
R102 VTAIL.n21 VTAIL.n6 9.69747
R103 VTAIL.n89 VTAIL.n74 9.69747
R104 VTAIL.n55 VTAIL.n40 9.69747
R105 VTAIL.n130 VTAIL.n102 9.45567
R106 VTAIL.n28 VTAIL.n0 9.45567
R107 VTAIL.n96 VTAIL.n68 9.45567
R108 VTAIL.n62 VTAIL.n34 9.45567
R109 VTAIL.n115 VTAIL.n114 9.3005
R110 VTAIL.n110 VTAIL.n109 9.3005
R111 VTAIL.n121 VTAIL.n120 9.3005
R112 VTAIL.n123 VTAIL.n122 9.3005
R113 VTAIL.n106 VTAIL.n105 9.3005
R114 VTAIL.n129 VTAIL.n128 9.3005
R115 VTAIL.n131 VTAIL.n130 9.3005
R116 VTAIL.n13 VTAIL.n12 9.3005
R117 VTAIL.n8 VTAIL.n7 9.3005
R118 VTAIL.n19 VTAIL.n18 9.3005
R119 VTAIL.n21 VTAIL.n20 9.3005
R120 VTAIL.n4 VTAIL.n3 9.3005
R121 VTAIL.n27 VTAIL.n26 9.3005
R122 VTAIL.n29 VTAIL.n28 9.3005
R123 VTAIL.n97 VTAIL.n96 9.3005
R124 VTAIL.n95 VTAIL.n94 9.3005
R125 VTAIL.n72 VTAIL.n71 9.3005
R126 VTAIL.n89 VTAIL.n88 9.3005
R127 VTAIL.n87 VTAIL.n86 9.3005
R128 VTAIL.n76 VTAIL.n75 9.3005
R129 VTAIL.n81 VTAIL.n80 9.3005
R130 VTAIL.n42 VTAIL.n41 9.3005
R131 VTAIL.n53 VTAIL.n52 9.3005
R132 VTAIL.n55 VTAIL.n54 9.3005
R133 VTAIL.n38 VTAIL.n37 9.3005
R134 VTAIL.n61 VTAIL.n60 9.3005
R135 VTAIL.n63 VTAIL.n62 9.3005
R136 VTAIL.n47 VTAIL.n46 9.3005
R137 VTAIL.n120 VTAIL.n119 8.92171
R138 VTAIL.n18 VTAIL.n17 8.92171
R139 VTAIL.n86 VTAIL.n85 8.92171
R140 VTAIL.n52 VTAIL.n51 8.92171
R141 VTAIL.n116 VTAIL.n110 8.14595
R142 VTAIL.n14 VTAIL.n8 8.14595
R143 VTAIL.n82 VTAIL.n76 8.14595
R144 VTAIL.n48 VTAIL.n42 8.14595
R145 VTAIL.n115 VTAIL.n112 7.3702
R146 VTAIL.n13 VTAIL.n10 7.3702
R147 VTAIL.n81 VTAIL.n78 7.3702
R148 VTAIL.n47 VTAIL.n44 7.3702
R149 VTAIL.n116 VTAIL.n115 5.81868
R150 VTAIL.n14 VTAIL.n13 5.81868
R151 VTAIL.n82 VTAIL.n81 5.81868
R152 VTAIL.n48 VTAIL.n47 5.81868
R153 VTAIL.n119 VTAIL.n110 5.04292
R154 VTAIL.n17 VTAIL.n8 5.04292
R155 VTAIL.n85 VTAIL.n76 5.04292
R156 VTAIL.n51 VTAIL.n42 5.04292
R157 VTAIL.n120 VTAIL.n108 4.26717
R158 VTAIL.n18 VTAIL.n6 4.26717
R159 VTAIL.n86 VTAIL.n74 4.26717
R160 VTAIL.n52 VTAIL.n40 4.26717
R161 VTAIL.n124 VTAIL.n123 3.49141
R162 VTAIL.n22 VTAIL.n21 3.49141
R163 VTAIL.n90 VTAIL.n89 3.49141
R164 VTAIL.n56 VTAIL.n55 3.49141
R165 VTAIL.n46 VTAIL.n45 2.84308
R166 VTAIL.n114 VTAIL.n113 2.84308
R167 VTAIL.n12 VTAIL.n11 2.84308
R168 VTAIL.n80 VTAIL.n79 2.84308
R169 VTAIL.n127 VTAIL.n106 2.71565
R170 VTAIL.n25 VTAIL.n4 2.71565
R171 VTAIL.n93 VTAIL.n72 2.71565
R172 VTAIL.n59 VTAIL.n38 2.71565
R173 VTAIL.n128 VTAIL.n104 1.93989
R174 VTAIL.n26 VTAIL.n2 1.93989
R175 VTAIL.n94 VTAIL.n70 1.93989
R176 VTAIL.n60 VTAIL.n36 1.93989
R177 VTAIL.n101 VTAIL.n67 1.28067
R178 VTAIL.n132 VTAIL.n131 1.16414
R179 VTAIL.n30 VTAIL.n29 1.16414
R180 VTAIL.n98 VTAIL.n97 1.16414
R181 VTAIL.n64 VTAIL.n63 1.16414
R182 VTAIL VTAIL.n33 0.93369
R183 VTAIL.n134 VTAIL.n102 0.388379
R184 VTAIL.n32 VTAIL.n0 0.388379
R185 VTAIL.n100 VTAIL.n68 0.388379
R186 VTAIL.n66 VTAIL.n34 0.388379
R187 VTAIL VTAIL.n135 0.347483
R188 VTAIL.n114 VTAIL.n109 0.155672
R189 VTAIL.n121 VTAIL.n109 0.155672
R190 VTAIL.n122 VTAIL.n121 0.155672
R191 VTAIL.n122 VTAIL.n105 0.155672
R192 VTAIL.n129 VTAIL.n105 0.155672
R193 VTAIL.n130 VTAIL.n129 0.155672
R194 VTAIL.n12 VTAIL.n7 0.155672
R195 VTAIL.n19 VTAIL.n7 0.155672
R196 VTAIL.n20 VTAIL.n19 0.155672
R197 VTAIL.n20 VTAIL.n3 0.155672
R198 VTAIL.n27 VTAIL.n3 0.155672
R199 VTAIL.n28 VTAIL.n27 0.155672
R200 VTAIL.n96 VTAIL.n95 0.155672
R201 VTAIL.n95 VTAIL.n71 0.155672
R202 VTAIL.n88 VTAIL.n71 0.155672
R203 VTAIL.n88 VTAIL.n87 0.155672
R204 VTAIL.n87 VTAIL.n75 0.155672
R205 VTAIL.n80 VTAIL.n75 0.155672
R206 VTAIL.n62 VTAIL.n61 0.155672
R207 VTAIL.n61 VTAIL.n37 0.155672
R208 VTAIL.n54 VTAIL.n37 0.155672
R209 VTAIL.n54 VTAIL.n53 0.155672
R210 VTAIL.n53 VTAIL.n41 0.155672
R211 VTAIL.n46 VTAIL.n41 0.155672
R212 VDD1.n32 VDD1.n31 289.615
R213 VDD1.n65 VDD1.n64 289.615
R214 VDD1.n31 VDD1.n30 185
R215 VDD1.n2 VDD1.n1 185
R216 VDD1.n25 VDD1.n24 185
R217 VDD1.n23 VDD1.n22 185
R218 VDD1.n6 VDD1.n5 185
R219 VDD1.n17 VDD1.n16 185
R220 VDD1.n15 VDD1.n14 185
R221 VDD1.n10 VDD1.n9 185
R222 VDD1.n43 VDD1.n42 185
R223 VDD1.n48 VDD1.n47 185
R224 VDD1.n50 VDD1.n49 185
R225 VDD1.n39 VDD1.n38 185
R226 VDD1.n56 VDD1.n55 185
R227 VDD1.n58 VDD1.n57 185
R228 VDD1.n35 VDD1.n34 185
R229 VDD1.n64 VDD1.n63 185
R230 VDD1.n11 VDD1.t0 149.525
R231 VDD1.n44 VDD1.t1 149.525
R232 VDD1.n31 VDD1.n1 104.615
R233 VDD1.n24 VDD1.n1 104.615
R234 VDD1.n24 VDD1.n23 104.615
R235 VDD1.n23 VDD1.n5 104.615
R236 VDD1.n16 VDD1.n5 104.615
R237 VDD1.n16 VDD1.n15 104.615
R238 VDD1.n15 VDD1.n9 104.615
R239 VDD1.n48 VDD1.n42 104.615
R240 VDD1.n49 VDD1.n48 104.615
R241 VDD1.n49 VDD1.n38 104.615
R242 VDD1.n56 VDD1.n38 104.615
R243 VDD1.n57 VDD1.n56 104.615
R244 VDD1.n57 VDD1.n34 104.615
R245 VDD1.n64 VDD1.n34 104.615
R246 VDD1 VDD1.n65 83.8154
R247 VDD1.t0 VDD1.n9 52.3082
R248 VDD1.t1 VDD1.n42 52.3082
R249 VDD1 VDD1.n32 50.879
R250 VDD1.n30 VDD1.n0 12.8005
R251 VDD1.n63 VDD1.n33 12.8005
R252 VDD1.n29 VDD1.n2 12.0247
R253 VDD1.n62 VDD1.n35 12.0247
R254 VDD1.n26 VDD1.n25 11.249
R255 VDD1.n59 VDD1.n58 11.249
R256 VDD1.n22 VDD1.n4 10.4732
R257 VDD1.n55 VDD1.n37 10.4732
R258 VDD1.n11 VDD1.n10 10.2746
R259 VDD1.n44 VDD1.n43 10.2746
R260 VDD1.n21 VDD1.n6 9.69747
R261 VDD1.n54 VDD1.n39 9.69747
R262 VDD1.n28 VDD1.n0 9.45567
R263 VDD1.n61 VDD1.n33 9.45567
R264 VDD1.n29 VDD1.n28 9.3005
R265 VDD1.n27 VDD1.n26 9.3005
R266 VDD1.n4 VDD1.n3 9.3005
R267 VDD1.n21 VDD1.n20 9.3005
R268 VDD1.n19 VDD1.n18 9.3005
R269 VDD1.n8 VDD1.n7 9.3005
R270 VDD1.n13 VDD1.n12 9.3005
R271 VDD1.n46 VDD1.n45 9.3005
R272 VDD1.n41 VDD1.n40 9.3005
R273 VDD1.n52 VDD1.n51 9.3005
R274 VDD1.n54 VDD1.n53 9.3005
R275 VDD1.n37 VDD1.n36 9.3005
R276 VDD1.n60 VDD1.n59 9.3005
R277 VDD1.n62 VDD1.n61 9.3005
R278 VDD1.n18 VDD1.n17 8.92171
R279 VDD1.n51 VDD1.n50 8.92171
R280 VDD1.n14 VDD1.n8 8.14595
R281 VDD1.n47 VDD1.n41 8.14595
R282 VDD1.n13 VDD1.n10 7.3702
R283 VDD1.n46 VDD1.n43 7.3702
R284 VDD1.n14 VDD1.n13 5.81868
R285 VDD1.n47 VDD1.n46 5.81868
R286 VDD1.n17 VDD1.n8 5.04292
R287 VDD1.n50 VDD1.n41 5.04292
R288 VDD1.n18 VDD1.n6 4.26717
R289 VDD1.n51 VDD1.n39 4.26717
R290 VDD1.n22 VDD1.n21 3.49141
R291 VDD1.n55 VDD1.n54 3.49141
R292 VDD1.n12 VDD1.n11 2.84308
R293 VDD1.n45 VDD1.n44 2.84308
R294 VDD1.n25 VDD1.n4 2.71565
R295 VDD1.n58 VDD1.n37 2.71565
R296 VDD1.n26 VDD1.n2 1.93989
R297 VDD1.n59 VDD1.n35 1.93989
R298 VDD1.n30 VDD1.n29 1.16414
R299 VDD1.n63 VDD1.n62 1.16414
R300 VDD1.n32 VDD1.n0 0.388379
R301 VDD1.n65 VDD1.n33 0.388379
R302 VDD1.n28 VDD1.n27 0.155672
R303 VDD1.n27 VDD1.n3 0.155672
R304 VDD1.n20 VDD1.n3 0.155672
R305 VDD1.n20 VDD1.n19 0.155672
R306 VDD1.n19 VDD1.n7 0.155672
R307 VDD1.n12 VDD1.n7 0.155672
R308 VDD1.n45 VDD1.n40 0.155672
R309 VDD1.n52 VDD1.n40 0.155672
R310 VDD1.n53 VDD1.n52 0.155672
R311 VDD1.n53 VDD1.n36 0.155672
R312 VDD1.n60 VDD1.n36 0.155672
R313 VDD1.n61 VDD1.n60 0.155672
R314 B.n462 B.n461 585
R315 B.n188 B.n68 585
R316 B.n187 B.n186 585
R317 B.n185 B.n184 585
R318 B.n183 B.n182 585
R319 B.n181 B.n180 585
R320 B.n179 B.n178 585
R321 B.n177 B.n176 585
R322 B.n175 B.n174 585
R323 B.n173 B.n172 585
R324 B.n171 B.n170 585
R325 B.n169 B.n168 585
R326 B.n167 B.n166 585
R327 B.n165 B.n164 585
R328 B.n163 B.n162 585
R329 B.n161 B.n160 585
R330 B.n159 B.n158 585
R331 B.n157 B.n156 585
R332 B.n155 B.n154 585
R333 B.n153 B.n152 585
R334 B.n151 B.n150 585
R335 B.n149 B.n148 585
R336 B.n147 B.n146 585
R337 B.n145 B.n144 585
R338 B.n143 B.n142 585
R339 B.n140 B.n139 585
R340 B.n138 B.n137 585
R341 B.n136 B.n135 585
R342 B.n134 B.n133 585
R343 B.n132 B.n131 585
R344 B.n130 B.n129 585
R345 B.n128 B.n127 585
R346 B.n126 B.n125 585
R347 B.n124 B.n123 585
R348 B.n122 B.n121 585
R349 B.n119 B.n118 585
R350 B.n117 B.n116 585
R351 B.n115 B.n114 585
R352 B.n113 B.n112 585
R353 B.n111 B.n110 585
R354 B.n109 B.n108 585
R355 B.n107 B.n106 585
R356 B.n105 B.n104 585
R357 B.n103 B.n102 585
R358 B.n101 B.n100 585
R359 B.n99 B.n98 585
R360 B.n97 B.n96 585
R361 B.n95 B.n94 585
R362 B.n93 B.n92 585
R363 B.n91 B.n90 585
R364 B.n89 B.n88 585
R365 B.n87 B.n86 585
R366 B.n85 B.n84 585
R367 B.n83 B.n82 585
R368 B.n81 B.n80 585
R369 B.n79 B.n78 585
R370 B.n77 B.n76 585
R371 B.n75 B.n74 585
R372 B.n39 B.n38 585
R373 B.n467 B.n466 585
R374 B.n460 B.n69 585
R375 B.n69 B.n36 585
R376 B.n459 B.n35 585
R377 B.n471 B.n35 585
R378 B.n458 B.n34 585
R379 B.n472 B.n34 585
R380 B.n457 B.n33 585
R381 B.n473 B.n33 585
R382 B.n456 B.n455 585
R383 B.n455 B.n29 585
R384 B.n454 B.n28 585
R385 B.n479 B.n28 585
R386 B.n453 B.n27 585
R387 B.n480 B.n27 585
R388 B.n452 B.n26 585
R389 B.n481 B.n26 585
R390 B.n451 B.n450 585
R391 B.n450 B.n22 585
R392 B.n449 B.n21 585
R393 B.n487 B.n21 585
R394 B.n448 B.n20 585
R395 B.n488 B.n20 585
R396 B.n447 B.n19 585
R397 B.n489 B.n19 585
R398 B.n446 B.n445 585
R399 B.n445 B.n15 585
R400 B.n444 B.n14 585
R401 B.n495 B.n14 585
R402 B.n443 B.n13 585
R403 B.n496 B.n13 585
R404 B.n442 B.n12 585
R405 B.n497 B.n12 585
R406 B.n441 B.n440 585
R407 B.n440 B.n8 585
R408 B.n439 B.n7 585
R409 B.n503 B.n7 585
R410 B.n438 B.n6 585
R411 B.n504 B.n6 585
R412 B.n437 B.n5 585
R413 B.n505 B.n5 585
R414 B.n436 B.n435 585
R415 B.n435 B.n4 585
R416 B.n434 B.n189 585
R417 B.n434 B.n433 585
R418 B.n424 B.n190 585
R419 B.n191 B.n190 585
R420 B.n426 B.n425 585
R421 B.n427 B.n426 585
R422 B.n423 B.n195 585
R423 B.n199 B.n195 585
R424 B.n422 B.n421 585
R425 B.n421 B.n420 585
R426 B.n197 B.n196 585
R427 B.n198 B.n197 585
R428 B.n413 B.n412 585
R429 B.n414 B.n413 585
R430 B.n411 B.n204 585
R431 B.n204 B.n203 585
R432 B.n410 B.n409 585
R433 B.n409 B.n408 585
R434 B.n206 B.n205 585
R435 B.n207 B.n206 585
R436 B.n401 B.n400 585
R437 B.n402 B.n401 585
R438 B.n399 B.n212 585
R439 B.n212 B.n211 585
R440 B.n398 B.n397 585
R441 B.n397 B.n396 585
R442 B.n214 B.n213 585
R443 B.n215 B.n214 585
R444 B.n389 B.n388 585
R445 B.n390 B.n389 585
R446 B.n387 B.n220 585
R447 B.n220 B.n219 585
R448 B.n386 B.n385 585
R449 B.n385 B.n384 585
R450 B.n222 B.n221 585
R451 B.n223 B.n222 585
R452 B.n380 B.n379 585
R453 B.n226 B.n225 585
R454 B.n376 B.n375 585
R455 B.n377 B.n376 585
R456 B.n374 B.n256 585
R457 B.n373 B.n372 585
R458 B.n371 B.n370 585
R459 B.n369 B.n368 585
R460 B.n367 B.n366 585
R461 B.n365 B.n364 585
R462 B.n363 B.n362 585
R463 B.n361 B.n360 585
R464 B.n359 B.n358 585
R465 B.n357 B.n356 585
R466 B.n355 B.n354 585
R467 B.n353 B.n352 585
R468 B.n351 B.n350 585
R469 B.n349 B.n348 585
R470 B.n347 B.n346 585
R471 B.n345 B.n344 585
R472 B.n343 B.n342 585
R473 B.n341 B.n340 585
R474 B.n339 B.n338 585
R475 B.n337 B.n336 585
R476 B.n335 B.n334 585
R477 B.n333 B.n332 585
R478 B.n331 B.n330 585
R479 B.n329 B.n328 585
R480 B.n327 B.n326 585
R481 B.n325 B.n324 585
R482 B.n323 B.n322 585
R483 B.n321 B.n320 585
R484 B.n319 B.n318 585
R485 B.n317 B.n316 585
R486 B.n315 B.n314 585
R487 B.n313 B.n312 585
R488 B.n311 B.n310 585
R489 B.n309 B.n308 585
R490 B.n307 B.n306 585
R491 B.n305 B.n304 585
R492 B.n303 B.n302 585
R493 B.n301 B.n300 585
R494 B.n299 B.n298 585
R495 B.n297 B.n296 585
R496 B.n295 B.n294 585
R497 B.n293 B.n292 585
R498 B.n291 B.n290 585
R499 B.n289 B.n288 585
R500 B.n287 B.n286 585
R501 B.n285 B.n284 585
R502 B.n283 B.n282 585
R503 B.n281 B.n280 585
R504 B.n279 B.n278 585
R505 B.n277 B.n276 585
R506 B.n275 B.n274 585
R507 B.n273 B.n272 585
R508 B.n271 B.n270 585
R509 B.n269 B.n268 585
R510 B.n267 B.n266 585
R511 B.n265 B.n264 585
R512 B.n263 B.n255 585
R513 B.n377 B.n255 585
R514 B.n381 B.n224 585
R515 B.n224 B.n223 585
R516 B.n383 B.n382 585
R517 B.n384 B.n383 585
R518 B.n218 B.n217 585
R519 B.n219 B.n218 585
R520 B.n392 B.n391 585
R521 B.n391 B.n390 585
R522 B.n393 B.n216 585
R523 B.n216 B.n215 585
R524 B.n395 B.n394 585
R525 B.n396 B.n395 585
R526 B.n210 B.n209 585
R527 B.n211 B.n210 585
R528 B.n404 B.n403 585
R529 B.n403 B.n402 585
R530 B.n405 B.n208 585
R531 B.n208 B.n207 585
R532 B.n407 B.n406 585
R533 B.n408 B.n407 585
R534 B.n202 B.n201 585
R535 B.n203 B.n202 585
R536 B.n416 B.n415 585
R537 B.n415 B.n414 585
R538 B.n417 B.n200 585
R539 B.n200 B.n198 585
R540 B.n419 B.n418 585
R541 B.n420 B.n419 585
R542 B.n194 B.n193 585
R543 B.n199 B.n194 585
R544 B.n429 B.n428 585
R545 B.n428 B.n427 585
R546 B.n430 B.n192 585
R547 B.n192 B.n191 585
R548 B.n432 B.n431 585
R549 B.n433 B.n432 585
R550 B.n2 B.n0 585
R551 B.n4 B.n2 585
R552 B.n3 B.n1 585
R553 B.n504 B.n3 585
R554 B.n502 B.n501 585
R555 B.n503 B.n502 585
R556 B.n500 B.n9 585
R557 B.n9 B.n8 585
R558 B.n499 B.n498 585
R559 B.n498 B.n497 585
R560 B.n11 B.n10 585
R561 B.n496 B.n11 585
R562 B.n494 B.n493 585
R563 B.n495 B.n494 585
R564 B.n492 B.n16 585
R565 B.n16 B.n15 585
R566 B.n491 B.n490 585
R567 B.n490 B.n489 585
R568 B.n18 B.n17 585
R569 B.n488 B.n18 585
R570 B.n486 B.n485 585
R571 B.n487 B.n486 585
R572 B.n484 B.n23 585
R573 B.n23 B.n22 585
R574 B.n483 B.n482 585
R575 B.n482 B.n481 585
R576 B.n25 B.n24 585
R577 B.n480 B.n25 585
R578 B.n478 B.n477 585
R579 B.n479 B.n478 585
R580 B.n476 B.n30 585
R581 B.n30 B.n29 585
R582 B.n475 B.n474 585
R583 B.n474 B.n473 585
R584 B.n32 B.n31 585
R585 B.n472 B.n32 585
R586 B.n470 B.n469 585
R587 B.n471 B.n470 585
R588 B.n468 B.n37 585
R589 B.n37 B.n36 585
R590 B.n507 B.n506 585
R591 B.n506 B.n505 585
R592 B.n379 B.n224 545.355
R593 B.n466 B.n37 545.355
R594 B.n255 B.n222 545.355
R595 B.n462 B.n69 545.355
R596 B.n260 B.t6 306.065
R597 B.n257 B.t2 306.065
R598 B.n72 B.t13 306.065
R599 B.n70 B.t9 306.065
R600 B.n464 B.n463 256.663
R601 B.n464 B.n67 256.663
R602 B.n464 B.n66 256.663
R603 B.n464 B.n65 256.663
R604 B.n464 B.n64 256.663
R605 B.n464 B.n63 256.663
R606 B.n464 B.n62 256.663
R607 B.n464 B.n61 256.663
R608 B.n464 B.n60 256.663
R609 B.n464 B.n59 256.663
R610 B.n464 B.n58 256.663
R611 B.n464 B.n57 256.663
R612 B.n464 B.n56 256.663
R613 B.n464 B.n55 256.663
R614 B.n464 B.n54 256.663
R615 B.n464 B.n53 256.663
R616 B.n464 B.n52 256.663
R617 B.n464 B.n51 256.663
R618 B.n464 B.n50 256.663
R619 B.n464 B.n49 256.663
R620 B.n464 B.n48 256.663
R621 B.n464 B.n47 256.663
R622 B.n464 B.n46 256.663
R623 B.n464 B.n45 256.663
R624 B.n464 B.n44 256.663
R625 B.n464 B.n43 256.663
R626 B.n464 B.n42 256.663
R627 B.n464 B.n41 256.663
R628 B.n464 B.n40 256.663
R629 B.n465 B.n464 256.663
R630 B.n378 B.n377 256.663
R631 B.n377 B.n227 256.663
R632 B.n377 B.n228 256.663
R633 B.n377 B.n229 256.663
R634 B.n377 B.n230 256.663
R635 B.n377 B.n231 256.663
R636 B.n377 B.n232 256.663
R637 B.n377 B.n233 256.663
R638 B.n377 B.n234 256.663
R639 B.n377 B.n235 256.663
R640 B.n377 B.n236 256.663
R641 B.n377 B.n237 256.663
R642 B.n377 B.n238 256.663
R643 B.n377 B.n239 256.663
R644 B.n377 B.n240 256.663
R645 B.n377 B.n241 256.663
R646 B.n377 B.n242 256.663
R647 B.n377 B.n243 256.663
R648 B.n377 B.n244 256.663
R649 B.n377 B.n245 256.663
R650 B.n377 B.n246 256.663
R651 B.n377 B.n247 256.663
R652 B.n377 B.n248 256.663
R653 B.n377 B.n249 256.663
R654 B.n377 B.n250 256.663
R655 B.n377 B.n251 256.663
R656 B.n377 B.n252 256.663
R657 B.n377 B.n253 256.663
R658 B.n377 B.n254 256.663
R659 B.n260 B.t8 222.858
R660 B.n70 B.t11 222.858
R661 B.n257 B.t5 222.858
R662 B.n72 B.t14 222.858
R663 B.n261 B.t7 186.399
R664 B.n71 B.t12 186.399
R665 B.n258 B.t4 186.399
R666 B.n73 B.t15 186.399
R667 B.n383 B.n224 163.367
R668 B.n383 B.n218 163.367
R669 B.n391 B.n218 163.367
R670 B.n391 B.n216 163.367
R671 B.n395 B.n216 163.367
R672 B.n395 B.n210 163.367
R673 B.n403 B.n210 163.367
R674 B.n403 B.n208 163.367
R675 B.n407 B.n208 163.367
R676 B.n407 B.n202 163.367
R677 B.n415 B.n202 163.367
R678 B.n415 B.n200 163.367
R679 B.n419 B.n200 163.367
R680 B.n419 B.n194 163.367
R681 B.n428 B.n194 163.367
R682 B.n428 B.n192 163.367
R683 B.n432 B.n192 163.367
R684 B.n432 B.n2 163.367
R685 B.n506 B.n2 163.367
R686 B.n506 B.n3 163.367
R687 B.n502 B.n3 163.367
R688 B.n502 B.n9 163.367
R689 B.n498 B.n9 163.367
R690 B.n498 B.n11 163.367
R691 B.n494 B.n11 163.367
R692 B.n494 B.n16 163.367
R693 B.n490 B.n16 163.367
R694 B.n490 B.n18 163.367
R695 B.n486 B.n18 163.367
R696 B.n486 B.n23 163.367
R697 B.n482 B.n23 163.367
R698 B.n482 B.n25 163.367
R699 B.n478 B.n25 163.367
R700 B.n478 B.n30 163.367
R701 B.n474 B.n30 163.367
R702 B.n474 B.n32 163.367
R703 B.n470 B.n32 163.367
R704 B.n470 B.n37 163.367
R705 B.n376 B.n226 163.367
R706 B.n376 B.n256 163.367
R707 B.n372 B.n371 163.367
R708 B.n368 B.n367 163.367
R709 B.n364 B.n363 163.367
R710 B.n360 B.n359 163.367
R711 B.n356 B.n355 163.367
R712 B.n352 B.n351 163.367
R713 B.n348 B.n347 163.367
R714 B.n344 B.n343 163.367
R715 B.n340 B.n339 163.367
R716 B.n336 B.n335 163.367
R717 B.n332 B.n331 163.367
R718 B.n328 B.n327 163.367
R719 B.n324 B.n323 163.367
R720 B.n320 B.n319 163.367
R721 B.n316 B.n315 163.367
R722 B.n312 B.n311 163.367
R723 B.n308 B.n307 163.367
R724 B.n304 B.n303 163.367
R725 B.n300 B.n299 163.367
R726 B.n296 B.n295 163.367
R727 B.n292 B.n291 163.367
R728 B.n288 B.n287 163.367
R729 B.n284 B.n283 163.367
R730 B.n280 B.n279 163.367
R731 B.n276 B.n275 163.367
R732 B.n272 B.n271 163.367
R733 B.n268 B.n267 163.367
R734 B.n264 B.n255 163.367
R735 B.n385 B.n222 163.367
R736 B.n385 B.n220 163.367
R737 B.n389 B.n220 163.367
R738 B.n389 B.n214 163.367
R739 B.n397 B.n214 163.367
R740 B.n397 B.n212 163.367
R741 B.n401 B.n212 163.367
R742 B.n401 B.n206 163.367
R743 B.n409 B.n206 163.367
R744 B.n409 B.n204 163.367
R745 B.n413 B.n204 163.367
R746 B.n413 B.n197 163.367
R747 B.n421 B.n197 163.367
R748 B.n421 B.n195 163.367
R749 B.n426 B.n195 163.367
R750 B.n426 B.n190 163.367
R751 B.n434 B.n190 163.367
R752 B.n435 B.n434 163.367
R753 B.n435 B.n5 163.367
R754 B.n6 B.n5 163.367
R755 B.n7 B.n6 163.367
R756 B.n440 B.n7 163.367
R757 B.n440 B.n12 163.367
R758 B.n13 B.n12 163.367
R759 B.n14 B.n13 163.367
R760 B.n445 B.n14 163.367
R761 B.n445 B.n19 163.367
R762 B.n20 B.n19 163.367
R763 B.n21 B.n20 163.367
R764 B.n450 B.n21 163.367
R765 B.n450 B.n26 163.367
R766 B.n27 B.n26 163.367
R767 B.n28 B.n27 163.367
R768 B.n455 B.n28 163.367
R769 B.n455 B.n33 163.367
R770 B.n34 B.n33 163.367
R771 B.n35 B.n34 163.367
R772 B.n69 B.n35 163.367
R773 B.n74 B.n39 163.367
R774 B.n78 B.n77 163.367
R775 B.n82 B.n81 163.367
R776 B.n86 B.n85 163.367
R777 B.n90 B.n89 163.367
R778 B.n94 B.n93 163.367
R779 B.n98 B.n97 163.367
R780 B.n102 B.n101 163.367
R781 B.n106 B.n105 163.367
R782 B.n110 B.n109 163.367
R783 B.n114 B.n113 163.367
R784 B.n118 B.n117 163.367
R785 B.n123 B.n122 163.367
R786 B.n127 B.n126 163.367
R787 B.n131 B.n130 163.367
R788 B.n135 B.n134 163.367
R789 B.n139 B.n138 163.367
R790 B.n144 B.n143 163.367
R791 B.n148 B.n147 163.367
R792 B.n152 B.n151 163.367
R793 B.n156 B.n155 163.367
R794 B.n160 B.n159 163.367
R795 B.n164 B.n163 163.367
R796 B.n168 B.n167 163.367
R797 B.n172 B.n171 163.367
R798 B.n176 B.n175 163.367
R799 B.n180 B.n179 163.367
R800 B.n184 B.n183 163.367
R801 B.n186 B.n68 163.367
R802 B.n377 B.n223 126.546
R803 B.n464 B.n36 126.546
R804 B.n379 B.n378 71.676
R805 B.n256 B.n227 71.676
R806 B.n371 B.n228 71.676
R807 B.n367 B.n229 71.676
R808 B.n363 B.n230 71.676
R809 B.n359 B.n231 71.676
R810 B.n355 B.n232 71.676
R811 B.n351 B.n233 71.676
R812 B.n347 B.n234 71.676
R813 B.n343 B.n235 71.676
R814 B.n339 B.n236 71.676
R815 B.n335 B.n237 71.676
R816 B.n331 B.n238 71.676
R817 B.n327 B.n239 71.676
R818 B.n323 B.n240 71.676
R819 B.n319 B.n241 71.676
R820 B.n315 B.n242 71.676
R821 B.n311 B.n243 71.676
R822 B.n307 B.n244 71.676
R823 B.n303 B.n245 71.676
R824 B.n299 B.n246 71.676
R825 B.n295 B.n247 71.676
R826 B.n291 B.n248 71.676
R827 B.n287 B.n249 71.676
R828 B.n283 B.n250 71.676
R829 B.n279 B.n251 71.676
R830 B.n275 B.n252 71.676
R831 B.n271 B.n253 71.676
R832 B.n267 B.n254 71.676
R833 B.n466 B.n465 71.676
R834 B.n74 B.n40 71.676
R835 B.n78 B.n41 71.676
R836 B.n82 B.n42 71.676
R837 B.n86 B.n43 71.676
R838 B.n90 B.n44 71.676
R839 B.n94 B.n45 71.676
R840 B.n98 B.n46 71.676
R841 B.n102 B.n47 71.676
R842 B.n106 B.n48 71.676
R843 B.n110 B.n49 71.676
R844 B.n114 B.n50 71.676
R845 B.n118 B.n51 71.676
R846 B.n123 B.n52 71.676
R847 B.n127 B.n53 71.676
R848 B.n131 B.n54 71.676
R849 B.n135 B.n55 71.676
R850 B.n139 B.n56 71.676
R851 B.n144 B.n57 71.676
R852 B.n148 B.n58 71.676
R853 B.n152 B.n59 71.676
R854 B.n156 B.n60 71.676
R855 B.n160 B.n61 71.676
R856 B.n164 B.n62 71.676
R857 B.n168 B.n63 71.676
R858 B.n172 B.n64 71.676
R859 B.n176 B.n65 71.676
R860 B.n180 B.n66 71.676
R861 B.n184 B.n67 71.676
R862 B.n463 B.n68 71.676
R863 B.n463 B.n462 71.676
R864 B.n186 B.n67 71.676
R865 B.n183 B.n66 71.676
R866 B.n179 B.n65 71.676
R867 B.n175 B.n64 71.676
R868 B.n171 B.n63 71.676
R869 B.n167 B.n62 71.676
R870 B.n163 B.n61 71.676
R871 B.n159 B.n60 71.676
R872 B.n155 B.n59 71.676
R873 B.n151 B.n58 71.676
R874 B.n147 B.n57 71.676
R875 B.n143 B.n56 71.676
R876 B.n138 B.n55 71.676
R877 B.n134 B.n54 71.676
R878 B.n130 B.n53 71.676
R879 B.n126 B.n52 71.676
R880 B.n122 B.n51 71.676
R881 B.n117 B.n50 71.676
R882 B.n113 B.n49 71.676
R883 B.n109 B.n48 71.676
R884 B.n105 B.n47 71.676
R885 B.n101 B.n46 71.676
R886 B.n97 B.n45 71.676
R887 B.n93 B.n44 71.676
R888 B.n89 B.n43 71.676
R889 B.n85 B.n42 71.676
R890 B.n81 B.n41 71.676
R891 B.n77 B.n40 71.676
R892 B.n465 B.n39 71.676
R893 B.n378 B.n226 71.676
R894 B.n372 B.n227 71.676
R895 B.n368 B.n228 71.676
R896 B.n364 B.n229 71.676
R897 B.n360 B.n230 71.676
R898 B.n356 B.n231 71.676
R899 B.n352 B.n232 71.676
R900 B.n348 B.n233 71.676
R901 B.n344 B.n234 71.676
R902 B.n340 B.n235 71.676
R903 B.n336 B.n236 71.676
R904 B.n332 B.n237 71.676
R905 B.n328 B.n238 71.676
R906 B.n324 B.n239 71.676
R907 B.n320 B.n240 71.676
R908 B.n316 B.n241 71.676
R909 B.n312 B.n242 71.676
R910 B.n308 B.n243 71.676
R911 B.n304 B.n244 71.676
R912 B.n300 B.n245 71.676
R913 B.n296 B.n246 71.676
R914 B.n292 B.n247 71.676
R915 B.n288 B.n248 71.676
R916 B.n284 B.n249 71.676
R917 B.n280 B.n250 71.676
R918 B.n276 B.n251 71.676
R919 B.n272 B.n252 71.676
R920 B.n268 B.n253 71.676
R921 B.n264 B.n254 71.676
R922 B.n384 B.n223 63.7414
R923 B.n384 B.n219 63.7414
R924 B.n390 B.n219 63.7414
R925 B.n390 B.n215 63.7414
R926 B.n396 B.n215 63.7414
R927 B.n402 B.n211 63.7414
R928 B.n402 B.n207 63.7414
R929 B.n408 B.n207 63.7414
R930 B.n408 B.n203 63.7414
R931 B.n414 B.n203 63.7414
R932 B.n414 B.n198 63.7414
R933 B.n420 B.n198 63.7414
R934 B.n420 B.n199 63.7414
R935 B.n427 B.n191 63.7414
R936 B.n433 B.n191 63.7414
R937 B.n433 B.n4 63.7414
R938 B.n505 B.n4 63.7414
R939 B.n505 B.n504 63.7414
R940 B.n504 B.n503 63.7414
R941 B.n503 B.n8 63.7414
R942 B.n497 B.n8 63.7414
R943 B.n496 B.n495 63.7414
R944 B.n495 B.n15 63.7414
R945 B.n489 B.n15 63.7414
R946 B.n489 B.n488 63.7414
R947 B.n488 B.n487 63.7414
R948 B.n487 B.n22 63.7414
R949 B.n481 B.n22 63.7414
R950 B.n481 B.n480 63.7414
R951 B.n479 B.n29 63.7414
R952 B.n473 B.n29 63.7414
R953 B.n473 B.n472 63.7414
R954 B.n472 B.n471 63.7414
R955 B.n471 B.n36 63.7414
R956 B.n262 B.n261 59.5399
R957 B.n259 B.n258 59.5399
R958 B.n120 B.n73 59.5399
R959 B.n141 B.n71 59.5399
R960 B.n396 B.t3 57.1799
R961 B.t10 B.n479 57.1799
R962 B.n199 B.t0 40.3073
R963 B.t1 B.n496 40.3073
R964 B.n261 B.n260 36.4611
R965 B.n258 B.n257 36.4611
R966 B.n73 B.n72 36.4611
R967 B.n71 B.n70 36.4611
R968 B.n461 B.n460 35.4346
R969 B.n468 B.n467 35.4346
R970 B.n263 B.n221 35.4346
R971 B.n381 B.n380 35.4346
R972 B.n427 B.t0 23.4347
R973 B.n497 B.t1 23.4347
R974 B B.n507 18.0485
R975 B.n467 B.n38 10.6151
R976 B.n75 B.n38 10.6151
R977 B.n76 B.n75 10.6151
R978 B.n79 B.n76 10.6151
R979 B.n80 B.n79 10.6151
R980 B.n83 B.n80 10.6151
R981 B.n84 B.n83 10.6151
R982 B.n87 B.n84 10.6151
R983 B.n88 B.n87 10.6151
R984 B.n91 B.n88 10.6151
R985 B.n92 B.n91 10.6151
R986 B.n95 B.n92 10.6151
R987 B.n96 B.n95 10.6151
R988 B.n99 B.n96 10.6151
R989 B.n100 B.n99 10.6151
R990 B.n103 B.n100 10.6151
R991 B.n104 B.n103 10.6151
R992 B.n107 B.n104 10.6151
R993 B.n108 B.n107 10.6151
R994 B.n111 B.n108 10.6151
R995 B.n112 B.n111 10.6151
R996 B.n115 B.n112 10.6151
R997 B.n116 B.n115 10.6151
R998 B.n119 B.n116 10.6151
R999 B.n124 B.n121 10.6151
R1000 B.n125 B.n124 10.6151
R1001 B.n128 B.n125 10.6151
R1002 B.n129 B.n128 10.6151
R1003 B.n132 B.n129 10.6151
R1004 B.n133 B.n132 10.6151
R1005 B.n136 B.n133 10.6151
R1006 B.n137 B.n136 10.6151
R1007 B.n140 B.n137 10.6151
R1008 B.n145 B.n142 10.6151
R1009 B.n146 B.n145 10.6151
R1010 B.n149 B.n146 10.6151
R1011 B.n150 B.n149 10.6151
R1012 B.n153 B.n150 10.6151
R1013 B.n154 B.n153 10.6151
R1014 B.n157 B.n154 10.6151
R1015 B.n158 B.n157 10.6151
R1016 B.n161 B.n158 10.6151
R1017 B.n162 B.n161 10.6151
R1018 B.n165 B.n162 10.6151
R1019 B.n166 B.n165 10.6151
R1020 B.n169 B.n166 10.6151
R1021 B.n170 B.n169 10.6151
R1022 B.n173 B.n170 10.6151
R1023 B.n174 B.n173 10.6151
R1024 B.n177 B.n174 10.6151
R1025 B.n178 B.n177 10.6151
R1026 B.n181 B.n178 10.6151
R1027 B.n182 B.n181 10.6151
R1028 B.n185 B.n182 10.6151
R1029 B.n187 B.n185 10.6151
R1030 B.n188 B.n187 10.6151
R1031 B.n461 B.n188 10.6151
R1032 B.n386 B.n221 10.6151
R1033 B.n387 B.n386 10.6151
R1034 B.n388 B.n387 10.6151
R1035 B.n388 B.n213 10.6151
R1036 B.n398 B.n213 10.6151
R1037 B.n399 B.n398 10.6151
R1038 B.n400 B.n399 10.6151
R1039 B.n400 B.n205 10.6151
R1040 B.n410 B.n205 10.6151
R1041 B.n411 B.n410 10.6151
R1042 B.n412 B.n411 10.6151
R1043 B.n412 B.n196 10.6151
R1044 B.n422 B.n196 10.6151
R1045 B.n423 B.n422 10.6151
R1046 B.n425 B.n423 10.6151
R1047 B.n425 B.n424 10.6151
R1048 B.n424 B.n189 10.6151
R1049 B.n436 B.n189 10.6151
R1050 B.n437 B.n436 10.6151
R1051 B.n438 B.n437 10.6151
R1052 B.n439 B.n438 10.6151
R1053 B.n441 B.n439 10.6151
R1054 B.n442 B.n441 10.6151
R1055 B.n443 B.n442 10.6151
R1056 B.n444 B.n443 10.6151
R1057 B.n446 B.n444 10.6151
R1058 B.n447 B.n446 10.6151
R1059 B.n448 B.n447 10.6151
R1060 B.n449 B.n448 10.6151
R1061 B.n451 B.n449 10.6151
R1062 B.n452 B.n451 10.6151
R1063 B.n453 B.n452 10.6151
R1064 B.n454 B.n453 10.6151
R1065 B.n456 B.n454 10.6151
R1066 B.n457 B.n456 10.6151
R1067 B.n458 B.n457 10.6151
R1068 B.n459 B.n458 10.6151
R1069 B.n460 B.n459 10.6151
R1070 B.n380 B.n225 10.6151
R1071 B.n375 B.n225 10.6151
R1072 B.n375 B.n374 10.6151
R1073 B.n374 B.n373 10.6151
R1074 B.n373 B.n370 10.6151
R1075 B.n370 B.n369 10.6151
R1076 B.n369 B.n366 10.6151
R1077 B.n366 B.n365 10.6151
R1078 B.n365 B.n362 10.6151
R1079 B.n362 B.n361 10.6151
R1080 B.n361 B.n358 10.6151
R1081 B.n358 B.n357 10.6151
R1082 B.n357 B.n354 10.6151
R1083 B.n354 B.n353 10.6151
R1084 B.n353 B.n350 10.6151
R1085 B.n350 B.n349 10.6151
R1086 B.n349 B.n346 10.6151
R1087 B.n346 B.n345 10.6151
R1088 B.n345 B.n342 10.6151
R1089 B.n342 B.n341 10.6151
R1090 B.n341 B.n338 10.6151
R1091 B.n338 B.n337 10.6151
R1092 B.n337 B.n334 10.6151
R1093 B.n334 B.n333 10.6151
R1094 B.n330 B.n329 10.6151
R1095 B.n329 B.n326 10.6151
R1096 B.n326 B.n325 10.6151
R1097 B.n325 B.n322 10.6151
R1098 B.n322 B.n321 10.6151
R1099 B.n321 B.n318 10.6151
R1100 B.n318 B.n317 10.6151
R1101 B.n317 B.n314 10.6151
R1102 B.n314 B.n313 10.6151
R1103 B.n310 B.n309 10.6151
R1104 B.n309 B.n306 10.6151
R1105 B.n306 B.n305 10.6151
R1106 B.n305 B.n302 10.6151
R1107 B.n302 B.n301 10.6151
R1108 B.n301 B.n298 10.6151
R1109 B.n298 B.n297 10.6151
R1110 B.n297 B.n294 10.6151
R1111 B.n294 B.n293 10.6151
R1112 B.n293 B.n290 10.6151
R1113 B.n290 B.n289 10.6151
R1114 B.n289 B.n286 10.6151
R1115 B.n286 B.n285 10.6151
R1116 B.n285 B.n282 10.6151
R1117 B.n282 B.n281 10.6151
R1118 B.n281 B.n278 10.6151
R1119 B.n278 B.n277 10.6151
R1120 B.n277 B.n274 10.6151
R1121 B.n274 B.n273 10.6151
R1122 B.n273 B.n270 10.6151
R1123 B.n270 B.n269 10.6151
R1124 B.n269 B.n266 10.6151
R1125 B.n266 B.n265 10.6151
R1126 B.n265 B.n263 10.6151
R1127 B.n382 B.n381 10.6151
R1128 B.n382 B.n217 10.6151
R1129 B.n392 B.n217 10.6151
R1130 B.n393 B.n392 10.6151
R1131 B.n394 B.n393 10.6151
R1132 B.n394 B.n209 10.6151
R1133 B.n404 B.n209 10.6151
R1134 B.n405 B.n404 10.6151
R1135 B.n406 B.n405 10.6151
R1136 B.n406 B.n201 10.6151
R1137 B.n416 B.n201 10.6151
R1138 B.n417 B.n416 10.6151
R1139 B.n418 B.n417 10.6151
R1140 B.n418 B.n193 10.6151
R1141 B.n429 B.n193 10.6151
R1142 B.n430 B.n429 10.6151
R1143 B.n431 B.n430 10.6151
R1144 B.n431 B.n0 10.6151
R1145 B.n501 B.n1 10.6151
R1146 B.n501 B.n500 10.6151
R1147 B.n500 B.n499 10.6151
R1148 B.n499 B.n10 10.6151
R1149 B.n493 B.n10 10.6151
R1150 B.n493 B.n492 10.6151
R1151 B.n492 B.n491 10.6151
R1152 B.n491 B.n17 10.6151
R1153 B.n485 B.n17 10.6151
R1154 B.n485 B.n484 10.6151
R1155 B.n484 B.n483 10.6151
R1156 B.n483 B.n24 10.6151
R1157 B.n477 B.n24 10.6151
R1158 B.n477 B.n476 10.6151
R1159 B.n476 B.n475 10.6151
R1160 B.n475 B.n31 10.6151
R1161 B.n469 B.n31 10.6151
R1162 B.n469 B.n468 10.6151
R1163 B.n120 B.n119 9.36635
R1164 B.n142 B.n141 9.36635
R1165 B.n333 B.n259 9.36635
R1166 B.n310 B.n262 9.36635
R1167 B.t3 B.n211 6.56207
R1168 B.n480 B.t10 6.56207
R1169 B.n507 B.n0 2.81026
R1170 B.n507 B.n1 2.81026
R1171 B.n121 B.n120 1.24928
R1172 B.n141 B.n140 1.24928
R1173 B.n330 B.n259 1.24928
R1174 B.n313 B.n262 1.24928
R1175 VN VN.t0 244.351
R1176 VN VN.t1 206.536
R1177 VDD2.n65 VDD2.n64 289.615
R1178 VDD2.n32 VDD2.n31 289.615
R1179 VDD2.n64 VDD2.n63 185
R1180 VDD2.n35 VDD2.n34 185
R1181 VDD2.n58 VDD2.n57 185
R1182 VDD2.n56 VDD2.n55 185
R1183 VDD2.n39 VDD2.n38 185
R1184 VDD2.n50 VDD2.n49 185
R1185 VDD2.n48 VDD2.n47 185
R1186 VDD2.n43 VDD2.n42 185
R1187 VDD2.n10 VDD2.n9 185
R1188 VDD2.n15 VDD2.n14 185
R1189 VDD2.n17 VDD2.n16 185
R1190 VDD2.n6 VDD2.n5 185
R1191 VDD2.n23 VDD2.n22 185
R1192 VDD2.n25 VDD2.n24 185
R1193 VDD2.n2 VDD2.n1 185
R1194 VDD2.n31 VDD2.n30 185
R1195 VDD2.n44 VDD2.t1 149.525
R1196 VDD2.n11 VDD2.t0 149.525
R1197 VDD2.n64 VDD2.n34 104.615
R1198 VDD2.n57 VDD2.n34 104.615
R1199 VDD2.n57 VDD2.n56 104.615
R1200 VDD2.n56 VDD2.n38 104.615
R1201 VDD2.n49 VDD2.n38 104.615
R1202 VDD2.n49 VDD2.n48 104.615
R1203 VDD2.n48 VDD2.n42 104.615
R1204 VDD2.n15 VDD2.n9 104.615
R1205 VDD2.n16 VDD2.n15 104.615
R1206 VDD2.n16 VDD2.n5 104.615
R1207 VDD2.n23 VDD2.n5 104.615
R1208 VDD2.n24 VDD2.n23 104.615
R1209 VDD2.n24 VDD2.n1 104.615
R1210 VDD2.n31 VDD2.n1 104.615
R1211 VDD2.n66 VDD2.n32 82.8854
R1212 VDD2.t1 VDD2.n42 52.3082
R1213 VDD2.t0 VDD2.n9 52.3082
R1214 VDD2.n66 VDD2.n65 50.4157
R1215 VDD2.n63 VDD2.n33 12.8005
R1216 VDD2.n30 VDD2.n0 12.8005
R1217 VDD2.n62 VDD2.n35 12.0247
R1218 VDD2.n29 VDD2.n2 12.0247
R1219 VDD2.n59 VDD2.n58 11.249
R1220 VDD2.n26 VDD2.n25 11.249
R1221 VDD2.n55 VDD2.n37 10.4732
R1222 VDD2.n22 VDD2.n4 10.4732
R1223 VDD2.n44 VDD2.n43 10.2746
R1224 VDD2.n11 VDD2.n10 10.2746
R1225 VDD2.n54 VDD2.n39 9.69747
R1226 VDD2.n21 VDD2.n6 9.69747
R1227 VDD2.n61 VDD2.n33 9.45567
R1228 VDD2.n28 VDD2.n0 9.45567
R1229 VDD2.n62 VDD2.n61 9.3005
R1230 VDD2.n60 VDD2.n59 9.3005
R1231 VDD2.n37 VDD2.n36 9.3005
R1232 VDD2.n54 VDD2.n53 9.3005
R1233 VDD2.n52 VDD2.n51 9.3005
R1234 VDD2.n41 VDD2.n40 9.3005
R1235 VDD2.n46 VDD2.n45 9.3005
R1236 VDD2.n13 VDD2.n12 9.3005
R1237 VDD2.n8 VDD2.n7 9.3005
R1238 VDD2.n19 VDD2.n18 9.3005
R1239 VDD2.n21 VDD2.n20 9.3005
R1240 VDD2.n4 VDD2.n3 9.3005
R1241 VDD2.n27 VDD2.n26 9.3005
R1242 VDD2.n29 VDD2.n28 9.3005
R1243 VDD2.n51 VDD2.n50 8.92171
R1244 VDD2.n18 VDD2.n17 8.92171
R1245 VDD2.n47 VDD2.n41 8.14595
R1246 VDD2.n14 VDD2.n8 8.14595
R1247 VDD2.n46 VDD2.n43 7.3702
R1248 VDD2.n13 VDD2.n10 7.3702
R1249 VDD2.n47 VDD2.n46 5.81868
R1250 VDD2.n14 VDD2.n13 5.81868
R1251 VDD2.n50 VDD2.n41 5.04292
R1252 VDD2.n17 VDD2.n8 5.04292
R1253 VDD2.n51 VDD2.n39 4.26717
R1254 VDD2.n18 VDD2.n6 4.26717
R1255 VDD2.n55 VDD2.n54 3.49141
R1256 VDD2.n22 VDD2.n21 3.49141
R1257 VDD2.n45 VDD2.n44 2.84308
R1258 VDD2.n12 VDD2.n11 2.84308
R1259 VDD2.n58 VDD2.n37 2.71565
R1260 VDD2.n25 VDD2.n4 2.71565
R1261 VDD2.n59 VDD2.n35 1.93989
R1262 VDD2.n26 VDD2.n2 1.93989
R1263 VDD2.n63 VDD2.n62 1.16414
R1264 VDD2.n30 VDD2.n29 1.16414
R1265 VDD2 VDD2.n66 0.463862
R1266 VDD2.n65 VDD2.n33 0.388379
R1267 VDD2.n32 VDD2.n0 0.388379
R1268 VDD2.n61 VDD2.n60 0.155672
R1269 VDD2.n60 VDD2.n36 0.155672
R1270 VDD2.n53 VDD2.n36 0.155672
R1271 VDD2.n53 VDD2.n52 0.155672
R1272 VDD2.n52 VDD2.n40 0.155672
R1273 VDD2.n45 VDD2.n40 0.155672
R1274 VDD2.n12 VDD2.n7 0.155672
R1275 VDD2.n19 VDD2.n7 0.155672
R1276 VDD2.n20 VDD2.n19 0.155672
R1277 VDD2.n20 VDD2.n3 0.155672
R1278 VDD2.n27 VDD2.n3 0.155672
R1279 VDD2.n28 VDD2.n27 0.155672
C0 VN VTAIL 1.36236f
C1 VN VDD1 0.147974f
C2 VTAIL VDD1 3.42468f
C3 VN VDD2 1.47018f
C4 VDD2 VTAIL 3.46867f
C5 VDD2 VDD1 0.550795f
C6 VN VP 3.93116f
C7 VP VTAIL 1.37663f
C8 VP VDD1 1.6091f
C9 VP VDD2 0.288799f
C10 VDD2 B 3.036266f
C11 VDD1 B 4.50249f
C12 VTAIL B 4.492227f
C13 VN B 6.72781f
C14 VP B 4.611297f
C15 VDD2.n0 B 0.008232f
C16 VDD2.n1 B 0.01862f
C17 VDD2.n2 B 0.008341f
C18 VDD2.n3 B 0.01466f
C19 VDD2.n4 B 0.007878f
C20 VDD2.n5 B 0.01862f
C21 VDD2.n6 B 0.008341f
C22 VDD2.n7 B 0.01466f
C23 VDD2.n8 B 0.007878f
C24 VDD2.n9 B 0.013965f
C25 VDD2.n10 B 0.013163f
C26 VDD2.t0 B 0.031044f
C27 VDD2.n11 B 0.074576f
C28 VDD2.n12 B 0.378252f
C29 VDD2.n13 B 0.007878f
C30 VDD2.n14 B 0.008341f
C31 VDD2.n15 B 0.01862f
C32 VDD2.n16 B 0.01862f
C33 VDD2.n17 B 0.008341f
C34 VDD2.n18 B 0.007878f
C35 VDD2.n19 B 0.01466f
C36 VDD2.n20 B 0.01466f
C37 VDD2.n21 B 0.007878f
C38 VDD2.n22 B 0.008341f
C39 VDD2.n23 B 0.01862f
C40 VDD2.n24 B 0.01862f
C41 VDD2.n25 B 0.008341f
C42 VDD2.n26 B 0.007878f
C43 VDD2.n27 B 0.01466f
C44 VDD2.n28 B 0.035889f
C45 VDD2.n29 B 0.007878f
C46 VDD2.n30 B 0.008341f
C47 VDD2.n31 B 0.036462f
C48 VDD2.n32 B 0.289498f
C49 VDD2.n33 B 0.008232f
C50 VDD2.n34 B 0.01862f
C51 VDD2.n35 B 0.008341f
C52 VDD2.n36 B 0.01466f
C53 VDD2.n37 B 0.007878f
C54 VDD2.n38 B 0.01862f
C55 VDD2.n39 B 0.008341f
C56 VDD2.n40 B 0.01466f
C57 VDD2.n41 B 0.007878f
C58 VDD2.n42 B 0.013965f
C59 VDD2.n43 B 0.013163f
C60 VDD2.t1 B 0.031044f
C61 VDD2.n44 B 0.074576f
C62 VDD2.n45 B 0.378252f
C63 VDD2.n46 B 0.007878f
C64 VDD2.n47 B 0.008341f
C65 VDD2.n48 B 0.01862f
C66 VDD2.n49 B 0.01862f
C67 VDD2.n50 B 0.008341f
C68 VDD2.n51 B 0.007878f
C69 VDD2.n52 B 0.01466f
C70 VDD2.n53 B 0.01466f
C71 VDD2.n54 B 0.007878f
C72 VDD2.n55 B 0.008341f
C73 VDD2.n56 B 0.01862f
C74 VDD2.n57 B 0.01862f
C75 VDD2.n58 B 0.008341f
C76 VDD2.n59 B 0.007878f
C77 VDD2.n60 B 0.01466f
C78 VDD2.n61 B 0.035889f
C79 VDD2.n62 B 0.007878f
C80 VDD2.n63 B 0.008341f
C81 VDD2.n64 B 0.036462f
C82 VDD2.n65 B 0.040138f
C83 VDD2.n66 B 1.3295f
C84 VN.t1 B 0.847697f
C85 VN.t0 B 1.01644f
C86 VDD1.n0 B 0.007875f
C87 VDD1.n1 B 0.017813f
C88 VDD1.n2 B 0.007979f
C89 VDD1.n3 B 0.014025f
C90 VDD1.n4 B 0.007536f
C91 VDD1.n5 B 0.017813f
C92 VDD1.n6 B 0.007979f
C93 VDD1.n7 B 0.014025f
C94 VDD1.n8 B 0.007536f
C95 VDD1.n9 B 0.01336f
C96 VDD1.n10 B 0.012592f
C97 VDD1.t0 B 0.029698f
C98 VDD1.n11 B 0.071342f
C99 VDD1.n12 B 0.361847f
C100 VDD1.n13 B 0.007536f
C101 VDD1.n14 B 0.007979f
C102 VDD1.n15 B 0.017813f
C103 VDD1.n16 B 0.017813f
C104 VDD1.n17 B 0.007979f
C105 VDD1.n18 B 0.007536f
C106 VDD1.n19 B 0.014025f
C107 VDD1.n20 B 0.014025f
C108 VDD1.n21 B 0.007536f
C109 VDD1.n22 B 0.007979f
C110 VDD1.n23 B 0.017813f
C111 VDD1.n24 B 0.017813f
C112 VDD1.n25 B 0.007979f
C113 VDD1.n26 B 0.007536f
C114 VDD1.n27 B 0.014025f
C115 VDD1.n28 B 0.034333f
C116 VDD1.n29 B 0.007536f
C117 VDD1.n30 B 0.007979f
C118 VDD1.n31 B 0.03488f
C119 VDD1.n32 B 0.038842f
C120 VDD1.n33 B 0.007875f
C121 VDD1.n34 B 0.017813f
C122 VDD1.n35 B 0.007979f
C123 VDD1.n36 B 0.014025f
C124 VDD1.n37 B 0.007536f
C125 VDD1.n38 B 0.017813f
C126 VDD1.n39 B 0.007979f
C127 VDD1.n40 B 0.014025f
C128 VDD1.n41 B 0.007536f
C129 VDD1.n42 B 0.01336f
C130 VDD1.n43 B 0.012592f
C131 VDD1.t1 B 0.029698f
C132 VDD1.n44 B 0.071342f
C133 VDD1.n45 B 0.361847f
C134 VDD1.n46 B 0.007536f
C135 VDD1.n47 B 0.007979f
C136 VDD1.n48 B 0.017813f
C137 VDD1.n49 B 0.017813f
C138 VDD1.n50 B 0.007979f
C139 VDD1.n51 B 0.007536f
C140 VDD1.n52 B 0.014025f
C141 VDD1.n53 B 0.014025f
C142 VDD1.n54 B 0.007536f
C143 VDD1.n55 B 0.007979f
C144 VDD1.n56 B 0.017813f
C145 VDD1.n57 B 0.017813f
C146 VDD1.n58 B 0.007979f
C147 VDD1.n59 B 0.007536f
C148 VDD1.n60 B 0.014025f
C149 VDD1.n61 B 0.034333f
C150 VDD1.n62 B 0.007536f
C151 VDD1.n63 B 0.007979f
C152 VDD1.n64 B 0.03488f
C153 VDD1.n65 B 0.296738f
C154 VTAIL.n0 B 0.009038f
C155 VTAIL.n1 B 0.020444f
C156 VTAIL.n2 B 0.009158f
C157 VTAIL.n3 B 0.016096f
C158 VTAIL.n4 B 0.008649f
C159 VTAIL.n5 B 0.020444f
C160 VTAIL.n6 B 0.009158f
C161 VTAIL.n7 B 0.016096f
C162 VTAIL.n8 B 0.008649f
C163 VTAIL.n9 B 0.015333f
C164 VTAIL.n10 B 0.014452f
C165 VTAIL.t3 B 0.034084f
C166 VTAIL.n11 B 0.08188f
C167 VTAIL.n12 B 0.415297f
C168 VTAIL.n13 B 0.008649f
C169 VTAIL.n14 B 0.009158f
C170 VTAIL.n15 B 0.020444f
C171 VTAIL.n16 B 0.020444f
C172 VTAIL.n17 B 0.009158f
C173 VTAIL.n18 B 0.008649f
C174 VTAIL.n19 B 0.016096f
C175 VTAIL.n20 B 0.016096f
C176 VTAIL.n21 B 0.008649f
C177 VTAIL.n22 B 0.009158f
C178 VTAIL.n23 B 0.020444f
C179 VTAIL.n24 B 0.020444f
C180 VTAIL.n25 B 0.009158f
C181 VTAIL.n26 B 0.008649f
C182 VTAIL.n27 B 0.016096f
C183 VTAIL.n28 B 0.039405f
C184 VTAIL.n29 B 0.008649f
C185 VTAIL.n30 B 0.009158f
C186 VTAIL.n31 B 0.040033f
C187 VTAIL.n32 B 0.032969f
C188 VTAIL.n33 B 0.738743f
C189 VTAIL.n34 B 0.009038f
C190 VTAIL.n35 B 0.020444f
C191 VTAIL.n36 B 0.009158f
C192 VTAIL.n37 B 0.016096f
C193 VTAIL.n38 B 0.008649f
C194 VTAIL.n39 B 0.020444f
C195 VTAIL.n40 B 0.009158f
C196 VTAIL.n41 B 0.016096f
C197 VTAIL.n42 B 0.008649f
C198 VTAIL.n43 B 0.015333f
C199 VTAIL.n44 B 0.014452f
C200 VTAIL.t0 B 0.034084f
C201 VTAIL.n45 B 0.08188f
C202 VTAIL.n46 B 0.415297f
C203 VTAIL.n47 B 0.008649f
C204 VTAIL.n48 B 0.009158f
C205 VTAIL.n49 B 0.020444f
C206 VTAIL.n50 B 0.020444f
C207 VTAIL.n51 B 0.009158f
C208 VTAIL.n52 B 0.008649f
C209 VTAIL.n53 B 0.016096f
C210 VTAIL.n54 B 0.016096f
C211 VTAIL.n55 B 0.008649f
C212 VTAIL.n56 B 0.009158f
C213 VTAIL.n57 B 0.020444f
C214 VTAIL.n58 B 0.020444f
C215 VTAIL.n59 B 0.009158f
C216 VTAIL.n60 B 0.008649f
C217 VTAIL.n61 B 0.016096f
C218 VTAIL.n62 B 0.039405f
C219 VTAIL.n63 B 0.008649f
C220 VTAIL.n64 B 0.009158f
C221 VTAIL.n65 B 0.040033f
C222 VTAIL.n66 B 0.032969f
C223 VTAIL.n67 B 0.756739f
C224 VTAIL.n68 B 0.009038f
C225 VTAIL.n69 B 0.020444f
C226 VTAIL.n70 B 0.009158f
C227 VTAIL.n71 B 0.016096f
C228 VTAIL.n72 B 0.008649f
C229 VTAIL.n73 B 0.020444f
C230 VTAIL.n74 B 0.009158f
C231 VTAIL.n75 B 0.016096f
C232 VTAIL.n76 B 0.008649f
C233 VTAIL.n77 B 0.015333f
C234 VTAIL.n78 B 0.014452f
C235 VTAIL.t2 B 0.034084f
C236 VTAIL.n79 B 0.08188f
C237 VTAIL.n80 B 0.415297f
C238 VTAIL.n81 B 0.008649f
C239 VTAIL.n82 B 0.009158f
C240 VTAIL.n83 B 0.020444f
C241 VTAIL.n84 B 0.020444f
C242 VTAIL.n85 B 0.009158f
C243 VTAIL.n86 B 0.008649f
C244 VTAIL.n87 B 0.016096f
C245 VTAIL.n88 B 0.016096f
C246 VTAIL.n89 B 0.008649f
C247 VTAIL.n90 B 0.009158f
C248 VTAIL.n91 B 0.020444f
C249 VTAIL.n92 B 0.020444f
C250 VTAIL.n93 B 0.009158f
C251 VTAIL.n94 B 0.008649f
C252 VTAIL.n95 B 0.016096f
C253 VTAIL.n96 B 0.039405f
C254 VTAIL.n97 B 0.008649f
C255 VTAIL.n98 B 0.009158f
C256 VTAIL.n99 B 0.040033f
C257 VTAIL.n100 B 0.032969f
C258 VTAIL.n101 B 0.672681f
C259 VTAIL.n102 B 0.009038f
C260 VTAIL.n103 B 0.020444f
C261 VTAIL.n104 B 0.009158f
C262 VTAIL.n105 B 0.016096f
C263 VTAIL.n106 B 0.008649f
C264 VTAIL.n107 B 0.020444f
C265 VTAIL.n108 B 0.009158f
C266 VTAIL.n109 B 0.016096f
C267 VTAIL.n110 B 0.008649f
C268 VTAIL.n111 B 0.015333f
C269 VTAIL.n112 B 0.014452f
C270 VTAIL.t1 B 0.034084f
C271 VTAIL.n113 B 0.08188f
C272 VTAIL.n114 B 0.415297f
C273 VTAIL.n115 B 0.008649f
C274 VTAIL.n116 B 0.009158f
C275 VTAIL.n117 B 0.020444f
C276 VTAIL.n118 B 0.020444f
C277 VTAIL.n119 B 0.009158f
C278 VTAIL.n120 B 0.008649f
C279 VTAIL.n121 B 0.016096f
C280 VTAIL.n122 B 0.016096f
C281 VTAIL.n123 B 0.008649f
C282 VTAIL.n124 B 0.009158f
C283 VTAIL.n125 B 0.020444f
C284 VTAIL.n126 B 0.020444f
C285 VTAIL.n127 B 0.009158f
C286 VTAIL.n128 B 0.008649f
C287 VTAIL.n129 B 0.016096f
C288 VTAIL.n130 B 0.039405f
C289 VTAIL.n131 B 0.008649f
C290 VTAIL.n132 B 0.009158f
C291 VTAIL.n133 B 0.040033f
C292 VTAIL.n134 B 0.032969f
C293 VTAIL.n135 B 0.624281f
C294 VP.t1 B 1.02236f
C295 VP.t0 B 0.855229f
C296 VP.n0 B 1.99549f
.ends

