* NGSPICE file created from diff_pair_sample_0381.ext - technology: sky130A

.subckt diff_pair_sample_0381 VTAIL VN VP B VDD2 VDD1
X0 B.t19 B.t17 B.t18 B.t14 sky130_fd_pr__nfet_01v8 ad=1.7901 pd=9.96 as=0 ps=0 w=4.59 l=1.54
X1 VDD1.t5 VP.t0 VTAIL.t7 B.t3 sky130_fd_pr__nfet_01v8 ad=1.7901 pd=9.96 as=0.75735 ps=4.92 w=4.59 l=1.54
X2 VTAIL.t5 VP.t1 VDD1.t4 B.t2 sky130_fd_pr__nfet_01v8 ad=0.75735 pd=4.92 as=0.75735 ps=4.92 w=4.59 l=1.54
X3 VDD1.t3 VP.t2 VTAIL.t9 B.t4 sky130_fd_pr__nfet_01v8 ad=0.75735 pd=4.92 as=1.7901 ps=9.96 w=4.59 l=1.54
X4 VDD2.t5 VN.t0 VTAIL.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=0.75735 pd=4.92 as=1.7901 ps=9.96 w=4.59 l=1.54
X5 VTAIL.t10 VP.t3 VDD1.t2 B.t5 sky130_fd_pr__nfet_01v8 ad=0.75735 pd=4.92 as=0.75735 ps=4.92 w=4.59 l=1.54
X6 B.t16 B.t13 B.t15 B.t14 sky130_fd_pr__nfet_01v8 ad=1.7901 pd=9.96 as=0 ps=0 w=4.59 l=1.54
X7 VTAIL.t11 VN.t1 VDD2.t4 B.t5 sky130_fd_pr__nfet_01v8 ad=0.75735 pd=4.92 as=0.75735 ps=4.92 w=4.59 l=1.54
X8 VDD2.t3 VN.t2 VTAIL.t2 B.t3 sky130_fd_pr__nfet_01v8 ad=1.7901 pd=9.96 as=0.75735 ps=4.92 w=4.59 l=1.54
X9 B.t12 B.t10 B.t11 B.t7 sky130_fd_pr__nfet_01v8 ad=1.7901 pd=9.96 as=0 ps=0 w=4.59 l=1.54
X10 VDD2.t2 VN.t3 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=0.75735 pd=4.92 as=1.7901 ps=9.96 w=4.59 l=1.54
X11 VDD1.t1 VP.t4 VTAIL.t6 B.t1 sky130_fd_pr__nfet_01v8 ad=1.7901 pd=9.96 as=0.75735 ps=4.92 w=4.59 l=1.54
X12 B.t9 B.t6 B.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=1.7901 pd=9.96 as=0 ps=0 w=4.59 l=1.54
X13 VDD2.t1 VN.t4 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=1.7901 pd=9.96 as=0.75735 ps=4.92 w=4.59 l=1.54
X14 VTAIL.t3 VN.t5 VDD2.t0 B.t2 sky130_fd_pr__nfet_01v8 ad=0.75735 pd=4.92 as=0.75735 ps=4.92 w=4.59 l=1.54
X15 VDD1.t0 VP.t5 VTAIL.t8 B.t0 sky130_fd_pr__nfet_01v8 ad=0.75735 pd=4.92 as=1.7901 ps=9.96 w=4.59 l=1.54
R0 B.n401 B.n86 585
R1 B.n86 B.n57 585
R2 B.n403 B.n402 585
R3 B.n405 B.n85 585
R4 B.n408 B.n407 585
R5 B.n409 B.n84 585
R6 B.n411 B.n410 585
R7 B.n413 B.n83 585
R8 B.n416 B.n415 585
R9 B.n417 B.n82 585
R10 B.n419 B.n418 585
R11 B.n421 B.n81 585
R12 B.n424 B.n423 585
R13 B.n425 B.n80 585
R14 B.n427 B.n426 585
R15 B.n429 B.n79 585
R16 B.n432 B.n431 585
R17 B.n433 B.n78 585
R18 B.n435 B.n434 585
R19 B.n437 B.n77 585
R20 B.n440 B.n439 585
R21 B.n442 B.n74 585
R22 B.n444 B.n443 585
R23 B.n446 B.n73 585
R24 B.n449 B.n448 585
R25 B.n450 B.n72 585
R26 B.n452 B.n451 585
R27 B.n454 B.n71 585
R28 B.n457 B.n456 585
R29 B.n458 B.n68 585
R30 B.n461 B.n460 585
R31 B.n463 B.n67 585
R32 B.n466 B.n465 585
R33 B.n467 B.n66 585
R34 B.n469 B.n468 585
R35 B.n471 B.n65 585
R36 B.n474 B.n473 585
R37 B.n475 B.n64 585
R38 B.n477 B.n476 585
R39 B.n479 B.n63 585
R40 B.n482 B.n481 585
R41 B.n483 B.n62 585
R42 B.n485 B.n484 585
R43 B.n487 B.n61 585
R44 B.n490 B.n489 585
R45 B.n491 B.n60 585
R46 B.n493 B.n492 585
R47 B.n495 B.n59 585
R48 B.n498 B.n497 585
R49 B.n499 B.n58 585
R50 B.n400 B.n56 585
R51 B.n502 B.n56 585
R52 B.n399 B.n55 585
R53 B.n503 B.n55 585
R54 B.n398 B.n54 585
R55 B.n504 B.n54 585
R56 B.n397 B.n396 585
R57 B.n396 B.n50 585
R58 B.n395 B.n49 585
R59 B.n510 B.n49 585
R60 B.n394 B.n48 585
R61 B.n511 B.n48 585
R62 B.n393 B.n47 585
R63 B.n512 B.n47 585
R64 B.n392 B.n391 585
R65 B.n391 B.n43 585
R66 B.n390 B.n42 585
R67 B.n518 B.n42 585
R68 B.n389 B.n41 585
R69 B.n519 B.n41 585
R70 B.n388 B.n40 585
R71 B.n520 B.n40 585
R72 B.n387 B.n386 585
R73 B.n386 B.n36 585
R74 B.n385 B.n35 585
R75 B.n526 B.n35 585
R76 B.n384 B.n34 585
R77 B.n527 B.n34 585
R78 B.n383 B.n33 585
R79 B.n528 B.n33 585
R80 B.n382 B.n381 585
R81 B.n381 B.n29 585
R82 B.n380 B.n28 585
R83 B.n534 B.n28 585
R84 B.n379 B.n27 585
R85 B.n535 B.n27 585
R86 B.n378 B.n26 585
R87 B.n536 B.n26 585
R88 B.n377 B.n376 585
R89 B.n376 B.n22 585
R90 B.n375 B.n21 585
R91 B.n542 B.n21 585
R92 B.n374 B.n20 585
R93 B.n543 B.n20 585
R94 B.n373 B.n19 585
R95 B.n544 B.n19 585
R96 B.n372 B.n371 585
R97 B.n371 B.n15 585
R98 B.n370 B.n14 585
R99 B.n550 B.n14 585
R100 B.n369 B.n13 585
R101 B.n551 B.n13 585
R102 B.n368 B.n12 585
R103 B.n552 B.n12 585
R104 B.n367 B.n366 585
R105 B.n366 B.n8 585
R106 B.n365 B.n7 585
R107 B.n558 B.n7 585
R108 B.n364 B.n6 585
R109 B.n559 B.n6 585
R110 B.n363 B.n5 585
R111 B.n560 B.n5 585
R112 B.n362 B.n361 585
R113 B.n361 B.n4 585
R114 B.n360 B.n87 585
R115 B.n360 B.n359 585
R116 B.n350 B.n88 585
R117 B.n89 B.n88 585
R118 B.n352 B.n351 585
R119 B.n353 B.n352 585
R120 B.n349 B.n93 585
R121 B.n97 B.n93 585
R122 B.n348 B.n347 585
R123 B.n347 B.n346 585
R124 B.n95 B.n94 585
R125 B.n96 B.n95 585
R126 B.n339 B.n338 585
R127 B.n340 B.n339 585
R128 B.n337 B.n102 585
R129 B.n102 B.n101 585
R130 B.n336 B.n335 585
R131 B.n335 B.n334 585
R132 B.n104 B.n103 585
R133 B.n105 B.n104 585
R134 B.n327 B.n326 585
R135 B.n328 B.n327 585
R136 B.n325 B.n110 585
R137 B.n110 B.n109 585
R138 B.n324 B.n323 585
R139 B.n323 B.n322 585
R140 B.n112 B.n111 585
R141 B.n113 B.n112 585
R142 B.n315 B.n314 585
R143 B.n316 B.n315 585
R144 B.n313 B.n118 585
R145 B.n118 B.n117 585
R146 B.n312 B.n311 585
R147 B.n311 B.n310 585
R148 B.n120 B.n119 585
R149 B.n121 B.n120 585
R150 B.n303 B.n302 585
R151 B.n304 B.n303 585
R152 B.n301 B.n126 585
R153 B.n126 B.n125 585
R154 B.n300 B.n299 585
R155 B.n299 B.n298 585
R156 B.n128 B.n127 585
R157 B.n129 B.n128 585
R158 B.n291 B.n290 585
R159 B.n292 B.n291 585
R160 B.n289 B.n133 585
R161 B.n137 B.n133 585
R162 B.n288 B.n287 585
R163 B.n287 B.n286 585
R164 B.n135 B.n134 585
R165 B.n136 B.n135 585
R166 B.n279 B.n278 585
R167 B.n280 B.n279 585
R168 B.n277 B.n142 585
R169 B.n142 B.n141 585
R170 B.n276 B.n275 585
R171 B.n275 B.n274 585
R172 B.n271 B.n146 585
R173 B.n270 B.n269 585
R174 B.n267 B.n147 585
R175 B.n267 B.n145 585
R176 B.n266 B.n265 585
R177 B.n264 B.n263 585
R178 B.n262 B.n149 585
R179 B.n260 B.n259 585
R180 B.n258 B.n150 585
R181 B.n257 B.n256 585
R182 B.n254 B.n151 585
R183 B.n252 B.n251 585
R184 B.n250 B.n152 585
R185 B.n249 B.n248 585
R186 B.n246 B.n153 585
R187 B.n244 B.n243 585
R188 B.n242 B.n154 585
R189 B.n241 B.n240 585
R190 B.n238 B.n155 585
R191 B.n236 B.n235 585
R192 B.n234 B.n156 585
R193 B.n232 B.n231 585
R194 B.n229 B.n159 585
R195 B.n227 B.n226 585
R196 B.n225 B.n160 585
R197 B.n224 B.n223 585
R198 B.n221 B.n161 585
R199 B.n219 B.n218 585
R200 B.n217 B.n162 585
R201 B.n216 B.n215 585
R202 B.n213 B.n212 585
R203 B.n211 B.n210 585
R204 B.n209 B.n167 585
R205 B.n207 B.n206 585
R206 B.n205 B.n168 585
R207 B.n204 B.n203 585
R208 B.n201 B.n169 585
R209 B.n199 B.n198 585
R210 B.n197 B.n170 585
R211 B.n196 B.n195 585
R212 B.n193 B.n171 585
R213 B.n191 B.n190 585
R214 B.n189 B.n172 585
R215 B.n188 B.n187 585
R216 B.n185 B.n173 585
R217 B.n183 B.n182 585
R218 B.n181 B.n174 585
R219 B.n180 B.n179 585
R220 B.n177 B.n175 585
R221 B.n144 B.n143 585
R222 B.n273 B.n272 585
R223 B.n274 B.n273 585
R224 B.n140 B.n139 585
R225 B.n141 B.n140 585
R226 B.n282 B.n281 585
R227 B.n281 B.n280 585
R228 B.n283 B.n138 585
R229 B.n138 B.n136 585
R230 B.n285 B.n284 585
R231 B.n286 B.n285 585
R232 B.n132 B.n131 585
R233 B.n137 B.n132 585
R234 B.n294 B.n293 585
R235 B.n293 B.n292 585
R236 B.n295 B.n130 585
R237 B.n130 B.n129 585
R238 B.n297 B.n296 585
R239 B.n298 B.n297 585
R240 B.n124 B.n123 585
R241 B.n125 B.n124 585
R242 B.n306 B.n305 585
R243 B.n305 B.n304 585
R244 B.n307 B.n122 585
R245 B.n122 B.n121 585
R246 B.n309 B.n308 585
R247 B.n310 B.n309 585
R248 B.n116 B.n115 585
R249 B.n117 B.n116 585
R250 B.n318 B.n317 585
R251 B.n317 B.n316 585
R252 B.n319 B.n114 585
R253 B.n114 B.n113 585
R254 B.n321 B.n320 585
R255 B.n322 B.n321 585
R256 B.n108 B.n107 585
R257 B.n109 B.n108 585
R258 B.n330 B.n329 585
R259 B.n329 B.n328 585
R260 B.n331 B.n106 585
R261 B.n106 B.n105 585
R262 B.n333 B.n332 585
R263 B.n334 B.n333 585
R264 B.n100 B.n99 585
R265 B.n101 B.n100 585
R266 B.n342 B.n341 585
R267 B.n341 B.n340 585
R268 B.n343 B.n98 585
R269 B.n98 B.n96 585
R270 B.n345 B.n344 585
R271 B.n346 B.n345 585
R272 B.n92 B.n91 585
R273 B.n97 B.n92 585
R274 B.n355 B.n354 585
R275 B.n354 B.n353 585
R276 B.n356 B.n90 585
R277 B.n90 B.n89 585
R278 B.n358 B.n357 585
R279 B.n359 B.n358 585
R280 B.n2 B.n0 585
R281 B.n4 B.n2 585
R282 B.n3 B.n1 585
R283 B.n559 B.n3 585
R284 B.n557 B.n556 585
R285 B.n558 B.n557 585
R286 B.n555 B.n9 585
R287 B.n9 B.n8 585
R288 B.n554 B.n553 585
R289 B.n553 B.n552 585
R290 B.n11 B.n10 585
R291 B.n551 B.n11 585
R292 B.n549 B.n548 585
R293 B.n550 B.n549 585
R294 B.n547 B.n16 585
R295 B.n16 B.n15 585
R296 B.n546 B.n545 585
R297 B.n545 B.n544 585
R298 B.n18 B.n17 585
R299 B.n543 B.n18 585
R300 B.n541 B.n540 585
R301 B.n542 B.n541 585
R302 B.n539 B.n23 585
R303 B.n23 B.n22 585
R304 B.n538 B.n537 585
R305 B.n537 B.n536 585
R306 B.n25 B.n24 585
R307 B.n535 B.n25 585
R308 B.n533 B.n532 585
R309 B.n534 B.n533 585
R310 B.n531 B.n30 585
R311 B.n30 B.n29 585
R312 B.n530 B.n529 585
R313 B.n529 B.n528 585
R314 B.n32 B.n31 585
R315 B.n527 B.n32 585
R316 B.n525 B.n524 585
R317 B.n526 B.n525 585
R318 B.n523 B.n37 585
R319 B.n37 B.n36 585
R320 B.n522 B.n521 585
R321 B.n521 B.n520 585
R322 B.n39 B.n38 585
R323 B.n519 B.n39 585
R324 B.n517 B.n516 585
R325 B.n518 B.n517 585
R326 B.n515 B.n44 585
R327 B.n44 B.n43 585
R328 B.n514 B.n513 585
R329 B.n513 B.n512 585
R330 B.n46 B.n45 585
R331 B.n511 B.n46 585
R332 B.n509 B.n508 585
R333 B.n510 B.n509 585
R334 B.n507 B.n51 585
R335 B.n51 B.n50 585
R336 B.n506 B.n505 585
R337 B.n505 B.n504 585
R338 B.n53 B.n52 585
R339 B.n503 B.n53 585
R340 B.n501 B.n500 585
R341 B.n502 B.n501 585
R342 B.n562 B.n561 585
R343 B.n561 B.n560 585
R344 B.n273 B.n146 535.745
R345 B.n501 B.n58 535.745
R346 B.n275 B.n144 535.745
R347 B.n86 B.n56 535.745
R348 B.n163 B.t10 277.416
R349 B.n157 B.t6 277.416
R350 B.n69 B.t17 277.416
R351 B.n75 B.t13 277.416
R352 B.n404 B.n57 256.663
R353 B.n406 B.n57 256.663
R354 B.n412 B.n57 256.663
R355 B.n414 B.n57 256.663
R356 B.n420 B.n57 256.663
R357 B.n422 B.n57 256.663
R358 B.n428 B.n57 256.663
R359 B.n430 B.n57 256.663
R360 B.n436 B.n57 256.663
R361 B.n438 B.n57 256.663
R362 B.n445 B.n57 256.663
R363 B.n447 B.n57 256.663
R364 B.n453 B.n57 256.663
R365 B.n455 B.n57 256.663
R366 B.n462 B.n57 256.663
R367 B.n464 B.n57 256.663
R368 B.n470 B.n57 256.663
R369 B.n472 B.n57 256.663
R370 B.n478 B.n57 256.663
R371 B.n480 B.n57 256.663
R372 B.n486 B.n57 256.663
R373 B.n488 B.n57 256.663
R374 B.n494 B.n57 256.663
R375 B.n496 B.n57 256.663
R376 B.n268 B.n145 256.663
R377 B.n148 B.n145 256.663
R378 B.n261 B.n145 256.663
R379 B.n255 B.n145 256.663
R380 B.n253 B.n145 256.663
R381 B.n247 B.n145 256.663
R382 B.n245 B.n145 256.663
R383 B.n239 B.n145 256.663
R384 B.n237 B.n145 256.663
R385 B.n230 B.n145 256.663
R386 B.n228 B.n145 256.663
R387 B.n222 B.n145 256.663
R388 B.n220 B.n145 256.663
R389 B.n214 B.n145 256.663
R390 B.n166 B.n145 256.663
R391 B.n208 B.n145 256.663
R392 B.n202 B.n145 256.663
R393 B.n200 B.n145 256.663
R394 B.n194 B.n145 256.663
R395 B.n192 B.n145 256.663
R396 B.n186 B.n145 256.663
R397 B.n184 B.n145 256.663
R398 B.n178 B.n145 256.663
R399 B.n176 B.n145 256.663
R400 B.n163 B.t12 191.103
R401 B.n75 B.t15 191.103
R402 B.n157 B.t9 191.103
R403 B.n69 B.t18 191.103
R404 B.n273 B.n140 163.367
R405 B.n281 B.n140 163.367
R406 B.n281 B.n138 163.367
R407 B.n285 B.n138 163.367
R408 B.n285 B.n132 163.367
R409 B.n293 B.n132 163.367
R410 B.n293 B.n130 163.367
R411 B.n297 B.n130 163.367
R412 B.n297 B.n124 163.367
R413 B.n305 B.n124 163.367
R414 B.n305 B.n122 163.367
R415 B.n309 B.n122 163.367
R416 B.n309 B.n116 163.367
R417 B.n317 B.n116 163.367
R418 B.n317 B.n114 163.367
R419 B.n321 B.n114 163.367
R420 B.n321 B.n108 163.367
R421 B.n329 B.n108 163.367
R422 B.n329 B.n106 163.367
R423 B.n333 B.n106 163.367
R424 B.n333 B.n100 163.367
R425 B.n341 B.n100 163.367
R426 B.n341 B.n98 163.367
R427 B.n345 B.n98 163.367
R428 B.n345 B.n92 163.367
R429 B.n354 B.n92 163.367
R430 B.n354 B.n90 163.367
R431 B.n358 B.n90 163.367
R432 B.n358 B.n2 163.367
R433 B.n561 B.n2 163.367
R434 B.n561 B.n3 163.367
R435 B.n557 B.n3 163.367
R436 B.n557 B.n9 163.367
R437 B.n553 B.n9 163.367
R438 B.n553 B.n11 163.367
R439 B.n549 B.n11 163.367
R440 B.n549 B.n16 163.367
R441 B.n545 B.n16 163.367
R442 B.n545 B.n18 163.367
R443 B.n541 B.n18 163.367
R444 B.n541 B.n23 163.367
R445 B.n537 B.n23 163.367
R446 B.n537 B.n25 163.367
R447 B.n533 B.n25 163.367
R448 B.n533 B.n30 163.367
R449 B.n529 B.n30 163.367
R450 B.n529 B.n32 163.367
R451 B.n525 B.n32 163.367
R452 B.n525 B.n37 163.367
R453 B.n521 B.n37 163.367
R454 B.n521 B.n39 163.367
R455 B.n517 B.n39 163.367
R456 B.n517 B.n44 163.367
R457 B.n513 B.n44 163.367
R458 B.n513 B.n46 163.367
R459 B.n509 B.n46 163.367
R460 B.n509 B.n51 163.367
R461 B.n505 B.n51 163.367
R462 B.n505 B.n53 163.367
R463 B.n501 B.n53 163.367
R464 B.n269 B.n267 163.367
R465 B.n267 B.n266 163.367
R466 B.n263 B.n262 163.367
R467 B.n260 B.n150 163.367
R468 B.n256 B.n254 163.367
R469 B.n252 B.n152 163.367
R470 B.n248 B.n246 163.367
R471 B.n244 B.n154 163.367
R472 B.n240 B.n238 163.367
R473 B.n236 B.n156 163.367
R474 B.n231 B.n229 163.367
R475 B.n227 B.n160 163.367
R476 B.n223 B.n221 163.367
R477 B.n219 B.n162 163.367
R478 B.n215 B.n213 163.367
R479 B.n210 B.n209 163.367
R480 B.n207 B.n168 163.367
R481 B.n203 B.n201 163.367
R482 B.n199 B.n170 163.367
R483 B.n195 B.n193 163.367
R484 B.n191 B.n172 163.367
R485 B.n187 B.n185 163.367
R486 B.n183 B.n174 163.367
R487 B.n179 B.n177 163.367
R488 B.n275 B.n142 163.367
R489 B.n279 B.n142 163.367
R490 B.n279 B.n135 163.367
R491 B.n287 B.n135 163.367
R492 B.n287 B.n133 163.367
R493 B.n291 B.n133 163.367
R494 B.n291 B.n128 163.367
R495 B.n299 B.n128 163.367
R496 B.n299 B.n126 163.367
R497 B.n303 B.n126 163.367
R498 B.n303 B.n120 163.367
R499 B.n311 B.n120 163.367
R500 B.n311 B.n118 163.367
R501 B.n315 B.n118 163.367
R502 B.n315 B.n112 163.367
R503 B.n323 B.n112 163.367
R504 B.n323 B.n110 163.367
R505 B.n327 B.n110 163.367
R506 B.n327 B.n104 163.367
R507 B.n335 B.n104 163.367
R508 B.n335 B.n102 163.367
R509 B.n339 B.n102 163.367
R510 B.n339 B.n95 163.367
R511 B.n347 B.n95 163.367
R512 B.n347 B.n93 163.367
R513 B.n352 B.n93 163.367
R514 B.n352 B.n88 163.367
R515 B.n360 B.n88 163.367
R516 B.n361 B.n360 163.367
R517 B.n361 B.n5 163.367
R518 B.n6 B.n5 163.367
R519 B.n7 B.n6 163.367
R520 B.n366 B.n7 163.367
R521 B.n366 B.n12 163.367
R522 B.n13 B.n12 163.367
R523 B.n14 B.n13 163.367
R524 B.n371 B.n14 163.367
R525 B.n371 B.n19 163.367
R526 B.n20 B.n19 163.367
R527 B.n21 B.n20 163.367
R528 B.n376 B.n21 163.367
R529 B.n376 B.n26 163.367
R530 B.n27 B.n26 163.367
R531 B.n28 B.n27 163.367
R532 B.n381 B.n28 163.367
R533 B.n381 B.n33 163.367
R534 B.n34 B.n33 163.367
R535 B.n35 B.n34 163.367
R536 B.n386 B.n35 163.367
R537 B.n386 B.n40 163.367
R538 B.n41 B.n40 163.367
R539 B.n42 B.n41 163.367
R540 B.n391 B.n42 163.367
R541 B.n391 B.n47 163.367
R542 B.n48 B.n47 163.367
R543 B.n49 B.n48 163.367
R544 B.n396 B.n49 163.367
R545 B.n396 B.n54 163.367
R546 B.n55 B.n54 163.367
R547 B.n56 B.n55 163.367
R548 B.n497 B.n495 163.367
R549 B.n493 B.n60 163.367
R550 B.n489 B.n487 163.367
R551 B.n485 B.n62 163.367
R552 B.n481 B.n479 163.367
R553 B.n477 B.n64 163.367
R554 B.n473 B.n471 163.367
R555 B.n469 B.n66 163.367
R556 B.n465 B.n463 163.367
R557 B.n461 B.n68 163.367
R558 B.n456 B.n454 163.367
R559 B.n452 B.n72 163.367
R560 B.n448 B.n446 163.367
R561 B.n444 B.n74 163.367
R562 B.n439 B.n437 163.367
R563 B.n435 B.n78 163.367
R564 B.n431 B.n429 163.367
R565 B.n427 B.n80 163.367
R566 B.n423 B.n421 163.367
R567 B.n419 B.n82 163.367
R568 B.n415 B.n413 163.367
R569 B.n411 B.n84 163.367
R570 B.n407 B.n405 163.367
R571 B.n403 B.n86 163.367
R572 B.n164 B.t11 154.837
R573 B.n76 B.t16 154.837
R574 B.n158 B.t8 154.837
R575 B.n70 B.t19 154.837
R576 B.n274 B.n145 146.072
R577 B.n502 B.n57 146.072
R578 B.n274 B.n141 75.8241
R579 B.n280 B.n141 75.8241
R580 B.n280 B.n136 75.8241
R581 B.n286 B.n136 75.8241
R582 B.n286 B.n137 75.8241
R583 B.n292 B.n129 75.8241
R584 B.n298 B.n129 75.8241
R585 B.n298 B.n125 75.8241
R586 B.n304 B.n125 75.8241
R587 B.n304 B.n121 75.8241
R588 B.n310 B.n121 75.8241
R589 B.n310 B.n117 75.8241
R590 B.n316 B.n117 75.8241
R591 B.n322 B.n113 75.8241
R592 B.n322 B.n109 75.8241
R593 B.n328 B.n109 75.8241
R594 B.n328 B.n105 75.8241
R595 B.n334 B.n105 75.8241
R596 B.n340 B.n101 75.8241
R597 B.n340 B.n96 75.8241
R598 B.n346 B.n96 75.8241
R599 B.n346 B.n97 75.8241
R600 B.n353 B.n89 75.8241
R601 B.n359 B.n89 75.8241
R602 B.n359 B.n4 75.8241
R603 B.n560 B.n4 75.8241
R604 B.n560 B.n559 75.8241
R605 B.n559 B.n558 75.8241
R606 B.n558 B.n8 75.8241
R607 B.n552 B.n8 75.8241
R608 B.n551 B.n550 75.8241
R609 B.n550 B.n15 75.8241
R610 B.n544 B.n15 75.8241
R611 B.n544 B.n543 75.8241
R612 B.n542 B.n22 75.8241
R613 B.n536 B.n22 75.8241
R614 B.n536 B.n535 75.8241
R615 B.n535 B.n534 75.8241
R616 B.n534 B.n29 75.8241
R617 B.n528 B.n527 75.8241
R618 B.n527 B.n526 75.8241
R619 B.n526 B.n36 75.8241
R620 B.n520 B.n36 75.8241
R621 B.n520 B.n519 75.8241
R622 B.n519 B.n518 75.8241
R623 B.n518 B.n43 75.8241
R624 B.n512 B.n43 75.8241
R625 B.n511 B.n510 75.8241
R626 B.n510 B.n50 75.8241
R627 B.n504 B.n50 75.8241
R628 B.n504 B.n503 75.8241
R629 B.n503 B.n502 75.8241
R630 B.n268 B.n146 71.676
R631 B.n266 B.n148 71.676
R632 B.n262 B.n261 71.676
R633 B.n255 B.n150 71.676
R634 B.n254 B.n253 71.676
R635 B.n247 B.n152 71.676
R636 B.n246 B.n245 71.676
R637 B.n239 B.n154 71.676
R638 B.n238 B.n237 71.676
R639 B.n230 B.n156 71.676
R640 B.n229 B.n228 71.676
R641 B.n222 B.n160 71.676
R642 B.n221 B.n220 71.676
R643 B.n214 B.n162 71.676
R644 B.n213 B.n166 71.676
R645 B.n209 B.n208 71.676
R646 B.n202 B.n168 71.676
R647 B.n201 B.n200 71.676
R648 B.n194 B.n170 71.676
R649 B.n193 B.n192 71.676
R650 B.n186 B.n172 71.676
R651 B.n185 B.n184 71.676
R652 B.n178 B.n174 71.676
R653 B.n177 B.n176 71.676
R654 B.n496 B.n58 71.676
R655 B.n495 B.n494 71.676
R656 B.n488 B.n60 71.676
R657 B.n487 B.n486 71.676
R658 B.n480 B.n62 71.676
R659 B.n479 B.n478 71.676
R660 B.n472 B.n64 71.676
R661 B.n471 B.n470 71.676
R662 B.n464 B.n66 71.676
R663 B.n463 B.n462 71.676
R664 B.n455 B.n68 71.676
R665 B.n454 B.n453 71.676
R666 B.n447 B.n72 71.676
R667 B.n446 B.n445 71.676
R668 B.n438 B.n74 71.676
R669 B.n437 B.n436 71.676
R670 B.n430 B.n78 71.676
R671 B.n429 B.n428 71.676
R672 B.n422 B.n80 71.676
R673 B.n421 B.n420 71.676
R674 B.n414 B.n82 71.676
R675 B.n413 B.n412 71.676
R676 B.n406 B.n84 71.676
R677 B.n405 B.n404 71.676
R678 B.n404 B.n403 71.676
R679 B.n407 B.n406 71.676
R680 B.n412 B.n411 71.676
R681 B.n415 B.n414 71.676
R682 B.n420 B.n419 71.676
R683 B.n423 B.n422 71.676
R684 B.n428 B.n427 71.676
R685 B.n431 B.n430 71.676
R686 B.n436 B.n435 71.676
R687 B.n439 B.n438 71.676
R688 B.n445 B.n444 71.676
R689 B.n448 B.n447 71.676
R690 B.n453 B.n452 71.676
R691 B.n456 B.n455 71.676
R692 B.n462 B.n461 71.676
R693 B.n465 B.n464 71.676
R694 B.n470 B.n469 71.676
R695 B.n473 B.n472 71.676
R696 B.n478 B.n477 71.676
R697 B.n481 B.n480 71.676
R698 B.n486 B.n485 71.676
R699 B.n489 B.n488 71.676
R700 B.n494 B.n493 71.676
R701 B.n497 B.n496 71.676
R702 B.n269 B.n268 71.676
R703 B.n263 B.n148 71.676
R704 B.n261 B.n260 71.676
R705 B.n256 B.n255 71.676
R706 B.n253 B.n252 71.676
R707 B.n248 B.n247 71.676
R708 B.n245 B.n244 71.676
R709 B.n240 B.n239 71.676
R710 B.n237 B.n236 71.676
R711 B.n231 B.n230 71.676
R712 B.n228 B.n227 71.676
R713 B.n223 B.n222 71.676
R714 B.n220 B.n219 71.676
R715 B.n215 B.n214 71.676
R716 B.n210 B.n166 71.676
R717 B.n208 B.n207 71.676
R718 B.n203 B.n202 71.676
R719 B.n200 B.n199 71.676
R720 B.n195 B.n194 71.676
R721 B.n192 B.n191 71.676
R722 B.n187 B.n186 71.676
R723 B.n184 B.n183 71.676
R724 B.n179 B.n178 71.676
R725 B.n176 B.n144 71.676
R726 B.n137 B.t7 71.3639
R727 B.t14 B.n511 71.3639
R728 B.t2 B.n101 64.6736
R729 B.n543 B.t5 64.6736
R730 B.n165 B.n164 59.5399
R731 B.n233 B.n158 59.5399
R732 B.n459 B.n70 59.5399
R733 B.n441 B.n76 59.5399
R734 B.n316 B.t1 49.0628
R735 B.n97 B.t0 49.0628
R736 B.t3 B.n551 49.0628
R737 B.n528 B.t4 49.0628
R738 B.n164 B.n163 36.2672
R739 B.n158 B.n157 36.2672
R740 B.n70 B.n69 36.2672
R741 B.n76 B.n75 36.2672
R742 B.n500 B.n499 34.8103
R743 B.n401 B.n400 34.8103
R744 B.n276 B.n143 34.8103
R745 B.n272 B.n271 34.8103
R746 B.t1 B.n113 26.7618
R747 B.n353 B.t0 26.7618
R748 B.n552 B.t3 26.7618
R749 B.t4 B.n29 26.7618
R750 B B.n562 18.0485
R751 B.n334 B.t2 11.151
R752 B.t5 B.n542 11.151
R753 B.n499 B.n498 10.6151
R754 B.n498 B.n59 10.6151
R755 B.n492 B.n59 10.6151
R756 B.n492 B.n491 10.6151
R757 B.n491 B.n490 10.6151
R758 B.n490 B.n61 10.6151
R759 B.n484 B.n61 10.6151
R760 B.n484 B.n483 10.6151
R761 B.n483 B.n482 10.6151
R762 B.n482 B.n63 10.6151
R763 B.n476 B.n63 10.6151
R764 B.n476 B.n475 10.6151
R765 B.n475 B.n474 10.6151
R766 B.n474 B.n65 10.6151
R767 B.n468 B.n65 10.6151
R768 B.n468 B.n467 10.6151
R769 B.n467 B.n466 10.6151
R770 B.n466 B.n67 10.6151
R771 B.n460 B.n67 10.6151
R772 B.n458 B.n457 10.6151
R773 B.n457 B.n71 10.6151
R774 B.n451 B.n71 10.6151
R775 B.n451 B.n450 10.6151
R776 B.n450 B.n449 10.6151
R777 B.n449 B.n73 10.6151
R778 B.n443 B.n73 10.6151
R779 B.n443 B.n442 10.6151
R780 B.n440 B.n77 10.6151
R781 B.n434 B.n77 10.6151
R782 B.n434 B.n433 10.6151
R783 B.n433 B.n432 10.6151
R784 B.n432 B.n79 10.6151
R785 B.n426 B.n79 10.6151
R786 B.n426 B.n425 10.6151
R787 B.n425 B.n424 10.6151
R788 B.n424 B.n81 10.6151
R789 B.n418 B.n81 10.6151
R790 B.n418 B.n417 10.6151
R791 B.n417 B.n416 10.6151
R792 B.n416 B.n83 10.6151
R793 B.n410 B.n83 10.6151
R794 B.n410 B.n409 10.6151
R795 B.n409 B.n408 10.6151
R796 B.n408 B.n85 10.6151
R797 B.n402 B.n85 10.6151
R798 B.n402 B.n401 10.6151
R799 B.n277 B.n276 10.6151
R800 B.n278 B.n277 10.6151
R801 B.n278 B.n134 10.6151
R802 B.n288 B.n134 10.6151
R803 B.n289 B.n288 10.6151
R804 B.n290 B.n289 10.6151
R805 B.n290 B.n127 10.6151
R806 B.n300 B.n127 10.6151
R807 B.n301 B.n300 10.6151
R808 B.n302 B.n301 10.6151
R809 B.n302 B.n119 10.6151
R810 B.n312 B.n119 10.6151
R811 B.n313 B.n312 10.6151
R812 B.n314 B.n313 10.6151
R813 B.n314 B.n111 10.6151
R814 B.n324 B.n111 10.6151
R815 B.n325 B.n324 10.6151
R816 B.n326 B.n325 10.6151
R817 B.n326 B.n103 10.6151
R818 B.n336 B.n103 10.6151
R819 B.n337 B.n336 10.6151
R820 B.n338 B.n337 10.6151
R821 B.n338 B.n94 10.6151
R822 B.n348 B.n94 10.6151
R823 B.n349 B.n348 10.6151
R824 B.n351 B.n349 10.6151
R825 B.n351 B.n350 10.6151
R826 B.n350 B.n87 10.6151
R827 B.n362 B.n87 10.6151
R828 B.n363 B.n362 10.6151
R829 B.n364 B.n363 10.6151
R830 B.n365 B.n364 10.6151
R831 B.n367 B.n365 10.6151
R832 B.n368 B.n367 10.6151
R833 B.n369 B.n368 10.6151
R834 B.n370 B.n369 10.6151
R835 B.n372 B.n370 10.6151
R836 B.n373 B.n372 10.6151
R837 B.n374 B.n373 10.6151
R838 B.n375 B.n374 10.6151
R839 B.n377 B.n375 10.6151
R840 B.n378 B.n377 10.6151
R841 B.n379 B.n378 10.6151
R842 B.n380 B.n379 10.6151
R843 B.n382 B.n380 10.6151
R844 B.n383 B.n382 10.6151
R845 B.n384 B.n383 10.6151
R846 B.n385 B.n384 10.6151
R847 B.n387 B.n385 10.6151
R848 B.n388 B.n387 10.6151
R849 B.n389 B.n388 10.6151
R850 B.n390 B.n389 10.6151
R851 B.n392 B.n390 10.6151
R852 B.n393 B.n392 10.6151
R853 B.n394 B.n393 10.6151
R854 B.n395 B.n394 10.6151
R855 B.n397 B.n395 10.6151
R856 B.n398 B.n397 10.6151
R857 B.n399 B.n398 10.6151
R858 B.n400 B.n399 10.6151
R859 B.n271 B.n270 10.6151
R860 B.n270 B.n147 10.6151
R861 B.n265 B.n147 10.6151
R862 B.n265 B.n264 10.6151
R863 B.n264 B.n149 10.6151
R864 B.n259 B.n149 10.6151
R865 B.n259 B.n258 10.6151
R866 B.n258 B.n257 10.6151
R867 B.n257 B.n151 10.6151
R868 B.n251 B.n151 10.6151
R869 B.n251 B.n250 10.6151
R870 B.n250 B.n249 10.6151
R871 B.n249 B.n153 10.6151
R872 B.n243 B.n153 10.6151
R873 B.n243 B.n242 10.6151
R874 B.n242 B.n241 10.6151
R875 B.n241 B.n155 10.6151
R876 B.n235 B.n155 10.6151
R877 B.n235 B.n234 10.6151
R878 B.n232 B.n159 10.6151
R879 B.n226 B.n159 10.6151
R880 B.n226 B.n225 10.6151
R881 B.n225 B.n224 10.6151
R882 B.n224 B.n161 10.6151
R883 B.n218 B.n161 10.6151
R884 B.n218 B.n217 10.6151
R885 B.n217 B.n216 10.6151
R886 B.n212 B.n211 10.6151
R887 B.n211 B.n167 10.6151
R888 B.n206 B.n167 10.6151
R889 B.n206 B.n205 10.6151
R890 B.n205 B.n204 10.6151
R891 B.n204 B.n169 10.6151
R892 B.n198 B.n169 10.6151
R893 B.n198 B.n197 10.6151
R894 B.n197 B.n196 10.6151
R895 B.n196 B.n171 10.6151
R896 B.n190 B.n171 10.6151
R897 B.n190 B.n189 10.6151
R898 B.n189 B.n188 10.6151
R899 B.n188 B.n173 10.6151
R900 B.n182 B.n173 10.6151
R901 B.n182 B.n181 10.6151
R902 B.n181 B.n180 10.6151
R903 B.n180 B.n175 10.6151
R904 B.n175 B.n143 10.6151
R905 B.n272 B.n139 10.6151
R906 B.n282 B.n139 10.6151
R907 B.n283 B.n282 10.6151
R908 B.n284 B.n283 10.6151
R909 B.n284 B.n131 10.6151
R910 B.n294 B.n131 10.6151
R911 B.n295 B.n294 10.6151
R912 B.n296 B.n295 10.6151
R913 B.n296 B.n123 10.6151
R914 B.n306 B.n123 10.6151
R915 B.n307 B.n306 10.6151
R916 B.n308 B.n307 10.6151
R917 B.n308 B.n115 10.6151
R918 B.n318 B.n115 10.6151
R919 B.n319 B.n318 10.6151
R920 B.n320 B.n319 10.6151
R921 B.n320 B.n107 10.6151
R922 B.n330 B.n107 10.6151
R923 B.n331 B.n330 10.6151
R924 B.n332 B.n331 10.6151
R925 B.n332 B.n99 10.6151
R926 B.n342 B.n99 10.6151
R927 B.n343 B.n342 10.6151
R928 B.n344 B.n343 10.6151
R929 B.n344 B.n91 10.6151
R930 B.n355 B.n91 10.6151
R931 B.n356 B.n355 10.6151
R932 B.n357 B.n356 10.6151
R933 B.n357 B.n0 10.6151
R934 B.n556 B.n1 10.6151
R935 B.n556 B.n555 10.6151
R936 B.n555 B.n554 10.6151
R937 B.n554 B.n10 10.6151
R938 B.n548 B.n10 10.6151
R939 B.n548 B.n547 10.6151
R940 B.n547 B.n546 10.6151
R941 B.n546 B.n17 10.6151
R942 B.n540 B.n17 10.6151
R943 B.n540 B.n539 10.6151
R944 B.n539 B.n538 10.6151
R945 B.n538 B.n24 10.6151
R946 B.n532 B.n24 10.6151
R947 B.n532 B.n531 10.6151
R948 B.n531 B.n530 10.6151
R949 B.n530 B.n31 10.6151
R950 B.n524 B.n31 10.6151
R951 B.n524 B.n523 10.6151
R952 B.n523 B.n522 10.6151
R953 B.n522 B.n38 10.6151
R954 B.n516 B.n38 10.6151
R955 B.n516 B.n515 10.6151
R956 B.n515 B.n514 10.6151
R957 B.n514 B.n45 10.6151
R958 B.n508 B.n45 10.6151
R959 B.n508 B.n507 10.6151
R960 B.n507 B.n506 10.6151
R961 B.n506 B.n52 10.6151
R962 B.n500 B.n52 10.6151
R963 B.n459 B.n458 6.5566
R964 B.n442 B.n441 6.5566
R965 B.n233 B.n232 6.5566
R966 B.n216 B.n165 6.5566
R967 B.n292 B.t7 4.46071
R968 B.n512 B.t14 4.46071
R969 B.n460 B.n459 4.05904
R970 B.n441 B.n440 4.05904
R971 B.n234 B.n233 4.05904
R972 B.n212 B.n165 4.05904
R973 B.n562 B.n0 2.81026
R974 B.n562 B.n1 2.81026
R975 VP.n17 VP.n16 179.895
R976 VP.n32 VP.n31 179.895
R977 VP.n15 VP.n14 179.895
R978 VP.n9 VP.n8 161.3
R979 VP.n10 VP.n5 161.3
R980 VP.n12 VP.n11 161.3
R981 VP.n13 VP.n4 161.3
R982 VP.n30 VP.n0 161.3
R983 VP.n29 VP.n28 161.3
R984 VP.n27 VP.n1 161.3
R985 VP.n26 VP.n25 161.3
R986 VP.n23 VP.n2 161.3
R987 VP.n22 VP.n21 161.3
R988 VP.n20 VP.n3 161.3
R989 VP.n19 VP.n18 161.3
R990 VP.n6 VP.t0 103.346
R991 VP.n17 VP.t4 71.831
R992 VP.n24 VP.t1 71.831
R993 VP.n31 VP.t5 71.831
R994 VP.n14 VP.t2 71.831
R995 VP.n7 VP.t3 71.831
R996 VP.n22 VP.n3 56.5193
R997 VP.n29 VP.n1 56.5193
R998 VP.n12 VP.n5 56.5193
R999 VP.n7 VP.n6 53.731
R1000 VP.n16 VP.n15 38.777
R1001 VP.n18 VP.n3 24.4675
R1002 VP.n23 VP.n22 24.4675
R1003 VP.n25 VP.n1 24.4675
R1004 VP.n30 VP.n29 24.4675
R1005 VP.n13 VP.n12 24.4675
R1006 VP.n8 VP.n5 24.4675
R1007 VP.n9 VP.n6 18.1923
R1008 VP.n24 VP.n23 12.234
R1009 VP.n25 VP.n24 12.234
R1010 VP.n8 VP.n7 12.234
R1011 VP.n18 VP.n17 5.87258
R1012 VP.n31 VP.n30 5.87258
R1013 VP.n14 VP.n13 5.87258
R1014 VP.n10 VP.n9 0.189894
R1015 VP.n11 VP.n10 0.189894
R1016 VP.n11 VP.n4 0.189894
R1017 VP.n15 VP.n4 0.189894
R1018 VP.n19 VP.n16 0.189894
R1019 VP.n20 VP.n19 0.189894
R1020 VP.n21 VP.n20 0.189894
R1021 VP.n21 VP.n2 0.189894
R1022 VP.n26 VP.n2 0.189894
R1023 VP.n27 VP.n26 0.189894
R1024 VP.n28 VP.n27 0.189894
R1025 VP.n28 VP.n0 0.189894
R1026 VP.n32 VP.n0 0.189894
R1027 VP VP.n32 0.0516364
R1028 VTAIL.n98 VTAIL.n80 289.615
R1029 VTAIL.n20 VTAIL.n2 289.615
R1030 VTAIL.n74 VTAIL.n56 289.615
R1031 VTAIL.n48 VTAIL.n30 289.615
R1032 VTAIL.n89 VTAIL.n88 185
R1033 VTAIL.n91 VTAIL.n90 185
R1034 VTAIL.n84 VTAIL.n83 185
R1035 VTAIL.n97 VTAIL.n96 185
R1036 VTAIL.n99 VTAIL.n98 185
R1037 VTAIL.n11 VTAIL.n10 185
R1038 VTAIL.n13 VTAIL.n12 185
R1039 VTAIL.n6 VTAIL.n5 185
R1040 VTAIL.n19 VTAIL.n18 185
R1041 VTAIL.n21 VTAIL.n20 185
R1042 VTAIL.n75 VTAIL.n74 185
R1043 VTAIL.n73 VTAIL.n72 185
R1044 VTAIL.n60 VTAIL.n59 185
R1045 VTAIL.n67 VTAIL.n66 185
R1046 VTAIL.n65 VTAIL.n64 185
R1047 VTAIL.n49 VTAIL.n48 185
R1048 VTAIL.n47 VTAIL.n46 185
R1049 VTAIL.n34 VTAIL.n33 185
R1050 VTAIL.n41 VTAIL.n40 185
R1051 VTAIL.n39 VTAIL.n38 185
R1052 VTAIL.n87 VTAIL.t4 147.714
R1053 VTAIL.n9 VTAIL.t8 147.714
R1054 VTAIL.n63 VTAIL.t9 147.714
R1055 VTAIL.n37 VTAIL.t0 147.714
R1056 VTAIL.n90 VTAIL.n89 104.615
R1057 VTAIL.n90 VTAIL.n83 104.615
R1058 VTAIL.n97 VTAIL.n83 104.615
R1059 VTAIL.n98 VTAIL.n97 104.615
R1060 VTAIL.n12 VTAIL.n11 104.615
R1061 VTAIL.n12 VTAIL.n5 104.615
R1062 VTAIL.n19 VTAIL.n5 104.615
R1063 VTAIL.n20 VTAIL.n19 104.615
R1064 VTAIL.n74 VTAIL.n73 104.615
R1065 VTAIL.n73 VTAIL.n59 104.615
R1066 VTAIL.n66 VTAIL.n59 104.615
R1067 VTAIL.n66 VTAIL.n65 104.615
R1068 VTAIL.n48 VTAIL.n47 104.615
R1069 VTAIL.n47 VTAIL.n33 104.615
R1070 VTAIL.n40 VTAIL.n33 104.615
R1071 VTAIL.n40 VTAIL.n39 104.615
R1072 VTAIL.n55 VTAIL.n54 54.5448
R1073 VTAIL.n29 VTAIL.n28 54.5448
R1074 VTAIL.n1 VTAIL.n0 54.5447
R1075 VTAIL.n27 VTAIL.n26 54.5447
R1076 VTAIL.n89 VTAIL.t4 52.3082
R1077 VTAIL.n11 VTAIL.t8 52.3082
R1078 VTAIL.n65 VTAIL.t9 52.3082
R1079 VTAIL.n39 VTAIL.t0 52.3082
R1080 VTAIL.n103 VTAIL.n102 32.7672
R1081 VTAIL.n25 VTAIL.n24 32.7672
R1082 VTAIL.n79 VTAIL.n78 32.7672
R1083 VTAIL.n53 VTAIL.n52 32.7672
R1084 VTAIL.n29 VTAIL.n27 19.5479
R1085 VTAIL.n103 VTAIL.n79 17.9358
R1086 VTAIL.n88 VTAIL.n87 15.6631
R1087 VTAIL.n10 VTAIL.n9 15.6631
R1088 VTAIL.n64 VTAIL.n63 15.6631
R1089 VTAIL.n38 VTAIL.n37 15.6631
R1090 VTAIL.n91 VTAIL.n86 12.8005
R1091 VTAIL.n13 VTAIL.n8 12.8005
R1092 VTAIL.n67 VTAIL.n62 12.8005
R1093 VTAIL.n41 VTAIL.n36 12.8005
R1094 VTAIL.n92 VTAIL.n84 12.0247
R1095 VTAIL.n14 VTAIL.n6 12.0247
R1096 VTAIL.n68 VTAIL.n60 12.0247
R1097 VTAIL.n42 VTAIL.n34 12.0247
R1098 VTAIL.n96 VTAIL.n95 11.249
R1099 VTAIL.n18 VTAIL.n17 11.249
R1100 VTAIL.n72 VTAIL.n71 11.249
R1101 VTAIL.n46 VTAIL.n45 11.249
R1102 VTAIL.n99 VTAIL.n82 10.4732
R1103 VTAIL.n21 VTAIL.n4 10.4732
R1104 VTAIL.n75 VTAIL.n58 10.4732
R1105 VTAIL.n49 VTAIL.n32 10.4732
R1106 VTAIL.n100 VTAIL.n80 9.69747
R1107 VTAIL.n22 VTAIL.n2 9.69747
R1108 VTAIL.n76 VTAIL.n56 9.69747
R1109 VTAIL.n50 VTAIL.n30 9.69747
R1110 VTAIL.n102 VTAIL.n101 9.45567
R1111 VTAIL.n24 VTAIL.n23 9.45567
R1112 VTAIL.n78 VTAIL.n77 9.45567
R1113 VTAIL.n52 VTAIL.n51 9.45567
R1114 VTAIL.n101 VTAIL.n100 9.3005
R1115 VTAIL.n82 VTAIL.n81 9.3005
R1116 VTAIL.n95 VTAIL.n94 9.3005
R1117 VTAIL.n93 VTAIL.n92 9.3005
R1118 VTAIL.n86 VTAIL.n85 9.3005
R1119 VTAIL.n23 VTAIL.n22 9.3005
R1120 VTAIL.n4 VTAIL.n3 9.3005
R1121 VTAIL.n17 VTAIL.n16 9.3005
R1122 VTAIL.n15 VTAIL.n14 9.3005
R1123 VTAIL.n8 VTAIL.n7 9.3005
R1124 VTAIL.n77 VTAIL.n76 9.3005
R1125 VTAIL.n58 VTAIL.n57 9.3005
R1126 VTAIL.n71 VTAIL.n70 9.3005
R1127 VTAIL.n69 VTAIL.n68 9.3005
R1128 VTAIL.n62 VTAIL.n61 9.3005
R1129 VTAIL.n51 VTAIL.n50 9.3005
R1130 VTAIL.n32 VTAIL.n31 9.3005
R1131 VTAIL.n45 VTAIL.n44 9.3005
R1132 VTAIL.n43 VTAIL.n42 9.3005
R1133 VTAIL.n36 VTAIL.n35 9.3005
R1134 VTAIL.n87 VTAIL.n85 4.39059
R1135 VTAIL.n9 VTAIL.n7 4.39059
R1136 VTAIL.n63 VTAIL.n61 4.39059
R1137 VTAIL.n37 VTAIL.n35 4.39059
R1138 VTAIL.n0 VTAIL.t2 4.31423
R1139 VTAIL.n0 VTAIL.t11 4.31423
R1140 VTAIL.n26 VTAIL.t6 4.31423
R1141 VTAIL.n26 VTAIL.t5 4.31423
R1142 VTAIL.n54 VTAIL.t7 4.31423
R1143 VTAIL.n54 VTAIL.t10 4.31423
R1144 VTAIL.n28 VTAIL.t1 4.31423
R1145 VTAIL.n28 VTAIL.t3 4.31423
R1146 VTAIL.n102 VTAIL.n80 4.26717
R1147 VTAIL.n24 VTAIL.n2 4.26717
R1148 VTAIL.n78 VTAIL.n56 4.26717
R1149 VTAIL.n52 VTAIL.n30 4.26717
R1150 VTAIL.n100 VTAIL.n99 3.49141
R1151 VTAIL.n22 VTAIL.n21 3.49141
R1152 VTAIL.n76 VTAIL.n75 3.49141
R1153 VTAIL.n50 VTAIL.n49 3.49141
R1154 VTAIL.n96 VTAIL.n82 2.71565
R1155 VTAIL.n18 VTAIL.n4 2.71565
R1156 VTAIL.n72 VTAIL.n58 2.71565
R1157 VTAIL.n46 VTAIL.n32 2.71565
R1158 VTAIL.n95 VTAIL.n84 1.93989
R1159 VTAIL.n17 VTAIL.n6 1.93989
R1160 VTAIL.n71 VTAIL.n60 1.93989
R1161 VTAIL.n45 VTAIL.n34 1.93989
R1162 VTAIL.n53 VTAIL.n29 1.61257
R1163 VTAIL.n79 VTAIL.n55 1.61257
R1164 VTAIL.n27 VTAIL.n25 1.61257
R1165 VTAIL.n55 VTAIL.n53 1.27636
R1166 VTAIL.n25 VTAIL.n1 1.27636
R1167 VTAIL.n92 VTAIL.n91 1.16414
R1168 VTAIL.n14 VTAIL.n13 1.16414
R1169 VTAIL.n68 VTAIL.n67 1.16414
R1170 VTAIL.n42 VTAIL.n41 1.16414
R1171 VTAIL VTAIL.n103 1.15136
R1172 VTAIL VTAIL.n1 0.461707
R1173 VTAIL.n88 VTAIL.n86 0.388379
R1174 VTAIL.n10 VTAIL.n8 0.388379
R1175 VTAIL.n64 VTAIL.n62 0.388379
R1176 VTAIL.n38 VTAIL.n36 0.388379
R1177 VTAIL.n93 VTAIL.n85 0.155672
R1178 VTAIL.n94 VTAIL.n93 0.155672
R1179 VTAIL.n94 VTAIL.n81 0.155672
R1180 VTAIL.n101 VTAIL.n81 0.155672
R1181 VTAIL.n15 VTAIL.n7 0.155672
R1182 VTAIL.n16 VTAIL.n15 0.155672
R1183 VTAIL.n16 VTAIL.n3 0.155672
R1184 VTAIL.n23 VTAIL.n3 0.155672
R1185 VTAIL.n77 VTAIL.n57 0.155672
R1186 VTAIL.n70 VTAIL.n57 0.155672
R1187 VTAIL.n70 VTAIL.n69 0.155672
R1188 VTAIL.n69 VTAIL.n61 0.155672
R1189 VTAIL.n51 VTAIL.n31 0.155672
R1190 VTAIL.n44 VTAIL.n31 0.155672
R1191 VTAIL.n44 VTAIL.n43 0.155672
R1192 VTAIL.n43 VTAIL.n35 0.155672
R1193 VDD1.n18 VDD1.n0 289.615
R1194 VDD1.n41 VDD1.n23 289.615
R1195 VDD1.n19 VDD1.n18 185
R1196 VDD1.n17 VDD1.n16 185
R1197 VDD1.n4 VDD1.n3 185
R1198 VDD1.n11 VDD1.n10 185
R1199 VDD1.n9 VDD1.n8 185
R1200 VDD1.n32 VDD1.n31 185
R1201 VDD1.n34 VDD1.n33 185
R1202 VDD1.n27 VDD1.n26 185
R1203 VDD1.n40 VDD1.n39 185
R1204 VDD1.n42 VDD1.n41 185
R1205 VDD1.n7 VDD1.t5 147.714
R1206 VDD1.n30 VDD1.t1 147.714
R1207 VDD1.n18 VDD1.n17 104.615
R1208 VDD1.n17 VDD1.n3 104.615
R1209 VDD1.n10 VDD1.n3 104.615
R1210 VDD1.n10 VDD1.n9 104.615
R1211 VDD1.n33 VDD1.n32 104.615
R1212 VDD1.n33 VDD1.n26 104.615
R1213 VDD1.n40 VDD1.n26 104.615
R1214 VDD1.n41 VDD1.n40 104.615
R1215 VDD1.n47 VDD1.n46 71.5711
R1216 VDD1.n49 VDD1.n48 71.2235
R1217 VDD1.n9 VDD1.t5 52.3082
R1218 VDD1.n32 VDD1.t1 52.3082
R1219 VDD1 VDD1.n22 50.7132
R1220 VDD1.n47 VDD1.n45 50.5997
R1221 VDD1.n49 VDD1.n47 34.3005
R1222 VDD1.n8 VDD1.n7 15.6631
R1223 VDD1.n31 VDD1.n30 15.6631
R1224 VDD1.n11 VDD1.n6 12.8005
R1225 VDD1.n34 VDD1.n29 12.8005
R1226 VDD1.n12 VDD1.n4 12.0247
R1227 VDD1.n35 VDD1.n27 12.0247
R1228 VDD1.n16 VDD1.n15 11.249
R1229 VDD1.n39 VDD1.n38 11.249
R1230 VDD1.n19 VDD1.n2 10.4732
R1231 VDD1.n42 VDD1.n25 10.4732
R1232 VDD1.n20 VDD1.n0 9.69747
R1233 VDD1.n43 VDD1.n23 9.69747
R1234 VDD1.n22 VDD1.n21 9.45567
R1235 VDD1.n45 VDD1.n44 9.45567
R1236 VDD1.n21 VDD1.n20 9.3005
R1237 VDD1.n2 VDD1.n1 9.3005
R1238 VDD1.n15 VDD1.n14 9.3005
R1239 VDD1.n13 VDD1.n12 9.3005
R1240 VDD1.n6 VDD1.n5 9.3005
R1241 VDD1.n44 VDD1.n43 9.3005
R1242 VDD1.n25 VDD1.n24 9.3005
R1243 VDD1.n38 VDD1.n37 9.3005
R1244 VDD1.n36 VDD1.n35 9.3005
R1245 VDD1.n29 VDD1.n28 9.3005
R1246 VDD1.n7 VDD1.n5 4.39059
R1247 VDD1.n30 VDD1.n28 4.39059
R1248 VDD1.n48 VDD1.t2 4.31423
R1249 VDD1.n48 VDD1.t3 4.31423
R1250 VDD1.n46 VDD1.t4 4.31423
R1251 VDD1.n46 VDD1.t0 4.31423
R1252 VDD1.n22 VDD1.n0 4.26717
R1253 VDD1.n45 VDD1.n23 4.26717
R1254 VDD1.n20 VDD1.n19 3.49141
R1255 VDD1.n43 VDD1.n42 3.49141
R1256 VDD1.n16 VDD1.n2 2.71565
R1257 VDD1.n39 VDD1.n25 2.71565
R1258 VDD1.n15 VDD1.n4 1.93989
R1259 VDD1.n38 VDD1.n27 1.93989
R1260 VDD1.n12 VDD1.n11 1.16414
R1261 VDD1.n35 VDD1.n34 1.16414
R1262 VDD1.n8 VDD1.n6 0.388379
R1263 VDD1.n31 VDD1.n29 0.388379
R1264 VDD1 VDD1.n49 0.345328
R1265 VDD1.n21 VDD1.n1 0.155672
R1266 VDD1.n14 VDD1.n1 0.155672
R1267 VDD1.n14 VDD1.n13 0.155672
R1268 VDD1.n13 VDD1.n5 0.155672
R1269 VDD1.n36 VDD1.n28 0.155672
R1270 VDD1.n37 VDD1.n36 0.155672
R1271 VDD1.n37 VDD1.n24 0.155672
R1272 VDD1.n44 VDD1.n24 0.155672
R1273 VN.n11 VN.n10 179.895
R1274 VN.n23 VN.n22 179.895
R1275 VN.n21 VN.n12 161.3
R1276 VN.n20 VN.n19 161.3
R1277 VN.n18 VN.n13 161.3
R1278 VN.n17 VN.n16 161.3
R1279 VN.n9 VN.n0 161.3
R1280 VN.n8 VN.n7 161.3
R1281 VN.n6 VN.n1 161.3
R1282 VN.n5 VN.n4 161.3
R1283 VN.n2 VN.t2 103.346
R1284 VN.n14 VN.t3 103.346
R1285 VN.n3 VN.t1 71.831
R1286 VN.n10 VN.t0 71.831
R1287 VN.n15 VN.t5 71.831
R1288 VN.n22 VN.t4 71.831
R1289 VN.n8 VN.n1 56.5193
R1290 VN.n20 VN.n13 56.5193
R1291 VN.n3 VN.n2 53.731
R1292 VN.n15 VN.n14 53.731
R1293 VN VN.n23 39.1577
R1294 VN.n4 VN.n1 24.4675
R1295 VN.n9 VN.n8 24.4675
R1296 VN.n16 VN.n13 24.4675
R1297 VN.n21 VN.n20 24.4675
R1298 VN.n17 VN.n14 18.1923
R1299 VN.n5 VN.n2 18.1923
R1300 VN.n4 VN.n3 12.234
R1301 VN.n16 VN.n15 12.234
R1302 VN.n10 VN.n9 5.87258
R1303 VN.n22 VN.n21 5.87258
R1304 VN.n23 VN.n12 0.189894
R1305 VN.n19 VN.n12 0.189894
R1306 VN.n19 VN.n18 0.189894
R1307 VN.n18 VN.n17 0.189894
R1308 VN.n6 VN.n5 0.189894
R1309 VN.n7 VN.n6 0.189894
R1310 VN.n7 VN.n0 0.189894
R1311 VN.n11 VN.n0 0.189894
R1312 VN VN.n11 0.0516364
R1313 VDD2.n43 VDD2.n25 289.615
R1314 VDD2.n18 VDD2.n0 289.615
R1315 VDD2.n44 VDD2.n43 185
R1316 VDD2.n42 VDD2.n41 185
R1317 VDD2.n29 VDD2.n28 185
R1318 VDD2.n36 VDD2.n35 185
R1319 VDD2.n34 VDD2.n33 185
R1320 VDD2.n9 VDD2.n8 185
R1321 VDD2.n11 VDD2.n10 185
R1322 VDD2.n4 VDD2.n3 185
R1323 VDD2.n17 VDD2.n16 185
R1324 VDD2.n19 VDD2.n18 185
R1325 VDD2.n32 VDD2.t1 147.714
R1326 VDD2.n7 VDD2.t3 147.714
R1327 VDD2.n43 VDD2.n42 104.615
R1328 VDD2.n42 VDD2.n28 104.615
R1329 VDD2.n35 VDD2.n28 104.615
R1330 VDD2.n35 VDD2.n34 104.615
R1331 VDD2.n10 VDD2.n9 104.615
R1332 VDD2.n10 VDD2.n3 104.615
R1333 VDD2.n17 VDD2.n3 104.615
R1334 VDD2.n18 VDD2.n17 104.615
R1335 VDD2.n24 VDD2.n23 71.5711
R1336 VDD2 VDD2.n49 71.5683
R1337 VDD2.n34 VDD2.t1 52.3082
R1338 VDD2.n9 VDD2.t3 52.3082
R1339 VDD2.n24 VDD2.n22 50.5997
R1340 VDD2.n48 VDD2.n47 49.446
R1341 VDD2.n48 VDD2.n24 32.9114
R1342 VDD2.n33 VDD2.n32 15.6631
R1343 VDD2.n8 VDD2.n7 15.6631
R1344 VDD2.n36 VDD2.n31 12.8005
R1345 VDD2.n11 VDD2.n6 12.8005
R1346 VDD2.n37 VDD2.n29 12.0247
R1347 VDD2.n12 VDD2.n4 12.0247
R1348 VDD2.n41 VDD2.n40 11.249
R1349 VDD2.n16 VDD2.n15 11.249
R1350 VDD2.n44 VDD2.n27 10.4732
R1351 VDD2.n19 VDD2.n2 10.4732
R1352 VDD2.n45 VDD2.n25 9.69747
R1353 VDD2.n20 VDD2.n0 9.69747
R1354 VDD2.n47 VDD2.n46 9.45567
R1355 VDD2.n22 VDD2.n21 9.45567
R1356 VDD2.n46 VDD2.n45 9.3005
R1357 VDD2.n27 VDD2.n26 9.3005
R1358 VDD2.n40 VDD2.n39 9.3005
R1359 VDD2.n38 VDD2.n37 9.3005
R1360 VDD2.n31 VDD2.n30 9.3005
R1361 VDD2.n21 VDD2.n20 9.3005
R1362 VDD2.n2 VDD2.n1 9.3005
R1363 VDD2.n15 VDD2.n14 9.3005
R1364 VDD2.n13 VDD2.n12 9.3005
R1365 VDD2.n6 VDD2.n5 9.3005
R1366 VDD2.n32 VDD2.n30 4.39059
R1367 VDD2.n7 VDD2.n5 4.39059
R1368 VDD2.n49 VDD2.t0 4.31423
R1369 VDD2.n49 VDD2.t2 4.31423
R1370 VDD2.n23 VDD2.t4 4.31423
R1371 VDD2.n23 VDD2.t5 4.31423
R1372 VDD2.n47 VDD2.n25 4.26717
R1373 VDD2.n22 VDD2.n0 4.26717
R1374 VDD2.n45 VDD2.n44 3.49141
R1375 VDD2.n20 VDD2.n19 3.49141
R1376 VDD2.n41 VDD2.n27 2.71565
R1377 VDD2.n16 VDD2.n2 2.71565
R1378 VDD2.n40 VDD2.n29 1.93989
R1379 VDD2.n15 VDD2.n4 1.93989
R1380 VDD2 VDD2.n48 1.26774
R1381 VDD2.n37 VDD2.n36 1.16414
R1382 VDD2.n12 VDD2.n11 1.16414
R1383 VDD2.n33 VDD2.n31 0.388379
R1384 VDD2.n8 VDD2.n6 0.388379
R1385 VDD2.n46 VDD2.n26 0.155672
R1386 VDD2.n39 VDD2.n26 0.155672
R1387 VDD2.n39 VDD2.n38 0.155672
R1388 VDD2.n38 VDD2.n30 0.155672
R1389 VDD2.n13 VDD2.n5 0.155672
R1390 VDD2.n14 VDD2.n13 0.155672
R1391 VDD2.n14 VDD2.n1 0.155672
R1392 VDD2.n21 VDD2.n1 0.155672
C0 VTAIL VP 2.82659f
C1 VN VP 4.53149f
C2 VDD1 VDD2 1.02136f
C3 VTAIL VN 2.81237f
C4 VDD1 VP 2.70587f
C5 VDD2 VP 0.372153f
C6 VDD1 VTAIL 4.60557f
C7 VDD1 VN 0.153328f
C8 VDD2 VTAIL 4.65038f
C9 VDD2 VN 2.4893f
C10 VDD2 B 3.815454f
C11 VDD1 B 3.887883f
C12 VTAIL B 3.983942f
C13 VN B 9.076851f
C14 VP B 7.648355f
C15 VDD2.n0 B 0.030691f
C16 VDD2.n1 B 0.022372f
C17 VDD2.n2 B 0.012022f
C18 VDD2.n3 B 0.028415f
C19 VDD2.n4 B 0.012729f
C20 VDD2.n5 B 0.386633f
C21 VDD2.n6 B 0.012022f
C22 VDD2.t3 B 0.046604f
C23 VDD2.n7 B 0.088559f
C24 VDD2.n8 B 0.016769f
C25 VDD2.n9 B 0.021311f
C26 VDD2.n10 B 0.028415f
C27 VDD2.n11 B 0.012729f
C28 VDD2.n12 B 0.012022f
C29 VDD2.n13 B 0.022372f
C30 VDD2.n14 B 0.022372f
C31 VDD2.n15 B 0.012022f
C32 VDD2.n16 B 0.012729f
C33 VDD2.n17 B 0.028415f
C34 VDD2.n18 B 0.060179f
C35 VDD2.n19 B 0.012729f
C36 VDD2.n20 B 0.012022f
C37 VDD2.n21 B 0.052628f
C38 VDD2.n22 B 0.051904f
C39 VDD2.t4 B 0.081146f
C40 VDD2.t5 B 0.081146f
C41 VDD2.n23 B 0.654089f
C42 VDD2.n24 B 1.58348f
C43 VDD2.n25 B 0.030691f
C44 VDD2.n26 B 0.022372f
C45 VDD2.n27 B 0.012022f
C46 VDD2.n28 B 0.028415f
C47 VDD2.n29 B 0.012729f
C48 VDD2.n30 B 0.386633f
C49 VDD2.n31 B 0.012022f
C50 VDD2.t1 B 0.046604f
C51 VDD2.n32 B 0.088559f
C52 VDD2.n33 B 0.016769f
C53 VDD2.n34 B 0.021311f
C54 VDD2.n35 B 0.028415f
C55 VDD2.n36 B 0.012729f
C56 VDD2.n37 B 0.012022f
C57 VDD2.n38 B 0.022372f
C58 VDD2.n39 B 0.022372f
C59 VDD2.n40 B 0.012022f
C60 VDD2.n41 B 0.012729f
C61 VDD2.n42 B 0.028415f
C62 VDD2.n43 B 0.060179f
C63 VDD2.n44 B 0.012729f
C64 VDD2.n45 B 0.012022f
C65 VDD2.n46 B 0.052628f
C66 VDD2.n47 B 0.049003f
C67 VDD2.n48 B 1.50809f
C68 VDD2.t0 B 0.081146f
C69 VDD2.t2 B 0.081146f
C70 VDD2.n49 B 0.654068f
C71 VN.n0 B 0.035173f
C72 VN.t0 B 0.64617f
C73 VN.n1 B 0.04498f
C74 VN.t2 B 0.768908f
C75 VN.n2 B 0.340061f
C76 VN.t1 B 0.64617f
C77 VN.n3 B 0.331214f
C78 VN.n4 B 0.049372f
C79 VN.n5 B 0.221285f
C80 VN.n6 B 0.035173f
C81 VN.n7 B 0.035173f
C82 VN.n8 B 0.057721f
C83 VN.n9 B 0.040957f
C84 VN.n10 B 0.332686f
C85 VN.n11 B 0.035105f
C86 VN.n12 B 0.035173f
C87 VN.t4 B 0.64617f
C88 VN.n13 B 0.04498f
C89 VN.t3 B 0.768908f
C90 VN.n14 B 0.340061f
C91 VN.t5 B 0.64617f
C92 VN.n15 B 0.331214f
C93 VN.n16 B 0.049372f
C94 VN.n17 B 0.221285f
C95 VN.n18 B 0.035173f
C96 VN.n19 B 0.035173f
C97 VN.n20 B 0.057721f
C98 VN.n21 B 0.040957f
C99 VN.n22 B 0.332686f
C100 VN.n23 B 1.29714f
C101 VDD1.n0 B 0.030764f
C102 VDD1.n1 B 0.022425f
C103 VDD1.n2 B 0.01205f
C104 VDD1.n3 B 0.028483f
C105 VDD1.n4 B 0.012759f
C106 VDD1.n5 B 0.387555f
C107 VDD1.n6 B 0.01205f
C108 VDD1.t5 B 0.046715f
C109 VDD1.n7 B 0.08877f
C110 VDD1.n8 B 0.016809f
C111 VDD1.n9 B 0.021362f
C112 VDD1.n10 B 0.028483f
C113 VDD1.n11 B 0.012759f
C114 VDD1.n12 B 0.01205f
C115 VDD1.n13 B 0.022425f
C116 VDD1.n14 B 0.022425f
C117 VDD1.n15 B 0.01205f
C118 VDD1.n16 B 0.012759f
C119 VDD1.n17 B 0.028483f
C120 VDD1.n18 B 0.060322f
C121 VDD1.n19 B 0.012759f
C122 VDD1.n20 B 0.01205f
C123 VDD1.n21 B 0.052754f
C124 VDD1.n22 B 0.0525f
C125 VDD1.n23 B 0.030764f
C126 VDD1.n24 B 0.022425f
C127 VDD1.n25 B 0.01205f
C128 VDD1.n26 B 0.028483f
C129 VDD1.n27 B 0.012759f
C130 VDD1.n28 B 0.387555f
C131 VDD1.n29 B 0.01205f
C132 VDD1.t1 B 0.046715f
C133 VDD1.n30 B 0.08877f
C134 VDD1.n31 B 0.016809f
C135 VDD1.n32 B 0.021362f
C136 VDD1.n33 B 0.028483f
C137 VDD1.n34 B 0.012759f
C138 VDD1.n35 B 0.01205f
C139 VDD1.n36 B 0.022425f
C140 VDD1.n37 B 0.022425f
C141 VDD1.n38 B 0.01205f
C142 VDD1.n39 B 0.012759f
C143 VDD1.n40 B 0.028483f
C144 VDD1.n41 B 0.060322f
C145 VDD1.n42 B 0.012759f
C146 VDD1.n43 B 0.01205f
C147 VDD1.n44 B 0.052754f
C148 VDD1.n45 B 0.052028f
C149 VDD1.t4 B 0.08134f
C150 VDD1.t0 B 0.08134f
C151 VDD1.n46 B 0.655649f
C152 VDD1.n47 B 1.66964f
C153 VDD1.t2 B 0.08134f
C154 VDD1.t3 B 0.08134f
C155 VDD1.n48 B 0.65405f
C156 VDD1.n49 B 1.70427f
C157 VTAIL.t2 B 0.0985f
C158 VTAIL.t11 B 0.0985f
C159 VTAIL.n0 B 0.728087f
C160 VTAIL.n1 B 0.393349f
C161 VTAIL.n2 B 0.037255f
C162 VTAIL.n3 B 0.027156f
C163 VTAIL.n4 B 0.014593f
C164 VTAIL.n5 B 0.034492f
C165 VTAIL.n6 B 0.015451f
C166 VTAIL.n7 B 0.469319f
C167 VTAIL.n8 B 0.014593f
C168 VTAIL.t8 B 0.05657f
C169 VTAIL.n9 B 0.107498f
C170 VTAIL.n10 B 0.020355f
C171 VTAIL.n11 B 0.025869f
C172 VTAIL.n12 B 0.034492f
C173 VTAIL.n13 B 0.015451f
C174 VTAIL.n14 B 0.014593f
C175 VTAIL.n15 B 0.027156f
C176 VTAIL.n16 B 0.027156f
C177 VTAIL.n17 B 0.014593f
C178 VTAIL.n18 B 0.015451f
C179 VTAIL.n19 B 0.034492f
C180 VTAIL.n20 B 0.073049f
C181 VTAIL.n21 B 0.015451f
C182 VTAIL.n22 B 0.014593f
C183 VTAIL.n23 B 0.063884f
C184 VTAIL.n24 B 0.040741f
C185 VTAIL.n25 B 0.276527f
C186 VTAIL.t6 B 0.0985f
C187 VTAIL.t5 B 0.0985f
C188 VTAIL.n26 B 0.728087f
C189 VTAIL.n27 B 1.37967f
C190 VTAIL.t1 B 0.0985f
C191 VTAIL.t3 B 0.0985f
C192 VTAIL.n28 B 0.728092f
C193 VTAIL.n29 B 1.37966f
C194 VTAIL.n30 B 0.037255f
C195 VTAIL.n31 B 0.027156f
C196 VTAIL.n32 B 0.014593f
C197 VTAIL.n33 B 0.034492f
C198 VTAIL.n34 B 0.015451f
C199 VTAIL.n35 B 0.469319f
C200 VTAIL.n36 B 0.014593f
C201 VTAIL.t0 B 0.05657f
C202 VTAIL.n37 B 0.107498f
C203 VTAIL.n38 B 0.020355f
C204 VTAIL.n39 B 0.025869f
C205 VTAIL.n40 B 0.034492f
C206 VTAIL.n41 B 0.015451f
C207 VTAIL.n42 B 0.014593f
C208 VTAIL.n43 B 0.027156f
C209 VTAIL.n44 B 0.027156f
C210 VTAIL.n45 B 0.014593f
C211 VTAIL.n46 B 0.015451f
C212 VTAIL.n47 B 0.034492f
C213 VTAIL.n48 B 0.073049f
C214 VTAIL.n49 B 0.015451f
C215 VTAIL.n50 B 0.014593f
C216 VTAIL.n51 B 0.063884f
C217 VTAIL.n52 B 0.040741f
C218 VTAIL.n53 B 0.276527f
C219 VTAIL.t7 B 0.0985f
C220 VTAIL.t10 B 0.0985f
C221 VTAIL.n54 B 0.728092f
C222 VTAIL.n55 B 0.494048f
C223 VTAIL.n56 B 0.037255f
C224 VTAIL.n57 B 0.027156f
C225 VTAIL.n58 B 0.014593f
C226 VTAIL.n59 B 0.034492f
C227 VTAIL.n60 B 0.015451f
C228 VTAIL.n61 B 0.469319f
C229 VTAIL.n62 B 0.014593f
C230 VTAIL.t9 B 0.05657f
C231 VTAIL.n63 B 0.107498f
C232 VTAIL.n64 B 0.020355f
C233 VTAIL.n65 B 0.025869f
C234 VTAIL.n66 B 0.034492f
C235 VTAIL.n67 B 0.015451f
C236 VTAIL.n68 B 0.014593f
C237 VTAIL.n69 B 0.027156f
C238 VTAIL.n70 B 0.027156f
C239 VTAIL.n71 B 0.014593f
C240 VTAIL.n72 B 0.015451f
C241 VTAIL.n73 B 0.034492f
C242 VTAIL.n74 B 0.073049f
C243 VTAIL.n75 B 0.015451f
C244 VTAIL.n76 B 0.014593f
C245 VTAIL.n77 B 0.063884f
C246 VTAIL.n78 B 0.040741f
C247 VTAIL.n79 B 1.02108f
C248 VTAIL.n80 B 0.037255f
C249 VTAIL.n81 B 0.027156f
C250 VTAIL.n82 B 0.014593f
C251 VTAIL.n83 B 0.034492f
C252 VTAIL.n84 B 0.015451f
C253 VTAIL.n85 B 0.469319f
C254 VTAIL.n86 B 0.014593f
C255 VTAIL.t4 B 0.05657f
C256 VTAIL.n87 B 0.107498f
C257 VTAIL.n88 B 0.020355f
C258 VTAIL.n89 B 0.025869f
C259 VTAIL.n90 B 0.034492f
C260 VTAIL.n91 B 0.015451f
C261 VTAIL.n92 B 0.014593f
C262 VTAIL.n93 B 0.027156f
C263 VTAIL.n94 B 0.027156f
C264 VTAIL.n95 B 0.014593f
C265 VTAIL.n96 B 0.015451f
C266 VTAIL.n97 B 0.034492f
C267 VTAIL.n98 B 0.073049f
C268 VTAIL.n99 B 0.015451f
C269 VTAIL.n100 B 0.014593f
C270 VTAIL.n101 B 0.063884f
C271 VTAIL.n102 B 0.040741f
C272 VTAIL.n103 B 0.98072f
C273 VP.n0 B 0.036073f
C274 VP.t5 B 0.662701f
C275 VP.n1 B 0.04613f
C276 VP.n2 B 0.036073f
C277 VP.t1 B 0.662701f
C278 VP.n3 B 0.059198f
C279 VP.n4 B 0.036073f
C280 VP.t2 B 0.662701f
C281 VP.n5 B 0.04613f
C282 VP.t0 B 0.788579f
C283 VP.n6 B 0.34876f
C284 VP.t3 B 0.662701f
C285 VP.n7 B 0.339687f
C286 VP.n8 B 0.050635f
C287 VP.n9 B 0.226946f
C288 VP.n10 B 0.036073f
C289 VP.n11 B 0.036073f
C290 VP.n12 B 0.059198f
C291 VP.n13 B 0.042005f
C292 VP.n14 B 0.341197f
C293 VP.n15 B 1.30652f
C294 VP.n16 B 1.33996f
C295 VP.t4 B 0.662701f
C296 VP.n17 B 0.341197f
C297 VP.n18 B 0.042005f
C298 VP.n19 B 0.036073f
C299 VP.n20 B 0.036073f
C300 VP.n21 B 0.036073f
C301 VP.n22 B 0.04613f
C302 VP.n23 B 0.050635f
C303 VP.n24 B 0.271391f
C304 VP.n25 B 0.050635f
C305 VP.n26 B 0.036073f
C306 VP.n27 B 0.036073f
C307 VP.n28 B 0.036073f
C308 VP.n29 B 0.059198f
C309 VP.n30 B 0.042005f
C310 VP.n31 B 0.341197f
C311 VP.n32 B 0.036003f
.ends

