* NGSPICE file created from diff_pair_sample_0884.ext - technology: sky130A

.subckt diff_pair_sample_0884 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t3 VN.t0 VTAIL.t7 w_n2782_n2174# sky130_fd_pr__pfet_01v8 ad=0.99495 pd=6.36 as=2.3517 ps=12.84 w=6.03 l=2.69
X1 VTAIL.t6 VN.t1 VDD2.t2 w_n2782_n2174# sky130_fd_pr__pfet_01v8 ad=2.3517 pd=12.84 as=0.99495 ps=6.36 w=6.03 l=2.69
X2 VDD1.t3 VP.t0 VTAIL.t3 w_n2782_n2174# sky130_fd_pr__pfet_01v8 ad=0.99495 pd=6.36 as=2.3517 ps=12.84 w=6.03 l=2.69
X3 VTAIL.t5 VN.t2 VDD2.t1 w_n2782_n2174# sky130_fd_pr__pfet_01v8 ad=2.3517 pd=12.84 as=0.99495 ps=6.36 w=6.03 l=2.69
X4 VDD2.t0 VN.t3 VTAIL.t4 w_n2782_n2174# sky130_fd_pr__pfet_01v8 ad=0.99495 pd=6.36 as=2.3517 ps=12.84 w=6.03 l=2.69
X5 VDD1.t2 VP.t1 VTAIL.t0 w_n2782_n2174# sky130_fd_pr__pfet_01v8 ad=0.99495 pd=6.36 as=2.3517 ps=12.84 w=6.03 l=2.69
X6 VTAIL.t2 VP.t2 VDD1.t1 w_n2782_n2174# sky130_fd_pr__pfet_01v8 ad=2.3517 pd=12.84 as=0.99495 ps=6.36 w=6.03 l=2.69
X7 B.t11 B.t9 B.t10 w_n2782_n2174# sky130_fd_pr__pfet_01v8 ad=2.3517 pd=12.84 as=0 ps=0 w=6.03 l=2.69
X8 VTAIL.t1 VP.t3 VDD1.t0 w_n2782_n2174# sky130_fd_pr__pfet_01v8 ad=2.3517 pd=12.84 as=0.99495 ps=6.36 w=6.03 l=2.69
X9 B.t8 B.t6 B.t7 w_n2782_n2174# sky130_fd_pr__pfet_01v8 ad=2.3517 pd=12.84 as=0 ps=0 w=6.03 l=2.69
X10 B.t5 B.t3 B.t4 w_n2782_n2174# sky130_fd_pr__pfet_01v8 ad=2.3517 pd=12.84 as=0 ps=0 w=6.03 l=2.69
X11 B.t2 B.t0 B.t1 w_n2782_n2174# sky130_fd_pr__pfet_01v8 ad=2.3517 pd=12.84 as=0 ps=0 w=6.03 l=2.69
R0 VN.n0 VN.t1 87.9394
R1 VN.n1 VN.t3 87.9394
R2 VN.n0 VN.t0 87.0709
R3 VN.n1 VN.t2 87.0709
R4 VN VN.n1 45.9062
R5 VN VN.n0 3.66761
R6 VTAIL.n250 VTAIL.n224 756.745
R7 VTAIL.n26 VTAIL.n0 756.745
R8 VTAIL.n58 VTAIL.n32 756.745
R9 VTAIL.n90 VTAIL.n64 756.745
R10 VTAIL.n218 VTAIL.n192 756.745
R11 VTAIL.n186 VTAIL.n160 756.745
R12 VTAIL.n154 VTAIL.n128 756.745
R13 VTAIL.n122 VTAIL.n96 756.745
R14 VTAIL.n235 VTAIL.n234 585
R15 VTAIL.n232 VTAIL.n231 585
R16 VTAIL.n241 VTAIL.n240 585
R17 VTAIL.n243 VTAIL.n242 585
R18 VTAIL.n228 VTAIL.n227 585
R19 VTAIL.n249 VTAIL.n248 585
R20 VTAIL.n251 VTAIL.n250 585
R21 VTAIL.n11 VTAIL.n10 585
R22 VTAIL.n8 VTAIL.n7 585
R23 VTAIL.n17 VTAIL.n16 585
R24 VTAIL.n19 VTAIL.n18 585
R25 VTAIL.n4 VTAIL.n3 585
R26 VTAIL.n25 VTAIL.n24 585
R27 VTAIL.n27 VTAIL.n26 585
R28 VTAIL.n43 VTAIL.n42 585
R29 VTAIL.n40 VTAIL.n39 585
R30 VTAIL.n49 VTAIL.n48 585
R31 VTAIL.n51 VTAIL.n50 585
R32 VTAIL.n36 VTAIL.n35 585
R33 VTAIL.n57 VTAIL.n56 585
R34 VTAIL.n59 VTAIL.n58 585
R35 VTAIL.n75 VTAIL.n74 585
R36 VTAIL.n72 VTAIL.n71 585
R37 VTAIL.n81 VTAIL.n80 585
R38 VTAIL.n83 VTAIL.n82 585
R39 VTAIL.n68 VTAIL.n67 585
R40 VTAIL.n89 VTAIL.n88 585
R41 VTAIL.n91 VTAIL.n90 585
R42 VTAIL.n219 VTAIL.n218 585
R43 VTAIL.n217 VTAIL.n216 585
R44 VTAIL.n196 VTAIL.n195 585
R45 VTAIL.n211 VTAIL.n210 585
R46 VTAIL.n209 VTAIL.n208 585
R47 VTAIL.n200 VTAIL.n199 585
R48 VTAIL.n203 VTAIL.n202 585
R49 VTAIL.n187 VTAIL.n186 585
R50 VTAIL.n185 VTAIL.n184 585
R51 VTAIL.n164 VTAIL.n163 585
R52 VTAIL.n179 VTAIL.n178 585
R53 VTAIL.n177 VTAIL.n176 585
R54 VTAIL.n168 VTAIL.n167 585
R55 VTAIL.n171 VTAIL.n170 585
R56 VTAIL.n155 VTAIL.n154 585
R57 VTAIL.n153 VTAIL.n152 585
R58 VTAIL.n132 VTAIL.n131 585
R59 VTAIL.n147 VTAIL.n146 585
R60 VTAIL.n145 VTAIL.n144 585
R61 VTAIL.n136 VTAIL.n135 585
R62 VTAIL.n139 VTAIL.n138 585
R63 VTAIL.n123 VTAIL.n122 585
R64 VTAIL.n121 VTAIL.n120 585
R65 VTAIL.n100 VTAIL.n99 585
R66 VTAIL.n115 VTAIL.n114 585
R67 VTAIL.n113 VTAIL.n112 585
R68 VTAIL.n104 VTAIL.n103 585
R69 VTAIL.n107 VTAIL.n106 585
R70 VTAIL.t7 VTAIL.n233 327.601
R71 VTAIL.t6 VTAIL.n9 327.601
R72 VTAIL.t0 VTAIL.n41 327.601
R73 VTAIL.t1 VTAIL.n73 327.601
R74 VTAIL.t3 VTAIL.n201 327.601
R75 VTAIL.t2 VTAIL.n169 327.601
R76 VTAIL.t4 VTAIL.n137 327.601
R77 VTAIL.t5 VTAIL.n105 327.601
R78 VTAIL.n234 VTAIL.n231 171.744
R79 VTAIL.n241 VTAIL.n231 171.744
R80 VTAIL.n242 VTAIL.n241 171.744
R81 VTAIL.n242 VTAIL.n227 171.744
R82 VTAIL.n249 VTAIL.n227 171.744
R83 VTAIL.n250 VTAIL.n249 171.744
R84 VTAIL.n10 VTAIL.n7 171.744
R85 VTAIL.n17 VTAIL.n7 171.744
R86 VTAIL.n18 VTAIL.n17 171.744
R87 VTAIL.n18 VTAIL.n3 171.744
R88 VTAIL.n25 VTAIL.n3 171.744
R89 VTAIL.n26 VTAIL.n25 171.744
R90 VTAIL.n42 VTAIL.n39 171.744
R91 VTAIL.n49 VTAIL.n39 171.744
R92 VTAIL.n50 VTAIL.n49 171.744
R93 VTAIL.n50 VTAIL.n35 171.744
R94 VTAIL.n57 VTAIL.n35 171.744
R95 VTAIL.n58 VTAIL.n57 171.744
R96 VTAIL.n74 VTAIL.n71 171.744
R97 VTAIL.n81 VTAIL.n71 171.744
R98 VTAIL.n82 VTAIL.n81 171.744
R99 VTAIL.n82 VTAIL.n67 171.744
R100 VTAIL.n89 VTAIL.n67 171.744
R101 VTAIL.n90 VTAIL.n89 171.744
R102 VTAIL.n218 VTAIL.n217 171.744
R103 VTAIL.n217 VTAIL.n195 171.744
R104 VTAIL.n210 VTAIL.n195 171.744
R105 VTAIL.n210 VTAIL.n209 171.744
R106 VTAIL.n209 VTAIL.n199 171.744
R107 VTAIL.n202 VTAIL.n199 171.744
R108 VTAIL.n186 VTAIL.n185 171.744
R109 VTAIL.n185 VTAIL.n163 171.744
R110 VTAIL.n178 VTAIL.n163 171.744
R111 VTAIL.n178 VTAIL.n177 171.744
R112 VTAIL.n177 VTAIL.n167 171.744
R113 VTAIL.n170 VTAIL.n167 171.744
R114 VTAIL.n154 VTAIL.n153 171.744
R115 VTAIL.n153 VTAIL.n131 171.744
R116 VTAIL.n146 VTAIL.n131 171.744
R117 VTAIL.n146 VTAIL.n145 171.744
R118 VTAIL.n145 VTAIL.n135 171.744
R119 VTAIL.n138 VTAIL.n135 171.744
R120 VTAIL.n122 VTAIL.n121 171.744
R121 VTAIL.n121 VTAIL.n99 171.744
R122 VTAIL.n114 VTAIL.n99 171.744
R123 VTAIL.n114 VTAIL.n113 171.744
R124 VTAIL.n113 VTAIL.n103 171.744
R125 VTAIL.n106 VTAIL.n103 171.744
R126 VTAIL.n234 VTAIL.t7 85.8723
R127 VTAIL.n10 VTAIL.t6 85.8723
R128 VTAIL.n42 VTAIL.t0 85.8723
R129 VTAIL.n74 VTAIL.t1 85.8723
R130 VTAIL.n202 VTAIL.t3 85.8723
R131 VTAIL.n170 VTAIL.t2 85.8723
R132 VTAIL.n138 VTAIL.t4 85.8723
R133 VTAIL.n106 VTAIL.t5 85.8723
R134 VTAIL.n255 VTAIL.n254 32.7672
R135 VTAIL.n31 VTAIL.n30 32.7672
R136 VTAIL.n63 VTAIL.n62 32.7672
R137 VTAIL.n95 VTAIL.n94 32.7672
R138 VTAIL.n223 VTAIL.n222 32.7672
R139 VTAIL.n191 VTAIL.n190 32.7672
R140 VTAIL.n159 VTAIL.n158 32.7672
R141 VTAIL.n127 VTAIL.n126 32.7672
R142 VTAIL.n255 VTAIL.n223 20.1686
R143 VTAIL.n127 VTAIL.n95 20.1686
R144 VTAIL.n235 VTAIL.n233 16.3865
R145 VTAIL.n11 VTAIL.n9 16.3865
R146 VTAIL.n43 VTAIL.n41 16.3865
R147 VTAIL.n75 VTAIL.n73 16.3865
R148 VTAIL.n203 VTAIL.n201 16.3865
R149 VTAIL.n171 VTAIL.n169 16.3865
R150 VTAIL.n139 VTAIL.n137 16.3865
R151 VTAIL.n107 VTAIL.n105 16.3865
R152 VTAIL.n236 VTAIL.n232 12.8005
R153 VTAIL.n12 VTAIL.n8 12.8005
R154 VTAIL.n44 VTAIL.n40 12.8005
R155 VTAIL.n76 VTAIL.n72 12.8005
R156 VTAIL.n204 VTAIL.n200 12.8005
R157 VTAIL.n172 VTAIL.n168 12.8005
R158 VTAIL.n140 VTAIL.n136 12.8005
R159 VTAIL.n108 VTAIL.n104 12.8005
R160 VTAIL.n240 VTAIL.n239 12.0247
R161 VTAIL.n16 VTAIL.n15 12.0247
R162 VTAIL.n48 VTAIL.n47 12.0247
R163 VTAIL.n80 VTAIL.n79 12.0247
R164 VTAIL.n208 VTAIL.n207 12.0247
R165 VTAIL.n176 VTAIL.n175 12.0247
R166 VTAIL.n144 VTAIL.n143 12.0247
R167 VTAIL.n112 VTAIL.n111 12.0247
R168 VTAIL.n243 VTAIL.n230 11.249
R169 VTAIL.n19 VTAIL.n6 11.249
R170 VTAIL.n51 VTAIL.n38 11.249
R171 VTAIL.n83 VTAIL.n70 11.249
R172 VTAIL.n211 VTAIL.n198 11.249
R173 VTAIL.n179 VTAIL.n166 11.249
R174 VTAIL.n147 VTAIL.n134 11.249
R175 VTAIL.n115 VTAIL.n102 11.249
R176 VTAIL.n244 VTAIL.n228 10.4732
R177 VTAIL.n20 VTAIL.n4 10.4732
R178 VTAIL.n52 VTAIL.n36 10.4732
R179 VTAIL.n84 VTAIL.n68 10.4732
R180 VTAIL.n212 VTAIL.n196 10.4732
R181 VTAIL.n180 VTAIL.n164 10.4732
R182 VTAIL.n148 VTAIL.n132 10.4732
R183 VTAIL.n116 VTAIL.n100 10.4732
R184 VTAIL.n248 VTAIL.n247 9.69747
R185 VTAIL.n24 VTAIL.n23 9.69747
R186 VTAIL.n56 VTAIL.n55 9.69747
R187 VTAIL.n88 VTAIL.n87 9.69747
R188 VTAIL.n216 VTAIL.n215 9.69747
R189 VTAIL.n184 VTAIL.n183 9.69747
R190 VTAIL.n152 VTAIL.n151 9.69747
R191 VTAIL.n120 VTAIL.n119 9.69747
R192 VTAIL.n254 VTAIL.n253 9.45567
R193 VTAIL.n30 VTAIL.n29 9.45567
R194 VTAIL.n62 VTAIL.n61 9.45567
R195 VTAIL.n94 VTAIL.n93 9.45567
R196 VTAIL.n222 VTAIL.n221 9.45567
R197 VTAIL.n190 VTAIL.n189 9.45567
R198 VTAIL.n158 VTAIL.n157 9.45567
R199 VTAIL.n126 VTAIL.n125 9.45567
R200 VTAIL.n253 VTAIL.n252 9.3005
R201 VTAIL.n226 VTAIL.n225 9.3005
R202 VTAIL.n247 VTAIL.n246 9.3005
R203 VTAIL.n245 VTAIL.n244 9.3005
R204 VTAIL.n230 VTAIL.n229 9.3005
R205 VTAIL.n239 VTAIL.n238 9.3005
R206 VTAIL.n237 VTAIL.n236 9.3005
R207 VTAIL.n29 VTAIL.n28 9.3005
R208 VTAIL.n2 VTAIL.n1 9.3005
R209 VTAIL.n23 VTAIL.n22 9.3005
R210 VTAIL.n21 VTAIL.n20 9.3005
R211 VTAIL.n6 VTAIL.n5 9.3005
R212 VTAIL.n15 VTAIL.n14 9.3005
R213 VTAIL.n13 VTAIL.n12 9.3005
R214 VTAIL.n61 VTAIL.n60 9.3005
R215 VTAIL.n34 VTAIL.n33 9.3005
R216 VTAIL.n55 VTAIL.n54 9.3005
R217 VTAIL.n53 VTAIL.n52 9.3005
R218 VTAIL.n38 VTAIL.n37 9.3005
R219 VTAIL.n47 VTAIL.n46 9.3005
R220 VTAIL.n45 VTAIL.n44 9.3005
R221 VTAIL.n93 VTAIL.n92 9.3005
R222 VTAIL.n66 VTAIL.n65 9.3005
R223 VTAIL.n87 VTAIL.n86 9.3005
R224 VTAIL.n85 VTAIL.n84 9.3005
R225 VTAIL.n70 VTAIL.n69 9.3005
R226 VTAIL.n79 VTAIL.n78 9.3005
R227 VTAIL.n77 VTAIL.n76 9.3005
R228 VTAIL.n221 VTAIL.n220 9.3005
R229 VTAIL.n194 VTAIL.n193 9.3005
R230 VTAIL.n215 VTAIL.n214 9.3005
R231 VTAIL.n213 VTAIL.n212 9.3005
R232 VTAIL.n198 VTAIL.n197 9.3005
R233 VTAIL.n207 VTAIL.n206 9.3005
R234 VTAIL.n205 VTAIL.n204 9.3005
R235 VTAIL.n189 VTAIL.n188 9.3005
R236 VTAIL.n162 VTAIL.n161 9.3005
R237 VTAIL.n183 VTAIL.n182 9.3005
R238 VTAIL.n181 VTAIL.n180 9.3005
R239 VTAIL.n166 VTAIL.n165 9.3005
R240 VTAIL.n175 VTAIL.n174 9.3005
R241 VTAIL.n173 VTAIL.n172 9.3005
R242 VTAIL.n157 VTAIL.n156 9.3005
R243 VTAIL.n130 VTAIL.n129 9.3005
R244 VTAIL.n151 VTAIL.n150 9.3005
R245 VTAIL.n149 VTAIL.n148 9.3005
R246 VTAIL.n134 VTAIL.n133 9.3005
R247 VTAIL.n143 VTAIL.n142 9.3005
R248 VTAIL.n141 VTAIL.n140 9.3005
R249 VTAIL.n125 VTAIL.n124 9.3005
R250 VTAIL.n98 VTAIL.n97 9.3005
R251 VTAIL.n119 VTAIL.n118 9.3005
R252 VTAIL.n117 VTAIL.n116 9.3005
R253 VTAIL.n102 VTAIL.n101 9.3005
R254 VTAIL.n111 VTAIL.n110 9.3005
R255 VTAIL.n109 VTAIL.n108 9.3005
R256 VTAIL.n251 VTAIL.n226 8.92171
R257 VTAIL.n27 VTAIL.n2 8.92171
R258 VTAIL.n59 VTAIL.n34 8.92171
R259 VTAIL.n91 VTAIL.n66 8.92171
R260 VTAIL.n219 VTAIL.n194 8.92171
R261 VTAIL.n187 VTAIL.n162 8.92171
R262 VTAIL.n155 VTAIL.n130 8.92171
R263 VTAIL.n123 VTAIL.n98 8.92171
R264 VTAIL.n252 VTAIL.n224 8.14595
R265 VTAIL.n28 VTAIL.n0 8.14595
R266 VTAIL.n60 VTAIL.n32 8.14595
R267 VTAIL.n92 VTAIL.n64 8.14595
R268 VTAIL.n220 VTAIL.n192 8.14595
R269 VTAIL.n188 VTAIL.n160 8.14595
R270 VTAIL.n156 VTAIL.n128 8.14595
R271 VTAIL.n124 VTAIL.n96 8.14595
R272 VTAIL.n254 VTAIL.n224 5.81868
R273 VTAIL.n30 VTAIL.n0 5.81868
R274 VTAIL.n62 VTAIL.n32 5.81868
R275 VTAIL.n94 VTAIL.n64 5.81868
R276 VTAIL.n222 VTAIL.n192 5.81868
R277 VTAIL.n190 VTAIL.n160 5.81868
R278 VTAIL.n158 VTAIL.n128 5.81868
R279 VTAIL.n126 VTAIL.n96 5.81868
R280 VTAIL.n252 VTAIL.n251 5.04292
R281 VTAIL.n28 VTAIL.n27 5.04292
R282 VTAIL.n60 VTAIL.n59 5.04292
R283 VTAIL.n92 VTAIL.n91 5.04292
R284 VTAIL.n220 VTAIL.n219 5.04292
R285 VTAIL.n188 VTAIL.n187 5.04292
R286 VTAIL.n156 VTAIL.n155 5.04292
R287 VTAIL.n124 VTAIL.n123 5.04292
R288 VTAIL.n248 VTAIL.n226 4.26717
R289 VTAIL.n24 VTAIL.n2 4.26717
R290 VTAIL.n56 VTAIL.n34 4.26717
R291 VTAIL.n88 VTAIL.n66 4.26717
R292 VTAIL.n216 VTAIL.n194 4.26717
R293 VTAIL.n184 VTAIL.n162 4.26717
R294 VTAIL.n152 VTAIL.n130 4.26717
R295 VTAIL.n120 VTAIL.n98 4.26717
R296 VTAIL.n205 VTAIL.n201 3.71286
R297 VTAIL.n173 VTAIL.n169 3.71286
R298 VTAIL.n141 VTAIL.n137 3.71286
R299 VTAIL.n109 VTAIL.n105 3.71286
R300 VTAIL.n237 VTAIL.n233 3.71286
R301 VTAIL.n13 VTAIL.n9 3.71286
R302 VTAIL.n45 VTAIL.n41 3.71286
R303 VTAIL.n77 VTAIL.n73 3.71286
R304 VTAIL.n247 VTAIL.n228 3.49141
R305 VTAIL.n23 VTAIL.n4 3.49141
R306 VTAIL.n55 VTAIL.n36 3.49141
R307 VTAIL.n87 VTAIL.n68 3.49141
R308 VTAIL.n215 VTAIL.n196 3.49141
R309 VTAIL.n183 VTAIL.n164 3.49141
R310 VTAIL.n151 VTAIL.n132 3.49141
R311 VTAIL.n119 VTAIL.n100 3.49141
R312 VTAIL.n244 VTAIL.n243 2.71565
R313 VTAIL.n20 VTAIL.n19 2.71565
R314 VTAIL.n52 VTAIL.n51 2.71565
R315 VTAIL.n84 VTAIL.n83 2.71565
R316 VTAIL.n212 VTAIL.n211 2.71565
R317 VTAIL.n180 VTAIL.n179 2.71565
R318 VTAIL.n148 VTAIL.n147 2.71565
R319 VTAIL.n116 VTAIL.n115 2.71565
R320 VTAIL.n159 VTAIL.n127 2.60395
R321 VTAIL.n223 VTAIL.n191 2.60395
R322 VTAIL.n95 VTAIL.n63 2.60395
R323 VTAIL.n240 VTAIL.n230 1.93989
R324 VTAIL.n16 VTAIL.n6 1.93989
R325 VTAIL.n48 VTAIL.n38 1.93989
R326 VTAIL.n80 VTAIL.n70 1.93989
R327 VTAIL.n208 VTAIL.n198 1.93989
R328 VTAIL.n176 VTAIL.n166 1.93989
R329 VTAIL.n144 VTAIL.n134 1.93989
R330 VTAIL.n112 VTAIL.n102 1.93989
R331 VTAIL VTAIL.n31 1.36041
R332 VTAIL VTAIL.n255 1.24403
R333 VTAIL.n239 VTAIL.n232 1.16414
R334 VTAIL.n15 VTAIL.n8 1.16414
R335 VTAIL.n47 VTAIL.n40 1.16414
R336 VTAIL.n79 VTAIL.n72 1.16414
R337 VTAIL.n207 VTAIL.n200 1.16414
R338 VTAIL.n175 VTAIL.n168 1.16414
R339 VTAIL.n143 VTAIL.n136 1.16414
R340 VTAIL.n111 VTAIL.n104 1.16414
R341 VTAIL.n191 VTAIL.n159 0.470328
R342 VTAIL.n63 VTAIL.n31 0.470328
R343 VTAIL.n236 VTAIL.n235 0.388379
R344 VTAIL.n12 VTAIL.n11 0.388379
R345 VTAIL.n44 VTAIL.n43 0.388379
R346 VTAIL.n76 VTAIL.n75 0.388379
R347 VTAIL.n204 VTAIL.n203 0.388379
R348 VTAIL.n172 VTAIL.n171 0.388379
R349 VTAIL.n140 VTAIL.n139 0.388379
R350 VTAIL.n108 VTAIL.n107 0.388379
R351 VTAIL.n238 VTAIL.n237 0.155672
R352 VTAIL.n238 VTAIL.n229 0.155672
R353 VTAIL.n245 VTAIL.n229 0.155672
R354 VTAIL.n246 VTAIL.n245 0.155672
R355 VTAIL.n246 VTAIL.n225 0.155672
R356 VTAIL.n253 VTAIL.n225 0.155672
R357 VTAIL.n14 VTAIL.n13 0.155672
R358 VTAIL.n14 VTAIL.n5 0.155672
R359 VTAIL.n21 VTAIL.n5 0.155672
R360 VTAIL.n22 VTAIL.n21 0.155672
R361 VTAIL.n22 VTAIL.n1 0.155672
R362 VTAIL.n29 VTAIL.n1 0.155672
R363 VTAIL.n46 VTAIL.n45 0.155672
R364 VTAIL.n46 VTAIL.n37 0.155672
R365 VTAIL.n53 VTAIL.n37 0.155672
R366 VTAIL.n54 VTAIL.n53 0.155672
R367 VTAIL.n54 VTAIL.n33 0.155672
R368 VTAIL.n61 VTAIL.n33 0.155672
R369 VTAIL.n78 VTAIL.n77 0.155672
R370 VTAIL.n78 VTAIL.n69 0.155672
R371 VTAIL.n85 VTAIL.n69 0.155672
R372 VTAIL.n86 VTAIL.n85 0.155672
R373 VTAIL.n86 VTAIL.n65 0.155672
R374 VTAIL.n93 VTAIL.n65 0.155672
R375 VTAIL.n221 VTAIL.n193 0.155672
R376 VTAIL.n214 VTAIL.n193 0.155672
R377 VTAIL.n214 VTAIL.n213 0.155672
R378 VTAIL.n213 VTAIL.n197 0.155672
R379 VTAIL.n206 VTAIL.n197 0.155672
R380 VTAIL.n206 VTAIL.n205 0.155672
R381 VTAIL.n189 VTAIL.n161 0.155672
R382 VTAIL.n182 VTAIL.n161 0.155672
R383 VTAIL.n182 VTAIL.n181 0.155672
R384 VTAIL.n181 VTAIL.n165 0.155672
R385 VTAIL.n174 VTAIL.n165 0.155672
R386 VTAIL.n174 VTAIL.n173 0.155672
R387 VTAIL.n157 VTAIL.n129 0.155672
R388 VTAIL.n150 VTAIL.n129 0.155672
R389 VTAIL.n150 VTAIL.n149 0.155672
R390 VTAIL.n149 VTAIL.n133 0.155672
R391 VTAIL.n142 VTAIL.n133 0.155672
R392 VTAIL.n142 VTAIL.n141 0.155672
R393 VTAIL.n125 VTAIL.n97 0.155672
R394 VTAIL.n118 VTAIL.n97 0.155672
R395 VTAIL.n118 VTAIL.n117 0.155672
R396 VTAIL.n117 VTAIL.n101 0.155672
R397 VTAIL.n110 VTAIL.n101 0.155672
R398 VTAIL.n110 VTAIL.n109 0.155672
R399 VDD2.n2 VDD2.n0 129.6
R400 VDD2.n2 VDD2.n1 92.8759
R401 VDD2.n1 VDD2.t1 5.39105
R402 VDD2.n1 VDD2.t0 5.39105
R403 VDD2.n0 VDD2.t2 5.39105
R404 VDD2.n0 VDD2.t3 5.39105
R405 VDD2 VDD2.n2 0.0586897
R406 VP.n16 VP.n0 161.3
R407 VP.n15 VP.n14 161.3
R408 VP.n13 VP.n1 161.3
R409 VP.n12 VP.n11 161.3
R410 VP.n10 VP.n2 161.3
R411 VP.n9 VP.n8 161.3
R412 VP.n7 VP.n3 161.3
R413 VP.n6 VP.n5 110.267
R414 VP.n18 VP.n17 110.267
R415 VP.n4 VP.t2 87.9394
R416 VP.n4 VP.t0 87.0709
R417 VP.n5 VP.t3 54.0239
R418 VP.n17 VP.t1 54.0239
R419 VP.n6 VP.n4 45.6274
R420 VP.n11 VP.n10 40.4934
R421 VP.n11 VP.n1 40.4934
R422 VP.n9 VP.n3 24.4675
R423 VP.n10 VP.n9 24.4675
R424 VP.n15 VP.n1 24.4675
R425 VP.n16 VP.n15 24.4675
R426 VP.n5 VP.n3 0.48984
R427 VP.n17 VP.n16 0.48984
R428 VP.n7 VP.n6 0.278367
R429 VP.n18 VP.n0 0.278367
R430 VP.n8 VP.n7 0.189894
R431 VP.n8 VP.n2 0.189894
R432 VP.n12 VP.n2 0.189894
R433 VP.n13 VP.n12 0.189894
R434 VP.n14 VP.n13 0.189894
R435 VP.n14 VP.n0 0.189894
R436 VP VP.n18 0.153454
R437 VDD1 VDD1.n1 130.125
R438 VDD1 VDD1.n0 92.9341
R439 VDD1.n0 VDD1.t1 5.39105
R440 VDD1.n0 VDD1.t3 5.39105
R441 VDD1.n1 VDD1.t0 5.39105
R442 VDD1.n1 VDD1.t2 5.39105
R443 B.n275 B.n274 585
R444 B.n273 B.n88 585
R445 B.n272 B.n271 585
R446 B.n270 B.n89 585
R447 B.n269 B.n268 585
R448 B.n267 B.n90 585
R449 B.n266 B.n265 585
R450 B.n264 B.n91 585
R451 B.n263 B.n262 585
R452 B.n261 B.n92 585
R453 B.n260 B.n259 585
R454 B.n258 B.n93 585
R455 B.n257 B.n256 585
R456 B.n255 B.n94 585
R457 B.n254 B.n253 585
R458 B.n252 B.n95 585
R459 B.n251 B.n250 585
R460 B.n249 B.n96 585
R461 B.n248 B.n247 585
R462 B.n246 B.n97 585
R463 B.n245 B.n244 585
R464 B.n243 B.n98 585
R465 B.n242 B.n241 585
R466 B.n240 B.n99 585
R467 B.n238 B.n237 585
R468 B.n236 B.n102 585
R469 B.n235 B.n234 585
R470 B.n233 B.n103 585
R471 B.n232 B.n231 585
R472 B.n230 B.n104 585
R473 B.n229 B.n228 585
R474 B.n227 B.n105 585
R475 B.n226 B.n225 585
R476 B.n224 B.n106 585
R477 B.n223 B.n222 585
R478 B.n218 B.n107 585
R479 B.n217 B.n216 585
R480 B.n215 B.n108 585
R481 B.n214 B.n213 585
R482 B.n212 B.n109 585
R483 B.n211 B.n210 585
R484 B.n209 B.n110 585
R485 B.n208 B.n207 585
R486 B.n206 B.n111 585
R487 B.n205 B.n204 585
R488 B.n203 B.n112 585
R489 B.n202 B.n201 585
R490 B.n200 B.n113 585
R491 B.n199 B.n198 585
R492 B.n197 B.n114 585
R493 B.n196 B.n195 585
R494 B.n194 B.n115 585
R495 B.n193 B.n192 585
R496 B.n191 B.n116 585
R497 B.n190 B.n189 585
R498 B.n188 B.n117 585
R499 B.n187 B.n186 585
R500 B.n185 B.n118 585
R501 B.n276 B.n87 585
R502 B.n278 B.n277 585
R503 B.n279 B.n86 585
R504 B.n281 B.n280 585
R505 B.n282 B.n85 585
R506 B.n284 B.n283 585
R507 B.n285 B.n84 585
R508 B.n287 B.n286 585
R509 B.n288 B.n83 585
R510 B.n290 B.n289 585
R511 B.n291 B.n82 585
R512 B.n293 B.n292 585
R513 B.n294 B.n81 585
R514 B.n296 B.n295 585
R515 B.n297 B.n80 585
R516 B.n299 B.n298 585
R517 B.n300 B.n79 585
R518 B.n302 B.n301 585
R519 B.n303 B.n78 585
R520 B.n305 B.n304 585
R521 B.n306 B.n77 585
R522 B.n308 B.n307 585
R523 B.n309 B.n76 585
R524 B.n311 B.n310 585
R525 B.n312 B.n75 585
R526 B.n314 B.n313 585
R527 B.n315 B.n74 585
R528 B.n317 B.n316 585
R529 B.n318 B.n73 585
R530 B.n320 B.n319 585
R531 B.n321 B.n72 585
R532 B.n323 B.n322 585
R533 B.n324 B.n71 585
R534 B.n326 B.n325 585
R535 B.n327 B.n70 585
R536 B.n329 B.n328 585
R537 B.n330 B.n69 585
R538 B.n332 B.n331 585
R539 B.n333 B.n68 585
R540 B.n335 B.n334 585
R541 B.n336 B.n67 585
R542 B.n338 B.n337 585
R543 B.n339 B.n66 585
R544 B.n341 B.n340 585
R545 B.n342 B.n65 585
R546 B.n344 B.n343 585
R547 B.n345 B.n64 585
R548 B.n347 B.n346 585
R549 B.n348 B.n63 585
R550 B.n350 B.n349 585
R551 B.n351 B.n62 585
R552 B.n353 B.n352 585
R553 B.n354 B.n61 585
R554 B.n356 B.n355 585
R555 B.n357 B.n60 585
R556 B.n359 B.n358 585
R557 B.n360 B.n59 585
R558 B.n362 B.n361 585
R559 B.n363 B.n58 585
R560 B.n365 B.n364 585
R561 B.n366 B.n57 585
R562 B.n368 B.n367 585
R563 B.n369 B.n56 585
R564 B.n371 B.n370 585
R565 B.n372 B.n55 585
R566 B.n374 B.n373 585
R567 B.n375 B.n54 585
R568 B.n377 B.n376 585
R569 B.n378 B.n53 585
R570 B.n380 B.n379 585
R571 B.n468 B.n19 585
R572 B.n467 B.n466 585
R573 B.n465 B.n20 585
R574 B.n464 B.n463 585
R575 B.n462 B.n21 585
R576 B.n461 B.n460 585
R577 B.n459 B.n22 585
R578 B.n458 B.n457 585
R579 B.n456 B.n23 585
R580 B.n455 B.n454 585
R581 B.n453 B.n24 585
R582 B.n452 B.n451 585
R583 B.n450 B.n25 585
R584 B.n449 B.n448 585
R585 B.n447 B.n26 585
R586 B.n446 B.n445 585
R587 B.n444 B.n27 585
R588 B.n443 B.n442 585
R589 B.n441 B.n28 585
R590 B.n440 B.n439 585
R591 B.n438 B.n29 585
R592 B.n437 B.n436 585
R593 B.n435 B.n30 585
R594 B.n434 B.n433 585
R595 B.n431 B.n31 585
R596 B.n430 B.n429 585
R597 B.n428 B.n34 585
R598 B.n427 B.n426 585
R599 B.n425 B.n35 585
R600 B.n424 B.n423 585
R601 B.n422 B.n36 585
R602 B.n421 B.n420 585
R603 B.n419 B.n37 585
R604 B.n418 B.n417 585
R605 B.n416 B.n415 585
R606 B.n414 B.n41 585
R607 B.n413 B.n412 585
R608 B.n411 B.n42 585
R609 B.n410 B.n409 585
R610 B.n408 B.n43 585
R611 B.n407 B.n406 585
R612 B.n405 B.n44 585
R613 B.n404 B.n403 585
R614 B.n402 B.n45 585
R615 B.n401 B.n400 585
R616 B.n399 B.n46 585
R617 B.n398 B.n397 585
R618 B.n396 B.n47 585
R619 B.n395 B.n394 585
R620 B.n393 B.n48 585
R621 B.n392 B.n391 585
R622 B.n390 B.n49 585
R623 B.n389 B.n388 585
R624 B.n387 B.n50 585
R625 B.n386 B.n385 585
R626 B.n384 B.n51 585
R627 B.n383 B.n382 585
R628 B.n381 B.n52 585
R629 B.n470 B.n469 585
R630 B.n471 B.n18 585
R631 B.n473 B.n472 585
R632 B.n474 B.n17 585
R633 B.n476 B.n475 585
R634 B.n477 B.n16 585
R635 B.n479 B.n478 585
R636 B.n480 B.n15 585
R637 B.n482 B.n481 585
R638 B.n483 B.n14 585
R639 B.n485 B.n484 585
R640 B.n486 B.n13 585
R641 B.n488 B.n487 585
R642 B.n489 B.n12 585
R643 B.n491 B.n490 585
R644 B.n492 B.n11 585
R645 B.n494 B.n493 585
R646 B.n495 B.n10 585
R647 B.n497 B.n496 585
R648 B.n498 B.n9 585
R649 B.n500 B.n499 585
R650 B.n501 B.n8 585
R651 B.n503 B.n502 585
R652 B.n504 B.n7 585
R653 B.n506 B.n505 585
R654 B.n507 B.n6 585
R655 B.n509 B.n508 585
R656 B.n510 B.n5 585
R657 B.n512 B.n511 585
R658 B.n513 B.n4 585
R659 B.n515 B.n514 585
R660 B.n516 B.n3 585
R661 B.n518 B.n517 585
R662 B.n519 B.n0 585
R663 B.n2 B.n1 585
R664 B.n136 B.n135 585
R665 B.n137 B.n134 585
R666 B.n139 B.n138 585
R667 B.n140 B.n133 585
R668 B.n142 B.n141 585
R669 B.n143 B.n132 585
R670 B.n145 B.n144 585
R671 B.n146 B.n131 585
R672 B.n148 B.n147 585
R673 B.n149 B.n130 585
R674 B.n151 B.n150 585
R675 B.n152 B.n129 585
R676 B.n154 B.n153 585
R677 B.n155 B.n128 585
R678 B.n157 B.n156 585
R679 B.n158 B.n127 585
R680 B.n160 B.n159 585
R681 B.n161 B.n126 585
R682 B.n163 B.n162 585
R683 B.n164 B.n125 585
R684 B.n166 B.n165 585
R685 B.n167 B.n124 585
R686 B.n169 B.n168 585
R687 B.n170 B.n123 585
R688 B.n172 B.n171 585
R689 B.n173 B.n122 585
R690 B.n175 B.n174 585
R691 B.n176 B.n121 585
R692 B.n178 B.n177 585
R693 B.n179 B.n120 585
R694 B.n181 B.n180 585
R695 B.n182 B.n119 585
R696 B.n184 B.n183 585
R697 B.n185 B.n184 516.524
R698 B.n274 B.n87 516.524
R699 B.n381 B.n380 516.524
R700 B.n470 B.n19 516.524
R701 B.n100 B.t10 327.344
R702 B.n38 B.t8 327.344
R703 B.n219 B.t4 327.344
R704 B.n32 B.t2 327.344
R705 B.n101 B.t11 268.774
R706 B.n39 B.t7 268.774
R707 B.n220 B.t5 268.774
R708 B.n33 B.t1 268.774
R709 B.n219 B.t3 262.202
R710 B.n100 B.t9 262.202
R711 B.n38 B.t6 262.202
R712 B.n32 B.t0 262.202
R713 B.n521 B.n520 256.663
R714 B.n520 B.n519 235.042
R715 B.n520 B.n2 235.042
R716 B.n186 B.n185 163.367
R717 B.n186 B.n117 163.367
R718 B.n190 B.n117 163.367
R719 B.n191 B.n190 163.367
R720 B.n192 B.n191 163.367
R721 B.n192 B.n115 163.367
R722 B.n196 B.n115 163.367
R723 B.n197 B.n196 163.367
R724 B.n198 B.n197 163.367
R725 B.n198 B.n113 163.367
R726 B.n202 B.n113 163.367
R727 B.n203 B.n202 163.367
R728 B.n204 B.n203 163.367
R729 B.n204 B.n111 163.367
R730 B.n208 B.n111 163.367
R731 B.n209 B.n208 163.367
R732 B.n210 B.n209 163.367
R733 B.n210 B.n109 163.367
R734 B.n214 B.n109 163.367
R735 B.n215 B.n214 163.367
R736 B.n216 B.n215 163.367
R737 B.n216 B.n107 163.367
R738 B.n223 B.n107 163.367
R739 B.n224 B.n223 163.367
R740 B.n225 B.n224 163.367
R741 B.n225 B.n105 163.367
R742 B.n229 B.n105 163.367
R743 B.n230 B.n229 163.367
R744 B.n231 B.n230 163.367
R745 B.n231 B.n103 163.367
R746 B.n235 B.n103 163.367
R747 B.n236 B.n235 163.367
R748 B.n237 B.n236 163.367
R749 B.n237 B.n99 163.367
R750 B.n242 B.n99 163.367
R751 B.n243 B.n242 163.367
R752 B.n244 B.n243 163.367
R753 B.n244 B.n97 163.367
R754 B.n248 B.n97 163.367
R755 B.n249 B.n248 163.367
R756 B.n250 B.n249 163.367
R757 B.n250 B.n95 163.367
R758 B.n254 B.n95 163.367
R759 B.n255 B.n254 163.367
R760 B.n256 B.n255 163.367
R761 B.n256 B.n93 163.367
R762 B.n260 B.n93 163.367
R763 B.n261 B.n260 163.367
R764 B.n262 B.n261 163.367
R765 B.n262 B.n91 163.367
R766 B.n266 B.n91 163.367
R767 B.n267 B.n266 163.367
R768 B.n268 B.n267 163.367
R769 B.n268 B.n89 163.367
R770 B.n272 B.n89 163.367
R771 B.n273 B.n272 163.367
R772 B.n274 B.n273 163.367
R773 B.n380 B.n53 163.367
R774 B.n376 B.n53 163.367
R775 B.n376 B.n375 163.367
R776 B.n375 B.n374 163.367
R777 B.n374 B.n55 163.367
R778 B.n370 B.n55 163.367
R779 B.n370 B.n369 163.367
R780 B.n369 B.n368 163.367
R781 B.n368 B.n57 163.367
R782 B.n364 B.n57 163.367
R783 B.n364 B.n363 163.367
R784 B.n363 B.n362 163.367
R785 B.n362 B.n59 163.367
R786 B.n358 B.n59 163.367
R787 B.n358 B.n357 163.367
R788 B.n357 B.n356 163.367
R789 B.n356 B.n61 163.367
R790 B.n352 B.n61 163.367
R791 B.n352 B.n351 163.367
R792 B.n351 B.n350 163.367
R793 B.n350 B.n63 163.367
R794 B.n346 B.n63 163.367
R795 B.n346 B.n345 163.367
R796 B.n345 B.n344 163.367
R797 B.n344 B.n65 163.367
R798 B.n340 B.n65 163.367
R799 B.n340 B.n339 163.367
R800 B.n339 B.n338 163.367
R801 B.n338 B.n67 163.367
R802 B.n334 B.n67 163.367
R803 B.n334 B.n333 163.367
R804 B.n333 B.n332 163.367
R805 B.n332 B.n69 163.367
R806 B.n328 B.n69 163.367
R807 B.n328 B.n327 163.367
R808 B.n327 B.n326 163.367
R809 B.n326 B.n71 163.367
R810 B.n322 B.n71 163.367
R811 B.n322 B.n321 163.367
R812 B.n321 B.n320 163.367
R813 B.n320 B.n73 163.367
R814 B.n316 B.n73 163.367
R815 B.n316 B.n315 163.367
R816 B.n315 B.n314 163.367
R817 B.n314 B.n75 163.367
R818 B.n310 B.n75 163.367
R819 B.n310 B.n309 163.367
R820 B.n309 B.n308 163.367
R821 B.n308 B.n77 163.367
R822 B.n304 B.n77 163.367
R823 B.n304 B.n303 163.367
R824 B.n303 B.n302 163.367
R825 B.n302 B.n79 163.367
R826 B.n298 B.n79 163.367
R827 B.n298 B.n297 163.367
R828 B.n297 B.n296 163.367
R829 B.n296 B.n81 163.367
R830 B.n292 B.n81 163.367
R831 B.n292 B.n291 163.367
R832 B.n291 B.n290 163.367
R833 B.n290 B.n83 163.367
R834 B.n286 B.n83 163.367
R835 B.n286 B.n285 163.367
R836 B.n285 B.n284 163.367
R837 B.n284 B.n85 163.367
R838 B.n280 B.n85 163.367
R839 B.n280 B.n279 163.367
R840 B.n279 B.n278 163.367
R841 B.n278 B.n87 163.367
R842 B.n466 B.n19 163.367
R843 B.n466 B.n465 163.367
R844 B.n465 B.n464 163.367
R845 B.n464 B.n21 163.367
R846 B.n460 B.n21 163.367
R847 B.n460 B.n459 163.367
R848 B.n459 B.n458 163.367
R849 B.n458 B.n23 163.367
R850 B.n454 B.n23 163.367
R851 B.n454 B.n453 163.367
R852 B.n453 B.n452 163.367
R853 B.n452 B.n25 163.367
R854 B.n448 B.n25 163.367
R855 B.n448 B.n447 163.367
R856 B.n447 B.n446 163.367
R857 B.n446 B.n27 163.367
R858 B.n442 B.n27 163.367
R859 B.n442 B.n441 163.367
R860 B.n441 B.n440 163.367
R861 B.n440 B.n29 163.367
R862 B.n436 B.n29 163.367
R863 B.n436 B.n435 163.367
R864 B.n435 B.n434 163.367
R865 B.n434 B.n31 163.367
R866 B.n429 B.n31 163.367
R867 B.n429 B.n428 163.367
R868 B.n428 B.n427 163.367
R869 B.n427 B.n35 163.367
R870 B.n423 B.n35 163.367
R871 B.n423 B.n422 163.367
R872 B.n422 B.n421 163.367
R873 B.n421 B.n37 163.367
R874 B.n417 B.n37 163.367
R875 B.n417 B.n416 163.367
R876 B.n416 B.n41 163.367
R877 B.n412 B.n41 163.367
R878 B.n412 B.n411 163.367
R879 B.n411 B.n410 163.367
R880 B.n410 B.n43 163.367
R881 B.n406 B.n43 163.367
R882 B.n406 B.n405 163.367
R883 B.n405 B.n404 163.367
R884 B.n404 B.n45 163.367
R885 B.n400 B.n45 163.367
R886 B.n400 B.n399 163.367
R887 B.n399 B.n398 163.367
R888 B.n398 B.n47 163.367
R889 B.n394 B.n47 163.367
R890 B.n394 B.n393 163.367
R891 B.n393 B.n392 163.367
R892 B.n392 B.n49 163.367
R893 B.n388 B.n49 163.367
R894 B.n388 B.n387 163.367
R895 B.n387 B.n386 163.367
R896 B.n386 B.n51 163.367
R897 B.n382 B.n51 163.367
R898 B.n382 B.n381 163.367
R899 B.n471 B.n470 163.367
R900 B.n472 B.n471 163.367
R901 B.n472 B.n17 163.367
R902 B.n476 B.n17 163.367
R903 B.n477 B.n476 163.367
R904 B.n478 B.n477 163.367
R905 B.n478 B.n15 163.367
R906 B.n482 B.n15 163.367
R907 B.n483 B.n482 163.367
R908 B.n484 B.n483 163.367
R909 B.n484 B.n13 163.367
R910 B.n488 B.n13 163.367
R911 B.n489 B.n488 163.367
R912 B.n490 B.n489 163.367
R913 B.n490 B.n11 163.367
R914 B.n494 B.n11 163.367
R915 B.n495 B.n494 163.367
R916 B.n496 B.n495 163.367
R917 B.n496 B.n9 163.367
R918 B.n500 B.n9 163.367
R919 B.n501 B.n500 163.367
R920 B.n502 B.n501 163.367
R921 B.n502 B.n7 163.367
R922 B.n506 B.n7 163.367
R923 B.n507 B.n506 163.367
R924 B.n508 B.n507 163.367
R925 B.n508 B.n5 163.367
R926 B.n512 B.n5 163.367
R927 B.n513 B.n512 163.367
R928 B.n514 B.n513 163.367
R929 B.n514 B.n3 163.367
R930 B.n518 B.n3 163.367
R931 B.n519 B.n518 163.367
R932 B.n136 B.n2 163.367
R933 B.n137 B.n136 163.367
R934 B.n138 B.n137 163.367
R935 B.n138 B.n133 163.367
R936 B.n142 B.n133 163.367
R937 B.n143 B.n142 163.367
R938 B.n144 B.n143 163.367
R939 B.n144 B.n131 163.367
R940 B.n148 B.n131 163.367
R941 B.n149 B.n148 163.367
R942 B.n150 B.n149 163.367
R943 B.n150 B.n129 163.367
R944 B.n154 B.n129 163.367
R945 B.n155 B.n154 163.367
R946 B.n156 B.n155 163.367
R947 B.n156 B.n127 163.367
R948 B.n160 B.n127 163.367
R949 B.n161 B.n160 163.367
R950 B.n162 B.n161 163.367
R951 B.n162 B.n125 163.367
R952 B.n166 B.n125 163.367
R953 B.n167 B.n166 163.367
R954 B.n168 B.n167 163.367
R955 B.n168 B.n123 163.367
R956 B.n172 B.n123 163.367
R957 B.n173 B.n172 163.367
R958 B.n174 B.n173 163.367
R959 B.n174 B.n121 163.367
R960 B.n178 B.n121 163.367
R961 B.n179 B.n178 163.367
R962 B.n180 B.n179 163.367
R963 B.n180 B.n119 163.367
R964 B.n184 B.n119 163.367
R965 B.n221 B.n220 59.5399
R966 B.n239 B.n101 59.5399
R967 B.n40 B.n39 59.5399
R968 B.n432 B.n33 59.5399
R969 B.n220 B.n219 58.5702
R970 B.n101 B.n100 58.5702
R971 B.n39 B.n38 58.5702
R972 B.n33 B.n32 58.5702
R973 B.n469 B.n468 33.5615
R974 B.n379 B.n52 33.5615
R975 B.n276 B.n275 33.5615
R976 B.n183 B.n118 33.5615
R977 B B.n521 18.0485
R978 B.n469 B.n18 10.6151
R979 B.n473 B.n18 10.6151
R980 B.n474 B.n473 10.6151
R981 B.n475 B.n474 10.6151
R982 B.n475 B.n16 10.6151
R983 B.n479 B.n16 10.6151
R984 B.n480 B.n479 10.6151
R985 B.n481 B.n480 10.6151
R986 B.n481 B.n14 10.6151
R987 B.n485 B.n14 10.6151
R988 B.n486 B.n485 10.6151
R989 B.n487 B.n486 10.6151
R990 B.n487 B.n12 10.6151
R991 B.n491 B.n12 10.6151
R992 B.n492 B.n491 10.6151
R993 B.n493 B.n492 10.6151
R994 B.n493 B.n10 10.6151
R995 B.n497 B.n10 10.6151
R996 B.n498 B.n497 10.6151
R997 B.n499 B.n498 10.6151
R998 B.n499 B.n8 10.6151
R999 B.n503 B.n8 10.6151
R1000 B.n504 B.n503 10.6151
R1001 B.n505 B.n504 10.6151
R1002 B.n505 B.n6 10.6151
R1003 B.n509 B.n6 10.6151
R1004 B.n510 B.n509 10.6151
R1005 B.n511 B.n510 10.6151
R1006 B.n511 B.n4 10.6151
R1007 B.n515 B.n4 10.6151
R1008 B.n516 B.n515 10.6151
R1009 B.n517 B.n516 10.6151
R1010 B.n517 B.n0 10.6151
R1011 B.n468 B.n467 10.6151
R1012 B.n467 B.n20 10.6151
R1013 B.n463 B.n20 10.6151
R1014 B.n463 B.n462 10.6151
R1015 B.n462 B.n461 10.6151
R1016 B.n461 B.n22 10.6151
R1017 B.n457 B.n22 10.6151
R1018 B.n457 B.n456 10.6151
R1019 B.n456 B.n455 10.6151
R1020 B.n455 B.n24 10.6151
R1021 B.n451 B.n24 10.6151
R1022 B.n451 B.n450 10.6151
R1023 B.n450 B.n449 10.6151
R1024 B.n449 B.n26 10.6151
R1025 B.n445 B.n26 10.6151
R1026 B.n445 B.n444 10.6151
R1027 B.n444 B.n443 10.6151
R1028 B.n443 B.n28 10.6151
R1029 B.n439 B.n28 10.6151
R1030 B.n439 B.n438 10.6151
R1031 B.n438 B.n437 10.6151
R1032 B.n437 B.n30 10.6151
R1033 B.n433 B.n30 10.6151
R1034 B.n431 B.n430 10.6151
R1035 B.n430 B.n34 10.6151
R1036 B.n426 B.n34 10.6151
R1037 B.n426 B.n425 10.6151
R1038 B.n425 B.n424 10.6151
R1039 B.n424 B.n36 10.6151
R1040 B.n420 B.n36 10.6151
R1041 B.n420 B.n419 10.6151
R1042 B.n419 B.n418 10.6151
R1043 B.n415 B.n414 10.6151
R1044 B.n414 B.n413 10.6151
R1045 B.n413 B.n42 10.6151
R1046 B.n409 B.n42 10.6151
R1047 B.n409 B.n408 10.6151
R1048 B.n408 B.n407 10.6151
R1049 B.n407 B.n44 10.6151
R1050 B.n403 B.n44 10.6151
R1051 B.n403 B.n402 10.6151
R1052 B.n402 B.n401 10.6151
R1053 B.n401 B.n46 10.6151
R1054 B.n397 B.n46 10.6151
R1055 B.n397 B.n396 10.6151
R1056 B.n396 B.n395 10.6151
R1057 B.n395 B.n48 10.6151
R1058 B.n391 B.n48 10.6151
R1059 B.n391 B.n390 10.6151
R1060 B.n390 B.n389 10.6151
R1061 B.n389 B.n50 10.6151
R1062 B.n385 B.n50 10.6151
R1063 B.n385 B.n384 10.6151
R1064 B.n384 B.n383 10.6151
R1065 B.n383 B.n52 10.6151
R1066 B.n379 B.n378 10.6151
R1067 B.n378 B.n377 10.6151
R1068 B.n377 B.n54 10.6151
R1069 B.n373 B.n54 10.6151
R1070 B.n373 B.n372 10.6151
R1071 B.n372 B.n371 10.6151
R1072 B.n371 B.n56 10.6151
R1073 B.n367 B.n56 10.6151
R1074 B.n367 B.n366 10.6151
R1075 B.n366 B.n365 10.6151
R1076 B.n365 B.n58 10.6151
R1077 B.n361 B.n58 10.6151
R1078 B.n361 B.n360 10.6151
R1079 B.n360 B.n359 10.6151
R1080 B.n359 B.n60 10.6151
R1081 B.n355 B.n60 10.6151
R1082 B.n355 B.n354 10.6151
R1083 B.n354 B.n353 10.6151
R1084 B.n353 B.n62 10.6151
R1085 B.n349 B.n62 10.6151
R1086 B.n349 B.n348 10.6151
R1087 B.n348 B.n347 10.6151
R1088 B.n347 B.n64 10.6151
R1089 B.n343 B.n64 10.6151
R1090 B.n343 B.n342 10.6151
R1091 B.n342 B.n341 10.6151
R1092 B.n341 B.n66 10.6151
R1093 B.n337 B.n66 10.6151
R1094 B.n337 B.n336 10.6151
R1095 B.n336 B.n335 10.6151
R1096 B.n335 B.n68 10.6151
R1097 B.n331 B.n68 10.6151
R1098 B.n331 B.n330 10.6151
R1099 B.n330 B.n329 10.6151
R1100 B.n329 B.n70 10.6151
R1101 B.n325 B.n70 10.6151
R1102 B.n325 B.n324 10.6151
R1103 B.n324 B.n323 10.6151
R1104 B.n323 B.n72 10.6151
R1105 B.n319 B.n72 10.6151
R1106 B.n319 B.n318 10.6151
R1107 B.n318 B.n317 10.6151
R1108 B.n317 B.n74 10.6151
R1109 B.n313 B.n74 10.6151
R1110 B.n313 B.n312 10.6151
R1111 B.n312 B.n311 10.6151
R1112 B.n311 B.n76 10.6151
R1113 B.n307 B.n76 10.6151
R1114 B.n307 B.n306 10.6151
R1115 B.n306 B.n305 10.6151
R1116 B.n305 B.n78 10.6151
R1117 B.n301 B.n78 10.6151
R1118 B.n301 B.n300 10.6151
R1119 B.n300 B.n299 10.6151
R1120 B.n299 B.n80 10.6151
R1121 B.n295 B.n80 10.6151
R1122 B.n295 B.n294 10.6151
R1123 B.n294 B.n293 10.6151
R1124 B.n293 B.n82 10.6151
R1125 B.n289 B.n82 10.6151
R1126 B.n289 B.n288 10.6151
R1127 B.n288 B.n287 10.6151
R1128 B.n287 B.n84 10.6151
R1129 B.n283 B.n84 10.6151
R1130 B.n283 B.n282 10.6151
R1131 B.n282 B.n281 10.6151
R1132 B.n281 B.n86 10.6151
R1133 B.n277 B.n86 10.6151
R1134 B.n277 B.n276 10.6151
R1135 B.n135 B.n1 10.6151
R1136 B.n135 B.n134 10.6151
R1137 B.n139 B.n134 10.6151
R1138 B.n140 B.n139 10.6151
R1139 B.n141 B.n140 10.6151
R1140 B.n141 B.n132 10.6151
R1141 B.n145 B.n132 10.6151
R1142 B.n146 B.n145 10.6151
R1143 B.n147 B.n146 10.6151
R1144 B.n147 B.n130 10.6151
R1145 B.n151 B.n130 10.6151
R1146 B.n152 B.n151 10.6151
R1147 B.n153 B.n152 10.6151
R1148 B.n153 B.n128 10.6151
R1149 B.n157 B.n128 10.6151
R1150 B.n158 B.n157 10.6151
R1151 B.n159 B.n158 10.6151
R1152 B.n159 B.n126 10.6151
R1153 B.n163 B.n126 10.6151
R1154 B.n164 B.n163 10.6151
R1155 B.n165 B.n164 10.6151
R1156 B.n165 B.n124 10.6151
R1157 B.n169 B.n124 10.6151
R1158 B.n170 B.n169 10.6151
R1159 B.n171 B.n170 10.6151
R1160 B.n171 B.n122 10.6151
R1161 B.n175 B.n122 10.6151
R1162 B.n176 B.n175 10.6151
R1163 B.n177 B.n176 10.6151
R1164 B.n177 B.n120 10.6151
R1165 B.n181 B.n120 10.6151
R1166 B.n182 B.n181 10.6151
R1167 B.n183 B.n182 10.6151
R1168 B.n187 B.n118 10.6151
R1169 B.n188 B.n187 10.6151
R1170 B.n189 B.n188 10.6151
R1171 B.n189 B.n116 10.6151
R1172 B.n193 B.n116 10.6151
R1173 B.n194 B.n193 10.6151
R1174 B.n195 B.n194 10.6151
R1175 B.n195 B.n114 10.6151
R1176 B.n199 B.n114 10.6151
R1177 B.n200 B.n199 10.6151
R1178 B.n201 B.n200 10.6151
R1179 B.n201 B.n112 10.6151
R1180 B.n205 B.n112 10.6151
R1181 B.n206 B.n205 10.6151
R1182 B.n207 B.n206 10.6151
R1183 B.n207 B.n110 10.6151
R1184 B.n211 B.n110 10.6151
R1185 B.n212 B.n211 10.6151
R1186 B.n213 B.n212 10.6151
R1187 B.n213 B.n108 10.6151
R1188 B.n217 B.n108 10.6151
R1189 B.n218 B.n217 10.6151
R1190 B.n222 B.n218 10.6151
R1191 B.n226 B.n106 10.6151
R1192 B.n227 B.n226 10.6151
R1193 B.n228 B.n227 10.6151
R1194 B.n228 B.n104 10.6151
R1195 B.n232 B.n104 10.6151
R1196 B.n233 B.n232 10.6151
R1197 B.n234 B.n233 10.6151
R1198 B.n234 B.n102 10.6151
R1199 B.n238 B.n102 10.6151
R1200 B.n241 B.n240 10.6151
R1201 B.n241 B.n98 10.6151
R1202 B.n245 B.n98 10.6151
R1203 B.n246 B.n245 10.6151
R1204 B.n247 B.n246 10.6151
R1205 B.n247 B.n96 10.6151
R1206 B.n251 B.n96 10.6151
R1207 B.n252 B.n251 10.6151
R1208 B.n253 B.n252 10.6151
R1209 B.n253 B.n94 10.6151
R1210 B.n257 B.n94 10.6151
R1211 B.n258 B.n257 10.6151
R1212 B.n259 B.n258 10.6151
R1213 B.n259 B.n92 10.6151
R1214 B.n263 B.n92 10.6151
R1215 B.n264 B.n263 10.6151
R1216 B.n265 B.n264 10.6151
R1217 B.n265 B.n90 10.6151
R1218 B.n269 B.n90 10.6151
R1219 B.n270 B.n269 10.6151
R1220 B.n271 B.n270 10.6151
R1221 B.n271 B.n88 10.6151
R1222 B.n275 B.n88 10.6151
R1223 B.n433 B.n432 9.36635
R1224 B.n415 B.n40 9.36635
R1225 B.n222 B.n221 9.36635
R1226 B.n240 B.n239 9.36635
R1227 B.n521 B.n0 8.11757
R1228 B.n521 B.n1 8.11757
R1229 B.n432 B.n431 1.24928
R1230 B.n418 B.n40 1.24928
R1231 B.n221 B.n106 1.24928
R1232 B.n239 B.n238 1.24928
C0 VDD2 VDD1 1.04143f
C1 VTAIL VP 2.88234f
C2 VDD1 B 1.11616f
C3 VDD2 w_n2782_n2174# 1.36572f
C4 B w_n2782_n2174# 7.69371f
C5 VDD1 VP 2.8168f
C6 VDD2 B 1.16979f
C7 VTAIL VN 2.86824f
C8 VP w_n2782_n2174# 4.98726f
C9 VDD2 VP 0.399868f
C10 VDD1 VN 0.148917f
C11 VP B 1.64539f
C12 VN w_n2782_n2174# 4.62939f
C13 VDD2 VN 2.56661f
C14 VDD1 VTAIL 4.02113f
C15 VTAIL w_n2782_n2174# 2.63515f
C16 VN B 1.05111f
C17 VDD2 VTAIL 4.07594f
C18 VDD1 w_n2782_n2174# 1.3076f
C19 VTAIL B 3.00706f
C20 VN VP 5.1539f
C21 VDD2 VSUBS 0.827403f
C22 VDD1 VSUBS 5.017149f
C23 VTAIL VSUBS 0.707706f
C24 VN VSUBS 5.36098f
C25 VP VSUBS 1.976365f
C26 B VSUBS 3.851212f
C27 w_n2782_n2174# VSUBS 75.4812f
C28 B.n0 VSUBS 0.007245f
C29 B.n1 VSUBS 0.007245f
C30 B.n2 VSUBS 0.010715f
C31 B.n3 VSUBS 0.008211f
C32 B.n4 VSUBS 0.008211f
C33 B.n5 VSUBS 0.008211f
C34 B.n6 VSUBS 0.008211f
C35 B.n7 VSUBS 0.008211f
C36 B.n8 VSUBS 0.008211f
C37 B.n9 VSUBS 0.008211f
C38 B.n10 VSUBS 0.008211f
C39 B.n11 VSUBS 0.008211f
C40 B.n12 VSUBS 0.008211f
C41 B.n13 VSUBS 0.008211f
C42 B.n14 VSUBS 0.008211f
C43 B.n15 VSUBS 0.008211f
C44 B.n16 VSUBS 0.008211f
C45 B.n17 VSUBS 0.008211f
C46 B.n18 VSUBS 0.008211f
C47 B.n19 VSUBS 0.020334f
C48 B.n20 VSUBS 0.008211f
C49 B.n21 VSUBS 0.008211f
C50 B.n22 VSUBS 0.008211f
C51 B.n23 VSUBS 0.008211f
C52 B.n24 VSUBS 0.008211f
C53 B.n25 VSUBS 0.008211f
C54 B.n26 VSUBS 0.008211f
C55 B.n27 VSUBS 0.008211f
C56 B.n28 VSUBS 0.008211f
C57 B.n29 VSUBS 0.008211f
C58 B.n30 VSUBS 0.008211f
C59 B.n31 VSUBS 0.008211f
C60 B.t1 VSUBS 0.105675f
C61 B.t2 VSUBS 0.136595f
C62 B.t0 VSUBS 0.901238f
C63 B.n32 VSUBS 0.231906f
C64 B.n33 VSUBS 0.184524f
C65 B.n34 VSUBS 0.008211f
C66 B.n35 VSUBS 0.008211f
C67 B.n36 VSUBS 0.008211f
C68 B.n37 VSUBS 0.008211f
C69 B.t7 VSUBS 0.105677f
C70 B.t8 VSUBS 0.136596f
C71 B.t6 VSUBS 0.901238f
C72 B.n38 VSUBS 0.231904f
C73 B.n39 VSUBS 0.184522f
C74 B.n40 VSUBS 0.019025f
C75 B.n41 VSUBS 0.008211f
C76 B.n42 VSUBS 0.008211f
C77 B.n43 VSUBS 0.008211f
C78 B.n44 VSUBS 0.008211f
C79 B.n45 VSUBS 0.008211f
C80 B.n46 VSUBS 0.008211f
C81 B.n47 VSUBS 0.008211f
C82 B.n48 VSUBS 0.008211f
C83 B.n49 VSUBS 0.008211f
C84 B.n50 VSUBS 0.008211f
C85 B.n51 VSUBS 0.008211f
C86 B.n52 VSUBS 0.020334f
C87 B.n53 VSUBS 0.008211f
C88 B.n54 VSUBS 0.008211f
C89 B.n55 VSUBS 0.008211f
C90 B.n56 VSUBS 0.008211f
C91 B.n57 VSUBS 0.008211f
C92 B.n58 VSUBS 0.008211f
C93 B.n59 VSUBS 0.008211f
C94 B.n60 VSUBS 0.008211f
C95 B.n61 VSUBS 0.008211f
C96 B.n62 VSUBS 0.008211f
C97 B.n63 VSUBS 0.008211f
C98 B.n64 VSUBS 0.008211f
C99 B.n65 VSUBS 0.008211f
C100 B.n66 VSUBS 0.008211f
C101 B.n67 VSUBS 0.008211f
C102 B.n68 VSUBS 0.008211f
C103 B.n69 VSUBS 0.008211f
C104 B.n70 VSUBS 0.008211f
C105 B.n71 VSUBS 0.008211f
C106 B.n72 VSUBS 0.008211f
C107 B.n73 VSUBS 0.008211f
C108 B.n74 VSUBS 0.008211f
C109 B.n75 VSUBS 0.008211f
C110 B.n76 VSUBS 0.008211f
C111 B.n77 VSUBS 0.008211f
C112 B.n78 VSUBS 0.008211f
C113 B.n79 VSUBS 0.008211f
C114 B.n80 VSUBS 0.008211f
C115 B.n81 VSUBS 0.008211f
C116 B.n82 VSUBS 0.008211f
C117 B.n83 VSUBS 0.008211f
C118 B.n84 VSUBS 0.008211f
C119 B.n85 VSUBS 0.008211f
C120 B.n86 VSUBS 0.008211f
C121 B.n87 VSUBS 0.018791f
C122 B.n88 VSUBS 0.008211f
C123 B.n89 VSUBS 0.008211f
C124 B.n90 VSUBS 0.008211f
C125 B.n91 VSUBS 0.008211f
C126 B.n92 VSUBS 0.008211f
C127 B.n93 VSUBS 0.008211f
C128 B.n94 VSUBS 0.008211f
C129 B.n95 VSUBS 0.008211f
C130 B.n96 VSUBS 0.008211f
C131 B.n97 VSUBS 0.008211f
C132 B.n98 VSUBS 0.008211f
C133 B.n99 VSUBS 0.008211f
C134 B.t11 VSUBS 0.105677f
C135 B.t10 VSUBS 0.136596f
C136 B.t9 VSUBS 0.901238f
C137 B.n100 VSUBS 0.231904f
C138 B.n101 VSUBS 0.184522f
C139 B.n102 VSUBS 0.008211f
C140 B.n103 VSUBS 0.008211f
C141 B.n104 VSUBS 0.008211f
C142 B.n105 VSUBS 0.008211f
C143 B.n106 VSUBS 0.004589f
C144 B.n107 VSUBS 0.008211f
C145 B.n108 VSUBS 0.008211f
C146 B.n109 VSUBS 0.008211f
C147 B.n110 VSUBS 0.008211f
C148 B.n111 VSUBS 0.008211f
C149 B.n112 VSUBS 0.008211f
C150 B.n113 VSUBS 0.008211f
C151 B.n114 VSUBS 0.008211f
C152 B.n115 VSUBS 0.008211f
C153 B.n116 VSUBS 0.008211f
C154 B.n117 VSUBS 0.008211f
C155 B.n118 VSUBS 0.020334f
C156 B.n119 VSUBS 0.008211f
C157 B.n120 VSUBS 0.008211f
C158 B.n121 VSUBS 0.008211f
C159 B.n122 VSUBS 0.008211f
C160 B.n123 VSUBS 0.008211f
C161 B.n124 VSUBS 0.008211f
C162 B.n125 VSUBS 0.008211f
C163 B.n126 VSUBS 0.008211f
C164 B.n127 VSUBS 0.008211f
C165 B.n128 VSUBS 0.008211f
C166 B.n129 VSUBS 0.008211f
C167 B.n130 VSUBS 0.008211f
C168 B.n131 VSUBS 0.008211f
C169 B.n132 VSUBS 0.008211f
C170 B.n133 VSUBS 0.008211f
C171 B.n134 VSUBS 0.008211f
C172 B.n135 VSUBS 0.008211f
C173 B.n136 VSUBS 0.008211f
C174 B.n137 VSUBS 0.008211f
C175 B.n138 VSUBS 0.008211f
C176 B.n139 VSUBS 0.008211f
C177 B.n140 VSUBS 0.008211f
C178 B.n141 VSUBS 0.008211f
C179 B.n142 VSUBS 0.008211f
C180 B.n143 VSUBS 0.008211f
C181 B.n144 VSUBS 0.008211f
C182 B.n145 VSUBS 0.008211f
C183 B.n146 VSUBS 0.008211f
C184 B.n147 VSUBS 0.008211f
C185 B.n148 VSUBS 0.008211f
C186 B.n149 VSUBS 0.008211f
C187 B.n150 VSUBS 0.008211f
C188 B.n151 VSUBS 0.008211f
C189 B.n152 VSUBS 0.008211f
C190 B.n153 VSUBS 0.008211f
C191 B.n154 VSUBS 0.008211f
C192 B.n155 VSUBS 0.008211f
C193 B.n156 VSUBS 0.008211f
C194 B.n157 VSUBS 0.008211f
C195 B.n158 VSUBS 0.008211f
C196 B.n159 VSUBS 0.008211f
C197 B.n160 VSUBS 0.008211f
C198 B.n161 VSUBS 0.008211f
C199 B.n162 VSUBS 0.008211f
C200 B.n163 VSUBS 0.008211f
C201 B.n164 VSUBS 0.008211f
C202 B.n165 VSUBS 0.008211f
C203 B.n166 VSUBS 0.008211f
C204 B.n167 VSUBS 0.008211f
C205 B.n168 VSUBS 0.008211f
C206 B.n169 VSUBS 0.008211f
C207 B.n170 VSUBS 0.008211f
C208 B.n171 VSUBS 0.008211f
C209 B.n172 VSUBS 0.008211f
C210 B.n173 VSUBS 0.008211f
C211 B.n174 VSUBS 0.008211f
C212 B.n175 VSUBS 0.008211f
C213 B.n176 VSUBS 0.008211f
C214 B.n177 VSUBS 0.008211f
C215 B.n178 VSUBS 0.008211f
C216 B.n179 VSUBS 0.008211f
C217 B.n180 VSUBS 0.008211f
C218 B.n181 VSUBS 0.008211f
C219 B.n182 VSUBS 0.008211f
C220 B.n183 VSUBS 0.018791f
C221 B.n184 VSUBS 0.018791f
C222 B.n185 VSUBS 0.020334f
C223 B.n186 VSUBS 0.008211f
C224 B.n187 VSUBS 0.008211f
C225 B.n188 VSUBS 0.008211f
C226 B.n189 VSUBS 0.008211f
C227 B.n190 VSUBS 0.008211f
C228 B.n191 VSUBS 0.008211f
C229 B.n192 VSUBS 0.008211f
C230 B.n193 VSUBS 0.008211f
C231 B.n194 VSUBS 0.008211f
C232 B.n195 VSUBS 0.008211f
C233 B.n196 VSUBS 0.008211f
C234 B.n197 VSUBS 0.008211f
C235 B.n198 VSUBS 0.008211f
C236 B.n199 VSUBS 0.008211f
C237 B.n200 VSUBS 0.008211f
C238 B.n201 VSUBS 0.008211f
C239 B.n202 VSUBS 0.008211f
C240 B.n203 VSUBS 0.008211f
C241 B.n204 VSUBS 0.008211f
C242 B.n205 VSUBS 0.008211f
C243 B.n206 VSUBS 0.008211f
C244 B.n207 VSUBS 0.008211f
C245 B.n208 VSUBS 0.008211f
C246 B.n209 VSUBS 0.008211f
C247 B.n210 VSUBS 0.008211f
C248 B.n211 VSUBS 0.008211f
C249 B.n212 VSUBS 0.008211f
C250 B.n213 VSUBS 0.008211f
C251 B.n214 VSUBS 0.008211f
C252 B.n215 VSUBS 0.008211f
C253 B.n216 VSUBS 0.008211f
C254 B.n217 VSUBS 0.008211f
C255 B.n218 VSUBS 0.008211f
C256 B.t5 VSUBS 0.105675f
C257 B.t4 VSUBS 0.136595f
C258 B.t3 VSUBS 0.901238f
C259 B.n219 VSUBS 0.231906f
C260 B.n220 VSUBS 0.184524f
C261 B.n221 VSUBS 0.019025f
C262 B.n222 VSUBS 0.007728f
C263 B.n223 VSUBS 0.008211f
C264 B.n224 VSUBS 0.008211f
C265 B.n225 VSUBS 0.008211f
C266 B.n226 VSUBS 0.008211f
C267 B.n227 VSUBS 0.008211f
C268 B.n228 VSUBS 0.008211f
C269 B.n229 VSUBS 0.008211f
C270 B.n230 VSUBS 0.008211f
C271 B.n231 VSUBS 0.008211f
C272 B.n232 VSUBS 0.008211f
C273 B.n233 VSUBS 0.008211f
C274 B.n234 VSUBS 0.008211f
C275 B.n235 VSUBS 0.008211f
C276 B.n236 VSUBS 0.008211f
C277 B.n237 VSUBS 0.008211f
C278 B.n238 VSUBS 0.004589f
C279 B.n239 VSUBS 0.019025f
C280 B.n240 VSUBS 0.007728f
C281 B.n241 VSUBS 0.008211f
C282 B.n242 VSUBS 0.008211f
C283 B.n243 VSUBS 0.008211f
C284 B.n244 VSUBS 0.008211f
C285 B.n245 VSUBS 0.008211f
C286 B.n246 VSUBS 0.008211f
C287 B.n247 VSUBS 0.008211f
C288 B.n248 VSUBS 0.008211f
C289 B.n249 VSUBS 0.008211f
C290 B.n250 VSUBS 0.008211f
C291 B.n251 VSUBS 0.008211f
C292 B.n252 VSUBS 0.008211f
C293 B.n253 VSUBS 0.008211f
C294 B.n254 VSUBS 0.008211f
C295 B.n255 VSUBS 0.008211f
C296 B.n256 VSUBS 0.008211f
C297 B.n257 VSUBS 0.008211f
C298 B.n258 VSUBS 0.008211f
C299 B.n259 VSUBS 0.008211f
C300 B.n260 VSUBS 0.008211f
C301 B.n261 VSUBS 0.008211f
C302 B.n262 VSUBS 0.008211f
C303 B.n263 VSUBS 0.008211f
C304 B.n264 VSUBS 0.008211f
C305 B.n265 VSUBS 0.008211f
C306 B.n266 VSUBS 0.008211f
C307 B.n267 VSUBS 0.008211f
C308 B.n268 VSUBS 0.008211f
C309 B.n269 VSUBS 0.008211f
C310 B.n270 VSUBS 0.008211f
C311 B.n271 VSUBS 0.008211f
C312 B.n272 VSUBS 0.008211f
C313 B.n273 VSUBS 0.008211f
C314 B.n274 VSUBS 0.020334f
C315 B.n275 VSUBS 0.01939f
C316 B.n276 VSUBS 0.019735f
C317 B.n277 VSUBS 0.008211f
C318 B.n278 VSUBS 0.008211f
C319 B.n279 VSUBS 0.008211f
C320 B.n280 VSUBS 0.008211f
C321 B.n281 VSUBS 0.008211f
C322 B.n282 VSUBS 0.008211f
C323 B.n283 VSUBS 0.008211f
C324 B.n284 VSUBS 0.008211f
C325 B.n285 VSUBS 0.008211f
C326 B.n286 VSUBS 0.008211f
C327 B.n287 VSUBS 0.008211f
C328 B.n288 VSUBS 0.008211f
C329 B.n289 VSUBS 0.008211f
C330 B.n290 VSUBS 0.008211f
C331 B.n291 VSUBS 0.008211f
C332 B.n292 VSUBS 0.008211f
C333 B.n293 VSUBS 0.008211f
C334 B.n294 VSUBS 0.008211f
C335 B.n295 VSUBS 0.008211f
C336 B.n296 VSUBS 0.008211f
C337 B.n297 VSUBS 0.008211f
C338 B.n298 VSUBS 0.008211f
C339 B.n299 VSUBS 0.008211f
C340 B.n300 VSUBS 0.008211f
C341 B.n301 VSUBS 0.008211f
C342 B.n302 VSUBS 0.008211f
C343 B.n303 VSUBS 0.008211f
C344 B.n304 VSUBS 0.008211f
C345 B.n305 VSUBS 0.008211f
C346 B.n306 VSUBS 0.008211f
C347 B.n307 VSUBS 0.008211f
C348 B.n308 VSUBS 0.008211f
C349 B.n309 VSUBS 0.008211f
C350 B.n310 VSUBS 0.008211f
C351 B.n311 VSUBS 0.008211f
C352 B.n312 VSUBS 0.008211f
C353 B.n313 VSUBS 0.008211f
C354 B.n314 VSUBS 0.008211f
C355 B.n315 VSUBS 0.008211f
C356 B.n316 VSUBS 0.008211f
C357 B.n317 VSUBS 0.008211f
C358 B.n318 VSUBS 0.008211f
C359 B.n319 VSUBS 0.008211f
C360 B.n320 VSUBS 0.008211f
C361 B.n321 VSUBS 0.008211f
C362 B.n322 VSUBS 0.008211f
C363 B.n323 VSUBS 0.008211f
C364 B.n324 VSUBS 0.008211f
C365 B.n325 VSUBS 0.008211f
C366 B.n326 VSUBS 0.008211f
C367 B.n327 VSUBS 0.008211f
C368 B.n328 VSUBS 0.008211f
C369 B.n329 VSUBS 0.008211f
C370 B.n330 VSUBS 0.008211f
C371 B.n331 VSUBS 0.008211f
C372 B.n332 VSUBS 0.008211f
C373 B.n333 VSUBS 0.008211f
C374 B.n334 VSUBS 0.008211f
C375 B.n335 VSUBS 0.008211f
C376 B.n336 VSUBS 0.008211f
C377 B.n337 VSUBS 0.008211f
C378 B.n338 VSUBS 0.008211f
C379 B.n339 VSUBS 0.008211f
C380 B.n340 VSUBS 0.008211f
C381 B.n341 VSUBS 0.008211f
C382 B.n342 VSUBS 0.008211f
C383 B.n343 VSUBS 0.008211f
C384 B.n344 VSUBS 0.008211f
C385 B.n345 VSUBS 0.008211f
C386 B.n346 VSUBS 0.008211f
C387 B.n347 VSUBS 0.008211f
C388 B.n348 VSUBS 0.008211f
C389 B.n349 VSUBS 0.008211f
C390 B.n350 VSUBS 0.008211f
C391 B.n351 VSUBS 0.008211f
C392 B.n352 VSUBS 0.008211f
C393 B.n353 VSUBS 0.008211f
C394 B.n354 VSUBS 0.008211f
C395 B.n355 VSUBS 0.008211f
C396 B.n356 VSUBS 0.008211f
C397 B.n357 VSUBS 0.008211f
C398 B.n358 VSUBS 0.008211f
C399 B.n359 VSUBS 0.008211f
C400 B.n360 VSUBS 0.008211f
C401 B.n361 VSUBS 0.008211f
C402 B.n362 VSUBS 0.008211f
C403 B.n363 VSUBS 0.008211f
C404 B.n364 VSUBS 0.008211f
C405 B.n365 VSUBS 0.008211f
C406 B.n366 VSUBS 0.008211f
C407 B.n367 VSUBS 0.008211f
C408 B.n368 VSUBS 0.008211f
C409 B.n369 VSUBS 0.008211f
C410 B.n370 VSUBS 0.008211f
C411 B.n371 VSUBS 0.008211f
C412 B.n372 VSUBS 0.008211f
C413 B.n373 VSUBS 0.008211f
C414 B.n374 VSUBS 0.008211f
C415 B.n375 VSUBS 0.008211f
C416 B.n376 VSUBS 0.008211f
C417 B.n377 VSUBS 0.008211f
C418 B.n378 VSUBS 0.008211f
C419 B.n379 VSUBS 0.018791f
C420 B.n380 VSUBS 0.018791f
C421 B.n381 VSUBS 0.020334f
C422 B.n382 VSUBS 0.008211f
C423 B.n383 VSUBS 0.008211f
C424 B.n384 VSUBS 0.008211f
C425 B.n385 VSUBS 0.008211f
C426 B.n386 VSUBS 0.008211f
C427 B.n387 VSUBS 0.008211f
C428 B.n388 VSUBS 0.008211f
C429 B.n389 VSUBS 0.008211f
C430 B.n390 VSUBS 0.008211f
C431 B.n391 VSUBS 0.008211f
C432 B.n392 VSUBS 0.008211f
C433 B.n393 VSUBS 0.008211f
C434 B.n394 VSUBS 0.008211f
C435 B.n395 VSUBS 0.008211f
C436 B.n396 VSUBS 0.008211f
C437 B.n397 VSUBS 0.008211f
C438 B.n398 VSUBS 0.008211f
C439 B.n399 VSUBS 0.008211f
C440 B.n400 VSUBS 0.008211f
C441 B.n401 VSUBS 0.008211f
C442 B.n402 VSUBS 0.008211f
C443 B.n403 VSUBS 0.008211f
C444 B.n404 VSUBS 0.008211f
C445 B.n405 VSUBS 0.008211f
C446 B.n406 VSUBS 0.008211f
C447 B.n407 VSUBS 0.008211f
C448 B.n408 VSUBS 0.008211f
C449 B.n409 VSUBS 0.008211f
C450 B.n410 VSUBS 0.008211f
C451 B.n411 VSUBS 0.008211f
C452 B.n412 VSUBS 0.008211f
C453 B.n413 VSUBS 0.008211f
C454 B.n414 VSUBS 0.008211f
C455 B.n415 VSUBS 0.007728f
C456 B.n416 VSUBS 0.008211f
C457 B.n417 VSUBS 0.008211f
C458 B.n418 VSUBS 0.004589f
C459 B.n419 VSUBS 0.008211f
C460 B.n420 VSUBS 0.008211f
C461 B.n421 VSUBS 0.008211f
C462 B.n422 VSUBS 0.008211f
C463 B.n423 VSUBS 0.008211f
C464 B.n424 VSUBS 0.008211f
C465 B.n425 VSUBS 0.008211f
C466 B.n426 VSUBS 0.008211f
C467 B.n427 VSUBS 0.008211f
C468 B.n428 VSUBS 0.008211f
C469 B.n429 VSUBS 0.008211f
C470 B.n430 VSUBS 0.008211f
C471 B.n431 VSUBS 0.004589f
C472 B.n432 VSUBS 0.019025f
C473 B.n433 VSUBS 0.007728f
C474 B.n434 VSUBS 0.008211f
C475 B.n435 VSUBS 0.008211f
C476 B.n436 VSUBS 0.008211f
C477 B.n437 VSUBS 0.008211f
C478 B.n438 VSUBS 0.008211f
C479 B.n439 VSUBS 0.008211f
C480 B.n440 VSUBS 0.008211f
C481 B.n441 VSUBS 0.008211f
C482 B.n442 VSUBS 0.008211f
C483 B.n443 VSUBS 0.008211f
C484 B.n444 VSUBS 0.008211f
C485 B.n445 VSUBS 0.008211f
C486 B.n446 VSUBS 0.008211f
C487 B.n447 VSUBS 0.008211f
C488 B.n448 VSUBS 0.008211f
C489 B.n449 VSUBS 0.008211f
C490 B.n450 VSUBS 0.008211f
C491 B.n451 VSUBS 0.008211f
C492 B.n452 VSUBS 0.008211f
C493 B.n453 VSUBS 0.008211f
C494 B.n454 VSUBS 0.008211f
C495 B.n455 VSUBS 0.008211f
C496 B.n456 VSUBS 0.008211f
C497 B.n457 VSUBS 0.008211f
C498 B.n458 VSUBS 0.008211f
C499 B.n459 VSUBS 0.008211f
C500 B.n460 VSUBS 0.008211f
C501 B.n461 VSUBS 0.008211f
C502 B.n462 VSUBS 0.008211f
C503 B.n463 VSUBS 0.008211f
C504 B.n464 VSUBS 0.008211f
C505 B.n465 VSUBS 0.008211f
C506 B.n466 VSUBS 0.008211f
C507 B.n467 VSUBS 0.008211f
C508 B.n468 VSUBS 0.020334f
C509 B.n469 VSUBS 0.018791f
C510 B.n470 VSUBS 0.018791f
C511 B.n471 VSUBS 0.008211f
C512 B.n472 VSUBS 0.008211f
C513 B.n473 VSUBS 0.008211f
C514 B.n474 VSUBS 0.008211f
C515 B.n475 VSUBS 0.008211f
C516 B.n476 VSUBS 0.008211f
C517 B.n477 VSUBS 0.008211f
C518 B.n478 VSUBS 0.008211f
C519 B.n479 VSUBS 0.008211f
C520 B.n480 VSUBS 0.008211f
C521 B.n481 VSUBS 0.008211f
C522 B.n482 VSUBS 0.008211f
C523 B.n483 VSUBS 0.008211f
C524 B.n484 VSUBS 0.008211f
C525 B.n485 VSUBS 0.008211f
C526 B.n486 VSUBS 0.008211f
C527 B.n487 VSUBS 0.008211f
C528 B.n488 VSUBS 0.008211f
C529 B.n489 VSUBS 0.008211f
C530 B.n490 VSUBS 0.008211f
C531 B.n491 VSUBS 0.008211f
C532 B.n492 VSUBS 0.008211f
C533 B.n493 VSUBS 0.008211f
C534 B.n494 VSUBS 0.008211f
C535 B.n495 VSUBS 0.008211f
C536 B.n496 VSUBS 0.008211f
C537 B.n497 VSUBS 0.008211f
C538 B.n498 VSUBS 0.008211f
C539 B.n499 VSUBS 0.008211f
C540 B.n500 VSUBS 0.008211f
C541 B.n501 VSUBS 0.008211f
C542 B.n502 VSUBS 0.008211f
C543 B.n503 VSUBS 0.008211f
C544 B.n504 VSUBS 0.008211f
C545 B.n505 VSUBS 0.008211f
C546 B.n506 VSUBS 0.008211f
C547 B.n507 VSUBS 0.008211f
C548 B.n508 VSUBS 0.008211f
C549 B.n509 VSUBS 0.008211f
C550 B.n510 VSUBS 0.008211f
C551 B.n511 VSUBS 0.008211f
C552 B.n512 VSUBS 0.008211f
C553 B.n513 VSUBS 0.008211f
C554 B.n514 VSUBS 0.008211f
C555 B.n515 VSUBS 0.008211f
C556 B.n516 VSUBS 0.008211f
C557 B.n517 VSUBS 0.008211f
C558 B.n518 VSUBS 0.008211f
C559 B.n519 VSUBS 0.010715f
C560 B.n520 VSUBS 0.011415f
C561 B.n521 VSUBS 0.022699f
C562 VDD1.t1 VSUBS 0.133002f
C563 VDD1.t3 VSUBS 0.133002f
C564 VDD1.n0 VSUBS 0.883497f
C565 VDD1.t0 VSUBS 0.133002f
C566 VDD1.t2 VSUBS 0.133002f
C567 VDD1.n1 VSUBS 1.34568f
C568 VP.n0 VSUBS 0.055648f
C569 VP.t1 VSUBS 1.81266f
C570 VP.n1 VSUBS 0.08389f
C571 VP.n2 VSUBS 0.042209f
C572 VP.n3 VSUBS 0.040605f
C573 VP.t0 VSUBS 2.17388f
C574 VP.t2 VSUBS 2.18322f
C575 VP.n4 VSUBS 3.40438f
C576 VP.t3 VSUBS 1.81266f
C577 VP.n5 VSUBS 0.803904f
C578 VP.n6 VSUBS 2.01878f
C579 VP.n7 VSUBS 0.055648f
C580 VP.n8 VSUBS 0.042209f
C581 VP.n9 VSUBS 0.078667f
C582 VP.n10 VSUBS 0.08389f
C583 VP.n11 VSUBS 0.034122f
C584 VP.n12 VSUBS 0.042209f
C585 VP.n13 VSUBS 0.042209f
C586 VP.n14 VSUBS 0.042209f
C587 VP.n15 VSUBS 0.078667f
C588 VP.n16 VSUBS 0.040605f
C589 VP.n17 VSUBS 0.803904f
C590 VP.n18 VSUBS 0.078758f
C591 VDD2.t2 VSUBS 0.133063f
C592 VDD2.t3 VSUBS 0.133063f
C593 VDD2.n0 VSUBS 1.32572f
C594 VDD2.t1 VSUBS 0.133063f
C595 VDD2.t0 VSUBS 0.133063f
C596 VDD2.n1 VSUBS 0.883464f
C597 VDD2.n2 VSUBS 3.7183f
C598 VTAIL.n0 VSUBS 0.030662f
C599 VTAIL.n1 VSUBS 0.02769f
C600 VTAIL.n2 VSUBS 0.014879f
C601 VTAIL.n3 VSUBS 0.035169f
C602 VTAIL.n4 VSUBS 0.015755f
C603 VTAIL.n5 VSUBS 0.02769f
C604 VTAIL.n6 VSUBS 0.014879f
C605 VTAIL.n7 VSUBS 0.035169f
C606 VTAIL.n8 VSUBS 0.015755f
C607 VTAIL.n9 VSUBS 0.12272f
C608 VTAIL.t6 VSUBS 0.075511f
C609 VTAIL.n10 VSUBS 0.026377f
C610 VTAIL.n11 VSUBS 0.022361f
C611 VTAIL.n12 VSUBS 0.014879f
C612 VTAIL.n13 VSUBS 0.638867f
C613 VTAIL.n14 VSUBS 0.02769f
C614 VTAIL.n15 VSUBS 0.014879f
C615 VTAIL.n16 VSUBS 0.015755f
C616 VTAIL.n17 VSUBS 0.035169f
C617 VTAIL.n18 VSUBS 0.035169f
C618 VTAIL.n19 VSUBS 0.015755f
C619 VTAIL.n20 VSUBS 0.014879f
C620 VTAIL.n21 VSUBS 0.02769f
C621 VTAIL.n22 VSUBS 0.02769f
C622 VTAIL.n23 VSUBS 0.014879f
C623 VTAIL.n24 VSUBS 0.015755f
C624 VTAIL.n25 VSUBS 0.035169f
C625 VTAIL.n26 VSUBS 0.085946f
C626 VTAIL.n27 VSUBS 0.015755f
C627 VTAIL.n28 VSUBS 0.014879f
C628 VTAIL.n29 VSUBS 0.065138f
C629 VTAIL.n30 VSUBS 0.043292f
C630 VTAIL.n31 VSUBS 0.187544f
C631 VTAIL.n32 VSUBS 0.030662f
C632 VTAIL.n33 VSUBS 0.02769f
C633 VTAIL.n34 VSUBS 0.014879f
C634 VTAIL.n35 VSUBS 0.035169f
C635 VTAIL.n36 VSUBS 0.015755f
C636 VTAIL.n37 VSUBS 0.02769f
C637 VTAIL.n38 VSUBS 0.014879f
C638 VTAIL.n39 VSUBS 0.035169f
C639 VTAIL.n40 VSUBS 0.015755f
C640 VTAIL.n41 VSUBS 0.12272f
C641 VTAIL.t0 VSUBS 0.075511f
C642 VTAIL.n42 VSUBS 0.026377f
C643 VTAIL.n43 VSUBS 0.022361f
C644 VTAIL.n44 VSUBS 0.014879f
C645 VTAIL.n45 VSUBS 0.638867f
C646 VTAIL.n46 VSUBS 0.02769f
C647 VTAIL.n47 VSUBS 0.014879f
C648 VTAIL.n48 VSUBS 0.015755f
C649 VTAIL.n49 VSUBS 0.035169f
C650 VTAIL.n50 VSUBS 0.035169f
C651 VTAIL.n51 VSUBS 0.015755f
C652 VTAIL.n52 VSUBS 0.014879f
C653 VTAIL.n53 VSUBS 0.02769f
C654 VTAIL.n54 VSUBS 0.02769f
C655 VTAIL.n55 VSUBS 0.014879f
C656 VTAIL.n56 VSUBS 0.015755f
C657 VTAIL.n57 VSUBS 0.035169f
C658 VTAIL.n58 VSUBS 0.085946f
C659 VTAIL.n59 VSUBS 0.015755f
C660 VTAIL.n60 VSUBS 0.014879f
C661 VTAIL.n61 VSUBS 0.065138f
C662 VTAIL.n62 VSUBS 0.043292f
C663 VTAIL.n63 VSUBS 0.298496f
C664 VTAIL.n64 VSUBS 0.030662f
C665 VTAIL.n65 VSUBS 0.02769f
C666 VTAIL.n66 VSUBS 0.014879f
C667 VTAIL.n67 VSUBS 0.035169f
C668 VTAIL.n68 VSUBS 0.015755f
C669 VTAIL.n69 VSUBS 0.02769f
C670 VTAIL.n70 VSUBS 0.014879f
C671 VTAIL.n71 VSUBS 0.035169f
C672 VTAIL.n72 VSUBS 0.015755f
C673 VTAIL.n73 VSUBS 0.12272f
C674 VTAIL.t1 VSUBS 0.075511f
C675 VTAIL.n74 VSUBS 0.026377f
C676 VTAIL.n75 VSUBS 0.022361f
C677 VTAIL.n76 VSUBS 0.014879f
C678 VTAIL.n77 VSUBS 0.638867f
C679 VTAIL.n78 VSUBS 0.02769f
C680 VTAIL.n79 VSUBS 0.014879f
C681 VTAIL.n80 VSUBS 0.015755f
C682 VTAIL.n81 VSUBS 0.035169f
C683 VTAIL.n82 VSUBS 0.035169f
C684 VTAIL.n83 VSUBS 0.015755f
C685 VTAIL.n84 VSUBS 0.014879f
C686 VTAIL.n85 VSUBS 0.02769f
C687 VTAIL.n86 VSUBS 0.02769f
C688 VTAIL.n87 VSUBS 0.014879f
C689 VTAIL.n88 VSUBS 0.015755f
C690 VTAIL.n89 VSUBS 0.035169f
C691 VTAIL.n90 VSUBS 0.085946f
C692 VTAIL.n91 VSUBS 0.015755f
C693 VTAIL.n92 VSUBS 0.014879f
C694 VTAIL.n93 VSUBS 0.065138f
C695 VTAIL.n94 VSUBS 0.043292f
C696 VTAIL.n95 VSUBS 1.3288f
C697 VTAIL.n96 VSUBS 0.030662f
C698 VTAIL.n97 VSUBS 0.02769f
C699 VTAIL.n98 VSUBS 0.014879f
C700 VTAIL.n99 VSUBS 0.035169f
C701 VTAIL.n100 VSUBS 0.015755f
C702 VTAIL.n101 VSUBS 0.02769f
C703 VTAIL.n102 VSUBS 0.014879f
C704 VTAIL.n103 VSUBS 0.035169f
C705 VTAIL.n104 VSUBS 0.015755f
C706 VTAIL.n105 VSUBS 0.12272f
C707 VTAIL.t5 VSUBS 0.075511f
C708 VTAIL.n106 VSUBS 0.026377f
C709 VTAIL.n107 VSUBS 0.022361f
C710 VTAIL.n108 VSUBS 0.014879f
C711 VTAIL.n109 VSUBS 0.638867f
C712 VTAIL.n110 VSUBS 0.02769f
C713 VTAIL.n111 VSUBS 0.014879f
C714 VTAIL.n112 VSUBS 0.015755f
C715 VTAIL.n113 VSUBS 0.035169f
C716 VTAIL.n114 VSUBS 0.035169f
C717 VTAIL.n115 VSUBS 0.015755f
C718 VTAIL.n116 VSUBS 0.014879f
C719 VTAIL.n117 VSUBS 0.02769f
C720 VTAIL.n118 VSUBS 0.02769f
C721 VTAIL.n119 VSUBS 0.014879f
C722 VTAIL.n120 VSUBS 0.015755f
C723 VTAIL.n121 VSUBS 0.035169f
C724 VTAIL.n122 VSUBS 0.085946f
C725 VTAIL.n123 VSUBS 0.015755f
C726 VTAIL.n124 VSUBS 0.014879f
C727 VTAIL.n125 VSUBS 0.065138f
C728 VTAIL.n126 VSUBS 0.043292f
C729 VTAIL.n127 VSUBS 1.3288f
C730 VTAIL.n128 VSUBS 0.030662f
C731 VTAIL.n129 VSUBS 0.02769f
C732 VTAIL.n130 VSUBS 0.014879f
C733 VTAIL.n131 VSUBS 0.035169f
C734 VTAIL.n132 VSUBS 0.015755f
C735 VTAIL.n133 VSUBS 0.02769f
C736 VTAIL.n134 VSUBS 0.014879f
C737 VTAIL.n135 VSUBS 0.035169f
C738 VTAIL.n136 VSUBS 0.015755f
C739 VTAIL.n137 VSUBS 0.12272f
C740 VTAIL.t4 VSUBS 0.075511f
C741 VTAIL.n138 VSUBS 0.026377f
C742 VTAIL.n139 VSUBS 0.022361f
C743 VTAIL.n140 VSUBS 0.014879f
C744 VTAIL.n141 VSUBS 0.638867f
C745 VTAIL.n142 VSUBS 0.02769f
C746 VTAIL.n143 VSUBS 0.014879f
C747 VTAIL.n144 VSUBS 0.015755f
C748 VTAIL.n145 VSUBS 0.035169f
C749 VTAIL.n146 VSUBS 0.035169f
C750 VTAIL.n147 VSUBS 0.015755f
C751 VTAIL.n148 VSUBS 0.014879f
C752 VTAIL.n149 VSUBS 0.02769f
C753 VTAIL.n150 VSUBS 0.02769f
C754 VTAIL.n151 VSUBS 0.014879f
C755 VTAIL.n152 VSUBS 0.015755f
C756 VTAIL.n153 VSUBS 0.035169f
C757 VTAIL.n154 VSUBS 0.085946f
C758 VTAIL.n155 VSUBS 0.015755f
C759 VTAIL.n156 VSUBS 0.014879f
C760 VTAIL.n157 VSUBS 0.065138f
C761 VTAIL.n158 VSUBS 0.043292f
C762 VTAIL.n159 VSUBS 0.298496f
C763 VTAIL.n160 VSUBS 0.030662f
C764 VTAIL.n161 VSUBS 0.02769f
C765 VTAIL.n162 VSUBS 0.014879f
C766 VTAIL.n163 VSUBS 0.035169f
C767 VTAIL.n164 VSUBS 0.015755f
C768 VTAIL.n165 VSUBS 0.02769f
C769 VTAIL.n166 VSUBS 0.014879f
C770 VTAIL.n167 VSUBS 0.035169f
C771 VTAIL.n168 VSUBS 0.015755f
C772 VTAIL.n169 VSUBS 0.12272f
C773 VTAIL.t2 VSUBS 0.075511f
C774 VTAIL.n170 VSUBS 0.026377f
C775 VTAIL.n171 VSUBS 0.022361f
C776 VTAIL.n172 VSUBS 0.014879f
C777 VTAIL.n173 VSUBS 0.638867f
C778 VTAIL.n174 VSUBS 0.02769f
C779 VTAIL.n175 VSUBS 0.014879f
C780 VTAIL.n176 VSUBS 0.015755f
C781 VTAIL.n177 VSUBS 0.035169f
C782 VTAIL.n178 VSUBS 0.035169f
C783 VTAIL.n179 VSUBS 0.015755f
C784 VTAIL.n180 VSUBS 0.014879f
C785 VTAIL.n181 VSUBS 0.02769f
C786 VTAIL.n182 VSUBS 0.02769f
C787 VTAIL.n183 VSUBS 0.014879f
C788 VTAIL.n184 VSUBS 0.015755f
C789 VTAIL.n185 VSUBS 0.035169f
C790 VTAIL.n186 VSUBS 0.085946f
C791 VTAIL.n187 VSUBS 0.015755f
C792 VTAIL.n188 VSUBS 0.014879f
C793 VTAIL.n189 VSUBS 0.065138f
C794 VTAIL.n190 VSUBS 0.043292f
C795 VTAIL.n191 VSUBS 0.298496f
C796 VTAIL.n192 VSUBS 0.030662f
C797 VTAIL.n193 VSUBS 0.02769f
C798 VTAIL.n194 VSUBS 0.014879f
C799 VTAIL.n195 VSUBS 0.035169f
C800 VTAIL.n196 VSUBS 0.015755f
C801 VTAIL.n197 VSUBS 0.02769f
C802 VTAIL.n198 VSUBS 0.014879f
C803 VTAIL.n199 VSUBS 0.035169f
C804 VTAIL.n200 VSUBS 0.015755f
C805 VTAIL.n201 VSUBS 0.12272f
C806 VTAIL.t3 VSUBS 0.075511f
C807 VTAIL.n202 VSUBS 0.026377f
C808 VTAIL.n203 VSUBS 0.022361f
C809 VTAIL.n204 VSUBS 0.014879f
C810 VTAIL.n205 VSUBS 0.638867f
C811 VTAIL.n206 VSUBS 0.02769f
C812 VTAIL.n207 VSUBS 0.014879f
C813 VTAIL.n208 VSUBS 0.015755f
C814 VTAIL.n209 VSUBS 0.035169f
C815 VTAIL.n210 VSUBS 0.035169f
C816 VTAIL.n211 VSUBS 0.015755f
C817 VTAIL.n212 VSUBS 0.014879f
C818 VTAIL.n213 VSUBS 0.02769f
C819 VTAIL.n214 VSUBS 0.02769f
C820 VTAIL.n215 VSUBS 0.014879f
C821 VTAIL.n216 VSUBS 0.015755f
C822 VTAIL.n217 VSUBS 0.035169f
C823 VTAIL.n218 VSUBS 0.085946f
C824 VTAIL.n219 VSUBS 0.015755f
C825 VTAIL.n220 VSUBS 0.014879f
C826 VTAIL.n221 VSUBS 0.065138f
C827 VTAIL.n222 VSUBS 0.043292f
C828 VTAIL.n223 VSUBS 1.3288f
C829 VTAIL.n224 VSUBS 0.030662f
C830 VTAIL.n225 VSUBS 0.02769f
C831 VTAIL.n226 VSUBS 0.014879f
C832 VTAIL.n227 VSUBS 0.035169f
C833 VTAIL.n228 VSUBS 0.015755f
C834 VTAIL.n229 VSUBS 0.02769f
C835 VTAIL.n230 VSUBS 0.014879f
C836 VTAIL.n231 VSUBS 0.035169f
C837 VTAIL.n232 VSUBS 0.015755f
C838 VTAIL.n233 VSUBS 0.12272f
C839 VTAIL.t7 VSUBS 0.075511f
C840 VTAIL.n234 VSUBS 0.026377f
C841 VTAIL.n235 VSUBS 0.022361f
C842 VTAIL.n236 VSUBS 0.014879f
C843 VTAIL.n237 VSUBS 0.638867f
C844 VTAIL.n238 VSUBS 0.02769f
C845 VTAIL.n239 VSUBS 0.014879f
C846 VTAIL.n240 VSUBS 0.015755f
C847 VTAIL.n241 VSUBS 0.035169f
C848 VTAIL.n242 VSUBS 0.035169f
C849 VTAIL.n243 VSUBS 0.015755f
C850 VTAIL.n244 VSUBS 0.014879f
C851 VTAIL.n245 VSUBS 0.02769f
C852 VTAIL.n246 VSUBS 0.02769f
C853 VTAIL.n247 VSUBS 0.014879f
C854 VTAIL.n248 VSUBS 0.015755f
C855 VTAIL.n249 VSUBS 0.035169f
C856 VTAIL.n250 VSUBS 0.085946f
C857 VTAIL.n251 VSUBS 0.015755f
C858 VTAIL.n252 VSUBS 0.014879f
C859 VTAIL.n253 VSUBS 0.065138f
C860 VTAIL.n254 VSUBS 0.043292f
C861 VTAIL.n255 VSUBS 1.20747f
C862 VN.t1 VSUBS 2.09302f
C863 VN.t0 VSUBS 2.08407f
C864 VN.n0 VSUBS 1.32402f
C865 VN.t3 VSUBS 2.09302f
C866 VN.t2 VSUBS 2.08407f
C867 VN.n1 VSUBS 3.28541f
.ends

