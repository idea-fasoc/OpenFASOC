* NGSPICE file created from diff_pair_sample_1659.ext - technology: sky130A

.subckt diff_pair_sample_1659 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t1 VN.t0 VTAIL.t2 B.t0 sky130_fd_pr__nfet_01v8 ad=2.7651 pd=14.96 as=2.7651 ps=14.96 w=7.09 l=0.35
X1 B.t15 B.t13 B.t14 B.t10 sky130_fd_pr__nfet_01v8 ad=2.7651 pd=14.96 as=0 ps=0 w=7.09 l=0.35
X2 VDD1.t1 VP.t0 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=2.7651 pd=14.96 as=2.7651 ps=14.96 w=7.09 l=0.35
X3 B.t12 B.t9 B.t11 B.t10 sky130_fd_pr__nfet_01v8 ad=2.7651 pd=14.96 as=0 ps=0 w=7.09 l=0.35
X4 VDD2.t0 VN.t1 VTAIL.t3 B.t1 sky130_fd_pr__nfet_01v8 ad=2.7651 pd=14.96 as=2.7651 ps=14.96 w=7.09 l=0.35
X5 VDD1.t0 VP.t1 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=2.7651 pd=14.96 as=2.7651 ps=14.96 w=7.09 l=0.35
X6 B.t8 B.t6 B.t7 B.t3 sky130_fd_pr__nfet_01v8 ad=2.7651 pd=14.96 as=0 ps=0 w=7.09 l=0.35
X7 B.t5 B.t2 B.t4 B.t3 sky130_fd_pr__nfet_01v8 ad=2.7651 pd=14.96 as=0 ps=0 w=7.09 l=0.35
R0 VN VN.t0 797.788
R1 VN VN.t1 762.475
R2 VTAIL.n1 VTAIL.t2 51.9191
R3 VTAIL.n2 VTAIL.t1 51.9188
R4 VTAIL.n3 VTAIL.t3 51.9188
R5 VTAIL.n0 VTAIL.t0 51.9188
R6 VTAIL.n1 VTAIL.n0 19.6686
R7 VTAIL.n3 VTAIL.n2 19.0824
R8 VTAIL.n2 VTAIL.n1 0.763431
R9 VTAIL VTAIL.n0 0.675069
R10 VTAIL VTAIL.n3 0.0888621
R11 VDD2.n0 VDD2.t0 99.5588
R12 VDD2.n0 VDD2.t1 68.5976
R13 VDD2 VDD2.n0 0.205241
R14 B.n224 B.t13 699.769
R15 B.n233 B.t9 699.769
R16 B.n61 B.t6 699.769
R17 B.n59 B.t2 699.769
R18 B.n428 B.n427 585
R19 B.n187 B.n58 585
R20 B.n186 B.n185 585
R21 B.n184 B.n183 585
R22 B.n182 B.n181 585
R23 B.n180 B.n179 585
R24 B.n178 B.n177 585
R25 B.n176 B.n175 585
R26 B.n174 B.n173 585
R27 B.n172 B.n171 585
R28 B.n170 B.n169 585
R29 B.n168 B.n167 585
R30 B.n166 B.n165 585
R31 B.n164 B.n163 585
R32 B.n162 B.n161 585
R33 B.n160 B.n159 585
R34 B.n158 B.n157 585
R35 B.n156 B.n155 585
R36 B.n154 B.n153 585
R37 B.n152 B.n151 585
R38 B.n150 B.n149 585
R39 B.n148 B.n147 585
R40 B.n146 B.n145 585
R41 B.n144 B.n143 585
R42 B.n142 B.n141 585
R43 B.n140 B.n139 585
R44 B.n138 B.n137 585
R45 B.n135 B.n134 585
R46 B.n133 B.n132 585
R47 B.n131 B.n130 585
R48 B.n129 B.n128 585
R49 B.n127 B.n126 585
R50 B.n125 B.n124 585
R51 B.n123 B.n122 585
R52 B.n121 B.n120 585
R53 B.n119 B.n118 585
R54 B.n117 B.n116 585
R55 B.n114 B.n113 585
R56 B.n112 B.n111 585
R57 B.n110 B.n109 585
R58 B.n108 B.n107 585
R59 B.n106 B.n105 585
R60 B.n104 B.n103 585
R61 B.n102 B.n101 585
R62 B.n100 B.n99 585
R63 B.n98 B.n97 585
R64 B.n96 B.n95 585
R65 B.n94 B.n93 585
R66 B.n92 B.n91 585
R67 B.n90 B.n89 585
R68 B.n88 B.n87 585
R69 B.n86 B.n85 585
R70 B.n84 B.n83 585
R71 B.n82 B.n81 585
R72 B.n80 B.n79 585
R73 B.n78 B.n77 585
R74 B.n76 B.n75 585
R75 B.n74 B.n73 585
R76 B.n72 B.n71 585
R77 B.n70 B.n69 585
R78 B.n68 B.n67 585
R79 B.n66 B.n65 585
R80 B.n64 B.n63 585
R81 B.n25 B.n24 585
R82 B.n426 B.n26 585
R83 B.n431 B.n26 585
R84 B.n425 B.n424 585
R85 B.n424 B.n22 585
R86 B.n423 B.n21 585
R87 B.n437 B.n21 585
R88 B.n422 B.n20 585
R89 B.n438 B.n20 585
R90 B.n421 B.n19 585
R91 B.n439 B.n19 585
R92 B.n420 B.n419 585
R93 B.n419 B.n15 585
R94 B.n418 B.n14 585
R95 B.n445 B.n14 585
R96 B.n417 B.n13 585
R97 B.n446 B.n13 585
R98 B.n416 B.n12 585
R99 B.n447 B.n12 585
R100 B.n415 B.n414 585
R101 B.n414 B.n11 585
R102 B.n413 B.n7 585
R103 B.n453 B.n7 585
R104 B.n412 B.n6 585
R105 B.n454 B.n6 585
R106 B.n411 B.n5 585
R107 B.n455 B.n5 585
R108 B.n410 B.n409 585
R109 B.n409 B.n4 585
R110 B.n408 B.n188 585
R111 B.n408 B.n407 585
R112 B.n397 B.n189 585
R113 B.n400 B.n189 585
R114 B.n399 B.n398 585
R115 B.n401 B.n399 585
R116 B.n396 B.n194 585
R117 B.n194 B.n193 585
R118 B.n395 B.n394 585
R119 B.n394 B.n393 585
R120 B.n196 B.n195 585
R121 B.n197 B.n196 585
R122 B.n386 B.n385 585
R123 B.n387 B.n386 585
R124 B.n384 B.n202 585
R125 B.n202 B.n201 585
R126 B.n383 B.n382 585
R127 B.n382 B.n381 585
R128 B.n204 B.n203 585
R129 B.n205 B.n204 585
R130 B.n374 B.n373 585
R131 B.n375 B.n374 585
R132 B.n208 B.n207 585
R133 B.n249 B.n248 585
R134 B.n250 B.n246 585
R135 B.n246 B.n209 585
R136 B.n252 B.n251 585
R137 B.n254 B.n245 585
R138 B.n257 B.n256 585
R139 B.n258 B.n244 585
R140 B.n260 B.n259 585
R141 B.n262 B.n243 585
R142 B.n265 B.n264 585
R143 B.n266 B.n242 585
R144 B.n268 B.n267 585
R145 B.n270 B.n241 585
R146 B.n273 B.n272 585
R147 B.n274 B.n240 585
R148 B.n276 B.n275 585
R149 B.n278 B.n239 585
R150 B.n281 B.n280 585
R151 B.n282 B.n238 585
R152 B.n284 B.n283 585
R153 B.n286 B.n237 585
R154 B.n289 B.n288 585
R155 B.n290 B.n236 585
R156 B.n292 B.n291 585
R157 B.n294 B.n235 585
R158 B.n297 B.n296 585
R159 B.n298 B.n232 585
R160 B.n301 B.n300 585
R161 B.n303 B.n231 585
R162 B.n306 B.n305 585
R163 B.n307 B.n230 585
R164 B.n309 B.n308 585
R165 B.n311 B.n229 585
R166 B.n314 B.n313 585
R167 B.n315 B.n228 585
R168 B.n317 B.n316 585
R169 B.n319 B.n227 585
R170 B.n322 B.n321 585
R171 B.n323 B.n223 585
R172 B.n325 B.n324 585
R173 B.n327 B.n222 585
R174 B.n330 B.n329 585
R175 B.n331 B.n221 585
R176 B.n333 B.n332 585
R177 B.n335 B.n220 585
R178 B.n338 B.n337 585
R179 B.n339 B.n219 585
R180 B.n341 B.n340 585
R181 B.n343 B.n218 585
R182 B.n346 B.n345 585
R183 B.n347 B.n217 585
R184 B.n349 B.n348 585
R185 B.n351 B.n216 585
R186 B.n354 B.n353 585
R187 B.n355 B.n215 585
R188 B.n357 B.n356 585
R189 B.n359 B.n214 585
R190 B.n362 B.n361 585
R191 B.n363 B.n213 585
R192 B.n365 B.n364 585
R193 B.n367 B.n212 585
R194 B.n368 B.n211 585
R195 B.n371 B.n370 585
R196 B.n372 B.n210 585
R197 B.n210 B.n209 585
R198 B.n377 B.n376 585
R199 B.n376 B.n375 585
R200 B.n378 B.n206 585
R201 B.n206 B.n205 585
R202 B.n380 B.n379 585
R203 B.n381 B.n380 585
R204 B.n200 B.n199 585
R205 B.n201 B.n200 585
R206 B.n389 B.n388 585
R207 B.n388 B.n387 585
R208 B.n390 B.n198 585
R209 B.n198 B.n197 585
R210 B.n392 B.n391 585
R211 B.n393 B.n392 585
R212 B.n192 B.n191 585
R213 B.n193 B.n192 585
R214 B.n403 B.n402 585
R215 B.n402 B.n401 585
R216 B.n404 B.n190 585
R217 B.n400 B.n190 585
R218 B.n406 B.n405 585
R219 B.n407 B.n406 585
R220 B.n2 B.n0 585
R221 B.n4 B.n2 585
R222 B.n3 B.n1 585
R223 B.n454 B.n3 585
R224 B.n452 B.n451 585
R225 B.n453 B.n452 585
R226 B.n450 B.n8 585
R227 B.n11 B.n8 585
R228 B.n449 B.n448 585
R229 B.n448 B.n447 585
R230 B.n10 B.n9 585
R231 B.n446 B.n10 585
R232 B.n444 B.n443 585
R233 B.n445 B.n444 585
R234 B.n442 B.n16 585
R235 B.n16 B.n15 585
R236 B.n441 B.n440 585
R237 B.n440 B.n439 585
R238 B.n18 B.n17 585
R239 B.n438 B.n18 585
R240 B.n436 B.n435 585
R241 B.n437 B.n436 585
R242 B.n434 B.n23 585
R243 B.n23 B.n22 585
R244 B.n433 B.n432 585
R245 B.n432 B.n431 585
R246 B.n457 B.n456 585
R247 B.n456 B.n455 585
R248 B.n376 B.n208 521.33
R249 B.n432 B.n25 521.33
R250 B.n374 B.n210 521.33
R251 B.n428 B.n26 521.33
R252 B.n430 B.n429 256.663
R253 B.n430 B.n57 256.663
R254 B.n430 B.n56 256.663
R255 B.n430 B.n55 256.663
R256 B.n430 B.n54 256.663
R257 B.n430 B.n53 256.663
R258 B.n430 B.n52 256.663
R259 B.n430 B.n51 256.663
R260 B.n430 B.n50 256.663
R261 B.n430 B.n49 256.663
R262 B.n430 B.n48 256.663
R263 B.n430 B.n47 256.663
R264 B.n430 B.n46 256.663
R265 B.n430 B.n45 256.663
R266 B.n430 B.n44 256.663
R267 B.n430 B.n43 256.663
R268 B.n430 B.n42 256.663
R269 B.n430 B.n41 256.663
R270 B.n430 B.n40 256.663
R271 B.n430 B.n39 256.663
R272 B.n430 B.n38 256.663
R273 B.n430 B.n37 256.663
R274 B.n430 B.n36 256.663
R275 B.n430 B.n35 256.663
R276 B.n430 B.n34 256.663
R277 B.n430 B.n33 256.663
R278 B.n430 B.n32 256.663
R279 B.n430 B.n31 256.663
R280 B.n430 B.n30 256.663
R281 B.n430 B.n29 256.663
R282 B.n430 B.n28 256.663
R283 B.n430 B.n27 256.663
R284 B.n247 B.n209 256.663
R285 B.n253 B.n209 256.663
R286 B.n255 B.n209 256.663
R287 B.n261 B.n209 256.663
R288 B.n263 B.n209 256.663
R289 B.n269 B.n209 256.663
R290 B.n271 B.n209 256.663
R291 B.n277 B.n209 256.663
R292 B.n279 B.n209 256.663
R293 B.n285 B.n209 256.663
R294 B.n287 B.n209 256.663
R295 B.n293 B.n209 256.663
R296 B.n295 B.n209 256.663
R297 B.n302 B.n209 256.663
R298 B.n304 B.n209 256.663
R299 B.n310 B.n209 256.663
R300 B.n312 B.n209 256.663
R301 B.n318 B.n209 256.663
R302 B.n320 B.n209 256.663
R303 B.n326 B.n209 256.663
R304 B.n328 B.n209 256.663
R305 B.n334 B.n209 256.663
R306 B.n336 B.n209 256.663
R307 B.n342 B.n209 256.663
R308 B.n344 B.n209 256.663
R309 B.n350 B.n209 256.663
R310 B.n352 B.n209 256.663
R311 B.n358 B.n209 256.663
R312 B.n360 B.n209 256.663
R313 B.n366 B.n209 256.663
R314 B.n369 B.n209 256.663
R315 B.n376 B.n206 163.367
R316 B.n380 B.n206 163.367
R317 B.n380 B.n200 163.367
R318 B.n388 B.n200 163.367
R319 B.n388 B.n198 163.367
R320 B.n392 B.n198 163.367
R321 B.n392 B.n192 163.367
R322 B.n402 B.n192 163.367
R323 B.n402 B.n190 163.367
R324 B.n406 B.n190 163.367
R325 B.n406 B.n2 163.367
R326 B.n456 B.n2 163.367
R327 B.n456 B.n3 163.367
R328 B.n452 B.n3 163.367
R329 B.n452 B.n8 163.367
R330 B.n448 B.n8 163.367
R331 B.n448 B.n10 163.367
R332 B.n444 B.n10 163.367
R333 B.n444 B.n16 163.367
R334 B.n440 B.n16 163.367
R335 B.n440 B.n18 163.367
R336 B.n436 B.n18 163.367
R337 B.n436 B.n23 163.367
R338 B.n432 B.n23 163.367
R339 B.n248 B.n246 163.367
R340 B.n252 B.n246 163.367
R341 B.n256 B.n254 163.367
R342 B.n260 B.n244 163.367
R343 B.n264 B.n262 163.367
R344 B.n268 B.n242 163.367
R345 B.n272 B.n270 163.367
R346 B.n276 B.n240 163.367
R347 B.n280 B.n278 163.367
R348 B.n284 B.n238 163.367
R349 B.n288 B.n286 163.367
R350 B.n292 B.n236 163.367
R351 B.n296 B.n294 163.367
R352 B.n301 B.n232 163.367
R353 B.n305 B.n303 163.367
R354 B.n309 B.n230 163.367
R355 B.n313 B.n311 163.367
R356 B.n317 B.n228 163.367
R357 B.n321 B.n319 163.367
R358 B.n325 B.n223 163.367
R359 B.n329 B.n327 163.367
R360 B.n333 B.n221 163.367
R361 B.n337 B.n335 163.367
R362 B.n341 B.n219 163.367
R363 B.n345 B.n343 163.367
R364 B.n349 B.n217 163.367
R365 B.n353 B.n351 163.367
R366 B.n357 B.n215 163.367
R367 B.n361 B.n359 163.367
R368 B.n365 B.n213 163.367
R369 B.n368 B.n367 163.367
R370 B.n370 B.n210 163.367
R371 B.n374 B.n204 163.367
R372 B.n382 B.n204 163.367
R373 B.n382 B.n202 163.367
R374 B.n386 B.n202 163.367
R375 B.n386 B.n196 163.367
R376 B.n394 B.n196 163.367
R377 B.n394 B.n194 163.367
R378 B.n399 B.n194 163.367
R379 B.n399 B.n189 163.367
R380 B.n408 B.n189 163.367
R381 B.n409 B.n408 163.367
R382 B.n409 B.n5 163.367
R383 B.n6 B.n5 163.367
R384 B.n7 B.n6 163.367
R385 B.n414 B.n7 163.367
R386 B.n414 B.n12 163.367
R387 B.n13 B.n12 163.367
R388 B.n14 B.n13 163.367
R389 B.n419 B.n14 163.367
R390 B.n419 B.n19 163.367
R391 B.n20 B.n19 163.367
R392 B.n21 B.n20 163.367
R393 B.n424 B.n21 163.367
R394 B.n424 B.n26 163.367
R395 B.n65 B.n64 163.367
R396 B.n69 B.n68 163.367
R397 B.n73 B.n72 163.367
R398 B.n77 B.n76 163.367
R399 B.n81 B.n80 163.367
R400 B.n85 B.n84 163.367
R401 B.n89 B.n88 163.367
R402 B.n93 B.n92 163.367
R403 B.n97 B.n96 163.367
R404 B.n101 B.n100 163.367
R405 B.n105 B.n104 163.367
R406 B.n109 B.n108 163.367
R407 B.n113 B.n112 163.367
R408 B.n118 B.n117 163.367
R409 B.n122 B.n121 163.367
R410 B.n126 B.n125 163.367
R411 B.n130 B.n129 163.367
R412 B.n134 B.n133 163.367
R413 B.n139 B.n138 163.367
R414 B.n143 B.n142 163.367
R415 B.n147 B.n146 163.367
R416 B.n151 B.n150 163.367
R417 B.n155 B.n154 163.367
R418 B.n159 B.n158 163.367
R419 B.n163 B.n162 163.367
R420 B.n167 B.n166 163.367
R421 B.n171 B.n170 163.367
R422 B.n175 B.n174 163.367
R423 B.n179 B.n178 163.367
R424 B.n183 B.n182 163.367
R425 B.n185 B.n58 163.367
R426 B.n375 B.n209 116.35
R427 B.n431 B.n430 116.35
R428 B.n224 B.t15 87.7412
R429 B.n59 B.t4 87.7412
R430 B.n233 B.t12 87.7335
R431 B.n61 B.t7 87.7335
R432 B.n225 B.t14 74.5534
R433 B.n60 B.t5 74.5534
R434 B.n234 B.t11 74.5456
R435 B.n62 B.t8 74.5456
R436 B.n247 B.n208 71.676
R437 B.n253 B.n252 71.676
R438 B.n256 B.n255 71.676
R439 B.n261 B.n260 71.676
R440 B.n264 B.n263 71.676
R441 B.n269 B.n268 71.676
R442 B.n272 B.n271 71.676
R443 B.n277 B.n276 71.676
R444 B.n280 B.n279 71.676
R445 B.n285 B.n284 71.676
R446 B.n288 B.n287 71.676
R447 B.n293 B.n292 71.676
R448 B.n296 B.n295 71.676
R449 B.n302 B.n301 71.676
R450 B.n305 B.n304 71.676
R451 B.n310 B.n309 71.676
R452 B.n313 B.n312 71.676
R453 B.n318 B.n317 71.676
R454 B.n321 B.n320 71.676
R455 B.n326 B.n325 71.676
R456 B.n329 B.n328 71.676
R457 B.n334 B.n333 71.676
R458 B.n337 B.n336 71.676
R459 B.n342 B.n341 71.676
R460 B.n345 B.n344 71.676
R461 B.n350 B.n349 71.676
R462 B.n353 B.n352 71.676
R463 B.n358 B.n357 71.676
R464 B.n361 B.n360 71.676
R465 B.n366 B.n365 71.676
R466 B.n369 B.n368 71.676
R467 B.n27 B.n25 71.676
R468 B.n65 B.n28 71.676
R469 B.n69 B.n29 71.676
R470 B.n73 B.n30 71.676
R471 B.n77 B.n31 71.676
R472 B.n81 B.n32 71.676
R473 B.n85 B.n33 71.676
R474 B.n89 B.n34 71.676
R475 B.n93 B.n35 71.676
R476 B.n97 B.n36 71.676
R477 B.n101 B.n37 71.676
R478 B.n105 B.n38 71.676
R479 B.n109 B.n39 71.676
R480 B.n113 B.n40 71.676
R481 B.n118 B.n41 71.676
R482 B.n122 B.n42 71.676
R483 B.n126 B.n43 71.676
R484 B.n130 B.n44 71.676
R485 B.n134 B.n45 71.676
R486 B.n139 B.n46 71.676
R487 B.n143 B.n47 71.676
R488 B.n147 B.n48 71.676
R489 B.n151 B.n49 71.676
R490 B.n155 B.n50 71.676
R491 B.n159 B.n51 71.676
R492 B.n163 B.n52 71.676
R493 B.n167 B.n53 71.676
R494 B.n171 B.n54 71.676
R495 B.n175 B.n55 71.676
R496 B.n179 B.n56 71.676
R497 B.n183 B.n57 71.676
R498 B.n429 B.n58 71.676
R499 B.n429 B.n428 71.676
R500 B.n185 B.n57 71.676
R501 B.n182 B.n56 71.676
R502 B.n178 B.n55 71.676
R503 B.n174 B.n54 71.676
R504 B.n170 B.n53 71.676
R505 B.n166 B.n52 71.676
R506 B.n162 B.n51 71.676
R507 B.n158 B.n50 71.676
R508 B.n154 B.n49 71.676
R509 B.n150 B.n48 71.676
R510 B.n146 B.n47 71.676
R511 B.n142 B.n46 71.676
R512 B.n138 B.n45 71.676
R513 B.n133 B.n44 71.676
R514 B.n129 B.n43 71.676
R515 B.n125 B.n42 71.676
R516 B.n121 B.n41 71.676
R517 B.n117 B.n40 71.676
R518 B.n112 B.n39 71.676
R519 B.n108 B.n38 71.676
R520 B.n104 B.n37 71.676
R521 B.n100 B.n36 71.676
R522 B.n96 B.n35 71.676
R523 B.n92 B.n34 71.676
R524 B.n88 B.n33 71.676
R525 B.n84 B.n32 71.676
R526 B.n80 B.n31 71.676
R527 B.n76 B.n30 71.676
R528 B.n72 B.n29 71.676
R529 B.n68 B.n28 71.676
R530 B.n64 B.n27 71.676
R531 B.n248 B.n247 71.676
R532 B.n254 B.n253 71.676
R533 B.n255 B.n244 71.676
R534 B.n262 B.n261 71.676
R535 B.n263 B.n242 71.676
R536 B.n270 B.n269 71.676
R537 B.n271 B.n240 71.676
R538 B.n278 B.n277 71.676
R539 B.n279 B.n238 71.676
R540 B.n286 B.n285 71.676
R541 B.n287 B.n236 71.676
R542 B.n294 B.n293 71.676
R543 B.n295 B.n232 71.676
R544 B.n303 B.n302 71.676
R545 B.n304 B.n230 71.676
R546 B.n311 B.n310 71.676
R547 B.n312 B.n228 71.676
R548 B.n319 B.n318 71.676
R549 B.n320 B.n223 71.676
R550 B.n327 B.n326 71.676
R551 B.n328 B.n221 71.676
R552 B.n335 B.n334 71.676
R553 B.n336 B.n219 71.676
R554 B.n343 B.n342 71.676
R555 B.n344 B.n217 71.676
R556 B.n351 B.n350 71.676
R557 B.n352 B.n215 71.676
R558 B.n359 B.n358 71.676
R559 B.n360 B.n213 71.676
R560 B.n367 B.n366 71.676
R561 B.n370 B.n369 71.676
R562 B.n375 B.n205 60.3961
R563 B.n381 B.n205 60.3961
R564 B.n381 B.n201 60.3961
R565 B.n387 B.n201 60.3961
R566 B.n393 B.n197 60.3961
R567 B.n393 B.n193 60.3961
R568 B.n401 B.n193 60.3961
R569 B.n401 B.n400 60.3961
R570 B.n407 B.n4 60.3961
R571 B.n455 B.n4 60.3961
R572 B.n455 B.n454 60.3961
R573 B.n454 B.n453 60.3961
R574 B.n447 B.n11 60.3961
R575 B.n447 B.n446 60.3961
R576 B.n446 B.n445 60.3961
R577 B.n445 B.n15 60.3961
R578 B.n439 B.n438 60.3961
R579 B.n438 B.n437 60.3961
R580 B.n437 B.n22 60.3961
R581 B.n431 B.n22 60.3961
R582 B.n226 B.n225 59.5399
R583 B.n299 B.n234 59.5399
R584 B.n115 B.n62 59.5399
R585 B.n136 B.n60 59.5399
R586 B.t10 B.n197 48.8499
R587 B.t3 B.n15 48.8499
R588 B.n407 B.t0 36.4155
R589 B.n453 B.t1 36.4155
R590 B.n433 B.n24 33.8737
R591 B.n427 B.n426 33.8737
R592 B.n373 B.n372 33.8737
R593 B.n377 B.n207 33.8737
R594 B.n400 B.t0 23.9811
R595 B.n11 B.t1 23.9811
R596 B B.n457 18.0485
R597 B.n225 B.n224 13.1884
R598 B.n234 B.n233 13.1884
R599 B.n62 B.n61 13.1884
R600 B.n60 B.n59 13.1884
R601 B.n387 B.t10 11.5467
R602 B.n439 B.t3 11.5467
R603 B.n63 B.n24 10.6151
R604 B.n66 B.n63 10.6151
R605 B.n67 B.n66 10.6151
R606 B.n70 B.n67 10.6151
R607 B.n71 B.n70 10.6151
R608 B.n74 B.n71 10.6151
R609 B.n75 B.n74 10.6151
R610 B.n78 B.n75 10.6151
R611 B.n79 B.n78 10.6151
R612 B.n82 B.n79 10.6151
R613 B.n83 B.n82 10.6151
R614 B.n86 B.n83 10.6151
R615 B.n87 B.n86 10.6151
R616 B.n90 B.n87 10.6151
R617 B.n91 B.n90 10.6151
R618 B.n94 B.n91 10.6151
R619 B.n95 B.n94 10.6151
R620 B.n98 B.n95 10.6151
R621 B.n99 B.n98 10.6151
R622 B.n102 B.n99 10.6151
R623 B.n103 B.n102 10.6151
R624 B.n106 B.n103 10.6151
R625 B.n107 B.n106 10.6151
R626 B.n110 B.n107 10.6151
R627 B.n111 B.n110 10.6151
R628 B.n114 B.n111 10.6151
R629 B.n119 B.n116 10.6151
R630 B.n120 B.n119 10.6151
R631 B.n123 B.n120 10.6151
R632 B.n124 B.n123 10.6151
R633 B.n127 B.n124 10.6151
R634 B.n128 B.n127 10.6151
R635 B.n131 B.n128 10.6151
R636 B.n132 B.n131 10.6151
R637 B.n135 B.n132 10.6151
R638 B.n140 B.n137 10.6151
R639 B.n141 B.n140 10.6151
R640 B.n144 B.n141 10.6151
R641 B.n145 B.n144 10.6151
R642 B.n148 B.n145 10.6151
R643 B.n149 B.n148 10.6151
R644 B.n152 B.n149 10.6151
R645 B.n153 B.n152 10.6151
R646 B.n156 B.n153 10.6151
R647 B.n157 B.n156 10.6151
R648 B.n160 B.n157 10.6151
R649 B.n161 B.n160 10.6151
R650 B.n164 B.n161 10.6151
R651 B.n165 B.n164 10.6151
R652 B.n168 B.n165 10.6151
R653 B.n169 B.n168 10.6151
R654 B.n172 B.n169 10.6151
R655 B.n173 B.n172 10.6151
R656 B.n176 B.n173 10.6151
R657 B.n177 B.n176 10.6151
R658 B.n180 B.n177 10.6151
R659 B.n181 B.n180 10.6151
R660 B.n184 B.n181 10.6151
R661 B.n186 B.n184 10.6151
R662 B.n187 B.n186 10.6151
R663 B.n427 B.n187 10.6151
R664 B.n373 B.n203 10.6151
R665 B.n383 B.n203 10.6151
R666 B.n384 B.n383 10.6151
R667 B.n385 B.n384 10.6151
R668 B.n385 B.n195 10.6151
R669 B.n395 B.n195 10.6151
R670 B.n396 B.n395 10.6151
R671 B.n398 B.n396 10.6151
R672 B.n398 B.n397 10.6151
R673 B.n397 B.n188 10.6151
R674 B.n410 B.n188 10.6151
R675 B.n411 B.n410 10.6151
R676 B.n412 B.n411 10.6151
R677 B.n413 B.n412 10.6151
R678 B.n415 B.n413 10.6151
R679 B.n416 B.n415 10.6151
R680 B.n417 B.n416 10.6151
R681 B.n418 B.n417 10.6151
R682 B.n420 B.n418 10.6151
R683 B.n421 B.n420 10.6151
R684 B.n422 B.n421 10.6151
R685 B.n423 B.n422 10.6151
R686 B.n425 B.n423 10.6151
R687 B.n426 B.n425 10.6151
R688 B.n249 B.n207 10.6151
R689 B.n250 B.n249 10.6151
R690 B.n251 B.n250 10.6151
R691 B.n251 B.n245 10.6151
R692 B.n257 B.n245 10.6151
R693 B.n258 B.n257 10.6151
R694 B.n259 B.n258 10.6151
R695 B.n259 B.n243 10.6151
R696 B.n265 B.n243 10.6151
R697 B.n266 B.n265 10.6151
R698 B.n267 B.n266 10.6151
R699 B.n267 B.n241 10.6151
R700 B.n273 B.n241 10.6151
R701 B.n274 B.n273 10.6151
R702 B.n275 B.n274 10.6151
R703 B.n275 B.n239 10.6151
R704 B.n281 B.n239 10.6151
R705 B.n282 B.n281 10.6151
R706 B.n283 B.n282 10.6151
R707 B.n283 B.n237 10.6151
R708 B.n289 B.n237 10.6151
R709 B.n290 B.n289 10.6151
R710 B.n291 B.n290 10.6151
R711 B.n291 B.n235 10.6151
R712 B.n297 B.n235 10.6151
R713 B.n298 B.n297 10.6151
R714 B.n300 B.n231 10.6151
R715 B.n306 B.n231 10.6151
R716 B.n307 B.n306 10.6151
R717 B.n308 B.n307 10.6151
R718 B.n308 B.n229 10.6151
R719 B.n314 B.n229 10.6151
R720 B.n315 B.n314 10.6151
R721 B.n316 B.n315 10.6151
R722 B.n316 B.n227 10.6151
R723 B.n323 B.n322 10.6151
R724 B.n324 B.n323 10.6151
R725 B.n324 B.n222 10.6151
R726 B.n330 B.n222 10.6151
R727 B.n331 B.n330 10.6151
R728 B.n332 B.n331 10.6151
R729 B.n332 B.n220 10.6151
R730 B.n338 B.n220 10.6151
R731 B.n339 B.n338 10.6151
R732 B.n340 B.n339 10.6151
R733 B.n340 B.n218 10.6151
R734 B.n346 B.n218 10.6151
R735 B.n347 B.n346 10.6151
R736 B.n348 B.n347 10.6151
R737 B.n348 B.n216 10.6151
R738 B.n354 B.n216 10.6151
R739 B.n355 B.n354 10.6151
R740 B.n356 B.n355 10.6151
R741 B.n356 B.n214 10.6151
R742 B.n362 B.n214 10.6151
R743 B.n363 B.n362 10.6151
R744 B.n364 B.n363 10.6151
R745 B.n364 B.n212 10.6151
R746 B.n212 B.n211 10.6151
R747 B.n371 B.n211 10.6151
R748 B.n372 B.n371 10.6151
R749 B.n378 B.n377 10.6151
R750 B.n379 B.n378 10.6151
R751 B.n379 B.n199 10.6151
R752 B.n389 B.n199 10.6151
R753 B.n390 B.n389 10.6151
R754 B.n391 B.n390 10.6151
R755 B.n391 B.n191 10.6151
R756 B.n403 B.n191 10.6151
R757 B.n404 B.n403 10.6151
R758 B.n405 B.n404 10.6151
R759 B.n405 B.n0 10.6151
R760 B.n451 B.n1 10.6151
R761 B.n451 B.n450 10.6151
R762 B.n450 B.n449 10.6151
R763 B.n449 B.n9 10.6151
R764 B.n443 B.n9 10.6151
R765 B.n443 B.n442 10.6151
R766 B.n442 B.n441 10.6151
R767 B.n441 B.n17 10.6151
R768 B.n435 B.n17 10.6151
R769 B.n435 B.n434 10.6151
R770 B.n434 B.n433 10.6151
R771 B.n115 B.n114 8.74196
R772 B.n137 B.n136 8.74196
R773 B.n299 B.n298 8.74196
R774 B.n322 B.n226 8.74196
R775 B.n457 B.n0 2.81026
R776 B.n457 B.n1 2.81026
R777 B.n116 B.n115 1.87367
R778 B.n136 B.n135 1.87367
R779 B.n300 B.n299 1.87367
R780 B.n227 B.n226 1.87367
R781 VP.n0 VP.t0 797.409
R782 VP.n0 VP.t1 762.423
R783 VP VP.n0 0.0516364
R784 VDD1 VDD1.t0 100.231
R785 VDD1 VDD1.t1 68.8024
C0 VDD2 VTAIL 4.44062f
C1 VTAIL VN 0.685777f
C2 VTAIL VP 0.700256f
C3 VDD1 VDD2 0.429231f
C4 VDD1 VN 0.148429f
C5 VDD1 VP 1.08292f
C6 VDD2 VN 0.994668f
C7 VDD2 VP 0.239634f
C8 VP VN 3.49406f
C9 VDD1 VTAIL 4.407279f
C10 VDD2 B 2.735787f
C11 VDD1 B 4.74236f
C12 VTAIL B 3.949302f
C13 VN B 6.09722f
C14 VP B 3.237105f
C15 VDD1.t1 B 1.09627f
C16 VDD1.t0 B 1.38704f
C17 VP.t0 B 0.399172f
C18 VP.t1 B 0.338219f
C19 VP.n0 B 2.75688f
C20 VDD2.t0 B 1.39078f
C21 VDD2.t1 B 1.11253f
C22 VDD2.n0 B 1.86671f
C23 VTAIL.t0 B 1.16154f
C24 VTAIL.n0 B 1.05185f
C25 VTAIL.t2 B 1.16154f
C26 VTAIL.n1 B 1.05762f
C27 VTAIL.t1 B 1.16154f
C28 VTAIL.n2 B 1.01929f
C29 VTAIL.t3 B 1.16154f
C30 VTAIL.n3 B 0.975179f
C31 VN.t1 B 0.332451f
C32 VN.t0 B 0.394231f
.ends

