* NGSPICE file created from diff_pair_sample_1032.ext - technology: sky130A

.subckt diff_pair_sample_1032 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t3 VP.t0 VTAIL.t7 w_n3562_n2922# sky130_fd_pr__pfet_01v8 ad=1.61205 pd=10.1 as=3.8103 ps=20.32 w=9.77 l=3.99
X1 VDD2.t3 VN.t0 VTAIL.t3 w_n3562_n2922# sky130_fd_pr__pfet_01v8 ad=1.61205 pd=10.1 as=3.8103 ps=20.32 w=9.77 l=3.99
X2 B.t11 B.t9 B.t10 w_n3562_n2922# sky130_fd_pr__pfet_01v8 ad=3.8103 pd=20.32 as=0 ps=0 w=9.77 l=3.99
X3 VDD2.t2 VN.t1 VTAIL.t1 w_n3562_n2922# sky130_fd_pr__pfet_01v8 ad=1.61205 pd=10.1 as=3.8103 ps=20.32 w=9.77 l=3.99
X4 VTAIL.t0 VN.t2 VDD2.t1 w_n3562_n2922# sky130_fd_pr__pfet_01v8 ad=3.8103 pd=20.32 as=1.61205 ps=10.1 w=9.77 l=3.99
X5 VDD1.t2 VP.t1 VTAIL.t5 w_n3562_n2922# sky130_fd_pr__pfet_01v8 ad=1.61205 pd=10.1 as=3.8103 ps=20.32 w=9.77 l=3.99
X6 VTAIL.t2 VN.t3 VDD2.t0 w_n3562_n2922# sky130_fd_pr__pfet_01v8 ad=3.8103 pd=20.32 as=1.61205 ps=10.1 w=9.77 l=3.99
X7 B.t8 B.t6 B.t7 w_n3562_n2922# sky130_fd_pr__pfet_01v8 ad=3.8103 pd=20.32 as=0 ps=0 w=9.77 l=3.99
X8 VTAIL.t4 VP.t2 VDD1.t1 w_n3562_n2922# sky130_fd_pr__pfet_01v8 ad=3.8103 pd=20.32 as=1.61205 ps=10.1 w=9.77 l=3.99
X9 B.t5 B.t3 B.t4 w_n3562_n2922# sky130_fd_pr__pfet_01v8 ad=3.8103 pd=20.32 as=0 ps=0 w=9.77 l=3.99
X10 B.t2 B.t0 B.t1 w_n3562_n2922# sky130_fd_pr__pfet_01v8 ad=3.8103 pd=20.32 as=0 ps=0 w=9.77 l=3.99
X11 VTAIL.t6 VP.t3 VDD1.t0 w_n3562_n2922# sky130_fd_pr__pfet_01v8 ad=3.8103 pd=20.32 as=1.61205 ps=10.1 w=9.77 l=3.99
R0 VP.n18 VP.n0 161.3
R1 VP.n17 VP.n16 161.3
R2 VP.n15 VP.n1 161.3
R3 VP.n14 VP.n13 161.3
R4 VP.n12 VP.n2 161.3
R5 VP.n11 VP.n10 161.3
R6 VP.n9 VP.n3 161.3
R7 VP.n8 VP.n7 161.3
R8 VP.n4 VP.t2 92.8018
R9 VP.n4 VP.t1 91.3581
R10 VP.n6 VP.n5 62.1188
R11 VP.n20 VP.n19 62.1188
R12 VP.n6 VP.t3 59.0123
R13 VP.n19 VP.t0 59.0123
R14 VP.n13 VP.n12 56.5193
R15 VP.n5 VP.n4 50.7423
R16 VP.n7 VP.n3 24.4675
R17 VP.n11 VP.n3 24.4675
R18 VP.n12 VP.n11 24.4675
R19 VP.n13 VP.n1 24.4675
R20 VP.n17 VP.n1 24.4675
R21 VP.n18 VP.n17 24.4675
R22 VP.n7 VP.n6 20.0634
R23 VP.n19 VP.n18 20.0634
R24 VP.n8 VP.n5 0.417535
R25 VP.n20 VP.n0 0.417535
R26 VP VP.n20 0.394291
R27 VP.n9 VP.n8 0.189894
R28 VP.n10 VP.n9 0.189894
R29 VP.n10 VP.n2 0.189894
R30 VP.n14 VP.n2 0.189894
R31 VP.n15 VP.n14 0.189894
R32 VP.n16 VP.n15 0.189894
R33 VP.n16 VP.n0 0.189894
R34 VTAIL.n5 VTAIL.t4 67.7655
R35 VTAIL.n4 VTAIL.t1 67.7655
R36 VTAIL.n3 VTAIL.t2 67.7655
R37 VTAIL.n7 VTAIL.t3 67.7654
R38 VTAIL.n0 VTAIL.t0 67.7654
R39 VTAIL.n1 VTAIL.t7 67.7654
R40 VTAIL.n2 VTAIL.t6 67.7654
R41 VTAIL.n6 VTAIL.t5 67.7654
R42 VTAIL.n7 VTAIL.n6 24.5134
R43 VTAIL.n3 VTAIL.n2 24.5134
R44 VTAIL.n4 VTAIL.n3 3.72464
R45 VTAIL.n6 VTAIL.n5 3.72464
R46 VTAIL.n2 VTAIL.n1 3.72464
R47 VTAIL VTAIL.n0 1.92076
R48 VTAIL VTAIL.n7 1.80438
R49 VTAIL.n5 VTAIL.n4 0.470328
R50 VTAIL.n1 VTAIL.n0 0.470328
R51 VDD1 VDD1.n1 124.951
R52 VDD1 VDD1.n0 81.1754
R53 VDD1.n0 VDD1.t1 3.32752
R54 VDD1.n0 VDD1.t2 3.32752
R55 VDD1.n1 VDD1.t0 3.32752
R56 VDD1.n1 VDD1.t3 3.32752
R57 VN.n0 VN.t2 92.8022
R58 VN.n1 VN.t1 92.8022
R59 VN.n0 VN.t0 91.3581
R60 VN.n1 VN.t3 91.3581
R61 VN VN.n1 50.7803
R62 VN VN.n0 1.73105
R63 VDD2.n2 VDD2.n0 124.427
R64 VDD2.n2 VDD2.n1 81.1172
R65 VDD2.n1 VDD2.t0 3.32752
R66 VDD2.n1 VDD2.t2 3.32752
R67 VDD2.n0 VDD2.t1 3.32752
R68 VDD2.n0 VDD2.t3 3.32752
R69 VDD2 VDD2.n2 0.0586897
R70 B.n513 B.n512 585
R71 B.n514 B.n69 585
R72 B.n516 B.n515 585
R73 B.n517 B.n68 585
R74 B.n519 B.n518 585
R75 B.n520 B.n67 585
R76 B.n522 B.n521 585
R77 B.n523 B.n66 585
R78 B.n525 B.n524 585
R79 B.n526 B.n65 585
R80 B.n528 B.n527 585
R81 B.n529 B.n64 585
R82 B.n531 B.n530 585
R83 B.n532 B.n63 585
R84 B.n534 B.n533 585
R85 B.n535 B.n62 585
R86 B.n537 B.n536 585
R87 B.n538 B.n61 585
R88 B.n540 B.n539 585
R89 B.n541 B.n60 585
R90 B.n543 B.n542 585
R91 B.n544 B.n59 585
R92 B.n546 B.n545 585
R93 B.n547 B.n58 585
R94 B.n549 B.n548 585
R95 B.n550 B.n57 585
R96 B.n552 B.n551 585
R97 B.n553 B.n56 585
R98 B.n555 B.n554 585
R99 B.n556 B.n55 585
R100 B.n558 B.n557 585
R101 B.n559 B.n54 585
R102 B.n561 B.n560 585
R103 B.n562 B.n53 585
R104 B.n564 B.n563 585
R105 B.n566 B.n50 585
R106 B.n568 B.n567 585
R107 B.n569 B.n49 585
R108 B.n571 B.n570 585
R109 B.n572 B.n48 585
R110 B.n574 B.n573 585
R111 B.n575 B.n47 585
R112 B.n577 B.n576 585
R113 B.n578 B.n43 585
R114 B.n580 B.n579 585
R115 B.n581 B.n42 585
R116 B.n583 B.n582 585
R117 B.n584 B.n41 585
R118 B.n586 B.n585 585
R119 B.n587 B.n40 585
R120 B.n589 B.n588 585
R121 B.n590 B.n39 585
R122 B.n592 B.n591 585
R123 B.n593 B.n38 585
R124 B.n595 B.n594 585
R125 B.n596 B.n37 585
R126 B.n598 B.n597 585
R127 B.n599 B.n36 585
R128 B.n601 B.n600 585
R129 B.n602 B.n35 585
R130 B.n604 B.n603 585
R131 B.n605 B.n34 585
R132 B.n607 B.n606 585
R133 B.n608 B.n33 585
R134 B.n610 B.n609 585
R135 B.n611 B.n32 585
R136 B.n613 B.n612 585
R137 B.n614 B.n31 585
R138 B.n616 B.n615 585
R139 B.n617 B.n30 585
R140 B.n619 B.n618 585
R141 B.n620 B.n29 585
R142 B.n622 B.n621 585
R143 B.n623 B.n28 585
R144 B.n625 B.n624 585
R145 B.n626 B.n27 585
R146 B.n628 B.n627 585
R147 B.n629 B.n26 585
R148 B.n631 B.n630 585
R149 B.n632 B.n25 585
R150 B.n511 B.n70 585
R151 B.n510 B.n509 585
R152 B.n508 B.n71 585
R153 B.n507 B.n506 585
R154 B.n505 B.n72 585
R155 B.n504 B.n503 585
R156 B.n502 B.n73 585
R157 B.n501 B.n500 585
R158 B.n499 B.n74 585
R159 B.n498 B.n497 585
R160 B.n496 B.n75 585
R161 B.n495 B.n494 585
R162 B.n493 B.n76 585
R163 B.n492 B.n491 585
R164 B.n490 B.n77 585
R165 B.n489 B.n488 585
R166 B.n487 B.n78 585
R167 B.n486 B.n485 585
R168 B.n484 B.n79 585
R169 B.n483 B.n482 585
R170 B.n481 B.n80 585
R171 B.n480 B.n479 585
R172 B.n478 B.n81 585
R173 B.n477 B.n476 585
R174 B.n475 B.n82 585
R175 B.n474 B.n473 585
R176 B.n472 B.n83 585
R177 B.n471 B.n470 585
R178 B.n469 B.n84 585
R179 B.n468 B.n467 585
R180 B.n466 B.n85 585
R181 B.n465 B.n464 585
R182 B.n463 B.n86 585
R183 B.n462 B.n461 585
R184 B.n460 B.n87 585
R185 B.n459 B.n458 585
R186 B.n457 B.n88 585
R187 B.n456 B.n455 585
R188 B.n454 B.n89 585
R189 B.n453 B.n452 585
R190 B.n451 B.n90 585
R191 B.n450 B.n449 585
R192 B.n448 B.n91 585
R193 B.n447 B.n446 585
R194 B.n445 B.n92 585
R195 B.n444 B.n443 585
R196 B.n442 B.n93 585
R197 B.n441 B.n440 585
R198 B.n439 B.n94 585
R199 B.n438 B.n437 585
R200 B.n436 B.n95 585
R201 B.n435 B.n434 585
R202 B.n433 B.n96 585
R203 B.n432 B.n431 585
R204 B.n430 B.n97 585
R205 B.n429 B.n428 585
R206 B.n427 B.n98 585
R207 B.n426 B.n425 585
R208 B.n424 B.n99 585
R209 B.n423 B.n422 585
R210 B.n421 B.n100 585
R211 B.n420 B.n419 585
R212 B.n418 B.n101 585
R213 B.n417 B.n416 585
R214 B.n415 B.n102 585
R215 B.n414 B.n413 585
R216 B.n412 B.n103 585
R217 B.n411 B.n410 585
R218 B.n409 B.n104 585
R219 B.n408 B.n407 585
R220 B.n406 B.n105 585
R221 B.n405 B.n404 585
R222 B.n403 B.n106 585
R223 B.n402 B.n401 585
R224 B.n400 B.n107 585
R225 B.n399 B.n398 585
R226 B.n397 B.n108 585
R227 B.n396 B.n395 585
R228 B.n394 B.n109 585
R229 B.n393 B.n392 585
R230 B.n391 B.n110 585
R231 B.n390 B.n389 585
R232 B.n388 B.n111 585
R233 B.n387 B.n386 585
R234 B.n385 B.n112 585
R235 B.n384 B.n383 585
R236 B.n382 B.n113 585
R237 B.n381 B.n380 585
R238 B.n379 B.n114 585
R239 B.n378 B.n377 585
R240 B.n376 B.n115 585
R241 B.n375 B.n374 585
R242 B.n373 B.n116 585
R243 B.n252 B.n251 585
R244 B.n253 B.n160 585
R245 B.n255 B.n254 585
R246 B.n256 B.n159 585
R247 B.n258 B.n257 585
R248 B.n259 B.n158 585
R249 B.n261 B.n260 585
R250 B.n262 B.n157 585
R251 B.n264 B.n263 585
R252 B.n265 B.n156 585
R253 B.n267 B.n266 585
R254 B.n268 B.n155 585
R255 B.n270 B.n269 585
R256 B.n271 B.n154 585
R257 B.n273 B.n272 585
R258 B.n274 B.n153 585
R259 B.n276 B.n275 585
R260 B.n277 B.n152 585
R261 B.n279 B.n278 585
R262 B.n280 B.n151 585
R263 B.n282 B.n281 585
R264 B.n283 B.n150 585
R265 B.n285 B.n284 585
R266 B.n286 B.n149 585
R267 B.n288 B.n287 585
R268 B.n289 B.n148 585
R269 B.n291 B.n290 585
R270 B.n292 B.n147 585
R271 B.n294 B.n293 585
R272 B.n295 B.n146 585
R273 B.n297 B.n296 585
R274 B.n298 B.n145 585
R275 B.n300 B.n299 585
R276 B.n301 B.n144 585
R277 B.n303 B.n302 585
R278 B.n305 B.n304 585
R279 B.n306 B.n140 585
R280 B.n308 B.n307 585
R281 B.n309 B.n139 585
R282 B.n311 B.n310 585
R283 B.n312 B.n138 585
R284 B.n314 B.n313 585
R285 B.n315 B.n137 585
R286 B.n317 B.n316 585
R287 B.n318 B.n134 585
R288 B.n321 B.n320 585
R289 B.n322 B.n133 585
R290 B.n324 B.n323 585
R291 B.n325 B.n132 585
R292 B.n327 B.n326 585
R293 B.n328 B.n131 585
R294 B.n330 B.n329 585
R295 B.n331 B.n130 585
R296 B.n333 B.n332 585
R297 B.n334 B.n129 585
R298 B.n336 B.n335 585
R299 B.n337 B.n128 585
R300 B.n339 B.n338 585
R301 B.n340 B.n127 585
R302 B.n342 B.n341 585
R303 B.n343 B.n126 585
R304 B.n345 B.n344 585
R305 B.n346 B.n125 585
R306 B.n348 B.n347 585
R307 B.n349 B.n124 585
R308 B.n351 B.n350 585
R309 B.n352 B.n123 585
R310 B.n354 B.n353 585
R311 B.n355 B.n122 585
R312 B.n357 B.n356 585
R313 B.n358 B.n121 585
R314 B.n360 B.n359 585
R315 B.n361 B.n120 585
R316 B.n363 B.n362 585
R317 B.n364 B.n119 585
R318 B.n366 B.n365 585
R319 B.n367 B.n118 585
R320 B.n369 B.n368 585
R321 B.n370 B.n117 585
R322 B.n372 B.n371 585
R323 B.n250 B.n161 585
R324 B.n249 B.n248 585
R325 B.n247 B.n162 585
R326 B.n246 B.n245 585
R327 B.n244 B.n163 585
R328 B.n243 B.n242 585
R329 B.n241 B.n164 585
R330 B.n240 B.n239 585
R331 B.n238 B.n165 585
R332 B.n237 B.n236 585
R333 B.n235 B.n166 585
R334 B.n234 B.n233 585
R335 B.n232 B.n167 585
R336 B.n231 B.n230 585
R337 B.n229 B.n168 585
R338 B.n228 B.n227 585
R339 B.n226 B.n169 585
R340 B.n225 B.n224 585
R341 B.n223 B.n170 585
R342 B.n222 B.n221 585
R343 B.n220 B.n171 585
R344 B.n219 B.n218 585
R345 B.n217 B.n172 585
R346 B.n216 B.n215 585
R347 B.n214 B.n173 585
R348 B.n213 B.n212 585
R349 B.n211 B.n174 585
R350 B.n210 B.n209 585
R351 B.n208 B.n175 585
R352 B.n207 B.n206 585
R353 B.n205 B.n176 585
R354 B.n204 B.n203 585
R355 B.n202 B.n177 585
R356 B.n201 B.n200 585
R357 B.n199 B.n178 585
R358 B.n198 B.n197 585
R359 B.n196 B.n179 585
R360 B.n195 B.n194 585
R361 B.n193 B.n180 585
R362 B.n192 B.n191 585
R363 B.n190 B.n181 585
R364 B.n189 B.n188 585
R365 B.n187 B.n182 585
R366 B.n186 B.n185 585
R367 B.n184 B.n183 585
R368 B.n2 B.n0 585
R369 B.n701 B.n1 585
R370 B.n700 B.n699 585
R371 B.n698 B.n3 585
R372 B.n697 B.n696 585
R373 B.n695 B.n4 585
R374 B.n694 B.n693 585
R375 B.n692 B.n5 585
R376 B.n691 B.n690 585
R377 B.n689 B.n6 585
R378 B.n688 B.n687 585
R379 B.n686 B.n7 585
R380 B.n685 B.n684 585
R381 B.n683 B.n8 585
R382 B.n682 B.n681 585
R383 B.n680 B.n9 585
R384 B.n679 B.n678 585
R385 B.n677 B.n10 585
R386 B.n676 B.n675 585
R387 B.n674 B.n11 585
R388 B.n673 B.n672 585
R389 B.n671 B.n12 585
R390 B.n670 B.n669 585
R391 B.n668 B.n13 585
R392 B.n667 B.n666 585
R393 B.n665 B.n14 585
R394 B.n664 B.n663 585
R395 B.n662 B.n15 585
R396 B.n661 B.n660 585
R397 B.n659 B.n16 585
R398 B.n658 B.n657 585
R399 B.n656 B.n17 585
R400 B.n655 B.n654 585
R401 B.n653 B.n18 585
R402 B.n652 B.n651 585
R403 B.n650 B.n19 585
R404 B.n649 B.n648 585
R405 B.n647 B.n20 585
R406 B.n646 B.n645 585
R407 B.n644 B.n21 585
R408 B.n643 B.n642 585
R409 B.n641 B.n22 585
R410 B.n640 B.n639 585
R411 B.n638 B.n23 585
R412 B.n637 B.n636 585
R413 B.n635 B.n24 585
R414 B.n634 B.n633 585
R415 B.n703 B.n702 585
R416 B.n251 B.n250 511.721
R417 B.n634 B.n25 511.721
R418 B.n371 B.n116 511.721
R419 B.n513 B.n70 511.721
R420 B.n135 B.t9 268.497
R421 B.n141 B.t3 268.497
R422 B.n44 B.t6 268.497
R423 B.n51 B.t0 268.497
R424 B.n135 B.t11 196.397
R425 B.n51 B.t1 196.397
R426 B.n141 B.t5 196.386
R427 B.n44 B.t7 196.386
R428 B.n250 B.n249 163.367
R429 B.n249 B.n162 163.367
R430 B.n245 B.n162 163.367
R431 B.n245 B.n244 163.367
R432 B.n244 B.n243 163.367
R433 B.n243 B.n164 163.367
R434 B.n239 B.n164 163.367
R435 B.n239 B.n238 163.367
R436 B.n238 B.n237 163.367
R437 B.n237 B.n166 163.367
R438 B.n233 B.n166 163.367
R439 B.n233 B.n232 163.367
R440 B.n232 B.n231 163.367
R441 B.n231 B.n168 163.367
R442 B.n227 B.n168 163.367
R443 B.n227 B.n226 163.367
R444 B.n226 B.n225 163.367
R445 B.n225 B.n170 163.367
R446 B.n221 B.n170 163.367
R447 B.n221 B.n220 163.367
R448 B.n220 B.n219 163.367
R449 B.n219 B.n172 163.367
R450 B.n215 B.n172 163.367
R451 B.n215 B.n214 163.367
R452 B.n214 B.n213 163.367
R453 B.n213 B.n174 163.367
R454 B.n209 B.n174 163.367
R455 B.n209 B.n208 163.367
R456 B.n208 B.n207 163.367
R457 B.n207 B.n176 163.367
R458 B.n203 B.n176 163.367
R459 B.n203 B.n202 163.367
R460 B.n202 B.n201 163.367
R461 B.n201 B.n178 163.367
R462 B.n197 B.n178 163.367
R463 B.n197 B.n196 163.367
R464 B.n196 B.n195 163.367
R465 B.n195 B.n180 163.367
R466 B.n191 B.n180 163.367
R467 B.n191 B.n190 163.367
R468 B.n190 B.n189 163.367
R469 B.n189 B.n182 163.367
R470 B.n185 B.n182 163.367
R471 B.n185 B.n184 163.367
R472 B.n184 B.n2 163.367
R473 B.n702 B.n2 163.367
R474 B.n702 B.n701 163.367
R475 B.n701 B.n700 163.367
R476 B.n700 B.n3 163.367
R477 B.n696 B.n3 163.367
R478 B.n696 B.n695 163.367
R479 B.n695 B.n694 163.367
R480 B.n694 B.n5 163.367
R481 B.n690 B.n5 163.367
R482 B.n690 B.n689 163.367
R483 B.n689 B.n688 163.367
R484 B.n688 B.n7 163.367
R485 B.n684 B.n7 163.367
R486 B.n684 B.n683 163.367
R487 B.n683 B.n682 163.367
R488 B.n682 B.n9 163.367
R489 B.n678 B.n9 163.367
R490 B.n678 B.n677 163.367
R491 B.n677 B.n676 163.367
R492 B.n676 B.n11 163.367
R493 B.n672 B.n11 163.367
R494 B.n672 B.n671 163.367
R495 B.n671 B.n670 163.367
R496 B.n670 B.n13 163.367
R497 B.n666 B.n13 163.367
R498 B.n666 B.n665 163.367
R499 B.n665 B.n664 163.367
R500 B.n664 B.n15 163.367
R501 B.n660 B.n15 163.367
R502 B.n660 B.n659 163.367
R503 B.n659 B.n658 163.367
R504 B.n658 B.n17 163.367
R505 B.n654 B.n17 163.367
R506 B.n654 B.n653 163.367
R507 B.n653 B.n652 163.367
R508 B.n652 B.n19 163.367
R509 B.n648 B.n19 163.367
R510 B.n648 B.n647 163.367
R511 B.n647 B.n646 163.367
R512 B.n646 B.n21 163.367
R513 B.n642 B.n21 163.367
R514 B.n642 B.n641 163.367
R515 B.n641 B.n640 163.367
R516 B.n640 B.n23 163.367
R517 B.n636 B.n23 163.367
R518 B.n636 B.n635 163.367
R519 B.n635 B.n634 163.367
R520 B.n251 B.n160 163.367
R521 B.n255 B.n160 163.367
R522 B.n256 B.n255 163.367
R523 B.n257 B.n256 163.367
R524 B.n257 B.n158 163.367
R525 B.n261 B.n158 163.367
R526 B.n262 B.n261 163.367
R527 B.n263 B.n262 163.367
R528 B.n263 B.n156 163.367
R529 B.n267 B.n156 163.367
R530 B.n268 B.n267 163.367
R531 B.n269 B.n268 163.367
R532 B.n269 B.n154 163.367
R533 B.n273 B.n154 163.367
R534 B.n274 B.n273 163.367
R535 B.n275 B.n274 163.367
R536 B.n275 B.n152 163.367
R537 B.n279 B.n152 163.367
R538 B.n280 B.n279 163.367
R539 B.n281 B.n280 163.367
R540 B.n281 B.n150 163.367
R541 B.n285 B.n150 163.367
R542 B.n286 B.n285 163.367
R543 B.n287 B.n286 163.367
R544 B.n287 B.n148 163.367
R545 B.n291 B.n148 163.367
R546 B.n292 B.n291 163.367
R547 B.n293 B.n292 163.367
R548 B.n293 B.n146 163.367
R549 B.n297 B.n146 163.367
R550 B.n298 B.n297 163.367
R551 B.n299 B.n298 163.367
R552 B.n299 B.n144 163.367
R553 B.n303 B.n144 163.367
R554 B.n304 B.n303 163.367
R555 B.n304 B.n140 163.367
R556 B.n308 B.n140 163.367
R557 B.n309 B.n308 163.367
R558 B.n310 B.n309 163.367
R559 B.n310 B.n138 163.367
R560 B.n314 B.n138 163.367
R561 B.n315 B.n314 163.367
R562 B.n316 B.n315 163.367
R563 B.n316 B.n134 163.367
R564 B.n321 B.n134 163.367
R565 B.n322 B.n321 163.367
R566 B.n323 B.n322 163.367
R567 B.n323 B.n132 163.367
R568 B.n327 B.n132 163.367
R569 B.n328 B.n327 163.367
R570 B.n329 B.n328 163.367
R571 B.n329 B.n130 163.367
R572 B.n333 B.n130 163.367
R573 B.n334 B.n333 163.367
R574 B.n335 B.n334 163.367
R575 B.n335 B.n128 163.367
R576 B.n339 B.n128 163.367
R577 B.n340 B.n339 163.367
R578 B.n341 B.n340 163.367
R579 B.n341 B.n126 163.367
R580 B.n345 B.n126 163.367
R581 B.n346 B.n345 163.367
R582 B.n347 B.n346 163.367
R583 B.n347 B.n124 163.367
R584 B.n351 B.n124 163.367
R585 B.n352 B.n351 163.367
R586 B.n353 B.n352 163.367
R587 B.n353 B.n122 163.367
R588 B.n357 B.n122 163.367
R589 B.n358 B.n357 163.367
R590 B.n359 B.n358 163.367
R591 B.n359 B.n120 163.367
R592 B.n363 B.n120 163.367
R593 B.n364 B.n363 163.367
R594 B.n365 B.n364 163.367
R595 B.n365 B.n118 163.367
R596 B.n369 B.n118 163.367
R597 B.n370 B.n369 163.367
R598 B.n371 B.n370 163.367
R599 B.n375 B.n116 163.367
R600 B.n376 B.n375 163.367
R601 B.n377 B.n376 163.367
R602 B.n377 B.n114 163.367
R603 B.n381 B.n114 163.367
R604 B.n382 B.n381 163.367
R605 B.n383 B.n382 163.367
R606 B.n383 B.n112 163.367
R607 B.n387 B.n112 163.367
R608 B.n388 B.n387 163.367
R609 B.n389 B.n388 163.367
R610 B.n389 B.n110 163.367
R611 B.n393 B.n110 163.367
R612 B.n394 B.n393 163.367
R613 B.n395 B.n394 163.367
R614 B.n395 B.n108 163.367
R615 B.n399 B.n108 163.367
R616 B.n400 B.n399 163.367
R617 B.n401 B.n400 163.367
R618 B.n401 B.n106 163.367
R619 B.n405 B.n106 163.367
R620 B.n406 B.n405 163.367
R621 B.n407 B.n406 163.367
R622 B.n407 B.n104 163.367
R623 B.n411 B.n104 163.367
R624 B.n412 B.n411 163.367
R625 B.n413 B.n412 163.367
R626 B.n413 B.n102 163.367
R627 B.n417 B.n102 163.367
R628 B.n418 B.n417 163.367
R629 B.n419 B.n418 163.367
R630 B.n419 B.n100 163.367
R631 B.n423 B.n100 163.367
R632 B.n424 B.n423 163.367
R633 B.n425 B.n424 163.367
R634 B.n425 B.n98 163.367
R635 B.n429 B.n98 163.367
R636 B.n430 B.n429 163.367
R637 B.n431 B.n430 163.367
R638 B.n431 B.n96 163.367
R639 B.n435 B.n96 163.367
R640 B.n436 B.n435 163.367
R641 B.n437 B.n436 163.367
R642 B.n437 B.n94 163.367
R643 B.n441 B.n94 163.367
R644 B.n442 B.n441 163.367
R645 B.n443 B.n442 163.367
R646 B.n443 B.n92 163.367
R647 B.n447 B.n92 163.367
R648 B.n448 B.n447 163.367
R649 B.n449 B.n448 163.367
R650 B.n449 B.n90 163.367
R651 B.n453 B.n90 163.367
R652 B.n454 B.n453 163.367
R653 B.n455 B.n454 163.367
R654 B.n455 B.n88 163.367
R655 B.n459 B.n88 163.367
R656 B.n460 B.n459 163.367
R657 B.n461 B.n460 163.367
R658 B.n461 B.n86 163.367
R659 B.n465 B.n86 163.367
R660 B.n466 B.n465 163.367
R661 B.n467 B.n466 163.367
R662 B.n467 B.n84 163.367
R663 B.n471 B.n84 163.367
R664 B.n472 B.n471 163.367
R665 B.n473 B.n472 163.367
R666 B.n473 B.n82 163.367
R667 B.n477 B.n82 163.367
R668 B.n478 B.n477 163.367
R669 B.n479 B.n478 163.367
R670 B.n479 B.n80 163.367
R671 B.n483 B.n80 163.367
R672 B.n484 B.n483 163.367
R673 B.n485 B.n484 163.367
R674 B.n485 B.n78 163.367
R675 B.n489 B.n78 163.367
R676 B.n490 B.n489 163.367
R677 B.n491 B.n490 163.367
R678 B.n491 B.n76 163.367
R679 B.n495 B.n76 163.367
R680 B.n496 B.n495 163.367
R681 B.n497 B.n496 163.367
R682 B.n497 B.n74 163.367
R683 B.n501 B.n74 163.367
R684 B.n502 B.n501 163.367
R685 B.n503 B.n502 163.367
R686 B.n503 B.n72 163.367
R687 B.n507 B.n72 163.367
R688 B.n508 B.n507 163.367
R689 B.n509 B.n508 163.367
R690 B.n509 B.n70 163.367
R691 B.n630 B.n25 163.367
R692 B.n630 B.n629 163.367
R693 B.n629 B.n628 163.367
R694 B.n628 B.n27 163.367
R695 B.n624 B.n27 163.367
R696 B.n624 B.n623 163.367
R697 B.n623 B.n622 163.367
R698 B.n622 B.n29 163.367
R699 B.n618 B.n29 163.367
R700 B.n618 B.n617 163.367
R701 B.n617 B.n616 163.367
R702 B.n616 B.n31 163.367
R703 B.n612 B.n31 163.367
R704 B.n612 B.n611 163.367
R705 B.n611 B.n610 163.367
R706 B.n610 B.n33 163.367
R707 B.n606 B.n33 163.367
R708 B.n606 B.n605 163.367
R709 B.n605 B.n604 163.367
R710 B.n604 B.n35 163.367
R711 B.n600 B.n35 163.367
R712 B.n600 B.n599 163.367
R713 B.n599 B.n598 163.367
R714 B.n598 B.n37 163.367
R715 B.n594 B.n37 163.367
R716 B.n594 B.n593 163.367
R717 B.n593 B.n592 163.367
R718 B.n592 B.n39 163.367
R719 B.n588 B.n39 163.367
R720 B.n588 B.n587 163.367
R721 B.n587 B.n586 163.367
R722 B.n586 B.n41 163.367
R723 B.n582 B.n41 163.367
R724 B.n582 B.n581 163.367
R725 B.n581 B.n580 163.367
R726 B.n580 B.n43 163.367
R727 B.n576 B.n43 163.367
R728 B.n576 B.n575 163.367
R729 B.n575 B.n574 163.367
R730 B.n574 B.n48 163.367
R731 B.n570 B.n48 163.367
R732 B.n570 B.n569 163.367
R733 B.n569 B.n568 163.367
R734 B.n568 B.n50 163.367
R735 B.n563 B.n50 163.367
R736 B.n563 B.n562 163.367
R737 B.n562 B.n561 163.367
R738 B.n561 B.n54 163.367
R739 B.n557 B.n54 163.367
R740 B.n557 B.n556 163.367
R741 B.n556 B.n555 163.367
R742 B.n555 B.n56 163.367
R743 B.n551 B.n56 163.367
R744 B.n551 B.n550 163.367
R745 B.n550 B.n549 163.367
R746 B.n549 B.n58 163.367
R747 B.n545 B.n58 163.367
R748 B.n545 B.n544 163.367
R749 B.n544 B.n543 163.367
R750 B.n543 B.n60 163.367
R751 B.n539 B.n60 163.367
R752 B.n539 B.n538 163.367
R753 B.n538 B.n537 163.367
R754 B.n537 B.n62 163.367
R755 B.n533 B.n62 163.367
R756 B.n533 B.n532 163.367
R757 B.n532 B.n531 163.367
R758 B.n531 B.n64 163.367
R759 B.n527 B.n64 163.367
R760 B.n527 B.n526 163.367
R761 B.n526 B.n525 163.367
R762 B.n525 B.n66 163.367
R763 B.n521 B.n66 163.367
R764 B.n521 B.n520 163.367
R765 B.n520 B.n519 163.367
R766 B.n519 B.n68 163.367
R767 B.n515 B.n68 163.367
R768 B.n515 B.n514 163.367
R769 B.n514 B.n513 163.367
R770 B.n136 B.t10 112.615
R771 B.n52 B.t2 112.615
R772 B.n142 B.t4 112.603
R773 B.n45 B.t8 112.603
R774 B.n136 B.n135 83.7823
R775 B.n142 B.n141 83.7823
R776 B.n45 B.n44 83.7823
R777 B.n52 B.n51 83.7823
R778 B.n319 B.n136 59.5399
R779 B.n143 B.n142 59.5399
R780 B.n46 B.n45 59.5399
R781 B.n565 B.n52 59.5399
R782 B.n633 B.n632 33.2493
R783 B.n512 B.n511 33.2493
R784 B.n373 B.n372 33.2493
R785 B.n252 B.n161 33.2493
R786 B B.n703 18.0485
R787 B.n632 B.n631 10.6151
R788 B.n631 B.n26 10.6151
R789 B.n627 B.n26 10.6151
R790 B.n627 B.n626 10.6151
R791 B.n626 B.n625 10.6151
R792 B.n625 B.n28 10.6151
R793 B.n621 B.n28 10.6151
R794 B.n621 B.n620 10.6151
R795 B.n620 B.n619 10.6151
R796 B.n619 B.n30 10.6151
R797 B.n615 B.n30 10.6151
R798 B.n615 B.n614 10.6151
R799 B.n614 B.n613 10.6151
R800 B.n613 B.n32 10.6151
R801 B.n609 B.n32 10.6151
R802 B.n609 B.n608 10.6151
R803 B.n608 B.n607 10.6151
R804 B.n607 B.n34 10.6151
R805 B.n603 B.n34 10.6151
R806 B.n603 B.n602 10.6151
R807 B.n602 B.n601 10.6151
R808 B.n601 B.n36 10.6151
R809 B.n597 B.n36 10.6151
R810 B.n597 B.n596 10.6151
R811 B.n596 B.n595 10.6151
R812 B.n595 B.n38 10.6151
R813 B.n591 B.n38 10.6151
R814 B.n591 B.n590 10.6151
R815 B.n590 B.n589 10.6151
R816 B.n589 B.n40 10.6151
R817 B.n585 B.n40 10.6151
R818 B.n585 B.n584 10.6151
R819 B.n584 B.n583 10.6151
R820 B.n583 B.n42 10.6151
R821 B.n579 B.n578 10.6151
R822 B.n578 B.n577 10.6151
R823 B.n577 B.n47 10.6151
R824 B.n573 B.n47 10.6151
R825 B.n573 B.n572 10.6151
R826 B.n572 B.n571 10.6151
R827 B.n571 B.n49 10.6151
R828 B.n567 B.n49 10.6151
R829 B.n567 B.n566 10.6151
R830 B.n564 B.n53 10.6151
R831 B.n560 B.n53 10.6151
R832 B.n560 B.n559 10.6151
R833 B.n559 B.n558 10.6151
R834 B.n558 B.n55 10.6151
R835 B.n554 B.n55 10.6151
R836 B.n554 B.n553 10.6151
R837 B.n553 B.n552 10.6151
R838 B.n552 B.n57 10.6151
R839 B.n548 B.n57 10.6151
R840 B.n548 B.n547 10.6151
R841 B.n547 B.n546 10.6151
R842 B.n546 B.n59 10.6151
R843 B.n542 B.n59 10.6151
R844 B.n542 B.n541 10.6151
R845 B.n541 B.n540 10.6151
R846 B.n540 B.n61 10.6151
R847 B.n536 B.n61 10.6151
R848 B.n536 B.n535 10.6151
R849 B.n535 B.n534 10.6151
R850 B.n534 B.n63 10.6151
R851 B.n530 B.n63 10.6151
R852 B.n530 B.n529 10.6151
R853 B.n529 B.n528 10.6151
R854 B.n528 B.n65 10.6151
R855 B.n524 B.n65 10.6151
R856 B.n524 B.n523 10.6151
R857 B.n523 B.n522 10.6151
R858 B.n522 B.n67 10.6151
R859 B.n518 B.n67 10.6151
R860 B.n518 B.n517 10.6151
R861 B.n517 B.n516 10.6151
R862 B.n516 B.n69 10.6151
R863 B.n512 B.n69 10.6151
R864 B.n374 B.n373 10.6151
R865 B.n374 B.n115 10.6151
R866 B.n378 B.n115 10.6151
R867 B.n379 B.n378 10.6151
R868 B.n380 B.n379 10.6151
R869 B.n380 B.n113 10.6151
R870 B.n384 B.n113 10.6151
R871 B.n385 B.n384 10.6151
R872 B.n386 B.n385 10.6151
R873 B.n386 B.n111 10.6151
R874 B.n390 B.n111 10.6151
R875 B.n391 B.n390 10.6151
R876 B.n392 B.n391 10.6151
R877 B.n392 B.n109 10.6151
R878 B.n396 B.n109 10.6151
R879 B.n397 B.n396 10.6151
R880 B.n398 B.n397 10.6151
R881 B.n398 B.n107 10.6151
R882 B.n402 B.n107 10.6151
R883 B.n403 B.n402 10.6151
R884 B.n404 B.n403 10.6151
R885 B.n404 B.n105 10.6151
R886 B.n408 B.n105 10.6151
R887 B.n409 B.n408 10.6151
R888 B.n410 B.n409 10.6151
R889 B.n410 B.n103 10.6151
R890 B.n414 B.n103 10.6151
R891 B.n415 B.n414 10.6151
R892 B.n416 B.n415 10.6151
R893 B.n416 B.n101 10.6151
R894 B.n420 B.n101 10.6151
R895 B.n421 B.n420 10.6151
R896 B.n422 B.n421 10.6151
R897 B.n422 B.n99 10.6151
R898 B.n426 B.n99 10.6151
R899 B.n427 B.n426 10.6151
R900 B.n428 B.n427 10.6151
R901 B.n428 B.n97 10.6151
R902 B.n432 B.n97 10.6151
R903 B.n433 B.n432 10.6151
R904 B.n434 B.n433 10.6151
R905 B.n434 B.n95 10.6151
R906 B.n438 B.n95 10.6151
R907 B.n439 B.n438 10.6151
R908 B.n440 B.n439 10.6151
R909 B.n440 B.n93 10.6151
R910 B.n444 B.n93 10.6151
R911 B.n445 B.n444 10.6151
R912 B.n446 B.n445 10.6151
R913 B.n446 B.n91 10.6151
R914 B.n450 B.n91 10.6151
R915 B.n451 B.n450 10.6151
R916 B.n452 B.n451 10.6151
R917 B.n452 B.n89 10.6151
R918 B.n456 B.n89 10.6151
R919 B.n457 B.n456 10.6151
R920 B.n458 B.n457 10.6151
R921 B.n458 B.n87 10.6151
R922 B.n462 B.n87 10.6151
R923 B.n463 B.n462 10.6151
R924 B.n464 B.n463 10.6151
R925 B.n464 B.n85 10.6151
R926 B.n468 B.n85 10.6151
R927 B.n469 B.n468 10.6151
R928 B.n470 B.n469 10.6151
R929 B.n470 B.n83 10.6151
R930 B.n474 B.n83 10.6151
R931 B.n475 B.n474 10.6151
R932 B.n476 B.n475 10.6151
R933 B.n476 B.n81 10.6151
R934 B.n480 B.n81 10.6151
R935 B.n481 B.n480 10.6151
R936 B.n482 B.n481 10.6151
R937 B.n482 B.n79 10.6151
R938 B.n486 B.n79 10.6151
R939 B.n487 B.n486 10.6151
R940 B.n488 B.n487 10.6151
R941 B.n488 B.n77 10.6151
R942 B.n492 B.n77 10.6151
R943 B.n493 B.n492 10.6151
R944 B.n494 B.n493 10.6151
R945 B.n494 B.n75 10.6151
R946 B.n498 B.n75 10.6151
R947 B.n499 B.n498 10.6151
R948 B.n500 B.n499 10.6151
R949 B.n500 B.n73 10.6151
R950 B.n504 B.n73 10.6151
R951 B.n505 B.n504 10.6151
R952 B.n506 B.n505 10.6151
R953 B.n506 B.n71 10.6151
R954 B.n510 B.n71 10.6151
R955 B.n511 B.n510 10.6151
R956 B.n253 B.n252 10.6151
R957 B.n254 B.n253 10.6151
R958 B.n254 B.n159 10.6151
R959 B.n258 B.n159 10.6151
R960 B.n259 B.n258 10.6151
R961 B.n260 B.n259 10.6151
R962 B.n260 B.n157 10.6151
R963 B.n264 B.n157 10.6151
R964 B.n265 B.n264 10.6151
R965 B.n266 B.n265 10.6151
R966 B.n266 B.n155 10.6151
R967 B.n270 B.n155 10.6151
R968 B.n271 B.n270 10.6151
R969 B.n272 B.n271 10.6151
R970 B.n272 B.n153 10.6151
R971 B.n276 B.n153 10.6151
R972 B.n277 B.n276 10.6151
R973 B.n278 B.n277 10.6151
R974 B.n278 B.n151 10.6151
R975 B.n282 B.n151 10.6151
R976 B.n283 B.n282 10.6151
R977 B.n284 B.n283 10.6151
R978 B.n284 B.n149 10.6151
R979 B.n288 B.n149 10.6151
R980 B.n289 B.n288 10.6151
R981 B.n290 B.n289 10.6151
R982 B.n290 B.n147 10.6151
R983 B.n294 B.n147 10.6151
R984 B.n295 B.n294 10.6151
R985 B.n296 B.n295 10.6151
R986 B.n296 B.n145 10.6151
R987 B.n300 B.n145 10.6151
R988 B.n301 B.n300 10.6151
R989 B.n302 B.n301 10.6151
R990 B.n306 B.n305 10.6151
R991 B.n307 B.n306 10.6151
R992 B.n307 B.n139 10.6151
R993 B.n311 B.n139 10.6151
R994 B.n312 B.n311 10.6151
R995 B.n313 B.n312 10.6151
R996 B.n313 B.n137 10.6151
R997 B.n317 B.n137 10.6151
R998 B.n318 B.n317 10.6151
R999 B.n320 B.n133 10.6151
R1000 B.n324 B.n133 10.6151
R1001 B.n325 B.n324 10.6151
R1002 B.n326 B.n325 10.6151
R1003 B.n326 B.n131 10.6151
R1004 B.n330 B.n131 10.6151
R1005 B.n331 B.n330 10.6151
R1006 B.n332 B.n331 10.6151
R1007 B.n332 B.n129 10.6151
R1008 B.n336 B.n129 10.6151
R1009 B.n337 B.n336 10.6151
R1010 B.n338 B.n337 10.6151
R1011 B.n338 B.n127 10.6151
R1012 B.n342 B.n127 10.6151
R1013 B.n343 B.n342 10.6151
R1014 B.n344 B.n343 10.6151
R1015 B.n344 B.n125 10.6151
R1016 B.n348 B.n125 10.6151
R1017 B.n349 B.n348 10.6151
R1018 B.n350 B.n349 10.6151
R1019 B.n350 B.n123 10.6151
R1020 B.n354 B.n123 10.6151
R1021 B.n355 B.n354 10.6151
R1022 B.n356 B.n355 10.6151
R1023 B.n356 B.n121 10.6151
R1024 B.n360 B.n121 10.6151
R1025 B.n361 B.n360 10.6151
R1026 B.n362 B.n361 10.6151
R1027 B.n362 B.n119 10.6151
R1028 B.n366 B.n119 10.6151
R1029 B.n367 B.n366 10.6151
R1030 B.n368 B.n367 10.6151
R1031 B.n368 B.n117 10.6151
R1032 B.n372 B.n117 10.6151
R1033 B.n248 B.n161 10.6151
R1034 B.n248 B.n247 10.6151
R1035 B.n247 B.n246 10.6151
R1036 B.n246 B.n163 10.6151
R1037 B.n242 B.n163 10.6151
R1038 B.n242 B.n241 10.6151
R1039 B.n241 B.n240 10.6151
R1040 B.n240 B.n165 10.6151
R1041 B.n236 B.n165 10.6151
R1042 B.n236 B.n235 10.6151
R1043 B.n235 B.n234 10.6151
R1044 B.n234 B.n167 10.6151
R1045 B.n230 B.n167 10.6151
R1046 B.n230 B.n229 10.6151
R1047 B.n229 B.n228 10.6151
R1048 B.n228 B.n169 10.6151
R1049 B.n224 B.n169 10.6151
R1050 B.n224 B.n223 10.6151
R1051 B.n223 B.n222 10.6151
R1052 B.n222 B.n171 10.6151
R1053 B.n218 B.n171 10.6151
R1054 B.n218 B.n217 10.6151
R1055 B.n217 B.n216 10.6151
R1056 B.n216 B.n173 10.6151
R1057 B.n212 B.n173 10.6151
R1058 B.n212 B.n211 10.6151
R1059 B.n211 B.n210 10.6151
R1060 B.n210 B.n175 10.6151
R1061 B.n206 B.n175 10.6151
R1062 B.n206 B.n205 10.6151
R1063 B.n205 B.n204 10.6151
R1064 B.n204 B.n177 10.6151
R1065 B.n200 B.n177 10.6151
R1066 B.n200 B.n199 10.6151
R1067 B.n199 B.n198 10.6151
R1068 B.n198 B.n179 10.6151
R1069 B.n194 B.n179 10.6151
R1070 B.n194 B.n193 10.6151
R1071 B.n193 B.n192 10.6151
R1072 B.n192 B.n181 10.6151
R1073 B.n188 B.n181 10.6151
R1074 B.n188 B.n187 10.6151
R1075 B.n187 B.n186 10.6151
R1076 B.n186 B.n183 10.6151
R1077 B.n183 B.n0 10.6151
R1078 B.n699 B.n1 10.6151
R1079 B.n699 B.n698 10.6151
R1080 B.n698 B.n697 10.6151
R1081 B.n697 B.n4 10.6151
R1082 B.n693 B.n4 10.6151
R1083 B.n693 B.n692 10.6151
R1084 B.n692 B.n691 10.6151
R1085 B.n691 B.n6 10.6151
R1086 B.n687 B.n6 10.6151
R1087 B.n687 B.n686 10.6151
R1088 B.n686 B.n685 10.6151
R1089 B.n685 B.n8 10.6151
R1090 B.n681 B.n8 10.6151
R1091 B.n681 B.n680 10.6151
R1092 B.n680 B.n679 10.6151
R1093 B.n679 B.n10 10.6151
R1094 B.n675 B.n10 10.6151
R1095 B.n675 B.n674 10.6151
R1096 B.n674 B.n673 10.6151
R1097 B.n673 B.n12 10.6151
R1098 B.n669 B.n12 10.6151
R1099 B.n669 B.n668 10.6151
R1100 B.n668 B.n667 10.6151
R1101 B.n667 B.n14 10.6151
R1102 B.n663 B.n14 10.6151
R1103 B.n663 B.n662 10.6151
R1104 B.n662 B.n661 10.6151
R1105 B.n661 B.n16 10.6151
R1106 B.n657 B.n16 10.6151
R1107 B.n657 B.n656 10.6151
R1108 B.n656 B.n655 10.6151
R1109 B.n655 B.n18 10.6151
R1110 B.n651 B.n18 10.6151
R1111 B.n651 B.n650 10.6151
R1112 B.n650 B.n649 10.6151
R1113 B.n649 B.n20 10.6151
R1114 B.n645 B.n20 10.6151
R1115 B.n645 B.n644 10.6151
R1116 B.n644 B.n643 10.6151
R1117 B.n643 B.n22 10.6151
R1118 B.n639 B.n22 10.6151
R1119 B.n639 B.n638 10.6151
R1120 B.n638 B.n637 10.6151
R1121 B.n637 B.n24 10.6151
R1122 B.n633 B.n24 10.6151
R1123 B.n46 B.n42 9.36635
R1124 B.n565 B.n564 9.36635
R1125 B.n302 B.n143 9.36635
R1126 B.n320 B.n319 9.36635
R1127 B.n703 B.n0 2.81026
R1128 B.n703 B.n1 2.81026
R1129 B.n579 B.n46 1.24928
R1130 B.n566 B.n565 1.24928
R1131 B.n305 B.n143 1.24928
R1132 B.n319 B.n318 1.24928
C0 w_n3562_n2922# B 10.33f
C1 VP VDD2 0.482912f
C2 VTAIL B 4.71703f
C3 VDD1 VN 0.150415f
C4 VDD2 B 1.52338f
C5 w_n3562_n2922# VDD1 1.6546f
C6 VP B 2.11829f
C7 w_n3562_n2922# VN 6.25104f
C8 VTAIL VDD1 5.3641f
C9 VTAIL VN 4.40849f
C10 w_n3562_n2922# VTAIL 3.53672f
C11 VDD2 VDD1 1.36932f
C12 VDD2 VN 4.180201f
C13 VP VDD1 4.51161f
C14 VP VN 6.78235f
C15 w_n3562_n2922# VDD2 1.74134f
C16 VP w_n3562_n2922# 6.71247f
C17 VDD2 VTAIL 5.42762f
C18 VDD1 B 1.44824f
C19 VP VTAIL 4.4226f
C20 B VN 1.34611f
C21 VDD2 VSUBS 1.11668f
C22 VDD1 VSUBS 6.30904f
C23 VTAIL VSUBS 1.311107f
C24 VN VSUBS 6.24454f
C25 VP VSUBS 2.965695f
C26 B VSUBS 5.284239f
C27 w_n3562_n2922# VSUBS 0.128617p
C28 B.n0 VSUBS 0.004696f
C29 B.n1 VSUBS 0.004696f
C30 B.n2 VSUBS 0.007426f
C31 B.n3 VSUBS 0.007426f
C32 B.n4 VSUBS 0.007426f
C33 B.n5 VSUBS 0.007426f
C34 B.n6 VSUBS 0.007426f
C35 B.n7 VSUBS 0.007426f
C36 B.n8 VSUBS 0.007426f
C37 B.n9 VSUBS 0.007426f
C38 B.n10 VSUBS 0.007426f
C39 B.n11 VSUBS 0.007426f
C40 B.n12 VSUBS 0.007426f
C41 B.n13 VSUBS 0.007426f
C42 B.n14 VSUBS 0.007426f
C43 B.n15 VSUBS 0.007426f
C44 B.n16 VSUBS 0.007426f
C45 B.n17 VSUBS 0.007426f
C46 B.n18 VSUBS 0.007426f
C47 B.n19 VSUBS 0.007426f
C48 B.n20 VSUBS 0.007426f
C49 B.n21 VSUBS 0.007426f
C50 B.n22 VSUBS 0.007426f
C51 B.n23 VSUBS 0.007426f
C52 B.n24 VSUBS 0.007426f
C53 B.n25 VSUBS 0.018265f
C54 B.n26 VSUBS 0.007426f
C55 B.n27 VSUBS 0.007426f
C56 B.n28 VSUBS 0.007426f
C57 B.n29 VSUBS 0.007426f
C58 B.n30 VSUBS 0.007426f
C59 B.n31 VSUBS 0.007426f
C60 B.n32 VSUBS 0.007426f
C61 B.n33 VSUBS 0.007426f
C62 B.n34 VSUBS 0.007426f
C63 B.n35 VSUBS 0.007426f
C64 B.n36 VSUBS 0.007426f
C65 B.n37 VSUBS 0.007426f
C66 B.n38 VSUBS 0.007426f
C67 B.n39 VSUBS 0.007426f
C68 B.n40 VSUBS 0.007426f
C69 B.n41 VSUBS 0.007426f
C70 B.n42 VSUBS 0.006989f
C71 B.n43 VSUBS 0.007426f
C72 B.t8 VSUBS 0.3295f
C73 B.t7 VSUBS 0.360002f
C74 B.t6 VSUBS 1.95324f
C75 B.n44 VSUBS 0.208076f
C76 B.n45 VSUBS 0.082087f
C77 B.n46 VSUBS 0.017205f
C78 B.n47 VSUBS 0.007426f
C79 B.n48 VSUBS 0.007426f
C80 B.n49 VSUBS 0.007426f
C81 B.n50 VSUBS 0.007426f
C82 B.t2 VSUBS 0.329496f
C83 B.t1 VSUBS 0.359998f
C84 B.t0 VSUBS 1.95324f
C85 B.n51 VSUBS 0.208081f
C86 B.n52 VSUBS 0.082092f
C87 B.n53 VSUBS 0.007426f
C88 B.n54 VSUBS 0.007426f
C89 B.n55 VSUBS 0.007426f
C90 B.n56 VSUBS 0.007426f
C91 B.n57 VSUBS 0.007426f
C92 B.n58 VSUBS 0.007426f
C93 B.n59 VSUBS 0.007426f
C94 B.n60 VSUBS 0.007426f
C95 B.n61 VSUBS 0.007426f
C96 B.n62 VSUBS 0.007426f
C97 B.n63 VSUBS 0.007426f
C98 B.n64 VSUBS 0.007426f
C99 B.n65 VSUBS 0.007426f
C100 B.n66 VSUBS 0.007426f
C101 B.n67 VSUBS 0.007426f
C102 B.n68 VSUBS 0.007426f
C103 B.n69 VSUBS 0.007426f
C104 B.n70 VSUBS 0.016898f
C105 B.n71 VSUBS 0.007426f
C106 B.n72 VSUBS 0.007426f
C107 B.n73 VSUBS 0.007426f
C108 B.n74 VSUBS 0.007426f
C109 B.n75 VSUBS 0.007426f
C110 B.n76 VSUBS 0.007426f
C111 B.n77 VSUBS 0.007426f
C112 B.n78 VSUBS 0.007426f
C113 B.n79 VSUBS 0.007426f
C114 B.n80 VSUBS 0.007426f
C115 B.n81 VSUBS 0.007426f
C116 B.n82 VSUBS 0.007426f
C117 B.n83 VSUBS 0.007426f
C118 B.n84 VSUBS 0.007426f
C119 B.n85 VSUBS 0.007426f
C120 B.n86 VSUBS 0.007426f
C121 B.n87 VSUBS 0.007426f
C122 B.n88 VSUBS 0.007426f
C123 B.n89 VSUBS 0.007426f
C124 B.n90 VSUBS 0.007426f
C125 B.n91 VSUBS 0.007426f
C126 B.n92 VSUBS 0.007426f
C127 B.n93 VSUBS 0.007426f
C128 B.n94 VSUBS 0.007426f
C129 B.n95 VSUBS 0.007426f
C130 B.n96 VSUBS 0.007426f
C131 B.n97 VSUBS 0.007426f
C132 B.n98 VSUBS 0.007426f
C133 B.n99 VSUBS 0.007426f
C134 B.n100 VSUBS 0.007426f
C135 B.n101 VSUBS 0.007426f
C136 B.n102 VSUBS 0.007426f
C137 B.n103 VSUBS 0.007426f
C138 B.n104 VSUBS 0.007426f
C139 B.n105 VSUBS 0.007426f
C140 B.n106 VSUBS 0.007426f
C141 B.n107 VSUBS 0.007426f
C142 B.n108 VSUBS 0.007426f
C143 B.n109 VSUBS 0.007426f
C144 B.n110 VSUBS 0.007426f
C145 B.n111 VSUBS 0.007426f
C146 B.n112 VSUBS 0.007426f
C147 B.n113 VSUBS 0.007426f
C148 B.n114 VSUBS 0.007426f
C149 B.n115 VSUBS 0.007426f
C150 B.n116 VSUBS 0.016898f
C151 B.n117 VSUBS 0.007426f
C152 B.n118 VSUBS 0.007426f
C153 B.n119 VSUBS 0.007426f
C154 B.n120 VSUBS 0.007426f
C155 B.n121 VSUBS 0.007426f
C156 B.n122 VSUBS 0.007426f
C157 B.n123 VSUBS 0.007426f
C158 B.n124 VSUBS 0.007426f
C159 B.n125 VSUBS 0.007426f
C160 B.n126 VSUBS 0.007426f
C161 B.n127 VSUBS 0.007426f
C162 B.n128 VSUBS 0.007426f
C163 B.n129 VSUBS 0.007426f
C164 B.n130 VSUBS 0.007426f
C165 B.n131 VSUBS 0.007426f
C166 B.n132 VSUBS 0.007426f
C167 B.n133 VSUBS 0.007426f
C168 B.n134 VSUBS 0.007426f
C169 B.t10 VSUBS 0.329496f
C170 B.t11 VSUBS 0.359998f
C171 B.t9 VSUBS 1.95324f
C172 B.n135 VSUBS 0.208081f
C173 B.n136 VSUBS 0.082092f
C174 B.n137 VSUBS 0.007426f
C175 B.n138 VSUBS 0.007426f
C176 B.n139 VSUBS 0.007426f
C177 B.n140 VSUBS 0.007426f
C178 B.t4 VSUBS 0.3295f
C179 B.t5 VSUBS 0.360002f
C180 B.t3 VSUBS 1.95324f
C181 B.n141 VSUBS 0.208076f
C182 B.n142 VSUBS 0.082087f
C183 B.n143 VSUBS 0.017205f
C184 B.n144 VSUBS 0.007426f
C185 B.n145 VSUBS 0.007426f
C186 B.n146 VSUBS 0.007426f
C187 B.n147 VSUBS 0.007426f
C188 B.n148 VSUBS 0.007426f
C189 B.n149 VSUBS 0.007426f
C190 B.n150 VSUBS 0.007426f
C191 B.n151 VSUBS 0.007426f
C192 B.n152 VSUBS 0.007426f
C193 B.n153 VSUBS 0.007426f
C194 B.n154 VSUBS 0.007426f
C195 B.n155 VSUBS 0.007426f
C196 B.n156 VSUBS 0.007426f
C197 B.n157 VSUBS 0.007426f
C198 B.n158 VSUBS 0.007426f
C199 B.n159 VSUBS 0.007426f
C200 B.n160 VSUBS 0.007426f
C201 B.n161 VSUBS 0.016898f
C202 B.n162 VSUBS 0.007426f
C203 B.n163 VSUBS 0.007426f
C204 B.n164 VSUBS 0.007426f
C205 B.n165 VSUBS 0.007426f
C206 B.n166 VSUBS 0.007426f
C207 B.n167 VSUBS 0.007426f
C208 B.n168 VSUBS 0.007426f
C209 B.n169 VSUBS 0.007426f
C210 B.n170 VSUBS 0.007426f
C211 B.n171 VSUBS 0.007426f
C212 B.n172 VSUBS 0.007426f
C213 B.n173 VSUBS 0.007426f
C214 B.n174 VSUBS 0.007426f
C215 B.n175 VSUBS 0.007426f
C216 B.n176 VSUBS 0.007426f
C217 B.n177 VSUBS 0.007426f
C218 B.n178 VSUBS 0.007426f
C219 B.n179 VSUBS 0.007426f
C220 B.n180 VSUBS 0.007426f
C221 B.n181 VSUBS 0.007426f
C222 B.n182 VSUBS 0.007426f
C223 B.n183 VSUBS 0.007426f
C224 B.n184 VSUBS 0.007426f
C225 B.n185 VSUBS 0.007426f
C226 B.n186 VSUBS 0.007426f
C227 B.n187 VSUBS 0.007426f
C228 B.n188 VSUBS 0.007426f
C229 B.n189 VSUBS 0.007426f
C230 B.n190 VSUBS 0.007426f
C231 B.n191 VSUBS 0.007426f
C232 B.n192 VSUBS 0.007426f
C233 B.n193 VSUBS 0.007426f
C234 B.n194 VSUBS 0.007426f
C235 B.n195 VSUBS 0.007426f
C236 B.n196 VSUBS 0.007426f
C237 B.n197 VSUBS 0.007426f
C238 B.n198 VSUBS 0.007426f
C239 B.n199 VSUBS 0.007426f
C240 B.n200 VSUBS 0.007426f
C241 B.n201 VSUBS 0.007426f
C242 B.n202 VSUBS 0.007426f
C243 B.n203 VSUBS 0.007426f
C244 B.n204 VSUBS 0.007426f
C245 B.n205 VSUBS 0.007426f
C246 B.n206 VSUBS 0.007426f
C247 B.n207 VSUBS 0.007426f
C248 B.n208 VSUBS 0.007426f
C249 B.n209 VSUBS 0.007426f
C250 B.n210 VSUBS 0.007426f
C251 B.n211 VSUBS 0.007426f
C252 B.n212 VSUBS 0.007426f
C253 B.n213 VSUBS 0.007426f
C254 B.n214 VSUBS 0.007426f
C255 B.n215 VSUBS 0.007426f
C256 B.n216 VSUBS 0.007426f
C257 B.n217 VSUBS 0.007426f
C258 B.n218 VSUBS 0.007426f
C259 B.n219 VSUBS 0.007426f
C260 B.n220 VSUBS 0.007426f
C261 B.n221 VSUBS 0.007426f
C262 B.n222 VSUBS 0.007426f
C263 B.n223 VSUBS 0.007426f
C264 B.n224 VSUBS 0.007426f
C265 B.n225 VSUBS 0.007426f
C266 B.n226 VSUBS 0.007426f
C267 B.n227 VSUBS 0.007426f
C268 B.n228 VSUBS 0.007426f
C269 B.n229 VSUBS 0.007426f
C270 B.n230 VSUBS 0.007426f
C271 B.n231 VSUBS 0.007426f
C272 B.n232 VSUBS 0.007426f
C273 B.n233 VSUBS 0.007426f
C274 B.n234 VSUBS 0.007426f
C275 B.n235 VSUBS 0.007426f
C276 B.n236 VSUBS 0.007426f
C277 B.n237 VSUBS 0.007426f
C278 B.n238 VSUBS 0.007426f
C279 B.n239 VSUBS 0.007426f
C280 B.n240 VSUBS 0.007426f
C281 B.n241 VSUBS 0.007426f
C282 B.n242 VSUBS 0.007426f
C283 B.n243 VSUBS 0.007426f
C284 B.n244 VSUBS 0.007426f
C285 B.n245 VSUBS 0.007426f
C286 B.n246 VSUBS 0.007426f
C287 B.n247 VSUBS 0.007426f
C288 B.n248 VSUBS 0.007426f
C289 B.n249 VSUBS 0.007426f
C290 B.n250 VSUBS 0.016898f
C291 B.n251 VSUBS 0.018265f
C292 B.n252 VSUBS 0.018265f
C293 B.n253 VSUBS 0.007426f
C294 B.n254 VSUBS 0.007426f
C295 B.n255 VSUBS 0.007426f
C296 B.n256 VSUBS 0.007426f
C297 B.n257 VSUBS 0.007426f
C298 B.n258 VSUBS 0.007426f
C299 B.n259 VSUBS 0.007426f
C300 B.n260 VSUBS 0.007426f
C301 B.n261 VSUBS 0.007426f
C302 B.n262 VSUBS 0.007426f
C303 B.n263 VSUBS 0.007426f
C304 B.n264 VSUBS 0.007426f
C305 B.n265 VSUBS 0.007426f
C306 B.n266 VSUBS 0.007426f
C307 B.n267 VSUBS 0.007426f
C308 B.n268 VSUBS 0.007426f
C309 B.n269 VSUBS 0.007426f
C310 B.n270 VSUBS 0.007426f
C311 B.n271 VSUBS 0.007426f
C312 B.n272 VSUBS 0.007426f
C313 B.n273 VSUBS 0.007426f
C314 B.n274 VSUBS 0.007426f
C315 B.n275 VSUBS 0.007426f
C316 B.n276 VSUBS 0.007426f
C317 B.n277 VSUBS 0.007426f
C318 B.n278 VSUBS 0.007426f
C319 B.n279 VSUBS 0.007426f
C320 B.n280 VSUBS 0.007426f
C321 B.n281 VSUBS 0.007426f
C322 B.n282 VSUBS 0.007426f
C323 B.n283 VSUBS 0.007426f
C324 B.n284 VSUBS 0.007426f
C325 B.n285 VSUBS 0.007426f
C326 B.n286 VSUBS 0.007426f
C327 B.n287 VSUBS 0.007426f
C328 B.n288 VSUBS 0.007426f
C329 B.n289 VSUBS 0.007426f
C330 B.n290 VSUBS 0.007426f
C331 B.n291 VSUBS 0.007426f
C332 B.n292 VSUBS 0.007426f
C333 B.n293 VSUBS 0.007426f
C334 B.n294 VSUBS 0.007426f
C335 B.n295 VSUBS 0.007426f
C336 B.n296 VSUBS 0.007426f
C337 B.n297 VSUBS 0.007426f
C338 B.n298 VSUBS 0.007426f
C339 B.n299 VSUBS 0.007426f
C340 B.n300 VSUBS 0.007426f
C341 B.n301 VSUBS 0.007426f
C342 B.n302 VSUBS 0.006989f
C343 B.n303 VSUBS 0.007426f
C344 B.n304 VSUBS 0.007426f
C345 B.n305 VSUBS 0.00415f
C346 B.n306 VSUBS 0.007426f
C347 B.n307 VSUBS 0.007426f
C348 B.n308 VSUBS 0.007426f
C349 B.n309 VSUBS 0.007426f
C350 B.n310 VSUBS 0.007426f
C351 B.n311 VSUBS 0.007426f
C352 B.n312 VSUBS 0.007426f
C353 B.n313 VSUBS 0.007426f
C354 B.n314 VSUBS 0.007426f
C355 B.n315 VSUBS 0.007426f
C356 B.n316 VSUBS 0.007426f
C357 B.n317 VSUBS 0.007426f
C358 B.n318 VSUBS 0.00415f
C359 B.n319 VSUBS 0.017205f
C360 B.n320 VSUBS 0.006989f
C361 B.n321 VSUBS 0.007426f
C362 B.n322 VSUBS 0.007426f
C363 B.n323 VSUBS 0.007426f
C364 B.n324 VSUBS 0.007426f
C365 B.n325 VSUBS 0.007426f
C366 B.n326 VSUBS 0.007426f
C367 B.n327 VSUBS 0.007426f
C368 B.n328 VSUBS 0.007426f
C369 B.n329 VSUBS 0.007426f
C370 B.n330 VSUBS 0.007426f
C371 B.n331 VSUBS 0.007426f
C372 B.n332 VSUBS 0.007426f
C373 B.n333 VSUBS 0.007426f
C374 B.n334 VSUBS 0.007426f
C375 B.n335 VSUBS 0.007426f
C376 B.n336 VSUBS 0.007426f
C377 B.n337 VSUBS 0.007426f
C378 B.n338 VSUBS 0.007426f
C379 B.n339 VSUBS 0.007426f
C380 B.n340 VSUBS 0.007426f
C381 B.n341 VSUBS 0.007426f
C382 B.n342 VSUBS 0.007426f
C383 B.n343 VSUBS 0.007426f
C384 B.n344 VSUBS 0.007426f
C385 B.n345 VSUBS 0.007426f
C386 B.n346 VSUBS 0.007426f
C387 B.n347 VSUBS 0.007426f
C388 B.n348 VSUBS 0.007426f
C389 B.n349 VSUBS 0.007426f
C390 B.n350 VSUBS 0.007426f
C391 B.n351 VSUBS 0.007426f
C392 B.n352 VSUBS 0.007426f
C393 B.n353 VSUBS 0.007426f
C394 B.n354 VSUBS 0.007426f
C395 B.n355 VSUBS 0.007426f
C396 B.n356 VSUBS 0.007426f
C397 B.n357 VSUBS 0.007426f
C398 B.n358 VSUBS 0.007426f
C399 B.n359 VSUBS 0.007426f
C400 B.n360 VSUBS 0.007426f
C401 B.n361 VSUBS 0.007426f
C402 B.n362 VSUBS 0.007426f
C403 B.n363 VSUBS 0.007426f
C404 B.n364 VSUBS 0.007426f
C405 B.n365 VSUBS 0.007426f
C406 B.n366 VSUBS 0.007426f
C407 B.n367 VSUBS 0.007426f
C408 B.n368 VSUBS 0.007426f
C409 B.n369 VSUBS 0.007426f
C410 B.n370 VSUBS 0.007426f
C411 B.n371 VSUBS 0.018265f
C412 B.n372 VSUBS 0.018265f
C413 B.n373 VSUBS 0.016898f
C414 B.n374 VSUBS 0.007426f
C415 B.n375 VSUBS 0.007426f
C416 B.n376 VSUBS 0.007426f
C417 B.n377 VSUBS 0.007426f
C418 B.n378 VSUBS 0.007426f
C419 B.n379 VSUBS 0.007426f
C420 B.n380 VSUBS 0.007426f
C421 B.n381 VSUBS 0.007426f
C422 B.n382 VSUBS 0.007426f
C423 B.n383 VSUBS 0.007426f
C424 B.n384 VSUBS 0.007426f
C425 B.n385 VSUBS 0.007426f
C426 B.n386 VSUBS 0.007426f
C427 B.n387 VSUBS 0.007426f
C428 B.n388 VSUBS 0.007426f
C429 B.n389 VSUBS 0.007426f
C430 B.n390 VSUBS 0.007426f
C431 B.n391 VSUBS 0.007426f
C432 B.n392 VSUBS 0.007426f
C433 B.n393 VSUBS 0.007426f
C434 B.n394 VSUBS 0.007426f
C435 B.n395 VSUBS 0.007426f
C436 B.n396 VSUBS 0.007426f
C437 B.n397 VSUBS 0.007426f
C438 B.n398 VSUBS 0.007426f
C439 B.n399 VSUBS 0.007426f
C440 B.n400 VSUBS 0.007426f
C441 B.n401 VSUBS 0.007426f
C442 B.n402 VSUBS 0.007426f
C443 B.n403 VSUBS 0.007426f
C444 B.n404 VSUBS 0.007426f
C445 B.n405 VSUBS 0.007426f
C446 B.n406 VSUBS 0.007426f
C447 B.n407 VSUBS 0.007426f
C448 B.n408 VSUBS 0.007426f
C449 B.n409 VSUBS 0.007426f
C450 B.n410 VSUBS 0.007426f
C451 B.n411 VSUBS 0.007426f
C452 B.n412 VSUBS 0.007426f
C453 B.n413 VSUBS 0.007426f
C454 B.n414 VSUBS 0.007426f
C455 B.n415 VSUBS 0.007426f
C456 B.n416 VSUBS 0.007426f
C457 B.n417 VSUBS 0.007426f
C458 B.n418 VSUBS 0.007426f
C459 B.n419 VSUBS 0.007426f
C460 B.n420 VSUBS 0.007426f
C461 B.n421 VSUBS 0.007426f
C462 B.n422 VSUBS 0.007426f
C463 B.n423 VSUBS 0.007426f
C464 B.n424 VSUBS 0.007426f
C465 B.n425 VSUBS 0.007426f
C466 B.n426 VSUBS 0.007426f
C467 B.n427 VSUBS 0.007426f
C468 B.n428 VSUBS 0.007426f
C469 B.n429 VSUBS 0.007426f
C470 B.n430 VSUBS 0.007426f
C471 B.n431 VSUBS 0.007426f
C472 B.n432 VSUBS 0.007426f
C473 B.n433 VSUBS 0.007426f
C474 B.n434 VSUBS 0.007426f
C475 B.n435 VSUBS 0.007426f
C476 B.n436 VSUBS 0.007426f
C477 B.n437 VSUBS 0.007426f
C478 B.n438 VSUBS 0.007426f
C479 B.n439 VSUBS 0.007426f
C480 B.n440 VSUBS 0.007426f
C481 B.n441 VSUBS 0.007426f
C482 B.n442 VSUBS 0.007426f
C483 B.n443 VSUBS 0.007426f
C484 B.n444 VSUBS 0.007426f
C485 B.n445 VSUBS 0.007426f
C486 B.n446 VSUBS 0.007426f
C487 B.n447 VSUBS 0.007426f
C488 B.n448 VSUBS 0.007426f
C489 B.n449 VSUBS 0.007426f
C490 B.n450 VSUBS 0.007426f
C491 B.n451 VSUBS 0.007426f
C492 B.n452 VSUBS 0.007426f
C493 B.n453 VSUBS 0.007426f
C494 B.n454 VSUBS 0.007426f
C495 B.n455 VSUBS 0.007426f
C496 B.n456 VSUBS 0.007426f
C497 B.n457 VSUBS 0.007426f
C498 B.n458 VSUBS 0.007426f
C499 B.n459 VSUBS 0.007426f
C500 B.n460 VSUBS 0.007426f
C501 B.n461 VSUBS 0.007426f
C502 B.n462 VSUBS 0.007426f
C503 B.n463 VSUBS 0.007426f
C504 B.n464 VSUBS 0.007426f
C505 B.n465 VSUBS 0.007426f
C506 B.n466 VSUBS 0.007426f
C507 B.n467 VSUBS 0.007426f
C508 B.n468 VSUBS 0.007426f
C509 B.n469 VSUBS 0.007426f
C510 B.n470 VSUBS 0.007426f
C511 B.n471 VSUBS 0.007426f
C512 B.n472 VSUBS 0.007426f
C513 B.n473 VSUBS 0.007426f
C514 B.n474 VSUBS 0.007426f
C515 B.n475 VSUBS 0.007426f
C516 B.n476 VSUBS 0.007426f
C517 B.n477 VSUBS 0.007426f
C518 B.n478 VSUBS 0.007426f
C519 B.n479 VSUBS 0.007426f
C520 B.n480 VSUBS 0.007426f
C521 B.n481 VSUBS 0.007426f
C522 B.n482 VSUBS 0.007426f
C523 B.n483 VSUBS 0.007426f
C524 B.n484 VSUBS 0.007426f
C525 B.n485 VSUBS 0.007426f
C526 B.n486 VSUBS 0.007426f
C527 B.n487 VSUBS 0.007426f
C528 B.n488 VSUBS 0.007426f
C529 B.n489 VSUBS 0.007426f
C530 B.n490 VSUBS 0.007426f
C531 B.n491 VSUBS 0.007426f
C532 B.n492 VSUBS 0.007426f
C533 B.n493 VSUBS 0.007426f
C534 B.n494 VSUBS 0.007426f
C535 B.n495 VSUBS 0.007426f
C536 B.n496 VSUBS 0.007426f
C537 B.n497 VSUBS 0.007426f
C538 B.n498 VSUBS 0.007426f
C539 B.n499 VSUBS 0.007426f
C540 B.n500 VSUBS 0.007426f
C541 B.n501 VSUBS 0.007426f
C542 B.n502 VSUBS 0.007426f
C543 B.n503 VSUBS 0.007426f
C544 B.n504 VSUBS 0.007426f
C545 B.n505 VSUBS 0.007426f
C546 B.n506 VSUBS 0.007426f
C547 B.n507 VSUBS 0.007426f
C548 B.n508 VSUBS 0.007426f
C549 B.n509 VSUBS 0.007426f
C550 B.n510 VSUBS 0.007426f
C551 B.n511 VSUBS 0.01776f
C552 B.n512 VSUBS 0.017403f
C553 B.n513 VSUBS 0.018265f
C554 B.n514 VSUBS 0.007426f
C555 B.n515 VSUBS 0.007426f
C556 B.n516 VSUBS 0.007426f
C557 B.n517 VSUBS 0.007426f
C558 B.n518 VSUBS 0.007426f
C559 B.n519 VSUBS 0.007426f
C560 B.n520 VSUBS 0.007426f
C561 B.n521 VSUBS 0.007426f
C562 B.n522 VSUBS 0.007426f
C563 B.n523 VSUBS 0.007426f
C564 B.n524 VSUBS 0.007426f
C565 B.n525 VSUBS 0.007426f
C566 B.n526 VSUBS 0.007426f
C567 B.n527 VSUBS 0.007426f
C568 B.n528 VSUBS 0.007426f
C569 B.n529 VSUBS 0.007426f
C570 B.n530 VSUBS 0.007426f
C571 B.n531 VSUBS 0.007426f
C572 B.n532 VSUBS 0.007426f
C573 B.n533 VSUBS 0.007426f
C574 B.n534 VSUBS 0.007426f
C575 B.n535 VSUBS 0.007426f
C576 B.n536 VSUBS 0.007426f
C577 B.n537 VSUBS 0.007426f
C578 B.n538 VSUBS 0.007426f
C579 B.n539 VSUBS 0.007426f
C580 B.n540 VSUBS 0.007426f
C581 B.n541 VSUBS 0.007426f
C582 B.n542 VSUBS 0.007426f
C583 B.n543 VSUBS 0.007426f
C584 B.n544 VSUBS 0.007426f
C585 B.n545 VSUBS 0.007426f
C586 B.n546 VSUBS 0.007426f
C587 B.n547 VSUBS 0.007426f
C588 B.n548 VSUBS 0.007426f
C589 B.n549 VSUBS 0.007426f
C590 B.n550 VSUBS 0.007426f
C591 B.n551 VSUBS 0.007426f
C592 B.n552 VSUBS 0.007426f
C593 B.n553 VSUBS 0.007426f
C594 B.n554 VSUBS 0.007426f
C595 B.n555 VSUBS 0.007426f
C596 B.n556 VSUBS 0.007426f
C597 B.n557 VSUBS 0.007426f
C598 B.n558 VSUBS 0.007426f
C599 B.n559 VSUBS 0.007426f
C600 B.n560 VSUBS 0.007426f
C601 B.n561 VSUBS 0.007426f
C602 B.n562 VSUBS 0.007426f
C603 B.n563 VSUBS 0.007426f
C604 B.n564 VSUBS 0.006989f
C605 B.n565 VSUBS 0.017205f
C606 B.n566 VSUBS 0.00415f
C607 B.n567 VSUBS 0.007426f
C608 B.n568 VSUBS 0.007426f
C609 B.n569 VSUBS 0.007426f
C610 B.n570 VSUBS 0.007426f
C611 B.n571 VSUBS 0.007426f
C612 B.n572 VSUBS 0.007426f
C613 B.n573 VSUBS 0.007426f
C614 B.n574 VSUBS 0.007426f
C615 B.n575 VSUBS 0.007426f
C616 B.n576 VSUBS 0.007426f
C617 B.n577 VSUBS 0.007426f
C618 B.n578 VSUBS 0.007426f
C619 B.n579 VSUBS 0.00415f
C620 B.n580 VSUBS 0.007426f
C621 B.n581 VSUBS 0.007426f
C622 B.n582 VSUBS 0.007426f
C623 B.n583 VSUBS 0.007426f
C624 B.n584 VSUBS 0.007426f
C625 B.n585 VSUBS 0.007426f
C626 B.n586 VSUBS 0.007426f
C627 B.n587 VSUBS 0.007426f
C628 B.n588 VSUBS 0.007426f
C629 B.n589 VSUBS 0.007426f
C630 B.n590 VSUBS 0.007426f
C631 B.n591 VSUBS 0.007426f
C632 B.n592 VSUBS 0.007426f
C633 B.n593 VSUBS 0.007426f
C634 B.n594 VSUBS 0.007426f
C635 B.n595 VSUBS 0.007426f
C636 B.n596 VSUBS 0.007426f
C637 B.n597 VSUBS 0.007426f
C638 B.n598 VSUBS 0.007426f
C639 B.n599 VSUBS 0.007426f
C640 B.n600 VSUBS 0.007426f
C641 B.n601 VSUBS 0.007426f
C642 B.n602 VSUBS 0.007426f
C643 B.n603 VSUBS 0.007426f
C644 B.n604 VSUBS 0.007426f
C645 B.n605 VSUBS 0.007426f
C646 B.n606 VSUBS 0.007426f
C647 B.n607 VSUBS 0.007426f
C648 B.n608 VSUBS 0.007426f
C649 B.n609 VSUBS 0.007426f
C650 B.n610 VSUBS 0.007426f
C651 B.n611 VSUBS 0.007426f
C652 B.n612 VSUBS 0.007426f
C653 B.n613 VSUBS 0.007426f
C654 B.n614 VSUBS 0.007426f
C655 B.n615 VSUBS 0.007426f
C656 B.n616 VSUBS 0.007426f
C657 B.n617 VSUBS 0.007426f
C658 B.n618 VSUBS 0.007426f
C659 B.n619 VSUBS 0.007426f
C660 B.n620 VSUBS 0.007426f
C661 B.n621 VSUBS 0.007426f
C662 B.n622 VSUBS 0.007426f
C663 B.n623 VSUBS 0.007426f
C664 B.n624 VSUBS 0.007426f
C665 B.n625 VSUBS 0.007426f
C666 B.n626 VSUBS 0.007426f
C667 B.n627 VSUBS 0.007426f
C668 B.n628 VSUBS 0.007426f
C669 B.n629 VSUBS 0.007426f
C670 B.n630 VSUBS 0.007426f
C671 B.n631 VSUBS 0.007426f
C672 B.n632 VSUBS 0.018265f
C673 B.n633 VSUBS 0.016898f
C674 B.n634 VSUBS 0.016898f
C675 B.n635 VSUBS 0.007426f
C676 B.n636 VSUBS 0.007426f
C677 B.n637 VSUBS 0.007426f
C678 B.n638 VSUBS 0.007426f
C679 B.n639 VSUBS 0.007426f
C680 B.n640 VSUBS 0.007426f
C681 B.n641 VSUBS 0.007426f
C682 B.n642 VSUBS 0.007426f
C683 B.n643 VSUBS 0.007426f
C684 B.n644 VSUBS 0.007426f
C685 B.n645 VSUBS 0.007426f
C686 B.n646 VSUBS 0.007426f
C687 B.n647 VSUBS 0.007426f
C688 B.n648 VSUBS 0.007426f
C689 B.n649 VSUBS 0.007426f
C690 B.n650 VSUBS 0.007426f
C691 B.n651 VSUBS 0.007426f
C692 B.n652 VSUBS 0.007426f
C693 B.n653 VSUBS 0.007426f
C694 B.n654 VSUBS 0.007426f
C695 B.n655 VSUBS 0.007426f
C696 B.n656 VSUBS 0.007426f
C697 B.n657 VSUBS 0.007426f
C698 B.n658 VSUBS 0.007426f
C699 B.n659 VSUBS 0.007426f
C700 B.n660 VSUBS 0.007426f
C701 B.n661 VSUBS 0.007426f
C702 B.n662 VSUBS 0.007426f
C703 B.n663 VSUBS 0.007426f
C704 B.n664 VSUBS 0.007426f
C705 B.n665 VSUBS 0.007426f
C706 B.n666 VSUBS 0.007426f
C707 B.n667 VSUBS 0.007426f
C708 B.n668 VSUBS 0.007426f
C709 B.n669 VSUBS 0.007426f
C710 B.n670 VSUBS 0.007426f
C711 B.n671 VSUBS 0.007426f
C712 B.n672 VSUBS 0.007426f
C713 B.n673 VSUBS 0.007426f
C714 B.n674 VSUBS 0.007426f
C715 B.n675 VSUBS 0.007426f
C716 B.n676 VSUBS 0.007426f
C717 B.n677 VSUBS 0.007426f
C718 B.n678 VSUBS 0.007426f
C719 B.n679 VSUBS 0.007426f
C720 B.n680 VSUBS 0.007426f
C721 B.n681 VSUBS 0.007426f
C722 B.n682 VSUBS 0.007426f
C723 B.n683 VSUBS 0.007426f
C724 B.n684 VSUBS 0.007426f
C725 B.n685 VSUBS 0.007426f
C726 B.n686 VSUBS 0.007426f
C727 B.n687 VSUBS 0.007426f
C728 B.n688 VSUBS 0.007426f
C729 B.n689 VSUBS 0.007426f
C730 B.n690 VSUBS 0.007426f
C731 B.n691 VSUBS 0.007426f
C732 B.n692 VSUBS 0.007426f
C733 B.n693 VSUBS 0.007426f
C734 B.n694 VSUBS 0.007426f
C735 B.n695 VSUBS 0.007426f
C736 B.n696 VSUBS 0.007426f
C737 B.n697 VSUBS 0.007426f
C738 B.n698 VSUBS 0.007426f
C739 B.n699 VSUBS 0.007426f
C740 B.n700 VSUBS 0.007426f
C741 B.n701 VSUBS 0.007426f
C742 B.n702 VSUBS 0.007426f
C743 B.n703 VSUBS 0.016814f
C744 VDD2.t1 VSUBS 0.213699f
C745 VDD2.t3 VSUBS 0.213699f
C746 VDD2.n0 VSUBS 2.28667f
C747 VDD2.t0 VSUBS 0.213699f
C748 VDD2.t2 VSUBS 0.213699f
C749 VDD2.n1 VSUBS 1.6161f
C750 VDD2.n2 VSUBS 4.50433f
C751 VN.t2 VSUBS 3.46487f
C752 VN.t0 VSUBS 3.4456f
C753 VN.n0 VSUBS 2.039f
C754 VN.t1 VSUBS 3.46487f
C755 VN.t3 VSUBS 3.4456f
C756 VN.n1 VSUBS 3.86472f
C757 VDD1.t1 VSUBS 0.218055f
C758 VDD1.t2 VSUBS 0.218055f
C759 VDD1.n0 VSUBS 1.64965f
C760 VDD1.t0 VSUBS 0.218055f
C761 VDD1.t3 VSUBS 0.218055f
C762 VDD1.n1 VSUBS 2.35821f
C763 VTAIL.t0 VSUBS 1.84629f
C764 VTAIL.n0 VSUBS 0.81895f
C765 VTAIL.t7 VSUBS 1.84629f
C766 VTAIL.n1 VSUBS 0.968766f
C767 VTAIL.t6 VSUBS 1.84629f
C768 VTAIL.n2 VSUBS 2.28866f
C769 VTAIL.t2 VSUBS 1.8463f
C770 VTAIL.n3 VSUBS 2.28865f
C771 VTAIL.t1 VSUBS 1.8463f
C772 VTAIL.n4 VSUBS 0.968753f
C773 VTAIL.t4 VSUBS 1.8463f
C774 VTAIL.n5 VSUBS 0.968753f
C775 VTAIL.t5 VSUBS 1.84629f
C776 VTAIL.n6 VSUBS 2.28866f
C777 VTAIL.t3 VSUBS 1.84629f
C778 VTAIL.n7 VSUBS 2.12918f
C779 VP.n0 VSUBS 0.060343f
C780 VP.t0 VSUBS 3.38507f
C781 VP.n1 VSUBS 0.059789f
C782 VP.n2 VSUBS 0.03208f
C783 VP.n3 VSUBS 0.059789f
C784 VP.t1 VSUBS 3.89736f
C785 VP.t2 VSUBS 3.91915f
C786 VP.n4 VSUBS 4.36314f
C787 VP.n5 VSUBS 1.91959f
C788 VP.t3 VSUBS 3.38507f
C789 VP.n6 VSUBS 1.33852f
C790 VP.n7 VSUBS 0.054476f
C791 VP.n8 VSUBS 0.060343f
C792 VP.n9 VSUBS 0.03208f
C793 VP.n10 VSUBS 0.03208f
C794 VP.n11 VSUBS 0.059789f
C795 VP.n12 VSUBS 0.046831f
C796 VP.n13 VSUBS 0.046831f
C797 VP.n14 VSUBS 0.03208f
C798 VP.n15 VSUBS 0.03208f
C799 VP.n16 VSUBS 0.03208f
C800 VP.n17 VSUBS 0.059789f
C801 VP.n18 VSUBS 0.054476f
C802 VP.n19 VSUBS 1.33852f
C803 VP.n20 VSUBS 0.102816f
.ends

